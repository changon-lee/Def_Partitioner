module aes_aes_die_0 ( clk, key, ld, rst, text_in, done, text_out, N100, N102, 
       N105, N114, N116, N132, N133, N134, N147, N148, N149, 
       N150, N169, N227, N228, N229, N230, N231, N233, N242, 
       N244, N245, N246, N247, N258, N261, N277, N278, N280, 
       N35, N36, N37, N38, N40, N41, N430, N434, N435, 
       N436, N437, N438, N439, N440, N441, N463, N52, N53, 
       N54, N57, N66, N67, N68, N73, N82, N83, N84, 
       N85, N86, N87, N88, N89, N98, N99, n1145, n1183, 
       n1212, n1213, n1214, n1215, n1216, n1217, n1219, n1220, n1221, 
       n342, n348, n354, n362, n394, n396, n414, n419, n433, 
       n462, n469, n481, n482, n500, n506, n515, n524, n534, 
       n547, n562, n590, n636, n657, n665, n786, n791, n817, 
       n823, n830, n861, n870, n900, n905, n911, n917, n923, 
       n927, n937, n957, sa00_sr_0, sa00_sr_1, sa00_sr_2, sa00_sr_3, sa00_sr_4, sa00_sr_5, 
       sa00_sr_6, sa00_sr_7, sa01_sr_0, sa01_sr_1, sa01_sr_2, sa01_sr_3, sa01_sr_4, sa01_sr_5, sa01_sr_6, 
       sa01_sr_7, sa02_sr_0, sa02_sr_1, sa02_sr_2, sa02_sr_3, sa02_sr_4, sa02_sr_5, sa02_sr_6, sa02_sr_7, 
       sa03_sr_0, sa03_sr_1, sa03_sr_2, sa03_sr_3, sa03_sr_4, sa03_sr_5, sa03_sr_6, sa03_sr_7, sa10_sr_0, 
       sa10_sr_1, sa10_sr_2, sa10_sr_3, sa10_sr_4, sa10_sr_5, sa10_sr_6, sa10_sr_7, sa11_sr_0, sa11_sr_1, 
       sa11_sr_2, sa11_sr_3, sa11_sr_4, sa11_sr_5, sa11_sr_6, sa11_sr_7, sa12_sr_0, sa12_sr_1, sa12_sr_2, 
       sa12_sr_4, sa12_sr_5, sa12_sr_6, sa12_sr_7, sa20_sr_0, sa20_sr_1, sa20_sr_2, sa20_sr_3, sa20_sr_4, 
       sa20_sr_5, sa20_sr_6, sa20_sr_7, sa21_sr_0, sa21_sr_1, sa21_sr_2, sa21_sr_3, sa21_sr_4, sa21_sr_5, 
       sa21_sr_6, sa21_sr_7, sa22_sr_0, sa22_sr_1, sa22_sr_3, sa22_sr_4, sa22_sr_5, sa22_sr_6, sa22_sr_7, 
       sa23_sr_0, sa23_sr_1, sa23_sr_2, sa23_sr_3, sa23_sr_4, sa23_sr_5, sa23_sr_6, sa23_sr_7, sa30_sr_0, 
       sa30_sr_1, sa30_sr_2, sa30_sr_3, sa30_sr_4, sa30_sr_5, sa30_sr_6, sa30_sr_7, sa31_sr_0, sa31_sr_1, 
       sa31_sr_2, sa31_sr_3, sa31_sr_4, sa31_sr_5, sa31_sr_6, sa31_sr_7, sa32_sr_0, sa32_sr_1, sa32_sr_2, 
       sa32_sr_3, sa32_sr_4, sa32_sr_5, sa32_sr_6, sa32_sr_7, sa33_sr_0, sa33_sr_1, sa33_sr_2, sa33_sr_3, 
       sa33_sr_4, sa33_sr_5, sa33_sr_6, sa33_sr_7, u0_n49, u0_n53, u0_n55, u0_n57, u0_n59, 
       u0_n61, u0_n63, u0_subword_10, u0_subword_11, u0_subword_12, u0_subword_13, u0_subword_14, u0_subword_15, u0_subword_16, 
       u0_subword_17, u0_subword_18, u0_subword_19, u0_subword_20, u0_subword_21, u0_subword_22, u0_subword_23, u0_subword_24, u0_subword_25, 
       u0_subword_26, u0_subword_27, u0_subword_28, u0_subword_29, u0_subword_30, u0_subword_31, u0_subword_6, u0_subword_8, u0_subword_9, n101, n103, n105, n1109, n1114, n115, n117, n119, n121, 
        n13, n143, n15, n195, n197, n199, n201, n203, n207, 
        n209, n21, n213, n215, n217, n219, n225, n23, n231, 
        n247, n249, n25, n253, n3, n31, n33, n35, n37, 
        n47, n49, n5, n51, n53, n55, n57, n59, n61, 
        n63, n65, n67, n69, n7, n73, n79, n81, n85, 
        n9, sa00_0, sa00_1, sa00_2, sa00_3, sa00_4, sa00_5, sa00_6, sa00_7, 
        sa01_0, sa01_1, sa01_2, sa01_3, sa01_4, sa01_5, sa01_6, sa01_7, sa02_0, 
        sa02_1, sa02_2, sa02_3, sa02_4, sa02_5, sa02_6, sa02_7, sa03_0, sa03_1, 
        sa03_2, sa03_3, sa03_4, sa03_5, sa03_6, sa03_7, sa10_0, sa10_1, sa10_2, 
        sa10_3, sa10_4, sa10_5, sa10_6, sa10_7, sa11_0, sa11_1, sa11_2, sa11_3, 
        sa11_4, sa11_5, sa11_6, sa11_7, sa12_0, sa12_1, sa12_2, sa12_3, sa12_4, 
        sa12_5, sa12_6, sa12_7, sa13_0, sa13_1, sa13_2, sa13_3, sa13_4, sa13_5, 
        sa13_6, sa13_7, sa20_0, sa20_1, sa20_2, sa20_3, sa20_4, sa20_5, sa20_6, 
        sa20_7, sa21_0, sa21_1, sa21_2, sa21_3, sa21_4, sa21_5, sa21_6, sa21_7, 
        sa22_0, sa22_1, sa22_2, sa22_3, sa22_4, sa22_5, sa22_6, sa22_7, sa23_0, 
        sa23_1, sa23_2, sa23_3, sa23_4, sa23_5, sa23_6, sa23_7, sa30_0, sa30_1, 
        sa30_2, sa30_3, sa30_4, sa30_5, sa30_6, sa30_7, sa31_0, sa31_1, sa31_2, 
        sa31_3, sa31_4, sa31_5, sa31_6, sa31_7, sa32_0, sa32_1, sa32_2, sa32_3, 
        sa32_4, sa32_5, sa32_6, sa32_7, sa33_0, sa33_1, sa33_2, sa33_3, sa33_4, 
        sa33_5, sa33_6, sa33_7, u0_n268, u0_n270, u0_n272, u0_n274, w0_0, w0_1, 
        w0_10, w0_11, w0_12, w0_13, w0_15, w0_16, w0_18, w0_19, w0_2, 
        w0_20, w0_25, w0_26, w0_27, w0_28, w0_3, w0_30, w0_4, w0_5, 
        w0_7, w0_8, w1_4, w1_7, w2_0, w2_1, w2_10, w2_11, w2_13, 
        w2_16, w2_18, w2_19, w2_2, w2_20, w2_25, w2_26, w2_27, w2_28, 
        w2_4, w2_7, w2_8, w2_9, w3_0, w3_1, w3_10, w3_11, w3_12, 
        w3_13, w3_15, w3_16, w3_17, w3_18, w3_19, w3_2, w3_20, w3_21, 
        w3_22, w3_23, w3_24, w3_25, w3_26, w3_27, w3_28, w3_29, w3_3, 
        w3_30, w3_31, w3_4, w3_5, w3_6, w3_7, w3_8, w3_9 );
  input clk;
  input [127:0] key;
  input ld;
  input rst;
  input [127:0] text_in;
  output done;
  output [127:0] text_out;
  input N100, N102, N105, N114, N116, N132, N133, N134, N147, 
        N148, N149, N150, N169, N227, N228, N229, N230, N231, 
        N233, N242, N244, N245, N246, N247, N258, N261, N277, 
        N278, N280, N35, N36, N37, N38, N40, N41, N430, 
        N434, N435, N436, N437, N438, N439, N440, N441, N463, 
        N52, N53, N54, N57, N66, N67, N68, N73, N82, 
        N83, N84, N85, N86, N87, N88, N89, N98, N99, 
        n1145, n1183, n1212, n1213, n1214, n1215, n1216, n1217, n1219, 
        n1220, n1221, n342, n348, n354, n362, n394, n396, n414, 
        n419, n433, n462, n469, n481, n482, n500, n506, n515, 
        n524, n534, n547, n562, n590, n636, n657, n665, n786, 
        n791, n817, n823, n830, n861, n870, n900, n905, n911, 
        n917, n923, n927, n937, n957, sa00_sr_0, sa00_sr_1, sa00_sr_2, sa00_sr_3, 
        sa00_sr_4, sa00_sr_5, sa00_sr_6, sa00_sr_7, sa01_sr_0, sa01_sr_1, sa01_sr_2, sa01_sr_3, sa01_sr_4, 
        sa01_sr_5, sa01_sr_6, sa01_sr_7, sa02_sr_0, sa02_sr_1, sa02_sr_2, sa02_sr_3, sa02_sr_4, sa02_sr_5, 
        sa02_sr_6, sa02_sr_7, sa03_sr_0, sa03_sr_1, sa03_sr_2, sa03_sr_3, sa03_sr_4, sa03_sr_5, sa03_sr_6, 
        sa03_sr_7, sa10_sr_0, sa10_sr_1, sa10_sr_2, sa10_sr_3, sa10_sr_4, sa10_sr_5, sa10_sr_6, sa10_sr_7, 
        sa11_sr_0, sa11_sr_1, sa11_sr_2, sa11_sr_3, sa11_sr_4, sa11_sr_5, sa11_sr_6, sa11_sr_7, sa12_sr_0, 
        sa12_sr_1, sa12_sr_2, sa12_sr_4, sa12_sr_5, sa12_sr_6, sa12_sr_7, sa20_sr_0, sa20_sr_1, sa20_sr_2, 
        sa20_sr_3, sa20_sr_4, sa20_sr_5, sa20_sr_6, sa20_sr_7, sa21_sr_0, sa21_sr_1, sa21_sr_2, sa21_sr_3, 
        sa21_sr_4, sa21_sr_5, sa21_sr_6, sa21_sr_7, sa22_sr_0, sa22_sr_1, sa22_sr_3, sa22_sr_4, sa22_sr_5, 
        sa22_sr_6, sa22_sr_7, sa23_sr_0, sa23_sr_1, sa23_sr_2, sa23_sr_3, sa23_sr_4, sa23_sr_5, sa23_sr_6, 
        sa23_sr_7, sa30_sr_0, sa30_sr_1, sa30_sr_2, sa30_sr_3, sa30_sr_4, sa30_sr_5, sa30_sr_6, sa30_sr_7, 
        sa31_sr_0, sa31_sr_1, sa31_sr_2, sa31_sr_3, sa31_sr_4, sa31_sr_5, sa31_sr_6, sa31_sr_7, sa32_sr_0, 
        sa32_sr_1, sa32_sr_2, sa32_sr_3, sa32_sr_4, sa32_sr_5, sa32_sr_6, sa32_sr_7, sa33_sr_0, sa33_sr_1, 
        sa33_sr_2, sa33_sr_3, sa33_sr_4, sa33_sr_5, sa33_sr_6, sa33_sr_7, u0_n49, u0_n53, u0_n55, 
        u0_n57, u0_n59, u0_n61, u0_n63, u0_subword_10, u0_subword_11, u0_subword_12, u0_subword_13, u0_subword_14, 
        u0_subword_15, u0_subword_16, u0_subword_17, u0_subword_18, u0_subword_19, u0_subword_20, u0_subword_21, u0_subword_22, u0_subword_23, 
        u0_subword_24, u0_subword_25, u0_subword_26, u0_subword_27, u0_subword_28, u0_subword_29, u0_subword_30, u0_subword_31, u0_subword_6, 
        u0_subword_8, u0_subword_9;
  output n101, n103, n105, n1109, n1114, n115, n117, n119, n121, 
        n13, n143, n15, n195, n197, n199, n201, n203, n207, 
        n209, n21, n213, n215, n217, n219, n225, n23, n231, 
        n247, n249, n25, n253, n3, n31, n33, n35, n37, 
        n47, n49, n5, n51, n53, n55, n57, n59, n61, 
        n63, n65, n67, n69, n7, n73, n79, n81, n85, 
        n9, sa00_0, sa00_1, sa00_2, sa00_3, sa00_4, sa00_5, sa00_6, sa00_7, 
        sa01_0, sa01_1, sa01_2, sa01_3, sa01_4, sa01_5, sa01_6, sa01_7, sa02_0, 
        sa02_1, sa02_2, sa02_3, sa02_4, sa02_5, sa02_6, sa02_7, sa03_0, sa03_1, 
        sa03_2, sa03_3, sa03_4, sa03_5, sa03_6, sa03_7, sa10_0, sa10_1, sa10_2, 
        sa10_3, sa10_4, sa10_5, sa10_6, sa10_7, sa11_0, sa11_1, sa11_2, sa11_3, 
        sa11_4, sa11_5, sa11_6, sa11_7, sa12_0, sa12_1, sa12_2, sa12_3, sa12_4, 
        sa12_5, sa12_6, sa12_7, sa13_0, sa13_1, sa13_2, sa13_3, sa13_4, sa13_5, 
        sa13_6, sa13_7, sa20_0, sa20_1, sa20_2, sa20_3, sa20_4, sa20_5, sa20_6, 
        sa20_7, sa21_0, sa21_1, sa21_2, sa21_3, sa21_4, sa21_5, sa21_6, sa21_7, 
        sa22_0, sa22_1, sa22_2, sa22_3, sa22_4, sa22_5, sa22_6, sa22_7, sa23_0, 
        sa23_1, sa23_2, sa23_3, sa23_4, sa23_5, sa23_6, sa23_7, sa30_0, sa30_1, 
        sa30_2, sa30_3, sa30_4, sa30_5, sa30_6, sa30_7, sa31_0, sa31_1, sa31_2, 
        sa31_3, sa31_4, sa31_5, sa31_6, sa31_7, sa32_0, sa32_1, sa32_2, sa32_3, 
        sa32_4, sa32_5, sa32_6, sa32_7, sa33_0, sa33_1, sa33_2, sa33_3, sa33_4, 
        sa33_5, sa33_6, sa33_7, u0_n268, u0_n270, u0_n272, u0_n274, w0_0, w0_1, 
        w0_10, w0_11, w0_12, w0_13, w0_15, w0_16, w0_18, w0_19, w0_2, 
        w0_20, w0_25, w0_26, w0_27, w0_28, w0_3, w0_30, w0_4, w0_5, 
        w0_7, w0_8, w1_4, w1_7, w2_0, w2_1, w2_10, w2_11, w2_13, 
        w2_16, w2_18, w2_19, w2_2, w2_20, w2_25, w2_26, w2_27, w2_28, 
        w2_4, w2_7, w2_8, w2_9, w3_0, w3_1, w3_10, w3_11, w3_12, 
        w3_13, w3_15, w3_16, w3_17, w3_18, w3_19, w3_2, w3_20, w3_21, 
        w3_22, w3_23, w3_24, w3_25, w3_26, w3_27, w3_28, w3_29, w3_3, 
        w3_30, w3_31, w3_4, w3_5, w3_6, w3_7, w3_8, w3_9;
  wire N101, N103, N104, N115, N117, N118, N119, N120, N121, 
       N130, N131, N135, N136, N137, N146, N151, N152, N153, 
       N162, N163, N164, N165, N166, N167, N168, N178, N179, 
       N180, N181, N182, N183, N184, N185, N194, N195, N196, 
       N197, N198, N199, N200, N201, N210, N211, N212, N213, 
       N214, N215, N216, N217, N226, N23, N232, N243, N248, 
       N249, N259, N260, N262, N263, N264, N265, N274, N275, 
       N276, N279, N281, N34, N378, N379, N380, N381, N382, 
       N383, N384, N385, N386, N387, N388, N389, N39, N390, 
       N391, N392, N393, N394, N395, N396, N397, N398, N399, 
       N400, N401, N402, N403, N404, N405, N406, N407, N408, 
       N409, N410, N411, N412, N413, N414, N415, N416, N417, 
       N418, N419, N420, N421, N422, N423, N424, N425, N426, 
       N427, N428, N429, N431, N432, N433, N442, N443, N444, 
       N445, N446, N447, N448, N449, N450, N451, N452, N453, 
       N454, N455, N456, N457, N458, N459, N460, N461, N462, 
       N464, N465, N466, N467, N468, N469, N470, N471, N472, 
       N473, N474, N475, N476, N477, N478, N479, N480, N481, 
       N482, N483, N484, N485, N486, N487, N488, N489, N490, 
       N491, N492, N493, N494, N495, N496, N497, N498, N499, 
       N50, N500, N501, N502, N503, N504, N505, N51, N55, 
       N56, N69, N70, N71, N72, n1, n10, n100, n1000, 
       n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, 
       n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, 
       n1019, n102, n1020, n1021, n1022, n1023, n1024, n1025, n1026, 
       n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, 
       n1036, n1037, n1038, n1039, n104, n1040, n1041, n1042, n1043, 
       n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, 
       n1053, n1054, n1055, n1056, n1057, n1058, n1059, n106, n1060, 
       n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, 
       n107, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, 
       n1078, n1079, n108, n1080, n1081, n1082, n1083, n1084, n1085, 
       n1086, n1087, n1088, n1089, n109, n1090, n1091, n1092, n1093, 
       n1094, n1095, n1096, n1097, n1098, n1099, n11, n110, n1100, 
       n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n111, 
       n1110, n1111, n1112, n1113, n112, n1121, n1125, n1129, n113, 
       n1131, n1132, n1136, n114, n1143, n1146, n1147, n1151, n1152, 
       n1154, n1156, n1157, n1158, n1159, n116, n1160, n1161, n1162, 
       n1163, n1164, n1167, n1169, n1170, n1171, n1174, n1176, n1177, 
       n118, n1184, n1185, n1186, n1187, n1189, n1191, n1192, n1197, 
       n1198, n12, n120, n1206, n1207, n1218, n122, n1222, n123, 
       n124, n125, n126, n127, n128, n129, n130, n131, n132, 
       n133, n134, n135, n136, n137, n138, n139, n14, n140, 
       n141, n142, n144, n145, n146, n147, n148, n149, n150, 
       n151, n152, n153, n154, n155, n156, n157, n158, n159, 
       n16, n160, n161, n162, n163, n164, n165, n166, n167, 
       n168, n169, n17, n170, n171, n172, n173, n174, n175, 
       n176, n177, n178, n179, n18, n180, n181, n182, n183, 
       n184, n185, n186, n187, n188, n189, n19, n190, n191, 
       n192, n193, n194, n196, n198, n2, n20, n200, n202, 
       n204, n205, n206, n208, n210, n211, n212, n214, n216, 
       n218, n22, n220, n221, n222, n223, n224, n226, n227, 
       n228, n229, n230, n232, n233, n234, n235, n236, n237, 
       n238, n239, n24, n240, n241, n242, n243, n244, n245, 
       n246, n248, n250, n251, n252, n254, n255, n256, n258, 
       n259, n26, n260, n261, n262, n263, n264, n265, n266, 
       n267, n268, n269, n27, n270, n28, n29, n30, n32, 
       n34, n341, n347, n353, n36, n361, n38, n39, n391, 
       n392, n395, n4, n40, n41, n413, n418, n42, n43, 
       n432, n44, n45, n46, n461, n465, n466, n468, n470, 
       n471, n478, n479, n48, n499, n50, n505, n512, n513, 
       n517, n518, n519, n52, n520, n521, n522, n523, n526, 
       n528, n529, n530, n531, n532, n533, n54, n546, n551, 
       n552, n554, n555, n56, n561, n565, n566, n568, n58, 
       n587, n588, n591, n6, n60, n601, n602, n603, n605, 
       n62, n635, n639, n64, n640, n642, n643, n644, n645, 
       n646, n647, n649, n650, n651, n652, n653, n655, n656, 
       n658, n659, n66, n660, n661, n662, n663, n664, n666, 
       n667, n669, n670, n671, n672, n673, n674, n676, n677, 
       n678, n679, n68, n680, n682, n683, n684, n685, n686, 
       n687, n689, n690, n691, n692, n693, n694, n696, n697, 
       n698, n70, n700, n702, n703, n704, n705, n706, n707, 
       n708, n709, n71, n710, n711, n712, n713, n714, n715, 
       n716, n718, n719, n72, n720, n721, n722, n724, n725, 
       n726, n728, n729, n730, n731, n732, n734, n735, n736, 
       n738, n739, n74, n740, n742, n743, n744, n745, n746, 
       n747, n748, n749, n75, n750, n751, n752, n753, n755, 
       n756, n757, n758, n76, n760, n761, n762, n764, n765, 
       n766, n767, n769, n77, n775, n776, n777, n778, n779, 
       n78, n780, n781, n782, n783, n784, n785, n792, n793, 
       n794, n796, n797, n798, n799, n8, n80, n800, n801, 
       n802, n803, n804, n806, n807, n808, n809, n810, n812, 
       n813, n814, n816, n818, n819, n82, n820, n821, n826, 
       n827, n828, n829, n83, n831, n84, n858, n859, n86, 
       n863, n864, n865, n866, n867, n868, n869, n87, n872, 
       n874, n875, n876, n877, n878, n88, n89, n898, n899, 
       n90, n901, n902, n904, n908, n909, n91, n912, n913, 
       n915, n916, n92, n920, n921, n922, n925, n926, n93, 
       n936, n94, n95, n950, n951, n952, n954, n955, n956, 
       n958, n959, n96, n966, n967, n969, n97, n970, n977, 
       n978, n979, n98, n980, n981, n982, n983, n984, n985, 
       n986, n987, n988, n989, n99, n990, n991, n992, n993, 
       n994, n995, n996, n997, n998, n999, u0_N108, u0_N109, u0_N110, 
       u0_N111, u0_N112, u0_N113, u0_N114, u0_N115, u0_N116, u0_N117, u0_N118, u0_N119, 
       u0_N120, u0_N121, u0_N122, u0_N123, u0_N124, u0_N125, u0_N126, u0_N127, u0_N128, 
       u0_N129, u0_N130, u0_N131, u0_N132, u0_N133, u0_N134, u0_N135, u0_N136, u0_N137, 
       u0_N138, u0_N139, u0_N174, u0_N175, u0_N176, u0_N177, u0_N178, u0_N179, u0_N180, 
       u0_N181, u0_N182, u0_N183, u0_N184, u0_N185, u0_N186, u0_N187, u0_N188, u0_N189, 
       u0_N190, u0_N191, u0_N192, u0_N193, u0_N194, u0_N195, u0_N196, u0_N197, u0_N198, 
       u0_N199, u0_N200, u0_N201, u0_N202, u0_N203, u0_N204, u0_N205, u0_N240, u0_N241, 
       u0_N242, u0_N243, u0_N244, u0_N245, u0_N246, u0_N247, u0_N248, u0_N249, u0_N250, 
       u0_N251, u0_N252, u0_N253, u0_N254, u0_N255, u0_N256, u0_N257, u0_N258, u0_N259, 
       u0_N260, u0_N261, u0_N262, u0_N263, u0_N264, u0_N265, u0_N266, u0_N267, u0_N268, 
       u0_N269, u0_N270, u0_N271, u0_N42, u0_N43, u0_N44, u0_N45, u0_N46, u0_N47, 
       u0_N48, u0_N49, u0_N50, u0_N51, u0_N52, u0_N53, u0_N54, u0_N55, u0_N56, 
       u0_N57, u0_N58, u0_N59, u0_N60, u0_N61, u0_N62, u0_N63, u0_N64, u0_N65, 
       u0_N66, u0_N67, u0_N68, u0_N69, u0_N70, u0_N71, u0_N72, u0_N73, u0_n1, 
       u0_n10, u0_n100, u0_n101, u0_n102, u0_n103, u0_n104, u0_n105, u0_n106, u0_n107, 
       u0_n108, u0_n109, u0_n11, u0_n110, u0_n111, u0_n112, u0_n113, u0_n114, u0_n115, 
       u0_n116, u0_n117, u0_n118, u0_n119, u0_n12, u0_n120, u0_n121, u0_n122, u0_n123, 
       u0_n124, u0_n125, u0_n126, u0_n127, u0_n128, u0_n129, u0_n13, u0_n130, u0_n131, 
       u0_n132, u0_n133, u0_n134, u0_n135, u0_n136, u0_n137, u0_n138, u0_n139, u0_n14, 
       u0_n140, u0_n141, u0_n142, u0_n143, u0_n144, u0_n145, u0_n146, u0_n147, u0_n148, 
       u0_n149, u0_n15, u0_n150, u0_n151, u0_n152, u0_n153, u0_n154, u0_n155, u0_n156, 
       u0_n157, u0_n158, u0_n159, u0_n16, u0_n160, u0_n161, u0_n162, u0_n163, u0_n164, 
       u0_n165, u0_n166, u0_n167, u0_n168, u0_n169, u0_n17, u0_n170, u0_n171, u0_n172, 
       u0_n173, u0_n174, u0_n175, u0_n176, u0_n177, u0_n178, u0_n179, u0_n18, u0_n180, 
       u0_n181, u0_n182, u0_n183, u0_n184, u0_n185, u0_n186, u0_n187, u0_n188, u0_n189, 
       u0_n19, u0_n190, u0_n191, u0_n192, u0_n193, u0_n194, u0_n195, u0_n196, u0_n197, 
       u0_n198, u0_n199, u0_n2, u0_n20, u0_n200, u0_n201, u0_n202, u0_n203, u0_n204, 
       u0_n205, u0_n206, u0_n207, u0_n208, u0_n209, u0_n21, u0_n210, u0_n211, u0_n212, 
       u0_n213, u0_n214, u0_n215, u0_n216, u0_n217, u0_n218, u0_n219, u0_n22, u0_n220, 
       u0_n221, u0_n222, u0_n223, u0_n224, u0_n225, u0_n226, u0_n227, u0_n228, u0_n229, 
       u0_n23, u0_n230, u0_n231, u0_n232, u0_n233, u0_n234, u0_n235, u0_n236, u0_n237, 
       u0_n238, u0_n239, u0_n24, u0_n240, u0_n241, u0_n242, u0_n243, u0_n244, u0_n245, 
       u0_n246, u0_n247, u0_n248, u0_n249, u0_n25, u0_n250, u0_n251, u0_n253, u0_n254, 
       u0_n255, u0_n257, u0_n258, u0_n259, u0_n26, u0_n261, u0_n262, u0_n263, u0_n264, 
       u0_n265, u0_n267, u0_n269, u0_n27, u0_n271, u0_n273, u0_n275, u0_n277, u0_n279, 
       u0_n28, u0_n281, u0_n283, u0_n285, u0_n287, u0_n29, u0_n3, u0_n30, u0_n31, 
       u0_n32, u0_n33, u0_n34, u0_n35, u0_n36, u0_n37, u0_n38, u0_n39, u0_n4, 
       u0_n40, u0_n41, u0_n42, u0_n43, u0_n44, u0_n45, u0_n46, u0_n47, u0_n48, 
       u0_n5, u0_n50, u0_n51, u0_n52, u0_n54, u0_n56, u0_n58, u0_n6, u0_n60, 
       u0_n62, u0_n64, u0_n65, u0_n66, u0_n67, u0_n68, u0_n69, u0_n7, u0_n70, 
       u0_n71, u0_n72, u0_n73, u0_n74, u0_n75, u0_n76, u0_n77, u0_n78, u0_n79, 
       u0_n8, u0_n80, u0_n81, u0_n82, u0_n83, u0_n84, u0_n85, u0_n86, u0_n87, 
       u0_n88, u0_n89, u0_n9, u0_n90, u0_n91, u0_n92, u0_n93, u0_n94, u0_n95, 
       u0_n96, u0_n97, u0_n98, u0_n99, u0_r0_N70, u0_r0_N71, u0_r0_N72, u0_r0_N73, u0_r0_N74, 
       u0_r0_N75, u0_r0_N76, u0_r0_N77, u0_r0_N78, u0_r0_N79, u0_r0_N80, u0_r0_N81, u0_r0_n1, u0_r0_n10, 
       u0_r0_n11, u0_r0_n12, u0_r0_n13, u0_r0_n14, u0_r0_n15, u0_r0_n16, u0_r0_n17, u0_r0_n18, u0_r0_n19, 
       u0_r0_n2, u0_r0_n20, u0_r0_n21, u0_r0_n22, u0_r0_n23, u0_r0_n24, u0_r0_n25, u0_r0_n3, u0_r0_n4, 
       u0_r0_n5, u0_r0_n6, u0_r0_n7, u0_r0_n8, u0_r0_n9, u0_r0_rcnt_0, u0_r0_rcnt_1, u0_r0_rcnt_2, u0_rcon_24, 
       u0_rcon_25, u0_rcon_26, u0_rcon_27, u0_rcon_28, u0_rcon_29, u0_rcon_30, u0_rcon_31, w0_14, w0_17, 
       w0_21, w0_22, w0_23, w0_24, w0_29, w0_31, w0_6, w0_9, w1_0, 
       w1_1, w1_10, w1_11, w1_12, w1_13, w1_14, w1_15, w1_16, w1_17, 
       w1_18, w1_19, w1_2, w1_20, w1_21, w1_22, w1_23, w1_24, w1_25, 
       w1_26, w1_27, w1_28, w1_29, w1_3, w1_30, w1_31, w1_5, w1_6, 
       w1_8, w1_9, w2_12, w2_14, w2_15, w2_17, w2_21, w2_22, w2_23, 
       w2_24, w2_29, w2_3, w2_30, w2_31, w2_5, w2_6,  w3_14;
  NAND2_X1 U10 (.A2( ld ) , .ZN( n8 ) , .A1( text_in[3] ) );
  NAND2_X1 U100 (.A2( ld ) , .ZN( n98 ) , .A1( text_in[48] ) );
  XOR2_X1 U1001 (.Z( n728 ) , .B( n729 ) , .A( sa11_sr_0 ) );
  XOR2_X1 U1002 (.Z( n729 ) , .B( sa21_sr_0 ) , .A( w1_17 ) );
  XNOR2_X1 U1004 (.B( n683 ) , .ZN( n730 ) , .A( sa01_sr_1 ) );
  XOR2_X1 U1005 (.A( n163 ) , .Z( n725 ) , .B( w1_17 ) );
  OAI22_X1 U1007 (.ZN( N194 ) , .A1( n1214 ) , .B2( n1221 ) , .A2( n731 ) , .B1( n732 ) );
  XOR2_X1 U1009 (.A( n690 ) , .B( n713 ) , .Z( n734 ) );
  OAI21_X1 U101 (.B1( ld ) , .A( n100 ) , .ZN( n1027 ) , .B2( n99 ) );
  XOR2_X1 U1010 (.Z( n713 ) , .A( sa11_sr_7 ) , .B( sa21_sr_7 ) );
  XOR2_X1 U1012 (.A( n161 ) , .Z( n731 ) , .B( w1_16 ) );
  OAI22_X1 U1014 (.ZN( N185 ) , .A1( n1214 ) , .B2( n1220 ) , .A2( n735 ) , .B1( n736 ) );
  XOR2_X1 U1016 (.A( n650 ) , .B( n665 ) , .Z( n738 ) );
  XOR2_X1 U1017 (.Z( n650 ) , .A( sa21_sr_6 ) , .B( sa31_sr_6 ) );
  XOR2_X1 U1019 (.A( n159 ) , .Z( n735 ) , .B( w1_15 ) );
  NAND2_X1 U102 (.A2( ld ) , .ZN( n100 ) , .A1( text_in[49] ) );
  OAI22_X1 U1021 (.ZN( N184 ) , .A1( n1214 ) , .B2( n1220 ) , .A2( n739 ) , .B1( n740 ) );
  XOR2_X1 U1023 (.A( n644 ) , .B( n656 ) , .Z( n742 ) );
  XOR2_X1 U1024 (.Z( n656 ) , .A( sa21_sr_5 ) , .B( sa31_sr_5 ) );
  XOR2_X1 U1026 (.A( n157 ) , .Z( n739 ) , .B( w1_14 ) );
  OAI22_X1 U1028 (.ZN( N183 ) , .A1( n1109 ) , .B2( n1221 ) , .A2( n743 ) , .B1( n744 ) );
  XOR2_X1 U1029 (.Z( n744 ) , .A( n745 ) , .B( n746 ) );
  OAI21_X1 U103 (.B1( ld ) , .B2( n101 ) , .A( n102 ) , .ZN( n1028 ) );
  XOR2_X1 U1030 (.A( n651 ) , .B( n663 ) , .Z( n746 ) );
  XOR2_X1 U1031 (.Z( n663 ) , .A( sa21_sr_4 ) , .B( sa31_sr_4 ) );
  XNOR2_X1 U1032 (.ZN( n745 ) , .B( sa31_sr_5 ) , .A( w1_13 ) );
  XOR2_X1 U1033 (.A( n155 ) , .Z( n743 ) , .B( w1_13 ) );
  OAI22_X1 U1035 (.ZN( N182 ) , .A1( n1213 ) , .B2( n1221 ) , .A2( n747 ) , .B1( n748 ) );
  XOR2_X1 U1036 (.Z( n748 ) , .A( n749 ) , .B( n750 ) );
  XOR2_X1 U1037 (.A( n657 ) , .B( n670 ) , .Z( n750 ) );
  XOR2_X1 U1038 (.Z( n670 ) , .A( sa21_sr_3 ) , .B( sa31_sr_3 ) );
  XOR2_X1 U1039 (.B( n643 ) , .Z( n749 ) , .A( n751 ) );
  NAND2_X1 U104 (.A2( ld ) , .ZN( n102 ) , .A1( text_in[50] ) );
  XNOR2_X1 U1040 (.ZN( n751 ) , .B( sa31_sr_4 ) , .A( w1_12 ) );
  XOR2_X1 U1041 (.A( n153 ) , .Z( n747 ) , .B( w1_12 ) );
  OAI22_X1 U1043 (.ZN( N181 ) , .A1( n1214 ) , .B2( n1220 ) , .A2( n752 ) , .B1( n753 ) );
  XOR2_X1 U1045 (.A( n662 ) , .B( n677 ) , .Z( n755 ) );
  XOR2_X1 U1046 (.Z( n677 ) , .A( sa21_sr_2 ) , .B( sa31_sr_2 ) );
  XNOR2_X1 U1048 (.ZN( n756 ) , .B( sa31_sr_3 ) , .A( w1_11 ) );
  XOR2_X1 U1049 (.A( n151 ) , .Z( n752 ) , .B( w1_11 ) );
  OAI21_X1 U105 (.B1( ld ) , .ZN( n1029 ) , .B2( n103 ) , .A( n104 ) );
  OAI22_X1 U1051 (.ZN( N180 ) , .A1( n1109 ) , .B2( n1217 ) , .A2( n757 ) , .B1( n758 ) );
  XOR2_X1 U1053 (.A( n671 ) , .B( n683 ) , .Z( n760 ) );
  XOR2_X1 U1054 (.Z( n683 ) , .A( sa21_sr_1 ) , .B( sa31_sr_1 ) );
  XOR2_X1 U1056 (.A( n149 ) , .Z( n757 ) , .B( w1_10 ) );
  OAI22_X1 U1058 (.ZN( N179 ) , .A1( n1214 ) , .B2( n1220 ) , .A2( n761 ) , .B1( n762 ) );
  NAND2_X1 U106 (.A2( ld ) , .ZN( n104 ) , .A1( text_in[51] ) );
  XOR2_X1 U1060 (.A( n678 ) , .B( n690 ) , .Z( n764 ) );
  XOR2_X1 U1061 (.Z( n690 ) , .A( sa21_sr_0 ) , .B( sa31_sr_0 ) );
  XNOR2_X1 U1063 (.ZN( n765 ) , .B( sa31_sr_1 ) , .A( w1_9 ) );
  XOR2_X1 U1064 (.A( n147 ) , .Z( n761 ) , .B( w1_9 ) );
  OAI22_X1 U1066 (.ZN( N178 ) , .A1( n1214 ) , .B2( n1218 ) , .A2( n766 ) , .B1( n767 ) );
  XOR2_X1 U1068 (.A( n643 ) , .B( n684 ) , .Z( n769 ) );
  XOR2_X1 U1069 (.Z( n643 ) , .A( sa21_sr_7 ) , .B( sa31_sr_7 ) );
  OAI21_X1 U107 (.B1( ld ) , .ZN( n1030 ) , .B2( n105 ) , .A( n106 ) );
  XOR2_X1 U1071 (.A( n145 ) , .Z( n766 ) , .B( w1_8 ) );
  NAND2_X1 U108 (.A2( ld ) , .ZN( n106 ) , .A1( text_in[52] ) );
  OAI22_X1 U1081 (.ZN( N168 ) , .A1( n1213 ) , .B2( n1218 ) , .A2( n775 ) , .B1( n776 ) );
  XOR2_X1 U1082 (.Z( n776 ) , .A( n777 ) , .B( n778 ) );
  XOR2_X1 U1083 (.Z( n778 ) , .B( n779 ) , .A( sa21_sr_6 ) );
  XOR2_X1 U1084 (.Z( n779 ) , .B( sa31_sr_5 ) , .A( w1_6 ) );
  XNOR2_X1 U1085 (.B( n644 ) , .ZN( n777 ) , .A( sa01_sr_5 ) );
  XOR2_X1 U1086 (.Z( n644 ) , .A( sa01_sr_6 ) , .B( sa11_sr_6 ) );
  XOR2_X1 U1087 (.A( n141 ) , .Z( n775 ) , .B( w1_6 ) );
  OAI22_X1 U1089 (.ZN( N167 ) , .A1( n1212 ) , .B2( n1217 ) , .A2( n780 ) , .B1( n781 ) );
  OAI21_X1 U109 (.B1( ld ) , .ZN( n1031 ) , .B2( n107 ) , .A( n108 ) );
  XOR2_X1 U1090 (.Z( n781 ) , .A( n782 ) , .B( n783 ) );
  XOR2_X1 U1091 (.Z( n783 ) , .B( n784 ) , .A( sa21_sr_5 ) );
  XOR2_X1 U1092 (.Z( n784 ) , .B( sa31_sr_4 ) , .A( w1_5 ) );
  XNOR2_X1 U1093 (.B( n651 ) , .ZN( n782 ) , .A( sa01_sr_4 ) );
  XOR2_X1 U1094 (.Z( n651 ) , .A( sa01_sr_5 ) , .B( sa11_sr_5 ) );
  XOR2_X1 U1095 (.A( n139 ) , .Z( n780 ) , .B( w1_5 ) );
  OAI22_X1 U1097 (.ZN( N166 ) , .A1( n1213 ) , .B2( n1220 ) , .A2( n785 ) , .B1( n786 ) );
  OAI21_X1 U11 (.B1( ld ) , .A( n10 ) , .B2( n9 ) , .ZN( n982 ) );
  NAND2_X1 U110 (.A2( ld ) , .ZN( n108 ) , .A1( text_in[53] ) );
  XOR2_X1 U1104 (.A( n137 ) , .Z( n785 ) , .B( w1_4 ) );
  OAI22_X1 U1106 (.ZN( N165 ) , .A1( n1216 ) , .B2( n1217 ) , .A2( n792 ) , .B1( n793 ) );
  XOR2_X1 U1109 (.Z( n796 ) , .B( sa31_sr_2 ) , .A( w1_3 ) );
  OAI21_X1 U111 (.B1( ld ) , .ZN( n1032 ) , .B2( n109 ) , .A( n110 ) );
  XOR2_X1 U1110 (.B( n791 ) , .Z( n794 ) , .A( n797 ) );
  XNOR2_X1 U1111 (.B( n662 ) , .ZN( n797 ) , .A( sa01_sr_2 ) );
  XOR2_X1 U1112 (.Z( n662 ) , .A( sa01_sr_3 ) , .B( sa11_sr_3 ) );
  XOR2_X1 U1113 (.A( n135 ) , .Z( n792 ) , .B( w1_3 ) );
  OAI22_X1 U1115 (.ZN( N164 ) , .A1( n1213 ) , .B2( n1218 ) , .A2( n798 ) , .B1( n799 ) );
  XOR2_X1 U1116 (.Z( n799 ) , .A( n800 ) , .B( n801 ) );
  XOR2_X1 U1117 (.Z( n801 ) , .B( n802 ) , .A( sa21_sr_2 ) );
  XOR2_X1 U1118 (.Z( n802 ) , .B( sa31_sr_1 ) , .A( w1_2 ) );
  XNOR2_X1 U1119 (.B( n671 ) , .ZN( n800 ) , .A( sa01_sr_1 ) );
  NAND2_X1 U112 (.A2( ld ) , .ZN( n110 ) , .A1( text_in[54] ) );
  XOR2_X1 U1120 (.Z( n671 ) , .A( sa01_sr_2 ) , .B( sa11_sr_2 ) );
  XOR2_X1 U1121 (.A( n133 ) , .Z( n798 ) , .B( w1_2 ) );
  OAI22_X1 U1123 (.ZN( N163 ) , .A1( n1215 ) , .B2( n1220 ) , .A2( n803 ) , .B1( n804 ) );
  XOR2_X1 U1125 (.Z( n806 ) , .B( n807 ) , .A( sa21_sr_1 ) );
  XOR2_X1 U1126 (.Z( n807 ) , .B( sa31_sr_0 ) , .A( w1_1 ) );
  XNOR2_X1 U1128 (.B( n678 ) , .ZN( n808 ) , .A( sa01_sr_0 ) );
  XOR2_X1 U1129 (.Z( n678 ) , .A( sa01_sr_1 ) , .B( sa11_sr_1 ) );
  OAI21_X1 U113 (.B1( ld ) , .ZN( n1033 ) , .B2( n111 ) , .A( n112 ) );
  XOR2_X1 U1130 (.A( n131 ) , .Z( n803 ) , .B( w1_1 ) );
  OAI22_X1 U1132 (.ZN( N162 ) , .A1( n1215 ) , .B2( n1217 ) , .A2( n809 ) , .B1( n810 ) );
  XOR2_X1 U1134 (.A( n684 ) , .B( n791 ) , .Z( n812 ) );
  XOR2_X1 U1136 (.Z( n684 ) , .A( sa01_sr_0 ) , .B( sa11_sr_0 ) );
  XOR2_X1 U1138 (.A( n129 ) , .Z( n809 ) , .B( w1_0 ) );
  NAND2_X1 U114 (.A2( ld ) , .ZN( n112 ) , .A1( text_in[55] ) );
  OAI22_X1 U1140 (.ZN( N153 ) , .A1( n1215 ) , .B2( n1218 ) , .A2( n813 ) , .B1( n814 ) );
  XOR2_X1 U1142 (.Z( n816 ) , .A( n817 ) , .B( n818 ) );
  INV_X1 U1144 (.ZN( n819 ) , .A( sa12_sr_7 ) );
  XOR2_X1 U1145 (.A( n127 ) , .Z( n813 ) , .B( w2_31 ) );
  OAI22_X1 U1147 (.ZN( N152 ) , .A1( n1215 ) , .B2( n1217 ) , .A2( n820 ) , .B1( n821 ) );
  OAI21_X1 U115 (.B1( ld ) , .ZN( n1034 ) , .B2( n113 ) , .A( n114 ) );
  XOR2_X1 U1151 (.A( n125 ) , .Z( n820 ) , .B( w2_30 ) );
  OAI22_X1 U1153 (.ZN( N151 ) , .A1( n1215 ) , .B2( n1218 ) , .A2( n826 ) , .B1( n827 ) );
  XOR2_X1 U1154 (.Z( n827 ) , .A( n828 ) , .B( n829 ) );
  XOR2_X1 U1155 (.Z( n829 ) , .A( n830 ) , .B( n831 ) );
  XNOR2_X1 U1156 (.ZN( n828 ) , .B( sa12_sr_5 ) , .A( w2_29 ) );
  XOR2_X1 U1157 (.A( n123 ) , .Z( n826 ) , .B( w2_29 ) );
  NAND2_X1 U116 (.A2( ld ) , .ZN( n114 ) , .A1( text_in[56] ) );
  OAI21_X1 U117 (.B1( ld ) , .ZN( n1035 ) , .B2( n115 ) , .A( n116 ) );
  NAND2_X1 U118 (.A2( ld ) , .ZN( n116 ) , .A1( text_in[57] ) );
  OAI22_X1 U1186 (.ZN( N146 ) , .A1( n1215 ) , .B2( n1217 ) , .A2( n858 ) , .B1( n859 ) );
  OAI21_X1 U119 (.B1( ld ) , .ZN( n1036 ) , .B2( n117 ) , .A( n118 ) );
  XOR2_X1 U1190 (.A( n113 ) , .Z( n858 ) , .B( w2_24 ) );
  OAI22_X1 U1192 (.ZN( N137 ) , .A1( n1215 ) , .B2( n1218 ) , .A2( n863 ) , .B1( n864 ) );
  XOR2_X1 U1193 (.Z( n864 ) , .A( n865 ) , .B( n866 ) );
  XOR2_X1 U1194 (.B( n817 ) , .Z( n866 ) , .A( sa02_sr_7 ) );
  XNOR2_X1 U1195 (.ZN( n865 ) , .B( n867 ) , .A( sa12_sr_6 ) );
  XOR2_X1 U1196 (.Z( n867 ) , .B( sa22_sr_6 ) , .A( w2_23 ) );
  XOR2_X1 U1197 (.A( n111 ) , .Z( n863 ) , .B( w2_23 ) );
  OAI22_X1 U1199 (.ZN( N136 ) , .A1( n1215 ) , .B2( n1219 ) , .A2( n868 ) , .B1( n869 ) );
  NAND2_X1 U12 (.A2( ld ) , .ZN( n10 ) , .A1( text_in[4] ) );
  NAND2_X1 U120 (.A2( ld ) , .ZN( n118 ) , .A1( text_in[58] ) );
  XOR2_X1 U1202 (.Z( n872 ) , .B( sa22_sr_5 ) , .A( w2_22 ) );
  XOR2_X1 U1205 (.A( n109 ) , .Z( n868 ) , .B( w2_22 ) );
  OAI22_X1 U1207 (.ZN( N135 ) , .A1( n1213 ) , .B2( n1219 ) , .A2( n874 ) , .B1( n875 ) );
  XOR2_X1 U1208 (.Z( n875 ) , .A( n876 ) , .B( n877 ) );
  XOR2_X1 U1209 (.Z( n877 ) , .B( n878 ) , .A( sa12_sr_4 ) );
  OAI21_X1 U121 (.B1( ld ) , .ZN( n1037 ) , .B2( n119 ) , .A( n120 ) );
  XOR2_X1 U1210 (.Z( n878 ) , .B( sa22_sr_4 ) , .A( w2_21 ) );
  XNOR2_X1 U1211 (.B( n831 ) , .ZN( n876 ) , .A( sa02_sr_5 ) );
  XOR2_X1 U1212 (.A( n107 ) , .Z( n874 ) , .B( w2_21 ) );
  NAND2_X1 U122 (.A2( ld ) , .ZN( n120 ) , .A1( text_in[59] ) );
  OAI21_X1 U123 (.B1( ld ) , .ZN( n1038 ) , .B2( n121 ) , .A( n122 ) );
  OAI22_X1 U1238 (.ZN( N131 ) , .A1( n1212 ) , .B2( n1219 ) , .A2( n898 ) , .B1( n899 ) );
  XOR2_X1 U1239 (.Z( n899 ) , .A( n900 ) , .B( n901 ) );
  NAND2_X1 U124 (.A2( ld ) , .ZN( n122 ) , .A1( text_in[60] ) );
  XOR2_X1 U1240 (.Z( n901 ) , .B( n902 ) , .A( sa12_sr_0 ) );
  XOR2_X1 U1241 (.Z( n902 ) , .B( sa22_sr_0 ) , .A( w2_17 ) );
  XOR2_X1 U1244 (.Z( n898 ) , .A( n99 ) , .B( w2_17 ) );
  OAI22_X1 U1246 (.ZN( N130 ) , .A1( n1213 ) , .B2( n1219 ) , .A2( n904 ) , .B1( n905 ) );
  OAI21_X1 U125 (.B1( ld ) , .ZN( n1039 ) , .B2( n123 ) , .A( n124 ) );
  XOR2_X1 U1251 (.Z( n904 ) , .A( n97 ) , .B( w2_16 ) );
  OAI22_X1 U1253 (.ZN( N121 ) , .A1( n1109 ) , .B2( n1219 ) , .A2( n908 ) , .B1( n909 ) );
  XOR2_X1 U1258 (.Z( n908 ) , .A( n95 ) , .B( w2_15 ) );
  NAND2_X1 U126 (.A2( ld ) , .ZN( n124 ) , .A1( text_in[61] ) );
  OAI22_X1 U1260 (.ZN( N120 ) , .A1( n1109 ) , .B2( n1220 ) , .A2( n912 ) , .B1( n913 ) );
  XOR2_X1 U1262 (.A( n818 ) , .B( n831 ) , .Z( n915 ) );
  XOR2_X1 U1263 (.Z( n831 ) , .A( sa22_sr_5 ) , .B( sa32_sr_5 ) );
  XOR2_X1 U1265 (.Z( n912 ) , .A( n93 ) , .B( w2_14 ) );
  OAI22_X1 U1267 (.ZN( N119 ) , .A1( n1109 ) , .B2( n1218 ) , .A2( n916 ) , .B1( n917 ) );
  OAI21_X1 U127 (.B1( ld ) , .ZN( n1040 ) , .B2( n125 ) , .A( n126 ) );
  XOR2_X1 U1272 (.A( n91 ) , .Z( n916 ) , .B( w2_13 ) );
  OAI22_X1 U1274 (.ZN( N118 ) , .A1( n1109 ) , .B2( n1220 ) , .A2( n920 ) , .B1( n921 ) );
  XOR2_X1 U1275 (.Z( n921 ) , .A( n922 ) , .B( n923 ) );
  XOR2_X1 U1279 (.B( n817 ) , .Z( n922 ) , .A( n925 ) );
  NAND2_X1 U128 (.A2( ld ) , .ZN( n126 ) , .A1( text_in[62] ) );
  XNOR2_X1 U1280 (.ZN( n925 ) , .B( sa32_sr_4 ) , .A( w2_12 ) );
  XOR2_X1 U1281 (.A( n89 ) , .Z( n920 ) , .B( w2_12 ) );
  OAI22_X1 U1283 (.ZN( N117 ) , .A1( n1212 ) , .B2( n1220 ) , .A2( n926 ) , .B1( n927 ) );
  OAI21_X1 U129 (.B1( ld ) , .ZN( n1041 ) , .B2( n127 ) , .A( n128 ) );
  XOR2_X1 U1290 (.A( n87 ) , .Z( n926 ) , .B( w2_11 ) );
  OAI22_X1 U1299 (.ZN( N115 ) , .B2( n1114 ) , .A1( n1216 ) , .A2( n936 ) , .B1( n937 ) );
  OAI21_X1 U13 (.B1( ld ) , .B2( n11 ) , .A( n12 ) , .ZN( n983 ) );
  NAND2_X1 U130 (.A2( ld ) , .ZN( n128 ) , .A1( text_in[63] ) );
  XOR2_X1 U1306 (.A( n83 ) , .Z( n936 ) , .B( w2_9 ) );
  OAI21_X1 U131 (.B1( ld ) , .ZN( n1042 ) , .B2( n129 ) , .A( n130 ) );
  NAND2_X1 U132 (.A2( ld ) , .ZN( n130 ) , .A1( text_in[64] ) );
  OAI22_X1 U1324 (.ZN( N104 ) , .B2( n1114 ) , .A1( n1216 ) , .A2( n950 ) , .B1( n951 ) );
  XOR2_X1 U1327 (.Z( n954 ) , .B( sa32_sr_5 ) , .A( w2_6 ) );
  XNOR2_X1 U1328 (.B( n818 ) , .ZN( n952 ) , .A( sa02_sr_5 ) );
  XOR2_X1 U1329 (.Z( n818 ) , .A( sa02_sr_6 ) , .B( sa12_sr_6 ) );
  OAI21_X1 U133 (.B1( ld ) , .ZN( n1043 ) , .B2( n131 ) , .A( n132 ) );
  XOR2_X1 U1330 (.A( n77 ) , .Z( n950 ) , .B( w2_6 ) );
  OAI22_X1 U1332 (.ZN( N103 ) , .B2( n1114 ) , .A1( n1216 ) , .A2( n955 ) , .B1( n956 ) );
  XOR2_X1 U1333 (.Z( n956 ) , .A( n957 ) , .B( n958 ) );
  XOR2_X1 U1334 (.Z( n958 ) , .B( n959 ) , .A( sa22_sr_5 ) );
  XOR2_X1 U1335 (.Z( n959 ) , .B( sa32_sr_4 ) , .A( w2_5 ) );
  XOR2_X1 U1338 (.A( n75 ) , .Z( n955 ) , .B( w2_5 ) );
  NAND2_X1 U134 (.A2( ld ) , .ZN( n132 ) , .A1( text_in[65] ) );
  OAI22_X1 U1349 (.ZN( N101 ) , .B2( n1114 ) , .A1( n1216 ) , .A2( n966 ) , .B1( n967 ) );
  OAI21_X1 U135 (.B1( ld ) , .ZN( n1044 ) , .B2( n133 ) , .A( n134 ) );
  XOR2_X1 U1351 (.Z( n969 ) , .B( n970 ) , .A( sa22_sr_3 ) );
  XOR2_X1 U1352 (.Z( n970 ) , .B( sa32_sr_2 ) , .A( w2_3 ) );
  XOR2_X1 U1357 (.A( n71 ) , .Z( n966 ) , .B( w2_3 ) );
  NAND2_X1 U136 (.A2( ld ) , .ZN( n134 ) , .A1( text_in[66] ) );
  OAI21_X1 U137 (.B1( ld ) , .ZN( n1045 ) , .B2( n135 ) , .A( n136 ) );
  XOR2_X1 U1374 (.Z( N495 ) , .B( sa32_sr_2 ) , .A( w2_2 ) );
  NAND2_X1 U138 (.A2( ld ) , .ZN( n136 ) , .A1( text_in[67] ) );
  XNOR2_X1 U1381 (.B( n650 ) , .ZN( n698 ) , .A( sa01_sr_6 ) );
  BUF_X1 U1386 (.Z( n1218 ) , .A( n1221 ) );
  OAI21_X1 U139 (.B1( ld ) , .ZN( n1046 ) , .B2( n137 ) , .A( n138 ) );
  XNOR2_X1 U1391 (.A( n1121 ) , .ZN( n392 ) , .B( n394 ) );
  XOR2_X1 U1392 (.Z( n1121 ) , .B( sa33_sr_6 ) , .A( w3_14 ) );
  NAND2_X1 U14 (.A2( ld ) , .ZN( n12 ) , .A1( text_in[5] ) );
  NAND2_X1 U140 (.A2( ld ) , .ZN( n138 ) , .A1( text_in[68] ) );
  XNOR2_X1 U1401 (.A( n1125 ) , .ZN( n753 ) , .B( n755 ) );
  XNOR2_X1 U1402 (.ZN( n1125 ) , .B( n643 ) , .A( n756 ) );
  XNOR2_X1 U1409 (.A( n1129 ) , .ZN( n667 ) , .B( n669 ) );
  OAI21_X1 U141 (.B1( ld ) , .ZN( n1047 ) , .B2( n139 ) , .A( n140 ) );
  XNOR2_X1 U1410 (.ZN( n1129 ) , .B( n665 ) , .A( n672 ) );
  XNOR2_X1 U1413 (.B( n1131 ) , .ZN( n602 ) , .A( n603 ) );
  XNOR2_X1 U1414 (.ZN( n1131 ) , .B( n605 ) , .A( sa20_sr_6 ) );
  XNOR2_X1 U1415 (.A( n1132 ) , .ZN( n479 ) , .B( n481 ) );
  XOR2_X1 U1416 (.Z( n1132 ) , .B( sa10_sr_5 ) , .A( w0_29 ) );
  NAND2_X1 U142 (.A2( ld ) , .ZN( n140 ) , .A1( text_in[69] ) );
  XNOR2_X1 U1423 (.A( n1136 ) , .ZN( n814 ) , .B( n816 ) );
  XNOR2_X1 U1424 (.ZN( n1136 ) , .B( n819 ) , .A( w2_31 ) );
  OAI21_X1 U143 (.B1( ld ) , .ZN( n1048 ) , .B2( n141 ) , .A( n142 ) );
  XNOR2_X1 U1437 (.B( n1143 ) , .ZN( n715 ) , .A( n716 ) );
  XNOR2_X1 U1438 (.ZN( n1143 ) , .B( n718 ) , .A( sa11_sr_2 ) );
  NAND2_X1 U144 (.A2( ld ) , .ZN( n142 ) , .A1( text_in[70] ) );
  XNOR2_X1 U1441 (.A( n1145 ) , .ZN( n967 ) , .B( n969 ) );
  XNOR2_X1 U1443 (.A( n1146 ) , .ZN( n640 ) , .B( n642 ) );
  XNOR2_X1 U1444 (.ZN( n1146 ) , .B( n645 ) , .A( w1_31 ) );
  XNOR2_X1 U1445 (.A( n1147 ) , .ZN( n687 ) , .B( n689 ) );
  XOR2_X1 U1446 (.Z( n1147 ) , .B( sa11_sr_0 ) , .A( w1_24 ) );
  OAI21_X1 U145 (.B1( ld ) , .ZN( n1049 ) , .B2( n143 ) , .A( n144 ) );
  XNOR2_X1 U1453 (.A( n1151 ) , .ZN( n859 ) , .B( n861 ) );
  XOR2_X1 U1454 (.Z( n1151 ) , .B( sa12_sr_0 ) , .A( w2_24 ) );
  XNOR2_X1 U1455 (.A( n1152 ) , .ZN( n736 ) , .B( n738 ) );
  XOR2_X1 U1456 (.Z( n1152 ) , .B( sa31_sr_7 ) , .A( w1_15 ) );
  XNOR2_X1 U1459 (.A( n1154 ) , .ZN( n909 ) , .B( n911 ) );
  NAND2_X1 U146 (.A2( ld ) , .ZN( n144 ) , .A1( text_in[71] ) );
  XOR2_X1 U1460 (.Z( n1154 ) , .B( sa32_sr_7 ) , .A( w2_15 ) );
  XNOR2_X1 U1463 (.A( n1156 ) , .ZN( n821 ) , .B( n823 ) );
  XOR2_X1 U1464 (.Z( n1156 ) , .B( sa12_sr_6 ) , .A( w2_30 ) );
  XNOR2_X1 U1465 (.A( n1157 ) , .ZN( n647 ) , .B( n649 ) );
  XOR2_X1 U1466 (.Z( n1157 ) , .B( sa11_sr_6 ) , .A( w1_30 ) );
  XNOR2_X1 U1467 (.A( n1158 ) , .ZN( n588 ) , .B( n590 ) );
  XNOR2_X1 U1468 (.ZN( n1158 ) , .B( n469 ) , .A( n591 ) );
  XNOR2_X1 U1469 (.A( n1159 ) , .ZN( n762 ) , .B( n764 ) );
  OAI21_X1 U147 (.B1( ld ) , .ZN( n1050 ) , .B2( n145 ) , .A( n146 ) );
  XNOR2_X1 U1470 (.ZN( n1159 ) , .B( n643 ) , .A( n765 ) );
  XNOR2_X1 U1471 (.B( n1160 ) , .ZN( n523 ) , .A( n524 ) );
  XNOR2_X1 U1472 (.ZN( n1160 ) , .B( n526 ) , .A( sa10_sr_5 ) );
  XNOR2_X1 U1473 (.B( n1161 ) , .ZN( n869 ) , .A( n870 ) );
  XNOR2_X1 U1474 (.ZN( n1161 ) , .B( n872 ) , .A( sa12_sr_5 ) );
  XNOR2_X1 U1475 (.B( n1162 ) , .ZN( n697 ) , .A( n698 ) );
  XNOR2_X1 U1476 (.ZN( n1162 ) , .B( n700 ) , .A( sa11_sr_5 ) );
  XNOR2_X1 U1477 (.A( n1163 ) , .ZN( n740 ) , .B( n742 ) );
  XOR2_X1 U1478 (.Z( n1163 ) , .B( sa31_sr_6 ) , .A( w1_14 ) );
  XNOR2_X1 U1479 (.A( n1164 ) , .ZN( n913 ) , .B( n915 ) );
  NAND2_X1 U148 (.A2( ld ) , .ZN( n146 ) , .A1( text_in[72] ) );
  XOR2_X1 U1480 (.Z( n1164 ) , .B( sa32_sr_6 ) , .A( w2_14 ) );
  XNOR2_X1 U1485 (.B( n1167 ) , .ZN( n793 ) , .A( n794 ) );
  XNOR2_X1 U1486 (.ZN( n1167 ) , .B( n796 ) , .A( sa21_sr_3 ) );
  XNOR2_X1 U1489 (.A( n1169 ) , .ZN( n566 ) , .B( n568 ) );
  OAI21_X1 U149 (.B1( ld ) , .ZN( n1051 ) , .B2( n147 ) , .A( n148 ) );
  XOR2_X1 U1490 (.Z( n1169 ) , .B( sa30_sr_6 ) , .A( w0_14 ) );
  XNOR2_X1 U1491 (.A( n1170 ) , .ZN( n767 ) , .B( n769 ) );
  XOR2_X1 U1492 (.Z( n1170 ) , .B( sa31_sr_0 ) , .A( w1_8 ) );
  XNOR2_X1 U1493 (.A( n1171 ) , .ZN( n732 ) , .B( n734 ) );
  XOR2_X1 U1494 (.Z( n1171 ) , .B( sa01_sr_0 ) , .A( w1_16 ) );
  XNOR2_X1 U1499 (.A( n1174 ) , .ZN( n653 ) , .B( n655 ) );
  OAI21_X1 U15 (.B1( ld ) , .B2( n13 ) , .A( n14 ) , .ZN( n984 ) );
  NAND2_X1 U150 (.A2( ld ) , .ZN( n148 ) , .A1( text_in[73] ) );
  XOR2_X1 U1500 (.Z( n1174 ) , .B( sa11_sr_5 ) , .A( w1_29 ) );
  XNOR2_X1 U1503 (.B( n1176 ) , .ZN( n721 ) , .A( n722 ) );
  XNOR2_X1 U1504 (.ZN( n1176 ) , .B( n724 ) , .A( sa11_sr_1 ) );
  XNOR2_X1 U1505 (.A( n1177 ) , .ZN( n680 ) , .B( n682 ) );
  XNOR2_X1 U1506 (.ZN( n1177 ) , .B( n665 ) , .A( n685 ) );
  OAI21_X1 U151 (.B1( ld ) , .ZN( n1052 ) , .B2( n149 ) , .A( n150 ) );
  XNOR2_X1 U1517 (.A( n1183 ) , .ZN( n552 ) , .B( n554 ) );
  XNOR2_X1 U1519 (.A( n1184 ) , .ZN( n810 ) , .B( n812 ) );
  NAND2_X1 U152 (.A2( ld ) , .ZN( n150 ) , .A1( text_in[74] ) );
  XOR2_X1 U1520 (.Z( n1184 ) , .B( sa21_sr_0 ) , .A( w1_0 ) );
  XNOR2_X1 U1521 (.A( n1185 ) , .ZN( n726 ) , .B( n728 ) );
  XNOR2_X1 U1522 (.ZN( n1185 ) , .B( n713 ) , .A( n730 ) );
  XNOR2_X1 U1523 (.B( n1186 ) , .ZN( n951 ) , .A( n952 ) );
  XNOR2_X1 U1524 (.ZN( n1186 ) , .B( n954 ) , .A( sa22_sr_6 ) );
  XNOR2_X1 U1525 (.A( n1187 ) , .ZN( n804 ) , .B( n806 ) );
  XNOR2_X1 U1526 (.ZN( n1187 ) , .B( n791 ) , .A( n808 ) );
  XOR2_X1 U1529 (.B( n1189 ) , .Z( n693 ) , .A( sa11_sr_6 ) );
  OAI21_X1 U153 (.B1( ld ) , .ZN( n1053 ) , .B2( n151 ) , .A( n152 ) );
  XNOR2_X1 U1530 (.ZN( n1189 ) , .B( sa21_sr_6 ) , .A( w1_23 ) );
  XNOR2_X1 U1533 (.A( n1191 ) , .ZN( n466 ) , .B( n468 ) );
  XNOR2_X1 U1534 (.ZN( n1191 ) , .B( n471 ) , .A( w0_31 ) );
  XNOR2_X1 U1535 (.A( n1192 ) , .ZN( n513 ) , .B( n515 ) );
  XOR2_X1 U1536 (.Z( n1192 ) , .B( sa10_sr_0 ) , .A( w0_24 ) );
  NAND2_X1 U154 (.A2( ld ) , .ZN( n152 ) , .A1( text_in[75] ) );
  XNOR2_X1 U1545 (.A( n1197 ) , .ZN( n674 ) , .B( n676 ) );
  XOR2_X1 U1546 (.Z( n1197 ) , .B( sa11_sr_2 ) , .A( w1_26 ) );
  XNOR2_X1 U1547 (.A( n1198 ) , .ZN( n758 ) , .B( n760 ) );
  XOR2_X1 U1548 (.Z( n1198 ) , .B( sa31_sr_2 ) , .A( w1_10 ) );
  OAI21_X1 U155 (.B1( ld ) , .ZN( n1054 ) , .B2( n153 ) , .A( n154 ) );
  NAND2_X1 U156 (.A2( ld ) , .ZN( n154 ) , .A1( text_in[76] ) );
  XNOR2_X1 U1563 (.ZN( N415 ) , .B( n1206 ) , .A( w0_18 ) );
  XNOR2_X1 U1566 (.ZN( N423 ) , .B( n1207 ) , .A( w1_18 ) );
  INV_X1 U1567 (.ZN( n1206 ) , .A( sa10_sr_2 ) );
  INV_X1 U1568 (.ZN( n1207 ) , .A( sa11_sr_2 ) );
  OAI21_X1 U157 (.B1( ld ) , .ZN( n1055 ) , .B2( n155 ) , .A( n156 ) );
  INV_X1 U1576 (.A( ld ) , .ZN( n1222 ) );
  NAND2_X1 U158 (.A2( ld ) , .ZN( n156 ) , .A1( text_in[77] ) );
  OAI21_X1 U159 (.B1( ld ) , .ZN( n1056 ) , .B2( n157 ) , .A( n158 ) );
  NAND2_X1 U16 (.A2( ld ) , .ZN( n14 ) , .A1( text_in[6] ) );
  NAND2_X1 U160 (.A2( ld ) , .ZN( n158 ) , .A1( text_in[78] ) );
  OAI21_X1 U161 (.B1( ld ) , .ZN( n1057 ) , .B2( n159 ) , .A( n160 ) );
  NAND2_X1 U162 (.A2( ld ) , .ZN( n160 ) , .A1( text_in[79] ) );
  OAI21_X1 U163 (.B1( ld ) , .ZN( n1058 ) , .B2( n161 ) , .A( n162 ) );
  NAND2_X1 U164 (.A2( ld ) , .ZN( n162 ) , .A1( text_in[80] ) );
  OAI21_X1 U165 (.B1( ld ) , .ZN( n1059 ) , .B2( n163 ) , .A( n164 ) );
  NAND2_X1 U166 (.A2( ld ) , .ZN( n164 ) , .A1( text_in[81] ) );
  OAI21_X1 U167 (.B1( ld ) , .ZN( n1060 ) , .B2( n165 ) , .A( n166 ) );
  NAND2_X1 U168 (.A2( ld ) , .ZN( n166 ) , .A1( text_in[82] ) );
  OAI21_X1 U169 (.B1( ld ) , .ZN( n1061 ) , .B2( n167 ) , .A( n168 ) );
  OAI21_X1 U17 (.B1( ld ) , .B2( n15 ) , .A( n16 ) , .ZN( n985 ) );
  NAND2_X1 U170 (.A2( ld ) , .ZN( n168 ) , .A1( text_in[83] ) );
  OAI21_X1 U171 (.B1( ld ) , .ZN( n1062 ) , .B2( n169 ) , .A( n170 ) );
  NAND2_X1 U172 (.A2( ld ) , .ZN( n170 ) , .A1( text_in[84] ) );
  OAI21_X1 U173 (.B1( ld ) , .ZN( n1063 ) , .B2( n171 ) , .A( n172 ) );
  NAND2_X1 U174 (.A2( ld ) , .ZN( n172 ) , .A1( text_in[85] ) );
  OAI21_X1 U175 (.B1( ld ) , .ZN( n1064 ) , .B2( n173 ) , .A( n174 ) );
  NAND2_X1 U176 (.A2( ld ) , .ZN( n174 ) , .A1( text_in[86] ) );
  OAI21_X1 U177 (.B1( ld ) , .ZN( n1065 ) , .B2( n175 ) , .A( n176 ) );
  NAND2_X1 U178 (.A2( ld ) , .ZN( n176 ) , .A1( text_in[87] ) );
  OAI21_X1 U179 (.B1( ld ) , .ZN( n1066 ) , .B2( n177 ) , .A( n178 ) );
  NAND2_X1 U18 (.A2( ld ) , .ZN( n16 ) , .A1( text_in[7] ) );
  NAND2_X1 U180 (.A2( ld ) , .ZN( n178 ) , .A1( text_in[88] ) );
  OAI21_X1 U181 (.B1( ld ) , .ZN( n1067 ) , .B2( n179 ) , .A( n180 ) );
  NAND2_X1 U182 (.A2( ld ) , .ZN( n180 ) , .A1( text_in[89] ) );
  OAI21_X1 U183 (.B1( ld ) , .ZN( n1068 ) , .B2( n181 ) , .A( n182 ) );
  NAND2_X1 U184 (.A2( ld ) , .ZN( n182 ) , .A1( text_in[90] ) );
  OAI21_X1 U185 (.B1( ld ) , .ZN( n1069 ) , .B2( n183 ) , .A( n184 ) );
  NAND2_X1 U186 (.A2( ld ) , .ZN( n184 ) , .A1( text_in[91] ) );
  OAI21_X1 U187 (.B1( ld ) , .ZN( n1070 ) , .B2( n185 ) , .A( n186 ) );
  NAND2_X1 U188 (.A2( ld ) , .ZN( n186 ) , .A1( text_in[92] ) );
  OAI21_X1 U189 (.B1( ld ) , .ZN( n1071 ) , .B2( n187 ) , .A( n188 ) );
  OAI21_X1 U19 (.B1( ld ) , .B2( n17 ) , .A( n18 ) , .ZN( n986 ) );
  NAND2_X1 U190 (.A2( ld ) , .ZN( n188 ) , .A1( text_in[93] ) );
  OAI21_X1 U191 (.B1( ld ) , .ZN( n1072 ) , .B2( n189 ) , .A( n190 ) );
  NAND2_X1 U192 (.A2( ld ) , .ZN( n190 ) , .A1( text_in[94] ) );
  OAI21_X1 U193 (.B1( ld ) , .ZN( n1073 ) , .B2( n191 ) , .A( n192 ) );
  NAND2_X1 U194 (.A2( ld ) , .ZN( n192 ) , .A1( text_in[95] ) );
  OAI21_X1 U195 (.B1( ld ) , .ZN( n1074 ) , .B2( n193 ) , .A( n194 ) );
  NAND2_X1 U196 (.A2( ld ) , .ZN( n194 ) , .A1( text_in[96] ) );
  OAI21_X1 U197 (.B1( ld ) , .ZN( n1075 ) , .B2( n195 ) , .A( n196 ) );
  NAND2_X1 U198 (.A2( ld ) , .ZN( n196 ) , .A1( text_in[97] ) );
  OAI21_X1 U199 (.B1( ld ) , .ZN( n1076 ) , .B2( n197 ) , .A( n198 ) );
  NAND2_X1 U20 (.A2( ld ) , .ZN( n18 ) , .A1( text_in[8] ) );
  NAND2_X1 U200 (.A2( ld ) , .ZN( n198 ) , .A1( text_in[98] ) );
  OAI21_X1 U201 (.B1( ld ) , .ZN( n1077 ) , .B2( n199 ) , .A( n200 ) );
  NAND2_X1 U202 (.A2( ld ) , .ZN( n200 ) , .A1( text_in[99] ) );
  OAI21_X1 U203 (.B1( ld ) , .ZN( n1078 ) , .B2( n201 ) , .A( n202 ) );
  NAND2_X1 U204 (.A2( ld ) , .ZN( n202 ) , .A1( text_in[100] ) );
  OAI21_X1 U205 (.B1( ld ) , .ZN( n1079 ) , .B2( n203 ) , .A( n204 ) );
  NAND2_X1 U206 (.A2( ld ) , .ZN( n204 ) , .A1( text_in[101] ) );
  OAI21_X1 U207 (.B1( ld ) , .ZN( n1080 ) , .B2( n205 ) , .A( n206 ) );
  NAND2_X1 U208 (.A2( ld ) , .ZN( n206 ) , .A1( text_in[102] ) );
  OAI21_X1 U209 (.B1( ld ) , .ZN( n1081 ) , .B2( n207 ) , .A( n208 ) );
  OAI21_X1 U21 (.B1( ld ) , .B2( n19 ) , .A( n20 ) , .ZN( n987 ) );
  NAND2_X1 U210 (.A2( ld ) , .ZN( n208 ) , .A1( text_in[103] ) );
  OAI21_X1 U211 (.B1( ld ) , .ZN( n1082 ) , .B2( n209 ) , .A( n210 ) );
  NAND2_X1 U212 (.A2( ld ) , .ZN( n210 ) , .A1( text_in[104] ) );
  OAI21_X1 U213 (.B1( ld ) , .ZN( n1083 ) , .B2( n211 ) , .A( n212 ) );
  NAND2_X1 U214 (.A2( ld ) , .ZN( n212 ) , .A1( text_in[105] ) );
  OAI21_X1 U215 (.B1( ld ) , .ZN( n1084 ) , .B2( n213 ) , .A( n214 ) );
  NAND2_X1 U216 (.A2( ld ) , .ZN( n214 ) , .A1( text_in[106] ) );
  OAI21_X1 U217 (.B1( ld ) , .ZN( n1085 ) , .B2( n215 ) , .A( n216 ) );
  NAND2_X1 U218 (.A2( ld ) , .ZN( n216 ) , .A1( text_in[107] ) );
  OAI21_X1 U219 (.B1( ld ) , .ZN( n1086 ) , .B2( n217 ) , .A( n218 ) );
  NAND2_X1 U22 (.A2( ld ) , .ZN( n20 ) , .A1( text_in[9] ) );
  NAND2_X1 U220 (.A2( ld ) , .ZN( n218 ) , .A1( text_in[108] ) );
  OAI21_X1 U221 (.B1( ld ) , .ZN( n1087 ) , .B2( n219 ) , .A( n220 ) );
  NAND2_X1 U222 (.A2( ld ) , .ZN( n220 ) , .A1( text_in[109] ) );
  OAI21_X1 U223 (.B1( ld ) , .ZN( n1088 ) , .B2( n221 ) , .A( n222 ) );
  NAND2_X1 U224 (.A2( ld ) , .ZN( n222 ) , .A1( text_in[110] ) );
  OAI21_X1 U225 (.B1( ld ) , .ZN( n1089 ) , .B2( n223 ) , .A( n224 ) );
  NAND2_X1 U226 (.A2( ld ) , .ZN( n224 ) , .A1( text_in[111] ) );
  OAI21_X1 U227 (.B1( ld ) , .ZN( n1090 ) , .B2( n225 ) , .A( n226 ) );
  NAND2_X1 U228 (.A2( ld ) , .ZN( n226 ) , .A1( text_in[112] ) );
  OAI21_X1 U229 (.B1( ld ) , .ZN( n1091 ) , .B2( n227 ) , .A( n228 ) );
  OAI21_X1 U23 (.B1( ld ) , .B2( n21 ) , .A( n22 ) , .ZN( n988 ) );
  NAND2_X1 U230 (.A2( ld ) , .ZN( n228 ) , .A1( text_in[113] ) );
  OAI21_X1 U231 (.B1( ld ) , .ZN( n1092 ) , .B2( n229 ) , .A( n230 ) );
  NAND2_X1 U232 (.A2( ld ) , .ZN( n230 ) , .A1( text_in[114] ) );
  OAI21_X1 U233 (.B1( ld ) , .ZN( n1093 ) , .B2( n231 ) , .A( n232 ) );
  NAND2_X1 U234 (.A2( ld ) , .ZN( n232 ) , .A1( text_in[115] ) );
  OAI21_X1 U235 (.B1( ld ) , .ZN( n1094 ) , .B2( n233 ) , .A( n234 ) );
  NAND2_X1 U236 (.A2( ld ) , .ZN( n234 ) , .A1( text_in[116] ) );
  OAI21_X1 U237 (.B1( ld ) , .ZN( n1095 ) , .B2( n235 ) , .A( n236 ) );
  NAND2_X1 U238 (.A2( ld ) , .ZN( n236 ) , .A1( text_in[117] ) );
  OAI21_X1 U239 (.B1( ld ) , .ZN( n1096 ) , .B2( n237 ) , .A( n238 ) );
  NAND2_X1 U24 (.A2( ld ) , .ZN( n22 ) , .A1( text_in[10] ) );
  NAND2_X1 U240 (.A2( ld ) , .ZN( n238 ) , .A1( text_in[118] ) );
  OAI21_X1 U241 (.B1( ld ) , .ZN( n1097 ) , .B2( n239 ) , .A( n240 ) );
  NAND2_X1 U242 (.A2( ld ) , .ZN( n240 ) , .A1( text_in[119] ) );
  OAI21_X1 U243 (.B1( ld ) , .ZN( n1098 ) , .B2( n241 ) , .A( n242 ) );
  NAND2_X1 U244 (.A2( ld ) , .ZN( n242 ) , .A1( text_in[120] ) );
  OAI21_X1 U245 (.B1( ld ) , .ZN( n1099 ) , .B2( n243 ) , .A( n244 ) );
  NAND2_X1 U246 (.A2( ld ) , .ZN( n244 ) , .A1( text_in[121] ) );
  OAI21_X1 U247 (.B1( ld ) , .ZN( n1100 ) , .B2( n245 ) , .A( n246 ) );
  NAND2_X1 U248 (.A2( ld ) , .ZN( n246 ) , .A1( text_in[122] ) );
  OAI21_X1 U249 (.B1( ld ) , .ZN( n1101 ) , .B2( n247 ) , .A( n248 ) );
  OAI21_X1 U25 (.B1( ld ) , .B2( n23 ) , .A( n24 ) , .ZN( n989 ) );
  NAND2_X1 U250 (.A2( ld ) , .ZN( n248 ) , .A1( text_in[123] ) );
  OAI21_X1 U251 (.B1( ld ) , .ZN( n1102 ) , .B2( n249 ) , .A( n250 ) );
  NAND2_X1 U252 (.A2( ld ) , .ZN( n250 ) , .A1( text_in[124] ) );
  OAI21_X1 U253 (.B1( ld ) , .ZN( n1103 ) , .B2( n251 ) , .A( n252 ) );
  NAND2_X1 U254 (.A2( ld ) , .ZN( n252 ) , .A1( text_in[125] ) );
  OAI21_X1 U255 (.B1( ld ) , .ZN( n1104 ) , .B2( n253 ) , .A( n254 ) );
  NAND2_X1 U256 (.A2( ld ) , .ZN( n254 ) , .A1( text_in[126] ) );
  OAI21_X1 U257 (.B1( ld ) , .ZN( n1105 ) , .B2( n255 ) , .A( n256 ) );
  NAND2_X1 U258 (.A2( ld ) , .ZN( n256 ) , .A1( text_in[127] ) );
  AOI21_X1 U259 (.ZN( n1110 ) , .B1( n1222 ) , .B2( n258 ) , .A( n259 ) );
  NAND2_X1 U26 (.A2( ld ) , .ZN( n24 ) , .A1( text_in[11] ) );
  OAI21_X1 U260 (.ZN( n258 ) , .B1( n260 ) , .B2( n261 ) , .A( n262 ) );
  NOR3_X1 U261 (.A2( ld ) , .ZN( n1111 ) , .A1( n259 ) , .A3( n263 ) );
  AOI22_X1 U262 (.ZN( n263 ) , .A1( n264 ) , .A2( n265 ) , .B1( n266 ) , .B2( n267 ) );
  NOR2_X1 U263 (.A1( n1106 ) , .ZN( n264 ) , .A2( n267 ) );
  INV_X1 U265 (.ZN( n1112 ) , .A( n268 ) );
  OAI21_X1 U266 (.B1( ld ) , .ZN( n268 ) , .B2( n269 ) , .A( rst ) );
  AOI21_X1 U267 (.A( n1106 ) , .B1( n1107 ) , .B2( n265 ) , .ZN( n269 ) );
  INV_X1 U268 (.ZN( n265 ) , .A( n266 ) );
  NAND2_X1 U269 (.A1( n1108 ) , .A2( n262 ) , .ZN( n266 ) );
  OAI21_X1 U27 (.B1( ld ) , .B2( n25 ) , .A( n26 ) , .ZN( n990 ) );
  XNOR2_X1 U270 (.B( n261 ) , .ZN( n262 ) , .A( n977 ) );
  AOI21_X1 U272 (.ZN( n1113 ) , .B1( n1222 ) , .A( n259 ) , .B2( n270 ) );
  INV_X1 U273 (.ZN( n259 ) , .A( rst ) );
  OAI21_X1 U274 (.A( n1108 ) , .B2( n260 ) , .ZN( n270 ) , .B1( n977 ) );
  NAND2_X1 U28 (.A2( ld ) , .ZN( n26 ) , .A1( text_in[12] ) );
  OAI21_X1 U29 (.B1( ld ) , .B2( n27 ) , .A( n28 ) , .ZN( n991 ) );
  OAI21_X1 U3 (.B1( ld ) , .B2( n1 ) , .A( n2 ) , .ZN( n978 ) );
  NAND2_X1 U30 (.A2( ld ) , .ZN( n28 ) , .A1( text_in[13] ) );
  OAI21_X1 U31 (.B1( ld ) , .B2( n29 ) , .A( n30 ) , .ZN( n992 ) );
  NAND2_X1 U32 (.A2( ld ) , .ZN( n30 ) , .A1( text_in[14] ) );
  OAI21_X1 U33 (.B1( ld ) , .B2( n31 ) , .A( n32 ) , .ZN( n993 ) );
  NAND2_X1 U34 (.A2( ld ) , .ZN( n32 ) , .A1( text_in[15] ) );
  OAI22_X1 U348 (.ZN( N72 ) , .A1( n1212 ) , .B2( n1217 ) , .A2( n341 ) , .B1( n342 ) );
  OAI21_X1 U35 (.B1( ld ) , .B2( n33 ) , .A( n34 ) , .ZN( n994 ) );
  XOR2_X1 U354 (.Z( n341 ) , .A( n45 ) , .B( w3_22 ) );
  OAI22_X1 U356 (.ZN( N71 ) , .A1( n1214 ) , .B2( n1221 ) , .A2( n347 ) , .B1( n348 ) );
  NAND2_X1 U36 (.A2( ld ) , .ZN( n34 ) , .A1( text_in[16] ) );
  XOR2_X1 U361 (.Z( n347 ) , .A( n43 ) , .B( w3_21 ) );
  OAI22_X1 U363 (.ZN( N70 ) , .B2( n1114 ) , .A1( n1213 ) , .A2( n353 ) , .B1( n354 ) );
  XOR2_X1 U369 (.Z( n353 ) , .A( n41 ) , .B( w3_20 ) );
  OAI21_X1 U37 (.B1( ld ) , .B2( n35 ) , .A( n36 ) , .ZN( n995 ) );
  OAI22_X1 U371 (.ZN( N69 ) , .B2( n1114 ) , .A1( n1212 ) , .A2( n361 ) , .B1( n362 ) );
  XOR2_X1 U377 (.Z( n361 ) , .A( n39 ) , .B( w3_19 ) );
  NAND2_X1 U38 (.A2( ld ) , .ZN( n36 ) , .A1( text_in[17] ) );
  OAI21_X1 U39 (.B1( ld ) , .B2( n37 ) , .A( n38 ) , .ZN( n996 ) );
  NAND2_X1 U4 (.A2( ld ) , .ZN( n2 ) , .A1( text_in[0] ) );
  NAND2_X1 U40 (.A2( ld ) , .ZN( n38 ) , .A1( text_in[18] ) );
  OAI22_X1 U408 (.ZN( N56 ) , .B2( n1114 ) , .A1( n1213 ) , .A2( n391 ) , .B1( n392 ) );
  OAI21_X1 U41 (.B1( ld ) , .B2( n39 ) , .A( n40 ) , .ZN( n997 ) );
  XOR2_X1 U413 (.A( n29 ) , .Z( n391 ) , .B( w3_14 ) );
  OAI22_X1 U415 (.ZN( N55 ) , .A1( n1216 ) , .B2( n1221 ) , .A2( n395 ) , .B1( n396 ) );
  NAND2_X1 U42 (.A2( ld ) , .ZN( n40 ) , .A1( text_in[19] ) );
  XOR2_X1 U420 (.A( n27 ) , .Z( n395 ) , .B( w3_13 ) );
  OAI21_X1 U43 (.B1( ld ) , .B2( n41 ) , .A( n42 ) , .ZN( n998 ) );
  NAND2_X1 U44 (.A2( ld ) , .ZN( n42 ) , .A1( text_in[20] ) );
  OAI22_X1 U445 (.ZN( N51 ) , .A1( n1214 ) , .B2( n1217 ) , .A2( n413 ) , .B1( n414 ) );
  OAI21_X1 U45 (.B1( ld ) , .B2( n43 ) , .A( n44 ) , .ZN( n999 ) );
  XOR2_X1 U451 (.A( n19 ) , .Z( n413 ) , .B( w3_9 ) );
  XOR2_X1 U453 (.Z( N505 ) , .B( sa33_sr_0 ) , .A( w3_0 ) );
  XOR2_X1 U454 (.Z( N504 ) , .B( sa33_sr_1 ) , .A( w3_1 ) );
  XOR2_X1 U455 (.Z( N503 ) , .B( sa33_sr_2 ) , .A( w3_2 ) );
  XOR2_X1 U456 (.Z( N502 ) , .B( sa33_sr_3 ) , .A( w3_3 ) );
  XOR2_X1 U457 (.Z( N501 ) , .B( sa33_sr_4 ) , .A( w3_4 ) );
  XOR2_X1 U458 (.Z( N500 ) , .B( sa33_sr_5 ) , .A( w3_5 ) );
  OAI22_X1 U459 (.ZN( N50 ) , .A1( n1214 ) , .B2( n1218 ) , .A2( n418 ) , .B1( n419 ) );
  NAND2_X1 U46 (.A2( ld ) , .ZN( n44 ) , .A1( text_in[21] ) );
  XOR2_X1 U464 (.A( n17 ) , .Z( n418 ) , .B( w3_8 ) );
  XOR2_X1 U466 (.Z( N499 ) , .B( sa33_sr_6 ) , .A( w3_6 ) );
  XOR2_X1 U467 (.Z( N498 ) , .B( sa33_sr_7 ) , .A( w3_7 ) );
  XOR2_X1 U468 (.Z( N497 ) , .B( sa32_sr_0 ) , .A( w2_0 ) );
  XOR2_X1 U469 (.Z( N496 ) , .B( sa32_sr_1 ) , .A( w2_1 ) );
  OAI21_X1 U47 (.B1( ld ) , .ZN( n1000 ) , .B2( n45 ) , .A( n46 ) );
  XOR2_X1 U471 (.Z( N494 ) , .B( sa32_sr_3 ) , .A( w2_3 ) );
  XOR2_X1 U472 (.Z( N493 ) , .B( sa32_sr_4 ) , .A( w2_4 ) );
  XOR2_X1 U473 (.Z( N492 ) , .B( sa32_sr_5 ) , .A( w2_5 ) );
  XOR2_X1 U474 (.Z( N491 ) , .B( sa32_sr_6 ) , .A( w2_6 ) );
  XOR2_X1 U475 (.Z( N490 ) , .B( sa32_sr_7 ) , .A( w2_7 ) );
  XOR2_X1 U476 (.Z( N489 ) , .B( sa31_sr_0 ) , .A( w1_0 ) );
  XOR2_X1 U477 (.Z( N488 ) , .B( sa31_sr_1 ) , .A( w1_1 ) );
  XOR2_X1 U478 (.Z( N487 ) , .B( sa31_sr_2 ) , .A( w1_2 ) );
  XOR2_X1 U479 (.Z( N486 ) , .B( sa31_sr_3 ) , .A( w1_3 ) );
  NAND2_X1 U48 (.A2( ld ) , .ZN( n46 ) , .A1( text_in[22] ) );
  XOR2_X1 U480 (.Z( N485 ) , .B( sa31_sr_4 ) , .A( w1_4 ) );
  XOR2_X1 U481 (.Z( N484 ) , .B( sa31_sr_5 ) , .A( w1_5 ) );
  XOR2_X1 U482 (.Z( N483 ) , .B( sa31_sr_6 ) , .A( w1_6 ) );
  XOR2_X1 U483 (.Z( N482 ) , .B( sa31_sr_7 ) , .A( w1_7 ) );
  XOR2_X1 U484 (.Z( N481 ) , .B( sa30_sr_0 ) , .A( w0_0 ) );
  XOR2_X1 U485 (.Z( N480 ) , .B( sa30_sr_1 ) , .A( w0_1 ) );
  XOR2_X1 U486 (.Z( N479 ) , .B( sa30_sr_2 ) , .A( w0_2 ) );
  XOR2_X1 U487 (.Z( N478 ) , .B( sa30_sr_3 ) , .A( w0_3 ) );
  XOR2_X1 U488 (.Z( N477 ) , .B( sa30_sr_4 ) , .A( w0_4 ) );
  XOR2_X1 U489 (.Z( N476 ) , .B( sa30_sr_5 ) , .A( w0_5 ) );
  OAI21_X1 U49 (.B1( ld ) , .ZN( n1001 ) , .B2( n47 ) , .A( n48 ) );
  XOR2_X1 U490 (.Z( N475 ) , .B( sa30_sr_6 ) , .A( w0_6 ) );
  XOR2_X1 U491 (.Z( N474 ) , .B( sa30_sr_7 ) , .A( w0_7 ) );
  XOR2_X1 U492 (.Z( N473 ) , .B( sa23_sr_0 ) , .A( w3_8 ) );
  XOR2_X1 U493 (.Z( N472 ) , .B( sa23_sr_1 ) , .A( w3_9 ) );
  XOR2_X1 U494 (.Z( N471 ) , .B( sa23_sr_2 ) , .A( w3_10 ) );
  XOR2_X1 U495 (.Z( N470 ) , .B( sa23_sr_3 ) , .A( w3_11 ) );
  XOR2_X1 U496 (.Z( N469 ) , .B( sa23_sr_4 ) , .A( w3_12 ) );
  XOR2_X1 U497 (.Z( N468 ) , .B( sa23_sr_5 ) , .A( w3_13 ) );
  XOR2_X1 U498 (.Z( N467 ) , .B( sa23_sr_6 ) , .A( w3_14 ) );
  XOR2_X1 U499 (.Z( N466 ) , .B( sa23_sr_7 ) , .A( w3_15 ) );
  OAI21_X1 U5 (.B1( ld ) , .B2( n3 ) , .A( n4 ) , .ZN( n979 ) );
  NAND2_X1 U50 (.A2( ld ) , .ZN( n48 ) , .A1( text_in[23] ) );
  XOR2_X1 U500 (.Z( N465 ) , .B( sa22_sr_0 ) , .A( w2_8 ) );
  XOR2_X1 U501 (.Z( N464 ) , .B( sa22_sr_1 ) , .A( w2_9 ) );
  XOR2_X1 U503 (.Z( N462 ) , .B( sa22_sr_3 ) , .A( w2_11 ) );
  XOR2_X1 U504 (.Z( N461 ) , .B( sa22_sr_4 ) , .A( w2_12 ) );
  XOR2_X1 U505 (.Z( N460 ) , .B( sa22_sr_5 ) , .A( w2_13 ) );
  XOR2_X1 U506 (.Z( N459 ) , .B( sa22_sr_6 ) , .A( w2_14 ) );
  XOR2_X1 U507 (.Z( N458 ) , .B( sa22_sr_7 ) , .A( w2_15 ) );
  XOR2_X1 U508 (.Z( N457 ) , .B( sa21_sr_0 ) , .A( w1_8 ) );
  XOR2_X1 U509 (.Z( N456 ) , .B( sa21_sr_1 ) , .A( w1_9 ) );
  OAI21_X1 U51 (.B1( ld ) , .ZN( n1002 ) , .B2( n49 ) , .A( n50 ) );
  XOR2_X1 U510 (.Z( N455 ) , .B( sa21_sr_2 ) , .A( w1_10 ) );
  XOR2_X1 U511 (.Z( N454 ) , .B( sa21_sr_3 ) , .A( w1_11 ) );
  XOR2_X1 U512 (.Z( N453 ) , .B( sa21_sr_4 ) , .A( w1_12 ) );
  XOR2_X1 U513 (.Z( N452 ) , .B( sa21_sr_5 ) , .A( w1_13 ) );
  XOR2_X1 U514 (.Z( N451 ) , .B( sa21_sr_6 ) , .A( w1_14 ) );
  XOR2_X1 U515 (.Z( N450 ) , .B( sa21_sr_7 ) , .A( w1_15 ) );
  XOR2_X1 U516 (.Z( N449 ) , .B( sa20_sr_0 ) , .A( w0_8 ) );
  XOR2_X1 U517 (.Z( N448 ) , .B( sa20_sr_1 ) , .A( w0_9 ) );
  XOR2_X1 U518 (.Z( N447 ) , .B( sa20_sr_2 ) , .A( w0_10 ) );
  XOR2_X1 U519 (.Z( N446 ) , .B( sa20_sr_3 ) , .A( w0_11 ) );
  NAND2_X1 U52 (.A2( ld ) , .ZN( n50 ) , .A1( text_in[24] ) );
  XOR2_X1 U520 (.Z( N445 ) , .B( sa20_sr_4 ) , .A( w0_12 ) );
  XOR2_X1 U521 (.Z( N444 ) , .B( sa20_sr_5 ) , .A( w0_13 ) );
  XOR2_X1 U522 (.Z( N443 ) , .B( sa20_sr_6 ) , .A( w0_14 ) );
  XOR2_X1 U523 (.Z( N442 ) , .B( sa20_sr_7 ) , .A( w0_15 ) );
  OAI21_X1 U53 (.B1( ld ) , .ZN( n1003 ) , .B2( n51 ) , .A( n52 ) );
  XOR2_X1 U532 (.Z( N433 ) , .B( sa12_sr_0 ) , .A( w2_16 ) );
  XOR2_X1 U533 (.Z( N432 ) , .B( sa12_sr_1 ) , .A( w2_17 ) );
  XOR2_X1 U534 (.Z( N431 ) , .B( sa12_sr_2 ) , .A( w2_18 ) );
  XOR2_X1 U536 (.Z( N429 ) , .B( sa12_sr_4 ) , .A( w2_20 ) );
  XOR2_X1 U537 (.Z( N428 ) , .B( sa12_sr_5 ) , .A( w2_21 ) );
  XOR2_X1 U538 (.Z( N427 ) , .B( sa12_sr_6 ) , .A( w2_22 ) );
  XOR2_X1 U539 (.Z( N426 ) , .B( sa12_sr_7 ) , .A( w2_23 ) );
  NAND2_X1 U54 (.A2( ld ) , .ZN( n52 ) , .A1( text_in[25] ) );
  XOR2_X1 U540 (.Z( N425 ) , .B( sa11_sr_0 ) , .A( w1_16 ) );
  XOR2_X1 U541 (.Z( N424 ) , .B( sa11_sr_1 ) , .A( w1_17 ) );
  XOR2_X1 U543 (.Z( N422 ) , .B( sa11_sr_3 ) , .A( w1_19 ) );
  XOR2_X1 U544 (.Z( N421 ) , .B( sa11_sr_4 ) , .A( w1_20 ) );
  XOR2_X1 U545 (.Z( N420 ) , .B( sa11_sr_5 ) , .A( w1_21 ) );
  XOR2_X1 U546 (.Z( N419 ) , .B( sa11_sr_6 ) , .A( w1_22 ) );
  XOR2_X1 U547 (.Z( N418 ) , .B( sa11_sr_7 ) , .A( w1_23 ) );
  XOR2_X1 U548 (.Z( N417 ) , .B( sa10_sr_0 ) , .A( w0_16 ) );
  XOR2_X1 U549 (.Z( N416 ) , .B( sa10_sr_1 ) , .A( w0_17 ) );
  OAI21_X1 U55 (.B1( ld ) , .ZN( n1004 ) , .B2( n53 ) , .A( n54 ) );
  XOR2_X1 U551 (.Z( N414 ) , .B( sa10_sr_3 ) , .A( w0_19 ) );
  XOR2_X1 U552 (.Z( N413 ) , .B( sa10_sr_4 ) , .A( w0_20 ) );
  XOR2_X1 U553 (.Z( N412 ) , .B( sa10_sr_5 ) , .A( w0_21 ) );
  XOR2_X1 U554 (.Z( N411 ) , .B( sa10_sr_6 ) , .A( w0_22 ) );
  XOR2_X1 U555 (.Z( N410 ) , .B( sa10_sr_7 ) , .A( w0_23 ) );
  NAND2_X1 U56 (.A2( ld ) , .ZN( n54 ) , .A1( text_in[26] ) );
  XOR2_X1 U565 (.Z( N409 ) , .B( sa03_sr_0 ) , .A( w3_24 ) );
  XOR2_X1 U566 (.Z( N408 ) , .B( sa03_sr_1 ) , .A( w3_25 ) );
  XOR2_X1 U567 (.Z( N407 ) , .B( sa03_sr_2 ) , .A( w3_26 ) );
  XOR2_X1 U568 (.Z( N406 ) , .B( sa03_sr_3 ) , .A( w3_27 ) );
  XOR2_X1 U569 (.Z( N405 ) , .B( sa03_sr_4 ) , .A( w3_28 ) );
  OAI21_X1 U57 (.B1( ld ) , .ZN( n1005 ) , .B2( n55 ) , .A( n56 ) );
  XOR2_X1 U570 (.Z( N404 ) , .B( sa03_sr_5 ) , .A( w3_29 ) );
  XOR2_X1 U571 (.Z( N403 ) , .B( sa03_sr_6 ) , .A( w3_30 ) );
  XOR2_X1 U572 (.Z( N402 ) , .B( sa03_sr_7 ) , .A( w3_31 ) );
  XOR2_X1 U573 (.Z( N401 ) , .B( sa02_sr_0 ) , .A( w2_24 ) );
  XOR2_X1 U574 (.Z( N400 ) , .B( sa02_sr_1 ) , .A( w2_25 ) );
  NAND2_X1 U58 (.A2( ld ) , .ZN( n56 ) , .A1( text_in[27] ) );
  XOR2_X1 U584 (.Z( N399 ) , .B( sa02_sr_2 ) , .A( w2_26 ) );
  XOR2_X1 U585 (.Z( N398 ) , .B( sa02_sr_3 ) , .A( w2_27 ) );
  XOR2_X1 U586 (.Z( N397 ) , .B( sa02_sr_4 ) , .A( w2_28 ) );
  XOR2_X1 U587 (.Z( N396 ) , .B( sa02_sr_5 ) , .A( w2_29 ) );
  XOR2_X1 U588 (.Z( N395 ) , .B( sa02_sr_6 ) , .A( w2_30 ) );
  XOR2_X1 U589 (.Z( N394 ) , .B( sa02_sr_7 ) , .A( w2_31 ) );
  OAI21_X1 U59 (.B1( ld ) , .ZN( n1006 ) , .B2( n57 ) , .A( n58 ) );
  XOR2_X1 U590 (.Z( N393 ) , .B( sa01_sr_0 ) , .A( w1_24 ) );
  XOR2_X1 U591 (.Z( N392 ) , .B( sa01_sr_1 ) , .A( w1_25 ) );
  XOR2_X1 U592 (.Z( N391 ) , .B( sa01_sr_2 ) , .A( w1_26 ) );
  XOR2_X1 U593 (.Z( N390 ) , .B( sa01_sr_3 ) , .A( w1_27 ) );
  OAI22_X1 U594 (.ZN( N39 ) , .A1( n1214 ) , .B2( n1218 ) , .A2( n432 ) , .B1( n433 ) );
  NAND2_X1 U6 (.A2( ld ) , .ZN( n4 ) , .A1( text_in[1] ) );
  NAND2_X1 U60 (.A2( ld ) , .ZN( n58 ) , .A1( text_in[28] ) );
  XOR2_X1 U601 (.A( n11 ) , .Z( n432 ) , .B( w3_5 ) );
  XOR2_X1 U603 (.Z( N389 ) , .B( sa01_sr_4 ) , .A( w1_28 ) );
  XOR2_X1 U604 (.Z( N388 ) , .B( sa01_sr_5 ) , .A( w1_29 ) );
  XOR2_X1 U605 (.Z( N387 ) , .B( sa01_sr_6 ) , .A( w1_30 ) );
  XOR2_X1 U606 (.Z( N386 ) , .B( sa01_sr_7 ) , .A( w1_31 ) );
  XOR2_X1 U607 (.Z( N385 ) , .B( sa00_sr_0 ) , .A( w0_24 ) );
  XOR2_X1 U608 (.Z( N384 ) , .B( sa00_sr_1 ) , .A( w0_25 ) );
  XOR2_X1 U609 (.Z( N383 ) , .B( sa00_sr_2 ) , .A( w0_26 ) );
  OAI21_X1 U61 (.B1( ld ) , .ZN( n1007 ) , .B2( n59 ) , .A( n60 ) );
  XOR2_X1 U610 (.Z( N382 ) , .B( sa00_sr_3 ) , .A( w0_27 ) );
  XOR2_X1 U611 (.Z( N381 ) , .B( sa00_sr_4 ) , .A( w0_28 ) );
  XOR2_X1 U612 (.Z( N380 ) , .B( sa00_sr_5 ) , .A( w0_29 ) );
  NAND2_X1 U62 (.A2( ld ) , .ZN( n60 ) , .A1( text_in[29] ) );
  XOR2_X1 U623 (.Z( N379 ) , .B( sa00_sr_6 ) , .A( w0_30 ) );
  XOR2_X1 U624 (.Z( N378 ) , .B( sa00_sr_7 ) , .A( w0_31 ) );
  OAI21_X1 U63 (.B1( ld ) , .ZN( n1008 ) , .B2( n61 ) , .A( n62 ) );
  NAND2_X1 U64 (.A2( ld ) , .ZN( n62 ) , .A1( text_in[30] ) );
  OAI21_X1 U65 (.B1( ld ) , .ZN( n1009 ) , .B2( n63 ) , .A( n64 ) );
  OAI22_X1 U654 (.ZN( N34 ) , .A1( n1214 ) , .B2( n1218 ) , .A2( n461 ) , .B1( n462 ) );
  NAND2_X1 U66 (.A2( ld ) , .ZN( n64 ) , .A1( text_in[31] ) );
  XOR2_X1 U660 (.A( n1 ) , .Z( n461 ) , .B( w3_0 ) );
  OAI22_X1 U662 (.ZN( N281 ) , .A1( n1214 ) , .B2( n1221 ) , .A2( n465 ) , .B1( n466 ) );
  XOR2_X1 U664 (.Z( n468 ) , .A( n469 ) , .B( n470 ) );
  INV_X1 U666 (.ZN( n471 ) , .A( sa10_sr_7 ) );
  XOR2_X1 U667 (.A( n255 ) , .Z( n465 ) , .B( w0_31 ) );
  OAI21_X1 U67 (.B1( ld ) , .ZN( n1010 ) , .B2( n65 ) , .A( n66 ) );
  OAI22_X1 U675 (.ZN( N279 ) , .A1( n1212 ) , .B2( n1218 ) , .A2( n478 ) , .B1( n479 ) );
  XOR2_X1 U679 (.A( n251 ) , .Z( n478 ) , .B( w0_29 ) );
  NAND2_X1 U68 (.A2( ld ) , .ZN( n66 ) , .A1( text_in[32] ) );
  OAI21_X1 U69 (.B1( ld ) , .ZN( n1011 ) , .B2( n67 ) , .A( n68 ) );
  OAI22_X1 U695 (.ZN( N276 ) , .A1( n1212 ) , .B2( n1220 ) , .A2( n499 ) , .B1( n500 ) );
  XOR2_X1 U699 (.A( n245 ) , .Z( n499 ) , .B( w0_26 ) );
  OAI21_X1 U7 (.B1( ld ) , .B2( n5 ) , .A( n6 ) , .ZN( n980 ) );
  NAND2_X1 U70 (.A2( ld ) , .ZN( n68 ) , .A1( text_in[33] ) );
  OAI22_X1 U701 (.ZN( N275 ) , .A1( n1213 ) , .B2( n1220 ) , .A2( n505 ) , .B1( n506 ) );
  XOR2_X1 U706 (.A( n243 ) , .Z( n505 ) , .B( w0_25 ) );
  OAI22_X1 U708 (.ZN( N274 ) , .A1( n1216 ) , .B2( n1221 ) , .A2( n512 ) , .B1( n513 ) );
  OAI21_X1 U71 (.B1( ld ) , .ZN( n1012 ) , .B2( n69 ) , .A( n70 ) );
  XOR2_X1 U712 (.A( n241 ) , .Z( n512 ) , .B( w0_24 ) );
  OAI22_X1 U714 (.ZN( N265 ) , .B2( n1114 ) , .A1( n1215 ) , .A2( n517 ) , .B1( n518 ) );
  XOR2_X1 U715 (.Z( n518 ) , .A( n519 ) , .B( n520 ) );
  XOR2_X1 U716 (.B( n469 ) , .Z( n520 ) , .A( sa00_sr_7 ) );
  XNOR2_X1 U717 (.ZN( n519 ) , .B( n521 ) , .A( sa10_sr_6 ) );
  XOR2_X1 U718 (.Z( n521 ) , .B( sa20_sr_6 ) , .A( w0_23 ) );
  XOR2_X1 U719 (.A( n239 ) , .Z( n517 ) , .B( w0_23 ) );
  NAND2_X1 U72 (.A2( ld ) , .ZN( n70 ) , .A1( text_in[34] ) );
  OAI22_X1 U721 (.ZN( N264 ) , .A1( n1213 ) , .B2( n1220 ) , .A2( n522 ) , .B1( n523 ) );
  XOR2_X1 U724 (.Z( n526 ) , .B( sa20_sr_5 ) , .A( w0_22 ) );
  XOR2_X1 U727 (.A( n237 ) , .Z( n522 ) , .B( w0_22 ) );
  OAI22_X1 U729 (.ZN( N263 ) , .A1( n1213 ) , .B2( n1221 ) , .A2( n528 ) , .B1( n529 ) );
  OAI21_X1 U73 (.B1( ld ) , .ZN( n1013 ) , .B2( n71 ) , .A( n72 ) );
  XOR2_X1 U730 (.Z( n529 ) , .A( n530 ) , .B( n531 ) );
  XOR2_X1 U731 (.Z( n531 ) , .B( n532 ) , .A( sa10_sr_4 ) );
  XOR2_X1 U732 (.Z( n532 ) , .B( sa20_sr_4 ) , .A( w0_21 ) );
  XNOR2_X1 U733 (.B( n482 ) , .ZN( n530 ) , .A( sa00_sr_5 ) );
  XOR2_X1 U734 (.A( n235 ) , .Z( n528 ) , .B( w0_21 ) );
  OAI22_X1 U736 (.ZN( N262 ) , .A1( n1213 ) , .B2( n1218 ) , .A2( n533 ) , .B1( n534 ) );
  NAND2_X1 U74 (.A2( ld ) , .ZN( n72 ) , .A1( text_in[35] ) );
  XOR2_X1 U742 (.A( n233 ) , .Z( n533 ) , .B( w0_20 ) );
  OAI21_X1 U75 (.B1( ld ) , .ZN( n1014 ) , .B2( n73 ) , .A( n74 ) );
  OAI22_X1 U752 (.ZN( N260 ) , .A1( n1213 ) , .B2( n1218 ) , .A2( n546 ) , .B1( n547 ) );
  XOR2_X1 U757 (.A( n229 ) , .Z( n546 ) , .B( w0_18 ) );
  OAI22_X1 U759 (.ZN( N259 ) , .A1( n1109 ) , .B2( n1218 ) , .A2( n551 ) , .B1( n552 ) );
  NAND2_X1 U76 (.A2( ld ) , .ZN( n74 ) , .A1( text_in[36] ) );
  XOR2_X1 U761 (.Z( n554 ) , .B( n555 ) , .A( sa10_sr_0 ) );
  XOR2_X1 U762 (.Z( n555 ) , .B( sa20_sr_0 ) , .A( w0_17 ) );
  XOR2_X1 U765 (.A( n227 ) , .Z( n551 ) , .B( w0_17 ) );
  OAI21_X1 U77 (.B1( ld ) , .ZN( n1015 ) , .B2( n75 ) , .A( n76 ) );
  OAI22_X1 U774 (.ZN( N249 ) , .A1( n1109 ) , .B2( n1217 ) , .A2( n561 ) , .B1( n562 ) );
  XOR2_X1 U779 (.A( n223 ) , .Z( n561 ) , .B( w0_15 ) );
  NAND2_X1 U78 (.A2( ld ) , .ZN( n76 ) , .A1( text_in[37] ) );
  OAI22_X1 U781 (.ZN( N248 ) , .A1( n1109 ) , .B2( n1220 ) , .A2( n565 ) , .B1( n566 ) );
  XOR2_X1 U783 (.A( n470 ) , .B( n482 ) , .Z( n568 ) );
  XOR2_X1 U786 (.A( n221 ) , .Z( n565 ) , .B( w0_14 ) );
  OAI21_X1 U79 (.B1( ld ) , .ZN( n1016 ) , .B2( n77 ) , .A( n78 ) );
  NAND2_X1 U8 (.A2( ld ) , .ZN( n6 ) , .A1( text_in[2] ) );
  NAND2_X1 U80 (.A2( ld ) , .ZN( n78 ) , .A1( text_in[38] ) );
  OAI21_X1 U81 (.B1( ld ) , .ZN( n1017 ) , .B2( n79 ) , .A( n80 ) );
  OAI22_X1 U818 (.ZN( N243 ) , .A1( n1212 ) , .B2( n1220 ) , .A2( n587 ) , .B1( n588 ) );
  NAND2_X1 U82 (.A2( ld ) , .ZN( n80 ) , .A1( text_in[39] ) );
  XNOR2_X1 U823 (.ZN( n591 ) , .B( sa30_sr_1 ) , .A( w0_9 ) );
  XOR2_X1 U824 (.A( n211 ) , .Z( n587 ) , .B( w0_9 ) );
  OAI21_X1 U83 (.B1( ld ) , .ZN( n1018 ) , .B2( n81 ) , .A( n82 ) );
  NAND2_X1 U84 (.A2( ld ) , .ZN( n82 ) , .A1( text_in[40] ) );
  OAI22_X1 U841 (.ZN( N232 ) , .A1( n1109 ) , .B2( n1217 ) , .A2( n601 ) , .B1( n602 ) );
  XOR2_X1 U844 (.Z( n605 ) , .B( sa30_sr_5 ) , .A( w0_6 ) );
  XNOR2_X1 U845 (.B( n470 ) , .ZN( n603 ) , .A( sa00_sr_5 ) );
  XOR2_X1 U846 (.Z( n470 ) , .A( sa00_sr_6 ) , .B( sa10_sr_6 ) );
  XOR2_X1 U847 (.A( n205 ) , .Z( n601 ) , .B( w0_6 ) );
  OAI21_X1 U85 (.B1( ld ) , .ZN( n1019 ) , .B2( n83 ) , .A( n84 ) );
  NAND2_X1 U86 (.A2( ld ) , .ZN( n84 ) , .A1( text_in[41] ) );
  NOR4_X1 U866 (.ZN( N23 ) , .A3( ld ) , .A2( n1108 ) , .A4( n260 ) , .A1( n977 ) );
  NAND2_X1 U867 (.A1( n1106 ) , .A2( n1107 ) , .ZN( n260 ) );
  OAI21_X1 U87 (.B1( ld ) , .ZN( n1020 ) , .B2( n85 ) , .A( n86 ) );
  NAND2_X1 U88 (.A2( ld ) , .ZN( n86 ) , .A1( text_in[42] ) );
  OAI21_X1 U89 (.B1( ld ) , .ZN( n1021 ) , .B2( n87 ) , .A( n88 ) );
  OAI22_X1 U894 (.ZN( N226 ) , .A1( n1109 ) , .B2( n1217 ) , .A2( n635 ) , .B1( n636 ) );
  OAI21_X1 U9 (.B1( ld ) , .B2( n7 ) , .A( n8 ) , .ZN( n981 ) );
  NAND2_X1 U90 (.A2( ld ) , .ZN( n88 ) , .A1( text_in[43] ) );
  XOR2_X1 U900 (.A( n193 ) , .Z( n635 ) , .B( w0_0 ) );
  OAI22_X1 U902 (.ZN( N217 ) , .A1( n1109 ) , .B2( n1218 ) , .A2( n639 ) , .B1( n640 ) );
  XOR2_X1 U904 (.Z( n642 ) , .A( n643 ) , .B( n644 ) );
  INV_X1 U906 (.ZN( n645 ) , .A( sa11_sr_7 ) );
  XOR2_X1 U907 (.A( n191 ) , .Z( n639 ) , .B( w1_31 ) );
  OAI22_X1 U909 (.ZN( N216 ) , .A1( n1109 ) , .B2( n1218 ) , .A2( n646 ) , .B1( n647 ) );
  OAI21_X1 U91 (.B1( ld ) , .ZN( n1022 ) , .B2( n89 ) , .A( n90 ) );
  XOR2_X1 U911 (.Z( n649 ) , .A( n650 ) , .B( n651 ) );
  XOR2_X1 U913 (.A( n189 ) , .Z( n646 ) , .B( w1_30 ) );
  OAI22_X1 U915 (.ZN( N215 ) , .A1( n1109 ) , .B2( n1218 ) , .A2( n652 ) , .B1( n653 ) );
  XOR2_X1 U917 (.Z( n655 ) , .A( n656 ) , .B( n657 ) );
  XOR2_X1 U919 (.A( n187 ) , .Z( n652 ) , .B( w1_29 ) );
  NAND2_X1 U92 (.A2( ld ) , .ZN( n90 ) , .A1( text_in[44] ) );
  OAI22_X1 U921 (.ZN( N214 ) , .A1( n1109 ) , .B2( n1218 ) , .A2( n658 ) , .B1( n659 ) );
  XOR2_X1 U922 (.Z( n659 ) , .A( n660 ) , .B( n661 ) );
  XOR2_X1 U923 (.Z( n661 ) , .A( n662 ) , .B( n663 ) );
  XOR2_X1 U924 (.Z( n660 ) , .A( n664 ) , .B( n665 ) );
  XNOR2_X1 U925 (.ZN( n664 ) , .B( sa11_sr_4 ) , .A( w1_28 ) );
  XOR2_X1 U926 (.A( n185 ) , .Z( n658 ) , .B( w1_28 ) );
  OAI22_X1 U928 (.ZN( N213 ) , .A1( n1213 ) , .B2( n1218 ) , .A2( n666 ) , .B1( n667 ) );
  OAI21_X1 U93 (.B1( ld ) , .ZN( n1023 ) , .B2( n91 ) , .A( n92 ) );
  XOR2_X1 U930 (.Z( n669 ) , .A( n670 ) , .B( n671 ) );
  XNOR2_X1 U932 (.ZN( n672 ) , .B( sa11_sr_3 ) , .A( w1_27 ) );
  XOR2_X1 U933 (.A( n183 ) , .Z( n666 ) , .B( w1_27 ) );
  OAI22_X1 U935 (.ZN( N212 ) , .A1( n1214 ) , .B2( n1218 ) , .A2( n673 ) , .B1( n674 ) );
  XOR2_X1 U937 (.Z( n676 ) , .A( n677 ) , .B( n678 ) );
  XOR2_X1 U939 (.A( n181 ) , .Z( n673 ) , .B( w1_26 ) );
  NAND2_X1 U94 (.A2( ld ) , .ZN( n92 ) , .A1( text_in[45] ) );
  OAI22_X1 U941 (.ZN( N211 ) , .A1( n1214 ) , .B2( n1218 ) , .A2( n679 ) , .B1( n680 ) );
  XOR2_X1 U943 (.Z( n682 ) , .A( n683 ) , .B( n684 ) );
  XNOR2_X1 U945 (.ZN( n685 ) , .B( sa11_sr_1 ) , .A( w1_25 ) );
  XOR2_X1 U946 (.A( n179 ) , .Z( n679 ) , .B( w1_25 ) );
  OAI22_X1 U948 (.ZN( N210 ) , .A1( n1109 ) , .B2( n1219 ) , .A2( n686 ) , .B1( n687 ) );
  OAI21_X1 U95 (.B1( ld ) , .ZN( n1024 ) , .B2( n93 ) , .A( n94 ) );
  XOR2_X1 U950 (.A( n665 ) , .Z( n689 ) , .B( n690 ) );
  XOR2_X1 U952 (.A( n177 ) , .Z( n686 ) , .B( w1_24 ) );
  OAI22_X1 U954 (.ZN( N201 ) , .A1( n1214 ) , .B2( n1217 ) , .A2( n691 ) , .B1( n692 ) );
  XOR2_X1 U955 (.Z( n692 ) , .A( n693 ) , .B( n694 ) );
  XOR2_X1 U956 (.B( n643 ) , .Z( n694 ) , .A( sa01_sr_7 ) );
  XOR2_X1 U959 (.A( n175 ) , .Z( n691 ) , .B( w1_23 ) );
  NAND2_X1 U96 (.A2( ld ) , .ZN( n94 ) , .A1( text_in[46] ) );
  OAI22_X1 U961 (.ZN( N200 ) , .A1( n1212 ) , .B2( n1219 ) , .A2( n696 ) , .B1( n697 ) );
  XOR2_X1 U964 (.Z( n700 ) , .B( sa21_sr_5 ) , .A( w1_22 ) );
  XOR2_X1 U967 (.A( n173 ) , .Z( n696 ) , .B( w1_22 ) );
  OAI22_X1 U969 (.ZN( N199 ) , .A1( n1215 ) , .B2( n1218 ) , .A2( n702 ) , .B1( n703 ) );
  OAI21_X1 U97 (.B1( ld ) , .ZN( n1025 ) , .B2( n95 ) , .A( n96 ) );
  XOR2_X1 U970 (.Z( n703 ) , .A( n704 ) , .B( n705 ) );
  XOR2_X1 U971 (.Z( n705 ) , .B( n706 ) , .A( sa11_sr_4 ) );
  XOR2_X1 U972 (.Z( n706 ) , .B( sa21_sr_4 ) , .A( w1_21 ) );
  XNOR2_X1 U973 (.B( n656 ) , .ZN( n704 ) , .A( sa01_sr_5 ) );
  XOR2_X1 U974 (.A( n171 ) , .Z( n702 ) , .B( w1_21 ) );
  OAI22_X1 U976 (.ZN( N198 ) , .A1( n1216 ) , .B2( n1217 ) , .A2( n707 ) , .B1( n708 ) );
  XOR2_X1 U977 (.Z( n708 ) , .A( n709 ) , .B( n710 ) );
  XOR2_X1 U978 (.Z( n710 ) , .B( n711 ) , .A( sa11_sr_3 ) );
  XOR2_X1 U979 (.Z( n711 ) , .B( sa21_sr_3 ) , .A( w1_20 ) );
  NAND2_X1 U98 (.A2( ld ) , .ZN( n96 ) , .A1( text_in[47] ) );
  XOR2_X1 U980 (.Z( n709 ) , .A( n712 ) , .B( n713 ) );
  XNOR2_X1 U981 (.B( n663 ) , .ZN( n712 ) , .A( sa01_sr_4 ) );
  XOR2_X1 U982 (.A( n169 ) , .Z( n707 ) , .B( w1_20 ) );
  OAI22_X1 U984 (.ZN( N197 ) , .A1( n1109 ) , .B2( n1220 ) , .A2( n714 ) , .B1( n715 ) );
  XOR2_X1 U987 (.Z( n718 ) , .B( sa21_sr_2 ) , .A( w1_19 ) );
  XOR2_X1 U988 (.B( n713 ) , .Z( n716 ) , .A( n719 ) );
  XNOR2_X1 U989 (.B( n670 ) , .ZN( n719 ) , .A( sa01_sr_3 ) );
  OAI21_X1 U99 (.B1( ld ) , .ZN( n1026 ) , .B2( n97 ) , .A( n98 ) );
  XOR2_X1 U990 (.A( n167 ) , .Z( n714 ) , .B( w1_19 ) );
  OAI22_X1 U992 (.ZN( N196 ) , .A1( n1212 ) , .B2( n1218 ) , .A2( n720 ) , .B1( n721 ) );
  XOR2_X1 U995 (.Z( n724 ) , .B( sa21_sr_1 ) , .A( w1_18 ) );
  XNOR2_X1 U996 (.B( n677 ) , .ZN( n722 ) , .A( sa01_sr_2 ) );
  XOR2_X1 U997 (.A( n165 ) , .Z( n720 ) , .B( w1_18 ) );
  OAI22_X1 U999 (.ZN( N195 ) , .A1( n1215 ) , .B2( n1221 ) , .A2( n725 ) , .B1( n726 ) );
  DFF_X1 dcnt_reg_0 (.CK( clk ) , .QN( n1108 ) , .D( n1113 ) , .Q( n261 ) );
  DFF_X1 dcnt_reg_1 (.CK( clk ) , .D( n1110 ) , .Q( n977 ) );
  DFF_X1 dcnt_reg_2 (.CK( clk ) , .QN( n1107 ) , .D( n1111 ) , .Q( n267 ) );
  DFF_X1 dcnt_reg_3 (.CK( clk ) , .QN( n1106 ) , .D( n1112 ) );
  DFF_X1 done_reg (.D( N23 ) , .CK( clk ) , .Q( done ) );
  DFF_X1 ld_r_reg (.CK( clk ) , .D( ld ) , .QN( n1109 ) , .Q( n1114 ) );
  DFF_X1 sa00_reg_0 (.D( N274 ) , .CK( clk ) , .Q( sa00_0 ) );
  DFF_X1 sa00_reg_1 (.D( N275 ) , .CK( clk ) , .Q( sa00_1 ) );
  DFF_X1 sa00_reg_2 (.D( N276 ) , .CK( clk ) , .Q( sa00_2 ) );
  DFF_X1 sa00_reg_3 (.D( N277 ) , .CK( clk ) , .Q( sa00_3 ) );
  DFF_X1 sa00_reg_4 (.D( N278 ) , .CK( clk ) , .Q( sa00_4 ) );
  DFF_X1 sa00_reg_5 (.D( N279 ) , .CK( clk ) , .Q( sa00_5 ) );
  DFF_X1 sa00_reg_6 (.D( N280 ) , .CK( clk ) , .Q( sa00_6 ) );
  DFF_X1 sa00_reg_7 (.D( N281 ) , .CK( clk ) , .Q( sa00_7 ) );
  DFF_X1 sa01_reg_0 (.D( N210 ) , .CK( clk ) , .Q( sa01_0 ) );
  DFF_X1 sa01_reg_1 (.D( N211 ) , .CK( clk ) , .Q( sa01_1 ) );
  DFF_X1 sa01_reg_2 (.D( N212 ) , .CK( clk ) , .Q( sa01_2 ) );
  DFF_X1 sa01_reg_3 (.D( N213 ) , .CK( clk ) , .Q( sa01_3 ) );
  DFF_X1 sa01_reg_4 (.D( N214 ) , .CK( clk ) , .Q( sa01_4 ) );
  DFF_X1 sa01_reg_5 (.D( N215 ) , .CK( clk ) , .Q( sa01_5 ) );
  DFF_X1 sa01_reg_6 (.D( N216 ) , .CK( clk ) , .Q( sa01_6 ) );
  DFF_X1 sa01_reg_7 (.D( N217 ) , .CK( clk ) , .Q( sa01_7 ) );
  DFF_X1 sa02_reg_0 (.D( N146 ) , .CK( clk ) , .Q( sa02_0 ) );
  DFF_X1 sa02_reg_1 (.D( N147 ) , .CK( clk ) , .Q( sa02_1 ) );
  DFF_X1 sa02_reg_2 (.D( N148 ) , .CK( clk ) , .Q( sa02_2 ) );
  DFF_X1 sa02_reg_3 (.D( N149 ) , .CK( clk ) , .Q( sa02_3 ) );
  DFF_X1 sa02_reg_4 (.D( N150 ) , .CK( clk ) , .Q( sa02_4 ) );
  DFF_X1 sa02_reg_5 (.D( N151 ) , .CK( clk ) , .Q( sa02_5 ) );
  DFF_X1 sa02_reg_6 (.D( N152 ) , .CK( clk ) , .Q( sa02_6 ) );
  DFF_X1 sa02_reg_7 (.D( N153 ) , .CK( clk ) , .Q( sa02_7 ) );
  DFF_X1 sa03_reg_0 (.D( N82 ) , .CK( clk ) , .Q( sa03_0 ) );
  DFF_X1 sa03_reg_1 (.D( N83 ) , .CK( clk ) , .Q( sa03_1 ) );
  DFF_X1 sa03_reg_2 (.D( N84 ) , .CK( clk ) , .Q( sa03_2 ) );
  DFF_X1 sa03_reg_3 (.D( N85 ) , .CK( clk ) , .Q( sa03_3 ) );
  DFF_X1 sa03_reg_4 (.D( N86 ) , .CK( clk ) , .Q( sa03_4 ) );
  DFF_X1 sa03_reg_5 (.D( N87 ) , .CK( clk ) , .Q( sa03_5 ) );
  DFF_X1 sa03_reg_6 (.D( N88 ) , .CK( clk ) , .Q( sa03_6 ) );
  DFF_X1 sa03_reg_7 (.D( N89 ) , .CK( clk ) , .Q( sa03_7 ) );
  DFF_X1 sa10_reg_0 (.D( N258 ) , .CK( clk ) , .Q( sa10_0 ) );
  DFF_X1 sa10_reg_1 (.D( N259 ) , .CK( clk ) , .Q( sa10_1 ) );
  DFF_X1 sa10_reg_2 (.D( N260 ) , .CK( clk ) , .Q( sa10_2 ) );
  DFF_X1 sa10_reg_3 (.D( N261 ) , .CK( clk ) , .Q( sa10_3 ) );
  DFF_X1 sa10_reg_4 (.D( N262 ) , .CK( clk ) , .Q( sa10_4 ) );
  DFF_X1 sa10_reg_5 (.D( N263 ) , .CK( clk ) , .Q( sa10_5 ) );
  DFF_X1 sa10_reg_6 (.D( N264 ) , .CK( clk ) , .Q( sa10_6 ) );
  DFF_X1 sa10_reg_7 (.D( N265 ) , .CK( clk ) , .Q( sa10_7 ) );
  DFF_X1 sa11_reg_0 (.D( N194 ) , .CK( clk ) , .Q( sa11_0 ) );
  DFF_X1 sa11_reg_1 (.D( N195 ) , .CK( clk ) , .Q( sa11_1 ) );
  DFF_X1 sa11_reg_2 (.D( N196 ) , .CK( clk ) , .Q( sa11_2 ) );
  DFF_X1 sa11_reg_3 (.D( N197 ) , .CK( clk ) , .Q( sa11_3 ) );
  DFF_X1 sa11_reg_4 (.D( N198 ) , .CK( clk ) , .Q( sa11_4 ) );
  DFF_X1 sa11_reg_5 (.D( N199 ) , .CK( clk ) , .Q( sa11_5 ) );
  DFF_X1 sa11_reg_6 (.D( N200 ) , .CK( clk ) , .Q( sa11_6 ) );
  DFF_X1 sa11_reg_7 (.D( N201 ) , .CK( clk ) , .Q( sa11_7 ) );
  DFF_X1 sa12_reg_0 (.D( N130 ) , .CK( clk ) , .Q( sa12_0 ) );
  DFF_X1 sa12_reg_1 (.D( N131 ) , .CK( clk ) , .Q( sa12_1 ) );
  DFF_X1 sa12_reg_2 (.D( N132 ) , .CK( clk ) , .Q( sa12_2 ) );
  DFF_X1 sa12_reg_3 (.D( N133 ) , .CK( clk ) , .Q( sa12_3 ) );
  DFF_X1 sa12_reg_4 (.D( N134 ) , .CK( clk ) , .Q( sa12_4 ) );
  DFF_X1 sa12_reg_5 (.D( N135 ) , .CK( clk ) , .Q( sa12_5 ) );
  DFF_X1 sa12_reg_6 (.D( N136 ) , .CK( clk ) , .Q( sa12_6 ) );
  DFF_X1 sa12_reg_7 (.D( N137 ) , .CK( clk ) , .Q( sa12_7 ) );
  DFF_X1 sa13_reg_0 (.D( N66 ) , .CK( clk ) , .Q( sa13_0 ) );
  DFF_X1 sa13_reg_1 (.D( N67 ) , .CK( clk ) , .Q( sa13_1 ) );
  DFF_X1 sa13_reg_2 (.D( N68 ) , .CK( clk ) , .Q( sa13_2 ) );
  DFF_X1 sa13_reg_3 (.D( N69 ) , .CK( clk ) , .Q( sa13_3 ) );
  DFF_X1 sa13_reg_4 (.D( N70 ) , .CK( clk ) , .Q( sa13_4 ) );
  DFF_X1 sa13_reg_5 (.D( N71 ) , .CK( clk ) , .Q( sa13_5 ) );
  DFF_X1 sa13_reg_6 (.D( N72 ) , .CK( clk ) , .Q( sa13_6 ) );
  DFF_X1 sa13_reg_7 (.D( N73 ) , .CK( clk ) , .Q( sa13_7 ) );
  DFF_X1 sa20_reg_0 (.D( N242 ) , .CK( clk ) , .Q( sa20_0 ) );
  DFF_X1 sa20_reg_1 (.D( N243 ) , .CK( clk ) , .Q( sa20_1 ) );
  DFF_X1 sa20_reg_2 (.D( N244 ) , .CK( clk ) , .Q( sa20_2 ) );
  DFF_X1 sa20_reg_3 (.D( N245 ) , .CK( clk ) , .Q( sa20_3 ) );
  DFF_X1 sa20_reg_4 (.D( N246 ) , .CK( clk ) , .Q( sa20_4 ) );
  DFF_X1 sa20_reg_5 (.D( N247 ) , .CK( clk ) , .Q( sa20_5 ) );
  DFF_X1 sa20_reg_6 (.D( N248 ) , .CK( clk ) , .Q( sa20_6 ) );
  DFF_X1 sa20_reg_7 (.D( N249 ) , .CK( clk ) , .Q( sa20_7 ) );
  DFF_X1 sa21_reg_0 (.D( N178 ) , .CK( clk ) , .Q( sa21_0 ) );
  DFF_X1 sa21_reg_1 (.D( N179 ) , .CK( clk ) , .Q( sa21_1 ) );
  DFF_X1 sa21_reg_2 (.D( N180 ) , .CK( clk ) , .Q( sa21_2 ) );
  DFF_X1 sa21_reg_3 (.D( N181 ) , .CK( clk ) , .Q( sa21_3 ) );
  DFF_X1 sa21_reg_4 (.D( N182 ) , .CK( clk ) , .Q( sa21_4 ) );
  DFF_X1 sa21_reg_5 (.D( N183 ) , .CK( clk ) , .Q( sa21_5 ) );
  DFF_X1 sa21_reg_6 (.D( N184 ) , .CK( clk ) , .Q( sa21_6 ) );
  DFF_X1 sa21_reg_7 (.D( N185 ) , .CK( clk ) , .Q( sa21_7 ) );
  DFF_X1 sa22_reg_0 (.D( N114 ) , .CK( clk ) , .Q( sa22_0 ) );
  DFF_X1 sa22_reg_1 (.D( N115 ) , .CK( clk ) , .Q( sa22_1 ) );
  DFF_X1 sa22_reg_2 (.D( N116 ) , .CK( clk ) , .Q( sa22_2 ) );
  DFF_X1 sa22_reg_3 (.D( N117 ) , .CK( clk ) , .Q( sa22_3 ) );
  DFF_X1 sa22_reg_4 (.D( N118 ) , .CK( clk ) , .Q( sa22_4 ) );
  DFF_X1 sa22_reg_5 (.D( N119 ) , .CK( clk ) , .Q( sa22_5 ) );
  DFF_X1 sa22_reg_6 (.D( N120 ) , .CK( clk ) , .Q( sa22_6 ) );
  DFF_X1 sa22_reg_7 (.D( N121 ) , .CK( clk ) , .Q( sa22_7 ) );
  DFF_X1 sa23_reg_0 (.D( N50 ) , .CK( clk ) , .Q( sa23_0 ) );
  DFF_X1 sa23_reg_1 (.D( N51 ) , .CK( clk ) , .Q( sa23_1 ) );
  DFF_X1 sa23_reg_2 (.D( N52 ) , .CK( clk ) , .Q( sa23_2 ) );
  DFF_X1 sa23_reg_3 (.D( N53 ) , .CK( clk ) , .Q( sa23_3 ) );
  DFF_X1 sa23_reg_4 (.D( N54 ) , .CK( clk ) , .Q( sa23_4 ) );
  DFF_X1 sa23_reg_5 (.D( N55 ) , .CK( clk ) , .Q( sa23_5 ) );
  DFF_X1 sa23_reg_6 (.D( N56 ) , .CK( clk ) , .Q( sa23_6 ) );
  DFF_X1 sa23_reg_7 (.D( N57 ) , .CK( clk ) , .Q( sa23_7 ) );
  DFF_X1 sa30_reg_0 (.D( N226 ) , .CK( clk ) , .Q( sa30_0 ) );
  DFF_X1 sa30_reg_1 (.D( N227 ) , .CK( clk ) , .Q( sa30_1 ) );
  DFF_X1 sa30_reg_2 (.D( N228 ) , .CK( clk ) , .Q( sa30_2 ) );
  DFF_X1 sa30_reg_3 (.D( N229 ) , .CK( clk ) , .Q( sa30_3 ) );
  DFF_X1 sa30_reg_4 (.D( N230 ) , .CK( clk ) , .Q( sa30_4 ) );
  DFF_X1 sa30_reg_5 (.D( N231 ) , .CK( clk ) , .Q( sa30_5 ) );
  DFF_X1 sa30_reg_6 (.D( N232 ) , .CK( clk ) , .Q( sa30_6 ) );
  DFF_X1 sa30_reg_7 (.D( N233 ) , .CK( clk ) , .Q( sa30_7 ) );
  DFF_X1 sa31_reg_0 (.D( N162 ) , .CK( clk ) , .Q( sa31_0 ) );
  DFF_X1 sa31_reg_1 (.D( N163 ) , .CK( clk ) , .Q( sa31_1 ) );
  DFF_X1 sa31_reg_2 (.D( N164 ) , .CK( clk ) , .Q( sa31_2 ) );
  DFF_X1 sa31_reg_3 (.D( N165 ) , .CK( clk ) , .Q( sa31_3 ) );
  DFF_X1 sa31_reg_4 (.D( N166 ) , .CK( clk ) , .Q( sa31_4 ) );
  DFF_X1 sa31_reg_5 (.D( N167 ) , .CK( clk ) , .Q( sa31_5 ) );
  DFF_X1 sa31_reg_6 (.D( N168 ) , .CK( clk ) , .Q( sa31_6 ) );
  DFF_X1 sa31_reg_7 (.D( N169 ) , .CK( clk ) , .Q( sa31_7 ) );
  DFF_X1 sa32_reg_0 (.D( N98 ) , .CK( clk ) , .Q( sa32_0 ) );
  DFF_X1 sa32_reg_1 (.D( N99 ) , .CK( clk ) , .Q( sa32_1 ) );
  DFF_X1 sa32_reg_2 (.D( N100 ) , .CK( clk ) , .Q( sa32_2 ) );
  DFF_X1 sa32_reg_3 (.D( N101 ) , .CK( clk ) , .Q( sa32_3 ) );
  DFF_X1 sa32_reg_4 (.D( N102 ) , .CK( clk ) , .Q( sa32_4 ) );
  DFF_X1 sa32_reg_5 (.D( N103 ) , .CK( clk ) , .Q( sa32_5 ) );
  DFF_X1 sa32_reg_6 (.D( N104 ) , .CK( clk ) , .Q( sa32_6 ) );
  DFF_X1 sa32_reg_7 (.D( N105 ) , .CK( clk ) , .Q( sa32_7 ) );
  DFF_X1 sa33_reg_0 (.D( N34 ) , .CK( clk ) , .Q( sa33_0 ) );
  DFF_X1 sa33_reg_1 (.D( N35 ) , .CK( clk ) , .Q( sa33_1 ) );
  DFF_X1 sa33_reg_2 (.D( N36 ) , .CK( clk ) , .Q( sa33_2 ) );
  DFF_X1 sa33_reg_3 (.D( N37 ) , .CK( clk ) , .Q( sa33_3 ) );
  DFF_X1 sa33_reg_4 (.D( N38 ) , .CK( clk ) , .Q( sa33_4 ) );
  DFF_X1 sa33_reg_5 (.D( N39 ) , .CK( clk ) , .Q( sa33_5 ) );
  DFF_X1 sa33_reg_6 (.D( N40 ) , .CK( clk ) , .Q( sa33_6 ) );
  DFF_X1 sa33_reg_7 (.D( N41 ) , .CK( clk ) , .Q( sa33_7 ) );
  DFF_X1 text_in_r_reg_0 (.CK( clk ) , .QN( n1 ) , .D( n978 ) );
  DFF_X1 text_in_r_reg_1 (.CK( clk ) , .QN( n3 ) , .D( n979 ) );
  DFF_X1 text_in_r_reg_10 (.CK( clk ) , .QN( n21 ) , .D( n988 ) );
  DFF_X1 text_in_r_reg_100 (.CK( clk ) , .D( n1078 ) , .QN( n201 ) );
  DFF_X1 text_in_r_reg_101 (.CK( clk ) , .D( n1079 ) , .QN( n203 ) );
  DFF_X1 text_in_r_reg_102 (.CK( clk ) , .D( n1080 ) , .QN( n205 ) );
  DFF_X1 text_in_r_reg_103 (.CK( clk ) , .D( n1081 ) , .QN( n207 ) );
  DFF_X1 text_in_r_reg_104 (.CK( clk ) , .D( n1082 ) , .QN( n209 ) );
  DFF_X1 text_in_r_reg_105 (.CK( clk ) , .D( n1083 ) , .QN( n211 ) );
  DFF_X1 text_in_r_reg_106 (.CK( clk ) , .D( n1084 ) , .QN( n213 ) );
  DFF_X1 text_in_r_reg_107 (.CK( clk ) , .D( n1085 ) , .QN( n215 ) );
  DFF_X1 text_in_r_reg_108 (.CK( clk ) , .D( n1086 ) , .QN( n217 ) );
  DFF_X1 text_in_r_reg_109 (.CK( clk ) , .D( n1087 ) , .QN( n219 ) );
  DFF_X1 text_in_r_reg_11 (.CK( clk ) , .QN( n23 ) , .D( n989 ) );
  DFF_X1 text_in_r_reg_110 (.CK( clk ) , .D( n1088 ) , .QN( n221 ) );
  DFF_X1 text_in_r_reg_111 (.CK( clk ) , .D( n1089 ) , .QN( n223 ) );
  DFF_X1 text_in_r_reg_112 (.CK( clk ) , .D( n1090 ) , .QN( n225 ) );
  DFF_X1 text_in_r_reg_113 (.CK( clk ) , .D( n1091 ) , .QN( n227 ) );
  DFF_X1 text_in_r_reg_114 (.CK( clk ) , .D( n1092 ) , .QN( n229 ) );
  DFF_X1 text_in_r_reg_115 (.CK( clk ) , .D( n1093 ) , .QN( n231 ) );
  DFF_X1 text_in_r_reg_116 (.CK( clk ) , .D( n1094 ) , .QN( n233 ) );
  DFF_X1 text_in_r_reg_117 (.CK( clk ) , .D( n1095 ) , .QN( n235 ) );
  DFF_X1 text_in_r_reg_118 (.CK( clk ) , .D( n1096 ) , .QN( n237 ) );
  DFF_X1 text_in_r_reg_119 (.CK( clk ) , .D( n1097 ) , .QN( n239 ) );
  DFF_X1 text_in_r_reg_12 (.CK( clk ) , .QN( n25 ) , .D( n990 ) );
  DFF_X1 text_in_r_reg_120 (.CK( clk ) , .D( n1098 ) , .QN( n241 ) );
  DFF_X1 text_in_r_reg_121 (.CK( clk ) , .D( n1099 ) , .QN( n243 ) );
  DFF_X1 text_in_r_reg_122 (.CK( clk ) , .D( n1100 ) , .QN( n245 ) );
  DFF_X1 text_in_r_reg_123 (.CK( clk ) , .D( n1101 ) , .QN( n247 ) );
  DFF_X1 text_in_r_reg_124 (.CK( clk ) , .D( n1102 ) , .QN( n249 ) );
  DFF_X1 text_in_r_reg_125 (.CK( clk ) , .D( n1103 ) , .QN( n251 ) );
  DFF_X1 text_in_r_reg_126 (.CK( clk ) , .D( n1104 ) , .QN( n253 ) );
  DFF_X1 text_in_r_reg_127 (.CK( clk ) , .D( n1105 ) , .QN( n255 ) );
  DFF_X1 text_in_r_reg_13 (.CK( clk ) , .QN( n27 ) , .D( n991 ) );
  DFF_X1 text_in_r_reg_14 (.CK( clk ) , .QN( n29 ) , .D( n992 ) );
  DFF_X1 text_in_r_reg_15 (.CK( clk ) , .QN( n31 ) , .D( n993 ) );
  DFF_X1 text_in_r_reg_16 (.CK( clk ) , .QN( n33 ) , .D( n994 ) );
  DFF_X1 text_in_r_reg_17 (.CK( clk ) , .QN( n35 ) , .D( n995 ) );
  DFF_X1 text_in_r_reg_18 (.CK( clk ) , .QN( n37 ) , .D( n996 ) );
  DFF_X1 text_in_r_reg_19 (.CK( clk ) , .QN( n39 ) , .D( n997 ) );
  DFF_X1 text_in_r_reg_2 (.CK( clk ) , .QN( n5 ) , .D( n980 ) );
  DFF_X1 text_in_r_reg_20 (.CK( clk ) , .QN( n41 ) , .D( n998 ) );
  DFF_X1 text_in_r_reg_21 (.CK( clk ) , .QN( n43 ) , .D( n999 ) );
  DFF_X1 text_in_r_reg_22 (.CK( clk ) , .D( n1000 ) , .QN( n45 ) );
  DFF_X1 text_in_r_reg_23 (.CK( clk ) , .D( n1001 ) , .QN( n47 ) );
  DFF_X1 text_in_r_reg_24 (.CK( clk ) , .D( n1002 ) , .QN( n49 ) );
  DFF_X1 text_in_r_reg_25 (.CK( clk ) , .D( n1003 ) , .QN( n51 ) );
  DFF_X1 text_in_r_reg_26 (.CK( clk ) , .D( n1004 ) , .QN( n53 ) );
  DFF_X1 text_in_r_reg_27 (.CK( clk ) , .D( n1005 ) , .QN( n55 ) );
  DFF_X1 text_in_r_reg_28 (.CK( clk ) , .D( n1006 ) , .QN( n57 ) );
  DFF_X1 text_in_r_reg_29 (.CK( clk ) , .D( n1007 ) , .QN( n59 ) );
  DFF_X1 text_in_r_reg_3 (.CK( clk ) , .QN( n7 ) , .D( n981 ) );
  DFF_X1 text_in_r_reg_30 (.CK( clk ) , .D( n1008 ) , .QN( n61 ) );
  DFF_X1 text_in_r_reg_31 (.CK( clk ) , .D( n1009 ) , .QN( n63 ) );
  DFF_X1 text_in_r_reg_32 (.CK( clk ) , .D( n1010 ) , .QN( n65 ) );
  DFF_X1 text_in_r_reg_33 (.CK( clk ) , .D( n1011 ) , .QN( n67 ) );
  DFF_X1 text_in_r_reg_34 (.CK( clk ) , .D( n1012 ) , .QN( n69 ) );
  DFF_X1 text_in_r_reg_35 (.CK( clk ) , .D( n1013 ) , .QN( n71 ) );
  DFF_X1 text_in_r_reg_36 (.CK( clk ) , .D( n1014 ) , .QN( n73 ) );
  DFF_X1 text_in_r_reg_37 (.CK( clk ) , .D( n1015 ) , .QN( n75 ) );
  DFF_X1 text_in_r_reg_38 (.CK( clk ) , .D( n1016 ) , .QN( n77 ) );
  DFF_X1 text_in_r_reg_39 (.CK( clk ) , .D( n1017 ) , .QN( n79 ) );
  DFF_X1 text_in_r_reg_4 (.CK( clk ) , .QN( n9 ) , .D( n982 ) );
  DFF_X1 text_in_r_reg_40 (.CK( clk ) , .D( n1018 ) , .QN( n81 ) );
  DFF_X1 text_in_r_reg_41 (.CK( clk ) , .D( n1019 ) , .QN( n83 ) );
  DFF_X1 text_in_r_reg_42 (.CK( clk ) , .D( n1020 ) , .QN( n85 ) );
  DFF_X1 text_in_r_reg_43 (.CK( clk ) , .D( n1021 ) , .QN( n87 ) );
  DFF_X1 text_in_r_reg_44 (.CK( clk ) , .D( n1022 ) , .QN( n89 ) );
  DFF_X1 text_in_r_reg_45 (.CK( clk ) , .D( n1023 ) , .QN( n91 ) );
  DFF_X1 text_in_r_reg_46 (.CK( clk ) , .D( n1024 ) , .QN( n93 ) );
  DFF_X1 text_in_r_reg_47 (.CK( clk ) , .D( n1025 ) , .QN( n95 ) );
  DFF_X1 text_in_r_reg_48 (.CK( clk ) , .D( n1026 ) , .QN( n97 ) );
  DFF_X1 text_in_r_reg_49 (.CK( clk ) , .D( n1027 ) , .QN( n99 ) );
  DFF_X1 text_in_r_reg_5 (.CK( clk ) , .QN( n11 ) , .D( n983 ) );
  DFF_X1 text_in_r_reg_50 (.CK( clk ) , .QN( n101 ) , .D( n1028 ) );
  DFF_X1 text_in_r_reg_51 (.CK( clk ) , .D( n1029 ) , .QN( n103 ) );
  DFF_X1 text_in_r_reg_52 (.CK( clk ) , .D( n1030 ) , .QN( n105 ) );
  DFF_X1 text_in_r_reg_53 (.CK( clk ) , .D( n1031 ) , .QN( n107 ) );
  DFF_X1 text_in_r_reg_54 (.CK( clk ) , .D( n1032 ) , .QN( n109 ) );
  DFF_X1 text_in_r_reg_55 (.CK( clk ) , .D( n1033 ) , .QN( n111 ) );
  DFF_X1 text_in_r_reg_56 (.CK( clk ) , .D( n1034 ) , .QN( n113 ) );
  DFF_X1 text_in_r_reg_57 (.CK( clk ) , .D( n1035 ) , .QN( n115 ) );
  DFF_X1 text_in_r_reg_58 (.CK( clk ) , .D( n1036 ) , .QN( n117 ) );
  DFF_X1 text_in_r_reg_59 (.CK( clk ) , .D( n1037 ) , .QN( n119 ) );
  DFF_X1 text_in_r_reg_6 (.CK( clk ) , .QN( n13 ) , .D( n984 ) );
  DFF_X1 text_in_r_reg_60 (.CK( clk ) , .D( n1038 ) , .QN( n121 ) );
  DFF_X1 text_in_r_reg_61 (.CK( clk ) , .D( n1039 ) , .QN( n123 ) );
  DFF_X1 text_in_r_reg_62 (.CK( clk ) , .D( n1040 ) , .QN( n125 ) );
  DFF_X1 text_in_r_reg_63 (.CK( clk ) , .D( n1041 ) , .QN( n127 ) );
  DFF_X1 text_in_r_reg_64 (.CK( clk ) , .D( n1042 ) , .QN( n129 ) );
  DFF_X1 text_in_r_reg_65 (.CK( clk ) , .D( n1043 ) , .QN( n131 ) );
  DFF_X1 text_in_r_reg_66 (.CK( clk ) , .D( n1044 ) , .QN( n133 ) );
  DFF_X1 text_in_r_reg_67 (.CK( clk ) , .D( n1045 ) , .QN( n135 ) );
  DFF_X1 text_in_r_reg_68 (.CK( clk ) , .D( n1046 ) , .QN( n137 ) );
  DFF_X1 text_in_r_reg_69 (.CK( clk ) , .D( n1047 ) , .QN( n139 ) );
  DFF_X1 text_in_r_reg_7 (.CK( clk ) , .QN( n15 ) , .D( n985 ) );
  DFF_X1 text_in_r_reg_70 (.CK( clk ) , .D( n1048 ) , .QN( n141 ) );
  DFF_X1 text_in_r_reg_71 (.CK( clk ) , .D( n1049 ) , .QN( n143 ) );
  DFF_X1 text_in_r_reg_72 (.CK( clk ) , .D( n1050 ) , .QN( n145 ) );
  DFF_X1 text_in_r_reg_73 (.CK( clk ) , .D( n1051 ) , .QN( n147 ) );
  DFF_X1 text_in_r_reg_74 (.CK( clk ) , .D( n1052 ) , .QN( n149 ) );
  DFF_X1 text_in_r_reg_75 (.CK( clk ) , .D( n1053 ) , .QN( n151 ) );
  DFF_X1 text_in_r_reg_76 (.CK( clk ) , .D( n1054 ) , .QN( n153 ) );
  DFF_X1 text_in_r_reg_77 (.CK( clk ) , .D( n1055 ) , .QN( n155 ) );
  DFF_X1 text_in_r_reg_78 (.CK( clk ) , .D( n1056 ) , .QN( n157 ) );
  DFF_X1 text_in_r_reg_79 (.CK( clk ) , .D( n1057 ) , .QN( n159 ) );
  DFF_X1 text_in_r_reg_8 (.CK( clk ) , .QN( n17 ) , .D( n986 ) );
  DFF_X1 text_in_r_reg_80 (.CK( clk ) , .D( n1058 ) , .QN( n161 ) );
  DFF_X1 text_in_r_reg_81 (.CK( clk ) , .D( n1059 ) , .QN( n163 ) );
  DFF_X1 text_in_r_reg_82 (.CK( clk ) , .D( n1060 ) , .QN( n165 ) );
  DFF_X1 text_in_r_reg_83 (.CK( clk ) , .D( n1061 ) , .QN( n167 ) );
  DFF_X1 text_in_r_reg_84 (.CK( clk ) , .D( n1062 ) , .QN( n169 ) );
  DFF_X1 text_in_r_reg_85 (.CK( clk ) , .D( n1063 ) , .QN( n171 ) );
  DFF_X1 text_in_r_reg_86 (.CK( clk ) , .D( n1064 ) , .QN( n173 ) );
  DFF_X1 text_in_r_reg_87 (.CK( clk ) , .D( n1065 ) , .QN( n175 ) );
  DFF_X1 text_in_r_reg_88 (.CK( clk ) , .D( n1066 ) , .QN( n177 ) );
  DFF_X1 text_in_r_reg_89 (.CK( clk ) , .D( n1067 ) , .QN( n179 ) );
  DFF_X1 text_in_r_reg_9 (.CK( clk ) , .QN( n19 ) , .D( n987 ) );
  DFF_X1 text_in_r_reg_90 (.CK( clk ) , .D( n1068 ) , .QN( n181 ) );
  DFF_X1 text_in_r_reg_91 (.CK( clk ) , .D( n1069 ) , .QN( n183 ) );
  DFF_X1 text_in_r_reg_92 (.CK( clk ) , .D( n1070 ) , .QN( n185 ) );
  DFF_X1 text_in_r_reg_93 (.CK( clk ) , .D( n1071 ) , .QN( n187 ) );
  DFF_X1 text_in_r_reg_94 (.CK( clk ) , .D( n1072 ) , .QN( n189 ) );
  DFF_X1 text_in_r_reg_95 (.CK( clk ) , .D( n1073 ) , .QN( n191 ) );
  DFF_X1 text_in_r_reg_96 (.CK( clk ) , .D( n1074 ) , .QN( n193 ) );
  DFF_X1 text_in_r_reg_97 (.CK( clk ) , .D( n1075 ) , .QN( n195 ) );
  DFF_X1 text_in_r_reg_98 (.CK( clk ) , .D( n1076 ) , .QN( n197 ) );
  DFF_X1 text_in_r_reg_99 (.CK( clk ) , .D( n1077 ) , .QN( n199 ) );
  DFF_X1 text_out_reg_0 (.D( N505 ) , .CK( clk ) , .Q( text_out[0] ) );
  DFF_X1 text_out_reg_1 (.D( N504 ) , .CK( clk ) , .Q( text_out[1] ) );
  DFF_X1 text_out_reg_10 (.D( N471 ) , .CK( clk ) , .Q( text_out[10] ) );
  DFF_X1 text_out_reg_100 (.D( N477 ) , .CK( clk ) , .Q( text_out[100] ) );
  DFF_X1 text_out_reg_101 (.D( N476 ) , .CK( clk ) , .Q( text_out[101] ) );
  DFF_X1 text_out_reg_102 (.D( N475 ) , .CK( clk ) , .Q( text_out[102] ) );
  DFF_X1 text_out_reg_103 (.D( N474 ) , .CK( clk ) , .Q( text_out[103] ) );
  DFF_X1 text_out_reg_104 (.D( N449 ) , .CK( clk ) , .Q( text_out[104] ) );
  DFF_X1 text_out_reg_105 (.D( N448 ) , .CK( clk ) , .Q( text_out[105] ) );
  DFF_X1 text_out_reg_106 (.D( N447 ) , .CK( clk ) , .Q( text_out[106] ) );
  DFF_X1 text_out_reg_107 (.D( N446 ) , .CK( clk ) , .Q( text_out[107] ) );
  DFF_X1 text_out_reg_108 (.D( N445 ) , .CK( clk ) , .Q( text_out[108] ) );
  DFF_X1 text_out_reg_109 (.D( N444 ) , .CK( clk ) , .Q( text_out[109] ) );
  DFF_X1 text_out_reg_11 (.D( N470 ) , .CK( clk ) , .Q( text_out[11] ) );
  DFF_X1 text_out_reg_110 (.D( N443 ) , .CK( clk ) , .Q( text_out[110] ) );
  DFF_X1 text_out_reg_111 (.D( N442 ) , .CK( clk ) , .Q( text_out[111] ) );
  DFF_X1 text_out_reg_112 (.D( N417 ) , .CK( clk ) , .Q( text_out[112] ) );
  DFF_X1 text_out_reg_113 (.D( N416 ) , .CK( clk ) , .Q( text_out[113] ) );
  DFF_X1 text_out_reg_114 (.D( N415 ) , .CK( clk ) , .Q( text_out[114] ) );
  DFF_X1 text_out_reg_115 (.D( N414 ) , .CK( clk ) , .Q( text_out[115] ) );
  DFF_X1 text_out_reg_116 (.D( N413 ) , .CK( clk ) , .Q( text_out[116] ) );
  DFF_X1 text_out_reg_117 (.D( N412 ) , .CK( clk ) , .Q( text_out[117] ) );
  DFF_X1 text_out_reg_118 (.D( N411 ) , .CK( clk ) , .Q( text_out[118] ) );
  DFF_X1 text_out_reg_119 (.D( N410 ) , .CK( clk ) , .Q( text_out[119] ) );
  DFF_X1 text_out_reg_12 (.D( N469 ) , .CK( clk ) , .Q( text_out[12] ) );
  DFF_X1 text_out_reg_120 (.D( N385 ) , .CK( clk ) , .Q( text_out[120] ) );
  DFF_X1 text_out_reg_121 (.D( N384 ) , .CK( clk ) , .Q( text_out[121] ) );
  DFF_X1 text_out_reg_122 (.D( N383 ) , .CK( clk ) , .Q( text_out[122] ) );
  DFF_X1 text_out_reg_123 (.D( N382 ) , .CK( clk ) , .Q( text_out[123] ) );
  DFF_X1 text_out_reg_124 (.D( N381 ) , .CK( clk ) , .Q( text_out[124] ) );
  DFF_X1 text_out_reg_125 (.D( N380 ) , .CK( clk ) , .Q( text_out[125] ) );
  DFF_X1 text_out_reg_126 (.D( N379 ) , .CK( clk ) , .Q( text_out[126] ) );
  DFF_X1 text_out_reg_127 (.D( N378 ) , .CK( clk ) , .Q( text_out[127] ) );
  DFF_X1 text_out_reg_13 (.D( N468 ) , .CK( clk ) , .Q( text_out[13] ) );
  DFF_X1 text_out_reg_14 (.D( N467 ) , .CK( clk ) , .Q( text_out[14] ) );
  DFF_X1 text_out_reg_15 (.D( N466 ) , .CK( clk ) , .Q( text_out[15] ) );
  DFF_X1 text_out_reg_16 (.D( N441 ) , .CK( clk ) , .Q( text_out[16] ) );
  DFF_X1 text_out_reg_17 (.D( N440 ) , .CK( clk ) , .Q( text_out[17] ) );
  DFF_X1 text_out_reg_18 (.D( N439 ) , .CK( clk ) , .Q( text_out[18] ) );
  DFF_X1 text_out_reg_19 (.D( N438 ) , .CK( clk ) , .Q( text_out[19] ) );
  DFF_X1 text_out_reg_2 (.D( N503 ) , .CK( clk ) , .Q( text_out[2] ) );
  DFF_X1 text_out_reg_20 (.D( N437 ) , .CK( clk ) , .Q( text_out[20] ) );
  DFF_X1 text_out_reg_21 (.D( N436 ) , .CK( clk ) , .Q( text_out[21] ) );
  DFF_X1 text_out_reg_22 (.D( N435 ) , .CK( clk ) , .Q( text_out[22] ) );
  DFF_X1 text_out_reg_23 (.D( N434 ) , .CK( clk ) , .Q( text_out[23] ) );
  DFF_X1 text_out_reg_24 (.D( N409 ) , .CK( clk ) , .Q( text_out[24] ) );
  DFF_X1 text_out_reg_25 (.D( N408 ) , .CK( clk ) , .Q( text_out[25] ) );
  DFF_X1 text_out_reg_26 (.D( N407 ) , .CK( clk ) , .Q( text_out[26] ) );
  DFF_X1 text_out_reg_27 (.D( N406 ) , .CK( clk ) , .Q( text_out[27] ) );
  DFF_X1 text_out_reg_28 (.D( N405 ) , .CK( clk ) , .Q( text_out[28] ) );
  DFF_X1 text_out_reg_29 (.D( N404 ) , .CK( clk ) , .Q( text_out[29] ) );
  DFF_X1 text_out_reg_3 (.D( N502 ) , .CK( clk ) , .Q( text_out[3] ) );
  DFF_X1 text_out_reg_30 (.D( N403 ) , .CK( clk ) , .Q( text_out[30] ) );
  DFF_X1 text_out_reg_31 (.D( N402 ) , .CK( clk ) , .Q( text_out[31] ) );
  DFF_X1 text_out_reg_32 (.D( N497 ) , .CK( clk ) , .Q( text_out[32] ) );
  DFF_X1 text_out_reg_33 (.D( N496 ) , .CK( clk ) , .Q( text_out[33] ) );
  DFF_X1 text_out_reg_34 (.D( N495 ) , .CK( clk ) , .Q( text_out[34] ) );
  DFF_X1 text_out_reg_35 (.D( N494 ) , .CK( clk ) , .Q( text_out[35] ) );
  DFF_X1 text_out_reg_36 (.D( N493 ) , .CK( clk ) , .Q( text_out[36] ) );
  DFF_X1 text_out_reg_37 (.D( N492 ) , .CK( clk ) , .Q( text_out[37] ) );
  DFF_X1 text_out_reg_38 (.D( N491 ) , .CK( clk ) , .Q( text_out[38] ) );
  DFF_X1 text_out_reg_39 (.D( N490 ) , .CK( clk ) , .Q( text_out[39] ) );
  DFF_X1 text_out_reg_4 (.D( N501 ) , .CK( clk ) , .Q( text_out[4] ) );
  DFF_X1 text_out_reg_40 (.D( N465 ) , .CK( clk ) , .Q( text_out[40] ) );
  DFF_X1 text_out_reg_41 (.D( N464 ) , .CK( clk ) , .Q( text_out[41] ) );
  DFF_X1 text_out_reg_42 (.D( N463 ) , .CK( clk ) , .Q( text_out[42] ) );
  DFF_X1 text_out_reg_43 (.D( N462 ) , .CK( clk ) , .Q( text_out[43] ) );
  DFF_X1 text_out_reg_44 (.D( N461 ) , .CK( clk ) , .Q( text_out[44] ) );
  DFF_X1 text_out_reg_45 (.D( N460 ) , .CK( clk ) , .Q( text_out[45] ) );
  DFF_X1 text_out_reg_46 (.D( N459 ) , .CK( clk ) , .Q( text_out[46] ) );
  DFF_X1 text_out_reg_47 (.D( N458 ) , .CK( clk ) , .Q( text_out[47] ) );
  DFF_X1 text_out_reg_48 (.D( N433 ) , .CK( clk ) , .Q( text_out[48] ) );
  DFF_X1 text_out_reg_49 (.D( N432 ) , .CK( clk ) , .Q( text_out[49] ) );
  DFF_X1 text_out_reg_5 (.D( N500 ) , .CK( clk ) , .Q( text_out[5] ) );
  DFF_X1 text_out_reg_50 (.D( N431 ) , .CK( clk ) , .Q( text_out[50] ) );
  DFF_X1 text_out_reg_51 (.D( N430 ) , .CK( clk ) , .Q( text_out[51] ) );
  DFF_X1 text_out_reg_52 (.D( N429 ) , .CK( clk ) , .Q( text_out[52] ) );
  DFF_X1 text_out_reg_53 (.D( N428 ) , .CK( clk ) , .Q( text_out[53] ) );
  DFF_X1 text_out_reg_54 (.D( N427 ) , .CK( clk ) , .Q( text_out[54] ) );
  DFF_X1 text_out_reg_55 (.D( N426 ) , .CK( clk ) , .Q( text_out[55] ) );
  DFF_X1 text_out_reg_56 (.D( N401 ) , .CK( clk ) , .Q( text_out[56] ) );
  DFF_X1 text_out_reg_57 (.D( N400 ) , .CK( clk ) , .Q( text_out[57] ) );
  DFF_X1 text_out_reg_58 (.D( N399 ) , .CK( clk ) , .Q( text_out[58] ) );
  DFF_X1 text_out_reg_59 (.D( N398 ) , .CK( clk ) , .Q( text_out[59] ) );
  DFF_X1 text_out_reg_6 (.D( N499 ) , .CK( clk ) , .Q( text_out[6] ) );
  DFF_X1 text_out_reg_60 (.D( N397 ) , .CK( clk ) , .Q( text_out[60] ) );
  DFF_X1 text_out_reg_61 (.D( N396 ) , .CK( clk ) , .Q( text_out[61] ) );
  DFF_X1 text_out_reg_62 (.D( N395 ) , .CK( clk ) , .Q( text_out[62] ) );
  DFF_X1 text_out_reg_63 (.D( N394 ) , .CK( clk ) , .Q( text_out[63] ) );
  DFF_X1 text_out_reg_64 (.D( N489 ) , .CK( clk ) , .Q( text_out[64] ) );
  DFF_X1 text_out_reg_65 (.D( N488 ) , .CK( clk ) , .Q( text_out[65] ) );
  DFF_X1 text_out_reg_66 (.D( N487 ) , .CK( clk ) , .Q( text_out[66] ) );
  DFF_X1 text_out_reg_67 (.D( N486 ) , .CK( clk ) , .Q( text_out[67] ) );
  DFF_X1 text_out_reg_68 (.D( N485 ) , .CK( clk ) , .Q( text_out[68] ) );
  DFF_X1 text_out_reg_69 (.D( N484 ) , .CK( clk ) , .Q( text_out[69] ) );
  DFF_X1 text_out_reg_7 (.D( N498 ) , .CK( clk ) , .Q( text_out[7] ) );
  DFF_X1 text_out_reg_70 (.D( N483 ) , .CK( clk ) , .Q( text_out[70] ) );
  DFF_X1 text_out_reg_71 (.D( N482 ) , .CK( clk ) , .Q( text_out[71] ) );
  DFF_X1 text_out_reg_72 (.D( N457 ) , .CK( clk ) , .Q( text_out[72] ) );
  DFF_X1 text_out_reg_73 (.D( N456 ) , .CK( clk ) , .Q( text_out[73] ) );
  DFF_X1 text_out_reg_74 (.D( N455 ) , .CK( clk ) , .Q( text_out[74] ) );
  DFF_X1 text_out_reg_75 (.D( N454 ) , .CK( clk ) , .Q( text_out[75] ) );
  DFF_X1 text_out_reg_76 (.D( N453 ) , .CK( clk ) , .Q( text_out[76] ) );
  DFF_X1 text_out_reg_77 (.D( N452 ) , .CK( clk ) , .Q( text_out[77] ) );
  DFF_X1 text_out_reg_78 (.D( N451 ) , .CK( clk ) , .Q( text_out[78] ) );
  DFF_X1 text_out_reg_79 (.D( N450 ) , .CK( clk ) , .Q( text_out[79] ) );
  DFF_X1 text_out_reg_8 (.D( N473 ) , .CK( clk ) , .Q( text_out[8] ) );
  DFF_X1 text_out_reg_80 (.D( N425 ) , .CK( clk ) , .Q( text_out[80] ) );
  DFF_X1 text_out_reg_81 (.D( N424 ) , .CK( clk ) , .Q( text_out[81] ) );
  DFF_X1 text_out_reg_82 (.D( N423 ) , .CK( clk ) , .Q( text_out[82] ) );
  DFF_X1 text_out_reg_83 (.D( N422 ) , .CK( clk ) , .Q( text_out[83] ) );
  DFF_X1 text_out_reg_84 (.D( N421 ) , .CK( clk ) , .Q( text_out[84] ) );
  DFF_X1 text_out_reg_85 (.D( N420 ) , .CK( clk ) , .Q( text_out[85] ) );
  DFF_X1 text_out_reg_86 (.D( N419 ) , .CK( clk ) , .Q( text_out[86] ) );
  DFF_X1 text_out_reg_87 (.D( N418 ) , .CK( clk ) , .Q( text_out[87] ) );
  DFF_X1 text_out_reg_88 (.D( N393 ) , .CK( clk ) , .Q( text_out[88] ) );
  DFF_X1 text_out_reg_89 (.D( N392 ) , .CK( clk ) , .Q( text_out[89] ) );
  DFF_X1 text_out_reg_9 (.D( N472 ) , .CK( clk ) , .Q( text_out[9] ) );
  DFF_X1 text_out_reg_90 (.D( N391 ) , .CK( clk ) , .Q( text_out[90] ) );
  DFF_X1 text_out_reg_91 (.D( N390 ) , .CK( clk ) , .Q( text_out[91] ) );
  DFF_X1 text_out_reg_92 (.D( N389 ) , .CK( clk ) , .Q( text_out[92] ) );
  DFF_X1 text_out_reg_93 (.D( N388 ) , .CK( clk ) , .Q( text_out[93] ) );
  DFF_X1 text_out_reg_94 (.D( N387 ) , .CK( clk ) , .Q( text_out[94] ) );
  DFF_X1 text_out_reg_95 (.D( N386 ) , .CK( clk ) , .Q( text_out[95] ) );
  DFF_X1 text_out_reg_96 (.D( N481 ) , .CK( clk ) , .Q( text_out[96] ) );
  DFF_X1 text_out_reg_97 (.D( N480 ) , .CK( clk ) , .Q( text_out[97] ) );
  DFF_X1 text_out_reg_98 (.D( N479 ) , .CK( clk ) , .Q( text_out[98] ) );
  DFF_X1 text_out_reg_99 (.D( N478 ) , .CK( clk ) , .Q( text_out[99] ) );
  NAND2_X1 u0_U100 (.A1( key[62] ) , .A2( ld ) , .ZN( u0_n163 ) );
  NAND2_X1 u0_U101 (.A1( key[15] ) , .A2( ld ) , .ZN( u0_n114 ) );
  NAND2_X1 u0_U102 (.A1( key[74] ) , .A2( ld ) , .ZN( u0_n267 ) );
  NAND2_X1 u0_U103 (.A1( key[10] ) , .A2( ld ) , .ZN( u0_n129 ) );
  NAND2_X1 u0_U104 (.A1( key[72] ) , .A2( ld ) , .ZN( u0_n271 ) );
  NAND2_X1 u0_U105 (.A2( key[127] ) , .A1( ld ) , .ZN( u0_n2 ) );
  NAND2_X1 u0_U106 (.A1( key[6] ) , .A2( ld ) , .ZN( u0_n141 ) );
  NAND2_X1 u0_U107 (.A1( key[2] ) , .A2( ld ) , .ZN( u0_n153 ) );
  NAND2_X1 u0_U108 (.A1( key[73] ) , .A2( ld ) , .ZN( u0_n269 ) );
  NAND2_X1 u0_U109 (.A1( key[30] ) , .A2( ld ) , .ZN( u0_n69 ) );
  XNOR2_X1 u0_U11 (.ZN( u0_n41 ) , .B( u0_subword_11 ) , .A( w0_11 ) );
  NAND2_X1 u0_U110 (.A1( key[29] ) , .A2( ld ) , .ZN( u0_n72 ) );
  NAND2_X1 u0_U111 (.A1( key[17] ) , .A2( ld ) , .ZN( u0_n108 ) );
  NAND2_X1 u0_U112 (.A1( key[18] ) , .A2( ld ) , .ZN( u0_n105 ) );
  NAND2_X1 u0_U113 (.A1( key[16] ) , .A2( ld ) , .ZN( u0_n111 ) );
  NAND2_X1 u0_U114 (.A1( key[9] ) , .A2( ld ) , .ZN( u0_n132 ) );
  NAND2_X1 u0_U115 (.A1( key[19] ) , .A2( ld ) , .ZN( u0_n102 ) );
  NAND2_X1 u0_U116 (.A1( key[8] ) , .A2( ld ) , .ZN( u0_n135 ) );
  NAND2_X1 u0_U117 (.A1( key[3] ) , .A2( ld ) , .ZN( u0_n150 ) );
  NAND2_X1 u0_U118 (.A1( key[0] ) , .A2( ld ) , .ZN( u0_n159 ) );
  NAND2_X1 u0_U119 (.A1( key[5] ) , .A2( ld ) , .ZN( u0_n144 ) );
  XNOR2_X1 u0_U12 (.ZN( u0_n33 ) , .B( u0_subword_15 ) , .A( w0_15 ) );
  NAND2_X1 u0_U120 (.A1( key[1] ) , .A2( ld ) , .ZN( u0_n156 ) );
  OAI21_X1 u0_U121 (.B1( ld ) , .ZN( u0_N181 ) , .B2( u0_n139 ) , .A( u0_n209 ) );
  NAND2_X1 u0_U122 (.A1( key[39] ) , .A2( ld ) , .ZN( u0_n209 ) );
  OAI21_X1 u0_U123 (.B1( ld ) , .ZN( u0_N135 ) , .B2( u0_n170 ) , .A( u0_n233 ) );
  NAND2_X1 u0_U124 (.A1( key[91] ) , .A2( ld ) , .ZN( u0_n233 ) );
  OAI21_X1 u0_U125 (.B1( ld ) , .ZN( u0_N57 ) , .B2( u0_n33 ) , .A( u0_n34 ) );
  NAND2_X1 u0_U126 (.A1( key[111] ) , .A2( ld ) , .ZN( u0_n34 ) );
  OAI21_X1 u0_U127 (.B1( ld ) , .ZN( u0_N46 ) , .B2( u0_n55 ) , .A( u0_n56 ) );
  NAND2_X1 u0_U128 (.A1( key[100] ) , .A2( ld ) , .ZN( u0_n56 ) );
  OAI21_X1 u0_U129 (.B1( ld ) , .ZN( u0_N45 ) , .B2( u0_n57 ) , .A( u0_n58 ) );
  XNOR2_X1 u0_U13 (.ZN( u0_n17 ) , .B( u0_subword_23 ) , .A( w0_23 ) );
  NAND2_X1 u0_U130 (.A1( key[99] ) , .A2( ld ) , .ZN( u0_n58 ) );
  OAI21_X1 u0_U131 (.B1( ld ) , .ZN( u0_N43 ) , .B2( u0_n61 ) , .A( u0_n62 ) );
  NAND2_X1 u0_U132 (.A1( key[97] ) , .A2( ld ) , .ZN( u0_n62 ) );
  OAI21_X1 u0_U133 (.B1( ld ) , .ZN( u0_N54 ) , .B2( u0_n39 ) , .A( u0_n40 ) );
  NAND2_X1 u0_U134 (.A1( key[108] ) , .A2( ld ) , .ZN( u0_n40 ) );
  OAI21_X1 u0_U135 (.B1( ld ) , .ZN( u0_N51 ) , .B2( u0_n45 ) , .A( u0_n46 ) );
  NAND2_X1 u0_U136 (.A1( key[105] ) , .A2( ld ) , .ZN( u0_n46 ) );
  OAI21_X1 u0_U137 (.B1( ld ) , .ZN( u0_N65 ) , .B2( u0_n17 ) , .A( u0_n18 ) );
  NAND2_X1 u0_U138 (.A1( key[119] ) , .A2( ld ) , .ZN( u0_n18 ) );
  OAI21_X1 u0_U139 (.B1( ld ) , .ZN( u0_N71 ) , .B2( u0_n5 ) , .A( u0_n6 ) );
  XNOR2_X1 u0_U14 (.ZN( u0_n45 ) , .B( u0_subword_9 ) , .A( w0_9 ) );
  NAND2_X1 u0_U140 (.A1( key[125] ) , .A2( ld ) , .ZN( u0_n6 ) );
  OAI21_X1 u0_U141 (.B1( ld ) , .ZN( u0_N70 ) , .B2( u0_n7 ) , .A( u0_n8 ) );
  NAND2_X1 u0_U142 (.A1( key[124] ) , .A2( ld ) , .ZN( u0_n8 ) );
  OAI21_X1 u0_U143 (.B1( ld ) , .ZN( u0_N69 ) , .A( u0_n10 ) , .B2( u0_n9 ) );
  NAND2_X1 u0_U144 (.A1( key[123] ) , .A2( ld ) , .ZN( u0_n10 ) );
  OAI21_X1 u0_U145 (.B1( ld ) , .ZN( u0_N123 ) , .B2( u0_n194 ) , .A( u0_n257 ) );
  NAND2_X1 u0_U146 (.A1( key[79] ) , .A2( ld ) , .ZN( u0_n257 ) );
  OAI21_X1 u0_U147 (.B1( ld ) , .ZN( u0_N131 ) , .B2( u0_n178 ) , .A( u0_n241 ) );
  NAND2_X1 u0_U148 (.A1( key[87] ) , .A2( ld ) , .ZN( u0_n241 ) );
  OAI21_X1 u0_U149 (.B1( ld ) , .ZN( u0_N121 ) , .B2( u0_n198 ) , .A( u0_n261 ) );
  XNOR2_X1 u0_U15 (.ZN( u0_n23 ) , .B( u0_subword_20 ) , .A( w0_20 ) );
  NAND2_X1 u0_U150 (.A1( key[77] ) , .A2( ld ) , .ZN( u0_n261 ) );
  OAI21_X1 u0_U151 (.B1( ld ) , .ZN( u0_N47 ) , .B2( u0_n53 ) , .A( u0_n54 ) );
  NAND2_X1 u0_U152 (.A1( key[101] ) , .A2( ld ) , .ZN( u0_n54 ) );
  OAI21_X1 u0_U153 (.B1( ld ) , .ZN( u0_N63 ) , .B2( u0_n21 ) , .A( u0_n22 ) );
  NAND2_X1 u0_U154 (.A1( key[117] ) , .A2( ld ) , .ZN( u0_n22 ) );
  OAI21_X1 u0_U155 (.B1( ld ) , .ZN( u0_N129 ) , .B2( u0_n182 ) , .A( u0_n245 ) );
  NAND2_X1 u0_U156 (.A1( key[85] ) , .A2( ld ) , .ZN( u0_n245 ) );
  OAI21_X1 u0_U157 (.B1( ld ) , .ZN( u0_N62 ) , .B2( u0_n23 ) , .A( u0_n24 ) );
  NAND2_X1 u0_U158 (.A1( key[116] ) , .A2( ld ) , .ZN( u0_n24 ) );
  OAI21_X1 u0_U159 (.B1( ld ) , .ZN( u0_N55 ) , .B2( u0_n37 ) , .A( u0_n38 ) );
  XNOR2_X1 u0_U16 (.ZN( u0_n37 ) , .B( u0_subword_13 ) , .A( w0_13 ) );
  NAND2_X1 u0_U160 (.A1( key[109] ) , .A2( ld ) , .ZN( u0_n38 ) );
  OAI21_X1 u0_U161 (.B1( ld ) , .ZN( u0_N120 ) , .B2( u0_n200 ) , .A( u0_n263 ) );
  NAND2_X1 u0_U162 (.A1( key[76] ) , .A2( ld ) , .ZN( u0_n263 ) );
  OAI21_X1 u0_U163 (.B1( ld ) , .ZN( u0_N53 ) , .B2( u0_n41 ) , .A( u0_n42 ) );
  NAND2_X1 u0_U164 (.A1( key[107] ) , .A2( ld ) , .ZN( u0_n42 ) );
  OAI21_X1 u0_U165 (.B1( ld ) , .ZN( u0_N268 ) , .B2( u0_n74 ) , .A( u0_n75 ) );
  NAND2_X1 u0_U166 (.A1( key[28] ) , .A2( ld ) , .ZN( u0_n75 ) );
  OAI21_X1 u0_U167 (.B1( ld ) , .ZN( u0_N271 ) , .B2( u0_n65 ) , .A( u0_n66 ) );
  NAND2_X1 u0_U168 (.A1( key[31] ) , .A2( ld ) , .ZN( u0_n66 ) );
  OAI21_X1 u0_U169 (.B1( ld ) , .ZN( u0_N260 ) , .B2( u0_n98 ) , .A( u0_n99 ) );
  NAND2_X1 u0_U170 (.A1( key[20] ) , .A2( ld ) , .ZN( u0_n99 ) );
  OAI21_X1 u0_U171 (.B1( ld ) , .ZN( u0_N251 ) , .B2( u0_n125 ) , .A( u0_n126 ) );
  NAND2_X1 u0_U172 (.A1( key[11] ) , .A2( ld ) , .ZN( u0_n126 ) );
  OAI21_X1 u0_U173 (.B1( ld ) , .ZN( u0_N244 ) , .B2( u0_n146 ) , .A( u0_n147 ) );
  NAND2_X1 u0_U174 (.A1( key[4] ) , .A2( ld ) , .ZN( u0_n147 ) );
  OAI21_X1 u0_U175 (.B1( ld ) , .ZN( u0_N115 ) , .B2( u0_n210 ) , .A( u0_n273 ) );
  NAND2_X1 u0_U176 (.A1( key[71] ) , .A2( ld ) , .ZN( u0_n273 ) );
  OAI21_X1 u0_U177 (.B1( ld ) , .ZN( u0_N113 ) , .B2( u0_n214 ) , .A( u0_n277 ) );
  NAND2_X1 u0_U178 (.A1( key[69] ) , .A2( ld ) , .ZN( u0_n277 ) );
  OAI21_X1 u0_U179 (.B1( ld ) , .ZN( u0_N111 ) , .B2( u0_n218 ) , .A( u0_n281 ) );
  XNOR2_X1 u0_U18 (.ZN( u0_n21 ) , .B( u0_subword_21 ) , .A( w0_21 ) );
  NAND2_X1 u0_U180 (.A1( key[67] ) , .A2( ld ) , .ZN( u0_n281 ) );
  XNOR2_X1 u0_U181 (.ZN( u0_n226 ) , .B( u0_subword_31 ) , .A( w0_31 ) );
  OAI21_X1 u0_U182 (.B1( ld ) , .ZN( u0_N42 ) , .B2( u0_n63 ) , .A( u0_n64 ) );
  OAI21_X1 u0_U184 (.B1( ld ) , .ZN( u0_N50 ) , .B2( u0_n47 ) , .A( u0_n48 ) );
  OAI21_X1 u0_U186 (.B1( ld ) , .ZN( u0_N44 ) , .B2( u0_n59 ) , .A( u0_n60 ) );
  OAI21_X1 u0_U187 (.B1( ld ) , .ZN( u0_N59 ) , .B2( u0_n29 ) , .A( u0_n30 ) );
  OAI21_X1 u0_U188 (.B1( ld ) , .ZN( u0_N247 ) , .B2( u0_n137 ) , .A( u0_n138 ) );
  OAI21_X1 u0_U189 (.B1( ld ) , .ZN( u0_N67 ) , .B2( u0_n13 ) , .A( u0_n14 ) );
  NAND2_X1 u0_U19 (.A1( key[22] ) , .A2( ld ) , .ZN( u0_n93 ) );
  OAI21_X1 u0_U190 (.B1( ld ) , .ZN( u0_N252 ) , .B2( u0_n122 ) , .A( u0_n123 ) );
  OAI21_X1 u0_U191 (.B1( ld ) , .ZN( u0_N186 ) , .B2( u0_n124 ) , .A( u0_n199 ) );
  OAI21_X1 u0_U192 (.B1( ld ) , .ZN( u0_N269 ) , .B2( u0_n71 ) , .A( u0_n72 ) );
  OAI21_X1 u0_U193 (.B1( ld ) , .ZN( u0_N73 ) , .B2( u0_n1 ) , .A( u0_n2 ) );
  XNOR2_X1 u0_U194 (.ZN( u0_n15 ) , .A( u0_n240 ) , .B( u0_n246 ) );
  XNOR2_X1 u0_U195 (.B( u0_n248 ) , .ZN( u0_n86 ) , .A( u0_n88 ) );
  OAI21_X1 u0_U196 (.B1( ld ) , .ZN( u0_N254 ) , .B2( u0_n116 ) , .A( u0_n117 ) );
  OAI21_X1 u0_U197 (.B1( ld ) , .ZN( u0_N109 ) , .B2( u0_n222 ) , .A( u0_n285 ) );
  OAI21_X1 u0_U198 (.B1( ld ) , .ZN( u0_N119 ) , .B2( u0_n202 ) , .A( u0_n265 ) );
  OAI21_X1 u0_U199 (.B1( ld ) , .ZN( u0_N185 ) , .B2( u0_n127 ) , .A( u0_n201 ) );
  XNOR2_X1 u0_U20 (.ZN( u0_n25 ) , .B( u0_subword_19 ) , .A( w0_19 ) );
  OAI21_X1 u0_U200 (.B1( ld ) , .ZN( u0_N136 ) , .B2( u0_n168 ) , .A( u0_n231 ) );
  OAI21_X1 u0_U201 (.B1( ld ) , .ZN( u0_N202 ) , .A( u0_n167 ) , .B2( u0_n76 ) );
  XNOR2_X1 u0_U202 (.ZN( u0_n31 ) , .B( u0_subword_16 ) , .A( w0_16 ) );
  INV_X1 u0_U203 (.A( u0_n250 ) , .ZN( w3_13 ) );
  OAI21_X1 u0_U204 (.B1( ld ) , .ZN( u0_N128 ) , .B2( u0_n184 ) , .A( u0_n247 ) );
  OAI21_X1 u0_U205 (.B1( ld ) , .ZN( u0_N194 ) , .B2( u0_n100 ) , .A( u0_n183 ) );
  INV_X1 u0_U206 (.A( u0_n254 ) , .ZN( w3_14 ) );
  OAI21_X1 u0_U207 (.B1( ld ) , .ZN( u0_N245 ) , .B2( u0_n143 ) , .A( u0_n144 ) );
  OAI21_X1 u0_U208 (.B1( ld ) , .ZN( u0_N179 ) , .B2( u0_n145 ) , .A( u0_n213 ) );
  OAI21_X1 u0_U209 (.B1( ld ) , .ZN( u0_N249 ) , .B2( u0_n131 ) , .A( u0_n132 ) );
  INV_X1 u0_U210 (.A( u0_n258 ) , .ZN( w3_12 ) );
  XNOR2_X1 u0_U211 (.ZN( u0_n43 ) , .B( u0_subword_10 ) , .A( w0_10 ) );
  OAI21_X1 u0_U213 (.B1( ld ) , .ZN( u0_N49 ) , .B2( u0_n49 ) , .A( u0_n50 ) );
  OAI21_X1 u0_U214 (.B1( ld ) , .ZN( u0_N125 ) , .B2( u0_n190 ) , .A( u0_n253 ) );
  XNOR2_X1 u0_U215 (.ZN( u0_n164 ) , .B( u0_n262 ) , .A( u0_n3 ) );
  OAI21_X1 u0_U216 (.B1( ld ) , .ZN( u0_N262 ) , .B2( u0_n92 ) , .A( u0_n93 ) );
  XNOR2_X1 u0_U217 (.ZN( u0_n27 ) , .B( u0_subword_18 ) , .A( w0_18 ) );
  OAI21_X1 u0_U218 (.B1( ld ) , .ZN( u0_N139 ) , .B2( u0_n162 ) , .A( u0_n225 ) );
  OAI21_X1 u0_U219 (.B1( ld ) , .ZN( u0_N205 ) , .A( u0_n161 ) , .B2( u0_n67 ) );
  XNOR2_X1 u0_U22 (.ZN( u0_n29 ) , .B( u0_subword_17 ) , .A( w0_17 ) );
  OAI21_X1 u0_U220 (.B1( ld ) , .ZN( u0_N112 ) , .B2( u0_n216 ) , .A( u0_n279 ) );
  OAI21_X1 u0_U221 (.B1( ld ) , .ZN( u0_N178 ) , .B2( u0_n148 ) , .A( u0_n215 ) );
  OAI21_X1 u0_U222 (.B1( ld ) , .ZN( u0_N246 ) , .B2( u0_n140 ) , .A( u0_n141 ) );
  OAI21_X1 u0_U223 (.B1( ld ) , .ZN( u0_N243 ) , .B2( u0_n149 ) , .A( u0_n150 ) );
  OAI21_X1 u0_U224 (.B1( ld ) , .ZN( u0_N177 ) , .B2( u0_n151 ) , .A( u0_n217 ) );
  OAI21_X1 u0_U225 (.B1( ld ) , .ZN( u0_N133 ) , .B2( u0_n174 ) , .A( u0_n237 ) );
  OAI21_X1 u0_U226 (.B1( ld ) , .ZN( u0_N259 ) , .B2( u0_n101 ) , .A( u0_n102 ) );
  OAI21_X1 u0_U227 (.B1( ld ) , .ZN( u0_N61 ) , .B2( u0_n25 ) , .A( u0_n26 ) );
  OAI21_X1 u0_U228 (.B1( ld ) , .ZN( u0_N255 ) , .B2( u0_n113 ) , .A( u0_n114 ) );
  OAI21_X1 u0_U229 (.B1( ld ) , .ZN( u0_N189 ) , .B2( u0_n115 ) , .A( u0_n193 ) );
  XNOR2_X1 u0_U23 (.ZN( u0_n39 ) , .B( u0_subword_12 ) , .A( w0_12 ) );
  INV_X1 u0_U230 (.A( u0_n264 ) , .ZN( w3_15 ) );
  OAI21_X1 u0_U231 (.B1( ld ) , .ZN( u0_N263 ) , .B2( u0_n89 ) , .A( u0_n90 ) );
  OAI21_X1 u0_U232 (.B1( ld ) , .ZN( u0_N197 ) , .A( u0_n177 ) , .B2( u0_n91 ) );
  OAI21_X1 u0_U233 (.B1( ld ) , .ZN( u0_N117 ) , .B2( u0_n206 ) , .A( u0_n269 ) );
  OAI21_X1 u0_U234 (.B1( ld ) , .ZN( u0_N183 ) , .B2( u0_n133 ) , .A( u0_n205 ) );
  XNOR2_X1 u0_U235 (.ZN( u0_n47 ) , .B( u0_subword_8 ) , .A( w0_8 ) );
  OAI21_X1 u0_U236 (.B1( ld ) , .ZN( u0_N127 ) , .B2( u0_n186 ) , .A( u0_n249 ) );
  OAI21_X1 u0_U237 (.B1( ld ) , .ZN( u0_N193 ) , .B2( u0_n103 ) , .A( u0_n185 ) );
  OAI21_X1 u0_U238 (.B1( ld ) , .ZN( u0_N241 ) , .B2( u0_n155 ) , .A( u0_n156 ) );
  OAI21_X1 u0_U239 (.B1( ld ) , .ZN( u0_N175 ) , .B2( u0_n157 ) , .A( u0_n221 ) );
  NAND2_X1 u0_U24 (.A1( key[47] ) , .A2( ld ) , .ZN( u0_n193 ) );
  XNOR2_X1 u0_U240 (.ZN( u0_n35 ) , .B( u0_subword_14 ) , .A( w0_14 ) );
  OAI21_X1 u0_U241 (.B1( ld ) , .ZN( u0_N257 ) , .B2( u0_n107 ) , .A( u0_n108 ) );
  OAI21_X1 u0_U242 (.B1( ld ) , .ZN( u0_N191 ) , .B2( u0_n109 ) , .A( u0_n189 ) );
  OAI21_X1 u0_U243 (.B1( ld ) , .ZN( u0_N48 ) , .B2( u0_n51 ) , .A( u0_n52 ) );
  OAI21_X1 u0_U244 (.B1( ld ) , .ZN( u0_N116 ) , .B2( u0_n208 ) , .A( u0_n271 ) );
  OAI21_X1 u0_U245 (.B1( ld ) , .ZN( u0_N264 ) , .B2( u0_n86 ) , .A( u0_n87 ) );
  OAI21_X1 u0_U246 (.B1( ld ) , .ZN( u0_N66 ) , .B2( u0_n15 ) , .A( u0_n16 ) );
  OAI21_X1 u0_U247 (.B1( ld ) , .ZN( u0_N64 ) , .B2( u0_n19 ) , .A( u0_n20 ) );
  OAI21_X1 u0_U249 (.B1( ld ) , .ZN( u0_N265 ) , .B2( u0_n83 ) , .A( u0_n84 ) );
  NAND2_X1 u0_U25 (.A1( key[55] ) , .A2( ld ) , .ZN( u0_n177 ) );
  OAI21_X1 u0_U250 (.B1( ld ) , .ZN( u0_N199 ) , .A( u0_n173 ) , .B2( u0_n85 ) );
  OAI21_X1 u0_U251 (.B1( ld ) , .ZN( u0_N108 ) , .B2( u0_n224 ) , .A( u0_n287 ) );
  OAI21_X1 u0_U252 (.B1( ld ) , .ZN( u0_N256 ) , .B2( u0_n110 ) , .A( u0_n111 ) );
  OAI21_X1 u0_U253 (.B1( ld ) , .ZN( u0_N58 ) , .B2( u0_n31 ) , .A( u0_n32 ) );
  XNOR2_X1 u0_U254 (.ZN( u0_n240 ) , .B( u0_subword_24 ) , .A( w0_24 ) );
  OAI21_X1 u0_U255 (.B1( ld ) , .ZN( u0_N267 ) , .B2( u0_n77 ) , .A( u0_n78 ) );
  OAI21_X1 u0_U256 (.B1( ld ) , .ZN( u0_N201 ) , .A( u0_n169 ) , .B2( u0_n79 ) );
  OAI21_X1 u0_U257 (.B1( ld ) , .ZN( u0_N72 ) , .B2( u0_n3 ) , .A( u0_n4 ) );
  OAI21_X1 u0_U258 (.B1( ld ) , .ZN( u0_N138 ) , .B2( u0_n164 ) , .A( u0_n227 ) );
  XNOR2_X1 u0_U259 (.ZN( u0_n51 ) , .B( u0_subword_6 ) , .A( w0_6 ) );
  NAND2_X1 u0_U26 (.A1( key[37] ) , .A2( ld ) , .ZN( u0_n213 ) );
  XNOR2_X1 u0_U260 (.ZN( u0_n230 ) , .B( u0_subword_29 ) , .A( w0_29 ) );
  OAI21_X1 u0_U261 (.B1( ld ) , .ZN( u0_N56 ) , .B2( u0_n35 ) , .A( u0_n36 ) );
  XNOR2_X1 u0_U262 (.ZN( u0_n19 ) , .B( u0_subword_22 ) , .A( w0_22 ) );
  OAI21_X1 u0_U263 (.B1( ld ) , .ZN( u0_N261 ) , .B2( u0_n95 ) , .A( u0_n96 ) );
  OAI21_X1 u0_U264 (.B1( ld ) , .ZN( u0_N195 ) , .A( u0_n181 ) , .B2( u0_n97 ) );
  OAI21_X1 u0_U265 (.B1( ld ) , .ZN( u0_N137 ) , .B2( u0_n166 ) , .A( u0_n229 ) );
  OAI21_X1 u0_U266 (.B1( ld ) , .ZN( u0_N203 ) , .A( u0_n165 ) , .B2( u0_n73 ) );
  OAI21_X1 u0_U267 (.B1( ld ) , .ZN( u0_N266 ) , .B2( u0_n80 ) , .A( u0_n81 ) );
  OAI21_X1 u0_U268 (.B1( ld ) , .ZN( u0_N114 ) , .B2( u0_n212 ) , .A( u0_n275 ) );
  OAI21_X1 u0_U269 (.B1( ld ) , .ZN( u0_N180 ) , .B2( u0_n142 ) , .A( u0_n211 ) );
  NAND2_X1 u0_U27 (.A1( key[35] ) , .A2( ld ) , .ZN( u0_n217 ) );
  OAI21_X1 u0_U270 (.B1( ld ) , .ZN( u0_N130 ) , .B2( u0_n180 ) , .A( u0_n243 ) );
  OAI21_X1 u0_U271 (.B1( ld ) , .ZN( u0_N196 ) , .A( u0_n179 ) , .B2( u0_n94 ) );
  OAI21_X1 u0_U272 (.B1( ld ) , .ZN( u0_N242 ) , .B2( u0_n152 ) , .A( u0_n153 ) );
  OAI21_X1 u0_U273 (.B1( ld ) , .ZN( u0_N122 ) , .B2( u0_n196 ) , .A( u0_n259 ) );
  OAI21_X1 u0_U274 (.B1( ld ) , .ZN( u0_N188 ) , .B2( u0_n118 ) , .A( u0_n195 ) );
  OAI21_X1 u0_U275 (.B1( ld ) , .ZN( u0_N253 ) , .B2( u0_n119 ) , .A( u0_n120 ) );
  OAI21_X1 u0_U276 (.B1( ld ) , .ZN( u0_N187 ) , .B2( u0_n121 ) , .A( u0_n197 ) );
  OAI21_X1 u0_U277 (.B1( ld ) , .ZN( u0_N270 ) , .B2( u0_n68 ) , .A( u0_n69 ) );
  OAI21_X1 u0_U278 (.B1( ld ) , .ZN( u0_N204 ) , .A( u0_n163 ) , .B2( u0_n70 ) );
  OAI21_X1 u0_U279 (.B1( ld ) , .ZN( u0_N124 ) , .B2( u0_n192 ) , .A( u0_n255 ) );
  NAND2_X1 u0_U28 (.A1( key[93] ) , .A2( ld ) , .ZN( u0_n229 ) );
  OAI21_X1 u0_U280 (.B1( ld ) , .ZN( u0_N190 ) , .B2( u0_n112 ) , .A( u0_n191 ) );
  OAI21_X1 u0_U281 (.B1( ld ) , .ZN( u0_N248 ) , .B2( u0_n134 ) , .A( u0_n135 ) );
  OAI21_X1 u0_U282 (.B1( ld ) , .ZN( u0_N182 ) , .B2( u0_n136 ) , .A( u0_n207 ) );
  OAI21_X1 u0_U283 (.B1( ld ) , .ZN( u0_N132 ) , .B2( u0_n176 ) , .A( u0_n239 ) );
  OAI21_X1 u0_U284 (.B1( ld ) , .ZN( u0_N198 ) , .A( u0_n175 ) , .B2( u0_n88 ) );
  OAI21_X1 u0_U285 (.B1( ld ) , .ZN( u0_N240 ) , .B2( u0_n158 ) , .A( u0_n159 ) );
  OAI21_X1 u0_U286 (.B1( ld ) , .ZN( u0_N174 ) , .B2( u0_n160 ) , .A( u0_n223 ) );
  XNOR2_X1 u0_U287 (.ZN( u0_n236 ) , .A( u0_subword_26 ) , .B( w0_26 ) );
  OAI21_X1 u0_U288 (.B1( ld ) , .ZN( u0_N52 ) , .B2( u0_n43 ) , .A( u0_n44 ) );
  OAI21_X1 u0_U289 (.B1( ld ) , .ZN( u0_N118 ) , .B2( u0_n204 ) , .A( u0_n267 ) );
  NAND2_X1 u0_U29 (.A1( key[92] ) , .A2( ld ) , .ZN( u0_n231 ) );
  OAI21_X1 u0_U290 (.B1( ld ) , .ZN( u0_N60 ) , .B2( u0_n27 ) , .A( u0_n28 ) );
  XOR2_X1 u0_U291 (.Z( u0_n65 ) , .A( u0_n67 ) , .B( w3_31 ) );
  XOR2_X1 u0_U292 (.Z( u0_n68 ) , .A( u0_n70 ) , .B( w3_30 ) );
  XOR2_X1 u0_U293 (.Z( u0_n71 ) , .A( u0_n73 ) , .B( w3_29 ) );
  XOR2_X1 u0_U294 (.Z( u0_n74 ) , .A( u0_n76 ) , .B( w3_28 ) );
  XOR2_X1 u0_U295 (.Z( u0_n77 ) , .A( u0_n79 ) , .B( w3_27 ) );
  XOR2_X1 u0_U296 (.Z( u0_n80 ) , .A( u0_n82 ) , .B( w3_26 ) );
  XOR2_X1 u0_U297 (.Z( u0_n83 ) , .A( u0_n85 ) , .B( w3_25 ) );
  OAI21_X1 u0_U298 (.B1( ld ) , .ZN( u0_N126 ) , .B2( u0_n188 ) , .A( u0_n251 ) );
  XOR2_X1 u0_U299 (.Z( u0_n89 ) , .A( u0_n91 ) , .B( w3_23 ) );
  XNOR2_X1 u0_U3 (.A( u0_n11 ) , .ZN( u0_n172 ) , .B( u0_n242 ) );
  NAND2_X1 u0_U30 (.A1( key[59] ) , .A2( ld ) , .ZN( u0_n169 ) );
  XOR2_X1 u0_U300 (.Z( u0_n92 ) , .A( u0_n94 ) , .B( w3_22 ) );
  XOR2_X1 u0_U301 (.Z( u0_n95 ) , .A( u0_n97 ) , .B( w3_21 ) );
  XOR2_X1 u0_U302 (.A( u0_n100 ) , .Z( u0_n98 ) , .B( w3_20 ) );
  XOR2_X1 u0_U303 (.Z( u0_n101 ) , .A( u0_n103 ) , .B( w3_19 ) );
  XOR2_X1 u0_U304 (.Z( u0_n104 ) , .A( u0_n106 ) , .B( w3_18 ) );
  XOR2_X1 u0_U305 (.Z( u0_n107 ) , .A( u0_n109 ) , .B( w3_17 ) );
  XOR2_X1 u0_U306 (.Z( u0_n110 ) , .A( u0_n112 ) , .B( w3_16 ) );
  XOR2_X1 u0_U307 (.Z( u0_n113 ) , .A( u0_n115 ) , .B( w3_15 ) );
  XOR2_X1 u0_U308 (.Z( u0_n116 ) , .A( u0_n118 ) , .B( w3_14 ) );
  XOR2_X1 u0_U309 (.Z( u0_n119 ) , .A( u0_n121 ) , .B( w3_13 ) );
  NAND2_X1 u0_U31 (.A1( key[53] ) , .A2( ld ) , .ZN( u0_n181 ) );
  XOR2_X1 u0_U310 (.Z( u0_n122 ) , .A( u0_n124 ) , .B( w3_12 ) );
  XOR2_X1 u0_U311 (.Z( u0_n125 ) , .A( u0_n127 ) , .B( w3_11 ) );
  XOR2_X1 u0_U312 (.Z( u0_n128 ) , .A( u0_n130 ) , .B( w3_10 ) );
  XOR2_X1 u0_U313 (.Z( u0_n131 ) , .A( u0_n133 ) , .B( w3_9 ) );
  XOR2_X1 u0_U314 (.Z( u0_n134 ) , .A( u0_n136 ) , .B( w3_8 ) );
  XOR2_X1 u0_U315 (.Z( u0_n137 ) , .A( u0_n139 ) , .B( w3_7 ) );
  XOR2_X1 u0_U316 (.Z( u0_n140 ) , .A( u0_n142 ) , .B( w3_6 ) );
  XOR2_X1 u0_U317 (.Z( u0_n143 ) , .A( u0_n145 ) , .B( w3_5 ) );
  XOR2_X1 u0_U318 (.Z( u0_n146 ) , .A( u0_n148 ) , .B( w3_4 ) );
  XOR2_X1 u0_U319 (.Z( u0_n149 ) , .A( u0_n151 ) , .B( w3_3 ) );
  NAND2_X1 u0_U32 (.A1( key[45] ) , .A2( ld ) , .ZN( u0_n197 ) );
  XOR2_X1 u0_U320 (.Z( u0_n152 ) , .A( u0_n154 ) , .B( w3_2 ) );
  XOR2_X1 u0_U321 (.Z( u0_n155 ) , .A( u0_n157 ) , .B( w3_1 ) );
  XOR2_X1 u0_U322 (.Z( u0_n158 ) , .A( u0_n160 ) , .B( w3_0 ) );
  XOR2_X1 u0_U323 (.A( u0_n162 ) , .Z( u0_n67 ) , .B( w2_31 ) );
  XOR2_X1 u0_U324 (.A( u0_n164 ) , .Z( u0_n70 ) , .B( w2_30 ) );
  XOR2_X1 u0_U325 (.A( u0_n166 ) , .Z( u0_n73 ) , .B( w2_29 ) );
  XOR2_X1 u0_U326 (.A( u0_n168 ) , .Z( u0_n76 ) , .B( w2_28 ) );
  XOR2_X1 u0_U327 (.A( u0_n170 ) , .Z( u0_n79 ) , .B( w2_27 ) );
  OAI21_X1 u0_U328 (.B1( ld ) , .ZN( u0_N68 ) , .B2( u0_n11 ) , .A( u0_n12 ) );
  XOR2_X1 u0_U329 (.A( u0_n174 ) , .Z( u0_n85 ) , .B( w2_25 ) );
  NAND2_X1 u0_U33 (.A1( key[44] ) , .A2( ld ) , .ZN( u0_n199 ) );
  XOR2_X1 u0_U330 (.A( u0_n176 ) , .Z( u0_n88 ) , .B( w2_24 ) );
  XOR2_X1 u0_U331 (.A( u0_n178 ) , .Z( u0_n91 ) , .B( w2_23 ) );
  XOR2_X1 u0_U332 (.A( u0_n180 ) , .Z( u0_n94 ) , .B( w2_22 ) );
  XOR2_X1 u0_U333 (.A( u0_n182 ) , .Z( u0_n97 ) , .B( w2_21 ) );
  XOR2_X1 u0_U334 (.Z( u0_n100 ) , .A( u0_n184 ) , .B( w2_20 ) );
  XOR2_X1 u0_U335 (.Z( u0_n103 ) , .A( u0_n186 ) , .B( w2_19 ) );
  XOR2_X1 u0_U336 (.Z( u0_n106 ) , .A( u0_n188 ) , .B( w2_18 ) );
  XOR2_X1 u0_U337 (.Z( u0_n109 ) , .A( u0_n190 ) , .B( w2_17 ) );
  XOR2_X1 u0_U338 (.Z( u0_n112 ) , .A( u0_n192 ) , .B( w2_16 ) );
  XOR2_X1 u0_U339 (.Z( u0_n115 ) , .A( u0_n194 ) , .B( w2_15 ) );
  NAND2_X1 u0_U34 (.A1( key[65] ) , .A2( ld ) , .ZN( u0_n285 ) );
  XOR2_X1 u0_U340 (.Z( u0_n118 ) , .A( u0_n196 ) , .B( w2_14 ) );
  XOR2_X1 u0_U341 (.Z( u0_n121 ) , .A( u0_n198 ) , .B( w2_13 ) );
  XOR2_X1 u0_U342 (.Z( u0_n124 ) , .A( u0_n200 ) , .B( w2_12 ) );
  XOR2_X1 u0_U343 (.Z( u0_n127 ) , .A( u0_n202 ) , .B( w2_11 ) );
  XOR2_X1 u0_U344 (.Z( u0_n130 ) , .A( u0_n204 ) , .B( w2_10 ) );
  XOR2_X1 u0_U345 (.Z( u0_n133 ) , .A( u0_n206 ) , .B( w2_9 ) );
  XOR2_X1 u0_U346 (.Z( u0_n136 ) , .A( u0_n208 ) , .B( w2_8 ) );
  XOR2_X1 u0_U347 (.Z( u0_n139 ) , .A( u0_n210 ) , .B( w2_7 ) );
  XOR2_X1 u0_U348 (.Z( u0_n142 ) , .A( u0_n212 ) , .B( w2_6 ) );
  XOR2_X1 u0_U349 (.Z( u0_n145 ) , .A( u0_n214 ) , .B( w2_5 ) );
  NAND2_X1 u0_U35 (.A1( key[68] ) , .A2( ld ) , .ZN( u0_n279 ) );
  XOR2_X1 u0_U350 (.Z( u0_n148 ) , .A( u0_n216 ) , .B( w2_4 ) );
  XOR2_X1 u0_U351 (.Z( u0_n151 ) , .A( u0_n218 ) , .B( w2_3 ) );
  XOR2_X1 u0_U352 (.Z( u0_n154 ) , .A( u0_n220 ) , .B( w2_2 ) );
  XOR2_X1 u0_U353 (.Z( u0_n157 ) , .A( u0_n222 ) , .B( w2_1 ) );
  XOR2_X1 u0_U354 (.Z( u0_n160 ) , .A( u0_n224 ) , .B( w2_0 ) );
  XOR2_X1 u0_U355 (.A( u0_n1 ) , .Z( u0_n162 ) , .B( w1_31 ) );
  XOR2_X1 u0_U356 (.Z( u0_n1 ) , .A( u0_n226 ) , .B( u0_rcon_31 ) );
  OAI21_X1 u0_U357 (.B1( ld ) , .ZN( u0_N258 ) , .B2( u0_n104 ) , .A( u0_n105 ) );
  XOR2_X1 u0_U358 (.A( u0_n228 ) , .Z( u0_n3 ) , .B( u0_rcon_30 ) );
  XOR2_X1 u0_U359 (.Z( u0_n166 ) , .A( u0_n5 ) , .B( w1_29 ) );
  NAND2_X1 u0_U36 (.A1( key[103] ) , .A2( ld ) , .ZN( u0_n50 ) );
  XOR2_X1 u0_U360 (.A( u0_n230 ) , .Z( u0_n5 ) , .B( u0_rcon_29 ) );
  XOR2_X1 u0_U361 (.Z( u0_n168 ) , .A( u0_n7 ) , .B( w1_28 ) );
  XOR2_X1 u0_U362 (.A( u0_n232 ) , .Z( u0_n7 ) , .B( u0_rcon_28 ) );
  XOR2_X1 u0_U363 (.Z( u0_n170 ) , .A( u0_n9 ) , .B( w1_27 ) );
  XOR2_X1 u0_U364 (.A( u0_n234 ) , .Z( u0_n9 ) , .B( u0_rcon_27 ) );
  OAI21_X1 u0_U365 (.B1( ld ) , .ZN( u0_N192 ) , .B2( u0_n106 ) , .A( u0_n187 ) );
  XOR2_X1 u0_U366 (.Z( u0_n11 ) , .A( u0_n236 ) , .B( u0_rcon_26 ) );
  XOR2_X1 u0_U367 (.A( u0_n13 ) , .Z( u0_n174 ) , .B( w1_25 ) );
  XOR2_X1 u0_U368 (.Z( u0_n13 ) , .A( u0_n238 ) , .B( u0_rcon_25 ) );
  XOR2_X1 u0_U369 (.A( u0_n15 ) , .Z( u0_n176 ) , .B( w1_24 ) );
  NAND2_X1 u0_U37 (.A1( key[102] ) , .A2( ld ) , .ZN( u0_n52 ) );
  OAI21_X1 u0_U370 (.B1( ld ) , .ZN( u0_N110 ) , .B2( u0_n220 ) , .A( u0_n283 ) );
  XOR2_X1 u0_U371 (.A( u0_n17 ) , .Z( u0_n178 ) , .B( w1_23 ) );
  OAI21_X1 u0_U372 (.B1( ld ) , .ZN( u0_N176 ) , .B2( u0_n154 ) , .A( u0_n219 ) );
  XOR2_X1 u0_U373 (.Z( u0_n180 ) , .A( u0_n19 ) , .B( w1_22 ) );
  OAI21_X1 u0_U374 (.B1( ld ) , .ZN( u0_N250 ) , .B2( u0_n128 ) , .A( u0_n129 ) );
  XOR2_X1 u0_U375 (.Z( u0_n182 ) , .A( u0_n21 ) , .B( w1_21 ) );
  OAI21_X1 u0_U376 (.B1( ld ) , .ZN( u0_N184 ) , .B2( u0_n130 ) , .A( u0_n203 ) );
  XOR2_X1 u0_U377 (.Z( u0_n184 ) , .A( u0_n23 ) , .B( w1_20 ) );
  OAI21_X1 u0_U378 (.B1( ld ) , .ZN( u0_N134 ) , .B2( u0_n172 ) , .A( u0_n235 ) );
  XOR2_X1 u0_U379 (.Z( u0_n186 ) , .A( u0_n25 ) , .B( w1_19 ) );
  NAND2_X1 u0_U38 (.A1( key[96] ) , .A2( ld ) , .ZN( u0_n64 ) );
  OAI21_X1 u0_U380 (.B1( ld ) , .ZN( u0_N200 ) , .A( u0_n171 ) , .B2( u0_n82 ) );
  XOR2_X1 u0_U381 (.Z( u0_n188 ) , .A( u0_n27 ) , .B( w1_18 ) );
  XOR2_X1 u0_U383 (.Z( u0_n190 ) , .A( u0_n29 ) , .B( w1_17 ) );
  XOR2_X1 u0_U385 (.Z( u0_n192 ) , .A( u0_n31 ) , .B( w1_16 ) );
  XOR2_X1 u0_U387 (.Z( u0_n194 ) , .A( u0_n33 ) , .B( w1_15 ) );
  XOR2_X1 u0_U389 (.Z( u0_n196 ) , .A( u0_n35 ) , .B( w1_14 ) );
  NAND2_X1 u0_U39 (.A1( key[115] ) , .A2( ld ) , .ZN( u0_n26 ) );
  XOR2_X1 u0_U391 (.Z( u0_n198 ) , .A( u0_n37 ) , .B( w1_13 ) );
  XOR2_X1 u0_U393 (.Z( u0_n200 ) , .A( u0_n39 ) , .B( w1_12 ) );
  XOR2_X1 u0_U395 (.Z( u0_n202 ) , .A( u0_n41 ) , .B( w1_11 ) );
  XOR2_X1 u0_U397 (.Z( u0_n204 ) , .A( u0_n43 ) , .B( w1_10 ) );
  XOR2_X1 u0_U399 (.Z( u0_n206 ) , .A( u0_n45 ) , .B( w1_9 ) );
  XNOR2_X1 u0_U4 (.A( u0_n172 ) , .B( u0_n244 ) , .ZN( u0_n82 ) );
  NAND2_X1 u0_U40 (.A1( key[114] ) , .A2( ld ) , .ZN( u0_n28 ) );
  XOR2_X1 u0_U401 (.Z( u0_n208 ) , .A( u0_n47 ) , .B( w1_8 ) );
  XOR2_X1 u0_U403 (.Z( u0_n210 ) , .A( u0_n49 ) , .B( w1_7 ) );
  XOR2_X1 u0_U405 (.Z( u0_n212 ) , .A( u0_n51 ) , .B( w1_6 ) );
  XOR2_X1 u0_U407 (.Z( u0_n214 ) , .A( u0_n53 ) , .B( w1_5 ) );
  XOR2_X1 u0_U409 (.Z( u0_n216 ) , .A( u0_n55 ) , .B( w1_4 ) );
  NAND2_X1 u0_U41 (.A1( key[112] ) , .A2( ld ) , .ZN( u0_n32 ) );
  XOR2_X1 u0_U411 (.Z( u0_n218 ) , .A( u0_n57 ) , .B( w1_3 ) );
  XOR2_X1 u0_U413 (.Z( u0_n220 ) , .A( u0_n59 ) , .B( w1_2 ) );
  XOR2_X1 u0_U415 (.Z( u0_n222 ) , .A( u0_n61 ) , .B( w1_1 ) );
  XOR2_X1 u0_U417 (.Z( u0_n224 ) , .A( u0_n63 ) , .B( w1_0 ) );
  NAND2_X1 u0_U42 (.A1( key[106] ) , .A2( ld ) , .ZN( u0_n44 ) );
  NAND2_X1 u0_U43 (.A1( key[64] ) , .A2( ld ) , .ZN( u0_n287 ) );
  NAND2_X1 u0_U44 (.A1( key[126] ) , .A2( ld ) , .ZN( u0_n4 ) );
  NAND2_X1 u0_U45 (.A1( key[23] ) , .A2( ld ) , .ZN( u0_n90 ) );
  NAND2_X1 u0_U46 (.A1( key[21] ) , .A2( ld ) , .ZN( u0_n96 ) );
  NAND2_X1 u0_U47 (.A1( key[24] ) , .A2( ld ) , .ZN( u0_n87 ) );
  NAND2_X1 u0_U48 (.A1( key[25] ) , .A2( ld ) , .ZN( u0_n84 ) );
  NAND2_X1 u0_U49 (.A1( key[122] ) , .A2( ld ) , .ZN( u0_n12 ) );
  XNOR2_X1 u0_U5 (.ZN( u0_n232 ) , .B( u0_subword_28 ) , .A( w0_28 ) );
  NAND2_X1 u0_U50 (.A1( key[118] ) , .A2( ld ) , .ZN( u0_n20 ) );
  NAND2_X1 u0_U51 (.A1( key[89] ) , .A2( ld ) , .ZN( u0_n237 ) );
  NAND2_X1 u0_U52 (.A1( key[120] ) , .A2( ld ) , .ZN( u0_n16 ) );
  NAND2_X1 u0_U53 (.A1( key[88] ) , .A2( ld ) , .ZN( u0_n239 ) );
  NAND2_X1 u0_U54 (.A1( key[86] ) , .A2( ld ) , .ZN( u0_n243 ) );
  NAND2_X1 u0_U55 (.A1( key[82] ) , .A2( ld ) , .ZN( u0_n251 ) );
  NAND2_X1 u0_U56 (.A1( key[80] ) , .A2( ld ) , .ZN( u0_n255 ) );
  NAND2_X1 u0_U57 (.A1( key[78] ) , .A2( ld ) , .ZN( u0_n259 ) );
  NAND2_X1 u0_U58 (.A1( key[26] ) , .A2( ld ) , .ZN( u0_n81 ) );
  NAND2_X1 u0_U59 (.A1( key[27] ) , .A2( ld ) , .ZN( u0_n78 ) );
  XNOR2_X1 u0_U6 (.ZN( u0_n234 ) , .B( u0_subword_27 ) , .A( w0_27 ) );
  NAND2_X1 u0_U60 (.A1( key[98] ) , .A2( ld ) , .ZN( u0_n60 ) );
  NAND2_X1 u0_U61 (.A1( key[121] ) , .A2( ld ) , .ZN( u0_n14 ) );
  NAND2_X1 u0_U62 (.A1( key[84] ) , .A2( ld ) , .ZN( u0_n247 ) );
  NAND2_X1 u0_U63 (.A1( key[83] ) , .A2( ld ) , .ZN( u0_n249 ) );
  NAND2_X1 u0_U64 (.A1( key[113] ) , .A2( ld ) , .ZN( u0_n30 ) );
  NAND2_X1 u0_U65 (.A1( key[81] ) , .A2( ld ) , .ZN( u0_n253 ) );
  NAND2_X1 u0_U66 (.A1( key[110] ) , .A2( ld ) , .ZN( u0_n36 ) );
  NAND2_X1 u0_U67 (.A1( key[75] ) , .A2( ld ) , .ZN( u0_n265 ) );
  NAND2_X1 u0_U68 (.A1( key[104] ) , .A2( ld ) , .ZN( u0_n48 ) );
  NAND2_X1 u0_U69 (.A1( key[95] ) , .A2( ld ) , .ZN( u0_n225 ) );
  XNOR2_X1 u0_U7 (.ZN( u0_n228 ) , .B( u0_subword_30 ) , .A( w0_30 ) );
  NAND2_X1 u0_U70 (.A1( key[63] ) , .A2( ld ) , .ZN( u0_n161 ) );
  NAND2_X1 u0_U71 (.A1( key[38] ) , .A2( ld ) , .ZN( u0_n211 ) );
  NAND2_X1 u0_U72 (.A1( key[36] ) , .A2( ld ) , .ZN( u0_n215 ) );
  NAND2_X1 u0_U73 (.A1( key[34] ) , .A2( ld ) , .ZN( u0_n219 ) );
  NAND2_X1 u0_U74 (.A1( key[33] ) , .A2( ld ) , .ZN( u0_n221 ) );
  NAND2_X1 u0_U75 (.A1( key[32] ) , .A2( ld ) , .ZN( u0_n223 ) );
  NAND2_X1 u0_U76 (.A1( key[94] ) , .A2( ld ) , .ZN( u0_n227 ) );
  NAND2_X1 u0_U77 (.A1( key[61] ) , .A2( ld ) , .ZN( u0_n165 ) );
  NAND2_X1 u0_U78 (.A1( key[60] ) , .A2( ld ) , .ZN( u0_n167 ) );
  NAND2_X1 u0_U79 (.A1( key[90] ) , .A2( ld ) , .ZN( u0_n235 ) );
  XNOR2_X1 u0_U8 (.ZN( u0_n238 ) , .B( u0_subword_25 ) , .A( w0_25 ) );
  NAND2_X1 u0_U80 (.A1( key[58] ) , .A2( ld ) , .ZN( u0_n171 ) );
  NAND2_X1 u0_U81 (.A1( key[57] ) , .A2( ld ) , .ZN( u0_n173 ) );
  NAND2_X1 u0_U82 (.A1( key[56] ) , .A2( ld ) , .ZN( u0_n175 ) );
  NAND2_X1 u0_U83 (.A1( key[54] ) , .A2( ld ) , .ZN( u0_n179 ) );
  NAND2_X1 u0_U84 (.A1( key[52] ) , .A2( ld ) , .ZN( u0_n183 ) );
  NAND2_X1 u0_U85 (.A1( key[51] ) , .A2( ld ) , .ZN( u0_n185 ) );
  NAND2_X1 u0_U86 (.A1( key[50] ) , .A2( ld ) , .ZN( u0_n187 ) );
  NAND2_X1 u0_U87 (.A1( key[49] ) , .A2( ld ) , .ZN( u0_n189 ) );
  NAND2_X1 u0_U88 (.A1( key[48] ) , .A2( ld ) , .ZN( u0_n191 ) );
  NAND2_X1 u0_U89 (.A1( key[46] ) , .A2( ld ) , .ZN( u0_n195 ) );
  INV_X1 u0_U9 (.ZN( u0_n246 ) , .A( u0_rcon_24 ) );
  NAND2_X1 u0_U90 (.A1( key[43] ) , .A2( ld ) , .ZN( u0_n201 ) );
  NAND2_X1 u0_U91 (.A1( key[42] ) , .A2( ld ) , .ZN( u0_n203 ) );
  NAND2_X1 u0_U92 (.A1( key[41] ) , .A2( ld ) , .ZN( u0_n205 ) );
  NAND2_X1 u0_U93 (.A1( key[40] ) , .A2( ld ) , .ZN( u0_n207 ) );
  NAND2_X1 u0_U94 (.A1( key[13] ) , .A2( ld ) , .ZN( u0_n120 ) );
  NAND2_X1 u0_U95 (.A1( key[14] ) , .A2( ld ) , .ZN( u0_n117 ) );
  NAND2_X1 u0_U96 (.A1( key[12] ) , .A2( ld ) , .ZN( u0_n123 ) );
  NAND2_X1 u0_U97 (.A1( key[7] ) , .A2( ld ) , .ZN( u0_n138 ) );
  NAND2_X1 u0_U98 (.A1( key[70] ) , .A2( ld ) , .ZN( u0_n275 ) );
  NAND2_X1 u0_U99 (.A1( key[66] ) , .A2( ld ) , .ZN( u0_n283 ) );
  OAI21_X1 u0_r0_U27 (.ZN( u0_r0_N70 ) , .B1( u0_r0_n4 ) , .B2( u0_r0_n5 ) , .A( u0_r0_n9 ) );
  NAND4_X1 u0_r0_U28 (.A3( u0_r0_N78 ) , .A2( u0_r0_n12 ) , .ZN( u0_r0_n14 ) , .A1( u0_r0_n18 ) , .A4( u0_r0_n2 ) );
  NAND2_X1 u0_r0_U29 (.A1( u0_r0_N80 ) , .ZN( u0_r0_n11 ) , .A2( u0_r0_n17 ) );
  NOR2_X1 u0_r0_U30 (.A2( ld ) , .ZN( u0_r0_N79 ) , .A1( u0_r0_n12 ) );
  NOR2_X1 u0_r0_U31 (.A2( ld ) , .ZN( u0_r0_N80 ) , .A1( u0_r0_n18 ) );
  NAND2_X1 u0_r0_U32 (.ZN( u0_r0_N71 ) , .A1( u0_r0_n10 ) , .A2( u0_r0_n23 ) );
  INV_X1 u0_r0_U33 (.A( u0_r0_n17 ) , .ZN( u0_r0_n2 ) );
  INV_X1 u0_r0_U34 (.A( u0_r0_n24 ) , .ZN( u0_r0_n5 ) );
  INV_X1 u0_r0_U35 (.A( u0_r0_n25 ) , .ZN( u0_r0_n4 ) );
  XNOR2_X1 u0_r0_U36 (.ZN( u0_r0_n12 ) , .B( u0_r0_rcnt_0 ) , .A( u0_r0_rcnt_1 ) );
  OAI21_X1 u0_r0_U37 (.B1( u0_r0_n12 ) , .A( u0_r0_n21 ) , .ZN( u0_r0_n25 ) , .B2( u0_r0_n6 ) );
  NAND4_X1 u0_r0_U38 (.ZN( u0_r0_n10 ) , .A1( u0_r0_n24 ) , .A2( u0_r0_n25 ) , .A4( u0_r0_n3 ) , .A3( u0_r0_n9 ) );
  OAI22_X1 u0_r0_U39 (.ZN( u0_r0_N73 ) , .B1( u0_r0_n16 ) , .A2( u0_r0_n19 ) , .B2( u0_r0_n20 ) , .A1( u0_r0_rcnt_0 ) );
  NAND2_X1 u0_r0_U40 (.A1( u0_r0_n12 ) , .ZN( u0_r0_n20 ) , .A2( u0_r0_rcnt_0 ) );
  NOR3_X1 u0_r0_U41 (.ZN( u0_r0_N76 ) , .A1( u0_r0_n11 ) , .A2( u0_r0_n12 ) , .A3( u0_r0_n8 ) );
  NOR3_X1 u0_r0_U42 (.ZN( u0_r0_N77 ) , .A1( u0_r0_n11 ) , .A3( u0_r0_n12 ) , .A2( u0_r0_rcnt_0 ) );
  NAND2_X1 u0_r0_U43 (.ZN( u0_r0_n21 ) , .A1( u0_r0_rcnt_0 ) , .A2( u0_r0_rcnt_1 ) );
  NOR2_X1 u0_r0_U44 (.A2( ld ) , .ZN( u0_r0_N78 ) , .A1( u0_r0_rcnt_0 ) );
  OAI21_X1 u0_r0_U45 (.ZN( u0_r0_N72 ) , .A( u0_r0_n14 ) , .B2( u0_r0_n19 ) , .B1( u0_r0_n8 ) );
  OAI21_X1 u0_r0_U46 (.ZN( u0_r0_N75 ) , .B1( u0_r0_n11 ) , .B2( u0_r0_n13 ) , .A( u0_r0_n14 ) );
  NAND2_X1 u0_r0_U47 (.A1( u0_r0_n12 ) , .ZN( u0_r0_n13 ) , .A2( u0_r0_n8 ) );
  NOR2_X1 u0_r0_U48 (.A2( u0_r0_n21 ) , .ZN( u0_r0_n22 ) , .A1( u0_r0_n6 ) );
  OAI21_X1 u0_r0_U49 (.B1( u0_r0_N70 ) , .ZN( u0_r0_N81 ) , .A( u0_r0_n10 ) , .B2( u0_r0_n3 ) );
  NAND2_X1 u0_r0_U50 (.ZN( u0_r0_N74 ) , .A2( u0_r0_n1 ) , .A1( u0_r0_n14 ) );
  INV_X1 u0_r0_U51 (.ZN( u0_r0_n1 ) , .A( u0_r0_n15 ) );
  AOI211_X1 u0_r0_U52 (.C2( u0_r0_n11 ) , .ZN( u0_r0_n15 ) , .C1( u0_r0_n16 ) , .B( u0_r0_n7 ) , .A( u0_r0_n8 ) );
  INV_X1 u0_r0_U53 (.A( u0_r0_n12 ) , .ZN( u0_r0_n7 ) );
  INV_X1 u0_r0_U54 (.A( ld ) , .ZN( u0_r0_n9 ) );
  NAND3_X1 u0_r0_U55 (.ZN( u0_r0_n16 ) , .A3( u0_r0_n18 ) , .A1( u0_r0_n2 ) , .A2( u0_r0_n9 ) );
  NAND3_X1 u0_r0_U56 (.A3( u0_r0_N79 ) , .A1( u0_r0_n17 ) , .A2( u0_r0_n18 ) , .ZN( u0_r0_n19 ) );
  XOR2_X1 u0_r0_U57 (.Z( u0_r0_n18 ) , .A( u0_r0_n21 ) , .B( u0_r0_rcnt_2 ) );
  XOR2_X1 u0_r0_U58 (.Z( u0_r0_n17 ) , .B( u0_r0_n22 ) , .A( u0_r0_n3 ) );
  NAND3_X1 u0_r0_U59 (.ZN( u0_r0_n23 ) , .A3( u0_r0_n4 ) , .A1( u0_r0_n5 ) , .A2( u0_r0_n9 ) );
  XOR2_X1 u0_r0_U60 (.B( u0_r0_n12 ) , .Z( u0_r0_n24 ) , .A( u0_r0_n6 ) );
  DFF_X1 u0_r0_out_reg_24 (.CK( clk ) , .D( u0_r0_N70 ) , .Q( u0_rcon_24 ) );
  DFF_X1 u0_r0_out_reg_25 (.CK( clk ) , .D( u0_r0_N71 ) , .Q( u0_rcon_25 ) );
  DFF_X1 u0_r0_out_reg_26 (.CK( clk ) , .D( u0_r0_N72 ) , .Q( u0_rcon_26 ) );
  DFF_X1 u0_r0_out_reg_27 (.CK( clk ) , .D( u0_r0_N73 ) , .Q( u0_rcon_27 ) );
  DFF_X1 u0_r0_out_reg_28 (.CK( clk ) , .D( u0_r0_N74 ) , .Q( u0_rcon_28 ) );
  DFF_X1 u0_r0_out_reg_29 (.CK( clk ) , .D( u0_r0_N75 ) , .Q( u0_rcon_29 ) );
  DFF_X1 u0_r0_out_reg_30 (.CK( clk ) , .D( u0_r0_N76 ) , .Q( u0_rcon_30 ) );
  DFF_X1 u0_r0_out_reg_31 (.CK( clk ) , .D( u0_r0_N77 ) , .Q( u0_rcon_31 ) );
  DFF_X1 u0_r0_rcnt_reg_0 (.CK( clk ) , .D( u0_r0_N78 ) , .QN( u0_r0_n8 ) , .Q( u0_r0_rcnt_0 ) );
  DFF_X1 u0_r0_rcnt_reg_1 (.CK( clk ) , .D( u0_r0_N79 ) , .Q( u0_r0_rcnt_1 ) );
  DFF_X1 u0_r0_rcnt_reg_2 (.CK( clk ) , .D( u0_r0_N80 ) , .QN( u0_r0_n6 ) , .Q( u0_r0_rcnt_2 ) );
  DFF_X1 u0_r0_rcnt_reg_3 (.CK( clk ) , .D( u0_r0_N81 ) , .QN( u0_r0_n3 ) );
  DFF_X1 u0_w_reg_0_0 (.CK( clk ) , .D( u0_N42 ) , .Q( w0_0 ) );
  DFF_X1 u0_w_reg_0_1 (.CK( clk ) , .D( u0_N43 ) , .Q( w0_1 ) );
  DFF_X1 u0_w_reg_0_10 (.CK( clk ) , .D( u0_N52 ) , .Q( w0_10 ) );
  DFF_X1 u0_w_reg_0_11 (.CK( clk ) , .D( u0_N53 ) , .Q( w0_11 ) );
  DFF_X1 u0_w_reg_0_12 (.CK( clk ) , .D( u0_N54 ) , .Q( w0_12 ) );
  DFF_X1 u0_w_reg_0_13 (.CK( clk ) , .D( u0_N55 ) , .Q( w0_13 ) );
  DFF_X1 u0_w_reg_0_14 (.CK( clk ) , .D( u0_N56 ) , .Q( w0_14 ) );
  DFF_X1 u0_w_reg_0_15 (.CK( clk ) , .D( u0_N57 ) , .Q( w0_15 ) );
  DFF_X1 u0_w_reg_0_16 (.CK( clk ) , .D( u0_N58 ) , .Q( w0_16 ) );
  DFF_X1 u0_w_reg_0_17 (.CK( clk ) , .D( u0_N59 ) , .Q( w0_17 ) );
  DFF_X1 u0_w_reg_0_18 (.CK( clk ) , .D( u0_N60 ) , .Q( w0_18 ) );
  DFF_X1 u0_w_reg_0_19 (.CK( clk ) , .D( u0_N61 ) , .Q( w0_19 ) );
  DFF_X1 u0_w_reg_0_2 (.CK( clk ) , .D( u0_N44 ) , .Q( w0_2 ) );
  DFF_X1 u0_w_reg_0_20 (.CK( clk ) , .D( u0_N62 ) , .Q( w0_20 ) );
  DFF_X1 u0_w_reg_0_21 (.CK( clk ) , .D( u0_N63 ) , .Q( w0_21 ) );
  DFF_X1 u0_w_reg_0_22 (.CK( clk ) , .D( u0_N64 ) , .Q( w0_22 ) );
  DFF_X1 u0_w_reg_0_23 (.CK( clk ) , .D( u0_N65 ) , .Q( w0_23 ) );
  DFF_X1 u0_w_reg_0_24 (.CK( clk ) , .D( u0_N66 ) , .Q( w0_24 ) );
  DFF_X1 u0_w_reg_0_25 (.CK( clk ) , .D( u0_N67 ) , .Q( w0_25 ) );
  DFF_X1 u0_w_reg_0_26 (.CK( clk ) , .D( u0_N68 ) , .Q( w0_26 ) );
  DFF_X1 u0_w_reg_0_27 (.CK( clk ) , .D( u0_N69 ) , .Q( w0_27 ) );
  DFF_X1 u0_w_reg_0_28 (.CK( clk ) , .D( u0_N70 ) , .Q( w0_28 ) );
  DFF_X1 u0_w_reg_0_29 (.CK( clk ) , .D( u0_N71 ) , .Q( w0_29 ) );
  DFF_X1 u0_w_reg_0_3 (.CK( clk ) , .D( u0_N45 ) , .Q( w0_3 ) );
  DFF_X1 u0_w_reg_0_30 (.CK( clk ) , .D( u0_N72 ) , .Q( w0_30 ) );
  DFF_X1 u0_w_reg_0_31 (.CK( clk ) , .D( u0_N73 ) , .Q( w0_31 ) );
  DFF_X1 u0_w_reg_0_4 (.CK( clk ) , .D( u0_N46 ) , .Q( w0_4 ) );
  DFF_X1 u0_w_reg_0_5 (.CK( clk ) , .D( u0_N47 ) , .Q( w0_5 ) );
  DFF_X1 u0_w_reg_0_6 (.CK( clk ) , .D( u0_N48 ) , .Q( w0_6 ) );
  DFF_X1 u0_w_reg_0_7 (.CK( clk ) , .D( u0_N49 ) , .Q( w0_7 ) );
  DFF_X1 u0_w_reg_0_8 (.CK( clk ) , .D( u0_N50 ) , .Q( w0_8 ) );
  DFF_X1 u0_w_reg_0_9 (.CK( clk ) , .D( u0_N51 ) , .Q( w0_9 ) );
  DFF_X1 u0_w_reg_1_0 (.CK( clk ) , .D( u0_N108 ) , .Q( w1_0 ) );
  DFF_X1 u0_w_reg_1_1 (.CK( clk ) , .D( u0_N109 ) , .Q( w1_1 ) );
  DFF_X1 u0_w_reg_1_10 (.CK( clk ) , .D( u0_N118 ) , .Q( w1_10 ) );
  DFF_X1 u0_w_reg_1_11 (.CK( clk ) , .D( u0_N119 ) , .Q( w1_11 ) );
  DFF_X1 u0_w_reg_1_12 (.CK( clk ) , .D( u0_N120 ) , .Q( w1_12 ) );
  DFF_X1 u0_w_reg_1_13 (.CK( clk ) , .D( u0_N121 ) , .Q( w1_13 ) );
  DFF_X1 u0_w_reg_1_14 (.CK( clk ) , .D( u0_N122 ) , .Q( w1_14 ) );
  DFF_X1 u0_w_reg_1_15 (.CK( clk ) , .D( u0_N123 ) , .Q( w1_15 ) );
  DFF_X1 u0_w_reg_1_16 (.CK( clk ) , .D( u0_N124 ) , .Q( w1_16 ) );
  DFF_X1 u0_w_reg_1_17 (.CK( clk ) , .D( u0_N125 ) , .Q( w1_17 ) );
  DFF_X1 u0_w_reg_1_18 (.CK( clk ) , .D( u0_N126 ) , .Q( w1_18 ) );
  DFF_X1 u0_w_reg_1_19 (.CK( clk ) , .D( u0_N127 ) , .Q( w1_19 ) );
  DFF_X1 u0_w_reg_1_2 (.CK( clk ) , .D( u0_N110 ) , .Q( w1_2 ) );
  DFF_X1 u0_w_reg_1_20 (.CK( clk ) , .D( u0_N128 ) , .Q( w1_20 ) );
  DFF_X1 u0_w_reg_1_21 (.CK( clk ) , .D( u0_N129 ) , .Q( w1_21 ) );
  DFF_X1 u0_w_reg_1_22 (.CK( clk ) , .D( u0_N130 ) , .Q( w1_22 ) );
  DFF_X1 u0_w_reg_1_23 (.CK( clk ) , .D( u0_N131 ) , .Q( w1_23 ) );
  DFF_X1 u0_w_reg_1_24 (.CK( clk ) , .D( u0_N132 ) , .Q( w1_24 ) );
  DFF_X1 u0_w_reg_1_25 (.CK( clk ) , .D( u0_N133 ) , .Q( w1_25 ) );
  DFF_X1 u0_w_reg_1_26 (.CK( clk ) , .D( u0_N134 ) , .QN( u0_n242 ) , .Q( w1_26 ) );
  DFF_X1 u0_w_reg_1_27 (.CK( clk ) , .D( u0_N135 ) , .Q( w1_27 ) );
  DFF_X1 u0_w_reg_1_28 (.CK( clk ) , .D( u0_N136 ) , .Q( w1_28 ) );
  DFF_X1 u0_w_reg_1_29 (.CK( clk ) , .D( u0_N137 ) , .Q( w1_29 ) );
  DFF_X1 u0_w_reg_1_3 (.CK( clk ) , .D( u0_N111 ) , .Q( w1_3 ) );
  DFF_X1 u0_w_reg_1_30 (.CK( clk ) , .D( u0_N138 ) , .QN( u0_n262 ) , .Q( w1_30 ) );
  DFF_X1 u0_w_reg_1_31 (.CK( clk ) , .D( u0_N139 ) , .Q( w1_31 ) );
  DFF_X1 u0_w_reg_1_4 (.CK( clk ) , .D( u0_N112 ) , .Q( w1_4 ) );
  DFF_X1 u0_w_reg_1_5 (.CK( clk ) , .D( u0_N113 ) , .Q( w1_5 ) );
  DFF_X1 u0_w_reg_1_6 (.CK( clk ) , .D( u0_N114 ) , .Q( w1_6 ) );
  DFF_X1 u0_w_reg_1_7 (.CK( clk ) , .D( u0_N115 ) , .Q( w1_7 ) );
  DFF_X1 u0_w_reg_1_8 (.CK( clk ) , .D( u0_N116 ) , .Q( w1_8 ) );
  DFF_X1 u0_w_reg_1_9 (.CK( clk ) , .D( u0_N117 ) , .Q( w1_9 ) );
  DFF_X1 u0_w_reg_2_0 (.CK( clk ) , .D( u0_N174 ) , .Q( w2_0 ) );
  DFF_X1 u0_w_reg_2_1 (.CK( clk ) , .D( u0_N175 ) , .Q( w2_1 ) );
  DFF_X1 u0_w_reg_2_10 (.CK( clk ) , .D( u0_N184 ) , .Q( w2_10 ) );
  DFF_X1 u0_w_reg_2_11 (.CK( clk ) , .D( u0_N185 ) , .Q( w2_11 ) );
  DFF_X1 u0_w_reg_2_12 (.CK( clk ) , .D( u0_N186 ) , .Q( w2_12 ) );
  DFF_X1 u0_w_reg_2_13 (.CK( clk ) , .D( u0_N187 ) , .Q( w2_13 ) );
  DFF_X1 u0_w_reg_2_14 (.CK( clk ) , .D( u0_N188 ) , .Q( w2_14 ) );
  DFF_X1 u0_w_reg_2_15 (.CK( clk ) , .D( u0_N189 ) , .Q( w2_15 ) );
  DFF_X1 u0_w_reg_2_16 (.CK( clk ) , .D( u0_N190 ) , .Q( w2_16 ) );
  DFF_X1 u0_w_reg_2_17 (.CK( clk ) , .D( u0_N191 ) , .Q( w2_17 ) );
  DFF_X1 u0_w_reg_2_18 (.CK( clk ) , .D( u0_N192 ) , .Q( w2_18 ) );
  DFF_X1 u0_w_reg_2_19 (.CK( clk ) , .D( u0_N193 ) , .Q( w2_19 ) );
  DFF_X1 u0_w_reg_2_2 (.CK( clk ) , .D( u0_N176 ) , .Q( w2_2 ) );
  DFF_X1 u0_w_reg_2_20 (.CK( clk ) , .D( u0_N194 ) , .Q( w2_20 ) );
  DFF_X1 u0_w_reg_2_21 (.CK( clk ) , .D( u0_N195 ) , .Q( w2_21 ) );
  DFF_X1 u0_w_reg_2_22 (.CK( clk ) , .D( u0_N196 ) , .Q( w2_22 ) );
  DFF_X1 u0_w_reg_2_23 (.CK( clk ) , .D( u0_N197 ) , .Q( w2_23 ) );
  DFF_X1 u0_w_reg_2_24 (.CK( clk ) , .D( u0_N198 ) , .Q( w2_24 ) );
  DFF_X1 u0_w_reg_2_25 (.CK( clk ) , .D( u0_N199 ) , .Q( w2_25 ) );
  DFF_X1 u0_w_reg_2_26 (.CK( clk ) , .D( u0_N200 ) , .QN( u0_n244 ) , .Q( w2_26 ) );
  DFF_X1 u0_w_reg_2_27 (.CK( clk ) , .D( u0_N201 ) , .Q( w2_27 ) );
  DFF_X1 u0_w_reg_2_28 (.CK( clk ) , .D( u0_N202 ) , .Q( w2_28 ) );
  DFF_X1 u0_w_reg_2_29 (.CK( clk ) , .D( u0_N203 ) , .Q( w2_29 ) );
  DFF_X1 u0_w_reg_2_3 (.CK( clk ) , .D( u0_N177 ) , .Q( w2_3 ) );
  DFF_X1 u0_w_reg_2_30 (.CK( clk ) , .D( u0_N204 ) , .Q( w2_30 ) );
  DFF_X1 u0_w_reg_2_31 (.CK( clk ) , .D( u0_N205 ) , .Q( w2_31 ) );
  DFF_X1 u0_w_reg_2_4 (.CK( clk ) , .D( u0_N178 ) , .Q( w2_4 ) );
  DFF_X1 u0_w_reg_2_5 (.CK( clk ) , .D( u0_N179 ) , .Q( w2_5 ) );
  DFF_X1 u0_w_reg_2_6 (.CK( clk ) , .D( u0_N180 ) , .Q( w2_6 ) );
  DFF_X1 u0_w_reg_2_7 (.CK( clk ) , .D( u0_N181 ) , .Q( w2_7 ) );
  DFF_X1 u0_w_reg_2_8 (.CK( clk ) , .D( u0_N182 ) , .Q( w2_8 ) );
  DFF_X1 u0_w_reg_2_9 (.CK( clk ) , .D( u0_N183 ) , .Q( w2_9 ) );
  DFF_X1 u0_w_reg_3_0 (.CK( clk ) , .D( u0_N240 ) , .Q( w3_0 ) );
  DFF_X1 u0_w_reg_3_1 (.CK( clk ) , .D( u0_N241 ) , .Q( w3_1 ) );
  DFF_X1 u0_w_reg_3_10 (.CK( clk ) , .D( u0_N250 ) , .Q( w3_10 ) );
  DFF_X1 u0_w_reg_3_11 (.CK( clk ) , .D( u0_N251 ) , .Q( w3_11 ) );
  DFF_X1 u0_w_reg_3_12 (.CK( clk ) , .D( u0_N252 ) , .QN( u0_n258 ) , .Q( u0_n274 ) );
  DFF_X1 u0_w_reg_3_13 (.CK( clk ) , .D( u0_N253 ) , .QN( u0_n250 ) , .Q( u0_n272 ) );
  DFF_X1 u0_w_reg_3_14 (.CK( clk ) , .D( u0_N254 ) , .QN( u0_n254 ) , .Q( u0_n270 ) );
  DFF_X1 u0_w_reg_3_15 (.CK( clk ) , .D( u0_N255 ) , .QN( u0_n264 ) , .Q( u0_n268 ) );
  DFF_X1 u0_w_reg_3_16 (.CK( clk ) , .D( u0_N256 ) , .Q( w3_16 ) );
  DFF_X1 u0_w_reg_3_17 (.CK( clk ) , .D( u0_N257 ) , .Q( w3_17 ) );
  DFF_X1 u0_w_reg_3_18 (.CK( clk ) , .D( u0_N258 ) , .Q( w3_18 ) );
  DFF_X1 u0_w_reg_3_19 (.CK( clk ) , .D( u0_N259 ) , .Q( w3_19 ) );
  DFF_X1 u0_w_reg_3_2 (.CK( clk ) , .D( u0_N242 ) , .Q( w3_2 ) );
  DFF_X1 u0_w_reg_3_20 (.CK( clk ) , .D( u0_N260 ) , .Q( w3_20 ) );
  DFF_X1 u0_w_reg_3_21 (.CK( clk ) , .D( u0_N261 ) , .Q( w3_21 ) );
  DFF_X1 u0_w_reg_3_22 (.CK( clk ) , .D( u0_N262 ) , .Q( w3_22 ) );
  DFF_X1 u0_w_reg_3_23 (.CK( clk ) , .D( u0_N263 ) , .Q( w3_23 ) );
  DFF_X1 u0_w_reg_3_24 (.CK( clk ) , .D( u0_N264 ) , .QN( u0_n248 ) , .Q( w3_24 ) );
  DFF_X1 u0_w_reg_3_25 (.CK( clk ) , .D( u0_N265 ) , .Q( w3_25 ) );
  DFF_X1 u0_w_reg_3_26 (.CK( clk ) , .D( u0_N266 ) , .Q( w3_26 ) );
  DFF_X1 u0_w_reg_3_27 (.CK( clk ) , .D( u0_N267 ) , .Q( w3_27 ) );
  DFF_X1 u0_w_reg_3_28 (.CK( clk ) , .D( u0_N268 ) , .Q( w3_28 ) );
  DFF_X1 u0_w_reg_3_29 (.CK( clk ) , .D( u0_N269 ) , .Q( w3_29 ) );
  DFF_X1 u0_w_reg_3_3 (.CK( clk ) , .D( u0_N243 ) , .Q( w3_3 ) );
  DFF_X1 u0_w_reg_3_30 (.CK( clk ) , .D( u0_N270 ) , .Q( w3_30 ) );
  DFF_X1 u0_w_reg_3_31 (.CK( clk ) , .D( u0_N271 ) , .Q( w3_31 ) );
  DFF_X1 u0_w_reg_3_4 (.CK( clk ) , .D( u0_N244 ) , .Q( w3_4 ) );
  DFF_X1 u0_w_reg_3_5 (.CK( clk ) , .D( u0_N245 ) , .Q( w3_5 ) );
  DFF_X1 u0_w_reg_3_6 (.CK( clk ) , .D( u0_N246 ) , .Q( w3_6 ) );
  DFF_X1 u0_w_reg_3_7 (.CK( clk ) , .D( u0_N247 ) , .Q( w3_7 ) );
  DFF_X1 u0_w_reg_3_8 (.CK( clk ) , .D( u0_N248 ) , .Q( w3_8 ) );
  DFF_X1 u0_w_reg_3_9 (.CK( clk ) , .D( u0_N249 ) , .Q( w3_9 ) );
endmodule
