module aes_aes_die_13 ( u0_n170, w2_27, w3_24, w3_25, w3_26, w3_27, w3_28, w3_29, w3_30, 
       w3_31, u0_n77, u0_n79, u0_subword_0, u0_subword_1, u0_subword_2, u0_subword_3, u0_subword_4, u0_subword_5, u0_subword_6, 
        u0_subword_7 );
  input u0_n170, w2_27, w3_24, w3_25, w3_26, w3_27, w3_28, w3_29, w3_30, 
        w3_31;
  output u0_n77, u0_n79, u0_subword_0, u0_subword_1, u0_subword_2, u0_subword_3, u0_subword_4, u0_subword_5, u0_subword_6, 
        u0_subword_7;
  wire u0_u3_n41, u0_u3_n438, u0_u3_n439, u0_u3_n440, u0_u3_n441, u0_u3_n442, u0_u3_n443, u0_u3_n444, u0_u3_n445, 
       u0_u3_n446, u0_u3_n447, u0_u3_n448, u0_u3_n449, u0_u3_n450, u0_u3_n451, u0_u3_n452, u0_u3_n453, u0_u3_n454, 
       u0_u3_n455, u0_u3_n456, u0_u3_n457, u0_u3_n458, u0_u3_n459, u0_u3_n460, u0_u3_n461, u0_u3_n462, u0_u3_n463, 
       u0_u3_n464, u0_u3_n465, u0_u3_n466, u0_u3_n467, u0_u3_n468, u0_u3_n469, u0_u3_n470, u0_u3_n471, u0_u3_n472, 
       u0_u3_n473, u0_u3_n474, u0_u3_n475, u0_u3_n476, u0_u3_n477, u0_u3_n478, u0_u3_n479, u0_u3_n480, u0_u3_n481, 
       u0_u3_n482, u0_u3_n483, u0_u3_n484, u0_u3_n485, u0_u3_n486, u0_u3_n487, u0_u3_n488, u0_u3_n489, u0_u3_n490, 
       u0_u3_n491, u0_u3_n492, u0_u3_n493, u0_u3_n494, u0_u3_n495, u0_u3_n496, u0_u3_n497, u0_u3_n498, u0_u3_n499, 
       u0_u3_n500, u0_u3_n501, u0_u3_n502, u0_u3_n503, u0_u3_n504, u0_u3_n505, u0_u3_n506, u0_u3_n507, u0_u3_n508, 
       u0_u3_n509, u0_u3_n510, u0_u3_n511, u0_u3_n512, u0_u3_n513, u0_u3_n514, u0_u3_n515, u0_u3_n516, u0_u3_n517, 
       u0_u3_n518, u0_u3_n519, u0_u3_n520, u0_u3_n521, u0_u3_n522, u0_u3_n523, u0_u3_n524, u0_u3_n525, u0_u3_n526, 
       u0_u3_n527, u0_u3_n528, u0_u3_n529, u0_u3_n530, u0_u3_n531, u0_u3_n532, u0_u3_n533, u0_u3_n534, u0_u3_n535, 
       u0_u3_n536, u0_u3_n537, u0_u3_n538, u0_u3_n539, u0_u3_n540, u0_u3_n541, u0_u3_n542, u0_u3_n543, u0_u3_n544, 
       u0_u3_n545, u0_u3_n546, u0_u3_n547, u0_u3_n548, u0_u3_n549, u0_u3_n550, u0_u3_n551, u0_u3_n552, u0_u3_n553, 
       u0_u3_n554, u0_u3_n555, u0_u3_n556, u0_u3_n557, u0_u3_n558, u0_u3_n559, u0_u3_n560, u0_u3_n561, u0_u3_n562, 
       u0_u3_n563, u0_u3_n564, u0_u3_n565, u0_u3_n566, u0_u3_n567, u0_u3_n568, u0_u3_n569, u0_u3_n570, u0_u3_n571, 
       u0_u3_n572, u0_u3_n573, u0_u3_n574, u0_u3_n575, u0_u3_n576, u0_u3_n577, u0_u3_n578, u0_u3_n579, u0_u3_n580, 
       u0_u3_n581, u0_u3_n582, u0_u3_n583, u0_u3_n584, u0_u3_n585, u0_u3_n586, u0_u3_n587, u0_u3_n588, u0_u3_n589, 
       u0_u3_n590, u0_u3_n591, u0_u3_n592, u0_u3_n593, u0_u3_n594, u0_u3_n595, u0_u3_n596, u0_u3_n597, u0_u3_n598, 
       u0_u3_n599, u0_u3_n600, u0_u3_n601, u0_u3_n602, u0_u3_n603, u0_u3_n604, u0_u3_n605, u0_u3_n606, u0_u3_n607, 
       u0_u3_n608, u0_u3_n609, u0_u3_n610, u0_u3_n611, u0_u3_n612, u0_u3_n613, u0_u3_n614, u0_u3_n615, u0_u3_n616, 
       u0_u3_n617, u0_u3_n618, u0_u3_n619, u0_u3_n620, u0_u3_n621, u0_u3_n622, u0_u3_n623, u0_u3_n624, u0_u3_n625, 
       u0_u3_n626, u0_u3_n627, u0_u3_n628, u0_u3_n629, u0_u3_n630, u0_u3_n631, u0_u3_n632, u0_u3_n633, u0_u3_n634, 
       u0_u3_n635, u0_u3_n636, u0_u3_n637, u0_u3_n638, u0_u3_n639, u0_u3_n640, u0_u3_n641, u0_u3_n642, u0_u3_n643, 
       u0_u3_n644, u0_u3_n645, u0_u3_n646, u0_u3_n647, u0_u3_n648, u0_u3_n649, u0_u3_n650, u0_u3_n651, u0_u3_n652, 
       u0_u3_n653, u0_u3_n654, u0_u3_n655, u0_u3_n656, u0_u3_n657, u0_u3_n658, u0_u3_n659, u0_u3_n660, u0_u3_n661, 
       u0_u3_n662, u0_u3_n663, u0_u3_n664, u0_u3_n665, u0_u3_n666, u0_u3_n667, u0_u3_n668, u0_u3_n669, u0_u3_n670, 
       u0_u3_n671, u0_u3_n672, u0_u3_n673, u0_u3_n674, u0_u3_n675, u0_u3_n676, u0_u3_n677, u0_u3_n678, u0_u3_n679, 
       u0_u3_n680, u0_u3_n681, u0_u3_n682, u0_u3_n683, u0_u3_n684, u0_u3_n685, u0_u3_n686, u0_u3_n687, u0_u3_n688, 
       u0_u3_n689, u0_u3_n690, u0_u3_n691, u0_u3_n692, u0_u3_n693, u0_u3_n694, u0_u3_n695, u0_u3_n696, u0_u3_n697, 
       u0_u3_n698, u0_u3_n699, u0_u3_n700, u0_u3_n701, u0_u3_n702, u0_u3_n703, u0_u3_n704, u0_u3_n705, u0_u3_n706, 
       u0_u3_n707, u0_u3_n708, u0_u3_n709, u0_u3_n710, u0_u3_n711, u0_u3_n712, u0_u3_n713, u0_u3_n714, u0_u3_n715, 
       u0_u3_n716, u0_u3_n717, u0_u3_n718, u0_u3_n719, u0_u3_n720, u0_u3_n721, u0_u3_n722, u0_u3_n723, u0_u3_n724, 
       u0_u3_n725, u0_u3_n726, u0_u3_n727, u0_u3_n728, u0_u3_n729, u0_u3_n730, u0_u3_n731, u0_u3_n732, u0_u3_n733, 
       u0_u3_n734, u0_u3_n735, u0_u3_n736, u0_u3_n737, u0_u3_n738, u0_u3_n739, u0_u3_n740, u0_u3_n741, u0_u3_n742, 
       u0_u3_n743, u0_u3_n744, u0_u3_n745, u0_u3_n746, u0_u3_n747, u0_u3_n748, u0_u3_n749, u0_u3_n750, u0_u3_n751, 
       u0_u3_n752, u0_u3_n753, u0_u3_n754, u0_u3_n755, u0_u3_n756, u0_u3_n757, u0_u3_n758, u0_u3_n759, u0_u3_n760, 
       u0_u3_n761, u0_u3_n762, u0_u3_n763, u0_u3_n764, u0_u3_n765, u0_u3_n766, u0_u3_n767, u0_u3_n768, u0_u3_n769, 
       u0_u3_n770, u0_u3_n771, u0_u3_n772, u0_u3_n773, u0_u3_n774, u0_u3_n775, u0_u3_n776, u0_u3_n777, u0_u3_n778, 
       u0_u3_n779, u0_u3_n780, u0_u3_n781, u0_u3_n782, u0_u3_n783, u0_u3_n784, u0_u3_n785, u0_u3_n786, u0_u3_n787, 
       u0_u3_n788, u0_u3_n789, u0_u3_n790, u0_u3_n791, u0_u3_n792, u0_u3_n793, u0_u3_n794, u0_u3_n795, u0_u3_n796, 
       u0_u3_n797, u0_u3_n798, u0_u3_n799, u0_u3_n800, u0_u3_n801, u0_u3_n802, u0_u3_n803, u0_u3_n804, u0_u3_n805, 
       u0_u3_n806, u0_u3_n807, u0_u3_n808, u0_u3_n809, u0_u3_n810, u0_u3_n811, u0_u3_n812, u0_u3_n813, u0_u3_n814, 
       u0_u3_n815, u0_u3_n816, u0_u3_n817, u0_u3_n818, u0_u3_n819, u0_u3_n820, u0_u3_n821, u0_u3_n822, u0_u3_n823, 
       u0_u3_n824, u0_u3_n825, u0_u3_n826, u0_u3_n827, u0_u3_n828, u0_u3_n829, u0_u3_n830, u0_u3_n831, u0_u3_n832, 
       u0_u3_n833, u0_u3_n834, u0_u3_n835, u0_u3_n836, u0_u3_n837, u0_u3_n838, u0_u3_n839, u0_u3_n840, u0_u3_n841, 
       u0_u3_n842, u0_u3_n843, u0_u3_n844, u0_u3_n845, u0_u3_n846, u0_u3_n847, u0_u3_n848, u0_u3_n849, u0_u3_n850, 
       u0_u3_n851, u0_u3_n852, u0_u3_n853, u0_u3_n854, u0_u3_n855, u0_u3_n856, u0_u3_n857, u0_u3_n858, u0_u3_n859, 
       u0_u3_n860, u0_u3_n861, u0_u3_n862, u0_u3_n863, u0_u3_n864, u0_u3_n865, u0_u3_n866, u0_u3_n867, u0_u3_n868, 
       u0_u3_n869, u0_u3_n870, u0_u3_n871, u0_u3_n872, u0_u3_n873, u0_u3_n874, u0_u3_n875, u0_u3_n876, u0_u3_n877, 
        u0_u3_n878;
  XOR2_X1 u0_U295 (.Z( u0_n77 ) , .A( u0_n79 ) , .B( w3_27 ) );
  XOR2_X1 u0_U327 (.A( u0_n170 ) , .Z( u0_n79 ) , .B( w2_27 ) );
  NOR2_X1 u0_u3_U10 (.ZN( u0_u3_n578 ) , .A1( u0_u3_n625 ) , .A2( u0_u3_n748 ) );
  NOR2_X1 u0_u3_U100 (.ZN( u0_u3_n669 ) , .A1( u0_u3_n731 ) , .A2( u0_u3_n806 ) );
  NOR2_X1 u0_u3_U101 (.ZN( u0_u3_n535 ) , .A2( u0_u3_n752 ) , .A1( u0_u3_n753 ) );
  NOR2_X1 u0_u3_U102 (.A2( u0_u3_n711 ) , .A1( u0_u3_n765 ) , .ZN( u0_u3_n797 ) );
  OAI22_X1 u0_u3_U103 (.B1( u0_u3_n493 ) , .ZN( u0_u3_n494 ) , .A1( u0_u3_n689 ) , .A2( u0_u3_n766 ) , .B2( u0_u3_n820 ) );
  NOR3_X1 u0_u3_U104 (.ZN( u0_u3_n493 ) , .A1( u0_u3_n785 ) , .A2( u0_u3_n852 ) , .A3( u0_u3_n865 ) );
  NOR2_X1 u0_u3_U105 (.ZN( u0_u3_n509 ) , .A2( u0_u3_n731 ) , .A1( u0_u3_n765 ) );
  NOR2_X1 u0_u3_U106 (.ZN( u0_u3_n520 ) , .A1( u0_u3_n711 ) , .A2( u0_u3_n806 ) );
  OAI21_X1 u0_u3_U107 (.ZN( u0_u3_n734 ) , .A( u0_u3_n836 ) , .B2( u0_u3_n854 ) , .B1( u0_u3_n875 ) );
  NOR2_X1 u0_u3_U108 (.ZN( u0_u3_n604 ) , .A2( u0_u3_n783 ) , .A1( u0_u3_n806 ) );
  NOR2_X1 u0_u3_U109 (.A2( u0_u3_n711 ) , .A1( u0_u3_n753 ) , .ZN( u0_u3_n774 ) );
  NOR2_X1 u0_u3_U11 (.A1( u0_u3_n681 ) , .ZN( u0_u3_n696 ) , .A2( u0_u3_n810 ) );
  NOR2_X1 u0_u3_U110 (.A2( u0_u3_n438 ) , .ZN( u0_u3_n670 ) , .A1( u0_u3_n753 ) );
  BUF_X2 u0_u3_U111 (.Z( u0_u3_n439 ) , .A( u0_u3_n794 ) );
  OAI21_X1 u0_u3_U112 (.ZN( u0_u3_n790 ) , .A( u0_u3_n841 ) , .B1( u0_u3_n865 ) , .B2( u0_u3_n875 ) );
  BUF_X2 u0_u3_U113 (.Z( u0_u3_n41 ) , .A( u0_u3_n700 ) );
  NOR2_X1 u0_u3_U114 (.ZN( u0_u3_n632 ) , .A2( u0_u3_n731 ) , .A1( u0_u3_n788 ) );
  NOR2_X1 u0_u3_U115 (.ZN( u0_u3_n512 ) , .A1( u0_u3_n732 ) , .A2( u0_u3_n782 ) );
  NOR2_X1 u0_u3_U116 (.ZN( u0_u3_n510 ) , .A1( u0_u3_n815 ) , .A2( u0_u3_n820 ) );
  NOR2_X1 u0_u3_U117 (.ZN( u0_u3_n666 ) , .A1( u0_u3_n732 ) , .A2( u0_u3_n788 ) );
  NOR2_X1 u0_u3_U118 (.ZN( u0_u3_n546 ) , .A2( u0_u3_n711 ) , .A1( u0_u3_n788 ) );
  NOR2_X1 u0_u3_U119 (.ZN( u0_u3_n511 ) , .A2( u0_u3_n783 ) , .A1( u0_u3_n788 ) );
  INV_X1 u0_u3_U12 (.A( u0_u3_n683 ) , .ZN( u0_u3_n842 ) );
  NOR2_X1 u0_u3_U120 (.ZN( u0_u3_n547 ) , .A2( u0_u3_n788 ) , .A1( u0_u3_n795 ) );
  NOR2_X1 u0_u3_U121 (.ZN( u0_u3_n685 ) , .A2( u0_u3_n711 ) , .A1( u0_u3_n820 ) );
  AOI21_X1 u0_u3_U122 (.ZN( u0_u3_n572 ) , .B1( u0_u3_n753 ) , .B2( u0_u3_n765 ) , .A( u0_u3_n783 ) );
  NOR2_X1 u0_u3_U123 (.ZN( u0_u3_n714 ) , .A1( u0_u3_n765 ) , .A2( u0_u3_n766 ) );
  NOR2_X1 u0_u3_U124 (.ZN( u0_u3_n532 ) , .A1( u0_u3_n711 ) , .A2( u0_u3_n782 ) );
  AOI21_X1 u0_u3_U125 (.ZN( u0_u3_n518 ) , .A( u0_u3_n732 ) , .B1( u0_u3_n753 ) , .B2( u0_u3_n806 ) );
  NOR2_X1 u0_u3_U126 (.ZN( u0_u3_n617 ) , .A1( u0_u3_n765 ) , .A2( u0_u3_n815 ) );
  INV_X1 u0_u3_U127 (.A( u0_u3_n753 ) , .ZN( u0_u3_n844 ) );
  AOI21_X1 u0_u3_U128 (.ZN( u0_u3_n594 ) , .B2( u0_u3_n766 ) , .A( u0_u3_n788 ) , .B1( u0_u3_n815 ) );
  AOI21_X1 u0_u3_U129 (.ZN( u0_u3_n517 ) , .A( u0_u3_n782 ) , .B2( u0_u3_n795 ) , .B1( u0_u3_n815 ) );
  INV_X1 u0_u3_U13 (.A( u0_u3_n650 ) , .ZN( u0_u3_n872 ) );
  AOI21_X1 u0_u3_U130 (.B1( u0_u3_n689 ) , .ZN( u0_u3_n690 ) , .A( u0_u3_n731 ) , .B2( u0_u3_n764 ) );
  INV_X1 u0_u3_U131 (.A( u0_u3_n731 ) , .ZN( u0_u3_n854 ) );
  NOR2_X1 u0_u3_U132 (.ZN( u0_u3_n571 ) , .A1( u0_u3_n732 ) , .A2( u0_u3_n765 ) );
  INV_X1 u0_u3_U133 (.A( u0_u3_n795 ) , .ZN( u0_u3_n853 ) );
  NOR2_X1 u0_u3_U134 (.A1( u0_u3_n752 ) , .ZN( u0_u3_n770 ) , .A2( u0_u3_n806 ) );
  NOR2_X1 u0_u3_U135 (.A2( u0_u3_n438 ) , .ZN( u0_u3_n618 ) , .A1( u0_u3_n788 ) );
  AOI211_X1 u0_u3_U136 (.C2( u0_u3_n440 ) , .B( u0_u3_n626 ) , .A( u0_u3_n627 ) , .ZN( u0_u3_n638 ) , .C1( u0_u3_n865 ) );
  NOR4_X1 u0_u3_U137 (.A4( u0_u3_n632 ) , .A3( u0_u3_n633 ) , .A2( u0_u3_n634 ) , .A1( u0_u3_n635 ) , .ZN( u0_u3_n636 ) );
  NOR4_X1 u0_u3_U138 (.A4( u0_u3_n629 ) , .A3( u0_u3_n630 ) , .A2( u0_u3_n631 ) , .ZN( u0_u3_n637 ) , .A1( u0_u3_n667 ) );
  INV_X1 u0_u3_U139 (.A( u0_u3_n783 ) , .ZN( u0_u3_n852 ) );
  NOR4_X1 u0_u3_U14 (.A4( u0_u3_n547 ) , .A3( u0_u3_n548 ) , .A2( u0_u3_n549 ) , .A1( u0_u3_n550 ) , .ZN( u0_u3_n551 ) );
  OAI21_X1 u0_u3_U140 (.A( u0_u3_n701 ) , .ZN( u0_u3_n705 ) , .B2( u0_u3_n753 ) , .B1( u0_u3_n807 ) );
  OAI21_X1 u0_u3_U141 (.ZN( u0_u3_n701 ) , .B2( u0_u3_n836 ) , .B1( u0_u3_n840 ) , .A( u0_u3_n862 ) );
  INV_X1 u0_u3_U142 (.A( u0_u3_n732 ) , .ZN( u0_u3_n870 ) );
  NOR2_X1 u0_u3_U143 (.A2( u0_u3_n440 ) , .ZN( u0_u3_n628 ) , .A1( u0_u3_n841 ) );
  INV_X1 u0_u3_U144 (.A( u0_u3_n766 ) , .ZN( u0_u3_n868 ) );
  NOR2_X1 u0_u3_U145 (.ZN( u0_u3_n473 ) , .A2( u0_u3_n782 ) , .A1( u0_u3_n818 ) );
  INV_X1 u0_u3_U146 (.A( u0_u3_n440 ) , .ZN( u0_u3_n816 ) );
  INV_X1 u0_u3_U147 (.A( u0_u3_n820 ) , .ZN( u0_u3_n846 ) );
  NAND2_X1 u0_u3_U148 (.ZN( u0_u3_n717 ) , .A1( u0_u3_n731 ) , .A2( u0_u3_n783 ) );
  INV_X1 u0_u3_U149 (.A( u0_u3_n788 ) , .ZN( u0_u3_n848 ) );
  NOR4_X1 u0_u3_U15 (.A4( u0_u3_n448 ) , .A3( u0_u3_n449 ) , .A2( u0_u3_n519 ) , .A1( u0_u3_n544 ) , .ZN( u0_u3_n709 ) );
  AOI221_X1 u0_u3_U150 (.A( u0_u3_n767 ) , .ZN( u0_u3_n777 ) , .C2( u0_u3_n813 ) , .B2( u0_u3_n838 ) , .C1( u0_u3_n857 ) , .B1( u0_u3_n868 ) );
  INV_X1 u0_u3_U151 (.A( u0_u3_n764 ) , .ZN( u0_u3_n838 ) );
  AND2_X1 u0_u3_U152 (.ZN( u0_u3_n735 ) , .A1( u0_u3_n782 ) , .A2( u0_u3_n788 ) );
  AOI221_X1 u0_u3_U153 (.A( u0_u3_n453 ) , .ZN( u0_u3_n462 ) , .C2( u0_u3_n756 ) , .B1( u0_u3_n835 ) , .C1( u0_u3_n844 ) , .B2( u0_u3_n863 ) );
  AOI21_X1 u0_u3_U154 (.ZN( u0_u3_n453 ) , .B2( u0_u3_n795 ) , .A( u0_u3_n806 ) , .B1( u0_u3_n818 ) );
  AOI211_X1 u0_u3_U155 (.A( u0_u3_n591 ) , .ZN( u0_u3_n600 ) , .B( u0_u3_n624 ) , .C1( u0_u3_n847 ) , .C2( u0_u3_n857 ) );
  OAI221_X1 u0_u3_U156 (.A( u0_u3_n730 ) , .C2( u0_u3_n731 ) , .B2( u0_u3_n732 ) , .B1( u0_u3_n733 ) , .ZN( u0_u3_n740 ) , .C1( u0_u3_n820 ) );
  NAND2_X1 u0_u3_U157 (.A1( u0_u3_n444 ) , .A2( u0_u3_n467 ) , .ZN( u0_u3_n711 ) );
  NAND2_X1 u0_u3_U158 (.A2( u0_u3_n474 ) , .A1( u0_u3_n475 ) , .ZN( u0_u3_n820 ) );
  NAND2_X1 u0_u3_U159 (.A2( u0_u3_n463 ) , .A1( u0_u3_n468 ) , .ZN( u0_u3_n783 ) );
  OR3_X1 u0_u3_U16 (.ZN( u0_u3_n449 ) , .A1( u0_u3_n531 ) , .A3( u0_u3_n580 ) , .A2( u0_u3_n877 ) );
  NAND2_X1 u0_u3_U160 (.A1( u0_u3_n458 ) , .A2( u0_u3_n474 ) , .ZN( u0_u3_n806 ) );
  NAND2_X1 u0_u3_U161 (.A2( u0_u3_n451 ) , .A1( u0_u3_n463 ) , .ZN( u0_u3_n731 ) );
  NAND2_X1 u0_u3_U162 (.A1( u0_u3_n452 ) , .A2( u0_u3_n467 ) , .ZN( u0_u3_n727 ) );
  NAND2_X1 u0_u3_U163 (.A2( u0_u3_n457 ) , .A1( u0_u3_n475 ) , .ZN( u0_u3_n782 ) );
  NOR2_X1 u0_u3_U164 (.ZN( u0_u3_n456 ) , .A1( u0_u3_n829 ) , .A2( u0_u3_n830 ) );
  NAND2_X1 u0_u3_U165 (.A2( u0_u3_n467 ) , .A1( u0_u3_n468 ) , .ZN( u0_u3_n815 ) );
  NAND2_X1 u0_u3_U166 (.A2( u0_u3_n451 ) , .A1( u0_u3_n455 ) , .ZN( u0_u3_n732 ) );
  NAND2_X1 u0_u3_U167 (.A2( u0_u3_n452 ) , .A1( u0_u3_n455 ) , .ZN( u0_u3_n766 ) );
  NAND2_X1 u0_u3_U168 (.A1( u0_u3_n454 ) , .A2( u0_u3_n474 ) , .ZN( u0_u3_n819 ) );
  NAND2_X1 u0_u3_U169 (.A1( u0_u3_n456 ) , .A2( u0_u3_n464 ) , .ZN( u0_u3_n747 ) );
  OR4_X1 u0_u3_U17 (.A4( u0_u3_n445 ) , .A2( u0_u3_n446 ) , .A1( u0_u3_n447 ) , .ZN( u0_u3_n448 ) , .A3( u0_u3_n556 ) );
  NAND2_X1 u0_u3_U170 (.A2( u0_u3_n444 ) , .A1( u0_u3_n450 ) , .ZN( u0_u3_n787 ) );
  NAND2_X1 u0_u3_U171 (.A1( u0_u3_n454 ) , .A2( u0_u3_n457 ) , .ZN( u0_u3_n817 ) );
  NAND2_X1 u0_u3_U172 (.A1( u0_u3_n450 ) , .A2( u0_u3_n452 ) , .ZN( u0_u3_n808 ) );
  NAND2_X1 u0_u3_U173 (.A2( u0_u3_n456 ) , .A1( u0_u3_n458 ) , .ZN( u0_u3_n809 ) );
  NAND2_X1 u0_u3_U174 (.A1( u0_u3_n450 ) , .A2( u0_u3_n451 ) , .ZN( u0_u3_n789 ) );
  NAND2_X1 u0_u3_U175 (.A2( u0_u3_n464 ) , .A1( u0_u3_n465 ) , .ZN( u0_u3_n750 ) );
  NAND2_X1 u0_u3_U176 (.A1( u0_u3_n465 ) , .A2( u0_u3_n475 ) , .ZN( u0_u3_n791 ) );
  NAND2_X1 u0_u3_U177 (.A2( u0_u3_n457 ) , .A1( u0_u3_n458 ) , .ZN( u0_u3_n733 ) );
  NAND2_X1 u0_u3_U178 (.A1( u0_u3_n454 ) , .A2( u0_u3_n465 ) , .ZN( u0_u3_n793 ) );
  AND2_X1 u0_u3_U179 (.ZN( u0_u3_n440 ) , .A1( u0_u3_n457 ) , .A2( u0_u3_n464 ) );
  INV_X1 u0_u3_U18 (.A( u0_u3_n616 ) , .ZN( u0_u3_n877 ) );
  NOR2_X1 u0_u3_U180 (.ZN( u0_u3_n452 ) , .A1( u0_u3_n850 ) , .A2( w3_28 ) );
  NAND4_X1 u0_u3_U181 (.ZN( u0_subword_1 ) , .A4( u0_u3_n598 ) , .A3( u0_u3_n599 ) , .A2( u0_u3_n600 ) , .A1( u0_u3_n601 ) );
  AOI211_X1 u0_u3_U182 (.B( u0_u3_n592 ) , .A( u0_u3_n593 ) , .ZN( u0_u3_n599 ) , .C2( u0_u3_n814 ) , .C1( u0_u3_n836 ) );
  NOR4_X1 u0_u3_U183 (.A4( u0_u3_n594 ) , .A3( u0_u3_n595 ) , .A2( u0_u3_n596 ) , .A1( u0_u3_n597 ) , .ZN( u0_u3_n598 ) );
  NOR4_X1 u0_u3_U184 (.A4( u0_u3_n737 ) , .A3( u0_u3_n738 ) , .A2( u0_u3_n739 ) , .A1( u0_u3_n740 ) , .ZN( u0_u3_n741 ) );
  AOI211_X1 u0_u3_U185 (.B( u0_u3_n728 ) , .A( u0_u3_n729 ) , .ZN( u0_u3_n742 ) , .C1( u0_u3_n845 ) , .C2( u0_u3_n857 ) );
  AOI222_X1 u0_u3_U186 (.B2( u0_u3_n641 ) , .ZN( u0_u3_n647 ) , .B1( u0_u3_n843 ) , .A1( u0_u3_n844 ) , .C2( u0_u3_n848 ) , .C1( u0_u3_n865 ) , .A2( u0_u3_n867 ) );
  NOR4_X1 u0_u3_U187 (.A4( u0_u3_n642 ) , .A3( u0_u3_n643 ) , .A2( u0_u3_n644 ) , .A1( u0_u3_n645 ) , .ZN( u0_u3_n646 ) );
  AOI221_X1 u0_u3_U188 (.A( u0_u3_n784 ) , .ZN( u0_u3_n801 ) , .C2( u0_u3_n839 ) , .B2( u0_u3_n840 ) , .B1( u0_u3_n867 ) , .C1( u0_u3_n868 ) );
  NOR4_X1 u0_u3_U189 (.A4( u0_u3_n796 ) , .A3( u0_u3_n797 ) , .A2( u0_u3_n798 ) , .A1( u0_u3_n799 ) , .ZN( u0_u3_n800 ) );
  NOR4_X1 u0_u3_U19 (.ZN( u0_u3_n478 ) , .A1( u0_u3_n534 ) , .A3( u0_u3_n571 ) , .A4( u0_u3_n603 ) , .A2( u0_u3_n645 ) );
  NAND4_X1 u0_u3_U190 (.ZN( u0_subword_0 ) , .A4( u0_u3_n504 ) , .A3( u0_u3_n505 ) , .A2( u0_u3_n506 ) , .A1( u0_u3_n507 ) );
  NOR4_X1 u0_u3_U191 (.A4( u0_u3_n501 ) , .A3( u0_u3_n502 ) , .A2( u0_u3_n503 ) , .ZN( u0_u3_n504 ) , .A1( u0_u3_n530 ) );
  AOI221_X1 u0_u3_U192 (.A( u0_u3_n500 ) , .ZN( u0_u3_n505 ) , .B2( u0_u3_n845 ) , .C1( u0_u3_n848 ) , .C2( u0_u3_n862 ) , .B1( u0_u3_n864 ) );
  NOR4_X1 u0_u3_U193 (.A4( u0_u3_n703 ) , .A3( u0_u3_n704 ) , .A2( u0_u3_n705 ) , .A1( u0_u3_n706 ) , .ZN( u0_u3_n707 ) );
  NOR4_X1 u0_u3_U194 (.A3( u0_u3_n758 ) , .A2( u0_u3_n759 ) , .A1( u0_u3_n760 ) , .ZN( u0_u3_n761 ) , .A4( u0_u3_n871 ) );
  AOI211_X1 u0_u3_U195 (.B( u0_u3_n748 ) , .A( u0_u3_n749 ) , .ZN( u0_u3_n762 ) , .C1( u0_u3_n835 ) , .C2( u0_u3_n855 ) );
  NAND4_X1 u0_u3_U196 (.ZN( u0_subword_7 ) , .A4( u0_u3_n825 ) , .A3( u0_u3_n826 ) , .A2( u0_u3_n827 ) , .A1( u0_u3_n828 ) );
  NOR4_X1 u0_u3_U197 (.A4( u0_u3_n821 ) , .A3( u0_u3_n822 ) , .A2( u0_u3_n823 ) , .A1( u0_u3_n824 ) , .ZN( u0_u3_n825 ) );
  NAND2_X1 u0_u3_U198 (.A2( u0_u3_n464 ) , .A1( u0_u3_n474 ) , .ZN( u0_u3_n700 ) );
  NAND2_X1 u0_u3_U199 (.A2( u0_u3_n451 ) , .A1( u0_u3_n467 ) , .ZN( u0_u3_n818 ) );
  INV_X1 u0_u3_U20 (.A( u0_u3_n752 ) , .ZN( u0_u3_n865 ) );
  OAI21_X1 u0_u3_U200 (.B1( u0_u3_n756 ) , .ZN( u0_u3_n757 ) , .A( u0_u3_n847 ) , .B2( u0_u3_n870 ) );
  AOI221_X1 u0_u3_U201 (.A( u0_u3_n567 ) , .C2( u0_u3_n568 ) , .ZN( u0_u3_n577 ) , .B2( u0_u3_n847 ) , .B1( u0_u3_n854 ) , .C1( u0_u3_n855 ) );
  AOI222_X1 u0_u3_U202 (.ZN( u0_u3_n663 ) , .A2( u0_u3_n841 ) , .B1( u0_u3_n843 ) , .C2( u0_u3_n847 ) , .A1( u0_u3_n862 ) , .C1( u0_u3_n865 ) , .B2( u0_u3_n872 ) );
  AOI221_X1 u0_u3_U203 (.A( u0_u3_n713 ) , .ZN( u0_u3_n724 ) , .C2( u0_u3_n846 ) , .B2( u0_u3_n847 ) , .C1( u0_u3_n863 ) , .B1( u0_u3_n864 ) );
  NAND4_X1 u0_u3_U204 (.A4( u0_u3_n538 ) , .A3( u0_u3_n539 ) , .A2( u0_u3_n540 ) , .A1( u0_u3_n541 ) , .ZN( u0_u3_n625 ) );
  NOR4_X1 u0_u3_U205 (.A1( u0_u3_n534 ) , .ZN( u0_u3_n539 ) , .A2( u0_u3_n657 ) , .A4( u0_u3_n671 ) , .A3( u0_u3_n768 ) );
  NAND4_X1 u0_u3_U206 (.A4( u0_u3_n496 ) , .A3( u0_u3_n497 ) , .A1( u0_u3_n498 ) , .ZN( u0_u3_n805 ) , .A2( u0_u3_n869 ) );
  NOR4_X1 u0_u3_U207 (.A2( u0_u3_n494 ) , .A1( u0_u3_n495 ) , .ZN( u0_u3_n496 ) , .A3( u0_u3_n583 ) , .A4( u0_u3_n615 ) );
  NAND2_X1 u0_u3_U208 (.A1( u0_u3_n444 ) , .A2( u0_u3_n463 ) , .ZN( u0_u3_n702 ) );
  NAND2_X1 u0_u3_U209 (.A1( u0_u3_n455 ) , .A2( u0_u3_n468 ) , .ZN( u0_u3_n672 ) );
  AOI222_X1 u0_u3_U21 (.ZN( u0_u3_n566 ) , .B1( u0_u3_n833 ) , .C1( u0_u3_n843 ) , .A2( u0_u3_n845 ) , .A1( u0_u3_n856 ) , .B2( u0_u3_n865 ) , .C2( u0_u3_n875 ) );
  NAND4_X1 u0_u3_U210 (.A4( u0_u3_n563 ) , .A3( u0_u3_n564 ) , .A2( u0_u3_n565 ) , .A1( u0_u3_n566 ) , .ZN( u0_u3_n610 ) );
  NOR4_X1 u0_u3_U211 (.ZN( u0_u3_n564 ) , .A1( u0_u3_n656 ) , .A3( u0_u3_n664 ) , .A4( u0_u3_n688 ) , .A2( u0_u3_n771 ) );
  NOR2_X1 u0_u3_U212 (.ZN( u0_u3_n454 ) , .A1( u0_u3_n831 ) , .A2( u0_u3_n832 ) );
  INV_X1 u0_u3_U213 (.ZN( u0_u3_n831 ) , .A( w3_26 ) );
  NOR2_X1 u0_u3_U214 (.ZN( u0_u3_n710 ) , .A2( u0_u3_n779 ) , .A1( u0_u3_n803 ) );
  OAI21_X1 u0_u3_U215 (.A( u0_u3_n734 ) , .B1( u0_u3_n735 ) , .ZN( u0_u3_n739 ) , .B2( u0_u3_n808 ) );
  AOI21_X1 u0_u3_U216 (.ZN( u0_u3_n653 ) , .A( u0_u3_n782 ) , .B1( u0_u3_n795 ) , .B2( u0_u3_n808 ) );
  INV_X1 u0_u3_U217 (.A( u0_u3_n808 ) , .ZN( u0_u3_n862 ) );
  NOR2_X1 u0_u3_U218 (.ZN( u0_u3_n738 ) , .A2( u0_u3_n806 ) , .A1( u0_u3_n808 ) );
  NAND2_X1 u0_u3_U219 (.ZN( u0_u3_n756 ) , .A1( u0_u3_n766 ) , .A2( u0_u3_n808 ) );
  NOR4_X1 u0_u3_U22 (.ZN( u0_u3_n482 ) , .A1( u0_u3_n523 ) , .A4( u0_u3_n560 ) , .A3( u0_u3_n585 ) , .A2( u0_u3_n633 ) );
  NOR2_X1 u0_u3_U220 (.ZN( u0_u3_n559 ) , .A1( u0_u3_n765 ) , .A2( u0_u3_n808 ) );
  OAI221_X1 u0_u3_U221 (.A( u0_u3_n699 ) , .ZN( u0_u3_n706 ) , .C2( u0_u3_n787 ) , .C1( u0_u3_n788 ) , .B1( u0_u3_n789 ) , .B2( u0_u3_n809 ) );
  OAI222_X1 u0_u3_U222 (.B1( u0_u3_n41 ) , .ZN( u0_u3_n620 ) , .C1( u0_u3_n727 ) , .C2( u0_u3_n750 ) , .B2( u0_u3_n789 ) , .A2( u0_u3_n795 ) , .A1( u0_u3_n819 ) );
  NAND2_X1 u0_u3_U223 (.A2( u0_u3_n444 ) , .A1( u0_u3_n455 ) , .ZN( u0_u3_n794 ) );
  OAI222_X1 u0_u3_U224 (.B2( u0_u3_n711 ) , .ZN( u0_u3_n712 ) , .C2( u0_u3_n727 ) , .B1( u0_u3_n750 ) , .A1( u0_u3_n809 ) , .C1( u0_u3_n817 ) , .A2( u0_u3_n818 ) );
  INV_X1 u0_u3_U225 (.A( u0_u3_n675 ) , .ZN( u0_u3_n861 ) );
  NOR2_X1 u0_u3_U226 (.ZN( u0_u3_n531 ) , .A2( u0_u3_n727 ) , .A1( u0_u3_n806 ) );
  NOR2_X1 u0_u3_U227 (.ZN( u0_u3_n529 ) , .A1( u0_u3_n727 ) , .A2( u0_u3_n753 ) );
  INV_X1 u0_u3_U228 (.A( u0_u3_n727 ) , .ZN( u0_u3_n858 ) );
  NOR2_X1 u0_u3_U229 (.ZN( u0_u3_n450 ) , .A2( u0_u3_n851 ) , .A1( u0_u3_n860 ) );
  NOR4_X1 u0_u3_U23 (.A4( u0_u3_n559 ) , .A3( u0_u3_n560 ) , .A2( u0_u3_n561 ) , .A1( u0_u3_n562 ) , .ZN( u0_u3_n563 ) );
  AOI222_X1 u0_u3_U230 (.ZN( u0_u3_n528 ) , .A1( u0_u3_n837 ) , .B2( u0_u3_n839 ) , .C1( u0_u3_n846 ) , .C2( u0_u3_n852 ) , .A2( u0_u3_n854 ) , .B1( u0_u3_n868 ) );
  NOR3_X1 u0_u3_U231 (.A2( u0_u3_n440 ) , .ZN( u0_u3_n443 ) , .A3( u0_u3_n839 ) , .A1( u0_u3_n848 ) );
  NAND2_X1 u0_u3_U232 (.ZN( u0_u3_n616 ) , .A2( u0_u3_n839 ) , .A1( u0_u3_n875 ) );
  NOR2_X1 u0_u3_U233 (.ZN( u0_u3_n498 ) , .A1( u0_u3_n681 ) , .A2( u0_u3_n697 ) );
  AOI211_X1 u0_u3_U234 (.B( u0_u3_n697 ) , .A( u0_u3_n698 ) , .ZN( u0_u3_n708 ) , .C2( u0_u3_n834 ) , .C1( u0_u3_n853 ) );
  NOR2_X1 u0_u3_U235 (.ZN( u0_u3_n586 ) , .A1( u0_u3_n795 ) , .A2( u0_u3_n820 ) );
  AOI21_X1 u0_u3_U236 (.ZN( u0_u3_n543 ) , .A( u0_u3_n766 ) , .B2( u0_u3_n782 ) , .B1( u0_u3_n820 ) );
  NOR2_X1 u0_u3_U237 (.ZN( u0_u3_n612 ) , .A2( u0_u3_n727 ) , .A1( u0_u3_n820 ) );
  NOR2_X1 u0_u3_U238 (.ZN( u0_u3_n718 ) , .A1( u0_u3_n808 ) , .A2( u0_u3_n820 ) );
  OAI21_X1 u0_u3_U239 (.A( u0_u3_n790 ) , .B2( u0_u3_n791 ) , .B1( u0_u3_n792 ) , .ZN( u0_u3_n798 ) );
  NOR4_X1 u0_u3_U24 (.A4( u0_u3_n555 ) , .A3( u0_u3_n556 ) , .A2( u0_u3_n557 ) , .A1( u0_u3_n558 ) , .ZN( u0_u3_n565 ) );
  AOI21_X1 u0_u3_U240 (.ZN( u0_u3_n642 ) , .B2( u0_u3_n752 ) , .A( u0_u3_n791 ) , .B1( u0_u3_n815 ) );
  AOI21_X1 u0_u3_U241 (.A( u0_u3_n736 ) , .ZN( u0_u3_n737 ) , .B2( u0_u3_n783 ) , .B1( u0_u3_n795 ) );
  AOI21_X1 u0_u3_U242 (.B2( u0_u3_n766 ) , .ZN( u0_u3_n767 ) , .A( u0_u3_n791 ) , .B1( u0_u3_n795 ) );
  NOR2_X1 u0_u3_U243 (.ZN( u0_u3_n521 ) , .A1( u0_u3_n711 ) , .A2( u0_u3_n791 ) );
  NOR2_X1 u0_u3_U244 (.ZN( u0_u3_n487 ) , .A1( u0_u3_n791 ) , .A2( u0_u3_n808 ) );
  NOR2_X1 u0_u3_U245 (.ZN( u0_u3_n537 ) , .A1( u0_u3_n727 ) , .A2( u0_u3_n791 ) );
  INV_X1 u0_u3_U246 (.A( u0_u3_n791 ) , .ZN( u0_u3_n847 ) );
  OAI22_X1 u0_u3_U247 (.B2( u0_u3_n782 ) , .B1( u0_u3_n783 ) , .ZN( u0_u3_n784 ) , .A2( u0_u3_n817 ) , .A1( u0_u3_n818 ) );
  AOI21_X1 u0_u3_U248 (.ZN( u0_u3_n501 ) , .A( u0_u3_n727 ) , .B2( u0_u3_n765 ) , .B1( u0_u3_n817 ) );
  NAND4_X1 u0_u3_U249 (.A4( u0_u3_n482 ) , .A3( u0_u3_n483 ) , .A2( u0_u3_n484 ) , .A1( u0_u3_n485 ) , .ZN( u0_u3_n697 ) );
  NOR4_X1 u0_u3_U25 (.A4( u0_u3_n771 ) , .A3( u0_u3_n772 ) , .A2( u0_u3_n773 ) , .A1( u0_u3_n774 ) , .ZN( u0_u3_n775 ) );
  AOI21_X1 u0_u3_U250 (.ZN( u0_u3_n542 ) , .B2( u0_u3_n815 ) , .A( u0_u3_n817 ) , .B1( u0_u3_n818 ) );
  NOR2_X1 u0_u3_U251 (.ZN( u0_u3_n523 ) , .A2( u0_u3_n711 ) , .A1( u0_u3_n817 ) );
  NOR2_X1 u0_u3_U252 (.ZN( u0_u3_n549 ) , .A2( u0_u3_n783 ) , .A1( u0_u3_n817 ) );
  INV_X1 u0_u3_U253 (.A( u0_u3_n817 ) , .ZN( u0_u3_n836 ) );
  NOR2_X1 u0_u3_U254 (.ZN( u0_u3_n548 ) , .A1( u0_u3_n752 ) , .A2( u0_u3_n817 ) );
  NOR2_X1 u0_u3_U255 (.ZN( u0_u3_n560 ) , .A1( u0_u3_n795 ) , .A2( u0_u3_n817 ) );
  AOI21_X1 u0_u3_U256 (.A( u0_u3_n673 ) , .B1( u0_u3_n674 ) , .ZN( u0_u3_n675 ) , .B2( u0_u3_n858 ) );
  AOI22_X1 u0_u3_U257 (.A2( u0_u3_n785 ) , .ZN( u0_u3_n786 ) , .B2( u0_u3_n834 ) , .A1( u0_u3_n837 ) , .B1( u0_u3_n865 ) );
  AOI21_X1 u0_u3_U258 (.ZN( u0_u3_n643 ) , .B2( u0_u3_n750 ) , .A( u0_u3_n795 ) , .B1( u0_u3_n806 ) );
  NAND4_X1 u0_u3_U259 (.A4( u0_u3_n775 ) , .A3( u0_u3_n776 ) , .A2( u0_u3_n777 ) , .A1( u0_u3_n778 ) , .ZN( u0_u3_n804 ) );
  NOR3_X1 u0_u3_U26 (.A3( u0_u3_n768 ) , .A2( u0_u3_n769 ) , .A1( u0_u3_n770 ) , .ZN( u0_u3_n776 ) );
  OAI21_X1 u0_u3_U260 (.ZN( u0_u3_n466 ) , .B1( u0_u3_n812 ) , .A( u0_u3_n837 ) , .B2( u0_u3_n853 ) );
  NOR2_X1 u0_u3_U261 (.ZN( u0_u3_n659 ) , .A1( u0_u3_n750 ) , .A2( u0_u3_n783 ) );
  NOR2_X1 u0_u3_U262 (.ZN( u0_u3_n683 ) , .A2( u0_u3_n837 ) , .A1( u0_u3_n841 ) );
  NOR2_X1 u0_u3_U263 (.ZN( u0_u3_n764 ) , .A1( u0_u3_n836 ) , .A2( u0_u3_n837 ) );
  NOR2_X1 u0_u3_U264 (.ZN( u0_u3_n570 ) , .A1( u0_u3_n750 ) , .A2( u0_u3_n808 ) );
  NOR2_X1 u0_u3_U265 (.A2( u0_u3_n438 ) , .ZN( u0_u3_n633 ) , .A1( u0_u3_n750 ) );
  INV_X1 u0_u3_U266 (.A( u0_u3_n750 ) , .ZN( u0_u3_n837 ) );
  NOR4_X1 u0_u3_U267 (.ZN( u0_u3_n488 ) , .A2( u0_u3_n536 ) , .A1( u0_u3_n561 ) , .A3( u0_u3_n634 ) , .A4( u0_u3_n721 ) );
  NAND4_X1 u0_u3_U268 (.A4( u0_u3_n488 ) , .A3( u0_u3_n489 ) , .A2( u0_u3_n490 ) , .A1( u0_u3_n491 ) , .ZN( u0_u3_n781 ) );
  AOI21_X1 u0_u3_U269 (.B1( u0_u3_n438 ) , .ZN( u0_u3_n592 ) , .B2( u0_u3_n702 ) , .A( u0_u3_n820 ) );
  NAND4_X1 u0_u3_U27 (.A4( u0_u3_n606 ) , .A3( u0_u3_n607 ) , .A2( u0_u3_n608 ) , .A1( u0_u3_n609 ) , .ZN( u0_u3_n725 ) );
  AOI21_X1 u0_u3_U270 (.B1( u0_u3_n702 ) , .ZN( u0_u3_n703 ) , .A( u0_u3_n735 ) , .B2( u0_u3_n766 ) );
  INV_X1 u0_u3_U271 (.A( u0_u3_n702 ) , .ZN( u0_u3_n855 ) );
  AOI21_X1 u0_u3_U272 (.ZN( u0_u3_n445 ) , .A( u0_u3_n702 ) , .B1( u0_u3_n736 ) , .B2( u0_u3_n753 ) );
  NOR2_X1 u0_u3_U273 (.ZN( u0_u3_n686 ) , .A2( u0_u3_n702 ) , .A1( u0_u3_n806 ) );
  NOR2_X1 u0_u3_U274 (.ZN( u0_u3_n580 ) , .A2( u0_u3_n702 ) , .A1( u0_u3_n817 ) );
  NAND2_X1 u0_u3_U275 (.A1( u0_u3_n702 ) , .A2( u0_u3_n732 ) , .ZN( u0_u3_n785 ) );
  NOR3_X1 u0_u3_U276 (.A3( u0_u3_n744 ) , .A2( u0_u3_n745 ) , .A1( u0_u3_n746 ) , .ZN( u0_u3_n763 ) );
  OAI22_X1 u0_u3_U277 (.ZN( u0_u3_n492 ) , .A1( u0_u3_n727 ) , .B2( u0_u3_n731 ) , .B1( u0_u3_n733 ) , .A2( u0_u3_n782 ) );
  NOR2_X1 u0_u3_U278 (.ZN( u0_u3_n582 ) , .A2( u0_u3_n711 ) , .A1( u0_u3_n733 ) );
  NOR2_X1 u0_u3_U279 (.ZN( u0_u3_n536 ) , .A2( u0_u3_n727 ) , .A1( u0_u3_n733 ) );
  NOR3_X1 u0_u3_U28 (.A1( u0_u3_n602 ) , .ZN( u0_u3_n607 ) , .A3( u0_u3_n666 ) , .A2( u0_u3_n773 ) );
  AOI222_X1 u0_u3_U280 (.ZN( u0_u3_n608 ) , .B2( u0_u3_n674 ) , .B1( u0_u3_n756 ) , .C2( u0_u3_n834 ) , .A1( u0_u3_n836 ) , .A2( u0_u3_n864 ) , .C1( u0_u3_n865 ) );
  AOI221_X1 u0_u3_U281 (.A( u0_u3_n486 ) , .ZN( u0_u3_n491 ) , .B1( u0_u3_n834 ) , .C2( u0_u3_n846 ) , .C1( u0_u3_n854 ) , .B2( u0_u3_n864 ) );
  NOR2_X1 u0_u3_U282 (.ZN( u0_u3_n792 ) , .A2( u0_u3_n864 ) , .A1( u0_u3_n870 ) );
  NOR2_X1 u0_u3_U283 (.ZN( u0_u3_n464 ) , .A1( u0_u3_n832 ) , .A2( w3_26 ) );
  NOR2_X1 u0_u3_U284 (.ZN( u0_u3_n474 ) , .A1( u0_u3_n829 ) , .A2( w3_25 ) );
  AOI21_X1 u0_u3_U285 (.A( u0_u3_n439 ) , .ZN( u0_u3_n644 ) , .B1( u0_u3_n683 ) , .B2( u0_u3_n820 ) );
  AOI21_X1 u0_u3_U286 (.B2( u0_u3_n439 ) , .ZN( u0_u3_n500 ) , .A( u0_u3_n782 ) , .B1( u0_u3_n807 ) );
  OAI22_X1 u0_u3_U287 (.B1( u0_u3_n439 ) , .ZN( u0_u3_n698 ) , .A2( u0_u3_n733 ) , .A1( u0_u3_n783 ) , .B2( u0_u3_n820 ) );
  AOI21_X1 u0_u3_U288 (.B2( u0_u3_n439 ) , .ZN( u0_u3_n567 ) , .B1( u0_u3_n727 ) , .A( u0_u3_n782 ) );
  AOI21_X1 u0_u3_U289 (.B2( u0_u3_n439 ) , .ZN( u0_u3_n446 ) , .B1( u0_u3_n792 ) , .A( u0_u3_n817 ) );
  NOR4_X1 u0_u3_U29 (.A3( u0_u3_n603 ) , .A2( u0_u3_n604 ) , .A1( u0_u3_n605 ) , .ZN( u0_u3_n606 ) , .A4( u0_u3_n658 ) );
  NOR2_X1 u0_u3_U290 (.A2( u0_u3_n439 ) , .ZN( u0_u3_n667 ) , .A1( u0_u3_n788 ) );
  NOR2_X1 u0_u3_U291 (.A2( u0_u3_n439 ) , .ZN( u0_u3_n558 ) , .A1( u0_u3_n753 ) );
  NOR2_X1 u0_u3_U292 (.A2( u0_u3_n439 ) , .ZN( u0_u3_n562 ) , .A1( u0_u3_n806 ) );
  NOR2_X1 u0_u3_U293 (.A1( u0_u3_n439 ) , .ZN( u0_u3_n645 ) , .A2( u0_u3_n791 ) );
  NOR2_X1 u0_u3_U294 (.A2( u0_u3_n439 ) , .ZN( u0_u3_n545 ) , .A1( u0_u3_n765 ) );
  INV_X1 u0_u3_U295 (.A( u0_u3_n794 ) , .ZN( u0_u3_n875 ) );
  NOR2_X1 u0_u3_U296 (.ZN( u0_u3_n463 ) , .A1( u0_u3_n851 ) , .A2( w3_31 ) );
  AOI21_X1 u0_u3_U297 (.B2( u0_u3_n439 ) , .A( u0_u3_n793 ) , .B1( u0_u3_n795 ) , .ZN( u0_u3_n796 ) );
  AOI222_X1 u0_u3_U298 (.C2( u0_u3_n812 ) , .B2( u0_u3_n813 ) , .A2( u0_u3_n814 ) , .ZN( u0_u3_n826 ) , .C1( u0_u3_n835 ) , .A1( u0_u3_n841 ) , .B1( u0_u3_n855 ) );
  AOI22_X1 u0_u3_U299 (.ZN( u0_u3_n730 ) , .B1( u0_u3_n835 ) , .A2( u0_u3_n840 ) , .A1( u0_u3_n865 ) , .B2( u0_u3_n868 ) );
  BUF_X1 u0_u3_U3 (.Z( u0_u3_n438 ) , .A( u0_u3_n818 ) );
  NOR4_X1 u0_u3_U30 (.A4( u0_u3_n487 ) , .ZN( u0_u3_n490 ) , .A1( u0_u3_n569 ) , .A2( u0_u3_n584 ) , .A3( u0_u3_n605 ) );
  AOI222_X1 u0_u3_U300 (.ZN( u0_u3_n516 ) , .C1( u0_u3_n835 ) , .B2( u0_u3_n839 ) , .A2( u0_u3_n845 ) , .C2( u0_u3_n864 ) , .B1( u0_u3_n865 ) , .A1( u0_u3_n868 ) );
  AOI222_X1 u0_u3_U301 (.ZN( u0_u3_n472 ) , .B1( u0_u3_n835 ) , .A1( u0_u3_n841 ) , .C1( u0_u3_n844 ) , .C2( u0_u3_n853 ) , .A2( u0_u3_n857 ) , .B2( u0_u3_n867 ) );
  NOR2_X1 u0_u3_U302 (.A2( u0_u3_n438 ) , .ZN( u0_u3_n658 ) , .A1( u0_u3_n793 ) );
  NOR2_X1 u0_u3_U303 (.ZN( u0_u3_n715 ) , .A2( u0_u3_n727 ) , .A1( u0_u3_n793 ) );
  NOR2_X1 u0_u3_U304 (.ZN( u0_u3_n689 ) , .A1( u0_u3_n834 ) , .A2( u0_u3_n835 ) );
  NOR2_X1 u0_u3_U305 (.ZN( u0_u3_n524 ) , .A1( u0_u3_n793 ) , .A2( u0_u3_n815 ) );
  NOR2_X1 u0_u3_U306 (.ZN( u0_u3_n664 ) , .A1( u0_u3_n732 ) , .A2( u0_u3_n793 ) );
  NOR2_X1 u0_u3_U307 (.ZN( u0_u3_n736 ) , .A2( u0_u3_n835 ) , .A1( u0_u3_n847 ) );
  NOR2_X1 u0_u3_U308 (.ZN( u0_u3_n671 ) , .A2( u0_u3_n711 ) , .A1( u0_u3_n793 ) );
  NOR2_X1 u0_u3_U309 (.ZN( u0_u3_n673 ) , .A1( u0_u3_n793 ) , .A2( u0_u3_n808 ) );
  NOR4_X1 u0_u3_U31 (.ZN( u0_u3_n489 ) , .A1( u0_u3_n510 ) , .A2( u0_u3_n522 ) , .A4( u0_u3_n549 ) , .A3( u0_u3_n614 ) );
  INV_X1 u0_u3_U310 (.A( u0_u3_n793 ) , .ZN( u0_u3_n835 ) );
  AOI21_X1 u0_u3_U311 (.B1( u0_u3_n438 ) , .ZN( u0_u3_n513 ) , .B2( u0_u3_n672 ) , .A( u0_u3_n733 ) );
  AOI21_X1 u0_u3_U312 (.B1( u0_u3_n439 ) , .ZN( u0_u3_n629 ) , .B2( u0_u3_n672 ) , .A( u0_u3_n793 ) );
  INV_X1 u0_u3_U313 (.A( u0_u3_n672 ) , .ZN( u0_u3_n867 ) );
  NOR2_X1 u0_u3_U314 (.ZN( u0_u3_n655 ) , .A1( u0_u3_n672 ) , .A2( u0_u3_n817 ) );
  NOR2_X1 u0_u3_U315 (.ZN( u0_u3_n631 ) , .A2( u0_u3_n672 ) , .A1( u0_u3_n788 ) );
  NOR2_X1 u0_u3_U316 (.ZN( u0_u3_n605 ) , .A1( u0_u3_n672 ) , .A2( u0_u3_n806 ) );
  NOR2_X1 u0_u3_U317 (.ZN( u0_u3_n530 ) , .A1( u0_u3_n672 ) , .A2( u0_u3_n782 ) );
  NOR2_X1 u0_u3_U318 (.ZN( u0_u3_n584 ) , .A1( u0_u3_n672 ) , .A2( u0_u3_n791 ) );
  NOR2_X1 u0_u3_U319 (.ZN( u0_u3_n444 ) , .A2( w3_28 ) , .A1( w3_29 ) );
  NOR4_X1 u0_u3_U32 (.A4( u0_u3_n529 ) , .A2( u0_u3_n530 ) , .A1( u0_u3_n531 ) , .ZN( u0_u3_n541 ) , .A3( u0_u3_n704 ) );
  NOR2_X1 u0_u3_U320 (.ZN( u0_u3_n468 ) , .A2( u0_u3_n849 ) , .A1( u0_u3_n850 ) );
  OAI222_X1 u0_u3_U321 (.B2( u0_u3_n750 ) , .B1( u0_u3_n751 ) , .A2( u0_u3_n752 ) , .ZN( u0_u3_n760 ) , .C2( u0_u3_n808 ) , .C1( u0_u3_n817 ) , .A1( u0_u3_n820 ) );
  INV_X1 u0_u3_U322 (.A( u0_u3_n789 ) , .ZN( u0_u3_n864 ) );
  NOR4_X1 u0_u3_U323 (.A4( u0_u3_n617 ) , .A3( u0_u3_n618 ) , .A1( u0_u3_n619 ) , .A2( u0_u3_n620 ) , .ZN( u0_u3_n621 ) );
  INV_X1 u0_u3_U324 (.ZN( u0_u3_n830 ) , .A( w3_25 ) );
  OAI22_X1 u0_u3_U325 (.B2( u0_u3_n753 ) , .B1( u0_u3_n754 ) , .A1( u0_u3_n755 ) , .ZN( u0_u3_n759 ) , .A2( u0_u3_n809 ) );
  OAI22_X1 u0_u3_U326 (.B2( u0_u3_n806 ) , .B1( u0_u3_n807 ) , .A2( u0_u3_n808 ) , .A1( u0_u3_n809 ) , .ZN( u0_u3_n811 ) );
  AOI21_X1 u0_u3_U327 (.ZN( u0_u3_n692 ) , .B2( u0_u3_n752 ) , .B1( u0_u3_n766 ) , .A( u0_u3_n809 ) );
  NAND2_X1 u0_u3_U328 (.A2( u0_u3_n765 ) , .A1( u0_u3_n809 ) , .ZN( u0_u3_n813 ) );
  NOR2_X1 u0_u3_U329 (.ZN( u0_u3_n573 ) , .A1( u0_u3_n731 ) , .A2( u0_u3_n809 ) );
  NOR4_X1 u0_u3_U33 (.A4( u0_u3_n535 ) , .A3( u0_u3_n536 ) , .A2( u0_u3_n537 ) , .ZN( u0_u3_n538 ) , .A1( u0_u3_n823 ) );
  NOR2_X1 u0_u3_U330 (.ZN( u0_u3_n614 ) , .A2( u0_u3_n783 ) , .A1( u0_u3_n809 ) );
  OAI22_X1 u0_u3_U331 (.ZN( u0_u3_n486 ) , .A1( u0_u3_n711 ) , .B2( u0_u3_n788 ) , .A2( u0_u3_n809 ) , .B1( u0_u3_n815 ) );
  AOI21_X1 u0_u3_U332 (.ZN( u0_u3_n480 ) , .A( u0_u3_n672 ) , .B1( u0_u3_n753 ) , .B2( u0_u3_n809 ) );
  INV_X1 u0_u3_U333 (.A( u0_u3_n809 ) , .ZN( u0_u3_n843 ) );
  OAI221_X1 u0_u3_U334 (.A( u0_u3_n786 ) , .C2( u0_u3_n787 ) , .B2( u0_u3_n788 ) , .B1( u0_u3_n789 ) , .ZN( u0_u3_n799 ) , .C1( u0_u3_n816 ) );
  NAND2_X1 u0_u3_U335 (.A1( u0_u3_n732 ) , .A2( u0_u3_n787 ) , .ZN( u0_u3_n814 ) );
  OAI22_X1 u0_u3_U336 (.ZN( u0_u3_n591 ) , .A2( u0_u3_n750 ) , .B2( u0_u3_n765 ) , .A1( u0_u3_n766 ) , .B1( u0_u3_n787 ) );
  AOI21_X1 u0_u3_U337 (.ZN( u0_u3_n595 ) , .B1( u0_u3_n731 ) , .B2( u0_u3_n787 ) , .A( u0_u3_n793 ) );
  NOR2_X1 u0_u3_U338 (.ZN( u0_u3_n807 ) , .A1( u0_u3_n856 ) , .A2( u0_u3_n863 ) );
  AOI21_X1 u0_u3_U339 (.ZN( u0_u3_n626 ) , .B1( u0_u3_n702 ) , .A( u0_u3_n782 ) , .B2( u0_u3_n787 ) );
  NOR4_X1 u0_u3_U34 (.A4( u0_u3_n532 ) , .A3( u0_u3_n533 ) , .ZN( u0_u3_n540 ) , .A2( u0_u3_n687 ) , .A1( u0_u3_n797 ) );
  NAND2_X2 u0_u3_U340 (.A1( u0_u3_n458 ) , .A2( u0_u3_n465 ) , .ZN( u0_u3_n753 ) );
  AOI222_X1 u0_u3_U341 (.ZN( u0_u3_n778 ) , .A1( u0_u3_n833 ) , .C1( u0_u3_n837 ) , .B2( u0_u3_n843 ) , .A2( u0_u3_n852 ) , .B1( u0_u3_n863 ) , .C2( u0_u3_n875 ) );
  AOI222_X1 u0_u3_U342 (.ZN( u0_u3_n609 ) , .A1( u0_u3_n833 ) , .C2( u0_u3_n839 ) , .B1( u0_u3_n844 ) , .A2( u0_u3_n858 ) , .B2( u0_u3_n863 ) , .C1( u0_u3_n870 ) );
  AOI21_X1 u0_u3_U343 (.ZN( u0_u3_n651 ) , .A( u0_u3_n765 ) , .B2( u0_u3_n787 ) , .B1( u0_u3_n795 ) );
  OAI22_X1 u0_u3_U344 (.ZN( u0_u3_n684 ) , .A1( u0_u3_n702 ) , .A2( u0_u3_n733 ) , .B2( u0_u3_n787 ) , .B1( u0_u3_n820 ) );
  NOR2_X1 u0_u3_U345 (.ZN( u0_u3_n654 ) , .A1( u0_u3_n787 ) , .A2( u0_u3_n791 ) );
  NOR2_X1 u0_u3_U346 (.ZN( u0_u3_n751 ) , .A1( u0_u3_n863 ) , .A2( u0_u3_n864 ) );
  NOR2_X1 u0_u3_U347 (.ZN( u0_u3_n455 ) , .A1( u0_u3_n860 ) , .A2( w3_30 ) );
  NOR2_X1 u0_u3_U348 (.ZN( u0_u3_n467 ) , .A2( w3_30 ) , .A1( w3_31 ) );
  AND2_X1 u0_u3_U349 (.ZN( u0_u3_n441 ) , .A2( u0_u3_n834 ) , .A1( u0_u3_n856 ) );
  NOR3_X1 u0_u3_U35 (.A3( u0_u3_n803 ) , .A2( u0_u3_n804 ) , .A1( u0_u3_n805 ) , .ZN( u0_u3_n828 ) );
  AND2_X1 u0_u3_U350 (.ZN( u0_u3_n442 ) , .A2( u0_u3_n845 ) , .A1( u0_u3_n863 ) );
  NOR3_X1 u0_u3_U351 (.A3( u0_u3_n441 ) , .A2( u0_u3_n442 ) , .A1( u0_u3_n579 ) , .ZN( u0_u3_n590 ) );
  INV_X1 u0_u3_U352 (.A( u0_u3_n815 ) , .ZN( u0_u3_n856 ) );
  INV_X1 u0_u3_U353 (.A( u0_u3_n787 ) , .ZN( u0_u3_n863 ) );
  INV_X1 u0_u3_U354 (.A( u0_u3_n806 ) , .ZN( u0_u3_n845 ) );
  INV_X1 u0_u3_U355 (.A( u0_u3_n41 ) , .ZN( u0_u3_n840 ) );
  NOR2_X1 u0_u3_U356 (.A1( u0_u3_n41 ) , .ZN( u0_u3_n773 ) , .A2( u0_u3_n818 ) );
  AOI21_X1 u0_u3_U357 (.B2( u0_u3_n41 ) , .ZN( u0_u3_n574 ) , .B1( u0_u3_n809 ) , .A( u0_u3_n815 ) );
  NOR2_X1 u0_u3_U358 (.A2( u0_u3_n41 ) , .ZN( u0_u3_n665 ) , .A1( u0_u3_n732 ) );
  NOR2_X1 u0_u3_U359 (.A2( u0_u3_n41 ) , .ZN( u0_u3_n635 ) , .A1( u0_u3_n727 ) );
  NAND4_X1 u0_u3_U36 (.A4( u0_u3_n660 ) , .A3( u0_u3_n661 ) , .A2( u0_u3_n662 ) , .A1( u0_u3_n663 ) , .ZN( u0_u3_n803 ) );
  NOR2_X1 u0_u3_U360 (.A2( u0_u3_n41 ) , .A1( u0_u3_n783 ) , .ZN( u0_u3_n823 ) );
  AOI21_X1 u0_u3_U361 (.B2( u0_u3_n41 ) , .ZN( u0_u3_n481 ) , .A( u0_u3_n752 ) , .B1( u0_u3_n782 ) );
  NOR2_X1 u0_u3_U362 (.A2( u0_u3_n41 ) , .ZN( u0_u3_n569 ) , .A1( u0_u3_n766 ) );
  NOR2_X1 u0_u3_U363 (.A2( u0_u3_n41 ) , .ZN( u0_u3_n719 ) , .A1( u0_u3_n795 ) );
  NOR2_X1 u0_u3_U364 (.A2( u0_u3_n41 ) , .ZN( u0_u3_n597 ) , .A1( u0_u3_n731 ) );
  AOI21_X1 u0_u3_U365 (.A( u0_u3_n41 ) , .ZN( u0_u3_n555 ) , .B1( u0_u3_n672 ) , .B2( u0_u3_n808 ) );
  NOR2_X1 u0_u3_U366 (.A2( u0_u3_n41 ) , .ZN( u0_u3_n544 ) , .A1( u0_u3_n702 ) );
  NOR2_X1 u0_u3_U367 (.ZN( u0_u3_n583 ) , .A2( u0_u3_n700 ) , .A1( u0_u3_n794 ) );
  NOR4_X1 u0_u3_U368 (.A4( u0_u3_n779 ) , .A3( u0_u3_n780 ) , .A1( u0_u3_n781 ) , .ZN( u0_u3_n802 ) , .A2( u0_u3_n804 ) );
  NAND4_X1 u0_u3_U369 (.A4( u0_u3_n694 ) , .A3( u0_u3_n695 ) , .A1( u0_u3_n696 ) , .ZN( u0_u3_n779 ) , .A2( u0_u3_n874 ) );
  NOR3_X1 u0_u3_U37 (.A3( u0_u3_n654 ) , .A2( u0_u3_n655 ) , .A1( u0_u3_n656 ) , .ZN( u0_u3_n661 ) );
  AOI21_X1 u0_u3_U370 (.ZN( u0_u3_n596 ) , .B1( u0_u3_n753 ) , .A( u0_u3_n795 ) , .B2( u0_u3_n816 ) );
  AOI21_X1 u0_u3_U371 (.A( u0_u3_n815 ) , .B2( u0_u3_n816 ) , .B1( u0_u3_n817 ) , .ZN( u0_u3_n822 ) );
  OAI222_X1 u0_u3_U372 (.ZN( u0_u3_n508 ) , .C2( u0_u3_n628 ) , .B2( u0_u3_n650 ) , .B1( u0_u3_n750 ) , .A2( u0_u3_n751 ) , .C1( u0_u3_n808 ) , .A1( u0_u3_n809 ) );
  AOI21_X1 u0_u3_U373 (.B1( u0_u3_n628 ) , .ZN( u0_u3_n630 ) , .A( u0_u3_n766 ) , .B2( u0_u3_n817 ) );
  AOI21_X1 u0_u3_U374 (.ZN( u0_u3_n652 ) , .B1( u0_u3_n732 ) , .B2( u0_u3_n766 ) , .A( u0_u3_n816 ) );
  OAI21_X1 u0_u3_U375 (.A( u0_u3_n616 ) , .ZN( u0_u3_n619 ) , .B1( u0_u3_n628 ) , .B2( u0_u3_n787 ) );
  NOR2_X1 u0_u3_U376 (.A1( u0_u3_n672 ) , .ZN( u0_u3_n769 ) , .A2( u0_u3_n816 ) );
  NOR2_X1 u0_u3_U377 (.A2( u0_u3_n816 ) , .A1( u0_u3_n818 ) , .ZN( u0_u3_n824 ) );
  NOR2_X1 u0_u3_U378 (.ZN( u0_u3_n581 ) , .A1( u0_u3_n711 ) , .A2( u0_u3_n816 ) );
  NOR2_X1 u0_u3_U379 (.A1( u0_u3_n439 ) , .ZN( u0_u3_n687 ) , .A2( u0_u3_n816 ) );
  NOR3_X1 u0_u3_U38 (.A3( u0_u3_n651 ) , .A2( u0_u3_n652 ) , .A1( u0_u3_n653 ) , .ZN( u0_u3_n662 ) );
  NOR2_X1 u0_u3_U380 (.ZN( u0_u3_n657 ) , .A1( u0_u3_n731 ) , .A2( u0_u3_n816 ) );
  NOR2_X1 u0_u3_U381 (.A1( u0_u3_n702 ) , .ZN( u0_u3_n771 ) , .A2( u0_u3_n816 ) );
  NOR2_X1 u0_u3_U382 (.ZN( u0_u3_n668 ) , .A1( u0_u3_n783 ) , .A2( u0_u3_n816 ) );
  NOR2_X1 u0_u3_U383 (.ZN( u0_u3_n634 ) , .A1( u0_u3_n727 ) , .A2( u0_u3_n816 ) );
  NOR2_X1 u0_u3_U384 (.ZN( u0_u3_n475 ) , .A2( w3_26 ) , .A1( w3_27 ) );
  NOR2_X1 u0_u3_U385 (.ZN( u0_u3_n458 ) , .A1( u0_u3_n831 ) , .A2( w3_27 ) );
  INV_X1 u0_u3_U386 (.ZN( u0_u3_n832 ) , .A( w3_27 ) );
  NOR3_X1 u0_u3_U387 (.A3( u0_u3_n624 ) , .A2( u0_u3_n625 ) , .ZN( u0_u3_n639 ) , .A1( u0_u3_n728 ) );
  NOR4_X1 u0_u3_U388 (.A1( u0_u3_n587 ) , .ZN( u0_u3_n588 ) , .A3( u0_u3_n655 ) , .A2( u0_u3_n665 ) , .A4( u0_u3_n770 ) );
  OAI22_X1 u0_u3_U389 (.ZN( u0_u3_n640 ) , .A1( u0_u3_n702 ) , .B2( u0_u3_n731 ) , .A2( u0_u3_n765 ) , .B1( u0_u3_n819 ) );
  NOR3_X1 u0_u3_U39 (.A3( u0_u3_n657 ) , .A2( u0_u3_n658 ) , .A1( u0_u3_n659 ) , .ZN( u0_u3_n660 ) );
  AOI21_X1 u0_u3_U390 (.ZN( u0_u3_n502 ) , .B1( u0_u3_n683 ) , .A( u0_u3_n815 ) , .B2( u0_u3_n819 ) );
  OAI22_X1 u0_u3_U391 (.A1( u0_u3_n727 ) , .ZN( u0_u3_n729 ) , .B2( u0_u3_n753 ) , .B1( u0_u3_n815 ) , .A2( u0_u3_n819 ) );
  AOI21_X1 u0_u3_U392 (.A( u0_u3_n438 ) , .B2( u0_u3_n819 ) , .B1( u0_u3_n820 ) , .ZN( u0_u3_n821 ) );
  OAI22_X1 u0_u3_U393 (.A1( u0_u3_n438 ) , .ZN( u0_u3_n627 ) , .B1( u0_u3_n672 ) , .B2( u0_u3_n750 ) , .A2( u0_u3_n819 ) );
  NOR2_X1 u0_u3_U394 (.ZN( u0_u3_n522 ) , .A2( u0_u3_n702 ) , .A1( u0_u3_n819 ) );
  NOR2_X1 u0_u3_U395 (.A1( u0_u3_n672 ) , .ZN( u0_u3_n691 ) , .A2( u0_u3_n819 ) );
  NOR2_X1 u0_u3_U396 (.A2( u0_u3_n439 ) , .ZN( u0_u3_n602 ) , .A1( u0_u3_n819 ) );
  NOR2_X1 u0_u3_U397 (.ZN( u0_u3_n534 ) , .A2( u0_u3_n783 ) , .A1( u0_u3_n819 ) );
  NOR2_X1 u0_u3_U398 (.ZN( u0_u3_n561 ) , .A1( u0_u3_n711 ) , .A2( u0_u3_n819 ) );
  NOR2_X1 u0_u3_U399 (.ZN( u0_u3_n688 ) , .A1( u0_u3_n732 ) , .A2( u0_u3_n819 ) );
  NAND2_X1 u0_u3_U4 (.A1( u0_u3_n452 ) , .A2( u0_u3_n463 ) , .ZN( u0_u3_n795 ) );
  NOR4_X1 u0_u3_U40 (.A4( u0_u3_n664 ) , .A3( u0_u3_n665 ) , .A2( u0_u3_n666 ) , .A1( u0_u3_n667 ) , .ZN( u0_u3_n680 ) );
  INV_X1 u0_u3_U400 (.A( u0_u3_n819 ) , .ZN( u0_u3_n834 ) );
  NAND2_X1 u0_u3_U401 (.ZN( u0_u3_n674 ) , .A1( u0_u3_n809 ) , .A2( u0_u3_n819 ) );
  NOR2_X1 u0_u3_U402 (.ZN( u0_u3_n465 ) , .A2( w3_24 ) , .A1( w3_25 ) );
  NOR2_X1 u0_u3_U403 (.ZN( u0_u3_n457 ) , .A1( u0_u3_n830 ) , .A2( w3_24 ) );
  INV_X1 u0_u3_U404 (.ZN( u0_u3_n829 ) , .A( w3_24 ) );
  INV_X1 u0_u3_U405 (.ZN( u0_u3_n850 ) , .A( w3_29 ) );
  NOR2_X1 u0_u3_U406 (.ZN( u0_u3_n451 ) , .A1( u0_u3_n849 ) , .A2( w3_29 ) );
  NAND4_X1 u0_u3_U407 (.ZN( u0_subword_3 ) , .A4( u0_u3_n707 ) , .A3( u0_u3_n708 ) , .A2( u0_u3_n709 ) , .A1( u0_u3_n710 ) );
  INV_X1 u0_u3_U408 (.A( u0_u3_n709 ) , .ZN( u0_u3_n878 ) );
  OAI22_X1 u0_u3_U409 (.B2( u0_u3_n747 ) , .ZN( u0_u3_n749 ) , .A2( u0_u3_n765 ) , .B1( u0_u3_n783 ) , .A1( u0_u3_n795 ) );
  NOR4_X1 u0_u3_U41 (.A4( u0_u3_n668 ) , .A3( u0_u3_n669 ) , .A2( u0_u3_n670 ) , .A1( u0_u3_n671 ) , .ZN( u0_u3_n679 ) );
  OAI22_X1 u0_u3_U410 (.B1( u0_u3_n439 ) , .ZN( u0_u3_n499 ) , .A2( u0_u3_n747 ) , .A1( u0_u3_n783 ) , .B2( u0_u3_n809 ) );
  NOR2_X1 u0_u3_U411 (.ZN( u0_u3_n519 ) , .A1( u0_u3_n711 ) , .A2( u0_u3_n747 ) );
  OAI22_X1 u0_u3_U412 (.ZN( u0_u3_n713 ) , .A2( u0_u3_n731 ) , .B2( u0_u3_n732 ) , .A1( u0_u3_n747 ) , .B1( u0_u3_n816 ) );
  NOR2_X1 u0_u3_U413 (.A2( u0_u3_n747 ) , .ZN( u0_u3_n772 ) , .A1( u0_u3_n815 ) );
  OAI22_X1 u0_u3_U414 (.B1( u0_u3_n443 ) , .ZN( u0_u3_n447 ) , .A2( u0_u3_n731 ) , .A1( u0_u3_n747 ) , .B2( u0_u3_n752 ) );
  NOR2_X1 u0_u3_U415 (.ZN( u0_u3_n550 ) , .A1( u0_u3_n702 ) , .A2( u0_u3_n747 ) );
  NOR2_X1 u0_u3_U416 (.ZN( u0_u3_n556 ) , .A2( u0_u3_n747 ) , .A1( u0_u3_n787 ) );
  NOR2_X1 u0_u3_U417 (.A2( u0_u3_n747 ) , .ZN( u0_u3_n758 ) , .A1( u0_u3_n808 ) );
  NOR2_X1 u0_u3_U418 (.A1( u0_u3_n672 ) , .ZN( u0_u3_n676 ) , .A2( u0_u3_n747 ) );
  NOR2_X1 u0_u3_U419 (.ZN( u0_u3_n533 ) , .A2( u0_u3_n747 ) , .A1( u0_u3_n795 ) );
  NOR4_X1 u0_u3_U42 (.A3( u0_u3_n676 ) , .A1( u0_u3_n677 ) , .ZN( u0_u3_n678 ) , .A4( u0_u3_n718 ) , .A2( u0_u3_n861 ) );
  NOR2_X1 u0_u3_U420 (.ZN( u0_u3_n721 ) , .A2( u0_u3_n727 ) , .A1( u0_u3_n747 ) );
  NOR2_X1 u0_u3_U421 (.ZN( u0_u3_n585 ) , .A1( u0_u3_n747 ) , .A2( u0_u3_n818 ) );
  INV_X1 u0_u3_U422 (.A( u0_u3_n747 ) , .ZN( u0_u3_n839 ) );
  AOI21_X1 u0_u3_U423 (.ZN( u0_u3_n579 ) , .B2( u0_u3_n727 ) , .B1( u0_u3_n751 ) , .A( u0_u3_n788 ) );
  NAND4_X1 u0_u3_U424 (.A4( u0_u3_n636 ) , .A3( u0_u3_n637 ) , .A2( u0_u3_n638 ) , .A1( u0_u3_n639 ) , .ZN( u0_u3_n746 ) );
  INV_X1 u0_u3_U425 (.ZN( u0_u3_n851 ) , .A( w3_30 ) );
  INV_X1 u0_u3_U426 (.ZN( u0_u3_n860 ) , .A( w3_31 ) );
  NAND4_X1 u0_u3_U427 (.ZN( u0_subword_2 ) , .A4( u0_u3_n646 ) , .A3( u0_u3_n647 ) , .A2( u0_u3_n648 ) , .A1( u0_u3_n649 ) );
  AOI211_X1 u0_u3_U428 (.A( u0_u3_n640 ) , .ZN( u0_u3_n648 ) , .B( u0_u3_n746 ) , .C2( u0_u3_n841 ) , .C1( u0_u3_n856 ) );
  NOR2_X1 u0_u3_U429 (.A2( u0_u3_n41 ) , .ZN( u0_u3_n603 ) , .A1( u0_u3_n787 ) );
  NOR4_X1 u0_u3_U43 (.A1( u0_u3_n469 ) , .ZN( u0_u3_n470 ) , .A4( u0_u3_n545 ) , .A2( u0_u3_n557 ) , .A3( u0_u3_n617 ) );
  OAI222_X1 u0_u3_U430 (.A2( u0_u3_n672 ) , .ZN( u0_u3_n677 ) , .B1( u0_u3_n750 ) , .B2( u0_u3_n787 ) , .C2( u0_u3_n791 ) , .C1( u0_u3_n818 ) , .A1( u0_u3_n820 ) );
  NOR2_X1 u0_u3_U431 (.ZN( u0_u3_n613 ) , .A1( u0_u3_n787 ) , .A2( u0_u3_n819 ) );
  AOI21_X1 u0_u3_U432 (.A( u0_u3_n41 ) , .ZN( u0_u3_n503 ) , .B1( u0_u3_n711 ) , .B2( u0_u3_n789 ) );
  OAI22_X1 u0_u3_U433 (.ZN( u0_u3_n593 ) , .B1( u0_u3_n733 ) , .B2( u0_u3_n752 ) , .A2( u0_u3_n789 ) , .A1( u0_u3_n806 ) );
  NOR2_X1 u0_u3_U434 (.ZN( u0_u3_n656 ) , .A1( u0_u3_n765 ) , .A2( u0_u3_n789 ) );
  NAND2_X1 u0_u3_U435 (.A2( u0_u3_n752 ) , .A1( u0_u3_n789 ) , .ZN( u0_u3_n812 ) );
  NOR2_X1 u0_u3_U436 (.ZN( u0_u3_n557 ) , .A1( u0_u3_n789 ) , .A2( u0_u3_n816 ) );
  NAND3_X1 u0_u3_U437 (.ZN( u0_subword_6 ) , .A3( u0_u3_n800 ) , .A2( u0_u3_n801 ) , .A1( u0_u3_n802 ) );
  NAND3_X1 u0_u3_U438 (.ZN( u0_subword_5 ) , .A3( u0_u3_n761 ) , .A2( u0_u3_n762 ) , .A1( u0_u3_n763 ) );
  NAND3_X1 u0_u3_U439 (.ZN( u0_subword_4 ) , .A3( u0_u3_n741 ) , .A2( u0_u3_n742 ) , .A1( u0_u3_n743 ) );
  AOI221_X1 u0_u3_U44 (.ZN( u0_u3_n471 ) , .C2( u0_u3_n717 ) , .B2( u0_u3_n834 ) , .C1( u0_u3_n847 ) , .B1( u0_u3_n862 ) , .A( u0_u3_n866 ) );
  NAND3_X1 u0_u3_U440 (.A3( u0_u3_n678 ) , .A2( u0_u3_n679 ) , .A1( u0_u3_n680 ) , .ZN( u0_u3_n810 ) );
  NAND3_X1 u0_u3_U441 (.ZN( u0_u3_n641 ) , .A3( u0_u3_n711 ) , .A2( u0_u3_n727 ) , .A1( u0_u3_n795 ) );
  NAND3_X1 u0_u3_U442 (.A3( u0_u3_n621 ) , .A2( u0_u3_n622 ) , .A1( u0_u3_n623 ) , .ZN( u0_u3_n728 ) );
  NAND3_X1 u0_u3_U443 (.A3( u0_u3_n588 ) , .A2( u0_u3_n589 ) , .A1( u0_u3_n590 ) , .ZN( u0_u3_n624 ) );
  NAND3_X1 u0_u3_U444 (.ZN( u0_u3_n568 ) , .A3( u0_u3_n683 ) , .A2( u0_u3_n753 ) , .A1( u0_u3_n788 ) );
  NAND3_X1 u0_u3_U445 (.A3( u0_u3_n526 ) , .A2( u0_u3_n527 ) , .A1( u0_u3_n528 ) , .ZN( u0_u3_n745 ) );
  NAND3_X1 u0_u3_U446 (.A3( u0_u3_n515 ) , .A1( u0_u3_n516 ) , .ZN( u0_u3_n611 ) , .A2( u0_u3_n873 ) );
  NAND3_X1 u0_u3_U447 (.A3( u0_u3_n470 ) , .A2( u0_u3_n471 ) , .A1( u0_u3_n472 ) , .ZN( u0_u3_n780 ) );
  NOR2_X1 u0_u3_U448 (.ZN( u0_u3_n615 ) , .A1( u0_u3_n782 ) , .A2( u0_u3_n789 ) );
  NOR2_X1 u0_u3_U449 (.ZN( u0_u3_n720 ) , .A2( u0_u3_n747 ) , .A1( u0_u3_n789 ) );
  NOR4_X1 u0_u3_U45 (.A4( u0_u3_n517 ) , .A3( u0_u3_n518 ) , .A2( u0_u3_n519 ) , .A1( u0_u3_n520 ) , .ZN( u0_u3_n527 ) );
  NOR2_X1 u0_u3_U450 (.ZN( u0_u3_n704 ) , .A2( u0_u3_n789 ) , .A1( u0_u3_n820 ) );
  NOR2_X1 u0_u3_U451 (.A1( u0_u3_n733 ) , .ZN( u0_u3_n768 ) , .A2( u0_u3_n789 ) );
  INV_X1 u0_u3_U452 (.ZN( u0_u3_n849 ) , .A( w3_28 ) );
  NOR4_X1 u0_u3_U46 (.A3( u0_u3_n524 ) , .A1( u0_u3_n525 ) , .ZN( u0_u3_n526 ) , .A2( u0_u3_n676 ) , .A4( u0_u3_n772 ) );
  NAND4_X1 u0_u3_U47 (.A4( u0_u3_n576 ) , .A3( u0_u3_n577 ) , .A1( u0_u3_n578 ) , .ZN( u0_u3_n726 ) , .A2( u0_u3_n876 ) );
  NOR4_X1 u0_u3_U48 (.A4( u0_u3_n572 ) , .A3( u0_u3_n573 ) , .A2( u0_u3_n574 ) , .A1( u0_u3_n575 ) , .ZN( u0_u3_n576 ) );
  INV_X1 u0_u3_U49 (.A( u0_u3_n610 ) , .ZN( u0_u3_n876 ) );
  NAND2_X1 u0_u3_U5 (.A1( u0_u3_n456 ) , .A2( u0_u3_n475 ) , .ZN( u0_u3_n788 ) );
  NAND4_X1 u0_u3_U50 (.A4( u0_u3_n459 ) , .A3( u0_u3_n460 ) , .A2( u0_u3_n461 ) , .A1( u0_u3_n462 ) , .ZN( u0_u3_n682 ) );
  NOR3_X1 u0_u3_U51 (.ZN( u0_u3_n460 ) , .A3( u0_u3_n533 ) , .A1( u0_u3_n558 ) , .A2( u0_u3_n573 ) );
  NOR4_X1 u0_u3_U52 (.ZN( u0_u3_n459 ) , .A2( u0_u3_n520 ) , .A1( u0_u3_n546 ) , .A3( u0_u3_n582 ) , .A4( u0_u3_n618 ) );
  NOR4_X1 u0_u3_U53 (.ZN( u0_u3_n461 ) , .A2( u0_u3_n512 ) , .A1( u0_u3_n602 ) , .A4( u0_u3_n631 ) , .A3( u0_u3_n714 ) );
  NAND4_X1 u0_u3_U54 (.A4( u0_u3_n722 ) , .A3( u0_u3_n723 ) , .A2( u0_u3_n724 ) , .ZN( u0_u3_n744 ) , .A1( u0_u3_n859 ) );
  INV_X1 u0_u3_U55 (.A( u0_u3_n712 ) , .ZN( u0_u3_n859 ) );
  NOR4_X1 u0_u3_U56 (.A4( u0_u3_n718 ) , .A3( u0_u3_n719 ) , .A2( u0_u3_n720 ) , .A1( u0_u3_n721 ) , .ZN( u0_u3_n722 ) );
  NOR3_X1 u0_u3_U57 (.ZN( u0_u3_n483 ) , .A2( u0_u3_n511 ) , .A3( u0_u3_n604 ) , .A1( u0_u3_n613 ) );
  NOR4_X1 u0_u3_U58 (.ZN( u0_u3_n484 ) , .A3( u0_u3_n535 ) , .A4( u0_u3_n548 ) , .A2( u0_u3_n570 ) , .A1( u0_u3_n720 ) );
  AOI211_X1 u0_u3_U59 (.B( u0_u3_n480 ) , .A( u0_u3_n481 ) , .ZN( u0_u3_n485 ) , .C2( u0_u3_n836 ) , .C1( u0_u3_n863 ) );
  NOR3_X1 u0_u3_U6 (.ZN( u0_u3_n601 ) , .A1( u0_u3_n611 ) , .A3( u0_u3_n726 ) , .A2( u0_u3_n745 ) );
  INV_X1 u0_u3_U60 (.A( u0_u3_n682 ) , .ZN( u0_u3_n874 ) );
  NOR4_X1 u0_u3_U61 (.A4( u0_u3_n690 ) , .A3( u0_u3_n691 ) , .A2( u0_u3_n692 ) , .A1( u0_u3_n693 ) , .ZN( u0_u3_n694 ) );
  AOI221_X1 u0_u3_U62 (.A( u0_u3_n684 ) , .ZN( u0_u3_n695 ) , .B2( u0_u3_n842 ) , .C1( u0_u3_n844 ) , .C2( u0_u3_n864 ) , .B1( u0_u3_n867 ) );
  NAND4_X1 u0_u3_U63 (.A4( u0_u3_n476 ) , .A3( u0_u3_n477 ) , .A2( u0_u3_n478 ) , .A1( u0_u3_n479 ) , .ZN( u0_u3_n681 ) );
  NOR4_X1 u0_u3_U64 (.A4( u0_u3_n473 ) , .ZN( u0_u3_n479 ) , .A3( u0_u3_n559 ) , .A1( u0_u3_n738 ) , .A2( u0_u3_n758 ) );
  NOR4_X1 u0_u3_U65 (.ZN( u0_u3_n477 ) , .A1( u0_u3_n509 ) , .A3( u0_u3_n547 ) , .A2( u0_u3_n586 ) , .A4( u0_u3_n719 ) );
  NOR4_X1 u0_u3_U66 (.ZN( u0_u3_n476 ) , .A2( u0_u3_n524 ) , .A4( u0_u3_n597 ) , .A1( u0_u3_n612 ) , .A3( u0_u3_n632 ) );
  NAND4_X1 u0_u3_U67 (.A4( u0_u3_n551 ) , .A3( u0_u3_n552 ) , .A2( u0_u3_n553 ) , .A1( u0_u3_n554 ) , .ZN( u0_u3_n748 ) );
  AOI211_X1 u0_u3_U68 (.B( u0_u3_n542 ) , .A( u0_u3_n543 ) , .ZN( u0_u3_n554 ) , .C2( u0_u3_n841 ) , .C1( u0_u3_n853 ) );
  NOR3_X1 u0_u3_U69 (.ZN( u0_u3_n552 ) , .A2( u0_u3_n654 ) , .A1( u0_u3_n670 ) , .A3( u0_u3_n774 ) );
  NOR3_X1 u0_u3_U7 (.ZN( u0_u3_n507 ) , .A2( u0_u3_n682 ) , .A3( u0_u3_n780 ) , .A1( u0_u3_n878 ) );
  NOR4_X1 u0_u3_U70 (.A4( u0_u3_n544 ) , .A3( u0_u3_n545 ) , .A2( u0_u3_n546 ) , .ZN( u0_u3_n553 ) , .A1( u0_u3_n691 ) );
  NOR4_X1 u0_u3_U71 (.A4( u0_u3_n612 ) , .A3( u0_u3_n613 ) , .A2( u0_u3_n614 ) , .A1( u0_u3_n615 ) , .ZN( u0_u3_n622 ) );
  NOR4_X1 u0_u3_U72 (.ZN( u0_u3_n623 ) , .A1( u0_u3_n659 ) , .A3( u0_u3_n669 ) , .A4( u0_u3_n685 ) , .A2( u0_u3_n769 ) );
  INV_X1 u0_u3_U73 (.A( u0_u3_n765 ) , .ZN( u0_u3_n833 ) );
  NOR2_X1 u0_u3_U74 (.ZN( u0_u3_n650 ) , .A1( u0_u3_n856 ) , .A2( u0_u3_n870 ) );
  NOR4_X1 u0_u3_U75 (.A4( u0_u3_n580 ) , .A3( u0_u3_n581 ) , .A2( u0_u3_n582 ) , .ZN( u0_u3_n589 ) , .A1( u0_u3_n686 ) );
  INV_X1 u0_u3_U76 (.A( u0_u3_n818 ) , .ZN( u0_u3_n857 ) );
  OR4_X1 u0_u3_U77 (.A4( u0_u3_n685 ) , .A3( u0_u3_n686 ) , .A2( u0_u3_n687 ) , .A1( u0_u3_n688 ) , .ZN( u0_u3_n693 ) );
  OR4_X1 u0_u3_U78 (.ZN( u0_u3_n469 ) , .A4( u0_u3_n521 ) , .A3( u0_u3_n532 ) , .A2( u0_u3_n581 ) , .A1( u0_u3_n715 ) );
  OR4_X1 u0_u3_U79 (.A4( u0_u3_n569 ) , .A3( u0_u3_n570 ) , .A2( u0_u3_n571 ) , .ZN( u0_u3_n575 ) , .A1( u0_u3_n668 ) );
  NOR3_X1 u0_u3_U8 (.A2( u0_u3_n610 ) , .A1( u0_u3_n611 ) , .ZN( u0_u3_n649 ) , .A3( u0_u3_n725 ) );
  OR4_X1 u0_u3_U80 (.A4( u0_u3_n521 ) , .A2( u0_u3_n522 ) , .A1( u0_u3_n523 ) , .ZN( u0_u3_n525 ) , .A3( u0_u3_n824 ) );
  OR4_X1 u0_u3_U81 (.A4( u0_u3_n583 ) , .A3( u0_u3_n584 ) , .A2( u0_u3_n585 ) , .A1( u0_u3_n586 ) , .ZN( u0_u3_n587 ) );
  OR4_X1 u0_u3_U82 (.ZN( u0_u3_n495 ) , .A4( u0_u3_n537 ) , .A2( u0_u3_n550 ) , .A1( u0_u3_n562 ) , .A3( u0_u3_n635 ) );
  NOR4_X1 u0_u3_U83 (.A4( u0_u3_n512 ) , .A2( u0_u3_n513 ) , .A1( u0_u3_n514 ) , .ZN( u0_u3_n515 ) , .A3( u0_u3_n673 ) );
  INV_X1 u0_u3_U84 (.A( u0_u3_n508 ) , .ZN( u0_u3_n873 ) );
  OR3_X1 u0_u3_U85 (.A3( u0_u3_n509 ) , .A2( u0_u3_n510 ) , .A1( u0_u3_n511 ) , .ZN( u0_u3_n514 ) );
  INV_X1 u0_u3_U86 (.A( u0_u3_n757 ) , .ZN( u0_u3_n871 ) );
  AOI221_X1 u0_u3_U87 (.A( u0_u3_n716 ) , .B2( u0_u3_n717 ) , .ZN( u0_u3_n723 ) , .C1( u0_u3_n835 ) , .B1( u0_u3_n841 ) , .C2( u0_u3_n865 ) );
  OR2_X1 u0_u3_U88 (.A2( u0_u3_n714 ) , .A1( u0_u3_n715 ) , .ZN( u0_u3_n716 ) );
  INV_X1 u0_u3_U89 (.A( u0_u3_n466 ) , .ZN( u0_u3_n866 ) );
  NOR3_X1 u0_u3_U9 (.A3( u0_u3_n725 ) , .A1( u0_u3_n726 ) , .ZN( u0_u3_n743 ) , .A2( u0_u3_n744 ) );
  NAND2_X1 u0_u3_U90 (.A1( u0_u3_n454 ) , .A2( u0_u3_n456 ) , .ZN( u0_u3_n765 ) );
  AOI22_X1 u0_u3_U91 (.ZN( u0_u3_n699 ) , .A1( u0_u3_n833 ) , .B2( u0_u3_n845 ) , .A2( u0_u3_n867 ) , .B1( u0_u3_n870 ) );
  NOR3_X1 u0_u3_U92 (.ZN( u0_u3_n755 ) , .A2( u0_u3_n855 ) , .A1( u0_u3_n865 ) , .A3( u0_u3_n867 ) );
  NOR2_X1 u0_u3_U93 (.ZN( u0_u3_n754 ) , .A2( u0_u3_n854 ) , .A1( u0_u3_n862 ) );
  AOI211_X1 u0_u3_U94 (.A( u0_u3_n499 ) , .ZN( u0_u3_n506 ) , .B( u0_u3_n805 ) , .C2( u0_u3_n841 ) , .C1( u0_u3_n853 ) );
  AOI211_X1 u0_u3_U95 (.B( u0_u3_n810 ) , .A( u0_u3_n811 ) , .ZN( u0_u3_n827 ) , .C1( u0_u3_n844 ) , .C2( u0_u3_n852 ) );
  NAND2_X1 u0_u3_U96 (.A1( u0_u3_n450 ) , .A2( u0_u3_n468 ) , .ZN( u0_u3_n752 ) );
  INV_X1 u0_u3_U97 (.A( u0_u3_n733 ) , .ZN( u0_u3_n841 ) );
  AOI221_X1 u0_u3_U98 (.B2( u0_u3_n440 ) , .A( u0_u3_n492 ) , .ZN( u0_u3_n497 ) , .C2( u0_u3_n843 ) , .C1( u0_u3_n853 ) , .B1( u0_u3_n862 ) );
  INV_X1 u0_u3_U99 (.A( u0_u3_n781 ) , .ZN( u0_u3_n869 ) );
endmodule

