module aes_aes_die_14 ( sa31_0, sa31_1, sa31_2, sa31_3, sa31_4, sa31_5, sa31_6, sa31_7, sa32_sr_0, sa32_sr_1, sa32_sr_2, sa32_sr_3, sa32_sr_4, sa32_sr_5, sa32_sr_6, sa32_sr_7 );
  input sa31_0, sa31_1, sa31_2, sa31_3, sa31_4, sa31_5, sa31_6, sa31_7;
  output sa32_sr_0, sa32_sr_1, sa32_sr_2, sa32_sr_3, sa32_sr_4, sa32_sr_5, sa32_sr_6, sa32_sr_7;
  wire us31_n438, us31_n439, us31_n440, us31_n441, us31_n442, us31_n443, us31_n444, us31_n445, us31_n446, 
       us31_n447, us31_n448, us31_n449, us31_n450, us31_n451, us31_n452, us31_n453, us31_n454, us31_n455, 
       us31_n456, us31_n457, us31_n458, us31_n459, us31_n460, us31_n461, us31_n462, us31_n463, us31_n464, 
       us31_n465, us31_n466, us31_n467, us31_n468, us31_n469, us31_n470, us31_n471, us31_n472, us31_n473, 
       us31_n474, us31_n475, us31_n476, us31_n477, us31_n478, us31_n479, us31_n480, us31_n481, us31_n482, 
       us31_n483, us31_n484, us31_n485, us31_n486, us31_n487, us31_n488, us31_n489, us31_n490, us31_n491, 
       us31_n492, us31_n493, us31_n494, us31_n495, us31_n496, us31_n497, us31_n498, us31_n499, us31_n500, 
       us31_n501, us31_n502, us31_n503, us31_n504, us31_n505, us31_n506, us31_n507, us31_n508, us31_n509, 
       us31_n510, us31_n511, us31_n512, us31_n513, us31_n514, us31_n515, us31_n516, us31_n517, us31_n518, 
       us31_n519, us31_n520, us31_n521, us31_n522, us31_n523, us31_n524, us31_n525, us31_n526, us31_n527, 
       us31_n528, us31_n529, us31_n530, us31_n531, us31_n532, us31_n533, us31_n534, us31_n535, us31_n536, 
       us31_n537, us31_n538, us31_n539, us31_n540, us31_n541, us31_n542, us31_n543, us31_n544, us31_n545, 
       us31_n546, us31_n547, us31_n548, us31_n549, us31_n550, us31_n551, us31_n552, us31_n553, us31_n554, 
       us31_n555, us31_n556, us31_n557, us31_n558, us31_n559, us31_n560, us31_n561, us31_n562, us31_n563, 
       us31_n564, us31_n565, us31_n566, us31_n567, us31_n568, us31_n569, us31_n570, us31_n571, us31_n572, 
       us31_n573, us31_n574, us31_n575, us31_n576, us31_n577, us31_n578, us31_n579, us31_n580, us31_n581, 
       us31_n582, us31_n583, us31_n584, us31_n585, us31_n586, us31_n587, us31_n588, us31_n589, us31_n590, 
       us31_n591, us31_n592, us31_n593, us31_n594, us31_n595, us31_n596, us31_n597, us31_n598, us31_n599, 
       us31_n600, us31_n601, us31_n602, us31_n603, us31_n604, us31_n605, us31_n606, us31_n607, us31_n608, 
       us31_n609, us31_n610, us31_n611, us31_n612, us31_n613, us31_n614, us31_n615, us31_n616, us31_n617, 
       us31_n618, us31_n619, us31_n620, us31_n621, us31_n622, us31_n623, us31_n624, us31_n625, us31_n626, 
       us31_n627, us31_n628, us31_n629, us31_n630, us31_n631, us31_n632, us31_n633, us31_n634, us31_n635, 
       us31_n636, us31_n637, us31_n638, us31_n639, us31_n640, us31_n641, us31_n642, us31_n643, us31_n644, 
       us31_n645, us31_n646, us31_n647, us31_n648, us31_n649, us31_n650, us31_n651, us31_n652, us31_n653, 
       us31_n654, us31_n655, us31_n656, us31_n657, us31_n658, us31_n659, us31_n660, us31_n661, us31_n662, 
       us31_n663, us31_n664, us31_n665, us31_n666, us31_n667, us31_n668, us31_n669, us31_n670, us31_n671, 
       us31_n672, us31_n673, us31_n674, us31_n675, us31_n676, us31_n677, us31_n678, us31_n679, us31_n680, 
       us31_n681, us31_n682, us31_n683, us31_n684, us31_n685, us31_n686, us31_n687, us31_n688, us31_n689, 
       us31_n690, us31_n691, us31_n692, us31_n693, us31_n694, us31_n695, us31_n696, us31_n697, us31_n698, 
       us31_n699, us31_n700, us31_n701, us31_n702, us31_n703, us31_n704, us31_n705, us31_n706, us31_n707, 
       us31_n708, us31_n709, us31_n710, us31_n711, us31_n712, us31_n713, us31_n714, us31_n715, us31_n716, 
       us31_n717, us31_n718, us31_n719, us31_n720, us31_n721, us31_n722, us31_n723, us31_n724, us31_n725, 
       us31_n726, us31_n727, us31_n728, us31_n729, us31_n730, us31_n731, us31_n732, us31_n733, us31_n734, 
       us31_n735, us31_n736, us31_n737, us31_n738, us31_n739, us31_n740, us31_n741, us31_n742, us31_n743, 
       us31_n744, us31_n745, us31_n746, us31_n747, us31_n748, us31_n749, us31_n750, us31_n751, us31_n752, 
       us31_n753, us31_n754, us31_n755, us31_n756, us31_n757, us31_n758, us31_n759, us31_n760, us31_n761, 
       us31_n762, us31_n763, us31_n764, us31_n765, us31_n766, us31_n767, us31_n768, us31_n769, us31_n770, 
       us31_n771, us31_n772, us31_n773, us31_n774, us31_n775, us31_n776, us31_n777, us31_n778, us31_n779, 
       us31_n780, us31_n781, us31_n782, us31_n783, us31_n784, us31_n785, us31_n786, us31_n787, us31_n788, 
       us31_n789, us31_n790, us31_n791, us31_n792, us31_n793, us31_n794, us31_n795, us31_n796, us31_n797, 
       us31_n798, us31_n799, us31_n800, us31_n801, us31_n802, us31_n803, us31_n804, us31_n805, us31_n806, 
       us31_n807, us31_n808, us31_n809, us31_n810, us31_n811, us31_n812, us31_n813, us31_n814, us31_n815, 
       us31_n816, us31_n817, us31_n818, us31_n819, us31_n820, us31_n821, us31_n822, us31_n823, us31_n824, 
       us31_n825, us31_n826, us31_n827, us31_n828, us31_n829, us31_n830, us31_n831, us31_n832, us31_n833, 
       us31_n834, us31_n835, us31_n836, us31_n837, us31_n838, us31_n839, us31_n840, us31_n841, us31_n842, 
       us31_n843, us31_n844, us31_n845, us31_n846, us31_n847, us31_n848, us31_n849, us31_n850, us31_n851, 
       us31_n852, us31_n853, us31_n854, us31_n855, us31_n856, us31_n857, us31_n858, us31_n859, us31_n860, 
       us31_n861, us31_n862, us31_n863, us31_n864, us31_n865, us31_n866, us31_n867, us31_n868, us31_n869, 
       us31_n870, us31_n871, us31_n872, us31_n873, us31_n874, us31_n875,  us31_n876;
  NOR3_X1 us31_U10 (.A3( us31_n621 ) , .A2( us31_n622 ) , .ZN( us31_n636 ) , .A1( us31_n725 ) );
  NOR4_X1 us31_U100 (.ZN( us31_n458 ) , .A2( us31_n509 ) , .A1( us31_n599 ) , .A4( us31_n628 ) , .A3( us31_n711 ) );
  NAND4_X1 us31_U101 (.A4( us31_n535 ) , .A3( us31_n536 ) , .A2( us31_n537 ) , .A1( us31_n538 ) , .ZN( us31_n622 ) );
  NOR4_X1 us31_U102 (.A4( us31_n526 ) , .A2( us31_n527 ) , .A1( us31_n528 ) , .ZN( us31_n538 ) , .A3( us31_n701 ) );
  NOR4_X1 us31_U103 (.A1( us31_n531 ) , .ZN( us31_n536 ) , .A2( us31_n654 ) , .A4( us31_n668 ) , .A3( us31_n765 ) );
  NOR4_X1 us31_U104 (.A4( us31_n529 ) , .A3( us31_n530 ) , .ZN( us31_n537 ) , .A2( us31_n684 ) , .A1( us31_n794 ) );
  NOR2_X1 us31_U105 (.ZN( us31_n647 ) , .A1( us31_n854 ) , .A2( us31_n868 ) );
  NAND4_X1 us31_U106 (.A4( us31_n548 ) , .A3( us31_n549 ) , .A2( us31_n550 ) , .A1( us31_n551 ) , .ZN( us31_n745 ) );
  NOR3_X1 us31_U107 (.ZN( us31_n549 ) , .A2( us31_n651 ) , .A1( us31_n667 ) , .A3( us31_n771 ) );
  AOI211_X1 us31_U108 (.B( us31_n539 ) , .A( us31_n540 ) , .ZN( us31_n551 ) , .C2( us31_n839 ) , .C1( us31_n851 ) );
  NOR4_X1 us31_U109 (.A4( us31_n541 ) , .A3( us31_n542 ) , .A2( us31_n543 ) , .ZN( us31_n550 ) , .A1( us31_n688 ) );
  NOR2_X1 us31_U11 (.A1( us31_n678 ) , .ZN( us31_n693 ) , .A2( us31_n807 ) );
  NAND4_X1 us31_U110 (.A4( us31_n479 ) , .A3( us31_n480 ) , .A2( us31_n481 ) , .A1( us31_n482 ) , .ZN( us31_n694 ) );
  NOR3_X1 us31_U111 (.ZN( us31_n480 ) , .A2( us31_n508 ) , .A3( us31_n601 ) , .A1( us31_n610 ) );
  AOI211_X1 us31_U112 (.B( us31_n477 ) , .A( us31_n478 ) , .ZN( us31_n482 ) , .C2( us31_n833 ) , .C1( us31_n861 ) );
  NOR4_X1 us31_U113 (.ZN( us31_n481 ) , .A3( us31_n532 ) , .A4( us31_n545 ) , .A2( us31_n567 ) , .A1( us31_n717 ) );
  NOR2_X1 us31_U114 (.ZN( us31_n686 ) , .A1( us31_n831 ) , .A2( us31_n832 ) );
  NAND4_X1 us31_U115 (.A4( us31_n485 ) , .A3( us31_n486 ) , .A2( us31_n487 ) , .A1( us31_n488 ) , .ZN( us31_n778 ) );
  NOR4_X1 us31_U116 (.A4( us31_n484 ) , .ZN( us31_n487 ) , .A1( us31_n566 ) , .A2( us31_n581 ) , .A3( us31_n602 ) );
  NOR4_X1 us31_U117 (.ZN( us31_n486 ) , .A1( us31_n507 ) , .A2( us31_n519 ) , .A4( us31_n546 ) , .A3( us31_n611 ) );
  NOR4_X1 us31_U118 (.ZN( us31_n485 ) , .A2( us31_n533 ) , .A1( us31_n558 ) , .A3( us31_n631 ) , .A4( us31_n718 ) );
  NAND4_X1 us31_U119 (.A4( us31_n691 ) , .A3( us31_n692 ) , .A1( us31_n693 ) , .ZN( us31_n776 ) , .A2( us31_n872 ) );
  NOR2_X1 us31_U12 (.ZN( us31_n495 ) , .A1( us31_n678 ) , .A2( us31_n694 ) );
  AOI221_X1 us31_U120 (.A( us31_n681 ) , .ZN( us31_n692 ) , .B2( us31_n840 ) , .C1( us31_n842 ) , .C2( us31_n862 ) , .B1( us31_n865 ) );
  INV_X1 us31_U121 (.A( us31_n679 ) , .ZN( us31_n872 ) );
  NOR4_X1 us31_U122 (.A4( us31_n687 ) , .A3( us31_n688 ) , .A2( us31_n689 ) , .A1( us31_n690 ) , .ZN( us31_n691 ) );
  NAND4_X1 us31_U123 (.A4( us31_n719 ) , .A3( us31_n720 ) , .A2( us31_n721 ) , .ZN( us31_n741 ) , .A1( us31_n857 ) );
  INV_X1 us31_U124 (.A( us31_n709 ) , .ZN( us31_n857 ) );
  AOI221_X1 us31_U125 (.A( us31_n710 ) , .ZN( us31_n721 ) , .C2( us31_n844 ) , .B2( us31_n845 ) , .C1( us31_n861 ) , .B1( us31_n862 ) );
  NOR4_X1 us31_U126 (.A4( us31_n715 ) , .A3( us31_n716 ) , .A2( us31_n717 ) , .A1( us31_n718 ) , .ZN( us31_n719 ) );
  NAND4_X1 us31_U127 (.A4( us31_n473 ) , .A3( us31_n474 ) , .A2( us31_n475 ) , .A1( us31_n476 ) , .ZN( us31_n678 ) );
  NOR4_X1 us31_U128 (.ZN( us31_n475 ) , .A1( us31_n531 ) , .A3( us31_n568 ) , .A4( us31_n600 ) , .A2( us31_n642 ) );
  NOR4_X1 us31_U129 (.ZN( us31_n473 ) , .A2( us31_n521 ) , .A4( us31_n594 ) , .A1( us31_n609 ) , .A3( us31_n629 ) );
  NOR3_X1 us31_U13 (.ZN( us31_n504 ) , .A2( us31_n679 ) , .A3( us31_n777 ) , .A1( us31_n876 ) );
  NOR4_X1 us31_U130 (.A4( us31_n470 ) , .ZN( us31_n476 ) , .A3( us31_n556 ) , .A1( us31_n735 ) , .A2( us31_n755 ) );
  NOR2_X1 us31_U131 (.ZN( us31_n733 ) , .A2( us31_n832 ) , .A1( us31_n845 ) );
  NOR2_X1 us31_U132 (.ZN( us31_n789 ) , .A2( us31_n862 ) , .A1( us31_n868 ) );
  NAND4_X1 us31_U133 (.A4( us31_n573 ) , .A3( us31_n574 ) , .A1( us31_n575 ) , .ZN( us31_n723 ) , .A2( us31_n874 ) );
  NOR4_X1 us31_U134 (.A4( us31_n569 ) , .A3( us31_n570 ) , .A2( us31_n571 ) , .A1( us31_n572 ) , .ZN( us31_n573 ) );
  AOI221_X1 us31_U135 (.A( us31_n564 ) , .C2( us31_n565 ) , .ZN( us31_n574 ) , .B2( us31_n845 ) , .B1( us31_n852 ) , .C1( us31_n853 ) );
  NOR2_X1 us31_U136 (.ZN( us31_n575 ) , .A1( us31_n622 ) , .A2( us31_n745 ) );
  NAND4_X1 us31_U137 (.A4( us31_n633 ) , .A3( us31_n634 ) , .A2( us31_n635 ) , .A1( us31_n636 ) , .ZN( us31_n743 ) );
  AOI211_X1 us31_U138 (.B( us31_n623 ) , .A( us31_n624 ) , .ZN( us31_n635 ) , .C2( us31_n836 ) , .C1( us31_n863 ) );
  NOR4_X1 us31_U139 (.A4( us31_n629 ) , .A3( us31_n630 ) , .A2( us31_n631 ) , .A1( us31_n632 ) , .ZN( us31_n633 ) );
  INV_X1 us31_U14 (.A( us31_n706 ) , .ZN( us31_n876 ) );
  NOR4_X1 us31_U140 (.A4( us31_n626 ) , .A3( us31_n627 ) , .A2( us31_n628 ) , .ZN( us31_n634 ) , .A1( us31_n664 ) );
  NAND4_X1 us31_U141 (.A4( us31_n493 ) , .A3( us31_n494 ) , .A1( us31_n495 ) , .ZN( us31_n802 ) , .A2( us31_n867 ) );
  AOI221_X1 us31_U142 (.A( us31_n489 ) , .ZN( us31_n494 ) , .B2( us31_n836 ) , .C2( us31_n841 ) , .C1( us31_n851 ) , .B1( us31_n860 ) );
  INV_X1 us31_U143 (.A( us31_n778 ) , .ZN( us31_n867 ) );
  NOR4_X1 us31_U144 (.A2( us31_n491 ) , .A1( us31_n492 ) , .ZN( us31_n493 ) , .A3( us31_n580 ) , .A4( us31_n612 ) );
  NOR4_X1 us31_U145 (.A4( us31_n734 ) , .A3( us31_n735 ) , .A2( us31_n736 ) , .A1( us31_n737 ) , .ZN( us31_n738 ) );
  AOI211_X1 us31_U146 (.B( us31_n725 ) , .A( us31_n726 ) , .ZN( us31_n739 ) , .C1( us31_n843 ) , .C2( us31_n855 ) );
  NOR3_X1 us31_U147 (.A3( us31_n722 ) , .A1( us31_n723 ) , .ZN( us31_n740 ) , .A2( us31_n741 ) );
  INV_X1 us31_U148 (.A( us31_n762 ) , .ZN( us31_n830 ) );
  INV_X1 us31_U149 (.A( us31_n697 ) , .ZN( us31_n838 ) );
  INV_X1 us31_U15 (.A( us31_n607 ) , .ZN( us31_n874 ) );
  OR4_X1 us31_U150 (.A4( us31_n566 ) , .A3( us31_n567 ) , .A2( us31_n568 ) , .ZN( us31_n572 ) , .A1( us31_n665 ) );
  OR4_X1 us31_U151 (.A4( us31_n682 ) , .A3( us31_n683 ) , .A2( us31_n684 ) , .A1( us31_n685 ) , .ZN( us31_n690 ) );
  OR4_X1 us31_U152 (.ZN( us31_n466 ) , .A4( us31_n518 ) , .A3( us31_n529 ) , .A2( us31_n578 ) , .A1( us31_n712 ) );
  OR4_X1 us31_U153 (.A4( us31_n518 ) , .A2( us31_n519 ) , .A1( us31_n520 ) , .ZN( us31_n522 ) , .A3( us31_n821 ) );
  OR4_X1 us31_U154 (.ZN( us31_n492 ) , .A4( us31_n534 ) , .A2( us31_n547 ) , .A1( us31_n559 ) , .A3( us31_n632 ) );
  OR4_X1 us31_U155 (.A4( us31_n580 ) , .A3( us31_n581 ) , .A2( us31_n582 ) , .A1( us31_n583 ) , .ZN( us31_n584 ) );
  NAND2_X1 us31_U156 (.ZN( us31_n613 ) , .A2( us31_n837 ) , .A1( us31_n873 ) );
  OR3_X1 us31_U157 (.A3( us31_n506 ) , .A2( us31_n507 ) , .A1( us31_n508 ) , .ZN( us31_n511 ) );
  INV_X1 us31_U158 (.A( us31_n463 ) , .ZN( us31_n864 ) );
  OAI21_X1 us31_U159 (.ZN( us31_n463 ) , .B1( us31_n809 ) , .A( us31_n834 ) , .B2( us31_n851 ) );
  INV_X1 us31_U16 (.A( us31_n680 ) , .ZN( us31_n840 ) );
  INV_X1 us31_U160 (.A( us31_n754 ) , .ZN( us31_n869 ) );
  OAI21_X1 us31_U161 (.B1( us31_n753 ) , .ZN( us31_n754 ) , .A( us31_n845 ) , .B2( us31_n868 ) );
  INV_X1 us31_U162 (.A( us31_n672 ) , .ZN( us31_n859 ) );
  AOI21_X1 us31_U163 (.A( us31_n670 ) , .B1( us31_n671 ) , .ZN( us31_n672 ) , .B2( us31_n856 ) );
  OAI222_X1 us31_U164 (.B2( us31_n747 ) , .B1( us31_n748 ) , .A2( us31_n749 ) , .ZN( us31_n757 ) , .C2( us31_n805 ) , .C1( us31_n814 ) , .A1( us31_n817 ) );
  OAI222_X1 us31_U165 (.ZN( us31_n505 ) , .C2( us31_n625 ) , .B2( us31_n647 ) , .B1( us31_n747 ) , .A2( us31_n748 ) , .C1( us31_n805 ) , .A1( us31_n806 ) );
  OAI222_X1 us31_U166 (.B2( us31_n708 ) , .ZN( us31_n709 ) , .C2( us31_n724 ) , .B1( us31_n747 ) , .A1( us31_n806 ) , .C1( us31_n814 ) , .A2( us31_n815 ) );
  NAND2_X1 us31_U167 (.A1( us31_n447 ) , .A2( us31_n465 ) , .ZN( us31_n749 ) );
  AOI22_X1 us31_U168 (.ZN( us31_n696 ) , .A1( us31_n830 ) , .B2( us31_n843 ) , .A2( us31_n865 ) , .B1( us31_n868 ) );
  AOI22_X1 us31_U169 (.A2( us31_n782 ) , .ZN( us31_n783 ) , .B2( us31_n831 ) , .A1( us31_n834 ) , .B1( us31_n863 ) );
  NOR4_X1 us31_U17 (.A4( us31_n445 ) , .A3( us31_n446 ) , .A2( us31_n516 ) , .A1( us31_n541 ) , .ZN( us31_n706 ) );
  INV_X1 us31_U170 (.A( us31_n730 ) , .ZN( us31_n839 ) );
  AOI221_X1 us31_U171 (.A( us31_n764 ) , .ZN( us31_n774 ) , .C2( us31_n810 ) , .B2( us31_n835 ) , .C1( us31_n855 ) , .B1( us31_n866 ) );
  AOI21_X1 us31_U172 (.B2( us31_n763 ) , .ZN( us31_n764 ) , .A( us31_n788 ) , .B1( us31_n792 ) );
  INV_X1 us31_U173 (.A( us31_n761 ) , .ZN( us31_n835 ) );
  AOI221_X1 us31_U174 (.A( us31_n483 ) , .ZN( us31_n488 ) , .B1( us31_n831 ) , .C2( us31_n844 ) , .C1( us31_n852 ) , .B2( us31_n862 ) );
  OAI22_X1 us31_U175 (.ZN( us31_n483 ) , .A1( us31_n708 ) , .B2( us31_n785 ) , .A2( us31_n806 ) , .B1( us31_n812 ) );
  INV_X1 us31_U176 (.A( us31_n790 ) , .ZN( us31_n832 ) );
  NAND2_X1 us31_U177 (.A1( us31_n451 ) , .A2( us31_n453 ) , .ZN( us31_n762 ) );
  AOI211_X1 us31_U178 (.A( us31_n637 ) , .ZN( us31_n645 ) , .B( us31_n743 ) , .C2( us31_n839 ) , .C1( us31_n854 ) );
  OAI22_X1 us31_U179 (.ZN( us31_n637 ) , .A1( us31_n699 ) , .B2( us31_n728 ) , .A2( us31_n762 ) , .B1( us31_n816 ) );
  OR3_X1 us31_U18 (.ZN( us31_n446 ) , .A1( us31_n528 ) , .A3( us31_n577 ) , .A2( us31_n875 ) );
  INV_X1 us31_U180 (.A( us31_n786 ) , .ZN( us31_n862 ) );
  OAI221_X1 us31_U181 (.A( us31_n727 ) , .C2( us31_n728 ) , .B2( us31_n729 ) , .B1( us31_n730 ) , .ZN( us31_n737 ) , .C1( us31_n817 ) );
  AOI22_X1 us31_U182 (.ZN( us31_n727 ) , .B1( us31_n832 ) , .A2( us31_n838 ) , .A1( us31_n863 ) , .B2( us31_n866 ) );
  OAI22_X1 us31_U183 (.ZN( us31_n710 ) , .A2( us31_n728 ) , .B2( us31_n729 ) , .A1( us31_n744 ) , .B1( us31_n813 ) );
  INV_X1 us31_U184 (.A( us31_n816 ) , .ZN( us31_n831 ) );
  OAI22_X1 us31_U185 (.ZN( us31_n624 ) , .B1( us31_n669 ) , .B2( us31_n747 ) , .A1( us31_n815 ) , .A2( us31_n816 ) );
  INV_X1 us31_U186 (.A( us31_n744 ) , .ZN( us31_n837 ) );
  INV_X1 us31_U187 (.A( us31_n788 ) , .ZN( us31_n845 ) );
  OAI22_X1 us31_U188 (.B2( us31_n779 ) , .B1( us31_n780 ) , .ZN( us31_n781 ) , .A2( us31_n814 ) , .A1( us31_n815 ) );
  OAI22_X1 us31_U189 (.A1( us31_n724 ) , .ZN( us31_n726 ) , .B2( us31_n750 ) , .B1( us31_n812 ) , .A2( us31_n816 ) );
  OR4_X1 us31_U19 (.A4( us31_n442 ) , .A2( us31_n443 ) , .A1( us31_n444 ) , .ZN( us31_n445 ) , .A3( us31_n553 ) );
  INV_X1 us31_U190 (.A( us31_n805 ) , .ZN( us31_n860 ) );
  INV_X1 us31_U191 (.A( us31_n814 ) , .ZN( us31_n833 ) );
  INV_X1 us31_U192 (.A( us31_n669 ) , .ZN( us31_n865 ) );
  OAI22_X1 us31_U193 (.B2( us31_n744 ) , .ZN( us31_n746 ) , .A2( us31_n762 ) , .B1( us31_n780 ) , .A1( us31_n792 ) );
  OAI22_X1 us31_U194 (.ZN( us31_n496 ) , .A2( us31_n744 ) , .A1( us31_n780 ) , .B1( us31_n791 ) , .B2( us31_n806 ) );
  OAI22_X1 us31_U195 (.B2( us31_n803 ) , .B1( us31_n804 ) , .A2( us31_n805 ) , .A1( us31_n806 ) , .ZN( us31_n808 ) );
  OAI22_X1 us31_U196 (.ZN( us31_n489 ) , .A1( us31_n724 ) , .B2( us31_n728 ) , .B1( us31_n730 ) , .A2( us31_n779 ) );
  OAI22_X1 us31_U197 (.ZN( us31_n695 ) , .A2( us31_n730 ) , .A1( us31_n780 ) , .B1( us31_n791 ) , .B2( us31_n817 ) );
  OAI22_X1 us31_U198 (.B1( us31_n490 ) , .ZN( us31_n491 ) , .A1( us31_n686 ) , .A2( us31_n763 ) , .B2( us31_n817 ) );
  NOR3_X1 us31_U199 (.ZN( us31_n490 ) , .A1( us31_n782 ) , .A2( us31_n850 ) , .A3( us31_n863 ) );
  INV_X1 us31_U20 (.A( us31_n613 ) , .ZN( us31_n875 ) );
  INV_X1 us31_U200 (.A( us31_n750 ) , .ZN( us31_n842 ) );
  NOR2_X1 us31_U201 (.ZN( us31_n715 ) , .A1( us31_n805 ) , .A2( us31_n817 ) );
  NOR2_X1 us31_U202 (.A2( us31_n744 ) , .ZN( us31_n755 ) , .A1( us31_n805 ) );
  NOR2_X1 us31_U203 (.ZN( us31_n735 ) , .A2( us31_n803 ) , .A1( us31_n805 ) );
  NOR2_X1 us31_U204 (.ZN( us31_n546 ) , .A2( us31_n780 ) , .A1( us31_n814 ) );
  NOR2_X1 us31_U205 (.ZN( us31_n577 ) , .A2( us31_n699 ) , .A1( us31_n814 ) );
  NOR2_X1 us31_U206 (.ZN( us31_n718 ) , .A2( us31_n724 ) , .A1( us31_n744 ) );
  NOR2_X1 us31_U207 (.ZN( us31_n532 ) , .A2( us31_n749 ) , .A1( us31_n750 ) );
  NOR2_X1 us31_U208 (.ZN( us31_n615 ) , .A1( us31_n785 ) , .A2( us31_n815 ) );
  NOR2_X1 us31_U209 (.ZN( us31_n629 ) , .A2( us31_n728 ) , .A1( us31_n785 ) );
  INV_X1 us31_U21 (.A( us31_n749 ) , .ZN( us31_n863 ) );
  NOR2_X1 us31_U210 (.ZN( us31_n611 ) , .A2( us31_n780 ) , .A1( us31_n806 ) );
  NOR2_X1 us31_U211 (.ZN( us31_n652 ) , .A1( us31_n669 ) , .A2( us31_n814 ) );
  NOR2_X1 us31_U212 (.A1( us31_n669 ) , .ZN( us31_n673 ) , .A2( us31_n744 ) );
  NOR2_X1 us31_U213 (.ZN( us31_n602 ) , .A1( us31_n669 ) , .A2( us31_n803 ) );
  NOR2_X1 us31_U214 (.A1( us31_n669 ) , .ZN( us31_n688 ) , .A2( us31_n816 ) );
  NOR2_X1 us31_U215 (.ZN( us31_n628 ) , .A2( us31_n669 ) , .A1( us31_n785 ) );
  INV_X1 us31_U216 (.A( us31_n747 ) , .ZN( us31_n834 ) );
  NOR2_X1 us31_U217 (.A1( us31_n669 ) , .ZN( us31_n766 ) , .A2( us31_n813 ) );
  NOR2_X1 us31_U218 (.A2( us31_n744 ) , .ZN( us31_n769 ) , .A1( us31_n812 ) );
  NOR2_X1 us31_U219 (.ZN( us31_n527 ) , .A1( us31_n669 ) , .A2( us31_n779 ) );
  AOI222_X1 us31_U22 (.ZN( us31_n605 ) , .B2( us31_n671 ) , .B1( us31_n753 ) , .C2( us31_n831 ) , .A1( us31_n833 ) , .A2( us31_n862 ) , .C1( us31_n863 ) );
  NOR2_X1 us31_U220 (.ZN( us31_n531 ) , .A2( us31_n780 ) , .A1( us31_n816 ) );
  INV_X1 us31_U221 (.A( us31_n792 ) , .ZN( us31_n851 ) );
  NOR2_X1 us31_U222 (.A2( us31_n708 ) , .A1( us31_n750 ) , .ZN( us31_n771 ) );
  NOR2_X1 us31_U223 (.ZN( us31_n599 ) , .A2( us31_n791 ) , .A1( us31_n816 ) );
  NOR2_X1 us31_U224 (.ZN( us31_n601 ) , .A2( us31_n780 ) , .A1( us31_n803 ) );
  NOR2_X1 us31_U225 (.A1( us31_n699 ) , .ZN( us31_n768 ) , .A2( us31_n813 ) );
  NOR2_X1 us31_U226 (.ZN( us31_n541 ) , .A2( us31_n697 ) , .A1( us31_n699 ) );
  NOR2_X1 us31_U227 (.ZN( us31_n667 ) , .A1( us31_n750 ) , .A2( us31_n815 ) );
  NOR2_X1 us31_U228 (.ZN( us31_n555 ) , .A1( us31_n750 ) , .A2( us31_n791 ) );
  NOR2_X1 us31_U229 (.ZN( us31_n508 ) , .A2( us31_n780 ) , .A1( us31_n785 ) );
  AOI222_X1 us31_U23 (.ZN( us31_n563 ) , .B1( us31_n830 ) , .C1( us31_n841 ) , .A2( us31_n843 ) , .A1( us31_n854 ) , .B2( us31_n863 ) , .C2( us31_n873 ) );
  NOR2_X1 us31_U230 (.ZN( us31_n543 ) , .A2( us31_n708 ) , .A1( us31_n785 ) );
  NOR2_X1 us31_U231 (.ZN( us31_n528 ) , .A2( us31_n724 ) , .A1( us31_n803 ) );
  NOR2_X1 us31_U232 (.ZN( us31_n664 ) , .A1( us31_n785 ) , .A2( us31_n791 ) );
  NOR2_X1 us31_U233 (.ZN( us31_n556 ) , .A1( us31_n762 ) , .A2( us31_n805 ) );
  INV_X1 us31_U234 (.A( us31_n806 ) , .ZN( us31_n841 ) );
  OAI22_X1 us31_U235 (.B1( us31_n440 ) , .ZN( us31_n444 ) , .A2( us31_n728 ) , .A1( us31_n744 ) , .B2( us31_n749 ) );
  NOR3_X1 us31_U236 (.ZN( us31_n440 ) , .A2( us31_n836 ) , .A3( us31_n837 ) , .A1( us31_n846 ) );
  NOR2_X1 us31_U237 (.ZN( us31_n507 ) , .A1( us31_n812 ) , .A2( us31_n817 ) );
  NOR2_X1 us31_U238 (.ZN( us31_n557 ) , .A1( us31_n792 ) , .A2( us31_n814 ) );
  NOR2_X1 us31_U239 (.ZN( us31_n545 ) , .A1( us31_n749 ) , .A2( us31_n814 ) );
  AOI222_X1 us31_U24 (.ZN( us31_n660 ) , .A2( us31_n839 ) , .B1( us31_n841 ) , .C2( us31_n845 ) , .A1( us31_n860 ) , .C1( us31_n863 ) , .B2( us31_n870 ) );
  OAI22_X1 us31_U240 (.B2( us31_n750 ) , .B1( us31_n751 ) , .A1( us31_n752 ) , .ZN( us31_n756 ) , .A2( us31_n806 ) );
  NOR2_X1 us31_U241 (.ZN( us31_n751 ) , .A2( us31_n852 ) , .A1( us31_n860 ) );
  NOR3_X1 us31_U242 (.ZN( us31_n752 ) , .A2( us31_n853 ) , .A1( us31_n863 ) , .A3( us31_n865 ) );
  NOR2_X1 us31_U243 (.ZN( us31_n544 ) , .A2( us31_n785 ) , .A1( us31_n792 ) );
  NOR2_X1 us31_U244 (.ZN( us31_n530 ) , .A2( us31_n744 ) , .A1( us31_n792 ) );
  NOR2_X1 us31_U245 (.ZN( us31_n509 ) , .A1( us31_n729 ) , .A2( us31_n779 ) );
  NOR2_X1 us31_U246 (.ZN( us31_n570 ) , .A1( us31_n728 ) , .A2( us31_n806 ) );
  NOR2_X1 us31_U247 (.ZN( us31_n666 ) , .A1( us31_n728 ) , .A2( us31_n803 ) );
  NOR2_X1 us31_U248 (.ZN( us31_n631 ) , .A1( us31_n724 ) , .A2( us31_n813 ) );
  NOR2_X1 us31_U249 (.ZN( us31_n614 ) , .A1( us31_n762 ) , .A2( us31_n812 ) );
  INV_X1 us31_U25 (.A( us31_n647 ) , .ZN( us31_n870 ) );
  NOR2_X1 us31_U250 (.A1( us31_n749 ) , .ZN( us31_n767 ) , .A2( us31_n803 ) );
  NOR2_X1 us31_U251 (.ZN( us31_n654 ) , .A1( us31_n728 ) , .A2( us31_n813 ) );
  NOR2_X1 us31_U252 (.ZN( us31_n516 ) , .A1( us31_n708 ) , .A2( us31_n744 ) );
  NOR2_X1 us31_U253 (.ZN( us31_n670 ) , .A1( us31_n790 ) , .A2( us31_n805 ) );
  NOR2_X1 us31_U254 (.ZN( us31_n558 ) , .A1( us31_n708 ) , .A2( us31_n816 ) );
  INV_X1 us31_U255 (.A( us31_n763 ) , .ZN( us31_n866 ) );
  NOR2_X1 us31_U256 (.ZN( us31_n663 ) , .A1( us31_n729 ) , .A2( us31_n785 ) );
  NOR2_X1 us31_U257 (.A2( us31_n697 ) , .ZN( us31_n716 ) , .A1( us31_n792 ) );
  NOR2_X1 us31_U258 (.ZN( us31_n517 ) , .A1( us31_n708 ) , .A2( us31_n803 ) );
  NOR2_X1 us31_U259 (.ZN( us31_n521 ) , .A1( us31_n790 ) , .A2( us31_n812 ) );
  NOR4_X1 us31_U26 (.A4( us31_n544 ) , .A3( us31_n545 ) , .A2( us31_n546 ) , .A1( us31_n547 ) , .ZN( us31_n548 ) );
  NOR2_X1 us31_U260 (.ZN( us31_n630 ) , .A1( us31_n747 ) , .A2( us31_n815 ) );
  NOR2_X1 us31_U261 (.ZN( us31_n655 ) , .A1( us31_n790 ) , .A2( us31_n815 ) );
  AOI21_X1 us31_U262 (.ZN( us31_n552 ) , .B1( us31_n669 ) , .A( us31_n697 ) , .B2( us31_n805 ) );
  NOR2_X1 us31_U263 (.ZN( us31_n668 ) , .A2( us31_n708 ) , .A1( us31_n790 ) );
  NOR2_X1 us31_U264 (.ZN( us31_n594 ) , .A2( us31_n697 ) , .A1( us31_n728 ) );
  NOR2_X1 us31_U265 (.ZN( us31_n542 ) , .A1( us31_n762 ) , .A2( us31_n791 ) );
  NOR2_X1 us31_U266 (.ZN( us31_n656 ) , .A1( us31_n747 ) , .A2( us31_n780 ) );
  NOR2_X1 us31_U267 (.ZN( us31_n609 ) , .A2( us31_n724 ) , .A1( us31_n817 ) );
  AOI21_X1 us31_U268 (.B1( us31_n625 ) , .ZN( us31_n627 ) , .A( us31_n763 ) , .B2( us31_n814 ) );
  NOR2_X1 us31_U269 (.ZN( us31_n661 ) , .A1( us31_n729 ) , .A2( us31_n790 ) );
  NOR4_X1 us31_U27 (.ZN( us31_n479 ) , .A1( us31_n520 ) , .A4( us31_n557 ) , .A3( us31_n582 ) , .A2( us31_n630 ) );
  NOR2_X1 us31_U270 (.ZN( us31_n642 ) , .A2( us31_n788 ) , .A1( us31_n791 ) );
  AOI21_X1 us31_U271 (.ZN( us31_n650 ) , .A( us31_n779 ) , .B1( us31_n792 ) , .B2( us31_n805 ) );
  AOI21_X1 us31_U272 (.ZN( us31_n626 ) , .B2( us31_n669 ) , .A( us31_n790 ) , .B1( us31_n791 ) );
  AOI21_X1 us31_U273 (.A( us31_n815 ) , .B2( us31_n816 ) , .B1( us31_n817 ) , .ZN( us31_n818 ) );
  NOR2_X1 us31_U274 (.ZN( us31_n579 ) , .A2( us31_n708 ) , .A1( us31_n730 ) );
  NOR2_X1 us31_U275 (.ZN( us31_n533 ) , .A2( us31_n724 ) , .A1( us31_n730 ) );
  AOI21_X1 us31_U276 (.A( us31_n812 ) , .B2( us31_n813 ) , .B1( us31_n814 ) , .ZN( us31_n819 ) );
  NOR2_X1 us31_U277 (.A2( us31_n708 ) , .A1( us31_n762 ) , .ZN( us31_n794 ) );
  NOR2_X1 us31_U278 (.A2( us31_n697 ) , .A1( us31_n780 ) , .ZN( us31_n820 ) );
  AOI21_X1 us31_U279 (.ZN( us31_n499 ) , .B1( us31_n680 ) , .A( us31_n812 ) , .B2( us31_n816 ) );
  NOR4_X1 us31_U28 (.ZN( us31_n456 ) , .A2( us31_n517 ) , .A1( us31_n543 ) , .A3( us31_n579 ) , .A4( us31_n615 ) );
  NOR2_X1 us31_U280 (.ZN( us31_n520 ) , .A2( us31_n708 ) , .A1( us31_n814 ) );
  AOI21_X1 us31_U281 (.ZN( us31_n477 ) , .A( us31_n669 ) , .B1( us31_n750 ) , .B2( us31_n806 ) );
  NOR2_X1 us31_U282 (.ZN( us31_n582 ) , .A1( us31_n744 ) , .A2( us31_n815 ) );
  NOR2_X1 us31_U283 (.ZN( us31_n662 ) , .A2( us31_n697 ) , .A1( us31_n729 ) );
  AOI21_X1 us31_U284 (.ZN( us31_n593 ) , .B1( us31_n750 ) , .A( us31_n792 ) , .B2( us31_n813 ) );
  AOI21_X1 us31_U285 (.ZN( us31_n515 ) , .A( us31_n729 ) , .B1( us31_n750 ) , .B2( us31_n803 ) );
  AOI21_X1 us31_U286 (.ZN( us31_n510 ) , .B2( us31_n669 ) , .A( us31_n730 ) , .B1( us31_n815 ) );
  NOR2_X1 us31_U287 (.ZN( us31_n506 ) , .A2( us31_n728 ) , .A1( us31_n762 ) );
  NOR2_X1 us31_U288 (.A1( us31_n697 ) , .ZN( us31_n770 ) , .A2( us31_n815 ) );
  NOR2_X1 us31_U289 (.ZN( us31_n519 ) , .A2( us31_n699 ) , .A1( us31_n816 ) );
  NOR4_X1 us31_U29 (.A4( us31_n532 ) , .A3( us31_n533 ) , .A2( us31_n534 ) , .ZN( us31_n535 ) , .A1( us31_n820 ) );
  NOR2_X1 us31_U290 (.ZN( us31_n581 ) , .A1( us31_n669 ) , .A2( us31_n788 ) );
  NOR2_X1 us31_U291 (.ZN( us31_n559 ) , .A2( us31_n791 ) , .A1( us31_n803 ) );
  AOI21_X1 us31_U292 (.B1( us31_n699 ) , .ZN( us31_n700 ) , .A( us31_n732 ) , .B2( us31_n763 ) );
  AOI21_X1 us31_U293 (.ZN( us31_n591 ) , .B2( us31_n763 ) , .A( us31_n785 ) , .B1( us31_n812 ) );
  INV_X1 us31_U294 (.A( us31_n813 ) , .ZN( us31_n836 ) );
  NOR2_X1 us31_U295 (.ZN( us31_n683 ) , .A2( us31_n699 ) , .A1( us31_n803 ) );
  AOI21_X1 us31_U296 (.ZN( us31_n589 ) , .B2( us31_n699 ) , .B1( us31_n815 ) , .A( us31_n817 ) );
  AOI21_X1 us31_U297 (.ZN( us31_n539 ) , .B2( us31_n812 ) , .A( us31_n814 ) , .B1( us31_n815 ) );
  INV_X1 us31_U298 (.A( us31_n728 ) , .ZN( us31_n852 ) );
  AOI21_X1 us31_U299 (.ZN( us31_n540 ) , .A( us31_n763 ) , .B2( us31_n779 ) , .B1( us31_n817 ) );
  NAND2_X1 us31_U3 (.A1( us31_n449 ) , .A2( us31_n460 ) , .ZN( us31_n792 ) );
  NOR4_X1 us31_U30 (.ZN( us31_n474 ) , .A1( us31_n506 ) , .A3( us31_n544 ) , .A2( us31_n583 ) , .A4( us31_n716 ) );
  INV_X1 us31_U300 (.A( us31_n791 ) , .ZN( us31_n873 ) );
  AOI21_X1 us31_U301 (.ZN( us31_n498 ) , .A( us31_n724 ) , .B2( us31_n762 ) , .B1( us31_n814 ) );
  AOI21_X1 us31_U302 (.ZN( us31_n649 ) , .B1( us31_n729 ) , .B2( us31_n763 ) , .A( us31_n813 ) );
  NOR2_X1 us31_U303 (.ZN( us31_n547 ) , .A1( us31_n699 ) , .A2( us31_n744 ) );
  NOR2_X1 us31_U304 (.ZN( us31_n566 ) , .A2( us31_n697 ) , .A1( us31_n763 ) );
  AOI21_X1 us31_U305 (.ZN( us31_n569 ) , .B1( us31_n750 ) , .B2( us31_n762 ) , .A( us31_n780 ) );
  AOI21_X1 us31_U306 (.ZN( us31_n571 ) , .B2( us31_n697 ) , .B1( us31_n806 ) , .A( us31_n812 ) );
  AOI21_X1 us31_U307 (.ZN( us31_n640 ) , .B2( us31_n747 ) , .A( us31_n792 ) , .B1( us31_n803 ) );
  INV_X1 us31_U308 (.A( us31_n699 ) , .ZN( us31_n853 ) );
  AOI21_X1 us31_U309 (.ZN( us31_n514 ) , .A( us31_n779 ) , .B2( us31_n792 ) , .B1( us31_n812 ) );
  AOI221_X1 us31_U31 (.A( us31_n713 ) , .B2( us31_n714 ) , .ZN( us31_n720 ) , .C1( us31_n832 ) , .B1( us31_n839 ) , .C2( us31_n863 ) );
  AOI21_X1 us31_U310 (.ZN( us31_n639 ) , .B2( us31_n749 ) , .A( us31_n788 ) , .B1( us31_n812 ) );
  NAND2_X1 us31_U311 (.ZN( us31_n753 ) , .A1( us31_n763 ) , .A2( us31_n805 ) );
  NOR2_X1 us31_U312 (.ZN( us31_n665 ) , .A1( us31_n780 ) , .A2( us31_n813 ) );
  INV_X1 us31_U313 (.A( us31_n729 ) , .ZN( us31_n868 ) );
  NOR2_X1 us31_U314 (.ZN( us31_n685 ) , .A1( us31_n729 ) , .A2( us31_n816 ) );
  AOI21_X1 us31_U315 (.ZN( us31_n564 ) , .B1( us31_n724 ) , .A( us31_n779 ) , .B2( us31_n791 ) );
  AOI21_X1 us31_U316 (.ZN( us31_n497 ) , .A( us31_n779 ) , .B2( us31_n791 ) , .B1( us31_n804 ) );
  AOI21_X1 us31_U317 (.ZN( us31_n689 ) , .B2( us31_n749 ) , .B1( us31_n763 ) , .A( us31_n806 ) );
  AOI21_X1 us31_U318 (.ZN( us31_n450 ) , .B2( us31_n792 ) , .A( us31_n803 ) , .B1( us31_n815 ) );
  NOR2_X1 us31_U319 (.ZN( us31_n567 ) , .A1( us31_n747 ) , .A2( us31_n805 ) );
  OR2_X1 us31_U32 (.A2( us31_n711 ) , .A1( us31_n712 ) , .ZN( us31_n713 ) );
  NOR2_X1 us31_U320 (.ZN( us31_n529 ) , .A1( us31_n708 ) , .A2( us31_n779 ) );
  NOR2_X1 us31_U321 (.ZN( us31_n578 ) , .A1( us31_n708 ) , .A2( us31_n813 ) );
  AOI21_X1 us31_U322 (.ZN( us31_n478 ) , .B2( us31_n697 ) , .A( us31_n749 ) , .B1( us31_n779 ) );
  AOI21_X1 us31_U323 (.A( us31_n790 ) , .B2( us31_n791 ) , .B1( us31_n792 ) , .ZN( us31_n793 ) );
  NOR2_X1 us31_U324 (.ZN( us31_n684 ) , .A1( us31_n791 ) , .A2( us31_n813 ) );
  AOI21_X1 us31_U325 (.A( us31_n733 ) , .ZN( us31_n734 ) , .B2( us31_n780 ) , .B1( us31_n792 ) );
  NOR2_X1 us31_U326 (.A2( us31_n813 ) , .A1( us31_n815 ) , .ZN( us31_n821 ) );
  NOR2_X1 us31_U327 (.ZN( us31_n711 ) , .A1( us31_n762 ) , .A2( us31_n763 ) );
  AOI21_X1 us31_U328 (.ZN( us31_n641 ) , .B1( us31_n680 ) , .A( us31_n791 ) , .B2( us31_n817 ) );
  NOR2_X1 us31_U329 (.ZN( us31_n580 ) , .A2( us31_n697 ) , .A1( us31_n791 ) );
  NOR2_X1 us31_U33 (.ZN( us31_n680 ) , .A2( us31_n834 ) , .A1( us31_n839 ) );
  NOR2_X1 us31_U330 (.ZN( us31_n583 ) , .A1( us31_n792 ) , .A2( us31_n817 ) );
  NOR2_X1 us31_U331 (.ZN( us31_n534 ) , .A1( us31_n724 ) , .A2( us31_n788 ) );
  NOR2_X1 us31_U332 (.ZN( us31_n632 ) , .A2( us31_n697 ) , .A1( us31_n724 ) );
  NOR2_X1 us31_U333 (.ZN( us31_n682 ) , .A2( us31_n708 ) , .A1( us31_n817 ) );
  AOI21_X1 us31_U334 (.B1( us31_n686 ) , .ZN( us31_n687 ) , .A( us31_n728 ) , .B2( us31_n761 ) );
  INV_X1 us31_U335 (.A( us31_n815 ) , .ZN( us31_n855 ) );
  AOI21_X1 us31_U336 (.ZN( us31_n442 ) , .A( us31_n699 ) , .B1( us31_n733 ) , .B2( us31_n750 ) );
  NOR2_X1 us31_U337 (.ZN( us31_n568 ) , .A1( us31_n729 ) , .A2( us31_n762 ) );
  INV_X1 us31_U338 (.A( us31_n780 ) , .ZN( us31_n850 ) );
  INV_X1 us31_U339 (.A( us31_n785 ) , .ZN( us31_n846 ) );
  AOI222_X1 us31_U34 (.ZN( us31_n469 ) , .B1( us31_n832 ) , .A1( us31_n839 ) , .C1( us31_n842 ) , .C2( us31_n851 ) , .A2( us31_n855 ) , .B2( us31_n865 ) );
  NAND2_X1 us31_U340 (.A2( us31_n762 ) , .A1( us31_n806 ) , .ZN( us31_n810 ) );
  AOI21_X1 us31_U341 (.ZN( us31_n443 ) , .B1( us31_n789 ) , .B2( us31_n791 ) , .A( us31_n814 ) );
  NAND2_X1 us31_U342 (.ZN( us31_n671 ) , .A1( us31_n806 ) , .A2( us31_n816 ) );
  NOR2_X1 us31_U343 (.ZN( us31_n484 ) , .A1( us31_n788 ) , .A2( us31_n805 ) );
  NOR2_X1 us31_U344 (.ZN( us31_n470 ) , .A2( us31_n779 ) , .A1( us31_n815 ) );
  NOR2_X1 us31_U345 (.ZN( us31_n712 ) , .A2( us31_n724 ) , .A1( us31_n790 ) );
  OAI21_X1 us31_U346 (.A( us31_n787 ) , .B2( us31_n788 ) , .B1( us31_n789 ) , .ZN( us31_n795 ) );
  OAI21_X1 us31_U347 (.ZN( us31_n787 ) , .A( us31_n839 ) , .B1( us31_n863 ) , .B2( us31_n873 ) );
  NOR2_X1 us31_U348 (.ZN( us31_n526 ) , .A1( us31_n724 ) , .A2( us31_n750 ) );
  NAND2_X1 us31_U349 (.A1( us31_n699 ) , .A2( us31_n729 ) , .ZN( us31_n782 ) );
  NOR4_X1 us31_U35 (.A1( us31_n466 ) , .ZN( us31_n467 ) , .A4( us31_n542 ) , .A2( us31_n554 ) , .A3( us31_n614 ) );
  NOR2_X1 us31_U350 (.ZN( us31_n518 ) , .A1( us31_n708 ) , .A2( us31_n788 ) );
  OAI21_X1 us31_U351 (.A( us31_n698 ) , .ZN( us31_n702 ) , .B2( us31_n750 ) , .B1( us31_n804 ) );
  OAI21_X1 us31_U352 (.ZN( us31_n698 ) , .B2( us31_n833 ) , .B1( us31_n838 ) , .A( us31_n860 ) );
  INV_X1 us31_U353 (.A( us31_n817 ) , .ZN( us31_n844 ) );
  OAI21_X1 us31_U354 (.A( us31_n731 ) , .B1( us31_n732 ) , .ZN( us31_n736 ) , .B2( us31_n805 ) );
  OAI21_X1 us31_U355 (.ZN( us31_n731 ) , .A( us31_n833 ) , .B2( us31_n852 ) , .B1( us31_n873 ) );
  NAND2_X1 us31_U356 (.ZN( us31_n714 ) , .A1( us31_n728 ) , .A2( us31_n780 ) );
  INV_X1 us31_U357 (.A( us31_n724 ) , .ZN( us31_n856 ) );
  AND2_X1 us31_U358 (.ZN( us31_n732 ) , .A1( us31_n779 ) , .A2( us31_n785 ) );
  NAND2_X1 us31_U359 (.A1( us31_n447 ) , .A2( us31_n449 ) , .ZN( us31_n805 ) );
  AOI221_X1 us31_U36 (.ZN( us31_n468 ) , .C2( us31_n714 ) , .B2( us31_n831 ) , .C1( us31_n845 ) , .B1( us31_n860 ) , .A( us31_n864 ) );
  NAND2_X1 us31_U360 (.A1( us31_n451 ) , .A2( us31_n454 ) , .ZN( us31_n814 ) );
  NAND2_X1 us31_U361 (.A1( us31_n452 ) , .A2( us31_n465 ) , .ZN( us31_n669 ) );
  NAND2_X1 us31_U362 (.A1( us31_n455 ) , .A2( us31_n462 ) , .ZN( us31_n750 ) );
  NAND2_X1 us31_U363 (.A2( us31_n453 ) , .A1( us31_n455 ) , .ZN( us31_n806 ) );
  NAND2_X1 us31_U364 (.A1( us31_n451 ) , .A2( us31_n471 ) , .ZN( us31_n816 ) );
  NAND2_X1 us31_U365 (.A1( us31_n454 ) , .A2( us31_n461 ) , .ZN( us31_n813 ) );
  NAND2_X1 us31_U366 (.A1( us31_n455 ) , .A2( us31_n471 ) , .ZN( us31_n803 ) );
  NAND2_X1 us31_U367 (.A1( us31_n453 ) , .A2( us31_n461 ) , .ZN( us31_n744 ) );
  NAND2_X1 us31_U368 (.A1( us31_n453 ) , .A2( us31_n472 ) , .ZN( us31_n785 ) );
  NAND2_X1 us31_U369 (.A2( us31_n454 ) , .A1( us31_n472 ) , .ZN( us31_n779 ) );
  NOR4_X1 us31_U37 (.A4( us31_n577 ) , .A3( us31_n578 ) , .A2( us31_n579 ) , .ZN( us31_n586 ) , .A1( us31_n683 ) );
  NAND2_X1 us31_U370 (.A2( us31_n464 ) , .A1( us31_n465 ) , .ZN( us31_n812 ) );
  NAND2_X1 us31_U371 (.A1( us31_n441 ) , .A2( us31_n460 ) , .ZN( us31_n699 ) );
  NAND2_X1 us31_U372 (.A2( us31_n449 ) , .A1( us31_n452 ) , .ZN( us31_n763 ) );
  NAND2_X1 us31_U373 (.A2( us31_n461 ) , .A1( us31_n462 ) , .ZN( us31_n747 ) );
  NAND2_X1 us31_U374 (.A1( us31_n462 ) , .A2( us31_n472 ) , .ZN( us31_n788 ) );
  NOR2_X1 us31_U375 (.ZN( us31_n465 ) , .A2( us31_n847 ) , .A1( us31_n848 ) );
  NOR2_X1 us31_U376 (.ZN( us31_n453 ) , .A1( us31_n826 ) , .A2( us31_n827 ) );
  NOR2_X1 us31_U377 (.ZN( us31_n451 ) , .A1( us31_n828 ) , .A2( us31_n829 ) );
  NAND2_X1 us31_U378 (.A1( us31_n451 ) , .A2( us31_n462 ) , .ZN( us31_n790 ) );
  NAND2_X1 us31_U379 (.A2( us31_n441 ) , .A1( us31_n447 ) , .ZN( us31_n784 ) );
  NOR4_X1 us31_U38 (.A1( us31_n584 ) , .ZN( us31_n585 ) , .A3( us31_n652 ) , .A2( us31_n662 ) , .A4( us31_n767 ) );
  NAND2_X1 us31_U380 (.A2( us31_n454 ) , .A1( us31_n455 ) , .ZN( us31_n730 ) );
  NAND2_X2 us31_U381 (.A1( us31_n449 ) , .A2( us31_n464 ) , .ZN( us31_n724 ) );
  NAND2_X2 us31_U382 (.A2( us31_n460 ) , .A1( us31_n465 ) , .ZN( us31_n780 ) );
  NOR2_X1 us31_U383 (.ZN( us31_n447 ) , .A2( us31_n849 ) , .A1( us31_n858 ) );
  NAND2_X1 us31_U384 (.A1( us31_n447 ) , .A2( us31_n448 ) , .ZN( us31_n786 ) );
  NAND2_X1 us31_U385 (.A2( us31_n448 ) , .A1( us31_n460 ) , .ZN( us31_n728 ) );
  NAND2_X1 us31_U386 (.A2( us31_n448 ) , .A1( us31_n452 ) , .ZN( us31_n729 ) );
  NOR2_X1 us31_U387 (.A2( sa31_5 ) , .ZN( us31_n448 ) , .A1( us31_n847 ) );
  NOR2_X1 us31_U388 (.A2( sa31_7 ) , .ZN( us31_n460 ) , .A1( us31_n849 ) );
  NOR2_X1 us31_U389 (.A2( sa31_6 ) , .A1( sa31_7 ) , .ZN( us31_n464 ) );
  NOR4_X1 us31_U39 (.ZN( us31_n620 ) , .A1( us31_n656 ) , .A3( us31_n666 ) , .A4( us31_n682 ) , .A2( us31_n766 ) );
  NOR2_X1 us31_U390 (.A2( sa31_4 ) , .ZN( us31_n449 ) , .A1( us31_n848 ) );
  NOR2_X1 us31_U391 (.A2( sa31_4 ) , .A1( sa31_5 ) , .ZN( us31_n441 ) );
  NOR2_X1 us31_U392 (.A2( sa31_6 ) , .ZN( us31_n452 ) , .A1( us31_n858 ) );
  NOR2_X1 us31_U393 (.A2( sa31_2 ) , .A1( sa31_3 ) , .ZN( us31_n472 ) );
  NOR2_X1 us31_U394 (.A2( sa31_1 ) , .ZN( us31_n471 ) , .A1( us31_n826 ) );
  NOR2_X1 us31_U395 (.A2( sa31_0 ) , .ZN( us31_n454 ) , .A1( us31_n827 ) );
  NOR2_X1 us31_U396 (.A2( sa31_0 ) , .A1( sa31_1 ) , .ZN( us31_n462 ) );
  NOR2_X1 us31_U397 (.A2( sa31_3 ) , .ZN( us31_n455 ) , .A1( us31_n828 ) );
  NOR2_X1 us31_U398 (.A2( sa31_2 ) , .ZN( us31_n461 ) , .A1( us31_n829 ) );
  INV_X1 us31_U399 (.A( sa31_4 ) , .ZN( us31_n847 ) );
  NAND2_X1 us31_U4 (.A2( us31_n448 ) , .A1( us31_n464 ) , .ZN( us31_n815 ) );
  NOR4_X1 us31_U40 (.A4( us31_n609 ) , .A3( us31_n610 ) , .A2( us31_n611 ) , .A1( us31_n612 ) , .ZN( us31_n619 ) );
  INV_X1 us31_U400 (.A( sa31_6 ) , .ZN( us31_n849 ) );
  INV_X1 us31_U401 (.A( sa31_3 ) , .ZN( us31_n829 ) );
  INV_X1 us31_U402 (.A( sa31_1 ) , .ZN( us31_n827 ) );
  INV_X1 us31_U403 (.A( sa31_0 ) , .ZN( us31_n826 ) );
  INV_X1 us31_U404 (.A( sa31_2 ) , .ZN( us31_n828 ) );
  INV_X1 us31_U405 (.A( sa31_5 ) , .ZN( us31_n848 ) );
  INV_X1 us31_U406 (.A( sa31_7 ) , .ZN( us31_n858 ) );
  NAND2_X1 us31_U407 (.A2( us31_n461 ) , .A1( us31_n471 ) , .ZN( us31_n697 ) );
  OAI22_X1 us31_U408 (.ZN( us31_n588 ) , .A2( us31_n747 ) , .B2( us31_n762 ) , .A1( us31_n763 ) , .B1( us31_n784 ) );
  AOI21_X1 us31_U409 (.ZN( us31_n592 ) , .B1( us31_n728 ) , .B2( us31_n784 ) , .A( us31_n790 ) );
  NOR4_X1 us31_U41 (.A4( us31_n614 ) , .A3( us31_n615 ) , .A2( us31_n616 ) , .A1( us31_n617 ) , .ZN( us31_n618 ) );
  NAND2_X1 us31_U410 (.A1( us31_n729 ) , .A2( us31_n784 ) , .ZN( us31_n811 ) );
  AOI21_X1 us31_U411 (.ZN( us31_n623 ) , .B1( us31_n699 ) , .A( us31_n779 ) , .B2( us31_n784 ) );
  OAI22_X1 us31_U412 (.ZN( us31_n681 ) , .A1( us31_n699 ) , .A2( us31_n730 ) , .B2( us31_n784 ) , .B1( us31_n817 ) );
  AOI21_X1 us31_U413 (.ZN( us31_n648 ) , .A( us31_n762 ) , .B2( us31_n784 ) , .B1( us31_n792 ) );
  OAI21_X1 us31_U414 (.A( us31_n613 ) , .ZN( us31_n616 ) , .B1( us31_n625 ) , .B2( us31_n784 ) );
  OAI222_X1 us31_U415 (.A2( us31_n669 ) , .ZN( us31_n674 ) , .B1( us31_n747 ) , .B2( us31_n784 ) , .C2( us31_n788 ) , .C1( us31_n815 ) , .A1( us31_n817 ) );
  NOR2_X1 us31_U416 (.ZN( us31_n610 ) , .A1( us31_n784 ) , .A2( us31_n816 ) );
  NOR2_X1 us31_U417 (.ZN( us31_n651 ) , .A1( us31_n784 ) , .A2( us31_n788 ) );
  NOR2_X1 us31_U418 (.ZN( us31_n553 ) , .A2( us31_n744 ) , .A1( us31_n784 ) );
  NOR2_X1 us31_U419 (.ZN( us31_n600 ) , .A2( us31_n697 ) , .A1( us31_n784 ) );
  NOR4_X1 us31_U42 (.A4( us31_n514 ) , .A3( us31_n515 ) , .A2( us31_n516 ) , .A1( us31_n517 ) , .ZN( us31_n524 ) );
  INV_X1 us31_U420 (.A( us31_n784 ) , .ZN( us31_n861 ) );
  AND2_X1 us31_U421 (.ZN( us31_n438 ) , .A2( us31_n831 ) , .A1( us31_n854 ) );
  AND2_X1 us31_U422 (.ZN( us31_n439 ) , .A2( us31_n843 ) , .A1( us31_n861 ) );
  NOR3_X1 us31_U423 (.A1( us31_n438 ) , .A2( us31_n439 ) , .A3( us31_n576 ) , .ZN( us31_n587 ) );
  INV_X1 us31_U424 (.A( us31_n812 ) , .ZN( us31_n854 ) );
  INV_X1 us31_U425 (.A( us31_n803 ) , .ZN( us31_n843 ) );
  AOI21_X1 us31_U426 (.ZN( us31_n576 ) , .B2( us31_n724 ) , .B1( us31_n748 ) , .A( us31_n785 ) );
  OAI221_X1 us31_U427 (.A( us31_n783 ) , .C2( us31_n784 ) , .B2( us31_n785 ) , .B1( us31_n786 ) , .ZN( us31_n796 ) , .C1( us31_n813 ) );
  AOI21_X1 us31_U428 (.ZN( us31_n500 ) , .A( us31_n697 ) , .B1( us31_n708 ) , .B2( us31_n786 ) );
  OAI221_X1 us31_U429 (.A( us31_n696 ) , .ZN( us31_n703 ) , .C2( us31_n784 ) , .C1( us31_n785 ) , .B1( us31_n786 ) , .B2( us31_n806 ) );
  AOI222_X1 us31_U43 (.ZN( us31_n525 ) , .A1( us31_n834 ) , .B2( us31_n837 ) , .C1( us31_n844 ) , .C2( us31_n850 ) , .A2( us31_n852 ) , .B1( us31_n866 ) );
  OAI22_X1 us31_U430 (.ZN( us31_n590 ) , .B1( us31_n730 ) , .B2( us31_n749 ) , .A2( us31_n786 ) , .A1( us31_n803 ) );
  NAND2_X1 us31_U431 (.A2( us31_n749 ) , .A1( us31_n786 ) , .ZN( us31_n809 ) );
  NOR2_X1 us31_U432 (.ZN( us31_n612 ) , .A1( us31_n779 ) , .A2( us31_n786 ) );
  OAI222_X1 us31_U433 (.ZN( us31_n617 ) , .B1( us31_n697 ) , .C1( us31_n724 ) , .C2( us31_n747 ) , .B2( us31_n786 ) , .A2( us31_n792 ) , .A1( us31_n816 ) );
  NOR2_X1 us31_U434 (.ZN( us31_n653 ) , .A1( us31_n762 ) , .A2( us31_n786 ) );
  NOR2_X1 us31_U435 (.ZN( us31_n554 ) , .A1( us31_n786 ) , .A2( us31_n813 ) );
  NOR2_X1 us31_U436 (.ZN( us31_n717 ) , .A2( us31_n744 ) , .A1( us31_n786 ) );
  NAND3_X1 us31_U437 (.ZN( sa32_sr_6 ) , .A3( us31_n797 ) , .A2( us31_n798 ) , .A1( us31_n799 ) );
  NAND3_X1 us31_U438 (.ZN( sa32_sr_5 ) , .A3( us31_n758 ) , .A2( us31_n759 ) , .A1( us31_n760 ) );
  NAND3_X1 us31_U439 (.ZN( sa32_sr_4 ) , .A3( us31_n738 ) , .A2( us31_n739 ) , .A1( us31_n740 ) );
  NOR4_X1 us31_U44 (.A3( us31_n521 ) , .A1( us31_n522 ) , .ZN( us31_n523 ) , .A2( us31_n673 ) , .A4( us31_n769 ) );
  NAND3_X1 us31_U440 (.A3( us31_n675 ) , .A2( us31_n676 ) , .A1( us31_n677 ) , .ZN( us31_n807 ) );
  NAND3_X1 us31_U441 (.ZN( us31_n638 ) , .A3( us31_n708 ) , .A2( us31_n724 ) , .A1( us31_n792 ) );
  NAND3_X1 us31_U442 (.A3( us31_n618 ) , .A2( us31_n619 ) , .A1( us31_n620 ) , .ZN( us31_n725 ) );
  NAND3_X1 us31_U443 (.A3( us31_n585 ) , .A2( us31_n586 ) , .A1( us31_n587 ) , .ZN( us31_n621 ) );
  NAND3_X1 us31_U444 (.ZN( us31_n565 ) , .A3( us31_n680 ) , .A2( us31_n750 ) , .A1( us31_n785 ) );
  NAND3_X1 us31_U445 (.A3( us31_n523 ) , .A2( us31_n524 ) , .A1( us31_n525 ) , .ZN( us31_n742 ) );
  NAND3_X1 us31_U446 (.A3( us31_n512 ) , .A1( us31_n513 ) , .ZN( us31_n608 ) , .A2( us31_n871 ) );
  NAND3_X1 us31_U447 (.A3( us31_n467 ) , .A2( us31_n468 ) , .A1( us31_n469 ) , .ZN( us31_n777 ) );
  NOR2_X1 us31_U448 (.ZN( us31_n701 ) , .A2( us31_n786 ) , .A1( us31_n817 ) );
  NOR2_X1 us31_U449 (.A1( us31_n730 ) , .ZN( us31_n765 ) , .A2( us31_n786 ) );
  AOI221_X1 us31_U45 (.A( us31_n781 ) , .ZN( us31_n798 ) , .C2( us31_n837 ) , .B2( us31_n838 ) , .B1( us31_n865 ) , .C1( us31_n866 ) );
  NOR4_X1 us31_U46 (.A4( us31_n793 ) , .A3( us31_n794 ) , .A2( us31_n795 ) , .A1( us31_n796 ) , .ZN( us31_n797 ) );
  NOR4_X1 us31_U47 (.A4( us31_n776 ) , .A3( us31_n777 ) , .A1( us31_n778 ) , .ZN( us31_n799 ) , .A2( us31_n801 ) );
  NOR4_X1 us31_U48 (.A3( us31_n755 ) , .A2( us31_n756 ) , .A1( us31_n757 ) , .ZN( us31_n758 ) , .A4( us31_n869 ) );
  AOI211_X1 us31_U49 (.B( us31_n745 ) , .A( us31_n746 ) , .ZN( us31_n759 ) , .C1( us31_n832 ) , .C2( us31_n853 ) );
  NAND2_X1 us31_U5 (.A1( us31_n441 ) , .A2( us31_n464 ) , .ZN( us31_n708 ) );
  NOR3_X1 us31_U50 (.A3( us31_n741 ) , .A2( us31_n742 ) , .A1( us31_n743 ) , .ZN( us31_n760 ) );
  NAND4_X1 us31_U51 (.ZN( sa32_sr_3 ) , .A4( us31_n704 ) , .A3( us31_n705 ) , .A2( us31_n706 ) , .A1( us31_n707 ) );
  NOR4_X1 us31_U52 (.A4( us31_n700 ) , .A3( us31_n701 ) , .A2( us31_n702 ) , .A1( us31_n703 ) , .ZN( us31_n704 ) );
  AOI211_X1 us31_U53 (.B( us31_n694 ) , .A( us31_n695 ) , .ZN( us31_n705 ) , .C2( us31_n831 ) , .C1( us31_n851 ) );
  NOR2_X1 us31_U54 (.ZN( us31_n707 ) , .A2( us31_n776 ) , .A1( us31_n800 ) );
  NOR2_X1 us31_U55 (.ZN( us31_n804 ) , .A1( us31_n854 ) , .A2( us31_n861 ) );
  NAND4_X1 us31_U56 (.ZN( sa32_sr_7 ) , .A4( us31_n822 ) , .A3( us31_n823 ) , .A2( us31_n824 ) , .A1( us31_n825 ) );
  NOR4_X1 us31_U57 (.A4( us31_n818 ) , .A3( us31_n819 ) , .A2( us31_n820 ) , .A1( us31_n821 ) , .ZN( us31_n822 ) );
  AOI222_X1 us31_U58 (.C2( us31_n809 ) , .B2( us31_n810 ) , .A2( us31_n811 ) , .ZN( us31_n823 ) , .C1( us31_n832 ) , .A1( us31_n839 ) , .B1( us31_n853 ) );
  AOI211_X1 us31_U59 (.B( us31_n807 ) , .A( us31_n808 ) , .ZN( us31_n824 ) , .C1( us31_n842 ) , .C2( us31_n850 ) );
  NAND2_X1 us31_U6 (.A2( us31_n441 ) , .A1( us31_n452 ) , .ZN( us31_n791 ) );
  NAND4_X1 us31_U60 (.ZN( sa32_sr_0 ) , .A4( us31_n501 ) , .A3( us31_n502 ) , .A2( us31_n503 ) , .A1( us31_n504 ) );
  AOI221_X1 us31_U61 (.A( us31_n497 ) , .ZN( us31_n502 ) , .B2( us31_n843 ) , .C1( us31_n846 ) , .C2( us31_n860 ) , .B1( us31_n862 ) );
  NOR4_X1 us31_U62 (.A4( us31_n498 ) , .A3( us31_n499 ) , .A2( us31_n500 ) , .ZN( us31_n501 ) , .A1( us31_n527 ) );
  AOI211_X1 us31_U63 (.A( us31_n496 ) , .ZN( us31_n503 ) , .B( us31_n802 ) , .C2( us31_n839 ) , .C1( us31_n851 ) );
  NAND4_X1 us31_U64 (.ZN( sa32_sr_1 ) , .A4( us31_n595 ) , .A3( us31_n596 ) , .A2( us31_n597 ) , .A1( us31_n598 ) );
  NOR4_X1 us31_U65 (.A4( us31_n591 ) , .A3( us31_n592 ) , .A2( us31_n593 ) , .A1( us31_n594 ) , .ZN( us31_n595 ) );
  AOI211_X1 us31_U66 (.B( us31_n589 ) , .A( us31_n590 ) , .ZN( us31_n596 ) , .C2( us31_n811 ) , .C1( us31_n833 ) );
  AOI211_X1 us31_U67 (.A( us31_n588 ) , .ZN( us31_n597 ) , .B( us31_n621 ) , .C1( us31_n845 ) , .C2( us31_n855 ) );
  NAND4_X1 us31_U68 (.ZN( sa32_sr_2 ) , .A4( us31_n643 ) , .A3( us31_n644 ) , .A2( us31_n645 ) , .A1( us31_n646 ) );
  AOI222_X1 us31_U69 (.B2( us31_n638 ) , .ZN( us31_n644 ) , .B1( us31_n841 ) , .A1( us31_n842 ) , .C2( us31_n846 ) , .C1( us31_n863 ) , .A2( us31_n865 ) );
  NAND2_X1 us31_U7 (.A2( us31_n471 ) , .A1( us31_n472 ) , .ZN( us31_n817 ) );
  NOR4_X1 us31_U70 (.A4( us31_n639 ) , .A3( us31_n640 ) , .A2( us31_n641 ) , .A1( us31_n642 ) , .ZN( us31_n643 ) );
  NOR3_X1 us31_U71 (.A2( us31_n607 ) , .A1( us31_n608 ) , .ZN( us31_n646 ) , .A3( us31_n722 ) );
  NOR2_X1 us31_U72 (.ZN( us31_n748 ) , .A1( us31_n861 ) , .A2( us31_n862 ) );
  NOR2_X1 us31_U73 (.ZN( us31_n625 ) , .A2( us31_n836 ) , .A1( us31_n839 ) );
  NAND4_X1 us31_U74 (.A4( us31_n603 ) , .A3( us31_n604 ) , .A2( us31_n605 ) , .A1( us31_n606 ) , .ZN( us31_n722 ) );
  NOR3_X1 us31_U75 (.A1( us31_n599 ) , .ZN( us31_n604 ) , .A3( us31_n663 ) , .A2( us31_n770 ) );
  NOR4_X1 us31_U76 (.A3( us31_n600 ) , .A2( us31_n601 ) , .A1( us31_n602 ) , .ZN( us31_n603 ) , .A4( us31_n655 ) );
  AOI222_X1 us31_U77 (.ZN( us31_n606 ) , .A1( us31_n830 ) , .C2( us31_n837 ) , .B1( us31_n842 ) , .A2( us31_n856 ) , .B2( us31_n861 ) , .C1( us31_n868 ) );
  NAND4_X1 us31_U78 (.A4( us31_n657 ) , .A3( us31_n658 ) , .A2( us31_n659 ) , .A1( us31_n660 ) , .ZN( us31_n800 ) );
  NOR3_X1 us31_U79 (.A3( us31_n648 ) , .A2( us31_n649 ) , .A1( us31_n650 ) , .ZN( us31_n659 ) );
  NOR3_X1 us31_U8 (.ZN( us31_n598 ) , .A1( us31_n608 ) , .A3( us31_n723 ) , .A2( us31_n742 ) );
  NOR3_X1 us31_U80 (.A3( us31_n651 ) , .A2( us31_n652 ) , .A1( us31_n653 ) , .ZN( us31_n658 ) );
  NOR3_X1 us31_U81 (.A3( us31_n654 ) , .A2( us31_n655 ) , .A1( us31_n656 ) , .ZN( us31_n657 ) );
  NAND4_X1 us31_U82 (.A4( us31_n560 ) , .A3( us31_n561 ) , .A2( us31_n562 ) , .A1( us31_n563 ) , .ZN( us31_n607 ) );
  NOR4_X1 us31_U83 (.ZN( us31_n561 ) , .A1( us31_n653 ) , .A3( us31_n661 ) , .A4( us31_n685 ) , .A2( us31_n768 ) );
  NOR4_X1 us31_U84 (.A4( us31_n552 ) , .A3( us31_n553 ) , .A2( us31_n554 ) , .A1( us31_n555 ) , .ZN( us31_n562 ) );
  NOR4_X1 us31_U85 (.A4( us31_n556 ) , .A3( us31_n557 ) , .A2( us31_n558 ) , .A1( us31_n559 ) , .ZN( us31_n560 ) );
  NAND4_X1 us31_U86 (.A4( us31_n772 ) , .A3( us31_n773 ) , .A2( us31_n774 ) , .A1( us31_n775 ) , .ZN( us31_n801 ) );
  NOR3_X1 us31_U87 (.A3( us31_n765 ) , .A2( us31_n766 ) , .A1( us31_n767 ) , .ZN( us31_n773 ) );
  NOR4_X1 us31_U88 (.A4( us31_n768 ) , .A3( us31_n769 ) , .A2( us31_n770 ) , .A1( us31_n771 ) , .ZN( us31_n772 ) );
  AOI222_X1 us31_U89 (.ZN( us31_n775 ) , .A1( us31_n830 ) , .C1( us31_n834 ) , .B2( us31_n841 ) , .A2( us31_n850 ) , .B1( us31_n861 ) , .C2( us31_n873 ) );
  NOR3_X1 us31_U9 (.A3( us31_n800 ) , .A2( us31_n801 ) , .A1( us31_n802 ) , .ZN( us31_n825 ) );
  NOR4_X1 us31_U90 (.A4( us31_n661 ) , .A3( us31_n662 ) , .A2( us31_n663 ) , .A1( us31_n664 ) , .ZN( us31_n677 ) );
  NOR4_X1 us31_U91 (.A4( us31_n665 ) , .A3( us31_n666 ) , .A2( us31_n667 ) , .A1( us31_n668 ) , .ZN( us31_n676 ) );
  NOR4_X1 us31_U92 (.A3( us31_n673 ) , .A1( us31_n674 ) , .ZN( us31_n675 ) , .A4( us31_n715 ) , .A2( us31_n859 ) );
  NOR2_X1 us31_U93 (.ZN( us31_n761 ) , .A1( us31_n833 ) , .A2( us31_n834 ) );
  AOI222_X1 us31_U94 (.ZN( us31_n513 ) , .C1( us31_n832 ) , .B2( us31_n837 ) , .A2( us31_n843 ) , .C2( us31_n862 ) , .B1( us31_n863 ) , .A1( us31_n866 ) );
  NOR4_X1 us31_U95 (.A4( us31_n509 ) , .A2( us31_n510 ) , .A1( us31_n511 ) , .ZN( us31_n512 ) , .A3( us31_n670 ) );
  INV_X1 us31_U96 (.A( us31_n505 ) , .ZN( us31_n871 ) );
  NAND4_X1 us31_U97 (.A4( us31_n456 ) , .A3( us31_n457 ) , .A2( us31_n458 ) , .A1( us31_n459 ) , .ZN( us31_n679 ) );
  NOR3_X1 us31_U98 (.ZN( us31_n457 ) , .A3( us31_n530 ) , .A1( us31_n555 ) , .A2( us31_n570 ) );
  AOI221_X1 us31_U99 (.A( us31_n450 ) , .ZN( us31_n459 ) , .C2( us31_n753 ) , .B1( us31_n832 ) , .C1( us31_n842 ) , .B2( us31_n861 ) );
endmodule

