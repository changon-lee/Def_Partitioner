module aes_aes_die_3 ( sa01_0, sa01_1, sa01_2, sa01_3, sa01_4, sa01_5, sa01_6, sa01_7, sa20_0, 
       sa20_1, sa20_2, sa20_3, sa20_4, sa20_5, sa20_6, sa20_7, sa32_0, sa32_1, 
       sa32_2, sa32_3, sa32_4, sa32_5, sa32_6, sa32_7, sa01_sr_0, sa01_sr_1, sa01_sr_2, sa01_sr_3, sa01_sr_4, sa01_sr_5, sa01_sr_6, sa01_sr_7, sa22_sr_0, 
        sa22_sr_1, sa22_sr_2, sa22_sr_3, sa22_sr_4, sa22_sr_5, sa22_sr_6, sa22_sr_7, sa33_sr_0, sa33_sr_1, 
        sa33_sr_2, sa33_sr_3, sa33_sr_4, sa33_sr_5, sa33_sr_6, sa33_sr_7 );
  input sa01_0, sa01_1, sa01_2, sa01_3, sa01_4, sa01_5, sa01_6, sa01_7, sa20_0, 
        sa20_1, sa20_2, sa20_3, sa20_4, sa20_5, sa20_6, sa20_7, sa32_0, sa32_1, 
        sa32_2, sa32_3, sa32_4, sa32_5, sa32_6, sa32_7;
  output sa01_sr_0, sa01_sr_1, sa01_sr_2, sa01_sr_3, sa01_sr_4, sa01_sr_5, sa01_sr_6, sa01_sr_7, sa22_sr_0, 
        sa22_sr_1, sa22_sr_2, sa22_sr_3, sa22_sr_4, sa22_sr_5, sa22_sr_6, sa22_sr_7, sa33_sr_0, sa33_sr_1, 
        sa33_sr_2, sa33_sr_3, sa33_sr_4, sa33_sr_5, sa33_sr_6, sa33_sr_7;
  wire us01_n438, us01_n439, us01_n440, us01_n441, us01_n442, us01_n443, us01_n444, us01_n445, us01_n446, 
       us01_n447, us01_n448, us01_n449, us01_n450, us01_n451, us01_n452, us01_n453, us01_n454, us01_n455, 
       us01_n456, us01_n457, us01_n458, us01_n459, us01_n460, us01_n461, us01_n462, us01_n463, us01_n464, 
       us01_n465, us01_n466, us01_n467, us01_n468, us01_n469, us01_n470, us01_n471, us01_n472, us01_n473, 
       us01_n474, us01_n475, us01_n476, us01_n477, us01_n478, us01_n479, us01_n480, us01_n481, us01_n482, 
       us01_n483, us01_n484, us01_n485, us01_n486, us01_n487, us01_n488, us01_n489, us01_n490, us01_n491, 
       us01_n492, us01_n493, us01_n494, us01_n495, us01_n496, us01_n497, us01_n498, us01_n499, us01_n500, 
       us01_n501, us01_n502, us01_n503, us01_n504, us01_n505, us01_n506, us01_n507, us01_n508, us01_n509, 
       us01_n510, us01_n511, us01_n512, us01_n513, us01_n514, us01_n515, us01_n516, us01_n517, us01_n518, 
       us01_n519, us01_n520, us01_n521, us01_n522, us01_n523, us01_n524, us01_n525, us01_n526, us01_n527, 
       us01_n528, us01_n529, us01_n530, us01_n531, us01_n532, us01_n533, us01_n534, us01_n535, us01_n536, 
       us01_n537, us01_n538, us01_n539, us01_n540, us01_n541, us01_n542, us01_n543, us01_n544, us01_n545, 
       us01_n546, us01_n547, us01_n548, us01_n549, us01_n550, us01_n551, us01_n552, us01_n553, us01_n554, 
       us01_n555, us01_n556, us01_n557, us01_n558, us01_n559, us01_n560, us01_n561, us01_n562, us01_n563, 
       us01_n564, us01_n565, us01_n566, us01_n567, us01_n568, us01_n569, us01_n570, us01_n571, us01_n572, 
       us01_n573, us01_n574, us01_n575, us01_n576, us01_n577, us01_n578, us01_n579, us01_n580, us01_n581, 
       us01_n582, us01_n583, us01_n584, us01_n585, us01_n586, us01_n587, us01_n588, us01_n589, us01_n590, 
       us01_n591, us01_n592, us01_n593, us01_n594, us01_n595, us01_n596, us01_n597, us01_n598, us01_n599, 
       us01_n600, us01_n601, us01_n602, us01_n603, us01_n604, us01_n605, us01_n606, us01_n607, us01_n608, 
       us01_n609, us01_n610, us01_n611, us01_n612, us01_n613, us01_n614, us01_n615, us01_n616, us01_n617, 
       us01_n618, us01_n619, us01_n620, us01_n621, us01_n622, us01_n623, us01_n624, us01_n625, us01_n626, 
       us01_n627, us01_n628, us01_n629, us01_n630, us01_n631, us01_n632, us01_n633, us01_n634, us01_n635, 
       us01_n636, us01_n637, us01_n638, us01_n639, us01_n640, us01_n641, us01_n642, us01_n643, us01_n644, 
       us01_n645, us01_n646, us01_n647, us01_n648, us01_n649, us01_n650, us01_n651, us01_n652, us01_n653, 
       us01_n654, us01_n655, us01_n656, us01_n657, us01_n658, us01_n659, us01_n660, us01_n661, us01_n662, 
       us01_n663, us01_n664, us01_n665, us01_n666, us01_n667, us01_n668, us01_n669, us01_n670, us01_n671, 
       us01_n672, us01_n673, us01_n674, us01_n675, us01_n676, us01_n677, us01_n678, us01_n679, us01_n680, 
       us01_n681, us01_n682, us01_n683, us01_n684, us01_n685, us01_n686, us01_n687, us01_n688, us01_n689, 
       us01_n690, us01_n691, us01_n692, us01_n693, us01_n694, us01_n695, us01_n696, us01_n697, us01_n698, 
       us01_n699, us01_n700, us01_n701, us01_n702, us01_n703, us01_n704, us01_n705, us01_n706, us01_n707, 
       us01_n708, us01_n709, us01_n710, us01_n711, us01_n712, us01_n713, us01_n714, us01_n715, us01_n716, 
       us01_n717, us01_n718, us01_n719, us01_n720, us01_n721, us01_n722, us01_n723, us01_n724, us01_n725, 
       us01_n726, us01_n727, us01_n728, us01_n729, us01_n730, us01_n731, us01_n732, us01_n733, us01_n734, 
       us01_n735, us01_n736, us01_n737, us01_n738, us01_n739, us01_n740, us01_n741, us01_n742, us01_n743, 
       us01_n744, us01_n745, us01_n746, us01_n747, us01_n748, us01_n749, us01_n750, us01_n751, us01_n752, 
       us01_n753, us01_n754, us01_n755, us01_n756, us01_n757, us01_n758, us01_n759, us01_n760, us01_n761, 
       us01_n762, us01_n763, us01_n764, us01_n765, us01_n766, us01_n767, us01_n768, us01_n769, us01_n770, 
       us01_n771, us01_n772, us01_n773, us01_n774, us01_n775, us01_n776, us01_n777, us01_n778, us01_n779, 
       us01_n780, us01_n781, us01_n782, us01_n783, us01_n784, us01_n785, us01_n786, us01_n787, us01_n788, 
       us01_n789, us01_n790, us01_n791, us01_n792, us01_n793, us01_n794, us01_n795, us01_n796, us01_n797, 
       us01_n798, us01_n799, us01_n800, us01_n801, us01_n802, us01_n803, us01_n804, us01_n805, us01_n806, 
       us01_n807, us01_n808, us01_n809, us01_n810, us01_n811, us01_n812, us01_n813, us01_n814, us01_n815, 
       us01_n816, us01_n817, us01_n818, us01_n819, us01_n820, us01_n821, us01_n822, us01_n823, us01_n824, 
       us01_n825, us01_n826, us01_n827, us01_n828, us01_n829, us01_n830, us01_n831, us01_n832, us01_n833, 
       us01_n834, us01_n835, us01_n836, us01_n837, us01_n838, us01_n839, us01_n840, us01_n841, us01_n842, 
       us01_n843, us01_n844, us01_n845, us01_n846, us01_n847, us01_n848, us01_n849, us01_n850, us01_n851, 
       us01_n852, us01_n853, us01_n854, us01_n855, us01_n856, us01_n857, us01_n858, us01_n859, us01_n860, 
       us01_n861, us01_n862, us01_n863, us01_n864, us01_n865, us01_n866, us01_n867, us01_n868, us01_n869, 
       us01_n870, us01_n871, us01_n872, us01_n873, us01_n874, us20_n438, us20_n439, us20_n440, us20_n441, 
       us20_n442, us20_n443, us20_n444, us20_n445, us20_n446, us20_n447, us20_n448, us20_n449, us20_n450, 
       us20_n451, us20_n452, us20_n453, us20_n454, us20_n455, us20_n456, us20_n457, us20_n458, us20_n459, 
       us20_n460, us20_n461, us20_n462, us20_n463, us20_n464, us20_n465, us20_n466, us20_n467, us20_n468, 
       us20_n469, us20_n470, us20_n471, us20_n472, us20_n473, us20_n474, us20_n475, us20_n476, us20_n477, 
       us20_n478, us20_n479, us20_n480, us20_n481, us20_n482, us20_n483, us20_n484, us20_n485, us20_n486, 
       us20_n487, us20_n488, us20_n489, us20_n490, us20_n491, us20_n492, us20_n493, us20_n494, us20_n495, 
       us20_n496, us20_n497, us20_n498, us20_n499, us20_n500, us20_n501, us20_n502, us20_n503, us20_n504, 
       us20_n505, us20_n506, us20_n507, us20_n508, us20_n509, us20_n510, us20_n511, us20_n512, us20_n513, 
       us20_n514, us20_n515, us20_n516, us20_n517, us20_n518, us20_n519, us20_n520, us20_n521, us20_n522, 
       us20_n523, us20_n524, us20_n525, us20_n526, us20_n527, us20_n528, us20_n529, us20_n530, us20_n531, 
       us20_n532, us20_n533, us20_n534, us20_n535, us20_n536, us20_n537, us20_n538, us20_n539, us20_n540, 
       us20_n541, us20_n542, us20_n543, us20_n544, us20_n545, us20_n546, us20_n547, us20_n548, us20_n549, 
       us20_n550, us20_n551, us20_n552, us20_n553, us20_n554, us20_n555, us20_n556, us20_n557, us20_n558, 
       us20_n559, us20_n560, us20_n561, us20_n562, us20_n563, us20_n564, us20_n565, us20_n566, us20_n567, 
       us20_n568, us20_n569, us20_n570, us20_n571, us20_n572, us20_n573, us20_n574, us20_n575, us20_n576, 
       us20_n577, us20_n578, us20_n579, us20_n580, us20_n581, us20_n582, us20_n583, us20_n584, us20_n585, 
       us20_n586, us20_n587, us20_n588, us20_n589, us20_n590, us20_n591, us20_n592, us20_n593, us20_n594, 
       us20_n595, us20_n596, us20_n597, us20_n598, us20_n599, us20_n600, us20_n601, us20_n602, us20_n603, 
       us20_n604, us20_n605, us20_n606, us20_n607, us20_n608, us20_n609, us20_n610, us20_n611, us20_n612, 
       us20_n613, us20_n614, us20_n615, us20_n616, us20_n617, us20_n618, us20_n619, us20_n620, us20_n621, 
       us20_n622, us20_n623, us20_n624, us20_n625, us20_n626, us20_n627, us20_n628, us20_n629, us20_n630, 
       us20_n631, us20_n632, us20_n633, us20_n634, us20_n635, us20_n636, us20_n637, us20_n638, us20_n639, 
       us20_n640, us20_n641, us20_n642, us20_n643, us20_n644, us20_n645, us20_n646, us20_n647, us20_n648, 
       us20_n649, us20_n650, us20_n651, us20_n652, us20_n653, us20_n654, us20_n655, us20_n656, us20_n657, 
       us20_n658, us20_n659, us20_n660, us20_n661, us20_n662, us20_n663, us20_n664, us20_n665, us20_n666, 
       us20_n667, us20_n668, us20_n669, us20_n670, us20_n671, us20_n672, us20_n673, us20_n674, us20_n675, 
       us20_n676, us20_n677, us20_n678, us20_n679, us20_n680, us20_n681, us20_n682, us20_n683, us20_n684, 
       us20_n685, us20_n686, us20_n687, us20_n688, us20_n689, us20_n690, us20_n691, us20_n692, us20_n693, 
       us20_n694, us20_n695, us20_n696, us20_n697, us20_n698, us20_n699, us20_n700, us20_n701, us20_n702, 
       us20_n703, us20_n704, us20_n705, us20_n706, us20_n707, us20_n708, us20_n709, us20_n710, us20_n711, 
       us20_n712, us20_n713, us20_n714, us20_n715, us20_n716, us20_n717, us20_n718, us20_n719, us20_n720, 
       us20_n721, us20_n722, us20_n723, us20_n724, us20_n725, us20_n726, us20_n727, us20_n728, us20_n729, 
       us20_n730, us20_n731, us20_n732, us20_n733, us20_n734, us20_n735, us20_n736, us20_n737, us20_n738, 
       us20_n739, us20_n740, us20_n741, us20_n742, us20_n743, us20_n744, us20_n745, us20_n746, us20_n747, 
       us20_n748, us20_n749, us20_n750, us20_n751, us20_n752, us20_n753, us20_n754, us20_n755, us20_n756, 
       us20_n757, us20_n758, us20_n759, us20_n760, us20_n761, us20_n762, us20_n763, us20_n764, us20_n765, 
       us20_n766, us20_n767, us20_n768, us20_n769, us20_n770, us20_n771, us20_n772, us20_n773, us20_n774, 
       us20_n775, us20_n776, us20_n777, us20_n778, us20_n779, us20_n780, us20_n781, us20_n782, us20_n783, 
       us20_n784, us20_n785, us20_n786, us20_n787, us20_n788, us20_n789, us20_n790, us20_n791, us20_n792, 
       us20_n793, us20_n794, us20_n795, us20_n796, us20_n797, us20_n798, us20_n799, us20_n800, us20_n801, 
       us20_n802, us20_n803, us20_n804, us20_n805, us20_n806, us20_n807, us20_n808, us20_n809, us20_n810, 
       us20_n811, us20_n812, us20_n813, us20_n814, us20_n815, us20_n816, us20_n817, us20_n818, us20_n819, 
       us20_n820, us20_n821, us20_n822, us20_n823, us20_n824, us20_n825, us20_n826, us20_n827, us20_n828, 
       us20_n829, us20_n830, us20_n831, us20_n832, us20_n833, us20_n834, us20_n835, us20_n836, us20_n837, 
       us20_n838, us20_n839, us20_n840, us20_n841, us20_n842, us20_n843, us20_n844, us20_n845, us20_n846, 
       us20_n847, us20_n848, us20_n849, us20_n850, us20_n851, us20_n852, us20_n853, us20_n854, us20_n855, 
       us20_n856, us20_n857, us20_n858, us20_n859, us20_n860, us20_n861, us20_n862, us20_n863, us20_n864, 
       us20_n865, us20_n866, us20_n867, us20_n868, us20_n869, us20_n870, us20_n871, us20_n872, us20_n873, 
       us20_n874, us20_n875, us20_n876, us32_n438, us32_n439, us32_n440, us32_n441, us32_n442, us32_n443, 
       us32_n444, us32_n445, us32_n446, us32_n447, us32_n448, us32_n449, us32_n450, us32_n451, us32_n452, 
       us32_n453, us32_n454, us32_n455, us32_n456, us32_n457, us32_n458, us32_n459, us32_n460, us32_n461, 
       us32_n462, us32_n463, us32_n464, us32_n465, us32_n466, us32_n467, us32_n468, us32_n469, us32_n470, 
       us32_n471, us32_n472, us32_n473, us32_n474, us32_n475, us32_n476, us32_n477, us32_n478, us32_n479, 
       us32_n480, us32_n481, us32_n482, us32_n483, us32_n484, us32_n485, us32_n486, us32_n487, us32_n488, 
       us32_n489, us32_n490, us32_n491, us32_n492, us32_n493, us32_n494, us32_n495, us32_n496, us32_n497, 
       us32_n498, us32_n499, us32_n500, us32_n501, us32_n502, us32_n503, us32_n504, us32_n505, us32_n506, 
       us32_n507, us32_n508, us32_n509, us32_n510, us32_n511, us32_n512, us32_n513, us32_n514, us32_n515, 
       us32_n516, us32_n517, us32_n518, us32_n519, us32_n520, us32_n521, us32_n522, us32_n523, us32_n524, 
       us32_n525, us32_n526, us32_n527, us32_n528, us32_n529, us32_n530, us32_n531, us32_n532, us32_n533, 
       us32_n534, us32_n535, us32_n536, us32_n537, us32_n538, us32_n539, us32_n540, us32_n541, us32_n542, 
       us32_n543, us32_n544, us32_n545, us32_n546, us32_n547, us32_n548, us32_n549, us32_n550, us32_n551, 
       us32_n552, us32_n553, us32_n554, us32_n555, us32_n556, us32_n557, us32_n558, us32_n559, us32_n560, 
       us32_n561, us32_n562, us32_n563, us32_n564, us32_n565, us32_n566, us32_n567, us32_n568, us32_n569, 
       us32_n570, us32_n571, us32_n572, us32_n573, us32_n574, us32_n575, us32_n576, us32_n577, us32_n578, 
       us32_n579, us32_n580, us32_n581, us32_n582, us32_n583, us32_n584, us32_n585, us32_n586, us32_n587, 
       us32_n588, us32_n589, us32_n590, us32_n591, us32_n592, us32_n593, us32_n594, us32_n595, us32_n596, 
       us32_n597, us32_n598, us32_n599, us32_n600, us32_n601, us32_n602, us32_n603, us32_n604, us32_n605, 
       us32_n606, us32_n607, us32_n608, us32_n609, us32_n610, us32_n611, us32_n612, us32_n613, us32_n614, 
       us32_n615, us32_n616, us32_n617, us32_n618, us32_n619, us32_n620, us32_n621, us32_n622, us32_n623, 
       us32_n624, us32_n625, us32_n626, us32_n627, us32_n628, us32_n629, us32_n630, us32_n631, us32_n632, 
       us32_n633, us32_n634, us32_n635, us32_n636, us32_n637, us32_n638, us32_n639, us32_n640, us32_n641, 
       us32_n642, us32_n643, us32_n644, us32_n645, us32_n646, us32_n647, us32_n648, us32_n649, us32_n650, 
       us32_n651, us32_n652, us32_n653, us32_n654, us32_n655, us32_n656, us32_n657, us32_n658, us32_n659, 
       us32_n660, us32_n661, us32_n662, us32_n663, us32_n664, us32_n665, us32_n666, us32_n667, us32_n668, 
       us32_n669, us32_n670, us32_n671, us32_n672, us32_n673, us32_n674, us32_n675, us32_n676, us32_n677, 
       us32_n678, us32_n679, us32_n680, us32_n681, us32_n682, us32_n683, us32_n684, us32_n685, us32_n686, 
       us32_n687, us32_n688, us32_n689, us32_n690, us32_n691, us32_n692, us32_n693, us32_n694, us32_n695, 
       us32_n696, us32_n697, us32_n698, us32_n699, us32_n700, us32_n701, us32_n702, us32_n703, us32_n704, 
       us32_n705, us32_n706, us32_n707, us32_n708, us32_n709, us32_n710, us32_n711, us32_n712, us32_n713, 
       us32_n714, us32_n715, us32_n716, us32_n717, us32_n718, us32_n719, us32_n720, us32_n721, us32_n722, 
       us32_n723, us32_n724, us32_n725, us32_n726, us32_n727, us32_n728, us32_n729, us32_n730, us32_n731, 
       us32_n732, us32_n733, us32_n734, us32_n735, us32_n736, us32_n737, us32_n738, us32_n739, us32_n740, 
       us32_n741, us32_n742, us32_n743, us32_n744, us32_n745, us32_n746, us32_n747, us32_n748, us32_n749, 
       us32_n750, us32_n751, us32_n752, us32_n753, us32_n754, us32_n755, us32_n756, us32_n757, us32_n758, 
       us32_n759, us32_n760, us32_n761, us32_n762, us32_n763, us32_n764, us32_n765, us32_n766, us32_n767, 
       us32_n768, us32_n769, us32_n770, us32_n771, us32_n772, us32_n773, us32_n774, us32_n775, us32_n776, 
       us32_n777, us32_n778, us32_n779, us32_n780, us32_n781, us32_n782, us32_n783, us32_n784, us32_n785, 
       us32_n786, us32_n787, us32_n788, us32_n789, us32_n790, us32_n791, us32_n792, us32_n793, us32_n794, 
       us32_n795, us32_n796, us32_n797, us32_n798, us32_n799, us32_n800, us32_n801, us32_n802, us32_n803, 
       us32_n804, us32_n805, us32_n806, us32_n807, us32_n808, us32_n809, us32_n810, us32_n811, us32_n812, 
       us32_n813, us32_n814, us32_n815, us32_n816, us32_n817, us32_n818, us32_n819, us32_n820, us32_n821, 
       us32_n822, us32_n823, us32_n824, us32_n825, us32_n826, us32_n827, us32_n828, us32_n829, us32_n830, 
       us32_n831, us32_n832, us32_n833, us32_n834, us32_n835, us32_n836, us32_n837, us32_n838, us32_n839, 
       us32_n840, us32_n841, us32_n842, us32_n843, us32_n844, us32_n845, us32_n846, us32_n847, us32_n848, 
       us32_n849, us32_n850, us32_n851, us32_n852, us32_n853, us32_n854, us32_n855, us32_n856, us32_n857, 
       us32_n858, us32_n859, us32_n860, us32_n861, us32_n862, us32_n863, us32_n864, us32_n865, us32_n866, 
       us32_n867, us32_n868, us32_n869, us32_n870, us32_n871, us32_n872, us32_n873, us32_n874, us32_n875, 
        us32_n876;
  NOR2_X1 us01_U10 (.ZN( us01_n573 ) , .A1( us01_n620 ) , .A2( us01_n743 ) );
  AOI211_X1 us01_U100 (.B( us01_n537 ) , .A( us01_n538 ) , .ZN( us01_n549 ) , .C2( us01_n837 ) , .C1( us01_n849 ) );
  NOR4_X1 us01_U101 (.A4( us01_n542 ) , .A3( us01_n543 ) , .A2( us01_n544 ) , .A1( us01_n545 ) , .ZN( us01_n546 ) );
  NOR4_X1 us01_U102 (.A4( us01_n607 ) , .A3( us01_n608 ) , .A2( us01_n609 ) , .A1( us01_n610 ) , .ZN( us01_n617 ) );
  NOR4_X1 us01_U103 (.ZN( us01_n618 ) , .A1( us01_n654 ) , .A3( us01_n664 ) , .A4( us01_n680 ) , .A2( us01_n764 ) );
  NOR4_X1 us01_U104 (.A4( us01_n612 ) , .A3( us01_n613 ) , .A2( us01_n614 ) , .A1( us01_n615 ) , .ZN( us01_n616 ) );
  NOR2_X1 us01_U105 (.ZN( us01_n684 ) , .A1( us01_n829 ) , .A2( us01_n830 ) );
  NAND4_X1 us01_U106 (.A4( us01_n471 ) , .A3( us01_n472 ) , .A2( us01_n473 ) , .A1( us01_n474 ) , .ZN( us01_n676 ) );
  NOR4_X1 us01_U107 (.A4( us01_n468 ) , .ZN( us01_n474 ) , .A3( us01_n554 ) , .A1( us01_n733 ) , .A2( us01_n753 ) );
  NOR4_X1 us01_U108 (.ZN( us01_n473 ) , .A1( us01_n529 ) , .A3( us01_n566 ) , .A4( us01_n598 ) , .A2( us01_n640 ) );
  NOR4_X1 us01_U109 (.ZN( us01_n472 ) , .A1( us01_n504 ) , .A3( us01_n542 ) , .A2( us01_n581 ) , .A4( us01_n714 ) );
  NOR2_X1 us01_U11 (.ZN( us01_n493 ) , .A1( us01_n676 ) , .A2( us01_n692 ) );
  NAND4_X1 us01_U110 (.A4( us01_n689 ) , .A3( us01_n690 ) , .A1( us01_n691 ) , .ZN( us01_n774 ) , .A2( us01_n870 ) );
  INV_X1 us01_U111 (.A( us01_n677 ) , .ZN( us01_n870 ) );
  AOI221_X1 us01_U112 (.A( us01_n679 ) , .ZN( us01_n690 ) , .B2( us01_n838 ) , .C1( us01_n840 ) , .C2( us01_n860 ) , .B1( us01_n863 ) );
  NOR4_X1 us01_U113 (.A4( us01_n685 ) , .A3( us01_n686 ) , .A2( us01_n687 ) , .A1( us01_n688 ) , .ZN( us01_n689 ) );
  NOR2_X1 us01_U114 (.ZN( us01_n731 ) , .A2( us01_n830 ) , .A1( us01_n843 ) );
  NAND4_X1 us01_U115 (.A4( us01_n717 ) , .A3( us01_n718 ) , .A2( us01_n719 ) , .ZN( us01_n739 ) , .A1( us01_n855 ) );
  AOI221_X1 us01_U116 (.A( us01_n708 ) , .ZN( us01_n719 ) , .C2( us01_n842 ) , .B2( us01_n843 ) , .C1( us01_n859 ) , .B1( us01_n860 ) );
  INV_X1 us01_U117 (.A( us01_n707 ) , .ZN( us01_n855 ) );
  NOR4_X1 us01_U118 (.A4( us01_n713 ) , .A3( us01_n714 ) , .A2( us01_n715 ) , .A1( us01_n716 ) , .ZN( us01_n717 ) );
  NOR2_X1 us01_U119 (.ZN( us01_n645 ) , .A1( us01_n852 ) , .A2( us01_n866 ) );
  NOR2_X1 us01_U12 (.A1( us01_n676 ) , .ZN( us01_n691 ) , .A2( us01_n805 ) );
  NAND4_X1 us01_U120 (.A4( us01_n571 ) , .A3( us01_n572 ) , .A1( us01_n573 ) , .ZN( us01_n721 ) , .A2( us01_n872 ) );
  AOI221_X1 us01_U121 (.A( us01_n562 ) , .C2( us01_n563 ) , .ZN( us01_n572 ) , .B2( us01_n843 ) , .B1( us01_n850 ) , .C1( us01_n851 ) );
  NOR4_X1 us01_U122 (.A4( us01_n567 ) , .A3( us01_n568 ) , .A2( us01_n569 ) , .A1( us01_n570 ) , .ZN( us01_n571 ) );
  INV_X1 us01_U123 (.A( us01_n605 ) , .ZN( us01_n872 ) );
  NAND4_X1 us01_U124 (.A4( us01_n491 ) , .A3( us01_n492 ) , .A1( us01_n493 ) , .ZN( us01_n800 ) , .A2( us01_n865 ) );
  AOI221_X1 us01_U125 (.A( us01_n487 ) , .ZN( us01_n492 ) , .B2( us01_n834 ) , .C2( us01_n839 ) , .C1( us01_n849 ) , .B1( us01_n858 ) );
  INV_X1 us01_U126 (.A( us01_n776 ) , .ZN( us01_n865 ) );
  NOR4_X1 us01_U127 (.A2( us01_n489 ) , .A1( us01_n490 ) , .ZN( us01_n491 ) , .A3( us01_n578 ) , .A4( us01_n610 ) );
  NOR4_X1 us01_U128 (.A3( us01_n753 ) , .A2( us01_n754 ) , .A1( us01_n755 ) , .ZN( us01_n756 ) , .A4( us01_n867 ) );
  AOI211_X1 us01_U129 (.B( us01_n743 ) , .A( us01_n744 ) , .ZN( us01_n757 ) , .C1( us01_n830 ) , .C2( us01_n851 ) );
  NOR3_X1 us01_U13 (.ZN( us01_n502 ) , .A2( us01_n677 ) , .A3( us01_n775 ) , .A1( us01_n874 ) );
  NOR3_X1 us01_U130 (.A3( us01_n739 ) , .A2( us01_n740 ) , .A1( us01_n741 ) , .ZN( us01_n758 ) );
  NOR4_X1 us01_U131 (.A4( us01_n732 ) , .A3( us01_n733 ) , .A2( us01_n734 ) , .A1( us01_n735 ) , .ZN( us01_n736 ) );
  AOI211_X1 us01_U132 (.B( us01_n723 ) , .A( us01_n724 ) , .ZN( us01_n737 ) , .C1( us01_n841 ) , .C2( us01_n853 ) );
  NOR3_X1 us01_U133 (.A3( us01_n720 ) , .A1( us01_n721 ) , .ZN( us01_n738 ) , .A2( us01_n739 ) );
  INV_X1 us01_U134 (.A( us01_n760 ) , .ZN( us01_n828 ) );
  NAND4_X1 us01_U135 (.ZN( sa01_sr_3 ) , .A4( us01_n702 ) , .A3( us01_n703 ) , .A2( us01_n704 ) , .A1( us01_n705 ) );
  NOR4_X1 us01_U136 (.A4( us01_n698 ) , .A3( us01_n699 ) , .A2( us01_n700 ) , .A1( us01_n701 ) , .ZN( us01_n702 ) );
  AOI211_X1 us01_U137 (.B( us01_n692 ) , .A( us01_n693 ) , .ZN( us01_n703 ) , .C2( us01_n829 ) , .C1( us01_n849 ) );
  NOR2_X1 us01_U138 (.ZN( us01_n705 ) , .A2( us01_n774 ) , .A1( us01_n798 ) );
  OR4_X1 us01_U139 (.A4( us01_n680 ) , .A3( us01_n681 ) , .A2( us01_n682 ) , .A1( us01_n683 ) , .ZN( us01_n688 ) );
  INV_X1 us01_U14 (.A( us01_n704 ) , .ZN( us01_n874 ) );
  OR4_X1 us01_U140 (.ZN( us01_n464 ) , .A4( us01_n516 ) , .A3( us01_n527 ) , .A2( us01_n576 ) , .A1( us01_n710 ) );
  OR4_X1 us01_U141 (.A4( us01_n564 ) , .A3( us01_n565 ) , .A2( us01_n566 ) , .ZN( us01_n570 ) , .A1( us01_n663 ) );
  OR4_X1 us01_U142 (.A4( us01_n516 ) , .A2( us01_n517 ) , .A1( us01_n518 ) , .ZN( us01_n520 ) , .A3( us01_n819 ) );
  OR4_X1 us01_U143 (.ZN( us01_n490 ) , .A4( us01_n532 ) , .A2( us01_n545 ) , .A1( us01_n557 ) , .A3( us01_n630 ) );
  OR4_X1 us01_U144 (.A4( us01_n578 ) , .A3( us01_n579 ) , .A2( us01_n580 ) , .A1( us01_n581 ) , .ZN( us01_n582 ) );
  INV_X1 us01_U145 (.A( us01_n695 ) , .ZN( us01_n836 ) );
  NAND2_X1 us01_U146 (.ZN( us01_n611 ) , .A2( us01_n835 ) , .A1( us01_n871 ) );
  OR3_X1 us01_U147 (.A3( us01_n504 ) , .A2( us01_n505 ) , .A1( us01_n506 ) , .ZN( us01_n509 ) );
  AOI221_X1 us01_U148 (.A( us01_n711 ) , .B2( us01_n712 ) , .ZN( us01_n718 ) , .C1( us01_n830 ) , .B1( us01_n837 ) , .C2( us01_n861 ) );
  OR2_X1 us01_U149 (.A2( us01_n709 ) , .A1( us01_n710 ) , .ZN( us01_n711 ) );
  INV_X1 us01_U15 (.A( us01_n678 ) , .ZN( us01_n838 ) );
  INV_X1 us01_U150 (.A( us01_n461 ) , .ZN( us01_n862 ) );
  OAI21_X1 us01_U151 (.ZN( us01_n461 ) , .B1( us01_n807 ) , .A( us01_n832 ) , .B2( us01_n849 ) );
  INV_X1 us01_U152 (.A( us01_n752 ) , .ZN( us01_n867 ) );
  OAI21_X1 us01_U153 (.B1( us01_n751 ) , .ZN( us01_n752 ) , .A( us01_n843 ) , .B2( us01_n866 ) );
  INV_X1 us01_U154 (.A( us01_n670 ) , .ZN( us01_n857 ) );
  AOI21_X1 us01_U155 (.A( us01_n668 ) , .B1( us01_n669 ) , .ZN( us01_n670 ) , .B2( us01_n854 ) );
  AOI222_X1 us01_U156 (.ZN( us01_n658 ) , .A2( us01_n837 ) , .B1( us01_n839 ) , .C2( us01_n843 ) , .A1( us01_n858 ) , .C1( us01_n861 ) , .B2( us01_n868 ) );
  INV_X1 us01_U157 (.A( us01_n645 ) , .ZN( us01_n868 ) );
  OAI22_X1 us01_U158 (.ZN( us01_n481 ) , .A1( us01_n706 ) , .B2( us01_n783 ) , .A2( us01_n804 ) , .B1( us01_n810 ) );
  OAI22_X1 us01_U159 (.ZN( us01_n635 ) , .A1( us01_n697 ) , .B2( us01_n726 ) , .A2( us01_n760 ) , .B1( us01_n814 ) );
  NOR4_X1 us01_U16 (.A4( us01_n443 ) , .A3( us01_n444 ) , .A2( us01_n514 ) , .A1( us01_n539 ) , .ZN( us01_n704 ) );
  OAI222_X1 us01_U160 (.ZN( us01_n503 ) , .C2( us01_n623 ) , .B2( us01_n645 ) , .B1( us01_n745 ) , .A2( us01_n746 ) , .C1( us01_n803 ) , .A1( us01_n804 ) );
  OAI222_X1 us01_U161 (.B2( us01_n745 ) , .B1( us01_n746 ) , .A2( us01_n747 ) , .ZN( us01_n755 ) , .C2( us01_n803 ) , .C1( us01_n812 ) , .A1( us01_n815 ) );
  OAI222_X1 us01_U162 (.B2( us01_n706 ) , .ZN( us01_n707 ) , .C2( us01_n722 ) , .B1( us01_n745 ) , .A1( us01_n804 ) , .C1( us01_n812 ) , .A2( us01_n813 ) );
  AOI22_X1 us01_U163 (.ZN( us01_n694 ) , .A1( us01_n828 ) , .B2( us01_n841 ) , .A2( us01_n863 ) , .B1( us01_n866 ) );
  AOI22_X1 us01_U164 (.A2( us01_n780 ) , .ZN( us01_n781 ) , .B2( us01_n829 ) , .A1( us01_n832 ) , .B1( us01_n861 ) );
  INV_X1 us01_U165 (.A( us01_n728 ) , .ZN( us01_n837 ) );
  AOI221_X1 us01_U166 (.A( us01_n762 ) , .ZN( us01_n772 ) , .C2( us01_n808 ) , .B2( us01_n833 ) , .C1( us01_n853 ) , .B1( us01_n864 ) );
  AOI21_X1 us01_U167 (.B2( us01_n761 ) , .ZN( us01_n762 ) , .A( us01_n786 ) , .B1( us01_n790 ) );
  INV_X1 us01_U168 (.A( us01_n759 ) , .ZN( us01_n833 ) );
  INV_X1 us01_U169 (.A( us01_n788 ) , .ZN( us01_n830 ) );
  OR3_X1 us01_U17 (.ZN( us01_n444 ) , .A1( us01_n526 ) , .A3( us01_n575 ) , .A2( us01_n873 ) );
  OAI221_X1 us01_U170 (.A( us01_n725 ) , .C2( us01_n726 ) , .B2( us01_n727 ) , .B1( us01_n728 ) , .ZN( us01_n735 ) , .C1( us01_n815 ) );
  AOI22_X1 us01_U171 (.ZN( us01_n725 ) , .B1( us01_n830 ) , .A2( us01_n836 ) , .A1( us01_n861 ) , .B2( us01_n864 ) );
  NAND2_X1 us01_U172 (.A1( us01_n449 ) , .A2( us01_n451 ) , .ZN( us01_n760 ) );
  OAI22_X1 us01_U173 (.ZN( us01_n622 ) , .B1( us01_n667 ) , .B2( us01_n745 ) , .A1( us01_n813 ) , .A2( us01_n814 ) );
  OAI22_X1 us01_U174 (.A1( us01_n722 ) , .ZN( us01_n724 ) , .B2( us01_n748 ) , .B1( us01_n810 ) , .A2( us01_n814 ) );
  OAI22_X1 us01_U175 (.ZN( us01_n487 ) , .A1( us01_n722 ) , .B2( us01_n726 ) , .B1( us01_n728 ) , .A2( us01_n777 ) );
  OAI22_X1 us01_U176 (.B2( us01_n777 ) , .B1( us01_n778 ) , .ZN( us01_n779 ) , .A2( us01_n812 ) , .A1( us01_n813 ) );
  OAI22_X1 us01_U177 (.B2( us01_n748 ) , .B1( us01_n749 ) , .A1( us01_n750 ) , .ZN( us01_n754 ) , .A2( us01_n804 ) );
  NOR3_X1 us01_U178 (.ZN( us01_n750 ) , .A2( us01_n851 ) , .A1( us01_n861 ) , .A3( us01_n863 ) );
  NOR2_X1 us01_U179 (.ZN( us01_n749 ) , .A2( us01_n850 ) , .A1( us01_n858 ) );
  OR4_X1 us01_U18 (.A4( us01_n440 ) , .A2( us01_n441 ) , .A1( us01_n442 ) , .ZN( us01_n443 ) , .A3( us01_n551 ) );
  INV_X1 us01_U180 (.A( us01_n803 ) , .ZN( us01_n858 ) );
  OAI22_X1 us01_U181 (.B2( us01_n742 ) , .ZN( us01_n744 ) , .A2( us01_n760 ) , .B1( us01_n778 ) , .A1( us01_n790 ) );
  OAI22_X1 us01_U182 (.ZN( us01_n494 ) , .A2( us01_n742 ) , .A1( us01_n778 ) , .B1( us01_n789 ) , .B2( us01_n804 ) );
  OAI22_X1 us01_U183 (.B2( us01_n801 ) , .B1( us01_n802 ) , .A2( us01_n803 ) , .A1( us01_n804 ) , .ZN( us01_n806 ) );
  OAI22_X1 us01_U184 (.ZN( us01_n693 ) , .A2( us01_n728 ) , .A1( us01_n778 ) , .B1( us01_n789 ) , .B2( us01_n815 ) );
  NOR2_X1 us01_U185 (.ZN( us01_n713 ) , .A1( us01_n803 ) , .A2( us01_n815 ) );
  NOR2_X1 us01_U186 (.A1( us01_n697 ) , .ZN( us01_n766 ) , .A2( us01_n811 ) );
  INV_X1 us01_U187 (.A( us01_n786 ) , .ZN( us01_n843 ) );
  NOR2_X1 us01_U188 (.ZN( us01_n539 ) , .A2( us01_n695 ) , .A1( us01_n697 ) );
  INV_X1 us01_U189 (.A( us01_n742 ) , .ZN( us01_n835 ) );
  INV_X1 us01_U19 (.A( us01_n611 ) , .ZN( us01_n873 ) );
  INV_X1 us01_U190 (.A( us01_n814 ) , .ZN( us01_n829 ) );
  INV_X1 us01_U191 (.A( us01_n812 ) , .ZN( us01_n831 ) );
  OAI22_X1 us01_U192 (.B1( us01_n488 ) , .ZN( us01_n489 ) , .A1( us01_n684 ) , .A2( us01_n761 ) , .B2( us01_n815 ) );
  NOR3_X1 us01_U193 (.ZN( us01_n488 ) , .A1( us01_n780 ) , .A2( us01_n848 ) , .A3( us01_n861 ) );
  NOR2_X1 us01_U194 (.A2( us01_n742 ) , .ZN( us01_n753 ) , .A1( us01_n803 ) );
  NOR2_X1 us01_U195 (.ZN( us01_n733 ) , .A2( us01_n801 ) , .A1( us01_n803 ) );
  INV_X1 us01_U196 (.A( us01_n790 ) , .ZN( us01_n849 ) );
  NOR2_X1 us01_U197 (.A2( us01_n742 ) , .ZN( us01_n767 ) , .A1( us01_n810 ) );
  NOR2_X1 us01_U198 (.ZN( us01_n664 ) , .A1( us01_n726 ) , .A2( us01_n801 ) );
  OAI22_X1 us01_U199 (.ZN( us01_n708 ) , .A2( us01_n726 ) , .B2( us01_n727 ) , .A1( us01_n742 ) , .B1( us01_n811 ) );
  AOI222_X1 us01_U20 (.ZN( us01_n561 ) , .B1( us01_n828 ) , .C1( us01_n839 ) , .A2( us01_n841 ) , .A1( us01_n852 ) , .B2( us01_n861 ) , .C2( us01_n871 ) );
  NOR2_X1 us01_U200 (.ZN( us01_n650 ) , .A1( us01_n667 ) , .A2( us01_n812 ) );
  NOR2_X1 us01_U201 (.ZN( us01_n592 ) , .A2( us01_n695 ) , .A1( us01_n726 ) );
  NOR2_X1 us01_U202 (.A1( us01_n667 ) , .ZN( us01_n671 ) , .A2( us01_n742 ) );
  NOR2_X1 us01_U203 (.ZN( us01_n600 ) , .A1( us01_n667 ) , .A2( us01_n801 ) );
  NOR2_X1 us01_U204 (.A1( us01_n667 ) , .ZN( us01_n686 ) , .A2( us01_n814 ) );
  NOR2_X1 us01_U205 (.ZN( us01_n568 ) , .A1( us01_n726 ) , .A2( us01_n804 ) );
  NOR2_X1 us01_U206 (.A1( us01_n667 ) , .ZN( us01_n764 ) , .A2( us01_n811 ) );
  NOR2_X1 us01_U207 (.ZN( us01_n525 ) , .A1( us01_n667 ) , .A2( us01_n777 ) );
  NOR2_X1 us01_U208 (.ZN( us01_n652 ) , .A1( us01_n726 ) , .A2( us01_n811 ) );
  NOR2_X1 us01_U209 (.ZN( us01_n505 ) , .A1( us01_n810 ) , .A2( us01_n815 ) );
  NOR4_X1 us01_U21 (.ZN( us01_n471 ) , .A2( us01_n519 ) , .A4( us01_n592 ) , .A1( us01_n607 ) , .A3( us01_n627 ) );
  NOR2_X1 us01_U210 (.ZN( us01_n659 ) , .A1( us01_n727 ) , .A2( us01_n788 ) );
  NOR2_X1 us01_U211 (.ZN( us01_n544 ) , .A2( us01_n778 ) , .A1( us01_n812 ) );
  NOR2_X1 us01_U212 (.ZN( us01_n575 ) , .A2( us01_n697 ) , .A1( us01_n812 ) );
  NOR2_X1 us01_U213 (.ZN( us01_n507 ) , .A1( us01_n727 ) , .A2( us01_n777 ) );
  NOR2_X1 us01_U214 (.ZN( us01_n716 ) , .A2( us01_n722 ) , .A1( us01_n742 ) );
  INV_X1 us01_U215 (.A( us01_n748 ) , .ZN( us01_n840 ) );
  NOR2_X1 us01_U216 (.ZN( us01_n530 ) , .A2( us01_n747 ) , .A1( us01_n748 ) );
  NOR2_X1 us01_U217 (.ZN( us01_n660 ) , .A2( us01_n695 ) , .A1( us01_n727 ) );
  NOR2_X1 us01_U218 (.ZN( us01_n613 ) , .A1( us01_n783 ) , .A2( us01_n813 ) );
  NOR2_X1 us01_U219 (.ZN( us01_n627 ) , .A2( us01_n726 ) , .A1( us01_n783 ) );
  NOR4_X1 us01_U22 (.ZN( us01_n477 ) , .A1( us01_n518 ) , .A4( us01_n555 ) , .A3( us01_n580 ) , .A2( us01_n628 ) );
  NOR2_X1 us01_U220 (.ZN( us01_n609 ) , .A2( us01_n778 ) , .A1( us01_n804 ) );
  NOR2_X1 us01_U221 (.ZN( us01_n661 ) , .A1( us01_n727 ) , .A2( us01_n783 ) );
  NOR2_X1 us01_U222 (.ZN( us01_n626 ) , .A2( us01_n667 ) , .A1( us01_n783 ) );
  NOR2_X1 us01_U223 (.ZN( us01_n599 ) , .A2( us01_n778 ) , .A1( us01_n801 ) );
  INV_X1 us01_U224 (.A( us01_n745 ) , .ZN( us01_n832 ) );
  NOR2_X1 us01_U225 (.ZN( us01_n554 ) , .A1( us01_n760 ) , .A2( us01_n803 ) );
  NOR2_X1 us01_U226 (.ZN( us01_n529 ) , .A2( us01_n778 ) , .A1( us01_n814 ) );
  NOR2_X1 us01_U227 (.ZN( us01_n526 ) , .A2( us01_n722 ) , .A1( us01_n801 ) );
  NOR2_X1 us01_U228 (.A2( us01_n706 ) , .A1( us01_n748 ) , .ZN( us01_n769 ) );
  NOR2_X1 us01_U229 (.ZN( us01_n597 ) , .A2( us01_n789 ) , .A1( us01_n814 ) );
  NOR4_X1 us01_U23 (.ZN( us01_n454 ) , .A2( us01_n515 ) , .A1( us01_n541 ) , .A3( us01_n577 ) , .A4( us01_n613 ) );
  NOR2_X1 us01_U230 (.ZN( us01_n555 ) , .A1( us01_n790 ) , .A2( us01_n812 ) );
  NOR2_X1 us01_U231 (.ZN( us01_n542 ) , .A2( us01_n783 ) , .A1( us01_n790 ) );
  NOR2_X1 us01_U232 (.A2( us01_n695 ) , .ZN( us01_n714 ) , .A1( us01_n790 ) );
  NOR2_X1 us01_U233 (.ZN( us01_n665 ) , .A1( us01_n748 ) , .A2( us01_n813 ) );
  NOR2_X1 us01_U234 (.ZN( us01_n543 ) , .A1( us01_n747 ) , .A2( us01_n812 ) );
  NOR2_X1 us01_U235 (.ZN( us01_n553 ) , .A1( us01_n748 ) , .A2( us01_n789 ) );
  NOR2_X1 us01_U236 (.ZN( us01_n506 ) , .A2( us01_n778 ) , .A1( us01_n783 ) );
  NOR2_X1 us01_U237 (.ZN( us01_n541 ) , .A2( us01_n706 ) , .A1( us01_n783 ) );
  NOR2_X1 us01_U238 (.ZN( us01_n514 ) , .A1( us01_n706 ) , .A2( us01_n742 ) );
  NOR2_X1 us01_U239 (.ZN( us01_n662 ) , .A1( us01_n783 ) , .A2( us01_n789 ) );
  NOR4_X1 us01_U24 (.A4( us01_n530 ) , .A3( us01_n531 ) , .A2( us01_n532 ) , .ZN( us01_n533 ) , .A1( us01_n818 ) );
  NOR2_X1 us01_U240 (.ZN( us01_n556 ) , .A1( us01_n706 ) , .A2( us01_n814 ) );
  NOR2_X1 us01_U241 (.ZN( us01_n515 ) , .A1( us01_n706 ) , .A2( us01_n801 ) );
  NOR2_X1 us01_U242 (.ZN( us01_n612 ) , .A1( us01_n760 ) , .A2( us01_n810 ) );
  NOR2_X1 us01_U243 (.ZN( us01_n629 ) , .A1( us01_n722 ) , .A2( us01_n811 ) );
  NOR2_X1 us01_U244 (.A1( us01_n747 ) , .ZN( us01_n765 ) , .A2( us01_n801 ) );
  NOR2_X1 us01_U245 (.ZN( us01_n528 ) , .A2( us01_n742 ) , .A1( us01_n790 ) );
  INV_X1 us01_U246 (.A( us01_n804 ) , .ZN( us01_n839 ) );
  OAI22_X1 us01_U247 (.B1( us01_n438 ) , .ZN( us01_n442 ) , .A2( us01_n726 ) , .A1( us01_n742 ) , .B2( us01_n747 ) );
  NOR3_X1 us01_U248 (.ZN( us01_n438 ) , .A2( us01_n834 ) , .A3( us01_n835 ) , .A1( us01_n844 ) );
  INV_X1 us01_U249 (.A( us01_n726 ) , .ZN( us01_n850 ) );
  NOR4_X1 us01_U25 (.A4( us01_n539 ) , .A3( us01_n540 ) , .A2( us01_n541 ) , .ZN( us01_n548 ) , .A1( us01_n686 ) );
  NOR2_X1 us01_U250 (.ZN( us01_n519 ) , .A1( us01_n788 ) , .A2( us01_n810 ) );
  NOR2_X1 us01_U251 (.ZN( us01_n668 ) , .A1( us01_n788 ) , .A2( us01_n803 ) );
  AOI21_X1 us01_U252 (.ZN( us01_n550 ) , .B1( us01_n667 ) , .A( us01_n695 ) , .B2( us01_n803 ) );
  AOI21_X1 us01_U253 (.ZN( us01_n587 ) , .B2( us01_n697 ) , .B1( us01_n813 ) , .A( us01_n815 ) );
  NOR2_X1 us01_U254 (.ZN( us01_n504 ) , .A2( us01_n726 ) , .A1( us01_n760 ) );
  NOR2_X1 us01_U255 (.ZN( us01_n653 ) , .A1( us01_n788 ) , .A2( us01_n813 ) );
  INV_X1 us01_U256 (.A( us01_n801 ) , .ZN( us01_n841 ) );
  NOR2_X1 us01_U257 (.ZN( us01_n628 ) , .A1( us01_n745 ) , .A2( us01_n813 ) );
  NOR2_X1 us01_U258 (.ZN( us01_n545 ) , .A1( us01_n697 ) , .A2( us01_n742 ) );
  INV_X1 us01_U259 (.A( us01_n697 ) , .ZN( us01_n851 ) );
  NOR2_X1 us01_U26 (.ZN( us01_n678 ) , .A2( us01_n832 ) , .A1( us01_n837 ) );
  NOR2_X1 us01_U260 (.ZN( us01_n640 ) , .A2( us01_n786 ) , .A1( us01_n789 ) );
  AOI21_X1 us01_U261 (.ZN( us01_n648 ) , .A( us01_n777 ) , .B1( us01_n790 ) , .B2( us01_n803 ) );
  NOR2_X1 us01_U262 (.ZN( us01_n666 ) , .A2( us01_n706 ) , .A1( us01_n788 ) );
  NOR2_X1 us01_U263 (.A2( us01_n695 ) , .A1( us01_n778 ) , .ZN( us01_n818 ) );
  NOR2_X1 us01_U264 (.A1( us01_n695 ) , .ZN( us01_n768 ) , .A2( us01_n813 ) );
  AOI21_X1 us01_U265 (.ZN( us01_n624 ) , .B2( us01_n667 ) , .A( us01_n788 ) , .B1( us01_n789 ) );
  NOR2_X1 us01_U266 (.ZN( us01_n577 ) , .A2( us01_n706 ) , .A1( us01_n728 ) );
  INV_X1 us01_U267 (.A( us01_n761 ) , .ZN( us01_n864 ) );
  NOR2_X1 us01_U268 (.A2( us01_n706 ) , .A1( us01_n760 ) , .ZN( us01_n792 ) );
  NOR2_X1 us01_U269 (.ZN( us01_n607 ) , .A2( us01_n722 ) , .A1( us01_n815 ) );
  AOI222_X1 us01_U27 (.ZN( us01_n467 ) , .B1( us01_n830 ) , .A1( us01_n837 ) , .C1( us01_n840 ) , .C2( us01_n849 ) , .A2( us01_n853 ) , .B2( us01_n863 ) );
  NOR2_X1 us01_U270 (.ZN( us01_n531 ) , .A2( us01_n722 ) , .A1( us01_n728 ) );
  AOI21_X1 us01_U271 (.ZN( us01_n508 ) , .B2( us01_n667 ) , .A( us01_n728 ) , .B1( us01_n813 ) );
  AOI21_X1 us01_U272 (.ZN( us01_n537 ) , .B2( us01_n810 ) , .A( us01_n812 ) , .B1( us01_n813 ) );
  INV_X1 us01_U273 (.A( us01_n727 ) , .ZN( us01_n866 ) );
  NOR2_X1 us01_U274 (.ZN( us01_n540 ) , .A1( us01_n760 ) , .A2( us01_n789 ) );
  INV_X1 us01_U275 (.A( us01_n810 ) , .ZN( us01_n852 ) );
  AOI21_X1 us01_U276 (.B1( us01_n697 ) , .ZN( us01_n698 ) , .A( us01_n730 ) , .B2( us01_n761 ) );
  NOR2_X1 us01_U277 (.ZN( us01_n579 ) , .A1( us01_n667 ) , .A2( us01_n786 ) );
  AOI21_X1 us01_U278 (.ZN( us01_n589 ) , .B2( us01_n761 ) , .A( us01_n783 ) , .B1( us01_n810 ) );
  NOR2_X1 us01_U279 (.ZN( us01_n654 ) , .A1( us01_n745 ) , .A2( us01_n778 ) );
  NOR4_X1 us01_U28 (.A1( us01_n464 ) , .ZN( us01_n465 ) , .A4( us01_n540 ) , .A2( us01_n552 ) , .A3( us01_n612 ) );
  INV_X1 us01_U280 (.A( us01_n789 ) , .ZN( us01_n871 ) );
  AOI21_X1 us01_U281 (.B1( us01_n623 ) , .ZN( us01_n625 ) , .A( us01_n761 ) , .B2( us01_n812 ) );
  NOR2_X1 us01_U282 (.ZN( us01_n683 ) , .A1( us01_n727 ) , .A2( us01_n814 ) );
  AOI21_X1 us01_U283 (.A( us01_n813 ) , .B2( us01_n814 ) , .B1( us01_n815 ) , .ZN( us01_n816 ) );
  AOI21_X1 us01_U284 (.ZN( us01_n647 ) , .B1( us01_n727 ) , .B2( us01_n761 ) , .A( us01_n811 ) );
  AOI21_X1 us01_U285 (.A( us01_n810 ) , .B2( us01_n811 ) , .B1( us01_n812 ) , .ZN( us01_n817 ) );
  AOI21_X1 us01_U286 (.ZN( us01_n513 ) , .A( us01_n727 ) , .B1( us01_n748 ) , .B2( us01_n801 ) );
  AOI21_X1 us01_U287 (.ZN( us01_n497 ) , .B1( us01_n678 ) , .A( us01_n810 ) , .B2( us01_n814 ) );
  NOR2_X1 us01_U288 (.ZN( us01_n518 ) , .A2( us01_n706 ) , .A1( us01_n812 ) );
  AOI21_X1 us01_U289 (.ZN( us01_n475 ) , .A( us01_n667 ) , .B1( us01_n748 ) , .B2( us01_n804 ) );
  AOI221_X1 us01_U29 (.ZN( us01_n466 ) , .C2( us01_n712 ) , .B2( us01_n829 ) , .C1( us01_n843 ) , .B1( us01_n858 ) , .A( us01_n862 ) );
  NOR2_X1 us01_U290 (.ZN( us01_n566 ) , .A1( us01_n727 ) , .A2( us01_n760 ) );
  NOR2_X1 us01_U291 (.ZN( us01_n580 ) , .A1( us01_n742 ) , .A2( us01_n813 ) );
  AOI21_X1 us01_U292 (.ZN( us01_n591 ) , .B1( us01_n748 ) , .A( us01_n790 ) , .B2( us01_n811 ) );
  NOR2_X1 us01_U293 (.ZN( us01_n564 ) , .A2( us01_n695 ) , .A1( us01_n761 ) );
  AOI21_X1 us01_U294 (.ZN( us01_n512 ) , .A( us01_n777 ) , .B2( us01_n790 ) , .B1( us01_n810 ) );
  NAND2_X2 us01_U295 (.A2( us01_n462 ) , .A1( us01_n463 ) , .ZN( us01_n810 ) );
  AOI21_X1 us01_U296 (.ZN( us01_n637 ) , .B2( us01_n747 ) , .A( us01_n786 ) , .B1( us01_n810 ) );
  NOR2_X1 us01_U297 (.ZN( us01_n557 ) , .A2( us01_n789 ) , .A1( us01_n801 ) );
  NOR2_X1 us01_U298 (.A2( us01_n811 ) , .A1( us01_n813 ) , .ZN( us01_n819 ) );
  NOR2_X1 us01_U299 (.ZN( us01_n527 ) , .A1( us01_n706 ) , .A2( us01_n777 ) );
  NAND2_X2 us01_U3 (.A1( us01_n447 ) , .A2( us01_n462 ) , .ZN( us01_n722 ) );
  NOR4_X1 us01_U30 (.A4( us01_n512 ) , .A3( us01_n513 ) , .A2( us01_n514 ) , .A1( us01_n515 ) , .ZN( us01_n522 ) );
  NOR2_X1 us01_U300 (.ZN( us01_n517 ) , .A2( us01_n697 ) , .A1( us01_n814 ) );
  NOR2_X1 us01_U301 (.ZN( us01_n681 ) , .A2( us01_n697 ) , .A1( us01_n801 ) );
  NOR2_X1 us01_U302 (.ZN( us01_n576 ) , .A1( us01_n706 ) , .A2( us01_n811 ) );
  INV_X1 us01_U303 (.A( us01_n813 ) , .ZN( us01_n853 ) );
  INV_X1 us01_U304 (.A( us01_n811 ) , .ZN( us01_n834 ) );
  AOI21_X1 us01_U305 (.ZN( us01_n448 ) , .B2( us01_n790 ) , .A( us01_n801 ) , .B1( us01_n813 ) );
  AOI21_X1 us01_U306 (.ZN( us01_n538 ) , .A( us01_n761 ) , .B2( us01_n777 ) , .B1( us01_n815 ) );
  AOI21_X1 us01_U307 (.ZN( us01_n496 ) , .A( us01_n722 ) , .B2( us01_n760 ) , .B1( us01_n812 ) );
  AOI21_X1 us01_U308 (.ZN( us01_n687 ) , .B2( us01_n747 ) , .B1( us01_n761 ) , .A( us01_n804 ) );
  AOI21_X1 us01_U309 (.B1( us01_n684 ) , .ZN( us01_n685 ) , .A( us01_n726 ) , .B2( us01_n759 ) );
  AOI222_X1 us01_U31 (.ZN( us01_n523 ) , .A1( us01_n832 ) , .B2( us01_n835 ) , .C1( us01_n842 ) , .C2( us01_n848 ) , .A2( us01_n850 ) , .B1( us01_n864 ) );
  NOR2_X1 us01_U310 (.ZN( us01_n581 ) , .A1( us01_n790 ) , .A2( us01_n815 ) );
  NOR2_X1 us01_U311 (.ZN( us01_n532 ) , .A1( us01_n722 ) , .A2( us01_n786 ) );
  NOR2_X1 us01_U312 (.ZN( us01_n630 ) , .A2( us01_n695 ) , .A1( us01_n722 ) );
  AOI21_X1 us01_U313 (.A( us01_n788 ) , .B2( us01_n789 ) , .B1( us01_n790 ) , .ZN( us01_n791 ) );
  AOI21_X1 us01_U314 (.A( us01_n731 ) , .ZN( us01_n732 ) , .B2( us01_n778 ) , .B1( us01_n790 ) );
  NOR2_X1 us01_U315 (.ZN( us01_n565 ) , .A1( us01_n745 ) , .A2( us01_n803 ) );
  AOI21_X1 us01_U316 (.ZN( us01_n567 ) , .B1( us01_n748 ) , .B2( us01_n760 ) , .A( us01_n778 ) );
  AOI21_X1 us01_U317 (.ZN( us01_n638 ) , .B2( us01_n745 ) , .A( us01_n790 ) , .B1( us01_n801 ) );
  AOI21_X1 us01_U318 (.ZN( us01_n562 ) , .B1( us01_n722 ) , .A( us01_n777 ) , .B2( us01_n789 ) );
  AOI21_X1 us01_U319 (.ZN( us01_n569 ) , .B2( us01_n695 ) , .B1( us01_n804 ) , .A( us01_n810 ) );
  NOR4_X1 us01_U32 (.A3( us01_n519 ) , .A1( us01_n520 ) , .ZN( us01_n521 ) , .A2( us01_n671 ) , .A4( us01_n767 ) );
  NOR2_X1 us01_U320 (.ZN( us01_n663 ) , .A1( us01_n778 ) , .A2( us01_n811 ) );
  NOR2_X1 us01_U321 (.ZN( us01_n578 ) , .A2( us01_n695 ) , .A1( us01_n789 ) );
  NOR2_X1 us01_U322 (.ZN( us01_n682 ) , .A1( us01_n789 ) , .A2( us01_n811 ) );
  NAND2_X2 us01_U323 (.A1( us01_n450 ) , .A2( us01_n463 ) , .ZN( us01_n667 ) );
  NAND2_X1 us01_U324 (.ZN( us01_n751 ) , .A1( us01_n761 ) , .A2( us01_n803 ) );
  NOR2_X1 us01_U325 (.ZN( us01_n709 ) , .A1( us01_n760 ) , .A2( us01_n761 ) );
  AOI21_X1 us01_U326 (.ZN( us01_n476 ) , .B2( us01_n695 ) , .A( us01_n747 ) , .B1( us01_n777 ) );
  NOR2_X1 us01_U327 (.ZN( us01_n680 ) , .A2( us01_n706 ) , .A1( us01_n815 ) );
  INV_X1 us01_U328 (.A( us01_n778 ) , .ZN( us01_n848 ) );
  OAI21_X1 us01_U329 (.A( us01_n729 ) , .B1( us01_n730 ) , .ZN( us01_n734 ) , .B2( us01_n803 ) );
  AOI221_X1 us01_U33 (.A( us01_n779 ) , .ZN( us01_n796 ) , .C2( us01_n835 ) , .B2( us01_n836 ) , .B1( us01_n863 ) , .C1( us01_n864 ) );
  OAI21_X1 us01_U330 (.ZN( us01_n729 ) , .A( us01_n831 ) , .B2( us01_n850 ) , .B1( us01_n871 ) );
  AOI21_X1 us01_U331 (.ZN( us01_n639 ) , .B1( us01_n678 ) , .A( us01_n789 ) , .B2( us01_n815 ) );
  AOI21_X1 us01_U332 (.ZN( us01_n440 ) , .A( us01_n697 ) , .B1( us01_n731 ) , .B2( us01_n748 ) );
  NAND2_X1 us01_U333 (.A1( us01_n697 ) , .A2( us01_n727 ) , .ZN( us01_n780 ) );
  NOR2_X1 us01_U334 (.ZN( us01_n468 ) , .A2( us01_n777 ) , .A1( us01_n813 ) );
  NOR2_X1 us01_U335 (.ZN( us01_n516 ) , .A1( us01_n706 ) , .A2( us01_n786 ) );
  NAND2_X2 us01_U336 (.A2( us01_n447 ) , .A1( us01_n450 ) , .ZN( us01_n761 ) );
  OAI21_X1 us01_U337 (.A( us01_n696 ) , .ZN( us01_n700 ) , .B2( us01_n748 ) , .B1( us01_n802 ) );
  OAI21_X1 us01_U338 (.ZN( us01_n696 ) , .B2( us01_n831 ) , .B1( us01_n836 ) , .A( us01_n858 ) );
  NOR2_X1 us01_U339 (.ZN( us01_n524 ) , .A1( us01_n722 ) , .A2( us01_n748 ) );
  NOR4_X1 us01_U34 (.A4( us01_n791 ) , .A3( us01_n792 ) , .A2( us01_n793 ) , .A1( us01_n794 ) , .ZN( us01_n795 ) );
  AOI21_X1 us01_U340 (.ZN( us01_n441 ) , .B1( us01_n787 ) , .B2( us01_n789 ) , .A( us01_n812 ) );
  AOI21_X1 us01_U341 (.ZN( us01_n495 ) , .A( us01_n777 ) , .B2( us01_n789 ) , .B1( us01_n802 ) );
  NAND2_X1 us01_U342 (.ZN( us01_n712 ) , .A1( us01_n726 ) , .A2( us01_n778 ) );
  NOR2_X1 us01_U343 (.ZN( us01_n482 ) , .A1( us01_n786 ) , .A2( us01_n803 ) );
  NAND2_X1 us01_U344 (.A2( us01_n760 ) , .A1( us01_n804 ) , .ZN( us01_n808 ) );
  OAI21_X1 us01_U345 (.A( us01_n785 ) , .B2( us01_n786 ) , .B1( us01_n787 ) , .ZN( us01_n793 ) );
  OAI21_X1 us01_U346 (.ZN( us01_n785 ) , .A( us01_n837 ) , .B1( us01_n861 ) , .B2( us01_n871 ) );
  INV_X1 us01_U347 (.A( us01_n783 ) , .ZN( us01_n844 ) );
  NOR2_X1 us01_U348 (.ZN( us01_n710 ) , .A2( us01_n722 ) , .A1( us01_n788 ) );
  NAND2_X1 us01_U349 (.ZN( us01_n669 ) , .A1( us01_n804 ) , .A2( us01_n814 ) );
  NOR4_X1 us01_U35 (.A4( us01_n774 ) , .A3( us01_n775 ) , .A1( us01_n776 ) , .ZN( us01_n797 ) , .A2( us01_n799 ) );
  NAND2_X2 us01_U350 (.A2( us01_n446 ) , .A1( us01_n450 ) , .ZN( us01_n727 ) );
  INV_X1 us01_U351 (.A( us01_n722 ) , .ZN( us01_n854 ) );
  NAND2_X2 us01_U352 (.A1( us01_n445 ) , .A2( us01_n463 ) , .ZN( us01_n747 ) );
  INV_X1 us01_U353 (.A( us01_n815 ) , .ZN( us01_n842 ) );
  AND2_X1 us01_U354 (.ZN( us01_n730 ) , .A1( us01_n777 ) , .A2( us01_n783 ) );
  NAND2_X1 us01_U355 (.A1( us01_n445 ) , .A2( us01_n447 ) , .ZN( us01_n803 ) );
  NAND2_X1 us01_U356 (.A1( us01_n449 ) , .A2( us01_n452 ) , .ZN( us01_n812 ) );
  NAND2_X1 us01_U357 (.A1( us01_n453 ) , .A2( us01_n469 ) , .ZN( us01_n801 ) );
  NAND2_X1 us01_U358 (.A1( us01_n453 ) , .A2( us01_n460 ) , .ZN( us01_n748 ) );
  NAND2_X2 us01_U359 (.A2( us01_n446 ) , .A1( us01_n458 ) , .ZN( us01_n726 ) );
  NOR2_X1 us01_U36 (.ZN( us01_n802 ) , .A1( us01_n852 ) , .A2( us01_n859 ) );
  NAND2_X1 us01_U360 (.A2( us01_n451 ) , .A1( us01_n453 ) , .ZN( us01_n804 ) );
  NAND2_X1 us01_U361 (.A1( us01_n449 ) , .A2( us01_n469 ) , .ZN( us01_n814 ) );
  NAND2_X1 us01_U362 (.A1( us01_n452 ) , .A2( us01_n459 ) , .ZN( us01_n811 ) );
  NAND2_X1 us01_U363 (.A1( us01_n451 ) , .A2( us01_n459 ) , .ZN( us01_n742 ) );
  NAND2_X1 us01_U364 (.A1( us01_n451 ) , .A2( us01_n470 ) , .ZN( us01_n783 ) );
  NAND2_X1 us01_U365 (.A2( us01_n452 ) , .A1( us01_n470 ) , .ZN( us01_n777 ) );
  NAND2_X1 us01_U366 (.A2( us01_n459 ) , .A1( us01_n460 ) , .ZN( us01_n745 ) );
  NAND2_X2 us01_U367 (.A2( us01_n446 ) , .A1( us01_n462 ) , .ZN( us01_n813 ) );
  NAND2_X1 us01_U368 (.A1( us01_n460 ) , .A2( us01_n470 ) , .ZN( us01_n786 ) );
  NOR2_X1 us01_U369 (.ZN( us01_n451 ) , .A1( us01_n824 ) , .A2( us01_n825 ) );
  NAND4_X1 us01_U37 (.ZN( sa01_sr_2 ) , .A4( us01_n641 ) , .A3( us01_n642 ) , .A2( us01_n643 ) , .A1( us01_n644 ) );
  NOR2_X1 us01_U370 (.ZN( us01_n449 ) , .A1( us01_n826 ) , .A2( us01_n827 ) );
  NAND2_X1 us01_U371 (.A1( us01_n449 ) , .A2( us01_n460 ) , .ZN( us01_n788 ) );
  NAND2_X2 us01_U372 (.A1( us01_n447 ) , .A2( us01_n458 ) , .ZN( us01_n790 ) );
  NAND2_X2 us01_U373 (.A2( us01_n439 ) , .A1( us01_n450 ) , .ZN( us01_n789 ) );
  NAND2_X1 us01_U374 (.A2( us01_n452 ) , .A1( us01_n453 ) , .ZN( us01_n728 ) );
  NAND2_X2 us01_U375 (.A2( us01_n469 ) , .A1( us01_n470 ) , .ZN( us01_n815 ) );
  NAND2_X1 us01_U376 (.A1( us01_n445 ) , .A2( us01_n446 ) , .ZN( us01_n784 ) );
  NAND2_X2 us01_U377 (.A2( us01_n439 ) , .A1( us01_n445 ) , .ZN( us01_n782 ) );
  NOR2_X1 us01_U378 (.A2( sa01_7 ) , .ZN( us01_n458 ) , .A1( us01_n847 ) );
  NOR2_X1 us01_U379 (.A2( sa01_2 ) , .A1( sa01_3 ) , .ZN( us01_n470 ) );
  AOI222_X1 us01_U38 (.B2( us01_n636 ) , .ZN( us01_n642 ) , .B1( us01_n839 ) , .A1( us01_n840 ) , .C2( us01_n844 ) , .C1( us01_n861 ) , .A2( us01_n863 ) );
  NOR2_X1 us01_U380 (.A2( sa01_1 ) , .ZN( us01_n469 ) , .A1( us01_n824 ) );
  NOR2_X1 us01_U381 (.A2( sa01_0 ) , .ZN( us01_n452 ) , .A1( us01_n825 ) );
  NOR2_X1 us01_U382 (.A2( sa01_0 ) , .A1( sa01_1 ) , .ZN( us01_n460 ) );
  NAND2_X2 us01_U383 (.A1( us01_n439 ) , .A2( us01_n458 ) , .ZN( us01_n697 ) );
  NOR2_X1 us01_U384 (.A2( sa01_3 ) , .ZN( us01_n453 ) , .A1( us01_n826 ) );
  NOR2_X1 us01_U385 (.A2( sa01_2 ) , .ZN( us01_n459 ) , .A1( us01_n827 ) );
  INV_X1 us01_U386 (.A( sa01_3 ) , .ZN( us01_n827 ) );
  INV_X1 us01_U387 (.A( sa01_1 ) , .ZN( us01_n825 ) );
  INV_X1 us01_U388 (.A( sa01_0 ) , .ZN( us01_n824 ) );
  INV_X1 us01_U389 (.A( sa01_2 ) , .ZN( us01_n826 ) );
  NOR4_X1 us01_U39 (.A4( us01_n637 ) , .A3( us01_n638 ) , .A2( us01_n639 ) , .A1( us01_n640 ) , .ZN( us01_n641 ) );
  INV_X1 us01_U390 (.A( sa01_5 ) , .ZN( us01_n846 ) );
  NAND2_X1 us01_U391 (.A1( us01_n727 ) , .A2( us01_n782 ) , .ZN( us01_n809 ) );
  OAI22_X1 us01_U392 (.ZN( us01_n586 ) , .A2( us01_n745 ) , .B2( us01_n760 ) , .A1( us01_n761 ) , .B1( us01_n782 ) );
  AOI21_X1 us01_U393 (.ZN( us01_n590 ) , .B1( us01_n726 ) , .B2( us01_n782 ) , .A( us01_n788 ) );
  AOI21_X1 us01_U394 (.ZN( us01_n646 ) , .A( us01_n760 ) , .B2( us01_n782 ) , .B1( us01_n790 ) );
  AOI21_X1 us01_U395 (.ZN( us01_n621 ) , .B1( us01_n697 ) , .A( us01_n777 ) , .B2( us01_n782 ) );
  OAI22_X1 us01_U396 (.ZN( us01_n679 ) , .A1( us01_n697 ) , .A2( us01_n728 ) , .B2( us01_n782 ) , .B1( us01_n815 ) );
  OAI21_X1 us01_U397 (.A( us01_n611 ) , .ZN( us01_n614 ) , .B1( us01_n623 ) , .B2( us01_n782 ) );
  NOR2_X1 us01_U398 (.ZN( us01_n608 ) , .A1( us01_n782 ) , .A2( us01_n814 ) );
  INV_X2 us01_U399 (.A( us01_n747 ) , .ZN( us01_n861 ) );
  NAND2_X2 us01_U4 (.A1( us01_n439 ) , .A2( us01_n462 ) , .ZN( us01_n706 ) );
  NOR3_X1 us01_U40 (.A2( us01_n605 ) , .A1( us01_n606 ) , .ZN( us01_n644 ) , .A3( us01_n720 ) );
  OAI222_X1 us01_U400 (.A2( us01_n667 ) , .ZN( us01_n672 ) , .B1( us01_n745 ) , .B2( us01_n782 ) , .C2( us01_n786 ) , .C1( us01_n813 ) , .A1( us01_n815 ) );
  NOR2_X1 us01_U401 (.ZN( us01_n649 ) , .A1( us01_n782 ) , .A2( us01_n786 ) );
  NOR2_X1 us01_U402 (.ZN( us01_n598 ) , .A2( us01_n695 ) , .A1( us01_n782 ) );
  NOR2_X1 us01_U403 (.ZN( us01_n551 ) , .A2( us01_n742 ) , .A1( us01_n782 ) );
  INV_X1 us01_U404 (.A( us01_n782 ) , .ZN( us01_n859 ) );
  NAND2_X1 us01_U405 (.A2( us01_n459 ) , .A1( us01_n469 ) , .ZN( us01_n695 ) );
  INV_X1 us01_U406 (.A( sa01_7 ) , .ZN( us01_n856 ) );
  OAI221_X1 us01_U407 (.A( us01_n781 ) , .C2( us01_n782 ) , .B2( us01_n783 ) , .B1( us01_n784 ) , .ZN( us01_n794 ) , .C1( us01_n811 ) );
  AOI21_X1 us01_U408 (.ZN( us01_n498 ) , .A( us01_n695 ) , .B1( us01_n706 ) , .B2( us01_n784 ) );
  OAI221_X1 us01_U409 (.A( us01_n694 ) , .ZN( us01_n701 ) , .C2( us01_n782 ) , .C1( us01_n783 ) , .B1( us01_n784 ) , .B2( us01_n804 ) );
  NAND4_X1 us01_U41 (.ZN( sa01_sr_7 ) , .A4( us01_n820 ) , .A3( us01_n821 ) , .A2( us01_n822 ) , .A1( us01_n823 ) );
  OAI22_X1 us01_U410 (.ZN( us01_n588 ) , .B1( us01_n728 ) , .B2( us01_n747 ) , .A2( us01_n784 ) , .A1( us01_n801 ) );
  AOI222_X1 us01_U411 (.ZN( us01_n511 ) , .C1( us01_n830 ) , .B2( us01_n835 ) , .A2( us01_n841 ) , .C2( us01_n860 ) , .B1( us01_n861 ) , .A1( us01_n864 ) );
  AOI222_X1 us01_U412 (.ZN( us01_n603 ) , .B2( us01_n669 ) , .B1( us01_n751 ) , .C2( us01_n829 ) , .A1( us01_n831 ) , .A2( us01_n860 ) , .C1( us01_n861 ) );
  AOI221_X1 us01_U413 (.A( us01_n481 ) , .ZN( us01_n486 ) , .B1( us01_n829 ) , .C2( us01_n842 ) , .C1( us01_n850 ) , .B2( us01_n860 ) );
  NAND2_X1 us01_U414 (.A2( us01_n747 ) , .A1( us01_n784 ) , .ZN( us01_n807 ) );
  NOR2_X1 us01_U415 (.ZN( us01_n610 ) , .A1( us01_n777 ) , .A2( us01_n784 ) );
  NOR2_X1 us01_U416 (.ZN( us01_n715 ) , .A2( us01_n742 ) , .A1( us01_n784 ) );
  OAI222_X1 us01_U417 (.ZN( us01_n615 ) , .B1( us01_n695 ) , .C1( us01_n722 ) , .C2( us01_n745 ) , .B2( us01_n784 ) , .A2( us01_n790 ) , .A1( us01_n814 ) );
  NOR2_X1 us01_U418 (.ZN( us01_n651 ) , .A1( us01_n760 ) , .A2( us01_n784 ) );
  NOR2_X1 us01_U419 (.ZN( us01_n552 ) , .A1( us01_n784 ) , .A2( us01_n811 ) );
  AOI222_X1 us01_U42 (.C2( us01_n807 ) , .B2( us01_n808 ) , .A2( us01_n809 ) , .ZN( us01_n821 ) , .C1( us01_n830 ) , .A1( us01_n837 ) , .B1( us01_n851 ) );
  NOR2_X1 us01_U420 (.ZN( us01_n787 ) , .A2( us01_n860 ) , .A1( us01_n866 ) );
  NOR2_X1 us01_U421 (.ZN( us01_n699 ) , .A2( us01_n784 ) , .A1( us01_n815 ) );
  NOR2_X1 us01_U422 (.A1( us01_n728 ) , .ZN( us01_n763 ) , .A2( us01_n784 ) );
  INV_X1 us01_U423 (.A( us01_n784 ) , .ZN( us01_n860 ) );
  NOR2_X1 us01_U424 (.A2( sa01_4 ) , .ZN( us01_n447 ) , .A1( us01_n846 ) );
  NOR2_X1 us01_U425 (.ZN( us01_n463 ) , .A2( us01_n845 ) , .A1( us01_n846 ) );
  NOR2_X1 us01_U426 (.A2( sa01_5 ) , .ZN( us01_n446 ) , .A1( us01_n845 ) );
  NOR2_X1 us01_U427 (.A2( sa01_4 ) , .A1( sa01_5 ) , .ZN( us01_n439 ) );
  INV_X1 us01_U428 (.A( sa01_6 ) , .ZN( us01_n847 ) );
  NOR2_X1 us01_U429 (.ZN( us01_n445 ) , .A2( us01_n847 ) , .A1( us01_n856 ) );
  NOR4_X1 us01_U43 (.A4( us01_n816 ) , .A3( us01_n817 ) , .A2( us01_n818 ) , .A1( us01_n819 ) , .ZN( us01_n820 ) );
  NOR2_X1 us01_U430 (.A2( sa01_6 ) , .ZN( us01_n450 ) , .A1( us01_n856 ) );
  NOR2_X1 us01_U431 (.A2( sa01_6 ) , .A1( sa01_7 ) , .ZN( us01_n462 ) );
  AOI221_X1 us01_U432 (.A( us01_n574 ) , .ZN( us01_n585 ) , .B2( us01_n829 ) , .C2( us01_n841 ) , .B1( us01_n852 ) , .C1( us01_n859 ) );
  AOI21_X1 us01_U433 (.ZN( us01_n574 ) , .B2( us01_n722 ) , .B1( us01_n746 ) , .A( us01_n783 ) );
  INV_X1 us01_U434 (.A( sa01_4 ) , .ZN( us01_n845 ) );
  AOI211_X1 us01_U435 (.A( us01_n635 ) , .ZN( us01_n643 ) , .B( us01_n741 ) , .C2( us01_n837 ) , .C1( us01_n852 ) );
  NAND4_X1 us01_U436 (.A4( us01_n631 ) , .A3( us01_n632 ) , .A2( us01_n633 ) , .A1( us01_n634 ) , .ZN( us01_n741 ) );
  NAND3_X1 us01_U437 (.ZN( sa01_sr_6 ) , .A3( us01_n795 ) , .A2( us01_n796 ) , .A1( us01_n797 ) );
  NAND3_X1 us01_U438 (.ZN( sa01_sr_5 ) , .A3( us01_n756 ) , .A2( us01_n757 ) , .A1( us01_n758 ) );
  NAND3_X1 us01_U439 (.ZN( sa01_sr_4 ) , .A3( us01_n736 ) , .A2( us01_n737 ) , .A1( us01_n738 ) );
  AOI211_X1 us01_U44 (.B( us01_n805 ) , .A( us01_n806 ) , .ZN( us01_n822 ) , .C1( us01_n840 ) , .C2( us01_n848 ) );
  NAND3_X1 us01_U440 (.A3( us01_n673 ) , .A2( us01_n674 ) , .A1( us01_n675 ) , .ZN( us01_n805 ) );
  NAND3_X1 us01_U441 (.ZN( us01_n636 ) , .A3( us01_n706 ) , .A2( us01_n722 ) , .A1( us01_n790 ) );
  NAND3_X1 us01_U442 (.A3( us01_n616 ) , .A2( us01_n617 ) , .A1( us01_n618 ) , .ZN( us01_n723 ) );
  NAND3_X1 us01_U443 (.A3( us01_n583 ) , .A2( us01_n584 ) , .A1( us01_n585 ) , .ZN( us01_n619 ) );
  NAND3_X1 us01_U444 (.ZN( us01_n563 ) , .A3( us01_n678 ) , .A2( us01_n748 ) , .A1( us01_n783 ) );
  NAND3_X1 us01_U445 (.A3( us01_n521 ) , .A2( us01_n522 ) , .A1( us01_n523 ) , .ZN( us01_n740 ) );
  NAND3_X1 us01_U446 (.A3( us01_n510 ) , .A1( us01_n511 ) , .ZN( us01_n606 ) , .A2( us01_n869 ) );
  NAND3_X1 us01_U447 (.A3( us01_n465 ) , .A2( us01_n466 ) , .A1( us01_n467 ) , .ZN( us01_n775 ) );
  NAND4_X1 us01_U45 (.ZN( sa01_sr_0 ) , .A4( us01_n499 ) , .A3( us01_n500 ) , .A2( us01_n501 ) , .A1( us01_n502 ) );
  NOR4_X1 us01_U46 (.A4( us01_n496 ) , .A3( us01_n497 ) , .A2( us01_n498 ) , .ZN( us01_n499 ) , .A1( us01_n525 ) );
  AOI221_X1 us01_U47 (.A( us01_n495 ) , .ZN( us01_n500 ) , .B2( us01_n841 ) , .C1( us01_n844 ) , .C2( us01_n858 ) , .B1( us01_n860 ) );
  AOI211_X1 us01_U48 (.A( us01_n494 ) , .ZN( us01_n501 ) , .B( us01_n800 ) , .C2( us01_n837 ) , .C1( us01_n849 ) );
  NOR2_X1 us01_U49 (.ZN( us01_n746 ) , .A1( us01_n859 ) , .A2( us01_n860 ) );
  NAND2_X2 us01_U5 (.A2( us01_n458 ) , .A1( us01_n463 ) , .ZN( us01_n778 ) );
  NAND4_X1 us01_U50 (.ZN( sa01_sr_1 ) , .A4( us01_n593 ) , .A3( us01_n594 ) , .A2( us01_n595 ) , .A1( us01_n596 ) );
  AOI211_X1 us01_U51 (.B( us01_n587 ) , .A( us01_n588 ) , .ZN( us01_n594 ) , .C2( us01_n809 ) , .C1( us01_n831 ) );
  NOR4_X1 us01_U52 (.A4( us01_n589 ) , .A3( us01_n590 ) , .A2( us01_n591 ) , .A1( us01_n592 ) , .ZN( us01_n593 ) );
  AOI211_X1 us01_U53 (.A( us01_n586 ) , .ZN( us01_n595 ) , .B( us01_n619 ) , .C1( us01_n843 ) , .C2( us01_n853 ) );
  NOR2_X1 us01_U54 (.ZN( us01_n623 ) , .A2( us01_n834 ) , .A1( us01_n837 ) );
  NAND4_X1 us01_U55 (.A4( us01_n601 ) , .A3( us01_n602 ) , .A2( us01_n603 ) , .A1( us01_n604 ) , .ZN( us01_n720 ) );
  NOR3_X1 us01_U56 (.A1( us01_n597 ) , .ZN( us01_n602 ) , .A3( us01_n661 ) , .A2( us01_n768 ) );
  NOR4_X1 us01_U57 (.A3( us01_n598 ) , .A2( us01_n599 ) , .A1( us01_n600 ) , .ZN( us01_n601 ) , .A4( us01_n653 ) );
  AOI222_X1 us01_U58 (.ZN( us01_n604 ) , .A1( us01_n828 ) , .C2( us01_n835 ) , .B1( us01_n840 ) , .A2( us01_n854 ) , .B2( us01_n859 ) , .C1( us01_n866 ) );
  NOR4_X1 us01_U59 (.A4( us01_n575 ) , .A3( us01_n576 ) , .A2( us01_n577 ) , .ZN( us01_n584 ) , .A1( us01_n681 ) );
  INV_X1 us01_U6 (.A( us01_n667 ) , .ZN( us01_n863 ) );
  NOR4_X1 us01_U60 (.A1( us01_n582 ) , .ZN( us01_n583 ) , .A3( us01_n650 ) , .A2( us01_n660 ) , .A4( us01_n765 ) );
  NAND4_X1 us01_U61 (.A4( us01_n483 ) , .A3( us01_n484 ) , .A2( us01_n485 ) , .A1( us01_n486 ) , .ZN( us01_n776 ) );
  NOR4_X1 us01_U62 (.A4( us01_n482 ) , .ZN( us01_n485 ) , .A1( us01_n564 ) , .A2( us01_n579 ) , .A3( us01_n600 ) );
  NOR4_X1 us01_U63 (.ZN( us01_n483 ) , .A2( us01_n531 ) , .A1( us01_n556 ) , .A3( us01_n629 ) , .A4( us01_n716 ) );
  NOR4_X1 us01_U64 (.ZN( us01_n484 ) , .A1( us01_n505 ) , .A2( us01_n517 ) , .A4( us01_n544 ) , .A3( us01_n609 ) );
  NOR4_X1 us01_U65 (.A4( us01_n627 ) , .A3( us01_n628 ) , .A2( us01_n629 ) , .A1( us01_n630 ) , .ZN( us01_n631 ) );
  AOI211_X1 us01_U66 (.B( us01_n621 ) , .A( us01_n622 ) , .ZN( us01_n633 ) , .C2( us01_n834 ) , .C1( us01_n861 ) );
  NOR4_X1 us01_U67 (.A4( us01_n624 ) , .A3( us01_n625 ) , .A2( us01_n626 ) , .ZN( us01_n632 ) , .A1( us01_n662 ) );
  NAND4_X1 us01_U68 (.A4( us01_n655 ) , .A3( us01_n656 ) , .A2( us01_n657 ) , .A1( us01_n658 ) , .ZN( us01_n798 ) );
  NOR3_X1 us01_U69 (.A3( us01_n649 ) , .A2( us01_n650 ) , .A1( us01_n651 ) , .ZN( us01_n656 ) );
  NOR3_X1 us01_U7 (.ZN( us01_n596 ) , .A1( us01_n606 ) , .A3( us01_n721 ) , .A2( us01_n740 ) );
  NOR3_X1 us01_U70 (.A3( us01_n652 ) , .A2( us01_n653 ) , .A1( us01_n654 ) , .ZN( us01_n655 ) );
  NOR3_X1 us01_U71 (.A3( us01_n646 ) , .A2( us01_n647 ) , .A1( us01_n648 ) , .ZN( us01_n657 ) );
  NAND4_X1 us01_U72 (.A4( us01_n558 ) , .A3( us01_n559 ) , .A2( us01_n560 ) , .A1( us01_n561 ) , .ZN( us01_n605 ) );
  NOR4_X1 us01_U73 (.ZN( us01_n559 ) , .A1( us01_n651 ) , .A3( us01_n659 ) , .A4( us01_n683 ) , .A2( us01_n766 ) );
  NOR4_X1 us01_U74 (.A4( us01_n550 ) , .A3( us01_n551 ) , .A2( us01_n552 ) , .A1( us01_n553 ) , .ZN( us01_n560 ) );
  NOR4_X1 us01_U75 (.A4( us01_n554 ) , .A3( us01_n555 ) , .A2( us01_n556 ) , .A1( us01_n557 ) , .ZN( us01_n558 ) );
  NAND4_X1 us01_U76 (.A4( us01_n770 ) , .A3( us01_n771 ) , .A2( us01_n772 ) , .A1( us01_n773 ) , .ZN( us01_n799 ) );
  NOR3_X1 us01_U77 (.A3( us01_n763 ) , .A2( us01_n764 ) , .A1( us01_n765 ) , .ZN( us01_n771 ) );
  NOR4_X1 us01_U78 (.A4( us01_n766 ) , .A3( us01_n767 ) , .A2( us01_n768 ) , .A1( us01_n769 ) , .ZN( us01_n770 ) );
  AOI222_X1 us01_U79 (.ZN( us01_n773 ) , .A1( us01_n828 ) , .C1( us01_n832 ) , .B2( us01_n839 ) , .A2( us01_n848 ) , .B1( us01_n859 ) , .C2( us01_n871 ) );
  NOR3_X1 us01_U8 (.A3( us01_n798 ) , .A2( us01_n799 ) , .A1( us01_n800 ) , .ZN( us01_n823 ) );
  NOR4_X1 us01_U80 (.A4( us01_n507 ) , .A2( us01_n508 ) , .A1( us01_n509 ) , .ZN( us01_n510 ) , .A3( us01_n668 ) );
  INV_X1 us01_U81 (.A( us01_n503 ) , .ZN( us01_n869 ) );
  NOR4_X1 us01_U82 (.A4( us01_n663 ) , .A3( us01_n664 ) , .A2( us01_n665 ) , .A1( us01_n666 ) , .ZN( us01_n674 ) );
  NOR4_X1 us01_U83 (.A4( us01_n659 ) , .A3( us01_n660 ) , .A2( us01_n661 ) , .A1( us01_n662 ) , .ZN( us01_n675 ) );
  NOR4_X1 us01_U84 (.A3( us01_n671 ) , .A1( us01_n672 ) , .ZN( us01_n673 ) , .A4( us01_n713 ) , .A2( us01_n857 ) );
  NOR2_X1 us01_U85 (.ZN( us01_n759 ) , .A1( us01_n831 ) , .A2( us01_n832 ) );
  NAND4_X1 us01_U86 (.A4( us01_n454 ) , .A3( us01_n455 ) , .A2( us01_n456 ) , .A1( us01_n457 ) , .ZN( us01_n677 ) );
  NOR3_X1 us01_U87 (.ZN( us01_n455 ) , .A3( us01_n528 ) , .A1( us01_n553 ) , .A2( us01_n568 ) );
  AOI221_X1 us01_U88 (.A( us01_n448 ) , .ZN( us01_n457 ) , .C2( us01_n751 ) , .B1( us01_n830 ) , .C1( us01_n840 ) , .B2( us01_n859 ) );
  NOR4_X1 us01_U89 (.ZN( us01_n456 ) , .A2( us01_n507 ) , .A1( us01_n597 ) , .A4( us01_n626 ) , .A3( us01_n709 ) );
  NOR3_X1 us01_U9 (.A3( us01_n619 ) , .A2( us01_n620 ) , .ZN( us01_n634 ) , .A1( us01_n723 ) );
  NAND4_X1 us01_U90 (.A4( us01_n533 ) , .A3( us01_n534 ) , .A2( us01_n535 ) , .A1( us01_n536 ) , .ZN( us01_n620 ) );
  NOR4_X1 us01_U91 (.A4( us01_n524 ) , .A2( us01_n525 ) , .A1( us01_n526 ) , .ZN( us01_n536 ) , .A3( us01_n699 ) );
  NOR4_X1 us01_U92 (.A1( us01_n529 ) , .ZN( us01_n534 ) , .A2( us01_n652 ) , .A4( us01_n666 ) , .A3( us01_n763 ) );
  NOR4_X1 us01_U93 (.A4( us01_n527 ) , .A3( us01_n528 ) , .ZN( us01_n535 ) , .A2( us01_n682 ) , .A1( us01_n792 ) );
  NAND4_X1 us01_U94 (.A4( us01_n477 ) , .A3( us01_n478 ) , .A2( us01_n479 ) , .A1( us01_n480 ) , .ZN( us01_n692 ) );
  NOR3_X1 us01_U95 (.ZN( us01_n478 ) , .A2( us01_n506 ) , .A3( us01_n599 ) , .A1( us01_n608 ) );
  AOI211_X1 us01_U96 (.B( us01_n475 ) , .A( us01_n476 ) , .ZN( us01_n480 ) , .C2( us01_n831 ) , .C1( us01_n859 ) );
  NOR4_X1 us01_U97 (.ZN( us01_n479 ) , .A3( us01_n530 ) , .A4( us01_n543 ) , .A2( us01_n565 ) , .A1( us01_n715 ) );
  NAND4_X1 us01_U98 (.A4( us01_n546 ) , .A3( us01_n547 ) , .A2( us01_n548 ) , .A1( us01_n549 ) , .ZN( us01_n743 ) );
  NOR3_X1 us01_U99 (.ZN( us01_n547 ) , .A2( us01_n649 ) , .A1( us01_n665 ) , .A3( us01_n769 ) );
  INV_X1 us20_U10 (.A( us20_n706 ) , .ZN( us20_n876 ) );
  NOR4_X1 us20_U100 (.A1( us20_n531 ) , .ZN( us20_n536 ) , .A2( us20_n654 ) , .A4( us20_n668 ) , .A3( us20_n765 ) );
  NOR4_X1 us20_U101 (.A4( us20_n529 ) , .A3( us20_n530 ) , .ZN( us20_n537 ) , .A2( us20_n684 ) , .A1( us20_n794 ) );
  NAND4_X1 us20_U102 (.A4( us20_n548 ) , .A3( us20_n549 ) , .A2( us20_n550 ) , .A1( us20_n551 ) , .ZN( us20_n745 ) );
  NOR3_X1 us20_U103 (.ZN( us20_n549 ) , .A2( us20_n651 ) , .A1( us20_n667 ) , .A3( us20_n771 ) );
  AOI211_X1 us20_U104 (.B( us20_n539 ) , .A( us20_n540 ) , .ZN( us20_n551 ) , .C2( us20_n839 ) , .C1( us20_n851 ) );
  NOR4_X1 us20_U105 (.A4( us20_n541 ) , .A3( us20_n542 ) , .A2( us20_n543 ) , .ZN( us20_n550 ) , .A1( us20_n688 ) );
  NAND4_X1 us20_U106 (.A4( us20_n479 ) , .A3( us20_n480 ) , .A2( us20_n481 ) , .A1( us20_n482 ) , .ZN( us20_n694 ) );
  NOR3_X1 us20_U107 (.ZN( us20_n480 ) , .A2( us20_n508 ) , .A3( us20_n601 ) , .A1( us20_n610 ) );
  AOI211_X1 us20_U108 (.B( us20_n477 ) , .A( us20_n478 ) , .ZN( us20_n482 ) , .C2( us20_n833 ) , .C1( us20_n861 ) );
  NOR4_X1 us20_U109 (.ZN( us20_n481 ) , .A3( us20_n532 ) , .A4( us20_n545 ) , .A2( us20_n567 ) , .A1( us20_n717 ) );
  INV_X1 us20_U11 (.A( us20_n607 ) , .ZN( us20_n874 ) );
  NOR2_X1 us20_U110 (.ZN( us20_n647 ) , .A1( us20_n854 ) , .A2( us20_n868 ) );
  NAND4_X1 us20_U111 (.A4( us20_n473 ) , .A3( us20_n474 ) , .A2( us20_n475 ) , .A1( us20_n476 ) , .ZN( us20_n678 ) );
  NOR4_X1 us20_U112 (.ZN( us20_n475 ) , .A1( us20_n531 ) , .A3( us20_n568 ) , .A4( us20_n600 ) , .A2( us20_n642 ) );
  NOR4_X1 us20_U113 (.A4( us20_n470 ) , .ZN( us20_n476 ) , .A3( us20_n556 ) , .A1( us20_n735 ) , .A2( us20_n755 ) );
  NOR4_X1 us20_U114 (.ZN( us20_n474 ) , .A1( us20_n506 ) , .A3( us20_n544 ) , .A2( us20_n583 ) , .A4( us20_n716 ) );
  NAND4_X1 us20_U115 (.A4( us20_n691 ) , .A3( us20_n692 ) , .A1( us20_n693 ) , .ZN( us20_n776 ) , .A2( us20_n872 ) );
  INV_X1 us20_U116 (.A( us20_n679 ) , .ZN( us20_n872 ) );
  AOI221_X1 us20_U117 (.A( us20_n681 ) , .ZN( us20_n692 ) , .B2( us20_n840 ) , .C1( us20_n842 ) , .C2( us20_n862 ) , .B1( us20_n865 ) );
  NOR4_X1 us20_U118 (.A4( us20_n687 ) , .A3( us20_n688 ) , .A2( us20_n689 ) , .A1( us20_n690 ) , .ZN( us20_n691 ) );
  NOR2_X1 us20_U119 (.ZN( us20_n733 ) , .A2( us20_n832 ) , .A1( us20_n845 ) );
  INV_X1 us20_U12 (.A( us20_n680 ) , .ZN( us20_n840 ) );
  NAND4_X1 us20_U120 (.A4( us20_n719 ) , .A3( us20_n720 ) , .A2( us20_n721 ) , .ZN( us20_n741 ) , .A1( us20_n857 ) );
  INV_X1 us20_U121 (.A( us20_n709 ) , .ZN( us20_n857 ) );
  NOR4_X1 us20_U122 (.A4( us20_n715 ) , .A3( us20_n716 ) , .A2( us20_n717 ) , .A1( us20_n718 ) , .ZN( us20_n719 ) );
  AOI221_X1 us20_U123 (.A( us20_n710 ) , .ZN( us20_n721 ) , .C2( us20_n844 ) , .B2( us20_n845 ) , .C1( us20_n861 ) , .B1( us20_n862 ) );
  NAND4_X1 us20_U124 (.A4( us20_n573 ) , .A3( us20_n574 ) , .A1( us20_n575 ) , .ZN( us20_n723 ) , .A2( us20_n874 ) );
  NOR4_X1 us20_U125 (.A4( us20_n569 ) , .A3( us20_n570 ) , .A2( us20_n571 ) , .A1( us20_n572 ) , .ZN( us20_n573 ) );
  AOI221_X1 us20_U126 (.A( us20_n564 ) , .C2( us20_n565 ) , .ZN( us20_n574 ) , .B2( us20_n845 ) , .B1( us20_n852 ) , .C1( us20_n853 ) );
  NOR2_X1 us20_U127 (.ZN( us20_n575 ) , .A1( us20_n622 ) , .A2( us20_n745 ) );
  NAND4_X1 us20_U128 (.A4( us20_n633 ) , .A3( us20_n634 ) , .A2( us20_n635 ) , .A1( us20_n636 ) , .ZN( us20_n743 ) );
  AOI211_X1 us20_U129 (.B( us20_n623 ) , .A( us20_n624 ) , .ZN( us20_n635 ) , .C2( us20_n836 ) , .C1( us20_n863 ) );
  NOR4_X1 us20_U13 (.A4( us20_n445 ) , .A3( us20_n446 ) , .A2( us20_n516 ) , .A1( us20_n541 ) , .ZN( us20_n706 ) );
  NOR4_X1 us20_U130 (.A4( us20_n629 ) , .A3( us20_n630 ) , .A2( us20_n631 ) , .A1( us20_n632 ) , .ZN( us20_n633 ) );
  NOR4_X1 us20_U131 (.A4( us20_n626 ) , .A3( us20_n627 ) , .A2( us20_n628 ) , .ZN( us20_n634 ) , .A1( us20_n664 ) );
  NAND4_X1 us20_U132 (.A4( us20_n493 ) , .A3( us20_n494 ) , .A1( us20_n495 ) , .ZN( us20_n802 ) , .A2( us20_n867 ) );
  AOI221_X1 us20_U133 (.A( us20_n489 ) , .ZN( us20_n494 ) , .B2( us20_n836 ) , .C2( us20_n841 ) , .C1( us20_n851 ) , .B1( us20_n860 ) );
  INV_X1 us20_U134 (.A( us20_n778 ) , .ZN( us20_n867 ) );
  NOR4_X1 us20_U135 (.A2( us20_n491 ) , .A1( us20_n492 ) , .ZN( us20_n493 ) , .A3( us20_n580 ) , .A4( us20_n612 ) );
  INV_X1 us20_U136 (.A( us20_n762 ) , .ZN( us20_n830 ) );
  OR4_X1 us20_U137 (.A4( us20_n580 ) , .A3( us20_n581 ) , .A2( us20_n582 ) , .A1( us20_n583 ) , .ZN( us20_n584 ) );
  OR4_X1 us20_U138 (.A4( us20_n566 ) , .A3( us20_n567 ) , .A2( us20_n568 ) , .ZN( us20_n572 ) , .A1( us20_n665 ) );
  OR4_X1 us20_U139 (.A4( us20_n682 ) , .A3( us20_n683 ) , .A2( us20_n684 ) , .A1( us20_n685 ) , .ZN( us20_n690 ) );
  OR3_X1 us20_U14 (.ZN( us20_n446 ) , .A1( us20_n528 ) , .A3( us20_n577 ) , .A2( us20_n875 ) );
  OR4_X1 us20_U140 (.ZN( us20_n466 ) , .A4( us20_n518 ) , .A3( us20_n529 ) , .A2( us20_n578 ) , .A1( us20_n712 ) );
  OR4_X1 us20_U141 (.A4( us20_n518 ) , .A2( us20_n519 ) , .A1( us20_n520 ) , .ZN( us20_n522 ) , .A3( us20_n821 ) );
  OR4_X1 us20_U142 (.ZN( us20_n492 ) , .A4( us20_n534 ) , .A2( us20_n547 ) , .A1( us20_n559 ) , .A3( us20_n632 ) );
  NAND2_X1 us20_U143 (.ZN( us20_n613 ) , .A2( us20_n837 ) , .A1( us20_n873 ) );
  OR3_X1 us20_U144 (.A3( us20_n506 ) , .A2( us20_n507 ) , .A1( us20_n508 ) , .ZN( us20_n511 ) );
  AOI221_X1 us20_U145 (.A( us20_n713 ) , .B2( us20_n714 ) , .ZN( us20_n720 ) , .C1( us20_n832 ) , .B1( us20_n839 ) , .C2( us20_n863 ) );
  OR2_X1 us20_U146 (.A2( us20_n711 ) , .A1( us20_n712 ) , .ZN( us20_n713 ) );
  INV_X1 us20_U147 (.A( us20_n463 ) , .ZN( us20_n864 ) );
  OAI21_X1 us20_U148 (.ZN( us20_n463 ) , .B1( us20_n809 ) , .A( us20_n834 ) , .B2( us20_n851 ) );
  INV_X1 us20_U149 (.A( us20_n754 ) , .ZN( us20_n869 ) );
  OR4_X1 us20_U15 (.A4( us20_n442 ) , .A2( us20_n443 ) , .A1( us20_n444 ) , .ZN( us20_n445 ) , .A3( us20_n553 ) );
  OAI21_X1 us20_U150 (.B1( us20_n753 ) , .ZN( us20_n754 ) , .A( us20_n845 ) , .B2( us20_n868 ) );
  AOI222_X1 us20_U151 (.ZN( us20_n660 ) , .A2( us20_n839 ) , .B1( us20_n841 ) , .C2( us20_n845 ) , .A1( us20_n860 ) , .C1( us20_n863 ) , .B2( us20_n870 ) );
  INV_X1 us20_U152 (.A( us20_n647 ) , .ZN( us20_n870 ) );
  INV_X1 us20_U153 (.A( us20_n672 ) , .ZN( us20_n859 ) );
  AOI21_X1 us20_U154 (.A( us20_n670 ) , .B1( us20_n671 ) , .ZN( us20_n672 ) , .B2( us20_n856 ) );
  OAI22_X1 us20_U155 (.ZN( us20_n483 ) , .A1( us20_n708 ) , .B2( us20_n785 ) , .A2( us20_n806 ) , .B1( us20_n812 ) );
  OAI222_X1 us20_U156 (.B2( us20_n747 ) , .B1( us20_n748 ) , .A2( us20_n749 ) , .ZN( us20_n757 ) , .C2( us20_n805 ) , .C1( us20_n814 ) , .A1( us20_n817 ) );
  OAI222_X1 us20_U157 (.B2( us20_n708 ) , .ZN( us20_n709 ) , .C2( us20_n724 ) , .B1( us20_n747 ) , .A1( us20_n806 ) , .C1( us20_n814 ) , .A2( us20_n815 ) );
  OAI222_X1 us20_U158 (.ZN( us20_n505 ) , .C2( us20_n625 ) , .B2( us20_n647 ) , .B1( us20_n747 ) , .A2( us20_n748 ) , .C1( us20_n805 ) , .A1( us20_n806 ) );
  NAND2_X1 us20_U159 (.A1( us20_n447 ) , .A2( us20_n465 ) , .ZN( us20_n749 ) );
  INV_X1 us20_U16 (.A( us20_n613 ) , .ZN( us20_n875 ) );
  AOI22_X1 us20_U160 (.ZN( us20_n696 ) , .A1( us20_n830 ) , .B2( us20_n843 ) , .A2( us20_n865 ) , .B1( us20_n868 ) );
  AOI22_X1 us20_U161 (.A2( us20_n782 ) , .ZN( us20_n783 ) , .B2( us20_n831 ) , .A1( us20_n834 ) , .B1( us20_n863 ) );
  INV_X1 us20_U162 (.A( us20_n730 ) , .ZN( us20_n839 ) );
  INV_X1 us20_U163 (.A( us20_n790 ) , .ZN( us20_n832 ) );
  NAND2_X1 us20_U164 (.A1( us20_n451 ) , .A2( us20_n453 ) , .ZN( us20_n762 ) );
  AOI211_X1 us20_U165 (.A( us20_n637 ) , .ZN( us20_n645 ) , .B( us20_n743 ) , .C2( us20_n839 ) , .C1( us20_n854 ) );
  OAI22_X1 us20_U166 (.ZN( us20_n637 ) , .A1( us20_n699 ) , .B2( us20_n728 ) , .A2( us20_n762 ) , .B1( us20_n816 ) );
  OAI221_X1 us20_U167 (.A( us20_n727 ) , .C2( us20_n728 ) , .B2( us20_n729 ) , .B1( us20_n730 ) , .ZN( us20_n737 ) , .C1( us20_n817 ) );
  AOI22_X1 us20_U168 (.ZN( us20_n727 ) , .B1( us20_n832 ) , .A2( us20_n838 ) , .A1( us20_n863 ) , .B2( us20_n866 ) );
  OAI22_X1 us20_U169 (.ZN( us20_n489 ) , .A1( us20_n724 ) , .B2( us20_n728 ) , .B1( us20_n730 ) , .A2( us20_n779 ) );
  INV_X1 us20_U17 (.A( us20_n749 ) , .ZN( us20_n863 ) );
  OAI22_X1 us20_U170 (.ZN( us20_n624 ) , .B1( us20_n669 ) , .B2( us20_n747 ) , .A1( us20_n815 ) , .A2( us20_n816 ) );
  OAI22_X1 us20_U171 (.B2( us20_n779 ) , .B1( us20_n780 ) , .ZN( us20_n781 ) , .A2( us20_n814 ) , .A1( us20_n815 ) );
  OAI22_X1 us20_U172 (.A1( us20_n724 ) , .ZN( us20_n726 ) , .B2( us20_n750 ) , .B1( us20_n812 ) , .A2( us20_n816 ) );
  OAI22_X1 us20_U173 (.B2( us20_n744 ) , .ZN( us20_n746 ) , .A2( us20_n762 ) , .B1( us20_n780 ) , .A1( us20_n792 ) );
  OAI22_X1 us20_U174 (.ZN( us20_n496 ) , .A2( us20_n744 ) , .A1( us20_n780 ) , .B1( us20_n791 ) , .B2( us20_n806 ) );
  OAI22_X1 us20_U175 (.B2( us20_n803 ) , .B1( us20_n804 ) , .A2( us20_n805 ) , .A1( us20_n806 ) , .ZN( us20_n808 ) );
  INV_X1 us20_U176 (.A( us20_n788 ) , .ZN( us20_n845 ) );
  INV_X1 us20_U177 (.A( us20_n744 ) , .ZN( us20_n837 ) );
  INV_X1 us20_U178 (.A( us20_n814 ) , .ZN( us20_n833 ) );
  OAI22_X1 us20_U179 (.B1( us20_n490 ) , .ZN( us20_n491 ) , .A1( us20_n686 ) , .A2( us20_n763 ) , .B2( us20_n817 ) );
  AOI222_X1 us20_U18 (.ZN( us20_n563 ) , .B1( us20_n830 ) , .C1( us20_n841 ) , .A2( us20_n843 ) , .A1( us20_n854 ) , .B2( us20_n863 ) , .C2( us20_n873 ) );
  NOR3_X1 us20_U180 (.ZN( us20_n490 ) , .A1( us20_n782 ) , .A2( us20_n850 ) , .A3( us20_n863 ) );
  OAI22_X1 us20_U181 (.ZN( us20_n695 ) , .A2( us20_n730 ) , .A1( us20_n780 ) , .B1( us20_n791 ) , .B2( us20_n817 ) );
  INV_X1 us20_U182 (.A( us20_n805 ) , .ZN( us20_n860 ) );
  INV_X1 us20_U183 (.A( us20_n669 ) , .ZN( us20_n865 ) );
  NOR2_X1 us20_U184 (.ZN( us20_n715 ) , .A1( us20_n805 ) , .A2( us20_n817 ) );
  NOR2_X1 us20_U185 (.ZN( us20_n666 ) , .A1( us20_n728 ) , .A2( us20_n803 ) );
  NOR2_X1 us20_U186 (.ZN( us20_n546 ) , .A2( us20_n780 ) , .A1( us20_n814 ) );
  NOR2_X1 us20_U187 (.ZN( us20_n577 ) , .A2( us20_n699 ) , .A1( us20_n814 ) );
  NOR2_X1 us20_U188 (.ZN( us20_n570 ) , .A1( us20_n728 ) , .A2( us20_n806 ) );
  NOR2_X1 us20_U189 (.A2( us20_n744 ) , .ZN( us20_n755 ) , .A1( us20_n805 ) );
  NOR4_X1 us20_U19 (.ZN( us20_n473 ) , .A2( us20_n521 ) , .A4( us20_n594 ) , .A1( us20_n609 ) , .A3( us20_n629 ) );
  NOR2_X1 us20_U190 (.ZN( us20_n718 ) , .A2( us20_n724 ) , .A1( us20_n744 ) );
  NOR2_X1 us20_U191 (.ZN( us20_n735 ) , .A2( us20_n803 ) , .A1( us20_n805 ) );
  INV_X1 us20_U192 (.A( us20_n750 ) , .ZN( us20_n842 ) );
  NOR2_X1 us20_U193 (.ZN( us20_n532 ) , .A2( us20_n749 ) , .A1( us20_n750 ) );
  NOR2_X1 us20_U194 (.ZN( us20_n654 ) , .A1( us20_n728 ) , .A2( us20_n813 ) );
  NOR2_X1 us20_U195 (.ZN( us20_n615 ) , .A1( us20_n785 ) , .A2( us20_n815 ) );
  NOR2_X1 us20_U196 (.ZN( us20_n629 ) , .A2( us20_n728 ) , .A1( us20_n785 ) );
  NOR2_X1 us20_U197 (.ZN( us20_n628 ) , .A2( us20_n669 ) , .A1( us20_n785 ) );
  NOR2_X1 us20_U198 (.ZN( us20_n611 ) , .A2( us20_n780 ) , .A1( us20_n806 ) );
  INV_X1 us20_U199 (.A( us20_n747 ) , .ZN( us20_n834 ) );
  NOR4_X1 us20_U20 (.A4( us20_n544 ) , .A3( us20_n545 ) , .A2( us20_n546 ) , .A1( us20_n547 ) , .ZN( us20_n548 ) );
  NOR2_X1 us20_U200 (.ZN( us20_n601 ) , .A2( us20_n780 ) , .A1( us20_n803 ) );
  NOR2_X1 us20_U201 (.A2( us20_n708 ) , .A1( us20_n750 ) , .ZN( us20_n771 ) );
  NOR2_X1 us20_U202 (.ZN( us20_n652 ) , .A1( us20_n669 ) , .A2( us20_n814 ) );
  INV_X1 us20_U203 (.A( us20_n792 ) , .ZN( us20_n851 ) );
  NOR2_X1 us20_U204 (.A1( us20_n669 ) , .ZN( us20_n673 ) , .A2( us20_n744 ) );
  NOR2_X1 us20_U205 (.ZN( us20_n602 ) , .A1( us20_n669 ) , .A2( us20_n803 ) );
  NOR2_X1 us20_U206 (.A1( us20_n669 ) , .ZN( us20_n688 ) , .A2( us20_n816 ) );
  NOR2_X1 us20_U207 (.ZN( us20_n667 ) , .A1( us20_n750 ) , .A2( us20_n815 ) );
  NOR2_X1 us20_U208 (.A2( us20_n744 ) , .ZN( us20_n769 ) , .A1( us20_n812 ) );
  NOR2_X1 us20_U209 (.ZN( us20_n555 ) , .A1( us20_n750 ) , .A2( us20_n791 ) );
  NOR4_X1 us20_U21 (.ZN( us20_n479 ) , .A1( us20_n520 ) , .A4( us20_n557 ) , .A3( us20_n582 ) , .A2( us20_n630 ) );
  NOR2_X1 us20_U210 (.ZN( us20_n528 ) , .A2( us20_n724 ) , .A1( us20_n803 ) );
  NOR2_X1 us20_U211 (.ZN( us20_n508 ) , .A2( us20_n780 ) , .A1( us20_n785 ) );
  NOR2_X1 us20_U212 (.ZN( us20_n543 ) , .A2( us20_n708 ) , .A1( us20_n785 ) );
  NOR2_X1 us20_U213 (.ZN( us20_n531 ) , .A2( us20_n780 ) , .A1( us20_n816 ) );
  NOR2_X1 us20_U214 (.ZN( us20_n664 ) , .A1( us20_n785 ) , .A2( us20_n791 ) );
  NOR2_X1 us20_U215 (.ZN( us20_n599 ) , .A2( us20_n791 ) , .A1( us20_n816 ) );
  NOR2_X1 us20_U216 (.A1( us20_n669 ) , .ZN( us20_n766 ) , .A2( us20_n813 ) );
  NOR2_X1 us20_U217 (.A1( us20_n699 ) , .ZN( us20_n768 ) , .A2( us20_n813 ) );
  NOR2_X1 us20_U218 (.ZN( us20_n527 ) , .A1( us20_n669 ) , .A2( us20_n779 ) );
  OAI22_X1 us20_U219 (.B1( us20_n440 ) , .ZN( us20_n444 ) , .A2( us20_n728 ) , .A1( us20_n744 ) , .B2( us20_n749 ) );
  NOR4_X1 us20_U22 (.A4( us20_n532 ) , .A3( us20_n533 ) , .A2( us20_n534 ) , .ZN( us20_n535 ) , .A1( us20_n820 ) );
  NOR3_X1 us20_U220 (.ZN( us20_n440 ) , .A2( us20_n836 ) , .A3( us20_n837 ) , .A1( us20_n846 ) );
  OAI22_X1 us20_U221 (.ZN( us20_n710 ) , .A2( us20_n728 ) , .B2( us20_n729 ) , .A1( us20_n744 ) , .B1( us20_n813 ) );
  NOR2_X1 us20_U222 (.ZN( us20_n557 ) , .A1( us20_n792 ) , .A2( us20_n814 ) );
  NOR2_X1 us20_U223 (.ZN( us20_n545 ) , .A1( us20_n749 ) , .A2( us20_n814 ) );
  NOR2_X1 us20_U224 (.ZN( us20_n556 ) , .A1( us20_n762 ) , .A2( us20_n805 ) );
  NOR2_X1 us20_U225 (.ZN( us20_n661 ) , .A1( us20_n729 ) , .A2( us20_n790 ) );
  NOR2_X1 us20_U226 (.ZN( us20_n507 ) , .A1( us20_n812 ) , .A2( us20_n817 ) );
  INV_X1 us20_U227 (.A( us20_n806 ) , .ZN( us20_n841 ) );
  NOR2_X1 us20_U228 (.ZN( us20_n509 ) , .A1( us20_n729 ) , .A2( us20_n779 ) );
  NOR2_X1 us20_U229 (.ZN( us20_n544 ) , .A2( us20_n785 ) , .A1( us20_n792 ) );
  NOR4_X1 us20_U23 (.ZN( us20_n456 ) , .A2( us20_n517 ) , .A1( us20_n543 ) , .A3( us20_n579 ) , .A4( us20_n615 ) );
  OAI22_X1 us20_U230 (.B2( us20_n750 ) , .B1( us20_n751 ) , .A1( us20_n752 ) , .ZN( us20_n756 ) , .A2( us20_n806 ) );
  NOR2_X1 us20_U231 (.ZN( us20_n751 ) , .A2( us20_n852 ) , .A1( us20_n860 ) );
  NOR3_X1 us20_U232 (.ZN( us20_n752 ) , .A2( us20_n853 ) , .A1( us20_n863 ) , .A3( us20_n865 ) );
  NOR2_X1 us20_U233 (.ZN( us20_n530 ) , .A2( us20_n744 ) , .A1( us20_n792 ) );
  NOR2_X1 us20_U234 (.ZN( us20_n663 ) , .A1( us20_n729 ) , .A2( us20_n785 ) );
  INV_X1 us20_U235 (.A( us20_n728 ) , .ZN( us20_n852 ) );
  NOR2_X1 us20_U236 (.A1( us20_n749 ) , .ZN( us20_n767 ) , .A2( us20_n803 ) );
  NOR2_X1 us20_U237 (.ZN( us20_n506 ) , .A2( us20_n728 ) , .A1( us20_n762 ) );
  NOR2_X1 us20_U238 (.ZN( us20_n516 ) , .A1( us20_n708 ) , .A2( us20_n744 ) );
  NOR2_X1 us20_U239 (.ZN( us20_n614 ) , .A1( us20_n762 ) , .A2( us20_n812 ) );
  NOR2_X1 us20_U24 (.ZN( us20_n680 ) , .A2( us20_n834 ) , .A1( us20_n839 ) );
  NOR2_X1 us20_U240 (.ZN( us20_n670 ) , .A1( us20_n790 ) , .A2( us20_n805 ) );
  NOR2_X1 us20_U241 (.ZN( us20_n517 ) , .A1( us20_n708 ) , .A2( us20_n803 ) );
  NOR2_X1 us20_U242 (.ZN( us20_n558 ) , .A1( us20_n708 ) , .A2( us20_n816 ) );
  NOR2_X1 us20_U243 (.ZN( us20_n630 ) , .A1( us20_n747 ) , .A2( us20_n815 ) );
  NOR2_X1 us20_U244 (.ZN( us20_n655 ) , .A1( us20_n790 ) , .A2( us20_n815 ) );
  NOR2_X1 us20_U245 (.ZN( us20_n521 ) , .A1( us20_n790 ) , .A2( us20_n812 ) );
  NOR2_X1 us20_U246 (.ZN( us20_n668 ) , .A2( us20_n708 ) , .A1( us20_n790 ) );
  NOR2_X1 us20_U247 (.ZN( us20_n631 ) , .A1( us20_n724 ) , .A2( us20_n813 ) );
  NOR2_X1 us20_U248 (.ZN( us20_n656 ) , .A1( us20_n747 ) , .A2( us20_n780 ) );
  NOR2_X1 us20_U249 (.ZN( us20_n542 ) , .A1( us20_n762 ) , .A2( us20_n791 ) );
  NOR4_X1 us20_U25 (.ZN( us20_n620 ) , .A1( us20_n656 ) , .A3( us20_n666 ) , .A4( us20_n682 ) , .A2( us20_n766 ) );
  NOR2_X1 us20_U250 (.ZN( us20_n609 ) , .A2( us20_n724 ) , .A1( us20_n817 ) );
  AOI21_X1 us20_U251 (.B1( us20_n625 ) , .ZN( us20_n627 ) , .A( us20_n763 ) , .B2( us20_n814 ) );
  NOR2_X1 us20_U252 (.ZN( us20_n579 ) , .A2( us20_n708 ) , .A1( us20_n730 ) );
  NOR2_X1 us20_U253 (.ZN( us20_n533 ) , .A2( us20_n724 ) , .A1( us20_n730 ) );
  NOR2_X1 us20_U254 (.ZN( us20_n642 ) , .A2( us20_n788 ) , .A1( us20_n791 ) );
  NOR2_X1 us20_U255 (.A2( us20_n708 ) , .A1( us20_n762 ) , .ZN( us20_n794 ) );
  AOI21_X1 us20_U256 (.ZN( us20_n650 ) , .A( us20_n779 ) , .B1( us20_n792 ) , .B2( us20_n805 ) );
  AOI21_X1 us20_U257 (.A( us20_n815 ) , .B2( us20_n816 ) , .B1( us20_n817 ) , .ZN( us20_n818 ) );
  NOR2_X1 us20_U258 (.ZN( us20_n520 ) , .A2( us20_n708 ) , .A1( us20_n814 ) );
  NOR2_X1 us20_U259 (.ZN( us20_n582 ) , .A1( us20_n744 ) , .A2( us20_n815 ) );
  NOR4_X1 us20_U26 (.A4( us20_n609 ) , .A3( us20_n610 ) , .A2( us20_n611 ) , .A1( us20_n612 ) , .ZN( us20_n619 ) );
  AOI21_X1 us20_U260 (.ZN( us20_n515 ) , .A( us20_n729 ) , .B1( us20_n750 ) , .B2( us20_n803 ) );
  AOI21_X1 us20_U261 (.ZN( us20_n626 ) , .B2( us20_n669 ) , .A( us20_n790 ) , .B1( us20_n791 ) );
  AOI21_X1 us20_U262 (.ZN( us20_n499 ) , .B1( us20_n680 ) , .A( us20_n812 ) , .B2( us20_n816 ) );
  AOI21_X1 us20_U263 (.ZN( us20_n477 ) , .A( us20_n669 ) , .B1( us20_n750 ) , .B2( us20_n806 ) );
  NOR2_X1 us20_U264 (.ZN( us20_n559 ) , .A2( us20_n791 ) , .A1( us20_n803 ) );
  AOI21_X1 us20_U265 (.ZN( us20_n510 ) , .B2( us20_n669 ) , .A( us20_n730 ) , .B1( us20_n815 ) );
  NOR2_X1 us20_U266 (.ZN( us20_n519 ) , .A2( us20_n699 ) , .A1( us20_n816 ) );
  NOR2_X1 us20_U267 (.ZN( us20_n683 ) , .A2( us20_n699 ) , .A1( us20_n803 ) );
  NOR2_X1 us20_U268 (.ZN( us20_n581 ) , .A1( us20_n669 ) , .A2( us20_n788 ) );
  AOI21_X1 us20_U269 (.ZN( us20_n589 ) , .B2( us20_n699 ) , .B1( us20_n815 ) , .A( us20_n817 ) );
  NOR4_X1 us20_U27 (.A4( us20_n614 ) , .A3( us20_n615 ) , .A2( us20_n616 ) , .A1( us20_n617 ) , .ZN( us20_n618 ) );
  INV_X1 us20_U270 (.A( us20_n763 ) , .ZN( us20_n866 ) );
  AOI21_X1 us20_U271 (.ZN( us20_n498 ) , .A( us20_n724 ) , .B2( us20_n762 ) , .B1( us20_n814 ) );
  AOI21_X1 us20_U272 (.ZN( us20_n539 ) , .B2( us20_n812 ) , .A( us20_n814 ) , .B1( us20_n815 ) );
  AOI21_X1 us20_U273 (.ZN( us20_n540 ) , .A( us20_n763 ) , .B2( us20_n779 ) , .B1( us20_n817 ) );
  AOI21_X1 us20_U274 (.B1( us20_n699 ) , .ZN( us20_n700 ) , .A( us20_n732 ) , .B2( us20_n763 ) );
  AOI21_X1 us20_U275 (.ZN( us20_n591 ) , .B2( us20_n763 ) , .A( us20_n785 ) , .B1( us20_n812 ) );
  AOI21_X1 us20_U276 (.A( us20_n812 ) , .B2( us20_n813 ) , .B1( us20_n814 ) , .ZN( us20_n819 ) );
  INV_X1 us20_U277 (.A( us20_n791 ) , .ZN( us20_n873 ) );
  NOR2_X1 us20_U278 (.ZN( us20_n547 ) , .A1( us20_n699 ) , .A2( us20_n744 ) );
  INV_X1 us20_U279 (.A( us20_n729 ) , .ZN( us20_n868 ) );
  NOR4_X1 us20_U28 (.A4( us20_n514 ) , .A3( us20_n515 ) , .A2( us20_n516 ) , .A1( us20_n517 ) , .ZN( us20_n524 ) );
  AOI21_X1 us20_U280 (.ZN( us20_n569 ) , .B1( us20_n750 ) , .B2( us20_n762 ) , .A( us20_n780 ) );
  AOI21_X1 us20_U281 (.ZN( us20_n649 ) , .B1( us20_n729 ) , .B2( us20_n763 ) , .A( us20_n813 ) );
  NOR2_X1 us20_U282 (.ZN( us20_n685 ) , .A1( us20_n729 ) , .A2( us20_n816 ) );
  AOI21_X1 us20_U283 (.B1( us20_n686 ) , .ZN( us20_n687 ) , .A( us20_n728 ) , .B2( us20_n761 ) );
  AOI21_X1 us20_U284 (.ZN( us20_n640 ) , .B2( us20_n747 ) , .A( us20_n792 ) , .B1( us20_n803 ) );
  NOR2_X1 us20_U285 (.ZN( us20_n568 ) , .A1( us20_n729 ) , .A2( us20_n762 ) );
  AOI21_X1 us20_U286 (.ZN( us20_n593 ) , .B1( us20_n750 ) , .A( us20_n792 ) , .B2( us20_n813 ) );
  AOI21_X1 us20_U287 (.ZN( us20_n514 ) , .A( us20_n779 ) , .B2( us20_n792 ) , .B1( us20_n812 ) );
  INV_X1 us20_U288 (.A( us20_n699 ) , .ZN( us20_n853 ) );
  AOI21_X1 us20_U289 (.ZN( us20_n450 ) , .B2( us20_n792 ) , .A( us20_n803 ) , .B1( us20_n815 ) );
  AOI222_X1 us20_U29 (.ZN( us20_n525 ) , .A1( us20_n834 ) , .B2( us20_n837 ) , .C1( us20_n844 ) , .C2( us20_n850 ) , .A2( us20_n852 ) , .B1( us20_n866 ) );
  AOI21_X1 us20_U290 (.ZN( us20_n639 ) , .B2( us20_n749 ) , .A( us20_n788 ) , .B1( us20_n812 ) );
  AOI21_X1 us20_U291 (.ZN( us20_n564 ) , .B1( us20_n724 ) , .A( us20_n779 ) , .B2( us20_n791 ) );
  AOI21_X1 us20_U292 (.ZN( us20_n689 ) , .B2( us20_n749 ) , .B1( us20_n763 ) , .A( us20_n806 ) );
  NOR2_X1 us20_U293 (.ZN( us20_n529 ) , .A1( us20_n708 ) , .A2( us20_n779 ) );
  NOR2_X1 us20_U294 (.ZN( us20_n567 ) , .A1( us20_n747 ) , .A2( us20_n805 ) );
  AOI21_X1 us20_U295 (.A( us20_n790 ) , .B2( us20_n791 ) , .B1( us20_n792 ) , .ZN( us20_n793 ) );
  AOI21_X1 us20_U296 (.A( us20_n733 ) , .ZN( us20_n734 ) , .B2( us20_n780 ) , .B1( us20_n792 ) );
  NOR2_X1 us20_U297 (.A2( us20_n813 ) , .A1( us20_n815 ) , .ZN( us20_n821 ) );
  AOI21_X1 us20_U298 (.ZN( us20_n641 ) , .B1( us20_n680 ) , .A( us20_n791 ) , .B2( us20_n817 ) );
  NOR2_X1 us20_U299 (.ZN( us20_n578 ) , .A1( us20_n708 ) , .A2( us20_n813 ) );
  NAND4_X1 us20_U3 (.ZN( sa22_sr_2 ) , .A4( us20_n643 ) , .A3( us20_n644 ) , .A2( us20_n645 ) , .A1( us20_n646 ) );
  NOR4_X1 us20_U30 (.A3( us20_n521 ) , .A1( us20_n522 ) , .ZN( us20_n523 ) , .A2( us20_n673 ) , .A4( us20_n769 ) );
  NOR2_X1 us20_U300 (.ZN( us20_n665 ) , .A1( us20_n780 ) , .A2( us20_n813 ) );
  NOR2_X1 us20_U301 (.ZN( us20_n711 ) , .A1( us20_n762 ) , .A2( us20_n763 ) );
  NOR2_X1 us20_U302 (.ZN( us20_n583 ) , .A1( us20_n792 ) , .A2( us20_n817 ) );
  NOR2_X1 us20_U303 (.ZN( us20_n682 ) , .A2( us20_n708 ) , .A1( us20_n817 ) );
  NOR2_X1 us20_U304 (.ZN( us20_n534 ) , .A1( us20_n724 ) , .A2( us20_n788 ) );
  NOR2_X1 us20_U305 (.ZN( us20_n684 ) , .A1( us20_n791 ) , .A2( us20_n813 ) );
  NAND2_X1 us20_U306 (.ZN( us20_n753 ) , .A1( us20_n763 ) , .A2( us20_n805 ) );
  INV_X1 us20_U307 (.A( us20_n815 ) , .ZN( us20_n855 ) );
  AOI21_X1 us20_U308 (.ZN( us20_n442 ) , .A( us20_n699 ) , .B1( us20_n733 ) , .B2( us20_n750 ) );
  OAI21_X1 us20_U309 (.A( us20_n731 ) , .B1( us20_n732 ) , .ZN( us20_n736 ) , .B2( us20_n805 ) );
  AOI221_X1 us20_U31 (.A( us20_n781 ) , .ZN( us20_n798 ) , .C2( us20_n837 ) , .B2( us20_n838 ) , .B1( us20_n865 ) , .C1( us20_n866 ) );
  OAI21_X1 us20_U310 (.ZN( us20_n731 ) , .A( us20_n833 ) , .B2( us20_n852 ) , .B1( us20_n873 ) );
  INV_X1 us20_U311 (.A( us20_n780 ) , .ZN( us20_n850 ) );
  AOI21_X1 us20_U312 (.ZN( us20_n443 ) , .B1( us20_n789 ) , .B2( us20_n791 ) , .A( us20_n814 ) );
  NAND2_X1 us20_U313 (.ZN( us20_n714 ) , .A1( us20_n728 ) , .A2( us20_n780 ) );
  NAND2_X1 us20_U314 (.A2( us20_n762 ) , .A1( us20_n806 ) , .ZN( us20_n810 ) );
  INV_X1 us20_U315 (.A( us20_n785 ) , .ZN( us20_n846 ) );
  NOR2_X1 us20_U316 (.ZN( us20_n484 ) , .A1( us20_n788 ) , .A2( us20_n805 ) );
  AOI21_X1 us20_U317 (.ZN( us20_n497 ) , .A( us20_n779 ) , .B2( us20_n791 ) , .B1( us20_n804 ) );
  NOR2_X1 us20_U318 (.ZN( us20_n470 ) , .A2( us20_n779 ) , .A1( us20_n815 ) );
  NOR2_X1 us20_U319 (.ZN( us20_n712 ) , .A2( us20_n724 ) , .A1( us20_n790 ) );
  NOR4_X1 us20_U32 (.A4( us20_n793 ) , .A3( us20_n794 ) , .A2( us20_n795 ) , .A1( us20_n796 ) , .ZN( us20_n797 ) );
  NOR2_X1 us20_U320 (.ZN( us20_n526 ) , .A1( us20_n724 ) , .A2( us20_n750 ) );
  OAI21_X1 us20_U321 (.A( us20_n787 ) , .B2( us20_n788 ) , .B1( us20_n789 ) , .ZN( us20_n795 ) );
  OAI21_X1 us20_U322 (.ZN( us20_n787 ) , .A( us20_n839 ) , .B1( us20_n863 ) , .B2( us20_n873 ) );
  NAND2_X1 us20_U323 (.A1( us20_n699 ) , .A2( us20_n729 ) , .ZN( us20_n782 ) );
  NOR2_X1 us20_U324 (.ZN( us20_n518 ) , .A1( us20_n708 ) , .A2( us20_n788 ) );
  INV_X1 us20_U325 (.A( us20_n813 ) , .ZN( us20_n836 ) );
  NAND2_X1 us20_U326 (.ZN( us20_n671 ) , .A1( us20_n806 ) , .A2( us20_n816 ) );
  OAI21_X1 us20_U327 (.A( us20_n698 ) , .ZN( us20_n702 ) , .B2( us20_n750 ) , .B1( us20_n804 ) );
  OAI21_X1 us20_U328 (.ZN( us20_n698 ) , .B2( us20_n833 ) , .B1( us20_n838 ) , .A( us20_n860 ) );
  INV_X1 us20_U329 (.A( us20_n724 ) , .ZN( us20_n856 ) );
  NOR4_X1 us20_U33 (.A4( us20_n776 ) , .A3( us20_n777 ) , .A1( us20_n778 ) , .ZN( us20_n799 ) , .A2( us20_n801 ) );
  INV_X1 us20_U330 (.A( us20_n817 ) , .ZN( us20_n844 ) );
  AND2_X1 us20_U331 (.ZN( us20_n732 ) , .A1( us20_n779 ) , .A2( us20_n785 ) );
  OAI222_X1 us20_U332 (.ZN( us20_n617 ) , .B1( us20_n697 ) , .C1( us20_n724 ) , .C2( us20_n747 ) , .B2( us20_n786 ) , .A2( us20_n792 ) , .A1( us20_n816 ) );
  AOI221_X1 us20_U333 (.A( us20_n764 ) , .ZN( us20_n774 ) , .C2( us20_n810 ) , .B2( us20_n835 ) , .C1( us20_n855 ) , .B1( us20_n866 ) );
  AOI21_X1 us20_U334 (.B2( us20_n763 ) , .ZN( us20_n764 ) , .A( us20_n788 ) , .B1( us20_n792 ) );
  INV_X1 us20_U335 (.A( us20_n761 ) , .ZN( us20_n835 ) );
  NAND2_X1 us20_U336 (.A1( us20_n451 ) , .A2( us20_n454 ) , .ZN( us20_n814 ) );
  NAND2_X1 us20_U337 (.A1( us20_n447 ) , .A2( us20_n449 ) , .ZN( us20_n805 ) );
  NAND2_X1 us20_U338 (.A1( us20_n455 ) , .A2( us20_n462 ) , .ZN( us20_n750 ) );
  NAND2_X1 us20_U339 (.A1( us20_n455 ) , .A2( us20_n471 ) , .ZN( us20_n803 ) );
  NOR4_X1 us20_U34 (.A4( us20_n734 ) , .A3( us20_n735 ) , .A2( us20_n736 ) , .A1( us20_n737 ) , .ZN( us20_n738 ) );
  NAND2_X1 us20_U340 (.A1( us20_n453 ) , .A2( us20_n461 ) , .ZN( us20_n744 ) );
  NAND2_X1 us20_U341 (.A1( us20_n452 ) , .A2( us20_n465 ) , .ZN( us20_n669 ) );
  NAND2_X1 us20_U342 (.A2( us20_n448 ) , .A1( us20_n460 ) , .ZN( us20_n728 ) );
  NAND2_X1 us20_U343 (.A2( us20_n453 ) , .A1( us20_n455 ) , .ZN( us20_n806 ) );
  NAND2_X1 us20_U344 (.A1( us20_n451 ) , .A2( us20_n471 ) , .ZN( us20_n816 ) );
  NAND2_X1 us20_U345 (.A1( us20_n453 ) , .A2( us20_n472 ) , .ZN( us20_n785 ) );
  NAND2_X1 us20_U346 (.A2( us20_n454 ) , .A1( us20_n472 ) , .ZN( us20_n779 ) );
  NAND2_X1 us20_U347 (.A2( us20_n464 ) , .A1( us20_n465 ) , .ZN( us20_n812 ) );
  NAND2_X1 us20_U348 (.A1( us20_n441 ) , .A2( us20_n460 ) , .ZN( us20_n699 ) );
  NAND2_X1 us20_U349 (.A2( us20_n449 ) , .A1( us20_n452 ) , .ZN( us20_n763 ) );
  AOI211_X1 us20_U35 (.B( us20_n725 ) , .A( us20_n726 ) , .ZN( us20_n739 ) , .C1( us20_n843 ) , .C2( us20_n855 ) );
  NAND2_X1 us20_U350 (.A2( us20_n448 ) , .A1( us20_n452 ) , .ZN( us20_n729 ) );
  NAND2_X1 us20_U351 (.A2( us20_n461 ) , .A1( us20_n462 ) , .ZN( us20_n747 ) );
  NAND2_X1 us20_U352 (.A1( us20_n462 ) , .A2( us20_n472 ) , .ZN( us20_n788 ) );
  NOR2_X1 us20_U353 (.ZN( us20_n465 ) , .A2( us20_n847 ) , .A1( us20_n848 ) );
  NOR2_X1 us20_U354 (.ZN( us20_n453 ) , .A1( us20_n826 ) , .A2( us20_n827 ) );
  NOR2_X1 us20_U355 (.ZN( us20_n451 ) , .A1( us20_n828 ) , .A2( us20_n829 ) );
  NAND2_X1 us20_U356 (.A2( us20_n461 ) , .A1( us20_n471 ) , .ZN( us20_n697 ) );
  NAND2_X1 us20_U357 (.A1( us20_n451 ) , .A2( us20_n462 ) , .ZN( us20_n790 ) );
  NAND2_X1 us20_U358 (.A2( us20_n441 ) , .A1( us20_n447 ) , .ZN( us20_n784 ) );
  NAND2_X2 us20_U359 (.A2( us20_n448 ) , .A1( us20_n464 ) , .ZN( us20_n815 ) );
  NOR3_X1 us20_U36 (.A3( us20_n722 ) , .A1( us20_n723 ) , .ZN( us20_n740 ) , .A2( us20_n741 ) );
  NAND2_X1 us20_U360 (.A2( us20_n454 ) , .A1( us20_n455 ) , .ZN( us20_n730 ) );
  NAND2_X2 us20_U361 (.A2( us20_n441 ) , .A1( us20_n452 ) , .ZN( us20_n791 ) );
  NAND2_X2 us20_U362 (.A1( us20_n449 ) , .A2( us20_n464 ) , .ZN( us20_n724 ) );
  NAND2_X2 us20_U363 (.A1( us20_n449 ) , .A2( us20_n460 ) , .ZN( us20_n792 ) );
  NAND2_X2 us20_U364 (.A1( us20_n441 ) , .A2( us20_n464 ) , .ZN( us20_n708 ) );
  NAND2_X2 us20_U365 (.A2( us20_n471 ) , .A1( us20_n472 ) , .ZN( us20_n817 ) );
  NAND2_X2 us20_U366 (.A2( us20_n460 ) , .A1( us20_n465 ) , .ZN( us20_n780 ) );
  NOR2_X1 us20_U367 (.ZN( us20_n447 ) , .A2( us20_n849 ) , .A1( us20_n858 ) );
  NAND2_X1 us20_U368 (.A1( us20_n447 ) , .A2( us20_n448 ) , .ZN( us20_n786 ) );
  NOR2_X1 us20_U369 (.A2( sa20_6 ) , .A1( sa20_7 ) , .ZN( us20_n464 ) );
  NOR4_X1 us20_U37 (.A3( us20_n755 ) , .A2( us20_n756 ) , .A1( us20_n757 ) , .ZN( us20_n758 ) , .A4( us20_n869 ) );
  NOR2_X1 us20_U370 (.A2( sa20_7 ) , .ZN( us20_n460 ) , .A1( us20_n849 ) );
  NOR2_X1 us20_U371 (.A2( sa20_4 ) , .ZN( us20_n449 ) , .A1( us20_n848 ) );
  NOR2_X1 us20_U372 (.A2( sa20_4 ) , .A1( sa20_5 ) , .ZN( us20_n441 ) );
  NOR2_X1 us20_U373 (.A2( sa20_5 ) , .ZN( us20_n448 ) , .A1( us20_n847 ) );
  NOR2_X1 us20_U374 (.A2( sa20_1 ) , .ZN( us20_n471 ) , .A1( us20_n826 ) );
  NOR2_X1 us20_U375 (.A2( sa20_2 ) , .A1( sa20_3 ) , .ZN( us20_n472 ) );
  NOR2_X1 us20_U376 (.A2( sa20_6 ) , .ZN( us20_n452 ) , .A1( us20_n858 ) );
  NOR2_X1 us20_U377 (.A2( sa20_0 ) , .A1( sa20_1 ) , .ZN( us20_n462 ) );
  NOR2_X1 us20_U378 (.A2( sa20_3 ) , .ZN( us20_n455 ) , .A1( us20_n828 ) );
  NOR2_X1 us20_U379 (.A2( sa20_2 ) , .ZN( us20_n461 ) , .A1( us20_n829 ) );
  AOI211_X1 us20_U38 (.B( us20_n745 ) , .A( us20_n746 ) , .ZN( us20_n759 ) , .C1( us20_n832 ) , .C2( us20_n853 ) );
  NOR2_X1 us20_U380 (.A2( sa20_0 ) , .ZN( us20_n454 ) , .A1( us20_n827 ) );
  INV_X1 us20_U381 (.A( sa20_4 ) , .ZN( us20_n847 ) );
  INV_X1 us20_U382 (.A( sa20_6 ) , .ZN( us20_n849 ) );
  INV_X1 us20_U383 (.A( sa20_3 ) , .ZN( us20_n829 ) );
  INV_X1 us20_U384 (.A( sa20_1 ) , .ZN( us20_n827 ) );
  INV_X1 us20_U385 (.A( sa20_2 ) , .ZN( us20_n828 ) );
  INV_X1 us20_U386 (.A( sa20_0 ) , .ZN( us20_n826 ) );
  INV_X1 us20_U387 (.A( sa20_5 ) , .ZN( us20_n848 ) );
  INV_X1 us20_U388 (.A( sa20_7 ) , .ZN( us20_n858 ) );
  NAND2_X1 us20_U389 (.A1( us20_n729 ) , .A2( us20_n784 ) , .ZN( us20_n811 ) );
  NOR3_X1 us20_U39 (.A3( us20_n741 ) , .A2( us20_n742 ) , .A1( us20_n743 ) , .ZN( us20_n760 ) );
  OAI22_X1 us20_U390 (.ZN( us20_n588 ) , .A2( us20_n747 ) , .B2( us20_n762 ) , .A1( us20_n763 ) , .B1( us20_n784 ) );
  AOI21_X1 us20_U391 (.ZN( us20_n592 ) , .B1( us20_n728 ) , .B2( us20_n784 ) , .A( us20_n790 ) );
  AOI21_X1 us20_U392 (.ZN( us20_n648 ) , .A( us20_n762 ) , .B2( us20_n784 ) , .B1( us20_n792 ) );
  AOI21_X1 us20_U393 (.ZN( us20_n623 ) , .B1( us20_n699 ) , .A( us20_n779 ) , .B2( us20_n784 ) );
  OAI22_X1 us20_U394 (.ZN( us20_n681 ) , .A1( us20_n699 ) , .A2( us20_n730 ) , .B2( us20_n784 ) , .B1( us20_n817 ) );
  OAI21_X1 us20_U395 (.A( us20_n613 ) , .ZN( us20_n616 ) , .B1( us20_n625 ) , .B2( us20_n784 ) );
  NOR2_X1 us20_U396 (.ZN( us20_n610 ) , .A1( us20_n784 ) , .A2( us20_n816 ) );
  OAI222_X1 us20_U397 (.A2( us20_n669 ) , .ZN( us20_n674 ) , .B1( us20_n747 ) , .B2( us20_n784 ) , .C2( us20_n788 ) , .C1( us20_n815 ) , .A1( us20_n817 ) );
  NOR2_X1 us20_U398 (.ZN( us20_n651 ) , .A1( us20_n784 ) , .A2( us20_n788 ) );
  NOR2_X1 us20_U399 (.ZN( us20_n553 ) , .A2( us20_n744 ) , .A1( us20_n784 ) );
  NOR3_X1 us20_U4 (.ZN( us20_n598 ) , .A1( us20_n608 ) , .A3( us20_n723 ) , .A2( us20_n742 ) );
  NOR2_X1 us20_U40 (.ZN( us20_n804 ) , .A1( us20_n854 ) , .A2( us20_n861 ) );
  INV_X1 us20_U400 (.A( us20_n784 ) , .ZN( us20_n861 ) );
  INV_X1 us20_U401 (.A( us20_n697 ) , .ZN( us20_n838 ) );
  NOR2_X1 us20_U402 (.A1( us20_n697 ) , .ZN( us20_n770 ) , .A2( us20_n815 ) );
  AOI21_X1 us20_U403 (.ZN( us20_n571 ) , .B2( us20_n697 ) , .B1( us20_n806 ) , .A( us20_n812 ) );
  NOR2_X1 us20_U404 (.ZN( us20_n632 ) , .A2( us20_n697 ) , .A1( us20_n724 ) );
  AOI21_X1 us20_U405 (.ZN( us20_n478 ) , .B2( us20_n697 ) , .A( us20_n749 ) , .B1( us20_n779 ) );
  NOR2_X1 us20_U406 (.ZN( us20_n662 ) , .A2( us20_n697 ) , .A1( us20_n729 ) );
  NOR2_X1 us20_U407 (.A2( us20_n697 ) , .A1( us20_n780 ) , .ZN( us20_n820 ) );
  NOR2_X1 us20_U408 (.ZN( us20_n600 ) , .A2( us20_n697 ) , .A1( us20_n784 ) );
  NOR2_X1 us20_U409 (.A2( us20_n697 ) , .ZN( us20_n716 ) , .A1( us20_n792 ) );
  NAND4_X1 us20_U41 (.ZN( sa22_sr_3 ) , .A4( us20_n704 ) , .A3( us20_n705 ) , .A2( us20_n706 ) , .A1( us20_n707 ) );
  NOR2_X1 us20_U410 (.ZN( us20_n566 ) , .A2( us20_n697 ) , .A1( us20_n763 ) );
  NOR2_X1 us20_U411 (.ZN( us20_n594 ) , .A2( us20_n697 ) , .A1( us20_n728 ) );
  AOI21_X1 us20_U412 (.ZN( us20_n552 ) , .B1( us20_n669 ) , .A( us20_n697 ) , .B2( us20_n805 ) );
  NOR2_X1 us20_U413 (.ZN( us20_n541 ) , .A2( us20_n697 ) , .A1( us20_n699 ) );
  NOR2_X1 us20_U414 (.ZN( us20_n580 ) , .A2( us20_n697 ) , .A1( us20_n791 ) );
  NAND2_X1 us20_U415 (.A1( us20_n454 ) , .A2( us20_n461 ) , .ZN( us20_n813 ) );
  AND2_X1 us20_U416 (.ZN( us20_n438 ) , .A2( us20_n831 ) , .A1( us20_n854 ) );
  AND2_X1 us20_U417 (.ZN( us20_n439 ) , .A2( us20_n843 ) , .A1( us20_n861 ) );
  NOR3_X1 us20_U418 (.A1( us20_n438 ) , .A2( us20_n439 ) , .A3( us20_n576 ) , .ZN( us20_n587 ) );
  INV_X1 us20_U419 (.A( us20_n812 ) , .ZN( us20_n854 ) );
  NOR4_X1 us20_U42 (.A4( us20_n700 ) , .A3( us20_n701 ) , .A2( us20_n702 ) , .A1( us20_n703 ) , .ZN( us20_n704 ) );
  INV_X1 us20_U420 (.A( us20_n816 ) , .ZN( us20_n831 ) );
  INV_X1 us20_U421 (.A( us20_n803 ) , .ZN( us20_n843 ) );
  AOI21_X1 us20_U422 (.ZN( us20_n576 ) , .B2( us20_n724 ) , .B1( us20_n748 ) , .A( us20_n785 ) );
  OAI221_X1 us20_U423 (.A( us20_n783 ) , .C2( us20_n784 ) , .B2( us20_n785 ) , .B1( us20_n786 ) , .ZN( us20_n796 ) , .C1( us20_n813 ) );
  AOI21_X1 us20_U424 (.ZN( us20_n500 ) , .A( us20_n697 ) , .B1( us20_n708 ) , .B2( us20_n786 ) );
  OAI221_X1 us20_U425 (.A( us20_n696 ) , .ZN( us20_n703 ) , .C2( us20_n784 ) , .C1( us20_n785 ) , .B1( us20_n786 ) , .B2( us20_n806 ) );
  OAI22_X1 us20_U426 (.ZN( us20_n590 ) , .B1( us20_n730 ) , .B2( us20_n749 ) , .A2( us20_n786 ) , .A1( us20_n803 ) );
  AOI222_X1 us20_U427 (.ZN( us20_n605 ) , .B2( us20_n671 ) , .B1( us20_n753 ) , .C2( us20_n831 ) , .A1( us20_n833 ) , .A2( us20_n862 ) , .C1( us20_n863 ) );
  AOI222_X1 us20_U428 (.ZN( us20_n513 ) , .C1( us20_n832 ) , .B2( us20_n837 ) , .A2( us20_n843 ) , .C2( us20_n862 ) , .B1( us20_n863 ) , .A1( us20_n866 ) );
  AOI221_X1 us20_U429 (.A( us20_n483 ) , .ZN( us20_n488 ) , .B1( us20_n831 ) , .C2( us20_n844 ) , .C1( us20_n852 ) , .B2( us20_n862 ) );
  AOI211_X1 us20_U43 (.B( us20_n694 ) , .A( us20_n695 ) , .ZN( us20_n705 ) , .C2( us20_n831 ) , .C1( us20_n851 ) );
  NAND2_X1 us20_U430 (.A2( us20_n749 ) , .A1( us20_n786 ) , .ZN( us20_n809 ) );
  NOR2_X1 us20_U431 (.ZN( us20_n612 ) , .A1( us20_n779 ) , .A2( us20_n786 ) );
  NOR2_X1 us20_U432 (.ZN( us20_n717 ) , .A2( us20_n744 ) , .A1( us20_n786 ) );
  NOR2_X1 us20_U433 (.ZN( us20_n653 ) , .A1( us20_n762 ) , .A2( us20_n786 ) );
  NOR2_X1 us20_U434 (.ZN( us20_n554 ) , .A1( us20_n786 ) , .A2( us20_n813 ) );
  NOR2_X1 us20_U435 (.ZN( us20_n789 ) , .A2( us20_n862 ) , .A1( us20_n868 ) );
  NOR2_X1 us20_U436 (.ZN( us20_n701 ) , .A2( us20_n786 ) , .A1( us20_n817 ) );
  NAND3_X1 us20_U437 (.ZN( sa22_sr_6 ) , .A3( us20_n797 ) , .A2( us20_n798 ) , .A1( us20_n799 ) );
  NAND3_X1 us20_U438 (.ZN( sa22_sr_5 ) , .A3( us20_n758 ) , .A2( us20_n759 ) , .A1( us20_n760 ) );
  NAND3_X1 us20_U439 (.ZN( sa22_sr_4 ) , .A3( us20_n738 ) , .A2( us20_n739 ) , .A1( us20_n740 ) );
  NOR2_X1 us20_U44 (.ZN( us20_n707 ) , .A2( us20_n776 ) , .A1( us20_n800 ) );
  NAND3_X1 us20_U440 (.A3( us20_n675 ) , .A2( us20_n676 ) , .A1( us20_n677 ) , .ZN( us20_n807 ) );
  NAND3_X1 us20_U441 (.ZN( us20_n638 ) , .A3( us20_n708 ) , .A2( us20_n724 ) , .A1( us20_n792 ) );
  NAND3_X1 us20_U442 (.A3( us20_n618 ) , .A2( us20_n619 ) , .A1( us20_n620 ) , .ZN( us20_n725 ) );
  NAND3_X1 us20_U443 (.A3( us20_n585 ) , .A2( us20_n586 ) , .A1( us20_n587 ) , .ZN( us20_n621 ) );
  NAND3_X1 us20_U444 (.ZN( us20_n565 ) , .A3( us20_n680 ) , .A2( us20_n750 ) , .A1( us20_n785 ) );
  NAND3_X1 us20_U445 (.A3( us20_n523 ) , .A2( us20_n524 ) , .A1( us20_n525 ) , .ZN( us20_n742 ) );
  NAND3_X1 us20_U446 (.A3( us20_n512 ) , .A1( us20_n513 ) , .ZN( us20_n608 ) , .A2( us20_n871 ) );
  NAND3_X1 us20_U447 (.A3( us20_n467 ) , .A2( us20_n468 ) , .A1( us20_n469 ) , .ZN( us20_n777 ) );
  NOR2_X1 us20_U448 (.A1( us20_n730 ) , .ZN( us20_n765 ) , .A2( us20_n786 ) );
  INV_X1 us20_U449 (.A( us20_n786 ) , .ZN( us20_n862 ) );
  NAND4_X1 us20_U45 (.ZN( sa22_sr_7 ) , .A4( us20_n822 ) , .A3( us20_n823 ) , .A2( us20_n824 ) , .A1( us20_n825 ) );
  NOR4_X1 us20_U46 (.A4( us20_n818 ) , .A3( us20_n819 ) , .A2( us20_n820 ) , .A1( us20_n821 ) , .ZN( us20_n822 ) );
  AOI222_X1 us20_U47 (.C2( us20_n809 ) , .B2( us20_n810 ) , .A2( us20_n811 ) , .ZN( us20_n823 ) , .C1( us20_n832 ) , .A1( us20_n839 ) , .B1( us20_n853 ) );
  AOI211_X1 us20_U48 (.B( us20_n807 ) , .A( us20_n808 ) , .ZN( us20_n824 ) , .C1( us20_n842 ) , .C2( us20_n850 ) );
  NAND4_X1 us20_U49 (.ZN( sa22_sr_0 ) , .A4( us20_n501 ) , .A3( us20_n502 ) , .A2( us20_n503 ) , .A1( us20_n504 ) );
  NOR3_X1 us20_U5 (.A3( us20_n800 ) , .A2( us20_n801 ) , .A1( us20_n802 ) , .ZN( us20_n825 ) );
  NOR4_X1 us20_U50 (.A4( us20_n498 ) , .A3( us20_n499 ) , .A2( us20_n500 ) , .ZN( us20_n501 ) , .A1( us20_n527 ) );
  AOI221_X1 us20_U51 (.A( us20_n497 ) , .ZN( us20_n502 ) , .B2( us20_n843 ) , .C1( us20_n846 ) , .C2( us20_n860 ) , .B1( us20_n862 ) );
  AOI211_X1 us20_U52 (.A( us20_n496 ) , .ZN( us20_n503 ) , .B( us20_n802 ) , .C2( us20_n839 ) , .C1( us20_n851 ) );
  NAND4_X1 us20_U53 (.ZN( sa22_sr_1 ) , .A4( us20_n595 ) , .A3( us20_n596 ) , .A2( us20_n597 ) , .A1( us20_n598 ) );
  NOR4_X1 us20_U54 (.A4( us20_n591 ) , .A3( us20_n592 ) , .A2( us20_n593 ) , .A1( us20_n594 ) , .ZN( us20_n595 ) );
  AOI211_X1 us20_U55 (.B( us20_n589 ) , .A( us20_n590 ) , .ZN( us20_n596 ) , .C2( us20_n811 ) , .C1( us20_n833 ) );
  AOI211_X1 us20_U56 (.A( us20_n588 ) , .ZN( us20_n597 ) , .B( us20_n621 ) , .C1( us20_n845 ) , .C2( us20_n855 ) );
  NOR2_X1 us20_U57 (.ZN( us20_n748 ) , .A1( us20_n861 ) , .A2( us20_n862 ) );
  NOR2_X1 us20_U58 (.ZN( us20_n625 ) , .A2( us20_n836 ) , .A1( us20_n839 ) );
  AOI222_X1 us20_U59 (.B2( us20_n638 ) , .ZN( us20_n644 ) , .B1( us20_n841 ) , .A1( us20_n842 ) , .C2( us20_n846 ) , .C1( us20_n863 ) , .A2( us20_n865 ) );
  NOR3_X1 us20_U6 (.A3( us20_n621 ) , .A2( us20_n622 ) , .ZN( us20_n636 ) , .A1( us20_n725 ) );
  NOR4_X1 us20_U60 (.A4( us20_n639 ) , .A3( us20_n640 ) , .A2( us20_n641 ) , .A1( us20_n642 ) , .ZN( us20_n643 ) );
  NOR3_X1 us20_U61 (.A2( us20_n607 ) , .A1( us20_n608 ) , .ZN( us20_n646 ) , .A3( us20_n722 ) );
  NAND4_X1 us20_U62 (.A4( us20_n603 ) , .A3( us20_n604 ) , .A2( us20_n605 ) , .A1( us20_n606 ) , .ZN( us20_n722 ) );
  NOR3_X1 us20_U63 (.A1( us20_n599 ) , .ZN( us20_n604 ) , .A3( us20_n663 ) , .A2( us20_n770 ) );
  NOR4_X1 us20_U64 (.A3( us20_n600 ) , .A2( us20_n601 ) , .A1( us20_n602 ) , .ZN( us20_n603 ) , .A4( us20_n655 ) );
  AOI222_X1 us20_U65 (.ZN( us20_n606 ) , .A1( us20_n830 ) , .C2( us20_n837 ) , .B1( us20_n842 ) , .A2( us20_n856 ) , .B2( us20_n861 ) , .C1( us20_n868 ) );
  AOI222_X1 us20_U66 (.ZN( us20_n469 ) , .B1( us20_n832 ) , .A1( us20_n839 ) , .C1( us20_n842 ) , .C2( us20_n851 ) , .A2( us20_n855 ) , .B2( us20_n865 ) );
  NOR4_X1 us20_U67 (.A1( us20_n466 ) , .ZN( us20_n467 ) , .A4( us20_n542 ) , .A2( us20_n554 ) , .A3( us20_n614 ) );
  AOI221_X1 us20_U68 (.ZN( us20_n468 ) , .C2( us20_n714 ) , .B2( us20_n831 ) , .C1( us20_n845 ) , .B1( us20_n860 ) , .A( us20_n864 ) );
  NAND4_X1 us20_U69 (.A4( us20_n485 ) , .A3( us20_n486 ) , .A2( us20_n487 ) , .A1( us20_n488 ) , .ZN( us20_n778 ) );
  NOR2_X1 us20_U7 (.ZN( us20_n495 ) , .A1( us20_n678 ) , .A2( us20_n694 ) );
  NOR4_X1 us20_U70 (.A4( us20_n484 ) , .ZN( us20_n487 ) , .A1( us20_n566 ) , .A2( us20_n581 ) , .A3( us20_n602 ) );
  NOR4_X1 us20_U71 (.ZN( us20_n486 ) , .A1( us20_n507 ) , .A2( us20_n519 ) , .A4( us20_n546 ) , .A3( us20_n611 ) );
  NOR4_X1 us20_U72 (.ZN( us20_n485 ) , .A2( us20_n533 ) , .A1( us20_n558 ) , .A3( us20_n631 ) , .A4( us20_n718 ) );
  NAND4_X1 us20_U73 (.A4( us20_n657 ) , .A3( us20_n658 ) , .A2( us20_n659 ) , .A1( us20_n660 ) , .ZN( us20_n800 ) );
  NOR3_X1 us20_U74 (.A3( us20_n648 ) , .A2( us20_n649 ) , .A1( us20_n650 ) , .ZN( us20_n659 ) );
  NOR3_X1 us20_U75 (.A3( us20_n651 ) , .A2( us20_n652 ) , .A1( us20_n653 ) , .ZN( us20_n658 ) );
  NOR3_X1 us20_U76 (.A3( us20_n654 ) , .A2( us20_n655 ) , .A1( us20_n656 ) , .ZN( us20_n657 ) );
  NAND4_X1 us20_U77 (.A4( us20_n560 ) , .A3( us20_n561 ) , .A2( us20_n562 ) , .A1( us20_n563 ) , .ZN( us20_n607 ) );
  NOR4_X1 us20_U78 (.A4( us20_n552 ) , .A3( us20_n553 ) , .A2( us20_n554 ) , .A1( us20_n555 ) , .ZN( us20_n562 ) );
  NOR4_X1 us20_U79 (.ZN( us20_n561 ) , .A1( us20_n653 ) , .A3( us20_n661 ) , .A4( us20_n685 ) , .A2( us20_n768 ) );
  NOR2_X1 us20_U8 (.A1( us20_n678 ) , .ZN( us20_n693 ) , .A2( us20_n807 ) );
  NOR4_X1 us20_U80 (.A4( us20_n556 ) , .A3( us20_n557 ) , .A2( us20_n558 ) , .A1( us20_n559 ) , .ZN( us20_n560 ) );
  NAND4_X1 us20_U81 (.A4( us20_n772 ) , .A3( us20_n773 ) , .A2( us20_n774 ) , .A1( us20_n775 ) , .ZN( us20_n801 ) );
  NOR3_X1 us20_U82 (.A3( us20_n765 ) , .A2( us20_n766 ) , .A1( us20_n767 ) , .ZN( us20_n773 ) );
  NOR4_X1 us20_U83 (.A4( us20_n768 ) , .A3( us20_n769 ) , .A2( us20_n770 ) , .A1( us20_n771 ) , .ZN( us20_n772 ) );
  AOI222_X1 us20_U84 (.ZN( us20_n775 ) , .A1( us20_n830 ) , .C1( us20_n834 ) , .B2( us20_n841 ) , .A2( us20_n850 ) , .B1( us20_n861 ) , .C2( us20_n873 ) );
  NOR4_X1 us20_U85 (.A4( us20_n509 ) , .A2( us20_n510 ) , .A1( us20_n511 ) , .ZN( us20_n512 ) , .A3( us20_n670 ) );
  INV_X1 us20_U86 (.A( us20_n505 ) , .ZN( us20_n871 ) );
  NOR4_X1 us20_U87 (.A4( us20_n661 ) , .A3( us20_n662 ) , .A2( us20_n663 ) , .A1( us20_n664 ) , .ZN( us20_n677 ) );
  NOR4_X1 us20_U88 (.A4( us20_n665 ) , .A3( us20_n666 ) , .A2( us20_n667 ) , .A1( us20_n668 ) , .ZN( us20_n676 ) );
  NOR4_X1 us20_U89 (.A3( us20_n673 ) , .A1( us20_n674 ) , .ZN( us20_n675 ) , .A4( us20_n715 ) , .A2( us20_n859 ) );
  NOR3_X1 us20_U9 (.ZN( us20_n504 ) , .A2( us20_n679 ) , .A3( us20_n777 ) , .A1( us20_n876 ) );
  NOR2_X1 us20_U90 (.ZN( us20_n761 ) , .A1( us20_n833 ) , .A2( us20_n834 ) );
  NOR2_X1 us20_U91 (.ZN( us20_n686 ) , .A1( us20_n831 ) , .A2( us20_n832 ) );
  NOR4_X1 us20_U92 (.A4( us20_n577 ) , .A3( us20_n578 ) , .A2( us20_n579 ) , .ZN( us20_n586 ) , .A1( us20_n683 ) );
  NOR4_X1 us20_U93 (.A1( us20_n584 ) , .ZN( us20_n585 ) , .A3( us20_n652 ) , .A2( us20_n662 ) , .A4( us20_n767 ) );
  NAND4_X1 us20_U94 (.A4( us20_n456 ) , .A3( us20_n457 ) , .A2( us20_n458 ) , .A1( us20_n459 ) , .ZN( us20_n679 ) );
  NOR3_X1 us20_U95 (.ZN( us20_n457 ) , .A3( us20_n530 ) , .A1( us20_n555 ) , .A2( us20_n570 ) );
  AOI221_X1 us20_U96 (.A( us20_n450 ) , .ZN( us20_n459 ) , .C2( us20_n753 ) , .B1( us20_n832 ) , .C1( us20_n842 ) , .B2( us20_n861 ) );
  NOR4_X1 us20_U97 (.ZN( us20_n458 ) , .A2( us20_n509 ) , .A1( us20_n599 ) , .A4( us20_n628 ) , .A3( us20_n711 ) );
  NAND4_X1 us20_U98 (.A4( us20_n535 ) , .A3( us20_n536 ) , .A2( us20_n537 ) , .A1( us20_n538 ) , .ZN( us20_n622 ) );
  NOR4_X1 us20_U99 (.A4( us20_n526 ) , .A2( us20_n527 ) , .A1( us20_n528 ) , .ZN( us20_n538 ) , .A3( us20_n701 ) );
  NOR2_X1 us32_U10 (.A1( us32_n678 ) , .ZN( us32_n693 ) , .A2( us32_n807 ) );
  AOI211_X1 us32_U100 (.B( us32_n477 ) , .A( us32_n478 ) , .ZN( us32_n482 ) , .C2( us32_n833 ) , .C1( us32_n861 ) );
  NOR4_X1 us32_U101 (.ZN( us32_n481 ) , .A3( us32_n532 ) , .A4( us32_n545 ) , .A2( us32_n567 ) , .A1( us32_n717 ) );
  NAND4_X1 us32_U102 (.A4( us32_n548 ) , .A3( us32_n549 ) , .A2( us32_n550 ) , .A1( us32_n551 ) , .ZN( us32_n745 ) );
  NOR3_X1 us32_U103 (.ZN( us32_n549 ) , .A2( us32_n651 ) , .A1( us32_n667 ) , .A3( us32_n771 ) );
  AOI211_X1 us32_U104 (.B( us32_n539 ) , .A( us32_n540 ) , .ZN( us32_n551 ) , .C2( us32_n839 ) , .C1( us32_n851 ) );
  NOR4_X1 us32_U105 (.A4( us32_n541 ) , .A3( us32_n542 ) , .A2( us32_n543 ) , .ZN( us32_n550 ) , .A1( us32_n688 ) );
  NOR4_X1 us32_U106 (.ZN( us32_n620 ) , .A1( us32_n656 ) , .A3( us32_n666 ) , .A4( us32_n682 ) , .A2( us32_n766 ) );
  NOR4_X1 us32_U107 (.A4( us32_n609 ) , .A3( us32_n610 ) , .A2( us32_n611 ) , .A1( us32_n612 ) , .ZN( us32_n619 ) );
  NOR4_X1 us32_U108 (.A4( us32_n614 ) , .A3( us32_n615 ) , .A2( us32_n616 ) , .A1( us32_n617 ) , .ZN( us32_n618 ) );
  NOR2_X1 us32_U109 (.ZN( us32_n686 ) , .A1( us32_n831 ) , .A2( us32_n832 ) );
  NOR3_X1 us32_U11 (.ZN( us32_n504 ) , .A2( us32_n679 ) , .A3( us32_n777 ) , .A1( us32_n876 ) );
  NAND4_X1 us32_U110 (.A4( us32_n485 ) , .A3( us32_n486 ) , .A2( us32_n487 ) , .A1( us32_n488 ) , .ZN( us32_n778 ) );
  NOR4_X1 us32_U111 (.A4( us32_n484 ) , .ZN( us32_n487 ) , .A1( us32_n566 ) , .A2( us32_n581 ) , .A3( us32_n602 ) );
  NOR4_X1 us32_U112 (.ZN( us32_n486 ) , .A1( us32_n507 ) , .A2( us32_n519 ) , .A4( us32_n546 ) , .A3( us32_n611 ) );
  NOR4_X1 us32_U113 (.ZN( us32_n485 ) , .A2( us32_n533 ) , .A1( us32_n558 ) , .A3( us32_n631 ) , .A4( us32_n718 ) );
  NAND4_X1 us32_U114 (.A4( us32_n691 ) , .A3( us32_n692 ) , .A1( us32_n693 ) , .ZN( us32_n776 ) , .A2( us32_n872 ) );
  AOI221_X1 us32_U115 (.A( us32_n681 ) , .ZN( us32_n692 ) , .B2( us32_n840 ) , .C1( us32_n842 ) , .C2( us32_n862 ) , .B1( us32_n865 ) );
  INV_X1 us32_U116 (.A( us32_n679 ) , .ZN( us32_n872 ) );
  NOR4_X1 us32_U117 (.A4( us32_n687 ) , .A3( us32_n688 ) , .A2( us32_n689 ) , .A1( us32_n690 ) , .ZN( us32_n691 ) );
  NAND4_X1 us32_U118 (.A4( us32_n473 ) , .A3( us32_n474 ) , .A2( us32_n475 ) , .A1( us32_n476 ) , .ZN( us32_n678 ) );
  NOR4_X1 us32_U119 (.ZN( us32_n475 ) , .A1( us32_n531 ) , .A3( us32_n568 ) , .A4( us32_n600 ) , .A2( us32_n642 ) );
  INV_X1 us32_U12 (.A( us32_n706 ) , .ZN( us32_n876 ) );
  NOR4_X1 us32_U120 (.A4( us32_n470 ) , .ZN( us32_n476 ) , .A3( us32_n556 ) , .A1( us32_n735 ) , .A2( us32_n755 ) );
  NOR4_X1 us32_U121 (.ZN( us32_n473 ) , .A2( us32_n521 ) , .A4( us32_n594 ) , .A1( us32_n609 ) , .A3( us32_n629 ) );
  NAND4_X1 us32_U122 (.A4( us32_n719 ) , .A3( us32_n720 ) , .A2( us32_n721 ) , .ZN( us32_n741 ) , .A1( us32_n857 ) );
  INV_X1 us32_U123 (.A( us32_n709 ) , .ZN( us32_n857 ) );
  AOI221_X1 us32_U124 (.A( us32_n710 ) , .ZN( us32_n721 ) , .C2( us32_n844 ) , .B2( us32_n845 ) , .C1( us32_n861 ) , .B1( us32_n862 ) );
  NOR4_X1 us32_U125 (.A4( us32_n715 ) , .A3( us32_n716 ) , .A2( us32_n717 ) , .A1( us32_n718 ) , .ZN( us32_n719 ) );
  NOR2_X1 us32_U126 (.ZN( us32_n733 ) , .A2( us32_n832 ) , .A1( us32_n845 ) );
  NOR2_X1 us32_U127 (.ZN( us32_n789 ) , .A2( us32_n862 ) , .A1( us32_n868 ) );
  NAND4_X1 us32_U128 (.A4( us32_n573 ) , .A3( us32_n574 ) , .A1( us32_n575 ) , .ZN( us32_n723 ) , .A2( us32_n874 ) );
  AOI221_X1 us32_U129 (.A( us32_n564 ) , .C2( us32_n565 ) , .ZN( us32_n574 ) , .B2( us32_n845 ) , .B1( us32_n852 ) , .C1( us32_n853 ) );
  INV_X1 us32_U13 (.A( us32_n607 ) , .ZN( us32_n874 ) );
  NOR4_X1 us32_U130 (.A4( us32_n569 ) , .A3( us32_n570 ) , .A2( us32_n571 ) , .A1( us32_n572 ) , .ZN( us32_n573 ) );
  NOR2_X1 us32_U131 (.ZN( us32_n575 ) , .A1( us32_n622 ) , .A2( us32_n745 ) );
  NOR2_X1 us32_U132 (.ZN( us32_n748 ) , .A1( us32_n861 ) , .A2( us32_n862 ) );
  NAND4_X1 us32_U133 (.A4( us32_n633 ) , .A3( us32_n634 ) , .A2( us32_n635 ) , .A1( us32_n636 ) , .ZN( us32_n743 ) );
  AOI211_X1 us32_U134 (.B( us32_n623 ) , .A( us32_n624 ) , .ZN( us32_n635 ) , .C2( us32_n836 ) , .C1( us32_n863 ) );
  NOR4_X1 us32_U135 (.A4( us32_n629 ) , .A3( us32_n630 ) , .A2( us32_n631 ) , .A1( us32_n632 ) , .ZN( us32_n633 ) );
  NOR4_X1 us32_U136 (.A4( us32_n626 ) , .A3( us32_n627 ) , .A2( us32_n628 ) , .ZN( us32_n634 ) , .A1( us32_n664 ) );
  NAND4_X1 us32_U137 (.A4( us32_n493 ) , .A3( us32_n494 ) , .A1( us32_n495 ) , .ZN( us32_n802 ) , .A2( us32_n867 ) );
  AOI221_X1 us32_U138 (.A( us32_n489 ) , .ZN( us32_n494 ) , .B2( us32_n836 ) , .C2( us32_n841 ) , .C1( us32_n851 ) , .B1( us32_n860 ) );
  INV_X1 us32_U139 (.A( us32_n778 ) , .ZN( us32_n867 ) );
  INV_X1 us32_U14 (.A( us32_n680 ) , .ZN( us32_n840 ) );
  NOR4_X1 us32_U140 (.A2( us32_n491 ) , .A1( us32_n492 ) , .ZN( us32_n493 ) , .A3( us32_n580 ) , .A4( us32_n612 ) );
  NOR4_X1 us32_U141 (.A4( us32_n734 ) , .A3( us32_n735 ) , .A2( us32_n736 ) , .A1( us32_n737 ) , .ZN( us32_n738 ) );
  AOI211_X1 us32_U142 (.B( us32_n725 ) , .A( us32_n726 ) , .ZN( us32_n739 ) , .C1( us32_n843 ) , .C2( us32_n855 ) );
  NOR3_X1 us32_U143 (.A3( us32_n722 ) , .A1( us32_n723 ) , .ZN( us32_n740 ) , .A2( us32_n741 ) );
  NOR2_X1 us32_U144 (.ZN( us32_n647 ) , .A1( us32_n854 ) , .A2( us32_n868 ) );
  INV_X1 us32_U145 (.A( us32_n762 ) , .ZN( us32_n830 ) );
  INV_X1 us32_U146 (.A( us32_n754 ) , .ZN( us32_n869 ) );
  OAI21_X1 us32_U147 (.B1( us32_n753 ) , .ZN( us32_n754 ) , .A( us32_n845 ) , .B2( us32_n868 ) );
  INV_X1 us32_U148 (.A( us32_n697 ) , .ZN( us32_n838 ) );
  OR4_X1 us32_U149 (.ZN( us32_n492 ) , .A4( us32_n534 ) , .A2( us32_n547 ) , .A1( us32_n559 ) , .A3( us32_n632 ) );
  NOR4_X1 us32_U15 (.A4( us32_n445 ) , .A3( us32_n446 ) , .A2( us32_n516 ) , .A1( us32_n541 ) , .ZN( us32_n706 ) );
  OR4_X1 us32_U150 (.A4( us32_n566 ) , .A3( us32_n567 ) , .A2( us32_n568 ) , .ZN( us32_n572 ) , .A1( us32_n665 ) );
  OR4_X1 us32_U151 (.A4( us32_n682 ) , .A3( us32_n683 ) , .A2( us32_n684 ) , .A1( us32_n685 ) , .ZN( us32_n690 ) );
  OR4_X1 us32_U152 (.ZN( us32_n466 ) , .A4( us32_n518 ) , .A3( us32_n529 ) , .A2( us32_n578 ) , .A1( us32_n712 ) );
  OR4_X1 us32_U153 (.A4( us32_n518 ) , .A2( us32_n519 ) , .A1( us32_n520 ) , .ZN( us32_n522 ) , .A3( us32_n821 ) );
  OR4_X1 us32_U154 (.A4( us32_n580 ) , .A3( us32_n581 ) , .A2( us32_n582 ) , .A1( us32_n583 ) , .ZN( us32_n584 ) );
  NAND2_X1 us32_U155 (.ZN( us32_n613 ) , .A2( us32_n837 ) , .A1( us32_n873 ) );
  OR3_X1 us32_U156 (.A3( us32_n506 ) , .A2( us32_n507 ) , .A1( us32_n508 ) , .ZN( us32_n511 ) );
  INV_X1 us32_U157 (.A( us32_n672 ) , .ZN( us32_n859 ) );
  AOI21_X1 us32_U158 (.A( us32_n670 ) , .B1( us32_n671 ) , .ZN( us32_n672 ) , .B2( us32_n856 ) );
  INV_X1 us32_U159 (.A( us32_n463 ) , .ZN( us32_n864 ) );
  OR3_X1 us32_U16 (.ZN( us32_n446 ) , .A1( us32_n528 ) , .A3( us32_n577 ) , .A2( us32_n875 ) );
  OAI21_X1 us32_U160 (.ZN( us32_n463 ) , .B1( us32_n809 ) , .A( us32_n834 ) , .B2( us32_n851 ) );
  OAI222_X1 us32_U161 (.B2( us32_n708 ) , .ZN( us32_n709 ) , .C2( us32_n724 ) , .B1( us32_n747 ) , .A1( us32_n806 ) , .C1( us32_n814 ) , .A2( us32_n815 ) );
  NAND2_X1 us32_U162 (.A1( us32_n447 ) , .A2( us32_n465 ) , .ZN( us32_n749 ) );
  AOI22_X1 us32_U163 (.A2( us32_n782 ) , .ZN( us32_n783 ) , .B2( us32_n831 ) , .A1( us32_n834 ) , .B1( us32_n863 ) );
  AOI22_X1 us32_U164 (.ZN( us32_n696 ) , .A1( us32_n830 ) , .B2( us32_n843 ) , .A2( us32_n865 ) , .B1( us32_n868 ) );
  INV_X1 us32_U165 (.A( us32_n730 ) , .ZN( us32_n839 ) );
  AOI221_X1 us32_U166 (.A( us32_n483 ) , .ZN( us32_n488 ) , .B1( us32_n831 ) , .C2( us32_n844 ) , .C1( us32_n852 ) , .B2( us32_n862 ) );
  OAI22_X1 us32_U167 (.ZN( us32_n483 ) , .A1( us32_n708 ) , .B2( us32_n785 ) , .A2( us32_n806 ) , .B1( us32_n812 ) );
  INV_X1 us32_U168 (.A( us32_n790 ) , .ZN( us32_n832 ) );
  OAI221_X1 us32_U169 (.A( us32_n727 ) , .C2( us32_n728 ) , .B2( us32_n729 ) , .B1( us32_n730 ) , .ZN( us32_n737 ) , .C1( us32_n817 ) );
  OR4_X1 us32_U17 (.A4( us32_n442 ) , .A2( us32_n443 ) , .A1( us32_n444 ) , .ZN( us32_n445 ) , .A3( us32_n553 ) );
  AOI22_X1 us32_U170 (.ZN( us32_n727 ) , .B1( us32_n832 ) , .A2( us32_n838 ) , .A1( us32_n863 ) , .B2( us32_n866 ) );
  NAND2_X1 us32_U171 (.A1( us32_n451 ) , .A2( us32_n453 ) , .ZN( us32_n762 ) );
  INV_X1 us32_U172 (.A( us32_n786 ) , .ZN( us32_n862 ) );
  OAI22_X1 us32_U173 (.ZN( us32_n710 ) , .A2( us32_n728 ) , .B2( us32_n729 ) , .A1( us32_n744 ) , .B1( us32_n813 ) );
  INV_X1 us32_U174 (.A( us32_n816 ) , .ZN( us32_n831 ) );
  OAI22_X1 us32_U175 (.ZN( us32_n489 ) , .A1( us32_n724 ) , .B2( us32_n728 ) , .B1( us32_n730 ) , .A2( us32_n779 ) );
  OAI22_X1 us32_U176 (.ZN( us32_n624 ) , .B1( us32_n669 ) , .B2( us32_n747 ) , .A1( us32_n815 ) , .A2( us32_n816 ) );
  INV_X1 us32_U177 (.A( us32_n788 ) , .ZN( us32_n845 ) );
  OAI22_X1 us32_U178 (.A1( us32_n724 ) , .ZN( us32_n726 ) , .B2( us32_n750 ) , .B1( us32_n812 ) , .A2( us32_n816 ) );
  INV_X1 us32_U179 (.A( us32_n744 ) , .ZN( us32_n837 ) );
  INV_X1 us32_U18 (.A( us32_n613 ) , .ZN( us32_n875 ) );
  OAI22_X1 us32_U180 (.B2( us32_n779 ) , .B1( us32_n780 ) , .ZN( us32_n781 ) , .A2( us32_n814 ) , .A1( us32_n815 ) );
  INV_X1 us32_U181 (.A( us32_n814 ) , .ZN( us32_n833 ) );
  INV_X1 us32_U182 (.A( us32_n669 ) , .ZN( us32_n865 ) );
  OAI22_X1 us32_U183 (.B2( us32_n744 ) , .ZN( us32_n746 ) , .A2( us32_n762 ) , .B1( us32_n780 ) , .A1( us32_n792 ) );
  OAI22_X1 us32_U184 (.ZN( us32_n496 ) , .A2( us32_n744 ) , .A1( us32_n780 ) , .B1( us32_n791 ) , .B2( us32_n806 ) );
  AOI211_X1 us32_U185 (.A( us32_n637 ) , .ZN( us32_n645 ) , .B( us32_n743 ) , .C2( us32_n839 ) , .C1( us32_n854 ) );
  OAI22_X1 us32_U186 (.ZN( us32_n637 ) , .A1( us32_n699 ) , .B2( us32_n728 ) , .A2( us32_n762 ) , .B1( us32_n816 ) );
  INV_X1 us32_U187 (.A( us32_n750 ) , .ZN( us32_n842 ) );
  OAI22_X1 us32_U188 (.B1( us32_n490 ) , .ZN( us32_n491 ) , .A1( us32_n686 ) , .A2( us32_n763 ) , .B2( us32_n817 ) );
  NOR3_X1 us32_U189 (.ZN( us32_n490 ) , .A1( us32_n782 ) , .A2( us32_n850 ) , .A3( us32_n863 ) );
  INV_X1 us32_U19 (.A( us32_n749 ) , .ZN( us32_n863 ) );
  OAI22_X1 us32_U190 (.ZN( us32_n695 ) , .A2( us32_n730 ) , .A1( us32_n780 ) , .B1( us32_n791 ) , .B2( us32_n817 ) );
  NOR2_X1 us32_U191 (.ZN( us32_n666 ) , .A1( us32_n728 ) , .A2( us32_n803 ) );
  NOR2_X1 us32_U192 (.ZN( us32_n594 ) , .A2( us32_n697 ) , .A1( us32_n728 ) );
  NOR2_X1 us32_U193 (.ZN( us32_n570 ) , .A1( us32_n728 ) , .A2( us32_n806 ) );
  NOR2_X1 us32_U194 (.ZN( us32_n654 ) , .A1( us32_n728 ) , .A2( us32_n813 ) );
  NOR2_X1 us32_U195 (.ZN( us32_n546 ) , .A2( us32_n780 ) , .A1( us32_n814 ) );
  NOR2_X1 us32_U196 (.ZN( us32_n532 ) , .A2( us32_n749 ) , .A1( us32_n750 ) );
  NOR2_X1 us32_U197 (.ZN( us32_n577 ) , .A2( us32_n699 ) , .A1( us32_n814 ) );
  NOR2_X1 us32_U198 (.ZN( us32_n615 ) , .A1( us32_n785 ) , .A2( us32_n815 ) );
  NOR2_X1 us32_U199 (.ZN( us32_n629 ) , .A2( us32_n728 ) , .A1( us32_n785 ) );
  AOI222_X1 us32_U20 (.ZN( us32_n605 ) , .B2( us32_n671 ) , .B1( us32_n753 ) , .C2( us32_n831 ) , .A1( us32_n833 ) , .A2( us32_n862 ) , .C1( us32_n863 ) );
  NOR2_X1 us32_U200 (.ZN( us32_n718 ) , .A2( us32_n724 ) , .A1( us32_n744 ) );
  NOR2_X1 us32_U201 (.ZN( us32_n628 ) , .A2( us32_n669 ) , .A1( us32_n785 ) );
  INV_X1 us32_U202 (.A( us32_n728 ) , .ZN( us32_n852 ) );
  NOR2_X1 us32_U203 (.A2( us32_n744 ) , .ZN( us32_n769 ) , .A1( us32_n812 ) );
  NOR2_X1 us32_U204 (.ZN( us32_n531 ) , .A2( us32_n780 ) , .A1( us32_n816 ) );
  NOR2_X1 us32_U205 (.A2( us32_n708 ) , .A1( us32_n750 ) , .ZN( us32_n771 ) );
  NOR2_X1 us32_U206 (.ZN( us32_n599 ) , .A2( us32_n791 ) , .A1( us32_n816 ) );
  NOR2_X1 us32_U207 (.ZN( us32_n611 ) , .A2( us32_n780 ) , .A1( us32_n806 ) );
  NOR2_X1 us32_U208 (.ZN( us32_n652 ) , .A1( us32_n669 ) , .A2( us32_n814 ) );
  INV_X1 us32_U209 (.A( us32_n792 ) , .ZN( us32_n851 ) );
  AOI222_X1 us32_U21 (.ZN( us32_n563 ) , .B1( us32_n830 ) , .C1( us32_n841 ) , .A2( us32_n843 ) , .A1( us32_n854 ) , .B2( us32_n863 ) , .C2( us32_n873 ) );
  NOR2_X1 us32_U210 (.A1( us32_n699 ) , .ZN( us32_n768 ) , .A2( us32_n813 ) );
  NOR2_X1 us32_U211 (.A1( us32_n669 ) , .ZN( us32_n673 ) , .A2( us32_n744 ) );
  NOR2_X1 us32_U212 (.ZN( us32_n541 ) , .A2( us32_n697 ) , .A1( us32_n699 ) );
  NOR2_X1 us32_U213 (.ZN( us32_n602 ) , .A1( us32_n669 ) , .A2( us32_n803 ) );
  NOR2_X1 us32_U214 (.A1( us32_n669 ) , .ZN( us32_n688 ) , .A2( us32_n816 ) );
  NOR2_X1 us32_U215 (.ZN( us32_n667 ) , .A1( us32_n750 ) , .A2( us32_n815 ) );
  NOR2_X1 us32_U216 (.ZN( us32_n555 ) , .A1( us32_n750 ) , .A2( us32_n791 ) );
  NOR2_X1 us32_U217 (.ZN( us32_n508 ) , .A2( us32_n780 ) , .A1( us32_n785 ) );
  NOR2_X1 us32_U218 (.ZN( us32_n543 ) , .A2( us32_n708 ) , .A1( us32_n785 ) );
  INV_X1 us32_U219 (.A( us32_n747 ) , .ZN( us32_n834 ) );
  AOI222_X1 us32_U22 (.ZN( us32_n660 ) , .A2( us32_n839 ) , .B1( us32_n841 ) , .C2( us32_n845 ) , .A1( us32_n860 ) , .C1( us32_n863 ) , .B2( us32_n870 ) );
  NOR2_X1 us32_U220 (.ZN( us32_n664 ) , .A1( us32_n785 ) , .A2( us32_n791 ) );
  NOR2_X1 us32_U221 (.A1( us32_n669 ) , .ZN( us32_n766 ) , .A2( us32_n813 ) );
  NOR2_X1 us32_U222 (.ZN( us32_n527 ) , .A1( us32_n669 ) , .A2( us32_n779 ) );
  NOR2_X1 us32_U223 (.ZN( us32_n661 ) , .A1( us32_n729 ) , .A2( us32_n790 ) );
  NOR2_X1 us32_U224 (.ZN( us32_n601 ) , .A2( us32_n780 ) , .A1( us32_n803 ) );
  NOR2_X1 us32_U225 (.ZN( us32_n507 ) , .A1( us32_n812 ) , .A2( us32_n817 ) );
  NOR2_X1 us32_U226 (.ZN( us32_n528 ) , .A2( us32_n724 ) , .A1( us32_n803 ) );
  NOR2_X1 us32_U227 (.ZN( us32_n509 ) , .A1( us32_n729 ) , .A2( us32_n779 ) );
  NOR2_X1 us32_U228 (.ZN( us32_n557 ) , .A1( us32_n792 ) , .A2( us32_n814 ) );
  NOR2_X1 us32_U229 (.ZN( us32_n545 ) , .A1( us32_n749 ) , .A2( us32_n814 ) );
  INV_X1 us32_U23 (.A( us32_n647 ) , .ZN( us32_n870 ) );
  OAI22_X1 us32_U230 (.B1( us32_n440 ) , .ZN( us32_n444 ) , .A2( us32_n728 ) , .A1( us32_n744 ) , .B2( us32_n749 ) );
  NOR3_X1 us32_U231 (.ZN( us32_n440 ) , .A2( us32_n836 ) , .A3( us32_n837 ) , .A1( us32_n846 ) );
  NOR2_X1 us32_U232 (.ZN( us32_n662 ) , .A2( us32_n697 ) , .A1( us32_n729 ) );
  OAI22_X1 us32_U233 (.B2( us32_n750 ) , .B1( us32_n751 ) , .A1( us32_n752 ) , .ZN( us32_n756 ) , .A2( us32_n806 ) );
  NOR2_X1 us32_U234 (.ZN( us32_n751 ) , .A2( us32_n852 ) , .A1( us32_n860 ) );
  NOR3_X1 us32_U235 (.ZN( us32_n752 ) , .A2( us32_n853 ) , .A1( us32_n863 ) , .A3( us32_n865 ) );
  NOR2_X1 us32_U236 (.ZN( us32_n544 ) , .A2( us32_n785 ) , .A1( us32_n792 ) );
  NOR2_X1 us32_U237 (.ZN( us32_n663 ) , .A1( us32_n729 ) , .A2( us32_n785 ) );
  INV_X1 us32_U238 (.A( us32_n806 ) , .ZN( us32_n841 ) );
  NOR2_X1 us32_U239 (.ZN( us32_n506 ) , .A2( us32_n728 ) , .A1( us32_n762 ) );
  NOR4_X1 us32_U24 (.A4( us32_n544 ) , .A3( us32_n545 ) , .A2( us32_n546 ) , .A1( us32_n547 ) , .ZN( us32_n548 ) );
  NOR2_X1 us32_U240 (.ZN( us32_n631 ) , .A1( us32_n724 ) , .A2( us32_n813 ) );
  NOR2_X1 us32_U241 (.ZN( us32_n614 ) , .A1( us32_n762 ) , .A2( us32_n812 ) );
  NOR2_X1 us32_U242 (.ZN( us32_n530 ) , .A2( us32_n744 ) , .A1( us32_n792 ) );
  NOR2_X1 us32_U243 (.ZN( us32_n558 ) , .A1( us32_n708 ) , .A2( us32_n816 ) );
  NOR2_X1 us32_U244 (.ZN( us32_n516 ) , .A1( us32_n708 ) , .A2( us32_n744 ) );
  NOR2_X1 us32_U245 (.A2( us32_n697 ) , .ZN( us32_n716 ) , .A1( us32_n792 ) );
  NOR2_X1 us32_U246 (.A1( us32_n749 ) , .ZN( us32_n767 ) , .A2( us32_n803 ) );
  NOR2_X1 us32_U247 (.ZN( us32_n521 ) , .A1( us32_n790 ) , .A2( us32_n812 ) );
  NOR2_X1 us32_U248 (.ZN( us32_n655 ) , .A1( us32_n790 ) , .A2( us32_n815 ) );
  NOR2_X1 us32_U249 (.ZN( us32_n668 ) , .A2( us32_n708 ) , .A1( us32_n790 ) );
  NOR4_X1 us32_U25 (.ZN( us32_n479 ) , .A1( us32_n520 ) , .A4( us32_n557 ) , .A3( us32_n582 ) , .A2( us32_n630 ) );
  NOR2_X1 us32_U250 (.ZN( us32_n517 ) , .A1( us32_n708 ) , .A2( us32_n803 ) );
  INV_X1 us32_U251 (.A( us32_n763 ) , .ZN( us32_n866 ) );
  NOR2_X1 us32_U252 (.ZN( us32_n542 ) , .A1( us32_n762 ) , .A2( us32_n791 ) );
  NOR2_X1 us32_U253 (.ZN( us32_n630 ) , .A1( us32_n747 ) , .A2( us32_n815 ) );
  INV_X1 us32_U254 (.A( us32_n729 ) , .ZN( us32_n868 ) );
  NOR2_X1 us32_U255 (.ZN( us32_n609 ) , .A2( us32_n724 ) , .A1( us32_n817 ) );
  AOI21_X1 us32_U256 (.A( us32_n815 ) , .B2( us32_n816 ) , .B1( us32_n817 ) , .ZN( us32_n818 ) );
  NOR2_X1 us32_U257 (.ZN( us32_n579 ) , .A2( us32_n708 ) , .A1( us32_n730 ) );
  NOR2_X1 us32_U258 (.ZN( us32_n533 ) , .A2( us32_n724 ) , .A1( us32_n730 ) );
  NOR2_X1 us32_U259 (.ZN( us32_n642 ) , .A2( us32_n788 ) , .A1( us32_n791 ) );
  NOR4_X1 us32_U26 (.ZN( us32_n456 ) , .A2( us32_n517 ) , .A1( us32_n543 ) , .A3( us32_n579 ) , .A4( us32_n615 ) );
  AOI21_X1 us32_U260 (.B1( us32_n625 ) , .ZN( us32_n627 ) , .A( us32_n763 ) , .B2( us32_n814 ) );
  NOR2_X1 us32_U261 (.ZN( us32_n656 ) , .A1( us32_n747 ) , .A2( us32_n780 ) );
  AOI21_X1 us32_U262 (.A( us32_n812 ) , .B2( us32_n813 ) , .B1( us32_n814 ) , .ZN( us32_n819 ) );
  NOR2_X1 us32_U263 (.A2( us32_n697 ) , .A1( us32_n780 ) , .ZN( us32_n820 ) );
  AOI21_X1 us32_U264 (.ZN( us32_n499 ) , .B1( us32_n680 ) , .A( us32_n812 ) , .B2( us32_n816 ) );
  NOR2_X1 us32_U265 (.A2( us32_n708 ) , .A1( us32_n762 ) , .ZN( us32_n794 ) );
  AOI21_X1 us32_U266 (.ZN( us32_n593 ) , .B1( us32_n750 ) , .A( us32_n792 ) , .B2( us32_n813 ) );
  AOI21_X1 us32_U267 (.ZN( us32_n626 ) , .B2( us32_n669 ) , .A( us32_n790 ) , .B1( us32_n791 ) );
  NOR2_X1 us32_U268 (.ZN( us32_n520 ) , .A2( us32_n708 ) , .A1( us32_n814 ) );
  NOR2_X1 us32_U269 (.A1( us32_n697 ) , .ZN( us32_n770 ) , .A2( us32_n815 ) );
  NOR4_X1 us32_U27 (.A4( us32_n532 ) , .A3( us32_n533 ) , .A2( us32_n534 ) , .ZN( us32_n535 ) , .A1( us32_n820 ) );
  NOR2_X1 us32_U270 (.ZN( us32_n582 ) , .A1( us32_n744 ) , .A2( us32_n815 ) );
  NOR2_X1 us32_U271 (.ZN( us32_n519 ) , .A2( us32_n699 ) , .A1( us32_n816 ) );
  AOI21_X1 us32_U272 (.ZN( us32_n477 ) , .A( us32_n669 ) , .B1( us32_n750 ) , .B2( us32_n806 ) );
  AOI21_X1 us32_U273 (.ZN( us32_n510 ) , .B2( us32_n669 ) , .A( us32_n730 ) , .B1( us32_n815 ) );
  INV_X1 us32_U274 (.A( us32_n813 ) , .ZN( us32_n836 ) );
  AOI21_X1 us32_U275 (.ZN( us32_n589 ) , .B2( us32_n699 ) , .B1( us32_n815 ) , .A( us32_n817 ) );
  AOI21_X1 us32_U276 (.ZN( us32_n515 ) , .A( us32_n729 ) , .B1( us32_n750 ) , .B2( us32_n803 ) );
  AOI21_X1 us32_U277 (.ZN( us32_n539 ) , .B2( us32_n812 ) , .A( us32_n814 ) , .B1( us32_n815 ) );
  NOR2_X1 us32_U278 (.ZN( us32_n581 ) , .A1( us32_n669 ) , .A2( us32_n788 ) );
  NOR2_X1 us32_U279 (.ZN( us32_n547 ) , .A1( us32_n699 ) , .A2( us32_n744 ) );
  NOR4_X1 us32_U28 (.ZN( us32_n474 ) , .A1( us32_n506 ) , .A3( us32_n544 ) , .A2( us32_n583 ) , .A4( us32_n716 ) );
  AOI21_X1 us32_U280 (.ZN( us32_n540 ) , .A( us32_n763 ) , .B2( us32_n779 ) , .B1( us32_n817 ) );
  AOI21_X1 us32_U281 (.B1( us32_n699 ) , .ZN( us32_n700 ) , .A( us32_n732 ) , .B2( us32_n763 ) );
  AOI21_X1 us32_U282 (.ZN( us32_n591 ) , .B2( us32_n763 ) , .A( us32_n785 ) , .B1( us32_n812 ) );
  INV_X1 us32_U283 (.A( us32_n791 ) , .ZN( us32_n873 ) );
  NOR2_X1 us32_U284 (.ZN( us32_n559 ) , .A2( us32_n791 ) , .A1( us32_n803 ) );
  AOI21_X1 us32_U285 (.ZN( us32_n498 ) , .A( us32_n724 ) , .B2( us32_n762 ) , .B1( us32_n814 ) );
  NOR2_X1 us32_U286 (.ZN( us32_n683 ) , .A2( us32_n699 ) , .A1( us32_n803 ) );
  NOR2_X1 us32_U287 (.ZN( us32_n685 ) , .A1( us32_n729 ) , .A2( us32_n816 ) );
  AOI21_X1 us32_U288 (.B1( us32_n686 ) , .ZN( us32_n687 ) , .A( us32_n728 ) , .B2( us32_n761 ) );
  AOI21_X1 us32_U289 (.ZN( us32_n569 ) , .B1( us32_n750 ) , .B2( us32_n762 ) , .A( us32_n780 ) );
  AOI221_X1 us32_U29 (.A( us32_n713 ) , .B2( us32_n714 ) , .ZN( us32_n720 ) , .C1( us32_n832 ) , .B1( us32_n839 ) , .C2( us32_n863 ) );
  AOI21_X1 us32_U290 (.ZN( us32_n649 ) , .B1( us32_n729 ) , .B2( us32_n763 ) , .A( us32_n813 ) );
  NOR2_X1 us32_U291 (.ZN( us32_n568 ) , .A1( us32_n729 ) , .A2( us32_n762 ) );
  INV_X1 us32_U292 (.A( us32_n699 ) , .ZN( us32_n853 ) );
  NOR2_X1 us32_U293 (.ZN( us32_n566 ) , .A2( us32_n697 ) , .A1( us32_n763 ) );
  AOI21_X1 us32_U294 (.ZN( us32_n514 ) , .A( us32_n779 ) , .B2( us32_n792 ) , .B1( us32_n812 ) );
  AOI21_X1 us32_U295 (.ZN( us32_n639 ) , .B2( us32_n749 ) , .A( us32_n788 ) , .B1( us32_n812 ) );
  NOR2_X1 us32_U296 (.ZN( us32_n665 ) , .A1( us32_n780 ) , .A2( us32_n813 ) );
  AOI21_X1 us32_U297 (.ZN( us32_n571 ) , .B2( us32_n697 ) , .B1( us32_n806 ) , .A( us32_n812 ) );
  AOI21_X1 us32_U298 (.ZN( us32_n564 ) , .B1( us32_n724 ) , .A( us32_n779 ) , .B2( us32_n791 ) );
  AOI21_X1 us32_U299 (.ZN( us32_n497 ) , .A( us32_n779 ) , .B2( us32_n791 ) , .B1( us32_n804 ) );
  NAND2_X1 us32_U3 (.A1( us32_n449 ) , .A2( us32_n464 ) , .ZN( us32_n724 ) );
  OR2_X1 us32_U30 (.A2( us32_n711 ) , .A1( us32_n712 ) , .ZN( us32_n713 ) );
  AOI21_X1 us32_U300 (.ZN( us32_n640 ) , .B2( us32_n747 ) , .A( us32_n792 ) , .B1( us32_n803 ) );
  NOR2_X1 us32_U301 (.ZN( us32_n578 ) , .A1( us32_n708 ) , .A2( us32_n813 ) );
  NOR2_X1 us32_U302 (.ZN( us32_n529 ) , .A1( us32_n708 ) , .A2( us32_n779 ) );
  AOI21_X1 us32_U303 (.ZN( us32_n689 ) , .B2( us32_n749 ) , .B1( us32_n763 ) , .A( us32_n806 ) );
  AOI21_X1 us32_U304 (.A( us32_n790 ) , .B2( us32_n791 ) , .B1( us32_n792 ) , .ZN( us32_n793 ) );
  AOI21_X1 us32_U305 (.ZN( us32_n478 ) , .B2( us32_n697 ) , .A( us32_n749 ) , .B1( us32_n779 ) );
  NOR2_X1 us32_U306 (.ZN( us32_n684 ) , .A1( us32_n791 ) , .A2( us32_n813 ) );
  AOI21_X1 us32_U307 (.ZN( us32_n450 ) , .B2( us32_n792 ) , .A( us32_n803 ) , .B1( us32_n815 ) );
  AOI21_X1 us32_U308 (.A( us32_n733 ) , .ZN( us32_n734 ) , .B2( us32_n780 ) , .B1( us32_n792 ) );
  NOR2_X1 us32_U309 (.A2( us32_n813 ) , .A1( us32_n815 ) , .ZN( us32_n821 ) );
  NOR2_X1 us32_U31 (.ZN( us32_n680 ) , .A2( us32_n834 ) , .A1( us32_n839 ) );
  AOI21_X1 us32_U310 (.ZN( us32_n641 ) , .B1( us32_n680 ) , .A( us32_n791 ) , .B2( us32_n817 ) );
  NOR2_X1 us32_U311 (.ZN( us32_n583 ) , .A1( us32_n792 ) , .A2( us32_n817 ) );
  NOR2_X1 us32_U312 (.ZN( us32_n711 ) , .A1( us32_n762 ) , .A2( us32_n763 ) );
  NOR2_X1 us32_U313 (.ZN( us32_n534 ) , .A1( us32_n724 ) , .A2( us32_n788 ) );
  NOR2_X1 us32_U314 (.ZN( us32_n632 ) , .A2( us32_n697 ) , .A1( us32_n724 ) );
  NOR2_X1 us32_U315 (.ZN( us32_n580 ) , .A2( us32_n697 ) , .A1( us32_n791 ) );
  NOR2_X1 us32_U316 (.ZN( us32_n682 ) , .A2( us32_n708 ) , .A1( us32_n817 ) );
  INV_X1 us32_U317 (.A( us32_n815 ) , .ZN( us32_n855 ) );
  AOI21_X1 us32_U318 (.ZN( us32_n442 ) , .A( us32_n699 ) , .B1( us32_n733 ) , .B2( us32_n750 ) );
  INV_X1 us32_U319 (.A( us32_n780 ) , .ZN( us32_n850 ) );
  NOR4_X1 us32_U32 (.A4( us32_n514 ) , .A3( us32_n515 ) , .A2( us32_n516 ) , .A1( us32_n517 ) , .ZN( us32_n524 ) );
  INV_X1 us32_U320 (.A( us32_n785 ) , .ZN( us32_n846 ) );
  NAND2_X1 us32_U321 (.ZN( us32_n714 ) , .A1( us32_n728 ) , .A2( us32_n780 ) );
  NAND2_X1 us32_U322 (.ZN( us32_n671 ) , .A1( us32_n806 ) , .A2( us32_n816 ) );
  AOI21_X1 us32_U323 (.ZN( us32_n443 ) , .B1( us32_n789 ) , .B2( us32_n791 ) , .A( us32_n814 ) );
  NOR2_X1 us32_U324 (.ZN( us32_n470 ) , .A2( us32_n779 ) , .A1( us32_n815 ) );
  NAND2_X1 us32_U325 (.A2( us32_n762 ) , .A1( us32_n806 ) , .ZN( us32_n810 ) );
  NOR2_X1 us32_U326 (.ZN( us32_n526 ) , .A1( us32_n724 ) , .A2( us32_n750 ) );
  OAI21_X1 us32_U327 (.A( us32_n787 ) , .B2( us32_n788 ) , .B1( us32_n789 ) , .ZN( us32_n795 ) );
  OAI21_X1 us32_U328 (.ZN( us32_n787 ) , .A( us32_n839 ) , .B1( us32_n863 ) , .B2( us32_n873 ) );
  NAND2_X1 us32_U329 (.A1( us32_n699 ) , .A2( us32_n729 ) , .ZN( us32_n782 ) );
  AOI222_X1 us32_U33 (.ZN( us32_n525 ) , .A1( us32_n834 ) , .B2( us32_n837 ) , .C1( us32_n844 ) , .C2( us32_n850 ) , .A2( us32_n852 ) , .B1( us32_n866 ) );
  NOR2_X1 us32_U330 (.ZN( us32_n712 ) , .A2( us32_n724 ) , .A1( us32_n790 ) );
  NOR2_X1 us32_U331 (.ZN( us32_n518 ) , .A1( us32_n708 ) , .A2( us32_n788 ) );
  OAI21_X1 us32_U332 (.A( us32_n698 ) , .ZN( us32_n702 ) , .B2( us32_n750 ) , .B1( us32_n804 ) );
  OAI21_X1 us32_U333 (.ZN( us32_n698 ) , .B2( us32_n833 ) , .B1( us32_n838 ) , .A( us32_n860 ) );
  INV_X1 us32_U334 (.A( us32_n817 ) , .ZN( us32_n844 ) );
  INV_X1 us32_U335 (.A( us32_n724 ) , .ZN( us32_n856 ) );
  OAI21_X1 us32_U336 (.ZN( us32_n731 ) , .A( us32_n833 ) , .B2( us32_n852 ) , .B1( us32_n873 ) );
  AND2_X1 us32_U337 (.ZN( us32_n732 ) , .A1( us32_n779 ) , .A2( us32_n785 ) );
  AOI221_X1 us32_U338 (.A( us32_n764 ) , .ZN( us32_n774 ) , .C2( us32_n810 ) , .B2( us32_n835 ) , .C1( us32_n855 ) , .B1( us32_n866 ) );
  AOI21_X1 us32_U339 (.B2( us32_n763 ) , .ZN( us32_n764 ) , .A( us32_n788 ) , .B1( us32_n792 ) );
  NOR4_X1 us32_U34 (.A3( us32_n521 ) , .A1( us32_n522 ) , .ZN( us32_n523 ) , .A2( us32_n673 ) , .A4( us32_n769 ) );
  INV_X1 us32_U340 (.A( us32_n761 ) , .ZN( us32_n835 ) );
  NAND2_X1 us32_U341 (.A2( us32_n448 ) , .A1( us32_n460 ) , .ZN( us32_n728 ) );
  NAND2_X1 us32_U342 (.A1( us32_n451 ) , .A2( us32_n454 ) , .ZN( us32_n814 ) );
  NAND2_X1 us32_U343 (.A1( us32_n455 ) , .A2( us32_n462 ) , .ZN( us32_n750 ) );
  NAND2_X1 us32_U344 (.A1( us32_n451 ) , .A2( us32_n471 ) , .ZN( us32_n816 ) );
  NAND2_X1 us32_U345 (.A1( us32_n454 ) , .A2( us32_n461 ) , .ZN( us32_n813 ) );
  NAND2_X1 us32_U346 (.A1( us32_n452 ) , .A2( us32_n465 ) , .ZN( us32_n669 ) );
  NAND2_X1 us32_U347 (.A1( us32_n453 ) , .A2( us32_n472 ) , .ZN( us32_n785 ) );
  NAND2_X1 us32_U348 (.A1( us32_n453 ) , .A2( us32_n461 ) , .ZN( us32_n744 ) );
  NAND2_X1 us32_U349 (.A2( us32_n453 ) , .A1( us32_n455 ) , .ZN( us32_n806 ) );
  AOI221_X1 us32_U35 (.A( us32_n781 ) , .ZN( us32_n798 ) , .C2( us32_n837 ) , .B2( us32_n838 ) , .B1( us32_n865 ) , .C1( us32_n866 ) );
  NAND2_X1 us32_U350 (.A1( us32_n455 ) , .A2( us32_n471 ) , .ZN( us32_n803 ) );
  NAND2_X1 us32_U351 (.A2( us32_n454 ) , .A1( us32_n472 ) , .ZN( us32_n779 ) );
  NAND2_X1 us32_U352 (.A2( us32_n464 ) , .A1( us32_n465 ) , .ZN( us32_n812 ) );
  NAND2_X1 us32_U353 (.A1( us32_n441 ) , .A2( us32_n460 ) , .ZN( us32_n699 ) );
  NAND2_X1 us32_U354 (.A2( us32_n448 ) , .A1( us32_n452 ) , .ZN( us32_n729 ) );
  NAND2_X1 us32_U355 (.A2( us32_n449 ) , .A1( us32_n452 ) , .ZN( us32_n763 ) );
  NOR2_X1 us32_U356 (.ZN( us32_n465 ) , .A2( us32_n847 ) , .A1( us32_n848 ) );
  NOR2_X1 us32_U357 (.ZN( us32_n453 ) , .A1( us32_n826 ) , .A2( us32_n827 ) );
  NAND2_X1 us32_U358 (.A1( us32_n462 ) , .A2( us32_n472 ) , .ZN( us32_n788 ) );
  NOR2_X1 us32_U359 (.ZN( us32_n451 ) , .A1( us32_n828 ) , .A2( us32_n829 ) );
  NOR4_X1 us32_U36 (.A4( us32_n793 ) , .A3( us32_n794 ) , .A2( us32_n795 ) , .A1( us32_n796 ) , .ZN( us32_n797 ) );
  NAND2_X1 us32_U360 (.A2( us32_n461 ) , .A1( us32_n462 ) , .ZN( us32_n747 ) );
  NAND2_X1 us32_U361 (.A1( us32_n451 ) , .A2( us32_n462 ) , .ZN( us32_n790 ) );
  NAND2_X2 us32_U362 (.A2( us32_n448 ) , .A1( us32_n464 ) , .ZN( us32_n815 ) );
  NAND2_X1 us32_U363 (.A2( us32_n441 ) , .A1( us32_n447 ) , .ZN( us32_n784 ) );
  NAND2_X1 us32_U364 (.A1( us32_n447 ) , .A2( us32_n449 ) , .ZN( us32_n805 ) );
  NAND2_X1 us32_U365 (.A2( us32_n454 ) , .A1( us32_n455 ) , .ZN( us32_n730 ) );
  NAND2_X2 us32_U366 (.A1( us32_n449 ) , .A2( us32_n460 ) , .ZN( us32_n792 ) );
  NAND2_X2 us32_U367 (.A2( us32_n460 ) , .A1( us32_n465 ) , .ZN( us32_n780 ) );
  NOR2_X1 us32_U368 (.ZN( us32_n447 ) , .A2( us32_n849 ) , .A1( us32_n858 ) );
  NAND2_X1 us32_U369 (.A1( us32_n447 ) , .A2( us32_n448 ) , .ZN( us32_n786 ) );
  NOR4_X1 us32_U37 (.A4( us32_n776 ) , .A3( us32_n777 ) , .A1( us32_n778 ) , .ZN( us32_n799 ) , .A2( us32_n801 ) );
  NAND2_X1 us32_U370 (.A2( us32_n471 ) , .A1( us32_n472 ) , .ZN( us32_n817 ) );
  NOR2_X1 us32_U371 (.A2( sa32_6 ) , .A1( sa32_7 ) , .ZN( us32_n464 ) );
  NOR2_X1 us32_U372 (.A2( sa32_7 ) , .ZN( us32_n460 ) , .A1( us32_n849 ) );
  NOR2_X1 us32_U373 (.A2( sa32_4 ) , .ZN( us32_n449 ) , .A1( us32_n848 ) );
  NOR2_X1 us32_U374 (.A2( sa32_4 ) , .A1( sa32_5 ) , .ZN( us32_n441 ) );
  NOR2_X1 us32_U375 (.A2( sa32_5 ) , .ZN( us32_n448 ) , .A1( us32_n847 ) );
  NOR2_X1 us32_U376 (.A2( sa32_2 ) , .A1( sa32_3 ) , .ZN( us32_n472 ) );
  NOR2_X1 us32_U377 (.A2( sa32_6 ) , .ZN( us32_n452 ) , .A1( us32_n858 ) );
  NOR2_X1 us32_U378 (.A2( sa32_1 ) , .ZN( us32_n471 ) , .A1( us32_n826 ) );
  NOR2_X1 us32_U379 (.A2( sa32_0 ) , .ZN( us32_n454 ) , .A1( us32_n827 ) );
  NOR4_X1 us32_U38 (.A3( us32_n755 ) , .A2( us32_n756 ) , .A1( us32_n757 ) , .ZN( us32_n758 ) , .A4( us32_n869 ) );
  NOR2_X1 us32_U380 (.A2( sa32_0 ) , .A1( sa32_1 ) , .ZN( us32_n462 ) );
  NOR2_X1 us32_U381 (.A2( sa32_3 ) , .ZN( us32_n455 ) , .A1( us32_n828 ) );
  NOR2_X1 us32_U382 (.A2( sa32_2 ) , .ZN( us32_n461 ) , .A1( us32_n829 ) );
  INV_X1 us32_U383 (.A( sa32_4 ) , .ZN( us32_n847 ) );
  INV_X1 us32_U384 (.A( sa32_6 ) , .ZN( us32_n849 ) );
  INV_X1 us32_U385 (.A( sa32_3 ) , .ZN( us32_n829 ) );
  INV_X1 us32_U386 (.A( sa32_1 ) , .ZN( us32_n827 ) );
  INV_X1 us32_U387 (.A( sa32_0 ) , .ZN( us32_n826 ) );
  INV_X1 us32_U388 (.A( sa32_2 ) , .ZN( us32_n828 ) );
  INV_X1 us32_U389 (.A( sa32_5 ) , .ZN( us32_n848 ) );
  AOI211_X1 us32_U39 (.B( us32_n745 ) , .A( us32_n746 ) , .ZN( us32_n759 ) , .C1( us32_n832 ) , .C2( us32_n853 ) );
  INV_X1 us32_U390 (.A( sa32_7 ) , .ZN( us32_n858 ) );
  NAND2_X1 us32_U391 (.A2( us32_n461 ) , .A1( us32_n471 ) , .ZN( us32_n697 ) );
  OAI222_X1 us32_U392 (.B2( us32_n747 ) , .B1( us32_n748 ) , .A2( us32_n749 ) , .ZN( us32_n757 ) , .C2( us32_n805 ) , .C1( us32_n814 ) , .A1( us32_n817 ) );
  OAI22_X1 us32_U393 (.B2( us32_n803 ) , .B1( us32_n804 ) , .A2( us32_n805 ) , .A1( us32_n806 ) , .ZN( us32_n808 ) );
  OAI21_X1 us32_U394 (.A( us32_n731 ) , .B1( us32_n732 ) , .ZN( us32_n736 ) , .B2( us32_n805 ) );
  OAI222_X1 us32_U395 (.ZN( us32_n505 ) , .C2( us32_n625 ) , .B2( us32_n647 ) , .B1( us32_n747 ) , .A2( us32_n748 ) , .C1( us32_n805 ) , .A1( us32_n806 ) );
  AOI21_X1 us32_U396 (.ZN( us32_n650 ) , .A( us32_n779 ) , .B1( us32_n792 ) , .B2( us32_n805 ) );
  INV_X1 us32_U397 (.A( us32_n805 ) , .ZN( us32_n860 ) );
  NOR2_X1 us32_U398 (.ZN( us32_n735 ) , .A2( us32_n803 ) , .A1( us32_n805 ) );
  NOR2_X1 us32_U399 (.ZN( us32_n484 ) , .A1( us32_n788 ) , .A2( us32_n805 ) );
  NAND2_X1 us32_U4 (.A1( us32_n441 ) , .A2( us32_n464 ) , .ZN( us32_n708 ) );
  NOR3_X1 us32_U40 (.A3( us32_n741 ) , .A2( us32_n742 ) , .A1( us32_n743 ) , .ZN( us32_n760 ) );
  NOR2_X1 us32_U400 (.A2( us32_n744 ) , .ZN( us32_n755 ) , .A1( us32_n805 ) );
  NAND2_X1 us32_U401 (.ZN( us32_n753 ) , .A1( us32_n763 ) , .A2( us32_n805 ) );
  NOR2_X1 us32_U402 (.ZN( us32_n715 ) , .A1( us32_n805 ) , .A2( us32_n817 ) );
  NOR2_X1 us32_U403 (.ZN( us32_n567 ) , .A1( us32_n747 ) , .A2( us32_n805 ) );
  AOI21_X1 us32_U404 (.ZN( us32_n552 ) , .B1( us32_n669 ) , .A( us32_n697 ) , .B2( us32_n805 ) );
  NOR2_X1 us32_U405 (.ZN( us32_n556 ) , .A1( us32_n762 ) , .A2( us32_n805 ) );
  NOR2_X1 us32_U406 (.ZN( us32_n670 ) , .A1( us32_n790 ) , .A2( us32_n805 ) );
  OAI221_X1 us32_U407 (.A( us32_n783 ) , .C2( us32_n784 ) , .B2( us32_n785 ) , .B1( us32_n786 ) , .ZN( us32_n796 ) , .C1( us32_n813 ) );
  NAND2_X1 us32_U408 (.A1( us32_n729 ) , .A2( us32_n784 ) , .ZN( us32_n811 ) );
  OAI22_X1 us32_U409 (.ZN( us32_n588 ) , .A2( us32_n747 ) , .B2( us32_n762 ) , .A1( us32_n763 ) , .B1( us32_n784 ) );
  NAND4_X1 us32_U41 (.ZN( sa33_sr_3 ) , .A4( us32_n704 ) , .A3( us32_n705 ) , .A2( us32_n706 ) , .A1( us32_n707 ) );
  AOI21_X1 us32_U410 (.ZN( us32_n592 ) , .B1( us32_n728 ) , .B2( us32_n784 ) , .A( us32_n790 ) );
  AOI21_X1 us32_U411 (.ZN( us32_n623 ) , .B1( us32_n699 ) , .A( us32_n779 ) , .B2( us32_n784 ) );
  AOI21_X1 us32_U412 (.ZN( us32_n648 ) , .A( us32_n762 ) , .B2( us32_n784 ) , .B1( us32_n792 ) );
  OAI22_X1 us32_U413 (.ZN( us32_n681 ) , .A1( us32_n699 ) , .A2( us32_n730 ) , .B2( us32_n784 ) , .B1( us32_n817 ) );
  OAI21_X1 us32_U414 (.A( us32_n613 ) , .ZN( us32_n616 ) , .B1( us32_n625 ) , .B2( us32_n784 ) );
  NOR2_X1 us32_U415 (.ZN( us32_n610 ) , .A1( us32_n784 ) , .A2( us32_n816 ) );
  OAI222_X1 us32_U416 (.A2( us32_n669 ) , .ZN( us32_n674 ) , .B1( us32_n747 ) , .B2( us32_n784 ) , .C2( us32_n788 ) , .C1( us32_n815 ) , .A1( us32_n817 ) );
  NOR2_X1 us32_U417 (.ZN( us32_n651 ) , .A1( us32_n784 ) , .A2( us32_n788 ) );
  NOR2_X1 us32_U418 (.ZN( us32_n600 ) , .A2( us32_n697 ) , .A1( us32_n784 ) );
  NOR2_X1 us32_U419 (.ZN( us32_n553 ) , .A2( us32_n744 ) , .A1( us32_n784 ) );
  NOR4_X1 us32_U42 (.A4( us32_n700 ) , .A3( us32_n701 ) , .A2( us32_n702 ) , .A1( us32_n703 ) , .ZN( us32_n704 ) );
  INV_X1 us32_U420 (.A( us32_n784 ) , .ZN( us32_n861 ) );
  AOI21_X1 us32_U421 (.ZN( us32_n500 ) , .A( us32_n697 ) , .B1( us32_n708 ) , .B2( us32_n786 ) );
  OAI221_X1 us32_U422 (.A( us32_n696 ) , .ZN( us32_n703 ) , .C2( us32_n784 ) , .C1( us32_n785 ) , .B1( us32_n786 ) , .B2( us32_n806 ) );
  OAI22_X1 us32_U423 (.ZN( us32_n590 ) , .B1( us32_n730 ) , .B2( us32_n749 ) , .A2( us32_n786 ) , .A1( us32_n803 ) );
  NOR2_X1 us32_U424 (.ZN( us32_n612 ) , .A1( us32_n779 ) , .A2( us32_n786 ) );
  NAND2_X1 us32_U425 (.A2( us32_n749 ) , .A1( us32_n786 ) , .ZN( us32_n809 ) );
  OAI222_X1 us32_U426 (.ZN( us32_n617 ) , .B1( us32_n697 ) , .C1( us32_n724 ) , .C2( us32_n747 ) , .B2( us32_n786 ) , .A2( us32_n792 ) , .A1( us32_n816 ) );
  NOR2_X1 us32_U427 (.ZN( us32_n717 ) , .A2( us32_n744 ) , .A1( us32_n786 ) );
  NOR2_X1 us32_U428 (.ZN( us32_n653 ) , .A1( us32_n762 ) , .A2( us32_n786 ) );
  NOR2_X1 us32_U429 (.ZN( us32_n554 ) , .A1( us32_n786 ) , .A2( us32_n813 ) );
  AOI211_X1 us32_U43 (.B( us32_n694 ) , .A( us32_n695 ) , .ZN( us32_n705 ) , .C2( us32_n831 ) , .C1( us32_n851 ) );
  NOR2_X1 us32_U430 (.ZN( us32_n701 ) , .A2( us32_n786 ) , .A1( us32_n817 ) );
  NOR2_X1 us32_U431 (.A1( us32_n730 ) , .ZN( us32_n765 ) , .A2( us32_n786 ) );
  AND2_X1 us32_U432 (.ZN( us32_n438 ) , .A2( us32_n831 ) , .A1( us32_n854 ) );
  AND2_X1 us32_U433 (.ZN( us32_n439 ) , .A2( us32_n843 ) , .A1( us32_n861 ) );
  NOR3_X1 us32_U434 (.A1( us32_n438 ) , .A2( us32_n439 ) , .A3( us32_n576 ) , .ZN( us32_n587 ) );
  NAND4_X1 us32_U435 (.ZN( sa33_sr_2 ) , .A4( us32_n643 ) , .A3( us32_n644 ) , .A2( us32_n645 ) , .A1( us32_n646 ) );
  INV_X1 us32_U436 (.A( us32_n812 ) , .ZN( us32_n854 ) );
  NAND3_X1 us32_U437 (.ZN( sa33_sr_6 ) , .A3( us32_n797 ) , .A2( us32_n798 ) , .A1( us32_n799 ) );
  NAND3_X1 us32_U438 (.ZN( sa33_sr_5 ) , .A3( us32_n758 ) , .A2( us32_n759 ) , .A1( us32_n760 ) );
  NAND3_X1 us32_U439 (.ZN( sa33_sr_4 ) , .A3( us32_n738 ) , .A2( us32_n739 ) , .A1( us32_n740 ) );
  NOR2_X1 us32_U44 (.ZN( us32_n707 ) , .A2( us32_n776 ) , .A1( us32_n800 ) );
  NAND3_X1 us32_U440 (.A3( us32_n675 ) , .A2( us32_n676 ) , .A1( us32_n677 ) , .ZN( us32_n807 ) );
  NAND3_X1 us32_U441 (.ZN( us32_n638 ) , .A3( us32_n708 ) , .A2( us32_n724 ) , .A1( us32_n792 ) );
  NAND3_X1 us32_U442 (.A3( us32_n618 ) , .A2( us32_n619 ) , .A1( us32_n620 ) , .ZN( us32_n725 ) );
  NAND3_X1 us32_U443 (.A3( us32_n585 ) , .A2( us32_n586 ) , .A1( us32_n587 ) , .ZN( us32_n621 ) );
  NAND3_X1 us32_U444 (.ZN( us32_n565 ) , .A3( us32_n680 ) , .A2( us32_n750 ) , .A1( us32_n785 ) );
  NAND3_X1 us32_U445 (.A3( us32_n523 ) , .A2( us32_n524 ) , .A1( us32_n525 ) , .ZN( us32_n742 ) );
  NAND3_X1 us32_U446 (.A3( us32_n512 ) , .A1( us32_n513 ) , .ZN( us32_n608 ) , .A2( us32_n871 ) );
  NAND3_X1 us32_U447 (.A3( us32_n467 ) , .A2( us32_n468 ) , .A1( us32_n469 ) , .ZN( us32_n777 ) );
  INV_X1 us32_U448 (.A( us32_n803 ) , .ZN( us32_n843 ) );
  AOI21_X1 us32_U449 (.ZN( us32_n576 ) , .B2( us32_n724 ) , .B1( us32_n748 ) , .A( us32_n785 ) );
  AOI222_X1 us32_U45 (.B2( us32_n638 ) , .ZN( us32_n644 ) , .B1( us32_n841 ) , .A1( us32_n842 ) , .C2( us32_n846 ) , .C1( us32_n863 ) , .A2( us32_n865 ) );
  NOR4_X1 us32_U46 (.A4( us32_n639 ) , .A3( us32_n640 ) , .A2( us32_n641 ) , .A1( us32_n642 ) , .ZN( us32_n643 ) );
  NOR3_X1 us32_U47 (.A2( us32_n607 ) , .A1( us32_n608 ) , .ZN( us32_n646 ) , .A3( us32_n722 ) );
  NAND4_X1 us32_U48 (.ZN( sa33_sr_7 ) , .A4( us32_n822 ) , .A3( us32_n823 ) , .A2( us32_n824 ) , .A1( us32_n825 ) );
  NOR4_X1 us32_U49 (.A4( us32_n818 ) , .A3( us32_n819 ) , .A2( us32_n820 ) , .A1( us32_n821 ) , .ZN( us32_n822 ) );
  NAND2_X1 us32_U5 (.A2( us32_n441 ) , .A1( us32_n452 ) , .ZN( us32_n791 ) );
  AOI222_X1 us32_U50 (.C2( us32_n809 ) , .B2( us32_n810 ) , .A2( us32_n811 ) , .ZN( us32_n823 ) , .C1( us32_n832 ) , .A1( us32_n839 ) , .B1( us32_n853 ) );
  AOI211_X1 us32_U51 (.B( us32_n807 ) , .A( us32_n808 ) , .ZN( us32_n824 ) , .C1( us32_n842 ) , .C2( us32_n850 ) );
  NAND4_X1 us32_U52 (.ZN( sa33_sr_0 ) , .A4( us32_n501 ) , .A3( us32_n502 ) , .A2( us32_n503 ) , .A1( us32_n504 ) );
  AOI221_X1 us32_U53 (.A( us32_n497 ) , .ZN( us32_n502 ) , .B2( us32_n843 ) , .C1( us32_n846 ) , .C2( us32_n860 ) , .B1( us32_n862 ) );
  NOR4_X1 us32_U54 (.A4( us32_n498 ) , .A3( us32_n499 ) , .A2( us32_n500 ) , .ZN( us32_n501 ) , .A1( us32_n527 ) );
  AOI211_X1 us32_U55 (.A( us32_n496 ) , .ZN( us32_n503 ) , .B( us32_n802 ) , .C2( us32_n839 ) , .C1( us32_n851 ) );
  NAND4_X1 us32_U56 (.ZN( sa33_sr_1 ) , .A4( us32_n595 ) , .A3( us32_n596 ) , .A2( us32_n597 ) , .A1( us32_n598 ) );
  NOR4_X1 us32_U57 (.A4( us32_n591 ) , .A3( us32_n592 ) , .A2( us32_n593 ) , .A1( us32_n594 ) , .ZN( us32_n595 ) );
  AOI211_X1 us32_U58 (.B( us32_n589 ) , .A( us32_n590 ) , .ZN( us32_n596 ) , .C2( us32_n811 ) , .C1( us32_n833 ) );
  AOI211_X1 us32_U59 (.A( us32_n588 ) , .ZN( us32_n597 ) , .B( us32_n621 ) , .C1( us32_n845 ) , .C2( us32_n855 ) );
  NOR3_X1 us32_U6 (.ZN( us32_n598 ) , .A1( us32_n608 ) , .A3( us32_n723 ) , .A2( us32_n742 ) );
  NOR2_X1 us32_U60 (.ZN( us32_n804 ) , .A1( us32_n854 ) , .A2( us32_n861 ) );
  AOI222_X1 us32_U61 (.ZN( us32_n469 ) , .B1( us32_n832 ) , .A1( us32_n839 ) , .C1( us32_n842 ) , .C2( us32_n851 ) , .A2( us32_n855 ) , .B2( us32_n865 ) );
  NOR4_X1 us32_U62 (.A1( us32_n466 ) , .ZN( us32_n467 ) , .A4( us32_n542 ) , .A2( us32_n554 ) , .A3( us32_n614 ) );
  AOI221_X1 us32_U63 (.ZN( us32_n468 ) , .C2( us32_n714 ) , .B2( us32_n831 ) , .C1( us32_n845 ) , .B1( us32_n860 ) , .A( us32_n864 ) );
  NAND4_X1 us32_U64 (.A4( us32_n603 ) , .A3( us32_n604 ) , .A2( us32_n605 ) , .A1( us32_n606 ) , .ZN( us32_n722 ) );
  NOR3_X1 us32_U65 (.A1( us32_n599 ) , .ZN( us32_n604 ) , .A3( us32_n663 ) , .A2( us32_n770 ) );
  NOR4_X1 us32_U66 (.A3( us32_n600 ) , .A2( us32_n601 ) , .A1( us32_n602 ) , .ZN( us32_n603 ) , .A4( us32_n655 ) );
  AOI222_X1 us32_U67 (.ZN( us32_n606 ) , .A1( us32_n830 ) , .C2( us32_n837 ) , .B1( us32_n842 ) , .A2( us32_n856 ) , .B2( us32_n861 ) , .C1( us32_n868 ) );
  NAND4_X1 us32_U68 (.A4( us32_n657 ) , .A3( us32_n658 ) , .A2( us32_n659 ) , .A1( us32_n660 ) , .ZN( us32_n800 ) );
  NOR3_X1 us32_U69 (.A3( us32_n648 ) , .A2( us32_n649 ) , .A1( us32_n650 ) , .ZN( us32_n659 ) );
  NOR3_X1 us32_U7 (.A3( us32_n800 ) , .A2( us32_n801 ) , .A1( us32_n802 ) , .ZN( us32_n825 ) );
  NOR3_X1 us32_U70 (.A3( us32_n651 ) , .A2( us32_n652 ) , .A1( us32_n653 ) , .ZN( us32_n658 ) );
  NOR3_X1 us32_U71 (.A3( us32_n654 ) , .A2( us32_n655 ) , .A1( us32_n656 ) , .ZN( us32_n657 ) );
  NAND4_X1 us32_U72 (.A4( us32_n560 ) , .A3( us32_n561 ) , .A2( us32_n562 ) , .A1( us32_n563 ) , .ZN( us32_n607 ) );
  NOR4_X1 us32_U73 (.A4( us32_n556 ) , .A3( us32_n557 ) , .A2( us32_n558 ) , .A1( us32_n559 ) , .ZN( us32_n560 ) );
  NOR4_X1 us32_U74 (.ZN( us32_n561 ) , .A1( us32_n653 ) , .A3( us32_n661 ) , .A4( us32_n685 ) , .A2( us32_n768 ) );
  NOR4_X1 us32_U75 (.A4( us32_n552 ) , .A3( us32_n553 ) , .A2( us32_n554 ) , .A1( us32_n555 ) , .ZN( us32_n562 ) );
  NAND4_X1 us32_U76 (.A4( us32_n772 ) , .A3( us32_n773 ) , .A2( us32_n774 ) , .A1( us32_n775 ) , .ZN( us32_n801 ) );
  NOR3_X1 us32_U77 (.A3( us32_n765 ) , .A2( us32_n766 ) , .A1( us32_n767 ) , .ZN( us32_n773 ) );
  NOR4_X1 us32_U78 (.A4( us32_n768 ) , .A3( us32_n769 ) , .A2( us32_n770 ) , .A1( us32_n771 ) , .ZN( us32_n772 ) );
  AOI222_X1 us32_U79 (.ZN( us32_n775 ) , .A1( us32_n830 ) , .C1( us32_n834 ) , .B2( us32_n841 ) , .A2( us32_n850 ) , .B1( us32_n861 ) , .C2( us32_n873 ) );
  NOR3_X1 us32_U8 (.A3( us32_n621 ) , .A2( us32_n622 ) , .ZN( us32_n636 ) , .A1( us32_n725 ) );
  NOR4_X1 us32_U80 (.A4( us32_n665 ) , .A3( us32_n666 ) , .A2( us32_n667 ) , .A1( us32_n668 ) , .ZN( us32_n676 ) );
  NOR4_X1 us32_U81 (.A4( us32_n661 ) , .A3( us32_n662 ) , .A2( us32_n663 ) , .A1( us32_n664 ) , .ZN( us32_n677 ) );
  NOR4_X1 us32_U82 (.A3( us32_n673 ) , .A1( us32_n674 ) , .ZN( us32_n675 ) , .A4( us32_n715 ) , .A2( us32_n859 ) );
  NOR2_X1 us32_U83 (.ZN( us32_n625 ) , .A2( us32_n836 ) , .A1( us32_n839 ) );
  NOR2_X1 us32_U84 (.ZN( us32_n761 ) , .A1( us32_n833 ) , .A2( us32_n834 ) );
  NOR4_X1 us32_U85 (.A4( us32_n577 ) , .A3( us32_n578 ) , .A2( us32_n579 ) , .ZN( us32_n586 ) , .A1( us32_n683 ) );
  NOR4_X1 us32_U86 (.A1( us32_n584 ) , .ZN( us32_n585 ) , .A3( us32_n652 ) , .A2( us32_n662 ) , .A4( us32_n767 ) );
  AOI222_X1 us32_U87 (.ZN( us32_n513 ) , .C1( us32_n832 ) , .B2( us32_n837 ) , .A2( us32_n843 ) , .C2( us32_n862 ) , .B1( us32_n863 ) , .A1( us32_n866 ) );
  NOR4_X1 us32_U88 (.A4( us32_n509 ) , .A2( us32_n510 ) , .A1( us32_n511 ) , .ZN( us32_n512 ) , .A3( us32_n670 ) );
  INV_X1 us32_U89 (.A( us32_n505 ) , .ZN( us32_n871 ) );
  NOR2_X1 us32_U9 (.ZN( us32_n495 ) , .A1( us32_n678 ) , .A2( us32_n694 ) );
  NAND4_X1 us32_U90 (.A4( us32_n456 ) , .A3( us32_n457 ) , .A2( us32_n458 ) , .A1( us32_n459 ) , .ZN( us32_n679 ) );
  NOR3_X1 us32_U91 (.ZN( us32_n457 ) , .A3( us32_n530 ) , .A1( us32_n555 ) , .A2( us32_n570 ) );
  AOI221_X1 us32_U92 (.A( us32_n450 ) , .ZN( us32_n459 ) , .C2( us32_n753 ) , .B1( us32_n832 ) , .C1( us32_n842 ) , .B2( us32_n861 ) );
  NOR4_X1 us32_U93 (.ZN( us32_n458 ) , .A2( us32_n509 ) , .A1( us32_n599 ) , .A4( us32_n628 ) , .A3( us32_n711 ) );
  NAND4_X1 us32_U94 (.A4( us32_n535 ) , .A3( us32_n536 ) , .A2( us32_n537 ) , .A1( us32_n538 ) , .ZN( us32_n622 ) );
  NOR4_X1 us32_U95 (.A4( us32_n526 ) , .A2( us32_n527 ) , .A1( us32_n528 ) , .ZN( us32_n538 ) , .A3( us32_n701 ) );
  NOR4_X1 us32_U96 (.A1( us32_n531 ) , .ZN( us32_n536 ) , .A2( us32_n654 ) , .A4( us32_n668 ) , .A3( us32_n765 ) );
  NOR4_X1 us32_U97 (.A4( us32_n529 ) , .A3( us32_n530 ) , .ZN( us32_n537 ) , .A2( us32_n684 ) , .A1( us32_n794 ) );
  NAND4_X1 us32_U98 (.A4( us32_n479 ) , .A3( us32_n480 ) , .A2( us32_n481 ) , .A1( us32_n482 ) , .ZN( us32_n694 ) );
  NOR3_X1 us32_U99 (.ZN( us32_n480 ) , .A2( us32_n508 ) , .A3( us32_n601 ) , .A1( us32_n610 ) );
endmodule

