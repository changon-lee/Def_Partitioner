module des_des_die_1 ( u0_K10_1, u0_K10_14, u0_K10_17, u0_K10_18, u0_K10_19, u0_K10_20, u0_K10_32, u0_K14_23, u0_K14_24, 
       u0_K14_25, u0_K14_26, u0_K14_29, u0_K14_5, u0_K14_7, u0_K4_36, u0_K4_43, u0_K4_48, u0_K4_6, 
       u0_K5_1, u0_K5_18, u0_K5_24, u0_K5_26, u0_K5_29, u0_K5_31, u0_K5_47, u0_K5_8, u0_K8_11, 
       u0_K8_13, u0_K8_19, u0_R11_16, u0_R11_20, u0_R12_16, u0_R12_17, u0_R12_19, u0_R12_20, u0_R12_22, 
       u0_R12_23, u0_R12_24, u0_R12_4, u0_R13_17, u0_R13_18, u0_R13_19, u0_R13_20, u0_R13_21, u0_R13_22, 
       u0_R13_23, u0_R13_24, u0_R13_25, u0_R13_26, u0_R13_27, u0_R13_28, u0_R13_29, u0_R13_30, u0_R13_31, 
       u0_R2_1, u0_R2_10, u0_R2_11, u0_R2_12, u0_R2_13, u0_R2_14, u0_R2_16, u0_R2_2, u0_R2_21, 
       u0_R2_22, u0_R2_25, u0_R2_28, u0_R2_3, u0_R2_32, u0_R2_4, u0_R2_5, u0_R2_6, u0_R2_7, 
       u0_R2_8, u0_R2_9, u0_R3_13, u0_R3_15, u0_R3_17, u0_R3_18, u0_R3_20, u0_R3_22, u0_R3_24, 
       u0_R3_25, u0_R3_32, u0_R3_5, u0_R5_12, u0_R5_13, u0_R5_2, u0_R5_25, u0_R5_3, u0_R5_32, 
       u0_R5_4, u0_R5_5, u0_R5_7, u0_R5_8, u0_R5_9, u0_R6_10, u0_R6_11, u0_R6_12, u0_R6_13, 
       u0_R6_14, u0_R6_17, u0_R6_4, u0_R6_5, u0_R6_7, u0_R6_8, u0_R6_9, u0_R8_1, u0_R8_12, 
       u0_R8_13, u0_R8_17, u0_R8_19, u0_R8_20, u0_R8_21, u0_R8_22, u0_R8_27, u0_R8_29, u0_R8_30, 
       u0_R8_32, u0_R8_5, u0_R8_6, u0_R8_9, u0_u12_X_26, u0_u12_X_27, u0_u12_X_28, u0_u12_X_30, u0_u12_X_32, 
       u0_u12_X_33, u0_u12_X_34, u0_u12_X_35, u0_u12_X_36, u0_u13_X_1, u0_u13_X_10, u0_u13_X_11, u0_u13_X_12, u0_u13_X_19, 
       u0_u13_X_2, u0_u13_X_20, u0_u13_X_21, u0_u13_X_22, u0_u13_X_27, u0_u13_X_3, u0_u13_X_30, u0_u13_X_32, u0_u13_X_36, 
       u0_u13_X_38, u0_u13_X_39, u0_u13_X_4, u0_u13_X_40, u0_u13_X_41, u0_u13_X_42, u0_u13_X_6, u0_u13_X_8, u0_u13_X_9, 
       u0_u14_X_25, u0_u14_X_47, u0_u14_X_48, u0_u3_X_22, u0_u3_X_24, u0_u3_X_26, u0_u3_X_27, u0_u3_X_28, u0_u3_X_29, 
       u0_u3_X_31, u0_u3_X_34, u0_u3_X_35, u0_u3_X_37, u0_u3_X_39, u0_u3_X_40, u0_u3_X_42, u0_u3_X_44, u0_u3_X_45, 
       u0_u3_X_46, u0_u4_X_10, u0_u4_X_11, u0_u4_X_12, u0_u4_X_13, u0_u4_X_14, u0_u4_X_15, u0_u4_X_16, u0_u4_X_17, 
       u0_u4_X_19, u0_u4_X_2, u0_u4_X_21, u0_u4_X_23, u0_u4_X_25, u0_u4_X_28, u0_u4_X_3, u0_u4_X_30, u0_u4_X_32, 
       u0_u4_X_34, u0_u4_X_4, u0_u4_X_43, u0_u4_X_44, u0_u4_X_45, u0_u4_X_46, u0_u4_X_48, u0_u4_X_5, u0_u4_X_7, 
       u0_u4_X_9, u0_u6_X_15, u0_u6_X_16, u0_u6_X_2, u0_u6_X_21, u0_u6_X_22, u0_u6_X_23, u0_u6_X_24, u0_u6_X_31, 
       u0_u6_X_32, u0_u6_X_33, u0_u6_X_34, u0_u6_X_35, u0_u6_X_9, u0_u7_X_1, u0_u7_X_2, u0_u7_X_22, u0_u7_X_23, 
       u0_u7_X_3, u0_u7_X_4, u0_u7_X_9, u0_u9_X_10, u0_u9_X_11, u0_u9_X_13, u0_u9_X_15, u0_u9_X_16, u0_u9_X_21, 
       u0_u9_X_22, u0_u9_X_23, u0_u9_X_25, u0_u9_X_27, u0_u9_X_3, u0_u9_X_34, u0_u9_X_35, u0_u9_X_36, u0_u9_X_37, 
       u0_u9_X_38, u0_u9_X_39, u0_u9_X_4, u0_u9_X_41, u0_u9_X_43, u0_u9_X_46, u0_u9_X_5, u0_u9_X_7, u0_uk_K_r13_0, 
       u0_uk_K_r13_38, u0_uk_K_r13_44, u0_uk_K_r2_13, u0_uk_K_r2_18, u0_uk_K_r2_20, u0_uk_K_r2_25, u0_uk_K_r2_26, u0_uk_K_r2_27, u0_uk_K_r2_28, 
       u0_uk_K_r2_33, u0_uk_K_r2_4, u0_uk_K_r2_41, u0_uk_K_r2_46, u0_uk_K_r2_50, u0_uk_K_r2_53, u0_uk_K_r2_55, u0_uk_K_r3_10, u0_uk_K_r3_14, 
       u0_uk_K_r5_10, u0_uk_K_r5_17, u0_uk_K_r5_39, u0_uk_K_r5_4, u0_uk_K_r6_26, u0_uk_K_r6_34, u0_uk_K_r6_46, u0_uk_K_r8_16, u0_uk_K_r8_40, 
       u0_uk_K_r8_41, u0_uk_n10, u0_uk_n100, u0_uk_n1005, u0_uk_n1006, u0_uk_n1012, u0_uk_n102, u0_uk_n1024, u0_uk_n109, 
       u0_uk_n11, u0_uk_n110, u0_uk_n113, u0_uk_n116, u0_uk_n117, u0_uk_n118, u0_uk_n12, u0_uk_n123, u0_uk_n128, 
       u0_uk_n129, u0_uk_n13, u0_uk_n141, u0_uk_n142, u0_uk_n145, u0_uk_n146, u0_uk_n147, u0_uk_n148, u0_uk_n155, 
       u0_uk_n161, u0_uk_n162, u0_uk_n163, u0_uk_n164, u0_uk_n17, u0_uk_n18, u0_uk_n182, u0_uk_n187, u0_uk_n188, 
       u0_uk_n202, u0_uk_n203, u0_uk_n207, u0_uk_n208, u0_uk_n209, u0_uk_n21, u0_uk_n214, u0_uk_n217, u0_uk_n22, 
       u0_uk_n220, u0_uk_n23, u0_uk_n230, u0_uk_n231, u0_uk_n232, u0_uk_n233, u0_uk_n238, u0_uk_n239, u0_uk_n240, 
       u0_uk_n241, u0_uk_n242, u0_uk_n243, u0_uk_n244, u0_uk_n248, u0_uk_n249, u0_uk_n250, u0_uk_n251, u0_uk_n252, 
       u0_uk_n253, u0_uk_n257, u0_uk_n259, u0_uk_n260, u0_uk_n261, u0_uk_n264, u0_uk_n266, u0_uk_n267, u0_uk_n269, 
       u0_uk_n27, u0_uk_n28, u0_uk_n3, u0_uk_n31, u0_uk_n318, u0_uk_n32, u0_uk_n324, u0_uk_n329, u0_uk_n33, 
       u0_uk_n330, u0_uk_n331, u0_uk_n336, u0_uk_n337, u0_uk_n339, u0_uk_n344, u0_uk_n352, u0_uk_n358, u0_uk_n361, 
       u0_uk_n370, u0_uk_n371, u0_uk_n383, u0_uk_n384, u0_uk_n39, u0_uk_n392, u0_uk_n393, u0_uk_n396, u0_uk_n4, 
       u0_uk_n40, u0_uk_n400, u0_uk_n401, u0_uk_n405, u0_uk_n41, u0_uk_n45, u0_uk_n457, u0_uk_n471, u0_uk_n497, 
       u0_uk_n499, u0_uk_n5, u0_uk_n502, u0_uk_n505, u0_uk_n508, u0_uk_n510, u0_uk_n511, u0_uk_n513, u0_uk_n517, 
       u0_uk_n519, u0_uk_n522, u0_uk_n523, u0_uk_n525, u0_uk_n529, u0_uk_n530, u0_uk_n531, u0_uk_n532, u0_uk_n534, 
       u0_uk_n535, u0_uk_n536, u0_uk_n539, u0_uk_n55, u0_uk_n60, u0_uk_n61, u0_uk_n63, u0_uk_n67, u0_uk_n73, 
       u0_uk_n759, u0_uk_n761, u0_uk_n763, u0_uk_n768, u0_uk_n780, u0_uk_n783, u0_uk_n809, u0_uk_n810, u0_uk_n813, 
       u0_uk_n815, u0_uk_n816, u0_uk_n83, u0_uk_n832, u0_uk_n839, u0_uk_n9, u0_uk_n915, u0_uk_n916, u0_uk_n917, 
       u0_uk_n918, u0_uk_n92, u0_uk_n93, u0_uk_n933, u0_uk_n934, u0_uk_n94, u0_uk_n98, u0_uk_n99, u2_K10_1, 
       u2_K10_36, u2_K10_42, u2_K10_43, u2_K10_44, u2_K10_48, u2_K10_5, u2_K11_24, u2_K11_26, u2_K11_29, 
       u2_K12_2, u2_K12_20, u2_K12_25, u2_K12_36, u2_K12_38, u2_K12_47, u2_K12_48, u2_K13_32, u2_K13_35, 
       u2_K13_37, u2_K13_48, u2_K14_38, u2_K15_1, u2_K15_12, u2_K15_17, u2_K15_2, u2_K15_23, u2_K15_29, 
       u2_K15_31, u2_K15_35, u2_K15_44, u2_K1_43, u2_K3_13, u2_K3_19, u2_K3_20, u2_K3_23, u2_K3_26, 
       u2_K3_42, u2_K3_43, u2_K3_47, u2_K3_48, u2_K4_14, u2_K4_18, u2_K4_19, u2_K4_24, u2_K4_48, 
       u2_K4_6, u2_K4_7, u2_K5_11, u2_K5_13, u2_K5_14, u2_K5_17, u2_K5_18, u2_K5_19, u2_K5_2, 
       u2_K5_23, u2_K5_24, u2_K5_25, u2_K5_26, u2_K5_29, u2_K5_30, u2_K5_31, u2_K5_32, u2_K5_37, 
       u2_K5_38, u2_K5_41, u2_K5_44, u2_K5_48, u2_K5_5, u2_K5_6, u2_K5_8, u2_K6_1, u2_K6_11, 
       u2_K6_13, u2_K6_14, u2_K6_19, u2_K6_20, u2_K6_24, u2_K6_32, u2_K6_47, u2_K6_6, u2_K6_8, 
       u2_K7_26, u2_K7_30, u2_K7_31, u2_K7_35, u2_K7_37, u2_K7_38, u2_K7_43, u2_K7_48, u2_K7_5, 
       u2_K7_7, u2_K9_12, u2_K9_14, u2_K9_23, u2_K9_25, u2_K9_5, u2_R10_1, u2_R10_12, u2_R10_13, 
       u2_R10_16, u2_R10_21, u2_R10_25, u2_R10_29, u2_R10_3, u2_R10_32, u2_R10_4, u2_R10_7, u2_R10_8, 
       u2_R10_9, u2_R11_1, u2_R11_21, u2_R11_24, u2_R11_4, u2_R12_20, u2_R12_21, u2_R12_22, u2_R12_25, 
       u2_R13_1, u2_R13_12, u2_R13_16, u2_R13_17, u2_R13_20, u2_R13_22, u2_R13_24, u2_R13_25, u2_R13_27, 
       u2_R13_29, u2_R13_32, u2_R13_5, u2_R13_9, u2_R1_1, u2_R1_12, u2_R1_13, u2_R1_14, u2_R1_15, 
       u2_R1_16, u2_R1_17, u2_R1_2, u2_R1_25, u2_R1_27, u2_R1_28, u2_R1_29, u2_R1_3, u2_R1_30, 
       u2_R1_31, u2_R1_32, u2_R1_5, u2_R1_6, u2_R1_7, u2_R1_8, u2_R1_9, u2_R2_1, u2_R2_10, 
       u2_R2_11, u2_R2_12, u2_R2_13, u2_R2_16, u2_R2_17, u2_R2_19, u2_R2_2, u2_R2_20, u2_R2_21, 
       u2_R2_25, u2_R2_3, u2_R2_32, u2_R2_4, u2_R2_5, u2_R2_6, u2_R2_7, u2_R2_8, u2_R2_9, 
       u2_R3_1, u2_R3_12, u2_R3_13, u2_R3_16, u2_R3_17, u2_R3_18, u2_R3_20, u2_R3_21, u2_R3_22, 
       u2_R3_24, u2_R3_25, u2_R3_28, u2_R3_29, u2_R3_30, u2_R3_4, u2_R3_5, u2_R3_8, u2_R3_9, 
       u2_R4_1, u2_R4_12, u2_R4_13, u2_R4_14, u2_R4_17, u2_R4_21, u2_R4_22, u2_R4_24, u2_R4_28, 
       u2_R4_29, u2_R4_31, u2_R4_32, u2_R4_4, u2_R4_5, u2_R4_6, u2_R4_8, u2_R4_9, u2_R5_1, 
       u2_R5_10, u2_R5_11, u2_R5_12, u2_R5_13, u2_R5_14, u2_R5_16, u2_R5_17, u2_R5_20, u2_R5_21, 
       u2_R5_23, u2_R5_24, u2_R5_25, u2_R5_26, u2_R5_28, u2_R5_29, u2_R5_32, u2_R5_4, u2_R5_5, 
       u2_R5_8, u2_R5_9, u2_R7_1, u2_R7_11, u2_R7_12, u2_R7_13, u2_R7_14, u2_R7_15, u2_R7_16, 
       u2_R7_17, u2_R7_3, u2_R7_4, u2_R7_5, u2_R7_6, u2_R7_7, u2_R7_8, u2_R7_9, u2_R8_1, 
       u2_R8_20, u2_R8_22, u2_R8_24, u2_R8_25, u2_R8_26, u2_R8_27, u2_R8_28, u2_R8_29, u2_R8_32, 
       u2_R8_4, u2_R9_12, u2_R9_13, u2_R9_17, u2_R9_20, u2_R9_32, u2_desIn_r_1, u2_desIn_r_25, u2_desIn_r_27, 
       u2_desIn_r_33, u2_desIn_r_57, u2_key_r_14, u2_key_r_23, u2_key_r_30, u2_key_r_7, u2_u0_X_10, u2_u0_X_11, u2_u0_X_12, 
       u2_u0_X_25, u2_u0_X_26, u2_u0_X_27, u2_u0_X_28, u2_u0_X_30, u2_u0_X_32, u2_u0_X_33, u2_u0_X_34, u2_u0_X_35, 
       u2_u0_X_37, u2_u0_X_39, u2_u0_X_40, u2_u0_X_45, u2_u0_X_46, u2_u0_X_48, u2_u0_X_7, u2_u0_X_8, u2_u0_X_9, 
       u2_u10_X_21, u2_u10_X_22, u2_u10_X_23, u2_u10_X_25, u2_u10_X_27, u2_u10_X_28, u2_u10_X_30, u2_u10_X_32, u2_u10_X_33, 
       u2_u10_X_34, u2_u10_X_35, u2_u10_X_36, u2_u10_X_37, u2_u10_X_38, u2_u10_X_39, u2_u10_X_40, u2_u10_X_41, u2_u10_X_42, 
       u2_u10_X_43, u2_u10_X_44, u2_u10_X_45, u2_u10_X_46, u2_u10_X_48, u2_u11_X_15, u2_u11_X_16, u2_u11_X_21, u2_u11_X_22, 
       u2_u11_X_24, u2_u11_X_26, u2_u11_X_27, u2_u11_X_28, u2_u11_X_29, u2_u11_X_3, u2_u11_X_31, u2_u11_X_33, u2_u11_X_34, 
       u2_u11_X_35, u2_u11_X_37, u2_u11_X_39, u2_u11_X_40, u2_u11_X_41, u2_u11_X_43, u2_u11_X_45, u2_u11_X_46, u2_u11_X_6, 
       u2_u11_X_8, u2_u11_X_9, u2_u12_X_1, u2_u12_X_10, u2_u12_X_11, u2_u12_X_12, u2_u12_X_25, u2_u12_X_26, u2_u12_X_27, 
       u2_u12_X_28, u2_u12_X_29, u2_u12_X_3, u2_u12_X_31, u2_u12_X_33, u2_u12_X_34, u2_u12_X_36, u2_u12_X_38, u2_u12_X_39, 
       u2_u12_X_4, u2_u12_X_40, u2_u12_X_41, u2_u12_X_42, u2_u12_X_43, u2_u12_X_44, u2_u12_X_45, u2_u12_X_46, u2_u12_X_47, 
       u2_u12_X_6, u2_u12_X_8, u2_u12_X_9, u2_u13_X_25, u2_u13_X_26, u2_u13_X_27, u2_u13_X_28, u2_u13_X_34, u2_u13_X_35, 
       u2_u13_X_37, u2_u13_X_39, u2_u13_X_40, u2_u13_X_41, u2_u13_X_42, u2_u13_X_43, u2_u13_X_44, u2_u13_X_45, u2_u13_X_46, 
       u2_u13_X_47, u2_u13_X_48, u2_u14_X_10, u2_u14_X_11, u2_u14_X_13, u2_u14_X_15, u2_u14_X_16, u2_u14_X_18, u2_u14_X_20, 
       u2_u14_X_21, u2_u14_X_22, u2_u14_X_27, u2_u14_X_28, u2_u14_X_3, u2_u14_X_30, u2_u14_X_32, u2_u14_X_34, u2_u14_X_39, 
       u2_u14_X_4, u2_u14_X_41, u2_u14_X_43, u2_u14_X_45, u2_u14_X_46, u2_u14_X_5, u2_u14_X_7, u2_u14_X_9, u2_u2_X_15, 
       u2_u2_X_16, u2_u2_X_27, u2_u2_X_28, u2_u2_X_29, u2_u2_X_30, u2_u2_X_31, u2_u2_X_32, u2_u2_X_33, u2_u2_X_34, 
       u2_u2_X_35, u2_u2_X_37, u2_u2_X_39, u2_u2_X_5, u2_u2_X_7, u2_u3_X_21, u2_u3_X_22, u2_u3_X_27, u2_u3_X_33, 
       u2_u3_X_34, u2_u3_X_35, u2_u3_X_43, u2_u3_X_44, u2_u3_X_45, u2_u3_X_46, u2_u4_X_1, u2_u4_X_10, u2_u4_X_15, 
       u2_u4_X_16, u2_u4_X_21, u2_u4_X_22, u2_u4_X_28, u2_u4_X_3, u2_u4_X_34, u2_u4_X_39, u2_u4_X_4, u2_u4_X_40, 
       u2_u4_X_46, u2_u4_X_47, u2_u4_X_9, u2_u5_X_10, u2_u5_X_15, u2_u5_X_16, u2_u5_X_22, u2_u5_X_23, u2_u5_X_25, 
       u2_u5_X_27, u2_u5_X_28, u2_u5_X_29, u2_u5_X_3, u2_u5_X_31, u2_u5_X_34, u2_u5_X_36, u2_u5_X_38, u2_u5_X_39, 
       u2_u5_X_4, u2_u5_X_40, u2_u5_X_45, u2_u6_X_10, u2_u6_X_22, u2_u6_X_27, u2_u6_X_28, u2_u6_X_3, u2_u6_X_33, 
       u2_u6_X_4, u2_u6_X_40, u2_u6_X_45, u2_u6_X_46, u2_u6_X_9, u2_u8_X_1, u2_u8_X_15, u2_u8_X_27, u2_u8_X_28, 
       u2_u8_X_29, u2_u8_X_3, u2_u8_X_30, u2_u9_X_3, u2_u9_X_32, u2_u9_X_34, u2_u9_X_4, u2_u9_X_45, u2_u9_X_46, 
       u2_u9_X_6, u2_uk_K_r11_28, u2_uk_K_r11_48, u2_uk_K_r11_53, u2_uk_K_r13_22, u2_uk_K_r13_32, u2_uk_K_r1_15, u2_uk_K_r1_16, u2_uk_K_r1_18, 
       u2_uk_K_r1_21, u2_uk_K_r1_22, u2_uk_K_r1_47, u2_uk_K_r2_13, u2_uk_K_r2_18, u2_uk_K_r2_21, u2_uk_K_r2_25, u2_uk_K_r2_27, u2_uk_K_r2_28, 
       u2_uk_K_r2_31, u2_uk_K_r2_36, u2_uk_K_r2_49, u2_uk_K_r2_55, u2_uk_K_r3_11, u2_uk_K_r3_14, u2_uk_K_r3_19, u2_uk_K_r3_43, u2_uk_K_r3_9, 
       u2_uk_K_r4_11, u2_uk_K_r4_17, u2_uk_K_r4_33, u2_uk_K_r4_35, u2_uk_K_r4_38, u2_uk_K_r4_4, u2_uk_K_r4_5, u2_uk_K_r4_55, u2_uk_K_r5_10, 
       u2_uk_K_r5_17, u2_uk_K_r5_19, u2_uk_K_r5_39, u2_uk_K_r5_4, u2_uk_K_r5_41, u2_uk_K_r7_25, u2_uk_K_r7_26, u2_uk_K_r7_32, u2_uk_K_r7_39, 
       u2_uk_K_r7_41, u2_uk_K_r7_48, u2_uk_K_r7_55, u2_uk_K_r8_16, u2_uk_K_r8_2, u2_uk_K_r8_22, u2_uk_K_r8_37, u2_uk_K_r8_41, u2_uk_K_r8_42, 
       u2_uk_K_r9_10, u2_uk_K_r9_4, u2_uk_K_r9_48, u2_uk_n1008, u2_uk_n1020, u2_uk_n1024, u2_uk_n1027, u2_uk_n1028, u2_uk_n1031, 
       u2_uk_n1035, u2_uk_n1038, u2_uk_n1040, u2_uk_n1043, u2_uk_n1046, u2_uk_n1049, u2_uk_n1050, u2_uk_n1053, u2_uk_n1069, 
       u2_uk_n1074, u2_uk_n1076, u2_uk_n1077, u2_uk_n1079, u2_uk_n1082, u2_uk_n1083, u2_uk_n1084, u2_uk_n1088, u2_uk_n1089, 
       u2_uk_n1091, u2_uk_n1093, u2_uk_n1096, u2_uk_n1120, u2_uk_n1123, u2_uk_n1124, u2_uk_n1128, u2_uk_n1130, u2_uk_n1141, 
       u2_uk_n1142, u2_uk_n1152, u2_uk_n1171, u2_uk_n1279, u2_uk_n1280, u2_uk_n1281, u2_uk_n1282, u2_uk_n1283, u2_uk_n1284, 
       u2_uk_n1285, u2_uk_n1286, u2_uk_n1287, u2_uk_n1288, u2_uk_n1290, u2_uk_n1291, u2_uk_n1293, u2_uk_n1295, u2_uk_n1296, 
       u2_uk_n1297, u2_uk_n1300, u2_uk_n1301, u2_uk_n1302, u2_uk_n1305, u2_uk_n1306, u2_uk_n1310, u2_uk_n1311, u2_uk_n1314, 
       u2_uk_n1316, u2_uk_n1317, u2_uk_n1318, u2_uk_n1323, u2_uk_n1324, u2_uk_n1326, u2_uk_n1328, u2_uk_n1329, u2_uk_n1333, 
       u2_uk_n1339, u2_uk_n1341, u2_uk_n1345, u2_uk_n1346, u2_uk_n1350, u2_uk_n1351, u2_uk_n1356, u2_uk_n1359, u2_uk_n1361, 
       u2_uk_n1370, u2_uk_n1375, u2_uk_n1382, u2_uk_n1401, u2_uk_n1405, u2_uk_n1408, u2_uk_n1410, u2_uk_n1413, u2_uk_n1422, 
       u2_uk_n1426, u2_uk_n1428, u2_uk_n1433, u2_uk_n1435, u2_uk_n1438, u2_uk_n1439, u2_uk_n1440, u2_uk_n1441, u2_uk_n1445, 
       u2_uk_n1446, u2_uk_n1447, u2_uk_n1453, u2_uk_n1454, u2_uk_n1456, u2_uk_n1458, u2_uk_n1459, u2_uk_n1462, u2_uk_n1465, 
       u2_uk_n1466, u2_uk_n1470, u2_uk_n1475, u2_uk_n1480, u2_uk_n1486, u2_uk_n1488, u2_uk_n1490, u2_uk_n1493, u2_uk_n1494, 
       u2_uk_n1496, u2_uk_n1497, u2_uk_n1544, u2_uk_n1548, u2_uk_n1549, u2_uk_n1555, u2_uk_n1556, u2_uk_n1563, u2_uk_n1568, 
       u2_uk_n1573, u2_uk_n1580, u2_uk_n1586, u2_uk_n1592, u2_uk_n1594, u2_uk_n1609, u2_uk_n1615, u2_uk_n1622, u2_uk_n1682, 
       u2_uk_n1683, u2_uk_n1688, u2_uk_n1689, u2_uk_n1693, u2_uk_n1708, u2_uk_n1709, u2_uk_n1720, u2_uk_n1721, u2_uk_n1746, 
       u2_uk_n1769, u2_uk_n1770, u2_uk_n1781, u2_uk_n1785, u2_uk_n1797, u2_uk_n1803, u2_uk_n1807, u2_uk_n1808, u2_uk_n1816, 
       u2_uk_n1817, u2_uk_n1819, u2_uk_n1821, u2_uk_n1824, u2_uk_n1826, u2_uk_n1834, u2_uk_n1840, u2_uk_n1846, u2_uk_n1849, 
       u2_uk_n1851, u2_uk_n1852, u2_uk_n1855, u2_uk_n1856, u2_uk_n238, u2_uk_n299, u2_uk_n301, u2_uk_n305, u2_uk_n373, 
       u2_uk_n386, u2_uk_n408, u2_uk_n415, u2_uk_n421, u2_uk_n454, u2_uk_n456, u2_uk_n467, u2_uk_n503, u2_uk_n504, 
       u2_uk_n515, u2_uk_n520, u2_uk_n665, u2_uk_n682, u2_uk_n689, u2_uk_n939, u2_uk_n942, u2_uk_n943, u2_uk_n945, 
       u2_uk_n946, u2_uk_n985, u2_uk_n986, u2_uk_n987, u0_out12_11, u0_out12_14, u0_out12_19, u0_out12_25, u0_out12_29, u0_out12_3, u0_out12_4, u0_out12_8, u0_out13_1, 
        u0_out13_10, u0_out13_11, u0_out13_12, u0_out13_13, u0_out13_14, u0_out13_17, u0_out13_18, u0_out13_19, u0_out13_2, 
        u0_out13_20, u0_out13_22, u0_out13_23, u0_out13_25, u0_out13_26, u0_out13_28, u0_out13_29, u0_out13_3, u0_out13_31, 
        u0_out13_32, u0_out13_4, u0_out13_7, u0_out13_8, u0_out13_9, u0_out14_11, u0_out14_12, u0_out14_14, u0_out14_15, 
        u0_out14_19, u0_out14_21, u0_out14_22, u0_out14_25, u0_out14_27, u0_out14_29, u0_out14_3, u0_out14_32, u0_out14_4, 
        u0_out14_5, u0_out14_7, u0_out14_8, u0_out3_1, u0_out3_10, u0_out3_11, u0_out3_12, u0_out3_13, u0_out3_14, 
        u0_out3_15, u0_out3_16, u0_out3_17, u0_out3_18, u0_out3_19, u0_out3_2, u0_out3_20, u0_out3_21, u0_out3_22, 
        u0_out3_23, u0_out3_24, u0_out3_25, u0_out3_26, u0_out3_27, u0_out3_28, u0_out3_29, u0_out3_3, u0_out3_30, 
        u0_out3_31, u0_out3_32, u0_out3_4, u0_out3_5, u0_out3_6, u0_out3_7, u0_out3_8, u0_out3_9, u0_out4_1, 
        u0_out4_10, u0_out4_11, u0_out4_13, u0_out4_14, u0_out4_15, u0_out4_16, u0_out4_17, u0_out4_18, u0_out4_19, 
        u0_out4_2, u0_out4_20, u0_out4_21, u0_out4_23, u0_out4_24, u0_out4_25, u0_out4_26, u0_out4_27, u0_out4_28, 
        u0_out4_29, u0_out4_3, u0_out4_30, u0_out4_31, u0_out4_4, u0_out4_5, u0_out4_6, u0_out4_8, u0_out4_9, 
        u0_out6_1, u0_out6_10, u0_out6_11, u0_out6_13, u0_out6_16, u0_out6_17, u0_out6_18, u0_out6_19, u0_out6_2, 
        u0_out6_20, u0_out6_23, u0_out6_24, u0_out6_26, u0_out6_28, u0_out6_29, u0_out6_30, u0_out6_31, u0_out6_4, 
        u0_out6_6, u0_out6_9, u0_out7_1, u0_out7_10, u0_out7_13, u0_out7_16, u0_out7_17, u0_out7_18, u0_out7_2, 
        u0_out7_20, u0_out7_23, u0_out7_24, u0_out7_26, u0_out7_28, u0_out7_30, u0_out7_31, u0_out7_6, u0_out7_9, 
        u0_out9_1, u0_out9_10, u0_out9_11, u0_out9_12, u0_out9_13, u0_out9_14, u0_out9_15, u0_out9_16, u0_out9_17, 
        u0_out9_18, u0_out9_19, u0_out9_2, u0_out9_20, u0_out9_21, u0_out9_22, u0_out9_23, u0_out9_24, u0_out9_25, 
        u0_out9_26, u0_out9_27, u0_out9_28, u0_out9_29, u0_out9_3, u0_out9_30, u0_out9_31, u0_out9_32, u0_out9_4, 
        u0_out9_5, u0_out9_6, u0_out9_7, u0_out9_8, u0_out9_9, u0_uk_n213, u0_uk_n223, u2_out0_11, u2_out0_12, 
        u2_out0_13, u2_out0_14, u2_out0_15, u2_out0_18, u2_out0_19, u2_out0_2, u2_out0_21, u2_out0_22, u2_out0_25, 
        u2_out0_27, u2_out0_28, u2_out0_29, u2_out0_3, u2_out0_32, u2_out0_4, u2_out0_5, u2_out0_7, u2_out0_8, 
        u2_out10_1, u2_out10_10, u2_out10_11, u2_out10_12, u2_out10_14, u2_out10_15, u2_out10_19, u2_out10_20, u2_out10_21, 
        u2_out10_22, u2_out10_25, u2_out10_26, u2_out10_27, u2_out10_29, u2_out10_3, u2_out10_32, u2_out10_4, u2_out10_5, 
        u2_out10_7, u2_out10_8, u2_out11_1, u2_out11_10, u2_out11_11, u2_out11_12, u2_out11_13, u2_out11_14, u2_out11_15, 
        u2_out11_16, u2_out11_17, u2_out11_18, u2_out11_19, u2_out11_2, u2_out11_20, u2_out11_21, u2_out11_22, u2_out11_23, 
        u2_out11_24, u2_out11_25, u2_out11_26, u2_out11_27, u2_out11_28, u2_out11_29, u2_out11_3, u2_out11_30, u2_out11_31, 
        u2_out11_32, u2_out11_4, u2_out11_5, u2_out11_6, u2_out11_7, u2_out11_8, u2_out11_9, u2_out12_11, u2_out12_12, 
        u2_out12_13, u2_out12_14, u2_out12_15, u2_out12_17, u2_out12_18, u2_out12_19, u2_out12_2, u2_out12_21, u2_out12_22, 
        u2_out12_23, u2_out12_25, u2_out12_27, u2_out12_28, u2_out12_29, u2_out12_3, u2_out12_31, u2_out12_32, u2_out12_4, 
        u2_out12_5, u2_out12_7, u2_out12_8, u2_out12_9, u2_out13_11, u2_out13_12, u2_out13_14, u2_out13_15, u2_out13_19, 
        u2_out13_21, u2_out13_22, u2_out13_25, u2_out13_27, u2_out13_29, u2_out13_3, u2_out13_32, u2_out13_4, u2_out13_5, 
        u2_out13_7, u2_out13_8, u2_out14_1, u2_out14_10, u2_out14_11, u2_out14_12, u2_out14_13, u2_out14_14, u2_out14_15, 
        u2_out14_16, u2_out14_17, u2_out14_18, u2_out14_19, u2_out14_2, u2_out14_20, u2_out14_21, u2_out14_22, u2_out14_23, 
        u2_out14_24, u2_out14_25, u2_out14_26, u2_out14_27, u2_out14_28, u2_out14_29, u2_out14_3, u2_out14_30, u2_out14_31, 
        u2_out14_32, u2_out14_4, u2_out14_5, u2_out14_6, u2_out14_7, u2_out14_8, u2_out14_9, u2_out2_1, u2_out2_10, 
        u2_out2_11, u2_out2_12, u2_out2_13, u2_out2_14, u2_out2_15, u2_out2_16, u2_out2_17, u2_out2_18, u2_out2_19, 
        u2_out2_2, u2_out2_20, u2_out2_21, u2_out2_22, u2_out2_23, u2_out2_24, u2_out2_25, u2_out2_26, u2_out2_27, 
        u2_out2_28, u2_out2_29, u2_out2_3, u2_out2_30, u2_out2_31, u2_out2_32, u2_out2_4, u2_out2_5, u2_out2_6, 
        u2_out2_7, u2_out2_8, u2_out2_9, u2_out3_1, u2_out3_10, u2_out3_11, u2_out3_13, u2_out3_14, u2_out3_15, 
        u2_out3_16, u2_out3_17, u2_out3_18, u2_out3_19, u2_out3_2, u2_out3_20, u2_out3_21, u2_out3_23, u2_out3_24, 
        u2_out3_25, u2_out3_26, u2_out3_27, u2_out3_28, u2_out3_29, u2_out3_3, u2_out3_30, u2_out3_31, u2_out3_4, 
        u2_out3_5, u2_out3_6, u2_out3_8, u2_out3_9, u2_out4_1, u2_out4_10, u2_out4_11, u2_out4_12, u2_out4_13, 
        u2_out4_14, u2_out4_15, u2_out4_16, u2_out4_17, u2_out4_18, u2_out4_19, u2_out4_2, u2_out4_20, u2_out4_21, 
        u2_out4_22, u2_out4_23, u2_out4_24, u2_out4_25, u2_out4_26, u2_out4_27, u2_out4_28, u2_out4_29, u2_out4_3, 
        u2_out4_30, u2_out4_31, u2_out4_32, u2_out4_4, u2_out4_5, u2_out4_6, u2_out4_7, u2_out4_8, u2_out4_9, 
        u2_out5_1, u2_out5_10, u2_out5_11, u2_out5_12, u2_out5_13, u2_out5_14, u2_out5_15, u2_out5_16, u2_out5_17, 
        u2_out5_18, u2_out5_19, u2_out5_2, u2_out5_20, u2_out5_21, u2_out5_22, u2_out5_23, u2_out5_24, u2_out5_25, 
        u2_out5_26, u2_out5_27, u2_out5_28, u2_out5_29, u2_out5_3, u2_out5_30, u2_out5_31, u2_out5_32, u2_out5_4, 
        u2_out5_5, u2_out5_6, u2_out5_7, u2_out5_8, u2_out5_9, u2_out6_1, u2_out6_10, u2_out6_11, u2_out6_12, 
        u2_out6_13, u2_out6_14, u2_out6_15, u2_out6_16, u2_out6_17, u2_out6_18, u2_out6_19, u2_out6_2, u2_out6_20, 
        u2_out6_21, u2_out6_22, u2_out6_23, u2_out6_24, u2_out6_25, u2_out6_26, u2_out6_27, u2_out6_28, u2_out6_29, 
        u2_out6_3, u2_out6_30, u2_out6_31, u2_out6_32, u2_out6_4, u2_out6_5, u2_out6_6, u2_out6_7, u2_out6_8, 
        u2_out6_9, u2_out8_1, u2_out8_10, u2_out8_13, u2_out8_14, u2_out8_16, u2_out8_17, u2_out8_18, u2_out8_2, 
        u2_out8_20, u2_out8_23, u2_out8_24, u2_out8_25, u2_out8_26, u2_out8_28, u2_out8_3, u2_out8_30, u2_out8_31, 
        u2_out8_6, u2_out8_8, u2_out8_9, u2_out9_11, u2_out9_12, u2_out9_15, u2_out9_17, u2_out9_19, u2_out9_21, 
        u2_out9_22, u2_out9_23, u2_out9_27, u2_out9_29, u2_out9_31, u2_out9_32, u2_out9_4, u2_out9_5, u2_out9_7, 
        u2_out9_9, u2_uk_n10, u2_uk_n100, u2_uk_n102, u2_uk_n109, u2_uk_n11, u2_uk_n110, u2_uk_n117, u2_uk_n118, 
        u2_uk_n128, u2_uk_n129, u2_uk_n141, u2_uk_n142, u2_uk_n145, u2_uk_n146, u2_uk_n147, u2_uk_n148, u2_uk_n155, 
        u2_uk_n161, u2_uk_n162, u2_uk_n163, u2_uk_n164, u2_uk_n17, u2_uk_n182, u2_uk_n187, u2_uk_n188, u2_uk_n191, 
        u2_uk_n202, u2_uk_n203, u2_uk_n207, u2_uk_n208, u2_uk_n209, u2_uk_n213, u2_uk_n214, u2_uk_n217, u2_uk_n220, 
        u2_uk_n222, u2_uk_n223, u2_uk_n230, u2_uk_n231, u2_uk_n27, u2_uk_n31, u2_uk_n60, u2_uk_n63, u2_uk_n83, 
        u2_uk_n92, u2_uk_n93, u2_uk_n94, u2_uk_n99 );
  input u0_K10_1, u0_K10_14, u0_K10_17, u0_K10_18, u0_K10_19, u0_K10_20, u0_K10_32, u0_K14_23, u0_K14_24, 
        u0_K14_25, u0_K14_26, u0_K14_29, u0_K14_5, u0_K14_7, u0_K4_36, u0_K4_43, u0_K4_48, u0_K4_6, 
        u0_K5_1, u0_K5_18, u0_K5_24, u0_K5_26, u0_K5_29, u0_K5_31, u0_K5_47, u0_K5_8, u0_K8_11, 
        u0_K8_13, u0_K8_19, u0_R11_16, u0_R11_20, u0_R12_16, u0_R12_17, u0_R12_19, u0_R12_20, u0_R12_22, 
        u0_R12_23, u0_R12_24, u0_R12_4, u0_R13_17, u0_R13_18, u0_R13_19, u0_R13_20, u0_R13_21, u0_R13_22, 
        u0_R13_23, u0_R13_24, u0_R13_25, u0_R13_26, u0_R13_27, u0_R13_28, u0_R13_29, u0_R13_30, u0_R13_31, 
        u0_R2_1, u0_R2_10, u0_R2_11, u0_R2_12, u0_R2_13, u0_R2_14, u0_R2_16, u0_R2_2, u0_R2_21, 
        u0_R2_22, u0_R2_25, u0_R2_28, u0_R2_3, u0_R2_32, u0_R2_4, u0_R2_5, u0_R2_6, u0_R2_7, 
        u0_R2_8, u0_R2_9, u0_R3_13, u0_R3_15, u0_R3_17, u0_R3_18, u0_R3_20, u0_R3_22, u0_R3_24, 
        u0_R3_25, u0_R3_32, u0_R3_5, u0_R5_12, u0_R5_13, u0_R5_2, u0_R5_25, u0_R5_3, u0_R5_32, 
        u0_R5_4, u0_R5_5, u0_R5_7, u0_R5_8, u0_R5_9, u0_R6_10, u0_R6_11, u0_R6_12, u0_R6_13, 
        u0_R6_14, u0_R6_17, u0_R6_4, u0_R6_5, u0_R6_7, u0_R6_8, u0_R6_9, u0_R8_1, u0_R8_12, 
        u0_R8_13, u0_R8_17, u0_R8_19, u0_R8_20, u0_R8_21, u0_R8_22, u0_R8_27, u0_R8_29, u0_R8_30, 
        u0_R8_32, u0_R8_5, u0_R8_6, u0_R8_9, u0_u12_X_26, u0_u12_X_27, u0_u12_X_28, u0_u12_X_30, u0_u12_X_32, 
        u0_u12_X_33, u0_u12_X_34, u0_u12_X_35, u0_u12_X_36, u0_u13_X_1, u0_u13_X_10, u0_u13_X_11, u0_u13_X_12, u0_u13_X_19, 
        u0_u13_X_2, u0_u13_X_20, u0_u13_X_21, u0_u13_X_22, u0_u13_X_27, u0_u13_X_3, u0_u13_X_30, u0_u13_X_32, u0_u13_X_36, 
        u0_u13_X_38, u0_u13_X_39, u0_u13_X_4, u0_u13_X_40, u0_u13_X_41, u0_u13_X_42, u0_u13_X_6, u0_u13_X_8, u0_u13_X_9, 
        u0_u14_X_25, u0_u14_X_47, u0_u14_X_48, u0_u3_X_22, u0_u3_X_24, u0_u3_X_26, u0_u3_X_27, u0_u3_X_28, u0_u3_X_29, 
        u0_u3_X_31, u0_u3_X_34, u0_u3_X_35, u0_u3_X_37, u0_u3_X_39, u0_u3_X_40, u0_u3_X_42, u0_u3_X_44, u0_u3_X_45, 
        u0_u3_X_46, u0_u4_X_10, u0_u4_X_11, u0_u4_X_12, u0_u4_X_13, u0_u4_X_14, u0_u4_X_15, u0_u4_X_16, u0_u4_X_17, 
        u0_u4_X_19, u0_u4_X_2, u0_u4_X_21, u0_u4_X_23, u0_u4_X_25, u0_u4_X_28, u0_u4_X_3, u0_u4_X_30, u0_u4_X_32, 
        u0_u4_X_34, u0_u4_X_4, u0_u4_X_43, u0_u4_X_44, u0_u4_X_45, u0_u4_X_46, u0_u4_X_48, u0_u4_X_5, u0_u4_X_7, 
        u0_u4_X_9, u0_u6_X_15, u0_u6_X_16, u0_u6_X_2, u0_u6_X_21, u0_u6_X_22, u0_u6_X_23, u0_u6_X_24, u0_u6_X_31, 
        u0_u6_X_32, u0_u6_X_33, u0_u6_X_34, u0_u6_X_35, u0_u6_X_9, u0_u7_X_1, u0_u7_X_2, u0_u7_X_22, u0_u7_X_23, 
        u0_u7_X_3, u0_u7_X_4, u0_u7_X_9, u0_u9_X_10, u0_u9_X_11, u0_u9_X_13, u0_u9_X_15, u0_u9_X_16, u0_u9_X_21, 
        u0_u9_X_22, u0_u9_X_23, u0_u9_X_25, u0_u9_X_27, u0_u9_X_3, u0_u9_X_34, u0_u9_X_35, u0_u9_X_36, u0_u9_X_37, 
        u0_u9_X_38, u0_u9_X_39, u0_u9_X_4, u0_u9_X_41, u0_u9_X_43, u0_u9_X_46, u0_u9_X_5, u0_u9_X_7, u0_uk_K_r13_0, 
        u0_uk_K_r13_38, u0_uk_K_r13_44, u0_uk_K_r2_13, u0_uk_K_r2_18, u0_uk_K_r2_20, u0_uk_K_r2_25, u0_uk_K_r2_26, u0_uk_K_r2_27, u0_uk_K_r2_28, 
        u0_uk_K_r2_33, u0_uk_K_r2_4, u0_uk_K_r2_41, u0_uk_K_r2_46, u0_uk_K_r2_50, u0_uk_K_r2_53, u0_uk_K_r2_55, u0_uk_K_r3_10, u0_uk_K_r3_14, 
        u0_uk_K_r5_10, u0_uk_K_r5_17, u0_uk_K_r5_39, u0_uk_K_r5_4, u0_uk_K_r6_26, u0_uk_K_r6_34, u0_uk_K_r6_46, u0_uk_K_r8_16, u0_uk_K_r8_40, 
        u0_uk_K_r8_41, u0_uk_n10, u0_uk_n100, u0_uk_n1005, u0_uk_n1006, u0_uk_n1012, u0_uk_n102, u0_uk_n1024, u0_uk_n109, 
        u0_uk_n11, u0_uk_n110, u0_uk_n113, u0_uk_n116, u0_uk_n117, u0_uk_n118, u0_uk_n12, u0_uk_n123, u0_uk_n128, 
        u0_uk_n129, u0_uk_n13, u0_uk_n141, u0_uk_n142, u0_uk_n145, u0_uk_n146, u0_uk_n147, u0_uk_n148, u0_uk_n155, 
        u0_uk_n161, u0_uk_n162, u0_uk_n163, u0_uk_n164, u0_uk_n17, u0_uk_n18, u0_uk_n182, u0_uk_n187, u0_uk_n188, 
        u0_uk_n202, u0_uk_n203, u0_uk_n207, u0_uk_n208, u0_uk_n209, u0_uk_n21, u0_uk_n214, u0_uk_n217, u0_uk_n22, 
        u0_uk_n220, u0_uk_n23, u0_uk_n230, u0_uk_n231, u0_uk_n232, u0_uk_n233, u0_uk_n238, u0_uk_n239, u0_uk_n240, 
        u0_uk_n241, u0_uk_n242, u0_uk_n243, u0_uk_n244, u0_uk_n248, u0_uk_n249, u0_uk_n250, u0_uk_n251, u0_uk_n252, 
        u0_uk_n253, u0_uk_n257, u0_uk_n259, u0_uk_n260, u0_uk_n261, u0_uk_n264, u0_uk_n266, u0_uk_n267, u0_uk_n269, 
        u0_uk_n27, u0_uk_n28, u0_uk_n3, u0_uk_n31, u0_uk_n318, u0_uk_n32, u0_uk_n324, u0_uk_n329, u0_uk_n33, 
        u0_uk_n330, u0_uk_n331, u0_uk_n336, u0_uk_n337, u0_uk_n339, u0_uk_n344, u0_uk_n352, u0_uk_n358, u0_uk_n361, 
        u0_uk_n370, u0_uk_n371, u0_uk_n383, u0_uk_n384, u0_uk_n39, u0_uk_n392, u0_uk_n393, u0_uk_n396, u0_uk_n4, 
        u0_uk_n40, u0_uk_n400, u0_uk_n401, u0_uk_n405, u0_uk_n41, u0_uk_n45, u0_uk_n457, u0_uk_n471, u0_uk_n497, 
        u0_uk_n499, u0_uk_n5, u0_uk_n502, u0_uk_n505, u0_uk_n508, u0_uk_n510, u0_uk_n511, u0_uk_n513, u0_uk_n517, 
        u0_uk_n519, u0_uk_n522, u0_uk_n523, u0_uk_n525, u0_uk_n529, u0_uk_n530, u0_uk_n531, u0_uk_n532, u0_uk_n534, 
        u0_uk_n535, u0_uk_n536, u0_uk_n539, u0_uk_n55, u0_uk_n60, u0_uk_n61, u0_uk_n63, u0_uk_n67, u0_uk_n73, 
        u0_uk_n759, u0_uk_n761, u0_uk_n763, u0_uk_n768, u0_uk_n780, u0_uk_n783, u0_uk_n809, u0_uk_n810, u0_uk_n813, 
        u0_uk_n815, u0_uk_n816, u0_uk_n83, u0_uk_n832, u0_uk_n839, u0_uk_n9, u0_uk_n915, u0_uk_n916, u0_uk_n917, 
        u0_uk_n918, u0_uk_n92, u0_uk_n93, u0_uk_n933, u0_uk_n934, u0_uk_n94, u0_uk_n98, u0_uk_n99, u2_K10_1, 
        u2_K10_36, u2_K10_42, u2_K10_43, u2_K10_44, u2_K10_48, u2_K10_5, u2_K11_24, u2_K11_26, u2_K11_29, 
        u2_K12_2, u2_K12_20, u2_K12_25, u2_K12_36, u2_K12_38, u2_K12_47, u2_K12_48, u2_K13_32, u2_K13_35, 
        u2_K13_37, u2_K13_48, u2_K14_38, u2_K15_1, u2_K15_12, u2_K15_17, u2_K15_2, u2_K15_23, u2_K15_29, 
        u2_K15_31, u2_K15_35, u2_K15_44, u2_K1_43, u2_K3_13, u2_K3_19, u2_K3_20, u2_K3_23, u2_K3_26, 
        u2_K3_42, u2_K3_43, u2_K3_47, u2_K3_48, u2_K4_14, u2_K4_18, u2_K4_19, u2_K4_24, u2_K4_48, 
        u2_K4_6, u2_K4_7, u2_K5_11, u2_K5_13, u2_K5_14, u2_K5_17, u2_K5_18, u2_K5_19, u2_K5_2, 
        u2_K5_23, u2_K5_24, u2_K5_25, u2_K5_26, u2_K5_29, u2_K5_30, u2_K5_31, u2_K5_32, u2_K5_37, 
        u2_K5_38, u2_K5_41, u2_K5_44, u2_K5_48, u2_K5_5, u2_K5_6, u2_K5_8, u2_K6_1, u2_K6_11, 
        u2_K6_13, u2_K6_14, u2_K6_19, u2_K6_20, u2_K6_24, u2_K6_32, u2_K6_47, u2_K6_6, u2_K6_8, 
        u2_K7_26, u2_K7_30, u2_K7_31, u2_K7_35, u2_K7_37, u2_K7_38, u2_K7_43, u2_K7_48, u2_K7_5, 
        u2_K7_7, u2_K9_12, u2_K9_14, u2_K9_23, u2_K9_25, u2_K9_5, u2_R10_1, u2_R10_12, u2_R10_13, 
        u2_R10_16, u2_R10_21, u2_R10_25, u2_R10_29, u2_R10_3, u2_R10_32, u2_R10_4, u2_R10_7, u2_R10_8, 
        u2_R10_9, u2_R11_1, u2_R11_21, u2_R11_24, u2_R11_4, u2_R12_20, u2_R12_21, u2_R12_22, u2_R12_25, 
        u2_R13_1, u2_R13_12, u2_R13_16, u2_R13_17, u2_R13_20, u2_R13_22, u2_R13_24, u2_R13_25, u2_R13_27, 
        u2_R13_29, u2_R13_32, u2_R13_5, u2_R13_9, u2_R1_1, u2_R1_12, u2_R1_13, u2_R1_14, u2_R1_15, 
        u2_R1_16, u2_R1_17, u2_R1_2, u2_R1_25, u2_R1_27, u2_R1_28, u2_R1_29, u2_R1_3, u2_R1_30, 
        u2_R1_31, u2_R1_32, u2_R1_5, u2_R1_6, u2_R1_7, u2_R1_8, u2_R1_9, u2_R2_1, u2_R2_10, 
        u2_R2_11, u2_R2_12, u2_R2_13, u2_R2_16, u2_R2_17, u2_R2_19, u2_R2_2, u2_R2_20, u2_R2_21, 
        u2_R2_25, u2_R2_3, u2_R2_32, u2_R2_4, u2_R2_5, u2_R2_6, u2_R2_7, u2_R2_8, u2_R2_9, 
        u2_R3_1, u2_R3_12, u2_R3_13, u2_R3_16, u2_R3_17, u2_R3_18, u2_R3_20, u2_R3_21, u2_R3_22, 
        u2_R3_24, u2_R3_25, u2_R3_28, u2_R3_29, u2_R3_30, u2_R3_4, u2_R3_5, u2_R3_8, u2_R3_9, 
        u2_R4_1, u2_R4_12, u2_R4_13, u2_R4_14, u2_R4_17, u2_R4_21, u2_R4_22, u2_R4_24, u2_R4_28, 
        u2_R4_29, u2_R4_31, u2_R4_32, u2_R4_4, u2_R4_5, u2_R4_6, u2_R4_8, u2_R4_9, u2_R5_1, 
        u2_R5_10, u2_R5_11, u2_R5_12, u2_R5_13, u2_R5_14, u2_R5_16, u2_R5_17, u2_R5_20, u2_R5_21, 
        u2_R5_23, u2_R5_24, u2_R5_25, u2_R5_26, u2_R5_28, u2_R5_29, u2_R5_32, u2_R5_4, u2_R5_5, 
        u2_R5_8, u2_R5_9, u2_R7_1, u2_R7_11, u2_R7_12, u2_R7_13, u2_R7_14, u2_R7_15, u2_R7_16, 
        u2_R7_17, u2_R7_3, u2_R7_4, u2_R7_5, u2_R7_6, u2_R7_7, u2_R7_8, u2_R7_9, u2_R8_1, 
        u2_R8_20, u2_R8_22, u2_R8_24, u2_R8_25, u2_R8_26, u2_R8_27, u2_R8_28, u2_R8_29, u2_R8_32, 
        u2_R8_4, u2_R9_12, u2_R9_13, u2_R9_17, u2_R9_20, u2_R9_32, u2_desIn_r_1, u2_desIn_r_25, u2_desIn_r_27, 
        u2_desIn_r_33, u2_desIn_r_57, u2_key_r_14, u2_key_r_23, u2_key_r_30, u2_key_r_7, u2_u0_X_10, u2_u0_X_11, u2_u0_X_12, 
        u2_u0_X_25, u2_u0_X_26, u2_u0_X_27, u2_u0_X_28, u2_u0_X_30, u2_u0_X_32, u2_u0_X_33, u2_u0_X_34, u2_u0_X_35, 
        u2_u0_X_37, u2_u0_X_39, u2_u0_X_40, u2_u0_X_45, u2_u0_X_46, u2_u0_X_48, u2_u0_X_7, u2_u0_X_8, u2_u0_X_9, 
        u2_u10_X_21, u2_u10_X_22, u2_u10_X_23, u2_u10_X_25, u2_u10_X_27, u2_u10_X_28, u2_u10_X_30, u2_u10_X_32, u2_u10_X_33, 
        u2_u10_X_34, u2_u10_X_35, u2_u10_X_36, u2_u10_X_37, u2_u10_X_38, u2_u10_X_39, u2_u10_X_40, u2_u10_X_41, u2_u10_X_42, 
        u2_u10_X_43, u2_u10_X_44, u2_u10_X_45, u2_u10_X_46, u2_u10_X_48, u2_u11_X_15, u2_u11_X_16, u2_u11_X_21, u2_u11_X_22, 
        u2_u11_X_24, u2_u11_X_26, u2_u11_X_27, u2_u11_X_28, u2_u11_X_29, u2_u11_X_3, u2_u11_X_31, u2_u11_X_33, u2_u11_X_34, 
        u2_u11_X_35, u2_u11_X_37, u2_u11_X_39, u2_u11_X_40, u2_u11_X_41, u2_u11_X_43, u2_u11_X_45, u2_u11_X_46, u2_u11_X_6, 
        u2_u11_X_8, u2_u11_X_9, u2_u12_X_1, u2_u12_X_10, u2_u12_X_11, u2_u12_X_12, u2_u12_X_25, u2_u12_X_26, u2_u12_X_27, 
        u2_u12_X_28, u2_u12_X_29, u2_u12_X_3, u2_u12_X_31, u2_u12_X_33, u2_u12_X_34, u2_u12_X_36, u2_u12_X_38, u2_u12_X_39, 
        u2_u12_X_4, u2_u12_X_40, u2_u12_X_41, u2_u12_X_42, u2_u12_X_43, u2_u12_X_44, u2_u12_X_45, u2_u12_X_46, u2_u12_X_47, 
        u2_u12_X_6, u2_u12_X_8, u2_u12_X_9, u2_u13_X_25, u2_u13_X_26, u2_u13_X_27, u2_u13_X_28, u2_u13_X_34, u2_u13_X_35, 
        u2_u13_X_37, u2_u13_X_39, u2_u13_X_40, u2_u13_X_41, u2_u13_X_42, u2_u13_X_43, u2_u13_X_44, u2_u13_X_45, u2_u13_X_46, 
        u2_u13_X_47, u2_u13_X_48, u2_u14_X_10, u2_u14_X_11, u2_u14_X_13, u2_u14_X_15, u2_u14_X_16, u2_u14_X_18, u2_u14_X_20, 
        u2_u14_X_21, u2_u14_X_22, u2_u14_X_27, u2_u14_X_28, u2_u14_X_3, u2_u14_X_30, u2_u14_X_32, u2_u14_X_34, u2_u14_X_39, 
        u2_u14_X_4, u2_u14_X_41, u2_u14_X_43, u2_u14_X_45, u2_u14_X_46, u2_u14_X_5, u2_u14_X_7, u2_u14_X_9, u2_u2_X_15, 
        u2_u2_X_16, u2_u2_X_27, u2_u2_X_28, u2_u2_X_29, u2_u2_X_30, u2_u2_X_31, u2_u2_X_32, u2_u2_X_33, u2_u2_X_34, 
        u2_u2_X_35, u2_u2_X_37, u2_u2_X_39, u2_u2_X_5, u2_u2_X_7, u2_u3_X_21, u2_u3_X_22, u2_u3_X_27, u2_u3_X_33, 
        u2_u3_X_34, u2_u3_X_35, u2_u3_X_43, u2_u3_X_44, u2_u3_X_45, u2_u3_X_46, u2_u4_X_1, u2_u4_X_10, u2_u4_X_15, 
        u2_u4_X_16, u2_u4_X_21, u2_u4_X_22, u2_u4_X_28, u2_u4_X_3, u2_u4_X_34, u2_u4_X_39, u2_u4_X_4, u2_u4_X_40, 
        u2_u4_X_46, u2_u4_X_47, u2_u4_X_9, u2_u5_X_10, u2_u5_X_15, u2_u5_X_16, u2_u5_X_22, u2_u5_X_23, u2_u5_X_25, 
        u2_u5_X_27, u2_u5_X_28, u2_u5_X_29, u2_u5_X_3, u2_u5_X_31, u2_u5_X_34, u2_u5_X_36, u2_u5_X_38, u2_u5_X_39, 
        u2_u5_X_4, u2_u5_X_40, u2_u5_X_45, u2_u6_X_10, u2_u6_X_22, u2_u6_X_27, u2_u6_X_28, u2_u6_X_3, u2_u6_X_33, 
        u2_u6_X_4, u2_u6_X_40, u2_u6_X_45, u2_u6_X_46, u2_u6_X_9, u2_u8_X_1, u2_u8_X_15, u2_u8_X_27, u2_u8_X_28, 
        u2_u8_X_29, u2_u8_X_3, u2_u8_X_30, u2_u9_X_3, u2_u9_X_32, u2_u9_X_34, u2_u9_X_4, u2_u9_X_45, u2_u9_X_46, 
        u2_u9_X_6, u2_uk_K_r11_28, u2_uk_K_r11_48, u2_uk_K_r11_53, u2_uk_K_r13_22, u2_uk_K_r13_32, u2_uk_K_r1_15, u2_uk_K_r1_16, u2_uk_K_r1_18, 
        u2_uk_K_r1_21, u2_uk_K_r1_22, u2_uk_K_r1_47, u2_uk_K_r2_13, u2_uk_K_r2_18, u2_uk_K_r2_21, u2_uk_K_r2_25, u2_uk_K_r2_27, u2_uk_K_r2_28, 
        u2_uk_K_r2_31, u2_uk_K_r2_36, u2_uk_K_r2_49, u2_uk_K_r2_55, u2_uk_K_r3_11, u2_uk_K_r3_14, u2_uk_K_r3_19, u2_uk_K_r3_43, u2_uk_K_r3_9, 
        u2_uk_K_r4_11, u2_uk_K_r4_17, u2_uk_K_r4_33, u2_uk_K_r4_35, u2_uk_K_r4_38, u2_uk_K_r4_4, u2_uk_K_r4_5, u2_uk_K_r4_55, u2_uk_K_r5_10, 
        u2_uk_K_r5_17, u2_uk_K_r5_19, u2_uk_K_r5_39, u2_uk_K_r5_4, u2_uk_K_r5_41, u2_uk_K_r7_25, u2_uk_K_r7_26, u2_uk_K_r7_32, u2_uk_K_r7_39, 
        u2_uk_K_r7_41, u2_uk_K_r7_48, u2_uk_K_r7_55, u2_uk_K_r8_16, u2_uk_K_r8_2, u2_uk_K_r8_22, u2_uk_K_r8_37, u2_uk_K_r8_41, u2_uk_K_r8_42, 
        u2_uk_K_r9_10, u2_uk_K_r9_4, u2_uk_K_r9_48, u2_uk_n1008, u2_uk_n1020, u2_uk_n1024, u2_uk_n1027, u2_uk_n1028, u2_uk_n1031, 
        u2_uk_n1035, u2_uk_n1038, u2_uk_n1040, u2_uk_n1043, u2_uk_n1046, u2_uk_n1049, u2_uk_n1050, u2_uk_n1053, u2_uk_n1069, 
        u2_uk_n1074, u2_uk_n1076, u2_uk_n1077, u2_uk_n1079, u2_uk_n1082, u2_uk_n1083, u2_uk_n1084, u2_uk_n1088, u2_uk_n1089, 
        u2_uk_n1091, u2_uk_n1093, u2_uk_n1096, u2_uk_n1120, u2_uk_n1123, u2_uk_n1124, u2_uk_n1128, u2_uk_n1130, u2_uk_n1141, 
        u2_uk_n1142, u2_uk_n1152, u2_uk_n1171, u2_uk_n1279, u2_uk_n1280, u2_uk_n1281, u2_uk_n1282, u2_uk_n1283, u2_uk_n1284, 
        u2_uk_n1285, u2_uk_n1286, u2_uk_n1287, u2_uk_n1288, u2_uk_n1290, u2_uk_n1291, u2_uk_n1293, u2_uk_n1295, u2_uk_n1296, 
        u2_uk_n1297, u2_uk_n1300, u2_uk_n1301, u2_uk_n1302, u2_uk_n1305, u2_uk_n1306, u2_uk_n1310, u2_uk_n1311, u2_uk_n1314, 
        u2_uk_n1316, u2_uk_n1317, u2_uk_n1318, u2_uk_n1323, u2_uk_n1324, u2_uk_n1326, u2_uk_n1328, u2_uk_n1329, u2_uk_n1333, 
        u2_uk_n1339, u2_uk_n1341, u2_uk_n1345, u2_uk_n1346, u2_uk_n1350, u2_uk_n1351, u2_uk_n1356, u2_uk_n1359, u2_uk_n1361, 
        u2_uk_n1370, u2_uk_n1375, u2_uk_n1382, u2_uk_n1401, u2_uk_n1405, u2_uk_n1408, u2_uk_n1410, u2_uk_n1413, u2_uk_n1422, 
        u2_uk_n1426, u2_uk_n1428, u2_uk_n1433, u2_uk_n1435, u2_uk_n1438, u2_uk_n1439, u2_uk_n1440, u2_uk_n1441, u2_uk_n1445, 
        u2_uk_n1446, u2_uk_n1447, u2_uk_n1453, u2_uk_n1454, u2_uk_n1456, u2_uk_n1458, u2_uk_n1459, u2_uk_n1462, u2_uk_n1465, 
        u2_uk_n1466, u2_uk_n1470, u2_uk_n1475, u2_uk_n1480, u2_uk_n1486, u2_uk_n1488, u2_uk_n1490, u2_uk_n1493, u2_uk_n1494, 
        u2_uk_n1496, u2_uk_n1497, u2_uk_n1544, u2_uk_n1548, u2_uk_n1549, u2_uk_n1555, u2_uk_n1556, u2_uk_n1563, u2_uk_n1568, 
        u2_uk_n1573, u2_uk_n1580, u2_uk_n1586, u2_uk_n1592, u2_uk_n1594, u2_uk_n1609, u2_uk_n1615, u2_uk_n1622, u2_uk_n1682, 
        u2_uk_n1683, u2_uk_n1688, u2_uk_n1689, u2_uk_n1693, u2_uk_n1708, u2_uk_n1709, u2_uk_n1720, u2_uk_n1721, u2_uk_n1746, 
        u2_uk_n1769, u2_uk_n1770, u2_uk_n1781, u2_uk_n1785, u2_uk_n1797, u2_uk_n1803, u2_uk_n1807, u2_uk_n1808, u2_uk_n1816, 
        u2_uk_n1817, u2_uk_n1819, u2_uk_n1821, u2_uk_n1824, u2_uk_n1826, u2_uk_n1834, u2_uk_n1840, u2_uk_n1846, u2_uk_n1849, 
        u2_uk_n1851, u2_uk_n1852, u2_uk_n1855, u2_uk_n1856, u2_uk_n238, u2_uk_n299, u2_uk_n301, u2_uk_n305, u2_uk_n373, 
        u2_uk_n386, u2_uk_n408, u2_uk_n415, u2_uk_n421, u2_uk_n454, u2_uk_n456, u2_uk_n467, u2_uk_n503, u2_uk_n504, 
        u2_uk_n515, u2_uk_n520, u2_uk_n665, u2_uk_n682, u2_uk_n689, u2_uk_n939, u2_uk_n942, u2_uk_n943, u2_uk_n945, 
        u2_uk_n946, u2_uk_n985, u2_uk_n986, u2_uk_n987;
  output u0_out12_11, u0_out12_14, u0_out12_19, u0_out12_25, u0_out12_29, u0_out12_3, u0_out12_4, u0_out12_8, u0_out13_1, 
        u0_out13_10, u0_out13_11, u0_out13_12, u0_out13_13, u0_out13_14, u0_out13_17, u0_out13_18, u0_out13_19, u0_out13_2, 
        u0_out13_20, u0_out13_22, u0_out13_23, u0_out13_25, u0_out13_26, u0_out13_28, u0_out13_29, u0_out13_3, u0_out13_31, 
        u0_out13_32, u0_out13_4, u0_out13_7, u0_out13_8, u0_out13_9, u0_out14_11, u0_out14_12, u0_out14_14, u0_out14_15, 
        u0_out14_19, u0_out14_21, u0_out14_22, u0_out14_25, u0_out14_27, u0_out14_29, u0_out14_3, u0_out14_32, u0_out14_4, 
        u0_out14_5, u0_out14_7, u0_out14_8, u0_out3_1, u0_out3_10, u0_out3_11, u0_out3_12, u0_out3_13, u0_out3_14, 
        u0_out3_15, u0_out3_16, u0_out3_17, u0_out3_18, u0_out3_19, u0_out3_2, u0_out3_20, u0_out3_21, u0_out3_22, 
        u0_out3_23, u0_out3_24, u0_out3_25, u0_out3_26, u0_out3_27, u0_out3_28, u0_out3_29, u0_out3_3, u0_out3_30, 
        u0_out3_31, u0_out3_32, u0_out3_4, u0_out3_5, u0_out3_6, u0_out3_7, u0_out3_8, u0_out3_9, u0_out4_1, 
        u0_out4_10, u0_out4_11, u0_out4_13, u0_out4_14, u0_out4_15, u0_out4_16, u0_out4_17, u0_out4_18, u0_out4_19, 
        u0_out4_2, u0_out4_20, u0_out4_21, u0_out4_23, u0_out4_24, u0_out4_25, u0_out4_26, u0_out4_27, u0_out4_28, 
        u0_out4_29, u0_out4_3, u0_out4_30, u0_out4_31, u0_out4_4, u0_out4_5, u0_out4_6, u0_out4_8, u0_out4_9, 
        u0_out6_1, u0_out6_10, u0_out6_11, u0_out6_13, u0_out6_16, u0_out6_17, u0_out6_18, u0_out6_19, u0_out6_2, 
        u0_out6_20, u0_out6_23, u0_out6_24, u0_out6_26, u0_out6_28, u0_out6_29, u0_out6_30, u0_out6_31, u0_out6_4, 
        u0_out6_6, u0_out6_9, u0_out7_1, u0_out7_10, u0_out7_13, u0_out7_16, u0_out7_17, u0_out7_18, u0_out7_2, 
        u0_out7_20, u0_out7_23, u0_out7_24, u0_out7_26, u0_out7_28, u0_out7_30, u0_out7_31, u0_out7_6, u0_out7_9, 
        u0_out9_1, u0_out9_10, u0_out9_11, u0_out9_12, u0_out9_13, u0_out9_14, u0_out9_15, u0_out9_16, u0_out9_17, 
        u0_out9_18, u0_out9_19, u0_out9_2, u0_out9_20, u0_out9_21, u0_out9_22, u0_out9_23, u0_out9_24, u0_out9_25, 
        u0_out9_26, u0_out9_27, u0_out9_28, u0_out9_29, u0_out9_3, u0_out9_30, u0_out9_31, u0_out9_32, u0_out9_4, 
        u0_out9_5, u0_out9_6, u0_out9_7, u0_out9_8, u0_out9_9, u0_uk_n213, u0_uk_n223, u2_out0_11, u2_out0_12, 
        u2_out0_13, u2_out0_14, u2_out0_15, u2_out0_18, u2_out0_19, u2_out0_2, u2_out0_21, u2_out0_22, u2_out0_25, 
        u2_out0_27, u2_out0_28, u2_out0_29, u2_out0_3, u2_out0_32, u2_out0_4, u2_out0_5, u2_out0_7, u2_out0_8, 
        u2_out10_1, u2_out10_10, u2_out10_11, u2_out10_12, u2_out10_14, u2_out10_15, u2_out10_19, u2_out10_20, u2_out10_21, 
        u2_out10_22, u2_out10_25, u2_out10_26, u2_out10_27, u2_out10_29, u2_out10_3, u2_out10_32, u2_out10_4, u2_out10_5, 
        u2_out10_7, u2_out10_8, u2_out11_1, u2_out11_10, u2_out11_11, u2_out11_12, u2_out11_13, u2_out11_14, u2_out11_15, 
        u2_out11_16, u2_out11_17, u2_out11_18, u2_out11_19, u2_out11_2, u2_out11_20, u2_out11_21, u2_out11_22, u2_out11_23, 
        u2_out11_24, u2_out11_25, u2_out11_26, u2_out11_27, u2_out11_28, u2_out11_29, u2_out11_3, u2_out11_30, u2_out11_31, 
        u2_out11_32, u2_out11_4, u2_out11_5, u2_out11_6, u2_out11_7, u2_out11_8, u2_out11_9, u2_out12_11, u2_out12_12, 
        u2_out12_13, u2_out12_14, u2_out12_15, u2_out12_17, u2_out12_18, u2_out12_19, u2_out12_2, u2_out12_21, u2_out12_22, 
        u2_out12_23, u2_out12_25, u2_out12_27, u2_out12_28, u2_out12_29, u2_out12_3, u2_out12_31, u2_out12_32, u2_out12_4, 
        u2_out12_5, u2_out12_7, u2_out12_8, u2_out12_9, u2_out13_11, u2_out13_12, u2_out13_14, u2_out13_15, u2_out13_19, 
        u2_out13_21, u2_out13_22, u2_out13_25, u2_out13_27, u2_out13_29, u2_out13_3, u2_out13_32, u2_out13_4, u2_out13_5, 
        u2_out13_7, u2_out13_8, u2_out14_1, u2_out14_10, u2_out14_11, u2_out14_12, u2_out14_13, u2_out14_14, u2_out14_15, 
        u2_out14_16, u2_out14_17, u2_out14_18, u2_out14_19, u2_out14_2, u2_out14_20, u2_out14_21, u2_out14_22, u2_out14_23, 
        u2_out14_24, u2_out14_25, u2_out14_26, u2_out14_27, u2_out14_28, u2_out14_29, u2_out14_3, u2_out14_30, u2_out14_31, 
        u2_out14_32, u2_out14_4, u2_out14_5, u2_out14_6, u2_out14_7, u2_out14_8, u2_out14_9, u2_out2_1, u2_out2_10, 
        u2_out2_11, u2_out2_12, u2_out2_13, u2_out2_14, u2_out2_15, u2_out2_16, u2_out2_17, u2_out2_18, u2_out2_19, 
        u2_out2_2, u2_out2_20, u2_out2_21, u2_out2_22, u2_out2_23, u2_out2_24, u2_out2_25, u2_out2_26, u2_out2_27, 
        u2_out2_28, u2_out2_29, u2_out2_3, u2_out2_30, u2_out2_31, u2_out2_32, u2_out2_4, u2_out2_5, u2_out2_6, 
        u2_out2_7, u2_out2_8, u2_out2_9, u2_out3_1, u2_out3_10, u2_out3_11, u2_out3_13, u2_out3_14, u2_out3_15, 
        u2_out3_16, u2_out3_17, u2_out3_18, u2_out3_19, u2_out3_2, u2_out3_20, u2_out3_21, u2_out3_23, u2_out3_24, 
        u2_out3_25, u2_out3_26, u2_out3_27, u2_out3_28, u2_out3_29, u2_out3_3, u2_out3_30, u2_out3_31, u2_out3_4, 
        u2_out3_5, u2_out3_6, u2_out3_8, u2_out3_9, u2_out4_1, u2_out4_10, u2_out4_11, u2_out4_12, u2_out4_13, 
        u2_out4_14, u2_out4_15, u2_out4_16, u2_out4_17, u2_out4_18, u2_out4_19, u2_out4_2, u2_out4_20, u2_out4_21, 
        u2_out4_22, u2_out4_23, u2_out4_24, u2_out4_25, u2_out4_26, u2_out4_27, u2_out4_28, u2_out4_29, u2_out4_3, 
        u2_out4_30, u2_out4_31, u2_out4_32, u2_out4_4, u2_out4_5, u2_out4_6, u2_out4_7, u2_out4_8, u2_out4_9, 
        u2_out5_1, u2_out5_10, u2_out5_11, u2_out5_12, u2_out5_13, u2_out5_14, u2_out5_15, u2_out5_16, u2_out5_17, 
        u2_out5_18, u2_out5_19, u2_out5_2, u2_out5_20, u2_out5_21, u2_out5_22, u2_out5_23, u2_out5_24, u2_out5_25, 
        u2_out5_26, u2_out5_27, u2_out5_28, u2_out5_29, u2_out5_3, u2_out5_30, u2_out5_31, u2_out5_32, u2_out5_4, 
        u2_out5_5, u2_out5_6, u2_out5_7, u2_out5_8, u2_out5_9, u2_out6_1, u2_out6_10, u2_out6_11, u2_out6_12, 
        u2_out6_13, u2_out6_14, u2_out6_15, u2_out6_16, u2_out6_17, u2_out6_18, u2_out6_19, u2_out6_2, u2_out6_20, 
        u2_out6_21, u2_out6_22, u2_out6_23, u2_out6_24, u2_out6_25, u2_out6_26, u2_out6_27, u2_out6_28, u2_out6_29, 
        u2_out6_3, u2_out6_30, u2_out6_31, u2_out6_32, u2_out6_4, u2_out6_5, u2_out6_6, u2_out6_7, u2_out6_8, 
        u2_out6_9, u2_out8_1, u2_out8_10, u2_out8_13, u2_out8_14, u2_out8_16, u2_out8_17, u2_out8_18, u2_out8_2, 
        u2_out8_20, u2_out8_23, u2_out8_24, u2_out8_25, u2_out8_26, u2_out8_28, u2_out8_3, u2_out8_30, u2_out8_31, 
        u2_out8_6, u2_out8_8, u2_out8_9, u2_out9_11, u2_out9_12, u2_out9_15, u2_out9_17, u2_out9_19, u2_out9_21, 
        u2_out9_22, u2_out9_23, u2_out9_27, u2_out9_29, u2_out9_31, u2_out9_32, u2_out9_4, u2_out9_5, u2_out9_7, 
        u2_out9_9, u2_uk_n10, u2_uk_n100, u2_uk_n102, u2_uk_n109, u2_uk_n11, u2_uk_n110, u2_uk_n117, u2_uk_n118, 
        u2_uk_n128, u2_uk_n129, u2_uk_n141, u2_uk_n142, u2_uk_n145, u2_uk_n146, u2_uk_n147, u2_uk_n148, u2_uk_n155, 
        u2_uk_n161, u2_uk_n162, u2_uk_n163, u2_uk_n164, u2_uk_n17, u2_uk_n182, u2_uk_n187, u2_uk_n188, u2_uk_n191, 
        u2_uk_n202, u2_uk_n203, u2_uk_n207, u2_uk_n208, u2_uk_n209, u2_uk_n213, u2_uk_n214, u2_uk_n217, u2_uk_n220, 
        u2_uk_n222, u2_uk_n223, u2_uk_n230, u2_uk_n231, u2_uk_n27, u2_uk_n31, u2_uk_n60, u2_uk_n63, u2_uk_n83, 
        u2_uk_n92, u2_uk_n93, u2_uk_n94, u2_uk_n99;
  wire u0_K10_12, u0_K10_2, u0_K10_24, u0_K10_26, u0_K10_28, u0_K10_29, u0_K10_30, u0_K10_31, u0_K10_33, 
       u0_K10_40, u0_K10_42, u0_K10_44, u0_K10_45, u0_K10_47, u0_K10_48, u0_K10_6, u0_K10_8, u0_K10_9, 
       u0_K13_25, u0_K13_29, u0_K13_31, u0_K14_28, u0_K14_31, u0_K14_33, u0_K14_34, u0_K14_35, u0_K14_37, 
       u0_K15_26, u0_K15_27, u0_K15_28, u0_K15_29, u0_K15_30, u0_K15_31, u0_K15_32, u0_K15_33, u0_K15_34, 
       u0_K15_35, u0_K15_36, u0_K15_37, u0_K15_38, u0_K15_39, u0_K15_40, u0_K15_41, u0_K15_42, u0_K15_43, 
       u0_K15_44, u0_K15_45, u0_K15_46, u0_K4_1, u0_K4_10, u0_K4_11, u0_K4_12, u0_K4_13, u0_K4_14, 
       u0_K4_15, u0_K4_16, u0_K4_17, u0_K4_18, u0_K4_19, u0_K4_2, u0_K4_20, u0_K4_21, u0_K4_23, 
       u0_K4_25, u0_K4_3, u0_K4_30, u0_K4_32, u0_K4_33, u0_K4_38, u0_K4_4, u0_K4_41, u0_K4_47, 
       u0_K4_5, u0_K4_7, u0_K4_8, u0_K4_9, u0_K5_20, u0_K5_22, u0_K5_27, u0_K5_33, u0_K5_35, 
       u0_K5_36, u0_K5_6, u0_K7_1, u0_K7_10, u0_K7_11, u0_K7_12, u0_K7_13, u0_K7_14, u0_K7_17, 
       u0_K7_18, u0_K7_19, u0_K7_20, u0_K7_3, u0_K7_36, u0_K7_4, u0_K7_5, u0_K7_6, u0_K7_7, 
       u0_K7_8, u0_K8_10, u0_K8_12, u0_K8_14, u0_K8_15, u0_K8_16, u0_K8_17, u0_K8_18, u0_K8_20, 
       u0_K8_21, u0_K8_24, u0_K8_5, u0_K8_6, u0_K8_7, u0_K8_8, u0_u12_X_25, u0_u12_X_29, u0_u12_X_31, 
       u0_u12_u4_n100, u0_u12_u4_n101, u0_u12_u4_n102, u0_u12_u4_n103, u0_u12_u4_n104, u0_u12_u4_n105, u0_u12_u4_n106, u0_u12_u4_n107, u0_u12_u4_n108, 
       u0_u12_u4_n109, u0_u12_u4_n110, u0_u12_u4_n111, u0_u12_u4_n112, u0_u12_u4_n113, u0_u12_u4_n114, u0_u12_u4_n115, u0_u12_u4_n116, u0_u12_u4_n117, 
       u0_u12_u4_n118, u0_u12_u4_n119, u0_u12_u4_n120, u0_u12_u4_n121, u0_u12_u4_n122, u0_u12_u4_n123, u0_u12_u4_n124, u0_u12_u4_n125, u0_u12_u4_n126, 
       u0_u12_u4_n127, u0_u12_u4_n128, u0_u12_u4_n129, u0_u12_u4_n130, u0_u12_u4_n131, u0_u12_u4_n132, u0_u12_u4_n133, u0_u12_u4_n134, u0_u12_u4_n135, 
       u0_u12_u4_n136, u0_u12_u4_n137, u0_u12_u4_n138, u0_u12_u4_n139, u0_u12_u4_n140, u0_u12_u4_n141, u0_u12_u4_n142, u0_u12_u4_n143, u0_u12_u4_n144, 
       u0_u12_u4_n145, u0_u12_u4_n146, u0_u12_u4_n147, u0_u12_u4_n148, u0_u12_u4_n149, u0_u12_u4_n150, u0_u12_u4_n151, u0_u12_u4_n152, u0_u12_u4_n153, 
       u0_u12_u4_n154, u0_u12_u4_n155, u0_u12_u4_n156, u0_u12_u4_n157, u0_u12_u4_n158, u0_u12_u4_n159, u0_u12_u4_n160, u0_u12_u4_n161, u0_u12_u4_n162, 
       u0_u12_u4_n163, u0_u12_u4_n164, u0_u12_u4_n165, u0_u12_u4_n166, u0_u12_u4_n167, u0_u12_u4_n168, u0_u12_u4_n169, u0_u12_u4_n170, u0_u12_u4_n171, 
       u0_u12_u4_n172, u0_u12_u4_n173, u0_u12_u4_n174, u0_u12_u4_n175, u0_u12_u4_n176, u0_u12_u4_n177, u0_u12_u4_n178, u0_u12_u4_n179, u0_u12_u4_n180, 
       u0_u12_u4_n181, u0_u12_u4_n182, u0_u12_u4_n183, u0_u12_u4_n184, u0_u12_u4_n185, u0_u12_u4_n186, u0_u12_u4_n94, u0_u12_u4_n95, u0_u12_u4_n96, 
       u0_u12_u4_n97, u0_u12_u4_n98, u0_u12_u4_n99, u0_u12_u5_n100, u0_u12_u5_n101, u0_u12_u5_n102, u0_u12_u5_n103, u0_u12_u5_n104, u0_u12_u5_n105, 
       u0_u12_u5_n106, u0_u12_u5_n107, u0_u12_u5_n108, u0_u12_u5_n109, u0_u12_u5_n110, u0_u12_u5_n111, u0_u12_u5_n112, u0_u12_u5_n113, u0_u12_u5_n114, 
       u0_u12_u5_n115, u0_u12_u5_n116, u0_u12_u5_n117, u0_u12_u5_n118, u0_u12_u5_n119, u0_u12_u5_n120, u0_u12_u5_n121, u0_u12_u5_n122, u0_u12_u5_n123, 
       u0_u12_u5_n124, u0_u12_u5_n125, u0_u12_u5_n126, u0_u12_u5_n127, u0_u12_u5_n128, u0_u12_u5_n129, u0_u12_u5_n130, u0_u12_u5_n131, u0_u12_u5_n132, 
       u0_u12_u5_n133, u0_u12_u5_n134, u0_u12_u5_n135, u0_u12_u5_n136, u0_u12_u5_n137, u0_u12_u5_n138, u0_u12_u5_n139, u0_u12_u5_n140, u0_u12_u5_n141, 
       u0_u12_u5_n142, u0_u12_u5_n143, u0_u12_u5_n144, u0_u12_u5_n145, u0_u12_u5_n146, u0_u12_u5_n147, u0_u12_u5_n148, u0_u12_u5_n149, u0_u12_u5_n150, 
       u0_u12_u5_n151, u0_u12_u5_n152, u0_u12_u5_n153, u0_u12_u5_n154, u0_u12_u5_n155, u0_u12_u5_n156, u0_u12_u5_n157, u0_u12_u5_n158, u0_u12_u5_n159, 
       u0_u12_u5_n160, u0_u12_u5_n161, u0_u12_u5_n162, u0_u12_u5_n163, u0_u12_u5_n164, u0_u12_u5_n165, u0_u12_u5_n166, u0_u12_u5_n167, u0_u12_u5_n168, 
       u0_u12_u5_n169, u0_u12_u5_n170, u0_u12_u5_n171, u0_u12_u5_n172, u0_u12_u5_n173, u0_u12_u5_n174, u0_u12_u5_n175, u0_u12_u5_n176, u0_u12_u5_n177, 
       u0_u12_u5_n178, u0_u12_u5_n179, u0_u12_u5_n180, u0_u12_u5_n181, u0_u12_u5_n182, u0_u12_u5_n183, u0_u12_u5_n184, u0_u12_u5_n185, u0_u12_u5_n186, 
       u0_u12_u5_n187, u0_u12_u5_n188, u0_u12_u5_n189, u0_u12_u5_n190, u0_u12_u5_n191, u0_u12_u5_n192, u0_u12_u5_n193, u0_u12_u5_n194, u0_u12_u5_n195, 
       u0_u12_u5_n196, u0_u12_u5_n99, u0_u13_X_23, u0_u13_X_24, u0_u13_X_25, u0_u13_X_26, u0_u13_X_28, u0_u13_X_29, u0_u13_X_31, 
       u0_u13_X_33, u0_u13_X_34, u0_u13_X_35, u0_u13_X_37, u0_u13_X_5, u0_u13_X_7, u0_u13_u0_n100, u0_u13_u0_n101, u0_u13_u0_n102, 
       u0_u13_u0_n103, u0_u13_u0_n104, u0_u13_u0_n105, u0_u13_u0_n106, u0_u13_u0_n107, u0_u13_u0_n108, u0_u13_u0_n109, u0_u13_u0_n110, u0_u13_u0_n111, 
       u0_u13_u0_n112, u0_u13_u0_n113, u0_u13_u0_n114, u0_u13_u0_n115, u0_u13_u0_n116, u0_u13_u0_n117, u0_u13_u0_n118, u0_u13_u0_n119, u0_u13_u0_n120, 
       u0_u13_u0_n121, u0_u13_u0_n122, u0_u13_u0_n123, u0_u13_u0_n124, u0_u13_u0_n125, u0_u13_u0_n126, u0_u13_u0_n127, u0_u13_u0_n128, u0_u13_u0_n129, 
       u0_u13_u0_n130, u0_u13_u0_n131, u0_u13_u0_n132, u0_u13_u0_n133, u0_u13_u0_n134, u0_u13_u0_n135, u0_u13_u0_n136, u0_u13_u0_n137, u0_u13_u0_n138, 
       u0_u13_u0_n139, u0_u13_u0_n140, u0_u13_u0_n141, u0_u13_u0_n142, u0_u13_u0_n143, u0_u13_u0_n144, u0_u13_u0_n145, u0_u13_u0_n146, u0_u13_u0_n147, 
       u0_u13_u0_n148, u0_u13_u0_n149, u0_u13_u0_n150, u0_u13_u0_n151, u0_u13_u0_n152, u0_u13_u0_n153, u0_u13_u0_n154, u0_u13_u0_n155, u0_u13_u0_n156, 
       u0_u13_u0_n157, u0_u13_u0_n158, u0_u13_u0_n159, u0_u13_u0_n160, u0_u13_u0_n161, u0_u13_u0_n162, u0_u13_u0_n163, u0_u13_u0_n164, u0_u13_u0_n165, 
       u0_u13_u0_n166, u0_u13_u0_n167, u0_u13_u0_n168, u0_u13_u0_n169, u0_u13_u0_n170, u0_u13_u0_n171, u0_u13_u0_n172, u0_u13_u0_n173, u0_u13_u0_n174, 
       u0_u13_u0_n88, u0_u13_u0_n89, u0_u13_u0_n90, u0_u13_u0_n91, u0_u13_u0_n92, u0_u13_u0_n93, u0_u13_u0_n94, u0_u13_u0_n95, u0_u13_u0_n96, 
       u0_u13_u0_n97, u0_u13_u0_n98, u0_u13_u0_n99, u0_u13_u1_n100, u0_u13_u1_n101, u0_u13_u1_n102, u0_u13_u1_n103, u0_u13_u1_n104, u0_u13_u1_n105, 
       u0_u13_u1_n106, u0_u13_u1_n107, u0_u13_u1_n108, u0_u13_u1_n109, u0_u13_u1_n110, u0_u13_u1_n111, u0_u13_u1_n112, u0_u13_u1_n113, u0_u13_u1_n114, 
       u0_u13_u1_n115, u0_u13_u1_n116, u0_u13_u1_n117, u0_u13_u1_n118, u0_u13_u1_n119, u0_u13_u1_n120, u0_u13_u1_n121, u0_u13_u1_n122, u0_u13_u1_n123, 
       u0_u13_u1_n124, u0_u13_u1_n125, u0_u13_u1_n126, u0_u13_u1_n127, u0_u13_u1_n128, u0_u13_u1_n129, u0_u13_u1_n130, u0_u13_u1_n131, u0_u13_u1_n132, 
       u0_u13_u1_n133, u0_u13_u1_n134, u0_u13_u1_n135, u0_u13_u1_n136, u0_u13_u1_n137, u0_u13_u1_n138, u0_u13_u1_n139, u0_u13_u1_n140, u0_u13_u1_n141, 
       u0_u13_u1_n142, u0_u13_u1_n143, u0_u13_u1_n144, u0_u13_u1_n145, u0_u13_u1_n146, u0_u13_u1_n147, u0_u13_u1_n148, u0_u13_u1_n149, u0_u13_u1_n150, 
       u0_u13_u1_n151, u0_u13_u1_n152, u0_u13_u1_n153, u0_u13_u1_n154, u0_u13_u1_n155, u0_u13_u1_n156, u0_u13_u1_n157, u0_u13_u1_n158, u0_u13_u1_n159, 
       u0_u13_u1_n160, u0_u13_u1_n161, u0_u13_u1_n162, u0_u13_u1_n163, u0_u13_u1_n164, u0_u13_u1_n165, u0_u13_u1_n166, u0_u13_u1_n167, u0_u13_u1_n168, 
       u0_u13_u1_n169, u0_u13_u1_n170, u0_u13_u1_n171, u0_u13_u1_n172, u0_u13_u1_n173, u0_u13_u1_n174, u0_u13_u1_n175, u0_u13_u1_n176, u0_u13_u1_n177, 
       u0_u13_u1_n178, u0_u13_u1_n179, u0_u13_u1_n180, u0_u13_u1_n181, u0_u13_u1_n182, u0_u13_u1_n183, u0_u13_u1_n184, u0_u13_u1_n185, u0_u13_u1_n186, 
       u0_u13_u1_n187, u0_u13_u1_n188, u0_u13_u1_n95, u0_u13_u1_n96, u0_u13_u1_n97, u0_u13_u1_n98, u0_u13_u1_n99, u0_u13_u3_n100, u0_u13_u3_n101, 
       u0_u13_u3_n102, u0_u13_u3_n103, u0_u13_u3_n104, u0_u13_u3_n105, u0_u13_u3_n106, u0_u13_u3_n107, u0_u13_u3_n108, u0_u13_u3_n109, u0_u13_u3_n110, 
       u0_u13_u3_n111, u0_u13_u3_n112, u0_u13_u3_n113, u0_u13_u3_n114, u0_u13_u3_n115, u0_u13_u3_n116, u0_u13_u3_n117, u0_u13_u3_n118, u0_u13_u3_n119, 
       u0_u13_u3_n120, u0_u13_u3_n121, u0_u13_u3_n122, u0_u13_u3_n123, u0_u13_u3_n124, u0_u13_u3_n125, u0_u13_u3_n126, u0_u13_u3_n127, u0_u13_u3_n128, 
       u0_u13_u3_n129, u0_u13_u3_n130, u0_u13_u3_n131, u0_u13_u3_n132, u0_u13_u3_n133, u0_u13_u3_n134, u0_u13_u3_n135, u0_u13_u3_n136, u0_u13_u3_n137, 
       u0_u13_u3_n138, u0_u13_u3_n139, u0_u13_u3_n140, u0_u13_u3_n141, u0_u13_u3_n142, u0_u13_u3_n143, u0_u13_u3_n144, u0_u13_u3_n145, u0_u13_u3_n146, 
       u0_u13_u3_n147, u0_u13_u3_n148, u0_u13_u3_n149, u0_u13_u3_n150, u0_u13_u3_n151, u0_u13_u3_n152, u0_u13_u3_n153, u0_u13_u3_n154, u0_u13_u3_n155, 
       u0_u13_u3_n156, u0_u13_u3_n157, u0_u13_u3_n158, u0_u13_u3_n159, u0_u13_u3_n160, u0_u13_u3_n161, u0_u13_u3_n162, u0_u13_u3_n163, u0_u13_u3_n164, 
       u0_u13_u3_n165, u0_u13_u3_n166, u0_u13_u3_n167, u0_u13_u3_n168, u0_u13_u3_n169, u0_u13_u3_n170, u0_u13_u3_n171, u0_u13_u3_n172, u0_u13_u3_n173, 
       u0_u13_u3_n174, u0_u13_u3_n175, u0_u13_u3_n176, u0_u13_u3_n177, u0_u13_u3_n178, u0_u13_u3_n179, u0_u13_u3_n180, u0_u13_u3_n181, u0_u13_u3_n182, 
       u0_u13_u3_n183, u0_u13_u3_n184, u0_u13_u3_n185, u0_u13_u3_n186, u0_u13_u3_n94, u0_u13_u3_n95, u0_u13_u3_n96, u0_u13_u3_n97, u0_u13_u3_n98, 
       u0_u13_u3_n99, u0_u13_u4_n100, u0_u13_u4_n101, u0_u13_u4_n102, u0_u13_u4_n103, u0_u13_u4_n104, u0_u13_u4_n105, u0_u13_u4_n106, u0_u13_u4_n107, 
       u0_u13_u4_n108, u0_u13_u4_n109, u0_u13_u4_n110, u0_u13_u4_n111, u0_u13_u4_n112, u0_u13_u4_n113, u0_u13_u4_n114, u0_u13_u4_n115, u0_u13_u4_n116, 
       u0_u13_u4_n117, u0_u13_u4_n118, u0_u13_u4_n119, u0_u13_u4_n120, u0_u13_u4_n121, u0_u13_u4_n122, u0_u13_u4_n123, u0_u13_u4_n124, u0_u13_u4_n125, 
       u0_u13_u4_n126, u0_u13_u4_n127, u0_u13_u4_n128, u0_u13_u4_n129, u0_u13_u4_n130, u0_u13_u4_n131, u0_u13_u4_n132, u0_u13_u4_n133, u0_u13_u4_n134, 
       u0_u13_u4_n135, u0_u13_u4_n136, u0_u13_u4_n137, u0_u13_u4_n138, u0_u13_u4_n139, u0_u13_u4_n140, u0_u13_u4_n141, u0_u13_u4_n142, u0_u13_u4_n143, 
       u0_u13_u4_n144, u0_u13_u4_n145, u0_u13_u4_n146, u0_u13_u4_n147, u0_u13_u4_n148, u0_u13_u4_n149, u0_u13_u4_n150, u0_u13_u4_n151, u0_u13_u4_n152, 
       u0_u13_u4_n153, u0_u13_u4_n154, u0_u13_u4_n155, u0_u13_u4_n156, u0_u13_u4_n157, u0_u13_u4_n158, u0_u13_u4_n159, u0_u13_u4_n160, u0_u13_u4_n161, 
       u0_u13_u4_n162, u0_u13_u4_n163, u0_u13_u4_n164, u0_u13_u4_n165, u0_u13_u4_n166, u0_u13_u4_n167, u0_u13_u4_n168, u0_u13_u4_n169, u0_u13_u4_n170, 
       u0_u13_u4_n171, u0_u13_u4_n172, u0_u13_u4_n173, u0_u13_u4_n174, u0_u13_u4_n175, u0_u13_u4_n176, u0_u13_u4_n177, u0_u13_u4_n178, u0_u13_u4_n179, 
       u0_u13_u4_n180, u0_u13_u4_n181, u0_u13_u4_n182, u0_u13_u4_n183, u0_u13_u4_n184, u0_u13_u4_n185, u0_u13_u4_n186, u0_u13_u4_n94, u0_u13_u4_n95, 
       u0_u13_u4_n96, u0_u13_u4_n97, u0_u13_u4_n98, u0_u13_u4_n99, u0_u13_u5_n100, u0_u13_u5_n101, u0_u13_u5_n102, u0_u13_u5_n103, u0_u13_u5_n104, 
       u0_u13_u5_n105, u0_u13_u5_n106, u0_u13_u5_n107, u0_u13_u5_n108, u0_u13_u5_n109, u0_u13_u5_n110, u0_u13_u5_n111, u0_u13_u5_n112, u0_u13_u5_n113, 
       u0_u13_u5_n114, u0_u13_u5_n115, u0_u13_u5_n116, u0_u13_u5_n117, u0_u13_u5_n118, u0_u13_u5_n119, u0_u13_u5_n120, u0_u13_u5_n121, u0_u13_u5_n122, 
       u0_u13_u5_n123, u0_u13_u5_n124, u0_u13_u5_n125, u0_u13_u5_n126, u0_u13_u5_n127, u0_u13_u5_n128, u0_u13_u5_n129, u0_u13_u5_n130, u0_u13_u5_n131, 
       u0_u13_u5_n132, u0_u13_u5_n133, u0_u13_u5_n134, u0_u13_u5_n135, u0_u13_u5_n136, u0_u13_u5_n137, u0_u13_u5_n138, u0_u13_u5_n139, u0_u13_u5_n140, 
       u0_u13_u5_n141, u0_u13_u5_n142, u0_u13_u5_n143, u0_u13_u5_n144, u0_u13_u5_n145, u0_u13_u5_n146, u0_u13_u5_n147, u0_u13_u5_n148, u0_u13_u5_n149, 
       u0_u13_u5_n150, u0_u13_u5_n151, u0_u13_u5_n152, u0_u13_u5_n153, u0_u13_u5_n154, u0_u13_u5_n155, u0_u13_u5_n156, u0_u13_u5_n157, u0_u13_u5_n158, 
       u0_u13_u5_n159, u0_u13_u5_n160, u0_u13_u5_n161, u0_u13_u5_n162, u0_u13_u5_n163, u0_u13_u5_n164, u0_u13_u5_n165, u0_u13_u5_n166, u0_u13_u5_n167, 
       u0_u13_u5_n168, u0_u13_u5_n169, u0_u13_u5_n170, u0_u13_u5_n171, u0_u13_u5_n172, u0_u13_u5_n173, u0_u13_u5_n174, u0_u13_u5_n175, u0_u13_u5_n176, 
       u0_u13_u5_n177, u0_u13_u5_n178, u0_u13_u5_n179, u0_u13_u5_n180, u0_u13_u5_n181, u0_u13_u5_n182, u0_u13_u5_n183, u0_u13_u5_n184, u0_u13_u5_n185, 
       u0_u13_u5_n186, u0_u13_u5_n187, u0_u13_u5_n188, u0_u13_u5_n189, u0_u13_u5_n190, u0_u13_u5_n191, u0_u13_u5_n192, u0_u13_u5_n193, u0_u13_u5_n194, 
       u0_u13_u5_n195, u0_u13_u5_n196, u0_u13_u5_n99, u0_u13_u6_n100, u0_u13_u6_n101, u0_u13_u6_n102, u0_u13_u6_n103, u0_u13_u6_n104, u0_u13_u6_n105, 
       u0_u13_u6_n106, u0_u13_u6_n107, u0_u13_u6_n108, u0_u13_u6_n109, u0_u13_u6_n110, u0_u13_u6_n111, u0_u13_u6_n112, u0_u13_u6_n113, u0_u13_u6_n114, 
       u0_u13_u6_n115, u0_u13_u6_n116, u0_u13_u6_n117, u0_u13_u6_n118, u0_u13_u6_n119, u0_u13_u6_n120, u0_u13_u6_n121, u0_u13_u6_n122, u0_u13_u6_n123, 
       u0_u13_u6_n124, u0_u13_u6_n125, u0_u13_u6_n126, u0_u13_u6_n127, u0_u13_u6_n128, u0_u13_u6_n129, u0_u13_u6_n130, u0_u13_u6_n131, u0_u13_u6_n132, 
       u0_u13_u6_n133, u0_u13_u6_n134, u0_u13_u6_n135, u0_u13_u6_n136, u0_u13_u6_n137, u0_u13_u6_n138, u0_u13_u6_n139, u0_u13_u6_n140, u0_u13_u6_n141, 
       u0_u13_u6_n142, u0_u13_u6_n143, u0_u13_u6_n144, u0_u13_u6_n145, u0_u13_u6_n146, u0_u13_u6_n147, u0_u13_u6_n148, u0_u13_u6_n149, u0_u13_u6_n150, 
       u0_u13_u6_n151, u0_u13_u6_n152, u0_u13_u6_n153, u0_u13_u6_n154, u0_u13_u6_n155, u0_u13_u6_n156, u0_u13_u6_n157, u0_u13_u6_n158, u0_u13_u6_n159, 
       u0_u13_u6_n160, u0_u13_u6_n161, u0_u13_u6_n162, u0_u13_u6_n163, u0_u13_u6_n164, u0_u13_u6_n165, u0_u13_u6_n166, u0_u13_u6_n167, u0_u13_u6_n168, 
       u0_u13_u6_n169, u0_u13_u6_n170, u0_u13_u6_n171, u0_u13_u6_n172, u0_u13_u6_n173, u0_u13_u6_n174, u0_u13_u6_n88, u0_u13_u6_n89, u0_u13_u6_n90, 
       u0_u13_u6_n91, u0_u13_u6_n92, u0_u13_u6_n93, u0_u13_u6_n94, u0_u13_u6_n95, u0_u13_u6_n96, u0_u13_u6_n97, u0_u13_u6_n98, u0_u13_u6_n99, 
       u0_u14_X_26, u0_u14_X_27, u0_u14_X_28, u0_u14_X_29, u0_u14_X_30, u0_u14_X_31, u0_u14_X_32, u0_u14_X_33, u0_u14_X_34, 
       u0_u14_X_35, u0_u14_X_36, u0_u14_X_37, u0_u14_X_38, u0_u14_X_39, u0_u14_X_40, u0_u14_X_41, u0_u14_X_42, u0_u14_X_43, 
       u0_u14_X_44, u0_u14_X_45, u0_u14_X_46, u0_u14_u4_n100, u0_u14_u4_n101, u0_u14_u4_n102, u0_u14_u4_n103, u0_u14_u4_n104, u0_u14_u4_n105, 
       u0_u14_u4_n106, u0_u14_u4_n107, u0_u14_u4_n108, u0_u14_u4_n109, u0_u14_u4_n110, u0_u14_u4_n111, u0_u14_u4_n112, u0_u14_u4_n113, u0_u14_u4_n114, 
       u0_u14_u4_n115, u0_u14_u4_n116, u0_u14_u4_n117, u0_u14_u4_n118, u0_u14_u4_n119, u0_u14_u4_n120, u0_u14_u4_n121, u0_u14_u4_n122, u0_u14_u4_n123, 
       u0_u14_u4_n124, u0_u14_u4_n125, u0_u14_u4_n126, u0_u14_u4_n127, u0_u14_u4_n128, u0_u14_u4_n129, u0_u14_u4_n130, u0_u14_u4_n131, u0_u14_u4_n132, 
       u0_u14_u4_n133, u0_u14_u4_n134, u0_u14_u4_n135, u0_u14_u4_n136, u0_u14_u4_n137, u0_u14_u4_n138, u0_u14_u4_n139, u0_u14_u4_n140, u0_u14_u4_n141, 
       u0_u14_u4_n142, u0_u14_u4_n143, u0_u14_u4_n144, u0_u14_u4_n145, u0_u14_u4_n146, u0_u14_u4_n147, u0_u14_u4_n148, u0_u14_u4_n149, u0_u14_u4_n150, 
       u0_u14_u4_n151, u0_u14_u4_n152, u0_u14_u4_n153, u0_u14_u4_n154, u0_u14_u4_n155, u0_u14_u4_n156, u0_u14_u4_n157, u0_u14_u4_n158, u0_u14_u4_n159, 
       u0_u14_u4_n160, u0_u14_u4_n161, u0_u14_u4_n162, u0_u14_u4_n163, u0_u14_u4_n164, u0_u14_u4_n165, u0_u14_u4_n166, u0_u14_u4_n167, u0_u14_u4_n168, 
       u0_u14_u4_n169, u0_u14_u4_n170, u0_u14_u4_n171, u0_u14_u4_n172, u0_u14_u4_n173, u0_u14_u4_n174, u0_u14_u4_n175, u0_u14_u4_n176, u0_u14_u4_n177, 
       u0_u14_u4_n178, u0_u14_u4_n179, u0_u14_u4_n180, u0_u14_u4_n181, u0_u14_u4_n182, u0_u14_u4_n183, u0_u14_u4_n184, u0_u14_u4_n185, u0_u14_u4_n186, 
       u0_u14_u4_n94, u0_u14_u4_n95, u0_u14_u4_n96, u0_u14_u4_n97, u0_u14_u4_n98, u0_u14_u4_n99, u0_u14_u5_n100, u0_u14_u5_n101, u0_u14_u5_n102, 
       u0_u14_u5_n103, u0_u14_u5_n104, u0_u14_u5_n105, u0_u14_u5_n106, u0_u14_u5_n107, u0_u14_u5_n108, u0_u14_u5_n109, u0_u14_u5_n110, u0_u14_u5_n111, 
       u0_u14_u5_n112, u0_u14_u5_n113, u0_u14_u5_n114, u0_u14_u5_n115, u0_u14_u5_n116, u0_u14_u5_n117, u0_u14_u5_n118, u0_u14_u5_n119, u0_u14_u5_n120, 
       u0_u14_u5_n121, u0_u14_u5_n122, u0_u14_u5_n123, u0_u14_u5_n124, u0_u14_u5_n125, u0_u14_u5_n126, u0_u14_u5_n127, u0_u14_u5_n128, u0_u14_u5_n129, 
       u0_u14_u5_n130, u0_u14_u5_n131, u0_u14_u5_n132, u0_u14_u5_n133, u0_u14_u5_n134, u0_u14_u5_n135, u0_u14_u5_n136, u0_u14_u5_n137, u0_u14_u5_n138, 
       u0_u14_u5_n139, u0_u14_u5_n140, u0_u14_u5_n141, u0_u14_u5_n142, u0_u14_u5_n143, u0_u14_u5_n144, u0_u14_u5_n145, u0_u14_u5_n146, u0_u14_u5_n147, 
       u0_u14_u5_n148, u0_u14_u5_n149, u0_u14_u5_n150, u0_u14_u5_n151, u0_u14_u5_n152, u0_u14_u5_n153, u0_u14_u5_n154, u0_u14_u5_n155, u0_u14_u5_n156, 
       u0_u14_u5_n157, u0_u14_u5_n158, u0_u14_u5_n159, u0_u14_u5_n160, u0_u14_u5_n161, u0_u14_u5_n162, u0_u14_u5_n163, u0_u14_u5_n164, u0_u14_u5_n165, 
       u0_u14_u5_n166, u0_u14_u5_n167, u0_u14_u5_n168, u0_u14_u5_n169, u0_u14_u5_n170, u0_u14_u5_n171, u0_u14_u5_n172, u0_u14_u5_n173, u0_u14_u5_n174, 
       u0_u14_u5_n175, u0_u14_u5_n176, u0_u14_u5_n177, u0_u14_u5_n178, u0_u14_u5_n179, u0_u14_u5_n180, u0_u14_u5_n181, u0_u14_u5_n182, u0_u14_u5_n183, 
       u0_u14_u5_n184, u0_u14_u5_n185, u0_u14_u5_n186, u0_u14_u5_n187, u0_u14_u5_n188, u0_u14_u5_n189, u0_u14_u5_n190, u0_u14_u5_n191, u0_u14_u5_n192, 
       u0_u14_u5_n193, u0_u14_u5_n194, u0_u14_u5_n195, u0_u14_u5_n196, u0_u14_u5_n99, u0_u14_u6_n100, u0_u14_u6_n101, u0_u14_u6_n102, u0_u14_u6_n103, 
       u0_u14_u6_n104, u0_u14_u6_n105, u0_u14_u6_n106, u0_u14_u6_n107, u0_u14_u6_n108, u0_u14_u6_n109, u0_u14_u6_n110, u0_u14_u6_n111, u0_u14_u6_n112, 
       u0_u14_u6_n113, u0_u14_u6_n114, u0_u14_u6_n115, u0_u14_u6_n116, u0_u14_u6_n117, u0_u14_u6_n118, u0_u14_u6_n119, u0_u14_u6_n120, u0_u14_u6_n121, 
       u0_u14_u6_n122, u0_u14_u6_n123, u0_u14_u6_n124, u0_u14_u6_n125, u0_u14_u6_n126, u0_u14_u6_n127, u0_u14_u6_n128, u0_u14_u6_n129, u0_u14_u6_n130, 
       u0_u14_u6_n131, u0_u14_u6_n132, u0_u14_u6_n133, u0_u14_u6_n134, u0_u14_u6_n135, u0_u14_u6_n136, u0_u14_u6_n137, u0_u14_u6_n138, u0_u14_u6_n139, 
       u0_u14_u6_n140, u0_u14_u6_n141, u0_u14_u6_n142, u0_u14_u6_n143, u0_u14_u6_n144, u0_u14_u6_n145, u0_u14_u6_n146, u0_u14_u6_n147, u0_u14_u6_n148, 
       u0_u14_u6_n149, u0_u14_u6_n150, u0_u14_u6_n151, u0_u14_u6_n152, u0_u14_u6_n153, u0_u14_u6_n154, u0_u14_u6_n155, u0_u14_u6_n156, u0_u14_u6_n157, 
       u0_u14_u6_n158, u0_u14_u6_n159, u0_u14_u6_n160, u0_u14_u6_n161, u0_u14_u6_n162, u0_u14_u6_n163, u0_u14_u6_n164, u0_u14_u6_n165, u0_u14_u6_n166, 
       u0_u14_u6_n167, u0_u14_u6_n168, u0_u14_u6_n169, u0_u14_u6_n170, u0_u14_u6_n171, u0_u14_u6_n172, u0_u14_u6_n173, u0_u14_u6_n174, u0_u14_u6_n88, 
       u0_u14_u6_n89, u0_u14_u6_n90, u0_u14_u6_n91, u0_u14_u6_n92, u0_u14_u6_n93, u0_u14_u6_n94, u0_u14_u6_n95, u0_u14_u6_n96, u0_u14_u6_n97, 
       u0_u14_u6_n98, u0_u14_u6_n99, u0_u14_u7_n100, u0_u14_u7_n101, u0_u14_u7_n102, u0_u14_u7_n103, u0_u14_u7_n104, u0_u14_u7_n105, u0_u14_u7_n106, 
       u0_u14_u7_n107, u0_u14_u7_n108, u0_u14_u7_n109, u0_u14_u7_n110, u0_u14_u7_n111, u0_u14_u7_n112, u0_u14_u7_n113, u0_u14_u7_n114, u0_u14_u7_n115, 
       u0_u14_u7_n116, u0_u14_u7_n117, u0_u14_u7_n118, u0_u14_u7_n119, u0_u14_u7_n120, u0_u14_u7_n121, u0_u14_u7_n122, u0_u14_u7_n123, u0_u14_u7_n124, 
       u0_u14_u7_n125, u0_u14_u7_n126, u0_u14_u7_n127, u0_u14_u7_n128, u0_u14_u7_n129, u0_u14_u7_n130, u0_u14_u7_n131, u0_u14_u7_n132, u0_u14_u7_n133, 
       u0_u14_u7_n134, u0_u14_u7_n135, u0_u14_u7_n136, u0_u14_u7_n137, u0_u14_u7_n138, u0_u14_u7_n139, u0_u14_u7_n140, u0_u14_u7_n141, u0_u14_u7_n142, 
       u0_u14_u7_n143, u0_u14_u7_n144, u0_u14_u7_n145, u0_u14_u7_n146, u0_u14_u7_n147, u0_u14_u7_n148, u0_u14_u7_n149, u0_u14_u7_n150, u0_u14_u7_n151, 
       u0_u14_u7_n152, u0_u14_u7_n153, u0_u14_u7_n154, u0_u14_u7_n155, u0_u14_u7_n156, u0_u14_u7_n157, u0_u14_u7_n158, u0_u14_u7_n159, u0_u14_u7_n160, 
       u0_u14_u7_n161, u0_u14_u7_n162, u0_u14_u7_n163, u0_u14_u7_n164, u0_u14_u7_n165, u0_u14_u7_n166, u0_u14_u7_n167, u0_u14_u7_n168, u0_u14_u7_n169, 
       u0_u14_u7_n170, u0_u14_u7_n171, u0_u14_u7_n172, u0_u14_u7_n173, u0_u14_u7_n174, u0_u14_u7_n175, u0_u14_u7_n176, u0_u14_u7_n177, u0_u14_u7_n178, 
       u0_u14_u7_n179, u0_u14_u7_n180, u0_u14_u7_n91, u0_u14_u7_n92, u0_u14_u7_n93, u0_u14_u7_n94, u0_u14_u7_n95, u0_u14_u7_n96, u0_u14_u7_n97, 
       u0_u14_u7_n98, u0_u14_u7_n99, u0_u3_X_1, u0_u3_X_10, u0_u3_X_11, u0_u3_X_12, u0_u3_X_13, u0_u3_X_14, u0_u3_X_15, 
       u0_u3_X_16, u0_u3_X_17, u0_u3_X_18, u0_u3_X_19, u0_u3_X_2, u0_u3_X_20, u0_u3_X_21, u0_u3_X_23, u0_u3_X_25, 
       u0_u3_X_3, u0_u3_X_30, u0_u3_X_32, u0_u3_X_33, u0_u3_X_36, u0_u3_X_38, u0_u3_X_4, u0_u3_X_41, u0_u3_X_43, 
       u0_u3_X_47, u0_u3_X_48, u0_u3_X_5, u0_u3_X_6, u0_u3_X_7, u0_u3_X_8, u0_u3_X_9, u0_u3_u0_n100, u0_u3_u0_n101, 
       u0_u3_u0_n102, u0_u3_u0_n103, u0_u3_u0_n104, u0_u3_u0_n105, u0_u3_u0_n106, u0_u3_u0_n107, u0_u3_u0_n108, u0_u3_u0_n109, u0_u3_u0_n110, 
       u0_u3_u0_n111, u0_u3_u0_n112, u0_u3_u0_n113, u0_u3_u0_n114, u0_u3_u0_n115, u0_u3_u0_n116, u0_u3_u0_n117, u0_u3_u0_n118, u0_u3_u0_n119, 
       u0_u3_u0_n120, u0_u3_u0_n121, u0_u3_u0_n122, u0_u3_u0_n123, u0_u3_u0_n124, u0_u3_u0_n125, u0_u3_u0_n126, u0_u3_u0_n127, u0_u3_u0_n128, 
       u0_u3_u0_n129, u0_u3_u0_n130, u0_u3_u0_n131, u0_u3_u0_n132, u0_u3_u0_n133, u0_u3_u0_n134, u0_u3_u0_n135, u0_u3_u0_n136, u0_u3_u0_n137, 
       u0_u3_u0_n138, u0_u3_u0_n139, u0_u3_u0_n140, u0_u3_u0_n141, u0_u3_u0_n142, u0_u3_u0_n143, u0_u3_u0_n144, u0_u3_u0_n145, u0_u3_u0_n146, 
       u0_u3_u0_n147, u0_u3_u0_n148, u0_u3_u0_n149, u0_u3_u0_n150, u0_u3_u0_n151, u0_u3_u0_n152, u0_u3_u0_n153, u0_u3_u0_n154, u0_u3_u0_n155, 
       u0_u3_u0_n156, u0_u3_u0_n157, u0_u3_u0_n158, u0_u3_u0_n159, u0_u3_u0_n160, u0_u3_u0_n161, u0_u3_u0_n162, u0_u3_u0_n163, u0_u3_u0_n164, 
       u0_u3_u0_n165, u0_u3_u0_n166, u0_u3_u0_n167, u0_u3_u0_n168, u0_u3_u0_n169, u0_u3_u0_n170, u0_u3_u0_n171, u0_u3_u0_n172, u0_u3_u0_n173, 
       u0_u3_u0_n174, u0_u3_u0_n175, u0_u3_u0_n176, u0_u3_u0_n88, u0_u3_u0_n89, u0_u3_u0_n90, u0_u3_u0_n91, u0_u3_u0_n92, u0_u3_u0_n93, 
       u0_u3_u0_n94, u0_u3_u0_n95, u0_u3_u0_n96, u0_u3_u0_n97, u0_u3_u0_n98, u0_u3_u0_n99, u0_u3_u1_n100, u0_u3_u1_n101, u0_u3_u1_n102, 
       u0_u3_u1_n103, u0_u3_u1_n104, u0_u3_u1_n105, u0_u3_u1_n106, u0_u3_u1_n107, u0_u3_u1_n108, u0_u3_u1_n109, u0_u3_u1_n110, u0_u3_u1_n111, 
       u0_u3_u1_n112, u0_u3_u1_n113, u0_u3_u1_n114, u0_u3_u1_n115, u0_u3_u1_n116, u0_u3_u1_n117, u0_u3_u1_n118, u0_u3_u1_n119, u0_u3_u1_n120, 
       u0_u3_u1_n121, u0_u3_u1_n122, u0_u3_u1_n123, u0_u3_u1_n124, u0_u3_u1_n125, u0_u3_u1_n126, u0_u3_u1_n127, u0_u3_u1_n128, u0_u3_u1_n129, 
       u0_u3_u1_n130, u0_u3_u1_n131, u0_u3_u1_n132, u0_u3_u1_n133, u0_u3_u1_n134, u0_u3_u1_n135, u0_u3_u1_n136, u0_u3_u1_n137, u0_u3_u1_n138, 
       u0_u3_u1_n139, u0_u3_u1_n140, u0_u3_u1_n141, u0_u3_u1_n142, u0_u3_u1_n143, u0_u3_u1_n144, u0_u3_u1_n145, u0_u3_u1_n146, u0_u3_u1_n147, 
       u0_u3_u1_n148, u0_u3_u1_n149, u0_u3_u1_n150, u0_u3_u1_n151, u0_u3_u1_n152, u0_u3_u1_n153, u0_u3_u1_n154, u0_u3_u1_n155, u0_u3_u1_n156, 
       u0_u3_u1_n157, u0_u3_u1_n158, u0_u3_u1_n159, u0_u3_u1_n160, u0_u3_u1_n161, u0_u3_u1_n162, u0_u3_u1_n163, u0_u3_u1_n164, u0_u3_u1_n165, 
       u0_u3_u1_n166, u0_u3_u1_n167, u0_u3_u1_n168, u0_u3_u1_n169, u0_u3_u1_n170, u0_u3_u1_n171, u0_u3_u1_n172, u0_u3_u1_n173, u0_u3_u1_n174, 
       u0_u3_u1_n175, u0_u3_u1_n176, u0_u3_u1_n177, u0_u3_u1_n178, u0_u3_u1_n179, u0_u3_u1_n180, u0_u3_u1_n181, u0_u3_u1_n182, u0_u3_u1_n183, 
       u0_u3_u1_n184, u0_u3_u1_n185, u0_u3_u1_n186, u0_u3_u1_n187, u0_u3_u1_n188, u0_u3_u1_n95, u0_u3_u1_n96, u0_u3_u1_n97, u0_u3_u1_n98, 
       u0_u3_u1_n99, u0_u3_u2_n100, u0_u3_u2_n101, u0_u3_u2_n102, u0_u3_u2_n103, u0_u3_u2_n104, u0_u3_u2_n105, u0_u3_u2_n106, u0_u3_u2_n107, 
       u0_u3_u2_n108, u0_u3_u2_n109, u0_u3_u2_n110, u0_u3_u2_n111, u0_u3_u2_n112, u0_u3_u2_n113, u0_u3_u2_n114, u0_u3_u2_n115, u0_u3_u2_n116, 
       u0_u3_u2_n117, u0_u3_u2_n118, u0_u3_u2_n119, u0_u3_u2_n120, u0_u3_u2_n121, u0_u3_u2_n122, u0_u3_u2_n123, u0_u3_u2_n124, u0_u3_u2_n125, 
       u0_u3_u2_n126, u0_u3_u2_n127, u0_u3_u2_n128, u0_u3_u2_n129, u0_u3_u2_n130, u0_u3_u2_n131, u0_u3_u2_n132, u0_u3_u2_n133, u0_u3_u2_n134, 
       u0_u3_u2_n135, u0_u3_u2_n136, u0_u3_u2_n137, u0_u3_u2_n138, u0_u3_u2_n139, u0_u3_u2_n140, u0_u3_u2_n141, u0_u3_u2_n142, u0_u3_u2_n143, 
       u0_u3_u2_n144, u0_u3_u2_n145, u0_u3_u2_n146, u0_u3_u2_n147, u0_u3_u2_n148, u0_u3_u2_n149, u0_u3_u2_n150, u0_u3_u2_n151, u0_u3_u2_n152, 
       u0_u3_u2_n153, u0_u3_u2_n154, u0_u3_u2_n155, u0_u3_u2_n156, u0_u3_u2_n157, u0_u3_u2_n158, u0_u3_u2_n159, u0_u3_u2_n160, u0_u3_u2_n161, 
       u0_u3_u2_n162, u0_u3_u2_n163, u0_u3_u2_n164, u0_u3_u2_n165, u0_u3_u2_n166, u0_u3_u2_n167, u0_u3_u2_n168, u0_u3_u2_n169, u0_u3_u2_n170, 
       u0_u3_u2_n171, u0_u3_u2_n172, u0_u3_u2_n173, u0_u3_u2_n174, u0_u3_u2_n175, u0_u3_u2_n176, u0_u3_u2_n177, u0_u3_u2_n178, u0_u3_u2_n179, 
       u0_u3_u2_n180, u0_u3_u2_n181, u0_u3_u2_n182, u0_u3_u2_n183, u0_u3_u2_n184, u0_u3_u2_n185, u0_u3_u2_n186, u0_u3_u2_n187, u0_u3_u2_n188, 
       u0_u3_u2_n95, u0_u3_u2_n96, u0_u3_u2_n97, u0_u3_u2_n98, u0_u3_u2_n99, u0_u3_u3_n100, u0_u3_u3_n101, u0_u3_u3_n102, u0_u3_u3_n103, 
       u0_u3_u3_n104, u0_u3_u3_n105, u0_u3_u3_n106, u0_u3_u3_n107, u0_u3_u3_n108, u0_u3_u3_n109, u0_u3_u3_n110, u0_u3_u3_n111, u0_u3_u3_n112, 
       u0_u3_u3_n113, u0_u3_u3_n114, u0_u3_u3_n115, u0_u3_u3_n116, u0_u3_u3_n117, u0_u3_u3_n118, u0_u3_u3_n119, u0_u3_u3_n120, u0_u3_u3_n121, 
       u0_u3_u3_n122, u0_u3_u3_n123, u0_u3_u3_n124, u0_u3_u3_n125, u0_u3_u3_n126, u0_u3_u3_n127, u0_u3_u3_n128, u0_u3_u3_n129, u0_u3_u3_n130, 
       u0_u3_u3_n131, u0_u3_u3_n132, u0_u3_u3_n133, u0_u3_u3_n134, u0_u3_u3_n135, u0_u3_u3_n136, u0_u3_u3_n137, u0_u3_u3_n138, u0_u3_u3_n139, 
       u0_u3_u3_n140, u0_u3_u3_n141, u0_u3_u3_n142, u0_u3_u3_n143, u0_u3_u3_n144, u0_u3_u3_n145, u0_u3_u3_n146, u0_u3_u3_n147, u0_u3_u3_n148, 
       u0_u3_u3_n149, u0_u3_u3_n150, u0_u3_u3_n151, u0_u3_u3_n152, u0_u3_u3_n153, u0_u3_u3_n154, u0_u3_u3_n155, u0_u3_u3_n156, u0_u3_u3_n157, 
       u0_u3_u3_n158, u0_u3_u3_n159, u0_u3_u3_n160, u0_u3_u3_n161, u0_u3_u3_n162, u0_u3_u3_n163, u0_u3_u3_n164, u0_u3_u3_n165, u0_u3_u3_n166, 
       u0_u3_u3_n167, u0_u3_u3_n168, u0_u3_u3_n169, u0_u3_u3_n170, u0_u3_u3_n171, u0_u3_u3_n172, u0_u3_u3_n173, u0_u3_u3_n174, u0_u3_u3_n175, 
       u0_u3_u3_n176, u0_u3_u3_n177, u0_u3_u3_n178, u0_u3_u3_n179, u0_u3_u3_n180, u0_u3_u3_n181, u0_u3_u3_n182, u0_u3_u3_n183, u0_u3_u3_n184, 
       u0_u3_u3_n185, u0_u3_u3_n186, u0_u3_u3_n94, u0_u3_u3_n95, u0_u3_u3_n96, u0_u3_u3_n97, u0_u3_u3_n98, u0_u3_u3_n99, u0_u3_u4_n100, 
       u0_u3_u4_n101, u0_u3_u4_n102, u0_u3_u4_n103, u0_u3_u4_n104, u0_u3_u4_n105, u0_u3_u4_n106, u0_u3_u4_n107, u0_u3_u4_n108, u0_u3_u4_n109, 
       u0_u3_u4_n110, u0_u3_u4_n111, u0_u3_u4_n112, u0_u3_u4_n113, u0_u3_u4_n114, u0_u3_u4_n115, u0_u3_u4_n116, u0_u3_u4_n117, u0_u3_u4_n118, 
       u0_u3_u4_n119, u0_u3_u4_n120, u0_u3_u4_n121, u0_u3_u4_n122, u0_u3_u4_n123, u0_u3_u4_n124, u0_u3_u4_n125, u0_u3_u4_n126, u0_u3_u4_n127, 
       u0_u3_u4_n128, u0_u3_u4_n129, u0_u3_u4_n130, u0_u3_u4_n131, u0_u3_u4_n132, u0_u3_u4_n133, u0_u3_u4_n134, u0_u3_u4_n135, u0_u3_u4_n136, 
       u0_u3_u4_n137, u0_u3_u4_n138, u0_u3_u4_n139, u0_u3_u4_n140, u0_u3_u4_n141, u0_u3_u4_n142, u0_u3_u4_n143, u0_u3_u4_n144, u0_u3_u4_n145, 
       u0_u3_u4_n146, u0_u3_u4_n147, u0_u3_u4_n148, u0_u3_u4_n149, u0_u3_u4_n150, u0_u3_u4_n151, u0_u3_u4_n152, u0_u3_u4_n153, u0_u3_u4_n154, 
       u0_u3_u4_n155, u0_u3_u4_n156, u0_u3_u4_n157, u0_u3_u4_n158, u0_u3_u4_n159, u0_u3_u4_n160, u0_u3_u4_n161, u0_u3_u4_n162, u0_u3_u4_n163, 
       u0_u3_u4_n164, u0_u3_u4_n165, u0_u3_u4_n166, u0_u3_u4_n167, u0_u3_u4_n168, u0_u3_u4_n169, u0_u3_u4_n170, u0_u3_u4_n171, u0_u3_u4_n172, 
       u0_u3_u4_n173, u0_u3_u4_n174, u0_u3_u4_n175, u0_u3_u4_n176, u0_u3_u4_n177, u0_u3_u4_n178, u0_u3_u4_n179, u0_u3_u4_n180, u0_u3_u4_n181, 
       u0_u3_u4_n182, u0_u3_u4_n183, u0_u3_u4_n184, u0_u3_u4_n185, u0_u3_u4_n186, u0_u3_u4_n94, u0_u3_u4_n95, u0_u3_u4_n96, u0_u3_u4_n97, 
       u0_u3_u4_n98, u0_u3_u4_n99, u0_u3_u5_n100, u0_u3_u5_n101, u0_u3_u5_n102, u0_u3_u5_n103, u0_u3_u5_n104, u0_u3_u5_n105, u0_u3_u5_n106, 
       u0_u3_u5_n107, u0_u3_u5_n108, u0_u3_u5_n109, u0_u3_u5_n110, u0_u3_u5_n111, u0_u3_u5_n112, u0_u3_u5_n113, u0_u3_u5_n114, u0_u3_u5_n115, 
       u0_u3_u5_n116, u0_u3_u5_n117, u0_u3_u5_n118, u0_u3_u5_n119, u0_u3_u5_n120, u0_u3_u5_n121, u0_u3_u5_n122, u0_u3_u5_n123, u0_u3_u5_n124, 
       u0_u3_u5_n125, u0_u3_u5_n126, u0_u3_u5_n127, u0_u3_u5_n128, u0_u3_u5_n129, u0_u3_u5_n130, u0_u3_u5_n131, u0_u3_u5_n132, u0_u3_u5_n133, 
       u0_u3_u5_n134, u0_u3_u5_n135, u0_u3_u5_n136, u0_u3_u5_n137, u0_u3_u5_n138, u0_u3_u5_n139, u0_u3_u5_n140, u0_u3_u5_n141, u0_u3_u5_n142, 
       u0_u3_u5_n143, u0_u3_u5_n144, u0_u3_u5_n145, u0_u3_u5_n146, u0_u3_u5_n147, u0_u3_u5_n148, u0_u3_u5_n149, u0_u3_u5_n150, u0_u3_u5_n151, 
       u0_u3_u5_n152, u0_u3_u5_n153, u0_u3_u5_n154, u0_u3_u5_n155, u0_u3_u5_n156, u0_u3_u5_n157, u0_u3_u5_n158, u0_u3_u5_n159, u0_u3_u5_n160, 
       u0_u3_u5_n161, u0_u3_u5_n162, u0_u3_u5_n163, u0_u3_u5_n164, u0_u3_u5_n165, u0_u3_u5_n166, u0_u3_u5_n167, u0_u3_u5_n168, u0_u3_u5_n169, 
       u0_u3_u5_n170, u0_u3_u5_n171, u0_u3_u5_n172, u0_u3_u5_n173, u0_u3_u5_n174, u0_u3_u5_n175, u0_u3_u5_n176, u0_u3_u5_n177, u0_u3_u5_n178, 
       u0_u3_u5_n179, u0_u3_u5_n180, u0_u3_u5_n181, u0_u3_u5_n182, u0_u3_u5_n183, u0_u3_u5_n184, u0_u3_u5_n185, u0_u3_u5_n186, u0_u3_u5_n187, 
       u0_u3_u5_n188, u0_u3_u5_n189, u0_u3_u5_n190, u0_u3_u5_n191, u0_u3_u5_n192, u0_u3_u5_n193, u0_u3_u5_n194, u0_u3_u5_n195, u0_u3_u5_n196, 
       u0_u3_u5_n99, u0_u3_u6_n100, u0_u3_u6_n101, u0_u3_u6_n102, u0_u3_u6_n103, u0_u3_u6_n104, u0_u3_u6_n105, u0_u3_u6_n106, u0_u3_u6_n107, 
       u0_u3_u6_n108, u0_u3_u6_n109, u0_u3_u6_n110, u0_u3_u6_n111, u0_u3_u6_n112, u0_u3_u6_n113, u0_u3_u6_n114, u0_u3_u6_n115, u0_u3_u6_n116, 
       u0_u3_u6_n117, u0_u3_u6_n118, u0_u3_u6_n119, u0_u3_u6_n120, u0_u3_u6_n121, u0_u3_u6_n122, u0_u3_u6_n123, u0_u3_u6_n124, u0_u3_u6_n125, 
       u0_u3_u6_n126, u0_u3_u6_n127, u0_u3_u6_n128, u0_u3_u6_n129, u0_u3_u6_n130, u0_u3_u6_n131, u0_u3_u6_n132, u0_u3_u6_n133, u0_u3_u6_n134, 
       u0_u3_u6_n135, u0_u3_u6_n136, u0_u3_u6_n137, u0_u3_u6_n138, u0_u3_u6_n139, u0_u3_u6_n140, u0_u3_u6_n141, u0_u3_u6_n142, u0_u3_u6_n143, 
       u0_u3_u6_n144, u0_u3_u6_n145, u0_u3_u6_n146, u0_u3_u6_n147, u0_u3_u6_n148, u0_u3_u6_n149, u0_u3_u6_n150, u0_u3_u6_n151, u0_u3_u6_n152, 
       u0_u3_u6_n153, u0_u3_u6_n154, u0_u3_u6_n155, u0_u3_u6_n156, u0_u3_u6_n157, u0_u3_u6_n158, u0_u3_u6_n159, u0_u3_u6_n160, u0_u3_u6_n161, 
       u0_u3_u6_n162, u0_u3_u6_n163, u0_u3_u6_n164, u0_u3_u6_n165, u0_u3_u6_n166, u0_u3_u6_n167, u0_u3_u6_n168, u0_u3_u6_n169, u0_u3_u6_n170, 
       u0_u3_u6_n171, u0_u3_u6_n172, u0_u3_u6_n173, u0_u3_u6_n174, u0_u3_u6_n88, u0_u3_u6_n89, u0_u3_u6_n90, u0_u3_u6_n91, u0_u3_u6_n92, 
       u0_u3_u6_n93, u0_u3_u6_n94, u0_u3_u6_n95, u0_u3_u6_n96, u0_u3_u6_n97, u0_u3_u6_n98, u0_u3_u6_n99, u0_u3_u7_n100, u0_u3_u7_n101, 
       u0_u3_u7_n102, u0_u3_u7_n103, u0_u3_u7_n104, u0_u3_u7_n105, u0_u3_u7_n106, u0_u3_u7_n107, u0_u3_u7_n108, u0_u3_u7_n109, u0_u3_u7_n110, 
       u0_u3_u7_n111, u0_u3_u7_n112, u0_u3_u7_n113, u0_u3_u7_n114, u0_u3_u7_n115, u0_u3_u7_n116, u0_u3_u7_n117, u0_u3_u7_n118, u0_u3_u7_n119, 
       u0_u3_u7_n120, u0_u3_u7_n121, u0_u3_u7_n122, u0_u3_u7_n123, u0_u3_u7_n124, u0_u3_u7_n125, u0_u3_u7_n126, u0_u3_u7_n127, u0_u3_u7_n128, 
       u0_u3_u7_n129, u0_u3_u7_n130, u0_u3_u7_n131, u0_u3_u7_n132, u0_u3_u7_n133, u0_u3_u7_n134, u0_u3_u7_n135, u0_u3_u7_n136, u0_u3_u7_n137, 
       u0_u3_u7_n138, u0_u3_u7_n139, u0_u3_u7_n140, u0_u3_u7_n141, u0_u3_u7_n142, u0_u3_u7_n143, u0_u3_u7_n144, u0_u3_u7_n145, u0_u3_u7_n146, 
       u0_u3_u7_n147, u0_u3_u7_n148, u0_u3_u7_n149, u0_u3_u7_n150, u0_u3_u7_n151, u0_u3_u7_n152, u0_u3_u7_n153, u0_u3_u7_n154, u0_u3_u7_n155, 
       u0_u3_u7_n156, u0_u3_u7_n157, u0_u3_u7_n158, u0_u3_u7_n159, u0_u3_u7_n160, u0_u3_u7_n161, u0_u3_u7_n162, u0_u3_u7_n163, u0_u3_u7_n164, 
       u0_u3_u7_n165, u0_u3_u7_n166, u0_u3_u7_n167, u0_u3_u7_n168, u0_u3_u7_n169, u0_u3_u7_n170, u0_u3_u7_n171, u0_u3_u7_n172, u0_u3_u7_n173, 
       u0_u3_u7_n174, u0_u3_u7_n175, u0_u3_u7_n176, u0_u3_u7_n177, u0_u3_u7_n178, u0_u3_u7_n179, u0_u3_u7_n180, u0_u3_u7_n91, u0_u3_u7_n92, 
       u0_u3_u7_n93, u0_u3_u7_n94, u0_u3_u7_n95, u0_u3_u7_n96, u0_u3_u7_n97, u0_u3_u7_n98, u0_u3_u7_n99, u0_u4_X_1, u0_u4_X_18, 
       u0_u4_X_20, u0_u4_X_22, u0_u4_X_24, u0_u4_X_26, u0_u4_X_27, u0_u4_X_29, u0_u4_X_31, u0_u4_X_33, u0_u4_X_35, 
       u0_u4_X_36, u0_u4_X_47, u0_u4_X_6, u0_u4_X_8, u0_u4_u0_n100, u0_u4_u0_n101, u0_u4_u0_n102, u0_u4_u0_n103, u0_u4_u0_n104, 
       u0_u4_u0_n105, u0_u4_u0_n106, u0_u4_u0_n107, u0_u4_u0_n108, u0_u4_u0_n109, u0_u4_u0_n110, u0_u4_u0_n111, u0_u4_u0_n112, u0_u4_u0_n113, 
       u0_u4_u0_n114, u0_u4_u0_n115, u0_u4_u0_n116, u0_u4_u0_n117, u0_u4_u0_n118, u0_u4_u0_n119, u0_u4_u0_n120, u0_u4_u0_n121, u0_u4_u0_n122, 
       u0_u4_u0_n123, u0_u4_u0_n124, u0_u4_u0_n125, u0_u4_u0_n126, u0_u4_u0_n127, u0_u4_u0_n128, u0_u4_u0_n129, u0_u4_u0_n130, u0_u4_u0_n131, 
       u0_u4_u0_n132, u0_u4_u0_n133, u0_u4_u0_n134, u0_u4_u0_n135, u0_u4_u0_n136, u0_u4_u0_n137, u0_u4_u0_n138, u0_u4_u0_n139, u0_u4_u0_n140, 
       u0_u4_u0_n141, u0_u4_u0_n142, u0_u4_u0_n143, u0_u4_u0_n144, u0_u4_u0_n145, u0_u4_u0_n146, u0_u4_u0_n147, u0_u4_u0_n148, u0_u4_u0_n149, 
       u0_u4_u0_n150, u0_u4_u0_n151, u0_u4_u0_n152, u0_u4_u0_n153, u0_u4_u0_n154, u0_u4_u0_n155, u0_u4_u0_n156, u0_u4_u0_n157, u0_u4_u0_n158, 
       u0_u4_u0_n159, u0_u4_u0_n160, u0_u4_u0_n161, u0_u4_u0_n162, u0_u4_u0_n163, u0_u4_u0_n164, u0_u4_u0_n165, u0_u4_u0_n166, u0_u4_u0_n167, 
       u0_u4_u0_n168, u0_u4_u0_n169, u0_u4_u0_n170, u0_u4_u0_n171, u0_u4_u0_n172, u0_u4_u0_n173, u0_u4_u0_n174, u0_u4_u0_n88, u0_u4_u0_n89, 
       u0_u4_u0_n90, u0_u4_u0_n91, u0_u4_u0_n92, u0_u4_u0_n93, u0_u4_u0_n94, u0_u4_u0_n95, u0_u4_u0_n96, u0_u4_u0_n97, u0_u4_u0_n98, 
       u0_u4_u0_n99, u0_u4_u1_n100, u0_u4_u1_n101, u0_u4_u1_n102, u0_u4_u1_n103, u0_u4_u1_n104, u0_u4_u1_n105, u0_u4_u1_n106, u0_u4_u1_n107, 
       u0_u4_u1_n108, u0_u4_u1_n109, u0_u4_u1_n110, u0_u4_u1_n111, u0_u4_u1_n112, u0_u4_u1_n113, u0_u4_u1_n114, u0_u4_u1_n115, u0_u4_u1_n116, 
       u0_u4_u1_n117, u0_u4_u1_n118, u0_u4_u1_n119, u0_u4_u1_n120, u0_u4_u1_n121, u0_u4_u1_n122, u0_u4_u1_n123, u0_u4_u1_n124, u0_u4_u1_n125, 
       u0_u4_u1_n126, u0_u4_u1_n127, u0_u4_u1_n128, u0_u4_u1_n129, u0_u4_u1_n130, u0_u4_u1_n131, u0_u4_u1_n132, u0_u4_u1_n133, u0_u4_u1_n134, 
       u0_u4_u1_n135, u0_u4_u1_n136, u0_u4_u1_n137, u0_u4_u1_n138, u0_u4_u1_n139, u0_u4_u1_n140, u0_u4_u1_n141, u0_u4_u1_n142, u0_u4_u1_n143, 
       u0_u4_u1_n144, u0_u4_u1_n145, u0_u4_u1_n146, u0_u4_u1_n147, u0_u4_u1_n148, u0_u4_u1_n149, u0_u4_u1_n150, u0_u4_u1_n151, u0_u4_u1_n152, 
       u0_u4_u1_n153, u0_u4_u1_n154, u0_u4_u1_n155, u0_u4_u1_n156, u0_u4_u1_n157, u0_u4_u1_n158, u0_u4_u1_n159, u0_u4_u1_n160, u0_u4_u1_n161, 
       u0_u4_u1_n162, u0_u4_u1_n163, u0_u4_u1_n164, u0_u4_u1_n165, u0_u4_u1_n166, u0_u4_u1_n167, u0_u4_u1_n168, u0_u4_u1_n169, u0_u4_u1_n170, 
       u0_u4_u1_n171, u0_u4_u1_n172, u0_u4_u1_n173, u0_u4_u1_n174, u0_u4_u1_n175, u0_u4_u1_n176, u0_u4_u1_n177, u0_u4_u1_n178, u0_u4_u1_n179, 
       u0_u4_u1_n180, u0_u4_u1_n181, u0_u4_u1_n182, u0_u4_u1_n183, u0_u4_u1_n184, u0_u4_u1_n185, u0_u4_u1_n186, u0_u4_u1_n187, u0_u4_u1_n188, 
       u0_u4_u1_n95, u0_u4_u1_n96, u0_u4_u1_n97, u0_u4_u1_n98, u0_u4_u1_n99, u0_u4_u2_n100, u0_u4_u2_n101, u0_u4_u2_n102, u0_u4_u2_n103, 
       u0_u4_u2_n104, u0_u4_u2_n105, u0_u4_u2_n106, u0_u4_u2_n107, u0_u4_u2_n108, u0_u4_u2_n109, u0_u4_u2_n110, u0_u4_u2_n111, u0_u4_u2_n112, 
       u0_u4_u2_n113, u0_u4_u2_n114, u0_u4_u2_n115, u0_u4_u2_n116, u0_u4_u2_n117, u0_u4_u2_n118, u0_u4_u2_n119, u0_u4_u2_n120, u0_u4_u2_n121, 
       u0_u4_u2_n122, u0_u4_u2_n123, u0_u4_u2_n124, u0_u4_u2_n125, u0_u4_u2_n126, u0_u4_u2_n127, u0_u4_u2_n128, u0_u4_u2_n129, u0_u4_u2_n130, 
       u0_u4_u2_n131, u0_u4_u2_n132, u0_u4_u2_n133, u0_u4_u2_n134, u0_u4_u2_n135, u0_u4_u2_n136, u0_u4_u2_n137, u0_u4_u2_n138, u0_u4_u2_n139, 
       u0_u4_u2_n140, u0_u4_u2_n141, u0_u4_u2_n142, u0_u4_u2_n143, u0_u4_u2_n144, u0_u4_u2_n145, u0_u4_u2_n146, u0_u4_u2_n147, u0_u4_u2_n148, 
       u0_u4_u2_n149, u0_u4_u2_n150, u0_u4_u2_n151, u0_u4_u2_n152, u0_u4_u2_n153, u0_u4_u2_n154, u0_u4_u2_n155, u0_u4_u2_n156, u0_u4_u2_n157, 
       u0_u4_u2_n158, u0_u4_u2_n159, u0_u4_u2_n160, u0_u4_u2_n161, u0_u4_u2_n162, u0_u4_u2_n163, u0_u4_u2_n164, u0_u4_u2_n165, u0_u4_u2_n166, 
       u0_u4_u2_n167, u0_u4_u2_n168, u0_u4_u2_n169, u0_u4_u2_n170, u0_u4_u2_n171, u0_u4_u2_n172, u0_u4_u2_n173, u0_u4_u2_n174, u0_u4_u2_n175, 
       u0_u4_u2_n176, u0_u4_u2_n177, u0_u4_u2_n178, u0_u4_u2_n179, u0_u4_u2_n180, u0_u4_u2_n181, u0_u4_u2_n182, u0_u4_u2_n183, u0_u4_u2_n184, 
       u0_u4_u2_n185, u0_u4_u2_n186, u0_u4_u2_n187, u0_u4_u2_n188, u0_u4_u2_n95, u0_u4_u2_n96, u0_u4_u2_n97, u0_u4_u2_n98, u0_u4_u2_n99, 
       u0_u4_u3_n100, u0_u4_u3_n101, u0_u4_u3_n102, u0_u4_u3_n103, u0_u4_u3_n104, u0_u4_u3_n105, u0_u4_u3_n106, u0_u4_u3_n107, u0_u4_u3_n108, 
       u0_u4_u3_n109, u0_u4_u3_n110, u0_u4_u3_n111, u0_u4_u3_n112, u0_u4_u3_n113, u0_u4_u3_n114, u0_u4_u3_n115, u0_u4_u3_n116, u0_u4_u3_n117, 
       u0_u4_u3_n118, u0_u4_u3_n119, u0_u4_u3_n120, u0_u4_u3_n121, u0_u4_u3_n122, u0_u4_u3_n123, u0_u4_u3_n124, u0_u4_u3_n125, u0_u4_u3_n126, 
       u0_u4_u3_n127, u0_u4_u3_n128, u0_u4_u3_n129, u0_u4_u3_n130, u0_u4_u3_n131, u0_u4_u3_n132, u0_u4_u3_n133, u0_u4_u3_n134, u0_u4_u3_n135, 
       u0_u4_u3_n136, u0_u4_u3_n137, u0_u4_u3_n138, u0_u4_u3_n139, u0_u4_u3_n140, u0_u4_u3_n141, u0_u4_u3_n142, u0_u4_u3_n143, u0_u4_u3_n144, 
       u0_u4_u3_n145, u0_u4_u3_n146, u0_u4_u3_n147, u0_u4_u3_n148, u0_u4_u3_n149, u0_u4_u3_n150, u0_u4_u3_n151, u0_u4_u3_n152, u0_u4_u3_n153, 
       u0_u4_u3_n154, u0_u4_u3_n155, u0_u4_u3_n156, u0_u4_u3_n157, u0_u4_u3_n158, u0_u4_u3_n159, u0_u4_u3_n160, u0_u4_u3_n161, u0_u4_u3_n162, 
       u0_u4_u3_n163, u0_u4_u3_n164, u0_u4_u3_n165, u0_u4_u3_n166, u0_u4_u3_n167, u0_u4_u3_n168, u0_u4_u3_n169, u0_u4_u3_n170, u0_u4_u3_n171, 
       u0_u4_u3_n172, u0_u4_u3_n173, u0_u4_u3_n174, u0_u4_u3_n175, u0_u4_u3_n176, u0_u4_u3_n177, u0_u4_u3_n178, u0_u4_u3_n179, u0_u4_u3_n180, 
       u0_u4_u3_n181, u0_u4_u3_n182, u0_u4_u3_n183, u0_u4_u3_n184, u0_u4_u3_n185, u0_u4_u3_n186, u0_u4_u3_n94, u0_u4_u3_n95, u0_u4_u3_n96, 
       u0_u4_u3_n97, u0_u4_u3_n98, u0_u4_u3_n99, u0_u4_u4_n100, u0_u4_u4_n101, u0_u4_u4_n102, u0_u4_u4_n103, u0_u4_u4_n104, u0_u4_u4_n105, 
       u0_u4_u4_n106, u0_u4_u4_n107, u0_u4_u4_n108, u0_u4_u4_n109, u0_u4_u4_n110, u0_u4_u4_n111, u0_u4_u4_n112, u0_u4_u4_n113, u0_u4_u4_n114, 
       u0_u4_u4_n115, u0_u4_u4_n116, u0_u4_u4_n117, u0_u4_u4_n118, u0_u4_u4_n119, u0_u4_u4_n120, u0_u4_u4_n121, u0_u4_u4_n122, u0_u4_u4_n123, 
       u0_u4_u4_n124, u0_u4_u4_n125, u0_u4_u4_n126, u0_u4_u4_n127, u0_u4_u4_n128, u0_u4_u4_n129, u0_u4_u4_n130, u0_u4_u4_n131, u0_u4_u4_n132, 
       u0_u4_u4_n133, u0_u4_u4_n134, u0_u4_u4_n135, u0_u4_u4_n136, u0_u4_u4_n137, u0_u4_u4_n138, u0_u4_u4_n139, u0_u4_u4_n140, u0_u4_u4_n141, 
       u0_u4_u4_n142, u0_u4_u4_n143, u0_u4_u4_n144, u0_u4_u4_n145, u0_u4_u4_n146, u0_u4_u4_n147, u0_u4_u4_n148, u0_u4_u4_n149, u0_u4_u4_n150, 
       u0_u4_u4_n151, u0_u4_u4_n152, u0_u4_u4_n153, u0_u4_u4_n154, u0_u4_u4_n155, u0_u4_u4_n156, u0_u4_u4_n157, u0_u4_u4_n158, u0_u4_u4_n159, 
       u0_u4_u4_n160, u0_u4_u4_n161, u0_u4_u4_n162, u0_u4_u4_n163, u0_u4_u4_n164, u0_u4_u4_n165, u0_u4_u4_n166, u0_u4_u4_n167, u0_u4_u4_n168, 
       u0_u4_u4_n169, u0_u4_u4_n170, u0_u4_u4_n171, u0_u4_u4_n172, u0_u4_u4_n173, u0_u4_u4_n174, u0_u4_u4_n175, u0_u4_u4_n176, u0_u4_u4_n177, 
       u0_u4_u4_n178, u0_u4_u4_n179, u0_u4_u4_n180, u0_u4_u4_n181, u0_u4_u4_n182, u0_u4_u4_n183, u0_u4_u4_n184, u0_u4_u4_n185, u0_u4_u4_n186, 
       u0_u4_u4_n94, u0_u4_u4_n95, u0_u4_u4_n96, u0_u4_u4_n97, u0_u4_u4_n98, u0_u4_u4_n99, u0_u4_u5_n100, u0_u4_u5_n101, u0_u4_u5_n102, 
       u0_u4_u5_n103, u0_u4_u5_n104, u0_u4_u5_n105, u0_u4_u5_n106, u0_u4_u5_n107, u0_u4_u5_n108, u0_u4_u5_n109, u0_u4_u5_n110, u0_u4_u5_n111, 
       u0_u4_u5_n112, u0_u4_u5_n113, u0_u4_u5_n114, u0_u4_u5_n115, u0_u4_u5_n116, u0_u4_u5_n117, u0_u4_u5_n118, u0_u4_u5_n119, u0_u4_u5_n120, 
       u0_u4_u5_n121, u0_u4_u5_n122, u0_u4_u5_n123, u0_u4_u5_n124, u0_u4_u5_n125, u0_u4_u5_n126, u0_u4_u5_n127, u0_u4_u5_n128, u0_u4_u5_n129, 
       u0_u4_u5_n130, u0_u4_u5_n131, u0_u4_u5_n132, u0_u4_u5_n133, u0_u4_u5_n134, u0_u4_u5_n135, u0_u4_u5_n136, u0_u4_u5_n137, u0_u4_u5_n138, 
       u0_u4_u5_n139, u0_u4_u5_n140, u0_u4_u5_n141, u0_u4_u5_n142, u0_u4_u5_n143, u0_u4_u5_n144, u0_u4_u5_n145, u0_u4_u5_n146, u0_u4_u5_n147, 
       u0_u4_u5_n148, u0_u4_u5_n149, u0_u4_u5_n150, u0_u4_u5_n151, u0_u4_u5_n152, u0_u4_u5_n153, u0_u4_u5_n154, u0_u4_u5_n155, u0_u4_u5_n156, 
       u0_u4_u5_n157, u0_u4_u5_n158, u0_u4_u5_n159, u0_u4_u5_n160, u0_u4_u5_n161, u0_u4_u5_n162, u0_u4_u5_n163, u0_u4_u5_n164, u0_u4_u5_n165, 
       u0_u4_u5_n166, u0_u4_u5_n167, u0_u4_u5_n168, u0_u4_u5_n169, u0_u4_u5_n170, u0_u4_u5_n171, u0_u4_u5_n172, u0_u4_u5_n173, u0_u4_u5_n174, 
       u0_u4_u5_n175, u0_u4_u5_n176, u0_u4_u5_n177, u0_u4_u5_n178, u0_u4_u5_n179, u0_u4_u5_n180, u0_u4_u5_n181, u0_u4_u5_n182, u0_u4_u5_n183, 
       u0_u4_u5_n184, u0_u4_u5_n185, u0_u4_u5_n186, u0_u4_u5_n187, u0_u4_u5_n188, u0_u4_u5_n189, u0_u4_u5_n190, u0_u4_u5_n191, u0_u4_u5_n192, 
       u0_u4_u5_n193, u0_u4_u5_n194, u0_u4_u5_n195, u0_u4_u5_n196, u0_u4_u5_n99, u0_u4_u7_n100, u0_u4_u7_n101, u0_u4_u7_n102, u0_u4_u7_n103, 
       u0_u4_u7_n104, u0_u4_u7_n105, u0_u4_u7_n106, u0_u4_u7_n107, u0_u4_u7_n108, u0_u4_u7_n109, u0_u4_u7_n110, u0_u4_u7_n111, u0_u4_u7_n112, 
       u0_u4_u7_n113, u0_u4_u7_n114, u0_u4_u7_n115, u0_u4_u7_n116, u0_u4_u7_n117, u0_u4_u7_n118, u0_u4_u7_n119, u0_u4_u7_n120, u0_u4_u7_n121, 
       u0_u4_u7_n122, u0_u4_u7_n123, u0_u4_u7_n124, u0_u4_u7_n125, u0_u4_u7_n126, u0_u4_u7_n127, u0_u4_u7_n128, u0_u4_u7_n129, u0_u4_u7_n130, 
       u0_u4_u7_n131, u0_u4_u7_n132, u0_u4_u7_n133, u0_u4_u7_n134, u0_u4_u7_n135, u0_u4_u7_n136, u0_u4_u7_n137, u0_u4_u7_n138, u0_u4_u7_n139, 
       u0_u4_u7_n140, u0_u4_u7_n141, u0_u4_u7_n142, u0_u4_u7_n143, u0_u4_u7_n144, u0_u4_u7_n145, u0_u4_u7_n146, u0_u4_u7_n147, u0_u4_u7_n148, 
       u0_u4_u7_n149, u0_u4_u7_n150, u0_u4_u7_n151, u0_u4_u7_n152, u0_u4_u7_n153, u0_u4_u7_n154, u0_u4_u7_n155, u0_u4_u7_n156, u0_u4_u7_n157, 
       u0_u4_u7_n158, u0_u4_u7_n159, u0_u4_u7_n160, u0_u4_u7_n161, u0_u4_u7_n162, u0_u4_u7_n163, u0_u4_u7_n164, u0_u4_u7_n165, u0_u4_u7_n166, 
       u0_u4_u7_n167, u0_u4_u7_n168, u0_u4_u7_n169, u0_u4_u7_n170, u0_u4_u7_n171, u0_u4_u7_n172, u0_u4_u7_n173, u0_u4_u7_n174, u0_u4_u7_n175, 
       u0_u4_u7_n176, u0_u4_u7_n177, u0_u4_u7_n178, u0_u4_u7_n179, u0_u4_u7_n180, u0_u4_u7_n91, u0_u4_u7_n92, u0_u4_u7_n93, u0_u4_u7_n94, 
       u0_u4_u7_n95, u0_u4_u7_n96, u0_u4_u7_n97, u0_u4_u7_n98, u0_u4_u7_n99, u0_u6_X_1, u0_u6_X_10, u0_u6_X_11, u0_u6_X_12, 
       u0_u6_X_13, u0_u6_X_14, u0_u6_X_17, u0_u6_X_18, u0_u6_X_19, u0_u6_X_20, u0_u6_X_3, u0_u6_X_36, u0_u6_X_4, 
       u0_u6_X_5, u0_u6_X_6, u0_u6_X_7, u0_u6_X_8, u0_u6_u0_n100, u0_u6_u0_n101, u0_u6_u0_n102, u0_u6_u0_n103, u0_u6_u0_n104, 
       u0_u6_u0_n105, u0_u6_u0_n106, u0_u6_u0_n107, u0_u6_u0_n108, u0_u6_u0_n109, u0_u6_u0_n110, u0_u6_u0_n111, u0_u6_u0_n112, u0_u6_u0_n113, 
       u0_u6_u0_n114, u0_u6_u0_n115, u0_u6_u0_n116, u0_u6_u0_n117, u0_u6_u0_n118, u0_u6_u0_n119, u0_u6_u0_n120, u0_u6_u0_n121, u0_u6_u0_n122, 
       u0_u6_u0_n123, u0_u6_u0_n124, u0_u6_u0_n125, u0_u6_u0_n126, u0_u6_u0_n127, u0_u6_u0_n128, u0_u6_u0_n129, u0_u6_u0_n130, u0_u6_u0_n131, 
       u0_u6_u0_n132, u0_u6_u0_n133, u0_u6_u0_n134, u0_u6_u0_n135, u0_u6_u0_n136, u0_u6_u0_n137, u0_u6_u0_n138, u0_u6_u0_n139, u0_u6_u0_n140, 
       u0_u6_u0_n141, u0_u6_u0_n142, u0_u6_u0_n143, u0_u6_u0_n144, u0_u6_u0_n145, u0_u6_u0_n146, u0_u6_u0_n147, u0_u6_u0_n148, u0_u6_u0_n149, 
       u0_u6_u0_n150, u0_u6_u0_n151, u0_u6_u0_n152, u0_u6_u0_n153, u0_u6_u0_n154, u0_u6_u0_n155, u0_u6_u0_n156, u0_u6_u0_n157, u0_u6_u0_n158, 
       u0_u6_u0_n159, u0_u6_u0_n160, u0_u6_u0_n161, u0_u6_u0_n162, u0_u6_u0_n163, u0_u6_u0_n164, u0_u6_u0_n165, u0_u6_u0_n166, u0_u6_u0_n167, 
       u0_u6_u0_n168, u0_u6_u0_n169, u0_u6_u0_n170, u0_u6_u0_n171, u0_u6_u0_n172, u0_u6_u0_n173, u0_u6_u0_n174, u0_u6_u0_n88, u0_u6_u0_n89, 
       u0_u6_u0_n90, u0_u6_u0_n91, u0_u6_u0_n92, u0_u6_u0_n93, u0_u6_u0_n94, u0_u6_u0_n95, u0_u6_u0_n96, u0_u6_u0_n97, u0_u6_u0_n98, 
       u0_u6_u0_n99, u0_u6_u1_n100, u0_u6_u1_n101, u0_u6_u1_n102, u0_u6_u1_n103, u0_u6_u1_n104, u0_u6_u1_n105, u0_u6_u1_n106, u0_u6_u1_n107, 
       u0_u6_u1_n108, u0_u6_u1_n109, u0_u6_u1_n110, u0_u6_u1_n111, u0_u6_u1_n112, u0_u6_u1_n113, u0_u6_u1_n114, u0_u6_u1_n115, u0_u6_u1_n116, 
       u0_u6_u1_n117, u0_u6_u1_n118, u0_u6_u1_n119, u0_u6_u1_n120, u0_u6_u1_n121, u0_u6_u1_n122, u0_u6_u1_n123, u0_u6_u1_n124, u0_u6_u1_n125, 
       u0_u6_u1_n126, u0_u6_u1_n127, u0_u6_u1_n128, u0_u6_u1_n129, u0_u6_u1_n130, u0_u6_u1_n131, u0_u6_u1_n132, u0_u6_u1_n133, u0_u6_u1_n134, 
       u0_u6_u1_n135, u0_u6_u1_n136, u0_u6_u1_n137, u0_u6_u1_n138, u0_u6_u1_n139, u0_u6_u1_n140, u0_u6_u1_n141, u0_u6_u1_n142, u0_u6_u1_n143, 
       u0_u6_u1_n144, u0_u6_u1_n145, u0_u6_u1_n146, u0_u6_u1_n147, u0_u6_u1_n148, u0_u6_u1_n149, u0_u6_u1_n150, u0_u6_u1_n151, u0_u6_u1_n152, 
       u0_u6_u1_n153, u0_u6_u1_n154, u0_u6_u1_n155, u0_u6_u1_n156, u0_u6_u1_n157, u0_u6_u1_n158, u0_u6_u1_n159, u0_u6_u1_n160, u0_u6_u1_n161, 
       u0_u6_u1_n162, u0_u6_u1_n163, u0_u6_u1_n164, u0_u6_u1_n165, u0_u6_u1_n166, u0_u6_u1_n167, u0_u6_u1_n168, u0_u6_u1_n169, u0_u6_u1_n170, 
       u0_u6_u1_n171, u0_u6_u1_n172, u0_u6_u1_n173, u0_u6_u1_n174, u0_u6_u1_n175, u0_u6_u1_n176, u0_u6_u1_n177, u0_u6_u1_n178, u0_u6_u1_n179, 
       u0_u6_u1_n180, u0_u6_u1_n181, u0_u6_u1_n182, u0_u6_u1_n183, u0_u6_u1_n184, u0_u6_u1_n185, u0_u6_u1_n186, u0_u6_u1_n187, u0_u6_u1_n188, 
       u0_u6_u1_n95, u0_u6_u1_n96, u0_u6_u1_n97, u0_u6_u1_n98, u0_u6_u1_n99, u0_u6_u2_n100, u0_u6_u2_n101, u0_u6_u2_n102, u0_u6_u2_n103, 
       u0_u6_u2_n104, u0_u6_u2_n105, u0_u6_u2_n106, u0_u6_u2_n107, u0_u6_u2_n108, u0_u6_u2_n109, u0_u6_u2_n110, u0_u6_u2_n111, u0_u6_u2_n112, 
       u0_u6_u2_n113, u0_u6_u2_n114, u0_u6_u2_n115, u0_u6_u2_n116, u0_u6_u2_n117, u0_u6_u2_n118, u0_u6_u2_n119, u0_u6_u2_n120, u0_u6_u2_n121, 
       u0_u6_u2_n122, u0_u6_u2_n123, u0_u6_u2_n124, u0_u6_u2_n125, u0_u6_u2_n126, u0_u6_u2_n127, u0_u6_u2_n128, u0_u6_u2_n129, u0_u6_u2_n130, 
       u0_u6_u2_n131, u0_u6_u2_n132, u0_u6_u2_n133, u0_u6_u2_n134, u0_u6_u2_n135, u0_u6_u2_n136, u0_u6_u2_n137, u0_u6_u2_n138, u0_u6_u2_n139, 
       u0_u6_u2_n140, u0_u6_u2_n141, u0_u6_u2_n142, u0_u6_u2_n143, u0_u6_u2_n144, u0_u6_u2_n145, u0_u6_u2_n146, u0_u6_u2_n147, u0_u6_u2_n148, 
       u0_u6_u2_n149, u0_u6_u2_n150, u0_u6_u2_n151, u0_u6_u2_n152, u0_u6_u2_n153, u0_u6_u2_n154, u0_u6_u2_n155, u0_u6_u2_n156, u0_u6_u2_n157, 
       u0_u6_u2_n158, u0_u6_u2_n159, u0_u6_u2_n160, u0_u6_u2_n161, u0_u6_u2_n162, u0_u6_u2_n163, u0_u6_u2_n164, u0_u6_u2_n165, u0_u6_u2_n166, 
       u0_u6_u2_n167, u0_u6_u2_n168, u0_u6_u2_n169, u0_u6_u2_n170, u0_u6_u2_n171, u0_u6_u2_n172, u0_u6_u2_n173, u0_u6_u2_n174, u0_u6_u2_n175, 
       u0_u6_u2_n176, u0_u6_u2_n177, u0_u6_u2_n178, u0_u6_u2_n179, u0_u6_u2_n180, u0_u6_u2_n181, u0_u6_u2_n182, u0_u6_u2_n183, u0_u6_u2_n184, 
       u0_u6_u2_n185, u0_u6_u2_n186, u0_u6_u2_n187, u0_u6_u2_n188, u0_u6_u2_n95, u0_u6_u2_n96, u0_u6_u2_n97, u0_u6_u2_n98, u0_u6_u2_n99, 
       u0_u6_u3_n100, u0_u6_u3_n101, u0_u6_u3_n102, u0_u6_u3_n103, u0_u6_u3_n104, u0_u6_u3_n105, u0_u6_u3_n106, u0_u6_u3_n107, u0_u6_u3_n108, 
       u0_u6_u3_n109, u0_u6_u3_n110, u0_u6_u3_n111, u0_u6_u3_n112, u0_u6_u3_n113, u0_u6_u3_n114, u0_u6_u3_n115, u0_u6_u3_n116, u0_u6_u3_n117, 
       u0_u6_u3_n118, u0_u6_u3_n119, u0_u6_u3_n120, u0_u6_u3_n121, u0_u6_u3_n122, u0_u6_u3_n123, u0_u6_u3_n124, u0_u6_u3_n125, u0_u6_u3_n126, 
       u0_u6_u3_n127, u0_u6_u3_n128, u0_u6_u3_n129, u0_u6_u3_n130, u0_u6_u3_n131, u0_u6_u3_n132, u0_u6_u3_n133, u0_u6_u3_n134, u0_u6_u3_n135, 
       u0_u6_u3_n136, u0_u6_u3_n137, u0_u6_u3_n138, u0_u6_u3_n139, u0_u6_u3_n140, u0_u6_u3_n141, u0_u6_u3_n142, u0_u6_u3_n143, u0_u6_u3_n144, 
       u0_u6_u3_n145, u0_u6_u3_n146, u0_u6_u3_n147, u0_u6_u3_n148, u0_u6_u3_n149, u0_u6_u3_n150, u0_u6_u3_n151, u0_u6_u3_n152, u0_u6_u3_n153, 
       u0_u6_u3_n154, u0_u6_u3_n155, u0_u6_u3_n156, u0_u6_u3_n157, u0_u6_u3_n158, u0_u6_u3_n159, u0_u6_u3_n160, u0_u6_u3_n161, u0_u6_u3_n162, 
       u0_u6_u3_n163, u0_u6_u3_n164, u0_u6_u3_n165, u0_u6_u3_n166, u0_u6_u3_n167, u0_u6_u3_n168, u0_u6_u3_n169, u0_u6_u3_n170, u0_u6_u3_n171, 
       u0_u6_u3_n172, u0_u6_u3_n173, u0_u6_u3_n174, u0_u6_u3_n175, u0_u6_u3_n176, u0_u6_u3_n177, u0_u6_u3_n178, u0_u6_u3_n179, u0_u6_u3_n180, 
       u0_u6_u3_n181, u0_u6_u3_n182, u0_u6_u3_n183, u0_u6_u3_n184, u0_u6_u3_n185, u0_u6_u3_n186, u0_u6_u3_n94, u0_u6_u3_n95, u0_u6_u3_n96, 
       u0_u6_u3_n97, u0_u6_u3_n98, u0_u6_u3_n99, u0_u6_u5_n100, u0_u6_u5_n101, u0_u6_u5_n102, u0_u6_u5_n103, u0_u6_u5_n104, u0_u6_u5_n105, 
       u0_u6_u5_n106, u0_u6_u5_n107, u0_u6_u5_n108, u0_u6_u5_n109, u0_u6_u5_n110, u0_u6_u5_n111, u0_u6_u5_n112, u0_u6_u5_n113, u0_u6_u5_n114, 
       u0_u6_u5_n115, u0_u6_u5_n116, u0_u6_u5_n117, u0_u6_u5_n118, u0_u6_u5_n119, u0_u6_u5_n120, u0_u6_u5_n121, u0_u6_u5_n122, u0_u6_u5_n123, 
       u0_u6_u5_n124, u0_u6_u5_n125, u0_u6_u5_n126, u0_u6_u5_n127, u0_u6_u5_n128, u0_u6_u5_n129, u0_u6_u5_n130, u0_u6_u5_n131, u0_u6_u5_n132, 
       u0_u6_u5_n133, u0_u6_u5_n134, u0_u6_u5_n135, u0_u6_u5_n136, u0_u6_u5_n137, u0_u6_u5_n138, u0_u6_u5_n139, u0_u6_u5_n140, u0_u6_u5_n141, 
       u0_u6_u5_n142, u0_u6_u5_n143, u0_u6_u5_n144, u0_u6_u5_n145, u0_u6_u5_n146, u0_u6_u5_n147, u0_u6_u5_n148, u0_u6_u5_n149, u0_u6_u5_n150, 
       u0_u6_u5_n151, u0_u6_u5_n152, u0_u6_u5_n153, u0_u6_u5_n154, u0_u6_u5_n155, u0_u6_u5_n156, u0_u6_u5_n157, u0_u6_u5_n158, u0_u6_u5_n159, 
       u0_u6_u5_n160, u0_u6_u5_n161, u0_u6_u5_n162, u0_u6_u5_n163, u0_u6_u5_n164, u0_u6_u5_n165, u0_u6_u5_n166, u0_u6_u5_n167, u0_u6_u5_n168, 
       u0_u6_u5_n169, u0_u6_u5_n170, u0_u6_u5_n171, u0_u6_u5_n172, u0_u6_u5_n173, u0_u6_u5_n174, u0_u6_u5_n175, u0_u6_u5_n176, u0_u6_u5_n177, 
       u0_u6_u5_n178, u0_u6_u5_n179, u0_u6_u5_n180, u0_u6_u5_n181, u0_u6_u5_n182, u0_u6_u5_n183, u0_u6_u5_n184, u0_u6_u5_n185, u0_u6_u5_n186, 
       u0_u6_u5_n187, u0_u6_u5_n188, u0_u6_u5_n189, u0_u6_u5_n190, u0_u6_u5_n191, u0_u6_u5_n192, u0_u6_u5_n193, u0_u6_u5_n194, u0_u6_u5_n195, 
       u0_u6_u5_n196, u0_u6_u5_n99, u0_u7_X_10, u0_u7_X_11, u0_u7_X_12, u0_u7_X_13, u0_u7_X_14, u0_u7_X_15, u0_u7_X_16, 
       u0_u7_X_17, u0_u7_X_18, u0_u7_X_19, u0_u7_X_20, u0_u7_X_21, u0_u7_X_24, u0_u7_X_5, u0_u7_X_6, u0_u7_X_7, 
       u0_u7_X_8, u0_u7_u0_n100, u0_u7_u0_n101, u0_u7_u0_n102, u0_u7_u0_n103, u0_u7_u0_n104, u0_u7_u0_n105, u0_u7_u0_n106, u0_u7_u0_n107, 
       u0_u7_u0_n108, u0_u7_u0_n109, u0_u7_u0_n110, u0_u7_u0_n111, u0_u7_u0_n112, u0_u7_u0_n113, u0_u7_u0_n114, u0_u7_u0_n115, u0_u7_u0_n116, 
       u0_u7_u0_n117, u0_u7_u0_n118, u0_u7_u0_n119, u0_u7_u0_n120, u0_u7_u0_n121, u0_u7_u0_n122, u0_u7_u0_n123, u0_u7_u0_n124, u0_u7_u0_n125, 
       u0_u7_u0_n126, u0_u7_u0_n127, u0_u7_u0_n128, u0_u7_u0_n129, u0_u7_u0_n130, u0_u7_u0_n131, u0_u7_u0_n132, u0_u7_u0_n133, u0_u7_u0_n134, 
       u0_u7_u0_n135, u0_u7_u0_n136, u0_u7_u0_n137, u0_u7_u0_n138, u0_u7_u0_n139, u0_u7_u0_n140, u0_u7_u0_n141, u0_u7_u0_n142, u0_u7_u0_n143, 
       u0_u7_u0_n144, u0_u7_u0_n145, u0_u7_u0_n146, u0_u7_u0_n147, u0_u7_u0_n148, u0_u7_u0_n149, u0_u7_u0_n150, u0_u7_u0_n151, u0_u7_u0_n152, 
       u0_u7_u0_n153, u0_u7_u0_n154, u0_u7_u0_n155, u0_u7_u0_n156, u0_u7_u0_n157, u0_u7_u0_n158, u0_u7_u0_n159, u0_u7_u0_n160, u0_u7_u0_n161, 
       u0_u7_u0_n162, u0_u7_u0_n163, u0_u7_u0_n164, u0_u7_u0_n165, u0_u7_u0_n166, u0_u7_u0_n167, u0_u7_u0_n168, u0_u7_u0_n169, u0_u7_u0_n170, 
       u0_u7_u0_n171, u0_u7_u0_n172, u0_u7_u0_n173, u0_u7_u0_n174, u0_u7_u0_n88, u0_u7_u0_n89, u0_u7_u0_n90, u0_u7_u0_n91, u0_u7_u0_n92, 
       u0_u7_u0_n93, u0_u7_u0_n94, u0_u7_u0_n95, u0_u7_u0_n96, u0_u7_u0_n97, u0_u7_u0_n98, u0_u7_u0_n99, u0_u7_u1_n100, u0_u7_u1_n101, 
       u0_u7_u1_n102, u0_u7_u1_n103, u0_u7_u1_n104, u0_u7_u1_n105, u0_u7_u1_n106, u0_u7_u1_n107, u0_u7_u1_n108, u0_u7_u1_n109, u0_u7_u1_n110, 
       u0_u7_u1_n111, u0_u7_u1_n112, u0_u7_u1_n113, u0_u7_u1_n114, u0_u7_u1_n115, u0_u7_u1_n116, u0_u7_u1_n117, u0_u7_u1_n118, u0_u7_u1_n119, 
       u0_u7_u1_n120, u0_u7_u1_n121, u0_u7_u1_n122, u0_u7_u1_n123, u0_u7_u1_n124, u0_u7_u1_n125, u0_u7_u1_n126, u0_u7_u1_n127, u0_u7_u1_n128, 
       u0_u7_u1_n129, u0_u7_u1_n130, u0_u7_u1_n131, u0_u7_u1_n132, u0_u7_u1_n133, u0_u7_u1_n134, u0_u7_u1_n135, u0_u7_u1_n136, u0_u7_u1_n137, 
       u0_u7_u1_n138, u0_u7_u1_n139, u0_u7_u1_n140, u0_u7_u1_n141, u0_u7_u1_n142, u0_u7_u1_n143, u0_u7_u1_n144, u0_u7_u1_n145, u0_u7_u1_n146, 
       u0_u7_u1_n147, u0_u7_u1_n148, u0_u7_u1_n149, u0_u7_u1_n150, u0_u7_u1_n151, u0_u7_u1_n152, u0_u7_u1_n153, u0_u7_u1_n154, u0_u7_u1_n155, 
       u0_u7_u1_n156, u0_u7_u1_n157, u0_u7_u1_n158, u0_u7_u1_n159, u0_u7_u1_n160, u0_u7_u1_n161, u0_u7_u1_n162, u0_u7_u1_n163, u0_u7_u1_n164, 
       u0_u7_u1_n165, u0_u7_u1_n166, u0_u7_u1_n167, u0_u7_u1_n168, u0_u7_u1_n169, u0_u7_u1_n170, u0_u7_u1_n171, u0_u7_u1_n172, u0_u7_u1_n173, 
       u0_u7_u1_n174, u0_u7_u1_n175, u0_u7_u1_n176, u0_u7_u1_n177, u0_u7_u1_n178, u0_u7_u1_n179, u0_u7_u1_n180, u0_u7_u1_n181, u0_u7_u1_n182, 
       u0_u7_u1_n183, u0_u7_u1_n184, u0_u7_u1_n185, u0_u7_u1_n186, u0_u7_u1_n187, u0_u7_u1_n188, u0_u7_u1_n95, u0_u7_u1_n96, u0_u7_u1_n97, 
       u0_u7_u1_n98, u0_u7_u1_n99, u0_u7_u2_n100, u0_u7_u2_n101, u0_u7_u2_n102, u0_u7_u2_n103, u0_u7_u2_n104, u0_u7_u2_n105, u0_u7_u2_n106, 
       u0_u7_u2_n107, u0_u7_u2_n108, u0_u7_u2_n109, u0_u7_u2_n110, u0_u7_u2_n111, u0_u7_u2_n112, u0_u7_u2_n113, u0_u7_u2_n114, u0_u7_u2_n115, 
       u0_u7_u2_n116, u0_u7_u2_n117, u0_u7_u2_n118, u0_u7_u2_n119, u0_u7_u2_n120, u0_u7_u2_n121, u0_u7_u2_n122, u0_u7_u2_n123, u0_u7_u2_n124, 
       u0_u7_u2_n125, u0_u7_u2_n126, u0_u7_u2_n127, u0_u7_u2_n128, u0_u7_u2_n129, u0_u7_u2_n130, u0_u7_u2_n131, u0_u7_u2_n132, u0_u7_u2_n133, 
       u0_u7_u2_n134, u0_u7_u2_n135, u0_u7_u2_n136, u0_u7_u2_n137, u0_u7_u2_n138, u0_u7_u2_n139, u0_u7_u2_n140, u0_u7_u2_n141, u0_u7_u2_n142, 
       u0_u7_u2_n143, u0_u7_u2_n144, u0_u7_u2_n145, u0_u7_u2_n146, u0_u7_u2_n147, u0_u7_u2_n148, u0_u7_u2_n149, u0_u7_u2_n150, u0_u7_u2_n151, 
       u0_u7_u2_n152, u0_u7_u2_n153, u0_u7_u2_n154, u0_u7_u2_n155, u0_u7_u2_n156, u0_u7_u2_n157, u0_u7_u2_n158, u0_u7_u2_n159, u0_u7_u2_n160, 
       u0_u7_u2_n161, u0_u7_u2_n162, u0_u7_u2_n163, u0_u7_u2_n164, u0_u7_u2_n165, u0_u7_u2_n166, u0_u7_u2_n167, u0_u7_u2_n168, u0_u7_u2_n169, 
       u0_u7_u2_n170, u0_u7_u2_n171, u0_u7_u2_n172, u0_u7_u2_n173, u0_u7_u2_n174, u0_u7_u2_n175, u0_u7_u2_n176, u0_u7_u2_n177, u0_u7_u2_n178, 
       u0_u7_u2_n179, u0_u7_u2_n180, u0_u7_u2_n181, u0_u7_u2_n182, u0_u7_u2_n183, u0_u7_u2_n184, u0_u7_u2_n185, u0_u7_u2_n186, u0_u7_u2_n187, 
       u0_u7_u2_n188, u0_u7_u2_n95, u0_u7_u2_n96, u0_u7_u2_n97, u0_u7_u2_n98, u0_u7_u2_n99, u0_u7_u3_n100, u0_u7_u3_n101, u0_u7_u3_n102, 
       u0_u7_u3_n103, u0_u7_u3_n104, u0_u7_u3_n105, u0_u7_u3_n106, u0_u7_u3_n107, u0_u7_u3_n108, u0_u7_u3_n109, u0_u7_u3_n110, u0_u7_u3_n111, 
       u0_u7_u3_n112, u0_u7_u3_n113, u0_u7_u3_n114, u0_u7_u3_n115, u0_u7_u3_n116, u0_u7_u3_n117, u0_u7_u3_n118, u0_u7_u3_n119, u0_u7_u3_n120, 
       u0_u7_u3_n121, u0_u7_u3_n122, u0_u7_u3_n123, u0_u7_u3_n124, u0_u7_u3_n125, u0_u7_u3_n126, u0_u7_u3_n127, u0_u7_u3_n128, u0_u7_u3_n129, 
       u0_u7_u3_n130, u0_u7_u3_n131, u0_u7_u3_n132, u0_u7_u3_n133, u0_u7_u3_n134, u0_u7_u3_n135, u0_u7_u3_n136, u0_u7_u3_n137, u0_u7_u3_n138, 
       u0_u7_u3_n139, u0_u7_u3_n140, u0_u7_u3_n141, u0_u7_u3_n142, u0_u7_u3_n143, u0_u7_u3_n144, u0_u7_u3_n145, u0_u7_u3_n146, u0_u7_u3_n147, 
       u0_u7_u3_n148, u0_u7_u3_n149, u0_u7_u3_n150, u0_u7_u3_n151, u0_u7_u3_n152, u0_u7_u3_n153, u0_u7_u3_n154, u0_u7_u3_n155, u0_u7_u3_n156, 
       u0_u7_u3_n157, u0_u7_u3_n158, u0_u7_u3_n159, u0_u7_u3_n160, u0_u7_u3_n161, u0_u7_u3_n162, u0_u7_u3_n163, u0_u7_u3_n164, u0_u7_u3_n165, 
       u0_u7_u3_n166, u0_u7_u3_n167, u0_u7_u3_n168, u0_u7_u3_n169, u0_u7_u3_n170, u0_u7_u3_n171, u0_u7_u3_n172, u0_u7_u3_n173, u0_u7_u3_n174, 
       u0_u7_u3_n175, u0_u7_u3_n176, u0_u7_u3_n177, u0_u7_u3_n178, u0_u7_u3_n179, u0_u7_u3_n180, u0_u7_u3_n181, u0_u7_u3_n182, u0_u7_u3_n183, 
       u0_u7_u3_n184, u0_u7_u3_n185, u0_u7_u3_n186, u0_u7_u3_n94, u0_u7_u3_n95, u0_u7_u3_n96, u0_u7_u3_n97, u0_u7_u3_n98, u0_u7_u3_n99, 
       u0_u9_X_1, u0_u9_X_12, u0_u9_X_14, u0_u9_X_17, u0_u9_X_18, u0_u9_X_19, u0_u9_X_2, u0_u9_X_20, u0_u9_X_24, 
       u0_u9_X_26, u0_u9_X_28, u0_u9_X_29, u0_u9_X_30, u0_u9_X_31, u0_u9_X_32, u0_u9_X_33, u0_u9_X_40, u0_u9_X_42, 
       u0_u9_X_44, u0_u9_X_45, u0_u9_X_47, u0_u9_X_48, u0_u9_X_6, u0_u9_X_8, u0_u9_X_9, u0_u9_u0_n100, u0_u9_u0_n101, 
       u0_u9_u0_n102, u0_u9_u0_n103, u0_u9_u0_n104, u0_u9_u0_n105, u0_u9_u0_n106, u0_u9_u0_n107, u0_u9_u0_n108, u0_u9_u0_n109, u0_u9_u0_n110, 
       u0_u9_u0_n111, u0_u9_u0_n112, u0_u9_u0_n113, u0_u9_u0_n114, u0_u9_u0_n115, u0_u9_u0_n116, u0_u9_u0_n117, u0_u9_u0_n118, u0_u9_u0_n119, 
       u0_u9_u0_n120, u0_u9_u0_n121, u0_u9_u0_n122, u0_u9_u0_n123, u0_u9_u0_n124, u0_u9_u0_n125, u0_u9_u0_n126, u0_u9_u0_n127, u0_u9_u0_n128, 
       u0_u9_u0_n129, u0_u9_u0_n130, u0_u9_u0_n131, u0_u9_u0_n132, u0_u9_u0_n133, u0_u9_u0_n134, u0_u9_u0_n135, u0_u9_u0_n136, u0_u9_u0_n137, 
       u0_u9_u0_n138, u0_u9_u0_n139, u0_u9_u0_n140, u0_u9_u0_n141, u0_u9_u0_n142, u0_u9_u0_n143, u0_u9_u0_n144, u0_u9_u0_n145, u0_u9_u0_n146, 
       u0_u9_u0_n147, u0_u9_u0_n148, u0_u9_u0_n149, u0_u9_u0_n150, u0_u9_u0_n151, u0_u9_u0_n152, u0_u9_u0_n153, u0_u9_u0_n154, u0_u9_u0_n155, 
       u0_u9_u0_n156, u0_u9_u0_n157, u0_u9_u0_n158, u0_u9_u0_n159, u0_u9_u0_n160, u0_u9_u0_n161, u0_u9_u0_n162, u0_u9_u0_n163, u0_u9_u0_n164, 
       u0_u9_u0_n165, u0_u9_u0_n166, u0_u9_u0_n167, u0_u9_u0_n168, u0_u9_u0_n169, u0_u9_u0_n170, u0_u9_u0_n171, u0_u9_u0_n172, u0_u9_u0_n173, 
       u0_u9_u0_n174, u0_u9_u0_n88, u0_u9_u0_n89, u0_u9_u0_n90, u0_u9_u0_n91, u0_u9_u0_n92, u0_u9_u0_n93, u0_u9_u0_n94, u0_u9_u0_n95, 
       u0_u9_u0_n96, u0_u9_u0_n97, u0_u9_u0_n98, u0_u9_u0_n99, u0_u9_u1_n100, u0_u9_u1_n101, u0_u9_u1_n102, u0_u9_u1_n103, u0_u9_u1_n104, 
       u0_u9_u1_n105, u0_u9_u1_n106, u0_u9_u1_n107, u0_u9_u1_n108, u0_u9_u1_n109, u0_u9_u1_n110, u0_u9_u1_n111, u0_u9_u1_n112, u0_u9_u1_n113, 
       u0_u9_u1_n114, u0_u9_u1_n115, u0_u9_u1_n116, u0_u9_u1_n117, u0_u9_u1_n118, u0_u9_u1_n119, u0_u9_u1_n120, u0_u9_u1_n121, u0_u9_u1_n122, 
       u0_u9_u1_n123, u0_u9_u1_n124, u0_u9_u1_n125, u0_u9_u1_n126, u0_u9_u1_n127, u0_u9_u1_n128, u0_u9_u1_n129, u0_u9_u1_n130, u0_u9_u1_n131, 
       u0_u9_u1_n132, u0_u9_u1_n133, u0_u9_u1_n134, u0_u9_u1_n135, u0_u9_u1_n136, u0_u9_u1_n137, u0_u9_u1_n138, u0_u9_u1_n139, u0_u9_u1_n140, 
       u0_u9_u1_n141, u0_u9_u1_n142, u0_u9_u1_n143, u0_u9_u1_n144, u0_u9_u1_n145, u0_u9_u1_n146, u0_u9_u1_n147, u0_u9_u1_n148, u0_u9_u1_n149, 
       u0_u9_u1_n150, u0_u9_u1_n151, u0_u9_u1_n152, u0_u9_u1_n153, u0_u9_u1_n154, u0_u9_u1_n155, u0_u9_u1_n156, u0_u9_u1_n157, u0_u9_u1_n158, 
       u0_u9_u1_n159, u0_u9_u1_n160, u0_u9_u1_n161, u0_u9_u1_n162, u0_u9_u1_n163, u0_u9_u1_n164, u0_u9_u1_n165, u0_u9_u1_n166, u0_u9_u1_n167, 
       u0_u9_u1_n168, u0_u9_u1_n169, u0_u9_u1_n170, u0_u9_u1_n171, u0_u9_u1_n172, u0_u9_u1_n173, u0_u9_u1_n174, u0_u9_u1_n175, u0_u9_u1_n176, 
       u0_u9_u1_n177, u0_u9_u1_n178, u0_u9_u1_n179, u0_u9_u1_n180, u0_u9_u1_n181, u0_u9_u1_n182, u0_u9_u1_n183, u0_u9_u1_n184, u0_u9_u1_n185, 
       u0_u9_u1_n186, u0_u9_u1_n187, u0_u9_u1_n188, u0_u9_u1_n95, u0_u9_u1_n96, u0_u9_u1_n97, u0_u9_u1_n98, u0_u9_u1_n99, u0_u9_u2_n100, 
       u0_u9_u2_n101, u0_u9_u2_n102, u0_u9_u2_n103, u0_u9_u2_n104, u0_u9_u2_n105, u0_u9_u2_n106, u0_u9_u2_n107, u0_u9_u2_n108, u0_u9_u2_n109, 
       u0_u9_u2_n110, u0_u9_u2_n111, u0_u9_u2_n112, u0_u9_u2_n113, u0_u9_u2_n114, u0_u9_u2_n115, u0_u9_u2_n116, u0_u9_u2_n117, u0_u9_u2_n118, 
       u0_u9_u2_n119, u0_u9_u2_n120, u0_u9_u2_n121, u0_u9_u2_n122, u0_u9_u2_n123, u0_u9_u2_n124, u0_u9_u2_n125, u0_u9_u2_n126, u0_u9_u2_n127, 
       u0_u9_u2_n128, u0_u9_u2_n129, u0_u9_u2_n130, u0_u9_u2_n131, u0_u9_u2_n132, u0_u9_u2_n133, u0_u9_u2_n134, u0_u9_u2_n135, u0_u9_u2_n136, 
       u0_u9_u2_n137, u0_u9_u2_n138, u0_u9_u2_n139, u0_u9_u2_n140, u0_u9_u2_n141, u0_u9_u2_n142, u0_u9_u2_n143, u0_u9_u2_n144, u0_u9_u2_n145, 
       u0_u9_u2_n146, u0_u9_u2_n147, u0_u9_u2_n148, u0_u9_u2_n149, u0_u9_u2_n150, u0_u9_u2_n151, u0_u9_u2_n152, u0_u9_u2_n153, u0_u9_u2_n154, 
       u0_u9_u2_n155, u0_u9_u2_n156, u0_u9_u2_n157, u0_u9_u2_n158, u0_u9_u2_n159, u0_u9_u2_n160, u0_u9_u2_n161, u0_u9_u2_n162, u0_u9_u2_n163, 
       u0_u9_u2_n164, u0_u9_u2_n165, u0_u9_u2_n166, u0_u9_u2_n167, u0_u9_u2_n168, u0_u9_u2_n169, u0_u9_u2_n170, u0_u9_u2_n171, u0_u9_u2_n172, 
       u0_u9_u2_n173, u0_u9_u2_n174, u0_u9_u2_n175, u0_u9_u2_n176, u0_u9_u2_n177, u0_u9_u2_n178, u0_u9_u2_n179, u0_u9_u2_n180, u0_u9_u2_n181, 
       u0_u9_u2_n182, u0_u9_u2_n183, u0_u9_u2_n184, u0_u9_u2_n185, u0_u9_u2_n186, u0_u9_u2_n187, u0_u9_u2_n188, u0_u9_u2_n95, u0_u9_u2_n96, 
       u0_u9_u2_n97, u0_u9_u2_n98, u0_u9_u2_n99, u0_u9_u3_n100, u0_u9_u3_n101, u0_u9_u3_n102, u0_u9_u3_n103, u0_u9_u3_n104, u0_u9_u3_n105, 
       u0_u9_u3_n106, u0_u9_u3_n107, u0_u9_u3_n108, u0_u9_u3_n109, u0_u9_u3_n110, u0_u9_u3_n111, u0_u9_u3_n112, u0_u9_u3_n113, u0_u9_u3_n114, 
       u0_u9_u3_n115, u0_u9_u3_n116, u0_u9_u3_n117, u0_u9_u3_n118, u0_u9_u3_n119, u0_u9_u3_n120, u0_u9_u3_n121, u0_u9_u3_n122, u0_u9_u3_n123, 
       u0_u9_u3_n124, u0_u9_u3_n125, u0_u9_u3_n126, u0_u9_u3_n127, u0_u9_u3_n128, u0_u9_u3_n129, u0_u9_u3_n130, u0_u9_u3_n131, u0_u9_u3_n132, 
       u0_u9_u3_n133, u0_u9_u3_n134, u0_u9_u3_n135, u0_u9_u3_n136, u0_u9_u3_n137, u0_u9_u3_n138, u0_u9_u3_n139, u0_u9_u3_n140, u0_u9_u3_n141, 
       u0_u9_u3_n142, u0_u9_u3_n143, u0_u9_u3_n144, u0_u9_u3_n145, u0_u9_u3_n146, u0_u9_u3_n147, u0_u9_u3_n148, u0_u9_u3_n149, u0_u9_u3_n150, 
       u0_u9_u3_n151, u0_u9_u3_n152, u0_u9_u3_n153, u0_u9_u3_n154, u0_u9_u3_n155, u0_u9_u3_n156, u0_u9_u3_n157, u0_u9_u3_n158, u0_u9_u3_n159, 
       u0_u9_u3_n160, u0_u9_u3_n161, u0_u9_u3_n162, u0_u9_u3_n163, u0_u9_u3_n164, u0_u9_u3_n165, u0_u9_u3_n166, u0_u9_u3_n167, u0_u9_u3_n168, 
       u0_u9_u3_n169, u0_u9_u3_n170, u0_u9_u3_n171, u0_u9_u3_n172, u0_u9_u3_n173, u0_u9_u3_n174, u0_u9_u3_n175, u0_u9_u3_n176, u0_u9_u3_n177, 
       u0_u9_u3_n178, u0_u9_u3_n179, u0_u9_u3_n180, u0_u9_u3_n181, u0_u9_u3_n182, u0_u9_u3_n183, u0_u9_u3_n184, u0_u9_u3_n185, u0_u9_u3_n186, 
       u0_u9_u3_n94, u0_u9_u3_n95, u0_u9_u3_n96, u0_u9_u3_n97, u0_u9_u3_n98, u0_u9_u3_n99, u0_u9_u4_n100, u0_u9_u4_n101, u0_u9_u4_n102, 
       u0_u9_u4_n103, u0_u9_u4_n104, u0_u9_u4_n105, u0_u9_u4_n106, u0_u9_u4_n107, u0_u9_u4_n108, u0_u9_u4_n109, u0_u9_u4_n110, u0_u9_u4_n111, 
       u0_u9_u4_n112, u0_u9_u4_n113, u0_u9_u4_n114, u0_u9_u4_n115, u0_u9_u4_n116, u0_u9_u4_n117, u0_u9_u4_n118, u0_u9_u4_n119, u0_u9_u4_n120, 
       u0_u9_u4_n121, u0_u9_u4_n122, u0_u9_u4_n123, u0_u9_u4_n124, u0_u9_u4_n125, u0_u9_u4_n126, u0_u9_u4_n127, u0_u9_u4_n128, u0_u9_u4_n129, 
       u0_u9_u4_n130, u0_u9_u4_n131, u0_u9_u4_n132, u0_u9_u4_n133, u0_u9_u4_n134, u0_u9_u4_n135, u0_u9_u4_n136, u0_u9_u4_n137, u0_u9_u4_n138, 
       u0_u9_u4_n139, u0_u9_u4_n140, u0_u9_u4_n141, u0_u9_u4_n142, u0_u9_u4_n143, u0_u9_u4_n144, u0_u9_u4_n145, u0_u9_u4_n146, u0_u9_u4_n147, 
       u0_u9_u4_n148, u0_u9_u4_n149, u0_u9_u4_n150, u0_u9_u4_n151, u0_u9_u4_n152, u0_u9_u4_n153, u0_u9_u4_n154, u0_u9_u4_n155, u0_u9_u4_n156, 
       u0_u9_u4_n157, u0_u9_u4_n158, u0_u9_u4_n159, u0_u9_u4_n160, u0_u9_u4_n161, u0_u9_u4_n162, u0_u9_u4_n163, u0_u9_u4_n164, u0_u9_u4_n165, 
       u0_u9_u4_n166, u0_u9_u4_n167, u0_u9_u4_n168, u0_u9_u4_n169, u0_u9_u4_n170, u0_u9_u4_n171, u0_u9_u4_n172, u0_u9_u4_n173, u0_u9_u4_n174, 
       u0_u9_u4_n175, u0_u9_u4_n176, u0_u9_u4_n177, u0_u9_u4_n178, u0_u9_u4_n179, u0_u9_u4_n180, u0_u9_u4_n181, u0_u9_u4_n182, u0_u9_u4_n183, 
       u0_u9_u4_n184, u0_u9_u4_n185, u0_u9_u4_n186, u0_u9_u4_n94, u0_u9_u4_n95, u0_u9_u4_n96, u0_u9_u4_n97, u0_u9_u4_n98, u0_u9_u4_n99, 
       u0_u9_u5_n100, u0_u9_u5_n101, u0_u9_u5_n102, u0_u9_u5_n103, u0_u9_u5_n104, u0_u9_u5_n105, u0_u9_u5_n106, u0_u9_u5_n107, u0_u9_u5_n108, 
       u0_u9_u5_n109, u0_u9_u5_n110, u0_u9_u5_n111, u0_u9_u5_n112, u0_u9_u5_n113, u0_u9_u5_n114, u0_u9_u5_n115, u0_u9_u5_n116, u0_u9_u5_n117, 
       u0_u9_u5_n118, u0_u9_u5_n119, u0_u9_u5_n120, u0_u9_u5_n121, u0_u9_u5_n122, u0_u9_u5_n123, u0_u9_u5_n124, u0_u9_u5_n125, u0_u9_u5_n126, 
       u0_u9_u5_n127, u0_u9_u5_n128, u0_u9_u5_n129, u0_u9_u5_n130, u0_u9_u5_n131, u0_u9_u5_n132, u0_u9_u5_n133, u0_u9_u5_n134, u0_u9_u5_n135, 
       u0_u9_u5_n136, u0_u9_u5_n137, u0_u9_u5_n138, u0_u9_u5_n139, u0_u9_u5_n140, u0_u9_u5_n141, u0_u9_u5_n142, u0_u9_u5_n143, u0_u9_u5_n144, 
       u0_u9_u5_n145, u0_u9_u5_n146, u0_u9_u5_n147, u0_u9_u5_n148, u0_u9_u5_n149, u0_u9_u5_n150, u0_u9_u5_n151, u0_u9_u5_n152, u0_u9_u5_n153, 
       u0_u9_u5_n154, u0_u9_u5_n155, u0_u9_u5_n156, u0_u9_u5_n157, u0_u9_u5_n158, u0_u9_u5_n159, u0_u9_u5_n160, u0_u9_u5_n161, u0_u9_u5_n162, 
       u0_u9_u5_n163, u0_u9_u5_n164, u0_u9_u5_n165, u0_u9_u5_n166, u0_u9_u5_n167, u0_u9_u5_n168, u0_u9_u5_n169, u0_u9_u5_n170, u0_u9_u5_n171, 
       u0_u9_u5_n172, u0_u9_u5_n173, u0_u9_u5_n174, u0_u9_u5_n175, u0_u9_u5_n176, u0_u9_u5_n177, u0_u9_u5_n178, u0_u9_u5_n179, u0_u9_u5_n180, 
       u0_u9_u5_n181, u0_u9_u5_n182, u0_u9_u5_n183, u0_u9_u5_n184, u0_u9_u5_n185, u0_u9_u5_n186, u0_u9_u5_n187, u0_u9_u5_n188, u0_u9_u5_n189, 
       u0_u9_u5_n190, u0_u9_u5_n191, u0_u9_u5_n192, u0_u9_u5_n193, u0_u9_u5_n194, u0_u9_u5_n195, u0_u9_u5_n196, u0_u9_u5_n99, u0_u9_u6_n100, 
       u0_u9_u6_n101, u0_u9_u6_n102, u0_u9_u6_n103, u0_u9_u6_n104, u0_u9_u6_n105, u0_u9_u6_n106, u0_u9_u6_n107, u0_u9_u6_n108, u0_u9_u6_n109, 
       u0_u9_u6_n110, u0_u9_u6_n111, u0_u9_u6_n112, u0_u9_u6_n113, u0_u9_u6_n114, u0_u9_u6_n115, u0_u9_u6_n116, u0_u9_u6_n117, u0_u9_u6_n118, 
       u0_u9_u6_n119, u0_u9_u6_n120, u0_u9_u6_n121, u0_u9_u6_n122, u0_u9_u6_n123, u0_u9_u6_n124, u0_u9_u6_n125, u0_u9_u6_n126, u0_u9_u6_n127, 
       u0_u9_u6_n128, u0_u9_u6_n129, u0_u9_u6_n130, u0_u9_u6_n131, u0_u9_u6_n132, u0_u9_u6_n133, u0_u9_u6_n134, u0_u9_u6_n135, u0_u9_u6_n136, 
       u0_u9_u6_n137, u0_u9_u6_n138, u0_u9_u6_n139, u0_u9_u6_n140, u0_u9_u6_n141, u0_u9_u6_n142, u0_u9_u6_n143, u0_u9_u6_n144, u0_u9_u6_n145, 
       u0_u9_u6_n146, u0_u9_u6_n147, u0_u9_u6_n148, u0_u9_u6_n149, u0_u9_u6_n150, u0_u9_u6_n151, u0_u9_u6_n152, u0_u9_u6_n153, u0_u9_u6_n154, 
       u0_u9_u6_n155, u0_u9_u6_n156, u0_u9_u6_n157, u0_u9_u6_n158, u0_u9_u6_n159, u0_u9_u6_n160, u0_u9_u6_n161, u0_u9_u6_n162, u0_u9_u6_n163, 
       u0_u9_u6_n164, u0_u9_u6_n165, u0_u9_u6_n166, u0_u9_u6_n167, u0_u9_u6_n168, u0_u9_u6_n169, u0_u9_u6_n170, u0_u9_u6_n171, u0_u9_u6_n172, 
       u0_u9_u6_n173, u0_u9_u6_n174, u0_u9_u6_n88, u0_u9_u6_n89, u0_u9_u6_n90, u0_u9_u6_n91, u0_u9_u6_n92, u0_u9_u6_n93, u0_u9_u6_n94, 
       u0_u9_u6_n95, u0_u9_u6_n96, u0_u9_u6_n97, u0_u9_u6_n98, u0_u9_u6_n99, u0_u9_u7_n100, u0_u9_u7_n101, u0_u9_u7_n102, u0_u9_u7_n103, 
       u0_u9_u7_n104, u0_u9_u7_n105, u0_u9_u7_n106, u0_u9_u7_n107, u0_u9_u7_n108, u0_u9_u7_n109, u0_u9_u7_n110, u0_u9_u7_n111, u0_u9_u7_n112, 
       u0_u9_u7_n113, u0_u9_u7_n114, u0_u9_u7_n115, u0_u9_u7_n116, u0_u9_u7_n117, u0_u9_u7_n118, u0_u9_u7_n119, u0_u9_u7_n120, u0_u9_u7_n121, 
       u0_u9_u7_n122, u0_u9_u7_n123, u0_u9_u7_n124, u0_u9_u7_n125, u0_u9_u7_n126, u0_u9_u7_n127, u0_u9_u7_n128, u0_u9_u7_n129, u0_u9_u7_n130, 
       u0_u9_u7_n131, u0_u9_u7_n132, u0_u9_u7_n133, u0_u9_u7_n134, u0_u9_u7_n135, u0_u9_u7_n136, u0_u9_u7_n137, u0_u9_u7_n138, u0_u9_u7_n139, 
       u0_u9_u7_n140, u0_u9_u7_n141, u0_u9_u7_n142, u0_u9_u7_n143, u0_u9_u7_n144, u0_u9_u7_n145, u0_u9_u7_n146, u0_u9_u7_n147, u0_u9_u7_n148, 
       u0_u9_u7_n149, u0_u9_u7_n150, u0_u9_u7_n151, u0_u9_u7_n152, u0_u9_u7_n153, u0_u9_u7_n154, u0_u9_u7_n155, u0_u9_u7_n156, u0_u9_u7_n157, 
       u0_u9_u7_n158, u0_u9_u7_n159, u0_u9_u7_n160, u0_u9_u7_n161, u0_u9_u7_n162, u0_u9_u7_n163, u0_u9_u7_n164, u0_u9_u7_n165, u0_u9_u7_n166, 
       u0_u9_u7_n167, u0_u9_u7_n168, u0_u9_u7_n169, u0_u9_u7_n170, u0_u9_u7_n171, u0_u9_u7_n172, u0_u9_u7_n173, u0_u9_u7_n174, u0_u9_u7_n175, 
       u0_u9_u7_n176, u0_u9_u7_n177, u0_u9_u7_n178, u0_u9_u7_n179, u0_u9_u7_n180, u0_u9_u7_n91, u0_u9_u7_n92, u0_u9_u7_n93, u0_u9_u7_n94, 
       u0_u9_u7_n95, u0_u9_u7_n96, u0_u9_u7_n97, u0_u9_u7_n98, u0_u9_u7_n99, u0_uk_n1014, u0_uk_n1015, u0_uk_n1017, u0_uk_n757, 
       u0_uk_n758, u0_uk_n760, u0_uk_n764, u0_uk_n781, u0_uk_n784, u0_uk_n803, u0_uk_n811, u0_uk_n819, u0_uk_n821, 
       u0_uk_n822, u0_uk_n824, u0_uk_n825, u0_uk_n827, u0_uk_n828, u0_uk_n833, u0_uk_n835, u0_uk_n836, u0_uk_n837, 
       u0_uk_n838, u0_uk_n919, u0_uk_n920, u2_K10_2, u2_K10_31, u2_K10_33, u2_K10_35, u2_K10_37, u2_K10_38, 
       u2_K10_39, u2_K10_40, u2_K10_41, u2_K10_47, u2_K11_19, u2_K11_20, u2_K11_31, u2_K11_47, u2_K12_1, 
       u2_K12_10, u2_K12_11, u2_K12_12, u2_K12_13, u2_K12_14, u2_K12_17, u2_K12_18, u2_K12_19, u2_K12_23, 
       u2_K12_30, u2_K12_32, u2_K12_4, u2_K12_42, u2_K12_44, u2_K12_5, u2_K12_7, u2_K13_2, u2_K13_30, 
       u2_K13_5, u2_K13_7, u2_K14_29, u2_K14_30, u2_K14_31, u2_K14_32, u2_K14_33, u2_K14_36, u2_K15_14, 
       u2_K15_19, u2_K15_24, u2_K15_25, u2_K15_26, u2_K15_33, u2_K15_36, u2_K15_37, u2_K15_38, u2_K15_40, 
       u2_K15_42, u2_K15_47, u2_K15_48, u2_K15_6, u2_K15_8, u2_K1_29, u2_K1_31, u2_K1_36, u2_K1_38, 
       u2_K1_41, u2_K1_42, u2_K1_44, u2_K1_47, u2_K3_1, u2_K3_10, u2_K3_11, u2_K3_12, u2_K3_14, 
       u2_K3_17, u2_K3_18, u2_K3_2, u2_K3_21, u2_K3_22, u2_K3_24, u2_K3_25, u2_K3_3, u2_K3_36, 
       u2_K3_38, u2_K3_4, u2_K3_40, u2_K3_41, u2_K3_44, u2_K3_45, u2_K3_46, u2_K3_6, u2_K3_8, 
       u2_K3_9, u2_K4_1, u2_K4_10, u2_K4_11, u2_K4_12, u2_K4_13, u2_K4_15, u2_K4_16, u2_K4_17, 
       u2_K4_2, u2_K4_20, u2_K4_23, u2_K4_25, u2_K4_26, u2_K4_28, u2_K4_29, u2_K4_3, u2_K4_30, 
       u2_K4_31, u2_K4_32, u2_K4_36, u2_K4_4, u2_K4_47, u2_K4_5, u2_K4_8, u2_K4_9, u2_K5_12, 
       u2_K5_20, u2_K5_27, u2_K5_33, u2_K5_35, u2_K5_36, u2_K5_42, u2_K5_43, u2_K5_45, u2_K5_7, 
       u2_K6_12, u2_K6_17, u2_K6_18, u2_K6_2, u2_K6_21, u2_K6_26, u2_K6_30, u2_K6_33, u2_K6_35, 
       u2_K6_37, u2_K6_41, u2_K6_42, u2_K6_43, u2_K6_44, u2_K6_46, u2_K6_48, u2_K6_5, u2_K6_7, 
       u2_K6_9, u2_K7_1, u2_K7_11, u2_K7_12, u2_K7_13, u2_K7_14, u2_K7_15, u2_K7_16, u2_K7_17, 
       u2_K7_18, u2_K7_19, u2_K7_2, u2_K7_20, u2_K7_21, u2_K7_23, u2_K7_24, u2_K7_25, u2_K7_29, 
       u2_K7_32, u2_K7_34, u2_K7_36, u2_K7_39, u2_K7_41, u2_K7_42, u2_K7_44, u2_K7_47, u2_K7_6, 
       u2_K7_8, u2_K9_10, u2_K9_11, u2_K9_13, u2_K9_16, u2_K9_17, u2_K9_18, u2_K9_19, u2_K9_2, 
       u2_K9_20, u2_K9_21, u2_K9_22, u2_K9_24, u2_K9_26, u2_K9_4, u2_K9_6, u2_K9_7, u2_K9_8, 
       u2_K9_9, u2_u0_X_29, u2_u0_X_31, u2_u0_X_36, u2_u0_X_38, u2_u0_X_41, u2_u0_X_42, u2_u0_X_43, u2_u0_X_44, 
       u2_u0_X_47, u2_u0_u1_n100, u2_u0_u1_n101, u2_u0_u1_n102, u2_u0_u1_n103, u2_u0_u1_n104, u2_u0_u1_n105, u2_u0_u1_n106, u2_u0_u1_n107, 
       u2_u0_u1_n108, u2_u0_u1_n109, u2_u0_u1_n110, u2_u0_u1_n111, u2_u0_u1_n112, u2_u0_u1_n113, u2_u0_u1_n114, u2_u0_u1_n115, u2_u0_u1_n116, 
       u2_u0_u1_n117, u2_u0_u1_n118, u2_u0_u1_n119, u2_u0_u1_n120, u2_u0_u1_n121, u2_u0_u1_n122, u2_u0_u1_n123, u2_u0_u1_n124, u2_u0_u1_n125, 
       u2_u0_u1_n126, u2_u0_u1_n127, u2_u0_u1_n128, u2_u0_u1_n129, u2_u0_u1_n130, u2_u0_u1_n131, u2_u0_u1_n132, u2_u0_u1_n133, u2_u0_u1_n134, 
       u2_u0_u1_n135, u2_u0_u1_n136, u2_u0_u1_n137, u2_u0_u1_n138, u2_u0_u1_n139, u2_u0_u1_n140, u2_u0_u1_n141, u2_u0_u1_n142, u2_u0_u1_n143, 
       u2_u0_u1_n144, u2_u0_u1_n145, u2_u0_u1_n146, u2_u0_u1_n147, u2_u0_u1_n148, u2_u0_u1_n149, u2_u0_u1_n150, u2_u0_u1_n151, u2_u0_u1_n152, 
       u2_u0_u1_n153, u2_u0_u1_n154, u2_u0_u1_n155, u2_u0_u1_n156, u2_u0_u1_n157, u2_u0_u1_n158, u2_u0_u1_n159, u2_u0_u1_n160, u2_u0_u1_n161, 
       u2_u0_u1_n162, u2_u0_u1_n163, u2_u0_u1_n164, u2_u0_u1_n165, u2_u0_u1_n166, u2_u0_u1_n167, u2_u0_u1_n168, u2_u0_u1_n169, u2_u0_u1_n170, 
       u2_u0_u1_n171, u2_u0_u1_n172, u2_u0_u1_n173, u2_u0_u1_n174, u2_u0_u1_n175, u2_u0_u1_n176, u2_u0_u1_n177, u2_u0_u1_n178, u2_u0_u1_n179, 
       u2_u0_u1_n180, u2_u0_u1_n181, u2_u0_u1_n182, u2_u0_u1_n183, u2_u0_u1_n184, u2_u0_u1_n185, u2_u0_u1_n186, u2_u0_u1_n187, u2_u0_u1_n188, 
       u2_u0_u1_n95, u2_u0_u1_n96, u2_u0_u1_n97, u2_u0_u1_n98, u2_u0_u1_n99, u2_u0_u4_n100, u2_u0_u4_n101, u2_u0_u4_n102, u2_u0_u4_n103, 
       u2_u0_u4_n104, u2_u0_u4_n105, u2_u0_u4_n106, u2_u0_u4_n107, u2_u0_u4_n108, u2_u0_u4_n109, u2_u0_u4_n110, u2_u0_u4_n111, u2_u0_u4_n112, 
       u2_u0_u4_n113, u2_u0_u4_n114, u2_u0_u4_n115, u2_u0_u4_n116, u2_u0_u4_n117, u2_u0_u4_n118, u2_u0_u4_n119, u2_u0_u4_n120, u2_u0_u4_n121, 
       u2_u0_u4_n122, u2_u0_u4_n123, u2_u0_u4_n124, u2_u0_u4_n125, u2_u0_u4_n126, u2_u0_u4_n127, u2_u0_u4_n128, u2_u0_u4_n129, u2_u0_u4_n130, 
       u2_u0_u4_n131, u2_u0_u4_n132, u2_u0_u4_n133, u2_u0_u4_n134, u2_u0_u4_n135, u2_u0_u4_n136, u2_u0_u4_n137, u2_u0_u4_n138, u2_u0_u4_n139, 
       u2_u0_u4_n140, u2_u0_u4_n141, u2_u0_u4_n142, u2_u0_u4_n143, u2_u0_u4_n144, u2_u0_u4_n145, u2_u0_u4_n146, u2_u0_u4_n147, u2_u0_u4_n148, 
       u2_u0_u4_n149, u2_u0_u4_n150, u2_u0_u4_n151, u2_u0_u4_n152, u2_u0_u4_n153, u2_u0_u4_n154, u2_u0_u4_n155, u2_u0_u4_n156, u2_u0_u4_n157, 
       u2_u0_u4_n158, u2_u0_u4_n159, u2_u0_u4_n160, u2_u0_u4_n161, u2_u0_u4_n162, u2_u0_u4_n163, u2_u0_u4_n164, u2_u0_u4_n165, u2_u0_u4_n166, 
       u2_u0_u4_n167, u2_u0_u4_n168, u2_u0_u4_n169, u2_u0_u4_n170, u2_u0_u4_n171, u2_u0_u4_n172, u2_u0_u4_n173, u2_u0_u4_n174, u2_u0_u4_n175, 
       u2_u0_u4_n176, u2_u0_u4_n177, u2_u0_u4_n178, u2_u0_u4_n179, u2_u0_u4_n180, u2_u0_u4_n181, u2_u0_u4_n182, u2_u0_u4_n183, u2_u0_u4_n184, 
       u2_u0_u4_n185, u2_u0_u4_n186, u2_u0_u4_n94, u2_u0_u4_n95, u2_u0_u4_n96, u2_u0_u4_n97, u2_u0_u4_n98, u2_u0_u4_n99, u2_u0_u5_n100, 
       u2_u0_u5_n101, u2_u0_u5_n102, u2_u0_u5_n103, u2_u0_u5_n104, u2_u0_u5_n105, u2_u0_u5_n106, u2_u0_u5_n107, u2_u0_u5_n108, u2_u0_u5_n109, 
       u2_u0_u5_n110, u2_u0_u5_n111, u2_u0_u5_n112, u2_u0_u5_n113, u2_u0_u5_n114, u2_u0_u5_n115, u2_u0_u5_n116, u2_u0_u5_n117, u2_u0_u5_n118, 
       u2_u0_u5_n119, u2_u0_u5_n120, u2_u0_u5_n121, u2_u0_u5_n122, u2_u0_u5_n123, u2_u0_u5_n124, u2_u0_u5_n125, u2_u0_u5_n126, u2_u0_u5_n127, 
       u2_u0_u5_n128, u2_u0_u5_n129, u2_u0_u5_n130, u2_u0_u5_n131, u2_u0_u5_n132, u2_u0_u5_n133, u2_u0_u5_n134, u2_u0_u5_n135, u2_u0_u5_n136, 
       u2_u0_u5_n137, u2_u0_u5_n138, u2_u0_u5_n139, u2_u0_u5_n140, u2_u0_u5_n141, u2_u0_u5_n142, u2_u0_u5_n143, u2_u0_u5_n144, u2_u0_u5_n145, 
       u2_u0_u5_n146, u2_u0_u5_n147, u2_u0_u5_n148, u2_u0_u5_n149, u2_u0_u5_n150, u2_u0_u5_n151, u2_u0_u5_n152, u2_u0_u5_n153, u2_u0_u5_n154, 
       u2_u0_u5_n155, u2_u0_u5_n156, u2_u0_u5_n157, u2_u0_u5_n158, u2_u0_u5_n159, u2_u0_u5_n160, u2_u0_u5_n161, u2_u0_u5_n162, u2_u0_u5_n163, 
       u2_u0_u5_n164, u2_u0_u5_n165, u2_u0_u5_n166, u2_u0_u5_n167, u2_u0_u5_n168, u2_u0_u5_n169, u2_u0_u5_n170, u2_u0_u5_n171, u2_u0_u5_n172, 
       u2_u0_u5_n173, u2_u0_u5_n174, u2_u0_u5_n175, u2_u0_u5_n176, u2_u0_u5_n177, u2_u0_u5_n178, u2_u0_u5_n179, u2_u0_u5_n180, u2_u0_u5_n181, 
       u2_u0_u5_n182, u2_u0_u5_n183, u2_u0_u5_n184, u2_u0_u5_n185, u2_u0_u5_n186, u2_u0_u5_n187, u2_u0_u5_n188, u2_u0_u5_n189, u2_u0_u5_n190, 
       u2_u0_u5_n191, u2_u0_u5_n192, u2_u0_u5_n193, u2_u0_u5_n194, u2_u0_u5_n195, u2_u0_u5_n196, u2_u0_u5_n99, u2_u0_u6_n100, u2_u0_u6_n101, 
       u2_u0_u6_n102, u2_u0_u6_n103, u2_u0_u6_n104, u2_u0_u6_n105, u2_u0_u6_n106, u2_u0_u6_n107, u2_u0_u6_n108, u2_u0_u6_n109, u2_u0_u6_n110, 
       u2_u0_u6_n111, u2_u0_u6_n112, u2_u0_u6_n113, u2_u0_u6_n114, u2_u0_u6_n115, u2_u0_u6_n116, u2_u0_u6_n117, u2_u0_u6_n118, u2_u0_u6_n119, 
       u2_u0_u6_n120, u2_u0_u6_n121, u2_u0_u6_n122, u2_u0_u6_n123, u2_u0_u6_n124, u2_u0_u6_n125, u2_u0_u6_n126, u2_u0_u6_n127, u2_u0_u6_n128, 
       u2_u0_u6_n129, u2_u0_u6_n130, u2_u0_u6_n131, u2_u0_u6_n132, u2_u0_u6_n133, u2_u0_u6_n134, u2_u0_u6_n135, u2_u0_u6_n136, u2_u0_u6_n137, 
       u2_u0_u6_n138, u2_u0_u6_n139, u2_u0_u6_n140, u2_u0_u6_n141, u2_u0_u6_n142, u2_u0_u6_n143, u2_u0_u6_n144, u2_u0_u6_n145, u2_u0_u6_n146, 
       u2_u0_u6_n147, u2_u0_u6_n148, u2_u0_u6_n149, u2_u0_u6_n150, u2_u0_u6_n151, u2_u0_u6_n152, u2_u0_u6_n153, u2_u0_u6_n154, u2_u0_u6_n155, 
       u2_u0_u6_n156, u2_u0_u6_n157, u2_u0_u6_n158, u2_u0_u6_n159, u2_u0_u6_n160, u2_u0_u6_n161, u2_u0_u6_n162, u2_u0_u6_n163, u2_u0_u6_n164, 
       u2_u0_u6_n165, u2_u0_u6_n166, u2_u0_u6_n167, u2_u0_u6_n168, u2_u0_u6_n169, u2_u0_u6_n170, u2_u0_u6_n171, u2_u0_u6_n172, u2_u0_u6_n173, 
       u2_u0_u6_n174, u2_u0_u6_n88, u2_u0_u6_n89, u2_u0_u6_n90, u2_u0_u6_n91, u2_u0_u6_n92, u2_u0_u6_n93, u2_u0_u6_n94, u2_u0_u6_n95, 
       u2_u0_u6_n96, u2_u0_u6_n97, u2_u0_u6_n98, u2_u0_u6_n99, u2_u0_u7_n100, u2_u0_u7_n101, u2_u0_u7_n102, u2_u0_u7_n103, u2_u0_u7_n104, 
       u2_u0_u7_n105, u2_u0_u7_n106, u2_u0_u7_n107, u2_u0_u7_n108, u2_u0_u7_n109, u2_u0_u7_n110, u2_u0_u7_n111, u2_u0_u7_n112, u2_u0_u7_n113, 
       u2_u0_u7_n114, u2_u0_u7_n115, u2_u0_u7_n116, u2_u0_u7_n117, u2_u0_u7_n118, u2_u0_u7_n119, u2_u0_u7_n120, u2_u0_u7_n121, u2_u0_u7_n122, 
       u2_u0_u7_n123, u2_u0_u7_n124, u2_u0_u7_n125, u2_u0_u7_n126, u2_u0_u7_n127, u2_u0_u7_n128, u2_u0_u7_n129, u2_u0_u7_n130, u2_u0_u7_n131, 
       u2_u0_u7_n132, u2_u0_u7_n133, u2_u0_u7_n134, u2_u0_u7_n135, u2_u0_u7_n136, u2_u0_u7_n137, u2_u0_u7_n138, u2_u0_u7_n139, u2_u0_u7_n140, 
       u2_u0_u7_n141, u2_u0_u7_n142, u2_u0_u7_n143, u2_u0_u7_n144, u2_u0_u7_n145, u2_u0_u7_n146, u2_u0_u7_n147, u2_u0_u7_n148, u2_u0_u7_n149, 
       u2_u0_u7_n150, u2_u0_u7_n151, u2_u0_u7_n152, u2_u0_u7_n153, u2_u0_u7_n154, u2_u0_u7_n155, u2_u0_u7_n156, u2_u0_u7_n157, u2_u0_u7_n158, 
       u2_u0_u7_n159, u2_u0_u7_n160, u2_u0_u7_n161, u2_u0_u7_n162, u2_u0_u7_n163, u2_u0_u7_n164, u2_u0_u7_n165, u2_u0_u7_n166, u2_u0_u7_n167, 
       u2_u0_u7_n168, u2_u0_u7_n169, u2_u0_u7_n170, u2_u0_u7_n171, u2_u0_u7_n172, u2_u0_u7_n173, u2_u0_u7_n174, u2_u0_u7_n175, u2_u0_u7_n176, 
       u2_u0_u7_n177, u2_u0_u7_n178, u2_u0_u7_n179, u2_u0_u7_n180, u2_u0_u7_n91, u2_u0_u7_n92, u2_u0_u7_n93, u2_u0_u7_n94, u2_u0_u7_n95, 
       u2_u0_u7_n96, u2_u0_u7_n97, u2_u0_u7_n98, u2_u0_u7_n99, u2_u10_X_19, u2_u10_X_20, u2_u10_X_24, u2_u10_X_26, u2_u10_X_29, 
       u2_u10_X_31, u2_u10_X_47, u2_u10_u3_n100, u2_u10_u3_n101, u2_u10_u3_n102, u2_u10_u3_n103, u2_u10_u3_n104, u2_u10_u3_n105, u2_u10_u3_n106, 
       u2_u10_u3_n107, u2_u10_u3_n108, u2_u10_u3_n109, u2_u10_u3_n110, u2_u10_u3_n111, u2_u10_u3_n112, u2_u10_u3_n113, u2_u10_u3_n114, u2_u10_u3_n115, 
       u2_u10_u3_n116, u2_u10_u3_n117, u2_u10_u3_n118, u2_u10_u3_n119, u2_u10_u3_n120, u2_u10_u3_n121, u2_u10_u3_n122, u2_u10_u3_n123, u2_u10_u3_n124, 
       u2_u10_u3_n125, u2_u10_u3_n126, u2_u10_u3_n127, u2_u10_u3_n128, u2_u10_u3_n129, u2_u10_u3_n130, u2_u10_u3_n131, u2_u10_u3_n132, u2_u10_u3_n133, 
       u2_u10_u3_n134, u2_u10_u3_n135, u2_u10_u3_n136, u2_u10_u3_n137, u2_u10_u3_n138, u2_u10_u3_n139, u2_u10_u3_n140, u2_u10_u3_n141, u2_u10_u3_n142, 
       u2_u10_u3_n143, u2_u10_u3_n144, u2_u10_u3_n145, u2_u10_u3_n146, u2_u10_u3_n147, u2_u10_u3_n148, u2_u10_u3_n149, u2_u10_u3_n150, u2_u10_u3_n151, 
       u2_u10_u3_n152, u2_u10_u3_n153, u2_u10_u3_n154, u2_u10_u3_n155, u2_u10_u3_n156, u2_u10_u3_n157, u2_u10_u3_n158, u2_u10_u3_n159, u2_u10_u3_n160, 
       u2_u10_u3_n161, u2_u10_u3_n162, u2_u10_u3_n163, u2_u10_u3_n164, u2_u10_u3_n165, u2_u10_u3_n166, u2_u10_u3_n167, u2_u10_u3_n168, u2_u10_u3_n169, 
       u2_u10_u3_n170, u2_u10_u3_n171, u2_u10_u3_n172, u2_u10_u3_n173, u2_u10_u3_n174, u2_u10_u3_n175, u2_u10_u3_n176, u2_u10_u3_n177, u2_u10_u3_n178, 
       u2_u10_u3_n179, u2_u10_u3_n180, u2_u10_u3_n181, u2_u10_u3_n182, u2_u10_u3_n183, u2_u10_u3_n184, u2_u10_u3_n185, u2_u10_u3_n186, u2_u10_u3_n94, 
       u2_u10_u3_n95, u2_u10_u3_n96, u2_u10_u3_n97, u2_u10_u3_n98, u2_u10_u3_n99, u2_u10_u4_n100, u2_u10_u4_n101, u2_u10_u4_n102, u2_u10_u4_n103, 
       u2_u10_u4_n104, u2_u10_u4_n105, u2_u10_u4_n106, u2_u10_u4_n107, u2_u10_u4_n108, u2_u10_u4_n109, u2_u10_u4_n110, u2_u10_u4_n111, u2_u10_u4_n112, 
       u2_u10_u4_n113, u2_u10_u4_n114, u2_u10_u4_n115, u2_u10_u4_n116, u2_u10_u4_n117, u2_u10_u4_n118, u2_u10_u4_n119, u2_u10_u4_n120, u2_u10_u4_n121, 
       u2_u10_u4_n122, u2_u10_u4_n123, u2_u10_u4_n124, u2_u10_u4_n125, u2_u10_u4_n126, u2_u10_u4_n127, u2_u10_u4_n128, u2_u10_u4_n129, u2_u10_u4_n130, 
       u2_u10_u4_n131, u2_u10_u4_n132, u2_u10_u4_n133, u2_u10_u4_n134, u2_u10_u4_n135, u2_u10_u4_n136, u2_u10_u4_n137, u2_u10_u4_n138, u2_u10_u4_n139, 
       u2_u10_u4_n140, u2_u10_u4_n141, u2_u10_u4_n142, u2_u10_u4_n143, u2_u10_u4_n144, u2_u10_u4_n145, u2_u10_u4_n146, u2_u10_u4_n147, u2_u10_u4_n148, 
       u2_u10_u4_n149, u2_u10_u4_n150, u2_u10_u4_n151, u2_u10_u4_n152, u2_u10_u4_n153, u2_u10_u4_n154, u2_u10_u4_n155, u2_u10_u4_n156, u2_u10_u4_n157, 
       u2_u10_u4_n158, u2_u10_u4_n159, u2_u10_u4_n160, u2_u10_u4_n161, u2_u10_u4_n162, u2_u10_u4_n163, u2_u10_u4_n164, u2_u10_u4_n165, u2_u10_u4_n166, 
       u2_u10_u4_n167, u2_u10_u4_n168, u2_u10_u4_n169, u2_u10_u4_n170, u2_u10_u4_n171, u2_u10_u4_n172, u2_u10_u4_n173, u2_u10_u4_n174, u2_u10_u4_n175, 
       u2_u10_u4_n176, u2_u10_u4_n177, u2_u10_u4_n178, u2_u10_u4_n179, u2_u10_u4_n180, u2_u10_u4_n181, u2_u10_u4_n182, u2_u10_u4_n183, u2_u10_u4_n184, 
       u2_u10_u4_n185, u2_u10_u4_n186, u2_u10_u4_n94, u2_u10_u4_n95, u2_u10_u4_n96, u2_u10_u4_n97, u2_u10_u4_n98, u2_u10_u4_n99, u2_u10_u5_n100, 
       u2_u10_u5_n101, u2_u10_u5_n102, u2_u10_u5_n103, u2_u10_u5_n104, u2_u10_u5_n105, u2_u10_u5_n106, u2_u10_u5_n107, u2_u10_u5_n108, u2_u10_u5_n109, 
       u2_u10_u5_n110, u2_u10_u5_n111, u2_u10_u5_n112, u2_u10_u5_n113, u2_u10_u5_n114, u2_u10_u5_n115, u2_u10_u5_n116, u2_u10_u5_n117, u2_u10_u5_n118, 
       u2_u10_u5_n119, u2_u10_u5_n120, u2_u10_u5_n121, u2_u10_u5_n122, u2_u10_u5_n123, u2_u10_u5_n124, u2_u10_u5_n125, u2_u10_u5_n126, u2_u10_u5_n127, 
       u2_u10_u5_n128, u2_u10_u5_n129, u2_u10_u5_n130, u2_u10_u5_n131, u2_u10_u5_n132, u2_u10_u5_n133, u2_u10_u5_n134, u2_u10_u5_n135, u2_u10_u5_n136, 
       u2_u10_u5_n137, u2_u10_u5_n138, u2_u10_u5_n139, u2_u10_u5_n140, u2_u10_u5_n141, u2_u10_u5_n142, u2_u10_u5_n143, u2_u10_u5_n144, u2_u10_u5_n145, 
       u2_u10_u5_n146, u2_u10_u5_n147, u2_u10_u5_n148, u2_u10_u5_n149, u2_u10_u5_n150, u2_u10_u5_n151, u2_u10_u5_n152, u2_u10_u5_n153, u2_u10_u5_n154, 
       u2_u10_u5_n155, u2_u10_u5_n156, u2_u10_u5_n157, u2_u10_u5_n158, u2_u10_u5_n159, u2_u10_u5_n160, u2_u10_u5_n161, u2_u10_u5_n162, u2_u10_u5_n163, 
       u2_u10_u5_n164, u2_u10_u5_n165, u2_u10_u5_n166, u2_u10_u5_n167, u2_u10_u5_n168, u2_u10_u5_n169, u2_u10_u5_n170, u2_u10_u5_n171, u2_u10_u5_n172, 
       u2_u10_u5_n173, u2_u10_u5_n174, u2_u10_u5_n175, u2_u10_u5_n176, u2_u10_u5_n177, u2_u10_u5_n178, u2_u10_u5_n179, u2_u10_u5_n180, u2_u10_u5_n181, 
       u2_u10_u5_n182, u2_u10_u5_n183, u2_u10_u5_n184, u2_u10_u5_n185, u2_u10_u5_n186, u2_u10_u5_n187, u2_u10_u5_n188, u2_u10_u5_n189, u2_u10_u5_n190, 
       u2_u10_u5_n191, u2_u10_u5_n192, u2_u10_u5_n193, u2_u10_u5_n194, u2_u10_u5_n195, u2_u10_u5_n196, u2_u10_u5_n99, u2_u10_u6_n100, u2_u10_u6_n101, 
       u2_u10_u6_n102, u2_u10_u6_n103, u2_u10_u6_n104, u2_u10_u6_n105, u2_u10_u6_n106, u2_u10_u6_n107, u2_u10_u6_n108, u2_u10_u6_n109, u2_u10_u6_n110, 
       u2_u10_u6_n111, u2_u10_u6_n112, u2_u10_u6_n113, u2_u10_u6_n114, u2_u10_u6_n115, u2_u10_u6_n116, u2_u10_u6_n117, u2_u10_u6_n118, u2_u10_u6_n119, 
       u2_u10_u6_n120, u2_u10_u6_n121, u2_u10_u6_n122, u2_u10_u6_n123, u2_u10_u6_n124, u2_u10_u6_n125, u2_u10_u6_n126, u2_u10_u6_n127, u2_u10_u6_n128, 
       u2_u10_u6_n129, u2_u10_u6_n130, u2_u10_u6_n131, u2_u10_u6_n132, u2_u10_u6_n133, u2_u10_u6_n134, u2_u10_u6_n135, u2_u10_u6_n136, u2_u10_u6_n137, 
       u2_u10_u6_n138, u2_u10_u6_n139, u2_u10_u6_n140, u2_u10_u6_n141, u2_u10_u6_n142, u2_u10_u6_n143, u2_u10_u6_n144, u2_u10_u6_n145, u2_u10_u6_n146, 
       u2_u10_u6_n147, u2_u10_u6_n148, u2_u10_u6_n149, u2_u10_u6_n150, u2_u10_u6_n151, u2_u10_u6_n152, u2_u10_u6_n153, u2_u10_u6_n154, u2_u10_u6_n155, 
       u2_u10_u6_n156, u2_u10_u6_n157, u2_u10_u6_n158, u2_u10_u6_n159, u2_u10_u6_n160, u2_u10_u6_n161, u2_u10_u6_n162, u2_u10_u6_n163, u2_u10_u6_n164, 
       u2_u10_u6_n165, u2_u10_u6_n166, u2_u10_u6_n167, u2_u10_u6_n168, u2_u10_u6_n169, u2_u10_u6_n170, u2_u10_u6_n171, u2_u10_u6_n172, u2_u10_u6_n173, 
       u2_u10_u6_n174, u2_u10_u6_n88, u2_u10_u6_n89, u2_u10_u6_n90, u2_u10_u6_n91, u2_u10_u6_n92, u2_u10_u6_n93, u2_u10_u6_n94, u2_u10_u6_n95, 
       u2_u10_u6_n96, u2_u10_u6_n97, u2_u10_u6_n98, u2_u10_u6_n99, u2_u10_u7_n100, u2_u10_u7_n101, u2_u10_u7_n102, u2_u10_u7_n103, u2_u10_u7_n104, 
       u2_u10_u7_n105, u2_u10_u7_n106, u2_u10_u7_n107, u2_u10_u7_n108, u2_u10_u7_n109, u2_u10_u7_n110, u2_u10_u7_n111, u2_u10_u7_n112, u2_u10_u7_n113, 
       u2_u10_u7_n114, u2_u10_u7_n115, u2_u10_u7_n116, u2_u10_u7_n117, u2_u10_u7_n118, u2_u10_u7_n119, u2_u10_u7_n120, u2_u10_u7_n121, u2_u10_u7_n122, 
       u2_u10_u7_n123, u2_u10_u7_n124, u2_u10_u7_n125, u2_u10_u7_n126, u2_u10_u7_n127, u2_u10_u7_n128, u2_u10_u7_n129, u2_u10_u7_n130, u2_u10_u7_n131, 
       u2_u10_u7_n132, u2_u10_u7_n133, u2_u10_u7_n134, u2_u10_u7_n135, u2_u10_u7_n136, u2_u10_u7_n137, u2_u10_u7_n138, u2_u10_u7_n139, u2_u10_u7_n140, 
       u2_u10_u7_n141, u2_u10_u7_n142, u2_u10_u7_n143, u2_u10_u7_n144, u2_u10_u7_n145, u2_u10_u7_n146, u2_u10_u7_n147, u2_u10_u7_n148, u2_u10_u7_n149, 
       u2_u10_u7_n150, u2_u10_u7_n151, u2_u10_u7_n152, u2_u10_u7_n153, u2_u10_u7_n154, u2_u10_u7_n155, u2_u10_u7_n156, u2_u10_u7_n157, u2_u10_u7_n158, 
       u2_u10_u7_n159, u2_u10_u7_n160, u2_u10_u7_n161, u2_u10_u7_n162, u2_u10_u7_n163, u2_u10_u7_n164, u2_u10_u7_n165, u2_u10_u7_n166, u2_u10_u7_n167, 
       u2_u10_u7_n168, u2_u10_u7_n169, u2_u10_u7_n170, u2_u10_u7_n171, u2_u10_u7_n172, u2_u10_u7_n173, u2_u10_u7_n174, u2_u10_u7_n175, u2_u10_u7_n176, 
       u2_u10_u7_n177, u2_u10_u7_n178, u2_u10_u7_n179, u2_u10_u7_n180, u2_u10_u7_n91, u2_u10_u7_n92, u2_u10_u7_n93, u2_u10_u7_n94, u2_u10_u7_n95, 
       u2_u10_u7_n96, u2_u10_u7_n97, u2_u10_u7_n98, u2_u10_u7_n99, u2_u11_X_1, u2_u11_X_10, u2_u11_X_11, u2_u11_X_12, u2_u11_X_13, 
       u2_u11_X_14, u2_u11_X_17, u2_u11_X_18, u2_u11_X_19, u2_u11_X_2, u2_u11_X_20, u2_u11_X_23, u2_u11_X_25, u2_u11_X_30, 
       u2_u11_X_32, u2_u11_X_36, u2_u11_X_38, u2_u11_X_4, u2_u11_X_42, u2_u11_X_44, u2_u11_X_47, u2_u11_X_48, u2_u11_X_5, 
       u2_u11_X_7, u2_u11_u0_n100, u2_u11_u0_n101, u2_u11_u0_n102, u2_u11_u0_n103, u2_u11_u0_n104, u2_u11_u0_n105, u2_u11_u0_n106, u2_u11_u0_n107, 
       u2_u11_u0_n108, u2_u11_u0_n109, u2_u11_u0_n110, u2_u11_u0_n111, u2_u11_u0_n112, u2_u11_u0_n113, u2_u11_u0_n114, u2_u11_u0_n115, u2_u11_u0_n116, 
       u2_u11_u0_n117, u2_u11_u0_n118, u2_u11_u0_n119, u2_u11_u0_n120, u2_u11_u0_n121, u2_u11_u0_n122, u2_u11_u0_n123, u2_u11_u0_n124, u2_u11_u0_n125, 
       u2_u11_u0_n126, u2_u11_u0_n127, u2_u11_u0_n128, u2_u11_u0_n129, u2_u11_u0_n130, u2_u11_u0_n131, u2_u11_u0_n132, u2_u11_u0_n133, u2_u11_u0_n134, 
       u2_u11_u0_n135, u2_u11_u0_n136, u2_u11_u0_n137, u2_u11_u0_n138, u2_u11_u0_n139, u2_u11_u0_n140, u2_u11_u0_n141, u2_u11_u0_n142, u2_u11_u0_n143, 
       u2_u11_u0_n144, u2_u11_u0_n145, u2_u11_u0_n146, u2_u11_u0_n147, u2_u11_u0_n148, u2_u11_u0_n149, u2_u11_u0_n150, u2_u11_u0_n151, u2_u11_u0_n152, 
       u2_u11_u0_n153, u2_u11_u0_n154, u2_u11_u0_n155, u2_u11_u0_n156, u2_u11_u0_n157, u2_u11_u0_n158, u2_u11_u0_n159, u2_u11_u0_n160, u2_u11_u0_n161, 
       u2_u11_u0_n162, u2_u11_u0_n163, u2_u11_u0_n164, u2_u11_u0_n165, u2_u11_u0_n166, u2_u11_u0_n167, u2_u11_u0_n168, u2_u11_u0_n169, u2_u11_u0_n170, 
       u2_u11_u0_n171, u2_u11_u0_n172, u2_u11_u0_n173, u2_u11_u0_n174, u2_u11_u0_n88, u2_u11_u0_n89, u2_u11_u0_n90, u2_u11_u0_n91, u2_u11_u0_n92, 
       u2_u11_u0_n93, u2_u11_u0_n94, u2_u11_u0_n95, u2_u11_u0_n96, u2_u11_u0_n97, u2_u11_u0_n98, u2_u11_u0_n99, u2_u11_u1_n100, u2_u11_u1_n101, 
       u2_u11_u1_n102, u2_u11_u1_n103, u2_u11_u1_n104, u2_u11_u1_n105, u2_u11_u1_n106, u2_u11_u1_n107, u2_u11_u1_n108, u2_u11_u1_n109, u2_u11_u1_n110, 
       u2_u11_u1_n111, u2_u11_u1_n112, u2_u11_u1_n113, u2_u11_u1_n114, u2_u11_u1_n115, u2_u11_u1_n116, u2_u11_u1_n117, u2_u11_u1_n118, u2_u11_u1_n119, 
       u2_u11_u1_n120, u2_u11_u1_n121, u2_u11_u1_n122, u2_u11_u1_n123, u2_u11_u1_n124, u2_u11_u1_n125, u2_u11_u1_n126, u2_u11_u1_n127, u2_u11_u1_n128, 
       u2_u11_u1_n129, u2_u11_u1_n130, u2_u11_u1_n131, u2_u11_u1_n132, u2_u11_u1_n133, u2_u11_u1_n134, u2_u11_u1_n135, u2_u11_u1_n136, u2_u11_u1_n137, 
       u2_u11_u1_n138, u2_u11_u1_n139, u2_u11_u1_n140, u2_u11_u1_n141, u2_u11_u1_n142, u2_u11_u1_n143, u2_u11_u1_n144, u2_u11_u1_n145, u2_u11_u1_n146, 
       u2_u11_u1_n147, u2_u11_u1_n148, u2_u11_u1_n149, u2_u11_u1_n150, u2_u11_u1_n151, u2_u11_u1_n152, u2_u11_u1_n153, u2_u11_u1_n154, u2_u11_u1_n155, 
       u2_u11_u1_n156, u2_u11_u1_n157, u2_u11_u1_n158, u2_u11_u1_n159, u2_u11_u1_n160, u2_u11_u1_n161, u2_u11_u1_n162, u2_u11_u1_n163, u2_u11_u1_n164, 
       u2_u11_u1_n165, u2_u11_u1_n166, u2_u11_u1_n167, u2_u11_u1_n168, u2_u11_u1_n169, u2_u11_u1_n170, u2_u11_u1_n171, u2_u11_u1_n172, u2_u11_u1_n173, 
       u2_u11_u1_n174, u2_u11_u1_n175, u2_u11_u1_n176, u2_u11_u1_n177, u2_u11_u1_n178, u2_u11_u1_n179, u2_u11_u1_n180, u2_u11_u1_n181, u2_u11_u1_n182, 
       u2_u11_u1_n183, u2_u11_u1_n184, u2_u11_u1_n185, u2_u11_u1_n186, u2_u11_u1_n187, u2_u11_u1_n188, u2_u11_u1_n95, u2_u11_u1_n96, u2_u11_u1_n97, 
       u2_u11_u1_n98, u2_u11_u1_n99, u2_u11_u2_n100, u2_u11_u2_n101, u2_u11_u2_n102, u2_u11_u2_n103, u2_u11_u2_n104, u2_u11_u2_n105, u2_u11_u2_n106, 
       u2_u11_u2_n107, u2_u11_u2_n108, u2_u11_u2_n109, u2_u11_u2_n110, u2_u11_u2_n111, u2_u11_u2_n112, u2_u11_u2_n113, u2_u11_u2_n114, u2_u11_u2_n115, 
       u2_u11_u2_n116, u2_u11_u2_n117, u2_u11_u2_n118, u2_u11_u2_n119, u2_u11_u2_n120, u2_u11_u2_n121, u2_u11_u2_n122, u2_u11_u2_n123, u2_u11_u2_n124, 
       u2_u11_u2_n125, u2_u11_u2_n126, u2_u11_u2_n127, u2_u11_u2_n128, u2_u11_u2_n129, u2_u11_u2_n130, u2_u11_u2_n131, u2_u11_u2_n132, u2_u11_u2_n133, 
       u2_u11_u2_n134, u2_u11_u2_n135, u2_u11_u2_n136, u2_u11_u2_n137, u2_u11_u2_n138, u2_u11_u2_n139, u2_u11_u2_n140, u2_u11_u2_n141, u2_u11_u2_n142, 
       u2_u11_u2_n143, u2_u11_u2_n144, u2_u11_u2_n145, u2_u11_u2_n146, u2_u11_u2_n147, u2_u11_u2_n148, u2_u11_u2_n149, u2_u11_u2_n150, u2_u11_u2_n151, 
       u2_u11_u2_n152, u2_u11_u2_n153, u2_u11_u2_n154, u2_u11_u2_n155, u2_u11_u2_n156, u2_u11_u2_n157, u2_u11_u2_n158, u2_u11_u2_n159, u2_u11_u2_n160, 
       u2_u11_u2_n161, u2_u11_u2_n162, u2_u11_u2_n163, u2_u11_u2_n164, u2_u11_u2_n165, u2_u11_u2_n166, u2_u11_u2_n167, u2_u11_u2_n168, u2_u11_u2_n169, 
       u2_u11_u2_n170, u2_u11_u2_n171, u2_u11_u2_n172, u2_u11_u2_n173, u2_u11_u2_n174, u2_u11_u2_n175, u2_u11_u2_n176, u2_u11_u2_n177, u2_u11_u2_n178, 
       u2_u11_u2_n179, u2_u11_u2_n180, u2_u11_u2_n181, u2_u11_u2_n182, u2_u11_u2_n183, u2_u11_u2_n184, u2_u11_u2_n185, u2_u11_u2_n186, u2_u11_u2_n187, 
       u2_u11_u2_n188, u2_u11_u2_n95, u2_u11_u2_n96, u2_u11_u2_n97, u2_u11_u2_n98, u2_u11_u2_n99, u2_u11_u3_n100, u2_u11_u3_n101, u2_u11_u3_n102, 
       u2_u11_u3_n103, u2_u11_u3_n104, u2_u11_u3_n105, u2_u11_u3_n106, u2_u11_u3_n107, u2_u11_u3_n108, u2_u11_u3_n109, u2_u11_u3_n110, u2_u11_u3_n111, 
       u2_u11_u3_n112, u2_u11_u3_n113, u2_u11_u3_n114, u2_u11_u3_n115, u2_u11_u3_n116, u2_u11_u3_n117, u2_u11_u3_n118, u2_u11_u3_n119, u2_u11_u3_n120, 
       u2_u11_u3_n121, u2_u11_u3_n122, u2_u11_u3_n123, u2_u11_u3_n124, u2_u11_u3_n125, u2_u11_u3_n126, u2_u11_u3_n127, u2_u11_u3_n128, u2_u11_u3_n129, 
       u2_u11_u3_n130, u2_u11_u3_n131, u2_u11_u3_n132, u2_u11_u3_n133, u2_u11_u3_n134, u2_u11_u3_n135, u2_u11_u3_n136, u2_u11_u3_n137, u2_u11_u3_n138, 
       u2_u11_u3_n139, u2_u11_u3_n140, u2_u11_u3_n141, u2_u11_u3_n142, u2_u11_u3_n143, u2_u11_u3_n144, u2_u11_u3_n145, u2_u11_u3_n146, u2_u11_u3_n147, 
       u2_u11_u3_n148, u2_u11_u3_n149, u2_u11_u3_n150, u2_u11_u3_n151, u2_u11_u3_n152, u2_u11_u3_n153, u2_u11_u3_n154, u2_u11_u3_n155, u2_u11_u3_n156, 
       u2_u11_u3_n157, u2_u11_u3_n158, u2_u11_u3_n159, u2_u11_u3_n160, u2_u11_u3_n161, u2_u11_u3_n162, u2_u11_u3_n163, u2_u11_u3_n164, u2_u11_u3_n165, 
       u2_u11_u3_n166, u2_u11_u3_n167, u2_u11_u3_n168, u2_u11_u3_n169, u2_u11_u3_n170, u2_u11_u3_n171, u2_u11_u3_n172, u2_u11_u3_n173, u2_u11_u3_n174, 
       u2_u11_u3_n175, u2_u11_u3_n176, u2_u11_u3_n177, u2_u11_u3_n178, u2_u11_u3_n179, u2_u11_u3_n180, u2_u11_u3_n181, u2_u11_u3_n182, u2_u11_u3_n183, 
       u2_u11_u3_n184, u2_u11_u3_n185, u2_u11_u3_n186, u2_u11_u3_n94, u2_u11_u3_n95, u2_u11_u3_n96, u2_u11_u3_n97, u2_u11_u3_n98, u2_u11_u3_n99, 
       u2_u11_u4_n100, u2_u11_u4_n101, u2_u11_u4_n102, u2_u11_u4_n103, u2_u11_u4_n104, u2_u11_u4_n105, u2_u11_u4_n106, u2_u11_u4_n107, u2_u11_u4_n108, 
       u2_u11_u4_n109, u2_u11_u4_n110, u2_u11_u4_n111, u2_u11_u4_n112, u2_u11_u4_n113, u2_u11_u4_n114, u2_u11_u4_n115, u2_u11_u4_n116, u2_u11_u4_n117, 
       u2_u11_u4_n118, u2_u11_u4_n119, u2_u11_u4_n120, u2_u11_u4_n121, u2_u11_u4_n122, u2_u11_u4_n123, u2_u11_u4_n124, u2_u11_u4_n125, u2_u11_u4_n126, 
       u2_u11_u4_n127, u2_u11_u4_n128, u2_u11_u4_n129, u2_u11_u4_n130, u2_u11_u4_n131, u2_u11_u4_n132, u2_u11_u4_n133, u2_u11_u4_n134, u2_u11_u4_n135, 
       u2_u11_u4_n136, u2_u11_u4_n137, u2_u11_u4_n138, u2_u11_u4_n139, u2_u11_u4_n140, u2_u11_u4_n141, u2_u11_u4_n142, u2_u11_u4_n143, u2_u11_u4_n144, 
       u2_u11_u4_n145, u2_u11_u4_n146, u2_u11_u4_n147, u2_u11_u4_n148, u2_u11_u4_n149, u2_u11_u4_n150, u2_u11_u4_n151, u2_u11_u4_n152, u2_u11_u4_n153, 
       u2_u11_u4_n154, u2_u11_u4_n155, u2_u11_u4_n156, u2_u11_u4_n157, u2_u11_u4_n158, u2_u11_u4_n159, u2_u11_u4_n160, u2_u11_u4_n161, u2_u11_u4_n162, 
       u2_u11_u4_n163, u2_u11_u4_n164, u2_u11_u4_n165, u2_u11_u4_n166, u2_u11_u4_n167, u2_u11_u4_n168, u2_u11_u4_n169, u2_u11_u4_n170, u2_u11_u4_n171, 
       u2_u11_u4_n172, u2_u11_u4_n173, u2_u11_u4_n174, u2_u11_u4_n175, u2_u11_u4_n176, u2_u11_u4_n177, u2_u11_u4_n178, u2_u11_u4_n179, u2_u11_u4_n180, 
       u2_u11_u4_n181, u2_u11_u4_n182, u2_u11_u4_n183, u2_u11_u4_n184, u2_u11_u4_n185, u2_u11_u4_n186, u2_u11_u4_n94, u2_u11_u4_n95, u2_u11_u4_n96, 
       u2_u11_u4_n97, u2_u11_u4_n98, u2_u11_u4_n99, u2_u11_u5_n100, u2_u11_u5_n101, u2_u11_u5_n102, u2_u11_u5_n103, u2_u11_u5_n104, u2_u11_u5_n105, 
       u2_u11_u5_n106, u2_u11_u5_n107, u2_u11_u5_n108, u2_u11_u5_n109, u2_u11_u5_n110, u2_u11_u5_n111, u2_u11_u5_n112, u2_u11_u5_n113, u2_u11_u5_n114, 
       u2_u11_u5_n115, u2_u11_u5_n116, u2_u11_u5_n117, u2_u11_u5_n118, u2_u11_u5_n119, u2_u11_u5_n120, u2_u11_u5_n121, u2_u11_u5_n122, u2_u11_u5_n123, 
       u2_u11_u5_n124, u2_u11_u5_n125, u2_u11_u5_n126, u2_u11_u5_n127, u2_u11_u5_n128, u2_u11_u5_n129, u2_u11_u5_n130, u2_u11_u5_n131, u2_u11_u5_n132, 
       u2_u11_u5_n133, u2_u11_u5_n134, u2_u11_u5_n135, u2_u11_u5_n136, u2_u11_u5_n137, u2_u11_u5_n138, u2_u11_u5_n139, u2_u11_u5_n140, u2_u11_u5_n141, 
       u2_u11_u5_n142, u2_u11_u5_n143, u2_u11_u5_n144, u2_u11_u5_n145, u2_u11_u5_n146, u2_u11_u5_n147, u2_u11_u5_n148, u2_u11_u5_n149, u2_u11_u5_n150, 
       u2_u11_u5_n151, u2_u11_u5_n152, u2_u11_u5_n153, u2_u11_u5_n154, u2_u11_u5_n155, u2_u11_u5_n156, u2_u11_u5_n157, u2_u11_u5_n158, u2_u11_u5_n159, 
       u2_u11_u5_n160, u2_u11_u5_n161, u2_u11_u5_n162, u2_u11_u5_n163, u2_u11_u5_n164, u2_u11_u5_n165, u2_u11_u5_n166, u2_u11_u5_n167, u2_u11_u5_n168, 
       u2_u11_u5_n169, u2_u11_u5_n170, u2_u11_u5_n171, u2_u11_u5_n172, u2_u11_u5_n173, u2_u11_u5_n174, u2_u11_u5_n175, u2_u11_u5_n176, u2_u11_u5_n177, 
       u2_u11_u5_n178, u2_u11_u5_n179, u2_u11_u5_n180, u2_u11_u5_n181, u2_u11_u5_n182, u2_u11_u5_n183, u2_u11_u5_n184, u2_u11_u5_n185, u2_u11_u5_n186, 
       u2_u11_u5_n187, u2_u11_u5_n188, u2_u11_u5_n189, u2_u11_u5_n190, u2_u11_u5_n191, u2_u11_u5_n192, u2_u11_u5_n193, u2_u11_u5_n194, u2_u11_u5_n195, 
       u2_u11_u5_n196, u2_u11_u5_n99, u2_u11_u6_n100, u2_u11_u6_n101, u2_u11_u6_n102, u2_u11_u6_n103, u2_u11_u6_n104, u2_u11_u6_n105, u2_u11_u6_n106, 
       u2_u11_u6_n107, u2_u11_u6_n108, u2_u11_u6_n109, u2_u11_u6_n110, u2_u11_u6_n111, u2_u11_u6_n112, u2_u11_u6_n113, u2_u11_u6_n114, u2_u11_u6_n115, 
       u2_u11_u6_n116, u2_u11_u6_n117, u2_u11_u6_n118, u2_u11_u6_n119, u2_u11_u6_n120, u2_u11_u6_n121, u2_u11_u6_n122, u2_u11_u6_n123, u2_u11_u6_n124, 
       u2_u11_u6_n125, u2_u11_u6_n126, u2_u11_u6_n127, u2_u11_u6_n128, u2_u11_u6_n129, u2_u11_u6_n130, u2_u11_u6_n131, u2_u11_u6_n132, u2_u11_u6_n133, 
       u2_u11_u6_n134, u2_u11_u6_n135, u2_u11_u6_n136, u2_u11_u6_n137, u2_u11_u6_n138, u2_u11_u6_n139, u2_u11_u6_n140, u2_u11_u6_n141, u2_u11_u6_n142, 
       u2_u11_u6_n143, u2_u11_u6_n144, u2_u11_u6_n145, u2_u11_u6_n146, u2_u11_u6_n147, u2_u11_u6_n148, u2_u11_u6_n149, u2_u11_u6_n150, u2_u11_u6_n151, 
       u2_u11_u6_n152, u2_u11_u6_n153, u2_u11_u6_n154, u2_u11_u6_n155, u2_u11_u6_n156, u2_u11_u6_n157, u2_u11_u6_n158, u2_u11_u6_n159, u2_u11_u6_n160, 
       u2_u11_u6_n161, u2_u11_u6_n162, u2_u11_u6_n163, u2_u11_u6_n164, u2_u11_u6_n165, u2_u11_u6_n166, u2_u11_u6_n167, u2_u11_u6_n168, u2_u11_u6_n169, 
       u2_u11_u6_n170, u2_u11_u6_n171, u2_u11_u6_n172, u2_u11_u6_n173, u2_u11_u6_n174, u2_u11_u6_n88, u2_u11_u6_n89, u2_u11_u6_n90, u2_u11_u6_n91, 
       u2_u11_u6_n92, u2_u11_u6_n93, u2_u11_u6_n94, u2_u11_u6_n95, u2_u11_u6_n96, u2_u11_u6_n97, u2_u11_u6_n98, u2_u11_u6_n99, u2_u11_u7_n100, 
       u2_u11_u7_n101, u2_u11_u7_n102, u2_u11_u7_n103, u2_u11_u7_n104, u2_u11_u7_n105, u2_u11_u7_n106, u2_u11_u7_n107, u2_u11_u7_n108, u2_u11_u7_n109, 
       u2_u11_u7_n110, u2_u11_u7_n111, u2_u11_u7_n112, u2_u11_u7_n113, u2_u11_u7_n114, u2_u11_u7_n115, u2_u11_u7_n116, u2_u11_u7_n117, u2_u11_u7_n118, 
       u2_u11_u7_n119, u2_u11_u7_n120, u2_u11_u7_n121, u2_u11_u7_n122, u2_u11_u7_n123, u2_u11_u7_n124, u2_u11_u7_n125, u2_u11_u7_n126, u2_u11_u7_n127, 
       u2_u11_u7_n128, u2_u11_u7_n129, u2_u11_u7_n130, u2_u11_u7_n131, u2_u11_u7_n132, u2_u11_u7_n133, u2_u11_u7_n134, u2_u11_u7_n135, u2_u11_u7_n136, 
       u2_u11_u7_n137, u2_u11_u7_n138, u2_u11_u7_n139, u2_u11_u7_n140, u2_u11_u7_n141, u2_u11_u7_n142, u2_u11_u7_n143, u2_u11_u7_n144, u2_u11_u7_n145, 
       u2_u11_u7_n146, u2_u11_u7_n147, u2_u11_u7_n148, u2_u11_u7_n149, u2_u11_u7_n150, u2_u11_u7_n151, u2_u11_u7_n152, u2_u11_u7_n153, u2_u11_u7_n154, 
       u2_u11_u7_n155, u2_u11_u7_n156, u2_u11_u7_n157, u2_u11_u7_n158, u2_u11_u7_n159, u2_u11_u7_n160, u2_u11_u7_n161, u2_u11_u7_n162, u2_u11_u7_n163, 
       u2_u11_u7_n164, u2_u11_u7_n165, u2_u11_u7_n166, u2_u11_u7_n167, u2_u11_u7_n168, u2_u11_u7_n169, u2_u11_u7_n170, u2_u11_u7_n171, u2_u11_u7_n172, 
       u2_u11_u7_n173, u2_u11_u7_n174, u2_u11_u7_n175, u2_u11_u7_n176, u2_u11_u7_n177, u2_u11_u7_n178, u2_u11_u7_n179, u2_u11_u7_n180, u2_u11_u7_n91, 
       u2_u11_u7_n92, u2_u11_u7_n93, u2_u11_u7_n94, u2_u11_u7_n95, u2_u11_u7_n96, u2_u11_u7_n97, u2_u11_u7_n98, u2_u11_u7_n99, u2_u12_X_2, 
       u2_u12_X_30, u2_u12_X_32, u2_u12_X_35, u2_u12_X_37, u2_u12_X_48, u2_u12_X_5, u2_u12_X_7, u2_u12_u0_n100, u2_u12_u0_n101, 
       u2_u12_u0_n102, u2_u12_u0_n103, u2_u12_u0_n104, u2_u12_u0_n105, u2_u12_u0_n106, u2_u12_u0_n107, u2_u12_u0_n108, u2_u12_u0_n109, u2_u12_u0_n110, 
       u2_u12_u0_n111, u2_u12_u0_n112, u2_u12_u0_n113, u2_u12_u0_n114, u2_u12_u0_n115, u2_u12_u0_n116, u2_u12_u0_n117, u2_u12_u0_n118, u2_u12_u0_n119, 
       u2_u12_u0_n120, u2_u12_u0_n121, u2_u12_u0_n122, u2_u12_u0_n123, u2_u12_u0_n124, u2_u12_u0_n125, u2_u12_u0_n126, u2_u12_u0_n127, u2_u12_u0_n128, 
       u2_u12_u0_n129, u2_u12_u0_n130, u2_u12_u0_n131, u2_u12_u0_n132, u2_u12_u0_n133, u2_u12_u0_n134, u2_u12_u0_n135, u2_u12_u0_n136, u2_u12_u0_n137, 
       u2_u12_u0_n138, u2_u12_u0_n139, u2_u12_u0_n140, u2_u12_u0_n141, u2_u12_u0_n142, u2_u12_u0_n143, u2_u12_u0_n144, u2_u12_u0_n145, u2_u12_u0_n146, 
       u2_u12_u0_n147, u2_u12_u0_n148, u2_u12_u0_n149, u2_u12_u0_n150, u2_u12_u0_n151, u2_u12_u0_n152, u2_u12_u0_n153, u2_u12_u0_n154, u2_u12_u0_n155, 
       u2_u12_u0_n156, u2_u12_u0_n157, u2_u12_u0_n158, u2_u12_u0_n159, u2_u12_u0_n160, u2_u12_u0_n161, u2_u12_u0_n162, u2_u12_u0_n163, u2_u12_u0_n164, 
       u2_u12_u0_n165, u2_u12_u0_n166, u2_u12_u0_n167, u2_u12_u0_n168, u2_u12_u0_n169, u2_u12_u0_n170, u2_u12_u0_n171, u2_u12_u0_n172, u2_u12_u0_n173, 
       u2_u12_u0_n174, u2_u12_u0_n88, u2_u12_u0_n89, u2_u12_u0_n90, u2_u12_u0_n91, u2_u12_u0_n92, u2_u12_u0_n93, u2_u12_u0_n94, u2_u12_u0_n95, 
       u2_u12_u0_n96, u2_u12_u0_n97, u2_u12_u0_n98, u2_u12_u0_n99, u2_u12_u1_n100, u2_u12_u1_n101, u2_u12_u1_n102, u2_u12_u1_n103, u2_u12_u1_n104, 
       u2_u12_u1_n105, u2_u12_u1_n106, u2_u12_u1_n107, u2_u12_u1_n108, u2_u12_u1_n109, u2_u12_u1_n110, u2_u12_u1_n111, u2_u12_u1_n112, u2_u12_u1_n113, 
       u2_u12_u1_n114, u2_u12_u1_n115, u2_u12_u1_n116, u2_u12_u1_n117, u2_u12_u1_n118, u2_u12_u1_n119, u2_u12_u1_n120, u2_u12_u1_n121, u2_u12_u1_n122, 
       u2_u12_u1_n123, u2_u12_u1_n124, u2_u12_u1_n125, u2_u12_u1_n126, u2_u12_u1_n127, u2_u12_u1_n128, u2_u12_u1_n129, u2_u12_u1_n130, u2_u12_u1_n131, 
       u2_u12_u1_n132, u2_u12_u1_n133, u2_u12_u1_n134, u2_u12_u1_n135, u2_u12_u1_n136, u2_u12_u1_n137, u2_u12_u1_n138, u2_u12_u1_n139, u2_u12_u1_n140, 
       u2_u12_u1_n141, u2_u12_u1_n142, u2_u12_u1_n143, u2_u12_u1_n144, u2_u12_u1_n145, u2_u12_u1_n146, u2_u12_u1_n147, u2_u12_u1_n148, u2_u12_u1_n149, 
       u2_u12_u1_n150, u2_u12_u1_n151, u2_u12_u1_n152, u2_u12_u1_n153, u2_u12_u1_n154, u2_u12_u1_n155, u2_u12_u1_n156, u2_u12_u1_n157, u2_u12_u1_n158, 
       u2_u12_u1_n159, u2_u12_u1_n160, u2_u12_u1_n161, u2_u12_u1_n162, u2_u12_u1_n163, u2_u12_u1_n164, u2_u12_u1_n165, u2_u12_u1_n166, u2_u12_u1_n167, 
       u2_u12_u1_n168, u2_u12_u1_n169, u2_u12_u1_n170, u2_u12_u1_n171, u2_u12_u1_n172, u2_u12_u1_n173, u2_u12_u1_n174, u2_u12_u1_n175, u2_u12_u1_n176, 
       u2_u12_u1_n177, u2_u12_u1_n178, u2_u12_u1_n179, u2_u12_u1_n180, u2_u12_u1_n181, u2_u12_u1_n182, u2_u12_u1_n183, u2_u12_u1_n184, u2_u12_u1_n185, 
       u2_u12_u1_n186, u2_u12_u1_n187, u2_u12_u1_n188, u2_u12_u1_n95, u2_u12_u1_n96, u2_u12_u1_n97, u2_u12_u1_n98, u2_u12_u1_n99, u2_u12_u4_n100, 
       u2_u12_u4_n101, u2_u12_u4_n102, u2_u12_u4_n103, u2_u12_u4_n104, u2_u12_u4_n105, u2_u12_u4_n106, u2_u12_u4_n107, u2_u12_u4_n108, u2_u12_u4_n109, 
       u2_u12_u4_n110, u2_u12_u4_n111, u2_u12_u4_n112, u2_u12_u4_n113, u2_u12_u4_n114, u2_u12_u4_n115, u2_u12_u4_n116, u2_u12_u4_n117, u2_u12_u4_n118, 
       u2_u12_u4_n119, u2_u12_u4_n120, u2_u12_u4_n121, u2_u12_u4_n122, u2_u12_u4_n123, u2_u12_u4_n124, u2_u12_u4_n125, u2_u12_u4_n126, u2_u12_u4_n127, 
       u2_u12_u4_n128, u2_u12_u4_n129, u2_u12_u4_n130, u2_u12_u4_n131, u2_u12_u4_n132, u2_u12_u4_n133, u2_u12_u4_n134, u2_u12_u4_n135, u2_u12_u4_n136, 
       u2_u12_u4_n137, u2_u12_u4_n138, u2_u12_u4_n139, u2_u12_u4_n140, u2_u12_u4_n141, u2_u12_u4_n142, u2_u12_u4_n143, u2_u12_u4_n144, u2_u12_u4_n145, 
       u2_u12_u4_n146, u2_u12_u4_n147, u2_u12_u4_n148, u2_u12_u4_n149, u2_u12_u4_n150, u2_u12_u4_n151, u2_u12_u4_n152, u2_u12_u4_n153, u2_u12_u4_n154, 
       u2_u12_u4_n155, u2_u12_u4_n156, u2_u12_u4_n157, u2_u12_u4_n158, u2_u12_u4_n159, u2_u12_u4_n160, u2_u12_u4_n161, u2_u12_u4_n162, u2_u12_u4_n163, 
       u2_u12_u4_n164, u2_u12_u4_n165, u2_u12_u4_n166, u2_u12_u4_n167, u2_u12_u4_n168, u2_u12_u4_n169, u2_u12_u4_n170, u2_u12_u4_n171, u2_u12_u4_n172, 
       u2_u12_u4_n173, u2_u12_u4_n174, u2_u12_u4_n175, u2_u12_u4_n176, u2_u12_u4_n177, u2_u12_u4_n178, u2_u12_u4_n179, u2_u12_u4_n180, u2_u12_u4_n181, 
       u2_u12_u4_n182, u2_u12_u4_n183, u2_u12_u4_n184, u2_u12_u4_n185, u2_u12_u4_n186, u2_u12_u4_n94, u2_u12_u4_n95, u2_u12_u4_n96, u2_u12_u4_n97, 
       u2_u12_u4_n98, u2_u12_u4_n99, u2_u12_u5_n100, u2_u12_u5_n101, u2_u12_u5_n102, u2_u12_u5_n103, u2_u12_u5_n104, u2_u12_u5_n105, u2_u12_u5_n106, 
       u2_u12_u5_n107, u2_u12_u5_n108, u2_u12_u5_n109, u2_u12_u5_n110, u2_u12_u5_n111, u2_u12_u5_n112, u2_u12_u5_n113, u2_u12_u5_n114, u2_u12_u5_n115, 
       u2_u12_u5_n116, u2_u12_u5_n117, u2_u12_u5_n118, u2_u12_u5_n119, u2_u12_u5_n120, u2_u12_u5_n121, u2_u12_u5_n122, u2_u12_u5_n123, u2_u12_u5_n124, 
       u2_u12_u5_n125, u2_u12_u5_n126, u2_u12_u5_n127, u2_u12_u5_n128, u2_u12_u5_n129, u2_u12_u5_n130, u2_u12_u5_n131, u2_u12_u5_n132, u2_u12_u5_n133, 
       u2_u12_u5_n134, u2_u12_u5_n135, u2_u12_u5_n136, u2_u12_u5_n137, u2_u12_u5_n138, u2_u12_u5_n139, u2_u12_u5_n140, u2_u12_u5_n141, u2_u12_u5_n142, 
       u2_u12_u5_n143, u2_u12_u5_n144, u2_u12_u5_n145, u2_u12_u5_n146, u2_u12_u5_n147, u2_u12_u5_n148, u2_u12_u5_n149, u2_u12_u5_n150, u2_u12_u5_n151, 
       u2_u12_u5_n152, u2_u12_u5_n153, u2_u12_u5_n154, u2_u12_u5_n155, u2_u12_u5_n156, u2_u12_u5_n157, u2_u12_u5_n158, u2_u12_u5_n159, u2_u12_u5_n160, 
       u2_u12_u5_n161, u2_u12_u5_n162, u2_u12_u5_n163, u2_u12_u5_n164, u2_u12_u5_n165, u2_u12_u5_n166, u2_u12_u5_n167, u2_u12_u5_n168, u2_u12_u5_n169, 
       u2_u12_u5_n170, u2_u12_u5_n171, u2_u12_u5_n172, u2_u12_u5_n173, u2_u12_u5_n174, u2_u12_u5_n175, u2_u12_u5_n176, u2_u12_u5_n177, u2_u12_u5_n178, 
       u2_u12_u5_n179, u2_u12_u5_n180, u2_u12_u5_n181, u2_u12_u5_n182, u2_u12_u5_n183, u2_u12_u5_n184, u2_u12_u5_n185, u2_u12_u5_n186, u2_u12_u5_n187, 
       u2_u12_u5_n188, u2_u12_u5_n189, u2_u12_u5_n190, u2_u12_u5_n191, u2_u12_u5_n192, u2_u12_u5_n193, u2_u12_u5_n194, u2_u12_u5_n195, u2_u12_u5_n196, 
       u2_u12_u5_n99, u2_u12_u6_n100, u2_u12_u6_n101, u2_u12_u6_n102, u2_u12_u6_n103, u2_u12_u6_n104, u2_u12_u6_n105, u2_u12_u6_n106, u2_u12_u6_n107, 
       u2_u12_u6_n108, u2_u12_u6_n109, u2_u12_u6_n110, u2_u12_u6_n111, u2_u12_u6_n112, u2_u12_u6_n113, u2_u12_u6_n114, u2_u12_u6_n115, u2_u12_u6_n116, 
       u2_u12_u6_n117, u2_u12_u6_n118, u2_u12_u6_n119, u2_u12_u6_n120, u2_u12_u6_n121, u2_u12_u6_n122, u2_u12_u6_n123, u2_u12_u6_n124, u2_u12_u6_n125, 
       u2_u12_u6_n126, u2_u12_u6_n127, u2_u12_u6_n128, u2_u12_u6_n129, u2_u12_u6_n130, u2_u12_u6_n131, u2_u12_u6_n132, u2_u12_u6_n133, u2_u12_u6_n134, 
       u2_u12_u6_n135, u2_u12_u6_n136, u2_u12_u6_n137, u2_u12_u6_n138, u2_u12_u6_n139, u2_u12_u6_n140, u2_u12_u6_n141, u2_u12_u6_n142, u2_u12_u6_n143, 
       u2_u12_u6_n144, u2_u12_u6_n145, u2_u12_u6_n146, u2_u12_u6_n147, u2_u12_u6_n148, u2_u12_u6_n149, u2_u12_u6_n150, u2_u12_u6_n151, u2_u12_u6_n152, 
       u2_u12_u6_n153, u2_u12_u6_n154, u2_u12_u6_n155, u2_u12_u6_n156, u2_u12_u6_n157, u2_u12_u6_n158, u2_u12_u6_n159, u2_u12_u6_n160, u2_u12_u6_n161, 
       u2_u12_u6_n162, u2_u12_u6_n163, u2_u12_u6_n164, u2_u12_u6_n165, u2_u12_u6_n166, u2_u12_u6_n167, u2_u12_u6_n168, u2_u12_u6_n169, u2_u12_u6_n170, 
       u2_u12_u6_n171, u2_u12_u6_n172, u2_u12_u6_n173, u2_u12_u6_n174, u2_u12_u6_n88, u2_u12_u6_n89, u2_u12_u6_n90, u2_u12_u6_n91, u2_u12_u6_n92, 
       u2_u12_u6_n93, u2_u12_u6_n94, u2_u12_u6_n95, u2_u12_u6_n96, u2_u12_u6_n97, u2_u12_u6_n98, u2_u12_u6_n99, u2_u12_u7_n100, u2_u12_u7_n101, 
       u2_u12_u7_n102, u2_u12_u7_n103, u2_u12_u7_n104, u2_u12_u7_n105, u2_u12_u7_n106, u2_u12_u7_n107, u2_u12_u7_n108, u2_u12_u7_n109, u2_u12_u7_n110, 
       u2_u12_u7_n111, u2_u12_u7_n112, u2_u12_u7_n113, u2_u12_u7_n114, u2_u12_u7_n115, u2_u12_u7_n116, u2_u12_u7_n117, u2_u12_u7_n118, u2_u12_u7_n119, 
       u2_u12_u7_n120, u2_u12_u7_n121, u2_u12_u7_n122, u2_u12_u7_n123, u2_u12_u7_n124, u2_u12_u7_n125, u2_u12_u7_n126, u2_u12_u7_n127, u2_u12_u7_n128, 
       u2_u12_u7_n129, u2_u12_u7_n130, u2_u12_u7_n131, u2_u12_u7_n132, u2_u12_u7_n133, u2_u12_u7_n134, u2_u12_u7_n135, u2_u12_u7_n136, u2_u12_u7_n137, 
       u2_u12_u7_n138, u2_u12_u7_n139, u2_u12_u7_n140, u2_u12_u7_n141, u2_u12_u7_n142, u2_u12_u7_n143, u2_u12_u7_n144, u2_u12_u7_n145, u2_u12_u7_n146, 
       u2_u12_u7_n147, u2_u12_u7_n148, u2_u12_u7_n149, u2_u12_u7_n150, u2_u12_u7_n151, u2_u12_u7_n152, u2_u12_u7_n153, u2_u12_u7_n154, u2_u12_u7_n155, 
       u2_u12_u7_n156, u2_u12_u7_n157, u2_u12_u7_n158, u2_u12_u7_n159, u2_u12_u7_n160, u2_u12_u7_n161, u2_u12_u7_n162, u2_u12_u7_n163, u2_u12_u7_n164, 
       u2_u12_u7_n165, u2_u12_u7_n166, u2_u12_u7_n167, u2_u12_u7_n168, u2_u12_u7_n169, u2_u12_u7_n170, u2_u12_u7_n171, u2_u12_u7_n172, u2_u12_u7_n173, 
       u2_u12_u7_n174, u2_u12_u7_n175, u2_u12_u7_n176, u2_u12_u7_n177, u2_u12_u7_n178, u2_u12_u7_n179, u2_u12_u7_n180, u2_u12_u7_n91, u2_u12_u7_n92, 
       u2_u12_u7_n93, u2_u12_u7_n94, u2_u12_u7_n95, u2_u12_u7_n96, u2_u12_u7_n97, u2_u12_u7_n98, u2_u12_u7_n99, u2_u13_X_29, u2_u13_X_30, 
       u2_u13_X_31, u2_u13_X_32, u2_u13_X_33, u2_u13_X_36, u2_u13_X_38, u2_u13_u4_n100, u2_u13_u4_n101, u2_u13_u4_n102, u2_u13_u4_n103, 
       u2_u13_u4_n104, u2_u13_u4_n105, u2_u13_u4_n106, u2_u13_u4_n107, u2_u13_u4_n108, u2_u13_u4_n109, u2_u13_u4_n110, u2_u13_u4_n111, u2_u13_u4_n112, 
       u2_u13_u4_n113, u2_u13_u4_n114, u2_u13_u4_n115, u2_u13_u4_n116, u2_u13_u4_n117, u2_u13_u4_n118, u2_u13_u4_n119, u2_u13_u4_n120, u2_u13_u4_n121, 
       u2_u13_u4_n122, u2_u13_u4_n123, u2_u13_u4_n124, u2_u13_u4_n125, u2_u13_u4_n126, u2_u13_u4_n127, u2_u13_u4_n128, u2_u13_u4_n129, u2_u13_u4_n130, 
       u2_u13_u4_n131, u2_u13_u4_n132, u2_u13_u4_n133, u2_u13_u4_n134, u2_u13_u4_n135, u2_u13_u4_n136, u2_u13_u4_n137, u2_u13_u4_n138, u2_u13_u4_n139, 
       u2_u13_u4_n140, u2_u13_u4_n141, u2_u13_u4_n142, u2_u13_u4_n143, u2_u13_u4_n144, u2_u13_u4_n145, u2_u13_u4_n146, u2_u13_u4_n147, u2_u13_u4_n148, 
       u2_u13_u4_n149, u2_u13_u4_n150, u2_u13_u4_n151, u2_u13_u4_n152, u2_u13_u4_n153, u2_u13_u4_n154, u2_u13_u4_n155, u2_u13_u4_n156, u2_u13_u4_n157, 
       u2_u13_u4_n158, u2_u13_u4_n159, u2_u13_u4_n160, u2_u13_u4_n161, u2_u13_u4_n162, u2_u13_u4_n163, u2_u13_u4_n164, u2_u13_u4_n165, u2_u13_u4_n166, 
       u2_u13_u4_n167, u2_u13_u4_n168, u2_u13_u4_n169, u2_u13_u4_n170, u2_u13_u4_n171, u2_u13_u4_n172, u2_u13_u4_n173, u2_u13_u4_n174, u2_u13_u4_n175, 
       u2_u13_u4_n176, u2_u13_u4_n177, u2_u13_u4_n178, u2_u13_u4_n179, u2_u13_u4_n180, u2_u13_u4_n181, u2_u13_u4_n182, u2_u13_u4_n183, u2_u13_u4_n184, 
       u2_u13_u4_n185, u2_u13_u4_n186, u2_u13_u4_n94, u2_u13_u4_n95, u2_u13_u4_n96, u2_u13_u4_n97, u2_u13_u4_n98, u2_u13_u4_n99, u2_u13_u5_n100, 
       u2_u13_u5_n101, u2_u13_u5_n102, u2_u13_u5_n103, u2_u13_u5_n104, u2_u13_u5_n105, u2_u13_u5_n106, u2_u13_u5_n107, u2_u13_u5_n108, u2_u13_u5_n109, 
       u2_u13_u5_n110, u2_u13_u5_n111, u2_u13_u5_n112, u2_u13_u5_n113, u2_u13_u5_n114, u2_u13_u5_n115, u2_u13_u5_n116, u2_u13_u5_n117, u2_u13_u5_n118, 
       u2_u13_u5_n119, u2_u13_u5_n120, u2_u13_u5_n121, u2_u13_u5_n122, u2_u13_u5_n123, u2_u13_u5_n124, u2_u13_u5_n125, u2_u13_u5_n126, u2_u13_u5_n127, 
       u2_u13_u5_n128, u2_u13_u5_n129, u2_u13_u5_n130, u2_u13_u5_n131, u2_u13_u5_n132, u2_u13_u5_n133, u2_u13_u5_n134, u2_u13_u5_n135, u2_u13_u5_n136, 
       u2_u13_u5_n137, u2_u13_u5_n138, u2_u13_u5_n139, u2_u13_u5_n140, u2_u13_u5_n141, u2_u13_u5_n142, u2_u13_u5_n143, u2_u13_u5_n144, u2_u13_u5_n145, 
       u2_u13_u5_n146, u2_u13_u5_n147, u2_u13_u5_n148, u2_u13_u5_n149, u2_u13_u5_n150, u2_u13_u5_n151, u2_u13_u5_n152, u2_u13_u5_n153, u2_u13_u5_n154, 
       u2_u13_u5_n155, u2_u13_u5_n156, u2_u13_u5_n157, u2_u13_u5_n158, u2_u13_u5_n159, u2_u13_u5_n160, u2_u13_u5_n161, u2_u13_u5_n162, u2_u13_u5_n163, 
       u2_u13_u5_n164, u2_u13_u5_n165, u2_u13_u5_n166, u2_u13_u5_n167, u2_u13_u5_n168, u2_u13_u5_n169, u2_u13_u5_n170, u2_u13_u5_n171, u2_u13_u5_n172, 
       u2_u13_u5_n173, u2_u13_u5_n174, u2_u13_u5_n175, u2_u13_u5_n176, u2_u13_u5_n177, u2_u13_u5_n178, u2_u13_u5_n179, u2_u13_u5_n180, u2_u13_u5_n181, 
       u2_u13_u5_n182, u2_u13_u5_n183, u2_u13_u5_n184, u2_u13_u5_n185, u2_u13_u5_n186, u2_u13_u5_n187, u2_u13_u5_n188, u2_u13_u5_n189, u2_u13_u5_n190, 
       u2_u13_u5_n191, u2_u13_u5_n192, u2_u13_u5_n193, u2_u13_u5_n194, u2_u13_u5_n195, u2_u13_u5_n196, u2_u13_u5_n99, u2_u13_u6_n100, u2_u13_u6_n101, 
       u2_u13_u6_n102, u2_u13_u6_n103, u2_u13_u6_n104, u2_u13_u6_n105, u2_u13_u6_n106, u2_u13_u6_n107, u2_u13_u6_n108, u2_u13_u6_n109, u2_u13_u6_n110, 
       u2_u13_u6_n111, u2_u13_u6_n112, u2_u13_u6_n113, u2_u13_u6_n114, u2_u13_u6_n115, u2_u13_u6_n116, u2_u13_u6_n117, u2_u13_u6_n118, u2_u13_u6_n119, 
       u2_u13_u6_n120, u2_u13_u6_n121, u2_u13_u6_n122, u2_u13_u6_n123, u2_u13_u6_n124, u2_u13_u6_n125, u2_u13_u6_n126, u2_u13_u6_n127, u2_u13_u6_n128, 
       u2_u13_u6_n129, u2_u13_u6_n130, u2_u13_u6_n131, u2_u13_u6_n132, u2_u13_u6_n133, u2_u13_u6_n134, u2_u13_u6_n135, u2_u13_u6_n136, u2_u13_u6_n137, 
       u2_u13_u6_n138, u2_u13_u6_n139, u2_u13_u6_n140, u2_u13_u6_n141, u2_u13_u6_n142, u2_u13_u6_n143, u2_u13_u6_n144, u2_u13_u6_n145, u2_u13_u6_n146, 
       u2_u13_u6_n147, u2_u13_u6_n148, u2_u13_u6_n149, u2_u13_u6_n150, u2_u13_u6_n151, u2_u13_u6_n152, u2_u13_u6_n153, u2_u13_u6_n154, u2_u13_u6_n155, 
       u2_u13_u6_n156, u2_u13_u6_n157, u2_u13_u6_n158, u2_u13_u6_n159, u2_u13_u6_n160, u2_u13_u6_n161, u2_u13_u6_n162, u2_u13_u6_n163, u2_u13_u6_n164, 
       u2_u13_u6_n165, u2_u13_u6_n166, u2_u13_u6_n167, u2_u13_u6_n168, u2_u13_u6_n169, u2_u13_u6_n170, u2_u13_u6_n171, u2_u13_u6_n172, u2_u13_u6_n173, 
       u2_u13_u6_n174, u2_u13_u6_n88, u2_u13_u6_n89, u2_u13_u6_n90, u2_u13_u6_n91, u2_u13_u6_n92, u2_u13_u6_n93, u2_u13_u6_n94, u2_u13_u6_n95, 
       u2_u13_u6_n96, u2_u13_u6_n97, u2_u13_u6_n98, u2_u13_u6_n99, u2_u13_u7_n100, u2_u13_u7_n101, u2_u13_u7_n102, u2_u13_u7_n103, u2_u13_u7_n104, 
       u2_u13_u7_n105, u2_u13_u7_n106, u2_u13_u7_n107, u2_u13_u7_n108, u2_u13_u7_n109, u2_u13_u7_n110, u2_u13_u7_n111, u2_u13_u7_n112, u2_u13_u7_n113, 
       u2_u13_u7_n114, u2_u13_u7_n115, u2_u13_u7_n116, u2_u13_u7_n117, u2_u13_u7_n118, u2_u13_u7_n119, u2_u13_u7_n120, u2_u13_u7_n121, u2_u13_u7_n122, 
       u2_u13_u7_n123, u2_u13_u7_n124, u2_u13_u7_n125, u2_u13_u7_n126, u2_u13_u7_n127, u2_u13_u7_n128, u2_u13_u7_n129, u2_u13_u7_n130, u2_u13_u7_n131, 
       u2_u13_u7_n132, u2_u13_u7_n133, u2_u13_u7_n134, u2_u13_u7_n135, u2_u13_u7_n136, u2_u13_u7_n137, u2_u13_u7_n138, u2_u13_u7_n139, u2_u13_u7_n140, 
       u2_u13_u7_n141, u2_u13_u7_n142, u2_u13_u7_n143, u2_u13_u7_n144, u2_u13_u7_n145, u2_u13_u7_n146, u2_u13_u7_n147, u2_u13_u7_n148, u2_u13_u7_n149, 
       u2_u13_u7_n150, u2_u13_u7_n151, u2_u13_u7_n152, u2_u13_u7_n153, u2_u13_u7_n154, u2_u13_u7_n155, u2_u13_u7_n156, u2_u13_u7_n157, u2_u13_u7_n158, 
       u2_u13_u7_n159, u2_u13_u7_n160, u2_u13_u7_n161, u2_u13_u7_n162, u2_u13_u7_n163, u2_u13_u7_n164, u2_u13_u7_n165, u2_u13_u7_n166, u2_u13_u7_n167, 
       u2_u13_u7_n168, u2_u13_u7_n169, u2_u13_u7_n170, u2_u13_u7_n171, u2_u13_u7_n172, u2_u13_u7_n173, u2_u13_u7_n174, u2_u13_u7_n175, u2_u13_u7_n176, 
       u2_u13_u7_n177, u2_u13_u7_n178, u2_u13_u7_n179, u2_u13_u7_n180, u2_u13_u7_n91, u2_u13_u7_n92, u2_u13_u7_n93, u2_u13_u7_n94, u2_u13_u7_n95, 
       u2_u13_u7_n96, u2_u13_u7_n97, u2_u13_u7_n98, u2_u13_u7_n99, u2_u14_X_1, u2_u14_X_12, u2_u14_X_14, u2_u14_X_17, u2_u14_X_19, 
       u2_u14_X_2, u2_u14_X_23, u2_u14_X_24, u2_u14_X_25, u2_u14_X_26, u2_u14_X_29, u2_u14_X_31, u2_u14_X_33, u2_u14_X_35, 
       u2_u14_X_36, u2_u14_X_37, u2_u14_X_38, u2_u14_X_40, u2_u14_X_42, u2_u14_X_44, u2_u14_X_47, u2_u14_X_48, u2_u14_X_6, 
       u2_u14_X_8, u2_u14_u0_n100, u2_u14_u0_n101, u2_u14_u0_n102, u2_u14_u0_n103, u2_u14_u0_n104, u2_u14_u0_n105, u2_u14_u0_n106, u2_u14_u0_n107, 
       u2_u14_u0_n108, u2_u14_u0_n109, u2_u14_u0_n110, u2_u14_u0_n111, u2_u14_u0_n112, u2_u14_u0_n113, u2_u14_u0_n114, u2_u14_u0_n115, u2_u14_u0_n116, 
       u2_u14_u0_n117, u2_u14_u0_n118, u2_u14_u0_n119, u2_u14_u0_n120, u2_u14_u0_n121, u2_u14_u0_n122, u2_u14_u0_n123, u2_u14_u0_n124, u2_u14_u0_n125, 
       u2_u14_u0_n126, u2_u14_u0_n127, u2_u14_u0_n128, u2_u14_u0_n129, u2_u14_u0_n130, u2_u14_u0_n131, u2_u14_u0_n132, u2_u14_u0_n133, u2_u14_u0_n134, 
       u2_u14_u0_n135, u2_u14_u0_n136, u2_u14_u0_n137, u2_u14_u0_n138, u2_u14_u0_n139, u2_u14_u0_n140, u2_u14_u0_n141, u2_u14_u0_n142, u2_u14_u0_n143, 
       u2_u14_u0_n144, u2_u14_u0_n145, u2_u14_u0_n146, u2_u14_u0_n147, u2_u14_u0_n148, u2_u14_u0_n149, u2_u14_u0_n150, u2_u14_u0_n151, u2_u14_u0_n152, 
       u2_u14_u0_n153, u2_u14_u0_n154, u2_u14_u0_n155, u2_u14_u0_n156, u2_u14_u0_n157, u2_u14_u0_n158, u2_u14_u0_n159, u2_u14_u0_n160, u2_u14_u0_n161, 
       u2_u14_u0_n162, u2_u14_u0_n163, u2_u14_u0_n164, u2_u14_u0_n165, u2_u14_u0_n166, u2_u14_u0_n167, u2_u14_u0_n168, u2_u14_u0_n169, u2_u14_u0_n170, 
       u2_u14_u0_n171, u2_u14_u0_n172, u2_u14_u0_n173, u2_u14_u0_n174, u2_u14_u0_n88, u2_u14_u0_n89, u2_u14_u0_n90, u2_u14_u0_n91, u2_u14_u0_n92, 
       u2_u14_u0_n93, u2_u14_u0_n94, u2_u14_u0_n95, u2_u14_u0_n96, u2_u14_u0_n97, u2_u14_u0_n98, u2_u14_u0_n99, u2_u14_u1_n100, u2_u14_u1_n101, 
       u2_u14_u1_n102, u2_u14_u1_n103, u2_u14_u1_n104, u2_u14_u1_n105, u2_u14_u1_n106, u2_u14_u1_n107, u2_u14_u1_n108, u2_u14_u1_n109, u2_u14_u1_n110, 
       u2_u14_u1_n111, u2_u14_u1_n112, u2_u14_u1_n113, u2_u14_u1_n114, u2_u14_u1_n115, u2_u14_u1_n116, u2_u14_u1_n117, u2_u14_u1_n118, u2_u14_u1_n119, 
       u2_u14_u1_n120, u2_u14_u1_n121, u2_u14_u1_n122, u2_u14_u1_n123, u2_u14_u1_n124, u2_u14_u1_n125, u2_u14_u1_n126, u2_u14_u1_n127, u2_u14_u1_n128, 
       u2_u14_u1_n129, u2_u14_u1_n130, u2_u14_u1_n131, u2_u14_u1_n132, u2_u14_u1_n133, u2_u14_u1_n134, u2_u14_u1_n135, u2_u14_u1_n136, u2_u14_u1_n137, 
       u2_u14_u1_n138, u2_u14_u1_n139, u2_u14_u1_n140, u2_u14_u1_n141, u2_u14_u1_n142, u2_u14_u1_n143, u2_u14_u1_n144, u2_u14_u1_n145, u2_u14_u1_n146, 
       u2_u14_u1_n147, u2_u14_u1_n148, u2_u14_u1_n149, u2_u14_u1_n150, u2_u14_u1_n151, u2_u14_u1_n152, u2_u14_u1_n153, u2_u14_u1_n154, u2_u14_u1_n155, 
       u2_u14_u1_n156, u2_u14_u1_n157, u2_u14_u1_n158, u2_u14_u1_n159, u2_u14_u1_n160, u2_u14_u1_n161, u2_u14_u1_n162, u2_u14_u1_n163, u2_u14_u1_n164, 
       u2_u14_u1_n165, u2_u14_u1_n166, u2_u14_u1_n167, u2_u14_u1_n168, u2_u14_u1_n169, u2_u14_u1_n170, u2_u14_u1_n171, u2_u14_u1_n172, u2_u14_u1_n173, 
       u2_u14_u1_n174, u2_u14_u1_n175, u2_u14_u1_n176, u2_u14_u1_n177, u2_u14_u1_n178, u2_u14_u1_n179, u2_u14_u1_n180, u2_u14_u1_n181, u2_u14_u1_n182, 
       u2_u14_u1_n183, u2_u14_u1_n184, u2_u14_u1_n185, u2_u14_u1_n186, u2_u14_u1_n187, u2_u14_u1_n188, u2_u14_u1_n95, u2_u14_u1_n96, u2_u14_u1_n97, 
       u2_u14_u1_n98, u2_u14_u1_n99, u2_u14_u2_n100, u2_u14_u2_n101, u2_u14_u2_n102, u2_u14_u2_n103, u2_u14_u2_n104, u2_u14_u2_n105, u2_u14_u2_n106, 
       u2_u14_u2_n107, u2_u14_u2_n108, u2_u14_u2_n109, u2_u14_u2_n110, u2_u14_u2_n111, u2_u14_u2_n112, u2_u14_u2_n113, u2_u14_u2_n114, u2_u14_u2_n115, 
       u2_u14_u2_n116, u2_u14_u2_n117, u2_u14_u2_n118, u2_u14_u2_n119, u2_u14_u2_n120, u2_u14_u2_n121, u2_u14_u2_n122, u2_u14_u2_n123, u2_u14_u2_n124, 
       u2_u14_u2_n125, u2_u14_u2_n126, u2_u14_u2_n127, u2_u14_u2_n128, u2_u14_u2_n129, u2_u14_u2_n130, u2_u14_u2_n131, u2_u14_u2_n132, u2_u14_u2_n133, 
       u2_u14_u2_n134, u2_u14_u2_n135, u2_u14_u2_n136, u2_u14_u2_n137, u2_u14_u2_n138, u2_u14_u2_n139, u2_u14_u2_n140, u2_u14_u2_n141, u2_u14_u2_n142, 
       u2_u14_u2_n143, u2_u14_u2_n144, u2_u14_u2_n145, u2_u14_u2_n146, u2_u14_u2_n147, u2_u14_u2_n148, u2_u14_u2_n149, u2_u14_u2_n150, u2_u14_u2_n151, 
       u2_u14_u2_n152, u2_u14_u2_n153, u2_u14_u2_n154, u2_u14_u2_n155, u2_u14_u2_n156, u2_u14_u2_n157, u2_u14_u2_n158, u2_u14_u2_n159, u2_u14_u2_n160, 
       u2_u14_u2_n161, u2_u14_u2_n162, u2_u14_u2_n163, u2_u14_u2_n164, u2_u14_u2_n165, u2_u14_u2_n166, u2_u14_u2_n167, u2_u14_u2_n168, u2_u14_u2_n169, 
       u2_u14_u2_n170, u2_u14_u2_n171, u2_u14_u2_n172, u2_u14_u2_n173, u2_u14_u2_n174, u2_u14_u2_n175, u2_u14_u2_n176, u2_u14_u2_n177, u2_u14_u2_n178, 
       u2_u14_u2_n179, u2_u14_u2_n180, u2_u14_u2_n181, u2_u14_u2_n182, u2_u14_u2_n183, u2_u14_u2_n184, u2_u14_u2_n185, u2_u14_u2_n186, u2_u14_u2_n187, 
       u2_u14_u2_n188, u2_u14_u2_n95, u2_u14_u2_n96, u2_u14_u2_n97, u2_u14_u2_n98, u2_u14_u2_n99, u2_u14_u3_n100, u2_u14_u3_n101, u2_u14_u3_n102, 
       u2_u14_u3_n103, u2_u14_u3_n104, u2_u14_u3_n105, u2_u14_u3_n106, u2_u14_u3_n107, u2_u14_u3_n108, u2_u14_u3_n109, u2_u14_u3_n110, u2_u14_u3_n111, 
       u2_u14_u3_n112, u2_u14_u3_n113, u2_u14_u3_n114, u2_u14_u3_n115, u2_u14_u3_n116, u2_u14_u3_n117, u2_u14_u3_n118, u2_u14_u3_n119, u2_u14_u3_n120, 
       u2_u14_u3_n121, u2_u14_u3_n122, u2_u14_u3_n123, u2_u14_u3_n124, u2_u14_u3_n125, u2_u14_u3_n126, u2_u14_u3_n127, u2_u14_u3_n128, u2_u14_u3_n129, 
       u2_u14_u3_n130, u2_u14_u3_n131, u2_u14_u3_n132, u2_u14_u3_n133, u2_u14_u3_n134, u2_u14_u3_n135, u2_u14_u3_n136, u2_u14_u3_n137, u2_u14_u3_n138, 
       u2_u14_u3_n139, u2_u14_u3_n140, u2_u14_u3_n141, u2_u14_u3_n142, u2_u14_u3_n143, u2_u14_u3_n144, u2_u14_u3_n145, u2_u14_u3_n146, u2_u14_u3_n147, 
       u2_u14_u3_n148, u2_u14_u3_n149, u2_u14_u3_n150, u2_u14_u3_n151, u2_u14_u3_n152, u2_u14_u3_n153, u2_u14_u3_n154, u2_u14_u3_n155, u2_u14_u3_n156, 
       u2_u14_u3_n157, u2_u14_u3_n158, u2_u14_u3_n159, u2_u14_u3_n160, u2_u14_u3_n161, u2_u14_u3_n162, u2_u14_u3_n163, u2_u14_u3_n164, u2_u14_u3_n165, 
       u2_u14_u3_n166, u2_u14_u3_n167, u2_u14_u3_n168, u2_u14_u3_n169, u2_u14_u3_n170, u2_u14_u3_n171, u2_u14_u3_n172, u2_u14_u3_n173, u2_u14_u3_n174, 
       u2_u14_u3_n175, u2_u14_u3_n176, u2_u14_u3_n177, u2_u14_u3_n178, u2_u14_u3_n179, u2_u14_u3_n180, u2_u14_u3_n181, u2_u14_u3_n182, u2_u14_u3_n183, 
       u2_u14_u3_n184, u2_u14_u3_n185, u2_u14_u3_n186, u2_u14_u3_n94, u2_u14_u3_n95, u2_u14_u3_n96, u2_u14_u3_n97, u2_u14_u3_n98, u2_u14_u3_n99, 
       u2_u14_u4_n100, u2_u14_u4_n101, u2_u14_u4_n102, u2_u14_u4_n103, u2_u14_u4_n104, u2_u14_u4_n105, u2_u14_u4_n106, u2_u14_u4_n107, u2_u14_u4_n108, 
       u2_u14_u4_n109, u2_u14_u4_n110, u2_u14_u4_n111, u2_u14_u4_n112, u2_u14_u4_n113, u2_u14_u4_n114, u2_u14_u4_n115, u2_u14_u4_n116, u2_u14_u4_n117, 
       u2_u14_u4_n118, u2_u14_u4_n119, u2_u14_u4_n120, u2_u14_u4_n121, u2_u14_u4_n122, u2_u14_u4_n123, u2_u14_u4_n124, u2_u14_u4_n125, u2_u14_u4_n126, 
       u2_u14_u4_n127, u2_u14_u4_n128, u2_u14_u4_n129, u2_u14_u4_n130, u2_u14_u4_n131, u2_u14_u4_n132, u2_u14_u4_n133, u2_u14_u4_n134, u2_u14_u4_n135, 
       u2_u14_u4_n136, u2_u14_u4_n137, u2_u14_u4_n138, u2_u14_u4_n139, u2_u14_u4_n140, u2_u14_u4_n141, u2_u14_u4_n142, u2_u14_u4_n143, u2_u14_u4_n144, 
       u2_u14_u4_n145, u2_u14_u4_n146, u2_u14_u4_n147, u2_u14_u4_n148, u2_u14_u4_n149, u2_u14_u4_n150, u2_u14_u4_n151, u2_u14_u4_n152, u2_u14_u4_n153, 
       u2_u14_u4_n154, u2_u14_u4_n155, u2_u14_u4_n156, u2_u14_u4_n157, u2_u14_u4_n158, u2_u14_u4_n159, u2_u14_u4_n160, u2_u14_u4_n161, u2_u14_u4_n162, 
       u2_u14_u4_n163, u2_u14_u4_n164, u2_u14_u4_n165, u2_u14_u4_n166, u2_u14_u4_n167, u2_u14_u4_n168, u2_u14_u4_n169, u2_u14_u4_n170, u2_u14_u4_n171, 
       u2_u14_u4_n172, u2_u14_u4_n173, u2_u14_u4_n174, u2_u14_u4_n175, u2_u14_u4_n176, u2_u14_u4_n177, u2_u14_u4_n178, u2_u14_u4_n179, u2_u14_u4_n180, 
       u2_u14_u4_n181, u2_u14_u4_n182, u2_u14_u4_n183, u2_u14_u4_n184, u2_u14_u4_n185, u2_u14_u4_n186, u2_u14_u4_n94, u2_u14_u4_n95, u2_u14_u4_n96, 
       u2_u14_u4_n97, u2_u14_u4_n98, u2_u14_u4_n99, u2_u14_u5_n100, u2_u14_u5_n101, u2_u14_u5_n102, u2_u14_u5_n103, u2_u14_u5_n104, u2_u14_u5_n105, 
       u2_u14_u5_n106, u2_u14_u5_n107, u2_u14_u5_n108, u2_u14_u5_n109, u2_u14_u5_n110, u2_u14_u5_n111, u2_u14_u5_n112, u2_u14_u5_n113, u2_u14_u5_n114, 
       u2_u14_u5_n115, u2_u14_u5_n116, u2_u14_u5_n117, u2_u14_u5_n118, u2_u14_u5_n119, u2_u14_u5_n120, u2_u14_u5_n121, u2_u14_u5_n122, u2_u14_u5_n123, 
       u2_u14_u5_n124, u2_u14_u5_n125, u2_u14_u5_n126, u2_u14_u5_n127, u2_u14_u5_n128, u2_u14_u5_n129, u2_u14_u5_n130, u2_u14_u5_n131, u2_u14_u5_n132, 
       u2_u14_u5_n133, u2_u14_u5_n134, u2_u14_u5_n135, u2_u14_u5_n136, u2_u14_u5_n137, u2_u14_u5_n138, u2_u14_u5_n139, u2_u14_u5_n140, u2_u14_u5_n141, 
       u2_u14_u5_n142, u2_u14_u5_n143, u2_u14_u5_n144, u2_u14_u5_n145, u2_u14_u5_n146, u2_u14_u5_n147, u2_u14_u5_n148, u2_u14_u5_n149, u2_u14_u5_n150, 
       u2_u14_u5_n151, u2_u14_u5_n152, u2_u14_u5_n153, u2_u14_u5_n154, u2_u14_u5_n155, u2_u14_u5_n156, u2_u14_u5_n157, u2_u14_u5_n158, u2_u14_u5_n159, 
       u2_u14_u5_n160, u2_u14_u5_n161, u2_u14_u5_n162, u2_u14_u5_n163, u2_u14_u5_n164, u2_u14_u5_n165, u2_u14_u5_n166, u2_u14_u5_n167, u2_u14_u5_n168, 
       u2_u14_u5_n169, u2_u14_u5_n170, u2_u14_u5_n171, u2_u14_u5_n172, u2_u14_u5_n173, u2_u14_u5_n174, u2_u14_u5_n175, u2_u14_u5_n176, u2_u14_u5_n177, 
       u2_u14_u5_n178, u2_u14_u5_n179, u2_u14_u5_n180, u2_u14_u5_n181, u2_u14_u5_n182, u2_u14_u5_n183, u2_u14_u5_n184, u2_u14_u5_n185, u2_u14_u5_n186, 
       u2_u14_u5_n187, u2_u14_u5_n188, u2_u14_u5_n189, u2_u14_u5_n190, u2_u14_u5_n191, u2_u14_u5_n192, u2_u14_u5_n193, u2_u14_u5_n194, u2_u14_u5_n195, 
       u2_u14_u5_n196, u2_u14_u5_n99, u2_u14_u6_n100, u2_u14_u6_n101, u2_u14_u6_n102, u2_u14_u6_n103, u2_u14_u6_n104, u2_u14_u6_n105, u2_u14_u6_n106, 
       u2_u14_u6_n107, u2_u14_u6_n108, u2_u14_u6_n109, u2_u14_u6_n110, u2_u14_u6_n111, u2_u14_u6_n112, u2_u14_u6_n113, u2_u14_u6_n114, u2_u14_u6_n115, 
       u2_u14_u6_n116, u2_u14_u6_n117, u2_u14_u6_n118, u2_u14_u6_n119, u2_u14_u6_n120, u2_u14_u6_n121, u2_u14_u6_n122, u2_u14_u6_n123, u2_u14_u6_n124, 
       u2_u14_u6_n125, u2_u14_u6_n126, u2_u14_u6_n127, u2_u14_u6_n128, u2_u14_u6_n129, u2_u14_u6_n130, u2_u14_u6_n131, u2_u14_u6_n132, u2_u14_u6_n133, 
       u2_u14_u6_n134, u2_u14_u6_n135, u2_u14_u6_n136, u2_u14_u6_n137, u2_u14_u6_n138, u2_u14_u6_n139, u2_u14_u6_n140, u2_u14_u6_n141, u2_u14_u6_n142, 
       u2_u14_u6_n143, u2_u14_u6_n144, u2_u14_u6_n145, u2_u14_u6_n146, u2_u14_u6_n147, u2_u14_u6_n148, u2_u14_u6_n149, u2_u14_u6_n150, u2_u14_u6_n151, 
       u2_u14_u6_n152, u2_u14_u6_n153, u2_u14_u6_n154, u2_u14_u6_n155, u2_u14_u6_n156, u2_u14_u6_n157, u2_u14_u6_n158, u2_u14_u6_n159, u2_u14_u6_n160, 
       u2_u14_u6_n161, u2_u14_u6_n162, u2_u14_u6_n163, u2_u14_u6_n164, u2_u14_u6_n165, u2_u14_u6_n166, u2_u14_u6_n167, u2_u14_u6_n168, u2_u14_u6_n169, 
       u2_u14_u6_n170, u2_u14_u6_n171, u2_u14_u6_n172, u2_u14_u6_n173, u2_u14_u6_n174, u2_u14_u6_n88, u2_u14_u6_n89, u2_u14_u6_n90, u2_u14_u6_n91, 
       u2_u14_u6_n92, u2_u14_u6_n93, u2_u14_u6_n94, u2_u14_u6_n95, u2_u14_u6_n96, u2_u14_u6_n97, u2_u14_u6_n98, u2_u14_u6_n99, u2_u14_u7_n100, 
       u2_u14_u7_n101, u2_u14_u7_n102, u2_u14_u7_n103, u2_u14_u7_n104, u2_u14_u7_n105, u2_u14_u7_n106, u2_u14_u7_n107, u2_u14_u7_n108, u2_u14_u7_n109, 
       u2_u14_u7_n110, u2_u14_u7_n111, u2_u14_u7_n112, u2_u14_u7_n113, u2_u14_u7_n114, u2_u14_u7_n115, u2_u14_u7_n116, u2_u14_u7_n117, u2_u14_u7_n118, 
       u2_u14_u7_n119, u2_u14_u7_n120, u2_u14_u7_n121, u2_u14_u7_n122, u2_u14_u7_n123, u2_u14_u7_n124, u2_u14_u7_n125, u2_u14_u7_n126, u2_u14_u7_n127, 
       u2_u14_u7_n128, u2_u14_u7_n129, u2_u14_u7_n130, u2_u14_u7_n131, u2_u14_u7_n132, u2_u14_u7_n133, u2_u14_u7_n134, u2_u14_u7_n135, u2_u14_u7_n136, 
       u2_u14_u7_n137, u2_u14_u7_n138, u2_u14_u7_n139, u2_u14_u7_n140, u2_u14_u7_n141, u2_u14_u7_n142, u2_u14_u7_n143, u2_u14_u7_n144, u2_u14_u7_n145, 
       u2_u14_u7_n146, u2_u14_u7_n147, u2_u14_u7_n148, u2_u14_u7_n149, u2_u14_u7_n150, u2_u14_u7_n151, u2_u14_u7_n152, u2_u14_u7_n153, u2_u14_u7_n154, 
       u2_u14_u7_n155, u2_u14_u7_n156, u2_u14_u7_n157, u2_u14_u7_n158, u2_u14_u7_n159, u2_u14_u7_n160, u2_u14_u7_n161, u2_u14_u7_n162, u2_u14_u7_n163, 
       u2_u14_u7_n164, u2_u14_u7_n165, u2_u14_u7_n166, u2_u14_u7_n167, u2_u14_u7_n168, u2_u14_u7_n169, u2_u14_u7_n170, u2_u14_u7_n171, u2_u14_u7_n172, 
       u2_u14_u7_n173, u2_u14_u7_n174, u2_u14_u7_n175, u2_u14_u7_n176, u2_u14_u7_n177, u2_u14_u7_n178, u2_u14_u7_n179, u2_u14_u7_n180, u2_u14_u7_n91, 
       u2_u14_u7_n92, u2_u14_u7_n93, u2_u14_u7_n94, u2_u14_u7_n95, u2_u14_u7_n96, u2_u14_u7_n97, u2_u14_u7_n98, u2_u14_u7_n99, u2_u2_X_1, 
       u2_u2_X_10, u2_u2_X_11, u2_u2_X_12, u2_u2_X_13, u2_u2_X_14, u2_u2_X_17, u2_u2_X_18, u2_u2_X_19, u2_u2_X_2, 
       u2_u2_X_20, u2_u2_X_21, u2_u2_X_22, u2_u2_X_23, u2_u2_X_24, u2_u2_X_25, u2_u2_X_26, u2_u2_X_3, u2_u2_X_36, 
       u2_u2_X_38, u2_u2_X_4, u2_u2_X_40, u2_u2_X_41, u2_u2_X_42, u2_u2_X_43, u2_u2_X_44, u2_u2_X_45, u2_u2_X_46, 
       u2_u2_X_47, u2_u2_X_48, u2_u2_X_6, u2_u2_X_8, u2_u2_X_9, u2_u2_u0_n100, u2_u2_u0_n101, u2_u2_u0_n102, u2_u2_u0_n103, 
       u2_u2_u0_n104, u2_u2_u0_n105, u2_u2_u0_n106, u2_u2_u0_n107, u2_u2_u0_n108, u2_u2_u0_n109, u2_u2_u0_n110, u2_u2_u0_n111, u2_u2_u0_n112, 
       u2_u2_u0_n113, u2_u2_u0_n114, u2_u2_u0_n115, u2_u2_u0_n116, u2_u2_u0_n117, u2_u2_u0_n118, u2_u2_u0_n119, u2_u2_u0_n120, u2_u2_u0_n121, 
       u2_u2_u0_n122, u2_u2_u0_n123, u2_u2_u0_n124, u2_u2_u0_n125, u2_u2_u0_n126, u2_u2_u0_n127, u2_u2_u0_n128, u2_u2_u0_n129, u2_u2_u0_n130, 
       u2_u2_u0_n131, u2_u2_u0_n132, u2_u2_u0_n133, u2_u2_u0_n134, u2_u2_u0_n135, u2_u2_u0_n136, u2_u2_u0_n137, u2_u2_u0_n138, u2_u2_u0_n139, 
       u2_u2_u0_n140, u2_u2_u0_n141, u2_u2_u0_n142, u2_u2_u0_n143, u2_u2_u0_n144, u2_u2_u0_n145, u2_u2_u0_n146, u2_u2_u0_n147, u2_u2_u0_n148, 
       u2_u2_u0_n149, u2_u2_u0_n150, u2_u2_u0_n151, u2_u2_u0_n152, u2_u2_u0_n153, u2_u2_u0_n154, u2_u2_u0_n155, u2_u2_u0_n156, u2_u2_u0_n157, 
       u2_u2_u0_n158, u2_u2_u0_n159, u2_u2_u0_n160, u2_u2_u0_n161, u2_u2_u0_n162, u2_u2_u0_n163, u2_u2_u0_n164, u2_u2_u0_n165, u2_u2_u0_n166, 
       u2_u2_u0_n167, u2_u2_u0_n168, u2_u2_u0_n169, u2_u2_u0_n170, u2_u2_u0_n171, u2_u2_u0_n172, u2_u2_u0_n173, u2_u2_u0_n174, u2_u2_u0_n88, 
       u2_u2_u0_n89, u2_u2_u0_n90, u2_u2_u0_n91, u2_u2_u0_n92, u2_u2_u0_n93, u2_u2_u0_n94, u2_u2_u0_n95, u2_u2_u0_n96, u2_u2_u0_n97, 
       u2_u2_u0_n98, u2_u2_u0_n99, u2_u2_u1_n100, u2_u2_u1_n101, u2_u2_u1_n102, u2_u2_u1_n103, u2_u2_u1_n104, u2_u2_u1_n105, u2_u2_u1_n106, 
       u2_u2_u1_n107, u2_u2_u1_n108, u2_u2_u1_n109, u2_u2_u1_n110, u2_u2_u1_n111, u2_u2_u1_n112, u2_u2_u1_n113, u2_u2_u1_n114, u2_u2_u1_n115, 
       u2_u2_u1_n116, u2_u2_u1_n117, u2_u2_u1_n118, u2_u2_u1_n119, u2_u2_u1_n120, u2_u2_u1_n121, u2_u2_u1_n122, u2_u2_u1_n123, u2_u2_u1_n124, 
       u2_u2_u1_n125, u2_u2_u1_n126, u2_u2_u1_n127, u2_u2_u1_n128, u2_u2_u1_n129, u2_u2_u1_n130, u2_u2_u1_n131, u2_u2_u1_n132, u2_u2_u1_n133, 
       u2_u2_u1_n134, u2_u2_u1_n135, u2_u2_u1_n136, u2_u2_u1_n137, u2_u2_u1_n138, u2_u2_u1_n139, u2_u2_u1_n140, u2_u2_u1_n141, u2_u2_u1_n142, 
       u2_u2_u1_n143, u2_u2_u1_n144, u2_u2_u1_n145, u2_u2_u1_n146, u2_u2_u1_n147, u2_u2_u1_n148, u2_u2_u1_n149, u2_u2_u1_n150, u2_u2_u1_n151, 
       u2_u2_u1_n152, u2_u2_u1_n153, u2_u2_u1_n154, u2_u2_u1_n155, u2_u2_u1_n156, u2_u2_u1_n157, u2_u2_u1_n158, u2_u2_u1_n159, u2_u2_u1_n160, 
       u2_u2_u1_n161, u2_u2_u1_n162, u2_u2_u1_n163, u2_u2_u1_n164, u2_u2_u1_n165, u2_u2_u1_n166, u2_u2_u1_n167, u2_u2_u1_n168, u2_u2_u1_n169, 
       u2_u2_u1_n170, u2_u2_u1_n171, u2_u2_u1_n172, u2_u2_u1_n173, u2_u2_u1_n174, u2_u2_u1_n175, u2_u2_u1_n176, u2_u2_u1_n177, u2_u2_u1_n178, 
       u2_u2_u1_n179, u2_u2_u1_n180, u2_u2_u1_n181, u2_u2_u1_n182, u2_u2_u1_n183, u2_u2_u1_n184, u2_u2_u1_n185, u2_u2_u1_n186, u2_u2_u1_n187, 
       u2_u2_u1_n188, u2_u2_u1_n95, u2_u2_u1_n96, u2_u2_u1_n97, u2_u2_u1_n98, u2_u2_u1_n99, u2_u2_u2_n100, u2_u2_u2_n101, u2_u2_u2_n102, 
       u2_u2_u2_n103, u2_u2_u2_n104, u2_u2_u2_n105, u2_u2_u2_n106, u2_u2_u2_n107, u2_u2_u2_n108, u2_u2_u2_n109, u2_u2_u2_n110, u2_u2_u2_n111, 
       u2_u2_u2_n112, u2_u2_u2_n113, u2_u2_u2_n114, u2_u2_u2_n115, u2_u2_u2_n116, u2_u2_u2_n117, u2_u2_u2_n118, u2_u2_u2_n119, u2_u2_u2_n120, 
       u2_u2_u2_n121, u2_u2_u2_n122, u2_u2_u2_n123, u2_u2_u2_n124, u2_u2_u2_n125, u2_u2_u2_n126, u2_u2_u2_n127, u2_u2_u2_n128, u2_u2_u2_n129, 
       u2_u2_u2_n130, u2_u2_u2_n131, u2_u2_u2_n132, u2_u2_u2_n133, u2_u2_u2_n134, u2_u2_u2_n135, u2_u2_u2_n136, u2_u2_u2_n137, u2_u2_u2_n138, 
       u2_u2_u2_n139, u2_u2_u2_n140, u2_u2_u2_n141, u2_u2_u2_n142, u2_u2_u2_n143, u2_u2_u2_n144, u2_u2_u2_n145, u2_u2_u2_n146, u2_u2_u2_n147, 
       u2_u2_u2_n148, u2_u2_u2_n149, u2_u2_u2_n150, u2_u2_u2_n151, u2_u2_u2_n152, u2_u2_u2_n153, u2_u2_u2_n154, u2_u2_u2_n155, u2_u2_u2_n156, 
       u2_u2_u2_n157, u2_u2_u2_n158, u2_u2_u2_n159, u2_u2_u2_n160, u2_u2_u2_n161, u2_u2_u2_n162, u2_u2_u2_n163, u2_u2_u2_n164, u2_u2_u2_n165, 
       u2_u2_u2_n166, u2_u2_u2_n167, u2_u2_u2_n168, u2_u2_u2_n169, u2_u2_u2_n170, u2_u2_u2_n171, u2_u2_u2_n172, u2_u2_u2_n173, u2_u2_u2_n174, 
       u2_u2_u2_n175, u2_u2_u2_n176, u2_u2_u2_n177, u2_u2_u2_n178, u2_u2_u2_n179, u2_u2_u2_n180, u2_u2_u2_n181, u2_u2_u2_n182, u2_u2_u2_n183, 
       u2_u2_u2_n184, u2_u2_u2_n185, u2_u2_u2_n186, u2_u2_u2_n187, u2_u2_u2_n188, u2_u2_u2_n95, u2_u2_u2_n96, u2_u2_u2_n97, u2_u2_u2_n98, 
       u2_u2_u2_n99, u2_u2_u3_n100, u2_u2_u3_n101, u2_u2_u3_n102, u2_u2_u3_n103, u2_u2_u3_n104, u2_u2_u3_n105, u2_u2_u3_n106, u2_u2_u3_n107, 
       u2_u2_u3_n108, u2_u2_u3_n109, u2_u2_u3_n110, u2_u2_u3_n111, u2_u2_u3_n112, u2_u2_u3_n113, u2_u2_u3_n114, u2_u2_u3_n115, u2_u2_u3_n116, 
       u2_u2_u3_n117, u2_u2_u3_n118, u2_u2_u3_n119, u2_u2_u3_n120, u2_u2_u3_n121, u2_u2_u3_n122, u2_u2_u3_n123, u2_u2_u3_n124, u2_u2_u3_n125, 
       u2_u2_u3_n126, u2_u2_u3_n127, u2_u2_u3_n128, u2_u2_u3_n129, u2_u2_u3_n130, u2_u2_u3_n131, u2_u2_u3_n132, u2_u2_u3_n133, u2_u2_u3_n134, 
       u2_u2_u3_n135, u2_u2_u3_n136, u2_u2_u3_n137, u2_u2_u3_n138, u2_u2_u3_n139, u2_u2_u3_n140, u2_u2_u3_n141, u2_u2_u3_n142, u2_u2_u3_n143, 
       u2_u2_u3_n144, u2_u2_u3_n145, u2_u2_u3_n146, u2_u2_u3_n147, u2_u2_u3_n148, u2_u2_u3_n149, u2_u2_u3_n150, u2_u2_u3_n151, u2_u2_u3_n152, 
       u2_u2_u3_n153, u2_u2_u3_n154, u2_u2_u3_n155, u2_u2_u3_n156, u2_u2_u3_n157, u2_u2_u3_n158, u2_u2_u3_n159, u2_u2_u3_n160, u2_u2_u3_n161, 
       u2_u2_u3_n162, u2_u2_u3_n163, u2_u2_u3_n164, u2_u2_u3_n165, u2_u2_u3_n166, u2_u2_u3_n167, u2_u2_u3_n168, u2_u2_u3_n169, u2_u2_u3_n170, 
       u2_u2_u3_n171, u2_u2_u3_n172, u2_u2_u3_n173, u2_u2_u3_n174, u2_u2_u3_n175, u2_u2_u3_n176, u2_u2_u3_n177, u2_u2_u3_n178, u2_u2_u3_n179, 
       u2_u2_u3_n180, u2_u2_u3_n181, u2_u2_u3_n182, u2_u2_u3_n183, u2_u2_u3_n184, u2_u2_u3_n185, u2_u2_u3_n186, u2_u2_u3_n94, u2_u2_u3_n95, 
       u2_u2_u3_n96, u2_u2_u3_n97, u2_u2_u3_n98, u2_u2_u3_n99, u2_u2_u4_n100, u2_u2_u4_n101, u2_u2_u4_n102, u2_u2_u4_n103, u2_u2_u4_n104, 
       u2_u2_u4_n105, u2_u2_u4_n106, u2_u2_u4_n107, u2_u2_u4_n108, u2_u2_u4_n109, u2_u2_u4_n110, u2_u2_u4_n111, u2_u2_u4_n112, u2_u2_u4_n113, 
       u2_u2_u4_n114, u2_u2_u4_n115, u2_u2_u4_n116, u2_u2_u4_n117, u2_u2_u4_n118, u2_u2_u4_n119, u2_u2_u4_n120, u2_u2_u4_n121, u2_u2_u4_n122, 
       u2_u2_u4_n123, u2_u2_u4_n124, u2_u2_u4_n125, u2_u2_u4_n126, u2_u2_u4_n127, u2_u2_u4_n128, u2_u2_u4_n129, u2_u2_u4_n130, u2_u2_u4_n131, 
       u2_u2_u4_n132, u2_u2_u4_n133, u2_u2_u4_n134, u2_u2_u4_n135, u2_u2_u4_n136, u2_u2_u4_n137, u2_u2_u4_n138, u2_u2_u4_n139, u2_u2_u4_n140, 
       u2_u2_u4_n141, u2_u2_u4_n142, u2_u2_u4_n143, u2_u2_u4_n144, u2_u2_u4_n145, u2_u2_u4_n146, u2_u2_u4_n147, u2_u2_u4_n148, u2_u2_u4_n149, 
       u2_u2_u4_n150, u2_u2_u4_n151, u2_u2_u4_n152, u2_u2_u4_n153, u2_u2_u4_n154, u2_u2_u4_n155, u2_u2_u4_n156, u2_u2_u4_n157, u2_u2_u4_n158, 
       u2_u2_u4_n159, u2_u2_u4_n160, u2_u2_u4_n161, u2_u2_u4_n162, u2_u2_u4_n163, u2_u2_u4_n164, u2_u2_u4_n165, u2_u2_u4_n166, u2_u2_u4_n167, 
       u2_u2_u4_n168, u2_u2_u4_n169, u2_u2_u4_n170, u2_u2_u4_n171, u2_u2_u4_n172, u2_u2_u4_n173, u2_u2_u4_n174, u2_u2_u4_n175, u2_u2_u4_n176, 
       u2_u2_u4_n177, u2_u2_u4_n178, u2_u2_u4_n179, u2_u2_u4_n180, u2_u2_u4_n181, u2_u2_u4_n182, u2_u2_u4_n183, u2_u2_u4_n184, u2_u2_u4_n185, 
       u2_u2_u4_n186, u2_u2_u4_n94, u2_u2_u4_n95, u2_u2_u4_n96, u2_u2_u4_n97, u2_u2_u4_n98, u2_u2_u4_n99, u2_u2_u5_n100, u2_u2_u5_n101, 
       u2_u2_u5_n102, u2_u2_u5_n103, u2_u2_u5_n104, u2_u2_u5_n105, u2_u2_u5_n106, u2_u2_u5_n107, u2_u2_u5_n108, u2_u2_u5_n109, u2_u2_u5_n110, 
       u2_u2_u5_n111, u2_u2_u5_n112, u2_u2_u5_n113, u2_u2_u5_n114, u2_u2_u5_n115, u2_u2_u5_n116, u2_u2_u5_n117, u2_u2_u5_n118, u2_u2_u5_n119, 
       u2_u2_u5_n120, u2_u2_u5_n121, u2_u2_u5_n122, u2_u2_u5_n123, u2_u2_u5_n124, u2_u2_u5_n125, u2_u2_u5_n126, u2_u2_u5_n127, u2_u2_u5_n128, 
       u2_u2_u5_n129, u2_u2_u5_n130, u2_u2_u5_n131, u2_u2_u5_n132, u2_u2_u5_n133, u2_u2_u5_n134, u2_u2_u5_n135, u2_u2_u5_n136, u2_u2_u5_n137, 
       u2_u2_u5_n138, u2_u2_u5_n139, u2_u2_u5_n140, u2_u2_u5_n141, u2_u2_u5_n142, u2_u2_u5_n143, u2_u2_u5_n144, u2_u2_u5_n145, u2_u2_u5_n146, 
       u2_u2_u5_n147, u2_u2_u5_n148, u2_u2_u5_n149, u2_u2_u5_n150, u2_u2_u5_n151, u2_u2_u5_n152, u2_u2_u5_n153, u2_u2_u5_n154, u2_u2_u5_n155, 
       u2_u2_u5_n156, u2_u2_u5_n157, u2_u2_u5_n158, u2_u2_u5_n159, u2_u2_u5_n160, u2_u2_u5_n161, u2_u2_u5_n162, u2_u2_u5_n163, u2_u2_u5_n164, 
       u2_u2_u5_n165, u2_u2_u5_n166, u2_u2_u5_n167, u2_u2_u5_n168, u2_u2_u5_n169, u2_u2_u5_n170, u2_u2_u5_n171, u2_u2_u5_n172, u2_u2_u5_n173, 
       u2_u2_u5_n174, u2_u2_u5_n175, u2_u2_u5_n176, u2_u2_u5_n177, u2_u2_u5_n178, u2_u2_u5_n179, u2_u2_u5_n180, u2_u2_u5_n181, u2_u2_u5_n182, 
       u2_u2_u5_n183, u2_u2_u5_n184, u2_u2_u5_n185, u2_u2_u5_n186, u2_u2_u5_n187, u2_u2_u5_n188, u2_u2_u5_n189, u2_u2_u5_n190, u2_u2_u5_n191, 
       u2_u2_u5_n192, u2_u2_u5_n193, u2_u2_u5_n194, u2_u2_u5_n195, u2_u2_u5_n196, u2_u2_u5_n99, u2_u2_u6_n100, u2_u2_u6_n101, u2_u2_u6_n102, 
       u2_u2_u6_n103, u2_u2_u6_n104, u2_u2_u6_n105, u2_u2_u6_n106, u2_u2_u6_n107, u2_u2_u6_n108, u2_u2_u6_n109, u2_u2_u6_n110, u2_u2_u6_n111, 
       u2_u2_u6_n112, u2_u2_u6_n113, u2_u2_u6_n114, u2_u2_u6_n115, u2_u2_u6_n116, u2_u2_u6_n117, u2_u2_u6_n118, u2_u2_u6_n119, u2_u2_u6_n120, 
       u2_u2_u6_n121, u2_u2_u6_n122, u2_u2_u6_n123, u2_u2_u6_n124, u2_u2_u6_n125, u2_u2_u6_n126, u2_u2_u6_n127, u2_u2_u6_n128, u2_u2_u6_n129, 
       u2_u2_u6_n130, u2_u2_u6_n131, u2_u2_u6_n132, u2_u2_u6_n133, u2_u2_u6_n134, u2_u2_u6_n135, u2_u2_u6_n136, u2_u2_u6_n137, u2_u2_u6_n138, 
       u2_u2_u6_n139, u2_u2_u6_n140, u2_u2_u6_n141, u2_u2_u6_n142, u2_u2_u6_n143, u2_u2_u6_n144, u2_u2_u6_n145, u2_u2_u6_n146, u2_u2_u6_n147, 
       u2_u2_u6_n148, u2_u2_u6_n149, u2_u2_u6_n150, u2_u2_u6_n151, u2_u2_u6_n152, u2_u2_u6_n153, u2_u2_u6_n154, u2_u2_u6_n155, u2_u2_u6_n156, 
       u2_u2_u6_n157, u2_u2_u6_n158, u2_u2_u6_n159, u2_u2_u6_n160, u2_u2_u6_n161, u2_u2_u6_n162, u2_u2_u6_n163, u2_u2_u6_n164, u2_u2_u6_n165, 
       u2_u2_u6_n166, u2_u2_u6_n167, u2_u2_u6_n168, u2_u2_u6_n169, u2_u2_u6_n170, u2_u2_u6_n171, u2_u2_u6_n172, u2_u2_u6_n173, u2_u2_u6_n174, 
       u2_u2_u6_n88, u2_u2_u6_n89, u2_u2_u6_n90, u2_u2_u6_n91, u2_u2_u6_n92, u2_u2_u6_n93, u2_u2_u6_n94, u2_u2_u6_n95, u2_u2_u6_n96, 
       u2_u2_u6_n97, u2_u2_u6_n98, u2_u2_u6_n99, u2_u2_u7_n100, u2_u2_u7_n101, u2_u2_u7_n102, u2_u2_u7_n103, u2_u2_u7_n104, u2_u2_u7_n105, 
       u2_u2_u7_n106, u2_u2_u7_n107, u2_u2_u7_n108, u2_u2_u7_n109, u2_u2_u7_n110, u2_u2_u7_n111, u2_u2_u7_n112, u2_u2_u7_n113, u2_u2_u7_n114, 
       u2_u2_u7_n115, u2_u2_u7_n116, u2_u2_u7_n117, u2_u2_u7_n118, u2_u2_u7_n119, u2_u2_u7_n120, u2_u2_u7_n121, u2_u2_u7_n122, u2_u2_u7_n123, 
       u2_u2_u7_n124, u2_u2_u7_n125, u2_u2_u7_n126, u2_u2_u7_n127, u2_u2_u7_n128, u2_u2_u7_n129, u2_u2_u7_n130, u2_u2_u7_n131, u2_u2_u7_n132, 
       u2_u2_u7_n133, u2_u2_u7_n134, u2_u2_u7_n135, u2_u2_u7_n136, u2_u2_u7_n137, u2_u2_u7_n138, u2_u2_u7_n139, u2_u2_u7_n140, u2_u2_u7_n141, 
       u2_u2_u7_n142, u2_u2_u7_n143, u2_u2_u7_n144, u2_u2_u7_n145, u2_u2_u7_n146, u2_u2_u7_n147, u2_u2_u7_n148, u2_u2_u7_n149, u2_u2_u7_n150, 
       u2_u2_u7_n151, u2_u2_u7_n152, u2_u2_u7_n153, u2_u2_u7_n154, u2_u2_u7_n155, u2_u2_u7_n156, u2_u2_u7_n157, u2_u2_u7_n158, u2_u2_u7_n159, 
       u2_u2_u7_n160, u2_u2_u7_n161, u2_u2_u7_n162, u2_u2_u7_n163, u2_u2_u7_n164, u2_u2_u7_n165, u2_u2_u7_n166, u2_u2_u7_n167, u2_u2_u7_n168, 
       u2_u2_u7_n169, u2_u2_u7_n170, u2_u2_u7_n171, u2_u2_u7_n172, u2_u2_u7_n173, u2_u2_u7_n174, u2_u2_u7_n175, u2_u2_u7_n176, u2_u2_u7_n177, 
       u2_u2_u7_n178, u2_u2_u7_n179, u2_u2_u7_n180, u2_u2_u7_n91, u2_u2_u7_n92, u2_u2_u7_n93, u2_u2_u7_n94, u2_u2_u7_n95, u2_u2_u7_n96, 
       u2_u2_u7_n97, u2_u2_u7_n98, u2_u2_u7_n99, u2_u3_X_1, u2_u3_X_10, u2_u3_X_11, u2_u3_X_12, u2_u3_X_13, u2_u3_X_14, 
       u2_u3_X_15, u2_u3_X_16, u2_u3_X_17, u2_u3_X_18, u2_u3_X_19, u2_u3_X_2, u2_u3_X_20, u2_u3_X_23, u2_u3_X_24, 
       u2_u3_X_25, u2_u3_X_26, u2_u3_X_28, u2_u3_X_29, u2_u3_X_3, u2_u3_X_30, u2_u3_X_31, u2_u3_X_32, u2_u3_X_36, 
       u2_u3_X_4, u2_u3_X_47, u2_u3_X_48, u2_u3_X_5, u2_u3_X_6, u2_u3_X_7, u2_u3_X_8, u2_u3_X_9, u2_u3_u0_n100, 
       u2_u3_u0_n101, u2_u3_u0_n102, u2_u3_u0_n103, u2_u3_u0_n104, u2_u3_u0_n105, u2_u3_u0_n106, u2_u3_u0_n107, u2_u3_u0_n108, u2_u3_u0_n109, 
       u2_u3_u0_n110, u2_u3_u0_n111, u2_u3_u0_n112, u2_u3_u0_n113, u2_u3_u0_n114, u2_u3_u0_n115, u2_u3_u0_n116, u2_u3_u0_n117, u2_u3_u0_n118, 
       u2_u3_u0_n119, u2_u3_u0_n120, u2_u3_u0_n121, u2_u3_u0_n122, u2_u3_u0_n123, u2_u3_u0_n124, u2_u3_u0_n125, u2_u3_u0_n126, u2_u3_u0_n127, 
       u2_u3_u0_n128, u2_u3_u0_n129, u2_u3_u0_n130, u2_u3_u0_n131, u2_u3_u0_n132, u2_u3_u0_n133, u2_u3_u0_n134, u2_u3_u0_n135, u2_u3_u0_n136, 
       u2_u3_u0_n137, u2_u3_u0_n138, u2_u3_u0_n139, u2_u3_u0_n140, u2_u3_u0_n141, u2_u3_u0_n142, u2_u3_u0_n143, u2_u3_u0_n144, u2_u3_u0_n145, 
       u2_u3_u0_n146, u2_u3_u0_n147, u2_u3_u0_n148, u2_u3_u0_n149, u2_u3_u0_n150, u2_u3_u0_n151, u2_u3_u0_n152, u2_u3_u0_n153, u2_u3_u0_n154, 
       u2_u3_u0_n155, u2_u3_u0_n156, u2_u3_u0_n157, u2_u3_u0_n158, u2_u3_u0_n159, u2_u3_u0_n160, u2_u3_u0_n161, u2_u3_u0_n162, u2_u3_u0_n163, 
       u2_u3_u0_n164, u2_u3_u0_n165, u2_u3_u0_n166, u2_u3_u0_n167, u2_u3_u0_n168, u2_u3_u0_n169, u2_u3_u0_n170, u2_u3_u0_n171, u2_u3_u0_n172, 
       u2_u3_u0_n173, u2_u3_u0_n174, u2_u3_u0_n88, u2_u3_u0_n89, u2_u3_u0_n90, u2_u3_u0_n91, u2_u3_u0_n92, u2_u3_u0_n93, u2_u3_u0_n94, 
       u2_u3_u0_n95, u2_u3_u0_n96, u2_u3_u0_n97, u2_u3_u0_n98, u2_u3_u0_n99, u2_u3_u1_n100, u2_u3_u1_n101, u2_u3_u1_n102, u2_u3_u1_n103, 
       u2_u3_u1_n104, u2_u3_u1_n105, u2_u3_u1_n106, u2_u3_u1_n107, u2_u3_u1_n108, u2_u3_u1_n109, u2_u3_u1_n110, u2_u3_u1_n111, u2_u3_u1_n112, 
       u2_u3_u1_n113, u2_u3_u1_n114, u2_u3_u1_n115, u2_u3_u1_n116, u2_u3_u1_n117, u2_u3_u1_n118, u2_u3_u1_n119, u2_u3_u1_n120, u2_u3_u1_n121, 
       u2_u3_u1_n122, u2_u3_u1_n123, u2_u3_u1_n124, u2_u3_u1_n125, u2_u3_u1_n126, u2_u3_u1_n127, u2_u3_u1_n128, u2_u3_u1_n129, u2_u3_u1_n130, 
       u2_u3_u1_n131, u2_u3_u1_n132, u2_u3_u1_n133, u2_u3_u1_n134, u2_u3_u1_n135, u2_u3_u1_n136, u2_u3_u1_n137, u2_u3_u1_n138, u2_u3_u1_n139, 
       u2_u3_u1_n140, u2_u3_u1_n141, u2_u3_u1_n142, u2_u3_u1_n143, u2_u3_u1_n144, u2_u3_u1_n145, u2_u3_u1_n146, u2_u3_u1_n147, u2_u3_u1_n148, 
       u2_u3_u1_n149, u2_u3_u1_n150, u2_u3_u1_n151, u2_u3_u1_n152, u2_u3_u1_n153, u2_u3_u1_n154, u2_u3_u1_n155, u2_u3_u1_n156, u2_u3_u1_n157, 
       u2_u3_u1_n158, u2_u3_u1_n159, u2_u3_u1_n160, u2_u3_u1_n161, u2_u3_u1_n162, u2_u3_u1_n163, u2_u3_u1_n164, u2_u3_u1_n165, u2_u3_u1_n166, 
       u2_u3_u1_n167, u2_u3_u1_n168, u2_u3_u1_n169, u2_u3_u1_n170, u2_u3_u1_n171, u2_u3_u1_n172, u2_u3_u1_n173, u2_u3_u1_n174, u2_u3_u1_n175, 
       u2_u3_u1_n176, u2_u3_u1_n177, u2_u3_u1_n178, u2_u3_u1_n179, u2_u3_u1_n180, u2_u3_u1_n181, u2_u3_u1_n182, u2_u3_u1_n183, u2_u3_u1_n184, 
       u2_u3_u1_n185, u2_u3_u1_n186, u2_u3_u1_n187, u2_u3_u1_n188, u2_u3_u1_n95, u2_u3_u1_n96, u2_u3_u1_n97, u2_u3_u1_n98, u2_u3_u1_n99, 
       u2_u3_u2_n100, u2_u3_u2_n101, u2_u3_u2_n102, u2_u3_u2_n103, u2_u3_u2_n104, u2_u3_u2_n105, u2_u3_u2_n106, u2_u3_u2_n107, u2_u3_u2_n108, 
       u2_u3_u2_n109, u2_u3_u2_n110, u2_u3_u2_n111, u2_u3_u2_n112, u2_u3_u2_n113, u2_u3_u2_n114, u2_u3_u2_n115, u2_u3_u2_n116, u2_u3_u2_n117, 
       u2_u3_u2_n118, u2_u3_u2_n119, u2_u3_u2_n120, u2_u3_u2_n121, u2_u3_u2_n122, u2_u3_u2_n123, u2_u3_u2_n124, u2_u3_u2_n125, u2_u3_u2_n126, 
       u2_u3_u2_n127, u2_u3_u2_n128, u2_u3_u2_n129, u2_u3_u2_n130, u2_u3_u2_n131, u2_u3_u2_n132, u2_u3_u2_n133, u2_u3_u2_n134, u2_u3_u2_n135, 
       u2_u3_u2_n136, u2_u3_u2_n137, u2_u3_u2_n138, u2_u3_u2_n139, u2_u3_u2_n140, u2_u3_u2_n141, u2_u3_u2_n142, u2_u3_u2_n143, u2_u3_u2_n144, 
       u2_u3_u2_n145, u2_u3_u2_n146, u2_u3_u2_n147, u2_u3_u2_n148, u2_u3_u2_n149, u2_u3_u2_n150, u2_u3_u2_n151, u2_u3_u2_n152, u2_u3_u2_n153, 
       u2_u3_u2_n154, u2_u3_u2_n155, u2_u3_u2_n156, u2_u3_u2_n157, u2_u3_u2_n158, u2_u3_u2_n159, u2_u3_u2_n160, u2_u3_u2_n161, u2_u3_u2_n162, 
       u2_u3_u2_n163, u2_u3_u2_n164, u2_u3_u2_n165, u2_u3_u2_n166, u2_u3_u2_n167, u2_u3_u2_n168, u2_u3_u2_n169, u2_u3_u2_n170, u2_u3_u2_n171, 
       u2_u3_u2_n172, u2_u3_u2_n173, u2_u3_u2_n174, u2_u3_u2_n175, u2_u3_u2_n176, u2_u3_u2_n177, u2_u3_u2_n178, u2_u3_u2_n179, u2_u3_u2_n180, 
       u2_u3_u2_n181, u2_u3_u2_n182, u2_u3_u2_n183, u2_u3_u2_n184, u2_u3_u2_n185, u2_u3_u2_n186, u2_u3_u2_n187, u2_u3_u2_n188, u2_u3_u2_n95, 
       u2_u3_u2_n96, u2_u3_u2_n97, u2_u3_u2_n98, u2_u3_u2_n99, u2_u3_u3_n100, u2_u3_u3_n101, u2_u3_u3_n102, u2_u3_u3_n103, u2_u3_u3_n104, 
       u2_u3_u3_n105, u2_u3_u3_n106, u2_u3_u3_n107, u2_u3_u3_n108, u2_u3_u3_n109, u2_u3_u3_n110, u2_u3_u3_n111, u2_u3_u3_n112, u2_u3_u3_n113, 
       u2_u3_u3_n114, u2_u3_u3_n115, u2_u3_u3_n116, u2_u3_u3_n117, u2_u3_u3_n118, u2_u3_u3_n119, u2_u3_u3_n120, u2_u3_u3_n121, u2_u3_u3_n122, 
       u2_u3_u3_n123, u2_u3_u3_n124, u2_u3_u3_n125, u2_u3_u3_n126, u2_u3_u3_n127, u2_u3_u3_n128, u2_u3_u3_n129, u2_u3_u3_n130, u2_u3_u3_n131, 
       u2_u3_u3_n132, u2_u3_u3_n133, u2_u3_u3_n134, u2_u3_u3_n135, u2_u3_u3_n136, u2_u3_u3_n137, u2_u3_u3_n138, u2_u3_u3_n139, u2_u3_u3_n140, 
       u2_u3_u3_n141, u2_u3_u3_n142, u2_u3_u3_n143, u2_u3_u3_n144, u2_u3_u3_n145, u2_u3_u3_n146, u2_u3_u3_n147, u2_u3_u3_n148, u2_u3_u3_n149, 
       u2_u3_u3_n150, u2_u3_u3_n151, u2_u3_u3_n152, u2_u3_u3_n153, u2_u3_u3_n154, u2_u3_u3_n155, u2_u3_u3_n156, u2_u3_u3_n157, u2_u3_u3_n158, 
       u2_u3_u3_n159, u2_u3_u3_n160, u2_u3_u3_n161, u2_u3_u3_n162, u2_u3_u3_n163, u2_u3_u3_n164, u2_u3_u3_n165, u2_u3_u3_n166, u2_u3_u3_n167, 
       u2_u3_u3_n168, u2_u3_u3_n169, u2_u3_u3_n170, u2_u3_u3_n171, u2_u3_u3_n172, u2_u3_u3_n173, u2_u3_u3_n174, u2_u3_u3_n175, u2_u3_u3_n176, 
       u2_u3_u3_n177, u2_u3_u3_n178, u2_u3_u3_n179, u2_u3_u3_n180, u2_u3_u3_n181, u2_u3_u3_n182, u2_u3_u3_n183, u2_u3_u3_n184, u2_u3_u3_n185, 
       u2_u3_u3_n186, u2_u3_u3_n94, u2_u3_u3_n95, u2_u3_u3_n96, u2_u3_u3_n97, u2_u3_u3_n98, u2_u3_u3_n99, u2_u3_u4_n100, u2_u3_u4_n101, 
       u2_u3_u4_n102, u2_u3_u4_n103, u2_u3_u4_n104, u2_u3_u4_n105, u2_u3_u4_n106, u2_u3_u4_n107, u2_u3_u4_n108, u2_u3_u4_n109, u2_u3_u4_n110, 
       u2_u3_u4_n111, u2_u3_u4_n112, u2_u3_u4_n113, u2_u3_u4_n114, u2_u3_u4_n115, u2_u3_u4_n116, u2_u3_u4_n117, u2_u3_u4_n118, u2_u3_u4_n119, 
       u2_u3_u4_n120, u2_u3_u4_n121, u2_u3_u4_n122, u2_u3_u4_n123, u2_u3_u4_n124, u2_u3_u4_n125, u2_u3_u4_n126, u2_u3_u4_n127, u2_u3_u4_n128, 
       u2_u3_u4_n129, u2_u3_u4_n130, u2_u3_u4_n131, u2_u3_u4_n132, u2_u3_u4_n133, u2_u3_u4_n134, u2_u3_u4_n135, u2_u3_u4_n136, u2_u3_u4_n137, 
       u2_u3_u4_n138, u2_u3_u4_n139, u2_u3_u4_n140, u2_u3_u4_n141, u2_u3_u4_n142, u2_u3_u4_n143, u2_u3_u4_n144, u2_u3_u4_n145, u2_u3_u4_n146, 
       u2_u3_u4_n147, u2_u3_u4_n148, u2_u3_u4_n149, u2_u3_u4_n150, u2_u3_u4_n151, u2_u3_u4_n152, u2_u3_u4_n153, u2_u3_u4_n154, u2_u3_u4_n155, 
       u2_u3_u4_n156, u2_u3_u4_n157, u2_u3_u4_n158, u2_u3_u4_n159, u2_u3_u4_n160, u2_u3_u4_n161, u2_u3_u4_n162, u2_u3_u4_n163, u2_u3_u4_n164, 
       u2_u3_u4_n165, u2_u3_u4_n166, u2_u3_u4_n167, u2_u3_u4_n168, u2_u3_u4_n169, u2_u3_u4_n170, u2_u3_u4_n171, u2_u3_u4_n172, u2_u3_u4_n173, 
       u2_u3_u4_n174, u2_u3_u4_n175, u2_u3_u4_n176, u2_u3_u4_n177, u2_u3_u4_n178, u2_u3_u4_n179, u2_u3_u4_n180, u2_u3_u4_n181, u2_u3_u4_n182, 
       u2_u3_u4_n183, u2_u3_u4_n184, u2_u3_u4_n185, u2_u3_u4_n186, u2_u3_u4_n94, u2_u3_u4_n95, u2_u3_u4_n96, u2_u3_u4_n97, u2_u3_u4_n98, 
       u2_u3_u4_n99, u2_u3_u5_n100, u2_u3_u5_n101, u2_u3_u5_n102, u2_u3_u5_n103, u2_u3_u5_n104, u2_u3_u5_n105, u2_u3_u5_n106, u2_u3_u5_n107, 
       u2_u3_u5_n108, u2_u3_u5_n109, u2_u3_u5_n110, u2_u3_u5_n111, u2_u3_u5_n112, u2_u3_u5_n113, u2_u3_u5_n114, u2_u3_u5_n115, u2_u3_u5_n116, 
       u2_u3_u5_n117, u2_u3_u5_n118, u2_u3_u5_n119, u2_u3_u5_n120, u2_u3_u5_n121, u2_u3_u5_n122, u2_u3_u5_n123, u2_u3_u5_n124, u2_u3_u5_n125, 
       u2_u3_u5_n126, u2_u3_u5_n127, u2_u3_u5_n128, u2_u3_u5_n129, u2_u3_u5_n130, u2_u3_u5_n131, u2_u3_u5_n132, u2_u3_u5_n133, u2_u3_u5_n134, 
       u2_u3_u5_n135, u2_u3_u5_n136, u2_u3_u5_n137, u2_u3_u5_n138, u2_u3_u5_n139, u2_u3_u5_n140, u2_u3_u5_n141, u2_u3_u5_n142, u2_u3_u5_n143, 
       u2_u3_u5_n144, u2_u3_u5_n145, u2_u3_u5_n146, u2_u3_u5_n147, u2_u3_u5_n148, u2_u3_u5_n149, u2_u3_u5_n150, u2_u3_u5_n151, u2_u3_u5_n152, 
       u2_u3_u5_n153, u2_u3_u5_n154, u2_u3_u5_n155, u2_u3_u5_n156, u2_u3_u5_n157, u2_u3_u5_n158, u2_u3_u5_n159, u2_u3_u5_n160, u2_u3_u5_n161, 
       u2_u3_u5_n162, u2_u3_u5_n163, u2_u3_u5_n164, u2_u3_u5_n165, u2_u3_u5_n166, u2_u3_u5_n167, u2_u3_u5_n168, u2_u3_u5_n169, u2_u3_u5_n170, 
       u2_u3_u5_n171, u2_u3_u5_n172, u2_u3_u5_n173, u2_u3_u5_n174, u2_u3_u5_n175, u2_u3_u5_n176, u2_u3_u5_n177, u2_u3_u5_n178, u2_u3_u5_n179, 
       u2_u3_u5_n180, u2_u3_u5_n181, u2_u3_u5_n182, u2_u3_u5_n183, u2_u3_u5_n184, u2_u3_u5_n185, u2_u3_u5_n186, u2_u3_u5_n187, u2_u3_u5_n188, 
       u2_u3_u5_n189, u2_u3_u5_n190, u2_u3_u5_n191, u2_u3_u5_n192, u2_u3_u5_n193, u2_u3_u5_n194, u2_u3_u5_n195, u2_u3_u5_n196, u2_u3_u5_n99, 
       u2_u3_u7_n100, u2_u3_u7_n101, u2_u3_u7_n102, u2_u3_u7_n103, u2_u3_u7_n104, u2_u3_u7_n105, u2_u3_u7_n106, u2_u3_u7_n107, u2_u3_u7_n108, 
       u2_u3_u7_n109, u2_u3_u7_n110, u2_u3_u7_n111, u2_u3_u7_n112, u2_u3_u7_n113, u2_u3_u7_n114, u2_u3_u7_n115, u2_u3_u7_n116, u2_u3_u7_n117, 
       u2_u3_u7_n118, u2_u3_u7_n119, u2_u3_u7_n120, u2_u3_u7_n121, u2_u3_u7_n122, u2_u3_u7_n123, u2_u3_u7_n124, u2_u3_u7_n125, u2_u3_u7_n126, 
       u2_u3_u7_n127, u2_u3_u7_n128, u2_u3_u7_n129, u2_u3_u7_n130, u2_u3_u7_n131, u2_u3_u7_n132, u2_u3_u7_n133, u2_u3_u7_n134, u2_u3_u7_n135, 
       u2_u3_u7_n136, u2_u3_u7_n137, u2_u3_u7_n138, u2_u3_u7_n139, u2_u3_u7_n140, u2_u3_u7_n141, u2_u3_u7_n142, u2_u3_u7_n143, u2_u3_u7_n144, 
       u2_u3_u7_n145, u2_u3_u7_n146, u2_u3_u7_n147, u2_u3_u7_n148, u2_u3_u7_n149, u2_u3_u7_n150, u2_u3_u7_n151, u2_u3_u7_n152, u2_u3_u7_n153, 
       u2_u3_u7_n154, u2_u3_u7_n155, u2_u3_u7_n156, u2_u3_u7_n157, u2_u3_u7_n158, u2_u3_u7_n159, u2_u3_u7_n160, u2_u3_u7_n161, u2_u3_u7_n162, 
       u2_u3_u7_n163, u2_u3_u7_n164, u2_u3_u7_n165, u2_u3_u7_n166, u2_u3_u7_n167, u2_u3_u7_n168, u2_u3_u7_n169, u2_u3_u7_n170, u2_u3_u7_n171, 
       u2_u3_u7_n172, u2_u3_u7_n173, u2_u3_u7_n174, u2_u3_u7_n175, u2_u3_u7_n176, u2_u3_u7_n177, u2_u3_u7_n178, u2_u3_u7_n179, u2_u3_u7_n180, 
       u2_u3_u7_n91, u2_u3_u7_n92, u2_u3_u7_n93, u2_u3_u7_n94, u2_u3_u7_n95, u2_u3_u7_n96, u2_u3_u7_n97, u2_u3_u7_n98, u2_u3_u7_n99, 
       u2_u4_X_11, u2_u4_X_12, u2_u4_X_13, u2_u4_X_14, u2_u4_X_17, u2_u4_X_18, u2_u4_X_19, u2_u4_X_2, u2_u4_X_20, 
       u2_u4_X_23, u2_u4_X_24, u2_u4_X_25, u2_u4_X_26, u2_u4_X_27, u2_u4_X_29, u2_u4_X_30, u2_u4_X_31, u2_u4_X_32, 
       u2_u4_X_33, u2_u4_X_35, u2_u4_X_36, u2_u4_X_37, u2_u4_X_38, u2_u4_X_41, u2_u4_X_42, u2_u4_X_43, u2_u4_X_44, 
       u2_u4_X_45, u2_u4_X_48, u2_u4_X_5, u2_u4_X_6, u2_u4_X_7, u2_u4_X_8, u2_u4_u0_n100, u2_u4_u0_n101, u2_u4_u0_n102, 
       u2_u4_u0_n103, u2_u4_u0_n104, u2_u4_u0_n105, u2_u4_u0_n106, u2_u4_u0_n107, u2_u4_u0_n108, u2_u4_u0_n109, u2_u4_u0_n110, u2_u4_u0_n111, 
       u2_u4_u0_n112, u2_u4_u0_n113, u2_u4_u0_n114, u2_u4_u0_n115, u2_u4_u0_n116, u2_u4_u0_n117, u2_u4_u0_n118, u2_u4_u0_n119, u2_u4_u0_n120, 
       u2_u4_u0_n121, u2_u4_u0_n122, u2_u4_u0_n123, u2_u4_u0_n124, u2_u4_u0_n125, u2_u4_u0_n126, u2_u4_u0_n127, u2_u4_u0_n128, u2_u4_u0_n129, 
       u2_u4_u0_n130, u2_u4_u0_n131, u2_u4_u0_n132, u2_u4_u0_n133, u2_u4_u0_n134, u2_u4_u0_n135, u2_u4_u0_n136, u2_u4_u0_n137, u2_u4_u0_n138, 
       u2_u4_u0_n139, u2_u4_u0_n140, u2_u4_u0_n141, u2_u4_u0_n142, u2_u4_u0_n143, u2_u4_u0_n144, u2_u4_u0_n145, u2_u4_u0_n146, u2_u4_u0_n147, 
       u2_u4_u0_n148, u2_u4_u0_n149, u2_u4_u0_n150, u2_u4_u0_n151, u2_u4_u0_n152, u2_u4_u0_n153, u2_u4_u0_n154, u2_u4_u0_n155, u2_u4_u0_n156, 
       u2_u4_u0_n157, u2_u4_u0_n158, u2_u4_u0_n159, u2_u4_u0_n160, u2_u4_u0_n161, u2_u4_u0_n162, u2_u4_u0_n163, u2_u4_u0_n164, u2_u4_u0_n165, 
       u2_u4_u0_n166, u2_u4_u0_n167, u2_u4_u0_n168, u2_u4_u0_n169, u2_u4_u0_n170, u2_u4_u0_n171, u2_u4_u0_n172, u2_u4_u0_n173, u2_u4_u0_n174, 
       u2_u4_u0_n88, u2_u4_u0_n89, u2_u4_u0_n90, u2_u4_u0_n91, u2_u4_u0_n92, u2_u4_u0_n93, u2_u4_u0_n94, u2_u4_u0_n95, u2_u4_u0_n96, 
       u2_u4_u0_n97, u2_u4_u0_n98, u2_u4_u0_n99, u2_u4_u1_n100, u2_u4_u1_n101, u2_u4_u1_n102, u2_u4_u1_n103, u2_u4_u1_n104, u2_u4_u1_n105, 
       u2_u4_u1_n106, u2_u4_u1_n107, u2_u4_u1_n108, u2_u4_u1_n109, u2_u4_u1_n110, u2_u4_u1_n111, u2_u4_u1_n112, u2_u4_u1_n113, u2_u4_u1_n114, 
       u2_u4_u1_n115, u2_u4_u1_n116, u2_u4_u1_n117, u2_u4_u1_n118, u2_u4_u1_n119, u2_u4_u1_n120, u2_u4_u1_n121, u2_u4_u1_n122, u2_u4_u1_n123, 
       u2_u4_u1_n124, u2_u4_u1_n125, u2_u4_u1_n126, u2_u4_u1_n127, u2_u4_u1_n128, u2_u4_u1_n129, u2_u4_u1_n130, u2_u4_u1_n131, u2_u4_u1_n132, 
       u2_u4_u1_n133, u2_u4_u1_n134, u2_u4_u1_n135, u2_u4_u1_n136, u2_u4_u1_n137, u2_u4_u1_n138, u2_u4_u1_n139, u2_u4_u1_n140, u2_u4_u1_n141, 
       u2_u4_u1_n142, u2_u4_u1_n143, u2_u4_u1_n144, u2_u4_u1_n145, u2_u4_u1_n146, u2_u4_u1_n147, u2_u4_u1_n148, u2_u4_u1_n149, u2_u4_u1_n150, 
       u2_u4_u1_n151, u2_u4_u1_n152, u2_u4_u1_n153, u2_u4_u1_n154, u2_u4_u1_n155, u2_u4_u1_n156, u2_u4_u1_n157, u2_u4_u1_n158, u2_u4_u1_n159, 
       u2_u4_u1_n160, u2_u4_u1_n161, u2_u4_u1_n162, u2_u4_u1_n163, u2_u4_u1_n164, u2_u4_u1_n165, u2_u4_u1_n166, u2_u4_u1_n167, u2_u4_u1_n168, 
       u2_u4_u1_n169, u2_u4_u1_n170, u2_u4_u1_n171, u2_u4_u1_n172, u2_u4_u1_n173, u2_u4_u1_n174, u2_u4_u1_n175, u2_u4_u1_n176, u2_u4_u1_n177, 
       u2_u4_u1_n178, u2_u4_u1_n179, u2_u4_u1_n180, u2_u4_u1_n181, u2_u4_u1_n182, u2_u4_u1_n183, u2_u4_u1_n184, u2_u4_u1_n185, u2_u4_u1_n186, 
       u2_u4_u1_n187, u2_u4_u1_n188, u2_u4_u1_n95, u2_u4_u1_n96, u2_u4_u1_n97, u2_u4_u1_n98, u2_u4_u1_n99, u2_u4_u2_n100, u2_u4_u2_n101, 
       u2_u4_u2_n102, u2_u4_u2_n103, u2_u4_u2_n104, u2_u4_u2_n105, u2_u4_u2_n106, u2_u4_u2_n107, u2_u4_u2_n108, u2_u4_u2_n109, u2_u4_u2_n110, 
       u2_u4_u2_n111, u2_u4_u2_n112, u2_u4_u2_n113, u2_u4_u2_n114, u2_u4_u2_n115, u2_u4_u2_n116, u2_u4_u2_n117, u2_u4_u2_n118, u2_u4_u2_n119, 
       u2_u4_u2_n120, u2_u4_u2_n121, u2_u4_u2_n122, u2_u4_u2_n123, u2_u4_u2_n124, u2_u4_u2_n125, u2_u4_u2_n126, u2_u4_u2_n127, u2_u4_u2_n128, 
       u2_u4_u2_n129, u2_u4_u2_n130, u2_u4_u2_n131, u2_u4_u2_n132, u2_u4_u2_n133, u2_u4_u2_n134, u2_u4_u2_n135, u2_u4_u2_n136, u2_u4_u2_n137, 
       u2_u4_u2_n138, u2_u4_u2_n139, u2_u4_u2_n140, u2_u4_u2_n141, u2_u4_u2_n142, u2_u4_u2_n143, u2_u4_u2_n144, u2_u4_u2_n145, u2_u4_u2_n146, 
       u2_u4_u2_n147, u2_u4_u2_n148, u2_u4_u2_n149, u2_u4_u2_n150, u2_u4_u2_n151, u2_u4_u2_n152, u2_u4_u2_n153, u2_u4_u2_n154, u2_u4_u2_n155, 
       u2_u4_u2_n156, u2_u4_u2_n157, u2_u4_u2_n158, u2_u4_u2_n159, u2_u4_u2_n160, u2_u4_u2_n161, u2_u4_u2_n162, u2_u4_u2_n163, u2_u4_u2_n164, 
       u2_u4_u2_n165, u2_u4_u2_n166, u2_u4_u2_n167, u2_u4_u2_n168, u2_u4_u2_n169, u2_u4_u2_n170, u2_u4_u2_n171, u2_u4_u2_n172, u2_u4_u2_n173, 
       u2_u4_u2_n174, u2_u4_u2_n175, u2_u4_u2_n176, u2_u4_u2_n177, u2_u4_u2_n178, u2_u4_u2_n179, u2_u4_u2_n180, u2_u4_u2_n181, u2_u4_u2_n182, 
       u2_u4_u2_n183, u2_u4_u2_n184, u2_u4_u2_n185, u2_u4_u2_n186, u2_u4_u2_n187, u2_u4_u2_n188, u2_u4_u2_n95, u2_u4_u2_n96, u2_u4_u2_n97, 
       u2_u4_u2_n98, u2_u4_u2_n99, u2_u4_u3_n100, u2_u4_u3_n101, u2_u4_u3_n102, u2_u4_u3_n103, u2_u4_u3_n104, u2_u4_u3_n105, u2_u4_u3_n106, 
       u2_u4_u3_n107, u2_u4_u3_n108, u2_u4_u3_n109, u2_u4_u3_n110, u2_u4_u3_n111, u2_u4_u3_n112, u2_u4_u3_n113, u2_u4_u3_n114, u2_u4_u3_n115, 
       u2_u4_u3_n116, u2_u4_u3_n117, u2_u4_u3_n118, u2_u4_u3_n119, u2_u4_u3_n120, u2_u4_u3_n121, u2_u4_u3_n122, u2_u4_u3_n123, u2_u4_u3_n124, 
       u2_u4_u3_n125, u2_u4_u3_n126, u2_u4_u3_n127, u2_u4_u3_n128, u2_u4_u3_n129, u2_u4_u3_n130, u2_u4_u3_n131, u2_u4_u3_n132, u2_u4_u3_n133, 
       u2_u4_u3_n134, u2_u4_u3_n135, u2_u4_u3_n136, u2_u4_u3_n137, u2_u4_u3_n138, u2_u4_u3_n139, u2_u4_u3_n140, u2_u4_u3_n141, u2_u4_u3_n142, 
       u2_u4_u3_n143, u2_u4_u3_n144, u2_u4_u3_n145, u2_u4_u3_n146, u2_u4_u3_n147, u2_u4_u3_n148, u2_u4_u3_n149, u2_u4_u3_n150, u2_u4_u3_n151, 
       u2_u4_u3_n152, u2_u4_u3_n153, u2_u4_u3_n154, u2_u4_u3_n155, u2_u4_u3_n156, u2_u4_u3_n157, u2_u4_u3_n158, u2_u4_u3_n159, u2_u4_u3_n160, 
       u2_u4_u3_n161, u2_u4_u3_n162, u2_u4_u3_n163, u2_u4_u3_n164, u2_u4_u3_n165, u2_u4_u3_n166, u2_u4_u3_n167, u2_u4_u3_n168, u2_u4_u3_n169, 
       u2_u4_u3_n170, u2_u4_u3_n171, u2_u4_u3_n172, u2_u4_u3_n173, u2_u4_u3_n174, u2_u4_u3_n175, u2_u4_u3_n176, u2_u4_u3_n177, u2_u4_u3_n178, 
       u2_u4_u3_n179, u2_u4_u3_n180, u2_u4_u3_n181, u2_u4_u3_n182, u2_u4_u3_n183, u2_u4_u3_n184, u2_u4_u3_n185, u2_u4_u3_n186, u2_u4_u3_n94, 
       u2_u4_u3_n95, u2_u4_u3_n96, u2_u4_u3_n97, u2_u4_u3_n98, u2_u4_u3_n99, u2_u4_u4_n100, u2_u4_u4_n101, u2_u4_u4_n102, u2_u4_u4_n103, 
       u2_u4_u4_n104, u2_u4_u4_n105, u2_u4_u4_n106, u2_u4_u4_n107, u2_u4_u4_n108, u2_u4_u4_n109, u2_u4_u4_n110, u2_u4_u4_n111, u2_u4_u4_n112, 
       u2_u4_u4_n113, u2_u4_u4_n114, u2_u4_u4_n115, u2_u4_u4_n116, u2_u4_u4_n117, u2_u4_u4_n118, u2_u4_u4_n119, u2_u4_u4_n120, u2_u4_u4_n121, 
       u2_u4_u4_n122, u2_u4_u4_n123, u2_u4_u4_n124, u2_u4_u4_n125, u2_u4_u4_n126, u2_u4_u4_n127, u2_u4_u4_n128, u2_u4_u4_n129, u2_u4_u4_n130, 
       u2_u4_u4_n131, u2_u4_u4_n132, u2_u4_u4_n133, u2_u4_u4_n134, u2_u4_u4_n135, u2_u4_u4_n136, u2_u4_u4_n137, u2_u4_u4_n138, u2_u4_u4_n139, 
       u2_u4_u4_n140, u2_u4_u4_n141, u2_u4_u4_n142, u2_u4_u4_n143, u2_u4_u4_n144, u2_u4_u4_n145, u2_u4_u4_n146, u2_u4_u4_n147, u2_u4_u4_n148, 
       u2_u4_u4_n149, u2_u4_u4_n150, u2_u4_u4_n151, u2_u4_u4_n152, u2_u4_u4_n153, u2_u4_u4_n154, u2_u4_u4_n155, u2_u4_u4_n156, u2_u4_u4_n157, 
       u2_u4_u4_n158, u2_u4_u4_n159, u2_u4_u4_n160, u2_u4_u4_n161, u2_u4_u4_n162, u2_u4_u4_n163, u2_u4_u4_n164, u2_u4_u4_n165, u2_u4_u4_n166, 
       u2_u4_u4_n167, u2_u4_u4_n168, u2_u4_u4_n169, u2_u4_u4_n170, u2_u4_u4_n171, u2_u4_u4_n172, u2_u4_u4_n173, u2_u4_u4_n174, u2_u4_u4_n175, 
       u2_u4_u4_n176, u2_u4_u4_n177, u2_u4_u4_n178, u2_u4_u4_n179, u2_u4_u4_n180, u2_u4_u4_n181, u2_u4_u4_n182, u2_u4_u4_n183, u2_u4_u4_n184, 
       u2_u4_u4_n185, u2_u4_u4_n186, u2_u4_u4_n94, u2_u4_u4_n95, u2_u4_u4_n96, u2_u4_u4_n97, u2_u4_u4_n98, u2_u4_u4_n99, u2_u4_u5_n100, 
       u2_u4_u5_n101, u2_u4_u5_n102, u2_u4_u5_n103, u2_u4_u5_n104, u2_u4_u5_n105, u2_u4_u5_n106, u2_u4_u5_n107, u2_u4_u5_n108, u2_u4_u5_n109, 
       u2_u4_u5_n110, u2_u4_u5_n111, u2_u4_u5_n112, u2_u4_u5_n113, u2_u4_u5_n114, u2_u4_u5_n115, u2_u4_u5_n116, u2_u4_u5_n117, u2_u4_u5_n118, 
       u2_u4_u5_n119, u2_u4_u5_n120, u2_u4_u5_n121, u2_u4_u5_n122, u2_u4_u5_n123, u2_u4_u5_n124, u2_u4_u5_n125, u2_u4_u5_n126, u2_u4_u5_n127, 
       u2_u4_u5_n128, u2_u4_u5_n129, u2_u4_u5_n130, u2_u4_u5_n131, u2_u4_u5_n132, u2_u4_u5_n133, u2_u4_u5_n134, u2_u4_u5_n135, u2_u4_u5_n136, 
       u2_u4_u5_n137, u2_u4_u5_n138, u2_u4_u5_n139, u2_u4_u5_n140, u2_u4_u5_n141, u2_u4_u5_n142, u2_u4_u5_n143, u2_u4_u5_n144, u2_u4_u5_n145, 
       u2_u4_u5_n146, u2_u4_u5_n147, u2_u4_u5_n148, u2_u4_u5_n149, u2_u4_u5_n150, u2_u4_u5_n151, u2_u4_u5_n152, u2_u4_u5_n153, u2_u4_u5_n154, 
       u2_u4_u5_n155, u2_u4_u5_n156, u2_u4_u5_n157, u2_u4_u5_n158, u2_u4_u5_n159, u2_u4_u5_n160, u2_u4_u5_n161, u2_u4_u5_n162, u2_u4_u5_n163, 
       u2_u4_u5_n164, u2_u4_u5_n165, u2_u4_u5_n166, u2_u4_u5_n167, u2_u4_u5_n168, u2_u4_u5_n169, u2_u4_u5_n170, u2_u4_u5_n171, u2_u4_u5_n172, 
       u2_u4_u5_n173, u2_u4_u5_n174, u2_u4_u5_n175, u2_u4_u5_n176, u2_u4_u5_n177, u2_u4_u5_n178, u2_u4_u5_n179, u2_u4_u5_n180, u2_u4_u5_n181, 
       u2_u4_u5_n182, u2_u4_u5_n183, u2_u4_u5_n184, u2_u4_u5_n185, u2_u4_u5_n186, u2_u4_u5_n187, u2_u4_u5_n188, u2_u4_u5_n189, u2_u4_u5_n190, 
       u2_u4_u5_n191, u2_u4_u5_n192, u2_u4_u5_n193, u2_u4_u5_n194, u2_u4_u5_n195, u2_u4_u5_n196, u2_u4_u5_n99, u2_u4_u6_n100, u2_u4_u6_n101, 
       u2_u4_u6_n102, u2_u4_u6_n103, u2_u4_u6_n104, u2_u4_u6_n105, u2_u4_u6_n106, u2_u4_u6_n107, u2_u4_u6_n108, u2_u4_u6_n109, u2_u4_u6_n110, 
       u2_u4_u6_n111, u2_u4_u6_n112, u2_u4_u6_n113, u2_u4_u6_n114, u2_u4_u6_n115, u2_u4_u6_n116, u2_u4_u6_n117, u2_u4_u6_n118, u2_u4_u6_n119, 
       u2_u4_u6_n120, u2_u4_u6_n121, u2_u4_u6_n122, u2_u4_u6_n123, u2_u4_u6_n124, u2_u4_u6_n125, u2_u4_u6_n126, u2_u4_u6_n127, u2_u4_u6_n128, 
       u2_u4_u6_n129, u2_u4_u6_n130, u2_u4_u6_n131, u2_u4_u6_n132, u2_u4_u6_n133, u2_u4_u6_n134, u2_u4_u6_n135, u2_u4_u6_n136, u2_u4_u6_n137, 
       u2_u4_u6_n138, u2_u4_u6_n139, u2_u4_u6_n140, u2_u4_u6_n141, u2_u4_u6_n142, u2_u4_u6_n143, u2_u4_u6_n144, u2_u4_u6_n145, u2_u4_u6_n146, 
       u2_u4_u6_n147, u2_u4_u6_n148, u2_u4_u6_n149, u2_u4_u6_n150, u2_u4_u6_n151, u2_u4_u6_n152, u2_u4_u6_n153, u2_u4_u6_n154, u2_u4_u6_n155, 
       u2_u4_u6_n156, u2_u4_u6_n157, u2_u4_u6_n158, u2_u4_u6_n159, u2_u4_u6_n160, u2_u4_u6_n161, u2_u4_u6_n162, u2_u4_u6_n163, u2_u4_u6_n164, 
       u2_u4_u6_n165, u2_u4_u6_n166, u2_u4_u6_n167, u2_u4_u6_n168, u2_u4_u6_n169, u2_u4_u6_n170, u2_u4_u6_n171, u2_u4_u6_n172, u2_u4_u6_n173, 
       u2_u4_u6_n174, u2_u4_u6_n88, u2_u4_u6_n89, u2_u4_u6_n90, u2_u4_u6_n91, u2_u4_u6_n92, u2_u4_u6_n93, u2_u4_u6_n94, u2_u4_u6_n95, 
       u2_u4_u6_n96, u2_u4_u6_n97, u2_u4_u6_n98, u2_u4_u6_n99, u2_u4_u7_n100, u2_u4_u7_n101, u2_u4_u7_n102, u2_u4_u7_n103, u2_u4_u7_n104, 
       u2_u4_u7_n105, u2_u4_u7_n106, u2_u4_u7_n107, u2_u4_u7_n108, u2_u4_u7_n109, u2_u4_u7_n110, u2_u4_u7_n111, u2_u4_u7_n112, u2_u4_u7_n113, 
       u2_u4_u7_n114, u2_u4_u7_n115, u2_u4_u7_n116, u2_u4_u7_n117, u2_u4_u7_n118, u2_u4_u7_n119, u2_u4_u7_n120, u2_u4_u7_n121, u2_u4_u7_n122, 
       u2_u4_u7_n123, u2_u4_u7_n124, u2_u4_u7_n125, u2_u4_u7_n126, u2_u4_u7_n127, u2_u4_u7_n128, u2_u4_u7_n129, u2_u4_u7_n130, u2_u4_u7_n131, 
       u2_u4_u7_n132, u2_u4_u7_n133, u2_u4_u7_n134, u2_u4_u7_n135, u2_u4_u7_n136, u2_u4_u7_n137, u2_u4_u7_n138, u2_u4_u7_n139, u2_u4_u7_n140, 
       u2_u4_u7_n141, u2_u4_u7_n142, u2_u4_u7_n143, u2_u4_u7_n144, u2_u4_u7_n145, u2_u4_u7_n146, u2_u4_u7_n147, u2_u4_u7_n148, u2_u4_u7_n149, 
       u2_u4_u7_n150, u2_u4_u7_n151, u2_u4_u7_n152, u2_u4_u7_n153, u2_u4_u7_n154, u2_u4_u7_n155, u2_u4_u7_n156, u2_u4_u7_n157, u2_u4_u7_n158, 
       u2_u4_u7_n159, u2_u4_u7_n160, u2_u4_u7_n161, u2_u4_u7_n162, u2_u4_u7_n163, u2_u4_u7_n164, u2_u4_u7_n165, u2_u4_u7_n166, u2_u4_u7_n167, 
       u2_u4_u7_n168, u2_u4_u7_n169, u2_u4_u7_n170, u2_u4_u7_n171, u2_u4_u7_n172, u2_u4_u7_n173, u2_u4_u7_n174, u2_u4_u7_n175, u2_u4_u7_n176, 
       u2_u4_u7_n177, u2_u4_u7_n178, u2_u4_u7_n179, u2_u4_u7_n180, u2_u4_u7_n91, u2_u4_u7_n92, u2_u4_u7_n93, u2_u4_u7_n94, u2_u4_u7_n95, 
       u2_u4_u7_n96, u2_u4_u7_n97, u2_u4_u7_n98, u2_u4_u7_n99, u2_u5_X_1, u2_u5_X_11, u2_u5_X_12, u2_u5_X_13, u2_u5_X_14, 
       u2_u5_X_17, u2_u5_X_18, u2_u5_X_19, u2_u5_X_2, u2_u5_X_20, u2_u5_X_21, u2_u5_X_24, u2_u5_X_26, u2_u5_X_30, 
       u2_u5_X_32, u2_u5_X_33, u2_u5_X_35, u2_u5_X_37, u2_u5_X_41, u2_u5_X_42, u2_u5_X_43, u2_u5_X_44, u2_u5_X_46, 
       u2_u5_X_47, u2_u5_X_48, u2_u5_X_5, u2_u5_X_6, u2_u5_X_7, u2_u5_X_8, u2_u5_X_9, u2_u5_u0_n100, u2_u5_u0_n101, 
       u2_u5_u0_n102, u2_u5_u0_n103, u2_u5_u0_n104, u2_u5_u0_n105, u2_u5_u0_n106, u2_u5_u0_n107, u2_u5_u0_n108, u2_u5_u0_n109, u2_u5_u0_n110, 
       u2_u5_u0_n111, u2_u5_u0_n112, u2_u5_u0_n113, u2_u5_u0_n114, u2_u5_u0_n115, u2_u5_u0_n116, u2_u5_u0_n117, u2_u5_u0_n118, u2_u5_u0_n119, 
       u2_u5_u0_n120, u2_u5_u0_n121, u2_u5_u0_n122, u2_u5_u0_n123, u2_u5_u0_n124, u2_u5_u0_n125, u2_u5_u0_n126, u2_u5_u0_n127, u2_u5_u0_n128, 
       u2_u5_u0_n129, u2_u5_u0_n130, u2_u5_u0_n131, u2_u5_u0_n132, u2_u5_u0_n133, u2_u5_u0_n134, u2_u5_u0_n135, u2_u5_u0_n136, u2_u5_u0_n137, 
       u2_u5_u0_n138, u2_u5_u0_n139, u2_u5_u0_n140, u2_u5_u0_n141, u2_u5_u0_n142, u2_u5_u0_n143, u2_u5_u0_n144, u2_u5_u0_n145, u2_u5_u0_n146, 
       u2_u5_u0_n147, u2_u5_u0_n148, u2_u5_u0_n149, u2_u5_u0_n150, u2_u5_u0_n151, u2_u5_u0_n152, u2_u5_u0_n153, u2_u5_u0_n154, u2_u5_u0_n155, 
       u2_u5_u0_n156, u2_u5_u0_n157, u2_u5_u0_n158, u2_u5_u0_n159, u2_u5_u0_n160, u2_u5_u0_n161, u2_u5_u0_n162, u2_u5_u0_n163, u2_u5_u0_n164, 
       u2_u5_u0_n165, u2_u5_u0_n166, u2_u5_u0_n167, u2_u5_u0_n168, u2_u5_u0_n169, u2_u5_u0_n170, u2_u5_u0_n171, u2_u5_u0_n172, u2_u5_u0_n173, 
       u2_u5_u0_n174, u2_u5_u0_n88, u2_u5_u0_n89, u2_u5_u0_n90, u2_u5_u0_n91, u2_u5_u0_n92, u2_u5_u0_n93, u2_u5_u0_n94, u2_u5_u0_n95, 
       u2_u5_u0_n96, u2_u5_u0_n97, u2_u5_u0_n98, u2_u5_u0_n99, u2_u5_u1_n100, u2_u5_u1_n101, u2_u5_u1_n102, u2_u5_u1_n103, u2_u5_u1_n104, 
       u2_u5_u1_n105, u2_u5_u1_n106, u2_u5_u1_n107, u2_u5_u1_n108, u2_u5_u1_n109, u2_u5_u1_n110, u2_u5_u1_n111, u2_u5_u1_n112, u2_u5_u1_n113, 
       u2_u5_u1_n114, u2_u5_u1_n115, u2_u5_u1_n116, u2_u5_u1_n117, u2_u5_u1_n118, u2_u5_u1_n119, u2_u5_u1_n120, u2_u5_u1_n121, u2_u5_u1_n122, 
       u2_u5_u1_n123, u2_u5_u1_n124, u2_u5_u1_n125, u2_u5_u1_n126, u2_u5_u1_n127, u2_u5_u1_n128, u2_u5_u1_n129, u2_u5_u1_n130, u2_u5_u1_n131, 
       u2_u5_u1_n132, u2_u5_u1_n133, u2_u5_u1_n134, u2_u5_u1_n135, u2_u5_u1_n136, u2_u5_u1_n137, u2_u5_u1_n138, u2_u5_u1_n139, u2_u5_u1_n140, 
       u2_u5_u1_n141, u2_u5_u1_n142, u2_u5_u1_n143, u2_u5_u1_n144, u2_u5_u1_n145, u2_u5_u1_n146, u2_u5_u1_n147, u2_u5_u1_n148, u2_u5_u1_n149, 
       u2_u5_u1_n150, u2_u5_u1_n151, u2_u5_u1_n152, u2_u5_u1_n153, u2_u5_u1_n154, u2_u5_u1_n155, u2_u5_u1_n156, u2_u5_u1_n157, u2_u5_u1_n158, 
       u2_u5_u1_n159, u2_u5_u1_n160, u2_u5_u1_n161, u2_u5_u1_n162, u2_u5_u1_n163, u2_u5_u1_n164, u2_u5_u1_n165, u2_u5_u1_n166, u2_u5_u1_n167, 
       u2_u5_u1_n168, u2_u5_u1_n169, u2_u5_u1_n170, u2_u5_u1_n171, u2_u5_u1_n172, u2_u5_u1_n173, u2_u5_u1_n174, u2_u5_u1_n175, u2_u5_u1_n176, 
       u2_u5_u1_n177, u2_u5_u1_n178, u2_u5_u1_n179, u2_u5_u1_n180, u2_u5_u1_n181, u2_u5_u1_n182, u2_u5_u1_n183, u2_u5_u1_n184, u2_u5_u1_n185, 
       u2_u5_u1_n186, u2_u5_u1_n187, u2_u5_u1_n188, u2_u5_u1_n95, u2_u5_u1_n96, u2_u5_u1_n97, u2_u5_u1_n98, u2_u5_u1_n99, u2_u5_u2_n100, 
       u2_u5_u2_n101, u2_u5_u2_n102, u2_u5_u2_n103, u2_u5_u2_n104, u2_u5_u2_n105, u2_u5_u2_n106, u2_u5_u2_n107, u2_u5_u2_n108, u2_u5_u2_n109, 
       u2_u5_u2_n110, u2_u5_u2_n111, u2_u5_u2_n112, u2_u5_u2_n113, u2_u5_u2_n114, u2_u5_u2_n115, u2_u5_u2_n116, u2_u5_u2_n117, u2_u5_u2_n118, 
       u2_u5_u2_n119, u2_u5_u2_n120, u2_u5_u2_n121, u2_u5_u2_n122, u2_u5_u2_n123, u2_u5_u2_n124, u2_u5_u2_n125, u2_u5_u2_n126, u2_u5_u2_n127, 
       u2_u5_u2_n128, u2_u5_u2_n129, u2_u5_u2_n130, u2_u5_u2_n131, u2_u5_u2_n132, u2_u5_u2_n133, u2_u5_u2_n134, u2_u5_u2_n135, u2_u5_u2_n136, 
       u2_u5_u2_n137, u2_u5_u2_n138, u2_u5_u2_n139, u2_u5_u2_n140, u2_u5_u2_n141, u2_u5_u2_n142, u2_u5_u2_n143, u2_u5_u2_n144, u2_u5_u2_n145, 
       u2_u5_u2_n146, u2_u5_u2_n147, u2_u5_u2_n148, u2_u5_u2_n149, u2_u5_u2_n150, u2_u5_u2_n151, u2_u5_u2_n152, u2_u5_u2_n153, u2_u5_u2_n154, 
       u2_u5_u2_n155, u2_u5_u2_n156, u2_u5_u2_n157, u2_u5_u2_n158, u2_u5_u2_n159, u2_u5_u2_n160, u2_u5_u2_n161, u2_u5_u2_n162, u2_u5_u2_n163, 
       u2_u5_u2_n164, u2_u5_u2_n165, u2_u5_u2_n166, u2_u5_u2_n167, u2_u5_u2_n168, u2_u5_u2_n169, u2_u5_u2_n170, u2_u5_u2_n171, u2_u5_u2_n172, 
       u2_u5_u2_n173, u2_u5_u2_n174, u2_u5_u2_n175, u2_u5_u2_n176, u2_u5_u2_n177, u2_u5_u2_n178, u2_u5_u2_n179, u2_u5_u2_n180, u2_u5_u2_n181, 
       u2_u5_u2_n182, u2_u5_u2_n183, u2_u5_u2_n184, u2_u5_u2_n185, u2_u5_u2_n186, u2_u5_u2_n187, u2_u5_u2_n188, u2_u5_u2_n95, u2_u5_u2_n96, 
       u2_u5_u2_n97, u2_u5_u2_n98, u2_u5_u2_n99, u2_u5_u3_n100, u2_u5_u3_n101, u2_u5_u3_n102, u2_u5_u3_n103, u2_u5_u3_n104, u2_u5_u3_n105, 
       u2_u5_u3_n106, u2_u5_u3_n107, u2_u5_u3_n108, u2_u5_u3_n109, u2_u5_u3_n110, u2_u5_u3_n111, u2_u5_u3_n112, u2_u5_u3_n113, u2_u5_u3_n114, 
       u2_u5_u3_n115, u2_u5_u3_n116, u2_u5_u3_n117, u2_u5_u3_n118, u2_u5_u3_n119, u2_u5_u3_n120, u2_u5_u3_n121, u2_u5_u3_n122, u2_u5_u3_n123, 
       u2_u5_u3_n124, u2_u5_u3_n125, u2_u5_u3_n126, u2_u5_u3_n127, u2_u5_u3_n128, u2_u5_u3_n129, u2_u5_u3_n130, u2_u5_u3_n131, u2_u5_u3_n132, 
       u2_u5_u3_n133, u2_u5_u3_n134, u2_u5_u3_n135, u2_u5_u3_n136, u2_u5_u3_n137, u2_u5_u3_n138, u2_u5_u3_n139, u2_u5_u3_n140, u2_u5_u3_n141, 
       u2_u5_u3_n142, u2_u5_u3_n143, u2_u5_u3_n144, u2_u5_u3_n145, u2_u5_u3_n146, u2_u5_u3_n147, u2_u5_u3_n148, u2_u5_u3_n149, u2_u5_u3_n150, 
       u2_u5_u3_n151, u2_u5_u3_n152, u2_u5_u3_n153, u2_u5_u3_n154, u2_u5_u3_n155, u2_u5_u3_n156, u2_u5_u3_n157, u2_u5_u3_n158, u2_u5_u3_n159, 
       u2_u5_u3_n160, u2_u5_u3_n161, u2_u5_u3_n162, u2_u5_u3_n163, u2_u5_u3_n164, u2_u5_u3_n165, u2_u5_u3_n166, u2_u5_u3_n167, u2_u5_u3_n168, 
       u2_u5_u3_n169, u2_u5_u3_n170, u2_u5_u3_n171, u2_u5_u3_n172, u2_u5_u3_n173, u2_u5_u3_n174, u2_u5_u3_n175, u2_u5_u3_n176, u2_u5_u3_n177, 
       u2_u5_u3_n178, u2_u5_u3_n179, u2_u5_u3_n180, u2_u5_u3_n181, u2_u5_u3_n182, u2_u5_u3_n183, u2_u5_u3_n184, u2_u5_u3_n185, u2_u5_u3_n186, 
       u2_u5_u3_n94, u2_u5_u3_n95, u2_u5_u3_n96, u2_u5_u3_n97, u2_u5_u3_n98, u2_u5_u3_n99, u2_u5_u4_n100, u2_u5_u4_n101, u2_u5_u4_n102, 
       u2_u5_u4_n103, u2_u5_u4_n104, u2_u5_u4_n105, u2_u5_u4_n106, u2_u5_u4_n107, u2_u5_u4_n108, u2_u5_u4_n109, u2_u5_u4_n110, u2_u5_u4_n111, 
       u2_u5_u4_n112, u2_u5_u4_n113, u2_u5_u4_n114, u2_u5_u4_n115, u2_u5_u4_n116, u2_u5_u4_n117, u2_u5_u4_n118, u2_u5_u4_n119, u2_u5_u4_n120, 
       u2_u5_u4_n121, u2_u5_u4_n122, u2_u5_u4_n123, u2_u5_u4_n124, u2_u5_u4_n125, u2_u5_u4_n126, u2_u5_u4_n127, u2_u5_u4_n128, u2_u5_u4_n129, 
       u2_u5_u4_n130, u2_u5_u4_n131, u2_u5_u4_n132, u2_u5_u4_n133, u2_u5_u4_n134, u2_u5_u4_n135, u2_u5_u4_n136, u2_u5_u4_n137, u2_u5_u4_n138, 
       u2_u5_u4_n139, u2_u5_u4_n140, u2_u5_u4_n141, u2_u5_u4_n142, u2_u5_u4_n143, u2_u5_u4_n144, u2_u5_u4_n145, u2_u5_u4_n146, u2_u5_u4_n147, 
       u2_u5_u4_n148, u2_u5_u4_n149, u2_u5_u4_n150, u2_u5_u4_n151, u2_u5_u4_n152, u2_u5_u4_n153, u2_u5_u4_n154, u2_u5_u4_n155, u2_u5_u4_n156, 
       u2_u5_u4_n157, u2_u5_u4_n158, u2_u5_u4_n159, u2_u5_u4_n160, u2_u5_u4_n161, u2_u5_u4_n162, u2_u5_u4_n163, u2_u5_u4_n164, u2_u5_u4_n165, 
       u2_u5_u4_n166, u2_u5_u4_n167, u2_u5_u4_n168, u2_u5_u4_n169, u2_u5_u4_n170, u2_u5_u4_n171, u2_u5_u4_n172, u2_u5_u4_n173, u2_u5_u4_n174, 
       u2_u5_u4_n175, u2_u5_u4_n176, u2_u5_u4_n177, u2_u5_u4_n178, u2_u5_u4_n179, u2_u5_u4_n180, u2_u5_u4_n181, u2_u5_u4_n182, u2_u5_u4_n183, 
       u2_u5_u4_n184, u2_u5_u4_n185, u2_u5_u4_n186, u2_u5_u4_n94, u2_u5_u4_n95, u2_u5_u4_n96, u2_u5_u4_n97, u2_u5_u4_n98, u2_u5_u4_n99, 
       u2_u5_u5_n100, u2_u5_u5_n101, u2_u5_u5_n102, u2_u5_u5_n103, u2_u5_u5_n104, u2_u5_u5_n105, u2_u5_u5_n106, u2_u5_u5_n107, u2_u5_u5_n108, 
       u2_u5_u5_n109, u2_u5_u5_n110, u2_u5_u5_n111, u2_u5_u5_n112, u2_u5_u5_n113, u2_u5_u5_n114, u2_u5_u5_n115, u2_u5_u5_n116, u2_u5_u5_n117, 
       u2_u5_u5_n118, u2_u5_u5_n119, u2_u5_u5_n120, u2_u5_u5_n121, u2_u5_u5_n122, u2_u5_u5_n123, u2_u5_u5_n124, u2_u5_u5_n125, u2_u5_u5_n126, 
       u2_u5_u5_n127, u2_u5_u5_n128, u2_u5_u5_n129, u2_u5_u5_n130, u2_u5_u5_n131, u2_u5_u5_n132, u2_u5_u5_n133, u2_u5_u5_n134, u2_u5_u5_n135, 
       u2_u5_u5_n136, u2_u5_u5_n137, u2_u5_u5_n138, u2_u5_u5_n139, u2_u5_u5_n140, u2_u5_u5_n141, u2_u5_u5_n142, u2_u5_u5_n143, u2_u5_u5_n144, 
       u2_u5_u5_n145, u2_u5_u5_n146, u2_u5_u5_n147, u2_u5_u5_n148, u2_u5_u5_n149, u2_u5_u5_n150, u2_u5_u5_n151, u2_u5_u5_n152, u2_u5_u5_n153, 
       u2_u5_u5_n154, u2_u5_u5_n155, u2_u5_u5_n156, u2_u5_u5_n157, u2_u5_u5_n158, u2_u5_u5_n159, u2_u5_u5_n160, u2_u5_u5_n161, u2_u5_u5_n162, 
       u2_u5_u5_n163, u2_u5_u5_n164, u2_u5_u5_n165, u2_u5_u5_n166, u2_u5_u5_n167, u2_u5_u5_n168, u2_u5_u5_n169, u2_u5_u5_n170, u2_u5_u5_n171, 
       u2_u5_u5_n172, u2_u5_u5_n173, u2_u5_u5_n174, u2_u5_u5_n175, u2_u5_u5_n176, u2_u5_u5_n177, u2_u5_u5_n178, u2_u5_u5_n179, u2_u5_u5_n180, 
       u2_u5_u5_n181, u2_u5_u5_n182, u2_u5_u5_n183, u2_u5_u5_n184, u2_u5_u5_n185, u2_u5_u5_n186, u2_u5_u5_n187, u2_u5_u5_n188, u2_u5_u5_n189, 
       u2_u5_u5_n190, u2_u5_u5_n191, u2_u5_u5_n192, u2_u5_u5_n193, u2_u5_u5_n194, u2_u5_u5_n195, u2_u5_u5_n196, u2_u5_u5_n99, u2_u5_u6_n100, 
       u2_u5_u6_n101, u2_u5_u6_n102, u2_u5_u6_n103, u2_u5_u6_n104, u2_u5_u6_n105, u2_u5_u6_n106, u2_u5_u6_n107, u2_u5_u6_n108, u2_u5_u6_n109, 
       u2_u5_u6_n110, u2_u5_u6_n111, u2_u5_u6_n112, u2_u5_u6_n113, u2_u5_u6_n114, u2_u5_u6_n115, u2_u5_u6_n116, u2_u5_u6_n117, u2_u5_u6_n118, 
       u2_u5_u6_n119, u2_u5_u6_n120, u2_u5_u6_n121, u2_u5_u6_n122, u2_u5_u6_n123, u2_u5_u6_n124, u2_u5_u6_n125, u2_u5_u6_n126, u2_u5_u6_n127, 
       u2_u5_u6_n128, u2_u5_u6_n129, u2_u5_u6_n130, u2_u5_u6_n131, u2_u5_u6_n132, u2_u5_u6_n133, u2_u5_u6_n134, u2_u5_u6_n135, u2_u5_u6_n136, 
       u2_u5_u6_n137, u2_u5_u6_n138, u2_u5_u6_n139, u2_u5_u6_n140, u2_u5_u6_n141, u2_u5_u6_n142, u2_u5_u6_n143, u2_u5_u6_n144, u2_u5_u6_n145, 
       u2_u5_u6_n146, u2_u5_u6_n147, u2_u5_u6_n148, u2_u5_u6_n149, u2_u5_u6_n150, u2_u5_u6_n151, u2_u5_u6_n152, u2_u5_u6_n153, u2_u5_u6_n154, 
       u2_u5_u6_n155, u2_u5_u6_n156, u2_u5_u6_n157, u2_u5_u6_n158, u2_u5_u6_n159, u2_u5_u6_n160, u2_u5_u6_n161, u2_u5_u6_n162, u2_u5_u6_n163, 
       u2_u5_u6_n164, u2_u5_u6_n165, u2_u5_u6_n166, u2_u5_u6_n167, u2_u5_u6_n168, u2_u5_u6_n169, u2_u5_u6_n170, u2_u5_u6_n171, u2_u5_u6_n172, 
       u2_u5_u6_n173, u2_u5_u6_n174, u2_u5_u6_n88, u2_u5_u6_n89, u2_u5_u6_n90, u2_u5_u6_n91, u2_u5_u6_n92, u2_u5_u6_n93, u2_u5_u6_n94, 
       u2_u5_u6_n95, u2_u5_u6_n96, u2_u5_u6_n97, u2_u5_u6_n98, u2_u5_u6_n99, u2_u5_u7_n100, u2_u5_u7_n101, u2_u5_u7_n102, u2_u5_u7_n103, 
       u2_u5_u7_n104, u2_u5_u7_n105, u2_u5_u7_n106, u2_u5_u7_n107, u2_u5_u7_n108, u2_u5_u7_n109, u2_u5_u7_n110, u2_u5_u7_n111, u2_u5_u7_n112, 
       u2_u5_u7_n113, u2_u5_u7_n114, u2_u5_u7_n115, u2_u5_u7_n116, u2_u5_u7_n117, u2_u5_u7_n118, u2_u5_u7_n119, u2_u5_u7_n120, u2_u5_u7_n121, 
       u2_u5_u7_n122, u2_u5_u7_n123, u2_u5_u7_n124, u2_u5_u7_n125, u2_u5_u7_n126, u2_u5_u7_n127, u2_u5_u7_n128, u2_u5_u7_n129, u2_u5_u7_n130, 
       u2_u5_u7_n131, u2_u5_u7_n132, u2_u5_u7_n133, u2_u5_u7_n134, u2_u5_u7_n135, u2_u5_u7_n136, u2_u5_u7_n137, u2_u5_u7_n138, u2_u5_u7_n139, 
       u2_u5_u7_n140, u2_u5_u7_n141, u2_u5_u7_n142, u2_u5_u7_n143, u2_u5_u7_n144, u2_u5_u7_n145, u2_u5_u7_n146, u2_u5_u7_n147, u2_u5_u7_n148, 
       u2_u5_u7_n149, u2_u5_u7_n150, u2_u5_u7_n151, u2_u5_u7_n152, u2_u5_u7_n153, u2_u5_u7_n154, u2_u5_u7_n155, u2_u5_u7_n156, u2_u5_u7_n157, 
       u2_u5_u7_n158, u2_u5_u7_n159, u2_u5_u7_n160, u2_u5_u7_n161, u2_u5_u7_n162, u2_u5_u7_n163, u2_u5_u7_n164, u2_u5_u7_n165, u2_u5_u7_n166, 
       u2_u5_u7_n167, u2_u5_u7_n168, u2_u5_u7_n169, u2_u5_u7_n170, u2_u5_u7_n171, u2_u5_u7_n172, u2_u5_u7_n173, u2_u5_u7_n174, u2_u5_u7_n175, 
       u2_u5_u7_n176, u2_u5_u7_n177, u2_u5_u7_n178, u2_u5_u7_n179, u2_u5_u7_n180, u2_u5_u7_n91, u2_u5_u7_n92, u2_u5_u7_n93, u2_u5_u7_n94, 
       u2_u5_u7_n95, u2_u5_u7_n96, u2_u5_u7_n97, u2_u5_u7_n98, u2_u5_u7_n99, u2_u6_X_1, u2_u6_X_11, u2_u6_X_12, u2_u6_X_13, 
       u2_u6_X_14, u2_u6_X_15, u2_u6_X_16, u2_u6_X_17, u2_u6_X_18, u2_u6_X_19, u2_u6_X_2, u2_u6_X_20, u2_u6_X_21, 
       u2_u6_X_23, u2_u6_X_24, u2_u6_X_25, u2_u6_X_26, u2_u6_X_29, u2_u6_X_30, u2_u6_X_31, u2_u6_X_32, u2_u6_X_34, 
       u2_u6_X_35, u2_u6_X_36, u2_u6_X_37, u2_u6_X_38, u2_u6_X_39, u2_u6_X_41, u2_u6_X_42, u2_u6_X_43, u2_u6_X_44, 
       u2_u6_X_47, u2_u6_X_48, u2_u6_X_5, u2_u6_X_6, u2_u6_X_7, u2_u6_X_8, u2_u6_u0_n100, u2_u6_u0_n101, u2_u6_u0_n102, 
       u2_u6_u0_n103, u2_u6_u0_n104, u2_u6_u0_n105, u2_u6_u0_n106, u2_u6_u0_n107, u2_u6_u0_n108, u2_u6_u0_n109, u2_u6_u0_n110, u2_u6_u0_n111, 
       u2_u6_u0_n112, u2_u6_u0_n113, u2_u6_u0_n114, u2_u6_u0_n115, u2_u6_u0_n116, u2_u6_u0_n117, u2_u6_u0_n118, u2_u6_u0_n119, u2_u6_u0_n120, 
       u2_u6_u0_n121, u2_u6_u0_n122, u2_u6_u0_n123, u2_u6_u0_n124, u2_u6_u0_n125, u2_u6_u0_n126, u2_u6_u0_n127, u2_u6_u0_n128, u2_u6_u0_n129, 
       u2_u6_u0_n130, u2_u6_u0_n131, u2_u6_u0_n132, u2_u6_u0_n133, u2_u6_u0_n134, u2_u6_u0_n135, u2_u6_u0_n136, u2_u6_u0_n137, u2_u6_u0_n138, 
       u2_u6_u0_n139, u2_u6_u0_n140, u2_u6_u0_n141, u2_u6_u0_n142, u2_u6_u0_n143, u2_u6_u0_n144, u2_u6_u0_n145, u2_u6_u0_n146, u2_u6_u0_n147, 
       u2_u6_u0_n148, u2_u6_u0_n149, u2_u6_u0_n150, u2_u6_u0_n151, u2_u6_u0_n152, u2_u6_u0_n153, u2_u6_u0_n154, u2_u6_u0_n155, u2_u6_u0_n156, 
       u2_u6_u0_n157, u2_u6_u0_n158, u2_u6_u0_n159, u2_u6_u0_n160, u2_u6_u0_n161, u2_u6_u0_n162, u2_u6_u0_n163, u2_u6_u0_n164, u2_u6_u0_n165, 
       u2_u6_u0_n166, u2_u6_u0_n167, u2_u6_u0_n168, u2_u6_u0_n169, u2_u6_u0_n170, u2_u6_u0_n171, u2_u6_u0_n172, u2_u6_u0_n173, u2_u6_u0_n174, 
       u2_u6_u0_n88, u2_u6_u0_n89, u2_u6_u0_n90, u2_u6_u0_n91, u2_u6_u0_n92, u2_u6_u0_n93, u2_u6_u0_n94, u2_u6_u0_n95, u2_u6_u0_n96, 
       u2_u6_u0_n97, u2_u6_u0_n98, u2_u6_u0_n99, u2_u6_u1_n100, u2_u6_u1_n101, u2_u6_u1_n102, u2_u6_u1_n103, u2_u6_u1_n104, u2_u6_u1_n105, 
       u2_u6_u1_n106, u2_u6_u1_n107, u2_u6_u1_n108, u2_u6_u1_n109, u2_u6_u1_n110, u2_u6_u1_n111, u2_u6_u1_n112, u2_u6_u1_n113, u2_u6_u1_n114, 
       u2_u6_u1_n115, u2_u6_u1_n116, u2_u6_u1_n117, u2_u6_u1_n118, u2_u6_u1_n119, u2_u6_u1_n120, u2_u6_u1_n121, u2_u6_u1_n122, u2_u6_u1_n123, 
       u2_u6_u1_n124, u2_u6_u1_n125, u2_u6_u1_n126, u2_u6_u1_n127, u2_u6_u1_n128, u2_u6_u1_n129, u2_u6_u1_n130, u2_u6_u1_n131, u2_u6_u1_n132, 
       u2_u6_u1_n133, u2_u6_u1_n134, u2_u6_u1_n135, u2_u6_u1_n136, u2_u6_u1_n137, u2_u6_u1_n138, u2_u6_u1_n139, u2_u6_u1_n140, u2_u6_u1_n141, 
       u2_u6_u1_n142, u2_u6_u1_n143, u2_u6_u1_n144, u2_u6_u1_n145, u2_u6_u1_n146, u2_u6_u1_n147, u2_u6_u1_n148, u2_u6_u1_n149, u2_u6_u1_n150, 
       u2_u6_u1_n151, u2_u6_u1_n152, u2_u6_u1_n153, u2_u6_u1_n154, u2_u6_u1_n155, u2_u6_u1_n156, u2_u6_u1_n157, u2_u6_u1_n158, u2_u6_u1_n159, 
       u2_u6_u1_n160, u2_u6_u1_n161, u2_u6_u1_n162, u2_u6_u1_n163, u2_u6_u1_n164, u2_u6_u1_n165, u2_u6_u1_n166, u2_u6_u1_n167, u2_u6_u1_n168, 
       u2_u6_u1_n169, u2_u6_u1_n170, u2_u6_u1_n171, u2_u6_u1_n172, u2_u6_u1_n173, u2_u6_u1_n174, u2_u6_u1_n175, u2_u6_u1_n176, u2_u6_u1_n177, 
       u2_u6_u1_n178, u2_u6_u1_n179, u2_u6_u1_n180, u2_u6_u1_n181, u2_u6_u1_n182, u2_u6_u1_n183, u2_u6_u1_n184, u2_u6_u1_n185, u2_u6_u1_n186, 
       u2_u6_u1_n187, u2_u6_u1_n188, u2_u6_u1_n95, u2_u6_u1_n96, u2_u6_u1_n97, u2_u6_u1_n98, u2_u6_u1_n99, u2_u6_u2_n100, u2_u6_u2_n101, 
       u2_u6_u2_n102, u2_u6_u2_n103, u2_u6_u2_n104, u2_u6_u2_n105, u2_u6_u2_n106, u2_u6_u2_n107, u2_u6_u2_n108, u2_u6_u2_n109, u2_u6_u2_n110, 
       u2_u6_u2_n111, u2_u6_u2_n112, u2_u6_u2_n113, u2_u6_u2_n114, u2_u6_u2_n115, u2_u6_u2_n116, u2_u6_u2_n117, u2_u6_u2_n118, u2_u6_u2_n119, 
       u2_u6_u2_n120, u2_u6_u2_n121, u2_u6_u2_n122, u2_u6_u2_n123, u2_u6_u2_n124, u2_u6_u2_n125, u2_u6_u2_n126, u2_u6_u2_n127, u2_u6_u2_n128, 
       u2_u6_u2_n129, u2_u6_u2_n130, u2_u6_u2_n131, u2_u6_u2_n132, u2_u6_u2_n133, u2_u6_u2_n134, u2_u6_u2_n135, u2_u6_u2_n136, u2_u6_u2_n137, 
       u2_u6_u2_n138, u2_u6_u2_n139, u2_u6_u2_n140, u2_u6_u2_n141, u2_u6_u2_n142, u2_u6_u2_n143, u2_u6_u2_n144, u2_u6_u2_n145, u2_u6_u2_n146, 
       u2_u6_u2_n147, u2_u6_u2_n148, u2_u6_u2_n149, u2_u6_u2_n150, u2_u6_u2_n151, u2_u6_u2_n152, u2_u6_u2_n153, u2_u6_u2_n154, u2_u6_u2_n155, 
       u2_u6_u2_n156, u2_u6_u2_n157, u2_u6_u2_n158, u2_u6_u2_n159, u2_u6_u2_n160, u2_u6_u2_n161, u2_u6_u2_n162, u2_u6_u2_n163, u2_u6_u2_n164, 
       u2_u6_u2_n165, u2_u6_u2_n166, u2_u6_u2_n167, u2_u6_u2_n168, u2_u6_u2_n169, u2_u6_u2_n170, u2_u6_u2_n171, u2_u6_u2_n172, u2_u6_u2_n173, 
       u2_u6_u2_n174, u2_u6_u2_n175, u2_u6_u2_n176, u2_u6_u2_n177, u2_u6_u2_n178, u2_u6_u2_n179, u2_u6_u2_n180, u2_u6_u2_n181, u2_u6_u2_n182, 
       u2_u6_u2_n183, u2_u6_u2_n184, u2_u6_u2_n185, u2_u6_u2_n186, u2_u6_u2_n187, u2_u6_u2_n188, u2_u6_u2_n95, u2_u6_u2_n96, u2_u6_u2_n97, 
       u2_u6_u2_n98, u2_u6_u2_n99, u2_u6_u3_n100, u2_u6_u3_n101, u2_u6_u3_n102, u2_u6_u3_n103, u2_u6_u3_n104, u2_u6_u3_n105, u2_u6_u3_n106, 
       u2_u6_u3_n107, u2_u6_u3_n108, u2_u6_u3_n109, u2_u6_u3_n110, u2_u6_u3_n111, u2_u6_u3_n112, u2_u6_u3_n113, u2_u6_u3_n114, u2_u6_u3_n115, 
       u2_u6_u3_n116, u2_u6_u3_n117, u2_u6_u3_n118, u2_u6_u3_n119, u2_u6_u3_n120, u2_u6_u3_n121, u2_u6_u3_n122, u2_u6_u3_n123, u2_u6_u3_n124, 
       u2_u6_u3_n125, u2_u6_u3_n126, u2_u6_u3_n127, u2_u6_u3_n128, u2_u6_u3_n129, u2_u6_u3_n130, u2_u6_u3_n131, u2_u6_u3_n132, u2_u6_u3_n133, 
       u2_u6_u3_n134, u2_u6_u3_n135, u2_u6_u3_n136, u2_u6_u3_n137, u2_u6_u3_n138, u2_u6_u3_n139, u2_u6_u3_n140, u2_u6_u3_n141, u2_u6_u3_n142, 
       u2_u6_u3_n143, u2_u6_u3_n144, u2_u6_u3_n145, u2_u6_u3_n146, u2_u6_u3_n147, u2_u6_u3_n148, u2_u6_u3_n149, u2_u6_u3_n150, u2_u6_u3_n151, 
       u2_u6_u3_n152, u2_u6_u3_n153, u2_u6_u3_n154, u2_u6_u3_n155, u2_u6_u3_n156, u2_u6_u3_n157, u2_u6_u3_n158, u2_u6_u3_n159, u2_u6_u3_n160, 
       u2_u6_u3_n161, u2_u6_u3_n162, u2_u6_u3_n163, u2_u6_u3_n164, u2_u6_u3_n165, u2_u6_u3_n166, u2_u6_u3_n167, u2_u6_u3_n168, u2_u6_u3_n169, 
       u2_u6_u3_n170, u2_u6_u3_n171, u2_u6_u3_n172, u2_u6_u3_n173, u2_u6_u3_n174, u2_u6_u3_n175, u2_u6_u3_n176, u2_u6_u3_n177, u2_u6_u3_n178, 
       u2_u6_u3_n179, u2_u6_u3_n180, u2_u6_u3_n181, u2_u6_u3_n182, u2_u6_u3_n183, u2_u6_u3_n184, u2_u6_u3_n185, u2_u6_u3_n186, u2_u6_u3_n94, 
       u2_u6_u3_n95, u2_u6_u3_n96, u2_u6_u3_n97, u2_u6_u3_n98, u2_u6_u3_n99, u2_u6_u4_n100, u2_u6_u4_n101, u2_u6_u4_n102, u2_u6_u4_n103, 
       u2_u6_u4_n104, u2_u6_u4_n105, u2_u6_u4_n106, u2_u6_u4_n107, u2_u6_u4_n108, u2_u6_u4_n109, u2_u6_u4_n110, u2_u6_u4_n111, u2_u6_u4_n112, 
       u2_u6_u4_n113, u2_u6_u4_n114, u2_u6_u4_n115, u2_u6_u4_n116, u2_u6_u4_n117, u2_u6_u4_n118, u2_u6_u4_n119, u2_u6_u4_n120, u2_u6_u4_n121, 
       u2_u6_u4_n122, u2_u6_u4_n123, u2_u6_u4_n124, u2_u6_u4_n125, u2_u6_u4_n126, u2_u6_u4_n127, u2_u6_u4_n128, u2_u6_u4_n129, u2_u6_u4_n130, 
       u2_u6_u4_n131, u2_u6_u4_n132, u2_u6_u4_n133, u2_u6_u4_n134, u2_u6_u4_n135, u2_u6_u4_n136, u2_u6_u4_n137, u2_u6_u4_n138, u2_u6_u4_n139, 
       u2_u6_u4_n140, u2_u6_u4_n141, u2_u6_u4_n142, u2_u6_u4_n143, u2_u6_u4_n144, u2_u6_u4_n145, u2_u6_u4_n146, u2_u6_u4_n147, u2_u6_u4_n148, 
       u2_u6_u4_n149, u2_u6_u4_n150, u2_u6_u4_n151, u2_u6_u4_n152, u2_u6_u4_n153, u2_u6_u4_n154, u2_u6_u4_n155, u2_u6_u4_n156, u2_u6_u4_n157, 
       u2_u6_u4_n158, u2_u6_u4_n159, u2_u6_u4_n160, u2_u6_u4_n161, u2_u6_u4_n162, u2_u6_u4_n163, u2_u6_u4_n164, u2_u6_u4_n165, u2_u6_u4_n166, 
       u2_u6_u4_n167, u2_u6_u4_n168, u2_u6_u4_n169, u2_u6_u4_n170, u2_u6_u4_n171, u2_u6_u4_n172, u2_u6_u4_n173, u2_u6_u4_n174, u2_u6_u4_n175, 
       u2_u6_u4_n176, u2_u6_u4_n177, u2_u6_u4_n178, u2_u6_u4_n179, u2_u6_u4_n180, u2_u6_u4_n181, u2_u6_u4_n182, u2_u6_u4_n183, u2_u6_u4_n184, 
       u2_u6_u4_n185, u2_u6_u4_n186, u2_u6_u4_n94, u2_u6_u4_n95, u2_u6_u4_n96, u2_u6_u4_n97, u2_u6_u4_n98, u2_u6_u4_n99, u2_u6_u5_n100, 
       u2_u6_u5_n101, u2_u6_u5_n102, u2_u6_u5_n103, u2_u6_u5_n104, u2_u6_u5_n105, u2_u6_u5_n106, u2_u6_u5_n107, u2_u6_u5_n108, u2_u6_u5_n109, 
       u2_u6_u5_n110, u2_u6_u5_n111, u2_u6_u5_n112, u2_u6_u5_n113, u2_u6_u5_n114, u2_u6_u5_n115, u2_u6_u5_n116, u2_u6_u5_n117, u2_u6_u5_n118, 
       u2_u6_u5_n119, u2_u6_u5_n120, u2_u6_u5_n121, u2_u6_u5_n122, u2_u6_u5_n123, u2_u6_u5_n124, u2_u6_u5_n125, u2_u6_u5_n126, u2_u6_u5_n127, 
       u2_u6_u5_n128, u2_u6_u5_n129, u2_u6_u5_n130, u2_u6_u5_n131, u2_u6_u5_n132, u2_u6_u5_n133, u2_u6_u5_n134, u2_u6_u5_n135, u2_u6_u5_n136, 
       u2_u6_u5_n137, u2_u6_u5_n138, u2_u6_u5_n139, u2_u6_u5_n140, u2_u6_u5_n141, u2_u6_u5_n142, u2_u6_u5_n143, u2_u6_u5_n144, u2_u6_u5_n145, 
       u2_u6_u5_n146, u2_u6_u5_n147, u2_u6_u5_n148, u2_u6_u5_n149, u2_u6_u5_n150, u2_u6_u5_n151, u2_u6_u5_n152, u2_u6_u5_n153, u2_u6_u5_n154, 
       u2_u6_u5_n155, u2_u6_u5_n156, u2_u6_u5_n157, u2_u6_u5_n158, u2_u6_u5_n159, u2_u6_u5_n160, u2_u6_u5_n161, u2_u6_u5_n162, u2_u6_u5_n163, 
       u2_u6_u5_n164, u2_u6_u5_n165, u2_u6_u5_n166, u2_u6_u5_n167, u2_u6_u5_n168, u2_u6_u5_n169, u2_u6_u5_n170, u2_u6_u5_n171, u2_u6_u5_n172, 
       u2_u6_u5_n173, u2_u6_u5_n174, u2_u6_u5_n175, u2_u6_u5_n176, u2_u6_u5_n177, u2_u6_u5_n178, u2_u6_u5_n179, u2_u6_u5_n180, u2_u6_u5_n181, 
       u2_u6_u5_n182, u2_u6_u5_n183, u2_u6_u5_n184, u2_u6_u5_n185, u2_u6_u5_n186, u2_u6_u5_n187, u2_u6_u5_n188, u2_u6_u5_n189, u2_u6_u5_n190, 
       u2_u6_u5_n191, u2_u6_u5_n192, u2_u6_u5_n193, u2_u6_u5_n194, u2_u6_u5_n195, u2_u6_u5_n196, u2_u6_u5_n99, u2_u6_u6_n100, u2_u6_u6_n101, 
       u2_u6_u6_n102, u2_u6_u6_n103, u2_u6_u6_n104, u2_u6_u6_n105, u2_u6_u6_n106, u2_u6_u6_n107, u2_u6_u6_n108, u2_u6_u6_n109, u2_u6_u6_n110, 
       u2_u6_u6_n111, u2_u6_u6_n112, u2_u6_u6_n113, u2_u6_u6_n114, u2_u6_u6_n115, u2_u6_u6_n116, u2_u6_u6_n117, u2_u6_u6_n118, u2_u6_u6_n119, 
       u2_u6_u6_n120, u2_u6_u6_n121, u2_u6_u6_n122, u2_u6_u6_n123, u2_u6_u6_n124, u2_u6_u6_n125, u2_u6_u6_n126, u2_u6_u6_n127, u2_u6_u6_n128, 
       u2_u6_u6_n129, u2_u6_u6_n130, u2_u6_u6_n131, u2_u6_u6_n132, u2_u6_u6_n133, u2_u6_u6_n134, u2_u6_u6_n135, u2_u6_u6_n136, u2_u6_u6_n137, 
       u2_u6_u6_n138, u2_u6_u6_n139, u2_u6_u6_n140, u2_u6_u6_n141, u2_u6_u6_n142, u2_u6_u6_n143, u2_u6_u6_n144, u2_u6_u6_n145, u2_u6_u6_n146, 
       u2_u6_u6_n147, u2_u6_u6_n148, u2_u6_u6_n149, u2_u6_u6_n150, u2_u6_u6_n151, u2_u6_u6_n152, u2_u6_u6_n153, u2_u6_u6_n154, u2_u6_u6_n155, 
       u2_u6_u6_n156, u2_u6_u6_n157, u2_u6_u6_n158, u2_u6_u6_n159, u2_u6_u6_n160, u2_u6_u6_n161, u2_u6_u6_n162, u2_u6_u6_n163, u2_u6_u6_n164, 
       u2_u6_u6_n165, u2_u6_u6_n166, u2_u6_u6_n167, u2_u6_u6_n168, u2_u6_u6_n169, u2_u6_u6_n170, u2_u6_u6_n171, u2_u6_u6_n172, u2_u6_u6_n173, 
       u2_u6_u6_n174, u2_u6_u6_n88, u2_u6_u6_n89, u2_u6_u6_n90, u2_u6_u6_n91, u2_u6_u6_n92, u2_u6_u6_n93, u2_u6_u6_n94, u2_u6_u6_n95, 
       u2_u6_u6_n96, u2_u6_u6_n97, u2_u6_u6_n98, u2_u6_u6_n99, u2_u6_u7_n100, u2_u6_u7_n101, u2_u6_u7_n102, u2_u6_u7_n103, u2_u6_u7_n104, 
       u2_u6_u7_n105, u2_u6_u7_n106, u2_u6_u7_n107, u2_u6_u7_n108, u2_u6_u7_n109, u2_u6_u7_n110, u2_u6_u7_n111, u2_u6_u7_n112, u2_u6_u7_n113, 
       u2_u6_u7_n114, u2_u6_u7_n115, u2_u6_u7_n116, u2_u6_u7_n117, u2_u6_u7_n118, u2_u6_u7_n119, u2_u6_u7_n120, u2_u6_u7_n121, u2_u6_u7_n122, 
       u2_u6_u7_n123, u2_u6_u7_n124, u2_u6_u7_n125, u2_u6_u7_n126, u2_u6_u7_n127, u2_u6_u7_n128, u2_u6_u7_n129, u2_u6_u7_n130, u2_u6_u7_n131, 
       u2_u6_u7_n132, u2_u6_u7_n133, u2_u6_u7_n134, u2_u6_u7_n135, u2_u6_u7_n136, u2_u6_u7_n137, u2_u6_u7_n138, u2_u6_u7_n139, u2_u6_u7_n140, 
       u2_u6_u7_n141, u2_u6_u7_n142, u2_u6_u7_n143, u2_u6_u7_n144, u2_u6_u7_n145, u2_u6_u7_n146, u2_u6_u7_n147, u2_u6_u7_n148, u2_u6_u7_n149, 
       u2_u6_u7_n150, u2_u6_u7_n151, u2_u6_u7_n152, u2_u6_u7_n153, u2_u6_u7_n154, u2_u6_u7_n155, u2_u6_u7_n156, u2_u6_u7_n157, u2_u6_u7_n158, 
       u2_u6_u7_n159, u2_u6_u7_n160, u2_u6_u7_n161, u2_u6_u7_n162, u2_u6_u7_n163, u2_u6_u7_n164, u2_u6_u7_n165, u2_u6_u7_n166, u2_u6_u7_n167, 
       u2_u6_u7_n168, u2_u6_u7_n169, u2_u6_u7_n170, u2_u6_u7_n171, u2_u6_u7_n172, u2_u6_u7_n173, u2_u6_u7_n174, u2_u6_u7_n175, u2_u6_u7_n176, 
       u2_u6_u7_n177, u2_u6_u7_n178, u2_u6_u7_n179, u2_u6_u7_n180, u2_u6_u7_n91, u2_u6_u7_n92, u2_u6_u7_n93, u2_u6_u7_n94, u2_u6_u7_n95, 
       u2_u6_u7_n96, u2_u6_u7_n97, u2_u6_u7_n98, u2_u6_u7_n99, u2_u8_X_10, u2_u8_X_11, u2_u8_X_12, u2_u8_X_13, u2_u8_X_14, 
       u2_u8_X_16, u2_u8_X_17, u2_u8_X_18, u2_u8_X_19, u2_u8_X_2, u2_u8_X_20, u2_u8_X_21, u2_u8_X_22, u2_u8_X_23, 
       u2_u8_X_24, u2_u8_X_25, u2_u8_X_26, u2_u8_X_4, u2_u8_X_5, u2_u8_X_6, u2_u8_X_7, u2_u8_X_8, u2_u8_X_9, 
       u2_u8_u0_n100, u2_u8_u0_n101, u2_u8_u0_n102, u2_u8_u0_n103, u2_u8_u0_n104, u2_u8_u0_n105, u2_u8_u0_n106, u2_u8_u0_n107, u2_u8_u0_n108, 
       u2_u8_u0_n109, u2_u8_u0_n110, u2_u8_u0_n111, u2_u8_u0_n112, u2_u8_u0_n113, u2_u8_u0_n114, u2_u8_u0_n115, u2_u8_u0_n116, u2_u8_u0_n117, 
       u2_u8_u0_n118, u2_u8_u0_n119, u2_u8_u0_n120, u2_u8_u0_n121, u2_u8_u0_n122, u2_u8_u0_n123, u2_u8_u0_n124, u2_u8_u0_n125, u2_u8_u0_n126, 
       u2_u8_u0_n127, u2_u8_u0_n128, u2_u8_u0_n129, u2_u8_u0_n130, u2_u8_u0_n131, u2_u8_u0_n132, u2_u8_u0_n133, u2_u8_u0_n134, u2_u8_u0_n135, 
       u2_u8_u0_n136, u2_u8_u0_n137, u2_u8_u0_n138, u2_u8_u0_n139, u2_u8_u0_n140, u2_u8_u0_n141, u2_u8_u0_n142, u2_u8_u0_n143, u2_u8_u0_n144, 
       u2_u8_u0_n145, u2_u8_u0_n146, u2_u8_u0_n147, u2_u8_u0_n148, u2_u8_u0_n149, u2_u8_u0_n150, u2_u8_u0_n151, u2_u8_u0_n152, u2_u8_u0_n153, 
       u2_u8_u0_n154, u2_u8_u0_n155, u2_u8_u0_n156, u2_u8_u0_n157, u2_u8_u0_n158, u2_u8_u0_n159, u2_u8_u0_n160, u2_u8_u0_n161, u2_u8_u0_n162, 
       u2_u8_u0_n163, u2_u8_u0_n164, u2_u8_u0_n165, u2_u8_u0_n166, u2_u8_u0_n167, u2_u8_u0_n168, u2_u8_u0_n169, u2_u8_u0_n170, u2_u8_u0_n171, 
       u2_u8_u0_n172, u2_u8_u0_n173, u2_u8_u0_n174, u2_u8_u0_n88, u2_u8_u0_n89, u2_u8_u0_n90, u2_u8_u0_n91, u2_u8_u0_n92, u2_u8_u0_n93, 
       u2_u8_u0_n94, u2_u8_u0_n95, u2_u8_u0_n96, u2_u8_u0_n97, u2_u8_u0_n98, u2_u8_u0_n99, u2_u8_u1_n100, u2_u8_u1_n101, u2_u8_u1_n102, 
       u2_u8_u1_n103, u2_u8_u1_n104, u2_u8_u1_n105, u2_u8_u1_n106, u2_u8_u1_n107, u2_u8_u1_n108, u2_u8_u1_n109, u2_u8_u1_n110, u2_u8_u1_n111, 
       u2_u8_u1_n112, u2_u8_u1_n113, u2_u8_u1_n114, u2_u8_u1_n115, u2_u8_u1_n116, u2_u8_u1_n117, u2_u8_u1_n118, u2_u8_u1_n119, u2_u8_u1_n120, 
       u2_u8_u1_n121, u2_u8_u1_n122, u2_u8_u1_n123, u2_u8_u1_n124, u2_u8_u1_n125, u2_u8_u1_n126, u2_u8_u1_n127, u2_u8_u1_n128, u2_u8_u1_n129, 
       u2_u8_u1_n130, u2_u8_u1_n131, u2_u8_u1_n132, u2_u8_u1_n133, u2_u8_u1_n134, u2_u8_u1_n135, u2_u8_u1_n136, u2_u8_u1_n137, u2_u8_u1_n138, 
       u2_u8_u1_n139, u2_u8_u1_n140, u2_u8_u1_n141, u2_u8_u1_n142, u2_u8_u1_n143, u2_u8_u1_n144, u2_u8_u1_n145, u2_u8_u1_n146, u2_u8_u1_n147, 
       u2_u8_u1_n148, u2_u8_u1_n149, u2_u8_u1_n150, u2_u8_u1_n151, u2_u8_u1_n152, u2_u8_u1_n153, u2_u8_u1_n154, u2_u8_u1_n155, u2_u8_u1_n156, 
       u2_u8_u1_n157, u2_u8_u1_n158, u2_u8_u1_n159, u2_u8_u1_n160, u2_u8_u1_n161, u2_u8_u1_n162, u2_u8_u1_n163, u2_u8_u1_n164, u2_u8_u1_n165, 
       u2_u8_u1_n166, u2_u8_u1_n167, u2_u8_u1_n168, u2_u8_u1_n169, u2_u8_u1_n170, u2_u8_u1_n171, u2_u8_u1_n172, u2_u8_u1_n173, u2_u8_u1_n174, 
       u2_u8_u1_n175, u2_u8_u1_n176, u2_u8_u1_n177, u2_u8_u1_n178, u2_u8_u1_n179, u2_u8_u1_n180, u2_u8_u1_n181, u2_u8_u1_n182, u2_u8_u1_n183, 
       u2_u8_u1_n184, u2_u8_u1_n185, u2_u8_u1_n186, u2_u8_u1_n187, u2_u8_u1_n188, u2_u8_u1_n95, u2_u8_u1_n96, u2_u8_u1_n97, u2_u8_u1_n98, 
       u2_u8_u1_n99, u2_u8_u2_n100, u2_u8_u2_n101, u2_u8_u2_n102, u2_u8_u2_n103, u2_u8_u2_n104, u2_u8_u2_n105, u2_u8_u2_n106, u2_u8_u2_n107, 
       u2_u8_u2_n108, u2_u8_u2_n109, u2_u8_u2_n110, u2_u8_u2_n111, u2_u8_u2_n112, u2_u8_u2_n113, u2_u8_u2_n114, u2_u8_u2_n115, u2_u8_u2_n116, 
       u2_u8_u2_n117, u2_u8_u2_n118, u2_u8_u2_n119, u2_u8_u2_n120, u2_u8_u2_n121, u2_u8_u2_n122, u2_u8_u2_n123, u2_u8_u2_n124, u2_u8_u2_n125, 
       u2_u8_u2_n126, u2_u8_u2_n127, u2_u8_u2_n128, u2_u8_u2_n129, u2_u8_u2_n130, u2_u8_u2_n131, u2_u8_u2_n132, u2_u8_u2_n133, u2_u8_u2_n134, 
       u2_u8_u2_n135, u2_u8_u2_n136, u2_u8_u2_n137, u2_u8_u2_n138, u2_u8_u2_n139, u2_u8_u2_n140, u2_u8_u2_n141, u2_u8_u2_n142, u2_u8_u2_n143, 
       u2_u8_u2_n144, u2_u8_u2_n145, u2_u8_u2_n146, u2_u8_u2_n147, u2_u8_u2_n148, u2_u8_u2_n149, u2_u8_u2_n150, u2_u8_u2_n151, u2_u8_u2_n152, 
       u2_u8_u2_n153, u2_u8_u2_n154, u2_u8_u2_n155, u2_u8_u2_n156, u2_u8_u2_n157, u2_u8_u2_n158, u2_u8_u2_n159, u2_u8_u2_n160, u2_u8_u2_n161, 
       u2_u8_u2_n162, u2_u8_u2_n163, u2_u8_u2_n164, u2_u8_u2_n165, u2_u8_u2_n166, u2_u8_u2_n167, u2_u8_u2_n168, u2_u8_u2_n169, u2_u8_u2_n170, 
       u2_u8_u2_n171, u2_u8_u2_n172, u2_u8_u2_n173, u2_u8_u2_n174, u2_u8_u2_n175, u2_u8_u2_n176, u2_u8_u2_n177, u2_u8_u2_n178, u2_u8_u2_n179, 
       u2_u8_u2_n180, u2_u8_u2_n181, u2_u8_u2_n182, u2_u8_u2_n183, u2_u8_u2_n184, u2_u8_u2_n185, u2_u8_u2_n186, u2_u8_u2_n187, u2_u8_u2_n188, 
       u2_u8_u2_n95, u2_u8_u2_n96, u2_u8_u2_n97, u2_u8_u2_n98, u2_u8_u2_n99, u2_u8_u3_n100, u2_u8_u3_n101, u2_u8_u3_n102, u2_u8_u3_n103, 
       u2_u8_u3_n104, u2_u8_u3_n105, u2_u8_u3_n106, u2_u8_u3_n107, u2_u8_u3_n108, u2_u8_u3_n109, u2_u8_u3_n110, u2_u8_u3_n111, u2_u8_u3_n112, 
       u2_u8_u3_n113, u2_u8_u3_n114, u2_u8_u3_n115, u2_u8_u3_n116, u2_u8_u3_n117, u2_u8_u3_n118, u2_u8_u3_n119, u2_u8_u3_n120, u2_u8_u3_n121, 
       u2_u8_u3_n122, u2_u8_u3_n123, u2_u8_u3_n124, u2_u8_u3_n125, u2_u8_u3_n126, u2_u8_u3_n127, u2_u8_u3_n128, u2_u8_u3_n129, u2_u8_u3_n130, 
       u2_u8_u3_n131, u2_u8_u3_n132, u2_u8_u3_n133, u2_u8_u3_n134, u2_u8_u3_n135, u2_u8_u3_n136, u2_u8_u3_n137, u2_u8_u3_n138, u2_u8_u3_n139, 
       u2_u8_u3_n140, u2_u8_u3_n141, u2_u8_u3_n142, u2_u8_u3_n143, u2_u8_u3_n144, u2_u8_u3_n145, u2_u8_u3_n146, u2_u8_u3_n147, u2_u8_u3_n148, 
       u2_u8_u3_n149, u2_u8_u3_n150, u2_u8_u3_n151, u2_u8_u3_n152, u2_u8_u3_n153, u2_u8_u3_n154, u2_u8_u3_n155, u2_u8_u3_n156, u2_u8_u3_n157, 
       u2_u8_u3_n158, u2_u8_u3_n159, u2_u8_u3_n160, u2_u8_u3_n161, u2_u8_u3_n162, u2_u8_u3_n163, u2_u8_u3_n164, u2_u8_u3_n165, u2_u8_u3_n166, 
       u2_u8_u3_n167, u2_u8_u3_n168, u2_u8_u3_n169, u2_u8_u3_n170, u2_u8_u3_n171, u2_u8_u3_n172, u2_u8_u3_n173, u2_u8_u3_n174, u2_u8_u3_n175, 
       u2_u8_u3_n176, u2_u8_u3_n177, u2_u8_u3_n178, u2_u8_u3_n179, u2_u8_u3_n180, u2_u8_u3_n181, u2_u8_u3_n182, u2_u8_u3_n183, u2_u8_u3_n184, 
       u2_u8_u3_n185, u2_u8_u3_n186, u2_u8_u3_n94, u2_u8_u3_n95, u2_u8_u3_n96, u2_u8_u3_n97, u2_u8_u3_n98, u2_u8_u3_n99, u2_u8_u4_n100, 
       u2_u8_u4_n101, u2_u8_u4_n102, u2_u8_u4_n103, u2_u8_u4_n104, u2_u8_u4_n105, u2_u8_u4_n106, u2_u8_u4_n107, u2_u8_u4_n108, u2_u8_u4_n109, 
       u2_u8_u4_n110, u2_u8_u4_n111, u2_u8_u4_n112, u2_u8_u4_n113, u2_u8_u4_n114, u2_u8_u4_n115, u2_u8_u4_n116, u2_u8_u4_n117, u2_u8_u4_n118, 
       u2_u8_u4_n119, u2_u8_u4_n120, u2_u8_u4_n121, u2_u8_u4_n122, u2_u8_u4_n123, u2_u8_u4_n124, u2_u8_u4_n125, u2_u8_u4_n126, u2_u8_u4_n127, 
       u2_u8_u4_n128, u2_u8_u4_n129, u2_u8_u4_n130, u2_u8_u4_n131, u2_u8_u4_n132, u2_u8_u4_n133, u2_u8_u4_n134, u2_u8_u4_n135, u2_u8_u4_n136, 
       u2_u8_u4_n137, u2_u8_u4_n138, u2_u8_u4_n139, u2_u8_u4_n140, u2_u8_u4_n141, u2_u8_u4_n142, u2_u8_u4_n143, u2_u8_u4_n144, u2_u8_u4_n145, 
       u2_u8_u4_n146, u2_u8_u4_n147, u2_u8_u4_n148, u2_u8_u4_n149, u2_u8_u4_n150, u2_u8_u4_n151, u2_u8_u4_n152, u2_u8_u4_n153, u2_u8_u4_n154, 
       u2_u8_u4_n155, u2_u8_u4_n156, u2_u8_u4_n157, u2_u8_u4_n158, u2_u8_u4_n159, u2_u8_u4_n160, u2_u8_u4_n161, u2_u8_u4_n162, u2_u8_u4_n163, 
       u2_u8_u4_n164, u2_u8_u4_n165, u2_u8_u4_n166, u2_u8_u4_n167, u2_u8_u4_n168, u2_u8_u4_n169, u2_u8_u4_n170, u2_u8_u4_n171, u2_u8_u4_n172, 
       u2_u8_u4_n173, u2_u8_u4_n174, u2_u8_u4_n175, u2_u8_u4_n176, u2_u8_u4_n177, u2_u8_u4_n178, u2_u8_u4_n179, u2_u8_u4_n180, u2_u8_u4_n181, 
       u2_u8_u4_n182, u2_u8_u4_n183, u2_u8_u4_n184, u2_u8_u4_n185, u2_u8_u4_n186, u2_u8_u4_n94, u2_u8_u4_n95, u2_u8_u4_n96, u2_u8_u4_n97, 
       u2_u8_u4_n98, u2_u8_u4_n99, u2_u9_X_1, u2_u9_X_2, u2_u9_X_31, u2_u9_X_33, u2_u9_X_35, u2_u9_X_36, u2_u9_X_37, 
       u2_u9_X_38, u2_u9_X_39, u2_u9_X_40, u2_u9_X_41, u2_u9_X_42, u2_u9_X_43, u2_u9_X_44, u2_u9_X_47, u2_u9_X_48, 
       u2_u9_X_5, u2_u9_u0_n100, u2_u9_u0_n101, u2_u9_u0_n102, u2_u9_u0_n103, u2_u9_u0_n104, u2_u9_u0_n105, u2_u9_u0_n106, u2_u9_u0_n107, 
       u2_u9_u0_n108, u2_u9_u0_n109, u2_u9_u0_n110, u2_u9_u0_n111, u2_u9_u0_n112, u2_u9_u0_n113, u2_u9_u0_n114, u2_u9_u0_n115, u2_u9_u0_n116, 
       u2_u9_u0_n117, u2_u9_u0_n118, u2_u9_u0_n119, u2_u9_u0_n120, u2_u9_u0_n121, u2_u9_u0_n122, u2_u9_u0_n123, u2_u9_u0_n124, u2_u9_u0_n125, 
       u2_u9_u0_n126, u2_u9_u0_n127, u2_u9_u0_n128, u2_u9_u0_n129, u2_u9_u0_n130, u2_u9_u0_n131, u2_u9_u0_n132, u2_u9_u0_n133, u2_u9_u0_n134, 
       u2_u9_u0_n135, u2_u9_u0_n136, u2_u9_u0_n137, u2_u9_u0_n138, u2_u9_u0_n139, u2_u9_u0_n140, u2_u9_u0_n141, u2_u9_u0_n142, u2_u9_u0_n143, 
       u2_u9_u0_n144, u2_u9_u0_n145, u2_u9_u0_n146, u2_u9_u0_n147, u2_u9_u0_n148, u2_u9_u0_n149, u2_u9_u0_n150, u2_u9_u0_n151, u2_u9_u0_n152, 
       u2_u9_u0_n153, u2_u9_u0_n154, u2_u9_u0_n155, u2_u9_u0_n156, u2_u9_u0_n157, u2_u9_u0_n158, u2_u9_u0_n159, u2_u9_u0_n160, u2_u9_u0_n161, 
       u2_u9_u0_n162, u2_u9_u0_n163, u2_u9_u0_n164, u2_u9_u0_n165, u2_u9_u0_n166, u2_u9_u0_n167, u2_u9_u0_n168, u2_u9_u0_n169, u2_u9_u0_n170, 
       u2_u9_u0_n171, u2_u9_u0_n172, u2_u9_u0_n173, u2_u9_u0_n174, u2_u9_u0_n88, u2_u9_u0_n89, u2_u9_u0_n90, u2_u9_u0_n91, u2_u9_u0_n92, 
       u2_u9_u0_n93, u2_u9_u0_n94, u2_u9_u0_n95, u2_u9_u0_n96, u2_u9_u0_n97, u2_u9_u0_n98, u2_u9_u0_n99, u2_u9_u5_n100, u2_u9_u5_n101, 
       u2_u9_u5_n102, u2_u9_u5_n103, u2_u9_u5_n104, u2_u9_u5_n105, u2_u9_u5_n106, u2_u9_u5_n107, u2_u9_u5_n108, u2_u9_u5_n109, u2_u9_u5_n110, 
       u2_u9_u5_n111, u2_u9_u5_n112, u2_u9_u5_n113, u2_u9_u5_n114, u2_u9_u5_n115, u2_u9_u5_n116, u2_u9_u5_n117, u2_u9_u5_n118, u2_u9_u5_n119, 
       u2_u9_u5_n120, u2_u9_u5_n121, u2_u9_u5_n122, u2_u9_u5_n123, u2_u9_u5_n124, u2_u9_u5_n125, u2_u9_u5_n126, u2_u9_u5_n127, u2_u9_u5_n128, 
       u2_u9_u5_n129, u2_u9_u5_n130, u2_u9_u5_n131, u2_u9_u5_n132, u2_u9_u5_n133, u2_u9_u5_n134, u2_u9_u5_n135, u2_u9_u5_n136, u2_u9_u5_n137, 
       u2_u9_u5_n138, u2_u9_u5_n139, u2_u9_u5_n140, u2_u9_u5_n141, u2_u9_u5_n142, u2_u9_u5_n143, u2_u9_u5_n144, u2_u9_u5_n145, u2_u9_u5_n146, 
       u2_u9_u5_n147, u2_u9_u5_n148, u2_u9_u5_n149, u2_u9_u5_n150, u2_u9_u5_n151, u2_u9_u5_n152, u2_u9_u5_n153, u2_u9_u5_n154, u2_u9_u5_n155, 
       u2_u9_u5_n156, u2_u9_u5_n157, u2_u9_u5_n158, u2_u9_u5_n159, u2_u9_u5_n160, u2_u9_u5_n161, u2_u9_u5_n162, u2_u9_u5_n163, u2_u9_u5_n164, 
       u2_u9_u5_n165, u2_u9_u5_n166, u2_u9_u5_n167, u2_u9_u5_n168, u2_u9_u5_n169, u2_u9_u5_n170, u2_u9_u5_n171, u2_u9_u5_n172, u2_u9_u5_n173, 
       u2_u9_u5_n174, u2_u9_u5_n175, u2_u9_u5_n176, u2_u9_u5_n177, u2_u9_u5_n178, u2_u9_u5_n179, u2_u9_u5_n180, u2_u9_u5_n181, u2_u9_u5_n182, 
       u2_u9_u5_n183, u2_u9_u5_n184, u2_u9_u5_n185, u2_u9_u5_n186, u2_u9_u5_n187, u2_u9_u5_n188, u2_u9_u5_n189, u2_u9_u5_n190, u2_u9_u5_n191, 
       u2_u9_u5_n192, u2_u9_u5_n193, u2_u9_u5_n194, u2_u9_u5_n195, u2_u9_u5_n196, u2_u9_u5_n99, u2_u9_u6_n100, u2_u9_u6_n101, u2_u9_u6_n102, 
       u2_u9_u6_n103, u2_u9_u6_n104, u2_u9_u6_n105, u2_u9_u6_n106, u2_u9_u6_n107, u2_u9_u6_n108, u2_u9_u6_n109, u2_u9_u6_n110, u2_u9_u6_n111, 
       u2_u9_u6_n112, u2_u9_u6_n113, u2_u9_u6_n114, u2_u9_u6_n115, u2_u9_u6_n116, u2_u9_u6_n117, u2_u9_u6_n118, u2_u9_u6_n119, u2_u9_u6_n120, 
       u2_u9_u6_n121, u2_u9_u6_n122, u2_u9_u6_n123, u2_u9_u6_n124, u2_u9_u6_n125, u2_u9_u6_n126, u2_u9_u6_n127, u2_u9_u6_n128, u2_u9_u6_n129, 
       u2_u9_u6_n130, u2_u9_u6_n131, u2_u9_u6_n132, u2_u9_u6_n133, u2_u9_u6_n134, u2_u9_u6_n135, u2_u9_u6_n136, u2_u9_u6_n137, u2_u9_u6_n138, 
       u2_u9_u6_n139, u2_u9_u6_n140, u2_u9_u6_n141, u2_u9_u6_n142, u2_u9_u6_n143, u2_u9_u6_n144, u2_u9_u6_n145, u2_u9_u6_n146, u2_u9_u6_n147, 
       u2_u9_u6_n148, u2_u9_u6_n149, u2_u9_u6_n150, u2_u9_u6_n151, u2_u9_u6_n152, u2_u9_u6_n153, u2_u9_u6_n154, u2_u9_u6_n155, u2_u9_u6_n156, 
       u2_u9_u6_n157, u2_u9_u6_n158, u2_u9_u6_n159, u2_u9_u6_n160, u2_u9_u6_n161, u2_u9_u6_n162, u2_u9_u6_n163, u2_u9_u6_n164, u2_u9_u6_n165, 
       u2_u9_u6_n166, u2_u9_u6_n167, u2_u9_u6_n168, u2_u9_u6_n169, u2_u9_u6_n170, u2_u9_u6_n171, u2_u9_u6_n172, u2_u9_u6_n173, u2_u9_u6_n174, 
       u2_u9_u6_n88, u2_u9_u6_n89, u2_u9_u6_n90, u2_u9_u6_n91, u2_u9_u6_n92, u2_u9_u6_n93, u2_u9_u6_n94, u2_u9_u6_n95, u2_u9_u6_n96, 
       u2_u9_u6_n97, u2_u9_u6_n98, u2_u9_u6_n99, u2_u9_u7_n100, u2_u9_u7_n101, u2_u9_u7_n102, u2_u9_u7_n103, u2_u9_u7_n104, u2_u9_u7_n105, 
       u2_u9_u7_n106, u2_u9_u7_n107, u2_u9_u7_n108, u2_u9_u7_n109, u2_u9_u7_n110, u2_u9_u7_n111, u2_u9_u7_n112, u2_u9_u7_n113, u2_u9_u7_n114, 
       u2_u9_u7_n115, u2_u9_u7_n116, u2_u9_u7_n117, u2_u9_u7_n118, u2_u9_u7_n119, u2_u9_u7_n120, u2_u9_u7_n121, u2_u9_u7_n122, u2_u9_u7_n123, 
       u2_u9_u7_n124, u2_u9_u7_n125, u2_u9_u7_n126, u2_u9_u7_n127, u2_u9_u7_n128, u2_u9_u7_n129, u2_u9_u7_n130, u2_u9_u7_n131, u2_u9_u7_n132, 
       u2_u9_u7_n133, u2_u9_u7_n134, u2_u9_u7_n135, u2_u9_u7_n136, u2_u9_u7_n137, u2_u9_u7_n138, u2_u9_u7_n139, u2_u9_u7_n140, u2_u9_u7_n141, 
       u2_u9_u7_n142, u2_u9_u7_n143, u2_u9_u7_n144, u2_u9_u7_n145, u2_u9_u7_n146, u2_u9_u7_n147, u2_u9_u7_n148, u2_u9_u7_n149, u2_u9_u7_n150, 
       u2_u9_u7_n151, u2_u9_u7_n152, u2_u9_u7_n153, u2_u9_u7_n154, u2_u9_u7_n155, u2_u9_u7_n156, u2_u9_u7_n157, u2_u9_u7_n158, u2_u9_u7_n159, 
       u2_u9_u7_n160, u2_u9_u7_n161, u2_u9_u7_n162, u2_u9_u7_n163, u2_u9_u7_n164, u2_u9_u7_n165, u2_u9_u7_n166, u2_u9_u7_n167, u2_u9_u7_n168, 
       u2_u9_u7_n169, u2_u9_u7_n170, u2_u9_u7_n171, u2_u9_u7_n172, u2_u9_u7_n173, u2_u9_u7_n174, u2_u9_u7_n175, u2_u9_u7_n176, u2_u9_u7_n177, 
       u2_u9_u7_n178, u2_u9_u7_n179, u2_u9_u7_n180, u2_u9_u7_n91, u2_u9_u7_n92, u2_u9_u7_n93, u2_u9_u7_n94, u2_u9_u7_n95, u2_u9_u7_n96, 
       u2_u9_u7_n97, u2_u9_u7_n98, u2_u9_u7_n99, u2_uk_n1013, u2_uk_n1014, u2_uk_n1015, u2_uk_n1016, u2_uk_n1017, u2_uk_n1019, 
       u2_uk_n1021, u2_uk_n1023, u2_uk_n1026, u2_uk_n1029, u2_uk_n1030, u2_uk_n1032, u2_uk_n1033, u2_uk_n1037, u2_uk_n1041, 
       u2_uk_n1048, u2_uk_n1052, u2_uk_n1054, u2_uk_n1057, u2_uk_n1059, u2_uk_n1060, u2_uk_n1062, u2_uk_n1064, u2_uk_n1066, 
       u2_uk_n1068, u2_uk_n1072, u2_uk_n1075, u2_uk_n1078, u2_uk_n1080, u2_uk_n1086, u2_uk_n1095, u2_uk_n1117, u2_uk_n1118, 
       u2_uk_n1122, u2_uk_n1126, u2_uk_n1127, u2_uk_n1147, u2_uk_n1151, u2_uk_n1158, u2_uk_n1165, u2_uk_n286, u2_uk_n291, 
       u2_uk_n294, u2_uk_n297, u2_uk_n306, u2_uk_n338, u2_uk_n342, u2_uk_n671, u2_uk_n678, u2_uk_n936,  u2_uk_n938;
  XOR2_X1 u0_u12_U25 (.B( u0_K13_31 ) , .A( u0_R11_20 ) , .Z( u0_u12_X_31 ) );
  XOR2_X1 u0_u12_U28 (.B( u0_K13_29 ) , .A( u0_R11_20 ) , .Z( u0_u12_X_29 ) );
  XOR2_X1 u0_u12_U32 (.B( u0_K13_25 ) , .A( u0_R11_16 ) , .Z( u0_u12_X_25 ) );
  OAI22_X1 u0_u12_u4_U10 (.B2( u0_u12_u4_n135 ) , .ZN( u0_u12_u4_n137 ) , .B1( u0_u12_u4_n153 ) , .A1( u0_u12_u4_n155 ) , .A2( u0_u12_u4_n171 ) );
  AND3_X1 u0_u12_u4_U11 (.A2( u0_u12_u4_n134 ) , .ZN( u0_u12_u4_n135 ) , .A3( u0_u12_u4_n145 ) , .A1( u0_u12_u4_n157 ) );
  NAND2_X1 u0_u12_u4_U12 (.ZN( u0_u12_u4_n132 ) , .A2( u0_u12_u4_n170 ) , .A1( u0_u12_u4_n173 ) );
  AOI21_X1 u0_u12_u4_U13 (.B2( u0_u12_u4_n160 ) , .B1( u0_u12_u4_n161 ) , .ZN( u0_u12_u4_n162 ) , .A( u0_u12_u4_n170 ) );
  AOI21_X1 u0_u12_u4_U14 (.ZN( u0_u12_u4_n107 ) , .B2( u0_u12_u4_n143 ) , .A( u0_u12_u4_n174 ) , .B1( u0_u12_u4_n184 ) );
  AOI21_X1 u0_u12_u4_U15 (.B2( u0_u12_u4_n158 ) , .B1( u0_u12_u4_n159 ) , .ZN( u0_u12_u4_n163 ) , .A( u0_u12_u4_n174 ) );
  AOI21_X1 u0_u12_u4_U16 (.A( u0_u12_u4_n153 ) , .B2( u0_u12_u4_n154 ) , .B1( u0_u12_u4_n155 ) , .ZN( u0_u12_u4_n165 ) );
  AOI21_X1 u0_u12_u4_U17 (.A( u0_u12_u4_n156 ) , .B2( u0_u12_u4_n157 ) , .ZN( u0_u12_u4_n164 ) , .B1( u0_u12_u4_n184 ) );
  INV_X1 u0_u12_u4_U18 (.A( u0_u12_u4_n138 ) , .ZN( u0_u12_u4_n170 ) );
  AND2_X1 u0_u12_u4_U19 (.A2( u0_u12_u4_n120 ) , .ZN( u0_u12_u4_n155 ) , .A1( u0_u12_u4_n160 ) );
  INV_X1 u0_u12_u4_U20 (.A( u0_u12_u4_n156 ) , .ZN( u0_u12_u4_n175 ) );
  NAND2_X1 u0_u12_u4_U21 (.A2( u0_u12_u4_n118 ) , .ZN( u0_u12_u4_n131 ) , .A1( u0_u12_u4_n147 ) );
  NAND2_X1 u0_u12_u4_U22 (.A1( u0_u12_u4_n119 ) , .A2( u0_u12_u4_n120 ) , .ZN( u0_u12_u4_n130 ) );
  NAND2_X1 u0_u12_u4_U23 (.ZN( u0_u12_u4_n117 ) , .A2( u0_u12_u4_n118 ) , .A1( u0_u12_u4_n148 ) );
  NAND2_X1 u0_u12_u4_U24 (.ZN( u0_u12_u4_n129 ) , .A1( u0_u12_u4_n134 ) , .A2( u0_u12_u4_n148 ) );
  AND3_X1 u0_u12_u4_U25 (.A1( u0_u12_u4_n119 ) , .A2( u0_u12_u4_n143 ) , .A3( u0_u12_u4_n154 ) , .ZN( u0_u12_u4_n161 ) );
  AND2_X1 u0_u12_u4_U26 (.A1( u0_u12_u4_n145 ) , .A2( u0_u12_u4_n147 ) , .ZN( u0_u12_u4_n159 ) );
  OR3_X1 u0_u12_u4_U27 (.A3( u0_u12_u4_n114 ) , .A2( u0_u12_u4_n115 ) , .A1( u0_u12_u4_n116 ) , .ZN( u0_u12_u4_n136 ) );
  AOI21_X1 u0_u12_u4_U28 (.A( u0_u12_u4_n113 ) , .ZN( u0_u12_u4_n116 ) , .B2( u0_u12_u4_n173 ) , .B1( u0_u12_u4_n174 ) );
  AOI21_X1 u0_u12_u4_U29 (.ZN( u0_u12_u4_n115 ) , .B2( u0_u12_u4_n145 ) , .B1( u0_u12_u4_n146 ) , .A( u0_u12_u4_n156 ) );
  NOR2_X1 u0_u12_u4_U3 (.ZN( u0_u12_u4_n121 ) , .A1( u0_u12_u4_n181 ) , .A2( u0_u12_u4_n182 ) );
  OAI22_X1 u0_u12_u4_U30 (.ZN( u0_u12_u4_n114 ) , .A2( u0_u12_u4_n121 ) , .B1( u0_u12_u4_n160 ) , .B2( u0_u12_u4_n170 ) , .A1( u0_u12_u4_n171 ) );
  INV_X1 u0_u12_u4_U31 (.A( u0_u12_u4_n158 ) , .ZN( u0_u12_u4_n182 ) );
  INV_X1 u0_u12_u4_U32 (.ZN( u0_u12_u4_n181 ) , .A( u0_u12_u4_n96 ) );
  INV_X1 u0_u12_u4_U33 (.A( u0_u12_u4_n144 ) , .ZN( u0_u12_u4_n179 ) );
  INV_X1 u0_u12_u4_U34 (.A( u0_u12_u4_n157 ) , .ZN( u0_u12_u4_n178 ) );
  NAND2_X1 u0_u12_u4_U35 (.A2( u0_u12_u4_n154 ) , .A1( u0_u12_u4_n96 ) , .ZN( u0_u12_u4_n97 ) );
  INV_X1 u0_u12_u4_U36 (.ZN( u0_u12_u4_n186 ) , .A( u0_u12_u4_n95 ) );
  OAI221_X1 u0_u12_u4_U37 (.C1( u0_u12_u4_n134 ) , .B1( u0_u12_u4_n158 ) , .B2( u0_u12_u4_n171 ) , .C2( u0_u12_u4_n173 ) , .A( u0_u12_u4_n94 ) , .ZN( u0_u12_u4_n95 ) );
  AOI222_X1 u0_u12_u4_U38 (.B2( u0_u12_u4_n132 ) , .A1( u0_u12_u4_n138 ) , .C2( u0_u12_u4_n175 ) , .A2( u0_u12_u4_n179 ) , .C1( u0_u12_u4_n181 ) , .B1( u0_u12_u4_n185 ) , .ZN( u0_u12_u4_n94 ) );
  INV_X1 u0_u12_u4_U39 (.A( u0_u12_u4_n113 ) , .ZN( u0_u12_u4_n185 ) );
  INV_X1 u0_u12_u4_U4 (.A( u0_u12_u4_n117 ) , .ZN( u0_u12_u4_n184 ) );
  INV_X1 u0_u12_u4_U40 (.A( u0_u12_u4_n143 ) , .ZN( u0_u12_u4_n183 ) );
  NOR2_X1 u0_u12_u4_U41 (.ZN( u0_u12_u4_n138 ) , .A1( u0_u12_u4_n168 ) , .A2( u0_u12_u4_n169 ) );
  NOR2_X1 u0_u12_u4_U42 (.A1( u0_u12_u4_n150 ) , .A2( u0_u12_u4_n152 ) , .ZN( u0_u12_u4_n153 ) );
  NOR2_X1 u0_u12_u4_U43 (.A2( u0_u12_u4_n128 ) , .A1( u0_u12_u4_n138 ) , .ZN( u0_u12_u4_n156 ) );
  AOI22_X1 u0_u12_u4_U44 (.B2( u0_u12_u4_n122 ) , .A1( u0_u12_u4_n123 ) , .ZN( u0_u12_u4_n124 ) , .B1( u0_u12_u4_n128 ) , .A2( u0_u12_u4_n172 ) );
  INV_X1 u0_u12_u4_U45 (.A( u0_u12_u4_n153 ) , .ZN( u0_u12_u4_n172 ) );
  NAND2_X1 u0_u12_u4_U46 (.A2( u0_u12_u4_n120 ) , .ZN( u0_u12_u4_n123 ) , .A1( u0_u12_u4_n161 ) );
  AOI22_X1 u0_u12_u4_U47 (.B2( u0_u12_u4_n132 ) , .A2( u0_u12_u4_n133 ) , .ZN( u0_u12_u4_n140 ) , .A1( u0_u12_u4_n150 ) , .B1( u0_u12_u4_n179 ) );
  NAND2_X1 u0_u12_u4_U48 (.ZN( u0_u12_u4_n133 ) , .A2( u0_u12_u4_n146 ) , .A1( u0_u12_u4_n154 ) );
  NAND2_X1 u0_u12_u4_U49 (.A1( u0_u12_u4_n103 ) , .ZN( u0_u12_u4_n154 ) , .A2( u0_u12_u4_n98 ) );
  NOR4_X1 u0_u12_u4_U5 (.A4( u0_u12_u4_n106 ) , .A3( u0_u12_u4_n107 ) , .A2( u0_u12_u4_n108 ) , .A1( u0_u12_u4_n109 ) , .ZN( u0_u12_u4_n110 ) );
  NAND2_X1 u0_u12_u4_U50 (.A1( u0_u12_u4_n101 ) , .ZN( u0_u12_u4_n158 ) , .A2( u0_u12_u4_n99 ) );
  AOI21_X1 u0_u12_u4_U51 (.ZN( u0_u12_u4_n127 ) , .A( u0_u12_u4_n136 ) , .B2( u0_u12_u4_n150 ) , .B1( u0_u12_u4_n180 ) );
  INV_X1 u0_u12_u4_U52 (.A( u0_u12_u4_n160 ) , .ZN( u0_u12_u4_n180 ) );
  NAND2_X1 u0_u12_u4_U53 (.A2( u0_u12_u4_n104 ) , .A1( u0_u12_u4_n105 ) , .ZN( u0_u12_u4_n146 ) );
  NAND2_X1 u0_u12_u4_U54 (.A2( u0_u12_u4_n101 ) , .A1( u0_u12_u4_n102 ) , .ZN( u0_u12_u4_n160 ) );
  NAND2_X1 u0_u12_u4_U55 (.ZN( u0_u12_u4_n134 ) , .A1( u0_u12_u4_n98 ) , .A2( u0_u12_u4_n99 ) );
  NAND2_X1 u0_u12_u4_U56 (.A1( u0_u12_u4_n103 ) , .A2( u0_u12_u4_n104 ) , .ZN( u0_u12_u4_n143 ) );
  NAND2_X1 u0_u12_u4_U57 (.A2( u0_u12_u4_n105 ) , .ZN( u0_u12_u4_n145 ) , .A1( u0_u12_u4_n98 ) );
  NAND2_X1 u0_u12_u4_U58 (.A1( u0_u12_u4_n100 ) , .A2( u0_u12_u4_n105 ) , .ZN( u0_u12_u4_n120 ) );
  NAND2_X1 u0_u12_u4_U59 (.A1( u0_u12_u4_n102 ) , .A2( u0_u12_u4_n104 ) , .ZN( u0_u12_u4_n148 ) );
  AOI21_X1 u0_u12_u4_U6 (.ZN( u0_u12_u4_n106 ) , .B2( u0_u12_u4_n146 ) , .B1( u0_u12_u4_n158 ) , .A( u0_u12_u4_n170 ) );
  NAND2_X1 u0_u12_u4_U60 (.A2( u0_u12_u4_n100 ) , .A1( u0_u12_u4_n103 ) , .ZN( u0_u12_u4_n157 ) );
  INV_X1 u0_u12_u4_U61 (.A( u0_u12_u4_n150 ) , .ZN( u0_u12_u4_n173 ) );
  INV_X1 u0_u12_u4_U62 (.A( u0_u12_u4_n152 ) , .ZN( u0_u12_u4_n171 ) );
  NAND2_X1 u0_u12_u4_U63 (.A1( u0_u12_u4_n100 ) , .ZN( u0_u12_u4_n118 ) , .A2( u0_u12_u4_n99 ) );
  NAND2_X1 u0_u12_u4_U64 (.A2( u0_u12_u4_n100 ) , .A1( u0_u12_u4_n102 ) , .ZN( u0_u12_u4_n144 ) );
  NAND2_X1 u0_u12_u4_U65 (.A2( u0_u12_u4_n101 ) , .A1( u0_u12_u4_n105 ) , .ZN( u0_u12_u4_n96 ) );
  INV_X1 u0_u12_u4_U66 (.A( u0_u12_u4_n128 ) , .ZN( u0_u12_u4_n174 ) );
  NAND2_X1 u0_u12_u4_U67 (.A2( u0_u12_u4_n102 ) , .ZN( u0_u12_u4_n119 ) , .A1( u0_u12_u4_n98 ) );
  NAND2_X1 u0_u12_u4_U68 (.A2( u0_u12_u4_n101 ) , .A1( u0_u12_u4_n103 ) , .ZN( u0_u12_u4_n147 ) );
  NAND2_X1 u0_u12_u4_U69 (.A2( u0_u12_u4_n104 ) , .ZN( u0_u12_u4_n113 ) , .A1( u0_u12_u4_n99 ) );
  AOI21_X1 u0_u12_u4_U7 (.ZN( u0_u12_u4_n108 ) , .B2( u0_u12_u4_n134 ) , .B1( u0_u12_u4_n155 ) , .A( u0_u12_u4_n156 ) );
  NOR2_X1 u0_u12_u4_U70 (.A2( u0_u12_X_28 ) , .ZN( u0_u12_u4_n150 ) , .A1( u0_u12_u4_n168 ) );
  NOR2_X1 u0_u12_u4_U71 (.A2( u0_u12_X_29 ) , .ZN( u0_u12_u4_n152 ) , .A1( u0_u12_u4_n169 ) );
  NOR2_X1 u0_u12_u4_U72 (.A2( u0_u12_X_30 ) , .ZN( u0_u12_u4_n105 ) , .A1( u0_u12_u4_n176 ) );
  NOR2_X1 u0_u12_u4_U73 (.A2( u0_u12_X_26 ) , .ZN( u0_u12_u4_n100 ) , .A1( u0_u12_u4_n177 ) );
  NOR2_X1 u0_u12_u4_U74 (.A2( u0_u12_X_28 ) , .A1( u0_u12_X_29 ) , .ZN( u0_u12_u4_n128 ) );
  NOR2_X1 u0_u12_u4_U75 (.A2( u0_u12_X_27 ) , .A1( u0_u12_X_30 ) , .ZN( u0_u12_u4_n102 ) );
  NOR2_X1 u0_u12_u4_U76 (.A2( u0_u12_X_25 ) , .A1( u0_u12_X_26 ) , .ZN( u0_u12_u4_n98 ) );
  AND2_X1 u0_u12_u4_U77 (.A2( u0_u12_X_25 ) , .A1( u0_u12_X_26 ) , .ZN( u0_u12_u4_n104 ) );
  AND2_X1 u0_u12_u4_U78 (.A1( u0_u12_X_30 ) , .A2( u0_u12_u4_n176 ) , .ZN( u0_u12_u4_n99 ) );
  AND2_X1 u0_u12_u4_U79 (.A1( u0_u12_X_26 ) , .ZN( u0_u12_u4_n101 ) , .A2( u0_u12_u4_n177 ) );
  AOI21_X1 u0_u12_u4_U8 (.ZN( u0_u12_u4_n109 ) , .A( u0_u12_u4_n153 ) , .B1( u0_u12_u4_n159 ) , .B2( u0_u12_u4_n184 ) );
  AND2_X1 u0_u12_u4_U80 (.A1( u0_u12_X_27 ) , .A2( u0_u12_X_30 ) , .ZN( u0_u12_u4_n103 ) );
  INV_X1 u0_u12_u4_U81 (.A( u0_u12_X_28 ) , .ZN( u0_u12_u4_n169 ) );
  INV_X1 u0_u12_u4_U82 (.A( u0_u12_X_29 ) , .ZN( u0_u12_u4_n168 ) );
  INV_X1 u0_u12_u4_U83 (.A( u0_u12_X_25 ) , .ZN( u0_u12_u4_n177 ) );
  INV_X1 u0_u12_u4_U84 (.A( u0_u12_X_27 ) , .ZN( u0_u12_u4_n176 ) );
  NAND4_X1 u0_u12_u4_U85 (.ZN( u0_out12_25 ) , .A4( u0_u12_u4_n139 ) , .A3( u0_u12_u4_n140 ) , .A2( u0_u12_u4_n141 ) , .A1( u0_u12_u4_n142 ) );
  OAI21_X1 u0_u12_u4_U86 (.A( u0_u12_u4_n128 ) , .B2( u0_u12_u4_n129 ) , .B1( u0_u12_u4_n130 ) , .ZN( u0_u12_u4_n142 ) );
  OAI21_X1 u0_u12_u4_U87 (.B2( u0_u12_u4_n131 ) , .ZN( u0_u12_u4_n141 ) , .A( u0_u12_u4_n175 ) , .B1( u0_u12_u4_n183 ) );
  NAND4_X1 u0_u12_u4_U88 (.ZN( u0_out12_14 ) , .A4( u0_u12_u4_n124 ) , .A3( u0_u12_u4_n125 ) , .A2( u0_u12_u4_n126 ) , .A1( u0_u12_u4_n127 ) );
  AOI22_X1 u0_u12_u4_U89 (.B2( u0_u12_u4_n117 ) , .ZN( u0_u12_u4_n126 ) , .A1( u0_u12_u4_n129 ) , .B1( u0_u12_u4_n152 ) , .A2( u0_u12_u4_n175 ) );
  AOI211_X1 u0_u12_u4_U9 (.B( u0_u12_u4_n136 ) , .A( u0_u12_u4_n137 ) , .C2( u0_u12_u4_n138 ) , .ZN( u0_u12_u4_n139 ) , .C1( u0_u12_u4_n182 ) );
  AOI22_X1 u0_u12_u4_U90 (.ZN( u0_u12_u4_n125 ) , .B2( u0_u12_u4_n131 ) , .A2( u0_u12_u4_n132 ) , .B1( u0_u12_u4_n138 ) , .A1( u0_u12_u4_n178 ) );
  NAND4_X1 u0_u12_u4_U91 (.ZN( u0_out12_8 ) , .A4( u0_u12_u4_n110 ) , .A3( u0_u12_u4_n111 ) , .A2( u0_u12_u4_n112 ) , .A1( u0_u12_u4_n186 ) );
  NAND2_X1 u0_u12_u4_U92 (.ZN( u0_u12_u4_n112 ) , .A2( u0_u12_u4_n130 ) , .A1( u0_u12_u4_n150 ) );
  AOI22_X1 u0_u12_u4_U93 (.ZN( u0_u12_u4_n111 ) , .B2( u0_u12_u4_n132 ) , .A1( u0_u12_u4_n152 ) , .B1( u0_u12_u4_n178 ) , .A2( u0_u12_u4_n97 ) );
  AOI22_X1 u0_u12_u4_U94 (.B2( u0_u12_u4_n149 ) , .B1( u0_u12_u4_n150 ) , .A2( u0_u12_u4_n151 ) , .A1( u0_u12_u4_n152 ) , .ZN( u0_u12_u4_n167 ) );
  NOR4_X1 u0_u12_u4_U95 (.A4( u0_u12_u4_n162 ) , .A3( u0_u12_u4_n163 ) , .A2( u0_u12_u4_n164 ) , .A1( u0_u12_u4_n165 ) , .ZN( u0_u12_u4_n166 ) );
  NAND3_X1 u0_u12_u4_U96 (.ZN( u0_out12_3 ) , .A3( u0_u12_u4_n166 ) , .A1( u0_u12_u4_n167 ) , .A2( u0_u12_u4_n186 ) );
  NAND3_X1 u0_u12_u4_U97 (.A3( u0_u12_u4_n146 ) , .A2( u0_u12_u4_n147 ) , .A1( u0_u12_u4_n148 ) , .ZN( u0_u12_u4_n149 ) );
  NAND3_X1 u0_u12_u4_U98 (.A3( u0_u12_u4_n143 ) , .A2( u0_u12_u4_n144 ) , .A1( u0_u12_u4_n145 ) , .ZN( u0_u12_u4_n151 ) );
  NAND3_X1 u0_u12_u4_U99 (.A3( u0_u12_u4_n121 ) , .ZN( u0_u12_u4_n122 ) , .A2( u0_u12_u4_n144 ) , .A1( u0_u12_u4_n154 ) );
  INV_X1 u0_u12_u5_U10 (.A( u0_u12_u5_n121 ) , .ZN( u0_u12_u5_n177 ) );
  NOR3_X1 u0_u12_u5_U100 (.A3( u0_u12_u5_n141 ) , .A1( u0_u12_u5_n142 ) , .ZN( u0_u12_u5_n143 ) , .A2( u0_u12_u5_n191 ) );
  NAND4_X1 u0_u12_u5_U101 (.ZN( u0_out12_4 ) , .A4( u0_u12_u5_n112 ) , .A2( u0_u12_u5_n113 ) , .A1( u0_u12_u5_n114 ) , .A3( u0_u12_u5_n195 ) );
  AOI211_X1 u0_u12_u5_U102 (.A( u0_u12_u5_n110 ) , .C1( u0_u12_u5_n111 ) , .ZN( u0_u12_u5_n112 ) , .B( u0_u12_u5_n118 ) , .C2( u0_u12_u5_n177 ) );
  AOI222_X1 u0_u12_u5_U103 (.ZN( u0_u12_u5_n113 ) , .A1( u0_u12_u5_n131 ) , .C1( u0_u12_u5_n148 ) , .B2( u0_u12_u5_n174 ) , .C2( u0_u12_u5_n178 ) , .A2( u0_u12_u5_n179 ) , .B1( u0_u12_u5_n99 ) );
  NAND3_X1 u0_u12_u5_U104 (.A2( u0_u12_u5_n154 ) , .A3( u0_u12_u5_n158 ) , .A1( u0_u12_u5_n161 ) , .ZN( u0_u12_u5_n99 ) );
  NOR2_X1 u0_u12_u5_U11 (.ZN( u0_u12_u5_n160 ) , .A2( u0_u12_u5_n173 ) , .A1( u0_u12_u5_n177 ) );
  INV_X1 u0_u12_u5_U12 (.A( u0_u12_u5_n150 ) , .ZN( u0_u12_u5_n174 ) );
  AOI21_X1 u0_u12_u5_U13 (.A( u0_u12_u5_n160 ) , .B2( u0_u12_u5_n161 ) , .ZN( u0_u12_u5_n162 ) , .B1( u0_u12_u5_n192 ) );
  INV_X1 u0_u12_u5_U14 (.A( u0_u12_u5_n159 ) , .ZN( u0_u12_u5_n192 ) );
  AOI21_X1 u0_u12_u5_U15 (.A( u0_u12_u5_n156 ) , .B2( u0_u12_u5_n157 ) , .B1( u0_u12_u5_n158 ) , .ZN( u0_u12_u5_n163 ) );
  AOI21_X1 u0_u12_u5_U16 (.B2( u0_u12_u5_n139 ) , .B1( u0_u12_u5_n140 ) , .ZN( u0_u12_u5_n141 ) , .A( u0_u12_u5_n150 ) );
  OAI21_X1 u0_u12_u5_U17 (.A( u0_u12_u5_n133 ) , .B2( u0_u12_u5_n134 ) , .B1( u0_u12_u5_n135 ) , .ZN( u0_u12_u5_n142 ) );
  OAI21_X1 u0_u12_u5_U18 (.ZN( u0_u12_u5_n133 ) , .B2( u0_u12_u5_n147 ) , .A( u0_u12_u5_n173 ) , .B1( u0_u12_u5_n188 ) );
  NAND2_X1 u0_u12_u5_U19 (.A2( u0_u12_u5_n119 ) , .A1( u0_u12_u5_n123 ) , .ZN( u0_u12_u5_n137 ) );
  INV_X1 u0_u12_u5_U20 (.A( u0_u12_u5_n155 ) , .ZN( u0_u12_u5_n194 ) );
  NAND2_X1 u0_u12_u5_U21 (.A1( u0_u12_u5_n121 ) , .ZN( u0_u12_u5_n132 ) , .A2( u0_u12_u5_n172 ) );
  NAND2_X1 u0_u12_u5_U22 (.A2( u0_u12_u5_n122 ) , .ZN( u0_u12_u5_n136 ) , .A1( u0_u12_u5_n154 ) );
  NAND2_X1 u0_u12_u5_U23 (.A2( u0_u12_u5_n119 ) , .A1( u0_u12_u5_n120 ) , .ZN( u0_u12_u5_n159 ) );
  INV_X1 u0_u12_u5_U24 (.A( u0_u12_u5_n156 ) , .ZN( u0_u12_u5_n175 ) );
  INV_X1 u0_u12_u5_U25 (.A( u0_u12_u5_n158 ) , .ZN( u0_u12_u5_n188 ) );
  INV_X1 u0_u12_u5_U26 (.A( u0_u12_u5_n152 ) , .ZN( u0_u12_u5_n179 ) );
  INV_X1 u0_u12_u5_U27 (.A( u0_u12_u5_n140 ) , .ZN( u0_u12_u5_n182 ) );
  INV_X1 u0_u12_u5_U28 (.A( u0_u12_u5_n151 ) , .ZN( u0_u12_u5_n183 ) );
  INV_X1 u0_u12_u5_U29 (.A( u0_u12_u5_n123 ) , .ZN( u0_u12_u5_n185 ) );
  NOR2_X1 u0_u12_u5_U3 (.ZN( u0_u12_u5_n134 ) , .A1( u0_u12_u5_n183 ) , .A2( u0_u12_u5_n190 ) );
  INV_X1 u0_u12_u5_U30 (.A( u0_u12_u5_n161 ) , .ZN( u0_u12_u5_n184 ) );
  INV_X1 u0_u12_u5_U31 (.A( u0_u12_u5_n139 ) , .ZN( u0_u12_u5_n189 ) );
  INV_X1 u0_u12_u5_U32 (.A( u0_u12_u5_n157 ) , .ZN( u0_u12_u5_n190 ) );
  INV_X1 u0_u12_u5_U33 (.A( u0_u12_u5_n120 ) , .ZN( u0_u12_u5_n193 ) );
  NAND2_X1 u0_u12_u5_U34 (.ZN( u0_u12_u5_n111 ) , .A1( u0_u12_u5_n140 ) , .A2( u0_u12_u5_n155 ) );
  NOR2_X1 u0_u12_u5_U35 (.ZN( u0_u12_u5_n100 ) , .A1( u0_u12_u5_n170 ) , .A2( u0_u12_u5_n180 ) );
  INV_X1 u0_u12_u5_U36 (.A( u0_u12_u5_n117 ) , .ZN( u0_u12_u5_n196 ) );
  OAI221_X1 u0_u12_u5_U37 (.A( u0_u12_u5_n116 ) , .ZN( u0_u12_u5_n117 ) , .B2( u0_u12_u5_n119 ) , .C1( u0_u12_u5_n153 ) , .C2( u0_u12_u5_n158 ) , .B1( u0_u12_u5_n172 ) );
  AOI222_X1 u0_u12_u5_U38 (.ZN( u0_u12_u5_n116 ) , .B2( u0_u12_u5_n145 ) , .C1( u0_u12_u5_n148 ) , .A2( u0_u12_u5_n174 ) , .C2( u0_u12_u5_n177 ) , .B1( u0_u12_u5_n187 ) , .A1( u0_u12_u5_n193 ) );
  INV_X1 u0_u12_u5_U39 (.A( u0_u12_u5_n115 ) , .ZN( u0_u12_u5_n187 ) );
  INV_X1 u0_u12_u5_U4 (.A( u0_u12_u5_n138 ) , .ZN( u0_u12_u5_n191 ) );
  AOI22_X1 u0_u12_u5_U40 (.B2( u0_u12_u5_n131 ) , .A2( u0_u12_u5_n146 ) , .ZN( u0_u12_u5_n169 ) , .B1( u0_u12_u5_n174 ) , .A1( u0_u12_u5_n185 ) );
  NOR2_X1 u0_u12_u5_U41 (.A1( u0_u12_u5_n146 ) , .ZN( u0_u12_u5_n150 ) , .A2( u0_u12_u5_n173 ) );
  AOI21_X1 u0_u12_u5_U42 (.A( u0_u12_u5_n118 ) , .B2( u0_u12_u5_n145 ) , .ZN( u0_u12_u5_n168 ) , .B1( u0_u12_u5_n186 ) );
  INV_X1 u0_u12_u5_U43 (.A( u0_u12_u5_n122 ) , .ZN( u0_u12_u5_n186 ) );
  NOR2_X1 u0_u12_u5_U44 (.A1( u0_u12_u5_n146 ) , .ZN( u0_u12_u5_n152 ) , .A2( u0_u12_u5_n176 ) );
  NOR2_X1 u0_u12_u5_U45 (.A1( u0_u12_u5_n115 ) , .ZN( u0_u12_u5_n118 ) , .A2( u0_u12_u5_n153 ) );
  NOR2_X1 u0_u12_u5_U46 (.A2( u0_u12_u5_n145 ) , .ZN( u0_u12_u5_n156 ) , .A1( u0_u12_u5_n174 ) );
  NOR2_X1 u0_u12_u5_U47 (.ZN( u0_u12_u5_n121 ) , .A2( u0_u12_u5_n145 ) , .A1( u0_u12_u5_n176 ) );
  AOI22_X1 u0_u12_u5_U48 (.ZN( u0_u12_u5_n114 ) , .A2( u0_u12_u5_n137 ) , .A1( u0_u12_u5_n145 ) , .B2( u0_u12_u5_n175 ) , .B1( u0_u12_u5_n193 ) );
  OAI211_X1 u0_u12_u5_U49 (.B( u0_u12_u5_n124 ) , .A( u0_u12_u5_n125 ) , .C2( u0_u12_u5_n126 ) , .C1( u0_u12_u5_n127 ) , .ZN( u0_u12_u5_n128 ) );
  OAI21_X1 u0_u12_u5_U5 (.B2( u0_u12_u5_n136 ) , .B1( u0_u12_u5_n137 ) , .ZN( u0_u12_u5_n138 ) , .A( u0_u12_u5_n177 ) );
  NOR3_X1 u0_u12_u5_U50 (.ZN( u0_u12_u5_n127 ) , .A1( u0_u12_u5_n136 ) , .A3( u0_u12_u5_n148 ) , .A2( u0_u12_u5_n182 ) );
  OAI21_X1 u0_u12_u5_U51 (.ZN( u0_u12_u5_n124 ) , .A( u0_u12_u5_n177 ) , .B2( u0_u12_u5_n183 ) , .B1( u0_u12_u5_n189 ) );
  OAI21_X1 u0_u12_u5_U52 (.ZN( u0_u12_u5_n125 ) , .A( u0_u12_u5_n174 ) , .B2( u0_u12_u5_n185 ) , .B1( u0_u12_u5_n190 ) );
  AOI21_X1 u0_u12_u5_U53 (.A( u0_u12_u5_n153 ) , .B2( u0_u12_u5_n154 ) , .B1( u0_u12_u5_n155 ) , .ZN( u0_u12_u5_n164 ) );
  AOI21_X1 u0_u12_u5_U54 (.ZN( u0_u12_u5_n110 ) , .B1( u0_u12_u5_n122 ) , .B2( u0_u12_u5_n139 ) , .A( u0_u12_u5_n153 ) );
  INV_X1 u0_u12_u5_U55 (.A( u0_u12_u5_n153 ) , .ZN( u0_u12_u5_n176 ) );
  INV_X1 u0_u12_u5_U56 (.A( u0_u12_u5_n126 ) , .ZN( u0_u12_u5_n173 ) );
  AND2_X1 u0_u12_u5_U57 (.A2( u0_u12_u5_n104 ) , .A1( u0_u12_u5_n107 ) , .ZN( u0_u12_u5_n147 ) );
  AND2_X1 u0_u12_u5_U58 (.A2( u0_u12_u5_n104 ) , .A1( u0_u12_u5_n108 ) , .ZN( u0_u12_u5_n148 ) );
  NAND2_X1 u0_u12_u5_U59 (.A1( u0_u12_u5_n105 ) , .A2( u0_u12_u5_n106 ) , .ZN( u0_u12_u5_n158 ) );
  INV_X1 u0_u12_u5_U6 (.A( u0_u12_u5_n135 ) , .ZN( u0_u12_u5_n178 ) );
  NAND2_X1 u0_u12_u5_U60 (.A2( u0_u12_u5_n108 ) , .A1( u0_u12_u5_n109 ) , .ZN( u0_u12_u5_n139 ) );
  NAND2_X1 u0_u12_u5_U61 (.A1( u0_u12_u5_n106 ) , .A2( u0_u12_u5_n108 ) , .ZN( u0_u12_u5_n119 ) );
  NAND2_X1 u0_u12_u5_U62 (.A2( u0_u12_u5_n103 ) , .A1( u0_u12_u5_n105 ) , .ZN( u0_u12_u5_n140 ) );
  NAND2_X1 u0_u12_u5_U63 (.A2( u0_u12_u5_n104 ) , .A1( u0_u12_u5_n105 ) , .ZN( u0_u12_u5_n155 ) );
  NAND2_X1 u0_u12_u5_U64 (.A2( u0_u12_u5_n106 ) , .A1( u0_u12_u5_n107 ) , .ZN( u0_u12_u5_n122 ) );
  NAND2_X1 u0_u12_u5_U65 (.A2( u0_u12_u5_n100 ) , .A1( u0_u12_u5_n106 ) , .ZN( u0_u12_u5_n115 ) );
  NAND2_X1 u0_u12_u5_U66 (.A2( u0_u12_u5_n100 ) , .A1( u0_u12_u5_n103 ) , .ZN( u0_u12_u5_n161 ) );
  NAND2_X1 u0_u12_u5_U67 (.A1( u0_u12_u5_n105 ) , .A2( u0_u12_u5_n109 ) , .ZN( u0_u12_u5_n154 ) );
  INV_X1 u0_u12_u5_U68 (.A( u0_u12_u5_n146 ) , .ZN( u0_u12_u5_n172 ) );
  NAND2_X1 u0_u12_u5_U69 (.A1( u0_u12_u5_n103 ) , .A2( u0_u12_u5_n108 ) , .ZN( u0_u12_u5_n123 ) );
  OAI22_X1 u0_u12_u5_U7 (.B2( u0_u12_u5_n149 ) , .B1( u0_u12_u5_n150 ) , .A2( u0_u12_u5_n151 ) , .A1( u0_u12_u5_n152 ) , .ZN( u0_u12_u5_n165 ) );
  NAND2_X1 u0_u12_u5_U70 (.A2( u0_u12_u5_n103 ) , .A1( u0_u12_u5_n107 ) , .ZN( u0_u12_u5_n151 ) );
  NAND2_X1 u0_u12_u5_U71 (.A2( u0_u12_u5_n107 ) , .A1( u0_u12_u5_n109 ) , .ZN( u0_u12_u5_n120 ) );
  NAND2_X1 u0_u12_u5_U72 (.A2( u0_u12_u5_n100 ) , .A1( u0_u12_u5_n109 ) , .ZN( u0_u12_u5_n157 ) );
  AND2_X1 u0_u12_u5_U73 (.A2( u0_u12_u5_n100 ) , .A1( u0_u12_u5_n104 ) , .ZN( u0_u12_u5_n131 ) );
  INV_X1 u0_u12_u5_U74 (.A( u0_u12_u5_n102 ) , .ZN( u0_u12_u5_n195 ) );
  OAI221_X1 u0_u12_u5_U75 (.A( u0_u12_u5_n101 ) , .ZN( u0_u12_u5_n102 ) , .C2( u0_u12_u5_n115 ) , .C1( u0_u12_u5_n126 ) , .B1( u0_u12_u5_n134 ) , .B2( u0_u12_u5_n160 ) );
  OAI21_X1 u0_u12_u5_U76 (.ZN( u0_u12_u5_n101 ) , .B1( u0_u12_u5_n137 ) , .A( u0_u12_u5_n146 ) , .B2( u0_u12_u5_n147 ) );
  NOR2_X1 u0_u12_u5_U77 (.A2( u0_u12_X_34 ) , .A1( u0_u12_X_35 ) , .ZN( u0_u12_u5_n145 ) );
  NOR2_X1 u0_u12_u5_U78 (.A2( u0_u12_X_34 ) , .ZN( u0_u12_u5_n146 ) , .A1( u0_u12_u5_n171 ) );
  NOR2_X1 u0_u12_u5_U79 (.A2( u0_u12_X_31 ) , .A1( u0_u12_X_32 ) , .ZN( u0_u12_u5_n103 ) );
  NOR3_X1 u0_u12_u5_U8 (.A2( u0_u12_u5_n147 ) , .A1( u0_u12_u5_n148 ) , .ZN( u0_u12_u5_n149 ) , .A3( u0_u12_u5_n194 ) );
  NOR2_X1 u0_u12_u5_U80 (.A2( u0_u12_X_36 ) , .ZN( u0_u12_u5_n105 ) , .A1( u0_u12_u5_n180 ) );
  NOR2_X1 u0_u12_u5_U81 (.A2( u0_u12_X_33 ) , .ZN( u0_u12_u5_n108 ) , .A1( u0_u12_u5_n170 ) );
  NOR2_X1 u0_u12_u5_U82 (.A2( u0_u12_X_33 ) , .A1( u0_u12_X_36 ) , .ZN( u0_u12_u5_n107 ) );
  NOR2_X1 u0_u12_u5_U83 (.A2( u0_u12_X_31 ) , .ZN( u0_u12_u5_n104 ) , .A1( u0_u12_u5_n181 ) );
  NAND2_X1 u0_u12_u5_U84 (.A2( u0_u12_X_34 ) , .A1( u0_u12_X_35 ) , .ZN( u0_u12_u5_n153 ) );
  NAND2_X1 u0_u12_u5_U85 (.A1( u0_u12_X_34 ) , .ZN( u0_u12_u5_n126 ) , .A2( u0_u12_u5_n171 ) );
  AND2_X1 u0_u12_u5_U86 (.A1( u0_u12_X_31 ) , .A2( u0_u12_X_32 ) , .ZN( u0_u12_u5_n106 ) );
  AND2_X1 u0_u12_u5_U87 (.A1( u0_u12_X_31 ) , .ZN( u0_u12_u5_n109 ) , .A2( u0_u12_u5_n181 ) );
  INV_X1 u0_u12_u5_U88 (.A( u0_u12_X_33 ) , .ZN( u0_u12_u5_n180 ) );
  INV_X1 u0_u12_u5_U89 (.A( u0_u12_X_35 ) , .ZN( u0_u12_u5_n171 ) );
  NOR2_X1 u0_u12_u5_U9 (.ZN( u0_u12_u5_n135 ) , .A1( u0_u12_u5_n173 ) , .A2( u0_u12_u5_n176 ) );
  INV_X1 u0_u12_u5_U90 (.A( u0_u12_X_36 ) , .ZN( u0_u12_u5_n170 ) );
  INV_X1 u0_u12_u5_U91 (.A( u0_u12_X_32 ) , .ZN( u0_u12_u5_n181 ) );
  NAND4_X1 u0_u12_u5_U92 (.ZN( u0_out12_29 ) , .A4( u0_u12_u5_n129 ) , .A3( u0_u12_u5_n130 ) , .A2( u0_u12_u5_n168 ) , .A1( u0_u12_u5_n196 ) );
  AOI221_X1 u0_u12_u5_U93 (.A( u0_u12_u5_n128 ) , .ZN( u0_u12_u5_n129 ) , .C2( u0_u12_u5_n132 ) , .B2( u0_u12_u5_n159 ) , .B1( u0_u12_u5_n176 ) , .C1( u0_u12_u5_n184 ) );
  AOI222_X1 u0_u12_u5_U94 (.ZN( u0_u12_u5_n130 ) , .A2( u0_u12_u5_n146 ) , .B1( u0_u12_u5_n147 ) , .C2( u0_u12_u5_n175 ) , .B2( u0_u12_u5_n179 ) , .A1( u0_u12_u5_n188 ) , .C1( u0_u12_u5_n194 ) );
  NAND4_X1 u0_u12_u5_U95 (.ZN( u0_out12_19 ) , .A4( u0_u12_u5_n166 ) , .A3( u0_u12_u5_n167 ) , .A2( u0_u12_u5_n168 ) , .A1( u0_u12_u5_n169 ) );
  AOI22_X1 u0_u12_u5_U96 (.B2( u0_u12_u5_n145 ) , .A2( u0_u12_u5_n146 ) , .ZN( u0_u12_u5_n167 ) , .B1( u0_u12_u5_n182 ) , .A1( u0_u12_u5_n189 ) );
  NOR4_X1 u0_u12_u5_U97 (.A4( u0_u12_u5_n162 ) , .A3( u0_u12_u5_n163 ) , .A2( u0_u12_u5_n164 ) , .A1( u0_u12_u5_n165 ) , .ZN( u0_u12_u5_n166 ) );
  NAND4_X1 u0_u12_u5_U98 (.ZN( u0_out12_11 ) , .A4( u0_u12_u5_n143 ) , .A3( u0_u12_u5_n144 ) , .A2( u0_u12_u5_n169 ) , .A1( u0_u12_u5_n196 ) );
  AOI22_X1 u0_u12_u5_U99 (.A2( u0_u12_u5_n132 ) , .ZN( u0_u12_u5_n144 ) , .B2( u0_u12_u5_n145 ) , .B1( u0_u12_u5_n184 ) , .A1( u0_u12_u5_n194 ) );
  XOR2_X1 u0_u13_U19 (.B( u0_K14_37 ) , .A( u0_R12_24 ) , .Z( u0_u13_X_37 ) );
  XOR2_X1 u0_u13_U21 (.B( u0_K14_35 ) , .A( u0_R12_24 ) , .Z( u0_u13_X_35 ) );
  XOR2_X1 u0_u13_U22 (.B( u0_K14_34 ) , .A( u0_R12_23 ) , .Z( u0_u13_X_34 ) );
  XOR2_X1 u0_u13_U23 (.B( u0_K14_33 ) , .A( u0_R12_22 ) , .Z( u0_u13_X_33 ) );
  XOR2_X1 u0_u13_U25 (.B( u0_K14_31 ) , .A( u0_R12_20 ) , .Z( u0_u13_X_31 ) );
  XOR2_X1 u0_u13_U28 (.B( u0_K14_29 ) , .A( u0_R12_20 ) , .Z( u0_u13_X_29 ) );
  XOR2_X1 u0_u13_U29 (.B( u0_K14_28 ) , .A( u0_R12_19 ) , .Z( u0_u13_X_28 ) );
  XOR2_X1 u0_u13_U3 (.B( u0_K14_7 ) , .A( u0_R12_4 ) , .Z( u0_u13_X_7 ) );
  XOR2_X1 u0_u13_U31 (.B( u0_K14_26 ) , .A( u0_R12_17 ) , .Z( u0_u13_X_26 ) );
  XOR2_X1 u0_u13_U32 (.B( u0_K14_25 ) , .A( u0_R12_16 ) , .Z( u0_u13_X_25 ) );
  XOR2_X1 u0_u13_U33 (.B( u0_K14_24 ) , .A( u0_R12_17 ) , .Z( u0_u13_X_24 ) );
  XOR2_X1 u0_u13_U34 (.B( u0_K14_23 ) , .A( u0_R12_16 ) , .Z( u0_u13_X_23 ) );
  XOR2_X1 u0_u13_U5 (.B( u0_K14_5 ) , .A( u0_R12_4 ) , .Z( u0_u13_X_5 ) );
  AND3_X1 u0_u13_u0_U10 (.A2( u0_u13_u0_n112 ) , .ZN( u0_u13_u0_n127 ) , .A3( u0_u13_u0_n130 ) , .A1( u0_u13_u0_n148 ) );
  NAND2_X1 u0_u13_u0_U11 (.ZN( u0_u13_u0_n113 ) , .A1( u0_u13_u0_n139 ) , .A2( u0_u13_u0_n149 ) );
  AND2_X1 u0_u13_u0_U12 (.ZN( u0_u13_u0_n107 ) , .A1( u0_u13_u0_n130 ) , .A2( u0_u13_u0_n140 ) );
  AND2_X1 u0_u13_u0_U13 (.A2( u0_u13_u0_n129 ) , .A1( u0_u13_u0_n130 ) , .ZN( u0_u13_u0_n151 ) );
  AND2_X1 u0_u13_u0_U14 (.A1( u0_u13_u0_n108 ) , .A2( u0_u13_u0_n125 ) , .ZN( u0_u13_u0_n145 ) );
  INV_X1 u0_u13_u0_U15 (.A( u0_u13_u0_n143 ) , .ZN( u0_u13_u0_n173 ) );
  NOR2_X1 u0_u13_u0_U16 (.A2( u0_u13_u0_n136 ) , .ZN( u0_u13_u0_n147 ) , .A1( u0_u13_u0_n160 ) );
  INV_X1 u0_u13_u0_U17 (.ZN( u0_u13_u0_n172 ) , .A( u0_u13_u0_n88 ) );
  OAI222_X1 u0_u13_u0_U18 (.C1( u0_u13_u0_n108 ) , .A1( u0_u13_u0_n125 ) , .B2( u0_u13_u0_n128 ) , .B1( u0_u13_u0_n144 ) , .A2( u0_u13_u0_n158 ) , .C2( u0_u13_u0_n161 ) , .ZN( u0_u13_u0_n88 ) );
  NOR2_X1 u0_u13_u0_U19 (.A1( u0_u13_u0_n163 ) , .A2( u0_u13_u0_n164 ) , .ZN( u0_u13_u0_n95 ) );
  AOI21_X1 u0_u13_u0_U20 (.B1( u0_u13_u0_n103 ) , .ZN( u0_u13_u0_n132 ) , .A( u0_u13_u0_n165 ) , .B2( u0_u13_u0_n93 ) );
  INV_X1 u0_u13_u0_U21 (.A( u0_u13_u0_n142 ) , .ZN( u0_u13_u0_n165 ) );
  OAI221_X1 u0_u13_u0_U22 (.C1( u0_u13_u0_n121 ) , .ZN( u0_u13_u0_n122 ) , .B2( u0_u13_u0_n127 ) , .A( u0_u13_u0_n143 ) , .B1( u0_u13_u0_n144 ) , .C2( u0_u13_u0_n147 ) );
  OAI22_X1 u0_u13_u0_U23 (.B1( u0_u13_u0_n125 ) , .ZN( u0_u13_u0_n126 ) , .A1( u0_u13_u0_n138 ) , .A2( u0_u13_u0_n146 ) , .B2( u0_u13_u0_n147 ) );
  OAI22_X1 u0_u13_u0_U24 (.B1( u0_u13_u0_n131 ) , .A1( u0_u13_u0_n144 ) , .B2( u0_u13_u0_n147 ) , .A2( u0_u13_u0_n90 ) , .ZN( u0_u13_u0_n91 ) );
  AND3_X1 u0_u13_u0_U25 (.A3( u0_u13_u0_n121 ) , .A2( u0_u13_u0_n125 ) , .A1( u0_u13_u0_n148 ) , .ZN( u0_u13_u0_n90 ) );
  INV_X1 u0_u13_u0_U26 (.A( u0_u13_u0_n136 ) , .ZN( u0_u13_u0_n161 ) );
  NOR2_X1 u0_u13_u0_U27 (.A1( u0_u13_u0_n120 ) , .ZN( u0_u13_u0_n143 ) , .A2( u0_u13_u0_n167 ) );
  OAI221_X1 u0_u13_u0_U28 (.C1( u0_u13_u0_n112 ) , .ZN( u0_u13_u0_n120 ) , .B1( u0_u13_u0_n138 ) , .B2( u0_u13_u0_n141 ) , .C2( u0_u13_u0_n147 ) , .A( u0_u13_u0_n172 ) );
  AOI211_X1 u0_u13_u0_U29 (.B( u0_u13_u0_n115 ) , .A( u0_u13_u0_n116 ) , .C2( u0_u13_u0_n117 ) , .C1( u0_u13_u0_n118 ) , .ZN( u0_u13_u0_n119 ) );
  INV_X1 u0_u13_u0_U3 (.A( u0_u13_u0_n113 ) , .ZN( u0_u13_u0_n166 ) );
  AOI22_X1 u0_u13_u0_U30 (.B2( u0_u13_u0_n109 ) , .A2( u0_u13_u0_n110 ) , .ZN( u0_u13_u0_n111 ) , .B1( u0_u13_u0_n118 ) , .A1( u0_u13_u0_n160 ) );
  INV_X1 u0_u13_u0_U31 (.A( u0_u13_u0_n118 ) , .ZN( u0_u13_u0_n158 ) );
  AOI21_X1 u0_u13_u0_U32 (.ZN( u0_u13_u0_n104 ) , .B1( u0_u13_u0_n107 ) , .B2( u0_u13_u0_n141 ) , .A( u0_u13_u0_n144 ) );
  AOI21_X1 u0_u13_u0_U33 (.B1( u0_u13_u0_n127 ) , .B2( u0_u13_u0_n129 ) , .A( u0_u13_u0_n138 ) , .ZN( u0_u13_u0_n96 ) );
  AOI21_X1 u0_u13_u0_U34 (.ZN( u0_u13_u0_n116 ) , .B2( u0_u13_u0_n142 ) , .A( u0_u13_u0_n144 ) , .B1( u0_u13_u0_n166 ) );
  NAND2_X1 u0_u13_u0_U35 (.A1( u0_u13_u0_n100 ) , .A2( u0_u13_u0_n103 ) , .ZN( u0_u13_u0_n125 ) );
  NAND2_X1 u0_u13_u0_U36 (.A1( u0_u13_u0_n101 ) , .A2( u0_u13_u0_n102 ) , .ZN( u0_u13_u0_n150 ) );
  INV_X1 u0_u13_u0_U37 (.A( u0_u13_u0_n138 ) , .ZN( u0_u13_u0_n160 ) );
  NAND2_X1 u0_u13_u0_U38 (.A1( u0_u13_u0_n102 ) , .ZN( u0_u13_u0_n128 ) , .A2( u0_u13_u0_n95 ) );
  NAND2_X1 u0_u13_u0_U39 (.A1( u0_u13_u0_n100 ) , .ZN( u0_u13_u0_n129 ) , .A2( u0_u13_u0_n95 ) );
  AOI21_X1 u0_u13_u0_U4 (.B1( u0_u13_u0_n114 ) , .ZN( u0_u13_u0_n115 ) , .B2( u0_u13_u0_n129 ) , .A( u0_u13_u0_n161 ) );
  NAND2_X1 u0_u13_u0_U40 (.A2( u0_u13_u0_n100 ) , .ZN( u0_u13_u0_n131 ) , .A1( u0_u13_u0_n92 ) );
  NAND2_X1 u0_u13_u0_U41 (.A2( u0_u13_u0_n100 ) , .A1( u0_u13_u0_n101 ) , .ZN( u0_u13_u0_n139 ) );
  NAND2_X1 u0_u13_u0_U42 (.ZN( u0_u13_u0_n148 ) , .A1( u0_u13_u0_n93 ) , .A2( u0_u13_u0_n95 ) );
  NAND2_X1 u0_u13_u0_U43 (.A2( u0_u13_u0_n102 ) , .A1( u0_u13_u0_n103 ) , .ZN( u0_u13_u0_n149 ) );
  NAND2_X1 u0_u13_u0_U44 (.A2( u0_u13_u0_n102 ) , .ZN( u0_u13_u0_n114 ) , .A1( u0_u13_u0_n92 ) );
  NAND2_X1 u0_u13_u0_U45 (.A2( u0_u13_u0_n101 ) , .ZN( u0_u13_u0_n121 ) , .A1( u0_u13_u0_n93 ) );
  NAND2_X1 u0_u13_u0_U46 (.ZN( u0_u13_u0_n112 ) , .A2( u0_u13_u0_n92 ) , .A1( u0_u13_u0_n93 ) );
  OR3_X1 u0_u13_u0_U47 (.A3( u0_u13_u0_n152 ) , .A2( u0_u13_u0_n153 ) , .A1( u0_u13_u0_n154 ) , .ZN( u0_u13_u0_n155 ) );
  AOI21_X1 u0_u13_u0_U48 (.B2( u0_u13_u0_n150 ) , .B1( u0_u13_u0_n151 ) , .ZN( u0_u13_u0_n152 ) , .A( u0_u13_u0_n158 ) );
  AOI21_X1 u0_u13_u0_U49 (.A( u0_u13_u0_n144 ) , .B2( u0_u13_u0_n145 ) , .B1( u0_u13_u0_n146 ) , .ZN( u0_u13_u0_n154 ) );
  AOI21_X1 u0_u13_u0_U5 (.B2( u0_u13_u0_n131 ) , .ZN( u0_u13_u0_n134 ) , .B1( u0_u13_u0_n151 ) , .A( u0_u13_u0_n158 ) );
  AOI21_X1 u0_u13_u0_U50 (.A( u0_u13_u0_n147 ) , .B2( u0_u13_u0_n148 ) , .B1( u0_u13_u0_n149 ) , .ZN( u0_u13_u0_n153 ) );
  INV_X1 u0_u13_u0_U51 (.ZN( u0_u13_u0_n171 ) , .A( u0_u13_u0_n99 ) );
  OAI211_X1 u0_u13_u0_U52 (.C2( u0_u13_u0_n140 ) , .C1( u0_u13_u0_n161 ) , .A( u0_u13_u0_n169 ) , .B( u0_u13_u0_n98 ) , .ZN( u0_u13_u0_n99 ) );
  AOI211_X1 u0_u13_u0_U53 (.C1( u0_u13_u0_n118 ) , .A( u0_u13_u0_n123 ) , .B( u0_u13_u0_n96 ) , .C2( u0_u13_u0_n97 ) , .ZN( u0_u13_u0_n98 ) );
  INV_X1 u0_u13_u0_U54 (.ZN( u0_u13_u0_n169 ) , .A( u0_u13_u0_n91 ) );
  NOR2_X1 u0_u13_u0_U55 (.A2( u0_u13_X_6 ) , .ZN( u0_u13_u0_n100 ) , .A1( u0_u13_u0_n162 ) );
  NOR2_X1 u0_u13_u0_U56 (.A2( u0_u13_X_4 ) , .A1( u0_u13_X_5 ) , .ZN( u0_u13_u0_n118 ) );
  NOR2_X1 u0_u13_u0_U57 (.A2( u0_u13_X_2 ) , .ZN( u0_u13_u0_n103 ) , .A1( u0_u13_u0_n164 ) );
  NOR2_X1 u0_u13_u0_U58 (.A2( u0_u13_X_1 ) , .A1( u0_u13_X_2 ) , .ZN( u0_u13_u0_n92 ) );
  NOR2_X1 u0_u13_u0_U59 (.A2( u0_u13_X_1 ) , .ZN( u0_u13_u0_n101 ) , .A1( u0_u13_u0_n163 ) );
  NOR2_X1 u0_u13_u0_U6 (.A1( u0_u13_u0_n108 ) , .ZN( u0_u13_u0_n123 ) , .A2( u0_u13_u0_n158 ) );
  NAND2_X1 u0_u13_u0_U60 (.A2( u0_u13_X_4 ) , .A1( u0_u13_X_5 ) , .ZN( u0_u13_u0_n144 ) );
  NOR2_X1 u0_u13_u0_U61 (.A2( u0_u13_X_5 ) , .ZN( u0_u13_u0_n136 ) , .A1( u0_u13_u0_n159 ) );
  NAND2_X1 u0_u13_u0_U62 (.A1( u0_u13_X_5 ) , .ZN( u0_u13_u0_n138 ) , .A2( u0_u13_u0_n159 ) );
  AND2_X1 u0_u13_u0_U63 (.A2( u0_u13_X_3 ) , .A1( u0_u13_X_6 ) , .ZN( u0_u13_u0_n102 ) );
  AND2_X1 u0_u13_u0_U64 (.A1( u0_u13_X_6 ) , .A2( u0_u13_u0_n162 ) , .ZN( u0_u13_u0_n93 ) );
  INV_X1 u0_u13_u0_U65 (.A( u0_u13_X_4 ) , .ZN( u0_u13_u0_n159 ) );
  INV_X1 u0_u13_u0_U66 (.A( u0_u13_X_1 ) , .ZN( u0_u13_u0_n164 ) );
  INV_X1 u0_u13_u0_U67 (.A( u0_u13_X_2 ) , .ZN( u0_u13_u0_n163 ) );
  INV_X1 u0_u13_u0_U68 (.A( u0_u13_u0_n126 ) , .ZN( u0_u13_u0_n168 ) );
  AOI211_X1 u0_u13_u0_U69 (.B( u0_u13_u0_n133 ) , .A( u0_u13_u0_n134 ) , .C2( u0_u13_u0_n135 ) , .C1( u0_u13_u0_n136 ) , .ZN( u0_u13_u0_n137 ) );
  OAI21_X1 u0_u13_u0_U7 (.B1( u0_u13_u0_n150 ) , .B2( u0_u13_u0_n158 ) , .A( u0_u13_u0_n172 ) , .ZN( u0_u13_u0_n89 ) );
  INV_X1 u0_u13_u0_U70 (.ZN( u0_u13_u0_n174 ) , .A( u0_u13_u0_n89 ) );
  AOI211_X1 u0_u13_u0_U71 (.B( u0_u13_u0_n104 ) , .A( u0_u13_u0_n105 ) , .ZN( u0_u13_u0_n106 ) , .C2( u0_u13_u0_n113 ) , .C1( u0_u13_u0_n160 ) );
  OR4_X1 u0_u13_u0_U72 (.ZN( u0_out13_17 ) , .A4( u0_u13_u0_n122 ) , .A2( u0_u13_u0_n123 ) , .A1( u0_u13_u0_n124 ) , .A3( u0_u13_u0_n170 ) );
  AOI21_X1 u0_u13_u0_U73 (.B2( u0_u13_u0_n107 ) , .ZN( u0_u13_u0_n124 ) , .B1( u0_u13_u0_n128 ) , .A( u0_u13_u0_n161 ) );
  INV_X1 u0_u13_u0_U74 (.A( u0_u13_u0_n111 ) , .ZN( u0_u13_u0_n170 ) );
  OR4_X1 u0_u13_u0_U75 (.ZN( u0_out13_31 ) , .A4( u0_u13_u0_n155 ) , .A2( u0_u13_u0_n156 ) , .A1( u0_u13_u0_n157 ) , .A3( u0_u13_u0_n173 ) );
  AOI21_X1 u0_u13_u0_U76 (.A( u0_u13_u0_n138 ) , .B2( u0_u13_u0_n139 ) , .B1( u0_u13_u0_n140 ) , .ZN( u0_u13_u0_n157 ) );
  AOI21_X1 u0_u13_u0_U77 (.B2( u0_u13_u0_n141 ) , .B1( u0_u13_u0_n142 ) , .ZN( u0_u13_u0_n156 ) , .A( u0_u13_u0_n161 ) );
  AOI21_X1 u0_u13_u0_U78 (.B1( u0_u13_u0_n132 ) , .ZN( u0_u13_u0_n133 ) , .A( u0_u13_u0_n144 ) , .B2( u0_u13_u0_n166 ) );
  OAI22_X1 u0_u13_u0_U79 (.ZN( u0_u13_u0_n105 ) , .A2( u0_u13_u0_n132 ) , .B1( u0_u13_u0_n146 ) , .A1( u0_u13_u0_n147 ) , .B2( u0_u13_u0_n161 ) );
  AND2_X1 u0_u13_u0_U8 (.A1( u0_u13_u0_n114 ) , .A2( u0_u13_u0_n121 ) , .ZN( u0_u13_u0_n146 ) );
  NAND2_X1 u0_u13_u0_U80 (.ZN( u0_u13_u0_n110 ) , .A2( u0_u13_u0_n132 ) , .A1( u0_u13_u0_n145 ) );
  INV_X1 u0_u13_u0_U81 (.A( u0_u13_u0_n119 ) , .ZN( u0_u13_u0_n167 ) );
  NAND2_X1 u0_u13_u0_U82 (.A2( u0_u13_u0_n103 ) , .ZN( u0_u13_u0_n140 ) , .A1( u0_u13_u0_n94 ) );
  NAND2_X1 u0_u13_u0_U83 (.A1( u0_u13_u0_n101 ) , .ZN( u0_u13_u0_n130 ) , .A2( u0_u13_u0_n94 ) );
  NAND2_X1 u0_u13_u0_U84 (.ZN( u0_u13_u0_n108 ) , .A1( u0_u13_u0_n92 ) , .A2( u0_u13_u0_n94 ) );
  NAND2_X1 u0_u13_u0_U85 (.ZN( u0_u13_u0_n142 ) , .A1( u0_u13_u0_n94 ) , .A2( u0_u13_u0_n95 ) );
  INV_X1 u0_u13_u0_U86 (.A( u0_u13_X_3 ) , .ZN( u0_u13_u0_n162 ) );
  NOR2_X1 u0_u13_u0_U87 (.A2( u0_u13_X_3 ) , .A1( u0_u13_X_6 ) , .ZN( u0_u13_u0_n94 ) );
  NAND3_X1 u0_u13_u0_U88 (.ZN( u0_out13_23 ) , .A3( u0_u13_u0_n137 ) , .A1( u0_u13_u0_n168 ) , .A2( u0_u13_u0_n171 ) );
  NAND3_X1 u0_u13_u0_U89 (.A3( u0_u13_u0_n127 ) , .A2( u0_u13_u0_n128 ) , .ZN( u0_u13_u0_n135 ) , .A1( u0_u13_u0_n150 ) );
  AND2_X1 u0_u13_u0_U9 (.A1( u0_u13_u0_n131 ) , .ZN( u0_u13_u0_n141 ) , .A2( u0_u13_u0_n150 ) );
  NAND3_X1 u0_u13_u0_U90 (.ZN( u0_u13_u0_n117 ) , .A3( u0_u13_u0_n132 ) , .A2( u0_u13_u0_n139 ) , .A1( u0_u13_u0_n148 ) );
  NAND3_X1 u0_u13_u0_U91 (.ZN( u0_u13_u0_n109 ) , .A2( u0_u13_u0_n114 ) , .A3( u0_u13_u0_n140 ) , .A1( u0_u13_u0_n149 ) );
  NAND3_X1 u0_u13_u0_U92 (.ZN( u0_out13_9 ) , .A3( u0_u13_u0_n106 ) , .A2( u0_u13_u0_n171 ) , .A1( u0_u13_u0_n174 ) );
  NAND3_X1 u0_u13_u0_U93 (.A2( u0_u13_u0_n128 ) , .A1( u0_u13_u0_n132 ) , .A3( u0_u13_u0_n146 ) , .ZN( u0_u13_u0_n97 ) );
  AOI21_X1 u0_u13_u1_U10 (.B2( u0_u13_u1_n155 ) , .B1( u0_u13_u1_n156 ) , .ZN( u0_u13_u1_n157 ) , .A( u0_u13_u1_n174 ) );
  NAND3_X1 u0_u13_u1_U100 (.ZN( u0_u13_u1_n113 ) , .A1( u0_u13_u1_n120 ) , .A3( u0_u13_u1_n133 ) , .A2( u0_u13_u1_n155 ) );
  NAND2_X1 u0_u13_u1_U11 (.ZN( u0_u13_u1_n140 ) , .A2( u0_u13_u1_n150 ) , .A1( u0_u13_u1_n155 ) );
  NAND2_X1 u0_u13_u1_U12 (.A1( u0_u13_u1_n131 ) , .ZN( u0_u13_u1_n147 ) , .A2( u0_u13_u1_n153 ) );
  INV_X1 u0_u13_u1_U13 (.A( u0_u13_u1_n139 ) , .ZN( u0_u13_u1_n174 ) );
  OR4_X1 u0_u13_u1_U14 (.A4( u0_u13_u1_n106 ) , .A3( u0_u13_u1_n107 ) , .ZN( u0_u13_u1_n108 ) , .A1( u0_u13_u1_n117 ) , .A2( u0_u13_u1_n184 ) );
  AOI21_X1 u0_u13_u1_U15 (.ZN( u0_u13_u1_n106 ) , .A( u0_u13_u1_n112 ) , .B1( u0_u13_u1_n154 ) , .B2( u0_u13_u1_n156 ) );
  AOI21_X1 u0_u13_u1_U16 (.ZN( u0_u13_u1_n107 ) , .B1( u0_u13_u1_n134 ) , .B2( u0_u13_u1_n149 ) , .A( u0_u13_u1_n174 ) );
  INV_X1 u0_u13_u1_U17 (.A( u0_u13_u1_n101 ) , .ZN( u0_u13_u1_n184 ) );
  INV_X1 u0_u13_u1_U18 (.A( u0_u13_u1_n112 ) , .ZN( u0_u13_u1_n171 ) );
  NAND2_X1 u0_u13_u1_U19 (.ZN( u0_u13_u1_n141 ) , .A1( u0_u13_u1_n153 ) , .A2( u0_u13_u1_n156 ) );
  AND2_X1 u0_u13_u1_U20 (.A1( u0_u13_u1_n123 ) , .ZN( u0_u13_u1_n134 ) , .A2( u0_u13_u1_n161 ) );
  NAND2_X1 u0_u13_u1_U21 (.A2( u0_u13_u1_n115 ) , .A1( u0_u13_u1_n116 ) , .ZN( u0_u13_u1_n148 ) );
  NAND2_X1 u0_u13_u1_U22 (.A2( u0_u13_u1_n133 ) , .A1( u0_u13_u1_n135 ) , .ZN( u0_u13_u1_n159 ) );
  NAND2_X1 u0_u13_u1_U23 (.A2( u0_u13_u1_n115 ) , .A1( u0_u13_u1_n120 ) , .ZN( u0_u13_u1_n132 ) );
  INV_X1 u0_u13_u1_U24 (.A( u0_u13_u1_n154 ) , .ZN( u0_u13_u1_n178 ) );
  AOI22_X1 u0_u13_u1_U25 (.B2( u0_u13_u1_n113 ) , .A2( u0_u13_u1_n114 ) , .ZN( u0_u13_u1_n125 ) , .A1( u0_u13_u1_n171 ) , .B1( u0_u13_u1_n173 ) );
  NAND2_X1 u0_u13_u1_U26 (.ZN( u0_u13_u1_n114 ) , .A1( u0_u13_u1_n134 ) , .A2( u0_u13_u1_n156 ) );
  INV_X1 u0_u13_u1_U27 (.A( u0_u13_u1_n151 ) , .ZN( u0_u13_u1_n183 ) );
  AND2_X1 u0_u13_u1_U28 (.A1( u0_u13_u1_n129 ) , .A2( u0_u13_u1_n133 ) , .ZN( u0_u13_u1_n149 ) );
  INV_X1 u0_u13_u1_U29 (.A( u0_u13_u1_n131 ) , .ZN( u0_u13_u1_n180 ) );
  INV_X1 u0_u13_u1_U3 (.A( u0_u13_u1_n159 ) , .ZN( u0_u13_u1_n182 ) );
  OAI221_X1 u0_u13_u1_U30 (.A( u0_u13_u1_n119 ) , .C2( u0_u13_u1_n129 ) , .ZN( u0_u13_u1_n138 ) , .B2( u0_u13_u1_n152 ) , .C1( u0_u13_u1_n174 ) , .B1( u0_u13_u1_n187 ) );
  INV_X1 u0_u13_u1_U31 (.A( u0_u13_u1_n148 ) , .ZN( u0_u13_u1_n187 ) );
  AOI211_X1 u0_u13_u1_U32 (.B( u0_u13_u1_n117 ) , .A( u0_u13_u1_n118 ) , .ZN( u0_u13_u1_n119 ) , .C2( u0_u13_u1_n146 ) , .C1( u0_u13_u1_n159 ) );
  NOR2_X1 u0_u13_u1_U33 (.A1( u0_u13_u1_n168 ) , .A2( u0_u13_u1_n176 ) , .ZN( u0_u13_u1_n98 ) );
  AOI211_X1 u0_u13_u1_U34 (.B( u0_u13_u1_n162 ) , .A( u0_u13_u1_n163 ) , .C2( u0_u13_u1_n164 ) , .ZN( u0_u13_u1_n165 ) , .C1( u0_u13_u1_n171 ) );
  AOI21_X1 u0_u13_u1_U35 (.A( u0_u13_u1_n160 ) , .B2( u0_u13_u1_n161 ) , .ZN( u0_u13_u1_n162 ) , .B1( u0_u13_u1_n182 ) );
  OR2_X1 u0_u13_u1_U36 (.A2( u0_u13_u1_n157 ) , .A1( u0_u13_u1_n158 ) , .ZN( u0_u13_u1_n163 ) );
  OAI21_X1 u0_u13_u1_U37 (.B2( u0_u13_u1_n123 ) , .ZN( u0_u13_u1_n145 ) , .B1( u0_u13_u1_n160 ) , .A( u0_u13_u1_n185 ) );
  INV_X1 u0_u13_u1_U38 (.A( u0_u13_u1_n122 ) , .ZN( u0_u13_u1_n185 ) );
  AOI21_X1 u0_u13_u1_U39 (.B2( u0_u13_u1_n120 ) , .B1( u0_u13_u1_n121 ) , .ZN( u0_u13_u1_n122 ) , .A( u0_u13_u1_n128 ) );
  AOI221_X1 u0_u13_u1_U4 (.A( u0_u13_u1_n138 ) , .C2( u0_u13_u1_n139 ) , .C1( u0_u13_u1_n140 ) , .B2( u0_u13_u1_n141 ) , .ZN( u0_u13_u1_n142 ) , .B1( u0_u13_u1_n175 ) );
  NAND2_X1 u0_u13_u1_U40 (.A1( u0_u13_u1_n128 ) , .ZN( u0_u13_u1_n146 ) , .A2( u0_u13_u1_n160 ) );
  NAND2_X1 u0_u13_u1_U41 (.A2( u0_u13_u1_n112 ) , .ZN( u0_u13_u1_n139 ) , .A1( u0_u13_u1_n152 ) );
  NAND2_X1 u0_u13_u1_U42 (.A1( u0_u13_u1_n105 ) , .ZN( u0_u13_u1_n156 ) , .A2( u0_u13_u1_n99 ) );
  AOI221_X1 u0_u13_u1_U43 (.B1( u0_u13_u1_n140 ) , .ZN( u0_u13_u1_n167 ) , .B2( u0_u13_u1_n172 ) , .C2( u0_u13_u1_n175 ) , .C1( u0_u13_u1_n178 ) , .A( u0_u13_u1_n188 ) );
  INV_X1 u0_u13_u1_U44 (.ZN( u0_u13_u1_n188 ) , .A( u0_u13_u1_n97 ) );
  AOI211_X1 u0_u13_u1_U45 (.A( u0_u13_u1_n118 ) , .C1( u0_u13_u1_n132 ) , .C2( u0_u13_u1_n139 ) , .B( u0_u13_u1_n96 ) , .ZN( u0_u13_u1_n97 ) );
  AOI21_X1 u0_u13_u1_U46 (.B2( u0_u13_u1_n121 ) , .B1( u0_u13_u1_n135 ) , .A( u0_u13_u1_n152 ) , .ZN( u0_u13_u1_n96 ) );
  NOR2_X1 u0_u13_u1_U47 (.ZN( u0_u13_u1_n117 ) , .A1( u0_u13_u1_n121 ) , .A2( u0_u13_u1_n160 ) );
  AOI21_X1 u0_u13_u1_U48 (.A( u0_u13_u1_n128 ) , .B2( u0_u13_u1_n129 ) , .ZN( u0_u13_u1_n130 ) , .B1( u0_u13_u1_n150 ) );
  NAND2_X1 u0_u13_u1_U49 (.ZN( u0_u13_u1_n112 ) , .A1( u0_u13_u1_n169 ) , .A2( u0_u13_u1_n170 ) );
  AOI211_X1 u0_u13_u1_U5 (.ZN( u0_u13_u1_n124 ) , .A( u0_u13_u1_n138 ) , .C2( u0_u13_u1_n139 ) , .B( u0_u13_u1_n145 ) , .C1( u0_u13_u1_n147 ) );
  NAND2_X1 u0_u13_u1_U50 (.ZN( u0_u13_u1_n129 ) , .A2( u0_u13_u1_n95 ) , .A1( u0_u13_u1_n98 ) );
  NAND2_X1 u0_u13_u1_U51 (.A1( u0_u13_u1_n102 ) , .ZN( u0_u13_u1_n154 ) , .A2( u0_u13_u1_n99 ) );
  NAND2_X1 u0_u13_u1_U52 (.A2( u0_u13_u1_n100 ) , .ZN( u0_u13_u1_n135 ) , .A1( u0_u13_u1_n99 ) );
  AOI21_X1 u0_u13_u1_U53 (.A( u0_u13_u1_n152 ) , .B2( u0_u13_u1_n153 ) , .B1( u0_u13_u1_n154 ) , .ZN( u0_u13_u1_n158 ) );
  INV_X1 u0_u13_u1_U54 (.A( u0_u13_u1_n160 ) , .ZN( u0_u13_u1_n175 ) );
  NAND2_X1 u0_u13_u1_U55 (.A1( u0_u13_u1_n100 ) , .ZN( u0_u13_u1_n116 ) , .A2( u0_u13_u1_n95 ) );
  NAND2_X1 u0_u13_u1_U56 (.A1( u0_u13_u1_n102 ) , .ZN( u0_u13_u1_n131 ) , .A2( u0_u13_u1_n95 ) );
  NAND2_X1 u0_u13_u1_U57 (.A2( u0_u13_u1_n104 ) , .ZN( u0_u13_u1_n121 ) , .A1( u0_u13_u1_n98 ) );
  NAND2_X1 u0_u13_u1_U58 (.A1( u0_u13_u1_n103 ) , .ZN( u0_u13_u1_n153 ) , .A2( u0_u13_u1_n98 ) );
  NAND2_X1 u0_u13_u1_U59 (.A2( u0_u13_u1_n104 ) , .A1( u0_u13_u1_n105 ) , .ZN( u0_u13_u1_n133 ) );
  AOI22_X1 u0_u13_u1_U6 (.B2( u0_u13_u1_n136 ) , .A2( u0_u13_u1_n137 ) , .ZN( u0_u13_u1_n143 ) , .A1( u0_u13_u1_n171 ) , .B1( u0_u13_u1_n173 ) );
  NAND2_X1 u0_u13_u1_U60 (.ZN( u0_u13_u1_n150 ) , .A2( u0_u13_u1_n98 ) , .A1( u0_u13_u1_n99 ) );
  NAND2_X1 u0_u13_u1_U61 (.A1( u0_u13_u1_n105 ) , .ZN( u0_u13_u1_n155 ) , .A2( u0_u13_u1_n95 ) );
  OAI21_X1 u0_u13_u1_U62 (.ZN( u0_u13_u1_n109 ) , .B1( u0_u13_u1_n129 ) , .B2( u0_u13_u1_n160 ) , .A( u0_u13_u1_n167 ) );
  NAND2_X1 u0_u13_u1_U63 (.A2( u0_u13_u1_n100 ) , .A1( u0_u13_u1_n103 ) , .ZN( u0_u13_u1_n120 ) );
  NAND2_X1 u0_u13_u1_U64 (.A1( u0_u13_u1_n102 ) , .A2( u0_u13_u1_n104 ) , .ZN( u0_u13_u1_n115 ) );
  NAND2_X1 u0_u13_u1_U65 (.A2( u0_u13_u1_n100 ) , .A1( u0_u13_u1_n104 ) , .ZN( u0_u13_u1_n151 ) );
  NAND2_X1 u0_u13_u1_U66 (.A2( u0_u13_u1_n103 ) , .A1( u0_u13_u1_n105 ) , .ZN( u0_u13_u1_n161 ) );
  INV_X1 u0_u13_u1_U67 (.A( u0_u13_u1_n152 ) , .ZN( u0_u13_u1_n173 ) );
  INV_X1 u0_u13_u1_U68 (.A( u0_u13_u1_n128 ) , .ZN( u0_u13_u1_n172 ) );
  NAND2_X1 u0_u13_u1_U69 (.A2( u0_u13_u1_n102 ) , .A1( u0_u13_u1_n103 ) , .ZN( u0_u13_u1_n123 ) );
  INV_X1 u0_u13_u1_U7 (.A( u0_u13_u1_n147 ) , .ZN( u0_u13_u1_n181 ) );
  NOR2_X1 u0_u13_u1_U70 (.A2( u0_u13_X_7 ) , .A1( u0_u13_X_8 ) , .ZN( u0_u13_u1_n95 ) );
  NOR2_X1 u0_u13_u1_U71 (.A1( u0_u13_X_12 ) , .A2( u0_u13_X_9 ) , .ZN( u0_u13_u1_n100 ) );
  NOR2_X1 u0_u13_u1_U72 (.A2( u0_u13_X_8 ) , .A1( u0_u13_u1_n177 ) , .ZN( u0_u13_u1_n99 ) );
  NOR2_X1 u0_u13_u1_U73 (.A2( u0_u13_X_12 ) , .ZN( u0_u13_u1_n102 ) , .A1( u0_u13_u1_n176 ) );
  NOR2_X1 u0_u13_u1_U74 (.A2( u0_u13_X_9 ) , .ZN( u0_u13_u1_n105 ) , .A1( u0_u13_u1_n168 ) );
  NAND2_X1 u0_u13_u1_U75 (.A1( u0_u13_X_10 ) , .ZN( u0_u13_u1_n160 ) , .A2( u0_u13_u1_n169 ) );
  NAND2_X1 u0_u13_u1_U76 (.A2( u0_u13_X_10 ) , .A1( u0_u13_X_11 ) , .ZN( u0_u13_u1_n152 ) );
  NAND2_X1 u0_u13_u1_U77 (.A1( u0_u13_X_11 ) , .ZN( u0_u13_u1_n128 ) , .A2( u0_u13_u1_n170 ) );
  AND2_X1 u0_u13_u1_U78 (.A2( u0_u13_X_7 ) , .A1( u0_u13_X_8 ) , .ZN( u0_u13_u1_n104 ) );
  AND2_X1 u0_u13_u1_U79 (.A1( u0_u13_X_8 ) , .ZN( u0_u13_u1_n103 ) , .A2( u0_u13_u1_n177 ) );
  NOR2_X1 u0_u13_u1_U8 (.A1( u0_u13_u1_n112 ) , .A2( u0_u13_u1_n116 ) , .ZN( u0_u13_u1_n118 ) );
  INV_X1 u0_u13_u1_U80 (.A( u0_u13_X_10 ) , .ZN( u0_u13_u1_n170 ) );
  INV_X1 u0_u13_u1_U81 (.A( u0_u13_X_9 ) , .ZN( u0_u13_u1_n176 ) );
  INV_X1 u0_u13_u1_U82 (.A( u0_u13_X_11 ) , .ZN( u0_u13_u1_n169 ) );
  INV_X1 u0_u13_u1_U83 (.A( u0_u13_X_12 ) , .ZN( u0_u13_u1_n168 ) );
  INV_X1 u0_u13_u1_U84 (.A( u0_u13_X_7 ) , .ZN( u0_u13_u1_n177 ) );
  NAND4_X1 u0_u13_u1_U85 (.ZN( u0_out13_28 ) , .A4( u0_u13_u1_n124 ) , .A3( u0_u13_u1_n125 ) , .A2( u0_u13_u1_n126 ) , .A1( u0_u13_u1_n127 ) );
  OAI21_X1 u0_u13_u1_U86 (.ZN( u0_u13_u1_n127 ) , .B2( u0_u13_u1_n139 ) , .B1( u0_u13_u1_n175 ) , .A( u0_u13_u1_n183 ) );
  OAI21_X1 u0_u13_u1_U87 (.ZN( u0_u13_u1_n126 ) , .B2( u0_u13_u1_n140 ) , .A( u0_u13_u1_n146 ) , .B1( u0_u13_u1_n178 ) );
  NAND4_X1 u0_u13_u1_U88 (.ZN( u0_out13_18 ) , .A4( u0_u13_u1_n165 ) , .A3( u0_u13_u1_n166 ) , .A1( u0_u13_u1_n167 ) , .A2( u0_u13_u1_n186 ) );
  AOI22_X1 u0_u13_u1_U89 (.B2( u0_u13_u1_n146 ) , .B1( u0_u13_u1_n147 ) , .A2( u0_u13_u1_n148 ) , .ZN( u0_u13_u1_n166 ) , .A1( u0_u13_u1_n172 ) );
  OAI21_X1 u0_u13_u1_U9 (.ZN( u0_u13_u1_n101 ) , .B1( u0_u13_u1_n141 ) , .A( u0_u13_u1_n146 ) , .B2( u0_u13_u1_n183 ) );
  INV_X1 u0_u13_u1_U90 (.A( u0_u13_u1_n145 ) , .ZN( u0_u13_u1_n186 ) );
  NAND4_X1 u0_u13_u1_U91 (.ZN( u0_out13_2 ) , .A4( u0_u13_u1_n142 ) , .A3( u0_u13_u1_n143 ) , .A2( u0_u13_u1_n144 ) , .A1( u0_u13_u1_n179 ) );
  OAI21_X1 u0_u13_u1_U92 (.B2( u0_u13_u1_n132 ) , .ZN( u0_u13_u1_n144 ) , .A( u0_u13_u1_n146 ) , .B1( u0_u13_u1_n180 ) );
  INV_X1 u0_u13_u1_U93 (.A( u0_u13_u1_n130 ) , .ZN( u0_u13_u1_n179 ) );
  OR4_X1 u0_u13_u1_U94 (.ZN( u0_out13_13 ) , .A4( u0_u13_u1_n108 ) , .A3( u0_u13_u1_n109 ) , .A2( u0_u13_u1_n110 ) , .A1( u0_u13_u1_n111 ) );
  AOI21_X1 u0_u13_u1_U95 (.ZN( u0_u13_u1_n111 ) , .A( u0_u13_u1_n128 ) , .B2( u0_u13_u1_n131 ) , .B1( u0_u13_u1_n135 ) );
  AOI21_X1 u0_u13_u1_U96 (.ZN( u0_u13_u1_n110 ) , .A( u0_u13_u1_n116 ) , .B1( u0_u13_u1_n152 ) , .B2( u0_u13_u1_n160 ) );
  NAND3_X1 u0_u13_u1_U97 (.A3( u0_u13_u1_n149 ) , .A2( u0_u13_u1_n150 ) , .A1( u0_u13_u1_n151 ) , .ZN( u0_u13_u1_n164 ) );
  NAND3_X1 u0_u13_u1_U98 (.A3( u0_u13_u1_n134 ) , .A2( u0_u13_u1_n135 ) , .ZN( u0_u13_u1_n136 ) , .A1( u0_u13_u1_n151 ) );
  NAND3_X1 u0_u13_u1_U99 (.A1( u0_u13_u1_n133 ) , .ZN( u0_u13_u1_n137 ) , .A2( u0_u13_u1_n154 ) , .A3( u0_u13_u1_n181 ) );
  OAI22_X1 u0_u13_u3_U10 (.B1( u0_u13_u3_n113 ) , .A2( u0_u13_u3_n135 ) , .A1( u0_u13_u3_n150 ) , .B2( u0_u13_u3_n164 ) , .ZN( u0_u13_u3_n98 ) );
  OAI211_X1 u0_u13_u3_U11 (.B( u0_u13_u3_n106 ) , .ZN( u0_u13_u3_n119 ) , .C2( u0_u13_u3_n128 ) , .C1( u0_u13_u3_n167 ) , .A( u0_u13_u3_n181 ) );
  AOI221_X1 u0_u13_u3_U12 (.C1( u0_u13_u3_n105 ) , .ZN( u0_u13_u3_n106 ) , .A( u0_u13_u3_n131 ) , .B2( u0_u13_u3_n132 ) , .C2( u0_u13_u3_n133 ) , .B1( u0_u13_u3_n169 ) );
  INV_X1 u0_u13_u3_U13 (.ZN( u0_u13_u3_n181 ) , .A( u0_u13_u3_n98 ) );
  NAND2_X1 u0_u13_u3_U14 (.ZN( u0_u13_u3_n105 ) , .A2( u0_u13_u3_n130 ) , .A1( u0_u13_u3_n155 ) );
  AOI22_X1 u0_u13_u3_U15 (.B1( u0_u13_u3_n115 ) , .A2( u0_u13_u3_n116 ) , .ZN( u0_u13_u3_n123 ) , .B2( u0_u13_u3_n133 ) , .A1( u0_u13_u3_n169 ) );
  NAND2_X1 u0_u13_u3_U16 (.ZN( u0_u13_u3_n116 ) , .A2( u0_u13_u3_n151 ) , .A1( u0_u13_u3_n182 ) );
  NOR2_X1 u0_u13_u3_U17 (.ZN( u0_u13_u3_n126 ) , .A2( u0_u13_u3_n150 ) , .A1( u0_u13_u3_n164 ) );
  AOI21_X1 u0_u13_u3_U18 (.ZN( u0_u13_u3_n112 ) , .B2( u0_u13_u3_n146 ) , .B1( u0_u13_u3_n155 ) , .A( u0_u13_u3_n167 ) );
  NAND2_X1 u0_u13_u3_U19 (.A1( u0_u13_u3_n135 ) , .ZN( u0_u13_u3_n142 ) , .A2( u0_u13_u3_n164 ) );
  NAND2_X1 u0_u13_u3_U20 (.ZN( u0_u13_u3_n132 ) , .A2( u0_u13_u3_n152 ) , .A1( u0_u13_u3_n156 ) );
  AND2_X1 u0_u13_u3_U21 (.A2( u0_u13_u3_n113 ) , .A1( u0_u13_u3_n114 ) , .ZN( u0_u13_u3_n151 ) );
  INV_X1 u0_u13_u3_U22 (.A( u0_u13_u3_n133 ) , .ZN( u0_u13_u3_n165 ) );
  INV_X1 u0_u13_u3_U23 (.A( u0_u13_u3_n135 ) , .ZN( u0_u13_u3_n170 ) );
  NAND2_X1 u0_u13_u3_U24 (.A1( u0_u13_u3_n107 ) , .A2( u0_u13_u3_n108 ) , .ZN( u0_u13_u3_n140 ) );
  NAND2_X1 u0_u13_u3_U25 (.ZN( u0_u13_u3_n117 ) , .A1( u0_u13_u3_n124 ) , .A2( u0_u13_u3_n148 ) );
  NAND2_X1 u0_u13_u3_U26 (.ZN( u0_u13_u3_n143 ) , .A1( u0_u13_u3_n165 ) , .A2( u0_u13_u3_n167 ) );
  INV_X1 u0_u13_u3_U27 (.A( u0_u13_u3_n130 ) , .ZN( u0_u13_u3_n177 ) );
  INV_X1 u0_u13_u3_U28 (.A( u0_u13_u3_n128 ) , .ZN( u0_u13_u3_n176 ) );
  INV_X1 u0_u13_u3_U29 (.A( u0_u13_u3_n155 ) , .ZN( u0_u13_u3_n174 ) );
  INV_X1 u0_u13_u3_U3 (.A( u0_u13_u3_n129 ) , .ZN( u0_u13_u3_n183 ) );
  INV_X1 u0_u13_u3_U30 (.A( u0_u13_u3_n139 ) , .ZN( u0_u13_u3_n185 ) );
  NOR2_X1 u0_u13_u3_U31 (.ZN( u0_u13_u3_n135 ) , .A2( u0_u13_u3_n141 ) , .A1( u0_u13_u3_n169 ) );
  OAI222_X1 u0_u13_u3_U32 (.C2( u0_u13_u3_n107 ) , .A2( u0_u13_u3_n108 ) , .B1( u0_u13_u3_n135 ) , .ZN( u0_u13_u3_n138 ) , .B2( u0_u13_u3_n146 ) , .C1( u0_u13_u3_n154 ) , .A1( u0_u13_u3_n164 ) );
  NOR4_X1 u0_u13_u3_U33 (.A4( u0_u13_u3_n157 ) , .A3( u0_u13_u3_n158 ) , .A2( u0_u13_u3_n159 ) , .A1( u0_u13_u3_n160 ) , .ZN( u0_u13_u3_n161 ) );
  AOI21_X1 u0_u13_u3_U34 (.B2( u0_u13_u3_n152 ) , .B1( u0_u13_u3_n153 ) , .ZN( u0_u13_u3_n158 ) , .A( u0_u13_u3_n164 ) );
  AOI21_X1 u0_u13_u3_U35 (.A( u0_u13_u3_n154 ) , .B2( u0_u13_u3_n155 ) , .B1( u0_u13_u3_n156 ) , .ZN( u0_u13_u3_n157 ) );
  AOI21_X1 u0_u13_u3_U36 (.A( u0_u13_u3_n149 ) , .B2( u0_u13_u3_n150 ) , .B1( u0_u13_u3_n151 ) , .ZN( u0_u13_u3_n159 ) );
  AOI211_X1 u0_u13_u3_U37 (.ZN( u0_u13_u3_n109 ) , .A( u0_u13_u3_n119 ) , .C2( u0_u13_u3_n129 ) , .B( u0_u13_u3_n138 ) , .C1( u0_u13_u3_n141 ) );
  AOI211_X1 u0_u13_u3_U38 (.B( u0_u13_u3_n119 ) , .A( u0_u13_u3_n120 ) , .C2( u0_u13_u3_n121 ) , .ZN( u0_u13_u3_n122 ) , .C1( u0_u13_u3_n179 ) );
  INV_X1 u0_u13_u3_U39 (.A( u0_u13_u3_n156 ) , .ZN( u0_u13_u3_n179 ) );
  INV_X1 u0_u13_u3_U4 (.A( u0_u13_u3_n140 ) , .ZN( u0_u13_u3_n182 ) );
  OAI22_X1 u0_u13_u3_U40 (.B1( u0_u13_u3_n118 ) , .ZN( u0_u13_u3_n120 ) , .A1( u0_u13_u3_n135 ) , .B2( u0_u13_u3_n154 ) , .A2( u0_u13_u3_n178 ) );
  AND3_X1 u0_u13_u3_U41 (.ZN( u0_u13_u3_n118 ) , .A2( u0_u13_u3_n124 ) , .A1( u0_u13_u3_n144 ) , .A3( u0_u13_u3_n152 ) );
  INV_X1 u0_u13_u3_U42 (.A( u0_u13_u3_n121 ) , .ZN( u0_u13_u3_n164 ) );
  NAND2_X1 u0_u13_u3_U43 (.ZN( u0_u13_u3_n133 ) , .A1( u0_u13_u3_n154 ) , .A2( u0_u13_u3_n164 ) );
  OAI211_X1 u0_u13_u3_U44 (.B( u0_u13_u3_n127 ) , .ZN( u0_u13_u3_n139 ) , .C1( u0_u13_u3_n150 ) , .C2( u0_u13_u3_n154 ) , .A( u0_u13_u3_n184 ) );
  INV_X1 u0_u13_u3_U45 (.A( u0_u13_u3_n125 ) , .ZN( u0_u13_u3_n184 ) );
  AOI221_X1 u0_u13_u3_U46 (.A( u0_u13_u3_n126 ) , .ZN( u0_u13_u3_n127 ) , .C2( u0_u13_u3_n132 ) , .C1( u0_u13_u3_n169 ) , .B2( u0_u13_u3_n170 ) , .B1( u0_u13_u3_n174 ) );
  OAI22_X1 u0_u13_u3_U47 (.A1( u0_u13_u3_n124 ) , .ZN( u0_u13_u3_n125 ) , .B2( u0_u13_u3_n145 ) , .A2( u0_u13_u3_n165 ) , .B1( u0_u13_u3_n167 ) );
  NOR2_X1 u0_u13_u3_U48 (.A1( u0_u13_u3_n113 ) , .ZN( u0_u13_u3_n131 ) , .A2( u0_u13_u3_n154 ) );
  NAND2_X1 u0_u13_u3_U49 (.A1( u0_u13_u3_n103 ) , .ZN( u0_u13_u3_n150 ) , .A2( u0_u13_u3_n99 ) );
  INV_X1 u0_u13_u3_U5 (.A( u0_u13_u3_n117 ) , .ZN( u0_u13_u3_n178 ) );
  NAND2_X1 u0_u13_u3_U50 (.A2( u0_u13_u3_n102 ) , .ZN( u0_u13_u3_n155 ) , .A1( u0_u13_u3_n97 ) );
  INV_X1 u0_u13_u3_U51 (.A( u0_u13_u3_n141 ) , .ZN( u0_u13_u3_n167 ) );
  AOI21_X1 u0_u13_u3_U52 (.B2( u0_u13_u3_n114 ) , .B1( u0_u13_u3_n146 ) , .A( u0_u13_u3_n154 ) , .ZN( u0_u13_u3_n94 ) );
  AOI21_X1 u0_u13_u3_U53 (.ZN( u0_u13_u3_n110 ) , .B2( u0_u13_u3_n142 ) , .B1( u0_u13_u3_n186 ) , .A( u0_u13_u3_n95 ) );
  INV_X1 u0_u13_u3_U54 (.A( u0_u13_u3_n145 ) , .ZN( u0_u13_u3_n186 ) );
  AOI21_X1 u0_u13_u3_U55 (.B1( u0_u13_u3_n124 ) , .A( u0_u13_u3_n149 ) , .B2( u0_u13_u3_n155 ) , .ZN( u0_u13_u3_n95 ) );
  INV_X1 u0_u13_u3_U56 (.A( u0_u13_u3_n149 ) , .ZN( u0_u13_u3_n169 ) );
  NAND2_X1 u0_u13_u3_U57 (.ZN( u0_u13_u3_n124 ) , .A1( u0_u13_u3_n96 ) , .A2( u0_u13_u3_n97 ) );
  NAND2_X1 u0_u13_u3_U58 (.A2( u0_u13_u3_n100 ) , .ZN( u0_u13_u3_n146 ) , .A1( u0_u13_u3_n96 ) );
  NAND2_X1 u0_u13_u3_U59 (.A1( u0_u13_u3_n101 ) , .ZN( u0_u13_u3_n145 ) , .A2( u0_u13_u3_n99 ) );
  AOI221_X1 u0_u13_u3_U6 (.A( u0_u13_u3_n131 ) , .C2( u0_u13_u3_n132 ) , .C1( u0_u13_u3_n133 ) , .ZN( u0_u13_u3_n134 ) , .B1( u0_u13_u3_n143 ) , .B2( u0_u13_u3_n177 ) );
  NAND2_X1 u0_u13_u3_U60 (.A1( u0_u13_u3_n100 ) , .ZN( u0_u13_u3_n156 ) , .A2( u0_u13_u3_n99 ) );
  NAND2_X1 u0_u13_u3_U61 (.A2( u0_u13_u3_n101 ) , .A1( u0_u13_u3_n104 ) , .ZN( u0_u13_u3_n148 ) );
  NAND2_X1 u0_u13_u3_U62 (.A1( u0_u13_u3_n100 ) , .A2( u0_u13_u3_n102 ) , .ZN( u0_u13_u3_n128 ) );
  NAND2_X1 u0_u13_u3_U63 (.A2( u0_u13_u3_n101 ) , .A1( u0_u13_u3_n102 ) , .ZN( u0_u13_u3_n152 ) );
  NAND2_X1 u0_u13_u3_U64 (.A2( u0_u13_u3_n101 ) , .ZN( u0_u13_u3_n114 ) , .A1( u0_u13_u3_n96 ) );
  NAND2_X1 u0_u13_u3_U65 (.ZN( u0_u13_u3_n107 ) , .A1( u0_u13_u3_n97 ) , .A2( u0_u13_u3_n99 ) );
  NAND2_X1 u0_u13_u3_U66 (.A2( u0_u13_u3_n100 ) , .A1( u0_u13_u3_n104 ) , .ZN( u0_u13_u3_n113 ) );
  NAND2_X1 u0_u13_u3_U67 (.A1( u0_u13_u3_n104 ) , .ZN( u0_u13_u3_n153 ) , .A2( u0_u13_u3_n97 ) );
  NAND2_X1 u0_u13_u3_U68 (.A2( u0_u13_u3_n103 ) , .A1( u0_u13_u3_n104 ) , .ZN( u0_u13_u3_n130 ) );
  NAND2_X1 u0_u13_u3_U69 (.A2( u0_u13_u3_n103 ) , .ZN( u0_u13_u3_n144 ) , .A1( u0_u13_u3_n96 ) );
  OAI22_X1 u0_u13_u3_U7 (.B2( u0_u13_u3_n147 ) , .A2( u0_u13_u3_n148 ) , .ZN( u0_u13_u3_n160 ) , .B1( u0_u13_u3_n165 ) , .A1( u0_u13_u3_n168 ) );
  NAND2_X1 u0_u13_u3_U70 (.A1( u0_u13_u3_n102 ) , .A2( u0_u13_u3_n103 ) , .ZN( u0_u13_u3_n108 ) );
  NOR2_X1 u0_u13_u3_U71 (.A2( u0_u13_X_19 ) , .A1( u0_u13_X_20 ) , .ZN( u0_u13_u3_n99 ) );
  NOR2_X1 u0_u13_u3_U72 (.A2( u0_u13_X_21 ) , .A1( u0_u13_X_24 ) , .ZN( u0_u13_u3_n103 ) );
  NOR2_X1 u0_u13_u3_U73 (.A2( u0_u13_X_24 ) , .A1( u0_u13_u3_n171 ) , .ZN( u0_u13_u3_n97 ) );
  NOR2_X1 u0_u13_u3_U74 (.A2( u0_u13_X_23 ) , .ZN( u0_u13_u3_n141 ) , .A1( u0_u13_u3_n166 ) );
  NOR2_X1 u0_u13_u3_U75 (.A2( u0_u13_X_19 ) , .A1( u0_u13_u3_n172 ) , .ZN( u0_u13_u3_n96 ) );
  NAND2_X1 u0_u13_u3_U76 (.A1( u0_u13_X_22 ) , .A2( u0_u13_X_23 ) , .ZN( u0_u13_u3_n154 ) );
  NAND2_X1 u0_u13_u3_U77 (.A1( u0_u13_X_23 ) , .ZN( u0_u13_u3_n149 ) , .A2( u0_u13_u3_n166 ) );
  NOR2_X1 u0_u13_u3_U78 (.A2( u0_u13_X_22 ) , .A1( u0_u13_X_23 ) , .ZN( u0_u13_u3_n121 ) );
  AND2_X1 u0_u13_u3_U79 (.A1( u0_u13_X_24 ) , .ZN( u0_u13_u3_n101 ) , .A2( u0_u13_u3_n171 ) );
  AND3_X1 u0_u13_u3_U8 (.A3( u0_u13_u3_n144 ) , .A2( u0_u13_u3_n145 ) , .A1( u0_u13_u3_n146 ) , .ZN( u0_u13_u3_n147 ) );
  AND2_X1 u0_u13_u3_U80 (.A1( u0_u13_X_19 ) , .ZN( u0_u13_u3_n102 ) , .A2( u0_u13_u3_n172 ) );
  AND2_X1 u0_u13_u3_U81 (.A1( u0_u13_X_21 ) , .A2( u0_u13_X_24 ) , .ZN( u0_u13_u3_n100 ) );
  AND2_X1 u0_u13_u3_U82 (.A2( u0_u13_X_19 ) , .A1( u0_u13_X_20 ) , .ZN( u0_u13_u3_n104 ) );
  INV_X1 u0_u13_u3_U83 (.A( u0_u13_X_22 ) , .ZN( u0_u13_u3_n166 ) );
  INV_X1 u0_u13_u3_U84 (.A( u0_u13_X_21 ) , .ZN( u0_u13_u3_n171 ) );
  INV_X1 u0_u13_u3_U85 (.A( u0_u13_X_20 ) , .ZN( u0_u13_u3_n172 ) );
  NAND4_X1 u0_u13_u3_U86 (.ZN( u0_out13_26 ) , .A4( u0_u13_u3_n109 ) , .A3( u0_u13_u3_n110 ) , .A2( u0_u13_u3_n111 ) , .A1( u0_u13_u3_n173 ) );
  INV_X1 u0_u13_u3_U87 (.ZN( u0_u13_u3_n173 ) , .A( u0_u13_u3_n94 ) );
  OAI21_X1 u0_u13_u3_U88 (.ZN( u0_u13_u3_n111 ) , .B2( u0_u13_u3_n117 ) , .A( u0_u13_u3_n133 ) , .B1( u0_u13_u3_n176 ) );
  NAND4_X1 u0_u13_u3_U89 (.ZN( u0_out13_20 ) , .A4( u0_u13_u3_n122 ) , .A3( u0_u13_u3_n123 ) , .A1( u0_u13_u3_n175 ) , .A2( u0_u13_u3_n180 ) );
  INV_X1 u0_u13_u3_U9 (.A( u0_u13_u3_n143 ) , .ZN( u0_u13_u3_n168 ) );
  INV_X1 u0_u13_u3_U90 (.A( u0_u13_u3_n112 ) , .ZN( u0_u13_u3_n175 ) );
  INV_X1 u0_u13_u3_U91 (.A( u0_u13_u3_n126 ) , .ZN( u0_u13_u3_n180 ) );
  NAND4_X1 u0_u13_u3_U92 (.ZN( u0_out13_1 ) , .A4( u0_u13_u3_n161 ) , .A3( u0_u13_u3_n162 ) , .A2( u0_u13_u3_n163 ) , .A1( u0_u13_u3_n185 ) );
  NAND2_X1 u0_u13_u3_U93 (.ZN( u0_u13_u3_n163 ) , .A2( u0_u13_u3_n170 ) , .A1( u0_u13_u3_n176 ) );
  AOI22_X1 u0_u13_u3_U94 (.B2( u0_u13_u3_n140 ) , .B1( u0_u13_u3_n141 ) , .A2( u0_u13_u3_n142 ) , .ZN( u0_u13_u3_n162 ) , .A1( u0_u13_u3_n177 ) );
  OR4_X1 u0_u13_u3_U95 (.ZN( u0_out13_10 ) , .A4( u0_u13_u3_n136 ) , .A3( u0_u13_u3_n137 ) , .A1( u0_u13_u3_n138 ) , .A2( u0_u13_u3_n139 ) );
  OAI222_X1 u0_u13_u3_U96 (.C1( u0_u13_u3_n128 ) , .ZN( u0_u13_u3_n137 ) , .B1( u0_u13_u3_n148 ) , .A2( u0_u13_u3_n150 ) , .B2( u0_u13_u3_n154 ) , .C2( u0_u13_u3_n164 ) , .A1( u0_u13_u3_n167 ) );
  OAI221_X1 u0_u13_u3_U97 (.A( u0_u13_u3_n134 ) , .B2( u0_u13_u3_n135 ) , .ZN( u0_u13_u3_n136 ) , .C1( u0_u13_u3_n149 ) , .B1( u0_u13_u3_n151 ) , .C2( u0_u13_u3_n183 ) );
  NAND3_X1 u0_u13_u3_U98 (.A1( u0_u13_u3_n114 ) , .ZN( u0_u13_u3_n115 ) , .A2( u0_u13_u3_n145 ) , .A3( u0_u13_u3_n153 ) );
  NAND3_X1 u0_u13_u3_U99 (.ZN( u0_u13_u3_n129 ) , .A2( u0_u13_u3_n144 ) , .A1( u0_u13_u3_n153 ) , .A3( u0_u13_u3_n182 ) );
  AOI21_X1 u0_u13_u4_U10 (.ZN( u0_u13_u4_n106 ) , .B2( u0_u13_u4_n146 ) , .B1( u0_u13_u4_n158 ) , .A( u0_u13_u4_n170 ) );
  AOI21_X1 u0_u13_u4_U11 (.ZN( u0_u13_u4_n108 ) , .B2( u0_u13_u4_n134 ) , .B1( u0_u13_u4_n155 ) , .A( u0_u13_u4_n156 ) );
  AOI21_X1 u0_u13_u4_U12 (.ZN( u0_u13_u4_n109 ) , .A( u0_u13_u4_n153 ) , .B1( u0_u13_u4_n159 ) , .B2( u0_u13_u4_n184 ) );
  AOI211_X1 u0_u13_u4_U13 (.B( u0_u13_u4_n136 ) , .A( u0_u13_u4_n137 ) , .C2( u0_u13_u4_n138 ) , .ZN( u0_u13_u4_n139 ) , .C1( u0_u13_u4_n182 ) );
  OAI22_X1 u0_u13_u4_U14 (.B2( u0_u13_u4_n135 ) , .ZN( u0_u13_u4_n137 ) , .B1( u0_u13_u4_n153 ) , .A1( u0_u13_u4_n155 ) , .A2( u0_u13_u4_n171 ) );
  AND3_X1 u0_u13_u4_U15 (.A2( u0_u13_u4_n134 ) , .ZN( u0_u13_u4_n135 ) , .A3( u0_u13_u4_n145 ) , .A1( u0_u13_u4_n157 ) );
  NAND2_X1 u0_u13_u4_U16 (.ZN( u0_u13_u4_n132 ) , .A2( u0_u13_u4_n170 ) , .A1( u0_u13_u4_n173 ) );
  AOI21_X1 u0_u13_u4_U17 (.B2( u0_u13_u4_n160 ) , .B1( u0_u13_u4_n161 ) , .ZN( u0_u13_u4_n162 ) , .A( u0_u13_u4_n170 ) );
  AOI21_X1 u0_u13_u4_U18 (.ZN( u0_u13_u4_n107 ) , .B2( u0_u13_u4_n143 ) , .A( u0_u13_u4_n174 ) , .B1( u0_u13_u4_n184 ) );
  AOI21_X1 u0_u13_u4_U19 (.B2( u0_u13_u4_n158 ) , .B1( u0_u13_u4_n159 ) , .ZN( u0_u13_u4_n163 ) , .A( u0_u13_u4_n174 ) );
  AOI21_X1 u0_u13_u4_U20 (.A( u0_u13_u4_n153 ) , .B2( u0_u13_u4_n154 ) , .B1( u0_u13_u4_n155 ) , .ZN( u0_u13_u4_n165 ) );
  AOI21_X1 u0_u13_u4_U21 (.A( u0_u13_u4_n156 ) , .B2( u0_u13_u4_n157 ) , .ZN( u0_u13_u4_n164 ) , .B1( u0_u13_u4_n184 ) );
  INV_X1 u0_u13_u4_U22 (.A( u0_u13_u4_n138 ) , .ZN( u0_u13_u4_n170 ) );
  AND2_X1 u0_u13_u4_U23 (.A2( u0_u13_u4_n120 ) , .ZN( u0_u13_u4_n155 ) , .A1( u0_u13_u4_n160 ) );
  INV_X1 u0_u13_u4_U24 (.A( u0_u13_u4_n156 ) , .ZN( u0_u13_u4_n175 ) );
  NAND2_X1 u0_u13_u4_U25 (.A2( u0_u13_u4_n118 ) , .ZN( u0_u13_u4_n131 ) , .A1( u0_u13_u4_n147 ) );
  NAND2_X1 u0_u13_u4_U26 (.A1( u0_u13_u4_n119 ) , .A2( u0_u13_u4_n120 ) , .ZN( u0_u13_u4_n130 ) );
  NAND2_X1 u0_u13_u4_U27 (.ZN( u0_u13_u4_n117 ) , .A2( u0_u13_u4_n118 ) , .A1( u0_u13_u4_n148 ) );
  NAND2_X1 u0_u13_u4_U28 (.ZN( u0_u13_u4_n129 ) , .A1( u0_u13_u4_n134 ) , .A2( u0_u13_u4_n148 ) );
  AND3_X1 u0_u13_u4_U29 (.A1( u0_u13_u4_n119 ) , .A2( u0_u13_u4_n143 ) , .A3( u0_u13_u4_n154 ) , .ZN( u0_u13_u4_n161 ) );
  NOR2_X1 u0_u13_u4_U3 (.ZN( u0_u13_u4_n121 ) , .A1( u0_u13_u4_n181 ) , .A2( u0_u13_u4_n182 ) );
  AND2_X1 u0_u13_u4_U30 (.A1( u0_u13_u4_n145 ) , .A2( u0_u13_u4_n147 ) , .ZN( u0_u13_u4_n159 ) );
  OR3_X1 u0_u13_u4_U31 (.A3( u0_u13_u4_n114 ) , .A2( u0_u13_u4_n115 ) , .A1( u0_u13_u4_n116 ) , .ZN( u0_u13_u4_n136 ) );
  AOI21_X1 u0_u13_u4_U32 (.A( u0_u13_u4_n113 ) , .ZN( u0_u13_u4_n116 ) , .B2( u0_u13_u4_n173 ) , .B1( u0_u13_u4_n174 ) );
  AOI21_X1 u0_u13_u4_U33 (.ZN( u0_u13_u4_n115 ) , .B2( u0_u13_u4_n145 ) , .B1( u0_u13_u4_n146 ) , .A( u0_u13_u4_n156 ) );
  OAI22_X1 u0_u13_u4_U34 (.ZN( u0_u13_u4_n114 ) , .A2( u0_u13_u4_n121 ) , .B1( u0_u13_u4_n160 ) , .B2( u0_u13_u4_n170 ) , .A1( u0_u13_u4_n171 ) );
  INV_X1 u0_u13_u4_U35 (.A( u0_u13_u4_n158 ) , .ZN( u0_u13_u4_n182 ) );
  INV_X1 u0_u13_u4_U36 (.ZN( u0_u13_u4_n181 ) , .A( u0_u13_u4_n96 ) );
  INV_X1 u0_u13_u4_U37 (.A( u0_u13_u4_n144 ) , .ZN( u0_u13_u4_n179 ) );
  INV_X1 u0_u13_u4_U38 (.A( u0_u13_u4_n157 ) , .ZN( u0_u13_u4_n178 ) );
  NAND2_X1 u0_u13_u4_U39 (.A2( u0_u13_u4_n154 ) , .A1( u0_u13_u4_n96 ) , .ZN( u0_u13_u4_n97 ) );
  INV_X1 u0_u13_u4_U4 (.A( u0_u13_u4_n117 ) , .ZN( u0_u13_u4_n184 ) );
  INV_X1 u0_u13_u4_U40 (.A( u0_u13_u4_n143 ) , .ZN( u0_u13_u4_n183 ) );
  NOR2_X1 u0_u13_u4_U41 (.ZN( u0_u13_u4_n138 ) , .A1( u0_u13_u4_n168 ) , .A2( u0_u13_u4_n169 ) );
  NOR2_X1 u0_u13_u4_U42 (.A1( u0_u13_u4_n150 ) , .A2( u0_u13_u4_n152 ) , .ZN( u0_u13_u4_n153 ) );
  NOR2_X1 u0_u13_u4_U43 (.A2( u0_u13_u4_n128 ) , .A1( u0_u13_u4_n138 ) , .ZN( u0_u13_u4_n156 ) );
  AOI22_X1 u0_u13_u4_U44 (.B2( u0_u13_u4_n122 ) , .A1( u0_u13_u4_n123 ) , .ZN( u0_u13_u4_n124 ) , .B1( u0_u13_u4_n128 ) , .A2( u0_u13_u4_n172 ) );
  NAND2_X1 u0_u13_u4_U45 (.A2( u0_u13_u4_n120 ) , .ZN( u0_u13_u4_n123 ) , .A1( u0_u13_u4_n161 ) );
  INV_X1 u0_u13_u4_U46 (.A( u0_u13_u4_n153 ) , .ZN( u0_u13_u4_n172 ) );
  AOI22_X1 u0_u13_u4_U47 (.B2( u0_u13_u4_n132 ) , .A2( u0_u13_u4_n133 ) , .ZN( u0_u13_u4_n140 ) , .A1( u0_u13_u4_n150 ) , .B1( u0_u13_u4_n179 ) );
  NAND2_X1 u0_u13_u4_U48 (.ZN( u0_u13_u4_n133 ) , .A2( u0_u13_u4_n146 ) , .A1( u0_u13_u4_n154 ) );
  NAND2_X1 u0_u13_u4_U49 (.A1( u0_u13_u4_n103 ) , .ZN( u0_u13_u4_n154 ) , .A2( u0_u13_u4_n98 ) );
  INV_X1 u0_u13_u4_U5 (.ZN( u0_u13_u4_n186 ) , .A( u0_u13_u4_n95 ) );
  NAND2_X1 u0_u13_u4_U50 (.A1( u0_u13_u4_n101 ) , .ZN( u0_u13_u4_n158 ) , .A2( u0_u13_u4_n99 ) );
  AOI21_X1 u0_u13_u4_U51 (.ZN( u0_u13_u4_n127 ) , .A( u0_u13_u4_n136 ) , .B2( u0_u13_u4_n150 ) , .B1( u0_u13_u4_n180 ) );
  INV_X1 u0_u13_u4_U52 (.A( u0_u13_u4_n160 ) , .ZN( u0_u13_u4_n180 ) );
  NAND2_X1 u0_u13_u4_U53 (.A2( u0_u13_u4_n104 ) , .A1( u0_u13_u4_n105 ) , .ZN( u0_u13_u4_n146 ) );
  NAND2_X1 u0_u13_u4_U54 (.A2( u0_u13_u4_n101 ) , .A1( u0_u13_u4_n102 ) , .ZN( u0_u13_u4_n160 ) );
  NAND2_X1 u0_u13_u4_U55 (.ZN( u0_u13_u4_n134 ) , .A1( u0_u13_u4_n98 ) , .A2( u0_u13_u4_n99 ) );
  NAND2_X1 u0_u13_u4_U56 (.A1( u0_u13_u4_n103 ) , .A2( u0_u13_u4_n104 ) , .ZN( u0_u13_u4_n143 ) );
  NAND2_X1 u0_u13_u4_U57 (.A2( u0_u13_u4_n105 ) , .ZN( u0_u13_u4_n145 ) , .A1( u0_u13_u4_n98 ) );
  NAND2_X1 u0_u13_u4_U58 (.A1( u0_u13_u4_n100 ) , .A2( u0_u13_u4_n105 ) , .ZN( u0_u13_u4_n120 ) );
  NAND2_X1 u0_u13_u4_U59 (.A1( u0_u13_u4_n102 ) , .A2( u0_u13_u4_n104 ) , .ZN( u0_u13_u4_n148 ) );
  OAI221_X1 u0_u13_u4_U6 (.C1( u0_u13_u4_n134 ) , .B1( u0_u13_u4_n158 ) , .B2( u0_u13_u4_n171 ) , .C2( u0_u13_u4_n173 ) , .A( u0_u13_u4_n94 ) , .ZN( u0_u13_u4_n95 ) );
  NAND2_X1 u0_u13_u4_U60 (.A2( u0_u13_u4_n100 ) , .A1( u0_u13_u4_n103 ) , .ZN( u0_u13_u4_n157 ) );
  INV_X1 u0_u13_u4_U61 (.A( u0_u13_u4_n150 ) , .ZN( u0_u13_u4_n173 ) );
  INV_X1 u0_u13_u4_U62 (.A( u0_u13_u4_n152 ) , .ZN( u0_u13_u4_n171 ) );
  NAND2_X1 u0_u13_u4_U63 (.A1( u0_u13_u4_n100 ) , .ZN( u0_u13_u4_n118 ) , .A2( u0_u13_u4_n99 ) );
  NAND2_X1 u0_u13_u4_U64 (.A2( u0_u13_u4_n100 ) , .A1( u0_u13_u4_n102 ) , .ZN( u0_u13_u4_n144 ) );
  NAND2_X1 u0_u13_u4_U65 (.A2( u0_u13_u4_n101 ) , .A1( u0_u13_u4_n105 ) , .ZN( u0_u13_u4_n96 ) );
  INV_X1 u0_u13_u4_U66 (.A( u0_u13_u4_n128 ) , .ZN( u0_u13_u4_n174 ) );
  NAND2_X1 u0_u13_u4_U67 (.A2( u0_u13_u4_n102 ) , .ZN( u0_u13_u4_n119 ) , .A1( u0_u13_u4_n98 ) );
  NAND2_X1 u0_u13_u4_U68 (.A2( u0_u13_u4_n101 ) , .A1( u0_u13_u4_n103 ) , .ZN( u0_u13_u4_n147 ) );
  NAND2_X1 u0_u13_u4_U69 (.A2( u0_u13_u4_n104 ) , .ZN( u0_u13_u4_n113 ) , .A1( u0_u13_u4_n99 ) );
  AOI222_X1 u0_u13_u4_U7 (.B2( u0_u13_u4_n132 ) , .A1( u0_u13_u4_n138 ) , .C2( u0_u13_u4_n175 ) , .A2( u0_u13_u4_n179 ) , .C1( u0_u13_u4_n181 ) , .B1( u0_u13_u4_n185 ) , .ZN( u0_u13_u4_n94 ) );
  NOR2_X1 u0_u13_u4_U70 (.A2( u0_u13_X_28 ) , .ZN( u0_u13_u4_n150 ) , .A1( u0_u13_u4_n168 ) );
  NOR2_X1 u0_u13_u4_U71 (.A2( u0_u13_X_29 ) , .ZN( u0_u13_u4_n152 ) , .A1( u0_u13_u4_n169 ) );
  NOR2_X1 u0_u13_u4_U72 (.A2( u0_u13_X_30 ) , .ZN( u0_u13_u4_n105 ) , .A1( u0_u13_u4_n176 ) );
  NOR2_X1 u0_u13_u4_U73 (.A2( u0_u13_X_26 ) , .ZN( u0_u13_u4_n100 ) , .A1( u0_u13_u4_n177 ) );
  NOR2_X1 u0_u13_u4_U74 (.A2( u0_u13_X_28 ) , .A1( u0_u13_X_29 ) , .ZN( u0_u13_u4_n128 ) );
  NOR2_X1 u0_u13_u4_U75 (.A2( u0_u13_X_27 ) , .A1( u0_u13_X_30 ) , .ZN( u0_u13_u4_n102 ) );
  NOR2_X1 u0_u13_u4_U76 (.A2( u0_u13_X_25 ) , .A1( u0_u13_X_26 ) , .ZN( u0_u13_u4_n98 ) );
  AND2_X1 u0_u13_u4_U77 (.A2( u0_u13_X_25 ) , .A1( u0_u13_X_26 ) , .ZN( u0_u13_u4_n104 ) );
  AND2_X1 u0_u13_u4_U78 (.A1( u0_u13_X_30 ) , .A2( u0_u13_u4_n176 ) , .ZN( u0_u13_u4_n99 ) );
  AND2_X1 u0_u13_u4_U79 (.A1( u0_u13_X_26 ) , .ZN( u0_u13_u4_n101 ) , .A2( u0_u13_u4_n177 ) );
  INV_X1 u0_u13_u4_U8 (.A( u0_u13_u4_n113 ) , .ZN( u0_u13_u4_n185 ) );
  AND2_X1 u0_u13_u4_U80 (.A1( u0_u13_X_27 ) , .A2( u0_u13_X_30 ) , .ZN( u0_u13_u4_n103 ) );
  INV_X1 u0_u13_u4_U81 (.A( u0_u13_X_28 ) , .ZN( u0_u13_u4_n169 ) );
  INV_X1 u0_u13_u4_U82 (.A( u0_u13_X_29 ) , .ZN( u0_u13_u4_n168 ) );
  INV_X1 u0_u13_u4_U83 (.A( u0_u13_X_25 ) , .ZN( u0_u13_u4_n177 ) );
  INV_X1 u0_u13_u4_U84 (.A( u0_u13_X_27 ) , .ZN( u0_u13_u4_n176 ) );
  NAND4_X1 u0_u13_u4_U85 (.ZN( u0_out13_25 ) , .A4( u0_u13_u4_n139 ) , .A3( u0_u13_u4_n140 ) , .A2( u0_u13_u4_n141 ) , .A1( u0_u13_u4_n142 ) );
  OAI21_X1 u0_u13_u4_U86 (.A( u0_u13_u4_n128 ) , .B2( u0_u13_u4_n129 ) , .B1( u0_u13_u4_n130 ) , .ZN( u0_u13_u4_n142 ) );
  OAI21_X1 u0_u13_u4_U87 (.B2( u0_u13_u4_n131 ) , .ZN( u0_u13_u4_n141 ) , .A( u0_u13_u4_n175 ) , .B1( u0_u13_u4_n183 ) );
  NAND4_X1 u0_u13_u4_U88 (.ZN( u0_out13_14 ) , .A4( u0_u13_u4_n124 ) , .A3( u0_u13_u4_n125 ) , .A2( u0_u13_u4_n126 ) , .A1( u0_u13_u4_n127 ) );
  AOI22_X1 u0_u13_u4_U89 (.B2( u0_u13_u4_n117 ) , .ZN( u0_u13_u4_n126 ) , .A1( u0_u13_u4_n129 ) , .B1( u0_u13_u4_n152 ) , .A2( u0_u13_u4_n175 ) );
  NOR4_X1 u0_u13_u4_U9 (.A4( u0_u13_u4_n106 ) , .A3( u0_u13_u4_n107 ) , .A2( u0_u13_u4_n108 ) , .A1( u0_u13_u4_n109 ) , .ZN( u0_u13_u4_n110 ) );
  AOI22_X1 u0_u13_u4_U90 (.ZN( u0_u13_u4_n125 ) , .B2( u0_u13_u4_n131 ) , .A2( u0_u13_u4_n132 ) , .B1( u0_u13_u4_n138 ) , .A1( u0_u13_u4_n178 ) );
  NAND4_X1 u0_u13_u4_U91 (.ZN( u0_out13_8 ) , .A4( u0_u13_u4_n110 ) , .A3( u0_u13_u4_n111 ) , .A2( u0_u13_u4_n112 ) , .A1( u0_u13_u4_n186 ) );
  NAND2_X1 u0_u13_u4_U92 (.ZN( u0_u13_u4_n112 ) , .A2( u0_u13_u4_n130 ) , .A1( u0_u13_u4_n150 ) );
  AOI22_X1 u0_u13_u4_U93 (.ZN( u0_u13_u4_n111 ) , .B2( u0_u13_u4_n132 ) , .A1( u0_u13_u4_n152 ) , .B1( u0_u13_u4_n178 ) , .A2( u0_u13_u4_n97 ) );
  AOI22_X1 u0_u13_u4_U94 (.B2( u0_u13_u4_n149 ) , .B1( u0_u13_u4_n150 ) , .A2( u0_u13_u4_n151 ) , .A1( u0_u13_u4_n152 ) , .ZN( u0_u13_u4_n167 ) );
  NOR4_X1 u0_u13_u4_U95 (.A4( u0_u13_u4_n162 ) , .A3( u0_u13_u4_n163 ) , .A2( u0_u13_u4_n164 ) , .A1( u0_u13_u4_n165 ) , .ZN( u0_u13_u4_n166 ) );
  NAND3_X1 u0_u13_u4_U96 (.ZN( u0_out13_3 ) , .A3( u0_u13_u4_n166 ) , .A1( u0_u13_u4_n167 ) , .A2( u0_u13_u4_n186 ) );
  NAND3_X1 u0_u13_u4_U97 (.A3( u0_u13_u4_n146 ) , .A2( u0_u13_u4_n147 ) , .A1( u0_u13_u4_n148 ) , .ZN( u0_u13_u4_n149 ) );
  NAND3_X1 u0_u13_u4_U98 (.A3( u0_u13_u4_n143 ) , .A2( u0_u13_u4_n144 ) , .A1( u0_u13_u4_n145 ) , .ZN( u0_u13_u4_n151 ) );
  NAND3_X1 u0_u13_u4_U99 (.A3( u0_u13_u4_n121 ) , .ZN( u0_u13_u4_n122 ) , .A2( u0_u13_u4_n144 ) , .A1( u0_u13_u4_n154 ) );
  INV_X1 u0_u13_u5_U10 (.A( u0_u13_u5_n121 ) , .ZN( u0_u13_u5_n177 ) );
  NOR3_X1 u0_u13_u5_U100 (.A3( u0_u13_u5_n141 ) , .A1( u0_u13_u5_n142 ) , .ZN( u0_u13_u5_n143 ) , .A2( u0_u13_u5_n191 ) );
  NAND4_X1 u0_u13_u5_U101 (.ZN( u0_out13_4 ) , .A4( u0_u13_u5_n112 ) , .A2( u0_u13_u5_n113 ) , .A1( u0_u13_u5_n114 ) , .A3( u0_u13_u5_n195 ) );
  AOI211_X1 u0_u13_u5_U102 (.A( u0_u13_u5_n110 ) , .C1( u0_u13_u5_n111 ) , .ZN( u0_u13_u5_n112 ) , .B( u0_u13_u5_n118 ) , .C2( u0_u13_u5_n177 ) );
  AOI222_X1 u0_u13_u5_U103 (.ZN( u0_u13_u5_n113 ) , .A1( u0_u13_u5_n131 ) , .C1( u0_u13_u5_n148 ) , .B2( u0_u13_u5_n174 ) , .C2( u0_u13_u5_n178 ) , .A2( u0_u13_u5_n179 ) , .B1( u0_u13_u5_n99 ) );
  NAND3_X1 u0_u13_u5_U104 (.A2( u0_u13_u5_n154 ) , .A3( u0_u13_u5_n158 ) , .A1( u0_u13_u5_n161 ) , .ZN( u0_u13_u5_n99 ) );
  NOR2_X1 u0_u13_u5_U11 (.ZN( u0_u13_u5_n160 ) , .A2( u0_u13_u5_n173 ) , .A1( u0_u13_u5_n177 ) );
  INV_X1 u0_u13_u5_U12 (.A( u0_u13_u5_n150 ) , .ZN( u0_u13_u5_n174 ) );
  AOI21_X1 u0_u13_u5_U13 (.A( u0_u13_u5_n160 ) , .B2( u0_u13_u5_n161 ) , .ZN( u0_u13_u5_n162 ) , .B1( u0_u13_u5_n192 ) );
  INV_X1 u0_u13_u5_U14 (.A( u0_u13_u5_n159 ) , .ZN( u0_u13_u5_n192 ) );
  AOI21_X1 u0_u13_u5_U15 (.A( u0_u13_u5_n156 ) , .B2( u0_u13_u5_n157 ) , .B1( u0_u13_u5_n158 ) , .ZN( u0_u13_u5_n163 ) );
  AOI21_X1 u0_u13_u5_U16 (.B2( u0_u13_u5_n139 ) , .B1( u0_u13_u5_n140 ) , .ZN( u0_u13_u5_n141 ) , .A( u0_u13_u5_n150 ) );
  OAI21_X1 u0_u13_u5_U17 (.A( u0_u13_u5_n133 ) , .B2( u0_u13_u5_n134 ) , .B1( u0_u13_u5_n135 ) , .ZN( u0_u13_u5_n142 ) );
  OAI21_X1 u0_u13_u5_U18 (.ZN( u0_u13_u5_n133 ) , .B2( u0_u13_u5_n147 ) , .A( u0_u13_u5_n173 ) , .B1( u0_u13_u5_n188 ) );
  NAND2_X1 u0_u13_u5_U19 (.A2( u0_u13_u5_n119 ) , .A1( u0_u13_u5_n123 ) , .ZN( u0_u13_u5_n137 ) );
  INV_X1 u0_u13_u5_U20 (.A( u0_u13_u5_n155 ) , .ZN( u0_u13_u5_n194 ) );
  NAND2_X1 u0_u13_u5_U21 (.A1( u0_u13_u5_n121 ) , .ZN( u0_u13_u5_n132 ) , .A2( u0_u13_u5_n172 ) );
  NAND2_X1 u0_u13_u5_U22 (.A2( u0_u13_u5_n122 ) , .ZN( u0_u13_u5_n136 ) , .A1( u0_u13_u5_n154 ) );
  NAND2_X1 u0_u13_u5_U23 (.A2( u0_u13_u5_n119 ) , .A1( u0_u13_u5_n120 ) , .ZN( u0_u13_u5_n159 ) );
  INV_X1 u0_u13_u5_U24 (.A( u0_u13_u5_n156 ) , .ZN( u0_u13_u5_n175 ) );
  INV_X1 u0_u13_u5_U25 (.A( u0_u13_u5_n158 ) , .ZN( u0_u13_u5_n188 ) );
  INV_X1 u0_u13_u5_U26 (.A( u0_u13_u5_n152 ) , .ZN( u0_u13_u5_n179 ) );
  INV_X1 u0_u13_u5_U27 (.A( u0_u13_u5_n140 ) , .ZN( u0_u13_u5_n182 ) );
  INV_X1 u0_u13_u5_U28 (.A( u0_u13_u5_n151 ) , .ZN( u0_u13_u5_n183 ) );
  INV_X1 u0_u13_u5_U29 (.A( u0_u13_u5_n123 ) , .ZN( u0_u13_u5_n185 ) );
  NOR2_X1 u0_u13_u5_U3 (.ZN( u0_u13_u5_n134 ) , .A1( u0_u13_u5_n183 ) , .A2( u0_u13_u5_n190 ) );
  INV_X1 u0_u13_u5_U30 (.A( u0_u13_u5_n161 ) , .ZN( u0_u13_u5_n184 ) );
  INV_X1 u0_u13_u5_U31 (.A( u0_u13_u5_n139 ) , .ZN( u0_u13_u5_n189 ) );
  INV_X1 u0_u13_u5_U32 (.A( u0_u13_u5_n157 ) , .ZN( u0_u13_u5_n190 ) );
  INV_X1 u0_u13_u5_U33 (.A( u0_u13_u5_n120 ) , .ZN( u0_u13_u5_n193 ) );
  NAND2_X1 u0_u13_u5_U34 (.ZN( u0_u13_u5_n111 ) , .A1( u0_u13_u5_n140 ) , .A2( u0_u13_u5_n155 ) );
  INV_X1 u0_u13_u5_U35 (.A( u0_u13_u5_n117 ) , .ZN( u0_u13_u5_n196 ) );
  OAI221_X1 u0_u13_u5_U36 (.A( u0_u13_u5_n116 ) , .ZN( u0_u13_u5_n117 ) , .B2( u0_u13_u5_n119 ) , .C1( u0_u13_u5_n153 ) , .C2( u0_u13_u5_n158 ) , .B1( u0_u13_u5_n172 ) );
  AOI222_X1 u0_u13_u5_U37 (.ZN( u0_u13_u5_n116 ) , .B2( u0_u13_u5_n145 ) , .C1( u0_u13_u5_n148 ) , .A2( u0_u13_u5_n174 ) , .C2( u0_u13_u5_n177 ) , .B1( u0_u13_u5_n187 ) , .A1( u0_u13_u5_n193 ) );
  INV_X1 u0_u13_u5_U38 (.A( u0_u13_u5_n115 ) , .ZN( u0_u13_u5_n187 ) );
  NOR2_X1 u0_u13_u5_U39 (.ZN( u0_u13_u5_n100 ) , .A1( u0_u13_u5_n170 ) , .A2( u0_u13_u5_n180 ) );
  INV_X1 u0_u13_u5_U4 (.A( u0_u13_u5_n138 ) , .ZN( u0_u13_u5_n191 ) );
  AOI22_X1 u0_u13_u5_U40 (.B2( u0_u13_u5_n131 ) , .A2( u0_u13_u5_n146 ) , .ZN( u0_u13_u5_n169 ) , .B1( u0_u13_u5_n174 ) , .A1( u0_u13_u5_n185 ) );
  NOR2_X1 u0_u13_u5_U41 (.A1( u0_u13_u5_n146 ) , .ZN( u0_u13_u5_n150 ) , .A2( u0_u13_u5_n173 ) );
  AOI21_X1 u0_u13_u5_U42 (.A( u0_u13_u5_n118 ) , .B2( u0_u13_u5_n145 ) , .ZN( u0_u13_u5_n168 ) , .B1( u0_u13_u5_n186 ) );
  INV_X1 u0_u13_u5_U43 (.A( u0_u13_u5_n122 ) , .ZN( u0_u13_u5_n186 ) );
  NOR2_X1 u0_u13_u5_U44 (.A1( u0_u13_u5_n146 ) , .ZN( u0_u13_u5_n152 ) , .A2( u0_u13_u5_n176 ) );
  NOR2_X1 u0_u13_u5_U45 (.A1( u0_u13_u5_n115 ) , .ZN( u0_u13_u5_n118 ) , .A2( u0_u13_u5_n153 ) );
  NOR2_X1 u0_u13_u5_U46 (.A2( u0_u13_u5_n145 ) , .ZN( u0_u13_u5_n156 ) , .A1( u0_u13_u5_n174 ) );
  NOR2_X1 u0_u13_u5_U47 (.ZN( u0_u13_u5_n121 ) , .A2( u0_u13_u5_n145 ) , .A1( u0_u13_u5_n176 ) );
  AOI22_X1 u0_u13_u5_U48 (.ZN( u0_u13_u5_n114 ) , .A2( u0_u13_u5_n137 ) , .A1( u0_u13_u5_n145 ) , .B2( u0_u13_u5_n175 ) , .B1( u0_u13_u5_n193 ) );
  OAI211_X1 u0_u13_u5_U49 (.B( u0_u13_u5_n124 ) , .A( u0_u13_u5_n125 ) , .C2( u0_u13_u5_n126 ) , .C1( u0_u13_u5_n127 ) , .ZN( u0_u13_u5_n128 ) );
  OAI21_X1 u0_u13_u5_U5 (.B2( u0_u13_u5_n136 ) , .B1( u0_u13_u5_n137 ) , .ZN( u0_u13_u5_n138 ) , .A( u0_u13_u5_n177 ) );
  NOR3_X1 u0_u13_u5_U50 (.ZN( u0_u13_u5_n127 ) , .A1( u0_u13_u5_n136 ) , .A3( u0_u13_u5_n148 ) , .A2( u0_u13_u5_n182 ) );
  OAI21_X1 u0_u13_u5_U51 (.ZN( u0_u13_u5_n124 ) , .A( u0_u13_u5_n177 ) , .B2( u0_u13_u5_n183 ) , .B1( u0_u13_u5_n189 ) );
  OAI21_X1 u0_u13_u5_U52 (.ZN( u0_u13_u5_n125 ) , .A( u0_u13_u5_n174 ) , .B2( u0_u13_u5_n185 ) , .B1( u0_u13_u5_n190 ) );
  AOI21_X1 u0_u13_u5_U53 (.A( u0_u13_u5_n153 ) , .B2( u0_u13_u5_n154 ) , .B1( u0_u13_u5_n155 ) , .ZN( u0_u13_u5_n164 ) );
  AOI21_X1 u0_u13_u5_U54 (.ZN( u0_u13_u5_n110 ) , .B1( u0_u13_u5_n122 ) , .B2( u0_u13_u5_n139 ) , .A( u0_u13_u5_n153 ) );
  INV_X1 u0_u13_u5_U55 (.A( u0_u13_u5_n153 ) , .ZN( u0_u13_u5_n176 ) );
  INV_X1 u0_u13_u5_U56 (.A( u0_u13_u5_n126 ) , .ZN( u0_u13_u5_n173 ) );
  AND2_X1 u0_u13_u5_U57 (.A2( u0_u13_u5_n104 ) , .A1( u0_u13_u5_n107 ) , .ZN( u0_u13_u5_n147 ) );
  AND2_X1 u0_u13_u5_U58 (.A2( u0_u13_u5_n104 ) , .A1( u0_u13_u5_n108 ) , .ZN( u0_u13_u5_n148 ) );
  NAND2_X1 u0_u13_u5_U59 (.A1( u0_u13_u5_n105 ) , .A2( u0_u13_u5_n106 ) , .ZN( u0_u13_u5_n158 ) );
  INV_X1 u0_u13_u5_U6 (.A( u0_u13_u5_n135 ) , .ZN( u0_u13_u5_n178 ) );
  NAND2_X1 u0_u13_u5_U60 (.A2( u0_u13_u5_n108 ) , .A1( u0_u13_u5_n109 ) , .ZN( u0_u13_u5_n139 ) );
  NAND2_X1 u0_u13_u5_U61 (.A1( u0_u13_u5_n106 ) , .A2( u0_u13_u5_n108 ) , .ZN( u0_u13_u5_n119 ) );
  NAND2_X1 u0_u13_u5_U62 (.A2( u0_u13_u5_n103 ) , .A1( u0_u13_u5_n105 ) , .ZN( u0_u13_u5_n140 ) );
  NAND2_X1 u0_u13_u5_U63 (.A2( u0_u13_u5_n104 ) , .A1( u0_u13_u5_n105 ) , .ZN( u0_u13_u5_n155 ) );
  NAND2_X1 u0_u13_u5_U64 (.A2( u0_u13_u5_n106 ) , .A1( u0_u13_u5_n107 ) , .ZN( u0_u13_u5_n122 ) );
  NAND2_X1 u0_u13_u5_U65 (.A2( u0_u13_u5_n100 ) , .A1( u0_u13_u5_n106 ) , .ZN( u0_u13_u5_n115 ) );
  NAND2_X1 u0_u13_u5_U66 (.A2( u0_u13_u5_n100 ) , .A1( u0_u13_u5_n103 ) , .ZN( u0_u13_u5_n161 ) );
  NAND2_X1 u0_u13_u5_U67 (.A1( u0_u13_u5_n105 ) , .A2( u0_u13_u5_n109 ) , .ZN( u0_u13_u5_n154 ) );
  INV_X1 u0_u13_u5_U68 (.A( u0_u13_u5_n146 ) , .ZN( u0_u13_u5_n172 ) );
  NAND2_X1 u0_u13_u5_U69 (.A1( u0_u13_u5_n103 ) , .A2( u0_u13_u5_n108 ) , .ZN( u0_u13_u5_n123 ) );
  OAI22_X1 u0_u13_u5_U7 (.B2( u0_u13_u5_n149 ) , .B1( u0_u13_u5_n150 ) , .A2( u0_u13_u5_n151 ) , .A1( u0_u13_u5_n152 ) , .ZN( u0_u13_u5_n165 ) );
  NAND2_X1 u0_u13_u5_U70 (.A2( u0_u13_u5_n103 ) , .A1( u0_u13_u5_n107 ) , .ZN( u0_u13_u5_n151 ) );
  NAND2_X1 u0_u13_u5_U71 (.A2( u0_u13_u5_n107 ) , .A1( u0_u13_u5_n109 ) , .ZN( u0_u13_u5_n120 ) );
  NAND2_X1 u0_u13_u5_U72 (.A2( u0_u13_u5_n100 ) , .A1( u0_u13_u5_n109 ) , .ZN( u0_u13_u5_n157 ) );
  AND2_X1 u0_u13_u5_U73 (.A2( u0_u13_u5_n100 ) , .A1( u0_u13_u5_n104 ) , .ZN( u0_u13_u5_n131 ) );
  INV_X1 u0_u13_u5_U74 (.A( u0_u13_u5_n102 ) , .ZN( u0_u13_u5_n195 ) );
  OAI221_X1 u0_u13_u5_U75 (.A( u0_u13_u5_n101 ) , .ZN( u0_u13_u5_n102 ) , .C2( u0_u13_u5_n115 ) , .C1( u0_u13_u5_n126 ) , .B1( u0_u13_u5_n134 ) , .B2( u0_u13_u5_n160 ) );
  OAI21_X1 u0_u13_u5_U76 (.ZN( u0_u13_u5_n101 ) , .B1( u0_u13_u5_n137 ) , .A( u0_u13_u5_n146 ) , .B2( u0_u13_u5_n147 ) );
  NOR2_X1 u0_u13_u5_U77 (.A2( u0_u13_X_34 ) , .A1( u0_u13_X_35 ) , .ZN( u0_u13_u5_n145 ) );
  NOR2_X1 u0_u13_u5_U78 (.A2( u0_u13_X_34 ) , .ZN( u0_u13_u5_n146 ) , .A1( u0_u13_u5_n171 ) );
  NOR2_X1 u0_u13_u5_U79 (.A2( u0_u13_X_31 ) , .A1( u0_u13_X_32 ) , .ZN( u0_u13_u5_n103 ) );
  NOR3_X1 u0_u13_u5_U8 (.A2( u0_u13_u5_n147 ) , .A1( u0_u13_u5_n148 ) , .ZN( u0_u13_u5_n149 ) , .A3( u0_u13_u5_n194 ) );
  NOR2_X1 u0_u13_u5_U80 (.A2( u0_u13_X_36 ) , .ZN( u0_u13_u5_n105 ) , .A1( u0_u13_u5_n180 ) );
  NOR2_X1 u0_u13_u5_U81 (.A2( u0_u13_X_33 ) , .ZN( u0_u13_u5_n108 ) , .A1( u0_u13_u5_n170 ) );
  NOR2_X1 u0_u13_u5_U82 (.A2( u0_u13_X_33 ) , .A1( u0_u13_X_36 ) , .ZN( u0_u13_u5_n107 ) );
  NOR2_X1 u0_u13_u5_U83 (.A2( u0_u13_X_31 ) , .ZN( u0_u13_u5_n104 ) , .A1( u0_u13_u5_n181 ) );
  NAND2_X1 u0_u13_u5_U84 (.A2( u0_u13_X_34 ) , .A1( u0_u13_X_35 ) , .ZN( u0_u13_u5_n153 ) );
  NAND2_X1 u0_u13_u5_U85 (.A1( u0_u13_X_34 ) , .ZN( u0_u13_u5_n126 ) , .A2( u0_u13_u5_n171 ) );
  AND2_X1 u0_u13_u5_U86 (.A1( u0_u13_X_31 ) , .A2( u0_u13_X_32 ) , .ZN( u0_u13_u5_n106 ) );
  AND2_X1 u0_u13_u5_U87 (.A1( u0_u13_X_31 ) , .ZN( u0_u13_u5_n109 ) , .A2( u0_u13_u5_n181 ) );
  INV_X1 u0_u13_u5_U88 (.A( u0_u13_X_33 ) , .ZN( u0_u13_u5_n180 ) );
  INV_X1 u0_u13_u5_U89 (.A( u0_u13_X_35 ) , .ZN( u0_u13_u5_n171 ) );
  NOR2_X1 u0_u13_u5_U9 (.ZN( u0_u13_u5_n135 ) , .A1( u0_u13_u5_n173 ) , .A2( u0_u13_u5_n176 ) );
  INV_X1 u0_u13_u5_U90 (.A( u0_u13_X_36 ) , .ZN( u0_u13_u5_n170 ) );
  INV_X1 u0_u13_u5_U91 (.A( u0_u13_X_32 ) , .ZN( u0_u13_u5_n181 ) );
  NAND4_X1 u0_u13_u5_U92 (.ZN( u0_out13_29 ) , .A4( u0_u13_u5_n129 ) , .A3( u0_u13_u5_n130 ) , .A2( u0_u13_u5_n168 ) , .A1( u0_u13_u5_n196 ) );
  AOI221_X1 u0_u13_u5_U93 (.A( u0_u13_u5_n128 ) , .ZN( u0_u13_u5_n129 ) , .C2( u0_u13_u5_n132 ) , .B2( u0_u13_u5_n159 ) , .B1( u0_u13_u5_n176 ) , .C1( u0_u13_u5_n184 ) );
  AOI222_X1 u0_u13_u5_U94 (.ZN( u0_u13_u5_n130 ) , .A2( u0_u13_u5_n146 ) , .B1( u0_u13_u5_n147 ) , .C2( u0_u13_u5_n175 ) , .B2( u0_u13_u5_n179 ) , .A1( u0_u13_u5_n188 ) , .C1( u0_u13_u5_n194 ) );
  NAND4_X1 u0_u13_u5_U95 (.ZN( u0_out13_19 ) , .A4( u0_u13_u5_n166 ) , .A3( u0_u13_u5_n167 ) , .A2( u0_u13_u5_n168 ) , .A1( u0_u13_u5_n169 ) );
  AOI22_X1 u0_u13_u5_U96 (.B2( u0_u13_u5_n145 ) , .A2( u0_u13_u5_n146 ) , .ZN( u0_u13_u5_n167 ) , .B1( u0_u13_u5_n182 ) , .A1( u0_u13_u5_n189 ) );
  NOR4_X1 u0_u13_u5_U97 (.A4( u0_u13_u5_n162 ) , .A3( u0_u13_u5_n163 ) , .A2( u0_u13_u5_n164 ) , .A1( u0_u13_u5_n165 ) , .ZN( u0_u13_u5_n166 ) );
  NAND4_X1 u0_u13_u5_U98 (.ZN( u0_out13_11 ) , .A4( u0_u13_u5_n143 ) , .A3( u0_u13_u5_n144 ) , .A2( u0_u13_u5_n169 ) , .A1( u0_u13_u5_n196 ) );
  AOI22_X1 u0_u13_u5_U99 (.A2( u0_u13_u5_n132 ) , .ZN( u0_u13_u5_n144 ) , .B2( u0_u13_u5_n145 ) , .B1( u0_u13_u5_n184 ) , .A1( u0_u13_u5_n194 ) );
  AOI22_X1 u0_u13_u6_U10 (.A2( u0_u13_u6_n151 ) , .B2( u0_u13_u6_n161 ) , .A1( u0_u13_u6_n167 ) , .B1( u0_u13_u6_n170 ) , .ZN( u0_u13_u6_n89 ) );
  AOI21_X1 u0_u13_u6_U11 (.B1( u0_u13_u6_n107 ) , .B2( u0_u13_u6_n132 ) , .A( u0_u13_u6_n158 ) , .ZN( u0_u13_u6_n88 ) );
  AOI21_X1 u0_u13_u6_U12 (.B2( u0_u13_u6_n147 ) , .B1( u0_u13_u6_n148 ) , .ZN( u0_u13_u6_n149 ) , .A( u0_u13_u6_n158 ) );
  AOI21_X1 u0_u13_u6_U13 (.ZN( u0_u13_u6_n106 ) , .A( u0_u13_u6_n142 ) , .B2( u0_u13_u6_n159 ) , .B1( u0_u13_u6_n164 ) );
  INV_X1 u0_u13_u6_U14 (.A( u0_u13_u6_n155 ) , .ZN( u0_u13_u6_n161 ) );
  INV_X1 u0_u13_u6_U15 (.A( u0_u13_u6_n128 ) , .ZN( u0_u13_u6_n164 ) );
  NAND2_X1 u0_u13_u6_U16 (.ZN( u0_u13_u6_n110 ) , .A1( u0_u13_u6_n122 ) , .A2( u0_u13_u6_n129 ) );
  NAND2_X1 u0_u13_u6_U17 (.ZN( u0_u13_u6_n124 ) , .A2( u0_u13_u6_n146 ) , .A1( u0_u13_u6_n148 ) );
  INV_X1 u0_u13_u6_U18 (.A( u0_u13_u6_n132 ) , .ZN( u0_u13_u6_n171 ) );
  AND2_X1 u0_u13_u6_U19 (.A1( u0_u13_u6_n100 ) , .ZN( u0_u13_u6_n130 ) , .A2( u0_u13_u6_n147 ) );
  INV_X1 u0_u13_u6_U20 (.A( u0_u13_u6_n127 ) , .ZN( u0_u13_u6_n173 ) );
  INV_X1 u0_u13_u6_U21 (.A( u0_u13_u6_n121 ) , .ZN( u0_u13_u6_n167 ) );
  INV_X1 u0_u13_u6_U22 (.A( u0_u13_u6_n100 ) , .ZN( u0_u13_u6_n169 ) );
  INV_X1 u0_u13_u6_U23 (.A( u0_u13_u6_n123 ) , .ZN( u0_u13_u6_n170 ) );
  INV_X1 u0_u13_u6_U24 (.A( u0_u13_u6_n113 ) , .ZN( u0_u13_u6_n168 ) );
  AND2_X1 u0_u13_u6_U25 (.A1( u0_u13_u6_n107 ) , .A2( u0_u13_u6_n119 ) , .ZN( u0_u13_u6_n133 ) );
  AND2_X1 u0_u13_u6_U26 (.A2( u0_u13_u6_n121 ) , .A1( u0_u13_u6_n122 ) , .ZN( u0_u13_u6_n131 ) );
  AND3_X1 u0_u13_u6_U27 (.ZN( u0_u13_u6_n120 ) , .A2( u0_u13_u6_n127 ) , .A1( u0_u13_u6_n132 ) , .A3( u0_u13_u6_n145 ) );
  INV_X1 u0_u13_u6_U28 (.A( u0_u13_u6_n146 ) , .ZN( u0_u13_u6_n163 ) );
  AOI222_X1 u0_u13_u6_U29 (.ZN( u0_u13_u6_n114 ) , .A1( u0_u13_u6_n118 ) , .A2( u0_u13_u6_n126 ) , .B2( u0_u13_u6_n151 ) , .C2( u0_u13_u6_n159 ) , .C1( u0_u13_u6_n168 ) , .B1( u0_u13_u6_n169 ) );
  INV_X1 u0_u13_u6_U3 (.A( u0_u13_u6_n110 ) , .ZN( u0_u13_u6_n166 ) );
  NOR2_X1 u0_u13_u6_U30 (.A1( u0_u13_u6_n162 ) , .A2( u0_u13_u6_n165 ) , .ZN( u0_u13_u6_n98 ) );
  AOI211_X1 u0_u13_u6_U31 (.B( u0_u13_u6_n134 ) , .A( u0_u13_u6_n135 ) , .C1( u0_u13_u6_n136 ) , .ZN( u0_u13_u6_n137 ) , .C2( u0_u13_u6_n151 ) );
  AOI21_X1 u0_u13_u6_U32 (.B2( u0_u13_u6_n132 ) , .B1( u0_u13_u6_n133 ) , .ZN( u0_u13_u6_n134 ) , .A( u0_u13_u6_n158 ) );
  AOI21_X1 u0_u13_u6_U33 (.B1( u0_u13_u6_n131 ) , .ZN( u0_u13_u6_n135 ) , .A( u0_u13_u6_n144 ) , .B2( u0_u13_u6_n146 ) );
  NAND4_X1 u0_u13_u6_U34 (.A4( u0_u13_u6_n127 ) , .A3( u0_u13_u6_n128 ) , .A2( u0_u13_u6_n129 ) , .A1( u0_u13_u6_n130 ) , .ZN( u0_u13_u6_n136 ) );
  NAND2_X1 u0_u13_u6_U35 (.A1( u0_u13_u6_n144 ) , .ZN( u0_u13_u6_n151 ) , .A2( u0_u13_u6_n158 ) );
  NAND2_X1 u0_u13_u6_U36 (.ZN( u0_u13_u6_n132 ) , .A1( u0_u13_u6_n91 ) , .A2( u0_u13_u6_n97 ) );
  AOI22_X1 u0_u13_u6_U37 (.B2( u0_u13_u6_n110 ) , .B1( u0_u13_u6_n111 ) , .A1( u0_u13_u6_n112 ) , .ZN( u0_u13_u6_n115 ) , .A2( u0_u13_u6_n161 ) );
  NAND4_X1 u0_u13_u6_U38 (.A3( u0_u13_u6_n109 ) , .ZN( u0_u13_u6_n112 ) , .A4( u0_u13_u6_n132 ) , .A2( u0_u13_u6_n147 ) , .A1( u0_u13_u6_n166 ) );
  NOR2_X1 u0_u13_u6_U39 (.ZN( u0_u13_u6_n109 ) , .A1( u0_u13_u6_n170 ) , .A2( u0_u13_u6_n173 ) );
  INV_X1 u0_u13_u6_U4 (.A( u0_u13_u6_n142 ) , .ZN( u0_u13_u6_n174 ) );
  NOR2_X1 u0_u13_u6_U40 (.A2( u0_u13_u6_n126 ) , .ZN( u0_u13_u6_n155 ) , .A1( u0_u13_u6_n160 ) );
  NAND2_X1 u0_u13_u6_U41 (.ZN( u0_u13_u6_n146 ) , .A2( u0_u13_u6_n94 ) , .A1( u0_u13_u6_n99 ) );
  AOI21_X1 u0_u13_u6_U42 (.A( u0_u13_u6_n144 ) , .B2( u0_u13_u6_n145 ) , .B1( u0_u13_u6_n146 ) , .ZN( u0_u13_u6_n150 ) );
  INV_X1 u0_u13_u6_U43 (.A( u0_u13_u6_n111 ) , .ZN( u0_u13_u6_n158 ) );
  NAND2_X1 u0_u13_u6_U44 (.ZN( u0_u13_u6_n127 ) , .A1( u0_u13_u6_n91 ) , .A2( u0_u13_u6_n92 ) );
  NAND2_X1 u0_u13_u6_U45 (.ZN( u0_u13_u6_n129 ) , .A2( u0_u13_u6_n95 ) , .A1( u0_u13_u6_n96 ) );
  INV_X1 u0_u13_u6_U46 (.A( u0_u13_u6_n144 ) , .ZN( u0_u13_u6_n159 ) );
  NAND2_X1 u0_u13_u6_U47 (.ZN( u0_u13_u6_n145 ) , .A2( u0_u13_u6_n97 ) , .A1( u0_u13_u6_n98 ) );
  NAND2_X1 u0_u13_u6_U48 (.ZN( u0_u13_u6_n148 ) , .A2( u0_u13_u6_n92 ) , .A1( u0_u13_u6_n94 ) );
  NAND2_X1 u0_u13_u6_U49 (.ZN( u0_u13_u6_n108 ) , .A2( u0_u13_u6_n139 ) , .A1( u0_u13_u6_n144 ) );
  NAND2_X1 u0_u13_u6_U5 (.A2( u0_u13_u6_n143 ) , .ZN( u0_u13_u6_n152 ) , .A1( u0_u13_u6_n166 ) );
  NAND2_X1 u0_u13_u6_U50 (.ZN( u0_u13_u6_n121 ) , .A2( u0_u13_u6_n95 ) , .A1( u0_u13_u6_n97 ) );
  NAND2_X1 u0_u13_u6_U51 (.ZN( u0_u13_u6_n107 ) , .A2( u0_u13_u6_n92 ) , .A1( u0_u13_u6_n95 ) );
  AND2_X1 u0_u13_u6_U52 (.ZN( u0_u13_u6_n118 ) , .A2( u0_u13_u6_n91 ) , .A1( u0_u13_u6_n99 ) );
  NAND2_X1 u0_u13_u6_U53 (.ZN( u0_u13_u6_n147 ) , .A2( u0_u13_u6_n98 ) , .A1( u0_u13_u6_n99 ) );
  NAND2_X1 u0_u13_u6_U54 (.ZN( u0_u13_u6_n128 ) , .A1( u0_u13_u6_n94 ) , .A2( u0_u13_u6_n96 ) );
  NAND2_X1 u0_u13_u6_U55 (.ZN( u0_u13_u6_n119 ) , .A2( u0_u13_u6_n95 ) , .A1( u0_u13_u6_n99 ) );
  NAND2_X1 u0_u13_u6_U56 (.ZN( u0_u13_u6_n123 ) , .A2( u0_u13_u6_n91 ) , .A1( u0_u13_u6_n96 ) );
  NAND2_X1 u0_u13_u6_U57 (.ZN( u0_u13_u6_n100 ) , .A2( u0_u13_u6_n92 ) , .A1( u0_u13_u6_n98 ) );
  NAND2_X1 u0_u13_u6_U58 (.ZN( u0_u13_u6_n122 ) , .A1( u0_u13_u6_n94 ) , .A2( u0_u13_u6_n97 ) );
  INV_X1 u0_u13_u6_U59 (.A( u0_u13_u6_n139 ) , .ZN( u0_u13_u6_n160 ) );
  AOI22_X1 u0_u13_u6_U6 (.B2( u0_u13_u6_n101 ) , .A1( u0_u13_u6_n102 ) , .ZN( u0_u13_u6_n103 ) , .B1( u0_u13_u6_n160 ) , .A2( u0_u13_u6_n161 ) );
  NAND2_X1 u0_u13_u6_U60 (.ZN( u0_u13_u6_n113 ) , .A1( u0_u13_u6_n96 ) , .A2( u0_u13_u6_n98 ) );
  NOR2_X1 u0_u13_u6_U61 (.A2( u0_u13_X_40 ) , .A1( u0_u13_X_41 ) , .ZN( u0_u13_u6_n126 ) );
  NOR2_X1 u0_u13_u6_U62 (.A2( u0_u13_X_39 ) , .A1( u0_u13_X_42 ) , .ZN( u0_u13_u6_n92 ) );
  NOR2_X1 u0_u13_u6_U63 (.A2( u0_u13_X_39 ) , .A1( u0_u13_u6_n156 ) , .ZN( u0_u13_u6_n97 ) );
  NOR2_X1 u0_u13_u6_U64 (.A2( u0_u13_X_38 ) , .A1( u0_u13_u6_n165 ) , .ZN( u0_u13_u6_n95 ) );
  NOR2_X1 u0_u13_u6_U65 (.A2( u0_u13_X_41 ) , .ZN( u0_u13_u6_n111 ) , .A1( u0_u13_u6_n157 ) );
  NOR2_X1 u0_u13_u6_U66 (.A2( u0_u13_X_37 ) , .A1( u0_u13_u6_n162 ) , .ZN( u0_u13_u6_n94 ) );
  NOR2_X1 u0_u13_u6_U67 (.A2( u0_u13_X_37 ) , .A1( u0_u13_X_38 ) , .ZN( u0_u13_u6_n91 ) );
  NAND2_X1 u0_u13_u6_U68 (.A1( u0_u13_X_41 ) , .ZN( u0_u13_u6_n144 ) , .A2( u0_u13_u6_n157 ) );
  NAND2_X1 u0_u13_u6_U69 (.A2( u0_u13_X_40 ) , .A1( u0_u13_X_41 ) , .ZN( u0_u13_u6_n139 ) );
  NOR2_X1 u0_u13_u6_U7 (.A1( u0_u13_u6_n118 ) , .ZN( u0_u13_u6_n143 ) , .A2( u0_u13_u6_n168 ) );
  AND2_X1 u0_u13_u6_U70 (.A1( u0_u13_X_39 ) , .A2( u0_u13_u6_n156 ) , .ZN( u0_u13_u6_n96 ) );
  AND2_X1 u0_u13_u6_U71 (.A1( u0_u13_X_39 ) , .A2( u0_u13_X_42 ) , .ZN( u0_u13_u6_n99 ) );
  INV_X1 u0_u13_u6_U72 (.A( u0_u13_X_40 ) , .ZN( u0_u13_u6_n157 ) );
  INV_X1 u0_u13_u6_U73 (.A( u0_u13_X_37 ) , .ZN( u0_u13_u6_n165 ) );
  INV_X1 u0_u13_u6_U74 (.A( u0_u13_X_38 ) , .ZN( u0_u13_u6_n162 ) );
  INV_X1 u0_u13_u6_U75 (.A( u0_u13_X_42 ) , .ZN( u0_u13_u6_n156 ) );
  NAND4_X1 u0_u13_u6_U76 (.ZN( u0_out13_32 ) , .A4( u0_u13_u6_n103 ) , .A3( u0_u13_u6_n104 ) , .A2( u0_u13_u6_n105 ) , .A1( u0_u13_u6_n106 ) );
  AOI22_X1 u0_u13_u6_U77 (.ZN( u0_u13_u6_n105 ) , .A2( u0_u13_u6_n108 ) , .A1( u0_u13_u6_n118 ) , .B2( u0_u13_u6_n126 ) , .B1( u0_u13_u6_n171 ) );
  AOI22_X1 u0_u13_u6_U78 (.ZN( u0_u13_u6_n104 ) , .A1( u0_u13_u6_n111 ) , .B1( u0_u13_u6_n124 ) , .B2( u0_u13_u6_n151 ) , .A2( u0_u13_u6_n93 ) );
  NAND4_X1 u0_u13_u6_U79 (.ZN( u0_out13_12 ) , .A4( u0_u13_u6_n114 ) , .A3( u0_u13_u6_n115 ) , .A2( u0_u13_u6_n116 ) , .A1( u0_u13_u6_n117 ) );
  OAI21_X1 u0_u13_u6_U8 (.A( u0_u13_u6_n159 ) , .B1( u0_u13_u6_n169 ) , .B2( u0_u13_u6_n173 ) , .ZN( u0_u13_u6_n90 ) );
  OAI22_X1 u0_u13_u6_U80 (.B2( u0_u13_u6_n111 ) , .ZN( u0_u13_u6_n116 ) , .B1( u0_u13_u6_n126 ) , .A2( u0_u13_u6_n164 ) , .A1( u0_u13_u6_n167 ) );
  OAI21_X1 u0_u13_u6_U81 (.A( u0_u13_u6_n108 ) , .ZN( u0_u13_u6_n117 ) , .B2( u0_u13_u6_n141 ) , .B1( u0_u13_u6_n163 ) );
  OAI211_X1 u0_u13_u6_U82 (.ZN( u0_out13_7 ) , .B( u0_u13_u6_n153 ) , .C2( u0_u13_u6_n154 ) , .C1( u0_u13_u6_n155 ) , .A( u0_u13_u6_n174 ) );
  NOR3_X1 u0_u13_u6_U83 (.A1( u0_u13_u6_n141 ) , .ZN( u0_u13_u6_n154 ) , .A3( u0_u13_u6_n164 ) , .A2( u0_u13_u6_n171 ) );
  AOI211_X1 u0_u13_u6_U84 (.B( u0_u13_u6_n149 ) , .A( u0_u13_u6_n150 ) , .C2( u0_u13_u6_n151 ) , .C1( u0_u13_u6_n152 ) , .ZN( u0_u13_u6_n153 ) );
  OAI211_X1 u0_u13_u6_U85 (.ZN( u0_out13_22 ) , .B( u0_u13_u6_n137 ) , .A( u0_u13_u6_n138 ) , .C2( u0_u13_u6_n139 ) , .C1( u0_u13_u6_n140 ) );
  AOI22_X1 u0_u13_u6_U86 (.B1( u0_u13_u6_n124 ) , .A2( u0_u13_u6_n125 ) , .A1( u0_u13_u6_n126 ) , .ZN( u0_u13_u6_n138 ) , .B2( u0_u13_u6_n161 ) );
  AND4_X1 u0_u13_u6_U87 (.A3( u0_u13_u6_n119 ) , .A1( u0_u13_u6_n120 ) , .A4( u0_u13_u6_n129 ) , .ZN( u0_u13_u6_n140 ) , .A2( u0_u13_u6_n143 ) );
  NAND3_X1 u0_u13_u6_U88 (.A2( u0_u13_u6_n123 ) , .ZN( u0_u13_u6_n125 ) , .A1( u0_u13_u6_n130 ) , .A3( u0_u13_u6_n131 ) );
  NAND3_X1 u0_u13_u6_U89 (.A3( u0_u13_u6_n133 ) , .ZN( u0_u13_u6_n141 ) , .A1( u0_u13_u6_n145 ) , .A2( u0_u13_u6_n148 ) );
  INV_X1 u0_u13_u6_U9 (.ZN( u0_u13_u6_n172 ) , .A( u0_u13_u6_n88 ) );
  NAND3_X1 u0_u13_u6_U90 (.ZN( u0_u13_u6_n101 ) , .A3( u0_u13_u6_n107 ) , .A2( u0_u13_u6_n121 ) , .A1( u0_u13_u6_n127 ) );
  NAND3_X1 u0_u13_u6_U91 (.ZN( u0_u13_u6_n102 ) , .A3( u0_u13_u6_n130 ) , .A2( u0_u13_u6_n145 ) , .A1( u0_u13_u6_n166 ) );
  NAND3_X1 u0_u13_u6_U92 (.A3( u0_u13_u6_n113 ) , .A1( u0_u13_u6_n119 ) , .A2( u0_u13_u6_n123 ) , .ZN( u0_u13_u6_n93 ) );
  NAND3_X1 u0_u13_u6_U93 (.ZN( u0_u13_u6_n142 ) , .A2( u0_u13_u6_n172 ) , .A3( u0_u13_u6_n89 ) , .A1( u0_u13_u6_n90 ) );
  XOR2_X1 u0_u14_U10 (.B( u0_K15_45 ) , .A( u0_R13_30 ) , .Z( u0_u14_X_45 ) );
  XOR2_X1 u0_u14_U11 (.B( u0_K15_44 ) , .A( u0_R13_29 ) , .Z( u0_u14_X_44 ) );
  XOR2_X1 u0_u14_U12 (.B( u0_K15_43 ) , .A( u0_R13_28 ) , .Z( u0_u14_X_43 ) );
  XOR2_X1 u0_u14_U13 (.B( u0_K15_42 ) , .A( u0_R13_29 ) , .Z( u0_u14_X_42 ) );
  XOR2_X1 u0_u14_U14 (.B( u0_K15_41 ) , .A( u0_R13_28 ) , .Z( u0_u14_X_41 ) );
  XOR2_X1 u0_u14_U15 (.B( u0_K15_40 ) , .A( u0_R13_27 ) , .Z( u0_u14_X_40 ) );
  XOR2_X1 u0_u14_U17 (.B( u0_K15_39 ) , .A( u0_R13_26 ) , .Z( u0_u14_X_39 ) );
  XOR2_X1 u0_u14_U18 (.B( u0_K15_38 ) , .A( u0_R13_25 ) , .Z( u0_u14_X_38 ) );
  XOR2_X1 u0_u14_U19 (.B( u0_K15_37 ) , .A( u0_R13_24 ) , .Z( u0_u14_X_37 ) );
  XOR2_X1 u0_u14_U20 (.B( u0_K15_36 ) , .A( u0_R13_25 ) , .Z( u0_u14_X_36 ) );
  XOR2_X1 u0_u14_U21 (.B( u0_K15_35 ) , .A( u0_R13_24 ) , .Z( u0_u14_X_35 ) );
  XOR2_X1 u0_u14_U22 (.B( u0_K15_34 ) , .A( u0_R13_23 ) , .Z( u0_u14_X_34 ) );
  XOR2_X1 u0_u14_U23 (.B( u0_K15_33 ) , .A( u0_R13_22 ) , .Z( u0_u14_X_33 ) );
  XOR2_X1 u0_u14_U24 (.B( u0_K15_32 ) , .A( u0_R13_21 ) , .Z( u0_u14_X_32 ) );
  XOR2_X1 u0_u14_U25 (.B( u0_K15_31 ) , .A( u0_R13_20 ) , .Z( u0_u14_X_31 ) );
  XOR2_X1 u0_u14_U26 (.B( u0_K15_30 ) , .A( u0_R13_21 ) , .Z( u0_u14_X_30 ) );
  XOR2_X1 u0_u14_U28 (.B( u0_K15_29 ) , .A( u0_R13_20 ) , .Z( u0_u14_X_29 ) );
  XOR2_X1 u0_u14_U29 (.B( u0_K15_28 ) , .A( u0_R13_19 ) , .Z( u0_u14_X_28 ) );
  XOR2_X1 u0_u14_U30 (.B( u0_K15_27 ) , .A( u0_R13_18 ) , .Z( u0_u14_X_27 ) );
  XOR2_X1 u0_u14_U31 (.B( u0_K15_26 ) , .A( u0_R13_17 ) , .Z( u0_u14_X_26 ) );
  XOR2_X1 u0_u14_U9 (.B( u0_K15_46 ) , .A( u0_R13_31 ) , .Z( u0_u14_X_46 ) );
  OAI22_X1 u0_u14_u4_U10 (.B2( u0_u14_u4_n135 ) , .ZN( u0_u14_u4_n137 ) , .B1( u0_u14_u4_n153 ) , .A1( u0_u14_u4_n155 ) , .A2( u0_u14_u4_n171 ) );
  AND3_X1 u0_u14_u4_U11 (.A2( u0_u14_u4_n134 ) , .ZN( u0_u14_u4_n135 ) , .A3( u0_u14_u4_n145 ) , .A1( u0_u14_u4_n157 ) );
  NAND2_X1 u0_u14_u4_U12 (.ZN( u0_u14_u4_n132 ) , .A2( u0_u14_u4_n170 ) , .A1( u0_u14_u4_n173 ) );
  AOI21_X1 u0_u14_u4_U13 (.B2( u0_u14_u4_n160 ) , .B1( u0_u14_u4_n161 ) , .ZN( u0_u14_u4_n162 ) , .A( u0_u14_u4_n170 ) );
  AOI21_X1 u0_u14_u4_U14 (.ZN( u0_u14_u4_n107 ) , .B2( u0_u14_u4_n143 ) , .A( u0_u14_u4_n174 ) , .B1( u0_u14_u4_n184 ) );
  AOI21_X1 u0_u14_u4_U15 (.B2( u0_u14_u4_n158 ) , .B1( u0_u14_u4_n159 ) , .ZN( u0_u14_u4_n163 ) , .A( u0_u14_u4_n174 ) );
  AOI21_X1 u0_u14_u4_U16 (.A( u0_u14_u4_n153 ) , .B2( u0_u14_u4_n154 ) , .B1( u0_u14_u4_n155 ) , .ZN( u0_u14_u4_n165 ) );
  AOI21_X1 u0_u14_u4_U17 (.A( u0_u14_u4_n156 ) , .B2( u0_u14_u4_n157 ) , .ZN( u0_u14_u4_n164 ) , .B1( u0_u14_u4_n184 ) );
  INV_X1 u0_u14_u4_U18 (.A( u0_u14_u4_n138 ) , .ZN( u0_u14_u4_n170 ) );
  AND2_X1 u0_u14_u4_U19 (.A2( u0_u14_u4_n120 ) , .ZN( u0_u14_u4_n155 ) , .A1( u0_u14_u4_n160 ) );
  INV_X1 u0_u14_u4_U20 (.A( u0_u14_u4_n156 ) , .ZN( u0_u14_u4_n175 ) );
  NAND2_X1 u0_u14_u4_U21 (.A2( u0_u14_u4_n118 ) , .ZN( u0_u14_u4_n131 ) , .A1( u0_u14_u4_n147 ) );
  NAND2_X1 u0_u14_u4_U22 (.A1( u0_u14_u4_n119 ) , .A2( u0_u14_u4_n120 ) , .ZN( u0_u14_u4_n130 ) );
  NAND2_X1 u0_u14_u4_U23 (.ZN( u0_u14_u4_n117 ) , .A2( u0_u14_u4_n118 ) , .A1( u0_u14_u4_n148 ) );
  NAND2_X1 u0_u14_u4_U24 (.ZN( u0_u14_u4_n129 ) , .A1( u0_u14_u4_n134 ) , .A2( u0_u14_u4_n148 ) );
  AND3_X1 u0_u14_u4_U25 (.A1( u0_u14_u4_n119 ) , .A2( u0_u14_u4_n143 ) , .A3( u0_u14_u4_n154 ) , .ZN( u0_u14_u4_n161 ) );
  AND2_X1 u0_u14_u4_U26 (.A1( u0_u14_u4_n145 ) , .A2( u0_u14_u4_n147 ) , .ZN( u0_u14_u4_n159 ) );
  OR3_X1 u0_u14_u4_U27 (.A3( u0_u14_u4_n114 ) , .A2( u0_u14_u4_n115 ) , .A1( u0_u14_u4_n116 ) , .ZN( u0_u14_u4_n136 ) );
  AOI21_X1 u0_u14_u4_U28 (.A( u0_u14_u4_n113 ) , .ZN( u0_u14_u4_n116 ) , .B2( u0_u14_u4_n173 ) , .B1( u0_u14_u4_n174 ) );
  AOI21_X1 u0_u14_u4_U29 (.ZN( u0_u14_u4_n115 ) , .B2( u0_u14_u4_n145 ) , .B1( u0_u14_u4_n146 ) , .A( u0_u14_u4_n156 ) );
  NOR2_X1 u0_u14_u4_U3 (.ZN( u0_u14_u4_n121 ) , .A1( u0_u14_u4_n181 ) , .A2( u0_u14_u4_n182 ) );
  OAI22_X1 u0_u14_u4_U30 (.ZN( u0_u14_u4_n114 ) , .A2( u0_u14_u4_n121 ) , .B1( u0_u14_u4_n160 ) , .B2( u0_u14_u4_n170 ) , .A1( u0_u14_u4_n171 ) );
  INV_X1 u0_u14_u4_U31 (.A( u0_u14_u4_n158 ) , .ZN( u0_u14_u4_n182 ) );
  INV_X1 u0_u14_u4_U32 (.ZN( u0_u14_u4_n181 ) , .A( u0_u14_u4_n96 ) );
  INV_X1 u0_u14_u4_U33 (.A( u0_u14_u4_n144 ) , .ZN( u0_u14_u4_n179 ) );
  INV_X1 u0_u14_u4_U34 (.A( u0_u14_u4_n157 ) , .ZN( u0_u14_u4_n178 ) );
  NAND2_X1 u0_u14_u4_U35 (.A2( u0_u14_u4_n154 ) , .A1( u0_u14_u4_n96 ) , .ZN( u0_u14_u4_n97 ) );
  INV_X1 u0_u14_u4_U36 (.ZN( u0_u14_u4_n186 ) , .A( u0_u14_u4_n95 ) );
  OAI221_X1 u0_u14_u4_U37 (.C1( u0_u14_u4_n134 ) , .B1( u0_u14_u4_n158 ) , .B2( u0_u14_u4_n171 ) , .C2( u0_u14_u4_n173 ) , .A( u0_u14_u4_n94 ) , .ZN( u0_u14_u4_n95 ) );
  AOI222_X1 u0_u14_u4_U38 (.B2( u0_u14_u4_n132 ) , .A1( u0_u14_u4_n138 ) , .C2( u0_u14_u4_n175 ) , .A2( u0_u14_u4_n179 ) , .C1( u0_u14_u4_n181 ) , .B1( u0_u14_u4_n185 ) , .ZN( u0_u14_u4_n94 ) );
  INV_X1 u0_u14_u4_U39 (.A( u0_u14_u4_n113 ) , .ZN( u0_u14_u4_n185 ) );
  INV_X1 u0_u14_u4_U4 (.A( u0_u14_u4_n117 ) , .ZN( u0_u14_u4_n184 ) );
  INV_X1 u0_u14_u4_U40 (.A( u0_u14_u4_n143 ) , .ZN( u0_u14_u4_n183 ) );
  NOR2_X1 u0_u14_u4_U41 (.ZN( u0_u14_u4_n138 ) , .A1( u0_u14_u4_n168 ) , .A2( u0_u14_u4_n169 ) );
  NOR2_X1 u0_u14_u4_U42 (.A1( u0_u14_u4_n150 ) , .A2( u0_u14_u4_n152 ) , .ZN( u0_u14_u4_n153 ) );
  NOR2_X1 u0_u14_u4_U43 (.A2( u0_u14_u4_n128 ) , .A1( u0_u14_u4_n138 ) , .ZN( u0_u14_u4_n156 ) );
  AOI22_X1 u0_u14_u4_U44 (.B2( u0_u14_u4_n122 ) , .A1( u0_u14_u4_n123 ) , .ZN( u0_u14_u4_n124 ) , .B1( u0_u14_u4_n128 ) , .A2( u0_u14_u4_n172 ) );
  INV_X1 u0_u14_u4_U45 (.A( u0_u14_u4_n153 ) , .ZN( u0_u14_u4_n172 ) );
  NAND2_X1 u0_u14_u4_U46 (.A2( u0_u14_u4_n120 ) , .ZN( u0_u14_u4_n123 ) , .A1( u0_u14_u4_n161 ) );
  AOI22_X1 u0_u14_u4_U47 (.B2( u0_u14_u4_n132 ) , .A2( u0_u14_u4_n133 ) , .ZN( u0_u14_u4_n140 ) , .A1( u0_u14_u4_n150 ) , .B1( u0_u14_u4_n179 ) );
  NAND2_X1 u0_u14_u4_U48 (.ZN( u0_u14_u4_n133 ) , .A2( u0_u14_u4_n146 ) , .A1( u0_u14_u4_n154 ) );
  NAND2_X1 u0_u14_u4_U49 (.A1( u0_u14_u4_n103 ) , .ZN( u0_u14_u4_n154 ) , .A2( u0_u14_u4_n98 ) );
  NOR4_X1 u0_u14_u4_U5 (.A4( u0_u14_u4_n106 ) , .A3( u0_u14_u4_n107 ) , .A2( u0_u14_u4_n108 ) , .A1( u0_u14_u4_n109 ) , .ZN( u0_u14_u4_n110 ) );
  NAND2_X1 u0_u14_u4_U50 (.A1( u0_u14_u4_n101 ) , .ZN( u0_u14_u4_n158 ) , .A2( u0_u14_u4_n99 ) );
  AOI21_X1 u0_u14_u4_U51 (.ZN( u0_u14_u4_n127 ) , .A( u0_u14_u4_n136 ) , .B2( u0_u14_u4_n150 ) , .B1( u0_u14_u4_n180 ) );
  INV_X1 u0_u14_u4_U52 (.A( u0_u14_u4_n160 ) , .ZN( u0_u14_u4_n180 ) );
  NAND2_X1 u0_u14_u4_U53 (.A2( u0_u14_u4_n104 ) , .A1( u0_u14_u4_n105 ) , .ZN( u0_u14_u4_n146 ) );
  NAND2_X1 u0_u14_u4_U54 (.A2( u0_u14_u4_n101 ) , .A1( u0_u14_u4_n102 ) , .ZN( u0_u14_u4_n160 ) );
  NAND2_X1 u0_u14_u4_U55 (.ZN( u0_u14_u4_n134 ) , .A1( u0_u14_u4_n98 ) , .A2( u0_u14_u4_n99 ) );
  NAND2_X1 u0_u14_u4_U56 (.A1( u0_u14_u4_n103 ) , .A2( u0_u14_u4_n104 ) , .ZN( u0_u14_u4_n143 ) );
  NAND2_X1 u0_u14_u4_U57 (.A2( u0_u14_u4_n105 ) , .ZN( u0_u14_u4_n145 ) , .A1( u0_u14_u4_n98 ) );
  NAND2_X1 u0_u14_u4_U58 (.A1( u0_u14_u4_n100 ) , .A2( u0_u14_u4_n105 ) , .ZN( u0_u14_u4_n120 ) );
  NAND2_X1 u0_u14_u4_U59 (.A1( u0_u14_u4_n102 ) , .A2( u0_u14_u4_n104 ) , .ZN( u0_u14_u4_n148 ) );
  AOI21_X1 u0_u14_u4_U6 (.ZN( u0_u14_u4_n106 ) , .B2( u0_u14_u4_n146 ) , .B1( u0_u14_u4_n158 ) , .A( u0_u14_u4_n170 ) );
  NAND2_X1 u0_u14_u4_U60 (.A2( u0_u14_u4_n100 ) , .A1( u0_u14_u4_n103 ) , .ZN( u0_u14_u4_n157 ) );
  INV_X1 u0_u14_u4_U61 (.A( u0_u14_u4_n150 ) , .ZN( u0_u14_u4_n173 ) );
  INV_X1 u0_u14_u4_U62 (.A( u0_u14_u4_n152 ) , .ZN( u0_u14_u4_n171 ) );
  NAND2_X1 u0_u14_u4_U63 (.A1( u0_u14_u4_n100 ) , .ZN( u0_u14_u4_n118 ) , .A2( u0_u14_u4_n99 ) );
  NAND2_X1 u0_u14_u4_U64 (.A2( u0_u14_u4_n100 ) , .A1( u0_u14_u4_n102 ) , .ZN( u0_u14_u4_n144 ) );
  NAND2_X1 u0_u14_u4_U65 (.A2( u0_u14_u4_n101 ) , .A1( u0_u14_u4_n105 ) , .ZN( u0_u14_u4_n96 ) );
  INV_X1 u0_u14_u4_U66 (.A( u0_u14_u4_n128 ) , .ZN( u0_u14_u4_n174 ) );
  NAND2_X1 u0_u14_u4_U67 (.A2( u0_u14_u4_n102 ) , .ZN( u0_u14_u4_n119 ) , .A1( u0_u14_u4_n98 ) );
  NAND2_X1 u0_u14_u4_U68 (.A2( u0_u14_u4_n101 ) , .A1( u0_u14_u4_n103 ) , .ZN( u0_u14_u4_n147 ) );
  NAND2_X1 u0_u14_u4_U69 (.A2( u0_u14_u4_n104 ) , .ZN( u0_u14_u4_n113 ) , .A1( u0_u14_u4_n99 ) );
  AOI21_X1 u0_u14_u4_U7 (.ZN( u0_u14_u4_n108 ) , .B2( u0_u14_u4_n134 ) , .B1( u0_u14_u4_n155 ) , .A( u0_u14_u4_n156 ) );
  NOR2_X1 u0_u14_u4_U70 (.A2( u0_u14_X_28 ) , .ZN( u0_u14_u4_n150 ) , .A1( u0_u14_u4_n168 ) );
  NOR2_X1 u0_u14_u4_U71 (.A2( u0_u14_X_29 ) , .ZN( u0_u14_u4_n152 ) , .A1( u0_u14_u4_n169 ) );
  NOR2_X1 u0_u14_u4_U72 (.A2( u0_u14_X_30 ) , .ZN( u0_u14_u4_n105 ) , .A1( u0_u14_u4_n176 ) );
  NOR2_X1 u0_u14_u4_U73 (.A2( u0_u14_X_26 ) , .ZN( u0_u14_u4_n100 ) , .A1( u0_u14_u4_n177 ) );
  NOR2_X1 u0_u14_u4_U74 (.A2( u0_u14_X_28 ) , .A1( u0_u14_X_29 ) , .ZN( u0_u14_u4_n128 ) );
  NOR2_X1 u0_u14_u4_U75 (.A2( u0_u14_X_27 ) , .A1( u0_u14_X_30 ) , .ZN( u0_u14_u4_n102 ) );
  NOR2_X1 u0_u14_u4_U76 (.A2( u0_u14_X_25 ) , .A1( u0_u14_X_26 ) , .ZN( u0_u14_u4_n98 ) );
  AND2_X1 u0_u14_u4_U77 (.A2( u0_u14_X_25 ) , .A1( u0_u14_X_26 ) , .ZN( u0_u14_u4_n104 ) );
  AND2_X1 u0_u14_u4_U78 (.A1( u0_u14_X_30 ) , .A2( u0_u14_u4_n176 ) , .ZN( u0_u14_u4_n99 ) );
  AND2_X1 u0_u14_u4_U79 (.A1( u0_u14_X_26 ) , .ZN( u0_u14_u4_n101 ) , .A2( u0_u14_u4_n177 ) );
  AOI21_X1 u0_u14_u4_U8 (.ZN( u0_u14_u4_n109 ) , .A( u0_u14_u4_n153 ) , .B1( u0_u14_u4_n159 ) , .B2( u0_u14_u4_n184 ) );
  AND2_X1 u0_u14_u4_U80 (.A1( u0_u14_X_27 ) , .A2( u0_u14_X_30 ) , .ZN( u0_u14_u4_n103 ) );
  INV_X1 u0_u14_u4_U81 (.A( u0_u14_X_28 ) , .ZN( u0_u14_u4_n169 ) );
  INV_X1 u0_u14_u4_U82 (.A( u0_u14_X_29 ) , .ZN( u0_u14_u4_n168 ) );
  INV_X1 u0_u14_u4_U83 (.A( u0_u14_X_25 ) , .ZN( u0_u14_u4_n177 ) );
  INV_X1 u0_u14_u4_U84 (.A( u0_u14_X_27 ) , .ZN( u0_u14_u4_n176 ) );
  NAND4_X1 u0_u14_u4_U85 (.ZN( u0_out14_25 ) , .A4( u0_u14_u4_n139 ) , .A3( u0_u14_u4_n140 ) , .A2( u0_u14_u4_n141 ) , .A1( u0_u14_u4_n142 ) );
  OAI21_X1 u0_u14_u4_U86 (.A( u0_u14_u4_n128 ) , .B2( u0_u14_u4_n129 ) , .B1( u0_u14_u4_n130 ) , .ZN( u0_u14_u4_n142 ) );
  OAI21_X1 u0_u14_u4_U87 (.B2( u0_u14_u4_n131 ) , .ZN( u0_u14_u4_n141 ) , .A( u0_u14_u4_n175 ) , .B1( u0_u14_u4_n183 ) );
  NAND4_X1 u0_u14_u4_U88 (.ZN( u0_out14_14 ) , .A4( u0_u14_u4_n124 ) , .A3( u0_u14_u4_n125 ) , .A2( u0_u14_u4_n126 ) , .A1( u0_u14_u4_n127 ) );
  AOI22_X1 u0_u14_u4_U89 (.B2( u0_u14_u4_n117 ) , .ZN( u0_u14_u4_n126 ) , .A1( u0_u14_u4_n129 ) , .B1( u0_u14_u4_n152 ) , .A2( u0_u14_u4_n175 ) );
  AOI211_X1 u0_u14_u4_U9 (.B( u0_u14_u4_n136 ) , .A( u0_u14_u4_n137 ) , .C2( u0_u14_u4_n138 ) , .ZN( u0_u14_u4_n139 ) , .C1( u0_u14_u4_n182 ) );
  AOI22_X1 u0_u14_u4_U90 (.ZN( u0_u14_u4_n125 ) , .B2( u0_u14_u4_n131 ) , .A2( u0_u14_u4_n132 ) , .B1( u0_u14_u4_n138 ) , .A1( u0_u14_u4_n178 ) );
  NAND4_X1 u0_u14_u4_U91 (.ZN( u0_out14_8 ) , .A4( u0_u14_u4_n110 ) , .A3( u0_u14_u4_n111 ) , .A2( u0_u14_u4_n112 ) , .A1( u0_u14_u4_n186 ) );
  NAND2_X1 u0_u14_u4_U92 (.ZN( u0_u14_u4_n112 ) , .A2( u0_u14_u4_n130 ) , .A1( u0_u14_u4_n150 ) );
  AOI22_X1 u0_u14_u4_U93 (.ZN( u0_u14_u4_n111 ) , .B2( u0_u14_u4_n132 ) , .A1( u0_u14_u4_n152 ) , .B1( u0_u14_u4_n178 ) , .A2( u0_u14_u4_n97 ) );
  AOI22_X1 u0_u14_u4_U94 (.B2( u0_u14_u4_n149 ) , .B1( u0_u14_u4_n150 ) , .A2( u0_u14_u4_n151 ) , .A1( u0_u14_u4_n152 ) , .ZN( u0_u14_u4_n167 ) );
  NOR4_X1 u0_u14_u4_U95 (.A4( u0_u14_u4_n162 ) , .A3( u0_u14_u4_n163 ) , .A2( u0_u14_u4_n164 ) , .A1( u0_u14_u4_n165 ) , .ZN( u0_u14_u4_n166 ) );
  NAND3_X1 u0_u14_u4_U96 (.ZN( u0_out14_3 ) , .A3( u0_u14_u4_n166 ) , .A1( u0_u14_u4_n167 ) , .A2( u0_u14_u4_n186 ) );
  NAND3_X1 u0_u14_u4_U97 (.A3( u0_u14_u4_n146 ) , .A2( u0_u14_u4_n147 ) , .A1( u0_u14_u4_n148 ) , .ZN( u0_u14_u4_n149 ) );
  NAND3_X1 u0_u14_u4_U98 (.A3( u0_u14_u4_n143 ) , .A2( u0_u14_u4_n144 ) , .A1( u0_u14_u4_n145 ) , .ZN( u0_u14_u4_n151 ) );
  NAND3_X1 u0_u14_u4_U99 (.A3( u0_u14_u4_n121 ) , .ZN( u0_u14_u4_n122 ) , .A2( u0_u14_u4_n144 ) , .A1( u0_u14_u4_n154 ) );
  INV_X1 u0_u14_u5_U10 (.A( u0_u14_u5_n121 ) , .ZN( u0_u14_u5_n177 ) );
  NOR3_X1 u0_u14_u5_U100 (.A3( u0_u14_u5_n141 ) , .A1( u0_u14_u5_n142 ) , .ZN( u0_u14_u5_n143 ) , .A2( u0_u14_u5_n191 ) );
  NAND4_X1 u0_u14_u5_U101 (.ZN( u0_out14_4 ) , .A4( u0_u14_u5_n112 ) , .A2( u0_u14_u5_n113 ) , .A1( u0_u14_u5_n114 ) , .A3( u0_u14_u5_n195 ) );
  AOI211_X1 u0_u14_u5_U102 (.A( u0_u14_u5_n110 ) , .C1( u0_u14_u5_n111 ) , .ZN( u0_u14_u5_n112 ) , .B( u0_u14_u5_n118 ) , .C2( u0_u14_u5_n177 ) );
  AOI222_X1 u0_u14_u5_U103 (.ZN( u0_u14_u5_n113 ) , .A1( u0_u14_u5_n131 ) , .C1( u0_u14_u5_n148 ) , .B2( u0_u14_u5_n174 ) , .C2( u0_u14_u5_n178 ) , .A2( u0_u14_u5_n179 ) , .B1( u0_u14_u5_n99 ) );
  NAND3_X1 u0_u14_u5_U104 (.A2( u0_u14_u5_n154 ) , .A3( u0_u14_u5_n158 ) , .A1( u0_u14_u5_n161 ) , .ZN( u0_u14_u5_n99 ) );
  NOR2_X1 u0_u14_u5_U11 (.ZN( u0_u14_u5_n160 ) , .A2( u0_u14_u5_n173 ) , .A1( u0_u14_u5_n177 ) );
  INV_X1 u0_u14_u5_U12 (.A( u0_u14_u5_n150 ) , .ZN( u0_u14_u5_n174 ) );
  AOI21_X1 u0_u14_u5_U13 (.A( u0_u14_u5_n160 ) , .B2( u0_u14_u5_n161 ) , .ZN( u0_u14_u5_n162 ) , .B1( u0_u14_u5_n192 ) );
  INV_X1 u0_u14_u5_U14 (.A( u0_u14_u5_n159 ) , .ZN( u0_u14_u5_n192 ) );
  AOI21_X1 u0_u14_u5_U15 (.A( u0_u14_u5_n156 ) , .B2( u0_u14_u5_n157 ) , .B1( u0_u14_u5_n158 ) , .ZN( u0_u14_u5_n163 ) );
  AOI21_X1 u0_u14_u5_U16 (.B2( u0_u14_u5_n139 ) , .B1( u0_u14_u5_n140 ) , .ZN( u0_u14_u5_n141 ) , .A( u0_u14_u5_n150 ) );
  OAI21_X1 u0_u14_u5_U17 (.A( u0_u14_u5_n133 ) , .B2( u0_u14_u5_n134 ) , .B1( u0_u14_u5_n135 ) , .ZN( u0_u14_u5_n142 ) );
  OAI21_X1 u0_u14_u5_U18 (.ZN( u0_u14_u5_n133 ) , .B2( u0_u14_u5_n147 ) , .A( u0_u14_u5_n173 ) , .B1( u0_u14_u5_n188 ) );
  NAND2_X1 u0_u14_u5_U19 (.A2( u0_u14_u5_n119 ) , .A1( u0_u14_u5_n123 ) , .ZN( u0_u14_u5_n137 ) );
  INV_X1 u0_u14_u5_U20 (.A( u0_u14_u5_n155 ) , .ZN( u0_u14_u5_n194 ) );
  NAND2_X1 u0_u14_u5_U21 (.A1( u0_u14_u5_n121 ) , .ZN( u0_u14_u5_n132 ) , .A2( u0_u14_u5_n172 ) );
  NAND2_X1 u0_u14_u5_U22 (.A2( u0_u14_u5_n122 ) , .ZN( u0_u14_u5_n136 ) , .A1( u0_u14_u5_n154 ) );
  NAND2_X1 u0_u14_u5_U23 (.A2( u0_u14_u5_n119 ) , .A1( u0_u14_u5_n120 ) , .ZN( u0_u14_u5_n159 ) );
  INV_X1 u0_u14_u5_U24 (.A( u0_u14_u5_n156 ) , .ZN( u0_u14_u5_n175 ) );
  INV_X1 u0_u14_u5_U25 (.A( u0_u14_u5_n158 ) , .ZN( u0_u14_u5_n188 ) );
  INV_X1 u0_u14_u5_U26 (.A( u0_u14_u5_n152 ) , .ZN( u0_u14_u5_n179 ) );
  INV_X1 u0_u14_u5_U27 (.A( u0_u14_u5_n140 ) , .ZN( u0_u14_u5_n182 ) );
  INV_X1 u0_u14_u5_U28 (.A( u0_u14_u5_n151 ) , .ZN( u0_u14_u5_n183 ) );
  INV_X1 u0_u14_u5_U29 (.A( u0_u14_u5_n123 ) , .ZN( u0_u14_u5_n185 ) );
  NOR2_X1 u0_u14_u5_U3 (.ZN( u0_u14_u5_n134 ) , .A1( u0_u14_u5_n183 ) , .A2( u0_u14_u5_n190 ) );
  INV_X1 u0_u14_u5_U30 (.A( u0_u14_u5_n161 ) , .ZN( u0_u14_u5_n184 ) );
  INV_X1 u0_u14_u5_U31 (.A( u0_u14_u5_n139 ) , .ZN( u0_u14_u5_n189 ) );
  INV_X1 u0_u14_u5_U32 (.A( u0_u14_u5_n157 ) , .ZN( u0_u14_u5_n190 ) );
  INV_X1 u0_u14_u5_U33 (.A( u0_u14_u5_n120 ) , .ZN( u0_u14_u5_n193 ) );
  NAND2_X1 u0_u14_u5_U34 (.ZN( u0_u14_u5_n111 ) , .A1( u0_u14_u5_n140 ) , .A2( u0_u14_u5_n155 ) );
  INV_X1 u0_u14_u5_U35 (.A( u0_u14_u5_n117 ) , .ZN( u0_u14_u5_n196 ) );
  OAI221_X1 u0_u14_u5_U36 (.A( u0_u14_u5_n116 ) , .ZN( u0_u14_u5_n117 ) , .B2( u0_u14_u5_n119 ) , .C1( u0_u14_u5_n153 ) , .C2( u0_u14_u5_n158 ) , .B1( u0_u14_u5_n172 ) );
  AOI222_X1 u0_u14_u5_U37 (.ZN( u0_u14_u5_n116 ) , .B2( u0_u14_u5_n145 ) , .C1( u0_u14_u5_n148 ) , .A2( u0_u14_u5_n174 ) , .C2( u0_u14_u5_n177 ) , .B1( u0_u14_u5_n187 ) , .A1( u0_u14_u5_n193 ) );
  INV_X1 u0_u14_u5_U38 (.A( u0_u14_u5_n115 ) , .ZN( u0_u14_u5_n187 ) );
  NOR2_X1 u0_u14_u5_U39 (.ZN( u0_u14_u5_n100 ) , .A1( u0_u14_u5_n170 ) , .A2( u0_u14_u5_n180 ) );
  INV_X1 u0_u14_u5_U4 (.A( u0_u14_u5_n138 ) , .ZN( u0_u14_u5_n191 ) );
  AOI22_X1 u0_u14_u5_U40 (.B2( u0_u14_u5_n131 ) , .A2( u0_u14_u5_n146 ) , .ZN( u0_u14_u5_n169 ) , .B1( u0_u14_u5_n174 ) , .A1( u0_u14_u5_n185 ) );
  NOR2_X1 u0_u14_u5_U41 (.A1( u0_u14_u5_n146 ) , .ZN( u0_u14_u5_n150 ) , .A2( u0_u14_u5_n173 ) );
  AOI21_X1 u0_u14_u5_U42 (.A( u0_u14_u5_n118 ) , .B2( u0_u14_u5_n145 ) , .ZN( u0_u14_u5_n168 ) , .B1( u0_u14_u5_n186 ) );
  INV_X1 u0_u14_u5_U43 (.A( u0_u14_u5_n122 ) , .ZN( u0_u14_u5_n186 ) );
  NOR2_X1 u0_u14_u5_U44 (.A1( u0_u14_u5_n146 ) , .ZN( u0_u14_u5_n152 ) , .A2( u0_u14_u5_n176 ) );
  NOR2_X1 u0_u14_u5_U45 (.A1( u0_u14_u5_n115 ) , .ZN( u0_u14_u5_n118 ) , .A2( u0_u14_u5_n153 ) );
  NOR2_X1 u0_u14_u5_U46 (.A2( u0_u14_u5_n145 ) , .ZN( u0_u14_u5_n156 ) , .A1( u0_u14_u5_n174 ) );
  NOR2_X1 u0_u14_u5_U47 (.ZN( u0_u14_u5_n121 ) , .A2( u0_u14_u5_n145 ) , .A1( u0_u14_u5_n176 ) );
  AOI22_X1 u0_u14_u5_U48 (.ZN( u0_u14_u5_n114 ) , .A2( u0_u14_u5_n137 ) , .A1( u0_u14_u5_n145 ) , .B2( u0_u14_u5_n175 ) , .B1( u0_u14_u5_n193 ) );
  OAI211_X1 u0_u14_u5_U49 (.B( u0_u14_u5_n124 ) , .A( u0_u14_u5_n125 ) , .C2( u0_u14_u5_n126 ) , .C1( u0_u14_u5_n127 ) , .ZN( u0_u14_u5_n128 ) );
  OAI21_X1 u0_u14_u5_U5 (.B2( u0_u14_u5_n136 ) , .B1( u0_u14_u5_n137 ) , .ZN( u0_u14_u5_n138 ) , .A( u0_u14_u5_n177 ) );
  NOR3_X1 u0_u14_u5_U50 (.ZN( u0_u14_u5_n127 ) , .A1( u0_u14_u5_n136 ) , .A3( u0_u14_u5_n148 ) , .A2( u0_u14_u5_n182 ) );
  OAI21_X1 u0_u14_u5_U51 (.ZN( u0_u14_u5_n124 ) , .A( u0_u14_u5_n177 ) , .B2( u0_u14_u5_n183 ) , .B1( u0_u14_u5_n189 ) );
  OAI21_X1 u0_u14_u5_U52 (.ZN( u0_u14_u5_n125 ) , .A( u0_u14_u5_n174 ) , .B2( u0_u14_u5_n185 ) , .B1( u0_u14_u5_n190 ) );
  AOI21_X1 u0_u14_u5_U53 (.A( u0_u14_u5_n153 ) , .B2( u0_u14_u5_n154 ) , .B1( u0_u14_u5_n155 ) , .ZN( u0_u14_u5_n164 ) );
  AOI21_X1 u0_u14_u5_U54 (.ZN( u0_u14_u5_n110 ) , .B1( u0_u14_u5_n122 ) , .B2( u0_u14_u5_n139 ) , .A( u0_u14_u5_n153 ) );
  INV_X1 u0_u14_u5_U55 (.A( u0_u14_u5_n153 ) , .ZN( u0_u14_u5_n176 ) );
  INV_X1 u0_u14_u5_U56 (.A( u0_u14_u5_n126 ) , .ZN( u0_u14_u5_n173 ) );
  AND2_X1 u0_u14_u5_U57 (.A2( u0_u14_u5_n104 ) , .A1( u0_u14_u5_n107 ) , .ZN( u0_u14_u5_n147 ) );
  AND2_X1 u0_u14_u5_U58 (.A2( u0_u14_u5_n104 ) , .A1( u0_u14_u5_n108 ) , .ZN( u0_u14_u5_n148 ) );
  NAND2_X1 u0_u14_u5_U59 (.A1( u0_u14_u5_n105 ) , .A2( u0_u14_u5_n106 ) , .ZN( u0_u14_u5_n158 ) );
  INV_X1 u0_u14_u5_U6 (.A( u0_u14_u5_n135 ) , .ZN( u0_u14_u5_n178 ) );
  NAND2_X1 u0_u14_u5_U60 (.A2( u0_u14_u5_n108 ) , .A1( u0_u14_u5_n109 ) , .ZN( u0_u14_u5_n139 ) );
  NAND2_X1 u0_u14_u5_U61 (.A1( u0_u14_u5_n106 ) , .A2( u0_u14_u5_n108 ) , .ZN( u0_u14_u5_n119 ) );
  NAND2_X1 u0_u14_u5_U62 (.A2( u0_u14_u5_n103 ) , .A1( u0_u14_u5_n105 ) , .ZN( u0_u14_u5_n140 ) );
  NAND2_X1 u0_u14_u5_U63 (.A2( u0_u14_u5_n104 ) , .A1( u0_u14_u5_n105 ) , .ZN( u0_u14_u5_n155 ) );
  NAND2_X1 u0_u14_u5_U64 (.A2( u0_u14_u5_n106 ) , .A1( u0_u14_u5_n107 ) , .ZN( u0_u14_u5_n122 ) );
  NAND2_X1 u0_u14_u5_U65 (.A2( u0_u14_u5_n100 ) , .A1( u0_u14_u5_n106 ) , .ZN( u0_u14_u5_n115 ) );
  NAND2_X1 u0_u14_u5_U66 (.A2( u0_u14_u5_n100 ) , .A1( u0_u14_u5_n103 ) , .ZN( u0_u14_u5_n161 ) );
  NAND2_X1 u0_u14_u5_U67 (.A1( u0_u14_u5_n105 ) , .A2( u0_u14_u5_n109 ) , .ZN( u0_u14_u5_n154 ) );
  INV_X1 u0_u14_u5_U68 (.A( u0_u14_u5_n146 ) , .ZN( u0_u14_u5_n172 ) );
  NAND2_X1 u0_u14_u5_U69 (.A1( u0_u14_u5_n103 ) , .A2( u0_u14_u5_n108 ) , .ZN( u0_u14_u5_n123 ) );
  OAI22_X1 u0_u14_u5_U7 (.B2( u0_u14_u5_n149 ) , .B1( u0_u14_u5_n150 ) , .A2( u0_u14_u5_n151 ) , .A1( u0_u14_u5_n152 ) , .ZN( u0_u14_u5_n165 ) );
  NAND2_X1 u0_u14_u5_U70 (.A2( u0_u14_u5_n103 ) , .A1( u0_u14_u5_n107 ) , .ZN( u0_u14_u5_n151 ) );
  NAND2_X1 u0_u14_u5_U71 (.A2( u0_u14_u5_n107 ) , .A1( u0_u14_u5_n109 ) , .ZN( u0_u14_u5_n120 ) );
  NAND2_X1 u0_u14_u5_U72 (.A2( u0_u14_u5_n100 ) , .A1( u0_u14_u5_n109 ) , .ZN( u0_u14_u5_n157 ) );
  AND2_X1 u0_u14_u5_U73 (.A2( u0_u14_u5_n100 ) , .A1( u0_u14_u5_n104 ) , .ZN( u0_u14_u5_n131 ) );
  INV_X1 u0_u14_u5_U74 (.A( u0_u14_u5_n102 ) , .ZN( u0_u14_u5_n195 ) );
  OAI221_X1 u0_u14_u5_U75 (.A( u0_u14_u5_n101 ) , .ZN( u0_u14_u5_n102 ) , .C2( u0_u14_u5_n115 ) , .C1( u0_u14_u5_n126 ) , .B1( u0_u14_u5_n134 ) , .B2( u0_u14_u5_n160 ) );
  OAI21_X1 u0_u14_u5_U76 (.ZN( u0_u14_u5_n101 ) , .B1( u0_u14_u5_n137 ) , .A( u0_u14_u5_n146 ) , .B2( u0_u14_u5_n147 ) );
  NOR2_X1 u0_u14_u5_U77 (.A2( u0_u14_X_34 ) , .A1( u0_u14_X_35 ) , .ZN( u0_u14_u5_n145 ) );
  NOR2_X1 u0_u14_u5_U78 (.A2( u0_u14_X_34 ) , .ZN( u0_u14_u5_n146 ) , .A1( u0_u14_u5_n171 ) );
  NOR2_X1 u0_u14_u5_U79 (.A2( u0_u14_X_31 ) , .A1( u0_u14_X_32 ) , .ZN( u0_u14_u5_n103 ) );
  NOR3_X1 u0_u14_u5_U8 (.A2( u0_u14_u5_n147 ) , .A1( u0_u14_u5_n148 ) , .ZN( u0_u14_u5_n149 ) , .A3( u0_u14_u5_n194 ) );
  NOR2_X1 u0_u14_u5_U80 (.A2( u0_u14_X_36 ) , .ZN( u0_u14_u5_n105 ) , .A1( u0_u14_u5_n180 ) );
  NOR2_X1 u0_u14_u5_U81 (.A2( u0_u14_X_33 ) , .ZN( u0_u14_u5_n108 ) , .A1( u0_u14_u5_n170 ) );
  NOR2_X1 u0_u14_u5_U82 (.A2( u0_u14_X_33 ) , .A1( u0_u14_X_36 ) , .ZN( u0_u14_u5_n107 ) );
  NOR2_X1 u0_u14_u5_U83 (.A2( u0_u14_X_31 ) , .ZN( u0_u14_u5_n104 ) , .A1( u0_u14_u5_n181 ) );
  NAND2_X1 u0_u14_u5_U84 (.A2( u0_u14_X_34 ) , .A1( u0_u14_X_35 ) , .ZN( u0_u14_u5_n153 ) );
  NAND2_X1 u0_u14_u5_U85 (.A1( u0_u14_X_34 ) , .ZN( u0_u14_u5_n126 ) , .A2( u0_u14_u5_n171 ) );
  AND2_X1 u0_u14_u5_U86 (.A1( u0_u14_X_31 ) , .A2( u0_u14_X_32 ) , .ZN( u0_u14_u5_n106 ) );
  AND2_X1 u0_u14_u5_U87 (.A1( u0_u14_X_31 ) , .ZN( u0_u14_u5_n109 ) , .A2( u0_u14_u5_n181 ) );
  INV_X1 u0_u14_u5_U88 (.A( u0_u14_X_33 ) , .ZN( u0_u14_u5_n180 ) );
  INV_X1 u0_u14_u5_U89 (.A( u0_u14_X_35 ) , .ZN( u0_u14_u5_n171 ) );
  NOR2_X1 u0_u14_u5_U9 (.ZN( u0_u14_u5_n135 ) , .A1( u0_u14_u5_n173 ) , .A2( u0_u14_u5_n176 ) );
  INV_X1 u0_u14_u5_U90 (.A( u0_u14_X_36 ) , .ZN( u0_u14_u5_n170 ) );
  INV_X1 u0_u14_u5_U91 (.A( u0_u14_X_32 ) , .ZN( u0_u14_u5_n181 ) );
  NAND4_X1 u0_u14_u5_U92 (.ZN( u0_out14_29 ) , .A4( u0_u14_u5_n129 ) , .A3( u0_u14_u5_n130 ) , .A2( u0_u14_u5_n168 ) , .A1( u0_u14_u5_n196 ) );
  AOI221_X1 u0_u14_u5_U93 (.A( u0_u14_u5_n128 ) , .ZN( u0_u14_u5_n129 ) , .C2( u0_u14_u5_n132 ) , .B2( u0_u14_u5_n159 ) , .B1( u0_u14_u5_n176 ) , .C1( u0_u14_u5_n184 ) );
  AOI222_X1 u0_u14_u5_U94 (.ZN( u0_u14_u5_n130 ) , .A2( u0_u14_u5_n146 ) , .B1( u0_u14_u5_n147 ) , .C2( u0_u14_u5_n175 ) , .B2( u0_u14_u5_n179 ) , .A1( u0_u14_u5_n188 ) , .C1( u0_u14_u5_n194 ) );
  NAND4_X1 u0_u14_u5_U95 (.ZN( u0_out14_19 ) , .A4( u0_u14_u5_n166 ) , .A3( u0_u14_u5_n167 ) , .A2( u0_u14_u5_n168 ) , .A1( u0_u14_u5_n169 ) );
  AOI22_X1 u0_u14_u5_U96 (.B2( u0_u14_u5_n145 ) , .A2( u0_u14_u5_n146 ) , .ZN( u0_u14_u5_n167 ) , .B1( u0_u14_u5_n182 ) , .A1( u0_u14_u5_n189 ) );
  NOR4_X1 u0_u14_u5_U97 (.A4( u0_u14_u5_n162 ) , .A3( u0_u14_u5_n163 ) , .A2( u0_u14_u5_n164 ) , .A1( u0_u14_u5_n165 ) , .ZN( u0_u14_u5_n166 ) );
  NAND4_X1 u0_u14_u5_U98 (.ZN( u0_out14_11 ) , .A4( u0_u14_u5_n143 ) , .A3( u0_u14_u5_n144 ) , .A2( u0_u14_u5_n169 ) , .A1( u0_u14_u5_n196 ) );
  AOI22_X1 u0_u14_u5_U99 (.A2( u0_u14_u5_n132 ) , .ZN( u0_u14_u5_n144 ) , .B2( u0_u14_u5_n145 ) , .B1( u0_u14_u5_n184 ) , .A1( u0_u14_u5_n194 ) );
  AOI21_X1 u0_u14_u6_U10 (.ZN( u0_u14_u6_n106 ) , .A( u0_u14_u6_n142 ) , .B2( u0_u14_u6_n159 ) , .B1( u0_u14_u6_n164 ) );
  INV_X1 u0_u14_u6_U11 (.A( u0_u14_u6_n155 ) , .ZN( u0_u14_u6_n161 ) );
  INV_X1 u0_u14_u6_U12 (.A( u0_u14_u6_n128 ) , .ZN( u0_u14_u6_n164 ) );
  NAND2_X1 u0_u14_u6_U13 (.ZN( u0_u14_u6_n110 ) , .A1( u0_u14_u6_n122 ) , .A2( u0_u14_u6_n129 ) );
  NAND2_X1 u0_u14_u6_U14 (.ZN( u0_u14_u6_n124 ) , .A2( u0_u14_u6_n146 ) , .A1( u0_u14_u6_n148 ) );
  INV_X1 u0_u14_u6_U15 (.A( u0_u14_u6_n132 ) , .ZN( u0_u14_u6_n171 ) );
  AND2_X1 u0_u14_u6_U16 (.A1( u0_u14_u6_n100 ) , .ZN( u0_u14_u6_n130 ) , .A2( u0_u14_u6_n147 ) );
  INV_X1 u0_u14_u6_U17 (.A( u0_u14_u6_n127 ) , .ZN( u0_u14_u6_n173 ) );
  INV_X1 u0_u14_u6_U18 (.A( u0_u14_u6_n121 ) , .ZN( u0_u14_u6_n167 ) );
  INV_X1 u0_u14_u6_U19 (.A( u0_u14_u6_n100 ) , .ZN( u0_u14_u6_n169 ) );
  INV_X1 u0_u14_u6_U20 (.A( u0_u14_u6_n123 ) , .ZN( u0_u14_u6_n170 ) );
  INV_X1 u0_u14_u6_U21 (.A( u0_u14_u6_n113 ) , .ZN( u0_u14_u6_n168 ) );
  AND2_X1 u0_u14_u6_U22 (.A1( u0_u14_u6_n107 ) , .A2( u0_u14_u6_n119 ) , .ZN( u0_u14_u6_n133 ) );
  AND2_X1 u0_u14_u6_U23 (.A2( u0_u14_u6_n121 ) , .A1( u0_u14_u6_n122 ) , .ZN( u0_u14_u6_n131 ) );
  AND3_X1 u0_u14_u6_U24 (.ZN( u0_u14_u6_n120 ) , .A2( u0_u14_u6_n127 ) , .A1( u0_u14_u6_n132 ) , .A3( u0_u14_u6_n145 ) );
  INV_X1 u0_u14_u6_U25 (.A( u0_u14_u6_n146 ) , .ZN( u0_u14_u6_n163 ) );
  AOI222_X1 u0_u14_u6_U26 (.ZN( u0_u14_u6_n114 ) , .A1( u0_u14_u6_n118 ) , .A2( u0_u14_u6_n126 ) , .B2( u0_u14_u6_n151 ) , .C2( u0_u14_u6_n159 ) , .C1( u0_u14_u6_n168 ) , .B1( u0_u14_u6_n169 ) );
  NOR2_X1 u0_u14_u6_U27 (.A1( u0_u14_u6_n162 ) , .A2( u0_u14_u6_n165 ) , .ZN( u0_u14_u6_n98 ) );
  AOI211_X1 u0_u14_u6_U28 (.B( u0_u14_u6_n149 ) , .A( u0_u14_u6_n150 ) , .C2( u0_u14_u6_n151 ) , .C1( u0_u14_u6_n152 ) , .ZN( u0_u14_u6_n153 ) );
  AOI21_X1 u0_u14_u6_U29 (.B2( u0_u14_u6_n147 ) , .B1( u0_u14_u6_n148 ) , .ZN( u0_u14_u6_n149 ) , .A( u0_u14_u6_n158 ) );
  INV_X1 u0_u14_u6_U3 (.A( u0_u14_u6_n110 ) , .ZN( u0_u14_u6_n166 ) );
  AOI21_X1 u0_u14_u6_U30 (.A( u0_u14_u6_n144 ) , .B2( u0_u14_u6_n145 ) , .B1( u0_u14_u6_n146 ) , .ZN( u0_u14_u6_n150 ) );
  NAND2_X1 u0_u14_u6_U31 (.A2( u0_u14_u6_n143 ) , .ZN( u0_u14_u6_n152 ) , .A1( u0_u14_u6_n166 ) );
  NAND2_X1 u0_u14_u6_U32 (.A1( u0_u14_u6_n144 ) , .ZN( u0_u14_u6_n151 ) , .A2( u0_u14_u6_n158 ) );
  NAND2_X1 u0_u14_u6_U33 (.ZN( u0_u14_u6_n132 ) , .A1( u0_u14_u6_n91 ) , .A2( u0_u14_u6_n97 ) );
  AOI22_X1 u0_u14_u6_U34 (.B2( u0_u14_u6_n110 ) , .B1( u0_u14_u6_n111 ) , .A1( u0_u14_u6_n112 ) , .ZN( u0_u14_u6_n115 ) , .A2( u0_u14_u6_n161 ) );
  NAND4_X1 u0_u14_u6_U35 (.A3( u0_u14_u6_n109 ) , .ZN( u0_u14_u6_n112 ) , .A4( u0_u14_u6_n132 ) , .A2( u0_u14_u6_n147 ) , .A1( u0_u14_u6_n166 ) );
  NOR2_X1 u0_u14_u6_U36 (.ZN( u0_u14_u6_n109 ) , .A1( u0_u14_u6_n170 ) , .A2( u0_u14_u6_n173 ) );
  NOR2_X1 u0_u14_u6_U37 (.A2( u0_u14_u6_n126 ) , .ZN( u0_u14_u6_n155 ) , .A1( u0_u14_u6_n160 ) );
  NAND2_X1 u0_u14_u6_U38 (.ZN( u0_u14_u6_n146 ) , .A2( u0_u14_u6_n94 ) , .A1( u0_u14_u6_n99 ) );
  AOI211_X1 u0_u14_u6_U39 (.B( u0_u14_u6_n134 ) , .A( u0_u14_u6_n135 ) , .C1( u0_u14_u6_n136 ) , .ZN( u0_u14_u6_n137 ) , .C2( u0_u14_u6_n151 ) );
  AOI22_X1 u0_u14_u6_U4 (.B2( u0_u14_u6_n101 ) , .A1( u0_u14_u6_n102 ) , .ZN( u0_u14_u6_n103 ) , .B1( u0_u14_u6_n160 ) , .A2( u0_u14_u6_n161 ) );
  AOI21_X1 u0_u14_u6_U40 (.B2( u0_u14_u6_n132 ) , .B1( u0_u14_u6_n133 ) , .ZN( u0_u14_u6_n134 ) , .A( u0_u14_u6_n158 ) );
  NAND4_X1 u0_u14_u6_U41 (.A4( u0_u14_u6_n127 ) , .A3( u0_u14_u6_n128 ) , .A2( u0_u14_u6_n129 ) , .A1( u0_u14_u6_n130 ) , .ZN( u0_u14_u6_n136 ) );
  AOI21_X1 u0_u14_u6_U42 (.B1( u0_u14_u6_n131 ) , .ZN( u0_u14_u6_n135 ) , .A( u0_u14_u6_n144 ) , .B2( u0_u14_u6_n146 ) );
  INV_X1 u0_u14_u6_U43 (.A( u0_u14_u6_n111 ) , .ZN( u0_u14_u6_n158 ) );
  NAND2_X1 u0_u14_u6_U44 (.ZN( u0_u14_u6_n127 ) , .A1( u0_u14_u6_n91 ) , .A2( u0_u14_u6_n92 ) );
  NAND2_X1 u0_u14_u6_U45 (.ZN( u0_u14_u6_n129 ) , .A2( u0_u14_u6_n95 ) , .A1( u0_u14_u6_n96 ) );
  INV_X1 u0_u14_u6_U46 (.A( u0_u14_u6_n144 ) , .ZN( u0_u14_u6_n159 ) );
  NAND2_X1 u0_u14_u6_U47 (.ZN( u0_u14_u6_n145 ) , .A2( u0_u14_u6_n97 ) , .A1( u0_u14_u6_n98 ) );
  NAND2_X1 u0_u14_u6_U48 (.ZN( u0_u14_u6_n148 ) , .A2( u0_u14_u6_n92 ) , .A1( u0_u14_u6_n94 ) );
  NAND2_X1 u0_u14_u6_U49 (.ZN( u0_u14_u6_n108 ) , .A2( u0_u14_u6_n139 ) , .A1( u0_u14_u6_n144 ) );
  NOR2_X1 u0_u14_u6_U5 (.A1( u0_u14_u6_n118 ) , .ZN( u0_u14_u6_n143 ) , .A2( u0_u14_u6_n168 ) );
  NAND2_X1 u0_u14_u6_U50 (.ZN( u0_u14_u6_n121 ) , .A2( u0_u14_u6_n95 ) , .A1( u0_u14_u6_n97 ) );
  NAND2_X1 u0_u14_u6_U51 (.ZN( u0_u14_u6_n107 ) , .A2( u0_u14_u6_n92 ) , .A1( u0_u14_u6_n95 ) );
  AND2_X1 u0_u14_u6_U52 (.ZN( u0_u14_u6_n118 ) , .A2( u0_u14_u6_n91 ) , .A1( u0_u14_u6_n99 ) );
  NAND2_X1 u0_u14_u6_U53 (.ZN( u0_u14_u6_n147 ) , .A2( u0_u14_u6_n98 ) , .A1( u0_u14_u6_n99 ) );
  NAND2_X1 u0_u14_u6_U54 (.ZN( u0_u14_u6_n128 ) , .A1( u0_u14_u6_n94 ) , .A2( u0_u14_u6_n96 ) );
  NAND2_X1 u0_u14_u6_U55 (.ZN( u0_u14_u6_n119 ) , .A2( u0_u14_u6_n95 ) , .A1( u0_u14_u6_n99 ) );
  NAND2_X1 u0_u14_u6_U56 (.ZN( u0_u14_u6_n123 ) , .A2( u0_u14_u6_n91 ) , .A1( u0_u14_u6_n96 ) );
  NAND2_X1 u0_u14_u6_U57 (.ZN( u0_u14_u6_n100 ) , .A2( u0_u14_u6_n92 ) , .A1( u0_u14_u6_n98 ) );
  NAND2_X1 u0_u14_u6_U58 (.ZN( u0_u14_u6_n122 ) , .A1( u0_u14_u6_n94 ) , .A2( u0_u14_u6_n97 ) );
  INV_X1 u0_u14_u6_U59 (.A( u0_u14_u6_n139 ) , .ZN( u0_u14_u6_n160 ) );
  INV_X1 u0_u14_u6_U6 (.ZN( u0_u14_u6_n172 ) , .A( u0_u14_u6_n88 ) );
  NAND2_X1 u0_u14_u6_U60 (.ZN( u0_u14_u6_n113 ) , .A1( u0_u14_u6_n96 ) , .A2( u0_u14_u6_n98 ) );
  NOR2_X1 u0_u14_u6_U61 (.A2( u0_u14_X_40 ) , .A1( u0_u14_X_41 ) , .ZN( u0_u14_u6_n126 ) );
  NOR2_X1 u0_u14_u6_U62 (.A2( u0_u14_X_39 ) , .A1( u0_u14_X_42 ) , .ZN( u0_u14_u6_n92 ) );
  NOR2_X1 u0_u14_u6_U63 (.A2( u0_u14_X_39 ) , .A1( u0_u14_u6_n156 ) , .ZN( u0_u14_u6_n97 ) );
  NOR2_X1 u0_u14_u6_U64 (.A2( u0_u14_X_38 ) , .A1( u0_u14_u6_n165 ) , .ZN( u0_u14_u6_n95 ) );
  NOR2_X1 u0_u14_u6_U65 (.A2( u0_u14_X_41 ) , .ZN( u0_u14_u6_n111 ) , .A1( u0_u14_u6_n157 ) );
  NOR2_X1 u0_u14_u6_U66 (.A2( u0_u14_X_37 ) , .A1( u0_u14_u6_n162 ) , .ZN( u0_u14_u6_n94 ) );
  NOR2_X1 u0_u14_u6_U67 (.A2( u0_u14_X_37 ) , .A1( u0_u14_X_38 ) , .ZN( u0_u14_u6_n91 ) );
  NAND2_X1 u0_u14_u6_U68 (.A1( u0_u14_X_41 ) , .ZN( u0_u14_u6_n144 ) , .A2( u0_u14_u6_n157 ) );
  NAND2_X1 u0_u14_u6_U69 (.A2( u0_u14_X_40 ) , .A1( u0_u14_X_41 ) , .ZN( u0_u14_u6_n139 ) );
  OAI21_X1 u0_u14_u6_U7 (.A( u0_u14_u6_n159 ) , .B1( u0_u14_u6_n169 ) , .B2( u0_u14_u6_n173 ) , .ZN( u0_u14_u6_n90 ) );
  AND2_X1 u0_u14_u6_U70 (.A1( u0_u14_X_39 ) , .A2( u0_u14_u6_n156 ) , .ZN( u0_u14_u6_n96 ) );
  AND2_X1 u0_u14_u6_U71 (.A1( u0_u14_X_39 ) , .A2( u0_u14_X_42 ) , .ZN( u0_u14_u6_n99 ) );
  INV_X1 u0_u14_u6_U72 (.A( u0_u14_X_40 ) , .ZN( u0_u14_u6_n157 ) );
  INV_X1 u0_u14_u6_U73 (.A( u0_u14_X_37 ) , .ZN( u0_u14_u6_n165 ) );
  INV_X1 u0_u14_u6_U74 (.A( u0_u14_X_38 ) , .ZN( u0_u14_u6_n162 ) );
  INV_X1 u0_u14_u6_U75 (.A( u0_u14_X_42 ) , .ZN( u0_u14_u6_n156 ) );
  NAND4_X1 u0_u14_u6_U76 (.ZN( u0_out14_32 ) , .A4( u0_u14_u6_n103 ) , .A3( u0_u14_u6_n104 ) , .A2( u0_u14_u6_n105 ) , .A1( u0_u14_u6_n106 ) );
  AOI22_X1 u0_u14_u6_U77 (.ZN( u0_u14_u6_n105 ) , .A2( u0_u14_u6_n108 ) , .A1( u0_u14_u6_n118 ) , .B2( u0_u14_u6_n126 ) , .B1( u0_u14_u6_n171 ) );
  AOI22_X1 u0_u14_u6_U78 (.ZN( u0_u14_u6_n104 ) , .A1( u0_u14_u6_n111 ) , .B1( u0_u14_u6_n124 ) , .B2( u0_u14_u6_n151 ) , .A2( u0_u14_u6_n93 ) );
  NAND4_X1 u0_u14_u6_U79 (.ZN( u0_out14_12 ) , .A4( u0_u14_u6_n114 ) , .A3( u0_u14_u6_n115 ) , .A2( u0_u14_u6_n116 ) , .A1( u0_u14_u6_n117 ) );
  AOI22_X1 u0_u14_u6_U8 (.A2( u0_u14_u6_n151 ) , .B2( u0_u14_u6_n161 ) , .A1( u0_u14_u6_n167 ) , .B1( u0_u14_u6_n170 ) , .ZN( u0_u14_u6_n89 ) );
  OAI22_X1 u0_u14_u6_U80 (.B2( u0_u14_u6_n111 ) , .ZN( u0_u14_u6_n116 ) , .B1( u0_u14_u6_n126 ) , .A2( u0_u14_u6_n164 ) , .A1( u0_u14_u6_n167 ) );
  OAI21_X1 u0_u14_u6_U81 (.A( u0_u14_u6_n108 ) , .ZN( u0_u14_u6_n117 ) , .B2( u0_u14_u6_n141 ) , .B1( u0_u14_u6_n163 ) );
  OAI211_X1 u0_u14_u6_U82 (.ZN( u0_out14_22 ) , .B( u0_u14_u6_n137 ) , .A( u0_u14_u6_n138 ) , .C2( u0_u14_u6_n139 ) , .C1( u0_u14_u6_n140 ) );
  AOI22_X1 u0_u14_u6_U83 (.B1( u0_u14_u6_n124 ) , .A2( u0_u14_u6_n125 ) , .A1( u0_u14_u6_n126 ) , .ZN( u0_u14_u6_n138 ) , .B2( u0_u14_u6_n161 ) );
  AND4_X1 u0_u14_u6_U84 (.A3( u0_u14_u6_n119 ) , .A1( u0_u14_u6_n120 ) , .A4( u0_u14_u6_n129 ) , .ZN( u0_u14_u6_n140 ) , .A2( u0_u14_u6_n143 ) );
  OAI211_X1 u0_u14_u6_U85 (.ZN( u0_out14_7 ) , .B( u0_u14_u6_n153 ) , .C2( u0_u14_u6_n154 ) , .C1( u0_u14_u6_n155 ) , .A( u0_u14_u6_n174 ) );
  NOR3_X1 u0_u14_u6_U86 (.A1( u0_u14_u6_n141 ) , .ZN( u0_u14_u6_n154 ) , .A3( u0_u14_u6_n164 ) , .A2( u0_u14_u6_n171 ) );
  INV_X1 u0_u14_u6_U87 (.A( u0_u14_u6_n142 ) , .ZN( u0_u14_u6_n174 ) );
  NAND3_X1 u0_u14_u6_U88 (.A2( u0_u14_u6_n123 ) , .ZN( u0_u14_u6_n125 ) , .A1( u0_u14_u6_n130 ) , .A3( u0_u14_u6_n131 ) );
  NAND3_X1 u0_u14_u6_U89 (.A3( u0_u14_u6_n133 ) , .ZN( u0_u14_u6_n141 ) , .A1( u0_u14_u6_n145 ) , .A2( u0_u14_u6_n148 ) );
  AOI21_X1 u0_u14_u6_U9 (.B1( u0_u14_u6_n107 ) , .B2( u0_u14_u6_n132 ) , .A( u0_u14_u6_n158 ) , .ZN( u0_u14_u6_n88 ) );
  NAND3_X1 u0_u14_u6_U90 (.ZN( u0_u14_u6_n101 ) , .A3( u0_u14_u6_n107 ) , .A2( u0_u14_u6_n121 ) , .A1( u0_u14_u6_n127 ) );
  NAND3_X1 u0_u14_u6_U91 (.ZN( u0_u14_u6_n102 ) , .A3( u0_u14_u6_n130 ) , .A2( u0_u14_u6_n145 ) , .A1( u0_u14_u6_n166 ) );
  NAND3_X1 u0_u14_u6_U92 (.A3( u0_u14_u6_n113 ) , .A1( u0_u14_u6_n119 ) , .A2( u0_u14_u6_n123 ) , .ZN( u0_u14_u6_n93 ) );
  NAND3_X1 u0_u14_u6_U93 (.ZN( u0_u14_u6_n142 ) , .A2( u0_u14_u6_n172 ) , .A3( u0_u14_u6_n89 ) , .A1( u0_u14_u6_n90 ) );
  AND3_X1 u0_u14_u7_U10 (.A3( u0_u14_u7_n110 ) , .A2( u0_u14_u7_n127 ) , .A1( u0_u14_u7_n132 ) , .ZN( u0_u14_u7_n92 ) );
  OAI21_X1 u0_u14_u7_U11 (.A( u0_u14_u7_n161 ) , .B1( u0_u14_u7_n168 ) , .B2( u0_u14_u7_n173 ) , .ZN( u0_u14_u7_n91 ) );
  AOI211_X1 u0_u14_u7_U12 (.A( u0_u14_u7_n117 ) , .ZN( u0_u14_u7_n118 ) , .C2( u0_u14_u7_n126 ) , .C1( u0_u14_u7_n177 ) , .B( u0_u14_u7_n180 ) );
  OAI22_X1 u0_u14_u7_U13 (.B1( u0_u14_u7_n115 ) , .ZN( u0_u14_u7_n117 ) , .A2( u0_u14_u7_n133 ) , .A1( u0_u14_u7_n137 ) , .B2( u0_u14_u7_n162 ) );
  INV_X1 u0_u14_u7_U14 (.A( u0_u14_u7_n116 ) , .ZN( u0_u14_u7_n180 ) );
  NOR3_X1 u0_u14_u7_U15 (.ZN( u0_u14_u7_n115 ) , .A3( u0_u14_u7_n145 ) , .A2( u0_u14_u7_n168 ) , .A1( u0_u14_u7_n169 ) );
  NOR3_X1 u0_u14_u7_U16 (.A2( u0_u14_u7_n134 ) , .A1( u0_u14_u7_n135 ) , .ZN( u0_u14_u7_n136 ) , .A3( u0_u14_u7_n171 ) );
  NOR2_X1 u0_u14_u7_U17 (.A1( u0_u14_u7_n130 ) , .A2( u0_u14_u7_n134 ) , .ZN( u0_u14_u7_n153 ) );
  NOR2_X1 u0_u14_u7_U18 (.ZN( u0_u14_u7_n111 ) , .A2( u0_u14_u7_n134 ) , .A1( u0_u14_u7_n169 ) );
  AOI21_X1 u0_u14_u7_U19 (.ZN( u0_u14_u7_n104 ) , .B2( u0_u14_u7_n112 ) , .B1( u0_u14_u7_n127 ) , .A( u0_u14_u7_n164 ) );
  AOI21_X1 u0_u14_u7_U20 (.ZN( u0_u14_u7_n106 ) , .B1( u0_u14_u7_n133 ) , .B2( u0_u14_u7_n146 ) , .A( u0_u14_u7_n162 ) );
  AOI21_X1 u0_u14_u7_U21 (.A( u0_u14_u7_n101 ) , .ZN( u0_u14_u7_n107 ) , .B2( u0_u14_u7_n128 ) , .B1( u0_u14_u7_n175 ) );
  INV_X1 u0_u14_u7_U22 (.A( u0_u14_u7_n101 ) , .ZN( u0_u14_u7_n165 ) );
  INV_X1 u0_u14_u7_U23 (.A( u0_u14_u7_n138 ) , .ZN( u0_u14_u7_n171 ) );
  INV_X1 u0_u14_u7_U24 (.A( u0_u14_u7_n131 ) , .ZN( u0_u14_u7_n177 ) );
  INV_X1 u0_u14_u7_U25 (.A( u0_u14_u7_n110 ) , .ZN( u0_u14_u7_n174 ) );
  NAND2_X1 u0_u14_u7_U26 (.A1( u0_u14_u7_n129 ) , .A2( u0_u14_u7_n132 ) , .ZN( u0_u14_u7_n149 ) );
  NAND2_X1 u0_u14_u7_U27 (.A1( u0_u14_u7_n113 ) , .A2( u0_u14_u7_n124 ) , .ZN( u0_u14_u7_n130 ) );
  INV_X1 u0_u14_u7_U28 (.A( u0_u14_u7_n128 ) , .ZN( u0_u14_u7_n168 ) );
  INV_X1 u0_u14_u7_U29 (.A( u0_u14_u7_n148 ) , .ZN( u0_u14_u7_n169 ) );
  INV_X1 u0_u14_u7_U3 (.A( u0_u14_u7_n149 ) , .ZN( u0_u14_u7_n175 ) );
  INV_X1 u0_u14_u7_U30 (.A( u0_u14_u7_n112 ) , .ZN( u0_u14_u7_n173 ) );
  INV_X1 u0_u14_u7_U31 (.A( u0_u14_u7_n127 ) , .ZN( u0_u14_u7_n179 ) );
  NOR2_X1 u0_u14_u7_U32 (.ZN( u0_u14_u7_n101 ) , .A2( u0_u14_u7_n150 ) , .A1( u0_u14_u7_n156 ) );
  AOI211_X1 u0_u14_u7_U33 (.B( u0_u14_u7_n154 ) , .A( u0_u14_u7_n155 ) , .C1( u0_u14_u7_n156 ) , .ZN( u0_u14_u7_n157 ) , .C2( u0_u14_u7_n172 ) );
  INV_X1 u0_u14_u7_U34 (.A( u0_u14_u7_n153 ) , .ZN( u0_u14_u7_n172 ) );
  AOI211_X1 u0_u14_u7_U35 (.B( u0_u14_u7_n139 ) , .A( u0_u14_u7_n140 ) , .C2( u0_u14_u7_n141 ) , .ZN( u0_u14_u7_n142 ) , .C1( u0_u14_u7_n156 ) );
  NAND4_X1 u0_u14_u7_U36 (.A3( u0_u14_u7_n127 ) , .A2( u0_u14_u7_n128 ) , .A1( u0_u14_u7_n129 ) , .ZN( u0_u14_u7_n141 ) , .A4( u0_u14_u7_n147 ) );
  AOI21_X1 u0_u14_u7_U37 (.A( u0_u14_u7_n137 ) , .B1( u0_u14_u7_n138 ) , .ZN( u0_u14_u7_n139 ) , .B2( u0_u14_u7_n146 ) );
  OAI22_X1 u0_u14_u7_U38 (.B1( u0_u14_u7_n136 ) , .ZN( u0_u14_u7_n140 ) , .A1( u0_u14_u7_n153 ) , .B2( u0_u14_u7_n162 ) , .A2( u0_u14_u7_n164 ) );
  INV_X1 u0_u14_u7_U39 (.A( u0_u14_u7_n125 ) , .ZN( u0_u14_u7_n161 ) );
  INV_X1 u0_u14_u7_U4 (.A( u0_u14_u7_n154 ) , .ZN( u0_u14_u7_n178 ) );
  AOI21_X1 u0_u14_u7_U40 (.ZN( u0_u14_u7_n123 ) , .B1( u0_u14_u7_n165 ) , .B2( u0_u14_u7_n177 ) , .A( u0_u14_u7_n97 ) );
  AOI21_X1 u0_u14_u7_U41 (.B2( u0_u14_u7_n113 ) , .B1( u0_u14_u7_n124 ) , .A( u0_u14_u7_n125 ) , .ZN( u0_u14_u7_n97 ) );
  INV_X1 u0_u14_u7_U42 (.A( u0_u14_u7_n152 ) , .ZN( u0_u14_u7_n162 ) );
  AOI22_X1 u0_u14_u7_U43 (.A2( u0_u14_u7_n114 ) , .ZN( u0_u14_u7_n119 ) , .B1( u0_u14_u7_n130 ) , .A1( u0_u14_u7_n156 ) , .B2( u0_u14_u7_n165 ) );
  NAND2_X1 u0_u14_u7_U44 (.A2( u0_u14_u7_n112 ) , .ZN( u0_u14_u7_n114 ) , .A1( u0_u14_u7_n175 ) );
  AOI22_X1 u0_u14_u7_U45 (.B2( u0_u14_u7_n149 ) , .B1( u0_u14_u7_n150 ) , .A2( u0_u14_u7_n151 ) , .A1( u0_u14_u7_n152 ) , .ZN( u0_u14_u7_n158 ) );
  NOR2_X1 u0_u14_u7_U46 (.ZN( u0_u14_u7_n137 ) , .A1( u0_u14_u7_n150 ) , .A2( u0_u14_u7_n161 ) );
  AND2_X1 u0_u14_u7_U47 (.ZN( u0_u14_u7_n145 ) , .A2( u0_u14_u7_n98 ) , .A1( u0_u14_u7_n99 ) );
  AOI21_X1 u0_u14_u7_U48 (.ZN( u0_u14_u7_n105 ) , .B2( u0_u14_u7_n110 ) , .A( u0_u14_u7_n125 ) , .B1( u0_u14_u7_n147 ) );
  NAND2_X1 u0_u14_u7_U49 (.ZN( u0_u14_u7_n146 ) , .A1( u0_u14_u7_n95 ) , .A2( u0_u14_u7_n98 ) );
  INV_X1 u0_u14_u7_U5 (.A( u0_u14_u7_n111 ) , .ZN( u0_u14_u7_n170 ) );
  NAND2_X1 u0_u14_u7_U50 (.A2( u0_u14_u7_n103 ) , .ZN( u0_u14_u7_n147 ) , .A1( u0_u14_u7_n93 ) );
  NAND2_X1 u0_u14_u7_U51 (.A1( u0_u14_u7_n103 ) , .ZN( u0_u14_u7_n127 ) , .A2( u0_u14_u7_n99 ) );
  NAND2_X1 u0_u14_u7_U52 (.A2( u0_u14_u7_n102 ) , .A1( u0_u14_u7_n103 ) , .ZN( u0_u14_u7_n133 ) );
  OR2_X1 u0_u14_u7_U53 (.ZN( u0_u14_u7_n126 ) , .A2( u0_u14_u7_n152 ) , .A1( u0_u14_u7_n156 ) );
  NAND2_X1 u0_u14_u7_U54 (.ZN( u0_u14_u7_n112 ) , .A2( u0_u14_u7_n96 ) , .A1( u0_u14_u7_n99 ) );
  NAND2_X1 u0_u14_u7_U55 (.A2( u0_u14_u7_n102 ) , .ZN( u0_u14_u7_n128 ) , .A1( u0_u14_u7_n98 ) );
  INV_X1 u0_u14_u7_U56 (.A( u0_u14_u7_n150 ) , .ZN( u0_u14_u7_n164 ) );
  AND2_X1 u0_u14_u7_U57 (.ZN( u0_u14_u7_n134 ) , .A1( u0_u14_u7_n93 ) , .A2( u0_u14_u7_n98 ) );
  NAND2_X1 u0_u14_u7_U58 (.ZN( u0_u14_u7_n110 ) , .A1( u0_u14_u7_n95 ) , .A2( u0_u14_u7_n96 ) );
  NAND2_X1 u0_u14_u7_U59 (.A2( u0_u14_u7_n102 ) , .ZN( u0_u14_u7_n124 ) , .A1( u0_u14_u7_n96 ) );
  AOI211_X1 u0_u14_u7_U6 (.ZN( u0_u14_u7_n116 ) , .A( u0_u14_u7_n155 ) , .C1( u0_u14_u7_n161 ) , .C2( u0_u14_u7_n171 ) , .B( u0_u14_u7_n94 ) );
  NAND2_X1 u0_u14_u7_U60 (.ZN( u0_u14_u7_n132 ) , .A1( u0_u14_u7_n93 ) , .A2( u0_u14_u7_n96 ) );
  NAND2_X1 u0_u14_u7_U61 (.A2( u0_u14_u7_n103 ) , .ZN( u0_u14_u7_n131 ) , .A1( u0_u14_u7_n95 ) );
  NOR2_X1 u0_u14_u7_U62 (.A2( u0_u14_X_47 ) , .ZN( u0_u14_u7_n150 ) , .A1( u0_u14_u7_n163 ) );
  NOR2_X1 u0_u14_u7_U63 (.A2( u0_u14_X_43 ) , .A1( u0_u14_X_44 ) , .ZN( u0_u14_u7_n103 ) );
  NOR2_X1 u0_u14_u7_U64 (.A2( u0_u14_X_48 ) , .A1( u0_u14_u7_n166 ) , .ZN( u0_u14_u7_n95 ) );
  NOR2_X1 u0_u14_u7_U65 (.A2( u0_u14_X_44 ) , .A1( u0_u14_u7_n167 ) , .ZN( u0_u14_u7_n98 ) );
  NOR2_X1 u0_u14_u7_U66 (.A2( u0_u14_X_45 ) , .A1( u0_u14_X_48 ) , .ZN( u0_u14_u7_n99 ) );
  NOR2_X1 u0_u14_u7_U67 (.A2( u0_u14_X_46 ) , .A1( u0_u14_X_47 ) , .ZN( u0_u14_u7_n152 ) );
  AND2_X1 u0_u14_u7_U68 (.A1( u0_u14_X_47 ) , .ZN( u0_u14_u7_n156 ) , .A2( u0_u14_u7_n163 ) );
  NAND2_X1 u0_u14_u7_U69 (.A2( u0_u14_X_46 ) , .A1( u0_u14_X_47 ) , .ZN( u0_u14_u7_n125 ) );
  OAI222_X1 u0_u14_u7_U7 (.C2( u0_u14_u7_n101 ) , .B2( u0_u14_u7_n111 ) , .A1( u0_u14_u7_n113 ) , .C1( u0_u14_u7_n146 ) , .A2( u0_u14_u7_n162 ) , .B1( u0_u14_u7_n164 ) , .ZN( u0_u14_u7_n94 ) );
  AND2_X1 u0_u14_u7_U70 (.A2( u0_u14_X_43 ) , .A1( u0_u14_X_44 ) , .ZN( u0_u14_u7_n96 ) );
  AND2_X1 u0_u14_u7_U71 (.A2( u0_u14_X_45 ) , .A1( u0_u14_X_48 ) , .ZN( u0_u14_u7_n102 ) );
  AND2_X1 u0_u14_u7_U72 (.A1( u0_u14_X_48 ) , .A2( u0_u14_u7_n166 ) , .ZN( u0_u14_u7_n93 ) );
  INV_X1 u0_u14_u7_U73 (.A( u0_u14_X_46 ) , .ZN( u0_u14_u7_n163 ) );
  AND2_X1 u0_u14_u7_U74 (.A1( u0_u14_X_44 ) , .ZN( u0_u14_u7_n100 ) , .A2( u0_u14_u7_n167 ) );
  INV_X1 u0_u14_u7_U75 (.A( u0_u14_X_43 ) , .ZN( u0_u14_u7_n167 ) );
  INV_X1 u0_u14_u7_U76 (.A( u0_u14_X_45 ) , .ZN( u0_u14_u7_n166 ) );
  NAND4_X1 u0_u14_u7_U77 (.ZN( u0_out14_27 ) , .A4( u0_u14_u7_n118 ) , .A3( u0_u14_u7_n119 ) , .A2( u0_u14_u7_n120 ) , .A1( u0_u14_u7_n121 ) );
  OAI21_X1 u0_u14_u7_U78 (.ZN( u0_u14_u7_n121 ) , .B2( u0_u14_u7_n145 ) , .A( u0_u14_u7_n150 ) , .B1( u0_u14_u7_n174 ) );
  OAI21_X1 u0_u14_u7_U79 (.ZN( u0_u14_u7_n120 ) , .A( u0_u14_u7_n161 ) , .B2( u0_u14_u7_n170 ) , .B1( u0_u14_u7_n179 ) );
  INV_X1 u0_u14_u7_U8 (.A( u0_u14_u7_n133 ) , .ZN( u0_u14_u7_n176 ) );
  NAND4_X1 u0_u14_u7_U80 (.ZN( u0_out14_21 ) , .A4( u0_u14_u7_n157 ) , .A3( u0_u14_u7_n158 ) , .A2( u0_u14_u7_n159 ) , .A1( u0_u14_u7_n160 ) );
  OAI21_X1 u0_u14_u7_U81 (.B1( u0_u14_u7_n145 ) , .ZN( u0_u14_u7_n160 ) , .A( u0_u14_u7_n161 ) , .B2( u0_u14_u7_n177 ) );
  OAI21_X1 u0_u14_u7_U82 (.ZN( u0_u14_u7_n159 ) , .A( u0_u14_u7_n165 ) , .B2( u0_u14_u7_n171 ) , .B1( u0_u14_u7_n174 ) );
  NAND4_X1 u0_u14_u7_U83 (.ZN( u0_out14_15 ) , .A4( u0_u14_u7_n142 ) , .A3( u0_u14_u7_n143 ) , .A2( u0_u14_u7_n144 ) , .A1( u0_u14_u7_n178 ) );
  OR2_X1 u0_u14_u7_U84 (.A2( u0_u14_u7_n125 ) , .A1( u0_u14_u7_n129 ) , .ZN( u0_u14_u7_n144 ) );
  AOI22_X1 u0_u14_u7_U85 (.A2( u0_u14_u7_n126 ) , .ZN( u0_u14_u7_n143 ) , .B2( u0_u14_u7_n165 ) , .B1( u0_u14_u7_n173 ) , .A1( u0_u14_u7_n174 ) );
  NAND4_X1 u0_u14_u7_U86 (.ZN( u0_out14_5 ) , .A4( u0_u14_u7_n108 ) , .A3( u0_u14_u7_n109 ) , .A1( u0_u14_u7_n116 ) , .A2( u0_u14_u7_n123 ) );
  AOI22_X1 u0_u14_u7_U87 (.ZN( u0_u14_u7_n109 ) , .A2( u0_u14_u7_n126 ) , .B2( u0_u14_u7_n145 ) , .B1( u0_u14_u7_n156 ) , .A1( u0_u14_u7_n171 ) );
  NOR4_X1 u0_u14_u7_U88 (.A4( u0_u14_u7_n104 ) , .A3( u0_u14_u7_n105 ) , .A2( u0_u14_u7_n106 ) , .A1( u0_u14_u7_n107 ) , .ZN( u0_u14_u7_n108 ) );
  NAND2_X1 u0_u14_u7_U89 (.A1( u0_u14_u7_n100 ) , .ZN( u0_u14_u7_n148 ) , .A2( u0_u14_u7_n95 ) );
  OAI221_X1 u0_u14_u7_U9 (.C1( u0_u14_u7_n101 ) , .C2( u0_u14_u7_n147 ) , .ZN( u0_u14_u7_n155 ) , .B2( u0_u14_u7_n162 ) , .A( u0_u14_u7_n91 ) , .B1( u0_u14_u7_n92 ) );
  NAND2_X1 u0_u14_u7_U90 (.A1( u0_u14_u7_n100 ) , .ZN( u0_u14_u7_n113 ) , .A2( u0_u14_u7_n93 ) );
  NAND2_X1 u0_u14_u7_U91 (.A1( u0_u14_u7_n100 ) , .ZN( u0_u14_u7_n138 ) , .A2( u0_u14_u7_n99 ) );
  NAND2_X1 u0_u14_u7_U92 (.A1( u0_u14_u7_n100 ) , .A2( u0_u14_u7_n102 ) , .ZN( u0_u14_u7_n129 ) );
  OAI211_X1 u0_u14_u7_U93 (.B( u0_u14_u7_n122 ) , .A( u0_u14_u7_n123 ) , .C2( u0_u14_u7_n124 ) , .ZN( u0_u14_u7_n154 ) , .C1( u0_u14_u7_n162 ) );
  AOI222_X1 u0_u14_u7_U94 (.ZN( u0_u14_u7_n122 ) , .C2( u0_u14_u7_n126 ) , .C1( u0_u14_u7_n145 ) , .B1( u0_u14_u7_n161 ) , .A2( u0_u14_u7_n165 ) , .B2( u0_u14_u7_n170 ) , .A1( u0_u14_u7_n176 ) );
  NAND3_X1 u0_u14_u7_U95 (.A3( u0_u14_u7_n146 ) , .A2( u0_u14_u7_n147 ) , .A1( u0_u14_u7_n148 ) , .ZN( u0_u14_u7_n151 ) );
  NAND3_X1 u0_u14_u7_U96 (.A3( u0_u14_u7_n131 ) , .A2( u0_u14_u7_n132 ) , .A1( u0_u14_u7_n133 ) , .ZN( u0_u14_u7_n135 ) );
  XOR2_X1 u0_u3_U1 (.B( u0_K4_9 ) , .A( u0_R2_6 ) , .Z( u0_u3_X_9 ) );
  XOR2_X1 u0_u3_U12 (.B( u0_K4_43 ) , .A( u0_R2_28 ) , .Z( u0_u3_X_43 ) );
  XOR2_X1 u0_u3_U14 (.B( u0_K4_41 ) , .A( u0_R2_28 ) , .Z( u0_u3_X_41 ) );
  XOR2_X1 u0_u3_U16 (.B( u0_K4_3 ) , .A( u0_R2_2 ) , .Z( u0_u3_X_3 ) );
  XOR2_X1 u0_u3_U18 (.B( u0_K4_38 ) , .A( u0_R2_25 ) , .Z( u0_u3_X_38 ) );
  XOR2_X1 u0_u3_U2 (.B( u0_K4_8 ) , .A( u0_R2_5 ) , .Z( u0_u3_X_8 ) );
  XOR2_X1 u0_u3_U20 (.B( u0_K4_36 ) , .A( u0_R2_25 ) , .Z( u0_u3_X_36 ) );
  XOR2_X1 u0_u3_U23 (.B( u0_K4_33 ) , .A( u0_R2_22 ) , .Z( u0_u3_X_33 ) );
  XOR2_X1 u0_u3_U24 (.B( u0_K4_32 ) , .A( u0_R2_21 ) , .Z( u0_u3_X_32 ) );
  XOR2_X1 u0_u3_U26 (.B( u0_K4_30 ) , .A( u0_R2_21 ) , .Z( u0_u3_X_30 ) );
  XOR2_X1 u0_u3_U27 (.B( u0_K4_2 ) , .A( u0_R2_1 ) , .Z( u0_u3_X_2 ) );
  XOR2_X1 u0_u3_U3 (.B( u0_K4_7 ) , .A( u0_R2_4 ) , .Z( u0_u3_X_7 ) );
  XOR2_X1 u0_u3_U32 (.B( u0_K4_25 ) , .A( u0_R2_16 ) , .Z( u0_u3_X_25 ) );
  XOR2_X1 u0_u3_U34 (.B( u0_K4_23 ) , .A( u0_R2_16 ) , .Z( u0_u3_X_23 ) );
  XOR2_X1 u0_u3_U36 (.B( u0_K4_21 ) , .A( u0_R2_14 ) , .Z( u0_u3_X_21 ) );
  XOR2_X1 u0_u3_U37 (.B( u0_K4_20 ) , .A( u0_R2_13 ) , .Z( u0_u3_X_20 ) );
  XOR2_X1 u0_u3_U38 (.B( u0_K4_1 ) , .A( u0_R2_32 ) , .Z( u0_u3_X_1 ) );
  XOR2_X1 u0_u3_U39 (.B( u0_K4_19 ) , .A( u0_R2_12 ) , .Z( u0_u3_X_19 ) );
  XOR2_X1 u0_u3_U4 (.B( u0_K4_6 ) , .A( u0_R2_5 ) , .Z( u0_u3_X_6 ) );
  XOR2_X1 u0_u3_U40 (.B( u0_K4_18 ) , .A( u0_R2_13 ) , .Z( u0_u3_X_18 ) );
  XOR2_X1 u0_u3_U41 (.B( u0_K4_17 ) , .A( u0_R2_12 ) , .Z( u0_u3_X_17 ) );
  XOR2_X1 u0_u3_U42 (.B( u0_K4_16 ) , .A( u0_R2_11 ) , .Z( u0_u3_X_16 ) );
  XOR2_X1 u0_u3_U43 (.B( u0_K4_15 ) , .A( u0_R2_10 ) , .Z( u0_u3_X_15 ) );
  XOR2_X1 u0_u3_U44 (.B( u0_K4_14 ) , .A( u0_R2_9 ) , .Z( u0_u3_X_14 ) );
  XOR2_X1 u0_u3_U45 (.B( u0_K4_13 ) , .A( u0_R2_8 ) , .Z( u0_u3_X_13 ) );
  XOR2_X1 u0_u3_U46 (.B( u0_K4_12 ) , .A( u0_R2_9 ) , .Z( u0_u3_X_12 ) );
  XOR2_X1 u0_u3_U47 (.B( u0_K4_11 ) , .A( u0_R2_8 ) , .Z( u0_u3_X_11 ) );
  XOR2_X1 u0_u3_U48 (.B( u0_K4_10 ) , .A( u0_R2_7 ) , .Z( u0_u3_X_10 ) );
  XOR2_X1 u0_u3_U5 (.B( u0_K4_5 ) , .A( u0_R2_4 ) , .Z( u0_u3_X_5 ) );
  XOR2_X1 u0_u3_U6 (.B( u0_K4_4 ) , .A( u0_R2_3 ) , .Z( u0_u3_X_4 ) );
  XOR2_X1 u0_u3_U7 (.B( u0_K4_48 ) , .A( u0_R2_1 ) , .Z( u0_u3_X_48 ) );
  XOR2_X1 u0_u3_U8 (.B( u0_K4_47 ) , .A( u0_R2_32 ) , .Z( u0_u3_X_47 ) );
  AND2_X1 u0_u3_u0_U10 (.A1( u0_u3_u0_n133 ) , .ZN( u0_u3_u0_n143 ) , .A2( u0_u3_u0_n152 ) );
  AND2_X1 u0_u3_u0_U11 (.ZN( u0_u3_u0_n109 ) , .A1( u0_u3_u0_n132 ) , .A2( u0_u3_u0_n142 ) );
  AND2_X1 u0_u3_u0_U12 (.A2( u0_u3_u0_n131 ) , .A1( u0_u3_u0_n132 ) , .ZN( u0_u3_u0_n153 ) );
  AND2_X1 u0_u3_u0_U13 (.A1( u0_u3_u0_n110 ) , .A2( u0_u3_u0_n127 ) , .ZN( u0_u3_u0_n147 ) );
  INV_X1 u0_u3_u0_U14 (.A( u0_u3_u0_n145 ) , .ZN( u0_u3_u0_n175 ) );
  NOR2_X1 u0_u3_u0_U15 (.A2( u0_u3_u0_n138 ) , .ZN( u0_u3_u0_n149 ) , .A1( u0_u3_u0_n162 ) );
  AOI21_X1 u0_u3_u0_U16 (.B1( u0_u3_u0_n105 ) , .ZN( u0_u3_u0_n134 ) , .A( u0_u3_u0_n167 ) , .B2( u0_u3_u0_n95 ) );
  OAI22_X1 u0_u3_u0_U17 (.B1( u0_u3_u0_n133 ) , .A1( u0_u3_u0_n146 ) , .B2( u0_u3_u0_n149 ) , .A2( u0_u3_u0_n92 ) , .ZN( u0_u3_u0_n93 ) );
  AND3_X1 u0_u3_u0_U18 (.A3( u0_u3_u0_n123 ) , .A2( u0_u3_u0_n127 ) , .A1( u0_u3_u0_n150 ) , .ZN( u0_u3_u0_n92 ) );
  OAI22_X1 u0_u3_u0_U19 (.B1( u0_u3_u0_n127 ) , .ZN( u0_u3_u0_n128 ) , .A1( u0_u3_u0_n140 ) , .A2( u0_u3_u0_n148 ) , .B2( u0_u3_u0_n149 ) );
  NOR2_X1 u0_u3_u0_U20 (.A1( u0_u3_u0_n165 ) , .A2( u0_u3_u0_n166 ) , .ZN( u0_u3_u0_n97 ) );
  AOI22_X1 u0_u3_u0_U21 (.B2( u0_u3_u0_n111 ) , .A2( u0_u3_u0_n112 ) , .ZN( u0_u3_u0_n113 ) , .B1( u0_u3_u0_n120 ) , .A1( u0_u3_u0_n162 ) );
  NAND2_X1 u0_u3_u0_U22 (.A2( u0_u3_u0_n104 ) , .A1( u0_u3_u0_n105 ) , .ZN( u0_u3_u0_n151 ) );
  INV_X1 u0_u3_u0_U23 (.A( u0_u3_u0_n138 ) , .ZN( u0_u3_u0_n163 ) );
  INV_X1 u0_u3_u0_U24 (.A( u0_u3_u0_n120 ) , .ZN( u0_u3_u0_n160 ) );
  NAND2_X1 u0_u3_u0_U25 (.A2( u0_u3_u0_n102 ) , .ZN( u0_u3_u0_n133 ) , .A1( u0_u3_u0_n94 ) );
  NAND2_X1 u0_u3_u0_U26 (.ZN( u0_u3_u0_n110 ) , .A1( u0_u3_u0_n94 ) , .A2( u0_u3_u0_n96 ) );
  AOI21_X1 u0_u3_u0_U27 (.ZN( u0_u3_u0_n106 ) , .B1( u0_u3_u0_n109 ) , .B2( u0_u3_u0_n143 ) , .A( u0_u3_u0_n146 ) );
  AOI21_X1 u0_u3_u0_U28 (.B1( u0_u3_u0_n129 ) , .B2( u0_u3_u0_n131 ) , .A( u0_u3_u0_n140 ) , .ZN( u0_u3_u0_n98 ) );
  NAND2_X1 u0_u3_u0_U29 (.A2( u0_u3_u0_n104 ) , .ZN( u0_u3_u0_n116 ) , .A1( u0_u3_u0_n94 ) );
  INV_X1 u0_u3_u0_U3 (.A( u0_u3_u0_n115 ) , .ZN( u0_u3_u0_n168 ) );
  NOR2_X1 u0_u3_u0_U30 (.A1( u0_u3_u0_n122 ) , .ZN( u0_u3_u0_n145 ) , .A2( u0_u3_u0_n169 ) );
  OAI221_X1 u0_u3_u0_U31 (.C1( u0_u3_u0_n114 ) , .ZN( u0_u3_u0_n122 ) , .B1( u0_u3_u0_n140 ) , .B2( u0_u3_u0_n143 ) , .C2( u0_u3_u0_n149 ) , .A( u0_u3_u0_n174 ) );
  AOI211_X1 u0_u3_u0_U32 (.B( u0_u3_u0_n117 ) , .A( u0_u3_u0_n118 ) , .C2( u0_u3_u0_n119 ) , .C1( u0_u3_u0_n120 ) , .ZN( u0_u3_u0_n121 ) );
  NAND2_X1 u0_u3_u0_U33 (.A2( u0_u3_u0_n105 ) , .ZN( u0_u3_u0_n142 ) , .A1( u0_u3_u0_n96 ) );
  NAND2_X1 u0_u3_u0_U34 (.A1( u0_u3_u0_n102 ) , .A2( u0_u3_u0_n105 ) , .ZN( u0_u3_u0_n127 ) );
  NAND2_X1 u0_u3_u0_U35 (.A1( u0_u3_u0_n103 ) , .A2( u0_u3_u0_n104 ) , .ZN( u0_u3_u0_n152 ) );
  INV_X1 u0_u3_u0_U36 (.A( u0_u3_u0_n140 ) , .ZN( u0_u3_u0_n162 ) );
  NAND2_X1 u0_u3_u0_U37 (.A2( u0_u3_u0_n102 ) , .A1( u0_u3_u0_n103 ) , .ZN( u0_u3_u0_n141 ) );
  NAND2_X1 u0_u3_u0_U38 (.ZN( u0_u3_u0_n114 ) , .A2( u0_u3_u0_n94 ) , .A1( u0_u3_u0_n95 ) );
  NAND2_X1 u0_u3_u0_U39 (.A1( u0_u3_u0_n103 ) , .ZN( u0_u3_u0_n132 ) , .A2( u0_u3_u0_n96 ) );
  AOI21_X1 u0_u3_u0_U4 (.B1( u0_u3_u0_n116 ) , .ZN( u0_u3_u0_n117 ) , .B2( u0_u3_u0_n131 ) , .A( u0_u3_u0_n163 ) );
  INV_X1 u0_u3_u0_U40 (.ZN( u0_u3_u0_n174 ) , .A( u0_u3_u0_n90 ) );
  OAI222_X1 u0_u3_u0_U41 (.C1( u0_u3_u0_n110 ) , .A1( u0_u3_u0_n127 ) , .B2( u0_u3_u0_n130 ) , .B1( u0_u3_u0_n146 ) , .A2( u0_u3_u0_n160 ) , .C2( u0_u3_u0_n163 ) , .ZN( u0_u3_u0_n90 ) );
  OR3_X1 u0_u3_u0_U42 (.A3( u0_u3_u0_n154 ) , .A2( u0_u3_u0_n155 ) , .A1( u0_u3_u0_n156 ) , .ZN( u0_u3_u0_n157 ) );
  AOI21_X1 u0_u3_u0_U43 (.A( u0_u3_u0_n146 ) , .B2( u0_u3_u0_n147 ) , .B1( u0_u3_u0_n148 ) , .ZN( u0_u3_u0_n156 ) );
  AOI21_X1 u0_u3_u0_U44 (.B2( u0_u3_u0_n152 ) , .B1( u0_u3_u0_n153 ) , .ZN( u0_u3_u0_n154 ) , .A( u0_u3_u0_n160 ) );
  AOI21_X1 u0_u3_u0_U45 (.A( u0_u3_u0_n149 ) , .B2( u0_u3_u0_n150 ) , .B1( u0_u3_u0_n151 ) , .ZN( u0_u3_u0_n155 ) );
  INV_X1 u0_u3_u0_U46 (.A( u0_u3_u0_n101 ) , .ZN( u0_u3_u0_n173 ) );
  OAI211_X1 u0_u3_u0_U47 (.B( u0_u3_u0_n100 ) , .ZN( u0_u3_u0_n101 ) , .C2( u0_u3_u0_n142 ) , .C1( u0_u3_u0_n163 ) , .A( u0_u3_u0_n171 ) );
  INV_X1 u0_u3_u0_U48 (.ZN( u0_u3_u0_n171 ) , .A( u0_u3_u0_n93 ) );
  AOI211_X1 u0_u3_u0_U49 (.ZN( u0_u3_u0_n100 ) , .C1( u0_u3_u0_n120 ) , .A( u0_u3_u0_n125 ) , .B( u0_u3_u0_n98 ) , .C2( u0_u3_u0_n99 ) );
  AOI21_X1 u0_u3_u0_U5 (.B2( u0_u3_u0_n133 ) , .ZN( u0_u3_u0_n136 ) , .B1( u0_u3_u0_n153 ) , .A( u0_u3_u0_n160 ) );
  NOR2_X1 u0_u3_u0_U50 (.A2( u0_u3_X_4 ) , .A1( u0_u3_X_5 ) , .ZN( u0_u3_u0_n120 ) );
  NOR2_X1 u0_u3_u0_U51 (.A2( u0_u3_X_3 ) , .A1( u0_u3_X_6 ) , .ZN( u0_u3_u0_n96 ) );
  NOR2_X1 u0_u3_u0_U52 (.A2( u0_u3_X_6 ) , .ZN( u0_u3_u0_n102 ) , .A1( u0_u3_u0_n164 ) );
  NOR2_X1 u0_u3_u0_U53 (.A2( u0_u3_X_1 ) , .ZN( u0_u3_u0_n103 ) , .A1( u0_u3_u0_n165 ) );
  NAND2_X1 u0_u3_u0_U54 (.A2( u0_u3_X_4 ) , .A1( u0_u3_X_5 ) , .ZN( u0_u3_u0_n146 ) );
  NOR2_X1 u0_u3_u0_U55 (.A2( u0_u3_X_5 ) , .ZN( u0_u3_u0_n138 ) , .A1( u0_u3_u0_n161 ) );
  NAND2_X1 u0_u3_u0_U56 (.A1( u0_u3_X_5 ) , .ZN( u0_u3_u0_n140 ) , .A2( u0_u3_u0_n161 ) );
  AND2_X1 u0_u3_u0_U57 (.A2( u0_u3_X_3 ) , .A1( u0_u3_X_6 ) , .ZN( u0_u3_u0_n104 ) );
  AND2_X1 u0_u3_u0_U58 (.A1( u0_u3_X_6 ) , .A2( u0_u3_u0_n164 ) , .ZN( u0_u3_u0_n95 ) );
  INV_X1 u0_u3_u0_U59 (.A( u0_u3_X_4 ) , .ZN( u0_u3_u0_n161 ) );
  NOR2_X1 u0_u3_u0_U6 (.A1( u0_u3_u0_n110 ) , .ZN( u0_u3_u0_n125 ) , .A2( u0_u3_u0_n160 ) );
  INV_X1 u0_u3_u0_U60 (.A( u0_u3_X_1 ) , .ZN( u0_u3_u0_n166 ) );
  INV_X1 u0_u3_u0_U61 (.A( u0_u3_X_3 ) , .ZN( u0_u3_u0_n164 ) );
  INV_X1 u0_u3_u0_U62 (.A( u0_u3_u0_n128 ) , .ZN( u0_u3_u0_n170 ) );
  AOI211_X1 u0_u3_u0_U63 (.B( u0_u3_u0_n135 ) , .A( u0_u3_u0_n136 ) , .C2( u0_u3_u0_n137 ) , .C1( u0_u3_u0_n138 ) , .ZN( u0_u3_u0_n139 ) );
  OR4_X1 u0_u3_u0_U64 (.ZN( u0_out3_31 ) , .A4( u0_u3_u0_n157 ) , .A2( u0_u3_u0_n158 ) , .A1( u0_u3_u0_n159 ) , .A3( u0_u3_u0_n175 ) );
  AOI21_X1 u0_u3_u0_U65 (.A( u0_u3_u0_n140 ) , .B2( u0_u3_u0_n141 ) , .B1( u0_u3_u0_n142 ) , .ZN( u0_u3_u0_n159 ) );
  OR4_X1 u0_u3_u0_U66 (.ZN( u0_out3_17 ) , .A4( u0_u3_u0_n124 ) , .A2( u0_u3_u0_n125 ) , .A1( u0_u3_u0_n126 ) , .A3( u0_u3_u0_n172 ) );
  AOI21_X1 u0_u3_u0_U67 (.B2( u0_u3_u0_n109 ) , .ZN( u0_u3_u0_n126 ) , .B1( u0_u3_u0_n130 ) , .A( u0_u3_u0_n163 ) );
  INV_X1 u0_u3_u0_U68 (.A( u0_u3_u0_n113 ) , .ZN( u0_u3_u0_n172 ) );
  INV_X1 u0_u3_u0_U69 (.ZN( u0_u3_u0_n176 ) , .A( u0_u3_u0_n91 ) );
  OAI21_X1 u0_u3_u0_U7 (.B1( u0_u3_u0_n152 ) , .B2( u0_u3_u0_n160 ) , .A( u0_u3_u0_n174 ) , .ZN( u0_u3_u0_n91 ) );
  AOI211_X1 u0_u3_u0_U70 (.B( u0_u3_u0_n106 ) , .A( u0_u3_u0_n107 ) , .ZN( u0_u3_u0_n108 ) , .C2( u0_u3_u0_n115 ) , .C1( u0_u3_u0_n162 ) );
  AOI21_X1 u0_u3_u0_U71 (.B2( u0_u3_u0_n143 ) , .B1( u0_u3_u0_n144 ) , .ZN( u0_u3_u0_n158 ) , .A( u0_u3_u0_n163 ) );
  AOI21_X1 u0_u3_u0_U72 (.ZN( u0_u3_u0_n118 ) , .B2( u0_u3_u0_n144 ) , .A( u0_u3_u0_n146 ) , .B1( u0_u3_u0_n168 ) );
  INV_X1 u0_u3_u0_U73 (.A( u0_u3_u0_n144 ) , .ZN( u0_u3_u0_n167 ) );
  NOR2_X1 u0_u3_u0_U74 (.A2( u0_u3_X_1 ) , .A1( u0_u3_X_2 ) , .ZN( u0_u3_u0_n94 ) );
  NOR2_X1 u0_u3_u0_U75 (.A2( u0_u3_X_2 ) , .ZN( u0_u3_u0_n105 ) , .A1( u0_u3_u0_n166 ) );
  INV_X1 u0_u3_u0_U76 (.A( u0_u3_X_2 ) , .ZN( u0_u3_u0_n165 ) );
  OR2_X1 u0_u3_u0_U77 (.A2( u0_u3_u0_n129 ) , .A1( u0_u3_u0_n146 ) , .ZN( u0_u3_u0_n88 ) );
  OR2_X1 u0_u3_u0_U78 (.A1( u0_u3_u0_n123 ) , .A2( u0_u3_u0_n149 ) , .ZN( u0_u3_u0_n89 ) );
  NAND3_X1 u0_u3_u0_U79 (.ZN( u0_u3_u0_n124 ) , .A3( u0_u3_u0_n145 ) , .A1( u0_u3_u0_n88 ) , .A2( u0_u3_u0_n89 ) );
  AND2_X1 u0_u3_u0_U8 (.A1( u0_u3_u0_n116 ) , .A2( u0_u3_u0_n123 ) , .ZN( u0_u3_u0_n148 ) );
  AND3_X1 u0_u3_u0_U80 (.A2( u0_u3_u0_n114 ) , .ZN( u0_u3_u0_n129 ) , .A3( u0_u3_u0_n132 ) , .A1( u0_u3_u0_n150 ) );
  NAND2_X1 u0_u3_u0_U81 (.A2( u0_u3_u0_n103 ) , .ZN( u0_u3_u0_n123 ) , .A1( u0_u3_u0_n95 ) );
  AOI21_X1 u0_u3_u0_U82 (.B1( u0_u3_u0_n134 ) , .ZN( u0_u3_u0_n135 ) , .A( u0_u3_u0_n146 ) , .B2( u0_u3_u0_n168 ) );
  OAI22_X1 u0_u3_u0_U83 (.ZN( u0_u3_u0_n107 ) , .A2( u0_u3_u0_n134 ) , .B1( u0_u3_u0_n148 ) , .A1( u0_u3_u0_n149 ) , .B2( u0_u3_u0_n163 ) );
  NAND2_X1 u0_u3_u0_U84 (.ZN( u0_u3_u0_n112 ) , .A2( u0_u3_u0_n134 ) , .A1( u0_u3_u0_n147 ) );
  INV_X1 u0_u3_u0_U85 (.A( u0_u3_u0_n121 ) , .ZN( u0_u3_u0_n169 ) );
  NAND2_X1 u0_u3_u0_U86 (.ZN( u0_u3_u0_n150 ) , .A1( u0_u3_u0_n95 ) , .A2( u0_u3_u0_n97 ) );
  NAND2_X1 u0_u3_u0_U87 (.A1( u0_u3_u0_n102 ) , .ZN( u0_u3_u0_n131 ) , .A2( u0_u3_u0_n97 ) );
  NAND3_X1 u0_u3_u0_U88 (.ZN( u0_out3_23 ) , .A3( u0_u3_u0_n139 ) , .A1( u0_u3_u0_n170 ) , .A2( u0_u3_u0_n173 ) );
  NAND3_X1 u0_u3_u0_U89 (.A3( u0_u3_u0_n129 ) , .A2( u0_u3_u0_n130 ) , .ZN( u0_u3_u0_n137 ) , .A1( u0_u3_u0_n152 ) );
  NAND2_X1 u0_u3_u0_U9 (.ZN( u0_u3_u0_n115 ) , .A1( u0_u3_u0_n141 ) , .A2( u0_u3_u0_n151 ) );
  NAND3_X1 u0_u3_u0_U90 (.ZN( u0_u3_u0_n119 ) , .A3( u0_u3_u0_n134 ) , .A2( u0_u3_u0_n141 ) , .A1( u0_u3_u0_n150 ) );
  NAND3_X1 u0_u3_u0_U91 (.ZN( u0_u3_u0_n111 ) , .A2( u0_u3_u0_n116 ) , .A3( u0_u3_u0_n142 ) , .A1( u0_u3_u0_n151 ) );
  NAND3_X1 u0_u3_u0_U92 (.ZN( u0_out3_9 ) , .A3( u0_u3_u0_n108 ) , .A2( u0_u3_u0_n173 ) , .A1( u0_u3_u0_n176 ) );
  NAND3_X1 u0_u3_u0_U93 (.A2( u0_u3_u0_n130 ) , .A1( u0_u3_u0_n134 ) , .A3( u0_u3_u0_n148 ) , .ZN( u0_u3_u0_n99 ) );
  NAND2_X1 u0_u3_u0_U94 (.A1( u0_u3_u0_n104 ) , .ZN( u0_u3_u0_n130 ) , .A2( u0_u3_u0_n97 ) );
  NAND2_X1 u0_u3_u0_U95 (.ZN( u0_u3_u0_n144 ) , .A1( u0_u3_u0_n96 ) , .A2( u0_u3_u0_n97 ) );
  NOR2_X1 u0_u3_u1_U10 (.A1( u0_u3_u1_n112 ) , .A2( u0_u3_u1_n116 ) , .ZN( u0_u3_u1_n118 ) );
  NAND3_X1 u0_u3_u1_U100 (.ZN( u0_u3_u1_n113 ) , .A1( u0_u3_u1_n120 ) , .A3( u0_u3_u1_n133 ) , .A2( u0_u3_u1_n155 ) );
  OAI21_X1 u0_u3_u1_U11 (.ZN( u0_u3_u1_n101 ) , .B1( u0_u3_u1_n141 ) , .A( u0_u3_u1_n146 ) , .B2( u0_u3_u1_n183 ) );
  AOI21_X1 u0_u3_u1_U12 (.B2( u0_u3_u1_n155 ) , .B1( u0_u3_u1_n156 ) , .ZN( u0_u3_u1_n157 ) , .A( u0_u3_u1_n174 ) );
  NAND2_X1 u0_u3_u1_U13 (.ZN( u0_u3_u1_n140 ) , .A2( u0_u3_u1_n150 ) , .A1( u0_u3_u1_n155 ) );
  NAND2_X1 u0_u3_u1_U14 (.A1( u0_u3_u1_n131 ) , .ZN( u0_u3_u1_n147 ) , .A2( u0_u3_u1_n153 ) );
  INV_X1 u0_u3_u1_U15 (.A( u0_u3_u1_n139 ) , .ZN( u0_u3_u1_n174 ) );
  OR4_X1 u0_u3_u1_U16 (.A4( u0_u3_u1_n106 ) , .A3( u0_u3_u1_n107 ) , .ZN( u0_u3_u1_n108 ) , .A1( u0_u3_u1_n117 ) , .A2( u0_u3_u1_n184 ) );
  AOI21_X1 u0_u3_u1_U17 (.ZN( u0_u3_u1_n106 ) , .A( u0_u3_u1_n112 ) , .B1( u0_u3_u1_n154 ) , .B2( u0_u3_u1_n156 ) );
  INV_X1 u0_u3_u1_U18 (.A( u0_u3_u1_n101 ) , .ZN( u0_u3_u1_n184 ) );
  AOI21_X1 u0_u3_u1_U19 (.ZN( u0_u3_u1_n107 ) , .B1( u0_u3_u1_n134 ) , .B2( u0_u3_u1_n149 ) , .A( u0_u3_u1_n174 ) );
  INV_X1 u0_u3_u1_U20 (.A( u0_u3_u1_n112 ) , .ZN( u0_u3_u1_n171 ) );
  NAND2_X1 u0_u3_u1_U21 (.ZN( u0_u3_u1_n141 ) , .A1( u0_u3_u1_n153 ) , .A2( u0_u3_u1_n156 ) );
  AND2_X1 u0_u3_u1_U22 (.A1( u0_u3_u1_n123 ) , .ZN( u0_u3_u1_n134 ) , .A2( u0_u3_u1_n161 ) );
  NAND2_X1 u0_u3_u1_U23 (.A2( u0_u3_u1_n115 ) , .A1( u0_u3_u1_n116 ) , .ZN( u0_u3_u1_n148 ) );
  NAND2_X1 u0_u3_u1_U24 (.A2( u0_u3_u1_n133 ) , .A1( u0_u3_u1_n135 ) , .ZN( u0_u3_u1_n159 ) );
  NAND2_X1 u0_u3_u1_U25 (.A2( u0_u3_u1_n115 ) , .A1( u0_u3_u1_n120 ) , .ZN( u0_u3_u1_n132 ) );
  INV_X1 u0_u3_u1_U26 (.A( u0_u3_u1_n154 ) , .ZN( u0_u3_u1_n178 ) );
  INV_X1 u0_u3_u1_U27 (.A( u0_u3_u1_n151 ) , .ZN( u0_u3_u1_n183 ) );
  AND2_X1 u0_u3_u1_U28 (.A1( u0_u3_u1_n129 ) , .A2( u0_u3_u1_n133 ) , .ZN( u0_u3_u1_n149 ) );
  INV_X1 u0_u3_u1_U29 (.A( u0_u3_u1_n131 ) , .ZN( u0_u3_u1_n180 ) );
  INV_X1 u0_u3_u1_U3 (.A( u0_u3_u1_n159 ) , .ZN( u0_u3_u1_n182 ) );
  AOI221_X1 u0_u3_u1_U30 (.B1( u0_u3_u1_n140 ) , .ZN( u0_u3_u1_n167 ) , .B2( u0_u3_u1_n172 ) , .C2( u0_u3_u1_n175 ) , .C1( u0_u3_u1_n178 ) , .A( u0_u3_u1_n188 ) );
  INV_X1 u0_u3_u1_U31 (.ZN( u0_u3_u1_n188 ) , .A( u0_u3_u1_n97 ) );
  AOI211_X1 u0_u3_u1_U32 (.A( u0_u3_u1_n118 ) , .C1( u0_u3_u1_n132 ) , .C2( u0_u3_u1_n139 ) , .B( u0_u3_u1_n96 ) , .ZN( u0_u3_u1_n97 ) );
  AOI21_X1 u0_u3_u1_U33 (.B2( u0_u3_u1_n121 ) , .B1( u0_u3_u1_n135 ) , .A( u0_u3_u1_n152 ) , .ZN( u0_u3_u1_n96 ) );
  OAI221_X1 u0_u3_u1_U34 (.A( u0_u3_u1_n119 ) , .C2( u0_u3_u1_n129 ) , .ZN( u0_u3_u1_n138 ) , .B2( u0_u3_u1_n152 ) , .C1( u0_u3_u1_n174 ) , .B1( u0_u3_u1_n187 ) );
  INV_X1 u0_u3_u1_U35 (.A( u0_u3_u1_n148 ) , .ZN( u0_u3_u1_n187 ) );
  AOI211_X1 u0_u3_u1_U36 (.B( u0_u3_u1_n117 ) , .A( u0_u3_u1_n118 ) , .ZN( u0_u3_u1_n119 ) , .C2( u0_u3_u1_n146 ) , .C1( u0_u3_u1_n159 ) );
  NOR2_X1 u0_u3_u1_U37 (.A1( u0_u3_u1_n168 ) , .A2( u0_u3_u1_n176 ) , .ZN( u0_u3_u1_n98 ) );
  NAND2_X1 u0_u3_u1_U38 (.A1( u0_u3_u1_n128 ) , .ZN( u0_u3_u1_n146 ) , .A2( u0_u3_u1_n160 ) );
  NAND2_X1 u0_u3_u1_U39 (.A2( u0_u3_u1_n112 ) , .ZN( u0_u3_u1_n139 ) , .A1( u0_u3_u1_n152 ) );
  AOI221_X1 u0_u3_u1_U4 (.A( u0_u3_u1_n138 ) , .C2( u0_u3_u1_n139 ) , .C1( u0_u3_u1_n140 ) , .B2( u0_u3_u1_n141 ) , .ZN( u0_u3_u1_n142 ) , .B1( u0_u3_u1_n175 ) );
  NAND2_X1 u0_u3_u1_U40 (.A1( u0_u3_u1_n105 ) , .ZN( u0_u3_u1_n156 ) , .A2( u0_u3_u1_n99 ) );
  NOR2_X1 u0_u3_u1_U41 (.ZN( u0_u3_u1_n117 ) , .A1( u0_u3_u1_n121 ) , .A2( u0_u3_u1_n160 ) );
  OAI21_X1 u0_u3_u1_U42 (.B2( u0_u3_u1_n123 ) , .ZN( u0_u3_u1_n145 ) , .B1( u0_u3_u1_n160 ) , .A( u0_u3_u1_n185 ) );
  INV_X1 u0_u3_u1_U43 (.A( u0_u3_u1_n122 ) , .ZN( u0_u3_u1_n185 ) );
  AOI21_X1 u0_u3_u1_U44 (.B2( u0_u3_u1_n120 ) , .B1( u0_u3_u1_n121 ) , .ZN( u0_u3_u1_n122 ) , .A( u0_u3_u1_n128 ) );
  AOI21_X1 u0_u3_u1_U45 (.A( u0_u3_u1_n128 ) , .B2( u0_u3_u1_n129 ) , .ZN( u0_u3_u1_n130 ) , .B1( u0_u3_u1_n150 ) );
  NAND2_X1 u0_u3_u1_U46 (.ZN( u0_u3_u1_n112 ) , .A1( u0_u3_u1_n169 ) , .A2( u0_u3_u1_n170 ) );
  NAND2_X1 u0_u3_u1_U47 (.ZN( u0_u3_u1_n129 ) , .A2( u0_u3_u1_n95 ) , .A1( u0_u3_u1_n98 ) );
  NAND2_X1 u0_u3_u1_U48 (.A1( u0_u3_u1_n102 ) , .ZN( u0_u3_u1_n154 ) , .A2( u0_u3_u1_n99 ) );
  NAND2_X1 u0_u3_u1_U49 (.A2( u0_u3_u1_n100 ) , .ZN( u0_u3_u1_n135 ) , .A1( u0_u3_u1_n99 ) );
  AOI211_X1 u0_u3_u1_U5 (.ZN( u0_u3_u1_n124 ) , .A( u0_u3_u1_n138 ) , .C2( u0_u3_u1_n139 ) , .B( u0_u3_u1_n145 ) , .C1( u0_u3_u1_n147 ) );
  AOI21_X1 u0_u3_u1_U50 (.A( u0_u3_u1_n152 ) , .B2( u0_u3_u1_n153 ) , .B1( u0_u3_u1_n154 ) , .ZN( u0_u3_u1_n158 ) );
  INV_X1 u0_u3_u1_U51 (.A( u0_u3_u1_n160 ) , .ZN( u0_u3_u1_n175 ) );
  NAND2_X1 u0_u3_u1_U52 (.A1( u0_u3_u1_n100 ) , .ZN( u0_u3_u1_n116 ) , .A2( u0_u3_u1_n95 ) );
  NAND2_X1 u0_u3_u1_U53 (.A1( u0_u3_u1_n102 ) , .ZN( u0_u3_u1_n131 ) , .A2( u0_u3_u1_n95 ) );
  NAND2_X1 u0_u3_u1_U54 (.A2( u0_u3_u1_n104 ) , .ZN( u0_u3_u1_n121 ) , .A1( u0_u3_u1_n98 ) );
  NAND2_X1 u0_u3_u1_U55 (.A1( u0_u3_u1_n103 ) , .ZN( u0_u3_u1_n153 ) , .A2( u0_u3_u1_n98 ) );
  NAND2_X1 u0_u3_u1_U56 (.A2( u0_u3_u1_n104 ) , .A1( u0_u3_u1_n105 ) , .ZN( u0_u3_u1_n133 ) );
  NAND2_X1 u0_u3_u1_U57 (.ZN( u0_u3_u1_n150 ) , .A2( u0_u3_u1_n98 ) , .A1( u0_u3_u1_n99 ) );
  NAND2_X1 u0_u3_u1_U58 (.A1( u0_u3_u1_n105 ) , .ZN( u0_u3_u1_n155 ) , .A2( u0_u3_u1_n95 ) );
  OAI21_X1 u0_u3_u1_U59 (.ZN( u0_u3_u1_n109 ) , .B1( u0_u3_u1_n129 ) , .B2( u0_u3_u1_n160 ) , .A( u0_u3_u1_n167 ) );
  AOI22_X1 u0_u3_u1_U6 (.B2( u0_u3_u1_n113 ) , .A2( u0_u3_u1_n114 ) , .ZN( u0_u3_u1_n125 ) , .A1( u0_u3_u1_n171 ) , .B1( u0_u3_u1_n173 ) );
  NAND2_X1 u0_u3_u1_U60 (.A2( u0_u3_u1_n100 ) , .A1( u0_u3_u1_n103 ) , .ZN( u0_u3_u1_n120 ) );
  NAND2_X1 u0_u3_u1_U61 (.A1( u0_u3_u1_n102 ) , .A2( u0_u3_u1_n104 ) , .ZN( u0_u3_u1_n115 ) );
  NAND2_X1 u0_u3_u1_U62 (.A2( u0_u3_u1_n100 ) , .A1( u0_u3_u1_n104 ) , .ZN( u0_u3_u1_n151 ) );
  NAND2_X1 u0_u3_u1_U63 (.A2( u0_u3_u1_n103 ) , .A1( u0_u3_u1_n105 ) , .ZN( u0_u3_u1_n161 ) );
  INV_X1 u0_u3_u1_U64 (.A( u0_u3_u1_n152 ) , .ZN( u0_u3_u1_n173 ) );
  INV_X1 u0_u3_u1_U65 (.A( u0_u3_u1_n128 ) , .ZN( u0_u3_u1_n172 ) );
  NAND2_X1 u0_u3_u1_U66 (.A2( u0_u3_u1_n102 ) , .A1( u0_u3_u1_n103 ) , .ZN( u0_u3_u1_n123 ) );
  AOI211_X1 u0_u3_u1_U67 (.B( u0_u3_u1_n162 ) , .A( u0_u3_u1_n163 ) , .C2( u0_u3_u1_n164 ) , .ZN( u0_u3_u1_n165 ) , .C1( u0_u3_u1_n171 ) );
  AOI21_X1 u0_u3_u1_U68 (.A( u0_u3_u1_n160 ) , .B2( u0_u3_u1_n161 ) , .ZN( u0_u3_u1_n162 ) , .B1( u0_u3_u1_n182 ) );
  OR2_X1 u0_u3_u1_U69 (.A2( u0_u3_u1_n157 ) , .A1( u0_u3_u1_n158 ) , .ZN( u0_u3_u1_n163 ) );
  NAND2_X1 u0_u3_u1_U7 (.ZN( u0_u3_u1_n114 ) , .A1( u0_u3_u1_n134 ) , .A2( u0_u3_u1_n156 ) );
  NOR2_X1 u0_u3_u1_U70 (.A2( u0_u3_X_7 ) , .A1( u0_u3_X_8 ) , .ZN( u0_u3_u1_n95 ) );
  NOR2_X1 u0_u3_u1_U71 (.A1( u0_u3_X_12 ) , .A2( u0_u3_X_9 ) , .ZN( u0_u3_u1_n100 ) );
  NOR2_X1 u0_u3_u1_U72 (.A2( u0_u3_X_8 ) , .A1( u0_u3_u1_n177 ) , .ZN( u0_u3_u1_n99 ) );
  NOR2_X1 u0_u3_u1_U73 (.A2( u0_u3_X_12 ) , .ZN( u0_u3_u1_n102 ) , .A1( u0_u3_u1_n176 ) );
  NOR2_X1 u0_u3_u1_U74 (.A2( u0_u3_X_9 ) , .ZN( u0_u3_u1_n105 ) , .A1( u0_u3_u1_n168 ) );
  NAND2_X1 u0_u3_u1_U75 (.A1( u0_u3_X_10 ) , .ZN( u0_u3_u1_n160 ) , .A2( u0_u3_u1_n169 ) );
  NAND2_X1 u0_u3_u1_U76 (.A2( u0_u3_X_10 ) , .A1( u0_u3_X_11 ) , .ZN( u0_u3_u1_n152 ) );
  NAND2_X1 u0_u3_u1_U77 (.A1( u0_u3_X_11 ) , .ZN( u0_u3_u1_n128 ) , .A2( u0_u3_u1_n170 ) );
  AND2_X1 u0_u3_u1_U78 (.A2( u0_u3_X_7 ) , .A1( u0_u3_X_8 ) , .ZN( u0_u3_u1_n104 ) );
  AND2_X1 u0_u3_u1_U79 (.A1( u0_u3_X_8 ) , .ZN( u0_u3_u1_n103 ) , .A2( u0_u3_u1_n177 ) );
  AOI22_X1 u0_u3_u1_U8 (.B2( u0_u3_u1_n136 ) , .A2( u0_u3_u1_n137 ) , .ZN( u0_u3_u1_n143 ) , .A1( u0_u3_u1_n171 ) , .B1( u0_u3_u1_n173 ) );
  INV_X1 u0_u3_u1_U80 (.A( u0_u3_X_10 ) , .ZN( u0_u3_u1_n170 ) );
  INV_X1 u0_u3_u1_U81 (.A( u0_u3_X_9 ) , .ZN( u0_u3_u1_n176 ) );
  INV_X1 u0_u3_u1_U82 (.A( u0_u3_X_11 ) , .ZN( u0_u3_u1_n169 ) );
  INV_X1 u0_u3_u1_U83 (.A( u0_u3_X_12 ) , .ZN( u0_u3_u1_n168 ) );
  INV_X1 u0_u3_u1_U84 (.A( u0_u3_X_7 ) , .ZN( u0_u3_u1_n177 ) );
  NAND4_X1 u0_u3_u1_U85 (.ZN( u0_out3_28 ) , .A4( u0_u3_u1_n124 ) , .A3( u0_u3_u1_n125 ) , .A2( u0_u3_u1_n126 ) , .A1( u0_u3_u1_n127 ) );
  OAI21_X1 u0_u3_u1_U86 (.ZN( u0_u3_u1_n127 ) , .B2( u0_u3_u1_n139 ) , .B1( u0_u3_u1_n175 ) , .A( u0_u3_u1_n183 ) );
  OAI21_X1 u0_u3_u1_U87 (.ZN( u0_u3_u1_n126 ) , .B2( u0_u3_u1_n140 ) , .A( u0_u3_u1_n146 ) , .B1( u0_u3_u1_n178 ) );
  NAND4_X1 u0_u3_u1_U88 (.ZN( u0_out3_18 ) , .A4( u0_u3_u1_n165 ) , .A3( u0_u3_u1_n166 ) , .A1( u0_u3_u1_n167 ) , .A2( u0_u3_u1_n186 ) );
  AOI22_X1 u0_u3_u1_U89 (.B2( u0_u3_u1_n146 ) , .B1( u0_u3_u1_n147 ) , .A2( u0_u3_u1_n148 ) , .ZN( u0_u3_u1_n166 ) , .A1( u0_u3_u1_n172 ) );
  INV_X1 u0_u3_u1_U9 (.A( u0_u3_u1_n147 ) , .ZN( u0_u3_u1_n181 ) );
  INV_X1 u0_u3_u1_U90 (.A( u0_u3_u1_n145 ) , .ZN( u0_u3_u1_n186 ) );
  NAND4_X1 u0_u3_u1_U91 (.ZN( u0_out3_2 ) , .A4( u0_u3_u1_n142 ) , .A3( u0_u3_u1_n143 ) , .A2( u0_u3_u1_n144 ) , .A1( u0_u3_u1_n179 ) );
  INV_X1 u0_u3_u1_U92 (.A( u0_u3_u1_n130 ) , .ZN( u0_u3_u1_n179 ) );
  OAI21_X1 u0_u3_u1_U93 (.B2( u0_u3_u1_n132 ) , .ZN( u0_u3_u1_n144 ) , .A( u0_u3_u1_n146 ) , .B1( u0_u3_u1_n180 ) );
  OR4_X1 u0_u3_u1_U94 (.ZN( u0_out3_13 ) , .A4( u0_u3_u1_n108 ) , .A3( u0_u3_u1_n109 ) , .A2( u0_u3_u1_n110 ) , .A1( u0_u3_u1_n111 ) );
  AOI21_X1 u0_u3_u1_U95 (.ZN( u0_u3_u1_n111 ) , .A( u0_u3_u1_n128 ) , .B2( u0_u3_u1_n131 ) , .B1( u0_u3_u1_n135 ) );
  AOI21_X1 u0_u3_u1_U96 (.ZN( u0_u3_u1_n110 ) , .A( u0_u3_u1_n116 ) , .B1( u0_u3_u1_n152 ) , .B2( u0_u3_u1_n160 ) );
  NAND3_X1 u0_u3_u1_U97 (.A3( u0_u3_u1_n149 ) , .A2( u0_u3_u1_n150 ) , .A1( u0_u3_u1_n151 ) , .ZN( u0_u3_u1_n164 ) );
  NAND3_X1 u0_u3_u1_U98 (.A3( u0_u3_u1_n134 ) , .A2( u0_u3_u1_n135 ) , .ZN( u0_u3_u1_n136 ) , .A1( u0_u3_u1_n151 ) );
  NAND3_X1 u0_u3_u1_U99 (.A1( u0_u3_u1_n133 ) , .ZN( u0_u3_u1_n137 ) , .A2( u0_u3_u1_n154 ) , .A3( u0_u3_u1_n181 ) );
  OAI22_X1 u0_u3_u2_U10 (.B1( u0_u3_u2_n151 ) , .A2( u0_u3_u2_n152 ) , .A1( u0_u3_u2_n153 ) , .ZN( u0_u3_u2_n160 ) , .B2( u0_u3_u2_n168 ) );
  NAND3_X1 u0_u3_u2_U100 (.A2( u0_u3_u2_n100 ) , .A1( u0_u3_u2_n104 ) , .A3( u0_u3_u2_n138 ) , .ZN( u0_u3_u2_n98 ) );
  NOR3_X1 u0_u3_u2_U11 (.A1( u0_u3_u2_n150 ) , .ZN( u0_u3_u2_n151 ) , .A3( u0_u3_u2_n175 ) , .A2( u0_u3_u2_n188 ) );
  AOI21_X1 u0_u3_u2_U12 (.B2( u0_u3_u2_n123 ) , .ZN( u0_u3_u2_n125 ) , .A( u0_u3_u2_n171 ) , .B1( u0_u3_u2_n184 ) );
  INV_X1 u0_u3_u2_U13 (.A( u0_u3_u2_n150 ) , .ZN( u0_u3_u2_n184 ) );
  AOI21_X1 u0_u3_u2_U14 (.ZN( u0_u3_u2_n144 ) , .B2( u0_u3_u2_n155 ) , .A( u0_u3_u2_n172 ) , .B1( u0_u3_u2_n185 ) );
  AOI21_X1 u0_u3_u2_U15 (.B2( u0_u3_u2_n143 ) , .ZN( u0_u3_u2_n145 ) , .B1( u0_u3_u2_n152 ) , .A( u0_u3_u2_n171 ) );
  INV_X1 u0_u3_u2_U16 (.A( u0_u3_u2_n156 ) , .ZN( u0_u3_u2_n171 ) );
  INV_X1 u0_u3_u2_U17 (.A( u0_u3_u2_n120 ) , .ZN( u0_u3_u2_n188 ) );
  NAND2_X1 u0_u3_u2_U18 (.A2( u0_u3_u2_n122 ) , .ZN( u0_u3_u2_n150 ) , .A1( u0_u3_u2_n152 ) );
  INV_X1 u0_u3_u2_U19 (.A( u0_u3_u2_n153 ) , .ZN( u0_u3_u2_n170 ) );
  INV_X1 u0_u3_u2_U20 (.A( u0_u3_u2_n137 ) , .ZN( u0_u3_u2_n173 ) );
  NAND2_X1 u0_u3_u2_U21 (.A1( u0_u3_u2_n132 ) , .A2( u0_u3_u2_n139 ) , .ZN( u0_u3_u2_n157 ) );
  INV_X1 u0_u3_u2_U22 (.A( u0_u3_u2_n113 ) , .ZN( u0_u3_u2_n178 ) );
  INV_X1 u0_u3_u2_U23 (.A( u0_u3_u2_n139 ) , .ZN( u0_u3_u2_n175 ) );
  INV_X1 u0_u3_u2_U24 (.A( u0_u3_u2_n155 ) , .ZN( u0_u3_u2_n181 ) );
  INV_X1 u0_u3_u2_U25 (.A( u0_u3_u2_n119 ) , .ZN( u0_u3_u2_n177 ) );
  INV_X1 u0_u3_u2_U26 (.A( u0_u3_u2_n116 ) , .ZN( u0_u3_u2_n180 ) );
  INV_X1 u0_u3_u2_U27 (.A( u0_u3_u2_n131 ) , .ZN( u0_u3_u2_n179 ) );
  INV_X1 u0_u3_u2_U28 (.A( u0_u3_u2_n154 ) , .ZN( u0_u3_u2_n176 ) );
  NAND2_X1 u0_u3_u2_U29 (.A2( u0_u3_u2_n116 ) , .A1( u0_u3_u2_n117 ) , .ZN( u0_u3_u2_n118 ) );
  NOR2_X1 u0_u3_u2_U3 (.ZN( u0_u3_u2_n121 ) , .A2( u0_u3_u2_n177 ) , .A1( u0_u3_u2_n180 ) );
  INV_X1 u0_u3_u2_U30 (.A( u0_u3_u2_n132 ) , .ZN( u0_u3_u2_n182 ) );
  INV_X1 u0_u3_u2_U31 (.A( u0_u3_u2_n158 ) , .ZN( u0_u3_u2_n183 ) );
  OAI21_X1 u0_u3_u2_U32 (.A( u0_u3_u2_n156 ) , .B1( u0_u3_u2_n157 ) , .ZN( u0_u3_u2_n158 ) , .B2( u0_u3_u2_n179 ) );
  NOR2_X1 u0_u3_u2_U33 (.ZN( u0_u3_u2_n156 ) , .A1( u0_u3_u2_n166 ) , .A2( u0_u3_u2_n169 ) );
  NOR2_X1 u0_u3_u2_U34 (.A2( u0_u3_u2_n114 ) , .ZN( u0_u3_u2_n137 ) , .A1( u0_u3_u2_n140 ) );
  NOR2_X1 u0_u3_u2_U35 (.A2( u0_u3_u2_n138 ) , .ZN( u0_u3_u2_n153 ) , .A1( u0_u3_u2_n156 ) );
  AOI211_X1 u0_u3_u2_U36 (.ZN( u0_u3_u2_n130 ) , .C1( u0_u3_u2_n138 ) , .C2( u0_u3_u2_n179 ) , .B( u0_u3_u2_n96 ) , .A( u0_u3_u2_n97 ) );
  OAI22_X1 u0_u3_u2_U37 (.B1( u0_u3_u2_n133 ) , .A2( u0_u3_u2_n137 ) , .A1( u0_u3_u2_n152 ) , .B2( u0_u3_u2_n168 ) , .ZN( u0_u3_u2_n97 ) );
  OAI221_X1 u0_u3_u2_U38 (.B1( u0_u3_u2_n113 ) , .C1( u0_u3_u2_n132 ) , .A( u0_u3_u2_n149 ) , .B2( u0_u3_u2_n171 ) , .C2( u0_u3_u2_n172 ) , .ZN( u0_u3_u2_n96 ) );
  OAI221_X1 u0_u3_u2_U39 (.A( u0_u3_u2_n115 ) , .C2( u0_u3_u2_n123 ) , .B2( u0_u3_u2_n143 ) , .B1( u0_u3_u2_n153 ) , .ZN( u0_u3_u2_n163 ) , .C1( u0_u3_u2_n168 ) );
  INV_X1 u0_u3_u2_U4 (.A( u0_u3_u2_n134 ) , .ZN( u0_u3_u2_n185 ) );
  OAI21_X1 u0_u3_u2_U40 (.A( u0_u3_u2_n114 ) , .ZN( u0_u3_u2_n115 ) , .B1( u0_u3_u2_n176 ) , .B2( u0_u3_u2_n178 ) );
  OAI221_X1 u0_u3_u2_U41 (.A( u0_u3_u2_n135 ) , .B2( u0_u3_u2_n136 ) , .B1( u0_u3_u2_n137 ) , .ZN( u0_u3_u2_n162 ) , .C2( u0_u3_u2_n167 ) , .C1( u0_u3_u2_n185 ) );
  AND3_X1 u0_u3_u2_U42 (.A3( u0_u3_u2_n131 ) , .A2( u0_u3_u2_n132 ) , .A1( u0_u3_u2_n133 ) , .ZN( u0_u3_u2_n136 ) );
  AOI22_X1 u0_u3_u2_U43 (.ZN( u0_u3_u2_n135 ) , .B1( u0_u3_u2_n140 ) , .A1( u0_u3_u2_n156 ) , .B2( u0_u3_u2_n180 ) , .A2( u0_u3_u2_n188 ) );
  AOI21_X1 u0_u3_u2_U44 (.ZN( u0_u3_u2_n149 ) , .B1( u0_u3_u2_n173 ) , .B2( u0_u3_u2_n188 ) , .A( u0_u3_u2_n95 ) );
  AND3_X1 u0_u3_u2_U45 (.A2( u0_u3_u2_n100 ) , .A1( u0_u3_u2_n104 ) , .A3( u0_u3_u2_n156 ) , .ZN( u0_u3_u2_n95 ) );
  OAI21_X1 u0_u3_u2_U46 (.A( u0_u3_u2_n141 ) , .B2( u0_u3_u2_n142 ) , .ZN( u0_u3_u2_n146 ) , .B1( u0_u3_u2_n153 ) );
  OAI21_X1 u0_u3_u2_U47 (.A( u0_u3_u2_n140 ) , .ZN( u0_u3_u2_n141 ) , .B1( u0_u3_u2_n176 ) , .B2( u0_u3_u2_n177 ) );
  NOR3_X1 u0_u3_u2_U48 (.ZN( u0_u3_u2_n142 ) , .A3( u0_u3_u2_n175 ) , .A2( u0_u3_u2_n178 ) , .A1( u0_u3_u2_n181 ) );
  OAI21_X1 u0_u3_u2_U49 (.A( u0_u3_u2_n101 ) , .B2( u0_u3_u2_n121 ) , .B1( u0_u3_u2_n153 ) , .ZN( u0_u3_u2_n164 ) );
  NOR4_X1 u0_u3_u2_U5 (.A4( u0_u3_u2_n124 ) , .A3( u0_u3_u2_n125 ) , .A2( u0_u3_u2_n126 ) , .A1( u0_u3_u2_n127 ) , .ZN( u0_u3_u2_n128 ) );
  NAND2_X1 u0_u3_u2_U50 (.A2( u0_u3_u2_n100 ) , .A1( u0_u3_u2_n107 ) , .ZN( u0_u3_u2_n155 ) );
  NAND2_X1 u0_u3_u2_U51 (.A2( u0_u3_u2_n105 ) , .A1( u0_u3_u2_n108 ) , .ZN( u0_u3_u2_n143 ) );
  NAND2_X1 u0_u3_u2_U52 (.A1( u0_u3_u2_n104 ) , .A2( u0_u3_u2_n106 ) , .ZN( u0_u3_u2_n152 ) );
  NAND2_X1 u0_u3_u2_U53 (.A1( u0_u3_u2_n100 ) , .A2( u0_u3_u2_n105 ) , .ZN( u0_u3_u2_n132 ) );
  INV_X1 u0_u3_u2_U54 (.A( u0_u3_u2_n140 ) , .ZN( u0_u3_u2_n168 ) );
  INV_X1 u0_u3_u2_U55 (.A( u0_u3_u2_n138 ) , .ZN( u0_u3_u2_n167 ) );
  INV_X1 u0_u3_u2_U56 (.ZN( u0_u3_u2_n187 ) , .A( u0_u3_u2_n99 ) );
  OAI21_X1 u0_u3_u2_U57 (.B1( u0_u3_u2_n137 ) , .B2( u0_u3_u2_n143 ) , .A( u0_u3_u2_n98 ) , .ZN( u0_u3_u2_n99 ) );
  NAND2_X1 u0_u3_u2_U58 (.A1( u0_u3_u2_n102 ) , .A2( u0_u3_u2_n106 ) , .ZN( u0_u3_u2_n113 ) );
  NAND2_X1 u0_u3_u2_U59 (.A1( u0_u3_u2_n106 ) , .A2( u0_u3_u2_n107 ) , .ZN( u0_u3_u2_n131 ) );
  AOI21_X1 u0_u3_u2_U6 (.B2( u0_u3_u2_n119 ) , .ZN( u0_u3_u2_n127 ) , .A( u0_u3_u2_n137 ) , .B1( u0_u3_u2_n155 ) );
  NAND2_X1 u0_u3_u2_U60 (.A1( u0_u3_u2_n103 ) , .A2( u0_u3_u2_n107 ) , .ZN( u0_u3_u2_n139 ) );
  NAND2_X1 u0_u3_u2_U61 (.A1( u0_u3_u2_n103 ) , .A2( u0_u3_u2_n105 ) , .ZN( u0_u3_u2_n133 ) );
  NAND2_X1 u0_u3_u2_U62 (.A1( u0_u3_u2_n102 ) , .A2( u0_u3_u2_n103 ) , .ZN( u0_u3_u2_n154 ) );
  NAND2_X1 u0_u3_u2_U63 (.A2( u0_u3_u2_n103 ) , .A1( u0_u3_u2_n104 ) , .ZN( u0_u3_u2_n119 ) );
  NAND2_X1 u0_u3_u2_U64 (.A2( u0_u3_u2_n107 ) , .A1( u0_u3_u2_n108 ) , .ZN( u0_u3_u2_n123 ) );
  NAND2_X1 u0_u3_u2_U65 (.A1( u0_u3_u2_n104 ) , .A2( u0_u3_u2_n108 ) , .ZN( u0_u3_u2_n122 ) );
  INV_X1 u0_u3_u2_U66 (.A( u0_u3_u2_n114 ) , .ZN( u0_u3_u2_n172 ) );
  NAND2_X1 u0_u3_u2_U67 (.A2( u0_u3_u2_n100 ) , .A1( u0_u3_u2_n102 ) , .ZN( u0_u3_u2_n116 ) );
  NAND2_X1 u0_u3_u2_U68 (.A1( u0_u3_u2_n102 ) , .A2( u0_u3_u2_n108 ) , .ZN( u0_u3_u2_n120 ) );
  NAND2_X1 u0_u3_u2_U69 (.A2( u0_u3_u2_n105 ) , .A1( u0_u3_u2_n106 ) , .ZN( u0_u3_u2_n117 ) );
  AOI21_X1 u0_u3_u2_U7 (.ZN( u0_u3_u2_n124 ) , .B1( u0_u3_u2_n131 ) , .B2( u0_u3_u2_n143 ) , .A( u0_u3_u2_n172 ) );
  NOR2_X1 u0_u3_u2_U70 (.A2( u0_u3_X_16 ) , .ZN( u0_u3_u2_n140 ) , .A1( u0_u3_u2_n166 ) );
  NOR2_X1 u0_u3_u2_U71 (.A2( u0_u3_X_13 ) , .A1( u0_u3_X_14 ) , .ZN( u0_u3_u2_n100 ) );
  NOR2_X1 u0_u3_u2_U72 (.A2( u0_u3_X_16 ) , .A1( u0_u3_X_17 ) , .ZN( u0_u3_u2_n138 ) );
  NOR2_X1 u0_u3_u2_U73 (.A2( u0_u3_X_15 ) , .A1( u0_u3_X_18 ) , .ZN( u0_u3_u2_n104 ) );
  NOR2_X1 u0_u3_u2_U74 (.A2( u0_u3_X_14 ) , .ZN( u0_u3_u2_n103 ) , .A1( u0_u3_u2_n174 ) );
  NOR2_X1 u0_u3_u2_U75 (.A2( u0_u3_X_15 ) , .ZN( u0_u3_u2_n102 ) , .A1( u0_u3_u2_n165 ) );
  NOR2_X1 u0_u3_u2_U76 (.A2( u0_u3_X_17 ) , .ZN( u0_u3_u2_n114 ) , .A1( u0_u3_u2_n169 ) );
  AND2_X1 u0_u3_u2_U77 (.A1( u0_u3_X_15 ) , .ZN( u0_u3_u2_n105 ) , .A2( u0_u3_u2_n165 ) );
  AND2_X1 u0_u3_u2_U78 (.A2( u0_u3_X_15 ) , .A1( u0_u3_X_18 ) , .ZN( u0_u3_u2_n107 ) );
  AND2_X1 u0_u3_u2_U79 (.A1( u0_u3_X_14 ) , .ZN( u0_u3_u2_n106 ) , .A2( u0_u3_u2_n174 ) );
  AOI21_X1 u0_u3_u2_U8 (.B2( u0_u3_u2_n120 ) , .B1( u0_u3_u2_n121 ) , .ZN( u0_u3_u2_n126 ) , .A( u0_u3_u2_n167 ) );
  AND2_X1 u0_u3_u2_U80 (.A1( u0_u3_X_13 ) , .A2( u0_u3_X_14 ) , .ZN( u0_u3_u2_n108 ) );
  INV_X1 u0_u3_u2_U81 (.A( u0_u3_X_16 ) , .ZN( u0_u3_u2_n169 ) );
  INV_X1 u0_u3_u2_U82 (.A( u0_u3_X_17 ) , .ZN( u0_u3_u2_n166 ) );
  INV_X1 u0_u3_u2_U83 (.A( u0_u3_X_13 ) , .ZN( u0_u3_u2_n174 ) );
  INV_X1 u0_u3_u2_U84 (.A( u0_u3_X_18 ) , .ZN( u0_u3_u2_n165 ) );
  NAND4_X1 u0_u3_u2_U85 (.ZN( u0_out3_24 ) , .A4( u0_u3_u2_n111 ) , .A3( u0_u3_u2_n112 ) , .A1( u0_u3_u2_n130 ) , .A2( u0_u3_u2_n187 ) );
  AOI221_X1 u0_u3_u2_U86 (.A( u0_u3_u2_n109 ) , .B1( u0_u3_u2_n110 ) , .ZN( u0_u3_u2_n111 ) , .C1( u0_u3_u2_n134 ) , .C2( u0_u3_u2_n170 ) , .B2( u0_u3_u2_n173 ) );
  AOI21_X1 u0_u3_u2_U87 (.ZN( u0_u3_u2_n112 ) , .B2( u0_u3_u2_n156 ) , .A( u0_u3_u2_n164 ) , .B1( u0_u3_u2_n181 ) );
  NAND4_X1 u0_u3_u2_U88 (.ZN( u0_out3_16 ) , .A4( u0_u3_u2_n128 ) , .A3( u0_u3_u2_n129 ) , .A1( u0_u3_u2_n130 ) , .A2( u0_u3_u2_n186 ) );
  AOI22_X1 u0_u3_u2_U89 (.A2( u0_u3_u2_n118 ) , .ZN( u0_u3_u2_n129 ) , .A1( u0_u3_u2_n140 ) , .B1( u0_u3_u2_n157 ) , .B2( u0_u3_u2_n170 ) );
  OAI22_X1 u0_u3_u2_U9 (.ZN( u0_u3_u2_n109 ) , .A2( u0_u3_u2_n113 ) , .B2( u0_u3_u2_n133 ) , .B1( u0_u3_u2_n167 ) , .A1( u0_u3_u2_n168 ) );
  INV_X1 u0_u3_u2_U90 (.A( u0_u3_u2_n163 ) , .ZN( u0_u3_u2_n186 ) );
  NAND4_X1 u0_u3_u2_U91 (.ZN( u0_out3_30 ) , .A4( u0_u3_u2_n147 ) , .A3( u0_u3_u2_n148 ) , .A2( u0_u3_u2_n149 ) , .A1( u0_u3_u2_n187 ) );
  AOI21_X1 u0_u3_u2_U92 (.B2( u0_u3_u2_n138 ) , .ZN( u0_u3_u2_n148 ) , .A( u0_u3_u2_n162 ) , .B1( u0_u3_u2_n182 ) );
  NOR3_X1 u0_u3_u2_U93 (.A3( u0_u3_u2_n144 ) , .A2( u0_u3_u2_n145 ) , .A1( u0_u3_u2_n146 ) , .ZN( u0_u3_u2_n147 ) );
  OR4_X1 u0_u3_u2_U94 (.ZN( u0_out3_6 ) , .A4( u0_u3_u2_n161 ) , .A3( u0_u3_u2_n162 ) , .A2( u0_u3_u2_n163 ) , .A1( u0_u3_u2_n164 ) );
  OR3_X1 u0_u3_u2_U95 (.A2( u0_u3_u2_n159 ) , .A1( u0_u3_u2_n160 ) , .ZN( u0_u3_u2_n161 ) , .A3( u0_u3_u2_n183 ) );
  AOI21_X1 u0_u3_u2_U96 (.B2( u0_u3_u2_n154 ) , .B1( u0_u3_u2_n155 ) , .ZN( u0_u3_u2_n159 ) , .A( u0_u3_u2_n167 ) );
  NAND3_X1 u0_u3_u2_U97 (.A2( u0_u3_u2_n117 ) , .A1( u0_u3_u2_n122 ) , .A3( u0_u3_u2_n123 ) , .ZN( u0_u3_u2_n134 ) );
  NAND3_X1 u0_u3_u2_U98 (.ZN( u0_u3_u2_n110 ) , .A2( u0_u3_u2_n131 ) , .A3( u0_u3_u2_n139 ) , .A1( u0_u3_u2_n154 ) );
  NAND3_X1 u0_u3_u2_U99 (.A2( u0_u3_u2_n100 ) , .ZN( u0_u3_u2_n101 ) , .A1( u0_u3_u2_n104 ) , .A3( u0_u3_u2_n114 ) );
  OAI22_X1 u0_u3_u3_U10 (.B1( u0_u3_u3_n113 ) , .A2( u0_u3_u3_n135 ) , .A1( u0_u3_u3_n150 ) , .B2( u0_u3_u3_n164 ) , .ZN( u0_u3_u3_n98 ) );
  OAI211_X1 u0_u3_u3_U11 (.B( u0_u3_u3_n106 ) , .ZN( u0_u3_u3_n119 ) , .C2( u0_u3_u3_n128 ) , .C1( u0_u3_u3_n167 ) , .A( u0_u3_u3_n181 ) );
  AOI221_X1 u0_u3_u3_U12 (.C1( u0_u3_u3_n105 ) , .ZN( u0_u3_u3_n106 ) , .A( u0_u3_u3_n131 ) , .B2( u0_u3_u3_n132 ) , .C2( u0_u3_u3_n133 ) , .B1( u0_u3_u3_n169 ) );
  INV_X1 u0_u3_u3_U13 (.ZN( u0_u3_u3_n181 ) , .A( u0_u3_u3_n98 ) );
  NAND2_X1 u0_u3_u3_U14 (.ZN( u0_u3_u3_n105 ) , .A2( u0_u3_u3_n130 ) , .A1( u0_u3_u3_n155 ) );
  AOI22_X1 u0_u3_u3_U15 (.B1( u0_u3_u3_n115 ) , .A2( u0_u3_u3_n116 ) , .ZN( u0_u3_u3_n123 ) , .B2( u0_u3_u3_n133 ) , .A1( u0_u3_u3_n169 ) );
  NAND2_X1 u0_u3_u3_U16 (.ZN( u0_u3_u3_n116 ) , .A2( u0_u3_u3_n151 ) , .A1( u0_u3_u3_n182 ) );
  NOR2_X1 u0_u3_u3_U17 (.ZN( u0_u3_u3_n126 ) , .A2( u0_u3_u3_n150 ) , .A1( u0_u3_u3_n164 ) );
  AOI21_X1 u0_u3_u3_U18 (.ZN( u0_u3_u3_n112 ) , .B2( u0_u3_u3_n146 ) , .B1( u0_u3_u3_n155 ) , .A( u0_u3_u3_n167 ) );
  NAND2_X1 u0_u3_u3_U19 (.A1( u0_u3_u3_n135 ) , .ZN( u0_u3_u3_n142 ) , .A2( u0_u3_u3_n164 ) );
  NAND2_X1 u0_u3_u3_U20 (.ZN( u0_u3_u3_n132 ) , .A2( u0_u3_u3_n152 ) , .A1( u0_u3_u3_n156 ) );
  INV_X1 u0_u3_u3_U21 (.A( u0_u3_u3_n133 ) , .ZN( u0_u3_u3_n165 ) );
  NAND2_X1 u0_u3_u3_U22 (.ZN( u0_u3_u3_n143 ) , .A1( u0_u3_u3_n165 ) , .A2( u0_u3_u3_n167 ) );
  AND2_X1 u0_u3_u3_U23 (.A2( u0_u3_u3_n113 ) , .A1( u0_u3_u3_n114 ) , .ZN( u0_u3_u3_n151 ) );
  INV_X1 u0_u3_u3_U24 (.A( u0_u3_u3_n135 ) , .ZN( u0_u3_u3_n170 ) );
  NAND2_X1 u0_u3_u3_U25 (.A1( u0_u3_u3_n107 ) , .A2( u0_u3_u3_n108 ) , .ZN( u0_u3_u3_n140 ) );
  NAND2_X1 u0_u3_u3_U26 (.ZN( u0_u3_u3_n117 ) , .A1( u0_u3_u3_n124 ) , .A2( u0_u3_u3_n148 ) );
  INV_X1 u0_u3_u3_U27 (.A( u0_u3_u3_n130 ) , .ZN( u0_u3_u3_n177 ) );
  INV_X1 u0_u3_u3_U28 (.A( u0_u3_u3_n128 ) , .ZN( u0_u3_u3_n176 ) );
  INV_X1 u0_u3_u3_U29 (.A( u0_u3_u3_n155 ) , .ZN( u0_u3_u3_n174 ) );
  INV_X1 u0_u3_u3_U3 (.A( u0_u3_u3_n140 ) , .ZN( u0_u3_u3_n182 ) );
  INV_X1 u0_u3_u3_U30 (.A( u0_u3_u3_n139 ) , .ZN( u0_u3_u3_n185 ) );
  NOR2_X1 u0_u3_u3_U31 (.ZN( u0_u3_u3_n135 ) , .A2( u0_u3_u3_n141 ) , .A1( u0_u3_u3_n169 ) );
  INV_X1 u0_u3_u3_U32 (.A( u0_u3_u3_n156 ) , .ZN( u0_u3_u3_n179 ) );
  OAI22_X1 u0_u3_u3_U33 (.B1( u0_u3_u3_n118 ) , .ZN( u0_u3_u3_n120 ) , .A1( u0_u3_u3_n135 ) , .B2( u0_u3_u3_n154 ) , .A2( u0_u3_u3_n178 ) );
  AND3_X1 u0_u3_u3_U34 (.ZN( u0_u3_u3_n118 ) , .A2( u0_u3_u3_n124 ) , .A1( u0_u3_u3_n144 ) , .A3( u0_u3_u3_n152 ) );
  OAI222_X1 u0_u3_u3_U35 (.C2( u0_u3_u3_n107 ) , .A2( u0_u3_u3_n108 ) , .B1( u0_u3_u3_n135 ) , .ZN( u0_u3_u3_n138 ) , .B2( u0_u3_u3_n146 ) , .C1( u0_u3_u3_n154 ) , .A1( u0_u3_u3_n164 ) );
  NOR4_X1 u0_u3_u3_U36 (.A4( u0_u3_u3_n157 ) , .A3( u0_u3_u3_n158 ) , .A2( u0_u3_u3_n159 ) , .A1( u0_u3_u3_n160 ) , .ZN( u0_u3_u3_n161 ) );
  AOI21_X1 u0_u3_u3_U37 (.B2( u0_u3_u3_n152 ) , .B1( u0_u3_u3_n153 ) , .ZN( u0_u3_u3_n158 ) , .A( u0_u3_u3_n164 ) );
  AOI21_X1 u0_u3_u3_U38 (.A( u0_u3_u3_n149 ) , .B2( u0_u3_u3_n150 ) , .B1( u0_u3_u3_n151 ) , .ZN( u0_u3_u3_n159 ) );
  AOI21_X1 u0_u3_u3_U39 (.A( u0_u3_u3_n154 ) , .B2( u0_u3_u3_n155 ) , .B1( u0_u3_u3_n156 ) , .ZN( u0_u3_u3_n157 ) );
  INV_X1 u0_u3_u3_U4 (.A( u0_u3_u3_n129 ) , .ZN( u0_u3_u3_n183 ) );
  AOI211_X1 u0_u3_u3_U40 (.ZN( u0_u3_u3_n109 ) , .A( u0_u3_u3_n119 ) , .C2( u0_u3_u3_n129 ) , .B( u0_u3_u3_n138 ) , .C1( u0_u3_u3_n141 ) );
  INV_X1 u0_u3_u3_U41 (.A( u0_u3_u3_n121 ) , .ZN( u0_u3_u3_n164 ) );
  NAND2_X1 u0_u3_u3_U42 (.ZN( u0_u3_u3_n133 ) , .A1( u0_u3_u3_n154 ) , .A2( u0_u3_u3_n164 ) );
  OAI211_X1 u0_u3_u3_U43 (.B( u0_u3_u3_n127 ) , .ZN( u0_u3_u3_n139 ) , .C1( u0_u3_u3_n150 ) , .C2( u0_u3_u3_n154 ) , .A( u0_u3_u3_n184 ) );
  INV_X1 u0_u3_u3_U44 (.A( u0_u3_u3_n125 ) , .ZN( u0_u3_u3_n184 ) );
  AOI221_X1 u0_u3_u3_U45 (.A( u0_u3_u3_n126 ) , .ZN( u0_u3_u3_n127 ) , .C2( u0_u3_u3_n132 ) , .C1( u0_u3_u3_n169 ) , .B2( u0_u3_u3_n170 ) , .B1( u0_u3_u3_n174 ) );
  OAI22_X1 u0_u3_u3_U46 (.A1( u0_u3_u3_n124 ) , .ZN( u0_u3_u3_n125 ) , .B2( u0_u3_u3_n145 ) , .A2( u0_u3_u3_n165 ) , .B1( u0_u3_u3_n167 ) );
  NOR2_X1 u0_u3_u3_U47 (.A1( u0_u3_u3_n113 ) , .ZN( u0_u3_u3_n131 ) , .A2( u0_u3_u3_n154 ) );
  NAND2_X1 u0_u3_u3_U48 (.A1( u0_u3_u3_n103 ) , .ZN( u0_u3_u3_n150 ) , .A2( u0_u3_u3_n99 ) );
  NAND2_X1 u0_u3_u3_U49 (.A2( u0_u3_u3_n102 ) , .ZN( u0_u3_u3_n155 ) , .A1( u0_u3_u3_n97 ) );
  INV_X1 u0_u3_u3_U5 (.A( u0_u3_u3_n117 ) , .ZN( u0_u3_u3_n178 ) );
  INV_X1 u0_u3_u3_U50 (.A( u0_u3_u3_n141 ) , .ZN( u0_u3_u3_n167 ) );
  AOI21_X1 u0_u3_u3_U51 (.B2( u0_u3_u3_n114 ) , .B1( u0_u3_u3_n146 ) , .A( u0_u3_u3_n154 ) , .ZN( u0_u3_u3_n94 ) );
  AOI21_X1 u0_u3_u3_U52 (.ZN( u0_u3_u3_n110 ) , .B2( u0_u3_u3_n142 ) , .B1( u0_u3_u3_n186 ) , .A( u0_u3_u3_n95 ) );
  INV_X1 u0_u3_u3_U53 (.A( u0_u3_u3_n145 ) , .ZN( u0_u3_u3_n186 ) );
  AOI21_X1 u0_u3_u3_U54 (.B1( u0_u3_u3_n124 ) , .A( u0_u3_u3_n149 ) , .B2( u0_u3_u3_n155 ) , .ZN( u0_u3_u3_n95 ) );
  INV_X1 u0_u3_u3_U55 (.A( u0_u3_u3_n149 ) , .ZN( u0_u3_u3_n169 ) );
  NAND2_X1 u0_u3_u3_U56 (.ZN( u0_u3_u3_n124 ) , .A1( u0_u3_u3_n96 ) , .A2( u0_u3_u3_n97 ) );
  NAND2_X1 u0_u3_u3_U57 (.A2( u0_u3_u3_n100 ) , .ZN( u0_u3_u3_n146 ) , .A1( u0_u3_u3_n96 ) );
  NAND2_X1 u0_u3_u3_U58 (.A1( u0_u3_u3_n101 ) , .ZN( u0_u3_u3_n145 ) , .A2( u0_u3_u3_n99 ) );
  NAND2_X1 u0_u3_u3_U59 (.A1( u0_u3_u3_n100 ) , .ZN( u0_u3_u3_n156 ) , .A2( u0_u3_u3_n99 ) );
  AOI221_X1 u0_u3_u3_U6 (.A( u0_u3_u3_n131 ) , .C2( u0_u3_u3_n132 ) , .C1( u0_u3_u3_n133 ) , .ZN( u0_u3_u3_n134 ) , .B1( u0_u3_u3_n143 ) , .B2( u0_u3_u3_n177 ) );
  NAND2_X1 u0_u3_u3_U60 (.A2( u0_u3_u3_n101 ) , .A1( u0_u3_u3_n104 ) , .ZN( u0_u3_u3_n148 ) );
  NAND2_X1 u0_u3_u3_U61 (.A1( u0_u3_u3_n100 ) , .A2( u0_u3_u3_n102 ) , .ZN( u0_u3_u3_n128 ) );
  NAND2_X1 u0_u3_u3_U62 (.A2( u0_u3_u3_n101 ) , .A1( u0_u3_u3_n102 ) , .ZN( u0_u3_u3_n152 ) );
  NAND2_X1 u0_u3_u3_U63 (.A2( u0_u3_u3_n101 ) , .ZN( u0_u3_u3_n114 ) , .A1( u0_u3_u3_n96 ) );
  NAND2_X1 u0_u3_u3_U64 (.ZN( u0_u3_u3_n107 ) , .A1( u0_u3_u3_n97 ) , .A2( u0_u3_u3_n99 ) );
  NAND2_X1 u0_u3_u3_U65 (.A2( u0_u3_u3_n100 ) , .A1( u0_u3_u3_n104 ) , .ZN( u0_u3_u3_n113 ) );
  NAND2_X1 u0_u3_u3_U66 (.A1( u0_u3_u3_n104 ) , .ZN( u0_u3_u3_n153 ) , .A2( u0_u3_u3_n97 ) );
  NAND2_X1 u0_u3_u3_U67 (.A2( u0_u3_u3_n103 ) , .A1( u0_u3_u3_n104 ) , .ZN( u0_u3_u3_n130 ) );
  NAND2_X1 u0_u3_u3_U68 (.A2( u0_u3_u3_n103 ) , .ZN( u0_u3_u3_n144 ) , .A1( u0_u3_u3_n96 ) );
  NAND2_X1 u0_u3_u3_U69 (.A1( u0_u3_u3_n102 ) , .A2( u0_u3_u3_n103 ) , .ZN( u0_u3_u3_n108 ) );
  OAI22_X1 u0_u3_u3_U7 (.B2( u0_u3_u3_n147 ) , .A2( u0_u3_u3_n148 ) , .ZN( u0_u3_u3_n160 ) , .B1( u0_u3_u3_n165 ) , .A1( u0_u3_u3_n168 ) );
  NOR2_X1 u0_u3_u3_U70 (.A2( u0_u3_X_19 ) , .A1( u0_u3_X_20 ) , .ZN( u0_u3_u3_n99 ) );
  NOR2_X1 u0_u3_u3_U71 (.A2( u0_u3_X_21 ) , .A1( u0_u3_X_24 ) , .ZN( u0_u3_u3_n103 ) );
  NOR2_X1 u0_u3_u3_U72 (.A2( u0_u3_X_24 ) , .A1( u0_u3_u3_n171 ) , .ZN( u0_u3_u3_n97 ) );
  NOR2_X1 u0_u3_u3_U73 (.A2( u0_u3_X_19 ) , .A1( u0_u3_u3_n172 ) , .ZN( u0_u3_u3_n96 ) );
  NAND2_X1 u0_u3_u3_U74 (.A1( u0_u3_X_22 ) , .A2( u0_u3_X_23 ) , .ZN( u0_u3_u3_n154 ) );
  AND2_X1 u0_u3_u3_U75 (.A1( u0_u3_X_24 ) , .ZN( u0_u3_u3_n101 ) , .A2( u0_u3_u3_n171 ) );
  AND2_X1 u0_u3_u3_U76 (.A1( u0_u3_X_19 ) , .ZN( u0_u3_u3_n102 ) , .A2( u0_u3_u3_n172 ) );
  AND2_X1 u0_u3_u3_U77 (.A1( u0_u3_X_21 ) , .A2( u0_u3_X_24 ) , .ZN( u0_u3_u3_n100 ) );
  AND2_X1 u0_u3_u3_U78 (.A2( u0_u3_X_19 ) , .A1( u0_u3_X_20 ) , .ZN( u0_u3_u3_n104 ) );
  INV_X1 u0_u3_u3_U79 (.A( u0_u3_X_21 ) , .ZN( u0_u3_u3_n171 ) );
  AND3_X1 u0_u3_u3_U8 (.A3( u0_u3_u3_n144 ) , .A2( u0_u3_u3_n145 ) , .A1( u0_u3_u3_n146 ) , .ZN( u0_u3_u3_n147 ) );
  INV_X1 u0_u3_u3_U80 (.A( u0_u3_X_20 ) , .ZN( u0_u3_u3_n172 ) );
  INV_X1 u0_u3_u3_U81 (.A( u0_u3_X_22 ) , .ZN( u0_u3_u3_n166 ) );
  NAND4_X1 u0_u3_u3_U82 (.ZN( u0_out3_26 ) , .A4( u0_u3_u3_n109 ) , .A3( u0_u3_u3_n110 ) , .A2( u0_u3_u3_n111 ) , .A1( u0_u3_u3_n173 ) );
  INV_X1 u0_u3_u3_U83 (.ZN( u0_u3_u3_n173 ) , .A( u0_u3_u3_n94 ) );
  OAI21_X1 u0_u3_u3_U84 (.ZN( u0_u3_u3_n111 ) , .B2( u0_u3_u3_n117 ) , .A( u0_u3_u3_n133 ) , .B1( u0_u3_u3_n176 ) );
  NAND4_X1 u0_u3_u3_U85 (.ZN( u0_out3_1 ) , .A4( u0_u3_u3_n161 ) , .A3( u0_u3_u3_n162 ) , .A2( u0_u3_u3_n163 ) , .A1( u0_u3_u3_n185 ) );
  NAND2_X1 u0_u3_u3_U86 (.ZN( u0_u3_u3_n163 ) , .A2( u0_u3_u3_n170 ) , .A1( u0_u3_u3_n176 ) );
  AOI22_X1 u0_u3_u3_U87 (.B2( u0_u3_u3_n140 ) , .B1( u0_u3_u3_n141 ) , .A2( u0_u3_u3_n142 ) , .ZN( u0_u3_u3_n162 ) , .A1( u0_u3_u3_n177 ) );
  NAND4_X1 u0_u3_u3_U88 (.ZN( u0_out3_20 ) , .A4( u0_u3_u3_n122 ) , .A3( u0_u3_u3_n123 ) , .A1( u0_u3_u3_n175 ) , .A2( u0_u3_u3_n180 ) );
  INV_X1 u0_u3_u3_U89 (.A( u0_u3_u3_n126 ) , .ZN( u0_u3_u3_n180 ) );
  INV_X1 u0_u3_u3_U9 (.A( u0_u3_u3_n143 ) , .ZN( u0_u3_u3_n168 ) );
  INV_X1 u0_u3_u3_U90 (.A( u0_u3_u3_n112 ) , .ZN( u0_u3_u3_n175 ) );
  OR4_X1 u0_u3_u3_U91 (.ZN( u0_out3_10 ) , .A4( u0_u3_u3_n136 ) , .A3( u0_u3_u3_n137 ) , .A1( u0_u3_u3_n138 ) , .A2( u0_u3_u3_n139 ) );
  OAI222_X1 u0_u3_u3_U92 (.C1( u0_u3_u3_n128 ) , .ZN( u0_u3_u3_n137 ) , .B1( u0_u3_u3_n148 ) , .A2( u0_u3_u3_n150 ) , .B2( u0_u3_u3_n154 ) , .C2( u0_u3_u3_n164 ) , .A1( u0_u3_u3_n167 ) );
  AOI211_X1 u0_u3_u3_U93 (.B( u0_u3_u3_n119 ) , .A( u0_u3_u3_n120 ) , .C2( u0_u3_u3_n121 ) , .ZN( u0_u3_u3_n122 ) , .C1( u0_u3_u3_n179 ) );
  OAI221_X1 u0_u3_u3_U94 (.A( u0_u3_u3_n134 ) , .B2( u0_u3_u3_n135 ) , .ZN( u0_u3_u3_n136 ) , .C1( u0_u3_u3_n149 ) , .B1( u0_u3_u3_n151 ) , .C2( u0_u3_u3_n183 ) );
  NOR2_X1 u0_u3_u3_U95 (.A2( u0_u3_X_23 ) , .ZN( u0_u3_u3_n141 ) , .A1( u0_u3_u3_n166 ) );
  NAND2_X1 u0_u3_u3_U96 (.A1( u0_u3_X_23 ) , .ZN( u0_u3_u3_n149 ) , .A2( u0_u3_u3_n166 ) );
  NOR2_X1 u0_u3_u3_U97 (.A2( u0_u3_X_22 ) , .A1( u0_u3_X_23 ) , .ZN( u0_u3_u3_n121 ) );
  NAND3_X1 u0_u3_u3_U98 (.A1( u0_u3_u3_n114 ) , .ZN( u0_u3_u3_n115 ) , .A2( u0_u3_u3_n145 ) , .A3( u0_u3_u3_n153 ) );
  NAND3_X1 u0_u3_u3_U99 (.ZN( u0_u3_u3_n129 ) , .A2( u0_u3_u3_n144 ) , .A1( u0_u3_u3_n153 ) , .A3( u0_u3_u3_n182 ) );
  OAI22_X1 u0_u3_u4_U10 (.B2( u0_u3_u4_n135 ) , .ZN( u0_u3_u4_n137 ) , .B1( u0_u3_u4_n153 ) , .A1( u0_u3_u4_n155 ) , .A2( u0_u3_u4_n171 ) );
  AND3_X1 u0_u3_u4_U11 (.A2( u0_u3_u4_n134 ) , .ZN( u0_u3_u4_n135 ) , .A3( u0_u3_u4_n145 ) , .A1( u0_u3_u4_n157 ) );
  OR3_X1 u0_u3_u4_U12 (.A3( u0_u3_u4_n114 ) , .A2( u0_u3_u4_n115 ) , .A1( u0_u3_u4_n116 ) , .ZN( u0_u3_u4_n136 ) );
  AOI21_X1 u0_u3_u4_U13 (.A( u0_u3_u4_n113 ) , .ZN( u0_u3_u4_n116 ) , .B2( u0_u3_u4_n173 ) , .B1( u0_u3_u4_n174 ) );
  AOI21_X1 u0_u3_u4_U14 (.ZN( u0_u3_u4_n115 ) , .B2( u0_u3_u4_n145 ) , .B1( u0_u3_u4_n146 ) , .A( u0_u3_u4_n156 ) );
  OAI22_X1 u0_u3_u4_U15 (.ZN( u0_u3_u4_n114 ) , .A2( u0_u3_u4_n121 ) , .B1( u0_u3_u4_n160 ) , .B2( u0_u3_u4_n170 ) , .A1( u0_u3_u4_n171 ) );
  NAND2_X1 u0_u3_u4_U16 (.ZN( u0_u3_u4_n132 ) , .A2( u0_u3_u4_n170 ) , .A1( u0_u3_u4_n173 ) );
  AOI21_X1 u0_u3_u4_U17 (.B2( u0_u3_u4_n160 ) , .B1( u0_u3_u4_n161 ) , .ZN( u0_u3_u4_n162 ) , .A( u0_u3_u4_n170 ) );
  AOI21_X1 u0_u3_u4_U18 (.ZN( u0_u3_u4_n107 ) , .B2( u0_u3_u4_n143 ) , .A( u0_u3_u4_n174 ) , .B1( u0_u3_u4_n184 ) );
  AOI21_X1 u0_u3_u4_U19 (.B2( u0_u3_u4_n158 ) , .B1( u0_u3_u4_n159 ) , .ZN( u0_u3_u4_n163 ) , .A( u0_u3_u4_n174 ) );
  AOI21_X1 u0_u3_u4_U20 (.A( u0_u3_u4_n153 ) , .B2( u0_u3_u4_n154 ) , .B1( u0_u3_u4_n155 ) , .ZN( u0_u3_u4_n165 ) );
  AOI21_X1 u0_u3_u4_U21 (.A( u0_u3_u4_n156 ) , .B2( u0_u3_u4_n157 ) , .ZN( u0_u3_u4_n164 ) , .B1( u0_u3_u4_n184 ) );
  INV_X1 u0_u3_u4_U22 (.A( u0_u3_u4_n138 ) , .ZN( u0_u3_u4_n170 ) );
  AND2_X1 u0_u3_u4_U23 (.A2( u0_u3_u4_n120 ) , .ZN( u0_u3_u4_n155 ) , .A1( u0_u3_u4_n160 ) );
  INV_X1 u0_u3_u4_U24 (.A( u0_u3_u4_n156 ) , .ZN( u0_u3_u4_n175 ) );
  NAND2_X1 u0_u3_u4_U25 (.A2( u0_u3_u4_n118 ) , .ZN( u0_u3_u4_n131 ) , .A1( u0_u3_u4_n147 ) );
  NAND2_X1 u0_u3_u4_U26 (.A1( u0_u3_u4_n119 ) , .A2( u0_u3_u4_n120 ) , .ZN( u0_u3_u4_n130 ) );
  NAND2_X1 u0_u3_u4_U27 (.ZN( u0_u3_u4_n117 ) , .A2( u0_u3_u4_n118 ) , .A1( u0_u3_u4_n148 ) );
  NAND2_X1 u0_u3_u4_U28 (.ZN( u0_u3_u4_n129 ) , .A1( u0_u3_u4_n134 ) , .A2( u0_u3_u4_n148 ) );
  AND3_X1 u0_u3_u4_U29 (.A1( u0_u3_u4_n119 ) , .A2( u0_u3_u4_n143 ) , .A3( u0_u3_u4_n154 ) , .ZN( u0_u3_u4_n161 ) );
  NOR2_X1 u0_u3_u4_U3 (.ZN( u0_u3_u4_n121 ) , .A1( u0_u3_u4_n181 ) , .A2( u0_u3_u4_n182 ) );
  AND2_X1 u0_u3_u4_U30 (.A1( u0_u3_u4_n145 ) , .A2( u0_u3_u4_n147 ) , .ZN( u0_u3_u4_n159 ) );
  INV_X1 u0_u3_u4_U31 (.A( u0_u3_u4_n158 ) , .ZN( u0_u3_u4_n182 ) );
  INV_X1 u0_u3_u4_U32 (.ZN( u0_u3_u4_n181 ) , .A( u0_u3_u4_n96 ) );
  INV_X1 u0_u3_u4_U33 (.A( u0_u3_u4_n144 ) , .ZN( u0_u3_u4_n179 ) );
  INV_X1 u0_u3_u4_U34 (.A( u0_u3_u4_n157 ) , .ZN( u0_u3_u4_n178 ) );
  NAND2_X1 u0_u3_u4_U35 (.A2( u0_u3_u4_n154 ) , .A1( u0_u3_u4_n96 ) , .ZN( u0_u3_u4_n97 ) );
  INV_X1 u0_u3_u4_U36 (.ZN( u0_u3_u4_n186 ) , .A( u0_u3_u4_n95 ) );
  OAI221_X1 u0_u3_u4_U37 (.C1( u0_u3_u4_n134 ) , .B1( u0_u3_u4_n158 ) , .B2( u0_u3_u4_n171 ) , .C2( u0_u3_u4_n173 ) , .A( u0_u3_u4_n94 ) , .ZN( u0_u3_u4_n95 ) );
  AOI222_X1 u0_u3_u4_U38 (.B2( u0_u3_u4_n132 ) , .A1( u0_u3_u4_n138 ) , .C2( u0_u3_u4_n175 ) , .A2( u0_u3_u4_n179 ) , .C1( u0_u3_u4_n181 ) , .B1( u0_u3_u4_n185 ) , .ZN( u0_u3_u4_n94 ) );
  INV_X1 u0_u3_u4_U39 (.A( u0_u3_u4_n113 ) , .ZN( u0_u3_u4_n185 ) );
  INV_X1 u0_u3_u4_U4 (.A( u0_u3_u4_n117 ) , .ZN( u0_u3_u4_n184 ) );
  INV_X1 u0_u3_u4_U40 (.A( u0_u3_u4_n143 ) , .ZN( u0_u3_u4_n183 ) );
  NOR2_X1 u0_u3_u4_U41 (.ZN( u0_u3_u4_n138 ) , .A1( u0_u3_u4_n168 ) , .A2( u0_u3_u4_n169 ) );
  NOR2_X1 u0_u3_u4_U42 (.A1( u0_u3_u4_n150 ) , .A2( u0_u3_u4_n152 ) , .ZN( u0_u3_u4_n153 ) );
  NOR2_X1 u0_u3_u4_U43 (.A2( u0_u3_u4_n128 ) , .A1( u0_u3_u4_n138 ) , .ZN( u0_u3_u4_n156 ) );
  AOI22_X1 u0_u3_u4_U44 (.B2( u0_u3_u4_n122 ) , .A1( u0_u3_u4_n123 ) , .ZN( u0_u3_u4_n124 ) , .B1( u0_u3_u4_n128 ) , .A2( u0_u3_u4_n172 ) );
  INV_X1 u0_u3_u4_U45 (.A( u0_u3_u4_n153 ) , .ZN( u0_u3_u4_n172 ) );
  NAND2_X1 u0_u3_u4_U46 (.A2( u0_u3_u4_n120 ) , .ZN( u0_u3_u4_n123 ) , .A1( u0_u3_u4_n161 ) );
  AOI22_X1 u0_u3_u4_U47 (.B2( u0_u3_u4_n132 ) , .A2( u0_u3_u4_n133 ) , .ZN( u0_u3_u4_n140 ) , .A1( u0_u3_u4_n150 ) , .B1( u0_u3_u4_n179 ) );
  NAND2_X1 u0_u3_u4_U48 (.ZN( u0_u3_u4_n133 ) , .A2( u0_u3_u4_n146 ) , .A1( u0_u3_u4_n154 ) );
  NAND2_X1 u0_u3_u4_U49 (.A1( u0_u3_u4_n103 ) , .ZN( u0_u3_u4_n154 ) , .A2( u0_u3_u4_n98 ) );
  NOR4_X1 u0_u3_u4_U5 (.A4( u0_u3_u4_n106 ) , .A3( u0_u3_u4_n107 ) , .A2( u0_u3_u4_n108 ) , .A1( u0_u3_u4_n109 ) , .ZN( u0_u3_u4_n110 ) );
  NAND2_X1 u0_u3_u4_U50 (.A1( u0_u3_u4_n101 ) , .ZN( u0_u3_u4_n158 ) , .A2( u0_u3_u4_n99 ) );
  AOI21_X1 u0_u3_u4_U51 (.ZN( u0_u3_u4_n127 ) , .A( u0_u3_u4_n136 ) , .B2( u0_u3_u4_n150 ) , .B1( u0_u3_u4_n180 ) );
  INV_X1 u0_u3_u4_U52 (.A( u0_u3_u4_n160 ) , .ZN( u0_u3_u4_n180 ) );
  NAND2_X1 u0_u3_u4_U53 (.A2( u0_u3_u4_n104 ) , .A1( u0_u3_u4_n105 ) , .ZN( u0_u3_u4_n146 ) );
  NAND2_X1 u0_u3_u4_U54 (.A2( u0_u3_u4_n101 ) , .A1( u0_u3_u4_n102 ) , .ZN( u0_u3_u4_n160 ) );
  NAND2_X1 u0_u3_u4_U55 (.ZN( u0_u3_u4_n134 ) , .A1( u0_u3_u4_n98 ) , .A2( u0_u3_u4_n99 ) );
  NAND2_X1 u0_u3_u4_U56 (.A1( u0_u3_u4_n103 ) , .A2( u0_u3_u4_n104 ) , .ZN( u0_u3_u4_n143 ) );
  NAND2_X1 u0_u3_u4_U57 (.A2( u0_u3_u4_n105 ) , .ZN( u0_u3_u4_n145 ) , .A1( u0_u3_u4_n98 ) );
  NAND2_X1 u0_u3_u4_U58 (.A1( u0_u3_u4_n100 ) , .A2( u0_u3_u4_n105 ) , .ZN( u0_u3_u4_n120 ) );
  NAND2_X1 u0_u3_u4_U59 (.A1( u0_u3_u4_n102 ) , .A2( u0_u3_u4_n104 ) , .ZN( u0_u3_u4_n148 ) );
  AOI21_X1 u0_u3_u4_U6 (.ZN( u0_u3_u4_n106 ) , .B2( u0_u3_u4_n146 ) , .B1( u0_u3_u4_n158 ) , .A( u0_u3_u4_n170 ) );
  NAND2_X1 u0_u3_u4_U60 (.A2( u0_u3_u4_n100 ) , .A1( u0_u3_u4_n103 ) , .ZN( u0_u3_u4_n157 ) );
  INV_X1 u0_u3_u4_U61 (.A( u0_u3_u4_n150 ) , .ZN( u0_u3_u4_n173 ) );
  INV_X1 u0_u3_u4_U62 (.A( u0_u3_u4_n152 ) , .ZN( u0_u3_u4_n171 ) );
  NAND2_X1 u0_u3_u4_U63 (.A1( u0_u3_u4_n100 ) , .ZN( u0_u3_u4_n118 ) , .A2( u0_u3_u4_n99 ) );
  NAND2_X1 u0_u3_u4_U64 (.A2( u0_u3_u4_n100 ) , .A1( u0_u3_u4_n102 ) , .ZN( u0_u3_u4_n144 ) );
  NAND2_X1 u0_u3_u4_U65 (.A2( u0_u3_u4_n101 ) , .A1( u0_u3_u4_n105 ) , .ZN( u0_u3_u4_n96 ) );
  INV_X1 u0_u3_u4_U66 (.A( u0_u3_u4_n128 ) , .ZN( u0_u3_u4_n174 ) );
  NAND2_X1 u0_u3_u4_U67 (.A2( u0_u3_u4_n102 ) , .ZN( u0_u3_u4_n119 ) , .A1( u0_u3_u4_n98 ) );
  NAND2_X1 u0_u3_u4_U68 (.A2( u0_u3_u4_n101 ) , .A1( u0_u3_u4_n103 ) , .ZN( u0_u3_u4_n147 ) );
  NAND2_X1 u0_u3_u4_U69 (.A2( u0_u3_u4_n104 ) , .ZN( u0_u3_u4_n113 ) , .A1( u0_u3_u4_n99 ) );
  AOI21_X1 u0_u3_u4_U7 (.ZN( u0_u3_u4_n109 ) , .A( u0_u3_u4_n153 ) , .B1( u0_u3_u4_n159 ) , .B2( u0_u3_u4_n184 ) );
  NOR2_X1 u0_u3_u4_U70 (.A2( u0_u3_X_28 ) , .ZN( u0_u3_u4_n150 ) , .A1( u0_u3_u4_n168 ) );
  NOR2_X1 u0_u3_u4_U71 (.A2( u0_u3_X_29 ) , .ZN( u0_u3_u4_n152 ) , .A1( u0_u3_u4_n169 ) );
  NOR2_X1 u0_u3_u4_U72 (.A2( u0_u3_X_30 ) , .ZN( u0_u3_u4_n105 ) , .A1( u0_u3_u4_n176 ) );
  NOR2_X1 u0_u3_u4_U73 (.A2( u0_u3_X_26 ) , .ZN( u0_u3_u4_n100 ) , .A1( u0_u3_u4_n177 ) );
  NOR2_X1 u0_u3_u4_U74 (.A2( u0_u3_X_28 ) , .A1( u0_u3_X_29 ) , .ZN( u0_u3_u4_n128 ) );
  NOR2_X1 u0_u3_u4_U75 (.A2( u0_u3_X_27 ) , .A1( u0_u3_X_30 ) , .ZN( u0_u3_u4_n102 ) );
  NOR2_X1 u0_u3_u4_U76 (.A2( u0_u3_X_25 ) , .A1( u0_u3_X_26 ) , .ZN( u0_u3_u4_n98 ) );
  AND2_X1 u0_u3_u4_U77 (.A2( u0_u3_X_25 ) , .A1( u0_u3_X_26 ) , .ZN( u0_u3_u4_n104 ) );
  AND2_X1 u0_u3_u4_U78 (.A1( u0_u3_X_30 ) , .A2( u0_u3_u4_n176 ) , .ZN( u0_u3_u4_n99 ) );
  AND2_X1 u0_u3_u4_U79 (.A1( u0_u3_X_26 ) , .ZN( u0_u3_u4_n101 ) , .A2( u0_u3_u4_n177 ) );
  AOI21_X1 u0_u3_u4_U8 (.ZN( u0_u3_u4_n108 ) , .B2( u0_u3_u4_n134 ) , .B1( u0_u3_u4_n155 ) , .A( u0_u3_u4_n156 ) );
  AND2_X1 u0_u3_u4_U80 (.A1( u0_u3_X_27 ) , .A2( u0_u3_X_30 ) , .ZN( u0_u3_u4_n103 ) );
  INV_X1 u0_u3_u4_U81 (.A( u0_u3_X_28 ) , .ZN( u0_u3_u4_n169 ) );
  INV_X1 u0_u3_u4_U82 (.A( u0_u3_X_29 ) , .ZN( u0_u3_u4_n168 ) );
  INV_X1 u0_u3_u4_U83 (.A( u0_u3_X_25 ) , .ZN( u0_u3_u4_n177 ) );
  INV_X1 u0_u3_u4_U84 (.A( u0_u3_X_27 ) , .ZN( u0_u3_u4_n176 ) );
  NAND4_X1 u0_u3_u4_U85 (.ZN( u0_out3_25 ) , .A4( u0_u3_u4_n139 ) , .A3( u0_u3_u4_n140 ) , .A2( u0_u3_u4_n141 ) , .A1( u0_u3_u4_n142 ) );
  OAI21_X1 u0_u3_u4_U86 (.A( u0_u3_u4_n128 ) , .B2( u0_u3_u4_n129 ) , .B1( u0_u3_u4_n130 ) , .ZN( u0_u3_u4_n142 ) );
  OAI21_X1 u0_u3_u4_U87 (.B2( u0_u3_u4_n131 ) , .ZN( u0_u3_u4_n141 ) , .A( u0_u3_u4_n175 ) , .B1( u0_u3_u4_n183 ) );
  NAND4_X1 u0_u3_u4_U88 (.ZN( u0_out3_14 ) , .A4( u0_u3_u4_n124 ) , .A3( u0_u3_u4_n125 ) , .A2( u0_u3_u4_n126 ) , .A1( u0_u3_u4_n127 ) );
  AOI22_X1 u0_u3_u4_U89 (.B2( u0_u3_u4_n117 ) , .ZN( u0_u3_u4_n126 ) , .A1( u0_u3_u4_n129 ) , .B1( u0_u3_u4_n152 ) , .A2( u0_u3_u4_n175 ) );
  AOI211_X1 u0_u3_u4_U9 (.B( u0_u3_u4_n136 ) , .A( u0_u3_u4_n137 ) , .C2( u0_u3_u4_n138 ) , .ZN( u0_u3_u4_n139 ) , .C1( u0_u3_u4_n182 ) );
  AOI22_X1 u0_u3_u4_U90 (.ZN( u0_u3_u4_n125 ) , .B2( u0_u3_u4_n131 ) , .A2( u0_u3_u4_n132 ) , .B1( u0_u3_u4_n138 ) , .A1( u0_u3_u4_n178 ) );
  AOI22_X1 u0_u3_u4_U91 (.B2( u0_u3_u4_n149 ) , .B1( u0_u3_u4_n150 ) , .A2( u0_u3_u4_n151 ) , .A1( u0_u3_u4_n152 ) , .ZN( u0_u3_u4_n167 ) );
  NOR4_X1 u0_u3_u4_U92 (.A4( u0_u3_u4_n162 ) , .A3( u0_u3_u4_n163 ) , .A2( u0_u3_u4_n164 ) , .A1( u0_u3_u4_n165 ) , .ZN( u0_u3_u4_n166 ) );
  NAND4_X1 u0_u3_u4_U93 (.ZN( u0_out3_8 ) , .A4( u0_u3_u4_n110 ) , .A3( u0_u3_u4_n111 ) , .A2( u0_u3_u4_n112 ) , .A1( u0_u3_u4_n186 ) );
  NAND2_X1 u0_u3_u4_U94 (.ZN( u0_u3_u4_n112 ) , .A2( u0_u3_u4_n130 ) , .A1( u0_u3_u4_n150 ) );
  AOI22_X1 u0_u3_u4_U95 (.ZN( u0_u3_u4_n111 ) , .B2( u0_u3_u4_n132 ) , .A1( u0_u3_u4_n152 ) , .B1( u0_u3_u4_n178 ) , .A2( u0_u3_u4_n97 ) );
  NAND3_X1 u0_u3_u4_U96 (.ZN( u0_out3_3 ) , .A3( u0_u3_u4_n166 ) , .A1( u0_u3_u4_n167 ) , .A2( u0_u3_u4_n186 ) );
  NAND3_X1 u0_u3_u4_U97 (.A3( u0_u3_u4_n146 ) , .A2( u0_u3_u4_n147 ) , .A1( u0_u3_u4_n148 ) , .ZN( u0_u3_u4_n149 ) );
  NAND3_X1 u0_u3_u4_U98 (.A3( u0_u3_u4_n143 ) , .A2( u0_u3_u4_n144 ) , .A1( u0_u3_u4_n145 ) , .ZN( u0_u3_u4_n151 ) );
  NAND3_X1 u0_u3_u4_U99 (.A3( u0_u3_u4_n121 ) , .ZN( u0_u3_u4_n122 ) , .A2( u0_u3_u4_n144 ) , .A1( u0_u3_u4_n154 ) );
  INV_X1 u0_u3_u5_U10 (.A( u0_u3_u5_n121 ) , .ZN( u0_u3_u5_n177 ) );
  NOR3_X1 u0_u3_u5_U100 (.A3( u0_u3_u5_n141 ) , .A1( u0_u3_u5_n142 ) , .ZN( u0_u3_u5_n143 ) , .A2( u0_u3_u5_n191 ) );
  NAND4_X1 u0_u3_u5_U101 (.ZN( u0_out3_4 ) , .A4( u0_u3_u5_n112 ) , .A2( u0_u3_u5_n113 ) , .A1( u0_u3_u5_n114 ) , .A3( u0_u3_u5_n195 ) );
  AOI211_X1 u0_u3_u5_U102 (.A( u0_u3_u5_n110 ) , .C1( u0_u3_u5_n111 ) , .ZN( u0_u3_u5_n112 ) , .B( u0_u3_u5_n118 ) , .C2( u0_u3_u5_n177 ) );
  AOI222_X1 u0_u3_u5_U103 (.ZN( u0_u3_u5_n113 ) , .A1( u0_u3_u5_n131 ) , .C1( u0_u3_u5_n148 ) , .B2( u0_u3_u5_n174 ) , .C2( u0_u3_u5_n178 ) , .A2( u0_u3_u5_n179 ) , .B1( u0_u3_u5_n99 ) );
  NAND3_X1 u0_u3_u5_U104 (.A2( u0_u3_u5_n154 ) , .A3( u0_u3_u5_n158 ) , .A1( u0_u3_u5_n161 ) , .ZN( u0_u3_u5_n99 ) );
  NOR2_X1 u0_u3_u5_U11 (.ZN( u0_u3_u5_n160 ) , .A2( u0_u3_u5_n173 ) , .A1( u0_u3_u5_n177 ) );
  INV_X1 u0_u3_u5_U12 (.A( u0_u3_u5_n150 ) , .ZN( u0_u3_u5_n174 ) );
  AOI21_X1 u0_u3_u5_U13 (.A( u0_u3_u5_n160 ) , .B2( u0_u3_u5_n161 ) , .ZN( u0_u3_u5_n162 ) , .B1( u0_u3_u5_n192 ) );
  INV_X1 u0_u3_u5_U14 (.A( u0_u3_u5_n159 ) , .ZN( u0_u3_u5_n192 ) );
  AOI21_X1 u0_u3_u5_U15 (.A( u0_u3_u5_n156 ) , .B2( u0_u3_u5_n157 ) , .B1( u0_u3_u5_n158 ) , .ZN( u0_u3_u5_n163 ) );
  AOI21_X1 u0_u3_u5_U16 (.B2( u0_u3_u5_n139 ) , .B1( u0_u3_u5_n140 ) , .ZN( u0_u3_u5_n141 ) , .A( u0_u3_u5_n150 ) );
  OAI21_X1 u0_u3_u5_U17 (.A( u0_u3_u5_n133 ) , .B2( u0_u3_u5_n134 ) , .B1( u0_u3_u5_n135 ) , .ZN( u0_u3_u5_n142 ) );
  OAI21_X1 u0_u3_u5_U18 (.ZN( u0_u3_u5_n133 ) , .B2( u0_u3_u5_n147 ) , .A( u0_u3_u5_n173 ) , .B1( u0_u3_u5_n188 ) );
  NAND2_X1 u0_u3_u5_U19 (.A2( u0_u3_u5_n119 ) , .A1( u0_u3_u5_n123 ) , .ZN( u0_u3_u5_n137 ) );
  INV_X1 u0_u3_u5_U20 (.A( u0_u3_u5_n155 ) , .ZN( u0_u3_u5_n194 ) );
  NAND2_X1 u0_u3_u5_U21 (.A1( u0_u3_u5_n121 ) , .ZN( u0_u3_u5_n132 ) , .A2( u0_u3_u5_n172 ) );
  NAND2_X1 u0_u3_u5_U22 (.A2( u0_u3_u5_n122 ) , .ZN( u0_u3_u5_n136 ) , .A1( u0_u3_u5_n154 ) );
  NAND2_X1 u0_u3_u5_U23 (.A2( u0_u3_u5_n119 ) , .A1( u0_u3_u5_n120 ) , .ZN( u0_u3_u5_n159 ) );
  INV_X1 u0_u3_u5_U24 (.A( u0_u3_u5_n156 ) , .ZN( u0_u3_u5_n175 ) );
  INV_X1 u0_u3_u5_U25 (.A( u0_u3_u5_n158 ) , .ZN( u0_u3_u5_n188 ) );
  INV_X1 u0_u3_u5_U26 (.A( u0_u3_u5_n152 ) , .ZN( u0_u3_u5_n179 ) );
  INV_X1 u0_u3_u5_U27 (.A( u0_u3_u5_n140 ) , .ZN( u0_u3_u5_n182 ) );
  INV_X1 u0_u3_u5_U28 (.A( u0_u3_u5_n151 ) , .ZN( u0_u3_u5_n183 ) );
  INV_X1 u0_u3_u5_U29 (.A( u0_u3_u5_n123 ) , .ZN( u0_u3_u5_n185 ) );
  NOR2_X1 u0_u3_u5_U3 (.ZN( u0_u3_u5_n134 ) , .A1( u0_u3_u5_n183 ) , .A2( u0_u3_u5_n190 ) );
  INV_X1 u0_u3_u5_U30 (.A( u0_u3_u5_n161 ) , .ZN( u0_u3_u5_n184 ) );
  INV_X1 u0_u3_u5_U31 (.A( u0_u3_u5_n139 ) , .ZN( u0_u3_u5_n189 ) );
  INV_X1 u0_u3_u5_U32 (.A( u0_u3_u5_n157 ) , .ZN( u0_u3_u5_n190 ) );
  INV_X1 u0_u3_u5_U33 (.A( u0_u3_u5_n120 ) , .ZN( u0_u3_u5_n193 ) );
  NAND2_X1 u0_u3_u5_U34 (.ZN( u0_u3_u5_n111 ) , .A1( u0_u3_u5_n140 ) , .A2( u0_u3_u5_n155 ) );
  INV_X1 u0_u3_u5_U35 (.A( u0_u3_u5_n117 ) , .ZN( u0_u3_u5_n196 ) );
  OAI221_X1 u0_u3_u5_U36 (.A( u0_u3_u5_n116 ) , .ZN( u0_u3_u5_n117 ) , .B2( u0_u3_u5_n119 ) , .C1( u0_u3_u5_n153 ) , .C2( u0_u3_u5_n158 ) , .B1( u0_u3_u5_n172 ) );
  AOI222_X1 u0_u3_u5_U37 (.ZN( u0_u3_u5_n116 ) , .B2( u0_u3_u5_n145 ) , .C1( u0_u3_u5_n148 ) , .A2( u0_u3_u5_n174 ) , .C2( u0_u3_u5_n177 ) , .B1( u0_u3_u5_n187 ) , .A1( u0_u3_u5_n193 ) );
  INV_X1 u0_u3_u5_U38 (.A( u0_u3_u5_n115 ) , .ZN( u0_u3_u5_n187 ) );
  NOR2_X1 u0_u3_u5_U39 (.ZN( u0_u3_u5_n100 ) , .A1( u0_u3_u5_n170 ) , .A2( u0_u3_u5_n180 ) );
  INV_X1 u0_u3_u5_U4 (.A( u0_u3_u5_n138 ) , .ZN( u0_u3_u5_n191 ) );
  AOI22_X1 u0_u3_u5_U40 (.B2( u0_u3_u5_n131 ) , .A2( u0_u3_u5_n146 ) , .ZN( u0_u3_u5_n169 ) , .B1( u0_u3_u5_n174 ) , .A1( u0_u3_u5_n185 ) );
  NOR2_X1 u0_u3_u5_U41 (.A1( u0_u3_u5_n146 ) , .ZN( u0_u3_u5_n150 ) , .A2( u0_u3_u5_n173 ) );
  AOI21_X1 u0_u3_u5_U42 (.A( u0_u3_u5_n118 ) , .B2( u0_u3_u5_n145 ) , .ZN( u0_u3_u5_n168 ) , .B1( u0_u3_u5_n186 ) );
  INV_X1 u0_u3_u5_U43 (.A( u0_u3_u5_n122 ) , .ZN( u0_u3_u5_n186 ) );
  NOR2_X1 u0_u3_u5_U44 (.A1( u0_u3_u5_n146 ) , .ZN( u0_u3_u5_n152 ) , .A2( u0_u3_u5_n176 ) );
  NOR2_X1 u0_u3_u5_U45 (.A1( u0_u3_u5_n115 ) , .ZN( u0_u3_u5_n118 ) , .A2( u0_u3_u5_n153 ) );
  NOR2_X1 u0_u3_u5_U46 (.A2( u0_u3_u5_n145 ) , .ZN( u0_u3_u5_n156 ) , .A1( u0_u3_u5_n174 ) );
  NOR2_X1 u0_u3_u5_U47 (.ZN( u0_u3_u5_n121 ) , .A2( u0_u3_u5_n145 ) , .A1( u0_u3_u5_n176 ) );
  AOI22_X1 u0_u3_u5_U48 (.ZN( u0_u3_u5_n114 ) , .A2( u0_u3_u5_n137 ) , .A1( u0_u3_u5_n145 ) , .B2( u0_u3_u5_n175 ) , .B1( u0_u3_u5_n193 ) );
  OAI211_X1 u0_u3_u5_U49 (.B( u0_u3_u5_n124 ) , .A( u0_u3_u5_n125 ) , .C2( u0_u3_u5_n126 ) , .C1( u0_u3_u5_n127 ) , .ZN( u0_u3_u5_n128 ) );
  OAI21_X1 u0_u3_u5_U5 (.B2( u0_u3_u5_n136 ) , .B1( u0_u3_u5_n137 ) , .ZN( u0_u3_u5_n138 ) , .A( u0_u3_u5_n177 ) );
  NOR3_X1 u0_u3_u5_U50 (.ZN( u0_u3_u5_n127 ) , .A1( u0_u3_u5_n136 ) , .A3( u0_u3_u5_n148 ) , .A2( u0_u3_u5_n182 ) );
  OAI21_X1 u0_u3_u5_U51 (.ZN( u0_u3_u5_n124 ) , .A( u0_u3_u5_n177 ) , .B2( u0_u3_u5_n183 ) , .B1( u0_u3_u5_n189 ) );
  OAI21_X1 u0_u3_u5_U52 (.ZN( u0_u3_u5_n125 ) , .A( u0_u3_u5_n174 ) , .B2( u0_u3_u5_n185 ) , .B1( u0_u3_u5_n190 ) );
  AOI21_X1 u0_u3_u5_U53 (.A( u0_u3_u5_n153 ) , .B2( u0_u3_u5_n154 ) , .B1( u0_u3_u5_n155 ) , .ZN( u0_u3_u5_n164 ) );
  AOI21_X1 u0_u3_u5_U54 (.ZN( u0_u3_u5_n110 ) , .B1( u0_u3_u5_n122 ) , .B2( u0_u3_u5_n139 ) , .A( u0_u3_u5_n153 ) );
  INV_X1 u0_u3_u5_U55 (.A( u0_u3_u5_n153 ) , .ZN( u0_u3_u5_n176 ) );
  INV_X1 u0_u3_u5_U56 (.A( u0_u3_u5_n126 ) , .ZN( u0_u3_u5_n173 ) );
  AND2_X1 u0_u3_u5_U57 (.A2( u0_u3_u5_n104 ) , .A1( u0_u3_u5_n107 ) , .ZN( u0_u3_u5_n147 ) );
  AND2_X1 u0_u3_u5_U58 (.A2( u0_u3_u5_n104 ) , .A1( u0_u3_u5_n108 ) , .ZN( u0_u3_u5_n148 ) );
  NAND2_X1 u0_u3_u5_U59 (.A1( u0_u3_u5_n105 ) , .A2( u0_u3_u5_n106 ) , .ZN( u0_u3_u5_n158 ) );
  INV_X1 u0_u3_u5_U6 (.A( u0_u3_u5_n135 ) , .ZN( u0_u3_u5_n178 ) );
  NAND2_X1 u0_u3_u5_U60 (.A2( u0_u3_u5_n108 ) , .A1( u0_u3_u5_n109 ) , .ZN( u0_u3_u5_n139 ) );
  NAND2_X1 u0_u3_u5_U61 (.A1( u0_u3_u5_n106 ) , .A2( u0_u3_u5_n108 ) , .ZN( u0_u3_u5_n119 ) );
  NAND2_X1 u0_u3_u5_U62 (.A2( u0_u3_u5_n103 ) , .A1( u0_u3_u5_n105 ) , .ZN( u0_u3_u5_n140 ) );
  NAND2_X1 u0_u3_u5_U63 (.A2( u0_u3_u5_n104 ) , .A1( u0_u3_u5_n105 ) , .ZN( u0_u3_u5_n155 ) );
  NAND2_X1 u0_u3_u5_U64 (.A2( u0_u3_u5_n106 ) , .A1( u0_u3_u5_n107 ) , .ZN( u0_u3_u5_n122 ) );
  NAND2_X1 u0_u3_u5_U65 (.A2( u0_u3_u5_n100 ) , .A1( u0_u3_u5_n106 ) , .ZN( u0_u3_u5_n115 ) );
  NAND2_X1 u0_u3_u5_U66 (.A2( u0_u3_u5_n100 ) , .A1( u0_u3_u5_n103 ) , .ZN( u0_u3_u5_n161 ) );
  NAND2_X1 u0_u3_u5_U67 (.A1( u0_u3_u5_n105 ) , .A2( u0_u3_u5_n109 ) , .ZN( u0_u3_u5_n154 ) );
  INV_X1 u0_u3_u5_U68 (.A( u0_u3_u5_n146 ) , .ZN( u0_u3_u5_n172 ) );
  NAND2_X1 u0_u3_u5_U69 (.A1( u0_u3_u5_n103 ) , .A2( u0_u3_u5_n108 ) , .ZN( u0_u3_u5_n123 ) );
  OAI22_X1 u0_u3_u5_U7 (.B2( u0_u3_u5_n149 ) , .B1( u0_u3_u5_n150 ) , .A2( u0_u3_u5_n151 ) , .A1( u0_u3_u5_n152 ) , .ZN( u0_u3_u5_n165 ) );
  NAND2_X1 u0_u3_u5_U70 (.A2( u0_u3_u5_n103 ) , .A1( u0_u3_u5_n107 ) , .ZN( u0_u3_u5_n151 ) );
  NAND2_X1 u0_u3_u5_U71 (.A2( u0_u3_u5_n107 ) , .A1( u0_u3_u5_n109 ) , .ZN( u0_u3_u5_n120 ) );
  NAND2_X1 u0_u3_u5_U72 (.A2( u0_u3_u5_n100 ) , .A1( u0_u3_u5_n109 ) , .ZN( u0_u3_u5_n157 ) );
  AND2_X1 u0_u3_u5_U73 (.A2( u0_u3_u5_n100 ) , .A1( u0_u3_u5_n104 ) , .ZN( u0_u3_u5_n131 ) );
  INV_X1 u0_u3_u5_U74 (.A( u0_u3_u5_n102 ) , .ZN( u0_u3_u5_n195 ) );
  OAI221_X1 u0_u3_u5_U75 (.A( u0_u3_u5_n101 ) , .ZN( u0_u3_u5_n102 ) , .C2( u0_u3_u5_n115 ) , .C1( u0_u3_u5_n126 ) , .B1( u0_u3_u5_n134 ) , .B2( u0_u3_u5_n160 ) );
  OAI21_X1 u0_u3_u5_U76 (.ZN( u0_u3_u5_n101 ) , .B1( u0_u3_u5_n137 ) , .A( u0_u3_u5_n146 ) , .B2( u0_u3_u5_n147 ) );
  NOR2_X1 u0_u3_u5_U77 (.A2( u0_u3_X_34 ) , .A1( u0_u3_X_35 ) , .ZN( u0_u3_u5_n145 ) );
  NOR2_X1 u0_u3_u5_U78 (.A2( u0_u3_X_34 ) , .ZN( u0_u3_u5_n146 ) , .A1( u0_u3_u5_n171 ) );
  NOR2_X1 u0_u3_u5_U79 (.A2( u0_u3_X_31 ) , .A1( u0_u3_X_32 ) , .ZN( u0_u3_u5_n103 ) );
  NOR3_X1 u0_u3_u5_U8 (.A2( u0_u3_u5_n147 ) , .A1( u0_u3_u5_n148 ) , .ZN( u0_u3_u5_n149 ) , .A3( u0_u3_u5_n194 ) );
  NOR2_X1 u0_u3_u5_U80 (.A2( u0_u3_X_36 ) , .ZN( u0_u3_u5_n105 ) , .A1( u0_u3_u5_n180 ) );
  NOR2_X1 u0_u3_u5_U81 (.A2( u0_u3_X_33 ) , .ZN( u0_u3_u5_n108 ) , .A1( u0_u3_u5_n170 ) );
  NOR2_X1 u0_u3_u5_U82 (.A2( u0_u3_X_33 ) , .A1( u0_u3_X_36 ) , .ZN( u0_u3_u5_n107 ) );
  NOR2_X1 u0_u3_u5_U83 (.A2( u0_u3_X_31 ) , .ZN( u0_u3_u5_n104 ) , .A1( u0_u3_u5_n181 ) );
  NAND2_X1 u0_u3_u5_U84 (.A2( u0_u3_X_34 ) , .A1( u0_u3_X_35 ) , .ZN( u0_u3_u5_n153 ) );
  NAND2_X1 u0_u3_u5_U85 (.A1( u0_u3_X_34 ) , .ZN( u0_u3_u5_n126 ) , .A2( u0_u3_u5_n171 ) );
  AND2_X1 u0_u3_u5_U86 (.A1( u0_u3_X_31 ) , .A2( u0_u3_X_32 ) , .ZN( u0_u3_u5_n106 ) );
  AND2_X1 u0_u3_u5_U87 (.A1( u0_u3_X_31 ) , .ZN( u0_u3_u5_n109 ) , .A2( u0_u3_u5_n181 ) );
  INV_X1 u0_u3_u5_U88 (.A( u0_u3_X_33 ) , .ZN( u0_u3_u5_n180 ) );
  INV_X1 u0_u3_u5_U89 (.A( u0_u3_X_35 ) , .ZN( u0_u3_u5_n171 ) );
  NOR2_X1 u0_u3_u5_U9 (.ZN( u0_u3_u5_n135 ) , .A1( u0_u3_u5_n173 ) , .A2( u0_u3_u5_n176 ) );
  INV_X1 u0_u3_u5_U90 (.A( u0_u3_X_36 ) , .ZN( u0_u3_u5_n170 ) );
  INV_X1 u0_u3_u5_U91 (.A( u0_u3_X_32 ) , .ZN( u0_u3_u5_n181 ) );
  NAND4_X1 u0_u3_u5_U92 (.ZN( u0_out3_29 ) , .A4( u0_u3_u5_n129 ) , .A3( u0_u3_u5_n130 ) , .A2( u0_u3_u5_n168 ) , .A1( u0_u3_u5_n196 ) );
  AOI221_X1 u0_u3_u5_U93 (.A( u0_u3_u5_n128 ) , .ZN( u0_u3_u5_n129 ) , .C2( u0_u3_u5_n132 ) , .B2( u0_u3_u5_n159 ) , .B1( u0_u3_u5_n176 ) , .C1( u0_u3_u5_n184 ) );
  AOI222_X1 u0_u3_u5_U94 (.ZN( u0_u3_u5_n130 ) , .A2( u0_u3_u5_n146 ) , .B1( u0_u3_u5_n147 ) , .C2( u0_u3_u5_n175 ) , .B2( u0_u3_u5_n179 ) , .A1( u0_u3_u5_n188 ) , .C1( u0_u3_u5_n194 ) );
  NAND4_X1 u0_u3_u5_U95 (.ZN( u0_out3_19 ) , .A4( u0_u3_u5_n166 ) , .A3( u0_u3_u5_n167 ) , .A2( u0_u3_u5_n168 ) , .A1( u0_u3_u5_n169 ) );
  AOI22_X1 u0_u3_u5_U96 (.B2( u0_u3_u5_n145 ) , .A2( u0_u3_u5_n146 ) , .ZN( u0_u3_u5_n167 ) , .B1( u0_u3_u5_n182 ) , .A1( u0_u3_u5_n189 ) );
  NOR4_X1 u0_u3_u5_U97 (.A4( u0_u3_u5_n162 ) , .A3( u0_u3_u5_n163 ) , .A2( u0_u3_u5_n164 ) , .A1( u0_u3_u5_n165 ) , .ZN( u0_u3_u5_n166 ) );
  NAND4_X1 u0_u3_u5_U98 (.ZN( u0_out3_11 ) , .A4( u0_u3_u5_n143 ) , .A3( u0_u3_u5_n144 ) , .A2( u0_u3_u5_n169 ) , .A1( u0_u3_u5_n196 ) );
  AOI22_X1 u0_u3_u5_U99 (.A2( u0_u3_u5_n132 ) , .ZN( u0_u3_u5_n144 ) , .B2( u0_u3_u5_n145 ) , .B1( u0_u3_u5_n184 ) , .A1( u0_u3_u5_n194 ) );
  INV_X1 u0_u3_u6_U10 (.ZN( u0_u3_u6_n172 ) , .A( u0_u3_u6_n88 ) );
  OAI21_X1 u0_u3_u6_U11 (.A( u0_u3_u6_n159 ) , .B1( u0_u3_u6_n169 ) , .B2( u0_u3_u6_n173 ) , .ZN( u0_u3_u6_n90 ) );
  AOI22_X1 u0_u3_u6_U12 (.A2( u0_u3_u6_n151 ) , .B2( u0_u3_u6_n161 ) , .A1( u0_u3_u6_n167 ) , .B1( u0_u3_u6_n170 ) , .ZN( u0_u3_u6_n89 ) );
  AOI21_X1 u0_u3_u6_U13 (.ZN( u0_u3_u6_n106 ) , .A( u0_u3_u6_n142 ) , .B2( u0_u3_u6_n159 ) , .B1( u0_u3_u6_n164 ) );
  INV_X1 u0_u3_u6_U14 (.A( u0_u3_u6_n155 ) , .ZN( u0_u3_u6_n161 ) );
  INV_X1 u0_u3_u6_U15 (.A( u0_u3_u6_n128 ) , .ZN( u0_u3_u6_n164 ) );
  NAND2_X1 u0_u3_u6_U16 (.ZN( u0_u3_u6_n110 ) , .A1( u0_u3_u6_n122 ) , .A2( u0_u3_u6_n129 ) );
  NAND2_X1 u0_u3_u6_U17 (.ZN( u0_u3_u6_n124 ) , .A2( u0_u3_u6_n146 ) , .A1( u0_u3_u6_n148 ) );
  INV_X1 u0_u3_u6_U18 (.A( u0_u3_u6_n132 ) , .ZN( u0_u3_u6_n171 ) );
  AND2_X1 u0_u3_u6_U19 (.A1( u0_u3_u6_n100 ) , .ZN( u0_u3_u6_n130 ) , .A2( u0_u3_u6_n147 ) );
  INV_X1 u0_u3_u6_U20 (.A( u0_u3_u6_n127 ) , .ZN( u0_u3_u6_n173 ) );
  INV_X1 u0_u3_u6_U21 (.A( u0_u3_u6_n121 ) , .ZN( u0_u3_u6_n167 ) );
  INV_X1 u0_u3_u6_U22 (.A( u0_u3_u6_n100 ) , .ZN( u0_u3_u6_n169 ) );
  INV_X1 u0_u3_u6_U23 (.A( u0_u3_u6_n123 ) , .ZN( u0_u3_u6_n170 ) );
  INV_X1 u0_u3_u6_U24 (.A( u0_u3_u6_n113 ) , .ZN( u0_u3_u6_n168 ) );
  AND2_X1 u0_u3_u6_U25 (.A1( u0_u3_u6_n107 ) , .A2( u0_u3_u6_n119 ) , .ZN( u0_u3_u6_n133 ) );
  AND2_X1 u0_u3_u6_U26 (.A2( u0_u3_u6_n121 ) , .A1( u0_u3_u6_n122 ) , .ZN( u0_u3_u6_n131 ) );
  AND3_X1 u0_u3_u6_U27 (.ZN( u0_u3_u6_n120 ) , .A2( u0_u3_u6_n127 ) , .A1( u0_u3_u6_n132 ) , .A3( u0_u3_u6_n145 ) );
  INV_X1 u0_u3_u6_U28 (.A( u0_u3_u6_n146 ) , .ZN( u0_u3_u6_n163 ) );
  AOI222_X1 u0_u3_u6_U29 (.ZN( u0_u3_u6_n114 ) , .A1( u0_u3_u6_n118 ) , .A2( u0_u3_u6_n126 ) , .B2( u0_u3_u6_n151 ) , .C2( u0_u3_u6_n159 ) , .C1( u0_u3_u6_n168 ) , .B1( u0_u3_u6_n169 ) );
  INV_X1 u0_u3_u6_U3 (.A( u0_u3_u6_n110 ) , .ZN( u0_u3_u6_n166 ) );
  NOR2_X1 u0_u3_u6_U30 (.A1( u0_u3_u6_n162 ) , .A2( u0_u3_u6_n165 ) , .ZN( u0_u3_u6_n98 ) );
  NAND2_X1 u0_u3_u6_U31 (.A1( u0_u3_u6_n144 ) , .ZN( u0_u3_u6_n151 ) , .A2( u0_u3_u6_n158 ) );
  NAND2_X1 u0_u3_u6_U32 (.ZN( u0_u3_u6_n132 ) , .A1( u0_u3_u6_n91 ) , .A2( u0_u3_u6_n97 ) );
  AOI22_X1 u0_u3_u6_U33 (.B2( u0_u3_u6_n110 ) , .B1( u0_u3_u6_n111 ) , .A1( u0_u3_u6_n112 ) , .ZN( u0_u3_u6_n115 ) , .A2( u0_u3_u6_n161 ) );
  NAND4_X1 u0_u3_u6_U34 (.A3( u0_u3_u6_n109 ) , .ZN( u0_u3_u6_n112 ) , .A4( u0_u3_u6_n132 ) , .A2( u0_u3_u6_n147 ) , .A1( u0_u3_u6_n166 ) );
  NOR2_X1 u0_u3_u6_U35 (.ZN( u0_u3_u6_n109 ) , .A1( u0_u3_u6_n170 ) , .A2( u0_u3_u6_n173 ) );
  NOR2_X1 u0_u3_u6_U36 (.A2( u0_u3_u6_n126 ) , .ZN( u0_u3_u6_n155 ) , .A1( u0_u3_u6_n160 ) );
  NAND2_X1 u0_u3_u6_U37 (.ZN( u0_u3_u6_n146 ) , .A2( u0_u3_u6_n94 ) , .A1( u0_u3_u6_n99 ) );
  AOI21_X1 u0_u3_u6_U38 (.A( u0_u3_u6_n144 ) , .B2( u0_u3_u6_n145 ) , .B1( u0_u3_u6_n146 ) , .ZN( u0_u3_u6_n150 ) );
  AOI211_X1 u0_u3_u6_U39 (.B( u0_u3_u6_n134 ) , .A( u0_u3_u6_n135 ) , .C1( u0_u3_u6_n136 ) , .ZN( u0_u3_u6_n137 ) , .C2( u0_u3_u6_n151 ) );
  INV_X1 u0_u3_u6_U4 (.A( u0_u3_u6_n142 ) , .ZN( u0_u3_u6_n174 ) );
  AOI21_X1 u0_u3_u6_U40 (.B2( u0_u3_u6_n132 ) , .B1( u0_u3_u6_n133 ) , .ZN( u0_u3_u6_n134 ) , .A( u0_u3_u6_n158 ) );
  NAND4_X1 u0_u3_u6_U41 (.A4( u0_u3_u6_n127 ) , .A3( u0_u3_u6_n128 ) , .A2( u0_u3_u6_n129 ) , .A1( u0_u3_u6_n130 ) , .ZN( u0_u3_u6_n136 ) );
  AOI21_X1 u0_u3_u6_U42 (.B1( u0_u3_u6_n131 ) , .ZN( u0_u3_u6_n135 ) , .A( u0_u3_u6_n144 ) , .B2( u0_u3_u6_n146 ) );
  INV_X1 u0_u3_u6_U43 (.A( u0_u3_u6_n111 ) , .ZN( u0_u3_u6_n158 ) );
  NAND2_X1 u0_u3_u6_U44 (.ZN( u0_u3_u6_n127 ) , .A1( u0_u3_u6_n91 ) , .A2( u0_u3_u6_n92 ) );
  NAND2_X1 u0_u3_u6_U45 (.ZN( u0_u3_u6_n129 ) , .A2( u0_u3_u6_n95 ) , .A1( u0_u3_u6_n96 ) );
  INV_X1 u0_u3_u6_U46 (.A( u0_u3_u6_n144 ) , .ZN( u0_u3_u6_n159 ) );
  NAND2_X1 u0_u3_u6_U47 (.ZN( u0_u3_u6_n145 ) , .A2( u0_u3_u6_n97 ) , .A1( u0_u3_u6_n98 ) );
  NAND2_X1 u0_u3_u6_U48 (.ZN( u0_u3_u6_n148 ) , .A2( u0_u3_u6_n92 ) , .A1( u0_u3_u6_n94 ) );
  NAND2_X1 u0_u3_u6_U49 (.ZN( u0_u3_u6_n108 ) , .A2( u0_u3_u6_n139 ) , .A1( u0_u3_u6_n144 ) );
  NAND2_X1 u0_u3_u6_U5 (.A2( u0_u3_u6_n143 ) , .ZN( u0_u3_u6_n152 ) , .A1( u0_u3_u6_n166 ) );
  NAND2_X1 u0_u3_u6_U50 (.ZN( u0_u3_u6_n121 ) , .A2( u0_u3_u6_n95 ) , .A1( u0_u3_u6_n97 ) );
  NAND2_X1 u0_u3_u6_U51 (.ZN( u0_u3_u6_n107 ) , .A2( u0_u3_u6_n92 ) , .A1( u0_u3_u6_n95 ) );
  AND2_X1 u0_u3_u6_U52 (.ZN( u0_u3_u6_n118 ) , .A2( u0_u3_u6_n91 ) , .A1( u0_u3_u6_n99 ) );
  NAND2_X1 u0_u3_u6_U53 (.ZN( u0_u3_u6_n147 ) , .A2( u0_u3_u6_n98 ) , .A1( u0_u3_u6_n99 ) );
  NAND2_X1 u0_u3_u6_U54 (.ZN( u0_u3_u6_n128 ) , .A1( u0_u3_u6_n94 ) , .A2( u0_u3_u6_n96 ) );
  NAND2_X1 u0_u3_u6_U55 (.ZN( u0_u3_u6_n119 ) , .A2( u0_u3_u6_n95 ) , .A1( u0_u3_u6_n99 ) );
  NAND2_X1 u0_u3_u6_U56 (.ZN( u0_u3_u6_n123 ) , .A2( u0_u3_u6_n91 ) , .A1( u0_u3_u6_n96 ) );
  NAND2_X1 u0_u3_u6_U57 (.ZN( u0_u3_u6_n100 ) , .A2( u0_u3_u6_n92 ) , .A1( u0_u3_u6_n98 ) );
  NAND2_X1 u0_u3_u6_U58 (.ZN( u0_u3_u6_n122 ) , .A1( u0_u3_u6_n94 ) , .A2( u0_u3_u6_n97 ) );
  INV_X1 u0_u3_u6_U59 (.A( u0_u3_u6_n139 ) , .ZN( u0_u3_u6_n160 ) );
  AOI22_X1 u0_u3_u6_U6 (.B2( u0_u3_u6_n101 ) , .A1( u0_u3_u6_n102 ) , .ZN( u0_u3_u6_n103 ) , .B1( u0_u3_u6_n160 ) , .A2( u0_u3_u6_n161 ) );
  NAND2_X1 u0_u3_u6_U60 (.ZN( u0_u3_u6_n113 ) , .A1( u0_u3_u6_n96 ) , .A2( u0_u3_u6_n98 ) );
  NOR2_X1 u0_u3_u6_U61 (.A2( u0_u3_X_40 ) , .A1( u0_u3_X_41 ) , .ZN( u0_u3_u6_n126 ) );
  NOR2_X1 u0_u3_u6_U62 (.A2( u0_u3_X_39 ) , .A1( u0_u3_X_42 ) , .ZN( u0_u3_u6_n92 ) );
  NOR2_X1 u0_u3_u6_U63 (.A2( u0_u3_X_39 ) , .A1( u0_u3_u6_n156 ) , .ZN( u0_u3_u6_n97 ) );
  NOR2_X1 u0_u3_u6_U64 (.A2( u0_u3_X_38 ) , .A1( u0_u3_u6_n165 ) , .ZN( u0_u3_u6_n95 ) );
  NOR2_X1 u0_u3_u6_U65 (.A2( u0_u3_X_41 ) , .ZN( u0_u3_u6_n111 ) , .A1( u0_u3_u6_n157 ) );
  NOR2_X1 u0_u3_u6_U66 (.A2( u0_u3_X_37 ) , .A1( u0_u3_u6_n162 ) , .ZN( u0_u3_u6_n94 ) );
  NOR2_X1 u0_u3_u6_U67 (.A2( u0_u3_X_37 ) , .A1( u0_u3_X_38 ) , .ZN( u0_u3_u6_n91 ) );
  NAND2_X1 u0_u3_u6_U68 (.A1( u0_u3_X_41 ) , .ZN( u0_u3_u6_n144 ) , .A2( u0_u3_u6_n157 ) );
  NAND2_X1 u0_u3_u6_U69 (.A2( u0_u3_X_40 ) , .A1( u0_u3_X_41 ) , .ZN( u0_u3_u6_n139 ) );
  NOR2_X1 u0_u3_u6_U7 (.A1( u0_u3_u6_n118 ) , .ZN( u0_u3_u6_n143 ) , .A2( u0_u3_u6_n168 ) );
  AND2_X1 u0_u3_u6_U70 (.A1( u0_u3_X_39 ) , .A2( u0_u3_u6_n156 ) , .ZN( u0_u3_u6_n96 ) );
  AND2_X1 u0_u3_u6_U71 (.A1( u0_u3_X_39 ) , .A2( u0_u3_X_42 ) , .ZN( u0_u3_u6_n99 ) );
  INV_X1 u0_u3_u6_U72 (.A( u0_u3_X_40 ) , .ZN( u0_u3_u6_n157 ) );
  INV_X1 u0_u3_u6_U73 (.A( u0_u3_X_37 ) , .ZN( u0_u3_u6_n165 ) );
  INV_X1 u0_u3_u6_U74 (.A( u0_u3_X_38 ) , .ZN( u0_u3_u6_n162 ) );
  INV_X1 u0_u3_u6_U75 (.A( u0_u3_X_42 ) , .ZN( u0_u3_u6_n156 ) );
  NAND4_X1 u0_u3_u6_U76 (.ZN( u0_out3_32 ) , .A4( u0_u3_u6_n103 ) , .A3( u0_u3_u6_n104 ) , .A2( u0_u3_u6_n105 ) , .A1( u0_u3_u6_n106 ) );
  AOI22_X1 u0_u3_u6_U77 (.ZN( u0_u3_u6_n105 ) , .A2( u0_u3_u6_n108 ) , .A1( u0_u3_u6_n118 ) , .B2( u0_u3_u6_n126 ) , .B1( u0_u3_u6_n171 ) );
  AOI22_X1 u0_u3_u6_U78 (.ZN( u0_u3_u6_n104 ) , .A1( u0_u3_u6_n111 ) , .B1( u0_u3_u6_n124 ) , .B2( u0_u3_u6_n151 ) , .A2( u0_u3_u6_n93 ) );
  NAND4_X1 u0_u3_u6_U79 (.ZN( u0_out3_12 ) , .A4( u0_u3_u6_n114 ) , .A3( u0_u3_u6_n115 ) , .A2( u0_u3_u6_n116 ) , .A1( u0_u3_u6_n117 ) );
  AOI21_X1 u0_u3_u6_U8 (.B1( u0_u3_u6_n107 ) , .B2( u0_u3_u6_n132 ) , .A( u0_u3_u6_n158 ) , .ZN( u0_u3_u6_n88 ) );
  OAI22_X1 u0_u3_u6_U80 (.B2( u0_u3_u6_n111 ) , .ZN( u0_u3_u6_n116 ) , .B1( u0_u3_u6_n126 ) , .A2( u0_u3_u6_n164 ) , .A1( u0_u3_u6_n167 ) );
  OAI21_X1 u0_u3_u6_U81 (.A( u0_u3_u6_n108 ) , .ZN( u0_u3_u6_n117 ) , .B2( u0_u3_u6_n141 ) , .B1( u0_u3_u6_n163 ) );
  OAI211_X1 u0_u3_u6_U82 (.ZN( u0_out3_22 ) , .B( u0_u3_u6_n137 ) , .A( u0_u3_u6_n138 ) , .C2( u0_u3_u6_n139 ) , .C1( u0_u3_u6_n140 ) );
  AOI22_X1 u0_u3_u6_U83 (.B1( u0_u3_u6_n124 ) , .A2( u0_u3_u6_n125 ) , .A1( u0_u3_u6_n126 ) , .ZN( u0_u3_u6_n138 ) , .B2( u0_u3_u6_n161 ) );
  AND4_X1 u0_u3_u6_U84 (.A3( u0_u3_u6_n119 ) , .A1( u0_u3_u6_n120 ) , .A4( u0_u3_u6_n129 ) , .ZN( u0_u3_u6_n140 ) , .A2( u0_u3_u6_n143 ) );
  OAI211_X1 u0_u3_u6_U85 (.ZN( u0_out3_7 ) , .B( u0_u3_u6_n153 ) , .C2( u0_u3_u6_n154 ) , .C1( u0_u3_u6_n155 ) , .A( u0_u3_u6_n174 ) );
  NOR3_X1 u0_u3_u6_U86 (.A1( u0_u3_u6_n141 ) , .ZN( u0_u3_u6_n154 ) , .A3( u0_u3_u6_n164 ) , .A2( u0_u3_u6_n171 ) );
  AOI211_X1 u0_u3_u6_U87 (.B( u0_u3_u6_n149 ) , .A( u0_u3_u6_n150 ) , .C2( u0_u3_u6_n151 ) , .C1( u0_u3_u6_n152 ) , .ZN( u0_u3_u6_n153 ) );
  NAND3_X1 u0_u3_u6_U88 (.A2( u0_u3_u6_n123 ) , .ZN( u0_u3_u6_n125 ) , .A1( u0_u3_u6_n130 ) , .A3( u0_u3_u6_n131 ) );
  NAND3_X1 u0_u3_u6_U89 (.A3( u0_u3_u6_n133 ) , .ZN( u0_u3_u6_n141 ) , .A1( u0_u3_u6_n145 ) , .A2( u0_u3_u6_n148 ) );
  AOI21_X1 u0_u3_u6_U9 (.B2( u0_u3_u6_n147 ) , .B1( u0_u3_u6_n148 ) , .ZN( u0_u3_u6_n149 ) , .A( u0_u3_u6_n158 ) );
  NAND3_X1 u0_u3_u6_U90 (.ZN( u0_u3_u6_n101 ) , .A3( u0_u3_u6_n107 ) , .A2( u0_u3_u6_n121 ) , .A1( u0_u3_u6_n127 ) );
  NAND3_X1 u0_u3_u6_U91 (.ZN( u0_u3_u6_n102 ) , .A3( u0_u3_u6_n130 ) , .A2( u0_u3_u6_n145 ) , .A1( u0_u3_u6_n166 ) );
  NAND3_X1 u0_u3_u6_U92 (.A3( u0_u3_u6_n113 ) , .A1( u0_u3_u6_n119 ) , .A2( u0_u3_u6_n123 ) , .ZN( u0_u3_u6_n93 ) );
  NAND3_X1 u0_u3_u6_U93 (.ZN( u0_u3_u6_n142 ) , .A2( u0_u3_u6_n172 ) , .A3( u0_u3_u6_n89 ) , .A1( u0_u3_u6_n90 ) );
  AND3_X1 u0_u3_u7_U10 (.A3( u0_u3_u7_n110 ) , .A2( u0_u3_u7_n127 ) , .A1( u0_u3_u7_n132 ) , .ZN( u0_u3_u7_n92 ) );
  OAI21_X1 u0_u3_u7_U11 (.A( u0_u3_u7_n161 ) , .B1( u0_u3_u7_n168 ) , .B2( u0_u3_u7_n173 ) , .ZN( u0_u3_u7_n91 ) );
  AOI211_X1 u0_u3_u7_U12 (.A( u0_u3_u7_n117 ) , .ZN( u0_u3_u7_n118 ) , .C2( u0_u3_u7_n126 ) , .C1( u0_u3_u7_n177 ) , .B( u0_u3_u7_n180 ) );
  OAI22_X1 u0_u3_u7_U13 (.B1( u0_u3_u7_n115 ) , .ZN( u0_u3_u7_n117 ) , .A2( u0_u3_u7_n133 ) , .A1( u0_u3_u7_n137 ) , .B2( u0_u3_u7_n162 ) );
  INV_X1 u0_u3_u7_U14 (.A( u0_u3_u7_n116 ) , .ZN( u0_u3_u7_n180 ) );
  NOR3_X1 u0_u3_u7_U15 (.ZN( u0_u3_u7_n115 ) , .A3( u0_u3_u7_n145 ) , .A2( u0_u3_u7_n168 ) , .A1( u0_u3_u7_n169 ) );
  OAI211_X1 u0_u3_u7_U16 (.B( u0_u3_u7_n122 ) , .A( u0_u3_u7_n123 ) , .C2( u0_u3_u7_n124 ) , .ZN( u0_u3_u7_n154 ) , .C1( u0_u3_u7_n162 ) );
  AOI222_X1 u0_u3_u7_U17 (.ZN( u0_u3_u7_n122 ) , .C2( u0_u3_u7_n126 ) , .C1( u0_u3_u7_n145 ) , .B1( u0_u3_u7_n161 ) , .A2( u0_u3_u7_n165 ) , .B2( u0_u3_u7_n170 ) , .A1( u0_u3_u7_n176 ) );
  INV_X1 u0_u3_u7_U18 (.A( u0_u3_u7_n133 ) , .ZN( u0_u3_u7_n176 ) );
  NOR3_X1 u0_u3_u7_U19 (.A2( u0_u3_u7_n134 ) , .A1( u0_u3_u7_n135 ) , .ZN( u0_u3_u7_n136 ) , .A3( u0_u3_u7_n171 ) );
  NOR2_X1 u0_u3_u7_U20 (.A1( u0_u3_u7_n130 ) , .A2( u0_u3_u7_n134 ) , .ZN( u0_u3_u7_n153 ) );
  INV_X1 u0_u3_u7_U21 (.A( u0_u3_u7_n101 ) , .ZN( u0_u3_u7_n165 ) );
  NOR2_X1 u0_u3_u7_U22 (.ZN( u0_u3_u7_n111 ) , .A2( u0_u3_u7_n134 ) , .A1( u0_u3_u7_n169 ) );
  AOI21_X1 u0_u3_u7_U23 (.ZN( u0_u3_u7_n104 ) , .B2( u0_u3_u7_n112 ) , .B1( u0_u3_u7_n127 ) , .A( u0_u3_u7_n164 ) );
  AOI21_X1 u0_u3_u7_U24 (.ZN( u0_u3_u7_n106 ) , .B1( u0_u3_u7_n133 ) , .B2( u0_u3_u7_n146 ) , .A( u0_u3_u7_n162 ) );
  AOI21_X1 u0_u3_u7_U25 (.A( u0_u3_u7_n101 ) , .ZN( u0_u3_u7_n107 ) , .B2( u0_u3_u7_n128 ) , .B1( u0_u3_u7_n175 ) );
  INV_X1 u0_u3_u7_U26 (.A( u0_u3_u7_n138 ) , .ZN( u0_u3_u7_n171 ) );
  INV_X1 u0_u3_u7_U27 (.A( u0_u3_u7_n131 ) , .ZN( u0_u3_u7_n177 ) );
  INV_X1 u0_u3_u7_U28 (.A( u0_u3_u7_n110 ) , .ZN( u0_u3_u7_n174 ) );
  NAND2_X1 u0_u3_u7_U29 (.A1( u0_u3_u7_n129 ) , .A2( u0_u3_u7_n132 ) , .ZN( u0_u3_u7_n149 ) );
  OAI21_X1 u0_u3_u7_U3 (.ZN( u0_u3_u7_n159 ) , .A( u0_u3_u7_n165 ) , .B2( u0_u3_u7_n171 ) , .B1( u0_u3_u7_n174 ) );
  NAND2_X1 u0_u3_u7_U30 (.A1( u0_u3_u7_n113 ) , .A2( u0_u3_u7_n124 ) , .ZN( u0_u3_u7_n130 ) );
  INV_X1 u0_u3_u7_U31 (.A( u0_u3_u7_n112 ) , .ZN( u0_u3_u7_n173 ) );
  INV_X1 u0_u3_u7_U32 (.A( u0_u3_u7_n128 ) , .ZN( u0_u3_u7_n168 ) );
  INV_X1 u0_u3_u7_U33 (.A( u0_u3_u7_n148 ) , .ZN( u0_u3_u7_n169 ) );
  INV_X1 u0_u3_u7_U34 (.A( u0_u3_u7_n127 ) , .ZN( u0_u3_u7_n179 ) );
  NOR2_X1 u0_u3_u7_U35 (.ZN( u0_u3_u7_n101 ) , .A2( u0_u3_u7_n150 ) , .A1( u0_u3_u7_n156 ) );
  AOI211_X1 u0_u3_u7_U36 (.B( u0_u3_u7_n154 ) , .A( u0_u3_u7_n155 ) , .C1( u0_u3_u7_n156 ) , .ZN( u0_u3_u7_n157 ) , .C2( u0_u3_u7_n172 ) );
  INV_X1 u0_u3_u7_U37 (.A( u0_u3_u7_n153 ) , .ZN( u0_u3_u7_n172 ) );
  AOI211_X1 u0_u3_u7_U38 (.B( u0_u3_u7_n139 ) , .A( u0_u3_u7_n140 ) , .C2( u0_u3_u7_n141 ) , .ZN( u0_u3_u7_n142 ) , .C1( u0_u3_u7_n156 ) );
  NAND4_X1 u0_u3_u7_U39 (.A3( u0_u3_u7_n127 ) , .A2( u0_u3_u7_n128 ) , .A1( u0_u3_u7_n129 ) , .ZN( u0_u3_u7_n141 ) , .A4( u0_u3_u7_n147 ) );
  INV_X1 u0_u3_u7_U4 (.A( u0_u3_u7_n111 ) , .ZN( u0_u3_u7_n170 ) );
  AOI21_X1 u0_u3_u7_U40 (.A( u0_u3_u7_n137 ) , .B1( u0_u3_u7_n138 ) , .ZN( u0_u3_u7_n139 ) , .B2( u0_u3_u7_n146 ) );
  OAI22_X1 u0_u3_u7_U41 (.B1( u0_u3_u7_n136 ) , .ZN( u0_u3_u7_n140 ) , .A1( u0_u3_u7_n153 ) , .B2( u0_u3_u7_n162 ) , .A2( u0_u3_u7_n164 ) );
  AOI21_X1 u0_u3_u7_U42 (.ZN( u0_u3_u7_n123 ) , .B1( u0_u3_u7_n165 ) , .B2( u0_u3_u7_n177 ) , .A( u0_u3_u7_n97 ) );
  AOI21_X1 u0_u3_u7_U43 (.B2( u0_u3_u7_n113 ) , .B1( u0_u3_u7_n124 ) , .A( u0_u3_u7_n125 ) , .ZN( u0_u3_u7_n97 ) );
  INV_X1 u0_u3_u7_U44 (.A( u0_u3_u7_n125 ) , .ZN( u0_u3_u7_n161 ) );
  INV_X1 u0_u3_u7_U45 (.A( u0_u3_u7_n152 ) , .ZN( u0_u3_u7_n162 ) );
  AOI22_X1 u0_u3_u7_U46 (.A2( u0_u3_u7_n114 ) , .ZN( u0_u3_u7_n119 ) , .B1( u0_u3_u7_n130 ) , .A1( u0_u3_u7_n156 ) , .B2( u0_u3_u7_n165 ) );
  NAND2_X1 u0_u3_u7_U47 (.A2( u0_u3_u7_n112 ) , .ZN( u0_u3_u7_n114 ) , .A1( u0_u3_u7_n175 ) );
  AND2_X1 u0_u3_u7_U48 (.ZN( u0_u3_u7_n145 ) , .A2( u0_u3_u7_n98 ) , .A1( u0_u3_u7_n99 ) );
  NOR2_X1 u0_u3_u7_U49 (.ZN( u0_u3_u7_n137 ) , .A1( u0_u3_u7_n150 ) , .A2( u0_u3_u7_n161 ) );
  INV_X1 u0_u3_u7_U5 (.A( u0_u3_u7_n149 ) , .ZN( u0_u3_u7_n175 ) );
  AOI21_X1 u0_u3_u7_U50 (.ZN( u0_u3_u7_n105 ) , .B2( u0_u3_u7_n110 ) , .A( u0_u3_u7_n125 ) , .B1( u0_u3_u7_n147 ) );
  NAND2_X1 u0_u3_u7_U51 (.ZN( u0_u3_u7_n146 ) , .A1( u0_u3_u7_n95 ) , .A2( u0_u3_u7_n98 ) );
  NAND2_X1 u0_u3_u7_U52 (.A2( u0_u3_u7_n103 ) , .ZN( u0_u3_u7_n147 ) , .A1( u0_u3_u7_n93 ) );
  NAND2_X1 u0_u3_u7_U53 (.A1( u0_u3_u7_n103 ) , .ZN( u0_u3_u7_n127 ) , .A2( u0_u3_u7_n99 ) );
  OR2_X1 u0_u3_u7_U54 (.ZN( u0_u3_u7_n126 ) , .A2( u0_u3_u7_n152 ) , .A1( u0_u3_u7_n156 ) );
  NAND2_X1 u0_u3_u7_U55 (.A2( u0_u3_u7_n102 ) , .A1( u0_u3_u7_n103 ) , .ZN( u0_u3_u7_n133 ) );
  NAND2_X1 u0_u3_u7_U56 (.ZN( u0_u3_u7_n112 ) , .A2( u0_u3_u7_n96 ) , .A1( u0_u3_u7_n99 ) );
  NAND2_X1 u0_u3_u7_U57 (.A2( u0_u3_u7_n102 ) , .ZN( u0_u3_u7_n128 ) , .A1( u0_u3_u7_n98 ) );
  NAND2_X1 u0_u3_u7_U58 (.A1( u0_u3_u7_n100 ) , .ZN( u0_u3_u7_n113 ) , .A2( u0_u3_u7_n93 ) );
  NAND2_X1 u0_u3_u7_U59 (.A2( u0_u3_u7_n102 ) , .ZN( u0_u3_u7_n124 ) , .A1( u0_u3_u7_n96 ) );
  INV_X1 u0_u3_u7_U6 (.A( u0_u3_u7_n154 ) , .ZN( u0_u3_u7_n178 ) );
  NAND2_X1 u0_u3_u7_U60 (.ZN( u0_u3_u7_n110 ) , .A1( u0_u3_u7_n95 ) , .A2( u0_u3_u7_n96 ) );
  INV_X1 u0_u3_u7_U61 (.A( u0_u3_u7_n150 ) , .ZN( u0_u3_u7_n164 ) );
  AND2_X1 u0_u3_u7_U62 (.ZN( u0_u3_u7_n134 ) , .A1( u0_u3_u7_n93 ) , .A2( u0_u3_u7_n98 ) );
  NAND2_X1 u0_u3_u7_U63 (.A1( u0_u3_u7_n100 ) , .A2( u0_u3_u7_n102 ) , .ZN( u0_u3_u7_n129 ) );
  NAND2_X1 u0_u3_u7_U64 (.A2( u0_u3_u7_n103 ) , .ZN( u0_u3_u7_n131 ) , .A1( u0_u3_u7_n95 ) );
  NAND2_X1 u0_u3_u7_U65 (.A1( u0_u3_u7_n100 ) , .ZN( u0_u3_u7_n138 ) , .A2( u0_u3_u7_n99 ) );
  NAND2_X1 u0_u3_u7_U66 (.ZN( u0_u3_u7_n132 ) , .A1( u0_u3_u7_n93 ) , .A2( u0_u3_u7_n96 ) );
  NAND2_X1 u0_u3_u7_U67 (.A1( u0_u3_u7_n100 ) , .ZN( u0_u3_u7_n148 ) , .A2( u0_u3_u7_n95 ) );
  NOR2_X1 u0_u3_u7_U68 (.A2( u0_u3_X_47 ) , .ZN( u0_u3_u7_n150 ) , .A1( u0_u3_u7_n163 ) );
  NOR2_X1 u0_u3_u7_U69 (.A2( u0_u3_X_43 ) , .A1( u0_u3_X_44 ) , .ZN( u0_u3_u7_n103 ) );
  AOI211_X1 u0_u3_u7_U7 (.ZN( u0_u3_u7_n116 ) , .A( u0_u3_u7_n155 ) , .C1( u0_u3_u7_n161 ) , .C2( u0_u3_u7_n171 ) , .B( u0_u3_u7_n94 ) );
  NOR2_X1 u0_u3_u7_U70 (.A2( u0_u3_X_48 ) , .A1( u0_u3_u7_n166 ) , .ZN( u0_u3_u7_n95 ) );
  NOR2_X1 u0_u3_u7_U71 (.A2( u0_u3_X_45 ) , .A1( u0_u3_X_48 ) , .ZN( u0_u3_u7_n99 ) );
  NOR2_X1 u0_u3_u7_U72 (.A2( u0_u3_X_44 ) , .A1( u0_u3_u7_n167 ) , .ZN( u0_u3_u7_n98 ) );
  NOR2_X1 u0_u3_u7_U73 (.A2( u0_u3_X_46 ) , .A1( u0_u3_X_47 ) , .ZN( u0_u3_u7_n152 ) );
  AND2_X1 u0_u3_u7_U74 (.A1( u0_u3_X_47 ) , .ZN( u0_u3_u7_n156 ) , .A2( u0_u3_u7_n163 ) );
  NAND2_X1 u0_u3_u7_U75 (.A2( u0_u3_X_46 ) , .A1( u0_u3_X_47 ) , .ZN( u0_u3_u7_n125 ) );
  AND2_X1 u0_u3_u7_U76 (.A2( u0_u3_X_45 ) , .A1( u0_u3_X_48 ) , .ZN( u0_u3_u7_n102 ) );
  AND2_X1 u0_u3_u7_U77 (.A2( u0_u3_X_43 ) , .A1( u0_u3_X_44 ) , .ZN( u0_u3_u7_n96 ) );
  AND2_X1 u0_u3_u7_U78 (.A1( u0_u3_X_44 ) , .ZN( u0_u3_u7_n100 ) , .A2( u0_u3_u7_n167 ) );
  AND2_X1 u0_u3_u7_U79 (.A1( u0_u3_X_48 ) , .A2( u0_u3_u7_n166 ) , .ZN( u0_u3_u7_n93 ) );
  OAI222_X1 u0_u3_u7_U8 (.C2( u0_u3_u7_n101 ) , .B2( u0_u3_u7_n111 ) , .A1( u0_u3_u7_n113 ) , .C1( u0_u3_u7_n146 ) , .A2( u0_u3_u7_n162 ) , .B1( u0_u3_u7_n164 ) , .ZN( u0_u3_u7_n94 ) );
  INV_X1 u0_u3_u7_U80 (.A( u0_u3_X_46 ) , .ZN( u0_u3_u7_n163 ) );
  INV_X1 u0_u3_u7_U81 (.A( u0_u3_X_43 ) , .ZN( u0_u3_u7_n167 ) );
  INV_X1 u0_u3_u7_U82 (.A( u0_u3_X_45 ) , .ZN( u0_u3_u7_n166 ) );
  NAND4_X1 u0_u3_u7_U83 (.ZN( u0_out3_5 ) , .A4( u0_u3_u7_n108 ) , .A3( u0_u3_u7_n109 ) , .A1( u0_u3_u7_n116 ) , .A2( u0_u3_u7_n123 ) );
  AOI22_X1 u0_u3_u7_U84 (.ZN( u0_u3_u7_n109 ) , .A2( u0_u3_u7_n126 ) , .B2( u0_u3_u7_n145 ) , .B1( u0_u3_u7_n156 ) , .A1( u0_u3_u7_n171 ) );
  NOR4_X1 u0_u3_u7_U85 (.A4( u0_u3_u7_n104 ) , .A3( u0_u3_u7_n105 ) , .A2( u0_u3_u7_n106 ) , .A1( u0_u3_u7_n107 ) , .ZN( u0_u3_u7_n108 ) );
  NAND4_X1 u0_u3_u7_U86 (.ZN( u0_out3_27 ) , .A4( u0_u3_u7_n118 ) , .A3( u0_u3_u7_n119 ) , .A2( u0_u3_u7_n120 ) , .A1( u0_u3_u7_n121 ) );
  OAI21_X1 u0_u3_u7_U87 (.ZN( u0_u3_u7_n121 ) , .B2( u0_u3_u7_n145 ) , .A( u0_u3_u7_n150 ) , .B1( u0_u3_u7_n174 ) );
  OAI21_X1 u0_u3_u7_U88 (.ZN( u0_u3_u7_n120 ) , .A( u0_u3_u7_n161 ) , .B2( u0_u3_u7_n170 ) , .B1( u0_u3_u7_n179 ) );
  NAND4_X1 u0_u3_u7_U89 (.ZN( u0_out3_21 ) , .A4( u0_u3_u7_n157 ) , .A3( u0_u3_u7_n158 ) , .A2( u0_u3_u7_n159 ) , .A1( u0_u3_u7_n160 ) );
  OAI221_X1 u0_u3_u7_U9 (.C1( u0_u3_u7_n101 ) , .C2( u0_u3_u7_n147 ) , .ZN( u0_u3_u7_n155 ) , .B2( u0_u3_u7_n162 ) , .A( u0_u3_u7_n91 ) , .B1( u0_u3_u7_n92 ) );
  OAI21_X1 u0_u3_u7_U90 (.B1( u0_u3_u7_n145 ) , .ZN( u0_u3_u7_n160 ) , .A( u0_u3_u7_n161 ) , .B2( u0_u3_u7_n177 ) );
  AOI22_X1 u0_u3_u7_U91 (.B2( u0_u3_u7_n149 ) , .B1( u0_u3_u7_n150 ) , .A2( u0_u3_u7_n151 ) , .A1( u0_u3_u7_n152 ) , .ZN( u0_u3_u7_n158 ) );
  NAND4_X1 u0_u3_u7_U92 (.ZN( u0_out3_15 ) , .A4( u0_u3_u7_n142 ) , .A3( u0_u3_u7_n143 ) , .A2( u0_u3_u7_n144 ) , .A1( u0_u3_u7_n178 ) );
  OR2_X1 u0_u3_u7_U93 (.A2( u0_u3_u7_n125 ) , .A1( u0_u3_u7_n129 ) , .ZN( u0_u3_u7_n144 ) );
  AOI22_X1 u0_u3_u7_U94 (.A2( u0_u3_u7_n126 ) , .ZN( u0_u3_u7_n143 ) , .B2( u0_u3_u7_n165 ) , .B1( u0_u3_u7_n173 ) , .A1( u0_u3_u7_n174 ) );
  NAND3_X1 u0_u3_u7_U95 (.A3( u0_u3_u7_n146 ) , .A2( u0_u3_u7_n147 ) , .A1( u0_u3_u7_n148 ) , .ZN( u0_u3_u7_n151 ) );
  NAND3_X1 u0_u3_u7_U96 (.A3( u0_u3_u7_n131 ) , .A2( u0_u3_u7_n132 ) , .A1( u0_u3_u7_n133 ) , .ZN( u0_u3_u7_n135 ) );
  XOR2_X1 u0_u4_U2 (.B( u0_K5_8 ) , .A( u0_R3_5 ) , .Z( u0_u4_X_8 ) );
  XOR2_X1 u0_u4_U20 (.B( u0_K5_36 ) , .A( u0_R3_25 ) , .Z( u0_u4_X_36 ) );
  XOR2_X1 u0_u4_U21 (.B( u0_K5_35 ) , .A( u0_R3_24 ) , .Z( u0_u4_X_35 ) );
  XOR2_X1 u0_u4_U23 (.B( u0_K5_33 ) , .A( u0_R3_22 ) , .Z( u0_u4_X_33 ) );
  XOR2_X1 u0_u4_U25 (.B( u0_K5_31 ) , .A( u0_R3_20 ) , .Z( u0_u4_X_31 ) );
  XOR2_X1 u0_u4_U28 (.B( u0_K5_29 ) , .A( u0_R3_20 ) , .Z( u0_u4_X_29 ) );
  XOR2_X1 u0_u4_U30 (.B( u0_K5_27 ) , .A( u0_R3_18 ) , .Z( u0_u4_X_27 ) );
  XOR2_X1 u0_u4_U31 (.B( u0_K5_26 ) , .A( u0_R3_17 ) , .Z( u0_u4_X_26 ) );
  XOR2_X1 u0_u4_U33 (.B( u0_K5_24 ) , .A( u0_R3_17 ) , .Z( u0_u4_X_24 ) );
  XOR2_X1 u0_u4_U35 (.B( u0_K5_22 ) , .A( u0_R3_15 ) , .Z( u0_u4_X_22 ) );
  XOR2_X1 u0_u4_U37 (.B( u0_K5_20 ) , .A( u0_R3_13 ) , .Z( u0_u4_X_20 ) );
  XOR2_X1 u0_u4_U38 (.B( u0_K5_1 ) , .A( u0_R3_32 ) , .Z( u0_u4_X_1 ) );
  XOR2_X1 u0_u4_U4 (.B( u0_K5_6 ) , .A( u0_R3_5 ) , .Z( u0_u4_X_6 ) );
  XOR2_X1 u0_u4_U40 (.B( u0_K5_18 ) , .A( u0_R3_13 ) , .Z( u0_u4_X_18 ) );
  XOR2_X1 u0_u4_U8 (.B( u0_K5_47 ) , .A( u0_R3_32 ) , .Z( u0_u4_X_47 ) );
  AND3_X1 u0_u4_u0_U10 (.A2( u0_u4_u0_n112 ) , .ZN( u0_u4_u0_n127 ) , .A3( u0_u4_u0_n130 ) , .A1( u0_u4_u0_n148 ) );
  NAND2_X1 u0_u4_u0_U11 (.ZN( u0_u4_u0_n113 ) , .A1( u0_u4_u0_n139 ) , .A2( u0_u4_u0_n149 ) );
  AND2_X1 u0_u4_u0_U12 (.ZN( u0_u4_u0_n107 ) , .A1( u0_u4_u0_n130 ) , .A2( u0_u4_u0_n140 ) );
  AND2_X1 u0_u4_u0_U13 (.A2( u0_u4_u0_n129 ) , .A1( u0_u4_u0_n130 ) , .ZN( u0_u4_u0_n151 ) );
  AND2_X1 u0_u4_u0_U14 (.A1( u0_u4_u0_n108 ) , .A2( u0_u4_u0_n125 ) , .ZN( u0_u4_u0_n145 ) );
  INV_X1 u0_u4_u0_U15 (.A( u0_u4_u0_n143 ) , .ZN( u0_u4_u0_n173 ) );
  NOR2_X1 u0_u4_u0_U16 (.A2( u0_u4_u0_n136 ) , .ZN( u0_u4_u0_n147 ) , .A1( u0_u4_u0_n160 ) );
  INV_X1 u0_u4_u0_U17 (.ZN( u0_u4_u0_n172 ) , .A( u0_u4_u0_n88 ) );
  OAI222_X1 u0_u4_u0_U18 (.C1( u0_u4_u0_n108 ) , .A1( u0_u4_u0_n125 ) , .B2( u0_u4_u0_n128 ) , .B1( u0_u4_u0_n144 ) , .A2( u0_u4_u0_n158 ) , .C2( u0_u4_u0_n161 ) , .ZN( u0_u4_u0_n88 ) );
  AOI21_X1 u0_u4_u0_U19 (.B1( u0_u4_u0_n103 ) , .ZN( u0_u4_u0_n132 ) , .A( u0_u4_u0_n165 ) , .B2( u0_u4_u0_n93 ) );
  INV_X1 u0_u4_u0_U20 (.A( u0_u4_u0_n142 ) , .ZN( u0_u4_u0_n165 ) );
  OAI221_X1 u0_u4_u0_U21 (.C1( u0_u4_u0_n112 ) , .ZN( u0_u4_u0_n120 ) , .B1( u0_u4_u0_n138 ) , .B2( u0_u4_u0_n141 ) , .C2( u0_u4_u0_n147 ) , .A( u0_u4_u0_n172 ) );
  AOI211_X1 u0_u4_u0_U22 (.B( u0_u4_u0_n115 ) , .A( u0_u4_u0_n116 ) , .C2( u0_u4_u0_n117 ) , .C1( u0_u4_u0_n118 ) , .ZN( u0_u4_u0_n119 ) );
  OAI22_X1 u0_u4_u0_U23 (.B1( u0_u4_u0_n125 ) , .ZN( u0_u4_u0_n126 ) , .A1( u0_u4_u0_n138 ) , .A2( u0_u4_u0_n146 ) , .B2( u0_u4_u0_n147 ) );
  OAI22_X1 u0_u4_u0_U24 (.B1( u0_u4_u0_n131 ) , .A1( u0_u4_u0_n144 ) , .B2( u0_u4_u0_n147 ) , .A2( u0_u4_u0_n90 ) , .ZN( u0_u4_u0_n91 ) );
  AND3_X1 u0_u4_u0_U25 (.A3( u0_u4_u0_n121 ) , .A2( u0_u4_u0_n125 ) , .A1( u0_u4_u0_n148 ) , .ZN( u0_u4_u0_n90 ) );
  INV_X1 u0_u4_u0_U26 (.A( u0_u4_u0_n136 ) , .ZN( u0_u4_u0_n161 ) );
  AOI22_X1 u0_u4_u0_U27 (.B2( u0_u4_u0_n109 ) , .A2( u0_u4_u0_n110 ) , .ZN( u0_u4_u0_n111 ) , .B1( u0_u4_u0_n118 ) , .A1( u0_u4_u0_n160 ) );
  INV_X1 u0_u4_u0_U28 (.A( u0_u4_u0_n118 ) , .ZN( u0_u4_u0_n158 ) );
  AOI21_X1 u0_u4_u0_U29 (.ZN( u0_u4_u0_n104 ) , .B1( u0_u4_u0_n107 ) , .B2( u0_u4_u0_n141 ) , .A( u0_u4_u0_n144 ) );
  INV_X1 u0_u4_u0_U3 (.A( u0_u4_u0_n113 ) , .ZN( u0_u4_u0_n166 ) );
  AOI21_X1 u0_u4_u0_U30 (.B1( u0_u4_u0_n127 ) , .B2( u0_u4_u0_n129 ) , .A( u0_u4_u0_n138 ) , .ZN( u0_u4_u0_n96 ) );
  AOI21_X1 u0_u4_u0_U31 (.ZN( u0_u4_u0_n116 ) , .B2( u0_u4_u0_n142 ) , .A( u0_u4_u0_n144 ) , .B1( u0_u4_u0_n166 ) );
  NAND2_X1 u0_u4_u0_U32 (.A1( u0_u4_u0_n102 ) , .ZN( u0_u4_u0_n128 ) , .A2( u0_u4_u0_n95 ) );
  NAND2_X1 u0_u4_u0_U33 (.A1( u0_u4_u0_n100 ) , .A2( u0_u4_u0_n103 ) , .ZN( u0_u4_u0_n125 ) );
  NAND2_X1 u0_u4_u0_U34 (.ZN( u0_u4_u0_n148 ) , .A1( u0_u4_u0_n93 ) , .A2( u0_u4_u0_n95 ) );
  NAND2_X1 u0_u4_u0_U35 (.A1( u0_u4_u0_n101 ) , .A2( u0_u4_u0_n102 ) , .ZN( u0_u4_u0_n150 ) );
  INV_X1 u0_u4_u0_U36 (.A( u0_u4_u0_n138 ) , .ZN( u0_u4_u0_n160 ) );
  NAND2_X1 u0_u4_u0_U37 (.A1( u0_u4_u0_n100 ) , .ZN( u0_u4_u0_n129 ) , .A2( u0_u4_u0_n95 ) );
  NAND2_X1 u0_u4_u0_U38 (.A2( u0_u4_u0_n102 ) , .A1( u0_u4_u0_n103 ) , .ZN( u0_u4_u0_n149 ) );
  NAND2_X1 u0_u4_u0_U39 (.A2( u0_u4_u0_n100 ) , .A1( u0_u4_u0_n101 ) , .ZN( u0_u4_u0_n139 ) );
  AOI21_X1 u0_u4_u0_U4 (.B1( u0_u4_u0_n114 ) , .ZN( u0_u4_u0_n115 ) , .B2( u0_u4_u0_n129 ) , .A( u0_u4_u0_n161 ) );
  NAND2_X1 u0_u4_u0_U40 (.A2( u0_u4_u0_n100 ) , .ZN( u0_u4_u0_n131 ) , .A1( u0_u4_u0_n92 ) );
  NAND2_X1 u0_u4_u0_U41 (.A2( u0_u4_u0_n102 ) , .ZN( u0_u4_u0_n114 ) , .A1( u0_u4_u0_n92 ) );
  NAND2_X1 u0_u4_u0_U42 (.A2( u0_u4_u0_n101 ) , .ZN( u0_u4_u0_n121 ) , .A1( u0_u4_u0_n93 ) );
  NAND2_X1 u0_u4_u0_U43 (.ZN( u0_u4_u0_n112 ) , .A2( u0_u4_u0_n92 ) , .A1( u0_u4_u0_n93 ) );
  OR3_X1 u0_u4_u0_U44 (.A3( u0_u4_u0_n152 ) , .A2( u0_u4_u0_n153 ) , .A1( u0_u4_u0_n154 ) , .ZN( u0_u4_u0_n155 ) );
  AOI21_X1 u0_u4_u0_U45 (.B2( u0_u4_u0_n150 ) , .B1( u0_u4_u0_n151 ) , .ZN( u0_u4_u0_n152 ) , .A( u0_u4_u0_n158 ) );
  AOI21_X1 u0_u4_u0_U46 (.A( u0_u4_u0_n144 ) , .B2( u0_u4_u0_n145 ) , .B1( u0_u4_u0_n146 ) , .ZN( u0_u4_u0_n154 ) );
  AOI21_X1 u0_u4_u0_U47 (.A( u0_u4_u0_n147 ) , .B2( u0_u4_u0_n148 ) , .B1( u0_u4_u0_n149 ) , .ZN( u0_u4_u0_n153 ) );
  INV_X1 u0_u4_u0_U48 (.ZN( u0_u4_u0_n171 ) , .A( u0_u4_u0_n99 ) );
  OAI211_X1 u0_u4_u0_U49 (.C2( u0_u4_u0_n140 ) , .C1( u0_u4_u0_n161 ) , .A( u0_u4_u0_n169 ) , .B( u0_u4_u0_n98 ) , .ZN( u0_u4_u0_n99 ) );
  AOI21_X1 u0_u4_u0_U5 (.B2( u0_u4_u0_n131 ) , .ZN( u0_u4_u0_n134 ) , .B1( u0_u4_u0_n151 ) , .A( u0_u4_u0_n158 ) );
  AOI211_X1 u0_u4_u0_U50 (.C1( u0_u4_u0_n118 ) , .A( u0_u4_u0_n123 ) , .B( u0_u4_u0_n96 ) , .C2( u0_u4_u0_n97 ) , .ZN( u0_u4_u0_n98 ) );
  INV_X1 u0_u4_u0_U51 (.ZN( u0_u4_u0_n169 ) , .A( u0_u4_u0_n91 ) );
  NOR2_X1 u0_u4_u0_U52 (.A2( u0_u4_X_6 ) , .ZN( u0_u4_u0_n100 ) , .A1( u0_u4_u0_n162 ) );
  NOR2_X1 u0_u4_u0_U53 (.A2( u0_u4_X_4 ) , .A1( u0_u4_X_5 ) , .ZN( u0_u4_u0_n118 ) );
  NOR2_X1 u0_u4_u0_U54 (.A2( u0_u4_X_2 ) , .ZN( u0_u4_u0_n103 ) , .A1( u0_u4_u0_n164 ) );
  NOR2_X1 u0_u4_u0_U55 (.A2( u0_u4_X_1 ) , .A1( u0_u4_X_2 ) , .ZN( u0_u4_u0_n92 ) );
  NOR2_X1 u0_u4_u0_U56 (.A2( u0_u4_X_1 ) , .ZN( u0_u4_u0_n101 ) , .A1( u0_u4_u0_n163 ) );
  NAND2_X1 u0_u4_u0_U57 (.A2( u0_u4_X_4 ) , .A1( u0_u4_X_5 ) , .ZN( u0_u4_u0_n144 ) );
  NOR2_X1 u0_u4_u0_U58 (.A2( u0_u4_X_5 ) , .ZN( u0_u4_u0_n136 ) , .A1( u0_u4_u0_n159 ) );
  NAND2_X1 u0_u4_u0_U59 (.A1( u0_u4_X_5 ) , .ZN( u0_u4_u0_n138 ) , .A2( u0_u4_u0_n159 ) );
  NOR2_X1 u0_u4_u0_U6 (.A1( u0_u4_u0_n108 ) , .ZN( u0_u4_u0_n123 ) , .A2( u0_u4_u0_n158 ) );
  AND2_X1 u0_u4_u0_U60 (.A2( u0_u4_X_3 ) , .A1( u0_u4_X_6 ) , .ZN( u0_u4_u0_n102 ) );
  AND2_X1 u0_u4_u0_U61 (.A1( u0_u4_X_6 ) , .A2( u0_u4_u0_n162 ) , .ZN( u0_u4_u0_n93 ) );
  INV_X1 u0_u4_u0_U62 (.A( u0_u4_X_4 ) , .ZN( u0_u4_u0_n159 ) );
  INV_X1 u0_u4_u0_U63 (.A( u0_u4_X_1 ) , .ZN( u0_u4_u0_n164 ) );
  INV_X1 u0_u4_u0_U64 (.A( u0_u4_X_2 ) , .ZN( u0_u4_u0_n163 ) );
  INV_X1 u0_u4_u0_U65 (.A( u0_u4_X_3 ) , .ZN( u0_u4_u0_n162 ) );
  INV_X1 u0_u4_u0_U66 (.A( u0_u4_u0_n126 ) , .ZN( u0_u4_u0_n168 ) );
  AOI211_X1 u0_u4_u0_U67 (.B( u0_u4_u0_n133 ) , .A( u0_u4_u0_n134 ) , .C2( u0_u4_u0_n135 ) , .C1( u0_u4_u0_n136 ) , .ZN( u0_u4_u0_n137 ) );
  OR4_X1 u0_u4_u0_U68 (.ZN( u0_out4_17 ) , .A4( u0_u4_u0_n122 ) , .A2( u0_u4_u0_n123 ) , .A1( u0_u4_u0_n124 ) , .A3( u0_u4_u0_n170 ) );
  AOI21_X1 u0_u4_u0_U69 (.B2( u0_u4_u0_n107 ) , .ZN( u0_u4_u0_n124 ) , .B1( u0_u4_u0_n128 ) , .A( u0_u4_u0_n161 ) );
  OAI21_X1 u0_u4_u0_U7 (.B1( u0_u4_u0_n150 ) , .B2( u0_u4_u0_n158 ) , .A( u0_u4_u0_n172 ) , .ZN( u0_u4_u0_n89 ) );
  INV_X1 u0_u4_u0_U70 (.A( u0_u4_u0_n111 ) , .ZN( u0_u4_u0_n170 ) );
  OR4_X1 u0_u4_u0_U71 (.ZN( u0_out4_31 ) , .A4( u0_u4_u0_n155 ) , .A2( u0_u4_u0_n156 ) , .A1( u0_u4_u0_n157 ) , .A3( u0_u4_u0_n173 ) );
  AOI21_X1 u0_u4_u0_U72 (.A( u0_u4_u0_n138 ) , .B2( u0_u4_u0_n139 ) , .B1( u0_u4_u0_n140 ) , .ZN( u0_u4_u0_n157 ) );
  AOI21_X1 u0_u4_u0_U73 (.B2( u0_u4_u0_n141 ) , .B1( u0_u4_u0_n142 ) , .ZN( u0_u4_u0_n156 ) , .A( u0_u4_u0_n161 ) );
  INV_X1 u0_u4_u0_U74 (.ZN( u0_u4_u0_n174 ) , .A( u0_u4_u0_n89 ) );
  AOI211_X1 u0_u4_u0_U75 (.B( u0_u4_u0_n104 ) , .A( u0_u4_u0_n105 ) , .ZN( u0_u4_u0_n106 ) , .C2( u0_u4_u0_n113 ) , .C1( u0_u4_u0_n160 ) );
  NOR2_X1 u0_u4_u0_U76 (.A2( u0_u4_X_3 ) , .A1( u0_u4_X_6 ) , .ZN( u0_u4_u0_n94 ) );
  NOR2_X1 u0_u4_u0_U77 (.A1( u0_u4_u0_n163 ) , .A2( u0_u4_u0_n164 ) , .ZN( u0_u4_u0_n95 ) );
  OAI221_X1 u0_u4_u0_U78 (.C1( u0_u4_u0_n121 ) , .ZN( u0_u4_u0_n122 ) , .B2( u0_u4_u0_n127 ) , .A( u0_u4_u0_n143 ) , .B1( u0_u4_u0_n144 ) , .C2( u0_u4_u0_n147 ) );
  NOR2_X1 u0_u4_u0_U79 (.A1( u0_u4_u0_n120 ) , .ZN( u0_u4_u0_n143 ) , .A2( u0_u4_u0_n167 ) );
  AND2_X1 u0_u4_u0_U8 (.A1( u0_u4_u0_n114 ) , .A2( u0_u4_u0_n121 ) , .ZN( u0_u4_u0_n146 ) );
  AOI21_X1 u0_u4_u0_U80 (.B1( u0_u4_u0_n132 ) , .ZN( u0_u4_u0_n133 ) , .A( u0_u4_u0_n144 ) , .B2( u0_u4_u0_n166 ) );
  OAI22_X1 u0_u4_u0_U81 (.ZN( u0_u4_u0_n105 ) , .A2( u0_u4_u0_n132 ) , .B1( u0_u4_u0_n146 ) , .A1( u0_u4_u0_n147 ) , .B2( u0_u4_u0_n161 ) );
  NAND2_X1 u0_u4_u0_U82 (.ZN( u0_u4_u0_n110 ) , .A2( u0_u4_u0_n132 ) , .A1( u0_u4_u0_n145 ) );
  INV_X1 u0_u4_u0_U83 (.A( u0_u4_u0_n119 ) , .ZN( u0_u4_u0_n167 ) );
  NAND2_X1 u0_u4_u0_U84 (.A2( u0_u4_u0_n103 ) , .ZN( u0_u4_u0_n140 ) , .A1( u0_u4_u0_n94 ) );
  NAND2_X1 u0_u4_u0_U85 (.A1( u0_u4_u0_n101 ) , .ZN( u0_u4_u0_n130 ) , .A2( u0_u4_u0_n94 ) );
  NAND2_X1 u0_u4_u0_U86 (.ZN( u0_u4_u0_n108 ) , .A1( u0_u4_u0_n92 ) , .A2( u0_u4_u0_n94 ) );
  NAND2_X1 u0_u4_u0_U87 (.ZN( u0_u4_u0_n142 ) , .A1( u0_u4_u0_n94 ) , .A2( u0_u4_u0_n95 ) );
  NAND3_X1 u0_u4_u0_U88 (.ZN( u0_out4_23 ) , .A3( u0_u4_u0_n137 ) , .A1( u0_u4_u0_n168 ) , .A2( u0_u4_u0_n171 ) );
  NAND3_X1 u0_u4_u0_U89 (.A3( u0_u4_u0_n127 ) , .A2( u0_u4_u0_n128 ) , .ZN( u0_u4_u0_n135 ) , .A1( u0_u4_u0_n150 ) );
  AND2_X1 u0_u4_u0_U9 (.A1( u0_u4_u0_n131 ) , .ZN( u0_u4_u0_n141 ) , .A2( u0_u4_u0_n150 ) );
  NAND3_X1 u0_u4_u0_U90 (.ZN( u0_u4_u0_n117 ) , .A3( u0_u4_u0_n132 ) , .A2( u0_u4_u0_n139 ) , .A1( u0_u4_u0_n148 ) );
  NAND3_X1 u0_u4_u0_U91 (.ZN( u0_u4_u0_n109 ) , .A2( u0_u4_u0_n114 ) , .A3( u0_u4_u0_n140 ) , .A1( u0_u4_u0_n149 ) );
  NAND3_X1 u0_u4_u0_U92 (.ZN( u0_out4_9 ) , .A3( u0_u4_u0_n106 ) , .A2( u0_u4_u0_n171 ) , .A1( u0_u4_u0_n174 ) );
  NAND3_X1 u0_u4_u0_U93 (.A2( u0_u4_u0_n128 ) , .A1( u0_u4_u0_n132 ) , .A3( u0_u4_u0_n146 ) , .ZN( u0_u4_u0_n97 ) );
  NOR2_X1 u0_u4_u1_U10 (.A1( u0_u4_u1_n112 ) , .A2( u0_u4_u1_n116 ) , .ZN( u0_u4_u1_n118 ) );
  NAND3_X1 u0_u4_u1_U100 (.ZN( u0_u4_u1_n113 ) , .A1( u0_u4_u1_n120 ) , .A3( u0_u4_u1_n133 ) , .A2( u0_u4_u1_n155 ) );
  OAI21_X1 u0_u4_u1_U11 (.ZN( u0_u4_u1_n101 ) , .B1( u0_u4_u1_n141 ) , .A( u0_u4_u1_n146 ) , .B2( u0_u4_u1_n183 ) );
  AOI21_X1 u0_u4_u1_U12 (.B2( u0_u4_u1_n155 ) , .B1( u0_u4_u1_n156 ) , .ZN( u0_u4_u1_n157 ) , .A( u0_u4_u1_n174 ) );
  NAND2_X1 u0_u4_u1_U13 (.ZN( u0_u4_u1_n140 ) , .A2( u0_u4_u1_n150 ) , .A1( u0_u4_u1_n155 ) );
  NAND2_X1 u0_u4_u1_U14 (.A1( u0_u4_u1_n131 ) , .ZN( u0_u4_u1_n147 ) , .A2( u0_u4_u1_n153 ) );
  INV_X1 u0_u4_u1_U15 (.A( u0_u4_u1_n139 ) , .ZN( u0_u4_u1_n174 ) );
  OR4_X1 u0_u4_u1_U16 (.A4( u0_u4_u1_n106 ) , .A3( u0_u4_u1_n107 ) , .ZN( u0_u4_u1_n108 ) , .A1( u0_u4_u1_n117 ) , .A2( u0_u4_u1_n184 ) );
  AOI21_X1 u0_u4_u1_U17 (.ZN( u0_u4_u1_n106 ) , .A( u0_u4_u1_n112 ) , .B1( u0_u4_u1_n154 ) , .B2( u0_u4_u1_n156 ) );
  AOI21_X1 u0_u4_u1_U18 (.ZN( u0_u4_u1_n107 ) , .B1( u0_u4_u1_n134 ) , .B2( u0_u4_u1_n149 ) , .A( u0_u4_u1_n174 ) );
  INV_X1 u0_u4_u1_U19 (.A( u0_u4_u1_n101 ) , .ZN( u0_u4_u1_n184 ) );
  INV_X1 u0_u4_u1_U20 (.A( u0_u4_u1_n112 ) , .ZN( u0_u4_u1_n171 ) );
  NAND2_X1 u0_u4_u1_U21 (.ZN( u0_u4_u1_n141 ) , .A1( u0_u4_u1_n153 ) , .A2( u0_u4_u1_n156 ) );
  AND2_X1 u0_u4_u1_U22 (.A1( u0_u4_u1_n123 ) , .ZN( u0_u4_u1_n134 ) , .A2( u0_u4_u1_n161 ) );
  NAND2_X1 u0_u4_u1_U23 (.A2( u0_u4_u1_n115 ) , .A1( u0_u4_u1_n116 ) , .ZN( u0_u4_u1_n148 ) );
  NAND2_X1 u0_u4_u1_U24 (.A2( u0_u4_u1_n133 ) , .A1( u0_u4_u1_n135 ) , .ZN( u0_u4_u1_n159 ) );
  NAND2_X1 u0_u4_u1_U25 (.A2( u0_u4_u1_n115 ) , .A1( u0_u4_u1_n120 ) , .ZN( u0_u4_u1_n132 ) );
  INV_X1 u0_u4_u1_U26 (.A( u0_u4_u1_n154 ) , .ZN( u0_u4_u1_n178 ) );
  INV_X1 u0_u4_u1_U27 (.A( u0_u4_u1_n151 ) , .ZN( u0_u4_u1_n183 ) );
  AND2_X1 u0_u4_u1_U28 (.A1( u0_u4_u1_n129 ) , .A2( u0_u4_u1_n133 ) , .ZN( u0_u4_u1_n149 ) );
  INV_X1 u0_u4_u1_U29 (.A( u0_u4_u1_n131 ) , .ZN( u0_u4_u1_n180 ) );
  INV_X1 u0_u4_u1_U3 (.A( u0_u4_u1_n159 ) , .ZN( u0_u4_u1_n182 ) );
  OAI221_X1 u0_u4_u1_U30 (.A( u0_u4_u1_n119 ) , .C2( u0_u4_u1_n129 ) , .ZN( u0_u4_u1_n138 ) , .B2( u0_u4_u1_n152 ) , .C1( u0_u4_u1_n174 ) , .B1( u0_u4_u1_n187 ) );
  INV_X1 u0_u4_u1_U31 (.A( u0_u4_u1_n148 ) , .ZN( u0_u4_u1_n187 ) );
  AOI211_X1 u0_u4_u1_U32 (.B( u0_u4_u1_n117 ) , .A( u0_u4_u1_n118 ) , .ZN( u0_u4_u1_n119 ) , .C2( u0_u4_u1_n146 ) , .C1( u0_u4_u1_n159 ) );
  NOR2_X1 u0_u4_u1_U33 (.A1( u0_u4_u1_n168 ) , .A2( u0_u4_u1_n176 ) , .ZN( u0_u4_u1_n98 ) );
  AOI211_X1 u0_u4_u1_U34 (.B( u0_u4_u1_n162 ) , .A( u0_u4_u1_n163 ) , .C2( u0_u4_u1_n164 ) , .ZN( u0_u4_u1_n165 ) , .C1( u0_u4_u1_n171 ) );
  AOI21_X1 u0_u4_u1_U35 (.A( u0_u4_u1_n160 ) , .B2( u0_u4_u1_n161 ) , .ZN( u0_u4_u1_n162 ) , .B1( u0_u4_u1_n182 ) );
  OR2_X1 u0_u4_u1_U36 (.A2( u0_u4_u1_n157 ) , .A1( u0_u4_u1_n158 ) , .ZN( u0_u4_u1_n163 ) );
  NAND2_X1 u0_u4_u1_U37 (.A1( u0_u4_u1_n128 ) , .ZN( u0_u4_u1_n146 ) , .A2( u0_u4_u1_n160 ) );
  NAND2_X1 u0_u4_u1_U38 (.A2( u0_u4_u1_n112 ) , .ZN( u0_u4_u1_n139 ) , .A1( u0_u4_u1_n152 ) );
  NAND2_X1 u0_u4_u1_U39 (.A1( u0_u4_u1_n105 ) , .ZN( u0_u4_u1_n156 ) , .A2( u0_u4_u1_n99 ) );
  AOI221_X1 u0_u4_u1_U4 (.A( u0_u4_u1_n138 ) , .C2( u0_u4_u1_n139 ) , .C1( u0_u4_u1_n140 ) , .B2( u0_u4_u1_n141 ) , .ZN( u0_u4_u1_n142 ) , .B1( u0_u4_u1_n175 ) );
  AOI221_X1 u0_u4_u1_U40 (.B1( u0_u4_u1_n140 ) , .ZN( u0_u4_u1_n167 ) , .B2( u0_u4_u1_n172 ) , .C2( u0_u4_u1_n175 ) , .C1( u0_u4_u1_n178 ) , .A( u0_u4_u1_n188 ) );
  INV_X1 u0_u4_u1_U41 (.ZN( u0_u4_u1_n188 ) , .A( u0_u4_u1_n97 ) );
  AOI211_X1 u0_u4_u1_U42 (.A( u0_u4_u1_n118 ) , .C1( u0_u4_u1_n132 ) , .C2( u0_u4_u1_n139 ) , .B( u0_u4_u1_n96 ) , .ZN( u0_u4_u1_n97 ) );
  AOI21_X1 u0_u4_u1_U43 (.B2( u0_u4_u1_n121 ) , .B1( u0_u4_u1_n135 ) , .A( u0_u4_u1_n152 ) , .ZN( u0_u4_u1_n96 ) );
  NOR2_X1 u0_u4_u1_U44 (.ZN( u0_u4_u1_n117 ) , .A1( u0_u4_u1_n121 ) , .A2( u0_u4_u1_n160 ) );
  OAI21_X1 u0_u4_u1_U45 (.B2( u0_u4_u1_n123 ) , .ZN( u0_u4_u1_n145 ) , .B1( u0_u4_u1_n160 ) , .A( u0_u4_u1_n185 ) );
  INV_X1 u0_u4_u1_U46 (.A( u0_u4_u1_n122 ) , .ZN( u0_u4_u1_n185 ) );
  AOI21_X1 u0_u4_u1_U47 (.B2( u0_u4_u1_n120 ) , .B1( u0_u4_u1_n121 ) , .ZN( u0_u4_u1_n122 ) , .A( u0_u4_u1_n128 ) );
  AOI21_X1 u0_u4_u1_U48 (.A( u0_u4_u1_n128 ) , .B2( u0_u4_u1_n129 ) , .ZN( u0_u4_u1_n130 ) , .B1( u0_u4_u1_n150 ) );
  NAND2_X1 u0_u4_u1_U49 (.ZN( u0_u4_u1_n112 ) , .A1( u0_u4_u1_n169 ) , .A2( u0_u4_u1_n170 ) );
  AOI211_X1 u0_u4_u1_U5 (.ZN( u0_u4_u1_n124 ) , .A( u0_u4_u1_n138 ) , .C2( u0_u4_u1_n139 ) , .B( u0_u4_u1_n145 ) , .C1( u0_u4_u1_n147 ) );
  NAND2_X1 u0_u4_u1_U50 (.ZN( u0_u4_u1_n129 ) , .A2( u0_u4_u1_n95 ) , .A1( u0_u4_u1_n98 ) );
  NAND2_X1 u0_u4_u1_U51 (.A1( u0_u4_u1_n102 ) , .ZN( u0_u4_u1_n154 ) , .A2( u0_u4_u1_n99 ) );
  NAND2_X1 u0_u4_u1_U52 (.A2( u0_u4_u1_n100 ) , .ZN( u0_u4_u1_n135 ) , .A1( u0_u4_u1_n99 ) );
  AOI21_X1 u0_u4_u1_U53 (.A( u0_u4_u1_n152 ) , .B2( u0_u4_u1_n153 ) , .B1( u0_u4_u1_n154 ) , .ZN( u0_u4_u1_n158 ) );
  INV_X1 u0_u4_u1_U54 (.A( u0_u4_u1_n160 ) , .ZN( u0_u4_u1_n175 ) );
  NAND2_X1 u0_u4_u1_U55 (.A1( u0_u4_u1_n100 ) , .ZN( u0_u4_u1_n116 ) , .A2( u0_u4_u1_n95 ) );
  NAND2_X1 u0_u4_u1_U56 (.A1( u0_u4_u1_n102 ) , .ZN( u0_u4_u1_n131 ) , .A2( u0_u4_u1_n95 ) );
  NAND2_X1 u0_u4_u1_U57 (.A2( u0_u4_u1_n104 ) , .ZN( u0_u4_u1_n121 ) , .A1( u0_u4_u1_n98 ) );
  NAND2_X1 u0_u4_u1_U58 (.A1( u0_u4_u1_n103 ) , .ZN( u0_u4_u1_n153 ) , .A2( u0_u4_u1_n98 ) );
  NAND2_X1 u0_u4_u1_U59 (.A2( u0_u4_u1_n104 ) , .A1( u0_u4_u1_n105 ) , .ZN( u0_u4_u1_n133 ) );
  AOI22_X1 u0_u4_u1_U6 (.B2( u0_u4_u1_n113 ) , .A2( u0_u4_u1_n114 ) , .ZN( u0_u4_u1_n125 ) , .A1( u0_u4_u1_n171 ) , .B1( u0_u4_u1_n173 ) );
  NAND2_X1 u0_u4_u1_U60 (.ZN( u0_u4_u1_n150 ) , .A2( u0_u4_u1_n98 ) , .A1( u0_u4_u1_n99 ) );
  NAND2_X1 u0_u4_u1_U61 (.A1( u0_u4_u1_n105 ) , .ZN( u0_u4_u1_n155 ) , .A2( u0_u4_u1_n95 ) );
  OAI21_X1 u0_u4_u1_U62 (.ZN( u0_u4_u1_n109 ) , .B1( u0_u4_u1_n129 ) , .B2( u0_u4_u1_n160 ) , .A( u0_u4_u1_n167 ) );
  NAND2_X1 u0_u4_u1_U63 (.A2( u0_u4_u1_n100 ) , .A1( u0_u4_u1_n103 ) , .ZN( u0_u4_u1_n120 ) );
  NAND2_X1 u0_u4_u1_U64 (.A1( u0_u4_u1_n102 ) , .A2( u0_u4_u1_n104 ) , .ZN( u0_u4_u1_n115 ) );
  NAND2_X1 u0_u4_u1_U65 (.A2( u0_u4_u1_n100 ) , .A1( u0_u4_u1_n104 ) , .ZN( u0_u4_u1_n151 ) );
  NAND2_X1 u0_u4_u1_U66 (.A2( u0_u4_u1_n103 ) , .A1( u0_u4_u1_n105 ) , .ZN( u0_u4_u1_n161 ) );
  INV_X1 u0_u4_u1_U67 (.A( u0_u4_u1_n152 ) , .ZN( u0_u4_u1_n173 ) );
  INV_X1 u0_u4_u1_U68 (.A( u0_u4_u1_n128 ) , .ZN( u0_u4_u1_n172 ) );
  NAND2_X1 u0_u4_u1_U69 (.A2( u0_u4_u1_n102 ) , .A1( u0_u4_u1_n103 ) , .ZN( u0_u4_u1_n123 ) );
  NAND2_X1 u0_u4_u1_U7 (.ZN( u0_u4_u1_n114 ) , .A1( u0_u4_u1_n134 ) , .A2( u0_u4_u1_n156 ) );
  NOR2_X1 u0_u4_u1_U70 (.A2( u0_u4_X_7 ) , .A1( u0_u4_X_8 ) , .ZN( u0_u4_u1_n95 ) );
  NOR2_X1 u0_u4_u1_U71 (.A1( u0_u4_X_12 ) , .A2( u0_u4_X_9 ) , .ZN( u0_u4_u1_n100 ) );
  NOR2_X1 u0_u4_u1_U72 (.A2( u0_u4_X_8 ) , .A1( u0_u4_u1_n177 ) , .ZN( u0_u4_u1_n99 ) );
  NOR2_X1 u0_u4_u1_U73 (.A2( u0_u4_X_12 ) , .ZN( u0_u4_u1_n102 ) , .A1( u0_u4_u1_n176 ) );
  NOR2_X1 u0_u4_u1_U74 (.A2( u0_u4_X_9 ) , .ZN( u0_u4_u1_n105 ) , .A1( u0_u4_u1_n168 ) );
  NAND2_X1 u0_u4_u1_U75 (.A1( u0_u4_X_10 ) , .ZN( u0_u4_u1_n160 ) , .A2( u0_u4_u1_n169 ) );
  NAND2_X1 u0_u4_u1_U76 (.A2( u0_u4_X_10 ) , .A1( u0_u4_X_11 ) , .ZN( u0_u4_u1_n152 ) );
  NAND2_X1 u0_u4_u1_U77 (.A1( u0_u4_X_11 ) , .ZN( u0_u4_u1_n128 ) , .A2( u0_u4_u1_n170 ) );
  AND2_X1 u0_u4_u1_U78 (.A2( u0_u4_X_7 ) , .A1( u0_u4_X_8 ) , .ZN( u0_u4_u1_n104 ) );
  AND2_X1 u0_u4_u1_U79 (.A1( u0_u4_X_8 ) , .ZN( u0_u4_u1_n103 ) , .A2( u0_u4_u1_n177 ) );
  AOI22_X1 u0_u4_u1_U8 (.B2( u0_u4_u1_n136 ) , .A2( u0_u4_u1_n137 ) , .ZN( u0_u4_u1_n143 ) , .A1( u0_u4_u1_n171 ) , .B1( u0_u4_u1_n173 ) );
  INV_X1 u0_u4_u1_U80 (.A( u0_u4_X_10 ) , .ZN( u0_u4_u1_n170 ) );
  INV_X1 u0_u4_u1_U81 (.A( u0_u4_X_9 ) , .ZN( u0_u4_u1_n176 ) );
  INV_X1 u0_u4_u1_U82 (.A( u0_u4_X_11 ) , .ZN( u0_u4_u1_n169 ) );
  INV_X1 u0_u4_u1_U83 (.A( u0_u4_X_12 ) , .ZN( u0_u4_u1_n168 ) );
  INV_X1 u0_u4_u1_U84 (.A( u0_u4_X_7 ) , .ZN( u0_u4_u1_n177 ) );
  NAND4_X1 u0_u4_u1_U85 (.ZN( u0_out4_28 ) , .A4( u0_u4_u1_n124 ) , .A3( u0_u4_u1_n125 ) , .A2( u0_u4_u1_n126 ) , .A1( u0_u4_u1_n127 ) );
  OAI21_X1 u0_u4_u1_U86 (.ZN( u0_u4_u1_n127 ) , .B2( u0_u4_u1_n139 ) , .B1( u0_u4_u1_n175 ) , .A( u0_u4_u1_n183 ) );
  OAI21_X1 u0_u4_u1_U87 (.ZN( u0_u4_u1_n126 ) , .B2( u0_u4_u1_n140 ) , .A( u0_u4_u1_n146 ) , .B1( u0_u4_u1_n178 ) );
  NAND4_X1 u0_u4_u1_U88 (.ZN( u0_out4_18 ) , .A4( u0_u4_u1_n165 ) , .A3( u0_u4_u1_n166 ) , .A1( u0_u4_u1_n167 ) , .A2( u0_u4_u1_n186 ) );
  AOI22_X1 u0_u4_u1_U89 (.B2( u0_u4_u1_n146 ) , .B1( u0_u4_u1_n147 ) , .A2( u0_u4_u1_n148 ) , .ZN( u0_u4_u1_n166 ) , .A1( u0_u4_u1_n172 ) );
  INV_X1 u0_u4_u1_U9 (.A( u0_u4_u1_n147 ) , .ZN( u0_u4_u1_n181 ) );
  INV_X1 u0_u4_u1_U90 (.A( u0_u4_u1_n145 ) , .ZN( u0_u4_u1_n186 ) );
  NAND4_X1 u0_u4_u1_U91 (.ZN( u0_out4_2 ) , .A4( u0_u4_u1_n142 ) , .A3( u0_u4_u1_n143 ) , .A2( u0_u4_u1_n144 ) , .A1( u0_u4_u1_n179 ) );
  OAI21_X1 u0_u4_u1_U92 (.B2( u0_u4_u1_n132 ) , .ZN( u0_u4_u1_n144 ) , .A( u0_u4_u1_n146 ) , .B1( u0_u4_u1_n180 ) );
  INV_X1 u0_u4_u1_U93 (.A( u0_u4_u1_n130 ) , .ZN( u0_u4_u1_n179 ) );
  OR4_X1 u0_u4_u1_U94 (.ZN( u0_out4_13 ) , .A4( u0_u4_u1_n108 ) , .A3( u0_u4_u1_n109 ) , .A2( u0_u4_u1_n110 ) , .A1( u0_u4_u1_n111 ) );
  AOI21_X1 u0_u4_u1_U95 (.ZN( u0_u4_u1_n111 ) , .A( u0_u4_u1_n128 ) , .B2( u0_u4_u1_n131 ) , .B1( u0_u4_u1_n135 ) );
  AOI21_X1 u0_u4_u1_U96 (.ZN( u0_u4_u1_n110 ) , .A( u0_u4_u1_n116 ) , .B1( u0_u4_u1_n152 ) , .B2( u0_u4_u1_n160 ) );
  NAND3_X1 u0_u4_u1_U97 (.A3( u0_u4_u1_n149 ) , .A2( u0_u4_u1_n150 ) , .A1( u0_u4_u1_n151 ) , .ZN( u0_u4_u1_n164 ) );
  NAND3_X1 u0_u4_u1_U98 (.A3( u0_u4_u1_n134 ) , .A2( u0_u4_u1_n135 ) , .ZN( u0_u4_u1_n136 ) , .A1( u0_u4_u1_n151 ) );
  NAND3_X1 u0_u4_u1_U99 (.A1( u0_u4_u1_n133 ) , .ZN( u0_u4_u1_n137 ) , .A2( u0_u4_u1_n154 ) , .A3( u0_u4_u1_n181 ) );
  OAI22_X1 u0_u4_u2_U10 (.ZN( u0_u4_u2_n109 ) , .A2( u0_u4_u2_n113 ) , .B2( u0_u4_u2_n133 ) , .B1( u0_u4_u2_n167 ) , .A1( u0_u4_u2_n168 ) );
  NAND3_X1 u0_u4_u2_U100 (.A2( u0_u4_u2_n100 ) , .A1( u0_u4_u2_n104 ) , .A3( u0_u4_u2_n138 ) , .ZN( u0_u4_u2_n98 ) );
  OAI22_X1 u0_u4_u2_U11 (.B1( u0_u4_u2_n151 ) , .A2( u0_u4_u2_n152 ) , .A1( u0_u4_u2_n153 ) , .ZN( u0_u4_u2_n160 ) , .B2( u0_u4_u2_n168 ) );
  NOR3_X1 u0_u4_u2_U12 (.A1( u0_u4_u2_n150 ) , .ZN( u0_u4_u2_n151 ) , .A3( u0_u4_u2_n175 ) , .A2( u0_u4_u2_n188 ) );
  AOI21_X1 u0_u4_u2_U13 (.ZN( u0_u4_u2_n144 ) , .B2( u0_u4_u2_n155 ) , .A( u0_u4_u2_n172 ) , .B1( u0_u4_u2_n185 ) );
  AOI21_X1 u0_u4_u2_U14 (.B2( u0_u4_u2_n143 ) , .ZN( u0_u4_u2_n145 ) , .B1( u0_u4_u2_n152 ) , .A( u0_u4_u2_n171 ) );
  AOI21_X1 u0_u4_u2_U15 (.B2( u0_u4_u2_n120 ) , .B1( u0_u4_u2_n121 ) , .ZN( u0_u4_u2_n126 ) , .A( u0_u4_u2_n167 ) );
  INV_X1 u0_u4_u2_U16 (.A( u0_u4_u2_n156 ) , .ZN( u0_u4_u2_n171 ) );
  INV_X1 u0_u4_u2_U17 (.A( u0_u4_u2_n120 ) , .ZN( u0_u4_u2_n188 ) );
  NAND2_X1 u0_u4_u2_U18 (.A2( u0_u4_u2_n122 ) , .ZN( u0_u4_u2_n150 ) , .A1( u0_u4_u2_n152 ) );
  INV_X1 u0_u4_u2_U19 (.A( u0_u4_u2_n153 ) , .ZN( u0_u4_u2_n170 ) );
  INV_X1 u0_u4_u2_U20 (.A( u0_u4_u2_n137 ) , .ZN( u0_u4_u2_n173 ) );
  NAND2_X1 u0_u4_u2_U21 (.A1( u0_u4_u2_n132 ) , .A2( u0_u4_u2_n139 ) , .ZN( u0_u4_u2_n157 ) );
  INV_X1 u0_u4_u2_U22 (.A( u0_u4_u2_n113 ) , .ZN( u0_u4_u2_n178 ) );
  INV_X1 u0_u4_u2_U23 (.A( u0_u4_u2_n139 ) , .ZN( u0_u4_u2_n175 ) );
  INV_X1 u0_u4_u2_U24 (.A( u0_u4_u2_n155 ) , .ZN( u0_u4_u2_n181 ) );
  INV_X1 u0_u4_u2_U25 (.A( u0_u4_u2_n119 ) , .ZN( u0_u4_u2_n177 ) );
  INV_X1 u0_u4_u2_U26 (.A( u0_u4_u2_n116 ) , .ZN( u0_u4_u2_n180 ) );
  INV_X1 u0_u4_u2_U27 (.A( u0_u4_u2_n131 ) , .ZN( u0_u4_u2_n179 ) );
  INV_X1 u0_u4_u2_U28 (.A( u0_u4_u2_n154 ) , .ZN( u0_u4_u2_n176 ) );
  NAND2_X1 u0_u4_u2_U29 (.A2( u0_u4_u2_n116 ) , .A1( u0_u4_u2_n117 ) , .ZN( u0_u4_u2_n118 ) );
  NOR2_X1 u0_u4_u2_U3 (.ZN( u0_u4_u2_n121 ) , .A2( u0_u4_u2_n177 ) , .A1( u0_u4_u2_n180 ) );
  INV_X1 u0_u4_u2_U30 (.A( u0_u4_u2_n132 ) , .ZN( u0_u4_u2_n182 ) );
  INV_X1 u0_u4_u2_U31 (.A( u0_u4_u2_n158 ) , .ZN( u0_u4_u2_n183 ) );
  OAI21_X1 u0_u4_u2_U32 (.A( u0_u4_u2_n156 ) , .B1( u0_u4_u2_n157 ) , .ZN( u0_u4_u2_n158 ) , .B2( u0_u4_u2_n179 ) );
  NOR2_X1 u0_u4_u2_U33 (.ZN( u0_u4_u2_n156 ) , .A1( u0_u4_u2_n166 ) , .A2( u0_u4_u2_n169 ) );
  NOR2_X1 u0_u4_u2_U34 (.A2( u0_u4_u2_n114 ) , .ZN( u0_u4_u2_n137 ) , .A1( u0_u4_u2_n140 ) );
  NOR2_X1 u0_u4_u2_U35 (.A2( u0_u4_u2_n138 ) , .ZN( u0_u4_u2_n153 ) , .A1( u0_u4_u2_n156 ) );
  AOI211_X1 u0_u4_u2_U36 (.ZN( u0_u4_u2_n130 ) , .C1( u0_u4_u2_n138 ) , .C2( u0_u4_u2_n179 ) , .B( u0_u4_u2_n96 ) , .A( u0_u4_u2_n97 ) );
  OAI22_X1 u0_u4_u2_U37 (.B1( u0_u4_u2_n133 ) , .A2( u0_u4_u2_n137 ) , .A1( u0_u4_u2_n152 ) , .B2( u0_u4_u2_n168 ) , .ZN( u0_u4_u2_n97 ) );
  OAI221_X1 u0_u4_u2_U38 (.B1( u0_u4_u2_n113 ) , .C1( u0_u4_u2_n132 ) , .A( u0_u4_u2_n149 ) , .B2( u0_u4_u2_n171 ) , .C2( u0_u4_u2_n172 ) , .ZN( u0_u4_u2_n96 ) );
  OAI221_X1 u0_u4_u2_U39 (.A( u0_u4_u2_n115 ) , .C2( u0_u4_u2_n123 ) , .B2( u0_u4_u2_n143 ) , .B1( u0_u4_u2_n153 ) , .ZN( u0_u4_u2_n163 ) , .C1( u0_u4_u2_n168 ) );
  INV_X1 u0_u4_u2_U4 (.A( u0_u4_u2_n134 ) , .ZN( u0_u4_u2_n185 ) );
  OAI21_X1 u0_u4_u2_U40 (.A( u0_u4_u2_n114 ) , .ZN( u0_u4_u2_n115 ) , .B1( u0_u4_u2_n176 ) , .B2( u0_u4_u2_n178 ) );
  OAI221_X1 u0_u4_u2_U41 (.A( u0_u4_u2_n135 ) , .B2( u0_u4_u2_n136 ) , .B1( u0_u4_u2_n137 ) , .ZN( u0_u4_u2_n162 ) , .C2( u0_u4_u2_n167 ) , .C1( u0_u4_u2_n185 ) );
  AND3_X1 u0_u4_u2_U42 (.A3( u0_u4_u2_n131 ) , .A2( u0_u4_u2_n132 ) , .A1( u0_u4_u2_n133 ) , .ZN( u0_u4_u2_n136 ) );
  AOI22_X1 u0_u4_u2_U43 (.ZN( u0_u4_u2_n135 ) , .B1( u0_u4_u2_n140 ) , .A1( u0_u4_u2_n156 ) , .B2( u0_u4_u2_n180 ) , .A2( u0_u4_u2_n188 ) );
  AOI21_X1 u0_u4_u2_U44 (.ZN( u0_u4_u2_n149 ) , .B1( u0_u4_u2_n173 ) , .B2( u0_u4_u2_n188 ) , .A( u0_u4_u2_n95 ) );
  AND3_X1 u0_u4_u2_U45 (.A2( u0_u4_u2_n100 ) , .A1( u0_u4_u2_n104 ) , .A3( u0_u4_u2_n156 ) , .ZN( u0_u4_u2_n95 ) );
  OAI21_X1 u0_u4_u2_U46 (.A( u0_u4_u2_n101 ) , .B2( u0_u4_u2_n121 ) , .B1( u0_u4_u2_n153 ) , .ZN( u0_u4_u2_n164 ) );
  NAND2_X1 u0_u4_u2_U47 (.A2( u0_u4_u2_n100 ) , .A1( u0_u4_u2_n107 ) , .ZN( u0_u4_u2_n155 ) );
  NAND2_X1 u0_u4_u2_U48 (.A2( u0_u4_u2_n105 ) , .A1( u0_u4_u2_n108 ) , .ZN( u0_u4_u2_n143 ) );
  NAND2_X1 u0_u4_u2_U49 (.A1( u0_u4_u2_n104 ) , .A2( u0_u4_u2_n106 ) , .ZN( u0_u4_u2_n152 ) );
  INV_X1 u0_u4_u2_U5 (.A( u0_u4_u2_n150 ) , .ZN( u0_u4_u2_n184 ) );
  NAND2_X1 u0_u4_u2_U50 (.A1( u0_u4_u2_n100 ) , .A2( u0_u4_u2_n105 ) , .ZN( u0_u4_u2_n132 ) );
  INV_X1 u0_u4_u2_U51 (.A( u0_u4_u2_n140 ) , .ZN( u0_u4_u2_n168 ) );
  INV_X1 u0_u4_u2_U52 (.A( u0_u4_u2_n138 ) , .ZN( u0_u4_u2_n167 ) );
  OAI21_X1 u0_u4_u2_U53 (.A( u0_u4_u2_n141 ) , .B2( u0_u4_u2_n142 ) , .ZN( u0_u4_u2_n146 ) , .B1( u0_u4_u2_n153 ) );
  OAI21_X1 u0_u4_u2_U54 (.A( u0_u4_u2_n140 ) , .ZN( u0_u4_u2_n141 ) , .B1( u0_u4_u2_n176 ) , .B2( u0_u4_u2_n177 ) );
  NOR3_X1 u0_u4_u2_U55 (.ZN( u0_u4_u2_n142 ) , .A3( u0_u4_u2_n175 ) , .A2( u0_u4_u2_n178 ) , .A1( u0_u4_u2_n181 ) );
  INV_X1 u0_u4_u2_U56 (.ZN( u0_u4_u2_n187 ) , .A( u0_u4_u2_n99 ) );
  OAI21_X1 u0_u4_u2_U57 (.B1( u0_u4_u2_n137 ) , .B2( u0_u4_u2_n143 ) , .A( u0_u4_u2_n98 ) , .ZN( u0_u4_u2_n99 ) );
  NAND2_X1 u0_u4_u2_U58 (.A1( u0_u4_u2_n102 ) , .A2( u0_u4_u2_n106 ) , .ZN( u0_u4_u2_n113 ) );
  NAND2_X1 u0_u4_u2_U59 (.A1( u0_u4_u2_n106 ) , .A2( u0_u4_u2_n107 ) , .ZN( u0_u4_u2_n131 ) );
  NOR4_X1 u0_u4_u2_U6 (.A4( u0_u4_u2_n124 ) , .A3( u0_u4_u2_n125 ) , .A2( u0_u4_u2_n126 ) , .A1( u0_u4_u2_n127 ) , .ZN( u0_u4_u2_n128 ) );
  NAND2_X1 u0_u4_u2_U60 (.A1( u0_u4_u2_n103 ) , .A2( u0_u4_u2_n107 ) , .ZN( u0_u4_u2_n139 ) );
  NAND2_X1 u0_u4_u2_U61 (.A1( u0_u4_u2_n103 ) , .A2( u0_u4_u2_n105 ) , .ZN( u0_u4_u2_n133 ) );
  NAND2_X1 u0_u4_u2_U62 (.A1( u0_u4_u2_n102 ) , .A2( u0_u4_u2_n103 ) , .ZN( u0_u4_u2_n154 ) );
  NAND2_X1 u0_u4_u2_U63 (.A2( u0_u4_u2_n103 ) , .A1( u0_u4_u2_n104 ) , .ZN( u0_u4_u2_n119 ) );
  NAND2_X1 u0_u4_u2_U64 (.A2( u0_u4_u2_n107 ) , .A1( u0_u4_u2_n108 ) , .ZN( u0_u4_u2_n123 ) );
  NAND2_X1 u0_u4_u2_U65 (.A1( u0_u4_u2_n104 ) , .A2( u0_u4_u2_n108 ) , .ZN( u0_u4_u2_n122 ) );
  INV_X1 u0_u4_u2_U66 (.A( u0_u4_u2_n114 ) , .ZN( u0_u4_u2_n172 ) );
  NAND2_X1 u0_u4_u2_U67 (.A2( u0_u4_u2_n100 ) , .A1( u0_u4_u2_n102 ) , .ZN( u0_u4_u2_n116 ) );
  NAND2_X1 u0_u4_u2_U68 (.A1( u0_u4_u2_n102 ) , .A2( u0_u4_u2_n108 ) , .ZN( u0_u4_u2_n120 ) );
  NAND2_X1 u0_u4_u2_U69 (.A2( u0_u4_u2_n105 ) , .A1( u0_u4_u2_n106 ) , .ZN( u0_u4_u2_n117 ) );
  AOI21_X1 u0_u4_u2_U7 (.B2( u0_u4_u2_n119 ) , .ZN( u0_u4_u2_n127 ) , .A( u0_u4_u2_n137 ) , .B1( u0_u4_u2_n155 ) );
  NOR2_X1 u0_u4_u2_U70 (.A2( u0_u4_X_16 ) , .ZN( u0_u4_u2_n140 ) , .A1( u0_u4_u2_n166 ) );
  NOR2_X1 u0_u4_u2_U71 (.A2( u0_u4_X_13 ) , .A1( u0_u4_X_14 ) , .ZN( u0_u4_u2_n100 ) );
  NOR2_X1 u0_u4_u2_U72 (.A2( u0_u4_X_16 ) , .A1( u0_u4_X_17 ) , .ZN( u0_u4_u2_n138 ) );
  NOR2_X1 u0_u4_u2_U73 (.A2( u0_u4_X_15 ) , .A1( u0_u4_X_18 ) , .ZN( u0_u4_u2_n104 ) );
  NOR2_X1 u0_u4_u2_U74 (.A2( u0_u4_X_14 ) , .ZN( u0_u4_u2_n103 ) , .A1( u0_u4_u2_n174 ) );
  NOR2_X1 u0_u4_u2_U75 (.A2( u0_u4_X_15 ) , .ZN( u0_u4_u2_n102 ) , .A1( u0_u4_u2_n165 ) );
  NOR2_X1 u0_u4_u2_U76 (.A2( u0_u4_X_17 ) , .ZN( u0_u4_u2_n114 ) , .A1( u0_u4_u2_n169 ) );
  AND2_X1 u0_u4_u2_U77 (.A1( u0_u4_X_15 ) , .ZN( u0_u4_u2_n105 ) , .A2( u0_u4_u2_n165 ) );
  AND2_X1 u0_u4_u2_U78 (.A2( u0_u4_X_15 ) , .A1( u0_u4_X_18 ) , .ZN( u0_u4_u2_n107 ) );
  AND2_X1 u0_u4_u2_U79 (.A1( u0_u4_X_14 ) , .ZN( u0_u4_u2_n106 ) , .A2( u0_u4_u2_n174 ) );
  AOI21_X1 u0_u4_u2_U8 (.ZN( u0_u4_u2_n124 ) , .B1( u0_u4_u2_n131 ) , .B2( u0_u4_u2_n143 ) , .A( u0_u4_u2_n172 ) );
  AND2_X1 u0_u4_u2_U80 (.A1( u0_u4_X_13 ) , .A2( u0_u4_X_14 ) , .ZN( u0_u4_u2_n108 ) );
  INV_X1 u0_u4_u2_U81 (.A( u0_u4_X_16 ) , .ZN( u0_u4_u2_n169 ) );
  INV_X1 u0_u4_u2_U82 (.A( u0_u4_X_17 ) , .ZN( u0_u4_u2_n166 ) );
  INV_X1 u0_u4_u2_U83 (.A( u0_u4_X_13 ) , .ZN( u0_u4_u2_n174 ) );
  INV_X1 u0_u4_u2_U84 (.A( u0_u4_X_18 ) , .ZN( u0_u4_u2_n165 ) );
  NAND4_X1 u0_u4_u2_U85 (.ZN( u0_out4_30 ) , .A4( u0_u4_u2_n147 ) , .A3( u0_u4_u2_n148 ) , .A2( u0_u4_u2_n149 ) , .A1( u0_u4_u2_n187 ) );
  NOR3_X1 u0_u4_u2_U86 (.A3( u0_u4_u2_n144 ) , .A2( u0_u4_u2_n145 ) , .A1( u0_u4_u2_n146 ) , .ZN( u0_u4_u2_n147 ) );
  AOI21_X1 u0_u4_u2_U87 (.B2( u0_u4_u2_n138 ) , .ZN( u0_u4_u2_n148 ) , .A( u0_u4_u2_n162 ) , .B1( u0_u4_u2_n182 ) );
  NAND4_X1 u0_u4_u2_U88 (.ZN( u0_out4_24 ) , .A4( u0_u4_u2_n111 ) , .A3( u0_u4_u2_n112 ) , .A1( u0_u4_u2_n130 ) , .A2( u0_u4_u2_n187 ) );
  AOI221_X1 u0_u4_u2_U89 (.A( u0_u4_u2_n109 ) , .B1( u0_u4_u2_n110 ) , .ZN( u0_u4_u2_n111 ) , .C1( u0_u4_u2_n134 ) , .C2( u0_u4_u2_n170 ) , .B2( u0_u4_u2_n173 ) );
  AOI21_X1 u0_u4_u2_U9 (.B2( u0_u4_u2_n123 ) , .ZN( u0_u4_u2_n125 ) , .A( u0_u4_u2_n171 ) , .B1( u0_u4_u2_n184 ) );
  AOI21_X1 u0_u4_u2_U90 (.ZN( u0_u4_u2_n112 ) , .B2( u0_u4_u2_n156 ) , .A( u0_u4_u2_n164 ) , .B1( u0_u4_u2_n181 ) );
  NAND4_X1 u0_u4_u2_U91 (.ZN( u0_out4_16 ) , .A4( u0_u4_u2_n128 ) , .A3( u0_u4_u2_n129 ) , .A1( u0_u4_u2_n130 ) , .A2( u0_u4_u2_n186 ) );
  AOI22_X1 u0_u4_u2_U92 (.A2( u0_u4_u2_n118 ) , .ZN( u0_u4_u2_n129 ) , .A1( u0_u4_u2_n140 ) , .B1( u0_u4_u2_n157 ) , .B2( u0_u4_u2_n170 ) );
  INV_X1 u0_u4_u2_U93 (.A( u0_u4_u2_n163 ) , .ZN( u0_u4_u2_n186 ) );
  OR4_X1 u0_u4_u2_U94 (.ZN( u0_out4_6 ) , .A4( u0_u4_u2_n161 ) , .A3( u0_u4_u2_n162 ) , .A2( u0_u4_u2_n163 ) , .A1( u0_u4_u2_n164 ) );
  OR3_X1 u0_u4_u2_U95 (.A2( u0_u4_u2_n159 ) , .A1( u0_u4_u2_n160 ) , .ZN( u0_u4_u2_n161 ) , .A3( u0_u4_u2_n183 ) );
  AOI21_X1 u0_u4_u2_U96 (.B2( u0_u4_u2_n154 ) , .B1( u0_u4_u2_n155 ) , .ZN( u0_u4_u2_n159 ) , .A( u0_u4_u2_n167 ) );
  NAND3_X1 u0_u4_u2_U97 (.A2( u0_u4_u2_n117 ) , .A1( u0_u4_u2_n122 ) , .A3( u0_u4_u2_n123 ) , .ZN( u0_u4_u2_n134 ) );
  NAND3_X1 u0_u4_u2_U98 (.ZN( u0_u4_u2_n110 ) , .A2( u0_u4_u2_n131 ) , .A3( u0_u4_u2_n139 ) , .A1( u0_u4_u2_n154 ) );
  NAND3_X1 u0_u4_u2_U99 (.A2( u0_u4_u2_n100 ) , .ZN( u0_u4_u2_n101 ) , .A1( u0_u4_u2_n104 ) , .A3( u0_u4_u2_n114 ) );
  OAI22_X1 u0_u4_u3_U10 (.B1( u0_u4_u3_n113 ) , .A2( u0_u4_u3_n135 ) , .A1( u0_u4_u3_n150 ) , .B2( u0_u4_u3_n164 ) , .ZN( u0_u4_u3_n98 ) );
  OAI211_X1 u0_u4_u3_U11 (.B( u0_u4_u3_n106 ) , .ZN( u0_u4_u3_n119 ) , .C2( u0_u4_u3_n128 ) , .C1( u0_u4_u3_n167 ) , .A( u0_u4_u3_n181 ) );
  AOI221_X1 u0_u4_u3_U12 (.C1( u0_u4_u3_n105 ) , .ZN( u0_u4_u3_n106 ) , .A( u0_u4_u3_n131 ) , .B2( u0_u4_u3_n132 ) , .C2( u0_u4_u3_n133 ) , .B1( u0_u4_u3_n169 ) );
  INV_X1 u0_u4_u3_U13 (.ZN( u0_u4_u3_n181 ) , .A( u0_u4_u3_n98 ) );
  NAND2_X1 u0_u4_u3_U14 (.ZN( u0_u4_u3_n105 ) , .A2( u0_u4_u3_n130 ) , .A1( u0_u4_u3_n155 ) );
  AOI22_X1 u0_u4_u3_U15 (.B1( u0_u4_u3_n115 ) , .A2( u0_u4_u3_n116 ) , .ZN( u0_u4_u3_n123 ) , .B2( u0_u4_u3_n133 ) , .A1( u0_u4_u3_n169 ) );
  NAND2_X1 u0_u4_u3_U16 (.ZN( u0_u4_u3_n116 ) , .A2( u0_u4_u3_n151 ) , .A1( u0_u4_u3_n182 ) );
  NOR2_X1 u0_u4_u3_U17 (.ZN( u0_u4_u3_n126 ) , .A2( u0_u4_u3_n150 ) , .A1( u0_u4_u3_n164 ) );
  AOI21_X1 u0_u4_u3_U18 (.ZN( u0_u4_u3_n112 ) , .B2( u0_u4_u3_n146 ) , .B1( u0_u4_u3_n155 ) , .A( u0_u4_u3_n167 ) );
  NAND2_X1 u0_u4_u3_U19 (.A1( u0_u4_u3_n135 ) , .ZN( u0_u4_u3_n142 ) , .A2( u0_u4_u3_n164 ) );
  NAND2_X1 u0_u4_u3_U20 (.ZN( u0_u4_u3_n132 ) , .A2( u0_u4_u3_n152 ) , .A1( u0_u4_u3_n156 ) );
  AND2_X1 u0_u4_u3_U21 (.A2( u0_u4_u3_n113 ) , .A1( u0_u4_u3_n114 ) , .ZN( u0_u4_u3_n151 ) );
  INV_X1 u0_u4_u3_U22 (.A( u0_u4_u3_n133 ) , .ZN( u0_u4_u3_n165 ) );
  INV_X1 u0_u4_u3_U23 (.A( u0_u4_u3_n135 ) , .ZN( u0_u4_u3_n170 ) );
  NAND2_X1 u0_u4_u3_U24 (.A1( u0_u4_u3_n107 ) , .A2( u0_u4_u3_n108 ) , .ZN( u0_u4_u3_n140 ) );
  NAND2_X1 u0_u4_u3_U25 (.ZN( u0_u4_u3_n117 ) , .A1( u0_u4_u3_n124 ) , .A2( u0_u4_u3_n148 ) );
  NAND2_X1 u0_u4_u3_U26 (.ZN( u0_u4_u3_n143 ) , .A1( u0_u4_u3_n165 ) , .A2( u0_u4_u3_n167 ) );
  INV_X1 u0_u4_u3_U27 (.A( u0_u4_u3_n130 ) , .ZN( u0_u4_u3_n177 ) );
  INV_X1 u0_u4_u3_U28 (.A( u0_u4_u3_n128 ) , .ZN( u0_u4_u3_n176 ) );
  INV_X1 u0_u4_u3_U29 (.A( u0_u4_u3_n155 ) , .ZN( u0_u4_u3_n174 ) );
  INV_X1 u0_u4_u3_U3 (.A( u0_u4_u3_n129 ) , .ZN( u0_u4_u3_n183 ) );
  INV_X1 u0_u4_u3_U30 (.A( u0_u4_u3_n139 ) , .ZN( u0_u4_u3_n185 ) );
  NOR2_X1 u0_u4_u3_U31 (.ZN( u0_u4_u3_n135 ) , .A2( u0_u4_u3_n141 ) , .A1( u0_u4_u3_n169 ) );
  OAI222_X1 u0_u4_u3_U32 (.C2( u0_u4_u3_n107 ) , .A2( u0_u4_u3_n108 ) , .B1( u0_u4_u3_n135 ) , .ZN( u0_u4_u3_n138 ) , .B2( u0_u4_u3_n146 ) , .C1( u0_u4_u3_n154 ) , .A1( u0_u4_u3_n164 ) );
  NOR4_X1 u0_u4_u3_U33 (.A4( u0_u4_u3_n157 ) , .A3( u0_u4_u3_n158 ) , .A2( u0_u4_u3_n159 ) , .A1( u0_u4_u3_n160 ) , .ZN( u0_u4_u3_n161 ) );
  AOI21_X1 u0_u4_u3_U34 (.B2( u0_u4_u3_n152 ) , .B1( u0_u4_u3_n153 ) , .ZN( u0_u4_u3_n158 ) , .A( u0_u4_u3_n164 ) );
  AOI21_X1 u0_u4_u3_U35 (.A( u0_u4_u3_n149 ) , .B2( u0_u4_u3_n150 ) , .B1( u0_u4_u3_n151 ) , .ZN( u0_u4_u3_n159 ) );
  AOI21_X1 u0_u4_u3_U36 (.A( u0_u4_u3_n154 ) , .B2( u0_u4_u3_n155 ) , .B1( u0_u4_u3_n156 ) , .ZN( u0_u4_u3_n157 ) );
  AOI211_X1 u0_u4_u3_U37 (.ZN( u0_u4_u3_n109 ) , .A( u0_u4_u3_n119 ) , .C2( u0_u4_u3_n129 ) , .B( u0_u4_u3_n138 ) , .C1( u0_u4_u3_n141 ) );
  AOI211_X1 u0_u4_u3_U38 (.B( u0_u4_u3_n119 ) , .A( u0_u4_u3_n120 ) , .C2( u0_u4_u3_n121 ) , .ZN( u0_u4_u3_n122 ) , .C1( u0_u4_u3_n179 ) );
  INV_X1 u0_u4_u3_U39 (.A( u0_u4_u3_n156 ) , .ZN( u0_u4_u3_n179 ) );
  INV_X1 u0_u4_u3_U4 (.A( u0_u4_u3_n140 ) , .ZN( u0_u4_u3_n182 ) );
  OAI22_X1 u0_u4_u3_U40 (.B1( u0_u4_u3_n118 ) , .ZN( u0_u4_u3_n120 ) , .A1( u0_u4_u3_n135 ) , .B2( u0_u4_u3_n154 ) , .A2( u0_u4_u3_n178 ) );
  AND3_X1 u0_u4_u3_U41 (.ZN( u0_u4_u3_n118 ) , .A2( u0_u4_u3_n124 ) , .A1( u0_u4_u3_n144 ) , .A3( u0_u4_u3_n152 ) );
  INV_X1 u0_u4_u3_U42 (.A( u0_u4_u3_n121 ) , .ZN( u0_u4_u3_n164 ) );
  NAND2_X1 u0_u4_u3_U43 (.ZN( u0_u4_u3_n133 ) , .A1( u0_u4_u3_n154 ) , .A2( u0_u4_u3_n164 ) );
  OAI211_X1 u0_u4_u3_U44 (.B( u0_u4_u3_n127 ) , .ZN( u0_u4_u3_n139 ) , .C1( u0_u4_u3_n150 ) , .C2( u0_u4_u3_n154 ) , .A( u0_u4_u3_n184 ) );
  INV_X1 u0_u4_u3_U45 (.A( u0_u4_u3_n125 ) , .ZN( u0_u4_u3_n184 ) );
  AOI221_X1 u0_u4_u3_U46 (.A( u0_u4_u3_n126 ) , .ZN( u0_u4_u3_n127 ) , .C2( u0_u4_u3_n132 ) , .C1( u0_u4_u3_n169 ) , .B2( u0_u4_u3_n170 ) , .B1( u0_u4_u3_n174 ) );
  OAI22_X1 u0_u4_u3_U47 (.A1( u0_u4_u3_n124 ) , .ZN( u0_u4_u3_n125 ) , .B2( u0_u4_u3_n145 ) , .A2( u0_u4_u3_n165 ) , .B1( u0_u4_u3_n167 ) );
  NOR2_X1 u0_u4_u3_U48 (.A1( u0_u4_u3_n113 ) , .ZN( u0_u4_u3_n131 ) , .A2( u0_u4_u3_n154 ) );
  NAND2_X1 u0_u4_u3_U49 (.A1( u0_u4_u3_n103 ) , .ZN( u0_u4_u3_n150 ) , .A2( u0_u4_u3_n99 ) );
  INV_X1 u0_u4_u3_U5 (.A( u0_u4_u3_n117 ) , .ZN( u0_u4_u3_n178 ) );
  NAND2_X1 u0_u4_u3_U50 (.A2( u0_u4_u3_n102 ) , .ZN( u0_u4_u3_n155 ) , .A1( u0_u4_u3_n97 ) );
  INV_X1 u0_u4_u3_U51 (.A( u0_u4_u3_n141 ) , .ZN( u0_u4_u3_n167 ) );
  AOI21_X1 u0_u4_u3_U52 (.B2( u0_u4_u3_n114 ) , .B1( u0_u4_u3_n146 ) , .A( u0_u4_u3_n154 ) , .ZN( u0_u4_u3_n94 ) );
  AOI21_X1 u0_u4_u3_U53 (.ZN( u0_u4_u3_n110 ) , .B2( u0_u4_u3_n142 ) , .B1( u0_u4_u3_n186 ) , .A( u0_u4_u3_n95 ) );
  INV_X1 u0_u4_u3_U54 (.A( u0_u4_u3_n145 ) , .ZN( u0_u4_u3_n186 ) );
  AOI21_X1 u0_u4_u3_U55 (.B1( u0_u4_u3_n124 ) , .A( u0_u4_u3_n149 ) , .B2( u0_u4_u3_n155 ) , .ZN( u0_u4_u3_n95 ) );
  INV_X1 u0_u4_u3_U56 (.A( u0_u4_u3_n149 ) , .ZN( u0_u4_u3_n169 ) );
  NAND2_X1 u0_u4_u3_U57 (.ZN( u0_u4_u3_n124 ) , .A1( u0_u4_u3_n96 ) , .A2( u0_u4_u3_n97 ) );
  NAND2_X1 u0_u4_u3_U58 (.A2( u0_u4_u3_n100 ) , .ZN( u0_u4_u3_n146 ) , .A1( u0_u4_u3_n96 ) );
  NAND2_X1 u0_u4_u3_U59 (.A1( u0_u4_u3_n101 ) , .ZN( u0_u4_u3_n145 ) , .A2( u0_u4_u3_n99 ) );
  AOI221_X1 u0_u4_u3_U6 (.A( u0_u4_u3_n131 ) , .C2( u0_u4_u3_n132 ) , .C1( u0_u4_u3_n133 ) , .ZN( u0_u4_u3_n134 ) , .B1( u0_u4_u3_n143 ) , .B2( u0_u4_u3_n177 ) );
  NAND2_X1 u0_u4_u3_U60 (.A1( u0_u4_u3_n100 ) , .ZN( u0_u4_u3_n156 ) , .A2( u0_u4_u3_n99 ) );
  NAND2_X1 u0_u4_u3_U61 (.A2( u0_u4_u3_n101 ) , .A1( u0_u4_u3_n104 ) , .ZN( u0_u4_u3_n148 ) );
  NAND2_X1 u0_u4_u3_U62 (.A1( u0_u4_u3_n100 ) , .A2( u0_u4_u3_n102 ) , .ZN( u0_u4_u3_n128 ) );
  NAND2_X1 u0_u4_u3_U63 (.A2( u0_u4_u3_n101 ) , .A1( u0_u4_u3_n102 ) , .ZN( u0_u4_u3_n152 ) );
  NAND2_X1 u0_u4_u3_U64 (.A2( u0_u4_u3_n101 ) , .ZN( u0_u4_u3_n114 ) , .A1( u0_u4_u3_n96 ) );
  NAND2_X1 u0_u4_u3_U65 (.ZN( u0_u4_u3_n107 ) , .A1( u0_u4_u3_n97 ) , .A2( u0_u4_u3_n99 ) );
  NAND2_X1 u0_u4_u3_U66 (.A2( u0_u4_u3_n100 ) , .A1( u0_u4_u3_n104 ) , .ZN( u0_u4_u3_n113 ) );
  NAND2_X1 u0_u4_u3_U67 (.A1( u0_u4_u3_n104 ) , .ZN( u0_u4_u3_n153 ) , .A2( u0_u4_u3_n97 ) );
  NAND2_X1 u0_u4_u3_U68 (.A2( u0_u4_u3_n103 ) , .A1( u0_u4_u3_n104 ) , .ZN( u0_u4_u3_n130 ) );
  NAND2_X1 u0_u4_u3_U69 (.A2( u0_u4_u3_n103 ) , .ZN( u0_u4_u3_n144 ) , .A1( u0_u4_u3_n96 ) );
  OAI22_X1 u0_u4_u3_U7 (.B2( u0_u4_u3_n147 ) , .A2( u0_u4_u3_n148 ) , .ZN( u0_u4_u3_n160 ) , .B1( u0_u4_u3_n165 ) , .A1( u0_u4_u3_n168 ) );
  NAND2_X1 u0_u4_u3_U70 (.A1( u0_u4_u3_n102 ) , .A2( u0_u4_u3_n103 ) , .ZN( u0_u4_u3_n108 ) );
  NOR2_X1 u0_u4_u3_U71 (.A2( u0_u4_X_19 ) , .A1( u0_u4_X_20 ) , .ZN( u0_u4_u3_n99 ) );
  NOR2_X1 u0_u4_u3_U72 (.A2( u0_u4_X_21 ) , .A1( u0_u4_X_24 ) , .ZN( u0_u4_u3_n103 ) );
  NOR2_X1 u0_u4_u3_U73 (.A2( u0_u4_X_24 ) , .A1( u0_u4_u3_n171 ) , .ZN( u0_u4_u3_n97 ) );
  NOR2_X1 u0_u4_u3_U74 (.A2( u0_u4_X_23 ) , .ZN( u0_u4_u3_n141 ) , .A1( u0_u4_u3_n166 ) );
  NOR2_X1 u0_u4_u3_U75 (.A2( u0_u4_X_19 ) , .A1( u0_u4_u3_n172 ) , .ZN( u0_u4_u3_n96 ) );
  NAND2_X1 u0_u4_u3_U76 (.A1( u0_u4_X_22 ) , .A2( u0_u4_X_23 ) , .ZN( u0_u4_u3_n154 ) );
  NAND2_X1 u0_u4_u3_U77 (.A1( u0_u4_X_23 ) , .ZN( u0_u4_u3_n149 ) , .A2( u0_u4_u3_n166 ) );
  NOR2_X1 u0_u4_u3_U78 (.A2( u0_u4_X_22 ) , .A1( u0_u4_X_23 ) , .ZN( u0_u4_u3_n121 ) );
  AND2_X1 u0_u4_u3_U79 (.A1( u0_u4_X_24 ) , .ZN( u0_u4_u3_n101 ) , .A2( u0_u4_u3_n171 ) );
  AND3_X1 u0_u4_u3_U8 (.A3( u0_u4_u3_n144 ) , .A2( u0_u4_u3_n145 ) , .A1( u0_u4_u3_n146 ) , .ZN( u0_u4_u3_n147 ) );
  AND2_X1 u0_u4_u3_U80 (.A1( u0_u4_X_19 ) , .ZN( u0_u4_u3_n102 ) , .A2( u0_u4_u3_n172 ) );
  AND2_X1 u0_u4_u3_U81 (.A1( u0_u4_X_21 ) , .A2( u0_u4_X_24 ) , .ZN( u0_u4_u3_n100 ) );
  AND2_X1 u0_u4_u3_U82 (.A2( u0_u4_X_19 ) , .A1( u0_u4_X_20 ) , .ZN( u0_u4_u3_n104 ) );
  INV_X1 u0_u4_u3_U83 (.A( u0_u4_X_22 ) , .ZN( u0_u4_u3_n166 ) );
  INV_X1 u0_u4_u3_U84 (.A( u0_u4_X_21 ) , .ZN( u0_u4_u3_n171 ) );
  INV_X1 u0_u4_u3_U85 (.A( u0_u4_X_20 ) , .ZN( u0_u4_u3_n172 ) );
  OR4_X1 u0_u4_u3_U86 (.ZN( u0_out4_10 ) , .A4( u0_u4_u3_n136 ) , .A3( u0_u4_u3_n137 ) , .A1( u0_u4_u3_n138 ) , .A2( u0_u4_u3_n139 ) );
  OAI222_X1 u0_u4_u3_U87 (.C1( u0_u4_u3_n128 ) , .ZN( u0_u4_u3_n137 ) , .B1( u0_u4_u3_n148 ) , .A2( u0_u4_u3_n150 ) , .B2( u0_u4_u3_n154 ) , .C2( u0_u4_u3_n164 ) , .A1( u0_u4_u3_n167 ) );
  OAI221_X1 u0_u4_u3_U88 (.A( u0_u4_u3_n134 ) , .B2( u0_u4_u3_n135 ) , .ZN( u0_u4_u3_n136 ) , .C1( u0_u4_u3_n149 ) , .B1( u0_u4_u3_n151 ) , .C2( u0_u4_u3_n183 ) );
  NAND4_X1 u0_u4_u3_U89 (.ZN( u0_out4_26 ) , .A4( u0_u4_u3_n109 ) , .A3( u0_u4_u3_n110 ) , .A2( u0_u4_u3_n111 ) , .A1( u0_u4_u3_n173 ) );
  INV_X1 u0_u4_u3_U9 (.A( u0_u4_u3_n143 ) , .ZN( u0_u4_u3_n168 ) );
  INV_X1 u0_u4_u3_U90 (.ZN( u0_u4_u3_n173 ) , .A( u0_u4_u3_n94 ) );
  OAI21_X1 u0_u4_u3_U91 (.ZN( u0_u4_u3_n111 ) , .B2( u0_u4_u3_n117 ) , .A( u0_u4_u3_n133 ) , .B1( u0_u4_u3_n176 ) );
  NAND4_X1 u0_u4_u3_U92 (.ZN( u0_out4_20 ) , .A4( u0_u4_u3_n122 ) , .A3( u0_u4_u3_n123 ) , .A1( u0_u4_u3_n175 ) , .A2( u0_u4_u3_n180 ) );
  INV_X1 u0_u4_u3_U93 (.A( u0_u4_u3_n126 ) , .ZN( u0_u4_u3_n180 ) );
  INV_X1 u0_u4_u3_U94 (.A( u0_u4_u3_n112 ) , .ZN( u0_u4_u3_n175 ) );
  NAND4_X1 u0_u4_u3_U95 (.ZN( u0_out4_1 ) , .A4( u0_u4_u3_n161 ) , .A3( u0_u4_u3_n162 ) , .A2( u0_u4_u3_n163 ) , .A1( u0_u4_u3_n185 ) );
  NAND2_X1 u0_u4_u3_U96 (.ZN( u0_u4_u3_n163 ) , .A2( u0_u4_u3_n170 ) , .A1( u0_u4_u3_n176 ) );
  AOI22_X1 u0_u4_u3_U97 (.B2( u0_u4_u3_n140 ) , .B1( u0_u4_u3_n141 ) , .A2( u0_u4_u3_n142 ) , .ZN( u0_u4_u3_n162 ) , .A1( u0_u4_u3_n177 ) );
  NAND3_X1 u0_u4_u3_U98 (.A1( u0_u4_u3_n114 ) , .ZN( u0_u4_u3_n115 ) , .A2( u0_u4_u3_n145 ) , .A3( u0_u4_u3_n153 ) );
  NAND3_X1 u0_u4_u3_U99 (.ZN( u0_u4_u3_n129 ) , .A2( u0_u4_u3_n144 ) , .A1( u0_u4_u3_n153 ) , .A3( u0_u4_u3_n182 ) );
  OAI22_X1 u0_u4_u4_U10 (.B2( u0_u4_u4_n135 ) , .ZN( u0_u4_u4_n137 ) , .B1( u0_u4_u4_n153 ) , .A1( u0_u4_u4_n155 ) , .A2( u0_u4_u4_n171 ) );
  AND3_X1 u0_u4_u4_U11 (.A2( u0_u4_u4_n134 ) , .ZN( u0_u4_u4_n135 ) , .A3( u0_u4_u4_n145 ) , .A1( u0_u4_u4_n157 ) );
  NAND2_X1 u0_u4_u4_U12 (.ZN( u0_u4_u4_n132 ) , .A2( u0_u4_u4_n170 ) , .A1( u0_u4_u4_n173 ) );
  AOI21_X1 u0_u4_u4_U13 (.B2( u0_u4_u4_n160 ) , .B1( u0_u4_u4_n161 ) , .ZN( u0_u4_u4_n162 ) , .A( u0_u4_u4_n170 ) );
  AOI21_X1 u0_u4_u4_U14 (.ZN( u0_u4_u4_n107 ) , .B2( u0_u4_u4_n143 ) , .A( u0_u4_u4_n174 ) , .B1( u0_u4_u4_n184 ) );
  AOI21_X1 u0_u4_u4_U15 (.B2( u0_u4_u4_n158 ) , .B1( u0_u4_u4_n159 ) , .ZN( u0_u4_u4_n163 ) , .A( u0_u4_u4_n174 ) );
  AOI21_X1 u0_u4_u4_U16 (.A( u0_u4_u4_n153 ) , .B2( u0_u4_u4_n154 ) , .B1( u0_u4_u4_n155 ) , .ZN( u0_u4_u4_n165 ) );
  AOI21_X1 u0_u4_u4_U17 (.A( u0_u4_u4_n156 ) , .B2( u0_u4_u4_n157 ) , .ZN( u0_u4_u4_n164 ) , .B1( u0_u4_u4_n184 ) );
  INV_X1 u0_u4_u4_U18 (.A( u0_u4_u4_n138 ) , .ZN( u0_u4_u4_n170 ) );
  AND2_X1 u0_u4_u4_U19 (.A2( u0_u4_u4_n120 ) , .ZN( u0_u4_u4_n155 ) , .A1( u0_u4_u4_n160 ) );
  INV_X1 u0_u4_u4_U20 (.A( u0_u4_u4_n156 ) , .ZN( u0_u4_u4_n175 ) );
  NAND2_X1 u0_u4_u4_U21 (.A2( u0_u4_u4_n118 ) , .ZN( u0_u4_u4_n131 ) , .A1( u0_u4_u4_n147 ) );
  NAND2_X1 u0_u4_u4_U22 (.A1( u0_u4_u4_n119 ) , .A2( u0_u4_u4_n120 ) , .ZN( u0_u4_u4_n130 ) );
  NAND2_X1 u0_u4_u4_U23 (.ZN( u0_u4_u4_n117 ) , .A2( u0_u4_u4_n118 ) , .A1( u0_u4_u4_n148 ) );
  NAND2_X1 u0_u4_u4_U24 (.ZN( u0_u4_u4_n129 ) , .A1( u0_u4_u4_n134 ) , .A2( u0_u4_u4_n148 ) );
  AND3_X1 u0_u4_u4_U25 (.A1( u0_u4_u4_n119 ) , .A2( u0_u4_u4_n143 ) , .A3( u0_u4_u4_n154 ) , .ZN( u0_u4_u4_n161 ) );
  AND2_X1 u0_u4_u4_U26 (.A1( u0_u4_u4_n145 ) , .A2( u0_u4_u4_n147 ) , .ZN( u0_u4_u4_n159 ) );
  OR3_X1 u0_u4_u4_U27 (.A3( u0_u4_u4_n114 ) , .A2( u0_u4_u4_n115 ) , .A1( u0_u4_u4_n116 ) , .ZN( u0_u4_u4_n136 ) );
  AOI21_X1 u0_u4_u4_U28 (.A( u0_u4_u4_n113 ) , .ZN( u0_u4_u4_n116 ) , .B2( u0_u4_u4_n173 ) , .B1( u0_u4_u4_n174 ) );
  AOI21_X1 u0_u4_u4_U29 (.ZN( u0_u4_u4_n115 ) , .B2( u0_u4_u4_n145 ) , .B1( u0_u4_u4_n146 ) , .A( u0_u4_u4_n156 ) );
  NOR2_X1 u0_u4_u4_U3 (.ZN( u0_u4_u4_n121 ) , .A1( u0_u4_u4_n181 ) , .A2( u0_u4_u4_n182 ) );
  OAI22_X1 u0_u4_u4_U30 (.ZN( u0_u4_u4_n114 ) , .A2( u0_u4_u4_n121 ) , .B1( u0_u4_u4_n160 ) , .B2( u0_u4_u4_n170 ) , .A1( u0_u4_u4_n171 ) );
  INV_X1 u0_u4_u4_U31 (.A( u0_u4_u4_n158 ) , .ZN( u0_u4_u4_n182 ) );
  INV_X1 u0_u4_u4_U32 (.ZN( u0_u4_u4_n181 ) , .A( u0_u4_u4_n96 ) );
  INV_X1 u0_u4_u4_U33 (.A( u0_u4_u4_n144 ) , .ZN( u0_u4_u4_n179 ) );
  INV_X1 u0_u4_u4_U34 (.A( u0_u4_u4_n157 ) , .ZN( u0_u4_u4_n178 ) );
  NAND2_X1 u0_u4_u4_U35 (.A2( u0_u4_u4_n154 ) , .A1( u0_u4_u4_n96 ) , .ZN( u0_u4_u4_n97 ) );
  INV_X1 u0_u4_u4_U36 (.ZN( u0_u4_u4_n186 ) , .A( u0_u4_u4_n95 ) );
  OAI221_X1 u0_u4_u4_U37 (.C1( u0_u4_u4_n134 ) , .B1( u0_u4_u4_n158 ) , .B2( u0_u4_u4_n171 ) , .C2( u0_u4_u4_n173 ) , .A( u0_u4_u4_n94 ) , .ZN( u0_u4_u4_n95 ) );
  AOI222_X1 u0_u4_u4_U38 (.B2( u0_u4_u4_n132 ) , .A1( u0_u4_u4_n138 ) , .C2( u0_u4_u4_n175 ) , .A2( u0_u4_u4_n179 ) , .C1( u0_u4_u4_n181 ) , .B1( u0_u4_u4_n185 ) , .ZN( u0_u4_u4_n94 ) );
  INV_X1 u0_u4_u4_U39 (.A( u0_u4_u4_n113 ) , .ZN( u0_u4_u4_n185 ) );
  INV_X1 u0_u4_u4_U4 (.A( u0_u4_u4_n117 ) , .ZN( u0_u4_u4_n184 ) );
  INV_X1 u0_u4_u4_U40 (.A( u0_u4_u4_n143 ) , .ZN( u0_u4_u4_n183 ) );
  NOR2_X1 u0_u4_u4_U41 (.ZN( u0_u4_u4_n138 ) , .A1( u0_u4_u4_n168 ) , .A2( u0_u4_u4_n169 ) );
  NOR2_X1 u0_u4_u4_U42 (.A1( u0_u4_u4_n150 ) , .A2( u0_u4_u4_n152 ) , .ZN( u0_u4_u4_n153 ) );
  NOR2_X1 u0_u4_u4_U43 (.A2( u0_u4_u4_n128 ) , .A1( u0_u4_u4_n138 ) , .ZN( u0_u4_u4_n156 ) );
  AOI22_X1 u0_u4_u4_U44 (.B2( u0_u4_u4_n122 ) , .A1( u0_u4_u4_n123 ) , .ZN( u0_u4_u4_n124 ) , .B1( u0_u4_u4_n128 ) , .A2( u0_u4_u4_n172 ) );
  INV_X1 u0_u4_u4_U45 (.A( u0_u4_u4_n153 ) , .ZN( u0_u4_u4_n172 ) );
  NAND2_X1 u0_u4_u4_U46 (.A2( u0_u4_u4_n120 ) , .ZN( u0_u4_u4_n123 ) , .A1( u0_u4_u4_n161 ) );
  AOI22_X1 u0_u4_u4_U47 (.B2( u0_u4_u4_n132 ) , .A2( u0_u4_u4_n133 ) , .ZN( u0_u4_u4_n140 ) , .A1( u0_u4_u4_n150 ) , .B1( u0_u4_u4_n179 ) );
  NAND2_X1 u0_u4_u4_U48 (.ZN( u0_u4_u4_n133 ) , .A2( u0_u4_u4_n146 ) , .A1( u0_u4_u4_n154 ) );
  NAND2_X1 u0_u4_u4_U49 (.A1( u0_u4_u4_n103 ) , .ZN( u0_u4_u4_n154 ) , .A2( u0_u4_u4_n98 ) );
  NOR4_X1 u0_u4_u4_U5 (.A4( u0_u4_u4_n106 ) , .A3( u0_u4_u4_n107 ) , .A2( u0_u4_u4_n108 ) , .A1( u0_u4_u4_n109 ) , .ZN( u0_u4_u4_n110 ) );
  NAND2_X1 u0_u4_u4_U50 (.A1( u0_u4_u4_n101 ) , .ZN( u0_u4_u4_n158 ) , .A2( u0_u4_u4_n99 ) );
  AOI21_X1 u0_u4_u4_U51 (.ZN( u0_u4_u4_n127 ) , .A( u0_u4_u4_n136 ) , .B2( u0_u4_u4_n150 ) , .B1( u0_u4_u4_n180 ) );
  INV_X1 u0_u4_u4_U52 (.A( u0_u4_u4_n160 ) , .ZN( u0_u4_u4_n180 ) );
  NAND2_X1 u0_u4_u4_U53 (.A2( u0_u4_u4_n104 ) , .A1( u0_u4_u4_n105 ) , .ZN( u0_u4_u4_n146 ) );
  NAND2_X1 u0_u4_u4_U54 (.A2( u0_u4_u4_n101 ) , .A1( u0_u4_u4_n102 ) , .ZN( u0_u4_u4_n160 ) );
  NAND2_X1 u0_u4_u4_U55 (.ZN( u0_u4_u4_n134 ) , .A1( u0_u4_u4_n98 ) , .A2( u0_u4_u4_n99 ) );
  NAND2_X1 u0_u4_u4_U56 (.A1( u0_u4_u4_n103 ) , .A2( u0_u4_u4_n104 ) , .ZN( u0_u4_u4_n143 ) );
  NAND2_X1 u0_u4_u4_U57 (.A2( u0_u4_u4_n105 ) , .ZN( u0_u4_u4_n145 ) , .A1( u0_u4_u4_n98 ) );
  NAND2_X1 u0_u4_u4_U58 (.A1( u0_u4_u4_n100 ) , .A2( u0_u4_u4_n105 ) , .ZN( u0_u4_u4_n120 ) );
  NAND2_X1 u0_u4_u4_U59 (.A1( u0_u4_u4_n102 ) , .A2( u0_u4_u4_n104 ) , .ZN( u0_u4_u4_n148 ) );
  AOI21_X1 u0_u4_u4_U6 (.ZN( u0_u4_u4_n106 ) , .B2( u0_u4_u4_n146 ) , .B1( u0_u4_u4_n158 ) , .A( u0_u4_u4_n170 ) );
  NAND2_X1 u0_u4_u4_U60 (.A2( u0_u4_u4_n100 ) , .A1( u0_u4_u4_n103 ) , .ZN( u0_u4_u4_n157 ) );
  INV_X1 u0_u4_u4_U61 (.A( u0_u4_u4_n150 ) , .ZN( u0_u4_u4_n173 ) );
  INV_X1 u0_u4_u4_U62 (.A( u0_u4_u4_n152 ) , .ZN( u0_u4_u4_n171 ) );
  NAND2_X1 u0_u4_u4_U63 (.A1( u0_u4_u4_n100 ) , .ZN( u0_u4_u4_n118 ) , .A2( u0_u4_u4_n99 ) );
  NAND2_X1 u0_u4_u4_U64 (.A2( u0_u4_u4_n100 ) , .A1( u0_u4_u4_n102 ) , .ZN( u0_u4_u4_n144 ) );
  NAND2_X1 u0_u4_u4_U65 (.A2( u0_u4_u4_n101 ) , .A1( u0_u4_u4_n105 ) , .ZN( u0_u4_u4_n96 ) );
  INV_X1 u0_u4_u4_U66 (.A( u0_u4_u4_n128 ) , .ZN( u0_u4_u4_n174 ) );
  NAND2_X1 u0_u4_u4_U67 (.A2( u0_u4_u4_n102 ) , .ZN( u0_u4_u4_n119 ) , .A1( u0_u4_u4_n98 ) );
  NAND2_X1 u0_u4_u4_U68 (.A2( u0_u4_u4_n101 ) , .A1( u0_u4_u4_n103 ) , .ZN( u0_u4_u4_n147 ) );
  NAND2_X1 u0_u4_u4_U69 (.A2( u0_u4_u4_n104 ) , .ZN( u0_u4_u4_n113 ) , .A1( u0_u4_u4_n99 ) );
  AOI21_X1 u0_u4_u4_U7 (.ZN( u0_u4_u4_n108 ) , .B2( u0_u4_u4_n134 ) , .B1( u0_u4_u4_n155 ) , .A( u0_u4_u4_n156 ) );
  NOR2_X1 u0_u4_u4_U70 (.A2( u0_u4_X_28 ) , .ZN( u0_u4_u4_n150 ) , .A1( u0_u4_u4_n168 ) );
  NOR2_X1 u0_u4_u4_U71 (.A2( u0_u4_X_29 ) , .ZN( u0_u4_u4_n152 ) , .A1( u0_u4_u4_n169 ) );
  NOR2_X1 u0_u4_u4_U72 (.A2( u0_u4_X_30 ) , .ZN( u0_u4_u4_n105 ) , .A1( u0_u4_u4_n176 ) );
  NOR2_X1 u0_u4_u4_U73 (.A2( u0_u4_X_26 ) , .ZN( u0_u4_u4_n100 ) , .A1( u0_u4_u4_n177 ) );
  NOR2_X1 u0_u4_u4_U74 (.A2( u0_u4_X_28 ) , .A1( u0_u4_X_29 ) , .ZN( u0_u4_u4_n128 ) );
  NOR2_X1 u0_u4_u4_U75 (.A2( u0_u4_X_27 ) , .A1( u0_u4_X_30 ) , .ZN( u0_u4_u4_n102 ) );
  NOR2_X1 u0_u4_u4_U76 (.A2( u0_u4_X_25 ) , .A1( u0_u4_X_26 ) , .ZN( u0_u4_u4_n98 ) );
  AND2_X1 u0_u4_u4_U77 (.A2( u0_u4_X_25 ) , .A1( u0_u4_X_26 ) , .ZN( u0_u4_u4_n104 ) );
  AND2_X1 u0_u4_u4_U78 (.A1( u0_u4_X_30 ) , .A2( u0_u4_u4_n176 ) , .ZN( u0_u4_u4_n99 ) );
  AND2_X1 u0_u4_u4_U79 (.A1( u0_u4_X_26 ) , .ZN( u0_u4_u4_n101 ) , .A2( u0_u4_u4_n177 ) );
  AOI21_X1 u0_u4_u4_U8 (.ZN( u0_u4_u4_n109 ) , .A( u0_u4_u4_n153 ) , .B1( u0_u4_u4_n159 ) , .B2( u0_u4_u4_n184 ) );
  AND2_X1 u0_u4_u4_U80 (.A1( u0_u4_X_27 ) , .A2( u0_u4_X_30 ) , .ZN( u0_u4_u4_n103 ) );
  INV_X1 u0_u4_u4_U81 (.A( u0_u4_X_28 ) , .ZN( u0_u4_u4_n169 ) );
  INV_X1 u0_u4_u4_U82 (.A( u0_u4_X_29 ) , .ZN( u0_u4_u4_n168 ) );
  INV_X1 u0_u4_u4_U83 (.A( u0_u4_X_25 ) , .ZN( u0_u4_u4_n177 ) );
  INV_X1 u0_u4_u4_U84 (.A( u0_u4_X_27 ) , .ZN( u0_u4_u4_n176 ) );
  NAND4_X1 u0_u4_u4_U85 (.ZN( u0_out4_25 ) , .A4( u0_u4_u4_n139 ) , .A3( u0_u4_u4_n140 ) , .A2( u0_u4_u4_n141 ) , .A1( u0_u4_u4_n142 ) );
  OAI21_X1 u0_u4_u4_U86 (.B2( u0_u4_u4_n131 ) , .ZN( u0_u4_u4_n141 ) , .A( u0_u4_u4_n175 ) , .B1( u0_u4_u4_n183 ) );
  OAI21_X1 u0_u4_u4_U87 (.A( u0_u4_u4_n128 ) , .B2( u0_u4_u4_n129 ) , .B1( u0_u4_u4_n130 ) , .ZN( u0_u4_u4_n142 ) );
  NAND4_X1 u0_u4_u4_U88 (.ZN( u0_out4_14 ) , .A4( u0_u4_u4_n124 ) , .A3( u0_u4_u4_n125 ) , .A2( u0_u4_u4_n126 ) , .A1( u0_u4_u4_n127 ) );
  AOI22_X1 u0_u4_u4_U89 (.B2( u0_u4_u4_n117 ) , .ZN( u0_u4_u4_n126 ) , .A1( u0_u4_u4_n129 ) , .B1( u0_u4_u4_n152 ) , .A2( u0_u4_u4_n175 ) );
  AOI211_X1 u0_u4_u4_U9 (.B( u0_u4_u4_n136 ) , .A( u0_u4_u4_n137 ) , .C2( u0_u4_u4_n138 ) , .ZN( u0_u4_u4_n139 ) , .C1( u0_u4_u4_n182 ) );
  AOI22_X1 u0_u4_u4_U90 (.ZN( u0_u4_u4_n125 ) , .B2( u0_u4_u4_n131 ) , .A2( u0_u4_u4_n132 ) , .B1( u0_u4_u4_n138 ) , .A1( u0_u4_u4_n178 ) );
  NAND4_X1 u0_u4_u4_U91 (.ZN( u0_out4_8 ) , .A4( u0_u4_u4_n110 ) , .A3( u0_u4_u4_n111 ) , .A2( u0_u4_u4_n112 ) , .A1( u0_u4_u4_n186 ) );
  NAND2_X1 u0_u4_u4_U92 (.ZN( u0_u4_u4_n112 ) , .A2( u0_u4_u4_n130 ) , .A1( u0_u4_u4_n150 ) );
  AOI22_X1 u0_u4_u4_U93 (.ZN( u0_u4_u4_n111 ) , .B2( u0_u4_u4_n132 ) , .A1( u0_u4_u4_n152 ) , .B1( u0_u4_u4_n178 ) , .A2( u0_u4_u4_n97 ) );
  AOI22_X1 u0_u4_u4_U94 (.B2( u0_u4_u4_n149 ) , .B1( u0_u4_u4_n150 ) , .A2( u0_u4_u4_n151 ) , .A1( u0_u4_u4_n152 ) , .ZN( u0_u4_u4_n167 ) );
  NOR4_X1 u0_u4_u4_U95 (.A4( u0_u4_u4_n162 ) , .A3( u0_u4_u4_n163 ) , .A2( u0_u4_u4_n164 ) , .A1( u0_u4_u4_n165 ) , .ZN( u0_u4_u4_n166 ) );
  NAND3_X1 u0_u4_u4_U96 (.ZN( u0_out4_3 ) , .A3( u0_u4_u4_n166 ) , .A1( u0_u4_u4_n167 ) , .A2( u0_u4_u4_n186 ) );
  NAND3_X1 u0_u4_u4_U97 (.A3( u0_u4_u4_n146 ) , .A2( u0_u4_u4_n147 ) , .A1( u0_u4_u4_n148 ) , .ZN( u0_u4_u4_n149 ) );
  NAND3_X1 u0_u4_u4_U98 (.A3( u0_u4_u4_n143 ) , .A2( u0_u4_u4_n144 ) , .A1( u0_u4_u4_n145 ) , .ZN( u0_u4_u4_n151 ) );
  NAND3_X1 u0_u4_u4_U99 (.A3( u0_u4_u4_n121 ) , .ZN( u0_u4_u4_n122 ) , .A2( u0_u4_u4_n144 ) , .A1( u0_u4_u4_n154 ) );
  NOR2_X1 u0_u4_u5_U10 (.ZN( u0_u4_u5_n135 ) , .A1( u0_u4_u5_n173 ) , .A2( u0_u4_u5_n176 ) );
  NOR3_X1 u0_u4_u5_U100 (.A3( u0_u4_u5_n141 ) , .A1( u0_u4_u5_n142 ) , .ZN( u0_u4_u5_n143 ) , .A2( u0_u4_u5_n191 ) );
  NAND4_X1 u0_u4_u5_U101 (.ZN( u0_out4_4 ) , .A4( u0_u4_u5_n112 ) , .A2( u0_u4_u5_n113 ) , .A1( u0_u4_u5_n114 ) , .A3( u0_u4_u5_n195 ) );
  AOI211_X1 u0_u4_u5_U102 (.A( u0_u4_u5_n110 ) , .C1( u0_u4_u5_n111 ) , .ZN( u0_u4_u5_n112 ) , .B( u0_u4_u5_n118 ) , .C2( u0_u4_u5_n177 ) );
  INV_X1 u0_u4_u5_U103 (.A( u0_u4_u5_n102 ) , .ZN( u0_u4_u5_n195 ) );
  NAND3_X1 u0_u4_u5_U104 (.A2( u0_u4_u5_n154 ) , .A3( u0_u4_u5_n158 ) , .A1( u0_u4_u5_n161 ) , .ZN( u0_u4_u5_n99 ) );
  INV_X1 u0_u4_u5_U11 (.A( u0_u4_u5_n121 ) , .ZN( u0_u4_u5_n177 ) );
  NOR2_X1 u0_u4_u5_U12 (.ZN( u0_u4_u5_n160 ) , .A2( u0_u4_u5_n173 ) , .A1( u0_u4_u5_n177 ) );
  INV_X1 u0_u4_u5_U13 (.A( u0_u4_u5_n150 ) , .ZN( u0_u4_u5_n174 ) );
  AOI21_X1 u0_u4_u5_U14 (.A( u0_u4_u5_n160 ) , .B2( u0_u4_u5_n161 ) , .ZN( u0_u4_u5_n162 ) , .B1( u0_u4_u5_n192 ) );
  INV_X1 u0_u4_u5_U15 (.A( u0_u4_u5_n159 ) , .ZN( u0_u4_u5_n192 ) );
  AOI21_X1 u0_u4_u5_U16 (.A( u0_u4_u5_n156 ) , .B2( u0_u4_u5_n157 ) , .B1( u0_u4_u5_n158 ) , .ZN( u0_u4_u5_n163 ) );
  AOI21_X1 u0_u4_u5_U17 (.B2( u0_u4_u5_n139 ) , .B1( u0_u4_u5_n140 ) , .ZN( u0_u4_u5_n141 ) , .A( u0_u4_u5_n150 ) );
  OAI21_X1 u0_u4_u5_U18 (.A( u0_u4_u5_n133 ) , .B2( u0_u4_u5_n134 ) , .B1( u0_u4_u5_n135 ) , .ZN( u0_u4_u5_n142 ) );
  OAI21_X1 u0_u4_u5_U19 (.ZN( u0_u4_u5_n133 ) , .B2( u0_u4_u5_n147 ) , .A( u0_u4_u5_n173 ) , .B1( u0_u4_u5_n188 ) );
  NAND2_X1 u0_u4_u5_U20 (.A2( u0_u4_u5_n119 ) , .A1( u0_u4_u5_n123 ) , .ZN( u0_u4_u5_n137 ) );
  INV_X1 u0_u4_u5_U21 (.A( u0_u4_u5_n155 ) , .ZN( u0_u4_u5_n194 ) );
  NAND2_X1 u0_u4_u5_U22 (.A1( u0_u4_u5_n121 ) , .ZN( u0_u4_u5_n132 ) , .A2( u0_u4_u5_n172 ) );
  NAND2_X1 u0_u4_u5_U23 (.A2( u0_u4_u5_n122 ) , .ZN( u0_u4_u5_n136 ) , .A1( u0_u4_u5_n154 ) );
  NAND2_X1 u0_u4_u5_U24 (.A2( u0_u4_u5_n119 ) , .A1( u0_u4_u5_n120 ) , .ZN( u0_u4_u5_n159 ) );
  INV_X1 u0_u4_u5_U25 (.A( u0_u4_u5_n156 ) , .ZN( u0_u4_u5_n175 ) );
  INV_X1 u0_u4_u5_U26 (.A( u0_u4_u5_n158 ) , .ZN( u0_u4_u5_n188 ) );
  INV_X1 u0_u4_u5_U27 (.A( u0_u4_u5_n152 ) , .ZN( u0_u4_u5_n179 ) );
  INV_X1 u0_u4_u5_U28 (.A( u0_u4_u5_n140 ) , .ZN( u0_u4_u5_n182 ) );
  INV_X1 u0_u4_u5_U29 (.A( u0_u4_u5_n151 ) , .ZN( u0_u4_u5_n183 ) );
  NOR2_X1 u0_u4_u5_U3 (.ZN( u0_u4_u5_n134 ) , .A1( u0_u4_u5_n183 ) , .A2( u0_u4_u5_n190 ) );
  INV_X1 u0_u4_u5_U30 (.A( u0_u4_u5_n123 ) , .ZN( u0_u4_u5_n185 ) );
  INV_X1 u0_u4_u5_U31 (.A( u0_u4_u5_n161 ) , .ZN( u0_u4_u5_n184 ) );
  INV_X1 u0_u4_u5_U32 (.A( u0_u4_u5_n139 ) , .ZN( u0_u4_u5_n189 ) );
  INV_X1 u0_u4_u5_U33 (.A( u0_u4_u5_n157 ) , .ZN( u0_u4_u5_n190 ) );
  INV_X1 u0_u4_u5_U34 (.A( u0_u4_u5_n120 ) , .ZN( u0_u4_u5_n193 ) );
  NAND2_X1 u0_u4_u5_U35 (.ZN( u0_u4_u5_n111 ) , .A1( u0_u4_u5_n140 ) , .A2( u0_u4_u5_n155 ) );
  INV_X1 u0_u4_u5_U36 (.A( u0_u4_u5_n117 ) , .ZN( u0_u4_u5_n196 ) );
  OAI221_X1 u0_u4_u5_U37 (.A( u0_u4_u5_n116 ) , .ZN( u0_u4_u5_n117 ) , .B2( u0_u4_u5_n119 ) , .C1( u0_u4_u5_n153 ) , .C2( u0_u4_u5_n158 ) , .B1( u0_u4_u5_n172 ) );
  AOI222_X1 u0_u4_u5_U38 (.ZN( u0_u4_u5_n116 ) , .B2( u0_u4_u5_n145 ) , .C1( u0_u4_u5_n148 ) , .A2( u0_u4_u5_n174 ) , .C2( u0_u4_u5_n177 ) , .B1( u0_u4_u5_n187 ) , .A1( u0_u4_u5_n193 ) );
  INV_X1 u0_u4_u5_U39 (.A( u0_u4_u5_n115 ) , .ZN( u0_u4_u5_n187 ) );
  INV_X1 u0_u4_u5_U4 (.A( u0_u4_u5_n138 ) , .ZN( u0_u4_u5_n191 ) );
  NOR2_X1 u0_u4_u5_U40 (.ZN( u0_u4_u5_n100 ) , .A1( u0_u4_u5_n170 ) , .A2( u0_u4_u5_n180 ) );
  OAI221_X1 u0_u4_u5_U41 (.A( u0_u4_u5_n101 ) , .ZN( u0_u4_u5_n102 ) , .C2( u0_u4_u5_n115 ) , .C1( u0_u4_u5_n126 ) , .B1( u0_u4_u5_n134 ) , .B2( u0_u4_u5_n160 ) );
  OAI21_X1 u0_u4_u5_U42 (.ZN( u0_u4_u5_n101 ) , .B1( u0_u4_u5_n137 ) , .A( u0_u4_u5_n146 ) , .B2( u0_u4_u5_n147 ) );
  AOI22_X1 u0_u4_u5_U43 (.B2( u0_u4_u5_n131 ) , .A2( u0_u4_u5_n146 ) , .ZN( u0_u4_u5_n169 ) , .B1( u0_u4_u5_n174 ) , .A1( u0_u4_u5_n185 ) );
  NOR2_X1 u0_u4_u5_U44 (.A1( u0_u4_u5_n146 ) , .ZN( u0_u4_u5_n150 ) , .A2( u0_u4_u5_n173 ) );
  AOI21_X1 u0_u4_u5_U45 (.A( u0_u4_u5_n118 ) , .B2( u0_u4_u5_n145 ) , .ZN( u0_u4_u5_n168 ) , .B1( u0_u4_u5_n186 ) );
  INV_X1 u0_u4_u5_U46 (.A( u0_u4_u5_n122 ) , .ZN( u0_u4_u5_n186 ) );
  NOR2_X1 u0_u4_u5_U47 (.A1( u0_u4_u5_n146 ) , .ZN( u0_u4_u5_n152 ) , .A2( u0_u4_u5_n176 ) );
  NOR2_X1 u0_u4_u5_U48 (.A1( u0_u4_u5_n115 ) , .ZN( u0_u4_u5_n118 ) , .A2( u0_u4_u5_n153 ) );
  NOR2_X1 u0_u4_u5_U49 (.A2( u0_u4_u5_n145 ) , .ZN( u0_u4_u5_n156 ) , .A1( u0_u4_u5_n174 ) );
  OAI21_X1 u0_u4_u5_U5 (.B2( u0_u4_u5_n136 ) , .B1( u0_u4_u5_n137 ) , .ZN( u0_u4_u5_n138 ) , .A( u0_u4_u5_n177 ) );
  NOR2_X1 u0_u4_u5_U50 (.ZN( u0_u4_u5_n121 ) , .A2( u0_u4_u5_n145 ) , .A1( u0_u4_u5_n176 ) );
  AOI22_X1 u0_u4_u5_U51 (.ZN( u0_u4_u5_n114 ) , .A2( u0_u4_u5_n137 ) , .A1( u0_u4_u5_n145 ) , .B2( u0_u4_u5_n175 ) , .B1( u0_u4_u5_n193 ) );
  OAI211_X1 u0_u4_u5_U52 (.B( u0_u4_u5_n124 ) , .A( u0_u4_u5_n125 ) , .C2( u0_u4_u5_n126 ) , .C1( u0_u4_u5_n127 ) , .ZN( u0_u4_u5_n128 ) );
  NOR3_X1 u0_u4_u5_U53 (.ZN( u0_u4_u5_n127 ) , .A1( u0_u4_u5_n136 ) , .A3( u0_u4_u5_n148 ) , .A2( u0_u4_u5_n182 ) );
  OAI21_X1 u0_u4_u5_U54 (.ZN( u0_u4_u5_n124 ) , .A( u0_u4_u5_n177 ) , .B2( u0_u4_u5_n183 ) , .B1( u0_u4_u5_n189 ) );
  OAI21_X1 u0_u4_u5_U55 (.ZN( u0_u4_u5_n125 ) , .A( u0_u4_u5_n174 ) , .B2( u0_u4_u5_n185 ) , .B1( u0_u4_u5_n190 ) );
  AOI21_X1 u0_u4_u5_U56 (.A( u0_u4_u5_n153 ) , .B2( u0_u4_u5_n154 ) , .B1( u0_u4_u5_n155 ) , .ZN( u0_u4_u5_n164 ) );
  AOI21_X1 u0_u4_u5_U57 (.ZN( u0_u4_u5_n110 ) , .B1( u0_u4_u5_n122 ) , .B2( u0_u4_u5_n139 ) , .A( u0_u4_u5_n153 ) );
  INV_X1 u0_u4_u5_U58 (.A( u0_u4_u5_n153 ) , .ZN( u0_u4_u5_n176 ) );
  INV_X1 u0_u4_u5_U59 (.A( u0_u4_u5_n126 ) , .ZN( u0_u4_u5_n173 ) );
  AOI222_X1 u0_u4_u5_U6 (.ZN( u0_u4_u5_n113 ) , .A1( u0_u4_u5_n131 ) , .C1( u0_u4_u5_n148 ) , .B2( u0_u4_u5_n174 ) , .C2( u0_u4_u5_n178 ) , .A2( u0_u4_u5_n179 ) , .B1( u0_u4_u5_n99 ) );
  AND2_X1 u0_u4_u5_U60 (.A2( u0_u4_u5_n104 ) , .A1( u0_u4_u5_n107 ) , .ZN( u0_u4_u5_n147 ) );
  AND2_X1 u0_u4_u5_U61 (.A2( u0_u4_u5_n104 ) , .A1( u0_u4_u5_n108 ) , .ZN( u0_u4_u5_n148 ) );
  NAND2_X1 u0_u4_u5_U62 (.A1( u0_u4_u5_n105 ) , .A2( u0_u4_u5_n106 ) , .ZN( u0_u4_u5_n158 ) );
  NAND2_X1 u0_u4_u5_U63 (.A2( u0_u4_u5_n108 ) , .A1( u0_u4_u5_n109 ) , .ZN( u0_u4_u5_n139 ) );
  NAND2_X1 u0_u4_u5_U64 (.A1( u0_u4_u5_n106 ) , .A2( u0_u4_u5_n108 ) , .ZN( u0_u4_u5_n119 ) );
  NAND2_X1 u0_u4_u5_U65 (.A2( u0_u4_u5_n103 ) , .A1( u0_u4_u5_n105 ) , .ZN( u0_u4_u5_n140 ) );
  NAND2_X1 u0_u4_u5_U66 (.A2( u0_u4_u5_n104 ) , .A1( u0_u4_u5_n105 ) , .ZN( u0_u4_u5_n155 ) );
  NAND2_X1 u0_u4_u5_U67 (.A2( u0_u4_u5_n106 ) , .A1( u0_u4_u5_n107 ) , .ZN( u0_u4_u5_n122 ) );
  NAND2_X1 u0_u4_u5_U68 (.A2( u0_u4_u5_n100 ) , .A1( u0_u4_u5_n106 ) , .ZN( u0_u4_u5_n115 ) );
  NAND2_X1 u0_u4_u5_U69 (.A2( u0_u4_u5_n100 ) , .A1( u0_u4_u5_n103 ) , .ZN( u0_u4_u5_n161 ) );
  INV_X1 u0_u4_u5_U7 (.A( u0_u4_u5_n135 ) , .ZN( u0_u4_u5_n178 ) );
  NAND2_X1 u0_u4_u5_U70 (.A1( u0_u4_u5_n105 ) , .A2( u0_u4_u5_n109 ) , .ZN( u0_u4_u5_n154 ) );
  INV_X1 u0_u4_u5_U71 (.A( u0_u4_u5_n146 ) , .ZN( u0_u4_u5_n172 ) );
  NAND2_X1 u0_u4_u5_U72 (.A1( u0_u4_u5_n103 ) , .A2( u0_u4_u5_n108 ) , .ZN( u0_u4_u5_n123 ) );
  NAND2_X1 u0_u4_u5_U73 (.A2( u0_u4_u5_n103 ) , .A1( u0_u4_u5_n107 ) , .ZN( u0_u4_u5_n151 ) );
  NAND2_X1 u0_u4_u5_U74 (.A2( u0_u4_u5_n107 ) , .A1( u0_u4_u5_n109 ) , .ZN( u0_u4_u5_n120 ) );
  NAND2_X1 u0_u4_u5_U75 (.A2( u0_u4_u5_n100 ) , .A1( u0_u4_u5_n109 ) , .ZN( u0_u4_u5_n157 ) );
  AND2_X1 u0_u4_u5_U76 (.A2( u0_u4_u5_n100 ) , .A1( u0_u4_u5_n104 ) , .ZN( u0_u4_u5_n131 ) );
  NOR2_X1 u0_u4_u5_U77 (.A2( u0_u4_X_34 ) , .A1( u0_u4_X_35 ) , .ZN( u0_u4_u5_n145 ) );
  NOR2_X1 u0_u4_u5_U78 (.A2( u0_u4_X_34 ) , .ZN( u0_u4_u5_n146 ) , .A1( u0_u4_u5_n171 ) );
  NOR2_X1 u0_u4_u5_U79 (.A2( u0_u4_X_31 ) , .A1( u0_u4_X_32 ) , .ZN( u0_u4_u5_n103 ) );
  OAI22_X1 u0_u4_u5_U8 (.B2( u0_u4_u5_n149 ) , .B1( u0_u4_u5_n150 ) , .A2( u0_u4_u5_n151 ) , .A1( u0_u4_u5_n152 ) , .ZN( u0_u4_u5_n165 ) );
  NOR2_X1 u0_u4_u5_U80 (.A2( u0_u4_X_36 ) , .ZN( u0_u4_u5_n105 ) , .A1( u0_u4_u5_n180 ) );
  NOR2_X1 u0_u4_u5_U81 (.A2( u0_u4_X_33 ) , .ZN( u0_u4_u5_n108 ) , .A1( u0_u4_u5_n170 ) );
  NOR2_X1 u0_u4_u5_U82 (.A2( u0_u4_X_33 ) , .A1( u0_u4_X_36 ) , .ZN( u0_u4_u5_n107 ) );
  NOR2_X1 u0_u4_u5_U83 (.A2( u0_u4_X_31 ) , .ZN( u0_u4_u5_n104 ) , .A1( u0_u4_u5_n181 ) );
  NAND2_X1 u0_u4_u5_U84 (.A2( u0_u4_X_34 ) , .A1( u0_u4_X_35 ) , .ZN( u0_u4_u5_n153 ) );
  NAND2_X1 u0_u4_u5_U85 (.A1( u0_u4_X_34 ) , .ZN( u0_u4_u5_n126 ) , .A2( u0_u4_u5_n171 ) );
  AND2_X1 u0_u4_u5_U86 (.A1( u0_u4_X_31 ) , .A2( u0_u4_X_32 ) , .ZN( u0_u4_u5_n106 ) );
  AND2_X1 u0_u4_u5_U87 (.A1( u0_u4_X_31 ) , .ZN( u0_u4_u5_n109 ) , .A2( u0_u4_u5_n181 ) );
  INV_X1 u0_u4_u5_U88 (.A( u0_u4_X_33 ) , .ZN( u0_u4_u5_n180 ) );
  INV_X1 u0_u4_u5_U89 (.A( u0_u4_X_35 ) , .ZN( u0_u4_u5_n171 ) );
  NOR3_X1 u0_u4_u5_U9 (.A2( u0_u4_u5_n147 ) , .A1( u0_u4_u5_n148 ) , .ZN( u0_u4_u5_n149 ) , .A3( u0_u4_u5_n194 ) );
  INV_X1 u0_u4_u5_U90 (.A( u0_u4_X_36 ) , .ZN( u0_u4_u5_n170 ) );
  INV_X1 u0_u4_u5_U91 (.A( u0_u4_X_32 ) , .ZN( u0_u4_u5_n181 ) );
  NAND4_X1 u0_u4_u5_U92 (.ZN( u0_out4_29 ) , .A4( u0_u4_u5_n129 ) , .A3( u0_u4_u5_n130 ) , .A2( u0_u4_u5_n168 ) , .A1( u0_u4_u5_n196 ) );
  AOI221_X1 u0_u4_u5_U93 (.A( u0_u4_u5_n128 ) , .ZN( u0_u4_u5_n129 ) , .C2( u0_u4_u5_n132 ) , .B2( u0_u4_u5_n159 ) , .B1( u0_u4_u5_n176 ) , .C1( u0_u4_u5_n184 ) );
  AOI222_X1 u0_u4_u5_U94 (.ZN( u0_u4_u5_n130 ) , .A2( u0_u4_u5_n146 ) , .B1( u0_u4_u5_n147 ) , .C2( u0_u4_u5_n175 ) , .B2( u0_u4_u5_n179 ) , .A1( u0_u4_u5_n188 ) , .C1( u0_u4_u5_n194 ) );
  NAND4_X1 u0_u4_u5_U95 (.ZN( u0_out4_19 ) , .A4( u0_u4_u5_n166 ) , .A3( u0_u4_u5_n167 ) , .A2( u0_u4_u5_n168 ) , .A1( u0_u4_u5_n169 ) );
  AOI22_X1 u0_u4_u5_U96 (.B2( u0_u4_u5_n145 ) , .A2( u0_u4_u5_n146 ) , .ZN( u0_u4_u5_n167 ) , .B1( u0_u4_u5_n182 ) , .A1( u0_u4_u5_n189 ) );
  NOR4_X1 u0_u4_u5_U97 (.A4( u0_u4_u5_n162 ) , .A3( u0_u4_u5_n163 ) , .A2( u0_u4_u5_n164 ) , .A1( u0_u4_u5_n165 ) , .ZN( u0_u4_u5_n166 ) );
  NAND4_X1 u0_u4_u5_U98 (.ZN( u0_out4_11 ) , .A4( u0_u4_u5_n143 ) , .A3( u0_u4_u5_n144 ) , .A2( u0_u4_u5_n169 ) , .A1( u0_u4_u5_n196 ) );
  AOI22_X1 u0_u4_u5_U99 (.A2( u0_u4_u5_n132 ) , .ZN( u0_u4_u5_n144 ) , .B2( u0_u4_u5_n145 ) , .B1( u0_u4_u5_n184 ) , .A1( u0_u4_u5_n194 ) );
  OAI21_X1 u0_u4_u7_U10 (.A( u0_u4_u7_n161 ) , .B1( u0_u4_u7_n168 ) , .B2( u0_u4_u7_n173 ) , .ZN( u0_u4_u7_n91 ) );
  AOI211_X1 u0_u4_u7_U11 (.A( u0_u4_u7_n117 ) , .ZN( u0_u4_u7_n118 ) , .C2( u0_u4_u7_n126 ) , .C1( u0_u4_u7_n177 ) , .B( u0_u4_u7_n180 ) );
  OAI22_X1 u0_u4_u7_U12 (.B1( u0_u4_u7_n115 ) , .ZN( u0_u4_u7_n117 ) , .A2( u0_u4_u7_n133 ) , .A1( u0_u4_u7_n137 ) , .B2( u0_u4_u7_n162 ) );
  INV_X1 u0_u4_u7_U13 (.A( u0_u4_u7_n116 ) , .ZN( u0_u4_u7_n180 ) );
  NOR3_X1 u0_u4_u7_U14 (.ZN( u0_u4_u7_n115 ) , .A3( u0_u4_u7_n145 ) , .A2( u0_u4_u7_n168 ) , .A1( u0_u4_u7_n169 ) );
  INV_X1 u0_u4_u7_U15 (.A( u0_u4_u7_n133 ) , .ZN( u0_u4_u7_n176 ) );
  NOR3_X1 u0_u4_u7_U16 (.A2( u0_u4_u7_n134 ) , .A1( u0_u4_u7_n135 ) , .ZN( u0_u4_u7_n136 ) , .A3( u0_u4_u7_n171 ) );
  NOR2_X1 u0_u4_u7_U17 (.A1( u0_u4_u7_n130 ) , .A2( u0_u4_u7_n134 ) , .ZN( u0_u4_u7_n153 ) );
  AOI21_X1 u0_u4_u7_U18 (.ZN( u0_u4_u7_n104 ) , .B2( u0_u4_u7_n112 ) , .B1( u0_u4_u7_n127 ) , .A( u0_u4_u7_n164 ) );
  AOI21_X1 u0_u4_u7_U19 (.ZN( u0_u4_u7_n106 ) , .B1( u0_u4_u7_n133 ) , .B2( u0_u4_u7_n146 ) , .A( u0_u4_u7_n162 ) );
  AOI21_X1 u0_u4_u7_U20 (.A( u0_u4_u7_n101 ) , .ZN( u0_u4_u7_n107 ) , .B2( u0_u4_u7_n128 ) , .B1( u0_u4_u7_n175 ) );
  INV_X1 u0_u4_u7_U21 (.A( u0_u4_u7_n101 ) , .ZN( u0_u4_u7_n165 ) );
  NOR2_X1 u0_u4_u7_U22 (.ZN( u0_u4_u7_n111 ) , .A2( u0_u4_u7_n134 ) , .A1( u0_u4_u7_n169 ) );
  INV_X1 u0_u4_u7_U23 (.A( u0_u4_u7_n138 ) , .ZN( u0_u4_u7_n171 ) );
  INV_X1 u0_u4_u7_U24 (.A( u0_u4_u7_n131 ) , .ZN( u0_u4_u7_n177 ) );
  INV_X1 u0_u4_u7_U25 (.A( u0_u4_u7_n110 ) , .ZN( u0_u4_u7_n174 ) );
  NAND2_X1 u0_u4_u7_U26 (.A1( u0_u4_u7_n129 ) , .A2( u0_u4_u7_n132 ) , .ZN( u0_u4_u7_n149 ) );
  NAND2_X1 u0_u4_u7_U27 (.A1( u0_u4_u7_n113 ) , .A2( u0_u4_u7_n124 ) , .ZN( u0_u4_u7_n130 ) );
  INV_X1 u0_u4_u7_U28 (.A( u0_u4_u7_n112 ) , .ZN( u0_u4_u7_n173 ) );
  INV_X1 u0_u4_u7_U29 (.A( u0_u4_u7_n128 ) , .ZN( u0_u4_u7_n168 ) );
  OAI21_X1 u0_u4_u7_U3 (.ZN( u0_u4_u7_n159 ) , .A( u0_u4_u7_n165 ) , .B2( u0_u4_u7_n171 ) , .B1( u0_u4_u7_n174 ) );
  INV_X1 u0_u4_u7_U30 (.A( u0_u4_u7_n148 ) , .ZN( u0_u4_u7_n169 ) );
  INV_X1 u0_u4_u7_U31 (.A( u0_u4_u7_n127 ) , .ZN( u0_u4_u7_n179 ) );
  NOR2_X1 u0_u4_u7_U32 (.ZN( u0_u4_u7_n101 ) , .A2( u0_u4_u7_n150 ) , .A1( u0_u4_u7_n156 ) );
  AOI211_X1 u0_u4_u7_U33 (.B( u0_u4_u7_n139 ) , .A( u0_u4_u7_n140 ) , .C2( u0_u4_u7_n141 ) , .ZN( u0_u4_u7_n142 ) , .C1( u0_u4_u7_n156 ) );
  AOI21_X1 u0_u4_u7_U34 (.A( u0_u4_u7_n137 ) , .B1( u0_u4_u7_n138 ) , .ZN( u0_u4_u7_n139 ) , .B2( u0_u4_u7_n146 ) );
  NAND4_X1 u0_u4_u7_U35 (.A3( u0_u4_u7_n127 ) , .A2( u0_u4_u7_n128 ) , .A1( u0_u4_u7_n129 ) , .ZN( u0_u4_u7_n141 ) , .A4( u0_u4_u7_n147 ) );
  OAI22_X1 u0_u4_u7_U36 (.B1( u0_u4_u7_n136 ) , .ZN( u0_u4_u7_n140 ) , .A1( u0_u4_u7_n153 ) , .B2( u0_u4_u7_n162 ) , .A2( u0_u4_u7_n164 ) );
  INV_X1 u0_u4_u7_U37 (.A( u0_u4_u7_n125 ) , .ZN( u0_u4_u7_n161 ) );
  AOI21_X1 u0_u4_u7_U38 (.ZN( u0_u4_u7_n123 ) , .B1( u0_u4_u7_n165 ) , .B2( u0_u4_u7_n177 ) , .A( u0_u4_u7_n97 ) );
  AOI21_X1 u0_u4_u7_U39 (.B2( u0_u4_u7_n113 ) , .B1( u0_u4_u7_n124 ) , .A( u0_u4_u7_n125 ) , .ZN( u0_u4_u7_n97 ) );
  INV_X1 u0_u4_u7_U4 (.A( u0_u4_u7_n149 ) , .ZN( u0_u4_u7_n175 ) );
  INV_X1 u0_u4_u7_U40 (.A( u0_u4_u7_n152 ) , .ZN( u0_u4_u7_n162 ) );
  AOI22_X1 u0_u4_u7_U41 (.A2( u0_u4_u7_n114 ) , .ZN( u0_u4_u7_n119 ) , .B1( u0_u4_u7_n130 ) , .A1( u0_u4_u7_n156 ) , .B2( u0_u4_u7_n165 ) );
  NAND2_X1 u0_u4_u7_U42 (.A2( u0_u4_u7_n112 ) , .ZN( u0_u4_u7_n114 ) , .A1( u0_u4_u7_n175 ) );
  NOR2_X1 u0_u4_u7_U43 (.ZN( u0_u4_u7_n137 ) , .A1( u0_u4_u7_n150 ) , .A2( u0_u4_u7_n161 ) );
  AND2_X1 u0_u4_u7_U44 (.ZN( u0_u4_u7_n145 ) , .A2( u0_u4_u7_n98 ) , .A1( u0_u4_u7_n99 ) );
  AOI21_X1 u0_u4_u7_U45 (.ZN( u0_u4_u7_n105 ) , .B2( u0_u4_u7_n110 ) , .A( u0_u4_u7_n125 ) , .B1( u0_u4_u7_n147 ) );
  NAND2_X1 u0_u4_u7_U46 (.ZN( u0_u4_u7_n146 ) , .A1( u0_u4_u7_n95 ) , .A2( u0_u4_u7_n98 ) );
  NAND2_X1 u0_u4_u7_U47 (.A2( u0_u4_u7_n103 ) , .ZN( u0_u4_u7_n147 ) , .A1( u0_u4_u7_n93 ) );
  NAND2_X1 u0_u4_u7_U48 (.A1( u0_u4_u7_n103 ) , .ZN( u0_u4_u7_n127 ) , .A2( u0_u4_u7_n99 ) );
  NAND2_X1 u0_u4_u7_U49 (.A2( u0_u4_u7_n102 ) , .A1( u0_u4_u7_n103 ) , .ZN( u0_u4_u7_n133 ) );
  INV_X1 u0_u4_u7_U5 (.A( u0_u4_u7_n154 ) , .ZN( u0_u4_u7_n178 ) );
  OR2_X1 u0_u4_u7_U50 (.ZN( u0_u4_u7_n126 ) , .A2( u0_u4_u7_n152 ) , .A1( u0_u4_u7_n156 ) );
  NAND2_X1 u0_u4_u7_U51 (.ZN( u0_u4_u7_n112 ) , .A2( u0_u4_u7_n96 ) , .A1( u0_u4_u7_n99 ) );
  NAND2_X1 u0_u4_u7_U52 (.A2( u0_u4_u7_n102 ) , .ZN( u0_u4_u7_n128 ) , .A1( u0_u4_u7_n98 ) );
  NAND2_X1 u0_u4_u7_U53 (.A1( u0_u4_u7_n100 ) , .ZN( u0_u4_u7_n113 ) , .A2( u0_u4_u7_n93 ) );
  NAND2_X1 u0_u4_u7_U54 (.ZN( u0_u4_u7_n110 ) , .A1( u0_u4_u7_n95 ) , .A2( u0_u4_u7_n96 ) );
  INV_X1 u0_u4_u7_U55 (.A( u0_u4_u7_n150 ) , .ZN( u0_u4_u7_n164 ) );
  AND2_X1 u0_u4_u7_U56 (.ZN( u0_u4_u7_n134 ) , .A1( u0_u4_u7_n93 ) , .A2( u0_u4_u7_n98 ) );
  NAND2_X1 u0_u4_u7_U57 (.A2( u0_u4_u7_n102 ) , .ZN( u0_u4_u7_n124 ) , .A1( u0_u4_u7_n96 ) );
  NAND2_X1 u0_u4_u7_U58 (.A1( u0_u4_u7_n100 ) , .A2( u0_u4_u7_n102 ) , .ZN( u0_u4_u7_n129 ) );
  NAND2_X1 u0_u4_u7_U59 (.A2( u0_u4_u7_n103 ) , .ZN( u0_u4_u7_n131 ) , .A1( u0_u4_u7_n95 ) );
  AOI211_X1 u0_u4_u7_U6 (.ZN( u0_u4_u7_n116 ) , .A( u0_u4_u7_n155 ) , .C1( u0_u4_u7_n161 ) , .C2( u0_u4_u7_n171 ) , .B( u0_u4_u7_n94 ) );
  NAND2_X1 u0_u4_u7_U60 (.A1( u0_u4_u7_n100 ) , .ZN( u0_u4_u7_n138 ) , .A2( u0_u4_u7_n99 ) );
  NAND2_X1 u0_u4_u7_U61 (.ZN( u0_u4_u7_n132 ) , .A1( u0_u4_u7_n93 ) , .A2( u0_u4_u7_n96 ) );
  NAND2_X1 u0_u4_u7_U62 (.A1( u0_u4_u7_n100 ) , .ZN( u0_u4_u7_n148 ) , .A2( u0_u4_u7_n95 ) );
  AOI211_X1 u0_u4_u7_U63 (.B( u0_u4_u7_n154 ) , .A( u0_u4_u7_n155 ) , .C1( u0_u4_u7_n156 ) , .ZN( u0_u4_u7_n157 ) , .C2( u0_u4_u7_n172 ) );
  INV_X1 u0_u4_u7_U64 (.A( u0_u4_u7_n153 ) , .ZN( u0_u4_u7_n172 ) );
  NOR2_X1 u0_u4_u7_U65 (.A2( u0_u4_X_47 ) , .ZN( u0_u4_u7_n150 ) , .A1( u0_u4_u7_n163 ) );
  NOR2_X1 u0_u4_u7_U66 (.A2( u0_u4_X_43 ) , .A1( u0_u4_X_44 ) , .ZN( u0_u4_u7_n103 ) );
  NOR2_X1 u0_u4_u7_U67 (.A2( u0_u4_X_48 ) , .A1( u0_u4_u7_n166 ) , .ZN( u0_u4_u7_n95 ) );
  NOR2_X1 u0_u4_u7_U68 (.A2( u0_u4_X_45 ) , .A1( u0_u4_X_48 ) , .ZN( u0_u4_u7_n99 ) );
  NOR2_X1 u0_u4_u7_U69 (.A2( u0_u4_X_44 ) , .A1( u0_u4_u7_n167 ) , .ZN( u0_u4_u7_n98 ) );
  OAI222_X1 u0_u4_u7_U7 (.C2( u0_u4_u7_n101 ) , .B2( u0_u4_u7_n111 ) , .A1( u0_u4_u7_n113 ) , .C1( u0_u4_u7_n146 ) , .A2( u0_u4_u7_n162 ) , .B1( u0_u4_u7_n164 ) , .ZN( u0_u4_u7_n94 ) );
  NOR2_X1 u0_u4_u7_U70 (.A2( u0_u4_X_46 ) , .A1( u0_u4_X_47 ) , .ZN( u0_u4_u7_n152 ) );
  NAND2_X1 u0_u4_u7_U71 (.A2( u0_u4_X_46 ) , .A1( u0_u4_X_47 ) , .ZN( u0_u4_u7_n125 ) );
  AND2_X1 u0_u4_u7_U72 (.A1( u0_u4_X_47 ) , .ZN( u0_u4_u7_n156 ) , .A2( u0_u4_u7_n163 ) );
  AND2_X1 u0_u4_u7_U73 (.A2( u0_u4_X_45 ) , .A1( u0_u4_X_48 ) , .ZN( u0_u4_u7_n102 ) );
  AND2_X1 u0_u4_u7_U74 (.A2( u0_u4_X_43 ) , .A1( u0_u4_X_44 ) , .ZN( u0_u4_u7_n96 ) );
  AND2_X1 u0_u4_u7_U75 (.A1( u0_u4_X_44 ) , .ZN( u0_u4_u7_n100 ) , .A2( u0_u4_u7_n167 ) );
  AND2_X1 u0_u4_u7_U76 (.A1( u0_u4_X_48 ) , .A2( u0_u4_u7_n166 ) , .ZN( u0_u4_u7_n93 ) );
  INV_X1 u0_u4_u7_U77 (.A( u0_u4_X_46 ) , .ZN( u0_u4_u7_n163 ) );
  INV_X1 u0_u4_u7_U78 (.A( u0_u4_X_43 ) , .ZN( u0_u4_u7_n167 ) );
  INV_X1 u0_u4_u7_U79 (.A( u0_u4_X_45 ) , .ZN( u0_u4_u7_n166 ) );
  OAI221_X1 u0_u4_u7_U8 (.C1( u0_u4_u7_n101 ) , .C2( u0_u4_u7_n147 ) , .ZN( u0_u4_u7_n155 ) , .B2( u0_u4_u7_n162 ) , .A( u0_u4_u7_n91 ) , .B1( u0_u4_u7_n92 ) );
  NAND4_X1 u0_u4_u7_U80 (.ZN( u0_out4_5 ) , .A4( u0_u4_u7_n108 ) , .A3( u0_u4_u7_n109 ) , .A1( u0_u4_u7_n116 ) , .A2( u0_u4_u7_n123 ) );
  AOI22_X1 u0_u4_u7_U81 (.ZN( u0_u4_u7_n109 ) , .A2( u0_u4_u7_n126 ) , .B2( u0_u4_u7_n145 ) , .B1( u0_u4_u7_n156 ) , .A1( u0_u4_u7_n171 ) );
  NOR4_X1 u0_u4_u7_U82 (.A4( u0_u4_u7_n104 ) , .A3( u0_u4_u7_n105 ) , .A2( u0_u4_u7_n106 ) , .A1( u0_u4_u7_n107 ) , .ZN( u0_u4_u7_n108 ) );
  NAND4_X1 u0_u4_u7_U83 (.ZN( u0_out4_27 ) , .A4( u0_u4_u7_n118 ) , .A3( u0_u4_u7_n119 ) , .A2( u0_u4_u7_n120 ) , .A1( u0_u4_u7_n121 ) );
  OAI21_X1 u0_u4_u7_U84 (.ZN( u0_u4_u7_n121 ) , .B2( u0_u4_u7_n145 ) , .A( u0_u4_u7_n150 ) , .B1( u0_u4_u7_n174 ) );
  OAI21_X1 u0_u4_u7_U85 (.ZN( u0_u4_u7_n120 ) , .A( u0_u4_u7_n161 ) , .B2( u0_u4_u7_n170 ) , .B1( u0_u4_u7_n179 ) );
  NAND4_X1 u0_u4_u7_U86 (.ZN( u0_out4_21 ) , .A4( u0_u4_u7_n157 ) , .A3( u0_u4_u7_n158 ) , .A2( u0_u4_u7_n159 ) , .A1( u0_u4_u7_n160 ) );
  OAI21_X1 u0_u4_u7_U87 (.B1( u0_u4_u7_n145 ) , .ZN( u0_u4_u7_n160 ) , .A( u0_u4_u7_n161 ) , .B2( u0_u4_u7_n177 ) );
  AOI22_X1 u0_u4_u7_U88 (.B2( u0_u4_u7_n149 ) , .B1( u0_u4_u7_n150 ) , .A2( u0_u4_u7_n151 ) , .A1( u0_u4_u7_n152 ) , .ZN( u0_u4_u7_n158 ) );
  NAND4_X1 u0_u4_u7_U89 (.ZN( u0_out4_15 ) , .A4( u0_u4_u7_n142 ) , .A3( u0_u4_u7_n143 ) , .A2( u0_u4_u7_n144 ) , .A1( u0_u4_u7_n178 ) );
  AND3_X1 u0_u4_u7_U9 (.A3( u0_u4_u7_n110 ) , .A2( u0_u4_u7_n127 ) , .A1( u0_u4_u7_n132 ) , .ZN( u0_u4_u7_n92 ) );
  OR2_X1 u0_u4_u7_U90 (.A2( u0_u4_u7_n125 ) , .A1( u0_u4_u7_n129 ) , .ZN( u0_u4_u7_n144 ) );
  AOI22_X1 u0_u4_u7_U91 (.A2( u0_u4_u7_n126 ) , .ZN( u0_u4_u7_n143 ) , .B2( u0_u4_u7_n165 ) , .B1( u0_u4_u7_n173 ) , .A1( u0_u4_u7_n174 ) );
  OAI211_X1 u0_u4_u7_U92 (.B( u0_u4_u7_n122 ) , .A( u0_u4_u7_n123 ) , .C2( u0_u4_u7_n124 ) , .ZN( u0_u4_u7_n154 ) , .C1( u0_u4_u7_n162 ) );
  AOI222_X1 u0_u4_u7_U93 (.ZN( u0_u4_u7_n122 ) , .C2( u0_u4_u7_n126 ) , .C1( u0_u4_u7_n145 ) , .B1( u0_u4_u7_n161 ) , .A2( u0_u4_u7_n165 ) , .B2( u0_u4_u7_n170 ) , .A1( u0_u4_u7_n176 ) );
  INV_X1 u0_u4_u7_U94 (.A( u0_u4_u7_n111 ) , .ZN( u0_u4_u7_n170 ) );
  NAND3_X1 u0_u4_u7_U95 (.A3( u0_u4_u7_n146 ) , .A2( u0_u4_u7_n147 ) , .A1( u0_u4_u7_n148 ) , .ZN( u0_u4_u7_n151 ) );
  NAND3_X1 u0_u4_u7_U96 (.A3( u0_u4_u7_n131 ) , .A2( u0_u4_u7_n132 ) , .A1( u0_u4_u7_n133 ) , .ZN( u0_u4_u7_n135 ) );
  XOR2_X1 u0_u6_U16 (.B( u0_K7_3 ) , .A( u0_R5_2 ) , .Z( u0_u6_X_3 ) );
  XOR2_X1 u0_u6_U2 (.B( u0_K7_8 ) , .A( u0_R5_5 ) , .Z( u0_u6_X_8 ) );
  XOR2_X1 u0_u6_U20 (.B( u0_K7_36 ) , .A( u0_R5_25 ) , .Z( u0_u6_X_36 ) );
  XOR2_X1 u0_u6_U3 (.B( u0_K7_7 ) , .A( u0_R5_4 ) , .Z( u0_u6_X_7 ) );
  XOR2_X1 u0_u6_U37 (.B( u0_K7_20 ) , .A( u0_R5_13 ) , .Z( u0_u6_X_20 ) );
  XOR2_X1 u0_u6_U38 (.B( u0_K7_1 ) , .A( u0_R5_32 ) , .Z( u0_u6_X_1 ) );
  XOR2_X1 u0_u6_U39 (.B( u0_K7_19 ) , .A( u0_R5_12 ) , .Z( u0_u6_X_19 ) );
  XOR2_X1 u0_u6_U4 (.B( u0_K7_6 ) , .A( u0_R5_5 ) , .Z( u0_u6_X_6 ) );
  XOR2_X1 u0_u6_U40 (.B( u0_K7_18 ) , .A( u0_R5_13 ) , .Z( u0_u6_X_18 ) );
  XOR2_X1 u0_u6_U41 (.B( u0_K7_17 ) , .A( u0_R5_12 ) , .Z( u0_u6_X_17 ) );
  XOR2_X1 u0_u6_U44 (.B( u0_K7_14 ) , .A( u0_R5_9 ) , .Z( u0_u6_X_14 ) );
  XOR2_X1 u0_u6_U45 (.B( u0_K7_13 ) , .A( u0_R5_8 ) , .Z( u0_u6_X_13 ) );
  XOR2_X1 u0_u6_U46 (.B( u0_K7_12 ) , .A( u0_R5_9 ) , .Z( u0_u6_X_12 ) );
  XOR2_X1 u0_u6_U47 (.B( u0_K7_11 ) , .A( u0_R5_8 ) , .Z( u0_u6_X_11 ) );
  XOR2_X1 u0_u6_U48 (.B( u0_K7_10 ) , .A( u0_R5_7 ) , .Z( u0_u6_X_10 ) );
  XOR2_X1 u0_u6_U5 (.B( u0_K7_5 ) , .A( u0_R5_4 ) , .Z( u0_u6_X_5 ) );
  XOR2_X1 u0_u6_U6 (.B( u0_K7_4 ) , .A( u0_R5_3 ) , .Z( u0_u6_X_4 ) );
  NAND2_X1 u0_u6_u0_U10 (.ZN( u0_u6_u0_n113 ) , .A1( u0_u6_u0_n139 ) , .A2( u0_u6_u0_n149 ) );
  AND2_X1 u0_u6_u0_U11 (.A1( u0_u6_u0_n131 ) , .ZN( u0_u6_u0_n141 ) , .A2( u0_u6_u0_n150 ) );
  AND2_X1 u0_u6_u0_U12 (.ZN( u0_u6_u0_n107 ) , .A1( u0_u6_u0_n130 ) , .A2( u0_u6_u0_n140 ) );
  AND2_X1 u0_u6_u0_U13 (.A2( u0_u6_u0_n129 ) , .A1( u0_u6_u0_n130 ) , .ZN( u0_u6_u0_n151 ) );
  AND2_X1 u0_u6_u0_U14 (.A1( u0_u6_u0_n108 ) , .A2( u0_u6_u0_n125 ) , .ZN( u0_u6_u0_n145 ) );
  INV_X1 u0_u6_u0_U15 (.A( u0_u6_u0_n143 ) , .ZN( u0_u6_u0_n173 ) );
  NOR2_X1 u0_u6_u0_U16 (.A2( u0_u6_u0_n136 ) , .ZN( u0_u6_u0_n147 ) , .A1( u0_u6_u0_n160 ) );
  AOI21_X1 u0_u6_u0_U17 (.B1( u0_u6_u0_n103 ) , .ZN( u0_u6_u0_n132 ) , .A( u0_u6_u0_n165 ) , .B2( u0_u6_u0_n93 ) );
  OAI221_X1 u0_u6_u0_U18 (.C1( u0_u6_u0_n121 ) , .ZN( u0_u6_u0_n122 ) , .B2( u0_u6_u0_n127 ) , .A( u0_u6_u0_n143 ) , .B1( u0_u6_u0_n144 ) , .C2( u0_u6_u0_n147 ) );
  OAI22_X1 u0_u6_u0_U19 (.B1( u0_u6_u0_n125 ) , .ZN( u0_u6_u0_n126 ) , .A1( u0_u6_u0_n138 ) , .A2( u0_u6_u0_n146 ) , .B2( u0_u6_u0_n147 ) );
  OAI22_X1 u0_u6_u0_U20 (.B1( u0_u6_u0_n131 ) , .A1( u0_u6_u0_n144 ) , .B2( u0_u6_u0_n147 ) , .A2( u0_u6_u0_n90 ) , .ZN( u0_u6_u0_n91 ) );
  AND3_X1 u0_u6_u0_U21 (.A3( u0_u6_u0_n121 ) , .A2( u0_u6_u0_n125 ) , .A1( u0_u6_u0_n148 ) , .ZN( u0_u6_u0_n90 ) );
  NOR2_X1 u0_u6_u0_U22 (.A1( u0_u6_u0_n163 ) , .A2( u0_u6_u0_n164 ) , .ZN( u0_u6_u0_n95 ) );
  NOR2_X1 u0_u6_u0_U23 (.A1( u0_u6_u0_n120 ) , .ZN( u0_u6_u0_n143 ) , .A2( u0_u6_u0_n167 ) );
  OAI221_X1 u0_u6_u0_U24 (.C1( u0_u6_u0_n112 ) , .ZN( u0_u6_u0_n120 ) , .B1( u0_u6_u0_n138 ) , .B2( u0_u6_u0_n141 ) , .C2( u0_u6_u0_n147 ) , .A( u0_u6_u0_n172 ) );
  AOI211_X1 u0_u6_u0_U25 (.B( u0_u6_u0_n115 ) , .A( u0_u6_u0_n116 ) , .C2( u0_u6_u0_n117 ) , .C1( u0_u6_u0_n118 ) , .ZN( u0_u6_u0_n119 ) );
  AOI22_X1 u0_u6_u0_U26 (.B2( u0_u6_u0_n109 ) , .A2( u0_u6_u0_n110 ) , .ZN( u0_u6_u0_n111 ) , .B1( u0_u6_u0_n118 ) , .A1( u0_u6_u0_n160 ) );
  NAND2_X1 u0_u6_u0_U27 (.A1( u0_u6_u0_n100 ) , .A2( u0_u6_u0_n103 ) , .ZN( u0_u6_u0_n125 ) );
  INV_X1 u0_u6_u0_U28 (.A( u0_u6_u0_n136 ) , .ZN( u0_u6_u0_n161 ) );
  INV_X1 u0_u6_u0_U29 (.A( u0_u6_u0_n118 ) , .ZN( u0_u6_u0_n158 ) );
  INV_X1 u0_u6_u0_U3 (.A( u0_u6_u0_n113 ) , .ZN( u0_u6_u0_n166 ) );
  AOI21_X1 u0_u6_u0_U30 (.B1( u0_u6_u0_n127 ) , .B2( u0_u6_u0_n129 ) , .A( u0_u6_u0_n138 ) , .ZN( u0_u6_u0_n96 ) );
  AOI21_X1 u0_u6_u0_U31 (.ZN( u0_u6_u0_n104 ) , .B1( u0_u6_u0_n107 ) , .B2( u0_u6_u0_n141 ) , .A( u0_u6_u0_n144 ) );
  NAND2_X1 u0_u6_u0_U32 (.A2( u0_u6_u0_n102 ) , .A1( u0_u6_u0_n103 ) , .ZN( u0_u6_u0_n149 ) );
  NAND2_X1 u0_u6_u0_U33 (.A2( u0_u6_u0_n100 ) , .ZN( u0_u6_u0_n131 ) , .A1( u0_u6_u0_n92 ) );
  NAND2_X1 u0_u6_u0_U34 (.A2( u0_u6_u0_n102 ) , .ZN( u0_u6_u0_n114 ) , .A1( u0_u6_u0_n92 ) );
  NAND2_X1 u0_u6_u0_U35 (.A1( u0_u6_u0_n101 ) , .A2( u0_u6_u0_n102 ) , .ZN( u0_u6_u0_n150 ) );
  INV_X1 u0_u6_u0_U36 (.A( u0_u6_u0_n138 ) , .ZN( u0_u6_u0_n160 ) );
  NAND2_X1 u0_u6_u0_U37 (.A2( u0_u6_u0_n100 ) , .A1( u0_u6_u0_n101 ) , .ZN( u0_u6_u0_n139 ) );
  NAND2_X1 u0_u6_u0_U38 (.ZN( u0_u6_u0_n112 ) , .A2( u0_u6_u0_n92 ) , .A1( u0_u6_u0_n93 ) );
  NAND2_X1 u0_u6_u0_U39 (.A2( u0_u6_u0_n101 ) , .ZN( u0_u6_u0_n121 ) , .A1( u0_u6_u0_n93 ) );
  AOI21_X1 u0_u6_u0_U4 (.B1( u0_u6_u0_n114 ) , .ZN( u0_u6_u0_n115 ) , .B2( u0_u6_u0_n129 ) , .A( u0_u6_u0_n161 ) );
  INV_X1 u0_u6_u0_U40 (.ZN( u0_u6_u0_n172 ) , .A( u0_u6_u0_n88 ) );
  OAI222_X1 u0_u6_u0_U41 (.C1( u0_u6_u0_n108 ) , .A1( u0_u6_u0_n125 ) , .B2( u0_u6_u0_n128 ) , .B1( u0_u6_u0_n144 ) , .A2( u0_u6_u0_n158 ) , .C2( u0_u6_u0_n161 ) , .ZN( u0_u6_u0_n88 ) );
  OR3_X1 u0_u6_u0_U42 (.A3( u0_u6_u0_n152 ) , .A2( u0_u6_u0_n153 ) , .A1( u0_u6_u0_n154 ) , .ZN( u0_u6_u0_n155 ) );
  AOI21_X1 u0_u6_u0_U43 (.A( u0_u6_u0_n144 ) , .B2( u0_u6_u0_n145 ) , .B1( u0_u6_u0_n146 ) , .ZN( u0_u6_u0_n154 ) );
  AOI21_X1 u0_u6_u0_U44 (.B2( u0_u6_u0_n150 ) , .B1( u0_u6_u0_n151 ) , .ZN( u0_u6_u0_n152 ) , .A( u0_u6_u0_n158 ) );
  AOI21_X1 u0_u6_u0_U45 (.A( u0_u6_u0_n147 ) , .B2( u0_u6_u0_n148 ) , .B1( u0_u6_u0_n149 ) , .ZN( u0_u6_u0_n153 ) );
  INV_X1 u0_u6_u0_U46 (.ZN( u0_u6_u0_n171 ) , .A( u0_u6_u0_n99 ) );
  OAI211_X1 u0_u6_u0_U47 (.C2( u0_u6_u0_n140 ) , .C1( u0_u6_u0_n161 ) , .A( u0_u6_u0_n169 ) , .B( u0_u6_u0_n98 ) , .ZN( u0_u6_u0_n99 ) );
  AOI211_X1 u0_u6_u0_U48 (.C1( u0_u6_u0_n118 ) , .A( u0_u6_u0_n123 ) , .B( u0_u6_u0_n96 ) , .C2( u0_u6_u0_n97 ) , .ZN( u0_u6_u0_n98 ) );
  INV_X1 u0_u6_u0_U49 (.ZN( u0_u6_u0_n169 ) , .A( u0_u6_u0_n91 ) );
  NOR2_X1 u0_u6_u0_U5 (.A1( u0_u6_u0_n108 ) , .ZN( u0_u6_u0_n123 ) , .A2( u0_u6_u0_n158 ) );
  NOR2_X1 u0_u6_u0_U50 (.A2( u0_u6_X_4 ) , .A1( u0_u6_X_5 ) , .ZN( u0_u6_u0_n118 ) );
  NOR2_X1 u0_u6_u0_U51 (.A2( u0_u6_X_1 ) , .ZN( u0_u6_u0_n101 ) , .A1( u0_u6_u0_n163 ) );
  NAND2_X1 u0_u6_u0_U52 (.A2( u0_u6_X_4 ) , .A1( u0_u6_X_5 ) , .ZN( u0_u6_u0_n144 ) );
  NOR2_X1 u0_u6_u0_U53 (.A2( u0_u6_X_5 ) , .ZN( u0_u6_u0_n136 ) , .A1( u0_u6_u0_n159 ) );
  NAND2_X1 u0_u6_u0_U54 (.A1( u0_u6_X_5 ) , .ZN( u0_u6_u0_n138 ) , .A2( u0_u6_u0_n159 ) );
  AND2_X1 u0_u6_u0_U55 (.A2( u0_u6_X_3 ) , .A1( u0_u6_X_6 ) , .ZN( u0_u6_u0_n102 ) );
  INV_X1 u0_u6_u0_U56 (.A( u0_u6_X_4 ) , .ZN( u0_u6_u0_n159 ) );
  INV_X1 u0_u6_u0_U57 (.A( u0_u6_X_1 ) , .ZN( u0_u6_u0_n164 ) );
  INV_X1 u0_u6_u0_U58 (.A( u0_u6_X_3 ) , .ZN( u0_u6_u0_n162 ) );
  INV_X1 u0_u6_u0_U59 (.A( u0_u6_u0_n126 ) , .ZN( u0_u6_u0_n168 ) );
  AOI21_X1 u0_u6_u0_U6 (.B2( u0_u6_u0_n131 ) , .ZN( u0_u6_u0_n134 ) , .B1( u0_u6_u0_n151 ) , .A( u0_u6_u0_n158 ) );
  AOI211_X1 u0_u6_u0_U60 (.B( u0_u6_u0_n133 ) , .A( u0_u6_u0_n134 ) , .C2( u0_u6_u0_n135 ) , .C1( u0_u6_u0_n136 ) , .ZN( u0_u6_u0_n137 ) );
  INV_X1 u0_u6_u0_U61 (.ZN( u0_u6_u0_n174 ) , .A( u0_u6_u0_n89 ) );
  AOI211_X1 u0_u6_u0_U62 (.B( u0_u6_u0_n104 ) , .A( u0_u6_u0_n105 ) , .ZN( u0_u6_u0_n106 ) , .C2( u0_u6_u0_n113 ) , .C1( u0_u6_u0_n160 ) );
  OR4_X1 u0_u6_u0_U63 (.ZN( u0_out6_31 ) , .A4( u0_u6_u0_n155 ) , .A2( u0_u6_u0_n156 ) , .A1( u0_u6_u0_n157 ) , .A3( u0_u6_u0_n173 ) );
  AOI21_X1 u0_u6_u0_U64 (.A( u0_u6_u0_n138 ) , .B2( u0_u6_u0_n139 ) , .B1( u0_u6_u0_n140 ) , .ZN( u0_u6_u0_n157 ) );
  OR4_X1 u0_u6_u0_U65 (.ZN( u0_out6_17 ) , .A4( u0_u6_u0_n122 ) , .A2( u0_u6_u0_n123 ) , .A1( u0_u6_u0_n124 ) , .A3( u0_u6_u0_n170 ) );
  AOI21_X1 u0_u6_u0_U66 (.B2( u0_u6_u0_n107 ) , .ZN( u0_u6_u0_n124 ) , .B1( u0_u6_u0_n128 ) , .A( u0_u6_u0_n161 ) );
  INV_X1 u0_u6_u0_U67 (.A( u0_u6_u0_n111 ) , .ZN( u0_u6_u0_n170 ) );
  AOI21_X1 u0_u6_u0_U68 (.B2( u0_u6_u0_n141 ) , .B1( u0_u6_u0_n142 ) , .ZN( u0_u6_u0_n156 ) , .A( u0_u6_u0_n161 ) );
  AOI21_X1 u0_u6_u0_U69 (.ZN( u0_u6_u0_n116 ) , .B2( u0_u6_u0_n142 ) , .A( u0_u6_u0_n144 ) , .B1( u0_u6_u0_n166 ) );
  OAI21_X1 u0_u6_u0_U7 (.B1( u0_u6_u0_n150 ) , .B2( u0_u6_u0_n158 ) , .A( u0_u6_u0_n172 ) , .ZN( u0_u6_u0_n89 ) );
  NAND2_X1 u0_u6_u0_U70 (.ZN( u0_u6_u0_n148 ) , .A1( u0_u6_u0_n93 ) , .A2( u0_u6_u0_n95 ) );
  NAND2_X1 u0_u6_u0_U71 (.A1( u0_u6_u0_n100 ) , .ZN( u0_u6_u0_n129 ) , .A2( u0_u6_u0_n95 ) );
  NAND2_X1 u0_u6_u0_U72 (.A1( u0_u6_u0_n102 ) , .ZN( u0_u6_u0_n128 ) , .A2( u0_u6_u0_n95 ) );
  INV_X1 u0_u6_u0_U73 (.A( u0_u6_u0_n142 ) , .ZN( u0_u6_u0_n165 ) );
  NOR2_X1 u0_u6_u0_U74 (.A2( u0_u6_X_1 ) , .A1( u0_u6_X_2 ) , .ZN( u0_u6_u0_n92 ) );
  NOR2_X1 u0_u6_u0_U75 (.A2( u0_u6_X_2 ) , .ZN( u0_u6_u0_n103 ) , .A1( u0_u6_u0_n164 ) );
  INV_X1 u0_u6_u0_U76 (.A( u0_u6_X_2 ) , .ZN( u0_u6_u0_n163 ) );
  AOI21_X1 u0_u6_u0_U77 (.B1( u0_u6_u0_n132 ) , .ZN( u0_u6_u0_n133 ) , .A( u0_u6_u0_n144 ) , .B2( u0_u6_u0_n166 ) );
  OAI22_X1 u0_u6_u0_U78 (.ZN( u0_u6_u0_n105 ) , .A2( u0_u6_u0_n132 ) , .B1( u0_u6_u0_n146 ) , .A1( u0_u6_u0_n147 ) , .B2( u0_u6_u0_n161 ) );
  NAND2_X1 u0_u6_u0_U79 (.ZN( u0_u6_u0_n110 ) , .A2( u0_u6_u0_n132 ) , .A1( u0_u6_u0_n145 ) );
  AND2_X1 u0_u6_u0_U8 (.A1( u0_u6_u0_n114 ) , .A2( u0_u6_u0_n121 ) , .ZN( u0_u6_u0_n146 ) );
  INV_X1 u0_u6_u0_U80 (.A( u0_u6_u0_n119 ) , .ZN( u0_u6_u0_n167 ) );
  NAND2_X1 u0_u6_u0_U81 (.A2( u0_u6_u0_n103 ) , .ZN( u0_u6_u0_n140 ) , .A1( u0_u6_u0_n94 ) );
  NAND2_X1 u0_u6_u0_U82 (.A1( u0_u6_u0_n101 ) , .ZN( u0_u6_u0_n130 ) , .A2( u0_u6_u0_n94 ) );
  NAND2_X1 u0_u6_u0_U83 (.ZN( u0_u6_u0_n108 ) , .A1( u0_u6_u0_n92 ) , .A2( u0_u6_u0_n94 ) );
  AND2_X1 u0_u6_u0_U84 (.A1( u0_u6_X_6 ) , .A2( u0_u6_u0_n162 ) , .ZN( u0_u6_u0_n93 ) );
  NAND2_X1 u0_u6_u0_U85 (.ZN( u0_u6_u0_n142 ) , .A1( u0_u6_u0_n94 ) , .A2( u0_u6_u0_n95 ) );
  NOR2_X1 u0_u6_u0_U86 (.A2( u0_u6_X_6 ) , .ZN( u0_u6_u0_n100 ) , .A1( u0_u6_u0_n162 ) );
  NOR2_X1 u0_u6_u0_U87 (.A2( u0_u6_X_3 ) , .A1( u0_u6_X_6 ) , .ZN( u0_u6_u0_n94 ) );
  NAND3_X1 u0_u6_u0_U88 (.ZN( u0_out6_23 ) , .A3( u0_u6_u0_n137 ) , .A1( u0_u6_u0_n168 ) , .A2( u0_u6_u0_n171 ) );
  NAND3_X1 u0_u6_u0_U89 (.A3( u0_u6_u0_n127 ) , .A2( u0_u6_u0_n128 ) , .ZN( u0_u6_u0_n135 ) , .A1( u0_u6_u0_n150 ) );
  AND3_X1 u0_u6_u0_U9 (.A2( u0_u6_u0_n112 ) , .ZN( u0_u6_u0_n127 ) , .A3( u0_u6_u0_n130 ) , .A1( u0_u6_u0_n148 ) );
  NAND3_X1 u0_u6_u0_U90 (.ZN( u0_u6_u0_n117 ) , .A3( u0_u6_u0_n132 ) , .A2( u0_u6_u0_n139 ) , .A1( u0_u6_u0_n148 ) );
  NAND3_X1 u0_u6_u0_U91 (.ZN( u0_u6_u0_n109 ) , .A2( u0_u6_u0_n114 ) , .A3( u0_u6_u0_n140 ) , .A1( u0_u6_u0_n149 ) );
  NAND3_X1 u0_u6_u0_U92 (.ZN( u0_out6_9 ) , .A3( u0_u6_u0_n106 ) , .A2( u0_u6_u0_n171 ) , .A1( u0_u6_u0_n174 ) );
  NAND3_X1 u0_u6_u0_U93 (.A2( u0_u6_u0_n128 ) , .A1( u0_u6_u0_n132 ) , .A3( u0_u6_u0_n146 ) , .ZN( u0_u6_u0_n97 ) );
  AOI21_X1 u0_u6_u1_U10 (.B2( u0_u6_u1_n155 ) , .B1( u0_u6_u1_n156 ) , .ZN( u0_u6_u1_n157 ) , .A( u0_u6_u1_n174 ) );
  NAND3_X1 u0_u6_u1_U100 (.ZN( u0_u6_u1_n113 ) , .A1( u0_u6_u1_n120 ) , .A3( u0_u6_u1_n133 ) , .A2( u0_u6_u1_n155 ) );
  NAND2_X1 u0_u6_u1_U11 (.ZN( u0_u6_u1_n140 ) , .A2( u0_u6_u1_n150 ) , .A1( u0_u6_u1_n155 ) );
  NAND2_X1 u0_u6_u1_U12 (.A1( u0_u6_u1_n131 ) , .ZN( u0_u6_u1_n147 ) , .A2( u0_u6_u1_n153 ) );
  INV_X1 u0_u6_u1_U13 (.A( u0_u6_u1_n139 ) , .ZN( u0_u6_u1_n174 ) );
  OR4_X1 u0_u6_u1_U14 (.A4( u0_u6_u1_n106 ) , .A3( u0_u6_u1_n107 ) , .ZN( u0_u6_u1_n108 ) , .A1( u0_u6_u1_n117 ) , .A2( u0_u6_u1_n184 ) );
  AOI21_X1 u0_u6_u1_U15 (.ZN( u0_u6_u1_n106 ) , .A( u0_u6_u1_n112 ) , .B1( u0_u6_u1_n154 ) , .B2( u0_u6_u1_n156 ) );
  AOI21_X1 u0_u6_u1_U16 (.ZN( u0_u6_u1_n107 ) , .B1( u0_u6_u1_n134 ) , .B2( u0_u6_u1_n149 ) , .A( u0_u6_u1_n174 ) );
  INV_X1 u0_u6_u1_U17 (.A( u0_u6_u1_n101 ) , .ZN( u0_u6_u1_n184 ) );
  INV_X1 u0_u6_u1_U18 (.A( u0_u6_u1_n112 ) , .ZN( u0_u6_u1_n171 ) );
  NAND2_X1 u0_u6_u1_U19 (.ZN( u0_u6_u1_n141 ) , .A1( u0_u6_u1_n153 ) , .A2( u0_u6_u1_n156 ) );
  AND2_X1 u0_u6_u1_U20 (.A1( u0_u6_u1_n123 ) , .ZN( u0_u6_u1_n134 ) , .A2( u0_u6_u1_n161 ) );
  NAND2_X1 u0_u6_u1_U21 (.A2( u0_u6_u1_n115 ) , .A1( u0_u6_u1_n116 ) , .ZN( u0_u6_u1_n148 ) );
  NAND2_X1 u0_u6_u1_U22 (.A2( u0_u6_u1_n133 ) , .A1( u0_u6_u1_n135 ) , .ZN( u0_u6_u1_n159 ) );
  NAND2_X1 u0_u6_u1_U23 (.A2( u0_u6_u1_n115 ) , .A1( u0_u6_u1_n120 ) , .ZN( u0_u6_u1_n132 ) );
  INV_X1 u0_u6_u1_U24 (.A( u0_u6_u1_n154 ) , .ZN( u0_u6_u1_n178 ) );
  AOI22_X1 u0_u6_u1_U25 (.B2( u0_u6_u1_n113 ) , .A2( u0_u6_u1_n114 ) , .ZN( u0_u6_u1_n125 ) , .A1( u0_u6_u1_n171 ) , .B1( u0_u6_u1_n173 ) );
  NAND2_X1 u0_u6_u1_U26 (.ZN( u0_u6_u1_n114 ) , .A1( u0_u6_u1_n134 ) , .A2( u0_u6_u1_n156 ) );
  INV_X1 u0_u6_u1_U27 (.A( u0_u6_u1_n151 ) , .ZN( u0_u6_u1_n183 ) );
  AND2_X1 u0_u6_u1_U28 (.A1( u0_u6_u1_n129 ) , .A2( u0_u6_u1_n133 ) , .ZN( u0_u6_u1_n149 ) );
  INV_X1 u0_u6_u1_U29 (.A( u0_u6_u1_n131 ) , .ZN( u0_u6_u1_n180 ) );
  INV_X1 u0_u6_u1_U3 (.A( u0_u6_u1_n159 ) , .ZN( u0_u6_u1_n182 ) );
  AOI221_X1 u0_u6_u1_U30 (.B1( u0_u6_u1_n140 ) , .ZN( u0_u6_u1_n167 ) , .B2( u0_u6_u1_n172 ) , .C2( u0_u6_u1_n175 ) , .C1( u0_u6_u1_n178 ) , .A( u0_u6_u1_n188 ) );
  INV_X1 u0_u6_u1_U31 (.ZN( u0_u6_u1_n188 ) , .A( u0_u6_u1_n97 ) );
  AOI211_X1 u0_u6_u1_U32 (.A( u0_u6_u1_n118 ) , .C1( u0_u6_u1_n132 ) , .C2( u0_u6_u1_n139 ) , .B( u0_u6_u1_n96 ) , .ZN( u0_u6_u1_n97 ) );
  AOI21_X1 u0_u6_u1_U33 (.B2( u0_u6_u1_n121 ) , .B1( u0_u6_u1_n135 ) , .A( u0_u6_u1_n152 ) , .ZN( u0_u6_u1_n96 ) );
  OAI221_X1 u0_u6_u1_U34 (.A( u0_u6_u1_n119 ) , .C2( u0_u6_u1_n129 ) , .ZN( u0_u6_u1_n138 ) , .B2( u0_u6_u1_n152 ) , .C1( u0_u6_u1_n174 ) , .B1( u0_u6_u1_n187 ) );
  INV_X1 u0_u6_u1_U35 (.A( u0_u6_u1_n148 ) , .ZN( u0_u6_u1_n187 ) );
  AOI211_X1 u0_u6_u1_U36 (.B( u0_u6_u1_n117 ) , .A( u0_u6_u1_n118 ) , .ZN( u0_u6_u1_n119 ) , .C2( u0_u6_u1_n146 ) , .C1( u0_u6_u1_n159 ) );
  NOR2_X1 u0_u6_u1_U37 (.A1( u0_u6_u1_n168 ) , .A2( u0_u6_u1_n176 ) , .ZN( u0_u6_u1_n98 ) );
  AOI211_X1 u0_u6_u1_U38 (.B( u0_u6_u1_n162 ) , .A( u0_u6_u1_n163 ) , .C2( u0_u6_u1_n164 ) , .ZN( u0_u6_u1_n165 ) , .C1( u0_u6_u1_n171 ) );
  AOI21_X1 u0_u6_u1_U39 (.A( u0_u6_u1_n160 ) , .B2( u0_u6_u1_n161 ) , .ZN( u0_u6_u1_n162 ) , .B1( u0_u6_u1_n182 ) );
  AOI221_X1 u0_u6_u1_U4 (.A( u0_u6_u1_n138 ) , .C2( u0_u6_u1_n139 ) , .C1( u0_u6_u1_n140 ) , .B2( u0_u6_u1_n141 ) , .ZN( u0_u6_u1_n142 ) , .B1( u0_u6_u1_n175 ) );
  OR2_X1 u0_u6_u1_U40 (.A2( u0_u6_u1_n157 ) , .A1( u0_u6_u1_n158 ) , .ZN( u0_u6_u1_n163 ) );
  NAND2_X1 u0_u6_u1_U41 (.A1( u0_u6_u1_n128 ) , .ZN( u0_u6_u1_n146 ) , .A2( u0_u6_u1_n160 ) );
  NAND2_X1 u0_u6_u1_U42 (.A2( u0_u6_u1_n112 ) , .ZN( u0_u6_u1_n139 ) , .A1( u0_u6_u1_n152 ) );
  NAND2_X1 u0_u6_u1_U43 (.A1( u0_u6_u1_n105 ) , .ZN( u0_u6_u1_n156 ) , .A2( u0_u6_u1_n99 ) );
  NOR2_X1 u0_u6_u1_U44 (.ZN( u0_u6_u1_n117 ) , .A1( u0_u6_u1_n121 ) , .A2( u0_u6_u1_n160 ) );
  OAI21_X1 u0_u6_u1_U45 (.B2( u0_u6_u1_n123 ) , .ZN( u0_u6_u1_n145 ) , .B1( u0_u6_u1_n160 ) , .A( u0_u6_u1_n185 ) );
  INV_X1 u0_u6_u1_U46 (.A( u0_u6_u1_n122 ) , .ZN( u0_u6_u1_n185 ) );
  AOI21_X1 u0_u6_u1_U47 (.B2( u0_u6_u1_n120 ) , .B1( u0_u6_u1_n121 ) , .ZN( u0_u6_u1_n122 ) , .A( u0_u6_u1_n128 ) );
  AOI21_X1 u0_u6_u1_U48 (.A( u0_u6_u1_n128 ) , .B2( u0_u6_u1_n129 ) , .ZN( u0_u6_u1_n130 ) , .B1( u0_u6_u1_n150 ) );
  NAND2_X1 u0_u6_u1_U49 (.ZN( u0_u6_u1_n112 ) , .A1( u0_u6_u1_n169 ) , .A2( u0_u6_u1_n170 ) );
  AOI211_X1 u0_u6_u1_U5 (.ZN( u0_u6_u1_n124 ) , .A( u0_u6_u1_n138 ) , .C2( u0_u6_u1_n139 ) , .B( u0_u6_u1_n145 ) , .C1( u0_u6_u1_n147 ) );
  NAND2_X1 u0_u6_u1_U50 (.ZN( u0_u6_u1_n129 ) , .A2( u0_u6_u1_n95 ) , .A1( u0_u6_u1_n98 ) );
  NAND2_X1 u0_u6_u1_U51 (.A1( u0_u6_u1_n102 ) , .ZN( u0_u6_u1_n154 ) , .A2( u0_u6_u1_n99 ) );
  NAND2_X1 u0_u6_u1_U52 (.A2( u0_u6_u1_n100 ) , .ZN( u0_u6_u1_n135 ) , .A1( u0_u6_u1_n99 ) );
  AOI21_X1 u0_u6_u1_U53 (.A( u0_u6_u1_n152 ) , .B2( u0_u6_u1_n153 ) , .B1( u0_u6_u1_n154 ) , .ZN( u0_u6_u1_n158 ) );
  INV_X1 u0_u6_u1_U54 (.A( u0_u6_u1_n160 ) , .ZN( u0_u6_u1_n175 ) );
  NAND2_X1 u0_u6_u1_U55 (.A1( u0_u6_u1_n100 ) , .ZN( u0_u6_u1_n116 ) , .A2( u0_u6_u1_n95 ) );
  NAND2_X1 u0_u6_u1_U56 (.A1( u0_u6_u1_n102 ) , .ZN( u0_u6_u1_n131 ) , .A2( u0_u6_u1_n95 ) );
  NAND2_X1 u0_u6_u1_U57 (.A2( u0_u6_u1_n104 ) , .ZN( u0_u6_u1_n121 ) , .A1( u0_u6_u1_n98 ) );
  NAND2_X1 u0_u6_u1_U58 (.A1( u0_u6_u1_n103 ) , .ZN( u0_u6_u1_n153 ) , .A2( u0_u6_u1_n98 ) );
  NAND2_X1 u0_u6_u1_U59 (.A2( u0_u6_u1_n104 ) , .A1( u0_u6_u1_n105 ) , .ZN( u0_u6_u1_n133 ) );
  AOI22_X1 u0_u6_u1_U6 (.B2( u0_u6_u1_n136 ) , .A2( u0_u6_u1_n137 ) , .ZN( u0_u6_u1_n143 ) , .A1( u0_u6_u1_n171 ) , .B1( u0_u6_u1_n173 ) );
  NAND2_X1 u0_u6_u1_U60 (.ZN( u0_u6_u1_n150 ) , .A2( u0_u6_u1_n98 ) , .A1( u0_u6_u1_n99 ) );
  NAND2_X1 u0_u6_u1_U61 (.A1( u0_u6_u1_n105 ) , .ZN( u0_u6_u1_n155 ) , .A2( u0_u6_u1_n95 ) );
  OAI21_X1 u0_u6_u1_U62 (.ZN( u0_u6_u1_n109 ) , .B1( u0_u6_u1_n129 ) , .B2( u0_u6_u1_n160 ) , .A( u0_u6_u1_n167 ) );
  NAND2_X1 u0_u6_u1_U63 (.A2( u0_u6_u1_n100 ) , .A1( u0_u6_u1_n103 ) , .ZN( u0_u6_u1_n120 ) );
  NAND2_X1 u0_u6_u1_U64 (.A1( u0_u6_u1_n102 ) , .A2( u0_u6_u1_n104 ) , .ZN( u0_u6_u1_n115 ) );
  NAND2_X1 u0_u6_u1_U65 (.A2( u0_u6_u1_n100 ) , .A1( u0_u6_u1_n104 ) , .ZN( u0_u6_u1_n151 ) );
  NAND2_X1 u0_u6_u1_U66 (.A2( u0_u6_u1_n103 ) , .A1( u0_u6_u1_n105 ) , .ZN( u0_u6_u1_n161 ) );
  INV_X1 u0_u6_u1_U67 (.A( u0_u6_u1_n152 ) , .ZN( u0_u6_u1_n173 ) );
  INV_X1 u0_u6_u1_U68 (.A( u0_u6_u1_n128 ) , .ZN( u0_u6_u1_n172 ) );
  NAND2_X1 u0_u6_u1_U69 (.A2( u0_u6_u1_n102 ) , .A1( u0_u6_u1_n103 ) , .ZN( u0_u6_u1_n123 ) );
  INV_X1 u0_u6_u1_U7 (.A( u0_u6_u1_n147 ) , .ZN( u0_u6_u1_n181 ) );
  NOR2_X1 u0_u6_u1_U70 (.A2( u0_u6_X_7 ) , .A1( u0_u6_X_8 ) , .ZN( u0_u6_u1_n95 ) );
  NOR2_X1 u0_u6_u1_U71 (.A1( u0_u6_X_12 ) , .A2( u0_u6_X_9 ) , .ZN( u0_u6_u1_n100 ) );
  NOR2_X1 u0_u6_u1_U72 (.A2( u0_u6_X_8 ) , .A1( u0_u6_u1_n177 ) , .ZN( u0_u6_u1_n99 ) );
  NOR2_X1 u0_u6_u1_U73 (.A2( u0_u6_X_12 ) , .ZN( u0_u6_u1_n102 ) , .A1( u0_u6_u1_n176 ) );
  NOR2_X1 u0_u6_u1_U74 (.A2( u0_u6_X_9 ) , .ZN( u0_u6_u1_n105 ) , .A1( u0_u6_u1_n168 ) );
  NAND2_X1 u0_u6_u1_U75 (.A1( u0_u6_X_10 ) , .ZN( u0_u6_u1_n160 ) , .A2( u0_u6_u1_n169 ) );
  NAND2_X1 u0_u6_u1_U76 (.A2( u0_u6_X_10 ) , .A1( u0_u6_X_11 ) , .ZN( u0_u6_u1_n152 ) );
  NAND2_X1 u0_u6_u1_U77 (.A1( u0_u6_X_11 ) , .ZN( u0_u6_u1_n128 ) , .A2( u0_u6_u1_n170 ) );
  AND2_X1 u0_u6_u1_U78 (.A2( u0_u6_X_7 ) , .A1( u0_u6_X_8 ) , .ZN( u0_u6_u1_n104 ) );
  AND2_X1 u0_u6_u1_U79 (.A1( u0_u6_X_8 ) , .ZN( u0_u6_u1_n103 ) , .A2( u0_u6_u1_n177 ) );
  NOR2_X1 u0_u6_u1_U8 (.A1( u0_u6_u1_n112 ) , .A2( u0_u6_u1_n116 ) , .ZN( u0_u6_u1_n118 ) );
  INV_X1 u0_u6_u1_U80 (.A( u0_u6_X_10 ) , .ZN( u0_u6_u1_n170 ) );
  INV_X1 u0_u6_u1_U81 (.A( u0_u6_X_9 ) , .ZN( u0_u6_u1_n176 ) );
  INV_X1 u0_u6_u1_U82 (.A( u0_u6_X_11 ) , .ZN( u0_u6_u1_n169 ) );
  INV_X1 u0_u6_u1_U83 (.A( u0_u6_X_12 ) , .ZN( u0_u6_u1_n168 ) );
  INV_X1 u0_u6_u1_U84 (.A( u0_u6_X_7 ) , .ZN( u0_u6_u1_n177 ) );
  NAND4_X1 u0_u6_u1_U85 (.ZN( u0_out6_28 ) , .A4( u0_u6_u1_n124 ) , .A3( u0_u6_u1_n125 ) , .A2( u0_u6_u1_n126 ) , .A1( u0_u6_u1_n127 ) );
  OAI21_X1 u0_u6_u1_U86 (.ZN( u0_u6_u1_n127 ) , .B2( u0_u6_u1_n139 ) , .B1( u0_u6_u1_n175 ) , .A( u0_u6_u1_n183 ) );
  OAI21_X1 u0_u6_u1_U87 (.ZN( u0_u6_u1_n126 ) , .B2( u0_u6_u1_n140 ) , .A( u0_u6_u1_n146 ) , .B1( u0_u6_u1_n178 ) );
  NAND4_X1 u0_u6_u1_U88 (.ZN( u0_out6_18 ) , .A4( u0_u6_u1_n165 ) , .A3( u0_u6_u1_n166 ) , .A1( u0_u6_u1_n167 ) , .A2( u0_u6_u1_n186 ) );
  AOI22_X1 u0_u6_u1_U89 (.B2( u0_u6_u1_n146 ) , .B1( u0_u6_u1_n147 ) , .A2( u0_u6_u1_n148 ) , .ZN( u0_u6_u1_n166 ) , .A1( u0_u6_u1_n172 ) );
  OAI21_X1 u0_u6_u1_U9 (.ZN( u0_u6_u1_n101 ) , .B1( u0_u6_u1_n141 ) , .A( u0_u6_u1_n146 ) , .B2( u0_u6_u1_n183 ) );
  INV_X1 u0_u6_u1_U90 (.A( u0_u6_u1_n145 ) , .ZN( u0_u6_u1_n186 ) );
  NAND4_X1 u0_u6_u1_U91 (.ZN( u0_out6_2 ) , .A4( u0_u6_u1_n142 ) , .A3( u0_u6_u1_n143 ) , .A2( u0_u6_u1_n144 ) , .A1( u0_u6_u1_n179 ) );
  OAI21_X1 u0_u6_u1_U92 (.B2( u0_u6_u1_n132 ) , .ZN( u0_u6_u1_n144 ) , .A( u0_u6_u1_n146 ) , .B1( u0_u6_u1_n180 ) );
  INV_X1 u0_u6_u1_U93 (.A( u0_u6_u1_n130 ) , .ZN( u0_u6_u1_n179 ) );
  OR4_X1 u0_u6_u1_U94 (.ZN( u0_out6_13 ) , .A4( u0_u6_u1_n108 ) , .A3( u0_u6_u1_n109 ) , .A2( u0_u6_u1_n110 ) , .A1( u0_u6_u1_n111 ) );
  AOI21_X1 u0_u6_u1_U95 (.ZN( u0_u6_u1_n111 ) , .A( u0_u6_u1_n128 ) , .B2( u0_u6_u1_n131 ) , .B1( u0_u6_u1_n135 ) );
  AOI21_X1 u0_u6_u1_U96 (.ZN( u0_u6_u1_n110 ) , .A( u0_u6_u1_n116 ) , .B1( u0_u6_u1_n152 ) , .B2( u0_u6_u1_n160 ) );
  NAND3_X1 u0_u6_u1_U97 (.A3( u0_u6_u1_n149 ) , .A2( u0_u6_u1_n150 ) , .A1( u0_u6_u1_n151 ) , .ZN( u0_u6_u1_n164 ) );
  NAND3_X1 u0_u6_u1_U98 (.A3( u0_u6_u1_n134 ) , .A2( u0_u6_u1_n135 ) , .ZN( u0_u6_u1_n136 ) , .A1( u0_u6_u1_n151 ) );
  NAND3_X1 u0_u6_u1_U99 (.A1( u0_u6_u1_n133 ) , .ZN( u0_u6_u1_n137 ) , .A2( u0_u6_u1_n154 ) , .A3( u0_u6_u1_n181 ) );
  OAI22_X1 u0_u6_u2_U10 (.B1( u0_u6_u2_n151 ) , .A2( u0_u6_u2_n152 ) , .A1( u0_u6_u2_n153 ) , .ZN( u0_u6_u2_n160 ) , .B2( u0_u6_u2_n168 ) );
  NAND3_X1 u0_u6_u2_U100 (.A2( u0_u6_u2_n100 ) , .A1( u0_u6_u2_n104 ) , .A3( u0_u6_u2_n138 ) , .ZN( u0_u6_u2_n98 ) );
  NOR3_X1 u0_u6_u2_U11 (.A1( u0_u6_u2_n150 ) , .ZN( u0_u6_u2_n151 ) , .A3( u0_u6_u2_n175 ) , .A2( u0_u6_u2_n188 ) );
  AOI21_X1 u0_u6_u2_U12 (.B2( u0_u6_u2_n123 ) , .ZN( u0_u6_u2_n125 ) , .A( u0_u6_u2_n171 ) , .B1( u0_u6_u2_n184 ) );
  INV_X1 u0_u6_u2_U13 (.A( u0_u6_u2_n150 ) , .ZN( u0_u6_u2_n184 ) );
  AOI21_X1 u0_u6_u2_U14 (.ZN( u0_u6_u2_n144 ) , .B2( u0_u6_u2_n155 ) , .A( u0_u6_u2_n172 ) , .B1( u0_u6_u2_n185 ) );
  AOI21_X1 u0_u6_u2_U15 (.B2( u0_u6_u2_n143 ) , .ZN( u0_u6_u2_n145 ) , .B1( u0_u6_u2_n152 ) , .A( u0_u6_u2_n171 ) );
  INV_X1 u0_u6_u2_U16 (.A( u0_u6_u2_n156 ) , .ZN( u0_u6_u2_n171 ) );
  INV_X1 u0_u6_u2_U17 (.A( u0_u6_u2_n120 ) , .ZN( u0_u6_u2_n188 ) );
  NAND2_X1 u0_u6_u2_U18 (.A2( u0_u6_u2_n122 ) , .ZN( u0_u6_u2_n150 ) , .A1( u0_u6_u2_n152 ) );
  INV_X1 u0_u6_u2_U19 (.A( u0_u6_u2_n153 ) , .ZN( u0_u6_u2_n170 ) );
  INV_X1 u0_u6_u2_U20 (.A( u0_u6_u2_n137 ) , .ZN( u0_u6_u2_n173 ) );
  NAND2_X1 u0_u6_u2_U21 (.A1( u0_u6_u2_n132 ) , .A2( u0_u6_u2_n139 ) , .ZN( u0_u6_u2_n157 ) );
  INV_X1 u0_u6_u2_U22 (.A( u0_u6_u2_n113 ) , .ZN( u0_u6_u2_n178 ) );
  INV_X1 u0_u6_u2_U23 (.A( u0_u6_u2_n139 ) , .ZN( u0_u6_u2_n175 ) );
  INV_X1 u0_u6_u2_U24 (.A( u0_u6_u2_n155 ) , .ZN( u0_u6_u2_n181 ) );
  INV_X1 u0_u6_u2_U25 (.A( u0_u6_u2_n119 ) , .ZN( u0_u6_u2_n177 ) );
  INV_X1 u0_u6_u2_U26 (.A( u0_u6_u2_n116 ) , .ZN( u0_u6_u2_n180 ) );
  INV_X1 u0_u6_u2_U27 (.A( u0_u6_u2_n131 ) , .ZN( u0_u6_u2_n179 ) );
  INV_X1 u0_u6_u2_U28 (.A( u0_u6_u2_n154 ) , .ZN( u0_u6_u2_n176 ) );
  NAND2_X1 u0_u6_u2_U29 (.A2( u0_u6_u2_n116 ) , .A1( u0_u6_u2_n117 ) , .ZN( u0_u6_u2_n118 ) );
  NOR2_X1 u0_u6_u2_U3 (.ZN( u0_u6_u2_n121 ) , .A2( u0_u6_u2_n177 ) , .A1( u0_u6_u2_n180 ) );
  INV_X1 u0_u6_u2_U30 (.A( u0_u6_u2_n132 ) , .ZN( u0_u6_u2_n182 ) );
  INV_X1 u0_u6_u2_U31 (.A( u0_u6_u2_n158 ) , .ZN( u0_u6_u2_n183 ) );
  OAI21_X1 u0_u6_u2_U32 (.A( u0_u6_u2_n156 ) , .B1( u0_u6_u2_n157 ) , .ZN( u0_u6_u2_n158 ) , .B2( u0_u6_u2_n179 ) );
  NOR2_X1 u0_u6_u2_U33 (.ZN( u0_u6_u2_n156 ) , .A1( u0_u6_u2_n166 ) , .A2( u0_u6_u2_n169 ) );
  NOR2_X1 u0_u6_u2_U34 (.A2( u0_u6_u2_n114 ) , .ZN( u0_u6_u2_n137 ) , .A1( u0_u6_u2_n140 ) );
  NOR2_X1 u0_u6_u2_U35 (.A2( u0_u6_u2_n138 ) , .ZN( u0_u6_u2_n153 ) , .A1( u0_u6_u2_n156 ) );
  AOI211_X1 u0_u6_u2_U36 (.ZN( u0_u6_u2_n130 ) , .C1( u0_u6_u2_n138 ) , .C2( u0_u6_u2_n179 ) , .B( u0_u6_u2_n96 ) , .A( u0_u6_u2_n97 ) );
  OAI22_X1 u0_u6_u2_U37 (.B1( u0_u6_u2_n133 ) , .A2( u0_u6_u2_n137 ) , .A1( u0_u6_u2_n152 ) , .B2( u0_u6_u2_n168 ) , .ZN( u0_u6_u2_n97 ) );
  OAI221_X1 u0_u6_u2_U38 (.B1( u0_u6_u2_n113 ) , .C1( u0_u6_u2_n132 ) , .A( u0_u6_u2_n149 ) , .B2( u0_u6_u2_n171 ) , .C2( u0_u6_u2_n172 ) , .ZN( u0_u6_u2_n96 ) );
  OAI221_X1 u0_u6_u2_U39 (.A( u0_u6_u2_n115 ) , .C2( u0_u6_u2_n123 ) , .B2( u0_u6_u2_n143 ) , .B1( u0_u6_u2_n153 ) , .ZN( u0_u6_u2_n163 ) , .C1( u0_u6_u2_n168 ) );
  INV_X1 u0_u6_u2_U4 (.A( u0_u6_u2_n134 ) , .ZN( u0_u6_u2_n185 ) );
  OAI21_X1 u0_u6_u2_U40 (.A( u0_u6_u2_n114 ) , .ZN( u0_u6_u2_n115 ) , .B1( u0_u6_u2_n176 ) , .B2( u0_u6_u2_n178 ) );
  OAI221_X1 u0_u6_u2_U41 (.A( u0_u6_u2_n135 ) , .B2( u0_u6_u2_n136 ) , .B1( u0_u6_u2_n137 ) , .ZN( u0_u6_u2_n162 ) , .C2( u0_u6_u2_n167 ) , .C1( u0_u6_u2_n185 ) );
  AND3_X1 u0_u6_u2_U42 (.A3( u0_u6_u2_n131 ) , .A2( u0_u6_u2_n132 ) , .A1( u0_u6_u2_n133 ) , .ZN( u0_u6_u2_n136 ) );
  AOI22_X1 u0_u6_u2_U43 (.ZN( u0_u6_u2_n135 ) , .B1( u0_u6_u2_n140 ) , .A1( u0_u6_u2_n156 ) , .B2( u0_u6_u2_n180 ) , .A2( u0_u6_u2_n188 ) );
  AOI21_X1 u0_u6_u2_U44 (.ZN( u0_u6_u2_n149 ) , .B1( u0_u6_u2_n173 ) , .B2( u0_u6_u2_n188 ) , .A( u0_u6_u2_n95 ) );
  AND3_X1 u0_u6_u2_U45 (.A2( u0_u6_u2_n100 ) , .A1( u0_u6_u2_n104 ) , .A3( u0_u6_u2_n156 ) , .ZN( u0_u6_u2_n95 ) );
  OAI21_X1 u0_u6_u2_U46 (.A( u0_u6_u2_n141 ) , .B2( u0_u6_u2_n142 ) , .ZN( u0_u6_u2_n146 ) , .B1( u0_u6_u2_n153 ) );
  OAI21_X1 u0_u6_u2_U47 (.A( u0_u6_u2_n140 ) , .ZN( u0_u6_u2_n141 ) , .B1( u0_u6_u2_n176 ) , .B2( u0_u6_u2_n177 ) );
  NOR3_X1 u0_u6_u2_U48 (.ZN( u0_u6_u2_n142 ) , .A3( u0_u6_u2_n175 ) , .A2( u0_u6_u2_n178 ) , .A1( u0_u6_u2_n181 ) );
  OAI21_X1 u0_u6_u2_U49 (.A( u0_u6_u2_n101 ) , .B2( u0_u6_u2_n121 ) , .B1( u0_u6_u2_n153 ) , .ZN( u0_u6_u2_n164 ) );
  NOR4_X1 u0_u6_u2_U5 (.A4( u0_u6_u2_n124 ) , .A3( u0_u6_u2_n125 ) , .A2( u0_u6_u2_n126 ) , .A1( u0_u6_u2_n127 ) , .ZN( u0_u6_u2_n128 ) );
  NAND2_X1 u0_u6_u2_U50 (.A2( u0_u6_u2_n100 ) , .A1( u0_u6_u2_n107 ) , .ZN( u0_u6_u2_n155 ) );
  NAND2_X1 u0_u6_u2_U51 (.A2( u0_u6_u2_n105 ) , .A1( u0_u6_u2_n108 ) , .ZN( u0_u6_u2_n143 ) );
  NAND2_X1 u0_u6_u2_U52 (.A1( u0_u6_u2_n104 ) , .A2( u0_u6_u2_n106 ) , .ZN( u0_u6_u2_n152 ) );
  NAND2_X1 u0_u6_u2_U53 (.A1( u0_u6_u2_n100 ) , .A2( u0_u6_u2_n105 ) , .ZN( u0_u6_u2_n132 ) );
  INV_X1 u0_u6_u2_U54 (.A( u0_u6_u2_n140 ) , .ZN( u0_u6_u2_n168 ) );
  INV_X1 u0_u6_u2_U55 (.A( u0_u6_u2_n138 ) , .ZN( u0_u6_u2_n167 ) );
  INV_X1 u0_u6_u2_U56 (.ZN( u0_u6_u2_n187 ) , .A( u0_u6_u2_n99 ) );
  OAI21_X1 u0_u6_u2_U57 (.B1( u0_u6_u2_n137 ) , .B2( u0_u6_u2_n143 ) , .A( u0_u6_u2_n98 ) , .ZN( u0_u6_u2_n99 ) );
  NAND2_X1 u0_u6_u2_U58 (.A1( u0_u6_u2_n102 ) , .A2( u0_u6_u2_n106 ) , .ZN( u0_u6_u2_n113 ) );
  NAND2_X1 u0_u6_u2_U59 (.A1( u0_u6_u2_n106 ) , .A2( u0_u6_u2_n107 ) , .ZN( u0_u6_u2_n131 ) );
  AOI21_X1 u0_u6_u2_U6 (.B2( u0_u6_u2_n119 ) , .ZN( u0_u6_u2_n127 ) , .A( u0_u6_u2_n137 ) , .B1( u0_u6_u2_n155 ) );
  NAND2_X1 u0_u6_u2_U60 (.A1( u0_u6_u2_n103 ) , .A2( u0_u6_u2_n107 ) , .ZN( u0_u6_u2_n139 ) );
  NAND2_X1 u0_u6_u2_U61 (.A1( u0_u6_u2_n103 ) , .A2( u0_u6_u2_n105 ) , .ZN( u0_u6_u2_n133 ) );
  NAND2_X1 u0_u6_u2_U62 (.A1( u0_u6_u2_n102 ) , .A2( u0_u6_u2_n103 ) , .ZN( u0_u6_u2_n154 ) );
  NAND2_X1 u0_u6_u2_U63 (.A2( u0_u6_u2_n103 ) , .A1( u0_u6_u2_n104 ) , .ZN( u0_u6_u2_n119 ) );
  NAND2_X1 u0_u6_u2_U64 (.A2( u0_u6_u2_n107 ) , .A1( u0_u6_u2_n108 ) , .ZN( u0_u6_u2_n123 ) );
  NAND2_X1 u0_u6_u2_U65 (.A1( u0_u6_u2_n104 ) , .A2( u0_u6_u2_n108 ) , .ZN( u0_u6_u2_n122 ) );
  INV_X1 u0_u6_u2_U66 (.A( u0_u6_u2_n114 ) , .ZN( u0_u6_u2_n172 ) );
  NAND2_X1 u0_u6_u2_U67 (.A2( u0_u6_u2_n100 ) , .A1( u0_u6_u2_n102 ) , .ZN( u0_u6_u2_n116 ) );
  NAND2_X1 u0_u6_u2_U68 (.A1( u0_u6_u2_n102 ) , .A2( u0_u6_u2_n108 ) , .ZN( u0_u6_u2_n120 ) );
  NAND2_X1 u0_u6_u2_U69 (.A2( u0_u6_u2_n105 ) , .A1( u0_u6_u2_n106 ) , .ZN( u0_u6_u2_n117 ) );
  AOI21_X1 u0_u6_u2_U7 (.ZN( u0_u6_u2_n124 ) , .B1( u0_u6_u2_n131 ) , .B2( u0_u6_u2_n143 ) , .A( u0_u6_u2_n172 ) );
  NOR2_X1 u0_u6_u2_U70 (.A2( u0_u6_X_16 ) , .ZN( u0_u6_u2_n140 ) , .A1( u0_u6_u2_n166 ) );
  NOR2_X1 u0_u6_u2_U71 (.A2( u0_u6_X_13 ) , .A1( u0_u6_X_14 ) , .ZN( u0_u6_u2_n100 ) );
  NOR2_X1 u0_u6_u2_U72 (.A2( u0_u6_X_16 ) , .A1( u0_u6_X_17 ) , .ZN( u0_u6_u2_n138 ) );
  NOR2_X1 u0_u6_u2_U73 (.A2( u0_u6_X_15 ) , .A1( u0_u6_X_18 ) , .ZN( u0_u6_u2_n104 ) );
  NOR2_X1 u0_u6_u2_U74 (.A2( u0_u6_X_14 ) , .ZN( u0_u6_u2_n103 ) , .A1( u0_u6_u2_n174 ) );
  NOR2_X1 u0_u6_u2_U75 (.A2( u0_u6_X_15 ) , .ZN( u0_u6_u2_n102 ) , .A1( u0_u6_u2_n165 ) );
  NOR2_X1 u0_u6_u2_U76 (.A2( u0_u6_X_17 ) , .ZN( u0_u6_u2_n114 ) , .A1( u0_u6_u2_n169 ) );
  AND2_X1 u0_u6_u2_U77 (.A1( u0_u6_X_15 ) , .ZN( u0_u6_u2_n105 ) , .A2( u0_u6_u2_n165 ) );
  AND2_X1 u0_u6_u2_U78 (.A2( u0_u6_X_15 ) , .A1( u0_u6_X_18 ) , .ZN( u0_u6_u2_n107 ) );
  AND2_X1 u0_u6_u2_U79 (.A1( u0_u6_X_14 ) , .ZN( u0_u6_u2_n106 ) , .A2( u0_u6_u2_n174 ) );
  AOI21_X1 u0_u6_u2_U8 (.B2( u0_u6_u2_n120 ) , .B1( u0_u6_u2_n121 ) , .ZN( u0_u6_u2_n126 ) , .A( u0_u6_u2_n167 ) );
  AND2_X1 u0_u6_u2_U80 (.A1( u0_u6_X_13 ) , .A2( u0_u6_X_14 ) , .ZN( u0_u6_u2_n108 ) );
  INV_X1 u0_u6_u2_U81 (.A( u0_u6_X_16 ) , .ZN( u0_u6_u2_n169 ) );
  INV_X1 u0_u6_u2_U82 (.A( u0_u6_X_17 ) , .ZN( u0_u6_u2_n166 ) );
  INV_X1 u0_u6_u2_U83 (.A( u0_u6_X_13 ) , .ZN( u0_u6_u2_n174 ) );
  INV_X1 u0_u6_u2_U84 (.A( u0_u6_X_18 ) , .ZN( u0_u6_u2_n165 ) );
  NAND4_X1 u0_u6_u2_U85 (.ZN( u0_out6_30 ) , .A4( u0_u6_u2_n147 ) , .A3( u0_u6_u2_n148 ) , .A2( u0_u6_u2_n149 ) , .A1( u0_u6_u2_n187 ) );
  AOI21_X1 u0_u6_u2_U86 (.B2( u0_u6_u2_n138 ) , .ZN( u0_u6_u2_n148 ) , .A( u0_u6_u2_n162 ) , .B1( u0_u6_u2_n182 ) );
  NOR3_X1 u0_u6_u2_U87 (.A3( u0_u6_u2_n144 ) , .A2( u0_u6_u2_n145 ) , .A1( u0_u6_u2_n146 ) , .ZN( u0_u6_u2_n147 ) );
  NAND4_X1 u0_u6_u2_U88 (.ZN( u0_out6_24 ) , .A4( u0_u6_u2_n111 ) , .A3( u0_u6_u2_n112 ) , .A1( u0_u6_u2_n130 ) , .A2( u0_u6_u2_n187 ) );
  AOI221_X1 u0_u6_u2_U89 (.A( u0_u6_u2_n109 ) , .B1( u0_u6_u2_n110 ) , .ZN( u0_u6_u2_n111 ) , .C1( u0_u6_u2_n134 ) , .C2( u0_u6_u2_n170 ) , .B2( u0_u6_u2_n173 ) );
  OAI22_X1 u0_u6_u2_U9 (.ZN( u0_u6_u2_n109 ) , .A2( u0_u6_u2_n113 ) , .B2( u0_u6_u2_n133 ) , .B1( u0_u6_u2_n167 ) , .A1( u0_u6_u2_n168 ) );
  AOI21_X1 u0_u6_u2_U90 (.ZN( u0_u6_u2_n112 ) , .B2( u0_u6_u2_n156 ) , .A( u0_u6_u2_n164 ) , .B1( u0_u6_u2_n181 ) );
  NAND4_X1 u0_u6_u2_U91 (.ZN( u0_out6_16 ) , .A4( u0_u6_u2_n128 ) , .A3( u0_u6_u2_n129 ) , .A1( u0_u6_u2_n130 ) , .A2( u0_u6_u2_n186 ) );
  AOI22_X1 u0_u6_u2_U92 (.A2( u0_u6_u2_n118 ) , .ZN( u0_u6_u2_n129 ) , .A1( u0_u6_u2_n140 ) , .B1( u0_u6_u2_n157 ) , .B2( u0_u6_u2_n170 ) );
  INV_X1 u0_u6_u2_U93 (.A( u0_u6_u2_n163 ) , .ZN( u0_u6_u2_n186 ) );
  OR4_X1 u0_u6_u2_U94 (.ZN( u0_out6_6 ) , .A4( u0_u6_u2_n161 ) , .A3( u0_u6_u2_n162 ) , .A2( u0_u6_u2_n163 ) , .A1( u0_u6_u2_n164 ) );
  OR3_X1 u0_u6_u2_U95 (.A2( u0_u6_u2_n159 ) , .A1( u0_u6_u2_n160 ) , .ZN( u0_u6_u2_n161 ) , .A3( u0_u6_u2_n183 ) );
  AOI21_X1 u0_u6_u2_U96 (.B2( u0_u6_u2_n154 ) , .B1( u0_u6_u2_n155 ) , .ZN( u0_u6_u2_n159 ) , .A( u0_u6_u2_n167 ) );
  NAND3_X1 u0_u6_u2_U97 (.A2( u0_u6_u2_n117 ) , .A1( u0_u6_u2_n122 ) , .A3( u0_u6_u2_n123 ) , .ZN( u0_u6_u2_n134 ) );
  NAND3_X1 u0_u6_u2_U98 (.ZN( u0_u6_u2_n110 ) , .A2( u0_u6_u2_n131 ) , .A3( u0_u6_u2_n139 ) , .A1( u0_u6_u2_n154 ) );
  NAND3_X1 u0_u6_u2_U99 (.A2( u0_u6_u2_n100 ) , .ZN( u0_u6_u2_n101 ) , .A1( u0_u6_u2_n104 ) , .A3( u0_u6_u2_n114 ) );
  OAI22_X1 u0_u6_u3_U10 (.B1( u0_u6_u3_n113 ) , .A2( u0_u6_u3_n135 ) , .A1( u0_u6_u3_n150 ) , .B2( u0_u6_u3_n164 ) , .ZN( u0_u6_u3_n98 ) );
  OAI211_X1 u0_u6_u3_U11 (.B( u0_u6_u3_n106 ) , .ZN( u0_u6_u3_n119 ) , .C2( u0_u6_u3_n128 ) , .C1( u0_u6_u3_n167 ) , .A( u0_u6_u3_n181 ) );
  AOI221_X1 u0_u6_u3_U12 (.C1( u0_u6_u3_n105 ) , .ZN( u0_u6_u3_n106 ) , .A( u0_u6_u3_n131 ) , .B2( u0_u6_u3_n132 ) , .C2( u0_u6_u3_n133 ) , .B1( u0_u6_u3_n169 ) );
  INV_X1 u0_u6_u3_U13 (.ZN( u0_u6_u3_n181 ) , .A( u0_u6_u3_n98 ) );
  NAND2_X1 u0_u6_u3_U14 (.ZN( u0_u6_u3_n105 ) , .A2( u0_u6_u3_n130 ) , .A1( u0_u6_u3_n155 ) );
  NOR2_X1 u0_u6_u3_U15 (.ZN( u0_u6_u3_n126 ) , .A2( u0_u6_u3_n150 ) , .A1( u0_u6_u3_n164 ) );
  AOI21_X1 u0_u6_u3_U16 (.ZN( u0_u6_u3_n112 ) , .B2( u0_u6_u3_n146 ) , .B1( u0_u6_u3_n155 ) , .A( u0_u6_u3_n167 ) );
  NAND2_X1 u0_u6_u3_U17 (.A1( u0_u6_u3_n135 ) , .ZN( u0_u6_u3_n142 ) , .A2( u0_u6_u3_n164 ) );
  NAND2_X1 u0_u6_u3_U18 (.ZN( u0_u6_u3_n132 ) , .A2( u0_u6_u3_n152 ) , .A1( u0_u6_u3_n156 ) );
  AND2_X1 u0_u6_u3_U19 (.A2( u0_u6_u3_n113 ) , .A1( u0_u6_u3_n114 ) , .ZN( u0_u6_u3_n151 ) );
  INV_X1 u0_u6_u3_U20 (.A( u0_u6_u3_n133 ) , .ZN( u0_u6_u3_n165 ) );
  INV_X1 u0_u6_u3_U21 (.A( u0_u6_u3_n135 ) , .ZN( u0_u6_u3_n170 ) );
  NAND2_X1 u0_u6_u3_U22 (.A1( u0_u6_u3_n107 ) , .A2( u0_u6_u3_n108 ) , .ZN( u0_u6_u3_n140 ) );
  NAND2_X1 u0_u6_u3_U23 (.ZN( u0_u6_u3_n117 ) , .A1( u0_u6_u3_n124 ) , .A2( u0_u6_u3_n148 ) );
  NAND2_X1 u0_u6_u3_U24 (.ZN( u0_u6_u3_n143 ) , .A1( u0_u6_u3_n165 ) , .A2( u0_u6_u3_n167 ) );
  INV_X1 u0_u6_u3_U25 (.A( u0_u6_u3_n130 ) , .ZN( u0_u6_u3_n177 ) );
  INV_X1 u0_u6_u3_U26 (.A( u0_u6_u3_n128 ) , .ZN( u0_u6_u3_n176 ) );
  INV_X1 u0_u6_u3_U27 (.A( u0_u6_u3_n155 ) , .ZN( u0_u6_u3_n174 ) );
  AOI22_X1 u0_u6_u3_U28 (.B1( u0_u6_u3_n115 ) , .A2( u0_u6_u3_n116 ) , .ZN( u0_u6_u3_n123 ) , .B2( u0_u6_u3_n133 ) , .A1( u0_u6_u3_n169 ) );
  NAND2_X1 u0_u6_u3_U29 (.ZN( u0_u6_u3_n116 ) , .A2( u0_u6_u3_n151 ) , .A1( u0_u6_u3_n182 ) );
  INV_X1 u0_u6_u3_U3 (.A( u0_u6_u3_n129 ) , .ZN( u0_u6_u3_n183 ) );
  INV_X1 u0_u6_u3_U30 (.A( u0_u6_u3_n139 ) , .ZN( u0_u6_u3_n185 ) );
  NOR2_X1 u0_u6_u3_U31 (.ZN( u0_u6_u3_n135 ) , .A2( u0_u6_u3_n141 ) , .A1( u0_u6_u3_n169 ) );
  OAI222_X1 u0_u6_u3_U32 (.C2( u0_u6_u3_n107 ) , .A2( u0_u6_u3_n108 ) , .B1( u0_u6_u3_n135 ) , .ZN( u0_u6_u3_n138 ) , .B2( u0_u6_u3_n146 ) , .C1( u0_u6_u3_n154 ) , .A1( u0_u6_u3_n164 ) );
  NOR4_X1 u0_u6_u3_U33 (.A4( u0_u6_u3_n157 ) , .A3( u0_u6_u3_n158 ) , .A2( u0_u6_u3_n159 ) , .A1( u0_u6_u3_n160 ) , .ZN( u0_u6_u3_n161 ) );
  AOI21_X1 u0_u6_u3_U34 (.B2( u0_u6_u3_n152 ) , .B1( u0_u6_u3_n153 ) , .ZN( u0_u6_u3_n158 ) , .A( u0_u6_u3_n164 ) );
  AOI21_X1 u0_u6_u3_U35 (.A( u0_u6_u3_n154 ) , .B2( u0_u6_u3_n155 ) , .B1( u0_u6_u3_n156 ) , .ZN( u0_u6_u3_n157 ) );
  AOI21_X1 u0_u6_u3_U36 (.A( u0_u6_u3_n149 ) , .B2( u0_u6_u3_n150 ) , .B1( u0_u6_u3_n151 ) , .ZN( u0_u6_u3_n159 ) );
  AOI211_X1 u0_u6_u3_U37 (.ZN( u0_u6_u3_n109 ) , .A( u0_u6_u3_n119 ) , .C2( u0_u6_u3_n129 ) , .B( u0_u6_u3_n138 ) , .C1( u0_u6_u3_n141 ) );
  AOI211_X1 u0_u6_u3_U38 (.B( u0_u6_u3_n119 ) , .A( u0_u6_u3_n120 ) , .C2( u0_u6_u3_n121 ) , .ZN( u0_u6_u3_n122 ) , .C1( u0_u6_u3_n179 ) );
  INV_X1 u0_u6_u3_U39 (.A( u0_u6_u3_n156 ) , .ZN( u0_u6_u3_n179 ) );
  INV_X1 u0_u6_u3_U4 (.A( u0_u6_u3_n140 ) , .ZN( u0_u6_u3_n182 ) );
  OAI22_X1 u0_u6_u3_U40 (.B1( u0_u6_u3_n118 ) , .ZN( u0_u6_u3_n120 ) , .A1( u0_u6_u3_n135 ) , .B2( u0_u6_u3_n154 ) , .A2( u0_u6_u3_n178 ) );
  AND3_X1 u0_u6_u3_U41 (.ZN( u0_u6_u3_n118 ) , .A2( u0_u6_u3_n124 ) , .A1( u0_u6_u3_n144 ) , .A3( u0_u6_u3_n152 ) );
  INV_X1 u0_u6_u3_U42 (.A( u0_u6_u3_n121 ) , .ZN( u0_u6_u3_n164 ) );
  NAND2_X1 u0_u6_u3_U43 (.ZN( u0_u6_u3_n133 ) , .A1( u0_u6_u3_n154 ) , .A2( u0_u6_u3_n164 ) );
  OAI211_X1 u0_u6_u3_U44 (.B( u0_u6_u3_n127 ) , .ZN( u0_u6_u3_n139 ) , .C1( u0_u6_u3_n150 ) , .C2( u0_u6_u3_n154 ) , .A( u0_u6_u3_n184 ) );
  INV_X1 u0_u6_u3_U45 (.A( u0_u6_u3_n125 ) , .ZN( u0_u6_u3_n184 ) );
  AOI221_X1 u0_u6_u3_U46 (.A( u0_u6_u3_n126 ) , .ZN( u0_u6_u3_n127 ) , .C2( u0_u6_u3_n132 ) , .C1( u0_u6_u3_n169 ) , .B2( u0_u6_u3_n170 ) , .B1( u0_u6_u3_n174 ) );
  OAI22_X1 u0_u6_u3_U47 (.A1( u0_u6_u3_n124 ) , .ZN( u0_u6_u3_n125 ) , .B2( u0_u6_u3_n145 ) , .A2( u0_u6_u3_n165 ) , .B1( u0_u6_u3_n167 ) );
  NOR2_X1 u0_u6_u3_U48 (.A1( u0_u6_u3_n113 ) , .ZN( u0_u6_u3_n131 ) , .A2( u0_u6_u3_n154 ) );
  NAND2_X1 u0_u6_u3_U49 (.A1( u0_u6_u3_n103 ) , .ZN( u0_u6_u3_n150 ) , .A2( u0_u6_u3_n99 ) );
  INV_X1 u0_u6_u3_U5 (.A( u0_u6_u3_n117 ) , .ZN( u0_u6_u3_n178 ) );
  NAND2_X1 u0_u6_u3_U50 (.A2( u0_u6_u3_n102 ) , .ZN( u0_u6_u3_n155 ) , .A1( u0_u6_u3_n97 ) );
  INV_X1 u0_u6_u3_U51 (.A( u0_u6_u3_n141 ) , .ZN( u0_u6_u3_n167 ) );
  AOI21_X1 u0_u6_u3_U52 (.B2( u0_u6_u3_n114 ) , .B1( u0_u6_u3_n146 ) , .A( u0_u6_u3_n154 ) , .ZN( u0_u6_u3_n94 ) );
  AOI21_X1 u0_u6_u3_U53 (.ZN( u0_u6_u3_n110 ) , .B2( u0_u6_u3_n142 ) , .B1( u0_u6_u3_n186 ) , .A( u0_u6_u3_n95 ) );
  INV_X1 u0_u6_u3_U54 (.A( u0_u6_u3_n145 ) , .ZN( u0_u6_u3_n186 ) );
  AOI21_X1 u0_u6_u3_U55 (.B1( u0_u6_u3_n124 ) , .A( u0_u6_u3_n149 ) , .B2( u0_u6_u3_n155 ) , .ZN( u0_u6_u3_n95 ) );
  INV_X1 u0_u6_u3_U56 (.A( u0_u6_u3_n149 ) , .ZN( u0_u6_u3_n169 ) );
  NAND2_X1 u0_u6_u3_U57 (.ZN( u0_u6_u3_n124 ) , .A1( u0_u6_u3_n96 ) , .A2( u0_u6_u3_n97 ) );
  NAND2_X1 u0_u6_u3_U58 (.A2( u0_u6_u3_n100 ) , .ZN( u0_u6_u3_n146 ) , .A1( u0_u6_u3_n96 ) );
  NAND2_X1 u0_u6_u3_U59 (.A1( u0_u6_u3_n101 ) , .ZN( u0_u6_u3_n145 ) , .A2( u0_u6_u3_n99 ) );
  AOI221_X1 u0_u6_u3_U6 (.A( u0_u6_u3_n131 ) , .C2( u0_u6_u3_n132 ) , .C1( u0_u6_u3_n133 ) , .ZN( u0_u6_u3_n134 ) , .B1( u0_u6_u3_n143 ) , .B2( u0_u6_u3_n177 ) );
  NAND2_X1 u0_u6_u3_U60 (.A1( u0_u6_u3_n100 ) , .ZN( u0_u6_u3_n156 ) , .A2( u0_u6_u3_n99 ) );
  NAND2_X1 u0_u6_u3_U61 (.A2( u0_u6_u3_n101 ) , .A1( u0_u6_u3_n104 ) , .ZN( u0_u6_u3_n148 ) );
  NAND2_X1 u0_u6_u3_U62 (.A1( u0_u6_u3_n100 ) , .A2( u0_u6_u3_n102 ) , .ZN( u0_u6_u3_n128 ) );
  NAND2_X1 u0_u6_u3_U63 (.A2( u0_u6_u3_n101 ) , .A1( u0_u6_u3_n102 ) , .ZN( u0_u6_u3_n152 ) );
  NAND2_X1 u0_u6_u3_U64 (.A2( u0_u6_u3_n101 ) , .ZN( u0_u6_u3_n114 ) , .A1( u0_u6_u3_n96 ) );
  NAND2_X1 u0_u6_u3_U65 (.ZN( u0_u6_u3_n107 ) , .A1( u0_u6_u3_n97 ) , .A2( u0_u6_u3_n99 ) );
  NAND2_X1 u0_u6_u3_U66 (.A2( u0_u6_u3_n100 ) , .A1( u0_u6_u3_n104 ) , .ZN( u0_u6_u3_n113 ) );
  NAND2_X1 u0_u6_u3_U67 (.A1( u0_u6_u3_n104 ) , .ZN( u0_u6_u3_n153 ) , .A2( u0_u6_u3_n97 ) );
  NAND2_X1 u0_u6_u3_U68 (.A2( u0_u6_u3_n103 ) , .A1( u0_u6_u3_n104 ) , .ZN( u0_u6_u3_n130 ) );
  NAND2_X1 u0_u6_u3_U69 (.A2( u0_u6_u3_n103 ) , .ZN( u0_u6_u3_n144 ) , .A1( u0_u6_u3_n96 ) );
  OAI22_X1 u0_u6_u3_U7 (.B2( u0_u6_u3_n147 ) , .A2( u0_u6_u3_n148 ) , .ZN( u0_u6_u3_n160 ) , .B1( u0_u6_u3_n165 ) , .A1( u0_u6_u3_n168 ) );
  NAND2_X1 u0_u6_u3_U70 (.A1( u0_u6_u3_n102 ) , .A2( u0_u6_u3_n103 ) , .ZN( u0_u6_u3_n108 ) );
  NOR2_X1 u0_u6_u3_U71 (.A2( u0_u6_X_19 ) , .A1( u0_u6_X_20 ) , .ZN( u0_u6_u3_n99 ) );
  NOR2_X1 u0_u6_u3_U72 (.A2( u0_u6_X_21 ) , .A1( u0_u6_X_24 ) , .ZN( u0_u6_u3_n103 ) );
  NOR2_X1 u0_u6_u3_U73 (.A2( u0_u6_X_24 ) , .A1( u0_u6_u3_n171 ) , .ZN( u0_u6_u3_n97 ) );
  NOR2_X1 u0_u6_u3_U74 (.A2( u0_u6_X_23 ) , .ZN( u0_u6_u3_n141 ) , .A1( u0_u6_u3_n166 ) );
  NOR2_X1 u0_u6_u3_U75 (.A2( u0_u6_X_19 ) , .A1( u0_u6_u3_n172 ) , .ZN( u0_u6_u3_n96 ) );
  NAND2_X1 u0_u6_u3_U76 (.A1( u0_u6_X_22 ) , .A2( u0_u6_X_23 ) , .ZN( u0_u6_u3_n154 ) );
  NAND2_X1 u0_u6_u3_U77 (.A1( u0_u6_X_23 ) , .ZN( u0_u6_u3_n149 ) , .A2( u0_u6_u3_n166 ) );
  NOR2_X1 u0_u6_u3_U78 (.A2( u0_u6_X_22 ) , .A1( u0_u6_X_23 ) , .ZN( u0_u6_u3_n121 ) );
  AND2_X1 u0_u6_u3_U79 (.A1( u0_u6_X_24 ) , .ZN( u0_u6_u3_n101 ) , .A2( u0_u6_u3_n171 ) );
  AND3_X1 u0_u6_u3_U8 (.A3( u0_u6_u3_n144 ) , .A2( u0_u6_u3_n145 ) , .A1( u0_u6_u3_n146 ) , .ZN( u0_u6_u3_n147 ) );
  AND2_X1 u0_u6_u3_U80 (.A1( u0_u6_X_19 ) , .ZN( u0_u6_u3_n102 ) , .A2( u0_u6_u3_n172 ) );
  AND2_X1 u0_u6_u3_U81 (.A1( u0_u6_X_21 ) , .A2( u0_u6_X_24 ) , .ZN( u0_u6_u3_n100 ) );
  AND2_X1 u0_u6_u3_U82 (.A2( u0_u6_X_19 ) , .A1( u0_u6_X_20 ) , .ZN( u0_u6_u3_n104 ) );
  INV_X1 u0_u6_u3_U83 (.A( u0_u6_X_22 ) , .ZN( u0_u6_u3_n166 ) );
  INV_X1 u0_u6_u3_U84 (.A( u0_u6_X_21 ) , .ZN( u0_u6_u3_n171 ) );
  INV_X1 u0_u6_u3_U85 (.A( u0_u6_X_20 ) , .ZN( u0_u6_u3_n172 ) );
  NAND4_X1 u0_u6_u3_U86 (.ZN( u0_out6_26 ) , .A4( u0_u6_u3_n109 ) , .A3( u0_u6_u3_n110 ) , .A2( u0_u6_u3_n111 ) , .A1( u0_u6_u3_n173 ) );
  INV_X1 u0_u6_u3_U87 (.ZN( u0_u6_u3_n173 ) , .A( u0_u6_u3_n94 ) );
  OAI21_X1 u0_u6_u3_U88 (.ZN( u0_u6_u3_n111 ) , .B2( u0_u6_u3_n117 ) , .A( u0_u6_u3_n133 ) , .B1( u0_u6_u3_n176 ) );
  NAND4_X1 u0_u6_u3_U89 (.ZN( u0_out6_20 ) , .A4( u0_u6_u3_n122 ) , .A3( u0_u6_u3_n123 ) , .A1( u0_u6_u3_n175 ) , .A2( u0_u6_u3_n180 ) );
  INV_X1 u0_u6_u3_U9 (.A( u0_u6_u3_n143 ) , .ZN( u0_u6_u3_n168 ) );
  INV_X1 u0_u6_u3_U90 (.A( u0_u6_u3_n126 ) , .ZN( u0_u6_u3_n180 ) );
  INV_X1 u0_u6_u3_U91 (.A( u0_u6_u3_n112 ) , .ZN( u0_u6_u3_n175 ) );
  NAND4_X1 u0_u6_u3_U92 (.ZN( u0_out6_1 ) , .A4( u0_u6_u3_n161 ) , .A3( u0_u6_u3_n162 ) , .A2( u0_u6_u3_n163 ) , .A1( u0_u6_u3_n185 ) );
  NAND2_X1 u0_u6_u3_U93 (.ZN( u0_u6_u3_n163 ) , .A2( u0_u6_u3_n170 ) , .A1( u0_u6_u3_n176 ) );
  AOI22_X1 u0_u6_u3_U94 (.B2( u0_u6_u3_n140 ) , .B1( u0_u6_u3_n141 ) , .A2( u0_u6_u3_n142 ) , .ZN( u0_u6_u3_n162 ) , .A1( u0_u6_u3_n177 ) );
  OR4_X1 u0_u6_u3_U95 (.ZN( u0_out6_10 ) , .A4( u0_u6_u3_n136 ) , .A3( u0_u6_u3_n137 ) , .A1( u0_u6_u3_n138 ) , .A2( u0_u6_u3_n139 ) );
  OAI222_X1 u0_u6_u3_U96 (.C1( u0_u6_u3_n128 ) , .ZN( u0_u6_u3_n137 ) , .B1( u0_u6_u3_n148 ) , .A2( u0_u6_u3_n150 ) , .B2( u0_u6_u3_n154 ) , .C2( u0_u6_u3_n164 ) , .A1( u0_u6_u3_n167 ) );
  OAI221_X1 u0_u6_u3_U97 (.A( u0_u6_u3_n134 ) , .B2( u0_u6_u3_n135 ) , .ZN( u0_u6_u3_n136 ) , .C1( u0_u6_u3_n149 ) , .B1( u0_u6_u3_n151 ) , .C2( u0_u6_u3_n183 ) );
  NAND3_X1 u0_u6_u3_U98 (.A1( u0_u6_u3_n114 ) , .ZN( u0_u6_u3_n115 ) , .A2( u0_u6_u3_n145 ) , .A3( u0_u6_u3_n153 ) );
  NAND3_X1 u0_u6_u3_U99 (.ZN( u0_u6_u3_n129 ) , .A2( u0_u6_u3_n144 ) , .A1( u0_u6_u3_n153 ) , .A3( u0_u6_u3_n182 ) );
  INV_X1 u0_u6_u5_U10 (.A( u0_u6_u5_n121 ) , .ZN( u0_u6_u5_n177 ) );
  NOR3_X1 u0_u6_u5_U100 (.A3( u0_u6_u5_n141 ) , .A1( u0_u6_u5_n142 ) , .ZN( u0_u6_u5_n143 ) , .A2( u0_u6_u5_n191 ) );
  NAND4_X1 u0_u6_u5_U101 (.ZN( u0_out6_4 ) , .A4( u0_u6_u5_n112 ) , .A2( u0_u6_u5_n113 ) , .A1( u0_u6_u5_n114 ) , .A3( u0_u6_u5_n195 ) );
  AOI211_X1 u0_u6_u5_U102 (.A( u0_u6_u5_n110 ) , .C1( u0_u6_u5_n111 ) , .ZN( u0_u6_u5_n112 ) , .B( u0_u6_u5_n118 ) , .C2( u0_u6_u5_n177 ) );
  AOI222_X1 u0_u6_u5_U103 (.ZN( u0_u6_u5_n113 ) , .A1( u0_u6_u5_n131 ) , .C1( u0_u6_u5_n148 ) , .B2( u0_u6_u5_n174 ) , .C2( u0_u6_u5_n178 ) , .A2( u0_u6_u5_n179 ) , .B1( u0_u6_u5_n99 ) );
  NAND3_X1 u0_u6_u5_U104 (.A2( u0_u6_u5_n154 ) , .A3( u0_u6_u5_n158 ) , .A1( u0_u6_u5_n161 ) , .ZN( u0_u6_u5_n99 ) );
  NOR2_X1 u0_u6_u5_U11 (.ZN( u0_u6_u5_n160 ) , .A2( u0_u6_u5_n173 ) , .A1( u0_u6_u5_n177 ) );
  INV_X1 u0_u6_u5_U12 (.A( u0_u6_u5_n150 ) , .ZN( u0_u6_u5_n174 ) );
  AOI21_X1 u0_u6_u5_U13 (.A( u0_u6_u5_n160 ) , .B2( u0_u6_u5_n161 ) , .ZN( u0_u6_u5_n162 ) , .B1( u0_u6_u5_n192 ) );
  INV_X1 u0_u6_u5_U14 (.A( u0_u6_u5_n159 ) , .ZN( u0_u6_u5_n192 ) );
  AOI21_X1 u0_u6_u5_U15 (.A( u0_u6_u5_n156 ) , .B2( u0_u6_u5_n157 ) , .B1( u0_u6_u5_n158 ) , .ZN( u0_u6_u5_n163 ) );
  AOI21_X1 u0_u6_u5_U16 (.B2( u0_u6_u5_n139 ) , .B1( u0_u6_u5_n140 ) , .ZN( u0_u6_u5_n141 ) , .A( u0_u6_u5_n150 ) );
  OAI21_X1 u0_u6_u5_U17 (.A( u0_u6_u5_n133 ) , .B2( u0_u6_u5_n134 ) , .B1( u0_u6_u5_n135 ) , .ZN( u0_u6_u5_n142 ) );
  OAI21_X1 u0_u6_u5_U18 (.ZN( u0_u6_u5_n133 ) , .B2( u0_u6_u5_n147 ) , .A( u0_u6_u5_n173 ) , .B1( u0_u6_u5_n188 ) );
  NAND2_X1 u0_u6_u5_U19 (.A2( u0_u6_u5_n119 ) , .A1( u0_u6_u5_n123 ) , .ZN( u0_u6_u5_n137 ) );
  INV_X1 u0_u6_u5_U20 (.A( u0_u6_u5_n155 ) , .ZN( u0_u6_u5_n194 ) );
  NAND2_X1 u0_u6_u5_U21 (.A1( u0_u6_u5_n121 ) , .ZN( u0_u6_u5_n132 ) , .A2( u0_u6_u5_n172 ) );
  NAND2_X1 u0_u6_u5_U22 (.A2( u0_u6_u5_n122 ) , .ZN( u0_u6_u5_n136 ) , .A1( u0_u6_u5_n154 ) );
  NAND2_X1 u0_u6_u5_U23 (.A2( u0_u6_u5_n119 ) , .A1( u0_u6_u5_n120 ) , .ZN( u0_u6_u5_n159 ) );
  INV_X1 u0_u6_u5_U24 (.A( u0_u6_u5_n156 ) , .ZN( u0_u6_u5_n175 ) );
  INV_X1 u0_u6_u5_U25 (.A( u0_u6_u5_n158 ) , .ZN( u0_u6_u5_n188 ) );
  INV_X1 u0_u6_u5_U26 (.A( u0_u6_u5_n152 ) , .ZN( u0_u6_u5_n179 ) );
  INV_X1 u0_u6_u5_U27 (.A( u0_u6_u5_n140 ) , .ZN( u0_u6_u5_n182 ) );
  INV_X1 u0_u6_u5_U28 (.A( u0_u6_u5_n151 ) , .ZN( u0_u6_u5_n183 ) );
  INV_X1 u0_u6_u5_U29 (.A( u0_u6_u5_n123 ) , .ZN( u0_u6_u5_n185 ) );
  NOR2_X1 u0_u6_u5_U3 (.ZN( u0_u6_u5_n134 ) , .A1( u0_u6_u5_n183 ) , .A2( u0_u6_u5_n190 ) );
  INV_X1 u0_u6_u5_U30 (.A( u0_u6_u5_n161 ) , .ZN( u0_u6_u5_n184 ) );
  INV_X1 u0_u6_u5_U31 (.A( u0_u6_u5_n139 ) , .ZN( u0_u6_u5_n189 ) );
  INV_X1 u0_u6_u5_U32 (.A( u0_u6_u5_n157 ) , .ZN( u0_u6_u5_n190 ) );
  INV_X1 u0_u6_u5_U33 (.A( u0_u6_u5_n120 ) , .ZN( u0_u6_u5_n193 ) );
  NAND2_X1 u0_u6_u5_U34 (.ZN( u0_u6_u5_n111 ) , .A1( u0_u6_u5_n140 ) , .A2( u0_u6_u5_n155 ) );
  INV_X1 u0_u6_u5_U35 (.A( u0_u6_u5_n117 ) , .ZN( u0_u6_u5_n196 ) );
  OAI221_X1 u0_u6_u5_U36 (.A( u0_u6_u5_n116 ) , .ZN( u0_u6_u5_n117 ) , .B2( u0_u6_u5_n119 ) , .C1( u0_u6_u5_n153 ) , .C2( u0_u6_u5_n158 ) , .B1( u0_u6_u5_n172 ) );
  AOI222_X1 u0_u6_u5_U37 (.ZN( u0_u6_u5_n116 ) , .B2( u0_u6_u5_n145 ) , .C1( u0_u6_u5_n148 ) , .A2( u0_u6_u5_n174 ) , .C2( u0_u6_u5_n177 ) , .B1( u0_u6_u5_n187 ) , .A1( u0_u6_u5_n193 ) );
  INV_X1 u0_u6_u5_U38 (.A( u0_u6_u5_n115 ) , .ZN( u0_u6_u5_n187 ) );
  NOR2_X1 u0_u6_u5_U39 (.ZN( u0_u6_u5_n100 ) , .A1( u0_u6_u5_n170 ) , .A2( u0_u6_u5_n180 ) );
  INV_X1 u0_u6_u5_U4 (.A( u0_u6_u5_n138 ) , .ZN( u0_u6_u5_n191 ) );
  AOI22_X1 u0_u6_u5_U40 (.B2( u0_u6_u5_n131 ) , .A2( u0_u6_u5_n146 ) , .ZN( u0_u6_u5_n169 ) , .B1( u0_u6_u5_n174 ) , .A1( u0_u6_u5_n185 ) );
  NOR2_X1 u0_u6_u5_U41 (.A1( u0_u6_u5_n146 ) , .ZN( u0_u6_u5_n150 ) , .A2( u0_u6_u5_n173 ) );
  AOI21_X1 u0_u6_u5_U42 (.A( u0_u6_u5_n118 ) , .B2( u0_u6_u5_n145 ) , .ZN( u0_u6_u5_n168 ) , .B1( u0_u6_u5_n186 ) );
  INV_X1 u0_u6_u5_U43 (.A( u0_u6_u5_n122 ) , .ZN( u0_u6_u5_n186 ) );
  NOR2_X1 u0_u6_u5_U44 (.A1( u0_u6_u5_n146 ) , .ZN( u0_u6_u5_n152 ) , .A2( u0_u6_u5_n176 ) );
  NOR2_X1 u0_u6_u5_U45 (.A1( u0_u6_u5_n115 ) , .ZN( u0_u6_u5_n118 ) , .A2( u0_u6_u5_n153 ) );
  NOR2_X1 u0_u6_u5_U46 (.A2( u0_u6_u5_n145 ) , .ZN( u0_u6_u5_n156 ) , .A1( u0_u6_u5_n174 ) );
  NOR2_X1 u0_u6_u5_U47 (.ZN( u0_u6_u5_n121 ) , .A2( u0_u6_u5_n145 ) , .A1( u0_u6_u5_n176 ) );
  AOI22_X1 u0_u6_u5_U48 (.ZN( u0_u6_u5_n114 ) , .A2( u0_u6_u5_n137 ) , .A1( u0_u6_u5_n145 ) , .B2( u0_u6_u5_n175 ) , .B1( u0_u6_u5_n193 ) );
  OAI211_X1 u0_u6_u5_U49 (.B( u0_u6_u5_n124 ) , .A( u0_u6_u5_n125 ) , .C2( u0_u6_u5_n126 ) , .C1( u0_u6_u5_n127 ) , .ZN( u0_u6_u5_n128 ) );
  OAI21_X1 u0_u6_u5_U5 (.B2( u0_u6_u5_n136 ) , .B1( u0_u6_u5_n137 ) , .ZN( u0_u6_u5_n138 ) , .A( u0_u6_u5_n177 ) );
  NOR3_X1 u0_u6_u5_U50 (.ZN( u0_u6_u5_n127 ) , .A1( u0_u6_u5_n136 ) , .A3( u0_u6_u5_n148 ) , .A2( u0_u6_u5_n182 ) );
  OAI21_X1 u0_u6_u5_U51 (.ZN( u0_u6_u5_n124 ) , .A( u0_u6_u5_n177 ) , .B2( u0_u6_u5_n183 ) , .B1( u0_u6_u5_n189 ) );
  OAI21_X1 u0_u6_u5_U52 (.ZN( u0_u6_u5_n125 ) , .A( u0_u6_u5_n174 ) , .B2( u0_u6_u5_n185 ) , .B1( u0_u6_u5_n190 ) );
  AOI21_X1 u0_u6_u5_U53 (.A( u0_u6_u5_n153 ) , .B2( u0_u6_u5_n154 ) , .B1( u0_u6_u5_n155 ) , .ZN( u0_u6_u5_n164 ) );
  AOI21_X1 u0_u6_u5_U54 (.ZN( u0_u6_u5_n110 ) , .B1( u0_u6_u5_n122 ) , .B2( u0_u6_u5_n139 ) , .A( u0_u6_u5_n153 ) );
  INV_X1 u0_u6_u5_U55 (.A( u0_u6_u5_n153 ) , .ZN( u0_u6_u5_n176 ) );
  INV_X1 u0_u6_u5_U56 (.A( u0_u6_u5_n126 ) , .ZN( u0_u6_u5_n173 ) );
  AND2_X1 u0_u6_u5_U57 (.A2( u0_u6_u5_n104 ) , .A1( u0_u6_u5_n107 ) , .ZN( u0_u6_u5_n147 ) );
  AND2_X1 u0_u6_u5_U58 (.A2( u0_u6_u5_n104 ) , .A1( u0_u6_u5_n108 ) , .ZN( u0_u6_u5_n148 ) );
  NAND2_X1 u0_u6_u5_U59 (.A1( u0_u6_u5_n105 ) , .A2( u0_u6_u5_n106 ) , .ZN( u0_u6_u5_n158 ) );
  INV_X1 u0_u6_u5_U6 (.A( u0_u6_u5_n135 ) , .ZN( u0_u6_u5_n178 ) );
  NAND2_X1 u0_u6_u5_U60 (.A2( u0_u6_u5_n108 ) , .A1( u0_u6_u5_n109 ) , .ZN( u0_u6_u5_n139 ) );
  NAND2_X1 u0_u6_u5_U61 (.A1( u0_u6_u5_n106 ) , .A2( u0_u6_u5_n108 ) , .ZN( u0_u6_u5_n119 ) );
  NAND2_X1 u0_u6_u5_U62 (.A2( u0_u6_u5_n103 ) , .A1( u0_u6_u5_n105 ) , .ZN( u0_u6_u5_n140 ) );
  NAND2_X1 u0_u6_u5_U63 (.A2( u0_u6_u5_n104 ) , .A1( u0_u6_u5_n105 ) , .ZN( u0_u6_u5_n155 ) );
  NAND2_X1 u0_u6_u5_U64 (.A2( u0_u6_u5_n106 ) , .A1( u0_u6_u5_n107 ) , .ZN( u0_u6_u5_n122 ) );
  NAND2_X1 u0_u6_u5_U65 (.A2( u0_u6_u5_n100 ) , .A1( u0_u6_u5_n106 ) , .ZN( u0_u6_u5_n115 ) );
  NAND2_X1 u0_u6_u5_U66 (.A2( u0_u6_u5_n100 ) , .A1( u0_u6_u5_n103 ) , .ZN( u0_u6_u5_n161 ) );
  NAND2_X1 u0_u6_u5_U67 (.A1( u0_u6_u5_n105 ) , .A2( u0_u6_u5_n109 ) , .ZN( u0_u6_u5_n154 ) );
  INV_X1 u0_u6_u5_U68 (.A( u0_u6_u5_n146 ) , .ZN( u0_u6_u5_n172 ) );
  NAND2_X1 u0_u6_u5_U69 (.A1( u0_u6_u5_n103 ) , .A2( u0_u6_u5_n108 ) , .ZN( u0_u6_u5_n123 ) );
  OAI22_X1 u0_u6_u5_U7 (.B2( u0_u6_u5_n149 ) , .B1( u0_u6_u5_n150 ) , .A2( u0_u6_u5_n151 ) , .A1( u0_u6_u5_n152 ) , .ZN( u0_u6_u5_n165 ) );
  NAND2_X1 u0_u6_u5_U70 (.A2( u0_u6_u5_n103 ) , .A1( u0_u6_u5_n107 ) , .ZN( u0_u6_u5_n151 ) );
  NAND2_X1 u0_u6_u5_U71 (.A2( u0_u6_u5_n107 ) , .A1( u0_u6_u5_n109 ) , .ZN( u0_u6_u5_n120 ) );
  NAND2_X1 u0_u6_u5_U72 (.A2( u0_u6_u5_n100 ) , .A1( u0_u6_u5_n109 ) , .ZN( u0_u6_u5_n157 ) );
  AND2_X1 u0_u6_u5_U73 (.A2( u0_u6_u5_n100 ) , .A1( u0_u6_u5_n104 ) , .ZN( u0_u6_u5_n131 ) );
  INV_X1 u0_u6_u5_U74 (.A( u0_u6_u5_n102 ) , .ZN( u0_u6_u5_n195 ) );
  OAI221_X1 u0_u6_u5_U75 (.A( u0_u6_u5_n101 ) , .ZN( u0_u6_u5_n102 ) , .C2( u0_u6_u5_n115 ) , .C1( u0_u6_u5_n126 ) , .B1( u0_u6_u5_n134 ) , .B2( u0_u6_u5_n160 ) );
  OAI21_X1 u0_u6_u5_U76 (.ZN( u0_u6_u5_n101 ) , .B1( u0_u6_u5_n137 ) , .A( u0_u6_u5_n146 ) , .B2( u0_u6_u5_n147 ) );
  NOR2_X1 u0_u6_u5_U77 (.A2( u0_u6_X_34 ) , .A1( u0_u6_X_35 ) , .ZN( u0_u6_u5_n145 ) );
  NOR2_X1 u0_u6_u5_U78 (.A2( u0_u6_X_34 ) , .ZN( u0_u6_u5_n146 ) , .A1( u0_u6_u5_n171 ) );
  NOR2_X1 u0_u6_u5_U79 (.A2( u0_u6_X_31 ) , .A1( u0_u6_X_32 ) , .ZN( u0_u6_u5_n103 ) );
  NOR3_X1 u0_u6_u5_U8 (.A2( u0_u6_u5_n147 ) , .A1( u0_u6_u5_n148 ) , .ZN( u0_u6_u5_n149 ) , .A3( u0_u6_u5_n194 ) );
  NOR2_X1 u0_u6_u5_U80 (.A2( u0_u6_X_36 ) , .ZN( u0_u6_u5_n105 ) , .A1( u0_u6_u5_n180 ) );
  NOR2_X1 u0_u6_u5_U81 (.A2( u0_u6_X_33 ) , .ZN( u0_u6_u5_n108 ) , .A1( u0_u6_u5_n170 ) );
  NOR2_X1 u0_u6_u5_U82 (.A2( u0_u6_X_33 ) , .A1( u0_u6_X_36 ) , .ZN( u0_u6_u5_n107 ) );
  NOR2_X1 u0_u6_u5_U83 (.A2( u0_u6_X_31 ) , .ZN( u0_u6_u5_n104 ) , .A1( u0_u6_u5_n181 ) );
  NAND2_X1 u0_u6_u5_U84 (.A2( u0_u6_X_34 ) , .A1( u0_u6_X_35 ) , .ZN( u0_u6_u5_n153 ) );
  NAND2_X1 u0_u6_u5_U85 (.A1( u0_u6_X_34 ) , .ZN( u0_u6_u5_n126 ) , .A2( u0_u6_u5_n171 ) );
  AND2_X1 u0_u6_u5_U86 (.A1( u0_u6_X_31 ) , .A2( u0_u6_X_32 ) , .ZN( u0_u6_u5_n106 ) );
  AND2_X1 u0_u6_u5_U87 (.A1( u0_u6_X_31 ) , .ZN( u0_u6_u5_n109 ) , .A2( u0_u6_u5_n181 ) );
  INV_X1 u0_u6_u5_U88 (.A( u0_u6_X_33 ) , .ZN( u0_u6_u5_n180 ) );
  INV_X1 u0_u6_u5_U89 (.A( u0_u6_X_35 ) , .ZN( u0_u6_u5_n171 ) );
  NOR2_X1 u0_u6_u5_U9 (.ZN( u0_u6_u5_n135 ) , .A1( u0_u6_u5_n173 ) , .A2( u0_u6_u5_n176 ) );
  INV_X1 u0_u6_u5_U90 (.A( u0_u6_X_36 ) , .ZN( u0_u6_u5_n170 ) );
  INV_X1 u0_u6_u5_U91 (.A( u0_u6_X_32 ) , .ZN( u0_u6_u5_n181 ) );
  NAND4_X1 u0_u6_u5_U92 (.ZN( u0_out6_29 ) , .A4( u0_u6_u5_n129 ) , .A3( u0_u6_u5_n130 ) , .A2( u0_u6_u5_n168 ) , .A1( u0_u6_u5_n196 ) );
  AOI221_X1 u0_u6_u5_U93 (.A( u0_u6_u5_n128 ) , .ZN( u0_u6_u5_n129 ) , .C2( u0_u6_u5_n132 ) , .B2( u0_u6_u5_n159 ) , .B1( u0_u6_u5_n176 ) , .C1( u0_u6_u5_n184 ) );
  AOI222_X1 u0_u6_u5_U94 (.ZN( u0_u6_u5_n130 ) , .A2( u0_u6_u5_n146 ) , .B1( u0_u6_u5_n147 ) , .C2( u0_u6_u5_n175 ) , .B2( u0_u6_u5_n179 ) , .A1( u0_u6_u5_n188 ) , .C1( u0_u6_u5_n194 ) );
  NAND4_X1 u0_u6_u5_U95 (.ZN( u0_out6_19 ) , .A4( u0_u6_u5_n166 ) , .A3( u0_u6_u5_n167 ) , .A2( u0_u6_u5_n168 ) , .A1( u0_u6_u5_n169 ) );
  AOI22_X1 u0_u6_u5_U96 (.B2( u0_u6_u5_n145 ) , .A2( u0_u6_u5_n146 ) , .ZN( u0_u6_u5_n167 ) , .B1( u0_u6_u5_n182 ) , .A1( u0_u6_u5_n189 ) );
  NOR4_X1 u0_u6_u5_U97 (.A4( u0_u6_u5_n162 ) , .A3( u0_u6_u5_n163 ) , .A2( u0_u6_u5_n164 ) , .A1( u0_u6_u5_n165 ) , .ZN( u0_u6_u5_n166 ) );
  NAND4_X1 u0_u6_u5_U98 (.ZN( u0_out6_11 ) , .A4( u0_u6_u5_n143 ) , .A3( u0_u6_u5_n144 ) , .A2( u0_u6_u5_n169 ) , .A1( u0_u6_u5_n196 ) );
  AOI22_X1 u0_u6_u5_U99 (.A2( u0_u6_u5_n132 ) , .ZN( u0_u6_u5_n144 ) , .B2( u0_u6_u5_n145 ) , .B1( u0_u6_u5_n184 ) , .A1( u0_u6_u5_n194 ) );
  XOR2_X1 u0_u7_U2 (.B( u0_K8_8 ) , .A( u0_R6_5 ) , .Z( u0_u7_X_8 ) );
  XOR2_X1 u0_u7_U3 (.B( u0_K8_7 ) , .A( u0_R6_4 ) , .Z( u0_u7_X_7 ) );
  XOR2_X1 u0_u7_U33 (.B( u0_K8_24 ) , .A( u0_R6_17 ) , .Z( u0_u7_X_24 ) );
  XOR2_X1 u0_u7_U36 (.B( u0_K8_21 ) , .A( u0_R6_14 ) , .Z( u0_u7_X_21 ) );
  XOR2_X1 u0_u7_U37 (.B( u0_K8_20 ) , .A( u0_R6_13 ) , .Z( u0_u7_X_20 ) );
  XOR2_X1 u0_u7_U39 (.B( u0_K8_19 ) , .A( u0_R6_12 ) , .Z( u0_u7_X_19 ) );
  XOR2_X1 u0_u7_U4 (.B( u0_K8_6 ) , .A( u0_R6_5 ) , .Z( u0_u7_X_6 ) );
  XOR2_X1 u0_u7_U40 (.B( u0_K8_18 ) , .A( u0_R6_13 ) , .Z( u0_u7_X_18 ) );
  XOR2_X1 u0_u7_U41 (.B( u0_K8_17 ) , .A( u0_R6_12 ) , .Z( u0_u7_X_17 ) );
  XOR2_X1 u0_u7_U42 (.B( u0_K8_16 ) , .A( u0_R6_11 ) , .Z( u0_u7_X_16 ) );
  XOR2_X1 u0_u7_U43 (.B( u0_K8_15 ) , .A( u0_R6_10 ) , .Z( u0_u7_X_15 ) );
  XOR2_X1 u0_u7_U44 (.B( u0_K8_14 ) , .A( u0_R6_9 ) , .Z( u0_u7_X_14 ) );
  XOR2_X1 u0_u7_U45 (.B( u0_K8_13 ) , .A( u0_R6_8 ) , .Z( u0_u7_X_13 ) );
  XOR2_X1 u0_u7_U46 (.B( u0_K8_12 ) , .A( u0_R6_9 ) , .Z( u0_u7_X_12 ) );
  XOR2_X1 u0_u7_U47 (.B( u0_K8_11 ) , .A( u0_R6_8 ) , .Z( u0_u7_X_11 ) );
  XOR2_X1 u0_u7_U48 (.B( u0_K8_10 ) , .A( u0_R6_7 ) , .Z( u0_u7_X_10 ) );
  XOR2_X1 u0_u7_U5 (.B( u0_K8_5 ) , .A( u0_R6_4 ) , .Z( u0_u7_X_5 ) );
  AND3_X1 u0_u7_u0_U10 (.A2( u0_u7_u0_n112 ) , .ZN( u0_u7_u0_n127 ) , .A3( u0_u7_u0_n130 ) , .A1( u0_u7_u0_n148 ) );
  NAND2_X1 u0_u7_u0_U11 (.ZN( u0_u7_u0_n113 ) , .A1( u0_u7_u0_n139 ) , .A2( u0_u7_u0_n149 ) );
  AND2_X1 u0_u7_u0_U12 (.ZN( u0_u7_u0_n107 ) , .A1( u0_u7_u0_n130 ) , .A2( u0_u7_u0_n140 ) );
  AND2_X1 u0_u7_u0_U13 (.A2( u0_u7_u0_n129 ) , .A1( u0_u7_u0_n130 ) , .ZN( u0_u7_u0_n151 ) );
  AND2_X1 u0_u7_u0_U14 (.A1( u0_u7_u0_n108 ) , .A2( u0_u7_u0_n125 ) , .ZN( u0_u7_u0_n145 ) );
  INV_X1 u0_u7_u0_U15 (.A( u0_u7_u0_n143 ) , .ZN( u0_u7_u0_n173 ) );
  NOR2_X1 u0_u7_u0_U16 (.A2( u0_u7_u0_n136 ) , .ZN( u0_u7_u0_n147 ) , .A1( u0_u7_u0_n160 ) );
  INV_X1 u0_u7_u0_U17 (.ZN( u0_u7_u0_n172 ) , .A( u0_u7_u0_n88 ) );
  OAI222_X1 u0_u7_u0_U18 (.C1( u0_u7_u0_n108 ) , .A1( u0_u7_u0_n125 ) , .B2( u0_u7_u0_n128 ) , .B1( u0_u7_u0_n144 ) , .A2( u0_u7_u0_n158 ) , .C2( u0_u7_u0_n161 ) , .ZN( u0_u7_u0_n88 ) );
  NOR2_X1 u0_u7_u0_U19 (.A1( u0_u7_u0_n163 ) , .A2( u0_u7_u0_n164 ) , .ZN( u0_u7_u0_n95 ) );
  AOI21_X1 u0_u7_u0_U20 (.B1( u0_u7_u0_n103 ) , .ZN( u0_u7_u0_n132 ) , .A( u0_u7_u0_n165 ) , .B2( u0_u7_u0_n93 ) );
  INV_X1 u0_u7_u0_U21 (.A( u0_u7_u0_n142 ) , .ZN( u0_u7_u0_n165 ) );
  OAI22_X1 u0_u7_u0_U22 (.B1( u0_u7_u0_n125 ) , .ZN( u0_u7_u0_n126 ) , .A1( u0_u7_u0_n138 ) , .A2( u0_u7_u0_n146 ) , .B2( u0_u7_u0_n147 ) );
  OAI22_X1 u0_u7_u0_U23 (.B1( u0_u7_u0_n131 ) , .A1( u0_u7_u0_n144 ) , .B2( u0_u7_u0_n147 ) , .A2( u0_u7_u0_n90 ) , .ZN( u0_u7_u0_n91 ) );
  AND3_X1 u0_u7_u0_U24 (.A3( u0_u7_u0_n121 ) , .A2( u0_u7_u0_n125 ) , .A1( u0_u7_u0_n148 ) , .ZN( u0_u7_u0_n90 ) );
  NAND2_X1 u0_u7_u0_U25 (.A1( u0_u7_u0_n100 ) , .A2( u0_u7_u0_n103 ) , .ZN( u0_u7_u0_n125 ) );
  INV_X1 u0_u7_u0_U26 (.A( u0_u7_u0_n136 ) , .ZN( u0_u7_u0_n161 ) );
  AOI22_X1 u0_u7_u0_U27 (.B2( u0_u7_u0_n109 ) , .A2( u0_u7_u0_n110 ) , .ZN( u0_u7_u0_n111 ) , .B1( u0_u7_u0_n118 ) , .A1( u0_u7_u0_n160 ) );
  NAND2_X1 u0_u7_u0_U28 (.A1( u0_u7_u0_n100 ) , .ZN( u0_u7_u0_n129 ) , .A2( u0_u7_u0_n95 ) );
  INV_X1 u0_u7_u0_U29 (.A( u0_u7_u0_n118 ) , .ZN( u0_u7_u0_n158 ) );
  INV_X1 u0_u7_u0_U3 (.A( u0_u7_u0_n113 ) , .ZN( u0_u7_u0_n166 ) );
  AOI21_X1 u0_u7_u0_U30 (.ZN( u0_u7_u0_n104 ) , .B1( u0_u7_u0_n107 ) , .B2( u0_u7_u0_n141 ) , .A( u0_u7_u0_n144 ) );
  AOI21_X1 u0_u7_u0_U31 (.B1( u0_u7_u0_n127 ) , .B2( u0_u7_u0_n129 ) , .A( u0_u7_u0_n138 ) , .ZN( u0_u7_u0_n96 ) );
  AOI21_X1 u0_u7_u0_U32 (.ZN( u0_u7_u0_n116 ) , .B2( u0_u7_u0_n142 ) , .A( u0_u7_u0_n144 ) , .B1( u0_u7_u0_n166 ) );
  NOR2_X1 u0_u7_u0_U33 (.A1( u0_u7_u0_n120 ) , .ZN( u0_u7_u0_n143 ) , .A2( u0_u7_u0_n167 ) );
  OAI221_X1 u0_u7_u0_U34 (.C1( u0_u7_u0_n112 ) , .ZN( u0_u7_u0_n120 ) , .B1( u0_u7_u0_n138 ) , .B2( u0_u7_u0_n141 ) , .C2( u0_u7_u0_n147 ) , .A( u0_u7_u0_n172 ) );
  AOI211_X1 u0_u7_u0_U35 (.B( u0_u7_u0_n115 ) , .A( u0_u7_u0_n116 ) , .C2( u0_u7_u0_n117 ) , .C1( u0_u7_u0_n118 ) , .ZN( u0_u7_u0_n119 ) );
  NAND2_X1 u0_u7_u0_U36 (.A2( u0_u7_u0_n100 ) , .A1( u0_u7_u0_n101 ) , .ZN( u0_u7_u0_n139 ) );
  NAND2_X1 u0_u7_u0_U37 (.A2( u0_u7_u0_n100 ) , .ZN( u0_u7_u0_n131 ) , .A1( u0_u7_u0_n92 ) );
  NAND2_X1 u0_u7_u0_U38 (.A1( u0_u7_u0_n101 ) , .A2( u0_u7_u0_n102 ) , .ZN( u0_u7_u0_n150 ) );
  INV_X1 u0_u7_u0_U39 (.A( u0_u7_u0_n138 ) , .ZN( u0_u7_u0_n160 ) );
  AOI21_X1 u0_u7_u0_U4 (.B1( u0_u7_u0_n114 ) , .ZN( u0_u7_u0_n115 ) , .B2( u0_u7_u0_n129 ) , .A( u0_u7_u0_n161 ) );
  NAND2_X1 u0_u7_u0_U40 (.A1( u0_u7_u0_n102 ) , .ZN( u0_u7_u0_n128 ) , .A2( u0_u7_u0_n95 ) );
  NAND2_X1 u0_u7_u0_U41 (.ZN( u0_u7_u0_n148 ) , .A1( u0_u7_u0_n93 ) , .A2( u0_u7_u0_n95 ) );
  NAND2_X1 u0_u7_u0_U42 (.A2( u0_u7_u0_n102 ) , .A1( u0_u7_u0_n103 ) , .ZN( u0_u7_u0_n149 ) );
  NAND2_X1 u0_u7_u0_U43 (.A2( u0_u7_u0_n102 ) , .ZN( u0_u7_u0_n114 ) , .A1( u0_u7_u0_n92 ) );
  NAND2_X1 u0_u7_u0_U44 (.A2( u0_u7_u0_n101 ) , .ZN( u0_u7_u0_n121 ) , .A1( u0_u7_u0_n93 ) );
  NAND2_X1 u0_u7_u0_U45 (.ZN( u0_u7_u0_n112 ) , .A2( u0_u7_u0_n92 ) , .A1( u0_u7_u0_n93 ) );
  OR3_X1 u0_u7_u0_U46 (.A3( u0_u7_u0_n152 ) , .A2( u0_u7_u0_n153 ) , .A1( u0_u7_u0_n154 ) , .ZN( u0_u7_u0_n155 ) );
  AOI21_X1 u0_u7_u0_U47 (.A( u0_u7_u0_n144 ) , .B2( u0_u7_u0_n145 ) , .B1( u0_u7_u0_n146 ) , .ZN( u0_u7_u0_n154 ) );
  AOI21_X1 u0_u7_u0_U48 (.B2( u0_u7_u0_n150 ) , .B1( u0_u7_u0_n151 ) , .ZN( u0_u7_u0_n152 ) , .A( u0_u7_u0_n158 ) );
  AOI21_X1 u0_u7_u0_U49 (.A( u0_u7_u0_n147 ) , .B2( u0_u7_u0_n148 ) , .B1( u0_u7_u0_n149 ) , .ZN( u0_u7_u0_n153 ) );
  AOI21_X1 u0_u7_u0_U5 (.B2( u0_u7_u0_n131 ) , .ZN( u0_u7_u0_n134 ) , .B1( u0_u7_u0_n151 ) , .A( u0_u7_u0_n158 ) );
  INV_X1 u0_u7_u0_U50 (.ZN( u0_u7_u0_n171 ) , .A( u0_u7_u0_n99 ) );
  OAI211_X1 u0_u7_u0_U51 (.C2( u0_u7_u0_n140 ) , .C1( u0_u7_u0_n161 ) , .A( u0_u7_u0_n169 ) , .B( u0_u7_u0_n98 ) , .ZN( u0_u7_u0_n99 ) );
  INV_X1 u0_u7_u0_U52 (.ZN( u0_u7_u0_n169 ) , .A( u0_u7_u0_n91 ) );
  AOI211_X1 u0_u7_u0_U53 (.C1( u0_u7_u0_n118 ) , .A( u0_u7_u0_n123 ) , .B( u0_u7_u0_n96 ) , .C2( u0_u7_u0_n97 ) , .ZN( u0_u7_u0_n98 ) );
  NOR2_X1 u0_u7_u0_U54 (.A2( u0_u7_X_4 ) , .A1( u0_u7_X_5 ) , .ZN( u0_u7_u0_n118 ) );
  NOR2_X1 u0_u7_u0_U55 (.A2( u0_u7_X_2 ) , .ZN( u0_u7_u0_n103 ) , .A1( u0_u7_u0_n164 ) );
  NOR2_X1 u0_u7_u0_U56 (.A2( u0_u7_X_1 ) , .A1( u0_u7_X_2 ) , .ZN( u0_u7_u0_n92 ) );
  NOR2_X1 u0_u7_u0_U57 (.A2( u0_u7_X_1 ) , .ZN( u0_u7_u0_n101 ) , .A1( u0_u7_u0_n163 ) );
  NAND2_X1 u0_u7_u0_U58 (.A2( u0_u7_X_4 ) , .A1( u0_u7_X_5 ) , .ZN( u0_u7_u0_n144 ) );
  NOR2_X1 u0_u7_u0_U59 (.A2( u0_u7_X_5 ) , .ZN( u0_u7_u0_n136 ) , .A1( u0_u7_u0_n159 ) );
  NOR2_X1 u0_u7_u0_U6 (.A1( u0_u7_u0_n108 ) , .ZN( u0_u7_u0_n123 ) , .A2( u0_u7_u0_n158 ) );
  NAND2_X1 u0_u7_u0_U60 (.A1( u0_u7_X_5 ) , .ZN( u0_u7_u0_n138 ) , .A2( u0_u7_u0_n159 ) );
  NOR2_X1 u0_u7_u0_U61 (.A2( u0_u7_X_3 ) , .A1( u0_u7_X_6 ) , .ZN( u0_u7_u0_n94 ) );
  AND2_X1 u0_u7_u0_U62 (.A2( u0_u7_X_3 ) , .A1( u0_u7_X_6 ) , .ZN( u0_u7_u0_n102 ) );
  AND2_X1 u0_u7_u0_U63 (.A1( u0_u7_X_6 ) , .A2( u0_u7_u0_n162 ) , .ZN( u0_u7_u0_n93 ) );
  INV_X1 u0_u7_u0_U64 (.A( u0_u7_X_4 ) , .ZN( u0_u7_u0_n159 ) );
  INV_X1 u0_u7_u0_U65 (.A( u0_u7_X_1 ) , .ZN( u0_u7_u0_n164 ) );
  INV_X1 u0_u7_u0_U66 (.A( u0_u7_X_2 ) , .ZN( u0_u7_u0_n163 ) );
  INV_X1 u0_u7_u0_U67 (.A( u0_u7_u0_n126 ) , .ZN( u0_u7_u0_n168 ) );
  AOI211_X1 u0_u7_u0_U68 (.B( u0_u7_u0_n133 ) , .A( u0_u7_u0_n134 ) , .C2( u0_u7_u0_n135 ) , .C1( u0_u7_u0_n136 ) , .ZN( u0_u7_u0_n137 ) );
  OR4_X1 u0_u7_u0_U69 (.ZN( u0_out7_17 ) , .A4( u0_u7_u0_n122 ) , .A2( u0_u7_u0_n123 ) , .A1( u0_u7_u0_n124 ) , .A3( u0_u7_u0_n170 ) );
  OAI21_X1 u0_u7_u0_U7 (.B1( u0_u7_u0_n150 ) , .B2( u0_u7_u0_n158 ) , .A( u0_u7_u0_n172 ) , .ZN( u0_u7_u0_n89 ) );
  AOI21_X1 u0_u7_u0_U70 (.B2( u0_u7_u0_n107 ) , .ZN( u0_u7_u0_n124 ) , .B1( u0_u7_u0_n128 ) , .A( u0_u7_u0_n161 ) );
  INV_X1 u0_u7_u0_U71 (.A( u0_u7_u0_n111 ) , .ZN( u0_u7_u0_n170 ) );
  OR4_X1 u0_u7_u0_U72 (.ZN( u0_out7_31 ) , .A4( u0_u7_u0_n155 ) , .A2( u0_u7_u0_n156 ) , .A1( u0_u7_u0_n157 ) , .A3( u0_u7_u0_n173 ) );
  AOI21_X1 u0_u7_u0_U73 (.A( u0_u7_u0_n138 ) , .B2( u0_u7_u0_n139 ) , .B1( u0_u7_u0_n140 ) , .ZN( u0_u7_u0_n157 ) );
  AOI21_X1 u0_u7_u0_U74 (.B2( u0_u7_u0_n141 ) , .B1( u0_u7_u0_n142 ) , .ZN( u0_u7_u0_n156 ) , .A( u0_u7_u0_n161 ) );
  INV_X1 u0_u7_u0_U75 (.ZN( u0_u7_u0_n174 ) , .A( u0_u7_u0_n89 ) );
  AOI211_X1 u0_u7_u0_U76 (.B( u0_u7_u0_n104 ) , .A( u0_u7_u0_n105 ) , .ZN( u0_u7_u0_n106 ) , .C2( u0_u7_u0_n113 ) , .C1( u0_u7_u0_n160 ) );
  OAI221_X1 u0_u7_u0_U77 (.C1( u0_u7_u0_n121 ) , .ZN( u0_u7_u0_n122 ) , .B2( u0_u7_u0_n127 ) , .A( u0_u7_u0_n143 ) , .B1( u0_u7_u0_n144 ) , .C2( u0_u7_u0_n147 ) );
  NOR2_X1 u0_u7_u0_U78 (.A2( u0_u7_X_6 ) , .ZN( u0_u7_u0_n100 ) , .A1( u0_u7_u0_n162 ) );
  INV_X1 u0_u7_u0_U79 (.A( u0_u7_X_3 ) , .ZN( u0_u7_u0_n162 ) );
  AND2_X1 u0_u7_u0_U8 (.A1( u0_u7_u0_n114 ) , .A2( u0_u7_u0_n121 ) , .ZN( u0_u7_u0_n146 ) );
  AOI21_X1 u0_u7_u0_U80 (.B1( u0_u7_u0_n132 ) , .ZN( u0_u7_u0_n133 ) , .A( u0_u7_u0_n144 ) , .B2( u0_u7_u0_n166 ) );
  OAI22_X1 u0_u7_u0_U81 (.ZN( u0_u7_u0_n105 ) , .A2( u0_u7_u0_n132 ) , .B1( u0_u7_u0_n146 ) , .A1( u0_u7_u0_n147 ) , .B2( u0_u7_u0_n161 ) );
  NAND2_X1 u0_u7_u0_U82 (.ZN( u0_u7_u0_n110 ) , .A2( u0_u7_u0_n132 ) , .A1( u0_u7_u0_n145 ) );
  INV_X1 u0_u7_u0_U83 (.A( u0_u7_u0_n119 ) , .ZN( u0_u7_u0_n167 ) );
  NAND2_X1 u0_u7_u0_U84 (.A2( u0_u7_u0_n103 ) , .ZN( u0_u7_u0_n140 ) , .A1( u0_u7_u0_n94 ) );
  NAND2_X1 u0_u7_u0_U85 (.A1( u0_u7_u0_n101 ) , .ZN( u0_u7_u0_n130 ) , .A2( u0_u7_u0_n94 ) );
  NAND2_X1 u0_u7_u0_U86 (.ZN( u0_u7_u0_n108 ) , .A1( u0_u7_u0_n92 ) , .A2( u0_u7_u0_n94 ) );
  NAND2_X1 u0_u7_u0_U87 (.ZN( u0_u7_u0_n142 ) , .A1( u0_u7_u0_n94 ) , .A2( u0_u7_u0_n95 ) );
  NAND3_X1 u0_u7_u0_U88 (.ZN( u0_out7_23 ) , .A3( u0_u7_u0_n137 ) , .A1( u0_u7_u0_n168 ) , .A2( u0_u7_u0_n171 ) );
  NAND3_X1 u0_u7_u0_U89 (.A3( u0_u7_u0_n127 ) , .A2( u0_u7_u0_n128 ) , .ZN( u0_u7_u0_n135 ) , .A1( u0_u7_u0_n150 ) );
  AND2_X1 u0_u7_u0_U9 (.A1( u0_u7_u0_n131 ) , .ZN( u0_u7_u0_n141 ) , .A2( u0_u7_u0_n150 ) );
  NAND3_X1 u0_u7_u0_U90 (.ZN( u0_u7_u0_n117 ) , .A3( u0_u7_u0_n132 ) , .A2( u0_u7_u0_n139 ) , .A1( u0_u7_u0_n148 ) );
  NAND3_X1 u0_u7_u0_U91 (.ZN( u0_u7_u0_n109 ) , .A2( u0_u7_u0_n114 ) , .A3( u0_u7_u0_n140 ) , .A1( u0_u7_u0_n149 ) );
  NAND3_X1 u0_u7_u0_U92 (.ZN( u0_out7_9 ) , .A3( u0_u7_u0_n106 ) , .A2( u0_u7_u0_n171 ) , .A1( u0_u7_u0_n174 ) );
  NAND3_X1 u0_u7_u0_U93 (.A2( u0_u7_u0_n128 ) , .A1( u0_u7_u0_n132 ) , .A3( u0_u7_u0_n146 ) , .ZN( u0_u7_u0_n97 ) );
  AOI21_X1 u0_u7_u1_U10 (.B2( u0_u7_u1_n155 ) , .B1( u0_u7_u1_n156 ) , .ZN( u0_u7_u1_n157 ) , .A( u0_u7_u1_n174 ) );
  NAND3_X1 u0_u7_u1_U100 (.ZN( u0_u7_u1_n113 ) , .A1( u0_u7_u1_n120 ) , .A3( u0_u7_u1_n133 ) , .A2( u0_u7_u1_n155 ) );
  NAND2_X1 u0_u7_u1_U11 (.ZN( u0_u7_u1_n140 ) , .A2( u0_u7_u1_n150 ) , .A1( u0_u7_u1_n155 ) );
  NAND2_X1 u0_u7_u1_U12 (.A1( u0_u7_u1_n131 ) , .ZN( u0_u7_u1_n147 ) , .A2( u0_u7_u1_n153 ) );
  AOI22_X1 u0_u7_u1_U13 (.B2( u0_u7_u1_n136 ) , .A2( u0_u7_u1_n137 ) , .ZN( u0_u7_u1_n143 ) , .A1( u0_u7_u1_n171 ) , .B1( u0_u7_u1_n173 ) );
  INV_X1 u0_u7_u1_U14 (.A( u0_u7_u1_n147 ) , .ZN( u0_u7_u1_n181 ) );
  INV_X1 u0_u7_u1_U15 (.A( u0_u7_u1_n139 ) , .ZN( u0_u7_u1_n174 ) );
  OR4_X1 u0_u7_u1_U16 (.A4( u0_u7_u1_n106 ) , .A3( u0_u7_u1_n107 ) , .ZN( u0_u7_u1_n108 ) , .A1( u0_u7_u1_n117 ) , .A2( u0_u7_u1_n184 ) );
  AOI21_X1 u0_u7_u1_U17 (.ZN( u0_u7_u1_n106 ) , .A( u0_u7_u1_n112 ) , .B1( u0_u7_u1_n154 ) , .B2( u0_u7_u1_n156 ) );
  AOI21_X1 u0_u7_u1_U18 (.ZN( u0_u7_u1_n107 ) , .B1( u0_u7_u1_n134 ) , .B2( u0_u7_u1_n149 ) , .A( u0_u7_u1_n174 ) );
  INV_X1 u0_u7_u1_U19 (.A( u0_u7_u1_n101 ) , .ZN( u0_u7_u1_n184 ) );
  INV_X1 u0_u7_u1_U20 (.A( u0_u7_u1_n112 ) , .ZN( u0_u7_u1_n171 ) );
  NAND2_X1 u0_u7_u1_U21 (.ZN( u0_u7_u1_n141 ) , .A1( u0_u7_u1_n153 ) , .A2( u0_u7_u1_n156 ) );
  AND2_X1 u0_u7_u1_U22 (.A1( u0_u7_u1_n123 ) , .ZN( u0_u7_u1_n134 ) , .A2( u0_u7_u1_n161 ) );
  NAND2_X1 u0_u7_u1_U23 (.A2( u0_u7_u1_n115 ) , .A1( u0_u7_u1_n116 ) , .ZN( u0_u7_u1_n148 ) );
  NAND2_X1 u0_u7_u1_U24 (.A2( u0_u7_u1_n133 ) , .A1( u0_u7_u1_n135 ) , .ZN( u0_u7_u1_n159 ) );
  NAND2_X1 u0_u7_u1_U25 (.A2( u0_u7_u1_n115 ) , .A1( u0_u7_u1_n120 ) , .ZN( u0_u7_u1_n132 ) );
  INV_X1 u0_u7_u1_U26 (.A( u0_u7_u1_n154 ) , .ZN( u0_u7_u1_n178 ) );
  INV_X1 u0_u7_u1_U27 (.A( u0_u7_u1_n151 ) , .ZN( u0_u7_u1_n183 ) );
  AND2_X1 u0_u7_u1_U28 (.A1( u0_u7_u1_n129 ) , .A2( u0_u7_u1_n133 ) , .ZN( u0_u7_u1_n149 ) );
  INV_X1 u0_u7_u1_U29 (.A( u0_u7_u1_n131 ) , .ZN( u0_u7_u1_n180 ) );
  INV_X1 u0_u7_u1_U3 (.A( u0_u7_u1_n159 ) , .ZN( u0_u7_u1_n182 ) );
  OAI221_X1 u0_u7_u1_U30 (.A( u0_u7_u1_n119 ) , .C2( u0_u7_u1_n129 ) , .ZN( u0_u7_u1_n138 ) , .B2( u0_u7_u1_n152 ) , .C1( u0_u7_u1_n174 ) , .B1( u0_u7_u1_n187 ) );
  INV_X1 u0_u7_u1_U31 (.A( u0_u7_u1_n148 ) , .ZN( u0_u7_u1_n187 ) );
  AOI211_X1 u0_u7_u1_U32 (.B( u0_u7_u1_n117 ) , .A( u0_u7_u1_n118 ) , .ZN( u0_u7_u1_n119 ) , .C2( u0_u7_u1_n146 ) , .C1( u0_u7_u1_n159 ) );
  NOR2_X1 u0_u7_u1_U33 (.A1( u0_u7_u1_n168 ) , .A2( u0_u7_u1_n176 ) , .ZN( u0_u7_u1_n98 ) );
  AOI211_X1 u0_u7_u1_U34 (.B( u0_u7_u1_n162 ) , .A( u0_u7_u1_n163 ) , .C2( u0_u7_u1_n164 ) , .ZN( u0_u7_u1_n165 ) , .C1( u0_u7_u1_n171 ) );
  AOI21_X1 u0_u7_u1_U35 (.A( u0_u7_u1_n160 ) , .B2( u0_u7_u1_n161 ) , .ZN( u0_u7_u1_n162 ) , .B1( u0_u7_u1_n182 ) );
  OR2_X1 u0_u7_u1_U36 (.A2( u0_u7_u1_n157 ) , .A1( u0_u7_u1_n158 ) , .ZN( u0_u7_u1_n163 ) );
  NAND2_X1 u0_u7_u1_U37 (.A1( u0_u7_u1_n128 ) , .ZN( u0_u7_u1_n146 ) , .A2( u0_u7_u1_n160 ) );
  NAND2_X1 u0_u7_u1_U38 (.A2( u0_u7_u1_n112 ) , .ZN( u0_u7_u1_n139 ) , .A1( u0_u7_u1_n152 ) );
  NAND2_X1 u0_u7_u1_U39 (.A1( u0_u7_u1_n105 ) , .ZN( u0_u7_u1_n156 ) , .A2( u0_u7_u1_n99 ) );
  AOI221_X1 u0_u7_u1_U4 (.A( u0_u7_u1_n138 ) , .C2( u0_u7_u1_n139 ) , .C1( u0_u7_u1_n140 ) , .B2( u0_u7_u1_n141 ) , .ZN( u0_u7_u1_n142 ) , .B1( u0_u7_u1_n175 ) );
  AOI221_X1 u0_u7_u1_U40 (.B1( u0_u7_u1_n140 ) , .ZN( u0_u7_u1_n167 ) , .B2( u0_u7_u1_n172 ) , .C2( u0_u7_u1_n175 ) , .C1( u0_u7_u1_n178 ) , .A( u0_u7_u1_n188 ) );
  INV_X1 u0_u7_u1_U41 (.ZN( u0_u7_u1_n188 ) , .A( u0_u7_u1_n97 ) );
  AOI211_X1 u0_u7_u1_U42 (.A( u0_u7_u1_n118 ) , .C1( u0_u7_u1_n132 ) , .C2( u0_u7_u1_n139 ) , .B( u0_u7_u1_n96 ) , .ZN( u0_u7_u1_n97 ) );
  AOI21_X1 u0_u7_u1_U43 (.B2( u0_u7_u1_n121 ) , .B1( u0_u7_u1_n135 ) , .A( u0_u7_u1_n152 ) , .ZN( u0_u7_u1_n96 ) );
  NOR2_X1 u0_u7_u1_U44 (.ZN( u0_u7_u1_n117 ) , .A1( u0_u7_u1_n121 ) , .A2( u0_u7_u1_n160 ) );
  OAI21_X1 u0_u7_u1_U45 (.B2( u0_u7_u1_n123 ) , .ZN( u0_u7_u1_n145 ) , .B1( u0_u7_u1_n160 ) , .A( u0_u7_u1_n185 ) );
  INV_X1 u0_u7_u1_U46 (.A( u0_u7_u1_n122 ) , .ZN( u0_u7_u1_n185 ) );
  AOI21_X1 u0_u7_u1_U47 (.B2( u0_u7_u1_n120 ) , .B1( u0_u7_u1_n121 ) , .ZN( u0_u7_u1_n122 ) , .A( u0_u7_u1_n128 ) );
  AOI21_X1 u0_u7_u1_U48 (.A( u0_u7_u1_n128 ) , .B2( u0_u7_u1_n129 ) , .ZN( u0_u7_u1_n130 ) , .B1( u0_u7_u1_n150 ) );
  NAND2_X1 u0_u7_u1_U49 (.ZN( u0_u7_u1_n112 ) , .A1( u0_u7_u1_n169 ) , .A2( u0_u7_u1_n170 ) );
  AOI211_X1 u0_u7_u1_U5 (.ZN( u0_u7_u1_n124 ) , .A( u0_u7_u1_n138 ) , .C2( u0_u7_u1_n139 ) , .B( u0_u7_u1_n145 ) , .C1( u0_u7_u1_n147 ) );
  NAND2_X1 u0_u7_u1_U50 (.ZN( u0_u7_u1_n129 ) , .A2( u0_u7_u1_n95 ) , .A1( u0_u7_u1_n98 ) );
  NAND2_X1 u0_u7_u1_U51 (.A1( u0_u7_u1_n102 ) , .ZN( u0_u7_u1_n154 ) , .A2( u0_u7_u1_n99 ) );
  NAND2_X1 u0_u7_u1_U52 (.A2( u0_u7_u1_n100 ) , .ZN( u0_u7_u1_n135 ) , .A1( u0_u7_u1_n99 ) );
  AOI21_X1 u0_u7_u1_U53 (.A( u0_u7_u1_n152 ) , .B2( u0_u7_u1_n153 ) , .B1( u0_u7_u1_n154 ) , .ZN( u0_u7_u1_n158 ) );
  INV_X1 u0_u7_u1_U54 (.A( u0_u7_u1_n160 ) , .ZN( u0_u7_u1_n175 ) );
  NAND2_X1 u0_u7_u1_U55 (.A1( u0_u7_u1_n100 ) , .ZN( u0_u7_u1_n116 ) , .A2( u0_u7_u1_n95 ) );
  NAND2_X1 u0_u7_u1_U56 (.A1( u0_u7_u1_n102 ) , .ZN( u0_u7_u1_n131 ) , .A2( u0_u7_u1_n95 ) );
  NAND2_X1 u0_u7_u1_U57 (.A2( u0_u7_u1_n104 ) , .ZN( u0_u7_u1_n121 ) , .A1( u0_u7_u1_n98 ) );
  NAND2_X1 u0_u7_u1_U58 (.A1( u0_u7_u1_n103 ) , .ZN( u0_u7_u1_n153 ) , .A2( u0_u7_u1_n98 ) );
  NAND2_X1 u0_u7_u1_U59 (.A2( u0_u7_u1_n104 ) , .A1( u0_u7_u1_n105 ) , .ZN( u0_u7_u1_n133 ) );
  AOI22_X1 u0_u7_u1_U6 (.B2( u0_u7_u1_n113 ) , .A2( u0_u7_u1_n114 ) , .ZN( u0_u7_u1_n125 ) , .A1( u0_u7_u1_n171 ) , .B1( u0_u7_u1_n173 ) );
  NAND2_X1 u0_u7_u1_U60 (.ZN( u0_u7_u1_n150 ) , .A2( u0_u7_u1_n98 ) , .A1( u0_u7_u1_n99 ) );
  NAND2_X1 u0_u7_u1_U61 (.A1( u0_u7_u1_n105 ) , .ZN( u0_u7_u1_n155 ) , .A2( u0_u7_u1_n95 ) );
  OAI21_X1 u0_u7_u1_U62 (.ZN( u0_u7_u1_n109 ) , .B1( u0_u7_u1_n129 ) , .B2( u0_u7_u1_n160 ) , .A( u0_u7_u1_n167 ) );
  NAND2_X1 u0_u7_u1_U63 (.A2( u0_u7_u1_n100 ) , .A1( u0_u7_u1_n103 ) , .ZN( u0_u7_u1_n120 ) );
  NAND2_X1 u0_u7_u1_U64 (.A1( u0_u7_u1_n102 ) , .A2( u0_u7_u1_n104 ) , .ZN( u0_u7_u1_n115 ) );
  NAND2_X1 u0_u7_u1_U65 (.A2( u0_u7_u1_n100 ) , .A1( u0_u7_u1_n104 ) , .ZN( u0_u7_u1_n151 ) );
  NAND2_X1 u0_u7_u1_U66 (.A2( u0_u7_u1_n103 ) , .A1( u0_u7_u1_n105 ) , .ZN( u0_u7_u1_n161 ) );
  INV_X1 u0_u7_u1_U67 (.A( u0_u7_u1_n152 ) , .ZN( u0_u7_u1_n173 ) );
  INV_X1 u0_u7_u1_U68 (.A( u0_u7_u1_n128 ) , .ZN( u0_u7_u1_n172 ) );
  NAND2_X1 u0_u7_u1_U69 (.A2( u0_u7_u1_n102 ) , .A1( u0_u7_u1_n103 ) , .ZN( u0_u7_u1_n123 ) );
  NAND2_X1 u0_u7_u1_U7 (.ZN( u0_u7_u1_n114 ) , .A1( u0_u7_u1_n134 ) , .A2( u0_u7_u1_n156 ) );
  NOR2_X1 u0_u7_u1_U70 (.A2( u0_u7_X_7 ) , .A1( u0_u7_X_8 ) , .ZN( u0_u7_u1_n95 ) );
  NOR2_X1 u0_u7_u1_U71 (.A1( u0_u7_X_12 ) , .A2( u0_u7_X_9 ) , .ZN( u0_u7_u1_n100 ) );
  NOR2_X1 u0_u7_u1_U72 (.A2( u0_u7_X_8 ) , .A1( u0_u7_u1_n177 ) , .ZN( u0_u7_u1_n99 ) );
  NOR2_X1 u0_u7_u1_U73 (.A2( u0_u7_X_12 ) , .ZN( u0_u7_u1_n102 ) , .A1( u0_u7_u1_n176 ) );
  NOR2_X1 u0_u7_u1_U74 (.A2( u0_u7_X_9 ) , .ZN( u0_u7_u1_n105 ) , .A1( u0_u7_u1_n168 ) );
  NAND2_X1 u0_u7_u1_U75 (.A1( u0_u7_X_10 ) , .ZN( u0_u7_u1_n160 ) , .A2( u0_u7_u1_n169 ) );
  NAND2_X1 u0_u7_u1_U76 (.A2( u0_u7_X_10 ) , .A1( u0_u7_X_11 ) , .ZN( u0_u7_u1_n152 ) );
  NAND2_X1 u0_u7_u1_U77 (.A1( u0_u7_X_11 ) , .ZN( u0_u7_u1_n128 ) , .A2( u0_u7_u1_n170 ) );
  AND2_X1 u0_u7_u1_U78 (.A2( u0_u7_X_7 ) , .A1( u0_u7_X_8 ) , .ZN( u0_u7_u1_n104 ) );
  AND2_X1 u0_u7_u1_U79 (.A1( u0_u7_X_8 ) , .ZN( u0_u7_u1_n103 ) , .A2( u0_u7_u1_n177 ) );
  NOR2_X1 u0_u7_u1_U8 (.A1( u0_u7_u1_n112 ) , .A2( u0_u7_u1_n116 ) , .ZN( u0_u7_u1_n118 ) );
  INV_X1 u0_u7_u1_U80 (.A( u0_u7_X_10 ) , .ZN( u0_u7_u1_n170 ) );
  INV_X1 u0_u7_u1_U81 (.A( u0_u7_X_9 ) , .ZN( u0_u7_u1_n176 ) );
  INV_X1 u0_u7_u1_U82 (.A( u0_u7_X_11 ) , .ZN( u0_u7_u1_n169 ) );
  INV_X1 u0_u7_u1_U83 (.A( u0_u7_X_12 ) , .ZN( u0_u7_u1_n168 ) );
  INV_X1 u0_u7_u1_U84 (.A( u0_u7_X_7 ) , .ZN( u0_u7_u1_n177 ) );
  NAND4_X1 u0_u7_u1_U85 (.ZN( u0_out7_28 ) , .A4( u0_u7_u1_n124 ) , .A3( u0_u7_u1_n125 ) , .A2( u0_u7_u1_n126 ) , .A1( u0_u7_u1_n127 ) );
  OAI21_X1 u0_u7_u1_U86 (.ZN( u0_u7_u1_n127 ) , .B2( u0_u7_u1_n139 ) , .B1( u0_u7_u1_n175 ) , .A( u0_u7_u1_n183 ) );
  OAI21_X1 u0_u7_u1_U87 (.ZN( u0_u7_u1_n126 ) , .B2( u0_u7_u1_n140 ) , .A( u0_u7_u1_n146 ) , .B1( u0_u7_u1_n178 ) );
  NAND4_X1 u0_u7_u1_U88 (.ZN( u0_out7_18 ) , .A4( u0_u7_u1_n165 ) , .A3( u0_u7_u1_n166 ) , .A1( u0_u7_u1_n167 ) , .A2( u0_u7_u1_n186 ) );
  AOI22_X1 u0_u7_u1_U89 (.B2( u0_u7_u1_n146 ) , .B1( u0_u7_u1_n147 ) , .A2( u0_u7_u1_n148 ) , .ZN( u0_u7_u1_n166 ) , .A1( u0_u7_u1_n172 ) );
  OAI21_X1 u0_u7_u1_U9 (.ZN( u0_u7_u1_n101 ) , .B1( u0_u7_u1_n141 ) , .A( u0_u7_u1_n146 ) , .B2( u0_u7_u1_n183 ) );
  INV_X1 u0_u7_u1_U90 (.A( u0_u7_u1_n145 ) , .ZN( u0_u7_u1_n186 ) );
  NAND4_X1 u0_u7_u1_U91 (.ZN( u0_out7_2 ) , .A4( u0_u7_u1_n142 ) , .A3( u0_u7_u1_n143 ) , .A2( u0_u7_u1_n144 ) , .A1( u0_u7_u1_n179 ) );
  OAI21_X1 u0_u7_u1_U92 (.B2( u0_u7_u1_n132 ) , .ZN( u0_u7_u1_n144 ) , .A( u0_u7_u1_n146 ) , .B1( u0_u7_u1_n180 ) );
  INV_X1 u0_u7_u1_U93 (.A( u0_u7_u1_n130 ) , .ZN( u0_u7_u1_n179 ) );
  OR4_X1 u0_u7_u1_U94 (.ZN( u0_out7_13 ) , .A4( u0_u7_u1_n108 ) , .A3( u0_u7_u1_n109 ) , .A2( u0_u7_u1_n110 ) , .A1( u0_u7_u1_n111 ) );
  AOI21_X1 u0_u7_u1_U95 (.ZN( u0_u7_u1_n111 ) , .A( u0_u7_u1_n128 ) , .B2( u0_u7_u1_n131 ) , .B1( u0_u7_u1_n135 ) );
  AOI21_X1 u0_u7_u1_U96 (.ZN( u0_u7_u1_n110 ) , .A( u0_u7_u1_n116 ) , .B1( u0_u7_u1_n152 ) , .B2( u0_u7_u1_n160 ) );
  NAND3_X1 u0_u7_u1_U97 (.A3( u0_u7_u1_n149 ) , .A2( u0_u7_u1_n150 ) , .A1( u0_u7_u1_n151 ) , .ZN( u0_u7_u1_n164 ) );
  NAND3_X1 u0_u7_u1_U98 (.A3( u0_u7_u1_n134 ) , .A2( u0_u7_u1_n135 ) , .ZN( u0_u7_u1_n136 ) , .A1( u0_u7_u1_n151 ) );
  NAND3_X1 u0_u7_u1_U99 (.A1( u0_u7_u1_n133 ) , .ZN( u0_u7_u1_n137 ) , .A2( u0_u7_u1_n154 ) , .A3( u0_u7_u1_n181 ) );
  OAI22_X1 u0_u7_u2_U10 (.ZN( u0_u7_u2_n109 ) , .A2( u0_u7_u2_n113 ) , .B2( u0_u7_u2_n133 ) , .B1( u0_u7_u2_n167 ) , .A1( u0_u7_u2_n168 ) );
  NAND3_X1 u0_u7_u2_U100 (.A2( u0_u7_u2_n100 ) , .A1( u0_u7_u2_n104 ) , .A3( u0_u7_u2_n138 ) , .ZN( u0_u7_u2_n98 ) );
  OAI22_X1 u0_u7_u2_U11 (.B1( u0_u7_u2_n151 ) , .A2( u0_u7_u2_n152 ) , .A1( u0_u7_u2_n153 ) , .ZN( u0_u7_u2_n160 ) , .B2( u0_u7_u2_n168 ) );
  NOR3_X1 u0_u7_u2_U12 (.A1( u0_u7_u2_n150 ) , .ZN( u0_u7_u2_n151 ) , .A3( u0_u7_u2_n175 ) , .A2( u0_u7_u2_n188 ) );
  AOI21_X1 u0_u7_u2_U13 (.ZN( u0_u7_u2_n144 ) , .B2( u0_u7_u2_n155 ) , .A( u0_u7_u2_n172 ) , .B1( u0_u7_u2_n185 ) );
  AOI21_X1 u0_u7_u2_U14 (.B2( u0_u7_u2_n143 ) , .ZN( u0_u7_u2_n145 ) , .B1( u0_u7_u2_n152 ) , .A( u0_u7_u2_n171 ) );
  AOI21_X1 u0_u7_u2_U15 (.B2( u0_u7_u2_n120 ) , .B1( u0_u7_u2_n121 ) , .ZN( u0_u7_u2_n126 ) , .A( u0_u7_u2_n167 ) );
  INV_X1 u0_u7_u2_U16 (.A( u0_u7_u2_n156 ) , .ZN( u0_u7_u2_n171 ) );
  INV_X1 u0_u7_u2_U17 (.A( u0_u7_u2_n120 ) , .ZN( u0_u7_u2_n188 ) );
  NAND2_X1 u0_u7_u2_U18 (.A2( u0_u7_u2_n122 ) , .ZN( u0_u7_u2_n150 ) , .A1( u0_u7_u2_n152 ) );
  INV_X1 u0_u7_u2_U19 (.A( u0_u7_u2_n153 ) , .ZN( u0_u7_u2_n170 ) );
  INV_X1 u0_u7_u2_U20 (.A( u0_u7_u2_n137 ) , .ZN( u0_u7_u2_n173 ) );
  NAND2_X1 u0_u7_u2_U21 (.A1( u0_u7_u2_n132 ) , .A2( u0_u7_u2_n139 ) , .ZN( u0_u7_u2_n157 ) );
  INV_X1 u0_u7_u2_U22 (.A( u0_u7_u2_n113 ) , .ZN( u0_u7_u2_n178 ) );
  INV_X1 u0_u7_u2_U23 (.A( u0_u7_u2_n139 ) , .ZN( u0_u7_u2_n175 ) );
  INV_X1 u0_u7_u2_U24 (.A( u0_u7_u2_n155 ) , .ZN( u0_u7_u2_n181 ) );
  INV_X1 u0_u7_u2_U25 (.A( u0_u7_u2_n119 ) , .ZN( u0_u7_u2_n177 ) );
  INV_X1 u0_u7_u2_U26 (.A( u0_u7_u2_n116 ) , .ZN( u0_u7_u2_n180 ) );
  INV_X1 u0_u7_u2_U27 (.A( u0_u7_u2_n131 ) , .ZN( u0_u7_u2_n179 ) );
  INV_X1 u0_u7_u2_U28 (.A( u0_u7_u2_n154 ) , .ZN( u0_u7_u2_n176 ) );
  NAND2_X1 u0_u7_u2_U29 (.A2( u0_u7_u2_n116 ) , .A1( u0_u7_u2_n117 ) , .ZN( u0_u7_u2_n118 ) );
  NOR2_X1 u0_u7_u2_U3 (.ZN( u0_u7_u2_n121 ) , .A2( u0_u7_u2_n177 ) , .A1( u0_u7_u2_n180 ) );
  INV_X1 u0_u7_u2_U30 (.A( u0_u7_u2_n132 ) , .ZN( u0_u7_u2_n182 ) );
  INV_X1 u0_u7_u2_U31 (.A( u0_u7_u2_n158 ) , .ZN( u0_u7_u2_n183 ) );
  OAI21_X1 u0_u7_u2_U32 (.A( u0_u7_u2_n156 ) , .B1( u0_u7_u2_n157 ) , .ZN( u0_u7_u2_n158 ) , .B2( u0_u7_u2_n179 ) );
  NOR2_X1 u0_u7_u2_U33 (.ZN( u0_u7_u2_n156 ) , .A1( u0_u7_u2_n166 ) , .A2( u0_u7_u2_n169 ) );
  NOR2_X1 u0_u7_u2_U34 (.A2( u0_u7_u2_n114 ) , .ZN( u0_u7_u2_n137 ) , .A1( u0_u7_u2_n140 ) );
  NOR2_X1 u0_u7_u2_U35 (.A2( u0_u7_u2_n138 ) , .ZN( u0_u7_u2_n153 ) , .A1( u0_u7_u2_n156 ) );
  AOI211_X1 u0_u7_u2_U36 (.ZN( u0_u7_u2_n130 ) , .C1( u0_u7_u2_n138 ) , .C2( u0_u7_u2_n179 ) , .B( u0_u7_u2_n96 ) , .A( u0_u7_u2_n97 ) );
  OAI22_X1 u0_u7_u2_U37 (.B1( u0_u7_u2_n133 ) , .A2( u0_u7_u2_n137 ) , .A1( u0_u7_u2_n152 ) , .B2( u0_u7_u2_n168 ) , .ZN( u0_u7_u2_n97 ) );
  OAI221_X1 u0_u7_u2_U38 (.B1( u0_u7_u2_n113 ) , .C1( u0_u7_u2_n132 ) , .A( u0_u7_u2_n149 ) , .B2( u0_u7_u2_n171 ) , .C2( u0_u7_u2_n172 ) , .ZN( u0_u7_u2_n96 ) );
  OAI221_X1 u0_u7_u2_U39 (.A( u0_u7_u2_n115 ) , .C2( u0_u7_u2_n123 ) , .B2( u0_u7_u2_n143 ) , .B1( u0_u7_u2_n153 ) , .ZN( u0_u7_u2_n163 ) , .C1( u0_u7_u2_n168 ) );
  INV_X1 u0_u7_u2_U4 (.A( u0_u7_u2_n134 ) , .ZN( u0_u7_u2_n185 ) );
  OAI21_X1 u0_u7_u2_U40 (.A( u0_u7_u2_n114 ) , .ZN( u0_u7_u2_n115 ) , .B1( u0_u7_u2_n176 ) , .B2( u0_u7_u2_n178 ) );
  OAI221_X1 u0_u7_u2_U41 (.A( u0_u7_u2_n135 ) , .B2( u0_u7_u2_n136 ) , .B1( u0_u7_u2_n137 ) , .ZN( u0_u7_u2_n162 ) , .C2( u0_u7_u2_n167 ) , .C1( u0_u7_u2_n185 ) );
  AND3_X1 u0_u7_u2_U42 (.A3( u0_u7_u2_n131 ) , .A2( u0_u7_u2_n132 ) , .A1( u0_u7_u2_n133 ) , .ZN( u0_u7_u2_n136 ) );
  AOI22_X1 u0_u7_u2_U43 (.ZN( u0_u7_u2_n135 ) , .B1( u0_u7_u2_n140 ) , .A1( u0_u7_u2_n156 ) , .B2( u0_u7_u2_n180 ) , .A2( u0_u7_u2_n188 ) );
  AOI21_X1 u0_u7_u2_U44 (.ZN( u0_u7_u2_n149 ) , .B1( u0_u7_u2_n173 ) , .B2( u0_u7_u2_n188 ) , .A( u0_u7_u2_n95 ) );
  AND3_X1 u0_u7_u2_U45 (.A2( u0_u7_u2_n100 ) , .A1( u0_u7_u2_n104 ) , .A3( u0_u7_u2_n156 ) , .ZN( u0_u7_u2_n95 ) );
  OAI21_X1 u0_u7_u2_U46 (.A( u0_u7_u2_n101 ) , .B2( u0_u7_u2_n121 ) , .B1( u0_u7_u2_n153 ) , .ZN( u0_u7_u2_n164 ) );
  NAND2_X1 u0_u7_u2_U47 (.A2( u0_u7_u2_n100 ) , .A1( u0_u7_u2_n107 ) , .ZN( u0_u7_u2_n155 ) );
  NAND2_X1 u0_u7_u2_U48 (.A2( u0_u7_u2_n105 ) , .A1( u0_u7_u2_n108 ) , .ZN( u0_u7_u2_n143 ) );
  NAND2_X1 u0_u7_u2_U49 (.A1( u0_u7_u2_n104 ) , .A2( u0_u7_u2_n106 ) , .ZN( u0_u7_u2_n152 ) );
  INV_X1 u0_u7_u2_U5 (.A( u0_u7_u2_n150 ) , .ZN( u0_u7_u2_n184 ) );
  NAND2_X1 u0_u7_u2_U50 (.A1( u0_u7_u2_n100 ) , .A2( u0_u7_u2_n105 ) , .ZN( u0_u7_u2_n132 ) );
  INV_X1 u0_u7_u2_U51 (.A( u0_u7_u2_n140 ) , .ZN( u0_u7_u2_n168 ) );
  INV_X1 u0_u7_u2_U52 (.A( u0_u7_u2_n138 ) , .ZN( u0_u7_u2_n167 ) );
  OAI21_X1 u0_u7_u2_U53 (.A( u0_u7_u2_n141 ) , .B2( u0_u7_u2_n142 ) , .ZN( u0_u7_u2_n146 ) , .B1( u0_u7_u2_n153 ) );
  OAI21_X1 u0_u7_u2_U54 (.A( u0_u7_u2_n140 ) , .ZN( u0_u7_u2_n141 ) , .B1( u0_u7_u2_n176 ) , .B2( u0_u7_u2_n177 ) );
  NOR3_X1 u0_u7_u2_U55 (.ZN( u0_u7_u2_n142 ) , .A3( u0_u7_u2_n175 ) , .A2( u0_u7_u2_n178 ) , .A1( u0_u7_u2_n181 ) );
  INV_X1 u0_u7_u2_U56 (.ZN( u0_u7_u2_n187 ) , .A( u0_u7_u2_n99 ) );
  OAI21_X1 u0_u7_u2_U57 (.B1( u0_u7_u2_n137 ) , .B2( u0_u7_u2_n143 ) , .A( u0_u7_u2_n98 ) , .ZN( u0_u7_u2_n99 ) );
  NAND2_X1 u0_u7_u2_U58 (.A1( u0_u7_u2_n102 ) , .A2( u0_u7_u2_n106 ) , .ZN( u0_u7_u2_n113 ) );
  NAND2_X1 u0_u7_u2_U59 (.A1( u0_u7_u2_n106 ) , .A2( u0_u7_u2_n107 ) , .ZN( u0_u7_u2_n131 ) );
  NOR4_X1 u0_u7_u2_U6 (.A4( u0_u7_u2_n124 ) , .A3( u0_u7_u2_n125 ) , .A2( u0_u7_u2_n126 ) , .A1( u0_u7_u2_n127 ) , .ZN( u0_u7_u2_n128 ) );
  NAND2_X1 u0_u7_u2_U60 (.A1( u0_u7_u2_n103 ) , .A2( u0_u7_u2_n107 ) , .ZN( u0_u7_u2_n139 ) );
  NAND2_X1 u0_u7_u2_U61 (.A1( u0_u7_u2_n103 ) , .A2( u0_u7_u2_n105 ) , .ZN( u0_u7_u2_n133 ) );
  NAND2_X1 u0_u7_u2_U62 (.A1( u0_u7_u2_n102 ) , .A2( u0_u7_u2_n103 ) , .ZN( u0_u7_u2_n154 ) );
  NAND2_X1 u0_u7_u2_U63 (.A2( u0_u7_u2_n103 ) , .A1( u0_u7_u2_n104 ) , .ZN( u0_u7_u2_n119 ) );
  NAND2_X1 u0_u7_u2_U64 (.A2( u0_u7_u2_n107 ) , .A1( u0_u7_u2_n108 ) , .ZN( u0_u7_u2_n123 ) );
  NAND2_X1 u0_u7_u2_U65 (.A1( u0_u7_u2_n104 ) , .A2( u0_u7_u2_n108 ) , .ZN( u0_u7_u2_n122 ) );
  INV_X1 u0_u7_u2_U66 (.A( u0_u7_u2_n114 ) , .ZN( u0_u7_u2_n172 ) );
  NAND2_X1 u0_u7_u2_U67 (.A2( u0_u7_u2_n100 ) , .A1( u0_u7_u2_n102 ) , .ZN( u0_u7_u2_n116 ) );
  NAND2_X1 u0_u7_u2_U68 (.A1( u0_u7_u2_n102 ) , .A2( u0_u7_u2_n108 ) , .ZN( u0_u7_u2_n120 ) );
  NAND2_X1 u0_u7_u2_U69 (.A2( u0_u7_u2_n105 ) , .A1( u0_u7_u2_n106 ) , .ZN( u0_u7_u2_n117 ) );
  AOI21_X1 u0_u7_u2_U7 (.B2( u0_u7_u2_n119 ) , .ZN( u0_u7_u2_n127 ) , .A( u0_u7_u2_n137 ) , .B1( u0_u7_u2_n155 ) );
  NOR2_X1 u0_u7_u2_U70 (.A2( u0_u7_X_16 ) , .ZN( u0_u7_u2_n140 ) , .A1( u0_u7_u2_n166 ) );
  NOR2_X1 u0_u7_u2_U71 (.A2( u0_u7_X_13 ) , .A1( u0_u7_X_14 ) , .ZN( u0_u7_u2_n100 ) );
  NOR2_X1 u0_u7_u2_U72 (.A2( u0_u7_X_16 ) , .A1( u0_u7_X_17 ) , .ZN( u0_u7_u2_n138 ) );
  NOR2_X1 u0_u7_u2_U73 (.A2( u0_u7_X_15 ) , .A1( u0_u7_X_18 ) , .ZN( u0_u7_u2_n104 ) );
  NOR2_X1 u0_u7_u2_U74 (.A2( u0_u7_X_14 ) , .ZN( u0_u7_u2_n103 ) , .A1( u0_u7_u2_n174 ) );
  NOR2_X1 u0_u7_u2_U75 (.A2( u0_u7_X_15 ) , .ZN( u0_u7_u2_n102 ) , .A1( u0_u7_u2_n165 ) );
  NOR2_X1 u0_u7_u2_U76 (.A2( u0_u7_X_17 ) , .ZN( u0_u7_u2_n114 ) , .A1( u0_u7_u2_n169 ) );
  AND2_X1 u0_u7_u2_U77 (.A1( u0_u7_X_15 ) , .ZN( u0_u7_u2_n105 ) , .A2( u0_u7_u2_n165 ) );
  AND2_X1 u0_u7_u2_U78 (.A2( u0_u7_X_15 ) , .A1( u0_u7_X_18 ) , .ZN( u0_u7_u2_n107 ) );
  AND2_X1 u0_u7_u2_U79 (.A1( u0_u7_X_14 ) , .ZN( u0_u7_u2_n106 ) , .A2( u0_u7_u2_n174 ) );
  AOI21_X1 u0_u7_u2_U8 (.ZN( u0_u7_u2_n124 ) , .B1( u0_u7_u2_n131 ) , .B2( u0_u7_u2_n143 ) , .A( u0_u7_u2_n172 ) );
  AND2_X1 u0_u7_u2_U80 (.A1( u0_u7_X_13 ) , .A2( u0_u7_X_14 ) , .ZN( u0_u7_u2_n108 ) );
  INV_X1 u0_u7_u2_U81 (.A( u0_u7_X_16 ) , .ZN( u0_u7_u2_n169 ) );
  INV_X1 u0_u7_u2_U82 (.A( u0_u7_X_17 ) , .ZN( u0_u7_u2_n166 ) );
  INV_X1 u0_u7_u2_U83 (.A( u0_u7_X_13 ) , .ZN( u0_u7_u2_n174 ) );
  INV_X1 u0_u7_u2_U84 (.A( u0_u7_X_18 ) , .ZN( u0_u7_u2_n165 ) );
  NAND4_X1 u0_u7_u2_U85 (.ZN( u0_out7_30 ) , .A4( u0_u7_u2_n147 ) , .A3( u0_u7_u2_n148 ) , .A2( u0_u7_u2_n149 ) , .A1( u0_u7_u2_n187 ) );
  NOR3_X1 u0_u7_u2_U86 (.A3( u0_u7_u2_n144 ) , .A2( u0_u7_u2_n145 ) , .A1( u0_u7_u2_n146 ) , .ZN( u0_u7_u2_n147 ) );
  AOI21_X1 u0_u7_u2_U87 (.B2( u0_u7_u2_n138 ) , .ZN( u0_u7_u2_n148 ) , .A( u0_u7_u2_n162 ) , .B1( u0_u7_u2_n182 ) );
  NAND4_X1 u0_u7_u2_U88 (.ZN( u0_out7_24 ) , .A4( u0_u7_u2_n111 ) , .A3( u0_u7_u2_n112 ) , .A1( u0_u7_u2_n130 ) , .A2( u0_u7_u2_n187 ) );
  AOI221_X1 u0_u7_u2_U89 (.A( u0_u7_u2_n109 ) , .B1( u0_u7_u2_n110 ) , .ZN( u0_u7_u2_n111 ) , .C1( u0_u7_u2_n134 ) , .C2( u0_u7_u2_n170 ) , .B2( u0_u7_u2_n173 ) );
  AOI21_X1 u0_u7_u2_U9 (.B2( u0_u7_u2_n123 ) , .ZN( u0_u7_u2_n125 ) , .A( u0_u7_u2_n171 ) , .B1( u0_u7_u2_n184 ) );
  AOI21_X1 u0_u7_u2_U90 (.ZN( u0_u7_u2_n112 ) , .B2( u0_u7_u2_n156 ) , .A( u0_u7_u2_n164 ) , .B1( u0_u7_u2_n181 ) );
  NAND4_X1 u0_u7_u2_U91 (.ZN( u0_out7_16 ) , .A4( u0_u7_u2_n128 ) , .A3( u0_u7_u2_n129 ) , .A1( u0_u7_u2_n130 ) , .A2( u0_u7_u2_n186 ) );
  AOI22_X1 u0_u7_u2_U92 (.A2( u0_u7_u2_n118 ) , .ZN( u0_u7_u2_n129 ) , .A1( u0_u7_u2_n140 ) , .B1( u0_u7_u2_n157 ) , .B2( u0_u7_u2_n170 ) );
  INV_X1 u0_u7_u2_U93 (.A( u0_u7_u2_n163 ) , .ZN( u0_u7_u2_n186 ) );
  OR4_X1 u0_u7_u2_U94 (.ZN( u0_out7_6 ) , .A4( u0_u7_u2_n161 ) , .A3( u0_u7_u2_n162 ) , .A2( u0_u7_u2_n163 ) , .A1( u0_u7_u2_n164 ) );
  OR3_X1 u0_u7_u2_U95 (.A2( u0_u7_u2_n159 ) , .A1( u0_u7_u2_n160 ) , .ZN( u0_u7_u2_n161 ) , .A3( u0_u7_u2_n183 ) );
  AOI21_X1 u0_u7_u2_U96 (.B2( u0_u7_u2_n154 ) , .B1( u0_u7_u2_n155 ) , .ZN( u0_u7_u2_n159 ) , .A( u0_u7_u2_n167 ) );
  NAND3_X1 u0_u7_u2_U97 (.A2( u0_u7_u2_n117 ) , .A1( u0_u7_u2_n122 ) , .A3( u0_u7_u2_n123 ) , .ZN( u0_u7_u2_n134 ) );
  NAND3_X1 u0_u7_u2_U98 (.ZN( u0_u7_u2_n110 ) , .A2( u0_u7_u2_n131 ) , .A3( u0_u7_u2_n139 ) , .A1( u0_u7_u2_n154 ) );
  NAND3_X1 u0_u7_u2_U99 (.A2( u0_u7_u2_n100 ) , .ZN( u0_u7_u2_n101 ) , .A1( u0_u7_u2_n104 ) , .A3( u0_u7_u2_n114 ) );
  OAI22_X1 u0_u7_u3_U10 (.B1( u0_u7_u3_n113 ) , .A2( u0_u7_u3_n135 ) , .A1( u0_u7_u3_n150 ) , .B2( u0_u7_u3_n164 ) , .ZN( u0_u7_u3_n98 ) );
  OAI211_X1 u0_u7_u3_U11 (.B( u0_u7_u3_n106 ) , .ZN( u0_u7_u3_n119 ) , .C2( u0_u7_u3_n128 ) , .C1( u0_u7_u3_n167 ) , .A( u0_u7_u3_n181 ) );
  AOI221_X1 u0_u7_u3_U12 (.C1( u0_u7_u3_n105 ) , .ZN( u0_u7_u3_n106 ) , .A( u0_u7_u3_n131 ) , .B2( u0_u7_u3_n132 ) , .C2( u0_u7_u3_n133 ) , .B1( u0_u7_u3_n169 ) );
  INV_X1 u0_u7_u3_U13 (.ZN( u0_u7_u3_n181 ) , .A( u0_u7_u3_n98 ) );
  NAND2_X1 u0_u7_u3_U14 (.ZN( u0_u7_u3_n105 ) , .A2( u0_u7_u3_n130 ) , .A1( u0_u7_u3_n155 ) );
  AOI22_X1 u0_u7_u3_U15 (.B1( u0_u7_u3_n115 ) , .A2( u0_u7_u3_n116 ) , .ZN( u0_u7_u3_n123 ) , .B2( u0_u7_u3_n133 ) , .A1( u0_u7_u3_n169 ) );
  NAND2_X1 u0_u7_u3_U16 (.ZN( u0_u7_u3_n116 ) , .A2( u0_u7_u3_n151 ) , .A1( u0_u7_u3_n182 ) );
  NOR2_X1 u0_u7_u3_U17 (.ZN( u0_u7_u3_n126 ) , .A2( u0_u7_u3_n150 ) , .A1( u0_u7_u3_n164 ) );
  AOI21_X1 u0_u7_u3_U18 (.ZN( u0_u7_u3_n112 ) , .B2( u0_u7_u3_n146 ) , .B1( u0_u7_u3_n155 ) , .A( u0_u7_u3_n167 ) );
  NAND2_X1 u0_u7_u3_U19 (.A1( u0_u7_u3_n135 ) , .ZN( u0_u7_u3_n142 ) , .A2( u0_u7_u3_n164 ) );
  NAND2_X1 u0_u7_u3_U20 (.ZN( u0_u7_u3_n132 ) , .A2( u0_u7_u3_n152 ) , .A1( u0_u7_u3_n156 ) );
  AND2_X1 u0_u7_u3_U21 (.A2( u0_u7_u3_n113 ) , .A1( u0_u7_u3_n114 ) , .ZN( u0_u7_u3_n151 ) );
  INV_X1 u0_u7_u3_U22 (.A( u0_u7_u3_n133 ) , .ZN( u0_u7_u3_n165 ) );
  INV_X1 u0_u7_u3_U23 (.A( u0_u7_u3_n135 ) , .ZN( u0_u7_u3_n170 ) );
  NAND2_X1 u0_u7_u3_U24 (.A1( u0_u7_u3_n107 ) , .A2( u0_u7_u3_n108 ) , .ZN( u0_u7_u3_n140 ) );
  NAND2_X1 u0_u7_u3_U25 (.ZN( u0_u7_u3_n117 ) , .A1( u0_u7_u3_n124 ) , .A2( u0_u7_u3_n148 ) );
  NAND2_X1 u0_u7_u3_U26 (.ZN( u0_u7_u3_n143 ) , .A1( u0_u7_u3_n165 ) , .A2( u0_u7_u3_n167 ) );
  INV_X1 u0_u7_u3_U27 (.A( u0_u7_u3_n130 ) , .ZN( u0_u7_u3_n177 ) );
  INV_X1 u0_u7_u3_U28 (.A( u0_u7_u3_n128 ) , .ZN( u0_u7_u3_n176 ) );
  INV_X1 u0_u7_u3_U29 (.A( u0_u7_u3_n155 ) , .ZN( u0_u7_u3_n174 ) );
  INV_X1 u0_u7_u3_U3 (.A( u0_u7_u3_n129 ) , .ZN( u0_u7_u3_n183 ) );
  INV_X1 u0_u7_u3_U30 (.A( u0_u7_u3_n139 ) , .ZN( u0_u7_u3_n185 ) );
  NOR2_X1 u0_u7_u3_U31 (.ZN( u0_u7_u3_n135 ) , .A2( u0_u7_u3_n141 ) , .A1( u0_u7_u3_n169 ) );
  OAI222_X1 u0_u7_u3_U32 (.C2( u0_u7_u3_n107 ) , .A2( u0_u7_u3_n108 ) , .B1( u0_u7_u3_n135 ) , .ZN( u0_u7_u3_n138 ) , .B2( u0_u7_u3_n146 ) , .C1( u0_u7_u3_n154 ) , .A1( u0_u7_u3_n164 ) );
  NOR4_X1 u0_u7_u3_U33 (.A4( u0_u7_u3_n157 ) , .A3( u0_u7_u3_n158 ) , .A2( u0_u7_u3_n159 ) , .A1( u0_u7_u3_n160 ) , .ZN( u0_u7_u3_n161 ) );
  AOI21_X1 u0_u7_u3_U34 (.B2( u0_u7_u3_n152 ) , .B1( u0_u7_u3_n153 ) , .ZN( u0_u7_u3_n158 ) , .A( u0_u7_u3_n164 ) );
  AOI21_X1 u0_u7_u3_U35 (.A( u0_u7_u3_n154 ) , .B2( u0_u7_u3_n155 ) , .B1( u0_u7_u3_n156 ) , .ZN( u0_u7_u3_n157 ) );
  AOI21_X1 u0_u7_u3_U36 (.A( u0_u7_u3_n149 ) , .B2( u0_u7_u3_n150 ) , .B1( u0_u7_u3_n151 ) , .ZN( u0_u7_u3_n159 ) );
  AOI211_X1 u0_u7_u3_U37 (.ZN( u0_u7_u3_n109 ) , .A( u0_u7_u3_n119 ) , .C2( u0_u7_u3_n129 ) , .B( u0_u7_u3_n138 ) , .C1( u0_u7_u3_n141 ) );
  AOI211_X1 u0_u7_u3_U38 (.B( u0_u7_u3_n119 ) , .A( u0_u7_u3_n120 ) , .C2( u0_u7_u3_n121 ) , .ZN( u0_u7_u3_n122 ) , .C1( u0_u7_u3_n179 ) );
  INV_X1 u0_u7_u3_U39 (.A( u0_u7_u3_n156 ) , .ZN( u0_u7_u3_n179 ) );
  INV_X1 u0_u7_u3_U4 (.A( u0_u7_u3_n140 ) , .ZN( u0_u7_u3_n182 ) );
  OAI22_X1 u0_u7_u3_U40 (.B1( u0_u7_u3_n118 ) , .ZN( u0_u7_u3_n120 ) , .A1( u0_u7_u3_n135 ) , .B2( u0_u7_u3_n154 ) , .A2( u0_u7_u3_n178 ) );
  AND3_X1 u0_u7_u3_U41 (.ZN( u0_u7_u3_n118 ) , .A2( u0_u7_u3_n124 ) , .A1( u0_u7_u3_n144 ) , .A3( u0_u7_u3_n152 ) );
  INV_X1 u0_u7_u3_U42 (.A( u0_u7_u3_n121 ) , .ZN( u0_u7_u3_n164 ) );
  NAND2_X1 u0_u7_u3_U43 (.ZN( u0_u7_u3_n133 ) , .A1( u0_u7_u3_n154 ) , .A2( u0_u7_u3_n164 ) );
  OAI211_X1 u0_u7_u3_U44 (.B( u0_u7_u3_n127 ) , .ZN( u0_u7_u3_n139 ) , .C1( u0_u7_u3_n150 ) , .C2( u0_u7_u3_n154 ) , .A( u0_u7_u3_n184 ) );
  INV_X1 u0_u7_u3_U45 (.A( u0_u7_u3_n125 ) , .ZN( u0_u7_u3_n184 ) );
  AOI221_X1 u0_u7_u3_U46 (.A( u0_u7_u3_n126 ) , .ZN( u0_u7_u3_n127 ) , .C2( u0_u7_u3_n132 ) , .C1( u0_u7_u3_n169 ) , .B2( u0_u7_u3_n170 ) , .B1( u0_u7_u3_n174 ) );
  OAI22_X1 u0_u7_u3_U47 (.A1( u0_u7_u3_n124 ) , .ZN( u0_u7_u3_n125 ) , .B2( u0_u7_u3_n145 ) , .A2( u0_u7_u3_n165 ) , .B1( u0_u7_u3_n167 ) );
  NOR2_X1 u0_u7_u3_U48 (.A1( u0_u7_u3_n113 ) , .ZN( u0_u7_u3_n131 ) , .A2( u0_u7_u3_n154 ) );
  NAND2_X1 u0_u7_u3_U49 (.A1( u0_u7_u3_n103 ) , .ZN( u0_u7_u3_n150 ) , .A2( u0_u7_u3_n99 ) );
  INV_X1 u0_u7_u3_U5 (.A( u0_u7_u3_n117 ) , .ZN( u0_u7_u3_n178 ) );
  NAND2_X1 u0_u7_u3_U50 (.A2( u0_u7_u3_n102 ) , .ZN( u0_u7_u3_n155 ) , .A1( u0_u7_u3_n97 ) );
  INV_X1 u0_u7_u3_U51 (.A( u0_u7_u3_n141 ) , .ZN( u0_u7_u3_n167 ) );
  AOI21_X1 u0_u7_u3_U52 (.B2( u0_u7_u3_n114 ) , .B1( u0_u7_u3_n146 ) , .A( u0_u7_u3_n154 ) , .ZN( u0_u7_u3_n94 ) );
  AOI21_X1 u0_u7_u3_U53 (.ZN( u0_u7_u3_n110 ) , .B2( u0_u7_u3_n142 ) , .B1( u0_u7_u3_n186 ) , .A( u0_u7_u3_n95 ) );
  INV_X1 u0_u7_u3_U54 (.A( u0_u7_u3_n145 ) , .ZN( u0_u7_u3_n186 ) );
  AOI21_X1 u0_u7_u3_U55 (.B1( u0_u7_u3_n124 ) , .A( u0_u7_u3_n149 ) , .B2( u0_u7_u3_n155 ) , .ZN( u0_u7_u3_n95 ) );
  INV_X1 u0_u7_u3_U56 (.A( u0_u7_u3_n149 ) , .ZN( u0_u7_u3_n169 ) );
  NAND2_X1 u0_u7_u3_U57 (.ZN( u0_u7_u3_n124 ) , .A1( u0_u7_u3_n96 ) , .A2( u0_u7_u3_n97 ) );
  NAND2_X1 u0_u7_u3_U58 (.A2( u0_u7_u3_n100 ) , .ZN( u0_u7_u3_n146 ) , .A1( u0_u7_u3_n96 ) );
  NAND2_X1 u0_u7_u3_U59 (.A1( u0_u7_u3_n101 ) , .ZN( u0_u7_u3_n145 ) , .A2( u0_u7_u3_n99 ) );
  AOI221_X1 u0_u7_u3_U6 (.A( u0_u7_u3_n131 ) , .C2( u0_u7_u3_n132 ) , .C1( u0_u7_u3_n133 ) , .ZN( u0_u7_u3_n134 ) , .B1( u0_u7_u3_n143 ) , .B2( u0_u7_u3_n177 ) );
  NAND2_X1 u0_u7_u3_U60 (.A1( u0_u7_u3_n100 ) , .ZN( u0_u7_u3_n156 ) , .A2( u0_u7_u3_n99 ) );
  NAND2_X1 u0_u7_u3_U61 (.A2( u0_u7_u3_n101 ) , .A1( u0_u7_u3_n104 ) , .ZN( u0_u7_u3_n148 ) );
  NAND2_X1 u0_u7_u3_U62 (.A1( u0_u7_u3_n100 ) , .A2( u0_u7_u3_n102 ) , .ZN( u0_u7_u3_n128 ) );
  NAND2_X1 u0_u7_u3_U63 (.A2( u0_u7_u3_n101 ) , .A1( u0_u7_u3_n102 ) , .ZN( u0_u7_u3_n152 ) );
  NAND2_X1 u0_u7_u3_U64 (.A2( u0_u7_u3_n101 ) , .ZN( u0_u7_u3_n114 ) , .A1( u0_u7_u3_n96 ) );
  NAND2_X1 u0_u7_u3_U65 (.ZN( u0_u7_u3_n107 ) , .A1( u0_u7_u3_n97 ) , .A2( u0_u7_u3_n99 ) );
  NAND2_X1 u0_u7_u3_U66 (.A2( u0_u7_u3_n100 ) , .A1( u0_u7_u3_n104 ) , .ZN( u0_u7_u3_n113 ) );
  NAND2_X1 u0_u7_u3_U67 (.A1( u0_u7_u3_n104 ) , .ZN( u0_u7_u3_n153 ) , .A2( u0_u7_u3_n97 ) );
  NAND2_X1 u0_u7_u3_U68 (.A2( u0_u7_u3_n103 ) , .A1( u0_u7_u3_n104 ) , .ZN( u0_u7_u3_n130 ) );
  NAND2_X1 u0_u7_u3_U69 (.A2( u0_u7_u3_n103 ) , .ZN( u0_u7_u3_n144 ) , .A1( u0_u7_u3_n96 ) );
  OAI22_X1 u0_u7_u3_U7 (.B2( u0_u7_u3_n147 ) , .A2( u0_u7_u3_n148 ) , .ZN( u0_u7_u3_n160 ) , .B1( u0_u7_u3_n165 ) , .A1( u0_u7_u3_n168 ) );
  NAND2_X1 u0_u7_u3_U70 (.A1( u0_u7_u3_n102 ) , .A2( u0_u7_u3_n103 ) , .ZN( u0_u7_u3_n108 ) );
  NOR2_X1 u0_u7_u3_U71 (.A2( u0_u7_X_19 ) , .A1( u0_u7_X_20 ) , .ZN( u0_u7_u3_n99 ) );
  NOR2_X1 u0_u7_u3_U72 (.A2( u0_u7_X_21 ) , .A1( u0_u7_X_24 ) , .ZN( u0_u7_u3_n103 ) );
  NOR2_X1 u0_u7_u3_U73 (.A2( u0_u7_X_24 ) , .A1( u0_u7_u3_n171 ) , .ZN( u0_u7_u3_n97 ) );
  NOR2_X1 u0_u7_u3_U74 (.A2( u0_u7_X_23 ) , .ZN( u0_u7_u3_n141 ) , .A1( u0_u7_u3_n166 ) );
  NOR2_X1 u0_u7_u3_U75 (.A2( u0_u7_X_19 ) , .A1( u0_u7_u3_n172 ) , .ZN( u0_u7_u3_n96 ) );
  NAND2_X1 u0_u7_u3_U76 (.A1( u0_u7_X_22 ) , .A2( u0_u7_X_23 ) , .ZN( u0_u7_u3_n154 ) );
  NAND2_X1 u0_u7_u3_U77 (.A1( u0_u7_X_23 ) , .ZN( u0_u7_u3_n149 ) , .A2( u0_u7_u3_n166 ) );
  NOR2_X1 u0_u7_u3_U78 (.A2( u0_u7_X_22 ) , .A1( u0_u7_X_23 ) , .ZN( u0_u7_u3_n121 ) );
  AND2_X1 u0_u7_u3_U79 (.A1( u0_u7_X_24 ) , .ZN( u0_u7_u3_n101 ) , .A2( u0_u7_u3_n171 ) );
  AND3_X1 u0_u7_u3_U8 (.A3( u0_u7_u3_n144 ) , .A2( u0_u7_u3_n145 ) , .A1( u0_u7_u3_n146 ) , .ZN( u0_u7_u3_n147 ) );
  AND2_X1 u0_u7_u3_U80 (.A1( u0_u7_X_19 ) , .ZN( u0_u7_u3_n102 ) , .A2( u0_u7_u3_n172 ) );
  AND2_X1 u0_u7_u3_U81 (.A1( u0_u7_X_21 ) , .A2( u0_u7_X_24 ) , .ZN( u0_u7_u3_n100 ) );
  AND2_X1 u0_u7_u3_U82 (.A2( u0_u7_X_19 ) , .A1( u0_u7_X_20 ) , .ZN( u0_u7_u3_n104 ) );
  INV_X1 u0_u7_u3_U83 (.A( u0_u7_X_22 ) , .ZN( u0_u7_u3_n166 ) );
  INV_X1 u0_u7_u3_U84 (.A( u0_u7_X_21 ) , .ZN( u0_u7_u3_n171 ) );
  INV_X1 u0_u7_u3_U85 (.A( u0_u7_X_20 ) , .ZN( u0_u7_u3_n172 ) );
  OR4_X1 u0_u7_u3_U86 (.ZN( u0_out7_10 ) , .A4( u0_u7_u3_n136 ) , .A3( u0_u7_u3_n137 ) , .A1( u0_u7_u3_n138 ) , .A2( u0_u7_u3_n139 ) );
  OAI222_X1 u0_u7_u3_U87 (.C1( u0_u7_u3_n128 ) , .ZN( u0_u7_u3_n137 ) , .B1( u0_u7_u3_n148 ) , .A2( u0_u7_u3_n150 ) , .B2( u0_u7_u3_n154 ) , .C2( u0_u7_u3_n164 ) , .A1( u0_u7_u3_n167 ) );
  OAI221_X1 u0_u7_u3_U88 (.A( u0_u7_u3_n134 ) , .B2( u0_u7_u3_n135 ) , .ZN( u0_u7_u3_n136 ) , .C1( u0_u7_u3_n149 ) , .B1( u0_u7_u3_n151 ) , .C2( u0_u7_u3_n183 ) );
  NAND4_X1 u0_u7_u3_U89 (.ZN( u0_out7_26 ) , .A4( u0_u7_u3_n109 ) , .A3( u0_u7_u3_n110 ) , .A2( u0_u7_u3_n111 ) , .A1( u0_u7_u3_n173 ) );
  INV_X1 u0_u7_u3_U9 (.A( u0_u7_u3_n143 ) , .ZN( u0_u7_u3_n168 ) );
  INV_X1 u0_u7_u3_U90 (.ZN( u0_u7_u3_n173 ) , .A( u0_u7_u3_n94 ) );
  OAI21_X1 u0_u7_u3_U91 (.ZN( u0_u7_u3_n111 ) , .B2( u0_u7_u3_n117 ) , .A( u0_u7_u3_n133 ) , .B1( u0_u7_u3_n176 ) );
  NAND4_X1 u0_u7_u3_U92 (.ZN( u0_out7_20 ) , .A4( u0_u7_u3_n122 ) , .A3( u0_u7_u3_n123 ) , .A1( u0_u7_u3_n175 ) , .A2( u0_u7_u3_n180 ) );
  INV_X1 u0_u7_u3_U93 (.A( u0_u7_u3_n126 ) , .ZN( u0_u7_u3_n180 ) );
  INV_X1 u0_u7_u3_U94 (.A( u0_u7_u3_n112 ) , .ZN( u0_u7_u3_n175 ) );
  NAND4_X1 u0_u7_u3_U95 (.ZN( u0_out7_1 ) , .A4( u0_u7_u3_n161 ) , .A3( u0_u7_u3_n162 ) , .A2( u0_u7_u3_n163 ) , .A1( u0_u7_u3_n185 ) );
  NAND2_X1 u0_u7_u3_U96 (.ZN( u0_u7_u3_n163 ) , .A2( u0_u7_u3_n170 ) , .A1( u0_u7_u3_n176 ) );
  AOI22_X1 u0_u7_u3_U97 (.B2( u0_u7_u3_n140 ) , .B1( u0_u7_u3_n141 ) , .A2( u0_u7_u3_n142 ) , .ZN( u0_u7_u3_n162 ) , .A1( u0_u7_u3_n177 ) );
  NAND3_X1 u0_u7_u3_U98 (.A1( u0_u7_u3_n114 ) , .ZN( u0_u7_u3_n115 ) , .A2( u0_u7_u3_n145 ) , .A3( u0_u7_u3_n153 ) );
  NAND3_X1 u0_u7_u3_U99 (.ZN( u0_u7_u3_n129 ) , .A2( u0_u7_u3_n144 ) , .A1( u0_u7_u3_n153 ) , .A3( u0_u7_u3_n182 ) );
  XOR2_X1 u0_u9_U1 (.B( u0_K10_9 ) , .A( u0_R8_6 ) , .Z( u0_u9_X_9 ) );
  XOR2_X1 u0_u9_U10 (.B( u0_K10_45 ) , .A( u0_R8_30 ) , .Z( u0_u9_X_45 ) );
  XOR2_X1 u0_u9_U11 (.B( u0_K10_44 ) , .A( u0_R8_29 ) , .Z( u0_u9_X_44 ) );
  XOR2_X1 u0_u9_U13 (.B( u0_K10_42 ) , .A( u0_R8_29 ) , .Z( u0_u9_X_42 ) );
  XOR2_X1 u0_u9_U15 (.B( u0_K10_40 ) , .A( u0_R8_27 ) , .Z( u0_u9_X_40 ) );
  XOR2_X1 u0_u9_U2 (.B( u0_K10_8 ) , .A( u0_R8_5 ) , .Z( u0_u9_X_8 ) );
  XOR2_X1 u0_u9_U23 (.B( u0_K10_33 ) , .A( u0_R8_22 ) , .Z( u0_u9_X_33 ) );
  XOR2_X1 u0_u9_U24 (.B( u0_K10_32 ) , .A( u0_R8_21 ) , .Z( u0_u9_X_32 ) );
  XOR2_X1 u0_u9_U25 (.B( u0_K10_31 ) , .A( u0_R8_20 ) , .Z( u0_u9_X_31 ) );
  XOR2_X1 u0_u9_U26 (.B( u0_K10_30 ) , .A( u0_R8_21 ) , .Z( u0_u9_X_30 ) );
  XOR2_X1 u0_u9_U27 (.B( u0_K10_2 ) , .A( u0_R8_1 ) , .Z( u0_u9_X_2 ) );
  XOR2_X1 u0_u9_U28 (.B( u0_K10_29 ) , .A( u0_R8_20 ) , .Z( u0_u9_X_29 ) );
  XOR2_X1 u0_u9_U29 (.B( u0_K10_28 ) , .A( u0_R8_19 ) , .Z( u0_u9_X_28 ) );
  XOR2_X1 u0_u9_U31 (.B( u0_K10_26 ) , .A( u0_R8_17 ) , .Z( u0_u9_X_26 ) );
  XOR2_X1 u0_u9_U33 (.B( u0_K10_24 ) , .A( u0_R8_17 ) , .Z( u0_u9_X_24 ) );
  XOR2_X1 u0_u9_U37 (.B( u0_K10_20 ) , .A( u0_R8_13 ) , .Z( u0_u9_X_20 ) );
  XOR2_X1 u0_u9_U38 (.B( u0_K10_1 ) , .A( u0_R8_32 ) , .Z( u0_u9_X_1 ) );
  XOR2_X1 u0_u9_U39 (.B( u0_K10_19 ) , .A( u0_R8_12 ) , .Z( u0_u9_X_19 ) );
  XOR2_X1 u0_u9_U4 (.B( u0_K10_6 ) , .A( u0_R8_5 ) , .Z( u0_u9_X_6 ) );
  XOR2_X1 u0_u9_U40 (.B( u0_K10_18 ) , .A( u0_R8_13 ) , .Z( u0_u9_X_18 ) );
  XOR2_X1 u0_u9_U41 (.B( u0_K10_17 ) , .A( u0_R8_12 ) , .Z( u0_u9_X_17 ) );
  XOR2_X1 u0_u9_U44 (.B( u0_K10_14 ) , .A( u0_R8_9 ) , .Z( u0_u9_X_14 ) );
  XOR2_X1 u0_u9_U46 (.B( u0_K10_12 ) , .A( u0_R8_9 ) , .Z( u0_u9_X_12 ) );
  XOR2_X1 u0_u9_U7 (.B( u0_K10_48 ) , .A( u0_R8_1 ) , .Z( u0_u9_X_48 ) );
  XOR2_X1 u0_u9_U8 (.B( u0_K10_47 ) , .A( u0_R8_32 ) , .Z( u0_u9_X_47 ) );
  AND3_X1 u0_u9_u0_U10 (.A2( u0_u9_u0_n112 ) , .ZN( u0_u9_u0_n127 ) , .A3( u0_u9_u0_n130 ) , .A1( u0_u9_u0_n148 ) );
  NAND2_X1 u0_u9_u0_U11 (.ZN( u0_u9_u0_n113 ) , .A1( u0_u9_u0_n139 ) , .A2( u0_u9_u0_n149 ) );
  AND2_X1 u0_u9_u0_U12 (.ZN( u0_u9_u0_n107 ) , .A1( u0_u9_u0_n130 ) , .A2( u0_u9_u0_n140 ) );
  AND2_X1 u0_u9_u0_U13 (.A2( u0_u9_u0_n129 ) , .A1( u0_u9_u0_n130 ) , .ZN( u0_u9_u0_n151 ) );
  AND2_X1 u0_u9_u0_U14 (.A1( u0_u9_u0_n108 ) , .A2( u0_u9_u0_n125 ) , .ZN( u0_u9_u0_n145 ) );
  INV_X1 u0_u9_u0_U15 (.A( u0_u9_u0_n143 ) , .ZN( u0_u9_u0_n173 ) );
  NOR2_X1 u0_u9_u0_U16 (.A2( u0_u9_u0_n136 ) , .ZN( u0_u9_u0_n147 ) , .A1( u0_u9_u0_n160 ) );
  AOI21_X1 u0_u9_u0_U17 (.B1( u0_u9_u0_n103 ) , .ZN( u0_u9_u0_n132 ) , .A( u0_u9_u0_n165 ) , .B2( u0_u9_u0_n93 ) );
  INV_X1 u0_u9_u0_U18 (.A( u0_u9_u0_n142 ) , .ZN( u0_u9_u0_n165 ) );
  OAI221_X1 u0_u9_u0_U19 (.C1( u0_u9_u0_n121 ) , .ZN( u0_u9_u0_n122 ) , .B2( u0_u9_u0_n127 ) , .A( u0_u9_u0_n143 ) , .B1( u0_u9_u0_n144 ) , .C2( u0_u9_u0_n147 ) );
  OAI22_X1 u0_u9_u0_U20 (.B1( u0_u9_u0_n131 ) , .A1( u0_u9_u0_n144 ) , .B2( u0_u9_u0_n147 ) , .A2( u0_u9_u0_n90 ) , .ZN( u0_u9_u0_n91 ) );
  AND3_X1 u0_u9_u0_U21 (.A3( u0_u9_u0_n121 ) , .A2( u0_u9_u0_n125 ) , .A1( u0_u9_u0_n148 ) , .ZN( u0_u9_u0_n90 ) );
  OAI22_X1 u0_u9_u0_U22 (.B1( u0_u9_u0_n125 ) , .ZN( u0_u9_u0_n126 ) , .A1( u0_u9_u0_n138 ) , .A2( u0_u9_u0_n146 ) , .B2( u0_u9_u0_n147 ) );
  NOR2_X1 u0_u9_u0_U23 (.A1( u0_u9_u0_n163 ) , .A2( u0_u9_u0_n164 ) , .ZN( u0_u9_u0_n95 ) );
  INV_X1 u0_u9_u0_U24 (.A( u0_u9_u0_n136 ) , .ZN( u0_u9_u0_n161 ) );
  NOR2_X1 u0_u9_u0_U25 (.A1( u0_u9_u0_n120 ) , .ZN( u0_u9_u0_n143 ) , .A2( u0_u9_u0_n167 ) );
  OAI221_X1 u0_u9_u0_U26 (.C1( u0_u9_u0_n112 ) , .ZN( u0_u9_u0_n120 ) , .B1( u0_u9_u0_n138 ) , .B2( u0_u9_u0_n141 ) , .C2( u0_u9_u0_n147 ) , .A( u0_u9_u0_n172 ) );
  AOI211_X1 u0_u9_u0_U27 (.B( u0_u9_u0_n115 ) , .A( u0_u9_u0_n116 ) , .C2( u0_u9_u0_n117 ) , .C1( u0_u9_u0_n118 ) , .ZN( u0_u9_u0_n119 ) );
  NAND2_X1 u0_u9_u0_U28 (.A1( u0_u9_u0_n101 ) , .A2( u0_u9_u0_n102 ) , .ZN( u0_u9_u0_n150 ) );
  AOI22_X1 u0_u9_u0_U29 (.B2( u0_u9_u0_n109 ) , .A2( u0_u9_u0_n110 ) , .ZN( u0_u9_u0_n111 ) , .B1( u0_u9_u0_n118 ) , .A1( u0_u9_u0_n160 ) );
  INV_X1 u0_u9_u0_U3 (.A( u0_u9_u0_n113 ) , .ZN( u0_u9_u0_n166 ) );
  INV_X1 u0_u9_u0_U30 (.A( u0_u9_u0_n118 ) , .ZN( u0_u9_u0_n158 ) );
  NAND2_X1 u0_u9_u0_U31 (.A2( u0_u9_u0_n100 ) , .A1( u0_u9_u0_n101 ) , .ZN( u0_u9_u0_n139 ) );
  NAND2_X1 u0_u9_u0_U32 (.A2( u0_u9_u0_n100 ) , .ZN( u0_u9_u0_n131 ) , .A1( u0_u9_u0_n92 ) );
  NAND2_X1 u0_u9_u0_U33 (.ZN( u0_u9_u0_n108 ) , .A1( u0_u9_u0_n92 ) , .A2( u0_u9_u0_n94 ) );
  AOI21_X1 u0_u9_u0_U34 (.ZN( u0_u9_u0_n104 ) , .B1( u0_u9_u0_n107 ) , .B2( u0_u9_u0_n141 ) , .A( u0_u9_u0_n144 ) );
  AOI21_X1 u0_u9_u0_U35 (.B1( u0_u9_u0_n127 ) , .B2( u0_u9_u0_n129 ) , .A( u0_u9_u0_n138 ) , .ZN( u0_u9_u0_n96 ) );
  NAND2_X1 u0_u9_u0_U36 (.A2( u0_u9_u0_n102 ) , .ZN( u0_u9_u0_n114 ) , .A1( u0_u9_u0_n92 ) );
  AOI21_X1 u0_u9_u0_U37 (.ZN( u0_u9_u0_n116 ) , .B2( u0_u9_u0_n142 ) , .A( u0_u9_u0_n144 ) , .B1( u0_u9_u0_n166 ) );
  NAND2_X1 u0_u9_u0_U38 (.A1( u0_u9_u0_n101 ) , .ZN( u0_u9_u0_n130 ) , .A2( u0_u9_u0_n94 ) );
  NAND2_X1 u0_u9_u0_U39 (.A1( u0_u9_u0_n100 ) , .A2( u0_u9_u0_n103 ) , .ZN( u0_u9_u0_n125 ) );
  AOI21_X1 u0_u9_u0_U4 (.B1( u0_u9_u0_n114 ) , .ZN( u0_u9_u0_n115 ) , .B2( u0_u9_u0_n129 ) , .A( u0_u9_u0_n161 ) );
  NAND2_X1 u0_u9_u0_U40 (.A2( u0_u9_u0_n103 ) , .ZN( u0_u9_u0_n140 ) , .A1( u0_u9_u0_n94 ) );
  INV_X1 u0_u9_u0_U41 (.A( u0_u9_u0_n138 ) , .ZN( u0_u9_u0_n160 ) );
  NAND2_X1 u0_u9_u0_U42 (.A2( u0_u9_u0_n102 ) , .A1( u0_u9_u0_n103 ) , .ZN( u0_u9_u0_n149 ) );
  NAND2_X1 u0_u9_u0_U43 (.A2( u0_u9_u0_n101 ) , .ZN( u0_u9_u0_n121 ) , .A1( u0_u9_u0_n93 ) );
  NAND2_X1 u0_u9_u0_U44 (.ZN( u0_u9_u0_n112 ) , .A2( u0_u9_u0_n92 ) , .A1( u0_u9_u0_n93 ) );
  INV_X1 u0_u9_u0_U45 (.ZN( u0_u9_u0_n172 ) , .A( u0_u9_u0_n88 ) );
  OAI222_X1 u0_u9_u0_U46 (.C1( u0_u9_u0_n108 ) , .A1( u0_u9_u0_n125 ) , .B2( u0_u9_u0_n128 ) , .B1( u0_u9_u0_n144 ) , .A2( u0_u9_u0_n158 ) , .C2( u0_u9_u0_n161 ) , .ZN( u0_u9_u0_n88 ) );
  OR3_X1 u0_u9_u0_U47 (.A3( u0_u9_u0_n152 ) , .A2( u0_u9_u0_n153 ) , .A1( u0_u9_u0_n154 ) , .ZN( u0_u9_u0_n155 ) );
  AOI21_X1 u0_u9_u0_U48 (.A( u0_u9_u0_n144 ) , .B2( u0_u9_u0_n145 ) , .B1( u0_u9_u0_n146 ) , .ZN( u0_u9_u0_n154 ) );
  AOI21_X1 u0_u9_u0_U49 (.B2( u0_u9_u0_n150 ) , .B1( u0_u9_u0_n151 ) , .ZN( u0_u9_u0_n152 ) , .A( u0_u9_u0_n158 ) );
  AOI21_X1 u0_u9_u0_U5 (.B2( u0_u9_u0_n131 ) , .ZN( u0_u9_u0_n134 ) , .B1( u0_u9_u0_n151 ) , .A( u0_u9_u0_n158 ) );
  AOI21_X1 u0_u9_u0_U50 (.A( u0_u9_u0_n147 ) , .B2( u0_u9_u0_n148 ) , .B1( u0_u9_u0_n149 ) , .ZN( u0_u9_u0_n153 ) );
  INV_X1 u0_u9_u0_U51 (.ZN( u0_u9_u0_n171 ) , .A( u0_u9_u0_n99 ) );
  OAI211_X1 u0_u9_u0_U52 (.C2( u0_u9_u0_n140 ) , .C1( u0_u9_u0_n161 ) , .A( u0_u9_u0_n169 ) , .B( u0_u9_u0_n98 ) , .ZN( u0_u9_u0_n99 ) );
  INV_X1 u0_u9_u0_U53 (.ZN( u0_u9_u0_n169 ) , .A( u0_u9_u0_n91 ) );
  AOI211_X1 u0_u9_u0_U54 (.C1( u0_u9_u0_n118 ) , .A( u0_u9_u0_n123 ) , .B( u0_u9_u0_n96 ) , .C2( u0_u9_u0_n97 ) , .ZN( u0_u9_u0_n98 ) );
  NOR2_X1 u0_u9_u0_U55 (.A2( u0_u9_X_2 ) , .ZN( u0_u9_u0_n103 ) , .A1( u0_u9_u0_n164 ) );
  NOR2_X1 u0_u9_u0_U56 (.A2( u0_u9_X_4 ) , .A1( u0_u9_X_5 ) , .ZN( u0_u9_u0_n118 ) );
  NOR2_X1 u0_u9_u0_U57 (.A2( u0_u9_X_3 ) , .A1( u0_u9_X_6 ) , .ZN( u0_u9_u0_n94 ) );
  NOR2_X1 u0_u9_u0_U58 (.A2( u0_u9_X_6 ) , .ZN( u0_u9_u0_n100 ) , .A1( u0_u9_u0_n162 ) );
  NAND2_X1 u0_u9_u0_U59 (.A2( u0_u9_X_4 ) , .A1( u0_u9_X_5 ) , .ZN( u0_u9_u0_n144 ) );
  NOR2_X1 u0_u9_u0_U6 (.A1( u0_u9_u0_n108 ) , .ZN( u0_u9_u0_n123 ) , .A2( u0_u9_u0_n158 ) );
  NOR2_X1 u0_u9_u0_U60 (.A2( u0_u9_X_5 ) , .ZN( u0_u9_u0_n136 ) , .A1( u0_u9_u0_n159 ) );
  NAND2_X1 u0_u9_u0_U61 (.A1( u0_u9_X_5 ) , .ZN( u0_u9_u0_n138 ) , .A2( u0_u9_u0_n159 ) );
  AND2_X1 u0_u9_u0_U62 (.A2( u0_u9_X_3 ) , .A1( u0_u9_X_6 ) , .ZN( u0_u9_u0_n102 ) );
  AND2_X1 u0_u9_u0_U63 (.A1( u0_u9_X_6 ) , .A2( u0_u9_u0_n162 ) , .ZN( u0_u9_u0_n93 ) );
  INV_X1 u0_u9_u0_U64 (.A( u0_u9_X_4 ) , .ZN( u0_u9_u0_n159 ) );
  INV_X1 u0_u9_u0_U65 (.A( u0_u9_X_3 ) , .ZN( u0_u9_u0_n162 ) );
  INV_X1 u0_u9_u0_U66 (.A( u0_u9_X_2 ) , .ZN( u0_u9_u0_n163 ) );
  INV_X1 u0_u9_u0_U67 (.A( u0_u9_u0_n126 ) , .ZN( u0_u9_u0_n168 ) );
  AOI211_X1 u0_u9_u0_U68 (.B( u0_u9_u0_n133 ) , .A( u0_u9_u0_n134 ) , .C2( u0_u9_u0_n135 ) , .C1( u0_u9_u0_n136 ) , .ZN( u0_u9_u0_n137 ) );
  INV_X1 u0_u9_u0_U69 (.ZN( u0_u9_u0_n174 ) , .A( u0_u9_u0_n89 ) );
  OAI21_X1 u0_u9_u0_U7 (.B1( u0_u9_u0_n150 ) , .B2( u0_u9_u0_n158 ) , .A( u0_u9_u0_n172 ) , .ZN( u0_u9_u0_n89 ) );
  AOI211_X1 u0_u9_u0_U70 (.B( u0_u9_u0_n104 ) , .A( u0_u9_u0_n105 ) , .ZN( u0_u9_u0_n106 ) , .C2( u0_u9_u0_n113 ) , .C1( u0_u9_u0_n160 ) );
  OR4_X1 u0_u9_u0_U71 (.ZN( u0_out9_17 ) , .A4( u0_u9_u0_n122 ) , .A2( u0_u9_u0_n123 ) , .A1( u0_u9_u0_n124 ) , .A3( u0_u9_u0_n170 ) );
  AOI21_X1 u0_u9_u0_U72 (.B2( u0_u9_u0_n107 ) , .ZN( u0_u9_u0_n124 ) , .B1( u0_u9_u0_n128 ) , .A( u0_u9_u0_n161 ) );
  INV_X1 u0_u9_u0_U73 (.A( u0_u9_u0_n111 ) , .ZN( u0_u9_u0_n170 ) );
  OR4_X1 u0_u9_u0_U74 (.ZN( u0_out9_31 ) , .A4( u0_u9_u0_n155 ) , .A2( u0_u9_u0_n156 ) , .A1( u0_u9_u0_n157 ) , .A3( u0_u9_u0_n173 ) );
  AOI21_X1 u0_u9_u0_U75 (.A( u0_u9_u0_n138 ) , .B2( u0_u9_u0_n139 ) , .B1( u0_u9_u0_n140 ) , .ZN( u0_u9_u0_n157 ) );
  AOI21_X1 u0_u9_u0_U76 (.B2( u0_u9_u0_n141 ) , .B1( u0_u9_u0_n142 ) , .ZN( u0_u9_u0_n156 ) , .A( u0_u9_u0_n161 ) );
  AOI21_X1 u0_u9_u0_U77 (.B1( u0_u9_u0_n132 ) , .ZN( u0_u9_u0_n133 ) , .A( u0_u9_u0_n144 ) , .B2( u0_u9_u0_n166 ) );
  OAI22_X1 u0_u9_u0_U78 (.ZN( u0_u9_u0_n105 ) , .A2( u0_u9_u0_n132 ) , .B1( u0_u9_u0_n146 ) , .A1( u0_u9_u0_n147 ) , .B2( u0_u9_u0_n161 ) );
  NAND2_X1 u0_u9_u0_U79 (.ZN( u0_u9_u0_n110 ) , .A2( u0_u9_u0_n132 ) , .A1( u0_u9_u0_n145 ) );
  AND2_X1 u0_u9_u0_U8 (.A1( u0_u9_u0_n114 ) , .A2( u0_u9_u0_n121 ) , .ZN( u0_u9_u0_n146 ) );
  INV_X1 u0_u9_u0_U80 (.A( u0_u9_u0_n119 ) , .ZN( u0_u9_u0_n167 ) );
  NAND2_X1 u0_u9_u0_U81 (.ZN( u0_u9_u0_n148 ) , .A1( u0_u9_u0_n93 ) , .A2( u0_u9_u0_n95 ) );
  NAND2_X1 u0_u9_u0_U82 (.A1( u0_u9_u0_n100 ) , .ZN( u0_u9_u0_n129 ) , .A2( u0_u9_u0_n95 ) );
  NAND2_X1 u0_u9_u0_U83 (.A1( u0_u9_u0_n102 ) , .ZN( u0_u9_u0_n128 ) , .A2( u0_u9_u0_n95 ) );
  NOR2_X1 u0_u9_u0_U84 (.A2( u0_u9_X_1 ) , .A1( u0_u9_X_2 ) , .ZN( u0_u9_u0_n92 ) );
  NAND2_X1 u0_u9_u0_U85 (.ZN( u0_u9_u0_n142 ) , .A1( u0_u9_u0_n94 ) , .A2( u0_u9_u0_n95 ) );
  NOR2_X1 u0_u9_u0_U86 (.A2( u0_u9_X_1 ) , .ZN( u0_u9_u0_n101 ) , .A1( u0_u9_u0_n163 ) );
  INV_X1 u0_u9_u0_U87 (.A( u0_u9_X_1 ) , .ZN( u0_u9_u0_n164 ) );
  NAND3_X1 u0_u9_u0_U88 (.ZN( u0_out9_23 ) , .A3( u0_u9_u0_n137 ) , .A1( u0_u9_u0_n168 ) , .A2( u0_u9_u0_n171 ) );
  NAND3_X1 u0_u9_u0_U89 (.A3( u0_u9_u0_n127 ) , .A2( u0_u9_u0_n128 ) , .ZN( u0_u9_u0_n135 ) , .A1( u0_u9_u0_n150 ) );
  AND2_X1 u0_u9_u0_U9 (.A1( u0_u9_u0_n131 ) , .ZN( u0_u9_u0_n141 ) , .A2( u0_u9_u0_n150 ) );
  NAND3_X1 u0_u9_u0_U90 (.ZN( u0_u9_u0_n117 ) , .A3( u0_u9_u0_n132 ) , .A2( u0_u9_u0_n139 ) , .A1( u0_u9_u0_n148 ) );
  NAND3_X1 u0_u9_u0_U91 (.ZN( u0_u9_u0_n109 ) , .A2( u0_u9_u0_n114 ) , .A3( u0_u9_u0_n140 ) , .A1( u0_u9_u0_n149 ) );
  NAND3_X1 u0_u9_u0_U92 (.ZN( u0_out9_9 ) , .A3( u0_u9_u0_n106 ) , .A2( u0_u9_u0_n171 ) , .A1( u0_u9_u0_n174 ) );
  NAND3_X1 u0_u9_u0_U93 (.A2( u0_u9_u0_n128 ) , .A1( u0_u9_u0_n132 ) , .A3( u0_u9_u0_n146 ) , .ZN( u0_u9_u0_n97 ) );
  NOR2_X1 u0_u9_u1_U10 (.A1( u0_u9_u1_n112 ) , .A2( u0_u9_u1_n116 ) , .ZN( u0_u9_u1_n118 ) );
  NAND3_X1 u0_u9_u1_U100 (.ZN( u0_u9_u1_n113 ) , .A1( u0_u9_u1_n120 ) , .A3( u0_u9_u1_n133 ) , .A2( u0_u9_u1_n155 ) );
  OAI21_X1 u0_u9_u1_U11 (.ZN( u0_u9_u1_n101 ) , .B1( u0_u9_u1_n141 ) , .A( u0_u9_u1_n146 ) , .B2( u0_u9_u1_n183 ) );
  AOI21_X1 u0_u9_u1_U12 (.B2( u0_u9_u1_n155 ) , .B1( u0_u9_u1_n156 ) , .ZN( u0_u9_u1_n157 ) , .A( u0_u9_u1_n174 ) );
  NAND2_X1 u0_u9_u1_U13 (.ZN( u0_u9_u1_n140 ) , .A2( u0_u9_u1_n150 ) , .A1( u0_u9_u1_n155 ) );
  NAND2_X1 u0_u9_u1_U14 (.A1( u0_u9_u1_n131 ) , .ZN( u0_u9_u1_n147 ) , .A2( u0_u9_u1_n153 ) );
  INV_X1 u0_u9_u1_U15 (.A( u0_u9_u1_n139 ) , .ZN( u0_u9_u1_n174 ) );
  OR4_X1 u0_u9_u1_U16 (.A4( u0_u9_u1_n106 ) , .A3( u0_u9_u1_n107 ) , .ZN( u0_u9_u1_n108 ) , .A1( u0_u9_u1_n117 ) , .A2( u0_u9_u1_n184 ) );
  AOI21_X1 u0_u9_u1_U17 (.ZN( u0_u9_u1_n106 ) , .A( u0_u9_u1_n112 ) , .B1( u0_u9_u1_n154 ) , .B2( u0_u9_u1_n156 ) );
  AOI21_X1 u0_u9_u1_U18 (.ZN( u0_u9_u1_n107 ) , .B1( u0_u9_u1_n134 ) , .B2( u0_u9_u1_n149 ) , .A( u0_u9_u1_n174 ) );
  INV_X1 u0_u9_u1_U19 (.A( u0_u9_u1_n101 ) , .ZN( u0_u9_u1_n184 ) );
  INV_X1 u0_u9_u1_U20 (.A( u0_u9_u1_n112 ) , .ZN( u0_u9_u1_n171 ) );
  NAND2_X1 u0_u9_u1_U21 (.ZN( u0_u9_u1_n141 ) , .A1( u0_u9_u1_n153 ) , .A2( u0_u9_u1_n156 ) );
  AND2_X1 u0_u9_u1_U22 (.A1( u0_u9_u1_n123 ) , .ZN( u0_u9_u1_n134 ) , .A2( u0_u9_u1_n161 ) );
  NAND2_X1 u0_u9_u1_U23 (.A2( u0_u9_u1_n115 ) , .A1( u0_u9_u1_n116 ) , .ZN( u0_u9_u1_n148 ) );
  NAND2_X1 u0_u9_u1_U24 (.A2( u0_u9_u1_n133 ) , .A1( u0_u9_u1_n135 ) , .ZN( u0_u9_u1_n159 ) );
  NAND2_X1 u0_u9_u1_U25 (.A2( u0_u9_u1_n115 ) , .A1( u0_u9_u1_n120 ) , .ZN( u0_u9_u1_n132 ) );
  INV_X1 u0_u9_u1_U26 (.A( u0_u9_u1_n154 ) , .ZN( u0_u9_u1_n178 ) );
  INV_X1 u0_u9_u1_U27 (.A( u0_u9_u1_n151 ) , .ZN( u0_u9_u1_n183 ) );
  AND2_X1 u0_u9_u1_U28 (.A1( u0_u9_u1_n129 ) , .A2( u0_u9_u1_n133 ) , .ZN( u0_u9_u1_n149 ) );
  INV_X1 u0_u9_u1_U29 (.A( u0_u9_u1_n131 ) , .ZN( u0_u9_u1_n180 ) );
  INV_X1 u0_u9_u1_U3 (.A( u0_u9_u1_n159 ) , .ZN( u0_u9_u1_n182 ) );
  OAI221_X1 u0_u9_u1_U30 (.A( u0_u9_u1_n119 ) , .C2( u0_u9_u1_n129 ) , .ZN( u0_u9_u1_n138 ) , .B2( u0_u9_u1_n152 ) , .C1( u0_u9_u1_n174 ) , .B1( u0_u9_u1_n187 ) );
  INV_X1 u0_u9_u1_U31 (.A( u0_u9_u1_n148 ) , .ZN( u0_u9_u1_n187 ) );
  AOI211_X1 u0_u9_u1_U32 (.B( u0_u9_u1_n117 ) , .A( u0_u9_u1_n118 ) , .ZN( u0_u9_u1_n119 ) , .C2( u0_u9_u1_n146 ) , .C1( u0_u9_u1_n159 ) );
  NOR2_X1 u0_u9_u1_U33 (.A1( u0_u9_u1_n168 ) , .A2( u0_u9_u1_n176 ) , .ZN( u0_u9_u1_n98 ) );
  AOI211_X1 u0_u9_u1_U34 (.B( u0_u9_u1_n162 ) , .A( u0_u9_u1_n163 ) , .C2( u0_u9_u1_n164 ) , .ZN( u0_u9_u1_n165 ) , .C1( u0_u9_u1_n171 ) );
  AOI21_X1 u0_u9_u1_U35 (.A( u0_u9_u1_n160 ) , .B2( u0_u9_u1_n161 ) , .ZN( u0_u9_u1_n162 ) , .B1( u0_u9_u1_n182 ) );
  OR2_X1 u0_u9_u1_U36 (.A2( u0_u9_u1_n157 ) , .A1( u0_u9_u1_n158 ) , .ZN( u0_u9_u1_n163 ) );
  NAND2_X1 u0_u9_u1_U37 (.A1( u0_u9_u1_n128 ) , .ZN( u0_u9_u1_n146 ) , .A2( u0_u9_u1_n160 ) );
  NAND2_X1 u0_u9_u1_U38 (.A2( u0_u9_u1_n112 ) , .ZN( u0_u9_u1_n139 ) , .A1( u0_u9_u1_n152 ) );
  NAND2_X1 u0_u9_u1_U39 (.A1( u0_u9_u1_n105 ) , .ZN( u0_u9_u1_n156 ) , .A2( u0_u9_u1_n99 ) );
  AOI221_X1 u0_u9_u1_U4 (.A( u0_u9_u1_n138 ) , .C2( u0_u9_u1_n139 ) , .C1( u0_u9_u1_n140 ) , .B2( u0_u9_u1_n141 ) , .ZN( u0_u9_u1_n142 ) , .B1( u0_u9_u1_n175 ) );
  AOI221_X1 u0_u9_u1_U40 (.B1( u0_u9_u1_n140 ) , .ZN( u0_u9_u1_n167 ) , .B2( u0_u9_u1_n172 ) , .C2( u0_u9_u1_n175 ) , .C1( u0_u9_u1_n178 ) , .A( u0_u9_u1_n188 ) );
  INV_X1 u0_u9_u1_U41 (.ZN( u0_u9_u1_n188 ) , .A( u0_u9_u1_n97 ) );
  AOI211_X1 u0_u9_u1_U42 (.A( u0_u9_u1_n118 ) , .C1( u0_u9_u1_n132 ) , .C2( u0_u9_u1_n139 ) , .B( u0_u9_u1_n96 ) , .ZN( u0_u9_u1_n97 ) );
  AOI21_X1 u0_u9_u1_U43 (.B2( u0_u9_u1_n121 ) , .B1( u0_u9_u1_n135 ) , .A( u0_u9_u1_n152 ) , .ZN( u0_u9_u1_n96 ) );
  NOR2_X1 u0_u9_u1_U44 (.ZN( u0_u9_u1_n117 ) , .A1( u0_u9_u1_n121 ) , .A2( u0_u9_u1_n160 ) );
  OAI21_X1 u0_u9_u1_U45 (.B2( u0_u9_u1_n123 ) , .ZN( u0_u9_u1_n145 ) , .B1( u0_u9_u1_n160 ) , .A( u0_u9_u1_n185 ) );
  INV_X1 u0_u9_u1_U46 (.A( u0_u9_u1_n122 ) , .ZN( u0_u9_u1_n185 ) );
  AOI21_X1 u0_u9_u1_U47 (.B2( u0_u9_u1_n120 ) , .B1( u0_u9_u1_n121 ) , .ZN( u0_u9_u1_n122 ) , .A( u0_u9_u1_n128 ) );
  AOI21_X1 u0_u9_u1_U48 (.A( u0_u9_u1_n128 ) , .B2( u0_u9_u1_n129 ) , .ZN( u0_u9_u1_n130 ) , .B1( u0_u9_u1_n150 ) );
  NAND2_X1 u0_u9_u1_U49 (.ZN( u0_u9_u1_n112 ) , .A1( u0_u9_u1_n169 ) , .A2( u0_u9_u1_n170 ) );
  AOI211_X1 u0_u9_u1_U5 (.ZN( u0_u9_u1_n124 ) , .A( u0_u9_u1_n138 ) , .C2( u0_u9_u1_n139 ) , .B( u0_u9_u1_n145 ) , .C1( u0_u9_u1_n147 ) );
  NAND2_X1 u0_u9_u1_U50 (.ZN( u0_u9_u1_n129 ) , .A2( u0_u9_u1_n95 ) , .A1( u0_u9_u1_n98 ) );
  NAND2_X1 u0_u9_u1_U51 (.A1( u0_u9_u1_n102 ) , .ZN( u0_u9_u1_n154 ) , .A2( u0_u9_u1_n99 ) );
  NAND2_X1 u0_u9_u1_U52 (.A2( u0_u9_u1_n100 ) , .ZN( u0_u9_u1_n135 ) , .A1( u0_u9_u1_n99 ) );
  AOI21_X1 u0_u9_u1_U53 (.A( u0_u9_u1_n152 ) , .B2( u0_u9_u1_n153 ) , .B1( u0_u9_u1_n154 ) , .ZN( u0_u9_u1_n158 ) );
  INV_X1 u0_u9_u1_U54 (.A( u0_u9_u1_n160 ) , .ZN( u0_u9_u1_n175 ) );
  NAND2_X1 u0_u9_u1_U55 (.A1( u0_u9_u1_n100 ) , .ZN( u0_u9_u1_n116 ) , .A2( u0_u9_u1_n95 ) );
  NAND2_X1 u0_u9_u1_U56 (.A1( u0_u9_u1_n102 ) , .ZN( u0_u9_u1_n131 ) , .A2( u0_u9_u1_n95 ) );
  NAND2_X1 u0_u9_u1_U57 (.A2( u0_u9_u1_n104 ) , .ZN( u0_u9_u1_n121 ) , .A1( u0_u9_u1_n98 ) );
  NAND2_X1 u0_u9_u1_U58 (.A1( u0_u9_u1_n103 ) , .ZN( u0_u9_u1_n153 ) , .A2( u0_u9_u1_n98 ) );
  NAND2_X1 u0_u9_u1_U59 (.A2( u0_u9_u1_n104 ) , .A1( u0_u9_u1_n105 ) , .ZN( u0_u9_u1_n133 ) );
  AOI22_X1 u0_u9_u1_U6 (.B2( u0_u9_u1_n136 ) , .A2( u0_u9_u1_n137 ) , .ZN( u0_u9_u1_n143 ) , .A1( u0_u9_u1_n171 ) , .B1( u0_u9_u1_n173 ) );
  NAND2_X1 u0_u9_u1_U60 (.ZN( u0_u9_u1_n150 ) , .A2( u0_u9_u1_n98 ) , .A1( u0_u9_u1_n99 ) );
  NAND2_X1 u0_u9_u1_U61 (.A1( u0_u9_u1_n105 ) , .ZN( u0_u9_u1_n155 ) , .A2( u0_u9_u1_n95 ) );
  OAI21_X1 u0_u9_u1_U62 (.ZN( u0_u9_u1_n109 ) , .B1( u0_u9_u1_n129 ) , .B2( u0_u9_u1_n160 ) , .A( u0_u9_u1_n167 ) );
  NAND2_X1 u0_u9_u1_U63 (.A2( u0_u9_u1_n100 ) , .A1( u0_u9_u1_n103 ) , .ZN( u0_u9_u1_n120 ) );
  NAND2_X1 u0_u9_u1_U64 (.A1( u0_u9_u1_n102 ) , .A2( u0_u9_u1_n104 ) , .ZN( u0_u9_u1_n115 ) );
  NAND2_X1 u0_u9_u1_U65 (.A2( u0_u9_u1_n100 ) , .A1( u0_u9_u1_n104 ) , .ZN( u0_u9_u1_n151 ) );
  NAND2_X1 u0_u9_u1_U66 (.A2( u0_u9_u1_n103 ) , .A1( u0_u9_u1_n105 ) , .ZN( u0_u9_u1_n161 ) );
  INV_X1 u0_u9_u1_U67 (.A( u0_u9_u1_n152 ) , .ZN( u0_u9_u1_n173 ) );
  INV_X1 u0_u9_u1_U68 (.A( u0_u9_u1_n128 ) , .ZN( u0_u9_u1_n172 ) );
  NAND2_X1 u0_u9_u1_U69 (.A2( u0_u9_u1_n102 ) , .A1( u0_u9_u1_n103 ) , .ZN( u0_u9_u1_n123 ) );
  INV_X1 u0_u9_u1_U7 (.A( u0_u9_u1_n147 ) , .ZN( u0_u9_u1_n181 ) );
  NOR2_X1 u0_u9_u1_U70 (.A2( u0_u9_X_7 ) , .A1( u0_u9_X_8 ) , .ZN( u0_u9_u1_n95 ) );
  NOR2_X1 u0_u9_u1_U71 (.A1( u0_u9_X_12 ) , .A2( u0_u9_X_9 ) , .ZN( u0_u9_u1_n100 ) );
  NOR2_X1 u0_u9_u1_U72 (.A2( u0_u9_X_8 ) , .A1( u0_u9_u1_n177 ) , .ZN( u0_u9_u1_n99 ) );
  NOR2_X1 u0_u9_u1_U73 (.A2( u0_u9_X_12 ) , .ZN( u0_u9_u1_n102 ) , .A1( u0_u9_u1_n176 ) );
  NOR2_X1 u0_u9_u1_U74 (.A2( u0_u9_X_9 ) , .ZN( u0_u9_u1_n105 ) , .A1( u0_u9_u1_n168 ) );
  NAND2_X1 u0_u9_u1_U75 (.A1( u0_u9_X_10 ) , .ZN( u0_u9_u1_n160 ) , .A2( u0_u9_u1_n169 ) );
  NAND2_X1 u0_u9_u1_U76 (.A2( u0_u9_X_10 ) , .A1( u0_u9_X_11 ) , .ZN( u0_u9_u1_n152 ) );
  NAND2_X1 u0_u9_u1_U77 (.A1( u0_u9_X_11 ) , .ZN( u0_u9_u1_n128 ) , .A2( u0_u9_u1_n170 ) );
  AND2_X1 u0_u9_u1_U78 (.A2( u0_u9_X_7 ) , .A1( u0_u9_X_8 ) , .ZN( u0_u9_u1_n104 ) );
  AND2_X1 u0_u9_u1_U79 (.A1( u0_u9_X_8 ) , .ZN( u0_u9_u1_n103 ) , .A2( u0_u9_u1_n177 ) );
  AOI22_X1 u0_u9_u1_U8 (.B2( u0_u9_u1_n113 ) , .A2( u0_u9_u1_n114 ) , .ZN( u0_u9_u1_n125 ) , .A1( u0_u9_u1_n171 ) , .B1( u0_u9_u1_n173 ) );
  INV_X1 u0_u9_u1_U80 (.A( u0_u9_X_10 ) , .ZN( u0_u9_u1_n170 ) );
  INV_X1 u0_u9_u1_U81 (.A( u0_u9_X_9 ) , .ZN( u0_u9_u1_n176 ) );
  INV_X1 u0_u9_u1_U82 (.A( u0_u9_X_11 ) , .ZN( u0_u9_u1_n169 ) );
  INV_X1 u0_u9_u1_U83 (.A( u0_u9_X_12 ) , .ZN( u0_u9_u1_n168 ) );
  INV_X1 u0_u9_u1_U84 (.A( u0_u9_X_7 ) , .ZN( u0_u9_u1_n177 ) );
  NAND4_X1 u0_u9_u1_U85 (.ZN( u0_out9_28 ) , .A4( u0_u9_u1_n124 ) , .A3( u0_u9_u1_n125 ) , .A2( u0_u9_u1_n126 ) , .A1( u0_u9_u1_n127 ) );
  OAI21_X1 u0_u9_u1_U86 (.ZN( u0_u9_u1_n127 ) , .B2( u0_u9_u1_n139 ) , .B1( u0_u9_u1_n175 ) , .A( u0_u9_u1_n183 ) );
  OAI21_X1 u0_u9_u1_U87 (.ZN( u0_u9_u1_n126 ) , .B2( u0_u9_u1_n140 ) , .A( u0_u9_u1_n146 ) , .B1( u0_u9_u1_n178 ) );
  NAND4_X1 u0_u9_u1_U88 (.ZN( u0_out9_18 ) , .A4( u0_u9_u1_n165 ) , .A3( u0_u9_u1_n166 ) , .A1( u0_u9_u1_n167 ) , .A2( u0_u9_u1_n186 ) );
  AOI22_X1 u0_u9_u1_U89 (.B2( u0_u9_u1_n146 ) , .B1( u0_u9_u1_n147 ) , .A2( u0_u9_u1_n148 ) , .ZN( u0_u9_u1_n166 ) , .A1( u0_u9_u1_n172 ) );
  NAND2_X1 u0_u9_u1_U9 (.ZN( u0_u9_u1_n114 ) , .A1( u0_u9_u1_n134 ) , .A2( u0_u9_u1_n156 ) );
  INV_X1 u0_u9_u1_U90 (.A( u0_u9_u1_n145 ) , .ZN( u0_u9_u1_n186 ) );
  NAND4_X1 u0_u9_u1_U91 (.ZN( u0_out9_2 ) , .A4( u0_u9_u1_n142 ) , .A3( u0_u9_u1_n143 ) , .A2( u0_u9_u1_n144 ) , .A1( u0_u9_u1_n179 ) );
  OAI21_X1 u0_u9_u1_U92 (.B2( u0_u9_u1_n132 ) , .ZN( u0_u9_u1_n144 ) , .A( u0_u9_u1_n146 ) , .B1( u0_u9_u1_n180 ) );
  INV_X1 u0_u9_u1_U93 (.A( u0_u9_u1_n130 ) , .ZN( u0_u9_u1_n179 ) );
  OR4_X1 u0_u9_u1_U94 (.ZN( u0_out9_13 ) , .A4( u0_u9_u1_n108 ) , .A3( u0_u9_u1_n109 ) , .A2( u0_u9_u1_n110 ) , .A1( u0_u9_u1_n111 ) );
  AOI21_X1 u0_u9_u1_U95 (.ZN( u0_u9_u1_n110 ) , .A( u0_u9_u1_n116 ) , .B1( u0_u9_u1_n152 ) , .B2( u0_u9_u1_n160 ) );
  AOI21_X1 u0_u9_u1_U96 (.ZN( u0_u9_u1_n111 ) , .A( u0_u9_u1_n128 ) , .B2( u0_u9_u1_n131 ) , .B1( u0_u9_u1_n135 ) );
  NAND3_X1 u0_u9_u1_U97 (.A3( u0_u9_u1_n149 ) , .A2( u0_u9_u1_n150 ) , .A1( u0_u9_u1_n151 ) , .ZN( u0_u9_u1_n164 ) );
  NAND3_X1 u0_u9_u1_U98 (.A3( u0_u9_u1_n134 ) , .A2( u0_u9_u1_n135 ) , .ZN( u0_u9_u1_n136 ) , .A1( u0_u9_u1_n151 ) );
  NAND3_X1 u0_u9_u1_U99 (.A1( u0_u9_u1_n133 ) , .ZN( u0_u9_u1_n137 ) , .A2( u0_u9_u1_n154 ) , .A3( u0_u9_u1_n181 ) );
  OAI22_X1 u0_u9_u2_U10 (.B1( u0_u9_u2_n151 ) , .A2( u0_u9_u2_n152 ) , .A1( u0_u9_u2_n153 ) , .ZN( u0_u9_u2_n160 ) , .B2( u0_u9_u2_n168 ) );
  NAND3_X1 u0_u9_u2_U100 (.A2( u0_u9_u2_n100 ) , .A1( u0_u9_u2_n104 ) , .A3( u0_u9_u2_n138 ) , .ZN( u0_u9_u2_n98 ) );
  NOR3_X1 u0_u9_u2_U11 (.A1( u0_u9_u2_n150 ) , .ZN( u0_u9_u2_n151 ) , .A3( u0_u9_u2_n175 ) , .A2( u0_u9_u2_n188 ) );
  AOI21_X1 u0_u9_u2_U12 (.B2( u0_u9_u2_n123 ) , .ZN( u0_u9_u2_n125 ) , .A( u0_u9_u2_n171 ) , .B1( u0_u9_u2_n184 ) );
  INV_X1 u0_u9_u2_U13 (.A( u0_u9_u2_n150 ) , .ZN( u0_u9_u2_n184 ) );
  AOI21_X1 u0_u9_u2_U14 (.ZN( u0_u9_u2_n144 ) , .B2( u0_u9_u2_n155 ) , .A( u0_u9_u2_n172 ) , .B1( u0_u9_u2_n185 ) );
  AOI21_X1 u0_u9_u2_U15 (.B2( u0_u9_u2_n143 ) , .ZN( u0_u9_u2_n145 ) , .B1( u0_u9_u2_n152 ) , .A( u0_u9_u2_n171 ) );
  INV_X1 u0_u9_u2_U16 (.A( u0_u9_u2_n156 ) , .ZN( u0_u9_u2_n171 ) );
  INV_X1 u0_u9_u2_U17 (.A( u0_u9_u2_n120 ) , .ZN( u0_u9_u2_n188 ) );
  NAND2_X1 u0_u9_u2_U18 (.A2( u0_u9_u2_n122 ) , .ZN( u0_u9_u2_n150 ) , .A1( u0_u9_u2_n152 ) );
  INV_X1 u0_u9_u2_U19 (.A( u0_u9_u2_n153 ) , .ZN( u0_u9_u2_n170 ) );
  INV_X1 u0_u9_u2_U20 (.A( u0_u9_u2_n137 ) , .ZN( u0_u9_u2_n173 ) );
  NAND2_X1 u0_u9_u2_U21 (.A1( u0_u9_u2_n132 ) , .A2( u0_u9_u2_n139 ) , .ZN( u0_u9_u2_n157 ) );
  INV_X1 u0_u9_u2_U22 (.A( u0_u9_u2_n113 ) , .ZN( u0_u9_u2_n178 ) );
  INV_X1 u0_u9_u2_U23 (.A( u0_u9_u2_n139 ) , .ZN( u0_u9_u2_n175 ) );
  INV_X1 u0_u9_u2_U24 (.A( u0_u9_u2_n155 ) , .ZN( u0_u9_u2_n181 ) );
  INV_X1 u0_u9_u2_U25 (.A( u0_u9_u2_n119 ) , .ZN( u0_u9_u2_n177 ) );
  INV_X1 u0_u9_u2_U26 (.A( u0_u9_u2_n116 ) , .ZN( u0_u9_u2_n180 ) );
  INV_X1 u0_u9_u2_U27 (.A( u0_u9_u2_n131 ) , .ZN( u0_u9_u2_n179 ) );
  INV_X1 u0_u9_u2_U28 (.A( u0_u9_u2_n154 ) , .ZN( u0_u9_u2_n176 ) );
  NAND2_X1 u0_u9_u2_U29 (.A2( u0_u9_u2_n116 ) , .A1( u0_u9_u2_n117 ) , .ZN( u0_u9_u2_n118 ) );
  NOR2_X1 u0_u9_u2_U3 (.ZN( u0_u9_u2_n121 ) , .A2( u0_u9_u2_n177 ) , .A1( u0_u9_u2_n180 ) );
  INV_X1 u0_u9_u2_U30 (.A( u0_u9_u2_n132 ) , .ZN( u0_u9_u2_n182 ) );
  INV_X1 u0_u9_u2_U31 (.A( u0_u9_u2_n158 ) , .ZN( u0_u9_u2_n183 ) );
  OAI21_X1 u0_u9_u2_U32 (.A( u0_u9_u2_n156 ) , .B1( u0_u9_u2_n157 ) , .ZN( u0_u9_u2_n158 ) , .B2( u0_u9_u2_n179 ) );
  NOR2_X1 u0_u9_u2_U33 (.ZN( u0_u9_u2_n156 ) , .A1( u0_u9_u2_n166 ) , .A2( u0_u9_u2_n169 ) );
  NOR2_X1 u0_u9_u2_U34 (.A2( u0_u9_u2_n114 ) , .ZN( u0_u9_u2_n137 ) , .A1( u0_u9_u2_n140 ) );
  NOR2_X1 u0_u9_u2_U35 (.A2( u0_u9_u2_n138 ) , .ZN( u0_u9_u2_n153 ) , .A1( u0_u9_u2_n156 ) );
  AOI211_X1 u0_u9_u2_U36 (.ZN( u0_u9_u2_n130 ) , .C1( u0_u9_u2_n138 ) , .C2( u0_u9_u2_n179 ) , .B( u0_u9_u2_n96 ) , .A( u0_u9_u2_n97 ) );
  OAI22_X1 u0_u9_u2_U37 (.B1( u0_u9_u2_n133 ) , .A2( u0_u9_u2_n137 ) , .A1( u0_u9_u2_n152 ) , .B2( u0_u9_u2_n168 ) , .ZN( u0_u9_u2_n97 ) );
  OAI221_X1 u0_u9_u2_U38 (.B1( u0_u9_u2_n113 ) , .C1( u0_u9_u2_n132 ) , .A( u0_u9_u2_n149 ) , .B2( u0_u9_u2_n171 ) , .C2( u0_u9_u2_n172 ) , .ZN( u0_u9_u2_n96 ) );
  OAI221_X1 u0_u9_u2_U39 (.A( u0_u9_u2_n115 ) , .C2( u0_u9_u2_n123 ) , .B2( u0_u9_u2_n143 ) , .B1( u0_u9_u2_n153 ) , .ZN( u0_u9_u2_n163 ) , .C1( u0_u9_u2_n168 ) );
  INV_X1 u0_u9_u2_U4 (.A( u0_u9_u2_n134 ) , .ZN( u0_u9_u2_n185 ) );
  OAI21_X1 u0_u9_u2_U40 (.A( u0_u9_u2_n114 ) , .ZN( u0_u9_u2_n115 ) , .B1( u0_u9_u2_n176 ) , .B2( u0_u9_u2_n178 ) );
  OAI221_X1 u0_u9_u2_U41 (.A( u0_u9_u2_n135 ) , .B2( u0_u9_u2_n136 ) , .B1( u0_u9_u2_n137 ) , .ZN( u0_u9_u2_n162 ) , .C2( u0_u9_u2_n167 ) , .C1( u0_u9_u2_n185 ) );
  AND3_X1 u0_u9_u2_U42 (.A3( u0_u9_u2_n131 ) , .A2( u0_u9_u2_n132 ) , .A1( u0_u9_u2_n133 ) , .ZN( u0_u9_u2_n136 ) );
  AOI22_X1 u0_u9_u2_U43 (.ZN( u0_u9_u2_n135 ) , .B1( u0_u9_u2_n140 ) , .A1( u0_u9_u2_n156 ) , .B2( u0_u9_u2_n180 ) , .A2( u0_u9_u2_n188 ) );
  AOI21_X1 u0_u9_u2_U44 (.ZN( u0_u9_u2_n149 ) , .B1( u0_u9_u2_n173 ) , .B2( u0_u9_u2_n188 ) , .A( u0_u9_u2_n95 ) );
  AND3_X1 u0_u9_u2_U45 (.A2( u0_u9_u2_n100 ) , .A1( u0_u9_u2_n104 ) , .A3( u0_u9_u2_n156 ) , .ZN( u0_u9_u2_n95 ) );
  OAI21_X1 u0_u9_u2_U46 (.A( u0_u9_u2_n141 ) , .B2( u0_u9_u2_n142 ) , .ZN( u0_u9_u2_n146 ) , .B1( u0_u9_u2_n153 ) );
  OAI21_X1 u0_u9_u2_U47 (.A( u0_u9_u2_n140 ) , .ZN( u0_u9_u2_n141 ) , .B1( u0_u9_u2_n176 ) , .B2( u0_u9_u2_n177 ) );
  NOR3_X1 u0_u9_u2_U48 (.ZN( u0_u9_u2_n142 ) , .A3( u0_u9_u2_n175 ) , .A2( u0_u9_u2_n178 ) , .A1( u0_u9_u2_n181 ) );
  OAI21_X1 u0_u9_u2_U49 (.A( u0_u9_u2_n101 ) , .B2( u0_u9_u2_n121 ) , .B1( u0_u9_u2_n153 ) , .ZN( u0_u9_u2_n164 ) );
  NOR4_X1 u0_u9_u2_U5 (.A4( u0_u9_u2_n124 ) , .A3( u0_u9_u2_n125 ) , .A2( u0_u9_u2_n126 ) , .A1( u0_u9_u2_n127 ) , .ZN( u0_u9_u2_n128 ) );
  NAND2_X1 u0_u9_u2_U50 (.A2( u0_u9_u2_n100 ) , .A1( u0_u9_u2_n107 ) , .ZN( u0_u9_u2_n155 ) );
  NAND2_X1 u0_u9_u2_U51 (.A2( u0_u9_u2_n105 ) , .A1( u0_u9_u2_n108 ) , .ZN( u0_u9_u2_n143 ) );
  NAND2_X1 u0_u9_u2_U52 (.A1( u0_u9_u2_n104 ) , .A2( u0_u9_u2_n106 ) , .ZN( u0_u9_u2_n152 ) );
  NAND2_X1 u0_u9_u2_U53 (.A1( u0_u9_u2_n100 ) , .A2( u0_u9_u2_n105 ) , .ZN( u0_u9_u2_n132 ) );
  INV_X1 u0_u9_u2_U54 (.A( u0_u9_u2_n140 ) , .ZN( u0_u9_u2_n168 ) );
  INV_X1 u0_u9_u2_U55 (.A( u0_u9_u2_n138 ) , .ZN( u0_u9_u2_n167 ) );
  NAND2_X1 u0_u9_u2_U56 (.A1( u0_u9_u2_n102 ) , .A2( u0_u9_u2_n106 ) , .ZN( u0_u9_u2_n113 ) );
  NAND2_X1 u0_u9_u2_U57 (.A1( u0_u9_u2_n106 ) , .A2( u0_u9_u2_n107 ) , .ZN( u0_u9_u2_n131 ) );
  NAND2_X1 u0_u9_u2_U58 (.A1( u0_u9_u2_n103 ) , .A2( u0_u9_u2_n107 ) , .ZN( u0_u9_u2_n139 ) );
  NAND2_X1 u0_u9_u2_U59 (.A1( u0_u9_u2_n103 ) , .A2( u0_u9_u2_n105 ) , .ZN( u0_u9_u2_n133 ) );
  AOI21_X1 u0_u9_u2_U6 (.B2( u0_u9_u2_n119 ) , .ZN( u0_u9_u2_n127 ) , .A( u0_u9_u2_n137 ) , .B1( u0_u9_u2_n155 ) );
  NAND2_X1 u0_u9_u2_U60 (.A1( u0_u9_u2_n102 ) , .A2( u0_u9_u2_n103 ) , .ZN( u0_u9_u2_n154 ) );
  NAND2_X1 u0_u9_u2_U61 (.A2( u0_u9_u2_n103 ) , .A1( u0_u9_u2_n104 ) , .ZN( u0_u9_u2_n119 ) );
  NAND2_X1 u0_u9_u2_U62 (.A2( u0_u9_u2_n107 ) , .A1( u0_u9_u2_n108 ) , .ZN( u0_u9_u2_n123 ) );
  NAND2_X1 u0_u9_u2_U63 (.A1( u0_u9_u2_n104 ) , .A2( u0_u9_u2_n108 ) , .ZN( u0_u9_u2_n122 ) );
  INV_X1 u0_u9_u2_U64 (.A( u0_u9_u2_n114 ) , .ZN( u0_u9_u2_n172 ) );
  NAND2_X1 u0_u9_u2_U65 (.A2( u0_u9_u2_n100 ) , .A1( u0_u9_u2_n102 ) , .ZN( u0_u9_u2_n116 ) );
  NAND2_X1 u0_u9_u2_U66 (.A1( u0_u9_u2_n102 ) , .A2( u0_u9_u2_n108 ) , .ZN( u0_u9_u2_n120 ) );
  NAND2_X1 u0_u9_u2_U67 (.A2( u0_u9_u2_n105 ) , .A1( u0_u9_u2_n106 ) , .ZN( u0_u9_u2_n117 ) );
  INV_X1 u0_u9_u2_U68 (.ZN( u0_u9_u2_n187 ) , .A( u0_u9_u2_n99 ) );
  OAI21_X1 u0_u9_u2_U69 (.B1( u0_u9_u2_n137 ) , .B2( u0_u9_u2_n143 ) , .A( u0_u9_u2_n98 ) , .ZN( u0_u9_u2_n99 ) );
  AOI21_X1 u0_u9_u2_U7 (.ZN( u0_u9_u2_n124 ) , .B1( u0_u9_u2_n131 ) , .B2( u0_u9_u2_n143 ) , .A( u0_u9_u2_n172 ) );
  NOR2_X1 u0_u9_u2_U70 (.A2( u0_u9_X_16 ) , .ZN( u0_u9_u2_n140 ) , .A1( u0_u9_u2_n166 ) );
  NOR2_X1 u0_u9_u2_U71 (.A2( u0_u9_X_13 ) , .A1( u0_u9_X_14 ) , .ZN( u0_u9_u2_n100 ) );
  NOR2_X1 u0_u9_u2_U72 (.A2( u0_u9_X_16 ) , .A1( u0_u9_X_17 ) , .ZN( u0_u9_u2_n138 ) );
  NOR2_X1 u0_u9_u2_U73 (.A2( u0_u9_X_15 ) , .A1( u0_u9_X_18 ) , .ZN( u0_u9_u2_n104 ) );
  NOR2_X1 u0_u9_u2_U74 (.A2( u0_u9_X_14 ) , .ZN( u0_u9_u2_n103 ) , .A1( u0_u9_u2_n174 ) );
  NOR2_X1 u0_u9_u2_U75 (.A2( u0_u9_X_15 ) , .ZN( u0_u9_u2_n102 ) , .A1( u0_u9_u2_n165 ) );
  NOR2_X1 u0_u9_u2_U76 (.A2( u0_u9_X_17 ) , .ZN( u0_u9_u2_n114 ) , .A1( u0_u9_u2_n169 ) );
  AND2_X1 u0_u9_u2_U77 (.A1( u0_u9_X_15 ) , .ZN( u0_u9_u2_n105 ) , .A2( u0_u9_u2_n165 ) );
  AND2_X1 u0_u9_u2_U78 (.A2( u0_u9_X_15 ) , .A1( u0_u9_X_18 ) , .ZN( u0_u9_u2_n107 ) );
  AND2_X1 u0_u9_u2_U79 (.A1( u0_u9_X_14 ) , .ZN( u0_u9_u2_n106 ) , .A2( u0_u9_u2_n174 ) );
  AOI21_X1 u0_u9_u2_U8 (.B2( u0_u9_u2_n120 ) , .B1( u0_u9_u2_n121 ) , .ZN( u0_u9_u2_n126 ) , .A( u0_u9_u2_n167 ) );
  AND2_X1 u0_u9_u2_U80 (.A1( u0_u9_X_13 ) , .A2( u0_u9_X_14 ) , .ZN( u0_u9_u2_n108 ) );
  INV_X1 u0_u9_u2_U81 (.A( u0_u9_X_16 ) , .ZN( u0_u9_u2_n169 ) );
  INV_X1 u0_u9_u2_U82 (.A( u0_u9_X_17 ) , .ZN( u0_u9_u2_n166 ) );
  INV_X1 u0_u9_u2_U83 (.A( u0_u9_X_13 ) , .ZN( u0_u9_u2_n174 ) );
  INV_X1 u0_u9_u2_U84 (.A( u0_u9_X_18 ) , .ZN( u0_u9_u2_n165 ) );
  NAND4_X1 u0_u9_u2_U85 (.ZN( u0_out9_30 ) , .A4( u0_u9_u2_n147 ) , .A3( u0_u9_u2_n148 ) , .A2( u0_u9_u2_n149 ) , .A1( u0_u9_u2_n187 ) );
  AOI21_X1 u0_u9_u2_U86 (.B2( u0_u9_u2_n138 ) , .ZN( u0_u9_u2_n148 ) , .A( u0_u9_u2_n162 ) , .B1( u0_u9_u2_n182 ) );
  NOR3_X1 u0_u9_u2_U87 (.A3( u0_u9_u2_n144 ) , .A2( u0_u9_u2_n145 ) , .A1( u0_u9_u2_n146 ) , .ZN( u0_u9_u2_n147 ) );
  NAND4_X1 u0_u9_u2_U88 (.ZN( u0_out9_24 ) , .A4( u0_u9_u2_n111 ) , .A3( u0_u9_u2_n112 ) , .A1( u0_u9_u2_n130 ) , .A2( u0_u9_u2_n187 ) );
  AOI221_X1 u0_u9_u2_U89 (.A( u0_u9_u2_n109 ) , .B1( u0_u9_u2_n110 ) , .ZN( u0_u9_u2_n111 ) , .C1( u0_u9_u2_n134 ) , .C2( u0_u9_u2_n170 ) , .B2( u0_u9_u2_n173 ) );
  OAI22_X1 u0_u9_u2_U9 (.ZN( u0_u9_u2_n109 ) , .A2( u0_u9_u2_n113 ) , .B2( u0_u9_u2_n133 ) , .B1( u0_u9_u2_n167 ) , .A1( u0_u9_u2_n168 ) );
  AOI21_X1 u0_u9_u2_U90 (.ZN( u0_u9_u2_n112 ) , .B2( u0_u9_u2_n156 ) , .A( u0_u9_u2_n164 ) , .B1( u0_u9_u2_n181 ) );
  NAND4_X1 u0_u9_u2_U91 (.ZN( u0_out9_16 ) , .A4( u0_u9_u2_n128 ) , .A3( u0_u9_u2_n129 ) , .A1( u0_u9_u2_n130 ) , .A2( u0_u9_u2_n186 ) );
  AOI22_X1 u0_u9_u2_U92 (.A2( u0_u9_u2_n118 ) , .ZN( u0_u9_u2_n129 ) , .A1( u0_u9_u2_n140 ) , .B1( u0_u9_u2_n157 ) , .B2( u0_u9_u2_n170 ) );
  INV_X1 u0_u9_u2_U93 (.A( u0_u9_u2_n163 ) , .ZN( u0_u9_u2_n186 ) );
  OR4_X1 u0_u9_u2_U94 (.ZN( u0_out9_6 ) , .A4( u0_u9_u2_n161 ) , .A3( u0_u9_u2_n162 ) , .A2( u0_u9_u2_n163 ) , .A1( u0_u9_u2_n164 ) );
  OR3_X1 u0_u9_u2_U95 (.A2( u0_u9_u2_n159 ) , .A1( u0_u9_u2_n160 ) , .ZN( u0_u9_u2_n161 ) , .A3( u0_u9_u2_n183 ) );
  AOI21_X1 u0_u9_u2_U96 (.B2( u0_u9_u2_n154 ) , .B1( u0_u9_u2_n155 ) , .ZN( u0_u9_u2_n159 ) , .A( u0_u9_u2_n167 ) );
  NAND3_X1 u0_u9_u2_U97 (.A2( u0_u9_u2_n117 ) , .A1( u0_u9_u2_n122 ) , .A3( u0_u9_u2_n123 ) , .ZN( u0_u9_u2_n134 ) );
  NAND3_X1 u0_u9_u2_U98 (.ZN( u0_u9_u2_n110 ) , .A2( u0_u9_u2_n131 ) , .A3( u0_u9_u2_n139 ) , .A1( u0_u9_u2_n154 ) );
  NAND3_X1 u0_u9_u2_U99 (.A2( u0_u9_u2_n100 ) , .ZN( u0_u9_u2_n101 ) , .A1( u0_u9_u2_n104 ) , .A3( u0_u9_u2_n114 ) );
  OAI22_X1 u0_u9_u3_U10 (.B1( u0_u9_u3_n113 ) , .A2( u0_u9_u3_n135 ) , .A1( u0_u9_u3_n150 ) , .B2( u0_u9_u3_n164 ) , .ZN( u0_u9_u3_n98 ) );
  OAI211_X1 u0_u9_u3_U11 (.B( u0_u9_u3_n106 ) , .ZN( u0_u9_u3_n119 ) , .C2( u0_u9_u3_n128 ) , .C1( u0_u9_u3_n167 ) , .A( u0_u9_u3_n181 ) );
  AOI221_X1 u0_u9_u3_U12 (.C1( u0_u9_u3_n105 ) , .ZN( u0_u9_u3_n106 ) , .A( u0_u9_u3_n131 ) , .B2( u0_u9_u3_n132 ) , .C2( u0_u9_u3_n133 ) , .B1( u0_u9_u3_n169 ) );
  INV_X1 u0_u9_u3_U13 (.ZN( u0_u9_u3_n181 ) , .A( u0_u9_u3_n98 ) );
  NAND2_X1 u0_u9_u3_U14 (.ZN( u0_u9_u3_n105 ) , .A2( u0_u9_u3_n130 ) , .A1( u0_u9_u3_n155 ) );
  AOI22_X1 u0_u9_u3_U15 (.B1( u0_u9_u3_n115 ) , .A2( u0_u9_u3_n116 ) , .ZN( u0_u9_u3_n123 ) , .B2( u0_u9_u3_n133 ) , .A1( u0_u9_u3_n169 ) );
  NAND2_X1 u0_u9_u3_U16 (.ZN( u0_u9_u3_n116 ) , .A2( u0_u9_u3_n151 ) , .A1( u0_u9_u3_n182 ) );
  NOR2_X1 u0_u9_u3_U17 (.ZN( u0_u9_u3_n126 ) , .A2( u0_u9_u3_n150 ) , .A1( u0_u9_u3_n164 ) );
  AOI21_X1 u0_u9_u3_U18 (.ZN( u0_u9_u3_n112 ) , .B2( u0_u9_u3_n146 ) , .B1( u0_u9_u3_n155 ) , .A( u0_u9_u3_n167 ) );
  NAND2_X1 u0_u9_u3_U19 (.A1( u0_u9_u3_n135 ) , .ZN( u0_u9_u3_n142 ) , .A2( u0_u9_u3_n164 ) );
  NAND2_X1 u0_u9_u3_U20 (.ZN( u0_u9_u3_n132 ) , .A2( u0_u9_u3_n152 ) , .A1( u0_u9_u3_n156 ) );
  AND2_X1 u0_u9_u3_U21 (.A2( u0_u9_u3_n113 ) , .A1( u0_u9_u3_n114 ) , .ZN( u0_u9_u3_n151 ) );
  INV_X1 u0_u9_u3_U22 (.A( u0_u9_u3_n133 ) , .ZN( u0_u9_u3_n165 ) );
  INV_X1 u0_u9_u3_U23 (.A( u0_u9_u3_n135 ) , .ZN( u0_u9_u3_n170 ) );
  NAND2_X1 u0_u9_u3_U24 (.A1( u0_u9_u3_n107 ) , .A2( u0_u9_u3_n108 ) , .ZN( u0_u9_u3_n140 ) );
  NAND2_X1 u0_u9_u3_U25 (.ZN( u0_u9_u3_n117 ) , .A1( u0_u9_u3_n124 ) , .A2( u0_u9_u3_n148 ) );
  NAND2_X1 u0_u9_u3_U26 (.ZN( u0_u9_u3_n143 ) , .A1( u0_u9_u3_n165 ) , .A2( u0_u9_u3_n167 ) );
  INV_X1 u0_u9_u3_U27 (.A( u0_u9_u3_n130 ) , .ZN( u0_u9_u3_n177 ) );
  INV_X1 u0_u9_u3_U28 (.A( u0_u9_u3_n128 ) , .ZN( u0_u9_u3_n176 ) );
  INV_X1 u0_u9_u3_U29 (.A( u0_u9_u3_n155 ) , .ZN( u0_u9_u3_n174 ) );
  INV_X1 u0_u9_u3_U3 (.A( u0_u9_u3_n129 ) , .ZN( u0_u9_u3_n183 ) );
  INV_X1 u0_u9_u3_U30 (.A( u0_u9_u3_n139 ) , .ZN( u0_u9_u3_n185 ) );
  NOR2_X1 u0_u9_u3_U31 (.ZN( u0_u9_u3_n135 ) , .A2( u0_u9_u3_n141 ) , .A1( u0_u9_u3_n169 ) );
  OAI222_X1 u0_u9_u3_U32 (.C2( u0_u9_u3_n107 ) , .A2( u0_u9_u3_n108 ) , .B1( u0_u9_u3_n135 ) , .ZN( u0_u9_u3_n138 ) , .B2( u0_u9_u3_n146 ) , .C1( u0_u9_u3_n154 ) , .A1( u0_u9_u3_n164 ) );
  NOR4_X1 u0_u9_u3_U33 (.A4( u0_u9_u3_n157 ) , .A3( u0_u9_u3_n158 ) , .A2( u0_u9_u3_n159 ) , .A1( u0_u9_u3_n160 ) , .ZN( u0_u9_u3_n161 ) );
  AOI21_X1 u0_u9_u3_U34 (.B2( u0_u9_u3_n152 ) , .B1( u0_u9_u3_n153 ) , .ZN( u0_u9_u3_n158 ) , .A( u0_u9_u3_n164 ) );
  AOI21_X1 u0_u9_u3_U35 (.A( u0_u9_u3_n154 ) , .B2( u0_u9_u3_n155 ) , .B1( u0_u9_u3_n156 ) , .ZN( u0_u9_u3_n157 ) );
  AOI21_X1 u0_u9_u3_U36 (.A( u0_u9_u3_n149 ) , .B2( u0_u9_u3_n150 ) , .B1( u0_u9_u3_n151 ) , .ZN( u0_u9_u3_n159 ) );
  AOI211_X1 u0_u9_u3_U37 (.ZN( u0_u9_u3_n109 ) , .A( u0_u9_u3_n119 ) , .C2( u0_u9_u3_n129 ) , .B( u0_u9_u3_n138 ) , .C1( u0_u9_u3_n141 ) );
  AOI211_X1 u0_u9_u3_U38 (.B( u0_u9_u3_n119 ) , .A( u0_u9_u3_n120 ) , .C2( u0_u9_u3_n121 ) , .ZN( u0_u9_u3_n122 ) , .C1( u0_u9_u3_n179 ) );
  INV_X1 u0_u9_u3_U39 (.A( u0_u9_u3_n156 ) , .ZN( u0_u9_u3_n179 ) );
  INV_X1 u0_u9_u3_U4 (.A( u0_u9_u3_n140 ) , .ZN( u0_u9_u3_n182 ) );
  OAI22_X1 u0_u9_u3_U40 (.B1( u0_u9_u3_n118 ) , .ZN( u0_u9_u3_n120 ) , .A1( u0_u9_u3_n135 ) , .B2( u0_u9_u3_n154 ) , .A2( u0_u9_u3_n178 ) );
  AND3_X1 u0_u9_u3_U41 (.ZN( u0_u9_u3_n118 ) , .A2( u0_u9_u3_n124 ) , .A1( u0_u9_u3_n144 ) , .A3( u0_u9_u3_n152 ) );
  INV_X1 u0_u9_u3_U42 (.A( u0_u9_u3_n121 ) , .ZN( u0_u9_u3_n164 ) );
  NAND2_X1 u0_u9_u3_U43 (.ZN( u0_u9_u3_n133 ) , .A1( u0_u9_u3_n154 ) , .A2( u0_u9_u3_n164 ) );
  OAI211_X1 u0_u9_u3_U44 (.B( u0_u9_u3_n127 ) , .ZN( u0_u9_u3_n139 ) , .C1( u0_u9_u3_n150 ) , .C2( u0_u9_u3_n154 ) , .A( u0_u9_u3_n184 ) );
  INV_X1 u0_u9_u3_U45 (.A( u0_u9_u3_n125 ) , .ZN( u0_u9_u3_n184 ) );
  AOI221_X1 u0_u9_u3_U46 (.A( u0_u9_u3_n126 ) , .ZN( u0_u9_u3_n127 ) , .C2( u0_u9_u3_n132 ) , .C1( u0_u9_u3_n169 ) , .B2( u0_u9_u3_n170 ) , .B1( u0_u9_u3_n174 ) );
  OAI22_X1 u0_u9_u3_U47 (.A1( u0_u9_u3_n124 ) , .ZN( u0_u9_u3_n125 ) , .B2( u0_u9_u3_n145 ) , .A2( u0_u9_u3_n165 ) , .B1( u0_u9_u3_n167 ) );
  NOR2_X1 u0_u9_u3_U48 (.A1( u0_u9_u3_n113 ) , .ZN( u0_u9_u3_n131 ) , .A2( u0_u9_u3_n154 ) );
  NAND2_X1 u0_u9_u3_U49 (.A1( u0_u9_u3_n103 ) , .ZN( u0_u9_u3_n150 ) , .A2( u0_u9_u3_n99 ) );
  INV_X1 u0_u9_u3_U5 (.A( u0_u9_u3_n117 ) , .ZN( u0_u9_u3_n178 ) );
  NAND2_X1 u0_u9_u3_U50 (.A2( u0_u9_u3_n102 ) , .ZN( u0_u9_u3_n155 ) , .A1( u0_u9_u3_n97 ) );
  INV_X1 u0_u9_u3_U51 (.A( u0_u9_u3_n141 ) , .ZN( u0_u9_u3_n167 ) );
  AOI21_X1 u0_u9_u3_U52 (.B2( u0_u9_u3_n114 ) , .B1( u0_u9_u3_n146 ) , .A( u0_u9_u3_n154 ) , .ZN( u0_u9_u3_n94 ) );
  AOI21_X1 u0_u9_u3_U53 (.ZN( u0_u9_u3_n110 ) , .B2( u0_u9_u3_n142 ) , .B1( u0_u9_u3_n186 ) , .A( u0_u9_u3_n95 ) );
  INV_X1 u0_u9_u3_U54 (.A( u0_u9_u3_n145 ) , .ZN( u0_u9_u3_n186 ) );
  AOI21_X1 u0_u9_u3_U55 (.B1( u0_u9_u3_n124 ) , .A( u0_u9_u3_n149 ) , .B2( u0_u9_u3_n155 ) , .ZN( u0_u9_u3_n95 ) );
  INV_X1 u0_u9_u3_U56 (.A( u0_u9_u3_n149 ) , .ZN( u0_u9_u3_n169 ) );
  NAND2_X1 u0_u9_u3_U57 (.ZN( u0_u9_u3_n124 ) , .A1( u0_u9_u3_n96 ) , .A2( u0_u9_u3_n97 ) );
  NAND2_X1 u0_u9_u3_U58 (.A2( u0_u9_u3_n100 ) , .ZN( u0_u9_u3_n146 ) , .A1( u0_u9_u3_n96 ) );
  NAND2_X1 u0_u9_u3_U59 (.A1( u0_u9_u3_n101 ) , .ZN( u0_u9_u3_n145 ) , .A2( u0_u9_u3_n99 ) );
  AOI221_X1 u0_u9_u3_U6 (.A( u0_u9_u3_n131 ) , .C2( u0_u9_u3_n132 ) , .C1( u0_u9_u3_n133 ) , .ZN( u0_u9_u3_n134 ) , .B1( u0_u9_u3_n143 ) , .B2( u0_u9_u3_n177 ) );
  NAND2_X1 u0_u9_u3_U60 (.A1( u0_u9_u3_n100 ) , .ZN( u0_u9_u3_n156 ) , .A2( u0_u9_u3_n99 ) );
  NAND2_X1 u0_u9_u3_U61 (.A2( u0_u9_u3_n101 ) , .A1( u0_u9_u3_n104 ) , .ZN( u0_u9_u3_n148 ) );
  NAND2_X1 u0_u9_u3_U62 (.A1( u0_u9_u3_n100 ) , .A2( u0_u9_u3_n102 ) , .ZN( u0_u9_u3_n128 ) );
  NAND2_X1 u0_u9_u3_U63 (.A2( u0_u9_u3_n101 ) , .A1( u0_u9_u3_n102 ) , .ZN( u0_u9_u3_n152 ) );
  NAND2_X1 u0_u9_u3_U64 (.A2( u0_u9_u3_n101 ) , .ZN( u0_u9_u3_n114 ) , .A1( u0_u9_u3_n96 ) );
  NAND2_X1 u0_u9_u3_U65 (.ZN( u0_u9_u3_n107 ) , .A1( u0_u9_u3_n97 ) , .A2( u0_u9_u3_n99 ) );
  NAND2_X1 u0_u9_u3_U66 (.A2( u0_u9_u3_n100 ) , .A1( u0_u9_u3_n104 ) , .ZN( u0_u9_u3_n113 ) );
  NAND2_X1 u0_u9_u3_U67 (.A1( u0_u9_u3_n104 ) , .ZN( u0_u9_u3_n153 ) , .A2( u0_u9_u3_n97 ) );
  NAND2_X1 u0_u9_u3_U68 (.A2( u0_u9_u3_n103 ) , .A1( u0_u9_u3_n104 ) , .ZN( u0_u9_u3_n130 ) );
  NAND2_X1 u0_u9_u3_U69 (.A2( u0_u9_u3_n103 ) , .ZN( u0_u9_u3_n144 ) , .A1( u0_u9_u3_n96 ) );
  OAI22_X1 u0_u9_u3_U7 (.B2( u0_u9_u3_n147 ) , .A2( u0_u9_u3_n148 ) , .ZN( u0_u9_u3_n160 ) , .B1( u0_u9_u3_n165 ) , .A1( u0_u9_u3_n168 ) );
  NAND2_X1 u0_u9_u3_U70 (.A1( u0_u9_u3_n102 ) , .A2( u0_u9_u3_n103 ) , .ZN( u0_u9_u3_n108 ) );
  NOR2_X1 u0_u9_u3_U71 (.A2( u0_u9_X_19 ) , .A1( u0_u9_X_20 ) , .ZN( u0_u9_u3_n99 ) );
  NOR2_X1 u0_u9_u3_U72 (.A2( u0_u9_X_21 ) , .A1( u0_u9_X_24 ) , .ZN( u0_u9_u3_n103 ) );
  NOR2_X1 u0_u9_u3_U73 (.A2( u0_u9_X_24 ) , .A1( u0_u9_u3_n171 ) , .ZN( u0_u9_u3_n97 ) );
  NOR2_X1 u0_u9_u3_U74 (.A2( u0_u9_X_23 ) , .ZN( u0_u9_u3_n141 ) , .A1( u0_u9_u3_n166 ) );
  NOR2_X1 u0_u9_u3_U75 (.A2( u0_u9_X_19 ) , .A1( u0_u9_u3_n172 ) , .ZN( u0_u9_u3_n96 ) );
  NAND2_X1 u0_u9_u3_U76 (.A1( u0_u9_X_22 ) , .A2( u0_u9_X_23 ) , .ZN( u0_u9_u3_n154 ) );
  NAND2_X1 u0_u9_u3_U77 (.A1( u0_u9_X_23 ) , .ZN( u0_u9_u3_n149 ) , .A2( u0_u9_u3_n166 ) );
  NOR2_X1 u0_u9_u3_U78 (.A2( u0_u9_X_22 ) , .A1( u0_u9_X_23 ) , .ZN( u0_u9_u3_n121 ) );
  AND2_X1 u0_u9_u3_U79 (.A1( u0_u9_X_24 ) , .ZN( u0_u9_u3_n101 ) , .A2( u0_u9_u3_n171 ) );
  AND3_X1 u0_u9_u3_U8 (.A3( u0_u9_u3_n144 ) , .A2( u0_u9_u3_n145 ) , .A1( u0_u9_u3_n146 ) , .ZN( u0_u9_u3_n147 ) );
  AND2_X1 u0_u9_u3_U80 (.A1( u0_u9_X_19 ) , .ZN( u0_u9_u3_n102 ) , .A2( u0_u9_u3_n172 ) );
  AND2_X1 u0_u9_u3_U81 (.A1( u0_u9_X_21 ) , .A2( u0_u9_X_24 ) , .ZN( u0_u9_u3_n100 ) );
  AND2_X1 u0_u9_u3_U82 (.A2( u0_u9_X_19 ) , .A1( u0_u9_X_20 ) , .ZN( u0_u9_u3_n104 ) );
  INV_X1 u0_u9_u3_U83 (.A( u0_u9_X_22 ) , .ZN( u0_u9_u3_n166 ) );
  INV_X1 u0_u9_u3_U84 (.A( u0_u9_X_21 ) , .ZN( u0_u9_u3_n171 ) );
  INV_X1 u0_u9_u3_U85 (.A( u0_u9_X_20 ) , .ZN( u0_u9_u3_n172 ) );
  OR4_X1 u0_u9_u3_U86 (.ZN( u0_out9_10 ) , .A4( u0_u9_u3_n136 ) , .A3( u0_u9_u3_n137 ) , .A1( u0_u9_u3_n138 ) , .A2( u0_u9_u3_n139 ) );
  OAI222_X1 u0_u9_u3_U87 (.C1( u0_u9_u3_n128 ) , .ZN( u0_u9_u3_n137 ) , .B1( u0_u9_u3_n148 ) , .A2( u0_u9_u3_n150 ) , .B2( u0_u9_u3_n154 ) , .C2( u0_u9_u3_n164 ) , .A1( u0_u9_u3_n167 ) );
  OAI221_X1 u0_u9_u3_U88 (.A( u0_u9_u3_n134 ) , .B2( u0_u9_u3_n135 ) , .ZN( u0_u9_u3_n136 ) , .C1( u0_u9_u3_n149 ) , .B1( u0_u9_u3_n151 ) , .C2( u0_u9_u3_n183 ) );
  NAND4_X1 u0_u9_u3_U89 (.ZN( u0_out9_26 ) , .A4( u0_u9_u3_n109 ) , .A3( u0_u9_u3_n110 ) , .A2( u0_u9_u3_n111 ) , .A1( u0_u9_u3_n173 ) );
  INV_X1 u0_u9_u3_U9 (.A( u0_u9_u3_n143 ) , .ZN( u0_u9_u3_n168 ) );
  INV_X1 u0_u9_u3_U90 (.ZN( u0_u9_u3_n173 ) , .A( u0_u9_u3_n94 ) );
  OAI21_X1 u0_u9_u3_U91 (.ZN( u0_u9_u3_n111 ) , .B2( u0_u9_u3_n117 ) , .A( u0_u9_u3_n133 ) , .B1( u0_u9_u3_n176 ) );
  NAND4_X1 u0_u9_u3_U92 (.ZN( u0_out9_20 ) , .A4( u0_u9_u3_n122 ) , .A3( u0_u9_u3_n123 ) , .A1( u0_u9_u3_n175 ) , .A2( u0_u9_u3_n180 ) );
  INV_X1 u0_u9_u3_U93 (.A( u0_u9_u3_n126 ) , .ZN( u0_u9_u3_n180 ) );
  INV_X1 u0_u9_u3_U94 (.A( u0_u9_u3_n112 ) , .ZN( u0_u9_u3_n175 ) );
  NAND4_X1 u0_u9_u3_U95 (.ZN( u0_out9_1 ) , .A4( u0_u9_u3_n161 ) , .A3( u0_u9_u3_n162 ) , .A2( u0_u9_u3_n163 ) , .A1( u0_u9_u3_n185 ) );
  NAND2_X1 u0_u9_u3_U96 (.ZN( u0_u9_u3_n163 ) , .A2( u0_u9_u3_n170 ) , .A1( u0_u9_u3_n176 ) );
  AOI22_X1 u0_u9_u3_U97 (.B2( u0_u9_u3_n140 ) , .B1( u0_u9_u3_n141 ) , .A2( u0_u9_u3_n142 ) , .ZN( u0_u9_u3_n162 ) , .A1( u0_u9_u3_n177 ) );
  NAND3_X1 u0_u9_u3_U98 (.A1( u0_u9_u3_n114 ) , .ZN( u0_u9_u3_n115 ) , .A2( u0_u9_u3_n145 ) , .A3( u0_u9_u3_n153 ) );
  NAND3_X1 u0_u9_u3_U99 (.ZN( u0_u9_u3_n129 ) , .A2( u0_u9_u3_n144 ) , .A1( u0_u9_u3_n153 ) , .A3( u0_u9_u3_n182 ) );
  OAI22_X1 u0_u9_u4_U10 (.B2( u0_u9_u4_n135 ) , .ZN( u0_u9_u4_n137 ) , .B1( u0_u9_u4_n153 ) , .A1( u0_u9_u4_n155 ) , .A2( u0_u9_u4_n171 ) );
  AND3_X1 u0_u9_u4_U11 (.A2( u0_u9_u4_n134 ) , .ZN( u0_u9_u4_n135 ) , .A3( u0_u9_u4_n145 ) , .A1( u0_u9_u4_n157 ) );
  NAND2_X1 u0_u9_u4_U12 (.ZN( u0_u9_u4_n132 ) , .A2( u0_u9_u4_n170 ) , .A1( u0_u9_u4_n173 ) );
  AOI21_X1 u0_u9_u4_U13 (.B2( u0_u9_u4_n160 ) , .B1( u0_u9_u4_n161 ) , .ZN( u0_u9_u4_n162 ) , .A( u0_u9_u4_n170 ) );
  AOI21_X1 u0_u9_u4_U14 (.ZN( u0_u9_u4_n107 ) , .B2( u0_u9_u4_n143 ) , .A( u0_u9_u4_n174 ) , .B1( u0_u9_u4_n184 ) );
  AOI21_X1 u0_u9_u4_U15 (.B2( u0_u9_u4_n158 ) , .B1( u0_u9_u4_n159 ) , .ZN( u0_u9_u4_n163 ) , .A( u0_u9_u4_n174 ) );
  AOI21_X1 u0_u9_u4_U16 (.A( u0_u9_u4_n153 ) , .B2( u0_u9_u4_n154 ) , .B1( u0_u9_u4_n155 ) , .ZN( u0_u9_u4_n165 ) );
  AOI21_X1 u0_u9_u4_U17 (.A( u0_u9_u4_n156 ) , .B2( u0_u9_u4_n157 ) , .ZN( u0_u9_u4_n164 ) , .B1( u0_u9_u4_n184 ) );
  INV_X1 u0_u9_u4_U18 (.A( u0_u9_u4_n138 ) , .ZN( u0_u9_u4_n170 ) );
  AND2_X1 u0_u9_u4_U19 (.A2( u0_u9_u4_n120 ) , .ZN( u0_u9_u4_n155 ) , .A1( u0_u9_u4_n160 ) );
  INV_X1 u0_u9_u4_U20 (.A( u0_u9_u4_n156 ) , .ZN( u0_u9_u4_n175 ) );
  NAND2_X1 u0_u9_u4_U21 (.A2( u0_u9_u4_n118 ) , .ZN( u0_u9_u4_n131 ) , .A1( u0_u9_u4_n147 ) );
  NAND2_X1 u0_u9_u4_U22 (.A1( u0_u9_u4_n119 ) , .A2( u0_u9_u4_n120 ) , .ZN( u0_u9_u4_n130 ) );
  NAND2_X1 u0_u9_u4_U23 (.ZN( u0_u9_u4_n117 ) , .A2( u0_u9_u4_n118 ) , .A1( u0_u9_u4_n148 ) );
  NAND2_X1 u0_u9_u4_U24 (.ZN( u0_u9_u4_n129 ) , .A1( u0_u9_u4_n134 ) , .A2( u0_u9_u4_n148 ) );
  AND3_X1 u0_u9_u4_U25 (.A1( u0_u9_u4_n119 ) , .A2( u0_u9_u4_n143 ) , .A3( u0_u9_u4_n154 ) , .ZN( u0_u9_u4_n161 ) );
  AND2_X1 u0_u9_u4_U26 (.A1( u0_u9_u4_n145 ) , .A2( u0_u9_u4_n147 ) , .ZN( u0_u9_u4_n159 ) );
  OR3_X1 u0_u9_u4_U27 (.A3( u0_u9_u4_n114 ) , .A2( u0_u9_u4_n115 ) , .A1( u0_u9_u4_n116 ) , .ZN( u0_u9_u4_n136 ) );
  AOI21_X1 u0_u9_u4_U28 (.A( u0_u9_u4_n113 ) , .ZN( u0_u9_u4_n116 ) , .B2( u0_u9_u4_n173 ) , .B1( u0_u9_u4_n174 ) );
  AOI21_X1 u0_u9_u4_U29 (.ZN( u0_u9_u4_n115 ) , .B2( u0_u9_u4_n145 ) , .B1( u0_u9_u4_n146 ) , .A( u0_u9_u4_n156 ) );
  NOR2_X1 u0_u9_u4_U3 (.ZN( u0_u9_u4_n121 ) , .A1( u0_u9_u4_n181 ) , .A2( u0_u9_u4_n182 ) );
  OAI22_X1 u0_u9_u4_U30 (.ZN( u0_u9_u4_n114 ) , .A2( u0_u9_u4_n121 ) , .B1( u0_u9_u4_n160 ) , .B2( u0_u9_u4_n170 ) , .A1( u0_u9_u4_n171 ) );
  INV_X1 u0_u9_u4_U31 (.A( u0_u9_u4_n158 ) , .ZN( u0_u9_u4_n182 ) );
  INV_X1 u0_u9_u4_U32 (.ZN( u0_u9_u4_n181 ) , .A( u0_u9_u4_n96 ) );
  INV_X1 u0_u9_u4_U33 (.A( u0_u9_u4_n144 ) , .ZN( u0_u9_u4_n179 ) );
  INV_X1 u0_u9_u4_U34 (.A( u0_u9_u4_n157 ) , .ZN( u0_u9_u4_n178 ) );
  NAND2_X1 u0_u9_u4_U35 (.A2( u0_u9_u4_n154 ) , .A1( u0_u9_u4_n96 ) , .ZN( u0_u9_u4_n97 ) );
  INV_X1 u0_u9_u4_U36 (.ZN( u0_u9_u4_n186 ) , .A( u0_u9_u4_n95 ) );
  OAI221_X1 u0_u9_u4_U37 (.C1( u0_u9_u4_n134 ) , .B1( u0_u9_u4_n158 ) , .B2( u0_u9_u4_n171 ) , .C2( u0_u9_u4_n173 ) , .A( u0_u9_u4_n94 ) , .ZN( u0_u9_u4_n95 ) );
  AOI222_X1 u0_u9_u4_U38 (.B2( u0_u9_u4_n132 ) , .A1( u0_u9_u4_n138 ) , .C2( u0_u9_u4_n175 ) , .A2( u0_u9_u4_n179 ) , .C1( u0_u9_u4_n181 ) , .B1( u0_u9_u4_n185 ) , .ZN( u0_u9_u4_n94 ) );
  INV_X1 u0_u9_u4_U39 (.A( u0_u9_u4_n113 ) , .ZN( u0_u9_u4_n185 ) );
  INV_X1 u0_u9_u4_U4 (.A( u0_u9_u4_n117 ) , .ZN( u0_u9_u4_n184 ) );
  INV_X1 u0_u9_u4_U40 (.A( u0_u9_u4_n143 ) , .ZN( u0_u9_u4_n183 ) );
  NOR2_X1 u0_u9_u4_U41 (.ZN( u0_u9_u4_n138 ) , .A1( u0_u9_u4_n168 ) , .A2( u0_u9_u4_n169 ) );
  NOR2_X1 u0_u9_u4_U42 (.A1( u0_u9_u4_n150 ) , .A2( u0_u9_u4_n152 ) , .ZN( u0_u9_u4_n153 ) );
  NOR2_X1 u0_u9_u4_U43 (.A2( u0_u9_u4_n128 ) , .A1( u0_u9_u4_n138 ) , .ZN( u0_u9_u4_n156 ) );
  AOI22_X1 u0_u9_u4_U44 (.B2( u0_u9_u4_n122 ) , .A1( u0_u9_u4_n123 ) , .ZN( u0_u9_u4_n124 ) , .B1( u0_u9_u4_n128 ) , .A2( u0_u9_u4_n172 ) );
  INV_X1 u0_u9_u4_U45 (.A( u0_u9_u4_n153 ) , .ZN( u0_u9_u4_n172 ) );
  NAND2_X1 u0_u9_u4_U46 (.A2( u0_u9_u4_n120 ) , .ZN( u0_u9_u4_n123 ) , .A1( u0_u9_u4_n161 ) );
  AOI22_X1 u0_u9_u4_U47 (.B2( u0_u9_u4_n132 ) , .A2( u0_u9_u4_n133 ) , .ZN( u0_u9_u4_n140 ) , .A1( u0_u9_u4_n150 ) , .B1( u0_u9_u4_n179 ) );
  NAND2_X1 u0_u9_u4_U48 (.ZN( u0_u9_u4_n133 ) , .A2( u0_u9_u4_n146 ) , .A1( u0_u9_u4_n154 ) );
  NAND2_X1 u0_u9_u4_U49 (.A1( u0_u9_u4_n103 ) , .ZN( u0_u9_u4_n154 ) , .A2( u0_u9_u4_n98 ) );
  NOR4_X1 u0_u9_u4_U5 (.A4( u0_u9_u4_n106 ) , .A3( u0_u9_u4_n107 ) , .A2( u0_u9_u4_n108 ) , .A1( u0_u9_u4_n109 ) , .ZN( u0_u9_u4_n110 ) );
  NAND2_X1 u0_u9_u4_U50 (.A1( u0_u9_u4_n101 ) , .ZN( u0_u9_u4_n158 ) , .A2( u0_u9_u4_n99 ) );
  AOI21_X1 u0_u9_u4_U51 (.ZN( u0_u9_u4_n127 ) , .A( u0_u9_u4_n136 ) , .B2( u0_u9_u4_n150 ) , .B1( u0_u9_u4_n180 ) );
  INV_X1 u0_u9_u4_U52 (.A( u0_u9_u4_n160 ) , .ZN( u0_u9_u4_n180 ) );
  NAND2_X1 u0_u9_u4_U53 (.A2( u0_u9_u4_n104 ) , .A1( u0_u9_u4_n105 ) , .ZN( u0_u9_u4_n146 ) );
  NAND2_X1 u0_u9_u4_U54 (.A2( u0_u9_u4_n101 ) , .A1( u0_u9_u4_n102 ) , .ZN( u0_u9_u4_n160 ) );
  NAND2_X1 u0_u9_u4_U55 (.ZN( u0_u9_u4_n134 ) , .A1( u0_u9_u4_n98 ) , .A2( u0_u9_u4_n99 ) );
  NAND2_X1 u0_u9_u4_U56 (.A1( u0_u9_u4_n103 ) , .A2( u0_u9_u4_n104 ) , .ZN( u0_u9_u4_n143 ) );
  NAND2_X1 u0_u9_u4_U57 (.A2( u0_u9_u4_n105 ) , .ZN( u0_u9_u4_n145 ) , .A1( u0_u9_u4_n98 ) );
  NAND2_X1 u0_u9_u4_U58 (.A1( u0_u9_u4_n100 ) , .A2( u0_u9_u4_n105 ) , .ZN( u0_u9_u4_n120 ) );
  NAND2_X1 u0_u9_u4_U59 (.A1( u0_u9_u4_n102 ) , .A2( u0_u9_u4_n104 ) , .ZN( u0_u9_u4_n148 ) );
  AOI21_X1 u0_u9_u4_U6 (.ZN( u0_u9_u4_n106 ) , .B2( u0_u9_u4_n146 ) , .B1( u0_u9_u4_n158 ) , .A( u0_u9_u4_n170 ) );
  NAND2_X1 u0_u9_u4_U60 (.A2( u0_u9_u4_n100 ) , .A1( u0_u9_u4_n103 ) , .ZN( u0_u9_u4_n157 ) );
  INV_X1 u0_u9_u4_U61 (.A( u0_u9_u4_n150 ) , .ZN( u0_u9_u4_n173 ) );
  INV_X1 u0_u9_u4_U62 (.A( u0_u9_u4_n152 ) , .ZN( u0_u9_u4_n171 ) );
  NAND2_X1 u0_u9_u4_U63 (.A1( u0_u9_u4_n100 ) , .ZN( u0_u9_u4_n118 ) , .A2( u0_u9_u4_n99 ) );
  NAND2_X1 u0_u9_u4_U64 (.A2( u0_u9_u4_n100 ) , .A1( u0_u9_u4_n102 ) , .ZN( u0_u9_u4_n144 ) );
  NAND2_X1 u0_u9_u4_U65 (.A2( u0_u9_u4_n101 ) , .A1( u0_u9_u4_n105 ) , .ZN( u0_u9_u4_n96 ) );
  INV_X1 u0_u9_u4_U66 (.A( u0_u9_u4_n128 ) , .ZN( u0_u9_u4_n174 ) );
  NAND2_X1 u0_u9_u4_U67 (.A2( u0_u9_u4_n102 ) , .ZN( u0_u9_u4_n119 ) , .A1( u0_u9_u4_n98 ) );
  NAND2_X1 u0_u9_u4_U68 (.A2( u0_u9_u4_n101 ) , .A1( u0_u9_u4_n103 ) , .ZN( u0_u9_u4_n147 ) );
  NAND2_X1 u0_u9_u4_U69 (.A2( u0_u9_u4_n104 ) , .ZN( u0_u9_u4_n113 ) , .A1( u0_u9_u4_n99 ) );
  AOI21_X1 u0_u9_u4_U7 (.ZN( u0_u9_u4_n108 ) , .B2( u0_u9_u4_n134 ) , .B1( u0_u9_u4_n155 ) , .A( u0_u9_u4_n156 ) );
  NOR2_X1 u0_u9_u4_U70 (.A2( u0_u9_X_28 ) , .ZN( u0_u9_u4_n150 ) , .A1( u0_u9_u4_n168 ) );
  NOR2_X1 u0_u9_u4_U71 (.A2( u0_u9_X_29 ) , .ZN( u0_u9_u4_n152 ) , .A1( u0_u9_u4_n169 ) );
  NOR2_X1 u0_u9_u4_U72 (.A2( u0_u9_X_30 ) , .ZN( u0_u9_u4_n105 ) , .A1( u0_u9_u4_n176 ) );
  NOR2_X1 u0_u9_u4_U73 (.A2( u0_u9_X_26 ) , .ZN( u0_u9_u4_n100 ) , .A1( u0_u9_u4_n177 ) );
  NOR2_X1 u0_u9_u4_U74 (.A2( u0_u9_X_28 ) , .A1( u0_u9_X_29 ) , .ZN( u0_u9_u4_n128 ) );
  NOR2_X1 u0_u9_u4_U75 (.A2( u0_u9_X_27 ) , .A1( u0_u9_X_30 ) , .ZN( u0_u9_u4_n102 ) );
  NOR2_X1 u0_u9_u4_U76 (.A2( u0_u9_X_25 ) , .A1( u0_u9_X_26 ) , .ZN( u0_u9_u4_n98 ) );
  AND2_X1 u0_u9_u4_U77 (.A2( u0_u9_X_25 ) , .A1( u0_u9_X_26 ) , .ZN( u0_u9_u4_n104 ) );
  AND2_X1 u0_u9_u4_U78 (.A1( u0_u9_X_30 ) , .A2( u0_u9_u4_n176 ) , .ZN( u0_u9_u4_n99 ) );
  AND2_X1 u0_u9_u4_U79 (.A1( u0_u9_X_26 ) , .ZN( u0_u9_u4_n101 ) , .A2( u0_u9_u4_n177 ) );
  AOI21_X1 u0_u9_u4_U8 (.ZN( u0_u9_u4_n109 ) , .A( u0_u9_u4_n153 ) , .B1( u0_u9_u4_n159 ) , .B2( u0_u9_u4_n184 ) );
  AND2_X1 u0_u9_u4_U80 (.A1( u0_u9_X_27 ) , .A2( u0_u9_X_30 ) , .ZN( u0_u9_u4_n103 ) );
  INV_X1 u0_u9_u4_U81 (.A( u0_u9_X_28 ) , .ZN( u0_u9_u4_n169 ) );
  INV_X1 u0_u9_u4_U82 (.A( u0_u9_X_29 ) , .ZN( u0_u9_u4_n168 ) );
  INV_X1 u0_u9_u4_U83 (.A( u0_u9_X_25 ) , .ZN( u0_u9_u4_n177 ) );
  INV_X1 u0_u9_u4_U84 (.A( u0_u9_X_27 ) , .ZN( u0_u9_u4_n176 ) );
  NAND4_X1 u0_u9_u4_U85 (.ZN( u0_out9_25 ) , .A4( u0_u9_u4_n139 ) , .A3( u0_u9_u4_n140 ) , .A2( u0_u9_u4_n141 ) , .A1( u0_u9_u4_n142 ) );
  OAI21_X1 u0_u9_u4_U86 (.A( u0_u9_u4_n128 ) , .B2( u0_u9_u4_n129 ) , .B1( u0_u9_u4_n130 ) , .ZN( u0_u9_u4_n142 ) );
  OAI21_X1 u0_u9_u4_U87 (.B2( u0_u9_u4_n131 ) , .ZN( u0_u9_u4_n141 ) , .A( u0_u9_u4_n175 ) , .B1( u0_u9_u4_n183 ) );
  NAND4_X1 u0_u9_u4_U88 (.ZN( u0_out9_14 ) , .A4( u0_u9_u4_n124 ) , .A3( u0_u9_u4_n125 ) , .A2( u0_u9_u4_n126 ) , .A1( u0_u9_u4_n127 ) );
  AOI22_X1 u0_u9_u4_U89 (.B2( u0_u9_u4_n117 ) , .ZN( u0_u9_u4_n126 ) , .A1( u0_u9_u4_n129 ) , .B1( u0_u9_u4_n152 ) , .A2( u0_u9_u4_n175 ) );
  AOI211_X1 u0_u9_u4_U9 (.B( u0_u9_u4_n136 ) , .A( u0_u9_u4_n137 ) , .C2( u0_u9_u4_n138 ) , .ZN( u0_u9_u4_n139 ) , .C1( u0_u9_u4_n182 ) );
  AOI22_X1 u0_u9_u4_U90 (.ZN( u0_u9_u4_n125 ) , .B2( u0_u9_u4_n131 ) , .A2( u0_u9_u4_n132 ) , .B1( u0_u9_u4_n138 ) , .A1( u0_u9_u4_n178 ) );
  NAND4_X1 u0_u9_u4_U91 (.ZN( u0_out9_8 ) , .A4( u0_u9_u4_n110 ) , .A3( u0_u9_u4_n111 ) , .A2( u0_u9_u4_n112 ) , .A1( u0_u9_u4_n186 ) );
  NAND2_X1 u0_u9_u4_U92 (.ZN( u0_u9_u4_n112 ) , .A2( u0_u9_u4_n130 ) , .A1( u0_u9_u4_n150 ) );
  AOI22_X1 u0_u9_u4_U93 (.ZN( u0_u9_u4_n111 ) , .B2( u0_u9_u4_n132 ) , .A1( u0_u9_u4_n152 ) , .B1( u0_u9_u4_n178 ) , .A2( u0_u9_u4_n97 ) );
  AOI22_X1 u0_u9_u4_U94 (.B2( u0_u9_u4_n149 ) , .B1( u0_u9_u4_n150 ) , .A2( u0_u9_u4_n151 ) , .A1( u0_u9_u4_n152 ) , .ZN( u0_u9_u4_n167 ) );
  NOR4_X1 u0_u9_u4_U95 (.A4( u0_u9_u4_n162 ) , .A3( u0_u9_u4_n163 ) , .A2( u0_u9_u4_n164 ) , .A1( u0_u9_u4_n165 ) , .ZN( u0_u9_u4_n166 ) );
  NAND3_X1 u0_u9_u4_U96 (.ZN( u0_out9_3 ) , .A3( u0_u9_u4_n166 ) , .A1( u0_u9_u4_n167 ) , .A2( u0_u9_u4_n186 ) );
  NAND3_X1 u0_u9_u4_U97 (.A3( u0_u9_u4_n146 ) , .A2( u0_u9_u4_n147 ) , .A1( u0_u9_u4_n148 ) , .ZN( u0_u9_u4_n149 ) );
  NAND3_X1 u0_u9_u4_U98 (.A3( u0_u9_u4_n143 ) , .A2( u0_u9_u4_n144 ) , .A1( u0_u9_u4_n145 ) , .ZN( u0_u9_u4_n151 ) );
  NAND3_X1 u0_u9_u4_U99 (.A3( u0_u9_u4_n121 ) , .ZN( u0_u9_u4_n122 ) , .A2( u0_u9_u4_n144 ) , .A1( u0_u9_u4_n154 ) );
  NOR2_X1 u0_u9_u5_U10 (.ZN( u0_u9_u5_n135 ) , .A1( u0_u9_u5_n173 ) , .A2( u0_u9_u5_n176 ) );
  NOR3_X1 u0_u9_u5_U100 (.A3( u0_u9_u5_n141 ) , .A1( u0_u9_u5_n142 ) , .ZN( u0_u9_u5_n143 ) , .A2( u0_u9_u5_n191 ) );
  NAND4_X1 u0_u9_u5_U101 (.ZN( u0_out9_4 ) , .A4( u0_u9_u5_n112 ) , .A2( u0_u9_u5_n113 ) , .A1( u0_u9_u5_n114 ) , .A3( u0_u9_u5_n195 ) );
  AOI211_X1 u0_u9_u5_U102 (.A( u0_u9_u5_n110 ) , .C1( u0_u9_u5_n111 ) , .ZN( u0_u9_u5_n112 ) , .B( u0_u9_u5_n118 ) , .C2( u0_u9_u5_n177 ) );
  INV_X1 u0_u9_u5_U103 (.A( u0_u9_u5_n102 ) , .ZN( u0_u9_u5_n195 ) );
  NAND3_X1 u0_u9_u5_U104 (.A2( u0_u9_u5_n154 ) , .A3( u0_u9_u5_n158 ) , .A1( u0_u9_u5_n161 ) , .ZN( u0_u9_u5_n99 ) );
  INV_X1 u0_u9_u5_U11 (.A( u0_u9_u5_n121 ) , .ZN( u0_u9_u5_n177 ) );
  NOR2_X1 u0_u9_u5_U12 (.ZN( u0_u9_u5_n160 ) , .A2( u0_u9_u5_n173 ) , .A1( u0_u9_u5_n177 ) );
  INV_X1 u0_u9_u5_U13 (.A( u0_u9_u5_n150 ) , .ZN( u0_u9_u5_n174 ) );
  AOI21_X1 u0_u9_u5_U14 (.A( u0_u9_u5_n160 ) , .B2( u0_u9_u5_n161 ) , .ZN( u0_u9_u5_n162 ) , .B1( u0_u9_u5_n192 ) );
  INV_X1 u0_u9_u5_U15 (.A( u0_u9_u5_n159 ) , .ZN( u0_u9_u5_n192 ) );
  AOI21_X1 u0_u9_u5_U16 (.A( u0_u9_u5_n156 ) , .B2( u0_u9_u5_n157 ) , .B1( u0_u9_u5_n158 ) , .ZN( u0_u9_u5_n163 ) );
  AOI21_X1 u0_u9_u5_U17 (.B2( u0_u9_u5_n139 ) , .B1( u0_u9_u5_n140 ) , .ZN( u0_u9_u5_n141 ) , .A( u0_u9_u5_n150 ) );
  OAI21_X1 u0_u9_u5_U18 (.A( u0_u9_u5_n133 ) , .B2( u0_u9_u5_n134 ) , .B1( u0_u9_u5_n135 ) , .ZN( u0_u9_u5_n142 ) );
  OAI21_X1 u0_u9_u5_U19 (.ZN( u0_u9_u5_n133 ) , .B2( u0_u9_u5_n147 ) , .A( u0_u9_u5_n173 ) , .B1( u0_u9_u5_n188 ) );
  NAND2_X1 u0_u9_u5_U20 (.A2( u0_u9_u5_n119 ) , .A1( u0_u9_u5_n123 ) , .ZN( u0_u9_u5_n137 ) );
  INV_X1 u0_u9_u5_U21 (.A( u0_u9_u5_n155 ) , .ZN( u0_u9_u5_n194 ) );
  NAND2_X1 u0_u9_u5_U22 (.A1( u0_u9_u5_n121 ) , .ZN( u0_u9_u5_n132 ) , .A2( u0_u9_u5_n172 ) );
  NAND2_X1 u0_u9_u5_U23 (.A2( u0_u9_u5_n122 ) , .ZN( u0_u9_u5_n136 ) , .A1( u0_u9_u5_n154 ) );
  NAND2_X1 u0_u9_u5_U24 (.A2( u0_u9_u5_n119 ) , .A1( u0_u9_u5_n120 ) , .ZN( u0_u9_u5_n159 ) );
  INV_X1 u0_u9_u5_U25 (.A( u0_u9_u5_n156 ) , .ZN( u0_u9_u5_n175 ) );
  INV_X1 u0_u9_u5_U26 (.A( u0_u9_u5_n158 ) , .ZN( u0_u9_u5_n188 ) );
  INV_X1 u0_u9_u5_U27 (.A( u0_u9_u5_n152 ) , .ZN( u0_u9_u5_n179 ) );
  INV_X1 u0_u9_u5_U28 (.A( u0_u9_u5_n140 ) , .ZN( u0_u9_u5_n182 ) );
  INV_X1 u0_u9_u5_U29 (.A( u0_u9_u5_n151 ) , .ZN( u0_u9_u5_n183 ) );
  NOR2_X1 u0_u9_u5_U3 (.ZN( u0_u9_u5_n134 ) , .A1( u0_u9_u5_n183 ) , .A2( u0_u9_u5_n190 ) );
  INV_X1 u0_u9_u5_U30 (.A( u0_u9_u5_n123 ) , .ZN( u0_u9_u5_n185 ) );
  INV_X1 u0_u9_u5_U31 (.A( u0_u9_u5_n161 ) , .ZN( u0_u9_u5_n184 ) );
  INV_X1 u0_u9_u5_U32 (.A( u0_u9_u5_n139 ) , .ZN( u0_u9_u5_n189 ) );
  INV_X1 u0_u9_u5_U33 (.A( u0_u9_u5_n157 ) , .ZN( u0_u9_u5_n190 ) );
  INV_X1 u0_u9_u5_U34 (.A( u0_u9_u5_n120 ) , .ZN( u0_u9_u5_n193 ) );
  NAND2_X1 u0_u9_u5_U35 (.ZN( u0_u9_u5_n111 ) , .A1( u0_u9_u5_n140 ) , .A2( u0_u9_u5_n155 ) );
  NOR2_X1 u0_u9_u5_U36 (.ZN( u0_u9_u5_n100 ) , .A1( u0_u9_u5_n170 ) , .A2( u0_u9_u5_n180 ) );
  INV_X1 u0_u9_u5_U37 (.A( u0_u9_u5_n117 ) , .ZN( u0_u9_u5_n196 ) );
  OAI221_X1 u0_u9_u5_U38 (.A( u0_u9_u5_n116 ) , .ZN( u0_u9_u5_n117 ) , .B2( u0_u9_u5_n119 ) , .C1( u0_u9_u5_n153 ) , .C2( u0_u9_u5_n158 ) , .B1( u0_u9_u5_n172 ) );
  AOI222_X1 u0_u9_u5_U39 (.ZN( u0_u9_u5_n116 ) , .B2( u0_u9_u5_n145 ) , .C1( u0_u9_u5_n148 ) , .A2( u0_u9_u5_n174 ) , .C2( u0_u9_u5_n177 ) , .B1( u0_u9_u5_n187 ) , .A1( u0_u9_u5_n193 ) );
  INV_X1 u0_u9_u5_U4 (.A( u0_u9_u5_n138 ) , .ZN( u0_u9_u5_n191 ) );
  INV_X1 u0_u9_u5_U40 (.A( u0_u9_u5_n115 ) , .ZN( u0_u9_u5_n187 ) );
  OAI221_X1 u0_u9_u5_U41 (.A( u0_u9_u5_n101 ) , .ZN( u0_u9_u5_n102 ) , .C2( u0_u9_u5_n115 ) , .C1( u0_u9_u5_n126 ) , .B1( u0_u9_u5_n134 ) , .B2( u0_u9_u5_n160 ) );
  OAI21_X1 u0_u9_u5_U42 (.ZN( u0_u9_u5_n101 ) , .B1( u0_u9_u5_n137 ) , .A( u0_u9_u5_n146 ) , .B2( u0_u9_u5_n147 ) );
  AOI22_X1 u0_u9_u5_U43 (.B2( u0_u9_u5_n131 ) , .A2( u0_u9_u5_n146 ) , .ZN( u0_u9_u5_n169 ) , .B1( u0_u9_u5_n174 ) , .A1( u0_u9_u5_n185 ) );
  NOR2_X1 u0_u9_u5_U44 (.A1( u0_u9_u5_n146 ) , .ZN( u0_u9_u5_n150 ) , .A2( u0_u9_u5_n173 ) );
  AOI21_X1 u0_u9_u5_U45 (.A( u0_u9_u5_n118 ) , .B2( u0_u9_u5_n145 ) , .ZN( u0_u9_u5_n168 ) , .B1( u0_u9_u5_n186 ) );
  INV_X1 u0_u9_u5_U46 (.A( u0_u9_u5_n122 ) , .ZN( u0_u9_u5_n186 ) );
  NOR2_X1 u0_u9_u5_U47 (.A1( u0_u9_u5_n146 ) , .ZN( u0_u9_u5_n152 ) , .A2( u0_u9_u5_n176 ) );
  NOR2_X1 u0_u9_u5_U48 (.A1( u0_u9_u5_n115 ) , .ZN( u0_u9_u5_n118 ) , .A2( u0_u9_u5_n153 ) );
  NOR2_X1 u0_u9_u5_U49 (.A2( u0_u9_u5_n145 ) , .ZN( u0_u9_u5_n156 ) , .A1( u0_u9_u5_n174 ) );
  OAI21_X1 u0_u9_u5_U5 (.B2( u0_u9_u5_n136 ) , .B1( u0_u9_u5_n137 ) , .ZN( u0_u9_u5_n138 ) , .A( u0_u9_u5_n177 ) );
  NOR2_X1 u0_u9_u5_U50 (.ZN( u0_u9_u5_n121 ) , .A2( u0_u9_u5_n145 ) , .A1( u0_u9_u5_n176 ) );
  AOI22_X1 u0_u9_u5_U51 (.ZN( u0_u9_u5_n114 ) , .A2( u0_u9_u5_n137 ) , .A1( u0_u9_u5_n145 ) , .B2( u0_u9_u5_n175 ) , .B1( u0_u9_u5_n193 ) );
  OAI211_X1 u0_u9_u5_U52 (.B( u0_u9_u5_n124 ) , .A( u0_u9_u5_n125 ) , .C2( u0_u9_u5_n126 ) , .C1( u0_u9_u5_n127 ) , .ZN( u0_u9_u5_n128 ) );
  NOR3_X1 u0_u9_u5_U53 (.ZN( u0_u9_u5_n127 ) , .A1( u0_u9_u5_n136 ) , .A3( u0_u9_u5_n148 ) , .A2( u0_u9_u5_n182 ) );
  OAI21_X1 u0_u9_u5_U54 (.ZN( u0_u9_u5_n124 ) , .A( u0_u9_u5_n177 ) , .B2( u0_u9_u5_n183 ) , .B1( u0_u9_u5_n189 ) );
  OAI21_X1 u0_u9_u5_U55 (.ZN( u0_u9_u5_n125 ) , .A( u0_u9_u5_n174 ) , .B2( u0_u9_u5_n185 ) , .B1( u0_u9_u5_n190 ) );
  AOI21_X1 u0_u9_u5_U56 (.A( u0_u9_u5_n153 ) , .B2( u0_u9_u5_n154 ) , .B1( u0_u9_u5_n155 ) , .ZN( u0_u9_u5_n164 ) );
  AOI21_X1 u0_u9_u5_U57 (.ZN( u0_u9_u5_n110 ) , .B1( u0_u9_u5_n122 ) , .B2( u0_u9_u5_n139 ) , .A( u0_u9_u5_n153 ) );
  INV_X1 u0_u9_u5_U58 (.A( u0_u9_u5_n153 ) , .ZN( u0_u9_u5_n176 ) );
  INV_X1 u0_u9_u5_U59 (.A( u0_u9_u5_n126 ) , .ZN( u0_u9_u5_n173 ) );
  AOI222_X1 u0_u9_u5_U6 (.ZN( u0_u9_u5_n113 ) , .A1( u0_u9_u5_n131 ) , .C1( u0_u9_u5_n148 ) , .B2( u0_u9_u5_n174 ) , .C2( u0_u9_u5_n178 ) , .A2( u0_u9_u5_n179 ) , .B1( u0_u9_u5_n99 ) );
  AND2_X1 u0_u9_u5_U60 (.A2( u0_u9_u5_n104 ) , .A1( u0_u9_u5_n107 ) , .ZN( u0_u9_u5_n147 ) );
  AND2_X1 u0_u9_u5_U61 (.A2( u0_u9_u5_n104 ) , .A1( u0_u9_u5_n108 ) , .ZN( u0_u9_u5_n148 ) );
  NAND2_X1 u0_u9_u5_U62 (.A1( u0_u9_u5_n105 ) , .A2( u0_u9_u5_n106 ) , .ZN( u0_u9_u5_n158 ) );
  NAND2_X1 u0_u9_u5_U63 (.A2( u0_u9_u5_n108 ) , .A1( u0_u9_u5_n109 ) , .ZN( u0_u9_u5_n139 ) );
  NAND2_X1 u0_u9_u5_U64 (.A1( u0_u9_u5_n106 ) , .A2( u0_u9_u5_n108 ) , .ZN( u0_u9_u5_n119 ) );
  NAND2_X1 u0_u9_u5_U65 (.A2( u0_u9_u5_n103 ) , .A1( u0_u9_u5_n105 ) , .ZN( u0_u9_u5_n140 ) );
  NAND2_X1 u0_u9_u5_U66 (.A2( u0_u9_u5_n104 ) , .A1( u0_u9_u5_n105 ) , .ZN( u0_u9_u5_n155 ) );
  NAND2_X1 u0_u9_u5_U67 (.A2( u0_u9_u5_n106 ) , .A1( u0_u9_u5_n107 ) , .ZN( u0_u9_u5_n122 ) );
  NAND2_X1 u0_u9_u5_U68 (.A2( u0_u9_u5_n100 ) , .A1( u0_u9_u5_n106 ) , .ZN( u0_u9_u5_n115 ) );
  NAND2_X1 u0_u9_u5_U69 (.A2( u0_u9_u5_n100 ) , .A1( u0_u9_u5_n103 ) , .ZN( u0_u9_u5_n161 ) );
  INV_X1 u0_u9_u5_U7 (.A( u0_u9_u5_n135 ) , .ZN( u0_u9_u5_n178 ) );
  NAND2_X1 u0_u9_u5_U70 (.A1( u0_u9_u5_n105 ) , .A2( u0_u9_u5_n109 ) , .ZN( u0_u9_u5_n154 ) );
  INV_X1 u0_u9_u5_U71 (.A( u0_u9_u5_n146 ) , .ZN( u0_u9_u5_n172 ) );
  NAND2_X1 u0_u9_u5_U72 (.A1( u0_u9_u5_n103 ) , .A2( u0_u9_u5_n108 ) , .ZN( u0_u9_u5_n123 ) );
  NAND2_X1 u0_u9_u5_U73 (.A2( u0_u9_u5_n103 ) , .A1( u0_u9_u5_n107 ) , .ZN( u0_u9_u5_n151 ) );
  NAND2_X1 u0_u9_u5_U74 (.A2( u0_u9_u5_n107 ) , .A1( u0_u9_u5_n109 ) , .ZN( u0_u9_u5_n120 ) );
  NAND2_X1 u0_u9_u5_U75 (.A2( u0_u9_u5_n100 ) , .A1( u0_u9_u5_n109 ) , .ZN( u0_u9_u5_n157 ) );
  AND2_X1 u0_u9_u5_U76 (.A2( u0_u9_u5_n100 ) , .A1( u0_u9_u5_n104 ) , .ZN( u0_u9_u5_n131 ) );
  NOR2_X1 u0_u9_u5_U77 (.A2( u0_u9_X_34 ) , .A1( u0_u9_X_35 ) , .ZN( u0_u9_u5_n145 ) );
  NOR2_X1 u0_u9_u5_U78 (.A2( u0_u9_X_34 ) , .ZN( u0_u9_u5_n146 ) , .A1( u0_u9_u5_n171 ) );
  NOR2_X1 u0_u9_u5_U79 (.A2( u0_u9_X_31 ) , .A1( u0_u9_X_32 ) , .ZN( u0_u9_u5_n103 ) );
  OAI22_X1 u0_u9_u5_U8 (.B2( u0_u9_u5_n149 ) , .B1( u0_u9_u5_n150 ) , .A2( u0_u9_u5_n151 ) , .A1( u0_u9_u5_n152 ) , .ZN( u0_u9_u5_n165 ) );
  NOR2_X1 u0_u9_u5_U80 (.A2( u0_u9_X_36 ) , .ZN( u0_u9_u5_n105 ) , .A1( u0_u9_u5_n180 ) );
  NOR2_X1 u0_u9_u5_U81 (.A2( u0_u9_X_33 ) , .ZN( u0_u9_u5_n108 ) , .A1( u0_u9_u5_n170 ) );
  NOR2_X1 u0_u9_u5_U82 (.A2( u0_u9_X_33 ) , .A1( u0_u9_X_36 ) , .ZN( u0_u9_u5_n107 ) );
  NOR2_X1 u0_u9_u5_U83 (.A2( u0_u9_X_31 ) , .ZN( u0_u9_u5_n104 ) , .A1( u0_u9_u5_n181 ) );
  NAND2_X1 u0_u9_u5_U84 (.A2( u0_u9_X_34 ) , .A1( u0_u9_X_35 ) , .ZN( u0_u9_u5_n153 ) );
  NAND2_X1 u0_u9_u5_U85 (.A1( u0_u9_X_34 ) , .ZN( u0_u9_u5_n126 ) , .A2( u0_u9_u5_n171 ) );
  AND2_X1 u0_u9_u5_U86 (.A1( u0_u9_X_31 ) , .A2( u0_u9_X_32 ) , .ZN( u0_u9_u5_n106 ) );
  AND2_X1 u0_u9_u5_U87 (.A1( u0_u9_X_31 ) , .ZN( u0_u9_u5_n109 ) , .A2( u0_u9_u5_n181 ) );
  INV_X1 u0_u9_u5_U88 (.A( u0_u9_X_33 ) , .ZN( u0_u9_u5_n180 ) );
  INV_X1 u0_u9_u5_U89 (.A( u0_u9_X_35 ) , .ZN( u0_u9_u5_n171 ) );
  NOR3_X1 u0_u9_u5_U9 (.A2( u0_u9_u5_n147 ) , .A1( u0_u9_u5_n148 ) , .ZN( u0_u9_u5_n149 ) , .A3( u0_u9_u5_n194 ) );
  INV_X1 u0_u9_u5_U90 (.A( u0_u9_X_36 ) , .ZN( u0_u9_u5_n170 ) );
  INV_X1 u0_u9_u5_U91 (.A( u0_u9_X_32 ) , .ZN( u0_u9_u5_n181 ) );
  NAND4_X1 u0_u9_u5_U92 (.ZN( u0_out9_29 ) , .A4( u0_u9_u5_n129 ) , .A3( u0_u9_u5_n130 ) , .A2( u0_u9_u5_n168 ) , .A1( u0_u9_u5_n196 ) );
  AOI221_X1 u0_u9_u5_U93 (.A( u0_u9_u5_n128 ) , .ZN( u0_u9_u5_n129 ) , .C2( u0_u9_u5_n132 ) , .B2( u0_u9_u5_n159 ) , .B1( u0_u9_u5_n176 ) , .C1( u0_u9_u5_n184 ) );
  AOI222_X1 u0_u9_u5_U94 (.ZN( u0_u9_u5_n130 ) , .A2( u0_u9_u5_n146 ) , .B1( u0_u9_u5_n147 ) , .C2( u0_u9_u5_n175 ) , .B2( u0_u9_u5_n179 ) , .A1( u0_u9_u5_n188 ) , .C1( u0_u9_u5_n194 ) );
  NAND4_X1 u0_u9_u5_U95 (.ZN( u0_out9_19 ) , .A4( u0_u9_u5_n166 ) , .A3( u0_u9_u5_n167 ) , .A2( u0_u9_u5_n168 ) , .A1( u0_u9_u5_n169 ) );
  AOI22_X1 u0_u9_u5_U96 (.B2( u0_u9_u5_n145 ) , .A2( u0_u9_u5_n146 ) , .ZN( u0_u9_u5_n167 ) , .B1( u0_u9_u5_n182 ) , .A1( u0_u9_u5_n189 ) );
  NOR4_X1 u0_u9_u5_U97 (.A4( u0_u9_u5_n162 ) , .A3( u0_u9_u5_n163 ) , .A2( u0_u9_u5_n164 ) , .A1( u0_u9_u5_n165 ) , .ZN( u0_u9_u5_n166 ) );
  NAND4_X1 u0_u9_u5_U98 (.ZN( u0_out9_11 ) , .A4( u0_u9_u5_n143 ) , .A3( u0_u9_u5_n144 ) , .A2( u0_u9_u5_n169 ) , .A1( u0_u9_u5_n196 ) );
  AOI22_X1 u0_u9_u5_U99 (.A2( u0_u9_u5_n132 ) , .ZN( u0_u9_u5_n144 ) , .B2( u0_u9_u5_n145 ) , .B1( u0_u9_u5_n184 ) , .A1( u0_u9_u5_n194 ) );
  AOI22_X1 u0_u9_u6_U10 (.A2( u0_u9_u6_n151 ) , .B2( u0_u9_u6_n161 ) , .A1( u0_u9_u6_n167 ) , .B1( u0_u9_u6_n170 ) , .ZN( u0_u9_u6_n89 ) );
  AOI21_X1 u0_u9_u6_U11 (.B1( u0_u9_u6_n107 ) , .B2( u0_u9_u6_n132 ) , .A( u0_u9_u6_n158 ) , .ZN( u0_u9_u6_n88 ) );
  AOI21_X1 u0_u9_u6_U12 (.B2( u0_u9_u6_n147 ) , .B1( u0_u9_u6_n148 ) , .ZN( u0_u9_u6_n149 ) , .A( u0_u9_u6_n158 ) );
  AOI21_X1 u0_u9_u6_U13 (.ZN( u0_u9_u6_n106 ) , .A( u0_u9_u6_n142 ) , .B2( u0_u9_u6_n159 ) , .B1( u0_u9_u6_n164 ) );
  INV_X1 u0_u9_u6_U14 (.A( u0_u9_u6_n155 ) , .ZN( u0_u9_u6_n161 ) );
  INV_X1 u0_u9_u6_U15 (.A( u0_u9_u6_n128 ) , .ZN( u0_u9_u6_n164 ) );
  NAND2_X1 u0_u9_u6_U16 (.ZN( u0_u9_u6_n110 ) , .A1( u0_u9_u6_n122 ) , .A2( u0_u9_u6_n129 ) );
  NAND2_X1 u0_u9_u6_U17 (.ZN( u0_u9_u6_n124 ) , .A2( u0_u9_u6_n146 ) , .A1( u0_u9_u6_n148 ) );
  INV_X1 u0_u9_u6_U18 (.A( u0_u9_u6_n132 ) , .ZN( u0_u9_u6_n171 ) );
  AND2_X1 u0_u9_u6_U19 (.A1( u0_u9_u6_n100 ) , .ZN( u0_u9_u6_n130 ) , .A2( u0_u9_u6_n147 ) );
  INV_X1 u0_u9_u6_U20 (.A( u0_u9_u6_n127 ) , .ZN( u0_u9_u6_n173 ) );
  INV_X1 u0_u9_u6_U21 (.A( u0_u9_u6_n121 ) , .ZN( u0_u9_u6_n167 ) );
  INV_X1 u0_u9_u6_U22 (.A( u0_u9_u6_n100 ) , .ZN( u0_u9_u6_n169 ) );
  INV_X1 u0_u9_u6_U23 (.A( u0_u9_u6_n123 ) , .ZN( u0_u9_u6_n170 ) );
  INV_X1 u0_u9_u6_U24 (.A( u0_u9_u6_n113 ) , .ZN( u0_u9_u6_n168 ) );
  AND2_X1 u0_u9_u6_U25 (.A1( u0_u9_u6_n107 ) , .A2( u0_u9_u6_n119 ) , .ZN( u0_u9_u6_n133 ) );
  AND2_X1 u0_u9_u6_U26 (.A2( u0_u9_u6_n121 ) , .A1( u0_u9_u6_n122 ) , .ZN( u0_u9_u6_n131 ) );
  AND3_X1 u0_u9_u6_U27 (.ZN( u0_u9_u6_n120 ) , .A2( u0_u9_u6_n127 ) , .A1( u0_u9_u6_n132 ) , .A3( u0_u9_u6_n145 ) );
  INV_X1 u0_u9_u6_U28 (.A( u0_u9_u6_n146 ) , .ZN( u0_u9_u6_n163 ) );
  AOI222_X1 u0_u9_u6_U29 (.ZN( u0_u9_u6_n114 ) , .A1( u0_u9_u6_n118 ) , .A2( u0_u9_u6_n126 ) , .B2( u0_u9_u6_n151 ) , .C2( u0_u9_u6_n159 ) , .C1( u0_u9_u6_n168 ) , .B1( u0_u9_u6_n169 ) );
  INV_X1 u0_u9_u6_U3 (.A( u0_u9_u6_n110 ) , .ZN( u0_u9_u6_n166 ) );
  NOR2_X1 u0_u9_u6_U30 (.A1( u0_u9_u6_n162 ) , .A2( u0_u9_u6_n165 ) , .ZN( u0_u9_u6_n98 ) );
  NAND2_X1 u0_u9_u6_U31 (.A1( u0_u9_u6_n144 ) , .ZN( u0_u9_u6_n151 ) , .A2( u0_u9_u6_n158 ) );
  NAND2_X1 u0_u9_u6_U32 (.ZN( u0_u9_u6_n132 ) , .A1( u0_u9_u6_n91 ) , .A2( u0_u9_u6_n97 ) );
  AOI22_X1 u0_u9_u6_U33 (.B2( u0_u9_u6_n110 ) , .B1( u0_u9_u6_n111 ) , .A1( u0_u9_u6_n112 ) , .ZN( u0_u9_u6_n115 ) , .A2( u0_u9_u6_n161 ) );
  NAND4_X1 u0_u9_u6_U34 (.A3( u0_u9_u6_n109 ) , .ZN( u0_u9_u6_n112 ) , .A4( u0_u9_u6_n132 ) , .A2( u0_u9_u6_n147 ) , .A1( u0_u9_u6_n166 ) );
  NOR2_X1 u0_u9_u6_U35 (.ZN( u0_u9_u6_n109 ) , .A1( u0_u9_u6_n170 ) , .A2( u0_u9_u6_n173 ) );
  NOR2_X1 u0_u9_u6_U36 (.A2( u0_u9_u6_n126 ) , .ZN( u0_u9_u6_n155 ) , .A1( u0_u9_u6_n160 ) );
  NAND2_X1 u0_u9_u6_U37 (.ZN( u0_u9_u6_n146 ) , .A2( u0_u9_u6_n94 ) , .A1( u0_u9_u6_n99 ) );
  AOI21_X1 u0_u9_u6_U38 (.A( u0_u9_u6_n144 ) , .B2( u0_u9_u6_n145 ) , .B1( u0_u9_u6_n146 ) , .ZN( u0_u9_u6_n150 ) );
  AOI211_X1 u0_u9_u6_U39 (.B( u0_u9_u6_n134 ) , .A( u0_u9_u6_n135 ) , .C1( u0_u9_u6_n136 ) , .ZN( u0_u9_u6_n137 ) , .C2( u0_u9_u6_n151 ) );
  INV_X1 u0_u9_u6_U4 (.A( u0_u9_u6_n142 ) , .ZN( u0_u9_u6_n174 ) );
  NAND4_X1 u0_u9_u6_U40 (.A4( u0_u9_u6_n127 ) , .A3( u0_u9_u6_n128 ) , .A2( u0_u9_u6_n129 ) , .A1( u0_u9_u6_n130 ) , .ZN( u0_u9_u6_n136 ) );
  AOI21_X1 u0_u9_u6_U41 (.B2( u0_u9_u6_n132 ) , .B1( u0_u9_u6_n133 ) , .ZN( u0_u9_u6_n134 ) , .A( u0_u9_u6_n158 ) );
  AOI21_X1 u0_u9_u6_U42 (.B1( u0_u9_u6_n131 ) , .ZN( u0_u9_u6_n135 ) , .A( u0_u9_u6_n144 ) , .B2( u0_u9_u6_n146 ) );
  INV_X1 u0_u9_u6_U43 (.A( u0_u9_u6_n111 ) , .ZN( u0_u9_u6_n158 ) );
  NAND2_X1 u0_u9_u6_U44 (.ZN( u0_u9_u6_n127 ) , .A1( u0_u9_u6_n91 ) , .A2( u0_u9_u6_n92 ) );
  NAND2_X1 u0_u9_u6_U45 (.ZN( u0_u9_u6_n129 ) , .A2( u0_u9_u6_n95 ) , .A1( u0_u9_u6_n96 ) );
  INV_X1 u0_u9_u6_U46 (.A( u0_u9_u6_n144 ) , .ZN( u0_u9_u6_n159 ) );
  NAND2_X1 u0_u9_u6_U47 (.ZN( u0_u9_u6_n145 ) , .A2( u0_u9_u6_n97 ) , .A1( u0_u9_u6_n98 ) );
  NAND2_X1 u0_u9_u6_U48 (.ZN( u0_u9_u6_n148 ) , .A2( u0_u9_u6_n92 ) , .A1( u0_u9_u6_n94 ) );
  NAND2_X1 u0_u9_u6_U49 (.ZN( u0_u9_u6_n108 ) , .A2( u0_u9_u6_n139 ) , .A1( u0_u9_u6_n144 ) );
  NAND2_X1 u0_u9_u6_U5 (.A2( u0_u9_u6_n143 ) , .ZN( u0_u9_u6_n152 ) , .A1( u0_u9_u6_n166 ) );
  NAND2_X1 u0_u9_u6_U50 (.ZN( u0_u9_u6_n121 ) , .A2( u0_u9_u6_n95 ) , .A1( u0_u9_u6_n97 ) );
  NAND2_X1 u0_u9_u6_U51 (.ZN( u0_u9_u6_n107 ) , .A2( u0_u9_u6_n92 ) , .A1( u0_u9_u6_n95 ) );
  AND2_X1 u0_u9_u6_U52 (.ZN( u0_u9_u6_n118 ) , .A2( u0_u9_u6_n91 ) , .A1( u0_u9_u6_n99 ) );
  NAND2_X1 u0_u9_u6_U53 (.ZN( u0_u9_u6_n147 ) , .A2( u0_u9_u6_n98 ) , .A1( u0_u9_u6_n99 ) );
  NAND2_X1 u0_u9_u6_U54 (.ZN( u0_u9_u6_n128 ) , .A1( u0_u9_u6_n94 ) , .A2( u0_u9_u6_n96 ) );
  NAND2_X1 u0_u9_u6_U55 (.ZN( u0_u9_u6_n119 ) , .A2( u0_u9_u6_n95 ) , .A1( u0_u9_u6_n99 ) );
  NAND2_X1 u0_u9_u6_U56 (.ZN( u0_u9_u6_n123 ) , .A2( u0_u9_u6_n91 ) , .A1( u0_u9_u6_n96 ) );
  NAND2_X1 u0_u9_u6_U57 (.ZN( u0_u9_u6_n100 ) , .A2( u0_u9_u6_n92 ) , .A1( u0_u9_u6_n98 ) );
  NAND2_X1 u0_u9_u6_U58 (.ZN( u0_u9_u6_n122 ) , .A1( u0_u9_u6_n94 ) , .A2( u0_u9_u6_n97 ) );
  INV_X1 u0_u9_u6_U59 (.A( u0_u9_u6_n139 ) , .ZN( u0_u9_u6_n160 ) );
  AOI22_X1 u0_u9_u6_U6 (.B2( u0_u9_u6_n101 ) , .A1( u0_u9_u6_n102 ) , .ZN( u0_u9_u6_n103 ) , .B1( u0_u9_u6_n160 ) , .A2( u0_u9_u6_n161 ) );
  NAND2_X1 u0_u9_u6_U60 (.ZN( u0_u9_u6_n113 ) , .A1( u0_u9_u6_n96 ) , .A2( u0_u9_u6_n98 ) );
  NOR2_X1 u0_u9_u6_U61 (.A2( u0_u9_X_40 ) , .A1( u0_u9_X_41 ) , .ZN( u0_u9_u6_n126 ) );
  NOR2_X1 u0_u9_u6_U62 (.A2( u0_u9_X_39 ) , .A1( u0_u9_X_42 ) , .ZN( u0_u9_u6_n92 ) );
  NOR2_X1 u0_u9_u6_U63 (.A2( u0_u9_X_39 ) , .A1( u0_u9_u6_n156 ) , .ZN( u0_u9_u6_n97 ) );
  NOR2_X1 u0_u9_u6_U64 (.A2( u0_u9_X_38 ) , .A1( u0_u9_u6_n165 ) , .ZN( u0_u9_u6_n95 ) );
  NOR2_X1 u0_u9_u6_U65 (.A2( u0_u9_X_41 ) , .ZN( u0_u9_u6_n111 ) , .A1( u0_u9_u6_n157 ) );
  NOR2_X1 u0_u9_u6_U66 (.A2( u0_u9_X_37 ) , .A1( u0_u9_u6_n162 ) , .ZN( u0_u9_u6_n94 ) );
  NOR2_X1 u0_u9_u6_U67 (.A2( u0_u9_X_37 ) , .A1( u0_u9_X_38 ) , .ZN( u0_u9_u6_n91 ) );
  NAND2_X1 u0_u9_u6_U68 (.A1( u0_u9_X_41 ) , .ZN( u0_u9_u6_n144 ) , .A2( u0_u9_u6_n157 ) );
  NAND2_X1 u0_u9_u6_U69 (.A2( u0_u9_X_40 ) , .A1( u0_u9_X_41 ) , .ZN( u0_u9_u6_n139 ) );
  NOR2_X1 u0_u9_u6_U7 (.A1( u0_u9_u6_n118 ) , .ZN( u0_u9_u6_n143 ) , .A2( u0_u9_u6_n168 ) );
  AND2_X1 u0_u9_u6_U70 (.A1( u0_u9_X_39 ) , .A2( u0_u9_u6_n156 ) , .ZN( u0_u9_u6_n96 ) );
  AND2_X1 u0_u9_u6_U71 (.A1( u0_u9_X_39 ) , .A2( u0_u9_X_42 ) , .ZN( u0_u9_u6_n99 ) );
  INV_X1 u0_u9_u6_U72 (.A( u0_u9_X_40 ) , .ZN( u0_u9_u6_n157 ) );
  INV_X1 u0_u9_u6_U73 (.A( u0_u9_X_37 ) , .ZN( u0_u9_u6_n165 ) );
  INV_X1 u0_u9_u6_U74 (.A( u0_u9_X_38 ) , .ZN( u0_u9_u6_n162 ) );
  INV_X1 u0_u9_u6_U75 (.A( u0_u9_X_42 ) , .ZN( u0_u9_u6_n156 ) );
  NAND4_X1 u0_u9_u6_U76 (.ZN( u0_out9_32 ) , .A4( u0_u9_u6_n103 ) , .A3( u0_u9_u6_n104 ) , .A2( u0_u9_u6_n105 ) , .A1( u0_u9_u6_n106 ) );
  AOI22_X1 u0_u9_u6_U77 (.ZN( u0_u9_u6_n105 ) , .A2( u0_u9_u6_n108 ) , .A1( u0_u9_u6_n118 ) , .B2( u0_u9_u6_n126 ) , .B1( u0_u9_u6_n171 ) );
  AOI22_X1 u0_u9_u6_U78 (.ZN( u0_u9_u6_n104 ) , .A1( u0_u9_u6_n111 ) , .B1( u0_u9_u6_n124 ) , .B2( u0_u9_u6_n151 ) , .A2( u0_u9_u6_n93 ) );
  NAND4_X1 u0_u9_u6_U79 (.ZN( u0_out9_12 ) , .A4( u0_u9_u6_n114 ) , .A3( u0_u9_u6_n115 ) , .A2( u0_u9_u6_n116 ) , .A1( u0_u9_u6_n117 ) );
  OAI21_X1 u0_u9_u6_U8 (.A( u0_u9_u6_n159 ) , .B1( u0_u9_u6_n169 ) , .B2( u0_u9_u6_n173 ) , .ZN( u0_u9_u6_n90 ) );
  OAI22_X1 u0_u9_u6_U80 (.B2( u0_u9_u6_n111 ) , .ZN( u0_u9_u6_n116 ) , .B1( u0_u9_u6_n126 ) , .A2( u0_u9_u6_n164 ) , .A1( u0_u9_u6_n167 ) );
  OAI21_X1 u0_u9_u6_U81 (.A( u0_u9_u6_n108 ) , .ZN( u0_u9_u6_n117 ) , .B2( u0_u9_u6_n141 ) , .B1( u0_u9_u6_n163 ) );
  OAI211_X1 u0_u9_u6_U82 (.ZN( u0_out9_7 ) , .B( u0_u9_u6_n153 ) , .C2( u0_u9_u6_n154 ) , .C1( u0_u9_u6_n155 ) , .A( u0_u9_u6_n174 ) );
  NOR3_X1 u0_u9_u6_U83 (.A1( u0_u9_u6_n141 ) , .ZN( u0_u9_u6_n154 ) , .A3( u0_u9_u6_n164 ) , .A2( u0_u9_u6_n171 ) );
  AOI211_X1 u0_u9_u6_U84 (.B( u0_u9_u6_n149 ) , .A( u0_u9_u6_n150 ) , .C2( u0_u9_u6_n151 ) , .C1( u0_u9_u6_n152 ) , .ZN( u0_u9_u6_n153 ) );
  OAI211_X1 u0_u9_u6_U85 (.ZN( u0_out9_22 ) , .B( u0_u9_u6_n137 ) , .A( u0_u9_u6_n138 ) , .C2( u0_u9_u6_n139 ) , .C1( u0_u9_u6_n140 ) );
  AOI22_X1 u0_u9_u6_U86 (.B1( u0_u9_u6_n124 ) , .A2( u0_u9_u6_n125 ) , .A1( u0_u9_u6_n126 ) , .ZN( u0_u9_u6_n138 ) , .B2( u0_u9_u6_n161 ) );
  AND4_X1 u0_u9_u6_U87 (.A3( u0_u9_u6_n119 ) , .A1( u0_u9_u6_n120 ) , .A4( u0_u9_u6_n129 ) , .ZN( u0_u9_u6_n140 ) , .A2( u0_u9_u6_n143 ) );
  NAND3_X1 u0_u9_u6_U88 (.A2( u0_u9_u6_n123 ) , .ZN( u0_u9_u6_n125 ) , .A1( u0_u9_u6_n130 ) , .A3( u0_u9_u6_n131 ) );
  NAND3_X1 u0_u9_u6_U89 (.A3( u0_u9_u6_n133 ) , .ZN( u0_u9_u6_n141 ) , .A1( u0_u9_u6_n145 ) , .A2( u0_u9_u6_n148 ) );
  INV_X1 u0_u9_u6_U9 (.ZN( u0_u9_u6_n172 ) , .A( u0_u9_u6_n88 ) );
  NAND3_X1 u0_u9_u6_U90 (.ZN( u0_u9_u6_n101 ) , .A3( u0_u9_u6_n107 ) , .A2( u0_u9_u6_n121 ) , .A1( u0_u9_u6_n127 ) );
  NAND3_X1 u0_u9_u6_U91 (.ZN( u0_u9_u6_n102 ) , .A3( u0_u9_u6_n130 ) , .A2( u0_u9_u6_n145 ) , .A1( u0_u9_u6_n166 ) );
  NAND3_X1 u0_u9_u6_U92 (.A3( u0_u9_u6_n113 ) , .A1( u0_u9_u6_n119 ) , .A2( u0_u9_u6_n123 ) , .ZN( u0_u9_u6_n93 ) );
  NAND3_X1 u0_u9_u6_U93 (.ZN( u0_u9_u6_n142 ) , .A2( u0_u9_u6_n172 ) , .A3( u0_u9_u6_n89 ) , .A1( u0_u9_u6_n90 ) );
  AND3_X1 u0_u9_u7_U10 (.A3( u0_u9_u7_n110 ) , .A2( u0_u9_u7_n127 ) , .A1( u0_u9_u7_n132 ) , .ZN( u0_u9_u7_n92 ) );
  OAI21_X1 u0_u9_u7_U11 (.A( u0_u9_u7_n161 ) , .B1( u0_u9_u7_n168 ) , .B2( u0_u9_u7_n173 ) , .ZN( u0_u9_u7_n91 ) );
  AOI211_X1 u0_u9_u7_U12 (.A( u0_u9_u7_n117 ) , .ZN( u0_u9_u7_n118 ) , .C2( u0_u9_u7_n126 ) , .C1( u0_u9_u7_n177 ) , .B( u0_u9_u7_n180 ) );
  OAI22_X1 u0_u9_u7_U13 (.B1( u0_u9_u7_n115 ) , .ZN( u0_u9_u7_n117 ) , .A2( u0_u9_u7_n133 ) , .A1( u0_u9_u7_n137 ) , .B2( u0_u9_u7_n162 ) );
  INV_X1 u0_u9_u7_U14 (.A( u0_u9_u7_n116 ) , .ZN( u0_u9_u7_n180 ) );
  NOR3_X1 u0_u9_u7_U15 (.ZN( u0_u9_u7_n115 ) , .A3( u0_u9_u7_n145 ) , .A2( u0_u9_u7_n168 ) , .A1( u0_u9_u7_n169 ) );
  OAI211_X1 u0_u9_u7_U16 (.B( u0_u9_u7_n122 ) , .A( u0_u9_u7_n123 ) , .C2( u0_u9_u7_n124 ) , .ZN( u0_u9_u7_n154 ) , .C1( u0_u9_u7_n162 ) );
  AOI222_X1 u0_u9_u7_U17 (.ZN( u0_u9_u7_n122 ) , .C2( u0_u9_u7_n126 ) , .C1( u0_u9_u7_n145 ) , .B1( u0_u9_u7_n161 ) , .A2( u0_u9_u7_n165 ) , .B2( u0_u9_u7_n170 ) , .A1( u0_u9_u7_n176 ) );
  INV_X1 u0_u9_u7_U18 (.A( u0_u9_u7_n133 ) , .ZN( u0_u9_u7_n176 ) );
  NOR3_X1 u0_u9_u7_U19 (.A2( u0_u9_u7_n134 ) , .A1( u0_u9_u7_n135 ) , .ZN( u0_u9_u7_n136 ) , .A3( u0_u9_u7_n171 ) );
  NOR2_X1 u0_u9_u7_U20 (.A1( u0_u9_u7_n130 ) , .A2( u0_u9_u7_n134 ) , .ZN( u0_u9_u7_n153 ) );
  INV_X1 u0_u9_u7_U21 (.A( u0_u9_u7_n101 ) , .ZN( u0_u9_u7_n165 ) );
  NOR2_X1 u0_u9_u7_U22 (.ZN( u0_u9_u7_n111 ) , .A2( u0_u9_u7_n134 ) , .A1( u0_u9_u7_n169 ) );
  AOI21_X1 u0_u9_u7_U23 (.ZN( u0_u9_u7_n104 ) , .B2( u0_u9_u7_n112 ) , .B1( u0_u9_u7_n127 ) , .A( u0_u9_u7_n164 ) );
  AOI21_X1 u0_u9_u7_U24 (.ZN( u0_u9_u7_n106 ) , .B1( u0_u9_u7_n133 ) , .B2( u0_u9_u7_n146 ) , .A( u0_u9_u7_n162 ) );
  AOI21_X1 u0_u9_u7_U25 (.A( u0_u9_u7_n101 ) , .ZN( u0_u9_u7_n107 ) , .B2( u0_u9_u7_n128 ) , .B1( u0_u9_u7_n175 ) );
  INV_X1 u0_u9_u7_U26 (.A( u0_u9_u7_n138 ) , .ZN( u0_u9_u7_n171 ) );
  INV_X1 u0_u9_u7_U27 (.A( u0_u9_u7_n131 ) , .ZN( u0_u9_u7_n177 ) );
  INV_X1 u0_u9_u7_U28 (.A( u0_u9_u7_n110 ) , .ZN( u0_u9_u7_n174 ) );
  NAND2_X1 u0_u9_u7_U29 (.A1( u0_u9_u7_n129 ) , .A2( u0_u9_u7_n132 ) , .ZN( u0_u9_u7_n149 ) );
  OAI21_X1 u0_u9_u7_U3 (.ZN( u0_u9_u7_n159 ) , .A( u0_u9_u7_n165 ) , .B2( u0_u9_u7_n171 ) , .B1( u0_u9_u7_n174 ) );
  NAND2_X1 u0_u9_u7_U30 (.A1( u0_u9_u7_n113 ) , .A2( u0_u9_u7_n124 ) , .ZN( u0_u9_u7_n130 ) );
  INV_X1 u0_u9_u7_U31 (.A( u0_u9_u7_n112 ) , .ZN( u0_u9_u7_n173 ) );
  INV_X1 u0_u9_u7_U32 (.A( u0_u9_u7_n128 ) , .ZN( u0_u9_u7_n168 ) );
  INV_X1 u0_u9_u7_U33 (.A( u0_u9_u7_n148 ) , .ZN( u0_u9_u7_n169 ) );
  INV_X1 u0_u9_u7_U34 (.A( u0_u9_u7_n127 ) , .ZN( u0_u9_u7_n179 ) );
  NOR2_X1 u0_u9_u7_U35 (.ZN( u0_u9_u7_n101 ) , .A2( u0_u9_u7_n150 ) , .A1( u0_u9_u7_n156 ) );
  AOI211_X1 u0_u9_u7_U36 (.B( u0_u9_u7_n154 ) , .A( u0_u9_u7_n155 ) , .C1( u0_u9_u7_n156 ) , .ZN( u0_u9_u7_n157 ) , .C2( u0_u9_u7_n172 ) );
  INV_X1 u0_u9_u7_U37 (.A( u0_u9_u7_n153 ) , .ZN( u0_u9_u7_n172 ) );
  AOI211_X1 u0_u9_u7_U38 (.B( u0_u9_u7_n139 ) , .A( u0_u9_u7_n140 ) , .C2( u0_u9_u7_n141 ) , .ZN( u0_u9_u7_n142 ) , .C1( u0_u9_u7_n156 ) );
  NAND4_X1 u0_u9_u7_U39 (.A3( u0_u9_u7_n127 ) , .A2( u0_u9_u7_n128 ) , .A1( u0_u9_u7_n129 ) , .ZN( u0_u9_u7_n141 ) , .A4( u0_u9_u7_n147 ) );
  INV_X1 u0_u9_u7_U4 (.A( u0_u9_u7_n111 ) , .ZN( u0_u9_u7_n170 ) );
  AOI21_X1 u0_u9_u7_U40 (.A( u0_u9_u7_n137 ) , .B1( u0_u9_u7_n138 ) , .ZN( u0_u9_u7_n139 ) , .B2( u0_u9_u7_n146 ) );
  OAI22_X1 u0_u9_u7_U41 (.B1( u0_u9_u7_n136 ) , .ZN( u0_u9_u7_n140 ) , .A1( u0_u9_u7_n153 ) , .B2( u0_u9_u7_n162 ) , .A2( u0_u9_u7_n164 ) );
  AOI21_X1 u0_u9_u7_U42 (.ZN( u0_u9_u7_n123 ) , .B1( u0_u9_u7_n165 ) , .B2( u0_u9_u7_n177 ) , .A( u0_u9_u7_n97 ) );
  AOI21_X1 u0_u9_u7_U43 (.B2( u0_u9_u7_n113 ) , .B1( u0_u9_u7_n124 ) , .A( u0_u9_u7_n125 ) , .ZN( u0_u9_u7_n97 ) );
  INV_X1 u0_u9_u7_U44 (.A( u0_u9_u7_n125 ) , .ZN( u0_u9_u7_n161 ) );
  INV_X1 u0_u9_u7_U45 (.A( u0_u9_u7_n152 ) , .ZN( u0_u9_u7_n162 ) );
  AOI22_X1 u0_u9_u7_U46 (.A2( u0_u9_u7_n114 ) , .ZN( u0_u9_u7_n119 ) , .B1( u0_u9_u7_n130 ) , .A1( u0_u9_u7_n156 ) , .B2( u0_u9_u7_n165 ) );
  NAND2_X1 u0_u9_u7_U47 (.A2( u0_u9_u7_n112 ) , .ZN( u0_u9_u7_n114 ) , .A1( u0_u9_u7_n175 ) );
  AND2_X1 u0_u9_u7_U48 (.ZN( u0_u9_u7_n145 ) , .A2( u0_u9_u7_n98 ) , .A1( u0_u9_u7_n99 ) );
  NOR2_X1 u0_u9_u7_U49 (.ZN( u0_u9_u7_n137 ) , .A1( u0_u9_u7_n150 ) , .A2( u0_u9_u7_n161 ) );
  INV_X1 u0_u9_u7_U5 (.A( u0_u9_u7_n149 ) , .ZN( u0_u9_u7_n175 ) );
  AOI21_X1 u0_u9_u7_U50 (.ZN( u0_u9_u7_n105 ) , .B2( u0_u9_u7_n110 ) , .A( u0_u9_u7_n125 ) , .B1( u0_u9_u7_n147 ) );
  NAND2_X1 u0_u9_u7_U51 (.ZN( u0_u9_u7_n146 ) , .A1( u0_u9_u7_n95 ) , .A2( u0_u9_u7_n98 ) );
  NAND2_X1 u0_u9_u7_U52 (.A2( u0_u9_u7_n103 ) , .ZN( u0_u9_u7_n147 ) , .A1( u0_u9_u7_n93 ) );
  NAND2_X1 u0_u9_u7_U53 (.A1( u0_u9_u7_n103 ) , .ZN( u0_u9_u7_n127 ) , .A2( u0_u9_u7_n99 ) );
  OR2_X1 u0_u9_u7_U54 (.ZN( u0_u9_u7_n126 ) , .A2( u0_u9_u7_n152 ) , .A1( u0_u9_u7_n156 ) );
  NAND2_X1 u0_u9_u7_U55 (.A2( u0_u9_u7_n102 ) , .A1( u0_u9_u7_n103 ) , .ZN( u0_u9_u7_n133 ) );
  NAND2_X1 u0_u9_u7_U56 (.ZN( u0_u9_u7_n112 ) , .A2( u0_u9_u7_n96 ) , .A1( u0_u9_u7_n99 ) );
  NAND2_X1 u0_u9_u7_U57 (.A2( u0_u9_u7_n102 ) , .ZN( u0_u9_u7_n128 ) , .A1( u0_u9_u7_n98 ) );
  NAND2_X1 u0_u9_u7_U58 (.A1( u0_u9_u7_n100 ) , .ZN( u0_u9_u7_n113 ) , .A2( u0_u9_u7_n93 ) );
  NAND2_X1 u0_u9_u7_U59 (.A2( u0_u9_u7_n102 ) , .ZN( u0_u9_u7_n124 ) , .A1( u0_u9_u7_n96 ) );
  INV_X1 u0_u9_u7_U6 (.A( u0_u9_u7_n154 ) , .ZN( u0_u9_u7_n178 ) );
  NAND2_X1 u0_u9_u7_U60 (.ZN( u0_u9_u7_n110 ) , .A1( u0_u9_u7_n95 ) , .A2( u0_u9_u7_n96 ) );
  INV_X1 u0_u9_u7_U61 (.A( u0_u9_u7_n150 ) , .ZN( u0_u9_u7_n164 ) );
  AND2_X1 u0_u9_u7_U62 (.ZN( u0_u9_u7_n134 ) , .A1( u0_u9_u7_n93 ) , .A2( u0_u9_u7_n98 ) );
  NAND2_X1 u0_u9_u7_U63 (.A1( u0_u9_u7_n100 ) , .A2( u0_u9_u7_n102 ) , .ZN( u0_u9_u7_n129 ) );
  NAND2_X1 u0_u9_u7_U64 (.A2( u0_u9_u7_n103 ) , .ZN( u0_u9_u7_n131 ) , .A1( u0_u9_u7_n95 ) );
  NAND2_X1 u0_u9_u7_U65 (.A1( u0_u9_u7_n100 ) , .ZN( u0_u9_u7_n138 ) , .A2( u0_u9_u7_n99 ) );
  NAND2_X1 u0_u9_u7_U66 (.ZN( u0_u9_u7_n132 ) , .A1( u0_u9_u7_n93 ) , .A2( u0_u9_u7_n96 ) );
  NAND2_X1 u0_u9_u7_U67 (.A1( u0_u9_u7_n100 ) , .ZN( u0_u9_u7_n148 ) , .A2( u0_u9_u7_n95 ) );
  NOR2_X1 u0_u9_u7_U68 (.A2( u0_u9_X_47 ) , .ZN( u0_u9_u7_n150 ) , .A1( u0_u9_u7_n163 ) );
  NOR2_X1 u0_u9_u7_U69 (.A2( u0_u9_X_43 ) , .A1( u0_u9_X_44 ) , .ZN( u0_u9_u7_n103 ) );
  AOI211_X1 u0_u9_u7_U7 (.ZN( u0_u9_u7_n116 ) , .A( u0_u9_u7_n155 ) , .C1( u0_u9_u7_n161 ) , .C2( u0_u9_u7_n171 ) , .B( u0_u9_u7_n94 ) );
  NOR2_X1 u0_u9_u7_U70 (.A2( u0_u9_X_48 ) , .A1( u0_u9_u7_n166 ) , .ZN( u0_u9_u7_n95 ) );
  NOR2_X1 u0_u9_u7_U71 (.A2( u0_u9_X_45 ) , .A1( u0_u9_X_48 ) , .ZN( u0_u9_u7_n99 ) );
  NOR2_X1 u0_u9_u7_U72 (.A2( u0_u9_X_44 ) , .A1( u0_u9_u7_n167 ) , .ZN( u0_u9_u7_n98 ) );
  NOR2_X1 u0_u9_u7_U73 (.A2( u0_u9_X_46 ) , .A1( u0_u9_X_47 ) , .ZN( u0_u9_u7_n152 ) );
  AND2_X1 u0_u9_u7_U74 (.A1( u0_u9_X_47 ) , .ZN( u0_u9_u7_n156 ) , .A2( u0_u9_u7_n163 ) );
  NAND2_X1 u0_u9_u7_U75 (.A2( u0_u9_X_46 ) , .A1( u0_u9_X_47 ) , .ZN( u0_u9_u7_n125 ) );
  AND2_X1 u0_u9_u7_U76 (.A2( u0_u9_X_45 ) , .A1( u0_u9_X_48 ) , .ZN( u0_u9_u7_n102 ) );
  AND2_X1 u0_u9_u7_U77 (.A2( u0_u9_X_43 ) , .A1( u0_u9_X_44 ) , .ZN( u0_u9_u7_n96 ) );
  AND2_X1 u0_u9_u7_U78 (.A1( u0_u9_X_44 ) , .ZN( u0_u9_u7_n100 ) , .A2( u0_u9_u7_n167 ) );
  AND2_X1 u0_u9_u7_U79 (.A1( u0_u9_X_48 ) , .A2( u0_u9_u7_n166 ) , .ZN( u0_u9_u7_n93 ) );
  OAI222_X1 u0_u9_u7_U8 (.C2( u0_u9_u7_n101 ) , .B2( u0_u9_u7_n111 ) , .A1( u0_u9_u7_n113 ) , .C1( u0_u9_u7_n146 ) , .A2( u0_u9_u7_n162 ) , .B1( u0_u9_u7_n164 ) , .ZN( u0_u9_u7_n94 ) );
  INV_X1 u0_u9_u7_U80 (.A( u0_u9_X_46 ) , .ZN( u0_u9_u7_n163 ) );
  INV_X1 u0_u9_u7_U81 (.A( u0_u9_X_45 ) , .ZN( u0_u9_u7_n166 ) );
  INV_X1 u0_u9_u7_U82 (.A( u0_u9_X_43 ) , .ZN( u0_u9_u7_n167 ) );
  NAND4_X1 u0_u9_u7_U83 (.ZN( u0_out9_27 ) , .A4( u0_u9_u7_n118 ) , .A3( u0_u9_u7_n119 ) , .A2( u0_u9_u7_n120 ) , .A1( u0_u9_u7_n121 ) );
  OAI21_X1 u0_u9_u7_U84 (.ZN( u0_u9_u7_n121 ) , .B2( u0_u9_u7_n145 ) , .A( u0_u9_u7_n150 ) , .B1( u0_u9_u7_n174 ) );
  OAI21_X1 u0_u9_u7_U85 (.ZN( u0_u9_u7_n120 ) , .A( u0_u9_u7_n161 ) , .B2( u0_u9_u7_n170 ) , .B1( u0_u9_u7_n179 ) );
  NAND4_X1 u0_u9_u7_U86 (.ZN( u0_out9_21 ) , .A4( u0_u9_u7_n157 ) , .A3( u0_u9_u7_n158 ) , .A2( u0_u9_u7_n159 ) , .A1( u0_u9_u7_n160 ) );
  OAI21_X1 u0_u9_u7_U87 (.B1( u0_u9_u7_n145 ) , .ZN( u0_u9_u7_n160 ) , .A( u0_u9_u7_n161 ) , .B2( u0_u9_u7_n177 ) );
  AOI22_X1 u0_u9_u7_U88 (.B2( u0_u9_u7_n149 ) , .B1( u0_u9_u7_n150 ) , .A2( u0_u9_u7_n151 ) , .A1( u0_u9_u7_n152 ) , .ZN( u0_u9_u7_n158 ) );
  NAND4_X1 u0_u9_u7_U89 (.ZN( u0_out9_15 ) , .A4( u0_u9_u7_n142 ) , .A3( u0_u9_u7_n143 ) , .A2( u0_u9_u7_n144 ) , .A1( u0_u9_u7_n178 ) );
  OAI221_X1 u0_u9_u7_U9 (.C1( u0_u9_u7_n101 ) , .C2( u0_u9_u7_n147 ) , .ZN( u0_u9_u7_n155 ) , .B2( u0_u9_u7_n162 ) , .A( u0_u9_u7_n91 ) , .B1( u0_u9_u7_n92 ) );
  OR2_X1 u0_u9_u7_U90 (.A2( u0_u9_u7_n125 ) , .A1( u0_u9_u7_n129 ) , .ZN( u0_u9_u7_n144 ) );
  AOI22_X1 u0_u9_u7_U91 (.A2( u0_u9_u7_n126 ) , .ZN( u0_u9_u7_n143 ) , .B2( u0_u9_u7_n165 ) , .B1( u0_u9_u7_n173 ) , .A1( u0_u9_u7_n174 ) );
  NAND4_X1 u0_u9_u7_U92 (.ZN( u0_out9_5 ) , .A4( u0_u9_u7_n108 ) , .A3( u0_u9_u7_n109 ) , .A1( u0_u9_u7_n116 ) , .A2( u0_u9_u7_n123 ) );
  AOI22_X1 u0_u9_u7_U93 (.ZN( u0_u9_u7_n109 ) , .A2( u0_u9_u7_n126 ) , .B2( u0_u9_u7_n145 ) , .B1( u0_u9_u7_n156 ) , .A1( u0_u9_u7_n171 ) );
  NOR4_X1 u0_u9_u7_U94 (.A4( u0_u9_u7_n104 ) , .A3( u0_u9_u7_n105 ) , .A2( u0_u9_u7_n106 ) , .A1( u0_u9_u7_n107 ) , .ZN( u0_u9_u7_n108 ) );
  NAND3_X1 u0_u9_u7_U95 (.A3( u0_u9_u7_n146 ) , .A2( u0_u9_u7_n147 ) , .A1( u0_u9_u7_n148 ) , .ZN( u0_u9_u7_n151 ) );
  NAND3_X1 u0_u9_u7_U96 (.A3( u0_u9_u7_n131 ) , .A2( u0_u9_u7_n132 ) , .A1( u0_u9_u7_n133 ) , .ZN( u0_u9_u7_n135 ) );
  OAI22_X1 u0_uk_U102 (.ZN( u0_K7_5 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n162 ) , .A2( u0_uk_n384 ) , .B2( u0_uk_n401 ) );
  OAI21_X1 u0_uk_U104 (.ZN( u0_K4_5 ) , .B1( u0_uk_n10 ) , .B2( u0_uk_n502 ) , .A( u0_uk_n821 ) );
  NAND2_X1 u0_uk_U105 (.A1( u0_uk_K_r2_53 ) , .ZN( u0_uk_n821 ) , .A2( u0_uk_n99 ) );
  OAI21_X1 u0_uk_U1050 (.ZN( u0_K15_32 ) , .B1( u0_uk_n31 ) , .B2( u0_uk_n33 ) , .A( u0_uk_n918 ) );
  OAI21_X1 u0_uk_U1058 (.ZN( u0_K4_38 ) , .B1( u0_uk_n27 ) , .B2( u0_uk_n505 ) , .A( u0_uk_n825 ) );
  NAND2_X1 u0_uk_U1059 (.A1( u0_uk_K_r2_50 ) , .A2( u0_uk_n63 ) , .ZN( u0_uk_n825 ) );
  OAI21_X1 u0_uk_U1087 (.ZN( u0_K8_14 ) , .B1( u0_uk_n250 ) , .B2( u0_uk_n329 ) , .A( u0_uk_n760 ) );
  NAND2_X1 u0_uk_U1088 (.A1( u0_uk_K_r6_34 ) , .A2( u0_uk_n202 ) , .ZN( u0_uk_n760 ) );
  INV_X1 u0_uk_U1113 (.ZN( u0_K8_12 ) , .A( u0_uk_n761 ) );
  INV_X1 u0_uk_U1121 (.ZN( u0_K5_20 ) , .A( u0_uk_n816 ) );
  INV_X1 u0_uk_U1123 (.ZN( u0_K7_13 ) , .A( u0_uk_n783 ) );
  INV_X1 u0_uk_U1135 (.ZN( u0_K4_2 ) , .A( u0_uk_n828 ) );
  AOI22_X1 u0_uk_U1136 (.B2( u0_uk_K_r2_26 ) , .A2( u0_uk_K_r2_46 ) , .B1( u0_uk_n129 ) , .A1( u0_uk_n148 ) , .ZN( u0_uk_n828 ) );
  INV_X1 u0_uk_U1137 (.ZN( u0_K4_20 ) , .A( u0_uk_n835 ) );
  AOI22_X1 u0_uk_U1138 (.B2( u0_uk_K_r2_13 ) , .A2( u0_uk_K_r2_33 ) , .B1( u0_uk_n129 ) , .A1( u0_uk_n208 ) , .ZN( u0_uk_n835 ) );
  INV_X1 u0_uk_U1141 (.ZN( u0_K10_12 ) , .A( u0_uk_n1024 ) );
  INV_X1 u0_uk_U1145 (.ZN( u0_K8_15 ) , .A( u0_uk_n759 ) );
  INV_X1 u0_uk_U1147 (.ZN( u0_K5_35 ) , .A( u0_uk_n810 ) );
  OAI21_X1 u0_uk_U1151 (.ZN( u0_K5_6 ) , .B1( u0_uk_n109 ) , .B2( u0_uk_n471 ) , .A( u0_uk_n803 ) );
  NAND2_X1 u0_uk_U1152 (.A1( u0_uk_K_r3_10 ) , .ZN( u0_uk_n803 ) , .A2( u0_uk_n93 ) );
  OAI22_X1 u0_uk_U117 (.ZN( u0_K10_47 ) , .A1( u0_uk_n109 ) , .B1( u0_uk_n214 ) , .B2( u0_uk_n249 ) , .A2( u0_uk_n264 ) );
  OAI22_X1 u0_uk_U123 (.ZN( u0_K4_47 ) , .A1( u0_uk_n161 ) , .A2( u0_uk_n499 ) , .B2( u0_uk_n508 ) , .B1( u0_uk_n93 ) );
  OAI22_X1 u0_uk_U127 (.ZN( u0_K4_15 ) , .A1( u0_uk_n242 ) , .A2( u0_uk_n502 ) , .B2( u0_uk_n530 ) , .B1( u0_uk_n83 ) );
  OAI22_X1 u0_uk_U155 (.ZN( u0_K7_19 ) , .A1( u0_uk_n162 ) , .B1( u0_uk_n31 ) , .A2( u0_uk_n383 ) , .B2( u0_uk_n393 ) );
  OAI22_X1 u0_uk_U156 (.ZN( u0_K4_19 ) , .A1( u0_uk_n129 ) , .B1( u0_uk_n148 ) , .A2( u0_uk_n511 ) , .B2( u0_uk_n523 ) );
  OAI22_X1 u0_uk_U169 (.ZN( u0_K10_30 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n214 ) , .A2( u0_uk_n232 ) , .B2( u0_uk_n260 ) );
  OAI21_X1 u0_uk_U182 (.ZN( u0_K10_24 ) , .A( u0_uk_n1017 ) , .B1( u0_uk_n11 ) , .B2( u0_uk_n259 ) );
  NAND2_X1 u0_uk_U183 (.A1( u0_uk_K_r8_40 ) , .ZN( u0_uk_n1017 ) , .A2( u0_uk_n11 ) );
  OAI21_X1 u0_uk_U205 (.ZN( u0_K4_30 ) , .B1( u0_uk_n252 ) , .B2( u0_uk_n513 ) , .A( u0_uk_n827 ) );
  NAND2_X1 u0_uk_U206 (.A1( u0_uk_K_r2_28 ) , .A2( u0_uk_n202 ) , .ZN( u0_uk_n827 ) );
  INV_X1 u0_uk_U207 (.ZN( u0_K15_30 ) , .A( u0_uk_n919 ) );
  AOI22_X1 u0_uk_U208 (.B2( u0_uk_K_r13_0 ) , .A2( u0_uk_K_r13_38 ) , .B1( u0_uk_n142 ) , .A1( u0_uk_n217 ) , .ZN( u0_uk_n919 ) );
  OAI22_X1 u0_uk_U225 (.ZN( u0_K13_31 ) , .B2( u0_uk_n116 ) , .A1( u0_uk_n209 ) , .B1( u0_uk_n92 ) , .A2( u0_uk_n98 ) );
  OAI21_X1 u0_uk_U226 (.ZN( u0_K10_31 ) , .A( u0_uk_n1014 ) , .B2( u0_uk_n243 ) , .B1( u0_uk_n250 ) );
  NAND2_X1 u0_uk_U227 (.A1( u0_uk_K_r8_16 ) , .ZN( u0_uk_n1014 ) , .A2( u0_uk_n207 ) );
  OAI22_X1 u0_uk_U230 (.ZN( u0_K15_31 ) , .A1( u0_uk_n187 ) , .A2( u0_uk_n28 ) , .B2( u0_uk_n45 ) , .B1( u0_uk_n92 ) );
  OAI22_X1 u0_uk_U234 (.ZN( u0_K14_31 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n240 ) , .A2( u0_uk_n55 ) , .B2( u0_uk_n61 ) );
  OAI22_X1 u0_uk_U236 (.ZN( u0_K15_39 ) , .A1( u0_uk_n128 ) , .B2( u0_uk_n22 ) , .B1( u0_uk_n220 ) , .A2( u0_uk_n40 ) );
  OAI22_X1 u0_uk_U244 (.ZN( u0_K15_44 ) , .A1( u0_uk_n155 ) , .B1( u0_uk_n17 ) , .B2( u0_uk_n22 ) , .A2( u0_uk_n4 ) );
  OAI22_X1 u0_uk_U262 (.ZN( u0_K10_44 ) , .A1( u0_uk_n162 ) , .A2( u0_uk_n241 ) , .B2( u0_uk_n261 ) , .B1( u0_uk_n83 ) );
  OAI22_X1 u0_uk_U263 (.ZN( u0_K10_48 ) , .A2( u0_uk_n232 ) , .A1( u0_uk_n240 ) , .B2( u0_uk_n248 ) , .B1( u0_uk_n94 ) );
  OAI22_X1 u0_uk_U278 (.ZN( u0_K10_6 ) , .B1( u0_uk_n102 ) , .A1( u0_uk_n162 ) , .B2( u0_uk_n239 ) , .A2( u0_uk_n267 ) );
  OAI22_X1 u0_uk_U287 (.ZN( u0_K8_8 ) , .A1( u0_uk_n162 ) , .B1( u0_uk_n27 ) , .A2( u0_uk_n324 ) , .B2( u0_uk_n330 ) );
  INV_X1 u0_uk_U288 (.ZN( u0_K7_8 ) , .A( u0_uk_n763 ) );
  INV_X1 u0_uk_U291 (.ZN( u0_K4_8 ) , .A( u0_uk_n819 ) );
  AOI22_X1 u0_uk_U292 (.B2( u0_uk_K_r2_41 ) , .A2( u0_uk_K_r2_46 ) , .A1( u0_uk_n146 ) , .B1( u0_uk_n203 ) , .ZN( u0_uk_n819 ) );
  INV_X1 u0_uk_U304 (.ZN( u0_K15_26 ) , .A( u0_uk_n920 ) );
  AOI22_X1 u0_uk_U305 (.B2( u0_uk_K_r13_38 ) , .A2( u0_uk_K_r13_44 ) , .B1( u0_uk_n129 ) , .A1( u0_uk_n251 ) , .ZN( u0_uk_n920 ) );
  OAI22_X1 u0_uk_U317 (.ZN( u0_K10_26 ) , .B1( u0_uk_n142 ) , .A1( u0_uk_n213 ) , .A2( u0_uk_n233 ) , .B2( u0_uk_n249 ) );
  OAI22_X1 u0_uk_U320 (.ZN( u0_K15_46 ) , .B2( u0_uk_n13 ) , .B1( u0_uk_n17 ) , .A1( u0_uk_n187 ) , .A2( u0_uk_n40 ) );
  OAI22_X1 u0_uk_U340 (.ZN( u0_K7_4 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n161 ) , .A2( u0_uk_n361 ) , .B2( u0_uk_n384 ) );
  INV_X1 u0_uk_U345 (.ZN( u0_K4_4 ) , .A( u0_uk_n822 ) );
  AOI22_X1 u0_uk_U346 (.B2( u0_uk_K_r2_13 ) , .A2( u0_uk_K_r2_18 ) , .B1( u0_uk_n203 ) , .ZN( u0_uk_n822 ) , .A1( u0_uk_n94 ) );
  INV_X1 u0_uk_U355 (.ZN( u0_K10_40 ) , .A( u0_uk_n1006 ) );
  OAI22_X1 u0_uk_U360 (.ZN( u0_K15_40 ) , .A1( u0_uk_n155 ) , .B1( u0_uk_n17 ) , .A2( u0_uk_n41 ) , .B2( u0_uk_n9 ) );
  OAI21_X1 u0_uk_U367 (.ZN( u0_K15_33 ) , .B2( u0_uk_n18 ) , .B1( u0_uk_n83 ) , .A( u0_uk_n917 ) );
  OAI22_X1 u0_uk_U373 (.ZN( u0_K14_28 ) , .A1( u0_uk_n109 ) , .B1( u0_uk_n203 ) , .A2( u0_uk_n61 ) , .B2( u0_uk_n67 ) );
  OAI21_X1 u0_uk_U379 (.ZN( u0_K5_33 ) , .B1( u0_uk_n250 ) , .B2( u0_uk_n457 ) , .A( u0_uk_n811 ) );
  NAND2_X1 u0_uk_U380 (.A1( u0_uk_K_r3_14 ) , .A2( u0_uk_n220 ) , .ZN( u0_uk_n811 ) );
  OAI22_X1 u0_uk_U381 (.ZN( u0_K15_28 ) , .A1( u0_uk_n128 ) , .B1( u0_uk_n230 ) , .B2( u0_uk_n33 ) , .A2( u0_uk_n5 ) );
  OAI22_X1 u0_uk_U383 (.ZN( u0_K10_28 ) , .A1( u0_uk_n100 ) , .B1( u0_uk_n182 ) , .A2( u0_uk_n241 ) , .B2( u0_uk_n248 ) );
  OAI22_X1 u0_uk_U396 (.ZN( u0_K8_16 ) , .A1( u0_uk_n213 ) , .A2( u0_uk_n344 ) , .B2( u0_uk_n352 ) , .B1( u0_uk_n63 ) );
  OAI22_X1 u0_uk_U401 (.ZN( u0_K4_16 ) , .B1( u0_uk_n128 ) , .A1( u0_uk_n238 ) , .A2( u0_uk_n525 ) , .B2( u0_uk_n529 ) );
  INV_X1 u0_uk_U416 (.ZN( u0_K10_9 ) , .A( u0_uk_n1005 ) );
  OAI22_X1 u0_uk_U421 (.ZN( u0_K4_9 ) , .A1( u0_uk_n146 ) , .B1( u0_uk_n217 ) , .A2( u0_uk_n519 ) , .B2( u0_uk_n529 ) );
  INV_X1 u0_uk_U439 (.ZN( u0_K10_33 ) , .A( u0_uk_n1012 ) );
  OAI22_X1 u0_uk_U444 (.ZN( u0_K14_33 ) , .A1( u0_uk_n230 ) , .A2( u0_uk_n55 ) , .B2( u0_uk_n73 ) , .B1( u0_uk_n94 ) );
  OAI22_X1 u0_uk_U449 (.ZN( u0_K4_33 ) , .B1( u0_uk_n110 ) , .A1( u0_uk_n148 ) , .A2( u0_uk_n532 ) , .B2( u0_uk_n539 ) );
  OAI22_X1 u0_uk_U451 (.ZN( u0_K14_37 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n231 ) , .A2( u0_uk_n67 ) , .B2( u0_uk_n73 ) );
  OAI22_X1 u0_uk_U454 (.ZN( u0_K15_37 ) , .B2( u0_uk_n12 ) , .A1( u0_uk_n187 ) , .B1( u0_uk_n27 ) , .A2( u0_uk_n39 ) );
  BUF_X1 u0_uk_U46 (.A( u0_uk_n162 ) , .Z( u0_uk_n223 ) );
  OAI22_X1 u0_uk_U474 (.ZN( u0_K13_29 ) , .A2( u0_uk_n113 ) , .B2( u0_uk_n116 ) , .A1( u0_uk_n118 ) , .B1( u0_uk_n161 ) );
  OAI22_X1 u0_uk_U482 (.ZN( u0_K15_29 ) , .A1( u0_uk_n128 ) , .B1( u0_uk_n188 ) , .B2( u0_uk_n21 ) , .A2( u0_uk_n39 ) );
  OAI22_X1 u0_uk_U483 (.ZN( u0_K10_29 ) , .A1( u0_uk_n100 ) , .B1( u0_uk_n214 ) , .A2( u0_uk_n233 ) , .B2( u0_uk_n261 ) );
  BUF_X1 u0_uk_U50 (.A( u0_uk_n162 ) , .Z( u0_uk_n213 ) );
  OAI21_X1 u0_uk_U510 (.ZN( u0_K8_17 ) , .B1( u0_uk_n252 ) , .B2( u0_uk_n336 ) , .A( u0_uk_n758 ) );
  NAND2_X1 u0_uk_U511 (.A1( u0_uk_K_r6_26 ) , .A2( u0_uk_n220 ) , .ZN( u0_uk_n758 ) );
  OAI22_X1 u0_uk_U512 (.ZN( u0_K7_17 ) , .A1( u0_uk_n161 ) , .B1( u0_uk_n31 ) , .A2( u0_uk_n370 ) , .B2( u0_uk_n400 ) );
  OAI21_X1 u0_uk_U513 (.ZN( u0_K4_17 ) , .B1( u0_uk_n250 ) , .B2( u0_uk_n519 ) , .A( u0_uk_n838 ) );
  NAND2_X1 u0_uk_U514 (.A1( u0_uk_K_r2_27 ) , .A2( u0_uk_n208 ) , .ZN( u0_uk_n838 ) );
  INV_X1 u0_uk_U522 (.ZN( u0_K7_12 ) , .A( u0_uk_n784 ) );
  AOI22_X1 u0_uk_U523 (.B2( u0_uk_K_r5_17 ) , .A2( u0_uk_K_r5_39 ) , .B1( u0_uk_n146 ) , .A1( u0_uk_n223 ) , .ZN( u0_uk_n784 ) );
  OAI22_X1 u0_uk_U526 (.ZN( u0_K4_12 ) , .A1( u0_uk_n10 ) , .B1( u0_uk_n161 ) , .A2( u0_uk_n497 ) , .B2( u0_uk_n517 ) );
  OAI22_X1 u0_uk_U544 (.ZN( u0_K15_36 ) , .A1( u0_uk_n155 ) , .A2( u0_uk_n18 ) , .B1( u0_uk_n27 ) , .B2( u0_uk_n32 ) );
  INV_X1 u0_uk_U550 (.ZN( u0_K5_36 ) , .A( u0_uk_n809 ) );
  INV_X1 u0_uk_U558 (.ZN( u0_K7_36 ) , .A( u0_uk_n768 ) );
  INV_X1 u0_uk_U562 (.ZN( u0_K15_38 ) , .A( u0_uk_n916 ) );
  OAI22_X1 u0_uk_U581 (.ZN( u0_K8_10 ) , .A1( u0_uk_n223 ) , .B1( u0_uk_n31 ) , .A2( u0_uk_n337 ) , .B2( u0_uk_n339 ) );
  INV_X1 u0_uk_U584 (.ZN( u0_K4_10 ) , .A( u0_uk_n839 ) );
  INV_X1 u0_uk_U599 (.ZN( u0_K5_22 ) , .A( u0_uk_n815 ) );
  OAI22_X1 u0_uk_U611 (.ZN( u0_K15_35 ) , .A2( u0_uk_n13 ) , .A1( u0_uk_n187 ) , .B1( u0_uk_n27 ) , .B2( u0_uk_n28 ) );
  INV_X1 u0_uk_U612 (.ZN( u0_K14_35 ) , .A( u0_uk_n933 ) );
  OAI22_X1 u0_uk_U633 (.ZN( u0_K7_11 ) , .A1( u0_uk_n109 ) , .B1( u0_uk_n214 ) , .A2( u0_uk_n383 ) , .B2( u0_uk_n400 ) );
  OAI22_X1 u0_uk_U64 (.ZN( u0_K15_34 ) , .A1( u0_uk_n128 ) , .B1( u0_uk_n230 ) , .B2( u0_uk_n32 ) , .A2( u0_uk_n4 ) );
  INV_X1 u0_uk_U643 (.ZN( u0_K4_23 ) , .A( u0_uk_n833 ) );
  AOI22_X1 u0_uk_U644 (.B2( u0_uk_K_r2_18 ) , .A2( u0_uk_K_r2_55 ) , .B1( u0_uk_n207 ) , .ZN( u0_uk_n833 ) , .A1( u0_uk_n94 ) );
  INV_X1 u0_uk_U65 (.ZN( u0_K14_34 ) , .A( u0_uk_n934 ) );
  INV_X1 u0_uk_U660 (.ZN( u0_K15_43 ) , .A( u0_uk_n915 ) );
  OAI22_X1 u0_uk_U670 (.ZN( u0_K10_45 ) , .A1( u0_uk_n223 ) , .A2( u0_uk_n244 ) , .B2( u0_uk_n260 ) , .B1( u0_uk_n94 ) );
  OAI22_X1 u0_uk_U684 (.ZN( u0_K4_7 ) , .B1( u0_uk_n202 ) , .B2( u0_uk_n531 ) , .A2( u0_uk_n535 ) , .A1( u0_uk_n99 ) );
  OAI22_X1 u0_uk_U689 (.ZN( u0_K13_25 ) , .A1( u0_uk_n118 ) , .B2( u0_uk_n123 ) , .B1( u0_uk_n242 ) , .A2( u0_uk_n98 ) );
  INV_X1 u0_uk_U702 (.ZN( u0_K4_3 ) , .A( u0_uk_n824 ) );
  AOI22_X1 u0_uk_U703 (.A2( u0_uk_K_r2_4 ) , .B2( u0_uk_K_r2_41 ) , .A1( u0_uk_n238 ) , .ZN( u0_uk_n824 ) , .B1( u0_uk_n99 ) );
  INV_X1 u0_uk_U712 (.ZN( u0_K4_25 ) , .A( u0_uk_n832 ) );
  OAI21_X1 u0_uk_U714 (.ZN( u0_K10_2 ) , .A( u0_uk_n1015 ) , .B1( u0_uk_n250 ) , .B2( u0_uk_n266 ) );
  NAND2_X1 u0_uk_U715 (.A1( u0_uk_K_r8_41 ) , .ZN( u0_uk_n1015 ) , .A2( u0_uk_n220 ) );
  OAI22_X1 u0_uk_U716 (.ZN( u0_K4_32 ) , .A1( u0_uk_n142 ) , .B1( u0_uk_n163 ) , .B2( u0_uk_n508 ) , .A2( u0_uk_n532 ) );
  OAI22_X1 u0_uk_U726 (.ZN( u0_K15_42 ) , .A1( u0_uk_n141 ) , .B1( u0_uk_n220 ) , .A2( u0_uk_n3 ) , .B2( u0_uk_n9 ) );
  OAI22_X1 u0_uk_U730 (.ZN( u0_K10_42 ) , .A1( u0_uk_n102 ) , .B1( u0_uk_n238 ) , .A2( u0_uk_n243 ) , .B2( u0_uk_n269 ) );
  OAI22_X1 u0_uk_U766 (.ZN( u0_K4_21 ) , .B1( u0_uk_n146 ) , .A1( u0_uk_n238 ) , .A2( u0_uk_n511 ) , .B2( u0_uk_n517 ) );
  OAI22_X1 u0_uk_U771 (.ZN( u0_K15_27 ) , .A1( u0_uk_n128 ) , .B1( u0_uk_n188 ) , .B2( u0_uk_n23 ) , .A2( u0_uk_n41 ) );
  OAI22_X1 u0_uk_U772 (.ZN( u0_K4_13 ) , .B1( u0_uk_n240 ) , .B2( u0_uk_n530 ) , .A2( u0_uk_n534 ) , .A1( u0_uk_n60 ) );
  INV_X1 u0_uk_U774 (.ZN( u0_K5_27 ) , .A( u0_uk_n813 ) );
  OAI21_X1 u0_uk_U800 (.ZN( u0_K7_1 ) , .B1( u0_uk_n250 ) , .B2( u0_uk_n396 ) , .A( u0_uk_n781 ) );
  NAND2_X1 u0_uk_U801 (.A1( u0_uk_K_r5_10 ) , .A2( u0_uk_n147 ) , .ZN( u0_uk_n781 ) );
  OAI21_X1 u0_uk_U802 (.ZN( u0_K4_1 ) , .B1( u0_uk_n252 ) , .B2( u0_uk_n535 ) , .A( u0_uk_n836 ) );
  NAND2_X1 u0_uk_U803 (.A1( u0_uk_K_r2_25 ) , .A2( u0_uk_n207 ) , .ZN( u0_uk_n836 ) );
  OAI21_X1 u0_uk_U804 (.ZN( u0_K4_18 ) , .B2( u0_uk_n510 ) , .A( u0_uk_n837 ) , .B1( u0_uk_n92 ) );
  NAND2_X1 u0_uk_U805 (.A1( u0_uk_K_r2_20 ) , .A2( u0_uk_n31 ) , .ZN( u0_uk_n837 ) );
  OAI22_X1 u0_uk_U807 (.ZN( u0_K7_18 ) , .A1( u0_uk_n213 ) , .B1( u0_uk_n31 ) , .B2( u0_uk_n392 ) , .A2( u0_uk_n405 ) );
  OAI21_X1 u0_uk_U812 (.ZN( u0_K8_18 ) , .B2( u0_uk_n331 ) , .A( u0_uk_n757 ) , .B1( u0_uk_n93 ) );
  NAND2_X1 u0_uk_U813 (.A1( u0_uk_K_r6_46 ) , .A2( u0_uk_n10 ) , .ZN( u0_uk_n757 ) );
  OAI22_X1 u0_uk_U824 (.ZN( u0_K8_20 ) , .B1( u0_uk_n110 ) , .A1( u0_uk_n213 ) , .A2( u0_uk_n331 ) , .B2( u0_uk_n337 ) );
  INV_X1 u0_uk_U833 (.ZN( u0_K7_20 ) , .A( u0_uk_n780 ) );
  OAI22_X1 u0_uk_U849 (.ZN( u0_K7_3 ) , .A1( u0_uk_n141 ) , .B1( u0_uk_n188 ) , .A2( u0_uk_n371 ) , .B2( u0_uk_n393 ) );
  INV_X1 u0_uk_U854 (.ZN( u0_K7_6 ) , .A( u0_uk_n764 ) );
  AOI22_X1 u0_uk_U855 (.B2( u0_uk_K_r5_39 ) , .A2( u0_uk_K_r5_4 ) , .B1( u0_uk_n145 ) , .A1( u0_uk_n213 ) , .ZN( u0_uk_n764 ) );
  OAI22_X1 u0_uk_U879 (.ZN( u0_K8_5 ) , .A1( u0_uk_n223 ) , .B1( u0_uk_n27 ) , .A2( u0_uk_n318 ) , .B2( u0_uk_n324 ) );
  OAI22_X1 u0_uk_U88 (.ZN( u0_K15_41 ) , .B1( u0_uk_n17 ) , .A1( u0_uk_n187 ) , .B2( u0_uk_n23 ) , .A2( u0_uk_n5 ) );
  OAI22_X1 u0_uk_U883 (.ZN( u0_K7_10 ) , .A1( u0_uk_n161 ) , .A2( u0_uk_n371 ) , .B2( u0_uk_n401 ) , .B1( u0_uk_n60 ) );
  OAI22_X1 u0_uk_U884 (.ZN( u0_K4_11 ) , .B1( u0_uk_n117 ) , .A1( u0_uk_n164 ) , .A2( u0_uk_n497 ) , .B2( u0_uk_n525 ) );
  OAI22_X1 u0_uk_U886 (.ZN( u0_K15_45 ) , .A1( u0_uk_n155 ) , .B1( u0_uk_n17 ) , .B2( u0_uk_n21 ) , .A2( u0_uk_n3 ) );
  OAI22_X1 u0_uk_U891 (.ZN( u0_K8_6 ) , .A1( u0_uk_n162 ) , .B1( u0_uk_n27 ) , .A2( u0_uk_n339 ) , .B2( u0_uk_n344 ) );
  OAI22_X1 u0_uk_U898 (.ZN( u0_K7_14 ) , .A1( u0_uk_n213 ) , .B1( u0_uk_n31 ) , .A2( u0_uk_n361 ) , .B2( u0_uk_n396 ) );
  OAI22_X1 u0_uk_U909 (.ZN( u0_K8_21 ) , .B1( u0_uk_n102 ) , .A1( u0_uk_n257 ) , .A2( u0_uk_n330 ) , .B2( u0_uk_n336 ) );
  OAI22_X1 u0_uk_U91 (.ZN( u0_K4_41 ) , .A1( u0_uk_n109 ) , .B1( u0_uk_n163 ) , .A2( u0_uk_n522 ) , .B2( u0_uk_n539 ) );
  OAI22_X1 u0_uk_U914 (.ZN( u0_K4_14 ) , .A1( u0_uk_n164 ) , .A2( u0_uk_n510 ) , .B2( u0_uk_n536 ) , .B1( u0_uk_n99 ) );
  OAI22_X1 u0_uk_U944 (.ZN( u0_K8_24 ) , .A1( u0_uk_n102 ) , .B1( u0_uk_n213 ) , .A2( u0_uk_n318 ) , .B2( u0_uk_n358 ) );
  OAI22_X1 u0_uk_U956 (.ZN( u0_K10_8 ) , .A1( u0_uk_n109 ) , .B1( u0_uk_n182 ) , .B2( u0_uk_n253 ) , .A2( u0_uk_n267 ) );
  OAI22_X1 u0_uk_U983 (.ZN( u0_K8_7 ) , .A1( u0_uk_n100 ) , .B1( u0_uk_n257 ) , .B2( u0_uk_n352 ) , .A2( u0_uk_n358 ) );
  OAI22_X1 u0_uk_U984 (.ZN( u0_K7_7 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n257 ) , .A2( u0_uk_n370 ) , .B2( u0_uk_n392 ) );
  XOR2_X1 u2_u0_U11 (.B( u2_K1_44 ) , .A( u2_desIn_r_33 ) , .Z( u2_u0_X_44 ) );
  XOR2_X1 u2_u0_U12 (.B( u2_K1_43 ) , .A( u2_desIn_r_25 ) , .Z( u2_u0_X_43 ) );
  XOR2_X1 u2_u0_U13 (.B( u2_K1_42 ) , .A( u2_desIn_r_33 ) , .Z( u2_u0_X_42 ) );
  XOR2_X1 u2_u0_U14 (.B( u2_K1_41 ) , .A( u2_desIn_r_25 ) , .Z( u2_u0_X_41 ) );
  XOR2_X1 u2_u0_U18 (.B( u2_K1_38 ) , .A( u2_desIn_r_1 ) , .Z( u2_u0_X_38 ) );
  XOR2_X1 u2_u0_U20 (.B( u2_K1_36 ) , .A( u2_desIn_r_1 ) , .Z( u2_u0_X_36 ) );
  XOR2_X1 u2_u0_U25 (.B( u2_K1_31 ) , .A( u2_desIn_r_27 ) , .Z( u2_u0_X_31 ) );
  XOR2_X1 u2_u0_U28 (.B( u2_K1_29 ) , .A( u2_desIn_r_27 ) , .Z( u2_u0_X_29 ) );
  XOR2_X1 u2_u0_U8 (.B( u2_K1_47 ) , .A( u2_desIn_r_57 ) , .Z( u2_u0_X_47 ) );
  AOI21_X1 u2_u0_u1_U10 (.B2( u2_u0_u1_n155 ) , .B1( u2_u0_u1_n156 ) , .ZN( u2_u0_u1_n157 ) , .A( u2_u0_u1_n174 ) );
  NAND3_X1 u2_u0_u1_U100 (.ZN( u2_u0_u1_n113 ) , .A1( u2_u0_u1_n120 ) , .A3( u2_u0_u1_n133 ) , .A2( u2_u0_u1_n155 ) );
  NAND2_X1 u2_u0_u1_U11 (.ZN( u2_u0_u1_n140 ) , .A2( u2_u0_u1_n150 ) , .A1( u2_u0_u1_n155 ) );
  NAND2_X1 u2_u0_u1_U12 (.A1( u2_u0_u1_n131 ) , .ZN( u2_u0_u1_n147 ) , .A2( u2_u0_u1_n153 ) );
  AOI22_X1 u2_u0_u1_U13 (.B2( u2_u0_u1_n136 ) , .A2( u2_u0_u1_n137 ) , .ZN( u2_u0_u1_n143 ) , .A1( u2_u0_u1_n171 ) , .B1( u2_u0_u1_n173 ) );
  INV_X1 u2_u0_u1_U14 (.A( u2_u0_u1_n147 ) , .ZN( u2_u0_u1_n181 ) );
  INV_X1 u2_u0_u1_U15 (.A( u2_u0_u1_n139 ) , .ZN( u2_u0_u1_n174 ) );
  OR4_X1 u2_u0_u1_U16 (.A4( u2_u0_u1_n106 ) , .A3( u2_u0_u1_n107 ) , .ZN( u2_u0_u1_n108 ) , .A1( u2_u0_u1_n117 ) , .A2( u2_u0_u1_n184 ) );
  AOI21_X1 u2_u0_u1_U17 (.ZN( u2_u0_u1_n106 ) , .A( u2_u0_u1_n112 ) , .B1( u2_u0_u1_n154 ) , .B2( u2_u0_u1_n156 ) );
  AOI21_X1 u2_u0_u1_U18 (.ZN( u2_u0_u1_n107 ) , .B1( u2_u0_u1_n134 ) , .B2( u2_u0_u1_n149 ) , .A( u2_u0_u1_n174 ) );
  INV_X1 u2_u0_u1_U19 (.A( u2_u0_u1_n101 ) , .ZN( u2_u0_u1_n184 ) );
  INV_X1 u2_u0_u1_U20 (.A( u2_u0_u1_n112 ) , .ZN( u2_u0_u1_n171 ) );
  NAND2_X1 u2_u0_u1_U21 (.ZN( u2_u0_u1_n141 ) , .A1( u2_u0_u1_n153 ) , .A2( u2_u0_u1_n156 ) );
  AND2_X1 u2_u0_u1_U22 (.A1( u2_u0_u1_n123 ) , .ZN( u2_u0_u1_n134 ) , .A2( u2_u0_u1_n161 ) );
  NAND2_X1 u2_u0_u1_U23 (.A2( u2_u0_u1_n115 ) , .A1( u2_u0_u1_n116 ) , .ZN( u2_u0_u1_n148 ) );
  NAND2_X1 u2_u0_u1_U24 (.A2( u2_u0_u1_n133 ) , .A1( u2_u0_u1_n135 ) , .ZN( u2_u0_u1_n159 ) );
  NAND2_X1 u2_u0_u1_U25 (.A2( u2_u0_u1_n115 ) , .A1( u2_u0_u1_n120 ) , .ZN( u2_u0_u1_n132 ) );
  INV_X1 u2_u0_u1_U26 (.A( u2_u0_u1_n154 ) , .ZN( u2_u0_u1_n178 ) );
  INV_X1 u2_u0_u1_U27 (.A( u2_u0_u1_n151 ) , .ZN( u2_u0_u1_n183 ) );
  AND2_X1 u2_u0_u1_U28 (.A1( u2_u0_u1_n129 ) , .A2( u2_u0_u1_n133 ) , .ZN( u2_u0_u1_n149 ) );
  INV_X1 u2_u0_u1_U29 (.A( u2_u0_u1_n131 ) , .ZN( u2_u0_u1_n180 ) );
  INV_X1 u2_u0_u1_U3 (.A( u2_u0_u1_n159 ) , .ZN( u2_u0_u1_n182 ) );
  AOI221_X1 u2_u0_u1_U30 (.B1( u2_u0_u1_n140 ) , .ZN( u2_u0_u1_n167 ) , .B2( u2_u0_u1_n172 ) , .C2( u2_u0_u1_n175 ) , .C1( u2_u0_u1_n178 ) , .A( u2_u0_u1_n188 ) );
  INV_X1 u2_u0_u1_U31 (.ZN( u2_u0_u1_n188 ) , .A( u2_u0_u1_n97 ) );
  AOI211_X1 u2_u0_u1_U32 (.A( u2_u0_u1_n118 ) , .C1( u2_u0_u1_n132 ) , .C2( u2_u0_u1_n139 ) , .B( u2_u0_u1_n96 ) , .ZN( u2_u0_u1_n97 ) );
  AOI21_X1 u2_u0_u1_U33 (.B2( u2_u0_u1_n121 ) , .B1( u2_u0_u1_n135 ) , .A( u2_u0_u1_n152 ) , .ZN( u2_u0_u1_n96 ) );
  OAI221_X1 u2_u0_u1_U34 (.A( u2_u0_u1_n119 ) , .C2( u2_u0_u1_n129 ) , .ZN( u2_u0_u1_n138 ) , .B2( u2_u0_u1_n152 ) , .C1( u2_u0_u1_n174 ) , .B1( u2_u0_u1_n187 ) );
  INV_X1 u2_u0_u1_U35 (.A( u2_u0_u1_n148 ) , .ZN( u2_u0_u1_n187 ) );
  AOI211_X1 u2_u0_u1_U36 (.B( u2_u0_u1_n117 ) , .A( u2_u0_u1_n118 ) , .ZN( u2_u0_u1_n119 ) , .C2( u2_u0_u1_n146 ) , .C1( u2_u0_u1_n159 ) );
  NOR2_X1 u2_u0_u1_U37 (.A1( u2_u0_u1_n168 ) , .A2( u2_u0_u1_n176 ) , .ZN( u2_u0_u1_n98 ) );
  AOI211_X1 u2_u0_u1_U38 (.B( u2_u0_u1_n162 ) , .A( u2_u0_u1_n163 ) , .C2( u2_u0_u1_n164 ) , .ZN( u2_u0_u1_n165 ) , .C1( u2_u0_u1_n171 ) );
  AOI21_X1 u2_u0_u1_U39 (.A( u2_u0_u1_n160 ) , .B2( u2_u0_u1_n161 ) , .ZN( u2_u0_u1_n162 ) , .B1( u2_u0_u1_n182 ) );
  AOI221_X1 u2_u0_u1_U4 (.A( u2_u0_u1_n138 ) , .C2( u2_u0_u1_n139 ) , .C1( u2_u0_u1_n140 ) , .B2( u2_u0_u1_n141 ) , .ZN( u2_u0_u1_n142 ) , .B1( u2_u0_u1_n175 ) );
  OR2_X1 u2_u0_u1_U40 (.A2( u2_u0_u1_n157 ) , .A1( u2_u0_u1_n158 ) , .ZN( u2_u0_u1_n163 ) );
  NAND2_X1 u2_u0_u1_U41 (.A1( u2_u0_u1_n128 ) , .ZN( u2_u0_u1_n146 ) , .A2( u2_u0_u1_n160 ) );
  NAND2_X1 u2_u0_u1_U42 (.A2( u2_u0_u1_n112 ) , .ZN( u2_u0_u1_n139 ) , .A1( u2_u0_u1_n152 ) );
  NAND2_X1 u2_u0_u1_U43 (.A1( u2_u0_u1_n105 ) , .ZN( u2_u0_u1_n156 ) , .A2( u2_u0_u1_n99 ) );
  NOR2_X1 u2_u0_u1_U44 (.ZN( u2_u0_u1_n117 ) , .A1( u2_u0_u1_n121 ) , .A2( u2_u0_u1_n160 ) );
  AOI21_X1 u2_u0_u1_U45 (.A( u2_u0_u1_n128 ) , .B2( u2_u0_u1_n129 ) , .ZN( u2_u0_u1_n130 ) , .B1( u2_u0_u1_n150 ) );
  NAND2_X1 u2_u0_u1_U46 (.ZN( u2_u0_u1_n112 ) , .A1( u2_u0_u1_n169 ) , .A2( u2_u0_u1_n170 ) );
  NAND2_X1 u2_u0_u1_U47 (.ZN( u2_u0_u1_n129 ) , .A2( u2_u0_u1_n95 ) , .A1( u2_u0_u1_n98 ) );
  NAND2_X1 u2_u0_u1_U48 (.A1( u2_u0_u1_n102 ) , .ZN( u2_u0_u1_n154 ) , .A2( u2_u0_u1_n99 ) );
  NAND2_X1 u2_u0_u1_U49 (.A2( u2_u0_u1_n100 ) , .ZN( u2_u0_u1_n135 ) , .A1( u2_u0_u1_n99 ) );
  AOI211_X1 u2_u0_u1_U5 (.ZN( u2_u0_u1_n124 ) , .A( u2_u0_u1_n138 ) , .C2( u2_u0_u1_n139 ) , .B( u2_u0_u1_n145 ) , .C1( u2_u0_u1_n147 ) );
  AOI21_X1 u2_u0_u1_U50 (.A( u2_u0_u1_n152 ) , .B2( u2_u0_u1_n153 ) , .B1( u2_u0_u1_n154 ) , .ZN( u2_u0_u1_n158 ) );
  INV_X1 u2_u0_u1_U51 (.A( u2_u0_u1_n160 ) , .ZN( u2_u0_u1_n175 ) );
  NAND2_X1 u2_u0_u1_U52 (.A1( u2_u0_u1_n100 ) , .ZN( u2_u0_u1_n116 ) , .A2( u2_u0_u1_n95 ) );
  NAND2_X1 u2_u0_u1_U53 (.A1( u2_u0_u1_n102 ) , .ZN( u2_u0_u1_n131 ) , .A2( u2_u0_u1_n95 ) );
  NAND2_X1 u2_u0_u1_U54 (.A2( u2_u0_u1_n104 ) , .ZN( u2_u0_u1_n121 ) , .A1( u2_u0_u1_n98 ) );
  NAND2_X1 u2_u0_u1_U55 (.A1( u2_u0_u1_n103 ) , .ZN( u2_u0_u1_n153 ) , .A2( u2_u0_u1_n98 ) );
  NAND2_X1 u2_u0_u1_U56 (.A2( u2_u0_u1_n104 ) , .A1( u2_u0_u1_n105 ) , .ZN( u2_u0_u1_n133 ) );
  NAND2_X1 u2_u0_u1_U57 (.ZN( u2_u0_u1_n150 ) , .A2( u2_u0_u1_n98 ) , .A1( u2_u0_u1_n99 ) );
  NAND2_X1 u2_u0_u1_U58 (.A1( u2_u0_u1_n105 ) , .ZN( u2_u0_u1_n155 ) , .A2( u2_u0_u1_n95 ) );
  OAI21_X1 u2_u0_u1_U59 (.ZN( u2_u0_u1_n109 ) , .B1( u2_u0_u1_n129 ) , .B2( u2_u0_u1_n160 ) , .A( u2_u0_u1_n167 ) );
  AOI22_X1 u2_u0_u1_U6 (.B2( u2_u0_u1_n113 ) , .A2( u2_u0_u1_n114 ) , .ZN( u2_u0_u1_n125 ) , .A1( u2_u0_u1_n171 ) , .B1( u2_u0_u1_n173 ) );
  NAND2_X1 u2_u0_u1_U60 (.A2( u2_u0_u1_n100 ) , .A1( u2_u0_u1_n103 ) , .ZN( u2_u0_u1_n120 ) );
  NAND2_X1 u2_u0_u1_U61 (.A1( u2_u0_u1_n102 ) , .A2( u2_u0_u1_n104 ) , .ZN( u2_u0_u1_n115 ) );
  NAND2_X1 u2_u0_u1_U62 (.A2( u2_u0_u1_n100 ) , .A1( u2_u0_u1_n104 ) , .ZN( u2_u0_u1_n151 ) );
  NAND2_X1 u2_u0_u1_U63 (.A2( u2_u0_u1_n103 ) , .A1( u2_u0_u1_n105 ) , .ZN( u2_u0_u1_n161 ) );
  INV_X1 u2_u0_u1_U64 (.A( u2_u0_u1_n152 ) , .ZN( u2_u0_u1_n173 ) );
  INV_X1 u2_u0_u1_U65 (.A( u2_u0_u1_n128 ) , .ZN( u2_u0_u1_n172 ) );
  NAND2_X1 u2_u0_u1_U66 (.A2( u2_u0_u1_n102 ) , .A1( u2_u0_u1_n103 ) , .ZN( u2_u0_u1_n123 ) );
  OAI21_X1 u2_u0_u1_U67 (.B2( u2_u0_u1_n123 ) , .ZN( u2_u0_u1_n145 ) , .B1( u2_u0_u1_n160 ) , .A( u2_u0_u1_n185 ) );
  INV_X1 u2_u0_u1_U68 (.A( u2_u0_u1_n122 ) , .ZN( u2_u0_u1_n185 ) );
  AOI21_X1 u2_u0_u1_U69 (.B2( u2_u0_u1_n120 ) , .B1( u2_u0_u1_n121 ) , .ZN( u2_u0_u1_n122 ) , .A( u2_u0_u1_n128 ) );
  NAND2_X1 u2_u0_u1_U7 (.ZN( u2_u0_u1_n114 ) , .A1( u2_u0_u1_n134 ) , .A2( u2_u0_u1_n156 ) );
  NOR2_X1 u2_u0_u1_U70 (.A2( u2_u0_X_7 ) , .A1( u2_u0_X_8 ) , .ZN( u2_u0_u1_n95 ) );
  NOR2_X1 u2_u0_u1_U71 (.A1( u2_u0_X_12 ) , .A2( u2_u0_X_9 ) , .ZN( u2_u0_u1_n100 ) );
  NOR2_X1 u2_u0_u1_U72 (.A2( u2_u0_X_8 ) , .A1( u2_u0_u1_n177 ) , .ZN( u2_u0_u1_n99 ) );
  NOR2_X1 u2_u0_u1_U73 (.A2( u2_u0_X_12 ) , .ZN( u2_u0_u1_n102 ) , .A1( u2_u0_u1_n176 ) );
  NOR2_X1 u2_u0_u1_U74 (.A2( u2_u0_X_9 ) , .ZN( u2_u0_u1_n105 ) , .A1( u2_u0_u1_n168 ) );
  NAND2_X1 u2_u0_u1_U75 (.A1( u2_u0_X_10 ) , .ZN( u2_u0_u1_n160 ) , .A2( u2_u0_u1_n169 ) );
  NAND2_X1 u2_u0_u1_U76 (.A2( u2_u0_X_10 ) , .A1( u2_u0_X_11 ) , .ZN( u2_u0_u1_n152 ) );
  NAND2_X1 u2_u0_u1_U77 (.A1( u2_u0_X_11 ) , .ZN( u2_u0_u1_n128 ) , .A2( u2_u0_u1_n170 ) );
  AND2_X1 u2_u0_u1_U78 (.A2( u2_u0_X_7 ) , .A1( u2_u0_X_8 ) , .ZN( u2_u0_u1_n104 ) );
  AND2_X1 u2_u0_u1_U79 (.A1( u2_u0_X_8 ) , .ZN( u2_u0_u1_n103 ) , .A2( u2_u0_u1_n177 ) );
  NOR2_X1 u2_u0_u1_U8 (.A1( u2_u0_u1_n112 ) , .A2( u2_u0_u1_n116 ) , .ZN( u2_u0_u1_n118 ) );
  INV_X1 u2_u0_u1_U80 (.A( u2_u0_X_10 ) , .ZN( u2_u0_u1_n170 ) );
  INV_X1 u2_u0_u1_U81 (.A( u2_u0_X_9 ) , .ZN( u2_u0_u1_n176 ) );
  INV_X1 u2_u0_u1_U82 (.A( u2_u0_X_11 ) , .ZN( u2_u0_u1_n169 ) );
  INV_X1 u2_u0_u1_U83 (.A( u2_u0_X_12 ) , .ZN( u2_u0_u1_n168 ) );
  INV_X1 u2_u0_u1_U84 (.A( u2_u0_X_7 ) , .ZN( u2_u0_u1_n177 ) );
  NAND4_X1 u2_u0_u1_U85 (.ZN( u2_out0_28 ) , .A4( u2_u0_u1_n124 ) , .A3( u2_u0_u1_n125 ) , .A2( u2_u0_u1_n126 ) , .A1( u2_u0_u1_n127 ) );
  OAI21_X1 u2_u0_u1_U86 (.ZN( u2_u0_u1_n127 ) , .B2( u2_u0_u1_n139 ) , .B1( u2_u0_u1_n175 ) , .A( u2_u0_u1_n183 ) );
  OAI21_X1 u2_u0_u1_U87 (.ZN( u2_u0_u1_n126 ) , .B2( u2_u0_u1_n140 ) , .A( u2_u0_u1_n146 ) , .B1( u2_u0_u1_n178 ) );
  NAND4_X1 u2_u0_u1_U88 (.ZN( u2_out0_18 ) , .A4( u2_u0_u1_n165 ) , .A3( u2_u0_u1_n166 ) , .A1( u2_u0_u1_n167 ) , .A2( u2_u0_u1_n186 ) );
  AOI22_X1 u2_u0_u1_U89 (.B2( u2_u0_u1_n146 ) , .B1( u2_u0_u1_n147 ) , .A2( u2_u0_u1_n148 ) , .ZN( u2_u0_u1_n166 ) , .A1( u2_u0_u1_n172 ) );
  OAI21_X1 u2_u0_u1_U9 (.ZN( u2_u0_u1_n101 ) , .B1( u2_u0_u1_n141 ) , .A( u2_u0_u1_n146 ) , .B2( u2_u0_u1_n183 ) );
  INV_X1 u2_u0_u1_U90 (.A( u2_u0_u1_n145 ) , .ZN( u2_u0_u1_n186 ) );
  NAND4_X1 u2_u0_u1_U91 (.ZN( u2_out0_2 ) , .A4( u2_u0_u1_n142 ) , .A3( u2_u0_u1_n143 ) , .A2( u2_u0_u1_n144 ) , .A1( u2_u0_u1_n179 ) );
  OAI21_X1 u2_u0_u1_U92 (.B2( u2_u0_u1_n132 ) , .ZN( u2_u0_u1_n144 ) , .A( u2_u0_u1_n146 ) , .B1( u2_u0_u1_n180 ) );
  INV_X1 u2_u0_u1_U93 (.A( u2_u0_u1_n130 ) , .ZN( u2_u0_u1_n179 ) );
  OR4_X1 u2_u0_u1_U94 (.ZN( u2_out0_13 ) , .A4( u2_u0_u1_n108 ) , .A3( u2_u0_u1_n109 ) , .A2( u2_u0_u1_n110 ) , .A1( u2_u0_u1_n111 ) );
  AOI21_X1 u2_u0_u1_U95 (.ZN( u2_u0_u1_n111 ) , .A( u2_u0_u1_n128 ) , .B2( u2_u0_u1_n131 ) , .B1( u2_u0_u1_n135 ) );
  AOI21_X1 u2_u0_u1_U96 (.ZN( u2_u0_u1_n110 ) , .A( u2_u0_u1_n116 ) , .B1( u2_u0_u1_n152 ) , .B2( u2_u0_u1_n160 ) );
  NAND3_X1 u2_u0_u1_U97 (.A3( u2_u0_u1_n149 ) , .A2( u2_u0_u1_n150 ) , .A1( u2_u0_u1_n151 ) , .ZN( u2_u0_u1_n164 ) );
  NAND3_X1 u2_u0_u1_U98 (.A3( u2_u0_u1_n134 ) , .A2( u2_u0_u1_n135 ) , .ZN( u2_u0_u1_n136 ) , .A1( u2_u0_u1_n151 ) );
  NAND3_X1 u2_u0_u1_U99 (.A1( u2_u0_u1_n133 ) , .ZN( u2_u0_u1_n137 ) , .A2( u2_u0_u1_n154 ) , .A3( u2_u0_u1_n181 ) );
  OAI22_X1 u2_u0_u4_U10 (.B2( u2_u0_u4_n135 ) , .ZN( u2_u0_u4_n137 ) , .B1( u2_u0_u4_n153 ) , .A1( u2_u0_u4_n155 ) , .A2( u2_u0_u4_n171 ) );
  AND3_X1 u2_u0_u4_U11 (.A2( u2_u0_u4_n134 ) , .ZN( u2_u0_u4_n135 ) , .A3( u2_u0_u4_n145 ) , .A1( u2_u0_u4_n157 ) );
  NAND2_X1 u2_u0_u4_U12 (.ZN( u2_u0_u4_n132 ) , .A2( u2_u0_u4_n170 ) , .A1( u2_u0_u4_n173 ) );
  AOI21_X1 u2_u0_u4_U13 (.B2( u2_u0_u4_n160 ) , .B1( u2_u0_u4_n161 ) , .ZN( u2_u0_u4_n162 ) , .A( u2_u0_u4_n170 ) );
  AOI21_X1 u2_u0_u4_U14 (.ZN( u2_u0_u4_n107 ) , .B2( u2_u0_u4_n143 ) , .A( u2_u0_u4_n174 ) , .B1( u2_u0_u4_n184 ) );
  AOI21_X1 u2_u0_u4_U15 (.B2( u2_u0_u4_n158 ) , .B1( u2_u0_u4_n159 ) , .ZN( u2_u0_u4_n163 ) , .A( u2_u0_u4_n174 ) );
  AOI21_X1 u2_u0_u4_U16 (.A( u2_u0_u4_n153 ) , .B2( u2_u0_u4_n154 ) , .B1( u2_u0_u4_n155 ) , .ZN( u2_u0_u4_n165 ) );
  AOI21_X1 u2_u0_u4_U17 (.A( u2_u0_u4_n156 ) , .B2( u2_u0_u4_n157 ) , .ZN( u2_u0_u4_n164 ) , .B1( u2_u0_u4_n184 ) );
  INV_X1 u2_u0_u4_U18 (.A( u2_u0_u4_n138 ) , .ZN( u2_u0_u4_n170 ) );
  AND2_X1 u2_u0_u4_U19 (.A2( u2_u0_u4_n120 ) , .ZN( u2_u0_u4_n155 ) , .A1( u2_u0_u4_n160 ) );
  INV_X1 u2_u0_u4_U20 (.A( u2_u0_u4_n156 ) , .ZN( u2_u0_u4_n175 ) );
  NAND2_X1 u2_u0_u4_U21 (.A2( u2_u0_u4_n118 ) , .ZN( u2_u0_u4_n131 ) , .A1( u2_u0_u4_n147 ) );
  NAND2_X1 u2_u0_u4_U22 (.A1( u2_u0_u4_n119 ) , .A2( u2_u0_u4_n120 ) , .ZN( u2_u0_u4_n130 ) );
  NAND2_X1 u2_u0_u4_U23 (.ZN( u2_u0_u4_n117 ) , .A2( u2_u0_u4_n118 ) , .A1( u2_u0_u4_n148 ) );
  NAND2_X1 u2_u0_u4_U24 (.ZN( u2_u0_u4_n129 ) , .A1( u2_u0_u4_n134 ) , .A2( u2_u0_u4_n148 ) );
  AND3_X1 u2_u0_u4_U25 (.A1( u2_u0_u4_n119 ) , .A2( u2_u0_u4_n143 ) , .A3( u2_u0_u4_n154 ) , .ZN( u2_u0_u4_n161 ) );
  AND2_X1 u2_u0_u4_U26 (.A1( u2_u0_u4_n145 ) , .A2( u2_u0_u4_n147 ) , .ZN( u2_u0_u4_n159 ) );
  OR3_X1 u2_u0_u4_U27 (.A3( u2_u0_u4_n114 ) , .A2( u2_u0_u4_n115 ) , .A1( u2_u0_u4_n116 ) , .ZN( u2_u0_u4_n136 ) );
  AOI21_X1 u2_u0_u4_U28 (.A( u2_u0_u4_n113 ) , .ZN( u2_u0_u4_n116 ) , .B2( u2_u0_u4_n173 ) , .B1( u2_u0_u4_n174 ) );
  AOI21_X1 u2_u0_u4_U29 (.ZN( u2_u0_u4_n115 ) , .B2( u2_u0_u4_n145 ) , .B1( u2_u0_u4_n146 ) , .A( u2_u0_u4_n156 ) );
  NOR2_X1 u2_u0_u4_U3 (.ZN( u2_u0_u4_n121 ) , .A1( u2_u0_u4_n181 ) , .A2( u2_u0_u4_n182 ) );
  OAI22_X1 u2_u0_u4_U30 (.ZN( u2_u0_u4_n114 ) , .A2( u2_u0_u4_n121 ) , .B1( u2_u0_u4_n160 ) , .B2( u2_u0_u4_n170 ) , .A1( u2_u0_u4_n171 ) );
  INV_X1 u2_u0_u4_U31 (.A( u2_u0_u4_n158 ) , .ZN( u2_u0_u4_n182 ) );
  INV_X1 u2_u0_u4_U32 (.ZN( u2_u0_u4_n181 ) , .A( u2_u0_u4_n96 ) );
  INV_X1 u2_u0_u4_U33 (.A( u2_u0_u4_n144 ) , .ZN( u2_u0_u4_n179 ) );
  INV_X1 u2_u0_u4_U34 (.A( u2_u0_u4_n157 ) , .ZN( u2_u0_u4_n178 ) );
  NAND2_X1 u2_u0_u4_U35 (.A2( u2_u0_u4_n154 ) , .A1( u2_u0_u4_n96 ) , .ZN( u2_u0_u4_n97 ) );
  INV_X1 u2_u0_u4_U36 (.ZN( u2_u0_u4_n186 ) , .A( u2_u0_u4_n95 ) );
  OAI221_X1 u2_u0_u4_U37 (.C1( u2_u0_u4_n134 ) , .B1( u2_u0_u4_n158 ) , .B2( u2_u0_u4_n171 ) , .C2( u2_u0_u4_n173 ) , .A( u2_u0_u4_n94 ) , .ZN( u2_u0_u4_n95 ) );
  AOI222_X1 u2_u0_u4_U38 (.B2( u2_u0_u4_n132 ) , .A1( u2_u0_u4_n138 ) , .C2( u2_u0_u4_n175 ) , .A2( u2_u0_u4_n179 ) , .C1( u2_u0_u4_n181 ) , .B1( u2_u0_u4_n185 ) , .ZN( u2_u0_u4_n94 ) );
  INV_X1 u2_u0_u4_U39 (.A( u2_u0_u4_n113 ) , .ZN( u2_u0_u4_n185 ) );
  INV_X1 u2_u0_u4_U4 (.A( u2_u0_u4_n117 ) , .ZN( u2_u0_u4_n184 ) );
  INV_X1 u2_u0_u4_U40 (.A( u2_u0_u4_n143 ) , .ZN( u2_u0_u4_n183 ) );
  NOR2_X1 u2_u0_u4_U41 (.ZN( u2_u0_u4_n138 ) , .A1( u2_u0_u4_n168 ) , .A2( u2_u0_u4_n169 ) );
  NOR2_X1 u2_u0_u4_U42 (.A1( u2_u0_u4_n150 ) , .A2( u2_u0_u4_n152 ) , .ZN( u2_u0_u4_n153 ) );
  NOR2_X1 u2_u0_u4_U43 (.A2( u2_u0_u4_n128 ) , .A1( u2_u0_u4_n138 ) , .ZN( u2_u0_u4_n156 ) );
  AOI22_X1 u2_u0_u4_U44 (.B2( u2_u0_u4_n122 ) , .A1( u2_u0_u4_n123 ) , .ZN( u2_u0_u4_n124 ) , .B1( u2_u0_u4_n128 ) , .A2( u2_u0_u4_n172 ) );
  INV_X1 u2_u0_u4_U45 (.A( u2_u0_u4_n153 ) , .ZN( u2_u0_u4_n172 ) );
  NAND2_X1 u2_u0_u4_U46 (.A2( u2_u0_u4_n120 ) , .ZN( u2_u0_u4_n123 ) , .A1( u2_u0_u4_n161 ) );
  AOI22_X1 u2_u0_u4_U47 (.B2( u2_u0_u4_n132 ) , .A2( u2_u0_u4_n133 ) , .ZN( u2_u0_u4_n140 ) , .A1( u2_u0_u4_n150 ) , .B1( u2_u0_u4_n179 ) );
  NAND2_X1 u2_u0_u4_U48 (.ZN( u2_u0_u4_n133 ) , .A2( u2_u0_u4_n146 ) , .A1( u2_u0_u4_n154 ) );
  NAND2_X1 u2_u0_u4_U49 (.A1( u2_u0_u4_n103 ) , .ZN( u2_u0_u4_n154 ) , .A2( u2_u0_u4_n98 ) );
  NOR4_X1 u2_u0_u4_U5 (.A4( u2_u0_u4_n106 ) , .A3( u2_u0_u4_n107 ) , .A2( u2_u0_u4_n108 ) , .A1( u2_u0_u4_n109 ) , .ZN( u2_u0_u4_n110 ) );
  NAND2_X1 u2_u0_u4_U50 (.A1( u2_u0_u4_n101 ) , .ZN( u2_u0_u4_n158 ) , .A2( u2_u0_u4_n99 ) );
  AOI21_X1 u2_u0_u4_U51 (.ZN( u2_u0_u4_n127 ) , .A( u2_u0_u4_n136 ) , .B2( u2_u0_u4_n150 ) , .B1( u2_u0_u4_n180 ) );
  INV_X1 u2_u0_u4_U52 (.A( u2_u0_u4_n160 ) , .ZN( u2_u0_u4_n180 ) );
  NAND2_X1 u2_u0_u4_U53 (.A2( u2_u0_u4_n104 ) , .A1( u2_u0_u4_n105 ) , .ZN( u2_u0_u4_n146 ) );
  NAND2_X1 u2_u0_u4_U54 (.A2( u2_u0_u4_n101 ) , .A1( u2_u0_u4_n102 ) , .ZN( u2_u0_u4_n160 ) );
  NAND2_X1 u2_u0_u4_U55 (.ZN( u2_u0_u4_n134 ) , .A1( u2_u0_u4_n98 ) , .A2( u2_u0_u4_n99 ) );
  NAND2_X1 u2_u0_u4_U56 (.A1( u2_u0_u4_n103 ) , .A2( u2_u0_u4_n104 ) , .ZN( u2_u0_u4_n143 ) );
  NAND2_X1 u2_u0_u4_U57 (.A2( u2_u0_u4_n105 ) , .ZN( u2_u0_u4_n145 ) , .A1( u2_u0_u4_n98 ) );
  NAND2_X1 u2_u0_u4_U58 (.A1( u2_u0_u4_n100 ) , .A2( u2_u0_u4_n105 ) , .ZN( u2_u0_u4_n120 ) );
  NAND2_X1 u2_u0_u4_U59 (.A1( u2_u0_u4_n102 ) , .A2( u2_u0_u4_n104 ) , .ZN( u2_u0_u4_n148 ) );
  AOI21_X1 u2_u0_u4_U6 (.ZN( u2_u0_u4_n106 ) , .B2( u2_u0_u4_n146 ) , .B1( u2_u0_u4_n158 ) , .A( u2_u0_u4_n170 ) );
  NAND2_X1 u2_u0_u4_U60 (.A2( u2_u0_u4_n100 ) , .A1( u2_u0_u4_n103 ) , .ZN( u2_u0_u4_n157 ) );
  INV_X1 u2_u0_u4_U61 (.A( u2_u0_u4_n150 ) , .ZN( u2_u0_u4_n173 ) );
  INV_X1 u2_u0_u4_U62 (.A( u2_u0_u4_n152 ) , .ZN( u2_u0_u4_n171 ) );
  NAND2_X1 u2_u0_u4_U63 (.A1( u2_u0_u4_n100 ) , .ZN( u2_u0_u4_n118 ) , .A2( u2_u0_u4_n99 ) );
  NAND2_X1 u2_u0_u4_U64 (.A2( u2_u0_u4_n100 ) , .A1( u2_u0_u4_n102 ) , .ZN( u2_u0_u4_n144 ) );
  NAND2_X1 u2_u0_u4_U65 (.A2( u2_u0_u4_n101 ) , .A1( u2_u0_u4_n105 ) , .ZN( u2_u0_u4_n96 ) );
  INV_X1 u2_u0_u4_U66 (.A( u2_u0_u4_n128 ) , .ZN( u2_u0_u4_n174 ) );
  NAND2_X1 u2_u0_u4_U67 (.A2( u2_u0_u4_n102 ) , .ZN( u2_u0_u4_n119 ) , .A1( u2_u0_u4_n98 ) );
  NAND2_X1 u2_u0_u4_U68 (.A2( u2_u0_u4_n101 ) , .A1( u2_u0_u4_n103 ) , .ZN( u2_u0_u4_n147 ) );
  NAND2_X1 u2_u0_u4_U69 (.A2( u2_u0_u4_n104 ) , .ZN( u2_u0_u4_n113 ) , .A1( u2_u0_u4_n99 ) );
  AOI21_X1 u2_u0_u4_U7 (.ZN( u2_u0_u4_n108 ) , .B2( u2_u0_u4_n134 ) , .B1( u2_u0_u4_n155 ) , .A( u2_u0_u4_n156 ) );
  NOR2_X1 u2_u0_u4_U70 (.A2( u2_u0_X_28 ) , .ZN( u2_u0_u4_n150 ) , .A1( u2_u0_u4_n168 ) );
  NOR2_X1 u2_u0_u4_U71 (.A2( u2_u0_X_29 ) , .ZN( u2_u0_u4_n152 ) , .A1( u2_u0_u4_n169 ) );
  NOR2_X1 u2_u0_u4_U72 (.A2( u2_u0_X_30 ) , .ZN( u2_u0_u4_n105 ) , .A1( u2_u0_u4_n176 ) );
  NOR2_X1 u2_u0_u4_U73 (.A2( u2_u0_X_26 ) , .ZN( u2_u0_u4_n100 ) , .A1( u2_u0_u4_n177 ) );
  NOR2_X1 u2_u0_u4_U74 (.A2( u2_u0_X_28 ) , .A1( u2_u0_X_29 ) , .ZN( u2_u0_u4_n128 ) );
  NOR2_X1 u2_u0_u4_U75 (.A2( u2_u0_X_27 ) , .A1( u2_u0_X_30 ) , .ZN( u2_u0_u4_n102 ) );
  NOR2_X1 u2_u0_u4_U76 (.A2( u2_u0_X_25 ) , .A1( u2_u0_X_26 ) , .ZN( u2_u0_u4_n98 ) );
  AND2_X1 u2_u0_u4_U77 (.A2( u2_u0_X_25 ) , .A1( u2_u0_X_26 ) , .ZN( u2_u0_u4_n104 ) );
  AND2_X1 u2_u0_u4_U78 (.A1( u2_u0_X_30 ) , .A2( u2_u0_u4_n176 ) , .ZN( u2_u0_u4_n99 ) );
  AND2_X1 u2_u0_u4_U79 (.A1( u2_u0_X_26 ) , .ZN( u2_u0_u4_n101 ) , .A2( u2_u0_u4_n177 ) );
  AOI21_X1 u2_u0_u4_U8 (.ZN( u2_u0_u4_n109 ) , .A( u2_u0_u4_n153 ) , .B1( u2_u0_u4_n159 ) , .B2( u2_u0_u4_n184 ) );
  AND2_X1 u2_u0_u4_U80 (.A1( u2_u0_X_27 ) , .A2( u2_u0_X_30 ) , .ZN( u2_u0_u4_n103 ) );
  INV_X1 u2_u0_u4_U81 (.A( u2_u0_X_28 ) , .ZN( u2_u0_u4_n169 ) );
  INV_X1 u2_u0_u4_U82 (.A( u2_u0_X_29 ) , .ZN( u2_u0_u4_n168 ) );
  INV_X1 u2_u0_u4_U83 (.A( u2_u0_X_25 ) , .ZN( u2_u0_u4_n177 ) );
  INV_X1 u2_u0_u4_U84 (.A( u2_u0_X_27 ) , .ZN( u2_u0_u4_n176 ) );
  NAND4_X1 u2_u0_u4_U85 (.ZN( u2_out0_25 ) , .A4( u2_u0_u4_n139 ) , .A3( u2_u0_u4_n140 ) , .A2( u2_u0_u4_n141 ) , .A1( u2_u0_u4_n142 ) );
  OAI21_X1 u2_u0_u4_U86 (.A( u2_u0_u4_n128 ) , .B2( u2_u0_u4_n129 ) , .B1( u2_u0_u4_n130 ) , .ZN( u2_u0_u4_n142 ) );
  OAI21_X1 u2_u0_u4_U87 (.B2( u2_u0_u4_n131 ) , .ZN( u2_u0_u4_n141 ) , .A( u2_u0_u4_n175 ) , .B1( u2_u0_u4_n183 ) );
  NAND4_X1 u2_u0_u4_U88 (.ZN( u2_out0_14 ) , .A4( u2_u0_u4_n124 ) , .A3( u2_u0_u4_n125 ) , .A2( u2_u0_u4_n126 ) , .A1( u2_u0_u4_n127 ) );
  AOI22_X1 u2_u0_u4_U89 (.B2( u2_u0_u4_n117 ) , .ZN( u2_u0_u4_n126 ) , .A1( u2_u0_u4_n129 ) , .B1( u2_u0_u4_n152 ) , .A2( u2_u0_u4_n175 ) );
  AOI211_X1 u2_u0_u4_U9 (.B( u2_u0_u4_n136 ) , .A( u2_u0_u4_n137 ) , .C2( u2_u0_u4_n138 ) , .ZN( u2_u0_u4_n139 ) , .C1( u2_u0_u4_n182 ) );
  AOI22_X1 u2_u0_u4_U90 (.ZN( u2_u0_u4_n125 ) , .B2( u2_u0_u4_n131 ) , .A2( u2_u0_u4_n132 ) , .B1( u2_u0_u4_n138 ) , .A1( u2_u0_u4_n178 ) );
  NAND4_X1 u2_u0_u4_U91 (.ZN( u2_out0_8 ) , .A4( u2_u0_u4_n110 ) , .A3( u2_u0_u4_n111 ) , .A2( u2_u0_u4_n112 ) , .A1( u2_u0_u4_n186 ) );
  NAND2_X1 u2_u0_u4_U92 (.ZN( u2_u0_u4_n112 ) , .A2( u2_u0_u4_n130 ) , .A1( u2_u0_u4_n150 ) );
  AOI22_X1 u2_u0_u4_U93 (.ZN( u2_u0_u4_n111 ) , .B2( u2_u0_u4_n132 ) , .A1( u2_u0_u4_n152 ) , .B1( u2_u0_u4_n178 ) , .A2( u2_u0_u4_n97 ) );
  AOI22_X1 u2_u0_u4_U94 (.B2( u2_u0_u4_n149 ) , .B1( u2_u0_u4_n150 ) , .A2( u2_u0_u4_n151 ) , .A1( u2_u0_u4_n152 ) , .ZN( u2_u0_u4_n167 ) );
  NOR4_X1 u2_u0_u4_U95 (.A4( u2_u0_u4_n162 ) , .A3( u2_u0_u4_n163 ) , .A2( u2_u0_u4_n164 ) , .A1( u2_u0_u4_n165 ) , .ZN( u2_u0_u4_n166 ) );
  NAND3_X1 u2_u0_u4_U96 (.ZN( u2_out0_3 ) , .A3( u2_u0_u4_n166 ) , .A1( u2_u0_u4_n167 ) , .A2( u2_u0_u4_n186 ) );
  NAND3_X1 u2_u0_u4_U97 (.A3( u2_u0_u4_n146 ) , .A2( u2_u0_u4_n147 ) , .A1( u2_u0_u4_n148 ) , .ZN( u2_u0_u4_n149 ) );
  NAND3_X1 u2_u0_u4_U98 (.A3( u2_u0_u4_n143 ) , .A2( u2_u0_u4_n144 ) , .A1( u2_u0_u4_n145 ) , .ZN( u2_u0_u4_n151 ) );
  NAND3_X1 u2_u0_u4_U99 (.A3( u2_u0_u4_n121 ) , .ZN( u2_u0_u4_n122 ) , .A2( u2_u0_u4_n144 ) , .A1( u2_u0_u4_n154 ) );
  INV_X1 u2_u0_u5_U10 (.A( u2_u0_u5_n121 ) , .ZN( u2_u0_u5_n177 ) );
  NOR3_X1 u2_u0_u5_U100 (.A3( u2_u0_u5_n141 ) , .A1( u2_u0_u5_n142 ) , .ZN( u2_u0_u5_n143 ) , .A2( u2_u0_u5_n191 ) );
  NAND4_X1 u2_u0_u5_U101 (.ZN( u2_out0_4 ) , .A4( u2_u0_u5_n112 ) , .A2( u2_u0_u5_n113 ) , .A1( u2_u0_u5_n114 ) , .A3( u2_u0_u5_n195 ) );
  AOI211_X1 u2_u0_u5_U102 (.A( u2_u0_u5_n110 ) , .C1( u2_u0_u5_n111 ) , .ZN( u2_u0_u5_n112 ) , .B( u2_u0_u5_n118 ) , .C2( u2_u0_u5_n177 ) );
  AOI222_X1 u2_u0_u5_U103 (.ZN( u2_u0_u5_n113 ) , .A1( u2_u0_u5_n131 ) , .C1( u2_u0_u5_n148 ) , .B2( u2_u0_u5_n174 ) , .C2( u2_u0_u5_n178 ) , .A2( u2_u0_u5_n179 ) , .B1( u2_u0_u5_n99 ) );
  NAND3_X1 u2_u0_u5_U104 (.A2( u2_u0_u5_n154 ) , .A3( u2_u0_u5_n158 ) , .A1( u2_u0_u5_n161 ) , .ZN( u2_u0_u5_n99 ) );
  NOR2_X1 u2_u0_u5_U11 (.ZN( u2_u0_u5_n160 ) , .A2( u2_u0_u5_n173 ) , .A1( u2_u0_u5_n177 ) );
  INV_X1 u2_u0_u5_U12 (.A( u2_u0_u5_n150 ) , .ZN( u2_u0_u5_n174 ) );
  AOI21_X1 u2_u0_u5_U13 (.A( u2_u0_u5_n160 ) , .B2( u2_u0_u5_n161 ) , .ZN( u2_u0_u5_n162 ) , .B1( u2_u0_u5_n192 ) );
  INV_X1 u2_u0_u5_U14 (.A( u2_u0_u5_n159 ) , .ZN( u2_u0_u5_n192 ) );
  AOI21_X1 u2_u0_u5_U15 (.A( u2_u0_u5_n156 ) , .B2( u2_u0_u5_n157 ) , .B1( u2_u0_u5_n158 ) , .ZN( u2_u0_u5_n163 ) );
  AOI21_X1 u2_u0_u5_U16 (.B2( u2_u0_u5_n139 ) , .B1( u2_u0_u5_n140 ) , .ZN( u2_u0_u5_n141 ) , .A( u2_u0_u5_n150 ) );
  OAI21_X1 u2_u0_u5_U17 (.A( u2_u0_u5_n133 ) , .B2( u2_u0_u5_n134 ) , .B1( u2_u0_u5_n135 ) , .ZN( u2_u0_u5_n142 ) );
  OAI21_X1 u2_u0_u5_U18 (.ZN( u2_u0_u5_n133 ) , .B2( u2_u0_u5_n147 ) , .A( u2_u0_u5_n173 ) , .B1( u2_u0_u5_n188 ) );
  NAND2_X1 u2_u0_u5_U19 (.A2( u2_u0_u5_n119 ) , .A1( u2_u0_u5_n123 ) , .ZN( u2_u0_u5_n137 ) );
  INV_X1 u2_u0_u5_U20 (.A( u2_u0_u5_n155 ) , .ZN( u2_u0_u5_n194 ) );
  NAND2_X1 u2_u0_u5_U21 (.A1( u2_u0_u5_n121 ) , .ZN( u2_u0_u5_n132 ) , .A2( u2_u0_u5_n172 ) );
  NAND2_X1 u2_u0_u5_U22 (.A2( u2_u0_u5_n122 ) , .ZN( u2_u0_u5_n136 ) , .A1( u2_u0_u5_n154 ) );
  NAND2_X1 u2_u0_u5_U23 (.A2( u2_u0_u5_n119 ) , .A1( u2_u0_u5_n120 ) , .ZN( u2_u0_u5_n159 ) );
  INV_X1 u2_u0_u5_U24 (.A( u2_u0_u5_n156 ) , .ZN( u2_u0_u5_n175 ) );
  INV_X1 u2_u0_u5_U25 (.A( u2_u0_u5_n158 ) , .ZN( u2_u0_u5_n188 ) );
  INV_X1 u2_u0_u5_U26 (.A( u2_u0_u5_n152 ) , .ZN( u2_u0_u5_n179 ) );
  INV_X1 u2_u0_u5_U27 (.A( u2_u0_u5_n140 ) , .ZN( u2_u0_u5_n182 ) );
  INV_X1 u2_u0_u5_U28 (.A( u2_u0_u5_n151 ) , .ZN( u2_u0_u5_n183 ) );
  INV_X1 u2_u0_u5_U29 (.A( u2_u0_u5_n123 ) , .ZN( u2_u0_u5_n185 ) );
  NOR2_X1 u2_u0_u5_U3 (.ZN( u2_u0_u5_n134 ) , .A1( u2_u0_u5_n183 ) , .A2( u2_u0_u5_n190 ) );
  INV_X1 u2_u0_u5_U30 (.A( u2_u0_u5_n161 ) , .ZN( u2_u0_u5_n184 ) );
  INV_X1 u2_u0_u5_U31 (.A( u2_u0_u5_n139 ) , .ZN( u2_u0_u5_n189 ) );
  INV_X1 u2_u0_u5_U32 (.A( u2_u0_u5_n157 ) , .ZN( u2_u0_u5_n190 ) );
  INV_X1 u2_u0_u5_U33 (.A( u2_u0_u5_n120 ) , .ZN( u2_u0_u5_n193 ) );
  NAND2_X1 u2_u0_u5_U34 (.ZN( u2_u0_u5_n111 ) , .A1( u2_u0_u5_n140 ) , .A2( u2_u0_u5_n155 ) );
  NOR2_X1 u2_u0_u5_U35 (.ZN( u2_u0_u5_n100 ) , .A1( u2_u0_u5_n170 ) , .A2( u2_u0_u5_n180 ) );
  INV_X1 u2_u0_u5_U36 (.A( u2_u0_u5_n117 ) , .ZN( u2_u0_u5_n196 ) );
  OAI221_X1 u2_u0_u5_U37 (.A( u2_u0_u5_n116 ) , .ZN( u2_u0_u5_n117 ) , .B2( u2_u0_u5_n119 ) , .C1( u2_u0_u5_n153 ) , .C2( u2_u0_u5_n158 ) , .B1( u2_u0_u5_n172 ) );
  AOI222_X1 u2_u0_u5_U38 (.ZN( u2_u0_u5_n116 ) , .B2( u2_u0_u5_n145 ) , .C1( u2_u0_u5_n148 ) , .A2( u2_u0_u5_n174 ) , .C2( u2_u0_u5_n177 ) , .B1( u2_u0_u5_n187 ) , .A1( u2_u0_u5_n193 ) );
  INV_X1 u2_u0_u5_U39 (.A( u2_u0_u5_n115 ) , .ZN( u2_u0_u5_n187 ) );
  INV_X1 u2_u0_u5_U4 (.A( u2_u0_u5_n138 ) , .ZN( u2_u0_u5_n191 ) );
  AOI22_X1 u2_u0_u5_U40 (.B2( u2_u0_u5_n131 ) , .A2( u2_u0_u5_n146 ) , .ZN( u2_u0_u5_n169 ) , .B1( u2_u0_u5_n174 ) , .A1( u2_u0_u5_n185 ) );
  NOR2_X1 u2_u0_u5_U41 (.A1( u2_u0_u5_n146 ) , .ZN( u2_u0_u5_n150 ) , .A2( u2_u0_u5_n173 ) );
  AOI21_X1 u2_u0_u5_U42 (.A( u2_u0_u5_n118 ) , .B2( u2_u0_u5_n145 ) , .ZN( u2_u0_u5_n168 ) , .B1( u2_u0_u5_n186 ) );
  INV_X1 u2_u0_u5_U43 (.A( u2_u0_u5_n122 ) , .ZN( u2_u0_u5_n186 ) );
  NOR2_X1 u2_u0_u5_U44 (.A1( u2_u0_u5_n146 ) , .ZN( u2_u0_u5_n152 ) , .A2( u2_u0_u5_n176 ) );
  NOR2_X1 u2_u0_u5_U45 (.A1( u2_u0_u5_n115 ) , .ZN( u2_u0_u5_n118 ) , .A2( u2_u0_u5_n153 ) );
  NOR2_X1 u2_u0_u5_U46 (.A2( u2_u0_u5_n145 ) , .ZN( u2_u0_u5_n156 ) , .A1( u2_u0_u5_n174 ) );
  NOR2_X1 u2_u0_u5_U47 (.ZN( u2_u0_u5_n121 ) , .A2( u2_u0_u5_n145 ) , .A1( u2_u0_u5_n176 ) );
  AOI22_X1 u2_u0_u5_U48 (.ZN( u2_u0_u5_n114 ) , .A2( u2_u0_u5_n137 ) , .A1( u2_u0_u5_n145 ) , .B2( u2_u0_u5_n175 ) , .B1( u2_u0_u5_n193 ) );
  OAI211_X1 u2_u0_u5_U49 (.B( u2_u0_u5_n124 ) , .A( u2_u0_u5_n125 ) , .C2( u2_u0_u5_n126 ) , .C1( u2_u0_u5_n127 ) , .ZN( u2_u0_u5_n128 ) );
  OAI21_X1 u2_u0_u5_U5 (.B2( u2_u0_u5_n136 ) , .B1( u2_u0_u5_n137 ) , .ZN( u2_u0_u5_n138 ) , .A( u2_u0_u5_n177 ) );
  NOR3_X1 u2_u0_u5_U50 (.ZN( u2_u0_u5_n127 ) , .A1( u2_u0_u5_n136 ) , .A3( u2_u0_u5_n148 ) , .A2( u2_u0_u5_n182 ) );
  OAI21_X1 u2_u0_u5_U51 (.ZN( u2_u0_u5_n124 ) , .A( u2_u0_u5_n177 ) , .B2( u2_u0_u5_n183 ) , .B1( u2_u0_u5_n189 ) );
  OAI21_X1 u2_u0_u5_U52 (.ZN( u2_u0_u5_n125 ) , .A( u2_u0_u5_n174 ) , .B2( u2_u0_u5_n185 ) , .B1( u2_u0_u5_n190 ) );
  AOI21_X1 u2_u0_u5_U53 (.A( u2_u0_u5_n153 ) , .B2( u2_u0_u5_n154 ) , .B1( u2_u0_u5_n155 ) , .ZN( u2_u0_u5_n164 ) );
  AOI21_X1 u2_u0_u5_U54 (.ZN( u2_u0_u5_n110 ) , .B1( u2_u0_u5_n122 ) , .B2( u2_u0_u5_n139 ) , .A( u2_u0_u5_n153 ) );
  INV_X1 u2_u0_u5_U55 (.A( u2_u0_u5_n153 ) , .ZN( u2_u0_u5_n176 ) );
  INV_X1 u2_u0_u5_U56 (.A( u2_u0_u5_n126 ) , .ZN( u2_u0_u5_n173 ) );
  AND2_X1 u2_u0_u5_U57 (.A2( u2_u0_u5_n104 ) , .A1( u2_u0_u5_n107 ) , .ZN( u2_u0_u5_n147 ) );
  AND2_X1 u2_u0_u5_U58 (.A2( u2_u0_u5_n104 ) , .A1( u2_u0_u5_n108 ) , .ZN( u2_u0_u5_n148 ) );
  NAND2_X1 u2_u0_u5_U59 (.A1( u2_u0_u5_n105 ) , .A2( u2_u0_u5_n106 ) , .ZN( u2_u0_u5_n158 ) );
  INV_X1 u2_u0_u5_U6 (.A( u2_u0_u5_n135 ) , .ZN( u2_u0_u5_n178 ) );
  NAND2_X1 u2_u0_u5_U60 (.A2( u2_u0_u5_n108 ) , .A1( u2_u0_u5_n109 ) , .ZN( u2_u0_u5_n139 ) );
  NAND2_X1 u2_u0_u5_U61 (.A1( u2_u0_u5_n106 ) , .A2( u2_u0_u5_n108 ) , .ZN( u2_u0_u5_n119 ) );
  NAND2_X1 u2_u0_u5_U62 (.A2( u2_u0_u5_n103 ) , .A1( u2_u0_u5_n105 ) , .ZN( u2_u0_u5_n140 ) );
  NAND2_X1 u2_u0_u5_U63 (.A2( u2_u0_u5_n104 ) , .A1( u2_u0_u5_n105 ) , .ZN( u2_u0_u5_n155 ) );
  NAND2_X1 u2_u0_u5_U64 (.A2( u2_u0_u5_n106 ) , .A1( u2_u0_u5_n107 ) , .ZN( u2_u0_u5_n122 ) );
  NAND2_X1 u2_u0_u5_U65 (.A2( u2_u0_u5_n100 ) , .A1( u2_u0_u5_n106 ) , .ZN( u2_u0_u5_n115 ) );
  NAND2_X1 u2_u0_u5_U66 (.A2( u2_u0_u5_n100 ) , .A1( u2_u0_u5_n103 ) , .ZN( u2_u0_u5_n161 ) );
  NAND2_X1 u2_u0_u5_U67 (.A1( u2_u0_u5_n105 ) , .A2( u2_u0_u5_n109 ) , .ZN( u2_u0_u5_n154 ) );
  INV_X1 u2_u0_u5_U68 (.A( u2_u0_u5_n146 ) , .ZN( u2_u0_u5_n172 ) );
  NAND2_X1 u2_u0_u5_U69 (.A1( u2_u0_u5_n103 ) , .A2( u2_u0_u5_n108 ) , .ZN( u2_u0_u5_n123 ) );
  OAI22_X1 u2_u0_u5_U7 (.B2( u2_u0_u5_n149 ) , .B1( u2_u0_u5_n150 ) , .A2( u2_u0_u5_n151 ) , .A1( u2_u0_u5_n152 ) , .ZN( u2_u0_u5_n165 ) );
  NAND2_X1 u2_u0_u5_U70 (.A2( u2_u0_u5_n103 ) , .A1( u2_u0_u5_n107 ) , .ZN( u2_u0_u5_n151 ) );
  NAND2_X1 u2_u0_u5_U71 (.A2( u2_u0_u5_n107 ) , .A1( u2_u0_u5_n109 ) , .ZN( u2_u0_u5_n120 ) );
  NAND2_X1 u2_u0_u5_U72 (.A2( u2_u0_u5_n100 ) , .A1( u2_u0_u5_n109 ) , .ZN( u2_u0_u5_n157 ) );
  AND2_X1 u2_u0_u5_U73 (.A2( u2_u0_u5_n100 ) , .A1( u2_u0_u5_n104 ) , .ZN( u2_u0_u5_n131 ) );
  INV_X1 u2_u0_u5_U74 (.A( u2_u0_u5_n102 ) , .ZN( u2_u0_u5_n195 ) );
  OAI221_X1 u2_u0_u5_U75 (.A( u2_u0_u5_n101 ) , .ZN( u2_u0_u5_n102 ) , .C2( u2_u0_u5_n115 ) , .C1( u2_u0_u5_n126 ) , .B1( u2_u0_u5_n134 ) , .B2( u2_u0_u5_n160 ) );
  OAI21_X1 u2_u0_u5_U76 (.ZN( u2_u0_u5_n101 ) , .B1( u2_u0_u5_n137 ) , .A( u2_u0_u5_n146 ) , .B2( u2_u0_u5_n147 ) );
  NOR2_X1 u2_u0_u5_U77 (.A2( u2_u0_X_34 ) , .A1( u2_u0_X_35 ) , .ZN( u2_u0_u5_n145 ) );
  NOR2_X1 u2_u0_u5_U78 (.A2( u2_u0_X_34 ) , .ZN( u2_u0_u5_n146 ) , .A1( u2_u0_u5_n171 ) );
  NOR2_X1 u2_u0_u5_U79 (.A2( u2_u0_X_31 ) , .A1( u2_u0_X_32 ) , .ZN( u2_u0_u5_n103 ) );
  NOR3_X1 u2_u0_u5_U8 (.A2( u2_u0_u5_n147 ) , .A1( u2_u0_u5_n148 ) , .ZN( u2_u0_u5_n149 ) , .A3( u2_u0_u5_n194 ) );
  NOR2_X1 u2_u0_u5_U80 (.A2( u2_u0_X_36 ) , .ZN( u2_u0_u5_n105 ) , .A1( u2_u0_u5_n180 ) );
  NOR2_X1 u2_u0_u5_U81 (.A2( u2_u0_X_33 ) , .ZN( u2_u0_u5_n108 ) , .A1( u2_u0_u5_n170 ) );
  NOR2_X1 u2_u0_u5_U82 (.A2( u2_u0_X_33 ) , .A1( u2_u0_X_36 ) , .ZN( u2_u0_u5_n107 ) );
  NOR2_X1 u2_u0_u5_U83 (.A2( u2_u0_X_31 ) , .ZN( u2_u0_u5_n104 ) , .A1( u2_u0_u5_n181 ) );
  NAND2_X1 u2_u0_u5_U84 (.A2( u2_u0_X_34 ) , .A1( u2_u0_X_35 ) , .ZN( u2_u0_u5_n153 ) );
  NAND2_X1 u2_u0_u5_U85 (.A1( u2_u0_X_34 ) , .ZN( u2_u0_u5_n126 ) , .A2( u2_u0_u5_n171 ) );
  AND2_X1 u2_u0_u5_U86 (.A1( u2_u0_X_31 ) , .A2( u2_u0_X_32 ) , .ZN( u2_u0_u5_n106 ) );
  AND2_X1 u2_u0_u5_U87 (.A1( u2_u0_X_31 ) , .ZN( u2_u0_u5_n109 ) , .A2( u2_u0_u5_n181 ) );
  INV_X1 u2_u0_u5_U88 (.A( u2_u0_X_33 ) , .ZN( u2_u0_u5_n180 ) );
  INV_X1 u2_u0_u5_U89 (.A( u2_u0_X_35 ) , .ZN( u2_u0_u5_n171 ) );
  NOR2_X1 u2_u0_u5_U9 (.ZN( u2_u0_u5_n135 ) , .A1( u2_u0_u5_n173 ) , .A2( u2_u0_u5_n176 ) );
  INV_X1 u2_u0_u5_U90 (.A( u2_u0_X_36 ) , .ZN( u2_u0_u5_n170 ) );
  INV_X1 u2_u0_u5_U91 (.A( u2_u0_X_32 ) , .ZN( u2_u0_u5_n181 ) );
  NAND4_X1 u2_u0_u5_U92 (.ZN( u2_out0_29 ) , .A4( u2_u0_u5_n129 ) , .A3( u2_u0_u5_n130 ) , .A2( u2_u0_u5_n168 ) , .A1( u2_u0_u5_n196 ) );
  AOI221_X1 u2_u0_u5_U93 (.A( u2_u0_u5_n128 ) , .ZN( u2_u0_u5_n129 ) , .C2( u2_u0_u5_n132 ) , .B2( u2_u0_u5_n159 ) , .B1( u2_u0_u5_n176 ) , .C1( u2_u0_u5_n184 ) );
  AOI222_X1 u2_u0_u5_U94 (.ZN( u2_u0_u5_n130 ) , .A2( u2_u0_u5_n146 ) , .B1( u2_u0_u5_n147 ) , .C2( u2_u0_u5_n175 ) , .B2( u2_u0_u5_n179 ) , .A1( u2_u0_u5_n188 ) , .C1( u2_u0_u5_n194 ) );
  NAND4_X1 u2_u0_u5_U95 (.ZN( u2_out0_19 ) , .A4( u2_u0_u5_n166 ) , .A3( u2_u0_u5_n167 ) , .A2( u2_u0_u5_n168 ) , .A1( u2_u0_u5_n169 ) );
  AOI22_X1 u2_u0_u5_U96 (.B2( u2_u0_u5_n145 ) , .A2( u2_u0_u5_n146 ) , .ZN( u2_u0_u5_n167 ) , .B1( u2_u0_u5_n182 ) , .A1( u2_u0_u5_n189 ) );
  NOR4_X1 u2_u0_u5_U97 (.A4( u2_u0_u5_n162 ) , .A3( u2_u0_u5_n163 ) , .A2( u2_u0_u5_n164 ) , .A1( u2_u0_u5_n165 ) , .ZN( u2_u0_u5_n166 ) );
  NAND4_X1 u2_u0_u5_U98 (.ZN( u2_out0_11 ) , .A4( u2_u0_u5_n143 ) , .A3( u2_u0_u5_n144 ) , .A2( u2_u0_u5_n169 ) , .A1( u2_u0_u5_n196 ) );
  AOI22_X1 u2_u0_u5_U99 (.A2( u2_u0_u5_n132 ) , .ZN( u2_u0_u5_n144 ) , .B2( u2_u0_u5_n145 ) , .B1( u2_u0_u5_n184 ) , .A1( u2_u0_u5_n194 ) );
  AOI22_X1 u2_u0_u6_U10 (.A2( u2_u0_u6_n151 ) , .B2( u2_u0_u6_n161 ) , .A1( u2_u0_u6_n167 ) , .B1( u2_u0_u6_n170 ) , .ZN( u2_u0_u6_n89 ) );
  AOI21_X1 u2_u0_u6_U11 (.B1( u2_u0_u6_n107 ) , .B2( u2_u0_u6_n132 ) , .A( u2_u0_u6_n158 ) , .ZN( u2_u0_u6_n88 ) );
  AOI21_X1 u2_u0_u6_U12 (.B2( u2_u0_u6_n147 ) , .B1( u2_u0_u6_n148 ) , .ZN( u2_u0_u6_n149 ) , .A( u2_u0_u6_n158 ) );
  AOI21_X1 u2_u0_u6_U13 (.ZN( u2_u0_u6_n106 ) , .A( u2_u0_u6_n142 ) , .B2( u2_u0_u6_n159 ) , .B1( u2_u0_u6_n164 ) );
  INV_X1 u2_u0_u6_U14 (.A( u2_u0_u6_n155 ) , .ZN( u2_u0_u6_n161 ) );
  INV_X1 u2_u0_u6_U15 (.A( u2_u0_u6_n128 ) , .ZN( u2_u0_u6_n164 ) );
  NAND2_X1 u2_u0_u6_U16 (.ZN( u2_u0_u6_n110 ) , .A1( u2_u0_u6_n122 ) , .A2( u2_u0_u6_n129 ) );
  NAND2_X1 u2_u0_u6_U17 (.ZN( u2_u0_u6_n124 ) , .A2( u2_u0_u6_n146 ) , .A1( u2_u0_u6_n148 ) );
  INV_X1 u2_u0_u6_U18 (.A( u2_u0_u6_n132 ) , .ZN( u2_u0_u6_n171 ) );
  AND2_X1 u2_u0_u6_U19 (.A1( u2_u0_u6_n100 ) , .ZN( u2_u0_u6_n130 ) , .A2( u2_u0_u6_n147 ) );
  INV_X1 u2_u0_u6_U20 (.A( u2_u0_u6_n127 ) , .ZN( u2_u0_u6_n173 ) );
  INV_X1 u2_u0_u6_U21 (.A( u2_u0_u6_n121 ) , .ZN( u2_u0_u6_n167 ) );
  INV_X1 u2_u0_u6_U22 (.A( u2_u0_u6_n100 ) , .ZN( u2_u0_u6_n169 ) );
  INV_X1 u2_u0_u6_U23 (.A( u2_u0_u6_n123 ) , .ZN( u2_u0_u6_n170 ) );
  INV_X1 u2_u0_u6_U24 (.A( u2_u0_u6_n113 ) , .ZN( u2_u0_u6_n168 ) );
  AND2_X1 u2_u0_u6_U25 (.A1( u2_u0_u6_n107 ) , .A2( u2_u0_u6_n119 ) , .ZN( u2_u0_u6_n133 ) );
  AND2_X1 u2_u0_u6_U26 (.A2( u2_u0_u6_n121 ) , .A1( u2_u0_u6_n122 ) , .ZN( u2_u0_u6_n131 ) );
  AND3_X1 u2_u0_u6_U27 (.ZN( u2_u0_u6_n120 ) , .A2( u2_u0_u6_n127 ) , .A1( u2_u0_u6_n132 ) , .A3( u2_u0_u6_n145 ) );
  INV_X1 u2_u0_u6_U28 (.A( u2_u0_u6_n146 ) , .ZN( u2_u0_u6_n163 ) );
  AOI222_X1 u2_u0_u6_U29 (.ZN( u2_u0_u6_n114 ) , .A1( u2_u0_u6_n118 ) , .A2( u2_u0_u6_n126 ) , .B2( u2_u0_u6_n151 ) , .C2( u2_u0_u6_n159 ) , .C1( u2_u0_u6_n168 ) , .B1( u2_u0_u6_n169 ) );
  INV_X1 u2_u0_u6_U3 (.A( u2_u0_u6_n110 ) , .ZN( u2_u0_u6_n166 ) );
  NOR2_X1 u2_u0_u6_U30 (.A1( u2_u0_u6_n162 ) , .A2( u2_u0_u6_n165 ) , .ZN( u2_u0_u6_n98 ) );
  AOI211_X1 u2_u0_u6_U31 (.B( u2_u0_u6_n134 ) , .A( u2_u0_u6_n135 ) , .C1( u2_u0_u6_n136 ) , .ZN( u2_u0_u6_n137 ) , .C2( u2_u0_u6_n151 ) );
  AOI21_X1 u2_u0_u6_U32 (.B2( u2_u0_u6_n132 ) , .B1( u2_u0_u6_n133 ) , .ZN( u2_u0_u6_n134 ) , .A( u2_u0_u6_n158 ) );
  NAND4_X1 u2_u0_u6_U33 (.A4( u2_u0_u6_n127 ) , .A3( u2_u0_u6_n128 ) , .A2( u2_u0_u6_n129 ) , .A1( u2_u0_u6_n130 ) , .ZN( u2_u0_u6_n136 ) );
  AOI21_X1 u2_u0_u6_U34 (.B1( u2_u0_u6_n131 ) , .ZN( u2_u0_u6_n135 ) , .A( u2_u0_u6_n144 ) , .B2( u2_u0_u6_n146 ) );
  NAND2_X1 u2_u0_u6_U35 (.A1( u2_u0_u6_n144 ) , .ZN( u2_u0_u6_n151 ) , .A2( u2_u0_u6_n158 ) );
  NAND2_X1 u2_u0_u6_U36 (.ZN( u2_u0_u6_n132 ) , .A1( u2_u0_u6_n91 ) , .A2( u2_u0_u6_n97 ) );
  AOI22_X1 u2_u0_u6_U37 (.B2( u2_u0_u6_n110 ) , .B1( u2_u0_u6_n111 ) , .A1( u2_u0_u6_n112 ) , .ZN( u2_u0_u6_n115 ) , .A2( u2_u0_u6_n161 ) );
  NAND4_X1 u2_u0_u6_U38 (.A3( u2_u0_u6_n109 ) , .ZN( u2_u0_u6_n112 ) , .A4( u2_u0_u6_n132 ) , .A2( u2_u0_u6_n147 ) , .A1( u2_u0_u6_n166 ) );
  NOR2_X1 u2_u0_u6_U39 (.ZN( u2_u0_u6_n109 ) , .A1( u2_u0_u6_n170 ) , .A2( u2_u0_u6_n173 ) );
  INV_X1 u2_u0_u6_U4 (.A( u2_u0_u6_n142 ) , .ZN( u2_u0_u6_n174 ) );
  NOR2_X1 u2_u0_u6_U40 (.A2( u2_u0_u6_n126 ) , .ZN( u2_u0_u6_n155 ) , .A1( u2_u0_u6_n160 ) );
  NAND2_X1 u2_u0_u6_U41 (.ZN( u2_u0_u6_n146 ) , .A2( u2_u0_u6_n94 ) , .A1( u2_u0_u6_n99 ) );
  AOI21_X1 u2_u0_u6_U42 (.A( u2_u0_u6_n144 ) , .B2( u2_u0_u6_n145 ) , .B1( u2_u0_u6_n146 ) , .ZN( u2_u0_u6_n150 ) );
  INV_X1 u2_u0_u6_U43 (.A( u2_u0_u6_n111 ) , .ZN( u2_u0_u6_n158 ) );
  NAND2_X1 u2_u0_u6_U44 (.ZN( u2_u0_u6_n127 ) , .A1( u2_u0_u6_n91 ) , .A2( u2_u0_u6_n92 ) );
  NAND2_X1 u2_u0_u6_U45 (.ZN( u2_u0_u6_n129 ) , .A2( u2_u0_u6_n95 ) , .A1( u2_u0_u6_n96 ) );
  INV_X1 u2_u0_u6_U46 (.A( u2_u0_u6_n144 ) , .ZN( u2_u0_u6_n159 ) );
  NAND2_X1 u2_u0_u6_U47 (.ZN( u2_u0_u6_n145 ) , .A2( u2_u0_u6_n97 ) , .A1( u2_u0_u6_n98 ) );
  NAND2_X1 u2_u0_u6_U48 (.ZN( u2_u0_u6_n148 ) , .A2( u2_u0_u6_n92 ) , .A1( u2_u0_u6_n94 ) );
  NAND2_X1 u2_u0_u6_U49 (.ZN( u2_u0_u6_n108 ) , .A2( u2_u0_u6_n139 ) , .A1( u2_u0_u6_n144 ) );
  NAND2_X1 u2_u0_u6_U5 (.A2( u2_u0_u6_n143 ) , .ZN( u2_u0_u6_n152 ) , .A1( u2_u0_u6_n166 ) );
  NAND2_X1 u2_u0_u6_U50 (.ZN( u2_u0_u6_n121 ) , .A2( u2_u0_u6_n95 ) , .A1( u2_u0_u6_n97 ) );
  NAND2_X1 u2_u0_u6_U51 (.ZN( u2_u0_u6_n107 ) , .A2( u2_u0_u6_n92 ) , .A1( u2_u0_u6_n95 ) );
  AND2_X1 u2_u0_u6_U52 (.ZN( u2_u0_u6_n118 ) , .A2( u2_u0_u6_n91 ) , .A1( u2_u0_u6_n99 ) );
  NAND2_X1 u2_u0_u6_U53 (.ZN( u2_u0_u6_n147 ) , .A2( u2_u0_u6_n98 ) , .A1( u2_u0_u6_n99 ) );
  NAND2_X1 u2_u0_u6_U54 (.ZN( u2_u0_u6_n128 ) , .A1( u2_u0_u6_n94 ) , .A2( u2_u0_u6_n96 ) );
  NAND2_X1 u2_u0_u6_U55 (.ZN( u2_u0_u6_n119 ) , .A2( u2_u0_u6_n95 ) , .A1( u2_u0_u6_n99 ) );
  NAND2_X1 u2_u0_u6_U56 (.ZN( u2_u0_u6_n123 ) , .A2( u2_u0_u6_n91 ) , .A1( u2_u0_u6_n96 ) );
  NAND2_X1 u2_u0_u6_U57 (.ZN( u2_u0_u6_n100 ) , .A2( u2_u0_u6_n92 ) , .A1( u2_u0_u6_n98 ) );
  NAND2_X1 u2_u0_u6_U58 (.ZN( u2_u0_u6_n122 ) , .A1( u2_u0_u6_n94 ) , .A2( u2_u0_u6_n97 ) );
  INV_X1 u2_u0_u6_U59 (.A( u2_u0_u6_n139 ) , .ZN( u2_u0_u6_n160 ) );
  AOI22_X1 u2_u0_u6_U6 (.B2( u2_u0_u6_n101 ) , .A1( u2_u0_u6_n102 ) , .ZN( u2_u0_u6_n103 ) , .B1( u2_u0_u6_n160 ) , .A2( u2_u0_u6_n161 ) );
  NAND2_X1 u2_u0_u6_U60 (.ZN( u2_u0_u6_n113 ) , .A1( u2_u0_u6_n96 ) , .A2( u2_u0_u6_n98 ) );
  NOR2_X1 u2_u0_u6_U61 (.A2( u2_u0_X_40 ) , .A1( u2_u0_X_41 ) , .ZN( u2_u0_u6_n126 ) );
  NOR2_X1 u2_u0_u6_U62 (.A2( u2_u0_X_39 ) , .A1( u2_u0_X_42 ) , .ZN( u2_u0_u6_n92 ) );
  NOR2_X1 u2_u0_u6_U63 (.A2( u2_u0_X_39 ) , .A1( u2_u0_u6_n156 ) , .ZN( u2_u0_u6_n97 ) );
  NOR2_X1 u2_u0_u6_U64 (.A2( u2_u0_X_38 ) , .A1( u2_u0_u6_n165 ) , .ZN( u2_u0_u6_n95 ) );
  NOR2_X1 u2_u0_u6_U65 (.A2( u2_u0_X_41 ) , .ZN( u2_u0_u6_n111 ) , .A1( u2_u0_u6_n157 ) );
  NOR2_X1 u2_u0_u6_U66 (.A2( u2_u0_X_37 ) , .A1( u2_u0_u6_n162 ) , .ZN( u2_u0_u6_n94 ) );
  NOR2_X1 u2_u0_u6_U67 (.A2( u2_u0_X_37 ) , .A1( u2_u0_X_38 ) , .ZN( u2_u0_u6_n91 ) );
  NAND2_X1 u2_u0_u6_U68 (.A1( u2_u0_X_41 ) , .ZN( u2_u0_u6_n144 ) , .A2( u2_u0_u6_n157 ) );
  NAND2_X1 u2_u0_u6_U69 (.A2( u2_u0_X_40 ) , .A1( u2_u0_X_41 ) , .ZN( u2_u0_u6_n139 ) );
  NOR2_X1 u2_u0_u6_U7 (.A1( u2_u0_u6_n118 ) , .ZN( u2_u0_u6_n143 ) , .A2( u2_u0_u6_n168 ) );
  AND2_X1 u2_u0_u6_U70 (.A1( u2_u0_X_39 ) , .A2( u2_u0_u6_n156 ) , .ZN( u2_u0_u6_n96 ) );
  AND2_X1 u2_u0_u6_U71 (.A1( u2_u0_X_39 ) , .A2( u2_u0_X_42 ) , .ZN( u2_u0_u6_n99 ) );
  INV_X1 u2_u0_u6_U72 (.A( u2_u0_X_40 ) , .ZN( u2_u0_u6_n157 ) );
  INV_X1 u2_u0_u6_U73 (.A( u2_u0_X_37 ) , .ZN( u2_u0_u6_n165 ) );
  INV_X1 u2_u0_u6_U74 (.A( u2_u0_X_38 ) , .ZN( u2_u0_u6_n162 ) );
  INV_X1 u2_u0_u6_U75 (.A( u2_u0_X_42 ) , .ZN( u2_u0_u6_n156 ) );
  NAND4_X1 u2_u0_u6_U76 (.ZN( u2_out0_32 ) , .A4( u2_u0_u6_n103 ) , .A3( u2_u0_u6_n104 ) , .A2( u2_u0_u6_n105 ) , .A1( u2_u0_u6_n106 ) );
  AOI22_X1 u2_u0_u6_U77 (.ZN( u2_u0_u6_n105 ) , .A2( u2_u0_u6_n108 ) , .A1( u2_u0_u6_n118 ) , .B2( u2_u0_u6_n126 ) , .B1( u2_u0_u6_n171 ) );
  AOI22_X1 u2_u0_u6_U78 (.ZN( u2_u0_u6_n104 ) , .A1( u2_u0_u6_n111 ) , .B1( u2_u0_u6_n124 ) , .B2( u2_u0_u6_n151 ) , .A2( u2_u0_u6_n93 ) );
  NAND4_X1 u2_u0_u6_U79 (.ZN( u2_out0_12 ) , .A4( u2_u0_u6_n114 ) , .A3( u2_u0_u6_n115 ) , .A2( u2_u0_u6_n116 ) , .A1( u2_u0_u6_n117 ) );
  OAI21_X1 u2_u0_u6_U8 (.A( u2_u0_u6_n159 ) , .B1( u2_u0_u6_n169 ) , .B2( u2_u0_u6_n173 ) , .ZN( u2_u0_u6_n90 ) );
  OAI22_X1 u2_u0_u6_U80 (.B2( u2_u0_u6_n111 ) , .ZN( u2_u0_u6_n116 ) , .B1( u2_u0_u6_n126 ) , .A2( u2_u0_u6_n164 ) , .A1( u2_u0_u6_n167 ) );
  OAI21_X1 u2_u0_u6_U81 (.A( u2_u0_u6_n108 ) , .ZN( u2_u0_u6_n117 ) , .B2( u2_u0_u6_n141 ) , .B1( u2_u0_u6_n163 ) );
  OAI211_X1 u2_u0_u6_U82 (.ZN( u2_out0_7 ) , .B( u2_u0_u6_n153 ) , .C2( u2_u0_u6_n154 ) , .C1( u2_u0_u6_n155 ) , .A( u2_u0_u6_n174 ) );
  NOR3_X1 u2_u0_u6_U83 (.A1( u2_u0_u6_n141 ) , .ZN( u2_u0_u6_n154 ) , .A3( u2_u0_u6_n164 ) , .A2( u2_u0_u6_n171 ) );
  AOI211_X1 u2_u0_u6_U84 (.B( u2_u0_u6_n149 ) , .A( u2_u0_u6_n150 ) , .C2( u2_u0_u6_n151 ) , .C1( u2_u0_u6_n152 ) , .ZN( u2_u0_u6_n153 ) );
  OAI211_X1 u2_u0_u6_U85 (.ZN( u2_out0_22 ) , .B( u2_u0_u6_n137 ) , .A( u2_u0_u6_n138 ) , .C2( u2_u0_u6_n139 ) , .C1( u2_u0_u6_n140 ) );
  AOI22_X1 u2_u0_u6_U86 (.B1( u2_u0_u6_n124 ) , .A2( u2_u0_u6_n125 ) , .A1( u2_u0_u6_n126 ) , .ZN( u2_u0_u6_n138 ) , .B2( u2_u0_u6_n161 ) );
  AND4_X1 u2_u0_u6_U87 (.A3( u2_u0_u6_n119 ) , .A1( u2_u0_u6_n120 ) , .A4( u2_u0_u6_n129 ) , .ZN( u2_u0_u6_n140 ) , .A2( u2_u0_u6_n143 ) );
  NAND3_X1 u2_u0_u6_U88 (.A2( u2_u0_u6_n123 ) , .ZN( u2_u0_u6_n125 ) , .A1( u2_u0_u6_n130 ) , .A3( u2_u0_u6_n131 ) );
  NAND3_X1 u2_u0_u6_U89 (.A3( u2_u0_u6_n133 ) , .ZN( u2_u0_u6_n141 ) , .A1( u2_u0_u6_n145 ) , .A2( u2_u0_u6_n148 ) );
  INV_X1 u2_u0_u6_U9 (.ZN( u2_u0_u6_n172 ) , .A( u2_u0_u6_n88 ) );
  NAND3_X1 u2_u0_u6_U90 (.ZN( u2_u0_u6_n101 ) , .A3( u2_u0_u6_n107 ) , .A2( u2_u0_u6_n121 ) , .A1( u2_u0_u6_n127 ) );
  NAND3_X1 u2_u0_u6_U91 (.ZN( u2_u0_u6_n102 ) , .A3( u2_u0_u6_n130 ) , .A2( u2_u0_u6_n145 ) , .A1( u2_u0_u6_n166 ) );
  NAND3_X1 u2_u0_u6_U92 (.A3( u2_u0_u6_n113 ) , .A1( u2_u0_u6_n119 ) , .A2( u2_u0_u6_n123 ) , .ZN( u2_u0_u6_n93 ) );
  NAND3_X1 u2_u0_u6_U93 (.ZN( u2_u0_u6_n142 ) , .A2( u2_u0_u6_n172 ) , .A3( u2_u0_u6_n89 ) , .A1( u2_u0_u6_n90 ) );
  INV_X1 u2_u0_u7_U10 (.A( u2_u0_u7_n133 ) , .ZN( u2_u0_u7_n176 ) );
  OAI221_X1 u2_u0_u7_U11 (.C1( u2_u0_u7_n101 ) , .C2( u2_u0_u7_n147 ) , .ZN( u2_u0_u7_n155 ) , .B2( u2_u0_u7_n162 ) , .A( u2_u0_u7_n91 ) , .B1( u2_u0_u7_n92 ) );
  AND3_X1 u2_u0_u7_U12 (.A3( u2_u0_u7_n110 ) , .A2( u2_u0_u7_n127 ) , .A1( u2_u0_u7_n132 ) , .ZN( u2_u0_u7_n92 ) );
  OAI21_X1 u2_u0_u7_U13 (.A( u2_u0_u7_n161 ) , .B1( u2_u0_u7_n168 ) , .B2( u2_u0_u7_n173 ) , .ZN( u2_u0_u7_n91 ) );
  AOI211_X1 u2_u0_u7_U14 (.A( u2_u0_u7_n117 ) , .ZN( u2_u0_u7_n118 ) , .C2( u2_u0_u7_n126 ) , .C1( u2_u0_u7_n177 ) , .B( u2_u0_u7_n180 ) );
  OAI22_X1 u2_u0_u7_U15 (.B1( u2_u0_u7_n115 ) , .ZN( u2_u0_u7_n117 ) , .A2( u2_u0_u7_n133 ) , .A1( u2_u0_u7_n137 ) , .B2( u2_u0_u7_n162 ) );
  INV_X1 u2_u0_u7_U16 (.A( u2_u0_u7_n116 ) , .ZN( u2_u0_u7_n180 ) );
  NOR3_X1 u2_u0_u7_U17 (.ZN( u2_u0_u7_n115 ) , .A3( u2_u0_u7_n145 ) , .A2( u2_u0_u7_n168 ) , .A1( u2_u0_u7_n169 ) );
  NOR3_X1 u2_u0_u7_U18 (.A2( u2_u0_u7_n134 ) , .A1( u2_u0_u7_n135 ) , .ZN( u2_u0_u7_n136 ) , .A3( u2_u0_u7_n171 ) );
  NOR2_X1 u2_u0_u7_U19 (.A1( u2_u0_u7_n130 ) , .A2( u2_u0_u7_n134 ) , .ZN( u2_u0_u7_n153 ) );
  INV_X1 u2_u0_u7_U20 (.A( u2_u0_u7_n101 ) , .ZN( u2_u0_u7_n165 ) );
  NOR2_X1 u2_u0_u7_U21 (.ZN( u2_u0_u7_n111 ) , .A2( u2_u0_u7_n134 ) , .A1( u2_u0_u7_n169 ) );
  AOI21_X1 u2_u0_u7_U22 (.ZN( u2_u0_u7_n104 ) , .B2( u2_u0_u7_n112 ) , .B1( u2_u0_u7_n127 ) , .A( u2_u0_u7_n164 ) );
  AOI21_X1 u2_u0_u7_U23 (.ZN( u2_u0_u7_n106 ) , .B1( u2_u0_u7_n133 ) , .B2( u2_u0_u7_n146 ) , .A( u2_u0_u7_n162 ) );
  AOI21_X1 u2_u0_u7_U24 (.A( u2_u0_u7_n101 ) , .ZN( u2_u0_u7_n107 ) , .B2( u2_u0_u7_n128 ) , .B1( u2_u0_u7_n175 ) );
  INV_X1 u2_u0_u7_U25 (.A( u2_u0_u7_n138 ) , .ZN( u2_u0_u7_n171 ) );
  INV_X1 u2_u0_u7_U26 (.A( u2_u0_u7_n131 ) , .ZN( u2_u0_u7_n177 ) );
  INV_X1 u2_u0_u7_U27 (.A( u2_u0_u7_n110 ) , .ZN( u2_u0_u7_n174 ) );
  NAND2_X1 u2_u0_u7_U28 (.A1( u2_u0_u7_n129 ) , .A2( u2_u0_u7_n132 ) , .ZN( u2_u0_u7_n149 ) );
  NAND2_X1 u2_u0_u7_U29 (.A1( u2_u0_u7_n113 ) , .A2( u2_u0_u7_n124 ) , .ZN( u2_u0_u7_n130 ) );
  OAI21_X1 u2_u0_u7_U3 (.ZN( u2_u0_u7_n159 ) , .A( u2_u0_u7_n165 ) , .B2( u2_u0_u7_n171 ) , .B1( u2_u0_u7_n174 ) );
  INV_X1 u2_u0_u7_U30 (.A( u2_u0_u7_n112 ) , .ZN( u2_u0_u7_n173 ) );
  INV_X1 u2_u0_u7_U31 (.A( u2_u0_u7_n128 ) , .ZN( u2_u0_u7_n168 ) );
  INV_X1 u2_u0_u7_U32 (.A( u2_u0_u7_n148 ) , .ZN( u2_u0_u7_n169 ) );
  INV_X1 u2_u0_u7_U33 (.A( u2_u0_u7_n127 ) , .ZN( u2_u0_u7_n179 ) );
  NOR2_X1 u2_u0_u7_U34 (.ZN( u2_u0_u7_n101 ) , .A2( u2_u0_u7_n150 ) , .A1( u2_u0_u7_n156 ) );
  AOI211_X1 u2_u0_u7_U35 (.B( u2_u0_u7_n139 ) , .A( u2_u0_u7_n140 ) , .C2( u2_u0_u7_n141 ) , .ZN( u2_u0_u7_n142 ) , .C1( u2_u0_u7_n156 ) );
  NAND4_X1 u2_u0_u7_U36 (.A3( u2_u0_u7_n127 ) , .A2( u2_u0_u7_n128 ) , .A1( u2_u0_u7_n129 ) , .ZN( u2_u0_u7_n141 ) , .A4( u2_u0_u7_n147 ) );
  AOI21_X1 u2_u0_u7_U37 (.A( u2_u0_u7_n137 ) , .B1( u2_u0_u7_n138 ) , .ZN( u2_u0_u7_n139 ) , .B2( u2_u0_u7_n146 ) );
  OAI22_X1 u2_u0_u7_U38 (.B1( u2_u0_u7_n136 ) , .ZN( u2_u0_u7_n140 ) , .A1( u2_u0_u7_n153 ) , .B2( u2_u0_u7_n162 ) , .A2( u2_u0_u7_n164 ) );
  AOI211_X1 u2_u0_u7_U39 (.B( u2_u0_u7_n154 ) , .A( u2_u0_u7_n155 ) , .C1( u2_u0_u7_n156 ) , .ZN( u2_u0_u7_n157 ) , .C2( u2_u0_u7_n172 ) );
  INV_X1 u2_u0_u7_U4 (.A( u2_u0_u7_n111 ) , .ZN( u2_u0_u7_n170 ) );
  INV_X1 u2_u0_u7_U40 (.A( u2_u0_u7_n153 ) , .ZN( u2_u0_u7_n172 ) );
  INV_X1 u2_u0_u7_U41 (.A( u2_u0_u7_n125 ) , .ZN( u2_u0_u7_n161 ) );
  NAND2_X1 u2_u0_u7_U42 (.A2( u2_u0_u7_n102 ) , .A1( u2_u0_u7_n103 ) , .ZN( u2_u0_u7_n133 ) );
  NAND2_X1 u2_u0_u7_U43 (.A1( u2_u0_u7_n103 ) , .ZN( u2_u0_u7_n127 ) , .A2( u2_u0_u7_n99 ) );
  AOI21_X1 u2_u0_u7_U44 (.ZN( u2_u0_u7_n123 ) , .B1( u2_u0_u7_n165 ) , .B2( u2_u0_u7_n177 ) , .A( u2_u0_u7_n97 ) );
  AOI21_X1 u2_u0_u7_U45 (.B2( u2_u0_u7_n113 ) , .B1( u2_u0_u7_n124 ) , .A( u2_u0_u7_n125 ) , .ZN( u2_u0_u7_n97 ) );
  INV_X1 u2_u0_u7_U46 (.A( u2_u0_u7_n152 ) , .ZN( u2_u0_u7_n162 ) );
  AND2_X1 u2_u0_u7_U47 (.ZN( u2_u0_u7_n145 ) , .A2( u2_u0_u7_n98 ) , .A1( u2_u0_u7_n99 ) );
  NOR2_X1 u2_u0_u7_U48 (.ZN( u2_u0_u7_n137 ) , .A1( u2_u0_u7_n150 ) , .A2( u2_u0_u7_n161 ) );
  AOI21_X1 u2_u0_u7_U49 (.ZN( u2_u0_u7_n105 ) , .B2( u2_u0_u7_n110 ) , .A( u2_u0_u7_n125 ) , .B1( u2_u0_u7_n147 ) );
  INV_X1 u2_u0_u7_U5 (.A( u2_u0_u7_n154 ) , .ZN( u2_u0_u7_n178 ) );
  NAND2_X1 u2_u0_u7_U50 (.A2( u2_u0_u7_n103 ) , .ZN( u2_u0_u7_n147 ) , .A1( u2_u0_u7_n93 ) );
  NAND2_X1 u2_u0_u7_U51 (.ZN( u2_u0_u7_n146 ) , .A1( u2_u0_u7_n95 ) , .A2( u2_u0_u7_n98 ) );
  OR2_X1 u2_u0_u7_U52 (.ZN( u2_u0_u7_n126 ) , .A2( u2_u0_u7_n152 ) , .A1( u2_u0_u7_n156 ) );
  NAND2_X1 u2_u0_u7_U53 (.ZN( u2_u0_u7_n112 ) , .A2( u2_u0_u7_n96 ) , .A1( u2_u0_u7_n99 ) );
  NAND2_X1 u2_u0_u7_U54 (.A2( u2_u0_u7_n102 ) , .ZN( u2_u0_u7_n128 ) , .A1( u2_u0_u7_n98 ) );
  NAND2_X1 u2_u0_u7_U55 (.A1( u2_u0_u7_n100 ) , .ZN( u2_u0_u7_n113 ) , .A2( u2_u0_u7_n93 ) );
  NAND2_X1 u2_u0_u7_U56 (.ZN( u2_u0_u7_n110 ) , .A1( u2_u0_u7_n95 ) , .A2( u2_u0_u7_n96 ) );
  INV_X1 u2_u0_u7_U57 (.A( u2_u0_u7_n150 ) , .ZN( u2_u0_u7_n164 ) );
  AND2_X1 u2_u0_u7_U58 (.ZN( u2_u0_u7_n134 ) , .A1( u2_u0_u7_n93 ) , .A2( u2_u0_u7_n98 ) );
  NAND2_X1 u2_u0_u7_U59 (.A2( u2_u0_u7_n103 ) , .ZN( u2_u0_u7_n131 ) , .A1( u2_u0_u7_n95 ) );
  INV_X1 u2_u0_u7_U6 (.A( u2_u0_u7_n149 ) , .ZN( u2_u0_u7_n175 ) );
  NAND2_X1 u2_u0_u7_U60 (.A2( u2_u0_u7_n102 ) , .ZN( u2_u0_u7_n124 ) , .A1( u2_u0_u7_n96 ) );
  NAND2_X1 u2_u0_u7_U61 (.A1( u2_u0_u7_n100 ) , .A2( u2_u0_u7_n102 ) , .ZN( u2_u0_u7_n129 ) );
  NAND2_X1 u2_u0_u7_U62 (.A1( u2_u0_u7_n100 ) , .ZN( u2_u0_u7_n138 ) , .A2( u2_u0_u7_n99 ) );
  NAND2_X1 u2_u0_u7_U63 (.ZN( u2_u0_u7_n132 ) , .A1( u2_u0_u7_n93 ) , .A2( u2_u0_u7_n96 ) );
  NAND2_X1 u2_u0_u7_U64 (.A1( u2_u0_u7_n100 ) , .ZN( u2_u0_u7_n148 ) , .A2( u2_u0_u7_n95 ) );
  AOI22_X1 u2_u0_u7_U65 (.A2( u2_u0_u7_n114 ) , .ZN( u2_u0_u7_n119 ) , .B1( u2_u0_u7_n130 ) , .A1( u2_u0_u7_n156 ) , .B2( u2_u0_u7_n165 ) );
  NAND2_X1 u2_u0_u7_U66 (.A2( u2_u0_u7_n112 ) , .ZN( u2_u0_u7_n114 ) , .A1( u2_u0_u7_n175 ) );
  NOR2_X1 u2_u0_u7_U67 (.A2( u2_u0_X_47 ) , .ZN( u2_u0_u7_n150 ) , .A1( u2_u0_u7_n163 ) );
  NOR2_X1 u2_u0_u7_U68 (.A2( u2_u0_X_48 ) , .A1( u2_u0_u7_n166 ) , .ZN( u2_u0_u7_n95 ) );
  NOR2_X1 u2_u0_u7_U69 (.A2( u2_u0_X_45 ) , .A1( u2_u0_X_48 ) , .ZN( u2_u0_u7_n99 ) );
  AOI211_X1 u2_u0_u7_U7 (.ZN( u2_u0_u7_n116 ) , .A( u2_u0_u7_n155 ) , .C1( u2_u0_u7_n161 ) , .C2( u2_u0_u7_n171 ) , .B( u2_u0_u7_n94 ) );
  NOR2_X1 u2_u0_u7_U70 (.A2( u2_u0_X_44 ) , .A1( u2_u0_u7_n167 ) , .ZN( u2_u0_u7_n98 ) );
  NOR2_X1 u2_u0_u7_U71 (.A2( u2_u0_X_46 ) , .A1( u2_u0_X_47 ) , .ZN( u2_u0_u7_n152 ) );
  AND2_X1 u2_u0_u7_U72 (.A1( u2_u0_X_47 ) , .ZN( u2_u0_u7_n156 ) , .A2( u2_u0_u7_n163 ) );
  NAND2_X1 u2_u0_u7_U73 (.A2( u2_u0_X_46 ) , .A1( u2_u0_X_47 ) , .ZN( u2_u0_u7_n125 ) );
  AND2_X1 u2_u0_u7_U74 (.A2( u2_u0_X_45 ) , .A1( u2_u0_X_48 ) , .ZN( u2_u0_u7_n102 ) );
  AND2_X1 u2_u0_u7_U75 (.A2( u2_u0_X_43 ) , .A1( u2_u0_X_44 ) , .ZN( u2_u0_u7_n96 ) );
  AND2_X1 u2_u0_u7_U76 (.A1( u2_u0_X_44 ) , .ZN( u2_u0_u7_n100 ) , .A2( u2_u0_u7_n167 ) );
  AND2_X1 u2_u0_u7_U77 (.A1( u2_u0_X_48 ) , .A2( u2_u0_u7_n166 ) , .ZN( u2_u0_u7_n93 ) );
  INV_X1 u2_u0_u7_U78 (.A( u2_u0_X_46 ) , .ZN( u2_u0_u7_n163 ) );
  INV_X1 u2_u0_u7_U79 (.A( u2_u0_X_45 ) , .ZN( u2_u0_u7_n166 ) );
  OAI222_X1 u2_u0_u7_U8 (.C2( u2_u0_u7_n101 ) , .B2( u2_u0_u7_n111 ) , .A1( u2_u0_u7_n113 ) , .C1( u2_u0_u7_n146 ) , .A2( u2_u0_u7_n162 ) , .B1( u2_u0_u7_n164 ) , .ZN( u2_u0_u7_n94 ) );
  OAI21_X1 u2_u0_u7_U80 (.B1( u2_u0_u7_n145 ) , .ZN( u2_u0_u7_n160 ) , .A( u2_u0_u7_n161 ) , .B2( u2_u0_u7_n177 ) );
  AOI22_X1 u2_u0_u7_U81 (.B2( u2_u0_u7_n149 ) , .B1( u2_u0_u7_n150 ) , .A2( u2_u0_u7_n151 ) , .A1( u2_u0_u7_n152 ) , .ZN( u2_u0_u7_n158 ) );
  NAND4_X1 u2_u0_u7_U82 (.ZN( u2_out0_27 ) , .A4( u2_u0_u7_n118 ) , .A3( u2_u0_u7_n119 ) , .A2( u2_u0_u7_n120 ) , .A1( u2_u0_u7_n121 ) );
  OAI21_X1 u2_u0_u7_U83 (.ZN( u2_u0_u7_n121 ) , .B2( u2_u0_u7_n145 ) , .A( u2_u0_u7_n150 ) , .B1( u2_u0_u7_n174 ) );
  OAI21_X1 u2_u0_u7_U84 (.ZN( u2_u0_u7_n120 ) , .A( u2_u0_u7_n161 ) , .B2( u2_u0_u7_n170 ) , .B1( u2_u0_u7_n179 ) );
  NAND4_X1 u2_u0_u7_U85 (.ZN( u2_out0_15 ) , .A4( u2_u0_u7_n142 ) , .A3( u2_u0_u7_n143 ) , .A2( u2_u0_u7_n144 ) , .A1( u2_u0_u7_n178 ) );
  OR2_X1 u2_u0_u7_U86 (.A2( u2_u0_u7_n125 ) , .A1( u2_u0_u7_n129 ) , .ZN( u2_u0_u7_n144 ) );
  AOI22_X1 u2_u0_u7_U87 (.A2( u2_u0_u7_n126 ) , .ZN( u2_u0_u7_n143 ) , .B2( u2_u0_u7_n165 ) , .B1( u2_u0_u7_n173 ) , .A1( u2_u0_u7_n174 ) );
  NAND4_X1 u2_u0_u7_U88 (.ZN( u2_out0_5 ) , .A4( u2_u0_u7_n108 ) , .A3( u2_u0_u7_n109 ) , .A1( u2_u0_u7_n116 ) , .A2( u2_u0_u7_n123 ) );
  AOI22_X1 u2_u0_u7_U89 (.ZN( u2_u0_u7_n109 ) , .A2( u2_u0_u7_n126 ) , .B2( u2_u0_u7_n145 ) , .B1( u2_u0_u7_n156 ) , .A1( u2_u0_u7_n171 ) );
  AOI222_X1 u2_u0_u7_U9 (.ZN( u2_u0_u7_n122 ) , .C2( u2_u0_u7_n126 ) , .C1( u2_u0_u7_n145 ) , .B1( u2_u0_u7_n161 ) , .A2( u2_u0_u7_n165 ) , .B2( u2_u0_u7_n170 ) , .A1( u2_u0_u7_n176 ) );
  NOR4_X1 u2_u0_u7_U90 (.A4( u2_u0_u7_n104 ) , .A3( u2_u0_u7_n105 ) , .A2( u2_u0_u7_n106 ) , .A1( u2_u0_u7_n107 ) , .ZN( u2_u0_u7_n108 ) );
  NAND4_X1 u2_u0_u7_U91 (.ZN( u2_out0_21 ) , .A4( u2_u0_u7_n157 ) , .A3( u2_u0_u7_n158 ) , .A2( u2_u0_u7_n159 ) , .A1( u2_u0_u7_n160 ) );
  OAI211_X1 u2_u0_u7_U92 (.B( u2_u0_u7_n122 ) , .A( u2_u0_u7_n123 ) , .C2( u2_u0_u7_n124 ) , .ZN( u2_u0_u7_n154 ) , .C1( u2_u0_u7_n162 ) );
  NOR2_X1 u2_u0_u7_U93 (.A2( u2_u0_X_43 ) , .A1( u2_u0_X_44 ) , .ZN( u2_u0_u7_n103 ) );
  INV_X1 u2_u0_u7_U94 (.A( u2_u0_X_43 ) , .ZN( u2_u0_u7_n167 ) );
  NAND3_X1 u2_u0_u7_U95 (.A3( u2_u0_u7_n146 ) , .A2( u2_u0_u7_n147 ) , .A1( u2_u0_u7_n148 ) , .ZN( u2_u0_u7_n151 ) );
  NAND3_X1 u2_u0_u7_U96 (.A3( u2_u0_u7_n131 ) , .A2( u2_u0_u7_n132 ) , .A1( u2_u0_u7_n133 ) , .ZN( u2_u0_u7_n135 ) );
  XOR2_X1 u2_u10_U25 (.B( u2_K11_31 ) , .A( u2_R9_20 ) , .Z( u2_u10_X_31 ) );
  XOR2_X1 u2_u10_U28 (.B( u2_K11_29 ) , .A( u2_R9_20 ) , .Z( u2_u10_X_29 ) );
  XOR2_X1 u2_u10_U31 (.B( u2_K11_26 ) , .A( u2_R9_17 ) , .Z( u2_u10_X_26 ) );
  XOR2_X1 u2_u10_U33 (.B( u2_K11_24 ) , .A( u2_R9_17 ) , .Z( u2_u10_X_24 ) );
  XOR2_X1 u2_u10_U37 (.B( u2_K11_20 ) , .A( u2_R9_13 ) , .Z( u2_u10_X_20 ) );
  XOR2_X1 u2_u10_U39 (.B( u2_K11_19 ) , .A( u2_R9_12 ) , .Z( u2_u10_X_19 ) );
  XOR2_X1 u2_u10_U8 (.B( u2_K11_47 ) , .A( u2_R9_32 ) , .Z( u2_u10_X_47 ) );
  OAI22_X1 u2_u10_u3_U10 (.B1( u2_u10_u3_n113 ) , .A2( u2_u10_u3_n135 ) , .A1( u2_u10_u3_n150 ) , .B2( u2_u10_u3_n164 ) , .ZN( u2_u10_u3_n98 ) );
  OAI211_X1 u2_u10_u3_U11 (.B( u2_u10_u3_n106 ) , .ZN( u2_u10_u3_n119 ) , .C2( u2_u10_u3_n128 ) , .C1( u2_u10_u3_n167 ) , .A( u2_u10_u3_n181 ) );
  AOI221_X1 u2_u10_u3_U12 (.C1( u2_u10_u3_n105 ) , .ZN( u2_u10_u3_n106 ) , .A( u2_u10_u3_n131 ) , .B2( u2_u10_u3_n132 ) , .C2( u2_u10_u3_n133 ) , .B1( u2_u10_u3_n169 ) );
  INV_X1 u2_u10_u3_U13 (.ZN( u2_u10_u3_n181 ) , .A( u2_u10_u3_n98 ) );
  NAND2_X1 u2_u10_u3_U14 (.ZN( u2_u10_u3_n105 ) , .A2( u2_u10_u3_n130 ) , .A1( u2_u10_u3_n155 ) );
  AOI22_X1 u2_u10_u3_U15 (.B1( u2_u10_u3_n115 ) , .A2( u2_u10_u3_n116 ) , .ZN( u2_u10_u3_n123 ) , .B2( u2_u10_u3_n133 ) , .A1( u2_u10_u3_n169 ) );
  NAND2_X1 u2_u10_u3_U16 (.ZN( u2_u10_u3_n116 ) , .A2( u2_u10_u3_n151 ) , .A1( u2_u10_u3_n182 ) );
  NOR2_X1 u2_u10_u3_U17 (.ZN( u2_u10_u3_n126 ) , .A2( u2_u10_u3_n150 ) , .A1( u2_u10_u3_n164 ) );
  AOI21_X1 u2_u10_u3_U18 (.ZN( u2_u10_u3_n112 ) , .B2( u2_u10_u3_n146 ) , .B1( u2_u10_u3_n155 ) , .A( u2_u10_u3_n167 ) );
  NAND2_X1 u2_u10_u3_U19 (.A1( u2_u10_u3_n135 ) , .ZN( u2_u10_u3_n142 ) , .A2( u2_u10_u3_n164 ) );
  NAND2_X1 u2_u10_u3_U20 (.ZN( u2_u10_u3_n132 ) , .A2( u2_u10_u3_n152 ) , .A1( u2_u10_u3_n156 ) );
  AND2_X1 u2_u10_u3_U21 (.A2( u2_u10_u3_n113 ) , .A1( u2_u10_u3_n114 ) , .ZN( u2_u10_u3_n151 ) );
  INV_X1 u2_u10_u3_U22 (.A( u2_u10_u3_n133 ) , .ZN( u2_u10_u3_n165 ) );
  INV_X1 u2_u10_u3_U23 (.A( u2_u10_u3_n135 ) , .ZN( u2_u10_u3_n170 ) );
  NAND2_X1 u2_u10_u3_U24 (.A1( u2_u10_u3_n107 ) , .A2( u2_u10_u3_n108 ) , .ZN( u2_u10_u3_n140 ) );
  NAND2_X1 u2_u10_u3_U25 (.ZN( u2_u10_u3_n117 ) , .A1( u2_u10_u3_n124 ) , .A2( u2_u10_u3_n148 ) );
  NAND2_X1 u2_u10_u3_U26 (.ZN( u2_u10_u3_n143 ) , .A1( u2_u10_u3_n165 ) , .A2( u2_u10_u3_n167 ) );
  INV_X1 u2_u10_u3_U27 (.A( u2_u10_u3_n130 ) , .ZN( u2_u10_u3_n177 ) );
  INV_X1 u2_u10_u3_U28 (.A( u2_u10_u3_n128 ) , .ZN( u2_u10_u3_n176 ) );
  INV_X1 u2_u10_u3_U29 (.A( u2_u10_u3_n155 ) , .ZN( u2_u10_u3_n174 ) );
  INV_X1 u2_u10_u3_U3 (.A( u2_u10_u3_n129 ) , .ZN( u2_u10_u3_n183 ) );
  INV_X1 u2_u10_u3_U30 (.A( u2_u10_u3_n139 ) , .ZN( u2_u10_u3_n185 ) );
  NOR2_X1 u2_u10_u3_U31 (.ZN( u2_u10_u3_n135 ) , .A2( u2_u10_u3_n141 ) , .A1( u2_u10_u3_n169 ) );
  OAI222_X1 u2_u10_u3_U32 (.C2( u2_u10_u3_n107 ) , .A2( u2_u10_u3_n108 ) , .B1( u2_u10_u3_n135 ) , .ZN( u2_u10_u3_n138 ) , .B2( u2_u10_u3_n146 ) , .C1( u2_u10_u3_n154 ) , .A1( u2_u10_u3_n164 ) );
  NOR4_X1 u2_u10_u3_U33 (.A4( u2_u10_u3_n157 ) , .A3( u2_u10_u3_n158 ) , .A2( u2_u10_u3_n159 ) , .A1( u2_u10_u3_n160 ) , .ZN( u2_u10_u3_n161 ) );
  AOI21_X1 u2_u10_u3_U34 (.B2( u2_u10_u3_n152 ) , .B1( u2_u10_u3_n153 ) , .ZN( u2_u10_u3_n158 ) , .A( u2_u10_u3_n164 ) );
  AOI21_X1 u2_u10_u3_U35 (.A( u2_u10_u3_n154 ) , .B2( u2_u10_u3_n155 ) , .B1( u2_u10_u3_n156 ) , .ZN( u2_u10_u3_n157 ) );
  AOI21_X1 u2_u10_u3_U36 (.A( u2_u10_u3_n149 ) , .B2( u2_u10_u3_n150 ) , .B1( u2_u10_u3_n151 ) , .ZN( u2_u10_u3_n159 ) );
  AOI211_X1 u2_u10_u3_U37 (.ZN( u2_u10_u3_n109 ) , .A( u2_u10_u3_n119 ) , .C2( u2_u10_u3_n129 ) , .B( u2_u10_u3_n138 ) , .C1( u2_u10_u3_n141 ) );
  AOI211_X1 u2_u10_u3_U38 (.B( u2_u10_u3_n119 ) , .A( u2_u10_u3_n120 ) , .C2( u2_u10_u3_n121 ) , .ZN( u2_u10_u3_n122 ) , .C1( u2_u10_u3_n179 ) );
  INV_X1 u2_u10_u3_U39 (.A( u2_u10_u3_n156 ) , .ZN( u2_u10_u3_n179 ) );
  INV_X1 u2_u10_u3_U4 (.A( u2_u10_u3_n140 ) , .ZN( u2_u10_u3_n182 ) );
  OAI22_X1 u2_u10_u3_U40 (.B1( u2_u10_u3_n118 ) , .ZN( u2_u10_u3_n120 ) , .A1( u2_u10_u3_n135 ) , .B2( u2_u10_u3_n154 ) , .A2( u2_u10_u3_n178 ) );
  AND3_X1 u2_u10_u3_U41 (.ZN( u2_u10_u3_n118 ) , .A2( u2_u10_u3_n124 ) , .A1( u2_u10_u3_n144 ) , .A3( u2_u10_u3_n152 ) );
  INV_X1 u2_u10_u3_U42 (.A( u2_u10_u3_n121 ) , .ZN( u2_u10_u3_n164 ) );
  NAND2_X1 u2_u10_u3_U43 (.ZN( u2_u10_u3_n133 ) , .A1( u2_u10_u3_n154 ) , .A2( u2_u10_u3_n164 ) );
  OAI211_X1 u2_u10_u3_U44 (.B( u2_u10_u3_n127 ) , .ZN( u2_u10_u3_n139 ) , .C1( u2_u10_u3_n150 ) , .C2( u2_u10_u3_n154 ) , .A( u2_u10_u3_n184 ) );
  INV_X1 u2_u10_u3_U45 (.A( u2_u10_u3_n125 ) , .ZN( u2_u10_u3_n184 ) );
  AOI221_X1 u2_u10_u3_U46 (.A( u2_u10_u3_n126 ) , .ZN( u2_u10_u3_n127 ) , .C2( u2_u10_u3_n132 ) , .C1( u2_u10_u3_n169 ) , .B2( u2_u10_u3_n170 ) , .B1( u2_u10_u3_n174 ) );
  OAI22_X1 u2_u10_u3_U47 (.A1( u2_u10_u3_n124 ) , .ZN( u2_u10_u3_n125 ) , .B2( u2_u10_u3_n145 ) , .A2( u2_u10_u3_n165 ) , .B1( u2_u10_u3_n167 ) );
  NOR2_X1 u2_u10_u3_U48 (.A1( u2_u10_u3_n113 ) , .ZN( u2_u10_u3_n131 ) , .A2( u2_u10_u3_n154 ) );
  NAND2_X1 u2_u10_u3_U49 (.A1( u2_u10_u3_n103 ) , .ZN( u2_u10_u3_n150 ) , .A2( u2_u10_u3_n99 ) );
  INV_X1 u2_u10_u3_U5 (.A( u2_u10_u3_n117 ) , .ZN( u2_u10_u3_n178 ) );
  NAND2_X1 u2_u10_u3_U50 (.A2( u2_u10_u3_n102 ) , .ZN( u2_u10_u3_n155 ) , .A1( u2_u10_u3_n97 ) );
  INV_X1 u2_u10_u3_U51 (.A( u2_u10_u3_n141 ) , .ZN( u2_u10_u3_n167 ) );
  AOI21_X1 u2_u10_u3_U52 (.B2( u2_u10_u3_n114 ) , .B1( u2_u10_u3_n146 ) , .A( u2_u10_u3_n154 ) , .ZN( u2_u10_u3_n94 ) );
  AOI21_X1 u2_u10_u3_U53 (.ZN( u2_u10_u3_n110 ) , .B2( u2_u10_u3_n142 ) , .B1( u2_u10_u3_n186 ) , .A( u2_u10_u3_n95 ) );
  INV_X1 u2_u10_u3_U54 (.A( u2_u10_u3_n145 ) , .ZN( u2_u10_u3_n186 ) );
  AOI21_X1 u2_u10_u3_U55 (.B1( u2_u10_u3_n124 ) , .A( u2_u10_u3_n149 ) , .B2( u2_u10_u3_n155 ) , .ZN( u2_u10_u3_n95 ) );
  INV_X1 u2_u10_u3_U56 (.A( u2_u10_u3_n149 ) , .ZN( u2_u10_u3_n169 ) );
  NAND2_X1 u2_u10_u3_U57 (.ZN( u2_u10_u3_n124 ) , .A1( u2_u10_u3_n96 ) , .A2( u2_u10_u3_n97 ) );
  NAND2_X1 u2_u10_u3_U58 (.A2( u2_u10_u3_n100 ) , .ZN( u2_u10_u3_n146 ) , .A1( u2_u10_u3_n96 ) );
  NAND2_X1 u2_u10_u3_U59 (.A1( u2_u10_u3_n101 ) , .ZN( u2_u10_u3_n145 ) , .A2( u2_u10_u3_n99 ) );
  AOI221_X1 u2_u10_u3_U6 (.A( u2_u10_u3_n131 ) , .C2( u2_u10_u3_n132 ) , .C1( u2_u10_u3_n133 ) , .ZN( u2_u10_u3_n134 ) , .B1( u2_u10_u3_n143 ) , .B2( u2_u10_u3_n177 ) );
  NAND2_X1 u2_u10_u3_U60 (.A1( u2_u10_u3_n100 ) , .ZN( u2_u10_u3_n156 ) , .A2( u2_u10_u3_n99 ) );
  NAND2_X1 u2_u10_u3_U61 (.A2( u2_u10_u3_n101 ) , .A1( u2_u10_u3_n104 ) , .ZN( u2_u10_u3_n148 ) );
  NAND2_X1 u2_u10_u3_U62 (.A1( u2_u10_u3_n100 ) , .A2( u2_u10_u3_n102 ) , .ZN( u2_u10_u3_n128 ) );
  NAND2_X1 u2_u10_u3_U63 (.A2( u2_u10_u3_n101 ) , .A1( u2_u10_u3_n102 ) , .ZN( u2_u10_u3_n152 ) );
  NAND2_X1 u2_u10_u3_U64 (.A2( u2_u10_u3_n101 ) , .ZN( u2_u10_u3_n114 ) , .A1( u2_u10_u3_n96 ) );
  NAND2_X1 u2_u10_u3_U65 (.ZN( u2_u10_u3_n107 ) , .A1( u2_u10_u3_n97 ) , .A2( u2_u10_u3_n99 ) );
  NAND2_X1 u2_u10_u3_U66 (.A2( u2_u10_u3_n100 ) , .A1( u2_u10_u3_n104 ) , .ZN( u2_u10_u3_n113 ) );
  NAND2_X1 u2_u10_u3_U67 (.A1( u2_u10_u3_n104 ) , .ZN( u2_u10_u3_n153 ) , .A2( u2_u10_u3_n97 ) );
  NAND2_X1 u2_u10_u3_U68 (.A2( u2_u10_u3_n103 ) , .A1( u2_u10_u3_n104 ) , .ZN( u2_u10_u3_n130 ) );
  NAND2_X1 u2_u10_u3_U69 (.A2( u2_u10_u3_n103 ) , .ZN( u2_u10_u3_n144 ) , .A1( u2_u10_u3_n96 ) );
  OAI22_X1 u2_u10_u3_U7 (.B2( u2_u10_u3_n147 ) , .A2( u2_u10_u3_n148 ) , .ZN( u2_u10_u3_n160 ) , .B1( u2_u10_u3_n165 ) , .A1( u2_u10_u3_n168 ) );
  NAND2_X1 u2_u10_u3_U70 (.A1( u2_u10_u3_n102 ) , .A2( u2_u10_u3_n103 ) , .ZN( u2_u10_u3_n108 ) );
  NOR2_X1 u2_u10_u3_U71 (.A2( u2_u10_X_19 ) , .A1( u2_u10_X_20 ) , .ZN( u2_u10_u3_n99 ) );
  NOR2_X1 u2_u10_u3_U72 (.A2( u2_u10_X_21 ) , .A1( u2_u10_X_24 ) , .ZN( u2_u10_u3_n103 ) );
  NOR2_X1 u2_u10_u3_U73 (.A2( u2_u10_X_24 ) , .A1( u2_u10_u3_n171 ) , .ZN( u2_u10_u3_n97 ) );
  NOR2_X1 u2_u10_u3_U74 (.A2( u2_u10_X_23 ) , .ZN( u2_u10_u3_n141 ) , .A1( u2_u10_u3_n166 ) );
  NOR2_X1 u2_u10_u3_U75 (.A2( u2_u10_X_19 ) , .A1( u2_u10_u3_n172 ) , .ZN( u2_u10_u3_n96 ) );
  NAND2_X1 u2_u10_u3_U76 (.A1( u2_u10_X_22 ) , .A2( u2_u10_X_23 ) , .ZN( u2_u10_u3_n154 ) );
  NAND2_X1 u2_u10_u3_U77 (.A1( u2_u10_X_23 ) , .ZN( u2_u10_u3_n149 ) , .A2( u2_u10_u3_n166 ) );
  NOR2_X1 u2_u10_u3_U78 (.A2( u2_u10_X_22 ) , .A1( u2_u10_X_23 ) , .ZN( u2_u10_u3_n121 ) );
  AND2_X1 u2_u10_u3_U79 (.A1( u2_u10_X_24 ) , .ZN( u2_u10_u3_n101 ) , .A2( u2_u10_u3_n171 ) );
  AND3_X1 u2_u10_u3_U8 (.A3( u2_u10_u3_n144 ) , .A2( u2_u10_u3_n145 ) , .A1( u2_u10_u3_n146 ) , .ZN( u2_u10_u3_n147 ) );
  AND2_X1 u2_u10_u3_U80 (.A1( u2_u10_X_19 ) , .ZN( u2_u10_u3_n102 ) , .A2( u2_u10_u3_n172 ) );
  AND2_X1 u2_u10_u3_U81 (.A1( u2_u10_X_21 ) , .A2( u2_u10_X_24 ) , .ZN( u2_u10_u3_n100 ) );
  AND2_X1 u2_u10_u3_U82 (.A2( u2_u10_X_19 ) , .A1( u2_u10_X_20 ) , .ZN( u2_u10_u3_n104 ) );
  INV_X1 u2_u10_u3_U83 (.A( u2_u10_X_22 ) , .ZN( u2_u10_u3_n166 ) );
  INV_X1 u2_u10_u3_U84 (.A( u2_u10_X_21 ) , .ZN( u2_u10_u3_n171 ) );
  INV_X1 u2_u10_u3_U85 (.A( u2_u10_X_20 ) , .ZN( u2_u10_u3_n172 ) );
  OR4_X1 u2_u10_u3_U86 (.ZN( u2_out10_10 ) , .A4( u2_u10_u3_n136 ) , .A3( u2_u10_u3_n137 ) , .A1( u2_u10_u3_n138 ) , .A2( u2_u10_u3_n139 ) );
  OAI222_X1 u2_u10_u3_U87 (.C1( u2_u10_u3_n128 ) , .ZN( u2_u10_u3_n137 ) , .B1( u2_u10_u3_n148 ) , .A2( u2_u10_u3_n150 ) , .B2( u2_u10_u3_n154 ) , .C2( u2_u10_u3_n164 ) , .A1( u2_u10_u3_n167 ) );
  OAI221_X1 u2_u10_u3_U88 (.A( u2_u10_u3_n134 ) , .B2( u2_u10_u3_n135 ) , .ZN( u2_u10_u3_n136 ) , .C1( u2_u10_u3_n149 ) , .B1( u2_u10_u3_n151 ) , .C2( u2_u10_u3_n183 ) );
  NAND4_X1 u2_u10_u3_U89 (.ZN( u2_out10_26 ) , .A4( u2_u10_u3_n109 ) , .A3( u2_u10_u3_n110 ) , .A2( u2_u10_u3_n111 ) , .A1( u2_u10_u3_n173 ) );
  INV_X1 u2_u10_u3_U9 (.A( u2_u10_u3_n143 ) , .ZN( u2_u10_u3_n168 ) );
  INV_X1 u2_u10_u3_U90 (.ZN( u2_u10_u3_n173 ) , .A( u2_u10_u3_n94 ) );
  OAI21_X1 u2_u10_u3_U91 (.ZN( u2_u10_u3_n111 ) , .B2( u2_u10_u3_n117 ) , .A( u2_u10_u3_n133 ) , .B1( u2_u10_u3_n176 ) );
  NAND4_X1 u2_u10_u3_U92 (.ZN( u2_out10_20 ) , .A4( u2_u10_u3_n122 ) , .A3( u2_u10_u3_n123 ) , .A1( u2_u10_u3_n175 ) , .A2( u2_u10_u3_n180 ) );
  INV_X1 u2_u10_u3_U93 (.A( u2_u10_u3_n126 ) , .ZN( u2_u10_u3_n180 ) );
  INV_X1 u2_u10_u3_U94 (.A( u2_u10_u3_n112 ) , .ZN( u2_u10_u3_n175 ) );
  NAND4_X1 u2_u10_u3_U95 (.ZN( u2_out10_1 ) , .A4( u2_u10_u3_n161 ) , .A3( u2_u10_u3_n162 ) , .A2( u2_u10_u3_n163 ) , .A1( u2_u10_u3_n185 ) );
  NAND2_X1 u2_u10_u3_U96 (.ZN( u2_u10_u3_n163 ) , .A2( u2_u10_u3_n170 ) , .A1( u2_u10_u3_n176 ) );
  AOI22_X1 u2_u10_u3_U97 (.B2( u2_u10_u3_n140 ) , .B1( u2_u10_u3_n141 ) , .A2( u2_u10_u3_n142 ) , .ZN( u2_u10_u3_n162 ) , .A1( u2_u10_u3_n177 ) );
  NAND3_X1 u2_u10_u3_U98 (.A1( u2_u10_u3_n114 ) , .ZN( u2_u10_u3_n115 ) , .A2( u2_u10_u3_n145 ) , .A3( u2_u10_u3_n153 ) );
  NAND3_X1 u2_u10_u3_U99 (.ZN( u2_u10_u3_n129 ) , .A2( u2_u10_u3_n144 ) , .A1( u2_u10_u3_n153 ) , .A3( u2_u10_u3_n182 ) );
  AOI21_X1 u2_u10_u4_U10 (.ZN( u2_u10_u4_n106 ) , .B2( u2_u10_u4_n146 ) , .B1( u2_u10_u4_n158 ) , .A( u2_u10_u4_n170 ) );
  AOI21_X1 u2_u10_u4_U11 (.ZN( u2_u10_u4_n108 ) , .B2( u2_u10_u4_n134 ) , .B1( u2_u10_u4_n155 ) , .A( u2_u10_u4_n156 ) );
  AOI21_X1 u2_u10_u4_U12 (.ZN( u2_u10_u4_n109 ) , .A( u2_u10_u4_n153 ) , .B1( u2_u10_u4_n159 ) , .B2( u2_u10_u4_n184 ) );
  AOI211_X1 u2_u10_u4_U13 (.B( u2_u10_u4_n136 ) , .A( u2_u10_u4_n137 ) , .C2( u2_u10_u4_n138 ) , .ZN( u2_u10_u4_n139 ) , .C1( u2_u10_u4_n182 ) );
  OAI22_X1 u2_u10_u4_U14 (.B2( u2_u10_u4_n135 ) , .ZN( u2_u10_u4_n137 ) , .B1( u2_u10_u4_n153 ) , .A1( u2_u10_u4_n155 ) , .A2( u2_u10_u4_n171 ) );
  AND3_X1 u2_u10_u4_U15 (.A2( u2_u10_u4_n134 ) , .ZN( u2_u10_u4_n135 ) , .A3( u2_u10_u4_n145 ) , .A1( u2_u10_u4_n157 ) );
  NAND2_X1 u2_u10_u4_U16 (.ZN( u2_u10_u4_n132 ) , .A2( u2_u10_u4_n170 ) , .A1( u2_u10_u4_n173 ) );
  AOI21_X1 u2_u10_u4_U17 (.B2( u2_u10_u4_n160 ) , .B1( u2_u10_u4_n161 ) , .ZN( u2_u10_u4_n162 ) , .A( u2_u10_u4_n170 ) );
  AOI21_X1 u2_u10_u4_U18 (.ZN( u2_u10_u4_n107 ) , .B2( u2_u10_u4_n143 ) , .A( u2_u10_u4_n174 ) , .B1( u2_u10_u4_n184 ) );
  AOI21_X1 u2_u10_u4_U19 (.B2( u2_u10_u4_n158 ) , .B1( u2_u10_u4_n159 ) , .ZN( u2_u10_u4_n163 ) , .A( u2_u10_u4_n174 ) );
  AOI21_X1 u2_u10_u4_U20 (.A( u2_u10_u4_n153 ) , .B2( u2_u10_u4_n154 ) , .B1( u2_u10_u4_n155 ) , .ZN( u2_u10_u4_n165 ) );
  AOI21_X1 u2_u10_u4_U21 (.A( u2_u10_u4_n156 ) , .B2( u2_u10_u4_n157 ) , .ZN( u2_u10_u4_n164 ) , .B1( u2_u10_u4_n184 ) );
  INV_X1 u2_u10_u4_U22 (.A( u2_u10_u4_n138 ) , .ZN( u2_u10_u4_n170 ) );
  AND2_X1 u2_u10_u4_U23 (.A2( u2_u10_u4_n120 ) , .ZN( u2_u10_u4_n155 ) , .A1( u2_u10_u4_n160 ) );
  INV_X1 u2_u10_u4_U24 (.A( u2_u10_u4_n156 ) , .ZN( u2_u10_u4_n175 ) );
  NAND2_X1 u2_u10_u4_U25 (.A2( u2_u10_u4_n118 ) , .ZN( u2_u10_u4_n131 ) , .A1( u2_u10_u4_n147 ) );
  NAND2_X1 u2_u10_u4_U26 (.A1( u2_u10_u4_n119 ) , .A2( u2_u10_u4_n120 ) , .ZN( u2_u10_u4_n130 ) );
  NAND2_X1 u2_u10_u4_U27 (.ZN( u2_u10_u4_n117 ) , .A2( u2_u10_u4_n118 ) , .A1( u2_u10_u4_n148 ) );
  NAND2_X1 u2_u10_u4_U28 (.ZN( u2_u10_u4_n129 ) , .A1( u2_u10_u4_n134 ) , .A2( u2_u10_u4_n148 ) );
  AND3_X1 u2_u10_u4_U29 (.A1( u2_u10_u4_n119 ) , .A2( u2_u10_u4_n143 ) , .A3( u2_u10_u4_n154 ) , .ZN( u2_u10_u4_n161 ) );
  NOR2_X1 u2_u10_u4_U3 (.ZN( u2_u10_u4_n121 ) , .A1( u2_u10_u4_n181 ) , .A2( u2_u10_u4_n182 ) );
  AND2_X1 u2_u10_u4_U30 (.A1( u2_u10_u4_n145 ) , .A2( u2_u10_u4_n147 ) , .ZN( u2_u10_u4_n159 ) );
  OR3_X1 u2_u10_u4_U31 (.A3( u2_u10_u4_n114 ) , .A2( u2_u10_u4_n115 ) , .A1( u2_u10_u4_n116 ) , .ZN( u2_u10_u4_n136 ) );
  AOI21_X1 u2_u10_u4_U32 (.A( u2_u10_u4_n113 ) , .ZN( u2_u10_u4_n116 ) , .B2( u2_u10_u4_n173 ) , .B1( u2_u10_u4_n174 ) );
  AOI21_X1 u2_u10_u4_U33 (.ZN( u2_u10_u4_n115 ) , .B2( u2_u10_u4_n145 ) , .B1( u2_u10_u4_n146 ) , .A( u2_u10_u4_n156 ) );
  OAI22_X1 u2_u10_u4_U34 (.ZN( u2_u10_u4_n114 ) , .A2( u2_u10_u4_n121 ) , .B1( u2_u10_u4_n160 ) , .B2( u2_u10_u4_n170 ) , .A1( u2_u10_u4_n171 ) );
  INV_X1 u2_u10_u4_U35 (.A( u2_u10_u4_n158 ) , .ZN( u2_u10_u4_n182 ) );
  INV_X1 u2_u10_u4_U36 (.ZN( u2_u10_u4_n181 ) , .A( u2_u10_u4_n96 ) );
  INV_X1 u2_u10_u4_U37 (.A( u2_u10_u4_n144 ) , .ZN( u2_u10_u4_n179 ) );
  INV_X1 u2_u10_u4_U38 (.A( u2_u10_u4_n157 ) , .ZN( u2_u10_u4_n178 ) );
  NAND2_X1 u2_u10_u4_U39 (.A2( u2_u10_u4_n154 ) , .A1( u2_u10_u4_n96 ) , .ZN( u2_u10_u4_n97 ) );
  INV_X1 u2_u10_u4_U4 (.A( u2_u10_u4_n117 ) , .ZN( u2_u10_u4_n184 ) );
  INV_X1 u2_u10_u4_U40 (.A( u2_u10_u4_n143 ) , .ZN( u2_u10_u4_n183 ) );
  NOR2_X1 u2_u10_u4_U41 (.ZN( u2_u10_u4_n138 ) , .A1( u2_u10_u4_n168 ) , .A2( u2_u10_u4_n169 ) );
  NOR2_X1 u2_u10_u4_U42 (.A1( u2_u10_u4_n150 ) , .A2( u2_u10_u4_n152 ) , .ZN( u2_u10_u4_n153 ) );
  NOR2_X1 u2_u10_u4_U43 (.A2( u2_u10_u4_n128 ) , .A1( u2_u10_u4_n138 ) , .ZN( u2_u10_u4_n156 ) );
  AOI22_X1 u2_u10_u4_U44 (.B2( u2_u10_u4_n122 ) , .A1( u2_u10_u4_n123 ) , .ZN( u2_u10_u4_n124 ) , .B1( u2_u10_u4_n128 ) , .A2( u2_u10_u4_n172 ) );
  INV_X1 u2_u10_u4_U45 (.A( u2_u10_u4_n153 ) , .ZN( u2_u10_u4_n172 ) );
  NAND2_X1 u2_u10_u4_U46 (.A2( u2_u10_u4_n120 ) , .ZN( u2_u10_u4_n123 ) , .A1( u2_u10_u4_n161 ) );
  AOI22_X1 u2_u10_u4_U47 (.B2( u2_u10_u4_n132 ) , .A2( u2_u10_u4_n133 ) , .ZN( u2_u10_u4_n140 ) , .A1( u2_u10_u4_n150 ) , .B1( u2_u10_u4_n179 ) );
  NAND2_X1 u2_u10_u4_U48 (.ZN( u2_u10_u4_n133 ) , .A2( u2_u10_u4_n146 ) , .A1( u2_u10_u4_n154 ) );
  NAND2_X1 u2_u10_u4_U49 (.A1( u2_u10_u4_n103 ) , .ZN( u2_u10_u4_n154 ) , .A2( u2_u10_u4_n98 ) );
  INV_X1 u2_u10_u4_U5 (.ZN( u2_u10_u4_n186 ) , .A( u2_u10_u4_n95 ) );
  NAND2_X1 u2_u10_u4_U50 (.A1( u2_u10_u4_n101 ) , .ZN( u2_u10_u4_n158 ) , .A2( u2_u10_u4_n99 ) );
  AOI21_X1 u2_u10_u4_U51 (.ZN( u2_u10_u4_n127 ) , .A( u2_u10_u4_n136 ) , .B2( u2_u10_u4_n150 ) , .B1( u2_u10_u4_n180 ) );
  INV_X1 u2_u10_u4_U52 (.A( u2_u10_u4_n160 ) , .ZN( u2_u10_u4_n180 ) );
  NAND2_X1 u2_u10_u4_U53 (.A2( u2_u10_u4_n104 ) , .A1( u2_u10_u4_n105 ) , .ZN( u2_u10_u4_n146 ) );
  NAND2_X1 u2_u10_u4_U54 (.A2( u2_u10_u4_n101 ) , .A1( u2_u10_u4_n102 ) , .ZN( u2_u10_u4_n160 ) );
  NAND2_X1 u2_u10_u4_U55 (.ZN( u2_u10_u4_n134 ) , .A1( u2_u10_u4_n98 ) , .A2( u2_u10_u4_n99 ) );
  NAND2_X1 u2_u10_u4_U56 (.A1( u2_u10_u4_n103 ) , .A2( u2_u10_u4_n104 ) , .ZN( u2_u10_u4_n143 ) );
  NAND2_X1 u2_u10_u4_U57 (.A2( u2_u10_u4_n105 ) , .ZN( u2_u10_u4_n145 ) , .A1( u2_u10_u4_n98 ) );
  NAND2_X1 u2_u10_u4_U58 (.A1( u2_u10_u4_n100 ) , .A2( u2_u10_u4_n105 ) , .ZN( u2_u10_u4_n120 ) );
  NAND2_X1 u2_u10_u4_U59 (.A1( u2_u10_u4_n102 ) , .A2( u2_u10_u4_n104 ) , .ZN( u2_u10_u4_n148 ) );
  OAI221_X1 u2_u10_u4_U6 (.C1( u2_u10_u4_n134 ) , .B1( u2_u10_u4_n158 ) , .B2( u2_u10_u4_n171 ) , .C2( u2_u10_u4_n173 ) , .A( u2_u10_u4_n94 ) , .ZN( u2_u10_u4_n95 ) );
  NAND2_X1 u2_u10_u4_U60 (.A2( u2_u10_u4_n100 ) , .A1( u2_u10_u4_n103 ) , .ZN( u2_u10_u4_n157 ) );
  INV_X1 u2_u10_u4_U61 (.A( u2_u10_u4_n150 ) , .ZN( u2_u10_u4_n173 ) );
  INV_X1 u2_u10_u4_U62 (.A( u2_u10_u4_n152 ) , .ZN( u2_u10_u4_n171 ) );
  NAND2_X1 u2_u10_u4_U63 (.A1( u2_u10_u4_n100 ) , .ZN( u2_u10_u4_n118 ) , .A2( u2_u10_u4_n99 ) );
  NAND2_X1 u2_u10_u4_U64 (.A2( u2_u10_u4_n100 ) , .A1( u2_u10_u4_n102 ) , .ZN( u2_u10_u4_n144 ) );
  NAND2_X1 u2_u10_u4_U65 (.A2( u2_u10_u4_n101 ) , .A1( u2_u10_u4_n105 ) , .ZN( u2_u10_u4_n96 ) );
  INV_X1 u2_u10_u4_U66 (.A( u2_u10_u4_n128 ) , .ZN( u2_u10_u4_n174 ) );
  NAND2_X1 u2_u10_u4_U67 (.A2( u2_u10_u4_n102 ) , .ZN( u2_u10_u4_n119 ) , .A1( u2_u10_u4_n98 ) );
  NAND2_X1 u2_u10_u4_U68 (.A2( u2_u10_u4_n101 ) , .A1( u2_u10_u4_n103 ) , .ZN( u2_u10_u4_n147 ) );
  NAND2_X1 u2_u10_u4_U69 (.A2( u2_u10_u4_n104 ) , .ZN( u2_u10_u4_n113 ) , .A1( u2_u10_u4_n99 ) );
  AOI222_X1 u2_u10_u4_U7 (.B2( u2_u10_u4_n132 ) , .A1( u2_u10_u4_n138 ) , .C2( u2_u10_u4_n175 ) , .A2( u2_u10_u4_n179 ) , .C1( u2_u10_u4_n181 ) , .B1( u2_u10_u4_n185 ) , .ZN( u2_u10_u4_n94 ) );
  NOR2_X1 u2_u10_u4_U70 (.A2( u2_u10_X_28 ) , .ZN( u2_u10_u4_n150 ) , .A1( u2_u10_u4_n168 ) );
  NOR2_X1 u2_u10_u4_U71 (.A2( u2_u10_X_29 ) , .ZN( u2_u10_u4_n152 ) , .A1( u2_u10_u4_n169 ) );
  NOR2_X1 u2_u10_u4_U72 (.A2( u2_u10_X_30 ) , .ZN( u2_u10_u4_n105 ) , .A1( u2_u10_u4_n176 ) );
  NOR2_X1 u2_u10_u4_U73 (.A2( u2_u10_X_26 ) , .ZN( u2_u10_u4_n100 ) , .A1( u2_u10_u4_n177 ) );
  NOR2_X1 u2_u10_u4_U74 (.A2( u2_u10_X_28 ) , .A1( u2_u10_X_29 ) , .ZN( u2_u10_u4_n128 ) );
  NOR2_X1 u2_u10_u4_U75 (.A2( u2_u10_X_27 ) , .A1( u2_u10_X_30 ) , .ZN( u2_u10_u4_n102 ) );
  NOR2_X1 u2_u10_u4_U76 (.A2( u2_u10_X_25 ) , .A1( u2_u10_X_26 ) , .ZN( u2_u10_u4_n98 ) );
  AND2_X1 u2_u10_u4_U77 (.A2( u2_u10_X_25 ) , .A1( u2_u10_X_26 ) , .ZN( u2_u10_u4_n104 ) );
  AND2_X1 u2_u10_u4_U78 (.A1( u2_u10_X_30 ) , .A2( u2_u10_u4_n176 ) , .ZN( u2_u10_u4_n99 ) );
  AND2_X1 u2_u10_u4_U79 (.A1( u2_u10_X_26 ) , .ZN( u2_u10_u4_n101 ) , .A2( u2_u10_u4_n177 ) );
  INV_X1 u2_u10_u4_U8 (.A( u2_u10_u4_n113 ) , .ZN( u2_u10_u4_n185 ) );
  AND2_X1 u2_u10_u4_U80 (.A1( u2_u10_X_27 ) , .A2( u2_u10_X_30 ) , .ZN( u2_u10_u4_n103 ) );
  INV_X1 u2_u10_u4_U81 (.A( u2_u10_X_28 ) , .ZN( u2_u10_u4_n169 ) );
  INV_X1 u2_u10_u4_U82 (.A( u2_u10_X_29 ) , .ZN( u2_u10_u4_n168 ) );
  INV_X1 u2_u10_u4_U83 (.A( u2_u10_X_25 ) , .ZN( u2_u10_u4_n177 ) );
  INV_X1 u2_u10_u4_U84 (.A( u2_u10_X_27 ) , .ZN( u2_u10_u4_n176 ) );
  NAND4_X1 u2_u10_u4_U85 (.ZN( u2_out10_25 ) , .A4( u2_u10_u4_n139 ) , .A3( u2_u10_u4_n140 ) , .A2( u2_u10_u4_n141 ) , .A1( u2_u10_u4_n142 ) );
  OAI21_X1 u2_u10_u4_U86 (.A( u2_u10_u4_n128 ) , .B2( u2_u10_u4_n129 ) , .B1( u2_u10_u4_n130 ) , .ZN( u2_u10_u4_n142 ) );
  OAI21_X1 u2_u10_u4_U87 (.B2( u2_u10_u4_n131 ) , .ZN( u2_u10_u4_n141 ) , .A( u2_u10_u4_n175 ) , .B1( u2_u10_u4_n183 ) );
  NAND4_X1 u2_u10_u4_U88 (.ZN( u2_out10_14 ) , .A4( u2_u10_u4_n124 ) , .A3( u2_u10_u4_n125 ) , .A2( u2_u10_u4_n126 ) , .A1( u2_u10_u4_n127 ) );
  AOI22_X1 u2_u10_u4_U89 (.B2( u2_u10_u4_n117 ) , .ZN( u2_u10_u4_n126 ) , .A1( u2_u10_u4_n129 ) , .B1( u2_u10_u4_n152 ) , .A2( u2_u10_u4_n175 ) );
  NOR4_X1 u2_u10_u4_U9 (.A4( u2_u10_u4_n106 ) , .A3( u2_u10_u4_n107 ) , .A2( u2_u10_u4_n108 ) , .A1( u2_u10_u4_n109 ) , .ZN( u2_u10_u4_n110 ) );
  AOI22_X1 u2_u10_u4_U90 (.ZN( u2_u10_u4_n125 ) , .B2( u2_u10_u4_n131 ) , .A2( u2_u10_u4_n132 ) , .B1( u2_u10_u4_n138 ) , .A1( u2_u10_u4_n178 ) );
  NAND4_X1 u2_u10_u4_U91 (.ZN( u2_out10_8 ) , .A4( u2_u10_u4_n110 ) , .A3( u2_u10_u4_n111 ) , .A2( u2_u10_u4_n112 ) , .A1( u2_u10_u4_n186 ) );
  NAND2_X1 u2_u10_u4_U92 (.ZN( u2_u10_u4_n112 ) , .A2( u2_u10_u4_n130 ) , .A1( u2_u10_u4_n150 ) );
  AOI22_X1 u2_u10_u4_U93 (.ZN( u2_u10_u4_n111 ) , .B2( u2_u10_u4_n132 ) , .A1( u2_u10_u4_n152 ) , .B1( u2_u10_u4_n178 ) , .A2( u2_u10_u4_n97 ) );
  AOI22_X1 u2_u10_u4_U94 (.B2( u2_u10_u4_n149 ) , .B1( u2_u10_u4_n150 ) , .A2( u2_u10_u4_n151 ) , .A1( u2_u10_u4_n152 ) , .ZN( u2_u10_u4_n167 ) );
  NOR4_X1 u2_u10_u4_U95 (.A4( u2_u10_u4_n162 ) , .A3( u2_u10_u4_n163 ) , .A2( u2_u10_u4_n164 ) , .A1( u2_u10_u4_n165 ) , .ZN( u2_u10_u4_n166 ) );
  NAND3_X1 u2_u10_u4_U96 (.ZN( u2_out10_3 ) , .A3( u2_u10_u4_n166 ) , .A1( u2_u10_u4_n167 ) , .A2( u2_u10_u4_n186 ) );
  NAND3_X1 u2_u10_u4_U97 (.A3( u2_u10_u4_n146 ) , .A2( u2_u10_u4_n147 ) , .A1( u2_u10_u4_n148 ) , .ZN( u2_u10_u4_n149 ) );
  NAND3_X1 u2_u10_u4_U98 (.A3( u2_u10_u4_n143 ) , .A2( u2_u10_u4_n144 ) , .A1( u2_u10_u4_n145 ) , .ZN( u2_u10_u4_n151 ) );
  NAND3_X1 u2_u10_u4_U99 (.A3( u2_u10_u4_n121 ) , .ZN( u2_u10_u4_n122 ) , .A2( u2_u10_u4_n144 ) , .A1( u2_u10_u4_n154 ) );
  INV_X1 u2_u10_u5_U10 (.A( u2_u10_u5_n121 ) , .ZN( u2_u10_u5_n177 ) );
  NOR3_X1 u2_u10_u5_U100 (.A3( u2_u10_u5_n141 ) , .A1( u2_u10_u5_n142 ) , .ZN( u2_u10_u5_n143 ) , .A2( u2_u10_u5_n191 ) );
  NAND4_X1 u2_u10_u5_U101 (.ZN( u2_out10_4 ) , .A4( u2_u10_u5_n112 ) , .A2( u2_u10_u5_n113 ) , .A1( u2_u10_u5_n114 ) , .A3( u2_u10_u5_n195 ) );
  AOI211_X1 u2_u10_u5_U102 (.A( u2_u10_u5_n110 ) , .C1( u2_u10_u5_n111 ) , .ZN( u2_u10_u5_n112 ) , .B( u2_u10_u5_n118 ) , .C2( u2_u10_u5_n177 ) );
  AOI222_X1 u2_u10_u5_U103 (.ZN( u2_u10_u5_n113 ) , .A1( u2_u10_u5_n131 ) , .C1( u2_u10_u5_n148 ) , .B2( u2_u10_u5_n174 ) , .C2( u2_u10_u5_n178 ) , .A2( u2_u10_u5_n179 ) , .B1( u2_u10_u5_n99 ) );
  NAND3_X1 u2_u10_u5_U104 (.A2( u2_u10_u5_n154 ) , .A3( u2_u10_u5_n158 ) , .A1( u2_u10_u5_n161 ) , .ZN( u2_u10_u5_n99 ) );
  NOR2_X1 u2_u10_u5_U11 (.ZN( u2_u10_u5_n160 ) , .A2( u2_u10_u5_n173 ) , .A1( u2_u10_u5_n177 ) );
  INV_X1 u2_u10_u5_U12 (.A( u2_u10_u5_n150 ) , .ZN( u2_u10_u5_n174 ) );
  AOI21_X1 u2_u10_u5_U13 (.A( u2_u10_u5_n160 ) , .B2( u2_u10_u5_n161 ) , .ZN( u2_u10_u5_n162 ) , .B1( u2_u10_u5_n192 ) );
  INV_X1 u2_u10_u5_U14 (.A( u2_u10_u5_n159 ) , .ZN( u2_u10_u5_n192 ) );
  AOI21_X1 u2_u10_u5_U15 (.A( u2_u10_u5_n156 ) , .B2( u2_u10_u5_n157 ) , .B1( u2_u10_u5_n158 ) , .ZN( u2_u10_u5_n163 ) );
  AOI21_X1 u2_u10_u5_U16 (.B2( u2_u10_u5_n139 ) , .B1( u2_u10_u5_n140 ) , .ZN( u2_u10_u5_n141 ) , .A( u2_u10_u5_n150 ) );
  OAI21_X1 u2_u10_u5_U17 (.A( u2_u10_u5_n133 ) , .B2( u2_u10_u5_n134 ) , .B1( u2_u10_u5_n135 ) , .ZN( u2_u10_u5_n142 ) );
  OAI21_X1 u2_u10_u5_U18 (.ZN( u2_u10_u5_n133 ) , .B2( u2_u10_u5_n147 ) , .A( u2_u10_u5_n173 ) , .B1( u2_u10_u5_n188 ) );
  NAND2_X1 u2_u10_u5_U19 (.A2( u2_u10_u5_n119 ) , .A1( u2_u10_u5_n123 ) , .ZN( u2_u10_u5_n137 ) );
  INV_X1 u2_u10_u5_U20 (.A( u2_u10_u5_n155 ) , .ZN( u2_u10_u5_n194 ) );
  NAND2_X1 u2_u10_u5_U21 (.A1( u2_u10_u5_n121 ) , .ZN( u2_u10_u5_n132 ) , .A2( u2_u10_u5_n172 ) );
  NAND2_X1 u2_u10_u5_U22 (.A2( u2_u10_u5_n122 ) , .ZN( u2_u10_u5_n136 ) , .A1( u2_u10_u5_n154 ) );
  NAND2_X1 u2_u10_u5_U23 (.A2( u2_u10_u5_n119 ) , .A1( u2_u10_u5_n120 ) , .ZN( u2_u10_u5_n159 ) );
  INV_X1 u2_u10_u5_U24 (.A( u2_u10_u5_n156 ) , .ZN( u2_u10_u5_n175 ) );
  INV_X1 u2_u10_u5_U25 (.A( u2_u10_u5_n158 ) , .ZN( u2_u10_u5_n188 ) );
  INV_X1 u2_u10_u5_U26 (.A( u2_u10_u5_n152 ) , .ZN( u2_u10_u5_n179 ) );
  INV_X1 u2_u10_u5_U27 (.A( u2_u10_u5_n140 ) , .ZN( u2_u10_u5_n182 ) );
  INV_X1 u2_u10_u5_U28 (.A( u2_u10_u5_n151 ) , .ZN( u2_u10_u5_n183 ) );
  INV_X1 u2_u10_u5_U29 (.A( u2_u10_u5_n123 ) , .ZN( u2_u10_u5_n185 ) );
  NOR2_X1 u2_u10_u5_U3 (.ZN( u2_u10_u5_n134 ) , .A1( u2_u10_u5_n183 ) , .A2( u2_u10_u5_n190 ) );
  INV_X1 u2_u10_u5_U30 (.A( u2_u10_u5_n161 ) , .ZN( u2_u10_u5_n184 ) );
  INV_X1 u2_u10_u5_U31 (.A( u2_u10_u5_n139 ) , .ZN( u2_u10_u5_n189 ) );
  INV_X1 u2_u10_u5_U32 (.A( u2_u10_u5_n157 ) , .ZN( u2_u10_u5_n190 ) );
  INV_X1 u2_u10_u5_U33 (.A( u2_u10_u5_n120 ) , .ZN( u2_u10_u5_n193 ) );
  NAND2_X1 u2_u10_u5_U34 (.ZN( u2_u10_u5_n111 ) , .A1( u2_u10_u5_n140 ) , .A2( u2_u10_u5_n155 ) );
  NOR2_X1 u2_u10_u5_U35 (.ZN( u2_u10_u5_n100 ) , .A1( u2_u10_u5_n170 ) , .A2( u2_u10_u5_n180 ) );
  INV_X1 u2_u10_u5_U36 (.A( u2_u10_u5_n117 ) , .ZN( u2_u10_u5_n196 ) );
  OAI221_X1 u2_u10_u5_U37 (.A( u2_u10_u5_n116 ) , .ZN( u2_u10_u5_n117 ) , .B2( u2_u10_u5_n119 ) , .C1( u2_u10_u5_n153 ) , .C2( u2_u10_u5_n158 ) , .B1( u2_u10_u5_n172 ) );
  AOI222_X1 u2_u10_u5_U38 (.ZN( u2_u10_u5_n116 ) , .B2( u2_u10_u5_n145 ) , .C1( u2_u10_u5_n148 ) , .A2( u2_u10_u5_n174 ) , .C2( u2_u10_u5_n177 ) , .B1( u2_u10_u5_n187 ) , .A1( u2_u10_u5_n193 ) );
  INV_X1 u2_u10_u5_U39 (.A( u2_u10_u5_n115 ) , .ZN( u2_u10_u5_n187 ) );
  INV_X1 u2_u10_u5_U4 (.A( u2_u10_u5_n138 ) , .ZN( u2_u10_u5_n191 ) );
  AOI22_X1 u2_u10_u5_U40 (.B2( u2_u10_u5_n131 ) , .A2( u2_u10_u5_n146 ) , .ZN( u2_u10_u5_n169 ) , .B1( u2_u10_u5_n174 ) , .A1( u2_u10_u5_n185 ) );
  NOR2_X1 u2_u10_u5_U41 (.A1( u2_u10_u5_n146 ) , .ZN( u2_u10_u5_n150 ) , .A2( u2_u10_u5_n173 ) );
  AOI21_X1 u2_u10_u5_U42 (.A( u2_u10_u5_n118 ) , .B2( u2_u10_u5_n145 ) , .ZN( u2_u10_u5_n168 ) , .B1( u2_u10_u5_n186 ) );
  INV_X1 u2_u10_u5_U43 (.A( u2_u10_u5_n122 ) , .ZN( u2_u10_u5_n186 ) );
  NOR2_X1 u2_u10_u5_U44 (.A1( u2_u10_u5_n146 ) , .ZN( u2_u10_u5_n152 ) , .A2( u2_u10_u5_n176 ) );
  NOR2_X1 u2_u10_u5_U45 (.A1( u2_u10_u5_n115 ) , .ZN( u2_u10_u5_n118 ) , .A2( u2_u10_u5_n153 ) );
  NOR2_X1 u2_u10_u5_U46 (.A2( u2_u10_u5_n145 ) , .ZN( u2_u10_u5_n156 ) , .A1( u2_u10_u5_n174 ) );
  NOR2_X1 u2_u10_u5_U47 (.ZN( u2_u10_u5_n121 ) , .A2( u2_u10_u5_n145 ) , .A1( u2_u10_u5_n176 ) );
  AOI22_X1 u2_u10_u5_U48 (.ZN( u2_u10_u5_n114 ) , .A2( u2_u10_u5_n137 ) , .A1( u2_u10_u5_n145 ) , .B2( u2_u10_u5_n175 ) , .B1( u2_u10_u5_n193 ) );
  OAI211_X1 u2_u10_u5_U49 (.B( u2_u10_u5_n124 ) , .A( u2_u10_u5_n125 ) , .C2( u2_u10_u5_n126 ) , .C1( u2_u10_u5_n127 ) , .ZN( u2_u10_u5_n128 ) );
  OAI21_X1 u2_u10_u5_U5 (.B2( u2_u10_u5_n136 ) , .B1( u2_u10_u5_n137 ) , .ZN( u2_u10_u5_n138 ) , .A( u2_u10_u5_n177 ) );
  NOR3_X1 u2_u10_u5_U50 (.ZN( u2_u10_u5_n127 ) , .A1( u2_u10_u5_n136 ) , .A3( u2_u10_u5_n148 ) , .A2( u2_u10_u5_n182 ) );
  OAI21_X1 u2_u10_u5_U51 (.ZN( u2_u10_u5_n124 ) , .A( u2_u10_u5_n177 ) , .B2( u2_u10_u5_n183 ) , .B1( u2_u10_u5_n189 ) );
  OAI21_X1 u2_u10_u5_U52 (.ZN( u2_u10_u5_n125 ) , .A( u2_u10_u5_n174 ) , .B2( u2_u10_u5_n185 ) , .B1( u2_u10_u5_n190 ) );
  AOI21_X1 u2_u10_u5_U53 (.A( u2_u10_u5_n153 ) , .B2( u2_u10_u5_n154 ) , .B1( u2_u10_u5_n155 ) , .ZN( u2_u10_u5_n164 ) );
  AOI21_X1 u2_u10_u5_U54 (.ZN( u2_u10_u5_n110 ) , .B1( u2_u10_u5_n122 ) , .B2( u2_u10_u5_n139 ) , .A( u2_u10_u5_n153 ) );
  INV_X1 u2_u10_u5_U55 (.A( u2_u10_u5_n153 ) , .ZN( u2_u10_u5_n176 ) );
  INV_X1 u2_u10_u5_U56 (.A( u2_u10_u5_n126 ) , .ZN( u2_u10_u5_n173 ) );
  AND2_X1 u2_u10_u5_U57 (.A2( u2_u10_u5_n104 ) , .A1( u2_u10_u5_n107 ) , .ZN( u2_u10_u5_n147 ) );
  AND2_X1 u2_u10_u5_U58 (.A2( u2_u10_u5_n104 ) , .A1( u2_u10_u5_n108 ) , .ZN( u2_u10_u5_n148 ) );
  NAND2_X1 u2_u10_u5_U59 (.A1( u2_u10_u5_n105 ) , .A2( u2_u10_u5_n106 ) , .ZN( u2_u10_u5_n158 ) );
  INV_X1 u2_u10_u5_U6 (.A( u2_u10_u5_n135 ) , .ZN( u2_u10_u5_n178 ) );
  NAND2_X1 u2_u10_u5_U60 (.A2( u2_u10_u5_n108 ) , .A1( u2_u10_u5_n109 ) , .ZN( u2_u10_u5_n139 ) );
  NAND2_X1 u2_u10_u5_U61 (.A1( u2_u10_u5_n106 ) , .A2( u2_u10_u5_n108 ) , .ZN( u2_u10_u5_n119 ) );
  NAND2_X1 u2_u10_u5_U62 (.A2( u2_u10_u5_n103 ) , .A1( u2_u10_u5_n105 ) , .ZN( u2_u10_u5_n140 ) );
  NAND2_X1 u2_u10_u5_U63 (.A2( u2_u10_u5_n104 ) , .A1( u2_u10_u5_n105 ) , .ZN( u2_u10_u5_n155 ) );
  NAND2_X1 u2_u10_u5_U64 (.A2( u2_u10_u5_n106 ) , .A1( u2_u10_u5_n107 ) , .ZN( u2_u10_u5_n122 ) );
  NAND2_X1 u2_u10_u5_U65 (.A2( u2_u10_u5_n100 ) , .A1( u2_u10_u5_n106 ) , .ZN( u2_u10_u5_n115 ) );
  NAND2_X1 u2_u10_u5_U66 (.A2( u2_u10_u5_n100 ) , .A1( u2_u10_u5_n103 ) , .ZN( u2_u10_u5_n161 ) );
  NAND2_X1 u2_u10_u5_U67 (.A1( u2_u10_u5_n105 ) , .A2( u2_u10_u5_n109 ) , .ZN( u2_u10_u5_n154 ) );
  INV_X1 u2_u10_u5_U68 (.A( u2_u10_u5_n146 ) , .ZN( u2_u10_u5_n172 ) );
  NAND2_X1 u2_u10_u5_U69 (.A1( u2_u10_u5_n103 ) , .A2( u2_u10_u5_n108 ) , .ZN( u2_u10_u5_n123 ) );
  OAI22_X1 u2_u10_u5_U7 (.B2( u2_u10_u5_n149 ) , .B1( u2_u10_u5_n150 ) , .A2( u2_u10_u5_n151 ) , .A1( u2_u10_u5_n152 ) , .ZN( u2_u10_u5_n165 ) );
  NAND2_X1 u2_u10_u5_U70 (.A2( u2_u10_u5_n103 ) , .A1( u2_u10_u5_n107 ) , .ZN( u2_u10_u5_n151 ) );
  NAND2_X1 u2_u10_u5_U71 (.A2( u2_u10_u5_n107 ) , .A1( u2_u10_u5_n109 ) , .ZN( u2_u10_u5_n120 ) );
  NAND2_X1 u2_u10_u5_U72 (.A2( u2_u10_u5_n100 ) , .A1( u2_u10_u5_n109 ) , .ZN( u2_u10_u5_n157 ) );
  AND2_X1 u2_u10_u5_U73 (.A2( u2_u10_u5_n100 ) , .A1( u2_u10_u5_n104 ) , .ZN( u2_u10_u5_n131 ) );
  INV_X1 u2_u10_u5_U74 (.A( u2_u10_u5_n102 ) , .ZN( u2_u10_u5_n195 ) );
  OAI221_X1 u2_u10_u5_U75 (.A( u2_u10_u5_n101 ) , .ZN( u2_u10_u5_n102 ) , .C2( u2_u10_u5_n115 ) , .C1( u2_u10_u5_n126 ) , .B1( u2_u10_u5_n134 ) , .B2( u2_u10_u5_n160 ) );
  OAI21_X1 u2_u10_u5_U76 (.ZN( u2_u10_u5_n101 ) , .B1( u2_u10_u5_n137 ) , .A( u2_u10_u5_n146 ) , .B2( u2_u10_u5_n147 ) );
  NOR2_X1 u2_u10_u5_U77 (.A2( u2_u10_X_34 ) , .A1( u2_u10_X_35 ) , .ZN( u2_u10_u5_n145 ) );
  NOR2_X1 u2_u10_u5_U78 (.A2( u2_u10_X_34 ) , .ZN( u2_u10_u5_n146 ) , .A1( u2_u10_u5_n171 ) );
  NOR2_X1 u2_u10_u5_U79 (.A2( u2_u10_X_31 ) , .A1( u2_u10_X_32 ) , .ZN( u2_u10_u5_n103 ) );
  NOR3_X1 u2_u10_u5_U8 (.A2( u2_u10_u5_n147 ) , .A1( u2_u10_u5_n148 ) , .ZN( u2_u10_u5_n149 ) , .A3( u2_u10_u5_n194 ) );
  NOR2_X1 u2_u10_u5_U80 (.A2( u2_u10_X_36 ) , .ZN( u2_u10_u5_n105 ) , .A1( u2_u10_u5_n180 ) );
  NOR2_X1 u2_u10_u5_U81 (.A2( u2_u10_X_33 ) , .ZN( u2_u10_u5_n108 ) , .A1( u2_u10_u5_n170 ) );
  NOR2_X1 u2_u10_u5_U82 (.A2( u2_u10_X_33 ) , .A1( u2_u10_X_36 ) , .ZN( u2_u10_u5_n107 ) );
  NOR2_X1 u2_u10_u5_U83 (.A2( u2_u10_X_31 ) , .ZN( u2_u10_u5_n104 ) , .A1( u2_u10_u5_n181 ) );
  NAND2_X1 u2_u10_u5_U84 (.A2( u2_u10_X_34 ) , .A1( u2_u10_X_35 ) , .ZN( u2_u10_u5_n153 ) );
  NAND2_X1 u2_u10_u5_U85 (.A1( u2_u10_X_34 ) , .ZN( u2_u10_u5_n126 ) , .A2( u2_u10_u5_n171 ) );
  AND2_X1 u2_u10_u5_U86 (.A1( u2_u10_X_31 ) , .A2( u2_u10_X_32 ) , .ZN( u2_u10_u5_n106 ) );
  AND2_X1 u2_u10_u5_U87 (.A1( u2_u10_X_31 ) , .ZN( u2_u10_u5_n109 ) , .A2( u2_u10_u5_n181 ) );
  INV_X1 u2_u10_u5_U88 (.A( u2_u10_X_33 ) , .ZN( u2_u10_u5_n180 ) );
  INV_X1 u2_u10_u5_U89 (.A( u2_u10_X_35 ) , .ZN( u2_u10_u5_n171 ) );
  NOR2_X1 u2_u10_u5_U9 (.ZN( u2_u10_u5_n135 ) , .A1( u2_u10_u5_n173 ) , .A2( u2_u10_u5_n176 ) );
  INV_X1 u2_u10_u5_U90 (.A( u2_u10_X_36 ) , .ZN( u2_u10_u5_n170 ) );
  INV_X1 u2_u10_u5_U91 (.A( u2_u10_X_32 ) , .ZN( u2_u10_u5_n181 ) );
  NAND4_X1 u2_u10_u5_U92 (.ZN( u2_out10_29 ) , .A4( u2_u10_u5_n129 ) , .A3( u2_u10_u5_n130 ) , .A2( u2_u10_u5_n168 ) , .A1( u2_u10_u5_n196 ) );
  AOI221_X1 u2_u10_u5_U93 (.A( u2_u10_u5_n128 ) , .ZN( u2_u10_u5_n129 ) , .C2( u2_u10_u5_n132 ) , .B2( u2_u10_u5_n159 ) , .B1( u2_u10_u5_n176 ) , .C1( u2_u10_u5_n184 ) );
  AOI222_X1 u2_u10_u5_U94 (.ZN( u2_u10_u5_n130 ) , .A2( u2_u10_u5_n146 ) , .B1( u2_u10_u5_n147 ) , .C2( u2_u10_u5_n175 ) , .B2( u2_u10_u5_n179 ) , .A1( u2_u10_u5_n188 ) , .C1( u2_u10_u5_n194 ) );
  NAND4_X1 u2_u10_u5_U95 (.ZN( u2_out10_19 ) , .A4( u2_u10_u5_n166 ) , .A3( u2_u10_u5_n167 ) , .A2( u2_u10_u5_n168 ) , .A1( u2_u10_u5_n169 ) );
  AOI22_X1 u2_u10_u5_U96 (.B2( u2_u10_u5_n145 ) , .A2( u2_u10_u5_n146 ) , .ZN( u2_u10_u5_n167 ) , .B1( u2_u10_u5_n182 ) , .A1( u2_u10_u5_n189 ) );
  NOR4_X1 u2_u10_u5_U97 (.A4( u2_u10_u5_n162 ) , .A3( u2_u10_u5_n163 ) , .A2( u2_u10_u5_n164 ) , .A1( u2_u10_u5_n165 ) , .ZN( u2_u10_u5_n166 ) );
  NAND4_X1 u2_u10_u5_U98 (.ZN( u2_out10_11 ) , .A4( u2_u10_u5_n143 ) , .A3( u2_u10_u5_n144 ) , .A2( u2_u10_u5_n169 ) , .A1( u2_u10_u5_n196 ) );
  AOI22_X1 u2_u10_u5_U99 (.A2( u2_u10_u5_n132 ) , .ZN( u2_u10_u5_n144 ) , .B2( u2_u10_u5_n145 ) , .B1( u2_u10_u5_n184 ) , .A1( u2_u10_u5_n194 ) );
  AOI22_X1 u2_u10_u6_U10 (.A2( u2_u10_u6_n151 ) , .B2( u2_u10_u6_n161 ) , .A1( u2_u10_u6_n167 ) , .B1( u2_u10_u6_n170 ) , .ZN( u2_u10_u6_n89 ) );
  AOI21_X1 u2_u10_u6_U11 (.B1( u2_u10_u6_n107 ) , .B2( u2_u10_u6_n132 ) , .A( u2_u10_u6_n158 ) , .ZN( u2_u10_u6_n88 ) );
  AOI21_X1 u2_u10_u6_U12 (.B2( u2_u10_u6_n147 ) , .B1( u2_u10_u6_n148 ) , .ZN( u2_u10_u6_n149 ) , .A( u2_u10_u6_n158 ) );
  AOI21_X1 u2_u10_u6_U13 (.ZN( u2_u10_u6_n106 ) , .A( u2_u10_u6_n142 ) , .B2( u2_u10_u6_n159 ) , .B1( u2_u10_u6_n164 ) );
  INV_X1 u2_u10_u6_U14 (.A( u2_u10_u6_n155 ) , .ZN( u2_u10_u6_n161 ) );
  INV_X1 u2_u10_u6_U15 (.A( u2_u10_u6_n128 ) , .ZN( u2_u10_u6_n164 ) );
  NAND2_X1 u2_u10_u6_U16 (.ZN( u2_u10_u6_n110 ) , .A1( u2_u10_u6_n122 ) , .A2( u2_u10_u6_n129 ) );
  NAND2_X1 u2_u10_u6_U17 (.ZN( u2_u10_u6_n124 ) , .A2( u2_u10_u6_n146 ) , .A1( u2_u10_u6_n148 ) );
  INV_X1 u2_u10_u6_U18 (.A( u2_u10_u6_n132 ) , .ZN( u2_u10_u6_n171 ) );
  AND2_X1 u2_u10_u6_U19 (.A1( u2_u10_u6_n100 ) , .ZN( u2_u10_u6_n130 ) , .A2( u2_u10_u6_n147 ) );
  INV_X1 u2_u10_u6_U20 (.A( u2_u10_u6_n127 ) , .ZN( u2_u10_u6_n173 ) );
  INV_X1 u2_u10_u6_U21 (.A( u2_u10_u6_n121 ) , .ZN( u2_u10_u6_n167 ) );
  INV_X1 u2_u10_u6_U22 (.A( u2_u10_u6_n100 ) , .ZN( u2_u10_u6_n169 ) );
  INV_X1 u2_u10_u6_U23 (.A( u2_u10_u6_n123 ) , .ZN( u2_u10_u6_n170 ) );
  INV_X1 u2_u10_u6_U24 (.A( u2_u10_u6_n113 ) , .ZN( u2_u10_u6_n168 ) );
  AND2_X1 u2_u10_u6_U25 (.A1( u2_u10_u6_n107 ) , .A2( u2_u10_u6_n119 ) , .ZN( u2_u10_u6_n133 ) );
  AND2_X1 u2_u10_u6_U26 (.A2( u2_u10_u6_n121 ) , .A1( u2_u10_u6_n122 ) , .ZN( u2_u10_u6_n131 ) );
  AND3_X1 u2_u10_u6_U27 (.ZN( u2_u10_u6_n120 ) , .A2( u2_u10_u6_n127 ) , .A1( u2_u10_u6_n132 ) , .A3( u2_u10_u6_n145 ) );
  INV_X1 u2_u10_u6_U28 (.A( u2_u10_u6_n146 ) , .ZN( u2_u10_u6_n163 ) );
  AOI222_X1 u2_u10_u6_U29 (.ZN( u2_u10_u6_n114 ) , .A1( u2_u10_u6_n118 ) , .A2( u2_u10_u6_n126 ) , .B2( u2_u10_u6_n151 ) , .C2( u2_u10_u6_n159 ) , .C1( u2_u10_u6_n168 ) , .B1( u2_u10_u6_n169 ) );
  INV_X1 u2_u10_u6_U3 (.A( u2_u10_u6_n110 ) , .ZN( u2_u10_u6_n166 ) );
  NOR2_X1 u2_u10_u6_U30 (.A1( u2_u10_u6_n162 ) , .A2( u2_u10_u6_n165 ) , .ZN( u2_u10_u6_n98 ) );
  AOI211_X1 u2_u10_u6_U31 (.B( u2_u10_u6_n134 ) , .A( u2_u10_u6_n135 ) , .C1( u2_u10_u6_n136 ) , .ZN( u2_u10_u6_n137 ) , .C2( u2_u10_u6_n151 ) );
  NAND4_X1 u2_u10_u6_U32 (.A4( u2_u10_u6_n127 ) , .A3( u2_u10_u6_n128 ) , .A2( u2_u10_u6_n129 ) , .A1( u2_u10_u6_n130 ) , .ZN( u2_u10_u6_n136 ) );
  AOI21_X1 u2_u10_u6_U33 (.B2( u2_u10_u6_n132 ) , .B1( u2_u10_u6_n133 ) , .ZN( u2_u10_u6_n134 ) , .A( u2_u10_u6_n158 ) );
  AOI21_X1 u2_u10_u6_U34 (.B1( u2_u10_u6_n131 ) , .ZN( u2_u10_u6_n135 ) , .A( u2_u10_u6_n144 ) , .B2( u2_u10_u6_n146 ) );
  NAND2_X1 u2_u10_u6_U35 (.A1( u2_u10_u6_n144 ) , .ZN( u2_u10_u6_n151 ) , .A2( u2_u10_u6_n158 ) );
  NAND2_X1 u2_u10_u6_U36 (.ZN( u2_u10_u6_n132 ) , .A1( u2_u10_u6_n91 ) , .A2( u2_u10_u6_n97 ) );
  AOI22_X1 u2_u10_u6_U37 (.B2( u2_u10_u6_n110 ) , .B1( u2_u10_u6_n111 ) , .A1( u2_u10_u6_n112 ) , .ZN( u2_u10_u6_n115 ) , .A2( u2_u10_u6_n161 ) );
  NAND4_X1 u2_u10_u6_U38 (.A3( u2_u10_u6_n109 ) , .ZN( u2_u10_u6_n112 ) , .A4( u2_u10_u6_n132 ) , .A2( u2_u10_u6_n147 ) , .A1( u2_u10_u6_n166 ) );
  NOR2_X1 u2_u10_u6_U39 (.ZN( u2_u10_u6_n109 ) , .A1( u2_u10_u6_n170 ) , .A2( u2_u10_u6_n173 ) );
  INV_X1 u2_u10_u6_U4 (.A( u2_u10_u6_n142 ) , .ZN( u2_u10_u6_n174 ) );
  NOR2_X1 u2_u10_u6_U40 (.A2( u2_u10_u6_n126 ) , .ZN( u2_u10_u6_n155 ) , .A1( u2_u10_u6_n160 ) );
  NAND2_X1 u2_u10_u6_U41 (.ZN( u2_u10_u6_n146 ) , .A2( u2_u10_u6_n94 ) , .A1( u2_u10_u6_n99 ) );
  AOI21_X1 u2_u10_u6_U42 (.A( u2_u10_u6_n144 ) , .B2( u2_u10_u6_n145 ) , .B1( u2_u10_u6_n146 ) , .ZN( u2_u10_u6_n150 ) );
  INV_X1 u2_u10_u6_U43 (.A( u2_u10_u6_n111 ) , .ZN( u2_u10_u6_n158 ) );
  NAND2_X1 u2_u10_u6_U44 (.ZN( u2_u10_u6_n127 ) , .A1( u2_u10_u6_n91 ) , .A2( u2_u10_u6_n92 ) );
  NAND2_X1 u2_u10_u6_U45 (.ZN( u2_u10_u6_n129 ) , .A2( u2_u10_u6_n95 ) , .A1( u2_u10_u6_n96 ) );
  INV_X1 u2_u10_u6_U46 (.A( u2_u10_u6_n144 ) , .ZN( u2_u10_u6_n159 ) );
  NAND2_X1 u2_u10_u6_U47 (.ZN( u2_u10_u6_n145 ) , .A2( u2_u10_u6_n97 ) , .A1( u2_u10_u6_n98 ) );
  NAND2_X1 u2_u10_u6_U48 (.ZN( u2_u10_u6_n148 ) , .A2( u2_u10_u6_n92 ) , .A1( u2_u10_u6_n94 ) );
  NAND2_X1 u2_u10_u6_U49 (.ZN( u2_u10_u6_n108 ) , .A2( u2_u10_u6_n139 ) , .A1( u2_u10_u6_n144 ) );
  NAND2_X1 u2_u10_u6_U5 (.A2( u2_u10_u6_n143 ) , .ZN( u2_u10_u6_n152 ) , .A1( u2_u10_u6_n166 ) );
  NAND2_X1 u2_u10_u6_U50 (.ZN( u2_u10_u6_n121 ) , .A2( u2_u10_u6_n95 ) , .A1( u2_u10_u6_n97 ) );
  NAND2_X1 u2_u10_u6_U51 (.ZN( u2_u10_u6_n107 ) , .A2( u2_u10_u6_n92 ) , .A1( u2_u10_u6_n95 ) );
  AND2_X1 u2_u10_u6_U52 (.ZN( u2_u10_u6_n118 ) , .A2( u2_u10_u6_n91 ) , .A1( u2_u10_u6_n99 ) );
  NAND2_X1 u2_u10_u6_U53 (.ZN( u2_u10_u6_n147 ) , .A2( u2_u10_u6_n98 ) , .A1( u2_u10_u6_n99 ) );
  NAND2_X1 u2_u10_u6_U54 (.ZN( u2_u10_u6_n128 ) , .A1( u2_u10_u6_n94 ) , .A2( u2_u10_u6_n96 ) );
  NAND2_X1 u2_u10_u6_U55 (.ZN( u2_u10_u6_n119 ) , .A2( u2_u10_u6_n95 ) , .A1( u2_u10_u6_n99 ) );
  NAND2_X1 u2_u10_u6_U56 (.ZN( u2_u10_u6_n123 ) , .A2( u2_u10_u6_n91 ) , .A1( u2_u10_u6_n96 ) );
  NAND2_X1 u2_u10_u6_U57 (.ZN( u2_u10_u6_n100 ) , .A2( u2_u10_u6_n92 ) , .A1( u2_u10_u6_n98 ) );
  NAND2_X1 u2_u10_u6_U58 (.ZN( u2_u10_u6_n122 ) , .A1( u2_u10_u6_n94 ) , .A2( u2_u10_u6_n97 ) );
  INV_X1 u2_u10_u6_U59 (.A( u2_u10_u6_n139 ) , .ZN( u2_u10_u6_n160 ) );
  AOI22_X1 u2_u10_u6_U6 (.B2( u2_u10_u6_n101 ) , .A1( u2_u10_u6_n102 ) , .ZN( u2_u10_u6_n103 ) , .B1( u2_u10_u6_n160 ) , .A2( u2_u10_u6_n161 ) );
  NAND2_X1 u2_u10_u6_U60 (.ZN( u2_u10_u6_n113 ) , .A1( u2_u10_u6_n96 ) , .A2( u2_u10_u6_n98 ) );
  NOR2_X1 u2_u10_u6_U61 (.A2( u2_u10_X_40 ) , .A1( u2_u10_X_41 ) , .ZN( u2_u10_u6_n126 ) );
  NOR2_X1 u2_u10_u6_U62 (.A2( u2_u10_X_39 ) , .A1( u2_u10_X_42 ) , .ZN( u2_u10_u6_n92 ) );
  NOR2_X1 u2_u10_u6_U63 (.A2( u2_u10_X_39 ) , .A1( u2_u10_u6_n156 ) , .ZN( u2_u10_u6_n97 ) );
  NOR2_X1 u2_u10_u6_U64 (.A2( u2_u10_X_38 ) , .A1( u2_u10_u6_n165 ) , .ZN( u2_u10_u6_n95 ) );
  NOR2_X1 u2_u10_u6_U65 (.A2( u2_u10_X_41 ) , .ZN( u2_u10_u6_n111 ) , .A1( u2_u10_u6_n157 ) );
  NOR2_X1 u2_u10_u6_U66 (.A2( u2_u10_X_37 ) , .A1( u2_u10_u6_n162 ) , .ZN( u2_u10_u6_n94 ) );
  NOR2_X1 u2_u10_u6_U67 (.A2( u2_u10_X_37 ) , .A1( u2_u10_X_38 ) , .ZN( u2_u10_u6_n91 ) );
  NAND2_X1 u2_u10_u6_U68 (.A1( u2_u10_X_41 ) , .ZN( u2_u10_u6_n144 ) , .A2( u2_u10_u6_n157 ) );
  NAND2_X1 u2_u10_u6_U69 (.A2( u2_u10_X_40 ) , .A1( u2_u10_X_41 ) , .ZN( u2_u10_u6_n139 ) );
  NOR2_X1 u2_u10_u6_U7 (.A1( u2_u10_u6_n118 ) , .ZN( u2_u10_u6_n143 ) , .A2( u2_u10_u6_n168 ) );
  AND2_X1 u2_u10_u6_U70 (.A1( u2_u10_X_39 ) , .A2( u2_u10_u6_n156 ) , .ZN( u2_u10_u6_n96 ) );
  AND2_X1 u2_u10_u6_U71 (.A1( u2_u10_X_39 ) , .A2( u2_u10_X_42 ) , .ZN( u2_u10_u6_n99 ) );
  INV_X1 u2_u10_u6_U72 (.A( u2_u10_X_40 ) , .ZN( u2_u10_u6_n157 ) );
  INV_X1 u2_u10_u6_U73 (.A( u2_u10_X_37 ) , .ZN( u2_u10_u6_n165 ) );
  INV_X1 u2_u10_u6_U74 (.A( u2_u10_X_38 ) , .ZN( u2_u10_u6_n162 ) );
  INV_X1 u2_u10_u6_U75 (.A( u2_u10_X_42 ) , .ZN( u2_u10_u6_n156 ) );
  NAND4_X1 u2_u10_u6_U76 (.ZN( u2_out10_12 ) , .A4( u2_u10_u6_n114 ) , .A3( u2_u10_u6_n115 ) , .A2( u2_u10_u6_n116 ) , .A1( u2_u10_u6_n117 ) );
  OAI22_X1 u2_u10_u6_U77 (.B2( u2_u10_u6_n111 ) , .ZN( u2_u10_u6_n116 ) , .B1( u2_u10_u6_n126 ) , .A2( u2_u10_u6_n164 ) , .A1( u2_u10_u6_n167 ) );
  OAI21_X1 u2_u10_u6_U78 (.A( u2_u10_u6_n108 ) , .ZN( u2_u10_u6_n117 ) , .B2( u2_u10_u6_n141 ) , .B1( u2_u10_u6_n163 ) );
  NAND4_X1 u2_u10_u6_U79 (.ZN( u2_out10_32 ) , .A4( u2_u10_u6_n103 ) , .A3( u2_u10_u6_n104 ) , .A2( u2_u10_u6_n105 ) , .A1( u2_u10_u6_n106 ) );
  INV_X1 u2_u10_u6_U8 (.ZN( u2_u10_u6_n172 ) , .A( u2_u10_u6_n88 ) );
  AOI22_X1 u2_u10_u6_U80 (.ZN( u2_u10_u6_n105 ) , .A2( u2_u10_u6_n108 ) , .A1( u2_u10_u6_n118 ) , .B2( u2_u10_u6_n126 ) , .B1( u2_u10_u6_n171 ) );
  AOI22_X1 u2_u10_u6_U81 (.ZN( u2_u10_u6_n104 ) , .A1( u2_u10_u6_n111 ) , .B1( u2_u10_u6_n124 ) , .B2( u2_u10_u6_n151 ) , .A2( u2_u10_u6_n93 ) );
  OAI211_X1 u2_u10_u6_U82 (.ZN( u2_out10_7 ) , .B( u2_u10_u6_n153 ) , .C2( u2_u10_u6_n154 ) , .C1( u2_u10_u6_n155 ) , .A( u2_u10_u6_n174 ) );
  NOR3_X1 u2_u10_u6_U83 (.A1( u2_u10_u6_n141 ) , .ZN( u2_u10_u6_n154 ) , .A3( u2_u10_u6_n164 ) , .A2( u2_u10_u6_n171 ) );
  AOI211_X1 u2_u10_u6_U84 (.B( u2_u10_u6_n149 ) , .A( u2_u10_u6_n150 ) , .C2( u2_u10_u6_n151 ) , .C1( u2_u10_u6_n152 ) , .ZN( u2_u10_u6_n153 ) );
  OAI211_X1 u2_u10_u6_U85 (.ZN( u2_out10_22 ) , .B( u2_u10_u6_n137 ) , .A( u2_u10_u6_n138 ) , .C2( u2_u10_u6_n139 ) , .C1( u2_u10_u6_n140 ) );
  AOI22_X1 u2_u10_u6_U86 (.B1( u2_u10_u6_n124 ) , .A2( u2_u10_u6_n125 ) , .A1( u2_u10_u6_n126 ) , .ZN( u2_u10_u6_n138 ) , .B2( u2_u10_u6_n161 ) );
  AND4_X1 u2_u10_u6_U87 (.A3( u2_u10_u6_n119 ) , .A1( u2_u10_u6_n120 ) , .A4( u2_u10_u6_n129 ) , .ZN( u2_u10_u6_n140 ) , .A2( u2_u10_u6_n143 ) );
  NAND3_X1 u2_u10_u6_U88 (.A2( u2_u10_u6_n123 ) , .ZN( u2_u10_u6_n125 ) , .A1( u2_u10_u6_n130 ) , .A3( u2_u10_u6_n131 ) );
  NAND3_X1 u2_u10_u6_U89 (.A3( u2_u10_u6_n133 ) , .ZN( u2_u10_u6_n141 ) , .A1( u2_u10_u6_n145 ) , .A2( u2_u10_u6_n148 ) );
  OAI21_X1 u2_u10_u6_U9 (.A( u2_u10_u6_n159 ) , .B1( u2_u10_u6_n169 ) , .B2( u2_u10_u6_n173 ) , .ZN( u2_u10_u6_n90 ) );
  NAND3_X1 u2_u10_u6_U90 (.ZN( u2_u10_u6_n101 ) , .A3( u2_u10_u6_n107 ) , .A2( u2_u10_u6_n121 ) , .A1( u2_u10_u6_n127 ) );
  NAND3_X1 u2_u10_u6_U91 (.ZN( u2_u10_u6_n102 ) , .A3( u2_u10_u6_n130 ) , .A2( u2_u10_u6_n145 ) , .A1( u2_u10_u6_n166 ) );
  NAND3_X1 u2_u10_u6_U92 (.A3( u2_u10_u6_n113 ) , .A1( u2_u10_u6_n119 ) , .A2( u2_u10_u6_n123 ) , .ZN( u2_u10_u6_n93 ) );
  NAND3_X1 u2_u10_u6_U93 (.ZN( u2_u10_u6_n142 ) , .A2( u2_u10_u6_n172 ) , .A3( u2_u10_u6_n89 ) , .A1( u2_u10_u6_n90 ) );
  AND3_X1 u2_u10_u7_U10 (.A3( u2_u10_u7_n110 ) , .A2( u2_u10_u7_n127 ) , .A1( u2_u10_u7_n132 ) , .ZN( u2_u10_u7_n92 ) );
  OAI21_X1 u2_u10_u7_U11 (.A( u2_u10_u7_n161 ) , .B1( u2_u10_u7_n168 ) , .B2( u2_u10_u7_n173 ) , .ZN( u2_u10_u7_n91 ) );
  AOI211_X1 u2_u10_u7_U12 (.A( u2_u10_u7_n117 ) , .ZN( u2_u10_u7_n118 ) , .C2( u2_u10_u7_n126 ) , .C1( u2_u10_u7_n177 ) , .B( u2_u10_u7_n180 ) );
  OAI22_X1 u2_u10_u7_U13 (.B1( u2_u10_u7_n115 ) , .ZN( u2_u10_u7_n117 ) , .A2( u2_u10_u7_n133 ) , .A1( u2_u10_u7_n137 ) , .B2( u2_u10_u7_n162 ) );
  INV_X1 u2_u10_u7_U14 (.A( u2_u10_u7_n116 ) , .ZN( u2_u10_u7_n180 ) );
  NOR3_X1 u2_u10_u7_U15 (.ZN( u2_u10_u7_n115 ) , .A3( u2_u10_u7_n145 ) , .A2( u2_u10_u7_n168 ) , .A1( u2_u10_u7_n169 ) );
  OAI211_X1 u2_u10_u7_U16 (.B( u2_u10_u7_n122 ) , .A( u2_u10_u7_n123 ) , .C2( u2_u10_u7_n124 ) , .ZN( u2_u10_u7_n154 ) , .C1( u2_u10_u7_n162 ) );
  AOI222_X1 u2_u10_u7_U17 (.ZN( u2_u10_u7_n122 ) , .C2( u2_u10_u7_n126 ) , .C1( u2_u10_u7_n145 ) , .B1( u2_u10_u7_n161 ) , .A2( u2_u10_u7_n165 ) , .B2( u2_u10_u7_n170 ) , .A1( u2_u10_u7_n176 ) );
  INV_X1 u2_u10_u7_U18 (.A( u2_u10_u7_n133 ) , .ZN( u2_u10_u7_n176 ) );
  NOR3_X1 u2_u10_u7_U19 (.A2( u2_u10_u7_n134 ) , .A1( u2_u10_u7_n135 ) , .ZN( u2_u10_u7_n136 ) , .A3( u2_u10_u7_n171 ) );
  NOR2_X1 u2_u10_u7_U20 (.A1( u2_u10_u7_n130 ) , .A2( u2_u10_u7_n134 ) , .ZN( u2_u10_u7_n153 ) );
  INV_X1 u2_u10_u7_U21 (.A( u2_u10_u7_n101 ) , .ZN( u2_u10_u7_n165 ) );
  NOR2_X1 u2_u10_u7_U22 (.ZN( u2_u10_u7_n111 ) , .A2( u2_u10_u7_n134 ) , .A1( u2_u10_u7_n169 ) );
  AOI21_X1 u2_u10_u7_U23 (.ZN( u2_u10_u7_n104 ) , .B2( u2_u10_u7_n112 ) , .B1( u2_u10_u7_n127 ) , .A( u2_u10_u7_n164 ) );
  AOI21_X1 u2_u10_u7_U24 (.ZN( u2_u10_u7_n106 ) , .B1( u2_u10_u7_n133 ) , .B2( u2_u10_u7_n146 ) , .A( u2_u10_u7_n162 ) );
  AOI21_X1 u2_u10_u7_U25 (.A( u2_u10_u7_n101 ) , .ZN( u2_u10_u7_n107 ) , .B2( u2_u10_u7_n128 ) , .B1( u2_u10_u7_n175 ) );
  INV_X1 u2_u10_u7_U26 (.A( u2_u10_u7_n138 ) , .ZN( u2_u10_u7_n171 ) );
  INV_X1 u2_u10_u7_U27 (.A( u2_u10_u7_n131 ) , .ZN( u2_u10_u7_n177 ) );
  INV_X1 u2_u10_u7_U28 (.A( u2_u10_u7_n110 ) , .ZN( u2_u10_u7_n174 ) );
  NAND2_X1 u2_u10_u7_U29 (.A1( u2_u10_u7_n129 ) , .A2( u2_u10_u7_n132 ) , .ZN( u2_u10_u7_n149 ) );
  OAI21_X1 u2_u10_u7_U3 (.ZN( u2_u10_u7_n159 ) , .A( u2_u10_u7_n165 ) , .B2( u2_u10_u7_n171 ) , .B1( u2_u10_u7_n174 ) );
  NAND2_X1 u2_u10_u7_U30 (.A1( u2_u10_u7_n113 ) , .A2( u2_u10_u7_n124 ) , .ZN( u2_u10_u7_n130 ) );
  INV_X1 u2_u10_u7_U31 (.A( u2_u10_u7_n112 ) , .ZN( u2_u10_u7_n173 ) );
  INV_X1 u2_u10_u7_U32 (.A( u2_u10_u7_n128 ) , .ZN( u2_u10_u7_n168 ) );
  INV_X1 u2_u10_u7_U33 (.A( u2_u10_u7_n148 ) , .ZN( u2_u10_u7_n169 ) );
  INV_X1 u2_u10_u7_U34 (.A( u2_u10_u7_n127 ) , .ZN( u2_u10_u7_n179 ) );
  NOR2_X1 u2_u10_u7_U35 (.ZN( u2_u10_u7_n101 ) , .A2( u2_u10_u7_n150 ) , .A1( u2_u10_u7_n156 ) );
  AOI211_X1 u2_u10_u7_U36 (.B( u2_u10_u7_n154 ) , .A( u2_u10_u7_n155 ) , .C1( u2_u10_u7_n156 ) , .ZN( u2_u10_u7_n157 ) , .C2( u2_u10_u7_n172 ) );
  INV_X1 u2_u10_u7_U37 (.A( u2_u10_u7_n153 ) , .ZN( u2_u10_u7_n172 ) );
  AOI211_X1 u2_u10_u7_U38 (.B( u2_u10_u7_n139 ) , .A( u2_u10_u7_n140 ) , .C2( u2_u10_u7_n141 ) , .ZN( u2_u10_u7_n142 ) , .C1( u2_u10_u7_n156 ) );
  NAND4_X1 u2_u10_u7_U39 (.A3( u2_u10_u7_n127 ) , .A2( u2_u10_u7_n128 ) , .A1( u2_u10_u7_n129 ) , .ZN( u2_u10_u7_n141 ) , .A4( u2_u10_u7_n147 ) );
  INV_X1 u2_u10_u7_U4 (.A( u2_u10_u7_n111 ) , .ZN( u2_u10_u7_n170 ) );
  AOI21_X1 u2_u10_u7_U40 (.A( u2_u10_u7_n137 ) , .B1( u2_u10_u7_n138 ) , .ZN( u2_u10_u7_n139 ) , .B2( u2_u10_u7_n146 ) );
  OAI22_X1 u2_u10_u7_U41 (.B1( u2_u10_u7_n136 ) , .ZN( u2_u10_u7_n140 ) , .A1( u2_u10_u7_n153 ) , .B2( u2_u10_u7_n162 ) , .A2( u2_u10_u7_n164 ) );
  AOI21_X1 u2_u10_u7_U42 (.ZN( u2_u10_u7_n123 ) , .B1( u2_u10_u7_n165 ) , .B2( u2_u10_u7_n177 ) , .A( u2_u10_u7_n97 ) );
  AOI21_X1 u2_u10_u7_U43 (.B2( u2_u10_u7_n113 ) , .B1( u2_u10_u7_n124 ) , .A( u2_u10_u7_n125 ) , .ZN( u2_u10_u7_n97 ) );
  INV_X1 u2_u10_u7_U44 (.A( u2_u10_u7_n125 ) , .ZN( u2_u10_u7_n161 ) );
  INV_X1 u2_u10_u7_U45 (.A( u2_u10_u7_n152 ) , .ZN( u2_u10_u7_n162 ) );
  AOI22_X1 u2_u10_u7_U46 (.A2( u2_u10_u7_n114 ) , .ZN( u2_u10_u7_n119 ) , .B1( u2_u10_u7_n130 ) , .A1( u2_u10_u7_n156 ) , .B2( u2_u10_u7_n165 ) );
  NAND2_X1 u2_u10_u7_U47 (.A2( u2_u10_u7_n112 ) , .ZN( u2_u10_u7_n114 ) , .A1( u2_u10_u7_n175 ) );
  AND2_X1 u2_u10_u7_U48 (.ZN( u2_u10_u7_n145 ) , .A2( u2_u10_u7_n98 ) , .A1( u2_u10_u7_n99 ) );
  NOR2_X1 u2_u10_u7_U49 (.ZN( u2_u10_u7_n137 ) , .A1( u2_u10_u7_n150 ) , .A2( u2_u10_u7_n161 ) );
  INV_X1 u2_u10_u7_U5 (.A( u2_u10_u7_n149 ) , .ZN( u2_u10_u7_n175 ) );
  AOI21_X1 u2_u10_u7_U50 (.ZN( u2_u10_u7_n105 ) , .B2( u2_u10_u7_n110 ) , .A( u2_u10_u7_n125 ) , .B1( u2_u10_u7_n147 ) );
  NAND2_X1 u2_u10_u7_U51 (.ZN( u2_u10_u7_n146 ) , .A1( u2_u10_u7_n95 ) , .A2( u2_u10_u7_n98 ) );
  NAND2_X1 u2_u10_u7_U52 (.A2( u2_u10_u7_n103 ) , .ZN( u2_u10_u7_n147 ) , .A1( u2_u10_u7_n93 ) );
  NAND2_X1 u2_u10_u7_U53 (.A1( u2_u10_u7_n103 ) , .ZN( u2_u10_u7_n127 ) , .A2( u2_u10_u7_n99 ) );
  OR2_X1 u2_u10_u7_U54 (.ZN( u2_u10_u7_n126 ) , .A2( u2_u10_u7_n152 ) , .A1( u2_u10_u7_n156 ) );
  NAND2_X1 u2_u10_u7_U55 (.A2( u2_u10_u7_n102 ) , .A1( u2_u10_u7_n103 ) , .ZN( u2_u10_u7_n133 ) );
  NAND2_X1 u2_u10_u7_U56 (.ZN( u2_u10_u7_n112 ) , .A2( u2_u10_u7_n96 ) , .A1( u2_u10_u7_n99 ) );
  NAND2_X1 u2_u10_u7_U57 (.A2( u2_u10_u7_n102 ) , .ZN( u2_u10_u7_n128 ) , .A1( u2_u10_u7_n98 ) );
  NAND2_X1 u2_u10_u7_U58 (.A1( u2_u10_u7_n100 ) , .ZN( u2_u10_u7_n113 ) , .A2( u2_u10_u7_n93 ) );
  NAND2_X1 u2_u10_u7_U59 (.A2( u2_u10_u7_n102 ) , .ZN( u2_u10_u7_n124 ) , .A1( u2_u10_u7_n96 ) );
  INV_X1 u2_u10_u7_U6 (.A( u2_u10_u7_n154 ) , .ZN( u2_u10_u7_n178 ) );
  NAND2_X1 u2_u10_u7_U60 (.ZN( u2_u10_u7_n110 ) , .A1( u2_u10_u7_n95 ) , .A2( u2_u10_u7_n96 ) );
  INV_X1 u2_u10_u7_U61 (.A( u2_u10_u7_n150 ) , .ZN( u2_u10_u7_n164 ) );
  AND2_X1 u2_u10_u7_U62 (.ZN( u2_u10_u7_n134 ) , .A1( u2_u10_u7_n93 ) , .A2( u2_u10_u7_n98 ) );
  NAND2_X1 u2_u10_u7_U63 (.A1( u2_u10_u7_n100 ) , .A2( u2_u10_u7_n102 ) , .ZN( u2_u10_u7_n129 ) );
  NAND2_X1 u2_u10_u7_U64 (.A2( u2_u10_u7_n103 ) , .ZN( u2_u10_u7_n131 ) , .A1( u2_u10_u7_n95 ) );
  NAND2_X1 u2_u10_u7_U65 (.A1( u2_u10_u7_n100 ) , .ZN( u2_u10_u7_n138 ) , .A2( u2_u10_u7_n99 ) );
  NAND2_X1 u2_u10_u7_U66 (.ZN( u2_u10_u7_n132 ) , .A1( u2_u10_u7_n93 ) , .A2( u2_u10_u7_n96 ) );
  NAND2_X1 u2_u10_u7_U67 (.A1( u2_u10_u7_n100 ) , .ZN( u2_u10_u7_n148 ) , .A2( u2_u10_u7_n95 ) );
  NOR2_X1 u2_u10_u7_U68 (.A2( u2_u10_X_47 ) , .ZN( u2_u10_u7_n150 ) , .A1( u2_u10_u7_n163 ) );
  NOR2_X1 u2_u10_u7_U69 (.A2( u2_u10_X_43 ) , .A1( u2_u10_X_44 ) , .ZN( u2_u10_u7_n103 ) );
  AOI211_X1 u2_u10_u7_U7 (.ZN( u2_u10_u7_n116 ) , .A( u2_u10_u7_n155 ) , .C1( u2_u10_u7_n161 ) , .C2( u2_u10_u7_n171 ) , .B( u2_u10_u7_n94 ) );
  NOR2_X1 u2_u10_u7_U70 (.A2( u2_u10_X_48 ) , .A1( u2_u10_u7_n166 ) , .ZN( u2_u10_u7_n95 ) );
  NOR2_X1 u2_u10_u7_U71 (.A2( u2_u10_X_45 ) , .A1( u2_u10_X_48 ) , .ZN( u2_u10_u7_n99 ) );
  NOR2_X1 u2_u10_u7_U72 (.A2( u2_u10_X_44 ) , .A1( u2_u10_u7_n167 ) , .ZN( u2_u10_u7_n98 ) );
  NOR2_X1 u2_u10_u7_U73 (.A2( u2_u10_X_46 ) , .A1( u2_u10_X_47 ) , .ZN( u2_u10_u7_n152 ) );
  AND2_X1 u2_u10_u7_U74 (.A1( u2_u10_X_47 ) , .ZN( u2_u10_u7_n156 ) , .A2( u2_u10_u7_n163 ) );
  NAND2_X1 u2_u10_u7_U75 (.A2( u2_u10_X_46 ) , .A1( u2_u10_X_47 ) , .ZN( u2_u10_u7_n125 ) );
  AND2_X1 u2_u10_u7_U76 (.A2( u2_u10_X_45 ) , .A1( u2_u10_X_48 ) , .ZN( u2_u10_u7_n102 ) );
  AND2_X1 u2_u10_u7_U77 (.A2( u2_u10_X_43 ) , .A1( u2_u10_X_44 ) , .ZN( u2_u10_u7_n96 ) );
  AND2_X1 u2_u10_u7_U78 (.A1( u2_u10_X_44 ) , .ZN( u2_u10_u7_n100 ) , .A2( u2_u10_u7_n167 ) );
  AND2_X1 u2_u10_u7_U79 (.A1( u2_u10_X_48 ) , .A2( u2_u10_u7_n166 ) , .ZN( u2_u10_u7_n93 ) );
  OAI222_X1 u2_u10_u7_U8 (.C2( u2_u10_u7_n101 ) , .B2( u2_u10_u7_n111 ) , .A1( u2_u10_u7_n113 ) , .C1( u2_u10_u7_n146 ) , .A2( u2_u10_u7_n162 ) , .B1( u2_u10_u7_n164 ) , .ZN( u2_u10_u7_n94 ) );
  INV_X1 u2_u10_u7_U80 (.A( u2_u10_X_46 ) , .ZN( u2_u10_u7_n163 ) );
  INV_X1 u2_u10_u7_U81 (.A( u2_u10_X_43 ) , .ZN( u2_u10_u7_n167 ) );
  INV_X1 u2_u10_u7_U82 (.A( u2_u10_X_45 ) , .ZN( u2_u10_u7_n166 ) );
  NAND4_X1 u2_u10_u7_U83 (.ZN( u2_out10_27 ) , .A4( u2_u10_u7_n118 ) , .A3( u2_u10_u7_n119 ) , .A2( u2_u10_u7_n120 ) , .A1( u2_u10_u7_n121 ) );
  OAI21_X1 u2_u10_u7_U84 (.ZN( u2_u10_u7_n121 ) , .B2( u2_u10_u7_n145 ) , .A( u2_u10_u7_n150 ) , .B1( u2_u10_u7_n174 ) );
  OAI21_X1 u2_u10_u7_U85 (.ZN( u2_u10_u7_n120 ) , .A( u2_u10_u7_n161 ) , .B2( u2_u10_u7_n170 ) , .B1( u2_u10_u7_n179 ) );
  NAND4_X1 u2_u10_u7_U86 (.ZN( u2_out10_21 ) , .A4( u2_u10_u7_n157 ) , .A3( u2_u10_u7_n158 ) , .A2( u2_u10_u7_n159 ) , .A1( u2_u10_u7_n160 ) );
  OAI21_X1 u2_u10_u7_U87 (.B1( u2_u10_u7_n145 ) , .ZN( u2_u10_u7_n160 ) , .A( u2_u10_u7_n161 ) , .B2( u2_u10_u7_n177 ) );
  AOI22_X1 u2_u10_u7_U88 (.B2( u2_u10_u7_n149 ) , .B1( u2_u10_u7_n150 ) , .A2( u2_u10_u7_n151 ) , .A1( u2_u10_u7_n152 ) , .ZN( u2_u10_u7_n158 ) );
  NAND4_X1 u2_u10_u7_U89 (.ZN( u2_out10_15 ) , .A4( u2_u10_u7_n142 ) , .A3( u2_u10_u7_n143 ) , .A2( u2_u10_u7_n144 ) , .A1( u2_u10_u7_n178 ) );
  OAI221_X1 u2_u10_u7_U9 (.C1( u2_u10_u7_n101 ) , .C2( u2_u10_u7_n147 ) , .ZN( u2_u10_u7_n155 ) , .B2( u2_u10_u7_n162 ) , .A( u2_u10_u7_n91 ) , .B1( u2_u10_u7_n92 ) );
  OR2_X1 u2_u10_u7_U90 (.A2( u2_u10_u7_n125 ) , .A1( u2_u10_u7_n129 ) , .ZN( u2_u10_u7_n144 ) );
  AOI22_X1 u2_u10_u7_U91 (.A2( u2_u10_u7_n126 ) , .ZN( u2_u10_u7_n143 ) , .B2( u2_u10_u7_n165 ) , .B1( u2_u10_u7_n173 ) , .A1( u2_u10_u7_n174 ) );
  NAND4_X1 u2_u10_u7_U92 (.ZN( u2_out10_5 ) , .A4( u2_u10_u7_n108 ) , .A3( u2_u10_u7_n109 ) , .A1( u2_u10_u7_n116 ) , .A2( u2_u10_u7_n123 ) );
  AOI22_X1 u2_u10_u7_U93 (.ZN( u2_u10_u7_n109 ) , .A2( u2_u10_u7_n126 ) , .B2( u2_u10_u7_n145 ) , .B1( u2_u10_u7_n156 ) , .A1( u2_u10_u7_n171 ) );
  NOR4_X1 u2_u10_u7_U94 (.A4( u2_u10_u7_n104 ) , .A3( u2_u10_u7_n105 ) , .A2( u2_u10_u7_n106 ) , .A1( u2_u10_u7_n107 ) , .ZN( u2_u10_u7_n108 ) );
  NAND3_X1 u2_u10_u7_U95 (.A3( u2_u10_u7_n146 ) , .A2( u2_u10_u7_n147 ) , .A1( u2_u10_u7_n148 ) , .ZN( u2_u10_u7_n151 ) );
  NAND3_X1 u2_u10_u7_U96 (.A3( u2_u10_u7_n131 ) , .A2( u2_u10_u7_n132 ) , .A1( u2_u10_u7_n133 ) , .ZN( u2_u10_u7_n135 ) );
  XOR2_X1 u2_u11_U11 (.B( u2_K12_44 ) , .A( u2_R10_29 ) , .Z( u2_u11_X_44 ) );
  XOR2_X1 u2_u11_U13 (.B( u2_K12_42 ) , .A( u2_R10_29 ) , .Z( u2_u11_X_42 ) );
  XOR2_X1 u2_u11_U18 (.B( u2_K12_38 ) , .A( u2_R10_25 ) , .Z( u2_u11_X_38 ) );
  XOR2_X1 u2_u11_U20 (.B( u2_K12_36 ) , .A( u2_R10_25 ) , .Z( u2_u11_X_36 ) );
  XOR2_X1 u2_u11_U24 (.B( u2_K12_32 ) , .A( u2_R10_21 ) , .Z( u2_u11_X_32 ) );
  XOR2_X1 u2_u11_U26 (.B( u2_K12_30 ) , .A( u2_R10_21 ) , .Z( u2_u11_X_30 ) );
  XOR2_X1 u2_u11_U27 (.B( u2_K12_2 ) , .A( u2_R10_1 ) , .Z( u2_u11_X_2 ) );
  XOR2_X1 u2_u11_U3 (.B( u2_K12_7 ) , .A( u2_R10_4 ) , .Z( u2_u11_X_7 ) );
  XOR2_X1 u2_u11_U32 (.B( u2_K12_25 ) , .A( u2_R10_16 ) , .Z( u2_u11_X_25 ) );
  XOR2_X1 u2_u11_U34 (.B( u2_K12_23 ) , .A( u2_R10_16 ) , .Z( u2_u11_X_23 ) );
  XOR2_X1 u2_u11_U37 (.B( u2_K12_20 ) , .A( u2_R10_13 ) , .Z( u2_u11_X_20 ) );
  XOR2_X1 u2_u11_U38 (.B( u2_K12_1 ) , .A( u2_R10_32 ) , .Z( u2_u11_X_1 ) );
  XOR2_X1 u2_u11_U39 (.B( u2_K12_19 ) , .A( u2_R10_12 ) , .Z( u2_u11_X_19 ) );
  XOR2_X1 u2_u11_U40 (.B( u2_K12_18 ) , .A( u2_R10_13 ) , .Z( u2_u11_X_18 ) );
  XOR2_X1 u2_u11_U41 (.B( u2_K12_17 ) , .A( u2_R10_12 ) , .Z( u2_u11_X_17 ) );
  XOR2_X1 u2_u11_U44 (.B( u2_K12_14 ) , .A( u2_R10_9 ) , .Z( u2_u11_X_14 ) );
  XOR2_X1 u2_u11_U45 (.B( u2_K12_13 ) , .A( u2_R10_8 ) , .Z( u2_u11_X_13 ) );
  XOR2_X1 u2_u11_U46 (.B( u2_K12_12 ) , .A( u2_R10_9 ) , .Z( u2_u11_X_12 ) );
  XOR2_X1 u2_u11_U47 (.B( u2_K12_11 ) , .A( u2_R10_8 ) , .Z( u2_u11_X_11 ) );
  XOR2_X1 u2_u11_U48 (.B( u2_K12_10 ) , .A( u2_R10_7 ) , .Z( u2_u11_X_10 ) );
  XOR2_X1 u2_u11_U5 (.B( u2_K12_5 ) , .A( u2_R10_4 ) , .Z( u2_u11_X_5 ) );
  XOR2_X1 u2_u11_U6 (.B( u2_K12_4 ) , .A( u2_R10_3 ) , .Z( u2_u11_X_4 ) );
  XOR2_X1 u2_u11_U7 (.B( u2_K12_48 ) , .A( u2_R10_1 ) , .Z( u2_u11_X_48 ) );
  XOR2_X1 u2_u11_U8 (.B( u2_K12_47 ) , .A( u2_R10_32 ) , .Z( u2_u11_X_47 ) );
  NAND2_X1 u2_u11_u0_U10 (.ZN( u2_u11_u0_n113 ) , .A1( u2_u11_u0_n139 ) , .A2( u2_u11_u0_n149 ) );
  AND3_X1 u2_u11_u0_U11 (.A2( u2_u11_u0_n112 ) , .ZN( u2_u11_u0_n127 ) , .A3( u2_u11_u0_n130 ) , .A1( u2_u11_u0_n148 ) );
  AND2_X1 u2_u11_u0_U12 (.ZN( u2_u11_u0_n107 ) , .A1( u2_u11_u0_n130 ) , .A2( u2_u11_u0_n140 ) );
  AND2_X1 u2_u11_u0_U13 (.A2( u2_u11_u0_n129 ) , .A1( u2_u11_u0_n130 ) , .ZN( u2_u11_u0_n151 ) );
  AND2_X1 u2_u11_u0_U14 (.A1( u2_u11_u0_n108 ) , .A2( u2_u11_u0_n125 ) , .ZN( u2_u11_u0_n145 ) );
  INV_X1 u2_u11_u0_U15 (.A( u2_u11_u0_n143 ) , .ZN( u2_u11_u0_n173 ) );
  NOR2_X1 u2_u11_u0_U16 (.A2( u2_u11_u0_n136 ) , .ZN( u2_u11_u0_n147 ) , .A1( u2_u11_u0_n160 ) );
  OAI22_X1 u2_u11_u0_U17 (.B1( u2_u11_u0_n125 ) , .ZN( u2_u11_u0_n126 ) , .A1( u2_u11_u0_n138 ) , .A2( u2_u11_u0_n146 ) , .B2( u2_u11_u0_n147 ) );
  OAI22_X1 u2_u11_u0_U18 (.B1( u2_u11_u0_n131 ) , .A1( u2_u11_u0_n144 ) , .B2( u2_u11_u0_n147 ) , .A2( u2_u11_u0_n90 ) , .ZN( u2_u11_u0_n91 ) );
  AND3_X1 u2_u11_u0_U19 (.A3( u2_u11_u0_n121 ) , .A2( u2_u11_u0_n125 ) , .A1( u2_u11_u0_n148 ) , .ZN( u2_u11_u0_n90 ) );
  NOR2_X1 u2_u11_u0_U20 (.A1( u2_u11_u0_n163 ) , .A2( u2_u11_u0_n164 ) , .ZN( u2_u11_u0_n95 ) );
  NAND2_X1 u2_u11_u0_U21 (.A1( u2_u11_u0_n101 ) , .A2( u2_u11_u0_n102 ) , .ZN( u2_u11_u0_n150 ) );
  AOI22_X1 u2_u11_u0_U22 (.B2( u2_u11_u0_n109 ) , .A2( u2_u11_u0_n110 ) , .ZN( u2_u11_u0_n111 ) , .B1( u2_u11_u0_n118 ) , .A1( u2_u11_u0_n160 ) );
  NAND2_X1 u2_u11_u0_U23 (.A1( u2_u11_u0_n100 ) , .A2( u2_u11_u0_n103 ) , .ZN( u2_u11_u0_n125 ) );
  INV_X1 u2_u11_u0_U24 (.A( u2_u11_u0_n136 ) , .ZN( u2_u11_u0_n161 ) );
  INV_X1 u2_u11_u0_U25 (.A( u2_u11_u0_n118 ) , .ZN( u2_u11_u0_n158 ) );
  NAND2_X1 u2_u11_u0_U26 (.A2( u2_u11_u0_n100 ) , .A1( u2_u11_u0_n101 ) , .ZN( u2_u11_u0_n139 ) );
  NAND2_X1 u2_u11_u0_U27 (.A2( u2_u11_u0_n100 ) , .ZN( u2_u11_u0_n131 ) , .A1( u2_u11_u0_n92 ) );
  NAND2_X1 u2_u11_u0_U28 (.ZN( u2_u11_u0_n108 ) , .A1( u2_u11_u0_n92 ) , .A2( u2_u11_u0_n94 ) );
  AOI21_X1 u2_u11_u0_U29 (.B1( u2_u11_u0_n127 ) , .B2( u2_u11_u0_n129 ) , .A( u2_u11_u0_n138 ) , .ZN( u2_u11_u0_n96 ) );
  INV_X1 u2_u11_u0_U3 (.A( u2_u11_u0_n113 ) , .ZN( u2_u11_u0_n166 ) );
  AOI21_X1 u2_u11_u0_U30 (.ZN( u2_u11_u0_n104 ) , .B1( u2_u11_u0_n107 ) , .B2( u2_u11_u0_n141 ) , .A( u2_u11_u0_n144 ) );
  NAND2_X1 u2_u11_u0_U31 (.A2( u2_u11_u0_n102 ) , .ZN( u2_u11_u0_n114 ) , .A1( u2_u11_u0_n92 ) );
  NAND2_X1 u2_u11_u0_U32 (.A1( u2_u11_u0_n101 ) , .ZN( u2_u11_u0_n130 ) , .A2( u2_u11_u0_n94 ) );
  NOR2_X1 u2_u11_u0_U33 (.A1( u2_u11_u0_n120 ) , .ZN( u2_u11_u0_n143 ) , .A2( u2_u11_u0_n167 ) );
  OAI221_X1 u2_u11_u0_U34 (.C1( u2_u11_u0_n112 ) , .ZN( u2_u11_u0_n120 ) , .B1( u2_u11_u0_n138 ) , .B2( u2_u11_u0_n141 ) , .C2( u2_u11_u0_n147 ) , .A( u2_u11_u0_n172 ) );
  AOI211_X1 u2_u11_u0_U35 (.B( u2_u11_u0_n115 ) , .A( u2_u11_u0_n116 ) , .C2( u2_u11_u0_n117 ) , .C1( u2_u11_u0_n118 ) , .ZN( u2_u11_u0_n119 ) );
  NAND2_X1 u2_u11_u0_U36 (.A2( u2_u11_u0_n103 ) , .ZN( u2_u11_u0_n140 ) , .A1( u2_u11_u0_n94 ) );
  INV_X1 u2_u11_u0_U37 (.A( u2_u11_u0_n138 ) , .ZN( u2_u11_u0_n160 ) );
  NAND2_X1 u2_u11_u0_U38 (.A2( u2_u11_u0_n102 ) , .A1( u2_u11_u0_n103 ) , .ZN( u2_u11_u0_n149 ) );
  NAND2_X1 u2_u11_u0_U39 (.A2( u2_u11_u0_n101 ) , .ZN( u2_u11_u0_n121 ) , .A1( u2_u11_u0_n93 ) );
  AOI21_X1 u2_u11_u0_U4 (.B1( u2_u11_u0_n114 ) , .ZN( u2_u11_u0_n115 ) , .B2( u2_u11_u0_n129 ) , .A( u2_u11_u0_n161 ) );
  NAND2_X1 u2_u11_u0_U40 (.ZN( u2_u11_u0_n112 ) , .A2( u2_u11_u0_n92 ) , .A1( u2_u11_u0_n93 ) );
  INV_X1 u2_u11_u0_U41 (.ZN( u2_u11_u0_n172 ) , .A( u2_u11_u0_n88 ) );
  OAI222_X1 u2_u11_u0_U42 (.C1( u2_u11_u0_n108 ) , .A1( u2_u11_u0_n125 ) , .B2( u2_u11_u0_n128 ) , .B1( u2_u11_u0_n144 ) , .A2( u2_u11_u0_n158 ) , .C2( u2_u11_u0_n161 ) , .ZN( u2_u11_u0_n88 ) );
  AOI21_X1 u2_u11_u0_U43 (.B1( u2_u11_u0_n103 ) , .ZN( u2_u11_u0_n132 ) , .A( u2_u11_u0_n165 ) , .B2( u2_u11_u0_n93 ) );
  OR3_X1 u2_u11_u0_U44 (.A3( u2_u11_u0_n152 ) , .A2( u2_u11_u0_n153 ) , .A1( u2_u11_u0_n154 ) , .ZN( u2_u11_u0_n155 ) );
  AOI21_X1 u2_u11_u0_U45 (.A( u2_u11_u0_n144 ) , .B2( u2_u11_u0_n145 ) , .B1( u2_u11_u0_n146 ) , .ZN( u2_u11_u0_n154 ) );
  AOI21_X1 u2_u11_u0_U46 (.B2( u2_u11_u0_n150 ) , .B1( u2_u11_u0_n151 ) , .ZN( u2_u11_u0_n152 ) , .A( u2_u11_u0_n158 ) );
  AOI21_X1 u2_u11_u0_U47 (.A( u2_u11_u0_n147 ) , .B2( u2_u11_u0_n148 ) , .B1( u2_u11_u0_n149 ) , .ZN( u2_u11_u0_n153 ) );
  INV_X1 u2_u11_u0_U48 (.ZN( u2_u11_u0_n171 ) , .A( u2_u11_u0_n99 ) );
  OAI211_X1 u2_u11_u0_U49 (.C2( u2_u11_u0_n140 ) , .C1( u2_u11_u0_n161 ) , .A( u2_u11_u0_n169 ) , .B( u2_u11_u0_n98 ) , .ZN( u2_u11_u0_n99 ) );
  AOI21_X1 u2_u11_u0_U5 (.B2( u2_u11_u0_n131 ) , .ZN( u2_u11_u0_n134 ) , .B1( u2_u11_u0_n151 ) , .A( u2_u11_u0_n158 ) );
  AOI211_X1 u2_u11_u0_U50 (.C1( u2_u11_u0_n118 ) , .A( u2_u11_u0_n123 ) , .B( u2_u11_u0_n96 ) , .C2( u2_u11_u0_n97 ) , .ZN( u2_u11_u0_n98 ) );
  INV_X1 u2_u11_u0_U51 (.ZN( u2_u11_u0_n169 ) , .A( u2_u11_u0_n91 ) );
  NOR2_X1 u2_u11_u0_U52 (.A2( u2_u11_X_2 ) , .ZN( u2_u11_u0_n103 ) , .A1( u2_u11_u0_n164 ) );
  NOR2_X1 u2_u11_u0_U53 (.A2( u2_u11_X_4 ) , .A1( u2_u11_X_5 ) , .ZN( u2_u11_u0_n118 ) );
  NOR2_X1 u2_u11_u0_U54 (.A2( u2_u11_X_3 ) , .A1( u2_u11_X_6 ) , .ZN( u2_u11_u0_n94 ) );
  NAND2_X1 u2_u11_u0_U55 (.A2( u2_u11_X_4 ) , .A1( u2_u11_X_5 ) , .ZN( u2_u11_u0_n144 ) );
  NOR2_X1 u2_u11_u0_U56 (.A2( u2_u11_X_5 ) , .ZN( u2_u11_u0_n136 ) , .A1( u2_u11_u0_n159 ) );
  NAND2_X1 u2_u11_u0_U57 (.A1( u2_u11_X_5 ) , .ZN( u2_u11_u0_n138 ) , .A2( u2_u11_u0_n159 ) );
  AND2_X1 u2_u11_u0_U58 (.A2( u2_u11_X_3 ) , .A1( u2_u11_X_6 ) , .ZN( u2_u11_u0_n102 ) );
  AND2_X1 u2_u11_u0_U59 (.A1( u2_u11_X_6 ) , .A2( u2_u11_u0_n162 ) , .ZN( u2_u11_u0_n93 ) );
  NOR2_X1 u2_u11_u0_U6 (.A1( u2_u11_u0_n108 ) , .ZN( u2_u11_u0_n123 ) , .A2( u2_u11_u0_n158 ) );
  INV_X1 u2_u11_u0_U60 (.A( u2_u11_X_4 ) , .ZN( u2_u11_u0_n159 ) );
  INV_X1 u2_u11_u0_U61 (.A( u2_u11_X_2 ) , .ZN( u2_u11_u0_n163 ) );
  INV_X1 u2_u11_u0_U62 (.A( u2_u11_u0_n126 ) , .ZN( u2_u11_u0_n168 ) );
  AOI211_X1 u2_u11_u0_U63 (.B( u2_u11_u0_n133 ) , .A( u2_u11_u0_n134 ) , .C2( u2_u11_u0_n135 ) , .C1( u2_u11_u0_n136 ) , .ZN( u2_u11_u0_n137 ) );
  OR4_X1 u2_u11_u0_U64 (.ZN( u2_out11_17 ) , .A4( u2_u11_u0_n122 ) , .A2( u2_u11_u0_n123 ) , .A1( u2_u11_u0_n124 ) , .A3( u2_u11_u0_n170 ) );
  AOI21_X1 u2_u11_u0_U65 (.B2( u2_u11_u0_n107 ) , .ZN( u2_u11_u0_n124 ) , .B1( u2_u11_u0_n128 ) , .A( u2_u11_u0_n161 ) );
  INV_X1 u2_u11_u0_U66 (.A( u2_u11_u0_n111 ) , .ZN( u2_u11_u0_n170 ) );
  OR4_X1 u2_u11_u0_U67 (.ZN( u2_out11_31 ) , .A4( u2_u11_u0_n155 ) , .A2( u2_u11_u0_n156 ) , .A1( u2_u11_u0_n157 ) , .A3( u2_u11_u0_n173 ) );
  AOI21_X1 u2_u11_u0_U68 (.A( u2_u11_u0_n138 ) , .B2( u2_u11_u0_n139 ) , .B1( u2_u11_u0_n140 ) , .ZN( u2_u11_u0_n157 ) );
  INV_X1 u2_u11_u0_U69 (.ZN( u2_u11_u0_n174 ) , .A( u2_u11_u0_n89 ) );
  OAI21_X1 u2_u11_u0_U7 (.B1( u2_u11_u0_n150 ) , .B2( u2_u11_u0_n158 ) , .A( u2_u11_u0_n172 ) , .ZN( u2_u11_u0_n89 ) );
  AOI211_X1 u2_u11_u0_U70 (.B( u2_u11_u0_n104 ) , .A( u2_u11_u0_n105 ) , .ZN( u2_u11_u0_n106 ) , .C2( u2_u11_u0_n113 ) , .C1( u2_u11_u0_n160 ) );
  INV_X1 u2_u11_u0_U71 (.A( u2_u11_u0_n142 ) , .ZN( u2_u11_u0_n165 ) );
  AOI21_X1 u2_u11_u0_U72 (.ZN( u2_u11_u0_n116 ) , .B2( u2_u11_u0_n142 ) , .A( u2_u11_u0_n144 ) , .B1( u2_u11_u0_n166 ) );
  AOI21_X1 u2_u11_u0_U73 (.B2( u2_u11_u0_n141 ) , .B1( u2_u11_u0_n142 ) , .ZN( u2_u11_u0_n156 ) , .A( u2_u11_u0_n161 ) );
  OAI221_X1 u2_u11_u0_U74 (.C1( u2_u11_u0_n121 ) , .ZN( u2_u11_u0_n122 ) , .B2( u2_u11_u0_n127 ) , .A( u2_u11_u0_n143 ) , .B1( u2_u11_u0_n144 ) , .C2( u2_u11_u0_n147 ) );
  NOR2_X1 u2_u11_u0_U75 (.A2( u2_u11_X_6 ) , .ZN( u2_u11_u0_n100 ) , .A1( u2_u11_u0_n162 ) );
  INV_X1 u2_u11_u0_U76 (.A( u2_u11_X_3 ) , .ZN( u2_u11_u0_n162 ) );
  AOI21_X1 u2_u11_u0_U77 (.B1( u2_u11_u0_n132 ) , .ZN( u2_u11_u0_n133 ) , .A( u2_u11_u0_n144 ) , .B2( u2_u11_u0_n166 ) );
  OAI22_X1 u2_u11_u0_U78 (.ZN( u2_u11_u0_n105 ) , .A2( u2_u11_u0_n132 ) , .B1( u2_u11_u0_n146 ) , .A1( u2_u11_u0_n147 ) , .B2( u2_u11_u0_n161 ) );
  NAND2_X1 u2_u11_u0_U79 (.ZN( u2_u11_u0_n110 ) , .A2( u2_u11_u0_n132 ) , .A1( u2_u11_u0_n145 ) );
  AND2_X1 u2_u11_u0_U8 (.A1( u2_u11_u0_n114 ) , .A2( u2_u11_u0_n121 ) , .ZN( u2_u11_u0_n146 ) );
  INV_X1 u2_u11_u0_U80 (.A( u2_u11_u0_n119 ) , .ZN( u2_u11_u0_n167 ) );
  NAND2_X1 u2_u11_u0_U81 (.ZN( u2_u11_u0_n148 ) , .A1( u2_u11_u0_n93 ) , .A2( u2_u11_u0_n95 ) );
  NAND2_X1 u2_u11_u0_U82 (.A1( u2_u11_u0_n100 ) , .ZN( u2_u11_u0_n129 ) , .A2( u2_u11_u0_n95 ) );
  NAND2_X1 u2_u11_u0_U83 (.A1( u2_u11_u0_n102 ) , .ZN( u2_u11_u0_n128 ) , .A2( u2_u11_u0_n95 ) );
  NOR2_X1 u2_u11_u0_U84 (.A2( u2_u11_X_1 ) , .A1( u2_u11_X_2 ) , .ZN( u2_u11_u0_n92 ) );
  NAND2_X1 u2_u11_u0_U85 (.ZN( u2_u11_u0_n142 ) , .A1( u2_u11_u0_n94 ) , .A2( u2_u11_u0_n95 ) );
  NOR2_X1 u2_u11_u0_U86 (.A2( u2_u11_X_1 ) , .ZN( u2_u11_u0_n101 ) , .A1( u2_u11_u0_n163 ) );
  INV_X1 u2_u11_u0_U87 (.A( u2_u11_X_1 ) , .ZN( u2_u11_u0_n164 ) );
  NAND3_X1 u2_u11_u0_U88 (.ZN( u2_out11_23 ) , .A3( u2_u11_u0_n137 ) , .A1( u2_u11_u0_n168 ) , .A2( u2_u11_u0_n171 ) );
  NAND3_X1 u2_u11_u0_U89 (.A3( u2_u11_u0_n127 ) , .A2( u2_u11_u0_n128 ) , .ZN( u2_u11_u0_n135 ) , .A1( u2_u11_u0_n150 ) );
  AND2_X1 u2_u11_u0_U9 (.A1( u2_u11_u0_n131 ) , .ZN( u2_u11_u0_n141 ) , .A2( u2_u11_u0_n150 ) );
  NAND3_X1 u2_u11_u0_U90 (.ZN( u2_u11_u0_n117 ) , .A3( u2_u11_u0_n132 ) , .A2( u2_u11_u0_n139 ) , .A1( u2_u11_u0_n148 ) );
  NAND3_X1 u2_u11_u0_U91 (.ZN( u2_u11_u0_n109 ) , .A2( u2_u11_u0_n114 ) , .A3( u2_u11_u0_n140 ) , .A1( u2_u11_u0_n149 ) );
  NAND3_X1 u2_u11_u0_U92 (.ZN( u2_out11_9 ) , .A3( u2_u11_u0_n106 ) , .A2( u2_u11_u0_n171 ) , .A1( u2_u11_u0_n174 ) );
  NAND3_X1 u2_u11_u0_U93 (.A2( u2_u11_u0_n128 ) , .A1( u2_u11_u0_n132 ) , .A3( u2_u11_u0_n146 ) , .ZN( u2_u11_u0_n97 ) );
  NOR2_X1 u2_u11_u1_U10 (.A1( u2_u11_u1_n112 ) , .A2( u2_u11_u1_n116 ) , .ZN( u2_u11_u1_n118 ) );
  NAND3_X1 u2_u11_u1_U100 (.ZN( u2_u11_u1_n113 ) , .A1( u2_u11_u1_n120 ) , .A3( u2_u11_u1_n133 ) , .A2( u2_u11_u1_n155 ) );
  OAI21_X1 u2_u11_u1_U11 (.ZN( u2_u11_u1_n101 ) , .B1( u2_u11_u1_n141 ) , .A( u2_u11_u1_n146 ) , .B2( u2_u11_u1_n183 ) );
  AOI21_X1 u2_u11_u1_U12 (.B2( u2_u11_u1_n155 ) , .B1( u2_u11_u1_n156 ) , .ZN( u2_u11_u1_n157 ) , .A( u2_u11_u1_n174 ) );
  NAND2_X1 u2_u11_u1_U13 (.ZN( u2_u11_u1_n140 ) , .A2( u2_u11_u1_n150 ) , .A1( u2_u11_u1_n155 ) );
  NAND2_X1 u2_u11_u1_U14 (.A1( u2_u11_u1_n131 ) , .ZN( u2_u11_u1_n147 ) , .A2( u2_u11_u1_n153 ) );
  INV_X1 u2_u11_u1_U15 (.A( u2_u11_u1_n139 ) , .ZN( u2_u11_u1_n174 ) );
  OR4_X1 u2_u11_u1_U16 (.A4( u2_u11_u1_n106 ) , .A3( u2_u11_u1_n107 ) , .ZN( u2_u11_u1_n108 ) , .A1( u2_u11_u1_n117 ) , .A2( u2_u11_u1_n184 ) );
  AOI21_X1 u2_u11_u1_U17 (.ZN( u2_u11_u1_n106 ) , .A( u2_u11_u1_n112 ) , .B1( u2_u11_u1_n154 ) , .B2( u2_u11_u1_n156 ) );
  AOI21_X1 u2_u11_u1_U18 (.ZN( u2_u11_u1_n107 ) , .B1( u2_u11_u1_n134 ) , .B2( u2_u11_u1_n149 ) , .A( u2_u11_u1_n174 ) );
  INV_X1 u2_u11_u1_U19 (.A( u2_u11_u1_n101 ) , .ZN( u2_u11_u1_n184 ) );
  INV_X1 u2_u11_u1_U20 (.A( u2_u11_u1_n112 ) , .ZN( u2_u11_u1_n171 ) );
  NAND2_X1 u2_u11_u1_U21 (.ZN( u2_u11_u1_n141 ) , .A1( u2_u11_u1_n153 ) , .A2( u2_u11_u1_n156 ) );
  AND2_X1 u2_u11_u1_U22 (.A1( u2_u11_u1_n123 ) , .ZN( u2_u11_u1_n134 ) , .A2( u2_u11_u1_n161 ) );
  NAND2_X1 u2_u11_u1_U23 (.A2( u2_u11_u1_n115 ) , .A1( u2_u11_u1_n116 ) , .ZN( u2_u11_u1_n148 ) );
  NAND2_X1 u2_u11_u1_U24 (.A2( u2_u11_u1_n133 ) , .A1( u2_u11_u1_n135 ) , .ZN( u2_u11_u1_n159 ) );
  NAND2_X1 u2_u11_u1_U25 (.A2( u2_u11_u1_n115 ) , .A1( u2_u11_u1_n120 ) , .ZN( u2_u11_u1_n132 ) );
  INV_X1 u2_u11_u1_U26 (.A( u2_u11_u1_n154 ) , .ZN( u2_u11_u1_n178 ) );
  INV_X1 u2_u11_u1_U27 (.A( u2_u11_u1_n151 ) , .ZN( u2_u11_u1_n183 ) );
  AND2_X1 u2_u11_u1_U28 (.A1( u2_u11_u1_n129 ) , .A2( u2_u11_u1_n133 ) , .ZN( u2_u11_u1_n149 ) );
  INV_X1 u2_u11_u1_U29 (.A( u2_u11_u1_n131 ) , .ZN( u2_u11_u1_n180 ) );
  INV_X1 u2_u11_u1_U3 (.A( u2_u11_u1_n159 ) , .ZN( u2_u11_u1_n182 ) );
  OAI221_X1 u2_u11_u1_U30 (.A( u2_u11_u1_n119 ) , .C2( u2_u11_u1_n129 ) , .ZN( u2_u11_u1_n138 ) , .B2( u2_u11_u1_n152 ) , .C1( u2_u11_u1_n174 ) , .B1( u2_u11_u1_n187 ) );
  INV_X1 u2_u11_u1_U31 (.A( u2_u11_u1_n148 ) , .ZN( u2_u11_u1_n187 ) );
  AOI211_X1 u2_u11_u1_U32 (.B( u2_u11_u1_n117 ) , .A( u2_u11_u1_n118 ) , .ZN( u2_u11_u1_n119 ) , .C2( u2_u11_u1_n146 ) , .C1( u2_u11_u1_n159 ) );
  NOR2_X1 u2_u11_u1_U33 (.A1( u2_u11_u1_n168 ) , .A2( u2_u11_u1_n176 ) , .ZN( u2_u11_u1_n98 ) );
  AOI211_X1 u2_u11_u1_U34 (.B( u2_u11_u1_n162 ) , .A( u2_u11_u1_n163 ) , .C2( u2_u11_u1_n164 ) , .ZN( u2_u11_u1_n165 ) , .C1( u2_u11_u1_n171 ) );
  AOI21_X1 u2_u11_u1_U35 (.A( u2_u11_u1_n160 ) , .B2( u2_u11_u1_n161 ) , .ZN( u2_u11_u1_n162 ) , .B1( u2_u11_u1_n182 ) );
  OR2_X1 u2_u11_u1_U36 (.A2( u2_u11_u1_n157 ) , .A1( u2_u11_u1_n158 ) , .ZN( u2_u11_u1_n163 ) );
  NAND2_X1 u2_u11_u1_U37 (.A1( u2_u11_u1_n128 ) , .ZN( u2_u11_u1_n146 ) , .A2( u2_u11_u1_n160 ) );
  NAND2_X1 u2_u11_u1_U38 (.A2( u2_u11_u1_n112 ) , .ZN( u2_u11_u1_n139 ) , .A1( u2_u11_u1_n152 ) );
  NAND2_X1 u2_u11_u1_U39 (.A1( u2_u11_u1_n105 ) , .ZN( u2_u11_u1_n156 ) , .A2( u2_u11_u1_n99 ) );
  AOI221_X1 u2_u11_u1_U4 (.A( u2_u11_u1_n138 ) , .C2( u2_u11_u1_n139 ) , .C1( u2_u11_u1_n140 ) , .B2( u2_u11_u1_n141 ) , .ZN( u2_u11_u1_n142 ) , .B1( u2_u11_u1_n175 ) );
  AOI221_X1 u2_u11_u1_U40 (.B1( u2_u11_u1_n140 ) , .ZN( u2_u11_u1_n167 ) , .B2( u2_u11_u1_n172 ) , .C2( u2_u11_u1_n175 ) , .C1( u2_u11_u1_n178 ) , .A( u2_u11_u1_n188 ) );
  INV_X1 u2_u11_u1_U41 (.ZN( u2_u11_u1_n188 ) , .A( u2_u11_u1_n97 ) );
  AOI211_X1 u2_u11_u1_U42 (.A( u2_u11_u1_n118 ) , .C1( u2_u11_u1_n132 ) , .C2( u2_u11_u1_n139 ) , .B( u2_u11_u1_n96 ) , .ZN( u2_u11_u1_n97 ) );
  AOI21_X1 u2_u11_u1_U43 (.B2( u2_u11_u1_n121 ) , .B1( u2_u11_u1_n135 ) , .A( u2_u11_u1_n152 ) , .ZN( u2_u11_u1_n96 ) );
  NOR2_X1 u2_u11_u1_U44 (.ZN( u2_u11_u1_n117 ) , .A1( u2_u11_u1_n121 ) , .A2( u2_u11_u1_n160 ) );
  OAI21_X1 u2_u11_u1_U45 (.B2( u2_u11_u1_n123 ) , .ZN( u2_u11_u1_n145 ) , .B1( u2_u11_u1_n160 ) , .A( u2_u11_u1_n185 ) );
  INV_X1 u2_u11_u1_U46 (.A( u2_u11_u1_n122 ) , .ZN( u2_u11_u1_n185 ) );
  AOI21_X1 u2_u11_u1_U47 (.B2( u2_u11_u1_n120 ) , .B1( u2_u11_u1_n121 ) , .ZN( u2_u11_u1_n122 ) , .A( u2_u11_u1_n128 ) );
  AOI21_X1 u2_u11_u1_U48 (.A( u2_u11_u1_n128 ) , .B2( u2_u11_u1_n129 ) , .ZN( u2_u11_u1_n130 ) , .B1( u2_u11_u1_n150 ) );
  NAND2_X1 u2_u11_u1_U49 (.ZN( u2_u11_u1_n112 ) , .A1( u2_u11_u1_n169 ) , .A2( u2_u11_u1_n170 ) );
  AOI211_X1 u2_u11_u1_U5 (.ZN( u2_u11_u1_n124 ) , .A( u2_u11_u1_n138 ) , .C2( u2_u11_u1_n139 ) , .B( u2_u11_u1_n145 ) , .C1( u2_u11_u1_n147 ) );
  NAND2_X1 u2_u11_u1_U50 (.ZN( u2_u11_u1_n129 ) , .A2( u2_u11_u1_n95 ) , .A1( u2_u11_u1_n98 ) );
  NAND2_X1 u2_u11_u1_U51 (.A1( u2_u11_u1_n102 ) , .ZN( u2_u11_u1_n154 ) , .A2( u2_u11_u1_n99 ) );
  NAND2_X1 u2_u11_u1_U52 (.A2( u2_u11_u1_n100 ) , .ZN( u2_u11_u1_n135 ) , .A1( u2_u11_u1_n99 ) );
  AOI21_X1 u2_u11_u1_U53 (.A( u2_u11_u1_n152 ) , .B2( u2_u11_u1_n153 ) , .B1( u2_u11_u1_n154 ) , .ZN( u2_u11_u1_n158 ) );
  INV_X1 u2_u11_u1_U54 (.A( u2_u11_u1_n160 ) , .ZN( u2_u11_u1_n175 ) );
  NAND2_X1 u2_u11_u1_U55 (.A1( u2_u11_u1_n100 ) , .ZN( u2_u11_u1_n116 ) , .A2( u2_u11_u1_n95 ) );
  NAND2_X1 u2_u11_u1_U56 (.A1( u2_u11_u1_n102 ) , .ZN( u2_u11_u1_n131 ) , .A2( u2_u11_u1_n95 ) );
  NAND2_X1 u2_u11_u1_U57 (.A2( u2_u11_u1_n104 ) , .ZN( u2_u11_u1_n121 ) , .A1( u2_u11_u1_n98 ) );
  NAND2_X1 u2_u11_u1_U58 (.A1( u2_u11_u1_n103 ) , .ZN( u2_u11_u1_n153 ) , .A2( u2_u11_u1_n98 ) );
  NAND2_X1 u2_u11_u1_U59 (.A2( u2_u11_u1_n104 ) , .A1( u2_u11_u1_n105 ) , .ZN( u2_u11_u1_n133 ) );
  AOI22_X1 u2_u11_u1_U6 (.B2( u2_u11_u1_n113 ) , .A2( u2_u11_u1_n114 ) , .ZN( u2_u11_u1_n125 ) , .A1( u2_u11_u1_n171 ) , .B1( u2_u11_u1_n173 ) );
  NAND2_X1 u2_u11_u1_U60 (.ZN( u2_u11_u1_n150 ) , .A2( u2_u11_u1_n98 ) , .A1( u2_u11_u1_n99 ) );
  NAND2_X1 u2_u11_u1_U61 (.A1( u2_u11_u1_n105 ) , .ZN( u2_u11_u1_n155 ) , .A2( u2_u11_u1_n95 ) );
  OAI21_X1 u2_u11_u1_U62 (.ZN( u2_u11_u1_n109 ) , .B1( u2_u11_u1_n129 ) , .B2( u2_u11_u1_n160 ) , .A( u2_u11_u1_n167 ) );
  NAND2_X1 u2_u11_u1_U63 (.A2( u2_u11_u1_n100 ) , .A1( u2_u11_u1_n103 ) , .ZN( u2_u11_u1_n120 ) );
  NAND2_X1 u2_u11_u1_U64 (.A1( u2_u11_u1_n102 ) , .A2( u2_u11_u1_n104 ) , .ZN( u2_u11_u1_n115 ) );
  NAND2_X1 u2_u11_u1_U65 (.A2( u2_u11_u1_n100 ) , .A1( u2_u11_u1_n104 ) , .ZN( u2_u11_u1_n151 ) );
  NAND2_X1 u2_u11_u1_U66 (.A2( u2_u11_u1_n103 ) , .A1( u2_u11_u1_n105 ) , .ZN( u2_u11_u1_n161 ) );
  INV_X1 u2_u11_u1_U67 (.A( u2_u11_u1_n152 ) , .ZN( u2_u11_u1_n173 ) );
  INV_X1 u2_u11_u1_U68 (.A( u2_u11_u1_n128 ) , .ZN( u2_u11_u1_n172 ) );
  NAND2_X1 u2_u11_u1_U69 (.A2( u2_u11_u1_n102 ) , .A1( u2_u11_u1_n103 ) , .ZN( u2_u11_u1_n123 ) );
  NAND2_X1 u2_u11_u1_U7 (.ZN( u2_u11_u1_n114 ) , .A1( u2_u11_u1_n134 ) , .A2( u2_u11_u1_n156 ) );
  NOR2_X1 u2_u11_u1_U70 (.A2( u2_u11_X_7 ) , .A1( u2_u11_X_8 ) , .ZN( u2_u11_u1_n95 ) );
  NOR2_X1 u2_u11_u1_U71 (.A1( u2_u11_X_12 ) , .A2( u2_u11_X_9 ) , .ZN( u2_u11_u1_n100 ) );
  NOR2_X1 u2_u11_u1_U72 (.A2( u2_u11_X_8 ) , .A1( u2_u11_u1_n177 ) , .ZN( u2_u11_u1_n99 ) );
  NOR2_X1 u2_u11_u1_U73 (.A2( u2_u11_X_12 ) , .ZN( u2_u11_u1_n102 ) , .A1( u2_u11_u1_n176 ) );
  NOR2_X1 u2_u11_u1_U74 (.A2( u2_u11_X_9 ) , .ZN( u2_u11_u1_n105 ) , .A1( u2_u11_u1_n168 ) );
  NAND2_X1 u2_u11_u1_U75 (.A1( u2_u11_X_10 ) , .ZN( u2_u11_u1_n160 ) , .A2( u2_u11_u1_n169 ) );
  NAND2_X1 u2_u11_u1_U76 (.A2( u2_u11_X_10 ) , .A1( u2_u11_X_11 ) , .ZN( u2_u11_u1_n152 ) );
  NAND2_X1 u2_u11_u1_U77 (.A1( u2_u11_X_11 ) , .ZN( u2_u11_u1_n128 ) , .A2( u2_u11_u1_n170 ) );
  AND2_X1 u2_u11_u1_U78 (.A2( u2_u11_X_7 ) , .A1( u2_u11_X_8 ) , .ZN( u2_u11_u1_n104 ) );
  AND2_X1 u2_u11_u1_U79 (.A1( u2_u11_X_8 ) , .ZN( u2_u11_u1_n103 ) , .A2( u2_u11_u1_n177 ) );
  AOI22_X1 u2_u11_u1_U8 (.B2( u2_u11_u1_n136 ) , .A2( u2_u11_u1_n137 ) , .ZN( u2_u11_u1_n143 ) , .A1( u2_u11_u1_n171 ) , .B1( u2_u11_u1_n173 ) );
  INV_X1 u2_u11_u1_U80 (.A( u2_u11_X_10 ) , .ZN( u2_u11_u1_n170 ) );
  INV_X1 u2_u11_u1_U81 (.A( u2_u11_X_9 ) , .ZN( u2_u11_u1_n176 ) );
  INV_X1 u2_u11_u1_U82 (.A( u2_u11_X_11 ) , .ZN( u2_u11_u1_n169 ) );
  INV_X1 u2_u11_u1_U83 (.A( u2_u11_X_12 ) , .ZN( u2_u11_u1_n168 ) );
  INV_X1 u2_u11_u1_U84 (.A( u2_u11_X_7 ) , .ZN( u2_u11_u1_n177 ) );
  NAND4_X1 u2_u11_u1_U85 (.ZN( u2_out11_28 ) , .A4( u2_u11_u1_n124 ) , .A3( u2_u11_u1_n125 ) , .A2( u2_u11_u1_n126 ) , .A1( u2_u11_u1_n127 ) );
  OAI21_X1 u2_u11_u1_U86 (.ZN( u2_u11_u1_n127 ) , .B2( u2_u11_u1_n139 ) , .B1( u2_u11_u1_n175 ) , .A( u2_u11_u1_n183 ) );
  OAI21_X1 u2_u11_u1_U87 (.ZN( u2_u11_u1_n126 ) , .B2( u2_u11_u1_n140 ) , .A( u2_u11_u1_n146 ) , .B1( u2_u11_u1_n178 ) );
  NAND4_X1 u2_u11_u1_U88 (.ZN( u2_out11_18 ) , .A4( u2_u11_u1_n165 ) , .A3( u2_u11_u1_n166 ) , .A1( u2_u11_u1_n167 ) , .A2( u2_u11_u1_n186 ) );
  AOI22_X1 u2_u11_u1_U89 (.B2( u2_u11_u1_n146 ) , .B1( u2_u11_u1_n147 ) , .A2( u2_u11_u1_n148 ) , .ZN( u2_u11_u1_n166 ) , .A1( u2_u11_u1_n172 ) );
  INV_X1 u2_u11_u1_U9 (.A( u2_u11_u1_n147 ) , .ZN( u2_u11_u1_n181 ) );
  INV_X1 u2_u11_u1_U90 (.A( u2_u11_u1_n145 ) , .ZN( u2_u11_u1_n186 ) );
  NAND4_X1 u2_u11_u1_U91 (.ZN( u2_out11_2 ) , .A4( u2_u11_u1_n142 ) , .A3( u2_u11_u1_n143 ) , .A2( u2_u11_u1_n144 ) , .A1( u2_u11_u1_n179 ) );
  OAI21_X1 u2_u11_u1_U92 (.B2( u2_u11_u1_n132 ) , .ZN( u2_u11_u1_n144 ) , .A( u2_u11_u1_n146 ) , .B1( u2_u11_u1_n180 ) );
  INV_X1 u2_u11_u1_U93 (.A( u2_u11_u1_n130 ) , .ZN( u2_u11_u1_n179 ) );
  OR4_X1 u2_u11_u1_U94 (.ZN( u2_out11_13 ) , .A4( u2_u11_u1_n108 ) , .A3( u2_u11_u1_n109 ) , .A2( u2_u11_u1_n110 ) , .A1( u2_u11_u1_n111 ) );
  AOI21_X1 u2_u11_u1_U95 (.ZN( u2_u11_u1_n111 ) , .A( u2_u11_u1_n128 ) , .B2( u2_u11_u1_n131 ) , .B1( u2_u11_u1_n135 ) );
  AOI21_X1 u2_u11_u1_U96 (.ZN( u2_u11_u1_n110 ) , .A( u2_u11_u1_n116 ) , .B1( u2_u11_u1_n152 ) , .B2( u2_u11_u1_n160 ) );
  NAND3_X1 u2_u11_u1_U97 (.A3( u2_u11_u1_n149 ) , .A2( u2_u11_u1_n150 ) , .A1( u2_u11_u1_n151 ) , .ZN( u2_u11_u1_n164 ) );
  NAND3_X1 u2_u11_u1_U98 (.A3( u2_u11_u1_n134 ) , .A2( u2_u11_u1_n135 ) , .ZN( u2_u11_u1_n136 ) , .A1( u2_u11_u1_n151 ) );
  NAND3_X1 u2_u11_u1_U99 (.A1( u2_u11_u1_n133 ) , .ZN( u2_u11_u1_n137 ) , .A2( u2_u11_u1_n154 ) , .A3( u2_u11_u1_n181 ) );
  OAI22_X1 u2_u11_u2_U10 (.ZN( u2_u11_u2_n109 ) , .A2( u2_u11_u2_n113 ) , .B2( u2_u11_u2_n133 ) , .B1( u2_u11_u2_n167 ) , .A1( u2_u11_u2_n168 ) );
  NAND3_X1 u2_u11_u2_U100 (.A2( u2_u11_u2_n100 ) , .A1( u2_u11_u2_n104 ) , .A3( u2_u11_u2_n138 ) , .ZN( u2_u11_u2_n98 ) );
  OAI22_X1 u2_u11_u2_U11 (.B1( u2_u11_u2_n151 ) , .A2( u2_u11_u2_n152 ) , .A1( u2_u11_u2_n153 ) , .ZN( u2_u11_u2_n160 ) , .B2( u2_u11_u2_n168 ) );
  NOR3_X1 u2_u11_u2_U12 (.A1( u2_u11_u2_n150 ) , .ZN( u2_u11_u2_n151 ) , .A3( u2_u11_u2_n175 ) , .A2( u2_u11_u2_n188 ) );
  AOI21_X1 u2_u11_u2_U13 (.ZN( u2_u11_u2_n144 ) , .B2( u2_u11_u2_n155 ) , .A( u2_u11_u2_n172 ) , .B1( u2_u11_u2_n185 ) );
  AOI21_X1 u2_u11_u2_U14 (.B2( u2_u11_u2_n143 ) , .ZN( u2_u11_u2_n145 ) , .B1( u2_u11_u2_n152 ) , .A( u2_u11_u2_n171 ) );
  AOI21_X1 u2_u11_u2_U15 (.B2( u2_u11_u2_n120 ) , .B1( u2_u11_u2_n121 ) , .ZN( u2_u11_u2_n126 ) , .A( u2_u11_u2_n167 ) );
  INV_X1 u2_u11_u2_U16 (.A( u2_u11_u2_n156 ) , .ZN( u2_u11_u2_n171 ) );
  INV_X1 u2_u11_u2_U17 (.A( u2_u11_u2_n120 ) , .ZN( u2_u11_u2_n188 ) );
  NAND2_X1 u2_u11_u2_U18 (.A2( u2_u11_u2_n122 ) , .ZN( u2_u11_u2_n150 ) , .A1( u2_u11_u2_n152 ) );
  INV_X1 u2_u11_u2_U19 (.A( u2_u11_u2_n153 ) , .ZN( u2_u11_u2_n170 ) );
  INV_X1 u2_u11_u2_U20 (.A( u2_u11_u2_n137 ) , .ZN( u2_u11_u2_n173 ) );
  NAND2_X1 u2_u11_u2_U21 (.A1( u2_u11_u2_n132 ) , .A2( u2_u11_u2_n139 ) , .ZN( u2_u11_u2_n157 ) );
  INV_X1 u2_u11_u2_U22 (.A( u2_u11_u2_n113 ) , .ZN( u2_u11_u2_n178 ) );
  INV_X1 u2_u11_u2_U23 (.A( u2_u11_u2_n139 ) , .ZN( u2_u11_u2_n175 ) );
  INV_X1 u2_u11_u2_U24 (.A( u2_u11_u2_n155 ) , .ZN( u2_u11_u2_n181 ) );
  INV_X1 u2_u11_u2_U25 (.A( u2_u11_u2_n119 ) , .ZN( u2_u11_u2_n177 ) );
  INV_X1 u2_u11_u2_U26 (.A( u2_u11_u2_n116 ) , .ZN( u2_u11_u2_n180 ) );
  INV_X1 u2_u11_u2_U27 (.A( u2_u11_u2_n131 ) , .ZN( u2_u11_u2_n179 ) );
  INV_X1 u2_u11_u2_U28 (.A( u2_u11_u2_n154 ) , .ZN( u2_u11_u2_n176 ) );
  NAND2_X1 u2_u11_u2_U29 (.A2( u2_u11_u2_n116 ) , .A1( u2_u11_u2_n117 ) , .ZN( u2_u11_u2_n118 ) );
  NOR2_X1 u2_u11_u2_U3 (.ZN( u2_u11_u2_n121 ) , .A2( u2_u11_u2_n177 ) , .A1( u2_u11_u2_n180 ) );
  INV_X1 u2_u11_u2_U30 (.A( u2_u11_u2_n132 ) , .ZN( u2_u11_u2_n182 ) );
  INV_X1 u2_u11_u2_U31 (.A( u2_u11_u2_n158 ) , .ZN( u2_u11_u2_n183 ) );
  OAI21_X1 u2_u11_u2_U32 (.A( u2_u11_u2_n156 ) , .B1( u2_u11_u2_n157 ) , .ZN( u2_u11_u2_n158 ) , .B2( u2_u11_u2_n179 ) );
  NOR2_X1 u2_u11_u2_U33 (.ZN( u2_u11_u2_n156 ) , .A1( u2_u11_u2_n166 ) , .A2( u2_u11_u2_n169 ) );
  NOR2_X1 u2_u11_u2_U34 (.A2( u2_u11_u2_n114 ) , .ZN( u2_u11_u2_n137 ) , .A1( u2_u11_u2_n140 ) );
  NOR2_X1 u2_u11_u2_U35 (.A2( u2_u11_u2_n138 ) , .ZN( u2_u11_u2_n153 ) , .A1( u2_u11_u2_n156 ) );
  AOI211_X1 u2_u11_u2_U36 (.ZN( u2_u11_u2_n130 ) , .C1( u2_u11_u2_n138 ) , .C2( u2_u11_u2_n179 ) , .B( u2_u11_u2_n96 ) , .A( u2_u11_u2_n97 ) );
  OAI22_X1 u2_u11_u2_U37 (.B1( u2_u11_u2_n133 ) , .A2( u2_u11_u2_n137 ) , .A1( u2_u11_u2_n152 ) , .B2( u2_u11_u2_n168 ) , .ZN( u2_u11_u2_n97 ) );
  OAI221_X1 u2_u11_u2_U38 (.B1( u2_u11_u2_n113 ) , .C1( u2_u11_u2_n132 ) , .A( u2_u11_u2_n149 ) , .B2( u2_u11_u2_n171 ) , .C2( u2_u11_u2_n172 ) , .ZN( u2_u11_u2_n96 ) );
  OAI221_X1 u2_u11_u2_U39 (.A( u2_u11_u2_n115 ) , .C2( u2_u11_u2_n123 ) , .B2( u2_u11_u2_n143 ) , .B1( u2_u11_u2_n153 ) , .ZN( u2_u11_u2_n163 ) , .C1( u2_u11_u2_n168 ) );
  INV_X1 u2_u11_u2_U4 (.A( u2_u11_u2_n134 ) , .ZN( u2_u11_u2_n185 ) );
  OAI21_X1 u2_u11_u2_U40 (.A( u2_u11_u2_n114 ) , .ZN( u2_u11_u2_n115 ) , .B1( u2_u11_u2_n176 ) , .B2( u2_u11_u2_n178 ) );
  OAI221_X1 u2_u11_u2_U41 (.A( u2_u11_u2_n135 ) , .B2( u2_u11_u2_n136 ) , .B1( u2_u11_u2_n137 ) , .ZN( u2_u11_u2_n162 ) , .C2( u2_u11_u2_n167 ) , .C1( u2_u11_u2_n185 ) );
  AND3_X1 u2_u11_u2_U42 (.A3( u2_u11_u2_n131 ) , .A2( u2_u11_u2_n132 ) , .A1( u2_u11_u2_n133 ) , .ZN( u2_u11_u2_n136 ) );
  AOI22_X1 u2_u11_u2_U43 (.ZN( u2_u11_u2_n135 ) , .B1( u2_u11_u2_n140 ) , .A1( u2_u11_u2_n156 ) , .B2( u2_u11_u2_n180 ) , .A2( u2_u11_u2_n188 ) );
  AOI21_X1 u2_u11_u2_U44 (.ZN( u2_u11_u2_n149 ) , .B1( u2_u11_u2_n173 ) , .B2( u2_u11_u2_n188 ) , .A( u2_u11_u2_n95 ) );
  AND3_X1 u2_u11_u2_U45 (.A2( u2_u11_u2_n100 ) , .A1( u2_u11_u2_n104 ) , .A3( u2_u11_u2_n156 ) , .ZN( u2_u11_u2_n95 ) );
  OAI21_X1 u2_u11_u2_U46 (.A( u2_u11_u2_n101 ) , .B2( u2_u11_u2_n121 ) , .B1( u2_u11_u2_n153 ) , .ZN( u2_u11_u2_n164 ) );
  NAND2_X1 u2_u11_u2_U47 (.A2( u2_u11_u2_n100 ) , .A1( u2_u11_u2_n107 ) , .ZN( u2_u11_u2_n155 ) );
  NAND2_X1 u2_u11_u2_U48 (.A2( u2_u11_u2_n105 ) , .A1( u2_u11_u2_n108 ) , .ZN( u2_u11_u2_n143 ) );
  NAND2_X1 u2_u11_u2_U49 (.A1( u2_u11_u2_n104 ) , .A2( u2_u11_u2_n106 ) , .ZN( u2_u11_u2_n152 ) );
  INV_X1 u2_u11_u2_U5 (.A( u2_u11_u2_n150 ) , .ZN( u2_u11_u2_n184 ) );
  NAND2_X1 u2_u11_u2_U50 (.A1( u2_u11_u2_n100 ) , .A2( u2_u11_u2_n105 ) , .ZN( u2_u11_u2_n132 ) );
  INV_X1 u2_u11_u2_U51 (.A( u2_u11_u2_n140 ) , .ZN( u2_u11_u2_n168 ) );
  INV_X1 u2_u11_u2_U52 (.A( u2_u11_u2_n138 ) , .ZN( u2_u11_u2_n167 ) );
  OAI21_X1 u2_u11_u2_U53 (.A( u2_u11_u2_n141 ) , .B2( u2_u11_u2_n142 ) , .ZN( u2_u11_u2_n146 ) , .B1( u2_u11_u2_n153 ) );
  OAI21_X1 u2_u11_u2_U54 (.A( u2_u11_u2_n140 ) , .ZN( u2_u11_u2_n141 ) , .B1( u2_u11_u2_n176 ) , .B2( u2_u11_u2_n177 ) );
  NOR3_X1 u2_u11_u2_U55 (.ZN( u2_u11_u2_n142 ) , .A3( u2_u11_u2_n175 ) , .A2( u2_u11_u2_n178 ) , .A1( u2_u11_u2_n181 ) );
  NAND2_X1 u2_u11_u2_U56 (.A1( u2_u11_u2_n102 ) , .A2( u2_u11_u2_n106 ) , .ZN( u2_u11_u2_n113 ) );
  NAND2_X1 u2_u11_u2_U57 (.A1( u2_u11_u2_n106 ) , .A2( u2_u11_u2_n107 ) , .ZN( u2_u11_u2_n131 ) );
  NAND2_X1 u2_u11_u2_U58 (.A1( u2_u11_u2_n103 ) , .A2( u2_u11_u2_n107 ) , .ZN( u2_u11_u2_n139 ) );
  NAND2_X1 u2_u11_u2_U59 (.A1( u2_u11_u2_n103 ) , .A2( u2_u11_u2_n105 ) , .ZN( u2_u11_u2_n133 ) );
  NOR4_X1 u2_u11_u2_U6 (.A4( u2_u11_u2_n124 ) , .A3( u2_u11_u2_n125 ) , .A2( u2_u11_u2_n126 ) , .A1( u2_u11_u2_n127 ) , .ZN( u2_u11_u2_n128 ) );
  NAND2_X1 u2_u11_u2_U60 (.A1( u2_u11_u2_n102 ) , .A2( u2_u11_u2_n103 ) , .ZN( u2_u11_u2_n154 ) );
  NAND2_X1 u2_u11_u2_U61 (.A2( u2_u11_u2_n103 ) , .A1( u2_u11_u2_n104 ) , .ZN( u2_u11_u2_n119 ) );
  NAND2_X1 u2_u11_u2_U62 (.A2( u2_u11_u2_n107 ) , .A1( u2_u11_u2_n108 ) , .ZN( u2_u11_u2_n123 ) );
  NAND2_X1 u2_u11_u2_U63 (.A1( u2_u11_u2_n104 ) , .A2( u2_u11_u2_n108 ) , .ZN( u2_u11_u2_n122 ) );
  INV_X1 u2_u11_u2_U64 (.A( u2_u11_u2_n114 ) , .ZN( u2_u11_u2_n172 ) );
  NAND2_X1 u2_u11_u2_U65 (.A2( u2_u11_u2_n100 ) , .A1( u2_u11_u2_n102 ) , .ZN( u2_u11_u2_n116 ) );
  NAND2_X1 u2_u11_u2_U66 (.A1( u2_u11_u2_n102 ) , .A2( u2_u11_u2_n108 ) , .ZN( u2_u11_u2_n120 ) );
  NAND2_X1 u2_u11_u2_U67 (.A2( u2_u11_u2_n105 ) , .A1( u2_u11_u2_n106 ) , .ZN( u2_u11_u2_n117 ) );
  INV_X1 u2_u11_u2_U68 (.ZN( u2_u11_u2_n187 ) , .A( u2_u11_u2_n99 ) );
  OAI21_X1 u2_u11_u2_U69 (.B1( u2_u11_u2_n137 ) , .B2( u2_u11_u2_n143 ) , .A( u2_u11_u2_n98 ) , .ZN( u2_u11_u2_n99 ) );
  AOI21_X1 u2_u11_u2_U7 (.ZN( u2_u11_u2_n124 ) , .B1( u2_u11_u2_n131 ) , .B2( u2_u11_u2_n143 ) , .A( u2_u11_u2_n172 ) );
  NOR2_X1 u2_u11_u2_U70 (.A2( u2_u11_X_16 ) , .ZN( u2_u11_u2_n140 ) , .A1( u2_u11_u2_n166 ) );
  NOR2_X1 u2_u11_u2_U71 (.A2( u2_u11_X_13 ) , .A1( u2_u11_X_14 ) , .ZN( u2_u11_u2_n100 ) );
  NOR2_X1 u2_u11_u2_U72 (.A2( u2_u11_X_16 ) , .A1( u2_u11_X_17 ) , .ZN( u2_u11_u2_n138 ) );
  NOR2_X1 u2_u11_u2_U73 (.A2( u2_u11_X_15 ) , .A1( u2_u11_X_18 ) , .ZN( u2_u11_u2_n104 ) );
  NOR2_X1 u2_u11_u2_U74 (.A2( u2_u11_X_14 ) , .ZN( u2_u11_u2_n103 ) , .A1( u2_u11_u2_n174 ) );
  NOR2_X1 u2_u11_u2_U75 (.A2( u2_u11_X_15 ) , .ZN( u2_u11_u2_n102 ) , .A1( u2_u11_u2_n165 ) );
  NOR2_X1 u2_u11_u2_U76 (.A2( u2_u11_X_17 ) , .ZN( u2_u11_u2_n114 ) , .A1( u2_u11_u2_n169 ) );
  AND2_X1 u2_u11_u2_U77 (.A1( u2_u11_X_15 ) , .ZN( u2_u11_u2_n105 ) , .A2( u2_u11_u2_n165 ) );
  AND2_X1 u2_u11_u2_U78 (.A2( u2_u11_X_15 ) , .A1( u2_u11_X_18 ) , .ZN( u2_u11_u2_n107 ) );
  AND2_X1 u2_u11_u2_U79 (.A1( u2_u11_X_14 ) , .ZN( u2_u11_u2_n106 ) , .A2( u2_u11_u2_n174 ) );
  AOI21_X1 u2_u11_u2_U8 (.B2( u2_u11_u2_n119 ) , .ZN( u2_u11_u2_n127 ) , .A( u2_u11_u2_n137 ) , .B1( u2_u11_u2_n155 ) );
  AND2_X1 u2_u11_u2_U80 (.A1( u2_u11_X_13 ) , .A2( u2_u11_X_14 ) , .ZN( u2_u11_u2_n108 ) );
  INV_X1 u2_u11_u2_U81 (.A( u2_u11_X_16 ) , .ZN( u2_u11_u2_n169 ) );
  INV_X1 u2_u11_u2_U82 (.A( u2_u11_X_17 ) , .ZN( u2_u11_u2_n166 ) );
  INV_X1 u2_u11_u2_U83 (.A( u2_u11_X_13 ) , .ZN( u2_u11_u2_n174 ) );
  INV_X1 u2_u11_u2_U84 (.A( u2_u11_X_18 ) , .ZN( u2_u11_u2_n165 ) );
  NAND4_X1 u2_u11_u2_U85 (.ZN( u2_out11_30 ) , .A4( u2_u11_u2_n147 ) , .A3( u2_u11_u2_n148 ) , .A2( u2_u11_u2_n149 ) , .A1( u2_u11_u2_n187 ) );
  NOR3_X1 u2_u11_u2_U86 (.A3( u2_u11_u2_n144 ) , .A2( u2_u11_u2_n145 ) , .A1( u2_u11_u2_n146 ) , .ZN( u2_u11_u2_n147 ) );
  AOI21_X1 u2_u11_u2_U87 (.B2( u2_u11_u2_n138 ) , .ZN( u2_u11_u2_n148 ) , .A( u2_u11_u2_n162 ) , .B1( u2_u11_u2_n182 ) );
  NAND4_X1 u2_u11_u2_U88 (.ZN( u2_out11_24 ) , .A4( u2_u11_u2_n111 ) , .A3( u2_u11_u2_n112 ) , .A1( u2_u11_u2_n130 ) , .A2( u2_u11_u2_n187 ) );
  AOI221_X1 u2_u11_u2_U89 (.A( u2_u11_u2_n109 ) , .B1( u2_u11_u2_n110 ) , .ZN( u2_u11_u2_n111 ) , .C1( u2_u11_u2_n134 ) , .C2( u2_u11_u2_n170 ) , .B2( u2_u11_u2_n173 ) );
  AOI21_X1 u2_u11_u2_U9 (.B2( u2_u11_u2_n123 ) , .ZN( u2_u11_u2_n125 ) , .A( u2_u11_u2_n171 ) , .B1( u2_u11_u2_n184 ) );
  AOI21_X1 u2_u11_u2_U90 (.ZN( u2_u11_u2_n112 ) , .B2( u2_u11_u2_n156 ) , .A( u2_u11_u2_n164 ) , .B1( u2_u11_u2_n181 ) );
  NAND4_X1 u2_u11_u2_U91 (.ZN( u2_out11_16 ) , .A4( u2_u11_u2_n128 ) , .A3( u2_u11_u2_n129 ) , .A1( u2_u11_u2_n130 ) , .A2( u2_u11_u2_n186 ) );
  AOI22_X1 u2_u11_u2_U92 (.A2( u2_u11_u2_n118 ) , .ZN( u2_u11_u2_n129 ) , .A1( u2_u11_u2_n140 ) , .B1( u2_u11_u2_n157 ) , .B2( u2_u11_u2_n170 ) );
  INV_X1 u2_u11_u2_U93 (.A( u2_u11_u2_n163 ) , .ZN( u2_u11_u2_n186 ) );
  OR4_X1 u2_u11_u2_U94 (.ZN( u2_out11_6 ) , .A4( u2_u11_u2_n161 ) , .A3( u2_u11_u2_n162 ) , .A2( u2_u11_u2_n163 ) , .A1( u2_u11_u2_n164 ) );
  OR3_X1 u2_u11_u2_U95 (.A2( u2_u11_u2_n159 ) , .A1( u2_u11_u2_n160 ) , .ZN( u2_u11_u2_n161 ) , .A3( u2_u11_u2_n183 ) );
  AOI21_X1 u2_u11_u2_U96 (.B2( u2_u11_u2_n154 ) , .B1( u2_u11_u2_n155 ) , .ZN( u2_u11_u2_n159 ) , .A( u2_u11_u2_n167 ) );
  NAND3_X1 u2_u11_u2_U97 (.A2( u2_u11_u2_n117 ) , .A1( u2_u11_u2_n122 ) , .A3( u2_u11_u2_n123 ) , .ZN( u2_u11_u2_n134 ) );
  NAND3_X1 u2_u11_u2_U98 (.ZN( u2_u11_u2_n110 ) , .A2( u2_u11_u2_n131 ) , .A3( u2_u11_u2_n139 ) , .A1( u2_u11_u2_n154 ) );
  NAND3_X1 u2_u11_u2_U99 (.A2( u2_u11_u2_n100 ) , .ZN( u2_u11_u2_n101 ) , .A1( u2_u11_u2_n104 ) , .A3( u2_u11_u2_n114 ) );
  OAI211_X1 u2_u11_u3_U10 (.B( u2_u11_u3_n106 ) , .ZN( u2_u11_u3_n119 ) , .C2( u2_u11_u3_n128 ) , .C1( u2_u11_u3_n167 ) , .A( u2_u11_u3_n181 ) );
  INV_X1 u2_u11_u3_U11 (.ZN( u2_u11_u3_n181 ) , .A( u2_u11_u3_n98 ) );
  AOI221_X1 u2_u11_u3_U12 (.C1( u2_u11_u3_n105 ) , .ZN( u2_u11_u3_n106 ) , .A( u2_u11_u3_n131 ) , .B2( u2_u11_u3_n132 ) , .C2( u2_u11_u3_n133 ) , .B1( u2_u11_u3_n169 ) );
  OAI22_X1 u2_u11_u3_U13 (.B1( u2_u11_u3_n113 ) , .A2( u2_u11_u3_n135 ) , .A1( u2_u11_u3_n150 ) , .B2( u2_u11_u3_n164 ) , .ZN( u2_u11_u3_n98 ) );
  AOI22_X1 u2_u11_u3_U14 (.B1( u2_u11_u3_n115 ) , .A2( u2_u11_u3_n116 ) , .ZN( u2_u11_u3_n123 ) , .B2( u2_u11_u3_n133 ) , .A1( u2_u11_u3_n169 ) );
  NAND2_X1 u2_u11_u3_U15 (.ZN( u2_u11_u3_n116 ) , .A2( u2_u11_u3_n151 ) , .A1( u2_u11_u3_n182 ) );
  NOR2_X1 u2_u11_u3_U16 (.ZN( u2_u11_u3_n126 ) , .A2( u2_u11_u3_n150 ) , .A1( u2_u11_u3_n164 ) );
  AOI21_X1 u2_u11_u3_U17 (.ZN( u2_u11_u3_n112 ) , .B2( u2_u11_u3_n146 ) , .B1( u2_u11_u3_n155 ) , .A( u2_u11_u3_n167 ) );
  NAND2_X1 u2_u11_u3_U18 (.A1( u2_u11_u3_n135 ) , .ZN( u2_u11_u3_n142 ) , .A2( u2_u11_u3_n164 ) );
  NAND2_X1 u2_u11_u3_U19 (.ZN( u2_u11_u3_n132 ) , .A2( u2_u11_u3_n152 ) , .A1( u2_u11_u3_n156 ) );
  INV_X1 u2_u11_u3_U20 (.A( u2_u11_u3_n133 ) , .ZN( u2_u11_u3_n165 ) );
  AND2_X1 u2_u11_u3_U21 (.A2( u2_u11_u3_n113 ) , .A1( u2_u11_u3_n114 ) , .ZN( u2_u11_u3_n151 ) );
  INV_X1 u2_u11_u3_U22 (.A( u2_u11_u3_n135 ) , .ZN( u2_u11_u3_n170 ) );
  NAND2_X1 u2_u11_u3_U23 (.A1( u2_u11_u3_n107 ) , .A2( u2_u11_u3_n108 ) , .ZN( u2_u11_u3_n140 ) );
  NAND2_X1 u2_u11_u3_U24 (.ZN( u2_u11_u3_n117 ) , .A1( u2_u11_u3_n124 ) , .A2( u2_u11_u3_n148 ) );
  NAND2_X1 u2_u11_u3_U25 (.ZN( u2_u11_u3_n143 ) , .A1( u2_u11_u3_n165 ) , .A2( u2_u11_u3_n167 ) );
  INV_X1 u2_u11_u3_U26 (.A( u2_u11_u3_n130 ) , .ZN( u2_u11_u3_n177 ) );
  INV_X1 u2_u11_u3_U27 (.A( u2_u11_u3_n128 ) , .ZN( u2_u11_u3_n176 ) );
  NAND2_X1 u2_u11_u3_U28 (.ZN( u2_u11_u3_n105 ) , .A2( u2_u11_u3_n130 ) , .A1( u2_u11_u3_n155 ) );
  INV_X1 u2_u11_u3_U29 (.A( u2_u11_u3_n155 ) , .ZN( u2_u11_u3_n174 ) );
  INV_X1 u2_u11_u3_U3 (.A( u2_u11_u3_n140 ) , .ZN( u2_u11_u3_n182 ) );
  INV_X1 u2_u11_u3_U30 (.A( u2_u11_u3_n139 ) , .ZN( u2_u11_u3_n185 ) );
  NOR2_X1 u2_u11_u3_U31 (.ZN( u2_u11_u3_n135 ) , .A2( u2_u11_u3_n141 ) , .A1( u2_u11_u3_n169 ) );
  OAI222_X1 u2_u11_u3_U32 (.C2( u2_u11_u3_n107 ) , .A2( u2_u11_u3_n108 ) , .B1( u2_u11_u3_n135 ) , .ZN( u2_u11_u3_n138 ) , .B2( u2_u11_u3_n146 ) , .C1( u2_u11_u3_n154 ) , .A1( u2_u11_u3_n164 ) );
  NOR4_X1 u2_u11_u3_U33 (.A4( u2_u11_u3_n157 ) , .A3( u2_u11_u3_n158 ) , .A2( u2_u11_u3_n159 ) , .A1( u2_u11_u3_n160 ) , .ZN( u2_u11_u3_n161 ) );
  AOI21_X1 u2_u11_u3_U34 (.B2( u2_u11_u3_n152 ) , .B1( u2_u11_u3_n153 ) , .ZN( u2_u11_u3_n158 ) , .A( u2_u11_u3_n164 ) );
  AOI21_X1 u2_u11_u3_U35 (.A( u2_u11_u3_n154 ) , .B2( u2_u11_u3_n155 ) , .B1( u2_u11_u3_n156 ) , .ZN( u2_u11_u3_n157 ) );
  AOI21_X1 u2_u11_u3_U36 (.A( u2_u11_u3_n149 ) , .B2( u2_u11_u3_n150 ) , .B1( u2_u11_u3_n151 ) , .ZN( u2_u11_u3_n159 ) );
  AOI211_X1 u2_u11_u3_U37 (.ZN( u2_u11_u3_n109 ) , .A( u2_u11_u3_n119 ) , .C2( u2_u11_u3_n129 ) , .B( u2_u11_u3_n138 ) , .C1( u2_u11_u3_n141 ) );
  AOI211_X1 u2_u11_u3_U38 (.B( u2_u11_u3_n119 ) , .A( u2_u11_u3_n120 ) , .C2( u2_u11_u3_n121 ) , .ZN( u2_u11_u3_n122 ) , .C1( u2_u11_u3_n179 ) );
  INV_X1 u2_u11_u3_U39 (.A( u2_u11_u3_n156 ) , .ZN( u2_u11_u3_n179 ) );
  INV_X1 u2_u11_u3_U4 (.A( u2_u11_u3_n129 ) , .ZN( u2_u11_u3_n183 ) );
  OAI22_X1 u2_u11_u3_U40 (.B1( u2_u11_u3_n118 ) , .ZN( u2_u11_u3_n120 ) , .A1( u2_u11_u3_n135 ) , .B2( u2_u11_u3_n154 ) , .A2( u2_u11_u3_n178 ) );
  AND3_X1 u2_u11_u3_U41 (.ZN( u2_u11_u3_n118 ) , .A2( u2_u11_u3_n124 ) , .A1( u2_u11_u3_n144 ) , .A3( u2_u11_u3_n152 ) );
  INV_X1 u2_u11_u3_U42 (.A( u2_u11_u3_n121 ) , .ZN( u2_u11_u3_n164 ) );
  NAND2_X1 u2_u11_u3_U43 (.ZN( u2_u11_u3_n133 ) , .A1( u2_u11_u3_n154 ) , .A2( u2_u11_u3_n164 ) );
  NOR2_X1 u2_u11_u3_U44 (.A1( u2_u11_u3_n113 ) , .ZN( u2_u11_u3_n131 ) , .A2( u2_u11_u3_n154 ) );
  NAND2_X1 u2_u11_u3_U45 (.A1( u2_u11_u3_n103 ) , .ZN( u2_u11_u3_n150 ) , .A2( u2_u11_u3_n99 ) );
  NAND2_X1 u2_u11_u3_U46 (.A2( u2_u11_u3_n102 ) , .ZN( u2_u11_u3_n155 ) , .A1( u2_u11_u3_n97 ) );
  OAI211_X1 u2_u11_u3_U47 (.B( u2_u11_u3_n127 ) , .ZN( u2_u11_u3_n139 ) , .C1( u2_u11_u3_n150 ) , .C2( u2_u11_u3_n154 ) , .A( u2_u11_u3_n184 ) );
  INV_X1 u2_u11_u3_U48 (.A( u2_u11_u3_n125 ) , .ZN( u2_u11_u3_n184 ) );
  AOI221_X1 u2_u11_u3_U49 (.A( u2_u11_u3_n126 ) , .ZN( u2_u11_u3_n127 ) , .C2( u2_u11_u3_n132 ) , .C1( u2_u11_u3_n169 ) , .B2( u2_u11_u3_n170 ) , .B1( u2_u11_u3_n174 ) );
  INV_X1 u2_u11_u3_U5 (.A( u2_u11_u3_n117 ) , .ZN( u2_u11_u3_n178 ) );
  OAI22_X1 u2_u11_u3_U50 (.A1( u2_u11_u3_n124 ) , .ZN( u2_u11_u3_n125 ) , .B2( u2_u11_u3_n145 ) , .A2( u2_u11_u3_n165 ) , .B1( u2_u11_u3_n167 ) );
  INV_X1 u2_u11_u3_U51 (.A( u2_u11_u3_n141 ) , .ZN( u2_u11_u3_n167 ) );
  AOI21_X1 u2_u11_u3_U52 (.B2( u2_u11_u3_n114 ) , .B1( u2_u11_u3_n146 ) , .A( u2_u11_u3_n154 ) , .ZN( u2_u11_u3_n94 ) );
  AOI21_X1 u2_u11_u3_U53 (.ZN( u2_u11_u3_n110 ) , .B2( u2_u11_u3_n142 ) , .B1( u2_u11_u3_n186 ) , .A( u2_u11_u3_n95 ) );
  INV_X1 u2_u11_u3_U54 (.A( u2_u11_u3_n145 ) , .ZN( u2_u11_u3_n186 ) );
  AOI21_X1 u2_u11_u3_U55 (.B1( u2_u11_u3_n124 ) , .A( u2_u11_u3_n149 ) , .B2( u2_u11_u3_n155 ) , .ZN( u2_u11_u3_n95 ) );
  INV_X1 u2_u11_u3_U56 (.A( u2_u11_u3_n149 ) , .ZN( u2_u11_u3_n169 ) );
  NAND2_X1 u2_u11_u3_U57 (.ZN( u2_u11_u3_n124 ) , .A1( u2_u11_u3_n96 ) , .A2( u2_u11_u3_n97 ) );
  NAND2_X1 u2_u11_u3_U58 (.A2( u2_u11_u3_n100 ) , .ZN( u2_u11_u3_n146 ) , .A1( u2_u11_u3_n96 ) );
  NAND2_X1 u2_u11_u3_U59 (.A1( u2_u11_u3_n101 ) , .ZN( u2_u11_u3_n145 ) , .A2( u2_u11_u3_n99 ) );
  AOI221_X1 u2_u11_u3_U6 (.A( u2_u11_u3_n131 ) , .C2( u2_u11_u3_n132 ) , .C1( u2_u11_u3_n133 ) , .ZN( u2_u11_u3_n134 ) , .B1( u2_u11_u3_n143 ) , .B2( u2_u11_u3_n177 ) );
  NAND2_X1 u2_u11_u3_U60 (.A1( u2_u11_u3_n100 ) , .ZN( u2_u11_u3_n156 ) , .A2( u2_u11_u3_n99 ) );
  NAND2_X1 u2_u11_u3_U61 (.A2( u2_u11_u3_n101 ) , .A1( u2_u11_u3_n104 ) , .ZN( u2_u11_u3_n148 ) );
  NAND2_X1 u2_u11_u3_U62 (.A1( u2_u11_u3_n100 ) , .A2( u2_u11_u3_n102 ) , .ZN( u2_u11_u3_n128 ) );
  NAND2_X1 u2_u11_u3_U63 (.A2( u2_u11_u3_n101 ) , .A1( u2_u11_u3_n102 ) , .ZN( u2_u11_u3_n152 ) );
  NAND2_X1 u2_u11_u3_U64 (.A2( u2_u11_u3_n101 ) , .ZN( u2_u11_u3_n114 ) , .A1( u2_u11_u3_n96 ) );
  NAND2_X1 u2_u11_u3_U65 (.ZN( u2_u11_u3_n107 ) , .A1( u2_u11_u3_n97 ) , .A2( u2_u11_u3_n99 ) );
  NAND2_X1 u2_u11_u3_U66 (.A2( u2_u11_u3_n100 ) , .A1( u2_u11_u3_n104 ) , .ZN( u2_u11_u3_n113 ) );
  NAND2_X1 u2_u11_u3_U67 (.A1( u2_u11_u3_n104 ) , .ZN( u2_u11_u3_n153 ) , .A2( u2_u11_u3_n97 ) );
  NAND2_X1 u2_u11_u3_U68 (.A2( u2_u11_u3_n103 ) , .A1( u2_u11_u3_n104 ) , .ZN( u2_u11_u3_n130 ) );
  NAND2_X1 u2_u11_u3_U69 (.A2( u2_u11_u3_n103 ) , .ZN( u2_u11_u3_n144 ) , .A1( u2_u11_u3_n96 ) );
  OAI22_X1 u2_u11_u3_U7 (.B2( u2_u11_u3_n147 ) , .A2( u2_u11_u3_n148 ) , .ZN( u2_u11_u3_n160 ) , .B1( u2_u11_u3_n165 ) , .A1( u2_u11_u3_n168 ) );
  NAND2_X1 u2_u11_u3_U70 (.A1( u2_u11_u3_n102 ) , .A2( u2_u11_u3_n103 ) , .ZN( u2_u11_u3_n108 ) );
  NOR2_X1 u2_u11_u3_U71 (.A2( u2_u11_X_19 ) , .A1( u2_u11_X_20 ) , .ZN( u2_u11_u3_n99 ) );
  NOR2_X1 u2_u11_u3_U72 (.A2( u2_u11_X_21 ) , .A1( u2_u11_X_24 ) , .ZN( u2_u11_u3_n103 ) );
  NOR2_X1 u2_u11_u3_U73 (.A2( u2_u11_X_24 ) , .A1( u2_u11_u3_n171 ) , .ZN( u2_u11_u3_n97 ) );
  NOR2_X1 u2_u11_u3_U74 (.A2( u2_u11_X_23 ) , .ZN( u2_u11_u3_n141 ) , .A1( u2_u11_u3_n166 ) );
  NOR2_X1 u2_u11_u3_U75 (.A2( u2_u11_X_19 ) , .A1( u2_u11_u3_n172 ) , .ZN( u2_u11_u3_n96 ) );
  NAND2_X1 u2_u11_u3_U76 (.A1( u2_u11_X_22 ) , .A2( u2_u11_X_23 ) , .ZN( u2_u11_u3_n154 ) );
  NAND2_X1 u2_u11_u3_U77 (.A1( u2_u11_X_23 ) , .ZN( u2_u11_u3_n149 ) , .A2( u2_u11_u3_n166 ) );
  NOR2_X1 u2_u11_u3_U78 (.A2( u2_u11_X_22 ) , .A1( u2_u11_X_23 ) , .ZN( u2_u11_u3_n121 ) );
  AND2_X1 u2_u11_u3_U79 (.A1( u2_u11_X_24 ) , .ZN( u2_u11_u3_n101 ) , .A2( u2_u11_u3_n171 ) );
  AND3_X1 u2_u11_u3_U8 (.A3( u2_u11_u3_n144 ) , .A2( u2_u11_u3_n145 ) , .A1( u2_u11_u3_n146 ) , .ZN( u2_u11_u3_n147 ) );
  AND2_X1 u2_u11_u3_U80 (.A1( u2_u11_X_19 ) , .ZN( u2_u11_u3_n102 ) , .A2( u2_u11_u3_n172 ) );
  AND2_X1 u2_u11_u3_U81 (.A1( u2_u11_X_21 ) , .A2( u2_u11_X_24 ) , .ZN( u2_u11_u3_n100 ) );
  AND2_X1 u2_u11_u3_U82 (.A2( u2_u11_X_19 ) , .A1( u2_u11_X_20 ) , .ZN( u2_u11_u3_n104 ) );
  INV_X1 u2_u11_u3_U83 (.A( u2_u11_X_22 ) , .ZN( u2_u11_u3_n166 ) );
  INV_X1 u2_u11_u3_U84 (.A( u2_u11_X_21 ) , .ZN( u2_u11_u3_n171 ) );
  INV_X1 u2_u11_u3_U85 (.A( u2_u11_X_20 ) , .ZN( u2_u11_u3_n172 ) );
  NAND4_X1 u2_u11_u3_U86 (.ZN( u2_out11_26 ) , .A4( u2_u11_u3_n109 ) , .A3( u2_u11_u3_n110 ) , .A2( u2_u11_u3_n111 ) , .A1( u2_u11_u3_n173 ) );
  INV_X1 u2_u11_u3_U87 (.ZN( u2_u11_u3_n173 ) , .A( u2_u11_u3_n94 ) );
  OAI21_X1 u2_u11_u3_U88 (.ZN( u2_u11_u3_n111 ) , .B2( u2_u11_u3_n117 ) , .A( u2_u11_u3_n133 ) , .B1( u2_u11_u3_n176 ) );
  NAND4_X1 u2_u11_u3_U89 (.ZN( u2_out11_20 ) , .A4( u2_u11_u3_n122 ) , .A3( u2_u11_u3_n123 ) , .A1( u2_u11_u3_n175 ) , .A2( u2_u11_u3_n180 ) );
  INV_X1 u2_u11_u3_U9 (.A( u2_u11_u3_n143 ) , .ZN( u2_u11_u3_n168 ) );
  INV_X1 u2_u11_u3_U90 (.A( u2_u11_u3_n126 ) , .ZN( u2_u11_u3_n180 ) );
  INV_X1 u2_u11_u3_U91 (.A( u2_u11_u3_n112 ) , .ZN( u2_u11_u3_n175 ) );
  NAND4_X1 u2_u11_u3_U92 (.ZN( u2_out11_1 ) , .A4( u2_u11_u3_n161 ) , .A3( u2_u11_u3_n162 ) , .A2( u2_u11_u3_n163 ) , .A1( u2_u11_u3_n185 ) );
  NAND2_X1 u2_u11_u3_U93 (.ZN( u2_u11_u3_n163 ) , .A2( u2_u11_u3_n170 ) , .A1( u2_u11_u3_n176 ) );
  AOI22_X1 u2_u11_u3_U94 (.B2( u2_u11_u3_n140 ) , .B1( u2_u11_u3_n141 ) , .A2( u2_u11_u3_n142 ) , .ZN( u2_u11_u3_n162 ) , .A1( u2_u11_u3_n177 ) );
  OAI222_X1 u2_u11_u3_U95 (.C1( u2_u11_u3_n128 ) , .ZN( u2_u11_u3_n137 ) , .B1( u2_u11_u3_n148 ) , .A2( u2_u11_u3_n150 ) , .B2( u2_u11_u3_n154 ) , .C2( u2_u11_u3_n164 ) , .A1( u2_u11_u3_n167 ) );
  OR4_X1 u2_u11_u3_U96 (.ZN( u2_out11_10 ) , .A4( u2_u11_u3_n136 ) , .A3( u2_u11_u3_n137 ) , .A1( u2_u11_u3_n138 ) , .A2( u2_u11_u3_n139 ) );
  OAI221_X1 u2_u11_u3_U97 (.A( u2_u11_u3_n134 ) , .B2( u2_u11_u3_n135 ) , .ZN( u2_u11_u3_n136 ) , .C1( u2_u11_u3_n149 ) , .B1( u2_u11_u3_n151 ) , .C2( u2_u11_u3_n183 ) );
  NAND3_X1 u2_u11_u3_U98 (.A1( u2_u11_u3_n114 ) , .ZN( u2_u11_u3_n115 ) , .A2( u2_u11_u3_n145 ) , .A3( u2_u11_u3_n153 ) );
  NAND3_X1 u2_u11_u3_U99 (.ZN( u2_u11_u3_n129 ) , .A2( u2_u11_u3_n144 ) , .A1( u2_u11_u3_n153 ) , .A3( u2_u11_u3_n182 ) );
  OAI22_X1 u2_u11_u4_U10 (.B2( u2_u11_u4_n135 ) , .ZN( u2_u11_u4_n137 ) , .B1( u2_u11_u4_n153 ) , .A1( u2_u11_u4_n155 ) , .A2( u2_u11_u4_n171 ) );
  AND3_X1 u2_u11_u4_U11 (.A2( u2_u11_u4_n134 ) , .ZN( u2_u11_u4_n135 ) , .A3( u2_u11_u4_n145 ) , .A1( u2_u11_u4_n157 ) );
  NAND2_X1 u2_u11_u4_U12 (.ZN( u2_u11_u4_n132 ) , .A2( u2_u11_u4_n170 ) , .A1( u2_u11_u4_n173 ) );
  AOI21_X1 u2_u11_u4_U13 (.B2( u2_u11_u4_n160 ) , .B1( u2_u11_u4_n161 ) , .ZN( u2_u11_u4_n162 ) , .A( u2_u11_u4_n170 ) );
  AOI21_X1 u2_u11_u4_U14 (.ZN( u2_u11_u4_n107 ) , .B2( u2_u11_u4_n143 ) , .A( u2_u11_u4_n174 ) , .B1( u2_u11_u4_n184 ) );
  AOI21_X1 u2_u11_u4_U15 (.B2( u2_u11_u4_n158 ) , .B1( u2_u11_u4_n159 ) , .ZN( u2_u11_u4_n163 ) , .A( u2_u11_u4_n174 ) );
  AOI21_X1 u2_u11_u4_U16 (.A( u2_u11_u4_n153 ) , .B2( u2_u11_u4_n154 ) , .B1( u2_u11_u4_n155 ) , .ZN( u2_u11_u4_n165 ) );
  AOI21_X1 u2_u11_u4_U17 (.A( u2_u11_u4_n156 ) , .B2( u2_u11_u4_n157 ) , .ZN( u2_u11_u4_n164 ) , .B1( u2_u11_u4_n184 ) );
  INV_X1 u2_u11_u4_U18 (.A( u2_u11_u4_n138 ) , .ZN( u2_u11_u4_n170 ) );
  AND2_X1 u2_u11_u4_U19 (.A2( u2_u11_u4_n120 ) , .ZN( u2_u11_u4_n155 ) , .A1( u2_u11_u4_n160 ) );
  INV_X1 u2_u11_u4_U20 (.A( u2_u11_u4_n156 ) , .ZN( u2_u11_u4_n175 ) );
  NAND2_X1 u2_u11_u4_U21 (.A2( u2_u11_u4_n118 ) , .ZN( u2_u11_u4_n131 ) , .A1( u2_u11_u4_n147 ) );
  NAND2_X1 u2_u11_u4_U22 (.A1( u2_u11_u4_n119 ) , .A2( u2_u11_u4_n120 ) , .ZN( u2_u11_u4_n130 ) );
  NAND2_X1 u2_u11_u4_U23 (.ZN( u2_u11_u4_n117 ) , .A2( u2_u11_u4_n118 ) , .A1( u2_u11_u4_n148 ) );
  NAND2_X1 u2_u11_u4_U24 (.ZN( u2_u11_u4_n129 ) , .A1( u2_u11_u4_n134 ) , .A2( u2_u11_u4_n148 ) );
  AND3_X1 u2_u11_u4_U25 (.A1( u2_u11_u4_n119 ) , .A2( u2_u11_u4_n143 ) , .A3( u2_u11_u4_n154 ) , .ZN( u2_u11_u4_n161 ) );
  AND2_X1 u2_u11_u4_U26 (.A1( u2_u11_u4_n145 ) , .A2( u2_u11_u4_n147 ) , .ZN( u2_u11_u4_n159 ) );
  OR3_X1 u2_u11_u4_U27 (.A3( u2_u11_u4_n114 ) , .A2( u2_u11_u4_n115 ) , .A1( u2_u11_u4_n116 ) , .ZN( u2_u11_u4_n136 ) );
  AOI21_X1 u2_u11_u4_U28 (.A( u2_u11_u4_n113 ) , .ZN( u2_u11_u4_n116 ) , .B2( u2_u11_u4_n173 ) , .B1( u2_u11_u4_n174 ) );
  AOI21_X1 u2_u11_u4_U29 (.ZN( u2_u11_u4_n115 ) , .B2( u2_u11_u4_n145 ) , .B1( u2_u11_u4_n146 ) , .A( u2_u11_u4_n156 ) );
  NOR2_X1 u2_u11_u4_U3 (.ZN( u2_u11_u4_n121 ) , .A1( u2_u11_u4_n181 ) , .A2( u2_u11_u4_n182 ) );
  OAI22_X1 u2_u11_u4_U30 (.ZN( u2_u11_u4_n114 ) , .A2( u2_u11_u4_n121 ) , .B1( u2_u11_u4_n160 ) , .B2( u2_u11_u4_n170 ) , .A1( u2_u11_u4_n171 ) );
  INV_X1 u2_u11_u4_U31 (.A( u2_u11_u4_n158 ) , .ZN( u2_u11_u4_n182 ) );
  INV_X1 u2_u11_u4_U32 (.ZN( u2_u11_u4_n181 ) , .A( u2_u11_u4_n96 ) );
  INV_X1 u2_u11_u4_U33 (.A( u2_u11_u4_n144 ) , .ZN( u2_u11_u4_n179 ) );
  INV_X1 u2_u11_u4_U34 (.A( u2_u11_u4_n157 ) , .ZN( u2_u11_u4_n178 ) );
  NAND2_X1 u2_u11_u4_U35 (.A2( u2_u11_u4_n154 ) , .A1( u2_u11_u4_n96 ) , .ZN( u2_u11_u4_n97 ) );
  INV_X1 u2_u11_u4_U36 (.ZN( u2_u11_u4_n186 ) , .A( u2_u11_u4_n95 ) );
  OAI221_X1 u2_u11_u4_U37 (.C1( u2_u11_u4_n134 ) , .B1( u2_u11_u4_n158 ) , .B2( u2_u11_u4_n171 ) , .C2( u2_u11_u4_n173 ) , .A( u2_u11_u4_n94 ) , .ZN( u2_u11_u4_n95 ) );
  AOI222_X1 u2_u11_u4_U38 (.B2( u2_u11_u4_n132 ) , .A1( u2_u11_u4_n138 ) , .C2( u2_u11_u4_n175 ) , .A2( u2_u11_u4_n179 ) , .C1( u2_u11_u4_n181 ) , .B1( u2_u11_u4_n185 ) , .ZN( u2_u11_u4_n94 ) );
  INV_X1 u2_u11_u4_U39 (.A( u2_u11_u4_n113 ) , .ZN( u2_u11_u4_n185 ) );
  INV_X1 u2_u11_u4_U4 (.A( u2_u11_u4_n117 ) , .ZN( u2_u11_u4_n184 ) );
  INV_X1 u2_u11_u4_U40 (.A( u2_u11_u4_n143 ) , .ZN( u2_u11_u4_n183 ) );
  NOR2_X1 u2_u11_u4_U41 (.ZN( u2_u11_u4_n138 ) , .A1( u2_u11_u4_n168 ) , .A2( u2_u11_u4_n169 ) );
  NOR2_X1 u2_u11_u4_U42 (.A1( u2_u11_u4_n150 ) , .A2( u2_u11_u4_n152 ) , .ZN( u2_u11_u4_n153 ) );
  NOR2_X1 u2_u11_u4_U43 (.A2( u2_u11_u4_n128 ) , .A1( u2_u11_u4_n138 ) , .ZN( u2_u11_u4_n156 ) );
  AOI22_X1 u2_u11_u4_U44 (.B2( u2_u11_u4_n122 ) , .A1( u2_u11_u4_n123 ) , .ZN( u2_u11_u4_n124 ) , .B1( u2_u11_u4_n128 ) , .A2( u2_u11_u4_n172 ) );
  INV_X1 u2_u11_u4_U45 (.A( u2_u11_u4_n153 ) , .ZN( u2_u11_u4_n172 ) );
  NAND2_X1 u2_u11_u4_U46 (.A2( u2_u11_u4_n120 ) , .ZN( u2_u11_u4_n123 ) , .A1( u2_u11_u4_n161 ) );
  AOI22_X1 u2_u11_u4_U47 (.B2( u2_u11_u4_n132 ) , .A2( u2_u11_u4_n133 ) , .ZN( u2_u11_u4_n140 ) , .A1( u2_u11_u4_n150 ) , .B1( u2_u11_u4_n179 ) );
  NAND2_X1 u2_u11_u4_U48 (.ZN( u2_u11_u4_n133 ) , .A2( u2_u11_u4_n146 ) , .A1( u2_u11_u4_n154 ) );
  NAND2_X1 u2_u11_u4_U49 (.A1( u2_u11_u4_n103 ) , .ZN( u2_u11_u4_n154 ) , .A2( u2_u11_u4_n98 ) );
  NOR4_X1 u2_u11_u4_U5 (.A4( u2_u11_u4_n106 ) , .A3( u2_u11_u4_n107 ) , .A2( u2_u11_u4_n108 ) , .A1( u2_u11_u4_n109 ) , .ZN( u2_u11_u4_n110 ) );
  NAND2_X1 u2_u11_u4_U50 (.A1( u2_u11_u4_n101 ) , .ZN( u2_u11_u4_n158 ) , .A2( u2_u11_u4_n99 ) );
  AOI21_X1 u2_u11_u4_U51 (.ZN( u2_u11_u4_n127 ) , .A( u2_u11_u4_n136 ) , .B2( u2_u11_u4_n150 ) , .B1( u2_u11_u4_n180 ) );
  INV_X1 u2_u11_u4_U52 (.A( u2_u11_u4_n160 ) , .ZN( u2_u11_u4_n180 ) );
  NAND2_X1 u2_u11_u4_U53 (.A2( u2_u11_u4_n104 ) , .A1( u2_u11_u4_n105 ) , .ZN( u2_u11_u4_n146 ) );
  NAND2_X1 u2_u11_u4_U54 (.A2( u2_u11_u4_n101 ) , .A1( u2_u11_u4_n102 ) , .ZN( u2_u11_u4_n160 ) );
  NAND2_X1 u2_u11_u4_U55 (.ZN( u2_u11_u4_n134 ) , .A1( u2_u11_u4_n98 ) , .A2( u2_u11_u4_n99 ) );
  NAND2_X1 u2_u11_u4_U56 (.A1( u2_u11_u4_n103 ) , .A2( u2_u11_u4_n104 ) , .ZN( u2_u11_u4_n143 ) );
  NAND2_X1 u2_u11_u4_U57 (.A2( u2_u11_u4_n105 ) , .ZN( u2_u11_u4_n145 ) , .A1( u2_u11_u4_n98 ) );
  NAND2_X1 u2_u11_u4_U58 (.A1( u2_u11_u4_n100 ) , .A2( u2_u11_u4_n105 ) , .ZN( u2_u11_u4_n120 ) );
  NAND2_X1 u2_u11_u4_U59 (.A1( u2_u11_u4_n102 ) , .A2( u2_u11_u4_n104 ) , .ZN( u2_u11_u4_n148 ) );
  AOI21_X1 u2_u11_u4_U6 (.ZN( u2_u11_u4_n106 ) , .B2( u2_u11_u4_n146 ) , .B1( u2_u11_u4_n158 ) , .A( u2_u11_u4_n170 ) );
  NAND2_X1 u2_u11_u4_U60 (.A2( u2_u11_u4_n100 ) , .A1( u2_u11_u4_n103 ) , .ZN( u2_u11_u4_n157 ) );
  INV_X1 u2_u11_u4_U61 (.A( u2_u11_u4_n150 ) , .ZN( u2_u11_u4_n173 ) );
  INV_X1 u2_u11_u4_U62 (.A( u2_u11_u4_n152 ) , .ZN( u2_u11_u4_n171 ) );
  NAND2_X1 u2_u11_u4_U63 (.A1( u2_u11_u4_n100 ) , .ZN( u2_u11_u4_n118 ) , .A2( u2_u11_u4_n99 ) );
  NAND2_X1 u2_u11_u4_U64 (.A2( u2_u11_u4_n100 ) , .A1( u2_u11_u4_n102 ) , .ZN( u2_u11_u4_n144 ) );
  NAND2_X1 u2_u11_u4_U65 (.A2( u2_u11_u4_n101 ) , .A1( u2_u11_u4_n105 ) , .ZN( u2_u11_u4_n96 ) );
  INV_X1 u2_u11_u4_U66 (.A( u2_u11_u4_n128 ) , .ZN( u2_u11_u4_n174 ) );
  NAND2_X1 u2_u11_u4_U67 (.A2( u2_u11_u4_n102 ) , .ZN( u2_u11_u4_n119 ) , .A1( u2_u11_u4_n98 ) );
  NAND2_X1 u2_u11_u4_U68 (.A2( u2_u11_u4_n101 ) , .A1( u2_u11_u4_n103 ) , .ZN( u2_u11_u4_n147 ) );
  NAND2_X1 u2_u11_u4_U69 (.A2( u2_u11_u4_n104 ) , .ZN( u2_u11_u4_n113 ) , .A1( u2_u11_u4_n99 ) );
  AOI21_X1 u2_u11_u4_U7 (.ZN( u2_u11_u4_n108 ) , .B2( u2_u11_u4_n134 ) , .B1( u2_u11_u4_n155 ) , .A( u2_u11_u4_n156 ) );
  NOR2_X1 u2_u11_u4_U70 (.A2( u2_u11_X_28 ) , .ZN( u2_u11_u4_n150 ) , .A1( u2_u11_u4_n168 ) );
  NOR2_X1 u2_u11_u4_U71 (.A2( u2_u11_X_29 ) , .ZN( u2_u11_u4_n152 ) , .A1( u2_u11_u4_n169 ) );
  NOR2_X1 u2_u11_u4_U72 (.A2( u2_u11_X_26 ) , .ZN( u2_u11_u4_n100 ) , .A1( u2_u11_u4_n177 ) );
  NOR2_X1 u2_u11_u4_U73 (.A2( u2_u11_X_30 ) , .ZN( u2_u11_u4_n105 ) , .A1( u2_u11_u4_n176 ) );
  NOR2_X1 u2_u11_u4_U74 (.A2( u2_u11_X_28 ) , .A1( u2_u11_X_29 ) , .ZN( u2_u11_u4_n128 ) );
  NOR2_X1 u2_u11_u4_U75 (.A2( u2_u11_X_25 ) , .A1( u2_u11_X_26 ) , .ZN( u2_u11_u4_n98 ) );
  NOR2_X1 u2_u11_u4_U76 (.A2( u2_u11_X_27 ) , .A1( u2_u11_X_30 ) , .ZN( u2_u11_u4_n102 ) );
  AND2_X1 u2_u11_u4_U77 (.A2( u2_u11_X_25 ) , .A1( u2_u11_X_26 ) , .ZN( u2_u11_u4_n104 ) );
  AND2_X1 u2_u11_u4_U78 (.A1( u2_u11_X_30 ) , .A2( u2_u11_u4_n176 ) , .ZN( u2_u11_u4_n99 ) );
  AND2_X1 u2_u11_u4_U79 (.A1( u2_u11_X_26 ) , .ZN( u2_u11_u4_n101 ) , .A2( u2_u11_u4_n177 ) );
  AOI21_X1 u2_u11_u4_U8 (.ZN( u2_u11_u4_n109 ) , .A( u2_u11_u4_n153 ) , .B1( u2_u11_u4_n159 ) , .B2( u2_u11_u4_n184 ) );
  AND2_X1 u2_u11_u4_U80 (.A1( u2_u11_X_27 ) , .A2( u2_u11_X_30 ) , .ZN( u2_u11_u4_n103 ) );
  INV_X1 u2_u11_u4_U81 (.A( u2_u11_X_28 ) , .ZN( u2_u11_u4_n169 ) );
  INV_X1 u2_u11_u4_U82 (.A( u2_u11_X_29 ) , .ZN( u2_u11_u4_n168 ) );
  INV_X1 u2_u11_u4_U83 (.A( u2_u11_X_25 ) , .ZN( u2_u11_u4_n177 ) );
  INV_X1 u2_u11_u4_U84 (.A( u2_u11_X_27 ) , .ZN( u2_u11_u4_n176 ) );
  NAND4_X1 u2_u11_u4_U85 (.ZN( u2_out11_25 ) , .A4( u2_u11_u4_n139 ) , .A3( u2_u11_u4_n140 ) , .A2( u2_u11_u4_n141 ) , .A1( u2_u11_u4_n142 ) );
  OAI21_X1 u2_u11_u4_U86 (.A( u2_u11_u4_n128 ) , .B2( u2_u11_u4_n129 ) , .B1( u2_u11_u4_n130 ) , .ZN( u2_u11_u4_n142 ) );
  OAI21_X1 u2_u11_u4_U87 (.B2( u2_u11_u4_n131 ) , .ZN( u2_u11_u4_n141 ) , .A( u2_u11_u4_n175 ) , .B1( u2_u11_u4_n183 ) );
  NAND4_X1 u2_u11_u4_U88 (.ZN( u2_out11_14 ) , .A4( u2_u11_u4_n124 ) , .A3( u2_u11_u4_n125 ) , .A2( u2_u11_u4_n126 ) , .A1( u2_u11_u4_n127 ) );
  AOI22_X1 u2_u11_u4_U89 (.B2( u2_u11_u4_n117 ) , .ZN( u2_u11_u4_n126 ) , .A1( u2_u11_u4_n129 ) , .B1( u2_u11_u4_n152 ) , .A2( u2_u11_u4_n175 ) );
  AOI211_X1 u2_u11_u4_U9 (.B( u2_u11_u4_n136 ) , .A( u2_u11_u4_n137 ) , .C2( u2_u11_u4_n138 ) , .ZN( u2_u11_u4_n139 ) , .C1( u2_u11_u4_n182 ) );
  AOI22_X1 u2_u11_u4_U90 (.ZN( u2_u11_u4_n125 ) , .B2( u2_u11_u4_n131 ) , .A2( u2_u11_u4_n132 ) , .B1( u2_u11_u4_n138 ) , .A1( u2_u11_u4_n178 ) );
  NAND4_X1 u2_u11_u4_U91 (.ZN( u2_out11_8 ) , .A4( u2_u11_u4_n110 ) , .A3( u2_u11_u4_n111 ) , .A2( u2_u11_u4_n112 ) , .A1( u2_u11_u4_n186 ) );
  NAND2_X1 u2_u11_u4_U92 (.ZN( u2_u11_u4_n112 ) , .A2( u2_u11_u4_n130 ) , .A1( u2_u11_u4_n150 ) );
  AOI22_X1 u2_u11_u4_U93 (.ZN( u2_u11_u4_n111 ) , .B2( u2_u11_u4_n132 ) , .A1( u2_u11_u4_n152 ) , .B1( u2_u11_u4_n178 ) , .A2( u2_u11_u4_n97 ) );
  AOI22_X1 u2_u11_u4_U94 (.B2( u2_u11_u4_n149 ) , .B1( u2_u11_u4_n150 ) , .A2( u2_u11_u4_n151 ) , .A1( u2_u11_u4_n152 ) , .ZN( u2_u11_u4_n167 ) );
  NOR4_X1 u2_u11_u4_U95 (.A4( u2_u11_u4_n162 ) , .A3( u2_u11_u4_n163 ) , .A2( u2_u11_u4_n164 ) , .A1( u2_u11_u4_n165 ) , .ZN( u2_u11_u4_n166 ) );
  NAND3_X1 u2_u11_u4_U96 (.ZN( u2_out11_3 ) , .A3( u2_u11_u4_n166 ) , .A1( u2_u11_u4_n167 ) , .A2( u2_u11_u4_n186 ) );
  NAND3_X1 u2_u11_u4_U97 (.A3( u2_u11_u4_n146 ) , .A2( u2_u11_u4_n147 ) , .A1( u2_u11_u4_n148 ) , .ZN( u2_u11_u4_n149 ) );
  NAND3_X1 u2_u11_u4_U98 (.A3( u2_u11_u4_n143 ) , .A2( u2_u11_u4_n144 ) , .A1( u2_u11_u4_n145 ) , .ZN( u2_u11_u4_n151 ) );
  NAND3_X1 u2_u11_u4_U99 (.A3( u2_u11_u4_n121 ) , .ZN( u2_u11_u4_n122 ) , .A2( u2_u11_u4_n144 ) , .A1( u2_u11_u4_n154 ) );
  INV_X1 u2_u11_u5_U10 (.A( u2_u11_u5_n121 ) , .ZN( u2_u11_u5_n177 ) );
  NOR3_X1 u2_u11_u5_U100 (.A3( u2_u11_u5_n141 ) , .A1( u2_u11_u5_n142 ) , .ZN( u2_u11_u5_n143 ) , .A2( u2_u11_u5_n191 ) );
  NAND4_X1 u2_u11_u5_U101 (.ZN( u2_out11_4 ) , .A4( u2_u11_u5_n112 ) , .A2( u2_u11_u5_n113 ) , .A1( u2_u11_u5_n114 ) , .A3( u2_u11_u5_n195 ) );
  AOI211_X1 u2_u11_u5_U102 (.A( u2_u11_u5_n110 ) , .C1( u2_u11_u5_n111 ) , .ZN( u2_u11_u5_n112 ) , .B( u2_u11_u5_n118 ) , .C2( u2_u11_u5_n177 ) );
  AOI222_X1 u2_u11_u5_U103 (.ZN( u2_u11_u5_n113 ) , .A1( u2_u11_u5_n131 ) , .C1( u2_u11_u5_n148 ) , .B2( u2_u11_u5_n174 ) , .C2( u2_u11_u5_n178 ) , .A2( u2_u11_u5_n179 ) , .B1( u2_u11_u5_n99 ) );
  NAND3_X1 u2_u11_u5_U104 (.A2( u2_u11_u5_n154 ) , .A3( u2_u11_u5_n158 ) , .A1( u2_u11_u5_n161 ) , .ZN( u2_u11_u5_n99 ) );
  NOR2_X1 u2_u11_u5_U11 (.ZN( u2_u11_u5_n160 ) , .A2( u2_u11_u5_n173 ) , .A1( u2_u11_u5_n177 ) );
  INV_X1 u2_u11_u5_U12 (.A( u2_u11_u5_n150 ) , .ZN( u2_u11_u5_n174 ) );
  AOI21_X1 u2_u11_u5_U13 (.A( u2_u11_u5_n160 ) , .B2( u2_u11_u5_n161 ) , .ZN( u2_u11_u5_n162 ) , .B1( u2_u11_u5_n192 ) );
  INV_X1 u2_u11_u5_U14 (.A( u2_u11_u5_n159 ) , .ZN( u2_u11_u5_n192 ) );
  AOI21_X1 u2_u11_u5_U15 (.A( u2_u11_u5_n156 ) , .B2( u2_u11_u5_n157 ) , .B1( u2_u11_u5_n158 ) , .ZN( u2_u11_u5_n163 ) );
  AOI21_X1 u2_u11_u5_U16 (.B2( u2_u11_u5_n139 ) , .B1( u2_u11_u5_n140 ) , .ZN( u2_u11_u5_n141 ) , .A( u2_u11_u5_n150 ) );
  OAI21_X1 u2_u11_u5_U17 (.A( u2_u11_u5_n133 ) , .B2( u2_u11_u5_n134 ) , .B1( u2_u11_u5_n135 ) , .ZN( u2_u11_u5_n142 ) );
  OAI21_X1 u2_u11_u5_U18 (.ZN( u2_u11_u5_n133 ) , .B2( u2_u11_u5_n147 ) , .A( u2_u11_u5_n173 ) , .B1( u2_u11_u5_n188 ) );
  NAND2_X1 u2_u11_u5_U19 (.A2( u2_u11_u5_n119 ) , .A1( u2_u11_u5_n123 ) , .ZN( u2_u11_u5_n137 ) );
  INV_X1 u2_u11_u5_U20 (.A( u2_u11_u5_n155 ) , .ZN( u2_u11_u5_n194 ) );
  NAND2_X1 u2_u11_u5_U21 (.A1( u2_u11_u5_n121 ) , .ZN( u2_u11_u5_n132 ) , .A2( u2_u11_u5_n172 ) );
  NAND2_X1 u2_u11_u5_U22 (.A2( u2_u11_u5_n122 ) , .ZN( u2_u11_u5_n136 ) , .A1( u2_u11_u5_n154 ) );
  NAND2_X1 u2_u11_u5_U23 (.A2( u2_u11_u5_n119 ) , .A1( u2_u11_u5_n120 ) , .ZN( u2_u11_u5_n159 ) );
  INV_X1 u2_u11_u5_U24 (.A( u2_u11_u5_n156 ) , .ZN( u2_u11_u5_n175 ) );
  INV_X1 u2_u11_u5_U25 (.A( u2_u11_u5_n158 ) , .ZN( u2_u11_u5_n188 ) );
  INV_X1 u2_u11_u5_U26 (.A( u2_u11_u5_n152 ) , .ZN( u2_u11_u5_n179 ) );
  INV_X1 u2_u11_u5_U27 (.A( u2_u11_u5_n140 ) , .ZN( u2_u11_u5_n182 ) );
  INV_X1 u2_u11_u5_U28 (.A( u2_u11_u5_n151 ) , .ZN( u2_u11_u5_n183 ) );
  INV_X1 u2_u11_u5_U29 (.A( u2_u11_u5_n123 ) , .ZN( u2_u11_u5_n185 ) );
  NOR2_X1 u2_u11_u5_U3 (.ZN( u2_u11_u5_n134 ) , .A1( u2_u11_u5_n183 ) , .A2( u2_u11_u5_n190 ) );
  INV_X1 u2_u11_u5_U30 (.A( u2_u11_u5_n161 ) , .ZN( u2_u11_u5_n184 ) );
  INV_X1 u2_u11_u5_U31 (.A( u2_u11_u5_n139 ) , .ZN( u2_u11_u5_n189 ) );
  INV_X1 u2_u11_u5_U32 (.A( u2_u11_u5_n157 ) , .ZN( u2_u11_u5_n190 ) );
  INV_X1 u2_u11_u5_U33 (.A( u2_u11_u5_n120 ) , .ZN( u2_u11_u5_n193 ) );
  NAND2_X1 u2_u11_u5_U34 (.ZN( u2_u11_u5_n111 ) , .A1( u2_u11_u5_n140 ) , .A2( u2_u11_u5_n155 ) );
  NOR2_X1 u2_u11_u5_U35 (.ZN( u2_u11_u5_n100 ) , .A1( u2_u11_u5_n170 ) , .A2( u2_u11_u5_n180 ) );
  INV_X1 u2_u11_u5_U36 (.A( u2_u11_u5_n117 ) , .ZN( u2_u11_u5_n196 ) );
  OAI221_X1 u2_u11_u5_U37 (.A( u2_u11_u5_n116 ) , .ZN( u2_u11_u5_n117 ) , .B2( u2_u11_u5_n119 ) , .C1( u2_u11_u5_n153 ) , .C2( u2_u11_u5_n158 ) , .B1( u2_u11_u5_n172 ) );
  AOI222_X1 u2_u11_u5_U38 (.ZN( u2_u11_u5_n116 ) , .B2( u2_u11_u5_n145 ) , .C1( u2_u11_u5_n148 ) , .A2( u2_u11_u5_n174 ) , .C2( u2_u11_u5_n177 ) , .B1( u2_u11_u5_n187 ) , .A1( u2_u11_u5_n193 ) );
  INV_X1 u2_u11_u5_U39 (.A( u2_u11_u5_n115 ) , .ZN( u2_u11_u5_n187 ) );
  INV_X1 u2_u11_u5_U4 (.A( u2_u11_u5_n138 ) , .ZN( u2_u11_u5_n191 ) );
  AOI22_X1 u2_u11_u5_U40 (.B2( u2_u11_u5_n131 ) , .A2( u2_u11_u5_n146 ) , .ZN( u2_u11_u5_n169 ) , .B1( u2_u11_u5_n174 ) , .A1( u2_u11_u5_n185 ) );
  NOR2_X1 u2_u11_u5_U41 (.A1( u2_u11_u5_n146 ) , .ZN( u2_u11_u5_n150 ) , .A2( u2_u11_u5_n173 ) );
  AOI21_X1 u2_u11_u5_U42 (.A( u2_u11_u5_n118 ) , .B2( u2_u11_u5_n145 ) , .ZN( u2_u11_u5_n168 ) , .B1( u2_u11_u5_n186 ) );
  INV_X1 u2_u11_u5_U43 (.A( u2_u11_u5_n122 ) , .ZN( u2_u11_u5_n186 ) );
  NOR2_X1 u2_u11_u5_U44 (.A1( u2_u11_u5_n146 ) , .ZN( u2_u11_u5_n152 ) , .A2( u2_u11_u5_n176 ) );
  NOR2_X1 u2_u11_u5_U45 (.A1( u2_u11_u5_n115 ) , .ZN( u2_u11_u5_n118 ) , .A2( u2_u11_u5_n153 ) );
  NOR2_X1 u2_u11_u5_U46 (.A2( u2_u11_u5_n145 ) , .ZN( u2_u11_u5_n156 ) , .A1( u2_u11_u5_n174 ) );
  NOR2_X1 u2_u11_u5_U47 (.ZN( u2_u11_u5_n121 ) , .A2( u2_u11_u5_n145 ) , .A1( u2_u11_u5_n176 ) );
  AOI22_X1 u2_u11_u5_U48 (.ZN( u2_u11_u5_n114 ) , .A2( u2_u11_u5_n137 ) , .A1( u2_u11_u5_n145 ) , .B2( u2_u11_u5_n175 ) , .B1( u2_u11_u5_n193 ) );
  OAI211_X1 u2_u11_u5_U49 (.B( u2_u11_u5_n124 ) , .A( u2_u11_u5_n125 ) , .C2( u2_u11_u5_n126 ) , .C1( u2_u11_u5_n127 ) , .ZN( u2_u11_u5_n128 ) );
  OAI21_X1 u2_u11_u5_U5 (.B2( u2_u11_u5_n136 ) , .B1( u2_u11_u5_n137 ) , .ZN( u2_u11_u5_n138 ) , .A( u2_u11_u5_n177 ) );
  OAI21_X1 u2_u11_u5_U50 (.ZN( u2_u11_u5_n124 ) , .A( u2_u11_u5_n177 ) , .B2( u2_u11_u5_n183 ) , .B1( u2_u11_u5_n189 ) );
  NOR3_X1 u2_u11_u5_U51 (.ZN( u2_u11_u5_n127 ) , .A1( u2_u11_u5_n136 ) , .A3( u2_u11_u5_n148 ) , .A2( u2_u11_u5_n182 ) );
  OAI21_X1 u2_u11_u5_U52 (.ZN( u2_u11_u5_n125 ) , .A( u2_u11_u5_n174 ) , .B2( u2_u11_u5_n185 ) , .B1( u2_u11_u5_n190 ) );
  AOI21_X1 u2_u11_u5_U53 (.A( u2_u11_u5_n153 ) , .B2( u2_u11_u5_n154 ) , .B1( u2_u11_u5_n155 ) , .ZN( u2_u11_u5_n164 ) );
  AOI21_X1 u2_u11_u5_U54 (.ZN( u2_u11_u5_n110 ) , .B1( u2_u11_u5_n122 ) , .B2( u2_u11_u5_n139 ) , .A( u2_u11_u5_n153 ) );
  INV_X1 u2_u11_u5_U55 (.A( u2_u11_u5_n153 ) , .ZN( u2_u11_u5_n176 ) );
  INV_X1 u2_u11_u5_U56 (.A( u2_u11_u5_n126 ) , .ZN( u2_u11_u5_n173 ) );
  AND2_X1 u2_u11_u5_U57 (.A2( u2_u11_u5_n104 ) , .A1( u2_u11_u5_n107 ) , .ZN( u2_u11_u5_n147 ) );
  AND2_X1 u2_u11_u5_U58 (.A2( u2_u11_u5_n104 ) , .A1( u2_u11_u5_n108 ) , .ZN( u2_u11_u5_n148 ) );
  NAND2_X1 u2_u11_u5_U59 (.A1( u2_u11_u5_n105 ) , .A2( u2_u11_u5_n106 ) , .ZN( u2_u11_u5_n158 ) );
  INV_X1 u2_u11_u5_U6 (.A( u2_u11_u5_n135 ) , .ZN( u2_u11_u5_n178 ) );
  NAND2_X1 u2_u11_u5_U60 (.A2( u2_u11_u5_n108 ) , .A1( u2_u11_u5_n109 ) , .ZN( u2_u11_u5_n139 ) );
  NAND2_X1 u2_u11_u5_U61 (.A1( u2_u11_u5_n106 ) , .A2( u2_u11_u5_n108 ) , .ZN( u2_u11_u5_n119 ) );
  NAND2_X1 u2_u11_u5_U62 (.A2( u2_u11_u5_n103 ) , .A1( u2_u11_u5_n105 ) , .ZN( u2_u11_u5_n140 ) );
  NAND2_X1 u2_u11_u5_U63 (.A2( u2_u11_u5_n104 ) , .A1( u2_u11_u5_n105 ) , .ZN( u2_u11_u5_n155 ) );
  NAND2_X1 u2_u11_u5_U64 (.A2( u2_u11_u5_n106 ) , .A1( u2_u11_u5_n107 ) , .ZN( u2_u11_u5_n122 ) );
  NAND2_X1 u2_u11_u5_U65 (.A2( u2_u11_u5_n100 ) , .A1( u2_u11_u5_n106 ) , .ZN( u2_u11_u5_n115 ) );
  NAND2_X1 u2_u11_u5_U66 (.A2( u2_u11_u5_n100 ) , .A1( u2_u11_u5_n103 ) , .ZN( u2_u11_u5_n161 ) );
  NAND2_X1 u2_u11_u5_U67 (.A1( u2_u11_u5_n105 ) , .A2( u2_u11_u5_n109 ) , .ZN( u2_u11_u5_n154 ) );
  INV_X1 u2_u11_u5_U68 (.A( u2_u11_u5_n146 ) , .ZN( u2_u11_u5_n172 ) );
  NAND2_X1 u2_u11_u5_U69 (.A1( u2_u11_u5_n103 ) , .A2( u2_u11_u5_n108 ) , .ZN( u2_u11_u5_n123 ) );
  OAI22_X1 u2_u11_u5_U7 (.B2( u2_u11_u5_n149 ) , .B1( u2_u11_u5_n150 ) , .A2( u2_u11_u5_n151 ) , .A1( u2_u11_u5_n152 ) , .ZN( u2_u11_u5_n165 ) );
  NAND2_X1 u2_u11_u5_U70 (.A2( u2_u11_u5_n103 ) , .A1( u2_u11_u5_n107 ) , .ZN( u2_u11_u5_n151 ) );
  NAND2_X1 u2_u11_u5_U71 (.A2( u2_u11_u5_n107 ) , .A1( u2_u11_u5_n109 ) , .ZN( u2_u11_u5_n120 ) );
  NAND2_X1 u2_u11_u5_U72 (.A2( u2_u11_u5_n100 ) , .A1( u2_u11_u5_n109 ) , .ZN( u2_u11_u5_n157 ) );
  AND2_X1 u2_u11_u5_U73 (.A2( u2_u11_u5_n100 ) , .A1( u2_u11_u5_n104 ) , .ZN( u2_u11_u5_n131 ) );
  INV_X1 u2_u11_u5_U74 (.A( u2_u11_u5_n102 ) , .ZN( u2_u11_u5_n195 ) );
  OAI221_X1 u2_u11_u5_U75 (.A( u2_u11_u5_n101 ) , .ZN( u2_u11_u5_n102 ) , .C2( u2_u11_u5_n115 ) , .C1( u2_u11_u5_n126 ) , .B1( u2_u11_u5_n134 ) , .B2( u2_u11_u5_n160 ) );
  OAI21_X1 u2_u11_u5_U76 (.ZN( u2_u11_u5_n101 ) , .B1( u2_u11_u5_n137 ) , .A( u2_u11_u5_n146 ) , .B2( u2_u11_u5_n147 ) );
  NOR2_X1 u2_u11_u5_U77 (.A2( u2_u11_X_34 ) , .A1( u2_u11_X_35 ) , .ZN( u2_u11_u5_n145 ) );
  NOR2_X1 u2_u11_u5_U78 (.A2( u2_u11_X_34 ) , .ZN( u2_u11_u5_n146 ) , .A1( u2_u11_u5_n171 ) );
  NOR2_X1 u2_u11_u5_U79 (.A2( u2_u11_X_31 ) , .A1( u2_u11_X_32 ) , .ZN( u2_u11_u5_n103 ) );
  NOR3_X1 u2_u11_u5_U8 (.A2( u2_u11_u5_n147 ) , .A1( u2_u11_u5_n148 ) , .ZN( u2_u11_u5_n149 ) , .A3( u2_u11_u5_n194 ) );
  NOR2_X1 u2_u11_u5_U80 (.A2( u2_u11_X_36 ) , .ZN( u2_u11_u5_n105 ) , .A1( u2_u11_u5_n180 ) );
  NOR2_X1 u2_u11_u5_U81 (.A2( u2_u11_X_33 ) , .ZN( u2_u11_u5_n108 ) , .A1( u2_u11_u5_n170 ) );
  NOR2_X1 u2_u11_u5_U82 (.A2( u2_u11_X_33 ) , .A1( u2_u11_X_36 ) , .ZN( u2_u11_u5_n107 ) );
  NOR2_X1 u2_u11_u5_U83 (.A2( u2_u11_X_31 ) , .ZN( u2_u11_u5_n104 ) , .A1( u2_u11_u5_n181 ) );
  NAND2_X1 u2_u11_u5_U84 (.A2( u2_u11_X_34 ) , .A1( u2_u11_X_35 ) , .ZN( u2_u11_u5_n153 ) );
  NAND2_X1 u2_u11_u5_U85 (.A1( u2_u11_X_34 ) , .ZN( u2_u11_u5_n126 ) , .A2( u2_u11_u5_n171 ) );
  AND2_X1 u2_u11_u5_U86 (.A1( u2_u11_X_31 ) , .A2( u2_u11_X_32 ) , .ZN( u2_u11_u5_n106 ) );
  AND2_X1 u2_u11_u5_U87 (.A1( u2_u11_X_31 ) , .ZN( u2_u11_u5_n109 ) , .A2( u2_u11_u5_n181 ) );
  INV_X1 u2_u11_u5_U88 (.A( u2_u11_X_33 ) , .ZN( u2_u11_u5_n180 ) );
  INV_X1 u2_u11_u5_U89 (.A( u2_u11_X_35 ) , .ZN( u2_u11_u5_n171 ) );
  NOR2_X1 u2_u11_u5_U9 (.ZN( u2_u11_u5_n135 ) , .A1( u2_u11_u5_n173 ) , .A2( u2_u11_u5_n176 ) );
  INV_X1 u2_u11_u5_U90 (.A( u2_u11_X_36 ) , .ZN( u2_u11_u5_n170 ) );
  INV_X1 u2_u11_u5_U91 (.A( u2_u11_X_32 ) , .ZN( u2_u11_u5_n181 ) );
  NAND4_X1 u2_u11_u5_U92 (.ZN( u2_out11_29 ) , .A4( u2_u11_u5_n129 ) , .A3( u2_u11_u5_n130 ) , .A2( u2_u11_u5_n168 ) , .A1( u2_u11_u5_n196 ) );
  AOI221_X1 u2_u11_u5_U93 (.A( u2_u11_u5_n128 ) , .ZN( u2_u11_u5_n129 ) , .C2( u2_u11_u5_n132 ) , .B2( u2_u11_u5_n159 ) , .B1( u2_u11_u5_n176 ) , .C1( u2_u11_u5_n184 ) );
  AOI222_X1 u2_u11_u5_U94 (.ZN( u2_u11_u5_n130 ) , .A2( u2_u11_u5_n146 ) , .B1( u2_u11_u5_n147 ) , .C2( u2_u11_u5_n175 ) , .B2( u2_u11_u5_n179 ) , .A1( u2_u11_u5_n188 ) , .C1( u2_u11_u5_n194 ) );
  NAND4_X1 u2_u11_u5_U95 (.ZN( u2_out11_19 ) , .A4( u2_u11_u5_n166 ) , .A3( u2_u11_u5_n167 ) , .A2( u2_u11_u5_n168 ) , .A1( u2_u11_u5_n169 ) );
  AOI22_X1 u2_u11_u5_U96 (.B2( u2_u11_u5_n145 ) , .A2( u2_u11_u5_n146 ) , .ZN( u2_u11_u5_n167 ) , .B1( u2_u11_u5_n182 ) , .A1( u2_u11_u5_n189 ) );
  NOR4_X1 u2_u11_u5_U97 (.A4( u2_u11_u5_n162 ) , .A3( u2_u11_u5_n163 ) , .A2( u2_u11_u5_n164 ) , .A1( u2_u11_u5_n165 ) , .ZN( u2_u11_u5_n166 ) );
  NAND4_X1 u2_u11_u5_U98 (.ZN( u2_out11_11 ) , .A4( u2_u11_u5_n143 ) , .A3( u2_u11_u5_n144 ) , .A2( u2_u11_u5_n169 ) , .A1( u2_u11_u5_n196 ) );
  AOI22_X1 u2_u11_u5_U99 (.A2( u2_u11_u5_n132 ) , .ZN( u2_u11_u5_n144 ) , .B2( u2_u11_u5_n145 ) , .B1( u2_u11_u5_n184 ) , .A1( u2_u11_u5_n194 ) );
  OAI21_X1 u2_u11_u6_U10 (.A( u2_u11_u6_n159 ) , .B1( u2_u11_u6_n169 ) , .B2( u2_u11_u6_n173 ) , .ZN( u2_u11_u6_n90 ) );
  INV_X1 u2_u11_u6_U11 (.ZN( u2_u11_u6_n172 ) , .A( u2_u11_u6_n88 ) );
  AOI22_X1 u2_u11_u6_U12 (.A2( u2_u11_u6_n151 ) , .B2( u2_u11_u6_n161 ) , .A1( u2_u11_u6_n167 ) , .B1( u2_u11_u6_n170 ) , .ZN( u2_u11_u6_n89 ) );
  AOI21_X1 u2_u11_u6_U13 (.ZN( u2_u11_u6_n106 ) , .A( u2_u11_u6_n142 ) , .B2( u2_u11_u6_n159 ) , .B1( u2_u11_u6_n164 ) );
  INV_X1 u2_u11_u6_U14 (.A( u2_u11_u6_n155 ) , .ZN( u2_u11_u6_n161 ) );
  INV_X1 u2_u11_u6_U15 (.A( u2_u11_u6_n128 ) , .ZN( u2_u11_u6_n164 ) );
  NAND2_X1 u2_u11_u6_U16 (.ZN( u2_u11_u6_n110 ) , .A1( u2_u11_u6_n122 ) , .A2( u2_u11_u6_n129 ) );
  NAND2_X1 u2_u11_u6_U17 (.ZN( u2_u11_u6_n124 ) , .A2( u2_u11_u6_n146 ) , .A1( u2_u11_u6_n148 ) );
  INV_X1 u2_u11_u6_U18 (.A( u2_u11_u6_n132 ) , .ZN( u2_u11_u6_n171 ) );
  AND2_X1 u2_u11_u6_U19 (.A1( u2_u11_u6_n100 ) , .ZN( u2_u11_u6_n130 ) , .A2( u2_u11_u6_n147 ) );
  INV_X1 u2_u11_u6_U20 (.A( u2_u11_u6_n127 ) , .ZN( u2_u11_u6_n173 ) );
  INV_X1 u2_u11_u6_U21 (.A( u2_u11_u6_n121 ) , .ZN( u2_u11_u6_n167 ) );
  INV_X1 u2_u11_u6_U22 (.A( u2_u11_u6_n100 ) , .ZN( u2_u11_u6_n169 ) );
  INV_X1 u2_u11_u6_U23 (.A( u2_u11_u6_n123 ) , .ZN( u2_u11_u6_n170 ) );
  INV_X1 u2_u11_u6_U24 (.A( u2_u11_u6_n113 ) , .ZN( u2_u11_u6_n168 ) );
  AND2_X1 u2_u11_u6_U25 (.A1( u2_u11_u6_n107 ) , .A2( u2_u11_u6_n119 ) , .ZN( u2_u11_u6_n133 ) );
  AND2_X1 u2_u11_u6_U26 (.A2( u2_u11_u6_n121 ) , .A1( u2_u11_u6_n122 ) , .ZN( u2_u11_u6_n131 ) );
  AND3_X1 u2_u11_u6_U27 (.ZN( u2_u11_u6_n120 ) , .A2( u2_u11_u6_n127 ) , .A1( u2_u11_u6_n132 ) , .A3( u2_u11_u6_n145 ) );
  INV_X1 u2_u11_u6_U28 (.A( u2_u11_u6_n146 ) , .ZN( u2_u11_u6_n163 ) );
  AOI222_X1 u2_u11_u6_U29 (.ZN( u2_u11_u6_n114 ) , .A1( u2_u11_u6_n118 ) , .A2( u2_u11_u6_n126 ) , .B2( u2_u11_u6_n151 ) , .C2( u2_u11_u6_n159 ) , .C1( u2_u11_u6_n168 ) , .B1( u2_u11_u6_n169 ) );
  INV_X1 u2_u11_u6_U3 (.A( u2_u11_u6_n110 ) , .ZN( u2_u11_u6_n166 ) );
  NOR2_X1 u2_u11_u6_U30 (.A1( u2_u11_u6_n162 ) , .A2( u2_u11_u6_n165 ) , .ZN( u2_u11_u6_n98 ) );
  NAND2_X1 u2_u11_u6_U31 (.A1( u2_u11_u6_n144 ) , .ZN( u2_u11_u6_n151 ) , .A2( u2_u11_u6_n158 ) );
  NAND2_X1 u2_u11_u6_U32 (.ZN( u2_u11_u6_n132 ) , .A1( u2_u11_u6_n91 ) , .A2( u2_u11_u6_n97 ) );
  AOI22_X1 u2_u11_u6_U33 (.B2( u2_u11_u6_n110 ) , .B1( u2_u11_u6_n111 ) , .A1( u2_u11_u6_n112 ) , .ZN( u2_u11_u6_n115 ) , .A2( u2_u11_u6_n161 ) );
  NAND4_X1 u2_u11_u6_U34 (.A3( u2_u11_u6_n109 ) , .ZN( u2_u11_u6_n112 ) , .A4( u2_u11_u6_n132 ) , .A2( u2_u11_u6_n147 ) , .A1( u2_u11_u6_n166 ) );
  NOR2_X1 u2_u11_u6_U35 (.ZN( u2_u11_u6_n109 ) , .A1( u2_u11_u6_n170 ) , .A2( u2_u11_u6_n173 ) );
  NOR2_X1 u2_u11_u6_U36 (.A2( u2_u11_u6_n126 ) , .ZN( u2_u11_u6_n155 ) , .A1( u2_u11_u6_n160 ) );
  NAND2_X1 u2_u11_u6_U37 (.ZN( u2_u11_u6_n146 ) , .A2( u2_u11_u6_n94 ) , .A1( u2_u11_u6_n99 ) );
  AOI21_X1 u2_u11_u6_U38 (.A( u2_u11_u6_n144 ) , .B2( u2_u11_u6_n145 ) , .B1( u2_u11_u6_n146 ) , .ZN( u2_u11_u6_n150 ) );
  AOI211_X1 u2_u11_u6_U39 (.B( u2_u11_u6_n134 ) , .A( u2_u11_u6_n135 ) , .C1( u2_u11_u6_n136 ) , .ZN( u2_u11_u6_n137 ) , .C2( u2_u11_u6_n151 ) );
  INV_X1 u2_u11_u6_U4 (.A( u2_u11_u6_n142 ) , .ZN( u2_u11_u6_n174 ) );
  NAND4_X1 u2_u11_u6_U40 (.A4( u2_u11_u6_n127 ) , .A3( u2_u11_u6_n128 ) , .A2( u2_u11_u6_n129 ) , .A1( u2_u11_u6_n130 ) , .ZN( u2_u11_u6_n136 ) );
  AOI21_X1 u2_u11_u6_U41 (.B2( u2_u11_u6_n132 ) , .B1( u2_u11_u6_n133 ) , .ZN( u2_u11_u6_n134 ) , .A( u2_u11_u6_n158 ) );
  AOI21_X1 u2_u11_u6_U42 (.B1( u2_u11_u6_n131 ) , .ZN( u2_u11_u6_n135 ) , .A( u2_u11_u6_n144 ) , .B2( u2_u11_u6_n146 ) );
  INV_X1 u2_u11_u6_U43 (.A( u2_u11_u6_n111 ) , .ZN( u2_u11_u6_n158 ) );
  NAND2_X1 u2_u11_u6_U44 (.ZN( u2_u11_u6_n127 ) , .A1( u2_u11_u6_n91 ) , .A2( u2_u11_u6_n92 ) );
  NAND2_X1 u2_u11_u6_U45 (.ZN( u2_u11_u6_n129 ) , .A2( u2_u11_u6_n95 ) , .A1( u2_u11_u6_n96 ) );
  INV_X1 u2_u11_u6_U46 (.A( u2_u11_u6_n144 ) , .ZN( u2_u11_u6_n159 ) );
  NAND2_X1 u2_u11_u6_U47 (.ZN( u2_u11_u6_n145 ) , .A2( u2_u11_u6_n97 ) , .A1( u2_u11_u6_n98 ) );
  NAND2_X1 u2_u11_u6_U48 (.ZN( u2_u11_u6_n148 ) , .A2( u2_u11_u6_n92 ) , .A1( u2_u11_u6_n94 ) );
  NAND2_X1 u2_u11_u6_U49 (.ZN( u2_u11_u6_n108 ) , .A2( u2_u11_u6_n139 ) , .A1( u2_u11_u6_n144 ) );
  NAND2_X1 u2_u11_u6_U5 (.A2( u2_u11_u6_n143 ) , .ZN( u2_u11_u6_n152 ) , .A1( u2_u11_u6_n166 ) );
  NAND2_X1 u2_u11_u6_U50 (.ZN( u2_u11_u6_n121 ) , .A2( u2_u11_u6_n95 ) , .A1( u2_u11_u6_n97 ) );
  NAND2_X1 u2_u11_u6_U51 (.ZN( u2_u11_u6_n107 ) , .A2( u2_u11_u6_n92 ) , .A1( u2_u11_u6_n95 ) );
  AND2_X1 u2_u11_u6_U52 (.ZN( u2_u11_u6_n118 ) , .A2( u2_u11_u6_n91 ) , .A1( u2_u11_u6_n99 ) );
  NAND2_X1 u2_u11_u6_U53 (.ZN( u2_u11_u6_n147 ) , .A2( u2_u11_u6_n98 ) , .A1( u2_u11_u6_n99 ) );
  NAND2_X1 u2_u11_u6_U54 (.ZN( u2_u11_u6_n128 ) , .A1( u2_u11_u6_n94 ) , .A2( u2_u11_u6_n96 ) );
  NAND2_X1 u2_u11_u6_U55 (.ZN( u2_u11_u6_n119 ) , .A2( u2_u11_u6_n95 ) , .A1( u2_u11_u6_n99 ) );
  NAND2_X1 u2_u11_u6_U56 (.ZN( u2_u11_u6_n123 ) , .A2( u2_u11_u6_n91 ) , .A1( u2_u11_u6_n96 ) );
  NAND2_X1 u2_u11_u6_U57 (.ZN( u2_u11_u6_n100 ) , .A2( u2_u11_u6_n92 ) , .A1( u2_u11_u6_n98 ) );
  NAND2_X1 u2_u11_u6_U58 (.ZN( u2_u11_u6_n122 ) , .A1( u2_u11_u6_n94 ) , .A2( u2_u11_u6_n97 ) );
  INV_X1 u2_u11_u6_U59 (.A( u2_u11_u6_n139 ) , .ZN( u2_u11_u6_n160 ) );
  AOI22_X1 u2_u11_u6_U6 (.B2( u2_u11_u6_n101 ) , .A1( u2_u11_u6_n102 ) , .ZN( u2_u11_u6_n103 ) , .B1( u2_u11_u6_n160 ) , .A2( u2_u11_u6_n161 ) );
  NAND2_X1 u2_u11_u6_U60 (.ZN( u2_u11_u6_n113 ) , .A1( u2_u11_u6_n96 ) , .A2( u2_u11_u6_n98 ) );
  NOR2_X1 u2_u11_u6_U61 (.A2( u2_u11_X_40 ) , .A1( u2_u11_X_41 ) , .ZN( u2_u11_u6_n126 ) );
  NOR2_X1 u2_u11_u6_U62 (.A2( u2_u11_X_39 ) , .A1( u2_u11_X_42 ) , .ZN( u2_u11_u6_n92 ) );
  NOR2_X1 u2_u11_u6_U63 (.A2( u2_u11_X_39 ) , .A1( u2_u11_u6_n156 ) , .ZN( u2_u11_u6_n97 ) );
  NOR2_X1 u2_u11_u6_U64 (.A2( u2_u11_X_38 ) , .A1( u2_u11_u6_n165 ) , .ZN( u2_u11_u6_n95 ) );
  NOR2_X1 u2_u11_u6_U65 (.A2( u2_u11_X_41 ) , .ZN( u2_u11_u6_n111 ) , .A1( u2_u11_u6_n157 ) );
  NOR2_X1 u2_u11_u6_U66 (.A2( u2_u11_X_37 ) , .A1( u2_u11_u6_n162 ) , .ZN( u2_u11_u6_n94 ) );
  NOR2_X1 u2_u11_u6_U67 (.A2( u2_u11_X_37 ) , .A1( u2_u11_X_38 ) , .ZN( u2_u11_u6_n91 ) );
  NAND2_X1 u2_u11_u6_U68 (.A1( u2_u11_X_41 ) , .ZN( u2_u11_u6_n144 ) , .A2( u2_u11_u6_n157 ) );
  NAND2_X1 u2_u11_u6_U69 (.A2( u2_u11_X_40 ) , .A1( u2_u11_X_41 ) , .ZN( u2_u11_u6_n139 ) );
  NOR2_X1 u2_u11_u6_U7 (.A1( u2_u11_u6_n118 ) , .ZN( u2_u11_u6_n143 ) , .A2( u2_u11_u6_n168 ) );
  AND2_X1 u2_u11_u6_U70 (.A1( u2_u11_X_39 ) , .A2( u2_u11_u6_n156 ) , .ZN( u2_u11_u6_n96 ) );
  AND2_X1 u2_u11_u6_U71 (.A1( u2_u11_X_39 ) , .A2( u2_u11_X_42 ) , .ZN( u2_u11_u6_n99 ) );
  INV_X1 u2_u11_u6_U72 (.A( u2_u11_X_40 ) , .ZN( u2_u11_u6_n157 ) );
  INV_X1 u2_u11_u6_U73 (.A( u2_u11_X_37 ) , .ZN( u2_u11_u6_n165 ) );
  INV_X1 u2_u11_u6_U74 (.A( u2_u11_X_38 ) , .ZN( u2_u11_u6_n162 ) );
  INV_X1 u2_u11_u6_U75 (.A( u2_u11_X_42 ) , .ZN( u2_u11_u6_n156 ) );
  NAND4_X1 u2_u11_u6_U76 (.ZN( u2_out11_32 ) , .A4( u2_u11_u6_n103 ) , .A3( u2_u11_u6_n104 ) , .A2( u2_u11_u6_n105 ) , .A1( u2_u11_u6_n106 ) );
  AOI22_X1 u2_u11_u6_U77 (.ZN( u2_u11_u6_n105 ) , .A2( u2_u11_u6_n108 ) , .A1( u2_u11_u6_n118 ) , .B2( u2_u11_u6_n126 ) , .B1( u2_u11_u6_n171 ) );
  AOI22_X1 u2_u11_u6_U78 (.ZN( u2_u11_u6_n104 ) , .A1( u2_u11_u6_n111 ) , .B1( u2_u11_u6_n124 ) , .B2( u2_u11_u6_n151 ) , .A2( u2_u11_u6_n93 ) );
  NAND4_X1 u2_u11_u6_U79 (.ZN( u2_out11_12 ) , .A4( u2_u11_u6_n114 ) , .A3( u2_u11_u6_n115 ) , .A2( u2_u11_u6_n116 ) , .A1( u2_u11_u6_n117 ) );
  AOI21_X1 u2_u11_u6_U8 (.B1( u2_u11_u6_n107 ) , .B2( u2_u11_u6_n132 ) , .A( u2_u11_u6_n158 ) , .ZN( u2_u11_u6_n88 ) );
  OAI22_X1 u2_u11_u6_U80 (.B2( u2_u11_u6_n111 ) , .ZN( u2_u11_u6_n116 ) , .B1( u2_u11_u6_n126 ) , .A2( u2_u11_u6_n164 ) , .A1( u2_u11_u6_n167 ) );
  OAI21_X1 u2_u11_u6_U81 (.A( u2_u11_u6_n108 ) , .ZN( u2_u11_u6_n117 ) , .B2( u2_u11_u6_n141 ) , .B1( u2_u11_u6_n163 ) );
  OAI211_X1 u2_u11_u6_U82 (.ZN( u2_out11_7 ) , .B( u2_u11_u6_n153 ) , .C2( u2_u11_u6_n154 ) , .C1( u2_u11_u6_n155 ) , .A( u2_u11_u6_n174 ) );
  NOR3_X1 u2_u11_u6_U83 (.A1( u2_u11_u6_n141 ) , .ZN( u2_u11_u6_n154 ) , .A3( u2_u11_u6_n164 ) , .A2( u2_u11_u6_n171 ) );
  AOI211_X1 u2_u11_u6_U84 (.B( u2_u11_u6_n149 ) , .A( u2_u11_u6_n150 ) , .C2( u2_u11_u6_n151 ) , .C1( u2_u11_u6_n152 ) , .ZN( u2_u11_u6_n153 ) );
  OAI211_X1 u2_u11_u6_U85 (.ZN( u2_out11_22 ) , .B( u2_u11_u6_n137 ) , .A( u2_u11_u6_n138 ) , .C2( u2_u11_u6_n139 ) , .C1( u2_u11_u6_n140 ) );
  AOI22_X1 u2_u11_u6_U86 (.B1( u2_u11_u6_n124 ) , .A2( u2_u11_u6_n125 ) , .A1( u2_u11_u6_n126 ) , .ZN( u2_u11_u6_n138 ) , .B2( u2_u11_u6_n161 ) );
  AND4_X1 u2_u11_u6_U87 (.A3( u2_u11_u6_n119 ) , .A1( u2_u11_u6_n120 ) , .A4( u2_u11_u6_n129 ) , .ZN( u2_u11_u6_n140 ) , .A2( u2_u11_u6_n143 ) );
  NAND3_X1 u2_u11_u6_U88 (.A2( u2_u11_u6_n123 ) , .ZN( u2_u11_u6_n125 ) , .A1( u2_u11_u6_n130 ) , .A3( u2_u11_u6_n131 ) );
  NAND3_X1 u2_u11_u6_U89 (.A3( u2_u11_u6_n133 ) , .ZN( u2_u11_u6_n141 ) , .A1( u2_u11_u6_n145 ) , .A2( u2_u11_u6_n148 ) );
  AOI21_X1 u2_u11_u6_U9 (.B2( u2_u11_u6_n147 ) , .B1( u2_u11_u6_n148 ) , .ZN( u2_u11_u6_n149 ) , .A( u2_u11_u6_n158 ) );
  NAND3_X1 u2_u11_u6_U90 (.ZN( u2_u11_u6_n101 ) , .A3( u2_u11_u6_n107 ) , .A2( u2_u11_u6_n121 ) , .A1( u2_u11_u6_n127 ) );
  NAND3_X1 u2_u11_u6_U91 (.ZN( u2_u11_u6_n102 ) , .A3( u2_u11_u6_n130 ) , .A2( u2_u11_u6_n145 ) , .A1( u2_u11_u6_n166 ) );
  NAND3_X1 u2_u11_u6_U92 (.A3( u2_u11_u6_n113 ) , .A1( u2_u11_u6_n119 ) , .A2( u2_u11_u6_n123 ) , .ZN( u2_u11_u6_n93 ) );
  NAND3_X1 u2_u11_u6_U93 (.ZN( u2_u11_u6_n142 ) , .A2( u2_u11_u6_n172 ) , .A3( u2_u11_u6_n89 ) , .A1( u2_u11_u6_n90 ) );
  AND3_X1 u2_u11_u7_U10 (.A3( u2_u11_u7_n110 ) , .A2( u2_u11_u7_n127 ) , .A1( u2_u11_u7_n132 ) , .ZN( u2_u11_u7_n92 ) );
  OAI21_X1 u2_u11_u7_U11 (.A( u2_u11_u7_n161 ) , .B1( u2_u11_u7_n168 ) , .B2( u2_u11_u7_n173 ) , .ZN( u2_u11_u7_n91 ) );
  AOI211_X1 u2_u11_u7_U12 (.A( u2_u11_u7_n117 ) , .ZN( u2_u11_u7_n118 ) , .C2( u2_u11_u7_n126 ) , .C1( u2_u11_u7_n177 ) , .B( u2_u11_u7_n180 ) );
  OAI22_X1 u2_u11_u7_U13 (.B1( u2_u11_u7_n115 ) , .ZN( u2_u11_u7_n117 ) , .A2( u2_u11_u7_n133 ) , .A1( u2_u11_u7_n137 ) , .B2( u2_u11_u7_n162 ) );
  INV_X1 u2_u11_u7_U14 (.A( u2_u11_u7_n116 ) , .ZN( u2_u11_u7_n180 ) );
  NOR3_X1 u2_u11_u7_U15 (.ZN( u2_u11_u7_n115 ) , .A3( u2_u11_u7_n145 ) , .A2( u2_u11_u7_n168 ) , .A1( u2_u11_u7_n169 ) );
  OAI211_X1 u2_u11_u7_U16 (.B( u2_u11_u7_n122 ) , .A( u2_u11_u7_n123 ) , .C2( u2_u11_u7_n124 ) , .ZN( u2_u11_u7_n154 ) , .C1( u2_u11_u7_n162 ) );
  AOI222_X1 u2_u11_u7_U17 (.ZN( u2_u11_u7_n122 ) , .C2( u2_u11_u7_n126 ) , .C1( u2_u11_u7_n145 ) , .B1( u2_u11_u7_n161 ) , .A2( u2_u11_u7_n165 ) , .B2( u2_u11_u7_n170 ) , .A1( u2_u11_u7_n176 ) );
  INV_X1 u2_u11_u7_U18 (.A( u2_u11_u7_n133 ) , .ZN( u2_u11_u7_n176 ) );
  NOR3_X1 u2_u11_u7_U19 (.A2( u2_u11_u7_n134 ) , .A1( u2_u11_u7_n135 ) , .ZN( u2_u11_u7_n136 ) , .A3( u2_u11_u7_n171 ) );
  NOR2_X1 u2_u11_u7_U20 (.A1( u2_u11_u7_n130 ) , .A2( u2_u11_u7_n134 ) , .ZN( u2_u11_u7_n153 ) );
  INV_X1 u2_u11_u7_U21 (.A( u2_u11_u7_n101 ) , .ZN( u2_u11_u7_n165 ) );
  NOR2_X1 u2_u11_u7_U22 (.ZN( u2_u11_u7_n111 ) , .A2( u2_u11_u7_n134 ) , .A1( u2_u11_u7_n169 ) );
  AOI21_X1 u2_u11_u7_U23 (.ZN( u2_u11_u7_n104 ) , .B2( u2_u11_u7_n112 ) , .B1( u2_u11_u7_n127 ) , .A( u2_u11_u7_n164 ) );
  AOI21_X1 u2_u11_u7_U24 (.ZN( u2_u11_u7_n106 ) , .B1( u2_u11_u7_n133 ) , .B2( u2_u11_u7_n146 ) , .A( u2_u11_u7_n162 ) );
  AOI21_X1 u2_u11_u7_U25 (.A( u2_u11_u7_n101 ) , .ZN( u2_u11_u7_n107 ) , .B2( u2_u11_u7_n128 ) , .B1( u2_u11_u7_n175 ) );
  INV_X1 u2_u11_u7_U26 (.A( u2_u11_u7_n138 ) , .ZN( u2_u11_u7_n171 ) );
  INV_X1 u2_u11_u7_U27 (.A( u2_u11_u7_n131 ) , .ZN( u2_u11_u7_n177 ) );
  INV_X1 u2_u11_u7_U28 (.A( u2_u11_u7_n110 ) , .ZN( u2_u11_u7_n174 ) );
  NAND2_X1 u2_u11_u7_U29 (.A1( u2_u11_u7_n129 ) , .A2( u2_u11_u7_n132 ) , .ZN( u2_u11_u7_n149 ) );
  OAI21_X1 u2_u11_u7_U3 (.ZN( u2_u11_u7_n159 ) , .A( u2_u11_u7_n165 ) , .B2( u2_u11_u7_n171 ) , .B1( u2_u11_u7_n174 ) );
  NAND2_X1 u2_u11_u7_U30 (.A1( u2_u11_u7_n113 ) , .A2( u2_u11_u7_n124 ) , .ZN( u2_u11_u7_n130 ) );
  INV_X1 u2_u11_u7_U31 (.A( u2_u11_u7_n112 ) , .ZN( u2_u11_u7_n173 ) );
  INV_X1 u2_u11_u7_U32 (.A( u2_u11_u7_n128 ) , .ZN( u2_u11_u7_n168 ) );
  INV_X1 u2_u11_u7_U33 (.A( u2_u11_u7_n148 ) , .ZN( u2_u11_u7_n169 ) );
  INV_X1 u2_u11_u7_U34 (.A( u2_u11_u7_n127 ) , .ZN( u2_u11_u7_n179 ) );
  NOR2_X1 u2_u11_u7_U35 (.ZN( u2_u11_u7_n101 ) , .A2( u2_u11_u7_n150 ) , .A1( u2_u11_u7_n156 ) );
  AOI211_X1 u2_u11_u7_U36 (.B( u2_u11_u7_n154 ) , .A( u2_u11_u7_n155 ) , .C1( u2_u11_u7_n156 ) , .ZN( u2_u11_u7_n157 ) , .C2( u2_u11_u7_n172 ) );
  INV_X1 u2_u11_u7_U37 (.A( u2_u11_u7_n153 ) , .ZN( u2_u11_u7_n172 ) );
  AOI211_X1 u2_u11_u7_U38 (.B( u2_u11_u7_n139 ) , .A( u2_u11_u7_n140 ) , .C2( u2_u11_u7_n141 ) , .ZN( u2_u11_u7_n142 ) , .C1( u2_u11_u7_n156 ) );
  AOI21_X1 u2_u11_u7_U39 (.A( u2_u11_u7_n137 ) , .B1( u2_u11_u7_n138 ) , .ZN( u2_u11_u7_n139 ) , .B2( u2_u11_u7_n146 ) );
  INV_X1 u2_u11_u7_U4 (.A( u2_u11_u7_n111 ) , .ZN( u2_u11_u7_n170 ) );
  NAND4_X1 u2_u11_u7_U40 (.A3( u2_u11_u7_n127 ) , .A2( u2_u11_u7_n128 ) , .A1( u2_u11_u7_n129 ) , .ZN( u2_u11_u7_n141 ) , .A4( u2_u11_u7_n147 ) );
  OAI22_X1 u2_u11_u7_U41 (.B1( u2_u11_u7_n136 ) , .ZN( u2_u11_u7_n140 ) , .A1( u2_u11_u7_n153 ) , .B2( u2_u11_u7_n162 ) , .A2( u2_u11_u7_n164 ) );
  AOI21_X1 u2_u11_u7_U42 (.ZN( u2_u11_u7_n123 ) , .B1( u2_u11_u7_n165 ) , .B2( u2_u11_u7_n177 ) , .A( u2_u11_u7_n97 ) );
  AOI21_X1 u2_u11_u7_U43 (.B2( u2_u11_u7_n113 ) , .B1( u2_u11_u7_n124 ) , .A( u2_u11_u7_n125 ) , .ZN( u2_u11_u7_n97 ) );
  INV_X1 u2_u11_u7_U44 (.A( u2_u11_u7_n125 ) , .ZN( u2_u11_u7_n161 ) );
  INV_X1 u2_u11_u7_U45 (.A( u2_u11_u7_n152 ) , .ZN( u2_u11_u7_n162 ) );
  AOI22_X1 u2_u11_u7_U46 (.A2( u2_u11_u7_n114 ) , .ZN( u2_u11_u7_n119 ) , .B1( u2_u11_u7_n130 ) , .A1( u2_u11_u7_n156 ) , .B2( u2_u11_u7_n165 ) );
  NAND2_X1 u2_u11_u7_U47 (.A2( u2_u11_u7_n112 ) , .ZN( u2_u11_u7_n114 ) , .A1( u2_u11_u7_n175 ) );
  AND2_X1 u2_u11_u7_U48 (.ZN( u2_u11_u7_n145 ) , .A2( u2_u11_u7_n98 ) , .A1( u2_u11_u7_n99 ) );
  NOR2_X1 u2_u11_u7_U49 (.ZN( u2_u11_u7_n137 ) , .A1( u2_u11_u7_n150 ) , .A2( u2_u11_u7_n161 ) );
  INV_X1 u2_u11_u7_U5 (.A( u2_u11_u7_n149 ) , .ZN( u2_u11_u7_n175 ) );
  AOI21_X1 u2_u11_u7_U50 (.ZN( u2_u11_u7_n105 ) , .B2( u2_u11_u7_n110 ) , .A( u2_u11_u7_n125 ) , .B1( u2_u11_u7_n147 ) );
  NAND2_X1 u2_u11_u7_U51 (.ZN( u2_u11_u7_n146 ) , .A1( u2_u11_u7_n95 ) , .A2( u2_u11_u7_n98 ) );
  NAND2_X1 u2_u11_u7_U52 (.A2( u2_u11_u7_n103 ) , .ZN( u2_u11_u7_n147 ) , .A1( u2_u11_u7_n93 ) );
  NAND2_X1 u2_u11_u7_U53 (.A1( u2_u11_u7_n103 ) , .ZN( u2_u11_u7_n127 ) , .A2( u2_u11_u7_n99 ) );
  OR2_X1 u2_u11_u7_U54 (.ZN( u2_u11_u7_n126 ) , .A2( u2_u11_u7_n152 ) , .A1( u2_u11_u7_n156 ) );
  NAND2_X1 u2_u11_u7_U55 (.A2( u2_u11_u7_n102 ) , .A1( u2_u11_u7_n103 ) , .ZN( u2_u11_u7_n133 ) );
  NAND2_X1 u2_u11_u7_U56 (.ZN( u2_u11_u7_n112 ) , .A2( u2_u11_u7_n96 ) , .A1( u2_u11_u7_n99 ) );
  NAND2_X1 u2_u11_u7_U57 (.A2( u2_u11_u7_n102 ) , .ZN( u2_u11_u7_n128 ) , .A1( u2_u11_u7_n98 ) );
  NAND2_X1 u2_u11_u7_U58 (.A1( u2_u11_u7_n100 ) , .ZN( u2_u11_u7_n113 ) , .A2( u2_u11_u7_n93 ) );
  NAND2_X1 u2_u11_u7_U59 (.A2( u2_u11_u7_n102 ) , .ZN( u2_u11_u7_n124 ) , .A1( u2_u11_u7_n96 ) );
  INV_X1 u2_u11_u7_U6 (.A( u2_u11_u7_n154 ) , .ZN( u2_u11_u7_n178 ) );
  NAND2_X1 u2_u11_u7_U60 (.ZN( u2_u11_u7_n110 ) , .A1( u2_u11_u7_n95 ) , .A2( u2_u11_u7_n96 ) );
  INV_X1 u2_u11_u7_U61 (.A( u2_u11_u7_n150 ) , .ZN( u2_u11_u7_n164 ) );
  AND2_X1 u2_u11_u7_U62 (.ZN( u2_u11_u7_n134 ) , .A1( u2_u11_u7_n93 ) , .A2( u2_u11_u7_n98 ) );
  NAND2_X1 u2_u11_u7_U63 (.A1( u2_u11_u7_n100 ) , .A2( u2_u11_u7_n102 ) , .ZN( u2_u11_u7_n129 ) );
  NAND2_X1 u2_u11_u7_U64 (.A2( u2_u11_u7_n103 ) , .ZN( u2_u11_u7_n131 ) , .A1( u2_u11_u7_n95 ) );
  NAND2_X1 u2_u11_u7_U65 (.A1( u2_u11_u7_n100 ) , .ZN( u2_u11_u7_n138 ) , .A2( u2_u11_u7_n99 ) );
  NAND2_X1 u2_u11_u7_U66 (.ZN( u2_u11_u7_n132 ) , .A1( u2_u11_u7_n93 ) , .A2( u2_u11_u7_n96 ) );
  NAND2_X1 u2_u11_u7_U67 (.A1( u2_u11_u7_n100 ) , .ZN( u2_u11_u7_n148 ) , .A2( u2_u11_u7_n95 ) );
  NOR2_X1 u2_u11_u7_U68 (.A2( u2_u11_X_47 ) , .ZN( u2_u11_u7_n150 ) , .A1( u2_u11_u7_n163 ) );
  NOR2_X1 u2_u11_u7_U69 (.A2( u2_u11_X_43 ) , .A1( u2_u11_X_44 ) , .ZN( u2_u11_u7_n103 ) );
  AOI211_X1 u2_u11_u7_U7 (.ZN( u2_u11_u7_n116 ) , .A( u2_u11_u7_n155 ) , .C1( u2_u11_u7_n161 ) , .C2( u2_u11_u7_n171 ) , .B( u2_u11_u7_n94 ) );
  NOR2_X1 u2_u11_u7_U70 (.A2( u2_u11_X_48 ) , .A1( u2_u11_u7_n166 ) , .ZN( u2_u11_u7_n95 ) );
  NOR2_X1 u2_u11_u7_U71 (.A2( u2_u11_X_45 ) , .A1( u2_u11_X_48 ) , .ZN( u2_u11_u7_n99 ) );
  NOR2_X1 u2_u11_u7_U72 (.A2( u2_u11_X_44 ) , .A1( u2_u11_u7_n167 ) , .ZN( u2_u11_u7_n98 ) );
  NOR2_X1 u2_u11_u7_U73 (.A2( u2_u11_X_46 ) , .A1( u2_u11_X_47 ) , .ZN( u2_u11_u7_n152 ) );
  AND2_X1 u2_u11_u7_U74 (.A1( u2_u11_X_47 ) , .ZN( u2_u11_u7_n156 ) , .A2( u2_u11_u7_n163 ) );
  NAND2_X1 u2_u11_u7_U75 (.A2( u2_u11_X_46 ) , .A1( u2_u11_X_47 ) , .ZN( u2_u11_u7_n125 ) );
  AND2_X1 u2_u11_u7_U76 (.A2( u2_u11_X_45 ) , .A1( u2_u11_X_48 ) , .ZN( u2_u11_u7_n102 ) );
  AND2_X1 u2_u11_u7_U77 (.A2( u2_u11_X_43 ) , .A1( u2_u11_X_44 ) , .ZN( u2_u11_u7_n96 ) );
  AND2_X1 u2_u11_u7_U78 (.A1( u2_u11_X_44 ) , .ZN( u2_u11_u7_n100 ) , .A2( u2_u11_u7_n167 ) );
  AND2_X1 u2_u11_u7_U79 (.A1( u2_u11_X_48 ) , .A2( u2_u11_u7_n166 ) , .ZN( u2_u11_u7_n93 ) );
  OAI222_X1 u2_u11_u7_U8 (.C2( u2_u11_u7_n101 ) , .B2( u2_u11_u7_n111 ) , .A1( u2_u11_u7_n113 ) , .C1( u2_u11_u7_n146 ) , .A2( u2_u11_u7_n162 ) , .B1( u2_u11_u7_n164 ) , .ZN( u2_u11_u7_n94 ) );
  INV_X1 u2_u11_u7_U80 (.A( u2_u11_X_46 ) , .ZN( u2_u11_u7_n163 ) );
  INV_X1 u2_u11_u7_U81 (.A( u2_u11_X_43 ) , .ZN( u2_u11_u7_n167 ) );
  INV_X1 u2_u11_u7_U82 (.A( u2_u11_X_45 ) , .ZN( u2_u11_u7_n166 ) );
  NAND4_X1 u2_u11_u7_U83 (.ZN( u2_out11_27 ) , .A4( u2_u11_u7_n118 ) , .A3( u2_u11_u7_n119 ) , .A2( u2_u11_u7_n120 ) , .A1( u2_u11_u7_n121 ) );
  OAI21_X1 u2_u11_u7_U84 (.ZN( u2_u11_u7_n121 ) , .B2( u2_u11_u7_n145 ) , .A( u2_u11_u7_n150 ) , .B1( u2_u11_u7_n174 ) );
  OAI21_X1 u2_u11_u7_U85 (.ZN( u2_u11_u7_n120 ) , .A( u2_u11_u7_n161 ) , .B2( u2_u11_u7_n170 ) , .B1( u2_u11_u7_n179 ) );
  NAND4_X1 u2_u11_u7_U86 (.ZN( u2_out11_21 ) , .A4( u2_u11_u7_n157 ) , .A3( u2_u11_u7_n158 ) , .A2( u2_u11_u7_n159 ) , .A1( u2_u11_u7_n160 ) );
  OAI21_X1 u2_u11_u7_U87 (.B1( u2_u11_u7_n145 ) , .ZN( u2_u11_u7_n160 ) , .A( u2_u11_u7_n161 ) , .B2( u2_u11_u7_n177 ) );
  AOI22_X1 u2_u11_u7_U88 (.B2( u2_u11_u7_n149 ) , .B1( u2_u11_u7_n150 ) , .A2( u2_u11_u7_n151 ) , .A1( u2_u11_u7_n152 ) , .ZN( u2_u11_u7_n158 ) );
  NAND4_X1 u2_u11_u7_U89 (.ZN( u2_out11_15 ) , .A4( u2_u11_u7_n142 ) , .A3( u2_u11_u7_n143 ) , .A2( u2_u11_u7_n144 ) , .A1( u2_u11_u7_n178 ) );
  OAI221_X1 u2_u11_u7_U9 (.C1( u2_u11_u7_n101 ) , .C2( u2_u11_u7_n147 ) , .ZN( u2_u11_u7_n155 ) , .B2( u2_u11_u7_n162 ) , .A( u2_u11_u7_n91 ) , .B1( u2_u11_u7_n92 ) );
  OR2_X1 u2_u11_u7_U90 (.A2( u2_u11_u7_n125 ) , .A1( u2_u11_u7_n129 ) , .ZN( u2_u11_u7_n144 ) );
  AOI22_X1 u2_u11_u7_U91 (.A2( u2_u11_u7_n126 ) , .ZN( u2_u11_u7_n143 ) , .B2( u2_u11_u7_n165 ) , .B1( u2_u11_u7_n173 ) , .A1( u2_u11_u7_n174 ) );
  NAND4_X1 u2_u11_u7_U92 (.ZN( u2_out11_5 ) , .A4( u2_u11_u7_n108 ) , .A3( u2_u11_u7_n109 ) , .A1( u2_u11_u7_n116 ) , .A2( u2_u11_u7_n123 ) );
  AOI22_X1 u2_u11_u7_U93 (.ZN( u2_u11_u7_n109 ) , .A2( u2_u11_u7_n126 ) , .B2( u2_u11_u7_n145 ) , .B1( u2_u11_u7_n156 ) , .A1( u2_u11_u7_n171 ) );
  NOR4_X1 u2_u11_u7_U94 (.A4( u2_u11_u7_n104 ) , .A3( u2_u11_u7_n105 ) , .A2( u2_u11_u7_n106 ) , .A1( u2_u11_u7_n107 ) , .ZN( u2_u11_u7_n108 ) );
  NAND3_X1 u2_u11_u7_U95 (.A3( u2_u11_u7_n146 ) , .A2( u2_u11_u7_n147 ) , .A1( u2_u11_u7_n148 ) , .ZN( u2_u11_u7_n151 ) );
  NAND3_X1 u2_u11_u7_U96 (.A3( u2_u11_u7_n131 ) , .A2( u2_u11_u7_n132 ) , .A1( u2_u11_u7_n133 ) , .ZN( u2_u11_u7_n135 ) );
  XOR2_X1 u2_u12_U19 (.B( u2_K13_37 ) , .A( u2_R11_24 ) , .Z( u2_u12_X_37 ) );
  XOR2_X1 u2_u12_U21 (.B( u2_K13_35 ) , .A( u2_R11_24 ) , .Z( u2_u12_X_35 ) );
  XOR2_X1 u2_u12_U24 (.B( u2_K13_32 ) , .A( u2_R11_21 ) , .Z( u2_u12_X_32 ) );
  XOR2_X1 u2_u12_U26 (.B( u2_K13_30 ) , .A( u2_R11_21 ) , .Z( u2_u12_X_30 ) );
  XOR2_X1 u2_u12_U27 (.B( u2_K13_2 ) , .A( u2_R11_1 ) , .Z( u2_u12_X_2 ) );
  XOR2_X1 u2_u12_U3 (.B( u2_K13_7 ) , .A( u2_R11_4 ) , .Z( u2_u12_X_7 ) );
  XOR2_X1 u2_u12_U5 (.B( u2_K13_5 ) , .A( u2_R11_4 ) , .Z( u2_u12_X_5 ) );
  XOR2_X1 u2_u12_U7 (.B( u2_K13_48 ) , .A( u2_R11_1 ) , .Z( u2_u12_X_48 ) );
  AND2_X1 u2_u12_u0_U10 (.A1( u2_u12_u0_n131 ) , .ZN( u2_u12_u0_n141 ) , .A2( u2_u12_u0_n150 ) );
  AND3_X1 u2_u12_u0_U11 (.A2( u2_u12_u0_n112 ) , .ZN( u2_u12_u0_n127 ) , .A3( u2_u12_u0_n130 ) , .A1( u2_u12_u0_n148 ) );
  AND2_X1 u2_u12_u0_U12 (.ZN( u2_u12_u0_n107 ) , .A1( u2_u12_u0_n130 ) , .A2( u2_u12_u0_n140 ) );
  AND2_X1 u2_u12_u0_U13 (.A2( u2_u12_u0_n129 ) , .A1( u2_u12_u0_n130 ) , .ZN( u2_u12_u0_n151 ) );
  AND2_X1 u2_u12_u0_U14 (.A1( u2_u12_u0_n108 ) , .A2( u2_u12_u0_n125 ) , .ZN( u2_u12_u0_n145 ) );
  INV_X1 u2_u12_u0_U15 (.A( u2_u12_u0_n143 ) , .ZN( u2_u12_u0_n173 ) );
  NOR2_X1 u2_u12_u0_U16 (.A2( u2_u12_u0_n136 ) , .ZN( u2_u12_u0_n147 ) , .A1( u2_u12_u0_n160 ) );
  AOI21_X1 u2_u12_u0_U17 (.B1( u2_u12_u0_n103 ) , .ZN( u2_u12_u0_n132 ) , .A( u2_u12_u0_n165 ) , .B2( u2_u12_u0_n93 ) );
  OAI22_X1 u2_u12_u0_U18 (.B1( u2_u12_u0_n125 ) , .ZN( u2_u12_u0_n126 ) , .A1( u2_u12_u0_n138 ) , .A2( u2_u12_u0_n146 ) , .B2( u2_u12_u0_n147 ) );
  OAI22_X1 u2_u12_u0_U19 (.B1( u2_u12_u0_n131 ) , .A1( u2_u12_u0_n144 ) , .B2( u2_u12_u0_n147 ) , .A2( u2_u12_u0_n90 ) , .ZN( u2_u12_u0_n91 ) );
  AND3_X1 u2_u12_u0_U20 (.A3( u2_u12_u0_n121 ) , .A2( u2_u12_u0_n125 ) , .A1( u2_u12_u0_n148 ) , .ZN( u2_u12_u0_n90 ) );
  NOR2_X1 u2_u12_u0_U21 (.A1( u2_u12_u0_n163 ) , .A2( u2_u12_u0_n164 ) , .ZN( u2_u12_u0_n95 ) );
  AOI22_X1 u2_u12_u0_U22 (.B2( u2_u12_u0_n109 ) , .A2( u2_u12_u0_n110 ) , .ZN( u2_u12_u0_n111 ) , .B1( u2_u12_u0_n118 ) , .A1( u2_u12_u0_n160 ) );
  NAND2_X1 u2_u12_u0_U23 (.A1( u2_u12_u0_n100 ) , .A2( u2_u12_u0_n103 ) , .ZN( u2_u12_u0_n125 ) );
  INV_X1 u2_u12_u0_U24 (.A( u2_u12_u0_n136 ) , .ZN( u2_u12_u0_n161 ) );
  INV_X1 u2_u12_u0_U25 (.A( u2_u12_u0_n118 ) , .ZN( u2_u12_u0_n158 ) );
  AOI21_X1 u2_u12_u0_U26 (.B1( u2_u12_u0_n127 ) , .B2( u2_u12_u0_n129 ) , .A( u2_u12_u0_n138 ) , .ZN( u2_u12_u0_n96 ) );
  AOI21_X1 u2_u12_u0_U27 (.ZN( u2_u12_u0_n104 ) , .B1( u2_u12_u0_n107 ) , .B2( u2_u12_u0_n141 ) , .A( u2_u12_u0_n144 ) );
  NAND2_X1 u2_u12_u0_U28 (.A2( u2_u12_u0_n102 ) , .A1( u2_u12_u0_n103 ) , .ZN( u2_u12_u0_n149 ) );
  NAND2_X1 u2_u12_u0_U29 (.A2( u2_u12_u0_n100 ) , .ZN( u2_u12_u0_n131 ) , .A1( u2_u12_u0_n92 ) );
  INV_X1 u2_u12_u0_U3 (.A( u2_u12_u0_n113 ) , .ZN( u2_u12_u0_n166 ) );
  NAND2_X1 u2_u12_u0_U30 (.A2( u2_u12_u0_n102 ) , .ZN( u2_u12_u0_n114 ) , .A1( u2_u12_u0_n92 ) );
  NOR2_X1 u2_u12_u0_U31 (.A1( u2_u12_u0_n120 ) , .ZN( u2_u12_u0_n143 ) , .A2( u2_u12_u0_n167 ) );
  OAI221_X1 u2_u12_u0_U32 (.C1( u2_u12_u0_n112 ) , .ZN( u2_u12_u0_n120 ) , .B1( u2_u12_u0_n138 ) , .B2( u2_u12_u0_n141 ) , .C2( u2_u12_u0_n147 ) , .A( u2_u12_u0_n172 ) );
  AOI211_X1 u2_u12_u0_U33 (.B( u2_u12_u0_n115 ) , .A( u2_u12_u0_n116 ) , .C2( u2_u12_u0_n117 ) , .C1( u2_u12_u0_n118 ) , .ZN( u2_u12_u0_n119 ) );
  NAND2_X1 u2_u12_u0_U34 (.A1( u2_u12_u0_n101 ) , .A2( u2_u12_u0_n102 ) , .ZN( u2_u12_u0_n150 ) );
  INV_X1 u2_u12_u0_U35 (.A( u2_u12_u0_n138 ) , .ZN( u2_u12_u0_n160 ) );
  NAND2_X1 u2_u12_u0_U36 (.A2( u2_u12_u0_n100 ) , .A1( u2_u12_u0_n101 ) , .ZN( u2_u12_u0_n139 ) );
  NAND2_X1 u2_u12_u0_U37 (.ZN( u2_u12_u0_n112 ) , .A2( u2_u12_u0_n92 ) , .A1( u2_u12_u0_n93 ) );
  INV_X1 u2_u12_u0_U38 (.ZN( u2_u12_u0_n172 ) , .A( u2_u12_u0_n88 ) );
  OAI222_X1 u2_u12_u0_U39 (.C1( u2_u12_u0_n108 ) , .A1( u2_u12_u0_n125 ) , .B2( u2_u12_u0_n128 ) , .B1( u2_u12_u0_n144 ) , .A2( u2_u12_u0_n158 ) , .C2( u2_u12_u0_n161 ) , .ZN( u2_u12_u0_n88 ) );
  AOI21_X1 u2_u12_u0_U4 (.B1( u2_u12_u0_n114 ) , .ZN( u2_u12_u0_n115 ) , .B2( u2_u12_u0_n129 ) , .A( u2_u12_u0_n161 ) );
  NAND2_X1 u2_u12_u0_U40 (.A2( u2_u12_u0_n101 ) , .ZN( u2_u12_u0_n121 ) , .A1( u2_u12_u0_n93 ) );
  OR3_X1 u2_u12_u0_U41 (.A3( u2_u12_u0_n152 ) , .A2( u2_u12_u0_n153 ) , .A1( u2_u12_u0_n154 ) , .ZN( u2_u12_u0_n155 ) );
  AOI21_X1 u2_u12_u0_U42 (.B2( u2_u12_u0_n150 ) , .B1( u2_u12_u0_n151 ) , .ZN( u2_u12_u0_n152 ) , .A( u2_u12_u0_n158 ) );
  AOI21_X1 u2_u12_u0_U43 (.A( u2_u12_u0_n144 ) , .B2( u2_u12_u0_n145 ) , .B1( u2_u12_u0_n146 ) , .ZN( u2_u12_u0_n154 ) );
  AOI21_X1 u2_u12_u0_U44 (.A( u2_u12_u0_n147 ) , .B2( u2_u12_u0_n148 ) , .B1( u2_u12_u0_n149 ) , .ZN( u2_u12_u0_n153 ) );
  INV_X1 u2_u12_u0_U45 (.ZN( u2_u12_u0_n171 ) , .A( u2_u12_u0_n99 ) );
  OAI211_X1 u2_u12_u0_U46 (.C2( u2_u12_u0_n140 ) , .C1( u2_u12_u0_n161 ) , .A( u2_u12_u0_n169 ) , .B( u2_u12_u0_n98 ) , .ZN( u2_u12_u0_n99 ) );
  INV_X1 u2_u12_u0_U47 (.ZN( u2_u12_u0_n169 ) , .A( u2_u12_u0_n91 ) );
  AOI211_X1 u2_u12_u0_U48 (.C1( u2_u12_u0_n118 ) , .A( u2_u12_u0_n123 ) , .B( u2_u12_u0_n96 ) , .C2( u2_u12_u0_n97 ) , .ZN( u2_u12_u0_n98 ) );
  NOR2_X1 u2_u12_u0_U49 (.A2( u2_u12_X_4 ) , .A1( u2_u12_X_5 ) , .ZN( u2_u12_u0_n118 ) );
  NOR2_X1 u2_u12_u0_U5 (.A1( u2_u12_u0_n108 ) , .ZN( u2_u12_u0_n123 ) , .A2( u2_u12_u0_n158 ) );
  NOR2_X1 u2_u12_u0_U50 (.A2( u2_u12_X_1 ) , .ZN( u2_u12_u0_n101 ) , .A1( u2_u12_u0_n163 ) );
  NAND2_X1 u2_u12_u0_U51 (.A2( u2_u12_X_4 ) , .A1( u2_u12_X_5 ) , .ZN( u2_u12_u0_n144 ) );
  NOR2_X1 u2_u12_u0_U52 (.A2( u2_u12_X_5 ) , .ZN( u2_u12_u0_n136 ) , .A1( u2_u12_u0_n159 ) );
  NAND2_X1 u2_u12_u0_U53 (.A1( u2_u12_X_5 ) , .ZN( u2_u12_u0_n138 ) , .A2( u2_u12_u0_n159 ) );
  AND2_X1 u2_u12_u0_U54 (.A2( u2_u12_X_3 ) , .A1( u2_u12_X_6 ) , .ZN( u2_u12_u0_n102 ) );
  INV_X1 u2_u12_u0_U55 (.A( u2_u12_X_4 ) , .ZN( u2_u12_u0_n159 ) );
  INV_X1 u2_u12_u0_U56 (.A( u2_u12_X_1 ) , .ZN( u2_u12_u0_n164 ) );
  INV_X1 u2_u12_u0_U57 (.A( u2_u12_X_3 ) , .ZN( u2_u12_u0_n162 ) );
  INV_X1 u2_u12_u0_U58 (.A( u2_u12_u0_n126 ) , .ZN( u2_u12_u0_n168 ) );
  AOI211_X1 u2_u12_u0_U59 (.B( u2_u12_u0_n133 ) , .A( u2_u12_u0_n134 ) , .C2( u2_u12_u0_n135 ) , .C1( u2_u12_u0_n136 ) , .ZN( u2_u12_u0_n137 ) );
  AOI21_X1 u2_u12_u0_U6 (.B2( u2_u12_u0_n131 ) , .ZN( u2_u12_u0_n134 ) , .B1( u2_u12_u0_n151 ) , .A( u2_u12_u0_n158 ) );
  OR4_X1 u2_u12_u0_U60 (.ZN( u2_out12_17 ) , .A4( u2_u12_u0_n122 ) , .A2( u2_u12_u0_n123 ) , .A1( u2_u12_u0_n124 ) , .A3( u2_u12_u0_n170 ) );
  AOI21_X1 u2_u12_u0_U61 (.B2( u2_u12_u0_n107 ) , .ZN( u2_u12_u0_n124 ) , .B1( u2_u12_u0_n128 ) , .A( u2_u12_u0_n161 ) );
  INV_X1 u2_u12_u0_U62 (.A( u2_u12_u0_n111 ) , .ZN( u2_u12_u0_n170 ) );
  OR4_X1 u2_u12_u0_U63 (.ZN( u2_out12_31 ) , .A4( u2_u12_u0_n155 ) , .A2( u2_u12_u0_n156 ) , .A1( u2_u12_u0_n157 ) , .A3( u2_u12_u0_n173 ) );
  AOI21_X1 u2_u12_u0_U64 (.A( u2_u12_u0_n138 ) , .B2( u2_u12_u0_n139 ) , .B1( u2_u12_u0_n140 ) , .ZN( u2_u12_u0_n157 ) );
  INV_X1 u2_u12_u0_U65 (.ZN( u2_u12_u0_n174 ) , .A( u2_u12_u0_n89 ) );
  AOI211_X1 u2_u12_u0_U66 (.B( u2_u12_u0_n104 ) , .A( u2_u12_u0_n105 ) , .ZN( u2_u12_u0_n106 ) , .C2( u2_u12_u0_n113 ) , .C1( u2_u12_u0_n160 ) );
  AOI21_X1 u2_u12_u0_U67 (.B2( u2_u12_u0_n141 ) , .B1( u2_u12_u0_n142 ) , .ZN( u2_u12_u0_n156 ) , .A( u2_u12_u0_n161 ) );
  AOI21_X1 u2_u12_u0_U68 (.ZN( u2_u12_u0_n116 ) , .B2( u2_u12_u0_n142 ) , .A( u2_u12_u0_n144 ) , .B1( u2_u12_u0_n166 ) );
  INV_X1 u2_u12_u0_U69 (.A( u2_u12_u0_n142 ) , .ZN( u2_u12_u0_n165 ) );
  OAI21_X1 u2_u12_u0_U7 (.B1( u2_u12_u0_n150 ) , .B2( u2_u12_u0_n158 ) , .A( u2_u12_u0_n172 ) , .ZN( u2_u12_u0_n89 ) );
  NAND2_X1 u2_u12_u0_U70 (.A2( u2_u12_u0_n103 ) , .ZN( u2_u12_u0_n140 ) , .A1( u2_u12_u0_n94 ) );
  NAND2_X1 u2_u12_u0_U71 (.A1( u2_u12_u0_n101 ) , .ZN( u2_u12_u0_n130 ) , .A2( u2_u12_u0_n94 ) );
  NAND2_X1 u2_u12_u0_U72 (.ZN( u2_u12_u0_n108 ) , .A1( u2_u12_u0_n92 ) , .A2( u2_u12_u0_n94 ) );
  AND2_X1 u2_u12_u0_U73 (.A1( u2_u12_X_6 ) , .A2( u2_u12_u0_n162 ) , .ZN( u2_u12_u0_n93 ) );
  NOR2_X1 u2_u12_u0_U74 (.A2( u2_u12_X_6 ) , .ZN( u2_u12_u0_n100 ) , .A1( u2_u12_u0_n162 ) );
  NOR2_X1 u2_u12_u0_U75 (.A2( u2_u12_X_3 ) , .A1( u2_u12_X_6 ) , .ZN( u2_u12_u0_n94 ) );
  OAI221_X1 u2_u12_u0_U76 (.C1( u2_u12_u0_n121 ) , .ZN( u2_u12_u0_n122 ) , .B2( u2_u12_u0_n127 ) , .A( u2_u12_u0_n143 ) , .B1( u2_u12_u0_n144 ) , .C2( u2_u12_u0_n147 ) );
  AOI21_X1 u2_u12_u0_U77 (.B1( u2_u12_u0_n132 ) , .ZN( u2_u12_u0_n133 ) , .A( u2_u12_u0_n144 ) , .B2( u2_u12_u0_n166 ) );
  OAI22_X1 u2_u12_u0_U78 (.ZN( u2_u12_u0_n105 ) , .A2( u2_u12_u0_n132 ) , .B1( u2_u12_u0_n146 ) , .A1( u2_u12_u0_n147 ) , .B2( u2_u12_u0_n161 ) );
  NAND2_X1 u2_u12_u0_U79 (.ZN( u2_u12_u0_n110 ) , .A2( u2_u12_u0_n132 ) , .A1( u2_u12_u0_n145 ) );
  AND2_X1 u2_u12_u0_U8 (.A1( u2_u12_u0_n114 ) , .A2( u2_u12_u0_n121 ) , .ZN( u2_u12_u0_n146 ) );
  INV_X1 u2_u12_u0_U80 (.A( u2_u12_u0_n119 ) , .ZN( u2_u12_u0_n167 ) );
  NAND2_X1 u2_u12_u0_U81 (.ZN( u2_u12_u0_n148 ) , .A1( u2_u12_u0_n93 ) , .A2( u2_u12_u0_n95 ) );
  NAND2_X1 u2_u12_u0_U82 (.A1( u2_u12_u0_n100 ) , .ZN( u2_u12_u0_n129 ) , .A2( u2_u12_u0_n95 ) );
  NAND2_X1 u2_u12_u0_U83 (.A1( u2_u12_u0_n102 ) , .ZN( u2_u12_u0_n128 ) , .A2( u2_u12_u0_n95 ) );
  NOR2_X1 u2_u12_u0_U84 (.A2( u2_u12_X_1 ) , .A1( u2_u12_X_2 ) , .ZN( u2_u12_u0_n92 ) );
  NAND2_X1 u2_u12_u0_U85 (.ZN( u2_u12_u0_n142 ) , .A1( u2_u12_u0_n94 ) , .A2( u2_u12_u0_n95 ) );
  NOR2_X1 u2_u12_u0_U86 (.A2( u2_u12_X_2 ) , .ZN( u2_u12_u0_n103 ) , .A1( u2_u12_u0_n164 ) );
  INV_X1 u2_u12_u0_U87 (.A( u2_u12_X_2 ) , .ZN( u2_u12_u0_n163 ) );
  NAND3_X1 u2_u12_u0_U88 (.ZN( u2_out12_23 ) , .A3( u2_u12_u0_n137 ) , .A1( u2_u12_u0_n168 ) , .A2( u2_u12_u0_n171 ) );
  NAND3_X1 u2_u12_u0_U89 (.A3( u2_u12_u0_n127 ) , .A2( u2_u12_u0_n128 ) , .ZN( u2_u12_u0_n135 ) , .A1( u2_u12_u0_n150 ) );
  NAND2_X1 u2_u12_u0_U9 (.ZN( u2_u12_u0_n113 ) , .A1( u2_u12_u0_n139 ) , .A2( u2_u12_u0_n149 ) );
  NAND3_X1 u2_u12_u0_U90 (.ZN( u2_u12_u0_n117 ) , .A3( u2_u12_u0_n132 ) , .A2( u2_u12_u0_n139 ) , .A1( u2_u12_u0_n148 ) );
  NAND3_X1 u2_u12_u0_U91 (.ZN( u2_u12_u0_n109 ) , .A2( u2_u12_u0_n114 ) , .A3( u2_u12_u0_n140 ) , .A1( u2_u12_u0_n149 ) );
  NAND3_X1 u2_u12_u0_U92 (.ZN( u2_out12_9 ) , .A3( u2_u12_u0_n106 ) , .A2( u2_u12_u0_n171 ) , .A1( u2_u12_u0_n174 ) );
  NAND3_X1 u2_u12_u0_U93 (.A2( u2_u12_u0_n128 ) , .A1( u2_u12_u0_n132 ) , .A3( u2_u12_u0_n146 ) , .ZN( u2_u12_u0_n97 ) );
  NOR2_X1 u2_u12_u1_U10 (.A1( u2_u12_u1_n112 ) , .A2( u2_u12_u1_n116 ) , .ZN( u2_u12_u1_n118 ) );
  NAND3_X1 u2_u12_u1_U100 (.ZN( u2_u12_u1_n113 ) , .A1( u2_u12_u1_n120 ) , .A3( u2_u12_u1_n133 ) , .A2( u2_u12_u1_n155 ) );
  OAI21_X1 u2_u12_u1_U11 (.ZN( u2_u12_u1_n101 ) , .B1( u2_u12_u1_n141 ) , .A( u2_u12_u1_n146 ) , .B2( u2_u12_u1_n183 ) );
  AOI21_X1 u2_u12_u1_U12 (.B2( u2_u12_u1_n155 ) , .B1( u2_u12_u1_n156 ) , .ZN( u2_u12_u1_n157 ) , .A( u2_u12_u1_n174 ) );
  NAND2_X1 u2_u12_u1_U13 (.ZN( u2_u12_u1_n140 ) , .A2( u2_u12_u1_n150 ) , .A1( u2_u12_u1_n155 ) );
  NAND2_X1 u2_u12_u1_U14 (.A1( u2_u12_u1_n131 ) , .ZN( u2_u12_u1_n147 ) , .A2( u2_u12_u1_n153 ) );
  INV_X1 u2_u12_u1_U15 (.A( u2_u12_u1_n139 ) , .ZN( u2_u12_u1_n174 ) );
  INV_X1 u2_u12_u1_U16 (.A( u2_u12_u1_n112 ) , .ZN( u2_u12_u1_n171 ) );
  NAND2_X1 u2_u12_u1_U17 (.ZN( u2_u12_u1_n141 ) , .A1( u2_u12_u1_n153 ) , .A2( u2_u12_u1_n156 ) );
  AND2_X1 u2_u12_u1_U18 (.A1( u2_u12_u1_n123 ) , .ZN( u2_u12_u1_n134 ) , .A2( u2_u12_u1_n161 ) );
  NAND2_X1 u2_u12_u1_U19 (.A2( u2_u12_u1_n115 ) , .A1( u2_u12_u1_n116 ) , .ZN( u2_u12_u1_n148 ) );
  NAND2_X1 u2_u12_u1_U20 (.A2( u2_u12_u1_n133 ) , .A1( u2_u12_u1_n135 ) , .ZN( u2_u12_u1_n159 ) );
  NAND2_X1 u2_u12_u1_U21 (.A2( u2_u12_u1_n115 ) , .A1( u2_u12_u1_n120 ) , .ZN( u2_u12_u1_n132 ) );
  INV_X1 u2_u12_u1_U22 (.A( u2_u12_u1_n154 ) , .ZN( u2_u12_u1_n178 ) );
  INV_X1 u2_u12_u1_U23 (.A( u2_u12_u1_n151 ) , .ZN( u2_u12_u1_n183 ) );
  AND2_X1 u2_u12_u1_U24 (.A1( u2_u12_u1_n129 ) , .A2( u2_u12_u1_n133 ) , .ZN( u2_u12_u1_n149 ) );
  INV_X1 u2_u12_u1_U25 (.A( u2_u12_u1_n131 ) , .ZN( u2_u12_u1_n180 ) );
  OR4_X1 u2_u12_u1_U26 (.A4( u2_u12_u1_n106 ) , .A3( u2_u12_u1_n107 ) , .ZN( u2_u12_u1_n108 ) , .A1( u2_u12_u1_n117 ) , .A2( u2_u12_u1_n184 ) );
  AOI21_X1 u2_u12_u1_U27 (.ZN( u2_u12_u1_n106 ) , .A( u2_u12_u1_n112 ) , .B1( u2_u12_u1_n154 ) , .B2( u2_u12_u1_n156 ) );
  AOI21_X1 u2_u12_u1_U28 (.ZN( u2_u12_u1_n107 ) , .B1( u2_u12_u1_n134 ) , .B2( u2_u12_u1_n149 ) , .A( u2_u12_u1_n174 ) );
  INV_X1 u2_u12_u1_U29 (.A( u2_u12_u1_n101 ) , .ZN( u2_u12_u1_n184 ) );
  INV_X1 u2_u12_u1_U3 (.A( u2_u12_u1_n159 ) , .ZN( u2_u12_u1_n182 ) );
  AOI221_X1 u2_u12_u1_U30 (.B1( u2_u12_u1_n140 ) , .ZN( u2_u12_u1_n167 ) , .B2( u2_u12_u1_n172 ) , .C2( u2_u12_u1_n175 ) , .C1( u2_u12_u1_n178 ) , .A( u2_u12_u1_n188 ) );
  INV_X1 u2_u12_u1_U31 (.ZN( u2_u12_u1_n188 ) , .A( u2_u12_u1_n97 ) );
  AOI211_X1 u2_u12_u1_U32 (.A( u2_u12_u1_n118 ) , .C1( u2_u12_u1_n132 ) , .C2( u2_u12_u1_n139 ) , .B( u2_u12_u1_n96 ) , .ZN( u2_u12_u1_n97 ) );
  AOI21_X1 u2_u12_u1_U33 (.B2( u2_u12_u1_n121 ) , .B1( u2_u12_u1_n135 ) , .A( u2_u12_u1_n152 ) , .ZN( u2_u12_u1_n96 ) );
  OAI221_X1 u2_u12_u1_U34 (.A( u2_u12_u1_n119 ) , .C2( u2_u12_u1_n129 ) , .ZN( u2_u12_u1_n138 ) , .B2( u2_u12_u1_n152 ) , .C1( u2_u12_u1_n174 ) , .B1( u2_u12_u1_n187 ) );
  INV_X1 u2_u12_u1_U35 (.A( u2_u12_u1_n148 ) , .ZN( u2_u12_u1_n187 ) );
  AOI211_X1 u2_u12_u1_U36 (.B( u2_u12_u1_n117 ) , .A( u2_u12_u1_n118 ) , .ZN( u2_u12_u1_n119 ) , .C2( u2_u12_u1_n146 ) , .C1( u2_u12_u1_n159 ) );
  NOR2_X1 u2_u12_u1_U37 (.A1( u2_u12_u1_n168 ) , .A2( u2_u12_u1_n176 ) , .ZN( u2_u12_u1_n98 ) );
  AOI211_X1 u2_u12_u1_U38 (.B( u2_u12_u1_n162 ) , .A( u2_u12_u1_n163 ) , .C2( u2_u12_u1_n164 ) , .ZN( u2_u12_u1_n165 ) , .C1( u2_u12_u1_n171 ) );
  AOI21_X1 u2_u12_u1_U39 (.A( u2_u12_u1_n160 ) , .B2( u2_u12_u1_n161 ) , .ZN( u2_u12_u1_n162 ) , .B1( u2_u12_u1_n182 ) );
  AOI221_X1 u2_u12_u1_U4 (.A( u2_u12_u1_n138 ) , .C2( u2_u12_u1_n139 ) , .C1( u2_u12_u1_n140 ) , .B2( u2_u12_u1_n141 ) , .ZN( u2_u12_u1_n142 ) , .B1( u2_u12_u1_n175 ) );
  OR2_X1 u2_u12_u1_U40 (.A2( u2_u12_u1_n157 ) , .A1( u2_u12_u1_n158 ) , .ZN( u2_u12_u1_n163 ) );
  NAND2_X1 u2_u12_u1_U41 (.A1( u2_u12_u1_n128 ) , .ZN( u2_u12_u1_n146 ) , .A2( u2_u12_u1_n160 ) );
  NAND2_X1 u2_u12_u1_U42 (.A2( u2_u12_u1_n112 ) , .ZN( u2_u12_u1_n139 ) , .A1( u2_u12_u1_n152 ) );
  NAND2_X1 u2_u12_u1_U43 (.A1( u2_u12_u1_n105 ) , .ZN( u2_u12_u1_n156 ) , .A2( u2_u12_u1_n99 ) );
  NOR2_X1 u2_u12_u1_U44 (.ZN( u2_u12_u1_n117 ) , .A1( u2_u12_u1_n121 ) , .A2( u2_u12_u1_n160 ) );
  OAI21_X1 u2_u12_u1_U45 (.B2( u2_u12_u1_n123 ) , .ZN( u2_u12_u1_n145 ) , .B1( u2_u12_u1_n160 ) , .A( u2_u12_u1_n185 ) );
  INV_X1 u2_u12_u1_U46 (.A( u2_u12_u1_n122 ) , .ZN( u2_u12_u1_n185 ) );
  AOI21_X1 u2_u12_u1_U47 (.B2( u2_u12_u1_n120 ) , .B1( u2_u12_u1_n121 ) , .ZN( u2_u12_u1_n122 ) , .A( u2_u12_u1_n128 ) );
  AOI21_X1 u2_u12_u1_U48 (.A( u2_u12_u1_n128 ) , .B2( u2_u12_u1_n129 ) , .ZN( u2_u12_u1_n130 ) , .B1( u2_u12_u1_n150 ) );
  NAND2_X1 u2_u12_u1_U49 (.ZN( u2_u12_u1_n112 ) , .A1( u2_u12_u1_n169 ) , .A2( u2_u12_u1_n170 ) );
  AOI211_X1 u2_u12_u1_U5 (.ZN( u2_u12_u1_n124 ) , .A( u2_u12_u1_n138 ) , .C2( u2_u12_u1_n139 ) , .B( u2_u12_u1_n145 ) , .C1( u2_u12_u1_n147 ) );
  NAND2_X1 u2_u12_u1_U50 (.ZN( u2_u12_u1_n129 ) , .A2( u2_u12_u1_n95 ) , .A1( u2_u12_u1_n98 ) );
  NAND2_X1 u2_u12_u1_U51 (.A1( u2_u12_u1_n102 ) , .ZN( u2_u12_u1_n154 ) , .A2( u2_u12_u1_n99 ) );
  NAND2_X1 u2_u12_u1_U52 (.A2( u2_u12_u1_n100 ) , .ZN( u2_u12_u1_n135 ) , .A1( u2_u12_u1_n99 ) );
  AOI21_X1 u2_u12_u1_U53 (.A( u2_u12_u1_n152 ) , .B2( u2_u12_u1_n153 ) , .B1( u2_u12_u1_n154 ) , .ZN( u2_u12_u1_n158 ) );
  INV_X1 u2_u12_u1_U54 (.A( u2_u12_u1_n160 ) , .ZN( u2_u12_u1_n175 ) );
  NAND2_X1 u2_u12_u1_U55 (.A1( u2_u12_u1_n100 ) , .ZN( u2_u12_u1_n116 ) , .A2( u2_u12_u1_n95 ) );
  NAND2_X1 u2_u12_u1_U56 (.A1( u2_u12_u1_n102 ) , .ZN( u2_u12_u1_n131 ) , .A2( u2_u12_u1_n95 ) );
  NAND2_X1 u2_u12_u1_U57 (.A2( u2_u12_u1_n104 ) , .ZN( u2_u12_u1_n121 ) , .A1( u2_u12_u1_n98 ) );
  NAND2_X1 u2_u12_u1_U58 (.A1( u2_u12_u1_n103 ) , .ZN( u2_u12_u1_n153 ) , .A2( u2_u12_u1_n98 ) );
  NAND2_X1 u2_u12_u1_U59 (.A2( u2_u12_u1_n104 ) , .A1( u2_u12_u1_n105 ) , .ZN( u2_u12_u1_n133 ) );
  AOI22_X1 u2_u12_u1_U6 (.B2( u2_u12_u1_n113 ) , .A2( u2_u12_u1_n114 ) , .ZN( u2_u12_u1_n125 ) , .A1( u2_u12_u1_n171 ) , .B1( u2_u12_u1_n173 ) );
  NAND2_X1 u2_u12_u1_U60 (.ZN( u2_u12_u1_n150 ) , .A2( u2_u12_u1_n98 ) , .A1( u2_u12_u1_n99 ) );
  NAND2_X1 u2_u12_u1_U61 (.A1( u2_u12_u1_n105 ) , .ZN( u2_u12_u1_n155 ) , .A2( u2_u12_u1_n95 ) );
  OAI21_X1 u2_u12_u1_U62 (.ZN( u2_u12_u1_n109 ) , .B1( u2_u12_u1_n129 ) , .B2( u2_u12_u1_n160 ) , .A( u2_u12_u1_n167 ) );
  NAND2_X1 u2_u12_u1_U63 (.A2( u2_u12_u1_n100 ) , .A1( u2_u12_u1_n103 ) , .ZN( u2_u12_u1_n120 ) );
  NAND2_X1 u2_u12_u1_U64 (.A1( u2_u12_u1_n102 ) , .A2( u2_u12_u1_n104 ) , .ZN( u2_u12_u1_n115 ) );
  NAND2_X1 u2_u12_u1_U65 (.A2( u2_u12_u1_n100 ) , .A1( u2_u12_u1_n104 ) , .ZN( u2_u12_u1_n151 ) );
  NAND2_X1 u2_u12_u1_U66 (.A2( u2_u12_u1_n103 ) , .A1( u2_u12_u1_n105 ) , .ZN( u2_u12_u1_n161 ) );
  INV_X1 u2_u12_u1_U67 (.A( u2_u12_u1_n152 ) , .ZN( u2_u12_u1_n173 ) );
  INV_X1 u2_u12_u1_U68 (.A( u2_u12_u1_n128 ) , .ZN( u2_u12_u1_n172 ) );
  NAND2_X1 u2_u12_u1_U69 (.A2( u2_u12_u1_n102 ) , .A1( u2_u12_u1_n103 ) , .ZN( u2_u12_u1_n123 ) );
  NAND2_X1 u2_u12_u1_U7 (.ZN( u2_u12_u1_n114 ) , .A1( u2_u12_u1_n134 ) , .A2( u2_u12_u1_n156 ) );
  NOR2_X1 u2_u12_u1_U70 (.A2( u2_u12_X_7 ) , .A1( u2_u12_X_8 ) , .ZN( u2_u12_u1_n95 ) );
  NOR2_X1 u2_u12_u1_U71 (.A1( u2_u12_X_12 ) , .A2( u2_u12_X_9 ) , .ZN( u2_u12_u1_n100 ) );
  NOR2_X1 u2_u12_u1_U72 (.A2( u2_u12_X_8 ) , .A1( u2_u12_u1_n177 ) , .ZN( u2_u12_u1_n99 ) );
  NOR2_X1 u2_u12_u1_U73 (.A2( u2_u12_X_12 ) , .ZN( u2_u12_u1_n102 ) , .A1( u2_u12_u1_n176 ) );
  NOR2_X1 u2_u12_u1_U74 (.A2( u2_u12_X_9 ) , .ZN( u2_u12_u1_n105 ) , .A1( u2_u12_u1_n168 ) );
  NAND2_X1 u2_u12_u1_U75 (.A1( u2_u12_X_10 ) , .ZN( u2_u12_u1_n160 ) , .A2( u2_u12_u1_n169 ) );
  NAND2_X1 u2_u12_u1_U76 (.A2( u2_u12_X_10 ) , .A1( u2_u12_X_11 ) , .ZN( u2_u12_u1_n152 ) );
  NAND2_X1 u2_u12_u1_U77 (.A1( u2_u12_X_11 ) , .ZN( u2_u12_u1_n128 ) , .A2( u2_u12_u1_n170 ) );
  AND2_X1 u2_u12_u1_U78 (.A2( u2_u12_X_7 ) , .A1( u2_u12_X_8 ) , .ZN( u2_u12_u1_n104 ) );
  AND2_X1 u2_u12_u1_U79 (.A1( u2_u12_X_8 ) , .ZN( u2_u12_u1_n103 ) , .A2( u2_u12_u1_n177 ) );
  AOI22_X1 u2_u12_u1_U8 (.B2( u2_u12_u1_n136 ) , .A2( u2_u12_u1_n137 ) , .ZN( u2_u12_u1_n143 ) , .A1( u2_u12_u1_n171 ) , .B1( u2_u12_u1_n173 ) );
  INV_X1 u2_u12_u1_U80 (.A( u2_u12_X_10 ) , .ZN( u2_u12_u1_n170 ) );
  INV_X1 u2_u12_u1_U81 (.A( u2_u12_X_9 ) , .ZN( u2_u12_u1_n176 ) );
  INV_X1 u2_u12_u1_U82 (.A( u2_u12_X_11 ) , .ZN( u2_u12_u1_n169 ) );
  INV_X1 u2_u12_u1_U83 (.A( u2_u12_X_12 ) , .ZN( u2_u12_u1_n168 ) );
  INV_X1 u2_u12_u1_U84 (.A( u2_u12_X_7 ) , .ZN( u2_u12_u1_n177 ) );
  NAND4_X1 u2_u12_u1_U85 (.ZN( u2_out12_28 ) , .A4( u2_u12_u1_n124 ) , .A3( u2_u12_u1_n125 ) , .A2( u2_u12_u1_n126 ) , .A1( u2_u12_u1_n127 ) );
  OAI21_X1 u2_u12_u1_U86 (.ZN( u2_u12_u1_n127 ) , .B2( u2_u12_u1_n139 ) , .B1( u2_u12_u1_n175 ) , .A( u2_u12_u1_n183 ) );
  OAI21_X1 u2_u12_u1_U87 (.ZN( u2_u12_u1_n126 ) , .B2( u2_u12_u1_n140 ) , .A( u2_u12_u1_n146 ) , .B1( u2_u12_u1_n178 ) );
  NAND4_X1 u2_u12_u1_U88 (.ZN( u2_out12_18 ) , .A4( u2_u12_u1_n165 ) , .A3( u2_u12_u1_n166 ) , .A1( u2_u12_u1_n167 ) , .A2( u2_u12_u1_n186 ) );
  AOI22_X1 u2_u12_u1_U89 (.B2( u2_u12_u1_n146 ) , .B1( u2_u12_u1_n147 ) , .A2( u2_u12_u1_n148 ) , .ZN( u2_u12_u1_n166 ) , .A1( u2_u12_u1_n172 ) );
  INV_X1 u2_u12_u1_U9 (.A( u2_u12_u1_n147 ) , .ZN( u2_u12_u1_n181 ) );
  INV_X1 u2_u12_u1_U90 (.A( u2_u12_u1_n145 ) , .ZN( u2_u12_u1_n186 ) );
  NAND4_X1 u2_u12_u1_U91 (.ZN( u2_out12_2 ) , .A4( u2_u12_u1_n142 ) , .A3( u2_u12_u1_n143 ) , .A2( u2_u12_u1_n144 ) , .A1( u2_u12_u1_n179 ) );
  OAI21_X1 u2_u12_u1_U92 (.B2( u2_u12_u1_n132 ) , .ZN( u2_u12_u1_n144 ) , .A( u2_u12_u1_n146 ) , .B1( u2_u12_u1_n180 ) );
  INV_X1 u2_u12_u1_U93 (.A( u2_u12_u1_n130 ) , .ZN( u2_u12_u1_n179 ) );
  OR4_X1 u2_u12_u1_U94 (.ZN( u2_out12_13 ) , .A4( u2_u12_u1_n108 ) , .A3( u2_u12_u1_n109 ) , .A2( u2_u12_u1_n110 ) , .A1( u2_u12_u1_n111 ) );
  AOI21_X1 u2_u12_u1_U95 (.ZN( u2_u12_u1_n111 ) , .A( u2_u12_u1_n128 ) , .B2( u2_u12_u1_n131 ) , .B1( u2_u12_u1_n135 ) );
  AOI21_X1 u2_u12_u1_U96 (.ZN( u2_u12_u1_n110 ) , .A( u2_u12_u1_n116 ) , .B1( u2_u12_u1_n152 ) , .B2( u2_u12_u1_n160 ) );
  NAND3_X1 u2_u12_u1_U97 (.A3( u2_u12_u1_n149 ) , .A2( u2_u12_u1_n150 ) , .A1( u2_u12_u1_n151 ) , .ZN( u2_u12_u1_n164 ) );
  NAND3_X1 u2_u12_u1_U98 (.A3( u2_u12_u1_n134 ) , .A2( u2_u12_u1_n135 ) , .ZN( u2_u12_u1_n136 ) , .A1( u2_u12_u1_n151 ) );
  NAND3_X1 u2_u12_u1_U99 (.A1( u2_u12_u1_n133 ) , .ZN( u2_u12_u1_n137 ) , .A2( u2_u12_u1_n154 ) , .A3( u2_u12_u1_n181 ) );
  OAI22_X1 u2_u12_u4_U10 (.B2( u2_u12_u4_n135 ) , .ZN( u2_u12_u4_n137 ) , .B1( u2_u12_u4_n153 ) , .A1( u2_u12_u4_n155 ) , .A2( u2_u12_u4_n171 ) );
  AND3_X1 u2_u12_u4_U11 (.A2( u2_u12_u4_n134 ) , .ZN( u2_u12_u4_n135 ) , .A3( u2_u12_u4_n145 ) , .A1( u2_u12_u4_n157 ) );
  NAND2_X1 u2_u12_u4_U12 (.ZN( u2_u12_u4_n132 ) , .A2( u2_u12_u4_n170 ) , .A1( u2_u12_u4_n173 ) );
  AOI21_X1 u2_u12_u4_U13 (.B2( u2_u12_u4_n160 ) , .B1( u2_u12_u4_n161 ) , .ZN( u2_u12_u4_n162 ) , .A( u2_u12_u4_n170 ) );
  AOI21_X1 u2_u12_u4_U14 (.ZN( u2_u12_u4_n107 ) , .B2( u2_u12_u4_n143 ) , .A( u2_u12_u4_n174 ) , .B1( u2_u12_u4_n184 ) );
  AOI21_X1 u2_u12_u4_U15 (.B2( u2_u12_u4_n158 ) , .B1( u2_u12_u4_n159 ) , .ZN( u2_u12_u4_n163 ) , .A( u2_u12_u4_n174 ) );
  AOI21_X1 u2_u12_u4_U16 (.A( u2_u12_u4_n153 ) , .B2( u2_u12_u4_n154 ) , .B1( u2_u12_u4_n155 ) , .ZN( u2_u12_u4_n165 ) );
  AOI21_X1 u2_u12_u4_U17 (.A( u2_u12_u4_n156 ) , .B2( u2_u12_u4_n157 ) , .ZN( u2_u12_u4_n164 ) , .B1( u2_u12_u4_n184 ) );
  INV_X1 u2_u12_u4_U18 (.A( u2_u12_u4_n138 ) , .ZN( u2_u12_u4_n170 ) );
  AND2_X1 u2_u12_u4_U19 (.A2( u2_u12_u4_n120 ) , .ZN( u2_u12_u4_n155 ) , .A1( u2_u12_u4_n160 ) );
  INV_X1 u2_u12_u4_U20 (.A( u2_u12_u4_n156 ) , .ZN( u2_u12_u4_n175 ) );
  NAND2_X1 u2_u12_u4_U21 (.A2( u2_u12_u4_n118 ) , .ZN( u2_u12_u4_n131 ) , .A1( u2_u12_u4_n147 ) );
  NAND2_X1 u2_u12_u4_U22 (.A1( u2_u12_u4_n119 ) , .A2( u2_u12_u4_n120 ) , .ZN( u2_u12_u4_n130 ) );
  NAND2_X1 u2_u12_u4_U23 (.ZN( u2_u12_u4_n117 ) , .A2( u2_u12_u4_n118 ) , .A1( u2_u12_u4_n148 ) );
  NAND2_X1 u2_u12_u4_U24 (.ZN( u2_u12_u4_n129 ) , .A1( u2_u12_u4_n134 ) , .A2( u2_u12_u4_n148 ) );
  AND3_X1 u2_u12_u4_U25 (.A1( u2_u12_u4_n119 ) , .A2( u2_u12_u4_n143 ) , .A3( u2_u12_u4_n154 ) , .ZN( u2_u12_u4_n161 ) );
  AND2_X1 u2_u12_u4_U26 (.A1( u2_u12_u4_n145 ) , .A2( u2_u12_u4_n147 ) , .ZN( u2_u12_u4_n159 ) );
  OR3_X1 u2_u12_u4_U27 (.A3( u2_u12_u4_n114 ) , .A2( u2_u12_u4_n115 ) , .A1( u2_u12_u4_n116 ) , .ZN( u2_u12_u4_n136 ) );
  AOI21_X1 u2_u12_u4_U28 (.A( u2_u12_u4_n113 ) , .ZN( u2_u12_u4_n116 ) , .B2( u2_u12_u4_n173 ) , .B1( u2_u12_u4_n174 ) );
  AOI21_X1 u2_u12_u4_U29 (.ZN( u2_u12_u4_n115 ) , .B2( u2_u12_u4_n145 ) , .B1( u2_u12_u4_n146 ) , .A( u2_u12_u4_n156 ) );
  NOR2_X1 u2_u12_u4_U3 (.ZN( u2_u12_u4_n121 ) , .A1( u2_u12_u4_n181 ) , .A2( u2_u12_u4_n182 ) );
  OAI22_X1 u2_u12_u4_U30 (.ZN( u2_u12_u4_n114 ) , .A2( u2_u12_u4_n121 ) , .B1( u2_u12_u4_n160 ) , .B2( u2_u12_u4_n170 ) , .A1( u2_u12_u4_n171 ) );
  INV_X1 u2_u12_u4_U31 (.A( u2_u12_u4_n158 ) , .ZN( u2_u12_u4_n182 ) );
  INV_X1 u2_u12_u4_U32 (.ZN( u2_u12_u4_n181 ) , .A( u2_u12_u4_n96 ) );
  INV_X1 u2_u12_u4_U33 (.A( u2_u12_u4_n144 ) , .ZN( u2_u12_u4_n179 ) );
  INV_X1 u2_u12_u4_U34 (.A( u2_u12_u4_n157 ) , .ZN( u2_u12_u4_n178 ) );
  NAND2_X1 u2_u12_u4_U35 (.A2( u2_u12_u4_n154 ) , .A1( u2_u12_u4_n96 ) , .ZN( u2_u12_u4_n97 ) );
  INV_X1 u2_u12_u4_U36 (.ZN( u2_u12_u4_n186 ) , .A( u2_u12_u4_n95 ) );
  OAI221_X1 u2_u12_u4_U37 (.C1( u2_u12_u4_n134 ) , .B1( u2_u12_u4_n158 ) , .B2( u2_u12_u4_n171 ) , .C2( u2_u12_u4_n173 ) , .A( u2_u12_u4_n94 ) , .ZN( u2_u12_u4_n95 ) );
  AOI222_X1 u2_u12_u4_U38 (.B2( u2_u12_u4_n132 ) , .A1( u2_u12_u4_n138 ) , .C2( u2_u12_u4_n175 ) , .A2( u2_u12_u4_n179 ) , .C1( u2_u12_u4_n181 ) , .B1( u2_u12_u4_n185 ) , .ZN( u2_u12_u4_n94 ) );
  INV_X1 u2_u12_u4_U39 (.A( u2_u12_u4_n113 ) , .ZN( u2_u12_u4_n185 ) );
  INV_X1 u2_u12_u4_U4 (.A( u2_u12_u4_n117 ) , .ZN( u2_u12_u4_n184 ) );
  INV_X1 u2_u12_u4_U40 (.A( u2_u12_u4_n143 ) , .ZN( u2_u12_u4_n183 ) );
  NOR2_X1 u2_u12_u4_U41 (.ZN( u2_u12_u4_n138 ) , .A1( u2_u12_u4_n168 ) , .A2( u2_u12_u4_n169 ) );
  NOR2_X1 u2_u12_u4_U42 (.A1( u2_u12_u4_n150 ) , .A2( u2_u12_u4_n152 ) , .ZN( u2_u12_u4_n153 ) );
  NOR2_X1 u2_u12_u4_U43 (.A2( u2_u12_u4_n128 ) , .A1( u2_u12_u4_n138 ) , .ZN( u2_u12_u4_n156 ) );
  AOI22_X1 u2_u12_u4_U44 (.B2( u2_u12_u4_n122 ) , .A1( u2_u12_u4_n123 ) , .ZN( u2_u12_u4_n124 ) , .B1( u2_u12_u4_n128 ) , .A2( u2_u12_u4_n172 ) );
  INV_X1 u2_u12_u4_U45 (.A( u2_u12_u4_n153 ) , .ZN( u2_u12_u4_n172 ) );
  NAND2_X1 u2_u12_u4_U46 (.A2( u2_u12_u4_n120 ) , .ZN( u2_u12_u4_n123 ) , .A1( u2_u12_u4_n161 ) );
  AOI22_X1 u2_u12_u4_U47 (.B2( u2_u12_u4_n132 ) , .A2( u2_u12_u4_n133 ) , .ZN( u2_u12_u4_n140 ) , .A1( u2_u12_u4_n150 ) , .B1( u2_u12_u4_n179 ) );
  NAND2_X1 u2_u12_u4_U48 (.ZN( u2_u12_u4_n133 ) , .A2( u2_u12_u4_n146 ) , .A1( u2_u12_u4_n154 ) );
  NAND2_X1 u2_u12_u4_U49 (.A1( u2_u12_u4_n103 ) , .ZN( u2_u12_u4_n154 ) , .A2( u2_u12_u4_n98 ) );
  NOR4_X1 u2_u12_u4_U5 (.A4( u2_u12_u4_n106 ) , .A3( u2_u12_u4_n107 ) , .A2( u2_u12_u4_n108 ) , .A1( u2_u12_u4_n109 ) , .ZN( u2_u12_u4_n110 ) );
  NAND2_X1 u2_u12_u4_U50 (.A1( u2_u12_u4_n101 ) , .ZN( u2_u12_u4_n158 ) , .A2( u2_u12_u4_n99 ) );
  AOI21_X1 u2_u12_u4_U51 (.ZN( u2_u12_u4_n127 ) , .A( u2_u12_u4_n136 ) , .B2( u2_u12_u4_n150 ) , .B1( u2_u12_u4_n180 ) );
  INV_X1 u2_u12_u4_U52 (.A( u2_u12_u4_n160 ) , .ZN( u2_u12_u4_n180 ) );
  NAND2_X1 u2_u12_u4_U53 (.A2( u2_u12_u4_n104 ) , .A1( u2_u12_u4_n105 ) , .ZN( u2_u12_u4_n146 ) );
  NAND2_X1 u2_u12_u4_U54 (.A2( u2_u12_u4_n101 ) , .A1( u2_u12_u4_n102 ) , .ZN( u2_u12_u4_n160 ) );
  NAND2_X1 u2_u12_u4_U55 (.ZN( u2_u12_u4_n134 ) , .A1( u2_u12_u4_n98 ) , .A2( u2_u12_u4_n99 ) );
  NAND2_X1 u2_u12_u4_U56 (.A1( u2_u12_u4_n103 ) , .A2( u2_u12_u4_n104 ) , .ZN( u2_u12_u4_n143 ) );
  NAND2_X1 u2_u12_u4_U57 (.A2( u2_u12_u4_n105 ) , .ZN( u2_u12_u4_n145 ) , .A1( u2_u12_u4_n98 ) );
  NAND2_X1 u2_u12_u4_U58 (.A1( u2_u12_u4_n100 ) , .A2( u2_u12_u4_n105 ) , .ZN( u2_u12_u4_n120 ) );
  NAND2_X1 u2_u12_u4_U59 (.A1( u2_u12_u4_n102 ) , .A2( u2_u12_u4_n104 ) , .ZN( u2_u12_u4_n148 ) );
  AOI21_X1 u2_u12_u4_U6 (.ZN( u2_u12_u4_n106 ) , .B2( u2_u12_u4_n146 ) , .B1( u2_u12_u4_n158 ) , .A( u2_u12_u4_n170 ) );
  NAND2_X1 u2_u12_u4_U60 (.A2( u2_u12_u4_n100 ) , .A1( u2_u12_u4_n103 ) , .ZN( u2_u12_u4_n157 ) );
  INV_X1 u2_u12_u4_U61 (.A( u2_u12_u4_n150 ) , .ZN( u2_u12_u4_n173 ) );
  INV_X1 u2_u12_u4_U62 (.A( u2_u12_u4_n152 ) , .ZN( u2_u12_u4_n171 ) );
  NAND2_X1 u2_u12_u4_U63 (.A1( u2_u12_u4_n100 ) , .ZN( u2_u12_u4_n118 ) , .A2( u2_u12_u4_n99 ) );
  NAND2_X1 u2_u12_u4_U64 (.A2( u2_u12_u4_n100 ) , .A1( u2_u12_u4_n102 ) , .ZN( u2_u12_u4_n144 ) );
  NAND2_X1 u2_u12_u4_U65 (.A2( u2_u12_u4_n101 ) , .A1( u2_u12_u4_n105 ) , .ZN( u2_u12_u4_n96 ) );
  INV_X1 u2_u12_u4_U66 (.A( u2_u12_u4_n128 ) , .ZN( u2_u12_u4_n174 ) );
  NAND2_X1 u2_u12_u4_U67 (.A2( u2_u12_u4_n102 ) , .ZN( u2_u12_u4_n119 ) , .A1( u2_u12_u4_n98 ) );
  NAND2_X1 u2_u12_u4_U68 (.A2( u2_u12_u4_n101 ) , .A1( u2_u12_u4_n103 ) , .ZN( u2_u12_u4_n147 ) );
  NAND2_X1 u2_u12_u4_U69 (.A2( u2_u12_u4_n104 ) , .ZN( u2_u12_u4_n113 ) , .A1( u2_u12_u4_n99 ) );
  AOI21_X1 u2_u12_u4_U7 (.ZN( u2_u12_u4_n108 ) , .B2( u2_u12_u4_n134 ) , .B1( u2_u12_u4_n155 ) , .A( u2_u12_u4_n156 ) );
  NOR2_X1 u2_u12_u4_U70 (.A2( u2_u12_X_28 ) , .ZN( u2_u12_u4_n150 ) , .A1( u2_u12_u4_n168 ) );
  NOR2_X1 u2_u12_u4_U71 (.A2( u2_u12_X_29 ) , .ZN( u2_u12_u4_n152 ) , .A1( u2_u12_u4_n169 ) );
  NOR2_X1 u2_u12_u4_U72 (.A2( u2_u12_X_30 ) , .ZN( u2_u12_u4_n105 ) , .A1( u2_u12_u4_n176 ) );
  NOR2_X1 u2_u12_u4_U73 (.A2( u2_u12_X_26 ) , .ZN( u2_u12_u4_n100 ) , .A1( u2_u12_u4_n177 ) );
  NOR2_X1 u2_u12_u4_U74 (.A2( u2_u12_X_28 ) , .A1( u2_u12_X_29 ) , .ZN( u2_u12_u4_n128 ) );
  NOR2_X1 u2_u12_u4_U75 (.A2( u2_u12_X_27 ) , .A1( u2_u12_X_30 ) , .ZN( u2_u12_u4_n102 ) );
  NOR2_X1 u2_u12_u4_U76 (.A2( u2_u12_X_25 ) , .A1( u2_u12_X_26 ) , .ZN( u2_u12_u4_n98 ) );
  AND2_X1 u2_u12_u4_U77 (.A2( u2_u12_X_25 ) , .A1( u2_u12_X_26 ) , .ZN( u2_u12_u4_n104 ) );
  AND2_X1 u2_u12_u4_U78 (.A1( u2_u12_X_30 ) , .A2( u2_u12_u4_n176 ) , .ZN( u2_u12_u4_n99 ) );
  AND2_X1 u2_u12_u4_U79 (.A1( u2_u12_X_26 ) , .ZN( u2_u12_u4_n101 ) , .A2( u2_u12_u4_n177 ) );
  AOI21_X1 u2_u12_u4_U8 (.ZN( u2_u12_u4_n109 ) , .A( u2_u12_u4_n153 ) , .B1( u2_u12_u4_n159 ) , .B2( u2_u12_u4_n184 ) );
  AND2_X1 u2_u12_u4_U80 (.A1( u2_u12_X_27 ) , .A2( u2_u12_X_30 ) , .ZN( u2_u12_u4_n103 ) );
  INV_X1 u2_u12_u4_U81 (.A( u2_u12_X_28 ) , .ZN( u2_u12_u4_n169 ) );
  INV_X1 u2_u12_u4_U82 (.A( u2_u12_X_29 ) , .ZN( u2_u12_u4_n168 ) );
  INV_X1 u2_u12_u4_U83 (.A( u2_u12_X_25 ) , .ZN( u2_u12_u4_n177 ) );
  INV_X1 u2_u12_u4_U84 (.A( u2_u12_X_27 ) , .ZN( u2_u12_u4_n176 ) );
  NAND4_X1 u2_u12_u4_U85 (.ZN( u2_out12_25 ) , .A4( u2_u12_u4_n139 ) , .A3( u2_u12_u4_n140 ) , .A2( u2_u12_u4_n141 ) , .A1( u2_u12_u4_n142 ) );
  OAI21_X1 u2_u12_u4_U86 (.A( u2_u12_u4_n128 ) , .B2( u2_u12_u4_n129 ) , .B1( u2_u12_u4_n130 ) , .ZN( u2_u12_u4_n142 ) );
  OAI21_X1 u2_u12_u4_U87 (.B2( u2_u12_u4_n131 ) , .ZN( u2_u12_u4_n141 ) , .A( u2_u12_u4_n175 ) , .B1( u2_u12_u4_n183 ) );
  NAND4_X1 u2_u12_u4_U88 (.ZN( u2_out12_14 ) , .A4( u2_u12_u4_n124 ) , .A3( u2_u12_u4_n125 ) , .A2( u2_u12_u4_n126 ) , .A1( u2_u12_u4_n127 ) );
  AOI22_X1 u2_u12_u4_U89 (.B2( u2_u12_u4_n117 ) , .ZN( u2_u12_u4_n126 ) , .A1( u2_u12_u4_n129 ) , .B1( u2_u12_u4_n152 ) , .A2( u2_u12_u4_n175 ) );
  AOI211_X1 u2_u12_u4_U9 (.B( u2_u12_u4_n136 ) , .A( u2_u12_u4_n137 ) , .C2( u2_u12_u4_n138 ) , .ZN( u2_u12_u4_n139 ) , .C1( u2_u12_u4_n182 ) );
  AOI22_X1 u2_u12_u4_U90 (.ZN( u2_u12_u4_n125 ) , .B2( u2_u12_u4_n131 ) , .A2( u2_u12_u4_n132 ) , .B1( u2_u12_u4_n138 ) , .A1( u2_u12_u4_n178 ) );
  NAND4_X1 u2_u12_u4_U91 (.ZN( u2_out12_8 ) , .A4( u2_u12_u4_n110 ) , .A3( u2_u12_u4_n111 ) , .A2( u2_u12_u4_n112 ) , .A1( u2_u12_u4_n186 ) );
  NAND2_X1 u2_u12_u4_U92 (.ZN( u2_u12_u4_n112 ) , .A2( u2_u12_u4_n130 ) , .A1( u2_u12_u4_n150 ) );
  AOI22_X1 u2_u12_u4_U93 (.ZN( u2_u12_u4_n111 ) , .B2( u2_u12_u4_n132 ) , .A1( u2_u12_u4_n152 ) , .B1( u2_u12_u4_n178 ) , .A2( u2_u12_u4_n97 ) );
  AOI22_X1 u2_u12_u4_U94 (.B2( u2_u12_u4_n149 ) , .B1( u2_u12_u4_n150 ) , .A2( u2_u12_u4_n151 ) , .A1( u2_u12_u4_n152 ) , .ZN( u2_u12_u4_n167 ) );
  NOR4_X1 u2_u12_u4_U95 (.A4( u2_u12_u4_n162 ) , .A3( u2_u12_u4_n163 ) , .A2( u2_u12_u4_n164 ) , .A1( u2_u12_u4_n165 ) , .ZN( u2_u12_u4_n166 ) );
  NAND3_X1 u2_u12_u4_U96 (.ZN( u2_out12_3 ) , .A3( u2_u12_u4_n166 ) , .A1( u2_u12_u4_n167 ) , .A2( u2_u12_u4_n186 ) );
  NAND3_X1 u2_u12_u4_U97 (.A3( u2_u12_u4_n146 ) , .A2( u2_u12_u4_n147 ) , .A1( u2_u12_u4_n148 ) , .ZN( u2_u12_u4_n149 ) );
  NAND3_X1 u2_u12_u4_U98 (.A3( u2_u12_u4_n143 ) , .A2( u2_u12_u4_n144 ) , .A1( u2_u12_u4_n145 ) , .ZN( u2_u12_u4_n151 ) );
  NAND3_X1 u2_u12_u4_U99 (.A3( u2_u12_u4_n121 ) , .ZN( u2_u12_u4_n122 ) , .A2( u2_u12_u4_n144 ) , .A1( u2_u12_u4_n154 ) );
  INV_X1 u2_u12_u5_U10 (.A( u2_u12_u5_n121 ) , .ZN( u2_u12_u5_n177 ) );
  NOR3_X1 u2_u12_u5_U100 (.A3( u2_u12_u5_n141 ) , .A1( u2_u12_u5_n142 ) , .ZN( u2_u12_u5_n143 ) , .A2( u2_u12_u5_n191 ) );
  NAND4_X1 u2_u12_u5_U101 (.ZN( u2_out12_4 ) , .A4( u2_u12_u5_n112 ) , .A2( u2_u12_u5_n113 ) , .A1( u2_u12_u5_n114 ) , .A3( u2_u12_u5_n195 ) );
  AOI211_X1 u2_u12_u5_U102 (.A( u2_u12_u5_n110 ) , .C1( u2_u12_u5_n111 ) , .ZN( u2_u12_u5_n112 ) , .B( u2_u12_u5_n118 ) , .C2( u2_u12_u5_n177 ) );
  AOI222_X1 u2_u12_u5_U103 (.ZN( u2_u12_u5_n113 ) , .A1( u2_u12_u5_n131 ) , .C1( u2_u12_u5_n148 ) , .B2( u2_u12_u5_n174 ) , .C2( u2_u12_u5_n178 ) , .A2( u2_u12_u5_n179 ) , .B1( u2_u12_u5_n99 ) );
  NAND3_X1 u2_u12_u5_U104 (.A2( u2_u12_u5_n154 ) , .A3( u2_u12_u5_n158 ) , .A1( u2_u12_u5_n161 ) , .ZN( u2_u12_u5_n99 ) );
  NOR2_X1 u2_u12_u5_U11 (.ZN( u2_u12_u5_n160 ) , .A2( u2_u12_u5_n173 ) , .A1( u2_u12_u5_n177 ) );
  INV_X1 u2_u12_u5_U12 (.A( u2_u12_u5_n150 ) , .ZN( u2_u12_u5_n174 ) );
  AOI21_X1 u2_u12_u5_U13 (.A( u2_u12_u5_n160 ) , .B2( u2_u12_u5_n161 ) , .ZN( u2_u12_u5_n162 ) , .B1( u2_u12_u5_n192 ) );
  INV_X1 u2_u12_u5_U14 (.A( u2_u12_u5_n159 ) , .ZN( u2_u12_u5_n192 ) );
  AOI21_X1 u2_u12_u5_U15 (.A( u2_u12_u5_n156 ) , .B2( u2_u12_u5_n157 ) , .B1( u2_u12_u5_n158 ) , .ZN( u2_u12_u5_n163 ) );
  AOI21_X1 u2_u12_u5_U16 (.B2( u2_u12_u5_n139 ) , .B1( u2_u12_u5_n140 ) , .ZN( u2_u12_u5_n141 ) , .A( u2_u12_u5_n150 ) );
  OAI21_X1 u2_u12_u5_U17 (.A( u2_u12_u5_n133 ) , .B2( u2_u12_u5_n134 ) , .B1( u2_u12_u5_n135 ) , .ZN( u2_u12_u5_n142 ) );
  OAI21_X1 u2_u12_u5_U18 (.ZN( u2_u12_u5_n133 ) , .B2( u2_u12_u5_n147 ) , .A( u2_u12_u5_n173 ) , .B1( u2_u12_u5_n188 ) );
  NAND2_X1 u2_u12_u5_U19 (.A2( u2_u12_u5_n119 ) , .A1( u2_u12_u5_n123 ) , .ZN( u2_u12_u5_n137 ) );
  INV_X1 u2_u12_u5_U20 (.A( u2_u12_u5_n155 ) , .ZN( u2_u12_u5_n194 ) );
  NAND2_X1 u2_u12_u5_U21 (.A1( u2_u12_u5_n121 ) , .ZN( u2_u12_u5_n132 ) , .A2( u2_u12_u5_n172 ) );
  NAND2_X1 u2_u12_u5_U22 (.A2( u2_u12_u5_n122 ) , .ZN( u2_u12_u5_n136 ) , .A1( u2_u12_u5_n154 ) );
  NAND2_X1 u2_u12_u5_U23 (.A2( u2_u12_u5_n119 ) , .A1( u2_u12_u5_n120 ) , .ZN( u2_u12_u5_n159 ) );
  INV_X1 u2_u12_u5_U24 (.A( u2_u12_u5_n156 ) , .ZN( u2_u12_u5_n175 ) );
  INV_X1 u2_u12_u5_U25 (.A( u2_u12_u5_n158 ) , .ZN( u2_u12_u5_n188 ) );
  INV_X1 u2_u12_u5_U26 (.A( u2_u12_u5_n152 ) , .ZN( u2_u12_u5_n179 ) );
  INV_X1 u2_u12_u5_U27 (.A( u2_u12_u5_n140 ) , .ZN( u2_u12_u5_n182 ) );
  INV_X1 u2_u12_u5_U28 (.A( u2_u12_u5_n151 ) , .ZN( u2_u12_u5_n183 ) );
  INV_X1 u2_u12_u5_U29 (.A( u2_u12_u5_n123 ) , .ZN( u2_u12_u5_n185 ) );
  NOR2_X1 u2_u12_u5_U3 (.ZN( u2_u12_u5_n134 ) , .A1( u2_u12_u5_n183 ) , .A2( u2_u12_u5_n190 ) );
  INV_X1 u2_u12_u5_U30 (.A( u2_u12_u5_n161 ) , .ZN( u2_u12_u5_n184 ) );
  INV_X1 u2_u12_u5_U31 (.A( u2_u12_u5_n139 ) , .ZN( u2_u12_u5_n189 ) );
  INV_X1 u2_u12_u5_U32 (.A( u2_u12_u5_n157 ) , .ZN( u2_u12_u5_n190 ) );
  INV_X1 u2_u12_u5_U33 (.A( u2_u12_u5_n120 ) , .ZN( u2_u12_u5_n193 ) );
  NAND2_X1 u2_u12_u5_U34 (.ZN( u2_u12_u5_n111 ) , .A1( u2_u12_u5_n140 ) , .A2( u2_u12_u5_n155 ) );
  NOR2_X1 u2_u12_u5_U35 (.ZN( u2_u12_u5_n100 ) , .A1( u2_u12_u5_n170 ) , .A2( u2_u12_u5_n180 ) );
  INV_X1 u2_u12_u5_U36 (.A( u2_u12_u5_n117 ) , .ZN( u2_u12_u5_n196 ) );
  OAI221_X1 u2_u12_u5_U37 (.A( u2_u12_u5_n116 ) , .ZN( u2_u12_u5_n117 ) , .B2( u2_u12_u5_n119 ) , .C1( u2_u12_u5_n153 ) , .C2( u2_u12_u5_n158 ) , .B1( u2_u12_u5_n172 ) );
  AOI222_X1 u2_u12_u5_U38 (.ZN( u2_u12_u5_n116 ) , .B2( u2_u12_u5_n145 ) , .C1( u2_u12_u5_n148 ) , .A2( u2_u12_u5_n174 ) , .C2( u2_u12_u5_n177 ) , .B1( u2_u12_u5_n187 ) , .A1( u2_u12_u5_n193 ) );
  INV_X1 u2_u12_u5_U39 (.A( u2_u12_u5_n115 ) , .ZN( u2_u12_u5_n187 ) );
  INV_X1 u2_u12_u5_U4 (.A( u2_u12_u5_n138 ) , .ZN( u2_u12_u5_n191 ) );
  AOI22_X1 u2_u12_u5_U40 (.B2( u2_u12_u5_n131 ) , .A2( u2_u12_u5_n146 ) , .ZN( u2_u12_u5_n169 ) , .B1( u2_u12_u5_n174 ) , .A1( u2_u12_u5_n185 ) );
  NOR2_X1 u2_u12_u5_U41 (.A1( u2_u12_u5_n146 ) , .ZN( u2_u12_u5_n150 ) , .A2( u2_u12_u5_n173 ) );
  AOI21_X1 u2_u12_u5_U42 (.A( u2_u12_u5_n118 ) , .B2( u2_u12_u5_n145 ) , .ZN( u2_u12_u5_n168 ) , .B1( u2_u12_u5_n186 ) );
  INV_X1 u2_u12_u5_U43 (.A( u2_u12_u5_n122 ) , .ZN( u2_u12_u5_n186 ) );
  NOR2_X1 u2_u12_u5_U44 (.A1( u2_u12_u5_n146 ) , .ZN( u2_u12_u5_n152 ) , .A2( u2_u12_u5_n176 ) );
  NOR2_X1 u2_u12_u5_U45 (.A1( u2_u12_u5_n115 ) , .ZN( u2_u12_u5_n118 ) , .A2( u2_u12_u5_n153 ) );
  NOR2_X1 u2_u12_u5_U46 (.A2( u2_u12_u5_n145 ) , .ZN( u2_u12_u5_n156 ) , .A1( u2_u12_u5_n174 ) );
  NOR2_X1 u2_u12_u5_U47 (.ZN( u2_u12_u5_n121 ) , .A2( u2_u12_u5_n145 ) , .A1( u2_u12_u5_n176 ) );
  AOI22_X1 u2_u12_u5_U48 (.ZN( u2_u12_u5_n114 ) , .A2( u2_u12_u5_n137 ) , .A1( u2_u12_u5_n145 ) , .B2( u2_u12_u5_n175 ) , .B1( u2_u12_u5_n193 ) );
  OAI211_X1 u2_u12_u5_U49 (.B( u2_u12_u5_n124 ) , .A( u2_u12_u5_n125 ) , .C2( u2_u12_u5_n126 ) , .C1( u2_u12_u5_n127 ) , .ZN( u2_u12_u5_n128 ) );
  OAI21_X1 u2_u12_u5_U5 (.B2( u2_u12_u5_n136 ) , .B1( u2_u12_u5_n137 ) , .ZN( u2_u12_u5_n138 ) , .A( u2_u12_u5_n177 ) );
  NOR3_X1 u2_u12_u5_U50 (.ZN( u2_u12_u5_n127 ) , .A1( u2_u12_u5_n136 ) , .A3( u2_u12_u5_n148 ) , .A2( u2_u12_u5_n182 ) );
  OAI21_X1 u2_u12_u5_U51 (.ZN( u2_u12_u5_n124 ) , .A( u2_u12_u5_n177 ) , .B2( u2_u12_u5_n183 ) , .B1( u2_u12_u5_n189 ) );
  OAI21_X1 u2_u12_u5_U52 (.ZN( u2_u12_u5_n125 ) , .A( u2_u12_u5_n174 ) , .B2( u2_u12_u5_n185 ) , .B1( u2_u12_u5_n190 ) );
  AOI21_X1 u2_u12_u5_U53 (.A( u2_u12_u5_n153 ) , .B2( u2_u12_u5_n154 ) , .B1( u2_u12_u5_n155 ) , .ZN( u2_u12_u5_n164 ) );
  AOI21_X1 u2_u12_u5_U54 (.ZN( u2_u12_u5_n110 ) , .B1( u2_u12_u5_n122 ) , .B2( u2_u12_u5_n139 ) , .A( u2_u12_u5_n153 ) );
  INV_X1 u2_u12_u5_U55 (.A( u2_u12_u5_n153 ) , .ZN( u2_u12_u5_n176 ) );
  INV_X1 u2_u12_u5_U56 (.A( u2_u12_u5_n126 ) , .ZN( u2_u12_u5_n173 ) );
  AND2_X1 u2_u12_u5_U57 (.A2( u2_u12_u5_n104 ) , .A1( u2_u12_u5_n107 ) , .ZN( u2_u12_u5_n147 ) );
  AND2_X1 u2_u12_u5_U58 (.A2( u2_u12_u5_n104 ) , .A1( u2_u12_u5_n108 ) , .ZN( u2_u12_u5_n148 ) );
  NAND2_X1 u2_u12_u5_U59 (.A1( u2_u12_u5_n105 ) , .A2( u2_u12_u5_n106 ) , .ZN( u2_u12_u5_n158 ) );
  INV_X1 u2_u12_u5_U6 (.A( u2_u12_u5_n135 ) , .ZN( u2_u12_u5_n178 ) );
  NAND2_X1 u2_u12_u5_U60 (.A2( u2_u12_u5_n108 ) , .A1( u2_u12_u5_n109 ) , .ZN( u2_u12_u5_n139 ) );
  NAND2_X1 u2_u12_u5_U61 (.A1( u2_u12_u5_n106 ) , .A2( u2_u12_u5_n108 ) , .ZN( u2_u12_u5_n119 ) );
  NAND2_X1 u2_u12_u5_U62 (.A2( u2_u12_u5_n103 ) , .A1( u2_u12_u5_n105 ) , .ZN( u2_u12_u5_n140 ) );
  NAND2_X1 u2_u12_u5_U63 (.A2( u2_u12_u5_n104 ) , .A1( u2_u12_u5_n105 ) , .ZN( u2_u12_u5_n155 ) );
  NAND2_X1 u2_u12_u5_U64 (.A2( u2_u12_u5_n106 ) , .A1( u2_u12_u5_n107 ) , .ZN( u2_u12_u5_n122 ) );
  NAND2_X1 u2_u12_u5_U65 (.A2( u2_u12_u5_n100 ) , .A1( u2_u12_u5_n106 ) , .ZN( u2_u12_u5_n115 ) );
  NAND2_X1 u2_u12_u5_U66 (.A2( u2_u12_u5_n100 ) , .A1( u2_u12_u5_n103 ) , .ZN( u2_u12_u5_n161 ) );
  NAND2_X1 u2_u12_u5_U67 (.A1( u2_u12_u5_n105 ) , .A2( u2_u12_u5_n109 ) , .ZN( u2_u12_u5_n154 ) );
  INV_X1 u2_u12_u5_U68 (.A( u2_u12_u5_n146 ) , .ZN( u2_u12_u5_n172 ) );
  NAND2_X1 u2_u12_u5_U69 (.A1( u2_u12_u5_n103 ) , .A2( u2_u12_u5_n108 ) , .ZN( u2_u12_u5_n123 ) );
  OAI22_X1 u2_u12_u5_U7 (.B2( u2_u12_u5_n149 ) , .B1( u2_u12_u5_n150 ) , .A2( u2_u12_u5_n151 ) , .A1( u2_u12_u5_n152 ) , .ZN( u2_u12_u5_n165 ) );
  NAND2_X1 u2_u12_u5_U70 (.A2( u2_u12_u5_n103 ) , .A1( u2_u12_u5_n107 ) , .ZN( u2_u12_u5_n151 ) );
  NAND2_X1 u2_u12_u5_U71 (.A2( u2_u12_u5_n107 ) , .A1( u2_u12_u5_n109 ) , .ZN( u2_u12_u5_n120 ) );
  NAND2_X1 u2_u12_u5_U72 (.A2( u2_u12_u5_n100 ) , .A1( u2_u12_u5_n109 ) , .ZN( u2_u12_u5_n157 ) );
  AND2_X1 u2_u12_u5_U73 (.A2( u2_u12_u5_n100 ) , .A1( u2_u12_u5_n104 ) , .ZN( u2_u12_u5_n131 ) );
  INV_X1 u2_u12_u5_U74 (.A( u2_u12_u5_n102 ) , .ZN( u2_u12_u5_n195 ) );
  OAI221_X1 u2_u12_u5_U75 (.A( u2_u12_u5_n101 ) , .ZN( u2_u12_u5_n102 ) , .C2( u2_u12_u5_n115 ) , .C1( u2_u12_u5_n126 ) , .B1( u2_u12_u5_n134 ) , .B2( u2_u12_u5_n160 ) );
  OAI21_X1 u2_u12_u5_U76 (.ZN( u2_u12_u5_n101 ) , .B1( u2_u12_u5_n137 ) , .A( u2_u12_u5_n146 ) , .B2( u2_u12_u5_n147 ) );
  NOR2_X1 u2_u12_u5_U77 (.A2( u2_u12_X_34 ) , .A1( u2_u12_X_35 ) , .ZN( u2_u12_u5_n145 ) );
  NOR2_X1 u2_u12_u5_U78 (.A2( u2_u12_X_34 ) , .ZN( u2_u12_u5_n146 ) , .A1( u2_u12_u5_n171 ) );
  NOR2_X1 u2_u12_u5_U79 (.A2( u2_u12_X_31 ) , .A1( u2_u12_X_32 ) , .ZN( u2_u12_u5_n103 ) );
  NOR3_X1 u2_u12_u5_U8 (.A2( u2_u12_u5_n147 ) , .A1( u2_u12_u5_n148 ) , .ZN( u2_u12_u5_n149 ) , .A3( u2_u12_u5_n194 ) );
  NOR2_X1 u2_u12_u5_U80 (.A2( u2_u12_X_36 ) , .ZN( u2_u12_u5_n105 ) , .A1( u2_u12_u5_n180 ) );
  NOR2_X1 u2_u12_u5_U81 (.A2( u2_u12_X_33 ) , .ZN( u2_u12_u5_n108 ) , .A1( u2_u12_u5_n170 ) );
  NOR2_X1 u2_u12_u5_U82 (.A2( u2_u12_X_33 ) , .A1( u2_u12_X_36 ) , .ZN( u2_u12_u5_n107 ) );
  NOR2_X1 u2_u12_u5_U83 (.A2( u2_u12_X_31 ) , .ZN( u2_u12_u5_n104 ) , .A1( u2_u12_u5_n181 ) );
  NAND2_X1 u2_u12_u5_U84 (.A2( u2_u12_X_34 ) , .A1( u2_u12_X_35 ) , .ZN( u2_u12_u5_n153 ) );
  NAND2_X1 u2_u12_u5_U85 (.A1( u2_u12_X_34 ) , .ZN( u2_u12_u5_n126 ) , .A2( u2_u12_u5_n171 ) );
  AND2_X1 u2_u12_u5_U86 (.A1( u2_u12_X_31 ) , .A2( u2_u12_X_32 ) , .ZN( u2_u12_u5_n106 ) );
  AND2_X1 u2_u12_u5_U87 (.A1( u2_u12_X_31 ) , .ZN( u2_u12_u5_n109 ) , .A2( u2_u12_u5_n181 ) );
  INV_X1 u2_u12_u5_U88 (.A( u2_u12_X_33 ) , .ZN( u2_u12_u5_n180 ) );
  INV_X1 u2_u12_u5_U89 (.A( u2_u12_X_35 ) , .ZN( u2_u12_u5_n171 ) );
  NOR2_X1 u2_u12_u5_U9 (.ZN( u2_u12_u5_n135 ) , .A1( u2_u12_u5_n173 ) , .A2( u2_u12_u5_n176 ) );
  INV_X1 u2_u12_u5_U90 (.A( u2_u12_X_36 ) , .ZN( u2_u12_u5_n170 ) );
  INV_X1 u2_u12_u5_U91 (.A( u2_u12_X_32 ) , .ZN( u2_u12_u5_n181 ) );
  NAND4_X1 u2_u12_u5_U92 (.ZN( u2_out12_29 ) , .A4( u2_u12_u5_n129 ) , .A3( u2_u12_u5_n130 ) , .A2( u2_u12_u5_n168 ) , .A1( u2_u12_u5_n196 ) );
  AOI221_X1 u2_u12_u5_U93 (.A( u2_u12_u5_n128 ) , .ZN( u2_u12_u5_n129 ) , .C2( u2_u12_u5_n132 ) , .B2( u2_u12_u5_n159 ) , .B1( u2_u12_u5_n176 ) , .C1( u2_u12_u5_n184 ) );
  AOI222_X1 u2_u12_u5_U94 (.ZN( u2_u12_u5_n130 ) , .A2( u2_u12_u5_n146 ) , .B1( u2_u12_u5_n147 ) , .C2( u2_u12_u5_n175 ) , .B2( u2_u12_u5_n179 ) , .A1( u2_u12_u5_n188 ) , .C1( u2_u12_u5_n194 ) );
  NAND4_X1 u2_u12_u5_U95 (.ZN( u2_out12_19 ) , .A4( u2_u12_u5_n166 ) , .A3( u2_u12_u5_n167 ) , .A2( u2_u12_u5_n168 ) , .A1( u2_u12_u5_n169 ) );
  AOI22_X1 u2_u12_u5_U96 (.B2( u2_u12_u5_n145 ) , .A2( u2_u12_u5_n146 ) , .ZN( u2_u12_u5_n167 ) , .B1( u2_u12_u5_n182 ) , .A1( u2_u12_u5_n189 ) );
  NOR4_X1 u2_u12_u5_U97 (.A4( u2_u12_u5_n162 ) , .A3( u2_u12_u5_n163 ) , .A2( u2_u12_u5_n164 ) , .A1( u2_u12_u5_n165 ) , .ZN( u2_u12_u5_n166 ) );
  NAND4_X1 u2_u12_u5_U98 (.ZN( u2_out12_11 ) , .A4( u2_u12_u5_n143 ) , .A3( u2_u12_u5_n144 ) , .A2( u2_u12_u5_n169 ) , .A1( u2_u12_u5_n196 ) );
  AOI22_X1 u2_u12_u5_U99 (.A2( u2_u12_u5_n132 ) , .ZN( u2_u12_u5_n144 ) , .B2( u2_u12_u5_n145 ) , .B1( u2_u12_u5_n184 ) , .A1( u2_u12_u5_n194 ) );
  AOI22_X1 u2_u12_u6_U10 (.A2( u2_u12_u6_n151 ) , .B2( u2_u12_u6_n161 ) , .A1( u2_u12_u6_n167 ) , .B1( u2_u12_u6_n170 ) , .ZN( u2_u12_u6_n89 ) );
  AOI21_X1 u2_u12_u6_U11 (.B1( u2_u12_u6_n107 ) , .B2( u2_u12_u6_n132 ) , .A( u2_u12_u6_n158 ) , .ZN( u2_u12_u6_n88 ) );
  AOI21_X1 u2_u12_u6_U12 (.B2( u2_u12_u6_n147 ) , .B1( u2_u12_u6_n148 ) , .ZN( u2_u12_u6_n149 ) , .A( u2_u12_u6_n158 ) );
  AOI21_X1 u2_u12_u6_U13 (.ZN( u2_u12_u6_n106 ) , .A( u2_u12_u6_n142 ) , .B2( u2_u12_u6_n159 ) , .B1( u2_u12_u6_n164 ) );
  INV_X1 u2_u12_u6_U14 (.A( u2_u12_u6_n155 ) , .ZN( u2_u12_u6_n161 ) );
  INV_X1 u2_u12_u6_U15 (.A( u2_u12_u6_n128 ) , .ZN( u2_u12_u6_n164 ) );
  NAND2_X1 u2_u12_u6_U16 (.ZN( u2_u12_u6_n110 ) , .A1( u2_u12_u6_n122 ) , .A2( u2_u12_u6_n129 ) );
  NAND2_X1 u2_u12_u6_U17 (.ZN( u2_u12_u6_n124 ) , .A2( u2_u12_u6_n146 ) , .A1( u2_u12_u6_n148 ) );
  INV_X1 u2_u12_u6_U18 (.A( u2_u12_u6_n132 ) , .ZN( u2_u12_u6_n171 ) );
  AND2_X1 u2_u12_u6_U19 (.A1( u2_u12_u6_n100 ) , .ZN( u2_u12_u6_n130 ) , .A2( u2_u12_u6_n147 ) );
  INV_X1 u2_u12_u6_U20 (.A( u2_u12_u6_n127 ) , .ZN( u2_u12_u6_n173 ) );
  INV_X1 u2_u12_u6_U21 (.A( u2_u12_u6_n121 ) , .ZN( u2_u12_u6_n167 ) );
  INV_X1 u2_u12_u6_U22 (.A( u2_u12_u6_n100 ) , .ZN( u2_u12_u6_n169 ) );
  INV_X1 u2_u12_u6_U23 (.A( u2_u12_u6_n123 ) , .ZN( u2_u12_u6_n170 ) );
  INV_X1 u2_u12_u6_U24 (.A( u2_u12_u6_n113 ) , .ZN( u2_u12_u6_n168 ) );
  AND2_X1 u2_u12_u6_U25 (.A1( u2_u12_u6_n107 ) , .A2( u2_u12_u6_n119 ) , .ZN( u2_u12_u6_n133 ) );
  AND2_X1 u2_u12_u6_U26 (.A2( u2_u12_u6_n121 ) , .A1( u2_u12_u6_n122 ) , .ZN( u2_u12_u6_n131 ) );
  AND3_X1 u2_u12_u6_U27 (.ZN( u2_u12_u6_n120 ) , .A2( u2_u12_u6_n127 ) , .A1( u2_u12_u6_n132 ) , .A3( u2_u12_u6_n145 ) );
  INV_X1 u2_u12_u6_U28 (.A( u2_u12_u6_n146 ) , .ZN( u2_u12_u6_n163 ) );
  AOI222_X1 u2_u12_u6_U29 (.ZN( u2_u12_u6_n114 ) , .A1( u2_u12_u6_n118 ) , .A2( u2_u12_u6_n126 ) , .B2( u2_u12_u6_n151 ) , .C2( u2_u12_u6_n159 ) , .C1( u2_u12_u6_n168 ) , .B1( u2_u12_u6_n169 ) );
  INV_X1 u2_u12_u6_U3 (.A( u2_u12_u6_n110 ) , .ZN( u2_u12_u6_n166 ) );
  NOR2_X1 u2_u12_u6_U30 (.A1( u2_u12_u6_n162 ) , .A2( u2_u12_u6_n165 ) , .ZN( u2_u12_u6_n98 ) );
  AOI211_X1 u2_u12_u6_U31 (.B( u2_u12_u6_n134 ) , .A( u2_u12_u6_n135 ) , .C1( u2_u12_u6_n136 ) , .ZN( u2_u12_u6_n137 ) , .C2( u2_u12_u6_n151 ) );
  AOI21_X1 u2_u12_u6_U32 (.B2( u2_u12_u6_n132 ) , .B1( u2_u12_u6_n133 ) , .ZN( u2_u12_u6_n134 ) , .A( u2_u12_u6_n158 ) );
  AOI21_X1 u2_u12_u6_U33 (.B1( u2_u12_u6_n131 ) , .ZN( u2_u12_u6_n135 ) , .A( u2_u12_u6_n144 ) , .B2( u2_u12_u6_n146 ) );
  NAND4_X1 u2_u12_u6_U34 (.A4( u2_u12_u6_n127 ) , .A3( u2_u12_u6_n128 ) , .A2( u2_u12_u6_n129 ) , .A1( u2_u12_u6_n130 ) , .ZN( u2_u12_u6_n136 ) );
  NAND2_X1 u2_u12_u6_U35 (.A1( u2_u12_u6_n144 ) , .ZN( u2_u12_u6_n151 ) , .A2( u2_u12_u6_n158 ) );
  NAND2_X1 u2_u12_u6_U36 (.ZN( u2_u12_u6_n132 ) , .A1( u2_u12_u6_n91 ) , .A2( u2_u12_u6_n97 ) );
  AOI22_X1 u2_u12_u6_U37 (.B2( u2_u12_u6_n110 ) , .B1( u2_u12_u6_n111 ) , .A1( u2_u12_u6_n112 ) , .ZN( u2_u12_u6_n115 ) , .A2( u2_u12_u6_n161 ) );
  NAND4_X1 u2_u12_u6_U38 (.A3( u2_u12_u6_n109 ) , .ZN( u2_u12_u6_n112 ) , .A4( u2_u12_u6_n132 ) , .A2( u2_u12_u6_n147 ) , .A1( u2_u12_u6_n166 ) );
  NOR2_X1 u2_u12_u6_U39 (.ZN( u2_u12_u6_n109 ) , .A1( u2_u12_u6_n170 ) , .A2( u2_u12_u6_n173 ) );
  INV_X1 u2_u12_u6_U4 (.A( u2_u12_u6_n142 ) , .ZN( u2_u12_u6_n174 ) );
  NOR2_X1 u2_u12_u6_U40 (.A2( u2_u12_u6_n126 ) , .ZN( u2_u12_u6_n155 ) , .A1( u2_u12_u6_n160 ) );
  NAND2_X1 u2_u12_u6_U41 (.ZN( u2_u12_u6_n146 ) , .A2( u2_u12_u6_n94 ) , .A1( u2_u12_u6_n99 ) );
  AOI21_X1 u2_u12_u6_U42 (.A( u2_u12_u6_n144 ) , .B2( u2_u12_u6_n145 ) , .B1( u2_u12_u6_n146 ) , .ZN( u2_u12_u6_n150 ) );
  INV_X1 u2_u12_u6_U43 (.A( u2_u12_u6_n111 ) , .ZN( u2_u12_u6_n158 ) );
  NAND2_X1 u2_u12_u6_U44 (.ZN( u2_u12_u6_n127 ) , .A1( u2_u12_u6_n91 ) , .A2( u2_u12_u6_n92 ) );
  NAND2_X1 u2_u12_u6_U45 (.ZN( u2_u12_u6_n129 ) , .A2( u2_u12_u6_n95 ) , .A1( u2_u12_u6_n96 ) );
  INV_X1 u2_u12_u6_U46 (.A( u2_u12_u6_n144 ) , .ZN( u2_u12_u6_n159 ) );
  NAND2_X1 u2_u12_u6_U47 (.ZN( u2_u12_u6_n145 ) , .A2( u2_u12_u6_n97 ) , .A1( u2_u12_u6_n98 ) );
  NAND2_X1 u2_u12_u6_U48 (.ZN( u2_u12_u6_n148 ) , .A2( u2_u12_u6_n92 ) , .A1( u2_u12_u6_n94 ) );
  NAND2_X1 u2_u12_u6_U49 (.ZN( u2_u12_u6_n108 ) , .A2( u2_u12_u6_n139 ) , .A1( u2_u12_u6_n144 ) );
  NAND2_X1 u2_u12_u6_U5 (.A2( u2_u12_u6_n143 ) , .ZN( u2_u12_u6_n152 ) , .A1( u2_u12_u6_n166 ) );
  NAND2_X1 u2_u12_u6_U50 (.ZN( u2_u12_u6_n121 ) , .A2( u2_u12_u6_n95 ) , .A1( u2_u12_u6_n97 ) );
  NAND2_X1 u2_u12_u6_U51 (.ZN( u2_u12_u6_n107 ) , .A2( u2_u12_u6_n92 ) , .A1( u2_u12_u6_n95 ) );
  AND2_X1 u2_u12_u6_U52 (.ZN( u2_u12_u6_n118 ) , .A2( u2_u12_u6_n91 ) , .A1( u2_u12_u6_n99 ) );
  NAND2_X1 u2_u12_u6_U53 (.ZN( u2_u12_u6_n147 ) , .A2( u2_u12_u6_n98 ) , .A1( u2_u12_u6_n99 ) );
  NAND2_X1 u2_u12_u6_U54 (.ZN( u2_u12_u6_n128 ) , .A1( u2_u12_u6_n94 ) , .A2( u2_u12_u6_n96 ) );
  NAND2_X1 u2_u12_u6_U55 (.ZN( u2_u12_u6_n119 ) , .A2( u2_u12_u6_n95 ) , .A1( u2_u12_u6_n99 ) );
  NAND2_X1 u2_u12_u6_U56 (.ZN( u2_u12_u6_n123 ) , .A2( u2_u12_u6_n91 ) , .A1( u2_u12_u6_n96 ) );
  NAND2_X1 u2_u12_u6_U57 (.ZN( u2_u12_u6_n100 ) , .A2( u2_u12_u6_n92 ) , .A1( u2_u12_u6_n98 ) );
  NAND2_X1 u2_u12_u6_U58 (.ZN( u2_u12_u6_n122 ) , .A1( u2_u12_u6_n94 ) , .A2( u2_u12_u6_n97 ) );
  INV_X1 u2_u12_u6_U59 (.A( u2_u12_u6_n139 ) , .ZN( u2_u12_u6_n160 ) );
  AOI22_X1 u2_u12_u6_U6 (.B2( u2_u12_u6_n101 ) , .A1( u2_u12_u6_n102 ) , .ZN( u2_u12_u6_n103 ) , .B1( u2_u12_u6_n160 ) , .A2( u2_u12_u6_n161 ) );
  NAND2_X1 u2_u12_u6_U60 (.ZN( u2_u12_u6_n113 ) , .A1( u2_u12_u6_n96 ) , .A2( u2_u12_u6_n98 ) );
  NOR2_X1 u2_u12_u6_U61 (.A2( u2_u12_X_40 ) , .A1( u2_u12_X_41 ) , .ZN( u2_u12_u6_n126 ) );
  NOR2_X1 u2_u12_u6_U62 (.A2( u2_u12_X_39 ) , .A1( u2_u12_X_42 ) , .ZN( u2_u12_u6_n92 ) );
  NOR2_X1 u2_u12_u6_U63 (.A2( u2_u12_X_39 ) , .A1( u2_u12_u6_n156 ) , .ZN( u2_u12_u6_n97 ) );
  NOR2_X1 u2_u12_u6_U64 (.A2( u2_u12_X_38 ) , .A1( u2_u12_u6_n165 ) , .ZN( u2_u12_u6_n95 ) );
  NOR2_X1 u2_u12_u6_U65 (.A2( u2_u12_X_41 ) , .ZN( u2_u12_u6_n111 ) , .A1( u2_u12_u6_n157 ) );
  NOR2_X1 u2_u12_u6_U66 (.A2( u2_u12_X_37 ) , .A1( u2_u12_u6_n162 ) , .ZN( u2_u12_u6_n94 ) );
  NOR2_X1 u2_u12_u6_U67 (.A2( u2_u12_X_37 ) , .A1( u2_u12_X_38 ) , .ZN( u2_u12_u6_n91 ) );
  NAND2_X1 u2_u12_u6_U68 (.A1( u2_u12_X_41 ) , .ZN( u2_u12_u6_n144 ) , .A2( u2_u12_u6_n157 ) );
  NAND2_X1 u2_u12_u6_U69 (.A2( u2_u12_X_40 ) , .A1( u2_u12_X_41 ) , .ZN( u2_u12_u6_n139 ) );
  NOR2_X1 u2_u12_u6_U7 (.A1( u2_u12_u6_n118 ) , .ZN( u2_u12_u6_n143 ) , .A2( u2_u12_u6_n168 ) );
  AND2_X1 u2_u12_u6_U70 (.A1( u2_u12_X_39 ) , .A2( u2_u12_u6_n156 ) , .ZN( u2_u12_u6_n96 ) );
  AND2_X1 u2_u12_u6_U71 (.A1( u2_u12_X_39 ) , .A2( u2_u12_X_42 ) , .ZN( u2_u12_u6_n99 ) );
  INV_X1 u2_u12_u6_U72 (.A( u2_u12_X_40 ) , .ZN( u2_u12_u6_n157 ) );
  INV_X1 u2_u12_u6_U73 (.A( u2_u12_X_37 ) , .ZN( u2_u12_u6_n165 ) );
  INV_X1 u2_u12_u6_U74 (.A( u2_u12_X_38 ) , .ZN( u2_u12_u6_n162 ) );
  INV_X1 u2_u12_u6_U75 (.A( u2_u12_X_42 ) , .ZN( u2_u12_u6_n156 ) );
  NAND4_X1 u2_u12_u6_U76 (.ZN( u2_out12_32 ) , .A4( u2_u12_u6_n103 ) , .A3( u2_u12_u6_n104 ) , .A2( u2_u12_u6_n105 ) , .A1( u2_u12_u6_n106 ) );
  AOI22_X1 u2_u12_u6_U77 (.ZN( u2_u12_u6_n105 ) , .A2( u2_u12_u6_n108 ) , .A1( u2_u12_u6_n118 ) , .B2( u2_u12_u6_n126 ) , .B1( u2_u12_u6_n171 ) );
  AOI22_X1 u2_u12_u6_U78 (.ZN( u2_u12_u6_n104 ) , .A1( u2_u12_u6_n111 ) , .B1( u2_u12_u6_n124 ) , .B2( u2_u12_u6_n151 ) , .A2( u2_u12_u6_n93 ) );
  NAND4_X1 u2_u12_u6_U79 (.ZN( u2_out12_12 ) , .A4( u2_u12_u6_n114 ) , .A3( u2_u12_u6_n115 ) , .A2( u2_u12_u6_n116 ) , .A1( u2_u12_u6_n117 ) );
  INV_X1 u2_u12_u6_U8 (.ZN( u2_u12_u6_n172 ) , .A( u2_u12_u6_n88 ) );
  OAI22_X1 u2_u12_u6_U80 (.B2( u2_u12_u6_n111 ) , .ZN( u2_u12_u6_n116 ) , .B1( u2_u12_u6_n126 ) , .A2( u2_u12_u6_n164 ) , .A1( u2_u12_u6_n167 ) );
  OAI21_X1 u2_u12_u6_U81 (.A( u2_u12_u6_n108 ) , .ZN( u2_u12_u6_n117 ) , .B2( u2_u12_u6_n141 ) , .B1( u2_u12_u6_n163 ) );
  OAI211_X1 u2_u12_u6_U82 (.ZN( u2_out12_22 ) , .B( u2_u12_u6_n137 ) , .A( u2_u12_u6_n138 ) , .C2( u2_u12_u6_n139 ) , .C1( u2_u12_u6_n140 ) );
  AOI22_X1 u2_u12_u6_U83 (.B1( u2_u12_u6_n124 ) , .A2( u2_u12_u6_n125 ) , .A1( u2_u12_u6_n126 ) , .ZN( u2_u12_u6_n138 ) , .B2( u2_u12_u6_n161 ) );
  AND4_X1 u2_u12_u6_U84 (.A3( u2_u12_u6_n119 ) , .A1( u2_u12_u6_n120 ) , .A4( u2_u12_u6_n129 ) , .ZN( u2_u12_u6_n140 ) , .A2( u2_u12_u6_n143 ) );
  OAI211_X1 u2_u12_u6_U85 (.ZN( u2_out12_7 ) , .B( u2_u12_u6_n153 ) , .C2( u2_u12_u6_n154 ) , .C1( u2_u12_u6_n155 ) , .A( u2_u12_u6_n174 ) );
  NOR3_X1 u2_u12_u6_U86 (.A1( u2_u12_u6_n141 ) , .ZN( u2_u12_u6_n154 ) , .A3( u2_u12_u6_n164 ) , .A2( u2_u12_u6_n171 ) );
  AOI211_X1 u2_u12_u6_U87 (.B( u2_u12_u6_n149 ) , .A( u2_u12_u6_n150 ) , .C2( u2_u12_u6_n151 ) , .C1( u2_u12_u6_n152 ) , .ZN( u2_u12_u6_n153 ) );
  NAND3_X1 u2_u12_u6_U88 (.A2( u2_u12_u6_n123 ) , .ZN( u2_u12_u6_n125 ) , .A1( u2_u12_u6_n130 ) , .A3( u2_u12_u6_n131 ) );
  NAND3_X1 u2_u12_u6_U89 (.A3( u2_u12_u6_n133 ) , .ZN( u2_u12_u6_n141 ) , .A1( u2_u12_u6_n145 ) , .A2( u2_u12_u6_n148 ) );
  OAI21_X1 u2_u12_u6_U9 (.A( u2_u12_u6_n159 ) , .B1( u2_u12_u6_n169 ) , .B2( u2_u12_u6_n173 ) , .ZN( u2_u12_u6_n90 ) );
  NAND3_X1 u2_u12_u6_U90 (.ZN( u2_u12_u6_n101 ) , .A3( u2_u12_u6_n107 ) , .A2( u2_u12_u6_n121 ) , .A1( u2_u12_u6_n127 ) );
  NAND3_X1 u2_u12_u6_U91 (.ZN( u2_u12_u6_n102 ) , .A3( u2_u12_u6_n130 ) , .A2( u2_u12_u6_n145 ) , .A1( u2_u12_u6_n166 ) );
  NAND3_X1 u2_u12_u6_U92 (.A3( u2_u12_u6_n113 ) , .A1( u2_u12_u6_n119 ) , .A2( u2_u12_u6_n123 ) , .ZN( u2_u12_u6_n93 ) );
  NAND3_X1 u2_u12_u6_U93 (.ZN( u2_u12_u6_n142 ) , .A2( u2_u12_u6_n172 ) , .A3( u2_u12_u6_n89 ) , .A1( u2_u12_u6_n90 ) );
  AND3_X1 u2_u12_u7_U10 (.A3( u2_u12_u7_n110 ) , .A2( u2_u12_u7_n127 ) , .A1( u2_u12_u7_n132 ) , .ZN( u2_u12_u7_n92 ) );
  OAI21_X1 u2_u12_u7_U11 (.A( u2_u12_u7_n161 ) , .B1( u2_u12_u7_n168 ) , .B2( u2_u12_u7_n173 ) , .ZN( u2_u12_u7_n91 ) );
  AOI211_X1 u2_u12_u7_U12 (.A( u2_u12_u7_n117 ) , .ZN( u2_u12_u7_n118 ) , .C2( u2_u12_u7_n126 ) , .C1( u2_u12_u7_n177 ) , .B( u2_u12_u7_n180 ) );
  OAI22_X1 u2_u12_u7_U13 (.B1( u2_u12_u7_n115 ) , .ZN( u2_u12_u7_n117 ) , .A2( u2_u12_u7_n133 ) , .A1( u2_u12_u7_n137 ) , .B2( u2_u12_u7_n162 ) );
  INV_X1 u2_u12_u7_U14 (.A( u2_u12_u7_n116 ) , .ZN( u2_u12_u7_n180 ) );
  NOR3_X1 u2_u12_u7_U15 (.ZN( u2_u12_u7_n115 ) , .A3( u2_u12_u7_n145 ) , .A2( u2_u12_u7_n168 ) , .A1( u2_u12_u7_n169 ) );
  OAI211_X1 u2_u12_u7_U16 (.B( u2_u12_u7_n122 ) , .A( u2_u12_u7_n123 ) , .C2( u2_u12_u7_n124 ) , .ZN( u2_u12_u7_n154 ) , .C1( u2_u12_u7_n162 ) );
  AOI222_X1 u2_u12_u7_U17 (.ZN( u2_u12_u7_n122 ) , .C2( u2_u12_u7_n126 ) , .C1( u2_u12_u7_n145 ) , .B1( u2_u12_u7_n161 ) , .A2( u2_u12_u7_n165 ) , .B2( u2_u12_u7_n170 ) , .A1( u2_u12_u7_n176 ) );
  INV_X1 u2_u12_u7_U18 (.A( u2_u12_u7_n133 ) , .ZN( u2_u12_u7_n176 ) );
  NOR3_X1 u2_u12_u7_U19 (.A2( u2_u12_u7_n134 ) , .A1( u2_u12_u7_n135 ) , .ZN( u2_u12_u7_n136 ) , .A3( u2_u12_u7_n171 ) );
  NOR2_X1 u2_u12_u7_U20 (.A1( u2_u12_u7_n130 ) , .A2( u2_u12_u7_n134 ) , .ZN( u2_u12_u7_n153 ) );
  INV_X1 u2_u12_u7_U21 (.A( u2_u12_u7_n101 ) , .ZN( u2_u12_u7_n165 ) );
  NOR2_X1 u2_u12_u7_U22 (.ZN( u2_u12_u7_n111 ) , .A2( u2_u12_u7_n134 ) , .A1( u2_u12_u7_n169 ) );
  AOI21_X1 u2_u12_u7_U23 (.ZN( u2_u12_u7_n104 ) , .B2( u2_u12_u7_n112 ) , .B1( u2_u12_u7_n127 ) , .A( u2_u12_u7_n164 ) );
  AOI21_X1 u2_u12_u7_U24 (.ZN( u2_u12_u7_n106 ) , .B1( u2_u12_u7_n133 ) , .B2( u2_u12_u7_n146 ) , .A( u2_u12_u7_n162 ) );
  AOI21_X1 u2_u12_u7_U25 (.A( u2_u12_u7_n101 ) , .ZN( u2_u12_u7_n107 ) , .B2( u2_u12_u7_n128 ) , .B1( u2_u12_u7_n175 ) );
  INV_X1 u2_u12_u7_U26 (.A( u2_u12_u7_n138 ) , .ZN( u2_u12_u7_n171 ) );
  INV_X1 u2_u12_u7_U27 (.A( u2_u12_u7_n131 ) , .ZN( u2_u12_u7_n177 ) );
  INV_X1 u2_u12_u7_U28 (.A( u2_u12_u7_n110 ) , .ZN( u2_u12_u7_n174 ) );
  NAND2_X1 u2_u12_u7_U29 (.A1( u2_u12_u7_n129 ) , .A2( u2_u12_u7_n132 ) , .ZN( u2_u12_u7_n149 ) );
  OAI21_X1 u2_u12_u7_U3 (.ZN( u2_u12_u7_n159 ) , .A( u2_u12_u7_n165 ) , .B2( u2_u12_u7_n171 ) , .B1( u2_u12_u7_n174 ) );
  NAND2_X1 u2_u12_u7_U30 (.A1( u2_u12_u7_n113 ) , .A2( u2_u12_u7_n124 ) , .ZN( u2_u12_u7_n130 ) );
  INV_X1 u2_u12_u7_U31 (.A( u2_u12_u7_n112 ) , .ZN( u2_u12_u7_n173 ) );
  INV_X1 u2_u12_u7_U32 (.A( u2_u12_u7_n128 ) , .ZN( u2_u12_u7_n168 ) );
  INV_X1 u2_u12_u7_U33 (.A( u2_u12_u7_n148 ) , .ZN( u2_u12_u7_n169 ) );
  INV_X1 u2_u12_u7_U34 (.A( u2_u12_u7_n127 ) , .ZN( u2_u12_u7_n179 ) );
  NOR2_X1 u2_u12_u7_U35 (.ZN( u2_u12_u7_n101 ) , .A2( u2_u12_u7_n150 ) , .A1( u2_u12_u7_n156 ) );
  AOI211_X1 u2_u12_u7_U36 (.B( u2_u12_u7_n154 ) , .A( u2_u12_u7_n155 ) , .C1( u2_u12_u7_n156 ) , .ZN( u2_u12_u7_n157 ) , .C2( u2_u12_u7_n172 ) );
  INV_X1 u2_u12_u7_U37 (.A( u2_u12_u7_n153 ) , .ZN( u2_u12_u7_n172 ) );
  AOI211_X1 u2_u12_u7_U38 (.B( u2_u12_u7_n139 ) , .A( u2_u12_u7_n140 ) , .C2( u2_u12_u7_n141 ) , .ZN( u2_u12_u7_n142 ) , .C1( u2_u12_u7_n156 ) );
  NAND4_X1 u2_u12_u7_U39 (.A3( u2_u12_u7_n127 ) , .A2( u2_u12_u7_n128 ) , .A1( u2_u12_u7_n129 ) , .ZN( u2_u12_u7_n141 ) , .A4( u2_u12_u7_n147 ) );
  INV_X1 u2_u12_u7_U4 (.A( u2_u12_u7_n111 ) , .ZN( u2_u12_u7_n170 ) );
  AOI21_X1 u2_u12_u7_U40 (.A( u2_u12_u7_n137 ) , .B1( u2_u12_u7_n138 ) , .ZN( u2_u12_u7_n139 ) , .B2( u2_u12_u7_n146 ) );
  OAI22_X1 u2_u12_u7_U41 (.B1( u2_u12_u7_n136 ) , .ZN( u2_u12_u7_n140 ) , .A1( u2_u12_u7_n153 ) , .B2( u2_u12_u7_n162 ) , .A2( u2_u12_u7_n164 ) );
  AOI21_X1 u2_u12_u7_U42 (.ZN( u2_u12_u7_n123 ) , .B1( u2_u12_u7_n165 ) , .B2( u2_u12_u7_n177 ) , .A( u2_u12_u7_n97 ) );
  AOI21_X1 u2_u12_u7_U43 (.B2( u2_u12_u7_n113 ) , .B1( u2_u12_u7_n124 ) , .A( u2_u12_u7_n125 ) , .ZN( u2_u12_u7_n97 ) );
  INV_X1 u2_u12_u7_U44 (.A( u2_u12_u7_n125 ) , .ZN( u2_u12_u7_n161 ) );
  INV_X1 u2_u12_u7_U45 (.A( u2_u12_u7_n152 ) , .ZN( u2_u12_u7_n162 ) );
  AOI22_X1 u2_u12_u7_U46 (.A2( u2_u12_u7_n114 ) , .ZN( u2_u12_u7_n119 ) , .B1( u2_u12_u7_n130 ) , .A1( u2_u12_u7_n156 ) , .B2( u2_u12_u7_n165 ) );
  NAND2_X1 u2_u12_u7_U47 (.A2( u2_u12_u7_n112 ) , .ZN( u2_u12_u7_n114 ) , .A1( u2_u12_u7_n175 ) );
  AND2_X1 u2_u12_u7_U48 (.ZN( u2_u12_u7_n145 ) , .A2( u2_u12_u7_n98 ) , .A1( u2_u12_u7_n99 ) );
  NOR2_X1 u2_u12_u7_U49 (.ZN( u2_u12_u7_n137 ) , .A1( u2_u12_u7_n150 ) , .A2( u2_u12_u7_n161 ) );
  INV_X1 u2_u12_u7_U5 (.A( u2_u12_u7_n149 ) , .ZN( u2_u12_u7_n175 ) );
  AOI21_X1 u2_u12_u7_U50 (.ZN( u2_u12_u7_n105 ) , .B2( u2_u12_u7_n110 ) , .A( u2_u12_u7_n125 ) , .B1( u2_u12_u7_n147 ) );
  NAND2_X1 u2_u12_u7_U51 (.ZN( u2_u12_u7_n146 ) , .A1( u2_u12_u7_n95 ) , .A2( u2_u12_u7_n98 ) );
  NAND2_X1 u2_u12_u7_U52 (.A2( u2_u12_u7_n103 ) , .ZN( u2_u12_u7_n147 ) , .A1( u2_u12_u7_n93 ) );
  NAND2_X1 u2_u12_u7_U53 (.A1( u2_u12_u7_n103 ) , .ZN( u2_u12_u7_n127 ) , .A2( u2_u12_u7_n99 ) );
  OR2_X1 u2_u12_u7_U54 (.ZN( u2_u12_u7_n126 ) , .A2( u2_u12_u7_n152 ) , .A1( u2_u12_u7_n156 ) );
  NAND2_X1 u2_u12_u7_U55 (.A2( u2_u12_u7_n102 ) , .A1( u2_u12_u7_n103 ) , .ZN( u2_u12_u7_n133 ) );
  NAND2_X1 u2_u12_u7_U56 (.ZN( u2_u12_u7_n112 ) , .A2( u2_u12_u7_n96 ) , .A1( u2_u12_u7_n99 ) );
  NAND2_X1 u2_u12_u7_U57 (.A2( u2_u12_u7_n102 ) , .ZN( u2_u12_u7_n128 ) , .A1( u2_u12_u7_n98 ) );
  NAND2_X1 u2_u12_u7_U58 (.A1( u2_u12_u7_n100 ) , .ZN( u2_u12_u7_n113 ) , .A2( u2_u12_u7_n93 ) );
  NAND2_X1 u2_u12_u7_U59 (.A2( u2_u12_u7_n102 ) , .ZN( u2_u12_u7_n124 ) , .A1( u2_u12_u7_n96 ) );
  INV_X1 u2_u12_u7_U6 (.A( u2_u12_u7_n154 ) , .ZN( u2_u12_u7_n178 ) );
  NAND2_X1 u2_u12_u7_U60 (.ZN( u2_u12_u7_n110 ) , .A1( u2_u12_u7_n95 ) , .A2( u2_u12_u7_n96 ) );
  INV_X1 u2_u12_u7_U61 (.A( u2_u12_u7_n150 ) , .ZN( u2_u12_u7_n164 ) );
  AND2_X1 u2_u12_u7_U62 (.ZN( u2_u12_u7_n134 ) , .A1( u2_u12_u7_n93 ) , .A2( u2_u12_u7_n98 ) );
  NAND2_X1 u2_u12_u7_U63 (.A1( u2_u12_u7_n100 ) , .A2( u2_u12_u7_n102 ) , .ZN( u2_u12_u7_n129 ) );
  NAND2_X1 u2_u12_u7_U64 (.A2( u2_u12_u7_n103 ) , .ZN( u2_u12_u7_n131 ) , .A1( u2_u12_u7_n95 ) );
  NAND2_X1 u2_u12_u7_U65 (.A1( u2_u12_u7_n100 ) , .ZN( u2_u12_u7_n138 ) , .A2( u2_u12_u7_n99 ) );
  NAND2_X1 u2_u12_u7_U66 (.ZN( u2_u12_u7_n132 ) , .A1( u2_u12_u7_n93 ) , .A2( u2_u12_u7_n96 ) );
  NAND2_X1 u2_u12_u7_U67 (.A1( u2_u12_u7_n100 ) , .ZN( u2_u12_u7_n148 ) , .A2( u2_u12_u7_n95 ) );
  NOR2_X1 u2_u12_u7_U68 (.A2( u2_u12_X_47 ) , .ZN( u2_u12_u7_n150 ) , .A1( u2_u12_u7_n163 ) );
  NOR2_X1 u2_u12_u7_U69 (.A2( u2_u12_X_43 ) , .A1( u2_u12_X_44 ) , .ZN( u2_u12_u7_n103 ) );
  AOI211_X1 u2_u12_u7_U7 (.ZN( u2_u12_u7_n116 ) , .A( u2_u12_u7_n155 ) , .C1( u2_u12_u7_n161 ) , .C2( u2_u12_u7_n171 ) , .B( u2_u12_u7_n94 ) );
  NOR2_X1 u2_u12_u7_U70 (.A2( u2_u12_X_48 ) , .A1( u2_u12_u7_n166 ) , .ZN( u2_u12_u7_n95 ) );
  NOR2_X1 u2_u12_u7_U71 (.A2( u2_u12_X_45 ) , .A1( u2_u12_X_48 ) , .ZN( u2_u12_u7_n99 ) );
  NOR2_X1 u2_u12_u7_U72 (.A2( u2_u12_X_44 ) , .A1( u2_u12_u7_n167 ) , .ZN( u2_u12_u7_n98 ) );
  NOR2_X1 u2_u12_u7_U73 (.A2( u2_u12_X_46 ) , .A1( u2_u12_X_47 ) , .ZN( u2_u12_u7_n152 ) );
  AND2_X1 u2_u12_u7_U74 (.A1( u2_u12_X_47 ) , .ZN( u2_u12_u7_n156 ) , .A2( u2_u12_u7_n163 ) );
  NAND2_X1 u2_u12_u7_U75 (.A2( u2_u12_X_46 ) , .A1( u2_u12_X_47 ) , .ZN( u2_u12_u7_n125 ) );
  AND2_X1 u2_u12_u7_U76 (.A2( u2_u12_X_45 ) , .A1( u2_u12_X_48 ) , .ZN( u2_u12_u7_n102 ) );
  AND2_X1 u2_u12_u7_U77 (.A2( u2_u12_X_43 ) , .A1( u2_u12_X_44 ) , .ZN( u2_u12_u7_n96 ) );
  AND2_X1 u2_u12_u7_U78 (.A1( u2_u12_X_44 ) , .ZN( u2_u12_u7_n100 ) , .A2( u2_u12_u7_n167 ) );
  AND2_X1 u2_u12_u7_U79 (.A1( u2_u12_X_48 ) , .A2( u2_u12_u7_n166 ) , .ZN( u2_u12_u7_n93 ) );
  OAI222_X1 u2_u12_u7_U8 (.C2( u2_u12_u7_n101 ) , .B2( u2_u12_u7_n111 ) , .A1( u2_u12_u7_n113 ) , .C1( u2_u12_u7_n146 ) , .A2( u2_u12_u7_n162 ) , .B1( u2_u12_u7_n164 ) , .ZN( u2_u12_u7_n94 ) );
  INV_X1 u2_u12_u7_U80 (.A( u2_u12_X_46 ) , .ZN( u2_u12_u7_n163 ) );
  INV_X1 u2_u12_u7_U81 (.A( u2_u12_X_43 ) , .ZN( u2_u12_u7_n167 ) );
  INV_X1 u2_u12_u7_U82 (.A( u2_u12_X_45 ) , .ZN( u2_u12_u7_n166 ) );
  NAND4_X1 u2_u12_u7_U83 (.ZN( u2_out12_27 ) , .A4( u2_u12_u7_n118 ) , .A3( u2_u12_u7_n119 ) , .A2( u2_u12_u7_n120 ) , .A1( u2_u12_u7_n121 ) );
  OAI21_X1 u2_u12_u7_U84 (.ZN( u2_u12_u7_n121 ) , .B2( u2_u12_u7_n145 ) , .A( u2_u12_u7_n150 ) , .B1( u2_u12_u7_n174 ) );
  OAI21_X1 u2_u12_u7_U85 (.ZN( u2_u12_u7_n120 ) , .A( u2_u12_u7_n161 ) , .B2( u2_u12_u7_n170 ) , .B1( u2_u12_u7_n179 ) );
  NAND4_X1 u2_u12_u7_U86 (.ZN( u2_out12_21 ) , .A4( u2_u12_u7_n157 ) , .A3( u2_u12_u7_n158 ) , .A2( u2_u12_u7_n159 ) , .A1( u2_u12_u7_n160 ) );
  OAI21_X1 u2_u12_u7_U87 (.B1( u2_u12_u7_n145 ) , .ZN( u2_u12_u7_n160 ) , .A( u2_u12_u7_n161 ) , .B2( u2_u12_u7_n177 ) );
  AOI22_X1 u2_u12_u7_U88 (.B2( u2_u12_u7_n149 ) , .B1( u2_u12_u7_n150 ) , .A2( u2_u12_u7_n151 ) , .A1( u2_u12_u7_n152 ) , .ZN( u2_u12_u7_n158 ) );
  NAND4_X1 u2_u12_u7_U89 (.ZN( u2_out12_15 ) , .A4( u2_u12_u7_n142 ) , .A3( u2_u12_u7_n143 ) , .A2( u2_u12_u7_n144 ) , .A1( u2_u12_u7_n178 ) );
  OAI221_X1 u2_u12_u7_U9 (.C1( u2_u12_u7_n101 ) , .C2( u2_u12_u7_n147 ) , .ZN( u2_u12_u7_n155 ) , .B2( u2_u12_u7_n162 ) , .A( u2_u12_u7_n91 ) , .B1( u2_u12_u7_n92 ) );
  OR2_X1 u2_u12_u7_U90 (.A2( u2_u12_u7_n125 ) , .A1( u2_u12_u7_n129 ) , .ZN( u2_u12_u7_n144 ) );
  AOI22_X1 u2_u12_u7_U91 (.A2( u2_u12_u7_n126 ) , .ZN( u2_u12_u7_n143 ) , .B2( u2_u12_u7_n165 ) , .B1( u2_u12_u7_n173 ) , .A1( u2_u12_u7_n174 ) );
  NAND4_X1 u2_u12_u7_U92 (.ZN( u2_out12_5 ) , .A4( u2_u12_u7_n108 ) , .A3( u2_u12_u7_n109 ) , .A1( u2_u12_u7_n116 ) , .A2( u2_u12_u7_n123 ) );
  AOI22_X1 u2_u12_u7_U93 (.ZN( u2_u12_u7_n109 ) , .A2( u2_u12_u7_n126 ) , .B2( u2_u12_u7_n145 ) , .B1( u2_u12_u7_n156 ) , .A1( u2_u12_u7_n171 ) );
  NOR4_X1 u2_u12_u7_U94 (.A4( u2_u12_u7_n104 ) , .A3( u2_u12_u7_n105 ) , .A2( u2_u12_u7_n106 ) , .A1( u2_u12_u7_n107 ) , .ZN( u2_u12_u7_n108 ) );
  NAND3_X1 u2_u12_u7_U95 (.A3( u2_u12_u7_n146 ) , .A2( u2_u12_u7_n147 ) , .A1( u2_u12_u7_n148 ) , .ZN( u2_u12_u7_n151 ) );
  NAND3_X1 u2_u12_u7_U96 (.A3( u2_u12_u7_n131 ) , .A2( u2_u12_u7_n132 ) , .A1( u2_u12_u7_n133 ) , .ZN( u2_u12_u7_n135 ) );
  XOR2_X1 u2_u13_U18 (.B( u2_K14_38 ) , .A( u2_R12_25 ) , .Z( u2_u13_X_38 ) );
  XOR2_X1 u2_u13_U20 (.B( u2_K14_36 ) , .A( u2_R12_25 ) , .Z( u2_u13_X_36 ) );
  XOR2_X1 u2_u13_U23 (.B( u2_K14_33 ) , .A( u2_R12_22 ) , .Z( u2_u13_X_33 ) );
  XOR2_X1 u2_u13_U24 (.B( u2_K14_32 ) , .A( u2_R12_21 ) , .Z( u2_u13_X_32 ) );
  XOR2_X1 u2_u13_U25 (.B( u2_K14_31 ) , .A( u2_R12_20 ) , .Z( u2_u13_X_31 ) );
  XOR2_X1 u2_u13_U26 (.B( u2_K14_30 ) , .A( u2_R12_21 ) , .Z( u2_u13_X_30 ) );
  XOR2_X1 u2_u13_U28 (.B( u2_K14_29 ) , .A( u2_R12_20 ) , .Z( u2_u13_X_29 ) );
  AOI21_X1 u2_u13_u4_U10 (.ZN( u2_u13_u4_n106 ) , .B2( u2_u13_u4_n146 ) , .B1( u2_u13_u4_n158 ) , .A( u2_u13_u4_n170 ) );
  AOI21_X1 u2_u13_u4_U11 (.ZN( u2_u13_u4_n108 ) , .B2( u2_u13_u4_n134 ) , .B1( u2_u13_u4_n155 ) , .A( u2_u13_u4_n156 ) );
  AOI21_X1 u2_u13_u4_U12 (.ZN( u2_u13_u4_n109 ) , .A( u2_u13_u4_n153 ) , .B1( u2_u13_u4_n159 ) , .B2( u2_u13_u4_n184 ) );
  AOI211_X1 u2_u13_u4_U13 (.B( u2_u13_u4_n136 ) , .A( u2_u13_u4_n137 ) , .C2( u2_u13_u4_n138 ) , .ZN( u2_u13_u4_n139 ) , .C1( u2_u13_u4_n182 ) );
  OAI22_X1 u2_u13_u4_U14 (.B2( u2_u13_u4_n135 ) , .ZN( u2_u13_u4_n137 ) , .B1( u2_u13_u4_n153 ) , .A1( u2_u13_u4_n155 ) , .A2( u2_u13_u4_n171 ) );
  AND3_X1 u2_u13_u4_U15 (.A2( u2_u13_u4_n134 ) , .ZN( u2_u13_u4_n135 ) , .A3( u2_u13_u4_n145 ) , .A1( u2_u13_u4_n157 ) );
  NAND2_X1 u2_u13_u4_U16 (.ZN( u2_u13_u4_n132 ) , .A2( u2_u13_u4_n170 ) , .A1( u2_u13_u4_n173 ) );
  AOI21_X1 u2_u13_u4_U17 (.B2( u2_u13_u4_n160 ) , .B1( u2_u13_u4_n161 ) , .ZN( u2_u13_u4_n162 ) , .A( u2_u13_u4_n170 ) );
  AOI21_X1 u2_u13_u4_U18 (.ZN( u2_u13_u4_n107 ) , .B2( u2_u13_u4_n143 ) , .A( u2_u13_u4_n174 ) , .B1( u2_u13_u4_n184 ) );
  AOI21_X1 u2_u13_u4_U19 (.B2( u2_u13_u4_n158 ) , .B1( u2_u13_u4_n159 ) , .ZN( u2_u13_u4_n163 ) , .A( u2_u13_u4_n174 ) );
  AOI21_X1 u2_u13_u4_U20 (.A( u2_u13_u4_n153 ) , .B2( u2_u13_u4_n154 ) , .B1( u2_u13_u4_n155 ) , .ZN( u2_u13_u4_n165 ) );
  AOI21_X1 u2_u13_u4_U21 (.A( u2_u13_u4_n156 ) , .B2( u2_u13_u4_n157 ) , .ZN( u2_u13_u4_n164 ) , .B1( u2_u13_u4_n184 ) );
  INV_X1 u2_u13_u4_U22 (.A( u2_u13_u4_n138 ) , .ZN( u2_u13_u4_n170 ) );
  AND2_X1 u2_u13_u4_U23 (.A2( u2_u13_u4_n120 ) , .ZN( u2_u13_u4_n155 ) , .A1( u2_u13_u4_n160 ) );
  INV_X1 u2_u13_u4_U24 (.A( u2_u13_u4_n156 ) , .ZN( u2_u13_u4_n175 ) );
  NAND2_X1 u2_u13_u4_U25 (.A2( u2_u13_u4_n118 ) , .ZN( u2_u13_u4_n131 ) , .A1( u2_u13_u4_n147 ) );
  NAND2_X1 u2_u13_u4_U26 (.A1( u2_u13_u4_n119 ) , .A2( u2_u13_u4_n120 ) , .ZN( u2_u13_u4_n130 ) );
  NAND2_X1 u2_u13_u4_U27 (.ZN( u2_u13_u4_n117 ) , .A2( u2_u13_u4_n118 ) , .A1( u2_u13_u4_n148 ) );
  NAND2_X1 u2_u13_u4_U28 (.ZN( u2_u13_u4_n129 ) , .A1( u2_u13_u4_n134 ) , .A2( u2_u13_u4_n148 ) );
  AND3_X1 u2_u13_u4_U29 (.A1( u2_u13_u4_n119 ) , .A2( u2_u13_u4_n143 ) , .A3( u2_u13_u4_n154 ) , .ZN( u2_u13_u4_n161 ) );
  NOR2_X1 u2_u13_u4_U3 (.ZN( u2_u13_u4_n121 ) , .A1( u2_u13_u4_n181 ) , .A2( u2_u13_u4_n182 ) );
  AND2_X1 u2_u13_u4_U30 (.A1( u2_u13_u4_n145 ) , .A2( u2_u13_u4_n147 ) , .ZN( u2_u13_u4_n159 ) );
  OR3_X1 u2_u13_u4_U31 (.A3( u2_u13_u4_n114 ) , .A2( u2_u13_u4_n115 ) , .A1( u2_u13_u4_n116 ) , .ZN( u2_u13_u4_n136 ) );
  AOI21_X1 u2_u13_u4_U32 (.A( u2_u13_u4_n113 ) , .ZN( u2_u13_u4_n116 ) , .B2( u2_u13_u4_n173 ) , .B1( u2_u13_u4_n174 ) );
  AOI21_X1 u2_u13_u4_U33 (.ZN( u2_u13_u4_n115 ) , .B2( u2_u13_u4_n145 ) , .B1( u2_u13_u4_n146 ) , .A( u2_u13_u4_n156 ) );
  OAI22_X1 u2_u13_u4_U34 (.ZN( u2_u13_u4_n114 ) , .A2( u2_u13_u4_n121 ) , .B1( u2_u13_u4_n160 ) , .B2( u2_u13_u4_n170 ) , .A1( u2_u13_u4_n171 ) );
  INV_X1 u2_u13_u4_U35 (.A( u2_u13_u4_n158 ) , .ZN( u2_u13_u4_n182 ) );
  INV_X1 u2_u13_u4_U36 (.ZN( u2_u13_u4_n181 ) , .A( u2_u13_u4_n96 ) );
  INV_X1 u2_u13_u4_U37 (.A( u2_u13_u4_n144 ) , .ZN( u2_u13_u4_n179 ) );
  INV_X1 u2_u13_u4_U38 (.A( u2_u13_u4_n157 ) , .ZN( u2_u13_u4_n178 ) );
  NAND2_X1 u2_u13_u4_U39 (.A2( u2_u13_u4_n154 ) , .A1( u2_u13_u4_n96 ) , .ZN( u2_u13_u4_n97 ) );
  INV_X1 u2_u13_u4_U4 (.A( u2_u13_u4_n117 ) , .ZN( u2_u13_u4_n184 ) );
  INV_X1 u2_u13_u4_U40 (.A( u2_u13_u4_n143 ) , .ZN( u2_u13_u4_n183 ) );
  NOR2_X1 u2_u13_u4_U41 (.ZN( u2_u13_u4_n138 ) , .A1( u2_u13_u4_n168 ) , .A2( u2_u13_u4_n169 ) );
  NOR2_X1 u2_u13_u4_U42 (.A1( u2_u13_u4_n150 ) , .A2( u2_u13_u4_n152 ) , .ZN( u2_u13_u4_n153 ) );
  NOR2_X1 u2_u13_u4_U43 (.A2( u2_u13_u4_n128 ) , .A1( u2_u13_u4_n138 ) , .ZN( u2_u13_u4_n156 ) );
  AOI22_X1 u2_u13_u4_U44 (.B2( u2_u13_u4_n122 ) , .A1( u2_u13_u4_n123 ) , .ZN( u2_u13_u4_n124 ) , .B1( u2_u13_u4_n128 ) , .A2( u2_u13_u4_n172 ) );
  NAND2_X1 u2_u13_u4_U45 (.A2( u2_u13_u4_n120 ) , .ZN( u2_u13_u4_n123 ) , .A1( u2_u13_u4_n161 ) );
  INV_X1 u2_u13_u4_U46 (.A( u2_u13_u4_n153 ) , .ZN( u2_u13_u4_n172 ) );
  AOI22_X1 u2_u13_u4_U47 (.B2( u2_u13_u4_n132 ) , .A2( u2_u13_u4_n133 ) , .ZN( u2_u13_u4_n140 ) , .A1( u2_u13_u4_n150 ) , .B1( u2_u13_u4_n179 ) );
  NAND2_X1 u2_u13_u4_U48 (.ZN( u2_u13_u4_n133 ) , .A2( u2_u13_u4_n146 ) , .A1( u2_u13_u4_n154 ) );
  NAND2_X1 u2_u13_u4_U49 (.A1( u2_u13_u4_n103 ) , .ZN( u2_u13_u4_n154 ) , .A2( u2_u13_u4_n98 ) );
  INV_X1 u2_u13_u4_U5 (.ZN( u2_u13_u4_n186 ) , .A( u2_u13_u4_n95 ) );
  NAND2_X1 u2_u13_u4_U50 (.A1( u2_u13_u4_n101 ) , .ZN( u2_u13_u4_n158 ) , .A2( u2_u13_u4_n99 ) );
  AOI21_X1 u2_u13_u4_U51 (.ZN( u2_u13_u4_n127 ) , .A( u2_u13_u4_n136 ) , .B2( u2_u13_u4_n150 ) , .B1( u2_u13_u4_n180 ) );
  INV_X1 u2_u13_u4_U52 (.A( u2_u13_u4_n160 ) , .ZN( u2_u13_u4_n180 ) );
  NAND2_X1 u2_u13_u4_U53 (.A2( u2_u13_u4_n104 ) , .A1( u2_u13_u4_n105 ) , .ZN( u2_u13_u4_n146 ) );
  NAND2_X1 u2_u13_u4_U54 (.A2( u2_u13_u4_n101 ) , .A1( u2_u13_u4_n102 ) , .ZN( u2_u13_u4_n160 ) );
  NAND2_X1 u2_u13_u4_U55 (.ZN( u2_u13_u4_n134 ) , .A1( u2_u13_u4_n98 ) , .A2( u2_u13_u4_n99 ) );
  NAND2_X1 u2_u13_u4_U56 (.A1( u2_u13_u4_n103 ) , .A2( u2_u13_u4_n104 ) , .ZN( u2_u13_u4_n143 ) );
  NAND2_X1 u2_u13_u4_U57 (.A2( u2_u13_u4_n105 ) , .ZN( u2_u13_u4_n145 ) , .A1( u2_u13_u4_n98 ) );
  NAND2_X1 u2_u13_u4_U58 (.A1( u2_u13_u4_n100 ) , .A2( u2_u13_u4_n105 ) , .ZN( u2_u13_u4_n120 ) );
  NAND2_X1 u2_u13_u4_U59 (.A1( u2_u13_u4_n102 ) , .A2( u2_u13_u4_n104 ) , .ZN( u2_u13_u4_n148 ) );
  OAI221_X1 u2_u13_u4_U6 (.C1( u2_u13_u4_n134 ) , .B1( u2_u13_u4_n158 ) , .B2( u2_u13_u4_n171 ) , .C2( u2_u13_u4_n173 ) , .A( u2_u13_u4_n94 ) , .ZN( u2_u13_u4_n95 ) );
  NAND2_X1 u2_u13_u4_U60 (.A2( u2_u13_u4_n100 ) , .A1( u2_u13_u4_n103 ) , .ZN( u2_u13_u4_n157 ) );
  INV_X1 u2_u13_u4_U61 (.A( u2_u13_u4_n150 ) , .ZN( u2_u13_u4_n173 ) );
  INV_X1 u2_u13_u4_U62 (.A( u2_u13_u4_n152 ) , .ZN( u2_u13_u4_n171 ) );
  NAND2_X1 u2_u13_u4_U63 (.A1( u2_u13_u4_n100 ) , .ZN( u2_u13_u4_n118 ) , .A2( u2_u13_u4_n99 ) );
  NAND2_X1 u2_u13_u4_U64 (.A2( u2_u13_u4_n100 ) , .A1( u2_u13_u4_n102 ) , .ZN( u2_u13_u4_n144 ) );
  NAND2_X1 u2_u13_u4_U65 (.A2( u2_u13_u4_n101 ) , .A1( u2_u13_u4_n105 ) , .ZN( u2_u13_u4_n96 ) );
  INV_X1 u2_u13_u4_U66 (.A( u2_u13_u4_n128 ) , .ZN( u2_u13_u4_n174 ) );
  NAND2_X1 u2_u13_u4_U67 (.A2( u2_u13_u4_n102 ) , .ZN( u2_u13_u4_n119 ) , .A1( u2_u13_u4_n98 ) );
  NAND2_X1 u2_u13_u4_U68 (.A2( u2_u13_u4_n101 ) , .A1( u2_u13_u4_n103 ) , .ZN( u2_u13_u4_n147 ) );
  NAND2_X1 u2_u13_u4_U69 (.A2( u2_u13_u4_n104 ) , .ZN( u2_u13_u4_n113 ) , .A1( u2_u13_u4_n99 ) );
  AOI222_X1 u2_u13_u4_U7 (.B2( u2_u13_u4_n132 ) , .A1( u2_u13_u4_n138 ) , .C2( u2_u13_u4_n175 ) , .A2( u2_u13_u4_n179 ) , .C1( u2_u13_u4_n181 ) , .B1( u2_u13_u4_n185 ) , .ZN( u2_u13_u4_n94 ) );
  NOR2_X1 u2_u13_u4_U70 (.A2( u2_u13_X_28 ) , .ZN( u2_u13_u4_n150 ) , .A1( u2_u13_u4_n168 ) );
  NOR2_X1 u2_u13_u4_U71 (.A2( u2_u13_X_29 ) , .ZN( u2_u13_u4_n152 ) , .A1( u2_u13_u4_n169 ) );
  NOR2_X1 u2_u13_u4_U72 (.A2( u2_u13_X_30 ) , .ZN( u2_u13_u4_n105 ) , .A1( u2_u13_u4_n176 ) );
  NOR2_X1 u2_u13_u4_U73 (.A2( u2_u13_X_26 ) , .ZN( u2_u13_u4_n100 ) , .A1( u2_u13_u4_n177 ) );
  NOR2_X1 u2_u13_u4_U74 (.A2( u2_u13_X_28 ) , .A1( u2_u13_X_29 ) , .ZN( u2_u13_u4_n128 ) );
  NOR2_X1 u2_u13_u4_U75 (.A2( u2_u13_X_27 ) , .A1( u2_u13_X_30 ) , .ZN( u2_u13_u4_n102 ) );
  NOR2_X1 u2_u13_u4_U76 (.A2( u2_u13_X_25 ) , .A1( u2_u13_X_26 ) , .ZN( u2_u13_u4_n98 ) );
  AND2_X1 u2_u13_u4_U77 (.A2( u2_u13_X_25 ) , .A1( u2_u13_X_26 ) , .ZN( u2_u13_u4_n104 ) );
  AND2_X1 u2_u13_u4_U78 (.A1( u2_u13_X_30 ) , .A2( u2_u13_u4_n176 ) , .ZN( u2_u13_u4_n99 ) );
  AND2_X1 u2_u13_u4_U79 (.A1( u2_u13_X_26 ) , .ZN( u2_u13_u4_n101 ) , .A2( u2_u13_u4_n177 ) );
  INV_X1 u2_u13_u4_U8 (.A( u2_u13_u4_n113 ) , .ZN( u2_u13_u4_n185 ) );
  AND2_X1 u2_u13_u4_U80 (.A1( u2_u13_X_27 ) , .A2( u2_u13_X_30 ) , .ZN( u2_u13_u4_n103 ) );
  INV_X1 u2_u13_u4_U81 (.A( u2_u13_X_28 ) , .ZN( u2_u13_u4_n169 ) );
  INV_X1 u2_u13_u4_U82 (.A( u2_u13_X_29 ) , .ZN( u2_u13_u4_n168 ) );
  INV_X1 u2_u13_u4_U83 (.A( u2_u13_X_25 ) , .ZN( u2_u13_u4_n177 ) );
  INV_X1 u2_u13_u4_U84 (.A( u2_u13_X_27 ) , .ZN( u2_u13_u4_n176 ) );
  NAND4_X1 u2_u13_u4_U85 (.ZN( u2_out13_25 ) , .A4( u2_u13_u4_n139 ) , .A3( u2_u13_u4_n140 ) , .A2( u2_u13_u4_n141 ) , .A1( u2_u13_u4_n142 ) );
  OAI21_X1 u2_u13_u4_U86 (.A( u2_u13_u4_n128 ) , .B2( u2_u13_u4_n129 ) , .B1( u2_u13_u4_n130 ) , .ZN( u2_u13_u4_n142 ) );
  OAI21_X1 u2_u13_u4_U87 (.B2( u2_u13_u4_n131 ) , .ZN( u2_u13_u4_n141 ) , .A( u2_u13_u4_n175 ) , .B1( u2_u13_u4_n183 ) );
  NAND4_X1 u2_u13_u4_U88 (.ZN( u2_out13_14 ) , .A4( u2_u13_u4_n124 ) , .A3( u2_u13_u4_n125 ) , .A2( u2_u13_u4_n126 ) , .A1( u2_u13_u4_n127 ) );
  AOI22_X1 u2_u13_u4_U89 (.B2( u2_u13_u4_n117 ) , .ZN( u2_u13_u4_n126 ) , .A1( u2_u13_u4_n129 ) , .B1( u2_u13_u4_n152 ) , .A2( u2_u13_u4_n175 ) );
  NOR4_X1 u2_u13_u4_U9 (.A4( u2_u13_u4_n106 ) , .A3( u2_u13_u4_n107 ) , .A2( u2_u13_u4_n108 ) , .A1( u2_u13_u4_n109 ) , .ZN( u2_u13_u4_n110 ) );
  AOI22_X1 u2_u13_u4_U90 (.ZN( u2_u13_u4_n125 ) , .B2( u2_u13_u4_n131 ) , .A2( u2_u13_u4_n132 ) , .B1( u2_u13_u4_n138 ) , .A1( u2_u13_u4_n178 ) );
  NAND4_X1 u2_u13_u4_U91 (.ZN( u2_out13_8 ) , .A4( u2_u13_u4_n110 ) , .A3( u2_u13_u4_n111 ) , .A2( u2_u13_u4_n112 ) , .A1( u2_u13_u4_n186 ) );
  NAND2_X1 u2_u13_u4_U92 (.ZN( u2_u13_u4_n112 ) , .A2( u2_u13_u4_n130 ) , .A1( u2_u13_u4_n150 ) );
  AOI22_X1 u2_u13_u4_U93 (.ZN( u2_u13_u4_n111 ) , .B2( u2_u13_u4_n132 ) , .A1( u2_u13_u4_n152 ) , .B1( u2_u13_u4_n178 ) , .A2( u2_u13_u4_n97 ) );
  AOI22_X1 u2_u13_u4_U94 (.B2( u2_u13_u4_n149 ) , .B1( u2_u13_u4_n150 ) , .A2( u2_u13_u4_n151 ) , .A1( u2_u13_u4_n152 ) , .ZN( u2_u13_u4_n167 ) );
  NOR4_X1 u2_u13_u4_U95 (.A4( u2_u13_u4_n162 ) , .A3( u2_u13_u4_n163 ) , .A2( u2_u13_u4_n164 ) , .A1( u2_u13_u4_n165 ) , .ZN( u2_u13_u4_n166 ) );
  NAND3_X1 u2_u13_u4_U96 (.ZN( u2_out13_3 ) , .A3( u2_u13_u4_n166 ) , .A1( u2_u13_u4_n167 ) , .A2( u2_u13_u4_n186 ) );
  NAND3_X1 u2_u13_u4_U97 (.A3( u2_u13_u4_n146 ) , .A2( u2_u13_u4_n147 ) , .A1( u2_u13_u4_n148 ) , .ZN( u2_u13_u4_n149 ) );
  NAND3_X1 u2_u13_u4_U98 (.A3( u2_u13_u4_n143 ) , .A2( u2_u13_u4_n144 ) , .A1( u2_u13_u4_n145 ) , .ZN( u2_u13_u4_n151 ) );
  NAND3_X1 u2_u13_u4_U99 (.A3( u2_u13_u4_n121 ) , .ZN( u2_u13_u4_n122 ) , .A2( u2_u13_u4_n144 ) , .A1( u2_u13_u4_n154 ) );
  INV_X1 u2_u13_u5_U10 (.A( u2_u13_u5_n121 ) , .ZN( u2_u13_u5_n177 ) );
  NOR3_X1 u2_u13_u5_U100 (.A3( u2_u13_u5_n141 ) , .A1( u2_u13_u5_n142 ) , .ZN( u2_u13_u5_n143 ) , .A2( u2_u13_u5_n191 ) );
  NAND4_X1 u2_u13_u5_U101 (.ZN( u2_out13_4 ) , .A4( u2_u13_u5_n112 ) , .A2( u2_u13_u5_n113 ) , .A1( u2_u13_u5_n114 ) , .A3( u2_u13_u5_n195 ) );
  AOI211_X1 u2_u13_u5_U102 (.A( u2_u13_u5_n110 ) , .C1( u2_u13_u5_n111 ) , .ZN( u2_u13_u5_n112 ) , .B( u2_u13_u5_n118 ) , .C2( u2_u13_u5_n177 ) );
  AOI222_X1 u2_u13_u5_U103 (.ZN( u2_u13_u5_n113 ) , .A1( u2_u13_u5_n131 ) , .C1( u2_u13_u5_n148 ) , .B2( u2_u13_u5_n174 ) , .C2( u2_u13_u5_n178 ) , .A2( u2_u13_u5_n179 ) , .B1( u2_u13_u5_n99 ) );
  NAND3_X1 u2_u13_u5_U104 (.A2( u2_u13_u5_n154 ) , .A3( u2_u13_u5_n158 ) , .A1( u2_u13_u5_n161 ) , .ZN( u2_u13_u5_n99 ) );
  NOR2_X1 u2_u13_u5_U11 (.ZN( u2_u13_u5_n160 ) , .A2( u2_u13_u5_n173 ) , .A1( u2_u13_u5_n177 ) );
  INV_X1 u2_u13_u5_U12 (.A( u2_u13_u5_n150 ) , .ZN( u2_u13_u5_n174 ) );
  AOI21_X1 u2_u13_u5_U13 (.A( u2_u13_u5_n160 ) , .B2( u2_u13_u5_n161 ) , .ZN( u2_u13_u5_n162 ) , .B1( u2_u13_u5_n192 ) );
  INV_X1 u2_u13_u5_U14 (.A( u2_u13_u5_n159 ) , .ZN( u2_u13_u5_n192 ) );
  AOI21_X1 u2_u13_u5_U15 (.A( u2_u13_u5_n156 ) , .B2( u2_u13_u5_n157 ) , .B1( u2_u13_u5_n158 ) , .ZN( u2_u13_u5_n163 ) );
  AOI21_X1 u2_u13_u5_U16 (.B2( u2_u13_u5_n139 ) , .B1( u2_u13_u5_n140 ) , .ZN( u2_u13_u5_n141 ) , .A( u2_u13_u5_n150 ) );
  OAI21_X1 u2_u13_u5_U17 (.A( u2_u13_u5_n133 ) , .B2( u2_u13_u5_n134 ) , .B1( u2_u13_u5_n135 ) , .ZN( u2_u13_u5_n142 ) );
  OAI21_X1 u2_u13_u5_U18 (.ZN( u2_u13_u5_n133 ) , .B2( u2_u13_u5_n147 ) , .A( u2_u13_u5_n173 ) , .B1( u2_u13_u5_n188 ) );
  NAND2_X1 u2_u13_u5_U19 (.A2( u2_u13_u5_n119 ) , .A1( u2_u13_u5_n123 ) , .ZN( u2_u13_u5_n137 ) );
  INV_X1 u2_u13_u5_U20 (.A( u2_u13_u5_n155 ) , .ZN( u2_u13_u5_n194 ) );
  NAND2_X1 u2_u13_u5_U21 (.A1( u2_u13_u5_n121 ) , .ZN( u2_u13_u5_n132 ) , .A2( u2_u13_u5_n172 ) );
  NAND2_X1 u2_u13_u5_U22 (.A2( u2_u13_u5_n122 ) , .ZN( u2_u13_u5_n136 ) , .A1( u2_u13_u5_n154 ) );
  NAND2_X1 u2_u13_u5_U23 (.A2( u2_u13_u5_n119 ) , .A1( u2_u13_u5_n120 ) , .ZN( u2_u13_u5_n159 ) );
  INV_X1 u2_u13_u5_U24 (.A( u2_u13_u5_n156 ) , .ZN( u2_u13_u5_n175 ) );
  INV_X1 u2_u13_u5_U25 (.A( u2_u13_u5_n158 ) , .ZN( u2_u13_u5_n188 ) );
  INV_X1 u2_u13_u5_U26 (.A( u2_u13_u5_n152 ) , .ZN( u2_u13_u5_n179 ) );
  INV_X1 u2_u13_u5_U27 (.A( u2_u13_u5_n140 ) , .ZN( u2_u13_u5_n182 ) );
  INV_X1 u2_u13_u5_U28 (.A( u2_u13_u5_n151 ) , .ZN( u2_u13_u5_n183 ) );
  INV_X1 u2_u13_u5_U29 (.A( u2_u13_u5_n123 ) , .ZN( u2_u13_u5_n185 ) );
  NOR2_X1 u2_u13_u5_U3 (.ZN( u2_u13_u5_n134 ) , .A1( u2_u13_u5_n183 ) , .A2( u2_u13_u5_n190 ) );
  INV_X1 u2_u13_u5_U30 (.A( u2_u13_u5_n161 ) , .ZN( u2_u13_u5_n184 ) );
  INV_X1 u2_u13_u5_U31 (.A( u2_u13_u5_n139 ) , .ZN( u2_u13_u5_n189 ) );
  INV_X1 u2_u13_u5_U32 (.A( u2_u13_u5_n157 ) , .ZN( u2_u13_u5_n190 ) );
  INV_X1 u2_u13_u5_U33 (.A( u2_u13_u5_n120 ) , .ZN( u2_u13_u5_n193 ) );
  NAND2_X1 u2_u13_u5_U34 (.ZN( u2_u13_u5_n111 ) , .A1( u2_u13_u5_n140 ) , .A2( u2_u13_u5_n155 ) );
  NOR2_X1 u2_u13_u5_U35 (.ZN( u2_u13_u5_n100 ) , .A1( u2_u13_u5_n170 ) , .A2( u2_u13_u5_n180 ) );
  INV_X1 u2_u13_u5_U36 (.A( u2_u13_u5_n117 ) , .ZN( u2_u13_u5_n196 ) );
  OAI221_X1 u2_u13_u5_U37 (.A( u2_u13_u5_n116 ) , .ZN( u2_u13_u5_n117 ) , .B2( u2_u13_u5_n119 ) , .C1( u2_u13_u5_n153 ) , .C2( u2_u13_u5_n158 ) , .B1( u2_u13_u5_n172 ) );
  AOI222_X1 u2_u13_u5_U38 (.ZN( u2_u13_u5_n116 ) , .B2( u2_u13_u5_n145 ) , .C1( u2_u13_u5_n148 ) , .A2( u2_u13_u5_n174 ) , .C2( u2_u13_u5_n177 ) , .B1( u2_u13_u5_n187 ) , .A1( u2_u13_u5_n193 ) );
  INV_X1 u2_u13_u5_U39 (.A( u2_u13_u5_n115 ) , .ZN( u2_u13_u5_n187 ) );
  INV_X1 u2_u13_u5_U4 (.A( u2_u13_u5_n138 ) , .ZN( u2_u13_u5_n191 ) );
  AOI22_X1 u2_u13_u5_U40 (.B2( u2_u13_u5_n131 ) , .A2( u2_u13_u5_n146 ) , .ZN( u2_u13_u5_n169 ) , .B1( u2_u13_u5_n174 ) , .A1( u2_u13_u5_n185 ) );
  NOR2_X1 u2_u13_u5_U41 (.A1( u2_u13_u5_n146 ) , .ZN( u2_u13_u5_n150 ) , .A2( u2_u13_u5_n173 ) );
  AOI21_X1 u2_u13_u5_U42 (.A( u2_u13_u5_n118 ) , .B2( u2_u13_u5_n145 ) , .ZN( u2_u13_u5_n168 ) , .B1( u2_u13_u5_n186 ) );
  INV_X1 u2_u13_u5_U43 (.A( u2_u13_u5_n122 ) , .ZN( u2_u13_u5_n186 ) );
  NOR2_X1 u2_u13_u5_U44 (.A1( u2_u13_u5_n146 ) , .ZN( u2_u13_u5_n152 ) , .A2( u2_u13_u5_n176 ) );
  NOR2_X1 u2_u13_u5_U45 (.A1( u2_u13_u5_n115 ) , .ZN( u2_u13_u5_n118 ) , .A2( u2_u13_u5_n153 ) );
  NOR2_X1 u2_u13_u5_U46 (.A2( u2_u13_u5_n145 ) , .ZN( u2_u13_u5_n156 ) , .A1( u2_u13_u5_n174 ) );
  NOR2_X1 u2_u13_u5_U47 (.ZN( u2_u13_u5_n121 ) , .A2( u2_u13_u5_n145 ) , .A1( u2_u13_u5_n176 ) );
  AOI22_X1 u2_u13_u5_U48 (.ZN( u2_u13_u5_n114 ) , .A2( u2_u13_u5_n137 ) , .A1( u2_u13_u5_n145 ) , .B2( u2_u13_u5_n175 ) , .B1( u2_u13_u5_n193 ) );
  OAI211_X1 u2_u13_u5_U49 (.B( u2_u13_u5_n124 ) , .A( u2_u13_u5_n125 ) , .C2( u2_u13_u5_n126 ) , .C1( u2_u13_u5_n127 ) , .ZN( u2_u13_u5_n128 ) );
  OAI21_X1 u2_u13_u5_U5 (.B2( u2_u13_u5_n136 ) , .B1( u2_u13_u5_n137 ) , .ZN( u2_u13_u5_n138 ) , .A( u2_u13_u5_n177 ) );
  NOR3_X1 u2_u13_u5_U50 (.ZN( u2_u13_u5_n127 ) , .A1( u2_u13_u5_n136 ) , .A3( u2_u13_u5_n148 ) , .A2( u2_u13_u5_n182 ) );
  OAI21_X1 u2_u13_u5_U51 (.ZN( u2_u13_u5_n124 ) , .A( u2_u13_u5_n177 ) , .B2( u2_u13_u5_n183 ) , .B1( u2_u13_u5_n189 ) );
  OAI21_X1 u2_u13_u5_U52 (.ZN( u2_u13_u5_n125 ) , .A( u2_u13_u5_n174 ) , .B2( u2_u13_u5_n185 ) , .B1( u2_u13_u5_n190 ) );
  AOI21_X1 u2_u13_u5_U53 (.A( u2_u13_u5_n153 ) , .B2( u2_u13_u5_n154 ) , .B1( u2_u13_u5_n155 ) , .ZN( u2_u13_u5_n164 ) );
  AOI21_X1 u2_u13_u5_U54 (.ZN( u2_u13_u5_n110 ) , .B1( u2_u13_u5_n122 ) , .B2( u2_u13_u5_n139 ) , .A( u2_u13_u5_n153 ) );
  INV_X1 u2_u13_u5_U55 (.A( u2_u13_u5_n153 ) , .ZN( u2_u13_u5_n176 ) );
  INV_X1 u2_u13_u5_U56 (.A( u2_u13_u5_n126 ) , .ZN( u2_u13_u5_n173 ) );
  AND2_X1 u2_u13_u5_U57 (.A2( u2_u13_u5_n104 ) , .A1( u2_u13_u5_n107 ) , .ZN( u2_u13_u5_n147 ) );
  AND2_X1 u2_u13_u5_U58 (.A2( u2_u13_u5_n104 ) , .A1( u2_u13_u5_n108 ) , .ZN( u2_u13_u5_n148 ) );
  NAND2_X1 u2_u13_u5_U59 (.A1( u2_u13_u5_n105 ) , .A2( u2_u13_u5_n106 ) , .ZN( u2_u13_u5_n158 ) );
  INV_X1 u2_u13_u5_U6 (.A( u2_u13_u5_n135 ) , .ZN( u2_u13_u5_n178 ) );
  NAND2_X1 u2_u13_u5_U60 (.A2( u2_u13_u5_n108 ) , .A1( u2_u13_u5_n109 ) , .ZN( u2_u13_u5_n139 ) );
  NAND2_X1 u2_u13_u5_U61 (.A1( u2_u13_u5_n106 ) , .A2( u2_u13_u5_n108 ) , .ZN( u2_u13_u5_n119 ) );
  NAND2_X1 u2_u13_u5_U62 (.A2( u2_u13_u5_n103 ) , .A1( u2_u13_u5_n105 ) , .ZN( u2_u13_u5_n140 ) );
  NAND2_X1 u2_u13_u5_U63 (.A2( u2_u13_u5_n104 ) , .A1( u2_u13_u5_n105 ) , .ZN( u2_u13_u5_n155 ) );
  NAND2_X1 u2_u13_u5_U64 (.A2( u2_u13_u5_n106 ) , .A1( u2_u13_u5_n107 ) , .ZN( u2_u13_u5_n122 ) );
  NAND2_X1 u2_u13_u5_U65 (.A2( u2_u13_u5_n100 ) , .A1( u2_u13_u5_n106 ) , .ZN( u2_u13_u5_n115 ) );
  NAND2_X1 u2_u13_u5_U66 (.A2( u2_u13_u5_n100 ) , .A1( u2_u13_u5_n103 ) , .ZN( u2_u13_u5_n161 ) );
  NAND2_X1 u2_u13_u5_U67 (.A1( u2_u13_u5_n105 ) , .A2( u2_u13_u5_n109 ) , .ZN( u2_u13_u5_n154 ) );
  INV_X1 u2_u13_u5_U68 (.A( u2_u13_u5_n146 ) , .ZN( u2_u13_u5_n172 ) );
  NAND2_X1 u2_u13_u5_U69 (.A1( u2_u13_u5_n103 ) , .A2( u2_u13_u5_n108 ) , .ZN( u2_u13_u5_n123 ) );
  OAI22_X1 u2_u13_u5_U7 (.B2( u2_u13_u5_n149 ) , .B1( u2_u13_u5_n150 ) , .A2( u2_u13_u5_n151 ) , .A1( u2_u13_u5_n152 ) , .ZN( u2_u13_u5_n165 ) );
  NAND2_X1 u2_u13_u5_U70 (.A2( u2_u13_u5_n103 ) , .A1( u2_u13_u5_n107 ) , .ZN( u2_u13_u5_n151 ) );
  NAND2_X1 u2_u13_u5_U71 (.A2( u2_u13_u5_n107 ) , .A1( u2_u13_u5_n109 ) , .ZN( u2_u13_u5_n120 ) );
  NAND2_X1 u2_u13_u5_U72 (.A2( u2_u13_u5_n100 ) , .A1( u2_u13_u5_n109 ) , .ZN( u2_u13_u5_n157 ) );
  AND2_X1 u2_u13_u5_U73 (.A2( u2_u13_u5_n100 ) , .A1( u2_u13_u5_n104 ) , .ZN( u2_u13_u5_n131 ) );
  INV_X1 u2_u13_u5_U74 (.A( u2_u13_u5_n102 ) , .ZN( u2_u13_u5_n195 ) );
  OAI221_X1 u2_u13_u5_U75 (.A( u2_u13_u5_n101 ) , .ZN( u2_u13_u5_n102 ) , .C2( u2_u13_u5_n115 ) , .C1( u2_u13_u5_n126 ) , .B1( u2_u13_u5_n134 ) , .B2( u2_u13_u5_n160 ) );
  OAI21_X1 u2_u13_u5_U76 (.ZN( u2_u13_u5_n101 ) , .B1( u2_u13_u5_n137 ) , .A( u2_u13_u5_n146 ) , .B2( u2_u13_u5_n147 ) );
  NOR2_X1 u2_u13_u5_U77 (.A2( u2_u13_X_34 ) , .A1( u2_u13_X_35 ) , .ZN( u2_u13_u5_n145 ) );
  NOR2_X1 u2_u13_u5_U78 (.A2( u2_u13_X_34 ) , .ZN( u2_u13_u5_n146 ) , .A1( u2_u13_u5_n171 ) );
  NOR2_X1 u2_u13_u5_U79 (.A2( u2_u13_X_31 ) , .A1( u2_u13_X_32 ) , .ZN( u2_u13_u5_n103 ) );
  NOR3_X1 u2_u13_u5_U8 (.A2( u2_u13_u5_n147 ) , .A1( u2_u13_u5_n148 ) , .ZN( u2_u13_u5_n149 ) , .A3( u2_u13_u5_n194 ) );
  NOR2_X1 u2_u13_u5_U80 (.A2( u2_u13_X_36 ) , .ZN( u2_u13_u5_n105 ) , .A1( u2_u13_u5_n180 ) );
  NOR2_X1 u2_u13_u5_U81 (.A2( u2_u13_X_33 ) , .ZN( u2_u13_u5_n108 ) , .A1( u2_u13_u5_n170 ) );
  NOR2_X1 u2_u13_u5_U82 (.A2( u2_u13_X_33 ) , .A1( u2_u13_X_36 ) , .ZN( u2_u13_u5_n107 ) );
  NOR2_X1 u2_u13_u5_U83 (.A2( u2_u13_X_31 ) , .ZN( u2_u13_u5_n104 ) , .A1( u2_u13_u5_n181 ) );
  NAND2_X1 u2_u13_u5_U84 (.A2( u2_u13_X_34 ) , .A1( u2_u13_X_35 ) , .ZN( u2_u13_u5_n153 ) );
  NAND2_X1 u2_u13_u5_U85 (.A1( u2_u13_X_34 ) , .ZN( u2_u13_u5_n126 ) , .A2( u2_u13_u5_n171 ) );
  AND2_X1 u2_u13_u5_U86 (.A1( u2_u13_X_31 ) , .A2( u2_u13_X_32 ) , .ZN( u2_u13_u5_n106 ) );
  AND2_X1 u2_u13_u5_U87 (.A1( u2_u13_X_31 ) , .ZN( u2_u13_u5_n109 ) , .A2( u2_u13_u5_n181 ) );
  INV_X1 u2_u13_u5_U88 (.A( u2_u13_X_33 ) , .ZN( u2_u13_u5_n180 ) );
  INV_X1 u2_u13_u5_U89 (.A( u2_u13_X_35 ) , .ZN( u2_u13_u5_n171 ) );
  NOR2_X1 u2_u13_u5_U9 (.ZN( u2_u13_u5_n135 ) , .A1( u2_u13_u5_n173 ) , .A2( u2_u13_u5_n176 ) );
  INV_X1 u2_u13_u5_U90 (.A( u2_u13_X_36 ) , .ZN( u2_u13_u5_n170 ) );
  INV_X1 u2_u13_u5_U91 (.A( u2_u13_X_32 ) , .ZN( u2_u13_u5_n181 ) );
  NAND4_X1 u2_u13_u5_U92 (.ZN( u2_out13_29 ) , .A4( u2_u13_u5_n129 ) , .A3( u2_u13_u5_n130 ) , .A2( u2_u13_u5_n168 ) , .A1( u2_u13_u5_n196 ) );
  AOI221_X1 u2_u13_u5_U93 (.A( u2_u13_u5_n128 ) , .ZN( u2_u13_u5_n129 ) , .C2( u2_u13_u5_n132 ) , .B2( u2_u13_u5_n159 ) , .B1( u2_u13_u5_n176 ) , .C1( u2_u13_u5_n184 ) );
  AOI222_X1 u2_u13_u5_U94 (.ZN( u2_u13_u5_n130 ) , .A2( u2_u13_u5_n146 ) , .B1( u2_u13_u5_n147 ) , .C2( u2_u13_u5_n175 ) , .B2( u2_u13_u5_n179 ) , .A1( u2_u13_u5_n188 ) , .C1( u2_u13_u5_n194 ) );
  NAND4_X1 u2_u13_u5_U95 (.ZN( u2_out13_19 ) , .A4( u2_u13_u5_n166 ) , .A3( u2_u13_u5_n167 ) , .A2( u2_u13_u5_n168 ) , .A1( u2_u13_u5_n169 ) );
  AOI22_X1 u2_u13_u5_U96 (.B2( u2_u13_u5_n145 ) , .A2( u2_u13_u5_n146 ) , .ZN( u2_u13_u5_n167 ) , .B1( u2_u13_u5_n182 ) , .A1( u2_u13_u5_n189 ) );
  NOR4_X1 u2_u13_u5_U97 (.A4( u2_u13_u5_n162 ) , .A3( u2_u13_u5_n163 ) , .A2( u2_u13_u5_n164 ) , .A1( u2_u13_u5_n165 ) , .ZN( u2_u13_u5_n166 ) );
  NAND4_X1 u2_u13_u5_U98 (.ZN( u2_out13_11 ) , .A4( u2_u13_u5_n143 ) , .A3( u2_u13_u5_n144 ) , .A2( u2_u13_u5_n169 ) , .A1( u2_u13_u5_n196 ) );
  AOI22_X1 u2_u13_u5_U99 (.A2( u2_u13_u5_n132 ) , .ZN( u2_u13_u5_n144 ) , .B2( u2_u13_u5_n145 ) , .B1( u2_u13_u5_n184 ) , .A1( u2_u13_u5_n194 ) );
  AOI22_X1 u2_u13_u6_U10 (.A2( u2_u13_u6_n151 ) , .B2( u2_u13_u6_n161 ) , .A1( u2_u13_u6_n167 ) , .B1( u2_u13_u6_n170 ) , .ZN( u2_u13_u6_n89 ) );
  AOI21_X1 u2_u13_u6_U11 (.B1( u2_u13_u6_n107 ) , .B2( u2_u13_u6_n132 ) , .A( u2_u13_u6_n158 ) , .ZN( u2_u13_u6_n88 ) );
  AOI21_X1 u2_u13_u6_U12 (.B2( u2_u13_u6_n147 ) , .B1( u2_u13_u6_n148 ) , .ZN( u2_u13_u6_n149 ) , .A( u2_u13_u6_n158 ) );
  AOI21_X1 u2_u13_u6_U13 (.ZN( u2_u13_u6_n106 ) , .A( u2_u13_u6_n142 ) , .B2( u2_u13_u6_n159 ) , .B1( u2_u13_u6_n164 ) );
  INV_X1 u2_u13_u6_U14 (.A( u2_u13_u6_n155 ) , .ZN( u2_u13_u6_n161 ) );
  INV_X1 u2_u13_u6_U15 (.A( u2_u13_u6_n128 ) , .ZN( u2_u13_u6_n164 ) );
  NAND2_X1 u2_u13_u6_U16 (.ZN( u2_u13_u6_n110 ) , .A1( u2_u13_u6_n122 ) , .A2( u2_u13_u6_n129 ) );
  NAND2_X1 u2_u13_u6_U17 (.ZN( u2_u13_u6_n124 ) , .A2( u2_u13_u6_n146 ) , .A1( u2_u13_u6_n148 ) );
  INV_X1 u2_u13_u6_U18 (.A( u2_u13_u6_n132 ) , .ZN( u2_u13_u6_n171 ) );
  AND2_X1 u2_u13_u6_U19 (.A1( u2_u13_u6_n100 ) , .ZN( u2_u13_u6_n130 ) , .A2( u2_u13_u6_n147 ) );
  INV_X1 u2_u13_u6_U20 (.A( u2_u13_u6_n127 ) , .ZN( u2_u13_u6_n173 ) );
  INV_X1 u2_u13_u6_U21 (.A( u2_u13_u6_n121 ) , .ZN( u2_u13_u6_n167 ) );
  INV_X1 u2_u13_u6_U22 (.A( u2_u13_u6_n100 ) , .ZN( u2_u13_u6_n169 ) );
  INV_X1 u2_u13_u6_U23 (.A( u2_u13_u6_n123 ) , .ZN( u2_u13_u6_n170 ) );
  INV_X1 u2_u13_u6_U24 (.A( u2_u13_u6_n113 ) , .ZN( u2_u13_u6_n168 ) );
  AND2_X1 u2_u13_u6_U25 (.A1( u2_u13_u6_n107 ) , .A2( u2_u13_u6_n119 ) , .ZN( u2_u13_u6_n133 ) );
  AND2_X1 u2_u13_u6_U26 (.A2( u2_u13_u6_n121 ) , .A1( u2_u13_u6_n122 ) , .ZN( u2_u13_u6_n131 ) );
  AND3_X1 u2_u13_u6_U27 (.ZN( u2_u13_u6_n120 ) , .A2( u2_u13_u6_n127 ) , .A1( u2_u13_u6_n132 ) , .A3( u2_u13_u6_n145 ) );
  INV_X1 u2_u13_u6_U28 (.A( u2_u13_u6_n146 ) , .ZN( u2_u13_u6_n163 ) );
  AOI222_X1 u2_u13_u6_U29 (.ZN( u2_u13_u6_n114 ) , .A1( u2_u13_u6_n118 ) , .A2( u2_u13_u6_n126 ) , .B2( u2_u13_u6_n151 ) , .C2( u2_u13_u6_n159 ) , .C1( u2_u13_u6_n168 ) , .B1( u2_u13_u6_n169 ) );
  INV_X1 u2_u13_u6_U3 (.A( u2_u13_u6_n110 ) , .ZN( u2_u13_u6_n166 ) );
  NOR2_X1 u2_u13_u6_U30 (.A1( u2_u13_u6_n162 ) , .A2( u2_u13_u6_n165 ) , .ZN( u2_u13_u6_n98 ) );
  AOI211_X1 u2_u13_u6_U31 (.B( u2_u13_u6_n134 ) , .A( u2_u13_u6_n135 ) , .C1( u2_u13_u6_n136 ) , .ZN( u2_u13_u6_n137 ) , .C2( u2_u13_u6_n151 ) );
  AOI21_X1 u2_u13_u6_U32 (.B2( u2_u13_u6_n132 ) , .B1( u2_u13_u6_n133 ) , .ZN( u2_u13_u6_n134 ) , .A( u2_u13_u6_n158 ) );
  AOI21_X1 u2_u13_u6_U33 (.B1( u2_u13_u6_n131 ) , .ZN( u2_u13_u6_n135 ) , .A( u2_u13_u6_n144 ) , .B2( u2_u13_u6_n146 ) );
  NAND4_X1 u2_u13_u6_U34 (.A4( u2_u13_u6_n127 ) , .A3( u2_u13_u6_n128 ) , .A2( u2_u13_u6_n129 ) , .A1( u2_u13_u6_n130 ) , .ZN( u2_u13_u6_n136 ) );
  NAND2_X1 u2_u13_u6_U35 (.A1( u2_u13_u6_n144 ) , .ZN( u2_u13_u6_n151 ) , .A2( u2_u13_u6_n158 ) );
  NAND2_X1 u2_u13_u6_U36 (.ZN( u2_u13_u6_n132 ) , .A1( u2_u13_u6_n91 ) , .A2( u2_u13_u6_n97 ) );
  AOI22_X1 u2_u13_u6_U37 (.B2( u2_u13_u6_n110 ) , .B1( u2_u13_u6_n111 ) , .A1( u2_u13_u6_n112 ) , .ZN( u2_u13_u6_n115 ) , .A2( u2_u13_u6_n161 ) );
  NAND4_X1 u2_u13_u6_U38 (.A3( u2_u13_u6_n109 ) , .ZN( u2_u13_u6_n112 ) , .A4( u2_u13_u6_n132 ) , .A2( u2_u13_u6_n147 ) , .A1( u2_u13_u6_n166 ) );
  NOR2_X1 u2_u13_u6_U39 (.ZN( u2_u13_u6_n109 ) , .A1( u2_u13_u6_n170 ) , .A2( u2_u13_u6_n173 ) );
  INV_X1 u2_u13_u6_U4 (.A( u2_u13_u6_n142 ) , .ZN( u2_u13_u6_n174 ) );
  NOR2_X1 u2_u13_u6_U40 (.A2( u2_u13_u6_n126 ) , .ZN( u2_u13_u6_n155 ) , .A1( u2_u13_u6_n160 ) );
  NAND2_X1 u2_u13_u6_U41 (.ZN( u2_u13_u6_n146 ) , .A2( u2_u13_u6_n94 ) , .A1( u2_u13_u6_n99 ) );
  AOI21_X1 u2_u13_u6_U42 (.A( u2_u13_u6_n144 ) , .B2( u2_u13_u6_n145 ) , .B1( u2_u13_u6_n146 ) , .ZN( u2_u13_u6_n150 ) );
  INV_X1 u2_u13_u6_U43 (.A( u2_u13_u6_n111 ) , .ZN( u2_u13_u6_n158 ) );
  NAND2_X1 u2_u13_u6_U44 (.ZN( u2_u13_u6_n127 ) , .A1( u2_u13_u6_n91 ) , .A2( u2_u13_u6_n92 ) );
  NAND2_X1 u2_u13_u6_U45 (.ZN( u2_u13_u6_n129 ) , .A2( u2_u13_u6_n95 ) , .A1( u2_u13_u6_n96 ) );
  INV_X1 u2_u13_u6_U46 (.A( u2_u13_u6_n144 ) , .ZN( u2_u13_u6_n159 ) );
  NAND2_X1 u2_u13_u6_U47 (.ZN( u2_u13_u6_n145 ) , .A2( u2_u13_u6_n97 ) , .A1( u2_u13_u6_n98 ) );
  NAND2_X1 u2_u13_u6_U48 (.ZN( u2_u13_u6_n148 ) , .A2( u2_u13_u6_n92 ) , .A1( u2_u13_u6_n94 ) );
  NAND2_X1 u2_u13_u6_U49 (.ZN( u2_u13_u6_n108 ) , .A2( u2_u13_u6_n139 ) , .A1( u2_u13_u6_n144 ) );
  NAND2_X1 u2_u13_u6_U5 (.A2( u2_u13_u6_n143 ) , .ZN( u2_u13_u6_n152 ) , .A1( u2_u13_u6_n166 ) );
  NAND2_X1 u2_u13_u6_U50 (.ZN( u2_u13_u6_n121 ) , .A2( u2_u13_u6_n95 ) , .A1( u2_u13_u6_n97 ) );
  NAND2_X1 u2_u13_u6_U51 (.ZN( u2_u13_u6_n107 ) , .A2( u2_u13_u6_n92 ) , .A1( u2_u13_u6_n95 ) );
  AND2_X1 u2_u13_u6_U52 (.ZN( u2_u13_u6_n118 ) , .A2( u2_u13_u6_n91 ) , .A1( u2_u13_u6_n99 ) );
  NAND2_X1 u2_u13_u6_U53 (.ZN( u2_u13_u6_n147 ) , .A2( u2_u13_u6_n98 ) , .A1( u2_u13_u6_n99 ) );
  NAND2_X1 u2_u13_u6_U54 (.ZN( u2_u13_u6_n128 ) , .A1( u2_u13_u6_n94 ) , .A2( u2_u13_u6_n96 ) );
  NAND2_X1 u2_u13_u6_U55 (.ZN( u2_u13_u6_n119 ) , .A2( u2_u13_u6_n95 ) , .A1( u2_u13_u6_n99 ) );
  NAND2_X1 u2_u13_u6_U56 (.ZN( u2_u13_u6_n123 ) , .A2( u2_u13_u6_n91 ) , .A1( u2_u13_u6_n96 ) );
  NAND2_X1 u2_u13_u6_U57 (.ZN( u2_u13_u6_n100 ) , .A2( u2_u13_u6_n92 ) , .A1( u2_u13_u6_n98 ) );
  NAND2_X1 u2_u13_u6_U58 (.ZN( u2_u13_u6_n122 ) , .A1( u2_u13_u6_n94 ) , .A2( u2_u13_u6_n97 ) );
  INV_X1 u2_u13_u6_U59 (.A( u2_u13_u6_n139 ) , .ZN( u2_u13_u6_n160 ) );
  AOI22_X1 u2_u13_u6_U6 (.B2( u2_u13_u6_n101 ) , .A1( u2_u13_u6_n102 ) , .ZN( u2_u13_u6_n103 ) , .B1( u2_u13_u6_n160 ) , .A2( u2_u13_u6_n161 ) );
  NAND2_X1 u2_u13_u6_U60 (.ZN( u2_u13_u6_n113 ) , .A1( u2_u13_u6_n96 ) , .A2( u2_u13_u6_n98 ) );
  NOR2_X1 u2_u13_u6_U61 (.A2( u2_u13_X_40 ) , .A1( u2_u13_X_41 ) , .ZN( u2_u13_u6_n126 ) );
  NOR2_X1 u2_u13_u6_U62 (.A2( u2_u13_X_39 ) , .A1( u2_u13_X_42 ) , .ZN( u2_u13_u6_n92 ) );
  NOR2_X1 u2_u13_u6_U63 (.A2( u2_u13_X_39 ) , .A1( u2_u13_u6_n156 ) , .ZN( u2_u13_u6_n97 ) );
  NOR2_X1 u2_u13_u6_U64 (.A2( u2_u13_X_38 ) , .A1( u2_u13_u6_n165 ) , .ZN( u2_u13_u6_n95 ) );
  NOR2_X1 u2_u13_u6_U65 (.A2( u2_u13_X_41 ) , .ZN( u2_u13_u6_n111 ) , .A1( u2_u13_u6_n157 ) );
  NOR2_X1 u2_u13_u6_U66 (.A2( u2_u13_X_37 ) , .A1( u2_u13_u6_n162 ) , .ZN( u2_u13_u6_n94 ) );
  NOR2_X1 u2_u13_u6_U67 (.A2( u2_u13_X_37 ) , .A1( u2_u13_X_38 ) , .ZN( u2_u13_u6_n91 ) );
  NAND2_X1 u2_u13_u6_U68 (.A1( u2_u13_X_41 ) , .ZN( u2_u13_u6_n144 ) , .A2( u2_u13_u6_n157 ) );
  NAND2_X1 u2_u13_u6_U69 (.A2( u2_u13_X_40 ) , .A1( u2_u13_X_41 ) , .ZN( u2_u13_u6_n139 ) );
  NOR2_X1 u2_u13_u6_U7 (.A1( u2_u13_u6_n118 ) , .ZN( u2_u13_u6_n143 ) , .A2( u2_u13_u6_n168 ) );
  AND2_X1 u2_u13_u6_U70 (.A1( u2_u13_X_39 ) , .A2( u2_u13_u6_n156 ) , .ZN( u2_u13_u6_n96 ) );
  AND2_X1 u2_u13_u6_U71 (.A1( u2_u13_X_39 ) , .A2( u2_u13_X_42 ) , .ZN( u2_u13_u6_n99 ) );
  INV_X1 u2_u13_u6_U72 (.A( u2_u13_X_40 ) , .ZN( u2_u13_u6_n157 ) );
  INV_X1 u2_u13_u6_U73 (.A( u2_u13_X_37 ) , .ZN( u2_u13_u6_n165 ) );
  INV_X1 u2_u13_u6_U74 (.A( u2_u13_X_38 ) , .ZN( u2_u13_u6_n162 ) );
  INV_X1 u2_u13_u6_U75 (.A( u2_u13_X_42 ) , .ZN( u2_u13_u6_n156 ) );
  NAND4_X1 u2_u13_u6_U76 (.ZN( u2_out13_32 ) , .A4( u2_u13_u6_n103 ) , .A3( u2_u13_u6_n104 ) , .A2( u2_u13_u6_n105 ) , .A1( u2_u13_u6_n106 ) );
  AOI22_X1 u2_u13_u6_U77 (.ZN( u2_u13_u6_n105 ) , .A2( u2_u13_u6_n108 ) , .A1( u2_u13_u6_n118 ) , .B2( u2_u13_u6_n126 ) , .B1( u2_u13_u6_n171 ) );
  AOI22_X1 u2_u13_u6_U78 (.ZN( u2_u13_u6_n104 ) , .A1( u2_u13_u6_n111 ) , .B1( u2_u13_u6_n124 ) , .B2( u2_u13_u6_n151 ) , .A2( u2_u13_u6_n93 ) );
  NAND4_X1 u2_u13_u6_U79 (.ZN( u2_out13_12 ) , .A4( u2_u13_u6_n114 ) , .A3( u2_u13_u6_n115 ) , .A2( u2_u13_u6_n116 ) , .A1( u2_u13_u6_n117 ) );
  OAI21_X1 u2_u13_u6_U8 (.A( u2_u13_u6_n159 ) , .B1( u2_u13_u6_n169 ) , .B2( u2_u13_u6_n173 ) , .ZN( u2_u13_u6_n90 ) );
  OAI22_X1 u2_u13_u6_U80 (.B2( u2_u13_u6_n111 ) , .ZN( u2_u13_u6_n116 ) , .B1( u2_u13_u6_n126 ) , .A2( u2_u13_u6_n164 ) , .A1( u2_u13_u6_n167 ) );
  OAI21_X1 u2_u13_u6_U81 (.A( u2_u13_u6_n108 ) , .ZN( u2_u13_u6_n117 ) , .B2( u2_u13_u6_n141 ) , .B1( u2_u13_u6_n163 ) );
  OAI211_X1 u2_u13_u6_U82 (.ZN( u2_out13_7 ) , .B( u2_u13_u6_n153 ) , .C2( u2_u13_u6_n154 ) , .C1( u2_u13_u6_n155 ) , .A( u2_u13_u6_n174 ) );
  NOR3_X1 u2_u13_u6_U83 (.A1( u2_u13_u6_n141 ) , .ZN( u2_u13_u6_n154 ) , .A3( u2_u13_u6_n164 ) , .A2( u2_u13_u6_n171 ) );
  AOI211_X1 u2_u13_u6_U84 (.B( u2_u13_u6_n149 ) , .A( u2_u13_u6_n150 ) , .C2( u2_u13_u6_n151 ) , .C1( u2_u13_u6_n152 ) , .ZN( u2_u13_u6_n153 ) );
  OAI211_X1 u2_u13_u6_U85 (.ZN( u2_out13_22 ) , .B( u2_u13_u6_n137 ) , .A( u2_u13_u6_n138 ) , .C2( u2_u13_u6_n139 ) , .C1( u2_u13_u6_n140 ) );
  AOI22_X1 u2_u13_u6_U86 (.B1( u2_u13_u6_n124 ) , .A2( u2_u13_u6_n125 ) , .A1( u2_u13_u6_n126 ) , .ZN( u2_u13_u6_n138 ) , .B2( u2_u13_u6_n161 ) );
  AND4_X1 u2_u13_u6_U87 (.A3( u2_u13_u6_n119 ) , .A1( u2_u13_u6_n120 ) , .A4( u2_u13_u6_n129 ) , .ZN( u2_u13_u6_n140 ) , .A2( u2_u13_u6_n143 ) );
  NAND3_X1 u2_u13_u6_U88 (.A2( u2_u13_u6_n123 ) , .ZN( u2_u13_u6_n125 ) , .A1( u2_u13_u6_n130 ) , .A3( u2_u13_u6_n131 ) );
  NAND3_X1 u2_u13_u6_U89 (.A3( u2_u13_u6_n133 ) , .ZN( u2_u13_u6_n141 ) , .A1( u2_u13_u6_n145 ) , .A2( u2_u13_u6_n148 ) );
  INV_X1 u2_u13_u6_U9 (.ZN( u2_u13_u6_n172 ) , .A( u2_u13_u6_n88 ) );
  NAND3_X1 u2_u13_u6_U90 (.ZN( u2_u13_u6_n101 ) , .A3( u2_u13_u6_n107 ) , .A2( u2_u13_u6_n121 ) , .A1( u2_u13_u6_n127 ) );
  NAND3_X1 u2_u13_u6_U91 (.ZN( u2_u13_u6_n102 ) , .A3( u2_u13_u6_n130 ) , .A2( u2_u13_u6_n145 ) , .A1( u2_u13_u6_n166 ) );
  NAND3_X1 u2_u13_u6_U92 (.A3( u2_u13_u6_n113 ) , .A1( u2_u13_u6_n119 ) , .A2( u2_u13_u6_n123 ) , .ZN( u2_u13_u6_n93 ) );
  NAND3_X1 u2_u13_u6_U93 (.ZN( u2_u13_u6_n142 ) , .A2( u2_u13_u6_n172 ) , .A3( u2_u13_u6_n89 ) , .A1( u2_u13_u6_n90 ) );
  AND3_X1 u2_u13_u7_U10 (.A3( u2_u13_u7_n110 ) , .A2( u2_u13_u7_n127 ) , .A1( u2_u13_u7_n132 ) , .ZN( u2_u13_u7_n92 ) );
  OAI21_X1 u2_u13_u7_U11 (.A( u2_u13_u7_n161 ) , .B1( u2_u13_u7_n168 ) , .B2( u2_u13_u7_n173 ) , .ZN( u2_u13_u7_n91 ) );
  AOI211_X1 u2_u13_u7_U12 (.A( u2_u13_u7_n117 ) , .ZN( u2_u13_u7_n118 ) , .C2( u2_u13_u7_n126 ) , .C1( u2_u13_u7_n177 ) , .B( u2_u13_u7_n180 ) );
  OAI22_X1 u2_u13_u7_U13 (.B1( u2_u13_u7_n115 ) , .ZN( u2_u13_u7_n117 ) , .A2( u2_u13_u7_n133 ) , .A1( u2_u13_u7_n137 ) , .B2( u2_u13_u7_n162 ) );
  INV_X1 u2_u13_u7_U14 (.A( u2_u13_u7_n116 ) , .ZN( u2_u13_u7_n180 ) );
  NOR3_X1 u2_u13_u7_U15 (.ZN( u2_u13_u7_n115 ) , .A3( u2_u13_u7_n145 ) , .A2( u2_u13_u7_n168 ) , .A1( u2_u13_u7_n169 ) );
  OAI211_X1 u2_u13_u7_U16 (.B( u2_u13_u7_n122 ) , .A( u2_u13_u7_n123 ) , .C2( u2_u13_u7_n124 ) , .ZN( u2_u13_u7_n154 ) , .C1( u2_u13_u7_n162 ) );
  AOI222_X1 u2_u13_u7_U17 (.ZN( u2_u13_u7_n122 ) , .C2( u2_u13_u7_n126 ) , .C1( u2_u13_u7_n145 ) , .B1( u2_u13_u7_n161 ) , .A2( u2_u13_u7_n165 ) , .B2( u2_u13_u7_n170 ) , .A1( u2_u13_u7_n176 ) );
  INV_X1 u2_u13_u7_U18 (.A( u2_u13_u7_n133 ) , .ZN( u2_u13_u7_n176 ) );
  NOR3_X1 u2_u13_u7_U19 (.A2( u2_u13_u7_n134 ) , .A1( u2_u13_u7_n135 ) , .ZN( u2_u13_u7_n136 ) , .A3( u2_u13_u7_n171 ) );
  NOR2_X1 u2_u13_u7_U20 (.A1( u2_u13_u7_n130 ) , .A2( u2_u13_u7_n134 ) , .ZN( u2_u13_u7_n153 ) );
  INV_X1 u2_u13_u7_U21 (.A( u2_u13_u7_n101 ) , .ZN( u2_u13_u7_n165 ) );
  NOR2_X1 u2_u13_u7_U22 (.ZN( u2_u13_u7_n111 ) , .A2( u2_u13_u7_n134 ) , .A1( u2_u13_u7_n169 ) );
  AOI21_X1 u2_u13_u7_U23 (.ZN( u2_u13_u7_n104 ) , .B2( u2_u13_u7_n112 ) , .B1( u2_u13_u7_n127 ) , .A( u2_u13_u7_n164 ) );
  AOI21_X1 u2_u13_u7_U24 (.ZN( u2_u13_u7_n106 ) , .B1( u2_u13_u7_n133 ) , .B2( u2_u13_u7_n146 ) , .A( u2_u13_u7_n162 ) );
  AOI21_X1 u2_u13_u7_U25 (.A( u2_u13_u7_n101 ) , .ZN( u2_u13_u7_n107 ) , .B2( u2_u13_u7_n128 ) , .B1( u2_u13_u7_n175 ) );
  INV_X1 u2_u13_u7_U26 (.A( u2_u13_u7_n138 ) , .ZN( u2_u13_u7_n171 ) );
  INV_X1 u2_u13_u7_U27 (.A( u2_u13_u7_n131 ) , .ZN( u2_u13_u7_n177 ) );
  INV_X1 u2_u13_u7_U28 (.A( u2_u13_u7_n110 ) , .ZN( u2_u13_u7_n174 ) );
  NAND2_X1 u2_u13_u7_U29 (.A1( u2_u13_u7_n129 ) , .A2( u2_u13_u7_n132 ) , .ZN( u2_u13_u7_n149 ) );
  OAI21_X1 u2_u13_u7_U3 (.ZN( u2_u13_u7_n159 ) , .A( u2_u13_u7_n165 ) , .B2( u2_u13_u7_n171 ) , .B1( u2_u13_u7_n174 ) );
  NAND2_X1 u2_u13_u7_U30 (.A1( u2_u13_u7_n113 ) , .A2( u2_u13_u7_n124 ) , .ZN( u2_u13_u7_n130 ) );
  INV_X1 u2_u13_u7_U31 (.A( u2_u13_u7_n112 ) , .ZN( u2_u13_u7_n173 ) );
  INV_X1 u2_u13_u7_U32 (.A( u2_u13_u7_n128 ) , .ZN( u2_u13_u7_n168 ) );
  INV_X1 u2_u13_u7_U33 (.A( u2_u13_u7_n148 ) , .ZN( u2_u13_u7_n169 ) );
  INV_X1 u2_u13_u7_U34 (.A( u2_u13_u7_n127 ) , .ZN( u2_u13_u7_n179 ) );
  NOR2_X1 u2_u13_u7_U35 (.ZN( u2_u13_u7_n101 ) , .A2( u2_u13_u7_n150 ) , .A1( u2_u13_u7_n156 ) );
  AOI211_X1 u2_u13_u7_U36 (.B( u2_u13_u7_n154 ) , .A( u2_u13_u7_n155 ) , .C1( u2_u13_u7_n156 ) , .ZN( u2_u13_u7_n157 ) , .C2( u2_u13_u7_n172 ) );
  INV_X1 u2_u13_u7_U37 (.A( u2_u13_u7_n153 ) , .ZN( u2_u13_u7_n172 ) );
  AOI211_X1 u2_u13_u7_U38 (.B( u2_u13_u7_n139 ) , .A( u2_u13_u7_n140 ) , .C2( u2_u13_u7_n141 ) , .ZN( u2_u13_u7_n142 ) , .C1( u2_u13_u7_n156 ) );
  NAND4_X1 u2_u13_u7_U39 (.A3( u2_u13_u7_n127 ) , .A2( u2_u13_u7_n128 ) , .A1( u2_u13_u7_n129 ) , .ZN( u2_u13_u7_n141 ) , .A4( u2_u13_u7_n147 ) );
  INV_X1 u2_u13_u7_U4 (.A( u2_u13_u7_n111 ) , .ZN( u2_u13_u7_n170 ) );
  AOI21_X1 u2_u13_u7_U40 (.A( u2_u13_u7_n137 ) , .B1( u2_u13_u7_n138 ) , .ZN( u2_u13_u7_n139 ) , .B2( u2_u13_u7_n146 ) );
  OAI22_X1 u2_u13_u7_U41 (.B1( u2_u13_u7_n136 ) , .ZN( u2_u13_u7_n140 ) , .A1( u2_u13_u7_n153 ) , .B2( u2_u13_u7_n162 ) , .A2( u2_u13_u7_n164 ) );
  AOI21_X1 u2_u13_u7_U42 (.ZN( u2_u13_u7_n123 ) , .B1( u2_u13_u7_n165 ) , .B2( u2_u13_u7_n177 ) , .A( u2_u13_u7_n97 ) );
  AOI21_X1 u2_u13_u7_U43 (.B2( u2_u13_u7_n113 ) , .B1( u2_u13_u7_n124 ) , .A( u2_u13_u7_n125 ) , .ZN( u2_u13_u7_n97 ) );
  INV_X1 u2_u13_u7_U44 (.A( u2_u13_u7_n125 ) , .ZN( u2_u13_u7_n161 ) );
  INV_X1 u2_u13_u7_U45 (.A( u2_u13_u7_n152 ) , .ZN( u2_u13_u7_n162 ) );
  AOI22_X1 u2_u13_u7_U46 (.A2( u2_u13_u7_n114 ) , .ZN( u2_u13_u7_n119 ) , .B1( u2_u13_u7_n130 ) , .A1( u2_u13_u7_n156 ) , .B2( u2_u13_u7_n165 ) );
  NAND2_X1 u2_u13_u7_U47 (.A2( u2_u13_u7_n112 ) , .ZN( u2_u13_u7_n114 ) , .A1( u2_u13_u7_n175 ) );
  AND2_X1 u2_u13_u7_U48 (.ZN( u2_u13_u7_n145 ) , .A2( u2_u13_u7_n98 ) , .A1( u2_u13_u7_n99 ) );
  NOR2_X1 u2_u13_u7_U49 (.ZN( u2_u13_u7_n137 ) , .A1( u2_u13_u7_n150 ) , .A2( u2_u13_u7_n161 ) );
  INV_X1 u2_u13_u7_U5 (.A( u2_u13_u7_n149 ) , .ZN( u2_u13_u7_n175 ) );
  AOI21_X1 u2_u13_u7_U50 (.ZN( u2_u13_u7_n105 ) , .B2( u2_u13_u7_n110 ) , .A( u2_u13_u7_n125 ) , .B1( u2_u13_u7_n147 ) );
  NAND2_X1 u2_u13_u7_U51 (.ZN( u2_u13_u7_n146 ) , .A1( u2_u13_u7_n95 ) , .A2( u2_u13_u7_n98 ) );
  NAND2_X1 u2_u13_u7_U52 (.A2( u2_u13_u7_n103 ) , .ZN( u2_u13_u7_n147 ) , .A1( u2_u13_u7_n93 ) );
  NAND2_X1 u2_u13_u7_U53 (.A1( u2_u13_u7_n103 ) , .ZN( u2_u13_u7_n127 ) , .A2( u2_u13_u7_n99 ) );
  OR2_X1 u2_u13_u7_U54 (.ZN( u2_u13_u7_n126 ) , .A2( u2_u13_u7_n152 ) , .A1( u2_u13_u7_n156 ) );
  NAND2_X1 u2_u13_u7_U55 (.A2( u2_u13_u7_n102 ) , .A1( u2_u13_u7_n103 ) , .ZN( u2_u13_u7_n133 ) );
  NAND2_X1 u2_u13_u7_U56 (.ZN( u2_u13_u7_n112 ) , .A2( u2_u13_u7_n96 ) , .A1( u2_u13_u7_n99 ) );
  NAND2_X1 u2_u13_u7_U57 (.A2( u2_u13_u7_n102 ) , .ZN( u2_u13_u7_n128 ) , .A1( u2_u13_u7_n98 ) );
  NAND2_X1 u2_u13_u7_U58 (.A1( u2_u13_u7_n100 ) , .ZN( u2_u13_u7_n113 ) , .A2( u2_u13_u7_n93 ) );
  NAND2_X1 u2_u13_u7_U59 (.A2( u2_u13_u7_n102 ) , .ZN( u2_u13_u7_n124 ) , .A1( u2_u13_u7_n96 ) );
  INV_X1 u2_u13_u7_U6 (.A( u2_u13_u7_n154 ) , .ZN( u2_u13_u7_n178 ) );
  NAND2_X1 u2_u13_u7_U60 (.ZN( u2_u13_u7_n110 ) , .A1( u2_u13_u7_n95 ) , .A2( u2_u13_u7_n96 ) );
  INV_X1 u2_u13_u7_U61 (.A( u2_u13_u7_n150 ) , .ZN( u2_u13_u7_n164 ) );
  AND2_X1 u2_u13_u7_U62 (.ZN( u2_u13_u7_n134 ) , .A1( u2_u13_u7_n93 ) , .A2( u2_u13_u7_n98 ) );
  NAND2_X1 u2_u13_u7_U63 (.A1( u2_u13_u7_n100 ) , .A2( u2_u13_u7_n102 ) , .ZN( u2_u13_u7_n129 ) );
  NAND2_X1 u2_u13_u7_U64 (.A2( u2_u13_u7_n103 ) , .ZN( u2_u13_u7_n131 ) , .A1( u2_u13_u7_n95 ) );
  NAND2_X1 u2_u13_u7_U65 (.A1( u2_u13_u7_n100 ) , .ZN( u2_u13_u7_n138 ) , .A2( u2_u13_u7_n99 ) );
  NAND2_X1 u2_u13_u7_U66 (.ZN( u2_u13_u7_n132 ) , .A1( u2_u13_u7_n93 ) , .A2( u2_u13_u7_n96 ) );
  NAND2_X1 u2_u13_u7_U67 (.A1( u2_u13_u7_n100 ) , .ZN( u2_u13_u7_n148 ) , .A2( u2_u13_u7_n95 ) );
  NOR2_X1 u2_u13_u7_U68 (.A2( u2_u13_X_47 ) , .ZN( u2_u13_u7_n150 ) , .A1( u2_u13_u7_n163 ) );
  NOR2_X1 u2_u13_u7_U69 (.A2( u2_u13_X_43 ) , .A1( u2_u13_X_44 ) , .ZN( u2_u13_u7_n103 ) );
  AOI211_X1 u2_u13_u7_U7 (.ZN( u2_u13_u7_n116 ) , .A( u2_u13_u7_n155 ) , .C1( u2_u13_u7_n161 ) , .C2( u2_u13_u7_n171 ) , .B( u2_u13_u7_n94 ) );
  NOR2_X1 u2_u13_u7_U70 (.A2( u2_u13_X_48 ) , .A1( u2_u13_u7_n166 ) , .ZN( u2_u13_u7_n95 ) );
  NOR2_X1 u2_u13_u7_U71 (.A2( u2_u13_X_45 ) , .A1( u2_u13_X_48 ) , .ZN( u2_u13_u7_n99 ) );
  NOR2_X1 u2_u13_u7_U72 (.A2( u2_u13_X_44 ) , .A1( u2_u13_u7_n167 ) , .ZN( u2_u13_u7_n98 ) );
  NOR2_X1 u2_u13_u7_U73 (.A2( u2_u13_X_46 ) , .A1( u2_u13_X_47 ) , .ZN( u2_u13_u7_n152 ) );
  AND2_X1 u2_u13_u7_U74 (.A1( u2_u13_X_47 ) , .ZN( u2_u13_u7_n156 ) , .A2( u2_u13_u7_n163 ) );
  NAND2_X1 u2_u13_u7_U75 (.A2( u2_u13_X_46 ) , .A1( u2_u13_X_47 ) , .ZN( u2_u13_u7_n125 ) );
  AND2_X1 u2_u13_u7_U76 (.A2( u2_u13_X_45 ) , .A1( u2_u13_X_48 ) , .ZN( u2_u13_u7_n102 ) );
  AND2_X1 u2_u13_u7_U77 (.A2( u2_u13_X_43 ) , .A1( u2_u13_X_44 ) , .ZN( u2_u13_u7_n96 ) );
  AND2_X1 u2_u13_u7_U78 (.A1( u2_u13_X_44 ) , .ZN( u2_u13_u7_n100 ) , .A2( u2_u13_u7_n167 ) );
  AND2_X1 u2_u13_u7_U79 (.A1( u2_u13_X_48 ) , .A2( u2_u13_u7_n166 ) , .ZN( u2_u13_u7_n93 ) );
  OAI222_X1 u2_u13_u7_U8 (.C2( u2_u13_u7_n101 ) , .B2( u2_u13_u7_n111 ) , .A1( u2_u13_u7_n113 ) , .C1( u2_u13_u7_n146 ) , .A2( u2_u13_u7_n162 ) , .B1( u2_u13_u7_n164 ) , .ZN( u2_u13_u7_n94 ) );
  INV_X1 u2_u13_u7_U80 (.A( u2_u13_X_46 ) , .ZN( u2_u13_u7_n163 ) );
  INV_X1 u2_u13_u7_U81 (.A( u2_u13_X_43 ) , .ZN( u2_u13_u7_n167 ) );
  INV_X1 u2_u13_u7_U82 (.A( u2_u13_X_45 ) , .ZN( u2_u13_u7_n166 ) );
  NAND4_X1 u2_u13_u7_U83 (.ZN( u2_out13_27 ) , .A4( u2_u13_u7_n118 ) , .A3( u2_u13_u7_n119 ) , .A2( u2_u13_u7_n120 ) , .A1( u2_u13_u7_n121 ) );
  OAI21_X1 u2_u13_u7_U84 (.ZN( u2_u13_u7_n121 ) , .B2( u2_u13_u7_n145 ) , .A( u2_u13_u7_n150 ) , .B1( u2_u13_u7_n174 ) );
  OAI21_X1 u2_u13_u7_U85 (.ZN( u2_u13_u7_n120 ) , .A( u2_u13_u7_n161 ) , .B2( u2_u13_u7_n170 ) , .B1( u2_u13_u7_n179 ) );
  NAND4_X1 u2_u13_u7_U86 (.ZN( u2_out13_21 ) , .A4( u2_u13_u7_n157 ) , .A3( u2_u13_u7_n158 ) , .A2( u2_u13_u7_n159 ) , .A1( u2_u13_u7_n160 ) );
  OAI21_X1 u2_u13_u7_U87 (.B1( u2_u13_u7_n145 ) , .ZN( u2_u13_u7_n160 ) , .A( u2_u13_u7_n161 ) , .B2( u2_u13_u7_n177 ) );
  AOI22_X1 u2_u13_u7_U88 (.B2( u2_u13_u7_n149 ) , .B1( u2_u13_u7_n150 ) , .A2( u2_u13_u7_n151 ) , .A1( u2_u13_u7_n152 ) , .ZN( u2_u13_u7_n158 ) );
  NAND4_X1 u2_u13_u7_U89 (.ZN( u2_out13_15 ) , .A4( u2_u13_u7_n142 ) , .A3( u2_u13_u7_n143 ) , .A2( u2_u13_u7_n144 ) , .A1( u2_u13_u7_n178 ) );
  OAI221_X1 u2_u13_u7_U9 (.C1( u2_u13_u7_n101 ) , .C2( u2_u13_u7_n147 ) , .ZN( u2_u13_u7_n155 ) , .B2( u2_u13_u7_n162 ) , .A( u2_u13_u7_n91 ) , .B1( u2_u13_u7_n92 ) );
  OR2_X1 u2_u13_u7_U90 (.A2( u2_u13_u7_n125 ) , .A1( u2_u13_u7_n129 ) , .ZN( u2_u13_u7_n144 ) );
  AOI22_X1 u2_u13_u7_U91 (.A2( u2_u13_u7_n126 ) , .ZN( u2_u13_u7_n143 ) , .B2( u2_u13_u7_n165 ) , .B1( u2_u13_u7_n173 ) , .A1( u2_u13_u7_n174 ) );
  NAND4_X1 u2_u13_u7_U92 (.ZN( u2_out13_5 ) , .A4( u2_u13_u7_n108 ) , .A3( u2_u13_u7_n109 ) , .A1( u2_u13_u7_n116 ) , .A2( u2_u13_u7_n123 ) );
  AOI22_X1 u2_u13_u7_U93 (.ZN( u2_u13_u7_n109 ) , .A2( u2_u13_u7_n126 ) , .B2( u2_u13_u7_n145 ) , .B1( u2_u13_u7_n156 ) , .A1( u2_u13_u7_n171 ) );
  NOR4_X1 u2_u13_u7_U94 (.A4( u2_u13_u7_n104 ) , .A3( u2_u13_u7_n105 ) , .A2( u2_u13_u7_n106 ) , .A1( u2_u13_u7_n107 ) , .ZN( u2_u13_u7_n108 ) );
  NAND3_X1 u2_u13_u7_U95 (.A3( u2_u13_u7_n146 ) , .A2( u2_u13_u7_n147 ) , .A1( u2_u13_u7_n148 ) , .ZN( u2_u13_u7_n151 ) );
  NAND3_X1 u2_u13_u7_U96 (.A3( u2_u13_u7_n131 ) , .A2( u2_u13_u7_n132 ) , .A1( u2_u13_u7_n133 ) , .ZN( u2_u13_u7_n135 ) );
  XOR2_X1 u2_u14_U11 (.B( u2_K15_44 ) , .A( u2_R13_29 ) , .Z( u2_u14_X_44 ) );
  XOR2_X1 u2_u14_U13 (.B( u2_K15_42 ) , .A( u2_R13_29 ) , .Z( u2_u14_X_42 ) );
  XOR2_X1 u2_u14_U15 (.B( u2_K15_40 ) , .A( u2_R13_27 ) , .Z( u2_u14_X_40 ) );
  XOR2_X1 u2_u14_U18 (.B( u2_K15_38 ) , .A( u2_R13_25 ) , .Z( u2_u14_X_38 ) );
  XOR2_X1 u2_u14_U19 (.B( u2_K15_37 ) , .A( u2_R13_24 ) , .Z( u2_u14_X_37 ) );
  XOR2_X1 u2_u14_U2 (.B( u2_K15_8 ) , .A( u2_R13_5 ) , .Z( u2_u14_X_8 ) );
  XOR2_X1 u2_u14_U20 (.B( u2_K15_36 ) , .A( u2_R13_25 ) , .Z( u2_u14_X_36 ) );
  XOR2_X1 u2_u14_U21 (.B( u2_K15_35 ) , .A( u2_R13_24 ) , .Z( u2_u14_X_35 ) );
  XOR2_X1 u2_u14_U23 (.B( u2_K15_33 ) , .A( u2_R13_22 ) , .Z( u2_u14_X_33 ) );
  XOR2_X1 u2_u14_U25 (.B( u2_K15_31 ) , .A( u2_R13_20 ) , .Z( u2_u14_X_31 ) );
  XOR2_X1 u2_u14_U27 (.B( u2_K15_2 ) , .A( u2_R13_1 ) , .Z( u2_u14_X_2 ) );
  XOR2_X1 u2_u14_U28 (.B( u2_K15_29 ) , .A( u2_R13_20 ) , .Z( u2_u14_X_29 ) );
  XOR2_X1 u2_u14_U31 (.B( u2_K15_26 ) , .A( u2_R13_17 ) , .Z( u2_u14_X_26 ) );
  XOR2_X1 u2_u14_U32 (.B( u2_K15_25 ) , .A( u2_R13_16 ) , .Z( u2_u14_X_25 ) );
  XOR2_X1 u2_u14_U33 (.B( u2_K15_24 ) , .A( u2_R13_17 ) , .Z( u2_u14_X_24 ) );
  XOR2_X1 u2_u14_U34 (.B( u2_K15_23 ) , .A( u2_R13_16 ) , .Z( u2_u14_X_23 ) );
  XOR2_X1 u2_u14_U38 (.B( u2_K15_1 ) , .A( u2_R13_32 ) , .Z( u2_u14_X_1 ) );
  XOR2_X1 u2_u14_U39 (.B( u2_K15_19 ) , .A( u2_R13_12 ) , .Z( u2_u14_X_19 ) );
  XOR2_X1 u2_u14_U4 (.B( u2_K15_6 ) , .A( u2_R13_5 ) , .Z( u2_u14_X_6 ) );
  XOR2_X1 u2_u14_U41 (.B( u2_K15_17 ) , .A( u2_R13_12 ) , .Z( u2_u14_X_17 ) );
  XOR2_X1 u2_u14_U44 (.B( u2_K15_14 ) , .A( u2_R13_9 ) , .Z( u2_u14_X_14 ) );
  XOR2_X1 u2_u14_U46 (.B( u2_K15_12 ) , .A( u2_R13_9 ) , .Z( u2_u14_X_12 ) );
  XOR2_X1 u2_u14_U7 (.B( u2_K15_48 ) , .A( u2_R13_1 ) , .Z( u2_u14_X_48 ) );
  XOR2_X1 u2_u14_U8 (.B( u2_K15_47 ) , .A( u2_R13_32 ) , .Z( u2_u14_X_47 ) );
  AND3_X1 u2_u14_u0_U10 (.A2( u2_u14_u0_n112 ) , .ZN( u2_u14_u0_n127 ) , .A3( u2_u14_u0_n130 ) , .A1( u2_u14_u0_n148 ) );
  NAND2_X1 u2_u14_u0_U11 (.ZN( u2_u14_u0_n113 ) , .A1( u2_u14_u0_n139 ) , .A2( u2_u14_u0_n149 ) );
  AND2_X1 u2_u14_u0_U12 (.ZN( u2_u14_u0_n107 ) , .A1( u2_u14_u0_n130 ) , .A2( u2_u14_u0_n140 ) );
  AND2_X1 u2_u14_u0_U13 (.A2( u2_u14_u0_n129 ) , .A1( u2_u14_u0_n130 ) , .ZN( u2_u14_u0_n151 ) );
  AND2_X1 u2_u14_u0_U14 (.A1( u2_u14_u0_n108 ) , .A2( u2_u14_u0_n125 ) , .ZN( u2_u14_u0_n145 ) );
  INV_X1 u2_u14_u0_U15 (.A( u2_u14_u0_n143 ) , .ZN( u2_u14_u0_n173 ) );
  NOR2_X1 u2_u14_u0_U16 (.A2( u2_u14_u0_n136 ) , .ZN( u2_u14_u0_n147 ) , .A1( u2_u14_u0_n160 ) );
  NOR2_X1 u2_u14_u0_U17 (.A1( u2_u14_u0_n163 ) , .A2( u2_u14_u0_n164 ) , .ZN( u2_u14_u0_n95 ) );
  AOI21_X1 u2_u14_u0_U18 (.B1( u2_u14_u0_n103 ) , .ZN( u2_u14_u0_n132 ) , .A( u2_u14_u0_n165 ) , .B2( u2_u14_u0_n93 ) );
  INV_X1 u2_u14_u0_U19 (.A( u2_u14_u0_n142 ) , .ZN( u2_u14_u0_n165 ) );
  OAI221_X1 u2_u14_u0_U20 (.C1( u2_u14_u0_n121 ) , .ZN( u2_u14_u0_n122 ) , .B2( u2_u14_u0_n127 ) , .A( u2_u14_u0_n143 ) , .B1( u2_u14_u0_n144 ) , .C2( u2_u14_u0_n147 ) );
  OAI22_X1 u2_u14_u0_U21 (.B1( u2_u14_u0_n125 ) , .ZN( u2_u14_u0_n126 ) , .A1( u2_u14_u0_n138 ) , .A2( u2_u14_u0_n146 ) , .B2( u2_u14_u0_n147 ) );
  OAI22_X1 u2_u14_u0_U22 (.B1( u2_u14_u0_n131 ) , .A1( u2_u14_u0_n144 ) , .B2( u2_u14_u0_n147 ) , .A2( u2_u14_u0_n90 ) , .ZN( u2_u14_u0_n91 ) );
  AND3_X1 u2_u14_u0_U23 (.A3( u2_u14_u0_n121 ) , .A2( u2_u14_u0_n125 ) , .A1( u2_u14_u0_n148 ) , .ZN( u2_u14_u0_n90 ) );
  INV_X1 u2_u14_u0_U24 (.A( u2_u14_u0_n136 ) , .ZN( u2_u14_u0_n161 ) );
  NOR2_X1 u2_u14_u0_U25 (.A1( u2_u14_u0_n120 ) , .ZN( u2_u14_u0_n143 ) , .A2( u2_u14_u0_n167 ) );
  OAI221_X1 u2_u14_u0_U26 (.C1( u2_u14_u0_n112 ) , .ZN( u2_u14_u0_n120 ) , .B1( u2_u14_u0_n138 ) , .B2( u2_u14_u0_n141 ) , .C2( u2_u14_u0_n147 ) , .A( u2_u14_u0_n172 ) );
  AOI211_X1 u2_u14_u0_U27 (.B( u2_u14_u0_n115 ) , .A( u2_u14_u0_n116 ) , .C2( u2_u14_u0_n117 ) , .C1( u2_u14_u0_n118 ) , .ZN( u2_u14_u0_n119 ) );
  AOI22_X1 u2_u14_u0_U28 (.B2( u2_u14_u0_n109 ) , .A2( u2_u14_u0_n110 ) , .ZN( u2_u14_u0_n111 ) , .B1( u2_u14_u0_n118 ) , .A1( u2_u14_u0_n160 ) );
  INV_X1 u2_u14_u0_U29 (.A( u2_u14_u0_n118 ) , .ZN( u2_u14_u0_n158 ) );
  INV_X1 u2_u14_u0_U3 (.A( u2_u14_u0_n113 ) , .ZN( u2_u14_u0_n166 ) );
  AOI21_X1 u2_u14_u0_U30 (.ZN( u2_u14_u0_n104 ) , .B1( u2_u14_u0_n107 ) , .B2( u2_u14_u0_n141 ) , .A( u2_u14_u0_n144 ) );
  AOI21_X1 u2_u14_u0_U31 (.B1( u2_u14_u0_n127 ) , .B2( u2_u14_u0_n129 ) , .A( u2_u14_u0_n138 ) , .ZN( u2_u14_u0_n96 ) );
  AOI21_X1 u2_u14_u0_U32 (.ZN( u2_u14_u0_n116 ) , .B2( u2_u14_u0_n142 ) , .A( u2_u14_u0_n144 ) , .B1( u2_u14_u0_n166 ) );
  NAND2_X1 u2_u14_u0_U33 (.A1( u2_u14_u0_n100 ) , .A2( u2_u14_u0_n103 ) , .ZN( u2_u14_u0_n125 ) );
  NAND2_X1 u2_u14_u0_U34 (.A2( u2_u14_u0_n103 ) , .ZN( u2_u14_u0_n140 ) , .A1( u2_u14_u0_n94 ) );
  NAND2_X1 u2_u14_u0_U35 (.A1( u2_u14_u0_n101 ) , .A2( u2_u14_u0_n102 ) , .ZN( u2_u14_u0_n150 ) );
  INV_X1 u2_u14_u0_U36 (.A( u2_u14_u0_n138 ) , .ZN( u2_u14_u0_n160 ) );
  NAND2_X1 u2_u14_u0_U37 (.ZN( u2_u14_u0_n142 ) , .A1( u2_u14_u0_n94 ) , .A2( u2_u14_u0_n95 ) );
  NAND2_X1 u2_u14_u0_U38 (.A1( u2_u14_u0_n102 ) , .ZN( u2_u14_u0_n128 ) , .A2( u2_u14_u0_n95 ) );
  NAND2_X1 u2_u14_u0_U39 (.A2( u2_u14_u0_n102 ) , .A1( u2_u14_u0_n103 ) , .ZN( u2_u14_u0_n149 ) );
  AOI21_X1 u2_u14_u0_U4 (.B1( u2_u14_u0_n114 ) , .ZN( u2_u14_u0_n115 ) , .B2( u2_u14_u0_n129 ) , .A( u2_u14_u0_n161 ) );
  NAND2_X1 u2_u14_u0_U40 (.A1( u2_u14_u0_n100 ) , .ZN( u2_u14_u0_n129 ) , .A2( u2_u14_u0_n95 ) );
  NAND2_X1 u2_u14_u0_U41 (.A2( u2_u14_u0_n100 ) , .A1( u2_u14_u0_n101 ) , .ZN( u2_u14_u0_n139 ) );
  NAND2_X1 u2_u14_u0_U42 (.A2( u2_u14_u0_n100 ) , .ZN( u2_u14_u0_n131 ) , .A1( u2_u14_u0_n92 ) );
  NAND2_X1 u2_u14_u0_U43 (.ZN( u2_u14_u0_n108 ) , .A1( u2_u14_u0_n92 ) , .A2( u2_u14_u0_n94 ) );
  NAND2_X1 u2_u14_u0_U44 (.ZN( u2_u14_u0_n148 ) , .A1( u2_u14_u0_n93 ) , .A2( u2_u14_u0_n95 ) );
  NAND2_X1 u2_u14_u0_U45 (.A2( u2_u14_u0_n102 ) , .ZN( u2_u14_u0_n114 ) , .A1( u2_u14_u0_n92 ) );
  NAND2_X1 u2_u14_u0_U46 (.A1( u2_u14_u0_n101 ) , .ZN( u2_u14_u0_n130 ) , .A2( u2_u14_u0_n94 ) );
  NAND2_X1 u2_u14_u0_U47 (.A2( u2_u14_u0_n101 ) , .ZN( u2_u14_u0_n121 ) , .A1( u2_u14_u0_n93 ) );
  INV_X1 u2_u14_u0_U48 (.ZN( u2_u14_u0_n172 ) , .A( u2_u14_u0_n88 ) );
  OAI222_X1 u2_u14_u0_U49 (.C1( u2_u14_u0_n108 ) , .A1( u2_u14_u0_n125 ) , .B2( u2_u14_u0_n128 ) , .B1( u2_u14_u0_n144 ) , .A2( u2_u14_u0_n158 ) , .C2( u2_u14_u0_n161 ) , .ZN( u2_u14_u0_n88 ) );
  AOI21_X1 u2_u14_u0_U5 (.B2( u2_u14_u0_n131 ) , .ZN( u2_u14_u0_n134 ) , .B1( u2_u14_u0_n151 ) , .A( u2_u14_u0_n158 ) );
  NAND2_X1 u2_u14_u0_U50 (.ZN( u2_u14_u0_n112 ) , .A2( u2_u14_u0_n92 ) , .A1( u2_u14_u0_n93 ) );
  OR3_X1 u2_u14_u0_U51 (.A3( u2_u14_u0_n152 ) , .A2( u2_u14_u0_n153 ) , .A1( u2_u14_u0_n154 ) , .ZN( u2_u14_u0_n155 ) );
  AOI21_X1 u2_u14_u0_U52 (.B2( u2_u14_u0_n150 ) , .B1( u2_u14_u0_n151 ) , .ZN( u2_u14_u0_n152 ) , .A( u2_u14_u0_n158 ) );
  AOI21_X1 u2_u14_u0_U53 (.A( u2_u14_u0_n144 ) , .B2( u2_u14_u0_n145 ) , .B1( u2_u14_u0_n146 ) , .ZN( u2_u14_u0_n154 ) );
  AOI21_X1 u2_u14_u0_U54 (.A( u2_u14_u0_n147 ) , .B2( u2_u14_u0_n148 ) , .B1( u2_u14_u0_n149 ) , .ZN( u2_u14_u0_n153 ) );
  INV_X1 u2_u14_u0_U55 (.ZN( u2_u14_u0_n171 ) , .A( u2_u14_u0_n99 ) );
  OAI211_X1 u2_u14_u0_U56 (.C2( u2_u14_u0_n140 ) , .C1( u2_u14_u0_n161 ) , .A( u2_u14_u0_n169 ) , .B( u2_u14_u0_n98 ) , .ZN( u2_u14_u0_n99 ) );
  INV_X1 u2_u14_u0_U57 (.ZN( u2_u14_u0_n169 ) , .A( u2_u14_u0_n91 ) );
  AOI211_X1 u2_u14_u0_U58 (.C1( u2_u14_u0_n118 ) , .A( u2_u14_u0_n123 ) , .B( u2_u14_u0_n96 ) , .C2( u2_u14_u0_n97 ) , .ZN( u2_u14_u0_n98 ) );
  NOR2_X1 u2_u14_u0_U59 (.A2( u2_u14_X_2 ) , .ZN( u2_u14_u0_n103 ) , .A1( u2_u14_u0_n164 ) );
  NOR2_X1 u2_u14_u0_U6 (.A1( u2_u14_u0_n108 ) , .ZN( u2_u14_u0_n123 ) , .A2( u2_u14_u0_n158 ) );
  NOR2_X1 u2_u14_u0_U60 (.A2( u2_u14_X_3 ) , .A1( u2_u14_X_6 ) , .ZN( u2_u14_u0_n94 ) );
  NOR2_X1 u2_u14_u0_U61 (.A2( u2_u14_X_6 ) , .ZN( u2_u14_u0_n100 ) , .A1( u2_u14_u0_n162 ) );
  NOR2_X1 u2_u14_u0_U62 (.A2( u2_u14_X_4 ) , .A1( u2_u14_X_5 ) , .ZN( u2_u14_u0_n118 ) );
  NOR2_X1 u2_u14_u0_U63 (.A2( u2_u14_X_1 ) , .A1( u2_u14_X_2 ) , .ZN( u2_u14_u0_n92 ) );
  NOR2_X1 u2_u14_u0_U64 (.A2( u2_u14_X_1 ) , .ZN( u2_u14_u0_n101 ) , .A1( u2_u14_u0_n163 ) );
  NAND2_X1 u2_u14_u0_U65 (.A2( u2_u14_X_4 ) , .A1( u2_u14_X_5 ) , .ZN( u2_u14_u0_n144 ) );
  NOR2_X1 u2_u14_u0_U66 (.A2( u2_u14_X_5 ) , .ZN( u2_u14_u0_n136 ) , .A1( u2_u14_u0_n159 ) );
  NAND2_X1 u2_u14_u0_U67 (.A1( u2_u14_X_5 ) , .ZN( u2_u14_u0_n138 ) , .A2( u2_u14_u0_n159 ) );
  AND2_X1 u2_u14_u0_U68 (.A2( u2_u14_X_3 ) , .A1( u2_u14_X_6 ) , .ZN( u2_u14_u0_n102 ) );
  AND2_X1 u2_u14_u0_U69 (.A1( u2_u14_X_6 ) , .A2( u2_u14_u0_n162 ) , .ZN( u2_u14_u0_n93 ) );
  OAI21_X1 u2_u14_u0_U7 (.B1( u2_u14_u0_n150 ) , .B2( u2_u14_u0_n158 ) , .A( u2_u14_u0_n172 ) , .ZN( u2_u14_u0_n89 ) );
  INV_X1 u2_u14_u0_U70 (.A( u2_u14_X_4 ) , .ZN( u2_u14_u0_n159 ) );
  INV_X1 u2_u14_u0_U71 (.A( u2_u14_X_1 ) , .ZN( u2_u14_u0_n164 ) );
  INV_X1 u2_u14_u0_U72 (.A( u2_u14_X_2 ) , .ZN( u2_u14_u0_n163 ) );
  INV_X1 u2_u14_u0_U73 (.A( u2_u14_X_3 ) , .ZN( u2_u14_u0_n162 ) );
  INV_X1 u2_u14_u0_U74 (.A( u2_u14_u0_n126 ) , .ZN( u2_u14_u0_n168 ) );
  AOI211_X1 u2_u14_u0_U75 (.B( u2_u14_u0_n133 ) , .A( u2_u14_u0_n134 ) , .C2( u2_u14_u0_n135 ) , .C1( u2_u14_u0_n136 ) , .ZN( u2_u14_u0_n137 ) );
  INV_X1 u2_u14_u0_U76 (.ZN( u2_u14_u0_n174 ) , .A( u2_u14_u0_n89 ) );
  AOI211_X1 u2_u14_u0_U77 (.B( u2_u14_u0_n104 ) , .A( u2_u14_u0_n105 ) , .ZN( u2_u14_u0_n106 ) , .C2( u2_u14_u0_n113 ) , .C1( u2_u14_u0_n160 ) );
  OR4_X1 u2_u14_u0_U78 (.ZN( u2_out14_17 ) , .A4( u2_u14_u0_n122 ) , .A2( u2_u14_u0_n123 ) , .A1( u2_u14_u0_n124 ) , .A3( u2_u14_u0_n170 ) );
  AOI21_X1 u2_u14_u0_U79 (.B2( u2_u14_u0_n107 ) , .ZN( u2_u14_u0_n124 ) , .B1( u2_u14_u0_n128 ) , .A( u2_u14_u0_n161 ) );
  AND2_X1 u2_u14_u0_U8 (.A1( u2_u14_u0_n114 ) , .A2( u2_u14_u0_n121 ) , .ZN( u2_u14_u0_n146 ) );
  INV_X1 u2_u14_u0_U80 (.A( u2_u14_u0_n111 ) , .ZN( u2_u14_u0_n170 ) );
  OR4_X1 u2_u14_u0_U81 (.ZN( u2_out14_31 ) , .A4( u2_u14_u0_n155 ) , .A2( u2_u14_u0_n156 ) , .A1( u2_u14_u0_n157 ) , .A3( u2_u14_u0_n173 ) );
  AOI21_X1 u2_u14_u0_U82 (.A( u2_u14_u0_n138 ) , .B2( u2_u14_u0_n139 ) , .B1( u2_u14_u0_n140 ) , .ZN( u2_u14_u0_n157 ) );
  AOI21_X1 u2_u14_u0_U83 (.B2( u2_u14_u0_n141 ) , .B1( u2_u14_u0_n142 ) , .ZN( u2_u14_u0_n156 ) , .A( u2_u14_u0_n161 ) );
  AOI21_X1 u2_u14_u0_U84 (.B1( u2_u14_u0_n132 ) , .ZN( u2_u14_u0_n133 ) , .A( u2_u14_u0_n144 ) , .B2( u2_u14_u0_n166 ) );
  OAI22_X1 u2_u14_u0_U85 (.ZN( u2_u14_u0_n105 ) , .A2( u2_u14_u0_n132 ) , .B1( u2_u14_u0_n146 ) , .A1( u2_u14_u0_n147 ) , .B2( u2_u14_u0_n161 ) );
  NAND2_X1 u2_u14_u0_U86 (.ZN( u2_u14_u0_n110 ) , .A2( u2_u14_u0_n132 ) , .A1( u2_u14_u0_n145 ) );
  INV_X1 u2_u14_u0_U87 (.A( u2_u14_u0_n119 ) , .ZN( u2_u14_u0_n167 ) );
  NAND3_X1 u2_u14_u0_U88 (.ZN( u2_out14_23 ) , .A3( u2_u14_u0_n137 ) , .A1( u2_u14_u0_n168 ) , .A2( u2_u14_u0_n171 ) );
  NAND3_X1 u2_u14_u0_U89 (.A3( u2_u14_u0_n127 ) , .A2( u2_u14_u0_n128 ) , .ZN( u2_u14_u0_n135 ) , .A1( u2_u14_u0_n150 ) );
  AND2_X1 u2_u14_u0_U9 (.A1( u2_u14_u0_n131 ) , .ZN( u2_u14_u0_n141 ) , .A2( u2_u14_u0_n150 ) );
  NAND3_X1 u2_u14_u0_U90 (.ZN( u2_u14_u0_n117 ) , .A3( u2_u14_u0_n132 ) , .A2( u2_u14_u0_n139 ) , .A1( u2_u14_u0_n148 ) );
  NAND3_X1 u2_u14_u0_U91 (.ZN( u2_u14_u0_n109 ) , .A2( u2_u14_u0_n114 ) , .A3( u2_u14_u0_n140 ) , .A1( u2_u14_u0_n149 ) );
  NAND3_X1 u2_u14_u0_U92 (.ZN( u2_out14_9 ) , .A3( u2_u14_u0_n106 ) , .A2( u2_u14_u0_n171 ) , .A1( u2_u14_u0_n174 ) );
  NAND3_X1 u2_u14_u0_U93 (.A2( u2_u14_u0_n128 ) , .A1( u2_u14_u0_n132 ) , .A3( u2_u14_u0_n146 ) , .ZN( u2_u14_u0_n97 ) );
  AOI21_X1 u2_u14_u1_U10 (.ZN( u2_u14_u1_n106 ) , .A( u2_u14_u1_n112 ) , .B1( u2_u14_u1_n154 ) , .B2( u2_u14_u1_n156 ) );
  NAND3_X1 u2_u14_u1_U100 (.ZN( u2_u14_u1_n113 ) , .A1( u2_u14_u1_n120 ) , .A3( u2_u14_u1_n133 ) , .A2( u2_u14_u1_n155 ) );
  INV_X1 u2_u14_u1_U11 (.A( u2_u14_u1_n101 ) , .ZN( u2_u14_u1_n184 ) );
  AOI21_X1 u2_u14_u1_U12 (.ZN( u2_u14_u1_n107 ) , .B1( u2_u14_u1_n134 ) , .B2( u2_u14_u1_n149 ) , .A( u2_u14_u1_n174 ) );
  NAND2_X1 u2_u14_u1_U13 (.ZN( u2_u14_u1_n140 ) , .A2( u2_u14_u1_n150 ) , .A1( u2_u14_u1_n155 ) );
  NAND2_X1 u2_u14_u1_U14 (.A1( u2_u14_u1_n131 ) , .ZN( u2_u14_u1_n147 ) , .A2( u2_u14_u1_n153 ) );
  AOI22_X1 u2_u14_u1_U15 (.B2( u2_u14_u1_n136 ) , .A2( u2_u14_u1_n137 ) , .ZN( u2_u14_u1_n143 ) , .A1( u2_u14_u1_n171 ) , .B1( u2_u14_u1_n173 ) );
  INV_X1 u2_u14_u1_U16 (.A( u2_u14_u1_n147 ) , .ZN( u2_u14_u1_n181 ) );
  INV_X1 u2_u14_u1_U17 (.A( u2_u14_u1_n139 ) , .ZN( u2_u14_u1_n174 ) );
  INV_X1 u2_u14_u1_U18 (.A( u2_u14_u1_n112 ) , .ZN( u2_u14_u1_n171 ) );
  NAND2_X1 u2_u14_u1_U19 (.ZN( u2_u14_u1_n141 ) , .A1( u2_u14_u1_n153 ) , .A2( u2_u14_u1_n156 ) );
  AND2_X1 u2_u14_u1_U20 (.A1( u2_u14_u1_n123 ) , .ZN( u2_u14_u1_n134 ) , .A2( u2_u14_u1_n161 ) );
  NAND2_X1 u2_u14_u1_U21 (.A2( u2_u14_u1_n115 ) , .A1( u2_u14_u1_n116 ) , .ZN( u2_u14_u1_n148 ) );
  NAND2_X1 u2_u14_u1_U22 (.A2( u2_u14_u1_n133 ) , .A1( u2_u14_u1_n135 ) , .ZN( u2_u14_u1_n159 ) );
  NAND2_X1 u2_u14_u1_U23 (.A2( u2_u14_u1_n115 ) , .A1( u2_u14_u1_n120 ) , .ZN( u2_u14_u1_n132 ) );
  INV_X1 u2_u14_u1_U24 (.A( u2_u14_u1_n154 ) , .ZN( u2_u14_u1_n178 ) );
  AOI22_X1 u2_u14_u1_U25 (.B2( u2_u14_u1_n113 ) , .A2( u2_u14_u1_n114 ) , .ZN( u2_u14_u1_n125 ) , .A1( u2_u14_u1_n171 ) , .B1( u2_u14_u1_n173 ) );
  NAND2_X1 u2_u14_u1_U26 (.ZN( u2_u14_u1_n114 ) , .A1( u2_u14_u1_n134 ) , .A2( u2_u14_u1_n156 ) );
  INV_X1 u2_u14_u1_U27 (.A( u2_u14_u1_n151 ) , .ZN( u2_u14_u1_n183 ) );
  AND2_X1 u2_u14_u1_U28 (.A1( u2_u14_u1_n129 ) , .A2( u2_u14_u1_n133 ) , .ZN( u2_u14_u1_n149 ) );
  INV_X1 u2_u14_u1_U29 (.A( u2_u14_u1_n131 ) , .ZN( u2_u14_u1_n180 ) );
  INV_X1 u2_u14_u1_U3 (.A( u2_u14_u1_n159 ) , .ZN( u2_u14_u1_n182 ) );
  AOI221_X1 u2_u14_u1_U30 (.B1( u2_u14_u1_n140 ) , .ZN( u2_u14_u1_n167 ) , .B2( u2_u14_u1_n172 ) , .C2( u2_u14_u1_n175 ) , .C1( u2_u14_u1_n178 ) , .A( u2_u14_u1_n188 ) );
  INV_X1 u2_u14_u1_U31 (.ZN( u2_u14_u1_n188 ) , .A( u2_u14_u1_n97 ) );
  AOI211_X1 u2_u14_u1_U32 (.A( u2_u14_u1_n118 ) , .C1( u2_u14_u1_n132 ) , .C2( u2_u14_u1_n139 ) , .B( u2_u14_u1_n96 ) , .ZN( u2_u14_u1_n97 ) );
  AOI21_X1 u2_u14_u1_U33 (.B2( u2_u14_u1_n121 ) , .B1( u2_u14_u1_n135 ) , .A( u2_u14_u1_n152 ) , .ZN( u2_u14_u1_n96 ) );
  OAI221_X1 u2_u14_u1_U34 (.A( u2_u14_u1_n119 ) , .C2( u2_u14_u1_n129 ) , .ZN( u2_u14_u1_n138 ) , .B2( u2_u14_u1_n152 ) , .C1( u2_u14_u1_n174 ) , .B1( u2_u14_u1_n187 ) );
  INV_X1 u2_u14_u1_U35 (.A( u2_u14_u1_n148 ) , .ZN( u2_u14_u1_n187 ) );
  AOI211_X1 u2_u14_u1_U36 (.B( u2_u14_u1_n117 ) , .A( u2_u14_u1_n118 ) , .ZN( u2_u14_u1_n119 ) , .C2( u2_u14_u1_n146 ) , .C1( u2_u14_u1_n159 ) );
  NOR2_X1 u2_u14_u1_U37 (.A1( u2_u14_u1_n168 ) , .A2( u2_u14_u1_n176 ) , .ZN( u2_u14_u1_n98 ) );
  AOI211_X1 u2_u14_u1_U38 (.B( u2_u14_u1_n162 ) , .A( u2_u14_u1_n163 ) , .C2( u2_u14_u1_n164 ) , .ZN( u2_u14_u1_n165 ) , .C1( u2_u14_u1_n171 ) );
  AOI21_X1 u2_u14_u1_U39 (.A( u2_u14_u1_n160 ) , .B2( u2_u14_u1_n161 ) , .ZN( u2_u14_u1_n162 ) , .B1( u2_u14_u1_n182 ) );
  AOI221_X1 u2_u14_u1_U4 (.A( u2_u14_u1_n138 ) , .C2( u2_u14_u1_n139 ) , .C1( u2_u14_u1_n140 ) , .B2( u2_u14_u1_n141 ) , .ZN( u2_u14_u1_n142 ) , .B1( u2_u14_u1_n175 ) );
  OR2_X1 u2_u14_u1_U40 (.A2( u2_u14_u1_n157 ) , .A1( u2_u14_u1_n158 ) , .ZN( u2_u14_u1_n163 ) );
  OAI21_X1 u2_u14_u1_U41 (.B2( u2_u14_u1_n123 ) , .ZN( u2_u14_u1_n145 ) , .B1( u2_u14_u1_n160 ) , .A( u2_u14_u1_n185 ) );
  INV_X1 u2_u14_u1_U42 (.A( u2_u14_u1_n122 ) , .ZN( u2_u14_u1_n185 ) );
  AOI21_X1 u2_u14_u1_U43 (.B2( u2_u14_u1_n120 ) , .B1( u2_u14_u1_n121 ) , .ZN( u2_u14_u1_n122 ) , .A( u2_u14_u1_n128 ) );
  NAND2_X1 u2_u14_u1_U44 (.A1( u2_u14_u1_n128 ) , .ZN( u2_u14_u1_n146 ) , .A2( u2_u14_u1_n160 ) );
  NAND2_X1 u2_u14_u1_U45 (.A2( u2_u14_u1_n112 ) , .ZN( u2_u14_u1_n139 ) , .A1( u2_u14_u1_n152 ) );
  NAND2_X1 u2_u14_u1_U46 (.A1( u2_u14_u1_n105 ) , .ZN( u2_u14_u1_n156 ) , .A2( u2_u14_u1_n99 ) );
  NOR2_X1 u2_u14_u1_U47 (.ZN( u2_u14_u1_n117 ) , .A1( u2_u14_u1_n121 ) , .A2( u2_u14_u1_n160 ) );
  AOI21_X1 u2_u14_u1_U48 (.A( u2_u14_u1_n128 ) , .B2( u2_u14_u1_n129 ) , .ZN( u2_u14_u1_n130 ) , .B1( u2_u14_u1_n150 ) );
  NAND2_X1 u2_u14_u1_U49 (.ZN( u2_u14_u1_n112 ) , .A1( u2_u14_u1_n169 ) , .A2( u2_u14_u1_n170 ) );
  AOI211_X1 u2_u14_u1_U5 (.ZN( u2_u14_u1_n124 ) , .A( u2_u14_u1_n138 ) , .C2( u2_u14_u1_n139 ) , .B( u2_u14_u1_n145 ) , .C1( u2_u14_u1_n147 ) );
  NAND2_X1 u2_u14_u1_U50 (.ZN( u2_u14_u1_n129 ) , .A2( u2_u14_u1_n95 ) , .A1( u2_u14_u1_n98 ) );
  NAND2_X1 u2_u14_u1_U51 (.A1( u2_u14_u1_n102 ) , .ZN( u2_u14_u1_n154 ) , .A2( u2_u14_u1_n99 ) );
  NAND2_X1 u2_u14_u1_U52 (.A2( u2_u14_u1_n100 ) , .ZN( u2_u14_u1_n135 ) , .A1( u2_u14_u1_n99 ) );
  AOI21_X1 u2_u14_u1_U53 (.A( u2_u14_u1_n152 ) , .B2( u2_u14_u1_n153 ) , .B1( u2_u14_u1_n154 ) , .ZN( u2_u14_u1_n158 ) );
  INV_X1 u2_u14_u1_U54 (.A( u2_u14_u1_n160 ) , .ZN( u2_u14_u1_n175 ) );
  NAND2_X1 u2_u14_u1_U55 (.A1( u2_u14_u1_n100 ) , .ZN( u2_u14_u1_n116 ) , .A2( u2_u14_u1_n95 ) );
  NAND2_X1 u2_u14_u1_U56 (.A1( u2_u14_u1_n102 ) , .ZN( u2_u14_u1_n131 ) , .A2( u2_u14_u1_n95 ) );
  NAND2_X1 u2_u14_u1_U57 (.A2( u2_u14_u1_n104 ) , .ZN( u2_u14_u1_n121 ) , .A1( u2_u14_u1_n98 ) );
  NAND2_X1 u2_u14_u1_U58 (.A1( u2_u14_u1_n103 ) , .ZN( u2_u14_u1_n153 ) , .A2( u2_u14_u1_n98 ) );
  NAND2_X1 u2_u14_u1_U59 (.A2( u2_u14_u1_n104 ) , .A1( u2_u14_u1_n105 ) , .ZN( u2_u14_u1_n133 ) );
  NOR2_X1 u2_u14_u1_U6 (.A1( u2_u14_u1_n112 ) , .A2( u2_u14_u1_n116 ) , .ZN( u2_u14_u1_n118 ) );
  NAND2_X1 u2_u14_u1_U60 (.ZN( u2_u14_u1_n150 ) , .A2( u2_u14_u1_n98 ) , .A1( u2_u14_u1_n99 ) );
  NAND2_X1 u2_u14_u1_U61 (.A1( u2_u14_u1_n105 ) , .ZN( u2_u14_u1_n155 ) , .A2( u2_u14_u1_n95 ) );
  OAI21_X1 u2_u14_u1_U62 (.ZN( u2_u14_u1_n109 ) , .B1( u2_u14_u1_n129 ) , .B2( u2_u14_u1_n160 ) , .A( u2_u14_u1_n167 ) );
  NAND2_X1 u2_u14_u1_U63 (.A2( u2_u14_u1_n100 ) , .A1( u2_u14_u1_n103 ) , .ZN( u2_u14_u1_n120 ) );
  NAND2_X1 u2_u14_u1_U64 (.A1( u2_u14_u1_n102 ) , .A2( u2_u14_u1_n104 ) , .ZN( u2_u14_u1_n115 ) );
  NAND2_X1 u2_u14_u1_U65 (.A2( u2_u14_u1_n100 ) , .A1( u2_u14_u1_n104 ) , .ZN( u2_u14_u1_n151 ) );
  NAND2_X1 u2_u14_u1_U66 (.A2( u2_u14_u1_n103 ) , .A1( u2_u14_u1_n105 ) , .ZN( u2_u14_u1_n161 ) );
  INV_X1 u2_u14_u1_U67 (.A( u2_u14_u1_n152 ) , .ZN( u2_u14_u1_n173 ) );
  INV_X1 u2_u14_u1_U68 (.A( u2_u14_u1_n128 ) , .ZN( u2_u14_u1_n172 ) );
  NAND2_X1 u2_u14_u1_U69 (.A2( u2_u14_u1_n102 ) , .A1( u2_u14_u1_n103 ) , .ZN( u2_u14_u1_n123 ) );
  OAI21_X1 u2_u14_u1_U7 (.ZN( u2_u14_u1_n101 ) , .B1( u2_u14_u1_n141 ) , .A( u2_u14_u1_n146 ) , .B2( u2_u14_u1_n183 ) );
  NOR2_X1 u2_u14_u1_U70 (.A2( u2_u14_X_7 ) , .A1( u2_u14_X_8 ) , .ZN( u2_u14_u1_n95 ) );
  NOR2_X1 u2_u14_u1_U71 (.A1( u2_u14_X_12 ) , .A2( u2_u14_X_9 ) , .ZN( u2_u14_u1_n100 ) );
  NOR2_X1 u2_u14_u1_U72 (.A2( u2_u14_X_8 ) , .A1( u2_u14_u1_n177 ) , .ZN( u2_u14_u1_n99 ) );
  NOR2_X1 u2_u14_u1_U73 (.A2( u2_u14_X_12 ) , .ZN( u2_u14_u1_n102 ) , .A1( u2_u14_u1_n176 ) );
  NOR2_X1 u2_u14_u1_U74 (.A2( u2_u14_X_9 ) , .ZN( u2_u14_u1_n105 ) , .A1( u2_u14_u1_n168 ) );
  NAND2_X1 u2_u14_u1_U75 (.A1( u2_u14_X_10 ) , .ZN( u2_u14_u1_n160 ) , .A2( u2_u14_u1_n169 ) );
  NAND2_X1 u2_u14_u1_U76 (.A2( u2_u14_X_10 ) , .A1( u2_u14_X_11 ) , .ZN( u2_u14_u1_n152 ) );
  NAND2_X1 u2_u14_u1_U77 (.A1( u2_u14_X_11 ) , .ZN( u2_u14_u1_n128 ) , .A2( u2_u14_u1_n170 ) );
  AND2_X1 u2_u14_u1_U78 (.A2( u2_u14_X_7 ) , .A1( u2_u14_X_8 ) , .ZN( u2_u14_u1_n104 ) );
  AND2_X1 u2_u14_u1_U79 (.A1( u2_u14_X_8 ) , .ZN( u2_u14_u1_n103 ) , .A2( u2_u14_u1_n177 ) );
  AOI21_X1 u2_u14_u1_U8 (.B2( u2_u14_u1_n155 ) , .B1( u2_u14_u1_n156 ) , .ZN( u2_u14_u1_n157 ) , .A( u2_u14_u1_n174 ) );
  INV_X1 u2_u14_u1_U80 (.A( u2_u14_X_10 ) , .ZN( u2_u14_u1_n170 ) );
  INV_X1 u2_u14_u1_U81 (.A( u2_u14_X_9 ) , .ZN( u2_u14_u1_n176 ) );
  INV_X1 u2_u14_u1_U82 (.A( u2_u14_X_11 ) , .ZN( u2_u14_u1_n169 ) );
  INV_X1 u2_u14_u1_U83 (.A( u2_u14_X_12 ) , .ZN( u2_u14_u1_n168 ) );
  INV_X1 u2_u14_u1_U84 (.A( u2_u14_X_7 ) , .ZN( u2_u14_u1_n177 ) );
  NAND4_X1 u2_u14_u1_U85 (.ZN( u2_out14_28 ) , .A4( u2_u14_u1_n124 ) , .A3( u2_u14_u1_n125 ) , .A2( u2_u14_u1_n126 ) , .A1( u2_u14_u1_n127 ) );
  OAI21_X1 u2_u14_u1_U86 (.ZN( u2_u14_u1_n127 ) , .B2( u2_u14_u1_n139 ) , .B1( u2_u14_u1_n175 ) , .A( u2_u14_u1_n183 ) );
  OAI21_X1 u2_u14_u1_U87 (.ZN( u2_u14_u1_n126 ) , .B2( u2_u14_u1_n140 ) , .A( u2_u14_u1_n146 ) , .B1( u2_u14_u1_n178 ) );
  NAND4_X1 u2_u14_u1_U88 (.ZN( u2_out14_18 ) , .A4( u2_u14_u1_n165 ) , .A3( u2_u14_u1_n166 ) , .A1( u2_u14_u1_n167 ) , .A2( u2_u14_u1_n186 ) );
  AOI22_X1 u2_u14_u1_U89 (.B2( u2_u14_u1_n146 ) , .B1( u2_u14_u1_n147 ) , .A2( u2_u14_u1_n148 ) , .ZN( u2_u14_u1_n166 ) , .A1( u2_u14_u1_n172 ) );
  OR4_X1 u2_u14_u1_U9 (.A4( u2_u14_u1_n106 ) , .A3( u2_u14_u1_n107 ) , .ZN( u2_u14_u1_n108 ) , .A1( u2_u14_u1_n117 ) , .A2( u2_u14_u1_n184 ) );
  INV_X1 u2_u14_u1_U90 (.A( u2_u14_u1_n145 ) , .ZN( u2_u14_u1_n186 ) );
  NAND4_X1 u2_u14_u1_U91 (.ZN( u2_out14_2 ) , .A4( u2_u14_u1_n142 ) , .A3( u2_u14_u1_n143 ) , .A2( u2_u14_u1_n144 ) , .A1( u2_u14_u1_n179 ) );
  OAI21_X1 u2_u14_u1_U92 (.B2( u2_u14_u1_n132 ) , .ZN( u2_u14_u1_n144 ) , .A( u2_u14_u1_n146 ) , .B1( u2_u14_u1_n180 ) );
  INV_X1 u2_u14_u1_U93 (.A( u2_u14_u1_n130 ) , .ZN( u2_u14_u1_n179 ) );
  OR4_X1 u2_u14_u1_U94 (.ZN( u2_out14_13 ) , .A4( u2_u14_u1_n108 ) , .A3( u2_u14_u1_n109 ) , .A2( u2_u14_u1_n110 ) , .A1( u2_u14_u1_n111 ) );
  AOI21_X1 u2_u14_u1_U95 (.ZN( u2_u14_u1_n111 ) , .A( u2_u14_u1_n128 ) , .B2( u2_u14_u1_n131 ) , .B1( u2_u14_u1_n135 ) );
  AOI21_X1 u2_u14_u1_U96 (.ZN( u2_u14_u1_n110 ) , .A( u2_u14_u1_n116 ) , .B1( u2_u14_u1_n152 ) , .B2( u2_u14_u1_n160 ) );
  NAND3_X1 u2_u14_u1_U97 (.A3( u2_u14_u1_n149 ) , .A2( u2_u14_u1_n150 ) , .A1( u2_u14_u1_n151 ) , .ZN( u2_u14_u1_n164 ) );
  NAND3_X1 u2_u14_u1_U98 (.A3( u2_u14_u1_n134 ) , .A2( u2_u14_u1_n135 ) , .ZN( u2_u14_u1_n136 ) , .A1( u2_u14_u1_n151 ) );
  NAND3_X1 u2_u14_u1_U99 (.A1( u2_u14_u1_n133 ) , .ZN( u2_u14_u1_n137 ) , .A2( u2_u14_u1_n154 ) , .A3( u2_u14_u1_n181 ) );
  OAI22_X1 u2_u14_u2_U10 (.ZN( u2_u14_u2_n109 ) , .A2( u2_u14_u2_n113 ) , .B2( u2_u14_u2_n133 ) , .B1( u2_u14_u2_n167 ) , .A1( u2_u14_u2_n168 ) );
  NAND3_X1 u2_u14_u2_U100 (.A2( u2_u14_u2_n100 ) , .A1( u2_u14_u2_n104 ) , .A3( u2_u14_u2_n138 ) , .ZN( u2_u14_u2_n98 ) );
  OAI22_X1 u2_u14_u2_U11 (.B1( u2_u14_u2_n151 ) , .A2( u2_u14_u2_n152 ) , .A1( u2_u14_u2_n153 ) , .ZN( u2_u14_u2_n160 ) , .B2( u2_u14_u2_n168 ) );
  NOR3_X1 u2_u14_u2_U12 (.A1( u2_u14_u2_n150 ) , .ZN( u2_u14_u2_n151 ) , .A3( u2_u14_u2_n175 ) , .A2( u2_u14_u2_n188 ) );
  AOI21_X1 u2_u14_u2_U13 (.ZN( u2_u14_u2_n144 ) , .B2( u2_u14_u2_n155 ) , .A( u2_u14_u2_n172 ) , .B1( u2_u14_u2_n185 ) );
  AOI21_X1 u2_u14_u2_U14 (.B2( u2_u14_u2_n143 ) , .ZN( u2_u14_u2_n145 ) , .B1( u2_u14_u2_n152 ) , .A( u2_u14_u2_n171 ) );
  AOI21_X1 u2_u14_u2_U15 (.B2( u2_u14_u2_n120 ) , .B1( u2_u14_u2_n121 ) , .ZN( u2_u14_u2_n126 ) , .A( u2_u14_u2_n167 ) );
  INV_X1 u2_u14_u2_U16 (.A( u2_u14_u2_n156 ) , .ZN( u2_u14_u2_n171 ) );
  INV_X1 u2_u14_u2_U17 (.A( u2_u14_u2_n120 ) , .ZN( u2_u14_u2_n188 ) );
  NAND2_X1 u2_u14_u2_U18 (.A2( u2_u14_u2_n122 ) , .ZN( u2_u14_u2_n150 ) , .A1( u2_u14_u2_n152 ) );
  INV_X1 u2_u14_u2_U19 (.A( u2_u14_u2_n153 ) , .ZN( u2_u14_u2_n170 ) );
  INV_X1 u2_u14_u2_U20 (.A( u2_u14_u2_n137 ) , .ZN( u2_u14_u2_n173 ) );
  NAND2_X1 u2_u14_u2_U21 (.A1( u2_u14_u2_n132 ) , .A2( u2_u14_u2_n139 ) , .ZN( u2_u14_u2_n157 ) );
  INV_X1 u2_u14_u2_U22 (.A( u2_u14_u2_n113 ) , .ZN( u2_u14_u2_n178 ) );
  INV_X1 u2_u14_u2_U23 (.A( u2_u14_u2_n139 ) , .ZN( u2_u14_u2_n175 ) );
  INV_X1 u2_u14_u2_U24 (.A( u2_u14_u2_n155 ) , .ZN( u2_u14_u2_n181 ) );
  INV_X1 u2_u14_u2_U25 (.A( u2_u14_u2_n119 ) , .ZN( u2_u14_u2_n177 ) );
  INV_X1 u2_u14_u2_U26 (.A( u2_u14_u2_n116 ) , .ZN( u2_u14_u2_n180 ) );
  INV_X1 u2_u14_u2_U27 (.A( u2_u14_u2_n131 ) , .ZN( u2_u14_u2_n179 ) );
  INV_X1 u2_u14_u2_U28 (.A( u2_u14_u2_n154 ) , .ZN( u2_u14_u2_n176 ) );
  NAND2_X1 u2_u14_u2_U29 (.A2( u2_u14_u2_n116 ) , .A1( u2_u14_u2_n117 ) , .ZN( u2_u14_u2_n118 ) );
  NOR2_X1 u2_u14_u2_U3 (.ZN( u2_u14_u2_n121 ) , .A2( u2_u14_u2_n177 ) , .A1( u2_u14_u2_n180 ) );
  INV_X1 u2_u14_u2_U30 (.A( u2_u14_u2_n132 ) , .ZN( u2_u14_u2_n182 ) );
  INV_X1 u2_u14_u2_U31 (.A( u2_u14_u2_n158 ) , .ZN( u2_u14_u2_n183 ) );
  OAI21_X1 u2_u14_u2_U32 (.A( u2_u14_u2_n156 ) , .B1( u2_u14_u2_n157 ) , .ZN( u2_u14_u2_n158 ) , .B2( u2_u14_u2_n179 ) );
  NOR2_X1 u2_u14_u2_U33 (.ZN( u2_u14_u2_n156 ) , .A1( u2_u14_u2_n166 ) , .A2( u2_u14_u2_n169 ) );
  NOR2_X1 u2_u14_u2_U34 (.A2( u2_u14_u2_n114 ) , .ZN( u2_u14_u2_n137 ) , .A1( u2_u14_u2_n140 ) );
  NOR2_X1 u2_u14_u2_U35 (.A2( u2_u14_u2_n138 ) , .ZN( u2_u14_u2_n153 ) , .A1( u2_u14_u2_n156 ) );
  AOI211_X1 u2_u14_u2_U36 (.ZN( u2_u14_u2_n130 ) , .C1( u2_u14_u2_n138 ) , .C2( u2_u14_u2_n179 ) , .B( u2_u14_u2_n96 ) , .A( u2_u14_u2_n97 ) );
  OAI22_X1 u2_u14_u2_U37 (.B1( u2_u14_u2_n133 ) , .A2( u2_u14_u2_n137 ) , .A1( u2_u14_u2_n152 ) , .B2( u2_u14_u2_n168 ) , .ZN( u2_u14_u2_n97 ) );
  OAI221_X1 u2_u14_u2_U38 (.B1( u2_u14_u2_n113 ) , .C1( u2_u14_u2_n132 ) , .A( u2_u14_u2_n149 ) , .B2( u2_u14_u2_n171 ) , .C2( u2_u14_u2_n172 ) , .ZN( u2_u14_u2_n96 ) );
  OAI221_X1 u2_u14_u2_U39 (.A( u2_u14_u2_n115 ) , .C2( u2_u14_u2_n123 ) , .B2( u2_u14_u2_n143 ) , .B1( u2_u14_u2_n153 ) , .ZN( u2_u14_u2_n163 ) , .C1( u2_u14_u2_n168 ) );
  INV_X1 u2_u14_u2_U4 (.A( u2_u14_u2_n134 ) , .ZN( u2_u14_u2_n185 ) );
  OAI21_X1 u2_u14_u2_U40 (.A( u2_u14_u2_n114 ) , .ZN( u2_u14_u2_n115 ) , .B1( u2_u14_u2_n176 ) , .B2( u2_u14_u2_n178 ) );
  OAI221_X1 u2_u14_u2_U41 (.A( u2_u14_u2_n135 ) , .B2( u2_u14_u2_n136 ) , .B1( u2_u14_u2_n137 ) , .ZN( u2_u14_u2_n162 ) , .C2( u2_u14_u2_n167 ) , .C1( u2_u14_u2_n185 ) );
  AND3_X1 u2_u14_u2_U42 (.A3( u2_u14_u2_n131 ) , .A2( u2_u14_u2_n132 ) , .A1( u2_u14_u2_n133 ) , .ZN( u2_u14_u2_n136 ) );
  AOI22_X1 u2_u14_u2_U43 (.ZN( u2_u14_u2_n135 ) , .B1( u2_u14_u2_n140 ) , .A1( u2_u14_u2_n156 ) , .B2( u2_u14_u2_n180 ) , .A2( u2_u14_u2_n188 ) );
  AOI21_X1 u2_u14_u2_U44 (.ZN( u2_u14_u2_n149 ) , .B1( u2_u14_u2_n173 ) , .B2( u2_u14_u2_n188 ) , .A( u2_u14_u2_n95 ) );
  AND3_X1 u2_u14_u2_U45 (.A2( u2_u14_u2_n100 ) , .A1( u2_u14_u2_n104 ) , .A3( u2_u14_u2_n156 ) , .ZN( u2_u14_u2_n95 ) );
  OAI21_X1 u2_u14_u2_U46 (.A( u2_u14_u2_n141 ) , .B2( u2_u14_u2_n142 ) , .ZN( u2_u14_u2_n146 ) , .B1( u2_u14_u2_n153 ) );
  OAI21_X1 u2_u14_u2_U47 (.A( u2_u14_u2_n140 ) , .ZN( u2_u14_u2_n141 ) , .B1( u2_u14_u2_n176 ) , .B2( u2_u14_u2_n177 ) );
  NOR3_X1 u2_u14_u2_U48 (.ZN( u2_u14_u2_n142 ) , .A3( u2_u14_u2_n175 ) , .A2( u2_u14_u2_n178 ) , .A1( u2_u14_u2_n181 ) );
  OAI21_X1 u2_u14_u2_U49 (.A( u2_u14_u2_n101 ) , .B2( u2_u14_u2_n121 ) , .B1( u2_u14_u2_n153 ) , .ZN( u2_u14_u2_n164 ) );
  INV_X1 u2_u14_u2_U5 (.A( u2_u14_u2_n150 ) , .ZN( u2_u14_u2_n184 ) );
  NAND2_X1 u2_u14_u2_U50 (.A2( u2_u14_u2_n100 ) , .A1( u2_u14_u2_n107 ) , .ZN( u2_u14_u2_n155 ) );
  NAND2_X1 u2_u14_u2_U51 (.A2( u2_u14_u2_n105 ) , .A1( u2_u14_u2_n108 ) , .ZN( u2_u14_u2_n143 ) );
  NAND2_X1 u2_u14_u2_U52 (.A1( u2_u14_u2_n104 ) , .A2( u2_u14_u2_n106 ) , .ZN( u2_u14_u2_n152 ) );
  NAND2_X1 u2_u14_u2_U53 (.A1( u2_u14_u2_n100 ) , .A2( u2_u14_u2_n105 ) , .ZN( u2_u14_u2_n132 ) );
  INV_X1 u2_u14_u2_U54 (.A( u2_u14_u2_n140 ) , .ZN( u2_u14_u2_n168 ) );
  INV_X1 u2_u14_u2_U55 (.A( u2_u14_u2_n138 ) , .ZN( u2_u14_u2_n167 ) );
  INV_X1 u2_u14_u2_U56 (.ZN( u2_u14_u2_n187 ) , .A( u2_u14_u2_n99 ) );
  OAI21_X1 u2_u14_u2_U57 (.B1( u2_u14_u2_n137 ) , .B2( u2_u14_u2_n143 ) , .A( u2_u14_u2_n98 ) , .ZN( u2_u14_u2_n99 ) );
  NAND2_X1 u2_u14_u2_U58 (.A1( u2_u14_u2_n102 ) , .A2( u2_u14_u2_n106 ) , .ZN( u2_u14_u2_n113 ) );
  NAND2_X1 u2_u14_u2_U59 (.A1( u2_u14_u2_n106 ) , .A2( u2_u14_u2_n107 ) , .ZN( u2_u14_u2_n131 ) );
  NOR4_X1 u2_u14_u2_U6 (.A4( u2_u14_u2_n124 ) , .A3( u2_u14_u2_n125 ) , .A2( u2_u14_u2_n126 ) , .A1( u2_u14_u2_n127 ) , .ZN( u2_u14_u2_n128 ) );
  NAND2_X1 u2_u14_u2_U60 (.A1( u2_u14_u2_n103 ) , .A2( u2_u14_u2_n107 ) , .ZN( u2_u14_u2_n139 ) );
  NAND2_X1 u2_u14_u2_U61 (.A1( u2_u14_u2_n103 ) , .A2( u2_u14_u2_n105 ) , .ZN( u2_u14_u2_n133 ) );
  NAND2_X1 u2_u14_u2_U62 (.A1( u2_u14_u2_n102 ) , .A2( u2_u14_u2_n103 ) , .ZN( u2_u14_u2_n154 ) );
  NAND2_X1 u2_u14_u2_U63 (.A2( u2_u14_u2_n103 ) , .A1( u2_u14_u2_n104 ) , .ZN( u2_u14_u2_n119 ) );
  NAND2_X1 u2_u14_u2_U64 (.A2( u2_u14_u2_n107 ) , .A1( u2_u14_u2_n108 ) , .ZN( u2_u14_u2_n123 ) );
  NAND2_X1 u2_u14_u2_U65 (.A1( u2_u14_u2_n104 ) , .A2( u2_u14_u2_n108 ) , .ZN( u2_u14_u2_n122 ) );
  INV_X1 u2_u14_u2_U66 (.A( u2_u14_u2_n114 ) , .ZN( u2_u14_u2_n172 ) );
  NAND2_X1 u2_u14_u2_U67 (.A2( u2_u14_u2_n100 ) , .A1( u2_u14_u2_n102 ) , .ZN( u2_u14_u2_n116 ) );
  NAND2_X1 u2_u14_u2_U68 (.A1( u2_u14_u2_n102 ) , .A2( u2_u14_u2_n108 ) , .ZN( u2_u14_u2_n120 ) );
  NAND2_X1 u2_u14_u2_U69 (.A2( u2_u14_u2_n105 ) , .A1( u2_u14_u2_n106 ) , .ZN( u2_u14_u2_n117 ) );
  AOI21_X1 u2_u14_u2_U7 (.B2( u2_u14_u2_n119 ) , .ZN( u2_u14_u2_n127 ) , .A( u2_u14_u2_n137 ) , .B1( u2_u14_u2_n155 ) );
  NOR2_X1 u2_u14_u2_U70 (.A2( u2_u14_X_16 ) , .ZN( u2_u14_u2_n140 ) , .A1( u2_u14_u2_n166 ) );
  NOR2_X1 u2_u14_u2_U71 (.A2( u2_u14_X_13 ) , .A1( u2_u14_X_14 ) , .ZN( u2_u14_u2_n100 ) );
  NOR2_X1 u2_u14_u2_U72 (.A2( u2_u14_X_16 ) , .A1( u2_u14_X_17 ) , .ZN( u2_u14_u2_n138 ) );
  NOR2_X1 u2_u14_u2_U73 (.A2( u2_u14_X_15 ) , .A1( u2_u14_X_18 ) , .ZN( u2_u14_u2_n104 ) );
  NOR2_X1 u2_u14_u2_U74 (.A2( u2_u14_X_14 ) , .ZN( u2_u14_u2_n103 ) , .A1( u2_u14_u2_n174 ) );
  NOR2_X1 u2_u14_u2_U75 (.A2( u2_u14_X_15 ) , .ZN( u2_u14_u2_n102 ) , .A1( u2_u14_u2_n165 ) );
  NOR2_X1 u2_u14_u2_U76 (.A2( u2_u14_X_17 ) , .ZN( u2_u14_u2_n114 ) , .A1( u2_u14_u2_n169 ) );
  AND2_X1 u2_u14_u2_U77 (.A1( u2_u14_X_15 ) , .ZN( u2_u14_u2_n105 ) , .A2( u2_u14_u2_n165 ) );
  AND2_X1 u2_u14_u2_U78 (.A2( u2_u14_X_15 ) , .A1( u2_u14_X_18 ) , .ZN( u2_u14_u2_n107 ) );
  AND2_X1 u2_u14_u2_U79 (.A1( u2_u14_X_14 ) , .ZN( u2_u14_u2_n106 ) , .A2( u2_u14_u2_n174 ) );
  AOI21_X1 u2_u14_u2_U8 (.ZN( u2_u14_u2_n124 ) , .B1( u2_u14_u2_n131 ) , .B2( u2_u14_u2_n143 ) , .A( u2_u14_u2_n172 ) );
  AND2_X1 u2_u14_u2_U80 (.A1( u2_u14_X_13 ) , .A2( u2_u14_X_14 ) , .ZN( u2_u14_u2_n108 ) );
  INV_X1 u2_u14_u2_U81 (.A( u2_u14_X_16 ) , .ZN( u2_u14_u2_n169 ) );
  INV_X1 u2_u14_u2_U82 (.A( u2_u14_X_17 ) , .ZN( u2_u14_u2_n166 ) );
  INV_X1 u2_u14_u2_U83 (.A( u2_u14_X_13 ) , .ZN( u2_u14_u2_n174 ) );
  INV_X1 u2_u14_u2_U84 (.A( u2_u14_X_18 ) , .ZN( u2_u14_u2_n165 ) );
  NAND4_X1 u2_u14_u2_U85 (.ZN( u2_out14_30 ) , .A4( u2_u14_u2_n147 ) , .A3( u2_u14_u2_n148 ) , .A2( u2_u14_u2_n149 ) , .A1( u2_u14_u2_n187 ) );
  NOR3_X1 u2_u14_u2_U86 (.A3( u2_u14_u2_n144 ) , .A2( u2_u14_u2_n145 ) , .A1( u2_u14_u2_n146 ) , .ZN( u2_u14_u2_n147 ) );
  AOI21_X1 u2_u14_u2_U87 (.B2( u2_u14_u2_n138 ) , .ZN( u2_u14_u2_n148 ) , .A( u2_u14_u2_n162 ) , .B1( u2_u14_u2_n182 ) );
  NAND4_X1 u2_u14_u2_U88 (.ZN( u2_out14_24 ) , .A4( u2_u14_u2_n111 ) , .A3( u2_u14_u2_n112 ) , .A1( u2_u14_u2_n130 ) , .A2( u2_u14_u2_n187 ) );
  AOI221_X1 u2_u14_u2_U89 (.A( u2_u14_u2_n109 ) , .B1( u2_u14_u2_n110 ) , .ZN( u2_u14_u2_n111 ) , .C1( u2_u14_u2_n134 ) , .C2( u2_u14_u2_n170 ) , .B2( u2_u14_u2_n173 ) );
  AOI21_X1 u2_u14_u2_U9 (.B2( u2_u14_u2_n123 ) , .ZN( u2_u14_u2_n125 ) , .A( u2_u14_u2_n171 ) , .B1( u2_u14_u2_n184 ) );
  AOI21_X1 u2_u14_u2_U90 (.ZN( u2_u14_u2_n112 ) , .B2( u2_u14_u2_n156 ) , .A( u2_u14_u2_n164 ) , .B1( u2_u14_u2_n181 ) );
  NAND4_X1 u2_u14_u2_U91 (.ZN( u2_out14_16 ) , .A4( u2_u14_u2_n128 ) , .A3( u2_u14_u2_n129 ) , .A1( u2_u14_u2_n130 ) , .A2( u2_u14_u2_n186 ) );
  AOI22_X1 u2_u14_u2_U92 (.A2( u2_u14_u2_n118 ) , .ZN( u2_u14_u2_n129 ) , .A1( u2_u14_u2_n140 ) , .B1( u2_u14_u2_n157 ) , .B2( u2_u14_u2_n170 ) );
  INV_X1 u2_u14_u2_U93 (.A( u2_u14_u2_n163 ) , .ZN( u2_u14_u2_n186 ) );
  OR4_X1 u2_u14_u2_U94 (.ZN( u2_out14_6 ) , .A4( u2_u14_u2_n161 ) , .A3( u2_u14_u2_n162 ) , .A2( u2_u14_u2_n163 ) , .A1( u2_u14_u2_n164 ) );
  OR3_X1 u2_u14_u2_U95 (.A2( u2_u14_u2_n159 ) , .A1( u2_u14_u2_n160 ) , .ZN( u2_u14_u2_n161 ) , .A3( u2_u14_u2_n183 ) );
  AOI21_X1 u2_u14_u2_U96 (.B2( u2_u14_u2_n154 ) , .B1( u2_u14_u2_n155 ) , .ZN( u2_u14_u2_n159 ) , .A( u2_u14_u2_n167 ) );
  NAND3_X1 u2_u14_u2_U97 (.A2( u2_u14_u2_n117 ) , .A1( u2_u14_u2_n122 ) , .A3( u2_u14_u2_n123 ) , .ZN( u2_u14_u2_n134 ) );
  NAND3_X1 u2_u14_u2_U98 (.ZN( u2_u14_u2_n110 ) , .A2( u2_u14_u2_n131 ) , .A3( u2_u14_u2_n139 ) , .A1( u2_u14_u2_n154 ) );
  NAND3_X1 u2_u14_u2_U99 (.A2( u2_u14_u2_n100 ) , .ZN( u2_u14_u2_n101 ) , .A1( u2_u14_u2_n104 ) , .A3( u2_u14_u2_n114 ) );
  OAI22_X1 u2_u14_u3_U10 (.B1( u2_u14_u3_n113 ) , .A2( u2_u14_u3_n135 ) , .A1( u2_u14_u3_n150 ) , .B2( u2_u14_u3_n164 ) , .ZN( u2_u14_u3_n98 ) );
  OAI211_X1 u2_u14_u3_U11 (.B( u2_u14_u3_n106 ) , .ZN( u2_u14_u3_n119 ) , .C2( u2_u14_u3_n128 ) , .C1( u2_u14_u3_n167 ) , .A( u2_u14_u3_n181 ) );
  AOI221_X1 u2_u14_u3_U12 (.C1( u2_u14_u3_n105 ) , .ZN( u2_u14_u3_n106 ) , .A( u2_u14_u3_n131 ) , .B2( u2_u14_u3_n132 ) , .C2( u2_u14_u3_n133 ) , .B1( u2_u14_u3_n169 ) );
  INV_X1 u2_u14_u3_U13 (.ZN( u2_u14_u3_n181 ) , .A( u2_u14_u3_n98 ) );
  NAND2_X1 u2_u14_u3_U14 (.ZN( u2_u14_u3_n105 ) , .A2( u2_u14_u3_n130 ) , .A1( u2_u14_u3_n155 ) );
  AOI22_X1 u2_u14_u3_U15 (.B1( u2_u14_u3_n115 ) , .A2( u2_u14_u3_n116 ) , .ZN( u2_u14_u3_n123 ) , .B2( u2_u14_u3_n133 ) , .A1( u2_u14_u3_n169 ) );
  NAND2_X1 u2_u14_u3_U16 (.ZN( u2_u14_u3_n116 ) , .A2( u2_u14_u3_n151 ) , .A1( u2_u14_u3_n182 ) );
  NOR2_X1 u2_u14_u3_U17 (.ZN( u2_u14_u3_n126 ) , .A2( u2_u14_u3_n150 ) , .A1( u2_u14_u3_n164 ) );
  AOI21_X1 u2_u14_u3_U18 (.ZN( u2_u14_u3_n112 ) , .B2( u2_u14_u3_n146 ) , .B1( u2_u14_u3_n155 ) , .A( u2_u14_u3_n167 ) );
  NAND2_X1 u2_u14_u3_U19 (.A1( u2_u14_u3_n135 ) , .ZN( u2_u14_u3_n142 ) , .A2( u2_u14_u3_n164 ) );
  NAND2_X1 u2_u14_u3_U20 (.ZN( u2_u14_u3_n132 ) , .A2( u2_u14_u3_n152 ) , .A1( u2_u14_u3_n156 ) );
  AND2_X1 u2_u14_u3_U21 (.A2( u2_u14_u3_n113 ) , .A1( u2_u14_u3_n114 ) , .ZN( u2_u14_u3_n151 ) );
  INV_X1 u2_u14_u3_U22 (.A( u2_u14_u3_n133 ) , .ZN( u2_u14_u3_n165 ) );
  INV_X1 u2_u14_u3_U23 (.A( u2_u14_u3_n135 ) , .ZN( u2_u14_u3_n170 ) );
  NAND2_X1 u2_u14_u3_U24 (.A1( u2_u14_u3_n107 ) , .A2( u2_u14_u3_n108 ) , .ZN( u2_u14_u3_n140 ) );
  NAND2_X1 u2_u14_u3_U25 (.ZN( u2_u14_u3_n117 ) , .A1( u2_u14_u3_n124 ) , .A2( u2_u14_u3_n148 ) );
  NAND2_X1 u2_u14_u3_U26 (.ZN( u2_u14_u3_n143 ) , .A1( u2_u14_u3_n165 ) , .A2( u2_u14_u3_n167 ) );
  INV_X1 u2_u14_u3_U27 (.A( u2_u14_u3_n130 ) , .ZN( u2_u14_u3_n177 ) );
  INV_X1 u2_u14_u3_U28 (.A( u2_u14_u3_n128 ) , .ZN( u2_u14_u3_n176 ) );
  INV_X1 u2_u14_u3_U29 (.A( u2_u14_u3_n155 ) , .ZN( u2_u14_u3_n174 ) );
  INV_X1 u2_u14_u3_U3 (.A( u2_u14_u3_n129 ) , .ZN( u2_u14_u3_n183 ) );
  INV_X1 u2_u14_u3_U30 (.A( u2_u14_u3_n139 ) , .ZN( u2_u14_u3_n185 ) );
  NOR2_X1 u2_u14_u3_U31 (.ZN( u2_u14_u3_n135 ) , .A2( u2_u14_u3_n141 ) , .A1( u2_u14_u3_n169 ) );
  OAI222_X1 u2_u14_u3_U32 (.C2( u2_u14_u3_n107 ) , .A2( u2_u14_u3_n108 ) , .B1( u2_u14_u3_n135 ) , .ZN( u2_u14_u3_n138 ) , .B2( u2_u14_u3_n146 ) , .C1( u2_u14_u3_n154 ) , .A1( u2_u14_u3_n164 ) );
  NOR4_X1 u2_u14_u3_U33 (.A4( u2_u14_u3_n157 ) , .A3( u2_u14_u3_n158 ) , .A2( u2_u14_u3_n159 ) , .A1( u2_u14_u3_n160 ) , .ZN( u2_u14_u3_n161 ) );
  AOI21_X1 u2_u14_u3_U34 (.B2( u2_u14_u3_n152 ) , .B1( u2_u14_u3_n153 ) , .ZN( u2_u14_u3_n158 ) , .A( u2_u14_u3_n164 ) );
  AOI21_X1 u2_u14_u3_U35 (.A( u2_u14_u3_n154 ) , .B2( u2_u14_u3_n155 ) , .B1( u2_u14_u3_n156 ) , .ZN( u2_u14_u3_n157 ) );
  AOI21_X1 u2_u14_u3_U36 (.A( u2_u14_u3_n149 ) , .B2( u2_u14_u3_n150 ) , .B1( u2_u14_u3_n151 ) , .ZN( u2_u14_u3_n159 ) );
  AOI211_X1 u2_u14_u3_U37 (.ZN( u2_u14_u3_n109 ) , .A( u2_u14_u3_n119 ) , .C2( u2_u14_u3_n129 ) , .B( u2_u14_u3_n138 ) , .C1( u2_u14_u3_n141 ) );
  AOI211_X1 u2_u14_u3_U38 (.B( u2_u14_u3_n119 ) , .A( u2_u14_u3_n120 ) , .C2( u2_u14_u3_n121 ) , .ZN( u2_u14_u3_n122 ) , .C1( u2_u14_u3_n179 ) );
  INV_X1 u2_u14_u3_U39 (.A( u2_u14_u3_n156 ) , .ZN( u2_u14_u3_n179 ) );
  INV_X1 u2_u14_u3_U4 (.A( u2_u14_u3_n140 ) , .ZN( u2_u14_u3_n182 ) );
  OAI22_X1 u2_u14_u3_U40 (.B1( u2_u14_u3_n118 ) , .ZN( u2_u14_u3_n120 ) , .A1( u2_u14_u3_n135 ) , .B2( u2_u14_u3_n154 ) , .A2( u2_u14_u3_n178 ) );
  AND3_X1 u2_u14_u3_U41 (.ZN( u2_u14_u3_n118 ) , .A2( u2_u14_u3_n124 ) , .A1( u2_u14_u3_n144 ) , .A3( u2_u14_u3_n152 ) );
  INV_X1 u2_u14_u3_U42 (.A( u2_u14_u3_n121 ) , .ZN( u2_u14_u3_n164 ) );
  NAND2_X1 u2_u14_u3_U43 (.ZN( u2_u14_u3_n133 ) , .A1( u2_u14_u3_n154 ) , .A2( u2_u14_u3_n164 ) );
  OAI211_X1 u2_u14_u3_U44 (.B( u2_u14_u3_n127 ) , .ZN( u2_u14_u3_n139 ) , .C1( u2_u14_u3_n150 ) , .C2( u2_u14_u3_n154 ) , .A( u2_u14_u3_n184 ) );
  INV_X1 u2_u14_u3_U45 (.A( u2_u14_u3_n125 ) , .ZN( u2_u14_u3_n184 ) );
  AOI221_X1 u2_u14_u3_U46 (.A( u2_u14_u3_n126 ) , .ZN( u2_u14_u3_n127 ) , .C2( u2_u14_u3_n132 ) , .C1( u2_u14_u3_n169 ) , .B2( u2_u14_u3_n170 ) , .B1( u2_u14_u3_n174 ) );
  OAI22_X1 u2_u14_u3_U47 (.A1( u2_u14_u3_n124 ) , .ZN( u2_u14_u3_n125 ) , .B2( u2_u14_u3_n145 ) , .A2( u2_u14_u3_n165 ) , .B1( u2_u14_u3_n167 ) );
  NOR2_X1 u2_u14_u3_U48 (.A1( u2_u14_u3_n113 ) , .ZN( u2_u14_u3_n131 ) , .A2( u2_u14_u3_n154 ) );
  NAND2_X1 u2_u14_u3_U49 (.A1( u2_u14_u3_n103 ) , .ZN( u2_u14_u3_n150 ) , .A2( u2_u14_u3_n99 ) );
  INV_X1 u2_u14_u3_U5 (.A( u2_u14_u3_n117 ) , .ZN( u2_u14_u3_n178 ) );
  NAND2_X1 u2_u14_u3_U50 (.A2( u2_u14_u3_n102 ) , .ZN( u2_u14_u3_n155 ) , .A1( u2_u14_u3_n97 ) );
  INV_X1 u2_u14_u3_U51 (.A( u2_u14_u3_n141 ) , .ZN( u2_u14_u3_n167 ) );
  AOI21_X1 u2_u14_u3_U52 (.B2( u2_u14_u3_n114 ) , .B1( u2_u14_u3_n146 ) , .A( u2_u14_u3_n154 ) , .ZN( u2_u14_u3_n94 ) );
  AOI21_X1 u2_u14_u3_U53 (.ZN( u2_u14_u3_n110 ) , .B2( u2_u14_u3_n142 ) , .B1( u2_u14_u3_n186 ) , .A( u2_u14_u3_n95 ) );
  INV_X1 u2_u14_u3_U54 (.A( u2_u14_u3_n145 ) , .ZN( u2_u14_u3_n186 ) );
  AOI21_X1 u2_u14_u3_U55 (.B1( u2_u14_u3_n124 ) , .A( u2_u14_u3_n149 ) , .B2( u2_u14_u3_n155 ) , .ZN( u2_u14_u3_n95 ) );
  INV_X1 u2_u14_u3_U56 (.A( u2_u14_u3_n149 ) , .ZN( u2_u14_u3_n169 ) );
  NAND2_X1 u2_u14_u3_U57 (.ZN( u2_u14_u3_n124 ) , .A1( u2_u14_u3_n96 ) , .A2( u2_u14_u3_n97 ) );
  NAND2_X1 u2_u14_u3_U58 (.A2( u2_u14_u3_n100 ) , .ZN( u2_u14_u3_n146 ) , .A1( u2_u14_u3_n96 ) );
  NAND2_X1 u2_u14_u3_U59 (.A1( u2_u14_u3_n101 ) , .ZN( u2_u14_u3_n145 ) , .A2( u2_u14_u3_n99 ) );
  AOI221_X1 u2_u14_u3_U6 (.A( u2_u14_u3_n131 ) , .C2( u2_u14_u3_n132 ) , .C1( u2_u14_u3_n133 ) , .ZN( u2_u14_u3_n134 ) , .B1( u2_u14_u3_n143 ) , .B2( u2_u14_u3_n177 ) );
  NAND2_X1 u2_u14_u3_U60 (.A1( u2_u14_u3_n100 ) , .ZN( u2_u14_u3_n156 ) , .A2( u2_u14_u3_n99 ) );
  NAND2_X1 u2_u14_u3_U61 (.A2( u2_u14_u3_n101 ) , .A1( u2_u14_u3_n104 ) , .ZN( u2_u14_u3_n148 ) );
  NAND2_X1 u2_u14_u3_U62 (.A1( u2_u14_u3_n100 ) , .A2( u2_u14_u3_n102 ) , .ZN( u2_u14_u3_n128 ) );
  NAND2_X1 u2_u14_u3_U63 (.A2( u2_u14_u3_n101 ) , .A1( u2_u14_u3_n102 ) , .ZN( u2_u14_u3_n152 ) );
  NAND2_X1 u2_u14_u3_U64 (.A2( u2_u14_u3_n101 ) , .ZN( u2_u14_u3_n114 ) , .A1( u2_u14_u3_n96 ) );
  NAND2_X1 u2_u14_u3_U65 (.ZN( u2_u14_u3_n107 ) , .A1( u2_u14_u3_n97 ) , .A2( u2_u14_u3_n99 ) );
  NAND2_X1 u2_u14_u3_U66 (.A2( u2_u14_u3_n100 ) , .A1( u2_u14_u3_n104 ) , .ZN( u2_u14_u3_n113 ) );
  NAND2_X1 u2_u14_u3_U67 (.A1( u2_u14_u3_n104 ) , .ZN( u2_u14_u3_n153 ) , .A2( u2_u14_u3_n97 ) );
  NAND2_X1 u2_u14_u3_U68 (.A2( u2_u14_u3_n103 ) , .A1( u2_u14_u3_n104 ) , .ZN( u2_u14_u3_n130 ) );
  NAND2_X1 u2_u14_u3_U69 (.A2( u2_u14_u3_n103 ) , .ZN( u2_u14_u3_n144 ) , .A1( u2_u14_u3_n96 ) );
  OAI22_X1 u2_u14_u3_U7 (.B2( u2_u14_u3_n147 ) , .A2( u2_u14_u3_n148 ) , .ZN( u2_u14_u3_n160 ) , .B1( u2_u14_u3_n165 ) , .A1( u2_u14_u3_n168 ) );
  NAND2_X1 u2_u14_u3_U70 (.A1( u2_u14_u3_n102 ) , .A2( u2_u14_u3_n103 ) , .ZN( u2_u14_u3_n108 ) );
  NOR2_X1 u2_u14_u3_U71 (.A2( u2_u14_X_19 ) , .A1( u2_u14_X_20 ) , .ZN( u2_u14_u3_n99 ) );
  NOR2_X1 u2_u14_u3_U72 (.A2( u2_u14_X_21 ) , .A1( u2_u14_X_24 ) , .ZN( u2_u14_u3_n103 ) );
  NOR2_X1 u2_u14_u3_U73 (.A2( u2_u14_X_24 ) , .A1( u2_u14_u3_n171 ) , .ZN( u2_u14_u3_n97 ) );
  NOR2_X1 u2_u14_u3_U74 (.A2( u2_u14_X_23 ) , .ZN( u2_u14_u3_n141 ) , .A1( u2_u14_u3_n166 ) );
  NOR2_X1 u2_u14_u3_U75 (.A2( u2_u14_X_19 ) , .A1( u2_u14_u3_n172 ) , .ZN( u2_u14_u3_n96 ) );
  NAND2_X1 u2_u14_u3_U76 (.A1( u2_u14_X_22 ) , .A2( u2_u14_X_23 ) , .ZN( u2_u14_u3_n154 ) );
  NAND2_X1 u2_u14_u3_U77 (.A1( u2_u14_X_23 ) , .ZN( u2_u14_u3_n149 ) , .A2( u2_u14_u3_n166 ) );
  NOR2_X1 u2_u14_u3_U78 (.A2( u2_u14_X_22 ) , .A1( u2_u14_X_23 ) , .ZN( u2_u14_u3_n121 ) );
  AND2_X1 u2_u14_u3_U79 (.A1( u2_u14_X_24 ) , .ZN( u2_u14_u3_n101 ) , .A2( u2_u14_u3_n171 ) );
  AND3_X1 u2_u14_u3_U8 (.A3( u2_u14_u3_n144 ) , .A2( u2_u14_u3_n145 ) , .A1( u2_u14_u3_n146 ) , .ZN( u2_u14_u3_n147 ) );
  AND2_X1 u2_u14_u3_U80 (.A1( u2_u14_X_19 ) , .ZN( u2_u14_u3_n102 ) , .A2( u2_u14_u3_n172 ) );
  AND2_X1 u2_u14_u3_U81 (.A1( u2_u14_X_21 ) , .A2( u2_u14_X_24 ) , .ZN( u2_u14_u3_n100 ) );
  AND2_X1 u2_u14_u3_U82 (.A2( u2_u14_X_19 ) , .A1( u2_u14_X_20 ) , .ZN( u2_u14_u3_n104 ) );
  INV_X1 u2_u14_u3_U83 (.A( u2_u14_X_22 ) , .ZN( u2_u14_u3_n166 ) );
  INV_X1 u2_u14_u3_U84 (.A( u2_u14_X_21 ) , .ZN( u2_u14_u3_n171 ) );
  INV_X1 u2_u14_u3_U85 (.A( u2_u14_X_20 ) , .ZN( u2_u14_u3_n172 ) );
  NAND4_X1 u2_u14_u3_U86 (.ZN( u2_out14_26 ) , .A4( u2_u14_u3_n109 ) , .A3( u2_u14_u3_n110 ) , .A2( u2_u14_u3_n111 ) , .A1( u2_u14_u3_n173 ) );
  INV_X1 u2_u14_u3_U87 (.ZN( u2_u14_u3_n173 ) , .A( u2_u14_u3_n94 ) );
  OAI21_X1 u2_u14_u3_U88 (.ZN( u2_u14_u3_n111 ) , .B2( u2_u14_u3_n117 ) , .A( u2_u14_u3_n133 ) , .B1( u2_u14_u3_n176 ) );
  NAND4_X1 u2_u14_u3_U89 (.ZN( u2_out14_20 ) , .A4( u2_u14_u3_n122 ) , .A3( u2_u14_u3_n123 ) , .A1( u2_u14_u3_n175 ) , .A2( u2_u14_u3_n180 ) );
  INV_X1 u2_u14_u3_U9 (.A( u2_u14_u3_n143 ) , .ZN( u2_u14_u3_n168 ) );
  INV_X1 u2_u14_u3_U90 (.A( u2_u14_u3_n126 ) , .ZN( u2_u14_u3_n180 ) );
  INV_X1 u2_u14_u3_U91 (.A( u2_u14_u3_n112 ) , .ZN( u2_u14_u3_n175 ) );
  NAND4_X1 u2_u14_u3_U92 (.ZN( u2_out14_1 ) , .A4( u2_u14_u3_n161 ) , .A3( u2_u14_u3_n162 ) , .A2( u2_u14_u3_n163 ) , .A1( u2_u14_u3_n185 ) );
  NAND2_X1 u2_u14_u3_U93 (.ZN( u2_u14_u3_n163 ) , .A2( u2_u14_u3_n170 ) , .A1( u2_u14_u3_n176 ) );
  AOI22_X1 u2_u14_u3_U94 (.B2( u2_u14_u3_n140 ) , .B1( u2_u14_u3_n141 ) , .A2( u2_u14_u3_n142 ) , .ZN( u2_u14_u3_n162 ) , .A1( u2_u14_u3_n177 ) );
  OR4_X1 u2_u14_u3_U95 (.ZN( u2_out14_10 ) , .A4( u2_u14_u3_n136 ) , .A3( u2_u14_u3_n137 ) , .A1( u2_u14_u3_n138 ) , .A2( u2_u14_u3_n139 ) );
  OAI222_X1 u2_u14_u3_U96 (.C1( u2_u14_u3_n128 ) , .ZN( u2_u14_u3_n137 ) , .B1( u2_u14_u3_n148 ) , .A2( u2_u14_u3_n150 ) , .B2( u2_u14_u3_n154 ) , .C2( u2_u14_u3_n164 ) , .A1( u2_u14_u3_n167 ) );
  OAI221_X1 u2_u14_u3_U97 (.A( u2_u14_u3_n134 ) , .B2( u2_u14_u3_n135 ) , .ZN( u2_u14_u3_n136 ) , .C1( u2_u14_u3_n149 ) , .B1( u2_u14_u3_n151 ) , .C2( u2_u14_u3_n183 ) );
  NAND3_X1 u2_u14_u3_U98 (.A1( u2_u14_u3_n114 ) , .ZN( u2_u14_u3_n115 ) , .A2( u2_u14_u3_n145 ) , .A3( u2_u14_u3_n153 ) );
  NAND3_X1 u2_u14_u3_U99 (.ZN( u2_u14_u3_n129 ) , .A2( u2_u14_u3_n144 ) , .A1( u2_u14_u3_n153 ) , .A3( u2_u14_u3_n182 ) );
  OAI22_X1 u2_u14_u4_U10 (.B2( u2_u14_u4_n135 ) , .ZN( u2_u14_u4_n137 ) , .B1( u2_u14_u4_n153 ) , .A1( u2_u14_u4_n155 ) , .A2( u2_u14_u4_n171 ) );
  AND3_X1 u2_u14_u4_U11 (.A2( u2_u14_u4_n134 ) , .ZN( u2_u14_u4_n135 ) , .A3( u2_u14_u4_n145 ) , .A1( u2_u14_u4_n157 ) );
  NAND2_X1 u2_u14_u4_U12 (.ZN( u2_u14_u4_n132 ) , .A2( u2_u14_u4_n170 ) , .A1( u2_u14_u4_n173 ) );
  AOI21_X1 u2_u14_u4_U13 (.B2( u2_u14_u4_n160 ) , .B1( u2_u14_u4_n161 ) , .ZN( u2_u14_u4_n162 ) , .A( u2_u14_u4_n170 ) );
  AOI21_X1 u2_u14_u4_U14 (.ZN( u2_u14_u4_n107 ) , .B2( u2_u14_u4_n143 ) , .A( u2_u14_u4_n174 ) , .B1( u2_u14_u4_n184 ) );
  AOI21_X1 u2_u14_u4_U15 (.B2( u2_u14_u4_n158 ) , .B1( u2_u14_u4_n159 ) , .ZN( u2_u14_u4_n163 ) , .A( u2_u14_u4_n174 ) );
  AOI21_X1 u2_u14_u4_U16 (.A( u2_u14_u4_n153 ) , .B2( u2_u14_u4_n154 ) , .B1( u2_u14_u4_n155 ) , .ZN( u2_u14_u4_n165 ) );
  AOI21_X1 u2_u14_u4_U17 (.A( u2_u14_u4_n156 ) , .B2( u2_u14_u4_n157 ) , .ZN( u2_u14_u4_n164 ) , .B1( u2_u14_u4_n184 ) );
  INV_X1 u2_u14_u4_U18 (.A( u2_u14_u4_n138 ) , .ZN( u2_u14_u4_n170 ) );
  AND2_X1 u2_u14_u4_U19 (.A2( u2_u14_u4_n120 ) , .ZN( u2_u14_u4_n155 ) , .A1( u2_u14_u4_n160 ) );
  INV_X1 u2_u14_u4_U20 (.A( u2_u14_u4_n156 ) , .ZN( u2_u14_u4_n175 ) );
  NAND2_X1 u2_u14_u4_U21 (.A2( u2_u14_u4_n118 ) , .ZN( u2_u14_u4_n131 ) , .A1( u2_u14_u4_n147 ) );
  NAND2_X1 u2_u14_u4_U22 (.A1( u2_u14_u4_n119 ) , .A2( u2_u14_u4_n120 ) , .ZN( u2_u14_u4_n130 ) );
  NAND2_X1 u2_u14_u4_U23 (.ZN( u2_u14_u4_n117 ) , .A2( u2_u14_u4_n118 ) , .A1( u2_u14_u4_n148 ) );
  NAND2_X1 u2_u14_u4_U24 (.ZN( u2_u14_u4_n129 ) , .A1( u2_u14_u4_n134 ) , .A2( u2_u14_u4_n148 ) );
  AND3_X1 u2_u14_u4_U25 (.A1( u2_u14_u4_n119 ) , .A2( u2_u14_u4_n143 ) , .A3( u2_u14_u4_n154 ) , .ZN( u2_u14_u4_n161 ) );
  AND2_X1 u2_u14_u4_U26 (.A1( u2_u14_u4_n145 ) , .A2( u2_u14_u4_n147 ) , .ZN( u2_u14_u4_n159 ) );
  OR3_X1 u2_u14_u4_U27 (.A3( u2_u14_u4_n114 ) , .A2( u2_u14_u4_n115 ) , .A1( u2_u14_u4_n116 ) , .ZN( u2_u14_u4_n136 ) );
  AOI21_X1 u2_u14_u4_U28 (.A( u2_u14_u4_n113 ) , .ZN( u2_u14_u4_n116 ) , .B2( u2_u14_u4_n173 ) , .B1( u2_u14_u4_n174 ) );
  AOI21_X1 u2_u14_u4_U29 (.ZN( u2_u14_u4_n115 ) , .B2( u2_u14_u4_n145 ) , .B1( u2_u14_u4_n146 ) , .A( u2_u14_u4_n156 ) );
  NOR2_X1 u2_u14_u4_U3 (.ZN( u2_u14_u4_n121 ) , .A1( u2_u14_u4_n181 ) , .A2( u2_u14_u4_n182 ) );
  OAI22_X1 u2_u14_u4_U30 (.ZN( u2_u14_u4_n114 ) , .A2( u2_u14_u4_n121 ) , .B1( u2_u14_u4_n160 ) , .B2( u2_u14_u4_n170 ) , .A1( u2_u14_u4_n171 ) );
  INV_X1 u2_u14_u4_U31 (.A( u2_u14_u4_n158 ) , .ZN( u2_u14_u4_n182 ) );
  INV_X1 u2_u14_u4_U32 (.ZN( u2_u14_u4_n181 ) , .A( u2_u14_u4_n96 ) );
  INV_X1 u2_u14_u4_U33 (.A( u2_u14_u4_n144 ) , .ZN( u2_u14_u4_n179 ) );
  INV_X1 u2_u14_u4_U34 (.A( u2_u14_u4_n157 ) , .ZN( u2_u14_u4_n178 ) );
  NAND2_X1 u2_u14_u4_U35 (.A2( u2_u14_u4_n154 ) , .A1( u2_u14_u4_n96 ) , .ZN( u2_u14_u4_n97 ) );
  INV_X1 u2_u14_u4_U36 (.ZN( u2_u14_u4_n186 ) , .A( u2_u14_u4_n95 ) );
  OAI221_X1 u2_u14_u4_U37 (.C1( u2_u14_u4_n134 ) , .B1( u2_u14_u4_n158 ) , .B2( u2_u14_u4_n171 ) , .C2( u2_u14_u4_n173 ) , .A( u2_u14_u4_n94 ) , .ZN( u2_u14_u4_n95 ) );
  AOI222_X1 u2_u14_u4_U38 (.B2( u2_u14_u4_n132 ) , .A1( u2_u14_u4_n138 ) , .C2( u2_u14_u4_n175 ) , .A2( u2_u14_u4_n179 ) , .C1( u2_u14_u4_n181 ) , .B1( u2_u14_u4_n185 ) , .ZN( u2_u14_u4_n94 ) );
  INV_X1 u2_u14_u4_U39 (.A( u2_u14_u4_n113 ) , .ZN( u2_u14_u4_n185 ) );
  INV_X1 u2_u14_u4_U4 (.A( u2_u14_u4_n117 ) , .ZN( u2_u14_u4_n184 ) );
  INV_X1 u2_u14_u4_U40 (.A( u2_u14_u4_n143 ) , .ZN( u2_u14_u4_n183 ) );
  NOR2_X1 u2_u14_u4_U41 (.ZN( u2_u14_u4_n138 ) , .A1( u2_u14_u4_n168 ) , .A2( u2_u14_u4_n169 ) );
  NOR2_X1 u2_u14_u4_U42 (.A1( u2_u14_u4_n150 ) , .A2( u2_u14_u4_n152 ) , .ZN( u2_u14_u4_n153 ) );
  NOR2_X1 u2_u14_u4_U43 (.A2( u2_u14_u4_n128 ) , .A1( u2_u14_u4_n138 ) , .ZN( u2_u14_u4_n156 ) );
  AOI22_X1 u2_u14_u4_U44 (.B2( u2_u14_u4_n122 ) , .A1( u2_u14_u4_n123 ) , .ZN( u2_u14_u4_n124 ) , .B1( u2_u14_u4_n128 ) , .A2( u2_u14_u4_n172 ) );
  INV_X1 u2_u14_u4_U45 (.A( u2_u14_u4_n153 ) , .ZN( u2_u14_u4_n172 ) );
  NAND2_X1 u2_u14_u4_U46 (.A2( u2_u14_u4_n120 ) , .ZN( u2_u14_u4_n123 ) , .A1( u2_u14_u4_n161 ) );
  AOI22_X1 u2_u14_u4_U47 (.B2( u2_u14_u4_n132 ) , .A2( u2_u14_u4_n133 ) , .ZN( u2_u14_u4_n140 ) , .A1( u2_u14_u4_n150 ) , .B1( u2_u14_u4_n179 ) );
  NAND2_X1 u2_u14_u4_U48 (.ZN( u2_u14_u4_n133 ) , .A2( u2_u14_u4_n146 ) , .A1( u2_u14_u4_n154 ) );
  NAND2_X1 u2_u14_u4_U49 (.A1( u2_u14_u4_n103 ) , .ZN( u2_u14_u4_n154 ) , .A2( u2_u14_u4_n98 ) );
  NOR4_X1 u2_u14_u4_U5 (.A4( u2_u14_u4_n106 ) , .A3( u2_u14_u4_n107 ) , .A2( u2_u14_u4_n108 ) , .A1( u2_u14_u4_n109 ) , .ZN( u2_u14_u4_n110 ) );
  NAND2_X1 u2_u14_u4_U50 (.A1( u2_u14_u4_n101 ) , .ZN( u2_u14_u4_n158 ) , .A2( u2_u14_u4_n99 ) );
  AOI21_X1 u2_u14_u4_U51 (.ZN( u2_u14_u4_n127 ) , .A( u2_u14_u4_n136 ) , .B2( u2_u14_u4_n150 ) , .B1( u2_u14_u4_n180 ) );
  INV_X1 u2_u14_u4_U52 (.A( u2_u14_u4_n160 ) , .ZN( u2_u14_u4_n180 ) );
  NAND2_X1 u2_u14_u4_U53 (.A2( u2_u14_u4_n104 ) , .A1( u2_u14_u4_n105 ) , .ZN( u2_u14_u4_n146 ) );
  NAND2_X1 u2_u14_u4_U54 (.A2( u2_u14_u4_n101 ) , .A1( u2_u14_u4_n102 ) , .ZN( u2_u14_u4_n160 ) );
  NAND2_X1 u2_u14_u4_U55 (.ZN( u2_u14_u4_n134 ) , .A1( u2_u14_u4_n98 ) , .A2( u2_u14_u4_n99 ) );
  NAND2_X1 u2_u14_u4_U56 (.A1( u2_u14_u4_n103 ) , .A2( u2_u14_u4_n104 ) , .ZN( u2_u14_u4_n143 ) );
  NAND2_X1 u2_u14_u4_U57 (.A2( u2_u14_u4_n105 ) , .ZN( u2_u14_u4_n145 ) , .A1( u2_u14_u4_n98 ) );
  NAND2_X1 u2_u14_u4_U58 (.A1( u2_u14_u4_n100 ) , .A2( u2_u14_u4_n105 ) , .ZN( u2_u14_u4_n120 ) );
  NAND2_X1 u2_u14_u4_U59 (.A1( u2_u14_u4_n102 ) , .A2( u2_u14_u4_n104 ) , .ZN( u2_u14_u4_n148 ) );
  AOI21_X1 u2_u14_u4_U6 (.ZN( u2_u14_u4_n106 ) , .B2( u2_u14_u4_n146 ) , .B1( u2_u14_u4_n158 ) , .A( u2_u14_u4_n170 ) );
  NAND2_X1 u2_u14_u4_U60 (.A2( u2_u14_u4_n100 ) , .A1( u2_u14_u4_n103 ) , .ZN( u2_u14_u4_n157 ) );
  INV_X1 u2_u14_u4_U61 (.A( u2_u14_u4_n150 ) , .ZN( u2_u14_u4_n173 ) );
  INV_X1 u2_u14_u4_U62 (.A( u2_u14_u4_n152 ) , .ZN( u2_u14_u4_n171 ) );
  NAND2_X1 u2_u14_u4_U63 (.A1( u2_u14_u4_n100 ) , .ZN( u2_u14_u4_n118 ) , .A2( u2_u14_u4_n99 ) );
  NAND2_X1 u2_u14_u4_U64 (.A2( u2_u14_u4_n100 ) , .A1( u2_u14_u4_n102 ) , .ZN( u2_u14_u4_n144 ) );
  NAND2_X1 u2_u14_u4_U65 (.A2( u2_u14_u4_n101 ) , .A1( u2_u14_u4_n105 ) , .ZN( u2_u14_u4_n96 ) );
  INV_X1 u2_u14_u4_U66 (.A( u2_u14_u4_n128 ) , .ZN( u2_u14_u4_n174 ) );
  NAND2_X1 u2_u14_u4_U67 (.A2( u2_u14_u4_n102 ) , .ZN( u2_u14_u4_n119 ) , .A1( u2_u14_u4_n98 ) );
  NAND2_X1 u2_u14_u4_U68 (.A2( u2_u14_u4_n101 ) , .A1( u2_u14_u4_n103 ) , .ZN( u2_u14_u4_n147 ) );
  NAND2_X1 u2_u14_u4_U69 (.A2( u2_u14_u4_n104 ) , .ZN( u2_u14_u4_n113 ) , .A1( u2_u14_u4_n99 ) );
  AOI21_X1 u2_u14_u4_U7 (.ZN( u2_u14_u4_n108 ) , .B2( u2_u14_u4_n134 ) , .B1( u2_u14_u4_n155 ) , .A( u2_u14_u4_n156 ) );
  NOR2_X1 u2_u14_u4_U70 (.A2( u2_u14_X_28 ) , .ZN( u2_u14_u4_n150 ) , .A1( u2_u14_u4_n168 ) );
  NOR2_X1 u2_u14_u4_U71 (.A2( u2_u14_X_29 ) , .ZN( u2_u14_u4_n152 ) , .A1( u2_u14_u4_n169 ) );
  NOR2_X1 u2_u14_u4_U72 (.A2( u2_u14_X_30 ) , .ZN( u2_u14_u4_n105 ) , .A1( u2_u14_u4_n176 ) );
  NOR2_X1 u2_u14_u4_U73 (.A2( u2_u14_X_26 ) , .ZN( u2_u14_u4_n100 ) , .A1( u2_u14_u4_n177 ) );
  NOR2_X1 u2_u14_u4_U74 (.A2( u2_u14_X_28 ) , .A1( u2_u14_X_29 ) , .ZN( u2_u14_u4_n128 ) );
  NOR2_X1 u2_u14_u4_U75 (.A2( u2_u14_X_27 ) , .A1( u2_u14_X_30 ) , .ZN( u2_u14_u4_n102 ) );
  NOR2_X1 u2_u14_u4_U76 (.A2( u2_u14_X_25 ) , .A1( u2_u14_X_26 ) , .ZN( u2_u14_u4_n98 ) );
  AND2_X1 u2_u14_u4_U77 (.A2( u2_u14_X_25 ) , .A1( u2_u14_X_26 ) , .ZN( u2_u14_u4_n104 ) );
  AND2_X1 u2_u14_u4_U78 (.A1( u2_u14_X_30 ) , .A2( u2_u14_u4_n176 ) , .ZN( u2_u14_u4_n99 ) );
  AND2_X1 u2_u14_u4_U79 (.A1( u2_u14_X_26 ) , .ZN( u2_u14_u4_n101 ) , .A2( u2_u14_u4_n177 ) );
  AOI21_X1 u2_u14_u4_U8 (.ZN( u2_u14_u4_n109 ) , .A( u2_u14_u4_n153 ) , .B1( u2_u14_u4_n159 ) , .B2( u2_u14_u4_n184 ) );
  AND2_X1 u2_u14_u4_U80 (.A1( u2_u14_X_27 ) , .A2( u2_u14_X_30 ) , .ZN( u2_u14_u4_n103 ) );
  INV_X1 u2_u14_u4_U81 (.A( u2_u14_X_28 ) , .ZN( u2_u14_u4_n169 ) );
  INV_X1 u2_u14_u4_U82 (.A( u2_u14_X_29 ) , .ZN( u2_u14_u4_n168 ) );
  INV_X1 u2_u14_u4_U83 (.A( u2_u14_X_25 ) , .ZN( u2_u14_u4_n177 ) );
  INV_X1 u2_u14_u4_U84 (.A( u2_u14_X_27 ) , .ZN( u2_u14_u4_n176 ) );
  NAND4_X1 u2_u14_u4_U85 (.ZN( u2_out14_25 ) , .A4( u2_u14_u4_n139 ) , .A3( u2_u14_u4_n140 ) , .A2( u2_u14_u4_n141 ) , .A1( u2_u14_u4_n142 ) );
  OAI21_X1 u2_u14_u4_U86 (.A( u2_u14_u4_n128 ) , .B2( u2_u14_u4_n129 ) , .B1( u2_u14_u4_n130 ) , .ZN( u2_u14_u4_n142 ) );
  OAI21_X1 u2_u14_u4_U87 (.B2( u2_u14_u4_n131 ) , .ZN( u2_u14_u4_n141 ) , .A( u2_u14_u4_n175 ) , .B1( u2_u14_u4_n183 ) );
  NAND4_X1 u2_u14_u4_U88 (.ZN( u2_out14_14 ) , .A4( u2_u14_u4_n124 ) , .A3( u2_u14_u4_n125 ) , .A2( u2_u14_u4_n126 ) , .A1( u2_u14_u4_n127 ) );
  AOI22_X1 u2_u14_u4_U89 (.B2( u2_u14_u4_n117 ) , .ZN( u2_u14_u4_n126 ) , .A1( u2_u14_u4_n129 ) , .B1( u2_u14_u4_n152 ) , .A2( u2_u14_u4_n175 ) );
  AOI211_X1 u2_u14_u4_U9 (.B( u2_u14_u4_n136 ) , .A( u2_u14_u4_n137 ) , .C2( u2_u14_u4_n138 ) , .ZN( u2_u14_u4_n139 ) , .C1( u2_u14_u4_n182 ) );
  AOI22_X1 u2_u14_u4_U90 (.ZN( u2_u14_u4_n125 ) , .B2( u2_u14_u4_n131 ) , .A2( u2_u14_u4_n132 ) , .B1( u2_u14_u4_n138 ) , .A1( u2_u14_u4_n178 ) );
  NAND4_X1 u2_u14_u4_U91 (.ZN( u2_out14_8 ) , .A4( u2_u14_u4_n110 ) , .A3( u2_u14_u4_n111 ) , .A2( u2_u14_u4_n112 ) , .A1( u2_u14_u4_n186 ) );
  NAND2_X1 u2_u14_u4_U92 (.ZN( u2_u14_u4_n112 ) , .A2( u2_u14_u4_n130 ) , .A1( u2_u14_u4_n150 ) );
  AOI22_X1 u2_u14_u4_U93 (.ZN( u2_u14_u4_n111 ) , .B2( u2_u14_u4_n132 ) , .A1( u2_u14_u4_n152 ) , .B1( u2_u14_u4_n178 ) , .A2( u2_u14_u4_n97 ) );
  AOI22_X1 u2_u14_u4_U94 (.B2( u2_u14_u4_n149 ) , .B1( u2_u14_u4_n150 ) , .A2( u2_u14_u4_n151 ) , .A1( u2_u14_u4_n152 ) , .ZN( u2_u14_u4_n167 ) );
  NOR4_X1 u2_u14_u4_U95 (.A4( u2_u14_u4_n162 ) , .A3( u2_u14_u4_n163 ) , .A2( u2_u14_u4_n164 ) , .A1( u2_u14_u4_n165 ) , .ZN( u2_u14_u4_n166 ) );
  NAND3_X1 u2_u14_u4_U96 (.ZN( u2_out14_3 ) , .A3( u2_u14_u4_n166 ) , .A1( u2_u14_u4_n167 ) , .A2( u2_u14_u4_n186 ) );
  NAND3_X1 u2_u14_u4_U97 (.A3( u2_u14_u4_n146 ) , .A2( u2_u14_u4_n147 ) , .A1( u2_u14_u4_n148 ) , .ZN( u2_u14_u4_n149 ) );
  NAND3_X1 u2_u14_u4_U98 (.A3( u2_u14_u4_n143 ) , .A2( u2_u14_u4_n144 ) , .A1( u2_u14_u4_n145 ) , .ZN( u2_u14_u4_n151 ) );
  NAND3_X1 u2_u14_u4_U99 (.A3( u2_u14_u4_n121 ) , .ZN( u2_u14_u4_n122 ) , .A2( u2_u14_u4_n144 ) , .A1( u2_u14_u4_n154 ) );
  INV_X1 u2_u14_u5_U10 (.A( u2_u14_u5_n121 ) , .ZN( u2_u14_u5_n177 ) );
  NOR3_X1 u2_u14_u5_U100 (.A3( u2_u14_u5_n141 ) , .A1( u2_u14_u5_n142 ) , .ZN( u2_u14_u5_n143 ) , .A2( u2_u14_u5_n191 ) );
  NAND4_X1 u2_u14_u5_U101 (.ZN( u2_out14_4 ) , .A4( u2_u14_u5_n112 ) , .A2( u2_u14_u5_n113 ) , .A1( u2_u14_u5_n114 ) , .A3( u2_u14_u5_n195 ) );
  AOI211_X1 u2_u14_u5_U102 (.A( u2_u14_u5_n110 ) , .C1( u2_u14_u5_n111 ) , .ZN( u2_u14_u5_n112 ) , .B( u2_u14_u5_n118 ) , .C2( u2_u14_u5_n177 ) );
  AOI222_X1 u2_u14_u5_U103 (.ZN( u2_u14_u5_n113 ) , .A1( u2_u14_u5_n131 ) , .C1( u2_u14_u5_n148 ) , .B2( u2_u14_u5_n174 ) , .C2( u2_u14_u5_n178 ) , .A2( u2_u14_u5_n179 ) , .B1( u2_u14_u5_n99 ) );
  NAND3_X1 u2_u14_u5_U104 (.A2( u2_u14_u5_n154 ) , .A3( u2_u14_u5_n158 ) , .A1( u2_u14_u5_n161 ) , .ZN( u2_u14_u5_n99 ) );
  NOR2_X1 u2_u14_u5_U11 (.ZN( u2_u14_u5_n160 ) , .A2( u2_u14_u5_n173 ) , .A1( u2_u14_u5_n177 ) );
  INV_X1 u2_u14_u5_U12 (.A( u2_u14_u5_n150 ) , .ZN( u2_u14_u5_n174 ) );
  AOI21_X1 u2_u14_u5_U13 (.A( u2_u14_u5_n160 ) , .B2( u2_u14_u5_n161 ) , .ZN( u2_u14_u5_n162 ) , .B1( u2_u14_u5_n192 ) );
  INV_X1 u2_u14_u5_U14 (.A( u2_u14_u5_n159 ) , .ZN( u2_u14_u5_n192 ) );
  AOI21_X1 u2_u14_u5_U15 (.A( u2_u14_u5_n156 ) , .B2( u2_u14_u5_n157 ) , .B1( u2_u14_u5_n158 ) , .ZN( u2_u14_u5_n163 ) );
  AOI21_X1 u2_u14_u5_U16 (.B2( u2_u14_u5_n139 ) , .B1( u2_u14_u5_n140 ) , .ZN( u2_u14_u5_n141 ) , .A( u2_u14_u5_n150 ) );
  OAI21_X1 u2_u14_u5_U17 (.A( u2_u14_u5_n133 ) , .B2( u2_u14_u5_n134 ) , .B1( u2_u14_u5_n135 ) , .ZN( u2_u14_u5_n142 ) );
  OAI21_X1 u2_u14_u5_U18 (.ZN( u2_u14_u5_n133 ) , .B2( u2_u14_u5_n147 ) , .A( u2_u14_u5_n173 ) , .B1( u2_u14_u5_n188 ) );
  NAND2_X1 u2_u14_u5_U19 (.A2( u2_u14_u5_n119 ) , .A1( u2_u14_u5_n123 ) , .ZN( u2_u14_u5_n137 ) );
  INV_X1 u2_u14_u5_U20 (.A( u2_u14_u5_n155 ) , .ZN( u2_u14_u5_n194 ) );
  NAND2_X1 u2_u14_u5_U21 (.A1( u2_u14_u5_n121 ) , .ZN( u2_u14_u5_n132 ) , .A2( u2_u14_u5_n172 ) );
  NAND2_X1 u2_u14_u5_U22 (.A2( u2_u14_u5_n122 ) , .ZN( u2_u14_u5_n136 ) , .A1( u2_u14_u5_n154 ) );
  NAND2_X1 u2_u14_u5_U23 (.A2( u2_u14_u5_n119 ) , .A1( u2_u14_u5_n120 ) , .ZN( u2_u14_u5_n159 ) );
  INV_X1 u2_u14_u5_U24 (.A( u2_u14_u5_n156 ) , .ZN( u2_u14_u5_n175 ) );
  INV_X1 u2_u14_u5_U25 (.A( u2_u14_u5_n158 ) , .ZN( u2_u14_u5_n188 ) );
  INV_X1 u2_u14_u5_U26 (.A( u2_u14_u5_n152 ) , .ZN( u2_u14_u5_n179 ) );
  INV_X1 u2_u14_u5_U27 (.A( u2_u14_u5_n140 ) , .ZN( u2_u14_u5_n182 ) );
  INV_X1 u2_u14_u5_U28 (.A( u2_u14_u5_n151 ) , .ZN( u2_u14_u5_n183 ) );
  INV_X1 u2_u14_u5_U29 (.A( u2_u14_u5_n123 ) , .ZN( u2_u14_u5_n185 ) );
  NOR2_X1 u2_u14_u5_U3 (.ZN( u2_u14_u5_n134 ) , .A1( u2_u14_u5_n183 ) , .A2( u2_u14_u5_n190 ) );
  INV_X1 u2_u14_u5_U30 (.A( u2_u14_u5_n161 ) , .ZN( u2_u14_u5_n184 ) );
  INV_X1 u2_u14_u5_U31 (.A( u2_u14_u5_n139 ) , .ZN( u2_u14_u5_n189 ) );
  INV_X1 u2_u14_u5_U32 (.A( u2_u14_u5_n157 ) , .ZN( u2_u14_u5_n190 ) );
  INV_X1 u2_u14_u5_U33 (.A( u2_u14_u5_n120 ) , .ZN( u2_u14_u5_n193 ) );
  NAND2_X1 u2_u14_u5_U34 (.ZN( u2_u14_u5_n111 ) , .A1( u2_u14_u5_n140 ) , .A2( u2_u14_u5_n155 ) );
  INV_X1 u2_u14_u5_U35 (.A( u2_u14_u5_n117 ) , .ZN( u2_u14_u5_n196 ) );
  OAI221_X1 u2_u14_u5_U36 (.A( u2_u14_u5_n116 ) , .ZN( u2_u14_u5_n117 ) , .B2( u2_u14_u5_n119 ) , .C1( u2_u14_u5_n153 ) , .C2( u2_u14_u5_n158 ) , .B1( u2_u14_u5_n172 ) );
  AOI222_X1 u2_u14_u5_U37 (.ZN( u2_u14_u5_n116 ) , .B2( u2_u14_u5_n145 ) , .C1( u2_u14_u5_n148 ) , .A2( u2_u14_u5_n174 ) , .C2( u2_u14_u5_n177 ) , .B1( u2_u14_u5_n187 ) , .A1( u2_u14_u5_n193 ) );
  INV_X1 u2_u14_u5_U38 (.A( u2_u14_u5_n115 ) , .ZN( u2_u14_u5_n187 ) );
  NOR2_X1 u2_u14_u5_U39 (.ZN( u2_u14_u5_n100 ) , .A1( u2_u14_u5_n170 ) , .A2( u2_u14_u5_n180 ) );
  INV_X1 u2_u14_u5_U4 (.A( u2_u14_u5_n138 ) , .ZN( u2_u14_u5_n191 ) );
  AOI22_X1 u2_u14_u5_U40 (.B2( u2_u14_u5_n131 ) , .A2( u2_u14_u5_n146 ) , .ZN( u2_u14_u5_n169 ) , .B1( u2_u14_u5_n174 ) , .A1( u2_u14_u5_n185 ) );
  NOR2_X1 u2_u14_u5_U41 (.A1( u2_u14_u5_n146 ) , .ZN( u2_u14_u5_n150 ) , .A2( u2_u14_u5_n173 ) );
  AOI21_X1 u2_u14_u5_U42 (.A( u2_u14_u5_n118 ) , .B2( u2_u14_u5_n145 ) , .ZN( u2_u14_u5_n168 ) , .B1( u2_u14_u5_n186 ) );
  INV_X1 u2_u14_u5_U43 (.A( u2_u14_u5_n122 ) , .ZN( u2_u14_u5_n186 ) );
  NOR2_X1 u2_u14_u5_U44 (.A1( u2_u14_u5_n146 ) , .ZN( u2_u14_u5_n152 ) , .A2( u2_u14_u5_n176 ) );
  NOR2_X1 u2_u14_u5_U45 (.A1( u2_u14_u5_n115 ) , .ZN( u2_u14_u5_n118 ) , .A2( u2_u14_u5_n153 ) );
  NOR2_X1 u2_u14_u5_U46 (.A2( u2_u14_u5_n145 ) , .ZN( u2_u14_u5_n156 ) , .A1( u2_u14_u5_n174 ) );
  NOR2_X1 u2_u14_u5_U47 (.ZN( u2_u14_u5_n121 ) , .A2( u2_u14_u5_n145 ) , .A1( u2_u14_u5_n176 ) );
  AOI22_X1 u2_u14_u5_U48 (.ZN( u2_u14_u5_n114 ) , .A2( u2_u14_u5_n137 ) , .A1( u2_u14_u5_n145 ) , .B2( u2_u14_u5_n175 ) , .B1( u2_u14_u5_n193 ) );
  OAI211_X1 u2_u14_u5_U49 (.B( u2_u14_u5_n124 ) , .A( u2_u14_u5_n125 ) , .C2( u2_u14_u5_n126 ) , .C1( u2_u14_u5_n127 ) , .ZN( u2_u14_u5_n128 ) );
  OAI21_X1 u2_u14_u5_U5 (.B2( u2_u14_u5_n136 ) , .B1( u2_u14_u5_n137 ) , .ZN( u2_u14_u5_n138 ) , .A( u2_u14_u5_n177 ) );
  NOR3_X1 u2_u14_u5_U50 (.ZN( u2_u14_u5_n127 ) , .A1( u2_u14_u5_n136 ) , .A3( u2_u14_u5_n148 ) , .A2( u2_u14_u5_n182 ) );
  OAI21_X1 u2_u14_u5_U51 (.ZN( u2_u14_u5_n124 ) , .A( u2_u14_u5_n177 ) , .B2( u2_u14_u5_n183 ) , .B1( u2_u14_u5_n189 ) );
  OAI21_X1 u2_u14_u5_U52 (.ZN( u2_u14_u5_n125 ) , .A( u2_u14_u5_n174 ) , .B2( u2_u14_u5_n185 ) , .B1( u2_u14_u5_n190 ) );
  AOI21_X1 u2_u14_u5_U53 (.A( u2_u14_u5_n153 ) , .B2( u2_u14_u5_n154 ) , .B1( u2_u14_u5_n155 ) , .ZN( u2_u14_u5_n164 ) );
  AOI21_X1 u2_u14_u5_U54 (.ZN( u2_u14_u5_n110 ) , .B1( u2_u14_u5_n122 ) , .B2( u2_u14_u5_n139 ) , .A( u2_u14_u5_n153 ) );
  INV_X1 u2_u14_u5_U55 (.A( u2_u14_u5_n153 ) , .ZN( u2_u14_u5_n176 ) );
  INV_X1 u2_u14_u5_U56 (.A( u2_u14_u5_n126 ) , .ZN( u2_u14_u5_n173 ) );
  AND2_X1 u2_u14_u5_U57 (.A2( u2_u14_u5_n104 ) , .A1( u2_u14_u5_n107 ) , .ZN( u2_u14_u5_n147 ) );
  AND2_X1 u2_u14_u5_U58 (.A2( u2_u14_u5_n104 ) , .A1( u2_u14_u5_n108 ) , .ZN( u2_u14_u5_n148 ) );
  NAND2_X1 u2_u14_u5_U59 (.A1( u2_u14_u5_n105 ) , .A2( u2_u14_u5_n106 ) , .ZN( u2_u14_u5_n158 ) );
  INV_X1 u2_u14_u5_U6 (.A( u2_u14_u5_n135 ) , .ZN( u2_u14_u5_n178 ) );
  NAND2_X1 u2_u14_u5_U60 (.A2( u2_u14_u5_n108 ) , .A1( u2_u14_u5_n109 ) , .ZN( u2_u14_u5_n139 ) );
  NAND2_X1 u2_u14_u5_U61 (.A1( u2_u14_u5_n106 ) , .A2( u2_u14_u5_n108 ) , .ZN( u2_u14_u5_n119 ) );
  NAND2_X1 u2_u14_u5_U62 (.A2( u2_u14_u5_n103 ) , .A1( u2_u14_u5_n105 ) , .ZN( u2_u14_u5_n140 ) );
  NAND2_X1 u2_u14_u5_U63 (.A2( u2_u14_u5_n104 ) , .A1( u2_u14_u5_n105 ) , .ZN( u2_u14_u5_n155 ) );
  NAND2_X1 u2_u14_u5_U64 (.A2( u2_u14_u5_n106 ) , .A1( u2_u14_u5_n107 ) , .ZN( u2_u14_u5_n122 ) );
  NAND2_X1 u2_u14_u5_U65 (.A2( u2_u14_u5_n100 ) , .A1( u2_u14_u5_n106 ) , .ZN( u2_u14_u5_n115 ) );
  NAND2_X1 u2_u14_u5_U66 (.A2( u2_u14_u5_n100 ) , .A1( u2_u14_u5_n103 ) , .ZN( u2_u14_u5_n161 ) );
  NAND2_X1 u2_u14_u5_U67 (.A1( u2_u14_u5_n105 ) , .A2( u2_u14_u5_n109 ) , .ZN( u2_u14_u5_n154 ) );
  INV_X1 u2_u14_u5_U68 (.A( u2_u14_u5_n146 ) , .ZN( u2_u14_u5_n172 ) );
  NAND2_X1 u2_u14_u5_U69 (.A1( u2_u14_u5_n103 ) , .A2( u2_u14_u5_n108 ) , .ZN( u2_u14_u5_n123 ) );
  OAI22_X1 u2_u14_u5_U7 (.B2( u2_u14_u5_n149 ) , .B1( u2_u14_u5_n150 ) , .A2( u2_u14_u5_n151 ) , .A1( u2_u14_u5_n152 ) , .ZN( u2_u14_u5_n165 ) );
  NAND2_X1 u2_u14_u5_U70 (.A2( u2_u14_u5_n103 ) , .A1( u2_u14_u5_n107 ) , .ZN( u2_u14_u5_n151 ) );
  NAND2_X1 u2_u14_u5_U71 (.A2( u2_u14_u5_n107 ) , .A1( u2_u14_u5_n109 ) , .ZN( u2_u14_u5_n120 ) );
  NAND2_X1 u2_u14_u5_U72 (.A2( u2_u14_u5_n100 ) , .A1( u2_u14_u5_n109 ) , .ZN( u2_u14_u5_n157 ) );
  AND2_X1 u2_u14_u5_U73 (.A2( u2_u14_u5_n100 ) , .A1( u2_u14_u5_n104 ) , .ZN( u2_u14_u5_n131 ) );
  INV_X1 u2_u14_u5_U74 (.A( u2_u14_u5_n102 ) , .ZN( u2_u14_u5_n195 ) );
  OAI221_X1 u2_u14_u5_U75 (.A( u2_u14_u5_n101 ) , .ZN( u2_u14_u5_n102 ) , .C2( u2_u14_u5_n115 ) , .C1( u2_u14_u5_n126 ) , .B1( u2_u14_u5_n134 ) , .B2( u2_u14_u5_n160 ) );
  OAI21_X1 u2_u14_u5_U76 (.ZN( u2_u14_u5_n101 ) , .B1( u2_u14_u5_n137 ) , .A( u2_u14_u5_n146 ) , .B2( u2_u14_u5_n147 ) );
  NOR2_X1 u2_u14_u5_U77 (.A2( u2_u14_X_34 ) , .A1( u2_u14_X_35 ) , .ZN( u2_u14_u5_n145 ) );
  NOR2_X1 u2_u14_u5_U78 (.A2( u2_u14_X_34 ) , .ZN( u2_u14_u5_n146 ) , .A1( u2_u14_u5_n171 ) );
  NOR2_X1 u2_u14_u5_U79 (.A2( u2_u14_X_31 ) , .A1( u2_u14_X_32 ) , .ZN( u2_u14_u5_n103 ) );
  NOR3_X1 u2_u14_u5_U8 (.A2( u2_u14_u5_n147 ) , .A1( u2_u14_u5_n148 ) , .ZN( u2_u14_u5_n149 ) , .A3( u2_u14_u5_n194 ) );
  NOR2_X1 u2_u14_u5_U80 (.A2( u2_u14_X_36 ) , .ZN( u2_u14_u5_n105 ) , .A1( u2_u14_u5_n180 ) );
  NOR2_X1 u2_u14_u5_U81 (.A2( u2_u14_X_33 ) , .ZN( u2_u14_u5_n108 ) , .A1( u2_u14_u5_n170 ) );
  NOR2_X1 u2_u14_u5_U82 (.A2( u2_u14_X_33 ) , .A1( u2_u14_X_36 ) , .ZN( u2_u14_u5_n107 ) );
  NOR2_X1 u2_u14_u5_U83 (.A2( u2_u14_X_31 ) , .ZN( u2_u14_u5_n104 ) , .A1( u2_u14_u5_n181 ) );
  NAND2_X1 u2_u14_u5_U84 (.A2( u2_u14_X_34 ) , .A1( u2_u14_X_35 ) , .ZN( u2_u14_u5_n153 ) );
  NAND2_X1 u2_u14_u5_U85 (.A1( u2_u14_X_34 ) , .ZN( u2_u14_u5_n126 ) , .A2( u2_u14_u5_n171 ) );
  AND2_X1 u2_u14_u5_U86 (.A1( u2_u14_X_31 ) , .A2( u2_u14_X_32 ) , .ZN( u2_u14_u5_n106 ) );
  AND2_X1 u2_u14_u5_U87 (.A1( u2_u14_X_31 ) , .ZN( u2_u14_u5_n109 ) , .A2( u2_u14_u5_n181 ) );
  INV_X1 u2_u14_u5_U88 (.A( u2_u14_X_33 ) , .ZN( u2_u14_u5_n180 ) );
  INV_X1 u2_u14_u5_U89 (.A( u2_u14_X_35 ) , .ZN( u2_u14_u5_n171 ) );
  NOR2_X1 u2_u14_u5_U9 (.ZN( u2_u14_u5_n135 ) , .A1( u2_u14_u5_n173 ) , .A2( u2_u14_u5_n176 ) );
  INV_X1 u2_u14_u5_U90 (.A( u2_u14_X_36 ) , .ZN( u2_u14_u5_n170 ) );
  INV_X1 u2_u14_u5_U91 (.A( u2_u14_X_32 ) , .ZN( u2_u14_u5_n181 ) );
  NAND4_X1 u2_u14_u5_U92 (.ZN( u2_out14_29 ) , .A4( u2_u14_u5_n129 ) , .A3( u2_u14_u5_n130 ) , .A2( u2_u14_u5_n168 ) , .A1( u2_u14_u5_n196 ) );
  AOI221_X1 u2_u14_u5_U93 (.A( u2_u14_u5_n128 ) , .ZN( u2_u14_u5_n129 ) , .C2( u2_u14_u5_n132 ) , .B2( u2_u14_u5_n159 ) , .B1( u2_u14_u5_n176 ) , .C1( u2_u14_u5_n184 ) );
  AOI222_X1 u2_u14_u5_U94 (.ZN( u2_u14_u5_n130 ) , .A2( u2_u14_u5_n146 ) , .B1( u2_u14_u5_n147 ) , .C2( u2_u14_u5_n175 ) , .B2( u2_u14_u5_n179 ) , .A1( u2_u14_u5_n188 ) , .C1( u2_u14_u5_n194 ) );
  NAND4_X1 u2_u14_u5_U95 (.ZN( u2_out14_19 ) , .A4( u2_u14_u5_n166 ) , .A3( u2_u14_u5_n167 ) , .A2( u2_u14_u5_n168 ) , .A1( u2_u14_u5_n169 ) );
  AOI22_X1 u2_u14_u5_U96 (.B2( u2_u14_u5_n145 ) , .A2( u2_u14_u5_n146 ) , .ZN( u2_u14_u5_n167 ) , .B1( u2_u14_u5_n182 ) , .A1( u2_u14_u5_n189 ) );
  NOR4_X1 u2_u14_u5_U97 (.A4( u2_u14_u5_n162 ) , .A3( u2_u14_u5_n163 ) , .A2( u2_u14_u5_n164 ) , .A1( u2_u14_u5_n165 ) , .ZN( u2_u14_u5_n166 ) );
  NAND4_X1 u2_u14_u5_U98 (.ZN( u2_out14_11 ) , .A4( u2_u14_u5_n143 ) , .A3( u2_u14_u5_n144 ) , .A2( u2_u14_u5_n169 ) , .A1( u2_u14_u5_n196 ) );
  AOI22_X1 u2_u14_u5_U99 (.A2( u2_u14_u5_n132 ) , .ZN( u2_u14_u5_n144 ) , .B2( u2_u14_u5_n145 ) , .B1( u2_u14_u5_n184 ) , .A1( u2_u14_u5_n194 ) );
  AOI22_X1 u2_u14_u6_U10 (.A2( u2_u14_u6_n151 ) , .B2( u2_u14_u6_n161 ) , .A1( u2_u14_u6_n167 ) , .B1( u2_u14_u6_n170 ) , .ZN( u2_u14_u6_n89 ) );
  AOI21_X1 u2_u14_u6_U11 (.B1( u2_u14_u6_n107 ) , .B2( u2_u14_u6_n132 ) , .A( u2_u14_u6_n158 ) , .ZN( u2_u14_u6_n88 ) );
  AOI21_X1 u2_u14_u6_U12 (.B2( u2_u14_u6_n147 ) , .B1( u2_u14_u6_n148 ) , .ZN( u2_u14_u6_n149 ) , .A( u2_u14_u6_n158 ) );
  AOI21_X1 u2_u14_u6_U13 (.ZN( u2_u14_u6_n106 ) , .A( u2_u14_u6_n142 ) , .B2( u2_u14_u6_n159 ) , .B1( u2_u14_u6_n164 ) );
  INV_X1 u2_u14_u6_U14 (.A( u2_u14_u6_n155 ) , .ZN( u2_u14_u6_n161 ) );
  INV_X1 u2_u14_u6_U15 (.A( u2_u14_u6_n128 ) , .ZN( u2_u14_u6_n164 ) );
  NAND2_X1 u2_u14_u6_U16 (.ZN( u2_u14_u6_n110 ) , .A1( u2_u14_u6_n122 ) , .A2( u2_u14_u6_n129 ) );
  NAND2_X1 u2_u14_u6_U17 (.ZN( u2_u14_u6_n124 ) , .A2( u2_u14_u6_n146 ) , .A1( u2_u14_u6_n148 ) );
  INV_X1 u2_u14_u6_U18 (.A( u2_u14_u6_n132 ) , .ZN( u2_u14_u6_n171 ) );
  AND2_X1 u2_u14_u6_U19 (.A1( u2_u14_u6_n100 ) , .ZN( u2_u14_u6_n130 ) , .A2( u2_u14_u6_n147 ) );
  INV_X1 u2_u14_u6_U20 (.A( u2_u14_u6_n127 ) , .ZN( u2_u14_u6_n173 ) );
  INV_X1 u2_u14_u6_U21 (.A( u2_u14_u6_n121 ) , .ZN( u2_u14_u6_n167 ) );
  INV_X1 u2_u14_u6_U22 (.A( u2_u14_u6_n100 ) , .ZN( u2_u14_u6_n169 ) );
  INV_X1 u2_u14_u6_U23 (.A( u2_u14_u6_n123 ) , .ZN( u2_u14_u6_n170 ) );
  INV_X1 u2_u14_u6_U24 (.A( u2_u14_u6_n113 ) , .ZN( u2_u14_u6_n168 ) );
  AND2_X1 u2_u14_u6_U25 (.A1( u2_u14_u6_n107 ) , .A2( u2_u14_u6_n119 ) , .ZN( u2_u14_u6_n133 ) );
  AND2_X1 u2_u14_u6_U26 (.A2( u2_u14_u6_n121 ) , .A1( u2_u14_u6_n122 ) , .ZN( u2_u14_u6_n131 ) );
  AND3_X1 u2_u14_u6_U27 (.ZN( u2_u14_u6_n120 ) , .A2( u2_u14_u6_n127 ) , .A1( u2_u14_u6_n132 ) , .A3( u2_u14_u6_n145 ) );
  INV_X1 u2_u14_u6_U28 (.A( u2_u14_u6_n146 ) , .ZN( u2_u14_u6_n163 ) );
  AOI222_X1 u2_u14_u6_U29 (.ZN( u2_u14_u6_n114 ) , .A1( u2_u14_u6_n118 ) , .A2( u2_u14_u6_n126 ) , .B2( u2_u14_u6_n151 ) , .C2( u2_u14_u6_n159 ) , .C1( u2_u14_u6_n168 ) , .B1( u2_u14_u6_n169 ) );
  INV_X1 u2_u14_u6_U3 (.A( u2_u14_u6_n110 ) , .ZN( u2_u14_u6_n166 ) );
  NOR2_X1 u2_u14_u6_U30 (.A1( u2_u14_u6_n162 ) , .A2( u2_u14_u6_n165 ) , .ZN( u2_u14_u6_n98 ) );
  NAND2_X1 u2_u14_u6_U31 (.A1( u2_u14_u6_n144 ) , .ZN( u2_u14_u6_n151 ) , .A2( u2_u14_u6_n158 ) );
  NAND2_X1 u2_u14_u6_U32 (.ZN( u2_u14_u6_n132 ) , .A1( u2_u14_u6_n91 ) , .A2( u2_u14_u6_n97 ) );
  AOI22_X1 u2_u14_u6_U33 (.B2( u2_u14_u6_n110 ) , .B1( u2_u14_u6_n111 ) , .A1( u2_u14_u6_n112 ) , .ZN( u2_u14_u6_n115 ) , .A2( u2_u14_u6_n161 ) );
  NAND4_X1 u2_u14_u6_U34 (.A3( u2_u14_u6_n109 ) , .ZN( u2_u14_u6_n112 ) , .A4( u2_u14_u6_n132 ) , .A2( u2_u14_u6_n147 ) , .A1( u2_u14_u6_n166 ) );
  NOR2_X1 u2_u14_u6_U35 (.ZN( u2_u14_u6_n109 ) , .A1( u2_u14_u6_n170 ) , .A2( u2_u14_u6_n173 ) );
  NOR2_X1 u2_u14_u6_U36 (.A2( u2_u14_u6_n126 ) , .ZN( u2_u14_u6_n155 ) , .A1( u2_u14_u6_n160 ) );
  NAND2_X1 u2_u14_u6_U37 (.ZN( u2_u14_u6_n146 ) , .A2( u2_u14_u6_n94 ) , .A1( u2_u14_u6_n99 ) );
  AOI21_X1 u2_u14_u6_U38 (.A( u2_u14_u6_n144 ) , .B2( u2_u14_u6_n145 ) , .B1( u2_u14_u6_n146 ) , .ZN( u2_u14_u6_n150 ) );
  AOI211_X1 u2_u14_u6_U39 (.B( u2_u14_u6_n134 ) , .A( u2_u14_u6_n135 ) , .C1( u2_u14_u6_n136 ) , .ZN( u2_u14_u6_n137 ) , .C2( u2_u14_u6_n151 ) );
  INV_X1 u2_u14_u6_U4 (.A( u2_u14_u6_n142 ) , .ZN( u2_u14_u6_n174 ) );
  AOI21_X1 u2_u14_u6_U40 (.B2( u2_u14_u6_n132 ) , .B1( u2_u14_u6_n133 ) , .ZN( u2_u14_u6_n134 ) , .A( u2_u14_u6_n158 ) );
  NAND4_X1 u2_u14_u6_U41 (.A4( u2_u14_u6_n127 ) , .A3( u2_u14_u6_n128 ) , .A2( u2_u14_u6_n129 ) , .A1( u2_u14_u6_n130 ) , .ZN( u2_u14_u6_n136 ) );
  AOI21_X1 u2_u14_u6_U42 (.B1( u2_u14_u6_n131 ) , .ZN( u2_u14_u6_n135 ) , .A( u2_u14_u6_n144 ) , .B2( u2_u14_u6_n146 ) );
  INV_X1 u2_u14_u6_U43 (.A( u2_u14_u6_n111 ) , .ZN( u2_u14_u6_n158 ) );
  NAND2_X1 u2_u14_u6_U44 (.ZN( u2_u14_u6_n127 ) , .A1( u2_u14_u6_n91 ) , .A2( u2_u14_u6_n92 ) );
  NAND2_X1 u2_u14_u6_U45 (.ZN( u2_u14_u6_n129 ) , .A2( u2_u14_u6_n95 ) , .A1( u2_u14_u6_n96 ) );
  INV_X1 u2_u14_u6_U46 (.A( u2_u14_u6_n144 ) , .ZN( u2_u14_u6_n159 ) );
  NAND2_X1 u2_u14_u6_U47 (.ZN( u2_u14_u6_n145 ) , .A2( u2_u14_u6_n97 ) , .A1( u2_u14_u6_n98 ) );
  NAND2_X1 u2_u14_u6_U48 (.ZN( u2_u14_u6_n148 ) , .A2( u2_u14_u6_n92 ) , .A1( u2_u14_u6_n94 ) );
  NAND2_X1 u2_u14_u6_U49 (.ZN( u2_u14_u6_n108 ) , .A2( u2_u14_u6_n139 ) , .A1( u2_u14_u6_n144 ) );
  NAND2_X1 u2_u14_u6_U5 (.A2( u2_u14_u6_n143 ) , .ZN( u2_u14_u6_n152 ) , .A1( u2_u14_u6_n166 ) );
  NAND2_X1 u2_u14_u6_U50 (.ZN( u2_u14_u6_n121 ) , .A2( u2_u14_u6_n95 ) , .A1( u2_u14_u6_n97 ) );
  NAND2_X1 u2_u14_u6_U51 (.ZN( u2_u14_u6_n107 ) , .A2( u2_u14_u6_n92 ) , .A1( u2_u14_u6_n95 ) );
  AND2_X1 u2_u14_u6_U52 (.ZN( u2_u14_u6_n118 ) , .A2( u2_u14_u6_n91 ) , .A1( u2_u14_u6_n99 ) );
  NAND2_X1 u2_u14_u6_U53 (.ZN( u2_u14_u6_n147 ) , .A2( u2_u14_u6_n98 ) , .A1( u2_u14_u6_n99 ) );
  NAND2_X1 u2_u14_u6_U54 (.ZN( u2_u14_u6_n128 ) , .A1( u2_u14_u6_n94 ) , .A2( u2_u14_u6_n96 ) );
  NAND2_X1 u2_u14_u6_U55 (.ZN( u2_u14_u6_n119 ) , .A2( u2_u14_u6_n95 ) , .A1( u2_u14_u6_n99 ) );
  NAND2_X1 u2_u14_u6_U56 (.ZN( u2_u14_u6_n123 ) , .A2( u2_u14_u6_n91 ) , .A1( u2_u14_u6_n96 ) );
  NAND2_X1 u2_u14_u6_U57 (.ZN( u2_u14_u6_n100 ) , .A2( u2_u14_u6_n92 ) , .A1( u2_u14_u6_n98 ) );
  NAND2_X1 u2_u14_u6_U58 (.ZN( u2_u14_u6_n122 ) , .A1( u2_u14_u6_n94 ) , .A2( u2_u14_u6_n97 ) );
  INV_X1 u2_u14_u6_U59 (.A( u2_u14_u6_n139 ) , .ZN( u2_u14_u6_n160 ) );
  AOI22_X1 u2_u14_u6_U6 (.B2( u2_u14_u6_n101 ) , .A1( u2_u14_u6_n102 ) , .ZN( u2_u14_u6_n103 ) , .B1( u2_u14_u6_n160 ) , .A2( u2_u14_u6_n161 ) );
  NAND2_X1 u2_u14_u6_U60 (.ZN( u2_u14_u6_n113 ) , .A1( u2_u14_u6_n96 ) , .A2( u2_u14_u6_n98 ) );
  NOR2_X1 u2_u14_u6_U61 (.A2( u2_u14_X_40 ) , .A1( u2_u14_X_41 ) , .ZN( u2_u14_u6_n126 ) );
  NOR2_X1 u2_u14_u6_U62 (.A2( u2_u14_X_39 ) , .A1( u2_u14_X_42 ) , .ZN( u2_u14_u6_n92 ) );
  NOR2_X1 u2_u14_u6_U63 (.A2( u2_u14_X_39 ) , .A1( u2_u14_u6_n156 ) , .ZN( u2_u14_u6_n97 ) );
  NOR2_X1 u2_u14_u6_U64 (.A2( u2_u14_X_38 ) , .A1( u2_u14_u6_n165 ) , .ZN( u2_u14_u6_n95 ) );
  NOR2_X1 u2_u14_u6_U65 (.A2( u2_u14_X_41 ) , .ZN( u2_u14_u6_n111 ) , .A1( u2_u14_u6_n157 ) );
  NOR2_X1 u2_u14_u6_U66 (.A2( u2_u14_X_37 ) , .A1( u2_u14_u6_n162 ) , .ZN( u2_u14_u6_n94 ) );
  NOR2_X1 u2_u14_u6_U67 (.A2( u2_u14_X_37 ) , .A1( u2_u14_X_38 ) , .ZN( u2_u14_u6_n91 ) );
  NAND2_X1 u2_u14_u6_U68 (.A1( u2_u14_X_41 ) , .ZN( u2_u14_u6_n144 ) , .A2( u2_u14_u6_n157 ) );
  NAND2_X1 u2_u14_u6_U69 (.A2( u2_u14_X_40 ) , .A1( u2_u14_X_41 ) , .ZN( u2_u14_u6_n139 ) );
  NOR2_X1 u2_u14_u6_U7 (.A1( u2_u14_u6_n118 ) , .ZN( u2_u14_u6_n143 ) , .A2( u2_u14_u6_n168 ) );
  AND2_X1 u2_u14_u6_U70 (.A1( u2_u14_X_39 ) , .A2( u2_u14_u6_n156 ) , .ZN( u2_u14_u6_n96 ) );
  AND2_X1 u2_u14_u6_U71 (.A1( u2_u14_X_39 ) , .A2( u2_u14_X_42 ) , .ZN( u2_u14_u6_n99 ) );
  INV_X1 u2_u14_u6_U72 (.A( u2_u14_X_40 ) , .ZN( u2_u14_u6_n157 ) );
  INV_X1 u2_u14_u6_U73 (.A( u2_u14_X_37 ) , .ZN( u2_u14_u6_n165 ) );
  INV_X1 u2_u14_u6_U74 (.A( u2_u14_X_38 ) , .ZN( u2_u14_u6_n162 ) );
  INV_X1 u2_u14_u6_U75 (.A( u2_u14_X_42 ) , .ZN( u2_u14_u6_n156 ) );
  NAND4_X1 u2_u14_u6_U76 (.ZN( u2_out14_32 ) , .A4( u2_u14_u6_n103 ) , .A3( u2_u14_u6_n104 ) , .A2( u2_u14_u6_n105 ) , .A1( u2_u14_u6_n106 ) );
  AOI22_X1 u2_u14_u6_U77 (.ZN( u2_u14_u6_n105 ) , .A2( u2_u14_u6_n108 ) , .A1( u2_u14_u6_n118 ) , .B2( u2_u14_u6_n126 ) , .B1( u2_u14_u6_n171 ) );
  AOI22_X1 u2_u14_u6_U78 (.ZN( u2_u14_u6_n104 ) , .A1( u2_u14_u6_n111 ) , .B1( u2_u14_u6_n124 ) , .B2( u2_u14_u6_n151 ) , .A2( u2_u14_u6_n93 ) );
  NAND4_X1 u2_u14_u6_U79 (.ZN( u2_out14_12 ) , .A4( u2_u14_u6_n114 ) , .A3( u2_u14_u6_n115 ) , .A2( u2_u14_u6_n116 ) , .A1( u2_u14_u6_n117 ) );
  INV_X1 u2_u14_u6_U8 (.ZN( u2_u14_u6_n172 ) , .A( u2_u14_u6_n88 ) );
  OAI22_X1 u2_u14_u6_U80 (.B2( u2_u14_u6_n111 ) , .ZN( u2_u14_u6_n116 ) , .B1( u2_u14_u6_n126 ) , .A2( u2_u14_u6_n164 ) , .A1( u2_u14_u6_n167 ) );
  OAI21_X1 u2_u14_u6_U81 (.A( u2_u14_u6_n108 ) , .ZN( u2_u14_u6_n117 ) , .B2( u2_u14_u6_n141 ) , .B1( u2_u14_u6_n163 ) );
  OAI211_X1 u2_u14_u6_U82 (.ZN( u2_out14_22 ) , .B( u2_u14_u6_n137 ) , .A( u2_u14_u6_n138 ) , .C2( u2_u14_u6_n139 ) , .C1( u2_u14_u6_n140 ) );
  AOI22_X1 u2_u14_u6_U83 (.B1( u2_u14_u6_n124 ) , .A2( u2_u14_u6_n125 ) , .A1( u2_u14_u6_n126 ) , .ZN( u2_u14_u6_n138 ) , .B2( u2_u14_u6_n161 ) );
  AND4_X1 u2_u14_u6_U84 (.A3( u2_u14_u6_n119 ) , .A1( u2_u14_u6_n120 ) , .A4( u2_u14_u6_n129 ) , .ZN( u2_u14_u6_n140 ) , .A2( u2_u14_u6_n143 ) );
  OAI211_X1 u2_u14_u6_U85 (.ZN( u2_out14_7 ) , .B( u2_u14_u6_n153 ) , .C2( u2_u14_u6_n154 ) , .C1( u2_u14_u6_n155 ) , .A( u2_u14_u6_n174 ) );
  NOR3_X1 u2_u14_u6_U86 (.A1( u2_u14_u6_n141 ) , .ZN( u2_u14_u6_n154 ) , .A3( u2_u14_u6_n164 ) , .A2( u2_u14_u6_n171 ) );
  AOI211_X1 u2_u14_u6_U87 (.B( u2_u14_u6_n149 ) , .A( u2_u14_u6_n150 ) , .C2( u2_u14_u6_n151 ) , .C1( u2_u14_u6_n152 ) , .ZN( u2_u14_u6_n153 ) );
  NAND3_X1 u2_u14_u6_U88 (.A2( u2_u14_u6_n123 ) , .ZN( u2_u14_u6_n125 ) , .A1( u2_u14_u6_n130 ) , .A3( u2_u14_u6_n131 ) );
  NAND3_X1 u2_u14_u6_U89 (.A3( u2_u14_u6_n133 ) , .ZN( u2_u14_u6_n141 ) , .A1( u2_u14_u6_n145 ) , .A2( u2_u14_u6_n148 ) );
  OAI21_X1 u2_u14_u6_U9 (.A( u2_u14_u6_n159 ) , .B1( u2_u14_u6_n169 ) , .B2( u2_u14_u6_n173 ) , .ZN( u2_u14_u6_n90 ) );
  NAND3_X1 u2_u14_u6_U90 (.ZN( u2_u14_u6_n101 ) , .A3( u2_u14_u6_n107 ) , .A2( u2_u14_u6_n121 ) , .A1( u2_u14_u6_n127 ) );
  NAND3_X1 u2_u14_u6_U91 (.ZN( u2_u14_u6_n102 ) , .A3( u2_u14_u6_n130 ) , .A2( u2_u14_u6_n145 ) , .A1( u2_u14_u6_n166 ) );
  NAND3_X1 u2_u14_u6_U92 (.A3( u2_u14_u6_n113 ) , .A1( u2_u14_u6_n119 ) , .A2( u2_u14_u6_n123 ) , .ZN( u2_u14_u6_n93 ) );
  NAND3_X1 u2_u14_u6_U93 (.ZN( u2_u14_u6_n142 ) , .A2( u2_u14_u6_n172 ) , .A3( u2_u14_u6_n89 ) , .A1( u2_u14_u6_n90 ) );
  OAI21_X1 u2_u14_u7_U10 (.A( u2_u14_u7_n161 ) , .B1( u2_u14_u7_n168 ) , .B2( u2_u14_u7_n173 ) , .ZN( u2_u14_u7_n91 ) );
  AOI211_X1 u2_u14_u7_U11 (.A( u2_u14_u7_n117 ) , .ZN( u2_u14_u7_n118 ) , .C2( u2_u14_u7_n126 ) , .C1( u2_u14_u7_n177 ) , .B( u2_u14_u7_n180 ) );
  OAI22_X1 u2_u14_u7_U12 (.B1( u2_u14_u7_n115 ) , .ZN( u2_u14_u7_n117 ) , .A2( u2_u14_u7_n133 ) , .A1( u2_u14_u7_n137 ) , .B2( u2_u14_u7_n162 ) );
  INV_X1 u2_u14_u7_U13 (.A( u2_u14_u7_n116 ) , .ZN( u2_u14_u7_n180 ) );
  NOR3_X1 u2_u14_u7_U14 (.ZN( u2_u14_u7_n115 ) , .A3( u2_u14_u7_n145 ) , .A2( u2_u14_u7_n168 ) , .A1( u2_u14_u7_n169 ) );
  INV_X1 u2_u14_u7_U15 (.A( u2_u14_u7_n133 ) , .ZN( u2_u14_u7_n176 ) );
  NOR3_X1 u2_u14_u7_U16 (.A2( u2_u14_u7_n134 ) , .A1( u2_u14_u7_n135 ) , .ZN( u2_u14_u7_n136 ) , .A3( u2_u14_u7_n171 ) );
  NOR2_X1 u2_u14_u7_U17 (.A1( u2_u14_u7_n130 ) , .A2( u2_u14_u7_n134 ) , .ZN( u2_u14_u7_n153 ) );
  AOI21_X1 u2_u14_u7_U18 (.ZN( u2_u14_u7_n104 ) , .B2( u2_u14_u7_n112 ) , .B1( u2_u14_u7_n127 ) , .A( u2_u14_u7_n164 ) );
  AOI21_X1 u2_u14_u7_U19 (.ZN( u2_u14_u7_n106 ) , .B1( u2_u14_u7_n133 ) , .B2( u2_u14_u7_n146 ) , .A( u2_u14_u7_n162 ) );
  AOI21_X1 u2_u14_u7_U20 (.A( u2_u14_u7_n101 ) , .ZN( u2_u14_u7_n107 ) , .B2( u2_u14_u7_n128 ) , .B1( u2_u14_u7_n175 ) );
  INV_X1 u2_u14_u7_U21 (.A( u2_u14_u7_n101 ) , .ZN( u2_u14_u7_n165 ) );
  NOR2_X1 u2_u14_u7_U22 (.ZN( u2_u14_u7_n111 ) , .A2( u2_u14_u7_n134 ) , .A1( u2_u14_u7_n169 ) );
  INV_X1 u2_u14_u7_U23 (.A( u2_u14_u7_n138 ) , .ZN( u2_u14_u7_n171 ) );
  INV_X1 u2_u14_u7_U24 (.A( u2_u14_u7_n131 ) , .ZN( u2_u14_u7_n177 ) );
  INV_X1 u2_u14_u7_U25 (.A( u2_u14_u7_n110 ) , .ZN( u2_u14_u7_n174 ) );
  NAND2_X1 u2_u14_u7_U26 (.A1( u2_u14_u7_n129 ) , .A2( u2_u14_u7_n132 ) , .ZN( u2_u14_u7_n149 ) );
  NAND2_X1 u2_u14_u7_U27 (.A1( u2_u14_u7_n113 ) , .A2( u2_u14_u7_n124 ) , .ZN( u2_u14_u7_n130 ) );
  INV_X1 u2_u14_u7_U28 (.A( u2_u14_u7_n112 ) , .ZN( u2_u14_u7_n173 ) );
  INV_X1 u2_u14_u7_U29 (.A( u2_u14_u7_n128 ) , .ZN( u2_u14_u7_n168 ) );
  OAI21_X1 u2_u14_u7_U3 (.ZN( u2_u14_u7_n159 ) , .A( u2_u14_u7_n165 ) , .B2( u2_u14_u7_n171 ) , .B1( u2_u14_u7_n174 ) );
  INV_X1 u2_u14_u7_U30 (.A( u2_u14_u7_n148 ) , .ZN( u2_u14_u7_n169 ) );
  INV_X1 u2_u14_u7_U31 (.A( u2_u14_u7_n127 ) , .ZN( u2_u14_u7_n179 ) );
  NOR2_X1 u2_u14_u7_U32 (.ZN( u2_u14_u7_n101 ) , .A2( u2_u14_u7_n150 ) , .A1( u2_u14_u7_n156 ) );
  AOI211_X1 u2_u14_u7_U33 (.B( u2_u14_u7_n139 ) , .A( u2_u14_u7_n140 ) , .C2( u2_u14_u7_n141 ) , .ZN( u2_u14_u7_n142 ) , .C1( u2_u14_u7_n156 ) );
  NAND4_X1 u2_u14_u7_U34 (.A3( u2_u14_u7_n127 ) , .A2( u2_u14_u7_n128 ) , .A1( u2_u14_u7_n129 ) , .ZN( u2_u14_u7_n141 ) , .A4( u2_u14_u7_n147 ) );
  AOI21_X1 u2_u14_u7_U35 (.A( u2_u14_u7_n137 ) , .B1( u2_u14_u7_n138 ) , .ZN( u2_u14_u7_n139 ) , .B2( u2_u14_u7_n146 ) );
  OAI22_X1 u2_u14_u7_U36 (.B1( u2_u14_u7_n136 ) , .ZN( u2_u14_u7_n140 ) , .A1( u2_u14_u7_n153 ) , .B2( u2_u14_u7_n162 ) , .A2( u2_u14_u7_n164 ) );
  INV_X1 u2_u14_u7_U37 (.A( u2_u14_u7_n125 ) , .ZN( u2_u14_u7_n161 ) );
  AOI21_X1 u2_u14_u7_U38 (.ZN( u2_u14_u7_n123 ) , .B1( u2_u14_u7_n165 ) , .B2( u2_u14_u7_n177 ) , .A( u2_u14_u7_n97 ) );
  AOI21_X1 u2_u14_u7_U39 (.B2( u2_u14_u7_n113 ) , .B1( u2_u14_u7_n124 ) , .A( u2_u14_u7_n125 ) , .ZN( u2_u14_u7_n97 ) );
  INV_X1 u2_u14_u7_U4 (.A( u2_u14_u7_n149 ) , .ZN( u2_u14_u7_n175 ) );
  INV_X1 u2_u14_u7_U40 (.A( u2_u14_u7_n152 ) , .ZN( u2_u14_u7_n162 ) );
  AOI22_X1 u2_u14_u7_U41 (.A2( u2_u14_u7_n114 ) , .ZN( u2_u14_u7_n119 ) , .B1( u2_u14_u7_n130 ) , .A1( u2_u14_u7_n156 ) , .B2( u2_u14_u7_n165 ) );
  NAND2_X1 u2_u14_u7_U42 (.A2( u2_u14_u7_n112 ) , .ZN( u2_u14_u7_n114 ) , .A1( u2_u14_u7_n175 ) );
  NOR2_X1 u2_u14_u7_U43 (.ZN( u2_u14_u7_n137 ) , .A1( u2_u14_u7_n150 ) , .A2( u2_u14_u7_n161 ) );
  AND2_X1 u2_u14_u7_U44 (.ZN( u2_u14_u7_n145 ) , .A2( u2_u14_u7_n98 ) , .A1( u2_u14_u7_n99 ) );
  AOI21_X1 u2_u14_u7_U45 (.ZN( u2_u14_u7_n105 ) , .B2( u2_u14_u7_n110 ) , .A( u2_u14_u7_n125 ) , .B1( u2_u14_u7_n147 ) );
  NAND2_X1 u2_u14_u7_U46 (.ZN( u2_u14_u7_n146 ) , .A1( u2_u14_u7_n95 ) , .A2( u2_u14_u7_n98 ) );
  NAND2_X1 u2_u14_u7_U47 (.A2( u2_u14_u7_n103 ) , .ZN( u2_u14_u7_n147 ) , .A1( u2_u14_u7_n93 ) );
  NAND2_X1 u2_u14_u7_U48 (.A1( u2_u14_u7_n103 ) , .ZN( u2_u14_u7_n127 ) , .A2( u2_u14_u7_n99 ) );
  NAND2_X1 u2_u14_u7_U49 (.A2( u2_u14_u7_n102 ) , .A1( u2_u14_u7_n103 ) , .ZN( u2_u14_u7_n133 ) );
  INV_X1 u2_u14_u7_U5 (.A( u2_u14_u7_n154 ) , .ZN( u2_u14_u7_n178 ) );
  OR2_X1 u2_u14_u7_U50 (.ZN( u2_u14_u7_n126 ) , .A2( u2_u14_u7_n152 ) , .A1( u2_u14_u7_n156 ) );
  NAND2_X1 u2_u14_u7_U51 (.ZN( u2_u14_u7_n112 ) , .A2( u2_u14_u7_n96 ) , .A1( u2_u14_u7_n99 ) );
  NAND2_X1 u2_u14_u7_U52 (.A2( u2_u14_u7_n102 ) , .ZN( u2_u14_u7_n128 ) , .A1( u2_u14_u7_n98 ) );
  NAND2_X1 u2_u14_u7_U53 (.A1( u2_u14_u7_n100 ) , .ZN( u2_u14_u7_n113 ) , .A2( u2_u14_u7_n93 ) );
  NAND2_X1 u2_u14_u7_U54 (.ZN( u2_u14_u7_n110 ) , .A1( u2_u14_u7_n95 ) , .A2( u2_u14_u7_n96 ) );
  INV_X1 u2_u14_u7_U55 (.A( u2_u14_u7_n150 ) , .ZN( u2_u14_u7_n164 ) );
  AND2_X1 u2_u14_u7_U56 (.ZN( u2_u14_u7_n134 ) , .A1( u2_u14_u7_n93 ) , .A2( u2_u14_u7_n98 ) );
  NAND2_X1 u2_u14_u7_U57 (.A2( u2_u14_u7_n102 ) , .ZN( u2_u14_u7_n124 ) , .A1( u2_u14_u7_n96 ) );
  NAND2_X1 u2_u14_u7_U58 (.A1( u2_u14_u7_n100 ) , .A2( u2_u14_u7_n102 ) , .ZN( u2_u14_u7_n129 ) );
  NAND2_X1 u2_u14_u7_U59 (.A2( u2_u14_u7_n103 ) , .ZN( u2_u14_u7_n131 ) , .A1( u2_u14_u7_n95 ) );
  AOI211_X1 u2_u14_u7_U6 (.ZN( u2_u14_u7_n116 ) , .A( u2_u14_u7_n155 ) , .C1( u2_u14_u7_n161 ) , .C2( u2_u14_u7_n171 ) , .B( u2_u14_u7_n94 ) );
  NAND2_X1 u2_u14_u7_U60 (.A1( u2_u14_u7_n100 ) , .ZN( u2_u14_u7_n138 ) , .A2( u2_u14_u7_n99 ) );
  NAND2_X1 u2_u14_u7_U61 (.ZN( u2_u14_u7_n132 ) , .A1( u2_u14_u7_n93 ) , .A2( u2_u14_u7_n96 ) );
  NAND2_X1 u2_u14_u7_U62 (.A1( u2_u14_u7_n100 ) , .ZN( u2_u14_u7_n148 ) , .A2( u2_u14_u7_n95 ) );
  AOI211_X1 u2_u14_u7_U63 (.B( u2_u14_u7_n154 ) , .A( u2_u14_u7_n155 ) , .C1( u2_u14_u7_n156 ) , .ZN( u2_u14_u7_n157 ) , .C2( u2_u14_u7_n172 ) );
  INV_X1 u2_u14_u7_U64 (.A( u2_u14_u7_n153 ) , .ZN( u2_u14_u7_n172 ) );
  NOR2_X1 u2_u14_u7_U65 (.A2( u2_u14_X_47 ) , .ZN( u2_u14_u7_n150 ) , .A1( u2_u14_u7_n163 ) );
  NOR2_X1 u2_u14_u7_U66 (.A2( u2_u14_X_43 ) , .A1( u2_u14_X_44 ) , .ZN( u2_u14_u7_n103 ) );
  NOR2_X1 u2_u14_u7_U67 (.A2( u2_u14_X_48 ) , .A1( u2_u14_u7_n166 ) , .ZN( u2_u14_u7_n95 ) );
  NOR2_X1 u2_u14_u7_U68 (.A2( u2_u14_X_45 ) , .A1( u2_u14_X_48 ) , .ZN( u2_u14_u7_n99 ) );
  NOR2_X1 u2_u14_u7_U69 (.A2( u2_u14_X_44 ) , .A1( u2_u14_u7_n167 ) , .ZN( u2_u14_u7_n98 ) );
  OAI222_X1 u2_u14_u7_U7 (.C2( u2_u14_u7_n101 ) , .B2( u2_u14_u7_n111 ) , .A1( u2_u14_u7_n113 ) , .C1( u2_u14_u7_n146 ) , .A2( u2_u14_u7_n162 ) , .B1( u2_u14_u7_n164 ) , .ZN( u2_u14_u7_n94 ) );
  NOR2_X1 u2_u14_u7_U70 (.A2( u2_u14_X_46 ) , .A1( u2_u14_X_47 ) , .ZN( u2_u14_u7_n152 ) );
  NAND2_X1 u2_u14_u7_U71 (.A2( u2_u14_X_46 ) , .A1( u2_u14_X_47 ) , .ZN( u2_u14_u7_n125 ) );
  AND2_X1 u2_u14_u7_U72 (.A1( u2_u14_X_47 ) , .ZN( u2_u14_u7_n156 ) , .A2( u2_u14_u7_n163 ) );
  AND2_X1 u2_u14_u7_U73 (.A2( u2_u14_X_45 ) , .A1( u2_u14_X_48 ) , .ZN( u2_u14_u7_n102 ) );
  AND2_X1 u2_u14_u7_U74 (.A2( u2_u14_X_43 ) , .A1( u2_u14_X_44 ) , .ZN( u2_u14_u7_n96 ) );
  AND2_X1 u2_u14_u7_U75 (.A1( u2_u14_X_44 ) , .ZN( u2_u14_u7_n100 ) , .A2( u2_u14_u7_n167 ) );
  AND2_X1 u2_u14_u7_U76 (.A1( u2_u14_X_48 ) , .A2( u2_u14_u7_n166 ) , .ZN( u2_u14_u7_n93 ) );
  INV_X1 u2_u14_u7_U77 (.A( u2_u14_X_46 ) , .ZN( u2_u14_u7_n163 ) );
  INV_X1 u2_u14_u7_U78 (.A( u2_u14_X_45 ) , .ZN( u2_u14_u7_n166 ) );
  INV_X1 u2_u14_u7_U79 (.A( u2_u14_X_43 ) , .ZN( u2_u14_u7_n167 ) );
  OAI221_X1 u2_u14_u7_U8 (.C1( u2_u14_u7_n101 ) , .C2( u2_u14_u7_n147 ) , .ZN( u2_u14_u7_n155 ) , .B2( u2_u14_u7_n162 ) , .A( u2_u14_u7_n91 ) , .B1( u2_u14_u7_n92 ) );
  NAND4_X1 u2_u14_u7_U80 (.ZN( u2_out14_27 ) , .A4( u2_u14_u7_n118 ) , .A3( u2_u14_u7_n119 ) , .A2( u2_u14_u7_n120 ) , .A1( u2_u14_u7_n121 ) );
  OAI21_X1 u2_u14_u7_U81 (.ZN( u2_u14_u7_n121 ) , .B2( u2_u14_u7_n145 ) , .A( u2_u14_u7_n150 ) , .B1( u2_u14_u7_n174 ) );
  OAI21_X1 u2_u14_u7_U82 (.ZN( u2_u14_u7_n120 ) , .A( u2_u14_u7_n161 ) , .B2( u2_u14_u7_n170 ) , .B1( u2_u14_u7_n179 ) );
  NAND4_X1 u2_u14_u7_U83 (.ZN( u2_out14_21 ) , .A4( u2_u14_u7_n157 ) , .A3( u2_u14_u7_n158 ) , .A2( u2_u14_u7_n159 ) , .A1( u2_u14_u7_n160 ) );
  OAI21_X1 u2_u14_u7_U84 (.B1( u2_u14_u7_n145 ) , .ZN( u2_u14_u7_n160 ) , .A( u2_u14_u7_n161 ) , .B2( u2_u14_u7_n177 ) );
  AOI22_X1 u2_u14_u7_U85 (.B2( u2_u14_u7_n149 ) , .B1( u2_u14_u7_n150 ) , .A2( u2_u14_u7_n151 ) , .A1( u2_u14_u7_n152 ) , .ZN( u2_u14_u7_n158 ) );
  NAND4_X1 u2_u14_u7_U86 (.ZN( u2_out14_15 ) , .A4( u2_u14_u7_n142 ) , .A3( u2_u14_u7_n143 ) , .A2( u2_u14_u7_n144 ) , .A1( u2_u14_u7_n178 ) );
  OR2_X1 u2_u14_u7_U87 (.A2( u2_u14_u7_n125 ) , .A1( u2_u14_u7_n129 ) , .ZN( u2_u14_u7_n144 ) );
  AOI22_X1 u2_u14_u7_U88 (.A2( u2_u14_u7_n126 ) , .ZN( u2_u14_u7_n143 ) , .B2( u2_u14_u7_n165 ) , .B1( u2_u14_u7_n173 ) , .A1( u2_u14_u7_n174 ) );
  NAND4_X1 u2_u14_u7_U89 (.ZN( u2_out14_5 ) , .A4( u2_u14_u7_n108 ) , .A3( u2_u14_u7_n109 ) , .A1( u2_u14_u7_n116 ) , .A2( u2_u14_u7_n123 ) );
  AND3_X1 u2_u14_u7_U9 (.A3( u2_u14_u7_n110 ) , .A2( u2_u14_u7_n127 ) , .A1( u2_u14_u7_n132 ) , .ZN( u2_u14_u7_n92 ) );
  AOI22_X1 u2_u14_u7_U90 (.ZN( u2_u14_u7_n109 ) , .A2( u2_u14_u7_n126 ) , .B2( u2_u14_u7_n145 ) , .B1( u2_u14_u7_n156 ) , .A1( u2_u14_u7_n171 ) );
  NOR4_X1 u2_u14_u7_U91 (.A4( u2_u14_u7_n104 ) , .A3( u2_u14_u7_n105 ) , .A2( u2_u14_u7_n106 ) , .A1( u2_u14_u7_n107 ) , .ZN( u2_u14_u7_n108 ) );
  OAI211_X1 u2_u14_u7_U92 (.B( u2_u14_u7_n122 ) , .A( u2_u14_u7_n123 ) , .C2( u2_u14_u7_n124 ) , .ZN( u2_u14_u7_n154 ) , .C1( u2_u14_u7_n162 ) );
  AOI222_X1 u2_u14_u7_U93 (.ZN( u2_u14_u7_n122 ) , .C2( u2_u14_u7_n126 ) , .C1( u2_u14_u7_n145 ) , .B1( u2_u14_u7_n161 ) , .A2( u2_u14_u7_n165 ) , .B2( u2_u14_u7_n170 ) , .A1( u2_u14_u7_n176 ) );
  INV_X1 u2_u14_u7_U94 (.A( u2_u14_u7_n111 ) , .ZN( u2_u14_u7_n170 ) );
  NAND3_X1 u2_u14_u7_U95 (.A3( u2_u14_u7_n146 ) , .A2( u2_u14_u7_n147 ) , .A1( u2_u14_u7_n148 ) , .ZN( u2_u14_u7_n151 ) );
  NAND3_X1 u2_u14_u7_U96 (.A3( u2_u14_u7_n131 ) , .A2( u2_u14_u7_n132 ) , .A1( u2_u14_u7_n133 ) , .ZN( u2_u14_u7_n135 ) );
  XOR2_X1 u2_u2_U1 (.B( u2_K3_9 ) , .A( u2_R1_6 ) , .Z( u2_u2_X_9 ) );
  XOR2_X1 u2_u2_U10 (.B( u2_K3_45 ) , .A( u2_R1_30 ) , .Z( u2_u2_X_45 ) );
  XOR2_X1 u2_u2_U11 (.B( u2_K3_44 ) , .A( u2_R1_29 ) , .Z( u2_u2_X_44 ) );
  XOR2_X1 u2_u2_U12 (.B( u2_K3_43 ) , .A( u2_R1_28 ) , .Z( u2_u2_X_43 ) );
  XOR2_X1 u2_u2_U13 (.B( u2_K3_42 ) , .A( u2_R1_29 ) , .Z( u2_u2_X_42 ) );
  XOR2_X1 u2_u2_U14 (.B( u2_K3_41 ) , .A( u2_R1_28 ) , .Z( u2_u2_X_41 ) );
  XOR2_X1 u2_u2_U15 (.B( u2_K3_40 ) , .A( u2_R1_27 ) , .Z( u2_u2_X_40 ) );
  XOR2_X1 u2_u2_U16 (.B( u2_K3_3 ) , .A( u2_R1_2 ) , .Z( u2_u2_X_3 ) );
  XOR2_X1 u2_u2_U18 (.B( u2_K3_38 ) , .A( u2_R1_25 ) , .Z( u2_u2_X_38 ) );
  XOR2_X1 u2_u2_U2 (.B( u2_K3_8 ) , .A( u2_R1_5 ) , .Z( u2_u2_X_8 ) );
  XOR2_X1 u2_u2_U20 (.B( u2_K3_36 ) , .A( u2_R1_25 ) , .Z( u2_u2_X_36 ) );
  XOR2_X1 u2_u2_U27 (.B( u2_K3_2 ) , .A( u2_R1_1 ) , .Z( u2_u2_X_2 ) );
  XOR2_X1 u2_u2_U31 (.B( u2_K3_26 ) , .A( u2_R1_17 ) , .Z( u2_u2_X_26 ) );
  XOR2_X1 u2_u2_U32 (.B( u2_K3_25 ) , .A( u2_R1_16 ) , .Z( u2_u2_X_25 ) );
  XOR2_X1 u2_u2_U33 (.B( u2_K3_24 ) , .A( u2_R1_17 ) , .Z( u2_u2_X_24 ) );
  XOR2_X1 u2_u2_U34 (.B( u2_K3_23 ) , .A( u2_R1_16 ) , .Z( u2_u2_X_23 ) );
  XOR2_X1 u2_u2_U35 (.B( u2_K3_22 ) , .A( u2_R1_15 ) , .Z( u2_u2_X_22 ) );
  XOR2_X1 u2_u2_U36 (.B( u2_K3_21 ) , .A( u2_R1_14 ) , .Z( u2_u2_X_21 ) );
  XOR2_X1 u2_u2_U37 (.B( u2_K3_20 ) , .A( u2_R1_13 ) , .Z( u2_u2_X_20 ) );
  XOR2_X1 u2_u2_U38 (.B( u2_K3_1 ) , .A( u2_R1_32 ) , .Z( u2_u2_X_1 ) );
  XOR2_X1 u2_u2_U39 (.B( u2_K3_19 ) , .A( u2_R1_12 ) , .Z( u2_u2_X_19 ) );
  XOR2_X1 u2_u2_U4 (.B( u2_K3_6 ) , .A( u2_R1_5 ) , .Z( u2_u2_X_6 ) );
  XOR2_X1 u2_u2_U40 (.B( u2_K3_18 ) , .A( u2_R1_13 ) , .Z( u2_u2_X_18 ) );
  XOR2_X1 u2_u2_U41 (.B( u2_K3_17 ) , .A( u2_R1_12 ) , .Z( u2_u2_X_17 ) );
  XOR2_X1 u2_u2_U44 (.B( u2_K3_14 ) , .A( u2_R1_9 ) , .Z( u2_u2_X_14 ) );
  XOR2_X1 u2_u2_U45 (.B( u2_K3_13 ) , .A( u2_R1_8 ) , .Z( u2_u2_X_13 ) );
  XOR2_X1 u2_u2_U46 (.B( u2_K3_12 ) , .A( u2_R1_9 ) , .Z( u2_u2_X_12 ) );
  XOR2_X1 u2_u2_U47 (.B( u2_K3_11 ) , .A( u2_R1_8 ) , .Z( u2_u2_X_11 ) );
  XOR2_X1 u2_u2_U48 (.B( u2_K3_10 ) , .A( u2_R1_7 ) , .Z( u2_u2_X_10 ) );
  XOR2_X1 u2_u2_U6 (.B( u2_K3_4 ) , .A( u2_R1_3 ) , .Z( u2_u2_X_4 ) );
  XOR2_X1 u2_u2_U7 (.B( u2_K3_48 ) , .A( u2_R1_1 ) , .Z( u2_u2_X_48 ) );
  XOR2_X1 u2_u2_U8 (.B( u2_K3_47 ) , .A( u2_R1_32 ) , .Z( u2_u2_X_47 ) );
  XOR2_X1 u2_u2_U9 (.B( u2_K3_46 ) , .A( u2_R1_31 ) , .Z( u2_u2_X_46 ) );
  AND3_X1 u2_u2_u0_U10 (.A2( u2_u2_u0_n112 ) , .ZN( u2_u2_u0_n127 ) , .A3( u2_u2_u0_n130 ) , .A1( u2_u2_u0_n148 ) );
  NAND2_X1 u2_u2_u0_U11 (.ZN( u2_u2_u0_n113 ) , .A1( u2_u2_u0_n139 ) , .A2( u2_u2_u0_n149 ) );
  AND2_X1 u2_u2_u0_U12 (.ZN( u2_u2_u0_n107 ) , .A1( u2_u2_u0_n130 ) , .A2( u2_u2_u0_n140 ) );
  AND2_X1 u2_u2_u0_U13 (.A2( u2_u2_u0_n129 ) , .A1( u2_u2_u0_n130 ) , .ZN( u2_u2_u0_n151 ) );
  AND2_X1 u2_u2_u0_U14 (.A1( u2_u2_u0_n108 ) , .A2( u2_u2_u0_n125 ) , .ZN( u2_u2_u0_n145 ) );
  INV_X1 u2_u2_u0_U15 (.A( u2_u2_u0_n143 ) , .ZN( u2_u2_u0_n173 ) );
  NOR2_X1 u2_u2_u0_U16 (.A2( u2_u2_u0_n136 ) , .ZN( u2_u2_u0_n147 ) , .A1( u2_u2_u0_n160 ) );
  INV_X1 u2_u2_u0_U17 (.ZN( u2_u2_u0_n172 ) , .A( u2_u2_u0_n88 ) );
  OAI222_X1 u2_u2_u0_U18 (.C1( u2_u2_u0_n108 ) , .A1( u2_u2_u0_n125 ) , .B2( u2_u2_u0_n128 ) , .B1( u2_u2_u0_n144 ) , .A2( u2_u2_u0_n158 ) , .C2( u2_u2_u0_n161 ) , .ZN( u2_u2_u0_n88 ) );
  NOR2_X1 u2_u2_u0_U19 (.A1( u2_u2_u0_n163 ) , .A2( u2_u2_u0_n164 ) , .ZN( u2_u2_u0_n95 ) );
  AOI21_X1 u2_u2_u0_U20 (.B1( u2_u2_u0_n103 ) , .ZN( u2_u2_u0_n132 ) , .A( u2_u2_u0_n165 ) , .B2( u2_u2_u0_n93 ) );
  INV_X1 u2_u2_u0_U21 (.A( u2_u2_u0_n142 ) , .ZN( u2_u2_u0_n165 ) );
  OAI221_X1 u2_u2_u0_U22 (.C1( u2_u2_u0_n121 ) , .ZN( u2_u2_u0_n122 ) , .B2( u2_u2_u0_n127 ) , .A( u2_u2_u0_n143 ) , .B1( u2_u2_u0_n144 ) , .C2( u2_u2_u0_n147 ) );
  OAI22_X1 u2_u2_u0_U23 (.B1( u2_u2_u0_n125 ) , .ZN( u2_u2_u0_n126 ) , .A1( u2_u2_u0_n138 ) , .A2( u2_u2_u0_n146 ) , .B2( u2_u2_u0_n147 ) );
  OAI22_X1 u2_u2_u0_U24 (.B1( u2_u2_u0_n131 ) , .A1( u2_u2_u0_n144 ) , .B2( u2_u2_u0_n147 ) , .A2( u2_u2_u0_n90 ) , .ZN( u2_u2_u0_n91 ) );
  AND3_X1 u2_u2_u0_U25 (.A3( u2_u2_u0_n121 ) , .A2( u2_u2_u0_n125 ) , .A1( u2_u2_u0_n148 ) , .ZN( u2_u2_u0_n90 ) );
  INV_X1 u2_u2_u0_U26 (.A( u2_u2_u0_n136 ) , .ZN( u2_u2_u0_n161 ) );
  NOR2_X1 u2_u2_u0_U27 (.A1( u2_u2_u0_n120 ) , .ZN( u2_u2_u0_n143 ) , .A2( u2_u2_u0_n167 ) );
  OAI221_X1 u2_u2_u0_U28 (.C1( u2_u2_u0_n112 ) , .ZN( u2_u2_u0_n120 ) , .B1( u2_u2_u0_n138 ) , .B2( u2_u2_u0_n141 ) , .C2( u2_u2_u0_n147 ) , .A( u2_u2_u0_n172 ) );
  AOI211_X1 u2_u2_u0_U29 (.B( u2_u2_u0_n115 ) , .A( u2_u2_u0_n116 ) , .C2( u2_u2_u0_n117 ) , .C1( u2_u2_u0_n118 ) , .ZN( u2_u2_u0_n119 ) );
  INV_X1 u2_u2_u0_U3 (.A( u2_u2_u0_n113 ) , .ZN( u2_u2_u0_n166 ) );
  AOI22_X1 u2_u2_u0_U30 (.B2( u2_u2_u0_n109 ) , .A2( u2_u2_u0_n110 ) , .ZN( u2_u2_u0_n111 ) , .B1( u2_u2_u0_n118 ) , .A1( u2_u2_u0_n160 ) );
  INV_X1 u2_u2_u0_U31 (.A( u2_u2_u0_n118 ) , .ZN( u2_u2_u0_n158 ) );
  AOI21_X1 u2_u2_u0_U32 (.ZN( u2_u2_u0_n104 ) , .B1( u2_u2_u0_n107 ) , .B2( u2_u2_u0_n141 ) , .A( u2_u2_u0_n144 ) );
  AOI21_X1 u2_u2_u0_U33 (.B1( u2_u2_u0_n127 ) , .B2( u2_u2_u0_n129 ) , .A( u2_u2_u0_n138 ) , .ZN( u2_u2_u0_n96 ) );
  AOI21_X1 u2_u2_u0_U34 (.ZN( u2_u2_u0_n116 ) , .B2( u2_u2_u0_n142 ) , .A( u2_u2_u0_n144 ) , .B1( u2_u2_u0_n166 ) );
  NAND2_X1 u2_u2_u0_U35 (.A1( u2_u2_u0_n100 ) , .A2( u2_u2_u0_n103 ) , .ZN( u2_u2_u0_n125 ) );
  NAND2_X1 u2_u2_u0_U36 (.A1( u2_u2_u0_n101 ) , .A2( u2_u2_u0_n102 ) , .ZN( u2_u2_u0_n150 ) );
  INV_X1 u2_u2_u0_U37 (.A( u2_u2_u0_n138 ) , .ZN( u2_u2_u0_n160 ) );
  NAND2_X1 u2_u2_u0_U38 (.A1( u2_u2_u0_n102 ) , .ZN( u2_u2_u0_n128 ) , .A2( u2_u2_u0_n95 ) );
  NAND2_X1 u2_u2_u0_U39 (.A1( u2_u2_u0_n100 ) , .ZN( u2_u2_u0_n129 ) , .A2( u2_u2_u0_n95 ) );
  AOI21_X1 u2_u2_u0_U4 (.B1( u2_u2_u0_n114 ) , .ZN( u2_u2_u0_n115 ) , .B2( u2_u2_u0_n129 ) , .A( u2_u2_u0_n161 ) );
  NAND2_X1 u2_u2_u0_U40 (.A2( u2_u2_u0_n100 ) , .ZN( u2_u2_u0_n131 ) , .A1( u2_u2_u0_n92 ) );
  NAND2_X1 u2_u2_u0_U41 (.A2( u2_u2_u0_n100 ) , .A1( u2_u2_u0_n101 ) , .ZN( u2_u2_u0_n139 ) );
  NAND2_X1 u2_u2_u0_U42 (.ZN( u2_u2_u0_n148 ) , .A1( u2_u2_u0_n93 ) , .A2( u2_u2_u0_n95 ) );
  NAND2_X1 u2_u2_u0_U43 (.A2( u2_u2_u0_n102 ) , .A1( u2_u2_u0_n103 ) , .ZN( u2_u2_u0_n149 ) );
  NAND2_X1 u2_u2_u0_U44 (.A2( u2_u2_u0_n102 ) , .ZN( u2_u2_u0_n114 ) , .A1( u2_u2_u0_n92 ) );
  NAND2_X1 u2_u2_u0_U45 (.A2( u2_u2_u0_n101 ) , .ZN( u2_u2_u0_n121 ) , .A1( u2_u2_u0_n93 ) );
  NAND2_X1 u2_u2_u0_U46 (.ZN( u2_u2_u0_n112 ) , .A2( u2_u2_u0_n92 ) , .A1( u2_u2_u0_n93 ) );
  OR3_X1 u2_u2_u0_U47 (.A3( u2_u2_u0_n152 ) , .A2( u2_u2_u0_n153 ) , .A1( u2_u2_u0_n154 ) , .ZN( u2_u2_u0_n155 ) );
  AOI21_X1 u2_u2_u0_U48 (.B2( u2_u2_u0_n150 ) , .B1( u2_u2_u0_n151 ) , .ZN( u2_u2_u0_n152 ) , .A( u2_u2_u0_n158 ) );
  AOI21_X1 u2_u2_u0_U49 (.A( u2_u2_u0_n144 ) , .B2( u2_u2_u0_n145 ) , .B1( u2_u2_u0_n146 ) , .ZN( u2_u2_u0_n154 ) );
  AOI21_X1 u2_u2_u0_U5 (.B2( u2_u2_u0_n131 ) , .ZN( u2_u2_u0_n134 ) , .B1( u2_u2_u0_n151 ) , .A( u2_u2_u0_n158 ) );
  AOI21_X1 u2_u2_u0_U50 (.A( u2_u2_u0_n147 ) , .B2( u2_u2_u0_n148 ) , .B1( u2_u2_u0_n149 ) , .ZN( u2_u2_u0_n153 ) );
  INV_X1 u2_u2_u0_U51 (.ZN( u2_u2_u0_n171 ) , .A( u2_u2_u0_n99 ) );
  OAI211_X1 u2_u2_u0_U52 (.C2( u2_u2_u0_n140 ) , .C1( u2_u2_u0_n161 ) , .A( u2_u2_u0_n169 ) , .B( u2_u2_u0_n98 ) , .ZN( u2_u2_u0_n99 ) );
  INV_X1 u2_u2_u0_U53 (.ZN( u2_u2_u0_n169 ) , .A( u2_u2_u0_n91 ) );
  AOI211_X1 u2_u2_u0_U54 (.C1( u2_u2_u0_n118 ) , .A( u2_u2_u0_n123 ) , .B( u2_u2_u0_n96 ) , .C2( u2_u2_u0_n97 ) , .ZN( u2_u2_u0_n98 ) );
  NOR2_X1 u2_u2_u0_U55 (.A2( u2_u2_X_6 ) , .ZN( u2_u2_u0_n100 ) , .A1( u2_u2_u0_n162 ) );
  NOR2_X1 u2_u2_u0_U56 (.A2( u2_u2_X_4 ) , .A1( u2_u2_X_5 ) , .ZN( u2_u2_u0_n118 ) );
  NOR2_X1 u2_u2_u0_U57 (.A2( u2_u2_X_2 ) , .ZN( u2_u2_u0_n103 ) , .A1( u2_u2_u0_n164 ) );
  NOR2_X1 u2_u2_u0_U58 (.A2( u2_u2_X_1 ) , .A1( u2_u2_X_2 ) , .ZN( u2_u2_u0_n92 ) );
  NOR2_X1 u2_u2_u0_U59 (.A2( u2_u2_X_1 ) , .ZN( u2_u2_u0_n101 ) , .A1( u2_u2_u0_n163 ) );
  NOR2_X1 u2_u2_u0_U6 (.A1( u2_u2_u0_n108 ) , .ZN( u2_u2_u0_n123 ) , .A2( u2_u2_u0_n158 ) );
  NAND2_X1 u2_u2_u0_U60 (.A2( u2_u2_X_4 ) , .A1( u2_u2_X_5 ) , .ZN( u2_u2_u0_n144 ) );
  NOR2_X1 u2_u2_u0_U61 (.A2( u2_u2_X_5 ) , .ZN( u2_u2_u0_n136 ) , .A1( u2_u2_u0_n159 ) );
  NAND2_X1 u2_u2_u0_U62 (.A1( u2_u2_X_5 ) , .ZN( u2_u2_u0_n138 ) , .A2( u2_u2_u0_n159 ) );
  NOR2_X1 u2_u2_u0_U63 (.A2( u2_u2_X_3 ) , .A1( u2_u2_X_6 ) , .ZN( u2_u2_u0_n94 ) );
  AND2_X1 u2_u2_u0_U64 (.A2( u2_u2_X_3 ) , .A1( u2_u2_X_6 ) , .ZN( u2_u2_u0_n102 ) );
  AND2_X1 u2_u2_u0_U65 (.A1( u2_u2_X_6 ) , .A2( u2_u2_u0_n162 ) , .ZN( u2_u2_u0_n93 ) );
  INV_X1 u2_u2_u0_U66 (.A( u2_u2_X_4 ) , .ZN( u2_u2_u0_n159 ) );
  INV_X1 u2_u2_u0_U67 (.A( u2_u2_X_1 ) , .ZN( u2_u2_u0_n164 ) );
  INV_X1 u2_u2_u0_U68 (.A( u2_u2_X_2 ) , .ZN( u2_u2_u0_n163 ) );
  INV_X1 u2_u2_u0_U69 (.A( u2_u2_X_3 ) , .ZN( u2_u2_u0_n162 ) );
  OAI21_X1 u2_u2_u0_U7 (.B1( u2_u2_u0_n150 ) , .B2( u2_u2_u0_n158 ) , .A( u2_u2_u0_n172 ) , .ZN( u2_u2_u0_n89 ) );
  INV_X1 u2_u2_u0_U70 (.A( u2_u2_u0_n126 ) , .ZN( u2_u2_u0_n168 ) );
  AOI211_X1 u2_u2_u0_U71 (.B( u2_u2_u0_n133 ) , .A( u2_u2_u0_n134 ) , .C2( u2_u2_u0_n135 ) , .C1( u2_u2_u0_n136 ) , .ZN( u2_u2_u0_n137 ) );
  INV_X1 u2_u2_u0_U72 (.ZN( u2_u2_u0_n174 ) , .A( u2_u2_u0_n89 ) );
  AOI211_X1 u2_u2_u0_U73 (.B( u2_u2_u0_n104 ) , .A( u2_u2_u0_n105 ) , .ZN( u2_u2_u0_n106 ) , .C2( u2_u2_u0_n113 ) , .C1( u2_u2_u0_n160 ) );
  OR4_X1 u2_u2_u0_U74 (.ZN( u2_out2_17 ) , .A4( u2_u2_u0_n122 ) , .A2( u2_u2_u0_n123 ) , .A1( u2_u2_u0_n124 ) , .A3( u2_u2_u0_n170 ) );
  AOI21_X1 u2_u2_u0_U75 (.B2( u2_u2_u0_n107 ) , .ZN( u2_u2_u0_n124 ) , .B1( u2_u2_u0_n128 ) , .A( u2_u2_u0_n161 ) );
  INV_X1 u2_u2_u0_U76 (.A( u2_u2_u0_n111 ) , .ZN( u2_u2_u0_n170 ) );
  OR4_X1 u2_u2_u0_U77 (.ZN( u2_out2_31 ) , .A4( u2_u2_u0_n155 ) , .A2( u2_u2_u0_n156 ) , .A1( u2_u2_u0_n157 ) , .A3( u2_u2_u0_n173 ) );
  AOI21_X1 u2_u2_u0_U78 (.A( u2_u2_u0_n138 ) , .B2( u2_u2_u0_n139 ) , .B1( u2_u2_u0_n140 ) , .ZN( u2_u2_u0_n157 ) );
  AOI21_X1 u2_u2_u0_U79 (.B2( u2_u2_u0_n141 ) , .B1( u2_u2_u0_n142 ) , .ZN( u2_u2_u0_n156 ) , .A( u2_u2_u0_n161 ) );
  AND2_X1 u2_u2_u0_U8 (.A1( u2_u2_u0_n114 ) , .A2( u2_u2_u0_n121 ) , .ZN( u2_u2_u0_n146 ) );
  AOI21_X1 u2_u2_u0_U80 (.B1( u2_u2_u0_n132 ) , .ZN( u2_u2_u0_n133 ) , .A( u2_u2_u0_n144 ) , .B2( u2_u2_u0_n166 ) );
  OAI22_X1 u2_u2_u0_U81 (.ZN( u2_u2_u0_n105 ) , .A2( u2_u2_u0_n132 ) , .B1( u2_u2_u0_n146 ) , .A1( u2_u2_u0_n147 ) , .B2( u2_u2_u0_n161 ) );
  NAND2_X1 u2_u2_u0_U82 (.ZN( u2_u2_u0_n110 ) , .A2( u2_u2_u0_n132 ) , .A1( u2_u2_u0_n145 ) );
  INV_X1 u2_u2_u0_U83 (.A( u2_u2_u0_n119 ) , .ZN( u2_u2_u0_n167 ) );
  NAND2_X1 u2_u2_u0_U84 (.A2( u2_u2_u0_n103 ) , .ZN( u2_u2_u0_n140 ) , .A1( u2_u2_u0_n94 ) );
  NAND2_X1 u2_u2_u0_U85 (.A1( u2_u2_u0_n101 ) , .ZN( u2_u2_u0_n130 ) , .A2( u2_u2_u0_n94 ) );
  NAND2_X1 u2_u2_u0_U86 (.ZN( u2_u2_u0_n108 ) , .A1( u2_u2_u0_n92 ) , .A2( u2_u2_u0_n94 ) );
  NAND2_X1 u2_u2_u0_U87 (.ZN( u2_u2_u0_n142 ) , .A1( u2_u2_u0_n94 ) , .A2( u2_u2_u0_n95 ) );
  NAND3_X1 u2_u2_u0_U88 (.ZN( u2_out2_23 ) , .A3( u2_u2_u0_n137 ) , .A1( u2_u2_u0_n168 ) , .A2( u2_u2_u0_n171 ) );
  NAND3_X1 u2_u2_u0_U89 (.A3( u2_u2_u0_n127 ) , .A2( u2_u2_u0_n128 ) , .ZN( u2_u2_u0_n135 ) , .A1( u2_u2_u0_n150 ) );
  AND2_X1 u2_u2_u0_U9 (.A1( u2_u2_u0_n131 ) , .ZN( u2_u2_u0_n141 ) , .A2( u2_u2_u0_n150 ) );
  NAND3_X1 u2_u2_u0_U90 (.ZN( u2_u2_u0_n117 ) , .A3( u2_u2_u0_n132 ) , .A2( u2_u2_u0_n139 ) , .A1( u2_u2_u0_n148 ) );
  NAND3_X1 u2_u2_u0_U91 (.ZN( u2_u2_u0_n109 ) , .A2( u2_u2_u0_n114 ) , .A3( u2_u2_u0_n140 ) , .A1( u2_u2_u0_n149 ) );
  NAND3_X1 u2_u2_u0_U92 (.ZN( u2_out2_9 ) , .A3( u2_u2_u0_n106 ) , .A2( u2_u2_u0_n171 ) , .A1( u2_u2_u0_n174 ) );
  NAND3_X1 u2_u2_u0_U93 (.A2( u2_u2_u0_n128 ) , .A1( u2_u2_u0_n132 ) , .A3( u2_u2_u0_n146 ) , .ZN( u2_u2_u0_n97 ) );
  NOR2_X1 u2_u2_u1_U10 (.A1( u2_u2_u1_n112 ) , .A2( u2_u2_u1_n116 ) , .ZN( u2_u2_u1_n118 ) );
  NAND3_X1 u2_u2_u1_U100 (.ZN( u2_u2_u1_n113 ) , .A1( u2_u2_u1_n120 ) , .A3( u2_u2_u1_n133 ) , .A2( u2_u2_u1_n155 ) );
  OAI21_X1 u2_u2_u1_U11 (.ZN( u2_u2_u1_n101 ) , .B1( u2_u2_u1_n141 ) , .A( u2_u2_u1_n146 ) , .B2( u2_u2_u1_n183 ) );
  AOI21_X1 u2_u2_u1_U12 (.B2( u2_u2_u1_n155 ) , .B1( u2_u2_u1_n156 ) , .ZN( u2_u2_u1_n157 ) , .A( u2_u2_u1_n174 ) );
  OR4_X1 u2_u2_u1_U13 (.A4( u2_u2_u1_n106 ) , .A3( u2_u2_u1_n107 ) , .ZN( u2_u2_u1_n108 ) , .A1( u2_u2_u1_n117 ) , .A2( u2_u2_u1_n184 ) );
  AOI21_X1 u2_u2_u1_U14 (.ZN( u2_u2_u1_n106 ) , .A( u2_u2_u1_n112 ) , .B1( u2_u2_u1_n154 ) , .B2( u2_u2_u1_n156 ) );
  INV_X1 u2_u2_u1_U15 (.A( u2_u2_u1_n101 ) , .ZN( u2_u2_u1_n184 ) );
  AOI21_X1 u2_u2_u1_U16 (.ZN( u2_u2_u1_n107 ) , .B1( u2_u2_u1_n134 ) , .B2( u2_u2_u1_n149 ) , .A( u2_u2_u1_n174 ) );
  NAND2_X1 u2_u2_u1_U17 (.ZN( u2_u2_u1_n140 ) , .A2( u2_u2_u1_n150 ) , .A1( u2_u2_u1_n155 ) );
  NAND2_X1 u2_u2_u1_U18 (.A1( u2_u2_u1_n131 ) , .ZN( u2_u2_u1_n147 ) , .A2( u2_u2_u1_n153 ) );
  INV_X1 u2_u2_u1_U19 (.A( u2_u2_u1_n139 ) , .ZN( u2_u2_u1_n174 ) );
  INV_X1 u2_u2_u1_U20 (.A( u2_u2_u1_n112 ) , .ZN( u2_u2_u1_n171 ) );
  NAND2_X1 u2_u2_u1_U21 (.ZN( u2_u2_u1_n141 ) , .A1( u2_u2_u1_n153 ) , .A2( u2_u2_u1_n156 ) );
  AND2_X1 u2_u2_u1_U22 (.A1( u2_u2_u1_n123 ) , .ZN( u2_u2_u1_n134 ) , .A2( u2_u2_u1_n161 ) );
  NAND2_X1 u2_u2_u1_U23 (.A2( u2_u2_u1_n115 ) , .A1( u2_u2_u1_n116 ) , .ZN( u2_u2_u1_n148 ) );
  NAND2_X1 u2_u2_u1_U24 (.A2( u2_u2_u1_n133 ) , .A1( u2_u2_u1_n135 ) , .ZN( u2_u2_u1_n159 ) );
  NAND2_X1 u2_u2_u1_U25 (.A2( u2_u2_u1_n115 ) , .A1( u2_u2_u1_n120 ) , .ZN( u2_u2_u1_n132 ) );
  INV_X1 u2_u2_u1_U26 (.A( u2_u2_u1_n154 ) , .ZN( u2_u2_u1_n178 ) );
  INV_X1 u2_u2_u1_U27 (.A( u2_u2_u1_n151 ) , .ZN( u2_u2_u1_n183 ) );
  AND2_X1 u2_u2_u1_U28 (.A1( u2_u2_u1_n129 ) , .A2( u2_u2_u1_n133 ) , .ZN( u2_u2_u1_n149 ) );
  INV_X1 u2_u2_u1_U29 (.A( u2_u2_u1_n131 ) , .ZN( u2_u2_u1_n180 ) );
  INV_X1 u2_u2_u1_U3 (.A( u2_u2_u1_n159 ) , .ZN( u2_u2_u1_n182 ) );
  OAI221_X1 u2_u2_u1_U30 (.A( u2_u2_u1_n119 ) , .C2( u2_u2_u1_n129 ) , .ZN( u2_u2_u1_n138 ) , .B2( u2_u2_u1_n152 ) , .C1( u2_u2_u1_n174 ) , .B1( u2_u2_u1_n187 ) );
  INV_X1 u2_u2_u1_U31 (.A( u2_u2_u1_n148 ) , .ZN( u2_u2_u1_n187 ) );
  AOI211_X1 u2_u2_u1_U32 (.B( u2_u2_u1_n117 ) , .A( u2_u2_u1_n118 ) , .ZN( u2_u2_u1_n119 ) , .C2( u2_u2_u1_n146 ) , .C1( u2_u2_u1_n159 ) );
  NOR2_X1 u2_u2_u1_U33 (.A1( u2_u2_u1_n168 ) , .A2( u2_u2_u1_n176 ) , .ZN( u2_u2_u1_n98 ) );
  AOI211_X1 u2_u2_u1_U34 (.B( u2_u2_u1_n162 ) , .A( u2_u2_u1_n163 ) , .C2( u2_u2_u1_n164 ) , .ZN( u2_u2_u1_n165 ) , .C1( u2_u2_u1_n171 ) );
  AOI21_X1 u2_u2_u1_U35 (.A( u2_u2_u1_n160 ) , .B2( u2_u2_u1_n161 ) , .ZN( u2_u2_u1_n162 ) , .B1( u2_u2_u1_n182 ) );
  OR2_X1 u2_u2_u1_U36 (.A2( u2_u2_u1_n157 ) , .A1( u2_u2_u1_n158 ) , .ZN( u2_u2_u1_n163 ) );
  OAI21_X1 u2_u2_u1_U37 (.B2( u2_u2_u1_n123 ) , .ZN( u2_u2_u1_n145 ) , .B1( u2_u2_u1_n160 ) , .A( u2_u2_u1_n185 ) );
  INV_X1 u2_u2_u1_U38 (.A( u2_u2_u1_n122 ) , .ZN( u2_u2_u1_n185 ) );
  AOI21_X1 u2_u2_u1_U39 (.B2( u2_u2_u1_n120 ) , .B1( u2_u2_u1_n121 ) , .ZN( u2_u2_u1_n122 ) , .A( u2_u2_u1_n128 ) );
  AOI221_X1 u2_u2_u1_U4 (.A( u2_u2_u1_n138 ) , .C2( u2_u2_u1_n139 ) , .C1( u2_u2_u1_n140 ) , .B2( u2_u2_u1_n141 ) , .ZN( u2_u2_u1_n142 ) , .B1( u2_u2_u1_n175 ) );
  NAND2_X1 u2_u2_u1_U40 (.A1( u2_u2_u1_n128 ) , .ZN( u2_u2_u1_n146 ) , .A2( u2_u2_u1_n160 ) );
  NAND2_X1 u2_u2_u1_U41 (.A2( u2_u2_u1_n112 ) , .ZN( u2_u2_u1_n139 ) , .A1( u2_u2_u1_n152 ) );
  NAND2_X1 u2_u2_u1_U42 (.A1( u2_u2_u1_n105 ) , .ZN( u2_u2_u1_n156 ) , .A2( u2_u2_u1_n99 ) );
  AOI221_X1 u2_u2_u1_U43 (.B1( u2_u2_u1_n140 ) , .ZN( u2_u2_u1_n167 ) , .B2( u2_u2_u1_n172 ) , .C2( u2_u2_u1_n175 ) , .C1( u2_u2_u1_n178 ) , .A( u2_u2_u1_n188 ) );
  INV_X1 u2_u2_u1_U44 (.ZN( u2_u2_u1_n188 ) , .A( u2_u2_u1_n97 ) );
  AOI211_X1 u2_u2_u1_U45 (.A( u2_u2_u1_n118 ) , .C1( u2_u2_u1_n132 ) , .C2( u2_u2_u1_n139 ) , .B( u2_u2_u1_n96 ) , .ZN( u2_u2_u1_n97 ) );
  AOI21_X1 u2_u2_u1_U46 (.B2( u2_u2_u1_n121 ) , .B1( u2_u2_u1_n135 ) , .A( u2_u2_u1_n152 ) , .ZN( u2_u2_u1_n96 ) );
  NOR2_X1 u2_u2_u1_U47 (.ZN( u2_u2_u1_n117 ) , .A1( u2_u2_u1_n121 ) , .A2( u2_u2_u1_n160 ) );
  AOI21_X1 u2_u2_u1_U48 (.A( u2_u2_u1_n128 ) , .B2( u2_u2_u1_n129 ) , .ZN( u2_u2_u1_n130 ) , .B1( u2_u2_u1_n150 ) );
  NAND2_X1 u2_u2_u1_U49 (.ZN( u2_u2_u1_n112 ) , .A1( u2_u2_u1_n169 ) , .A2( u2_u2_u1_n170 ) );
  AOI211_X1 u2_u2_u1_U5 (.ZN( u2_u2_u1_n124 ) , .A( u2_u2_u1_n138 ) , .C2( u2_u2_u1_n139 ) , .B( u2_u2_u1_n145 ) , .C1( u2_u2_u1_n147 ) );
  NAND2_X1 u2_u2_u1_U50 (.ZN( u2_u2_u1_n129 ) , .A2( u2_u2_u1_n95 ) , .A1( u2_u2_u1_n98 ) );
  NAND2_X1 u2_u2_u1_U51 (.A1( u2_u2_u1_n102 ) , .ZN( u2_u2_u1_n154 ) , .A2( u2_u2_u1_n99 ) );
  NAND2_X1 u2_u2_u1_U52 (.A2( u2_u2_u1_n100 ) , .ZN( u2_u2_u1_n135 ) , .A1( u2_u2_u1_n99 ) );
  AOI21_X1 u2_u2_u1_U53 (.A( u2_u2_u1_n152 ) , .B2( u2_u2_u1_n153 ) , .B1( u2_u2_u1_n154 ) , .ZN( u2_u2_u1_n158 ) );
  INV_X1 u2_u2_u1_U54 (.A( u2_u2_u1_n160 ) , .ZN( u2_u2_u1_n175 ) );
  NAND2_X1 u2_u2_u1_U55 (.A1( u2_u2_u1_n100 ) , .ZN( u2_u2_u1_n116 ) , .A2( u2_u2_u1_n95 ) );
  NAND2_X1 u2_u2_u1_U56 (.A1( u2_u2_u1_n102 ) , .ZN( u2_u2_u1_n131 ) , .A2( u2_u2_u1_n95 ) );
  NAND2_X1 u2_u2_u1_U57 (.A2( u2_u2_u1_n104 ) , .ZN( u2_u2_u1_n121 ) , .A1( u2_u2_u1_n98 ) );
  NAND2_X1 u2_u2_u1_U58 (.A1( u2_u2_u1_n103 ) , .ZN( u2_u2_u1_n153 ) , .A2( u2_u2_u1_n98 ) );
  NAND2_X1 u2_u2_u1_U59 (.A2( u2_u2_u1_n104 ) , .A1( u2_u2_u1_n105 ) , .ZN( u2_u2_u1_n133 ) );
  AOI22_X1 u2_u2_u1_U6 (.B2( u2_u2_u1_n113 ) , .A2( u2_u2_u1_n114 ) , .ZN( u2_u2_u1_n125 ) , .A1( u2_u2_u1_n171 ) , .B1( u2_u2_u1_n173 ) );
  NAND2_X1 u2_u2_u1_U60 (.ZN( u2_u2_u1_n150 ) , .A2( u2_u2_u1_n98 ) , .A1( u2_u2_u1_n99 ) );
  NAND2_X1 u2_u2_u1_U61 (.A1( u2_u2_u1_n105 ) , .ZN( u2_u2_u1_n155 ) , .A2( u2_u2_u1_n95 ) );
  OAI21_X1 u2_u2_u1_U62 (.ZN( u2_u2_u1_n109 ) , .B1( u2_u2_u1_n129 ) , .B2( u2_u2_u1_n160 ) , .A( u2_u2_u1_n167 ) );
  NAND2_X1 u2_u2_u1_U63 (.A2( u2_u2_u1_n100 ) , .A1( u2_u2_u1_n103 ) , .ZN( u2_u2_u1_n120 ) );
  NAND2_X1 u2_u2_u1_U64 (.A1( u2_u2_u1_n102 ) , .A2( u2_u2_u1_n104 ) , .ZN( u2_u2_u1_n115 ) );
  NAND2_X1 u2_u2_u1_U65 (.A2( u2_u2_u1_n100 ) , .A1( u2_u2_u1_n104 ) , .ZN( u2_u2_u1_n151 ) );
  NAND2_X1 u2_u2_u1_U66 (.A2( u2_u2_u1_n103 ) , .A1( u2_u2_u1_n105 ) , .ZN( u2_u2_u1_n161 ) );
  INV_X1 u2_u2_u1_U67 (.A( u2_u2_u1_n152 ) , .ZN( u2_u2_u1_n173 ) );
  INV_X1 u2_u2_u1_U68 (.A( u2_u2_u1_n128 ) , .ZN( u2_u2_u1_n172 ) );
  NAND2_X1 u2_u2_u1_U69 (.A2( u2_u2_u1_n102 ) , .A1( u2_u2_u1_n103 ) , .ZN( u2_u2_u1_n123 ) );
  NAND2_X1 u2_u2_u1_U7 (.ZN( u2_u2_u1_n114 ) , .A1( u2_u2_u1_n134 ) , .A2( u2_u2_u1_n156 ) );
  NOR2_X1 u2_u2_u1_U70 (.A2( u2_u2_X_7 ) , .A1( u2_u2_X_8 ) , .ZN( u2_u2_u1_n95 ) );
  NOR2_X1 u2_u2_u1_U71 (.A1( u2_u2_X_12 ) , .A2( u2_u2_X_9 ) , .ZN( u2_u2_u1_n100 ) );
  NOR2_X1 u2_u2_u1_U72 (.A2( u2_u2_X_8 ) , .A1( u2_u2_u1_n177 ) , .ZN( u2_u2_u1_n99 ) );
  NOR2_X1 u2_u2_u1_U73 (.A2( u2_u2_X_12 ) , .ZN( u2_u2_u1_n102 ) , .A1( u2_u2_u1_n176 ) );
  NOR2_X1 u2_u2_u1_U74 (.A2( u2_u2_X_9 ) , .ZN( u2_u2_u1_n105 ) , .A1( u2_u2_u1_n168 ) );
  NAND2_X1 u2_u2_u1_U75 (.A1( u2_u2_X_10 ) , .ZN( u2_u2_u1_n160 ) , .A2( u2_u2_u1_n169 ) );
  NAND2_X1 u2_u2_u1_U76 (.A2( u2_u2_X_10 ) , .A1( u2_u2_X_11 ) , .ZN( u2_u2_u1_n152 ) );
  NAND2_X1 u2_u2_u1_U77 (.A1( u2_u2_X_11 ) , .ZN( u2_u2_u1_n128 ) , .A2( u2_u2_u1_n170 ) );
  AND2_X1 u2_u2_u1_U78 (.A2( u2_u2_X_7 ) , .A1( u2_u2_X_8 ) , .ZN( u2_u2_u1_n104 ) );
  AND2_X1 u2_u2_u1_U79 (.A1( u2_u2_X_8 ) , .ZN( u2_u2_u1_n103 ) , .A2( u2_u2_u1_n177 ) );
  AOI22_X1 u2_u2_u1_U8 (.B2( u2_u2_u1_n136 ) , .A2( u2_u2_u1_n137 ) , .ZN( u2_u2_u1_n143 ) , .A1( u2_u2_u1_n171 ) , .B1( u2_u2_u1_n173 ) );
  INV_X1 u2_u2_u1_U80 (.A( u2_u2_X_10 ) , .ZN( u2_u2_u1_n170 ) );
  INV_X1 u2_u2_u1_U81 (.A( u2_u2_X_9 ) , .ZN( u2_u2_u1_n176 ) );
  INV_X1 u2_u2_u1_U82 (.A( u2_u2_X_11 ) , .ZN( u2_u2_u1_n169 ) );
  INV_X1 u2_u2_u1_U83 (.A( u2_u2_X_12 ) , .ZN( u2_u2_u1_n168 ) );
  INV_X1 u2_u2_u1_U84 (.A( u2_u2_X_7 ) , .ZN( u2_u2_u1_n177 ) );
  NAND4_X1 u2_u2_u1_U85 (.ZN( u2_out2_28 ) , .A4( u2_u2_u1_n124 ) , .A3( u2_u2_u1_n125 ) , .A2( u2_u2_u1_n126 ) , .A1( u2_u2_u1_n127 ) );
  OAI21_X1 u2_u2_u1_U86 (.ZN( u2_u2_u1_n127 ) , .B2( u2_u2_u1_n139 ) , .B1( u2_u2_u1_n175 ) , .A( u2_u2_u1_n183 ) );
  OAI21_X1 u2_u2_u1_U87 (.ZN( u2_u2_u1_n126 ) , .B2( u2_u2_u1_n140 ) , .A( u2_u2_u1_n146 ) , .B1( u2_u2_u1_n178 ) );
  NAND4_X1 u2_u2_u1_U88 (.ZN( u2_out2_18 ) , .A4( u2_u2_u1_n165 ) , .A3( u2_u2_u1_n166 ) , .A1( u2_u2_u1_n167 ) , .A2( u2_u2_u1_n186 ) );
  AOI22_X1 u2_u2_u1_U89 (.B2( u2_u2_u1_n146 ) , .B1( u2_u2_u1_n147 ) , .A2( u2_u2_u1_n148 ) , .ZN( u2_u2_u1_n166 ) , .A1( u2_u2_u1_n172 ) );
  INV_X1 u2_u2_u1_U9 (.A( u2_u2_u1_n147 ) , .ZN( u2_u2_u1_n181 ) );
  INV_X1 u2_u2_u1_U90 (.A( u2_u2_u1_n145 ) , .ZN( u2_u2_u1_n186 ) );
  NAND4_X1 u2_u2_u1_U91 (.ZN( u2_out2_2 ) , .A4( u2_u2_u1_n142 ) , .A3( u2_u2_u1_n143 ) , .A2( u2_u2_u1_n144 ) , .A1( u2_u2_u1_n179 ) );
  OAI21_X1 u2_u2_u1_U92 (.B2( u2_u2_u1_n132 ) , .ZN( u2_u2_u1_n144 ) , .A( u2_u2_u1_n146 ) , .B1( u2_u2_u1_n180 ) );
  INV_X1 u2_u2_u1_U93 (.A( u2_u2_u1_n130 ) , .ZN( u2_u2_u1_n179 ) );
  OR4_X1 u2_u2_u1_U94 (.ZN( u2_out2_13 ) , .A4( u2_u2_u1_n108 ) , .A3( u2_u2_u1_n109 ) , .A2( u2_u2_u1_n110 ) , .A1( u2_u2_u1_n111 ) );
  AOI21_X1 u2_u2_u1_U95 (.ZN( u2_u2_u1_n111 ) , .A( u2_u2_u1_n128 ) , .B2( u2_u2_u1_n131 ) , .B1( u2_u2_u1_n135 ) );
  AOI21_X1 u2_u2_u1_U96 (.ZN( u2_u2_u1_n110 ) , .A( u2_u2_u1_n116 ) , .B1( u2_u2_u1_n152 ) , .B2( u2_u2_u1_n160 ) );
  NAND3_X1 u2_u2_u1_U97 (.A3( u2_u2_u1_n149 ) , .A2( u2_u2_u1_n150 ) , .A1( u2_u2_u1_n151 ) , .ZN( u2_u2_u1_n164 ) );
  NAND3_X1 u2_u2_u1_U98 (.A3( u2_u2_u1_n134 ) , .A2( u2_u2_u1_n135 ) , .ZN( u2_u2_u1_n136 ) , .A1( u2_u2_u1_n151 ) );
  NAND3_X1 u2_u2_u1_U99 (.A1( u2_u2_u1_n133 ) , .ZN( u2_u2_u1_n137 ) , .A2( u2_u2_u1_n154 ) , .A3( u2_u2_u1_n181 ) );
  OAI22_X1 u2_u2_u2_U10 (.B1( u2_u2_u2_n151 ) , .A2( u2_u2_u2_n152 ) , .A1( u2_u2_u2_n153 ) , .ZN( u2_u2_u2_n160 ) , .B2( u2_u2_u2_n168 ) );
  NAND3_X1 u2_u2_u2_U100 (.A2( u2_u2_u2_n100 ) , .A1( u2_u2_u2_n104 ) , .A3( u2_u2_u2_n138 ) , .ZN( u2_u2_u2_n98 ) );
  NOR3_X1 u2_u2_u2_U11 (.A1( u2_u2_u2_n150 ) , .ZN( u2_u2_u2_n151 ) , .A3( u2_u2_u2_n175 ) , .A2( u2_u2_u2_n188 ) );
  AOI21_X1 u2_u2_u2_U12 (.B2( u2_u2_u2_n123 ) , .ZN( u2_u2_u2_n125 ) , .A( u2_u2_u2_n171 ) , .B1( u2_u2_u2_n184 ) );
  INV_X1 u2_u2_u2_U13 (.A( u2_u2_u2_n150 ) , .ZN( u2_u2_u2_n184 ) );
  AOI21_X1 u2_u2_u2_U14 (.ZN( u2_u2_u2_n144 ) , .B2( u2_u2_u2_n155 ) , .A( u2_u2_u2_n172 ) , .B1( u2_u2_u2_n185 ) );
  AOI21_X1 u2_u2_u2_U15 (.B2( u2_u2_u2_n143 ) , .ZN( u2_u2_u2_n145 ) , .B1( u2_u2_u2_n152 ) , .A( u2_u2_u2_n171 ) );
  INV_X1 u2_u2_u2_U16 (.A( u2_u2_u2_n156 ) , .ZN( u2_u2_u2_n171 ) );
  INV_X1 u2_u2_u2_U17 (.A( u2_u2_u2_n120 ) , .ZN( u2_u2_u2_n188 ) );
  NAND2_X1 u2_u2_u2_U18 (.A2( u2_u2_u2_n122 ) , .ZN( u2_u2_u2_n150 ) , .A1( u2_u2_u2_n152 ) );
  INV_X1 u2_u2_u2_U19 (.A( u2_u2_u2_n153 ) , .ZN( u2_u2_u2_n170 ) );
  INV_X1 u2_u2_u2_U20 (.A( u2_u2_u2_n137 ) , .ZN( u2_u2_u2_n173 ) );
  NAND2_X1 u2_u2_u2_U21 (.A1( u2_u2_u2_n132 ) , .A2( u2_u2_u2_n139 ) , .ZN( u2_u2_u2_n157 ) );
  INV_X1 u2_u2_u2_U22 (.A( u2_u2_u2_n113 ) , .ZN( u2_u2_u2_n178 ) );
  INV_X1 u2_u2_u2_U23 (.A( u2_u2_u2_n139 ) , .ZN( u2_u2_u2_n175 ) );
  INV_X1 u2_u2_u2_U24 (.A( u2_u2_u2_n155 ) , .ZN( u2_u2_u2_n181 ) );
  INV_X1 u2_u2_u2_U25 (.A( u2_u2_u2_n119 ) , .ZN( u2_u2_u2_n177 ) );
  INV_X1 u2_u2_u2_U26 (.A( u2_u2_u2_n116 ) , .ZN( u2_u2_u2_n180 ) );
  INV_X1 u2_u2_u2_U27 (.A( u2_u2_u2_n131 ) , .ZN( u2_u2_u2_n179 ) );
  INV_X1 u2_u2_u2_U28 (.A( u2_u2_u2_n154 ) , .ZN( u2_u2_u2_n176 ) );
  NAND2_X1 u2_u2_u2_U29 (.A2( u2_u2_u2_n116 ) , .A1( u2_u2_u2_n117 ) , .ZN( u2_u2_u2_n118 ) );
  NOR2_X1 u2_u2_u2_U3 (.ZN( u2_u2_u2_n121 ) , .A2( u2_u2_u2_n177 ) , .A1( u2_u2_u2_n180 ) );
  INV_X1 u2_u2_u2_U30 (.A( u2_u2_u2_n132 ) , .ZN( u2_u2_u2_n182 ) );
  INV_X1 u2_u2_u2_U31 (.A( u2_u2_u2_n158 ) , .ZN( u2_u2_u2_n183 ) );
  OAI21_X1 u2_u2_u2_U32 (.A( u2_u2_u2_n156 ) , .B1( u2_u2_u2_n157 ) , .ZN( u2_u2_u2_n158 ) , .B2( u2_u2_u2_n179 ) );
  NOR2_X1 u2_u2_u2_U33 (.ZN( u2_u2_u2_n156 ) , .A1( u2_u2_u2_n166 ) , .A2( u2_u2_u2_n169 ) );
  NOR2_X1 u2_u2_u2_U34 (.A2( u2_u2_u2_n114 ) , .ZN( u2_u2_u2_n137 ) , .A1( u2_u2_u2_n140 ) );
  NOR2_X1 u2_u2_u2_U35 (.A2( u2_u2_u2_n138 ) , .ZN( u2_u2_u2_n153 ) , .A1( u2_u2_u2_n156 ) );
  AOI211_X1 u2_u2_u2_U36 (.ZN( u2_u2_u2_n130 ) , .C1( u2_u2_u2_n138 ) , .C2( u2_u2_u2_n179 ) , .B( u2_u2_u2_n96 ) , .A( u2_u2_u2_n97 ) );
  OAI22_X1 u2_u2_u2_U37 (.B1( u2_u2_u2_n133 ) , .A2( u2_u2_u2_n137 ) , .A1( u2_u2_u2_n152 ) , .B2( u2_u2_u2_n168 ) , .ZN( u2_u2_u2_n97 ) );
  OAI221_X1 u2_u2_u2_U38 (.B1( u2_u2_u2_n113 ) , .C1( u2_u2_u2_n132 ) , .A( u2_u2_u2_n149 ) , .B2( u2_u2_u2_n171 ) , .C2( u2_u2_u2_n172 ) , .ZN( u2_u2_u2_n96 ) );
  OAI221_X1 u2_u2_u2_U39 (.A( u2_u2_u2_n115 ) , .C2( u2_u2_u2_n123 ) , .B2( u2_u2_u2_n143 ) , .B1( u2_u2_u2_n153 ) , .ZN( u2_u2_u2_n163 ) , .C1( u2_u2_u2_n168 ) );
  INV_X1 u2_u2_u2_U4 (.A( u2_u2_u2_n134 ) , .ZN( u2_u2_u2_n185 ) );
  OAI21_X1 u2_u2_u2_U40 (.A( u2_u2_u2_n114 ) , .ZN( u2_u2_u2_n115 ) , .B1( u2_u2_u2_n176 ) , .B2( u2_u2_u2_n178 ) );
  OAI221_X1 u2_u2_u2_U41 (.A( u2_u2_u2_n135 ) , .B2( u2_u2_u2_n136 ) , .B1( u2_u2_u2_n137 ) , .ZN( u2_u2_u2_n162 ) , .C2( u2_u2_u2_n167 ) , .C1( u2_u2_u2_n185 ) );
  AND3_X1 u2_u2_u2_U42 (.A3( u2_u2_u2_n131 ) , .A2( u2_u2_u2_n132 ) , .A1( u2_u2_u2_n133 ) , .ZN( u2_u2_u2_n136 ) );
  AOI22_X1 u2_u2_u2_U43 (.ZN( u2_u2_u2_n135 ) , .B1( u2_u2_u2_n140 ) , .A1( u2_u2_u2_n156 ) , .B2( u2_u2_u2_n180 ) , .A2( u2_u2_u2_n188 ) );
  AOI21_X1 u2_u2_u2_U44 (.ZN( u2_u2_u2_n149 ) , .B1( u2_u2_u2_n173 ) , .B2( u2_u2_u2_n188 ) , .A( u2_u2_u2_n95 ) );
  AND3_X1 u2_u2_u2_U45 (.A2( u2_u2_u2_n100 ) , .A1( u2_u2_u2_n104 ) , .A3( u2_u2_u2_n156 ) , .ZN( u2_u2_u2_n95 ) );
  OAI21_X1 u2_u2_u2_U46 (.A( u2_u2_u2_n141 ) , .B2( u2_u2_u2_n142 ) , .ZN( u2_u2_u2_n146 ) , .B1( u2_u2_u2_n153 ) );
  OAI21_X1 u2_u2_u2_U47 (.A( u2_u2_u2_n140 ) , .ZN( u2_u2_u2_n141 ) , .B1( u2_u2_u2_n176 ) , .B2( u2_u2_u2_n177 ) );
  NOR3_X1 u2_u2_u2_U48 (.ZN( u2_u2_u2_n142 ) , .A3( u2_u2_u2_n175 ) , .A2( u2_u2_u2_n178 ) , .A1( u2_u2_u2_n181 ) );
  OAI21_X1 u2_u2_u2_U49 (.A( u2_u2_u2_n101 ) , .B2( u2_u2_u2_n121 ) , .B1( u2_u2_u2_n153 ) , .ZN( u2_u2_u2_n164 ) );
  NOR4_X1 u2_u2_u2_U5 (.A4( u2_u2_u2_n124 ) , .A3( u2_u2_u2_n125 ) , .A2( u2_u2_u2_n126 ) , .A1( u2_u2_u2_n127 ) , .ZN( u2_u2_u2_n128 ) );
  NAND2_X1 u2_u2_u2_U50 (.A2( u2_u2_u2_n100 ) , .A1( u2_u2_u2_n107 ) , .ZN( u2_u2_u2_n155 ) );
  NAND2_X1 u2_u2_u2_U51 (.A2( u2_u2_u2_n105 ) , .A1( u2_u2_u2_n108 ) , .ZN( u2_u2_u2_n143 ) );
  NAND2_X1 u2_u2_u2_U52 (.A1( u2_u2_u2_n104 ) , .A2( u2_u2_u2_n106 ) , .ZN( u2_u2_u2_n152 ) );
  NAND2_X1 u2_u2_u2_U53 (.A1( u2_u2_u2_n100 ) , .A2( u2_u2_u2_n105 ) , .ZN( u2_u2_u2_n132 ) );
  INV_X1 u2_u2_u2_U54 (.A( u2_u2_u2_n140 ) , .ZN( u2_u2_u2_n168 ) );
  INV_X1 u2_u2_u2_U55 (.A( u2_u2_u2_n138 ) , .ZN( u2_u2_u2_n167 ) );
  INV_X1 u2_u2_u2_U56 (.ZN( u2_u2_u2_n187 ) , .A( u2_u2_u2_n99 ) );
  OAI21_X1 u2_u2_u2_U57 (.B1( u2_u2_u2_n137 ) , .B2( u2_u2_u2_n143 ) , .A( u2_u2_u2_n98 ) , .ZN( u2_u2_u2_n99 ) );
  NAND2_X1 u2_u2_u2_U58 (.A1( u2_u2_u2_n102 ) , .A2( u2_u2_u2_n106 ) , .ZN( u2_u2_u2_n113 ) );
  NAND2_X1 u2_u2_u2_U59 (.A1( u2_u2_u2_n106 ) , .A2( u2_u2_u2_n107 ) , .ZN( u2_u2_u2_n131 ) );
  AOI21_X1 u2_u2_u2_U6 (.B2( u2_u2_u2_n119 ) , .ZN( u2_u2_u2_n127 ) , .A( u2_u2_u2_n137 ) , .B1( u2_u2_u2_n155 ) );
  NAND2_X1 u2_u2_u2_U60 (.A1( u2_u2_u2_n103 ) , .A2( u2_u2_u2_n107 ) , .ZN( u2_u2_u2_n139 ) );
  NAND2_X1 u2_u2_u2_U61 (.A1( u2_u2_u2_n103 ) , .A2( u2_u2_u2_n105 ) , .ZN( u2_u2_u2_n133 ) );
  NAND2_X1 u2_u2_u2_U62 (.A1( u2_u2_u2_n102 ) , .A2( u2_u2_u2_n103 ) , .ZN( u2_u2_u2_n154 ) );
  NAND2_X1 u2_u2_u2_U63 (.A2( u2_u2_u2_n103 ) , .A1( u2_u2_u2_n104 ) , .ZN( u2_u2_u2_n119 ) );
  NAND2_X1 u2_u2_u2_U64 (.A2( u2_u2_u2_n107 ) , .A1( u2_u2_u2_n108 ) , .ZN( u2_u2_u2_n123 ) );
  NAND2_X1 u2_u2_u2_U65 (.A1( u2_u2_u2_n104 ) , .A2( u2_u2_u2_n108 ) , .ZN( u2_u2_u2_n122 ) );
  INV_X1 u2_u2_u2_U66 (.A( u2_u2_u2_n114 ) , .ZN( u2_u2_u2_n172 ) );
  NAND2_X1 u2_u2_u2_U67 (.A2( u2_u2_u2_n100 ) , .A1( u2_u2_u2_n102 ) , .ZN( u2_u2_u2_n116 ) );
  NAND2_X1 u2_u2_u2_U68 (.A1( u2_u2_u2_n102 ) , .A2( u2_u2_u2_n108 ) , .ZN( u2_u2_u2_n120 ) );
  NAND2_X1 u2_u2_u2_U69 (.A2( u2_u2_u2_n105 ) , .A1( u2_u2_u2_n106 ) , .ZN( u2_u2_u2_n117 ) );
  AOI21_X1 u2_u2_u2_U7 (.ZN( u2_u2_u2_n124 ) , .B1( u2_u2_u2_n131 ) , .B2( u2_u2_u2_n143 ) , .A( u2_u2_u2_n172 ) );
  NOR2_X1 u2_u2_u2_U70 (.A2( u2_u2_X_16 ) , .ZN( u2_u2_u2_n140 ) , .A1( u2_u2_u2_n166 ) );
  NOR2_X1 u2_u2_u2_U71 (.A2( u2_u2_X_13 ) , .A1( u2_u2_X_14 ) , .ZN( u2_u2_u2_n100 ) );
  NOR2_X1 u2_u2_u2_U72 (.A2( u2_u2_X_16 ) , .A1( u2_u2_X_17 ) , .ZN( u2_u2_u2_n138 ) );
  NOR2_X1 u2_u2_u2_U73 (.A2( u2_u2_X_15 ) , .A1( u2_u2_X_18 ) , .ZN( u2_u2_u2_n104 ) );
  NOR2_X1 u2_u2_u2_U74 (.A2( u2_u2_X_14 ) , .ZN( u2_u2_u2_n103 ) , .A1( u2_u2_u2_n174 ) );
  NOR2_X1 u2_u2_u2_U75 (.A2( u2_u2_X_15 ) , .ZN( u2_u2_u2_n102 ) , .A1( u2_u2_u2_n165 ) );
  NOR2_X1 u2_u2_u2_U76 (.A2( u2_u2_X_17 ) , .ZN( u2_u2_u2_n114 ) , .A1( u2_u2_u2_n169 ) );
  AND2_X1 u2_u2_u2_U77 (.A1( u2_u2_X_15 ) , .ZN( u2_u2_u2_n105 ) , .A2( u2_u2_u2_n165 ) );
  AND2_X1 u2_u2_u2_U78 (.A2( u2_u2_X_15 ) , .A1( u2_u2_X_18 ) , .ZN( u2_u2_u2_n107 ) );
  AND2_X1 u2_u2_u2_U79 (.A1( u2_u2_X_14 ) , .ZN( u2_u2_u2_n106 ) , .A2( u2_u2_u2_n174 ) );
  AOI21_X1 u2_u2_u2_U8 (.B2( u2_u2_u2_n120 ) , .B1( u2_u2_u2_n121 ) , .ZN( u2_u2_u2_n126 ) , .A( u2_u2_u2_n167 ) );
  AND2_X1 u2_u2_u2_U80 (.A1( u2_u2_X_13 ) , .A2( u2_u2_X_14 ) , .ZN( u2_u2_u2_n108 ) );
  INV_X1 u2_u2_u2_U81 (.A( u2_u2_X_16 ) , .ZN( u2_u2_u2_n169 ) );
  INV_X1 u2_u2_u2_U82 (.A( u2_u2_X_17 ) , .ZN( u2_u2_u2_n166 ) );
  INV_X1 u2_u2_u2_U83 (.A( u2_u2_X_13 ) , .ZN( u2_u2_u2_n174 ) );
  INV_X1 u2_u2_u2_U84 (.A( u2_u2_X_18 ) , .ZN( u2_u2_u2_n165 ) );
  NAND4_X1 u2_u2_u2_U85 (.ZN( u2_out2_24 ) , .A4( u2_u2_u2_n111 ) , .A3( u2_u2_u2_n112 ) , .A1( u2_u2_u2_n130 ) , .A2( u2_u2_u2_n187 ) );
  AOI21_X1 u2_u2_u2_U86 (.ZN( u2_u2_u2_n112 ) , .B2( u2_u2_u2_n156 ) , .A( u2_u2_u2_n164 ) , .B1( u2_u2_u2_n181 ) );
  AOI221_X1 u2_u2_u2_U87 (.A( u2_u2_u2_n109 ) , .B1( u2_u2_u2_n110 ) , .ZN( u2_u2_u2_n111 ) , .C1( u2_u2_u2_n134 ) , .C2( u2_u2_u2_n170 ) , .B2( u2_u2_u2_n173 ) );
  NAND4_X1 u2_u2_u2_U88 (.ZN( u2_out2_16 ) , .A4( u2_u2_u2_n128 ) , .A3( u2_u2_u2_n129 ) , .A1( u2_u2_u2_n130 ) , .A2( u2_u2_u2_n186 ) );
  AOI22_X1 u2_u2_u2_U89 (.A2( u2_u2_u2_n118 ) , .ZN( u2_u2_u2_n129 ) , .A1( u2_u2_u2_n140 ) , .B1( u2_u2_u2_n157 ) , .B2( u2_u2_u2_n170 ) );
  OAI22_X1 u2_u2_u2_U9 (.ZN( u2_u2_u2_n109 ) , .A2( u2_u2_u2_n113 ) , .B2( u2_u2_u2_n133 ) , .B1( u2_u2_u2_n167 ) , .A1( u2_u2_u2_n168 ) );
  INV_X1 u2_u2_u2_U90 (.A( u2_u2_u2_n163 ) , .ZN( u2_u2_u2_n186 ) );
  NAND4_X1 u2_u2_u2_U91 (.ZN( u2_out2_30 ) , .A4( u2_u2_u2_n147 ) , .A3( u2_u2_u2_n148 ) , .A2( u2_u2_u2_n149 ) , .A1( u2_u2_u2_n187 ) );
  NOR3_X1 u2_u2_u2_U92 (.A3( u2_u2_u2_n144 ) , .A2( u2_u2_u2_n145 ) , .A1( u2_u2_u2_n146 ) , .ZN( u2_u2_u2_n147 ) );
  AOI21_X1 u2_u2_u2_U93 (.B2( u2_u2_u2_n138 ) , .ZN( u2_u2_u2_n148 ) , .A( u2_u2_u2_n162 ) , .B1( u2_u2_u2_n182 ) );
  OR4_X1 u2_u2_u2_U94 (.ZN( u2_out2_6 ) , .A4( u2_u2_u2_n161 ) , .A3( u2_u2_u2_n162 ) , .A2( u2_u2_u2_n163 ) , .A1( u2_u2_u2_n164 ) );
  OR3_X1 u2_u2_u2_U95 (.A2( u2_u2_u2_n159 ) , .A1( u2_u2_u2_n160 ) , .ZN( u2_u2_u2_n161 ) , .A3( u2_u2_u2_n183 ) );
  AOI21_X1 u2_u2_u2_U96 (.B2( u2_u2_u2_n154 ) , .B1( u2_u2_u2_n155 ) , .ZN( u2_u2_u2_n159 ) , .A( u2_u2_u2_n167 ) );
  NAND3_X1 u2_u2_u2_U97 (.A2( u2_u2_u2_n117 ) , .A1( u2_u2_u2_n122 ) , .A3( u2_u2_u2_n123 ) , .ZN( u2_u2_u2_n134 ) );
  NAND3_X1 u2_u2_u2_U98 (.ZN( u2_u2_u2_n110 ) , .A2( u2_u2_u2_n131 ) , .A3( u2_u2_u2_n139 ) , .A1( u2_u2_u2_n154 ) );
  NAND3_X1 u2_u2_u2_U99 (.A2( u2_u2_u2_n100 ) , .ZN( u2_u2_u2_n101 ) , .A1( u2_u2_u2_n104 ) , .A3( u2_u2_u2_n114 ) );
  OAI22_X1 u2_u2_u3_U10 (.B1( u2_u2_u3_n113 ) , .A2( u2_u2_u3_n135 ) , .A1( u2_u2_u3_n150 ) , .B2( u2_u2_u3_n164 ) , .ZN( u2_u2_u3_n98 ) );
  OAI211_X1 u2_u2_u3_U11 (.B( u2_u2_u3_n106 ) , .ZN( u2_u2_u3_n119 ) , .C2( u2_u2_u3_n128 ) , .C1( u2_u2_u3_n167 ) , .A( u2_u2_u3_n181 ) );
  AOI221_X1 u2_u2_u3_U12 (.C1( u2_u2_u3_n105 ) , .ZN( u2_u2_u3_n106 ) , .A( u2_u2_u3_n131 ) , .B2( u2_u2_u3_n132 ) , .C2( u2_u2_u3_n133 ) , .B1( u2_u2_u3_n169 ) );
  INV_X1 u2_u2_u3_U13 (.ZN( u2_u2_u3_n181 ) , .A( u2_u2_u3_n98 ) );
  NAND2_X1 u2_u2_u3_U14 (.ZN( u2_u2_u3_n105 ) , .A2( u2_u2_u3_n130 ) , .A1( u2_u2_u3_n155 ) );
  AOI22_X1 u2_u2_u3_U15 (.B1( u2_u2_u3_n115 ) , .A2( u2_u2_u3_n116 ) , .ZN( u2_u2_u3_n123 ) , .B2( u2_u2_u3_n133 ) , .A1( u2_u2_u3_n169 ) );
  NAND2_X1 u2_u2_u3_U16 (.ZN( u2_u2_u3_n116 ) , .A2( u2_u2_u3_n151 ) , .A1( u2_u2_u3_n182 ) );
  NOR2_X1 u2_u2_u3_U17 (.ZN( u2_u2_u3_n126 ) , .A2( u2_u2_u3_n150 ) , .A1( u2_u2_u3_n164 ) );
  AOI21_X1 u2_u2_u3_U18 (.ZN( u2_u2_u3_n112 ) , .B2( u2_u2_u3_n146 ) , .B1( u2_u2_u3_n155 ) , .A( u2_u2_u3_n167 ) );
  NAND2_X1 u2_u2_u3_U19 (.A1( u2_u2_u3_n135 ) , .ZN( u2_u2_u3_n142 ) , .A2( u2_u2_u3_n164 ) );
  NAND2_X1 u2_u2_u3_U20 (.ZN( u2_u2_u3_n132 ) , .A2( u2_u2_u3_n152 ) , .A1( u2_u2_u3_n156 ) );
  AND2_X1 u2_u2_u3_U21 (.A2( u2_u2_u3_n113 ) , .A1( u2_u2_u3_n114 ) , .ZN( u2_u2_u3_n151 ) );
  INV_X1 u2_u2_u3_U22 (.A( u2_u2_u3_n133 ) , .ZN( u2_u2_u3_n165 ) );
  INV_X1 u2_u2_u3_U23 (.A( u2_u2_u3_n135 ) , .ZN( u2_u2_u3_n170 ) );
  NAND2_X1 u2_u2_u3_U24 (.A1( u2_u2_u3_n107 ) , .A2( u2_u2_u3_n108 ) , .ZN( u2_u2_u3_n140 ) );
  NAND2_X1 u2_u2_u3_U25 (.ZN( u2_u2_u3_n117 ) , .A1( u2_u2_u3_n124 ) , .A2( u2_u2_u3_n148 ) );
  NAND2_X1 u2_u2_u3_U26 (.ZN( u2_u2_u3_n143 ) , .A1( u2_u2_u3_n165 ) , .A2( u2_u2_u3_n167 ) );
  INV_X1 u2_u2_u3_U27 (.A( u2_u2_u3_n130 ) , .ZN( u2_u2_u3_n177 ) );
  INV_X1 u2_u2_u3_U28 (.A( u2_u2_u3_n128 ) , .ZN( u2_u2_u3_n176 ) );
  INV_X1 u2_u2_u3_U29 (.A( u2_u2_u3_n155 ) , .ZN( u2_u2_u3_n174 ) );
  INV_X1 u2_u2_u3_U3 (.A( u2_u2_u3_n129 ) , .ZN( u2_u2_u3_n183 ) );
  INV_X1 u2_u2_u3_U30 (.A( u2_u2_u3_n139 ) , .ZN( u2_u2_u3_n185 ) );
  NOR2_X1 u2_u2_u3_U31 (.ZN( u2_u2_u3_n135 ) , .A2( u2_u2_u3_n141 ) , .A1( u2_u2_u3_n169 ) );
  OAI222_X1 u2_u2_u3_U32 (.C2( u2_u2_u3_n107 ) , .A2( u2_u2_u3_n108 ) , .B1( u2_u2_u3_n135 ) , .ZN( u2_u2_u3_n138 ) , .B2( u2_u2_u3_n146 ) , .C1( u2_u2_u3_n154 ) , .A1( u2_u2_u3_n164 ) );
  NOR4_X1 u2_u2_u3_U33 (.A4( u2_u2_u3_n157 ) , .A3( u2_u2_u3_n158 ) , .A2( u2_u2_u3_n159 ) , .A1( u2_u2_u3_n160 ) , .ZN( u2_u2_u3_n161 ) );
  AOI21_X1 u2_u2_u3_U34 (.B2( u2_u2_u3_n152 ) , .B1( u2_u2_u3_n153 ) , .ZN( u2_u2_u3_n158 ) , .A( u2_u2_u3_n164 ) );
  AOI21_X1 u2_u2_u3_U35 (.A( u2_u2_u3_n154 ) , .B2( u2_u2_u3_n155 ) , .B1( u2_u2_u3_n156 ) , .ZN( u2_u2_u3_n157 ) );
  AOI21_X1 u2_u2_u3_U36 (.A( u2_u2_u3_n149 ) , .B2( u2_u2_u3_n150 ) , .B1( u2_u2_u3_n151 ) , .ZN( u2_u2_u3_n159 ) );
  AOI211_X1 u2_u2_u3_U37 (.ZN( u2_u2_u3_n109 ) , .A( u2_u2_u3_n119 ) , .C2( u2_u2_u3_n129 ) , .B( u2_u2_u3_n138 ) , .C1( u2_u2_u3_n141 ) );
  AOI211_X1 u2_u2_u3_U38 (.B( u2_u2_u3_n119 ) , .A( u2_u2_u3_n120 ) , .C2( u2_u2_u3_n121 ) , .ZN( u2_u2_u3_n122 ) , .C1( u2_u2_u3_n179 ) );
  INV_X1 u2_u2_u3_U39 (.A( u2_u2_u3_n156 ) , .ZN( u2_u2_u3_n179 ) );
  INV_X1 u2_u2_u3_U4 (.A( u2_u2_u3_n140 ) , .ZN( u2_u2_u3_n182 ) );
  OAI22_X1 u2_u2_u3_U40 (.B1( u2_u2_u3_n118 ) , .ZN( u2_u2_u3_n120 ) , .A1( u2_u2_u3_n135 ) , .B2( u2_u2_u3_n154 ) , .A2( u2_u2_u3_n178 ) );
  AND3_X1 u2_u2_u3_U41 (.ZN( u2_u2_u3_n118 ) , .A2( u2_u2_u3_n124 ) , .A1( u2_u2_u3_n144 ) , .A3( u2_u2_u3_n152 ) );
  INV_X1 u2_u2_u3_U42 (.A( u2_u2_u3_n121 ) , .ZN( u2_u2_u3_n164 ) );
  NAND2_X1 u2_u2_u3_U43 (.ZN( u2_u2_u3_n133 ) , .A1( u2_u2_u3_n154 ) , .A2( u2_u2_u3_n164 ) );
  OAI211_X1 u2_u2_u3_U44 (.B( u2_u2_u3_n127 ) , .ZN( u2_u2_u3_n139 ) , .C1( u2_u2_u3_n150 ) , .C2( u2_u2_u3_n154 ) , .A( u2_u2_u3_n184 ) );
  INV_X1 u2_u2_u3_U45 (.A( u2_u2_u3_n125 ) , .ZN( u2_u2_u3_n184 ) );
  AOI221_X1 u2_u2_u3_U46 (.A( u2_u2_u3_n126 ) , .ZN( u2_u2_u3_n127 ) , .C2( u2_u2_u3_n132 ) , .C1( u2_u2_u3_n169 ) , .B2( u2_u2_u3_n170 ) , .B1( u2_u2_u3_n174 ) );
  OAI22_X1 u2_u2_u3_U47 (.A1( u2_u2_u3_n124 ) , .ZN( u2_u2_u3_n125 ) , .B2( u2_u2_u3_n145 ) , .A2( u2_u2_u3_n165 ) , .B1( u2_u2_u3_n167 ) );
  NOR2_X1 u2_u2_u3_U48 (.A1( u2_u2_u3_n113 ) , .ZN( u2_u2_u3_n131 ) , .A2( u2_u2_u3_n154 ) );
  NAND2_X1 u2_u2_u3_U49 (.A1( u2_u2_u3_n103 ) , .ZN( u2_u2_u3_n150 ) , .A2( u2_u2_u3_n99 ) );
  INV_X1 u2_u2_u3_U5 (.A( u2_u2_u3_n117 ) , .ZN( u2_u2_u3_n178 ) );
  NAND2_X1 u2_u2_u3_U50 (.A2( u2_u2_u3_n102 ) , .ZN( u2_u2_u3_n155 ) , .A1( u2_u2_u3_n97 ) );
  INV_X1 u2_u2_u3_U51 (.A( u2_u2_u3_n141 ) , .ZN( u2_u2_u3_n167 ) );
  AOI21_X1 u2_u2_u3_U52 (.B2( u2_u2_u3_n114 ) , .B1( u2_u2_u3_n146 ) , .A( u2_u2_u3_n154 ) , .ZN( u2_u2_u3_n94 ) );
  AOI21_X1 u2_u2_u3_U53 (.ZN( u2_u2_u3_n110 ) , .B2( u2_u2_u3_n142 ) , .B1( u2_u2_u3_n186 ) , .A( u2_u2_u3_n95 ) );
  INV_X1 u2_u2_u3_U54 (.A( u2_u2_u3_n145 ) , .ZN( u2_u2_u3_n186 ) );
  AOI21_X1 u2_u2_u3_U55 (.B1( u2_u2_u3_n124 ) , .A( u2_u2_u3_n149 ) , .B2( u2_u2_u3_n155 ) , .ZN( u2_u2_u3_n95 ) );
  INV_X1 u2_u2_u3_U56 (.A( u2_u2_u3_n149 ) , .ZN( u2_u2_u3_n169 ) );
  NAND2_X1 u2_u2_u3_U57 (.ZN( u2_u2_u3_n124 ) , .A1( u2_u2_u3_n96 ) , .A2( u2_u2_u3_n97 ) );
  NAND2_X1 u2_u2_u3_U58 (.A2( u2_u2_u3_n100 ) , .ZN( u2_u2_u3_n146 ) , .A1( u2_u2_u3_n96 ) );
  NAND2_X1 u2_u2_u3_U59 (.A1( u2_u2_u3_n101 ) , .ZN( u2_u2_u3_n145 ) , .A2( u2_u2_u3_n99 ) );
  AOI221_X1 u2_u2_u3_U6 (.A( u2_u2_u3_n131 ) , .C2( u2_u2_u3_n132 ) , .C1( u2_u2_u3_n133 ) , .ZN( u2_u2_u3_n134 ) , .B1( u2_u2_u3_n143 ) , .B2( u2_u2_u3_n177 ) );
  NAND2_X1 u2_u2_u3_U60 (.A1( u2_u2_u3_n100 ) , .ZN( u2_u2_u3_n156 ) , .A2( u2_u2_u3_n99 ) );
  NAND2_X1 u2_u2_u3_U61 (.A2( u2_u2_u3_n101 ) , .A1( u2_u2_u3_n104 ) , .ZN( u2_u2_u3_n148 ) );
  NAND2_X1 u2_u2_u3_U62 (.A1( u2_u2_u3_n100 ) , .A2( u2_u2_u3_n102 ) , .ZN( u2_u2_u3_n128 ) );
  NAND2_X1 u2_u2_u3_U63 (.A2( u2_u2_u3_n101 ) , .A1( u2_u2_u3_n102 ) , .ZN( u2_u2_u3_n152 ) );
  NAND2_X1 u2_u2_u3_U64 (.A2( u2_u2_u3_n101 ) , .ZN( u2_u2_u3_n114 ) , .A1( u2_u2_u3_n96 ) );
  NAND2_X1 u2_u2_u3_U65 (.ZN( u2_u2_u3_n107 ) , .A1( u2_u2_u3_n97 ) , .A2( u2_u2_u3_n99 ) );
  NAND2_X1 u2_u2_u3_U66 (.A2( u2_u2_u3_n100 ) , .A1( u2_u2_u3_n104 ) , .ZN( u2_u2_u3_n113 ) );
  NAND2_X1 u2_u2_u3_U67 (.A1( u2_u2_u3_n104 ) , .ZN( u2_u2_u3_n153 ) , .A2( u2_u2_u3_n97 ) );
  NAND2_X1 u2_u2_u3_U68 (.A2( u2_u2_u3_n103 ) , .A1( u2_u2_u3_n104 ) , .ZN( u2_u2_u3_n130 ) );
  NAND2_X1 u2_u2_u3_U69 (.A2( u2_u2_u3_n103 ) , .ZN( u2_u2_u3_n144 ) , .A1( u2_u2_u3_n96 ) );
  OAI22_X1 u2_u2_u3_U7 (.B2( u2_u2_u3_n147 ) , .A2( u2_u2_u3_n148 ) , .ZN( u2_u2_u3_n160 ) , .B1( u2_u2_u3_n165 ) , .A1( u2_u2_u3_n168 ) );
  NAND2_X1 u2_u2_u3_U70 (.A1( u2_u2_u3_n102 ) , .A2( u2_u2_u3_n103 ) , .ZN( u2_u2_u3_n108 ) );
  NOR2_X1 u2_u2_u3_U71 (.A2( u2_u2_X_19 ) , .A1( u2_u2_X_20 ) , .ZN( u2_u2_u3_n99 ) );
  NOR2_X1 u2_u2_u3_U72 (.A2( u2_u2_X_21 ) , .A1( u2_u2_X_24 ) , .ZN( u2_u2_u3_n103 ) );
  NOR2_X1 u2_u2_u3_U73 (.A2( u2_u2_X_24 ) , .A1( u2_u2_u3_n171 ) , .ZN( u2_u2_u3_n97 ) );
  NOR2_X1 u2_u2_u3_U74 (.A2( u2_u2_X_23 ) , .ZN( u2_u2_u3_n141 ) , .A1( u2_u2_u3_n166 ) );
  NOR2_X1 u2_u2_u3_U75 (.A2( u2_u2_X_19 ) , .A1( u2_u2_u3_n172 ) , .ZN( u2_u2_u3_n96 ) );
  NAND2_X1 u2_u2_u3_U76 (.A1( u2_u2_X_22 ) , .A2( u2_u2_X_23 ) , .ZN( u2_u2_u3_n154 ) );
  NAND2_X1 u2_u2_u3_U77 (.A1( u2_u2_X_23 ) , .ZN( u2_u2_u3_n149 ) , .A2( u2_u2_u3_n166 ) );
  NOR2_X1 u2_u2_u3_U78 (.A2( u2_u2_X_22 ) , .A1( u2_u2_X_23 ) , .ZN( u2_u2_u3_n121 ) );
  AND2_X1 u2_u2_u3_U79 (.A1( u2_u2_X_24 ) , .ZN( u2_u2_u3_n101 ) , .A2( u2_u2_u3_n171 ) );
  AND3_X1 u2_u2_u3_U8 (.A3( u2_u2_u3_n144 ) , .A2( u2_u2_u3_n145 ) , .A1( u2_u2_u3_n146 ) , .ZN( u2_u2_u3_n147 ) );
  AND2_X1 u2_u2_u3_U80 (.A1( u2_u2_X_19 ) , .ZN( u2_u2_u3_n102 ) , .A2( u2_u2_u3_n172 ) );
  AND2_X1 u2_u2_u3_U81 (.A1( u2_u2_X_21 ) , .A2( u2_u2_X_24 ) , .ZN( u2_u2_u3_n100 ) );
  AND2_X1 u2_u2_u3_U82 (.A2( u2_u2_X_19 ) , .A1( u2_u2_X_20 ) , .ZN( u2_u2_u3_n104 ) );
  INV_X1 u2_u2_u3_U83 (.A( u2_u2_X_22 ) , .ZN( u2_u2_u3_n166 ) );
  INV_X1 u2_u2_u3_U84 (.A( u2_u2_X_21 ) , .ZN( u2_u2_u3_n171 ) );
  INV_X1 u2_u2_u3_U85 (.A( u2_u2_X_20 ) , .ZN( u2_u2_u3_n172 ) );
  OR4_X1 u2_u2_u3_U86 (.ZN( u2_out2_10 ) , .A4( u2_u2_u3_n136 ) , .A3( u2_u2_u3_n137 ) , .A1( u2_u2_u3_n138 ) , .A2( u2_u2_u3_n139 ) );
  OAI222_X1 u2_u2_u3_U87 (.C1( u2_u2_u3_n128 ) , .ZN( u2_u2_u3_n137 ) , .B1( u2_u2_u3_n148 ) , .A2( u2_u2_u3_n150 ) , .B2( u2_u2_u3_n154 ) , .C2( u2_u2_u3_n164 ) , .A1( u2_u2_u3_n167 ) );
  OAI221_X1 u2_u2_u3_U88 (.A( u2_u2_u3_n134 ) , .B2( u2_u2_u3_n135 ) , .ZN( u2_u2_u3_n136 ) , .C1( u2_u2_u3_n149 ) , .B1( u2_u2_u3_n151 ) , .C2( u2_u2_u3_n183 ) );
  NAND4_X1 u2_u2_u3_U89 (.ZN( u2_out2_26 ) , .A4( u2_u2_u3_n109 ) , .A3( u2_u2_u3_n110 ) , .A2( u2_u2_u3_n111 ) , .A1( u2_u2_u3_n173 ) );
  INV_X1 u2_u2_u3_U9 (.A( u2_u2_u3_n143 ) , .ZN( u2_u2_u3_n168 ) );
  INV_X1 u2_u2_u3_U90 (.ZN( u2_u2_u3_n173 ) , .A( u2_u2_u3_n94 ) );
  OAI21_X1 u2_u2_u3_U91 (.ZN( u2_u2_u3_n111 ) , .B2( u2_u2_u3_n117 ) , .A( u2_u2_u3_n133 ) , .B1( u2_u2_u3_n176 ) );
  NAND4_X1 u2_u2_u3_U92 (.ZN( u2_out2_20 ) , .A4( u2_u2_u3_n122 ) , .A3( u2_u2_u3_n123 ) , .A1( u2_u2_u3_n175 ) , .A2( u2_u2_u3_n180 ) );
  INV_X1 u2_u2_u3_U93 (.A( u2_u2_u3_n112 ) , .ZN( u2_u2_u3_n175 ) );
  INV_X1 u2_u2_u3_U94 (.A( u2_u2_u3_n126 ) , .ZN( u2_u2_u3_n180 ) );
  NAND4_X1 u2_u2_u3_U95 (.ZN( u2_out2_1 ) , .A4( u2_u2_u3_n161 ) , .A3( u2_u2_u3_n162 ) , .A2( u2_u2_u3_n163 ) , .A1( u2_u2_u3_n185 ) );
  NAND2_X1 u2_u2_u3_U96 (.ZN( u2_u2_u3_n163 ) , .A2( u2_u2_u3_n170 ) , .A1( u2_u2_u3_n176 ) );
  AOI22_X1 u2_u2_u3_U97 (.B2( u2_u2_u3_n140 ) , .B1( u2_u2_u3_n141 ) , .A2( u2_u2_u3_n142 ) , .ZN( u2_u2_u3_n162 ) , .A1( u2_u2_u3_n177 ) );
  NAND3_X1 u2_u2_u3_U98 (.A1( u2_u2_u3_n114 ) , .ZN( u2_u2_u3_n115 ) , .A2( u2_u2_u3_n145 ) , .A3( u2_u2_u3_n153 ) );
  NAND3_X1 u2_u2_u3_U99 (.ZN( u2_u2_u3_n129 ) , .A2( u2_u2_u3_n144 ) , .A1( u2_u2_u3_n153 ) , .A3( u2_u2_u3_n182 ) );
  OAI22_X1 u2_u2_u4_U10 (.B2( u2_u2_u4_n135 ) , .ZN( u2_u2_u4_n137 ) , .B1( u2_u2_u4_n153 ) , .A1( u2_u2_u4_n155 ) , .A2( u2_u2_u4_n171 ) );
  AND3_X1 u2_u2_u4_U11 (.A2( u2_u2_u4_n134 ) , .ZN( u2_u2_u4_n135 ) , .A3( u2_u2_u4_n145 ) , .A1( u2_u2_u4_n157 ) );
  NAND2_X1 u2_u2_u4_U12 (.ZN( u2_u2_u4_n132 ) , .A2( u2_u2_u4_n170 ) , .A1( u2_u2_u4_n173 ) );
  AOI21_X1 u2_u2_u4_U13 (.B2( u2_u2_u4_n160 ) , .B1( u2_u2_u4_n161 ) , .ZN( u2_u2_u4_n162 ) , .A( u2_u2_u4_n170 ) );
  AOI21_X1 u2_u2_u4_U14 (.ZN( u2_u2_u4_n107 ) , .B2( u2_u2_u4_n143 ) , .A( u2_u2_u4_n174 ) , .B1( u2_u2_u4_n184 ) );
  AOI21_X1 u2_u2_u4_U15 (.B2( u2_u2_u4_n158 ) , .B1( u2_u2_u4_n159 ) , .ZN( u2_u2_u4_n163 ) , .A( u2_u2_u4_n174 ) );
  AOI21_X1 u2_u2_u4_U16 (.A( u2_u2_u4_n153 ) , .B2( u2_u2_u4_n154 ) , .B1( u2_u2_u4_n155 ) , .ZN( u2_u2_u4_n165 ) );
  AOI21_X1 u2_u2_u4_U17 (.A( u2_u2_u4_n156 ) , .B2( u2_u2_u4_n157 ) , .ZN( u2_u2_u4_n164 ) , .B1( u2_u2_u4_n184 ) );
  INV_X1 u2_u2_u4_U18 (.A( u2_u2_u4_n138 ) , .ZN( u2_u2_u4_n170 ) );
  AND2_X1 u2_u2_u4_U19 (.A2( u2_u2_u4_n120 ) , .ZN( u2_u2_u4_n155 ) , .A1( u2_u2_u4_n160 ) );
  INV_X1 u2_u2_u4_U20 (.A( u2_u2_u4_n156 ) , .ZN( u2_u2_u4_n175 ) );
  NAND2_X1 u2_u2_u4_U21 (.A2( u2_u2_u4_n118 ) , .ZN( u2_u2_u4_n131 ) , .A1( u2_u2_u4_n147 ) );
  NAND2_X1 u2_u2_u4_U22 (.A1( u2_u2_u4_n119 ) , .A2( u2_u2_u4_n120 ) , .ZN( u2_u2_u4_n130 ) );
  NAND2_X1 u2_u2_u4_U23 (.ZN( u2_u2_u4_n117 ) , .A2( u2_u2_u4_n118 ) , .A1( u2_u2_u4_n148 ) );
  NAND2_X1 u2_u2_u4_U24 (.ZN( u2_u2_u4_n129 ) , .A1( u2_u2_u4_n134 ) , .A2( u2_u2_u4_n148 ) );
  AND3_X1 u2_u2_u4_U25 (.A1( u2_u2_u4_n119 ) , .A2( u2_u2_u4_n143 ) , .A3( u2_u2_u4_n154 ) , .ZN( u2_u2_u4_n161 ) );
  AND2_X1 u2_u2_u4_U26 (.A1( u2_u2_u4_n145 ) , .A2( u2_u2_u4_n147 ) , .ZN( u2_u2_u4_n159 ) );
  OR3_X1 u2_u2_u4_U27 (.A3( u2_u2_u4_n114 ) , .A2( u2_u2_u4_n115 ) , .A1( u2_u2_u4_n116 ) , .ZN( u2_u2_u4_n136 ) );
  AOI21_X1 u2_u2_u4_U28 (.A( u2_u2_u4_n113 ) , .ZN( u2_u2_u4_n116 ) , .B2( u2_u2_u4_n173 ) , .B1( u2_u2_u4_n174 ) );
  AOI21_X1 u2_u2_u4_U29 (.ZN( u2_u2_u4_n115 ) , .B2( u2_u2_u4_n145 ) , .B1( u2_u2_u4_n146 ) , .A( u2_u2_u4_n156 ) );
  NOR2_X1 u2_u2_u4_U3 (.ZN( u2_u2_u4_n121 ) , .A1( u2_u2_u4_n181 ) , .A2( u2_u2_u4_n182 ) );
  OAI22_X1 u2_u2_u4_U30 (.ZN( u2_u2_u4_n114 ) , .A2( u2_u2_u4_n121 ) , .B1( u2_u2_u4_n160 ) , .B2( u2_u2_u4_n170 ) , .A1( u2_u2_u4_n171 ) );
  INV_X1 u2_u2_u4_U31 (.A( u2_u2_u4_n158 ) , .ZN( u2_u2_u4_n182 ) );
  INV_X1 u2_u2_u4_U32 (.ZN( u2_u2_u4_n181 ) , .A( u2_u2_u4_n96 ) );
  INV_X1 u2_u2_u4_U33 (.A( u2_u2_u4_n144 ) , .ZN( u2_u2_u4_n179 ) );
  INV_X1 u2_u2_u4_U34 (.A( u2_u2_u4_n157 ) , .ZN( u2_u2_u4_n178 ) );
  NAND2_X1 u2_u2_u4_U35 (.A2( u2_u2_u4_n154 ) , .A1( u2_u2_u4_n96 ) , .ZN( u2_u2_u4_n97 ) );
  INV_X1 u2_u2_u4_U36 (.ZN( u2_u2_u4_n186 ) , .A( u2_u2_u4_n95 ) );
  OAI221_X1 u2_u2_u4_U37 (.C1( u2_u2_u4_n134 ) , .B1( u2_u2_u4_n158 ) , .B2( u2_u2_u4_n171 ) , .C2( u2_u2_u4_n173 ) , .A( u2_u2_u4_n94 ) , .ZN( u2_u2_u4_n95 ) );
  AOI222_X1 u2_u2_u4_U38 (.B2( u2_u2_u4_n132 ) , .A1( u2_u2_u4_n138 ) , .C2( u2_u2_u4_n175 ) , .A2( u2_u2_u4_n179 ) , .C1( u2_u2_u4_n181 ) , .B1( u2_u2_u4_n185 ) , .ZN( u2_u2_u4_n94 ) );
  INV_X1 u2_u2_u4_U39 (.A( u2_u2_u4_n113 ) , .ZN( u2_u2_u4_n185 ) );
  INV_X1 u2_u2_u4_U4 (.A( u2_u2_u4_n117 ) , .ZN( u2_u2_u4_n184 ) );
  INV_X1 u2_u2_u4_U40 (.A( u2_u2_u4_n143 ) , .ZN( u2_u2_u4_n183 ) );
  NOR2_X1 u2_u2_u4_U41 (.ZN( u2_u2_u4_n138 ) , .A1( u2_u2_u4_n168 ) , .A2( u2_u2_u4_n169 ) );
  NOR2_X1 u2_u2_u4_U42 (.A1( u2_u2_u4_n150 ) , .A2( u2_u2_u4_n152 ) , .ZN( u2_u2_u4_n153 ) );
  NOR2_X1 u2_u2_u4_U43 (.A2( u2_u2_u4_n128 ) , .A1( u2_u2_u4_n138 ) , .ZN( u2_u2_u4_n156 ) );
  AOI22_X1 u2_u2_u4_U44 (.B2( u2_u2_u4_n122 ) , .A1( u2_u2_u4_n123 ) , .ZN( u2_u2_u4_n124 ) , .B1( u2_u2_u4_n128 ) , .A2( u2_u2_u4_n172 ) );
  INV_X1 u2_u2_u4_U45 (.A( u2_u2_u4_n153 ) , .ZN( u2_u2_u4_n172 ) );
  NAND2_X1 u2_u2_u4_U46 (.A2( u2_u2_u4_n120 ) , .ZN( u2_u2_u4_n123 ) , .A1( u2_u2_u4_n161 ) );
  AOI22_X1 u2_u2_u4_U47 (.B2( u2_u2_u4_n132 ) , .A2( u2_u2_u4_n133 ) , .ZN( u2_u2_u4_n140 ) , .A1( u2_u2_u4_n150 ) , .B1( u2_u2_u4_n179 ) );
  NAND2_X1 u2_u2_u4_U48 (.ZN( u2_u2_u4_n133 ) , .A2( u2_u2_u4_n146 ) , .A1( u2_u2_u4_n154 ) );
  NAND2_X1 u2_u2_u4_U49 (.A1( u2_u2_u4_n103 ) , .ZN( u2_u2_u4_n154 ) , .A2( u2_u2_u4_n98 ) );
  NOR4_X1 u2_u2_u4_U5 (.A4( u2_u2_u4_n106 ) , .A3( u2_u2_u4_n107 ) , .A2( u2_u2_u4_n108 ) , .A1( u2_u2_u4_n109 ) , .ZN( u2_u2_u4_n110 ) );
  NAND2_X1 u2_u2_u4_U50 (.A1( u2_u2_u4_n101 ) , .ZN( u2_u2_u4_n158 ) , .A2( u2_u2_u4_n99 ) );
  AOI21_X1 u2_u2_u4_U51 (.ZN( u2_u2_u4_n127 ) , .A( u2_u2_u4_n136 ) , .B2( u2_u2_u4_n150 ) , .B1( u2_u2_u4_n180 ) );
  INV_X1 u2_u2_u4_U52 (.A( u2_u2_u4_n160 ) , .ZN( u2_u2_u4_n180 ) );
  NAND2_X1 u2_u2_u4_U53 (.A2( u2_u2_u4_n104 ) , .A1( u2_u2_u4_n105 ) , .ZN( u2_u2_u4_n146 ) );
  NAND2_X1 u2_u2_u4_U54 (.A2( u2_u2_u4_n101 ) , .A1( u2_u2_u4_n102 ) , .ZN( u2_u2_u4_n160 ) );
  NAND2_X1 u2_u2_u4_U55 (.ZN( u2_u2_u4_n134 ) , .A1( u2_u2_u4_n98 ) , .A2( u2_u2_u4_n99 ) );
  NAND2_X1 u2_u2_u4_U56 (.A1( u2_u2_u4_n103 ) , .A2( u2_u2_u4_n104 ) , .ZN( u2_u2_u4_n143 ) );
  NAND2_X1 u2_u2_u4_U57 (.A2( u2_u2_u4_n105 ) , .ZN( u2_u2_u4_n145 ) , .A1( u2_u2_u4_n98 ) );
  NAND2_X1 u2_u2_u4_U58 (.A1( u2_u2_u4_n100 ) , .A2( u2_u2_u4_n105 ) , .ZN( u2_u2_u4_n120 ) );
  NAND2_X1 u2_u2_u4_U59 (.A1( u2_u2_u4_n102 ) , .A2( u2_u2_u4_n104 ) , .ZN( u2_u2_u4_n148 ) );
  AOI21_X1 u2_u2_u4_U6 (.ZN( u2_u2_u4_n106 ) , .B2( u2_u2_u4_n146 ) , .B1( u2_u2_u4_n158 ) , .A( u2_u2_u4_n170 ) );
  NAND2_X1 u2_u2_u4_U60 (.A2( u2_u2_u4_n100 ) , .A1( u2_u2_u4_n103 ) , .ZN( u2_u2_u4_n157 ) );
  INV_X1 u2_u2_u4_U61 (.A( u2_u2_u4_n150 ) , .ZN( u2_u2_u4_n173 ) );
  INV_X1 u2_u2_u4_U62 (.A( u2_u2_u4_n152 ) , .ZN( u2_u2_u4_n171 ) );
  NAND2_X1 u2_u2_u4_U63 (.A1( u2_u2_u4_n100 ) , .ZN( u2_u2_u4_n118 ) , .A2( u2_u2_u4_n99 ) );
  NAND2_X1 u2_u2_u4_U64 (.A2( u2_u2_u4_n100 ) , .A1( u2_u2_u4_n102 ) , .ZN( u2_u2_u4_n144 ) );
  NAND2_X1 u2_u2_u4_U65 (.A2( u2_u2_u4_n101 ) , .A1( u2_u2_u4_n105 ) , .ZN( u2_u2_u4_n96 ) );
  INV_X1 u2_u2_u4_U66 (.A( u2_u2_u4_n128 ) , .ZN( u2_u2_u4_n174 ) );
  NAND2_X1 u2_u2_u4_U67 (.A2( u2_u2_u4_n102 ) , .ZN( u2_u2_u4_n119 ) , .A1( u2_u2_u4_n98 ) );
  NAND2_X1 u2_u2_u4_U68 (.A2( u2_u2_u4_n101 ) , .A1( u2_u2_u4_n103 ) , .ZN( u2_u2_u4_n147 ) );
  NAND2_X1 u2_u2_u4_U69 (.A2( u2_u2_u4_n104 ) , .ZN( u2_u2_u4_n113 ) , .A1( u2_u2_u4_n99 ) );
  AOI21_X1 u2_u2_u4_U7 (.ZN( u2_u2_u4_n108 ) , .B2( u2_u2_u4_n134 ) , .B1( u2_u2_u4_n155 ) , .A( u2_u2_u4_n156 ) );
  NOR2_X1 u2_u2_u4_U70 (.A2( u2_u2_X_28 ) , .ZN( u2_u2_u4_n150 ) , .A1( u2_u2_u4_n168 ) );
  NOR2_X1 u2_u2_u4_U71 (.A2( u2_u2_X_29 ) , .ZN( u2_u2_u4_n152 ) , .A1( u2_u2_u4_n169 ) );
  NOR2_X1 u2_u2_u4_U72 (.A2( u2_u2_X_30 ) , .ZN( u2_u2_u4_n105 ) , .A1( u2_u2_u4_n176 ) );
  NOR2_X1 u2_u2_u4_U73 (.A2( u2_u2_X_26 ) , .ZN( u2_u2_u4_n100 ) , .A1( u2_u2_u4_n177 ) );
  NOR2_X1 u2_u2_u4_U74 (.A2( u2_u2_X_28 ) , .A1( u2_u2_X_29 ) , .ZN( u2_u2_u4_n128 ) );
  NOR2_X1 u2_u2_u4_U75 (.A2( u2_u2_X_27 ) , .A1( u2_u2_X_30 ) , .ZN( u2_u2_u4_n102 ) );
  NOR2_X1 u2_u2_u4_U76 (.A2( u2_u2_X_25 ) , .A1( u2_u2_X_26 ) , .ZN( u2_u2_u4_n98 ) );
  AND2_X1 u2_u2_u4_U77 (.A2( u2_u2_X_25 ) , .A1( u2_u2_X_26 ) , .ZN( u2_u2_u4_n104 ) );
  AND2_X1 u2_u2_u4_U78 (.A1( u2_u2_X_30 ) , .A2( u2_u2_u4_n176 ) , .ZN( u2_u2_u4_n99 ) );
  AND2_X1 u2_u2_u4_U79 (.A1( u2_u2_X_26 ) , .ZN( u2_u2_u4_n101 ) , .A2( u2_u2_u4_n177 ) );
  AOI21_X1 u2_u2_u4_U8 (.ZN( u2_u2_u4_n109 ) , .A( u2_u2_u4_n153 ) , .B1( u2_u2_u4_n159 ) , .B2( u2_u2_u4_n184 ) );
  AND2_X1 u2_u2_u4_U80 (.A1( u2_u2_X_27 ) , .A2( u2_u2_X_30 ) , .ZN( u2_u2_u4_n103 ) );
  INV_X1 u2_u2_u4_U81 (.A( u2_u2_X_28 ) , .ZN( u2_u2_u4_n169 ) );
  INV_X1 u2_u2_u4_U82 (.A( u2_u2_X_29 ) , .ZN( u2_u2_u4_n168 ) );
  INV_X1 u2_u2_u4_U83 (.A( u2_u2_X_25 ) , .ZN( u2_u2_u4_n177 ) );
  INV_X1 u2_u2_u4_U84 (.A( u2_u2_X_27 ) , .ZN( u2_u2_u4_n176 ) );
  NAND4_X1 u2_u2_u4_U85 (.ZN( u2_out2_25 ) , .A4( u2_u2_u4_n139 ) , .A3( u2_u2_u4_n140 ) , .A2( u2_u2_u4_n141 ) , .A1( u2_u2_u4_n142 ) );
  OAI21_X1 u2_u2_u4_U86 (.A( u2_u2_u4_n128 ) , .B2( u2_u2_u4_n129 ) , .B1( u2_u2_u4_n130 ) , .ZN( u2_u2_u4_n142 ) );
  OAI21_X1 u2_u2_u4_U87 (.B2( u2_u2_u4_n131 ) , .ZN( u2_u2_u4_n141 ) , .A( u2_u2_u4_n175 ) , .B1( u2_u2_u4_n183 ) );
  NAND4_X1 u2_u2_u4_U88 (.ZN( u2_out2_14 ) , .A4( u2_u2_u4_n124 ) , .A3( u2_u2_u4_n125 ) , .A2( u2_u2_u4_n126 ) , .A1( u2_u2_u4_n127 ) );
  AOI22_X1 u2_u2_u4_U89 (.B2( u2_u2_u4_n117 ) , .ZN( u2_u2_u4_n126 ) , .A1( u2_u2_u4_n129 ) , .B1( u2_u2_u4_n152 ) , .A2( u2_u2_u4_n175 ) );
  AOI211_X1 u2_u2_u4_U9 (.B( u2_u2_u4_n136 ) , .A( u2_u2_u4_n137 ) , .C2( u2_u2_u4_n138 ) , .ZN( u2_u2_u4_n139 ) , .C1( u2_u2_u4_n182 ) );
  AOI22_X1 u2_u2_u4_U90 (.ZN( u2_u2_u4_n125 ) , .B2( u2_u2_u4_n131 ) , .A2( u2_u2_u4_n132 ) , .B1( u2_u2_u4_n138 ) , .A1( u2_u2_u4_n178 ) );
  NAND4_X1 u2_u2_u4_U91 (.ZN( u2_out2_8 ) , .A4( u2_u2_u4_n110 ) , .A3( u2_u2_u4_n111 ) , .A2( u2_u2_u4_n112 ) , .A1( u2_u2_u4_n186 ) );
  NAND2_X1 u2_u2_u4_U92 (.ZN( u2_u2_u4_n112 ) , .A2( u2_u2_u4_n130 ) , .A1( u2_u2_u4_n150 ) );
  AOI22_X1 u2_u2_u4_U93 (.ZN( u2_u2_u4_n111 ) , .B2( u2_u2_u4_n132 ) , .A1( u2_u2_u4_n152 ) , .B1( u2_u2_u4_n178 ) , .A2( u2_u2_u4_n97 ) );
  AOI22_X1 u2_u2_u4_U94 (.B2( u2_u2_u4_n149 ) , .B1( u2_u2_u4_n150 ) , .A2( u2_u2_u4_n151 ) , .A1( u2_u2_u4_n152 ) , .ZN( u2_u2_u4_n167 ) );
  NOR4_X1 u2_u2_u4_U95 (.A4( u2_u2_u4_n162 ) , .A3( u2_u2_u4_n163 ) , .A2( u2_u2_u4_n164 ) , .A1( u2_u2_u4_n165 ) , .ZN( u2_u2_u4_n166 ) );
  NAND3_X1 u2_u2_u4_U96 (.ZN( u2_out2_3 ) , .A3( u2_u2_u4_n166 ) , .A1( u2_u2_u4_n167 ) , .A2( u2_u2_u4_n186 ) );
  NAND3_X1 u2_u2_u4_U97 (.A3( u2_u2_u4_n146 ) , .A2( u2_u2_u4_n147 ) , .A1( u2_u2_u4_n148 ) , .ZN( u2_u2_u4_n149 ) );
  NAND3_X1 u2_u2_u4_U98 (.A3( u2_u2_u4_n143 ) , .A2( u2_u2_u4_n144 ) , .A1( u2_u2_u4_n145 ) , .ZN( u2_u2_u4_n151 ) );
  NAND3_X1 u2_u2_u4_U99 (.A3( u2_u2_u4_n121 ) , .ZN( u2_u2_u4_n122 ) , .A2( u2_u2_u4_n144 ) , .A1( u2_u2_u4_n154 ) );
  INV_X1 u2_u2_u5_U10 (.A( u2_u2_u5_n121 ) , .ZN( u2_u2_u5_n177 ) );
  NOR3_X1 u2_u2_u5_U100 (.A3( u2_u2_u5_n141 ) , .A1( u2_u2_u5_n142 ) , .ZN( u2_u2_u5_n143 ) , .A2( u2_u2_u5_n191 ) );
  NAND4_X1 u2_u2_u5_U101 (.ZN( u2_out2_4 ) , .A4( u2_u2_u5_n112 ) , .A2( u2_u2_u5_n113 ) , .A1( u2_u2_u5_n114 ) , .A3( u2_u2_u5_n195 ) );
  AOI211_X1 u2_u2_u5_U102 (.A( u2_u2_u5_n110 ) , .C1( u2_u2_u5_n111 ) , .ZN( u2_u2_u5_n112 ) , .B( u2_u2_u5_n118 ) , .C2( u2_u2_u5_n177 ) );
  AOI222_X1 u2_u2_u5_U103 (.ZN( u2_u2_u5_n113 ) , .A1( u2_u2_u5_n131 ) , .C1( u2_u2_u5_n148 ) , .B2( u2_u2_u5_n174 ) , .C2( u2_u2_u5_n178 ) , .A2( u2_u2_u5_n179 ) , .B1( u2_u2_u5_n99 ) );
  NAND3_X1 u2_u2_u5_U104 (.A2( u2_u2_u5_n154 ) , .A3( u2_u2_u5_n158 ) , .A1( u2_u2_u5_n161 ) , .ZN( u2_u2_u5_n99 ) );
  NOR2_X1 u2_u2_u5_U11 (.ZN( u2_u2_u5_n160 ) , .A2( u2_u2_u5_n173 ) , .A1( u2_u2_u5_n177 ) );
  INV_X1 u2_u2_u5_U12 (.A( u2_u2_u5_n150 ) , .ZN( u2_u2_u5_n174 ) );
  AOI21_X1 u2_u2_u5_U13 (.A( u2_u2_u5_n160 ) , .B2( u2_u2_u5_n161 ) , .ZN( u2_u2_u5_n162 ) , .B1( u2_u2_u5_n192 ) );
  INV_X1 u2_u2_u5_U14 (.A( u2_u2_u5_n159 ) , .ZN( u2_u2_u5_n192 ) );
  AOI21_X1 u2_u2_u5_U15 (.A( u2_u2_u5_n156 ) , .B2( u2_u2_u5_n157 ) , .B1( u2_u2_u5_n158 ) , .ZN( u2_u2_u5_n163 ) );
  AOI21_X1 u2_u2_u5_U16 (.B2( u2_u2_u5_n139 ) , .B1( u2_u2_u5_n140 ) , .ZN( u2_u2_u5_n141 ) , .A( u2_u2_u5_n150 ) );
  OAI21_X1 u2_u2_u5_U17 (.A( u2_u2_u5_n133 ) , .B2( u2_u2_u5_n134 ) , .B1( u2_u2_u5_n135 ) , .ZN( u2_u2_u5_n142 ) );
  OAI21_X1 u2_u2_u5_U18 (.ZN( u2_u2_u5_n133 ) , .B2( u2_u2_u5_n147 ) , .A( u2_u2_u5_n173 ) , .B1( u2_u2_u5_n188 ) );
  NAND2_X1 u2_u2_u5_U19 (.A2( u2_u2_u5_n119 ) , .A1( u2_u2_u5_n123 ) , .ZN( u2_u2_u5_n137 ) );
  INV_X1 u2_u2_u5_U20 (.A( u2_u2_u5_n155 ) , .ZN( u2_u2_u5_n194 ) );
  NAND2_X1 u2_u2_u5_U21 (.A1( u2_u2_u5_n121 ) , .ZN( u2_u2_u5_n132 ) , .A2( u2_u2_u5_n172 ) );
  NAND2_X1 u2_u2_u5_U22 (.A2( u2_u2_u5_n122 ) , .ZN( u2_u2_u5_n136 ) , .A1( u2_u2_u5_n154 ) );
  NAND2_X1 u2_u2_u5_U23 (.A2( u2_u2_u5_n119 ) , .A1( u2_u2_u5_n120 ) , .ZN( u2_u2_u5_n159 ) );
  INV_X1 u2_u2_u5_U24 (.A( u2_u2_u5_n156 ) , .ZN( u2_u2_u5_n175 ) );
  INV_X1 u2_u2_u5_U25 (.A( u2_u2_u5_n158 ) , .ZN( u2_u2_u5_n188 ) );
  INV_X1 u2_u2_u5_U26 (.A( u2_u2_u5_n152 ) , .ZN( u2_u2_u5_n179 ) );
  INV_X1 u2_u2_u5_U27 (.A( u2_u2_u5_n140 ) , .ZN( u2_u2_u5_n182 ) );
  INV_X1 u2_u2_u5_U28 (.A( u2_u2_u5_n151 ) , .ZN( u2_u2_u5_n183 ) );
  INV_X1 u2_u2_u5_U29 (.A( u2_u2_u5_n123 ) , .ZN( u2_u2_u5_n185 ) );
  NOR2_X1 u2_u2_u5_U3 (.ZN( u2_u2_u5_n134 ) , .A1( u2_u2_u5_n183 ) , .A2( u2_u2_u5_n190 ) );
  INV_X1 u2_u2_u5_U30 (.A( u2_u2_u5_n161 ) , .ZN( u2_u2_u5_n184 ) );
  INV_X1 u2_u2_u5_U31 (.A( u2_u2_u5_n139 ) , .ZN( u2_u2_u5_n189 ) );
  INV_X1 u2_u2_u5_U32 (.A( u2_u2_u5_n157 ) , .ZN( u2_u2_u5_n190 ) );
  INV_X1 u2_u2_u5_U33 (.A( u2_u2_u5_n120 ) , .ZN( u2_u2_u5_n193 ) );
  NAND2_X1 u2_u2_u5_U34 (.ZN( u2_u2_u5_n111 ) , .A1( u2_u2_u5_n140 ) , .A2( u2_u2_u5_n155 ) );
  INV_X1 u2_u2_u5_U35 (.A( u2_u2_u5_n117 ) , .ZN( u2_u2_u5_n196 ) );
  OAI221_X1 u2_u2_u5_U36 (.A( u2_u2_u5_n116 ) , .ZN( u2_u2_u5_n117 ) , .B2( u2_u2_u5_n119 ) , .C1( u2_u2_u5_n153 ) , .C2( u2_u2_u5_n158 ) , .B1( u2_u2_u5_n172 ) );
  AOI222_X1 u2_u2_u5_U37 (.ZN( u2_u2_u5_n116 ) , .B2( u2_u2_u5_n145 ) , .C1( u2_u2_u5_n148 ) , .A2( u2_u2_u5_n174 ) , .C2( u2_u2_u5_n177 ) , .B1( u2_u2_u5_n187 ) , .A1( u2_u2_u5_n193 ) );
  INV_X1 u2_u2_u5_U38 (.A( u2_u2_u5_n115 ) , .ZN( u2_u2_u5_n187 ) );
  NOR2_X1 u2_u2_u5_U39 (.ZN( u2_u2_u5_n100 ) , .A1( u2_u2_u5_n170 ) , .A2( u2_u2_u5_n180 ) );
  INV_X1 u2_u2_u5_U4 (.A( u2_u2_u5_n138 ) , .ZN( u2_u2_u5_n191 ) );
  AOI22_X1 u2_u2_u5_U40 (.B2( u2_u2_u5_n131 ) , .A2( u2_u2_u5_n146 ) , .ZN( u2_u2_u5_n169 ) , .B1( u2_u2_u5_n174 ) , .A1( u2_u2_u5_n185 ) );
  NOR2_X1 u2_u2_u5_U41 (.A1( u2_u2_u5_n146 ) , .ZN( u2_u2_u5_n150 ) , .A2( u2_u2_u5_n173 ) );
  AOI21_X1 u2_u2_u5_U42 (.A( u2_u2_u5_n118 ) , .B2( u2_u2_u5_n145 ) , .ZN( u2_u2_u5_n168 ) , .B1( u2_u2_u5_n186 ) );
  INV_X1 u2_u2_u5_U43 (.A( u2_u2_u5_n122 ) , .ZN( u2_u2_u5_n186 ) );
  NOR2_X1 u2_u2_u5_U44 (.A1( u2_u2_u5_n146 ) , .ZN( u2_u2_u5_n152 ) , .A2( u2_u2_u5_n176 ) );
  NOR2_X1 u2_u2_u5_U45 (.A1( u2_u2_u5_n115 ) , .ZN( u2_u2_u5_n118 ) , .A2( u2_u2_u5_n153 ) );
  NOR2_X1 u2_u2_u5_U46 (.A2( u2_u2_u5_n145 ) , .ZN( u2_u2_u5_n156 ) , .A1( u2_u2_u5_n174 ) );
  NOR2_X1 u2_u2_u5_U47 (.ZN( u2_u2_u5_n121 ) , .A2( u2_u2_u5_n145 ) , .A1( u2_u2_u5_n176 ) );
  AOI22_X1 u2_u2_u5_U48 (.ZN( u2_u2_u5_n114 ) , .A2( u2_u2_u5_n137 ) , .A1( u2_u2_u5_n145 ) , .B2( u2_u2_u5_n175 ) , .B1( u2_u2_u5_n193 ) );
  AOI21_X1 u2_u2_u5_U49 (.A( u2_u2_u5_n153 ) , .B2( u2_u2_u5_n154 ) , .B1( u2_u2_u5_n155 ) , .ZN( u2_u2_u5_n164 ) );
  OAI21_X1 u2_u2_u5_U5 (.B2( u2_u2_u5_n136 ) , .B1( u2_u2_u5_n137 ) , .ZN( u2_u2_u5_n138 ) , .A( u2_u2_u5_n177 ) );
  AOI21_X1 u2_u2_u5_U50 (.ZN( u2_u2_u5_n110 ) , .B1( u2_u2_u5_n122 ) , .B2( u2_u2_u5_n139 ) , .A( u2_u2_u5_n153 ) );
  INV_X1 u2_u2_u5_U51 (.A( u2_u2_u5_n153 ) , .ZN( u2_u2_u5_n176 ) );
  INV_X1 u2_u2_u5_U52 (.A( u2_u2_u5_n126 ) , .ZN( u2_u2_u5_n173 ) );
  AND2_X1 u2_u2_u5_U53 (.A2( u2_u2_u5_n104 ) , .A1( u2_u2_u5_n107 ) , .ZN( u2_u2_u5_n147 ) );
  AND2_X1 u2_u2_u5_U54 (.A2( u2_u2_u5_n104 ) , .A1( u2_u2_u5_n108 ) , .ZN( u2_u2_u5_n148 ) );
  NAND2_X1 u2_u2_u5_U55 (.A1( u2_u2_u5_n105 ) , .A2( u2_u2_u5_n106 ) , .ZN( u2_u2_u5_n158 ) );
  NAND2_X1 u2_u2_u5_U56 (.A2( u2_u2_u5_n108 ) , .A1( u2_u2_u5_n109 ) , .ZN( u2_u2_u5_n139 ) );
  NAND2_X1 u2_u2_u5_U57 (.A1( u2_u2_u5_n106 ) , .A2( u2_u2_u5_n108 ) , .ZN( u2_u2_u5_n119 ) );
  OAI211_X1 u2_u2_u5_U58 (.B( u2_u2_u5_n124 ) , .A( u2_u2_u5_n125 ) , .C2( u2_u2_u5_n126 ) , .C1( u2_u2_u5_n127 ) , .ZN( u2_u2_u5_n128 ) );
  NOR3_X1 u2_u2_u5_U59 (.ZN( u2_u2_u5_n127 ) , .A1( u2_u2_u5_n136 ) , .A3( u2_u2_u5_n148 ) , .A2( u2_u2_u5_n182 ) );
  INV_X1 u2_u2_u5_U6 (.A( u2_u2_u5_n135 ) , .ZN( u2_u2_u5_n178 ) );
  OAI21_X1 u2_u2_u5_U60 (.ZN( u2_u2_u5_n124 ) , .A( u2_u2_u5_n177 ) , .B2( u2_u2_u5_n183 ) , .B1( u2_u2_u5_n189 ) );
  OAI21_X1 u2_u2_u5_U61 (.ZN( u2_u2_u5_n125 ) , .A( u2_u2_u5_n174 ) , .B2( u2_u2_u5_n185 ) , .B1( u2_u2_u5_n190 ) );
  NAND2_X1 u2_u2_u5_U62 (.A2( u2_u2_u5_n103 ) , .A1( u2_u2_u5_n105 ) , .ZN( u2_u2_u5_n140 ) );
  NAND2_X1 u2_u2_u5_U63 (.A2( u2_u2_u5_n104 ) , .A1( u2_u2_u5_n105 ) , .ZN( u2_u2_u5_n155 ) );
  NAND2_X1 u2_u2_u5_U64 (.A2( u2_u2_u5_n106 ) , .A1( u2_u2_u5_n107 ) , .ZN( u2_u2_u5_n122 ) );
  NAND2_X1 u2_u2_u5_U65 (.A2( u2_u2_u5_n100 ) , .A1( u2_u2_u5_n106 ) , .ZN( u2_u2_u5_n115 ) );
  NAND2_X1 u2_u2_u5_U66 (.A2( u2_u2_u5_n100 ) , .A1( u2_u2_u5_n103 ) , .ZN( u2_u2_u5_n161 ) );
  NAND2_X1 u2_u2_u5_U67 (.A1( u2_u2_u5_n105 ) , .A2( u2_u2_u5_n109 ) , .ZN( u2_u2_u5_n154 ) );
  INV_X1 u2_u2_u5_U68 (.A( u2_u2_u5_n146 ) , .ZN( u2_u2_u5_n172 ) );
  NAND2_X1 u2_u2_u5_U69 (.A1( u2_u2_u5_n103 ) , .A2( u2_u2_u5_n108 ) , .ZN( u2_u2_u5_n123 ) );
  OAI22_X1 u2_u2_u5_U7 (.B2( u2_u2_u5_n149 ) , .B1( u2_u2_u5_n150 ) , .A2( u2_u2_u5_n151 ) , .A1( u2_u2_u5_n152 ) , .ZN( u2_u2_u5_n165 ) );
  NAND2_X1 u2_u2_u5_U70 (.A2( u2_u2_u5_n103 ) , .A1( u2_u2_u5_n107 ) , .ZN( u2_u2_u5_n151 ) );
  NAND2_X1 u2_u2_u5_U71 (.A2( u2_u2_u5_n107 ) , .A1( u2_u2_u5_n109 ) , .ZN( u2_u2_u5_n120 ) );
  NAND2_X1 u2_u2_u5_U72 (.A2( u2_u2_u5_n100 ) , .A1( u2_u2_u5_n109 ) , .ZN( u2_u2_u5_n157 ) );
  AND2_X1 u2_u2_u5_U73 (.A2( u2_u2_u5_n100 ) , .A1( u2_u2_u5_n104 ) , .ZN( u2_u2_u5_n131 ) );
  INV_X1 u2_u2_u5_U74 (.A( u2_u2_u5_n102 ) , .ZN( u2_u2_u5_n195 ) );
  OAI221_X1 u2_u2_u5_U75 (.A( u2_u2_u5_n101 ) , .ZN( u2_u2_u5_n102 ) , .C2( u2_u2_u5_n115 ) , .C1( u2_u2_u5_n126 ) , .B1( u2_u2_u5_n134 ) , .B2( u2_u2_u5_n160 ) );
  OAI21_X1 u2_u2_u5_U76 (.ZN( u2_u2_u5_n101 ) , .B1( u2_u2_u5_n137 ) , .A( u2_u2_u5_n146 ) , .B2( u2_u2_u5_n147 ) );
  NOR2_X1 u2_u2_u5_U77 (.A2( u2_u2_X_34 ) , .A1( u2_u2_X_35 ) , .ZN( u2_u2_u5_n145 ) );
  NOR2_X1 u2_u2_u5_U78 (.A2( u2_u2_X_34 ) , .ZN( u2_u2_u5_n146 ) , .A1( u2_u2_u5_n171 ) );
  NOR2_X1 u2_u2_u5_U79 (.A2( u2_u2_X_31 ) , .A1( u2_u2_X_32 ) , .ZN( u2_u2_u5_n103 ) );
  NOR3_X1 u2_u2_u5_U8 (.A2( u2_u2_u5_n147 ) , .A1( u2_u2_u5_n148 ) , .ZN( u2_u2_u5_n149 ) , .A3( u2_u2_u5_n194 ) );
  NOR2_X1 u2_u2_u5_U80 (.A2( u2_u2_X_36 ) , .ZN( u2_u2_u5_n105 ) , .A1( u2_u2_u5_n180 ) );
  NOR2_X1 u2_u2_u5_U81 (.A2( u2_u2_X_33 ) , .ZN( u2_u2_u5_n108 ) , .A1( u2_u2_u5_n170 ) );
  NOR2_X1 u2_u2_u5_U82 (.A2( u2_u2_X_33 ) , .A1( u2_u2_X_36 ) , .ZN( u2_u2_u5_n107 ) );
  NOR2_X1 u2_u2_u5_U83 (.A2( u2_u2_X_31 ) , .ZN( u2_u2_u5_n104 ) , .A1( u2_u2_u5_n181 ) );
  NAND2_X1 u2_u2_u5_U84 (.A2( u2_u2_X_34 ) , .A1( u2_u2_X_35 ) , .ZN( u2_u2_u5_n153 ) );
  NAND2_X1 u2_u2_u5_U85 (.A1( u2_u2_X_34 ) , .ZN( u2_u2_u5_n126 ) , .A2( u2_u2_u5_n171 ) );
  AND2_X1 u2_u2_u5_U86 (.A1( u2_u2_X_31 ) , .A2( u2_u2_X_32 ) , .ZN( u2_u2_u5_n106 ) );
  AND2_X1 u2_u2_u5_U87 (.A1( u2_u2_X_31 ) , .ZN( u2_u2_u5_n109 ) , .A2( u2_u2_u5_n181 ) );
  INV_X1 u2_u2_u5_U88 (.A( u2_u2_X_33 ) , .ZN( u2_u2_u5_n180 ) );
  INV_X1 u2_u2_u5_U89 (.A( u2_u2_X_35 ) , .ZN( u2_u2_u5_n171 ) );
  NOR2_X1 u2_u2_u5_U9 (.ZN( u2_u2_u5_n135 ) , .A1( u2_u2_u5_n173 ) , .A2( u2_u2_u5_n176 ) );
  INV_X1 u2_u2_u5_U90 (.A( u2_u2_X_36 ) , .ZN( u2_u2_u5_n170 ) );
  INV_X1 u2_u2_u5_U91 (.A( u2_u2_X_32 ) , .ZN( u2_u2_u5_n181 ) );
  NAND4_X1 u2_u2_u5_U92 (.ZN( u2_out2_29 ) , .A4( u2_u2_u5_n129 ) , .A3( u2_u2_u5_n130 ) , .A2( u2_u2_u5_n168 ) , .A1( u2_u2_u5_n196 ) );
  AOI221_X1 u2_u2_u5_U93 (.A( u2_u2_u5_n128 ) , .ZN( u2_u2_u5_n129 ) , .C2( u2_u2_u5_n132 ) , .B2( u2_u2_u5_n159 ) , .B1( u2_u2_u5_n176 ) , .C1( u2_u2_u5_n184 ) );
  AOI222_X1 u2_u2_u5_U94 (.ZN( u2_u2_u5_n130 ) , .A2( u2_u2_u5_n146 ) , .B1( u2_u2_u5_n147 ) , .C2( u2_u2_u5_n175 ) , .B2( u2_u2_u5_n179 ) , .A1( u2_u2_u5_n188 ) , .C1( u2_u2_u5_n194 ) );
  NAND4_X1 u2_u2_u5_U95 (.ZN( u2_out2_19 ) , .A4( u2_u2_u5_n166 ) , .A3( u2_u2_u5_n167 ) , .A2( u2_u2_u5_n168 ) , .A1( u2_u2_u5_n169 ) );
  AOI22_X1 u2_u2_u5_U96 (.B2( u2_u2_u5_n145 ) , .A2( u2_u2_u5_n146 ) , .ZN( u2_u2_u5_n167 ) , .B1( u2_u2_u5_n182 ) , .A1( u2_u2_u5_n189 ) );
  NOR4_X1 u2_u2_u5_U97 (.A4( u2_u2_u5_n162 ) , .A3( u2_u2_u5_n163 ) , .A2( u2_u2_u5_n164 ) , .A1( u2_u2_u5_n165 ) , .ZN( u2_u2_u5_n166 ) );
  NAND4_X1 u2_u2_u5_U98 (.ZN( u2_out2_11 ) , .A4( u2_u2_u5_n143 ) , .A3( u2_u2_u5_n144 ) , .A2( u2_u2_u5_n169 ) , .A1( u2_u2_u5_n196 ) );
  AOI22_X1 u2_u2_u5_U99 (.A2( u2_u2_u5_n132 ) , .ZN( u2_u2_u5_n144 ) , .B2( u2_u2_u5_n145 ) , .B1( u2_u2_u5_n184 ) , .A1( u2_u2_u5_n194 ) );
  OAI21_X1 u2_u2_u6_U10 (.A( u2_u2_u6_n159 ) , .B1( u2_u2_u6_n169 ) , .B2( u2_u2_u6_n173 ) , .ZN( u2_u2_u6_n90 ) );
  INV_X1 u2_u2_u6_U11 (.ZN( u2_u2_u6_n172 ) , .A( u2_u2_u6_n88 ) );
  AOI22_X1 u2_u2_u6_U12 (.A2( u2_u2_u6_n151 ) , .B2( u2_u2_u6_n161 ) , .A1( u2_u2_u6_n167 ) , .B1( u2_u2_u6_n170 ) , .ZN( u2_u2_u6_n89 ) );
  AOI21_X1 u2_u2_u6_U13 (.ZN( u2_u2_u6_n106 ) , .A( u2_u2_u6_n142 ) , .B2( u2_u2_u6_n159 ) , .B1( u2_u2_u6_n164 ) );
  INV_X1 u2_u2_u6_U14 (.A( u2_u2_u6_n155 ) , .ZN( u2_u2_u6_n161 ) );
  INV_X1 u2_u2_u6_U15 (.A( u2_u2_u6_n128 ) , .ZN( u2_u2_u6_n164 ) );
  NAND2_X1 u2_u2_u6_U16 (.ZN( u2_u2_u6_n110 ) , .A1( u2_u2_u6_n122 ) , .A2( u2_u2_u6_n129 ) );
  NAND2_X1 u2_u2_u6_U17 (.ZN( u2_u2_u6_n124 ) , .A2( u2_u2_u6_n146 ) , .A1( u2_u2_u6_n148 ) );
  INV_X1 u2_u2_u6_U18 (.A( u2_u2_u6_n132 ) , .ZN( u2_u2_u6_n171 ) );
  AND2_X1 u2_u2_u6_U19 (.A1( u2_u2_u6_n100 ) , .ZN( u2_u2_u6_n130 ) , .A2( u2_u2_u6_n147 ) );
  INV_X1 u2_u2_u6_U20 (.A( u2_u2_u6_n127 ) , .ZN( u2_u2_u6_n173 ) );
  INV_X1 u2_u2_u6_U21 (.A( u2_u2_u6_n121 ) , .ZN( u2_u2_u6_n167 ) );
  INV_X1 u2_u2_u6_U22 (.A( u2_u2_u6_n100 ) , .ZN( u2_u2_u6_n169 ) );
  INV_X1 u2_u2_u6_U23 (.A( u2_u2_u6_n123 ) , .ZN( u2_u2_u6_n170 ) );
  INV_X1 u2_u2_u6_U24 (.A( u2_u2_u6_n113 ) , .ZN( u2_u2_u6_n168 ) );
  AND2_X1 u2_u2_u6_U25 (.A1( u2_u2_u6_n107 ) , .A2( u2_u2_u6_n119 ) , .ZN( u2_u2_u6_n133 ) );
  AND2_X1 u2_u2_u6_U26 (.A2( u2_u2_u6_n121 ) , .A1( u2_u2_u6_n122 ) , .ZN( u2_u2_u6_n131 ) );
  AND3_X1 u2_u2_u6_U27 (.ZN( u2_u2_u6_n120 ) , .A2( u2_u2_u6_n127 ) , .A1( u2_u2_u6_n132 ) , .A3( u2_u2_u6_n145 ) );
  INV_X1 u2_u2_u6_U28 (.A( u2_u2_u6_n146 ) , .ZN( u2_u2_u6_n163 ) );
  AOI222_X1 u2_u2_u6_U29 (.ZN( u2_u2_u6_n114 ) , .A1( u2_u2_u6_n118 ) , .A2( u2_u2_u6_n126 ) , .B2( u2_u2_u6_n151 ) , .C2( u2_u2_u6_n159 ) , .C1( u2_u2_u6_n168 ) , .B1( u2_u2_u6_n169 ) );
  INV_X1 u2_u2_u6_U3 (.A( u2_u2_u6_n110 ) , .ZN( u2_u2_u6_n166 ) );
  NOR2_X1 u2_u2_u6_U30 (.A1( u2_u2_u6_n162 ) , .A2( u2_u2_u6_n165 ) , .ZN( u2_u2_u6_n98 ) );
  NAND2_X1 u2_u2_u6_U31 (.A1( u2_u2_u6_n144 ) , .ZN( u2_u2_u6_n151 ) , .A2( u2_u2_u6_n158 ) );
  NAND2_X1 u2_u2_u6_U32 (.ZN( u2_u2_u6_n132 ) , .A1( u2_u2_u6_n91 ) , .A2( u2_u2_u6_n97 ) );
  AOI22_X1 u2_u2_u6_U33 (.B2( u2_u2_u6_n110 ) , .B1( u2_u2_u6_n111 ) , .A1( u2_u2_u6_n112 ) , .ZN( u2_u2_u6_n115 ) , .A2( u2_u2_u6_n161 ) );
  NAND4_X1 u2_u2_u6_U34 (.A3( u2_u2_u6_n109 ) , .ZN( u2_u2_u6_n112 ) , .A4( u2_u2_u6_n132 ) , .A2( u2_u2_u6_n147 ) , .A1( u2_u2_u6_n166 ) );
  NOR2_X1 u2_u2_u6_U35 (.ZN( u2_u2_u6_n109 ) , .A1( u2_u2_u6_n170 ) , .A2( u2_u2_u6_n173 ) );
  NOR2_X1 u2_u2_u6_U36 (.A2( u2_u2_u6_n126 ) , .ZN( u2_u2_u6_n155 ) , .A1( u2_u2_u6_n160 ) );
  NAND2_X1 u2_u2_u6_U37 (.ZN( u2_u2_u6_n146 ) , .A2( u2_u2_u6_n94 ) , .A1( u2_u2_u6_n99 ) );
  AOI21_X1 u2_u2_u6_U38 (.A( u2_u2_u6_n144 ) , .B2( u2_u2_u6_n145 ) , .B1( u2_u2_u6_n146 ) , .ZN( u2_u2_u6_n150 ) );
  INV_X1 u2_u2_u6_U39 (.A( u2_u2_u6_n111 ) , .ZN( u2_u2_u6_n158 ) );
  INV_X1 u2_u2_u6_U4 (.A( u2_u2_u6_n142 ) , .ZN( u2_u2_u6_n174 ) );
  NAND2_X1 u2_u2_u6_U40 (.ZN( u2_u2_u6_n127 ) , .A1( u2_u2_u6_n91 ) , .A2( u2_u2_u6_n92 ) );
  NAND2_X1 u2_u2_u6_U41 (.ZN( u2_u2_u6_n129 ) , .A2( u2_u2_u6_n95 ) , .A1( u2_u2_u6_n96 ) );
  INV_X1 u2_u2_u6_U42 (.A( u2_u2_u6_n144 ) , .ZN( u2_u2_u6_n159 ) );
  NAND2_X1 u2_u2_u6_U43 (.ZN( u2_u2_u6_n145 ) , .A2( u2_u2_u6_n97 ) , .A1( u2_u2_u6_n98 ) );
  NAND2_X1 u2_u2_u6_U44 (.ZN( u2_u2_u6_n148 ) , .A2( u2_u2_u6_n92 ) , .A1( u2_u2_u6_n94 ) );
  NAND2_X1 u2_u2_u6_U45 (.ZN( u2_u2_u6_n108 ) , .A2( u2_u2_u6_n139 ) , .A1( u2_u2_u6_n144 ) );
  NAND2_X1 u2_u2_u6_U46 (.ZN( u2_u2_u6_n121 ) , .A2( u2_u2_u6_n95 ) , .A1( u2_u2_u6_n97 ) );
  NAND2_X1 u2_u2_u6_U47 (.ZN( u2_u2_u6_n107 ) , .A2( u2_u2_u6_n92 ) , .A1( u2_u2_u6_n95 ) );
  AND2_X1 u2_u2_u6_U48 (.ZN( u2_u2_u6_n118 ) , .A2( u2_u2_u6_n91 ) , .A1( u2_u2_u6_n99 ) );
  NAND2_X1 u2_u2_u6_U49 (.ZN( u2_u2_u6_n147 ) , .A2( u2_u2_u6_n98 ) , .A1( u2_u2_u6_n99 ) );
  NAND2_X1 u2_u2_u6_U5 (.A2( u2_u2_u6_n143 ) , .ZN( u2_u2_u6_n152 ) , .A1( u2_u2_u6_n166 ) );
  NAND2_X1 u2_u2_u6_U50 (.ZN( u2_u2_u6_n128 ) , .A1( u2_u2_u6_n94 ) , .A2( u2_u2_u6_n96 ) );
  AOI211_X1 u2_u2_u6_U51 (.B( u2_u2_u6_n134 ) , .A( u2_u2_u6_n135 ) , .C1( u2_u2_u6_n136 ) , .ZN( u2_u2_u6_n137 ) , .C2( u2_u2_u6_n151 ) );
  AOI21_X1 u2_u2_u6_U52 (.B2( u2_u2_u6_n132 ) , .B1( u2_u2_u6_n133 ) , .ZN( u2_u2_u6_n134 ) , .A( u2_u2_u6_n158 ) );
  AOI21_X1 u2_u2_u6_U53 (.B1( u2_u2_u6_n131 ) , .ZN( u2_u2_u6_n135 ) , .A( u2_u2_u6_n144 ) , .B2( u2_u2_u6_n146 ) );
  NAND4_X1 u2_u2_u6_U54 (.A4( u2_u2_u6_n127 ) , .A3( u2_u2_u6_n128 ) , .A2( u2_u2_u6_n129 ) , .A1( u2_u2_u6_n130 ) , .ZN( u2_u2_u6_n136 ) );
  NAND2_X1 u2_u2_u6_U55 (.ZN( u2_u2_u6_n119 ) , .A2( u2_u2_u6_n95 ) , .A1( u2_u2_u6_n99 ) );
  NAND2_X1 u2_u2_u6_U56 (.ZN( u2_u2_u6_n123 ) , .A2( u2_u2_u6_n91 ) , .A1( u2_u2_u6_n96 ) );
  NAND2_X1 u2_u2_u6_U57 (.ZN( u2_u2_u6_n100 ) , .A2( u2_u2_u6_n92 ) , .A1( u2_u2_u6_n98 ) );
  NAND2_X1 u2_u2_u6_U58 (.ZN( u2_u2_u6_n122 ) , .A1( u2_u2_u6_n94 ) , .A2( u2_u2_u6_n97 ) );
  INV_X1 u2_u2_u6_U59 (.A( u2_u2_u6_n139 ) , .ZN( u2_u2_u6_n160 ) );
  AOI22_X1 u2_u2_u6_U6 (.B2( u2_u2_u6_n101 ) , .A1( u2_u2_u6_n102 ) , .ZN( u2_u2_u6_n103 ) , .B1( u2_u2_u6_n160 ) , .A2( u2_u2_u6_n161 ) );
  NAND2_X1 u2_u2_u6_U60 (.ZN( u2_u2_u6_n113 ) , .A1( u2_u2_u6_n96 ) , .A2( u2_u2_u6_n98 ) );
  NOR2_X1 u2_u2_u6_U61 (.A2( u2_u2_X_40 ) , .A1( u2_u2_X_41 ) , .ZN( u2_u2_u6_n126 ) );
  NOR2_X1 u2_u2_u6_U62 (.A2( u2_u2_X_39 ) , .A1( u2_u2_X_42 ) , .ZN( u2_u2_u6_n92 ) );
  NOR2_X1 u2_u2_u6_U63 (.A2( u2_u2_X_39 ) , .A1( u2_u2_u6_n156 ) , .ZN( u2_u2_u6_n97 ) );
  NOR2_X1 u2_u2_u6_U64 (.A2( u2_u2_X_38 ) , .A1( u2_u2_u6_n165 ) , .ZN( u2_u2_u6_n95 ) );
  NOR2_X1 u2_u2_u6_U65 (.A2( u2_u2_X_41 ) , .ZN( u2_u2_u6_n111 ) , .A1( u2_u2_u6_n157 ) );
  NOR2_X1 u2_u2_u6_U66 (.A2( u2_u2_X_37 ) , .A1( u2_u2_u6_n162 ) , .ZN( u2_u2_u6_n94 ) );
  NOR2_X1 u2_u2_u6_U67 (.A2( u2_u2_X_37 ) , .A1( u2_u2_X_38 ) , .ZN( u2_u2_u6_n91 ) );
  NAND2_X1 u2_u2_u6_U68 (.A1( u2_u2_X_41 ) , .ZN( u2_u2_u6_n144 ) , .A2( u2_u2_u6_n157 ) );
  NAND2_X1 u2_u2_u6_U69 (.A2( u2_u2_X_40 ) , .A1( u2_u2_X_41 ) , .ZN( u2_u2_u6_n139 ) );
  NOR2_X1 u2_u2_u6_U7 (.A1( u2_u2_u6_n118 ) , .ZN( u2_u2_u6_n143 ) , .A2( u2_u2_u6_n168 ) );
  AND2_X1 u2_u2_u6_U70 (.A1( u2_u2_X_39 ) , .A2( u2_u2_u6_n156 ) , .ZN( u2_u2_u6_n96 ) );
  AND2_X1 u2_u2_u6_U71 (.A1( u2_u2_X_39 ) , .A2( u2_u2_X_42 ) , .ZN( u2_u2_u6_n99 ) );
  INV_X1 u2_u2_u6_U72 (.A( u2_u2_X_40 ) , .ZN( u2_u2_u6_n157 ) );
  INV_X1 u2_u2_u6_U73 (.A( u2_u2_X_37 ) , .ZN( u2_u2_u6_n165 ) );
  INV_X1 u2_u2_u6_U74 (.A( u2_u2_X_38 ) , .ZN( u2_u2_u6_n162 ) );
  INV_X1 u2_u2_u6_U75 (.A( u2_u2_X_42 ) , .ZN( u2_u2_u6_n156 ) );
  NAND4_X1 u2_u2_u6_U76 (.ZN( u2_out2_32 ) , .A4( u2_u2_u6_n103 ) , .A3( u2_u2_u6_n104 ) , .A2( u2_u2_u6_n105 ) , .A1( u2_u2_u6_n106 ) );
  AOI22_X1 u2_u2_u6_U77 (.ZN( u2_u2_u6_n105 ) , .A2( u2_u2_u6_n108 ) , .A1( u2_u2_u6_n118 ) , .B2( u2_u2_u6_n126 ) , .B1( u2_u2_u6_n171 ) );
  AOI22_X1 u2_u2_u6_U78 (.ZN( u2_u2_u6_n104 ) , .A1( u2_u2_u6_n111 ) , .B1( u2_u2_u6_n124 ) , .B2( u2_u2_u6_n151 ) , .A2( u2_u2_u6_n93 ) );
  NAND4_X1 u2_u2_u6_U79 (.ZN( u2_out2_12 ) , .A4( u2_u2_u6_n114 ) , .A3( u2_u2_u6_n115 ) , .A2( u2_u2_u6_n116 ) , .A1( u2_u2_u6_n117 ) );
  AOI21_X1 u2_u2_u6_U8 (.B1( u2_u2_u6_n107 ) , .B2( u2_u2_u6_n132 ) , .A( u2_u2_u6_n158 ) , .ZN( u2_u2_u6_n88 ) );
  OAI22_X1 u2_u2_u6_U80 (.B2( u2_u2_u6_n111 ) , .ZN( u2_u2_u6_n116 ) , .B1( u2_u2_u6_n126 ) , .A2( u2_u2_u6_n164 ) , .A1( u2_u2_u6_n167 ) );
  OAI21_X1 u2_u2_u6_U81 (.A( u2_u2_u6_n108 ) , .ZN( u2_u2_u6_n117 ) , .B2( u2_u2_u6_n141 ) , .B1( u2_u2_u6_n163 ) );
  OAI211_X1 u2_u2_u6_U82 (.ZN( u2_out2_7 ) , .B( u2_u2_u6_n153 ) , .C2( u2_u2_u6_n154 ) , .C1( u2_u2_u6_n155 ) , .A( u2_u2_u6_n174 ) );
  NOR3_X1 u2_u2_u6_U83 (.A1( u2_u2_u6_n141 ) , .ZN( u2_u2_u6_n154 ) , .A3( u2_u2_u6_n164 ) , .A2( u2_u2_u6_n171 ) );
  AOI211_X1 u2_u2_u6_U84 (.B( u2_u2_u6_n149 ) , .A( u2_u2_u6_n150 ) , .C2( u2_u2_u6_n151 ) , .C1( u2_u2_u6_n152 ) , .ZN( u2_u2_u6_n153 ) );
  OAI211_X1 u2_u2_u6_U85 (.ZN( u2_out2_22 ) , .B( u2_u2_u6_n137 ) , .A( u2_u2_u6_n138 ) , .C2( u2_u2_u6_n139 ) , .C1( u2_u2_u6_n140 ) );
  AOI22_X1 u2_u2_u6_U86 (.B1( u2_u2_u6_n124 ) , .A2( u2_u2_u6_n125 ) , .A1( u2_u2_u6_n126 ) , .ZN( u2_u2_u6_n138 ) , .B2( u2_u2_u6_n161 ) );
  AND4_X1 u2_u2_u6_U87 (.A3( u2_u2_u6_n119 ) , .A1( u2_u2_u6_n120 ) , .A4( u2_u2_u6_n129 ) , .ZN( u2_u2_u6_n140 ) , .A2( u2_u2_u6_n143 ) );
  NAND3_X1 u2_u2_u6_U88 (.A2( u2_u2_u6_n123 ) , .ZN( u2_u2_u6_n125 ) , .A1( u2_u2_u6_n130 ) , .A3( u2_u2_u6_n131 ) );
  NAND3_X1 u2_u2_u6_U89 (.A3( u2_u2_u6_n133 ) , .ZN( u2_u2_u6_n141 ) , .A1( u2_u2_u6_n145 ) , .A2( u2_u2_u6_n148 ) );
  AOI21_X1 u2_u2_u6_U9 (.B2( u2_u2_u6_n147 ) , .B1( u2_u2_u6_n148 ) , .ZN( u2_u2_u6_n149 ) , .A( u2_u2_u6_n158 ) );
  NAND3_X1 u2_u2_u6_U90 (.ZN( u2_u2_u6_n101 ) , .A3( u2_u2_u6_n107 ) , .A2( u2_u2_u6_n121 ) , .A1( u2_u2_u6_n127 ) );
  NAND3_X1 u2_u2_u6_U91 (.ZN( u2_u2_u6_n102 ) , .A3( u2_u2_u6_n130 ) , .A2( u2_u2_u6_n145 ) , .A1( u2_u2_u6_n166 ) );
  NAND3_X1 u2_u2_u6_U92 (.A3( u2_u2_u6_n113 ) , .A1( u2_u2_u6_n119 ) , .A2( u2_u2_u6_n123 ) , .ZN( u2_u2_u6_n93 ) );
  NAND3_X1 u2_u2_u6_U93 (.ZN( u2_u2_u6_n142 ) , .A2( u2_u2_u6_n172 ) , .A3( u2_u2_u6_n89 ) , .A1( u2_u2_u6_n90 ) );
  AND3_X1 u2_u2_u7_U10 (.A3( u2_u2_u7_n110 ) , .A2( u2_u2_u7_n127 ) , .A1( u2_u2_u7_n132 ) , .ZN( u2_u2_u7_n92 ) );
  OAI21_X1 u2_u2_u7_U11 (.A( u2_u2_u7_n161 ) , .B1( u2_u2_u7_n168 ) , .B2( u2_u2_u7_n173 ) , .ZN( u2_u2_u7_n91 ) );
  AOI211_X1 u2_u2_u7_U12 (.A( u2_u2_u7_n117 ) , .ZN( u2_u2_u7_n118 ) , .C2( u2_u2_u7_n126 ) , .C1( u2_u2_u7_n177 ) , .B( u2_u2_u7_n180 ) );
  OAI22_X1 u2_u2_u7_U13 (.B1( u2_u2_u7_n115 ) , .ZN( u2_u2_u7_n117 ) , .A2( u2_u2_u7_n133 ) , .A1( u2_u2_u7_n137 ) , .B2( u2_u2_u7_n162 ) );
  INV_X1 u2_u2_u7_U14 (.A( u2_u2_u7_n116 ) , .ZN( u2_u2_u7_n180 ) );
  NOR3_X1 u2_u2_u7_U15 (.ZN( u2_u2_u7_n115 ) , .A3( u2_u2_u7_n145 ) , .A2( u2_u2_u7_n168 ) , .A1( u2_u2_u7_n169 ) );
  OAI211_X1 u2_u2_u7_U16 (.B( u2_u2_u7_n122 ) , .A( u2_u2_u7_n123 ) , .C2( u2_u2_u7_n124 ) , .ZN( u2_u2_u7_n154 ) , .C1( u2_u2_u7_n162 ) );
  AOI222_X1 u2_u2_u7_U17 (.ZN( u2_u2_u7_n122 ) , .C2( u2_u2_u7_n126 ) , .C1( u2_u2_u7_n145 ) , .B1( u2_u2_u7_n161 ) , .A2( u2_u2_u7_n165 ) , .B2( u2_u2_u7_n170 ) , .A1( u2_u2_u7_n176 ) );
  INV_X1 u2_u2_u7_U18 (.A( u2_u2_u7_n133 ) , .ZN( u2_u2_u7_n176 ) );
  NOR3_X1 u2_u2_u7_U19 (.A2( u2_u2_u7_n134 ) , .A1( u2_u2_u7_n135 ) , .ZN( u2_u2_u7_n136 ) , .A3( u2_u2_u7_n171 ) );
  NOR2_X1 u2_u2_u7_U20 (.A1( u2_u2_u7_n130 ) , .A2( u2_u2_u7_n134 ) , .ZN( u2_u2_u7_n153 ) );
  INV_X1 u2_u2_u7_U21 (.A( u2_u2_u7_n101 ) , .ZN( u2_u2_u7_n165 ) );
  NOR2_X1 u2_u2_u7_U22 (.ZN( u2_u2_u7_n111 ) , .A2( u2_u2_u7_n134 ) , .A1( u2_u2_u7_n169 ) );
  AOI21_X1 u2_u2_u7_U23 (.ZN( u2_u2_u7_n104 ) , .B2( u2_u2_u7_n112 ) , .B1( u2_u2_u7_n127 ) , .A( u2_u2_u7_n164 ) );
  AOI21_X1 u2_u2_u7_U24 (.ZN( u2_u2_u7_n106 ) , .B1( u2_u2_u7_n133 ) , .B2( u2_u2_u7_n146 ) , .A( u2_u2_u7_n162 ) );
  AOI21_X1 u2_u2_u7_U25 (.A( u2_u2_u7_n101 ) , .ZN( u2_u2_u7_n107 ) , .B2( u2_u2_u7_n128 ) , .B1( u2_u2_u7_n175 ) );
  INV_X1 u2_u2_u7_U26 (.A( u2_u2_u7_n138 ) , .ZN( u2_u2_u7_n171 ) );
  INV_X1 u2_u2_u7_U27 (.A( u2_u2_u7_n131 ) , .ZN( u2_u2_u7_n177 ) );
  INV_X1 u2_u2_u7_U28 (.A( u2_u2_u7_n110 ) , .ZN( u2_u2_u7_n174 ) );
  NAND2_X1 u2_u2_u7_U29 (.A1( u2_u2_u7_n129 ) , .A2( u2_u2_u7_n132 ) , .ZN( u2_u2_u7_n149 ) );
  OAI21_X1 u2_u2_u7_U3 (.ZN( u2_u2_u7_n159 ) , .A( u2_u2_u7_n165 ) , .B2( u2_u2_u7_n171 ) , .B1( u2_u2_u7_n174 ) );
  NAND2_X1 u2_u2_u7_U30 (.A1( u2_u2_u7_n113 ) , .A2( u2_u2_u7_n124 ) , .ZN( u2_u2_u7_n130 ) );
  INV_X1 u2_u2_u7_U31 (.A( u2_u2_u7_n112 ) , .ZN( u2_u2_u7_n173 ) );
  INV_X1 u2_u2_u7_U32 (.A( u2_u2_u7_n128 ) , .ZN( u2_u2_u7_n168 ) );
  INV_X1 u2_u2_u7_U33 (.A( u2_u2_u7_n148 ) , .ZN( u2_u2_u7_n169 ) );
  INV_X1 u2_u2_u7_U34 (.A( u2_u2_u7_n127 ) , .ZN( u2_u2_u7_n179 ) );
  NOR2_X1 u2_u2_u7_U35 (.ZN( u2_u2_u7_n101 ) , .A2( u2_u2_u7_n150 ) , .A1( u2_u2_u7_n156 ) );
  AOI211_X1 u2_u2_u7_U36 (.B( u2_u2_u7_n154 ) , .A( u2_u2_u7_n155 ) , .C1( u2_u2_u7_n156 ) , .ZN( u2_u2_u7_n157 ) , .C2( u2_u2_u7_n172 ) );
  INV_X1 u2_u2_u7_U37 (.A( u2_u2_u7_n153 ) , .ZN( u2_u2_u7_n172 ) );
  AOI211_X1 u2_u2_u7_U38 (.B( u2_u2_u7_n139 ) , .A( u2_u2_u7_n140 ) , .C2( u2_u2_u7_n141 ) , .ZN( u2_u2_u7_n142 ) , .C1( u2_u2_u7_n156 ) );
  NAND4_X1 u2_u2_u7_U39 (.A3( u2_u2_u7_n127 ) , .A2( u2_u2_u7_n128 ) , .A1( u2_u2_u7_n129 ) , .ZN( u2_u2_u7_n141 ) , .A4( u2_u2_u7_n147 ) );
  INV_X1 u2_u2_u7_U4 (.A( u2_u2_u7_n111 ) , .ZN( u2_u2_u7_n170 ) );
  AOI21_X1 u2_u2_u7_U40 (.A( u2_u2_u7_n137 ) , .B1( u2_u2_u7_n138 ) , .ZN( u2_u2_u7_n139 ) , .B2( u2_u2_u7_n146 ) );
  OAI22_X1 u2_u2_u7_U41 (.B1( u2_u2_u7_n136 ) , .ZN( u2_u2_u7_n140 ) , .A1( u2_u2_u7_n153 ) , .B2( u2_u2_u7_n162 ) , .A2( u2_u2_u7_n164 ) );
  AOI21_X1 u2_u2_u7_U42 (.ZN( u2_u2_u7_n123 ) , .B1( u2_u2_u7_n165 ) , .B2( u2_u2_u7_n177 ) , .A( u2_u2_u7_n97 ) );
  AOI21_X1 u2_u2_u7_U43 (.B2( u2_u2_u7_n113 ) , .B1( u2_u2_u7_n124 ) , .A( u2_u2_u7_n125 ) , .ZN( u2_u2_u7_n97 ) );
  INV_X1 u2_u2_u7_U44 (.A( u2_u2_u7_n125 ) , .ZN( u2_u2_u7_n161 ) );
  INV_X1 u2_u2_u7_U45 (.A( u2_u2_u7_n152 ) , .ZN( u2_u2_u7_n162 ) );
  AOI22_X1 u2_u2_u7_U46 (.A2( u2_u2_u7_n114 ) , .ZN( u2_u2_u7_n119 ) , .B1( u2_u2_u7_n130 ) , .A1( u2_u2_u7_n156 ) , .B2( u2_u2_u7_n165 ) );
  NAND2_X1 u2_u2_u7_U47 (.A2( u2_u2_u7_n112 ) , .ZN( u2_u2_u7_n114 ) , .A1( u2_u2_u7_n175 ) );
  AND2_X1 u2_u2_u7_U48 (.ZN( u2_u2_u7_n145 ) , .A2( u2_u2_u7_n98 ) , .A1( u2_u2_u7_n99 ) );
  NOR2_X1 u2_u2_u7_U49 (.ZN( u2_u2_u7_n137 ) , .A1( u2_u2_u7_n150 ) , .A2( u2_u2_u7_n161 ) );
  INV_X1 u2_u2_u7_U5 (.A( u2_u2_u7_n149 ) , .ZN( u2_u2_u7_n175 ) );
  AOI21_X1 u2_u2_u7_U50 (.ZN( u2_u2_u7_n105 ) , .B2( u2_u2_u7_n110 ) , .A( u2_u2_u7_n125 ) , .B1( u2_u2_u7_n147 ) );
  NAND2_X1 u2_u2_u7_U51 (.ZN( u2_u2_u7_n146 ) , .A1( u2_u2_u7_n95 ) , .A2( u2_u2_u7_n98 ) );
  NAND2_X1 u2_u2_u7_U52 (.A2( u2_u2_u7_n103 ) , .ZN( u2_u2_u7_n147 ) , .A1( u2_u2_u7_n93 ) );
  NAND2_X1 u2_u2_u7_U53 (.A1( u2_u2_u7_n103 ) , .ZN( u2_u2_u7_n127 ) , .A2( u2_u2_u7_n99 ) );
  OR2_X1 u2_u2_u7_U54 (.ZN( u2_u2_u7_n126 ) , .A2( u2_u2_u7_n152 ) , .A1( u2_u2_u7_n156 ) );
  NAND2_X1 u2_u2_u7_U55 (.A2( u2_u2_u7_n102 ) , .A1( u2_u2_u7_n103 ) , .ZN( u2_u2_u7_n133 ) );
  NAND2_X1 u2_u2_u7_U56 (.ZN( u2_u2_u7_n112 ) , .A2( u2_u2_u7_n96 ) , .A1( u2_u2_u7_n99 ) );
  NAND2_X1 u2_u2_u7_U57 (.A2( u2_u2_u7_n102 ) , .ZN( u2_u2_u7_n128 ) , .A1( u2_u2_u7_n98 ) );
  NAND2_X1 u2_u2_u7_U58 (.A1( u2_u2_u7_n100 ) , .ZN( u2_u2_u7_n113 ) , .A2( u2_u2_u7_n93 ) );
  NAND2_X1 u2_u2_u7_U59 (.A2( u2_u2_u7_n102 ) , .ZN( u2_u2_u7_n124 ) , .A1( u2_u2_u7_n96 ) );
  INV_X1 u2_u2_u7_U6 (.A( u2_u2_u7_n154 ) , .ZN( u2_u2_u7_n178 ) );
  NAND2_X1 u2_u2_u7_U60 (.ZN( u2_u2_u7_n110 ) , .A1( u2_u2_u7_n95 ) , .A2( u2_u2_u7_n96 ) );
  INV_X1 u2_u2_u7_U61 (.A( u2_u2_u7_n150 ) , .ZN( u2_u2_u7_n164 ) );
  AND2_X1 u2_u2_u7_U62 (.ZN( u2_u2_u7_n134 ) , .A1( u2_u2_u7_n93 ) , .A2( u2_u2_u7_n98 ) );
  NAND2_X1 u2_u2_u7_U63 (.A1( u2_u2_u7_n100 ) , .A2( u2_u2_u7_n102 ) , .ZN( u2_u2_u7_n129 ) );
  NAND2_X1 u2_u2_u7_U64 (.A2( u2_u2_u7_n103 ) , .ZN( u2_u2_u7_n131 ) , .A1( u2_u2_u7_n95 ) );
  NAND2_X1 u2_u2_u7_U65 (.A1( u2_u2_u7_n100 ) , .ZN( u2_u2_u7_n138 ) , .A2( u2_u2_u7_n99 ) );
  NAND2_X1 u2_u2_u7_U66 (.ZN( u2_u2_u7_n132 ) , .A1( u2_u2_u7_n93 ) , .A2( u2_u2_u7_n96 ) );
  NAND2_X1 u2_u2_u7_U67 (.A1( u2_u2_u7_n100 ) , .ZN( u2_u2_u7_n148 ) , .A2( u2_u2_u7_n95 ) );
  NOR2_X1 u2_u2_u7_U68 (.A2( u2_u2_X_47 ) , .ZN( u2_u2_u7_n150 ) , .A1( u2_u2_u7_n163 ) );
  NOR2_X1 u2_u2_u7_U69 (.A2( u2_u2_X_43 ) , .A1( u2_u2_X_44 ) , .ZN( u2_u2_u7_n103 ) );
  AOI211_X1 u2_u2_u7_U7 (.ZN( u2_u2_u7_n116 ) , .A( u2_u2_u7_n155 ) , .C1( u2_u2_u7_n161 ) , .C2( u2_u2_u7_n171 ) , .B( u2_u2_u7_n94 ) );
  NOR2_X1 u2_u2_u7_U70 (.A2( u2_u2_X_48 ) , .A1( u2_u2_u7_n166 ) , .ZN( u2_u2_u7_n95 ) );
  NOR2_X1 u2_u2_u7_U71 (.A2( u2_u2_X_45 ) , .A1( u2_u2_X_48 ) , .ZN( u2_u2_u7_n99 ) );
  NOR2_X1 u2_u2_u7_U72 (.A2( u2_u2_X_44 ) , .A1( u2_u2_u7_n167 ) , .ZN( u2_u2_u7_n98 ) );
  NOR2_X1 u2_u2_u7_U73 (.A2( u2_u2_X_46 ) , .A1( u2_u2_X_47 ) , .ZN( u2_u2_u7_n152 ) );
  AND2_X1 u2_u2_u7_U74 (.A1( u2_u2_X_47 ) , .ZN( u2_u2_u7_n156 ) , .A2( u2_u2_u7_n163 ) );
  NAND2_X1 u2_u2_u7_U75 (.A2( u2_u2_X_46 ) , .A1( u2_u2_X_47 ) , .ZN( u2_u2_u7_n125 ) );
  AND2_X1 u2_u2_u7_U76 (.A2( u2_u2_X_45 ) , .A1( u2_u2_X_48 ) , .ZN( u2_u2_u7_n102 ) );
  AND2_X1 u2_u2_u7_U77 (.A2( u2_u2_X_43 ) , .A1( u2_u2_X_44 ) , .ZN( u2_u2_u7_n96 ) );
  AND2_X1 u2_u2_u7_U78 (.A1( u2_u2_X_44 ) , .ZN( u2_u2_u7_n100 ) , .A2( u2_u2_u7_n167 ) );
  AND2_X1 u2_u2_u7_U79 (.A1( u2_u2_X_48 ) , .A2( u2_u2_u7_n166 ) , .ZN( u2_u2_u7_n93 ) );
  OAI222_X1 u2_u2_u7_U8 (.C2( u2_u2_u7_n101 ) , .B2( u2_u2_u7_n111 ) , .A1( u2_u2_u7_n113 ) , .C1( u2_u2_u7_n146 ) , .A2( u2_u2_u7_n162 ) , .B1( u2_u2_u7_n164 ) , .ZN( u2_u2_u7_n94 ) );
  INV_X1 u2_u2_u7_U80 (.A( u2_u2_X_46 ) , .ZN( u2_u2_u7_n163 ) );
  INV_X1 u2_u2_u7_U81 (.A( u2_u2_X_43 ) , .ZN( u2_u2_u7_n167 ) );
  INV_X1 u2_u2_u7_U82 (.A( u2_u2_X_45 ) , .ZN( u2_u2_u7_n166 ) );
  NAND4_X1 u2_u2_u7_U83 (.ZN( u2_out2_5 ) , .A4( u2_u2_u7_n108 ) , .A3( u2_u2_u7_n109 ) , .A1( u2_u2_u7_n116 ) , .A2( u2_u2_u7_n123 ) );
  AOI22_X1 u2_u2_u7_U84 (.ZN( u2_u2_u7_n109 ) , .A2( u2_u2_u7_n126 ) , .B2( u2_u2_u7_n145 ) , .B1( u2_u2_u7_n156 ) , .A1( u2_u2_u7_n171 ) );
  NOR4_X1 u2_u2_u7_U85 (.A4( u2_u2_u7_n104 ) , .A3( u2_u2_u7_n105 ) , .A2( u2_u2_u7_n106 ) , .A1( u2_u2_u7_n107 ) , .ZN( u2_u2_u7_n108 ) );
  NAND4_X1 u2_u2_u7_U86 (.ZN( u2_out2_27 ) , .A4( u2_u2_u7_n118 ) , .A3( u2_u2_u7_n119 ) , .A2( u2_u2_u7_n120 ) , .A1( u2_u2_u7_n121 ) );
  OAI21_X1 u2_u2_u7_U87 (.ZN( u2_u2_u7_n121 ) , .B2( u2_u2_u7_n145 ) , .A( u2_u2_u7_n150 ) , .B1( u2_u2_u7_n174 ) );
  OAI21_X1 u2_u2_u7_U88 (.ZN( u2_u2_u7_n120 ) , .A( u2_u2_u7_n161 ) , .B2( u2_u2_u7_n170 ) , .B1( u2_u2_u7_n179 ) );
  NAND4_X1 u2_u2_u7_U89 (.ZN( u2_out2_21 ) , .A4( u2_u2_u7_n157 ) , .A3( u2_u2_u7_n158 ) , .A2( u2_u2_u7_n159 ) , .A1( u2_u2_u7_n160 ) );
  OAI221_X1 u2_u2_u7_U9 (.C1( u2_u2_u7_n101 ) , .C2( u2_u2_u7_n147 ) , .ZN( u2_u2_u7_n155 ) , .B2( u2_u2_u7_n162 ) , .A( u2_u2_u7_n91 ) , .B1( u2_u2_u7_n92 ) );
  OAI21_X1 u2_u2_u7_U90 (.B1( u2_u2_u7_n145 ) , .ZN( u2_u2_u7_n160 ) , .A( u2_u2_u7_n161 ) , .B2( u2_u2_u7_n177 ) );
  AOI22_X1 u2_u2_u7_U91 (.B2( u2_u2_u7_n149 ) , .B1( u2_u2_u7_n150 ) , .A2( u2_u2_u7_n151 ) , .A1( u2_u2_u7_n152 ) , .ZN( u2_u2_u7_n158 ) );
  NAND4_X1 u2_u2_u7_U92 (.ZN( u2_out2_15 ) , .A4( u2_u2_u7_n142 ) , .A3( u2_u2_u7_n143 ) , .A2( u2_u2_u7_n144 ) , .A1( u2_u2_u7_n178 ) );
  OR2_X1 u2_u2_u7_U93 (.A2( u2_u2_u7_n125 ) , .A1( u2_u2_u7_n129 ) , .ZN( u2_u2_u7_n144 ) );
  AOI22_X1 u2_u2_u7_U94 (.A2( u2_u2_u7_n126 ) , .ZN( u2_u2_u7_n143 ) , .B2( u2_u2_u7_n165 ) , .B1( u2_u2_u7_n173 ) , .A1( u2_u2_u7_n174 ) );
  NAND3_X1 u2_u2_u7_U95 (.A3( u2_u2_u7_n146 ) , .A2( u2_u2_u7_n147 ) , .A1( u2_u2_u7_n148 ) , .ZN( u2_u2_u7_n151 ) );
  NAND3_X1 u2_u2_u7_U96 (.A3( u2_u2_u7_n131 ) , .A2( u2_u2_u7_n132 ) , .A1( u2_u2_u7_n133 ) , .ZN( u2_u2_u7_n135 ) );
  XOR2_X1 u2_u3_U1 (.B( u2_K4_9 ) , .A( u2_R2_6 ) , .Z( u2_u3_X_9 ) );
  XOR2_X1 u2_u3_U16 (.B( u2_K4_3 ) , .A( u2_R2_2 ) , .Z( u2_u3_X_3 ) );
  XOR2_X1 u2_u3_U2 (.B( u2_K4_8 ) , .A( u2_R2_5 ) , .Z( u2_u3_X_8 ) );
  XOR2_X1 u2_u3_U20 (.B( u2_K4_36 ) , .A( u2_R2_25 ) , .Z( u2_u3_X_36 ) );
  XOR2_X1 u2_u3_U24 (.B( u2_K4_32 ) , .A( u2_R2_21 ) , .Z( u2_u3_X_32 ) );
  XOR2_X1 u2_u3_U25 (.B( u2_K4_31 ) , .A( u2_R2_20 ) , .Z( u2_u3_X_31 ) );
  XOR2_X1 u2_u3_U26 (.B( u2_K4_30 ) , .A( u2_R2_21 ) , .Z( u2_u3_X_30 ) );
  XOR2_X1 u2_u3_U27 (.B( u2_K4_2 ) , .A( u2_R2_1 ) , .Z( u2_u3_X_2 ) );
  XOR2_X1 u2_u3_U28 (.B( u2_K4_29 ) , .A( u2_R2_20 ) , .Z( u2_u3_X_29 ) );
  XOR2_X1 u2_u3_U29 (.B( u2_K4_28 ) , .A( u2_R2_19 ) , .Z( u2_u3_X_28 ) );
  XOR2_X1 u2_u3_U3 (.B( u2_K4_7 ) , .A( u2_R2_4 ) , .Z( u2_u3_X_7 ) );
  XOR2_X1 u2_u3_U31 (.B( u2_K4_26 ) , .A( u2_R2_17 ) , .Z( u2_u3_X_26 ) );
  XOR2_X1 u2_u3_U32 (.B( u2_K4_25 ) , .A( u2_R2_16 ) , .Z( u2_u3_X_25 ) );
  XOR2_X1 u2_u3_U33 (.B( u2_K4_24 ) , .A( u2_R2_17 ) , .Z( u2_u3_X_24 ) );
  XOR2_X1 u2_u3_U34 (.B( u2_K4_23 ) , .A( u2_R2_16 ) , .Z( u2_u3_X_23 ) );
  XOR2_X1 u2_u3_U37 (.B( u2_K4_20 ) , .A( u2_R2_13 ) , .Z( u2_u3_X_20 ) );
  XOR2_X1 u2_u3_U38 (.B( u2_K4_1 ) , .A( u2_R2_32 ) , .Z( u2_u3_X_1 ) );
  XOR2_X1 u2_u3_U39 (.B( u2_K4_19 ) , .A( u2_R2_12 ) , .Z( u2_u3_X_19 ) );
  XOR2_X1 u2_u3_U4 (.B( u2_K4_6 ) , .A( u2_R2_5 ) , .Z( u2_u3_X_6 ) );
  XOR2_X1 u2_u3_U40 (.B( u2_K4_18 ) , .A( u2_R2_13 ) , .Z( u2_u3_X_18 ) );
  XOR2_X1 u2_u3_U41 (.B( u2_K4_17 ) , .A( u2_R2_12 ) , .Z( u2_u3_X_17 ) );
  XOR2_X1 u2_u3_U42 (.B( u2_K4_16 ) , .A( u2_R2_11 ) , .Z( u2_u3_X_16 ) );
  XOR2_X1 u2_u3_U43 (.B( u2_K4_15 ) , .A( u2_R2_10 ) , .Z( u2_u3_X_15 ) );
  XOR2_X1 u2_u3_U44 (.B( u2_K4_14 ) , .A( u2_R2_9 ) , .Z( u2_u3_X_14 ) );
  XOR2_X1 u2_u3_U45 (.B( u2_K4_13 ) , .A( u2_R2_8 ) , .Z( u2_u3_X_13 ) );
  XOR2_X1 u2_u3_U46 (.B( u2_K4_12 ) , .A( u2_R2_9 ) , .Z( u2_u3_X_12 ) );
  XOR2_X1 u2_u3_U47 (.B( u2_K4_11 ) , .A( u2_R2_8 ) , .Z( u2_u3_X_11 ) );
  XOR2_X1 u2_u3_U48 (.B( u2_K4_10 ) , .A( u2_R2_7 ) , .Z( u2_u3_X_10 ) );
  XOR2_X1 u2_u3_U5 (.B( u2_K4_5 ) , .A( u2_R2_4 ) , .Z( u2_u3_X_5 ) );
  XOR2_X1 u2_u3_U6 (.B( u2_K4_4 ) , .A( u2_R2_3 ) , .Z( u2_u3_X_4 ) );
  XOR2_X1 u2_u3_U7 (.B( u2_K4_48 ) , .A( u2_R2_1 ) , .Z( u2_u3_X_48 ) );
  XOR2_X1 u2_u3_U8 (.B( u2_K4_47 ) , .A( u2_R2_32 ) , .Z( u2_u3_X_47 ) );
  AND3_X1 u2_u3_u0_U10 (.A2( u2_u3_u0_n112 ) , .ZN( u2_u3_u0_n127 ) , .A3( u2_u3_u0_n130 ) , .A1( u2_u3_u0_n148 ) );
  NAND2_X1 u2_u3_u0_U11 (.ZN( u2_u3_u0_n113 ) , .A1( u2_u3_u0_n139 ) , .A2( u2_u3_u0_n149 ) );
  AND2_X1 u2_u3_u0_U12 (.ZN( u2_u3_u0_n107 ) , .A1( u2_u3_u0_n130 ) , .A2( u2_u3_u0_n140 ) );
  AND2_X1 u2_u3_u0_U13 (.A2( u2_u3_u0_n129 ) , .A1( u2_u3_u0_n130 ) , .ZN( u2_u3_u0_n151 ) );
  AND2_X1 u2_u3_u0_U14 (.A1( u2_u3_u0_n108 ) , .A2( u2_u3_u0_n125 ) , .ZN( u2_u3_u0_n145 ) );
  INV_X1 u2_u3_u0_U15 (.A( u2_u3_u0_n143 ) , .ZN( u2_u3_u0_n173 ) );
  NOR2_X1 u2_u3_u0_U16 (.A2( u2_u3_u0_n136 ) , .ZN( u2_u3_u0_n147 ) , .A1( u2_u3_u0_n160 ) );
  INV_X1 u2_u3_u0_U17 (.ZN( u2_u3_u0_n172 ) , .A( u2_u3_u0_n88 ) );
  OAI222_X1 u2_u3_u0_U18 (.C1( u2_u3_u0_n108 ) , .A1( u2_u3_u0_n125 ) , .B2( u2_u3_u0_n128 ) , .B1( u2_u3_u0_n144 ) , .A2( u2_u3_u0_n158 ) , .C2( u2_u3_u0_n161 ) , .ZN( u2_u3_u0_n88 ) );
  AOI21_X1 u2_u3_u0_U19 (.B1( u2_u3_u0_n103 ) , .ZN( u2_u3_u0_n132 ) , .A( u2_u3_u0_n165 ) , .B2( u2_u3_u0_n93 ) );
  INV_X1 u2_u3_u0_U20 (.A( u2_u3_u0_n142 ) , .ZN( u2_u3_u0_n165 ) );
  OAI22_X1 u2_u3_u0_U21 (.B1( u2_u3_u0_n125 ) , .ZN( u2_u3_u0_n126 ) , .A1( u2_u3_u0_n138 ) , .A2( u2_u3_u0_n146 ) , .B2( u2_u3_u0_n147 ) );
  OAI22_X1 u2_u3_u0_U22 (.B1( u2_u3_u0_n131 ) , .A1( u2_u3_u0_n144 ) , .B2( u2_u3_u0_n147 ) , .A2( u2_u3_u0_n90 ) , .ZN( u2_u3_u0_n91 ) );
  AND3_X1 u2_u3_u0_U23 (.A3( u2_u3_u0_n121 ) , .A2( u2_u3_u0_n125 ) , .A1( u2_u3_u0_n148 ) , .ZN( u2_u3_u0_n90 ) );
  INV_X1 u2_u3_u0_U24 (.A( u2_u3_u0_n136 ) , .ZN( u2_u3_u0_n161 ) );
  AOI22_X1 u2_u3_u0_U25 (.B2( u2_u3_u0_n109 ) , .A2( u2_u3_u0_n110 ) , .ZN( u2_u3_u0_n111 ) , .B1( u2_u3_u0_n118 ) , .A1( u2_u3_u0_n160 ) );
  NAND2_X1 u2_u3_u0_U26 (.A2( u2_u3_u0_n103 ) , .ZN( u2_u3_u0_n140 ) , .A1( u2_u3_u0_n94 ) );
  INV_X1 u2_u3_u0_U27 (.A( u2_u3_u0_n118 ) , .ZN( u2_u3_u0_n158 ) );
  AOI21_X1 u2_u3_u0_U28 (.ZN( u2_u3_u0_n104 ) , .B1( u2_u3_u0_n107 ) , .B2( u2_u3_u0_n141 ) , .A( u2_u3_u0_n144 ) );
  AOI21_X1 u2_u3_u0_U29 (.B1( u2_u3_u0_n127 ) , .B2( u2_u3_u0_n129 ) , .A( u2_u3_u0_n138 ) , .ZN( u2_u3_u0_n96 ) );
  INV_X1 u2_u3_u0_U3 (.A( u2_u3_u0_n113 ) , .ZN( u2_u3_u0_n166 ) );
  NOR2_X1 u2_u3_u0_U30 (.A1( u2_u3_u0_n120 ) , .ZN( u2_u3_u0_n143 ) , .A2( u2_u3_u0_n167 ) );
  OAI221_X1 u2_u3_u0_U31 (.C1( u2_u3_u0_n112 ) , .ZN( u2_u3_u0_n120 ) , .B1( u2_u3_u0_n138 ) , .B2( u2_u3_u0_n141 ) , .C2( u2_u3_u0_n147 ) , .A( u2_u3_u0_n172 ) );
  AOI21_X1 u2_u3_u0_U32 (.ZN( u2_u3_u0_n116 ) , .B2( u2_u3_u0_n142 ) , .A( u2_u3_u0_n144 ) , .B1( u2_u3_u0_n166 ) );
  NAND2_X1 u2_u3_u0_U33 (.A1( u2_u3_u0_n101 ) , .A2( u2_u3_u0_n102 ) , .ZN( u2_u3_u0_n150 ) );
  INV_X1 u2_u3_u0_U34 (.A( u2_u3_u0_n138 ) , .ZN( u2_u3_u0_n160 ) );
  NAND2_X1 u2_u3_u0_U35 (.ZN( u2_u3_u0_n108 ) , .A1( u2_u3_u0_n92 ) , .A2( u2_u3_u0_n94 ) );
  NAND2_X1 u2_u3_u0_U36 (.A2( u2_u3_u0_n102 ) , .A1( u2_u3_u0_n103 ) , .ZN( u2_u3_u0_n149 ) );
  NAND2_X1 u2_u3_u0_U37 (.A1( u2_u3_u0_n101 ) , .ZN( u2_u3_u0_n130 ) , .A2( u2_u3_u0_n94 ) );
  NAND2_X1 u2_u3_u0_U38 (.A2( u2_u3_u0_n102 ) , .ZN( u2_u3_u0_n114 ) , .A1( u2_u3_u0_n92 ) );
  NAND2_X1 u2_u3_u0_U39 (.A2( u2_u3_u0_n101 ) , .ZN( u2_u3_u0_n121 ) , .A1( u2_u3_u0_n93 ) );
  AOI21_X1 u2_u3_u0_U4 (.B2( u2_u3_u0_n131 ) , .ZN( u2_u3_u0_n134 ) , .B1( u2_u3_u0_n151 ) , .A( u2_u3_u0_n158 ) );
  NAND2_X1 u2_u3_u0_U40 (.ZN( u2_u3_u0_n112 ) , .A2( u2_u3_u0_n92 ) , .A1( u2_u3_u0_n93 ) );
  OR3_X1 u2_u3_u0_U41 (.A3( u2_u3_u0_n152 ) , .A2( u2_u3_u0_n153 ) , .A1( u2_u3_u0_n154 ) , .ZN( u2_u3_u0_n155 ) );
  AOI21_X1 u2_u3_u0_U42 (.A( u2_u3_u0_n144 ) , .B2( u2_u3_u0_n145 ) , .B1( u2_u3_u0_n146 ) , .ZN( u2_u3_u0_n154 ) );
  AOI21_X1 u2_u3_u0_U43 (.B2( u2_u3_u0_n150 ) , .B1( u2_u3_u0_n151 ) , .ZN( u2_u3_u0_n152 ) , .A( u2_u3_u0_n158 ) );
  AOI21_X1 u2_u3_u0_U44 (.A( u2_u3_u0_n147 ) , .B2( u2_u3_u0_n148 ) , .B1( u2_u3_u0_n149 ) , .ZN( u2_u3_u0_n153 ) );
  INV_X1 u2_u3_u0_U45 (.ZN( u2_u3_u0_n171 ) , .A( u2_u3_u0_n99 ) );
  OAI211_X1 u2_u3_u0_U46 (.C2( u2_u3_u0_n140 ) , .C1( u2_u3_u0_n161 ) , .A( u2_u3_u0_n169 ) , .B( u2_u3_u0_n98 ) , .ZN( u2_u3_u0_n99 ) );
  AOI211_X1 u2_u3_u0_U47 (.C1( u2_u3_u0_n118 ) , .A( u2_u3_u0_n123 ) , .B( u2_u3_u0_n96 ) , .C2( u2_u3_u0_n97 ) , .ZN( u2_u3_u0_n98 ) );
  INV_X1 u2_u3_u0_U48 (.ZN( u2_u3_u0_n169 ) , .A( u2_u3_u0_n91 ) );
  NOR2_X1 u2_u3_u0_U49 (.A2( u2_u3_X_2 ) , .ZN( u2_u3_u0_n103 ) , .A1( u2_u3_u0_n164 ) );
  NOR2_X1 u2_u3_u0_U5 (.A1( u2_u3_u0_n108 ) , .ZN( u2_u3_u0_n123 ) , .A2( u2_u3_u0_n158 ) );
  NOR2_X1 u2_u3_u0_U50 (.A2( u2_u3_X_1 ) , .A1( u2_u3_X_2 ) , .ZN( u2_u3_u0_n92 ) );
  NOR2_X1 u2_u3_u0_U51 (.A2( u2_u3_X_4 ) , .A1( u2_u3_X_5 ) , .ZN( u2_u3_u0_n118 ) );
  NOR2_X1 u2_u3_u0_U52 (.A2( u2_u3_X_1 ) , .ZN( u2_u3_u0_n101 ) , .A1( u2_u3_u0_n163 ) );
  NAND2_X1 u2_u3_u0_U53 (.A2( u2_u3_X_4 ) , .A1( u2_u3_X_5 ) , .ZN( u2_u3_u0_n144 ) );
  NOR2_X1 u2_u3_u0_U54 (.A2( u2_u3_X_5 ) , .ZN( u2_u3_u0_n136 ) , .A1( u2_u3_u0_n159 ) );
  NAND2_X1 u2_u3_u0_U55 (.A1( u2_u3_X_5 ) , .ZN( u2_u3_u0_n138 ) , .A2( u2_u3_u0_n159 ) );
  NOR2_X1 u2_u3_u0_U56 (.A2( u2_u3_X_6 ) , .ZN( u2_u3_u0_n100 ) , .A1( u2_u3_u0_n162 ) );
  AND2_X1 u2_u3_u0_U57 (.A2( u2_u3_X_3 ) , .A1( u2_u3_X_6 ) , .ZN( u2_u3_u0_n102 ) );
  AND2_X1 u2_u3_u0_U58 (.A1( u2_u3_X_6 ) , .A2( u2_u3_u0_n162 ) , .ZN( u2_u3_u0_n93 ) );
  INV_X1 u2_u3_u0_U59 (.A( u2_u3_X_4 ) , .ZN( u2_u3_u0_n159 ) );
  OAI21_X1 u2_u3_u0_U6 (.B1( u2_u3_u0_n150 ) , .B2( u2_u3_u0_n158 ) , .A( u2_u3_u0_n172 ) , .ZN( u2_u3_u0_n89 ) );
  INV_X1 u2_u3_u0_U60 (.A( u2_u3_X_1 ) , .ZN( u2_u3_u0_n164 ) );
  INV_X1 u2_u3_u0_U61 (.A( u2_u3_X_2 ) , .ZN( u2_u3_u0_n163 ) );
  INV_X1 u2_u3_u0_U62 (.A( u2_u3_u0_n126 ) , .ZN( u2_u3_u0_n168 ) );
  AOI211_X1 u2_u3_u0_U63 (.B( u2_u3_u0_n133 ) , .A( u2_u3_u0_n134 ) , .C2( u2_u3_u0_n135 ) , .C1( u2_u3_u0_n136 ) , .ZN( u2_u3_u0_n137 ) );
  OR4_X1 u2_u3_u0_U64 (.ZN( u2_out3_17 ) , .A4( u2_u3_u0_n122 ) , .A2( u2_u3_u0_n123 ) , .A1( u2_u3_u0_n124 ) , .A3( u2_u3_u0_n170 ) );
  AOI21_X1 u2_u3_u0_U65 (.B2( u2_u3_u0_n107 ) , .ZN( u2_u3_u0_n124 ) , .B1( u2_u3_u0_n128 ) , .A( u2_u3_u0_n161 ) );
  INV_X1 u2_u3_u0_U66 (.A( u2_u3_u0_n111 ) , .ZN( u2_u3_u0_n170 ) );
  OR4_X1 u2_u3_u0_U67 (.ZN( u2_out3_31 ) , .A4( u2_u3_u0_n155 ) , .A2( u2_u3_u0_n156 ) , .A1( u2_u3_u0_n157 ) , .A3( u2_u3_u0_n173 ) );
  AOI21_X1 u2_u3_u0_U68 (.A( u2_u3_u0_n138 ) , .B2( u2_u3_u0_n139 ) , .B1( u2_u3_u0_n140 ) , .ZN( u2_u3_u0_n157 ) );
  AOI21_X1 u2_u3_u0_U69 (.B2( u2_u3_u0_n141 ) , .B1( u2_u3_u0_n142 ) , .ZN( u2_u3_u0_n156 ) , .A( u2_u3_u0_n161 ) );
  AOI21_X1 u2_u3_u0_U7 (.B1( u2_u3_u0_n114 ) , .ZN( u2_u3_u0_n115 ) , .B2( u2_u3_u0_n129 ) , .A( u2_u3_u0_n161 ) );
  INV_X1 u2_u3_u0_U70 (.ZN( u2_u3_u0_n174 ) , .A( u2_u3_u0_n89 ) );
  AOI211_X1 u2_u3_u0_U71 (.B( u2_u3_u0_n104 ) , .A( u2_u3_u0_n105 ) , .ZN( u2_u3_u0_n106 ) , .C2( u2_u3_u0_n113 ) , .C1( u2_u3_u0_n160 ) );
  AOI211_X1 u2_u3_u0_U72 (.B( u2_u3_u0_n115 ) , .A( u2_u3_u0_n116 ) , .C2( u2_u3_u0_n117 ) , .C1( u2_u3_u0_n118 ) , .ZN( u2_u3_u0_n119 ) );
  NAND2_X1 u2_u3_u0_U73 (.A2( u2_u3_u0_n100 ) , .ZN( u2_u3_u0_n131 ) , .A1( u2_u3_u0_n92 ) );
  NAND2_X1 u2_u3_u0_U74 (.A1( u2_u3_u0_n100 ) , .A2( u2_u3_u0_n103 ) , .ZN( u2_u3_u0_n125 ) );
  NAND2_X1 u2_u3_u0_U75 (.A2( u2_u3_u0_n100 ) , .A1( u2_u3_u0_n101 ) , .ZN( u2_u3_u0_n139 ) );
  NOR2_X1 u2_u3_u0_U76 (.A2( u2_u3_X_3 ) , .A1( u2_u3_X_6 ) , .ZN( u2_u3_u0_n94 ) );
  INV_X1 u2_u3_u0_U77 (.A( u2_u3_X_3 ) , .ZN( u2_u3_u0_n162 ) );
  NOR2_X1 u2_u3_u0_U78 (.A1( u2_u3_u0_n163 ) , .A2( u2_u3_u0_n164 ) , .ZN( u2_u3_u0_n95 ) );
  OAI221_X1 u2_u3_u0_U79 (.C1( u2_u3_u0_n121 ) , .ZN( u2_u3_u0_n122 ) , .B2( u2_u3_u0_n127 ) , .A( u2_u3_u0_n143 ) , .B1( u2_u3_u0_n144 ) , .C2( u2_u3_u0_n147 ) );
  AND2_X1 u2_u3_u0_U8 (.A1( u2_u3_u0_n114 ) , .A2( u2_u3_u0_n121 ) , .ZN( u2_u3_u0_n146 ) );
  AOI21_X1 u2_u3_u0_U80 (.B1( u2_u3_u0_n132 ) , .ZN( u2_u3_u0_n133 ) , .A( u2_u3_u0_n144 ) , .B2( u2_u3_u0_n166 ) );
  OAI22_X1 u2_u3_u0_U81 (.ZN( u2_u3_u0_n105 ) , .A2( u2_u3_u0_n132 ) , .B1( u2_u3_u0_n146 ) , .A1( u2_u3_u0_n147 ) , .B2( u2_u3_u0_n161 ) );
  NAND2_X1 u2_u3_u0_U82 (.ZN( u2_u3_u0_n110 ) , .A2( u2_u3_u0_n132 ) , .A1( u2_u3_u0_n145 ) );
  INV_X1 u2_u3_u0_U83 (.A( u2_u3_u0_n119 ) , .ZN( u2_u3_u0_n167 ) );
  NAND2_X1 u2_u3_u0_U84 (.ZN( u2_u3_u0_n148 ) , .A1( u2_u3_u0_n93 ) , .A2( u2_u3_u0_n95 ) );
  NAND2_X1 u2_u3_u0_U85 (.A1( u2_u3_u0_n100 ) , .ZN( u2_u3_u0_n129 ) , .A2( u2_u3_u0_n95 ) );
  NAND2_X1 u2_u3_u0_U86 (.A1( u2_u3_u0_n102 ) , .ZN( u2_u3_u0_n128 ) , .A2( u2_u3_u0_n95 ) );
  NAND2_X1 u2_u3_u0_U87 (.ZN( u2_u3_u0_n142 ) , .A1( u2_u3_u0_n94 ) , .A2( u2_u3_u0_n95 ) );
  NAND3_X1 u2_u3_u0_U88 (.ZN( u2_out3_23 ) , .A3( u2_u3_u0_n137 ) , .A1( u2_u3_u0_n168 ) , .A2( u2_u3_u0_n171 ) );
  NAND3_X1 u2_u3_u0_U89 (.A3( u2_u3_u0_n127 ) , .A2( u2_u3_u0_n128 ) , .ZN( u2_u3_u0_n135 ) , .A1( u2_u3_u0_n150 ) );
  AND2_X1 u2_u3_u0_U9 (.A1( u2_u3_u0_n131 ) , .ZN( u2_u3_u0_n141 ) , .A2( u2_u3_u0_n150 ) );
  NAND3_X1 u2_u3_u0_U90 (.ZN( u2_u3_u0_n117 ) , .A3( u2_u3_u0_n132 ) , .A2( u2_u3_u0_n139 ) , .A1( u2_u3_u0_n148 ) );
  NAND3_X1 u2_u3_u0_U91 (.ZN( u2_u3_u0_n109 ) , .A2( u2_u3_u0_n114 ) , .A3( u2_u3_u0_n140 ) , .A1( u2_u3_u0_n149 ) );
  NAND3_X1 u2_u3_u0_U92 (.ZN( u2_out3_9 ) , .A3( u2_u3_u0_n106 ) , .A2( u2_u3_u0_n171 ) , .A1( u2_u3_u0_n174 ) );
  NAND3_X1 u2_u3_u0_U93 (.A2( u2_u3_u0_n128 ) , .A1( u2_u3_u0_n132 ) , .A3( u2_u3_u0_n146 ) , .ZN( u2_u3_u0_n97 ) );
  NOR2_X1 u2_u3_u1_U10 (.A1( u2_u3_u1_n112 ) , .A2( u2_u3_u1_n116 ) , .ZN( u2_u3_u1_n118 ) );
  NAND3_X1 u2_u3_u1_U100 (.ZN( u2_u3_u1_n113 ) , .A1( u2_u3_u1_n120 ) , .A3( u2_u3_u1_n133 ) , .A2( u2_u3_u1_n155 ) );
  OAI21_X1 u2_u3_u1_U11 (.ZN( u2_u3_u1_n101 ) , .B1( u2_u3_u1_n141 ) , .A( u2_u3_u1_n146 ) , .B2( u2_u3_u1_n183 ) );
  AOI21_X1 u2_u3_u1_U12 (.B2( u2_u3_u1_n155 ) , .B1( u2_u3_u1_n156 ) , .ZN( u2_u3_u1_n157 ) , .A( u2_u3_u1_n174 ) );
  NAND2_X1 u2_u3_u1_U13 (.ZN( u2_u3_u1_n140 ) , .A2( u2_u3_u1_n150 ) , .A1( u2_u3_u1_n155 ) );
  NAND2_X1 u2_u3_u1_U14 (.A1( u2_u3_u1_n131 ) , .ZN( u2_u3_u1_n147 ) , .A2( u2_u3_u1_n153 ) );
  INV_X1 u2_u3_u1_U15 (.A( u2_u3_u1_n139 ) , .ZN( u2_u3_u1_n174 ) );
  OR4_X1 u2_u3_u1_U16 (.A4( u2_u3_u1_n106 ) , .A3( u2_u3_u1_n107 ) , .ZN( u2_u3_u1_n108 ) , .A1( u2_u3_u1_n117 ) , .A2( u2_u3_u1_n184 ) );
  AOI21_X1 u2_u3_u1_U17 (.ZN( u2_u3_u1_n106 ) , .A( u2_u3_u1_n112 ) , .B1( u2_u3_u1_n154 ) , .B2( u2_u3_u1_n156 ) );
  INV_X1 u2_u3_u1_U18 (.A( u2_u3_u1_n101 ) , .ZN( u2_u3_u1_n184 ) );
  AOI21_X1 u2_u3_u1_U19 (.ZN( u2_u3_u1_n107 ) , .B1( u2_u3_u1_n134 ) , .B2( u2_u3_u1_n149 ) , .A( u2_u3_u1_n174 ) );
  INV_X1 u2_u3_u1_U20 (.A( u2_u3_u1_n112 ) , .ZN( u2_u3_u1_n171 ) );
  NAND2_X1 u2_u3_u1_U21 (.ZN( u2_u3_u1_n141 ) , .A1( u2_u3_u1_n153 ) , .A2( u2_u3_u1_n156 ) );
  AND2_X1 u2_u3_u1_U22 (.A1( u2_u3_u1_n123 ) , .ZN( u2_u3_u1_n134 ) , .A2( u2_u3_u1_n161 ) );
  NAND2_X1 u2_u3_u1_U23 (.A2( u2_u3_u1_n115 ) , .A1( u2_u3_u1_n116 ) , .ZN( u2_u3_u1_n148 ) );
  NAND2_X1 u2_u3_u1_U24 (.A2( u2_u3_u1_n133 ) , .A1( u2_u3_u1_n135 ) , .ZN( u2_u3_u1_n159 ) );
  NAND2_X1 u2_u3_u1_U25 (.A2( u2_u3_u1_n115 ) , .A1( u2_u3_u1_n120 ) , .ZN( u2_u3_u1_n132 ) );
  INV_X1 u2_u3_u1_U26 (.A( u2_u3_u1_n154 ) , .ZN( u2_u3_u1_n178 ) );
  INV_X1 u2_u3_u1_U27 (.A( u2_u3_u1_n151 ) , .ZN( u2_u3_u1_n183 ) );
  AND2_X1 u2_u3_u1_U28 (.A1( u2_u3_u1_n129 ) , .A2( u2_u3_u1_n133 ) , .ZN( u2_u3_u1_n149 ) );
  INV_X1 u2_u3_u1_U29 (.A( u2_u3_u1_n131 ) , .ZN( u2_u3_u1_n180 ) );
  INV_X1 u2_u3_u1_U3 (.A( u2_u3_u1_n159 ) , .ZN( u2_u3_u1_n182 ) );
  AOI221_X1 u2_u3_u1_U30 (.B1( u2_u3_u1_n140 ) , .ZN( u2_u3_u1_n167 ) , .B2( u2_u3_u1_n172 ) , .C2( u2_u3_u1_n175 ) , .C1( u2_u3_u1_n178 ) , .A( u2_u3_u1_n188 ) );
  INV_X1 u2_u3_u1_U31 (.ZN( u2_u3_u1_n188 ) , .A( u2_u3_u1_n97 ) );
  AOI211_X1 u2_u3_u1_U32 (.A( u2_u3_u1_n118 ) , .C1( u2_u3_u1_n132 ) , .C2( u2_u3_u1_n139 ) , .B( u2_u3_u1_n96 ) , .ZN( u2_u3_u1_n97 ) );
  AOI21_X1 u2_u3_u1_U33 (.B2( u2_u3_u1_n121 ) , .B1( u2_u3_u1_n135 ) , .A( u2_u3_u1_n152 ) , .ZN( u2_u3_u1_n96 ) );
  OAI221_X1 u2_u3_u1_U34 (.A( u2_u3_u1_n119 ) , .C2( u2_u3_u1_n129 ) , .ZN( u2_u3_u1_n138 ) , .B2( u2_u3_u1_n152 ) , .C1( u2_u3_u1_n174 ) , .B1( u2_u3_u1_n187 ) );
  INV_X1 u2_u3_u1_U35 (.A( u2_u3_u1_n148 ) , .ZN( u2_u3_u1_n187 ) );
  AOI211_X1 u2_u3_u1_U36 (.B( u2_u3_u1_n117 ) , .A( u2_u3_u1_n118 ) , .ZN( u2_u3_u1_n119 ) , .C2( u2_u3_u1_n146 ) , .C1( u2_u3_u1_n159 ) );
  NOR2_X1 u2_u3_u1_U37 (.A1( u2_u3_u1_n168 ) , .A2( u2_u3_u1_n176 ) , .ZN( u2_u3_u1_n98 ) );
  NAND2_X1 u2_u3_u1_U38 (.A1( u2_u3_u1_n128 ) , .ZN( u2_u3_u1_n146 ) , .A2( u2_u3_u1_n160 ) );
  NAND2_X1 u2_u3_u1_U39 (.A2( u2_u3_u1_n112 ) , .ZN( u2_u3_u1_n139 ) , .A1( u2_u3_u1_n152 ) );
  AOI221_X1 u2_u3_u1_U4 (.A( u2_u3_u1_n138 ) , .C2( u2_u3_u1_n139 ) , .C1( u2_u3_u1_n140 ) , .B2( u2_u3_u1_n141 ) , .ZN( u2_u3_u1_n142 ) , .B1( u2_u3_u1_n175 ) );
  NAND2_X1 u2_u3_u1_U40 (.A1( u2_u3_u1_n105 ) , .ZN( u2_u3_u1_n156 ) , .A2( u2_u3_u1_n99 ) );
  NOR2_X1 u2_u3_u1_U41 (.ZN( u2_u3_u1_n117 ) , .A1( u2_u3_u1_n121 ) , .A2( u2_u3_u1_n160 ) );
  OAI21_X1 u2_u3_u1_U42 (.B2( u2_u3_u1_n123 ) , .ZN( u2_u3_u1_n145 ) , .B1( u2_u3_u1_n160 ) , .A( u2_u3_u1_n185 ) );
  INV_X1 u2_u3_u1_U43 (.A( u2_u3_u1_n122 ) , .ZN( u2_u3_u1_n185 ) );
  AOI21_X1 u2_u3_u1_U44 (.B2( u2_u3_u1_n120 ) , .B1( u2_u3_u1_n121 ) , .ZN( u2_u3_u1_n122 ) , .A( u2_u3_u1_n128 ) );
  AOI21_X1 u2_u3_u1_U45 (.A( u2_u3_u1_n128 ) , .B2( u2_u3_u1_n129 ) , .ZN( u2_u3_u1_n130 ) , .B1( u2_u3_u1_n150 ) );
  NAND2_X1 u2_u3_u1_U46 (.ZN( u2_u3_u1_n112 ) , .A1( u2_u3_u1_n169 ) , .A2( u2_u3_u1_n170 ) );
  NAND2_X1 u2_u3_u1_U47 (.ZN( u2_u3_u1_n129 ) , .A2( u2_u3_u1_n95 ) , .A1( u2_u3_u1_n98 ) );
  NAND2_X1 u2_u3_u1_U48 (.A1( u2_u3_u1_n102 ) , .ZN( u2_u3_u1_n154 ) , .A2( u2_u3_u1_n99 ) );
  NAND2_X1 u2_u3_u1_U49 (.A2( u2_u3_u1_n100 ) , .ZN( u2_u3_u1_n135 ) , .A1( u2_u3_u1_n99 ) );
  AOI211_X1 u2_u3_u1_U5 (.ZN( u2_u3_u1_n124 ) , .A( u2_u3_u1_n138 ) , .C2( u2_u3_u1_n139 ) , .B( u2_u3_u1_n145 ) , .C1( u2_u3_u1_n147 ) );
  AOI21_X1 u2_u3_u1_U50 (.A( u2_u3_u1_n152 ) , .B2( u2_u3_u1_n153 ) , .B1( u2_u3_u1_n154 ) , .ZN( u2_u3_u1_n158 ) );
  INV_X1 u2_u3_u1_U51 (.A( u2_u3_u1_n160 ) , .ZN( u2_u3_u1_n175 ) );
  NAND2_X1 u2_u3_u1_U52 (.A1( u2_u3_u1_n100 ) , .ZN( u2_u3_u1_n116 ) , .A2( u2_u3_u1_n95 ) );
  NAND2_X1 u2_u3_u1_U53 (.A1( u2_u3_u1_n102 ) , .ZN( u2_u3_u1_n131 ) , .A2( u2_u3_u1_n95 ) );
  NAND2_X1 u2_u3_u1_U54 (.A2( u2_u3_u1_n104 ) , .ZN( u2_u3_u1_n121 ) , .A1( u2_u3_u1_n98 ) );
  NAND2_X1 u2_u3_u1_U55 (.A1( u2_u3_u1_n103 ) , .ZN( u2_u3_u1_n153 ) , .A2( u2_u3_u1_n98 ) );
  NAND2_X1 u2_u3_u1_U56 (.A2( u2_u3_u1_n104 ) , .A1( u2_u3_u1_n105 ) , .ZN( u2_u3_u1_n133 ) );
  NAND2_X1 u2_u3_u1_U57 (.ZN( u2_u3_u1_n150 ) , .A2( u2_u3_u1_n98 ) , .A1( u2_u3_u1_n99 ) );
  NAND2_X1 u2_u3_u1_U58 (.A1( u2_u3_u1_n105 ) , .ZN( u2_u3_u1_n155 ) , .A2( u2_u3_u1_n95 ) );
  OAI21_X1 u2_u3_u1_U59 (.ZN( u2_u3_u1_n109 ) , .B1( u2_u3_u1_n129 ) , .B2( u2_u3_u1_n160 ) , .A( u2_u3_u1_n167 ) );
  AOI22_X1 u2_u3_u1_U6 (.B2( u2_u3_u1_n113 ) , .A2( u2_u3_u1_n114 ) , .ZN( u2_u3_u1_n125 ) , .A1( u2_u3_u1_n171 ) , .B1( u2_u3_u1_n173 ) );
  NAND2_X1 u2_u3_u1_U60 (.A2( u2_u3_u1_n100 ) , .A1( u2_u3_u1_n103 ) , .ZN( u2_u3_u1_n120 ) );
  NAND2_X1 u2_u3_u1_U61 (.A1( u2_u3_u1_n102 ) , .A2( u2_u3_u1_n104 ) , .ZN( u2_u3_u1_n115 ) );
  NAND2_X1 u2_u3_u1_U62 (.A2( u2_u3_u1_n100 ) , .A1( u2_u3_u1_n104 ) , .ZN( u2_u3_u1_n151 ) );
  NAND2_X1 u2_u3_u1_U63 (.A2( u2_u3_u1_n103 ) , .A1( u2_u3_u1_n105 ) , .ZN( u2_u3_u1_n161 ) );
  INV_X1 u2_u3_u1_U64 (.A( u2_u3_u1_n152 ) , .ZN( u2_u3_u1_n173 ) );
  INV_X1 u2_u3_u1_U65 (.A( u2_u3_u1_n128 ) , .ZN( u2_u3_u1_n172 ) );
  NAND2_X1 u2_u3_u1_U66 (.A2( u2_u3_u1_n102 ) , .A1( u2_u3_u1_n103 ) , .ZN( u2_u3_u1_n123 ) );
  AOI211_X1 u2_u3_u1_U67 (.B( u2_u3_u1_n162 ) , .A( u2_u3_u1_n163 ) , .C2( u2_u3_u1_n164 ) , .ZN( u2_u3_u1_n165 ) , .C1( u2_u3_u1_n171 ) );
  AOI21_X1 u2_u3_u1_U68 (.A( u2_u3_u1_n160 ) , .B2( u2_u3_u1_n161 ) , .ZN( u2_u3_u1_n162 ) , .B1( u2_u3_u1_n182 ) );
  OR2_X1 u2_u3_u1_U69 (.A2( u2_u3_u1_n157 ) , .A1( u2_u3_u1_n158 ) , .ZN( u2_u3_u1_n163 ) );
  NAND2_X1 u2_u3_u1_U7 (.ZN( u2_u3_u1_n114 ) , .A1( u2_u3_u1_n134 ) , .A2( u2_u3_u1_n156 ) );
  NOR2_X1 u2_u3_u1_U70 (.A2( u2_u3_X_7 ) , .A1( u2_u3_X_8 ) , .ZN( u2_u3_u1_n95 ) );
  NOR2_X1 u2_u3_u1_U71 (.A1( u2_u3_X_12 ) , .A2( u2_u3_X_9 ) , .ZN( u2_u3_u1_n100 ) );
  NOR2_X1 u2_u3_u1_U72 (.A2( u2_u3_X_8 ) , .A1( u2_u3_u1_n177 ) , .ZN( u2_u3_u1_n99 ) );
  NOR2_X1 u2_u3_u1_U73 (.A2( u2_u3_X_12 ) , .ZN( u2_u3_u1_n102 ) , .A1( u2_u3_u1_n176 ) );
  NOR2_X1 u2_u3_u1_U74 (.A2( u2_u3_X_9 ) , .ZN( u2_u3_u1_n105 ) , .A1( u2_u3_u1_n168 ) );
  NAND2_X1 u2_u3_u1_U75 (.A1( u2_u3_X_10 ) , .ZN( u2_u3_u1_n160 ) , .A2( u2_u3_u1_n169 ) );
  NAND2_X1 u2_u3_u1_U76 (.A2( u2_u3_X_10 ) , .A1( u2_u3_X_11 ) , .ZN( u2_u3_u1_n152 ) );
  NAND2_X1 u2_u3_u1_U77 (.A1( u2_u3_X_11 ) , .ZN( u2_u3_u1_n128 ) , .A2( u2_u3_u1_n170 ) );
  AND2_X1 u2_u3_u1_U78 (.A2( u2_u3_X_7 ) , .A1( u2_u3_X_8 ) , .ZN( u2_u3_u1_n104 ) );
  AND2_X1 u2_u3_u1_U79 (.A1( u2_u3_X_8 ) , .ZN( u2_u3_u1_n103 ) , .A2( u2_u3_u1_n177 ) );
  AOI22_X1 u2_u3_u1_U8 (.B2( u2_u3_u1_n136 ) , .A2( u2_u3_u1_n137 ) , .ZN( u2_u3_u1_n143 ) , .A1( u2_u3_u1_n171 ) , .B1( u2_u3_u1_n173 ) );
  INV_X1 u2_u3_u1_U80 (.A( u2_u3_X_10 ) , .ZN( u2_u3_u1_n170 ) );
  INV_X1 u2_u3_u1_U81 (.A( u2_u3_X_9 ) , .ZN( u2_u3_u1_n176 ) );
  INV_X1 u2_u3_u1_U82 (.A( u2_u3_X_11 ) , .ZN( u2_u3_u1_n169 ) );
  INV_X1 u2_u3_u1_U83 (.A( u2_u3_X_12 ) , .ZN( u2_u3_u1_n168 ) );
  INV_X1 u2_u3_u1_U84 (.A( u2_u3_X_7 ) , .ZN( u2_u3_u1_n177 ) );
  NAND4_X1 u2_u3_u1_U85 (.ZN( u2_out3_28 ) , .A4( u2_u3_u1_n124 ) , .A3( u2_u3_u1_n125 ) , .A2( u2_u3_u1_n126 ) , .A1( u2_u3_u1_n127 ) );
  OAI21_X1 u2_u3_u1_U86 (.ZN( u2_u3_u1_n127 ) , .B2( u2_u3_u1_n139 ) , .B1( u2_u3_u1_n175 ) , .A( u2_u3_u1_n183 ) );
  OAI21_X1 u2_u3_u1_U87 (.ZN( u2_u3_u1_n126 ) , .B2( u2_u3_u1_n140 ) , .A( u2_u3_u1_n146 ) , .B1( u2_u3_u1_n178 ) );
  NAND4_X1 u2_u3_u1_U88 (.ZN( u2_out3_18 ) , .A4( u2_u3_u1_n165 ) , .A3( u2_u3_u1_n166 ) , .A1( u2_u3_u1_n167 ) , .A2( u2_u3_u1_n186 ) );
  AOI22_X1 u2_u3_u1_U89 (.B2( u2_u3_u1_n146 ) , .B1( u2_u3_u1_n147 ) , .A2( u2_u3_u1_n148 ) , .ZN( u2_u3_u1_n166 ) , .A1( u2_u3_u1_n172 ) );
  INV_X1 u2_u3_u1_U9 (.A( u2_u3_u1_n147 ) , .ZN( u2_u3_u1_n181 ) );
  INV_X1 u2_u3_u1_U90 (.A( u2_u3_u1_n145 ) , .ZN( u2_u3_u1_n186 ) );
  NAND4_X1 u2_u3_u1_U91 (.ZN( u2_out3_2 ) , .A4( u2_u3_u1_n142 ) , .A3( u2_u3_u1_n143 ) , .A2( u2_u3_u1_n144 ) , .A1( u2_u3_u1_n179 ) );
  OAI21_X1 u2_u3_u1_U92 (.B2( u2_u3_u1_n132 ) , .ZN( u2_u3_u1_n144 ) , .A( u2_u3_u1_n146 ) , .B1( u2_u3_u1_n180 ) );
  INV_X1 u2_u3_u1_U93 (.A( u2_u3_u1_n130 ) , .ZN( u2_u3_u1_n179 ) );
  OR4_X1 u2_u3_u1_U94 (.ZN( u2_out3_13 ) , .A4( u2_u3_u1_n108 ) , .A3( u2_u3_u1_n109 ) , .A2( u2_u3_u1_n110 ) , .A1( u2_u3_u1_n111 ) );
  AOI21_X1 u2_u3_u1_U95 (.ZN( u2_u3_u1_n111 ) , .A( u2_u3_u1_n128 ) , .B2( u2_u3_u1_n131 ) , .B1( u2_u3_u1_n135 ) );
  AOI21_X1 u2_u3_u1_U96 (.ZN( u2_u3_u1_n110 ) , .A( u2_u3_u1_n116 ) , .B1( u2_u3_u1_n152 ) , .B2( u2_u3_u1_n160 ) );
  NAND3_X1 u2_u3_u1_U97 (.A3( u2_u3_u1_n149 ) , .A2( u2_u3_u1_n150 ) , .A1( u2_u3_u1_n151 ) , .ZN( u2_u3_u1_n164 ) );
  NAND3_X1 u2_u3_u1_U98 (.A3( u2_u3_u1_n134 ) , .A2( u2_u3_u1_n135 ) , .ZN( u2_u3_u1_n136 ) , .A1( u2_u3_u1_n151 ) );
  NAND3_X1 u2_u3_u1_U99 (.A1( u2_u3_u1_n133 ) , .ZN( u2_u3_u1_n137 ) , .A2( u2_u3_u1_n154 ) , .A3( u2_u3_u1_n181 ) );
  OAI22_X1 u2_u3_u2_U10 (.B1( u2_u3_u2_n151 ) , .A2( u2_u3_u2_n152 ) , .A1( u2_u3_u2_n153 ) , .ZN( u2_u3_u2_n160 ) , .B2( u2_u3_u2_n168 ) );
  NAND3_X1 u2_u3_u2_U100 (.A2( u2_u3_u2_n100 ) , .A1( u2_u3_u2_n104 ) , .A3( u2_u3_u2_n138 ) , .ZN( u2_u3_u2_n98 ) );
  NOR3_X1 u2_u3_u2_U11 (.A1( u2_u3_u2_n150 ) , .ZN( u2_u3_u2_n151 ) , .A3( u2_u3_u2_n175 ) , .A2( u2_u3_u2_n188 ) );
  AOI21_X1 u2_u3_u2_U12 (.B2( u2_u3_u2_n123 ) , .ZN( u2_u3_u2_n125 ) , .A( u2_u3_u2_n171 ) , .B1( u2_u3_u2_n184 ) );
  INV_X1 u2_u3_u2_U13 (.A( u2_u3_u2_n150 ) , .ZN( u2_u3_u2_n184 ) );
  AOI21_X1 u2_u3_u2_U14 (.ZN( u2_u3_u2_n144 ) , .B2( u2_u3_u2_n155 ) , .A( u2_u3_u2_n172 ) , .B1( u2_u3_u2_n185 ) );
  AOI21_X1 u2_u3_u2_U15 (.B2( u2_u3_u2_n143 ) , .ZN( u2_u3_u2_n145 ) , .B1( u2_u3_u2_n152 ) , .A( u2_u3_u2_n171 ) );
  INV_X1 u2_u3_u2_U16 (.A( u2_u3_u2_n156 ) , .ZN( u2_u3_u2_n171 ) );
  INV_X1 u2_u3_u2_U17 (.A( u2_u3_u2_n120 ) , .ZN( u2_u3_u2_n188 ) );
  NAND2_X1 u2_u3_u2_U18 (.A2( u2_u3_u2_n122 ) , .ZN( u2_u3_u2_n150 ) , .A1( u2_u3_u2_n152 ) );
  INV_X1 u2_u3_u2_U19 (.A( u2_u3_u2_n153 ) , .ZN( u2_u3_u2_n170 ) );
  INV_X1 u2_u3_u2_U20 (.A( u2_u3_u2_n137 ) , .ZN( u2_u3_u2_n173 ) );
  NAND2_X1 u2_u3_u2_U21 (.A1( u2_u3_u2_n132 ) , .A2( u2_u3_u2_n139 ) , .ZN( u2_u3_u2_n157 ) );
  INV_X1 u2_u3_u2_U22 (.A( u2_u3_u2_n113 ) , .ZN( u2_u3_u2_n178 ) );
  INV_X1 u2_u3_u2_U23 (.A( u2_u3_u2_n139 ) , .ZN( u2_u3_u2_n175 ) );
  INV_X1 u2_u3_u2_U24 (.A( u2_u3_u2_n155 ) , .ZN( u2_u3_u2_n181 ) );
  INV_X1 u2_u3_u2_U25 (.A( u2_u3_u2_n119 ) , .ZN( u2_u3_u2_n177 ) );
  INV_X1 u2_u3_u2_U26 (.A( u2_u3_u2_n116 ) , .ZN( u2_u3_u2_n180 ) );
  INV_X1 u2_u3_u2_U27 (.A( u2_u3_u2_n131 ) , .ZN( u2_u3_u2_n179 ) );
  INV_X1 u2_u3_u2_U28 (.A( u2_u3_u2_n154 ) , .ZN( u2_u3_u2_n176 ) );
  NAND2_X1 u2_u3_u2_U29 (.A2( u2_u3_u2_n116 ) , .A1( u2_u3_u2_n117 ) , .ZN( u2_u3_u2_n118 ) );
  NOR2_X1 u2_u3_u2_U3 (.ZN( u2_u3_u2_n121 ) , .A2( u2_u3_u2_n177 ) , .A1( u2_u3_u2_n180 ) );
  INV_X1 u2_u3_u2_U30 (.A( u2_u3_u2_n132 ) , .ZN( u2_u3_u2_n182 ) );
  INV_X1 u2_u3_u2_U31 (.A( u2_u3_u2_n158 ) , .ZN( u2_u3_u2_n183 ) );
  OAI21_X1 u2_u3_u2_U32 (.A( u2_u3_u2_n156 ) , .B1( u2_u3_u2_n157 ) , .ZN( u2_u3_u2_n158 ) , .B2( u2_u3_u2_n179 ) );
  NOR2_X1 u2_u3_u2_U33 (.ZN( u2_u3_u2_n156 ) , .A1( u2_u3_u2_n166 ) , .A2( u2_u3_u2_n169 ) );
  NOR2_X1 u2_u3_u2_U34 (.A2( u2_u3_u2_n114 ) , .ZN( u2_u3_u2_n137 ) , .A1( u2_u3_u2_n140 ) );
  NOR2_X1 u2_u3_u2_U35 (.A2( u2_u3_u2_n138 ) , .ZN( u2_u3_u2_n153 ) , .A1( u2_u3_u2_n156 ) );
  AOI211_X1 u2_u3_u2_U36 (.ZN( u2_u3_u2_n130 ) , .C1( u2_u3_u2_n138 ) , .C2( u2_u3_u2_n179 ) , .B( u2_u3_u2_n96 ) , .A( u2_u3_u2_n97 ) );
  OAI22_X1 u2_u3_u2_U37 (.B1( u2_u3_u2_n133 ) , .A2( u2_u3_u2_n137 ) , .A1( u2_u3_u2_n152 ) , .B2( u2_u3_u2_n168 ) , .ZN( u2_u3_u2_n97 ) );
  OAI221_X1 u2_u3_u2_U38 (.B1( u2_u3_u2_n113 ) , .C1( u2_u3_u2_n132 ) , .A( u2_u3_u2_n149 ) , .B2( u2_u3_u2_n171 ) , .C2( u2_u3_u2_n172 ) , .ZN( u2_u3_u2_n96 ) );
  OAI221_X1 u2_u3_u2_U39 (.A( u2_u3_u2_n115 ) , .C2( u2_u3_u2_n123 ) , .B2( u2_u3_u2_n143 ) , .B1( u2_u3_u2_n153 ) , .ZN( u2_u3_u2_n163 ) , .C1( u2_u3_u2_n168 ) );
  INV_X1 u2_u3_u2_U4 (.A( u2_u3_u2_n134 ) , .ZN( u2_u3_u2_n185 ) );
  OAI21_X1 u2_u3_u2_U40 (.A( u2_u3_u2_n114 ) , .ZN( u2_u3_u2_n115 ) , .B1( u2_u3_u2_n176 ) , .B2( u2_u3_u2_n178 ) );
  OAI221_X1 u2_u3_u2_U41 (.A( u2_u3_u2_n135 ) , .B2( u2_u3_u2_n136 ) , .B1( u2_u3_u2_n137 ) , .ZN( u2_u3_u2_n162 ) , .C2( u2_u3_u2_n167 ) , .C1( u2_u3_u2_n185 ) );
  AND3_X1 u2_u3_u2_U42 (.A3( u2_u3_u2_n131 ) , .A2( u2_u3_u2_n132 ) , .A1( u2_u3_u2_n133 ) , .ZN( u2_u3_u2_n136 ) );
  AOI22_X1 u2_u3_u2_U43 (.ZN( u2_u3_u2_n135 ) , .B1( u2_u3_u2_n140 ) , .A1( u2_u3_u2_n156 ) , .B2( u2_u3_u2_n180 ) , .A2( u2_u3_u2_n188 ) );
  AOI21_X1 u2_u3_u2_U44 (.ZN( u2_u3_u2_n149 ) , .B1( u2_u3_u2_n173 ) , .B2( u2_u3_u2_n188 ) , .A( u2_u3_u2_n95 ) );
  AND3_X1 u2_u3_u2_U45 (.A2( u2_u3_u2_n100 ) , .A1( u2_u3_u2_n104 ) , .A3( u2_u3_u2_n156 ) , .ZN( u2_u3_u2_n95 ) );
  OAI21_X1 u2_u3_u2_U46 (.A( u2_u3_u2_n141 ) , .B2( u2_u3_u2_n142 ) , .ZN( u2_u3_u2_n146 ) , .B1( u2_u3_u2_n153 ) );
  OAI21_X1 u2_u3_u2_U47 (.A( u2_u3_u2_n140 ) , .ZN( u2_u3_u2_n141 ) , .B1( u2_u3_u2_n176 ) , .B2( u2_u3_u2_n177 ) );
  NOR3_X1 u2_u3_u2_U48 (.ZN( u2_u3_u2_n142 ) , .A3( u2_u3_u2_n175 ) , .A2( u2_u3_u2_n178 ) , .A1( u2_u3_u2_n181 ) );
  OAI21_X1 u2_u3_u2_U49 (.A( u2_u3_u2_n101 ) , .B2( u2_u3_u2_n121 ) , .B1( u2_u3_u2_n153 ) , .ZN( u2_u3_u2_n164 ) );
  NOR4_X1 u2_u3_u2_U5 (.A4( u2_u3_u2_n124 ) , .A3( u2_u3_u2_n125 ) , .A2( u2_u3_u2_n126 ) , .A1( u2_u3_u2_n127 ) , .ZN( u2_u3_u2_n128 ) );
  NAND2_X1 u2_u3_u2_U50 (.A2( u2_u3_u2_n100 ) , .A1( u2_u3_u2_n107 ) , .ZN( u2_u3_u2_n155 ) );
  NAND2_X1 u2_u3_u2_U51 (.A2( u2_u3_u2_n105 ) , .A1( u2_u3_u2_n108 ) , .ZN( u2_u3_u2_n143 ) );
  NAND2_X1 u2_u3_u2_U52 (.A1( u2_u3_u2_n104 ) , .A2( u2_u3_u2_n106 ) , .ZN( u2_u3_u2_n152 ) );
  NAND2_X1 u2_u3_u2_U53 (.A1( u2_u3_u2_n100 ) , .A2( u2_u3_u2_n105 ) , .ZN( u2_u3_u2_n132 ) );
  INV_X1 u2_u3_u2_U54 (.A( u2_u3_u2_n140 ) , .ZN( u2_u3_u2_n168 ) );
  INV_X1 u2_u3_u2_U55 (.A( u2_u3_u2_n138 ) , .ZN( u2_u3_u2_n167 ) );
  INV_X1 u2_u3_u2_U56 (.ZN( u2_u3_u2_n187 ) , .A( u2_u3_u2_n99 ) );
  OAI21_X1 u2_u3_u2_U57 (.B1( u2_u3_u2_n137 ) , .B2( u2_u3_u2_n143 ) , .A( u2_u3_u2_n98 ) , .ZN( u2_u3_u2_n99 ) );
  NAND2_X1 u2_u3_u2_U58 (.A1( u2_u3_u2_n102 ) , .A2( u2_u3_u2_n106 ) , .ZN( u2_u3_u2_n113 ) );
  NAND2_X1 u2_u3_u2_U59 (.A1( u2_u3_u2_n106 ) , .A2( u2_u3_u2_n107 ) , .ZN( u2_u3_u2_n131 ) );
  AOI21_X1 u2_u3_u2_U6 (.B2( u2_u3_u2_n119 ) , .ZN( u2_u3_u2_n127 ) , .A( u2_u3_u2_n137 ) , .B1( u2_u3_u2_n155 ) );
  NAND2_X1 u2_u3_u2_U60 (.A1( u2_u3_u2_n103 ) , .A2( u2_u3_u2_n107 ) , .ZN( u2_u3_u2_n139 ) );
  NAND2_X1 u2_u3_u2_U61 (.A1( u2_u3_u2_n103 ) , .A2( u2_u3_u2_n105 ) , .ZN( u2_u3_u2_n133 ) );
  NAND2_X1 u2_u3_u2_U62 (.A1( u2_u3_u2_n102 ) , .A2( u2_u3_u2_n103 ) , .ZN( u2_u3_u2_n154 ) );
  NAND2_X1 u2_u3_u2_U63 (.A2( u2_u3_u2_n103 ) , .A1( u2_u3_u2_n104 ) , .ZN( u2_u3_u2_n119 ) );
  NAND2_X1 u2_u3_u2_U64 (.A2( u2_u3_u2_n107 ) , .A1( u2_u3_u2_n108 ) , .ZN( u2_u3_u2_n123 ) );
  NAND2_X1 u2_u3_u2_U65 (.A1( u2_u3_u2_n104 ) , .A2( u2_u3_u2_n108 ) , .ZN( u2_u3_u2_n122 ) );
  INV_X1 u2_u3_u2_U66 (.A( u2_u3_u2_n114 ) , .ZN( u2_u3_u2_n172 ) );
  NAND2_X1 u2_u3_u2_U67 (.A2( u2_u3_u2_n100 ) , .A1( u2_u3_u2_n102 ) , .ZN( u2_u3_u2_n116 ) );
  NAND2_X1 u2_u3_u2_U68 (.A1( u2_u3_u2_n102 ) , .A2( u2_u3_u2_n108 ) , .ZN( u2_u3_u2_n120 ) );
  NAND2_X1 u2_u3_u2_U69 (.A2( u2_u3_u2_n105 ) , .A1( u2_u3_u2_n106 ) , .ZN( u2_u3_u2_n117 ) );
  AOI21_X1 u2_u3_u2_U7 (.ZN( u2_u3_u2_n124 ) , .B1( u2_u3_u2_n131 ) , .B2( u2_u3_u2_n143 ) , .A( u2_u3_u2_n172 ) );
  NOR2_X1 u2_u3_u2_U70 (.A2( u2_u3_X_16 ) , .ZN( u2_u3_u2_n140 ) , .A1( u2_u3_u2_n166 ) );
  NOR2_X1 u2_u3_u2_U71 (.A2( u2_u3_X_13 ) , .A1( u2_u3_X_14 ) , .ZN( u2_u3_u2_n100 ) );
  NOR2_X1 u2_u3_u2_U72 (.A2( u2_u3_X_16 ) , .A1( u2_u3_X_17 ) , .ZN( u2_u3_u2_n138 ) );
  NOR2_X1 u2_u3_u2_U73 (.A2( u2_u3_X_15 ) , .A1( u2_u3_X_18 ) , .ZN( u2_u3_u2_n104 ) );
  NOR2_X1 u2_u3_u2_U74 (.A2( u2_u3_X_14 ) , .ZN( u2_u3_u2_n103 ) , .A1( u2_u3_u2_n174 ) );
  NOR2_X1 u2_u3_u2_U75 (.A2( u2_u3_X_15 ) , .ZN( u2_u3_u2_n102 ) , .A1( u2_u3_u2_n165 ) );
  NOR2_X1 u2_u3_u2_U76 (.A2( u2_u3_X_17 ) , .ZN( u2_u3_u2_n114 ) , .A1( u2_u3_u2_n169 ) );
  AND2_X1 u2_u3_u2_U77 (.A1( u2_u3_X_15 ) , .ZN( u2_u3_u2_n105 ) , .A2( u2_u3_u2_n165 ) );
  AND2_X1 u2_u3_u2_U78 (.A2( u2_u3_X_15 ) , .A1( u2_u3_X_18 ) , .ZN( u2_u3_u2_n107 ) );
  AND2_X1 u2_u3_u2_U79 (.A1( u2_u3_X_14 ) , .ZN( u2_u3_u2_n106 ) , .A2( u2_u3_u2_n174 ) );
  AOI21_X1 u2_u3_u2_U8 (.B2( u2_u3_u2_n120 ) , .B1( u2_u3_u2_n121 ) , .ZN( u2_u3_u2_n126 ) , .A( u2_u3_u2_n167 ) );
  AND2_X1 u2_u3_u2_U80 (.A1( u2_u3_X_13 ) , .A2( u2_u3_X_14 ) , .ZN( u2_u3_u2_n108 ) );
  INV_X1 u2_u3_u2_U81 (.A( u2_u3_X_16 ) , .ZN( u2_u3_u2_n169 ) );
  INV_X1 u2_u3_u2_U82 (.A( u2_u3_X_17 ) , .ZN( u2_u3_u2_n166 ) );
  INV_X1 u2_u3_u2_U83 (.A( u2_u3_X_13 ) , .ZN( u2_u3_u2_n174 ) );
  INV_X1 u2_u3_u2_U84 (.A( u2_u3_X_18 ) , .ZN( u2_u3_u2_n165 ) );
  NAND4_X1 u2_u3_u2_U85 (.ZN( u2_out3_24 ) , .A4( u2_u3_u2_n111 ) , .A3( u2_u3_u2_n112 ) , .A1( u2_u3_u2_n130 ) , .A2( u2_u3_u2_n187 ) );
  AOI221_X1 u2_u3_u2_U86 (.A( u2_u3_u2_n109 ) , .B1( u2_u3_u2_n110 ) , .ZN( u2_u3_u2_n111 ) , .C1( u2_u3_u2_n134 ) , .C2( u2_u3_u2_n170 ) , .B2( u2_u3_u2_n173 ) );
  AOI21_X1 u2_u3_u2_U87 (.ZN( u2_u3_u2_n112 ) , .B2( u2_u3_u2_n156 ) , .A( u2_u3_u2_n164 ) , .B1( u2_u3_u2_n181 ) );
  NAND4_X1 u2_u3_u2_U88 (.ZN( u2_out3_16 ) , .A4( u2_u3_u2_n128 ) , .A3( u2_u3_u2_n129 ) , .A1( u2_u3_u2_n130 ) , .A2( u2_u3_u2_n186 ) );
  AOI22_X1 u2_u3_u2_U89 (.A2( u2_u3_u2_n118 ) , .ZN( u2_u3_u2_n129 ) , .A1( u2_u3_u2_n140 ) , .B1( u2_u3_u2_n157 ) , .B2( u2_u3_u2_n170 ) );
  OAI22_X1 u2_u3_u2_U9 (.ZN( u2_u3_u2_n109 ) , .A2( u2_u3_u2_n113 ) , .B2( u2_u3_u2_n133 ) , .B1( u2_u3_u2_n167 ) , .A1( u2_u3_u2_n168 ) );
  INV_X1 u2_u3_u2_U90 (.A( u2_u3_u2_n163 ) , .ZN( u2_u3_u2_n186 ) );
  NAND4_X1 u2_u3_u2_U91 (.ZN( u2_out3_30 ) , .A4( u2_u3_u2_n147 ) , .A3( u2_u3_u2_n148 ) , .A2( u2_u3_u2_n149 ) , .A1( u2_u3_u2_n187 ) );
  AOI21_X1 u2_u3_u2_U92 (.B2( u2_u3_u2_n138 ) , .ZN( u2_u3_u2_n148 ) , .A( u2_u3_u2_n162 ) , .B1( u2_u3_u2_n182 ) );
  NOR3_X1 u2_u3_u2_U93 (.A3( u2_u3_u2_n144 ) , .A2( u2_u3_u2_n145 ) , .A1( u2_u3_u2_n146 ) , .ZN( u2_u3_u2_n147 ) );
  OR4_X1 u2_u3_u2_U94 (.ZN( u2_out3_6 ) , .A4( u2_u3_u2_n161 ) , .A3( u2_u3_u2_n162 ) , .A2( u2_u3_u2_n163 ) , .A1( u2_u3_u2_n164 ) );
  OR3_X1 u2_u3_u2_U95 (.A2( u2_u3_u2_n159 ) , .A1( u2_u3_u2_n160 ) , .ZN( u2_u3_u2_n161 ) , .A3( u2_u3_u2_n183 ) );
  AOI21_X1 u2_u3_u2_U96 (.B2( u2_u3_u2_n154 ) , .B1( u2_u3_u2_n155 ) , .ZN( u2_u3_u2_n159 ) , .A( u2_u3_u2_n167 ) );
  NAND3_X1 u2_u3_u2_U97 (.A2( u2_u3_u2_n117 ) , .A1( u2_u3_u2_n122 ) , .A3( u2_u3_u2_n123 ) , .ZN( u2_u3_u2_n134 ) );
  NAND3_X1 u2_u3_u2_U98 (.ZN( u2_u3_u2_n110 ) , .A2( u2_u3_u2_n131 ) , .A3( u2_u3_u2_n139 ) , .A1( u2_u3_u2_n154 ) );
  NAND3_X1 u2_u3_u2_U99 (.A2( u2_u3_u2_n100 ) , .ZN( u2_u3_u2_n101 ) , .A1( u2_u3_u2_n104 ) , .A3( u2_u3_u2_n114 ) );
  OAI22_X1 u2_u3_u3_U10 (.B1( u2_u3_u3_n113 ) , .A2( u2_u3_u3_n135 ) , .A1( u2_u3_u3_n150 ) , .B2( u2_u3_u3_n164 ) , .ZN( u2_u3_u3_n98 ) );
  OAI211_X1 u2_u3_u3_U11 (.B( u2_u3_u3_n106 ) , .ZN( u2_u3_u3_n119 ) , .C2( u2_u3_u3_n128 ) , .C1( u2_u3_u3_n167 ) , .A( u2_u3_u3_n181 ) );
  AOI221_X1 u2_u3_u3_U12 (.C1( u2_u3_u3_n105 ) , .ZN( u2_u3_u3_n106 ) , .A( u2_u3_u3_n131 ) , .B2( u2_u3_u3_n132 ) , .C2( u2_u3_u3_n133 ) , .B1( u2_u3_u3_n169 ) );
  INV_X1 u2_u3_u3_U13 (.ZN( u2_u3_u3_n181 ) , .A( u2_u3_u3_n98 ) );
  NAND2_X1 u2_u3_u3_U14 (.ZN( u2_u3_u3_n105 ) , .A2( u2_u3_u3_n130 ) , .A1( u2_u3_u3_n155 ) );
  AOI22_X1 u2_u3_u3_U15 (.B1( u2_u3_u3_n115 ) , .A2( u2_u3_u3_n116 ) , .ZN( u2_u3_u3_n123 ) , .B2( u2_u3_u3_n133 ) , .A1( u2_u3_u3_n169 ) );
  NAND2_X1 u2_u3_u3_U16 (.ZN( u2_u3_u3_n116 ) , .A2( u2_u3_u3_n151 ) , .A1( u2_u3_u3_n182 ) );
  NOR2_X1 u2_u3_u3_U17 (.ZN( u2_u3_u3_n126 ) , .A2( u2_u3_u3_n150 ) , .A1( u2_u3_u3_n164 ) );
  AOI21_X1 u2_u3_u3_U18 (.ZN( u2_u3_u3_n112 ) , .B2( u2_u3_u3_n146 ) , .B1( u2_u3_u3_n155 ) , .A( u2_u3_u3_n167 ) );
  NAND2_X1 u2_u3_u3_U19 (.A1( u2_u3_u3_n135 ) , .ZN( u2_u3_u3_n142 ) , .A2( u2_u3_u3_n164 ) );
  NAND2_X1 u2_u3_u3_U20 (.ZN( u2_u3_u3_n132 ) , .A2( u2_u3_u3_n152 ) , .A1( u2_u3_u3_n156 ) );
  INV_X1 u2_u3_u3_U21 (.A( u2_u3_u3_n133 ) , .ZN( u2_u3_u3_n165 ) );
  AND2_X1 u2_u3_u3_U22 (.A2( u2_u3_u3_n113 ) , .A1( u2_u3_u3_n114 ) , .ZN( u2_u3_u3_n151 ) );
  INV_X1 u2_u3_u3_U23 (.A( u2_u3_u3_n135 ) , .ZN( u2_u3_u3_n170 ) );
  NAND2_X1 u2_u3_u3_U24 (.A1( u2_u3_u3_n107 ) , .A2( u2_u3_u3_n108 ) , .ZN( u2_u3_u3_n140 ) );
  NAND2_X1 u2_u3_u3_U25 (.ZN( u2_u3_u3_n117 ) , .A1( u2_u3_u3_n124 ) , .A2( u2_u3_u3_n148 ) );
  NAND2_X1 u2_u3_u3_U26 (.ZN( u2_u3_u3_n143 ) , .A1( u2_u3_u3_n165 ) , .A2( u2_u3_u3_n167 ) );
  INV_X1 u2_u3_u3_U27 (.A( u2_u3_u3_n130 ) , .ZN( u2_u3_u3_n177 ) );
  INV_X1 u2_u3_u3_U28 (.A( u2_u3_u3_n128 ) , .ZN( u2_u3_u3_n176 ) );
  INV_X1 u2_u3_u3_U29 (.A( u2_u3_u3_n155 ) , .ZN( u2_u3_u3_n174 ) );
  INV_X1 u2_u3_u3_U3 (.A( u2_u3_u3_n140 ) , .ZN( u2_u3_u3_n182 ) );
  INV_X1 u2_u3_u3_U30 (.A( u2_u3_u3_n139 ) , .ZN( u2_u3_u3_n185 ) );
  NOR2_X1 u2_u3_u3_U31 (.ZN( u2_u3_u3_n135 ) , .A2( u2_u3_u3_n141 ) , .A1( u2_u3_u3_n169 ) );
  OAI222_X1 u2_u3_u3_U32 (.C2( u2_u3_u3_n107 ) , .A2( u2_u3_u3_n108 ) , .B1( u2_u3_u3_n135 ) , .ZN( u2_u3_u3_n138 ) , .B2( u2_u3_u3_n146 ) , .C1( u2_u3_u3_n154 ) , .A1( u2_u3_u3_n164 ) );
  NOR4_X1 u2_u3_u3_U33 (.A4( u2_u3_u3_n157 ) , .A3( u2_u3_u3_n158 ) , .A2( u2_u3_u3_n159 ) , .A1( u2_u3_u3_n160 ) , .ZN( u2_u3_u3_n161 ) );
  AOI21_X1 u2_u3_u3_U34 (.B2( u2_u3_u3_n152 ) , .B1( u2_u3_u3_n153 ) , .ZN( u2_u3_u3_n158 ) , .A( u2_u3_u3_n164 ) );
  AOI21_X1 u2_u3_u3_U35 (.A( u2_u3_u3_n149 ) , .B2( u2_u3_u3_n150 ) , .B1( u2_u3_u3_n151 ) , .ZN( u2_u3_u3_n159 ) );
  AOI21_X1 u2_u3_u3_U36 (.A( u2_u3_u3_n154 ) , .B2( u2_u3_u3_n155 ) , .B1( u2_u3_u3_n156 ) , .ZN( u2_u3_u3_n157 ) );
  AOI211_X1 u2_u3_u3_U37 (.ZN( u2_u3_u3_n109 ) , .A( u2_u3_u3_n119 ) , .C2( u2_u3_u3_n129 ) , .B( u2_u3_u3_n138 ) , .C1( u2_u3_u3_n141 ) );
  AOI211_X1 u2_u3_u3_U38 (.B( u2_u3_u3_n119 ) , .A( u2_u3_u3_n120 ) , .C2( u2_u3_u3_n121 ) , .ZN( u2_u3_u3_n122 ) , .C1( u2_u3_u3_n179 ) );
  INV_X1 u2_u3_u3_U39 (.A( u2_u3_u3_n156 ) , .ZN( u2_u3_u3_n179 ) );
  INV_X1 u2_u3_u3_U4 (.A( u2_u3_u3_n129 ) , .ZN( u2_u3_u3_n183 ) );
  OAI22_X1 u2_u3_u3_U40 (.B1( u2_u3_u3_n118 ) , .ZN( u2_u3_u3_n120 ) , .A1( u2_u3_u3_n135 ) , .B2( u2_u3_u3_n154 ) , .A2( u2_u3_u3_n178 ) );
  AND3_X1 u2_u3_u3_U41 (.ZN( u2_u3_u3_n118 ) , .A2( u2_u3_u3_n124 ) , .A1( u2_u3_u3_n144 ) , .A3( u2_u3_u3_n152 ) );
  INV_X1 u2_u3_u3_U42 (.A( u2_u3_u3_n121 ) , .ZN( u2_u3_u3_n164 ) );
  NAND2_X1 u2_u3_u3_U43 (.ZN( u2_u3_u3_n133 ) , .A1( u2_u3_u3_n154 ) , .A2( u2_u3_u3_n164 ) );
  NOR2_X1 u2_u3_u3_U44 (.A1( u2_u3_u3_n113 ) , .ZN( u2_u3_u3_n131 ) , .A2( u2_u3_u3_n154 ) );
  NAND2_X1 u2_u3_u3_U45 (.A1( u2_u3_u3_n103 ) , .ZN( u2_u3_u3_n150 ) , .A2( u2_u3_u3_n99 ) );
  NAND2_X1 u2_u3_u3_U46 (.A2( u2_u3_u3_n102 ) , .ZN( u2_u3_u3_n155 ) , .A1( u2_u3_u3_n97 ) );
  OAI211_X1 u2_u3_u3_U47 (.B( u2_u3_u3_n127 ) , .ZN( u2_u3_u3_n139 ) , .C1( u2_u3_u3_n150 ) , .C2( u2_u3_u3_n154 ) , .A( u2_u3_u3_n184 ) );
  INV_X1 u2_u3_u3_U48 (.A( u2_u3_u3_n125 ) , .ZN( u2_u3_u3_n184 ) );
  AOI221_X1 u2_u3_u3_U49 (.A( u2_u3_u3_n126 ) , .ZN( u2_u3_u3_n127 ) , .C2( u2_u3_u3_n132 ) , .C1( u2_u3_u3_n169 ) , .B2( u2_u3_u3_n170 ) , .B1( u2_u3_u3_n174 ) );
  INV_X1 u2_u3_u3_U5 (.A( u2_u3_u3_n117 ) , .ZN( u2_u3_u3_n178 ) );
  OAI22_X1 u2_u3_u3_U50 (.A1( u2_u3_u3_n124 ) , .ZN( u2_u3_u3_n125 ) , .B2( u2_u3_u3_n145 ) , .A2( u2_u3_u3_n165 ) , .B1( u2_u3_u3_n167 ) );
  INV_X1 u2_u3_u3_U51 (.A( u2_u3_u3_n141 ) , .ZN( u2_u3_u3_n167 ) );
  AOI21_X1 u2_u3_u3_U52 (.B2( u2_u3_u3_n114 ) , .B1( u2_u3_u3_n146 ) , .A( u2_u3_u3_n154 ) , .ZN( u2_u3_u3_n94 ) );
  AOI21_X1 u2_u3_u3_U53 (.ZN( u2_u3_u3_n110 ) , .B2( u2_u3_u3_n142 ) , .B1( u2_u3_u3_n186 ) , .A( u2_u3_u3_n95 ) );
  INV_X1 u2_u3_u3_U54 (.A( u2_u3_u3_n145 ) , .ZN( u2_u3_u3_n186 ) );
  AOI21_X1 u2_u3_u3_U55 (.B1( u2_u3_u3_n124 ) , .A( u2_u3_u3_n149 ) , .B2( u2_u3_u3_n155 ) , .ZN( u2_u3_u3_n95 ) );
  INV_X1 u2_u3_u3_U56 (.A( u2_u3_u3_n149 ) , .ZN( u2_u3_u3_n169 ) );
  NAND2_X1 u2_u3_u3_U57 (.ZN( u2_u3_u3_n124 ) , .A1( u2_u3_u3_n96 ) , .A2( u2_u3_u3_n97 ) );
  NAND2_X1 u2_u3_u3_U58 (.A2( u2_u3_u3_n100 ) , .ZN( u2_u3_u3_n146 ) , .A1( u2_u3_u3_n96 ) );
  NAND2_X1 u2_u3_u3_U59 (.A1( u2_u3_u3_n101 ) , .ZN( u2_u3_u3_n145 ) , .A2( u2_u3_u3_n99 ) );
  AOI221_X1 u2_u3_u3_U6 (.A( u2_u3_u3_n131 ) , .C2( u2_u3_u3_n132 ) , .C1( u2_u3_u3_n133 ) , .ZN( u2_u3_u3_n134 ) , .B1( u2_u3_u3_n143 ) , .B2( u2_u3_u3_n177 ) );
  NAND2_X1 u2_u3_u3_U60 (.A1( u2_u3_u3_n100 ) , .ZN( u2_u3_u3_n156 ) , .A2( u2_u3_u3_n99 ) );
  NAND2_X1 u2_u3_u3_U61 (.A2( u2_u3_u3_n101 ) , .A1( u2_u3_u3_n104 ) , .ZN( u2_u3_u3_n148 ) );
  NAND2_X1 u2_u3_u3_U62 (.A1( u2_u3_u3_n100 ) , .A2( u2_u3_u3_n102 ) , .ZN( u2_u3_u3_n128 ) );
  NAND2_X1 u2_u3_u3_U63 (.A2( u2_u3_u3_n101 ) , .A1( u2_u3_u3_n102 ) , .ZN( u2_u3_u3_n152 ) );
  NAND2_X1 u2_u3_u3_U64 (.A2( u2_u3_u3_n101 ) , .ZN( u2_u3_u3_n114 ) , .A1( u2_u3_u3_n96 ) );
  NAND2_X1 u2_u3_u3_U65 (.ZN( u2_u3_u3_n107 ) , .A1( u2_u3_u3_n97 ) , .A2( u2_u3_u3_n99 ) );
  NAND2_X1 u2_u3_u3_U66 (.A2( u2_u3_u3_n100 ) , .A1( u2_u3_u3_n104 ) , .ZN( u2_u3_u3_n113 ) );
  NAND2_X1 u2_u3_u3_U67 (.A1( u2_u3_u3_n104 ) , .ZN( u2_u3_u3_n153 ) , .A2( u2_u3_u3_n97 ) );
  NAND2_X1 u2_u3_u3_U68 (.A2( u2_u3_u3_n103 ) , .A1( u2_u3_u3_n104 ) , .ZN( u2_u3_u3_n130 ) );
  NAND2_X1 u2_u3_u3_U69 (.A2( u2_u3_u3_n103 ) , .ZN( u2_u3_u3_n144 ) , .A1( u2_u3_u3_n96 ) );
  OAI22_X1 u2_u3_u3_U7 (.B2( u2_u3_u3_n147 ) , .A2( u2_u3_u3_n148 ) , .ZN( u2_u3_u3_n160 ) , .B1( u2_u3_u3_n165 ) , .A1( u2_u3_u3_n168 ) );
  NAND2_X1 u2_u3_u3_U70 (.A1( u2_u3_u3_n102 ) , .A2( u2_u3_u3_n103 ) , .ZN( u2_u3_u3_n108 ) );
  NOR2_X1 u2_u3_u3_U71 (.A2( u2_u3_X_19 ) , .A1( u2_u3_X_20 ) , .ZN( u2_u3_u3_n99 ) );
  NOR2_X1 u2_u3_u3_U72 (.A2( u2_u3_X_21 ) , .A1( u2_u3_X_24 ) , .ZN( u2_u3_u3_n103 ) );
  NOR2_X1 u2_u3_u3_U73 (.A2( u2_u3_X_24 ) , .A1( u2_u3_u3_n171 ) , .ZN( u2_u3_u3_n97 ) );
  NOR2_X1 u2_u3_u3_U74 (.A2( u2_u3_X_23 ) , .ZN( u2_u3_u3_n141 ) , .A1( u2_u3_u3_n166 ) );
  NOR2_X1 u2_u3_u3_U75 (.A2( u2_u3_X_19 ) , .A1( u2_u3_u3_n172 ) , .ZN( u2_u3_u3_n96 ) );
  NAND2_X1 u2_u3_u3_U76 (.A1( u2_u3_X_22 ) , .A2( u2_u3_X_23 ) , .ZN( u2_u3_u3_n154 ) );
  NAND2_X1 u2_u3_u3_U77 (.A1( u2_u3_X_23 ) , .ZN( u2_u3_u3_n149 ) , .A2( u2_u3_u3_n166 ) );
  NOR2_X1 u2_u3_u3_U78 (.A2( u2_u3_X_22 ) , .A1( u2_u3_X_23 ) , .ZN( u2_u3_u3_n121 ) );
  AND2_X1 u2_u3_u3_U79 (.A1( u2_u3_X_24 ) , .ZN( u2_u3_u3_n101 ) , .A2( u2_u3_u3_n171 ) );
  AND3_X1 u2_u3_u3_U8 (.A3( u2_u3_u3_n144 ) , .A2( u2_u3_u3_n145 ) , .A1( u2_u3_u3_n146 ) , .ZN( u2_u3_u3_n147 ) );
  AND2_X1 u2_u3_u3_U80 (.A1( u2_u3_X_19 ) , .ZN( u2_u3_u3_n102 ) , .A2( u2_u3_u3_n172 ) );
  AND2_X1 u2_u3_u3_U81 (.A1( u2_u3_X_21 ) , .A2( u2_u3_X_24 ) , .ZN( u2_u3_u3_n100 ) );
  AND2_X1 u2_u3_u3_U82 (.A2( u2_u3_X_19 ) , .A1( u2_u3_X_20 ) , .ZN( u2_u3_u3_n104 ) );
  INV_X1 u2_u3_u3_U83 (.A( u2_u3_X_22 ) , .ZN( u2_u3_u3_n166 ) );
  INV_X1 u2_u3_u3_U84 (.A( u2_u3_X_21 ) , .ZN( u2_u3_u3_n171 ) );
  INV_X1 u2_u3_u3_U85 (.A( u2_u3_X_20 ) , .ZN( u2_u3_u3_n172 ) );
  NAND4_X1 u2_u3_u3_U86 (.ZN( u2_out3_26 ) , .A4( u2_u3_u3_n109 ) , .A3( u2_u3_u3_n110 ) , .A2( u2_u3_u3_n111 ) , .A1( u2_u3_u3_n173 ) );
  INV_X1 u2_u3_u3_U87 (.ZN( u2_u3_u3_n173 ) , .A( u2_u3_u3_n94 ) );
  OAI21_X1 u2_u3_u3_U88 (.ZN( u2_u3_u3_n111 ) , .B2( u2_u3_u3_n117 ) , .A( u2_u3_u3_n133 ) , .B1( u2_u3_u3_n176 ) );
  NAND4_X1 u2_u3_u3_U89 (.ZN( u2_out3_20 ) , .A4( u2_u3_u3_n122 ) , .A3( u2_u3_u3_n123 ) , .A1( u2_u3_u3_n175 ) , .A2( u2_u3_u3_n180 ) );
  INV_X1 u2_u3_u3_U9 (.A( u2_u3_u3_n143 ) , .ZN( u2_u3_u3_n168 ) );
  INV_X1 u2_u3_u3_U90 (.A( u2_u3_u3_n126 ) , .ZN( u2_u3_u3_n180 ) );
  INV_X1 u2_u3_u3_U91 (.A( u2_u3_u3_n112 ) , .ZN( u2_u3_u3_n175 ) );
  NAND4_X1 u2_u3_u3_U92 (.ZN( u2_out3_1 ) , .A4( u2_u3_u3_n161 ) , .A3( u2_u3_u3_n162 ) , .A2( u2_u3_u3_n163 ) , .A1( u2_u3_u3_n185 ) );
  NAND2_X1 u2_u3_u3_U93 (.ZN( u2_u3_u3_n163 ) , .A2( u2_u3_u3_n170 ) , .A1( u2_u3_u3_n176 ) );
  AOI22_X1 u2_u3_u3_U94 (.B2( u2_u3_u3_n140 ) , .B1( u2_u3_u3_n141 ) , .A2( u2_u3_u3_n142 ) , .ZN( u2_u3_u3_n162 ) , .A1( u2_u3_u3_n177 ) );
  OAI222_X1 u2_u3_u3_U95 (.C1( u2_u3_u3_n128 ) , .ZN( u2_u3_u3_n137 ) , .B1( u2_u3_u3_n148 ) , .A2( u2_u3_u3_n150 ) , .B2( u2_u3_u3_n154 ) , .C2( u2_u3_u3_n164 ) , .A1( u2_u3_u3_n167 ) );
  OR4_X1 u2_u3_u3_U96 (.ZN( u2_out3_10 ) , .A4( u2_u3_u3_n136 ) , .A3( u2_u3_u3_n137 ) , .A1( u2_u3_u3_n138 ) , .A2( u2_u3_u3_n139 ) );
  OAI221_X1 u2_u3_u3_U97 (.A( u2_u3_u3_n134 ) , .B2( u2_u3_u3_n135 ) , .ZN( u2_u3_u3_n136 ) , .C1( u2_u3_u3_n149 ) , .B1( u2_u3_u3_n151 ) , .C2( u2_u3_u3_n183 ) );
  NAND3_X1 u2_u3_u3_U98 (.A1( u2_u3_u3_n114 ) , .ZN( u2_u3_u3_n115 ) , .A2( u2_u3_u3_n145 ) , .A3( u2_u3_u3_n153 ) );
  NAND3_X1 u2_u3_u3_U99 (.ZN( u2_u3_u3_n129 ) , .A2( u2_u3_u3_n144 ) , .A1( u2_u3_u3_n153 ) , .A3( u2_u3_u3_n182 ) );
  OAI22_X1 u2_u3_u4_U10 (.B2( u2_u3_u4_n135 ) , .ZN( u2_u3_u4_n137 ) , .B1( u2_u3_u4_n153 ) , .A1( u2_u3_u4_n155 ) , .A2( u2_u3_u4_n171 ) );
  AND3_X1 u2_u3_u4_U11 (.A2( u2_u3_u4_n134 ) , .ZN( u2_u3_u4_n135 ) , .A3( u2_u3_u4_n145 ) , .A1( u2_u3_u4_n157 ) );
  OR3_X1 u2_u3_u4_U12 (.A3( u2_u3_u4_n114 ) , .A2( u2_u3_u4_n115 ) , .A1( u2_u3_u4_n116 ) , .ZN( u2_u3_u4_n136 ) );
  AOI21_X1 u2_u3_u4_U13 (.A( u2_u3_u4_n113 ) , .ZN( u2_u3_u4_n116 ) , .B2( u2_u3_u4_n173 ) , .B1( u2_u3_u4_n174 ) );
  AOI21_X1 u2_u3_u4_U14 (.ZN( u2_u3_u4_n115 ) , .B2( u2_u3_u4_n145 ) , .B1( u2_u3_u4_n146 ) , .A( u2_u3_u4_n156 ) );
  OAI22_X1 u2_u3_u4_U15 (.ZN( u2_u3_u4_n114 ) , .A2( u2_u3_u4_n121 ) , .B1( u2_u3_u4_n160 ) , .B2( u2_u3_u4_n170 ) , .A1( u2_u3_u4_n171 ) );
  NAND2_X1 u2_u3_u4_U16 (.ZN( u2_u3_u4_n132 ) , .A2( u2_u3_u4_n170 ) , .A1( u2_u3_u4_n173 ) );
  AOI21_X1 u2_u3_u4_U17 (.B2( u2_u3_u4_n160 ) , .B1( u2_u3_u4_n161 ) , .ZN( u2_u3_u4_n162 ) , .A( u2_u3_u4_n170 ) );
  AOI21_X1 u2_u3_u4_U18 (.ZN( u2_u3_u4_n107 ) , .B2( u2_u3_u4_n143 ) , .A( u2_u3_u4_n174 ) , .B1( u2_u3_u4_n184 ) );
  AOI21_X1 u2_u3_u4_U19 (.B2( u2_u3_u4_n158 ) , .B1( u2_u3_u4_n159 ) , .ZN( u2_u3_u4_n163 ) , .A( u2_u3_u4_n174 ) );
  AOI21_X1 u2_u3_u4_U20 (.A( u2_u3_u4_n153 ) , .B2( u2_u3_u4_n154 ) , .B1( u2_u3_u4_n155 ) , .ZN( u2_u3_u4_n165 ) );
  AOI21_X1 u2_u3_u4_U21 (.A( u2_u3_u4_n156 ) , .B2( u2_u3_u4_n157 ) , .ZN( u2_u3_u4_n164 ) , .B1( u2_u3_u4_n184 ) );
  INV_X1 u2_u3_u4_U22 (.A( u2_u3_u4_n138 ) , .ZN( u2_u3_u4_n170 ) );
  AND2_X1 u2_u3_u4_U23 (.A2( u2_u3_u4_n120 ) , .ZN( u2_u3_u4_n155 ) , .A1( u2_u3_u4_n160 ) );
  INV_X1 u2_u3_u4_U24 (.A( u2_u3_u4_n156 ) , .ZN( u2_u3_u4_n175 ) );
  NAND2_X1 u2_u3_u4_U25 (.A2( u2_u3_u4_n118 ) , .ZN( u2_u3_u4_n131 ) , .A1( u2_u3_u4_n147 ) );
  NAND2_X1 u2_u3_u4_U26 (.A1( u2_u3_u4_n119 ) , .A2( u2_u3_u4_n120 ) , .ZN( u2_u3_u4_n130 ) );
  NAND2_X1 u2_u3_u4_U27 (.ZN( u2_u3_u4_n117 ) , .A2( u2_u3_u4_n118 ) , .A1( u2_u3_u4_n148 ) );
  NAND2_X1 u2_u3_u4_U28 (.ZN( u2_u3_u4_n129 ) , .A1( u2_u3_u4_n134 ) , .A2( u2_u3_u4_n148 ) );
  AND3_X1 u2_u3_u4_U29 (.A1( u2_u3_u4_n119 ) , .A2( u2_u3_u4_n143 ) , .A3( u2_u3_u4_n154 ) , .ZN( u2_u3_u4_n161 ) );
  NOR2_X1 u2_u3_u4_U3 (.ZN( u2_u3_u4_n121 ) , .A1( u2_u3_u4_n181 ) , .A2( u2_u3_u4_n182 ) );
  AND2_X1 u2_u3_u4_U30 (.A1( u2_u3_u4_n145 ) , .A2( u2_u3_u4_n147 ) , .ZN( u2_u3_u4_n159 ) );
  INV_X1 u2_u3_u4_U31 (.A( u2_u3_u4_n158 ) , .ZN( u2_u3_u4_n182 ) );
  INV_X1 u2_u3_u4_U32 (.ZN( u2_u3_u4_n181 ) , .A( u2_u3_u4_n96 ) );
  INV_X1 u2_u3_u4_U33 (.A( u2_u3_u4_n144 ) , .ZN( u2_u3_u4_n179 ) );
  INV_X1 u2_u3_u4_U34 (.A( u2_u3_u4_n157 ) , .ZN( u2_u3_u4_n178 ) );
  NAND2_X1 u2_u3_u4_U35 (.A2( u2_u3_u4_n154 ) , .A1( u2_u3_u4_n96 ) , .ZN( u2_u3_u4_n97 ) );
  INV_X1 u2_u3_u4_U36 (.ZN( u2_u3_u4_n186 ) , .A( u2_u3_u4_n95 ) );
  OAI221_X1 u2_u3_u4_U37 (.C1( u2_u3_u4_n134 ) , .B1( u2_u3_u4_n158 ) , .B2( u2_u3_u4_n171 ) , .C2( u2_u3_u4_n173 ) , .A( u2_u3_u4_n94 ) , .ZN( u2_u3_u4_n95 ) );
  AOI222_X1 u2_u3_u4_U38 (.B2( u2_u3_u4_n132 ) , .A1( u2_u3_u4_n138 ) , .C2( u2_u3_u4_n175 ) , .A2( u2_u3_u4_n179 ) , .C1( u2_u3_u4_n181 ) , .B1( u2_u3_u4_n185 ) , .ZN( u2_u3_u4_n94 ) );
  INV_X1 u2_u3_u4_U39 (.A( u2_u3_u4_n113 ) , .ZN( u2_u3_u4_n185 ) );
  INV_X1 u2_u3_u4_U4 (.A( u2_u3_u4_n117 ) , .ZN( u2_u3_u4_n184 ) );
  INV_X1 u2_u3_u4_U40 (.A( u2_u3_u4_n143 ) , .ZN( u2_u3_u4_n183 ) );
  NOR2_X1 u2_u3_u4_U41 (.ZN( u2_u3_u4_n138 ) , .A1( u2_u3_u4_n168 ) , .A2( u2_u3_u4_n169 ) );
  NOR2_X1 u2_u3_u4_U42 (.A1( u2_u3_u4_n150 ) , .A2( u2_u3_u4_n152 ) , .ZN( u2_u3_u4_n153 ) );
  NOR2_X1 u2_u3_u4_U43 (.A2( u2_u3_u4_n128 ) , .A1( u2_u3_u4_n138 ) , .ZN( u2_u3_u4_n156 ) );
  AOI22_X1 u2_u3_u4_U44 (.B2( u2_u3_u4_n122 ) , .A1( u2_u3_u4_n123 ) , .ZN( u2_u3_u4_n124 ) , .B1( u2_u3_u4_n128 ) , .A2( u2_u3_u4_n172 ) );
  INV_X1 u2_u3_u4_U45 (.A( u2_u3_u4_n153 ) , .ZN( u2_u3_u4_n172 ) );
  NAND2_X1 u2_u3_u4_U46 (.A2( u2_u3_u4_n120 ) , .ZN( u2_u3_u4_n123 ) , .A1( u2_u3_u4_n161 ) );
  AOI22_X1 u2_u3_u4_U47 (.B2( u2_u3_u4_n132 ) , .A2( u2_u3_u4_n133 ) , .ZN( u2_u3_u4_n140 ) , .A1( u2_u3_u4_n150 ) , .B1( u2_u3_u4_n179 ) );
  NAND2_X1 u2_u3_u4_U48 (.ZN( u2_u3_u4_n133 ) , .A2( u2_u3_u4_n146 ) , .A1( u2_u3_u4_n154 ) );
  NAND2_X1 u2_u3_u4_U49 (.A1( u2_u3_u4_n103 ) , .ZN( u2_u3_u4_n154 ) , .A2( u2_u3_u4_n98 ) );
  NOR4_X1 u2_u3_u4_U5 (.A4( u2_u3_u4_n106 ) , .A3( u2_u3_u4_n107 ) , .A2( u2_u3_u4_n108 ) , .A1( u2_u3_u4_n109 ) , .ZN( u2_u3_u4_n110 ) );
  NAND2_X1 u2_u3_u4_U50 (.A1( u2_u3_u4_n101 ) , .ZN( u2_u3_u4_n158 ) , .A2( u2_u3_u4_n99 ) );
  AOI21_X1 u2_u3_u4_U51 (.ZN( u2_u3_u4_n127 ) , .A( u2_u3_u4_n136 ) , .B2( u2_u3_u4_n150 ) , .B1( u2_u3_u4_n180 ) );
  INV_X1 u2_u3_u4_U52 (.A( u2_u3_u4_n160 ) , .ZN( u2_u3_u4_n180 ) );
  NAND2_X1 u2_u3_u4_U53 (.A2( u2_u3_u4_n104 ) , .A1( u2_u3_u4_n105 ) , .ZN( u2_u3_u4_n146 ) );
  NAND2_X1 u2_u3_u4_U54 (.A2( u2_u3_u4_n101 ) , .A1( u2_u3_u4_n102 ) , .ZN( u2_u3_u4_n160 ) );
  NAND2_X1 u2_u3_u4_U55 (.ZN( u2_u3_u4_n134 ) , .A1( u2_u3_u4_n98 ) , .A2( u2_u3_u4_n99 ) );
  NAND2_X1 u2_u3_u4_U56 (.A1( u2_u3_u4_n103 ) , .A2( u2_u3_u4_n104 ) , .ZN( u2_u3_u4_n143 ) );
  NAND2_X1 u2_u3_u4_U57 (.A2( u2_u3_u4_n105 ) , .ZN( u2_u3_u4_n145 ) , .A1( u2_u3_u4_n98 ) );
  NAND2_X1 u2_u3_u4_U58 (.A1( u2_u3_u4_n100 ) , .A2( u2_u3_u4_n105 ) , .ZN( u2_u3_u4_n120 ) );
  NAND2_X1 u2_u3_u4_U59 (.A1( u2_u3_u4_n102 ) , .A2( u2_u3_u4_n104 ) , .ZN( u2_u3_u4_n148 ) );
  AOI21_X1 u2_u3_u4_U6 (.ZN( u2_u3_u4_n106 ) , .B2( u2_u3_u4_n146 ) , .B1( u2_u3_u4_n158 ) , .A( u2_u3_u4_n170 ) );
  NAND2_X1 u2_u3_u4_U60 (.A2( u2_u3_u4_n100 ) , .A1( u2_u3_u4_n103 ) , .ZN( u2_u3_u4_n157 ) );
  INV_X1 u2_u3_u4_U61 (.A( u2_u3_u4_n150 ) , .ZN( u2_u3_u4_n173 ) );
  INV_X1 u2_u3_u4_U62 (.A( u2_u3_u4_n152 ) , .ZN( u2_u3_u4_n171 ) );
  NAND2_X1 u2_u3_u4_U63 (.A1( u2_u3_u4_n100 ) , .ZN( u2_u3_u4_n118 ) , .A2( u2_u3_u4_n99 ) );
  NAND2_X1 u2_u3_u4_U64 (.A2( u2_u3_u4_n100 ) , .A1( u2_u3_u4_n102 ) , .ZN( u2_u3_u4_n144 ) );
  NAND2_X1 u2_u3_u4_U65 (.A2( u2_u3_u4_n101 ) , .A1( u2_u3_u4_n105 ) , .ZN( u2_u3_u4_n96 ) );
  INV_X1 u2_u3_u4_U66 (.A( u2_u3_u4_n128 ) , .ZN( u2_u3_u4_n174 ) );
  NAND2_X1 u2_u3_u4_U67 (.A2( u2_u3_u4_n102 ) , .ZN( u2_u3_u4_n119 ) , .A1( u2_u3_u4_n98 ) );
  NAND2_X1 u2_u3_u4_U68 (.A2( u2_u3_u4_n101 ) , .A1( u2_u3_u4_n103 ) , .ZN( u2_u3_u4_n147 ) );
  NAND2_X1 u2_u3_u4_U69 (.A2( u2_u3_u4_n104 ) , .ZN( u2_u3_u4_n113 ) , .A1( u2_u3_u4_n99 ) );
  AOI21_X1 u2_u3_u4_U7 (.ZN( u2_u3_u4_n109 ) , .A( u2_u3_u4_n153 ) , .B1( u2_u3_u4_n159 ) , .B2( u2_u3_u4_n184 ) );
  NOR2_X1 u2_u3_u4_U70 (.A2( u2_u3_X_28 ) , .ZN( u2_u3_u4_n150 ) , .A1( u2_u3_u4_n168 ) );
  NOR2_X1 u2_u3_u4_U71 (.A2( u2_u3_X_29 ) , .ZN( u2_u3_u4_n152 ) , .A1( u2_u3_u4_n169 ) );
  NOR2_X1 u2_u3_u4_U72 (.A2( u2_u3_X_30 ) , .ZN( u2_u3_u4_n105 ) , .A1( u2_u3_u4_n176 ) );
  NOR2_X1 u2_u3_u4_U73 (.A2( u2_u3_X_26 ) , .ZN( u2_u3_u4_n100 ) , .A1( u2_u3_u4_n177 ) );
  NOR2_X1 u2_u3_u4_U74 (.A2( u2_u3_X_28 ) , .A1( u2_u3_X_29 ) , .ZN( u2_u3_u4_n128 ) );
  NOR2_X1 u2_u3_u4_U75 (.A2( u2_u3_X_27 ) , .A1( u2_u3_X_30 ) , .ZN( u2_u3_u4_n102 ) );
  NOR2_X1 u2_u3_u4_U76 (.A2( u2_u3_X_25 ) , .A1( u2_u3_X_26 ) , .ZN( u2_u3_u4_n98 ) );
  AND2_X1 u2_u3_u4_U77 (.A2( u2_u3_X_25 ) , .A1( u2_u3_X_26 ) , .ZN( u2_u3_u4_n104 ) );
  AND2_X1 u2_u3_u4_U78 (.A1( u2_u3_X_30 ) , .A2( u2_u3_u4_n176 ) , .ZN( u2_u3_u4_n99 ) );
  AND2_X1 u2_u3_u4_U79 (.A1( u2_u3_X_26 ) , .ZN( u2_u3_u4_n101 ) , .A2( u2_u3_u4_n177 ) );
  AOI21_X1 u2_u3_u4_U8 (.ZN( u2_u3_u4_n108 ) , .B2( u2_u3_u4_n134 ) , .B1( u2_u3_u4_n155 ) , .A( u2_u3_u4_n156 ) );
  AND2_X1 u2_u3_u4_U80 (.A1( u2_u3_X_27 ) , .A2( u2_u3_X_30 ) , .ZN( u2_u3_u4_n103 ) );
  INV_X1 u2_u3_u4_U81 (.A( u2_u3_X_28 ) , .ZN( u2_u3_u4_n169 ) );
  INV_X1 u2_u3_u4_U82 (.A( u2_u3_X_29 ) , .ZN( u2_u3_u4_n168 ) );
  INV_X1 u2_u3_u4_U83 (.A( u2_u3_X_25 ) , .ZN( u2_u3_u4_n177 ) );
  INV_X1 u2_u3_u4_U84 (.A( u2_u3_X_27 ) , .ZN( u2_u3_u4_n176 ) );
  NAND4_X1 u2_u3_u4_U85 (.ZN( u2_out3_25 ) , .A4( u2_u3_u4_n139 ) , .A3( u2_u3_u4_n140 ) , .A2( u2_u3_u4_n141 ) , .A1( u2_u3_u4_n142 ) );
  OAI21_X1 u2_u3_u4_U86 (.A( u2_u3_u4_n128 ) , .B2( u2_u3_u4_n129 ) , .B1( u2_u3_u4_n130 ) , .ZN( u2_u3_u4_n142 ) );
  OAI21_X1 u2_u3_u4_U87 (.B2( u2_u3_u4_n131 ) , .ZN( u2_u3_u4_n141 ) , .A( u2_u3_u4_n175 ) , .B1( u2_u3_u4_n183 ) );
  NAND4_X1 u2_u3_u4_U88 (.ZN( u2_out3_14 ) , .A4( u2_u3_u4_n124 ) , .A3( u2_u3_u4_n125 ) , .A2( u2_u3_u4_n126 ) , .A1( u2_u3_u4_n127 ) );
  AOI22_X1 u2_u3_u4_U89 (.B2( u2_u3_u4_n117 ) , .ZN( u2_u3_u4_n126 ) , .A1( u2_u3_u4_n129 ) , .B1( u2_u3_u4_n152 ) , .A2( u2_u3_u4_n175 ) );
  AOI211_X1 u2_u3_u4_U9 (.B( u2_u3_u4_n136 ) , .A( u2_u3_u4_n137 ) , .C2( u2_u3_u4_n138 ) , .ZN( u2_u3_u4_n139 ) , .C1( u2_u3_u4_n182 ) );
  AOI22_X1 u2_u3_u4_U90 (.ZN( u2_u3_u4_n125 ) , .B2( u2_u3_u4_n131 ) , .A2( u2_u3_u4_n132 ) , .B1( u2_u3_u4_n138 ) , .A1( u2_u3_u4_n178 ) );
  NAND4_X1 u2_u3_u4_U91 (.ZN( u2_out3_8 ) , .A4( u2_u3_u4_n110 ) , .A3( u2_u3_u4_n111 ) , .A2( u2_u3_u4_n112 ) , .A1( u2_u3_u4_n186 ) );
  NAND2_X1 u2_u3_u4_U92 (.ZN( u2_u3_u4_n112 ) , .A2( u2_u3_u4_n130 ) , .A1( u2_u3_u4_n150 ) );
  AOI22_X1 u2_u3_u4_U93 (.ZN( u2_u3_u4_n111 ) , .B2( u2_u3_u4_n132 ) , .A1( u2_u3_u4_n152 ) , .B1( u2_u3_u4_n178 ) , .A2( u2_u3_u4_n97 ) );
  AOI22_X1 u2_u3_u4_U94 (.B2( u2_u3_u4_n149 ) , .B1( u2_u3_u4_n150 ) , .A2( u2_u3_u4_n151 ) , .A1( u2_u3_u4_n152 ) , .ZN( u2_u3_u4_n167 ) );
  NOR4_X1 u2_u3_u4_U95 (.A4( u2_u3_u4_n162 ) , .A3( u2_u3_u4_n163 ) , .A2( u2_u3_u4_n164 ) , .A1( u2_u3_u4_n165 ) , .ZN( u2_u3_u4_n166 ) );
  NAND3_X1 u2_u3_u4_U96 (.ZN( u2_out3_3 ) , .A3( u2_u3_u4_n166 ) , .A1( u2_u3_u4_n167 ) , .A2( u2_u3_u4_n186 ) );
  NAND3_X1 u2_u3_u4_U97 (.A3( u2_u3_u4_n146 ) , .A2( u2_u3_u4_n147 ) , .A1( u2_u3_u4_n148 ) , .ZN( u2_u3_u4_n149 ) );
  NAND3_X1 u2_u3_u4_U98 (.A3( u2_u3_u4_n143 ) , .A2( u2_u3_u4_n144 ) , .A1( u2_u3_u4_n145 ) , .ZN( u2_u3_u4_n151 ) );
  NAND3_X1 u2_u3_u4_U99 (.A3( u2_u3_u4_n121 ) , .ZN( u2_u3_u4_n122 ) , .A2( u2_u3_u4_n144 ) , .A1( u2_u3_u4_n154 ) );
  INV_X1 u2_u3_u5_U10 (.A( u2_u3_u5_n121 ) , .ZN( u2_u3_u5_n177 ) );
  NOR3_X1 u2_u3_u5_U100 (.A3( u2_u3_u5_n141 ) , .A1( u2_u3_u5_n142 ) , .ZN( u2_u3_u5_n143 ) , .A2( u2_u3_u5_n191 ) );
  NAND4_X1 u2_u3_u5_U101 (.ZN( u2_out3_4 ) , .A4( u2_u3_u5_n112 ) , .A2( u2_u3_u5_n113 ) , .A1( u2_u3_u5_n114 ) , .A3( u2_u3_u5_n195 ) );
  AOI211_X1 u2_u3_u5_U102 (.A( u2_u3_u5_n110 ) , .C1( u2_u3_u5_n111 ) , .ZN( u2_u3_u5_n112 ) , .B( u2_u3_u5_n118 ) , .C2( u2_u3_u5_n177 ) );
  AOI222_X1 u2_u3_u5_U103 (.ZN( u2_u3_u5_n113 ) , .A1( u2_u3_u5_n131 ) , .C1( u2_u3_u5_n148 ) , .B2( u2_u3_u5_n174 ) , .C2( u2_u3_u5_n178 ) , .A2( u2_u3_u5_n179 ) , .B1( u2_u3_u5_n99 ) );
  NAND3_X1 u2_u3_u5_U104 (.A2( u2_u3_u5_n154 ) , .A3( u2_u3_u5_n158 ) , .A1( u2_u3_u5_n161 ) , .ZN( u2_u3_u5_n99 ) );
  NOR2_X1 u2_u3_u5_U11 (.ZN( u2_u3_u5_n160 ) , .A2( u2_u3_u5_n173 ) , .A1( u2_u3_u5_n177 ) );
  INV_X1 u2_u3_u5_U12 (.A( u2_u3_u5_n150 ) , .ZN( u2_u3_u5_n174 ) );
  AOI21_X1 u2_u3_u5_U13 (.A( u2_u3_u5_n160 ) , .B2( u2_u3_u5_n161 ) , .ZN( u2_u3_u5_n162 ) , .B1( u2_u3_u5_n192 ) );
  INV_X1 u2_u3_u5_U14 (.A( u2_u3_u5_n159 ) , .ZN( u2_u3_u5_n192 ) );
  AOI21_X1 u2_u3_u5_U15 (.A( u2_u3_u5_n156 ) , .B2( u2_u3_u5_n157 ) , .B1( u2_u3_u5_n158 ) , .ZN( u2_u3_u5_n163 ) );
  AOI21_X1 u2_u3_u5_U16 (.B2( u2_u3_u5_n139 ) , .B1( u2_u3_u5_n140 ) , .ZN( u2_u3_u5_n141 ) , .A( u2_u3_u5_n150 ) );
  OAI21_X1 u2_u3_u5_U17 (.A( u2_u3_u5_n133 ) , .B2( u2_u3_u5_n134 ) , .B1( u2_u3_u5_n135 ) , .ZN( u2_u3_u5_n142 ) );
  OAI21_X1 u2_u3_u5_U18 (.ZN( u2_u3_u5_n133 ) , .B2( u2_u3_u5_n147 ) , .A( u2_u3_u5_n173 ) , .B1( u2_u3_u5_n188 ) );
  NAND2_X1 u2_u3_u5_U19 (.A2( u2_u3_u5_n119 ) , .A1( u2_u3_u5_n123 ) , .ZN( u2_u3_u5_n137 ) );
  INV_X1 u2_u3_u5_U20 (.A( u2_u3_u5_n155 ) , .ZN( u2_u3_u5_n194 ) );
  NAND2_X1 u2_u3_u5_U21 (.A1( u2_u3_u5_n121 ) , .ZN( u2_u3_u5_n132 ) , .A2( u2_u3_u5_n172 ) );
  NAND2_X1 u2_u3_u5_U22 (.A2( u2_u3_u5_n122 ) , .ZN( u2_u3_u5_n136 ) , .A1( u2_u3_u5_n154 ) );
  NAND2_X1 u2_u3_u5_U23 (.A2( u2_u3_u5_n119 ) , .A1( u2_u3_u5_n120 ) , .ZN( u2_u3_u5_n159 ) );
  INV_X1 u2_u3_u5_U24 (.A( u2_u3_u5_n156 ) , .ZN( u2_u3_u5_n175 ) );
  INV_X1 u2_u3_u5_U25 (.A( u2_u3_u5_n158 ) , .ZN( u2_u3_u5_n188 ) );
  INV_X1 u2_u3_u5_U26 (.A( u2_u3_u5_n152 ) , .ZN( u2_u3_u5_n179 ) );
  INV_X1 u2_u3_u5_U27 (.A( u2_u3_u5_n140 ) , .ZN( u2_u3_u5_n182 ) );
  INV_X1 u2_u3_u5_U28 (.A( u2_u3_u5_n151 ) , .ZN( u2_u3_u5_n183 ) );
  INV_X1 u2_u3_u5_U29 (.A( u2_u3_u5_n123 ) , .ZN( u2_u3_u5_n185 ) );
  NOR2_X1 u2_u3_u5_U3 (.ZN( u2_u3_u5_n134 ) , .A1( u2_u3_u5_n183 ) , .A2( u2_u3_u5_n190 ) );
  INV_X1 u2_u3_u5_U30 (.A( u2_u3_u5_n161 ) , .ZN( u2_u3_u5_n184 ) );
  INV_X1 u2_u3_u5_U31 (.A( u2_u3_u5_n139 ) , .ZN( u2_u3_u5_n189 ) );
  INV_X1 u2_u3_u5_U32 (.A( u2_u3_u5_n157 ) , .ZN( u2_u3_u5_n190 ) );
  INV_X1 u2_u3_u5_U33 (.A( u2_u3_u5_n120 ) , .ZN( u2_u3_u5_n193 ) );
  NAND2_X1 u2_u3_u5_U34 (.ZN( u2_u3_u5_n111 ) , .A1( u2_u3_u5_n140 ) , .A2( u2_u3_u5_n155 ) );
  INV_X1 u2_u3_u5_U35 (.A( u2_u3_u5_n117 ) , .ZN( u2_u3_u5_n196 ) );
  OAI221_X1 u2_u3_u5_U36 (.A( u2_u3_u5_n116 ) , .ZN( u2_u3_u5_n117 ) , .B2( u2_u3_u5_n119 ) , .C1( u2_u3_u5_n153 ) , .C2( u2_u3_u5_n158 ) , .B1( u2_u3_u5_n172 ) );
  AOI222_X1 u2_u3_u5_U37 (.ZN( u2_u3_u5_n116 ) , .B2( u2_u3_u5_n145 ) , .C1( u2_u3_u5_n148 ) , .A2( u2_u3_u5_n174 ) , .C2( u2_u3_u5_n177 ) , .B1( u2_u3_u5_n187 ) , .A1( u2_u3_u5_n193 ) );
  INV_X1 u2_u3_u5_U38 (.A( u2_u3_u5_n115 ) , .ZN( u2_u3_u5_n187 ) );
  NOR2_X1 u2_u3_u5_U39 (.ZN( u2_u3_u5_n100 ) , .A1( u2_u3_u5_n170 ) , .A2( u2_u3_u5_n180 ) );
  INV_X1 u2_u3_u5_U4 (.A( u2_u3_u5_n138 ) , .ZN( u2_u3_u5_n191 ) );
  AOI22_X1 u2_u3_u5_U40 (.B2( u2_u3_u5_n131 ) , .A2( u2_u3_u5_n146 ) , .ZN( u2_u3_u5_n169 ) , .B1( u2_u3_u5_n174 ) , .A1( u2_u3_u5_n185 ) );
  NOR2_X1 u2_u3_u5_U41 (.A1( u2_u3_u5_n146 ) , .ZN( u2_u3_u5_n150 ) , .A2( u2_u3_u5_n173 ) );
  AOI21_X1 u2_u3_u5_U42 (.A( u2_u3_u5_n118 ) , .B2( u2_u3_u5_n145 ) , .ZN( u2_u3_u5_n168 ) , .B1( u2_u3_u5_n186 ) );
  INV_X1 u2_u3_u5_U43 (.A( u2_u3_u5_n122 ) , .ZN( u2_u3_u5_n186 ) );
  NOR2_X1 u2_u3_u5_U44 (.A1( u2_u3_u5_n146 ) , .ZN( u2_u3_u5_n152 ) , .A2( u2_u3_u5_n176 ) );
  NOR2_X1 u2_u3_u5_U45 (.A1( u2_u3_u5_n115 ) , .ZN( u2_u3_u5_n118 ) , .A2( u2_u3_u5_n153 ) );
  NOR2_X1 u2_u3_u5_U46 (.A2( u2_u3_u5_n145 ) , .ZN( u2_u3_u5_n156 ) , .A1( u2_u3_u5_n174 ) );
  NOR2_X1 u2_u3_u5_U47 (.ZN( u2_u3_u5_n121 ) , .A2( u2_u3_u5_n145 ) , .A1( u2_u3_u5_n176 ) );
  AOI22_X1 u2_u3_u5_U48 (.ZN( u2_u3_u5_n114 ) , .A2( u2_u3_u5_n137 ) , .A1( u2_u3_u5_n145 ) , .B2( u2_u3_u5_n175 ) , .B1( u2_u3_u5_n193 ) );
  OAI211_X1 u2_u3_u5_U49 (.B( u2_u3_u5_n124 ) , .A( u2_u3_u5_n125 ) , .C2( u2_u3_u5_n126 ) , .C1( u2_u3_u5_n127 ) , .ZN( u2_u3_u5_n128 ) );
  OAI21_X1 u2_u3_u5_U5 (.B2( u2_u3_u5_n136 ) , .B1( u2_u3_u5_n137 ) , .ZN( u2_u3_u5_n138 ) , .A( u2_u3_u5_n177 ) );
  NOR3_X1 u2_u3_u5_U50 (.ZN( u2_u3_u5_n127 ) , .A1( u2_u3_u5_n136 ) , .A3( u2_u3_u5_n148 ) , .A2( u2_u3_u5_n182 ) );
  OAI21_X1 u2_u3_u5_U51 (.ZN( u2_u3_u5_n124 ) , .A( u2_u3_u5_n177 ) , .B2( u2_u3_u5_n183 ) , .B1( u2_u3_u5_n189 ) );
  OAI21_X1 u2_u3_u5_U52 (.ZN( u2_u3_u5_n125 ) , .A( u2_u3_u5_n174 ) , .B2( u2_u3_u5_n185 ) , .B1( u2_u3_u5_n190 ) );
  AOI21_X1 u2_u3_u5_U53 (.A( u2_u3_u5_n153 ) , .B2( u2_u3_u5_n154 ) , .B1( u2_u3_u5_n155 ) , .ZN( u2_u3_u5_n164 ) );
  AOI21_X1 u2_u3_u5_U54 (.ZN( u2_u3_u5_n110 ) , .B1( u2_u3_u5_n122 ) , .B2( u2_u3_u5_n139 ) , .A( u2_u3_u5_n153 ) );
  INV_X1 u2_u3_u5_U55 (.A( u2_u3_u5_n153 ) , .ZN( u2_u3_u5_n176 ) );
  INV_X1 u2_u3_u5_U56 (.A( u2_u3_u5_n126 ) , .ZN( u2_u3_u5_n173 ) );
  AND2_X1 u2_u3_u5_U57 (.A2( u2_u3_u5_n104 ) , .A1( u2_u3_u5_n107 ) , .ZN( u2_u3_u5_n147 ) );
  AND2_X1 u2_u3_u5_U58 (.A2( u2_u3_u5_n104 ) , .A1( u2_u3_u5_n108 ) , .ZN( u2_u3_u5_n148 ) );
  NAND2_X1 u2_u3_u5_U59 (.A1( u2_u3_u5_n105 ) , .A2( u2_u3_u5_n106 ) , .ZN( u2_u3_u5_n158 ) );
  INV_X1 u2_u3_u5_U6 (.A( u2_u3_u5_n135 ) , .ZN( u2_u3_u5_n178 ) );
  NAND2_X1 u2_u3_u5_U60 (.A2( u2_u3_u5_n108 ) , .A1( u2_u3_u5_n109 ) , .ZN( u2_u3_u5_n139 ) );
  NAND2_X1 u2_u3_u5_U61 (.A1( u2_u3_u5_n106 ) , .A2( u2_u3_u5_n108 ) , .ZN( u2_u3_u5_n119 ) );
  NAND2_X1 u2_u3_u5_U62 (.A2( u2_u3_u5_n103 ) , .A1( u2_u3_u5_n105 ) , .ZN( u2_u3_u5_n140 ) );
  NAND2_X1 u2_u3_u5_U63 (.A2( u2_u3_u5_n104 ) , .A1( u2_u3_u5_n105 ) , .ZN( u2_u3_u5_n155 ) );
  NAND2_X1 u2_u3_u5_U64 (.A2( u2_u3_u5_n106 ) , .A1( u2_u3_u5_n107 ) , .ZN( u2_u3_u5_n122 ) );
  NAND2_X1 u2_u3_u5_U65 (.A2( u2_u3_u5_n100 ) , .A1( u2_u3_u5_n106 ) , .ZN( u2_u3_u5_n115 ) );
  NAND2_X1 u2_u3_u5_U66 (.A2( u2_u3_u5_n100 ) , .A1( u2_u3_u5_n103 ) , .ZN( u2_u3_u5_n161 ) );
  NAND2_X1 u2_u3_u5_U67 (.A1( u2_u3_u5_n105 ) , .A2( u2_u3_u5_n109 ) , .ZN( u2_u3_u5_n154 ) );
  INV_X1 u2_u3_u5_U68 (.A( u2_u3_u5_n146 ) , .ZN( u2_u3_u5_n172 ) );
  NAND2_X1 u2_u3_u5_U69 (.A1( u2_u3_u5_n103 ) , .A2( u2_u3_u5_n108 ) , .ZN( u2_u3_u5_n123 ) );
  OAI22_X1 u2_u3_u5_U7 (.B2( u2_u3_u5_n149 ) , .B1( u2_u3_u5_n150 ) , .A2( u2_u3_u5_n151 ) , .A1( u2_u3_u5_n152 ) , .ZN( u2_u3_u5_n165 ) );
  NAND2_X1 u2_u3_u5_U70 (.A2( u2_u3_u5_n103 ) , .A1( u2_u3_u5_n107 ) , .ZN( u2_u3_u5_n151 ) );
  NAND2_X1 u2_u3_u5_U71 (.A2( u2_u3_u5_n107 ) , .A1( u2_u3_u5_n109 ) , .ZN( u2_u3_u5_n120 ) );
  NAND2_X1 u2_u3_u5_U72 (.A2( u2_u3_u5_n100 ) , .A1( u2_u3_u5_n109 ) , .ZN( u2_u3_u5_n157 ) );
  AND2_X1 u2_u3_u5_U73 (.A2( u2_u3_u5_n100 ) , .A1( u2_u3_u5_n104 ) , .ZN( u2_u3_u5_n131 ) );
  INV_X1 u2_u3_u5_U74 (.A( u2_u3_u5_n102 ) , .ZN( u2_u3_u5_n195 ) );
  OAI221_X1 u2_u3_u5_U75 (.A( u2_u3_u5_n101 ) , .ZN( u2_u3_u5_n102 ) , .C2( u2_u3_u5_n115 ) , .C1( u2_u3_u5_n126 ) , .B1( u2_u3_u5_n134 ) , .B2( u2_u3_u5_n160 ) );
  OAI21_X1 u2_u3_u5_U76 (.ZN( u2_u3_u5_n101 ) , .B1( u2_u3_u5_n137 ) , .A( u2_u3_u5_n146 ) , .B2( u2_u3_u5_n147 ) );
  NOR2_X1 u2_u3_u5_U77 (.A2( u2_u3_X_34 ) , .A1( u2_u3_X_35 ) , .ZN( u2_u3_u5_n145 ) );
  NOR2_X1 u2_u3_u5_U78 (.A2( u2_u3_X_34 ) , .ZN( u2_u3_u5_n146 ) , .A1( u2_u3_u5_n171 ) );
  NOR2_X1 u2_u3_u5_U79 (.A2( u2_u3_X_31 ) , .A1( u2_u3_X_32 ) , .ZN( u2_u3_u5_n103 ) );
  NOR3_X1 u2_u3_u5_U8 (.A2( u2_u3_u5_n147 ) , .A1( u2_u3_u5_n148 ) , .ZN( u2_u3_u5_n149 ) , .A3( u2_u3_u5_n194 ) );
  NOR2_X1 u2_u3_u5_U80 (.A2( u2_u3_X_36 ) , .ZN( u2_u3_u5_n105 ) , .A1( u2_u3_u5_n180 ) );
  NOR2_X1 u2_u3_u5_U81 (.A2( u2_u3_X_33 ) , .ZN( u2_u3_u5_n108 ) , .A1( u2_u3_u5_n170 ) );
  NOR2_X1 u2_u3_u5_U82 (.A2( u2_u3_X_33 ) , .A1( u2_u3_X_36 ) , .ZN( u2_u3_u5_n107 ) );
  NOR2_X1 u2_u3_u5_U83 (.A2( u2_u3_X_31 ) , .ZN( u2_u3_u5_n104 ) , .A1( u2_u3_u5_n181 ) );
  NAND2_X1 u2_u3_u5_U84 (.A2( u2_u3_X_34 ) , .A1( u2_u3_X_35 ) , .ZN( u2_u3_u5_n153 ) );
  NAND2_X1 u2_u3_u5_U85 (.A1( u2_u3_X_34 ) , .ZN( u2_u3_u5_n126 ) , .A2( u2_u3_u5_n171 ) );
  AND2_X1 u2_u3_u5_U86 (.A1( u2_u3_X_31 ) , .A2( u2_u3_X_32 ) , .ZN( u2_u3_u5_n106 ) );
  AND2_X1 u2_u3_u5_U87 (.A1( u2_u3_X_31 ) , .ZN( u2_u3_u5_n109 ) , .A2( u2_u3_u5_n181 ) );
  INV_X1 u2_u3_u5_U88 (.A( u2_u3_X_33 ) , .ZN( u2_u3_u5_n180 ) );
  INV_X1 u2_u3_u5_U89 (.A( u2_u3_X_35 ) , .ZN( u2_u3_u5_n171 ) );
  NOR2_X1 u2_u3_u5_U9 (.ZN( u2_u3_u5_n135 ) , .A1( u2_u3_u5_n173 ) , .A2( u2_u3_u5_n176 ) );
  INV_X1 u2_u3_u5_U90 (.A( u2_u3_X_36 ) , .ZN( u2_u3_u5_n170 ) );
  INV_X1 u2_u3_u5_U91 (.A( u2_u3_X_32 ) , .ZN( u2_u3_u5_n181 ) );
  NAND4_X1 u2_u3_u5_U92 (.ZN( u2_out3_29 ) , .A4( u2_u3_u5_n129 ) , .A3( u2_u3_u5_n130 ) , .A2( u2_u3_u5_n168 ) , .A1( u2_u3_u5_n196 ) );
  AOI221_X1 u2_u3_u5_U93 (.A( u2_u3_u5_n128 ) , .ZN( u2_u3_u5_n129 ) , .C2( u2_u3_u5_n132 ) , .B2( u2_u3_u5_n159 ) , .B1( u2_u3_u5_n176 ) , .C1( u2_u3_u5_n184 ) );
  AOI222_X1 u2_u3_u5_U94 (.ZN( u2_u3_u5_n130 ) , .A2( u2_u3_u5_n146 ) , .B1( u2_u3_u5_n147 ) , .C2( u2_u3_u5_n175 ) , .B2( u2_u3_u5_n179 ) , .A1( u2_u3_u5_n188 ) , .C1( u2_u3_u5_n194 ) );
  NAND4_X1 u2_u3_u5_U95 (.ZN( u2_out3_19 ) , .A4( u2_u3_u5_n166 ) , .A3( u2_u3_u5_n167 ) , .A2( u2_u3_u5_n168 ) , .A1( u2_u3_u5_n169 ) );
  AOI22_X1 u2_u3_u5_U96 (.B2( u2_u3_u5_n145 ) , .A2( u2_u3_u5_n146 ) , .ZN( u2_u3_u5_n167 ) , .B1( u2_u3_u5_n182 ) , .A1( u2_u3_u5_n189 ) );
  NOR4_X1 u2_u3_u5_U97 (.A4( u2_u3_u5_n162 ) , .A3( u2_u3_u5_n163 ) , .A2( u2_u3_u5_n164 ) , .A1( u2_u3_u5_n165 ) , .ZN( u2_u3_u5_n166 ) );
  NAND4_X1 u2_u3_u5_U98 (.ZN( u2_out3_11 ) , .A4( u2_u3_u5_n143 ) , .A3( u2_u3_u5_n144 ) , .A2( u2_u3_u5_n169 ) , .A1( u2_u3_u5_n196 ) );
  AOI22_X1 u2_u3_u5_U99 (.A2( u2_u3_u5_n132 ) , .ZN( u2_u3_u5_n144 ) , .B2( u2_u3_u5_n145 ) , .B1( u2_u3_u5_n184 ) , .A1( u2_u3_u5_n194 ) );
  AND3_X1 u2_u3_u7_U10 (.A3( u2_u3_u7_n110 ) , .A2( u2_u3_u7_n127 ) , .A1( u2_u3_u7_n132 ) , .ZN( u2_u3_u7_n92 ) );
  OAI21_X1 u2_u3_u7_U11 (.A( u2_u3_u7_n161 ) , .B1( u2_u3_u7_n168 ) , .B2( u2_u3_u7_n173 ) , .ZN( u2_u3_u7_n91 ) );
  AOI211_X1 u2_u3_u7_U12 (.A( u2_u3_u7_n117 ) , .ZN( u2_u3_u7_n118 ) , .C2( u2_u3_u7_n126 ) , .C1( u2_u3_u7_n177 ) , .B( u2_u3_u7_n180 ) );
  OAI22_X1 u2_u3_u7_U13 (.B1( u2_u3_u7_n115 ) , .ZN( u2_u3_u7_n117 ) , .A2( u2_u3_u7_n133 ) , .A1( u2_u3_u7_n137 ) , .B2( u2_u3_u7_n162 ) );
  INV_X1 u2_u3_u7_U14 (.A( u2_u3_u7_n116 ) , .ZN( u2_u3_u7_n180 ) );
  NOR3_X1 u2_u3_u7_U15 (.ZN( u2_u3_u7_n115 ) , .A3( u2_u3_u7_n145 ) , .A2( u2_u3_u7_n168 ) , .A1( u2_u3_u7_n169 ) );
  OAI211_X1 u2_u3_u7_U16 (.B( u2_u3_u7_n122 ) , .A( u2_u3_u7_n123 ) , .C2( u2_u3_u7_n124 ) , .ZN( u2_u3_u7_n154 ) , .C1( u2_u3_u7_n162 ) );
  AOI222_X1 u2_u3_u7_U17 (.ZN( u2_u3_u7_n122 ) , .C2( u2_u3_u7_n126 ) , .C1( u2_u3_u7_n145 ) , .B1( u2_u3_u7_n161 ) , .A2( u2_u3_u7_n165 ) , .B2( u2_u3_u7_n170 ) , .A1( u2_u3_u7_n176 ) );
  INV_X1 u2_u3_u7_U18 (.A( u2_u3_u7_n133 ) , .ZN( u2_u3_u7_n176 ) );
  NOR3_X1 u2_u3_u7_U19 (.A2( u2_u3_u7_n134 ) , .A1( u2_u3_u7_n135 ) , .ZN( u2_u3_u7_n136 ) , .A3( u2_u3_u7_n171 ) );
  NOR2_X1 u2_u3_u7_U20 (.A1( u2_u3_u7_n130 ) , .A2( u2_u3_u7_n134 ) , .ZN( u2_u3_u7_n153 ) );
  INV_X1 u2_u3_u7_U21 (.A( u2_u3_u7_n101 ) , .ZN( u2_u3_u7_n165 ) );
  NOR2_X1 u2_u3_u7_U22 (.ZN( u2_u3_u7_n111 ) , .A2( u2_u3_u7_n134 ) , .A1( u2_u3_u7_n169 ) );
  AOI21_X1 u2_u3_u7_U23 (.ZN( u2_u3_u7_n104 ) , .B2( u2_u3_u7_n112 ) , .B1( u2_u3_u7_n127 ) , .A( u2_u3_u7_n164 ) );
  AOI21_X1 u2_u3_u7_U24 (.ZN( u2_u3_u7_n106 ) , .B1( u2_u3_u7_n133 ) , .B2( u2_u3_u7_n146 ) , .A( u2_u3_u7_n162 ) );
  AOI21_X1 u2_u3_u7_U25 (.A( u2_u3_u7_n101 ) , .ZN( u2_u3_u7_n107 ) , .B2( u2_u3_u7_n128 ) , .B1( u2_u3_u7_n175 ) );
  INV_X1 u2_u3_u7_U26 (.A( u2_u3_u7_n138 ) , .ZN( u2_u3_u7_n171 ) );
  INV_X1 u2_u3_u7_U27 (.A( u2_u3_u7_n131 ) , .ZN( u2_u3_u7_n177 ) );
  INV_X1 u2_u3_u7_U28 (.A( u2_u3_u7_n110 ) , .ZN( u2_u3_u7_n174 ) );
  NAND2_X1 u2_u3_u7_U29 (.A1( u2_u3_u7_n129 ) , .A2( u2_u3_u7_n132 ) , .ZN( u2_u3_u7_n149 ) );
  OAI21_X1 u2_u3_u7_U3 (.ZN( u2_u3_u7_n159 ) , .A( u2_u3_u7_n165 ) , .B2( u2_u3_u7_n171 ) , .B1( u2_u3_u7_n174 ) );
  NAND2_X1 u2_u3_u7_U30 (.A1( u2_u3_u7_n113 ) , .A2( u2_u3_u7_n124 ) , .ZN( u2_u3_u7_n130 ) );
  INV_X1 u2_u3_u7_U31 (.A( u2_u3_u7_n112 ) , .ZN( u2_u3_u7_n173 ) );
  INV_X1 u2_u3_u7_U32 (.A( u2_u3_u7_n128 ) , .ZN( u2_u3_u7_n168 ) );
  INV_X1 u2_u3_u7_U33 (.A( u2_u3_u7_n148 ) , .ZN( u2_u3_u7_n169 ) );
  INV_X1 u2_u3_u7_U34 (.A( u2_u3_u7_n127 ) , .ZN( u2_u3_u7_n179 ) );
  NOR2_X1 u2_u3_u7_U35 (.ZN( u2_u3_u7_n101 ) , .A2( u2_u3_u7_n150 ) , .A1( u2_u3_u7_n156 ) );
  AOI211_X1 u2_u3_u7_U36 (.B( u2_u3_u7_n154 ) , .A( u2_u3_u7_n155 ) , .C1( u2_u3_u7_n156 ) , .ZN( u2_u3_u7_n157 ) , .C2( u2_u3_u7_n172 ) );
  INV_X1 u2_u3_u7_U37 (.A( u2_u3_u7_n153 ) , .ZN( u2_u3_u7_n172 ) );
  AOI211_X1 u2_u3_u7_U38 (.B( u2_u3_u7_n139 ) , .A( u2_u3_u7_n140 ) , .C2( u2_u3_u7_n141 ) , .ZN( u2_u3_u7_n142 ) , .C1( u2_u3_u7_n156 ) );
  NAND4_X1 u2_u3_u7_U39 (.A3( u2_u3_u7_n127 ) , .A2( u2_u3_u7_n128 ) , .A1( u2_u3_u7_n129 ) , .ZN( u2_u3_u7_n141 ) , .A4( u2_u3_u7_n147 ) );
  INV_X1 u2_u3_u7_U4 (.A( u2_u3_u7_n111 ) , .ZN( u2_u3_u7_n170 ) );
  AOI21_X1 u2_u3_u7_U40 (.A( u2_u3_u7_n137 ) , .B1( u2_u3_u7_n138 ) , .ZN( u2_u3_u7_n139 ) , .B2( u2_u3_u7_n146 ) );
  OAI22_X1 u2_u3_u7_U41 (.B1( u2_u3_u7_n136 ) , .ZN( u2_u3_u7_n140 ) , .A1( u2_u3_u7_n153 ) , .B2( u2_u3_u7_n162 ) , .A2( u2_u3_u7_n164 ) );
  AOI21_X1 u2_u3_u7_U42 (.ZN( u2_u3_u7_n123 ) , .B1( u2_u3_u7_n165 ) , .B2( u2_u3_u7_n177 ) , .A( u2_u3_u7_n97 ) );
  AOI21_X1 u2_u3_u7_U43 (.B2( u2_u3_u7_n113 ) , .B1( u2_u3_u7_n124 ) , .A( u2_u3_u7_n125 ) , .ZN( u2_u3_u7_n97 ) );
  INV_X1 u2_u3_u7_U44 (.A( u2_u3_u7_n125 ) , .ZN( u2_u3_u7_n161 ) );
  INV_X1 u2_u3_u7_U45 (.A( u2_u3_u7_n152 ) , .ZN( u2_u3_u7_n162 ) );
  AOI22_X1 u2_u3_u7_U46 (.A2( u2_u3_u7_n114 ) , .ZN( u2_u3_u7_n119 ) , .B1( u2_u3_u7_n130 ) , .A1( u2_u3_u7_n156 ) , .B2( u2_u3_u7_n165 ) );
  NAND2_X1 u2_u3_u7_U47 (.A2( u2_u3_u7_n112 ) , .ZN( u2_u3_u7_n114 ) , .A1( u2_u3_u7_n175 ) );
  AND2_X1 u2_u3_u7_U48 (.ZN( u2_u3_u7_n145 ) , .A2( u2_u3_u7_n98 ) , .A1( u2_u3_u7_n99 ) );
  NOR2_X1 u2_u3_u7_U49 (.ZN( u2_u3_u7_n137 ) , .A1( u2_u3_u7_n150 ) , .A2( u2_u3_u7_n161 ) );
  INV_X1 u2_u3_u7_U5 (.A( u2_u3_u7_n149 ) , .ZN( u2_u3_u7_n175 ) );
  AOI21_X1 u2_u3_u7_U50 (.ZN( u2_u3_u7_n105 ) , .B2( u2_u3_u7_n110 ) , .A( u2_u3_u7_n125 ) , .B1( u2_u3_u7_n147 ) );
  NAND2_X1 u2_u3_u7_U51 (.ZN( u2_u3_u7_n146 ) , .A1( u2_u3_u7_n95 ) , .A2( u2_u3_u7_n98 ) );
  NAND2_X1 u2_u3_u7_U52 (.A2( u2_u3_u7_n103 ) , .ZN( u2_u3_u7_n147 ) , .A1( u2_u3_u7_n93 ) );
  NAND2_X1 u2_u3_u7_U53 (.A1( u2_u3_u7_n103 ) , .ZN( u2_u3_u7_n127 ) , .A2( u2_u3_u7_n99 ) );
  OR2_X1 u2_u3_u7_U54 (.ZN( u2_u3_u7_n126 ) , .A2( u2_u3_u7_n152 ) , .A1( u2_u3_u7_n156 ) );
  NAND2_X1 u2_u3_u7_U55 (.A2( u2_u3_u7_n102 ) , .A1( u2_u3_u7_n103 ) , .ZN( u2_u3_u7_n133 ) );
  NAND2_X1 u2_u3_u7_U56 (.ZN( u2_u3_u7_n112 ) , .A2( u2_u3_u7_n96 ) , .A1( u2_u3_u7_n99 ) );
  NAND2_X1 u2_u3_u7_U57 (.A2( u2_u3_u7_n102 ) , .ZN( u2_u3_u7_n128 ) , .A1( u2_u3_u7_n98 ) );
  NAND2_X1 u2_u3_u7_U58 (.A1( u2_u3_u7_n100 ) , .ZN( u2_u3_u7_n113 ) , .A2( u2_u3_u7_n93 ) );
  NAND2_X1 u2_u3_u7_U59 (.A2( u2_u3_u7_n102 ) , .ZN( u2_u3_u7_n124 ) , .A1( u2_u3_u7_n96 ) );
  INV_X1 u2_u3_u7_U6 (.A( u2_u3_u7_n154 ) , .ZN( u2_u3_u7_n178 ) );
  NAND2_X1 u2_u3_u7_U60 (.ZN( u2_u3_u7_n110 ) , .A1( u2_u3_u7_n95 ) , .A2( u2_u3_u7_n96 ) );
  INV_X1 u2_u3_u7_U61 (.A( u2_u3_u7_n150 ) , .ZN( u2_u3_u7_n164 ) );
  AND2_X1 u2_u3_u7_U62 (.ZN( u2_u3_u7_n134 ) , .A1( u2_u3_u7_n93 ) , .A2( u2_u3_u7_n98 ) );
  NAND2_X1 u2_u3_u7_U63 (.A1( u2_u3_u7_n100 ) , .A2( u2_u3_u7_n102 ) , .ZN( u2_u3_u7_n129 ) );
  NAND2_X1 u2_u3_u7_U64 (.A2( u2_u3_u7_n103 ) , .ZN( u2_u3_u7_n131 ) , .A1( u2_u3_u7_n95 ) );
  NAND2_X1 u2_u3_u7_U65 (.A1( u2_u3_u7_n100 ) , .ZN( u2_u3_u7_n138 ) , .A2( u2_u3_u7_n99 ) );
  NAND2_X1 u2_u3_u7_U66 (.ZN( u2_u3_u7_n132 ) , .A1( u2_u3_u7_n93 ) , .A2( u2_u3_u7_n96 ) );
  NAND2_X1 u2_u3_u7_U67 (.A1( u2_u3_u7_n100 ) , .ZN( u2_u3_u7_n148 ) , .A2( u2_u3_u7_n95 ) );
  NOR2_X1 u2_u3_u7_U68 (.A2( u2_u3_X_47 ) , .ZN( u2_u3_u7_n150 ) , .A1( u2_u3_u7_n163 ) );
  NOR2_X1 u2_u3_u7_U69 (.A2( u2_u3_X_43 ) , .A1( u2_u3_X_44 ) , .ZN( u2_u3_u7_n103 ) );
  AOI211_X1 u2_u3_u7_U7 (.ZN( u2_u3_u7_n116 ) , .A( u2_u3_u7_n155 ) , .C1( u2_u3_u7_n161 ) , .C2( u2_u3_u7_n171 ) , .B( u2_u3_u7_n94 ) );
  NOR2_X1 u2_u3_u7_U70 (.A2( u2_u3_X_48 ) , .A1( u2_u3_u7_n166 ) , .ZN( u2_u3_u7_n95 ) );
  NOR2_X1 u2_u3_u7_U71 (.A2( u2_u3_X_45 ) , .A1( u2_u3_X_48 ) , .ZN( u2_u3_u7_n99 ) );
  NOR2_X1 u2_u3_u7_U72 (.A2( u2_u3_X_44 ) , .A1( u2_u3_u7_n167 ) , .ZN( u2_u3_u7_n98 ) );
  NOR2_X1 u2_u3_u7_U73 (.A2( u2_u3_X_46 ) , .A1( u2_u3_X_47 ) , .ZN( u2_u3_u7_n152 ) );
  AND2_X1 u2_u3_u7_U74 (.A1( u2_u3_X_47 ) , .ZN( u2_u3_u7_n156 ) , .A2( u2_u3_u7_n163 ) );
  NAND2_X1 u2_u3_u7_U75 (.A2( u2_u3_X_46 ) , .A1( u2_u3_X_47 ) , .ZN( u2_u3_u7_n125 ) );
  AND2_X1 u2_u3_u7_U76 (.A2( u2_u3_X_45 ) , .A1( u2_u3_X_48 ) , .ZN( u2_u3_u7_n102 ) );
  AND2_X1 u2_u3_u7_U77 (.A2( u2_u3_X_43 ) , .A1( u2_u3_X_44 ) , .ZN( u2_u3_u7_n96 ) );
  AND2_X1 u2_u3_u7_U78 (.A1( u2_u3_X_44 ) , .ZN( u2_u3_u7_n100 ) , .A2( u2_u3_u7_n167 ) );
  AND2_X1 u2_u3_u7_U79 (.A1( u2_u3_X_48 ) , .A2( u2_u3_u7_n166 ) , .ZN( u2_u3_u7_n93 ) );
  OAI222_X1 u2_u3_u7_U8 (.C2( u2_u3_u7_n101 ) , .B2( u2_u3_u7_n111 ) , .A1( u2_u3_u7_n113 ) , .C1( u2_u3_u7_n146 ) , .A2( u2_u3_u7_n162 ) , .B1( u2_u3_u7_n164 ) , .ZN( u2_u3_u7_n94 ) );
  INV_X1 u2_u3_u7_U80 (.A( u2_u3_X_46 ) , .ZN( u2_u3_u7_n163 ) );
  INV_X1 u2_u3_u7_U81 (.A( u2_u3_X_43 ) , .ZN( u2_u3_u7_n167 ) );
  INV_X1 u2_u3_u7_U82 (.A( u2_u3_X_45 ) , .ZN( u2_u3_u7_n166 ) );
  NAND4_X1 u2_u3_u7_U83 (.ZN( u2_out3_5 ) , .A4( u2_u3_u7_n108 ) , .A3( u2_u3_u7_n109 ) , .A1( u2_u3_u7_n116 ) , .A2( u2_u3_u7_n123 ) );
  AOI22_X1 u2_u3_u7_U84 (.ZN( u2_u3_u7_n109 ) , .A2( u2_u3_u7_n126 ) , .B2( u2_u3_u7_n145 ) , .B1( u2_u3_u7_n156 ) , .A1( u2_u3_u7_n171 ) );
  NOR4_X1 u2_u3_u7_U85 (.A4( u2_u3_u7_n104 ) , .A3( u2_u3_u7_n105 ) , .A2( u2_u3_u7_n106 ) , .A1( u2_u3_u7_n107 ) , .ZN( u2_u3_u7_n108 ) );
  NAND4_X1 u2_u3_u7_U86 (.ZN( u2_out3_27 ) , .A4( u2_u3_u7_n118 ) , .A3( u2_u3_u7_n119 ) , .A2( u2_u3_u7_n120 ) , .A1( u2_u3_u7_n121 ) );
  OAI21_X1 u2_u3_u7_U87 (.ZN( u2_u3_u7_n121 ) , .B2( u2_u3_u7_n145 ) , .A( u2_u3_u7_n150 ) , .B1( u2_u3_u7_n174 ) );
  OAI21_X1 u2_u3_u7_U88 (.ZN( u2_u3_u7_n120 ) , .A( u2_u3_u7_n161 ) , .B2( u2_u3_u7_n170 ) , .B1( u2_u3_u7_n179 ) );
  NAND4_X1 u2_u3_u7_U89 (.ZN( u2_out3_21 ) , .A4( u2_u3_u7_n157 ) , .A3( u2_u3_u7_n158 ) , .A2( u2_u3_u7_n159 ) , .A1( u2_u3_u7_n160 ) );
  OAI221_X1 u2_u3_u7_U9 (.C1( u2_u3_u7_n101 ) , .C2( u2_u3_u7_n147 ) , .ZN( u2_u3_u7_n155 ) , .B2( u2_u3_u7_n162 ) , .A( u2_u3_u7_n91 ) , .B1( u2_u3_u7_n92 ) );
  OAI21_X1 u2_u3_u7_U90 (.B1( u2_u3_u7_n145 ) , .ZN( u2_u3_u7_n160 ) , .A( u2_u3_u7_n161 ) , .B2( u2_u3_u7_n177 ) );
  AOI22_X1 u2_u3_u7_U91 (.B2( u2_u3_u7_n149 ) , .B1( u2_u3_u7_n150 ) , .A2( u2_u3_u7_n151 ) , .A1( u2_u3_u7_n152 ) , .ZN( u2_u3_u7_n158 ) );
  NAND4_X1 u2_u3_u7_U92 (.ZN( u2_out3_15 ) , .A4( u2_u3_u7_n142 ) , .A3( u2_u3_u7_n143 ) , .A2( u2_u3_u7_n144 ) , .A1( u2_u3_u7_n178 ) );
  OR2_X1 u2_u3_u7_U93 (.A2( u2_u3_u7_n125 ) , .A1( u2_u3_u7_n129 ) , .ZN( u2_u3_u7_n144 ) );
  AOI22_X1 u2_u3_u7_U94 (.A2( u2_u3_u7_n126 ) , .ZN( u2_u3_u7_n143 ) , .B2( u2_u3_u7_n165 ) , .B1( u2_u3_u7_n173 ) , .A1( u2_u3_u7_n174 ) );
  NAND3_X1 u2_u3_u7_U95 (.A3( u2_u3_u7_n146 ) , .A2( u2_u3_u7_n147 ) , .A1( u2_u3_u7_n148 ) , .ZN( u2_u3_u7_n151 ) );
  NAND3_X1 u2_u3_u7_U96 (.A3( u2_u3_u7_n131 ) , .A2( u2_u3_u7_n132 ) , .A1( u2_u3_u7_n133 ) , .ZN( u2_u3_u7_n135 ) );
  XOR2_X1 u2_u4_U10 (.B( u2_K5_45 ) , .A( u2_R3_30 ) , .Z( u2_u4_X_45 ) );
  XOR2_X1 u2_u4_U11 (.B( u2_K5_44 ) , .A( u2_R3_29 ) , .Z( u2_u4_X_44 ) );
  XOR2_X1 u2_u4_U12 (.B( u2_K5_43 ) , .A( u2_R3_28 ) , .Z( u2_u4_X_43 ) );
  XOR2_X1 u2_u4_U13 (.B( u2_K5_42 ) , .A( u2_R3_29 ) , .Z( u2_u4_X_42 ) );
  XOR2_X1 u2_u4_U14 (.B( u2_K5_41 ) , .A( u2_R3_28 ) , .Z( u2_u4_X_41 ) );
  XOR2_X1 u2_u4_U18 (.B( u2_K5_38 ) , .A( u2_R3_25 ) , .Z( u2_u4_X_38 ) );
  XOR2_X1 u2_u4_U19 (.B( u2_K5_37 ) , .A( u2_R3_24 ) , .Z( u2_u4_X_37 ) );
  XOR2_X1 u2_u4_U2 (.B( u2_K5_8 ) , .A( u2_R3_5 ) , .Z( u2_u4_X_8 ) );
  XOR2_X1 u2_u4_U20 (.B( u2_K5_36 ) , .A( u2_R3_25 ) , .Z( u2_u4_X_36 ) );
  XOR2_X1 u2_u4_U21 (.B( u2_K5_35 ) , .A( u2_R3_24 ) , .Z( u2_u4_X_35 ) );
  XOR2_X1 u2_u4_U23 (.B( u2_K5_33 ) , .A( u2_R3_22 ) , .Z( u2_u4_X_33 ) );
  XOR2_X1 u2_u4_U24 (.B( u2_K5_32 ) , .A( u2_R3_21 ) , .Z( u2_u4_X_32 ) );
  XOR2_X1 u2_u4_U25 (.B( u2_K5_31 ) , .A( u2_R3_20 ) , .Z( u2_u4_X_31 ) );
  XOR2_X1 u2_u4_U26 (.B( u2_K5_30 ) , .A( u2_R3_21 ) , .Z( u2_u4_X_30 ) );
  XOR2_X1 u2_u4_U27 (.B( u2_K5_2 ) , .A( u2_R3_1 ) , .Z( u2_u4_X_2 ) );
  XOR2_X1 u2_u4_U28 (.B( u2_K5_29 ) , .A( u2_R3_20 ) , .Z( u2_u4_X_29 ) );
  XOR2_X1 u2_u4_U3 (.B( u2_K5_7 ) , .A( u2_R3_4 ) , .Z( u2_u4_X_7 ) );
  XOR2_X1 u2_u4_U30 (.B( u2_K5_27 ) , .A( u2_R3_18 ) , .Z( u2_u4_X_27 ) );
  XOR2_X1 u2_u4_U31 (.B( u2_K5_26 ) , .A( u2_R3_17 ) , .Z( u2_u4_X_26 ) );
  XOR2_X1 u2_u4_U32 (.B( u2_K5_25 ) , .A( u2_R3_16 ) , .Z( u2_u4_X_25 ) );
  XOR2_X1 u2_u4_U33 (.B( u2_K5_24 ) , .A( u2_R3_17 ) , .Z( u2_u4_X_24 ) );
  XOR2_X1 u2_u4_U34 (.B( u2_K5_23 ) , .A( u2_R3_16 ) , .Z( u2_u4_X_23 ) );
  XOR2_X1 u2_u4_U37 (.B( u2_K5_20 ) , .A( u2_R3_13 ) , .Z( u2_u4_X_20 ) );
  XOR2_X1 u2_u4_U39 (.B( u2_K5_19 ) , .A( u2_R3_12 ) , .Z( u2_u4_X_19 ) );
  XOR2_X1 u2_u4_U4 (.B( u2_K5_6 ) , .A( u2_R3_5 ) , .Z( u2_u4_X_6 ) );
  XOR2_X1 u2_u4_U40 (.B( u2_K5_18 ) , .A( u2_R3_13 ) , .Z( u2_u4_X_18 ) );
  XOR2_X1 u2_u4_U41 (.B( u2_K5_17 ) , .A( u2_R3_12 ) , .Z( u2_u4_X_17 ) );
  XOR2_X1 u2_u4_U44 (.B( u2_K5_14 ) , .A( u2_R3_9 ) , .Z( u2_u4_X_14 ) );
  XOR2_X1 u2_u4_U45 (.B( u2_K5_13 ) , .A( u2_R3_8 ) , .Z( u2_u4_X_13 ) );
  XOR2_X1 u2_u4_U46 (.B( u2_K5_12 ) , .A( u2_R3_9 ) , .Z( u2_u4_X_12 ) );
  XOR2_X1 u2_u4_U47 (.B( u2_K5_11 ) , .A( u2_R3_8 ) , .Z( u2_u4_X_11 ) );
  XOR2_X1 u2_u4_U5 (.B( u2_K5_5 ) , .A( u2_R3_4 ) , .Z( u2_u4_X_5 ) );
  XOR2_X1 u2_u4_U7 (.B( u2_K5_48 ) , .A( u2_R3_1 ) , .Z( u2_u4_X_48 ) );
  AND3_X1 u2_u4_u0_U10 (.A2( u2_u4_u0_n112 ) , .ZN( u2_u4_u0_n127 ) , .A3( u2_u4_u0_n130 ) , .A1( u2_u4_u0_n148 ) );
  NAND2_X1 u2_u4_u0_U11 (.ZN( u2_u4_u0_n113 ) , .A1( u2_u4_u0_n139 ) , .A2( u2_u4_u0_n149 ) );
  AND2_X1 u2_u4_u0_U12 (.ZN( u2_u4_u0_n107 ) , .A1( u2_u4_u0_n130 ) , .A2( u2_u4_u0_n140 ) );
  AND2_X1 u2_u4_u0_U13 (.A2( u2_u4_u0_n129 ) , .A1( u2_u4_u0_n130 ) , .ZN( u2_u4_u0_n151 ) );
  AND2_X1 u2_u4_u0_U14 (.A1( u2_u4_u0_n108 ) , .A2( u2_u4_u0_n125 ) , .ZN( u2_u4_u0_n145 ) );
  INV_X1 u2_u4_u0_U15 (.A( u2_u4_u0_n143 ) , .ZN( u2_u4_u0_n173 ) );
  NOR2_X1 u2_u4_u0_U16 (.A2( u2_u4_u0_n136 ) , .ZN( u2_u4_u0_n147 ) , .A1( u2_u4_u0_n160 ) );
  NOR2_X1 u2_u4_u0_U17 (.A1( u2_u4_u0_n163 ) , .A2( u2_u4_u0_n164 ) , .ZN( u2_u4_u0_n95 ) );
  AOI21_X1 u2_u4_u0_U18 (.B1( u2_u4_u0_n103 ) , .ZN( u2_u4_u0_n132 ) , .A( u2_u4_u0_n165 ) , .B2( u2_u4_u0_n93 ) );
  INV_X1 u2_u4_u0_U19 (.A( u2_u4_u0_n142 ) , .ZN( u2_u4_u0_n165 ) );
  OAI221_X1 u2_u4_u0_U20 (.C1( u2_u4_u0_n121 ) , .ZN( u2_u4_u0_n122 ) , .B2( u2_u4_u0_n127 ) , .A( u2_u4_u0_n143 ) , .B1( u2_u4_u0_n144 ) , .C2( u2_u4_u0_n147 ) );
  OAI22_X1 u2_u4_u0_U21 (.B1( u2_u4_u0_n125 ) , .ZN( u2_u4_u0_n126 ) , .A1( u2_u4_u0_n138 ) , .A2( u2_u4_u0_n146 ) , .B2( u2_u4_u0_n147 ) );
  OAI22_X1 u2_u4_u0_U22 (.B1( u2_u4_u0_n131 ) , .A1( u2_u4_u0_n144 ) , .B2( u2_u4_u0_n147 ) , .A2( u2_u4_u0_n90 ) , .ZN( u2_u4_u0_n91 ) );
  AND3_X1 u2_u4_u0_U23 (.A3( u2_u4_u0_n121 ) , .A2( u2_u4_u0_n125 ) , .A1( u2_u4_u0_n148 ) , .ZN( u2_u4_u0_n90 ) );
  NAND2_X1 u2_u4_u0_U24 (.A1( u2_u4_u0_n100 ) , .A2( u2_u4_u0_n103 ) , .ZN( u2_u4_u0_n125 ) );
  INV_X1 u2_u4_u0_U25 (.A( u2_u4_u0_n136 ) , .ZN( u2_u4_u0_n161 ) );
  NOR2_X1 u2_u4_u0_U26 (.A1( u2_u4_u0_n120 ) , .ZN( u2_u4_u0_n143 ) , .A2( u2_u4_u0_n167 ) );
  OAI221_X1 u2_u4_u0_U27 (.C1( u2_u4_u0_n112 ) , .ZN( u2_u4_u0_n120 ) , .B1( u2_u4_u0_n138 ) , .B2( u2_u4_u0_n141 ) , .C2( u2_u4_u0_n147 ) , .A( u2_u4_u0_n172 ) );
  AOI211_X1 u2_u4_u0_U28 (.B( u2_u4_u0_n115 ) , .A( u2_u4_u0_n116 ) , .C2( u2_u4_u0_n117 ) , .C1( u2_u4_u0_n118 ) , .ZN( u2_u4_u0_n119 ) );
  AOI22_X1 u2_u4_u0_U29 (.B2( u2_u4_u0_n109 ) , .A2( u2_u4_u0_n110 ) , .ZN( u2_u4_u0_n111 ) , .B1( u2_u4_u0_n118 ) , .A1( u2_u4_u0_n160 ) );
  INV_X1 u2_u4_u0_U3 (.A( u2_u4_u0_n113 ) , .ZN( u2_u4_u0_n166 ) );
  NAND2_X1 u2_u4_u0_U30 (.A1( u2_u4_u0_n100 ) , .ZN( u2_u4_u0_n129 ) , .A2( u2_u4_u0_n95 ) );
  INV_X1 u2_u4_u0_U31 (.A( u2_u4_u0_n118 ) , .ZN( u2_u4_u0_n158 ) );
  AOI21_X1 u2_u4_u0_U32 (.ZN( u2_u4_u0_n104 ) , .B1( u2_u4_u0_n107 ) , .B2( u2_u4_u0_n141 ) , .A( u2_u4_u0_n144 ) );
  AOI21_X1 u2_u4_u0_U33 (.B1( u2_u4_u0_n127 ) , .B2( u2_u4_u0_n129 ) , .A( u2_u4_u0_n138 ) , .ZN( u2_u4_u0_n96 ) );
  AOI21_X1 u2_u4_u0_U34 (.ZN( u2_u4_u0_n116 ) , .B2( u2_u4_u0_n142 ) , .A( u2_u4_u0_n144 ) , .B1( u2_u4_u0_n166 ) );
  NAND2_X1 u2_u4_u0_U35 (.A2( u2_u4_u0_n100 ) , .A1( u2_u4_u0_n101 ) , .ZN( u2_u4_u0_n139 ) );
  NAND2_X1 u2_u4_u0_U36 (.A2( u2_u4_u0_n100 ) , .ZN( u2_u4_u0_n131 ) , .A1( u2_u4_u0_n92 ) );
  NAND2_X1 u2_u4_u0_U37 (.A1( u2_u4_u0_n101 ) , .A2( u2_u4_u0_n102 ) , .ZN( u2_u4_u0_n150 ) );
  INV_X1 u2_u4_u0_U38 (.A( u2_u4_u0_n138 ) , .ZN( u2_u4_u0_n160 ) );
  NAND2_X1 u2_u4_u0_U39 (.A1( u2_u4_u0_n102 ) , .ZN( u2_u4_u0_n128 ) , .A2( u2_u4_u0_n95 ) );
  AOI21_X1 u2_u4_u0_U4 (.B1( u2_u4_u0_n114 ) , .ZN( u2_u4_u0_n115 ) , .B2( u2_u4_u0_n129 ) , .A( u2_u4_u0_n161 ) );
  NAND2_X1 u2_u4_u0_U40 (.ZN( u2_u4_u0_n148 ) , .A1( u2_u4_u0_n93 ) , .A2( u2_u4_u0_n95 ) );
  NAND2_X1 u2_u4_u0_U41 (.A2( u2_u4_u0_n102 ) , .A1( u2_u4_u0_n103 ) , .ZN( u2_u4_u0_n149 ) );
  NAND2_X1 u2_u4_u0_U42 (.A2( u2_u4_u0_n102 ) , .ZN( u2_u4_u0_n114 ) , .A1( u2_u4_u0_n92 ) );
  NAND2_X1 u2_u4_u0_U43 (.A2( u2_u4_u0_n101 ) , .ZN( u2_u4_u0_n121 ) , .A1( u2_u4_u0_n93 ) );
  NAND2_X1 u2_u4_u0_U44 (.ZN( u2_u4_u0_n112 ) , .A2( u2_u4_u0_n92 ) , .A1( u2_u4_u0_n93 ) );
  INV_X1 u2_u4_u0_U45 (.ZN( u2_u4_u0_n172 ) , .A( u2_u4_u0_n88 ) );
  OAI222_X1 u2_u4_u0_U46 (.C1( u2_u4_u0_n108 ) , .A1( u2_u4_u0_n125 ) , .B2( u2_u4_u0_n128 ) , .B1( u2_u4_u0_n144 ) , .A2( u2_u4_u0_n158 ) , .C2( u2_u4_u0_n161 ) , .ZN( u2_u4_u0_n88 ) );
  OR3_X1 u2_u4_u0_U47 (.A3( u2_u4_u0_n152 ) , .A2( u2_u4_u0_n153 ) , .A1( u2_u4_u0_n154 ) , .ZN( u2_u4_u0_n155 ) );
  AOI21_X1 u2_u4_u0_U48 (.B2( u2_u4_u0_n150 ) , .B1( u2_u4_u0_n151 ) , .ZN( u2_u4_u0_n152 ) , .A( u2_u4_u0_n158 ) );
  AOI21_X1 u2_u4_u0_U49 (.A( u2_u4_u0_n144 ) , .B2( u2_u4_u0_n145 ) , .B1( u2_u4_u0_n146 ) , .ZN( u2_u4_u0_n154 ) );
  AOI21_X1 u2_u4_u0_U5 (.B2( u2_u4_u0_n131 ) , .ZN( u2_u4_u0_n134 ) , .B1( u2_u4_u0_n151 ) , .A( u2_u4_u0_n158 ) );
  AOI21_X1 u2_u4_u0_U50 (.A( u2_u4_u0_n147 ) , .B2( u2_u4_u0_n148 ) , .B1( u2_u4_u0_n149 ) , .ZN( u2_u4_u0_n153 ) );
  INV_X1 u2_u4_u0_U51 (.ZN( u2_u4_u0_n171 ) , .A( u2_u4_u0_n99 ) );
  OAI211_X1 u2_u4_u0_U52 (.C2( u2_u4_u0_n140 ) , .C1( u2_u4_u0_n161 ) , .A( u2_u4_u0_n169 ) , .B( u2_u4_u0_n98 ) , .ZN( u2_u4_u0_n99 ) );
  AOI211_X1 u2_u4_u0_U53 (.C1( u2_u4_u0_n118 ) , .A( u2_u4_u0_n123 ) , .B( u2_u4_u0_n96 ) , .C2( u2_u4_u0_n97 ) , .ZN( u2_u4_u0_n98 ) );
  INV_X1 u2_u4_u0_U54 (.ZN( u2_u4_u0_n169 ) , .A( u2_u4_u0_n91 ) );
  NOR2_X1 u2_u4_u0_U55 (.A2( u2_u4_X_4 ) , .A1( u2_u4_X_5 ) , .ZN( u2_u4_u0_n118 ) );
  NOR2_X1 u2_u4_u0_U56 (.A2( u2_u4_X_2 ) , .ZN( u2_u4_u0_n103 ) , .A1( u2_u4_u0_n164 ) );
  NOR2_X1 u2_u4_u0_U57 (.A2( u2_u4_X_1 ) , .A1( u2_u4_X_2 ) , .ZN( u2_u4_u0_n92 ) );
  NOR2_X1 u2_u4_u0_U58 (.A2( u2_u4_X_1 ) , .ZN( u2_u4_u0_n101 ) , .A1( u2_u4_u0_n163 ) );
  NAND2_X1 u2_u4_u0_U59 (.A2( u2_u4_X_4 ) , .A1( u2_u4_X_5 ) , .ZN( u2_u4_u0_n144 ) );
  NOR2_X1 u2_u4_u0_U6 (.A1( u2_u4_u0_n108 ) , .ZN( u2_u4_u0_n123 ) , .A2( u2_u4_u0_n158 ) );
  NOR2_X1 u2_u4_u0_U60 (.A2( u2_u4_X_5 ) , .ZN( u2_u4_u0_n136 ) , .A1( u2_u4_u0_n159 ) );
  NAND2_X1 u2_u4_u0_U61 (.A1( u2_u4_X_5 ) , .ZN( u2_u4_u0_n138 ) , .A2( u2_u4_u0_n159 ) );
  AND2_X1 u2_u4_u0_U62 (.A2( u2_u4_X_3 ) , .A1( u2_u4_X_6 ) , .ZN( u2_u4_u0_n102 ) );
  INV_X1 u2_u4_u0_U63 (.A( u2_u4_X_4 ) , .ZN( u2_u4_u0_n159 ) );
  INV_X1 u2_u4_u0_U64 (.A( u2_u4_X_1 ) , .ZN( u2_u4_u0_n164 ) );
  INV_X1 u2_u4_u0_U65 (.A( u2_u4_X_2 ) , .ZN( u2_u4_u0_n163 ) );
  INV_X1 u2_u4_u0_U66 (.A( u2_u4_X_3 ) , .ZN( u2_u4_u0_n162 ) );
  AOI211_X1 u2_u4_u0_U67 (.B( u2_u4_u0_n133 ) , .A( u2_u4_u0_n134 ) , .C2( u2_u4_u0_n135 ) , .C1( u2_u4_u0_n136 ) , .ZN( u2_u4_u0_n137 ) );
  INV_X1 u2_u4_u0_U68 (.A( u2_u4_u0_n126 ) , .ZN( u2_u4_u0_n168 ) );
  INV_X1 u2_u4_u0_U69 (.ZN( u2_u4_u0_n174 ) , .A( u2_u4_u0_n89 ) );
  OAI21_X1 u2_u4_u0_U7 (.B1( u2_u4_u0_n150 ) , .B2( u2_u4_u0_n158 ) , .A( u2_u4_u0_n172 ) , .ZN( u2_u4_u0_n89 ) );
  AOI211_X1 u2_u4_u0_U70 (.B( u2_u4_u0_n104 ) , .A( u2_u4_u0_n105 ) , .ZN( u2_u4_u0_n106 ) , .C2( u2_u4_u0_n113 ) , .C1( u2_u4_u0_n160 ) );
  OR4_X1 u2_u4_u0_U71 (.ZN( u2_out4_31 ) , .A4( u2_u4_u0_n155 ) , .A2( u2_u4_u0_n156 ) , .A1( u2_u4_u0_n157 ) , .A3( u2_u4_u0_n173 ) );
  AOI21_X1 u2_u4_u0_U72 (.A( u2_u4_u0_n138 ) , .B2( u2_u4_u0_n139 ) , .B1( u2_u4_u0_n140 ) , .ZN( u2_u4_u0_n157 ) );
  AOI21_X1 u2_u4_u0_U73 (.B2( u2_u4_u0_n141 ) , .B1( u2_u4_u0_n142 ) , .ZN( u2_u4_u0_n156 ) , .A( u2_u4_u0_n161 ) );
  OR4_X1 u2_u4_u0_U74 (.ZN( u2_out4_17 ) , .A4( u2_u4_u0_n122 ) , .A2( u2_u4_u0_n123 ) , .A1( u2_u4_u0_n124 ) , .A3( u2_u4_u0_n170 ) );
  AOI21_X1 u2_u4_u0_U75 (.B2( u2_u4_u0_n107 ) , .ZN( u2_u4_u0_n124 ) , .B1( u2_u4_u0_n128 ) , .A( u2_u4_u0_n161 ) );
  INV_X1 u2_u4_u0_U76 (.A( u2_u4_u0_n111 ) , .ZN( u2_u4_u0_n170 ) );
  AOI21_X1 u2_u4_u0_U77 (.B1( u2_u4_u0_n132 ) , .ZN( u2_u4_u0_n133 ) , .A( u2_u4_u0_n144 ) , .B2( u2_u4_u0_n166 ) );
  OAI22_X1 u2_u4_u0_U78 (.ZN( u2_u4_u0_n105 ) , .A2( u2_u4_u0_n132 ) , .B1( u2_u4_u0_n146 ) , .A1( u2_u4_u0_n147 ) , .B2( u2_u4_u0_n161 ) );
  NAND2_X1 u2_u4_u0_U79 (.ZN( u2_u4_u0_n110 ) , .A2( u2_u4_u0_n132 ) , .A1( u2_u4_u0_n145 ) );
  AND2_X1 u2_u4_u0_U8 (.A1( u2_u4_u0_n114 ) , .A2( u2_u4_u0_n121 ) , .ZN( u2_u4_u0_n146 ) );
  INV_X1 u2_u4_u0_U80 (.A( u2_u4_u0_n119 ) , .ZN( u2_u4_u0_n167 ) );
  NAND2_X1 u2_u4_u0_U81 (.A2( u2_u4_u0_n103 ) , .ZN( u2_u4_u0_n140 ) , .A1( u2_u4_u0_n94 ) );
  NAND2_X1 u2_u4_u0_U82 (.A1( u2_u4_u0_n101 ) , .ZN( u2_u4_u0_n130 ) , .A2( u2_u4_u0_n94 ) );
  NAND2_X1 u2_u4_u0_U83 (.ZN( u2_u4_u0_n108 ) , .A1( u2_u4_u0_n92 ) , .A2( u2_u4_u0_n94 ) );
  AND2_X1 u2_u4_u0_U84 (.A1( u2_u4_X_6 ) , .A2( u2_u4_u0_n162 ) , .ZN( u2_u4_u0_n93 ) );
  NAND2_X1 u2_u4_u0_U85 (.ZN( u2_u4_u0_n142 ) , .A1( u2_u4_u0_n94 ) , .A2( u2_u4_u0_n95 ) );
  NOR2_X1 u2_u4_u0_U86 (.A2( u2_u4_X_6 ) , .ZN( u2_u4_u0_n100 ) , .A1( u2_u4_u0_n162 ) );
  NOR2_X1 u2_u4_u0_U87 (.A2( u2_u4_X_3 ) , .A1( u2_u4_X_6 ) , .ZN( u2_u4_u0_n94 ) );
  NAND3_X1 u2_u4_u0_U88 (.ZN( u2_out4_23 ) , .A3( u2_u4_u0_n137 ) , .A1( u2_u4_u0_n168 ) , .A2( u2_u4_u0_n171 ) );
  NAND3_X1 u2_u4_u0_U89 (.A3( u2_u4_u0_n127 ) , .A2( u2_u4_u0_n128 ) , .ZN( u2_u4_u0_n135 ) , .A1( u2_u4_u0_n150 ) );
  AND2_X1 u2_u4_u0_U9 (.A1( u2_u4_u0_n131 ) , .ZN( u2_u4_u0_n141 ) , .A2( u2_u4_u0_n150 ) );
  NAND3_X1 u2_u4_u0_U90 (.ZN( u2_u4_u0_n117 ) , .A3( u2_u4_u0_n132 ) , .A2( u2_u4_u0_n139 ) , .A1( u2_u4_u0_n148 ) );
  NAND3_X1 u2_u4_u0_U91 (.ZN( u2_u4_u0_n109 ) , .A2( u2_u4_u0_n114 ) , .A3( u2_u4_u0_n140 ) , .A1( u2_u4_u0_n149 ) );
  NAND3_X1 u2_u4_u0_U92 (.ZN( u2_out4_9 ) , .A3( u2_u4_u0_n106 ) , .A2( u2_u4_u0_n171 ) , .A1( u2_u4_u0_n174 ) );
  NAND3_X1 u2_u4_u0_U93 (.A2( u2_u4_u0_n128 ) , .A1( u2_u4_u0_n132 ) , .A3( u2_u4_u0_n146 ) , .ZN( u2_u4_u0_n97 ) );
  NOR2_X1 u2_u4_u1_U10 (.A1( u2_u4_u1_n112 ) , .A2( u2_u4_u1_n116 ) , .ZN( u2_u4_u1_n118 ) );
  NAND3_X1 u2_u4_u1_U100 (.ZN( u2_u4_u1_n113 ) , .A1( u2_u4_u1_n120 ) , .A3( u2_u4_u1_n133 ) , .A2( u2_u4_u1_n155 ) );
  OAI21_X1 u2_u4_u1_U11 (.ZN( u2_u4_u1_n101 ) , .B1( u2_u4_u1_n141 ) , .A( u2_u4_u1_n146 ) , .B2( u2_u4_u1_n183 ) );
  AOI21_X1 u2_u4_u1_U12 (.B2( u2_u4_u1_n155 ) , .B1( u2_u4_u1_n156 ) , .ZN( u2_u4_u1_n157 ) , .A( u2_u4_u1_n174 ) );
  NAND2_X1 u2_u4_u1_U13 (.ZN( u2_u4_u1_n140 ) , .A2( u2_u4_u1_n150 ) , .A1( u2_u4_u1_n155 ) );
  NAND2_X1 u2_u4_u1_U14 (.A1( u2_u4_u1_n131 ) , .ZN( u2_u4_u1_n147 ) , .A2( u2_u4_u1_n153 ) );
  INV_X1 u2_u4_u1_U15 (.A( u2_u4_u1_n139 ) , .ZN( u2_u4_u1_n174 ) );
  OR4_X1 u2_u4_u1_U16 (.A4( u2_u4_u1_n106 ) , .A3( u2_u4_u1_n107 ) , .ZN( u2_u4_u1_n108 ) , .A1( u2_u4_u1_n117 ) , .A2( u2_u4_u1_n184 ) );
  AOI21_X1 u2_u4_u1_U17 (.ZN( u2_u4_u1_n106 ) , .A( u2_u4_u1_n112 ) , .B1( u2_u4_u1_n154 ) , .B2( u2_u4_u1_n156 ) );
  AOI21_X1 u2_u4_u1_U18 (.ZN( u2_u4_u1_n107 ) , .B1( u2_u4_u1_n134 ) , .B2( u2_u4_u1_n149 ) , .A( u2_u4_u1_n174 ) );
  INV_X1 u2_u4_u1_U19 (.A( u2_u4_u1_n101 ) , .ZN( u2_u4_u1_n184 ) );
  INV_X1 u2_u4_u1_U20 (.A( u2_u4_u1_n112 ) , .ZN( u2_u4_u1_n171 ) );
  NAND2_X1 u2_u4_u1_U21 (.ZN( u2_u4_u1_n141 ) , .A1( u2_u4_u1_n153 ) , .A2( u2_u4_u1_n156 ) );
  AND2_X1 u2_u4_u1_U22 (.A1( u2_u4_u1_n123 ) , .ZN( u2_u4_u1_n134 ) , .A2( u2_u4_u1_n161 ) );
  NAND2_X1 u2_u4_u1_U23 (.A2( u2_u4_u1_n115 ) , .A1( u2_u4_u1_n116 ) , .ZN( u2_u4_u1_n148 ) );
  NAND2_X1 u2_u4_u1_U24 (.A2( u2_u4_u1_n133 ) , .A1( u2_u4_u1_n135 ) , .ZN( u2_u4_u1_n159 ) );
  NAND2_X1 u2_u4_u1_U25 (.A2( u2_u4_u1_n115 ) , .A1( u2_u4_u1_n120 ) , .ZN( u2_u4_u1_n132 ) );
  INV_X1 u2_u4_u1_U26 (.A( u2_u4_u1_n154 ) , .ZN( u2_u4_u1_n178 ) );
  INV_X1 u2_u4_u1_U27 (.A( u2_u4_u1_n151 ) , .ZN( u2_u4_u1_n183 ) );
  AND2_X1 u2_u4_u1_U28 (.A1( u2_u4_u1_n129 ) , .A2( u2_u4_u1_n133 ) , .ZN( u2_u4_u1_n149 ) );
  INV_X1 u2_u4_u1_U29 (.A( u2_u4_u1_n131 ) , .ZN( u2_u4_u1_n180 ) );
  INV_X1 u2_u4_u1_U3 (.A( u2_u4_u1_n159 ) , .ZN( u2_u4_u1_n182 ) );
  OAI221_X1 u2_u4_u1_U30 (.A( u2_u4_u1_n119 ) , .C2( u2_u4_u1_n129 ) , .ZN( u2_u4_u1_n138 ) , .B2( u2_u4_u1_n152 ) , .C1( u2_u4_u1_n174 ) , .B1( u2_u4_u1_n187 ) );
  INV_X1 u2_u4_u1_U31 (.A( u2_u4_u1_n148 ) , .ZN( u2_u4_u1_n187 ) );
  AOI211_X1 u2_u4_u1_U32 (.B( u2_u4_u1_n117 ) , .A( u2_u4_u1_n118 ) , .ZN( u2_u4_u1_n119 ) , .C2( u2_u4_u1_n146 ) , .C1( u2_u4_u1_n159 ) );
  NOR2_X1 u2_u4_u1_U33 (.A1( u2_u4_u1_n168 ) , .A2( u2_u4_u1_n176 ) , .ZN( u2_u4_u1_n98 ) );
  AOI211_X1 u2_u4_u1_U34 (.B( u2_u4_u1_n162 ) , .A( u2_u4_u1_n163 ) , .C2( u2_u4_u1_n164 ) , .ZN( u2_u4_u1_n165 ) , .C1( u2_u4_u1_n171 ) );
  AOI21_X1 u2_u4_u1_U35 (.A( u2_u4_u1_n160 ) , .B2( u2_u4_u1_n161 ) , .ZN( u2_u4_u1_n162 ) , .B1( u2_u4_u1_n182 ) );
  OR2_X1 u2_u4_u1_U36 (.A2( u2_u4_u1_n157 ) , .A1( u2_u4_u1_n158 ) , .ZN( u2_u4_u1_n163 ) );
  NAND2_X1 u2_u4_u1_U37 (.A1( u2_u4_u1_n128 ) , .ZN( u2_u4_u1_n146 ) , .A2( u2_u4_u1_n160 ) );
  NAND2_X1 u2_u4_u1_U38 (.A2( u2_u4_u1_n112 ) , .ZN( u2_u4_u1_n139 ) , .A1( u2_u4_u1_n152 ) );
  NAND2_X1 u2_u4_u1_U39 (.A1( u2_u4_u1_n105 ) , .ZN( u2_u4_u1_n156 ) , .A2( u2_u4_u1_n99 ) );
  AOI221_X1 u2_u4_u1_U4 (.A( u2_u4_u1_n138 ) , .C2( u2_u4_u1_n139 ) , .C1( u2_u4_u1_n140 ) , .B2( u2_u4_u1_n141 ) , .ZN( u2_u4_u1_n142 ) , .B1( u2_u4_u1_n175 ) );
  AOI221_X1 u2_u4_u1_U40 (.B1( u2_u4_u1_n140 ) , .ZN( u2_u4_u1_n167 ) , .B2( u2_u4_u1_n172 ) , .C2( u2_u4_u1_n175 ) , .C1( u2_u4_u1_n178 ) , .A( u2_u4_u1_n188 ) );
  INV_X1 u2_u4_u1_U41 (.ZN( u2_u4_u1_n188 ) , .A( u2_u4_u1_n97 ) );
  AOI211_X1 u2_u4_u1_U42 (.A( u2_u4_u1_n118 ) , .C1( u2_u4_u1_n132 ) , .C2( u2_u4_u1_n139 ) , .B( u2_u4_u1_n96 ) , .ZN( u2_u4_u1_n97 ) );
  AOI21_X1 u2_u4_u1_U43 (.B2( u2_u4_u1_n121 ) , .B1( u2_u4_u1_n135 ) , .A( u2_u4_u1_n152 ) , .ZN( u2_u4_u1_n96 ) );
  NOR2_X1 u2_u4_u1_U44 (.ZN( u2_u4_u1_n117 ) , .A1( u2_u4_u1_n121 ) , .A2( u2_u4_u1_n160 ) );
  OAI21_X1 u2_u4_u1_U45 (.B2( u2_u4_u1_n123 ) , .ZN( u2_u4_u1_n145 ) , .B1( u2_u4_u1_n160 ) , .A( u2_u4_u1_n185 ) );
  INV_X1 u2_u4_u1_U46 (.A( u2_u4_u1_n122 ) , .ZN( u2_u4_u1_n185 ) );
  AOI21_X1 u2_u4_u1_U47 (.B2( u2_u4_u1_n120 ) , .B1( u2_u4_u1_n121 ) , .ZN( u2_u4_u1_n122 ) , .A( u2_u4_u1_n128 ) );
  AOI21_X1 u2_u4_u1_U48 (.A( u2_u4_u1_n128 ) , .B2( u2_u4_u1_n129 ) , .ZN( u2_u4_u1_n130 ) , .B1( u2_u4_u1_n150 ) );
  NAND2_X1 u2_u4_u1_U49 (.ZN( u2_u4_u1_n112 ) , .A1( u2_u4_u1_n169 ) , .A2( u2_u4_u1_n170 ) );
  AOI211_X1 u2_u4_u1_U5 (.ZN( u2_u4_u1_n124 ) , .A( u2_u4_u1_n138 ) , .C2( u2_u4_u1_n139 ) , .B( u2_u4_u1_n145 ) , .C1( u2_u4_u1_n147 ) );
  NAND2_X1 u2_u4_u1_U50 (.ZN( u2_u4_u1_n129 ) , .A2( u2_u4_u1_n95 ) , .A1( u2_u4_u1_n98 ) );
  NAND2_X1 u2_u4_u1_U51 (.A1( u2_u4_u1_n102 ) , .ZN( u2_u4_u1_n154 ) , .A2( u2_u4_u1_n99 ) );
  NAND2_X1 u2_u4_u1_U52 (.A2( u2_u4_u1_n100 ) , .ZN( u2_u4_u1_n135 ) , .A1( u2_u4_u1_n99 ) );
  AOI21_X1 u2_u4_u1_U53 (.A( u2_u4_u1_n152 ) , .B2( u2_u4_u1_n153 ) , .B1( u2_u4_u1_n154 ) , .ZN( u2_u4_u1_n158 ) );
  INV_X1 u2_u4_u1_U54 (.A( u2_u4_u1_n160 ) , .ZN( u2_u4_u1_n175 ) );
  NAND2_X1 u2_u4_u1_U55 (.A1( u2_u4_u1_n100 ) , .ZN( u2_u4_u1_n116 ) , .A2( u2_u4_u1_n95 ) );
  NAND2_X1 u2_u4_u1_U56 (.A1( u2_u4_u1_n102 ) , .ZN( u2_u4_u1_n131 ) , .A2( u2_u4_u1_n95 ) );
  NAND2_X1 u2_u4_u1_U57 (.A2( u2_u4_u1_n104 ) , .ZN( u2_u4_u1_n121 ) , .A1( u2_u4_u1_n98 ) );
  NAND2_X1 u2_u4_u1_U58 (.A1( u2_u4_u1_n103 ) , .ZN( u2_u4_u1_n153 ) , .A2( u2_u4_u1_n98 ) );
  NAND2_X1 u2_u4_u1_U59 (.A2( u2_u4_u1_n104 ) , .A1( u2_u4_u1_n105 ) , .ZN( u2_u4_u1_n133 ) );
  AOI22_X1 u2_u4_u1_U6 (.B2( u2_u4_u1_n113 ) , .A2( u2_u4_u1_n114 ) , .ZN( u2_u4_u1_n125 ) , .A1( u2_u4_u1_n171 ) , .B1( u2_u4_u1_n173 ) );
  NAND2_X1 u2_u4_u1_U60 (.ZN( u2_u4_u1_n150 ) , .A2( u2_u4_u1_n98 ) , .A1( u2_u4_u1_n99 ) );
  NAND2_X1 u2_u4_u1_U61 (.A1( u2_u4_u1_n105 ) , .ZN( u2_u4_u1_n155 ) , .A2( u2_u4_u1_n95 ) );
  OAI21_X1 u2_u4_u1_U62 (.ZN( u2_u4_u1_n109 ) , .B1( u2_u4_u1_n129 ) , .B2( u2_u4_u1_n160 ) , .A( u2_u4_u1_n167 ) );
  NAND2_X1 u2_u4_u1_U63 (.A2( u2_u4_u1_n100 ) , .A1( u2_u4_u1_n103 ) , .ZN( u2_u4_u1_n120 ) );
  NAND2_X1 u2_u4_u1_U64 (.A1( u2_u4_u1_n102 ) , .A2( u2_u4_u1_n104 ) , .ZN( u2_u4_u1_n115 ) );
  NAND2_X1 u2_u4_u1_U65 (.A2( u2_u4_u1_n100 ) , .A1( u2_u4_u1_n104 ) , .ZN( u2_u4_u1_n151 ) );
  NAND2_X1 u2_u4_u1_U66 (.A2( u2_u4_u1_n103 ) , .A1( u2_u4_u1_n105 ) , .ZN( u2_u4_u1_n161 ) );
  INV_X1 u2_u4_u1_U67 (.A( u2_u4_u1_n152 ) , .ZN( u2_u4_u1_n173 ) );
  INV_X1 u2_u4_u1_U68 (.A( u2_u4_u1_n128 ) , .ZN( u2_u4_u1_n172 ) );
  NAND2_X1 u2_u4_u1_U69 (.A2( u2_u4_u1_n102 ) , .A1( u2_u4_u1_n103 ) , .ZN( u2_u4_u1_n123 ) );
  NAND2_X1 u2_u4_u1_U7 (.ZN( u2_u4_u1_n114 ) , .A1( u2_u4_u1_n134 ) , .A2( u2_u4_u1_n156 ) );
  NOR2_X1 u2_u4_u1_U70 (.A2( u2_u4_X_7 ) , .A1( u2_u4_X_8 ) , .ZN( u2_u4_u1_n95 ) );
  NOR2_X1 u2_u4_u1_U71 (.A1( u2_u4_X_12 ) , .A2( u2_u4_X_9 ) , .ZN( u2_u4_u1_n100 ) );
  NOR2_X1 u2_u4_u1_U72 (.A2( u2_u4_X_8 ) , .A1( u2_u4_u1_n177 ) , .ZN( u2_u4_u1_n99 ) );
  NOR2_X1 u2_u4_u1_U73 (.A2( u2_u4_X_12 ) , .ZN( u2_u4_u1_n102 ) , .A1( u2_u4_u1_n176 ) );
  NOR2_X1 u2_u4_u1_U74 (.A2( u2_u4_X_9 ) , .ZN( u2_u4_u1_n105 ) , .A1( u2_u4_u1_n168 ) );
  NAND2_X1 u2_u4_u1_U75 (.A1( u2_u4_X_10 ) , .ZN( u2_u4_u1_n160 ) , .A2( u2_u4_u1_n169 ) );
  NAND2_X1 u2_u4_u1_U76 (.A2( u2_u4_X_10 ) , .A1( u2_u4_X_11 ) , .ZN( u2_u4_u1_n152 ) );
  NAND2_X1 u2_u4_u1_U77 (.A1( u2_u4_X_11 ) , .ZN( u2_u4_u1_n128 ) , .A2( u2_u4_u1_n170 ) );
  AND2_X1 u2_u4_u1_U78 (.A2( u2_u4_X_7 ) , .A1( u2_u4_X_8 ) , .ZN( u2_u4_u1_n104 ) );
  AND2_X1 u2_u4_u1_U79 (.A1( u2_u4_X_8 ) , .ZN( u2_u4_u1_n103 ) , .A2( u2_u4_u1_n177 ) );
  AOI22_X1 u2_u4_u1_U8 (.B2( u2_u4_u1_n136 ) , .A2( u2_u4_u1_n137 ) , .ZN( u2_u4_u1_n143 ) , .A1( u2_u4_u1_n171 ) , .B1( u2_u4_u1_n173 ) );
  INV_X1 u2_u4_u1_U80 (.A( u2_u4_X_10 ) , .ZN( u2_u4_u1_n170 ) );
  INV_X1 u2_u4_u1_U81 (.A( u2_u4_X_9 ) , .ZN( u2_u4_u1_n176 ) );
  INV_X1 u2_u4_u1_U82 (.A( u2_u4_X_11 ) , .ZN( u2_u4_u1_n169 ) );
  INV_X1 u2_u4_u1_U83 (.A( u2_u4_X_12 ) , .ZN( u2_u4_u1_n168 ) );
  INV_X1 u2_u4_u1_U84 (.A( u2_u4_X_7 ) , .ZN( u2_u4_u1_n177 ) );
  NAND4_X1 u2_u4_u1_U85 (.ZN( u2_out4_28 ) , .A4( u2_u4_u1_n124 ) , .A3( u2_u4_u1_n125 ) , .A2( u2_u4_u1_n126 ) , .A1( u2_u4_u1_n127 ) );
  OAI21_X1 u2_u4_u1_U86 (.ZN( u2_u4_u1_n127 ) , .B2( u2_u4_u1_n139 ) , .B1( u2_u4_u1_n175 ) , .A( u2_u4_u1_n183 ) );
  OAI21_X1 u2_u4_u1_U87 (.ZN( u2_u4_u1_n126 ) , .B2( u2_u4_u1_n140 ) , .A( u2_u4_u1_n146 ) , .B1( u2_u4_u1_n178 ) );
  NAND4_X1 u2_u4_u1_U88 (.ZN( u2_out4_18 ) , .A4( u2_u4_u1_n165 ) , .A3( u2_u4_u1_n166 ) , .A1( u2_u4_u1_n167 ) , .A2( u2_u4_u1_n186 ) );
  AOI22_X1 u2_u4_u1_U89 (.B2( u2_u4_u1_n146 ) , .B1( u2_u4_u1_n147 ) , .A2( u2_u4_u1_n148 ) , .ZN( u2_u4_u1_n166 ) , .A1( u2_u4_u1_n172 ) );
  INV_X1 u2_u4_u1_U9 (.A( u2_u4_u1_n147 ) , .ZN( u2_u4_u1_n181 ) );
  INV_X1 u2_u4_u1_U90 (.A( u2_u4_u1_n145 ) , .ZN( u2_u4_u1_n186 ) );
  NAND4_X1 u2_u4_u1_U91 (.ZN( u2_out4_2 ) , .A4( u2_u4_u1_n142 ) , .A3( u2_u4_u1_n143 ) , .A2( u2_u4_u1_n144 ) , .A1( u2_u4_u1_n179 ) );
  OAI21_X1 u2_u4_u1_U92 (.B2( u2_u4_u1_n132 ) , .ZN( u2_u4_u1_n144 ) , .A( u2_u4_u1_n146 ) , .B1( u2_u4_u1_n180 ) );
  INV_X1 u2_u4_u1_U93 (.A( u2_u4_u1_n130 ) , .ZN( u2_u4_u1_n179 ) );
  OR4_X1 u2_u4_u1_U94 (.ZN( u2_out4_13 ) , .A4( u2_u4_u1_n108 ) , .A3( u2_u4_u1_n109 ) , .A2( u2_u4_u1_n110 ) , .A1( u2_u4_u1_n111 ) );
  AOI21_X1 u2_u4_u1_U95 (.ZN( u2_u4_u1_n111 ) , .A( u2_u4_u1_n128 ) , .B2( u2_u4_u1_n131 ) , .B1( u2_u4_u1_n135 ) );
  AOI21_X1 u2_u4_u1_U96 (.ZN( u2_u4_u1_n110 ) , .A( u2_u4_u1_n116 ) , .B1( u2_u4_u1_n152 ) , .B2( u2_u4_u1_n160 ) );
  NAND3_X1 u2_u4_u1_U97 (.A3( u2_u4_u1_n149 ) , .A2( u2_u4_u1_n150 ) , .A1( u2_u4_u1_n151 ) , .ZN( u2_u4_u1_n164 ) );
  NAND3_X1 u2_u4_u1_U98 (.A3( u2_u4_u1_n134 ) , .A2( u2_u4_u1_n135 ) , .ZN( u2_u4_u1_n136 ) , .A1( u2_u4_u1_n151 ) );
  NAND3_X1 u2_u4_u1_U99 (.A1( u2_u4_u1_n133 ) , .ZN( u2_u4_u1_n137 ) , .A2( u2_u4_u1_n154 ) , .A3( u2_u4_u1_n181 ) );
  OAI22_X1 u2_u4_u2_U10 (.ZN( u2_u4_u2_n109 ) , .A2( u2_u4_u2_n113 ) , .B2( u2_u4_u2_n133 ) , .B1( u2_u4_u2_n167 ) , .A1( u2_u4_u2_n168 ) );
  NAND3_X1 u2_u4_u2_U100 (.A2( u2_u4_u2_n100 ) , .A1( u2_u4_u2_n104 ) , .A3( u2_u4_u2_n138 ) , .ZN( u2_u4_u2_n98 ) );
  OAI22_X1 u2_u4_u2_U11 (.B1( u2_u4_u2_n151 ) , .A2( u2_u4_u2_n152 ) , .A1( u2_u4_u2_n153 ) , .ZN( u2_u4_u2_n160 ) , .B2( u2_u4_u2_n168 ) );
  NOR3_X1 u2_u4_u2_U12 (.A1( u2_u4_u2_n150 ) , .ZN( u2_u4_u2_n151 ) , .A3( u2_u4_u2_n175 ) , .A2( u2_u4_u2_n188 ) );
  AOI21_X1 u2_u4_u2_U13 (.ZN( u2_u4_u2_n144 ) , .B2( u2_u4_u2_n155 ) , .A( u2_u4_u2_n172 ) , .B1( u2_u4_u2_n185 ) );
  AOI21_X1 u2_u4_u2_U14 (.B2( u2_u4_u2_n143 ) , .ZN( u2_u4_u2_n145 ) , .B1( u2_u4_u2_n152 ) , .A( u2_u4_u2_n171 ) );
  AOI21_X1 u2_u4_u2_U15 (.B2( u2_u4_u2_n120 ) , .B1( u2_u4_u2_n121 ) , .ZN( u2_u4_u2_n126 ) , .A( u2_u4_u2_n167 ) );
  INV_X1 u2_u4_u2_U16 (.A( u2_u4_u2_n156 ) , .ZN( u2_u4_u2_n171 ) );
  INV_X1 u2_u4_u2_U17 (.A( u2_u4_u2_n120 ) , .ZN( u2_u4_u2_n188 ) );
  NAND2_X1 u2_u4_u2_U18 (.A2( u2_u4_u2_n122 ) , .ZN( u2_u4_u2_n150 ) , .A1( u2_u4_u2_n152 ) );
  INV_X1 u2_u4_u2_U19 (.A( u2_u4_u2_n153 ) , .ZN( u2_u4_u2_n170 ) );
  INV_X1 u2_u4_u2_U20 (.A( u2_u4_u2_n137 ) , .ZN( u2_u4_u2_n173 ) );
  NAND2_X1 u2_u4_u2_U21 (.A1( u2_u4_u2_n132 ) , .A2( u2_u4_u2_n139 ) , .ZN( u2_u4_u2_n157 ) );
  INV_X1 u2_u4_u2_U22 (.A( u2_u4_u2_n113 ) , .ZN( u2_u4_u2_n178 ) );
  INV_X1 u2_u4_u2_U23 (.A( u2_u4_u2_n139 ) , .ZN( u2_u4_u2_n175 ) );
  INV_X1 u2_u4_u2_U24 (.A( u2_u4_u2_n155 ) , .ZN( u2_u4_u2_n181 ) );
  INV_X1 u2_u4_u2_U25 (.A( u2_u4_u2_n119 ) , .ZN( u2_u4_u2_n177 ) );
  INV_X1 u2_u4_u2_U26 (.A( u2_u4_u2_n116 ) , .ZN( u2_u4_u2_n180 ) );
  INV_X1 u2_u4_u2_U27 (.A( u2_u4_u2_n131 ) , .ZN( u2_u4_u2_n179 ) );
  INV_X1 u2_u4_u2_U28 (.A( u2_u4_u2_n154 ) , .ZN( u2_u4_u2_n176 ) );
  NAND2_X1 u2_u4_u2_U29 (.A2( u2_u4_u2_n116 ) , .A1( u2_u4_u2_n117 ) , .ZN( u2_u4_u2_n118 ) );
  NOR2_X1 u2_u4_u2_U3 (.ZN( u2_u4_u2_n121 ) , .A2( u2_u4_u2_n177 ) , .A1( u2_u4_u2_n180 ) );
  INV_X1 u2_u4_u2_U30 (.A( u2_u4_u2_n132 ) , .ZN( u2_u4_u2_n182 ) );
  INV_X1 u2_u4_u2_U31 (.A( u2_u4_u2_n158 ) , .ZN( u2_u4_u2_n183 ) );
  OAI21_X1 u2_u4_u2_U32 (.A( u2_u4_u2_n156 ) , .B1( u2_u4_u2_n157 ) , .ZN( u2_u4_u2_n158 ) , .B2( u2_u4_u2_n179 ) );
  NOR2_X1 u2_u4_u2_U33 (.ZN( u2_u4_u2_n156 ) , .A1( u2_u4_u2_n166 ) , .A2( u2_u4_u2_n169 ) );
  NOR2_X1 u2_u4_u2_U34 (.A2( u2_u4_u2_n114 ) , .ZN( u2_u4_u2_n137 ) , .A1( u2_u4_u2_n140 ) );
  NOR2_X1 u2_u4_u2_U35 (.A2( u2_u4_u2_n138 ) , .ZN( u2_u4_u2_n153 ) , .A1( u2_u4_u2_n156 ) );
  AOI211_X1 u2_u4_u2_U36 (.ZN( u2_u4_u2_n130 ) , .C1( u2_u4_u2_n138 ) , .C2( u2_u4_u2_n179 ) , .B( u2_u4_u2_n96 ) , .A( u2_u4_u2_n97 ) );
  OAI22_X1 u2_u4_u2_U37 (.B1( u2_u4_u2_n133 ) , .A2( u2_u4_u2_n137 ) , .A1( u2_u4_u2_n152 ) , .B2( u2_u4_u2_n168 ) , .ZN( u2_u4_u2_n97 ) );
  OAI221_X1 u2_u4_u2_U38 (.B1( u2_u4_u2_n113 ) , .C1( u2_u4_u2_n132 ) , .A( u2_u4_u2_n149 ) , .B2( u2_u4_u2_n171 ) , .C2( u2_u4_u2_n172 ) , .ZN( u2_u4_u2_n96 ) );
  OAI221_X1 u2_u4_u2_U39 (.A( u2_u4_u2_n115 ) , .C2( u2_u4_u2_n123 ) , .B2( u2_u4_u2_n143 ) , .B1( u2_u4_u2_n153 ) , .ZN( u2_u4_u2_n163 ) , .C1( u2_u4_u2_n168 ) );
  INV_X1 u2_u4_u2_U4 (.A( u2_u4_u2_n134 ) , .ZN( u2_u4_u2_n185 ) );
  OAI21_X1 u2_u4_u2_U40 (.A( u2_u4_u2_n114 ) , .ZN( u2_u4_u2_n115 ) , .B1( u2_u4_u2_n176 ) , .B2( u2_u4_u2_n178 ) );
  OAI221_X1 u2_u4_u2_U41 (.A( u2_u4_u2_n135 ) , .B2( u2_u4_u2_n136 ) , .B1( u2_u4_u2_n137 ) , .ZN( u2_u4_u2_n162 ) , .C2( u2_u4_u2_n167 ) , .C1( u2_u4_u2_n185 ) );
  AND3_X1 u2_u4_u2_U42 (.A3( u2_u4_u2_n131 ) , .A2( u2_u4_u2_n132 ) , .A1( u2_u4_u2_n133 ) , .ZN( u2_u4_u2_n136 ) );
  AOI22_X1 u2_u4_u2_U43 (.ZN( u2_u4_u2_n135 ) , .B1( u2_u4_u2_n140 ) , .A1( u2_u4_u2_n156 ) , .B2( u2_u4_u2_n180 ) , .A2( u2_u4_u2_n188 ) );
  AOI21_X1 u2_u4_u2_U44 (.ZN( u2_u4_u2_n149 ) , .B1( u2_u4_u2_n173 ) , .B2( u2_u4_u2_n188 ) , .A( u2_u4_u2_n95 ) );
  AND3_X1 u2_u4_u2_U45 (.A2( u2_u4_u2_n100 ) , .A1( u2_u4_u2_n104 ) , .A3( u2_u4_u2_n156 ) , .ZN( u2_u4_u2_n95 ) );
  OAI21_X1 u2_u4_u2_U46 (.A( u2_u4_u2_n101 ) , .B2( u2_u4_u2_n121 ) , .B1( u2_u4_u2_n153 ) , .ZN( u2_u4_u2_n164 ) );
  NAND2_X1 u2_u4_u2_U47 (.A2( u2_u4_u2_n100 ) , .A1( u2_u4_u2_n107 ) , .ZN( u2_u4_u2_n155 ) );
  NAND2_X1 u2_u4_u2_U48 (.A2( u2_u4_u2_n105 ) , .A1( u2_u4_u2_n108 ) , .ZN( u2_u4_u2_n143 ) );
  NAND2_X1 u2_u4_u2_U49 (.A1( u2_u4_u2_n104 ) , .A2( u2_u4_u2_n106 ) , .ZN( u2_u4_u2_n152 ) );
  INV_X1 u2_u4_u2_U5 (.A( u2_u4_u2_n150 ) , .ZN( u2_u4_u2_n184 ) );
  NAND2_X1 u2_u4_u2_U50 (.A1( u2_u4_u2_n100 ) , .A2( u2_u4_u2_n105 ) , .ZN( u2_u4_u2_n132 ) );
  INV_X1 u2_u4_u2_U51 (.A( u2_u4_u2_n140 ) , .ZN( u2_u4_u2_n168 ) );
  INV_X1 u2_u4_u2_U52 (.A( u2_u4_u2_n138 ) , .ZN( u2_u4_u2_n167 ) );
  OAI21_X1 u2_u4_u2_U53 (.A( u2_u4_u2_n141 ) , .B2( u2_u4_u2_n142 ) , .ZN( u2_u4_u2_n146 ) , .B1( u2_u4_u2_n153 ) );
  OAI21_X1 u2_u4_u2_U54 (.A( u2_u4_u2_n140 ) , .ZN( u2_u4_u2_n141 ) , .B1( u2_u4_u2_n176 ) , .B2( u2_u4_u2_n177 ) );
  NOR3_X1 u2_u4_u2_U55 (.ZN( u2_u4_u2_n142 ) , .A3( u2_u4_u2_n175 ) , .A2( u2_u4_u2_n178 ) , .A1( u2_u4_u2_n181 ) );
  INV_X1 u2_u4_u2_U56 (.ZN( u2_u4_u2_n187 ) , .A( u2_u4_u2_n99 ) );
  OAI21_X1 u2_u4_u2_U57 (.B1( u2_u4_u2_n137 ) , .B2( u2_u4_u2_n143 ) , .A( u2_u4_u2_n98 ) , .ZN( u2_u4_u2_n99 ) );
  NAND2_X1 u2_u4_u2_U58 (.A1( u2_u4_u2_n102 ) , .A2( u2_u4_u2_n106 ) , .ZN( u2_u4_u2_n113 ) );
  NAND2_X1 u2_u4_u2_U59 (.A1( u2_u4_u2_n106 ) , .A2( u2_u4_u2_n107 ) , .ZN( u2_u4_u2_n131 ) );
  NOR4_X1 u2_u4_u2_U6 (.A4( u2_u4_u2_n124 ) , .A3( u2_u4_u2_n125 ) , .A2( u2_u4_u2_n126 ) , .A1( u2_u4_u2_n127 ) , .ZN( u2_u4_u2_n128 ) );
  NAND2_X1 u2_u4_u2_U60 (.A1( u2_u4_u2_n103 ) , .A2( u2_u4_u2_n107 ) , .ZN( u2_u4_u2_n139 ) );
  NAND2_X1 u2_u4_u2_U61 (.A1( u2_u4_u2_n103 ) , .A2( u2_u4_u2_n105 ) , .ZN( u2_u4_u2_n133 ) );
  NAND2_X1 u2_u4_u2_U62 (.A1( u2_u4_u2_n102 ) , .A2( u2_u4_u2_n103 ) , .ZN( u2_u4_u2_n154 ) );
  NAND2_X1 u2_u4_u2_U63 (.A2( u2_u4_u2_n103 ) , .A1( u2_u4_u2_n104 ) , .ZN( u2_u4_u2_n119 ) );
  NAND2_X1 u2_u4_u2_U64 (.A2( u2_u4_u2_n107 ) , .A1( u2_u4_u2_n108 ) , .ZN( u2_u4_u2_n123 ) );
  NAND2_X1 u2_u4_u2_U65 (.A1( u2_u4_u2_n104 ) , .A2( u2_u4_u2_n108 ) , .ZN( u2_u4_u2_n122 ) );
  INV_X1 u2_u4_u2_U66 (.A( u2_u4_u2_n114 ) , .ZN( u2_u4_u2_n172 ) );
  NAND2_X1 u2_u4_u2_U67 (.A2( u2_u4_u2_n100 ) , .A1( u2_u4_u2_n102 ) , .ZN( u2_u4_u2_n116 ) );
  NAND2_X1 u2_u4_u2_U68 (.A1( u2_u4_u2_n102 ) , .A2( u2_u4_u2_n108 ) , .ZN( u2_u4_u2_n120 ) );
  NAND2_X1 u2_u4_u2_U69 (.A2( u2_u4_u2_n105 ) , .A1( u2_u4_u2_n106 ) , .ZN( u2_u4_u2_n117 ) );
  AOI21_X1 u2_u4_u2_U7 (.B2( u2_u4_u2_n119 ) , .ZN( u2_u4_u2_n127 ) , .A( u2_u4_u2_n137 ) , .B1( u2_u4_u2_n155 ) );
  NOR2_X1 u2_u4_u2_U70 (.A2( u2_u4_X_16 ) , .ZN( u2_u4_u2_n140 ) , .A1( u2_u4_u2_n166 ) );
  NOR2_X1 u2_u4_u2_U71 (.A2( u2_u4_X_13 ) , .A1( u2_u4_X_14 ) , .ZN( u2_u4_u2_n100 ) );
  NOR2_X1 u2_u4_u2_U72 (.A2( u2_u4_X_16 ) , .A1( u2_u4_X_17 ) , .ZN( u2_u4_u2_n138 ) );
  NOR2_X1 u2_u4_u2_U73 (.A2( u2_u4_X_15 ) , .A1( u2_u4_X_18 ) , .ZN( u2_u4_u2_n104 ) );
  NOR2_X1 u2_u4_u2_U74 (.A2( u2_u4_X_14 ) , .ZN( u2_u4_u2_n103 ) , .A1( u2_u4_u2_n174 ) );
  NOR2_X1 u2_u4_u2_U75 (.A2( u2_u4_X_15 ) , .ZN( u2_u4_u2_n102 ) , .A1( u2_u4_u2_n165 ) );
  NOR2_X1 u2_u4_u2_U76 (.A2( u2_u4_X_17 ) , .ZN( u2_u4_u2_n114 ) , .A1( u2_u4_u2_n169 ) );
  AND2_X1 u2_u4_u2_U77 (.A1( u2_u4_X_15 ) , .ZN( u2_u4_u2_n105 ) , .A2( u2_u4_u2_n165 ) );
  AND2_X1 u2_u4_u2_U78 (.A2( u2_u4_X_15 ) , .A1( u2_u4_X_18 ) , .ZN( u2_u4_u2_n107 ) );
  AND2_X1 u2_u4_u2_U79 (.A1( u2_u4_X_14 ) , .ZN( u2_u4_u2_n106 ) , .A2( u2_u4_u2_n174 ) );
  AOI21_X1 u2_u4_u2_U8 (.ZN( u2_u4_u2_n124 ) , .B1( u2_u4_u2_n131 ) , .B2( u2_u4_u2_n143 ) , .A( u2_u4_u2_n172 ) );
  AND2_X1 u2_u4_u2_U80 (.A1( u2_u4_X_13 ) , .A2( u2_u4_X_14 ) , .ZN( u2_u4_u2_n108 ) );
  INV_X1 u2_u4_u2_U81 (.A( u2_u4_X_16 ) , .ZN( u2_u4_u2_n169 ) );
  INV_X1 u2_u4_u2_U82 (.A( u2_u4_X_17 ) , .ZN( u2_u4_u2_n166 ) );
  INV_X1 u2_u4_u2_U83 (.A( u2_u4_X_13 ) , .ZN( u2_u4_u2_n174 ) );
  INV_X1 u2_u4_u2_U84 (.A( u2_u4_X_18 ) , .ZN( u2_u4_u2_n165 ) );
  NAND4_X1 u2_u4_u2_U85 (.ZN( u2_out4_30 ) , .A4( u2_u4_u2_n147 ) , .A3( u2_u4_u2_n148 ) , .A2( u2_u4_u2_n149 ) , .A1( u2_u4_u2_n187 ) );
  NOR3_X1 u2_u4_u2_U86 (.A3( u2_u4_u2_n144 ) , .A2( u2_u4_u2_n145 ) , .A1( u2_u4_u2_n146 ) , .ZN( u2_u4_u2_n147 ) );
  AOI21_X1 u2_u4_u2_U87 (.B2( u2_u4_u2_n138 ) , .ZN( u2_u4_u2_n148 ) , .A( u2_u4_u2_n162 ) , .B1( u2_u4_u2_n182 ) );
  NAND4_X1 u2_u4_u2_U88 (.ZN( u2_out4_24 ) , .A4( u2_u4_u2_n111 ) , .A3( u2_u4_u2_n112 ) , .A1( u2_u4_u2_n130 ) , .A2( u2_u4_u2_n187 ) );
  AOI221_X1 u2_u4_u2_U89 (.A( u2_u4_u2_n109 ) , .B1( u2_u4_u2_n110 ) , .ZN( u2_u4_u2_n111 ) , .C1( u2_u4_u2_n134 ) , .C2( u2_u4_u2_n170 ) , .B2( u2_u4_u2_n173 ) );
  AOI21_X1 u2_u4_u2_U9 (.B2( u2_u4_u2_n123 ) , .ZN( u2_u4_u2_n125 ) , .A( u2_u4_u2_n171 ) , .B1( u2_u4_u2_n184 ) );
  AOI21_X1 u2_u4_u2_U90 (.ZN( u2_u4_u2_n112 ) , .B2( u2_u4_u2_n156 ) , .A( u2_u4_u2_n164 ) , .B1( u2_u4_u2_n181 ) );
  NAND4_X1 u2_u4_u2_U91 (.ZN( u2_out4_16 ) , .A4( u2_u4_u2_n128 ) , .A3( u2_u4_u2_n129 ) , .A1( u2_u4_u2_n130 ) , .A2( u2_u4_u2_n186 ) );
  AOI22_X1 u2_u4_u2_U92 (.A2( u2_u4_u2_n118 ) , .ZN( u2_u4_u2_n129 ) , .A1( u2_u4_u2_n140 ) , .B1( u2_u4_u2_n157 ) , .B2( u2_u4_u2_n170 ) );
  INV_X1 u2_u4_u2_U93 (.A( u2_u4_u2_n163 ) , .ZN( u2_u4_u2_n186 ) );
  OR4_X1 u2_u4_u2_U94 (.ZN( u2_out4_6 ) , .A4( u2_u4_u2_n161 ) , .A3( u2_u4_u2_n162 ) , .A2( u2_u4_u2_n163 ) , .A1( u2_u4_u2_n164 ) );
  OR3_X1 u2_u4_u2_U95 (.A2( u2_u4_u2_n159 ) , .A1( u2_u4_u2_n160 ) , .ZN( u2_u4_u2_n161 ) , .A3( u2_u4_u2_n183 ) );
  AOI21_X1 u2_u4_u2_U96 (.B2( u2_u4_u2_n154 ) , .B1( u2_u4_u2_n155 ) , .ZN( u2_u4_u2_n159 ) , .A( u2_u4_u2_n167 ) );
  NAND3_X1 u2_u4_u2_U97 (.A2( u2_u4_u2_n117 ) , .A1( u2_u4_u2_n122 ) , .A3( u2_u4_u2_n123 ) , .ZN( u2_u4_u2_n134 ) );
  NAND3_X1 u2_u4_u2_U98 (.ZN( u2_u4_u2_n110 ) , .A2( u2_u4_u2_n131 ) , .A3( u2_u4_u2_n139 ) , .A1( u2_u4_u2_n154 ) );
  NAND3_X1 u2_u4_u2_U99 (.A2( u2_u4_u2_n100 ) , .ZN( u2_u4_u2_n101 ) , .A1( u2_u4_u2_n104 ) , .A3( u2_u4_u2_n114 ) );
  OAI22_X1 u2_u4_u3_U10 (.B1( u2_u4_u3_n113 ) , .A2( u2_u4_u3_n135 ) , .A1( u2_u4_u3_n150 ) , .B2( u2_u4_u3_n164 ) , .ZN( u2_u4_u3_n98 ) );
  OAI211_X1 u2_u4_u3_U11 (.B( u2_u4_u3_n106 ) , .ZN( u2_u4_u3_n119 ) , .C2( u2_u4_u3_n128 ) , .C1( u2_u4_u3_n167 ) , .A( u2_u4_u3_n181 ) );
  AOI221_X1 u2_u4_u3_U12 (.C1( u2_u4_u3_n105 ) , .ZN( u2_u4_u3_n106 ) , .A( u2_u4_u3_n131 ) , .B2( u2_u4_u3_n132 ) , .C2( u2_u4_u3_n133 ) , .B1( u2_u4_u3_n169 ) );
  INV_X1 u2_u4_u3_U13 (.ZN( u2_u4_u3_n181 ) , .A( u2_u4_u3_n98 ) );
  NAND2_X1 u2_u4_u3_U14 (.ZN( u2_u4_u3_n105 ) , .A2( u2_u4_u3_n130 ) , .A1( u2_u4_u3_n155 ) );
  AOI22_X1 u2_u4_u3_U15 (.B1( u2_u4_u3_n115 ) , .A2( u2_u4_u3_n116 ) , .ZN( u2_u4_u3_n123 ) , .B2( u2_u4_u3_n133 ) , .A1( u2_u4_u3_n169 ) );
  NAND2_X1 u2_u4_u3_U16 (.ZN( u2_u4_u3_n116 ) , .A2( u2_u4_u3_n151 ) , .A1( u2_u4_u3_n182 ) );
  NOR2_X1 u2_u4_u3_U17 (.ZN( u2_u4_u3_n126 ) , .A2( u2_u4_u3_n150 ) , .A1( u2_u4_u3_n164 ) );
  AOI21_X1 u2_u4_u3_U18 (.ZN( u2_u4_u3_n112 ) , .B2( u2_u4_u3_n146 ) , .B1( u2_u4_u3_n155 ) , .A( u2_u4_u3_n167 ) );
  NAND2_X1 u2_u4_u3_U19 (.A1( u2_u4_u3_n135 ) , .ZN( u2_u4_u3_n142 ) , .A2( u2_u4_u3_n164 ) );
  NAND2_X1 u2_u4_u3_U20 (.ZN( u2_u4_u3_n132 ) , .A2( u2_u4_u3_n152 ) , .A1( u2_u4_u3_n156 ) );
  AND2_X1 u2_u4_u3_U21 (.A2( u2_u4_u3_n113 ) , .A1( u2_u4_u3_n114 ) , .ZN( u2_u4_u3_n151 ) );
  INV_X1 u2_u4_u3_U22 (.A( u2_u4_u3_n133 ) , .ZN( u2_u4_u3_n165 ) );
  INV_X1 u2_u4_u3_U23 (.A( u2_u4_u3_n135 ) , .ZN( u2_u4_u3_n170 ) );
  NAND2_X1 u2_u4_u3_U24 (.A1( u2_u4_u3_n107 ) , .A2( u2_u4_u3_n108 ) , .ZN( u2_u4_u3_n140 ) );
  NAND2_X1 u2_u4_u3_U25 (.ZN( u2_u4_u3_n117 ) , .A1( u2_u4_u3_n124 ) , .A2( u2_u4_u3_n148 ) );
  NAND2_X1 u2_u4_u3_U26 (.ZN( u2_u4_u3_n143 ) , .A1( u2_u4_u3_n165 ) , .A2( u2_u4_u3_n167 ) );
  INV_X1 u2_u4_u3_U27 (.A( u2_u4_u3_n130 ) , .ZN( u2_u4_u3_n177 ) );
  INV_X1 u2_u4_u3_U28 (.A( u2_u4_u3_n128 ) , .ZN( u2_u4_u3_n176 ) );
  INV_X1 u2_u4_u3_U29 (.A( u2_u4_u3_n155 ) , .ZN( u2_u4_u3_n174 ) );
  INV_X1 u2_u4_u3_U3 (.A( u2_u4_u3_n129 ) , .ZN( u2_u4_u3_n183 ) );
  INV_X1 u2_u4_u3_U30 (.A( u2_u4_u3_n139 ) , .ZN( u2_u4_u3_n185 ) );
  NOR2_X1 u2_u4_u3_U31 (.ZN( u2_u4_u3_n135 ) , .A2( u2_u4_u3_n141 ) , .A1( u2_u4_u3_n169 ) );
  OAI222_X1 u2_u4_u3_U32 (.C2( u2_u4_u3_n107 ) , .A2( u2_u4_u3_n108 ) , .B1( u2_u4_u3_n135 ) , .ZN( u2_u4_u3_n138 ) , .B2( u2_u4_u3_n146 ) , .C1( u2_u4_u3_n154 ) , .A1( u2_u4_u3_n164 ) );
  NOR4_X1 u2_u4_u3_U33 (.A4( u2_u4_u3_n157 ) , .A3( u2_u4_u3_n158 ) , .A2( u2_u4_u3_n159 ) , .A1( u2_u4_u3_n160 ) , .ZN( u2_u4_u3_n161 ) );
  AOI21_X1 u2_u4_u3_U34 (.B2( u2_u4_u3_n152 ) , .B1( u2_u4_u3_n153 ) , .ZN( u2_u4_u3_n158 ) , .A( u2_u4_u3_n164 ) );
  AOI21_X1 u2_u4_u3_U35 (.A( u2_u4_u3_n149 ) , .B2( u2_u4_u3_n150 ) , .B1( u2_u4_u3_n151 ) , .ZN( u2_u4_u3_n159 ) );
  AOI21_X1 u2_u4_u3_U36 (.A( u2_u4_u3_n154 ) , .B2( u2_u4_u3_n155 ) , .B1( u2_u4_u3_n156 ) , .ZN( u2_u4_u3_n157 ) );
  AOI211_X1 u2_u4_u3_U37 (.ZN( u2_u4_u3_n109 ) , .A( u2_u4_u3_n119 ) , .C2( u2_u4_u3_n129 ) , .B( u2_u4_u3_n138 ) , .C1( u2_u4_u3_n141 ) );
  AOI211_X1 u2_u4_u3_U38 (.B( u2_u4_u3_n119 ) , .A( u2_u4_u3_n120 ) , .C2( u2_u4_u3_n121 ) , .ZN( u2_u4_u3_n122 ) , .C1( u2_u4_u3_n179 ) );
  INV_X1 u2_u4_u3_U39 (.A( u2_u4_u3_n156 ) , .ZN( u2_u4_u3_n179 ) );
  INV_X1 u2_u4_u3_U4 (.A( u2_u4_u3_n140 ) , .ZN( u2_u4_u3_n182 ) );
  OAI22_X1 u2_u4_u3_U40 (.B1( u2_u4_u3_n118 ) , .ZN( u2_u4_u3_n120 ) , .A1( u2_u4_u3_n135 ) , .B2( u2_u4_u3_n154 ) , .A2( u2_u4_u3_n178 ) );
  AND3_X1 u2_u4_u3_U41 (.ZN( u2_u4_u3_n118 ) , .A2( u2_u4_u3_n124 ) , .A1( u2_u4_u3_n144 ) , .A3( u2_u4_u3_n152 ) );
  INV_X1 u2_u4_u3_U42 (.A( u2_u4_u3_n121 ) , .ZN( u2_u4_u3_n164 ) );
  NAND2_X1 u2_u4_u3_U43 (.ZN( u2_u4_u3_n133 ) , .A1( u2_u4_u3_n154 ) , .A2( u2_u4_u3_n164 ) );
  OAI211_X1 u2_u4_u3_U44 (.B( u2_u4_u3_n127 ) , .ZN( u2_u4_u3_n139 ) , .C1( u2_u4_u3_n150 ) , .C2( u2_u4_u3_n154 ) , .A( u2_u4_u3_n184 ) );
  INV_X1 u2_u4_u3_U45 (.A( u2_u4_u3_n125 ) , .ZN( u2_u4_u3_n184 ) );
  AOI221_X1 u2_u4_u3_U46 (.A( u2_u4_u3_n126 ) , .ZN( u2_u4_u3_n127 ) , .C2( u2_u4_u3_n132 ) , .C1( u2_u4_u3_n169 ) , .B2( u2_u4_u3_n170 ) , .B1( u2_u4_u3_n174 ) );
  OAI22_X1 u2_u4_u3_U47 (.A1( u2_u4_u3_n124 ) , .ZN( u2_u4_u3_n125 ) , .B2( u2_u4_u3_n145 ) , .A2( u2_u4_u3_n165 ) , .B1( u2_u4_u3_n167 ) );
  NOR2_X1 u2_u4_u3_U48 (.A1( u2_u4_u3_n113 ) , .ZN( u2_u4_u3_n131 ) , .A2( u2_u4_u3_n154 ) );
  NAND2_X1 u2_u4_u3_U49 (.A1( u2_u4_u3_n103 ) , .ZN( u2_u4_u3_n150 ) , .A2( u2_u4_u3_n99 ) );
  INV_X1 u2_u4_u3_U5 (.A( u2_u4_u3_n117 ) , .ZN( u2_u4_u3_n178 ) );
  NAND2_X1 u2_u4_u3_U50 (.A2( u2_u4_u3_n102 ) , .ZN( u2_u4_u3_n155 ) , .A1( u2_u4_u3_n97 ) );
  INV_X1 u2_u4_u3_U51 (.A( u2_u4_u3_n141 ) , .ZN( u2_u4_u3_n167 ) );
  AOI21_X1 u2_u4_u3_U52 (.B2( u2_u4_u3_n114 ) , .B1( u2_u4_u3_n146 ) , .A( u2_u4_u3_n154 ) , .ZN( u2_u4_u3_n94 ) );
  AOI21_X1 u2_u4_u3_U53 (.ZN( u2_u4_u3_n110 ) , .B2( u2_u4_u3_n142 ) , .B1( u2_u4_u3_n186 ) , .A( u2_u4_u3_n95 ) );
  INV_X1 u2_u4_u3_U54 (.A( u2_u4_u3_n145 ) , .ZN( u2_u4_u3_n186 ) );
  AOI21_X1 u2_u4_u3_U55 (.B1( u2_u4_u3_n124 ) , .A( u2_u4_u3_n149 ) , .B2( u2_u4_u3_n155 ) , .ZN( u2_u4_u3_n95 ) );
  INV_X1 u2_u4_u3_U56 (.A( u2_u4_u3_n149 ) , .ZN( u2_u4_u3_n169 ) );
  NAND2_X1 u2_u4_u3_U57 (.ZN( u2_u4_u3_n124 ) , .A1( u2_u4_u3_n96 ) , .A2( u2_u4_u3_n97 ) );
  NAND2_X1 u2_u4_u3_U58 (.A2( u2_u4_u3_n100 ) , .ZN( u2_u4_u3_n146 ) , .A1( u2_u4_u3_n96 ) );
  NAND2_X1 u2_u4_u3_U59 (.A1( u2_u4_u3_n101 ) , .ZN( u2_u4_u3_n145 ) , .A2( u2_u4_u3_n99 ) );
  AOI221_X1 u2_u4_u3_U6 (.A( u2_u4_u3_n131 ) , .C2( u2_u4_u3_n132 ) , .C1( u2_u4_u3_n133 ) , .ZN( u2_u4_u3_n134 ) , .B1( u2_u4_u3_n143 ) , .B2( u2_u4_u3_n177 ) );
  NAND2_X1 u2_u4_u3_U60 (.A1( u2_u4_u3_n100 ) , .ZN( u2_u4_u3_n156 ) , .A2( u2_u4_u3_n99 ) );
  NAND2_X1 u2_u4_u3_U61 (.A2( u2_u4_u3_n101 ) , .A1( u2_u4_u3_n104 ) , .ZN( u2_u4_u3_n148 ) );
  NAND2_X1 u2_u4_u3_U62 (.A1( u2_u4_u3_n100 ) , .A2( u2_u4_u3_n102 ) , .ZN( u2_u4_u3_n128 ) );
  NAND2_X1 u2_u4_u3_U63 (.A2( u2_u4_u3_n101 ) , .A1( u2_u4_u3_n102 ) , .ZN( u2_u4_u3_n152 ) );
  NAND2_X1 u2_u4_u3_U64 (.A2( u2_u4_u3_n101 ) , .ZN( u2_u4_u3_n114 ) , .A1( u2_u4_u3_n96 ) );
  NAND2_X1 u2_u4_u3_U65 (.ZN( u2_u4_u3_n107 ) , .A1( u2_u4_u3_n97 ) , .A2( u2_u4_u3_n99 ) );
  NAND2_X1 u2_u4_u3_U66 (.A2( u2_u4_u3_n100 ) , .A1( u2_u4_u3_n104 ) , .ZN( u2_u4_u3_n113 ) );
  NAND2_X1 u2_u4_u3_U67 (.A1( u2_u4_u3_n104 ) , .ZN( u2_u4_u3_n153 ) , .A2( u2_u4_u3_n97 ) );
  NAND2_X1 u2_u4_u3_U68 (.A2( u2_u4_u3_n103 ) , .A1( u2_u4_u3_n104 ) , .ZN( u2_u4_u3_n130 ) );
  NAND2_X1 u2_u4_u3_U69 (.A2( u2_u4_u3_n103 ) , .ZN( u2_u4_u3_n144 ) , .A1( u2_u4_u3_n96 ) );
  OAI22_X1 u2_u4_u3_U7 (.B2( u2_u4_u3_n147 ) , .A2( u2_u4_u3_n148 ) , .ZN( u2_u4_u3_n160 ) , .B1( u2_u4_u3_n165 ) , .A1( u2_u4_u3_n168 ) );
  NAND2_X1 u2_u4_u3_U70 (.A1( u2_u4_u3_n102 ) , .A2( u2_u4_u3_n103 ) , .ZN( u2_u4_u3_n108 ) );
  NOR2_X1 u2_u4_u3_U71 (.A2( u2_u4_X_19 ) , .A1( u2_u4_X_20 ) , .ZN( u2_u4_u3_n99 ) );
  NOR2_X1 u2_u4_u3_U72 (.A2( u2_u4_X_21 ) , .A1( u2_u4_X_24 ) , .ZN( u2_u4_u3_n103 ) );
  NOR2_X1 u2_u4_u3_U73 (.A2( u2_u4_X_24 ) , .A1( u2_u4_u3_n171 ) , .ZN( u2_u4_u3_n97 ) );
  NOR2_X1 u2_u4_u3_U74 (.A2( u2_u4_X_23 ) , .ZN( u2_u4_u3_n141 ) , .A1( u2_u4_u3_n166 ) );
  NOR2_X1 u2_u4_u3_U75 (.A2( u2_u4_X_19 ) , .A1( u2_u4_u3_n172 ) , .ZN( u2_u4_u3_n96 ) );
  NAND2_X1 u2_u4_u3_U76 (.A1( u2_u4_X_22 ) , .A2( u2_u4_X_23 ) , .ZN( u2_u4_u3_n154 ) );
  NAND2_X1 u2_u4_u3_U77 (.A1( u2_u4_X_23 ) , .ZN( u2_u4_u3_n149 ) , .A2( u2_u4_u3_n166 ) );
  NOR2_X1 u2_u4_u3_U78 (.A2( u2_u4_X_22 ) , .A1( u2_u4_X_23 ) , .ZN( u2_u4_u3_n121 ) );
  AND2_X1 u2_u4_u3_U79 (.A1( u2_u4_X_24 ) , .ZN( u2_u4_u3_n101 ) , .A2( u2_u4_u3_n171 ) );
  AND3_X1 u2_u4_u3_U8 (.A3( u2_u4_u3_n144 ) , .A2( u2_u4_u3_n145 ) , .A1( u2_u4_u3_n146 ) , .ZN( u2_u4_u3_n147 ) );
  AND2_X1 u2_u4_u3_U80 (.A1( u2_u4_X_19 ) , .ZN( u2_u4_u3_n102 ) , .A2( u2_u4_u3_n172 ) );
  AND2_X1 u2_u4_u3_U81 (.A1( u2_u4_X_21 ) , .A2( u2_u4_X_24 ) , .ZN( u2_u4_u3_n100 ) );
  AND2_X1 u2_u4_u3_U82 (.A2( u2_u4_X_19 ) , .A1( u2_u4_X_20 ) , .ZN( u2_u4_u3_n104 ) );
  INV_X1 u2_u4_u3_U83 (.A( u2_u4_X_22 ) , .ZN( u2_u4_u3_n166 ) );
  INV_X1 u2_u4_u3_U84 (.A( u2_u4_X_21 ) , .ZN( u2_u4_u3_n171 ) );
  INV_X1 u2_u4_u3_U85 (.A( u2_u4_X_20 ) , .ZN( u2_u4_u3_n172 ) );
  OR4_X1 u2_u4_u3_U86 (.ZN( u2_out4_10 ) , .A4( u2_u4_u3_n136 ) , .A3( u2_u4_u3_n137 ) , .A1( u2_u4_u3_n138 ) , .A2( u2_u4_u3_n139 ) );
  OAI222_X1 u2_u4_u3_U87 (.C1( u2_u4_u3_n128 ) , .ZN( u2_u4_u3_n137 ) , .B1( u2_u4_u3_n148 ) , .A2( u2_u4_u3_n150 ) , .B2( u2_u4_u3_n154 ) , .C2( u2_u4_u3_n164 ) , .A1( u2_u4_u3_n167 ) );
  OAI221_X1 u2_u4_u3_U88 (.A( u2_u4_u3_n134 ) , .B2( u2_u4_u3_n135 ) , .ZN( u2_u4_u3_n136 ) , .C1( u2_u4_u3_n149 ) , .B1( u2_u4_u3_n151 ) , .C2( u2_u4_u3_n183 ) );
  NAND4_X1 u2_u4_u3_U89 (.ZN( u2_out4_26 ) , .A4( u2_u4_u3_n109 ) , .A3( u2_u4_u3_n110 ) , .A2( u2_u4_u3_n111 ) , .A1( u2_u4_u3_n173 ) );
  INV_X1 u2_u4_u3_U9 (.A( u2_u4_u3_n143 ) , .ZN( u2_u4_u3_n168 ) );
  INV_X1 u2_u4_u3_U90 (.ZN( u2_u4_u3_n173 ) , .A( u2_u4_u3_n94 ) );
  OAI21_X1 u2_u4_u3_U91 (.ZN( u2_u4_u3_n111 ) , .B2( u2_u4_u3_n117 ) , .A( u2_u4_u3_n133 ) , .B1( u2_u4_u3_n176 ) );
  NAND4_X1 u2_u4_u3_U92 (.ZN( u2_out4_20 ) , .A4( u2_u4_u3_n122 ) , .A3( u2_u4_u3_n123 ) , .A1( u2_u4_u3_n175 ) , .A2( u2_u4_u3_n180 ) );
  INV_X1 u2_u4_u3_U93 (.A( u2_u4_u3_n126 ) , .ZN( u2_u4_u3_n180 ) );
  INV_X1 u2_u4_u3_U94 (.A( u2_u4_u3_n112 ) , .ZN( u2_u4_u3_n175 ) );
  NAND4_X1 u2_u4_u3_U95 (.ZN( u2_out4_1 ) , .A4( u2_u4_u3_n161 ) , .A3( u2_u4_u3_n162 ) , .A2( u2_u4_u3_n163 ) , .A1( u2_u4_u3_n185 ) );
  NAND2_X1 u2_u4_u3_U96 (.ZN( u2_u4_u3_n163 ) , .A2( u2_u4_u3_n170 ) , .A1( u2_u4_u3_n176 ) );
  AOI22_X1 u2_u4_u3_U97 (.B2( u2_u4_u3_n140 ) , .B1( u2_u4_u3_n141 ) , .A2( u2_u4_u3_n142 ) , .ZN( u2_u4_u3_n162 ) , .A1( u2_u4_u3_n177 ) );
  NAND3_X1 u2_u4_u3_U98 (.A1( u2_u4_u3_n114 ) , .ZN( u2_u4_u3_n115 ) , .A2( u2_u4_u3_n145 ) , .A3( u2_u4_u3_n153 ) );
  NAND3_X1 u2_u4_u3_U99 (.ZN( u2_u4_u3_n129 ) , .A2( u2_u4_u3_n144 ) , .A1( u2_u4_u3_n153 ) , .A3( u2_u4_u3_n182 ) );
  OAI22_X1 u2_u4_u4_U10 (.B2( u2_u4_u4_n135 ) , .ZN( u2_u4_u4_n137 ) , .B1( u2_u4_u4_n153 ) , .A1( u2_u4_u4_n155 ) , .A2( u2_u4_u4_n171 ) );
  AND3_X1 u2_u4_u4_U11 (.A2( u2_u4_u4_n134 ) , .ZN( u2_u4_u4_n135 ) , .A3( u2_u4_u4_n145 ) , .A1( u2_u4_u4_n157 ) );
  NAND2_X1 u2_u4_u4_U12 (.ZN( u2_u4_u4_n132 ) , .A2( u2_u4_u4_n170 ) , .A1( u2_u4_u4_n173 ) );
  AOI21_X1 u2_u4_u4_U13 (.B2( u2_u4_u4_n160 ) , .B1( u2_u4_u4_n161 ) , .ZN( u2_u4_u4_n162 ) , .A( u2_u4_u4_n170 ) );
  AOI21_X1 u2_u4_u4_U14 (.ZN( u2_u4_u4_n107 ) , .B2( u2_u4_u4_n143 ) , .A( u2_u4_u4_n174 ) , .B1( u2_u4_u4_n184 ) );
  AOI21_X1 u2_u4_u4_U15 (.B2( u2_u4_u4_n158 ) , .B1( u2_u4_u4_n159 ) , .ZN( u2_u4_u4_n163 ) , .A( u2_u4_u4_n174 ) );
  AOI21_X1 u2_u4_u4_U16 (.A( u2_u4_u4_n153 ) , .B2( u2_u4_u4_n154 ) , .B1( u2_u4_u4_n155 ) , .ZN( u2_u4_u4_n165 ) );
  AOI21_X1 u2_u4_u4_U17 (.A( u2_u4_u4_n156 ) , .B2( u2_u4_u4_n157 ) , .ZN( u2_u4_u4_n164 ) , .B1( u2_u4_u4_n184 ) );
  INV_X1 u2_u4_u4_U18 (.A( u2_u4_u4_n138 ) , .ZN( u2_u4_u4_n170 ) );
  AND2_X1 u2_u4_u4_U19 (.A2( u2_u4_u4_n120 ) , .ZN( u2_u4_u4_n155 ) , .A1( u2_u4_u4_n160 ) );
  INV_X1 u2_u4_u4_U20 (.A( u2_u4_u4_n156 ) , .ZN( u2_u4_u4_n175 ) );
  NAND2_X1 u2_u4_u4_U21 (.A2( u2_u4_u4_n118 ) , .ZN( u2_u4_u4_n131 ) , .A1( u2_u4_u4_n147 ) );
  NAND2_X1 u2_u4_u4_U22 (.A1( u2_u4_u4_n119 ) , .A2( u2_u4_u4_n120 ) , .ZN( u2_u4_u4_n130 ) );
  NAND2_X1 u2_u4_u4_U23 (.ZN( u2_u4_u4_n117 ) , .A2( u2_u4_u4_n118 ) , .A1( u2_u4_u4_n148 ) );
  NAND2_X1 u2_u4_u4_U24 (.ZN( u2_u4_u4_n129 ) , .A1( u2_u4_u4_n134 ) , .A2( u2_u4_u4_n148 ) );
  AND3_X1 u2_u4_u4_U25 (.A1( u2_u4_u4_n119 ) , .A2( u2_u4_u4_n143 ) , .A3( u2_u4_u4_n154 ) , .ZN( u2_u4_u4_n161 ) );
  AND2_X1 u2_u4_u4_U26 (.A1( u2_u4_u4_n145 ) , .A2( u2_u4_u4_n147 ) , .ZN( u2_u4_u4_n159 ) );
  OR3_X1 u2_u4_u4_U27 (.A3( u2_u4_u4_n114 ) , .A2( u2_u4_u4_n115 ) , .A1( u2_u4_u4_n116 ) , .ZN( u2_u4_u4_n136 ) );
  AOI21_X1 u2_u4_u4_U28 (.A( u2_u4_u4_n113 ) , .ZN( u2_u4_u4_n116 ) , .B2( u2_u4_u4_n173 ) , .B1( u2_u4_u4_n174 ) );
  AOI21_X1 u2_u4_u4_U29 (.ZN( u2_u4_u4_n115 ) , .B2( u2_u4_u4_n145 ) , .B1( u2_u4_u4_n146 ) , .A( u2_u4_u4_n156 ) );
  NOR2_X1 u2_u4_u4_U3 (.ZN( u2_u4_u4_n121 ) , .A1( u2_u4_u4_n181 ) , .A2( u2_u4_u4_n182 ) );
  OAI22_X1 u2_u4_u4_U30 (.ZN( u2_u4_u4_n114 ) , .A2( u2_u4_u4_n121 ) , .B1( u2_u4_u4_n160 ) , .B2( u2_u4_u4_n170 ) , .A1( u2_u4_u4_n171 ) );
  INV_X1 u2_u4_u4_U31 (.A( u2_u4_u4_n158 ) , .ZN( u2_u4_u4_n182 ) );
  INV_X1 u2_u4_u4_U32 (.ZN( u2_u4_u4_n181 ) , .A( u2_u4_u4_n96 ) );
  INV_X1 u2_u4_u4_U33 (.A( u2_u4_u4_n144 ) , .ZN( u2_u4_u4_n179 ) );
  INV_X1 u2_u4_u4_U34 (.A( u2_u4_u4_n157 ) , .ZN( u2_u4_u4_n178 ) );
  NAND2_X1 u2_u4_u4_U35 (.A2( u2_u4_u4_n154 ) , .A1( u2_u4_u4_n96 ) , .ZN( u2_u4_u4_n97 ) );
  INV_X1 u2_u4_u4_U36 (.ZN( u2_u4_u4_n186 ) , .A( u2_u4_u4_n95 ) );
  OAI221_X1 u2_u4_u4_U37 (.C1( u2_u4_u4_n134 ) , .B1( u2_u4_u4_n158 ) , .B2( u2_u4_u4_n171 ) , .C2( u2_u4_u4_n173 ) , .A( u2_u4_u4_n94 ) , .ZN( u2_u4_u4_n95 ) );
  AOI222_X1 u2_u4_u4_U38 (.B2( u2_u4_u4_n132 ) , .A1( u2_u4_u4_n138 ) , .C2( u2_u4_u4_n175 ) , .A2( u2_u4_u4_n179 ) , .C1( u2_u4_u4_n181 ) , .B1( u2_u4_u4_n185 ) , .ZN( u2_u4_u4_n94 ) );
  INV_X1 u2_u4_u4_U39 (.A( u2_u4_u4_n113 ) , .ZN( u2_u4_u4_n185 ) );
  INV_X1 u2_u4_u4_U4 (.A( u2_u4_u4_n117 ) , .ZN( u2_u4_u4_n184 ) );
  INV_X1 u2_u4_u4_U40 (.A( u2_u4_u4_n143 ) , .ZN( u2_u4_u4_n183 ) );
  NOR2_X1 u2_u4_u4_U41 (.ZN( u2_u4_u4_n138 ) , .A1( u2_u4_u4_n168 ) , .A2( u2_u4_u4_n169 ) );
  NOR2_X1 u2_u4_u4_U42 (.A1( u2_u4_u4_n150 ) , .A2( u2_u4_u4_n152 ) , .ZN( u2_u4_u4_n153 ) );
  NOR2_X1 u2_u4_u4_U43 (.A2( u2_u4_u4_n128 ) , .A1( u2_u4_u4_n138 ) , .ZN( u2_u4_u4_n156 ) );
  AOI22_X1 u2_u4_u4_U44 (.B2( u2_u4_u4_n122 ) , .A1( u2_u4_u4_n123 ) , .ZN( u2_u4_u4_n124 ) , .B1( u2_u4_u4_n128 ) , .A2( u2_u4_u4_n172 ) );
  INV_X1 u2_u4_u4_U45 (.A( u2_u4_u4_n153 ) , .ZN( u2_u4_u4_n172 ) );
  NAND2_X1 u2_u4_u4_U46 (.A2( u2_u4_u4_n120 ) , .ZN( u2_u4_u4_n123 ) , .A1( u2_u4_u4_n161 ) );
  AOI22_X1 u2_u4_u4_U47 (.B2( u2_u4_u4_n132 ) , .A2( u2_u4_u4_n133 ) , .ZN( u2_u4_u4_n140 ) , .A1( u2_u4_u4_n150 ) , .B1( u2_u4_u4_n179 ) );
  NAND2_X1 u2_u4_u4_U48 (.ZN( u2_u4_u4_n133 ) , .A2( u2_u4_u4_n146 ) , .A1( u2_u4_u4_n154 ) );
  NAND2_X1 u2_u4_u4_U49 (.A1( u2_u4_u4_n103 ) , .ZN( u2_u4_u4_n154 ) , .A2( u2_u4_u4_n98 ) );
  NOR4_X1 u2_u4_u4_U5 (.A4( u2_u4_u4_n106 ) , .A3( u2_u4_u4_n107 ) , .A2( u2_u4_u4_n108 ) , .A1( u2_u4_u4_n109 ) , .ZN( u2_u4_u4_n110 ) );
  NAND2_X1 u2_u4_u4_U50 (.A1( u2_u4_u4_n101 ) , .ZN( u2_u4_u4_n158 ) , .A2( u2_u4_u4_n99 ) );
  AOI21_X1 u2_u4_u4_U51 (.ZN( u2_u4_u4_n127 ) , .A( u2_u4_u4_n136 ) , .B2( u2_u4_u4_n150 ) , .B1( u2_u4_u4_n180 ) );
  INV_X1 u2_u4_u4_U52 (.A( u2_u4_u4_n160 ) , .ZN( u2_u4_u4_n180 ) );
  NAND2_X1 u2_u4_u4_U53 (.A2( u2_u4_u4_n104 ) , .A1( u2_u4_u4_n105 ) , .ZN( u2_u4_u4_n146 ) );
  NAND2_X1 u2_u4_u4_U54 (.A2( u2_u4_u4_n101 ) , .A1( u2_u4_u4_n102 ) , .ZN( u2_u4_u4_n160 ) );
  NAND2_X1 u2_u4_u4_U55 (.ZN( u2_u4_u4_n134 ) , .A1( u2_u4_u4_n98 ) , .A2( u2_u4_u4_n99 ) );
  NAND2_X1 u2_u4_u4_U56 (.A1( u2_u4_u4_n103 ) , .A2( u2_u4_u4_n104 ) , .ZN( u2_u4_u4_n143 ) );
  NAND2_X1 u2_u4_u4_U57 (.A2( u2_u4_u4_n105 ) , .ZN( u2_u4_u4_n145 ) , .A1( u2_u4_u4_n98 ) );
  NAND2_X1 u2_u4_u4_U58 (.A1( u2_u4_u4_n100 ) , .A2( u2_u4_u4_n105 ) , .ZN( u2_u4_u4_n120 ) );
  NAND2_X1 u2_u4_u4_U59 (.A1( u2_u4_u4_n102 ) , .A2( u2_u4_u4_n104 ) , .ZN( u2_u4_u4_n148 ) );
  AOI21_X1 u2_u4_u4_U6 (.ZN( u2_u4_u4_n106 ) , .B2( u2_u4_u4_n146 ) , .B1( u2_u4_u4_n158 ) , .A( u2_u4_u4_n170 ) );
  NAND2_X1 u2_u4_u4_U60 (.A2( u2_u4_u4_n100 ) , .A1( u2_u4_u4_n103 ) , .ZN( u2_u4_u4_n157 ) );
  INV_X1 u2_u4_u4_U61 (.A( u2_u4_u4_n150 ) , .ZN( u2_u4_u4_n173 ) );
  INV_X1 u2_u4_u4_U62 (.A( u2_u4_u4_n152 ) , .ZN( u2_u4_u4_n171 ) );
  NAND2_X1 u2_u4_u4_U63 (.A1( u2_u4_u4_n100 ) , .ZN( u2_u4_u4_n118 ) , .A2( u2_u4_u4_n99 ) );
  NAND2_X1 u2_u4_u4_U64 (.A2( u2_u4_u4_n100 ) , .A1( u2_u4_u4_n102 ) , .ZN( u2_u4_u4_n144 ) );
  NAND2_X1 u2_u4_u4_U65 (.A2( u2_u4_u4_n101 ) , .A1( u2_u4_u4_n105 ) , .ZN( u2_u4_u4_n96 ) );
  INV_X1 u2_u4_u4_U66 (.A( u2_u4_u4_n128 ) , .ZN( u2_u4_u4_n174 ) );
  NAND2_X1 u2_u4_u4_U67 (.A2( u2_u4_u4_n102 ) , .ZN( u2_u4_u4_n119 ) , .A1( u2_u4_u4_n98 ) );
  NAND2_X1 u2_u4_u4_U68 (.A2( u2_u4_u4_n101 ) , .A1( u2_u4_u4_n103 ) , .ZN( u2_u4_u4_n147 ) );
  NAND2_X1 u2_u4_u4_U69 (.A2( u2_u4_u4_n104 ) , .ZN( u2_u4_u4_n113 ) , .A1( u2_u4_u4_n99 ) );
  AOI21_X1 u2_u4_u4_U7 (.ZN( u2_u4_u4_n108 ) , .B2( u2_u4_u4_n134 ) , .B1( u2_u4_u4_n155 ) , .A( u2_u4_u4_n156 ) );
  NOR2_X1 u2_u4_u4_U70 (.A2( u2_u4_X_28 ) , .ZN( u2_u4_u4_n150 ) , .A1( u2_u4_u4_n168 ) );
  NOR2_X1 u2_u4_u4_U71 (.A2( u2_u4_X_29 ) , .ZN( u2_u4_u4_n152 ) , .A1( u2_u4_u4_n169 ) );
  NOR2_X1 u2_u4_u4_U72 (.A2( u2_u4_X_30 ) , .ZN( u2_u4_u4_n105 ) , .A1( u2_u4_u4_n176 ) );
  NOR2_X1 u2_u4_u4_U73 (.A2( u2_u4_X_26 ) , .ZN( u2_u4_u4_n100 ) , .A1( u2_u4_u4_n177 ) );
  NOR2_X1 u2_u4_u4_U74 (.A2( u2_u4_X_28 ) , .A1( u2_u4_X_29 ) , .ZN( u2_u4_u4_n128 ) );
  NOR2_X1 u2_u4_u4_U75 (.A2( u2_u4_X_27 ) , .A1( u2_u4_X_30 ) , .ZN( u2_u4_u4_n102 ) );
  NOR2_X1 u2_u4_u4_U76 (.A2( u2_u4_X_25 ) , .A1( u2_u4_X_26 ) , .ZN( u2_u4_u4_n98 ) );
  AND2_X1 u2_u4_u4_U77 (.A2( u2_u4_X_25 ) , .A1( u2_u4_X_26 ) , .ZN( u2_u4_u4_n104 ) );
  AND2_X1 u2_u4_u4_U78 (.A1( u2_u4_X_30 ) , .A2( u2_u4_u4_n176 ) , .ZN( u2_u4_u4_n99 ) );
  AND2_X1 u2_u4_u4_U79 (.A1( u2_u4_X_26 ) , .ZN( u2_u4_u4_n101 ) , .A2( u2_u4_u4_n177 ) );
  AOI21_X1 u2_u4_u4_U8 (.ZN( u2_u4_u4_n109 ) , .A( u2_u4_u4_n153 ) , .B1( u2_u4_u4_n159 ) , .B2( u2_u4_u4_n184 ) );
  AND2_X1 u2_u4_u4_U80 (.A1( u2_u4_X_27 ) , .A2( u2_u4_X_30 ) , .ZN( u2_u4_u4_n103 ) );
  INV_X1 u2_u4_u4_U81 (.A( u2_u4_X_28 ) , .ZN( u2_u4_u4_n169 ) );
  INV_X1 u2_u4_u4_U82 (.A( u2_u4_X_29 ) , .ZN( u2_u4_u4_n168 ) );
  INV_X1 u2_u4_u4_U83 (.A( u2_u4_X_25 ) , .ZN( u2_u4_u4_n177 ) );
  INV_X1 u2_u4_u4_U84 (.A( u2_u4_X_27 ) , .ZN( u2_u4_u4_n176 ) );
  NAND4_X1 u2_u4_u4_U85 (.ZN( u2_out4_25 ) , .A4( u2_u4_u4_n139 ) , .A3( u2_u4_u4_n140 ) , .A2( u2_u4_u4_n141 ) , .A1( u2_u4_u4_n142 ) );
  OAI21_X1 u2_u4_u4_U86 (.B2( u2_u4_u4_n131 ) , .ZN( u2_u4_u4_n141 ) , .A( u2_u4_u4_n175 ) , .B1( u2_u4_u4_n183 ) );
  OAI21_X1 u2_u4_u4_U87 (.A( u2_u4_u4_n128 ) , .B2( u2_u4_u4_n129 ) , .B1( u2_u4_u4_n130 ) , .ZN( u2_u4_u4_n142 ) );
  NAND4_X1 u2_u4_u4_U88 (.ZN( u2_out4_14 ) , .A4( u2_u4_u4_n124 ) , .A3( u2_u4_u4_n125 ) , .A2( u2_u4_u4_n126 ) , .A1( u2_u4_u4_n127 ) );
  AOI22_X1 u2_u4_u4_U89 (.B2( u2_u4_u4_n117 ) , .ZN( u2_u4_u4_n126 ) , .A1( u2_u4_u4_n129 ) , .B1( u2_u4_u4_n152 ) , .A2( u2_u4_u4_n175 ) );
  AOI211_X1 u2_u4_u4_U9 (.B( u2_u4_u4_n136 ) , .A( u2_u4_u4_n137 ) , .C2( u2_u4_u4_n138 ) , .ZN( u2_u4_u4_n139 ) , .C1( u2_u4_u4_n182 ) );
  AOI22_X1 u2_u4_u4_U90 (.ZN( u2_u4_u4_n125 ) , .B2( u2_u4_u4_n131 ) , .A2( u2_u4_u4_n132 ) , .B1( u2_u4_u4_n138 ) , .A1( u2_u4_u4_n178 ) );
  NAND4_X1 u2_u4_u4_U91 (.ZN( u2_out4_8 ) , .A4( u2_u4_u4_n110 ) , .A3( u2_u4_u4_n111 ) , .A2( u2_u4_u4_n112 ) , .A1( u2_u4_u4_n186 ) );
  NAND2_X1 u2_u4_u4_U92 (.ZN( u2_u4_u4_n112 ) , .A2( u2_u4_u4_n130 ) , .A1( u2_u4_u4_n150 ) );
  AOI22_X1 u2_u4_u4_U93 (.ZN( u2_u4_u4_n111 ) , .B2( u2_u4_u4_n132 ) , .A1( u2_u4_u4_n152 ) , .B1( u2_u4_u4_n178 ) , .A2( u2_u4_u4_n97 ) );
  AOI22_X1 u2_u4_u4_U94 (.B2( u2_u4_u4_n149 ) , .B1( u2_u4_u4_n150 ) , .A2( u2_u4_u4_n151 ) , .A1( u2_u4_u4_n152 ) , .ZN( u2_u4_u4_n167 ) );
  NOR4_X1 u2_u4_u4_U95 (.A4( u2_u4_u4_n162 ) , .A3( u2_u4_u4_n163 ) , .A2( u2_u4_u4_n164 ) , .A1( u2_u4_u4_n165 ) , .ZN( u2_u4_u4_n166 ) );
  NAND3_X1 u2_u4_u4_U96 (.ZN( u2_out4_3 ) , .A3( u2_u4_u4_n166 ) , .A1( u2_u4_u4_n167 ) , .A2( u2_u4_u4_n186 ) );
  NAND3_X1 u2_u4_u4_U97 (.A3( u2_u4_u4_n146 ) , .A2( u2_u4_u4_n147 ) , .A1( u2_u4_u4_n148 ) , .ZN( u2_u4_u4_n149 ) );
  NAND3_X1 u2_u4_u4_U98 (.A3( u2_u4_u4_n143 ) , .A2( u2_u4_u4_n144 ) , .A1( u2_u4_u4_n145 ) , .ZN( u2_u4_u4_n151 ) );
  NAND3_X1 u2_u4_u4_U99 (.A3( u2_u4_u4_n121 ) , .ZN( u2_u4_u4_n122 ) , .A2( u2_u4_u4_n144 ) , .A1( u2_u4_u4_n154 ) );
  NOR2_X1 u2_u4_u5_U10 (.ZN( u2_u4_u5_n135 ) , .A1( u2_u4_u5_n173 ) , .A2( u2_u4_u5_n176 ) );
  NOR3_X1 u2_u4_u5_U100 (.A3( u2_u4_u5_n141 ) , .A1( u2_u4_u5_n142 ) , .ZN( u2_u4_u5_n143 ) , .A2( u2_u4_u5_n191 ) );
  NAND4_X1 u2_u4_u5_U101 (.ZN( u2_out4_4 ) , .A4( u2_u4_u5_n112 ) , .A2( u2_u4_u5_n113 ) , .A1( u2_u4_u5_n114 ) , .A3( u2_u4_u5_n195 ) );
  AOI211_X1 u2_u4_u5_U102 (.A( u2_u4_u5_n110 ) , .C1( u2_u4_u5_n111 ) , .ZN( u2_u4_u5_n112 ) , .B( u2_u4_u5_n118 ) , .C2( u2_u4_u5_n177 ) );
  INV_X1 u2_u4_u5_U103 (.A( u2_u4_u5_n102 ) , .ZN( u2_u4_u5_n195 ) );
  NAND3_X1 u2_u4_u5_U104 (.A2( u2_u4_u5_n154 ) , .A3( u2_u4_u5_n158 ) , .A1( u2_u4_u5_n161 ) , .ZN( u2_u4_u5_n99 ) );
  INV_X1 u2_u4_u5_U11 (.A( u2_u4_u5_n121 ) , .ZN( u2_u4_u5_n177 ) );
  NOR2_X1 u2_u4_u5_U12 (.ZN( u2_u4_u5_n160 ) , .A2( u2_u4_u5_n173 ) , .A1( u2_u4_u5_n177 ) );
  INV_X1 u2_u4_u5_U13 (.A( u2_u4_u5_n150 ) , .ZN( u2_u4_u5_n174 ) );
  AOI21_X1 u2_u4_u5_U14 (.A( u2_u4_u5_n160 ) , .B2( u2_u4_u5_n161 ) , .ZN( u2_u4_u5_n162 ) , .B1( u2_u4_u5_n192 ) );
  INV_X1 u2_u4_u5_U15 (.A( u2_u4_u5_n159 ) , .ZN( u2_u4_u5_n192 ) );
  AOI21_X1 u2_u4_u5_U16 (.A( u2_u4_u5_n156 ) , .B2( u2_u4_u5_n157 ) , .B1( u2_u4_u5_n158 ) , .ZN( u2_u4_u5_n163 ) );
  AOI21_X1 u2_u4_u5_U17 (.B2( u2_u4_u5_n139 ) , .B1( u2_u4_u5_n140 ) , .ZN( u2_u4_u5_n141 ) , .A( u2_u4_u5_n150 ) );
  OAI21_X1 u2_u4_u5_U18 (.A( u2_u4_u5_n133 ) , .B2( u2_u4_u5_n134 ) , .B1( u2_u4_u5_n135 ) , .ZN( u2_u4_u5_n142 ) );
  OAI21_X1 u2_u4_u5_U19 (.ZN( u2_u4_u5_n133 ) , .B2( u2_u4_u5_n147 ) , .A( u2_u4_u5_n173 ) , .B1( u2_u4_u5_n188 ) );
  NAND2_X1 u2_u4_u5_U20 (.A2( u2_u4_u5_n119 ) , .A1( u2_u4_u5_n123 ) , .ZN( u2_u4_u5_n137 ) );
  INV_X1 u2_u4_u5_U21 (.A( u2_u4_u5_n155 ) , .ZN( u2_u4_u5_n194 ) );
  NAND2_X1 u2_u4_u5_U22 (.A1( u2_u4_u5_n121 ) , .ZN( u2_u4_u5_n132 ) , .A2( u2_u4_u5_n172 ) );
  NAND2_X1 u2_u4_u5_U23 (.A2( u2_u4_u5_n122 ) , .ZN( u2_u4_u5_n136 ) , .A1( u2_u4_u5_n154 ) );
  NAND2_X1 u2_u4_u5_U24 (.A2( u2_u4_u5_n119 ) , .A1( u2_u4_u5_n120 ) , .ZN( u2_u4_u5_n159 ) );
  INV_X1 u2_u4_u5_U25 (.A( u2_u4_u5_n156 ) , .ZN( u2_u4_u5_n175 ) );
  INV_X1 u2_u4_u5_U26 (.A( u2_u4_u5_n158 ) , .ZN( u2_u4_u5_n188 ) );
  INV_X1 u2_u4_u5_U27 (.A( u2_u4_u5_n152 ) , .ZN( u2_u4_u5_n179 ) );
  INV_X1 u2_u4_u5_U28 (.A( u2_u4_u5_n140 ) , .ZN( u2_u4_u5_n182 ) );
  INV_X1 u2_u4_u5_U29 (.A( u2_u4_u5_n151 ) , .ZN( u2_u4_u5_n183 ) );
  NOR2_X1 u2_u4_u5_U3 (.ZN( u2_u4_u5_n134 ) , .A1( u2_u4_u5_n183 ) , .A2( u2_u4_u5_n190 ) );
  INV_X1 u2_u4_u5_U30 (.A( u2_u4_u5_n123 ) , .ZN( u2_u4_u5_n185 ) );
  INV_X1 u2_u4_u5_U31 (.A( u2_u4_u5_n161 ) , .ZN( u2_u4_u5_n184 ) );
  INV_X1 u2_u4_u5_U32 (.A( u2_u4_u5_n139 ) , .ZN( u2_u4_u5_n189 ) );
  INV_X1 u2_u4_u5_U33 (.A( u2_u4_u5_n157 ) , .ZN( u2_u4_u5_n190 ) );
  INV_X1 u2_u4_u5_U34 (.A( u2_u4_u5_n120 ) , .ZN( u2_u4_u5_n193 ) );
  NAND2_X1 u2_u4_u5_U35 (.ZN( u2_u4_u5_n111 ) , .A1( u2_u4_u5_n140 ) , .A2( u2_u4_u5_n155 ) );
  INV_X1 u2_u4_u5_U36 (.A( u2_u4_u5_n117 ) , .ZN( u2_u4_u5_n196 ) );
  OAI221_X1 u2_u4_u5_U37 (.A( u2_u4_u5_n116 ) , .ZN( u2_u4_u5_n117 ) , .B2( u2_u4_u5_n119 ) , .C1( u2_u4_u5_n153 ) , .C2( u2_u4_u5_n158 ) , .B1( u2_u4_u5_n172 ) );
  AOI222_X1 u2_u4_u5_U38 (.ZN( u2_u4_u5_n116 ) , .B2( u2_u4_u5_n145 ) , .C1( u2_u4_u5_n148 ) , .A2( u2_u4_u5_n174 ) , .C2( u2_u4_u5_n177 ) , .B1( u2_u4_u5_n187 ) , .A1( u2_u4_u5_n193 ) );
  INV_X1 u2_u4_u5_U39 (.A( u2_u4_u5_n115 ) , .ZN( u2_u4_u5_n187 ) );
  INV_X1 u2_u4_u5_U4 (.A( u2_u4_u5_n138 ) , .ZN( u2_u4_u5_n191 ) );
  NOR2_X1 u2_u4_u5_U40 (.ZN( u2_u4_u5_n100 ) , .A1( u2_u4_u5_n170 ) , .A2( u2_u4_u5_n180 ) );
  OAI221_X1 u2_u4_u5_U41 (.A( u2_u4_u5_n101 ) , .ZN( u2_u4_u5_n102 ) , .C2( u2_u4_u5_n115 ) , .C1( u2_u4_u5_n126 ) , .B1( u2_u4_u5_n134 ) , .B2( u2_u4_u5_n160 ) );
  OAI21_X1 u2_u4_u5_U42 (.ZN( u2_u4_u5_n101 ) , .B1( u2_u4_u5_n137 ) , .A( u2_u4_u5_n146 ) , .B2( u2_u4_u5_n147 ) );
  AOI22_X1 u2_u4_u5_U43 (.B2( u2_u4_u5_n131 ) , .A2( u2_u4_u5_n146 ) , .ZN( u2_u4_u5_n169 ) , .B1( u2_u4_u5_n174 ) , .A1( u2_u4_u5_n185 ) );
  NOR2_X1 u2_u4_u5_U44 (.A1( u2_u4_u5_n146 ) , .ZN( u2_u4_u5_n150 ) , .A2( u2_u4_u5_n173 ) );
  AOI21_X1 u2_u4_u5_U45 (.A( u2_u4_u5_n118 ) , .B2( u2_u4_u5_n145 ) , .ZN( u2_u4_u5_n168 ) , .B1( u2_u4_u5_n186 ) );
  INV_X1 u2_u4_u5_U46 (.A( u2_u4_u5_n122 ) , .ZN( u2_u4_u5_n186 ) );
  NOR2_X1 u2_u4_u5_U47 (.A1( u2_u4_u5_n146 ) , .ZN( u2_u4_u5_n152 ) , .A2( u2_u4_u5_n176 ) );
  NOR2_X1 u2_u4_u5_U48 (.A1( u2_u4_u5_n115 ) , .ZN( u2_u4_u5_n118 ) , .A2( u2_u4_u5_n153 ) );
  NOR2_X1 u2_u4_u5_U49 (.A2( u2_u4_u5_n145 ) , .ZN( u2_u4_u5_n156 ) , .A1( u2_u4_u5_n174 ) );
  OAI21_X1 u2_u4_u5_U5 (.B2( u2_u4_u5_n136 ) , .B1( u2_u4_u5_n137 ) , .ZN( u2_u4_u5_n138 ) , .A( u2_u4_u5_n177 ) );
  NOR2_X1 u2_u4_u5_U50 (.ZN( u2_u4_u5_n121 ) , .A2( u2_u4_u5_n145 ) , .A1( u2_u4_u5_n176 ) );
  AOI22_X1 u2_u4_u5_U51 (.ZN( u2_u4_u5_n114 ) , .A2( u2_u4_u5_n137 ) , .A1( u2_u4_u5_n145 ) , .B2( u2_u4_u5_n175 ) , .B1( u2_u4_u5_n193 ) );
  OAI211_X1 u2_u4_u5_U52 (.B( u2_u4_u5_n124 ) , .A( u2_u4_u5_n125 ) , .C2( u2_u4_u5_n126 ) , .C1( u2_u4_u5_n127 ) , .ZN( u2_u4_u5_n128 ) );
  NOR3_X1 u2_u4_u5_U53 (.ZN( u2_u4_u5_n127 ) , .A1( u2_u4_u5_n136 ) , .A3( u2_u4_u5_n148 ) , .A2( u2_u4_u5_n182 ) );
  OAI21_X1 u2_u4_u5_U54 (.ZN( u2_u4_u5_n124 ) , .A( u2_u4_u5_n177 ) , .B2( u2_u4_u5_n183 ) , .B1( u2_u4_u5_n189 ) );
  OAI21_X1 u2_u4_u5_U55 (.ZN( u2_u4_u5_n125 ) , .A( u2_u4_u5_n174 ) , .B2( u2_u4_u5_n185 ) , .B1( u2_u4_u5_n190 ) );
  AOI21_X1 u2_u4_u5_U56 (.A( u2_u4_u5_n153 ) , .B2( u2_u4_u5_n154 ) , .B1( u2_u4_u5_n155 ) , .ZN( u2_u4_u5_n164 ) );
  AOI21_X1 u2_u4_u5_U57 (.ZN( u2_u4_u5_n110 ) , .B1( u2_u4_u5_n122 ) , .B2( u2_u4_u5_n139 ) , .A( u2_u4_u5_n153 ) );
  INV_X1 u2_u4_u5_U58 (.A( u2_u4_u5_n153 ) , .ZN( u2_u4_u5_n176 ) );
  INV_X1 u2_u4_u5_U59 (.A( u2_u4_u5_n126 ) , .ZN( u2_u4_u5_n173 ) );
  AOI222_X1 u2_u4_u5_U6 (.ZN( u2_u4_u5_n113 ) , .A1( u2_u4_u5_n131 ) , .C1( u2_u4_u5_n148 ) , .B2( u2_u4_u5_n174 ) , .C2( u2_u4_u5_n178 ) , .A2( u2_u4_u5_n179 ) , .B1( u2_u4_u5_n99 ) );
  AND2_X1 u2_u4_u5_U60 (.A2( u2_u4_u5_n104 ) , .A1( u2_u4_u5_n107 ) , .ZN( u2_u4_u5_n147 ) );
  AND2_X1 u2_u4_u5_U61 (.A2( u2_u4_u5_n104 ) , .A1( u2_u4_u5_n108 ) , .ZN( u2_u4_u5_n148 ) );
  NAND2_X1 u2_u4_u5_U62 (.A1( u2_u4_u5_n105 ) , .A2( u2_u4_u5_n106 ) , .ZN( u2_u4_u5_n158 ) );
  NAND2_X1 u2_u4_u5_U63 (.A2( u2_u4_u5_n108 ) , .A1( u2_u4_u5_n109 ) , .ZN( u2_u4_u5_n139 ) );
  NAND2_X1 u2_u4_u5_U64 (.A1( u2_u4_u5_n106 ) , .A2( u2_u4_u5_n108 ) , .ZN( u2_u4_u5_n119 ) );
  NAND2_X1 u2_u4_u5_U65 (.A2( u2_u4_u5_n103 ) , .A1( u2_u4_u5_n105 ) , .ZN( u2_u4_u5_n140 ) );
  NAND2_X1 u2_u4_u5_U66 (.A2( u2_u4_u5_n104 ) , .A1( u2_u4_u5_n105 ) , .ZN( u2_u4_u5_n155 ) );
  NAND2_X1 u2_u4_u5_U67 (.A2( u2_u4_u5_n106 ) , .A1( u2_u4_u5_n107 ) , .ZN( u2_u4_u5_n122 ) );
  NAND2_X1 u2_u4_u5_U68 (.A2( u2_u4_u5_n100 ) , .A1( u2_u4_u5_n106 ) , .ZN( u2_u4_u5_n115 ) );
  NAND2_X1 u2_u4_u5_U69 (.A2( u2_u4_u5_n100 ) , .A1( u2_u4_u5_n103 ) , .ZN( u2_u4_u5_n161 ) );
  INV_X1 u2_u4_u5_U7 (.A( u2_u4_u5_n135 ) , .ZN( u2_u4_u5_n178 ) );
  NAND2_X1 u2_u4_u5_U70 (.A1( u2_u4_u5_n105 ) , .A2( u2_u4_u5_n109 ) , .ZN( u2_u4_u5_n154 ) );
  INV_X1 u2_u4_u5_U71 (.A( u2_u4_u5_n146 ) , .ZN( u2_u4_u5_n172 ) );
  NAND2_X1 u2_u4_u5_U72 (.A1( u2_u4_u5_n103 ) , .A2( u2_u4_u5_n108 ) , .ZN( u2_u4_u5_n123 ) );
  NAND2_X1 u2_u4_u5_U73 (.A2( u2_u4_u5_n103 ) , .A1( u2_u4_u5_n107 ) , .ZN( u2_u4_u5_n151 ) );
  NAND2_X1 u2_u4_u5_U74 (.A2( u2_u4_u5_n107 ) , .A1( u2_u4_u5_n109 ) , .ZN( u2_u4_u5_n120 ) );
  NAND2_X1 u2_u4_u5_U75 (.A2( u2_u4_u5_n100 ) , .A1( u2_u4_u5_n109 ) , .ZN( u2_u4_u5_n157 ) );
  AND2_X1 u2_u4_u5_U76 (.A2( u2_u4_u5_n100 ) , .A1( u2_u4_u5_n104 ) , .ZN( u2_u4_u5_n131 ) );
  NOR2_X1 u2_u4_u5_U77 (.A2( u2_u4_X_34 ) , .A1( u2_u4_X_35 ) , .ZN( u2_u4_u5_n145 ) );
  NOR2_X1 u2_u4_u5_U78 (.A2( u2_u4_X_34 ) , .ZN( u2_u4_u5_n146 ) , .A1( u2_u4_u5_n171 ) );
  NOR2_X1 u2_u4_u5_U79 (.A2( u2_u4_X_31 ) , .A1( u2_u4_X_32 ) , .ZN( u2_u4_u5_n103 ) );
  OAI22_X1 u2_u4_u5_U8 (.B2( u2_u4_u5_n149 ) , .B1( u2_u4_u5_n150 ) , .A2( u2_u4_u5_n151 ) , .A1( u2_u4_u5_n152 ) , .ZN( u2_u4_u5_n165 ) );
  NOR2_X1 u2_u4_u5_U80 (.A2( u2_u4_X_36 ) , .ZN( u2_u4_u5_n105 ) , .A1( u2_u4_u5_n180 ) );
  NOR2_X1 u2_u4_u5_U81 (.A2( u2_u4_X_33 ) , .ZN( u2_u4_u5_n108 ) , .A1( u2_u4_u5_n170 ) );
  NOR2_X1 u2_u4_u5_U82 (.A2( u2_u4_X_33 ) , .A1( u2_u4_X_36 ) , .ZN( u2_u4_u5_n107 ) );
  NOR2_X1 u2_u4_u5_U83 (.A2( u2_u4_X_31 ) , .ZN( u2_u4_u5_n104 ) , .A1( u2_u4_u5_n181 ) );
  NAND2_X1 u2_u4_u5_U84 (.A2( u2_u4_X_34 ) , .A1( u2_u4_X_35 ) , .ZN( u2_u4_u5_n153 ) );
  NAND2_X1 u2_u4_u5_U85 (.A1( u2_u4_X_34 ) , .ZN( u2_u4_u5_n126 ) , .A2( u2_u4_u5_n171 ) );
  AND2_X1 u2_u4_u5_U86 (.A1( u2_u4_X_31 ) , .A2( u2_u4_X_32 ) , .ZN( u2_u4_u5_n106 ) );
  AND2_X1 u2_u4_u5_U87 (.A1( u2_u4_X_31 ) , .ZN( u2_u4_u5_n109 ) , .A2( u2_u4_u5_n181 ) );
  INV_X1 u2_u4_u5_U88 (.A( u2_u4_X_33 ) , .ZN( u2_u4_u5_n180 ) );
  INV_X1 u2_u4_u5_U89 (.A( u2_u4_X_35 ) , .ZN( u2_u4_u5_n171 ) );
  NOR3_X1 u2_u4_u5_U9 (.A2( u2_u4_u5_n147 ) , .A1( u2_u4_u5_n148 ) , .ZN( u2_u4_u5_n149 ) , .A3( u2_u4_u5_n194 ) );
  INV_X1 u2_u4_u5_U90 (.A( u2_u4_X_36 ) , .ZN( u2_u4_u5_n170 ) );
  INV_X1 u2_u4_u5_U91 (.A( u2_u4_X_32 ) , .ZN( u2_u4_u5_n181 ) );
  NAND4_X1 u2_u4_u5_U92 (.ZN( u2_out4_29 ) , .A4( u2_u4_u5_n129 ) , .A3( u2_u4_u5_n130 ) , .A2( u2_u4_u5_n168 ) , .A1( u2_u4_u5_n196 ) );
  AOI221_X1 u2_u4_u5_U93 (.A( u2_u4_u5_n128 ) , .ZN( u2_u4_u5_n129 ) , .C2( u2_u4_u5_n132 ) , .B2( u2_u4_u5_n159 ) , .B1( u2_u4_u5_n176 ) , .C1( u2_u4_u5_n184 ) );
  AOI222_X1 u2_u4_u5_U94 (.ZN( u2_u4_u5_n130 ) , .A2( u2_u4_u5_n146 ) , .B1( u2_u4_u5_n147 ) , .C2( u2_u4_u5_n175 ) , .B2( u2_u4_u5_n179 ) , .A1( u2_u4_u5_n188 ) , .C1( u2_u4_u5_n194 ) );
  NAND4_X1 u2_u4_u5_U95 (.ZN( u2_out4_19 ) , .A4( u2_u4_u5_n166 ) , .A3( u2_u4_u5_n167 ) , .A2( u2_u4_u5_n168 ) , .A1( u2_u4_u5_n169 ) );
  AOI22_X1 u2_u4_u5_U96 (.B2( u2_u4_u5_n145 ) , .A2( u2_u4_u5_n146 ) , .ZN( u2_u4_u5_n167 ) , .B1( u2_u4_u5_n182 ) , .A1( u2_u4_u5_n189 ) );
  NOR4_X1 u2_u4_u5_U97 (.A4( u2_u4_u5_n162 ) , .A3( u2_u4_u5_n163 ) , .A2( u2_u4_u5_n164 ) , .A1( u2_u4_u5_n165 ) , .ZN( u2_u4_u5_n166 ) );
  NAND4_X1 u2_u4_u5_U98 (.ZN( u2_out4_11 ) , .A4( u2_u4_u5_n143 ) , .A3( u2_u4_u5_n144 ) , .A2( u2_u4_u5_n169 ) , .A1( u2_u4_u5_n196 ) );
  AOI22_X1 u2_u4_u5_U99 (.A2( u2_u4_u5_n132 ) , .ZN( u2_u4_u5_n144 ) , .B2( u2_u4_u5_n145 ) , .B1( u2_u4_u5_n184 ) , .A1( u2_u4_u5_n194 ) );
  AOI22_X1 u2_u4_u6_U10 (.A2( u2_u4_u6_n151 ) , .B2( u2_u4_u6_n161 ) , .A1( u2_u4_u6_n167 ) , .B1( u2_u4_u6_n170 ) , .ZN( u2_u4_u6_n89 ) );
  AOI21_X1 u2_u4_u6_U11 (.B1( u2_u4_u6_n107 ) , .B2( u2_u4_u6_n132 ) , .A( u2_u4_u6_n158 ) , .ZN( u2_u4_u6_n88 ) );
  AOI21_X1 u2_u4_u6_U12 (.B2( u2_u4_u6_n147 ) , .B1( u2_u4_u6_n148 ) , .ZN( u2_u4_u6_n149 ) , .A( u2_u4_u6_n158 ) );
  AOI21_X1 u2_u4_u6_U13 (.ZN( u2_u4_u6_n106 ) , .A( u2_u4_u6_n142 ) , .B2( u2_u4_u6_n159 ) , .B1( u2_u4_u6_n164 ) );
  INV_X1 u2_u4_u6_U14 (.A( u2_u4_u6_n155 ) , .ZN( u2_u4_u6_n161 ) );
  INV_X1 u2_u4_u6_U15 (.A( u2_u4_u6_n128 ) , .ZN( u2_u4_u6_n164 ) );
  NAND2_X1 u2_u4_u6_U16 (.ZN( u2_u4_u6_n110 ) , .A1( u2_u4_u6_n122 ) , .A2( u2_u4_u6_n129 ) );
  NAND2_X1 u2_u4_u6_U17 (.ZN( u2_u4_u6_n124 ) , .A2( u2_u4_u6_n146 ) , .A1( u2_u4_u6_n148 ) );
  INV_X1 u2_u4_u6_U18 (.A( u2_u4_u6_n132 ) , .ZN( u2_u4_u6_n171 ) );
  AND2_X1 u2_u4_u6_U19 (.A1( u2_u4_u6_n100 ) , .ZN( u2_u4_u6_n130 ) , .A2( u2_u4_u6_n147 ) );
  INV_X1 u2_u4_u6_U20 (.A( u2_u4_u6_n127 ) , .ZN( u2_u4_u6_n173 ) );
  INV_X1 u2_u4_u6_U21 (.A( u2_u4_u6_n121 ) , .ZN( u2_u4_u6_n167 ) );
  INV_X1 u2_u4_u6_U22 (.A( u2_u4_u6_n100 ) , .ZN( u2_u4_u6_n169 ) );
  INV_X1 u2_u4_u6_U23 (.A( u2_u4_u6_n123 ) , .ZN( u2_u4_u6_n170 ) );
  INV_X1 u2_u4_u6_U24 (.A( u2_u4_u6_n113 ) , .ZN( u2_u4_u6_n168 ) );
  AND2_X1 u2_u4_u6_U25 (.A1( u2_u4_u6_n107 ) , .A2( u2_u4_u6_n119 ) , .ZN( u2_u4_u6_n133 ) );
  AND2_X1 u2_u4_u6_U26 (.A2( u2_u4_u6_n121 ) , .A1( u2_u4_u6_n122 ) , .ZN( u2_u4_u6_n131 ) );
  AND3_X1 u2_u4_u6_U27 (.ZN( u2_u4_u6_n120 ) , .A2( u2_u4_u6_n127 ) , .A1( u2_u4_u6_n132 ) , .A3( u2_u4_u6_n145 ) );
  INV_X1 u2_u4_u6_U28 (.A( u2_u4_u6_n146 ) , .ZN( u2_u4_u6_n163 ) );
  AOI222_X1 u2_u4_u6_U29 (.ZN( u2_u4_u6_n114 ) , .A1( u2_u4_u6_n118 ) , .A2( u2_u4_u6_n126 ) , .B2( u2_u4_u6_n151 ) , .C2( u2_u4_u6_n159 ) , .C1( u2_u4_u6_n168 ) , .B1( u2_u4_u6_n169 ) );
  INV_X1 u2_u4_u6_U3 (.A( u2_u4_u6_n110 ) , .ZN( u2_u4_u6_n166 ) );
  NOR2_X1 u2_u4_u6_U30 (.A1( u2_u4_u6_n162 ) , .A2( u2_u4_u6_n165 ) , .ZN( u2_u4_u6_n98 ) );
  NAND2_X1 u2_u4_u6_U31 (.A1( u2_u4_u6_n144 ) , .ZN( u2_u4_u6_n151 ) , .A2( u2_u4_u6_n158 ) );
  NAND2_X1 u2_u4_u6_U32 (.ZN( u2_u4_u6_n132 ) , .A1( u2_u4_u6_n91 ) , .A2( u2_u4_u6_n97 ) );
  AOI22_X1 u2_u4_u6_U33 (.B2( u2_u4_u6_n110 ) , .B1( u2_u4_u6_n111 ) , .A1( u2_u4_u6_n112 ) , .ZN( u2_u4_u6_n115 ) , .A2( u2_u4_u6_n161 ) );
  NAND4_X1 u2_u4_u6_U34 (.A3( u2_u4_u6_n109 ) , .ZN( u2_u4_u6_n112 ) , .A4( u2_u4_u6_n132 ) , .A2( u2_u4_u6_n147 ) , .A1( u2_u4_u6_n166 ) );
  NOR2_X1 u2_u4_u6_U35 (.ZN( u2_u4_u6_n109 ) , .A1( u2_u4_u6_n170 ) , .A2( u2_u4_u6_n173 ) );
  NOR2_X1 u2_u4_u6_U36 (.A2( u2_u4_u6_n126 ) , .ZN( u2_u4_u6_n155 ) , .A1( u2_u4_u6_n160 ) );
  NAND2_X1 u2_u4_u6_U37 (.ZN( u2_u4_u6_n146 ) , .A2( u2_u4_u6_n94 ) , .A1( u2_u4_u6_n99 ) );
  AOI21_X1 u2_u4_u6_U38 (.A( u2_u4_u6_n144 ) , .B2( u2_u4_u6_n145 ) , .B1( u2_u4_u6_n146 ) , .ZN( u2_u4_u6_n150 ) );
  AOI211_X1 u2_u4_u6_U39 (.B( u2_u4_u6_n134 ) , .A( u2_u4_u6_n135 ) , .C1( u2_u4_u6_n136 ) , .ZN( u2_u4_u6_n137 ) , .C2( u2_u4_u6_n151 ) );
  INV_X1 u2_u4_u6_U4 (.A( u2_u4_u6_n142 ) , .ZN( u2_u4_u6_n174 ) );
  NAND4_X1 u2_u4_u6_U40 (.A4( u2_u4_u6_n127 ) , .A3( u2_u4_u6_n128 ) , .A2( u2_u4_u6_n129 ) , .A1( u2_u4_u6_n130 ) , .ZN( u2_u4_u6_n136 ) );
  AOI21_X1 u2_u4_u6_U41 (.B2( u2_u4_u6_n132 ) , .B1( u2_u4_u6_n133 ) , .ZN( u2_u4_u6_n134 ) , .A( u2_u4_u6_n158 ) );
  AOI21_X1 u2_u4_u6_U42 (.B1( u2_u4_u6_n131 ) , .ZN( u2_u4_u6_n135 ) , .A( u2_u4_u6_n144 ) , .B2( u2_u4_u6_n146 ) );
  INV_X1 u2_u4_u6_U43 (.A( u2_u4_u6_n111 ) , .ZN( u2_u4_u6_n158 ) );
  NAND2_X1 u2_u4_u6_U44 (.ZN( u2_u4_u6_n127 ) , .A1( u2_u4_u6_n91 ) , .A2( u2_u4_u6_n92 ) );
  NAND2_X1 u2_u4_u6_U45 (.ZN( u2_u4_u6_n129 ) , .A2( u2_u4_u6_n95 ) , .A1( u2_u4_u6_n96 ) );
  INV_X1 u2_u4_u6_U46 (.A( u2_u4_u6_n144 ) , .ZN( u2_u4_u6_n159 ) );
  NAND2_X1 u2_u4_u6_U47 (.ZN( u2_u4_u6_n145 ) , .A2( u2_u4_u6_n97 ) , .A1( u2_u4_u6_n98 ) );
  NAND2_X1 u2_u4_u6_U48 (.ZN( u2_u4_u6_n148 ) , .A2( u2_u4_u6_n92 ) , .A1( u2_u4_u6_n94 ) );
  NAND2_X1 u2_u4_u6_U49 (.ZN( u2_u4_u6_n108 ) , .A2( u2_u4_u6_n139 ) , .A1( u2_u4_u6_n144 ) );
  NAND2_X1 u2_u4_u6_U5 (.A2( u2_u4_u6_n143 ) , .ZN( u2_u4_u6_n152 ) , .A1( u2_u4_u6_n166 ) );
  NAND2_X1 u2_u4_u6_U50 (.ZN( u2_u4_u6_n121 ) , .A2( u2_u4_u6_n95 ) , .A1( u2_u4_u6_n97 ) );
  NAND2_X1 u2_u4_u6_U51 (.ZN( u2_u4_u6_n107 ) , .A2( u2_u4_u6_n92 ) , .A1( u2_u4_u6_n95 ) );
  AND2_X1 u2_u4_u6_U52 (.ZN( u2_u4_u6_n118 ) , .A2( u2_u4_u6_n91 ) , .A1( u2_u4_u6_n99 ) );
  NAND2_X1 u2_u4_u6_U53 (.ZN( u2_u4_u6_n147 ) , .A2( u2_u4_u6_n98 ) , .A1( u2_u4_u6_n99 ) );
  NAND2_X1 u2_u4_u6_U54 (.ZN( u2_u4_u6_n128 ) , .A1( u2_u4_u6_n94 ) , .A2( u2_u4_u6_n96 ) );
  NAND2_X1 u2_u4_u6_U55 (.ZN( u2_u4_u6_n119 ) , .A2( u2_u4_u6_n95 ) , .A1( u2_u4_u6_n99 ) );
  NAND2_X1 u2_u4_u6_U56 (.ZN( u2_u4_u6_n123 ) , .A2( u2_u4_u6_n91 ) , .A1( u2_u4_u6_n96 ) );
  NAND2_X1 u2_u4_u6_U57 (.ZN( u2_u4_u6_n100 ) , .A2( u2_u4_u6_n92 ) , .A1( u2_u4_u6_n98 ) );
  NAND2_X1 u2_u4_u6_U58 (.ZN( u2_u4_u6_n122 ) , .A1( u2_u4_u6_n94 ) , .A2( u2_u4_u6_n97 ) );
  INV_X1 u2_u4_u6_U59 (.A( u2_u4_u6_n139 ) , .ZN( u2_u4_u6_n160 ) );
  AOI22_X1 u2_u4_u6_U6 (.B2( u2_u4_u6_n101 ) , .A1( u2_u4_u6_n102 ) , .ZN( u2_u4_u6_n103 ) , .B1( u2_u4_u6_n160 ) , .A2( u2_u4_u6_n161 ) );
  NAND2_X1 u2_u4_u6_U60 (.ZN( u2_u4_u6_n113 ) , .A1( u2_u4_u6_n96 ) , .A2( u2_u4_u6_n98 ) );
  NOR2_X1 u2_u4_u6_U61 (.A2( u2_u4_X_40 ) , .A1( u2_u4_X_41 ) , .ZN( u2_u4_u6_n126 ) );
  NOR2_X1 u2_u4_u6_U62 (.A2( u2_u4_X_39 ) , .A1( u2_u4_X_42 ) , .ZN( u2_u4_u6_n92 ) );
  NOR2_X1 u2_u4_u6_U63 (.A2( u2_u4_X_39 ) , .A1( u2_u4_u6_n156 ) , .ZN( u2_u4_u6_n97 ) );
  NOR2_X1 u2_u4_u6_U64 (.A2( u2_u4_X_38 ) , .A1( u2_u4_u6_n165 ) , .ZN( u2_u4_u6_n95 ) );
  NOR2_X1 u2_u4_u6_U65 (.A2( u2_u4_X_41 ) , .ZN( u2_u4_u6_n111 ) , .A1( u2_u4_u6_n157 ) );
  NOR2_X1 u2_u4_u6_U66 (.A2( u2_u4_X_37 ) , .A1( u2_u4_u6_n162 ) , .ZN( u2_u4_u6_n94 ) );
  NOR2_X1 u2_u4_u6_U67 (.A2( u2_u4_X_37 ) , .A1( u2_u4_X_38 ) , .ZN( u2_u4_u6_n91 ) );
  NAND2_X1 u2_u4_u6_U68 (.A1( u2_u4_X_41 ) , .ZN( u2_u4_u6_n144 ) , .A2( u2_u4_u6_n157 ) );
  NAND2_X1 u2_u4_u6_U69 (.A2( u2_u4_X_40 ) , .A1( u2_u4_X_41 ) , .ZN( u2_u4_u6_n139 ) );
  NOR2_X1 u2_u4_u6_U7 (.A1( u2_u4_u6_n118 ) , .ZN( u2_u4_u6_n143 ) , .A2( u2_u4_u6_n168 ) );
  AND2_X1 u2_u4_u6_U70 (.A1( u2_u4_X_39 ) , .A2( u2_u4_u6_n156 ) , .ZN( u2_u4_u6_n96 ) );
  AND2_X1 u2_u4_u6_U71 (.A1( u2_u4_X_39 ) , .A2( u2_u4_X_42 ) , .ZN( u2_u4_u6_n99 ) );
  INV_X1 u2_u4_u6_U72 (.A( u2_u4_X_40 ) , .ZN( u2_u4_u6_n157 ) );
  INV_X1 u2_u4_u6_U73 (.A( u2_u4_X_37 ) , .ZN( u2_u4_u6_n165 ) );
  INV_X1 u2_u4_u6_U74 (.A( u2_u4_X_38 ) , .ZN( u2_u4_u6_n162 ) );
  INV_X1 u2_u4_u6_U75 (.A( u2_u4_X_42 ) , .ZN( u2_u4_u6_n156 ) );
  NAND4_X1 u2_u4_u6_U76 (.ZN( u2_out4_32 ) , .A4( u2_u4_u6_n103 ) , .A3( u2_u4_u6_n104 ) , .A2( u2_u4_u6_n105 ) , .A1( u2_u4_u6_n106 ) );
  AOI22_X1 u2_u4_u6_U77 (.ZN( u2_u4_u6_n105 ) , .A2( u2_u4_u6_n108 ) , .A1( u2_u4_u6_n118 ) , .B2( u2_u4_u6_n126 ) , .B1( u2_u4_u6_n171 ) );
  AOI22_X1 u2_u4_u6_U78 (.ZN( u2_u4_u6_n104 ) , .A1( u2_u4_u6_n111 ) , .B1( u2_u4_u6_n124 ) , .B2( u2_u4_u6_n151 ) , .A2( u2_u4_u6_n93 ) );
  NAND4_X1 u2_u4_u6_U79 (.ZN( u2_out4_12 ) , .A4( u2_u4_u6_n114 ) , .A3( u2_u4_u6_n115 ) , .A2( u2_u4_u6_n116 ) , .A1( u2_u4_u6_n117 ) );
  INV_X1 u2_u4_u6_U8 (.ZN( u2_u4_u6_n172 ) , .A( u2_u4_u6_n88 ) );
  OAI22_X1 u2_u4_u6_U80 (.B2( u2_u4_u6_n111 ) , .ZN( u2_u4_u6_n116 ) , .B1( u2_u4_u6_n126 ) , .A2( u2_u4_u6_n164 ) , .A1( u2_u4_u6_n167 ) );
  OAI21_X1 u2_u4_u6_U81 (.A( u2_u4_u6_n108 ) , .ZN( u2_u4_u6_n117 ) , .B2( u2_u4_u6_n141 ) , .B1( u2_u4_u6_n163 ) );
  OAI211_X1 u2_u4_u6_U82 (.ZN( u2_out4_22 ) , .B( u2_u4_u6_n137 ) , .A( u2_u4_u6_n138 ) , .C2( u2_u4_u6_n139 ) , .C1( u2_u4_u6_n140 ) );
  AOI22_X1 u2_u4_u6_U83 (.B1( u2_u4_u6_n124 ) , .A2( u2_u4_u6_n125 ) , .A1( u2_u4_u6_n126 ) , .ZN( u2_u4_u6_n138 ) , .B2( u2_u4_u6_n161 ) );
  AND4_X1 u2_u4_u6_U84 (.A3( u2_u4_u6_n119 ) , .A1( u2_u4_u6_n120 ) , .A4( u2_u4_u6_n129 ) , .ZN( u2_u4_u6_n140 ) , .A2( u2_u4_u6_n143 ) );
  OAI211_X1 u2_u4_u6_U85 (.ZN( u2_out4_7 ) , .B( u2_u4_u6_n153 ) , .C2( u2_u4_u6_n154 ) , .C1( u2_u4_u6_n155 ) , .A( u2_u4_u6_n174 ) );
  NOR3_X1 u2_u4_u6_U86 (.A1( u2_u4_u6_n141 ) , .ZN( u2_u4_u6_n154 ) , .A3( u2_u4_u6_n164 ) , .A2( u2_u4_u6_n171 ) );
  AOI211_X1 u2_u4_u6_U87 (.B( u2_u4_u6_n149 ) , .A( u2_u4_u6_n150 ) , .C2( u2_u4_u6_n151 ) , .C1( u2_u4_u6_n152 ) , .ZN( u2_u4_u6_n153 ) );
  NAND3_X1 u2_u4_u6_U88 (.A2( u2_u4_u6_n123 ) , .ZN( u2_u4_u6_n125 ) , .A1( u2_u4_u6_n130 ) , .A3( u2_u4_u6_n131 ) );
  NAND3_X1 u2_u4_u6_U89 (.A3( u2_u4_u6_n133 ) , .ZN( u2_u4_u6_n141 ) , .A1( u2_u4_u6_n145 ) , .A2( u2_u4_u6_n148 ) );
  OAI21_X1 u2_u4_u6_U9 (.A( u2_u4_u6_n159 ) , .B1( u2_u4_u6_n169 ) , .B2( u2_u4_u6_n173 ) , .ZN( u2_u4_u6_n90 ) );
  NAND3_X1 u2_u4_u6_U90 (.ZN( u2_u4_u6_n101 ) , .A3( u2_u4_u6_n107 ) , .A2( u2_u4_u6_n121 ) , .A1( u2_u4_u6_n127 ) );
  NAND3_X1 u2_u4_u6_U91 (.ZN( u2_u4_u6_n102 ) , .A3( u2_u4_u6_n130 ) , .A2( u2_u4_u6_n145 ) , .A1( u2_u4_u6_n166 ) );
  NAND3_X1 u2_u4_u6_U92 (.A3( u2_u4_u6_n113 ) , .A1( u2_u4_u6_n119 ) , .A2( u2_u4_u6_n123 ) , .ZN( u2_u4_u6_n93 ) );
  NAND3_X1 u2_u4_u6_U93 (.ZN( u2_u4_u6_n142 ) , .A2( u2_u4_u6_n172 ) , .A3( u2_u4_u6_n89 ) , .A1( u2_u4_u6_n90 ) );
  AND3_X1 u2_u4_u7_U10 (.A3( u2_u4_u7_n110 ) , .A2( u2_u4_u7_n127 ) , .A1( u2_u4_u7_n132 ) , .ZN( u2_u4_u7_n92 ) );
  OAI21_X1 u2_u4_u7_U11 (.A( u2_u4_u7_n161 ) , .B1( u2_u4_u7_n168 ) , .B2( u2_u4_u7_n173 ) , .ZN( u2_u4_u7_n91 ) );
  AOI211_X1 u2_u4_u7_U12 (.A( u2_u4_u7_n117 ) , .ZN( u2_u4_u7_n118 ) , .C2( u2_u4_u7_n126 ) , .C1( u2_u4_u7_n177 ) , .B( u2_u4_u7_n180 ) );
  OAI22_X1 u2_u4_u7_U13 (.B1( u2_u4_u7_n115 ) , .ZN( u2_u4_u7_n117 ) , .A2( u2_u4_u7_n133 ) , .A1( u2_u4_u7_n137 ) , .B2( u2_u4_u7_n162 ) );
  INV_X1 u2_u4_u7_U14 (.A( u2_u4_u7_n116 ) , .ZN( u2_u4_u7_n180 ) );
  NOR3_X1 u2_u4_u7_U15 (.ZN( u2_u4_u7_n115 ) , .A3( u2_u4_u7_n145 ) , .A2( u2_u4_u7_n168 ) , .A1( u2_u4_u7_n169 ) );
  NOR3_X1 u2_u4_u7_U16 (.A2( u2_u4_u7_n134 ) , .A1( u2_u4_u7_n135 ) , .ZN( u2_u4_u7_n136 ) , .A3( u2_u4_u7_n171 ) );
  NOR2_X1 u2_u4_u7_U17 (.A1( u2_u4_u7_n130 ) , .A2( u2_u4_u7_n134 ) , .ZN( u2_u4_u7_n153 ) );
  NOR2_X1 u2_u4_u7_U18 (.ZN( u2_u4_u7_n111 ) , .A2( u2_u4_u7_n134 ) , .A1( u2_u4_u7_n169 ) );
  AOI21_X1 u2_u4_u7_U19 (.ZN( u2_u4_u7_n104 ) , .B2( u2_u4_u7_n112 ) , .B1( u2_u4_u7_n127 ) , .A( u2_u4_u7_n164 ) );
  AOI21_X1 u2_u4_u7_U20 (.ZN( u2_u4_u7_n106 ) , .B1( u2_u4_u7_n133 ) , .B2( u2_u4_u7_n146 ) , .A( u2_u4_u7_n162 ) );
  AOI21_X1 u2_u4_u7_U21 (.A( u2_u4_u7_n101 ) , .ZN( u2_u4_u7_n107 ) , .B2( u2_u4_u7_n128 ) , .B1( u2_u4_u7_n175 ) );
  INV_X1 u2_u4_u7_U22 (.A( u2_u4_u7_n101 ) , .ZN( u2_u4_u7_n165 ) );
  INV_X1 u2_u4_u7_U23 (.A( u2_u4_u7_n138 ) , .ZN( u2_u4_u7_n171 ) );
  INV_X1 u2_u4_u7_U24 (.A( u2_u4_u7_n131 ) , .ZN( u2_u4_u7_n177 ) );
  INV_X1 u2_u4_u7_U25 (.A( u2_u4_u7_n110 ) , .ZN( u2_u4_u7_n174 ) );
  NAND2_X1 u2_u4_u7_U26 (.A1( u2_u4_u7_n129 ) , .A2( u2_u4_u7_n132 ) , .ZN( u2_u4_u7_n149 ) );
  NAND2_X1 u2_u4_u7_U27 (.A1( u2_u4_u7_n113 ) , .A2( u2_u4_u7_n124 ) , .ZN( u2_u4_u7_n130 ) );
  INV_X1 u2_u4_u7_U28 (.A( u2_u4_u7_n128 ) , .ZN( u2_u4_u7_n168 ) );
  INV_X1 u2_u4_u7_U29 (.A( u2_u4_u7_n148 ) , .ZN( u2_u4_u7_n169 ) );
  INV_X1 u2_u4_u7_U3 (.A( u2_u4_u7_n149 ) , .ZN( u2_u4_u7_n175 ) );
  INV_X1 u2_u4_u7_U30 (.A( u2_u4_u7_n112 ) , .ZN( u2_u4_u7_n173 ) );
  INV_X1 u2_u4_u7_U31 (.A( u2_u4_u7_n127 ) , .ZN( u2_u4_u7_n179 ) );
  NOR2_X1 u2_u4_u7_U32 (.ZN( u2_u4_u7_n101 ) , .A2( u2_u4_u7_n150 ) , .A1( u2_u4_u7_n156 ) );
  AOI211_X1 u2_u4_u7_U33 (.B( u2_u4_u7_n154 ) , .A( u2_u4_u7_n155 ) , .C1( u2_u4_u7_n156 ) , .ZN( u2_u4_u7_n157 ) , .C2( u2_u4_u7_n172 ) );
  INV_X1 u2_u4_u7_U34 (.A( u2_u4_u7_n153 ) , .ZN( u2_u4_u7_n172 ) );
  AOI211_X1 u2_u4_u7_U35 (.B( u2_u4_u7_n139 ) , .A( u2_u4_u7_n140 ) , .C2( u2_u4_u7_n141 ) , .ZN( u2_u4_u7_n142 ) , .C1( u2_u4_u7_n156 ) );
  NAND4_X1 u2_u4_u7_U36 (.A3( u2_u4_u7_n127 ) , .A2( u2_u4_u7_n128 ) , .A1( u2_u4_u7_n129 ) , .ZN( u2_u4_u7_n141 ) , .A4( u2_u4_u7_n147 ) );
  AOI21_X1 u2_u4_u7_U37 (.A( u2_u4_u7_n137 ) , .B1( u2_u4_u7_n138 ) , .ZN( u2_u4_u7_n139 ) , .B2( u2_u4_u7_n146 ) );
  OAI22_X1 u2_u4_u7_U38 (.B1( u2_u4_u7_n136 ) , .ZN( u2_u4_u7_n140 ) , .A1( u2_u4_u7_n153 ) , .B2( u2_u4_u7_n162 ) , .A2( u2_u4_u7_n164 ) );
  INV_X1 u2_u4_u7_U39 (.A( u2_u4_u7_n125 ) , .ZN( u2_u4_u7_n161 ) );
  INV_X1 u2_u4_u7_U4 (.A( u2_u4_u7_n154 ) , .ZN( u2_u4_u7_n178 ) );
  AOI21_X1 u2_u4_u7_U40 (.ZN( u2_u4_u7_n123 ) , .B1( u2_u4_u7_n165 ) , .B2( u2_u4_u7_n177 ) , .A( u2_u4_u7_n97 ) );
  AOI21_X1 u2_u4_u7_U41 (.B2( u2_u4_u7_n113 ) , .B1( u2_u4_u7_n124 ) , .A( u2_u4_u7_n125 ) , .ZN( u2_u4_u7_n97 ) );
  INV_X1 u2_u4_u7_U42 (.A( u2_u4_u7_n152 ) , .ZN( u2_u4_u7_n162 ) );
  AOI22_X1 u2_u4_u7_U43 (.A2( u2_u4_u7_n114 ) , .ZN( u2_u4_u7_n119 ) , .B1( u2_u4_u7_n130 ) , .A1( u2_u4_u7_n156 ) , .B2( u2_u4_u7_n165 ) );
  NAND2_X1 u2_u4_u7_U44 (.A2( u2_u4_u7_n112 ) , .ZN( u2_u4_u7_n114 ) , .A1( u2_u4_u7_n175 ) );
  AOI22_X1 u2_u4_u7_U45 (.B2( u2_u4_u7_n149 ) , .B1( u2_u4_u7_n150 ) , .A2( u2_u4_u7_n151 ) , .A1( u2_u4_u7_n152 ) , .ZN( u2_u4_u7_n158 ) );
  NOR2_X1 u2_u4_u7_U46 (.ZN( u2_u4_u7_n137 ) , .A1( u2_u4_u7_n150 ) , .A2( u2_u4_u7_n161 ) );
  AND2_X1 u2_u4_u7_U47 (.ZN( u2_u4_u7_n145 ) , .A2( u2_u4_u7_n98 ) , .A1( u2_u4_u7_n99 ) );
  AOI21_X1 u2_u4_u7_U48 (.ZN( u2_u4_u7_n105 ) , .B2( u2_u4_u7_n110 ) , .A( u2_u4_u7_n125 ) , .B1( u2_u4_u7_n147 ) );
  NAND2_X1 u2_u4_u7_U49 (.ZN( u2_u4_u7_n146 ) , .A1( u2_u4_u7_n95 ) , .A2( u2_u4_u7_n98 ) );
  INV_X1 u2_u4_u7_U5 (.A( u2_u4_u7_n111 ) , .ZN( u2_u4_u7_n170 ) );
  NAND2_X1 u2_u4_u7_U50 (.A2( u2_u4_u7_n103 ) , .ZN( u2_u4_u7_n147 ) , .A1( u2_u4_u7_n93 ) );
  NAND2_X1 u2_u4_u7_U51 (.A1( u2_u4_u7_n103 ) , .ZN( u2_u4_u7_n127 ) , .A2( u2_u4_u7_n99 ) );
  NAND2_X1 u2_u4_u7_U52 (.A2( u2_u4_u7_n102 ) , .A1( u2_u4_u7_n103 ) , .ZN( u2_u4_u7_n133 ) );
  OR2_X1 u2_u4_u7_U53 (.ZN( u2_u4_u7_n126 ) , .A2( u2_u4_u7_n152 ) , .A1( u2_u4_u7_n156 ) );
  NAND2_X1 u2_u4_u7_U54 (.ZN( u2_u4_u7_n112 ) , .A2( u2_u4_u7_n96 ) , .A1( u2_u4_u7_n99 ) );
  NAND2_X1 u2_u4_u7_U55 (.A2( u2_u4_u7_n102 ) , .ZN( u2_u4_u7_n128 ) , .A1( u2_u4_u7_n98 ) );
  INV_X1 u2_u4_u7_U56 (.A( u2_u4_u7_n150 ) , .ZN( u2_u4_u7_n164 ) );
  AND2_X1 u2_u4_u7_U57 (.ZN( u2_u4_u7_n134 ) , .A1( u2_u4_u7_n93 ) , .A2( u2_u4_u7_n98 ) );
  NAND2_X1 u2_u4_u7_U58 (.ZN( u2_u4_u7_n110 ) , .A1( u2_u4_u7_n95 ) , .A2( u2_u4_u7_n96 ) );
  NAND2_X1 u2_u4_u7_U59 (.A2( u2_u4_u7_n102 ) , .ZN( u2_u4_u7_n124 ) , .A1( u2_u4_u7_n96 ) );
  AOI211_X1 u2_u4_u7_U6 (.ZN( u2_u4_u7_n116 ) , .A( u2_u4_u7_n155 ) , .C1( u2_u4_u7_n161 ) , .C2( u2_u4_u7_n171 ) , .B( u2_u4_u7_n94 ) );
  NAND2_X1 u2_u4_u7_U60 (.ZN( u2_u4_u7_n132 ) , .A1( u2_u4_u7_n93 ) , .A2( u2_u4_u7_n96 ) );
  NAND2_X1 u2_u4_u7_U61 (.A2( u2_u4_u7_n103 ) , .ZN( u2_u4_u7_n131 ) , .A1( u2_u4_u7_n95 ) );
  NOR2_X1 u2_u4_u7_U62 (.A2( u2_u4_X_47 ) , .ZN( u2_u4_u7_n150 ) , .A1( u2_u4_u7_n163 ) );
  NOR2_X1 u2_u4_u7_U63 (.A2( u2_u4_X_43 ) , .A1( u2_u4_X_44 ) , .ZN( u2_u4_u7_n103 ) );
  NOR2_X1 u2_u4_u7_U64 (.A2( u2_u4_X_48 ) , .A1( u2_u4_u7_n166 ) , .ZN( u2_u4_u7_n95 ) );
  NOR2_X1 u2_u4_u7_U65 (.A2( u2_u4_X_44 ) , .A1( u2_u4_u7_n167 ) , .ZN( u2_u4_u7_n98 ) );
  NOR2_X1 u2_u4_u7_U66 (.A2( u2_u4_X_45 ) , .A1( u2_u4_X_48 ) , .ZN( u2_u4_u7_n99 ) );
  NOR2_X1 u2_u4_u7_U67 (.A2( u2_u4_X_46 ) , .A1( u2_u4_X_47 ) , .ZN( u2_u4_u7_n152 ) );
  AND2_X1 u2_u4_u7_U68 (.A1( u2_u4_X_47 ) , .ZN( u2_u4_u7_n156 ) , .A2( u2_u4_u7_n163 ) );
  NAND2_X1 u2_u4_u7_U69 (.A2( u2_u4_X_46 ) , .A1( u2_u4_X_47 ) , .ZN( u2_u4_u7_n125 ) );
  OAI222_X1 u2_u4_u7_U7 (.C2( u2_u4_u7_n101 ) , .B2( u2_u4_u7_n111 ) , .A1( u2_u4_u7_n113 ) , .C1( u2_u4_u7_n146 ) , .A2( u2_u4_u7_n162 ) , .B1( u2_u4_u7_n164 ) , .ZN( u2_u4_u7_n94 ) );
  AND2_X1 u2_u4_u7_U70 (.A2( u2_u4_X_43 ) , .A1( u2_u4_X_44 ) , .ZN( u2_u4_u7_n96 ) );
  AND2_X1 u2_u4_u7_U71 (.A2( u2_u4_X_45 ) , .A1( u2_u4_X_48 ) , .ZN( u2_u4_u7_n102 ) );
  AND2_X1 u2_u4_u7_U72 (.A1( u2_u4_X_48 ) , .A2( u2_u4_u7_n166 ) , .ZN( u2_u4_u7_n93 ) );
  INV_X1 u2_u4_u7_U73 (.A( u2_u4_X_46 ) , .ZN( u2_u4_u7_n163 ) );
  AND2_X1 u2_u4_u7_U74 (.A1( u2_u4_X_44 ) , .ZN( u2_u4_u7_n100 ) , .A2( u2_u4_u7_n167 ) );
  INV_X1 u2_u4_u7_U75 (.A( u2_u4_X_45 ) , .ZN( u2_u4_u7_n166 ) );
  INV_X1 u2_u4_u7_U76 (.A( u2_u4_X_43 ) , .ZN( u2_u4_u7_n167 ) );
  NAND4_X1 u2_u4_u7_U77 (.ZN( u2_out4_5 ) , .A4( u2_u4_u7_n108 ) , .A3( u2_u4_u7_n109 ) , .A1( u2_u4_u7_n116 ) , .A2( u2_u4_u7_n123 ) );
  AOI22_X1 u2_u4_u7_U78 (.ZN( u2_u4_u7_n109 ) , .A2( u2_u4_u7_n126 ) , .B2( u2_u4_u7_n145 ) , .B1( u2_u4_u7_n156 ) , .A1( u2_u4_u7_n171 ) );
  NOR4_X1 u2_u4_u7_U79 (.A4( u2_u4_u7_n104 ) , .A3( u2_u4_u7_n105 ) , .A2( u2_u4_u7_n106 ) , .A1( u2_u4_u7_n107 ) , .ZN( u2_u4_u7_n108 ) );
  INV_X1 u2_u4_u7_U8 (.A( u2_u4_u7_n133 ) , .ZN( u2_u4_u7_n176 ) );
  NAND4_X1 u2_u4_u7_U80 (.ZN( u2_out4_27 ) , .A4( u2_u4_u7_n118 ) , .A3( u2_u4_u7_n119 ) , .A2( u2_u4_u7_n120 ) , .A1( u2_u4_u7_n121 ) );
  OAI21_X1 u2_u4_u7_U81 (.ZN( u2_u4_u7_n121 ) , .B2( u2_u4_u7_n145 ) , .A( u2_u4_u7_n150 ) , .B1( u2_u4_u7_n174 ) );
  OAI21_X1 u2_u4_u7_U82 (.ZN( u2_u4_u7_n120 ) , .A( u2_u4_u7_n161 ) , .B2( u2_u4_u7_n170 ) , .B1( u2_u4_u7_n179 ) );
  NAND4_X1 u2_u4_u7_U83 (.ZN( u2_out4_21 ) , .A4( u2_u4_u7_n157 ) , .A3( u2_u4_u7_n158 ) , .A2( u2_u4_u7_n159 ) , .A1( u2_u4_u7_n160 ) );
  OAI21_X1 u2_u4_u7_U84 (.B1( u2_u4_u7_n145 ) , .ZN( u2_u4_u7_n160 ) , .A( u2_u4_u7_n161 ) , .B2( u2_u4_u7_n177 ) );
  OAI21_X1 u2_u4_u7_U85 (.ZN( u2_u4_u7_n159 ) , .A( u2_u4_u7_n165 ) , .B2( u2_u4_u7_n171 ) , .B1( u2_u4_u7_n174 ) );
  NAND4_X1 u2_u4_u7_U86 (.ZN( u2_out4_15 ) , .A4( u2_u4_u7_n142 ) , .A3( u2_u4_u7_n143 ) , .A2( u2_u4_u7_n144 ) , .A1( u2_u4_u7_n178 ) );
  OR2_X1 u2_u4_u7_U87 (.A2( u2_u4_u7_n125 ) , .A1( u2_u4_u7_n129 ) , .ZN( u2_u4_u7_n144 ) );
  AOI22_X1 u2_u4_u7_U88 (.A2( u2_u4_u7_n126 ) , .ZN( u2_u4_u7_n143 ) , .B2( u2_u4_u7_n165 ) , .B1( u2_u4_u7_n173 ) , .A1( u2_u4_u7_n174 ) );
  NAND2_X1 u2_u4_u7_U89 (.A1( u2_u4_u7_n100 ) , .ZN( u2_u4_u7_n148 ) , .A2( u2_u4_u7_n95 ) );
  OAI221_X1 u2_u4_u7_U9 (.C1( u2_u4_u7_n101 ) , .C2( u2_u4_u7_n147 ) , .ZN( u2_u4_u7_n155 ) , .B2( u2_u4_u7_n162 ) , .A( u2_u4_u7_n91 ) , .B1( u2_u4_u7_n92 ) );
  NAND2_X1 u2_u4_u7_U90 (.A1( u2_u4_u7_n100 ) , .ZN( u2_u4_u7_n113 ) , .A2( u2_u4_u7_n93 ) );
  NAND2_X1 u2_u4_u7_U91 (.A1( u2_u4_u7_n100 ) , .ZN( u2_u4_u7_n138 ) , .A2( u2_u4_u7_n99 ) );
  NAND2_X1 u2_u4_u7_U92 (.A1( u2_u4_u7_n100 ) , .A2( u2_u4_u7_n102 ) , .ZN( u2_u4_u7_n129 ) );
  OAI211_X1 u2_u4_u7_U93 (.B( u2_u4_u7_n122 ) , .A( u2_u4_u7_n123 ) , .C2( u2_u4_u7_n124 ) , .ZN( u2_u4_u7_n154 ) , .C1( u2_u4_u7_n162 ) );
  AOI222_X1 u2_u4_u7_U94 (.ZN( u2_u4_u7_n122 ) , .C2( u2_u4_u7_n126 ) , .C1( u2_u4_u7_n145 ) , .B1( u2_u4_u7_n161 ) , .A2( u2_u4_u7_n165 ) , .B2( u2_u4_u7_n170 ) , .A1( u2_u4_u7_n176 ) );
  NAND3_X1 u2_u4_u7_U95 (.A3( u2_u4_u7_n146 ) , .A2( u2_u4_u7_n147 ) , .A1( u2_u4_u7_n148 ) , .ZN( u2_u4_u7_n151 ) );
  NAND3_X1 u2_u4_u7_U96 (.A3( u2_u4_u7_n131 ) , .A2( u2_u4_u7_n132 ) , .A1( u2_u4_u7_n133 ) , .ZN( u2_u4_u7_n135 ) );
  XOR2_X1 u2_u5_U1 (.B( u2_K6_9 ) , .A( u2_R4_6 ) , .Z( u2_u5_X_9 ) );
  XOR2_X1 u2_u5_U11 (.B( u2_K6_44 ) , .A( u2_R4_29 ) , .Z( u2_u5_X_44 ) );
  XOR2_X1 u2_u5_U12 (.B( u2_K6_43 ) , .A( u2_R4_28 ) , .Z( u2_u5_X_43 ) );
  XOR2_X1 u2_u5_U13 (.B( u2_K6_42 ) , .A( u2_R4_29 ) , .Z( u2_u5_X_42 ) );
  XOR2_X1 u2_u5_U14 (.B( u2_K6_41 ) , .A( u2_R4_28 ) , .Z( u2_u5_X_41 ) );
  XOR2_X1 u2_u5_U19 (.B( u2_K6_37 ) , .A( u2_R4_24 ) , .Z( u2_u5_X_37 ) );
  XOR2_X1 u2_u5_U2 (.B( u2_K6_8 ) , .A( u2_R4_5 ) , .Z( u2_u5_X_8 ) );
  XOR2_X1 u2_u5_U21 (.B( u2_K6_35 ) , .A( u2_R4_24 ) , .Z( u2_u5_X_35 ) );
  XOR2_X1 u2_u5_U23 (.B( u2_K6_33 ) , .A( u2_R4_22 ) , .Z( u2_u5_X_33 ) );
  XOR2_X1 u2_u5_U24 (.B( u2_K6_32 ) , .A( u2_R4_21 ) , .Z( u2_u5_X_32 ) );
  XOR2_X1 u2_u5_U26 (.B( u2_K6_30 ) , .A( u2_R4_21 ) , .Z( u2_u5_X_30 ) );
  XOR2_X1 u2_u5_U27 (.B( u2_K6_2 ) , .A( u2_R4_1 ) , .Z( u2_u5_X_2 ) );
  XOR2_X1 u2_u5_U3 (.B( u2_K6_7 ) , .A( u2_R4_4 ) , .Z( u2_u5_X_7 ) );
  XOR2_X1 u2_u5_U31 (.B( u2_K6_26 ) , .A( u2_R4_17 ) , .Z( u2_u5_X_26 ) );
  XOR2_X1 u2_u5_U33 (.B( u2_K6_24 ) , .A( u2_R4_17 ) , .Z( u2_u5_X_24 ) );
  XOR2_X1 u2_u5_U36 (.B( u2_K6_21 ) , .A( u2_R4_14 ) , .Z( u2_u5_X_21 ) );
  XOR2_X1 u2_u5_U37 (.B( u2_K6_20 ) , .A( u2_R4_13 ) , .Z( u2_u5_X_20 ) );
  XOR2_X1 u2_u5_U38 (.B( u2_K6_1 ) , .A( u2_R4_32 ) , .Z( u2_u5_X_1 ) );
  XOR2_X1 u2_u5_U39 (.B( u2_K6_19 ) , .A( u2_R4_12 ) , .Z( u2_u5_X_19 ) );
  XOR2_X1 u2_u5_U4 (.B( u2_K6_6 ) , .A( u2_R4_5 ) , .Z( u2_u5_X_6 ) );
  XOR2_X1 u2_u5_U40 (.B( u2_K6_18 ) , .A( u2_R4_13 ) , .Z( u2_u5_X_18 ) );
  XOR2_X1 u2_u5_U41 (.B( u2_K6_17 ) , .A( u2_R4_12 ) , .Z( u2_u5_X_17 ) );
  XOR2_X1 u2_u5_U44 (.B( u2_K6_14 ) , .A( u2_R4_9 ) , .Z( u2_u5_X_14 ) );
  XOR2_X1 u2_u5_U45 (.B( u2_K6_13 ) , .A( u2_R4_8 ) , .Z( u2_u5_X_13 ) );
  XOR2_X1 u2_u5_U46 (.B( u2_K6_12 ) , .A( u2_R4_9 ) , .Z( u2_u5_X_12 ) );
  XOR2_X1 u2_u5_U47 (.B( u2_K6_11 ) , .A( u2_R4_8 ) , .Z( u2_u5_X_11 ) );
  XOR2_X1 u2_u5_U5 (.B( u2_K6_5 ) , .A( u2_R4_4 ) , .Z( u2_u5_X_5 ) );
  XOR2_X1 u2_u5_U7 (.B( u2_K6_48 ) , .A( u2_R4_1 ) , .Z( u2_u5_X_48 ) );
  XOR2_X1 u2_u5_U8 (.B( u2_K6_47 ) , .A( u2_R4_32 ) , .Z( u2_u5_X_47 ) );
  XOR2_X1 u2_u5_U9 (.B( u2_K6_46 ) , .A( u2_R4_31 ) , .Z( u2_u5_X_46 ) );
  AND3_X1 u2_u5_u0_U10 (.A2( u2_u5_u0_n112 ) , .ZN( u2_u5_u0_n127 ) , .A3( u2_u5_u0_n130 ) , .A1( u2_u5_u0_n148 ) );
  NAND2_X1 u2_u5_u0_U11 (.ZN( u2_u5_u0_n113 ) , .A1( u2_u5_u0_n139 ) , .A2( u2_u5_u0_n149 ) );
  AND2_X1 u2_u5_u0_U12 (.ZN( u2_u5_u0_n107 ) , .A1( u2_u5_u0_n130 ) , .A2( u2_u5_u0_n140 ) );
  AND2_X1 u2_u5_u0_U13 (.A2( u2_u5_u0_n129 ) , .A1( u2_u5_u0_n130 ) , .ZN( u2_u5_u0_n151 ) );
  AND2_X1 u2_u5_u0_U14 (.A1( u2_u5_u0_n108 ) , .A2( u2_u5_u0_n125 ) , .ZN( u2_u5_u0_n145 ) );
  INV_X1 u2_u5_u0_U15 (.A( u2_u5_u0_n143 ) , .ZN( u2_u5_u0_n173 ) );
  NOR2_X1 u2_u5_u0_U16 (.A2( u2_u5_u0_n136 ) , .ZN( u2_u5_u0_n147 ) , .A1( u2_u5_u0_n160 ) );
  AOI21_X1 u2_u5_u0_U17 (.B1( u2_u5_u0_n103 ) , .ZN( u2_u5_u0_n132 ) , .A( u2_u5_u0_n165 ) , .B2( u2_u5_u0_n93 ) );
  INV_X1 u2_u5_u0_U18 (.A( u2_u5_u0_n142 ) , .ZN( u2_u5_u0_n165 ) );
  OAI22_X1 u2_u5_u0_U19 (.B1( u2_u5_u0_n125 ) , .ZN( u2_u5_u0_n126 ) , .A1( u2_u5_u0_n138 ) , .A2( u2_u5_u0_n146 ) , .B2( u2_u5_u0_n147 ) );
  OAI22_X1 u2_u5_u0_U20 (.B1( u2_u5_u0_n131 ) , .A1( u2_u5_u0_n144 ) , .B2( u2_u5_u0_n147 ) , .A2( u2_u5_u0_n90 ) , .ZN( u2_u5_u0_n91 ) );
  AND3_X1 u2_u5_u0_U21 (.A3( u2_u5_u0_n121 ) , .A2( u2_u5_u0_n125 ) , .A1( u2_u5_u0_n148 ) , .ZN( u2_u5_u0_n90 ) );
  INV_X1 u2_u5_u0_U22 (.A( u2_u5_u0_n136 ) , .ZN( u2_u5_u0_n161 ) );
  AOI22_X1 u2_u5_u0_U23 (.B2( u2_u5_u0_n109 ) , .A2( u2_u5_u0_n110 ) , .ZN( u2_u5_u0_n111 ) , .B1( u2_u5_u0_n118 ) , .A1( u2_u5_u0_n160 ) );
  INV_X1 u2_u5_u0_U24 (.A( u2_u5_u0_n118 ) , .ZN( u2_u5_u0_n158 ) );
  AOI21_X1 u2_u5_u0_U25 (.ZN( u2_u5_u0_n104 ) , .B1( u2_u5_u0_n107 ) , .B2( u2_u5_u0_n141 ) , .A( u2_u5_u0_n144 ) );
  AOI21_X1 u2_u5_u0_U26 (.B1( u2_u5_u0_n127 ) , .B2( u2_u5_u0_n129 ) , .A( u2_u5_u0_n138 ) , .ZN( u2_u5_u0_n96 ) );
  AOI21_X1 u2_u5_u0_U27 (.ZN( u2_u5_u0_n116 ) , .B2( u2_u5_u0_n142 ) , .A( u2_u5_u0_n144 ) , .B1( u2_u5_u0_n166 ) );
  NOR2_X1 u2_u5_u0_U28 (.A1( u2_u5_u0_n120 ) , .ZN( u2_u5_u0_n143 ) , .A2( u2_u5_u0_n167 ) );
  OAI221_X1 u2_u5_u0_U29 (.C1( u2_u5_u0_n112 ) , .ZN( u2_u5_u0_n120 ) , .B1( u2_u5_u0_n138 ) , .B2( u2_u5_u0_n141 ) , .C2( u2_u5_u0_n147 ) , .A( u2_u5_u0_n172 ) );
  INV_X1 u2_u5_u0_U3 (.A( u2_u5_u0_n113 ) , .ZN( u2_u5_u0_n166 ) );
  AOI211_X1 u2_u5_u0_U30 (.B( u2_u5_u0_n115 ) , .A( u2_u5_u0_n116 ) , .C2( u2_u5_u0_n117 ) , .C1( u2_u5_u0_n118 ) , .ZN( u2_u5_u0_n119 ) );
  NAND2_X1 u2_u5_u0_U31 (.A1( u2_u5_u0_n100 ) , .A2( u2_u5_u0_n103 ) , .ZN( u2_u5_u0_n125 ) );
  NAND2_X1 u2_u5_u0_U32 (.A2( u2_u5_u0_n103 ) , .ZN( u2_u5_u0_n140 ) , .A1( u2_u5_u0_n94 ) );
  NAND2_X1 u2_u5_u0_U33 (.A1( u2_u5_u0_n101 ) , .A2( u2_u5_u0_n102 ) , .ZN( u2_u5_u0_n150 ) );
  INV_X1 u2_u5_u0_U34 (.A( u2_u5_u0_n138 ) , .ZN( u2_u5_u0_n160 ) );
  NAND2_X1 u2_u5_u0_U35 (.A2( u2_u5_u0_n102 ) , .A1( u2_u5_u0_n103 ) , .ZN( u2_u5_u0_n149 ) );
  NAND2_X1 u2_u5_u0_U36 (.A2( u2_u5_u0_n100 ) , .A1( u2_u5_u0_n101 ) , .ZN( u2_u5_u0_n139 ) );
  NAND2_X1 u2_u5_u0_U37 (.A2( u2_u5_u0_n100 ) , .ZN( u2_u5_u0_n131 ) , .A1( u2_u5_u0_n92 ) );
  NAND2_X1 u2_u5_u0_U38 (.ZN( u2_u5_u0_n108 ) , .A1( u2_u5_u0_n92 ) , .A2( u2_u5_u0_n94 ) );
  NAND2_X1 u2_u5_u0_U39 (.A2( u2_u5_u0_n102 ) , .ZN( u2_u5_u0_n114 ) , .A1( u2_u5_u0_n92 ) );
  AOI21_X1 u2_u5_u0_U4 (.B1( u2_u5_u0_n114 ) , .ZN( u2_u5_u0_n115 ) , .B2( u2_u5_u0_n129 ) , .A( u2_u5_u0_n161 ) );
  NAND2_X1 u2_u5_u0_U40 (.A1( u2_u5_u0_n101 ) , .ZN( u2_u5_u0_n130 ) , .A2( u2_u5_u0_n94 ) );
  NAND2_X1 u2_u5_u0_U41 (.A2( u2_u5_u0_n101 ) , .ZN( u2_u5_u0_n121 ) , .A1( u2_u5_u0_n93 ) );
  INV_X1 u2_u5_u0_U42 (.ZN( u2_u5_u0_n172 ) , .A( u2_u5_u0_n88 ) );
  OAI222_X1 u2_u5_u0_U43 (.C1( u2_u5_u0_n108 ) , .A1( u2_u5_u0_n125 ) , .B2( u2_u5_u0_n128 ) , .B1( u2_u5_u0_n144 ) , .A2( u2_u5_u0_n158 ) , .C2( u2_u5_u0_n161 ) , .ZN( u2_u5_u0_n88 ) );
  NAND2_X1 u2_u5_u0_U44 (.ZN( u2_u5_u0_n112 ) , .A2( u2_u5_u0_n92 ) , .A1( u2_u5_u0_n93 ) );
  OR3_X1 u2_u5_u0_U45 (.A3( u2_u5_u0_n152 ) , .A2( u2_u5_u0_n153 ) , .A1( u2_u5_u0_n154 ) , .ZN( u2_u5_u0_n155 ) );
  AOI21_X1 u2_u5_u0_U46 (.A( u2_u5_u0_n144 ) , .B2( u2_u5_u0_n145 ) , .B1( u2_u5_u0_n146 ) , .ZN( u2_u5_u0_n154 ) );
  AOI21_X1 u2_u5_u0_U47 (.B2( u2_u5_u0_n150 ) , .B1( u2_u5_u0_n151 ) , .ZN( u2_u5_u0_n152 ) , .A( u2_u5_u0_n158 ) );
  AOI21_X1 u2_u5_u0_U48 (.A( u2_u5_u0_n147 ) , .B2( u2_u5_u0_n148 ) , .B1( u2_u5_u0_n149 ) , .ZN( u2_u5_u0_n153 ) );
  INV_X1 u2_u5_u0_U49 (.ZN( u2_u5_u0_n171 ) , .A( u2_u5_u0_n99 ) );
  AOI21_X1 u2_u5_u0_U5 (.B2( u2_u5_u0_n131 ) , .ZN( u2_u5_u0_n134 ) , .B1( u2_u5_u0_n151 ) , .A( u2_u5_u0_n158 ) );
  OAI211_X1 u2_u5_u0_U50 (.C2( u2_u5_u0_n140 ) , .C1( u2_u5_u0_n161 ) , .A( u2_u5_u0_n169 ) , .B( u2_u5_u0_n98 ) , .ZN( u2_u5_u0_n99 ) );
  AOI211_X1 u2_u5_u0_U51 (.C1( u2_u5_u0_n118 ) , .A( u2_u5_u0_n123 ) , .B( u2_u5_u0_n96 ) , .C2( u2_u5_u0_n97 ) , .ZN( u2_u5_u0_n98 ) );
  INV_X1 u2_u5_u0_U52 (.ZN( u2_u5_u0_n169 ) , .A( u2_u5_u0_n91 ) );
  NOR2_X1 u2_u5_u0_U53 (.A2( u2_u5_X_2 ) , .ZN( u2_u5_u0_n103 ) , .A1( u2_u5_u0_n164 ) );
  NOR2_X1 u2_u5_u0_U54 (.A2( u2_u5_X_4 ) , .A1( u2_u5_X_5 ) , .ZN( u2_u5_u0_n118 ) );
  NOR2_X1 u2_u5_u0_U55 (.A2( u2_u5_X_1 ) , .A1( u2_u5_X_2 ) , .ZN( u2_u5_u0_n92 ) );
  NOR2_X1 u2_u5_u0_U56 (.A2( u2_u5_X_1 ) , .ZN( u2_u5_u0_n101 ) , .A1( u2_u5_u0_n163 ) );
  NOR2_X1 u2_u5_u0_U57 (.A2( u2_u5_X_3 ) , .A1( u2_u5_X_6 ) , .ZN( u2_u5_u0_n94 ) );
  NOR2_X1 u2_u5_u0_U58 (.A2( u2_u5_X_6 ) , .ZN( u2_u5_u0_n100 ) , .A1( u2_u5_u0_n162 ) );
  NAND2_X1 u2_u5_u0_U59 (.A2( u2_u5_X_4 ) , .A1( u2_u5_X_5 ) , .ZN( u2_u5_u0_n144 ) );
  NOR2_X1 u2_u5_u0_U6 (.A1( u2_u5_u0_n108 ) , .ZN( u2_u5_u0_n123 ) , .A2( u2_u5_u0_n158 ) );
  NOR2_X1 u2_u5_u0_U60 (.A2( u2_u5_X_5 ) , .ZN( u2_u5_u0_n136 ) , .A1( u2_u5_u0_n159 ) );
  NAND2_X1 u2_u5_u0_U61 (.A1( u2_u5_X_5 ) , .ZN( u2_u5_u0_n138 ) , .A2( u2_u5_u0_n159 ) );
  AND2_X1 u2_u5_u0_U62 (.A2( u2_u5_X_3 ) , .A1( u2_u5_X_6 ) , .ZN( u2_u5_u0_n102 ) );
  AND2_X1 u2_u5_u0_U63 (.A1( u2_u5_X_6 ) , .A2( u2_u5_u0_n162 ) , .ZN( u2_u5_u0_n93 ) );
  INV_X1 u2_u5_u0_U64 (.A( u2_u5_X_4 ) , .ZN( u2_u5_u0_n159 ) );
  INV_X1 u2_u5_u0_U65 (.A( u2_u5_X_1 ) , .ZN( u2_u5_u0_n164 ) );
  INV_X1 u2_u5_u0_U66 (.A( u2_u5_X_2 ) , .ZN( u2_u5_u0_n163 ) );
  INV_X1 u2_u5_u0_U67 (.A( u2_u5_X_3 ) , .ZN( u2_u5_u0_n162 ) );
  INV_X1 u2_u5_u0_U68 (.A( u2_u5_u0_n126 ) , .ZN( u2_u5_u0_n168 ) );
  AOI211_X1 u2_u5_u0_U69 (.B( u2_u5_u0_n133 ) , .A( u2_u5_u0_n134 ) , .C2( u2_u5_u0_n135 ) , .C1( u2_u5_u0_n136 ) , .ZN( u2_u5_u0_n137 ) );
  OAI21_X1 u2_u5_u0_U7 (.B1( u2_u5_u0_n150 ) , .B2( u2_u5_u0_n158 ) , .A( u2_u5_u0_n172 ) , .ZN( u2_u5_u0_n89 ) );
  OR4_X1 u2_u5_u0_U70 (.ZN( u2_out5_17 ) , .A4( u2_u5_u0_n122 ) , .A2( u2_u5_u0_n123 ) , .A1( u2_u5_u0_n124 ) , .A3( u2_u5_u0_n170 ) );
  AOI21_X1 u2_u5_u0_U71 (.B2( u2_u5_u0_n107 ) , .ZN( u2_u5_u0_n124 ) , .B1( u2_u5_u0_n128 ) , .A( u2_u5_u0_n161 ) );
  INV_X1 u2_u5_u0_U72 (.A( u2_u5_u0_n111 ) , .ZN( u2_u5_u0_n170 ) );
  OR4_X1 u2_u5_u0_U73 (.ZN( u2_out5_31 ) , .A4( u2_u5_u0_n155 ) , .A2( u2_u5_u0_n156 ) , .A1( u2_u5_u0_n157 ) , .A3( u2_u5_u0_n173 ) );
  AOI21_X1 u2_u5_u0_U74 (.A( u2_u5_u0_n138 ) , .B2( u2_u5_u0_n139 ) , .B1( u2_u5_u0_n140 ) , .ZN( u2_u5_u0_n157 ) );
  AOI21_X1 u2_u5_u0_U75 (.B2( u2_u5_u0_n141 ) , .B1( u2_u5_u0_n142 ) , .ZN( u2_u5_u0_n156 ) , .A( u2_u5_u0_n161 ) );
  INV_X1 u2_u5_u0_U76 (.ZN( u2_u5_u0_n174 ) , .A( u2_u5_u0_n89 ) );
  AOI211_X1 u2_u5_u0_U77 (.B( u2_u5_u0_n104 ) , .A( u2_u5_u0_n105 ) , .ZN( u2_u5_u0_n106 ) , .C2( u2_u5_u0_n113 ) , .C1( u2_u5_u0_n160 ) );
  NOR2_X1 u2_u5_u0_U78 (.A1( u2_u5_u0_n163 ) , .A2( u2_u5_u0_n164 ) , .ZN( u2_u5_u0_n95 ) );
  OAI221_X1 u2_u5_u0_U79 (.C1( u2_u5_u0_n121 ) , .ZN( u2_u5_u0_n122 ) , .B2( u2_u5_u0_n127 ) , .A( u2_u5_u0_n143 ) , .B1( u2_u5_u0_n144 ) , .C2( u2_u5_u0_n147 ) );
  AND2_X1 u2_u5_u0_U8 (.A1( u2_u5_u0_n114 ) , .A2( u2_u5_u0_n121 ) , .ZN( u2_u5_u0_n146 ) );
  AOI21_X1 u2_u5_u0_U80 (.B1( u2_u5_u0_n132 ) , .ZN( u2_u5_u0_n133 ) , .A( u2_u5_u0_n144 ) , .B2( u2_u5_u0_n166 ) );
  OAI22_X1 u2_u5_u0_U81 (.ZN( u2_u5_u0_n105 ) , .A2( u2_u5_u0_n132 ) , .B1( u2_u5_u0_n146 ) , .A1( u2_u5_u0_n147 ) , .B2( u2_u5_u0_n161 ) );
  NAND2_X1 u2_u5_u0_U82 (.ZN( u2_u5_u0_n110 ) , .A2( u2_u5_u0_n132 ) , .A1( u2_u5_u0_n145 ) );
  INV_X1 u2_u5_u0_U83 (.A( u2_u5_u0_n119 ) , .ZN( u2_u5_u0_n167 ) );
  NAND2_X1 u2_u5_u0_U84 (.ZN( u2_u5_u0_n148 ) , .A1( u2_u5_u0_n93 ) , .A2( u2_u5_u0_n95 ) );
  NAND2_X1 u2_u5_u0_U85 (.A1( u2_u5_u0_n100 ) , .ZN( u2_u5_u0_n129 ) , .A2( u2_u5_u0_n95 ) );
  NAND2_X1 u2_u5_u0_U86 (.A1( u2_u5_u0_n102 ) , .ZN( u2_u5_u0_n128 ) , .A2( u2_u5_u0_n95 ) );
  NAND2_X1 u2_u5_u0_U87 (.ZN( u2_u5_u0_n142 ) , .A1( u2_u5_u0_n94 ) , .A2( u2_u5_u0_n95 ) );
  NAND3_X1 u2_u5_u0_U88 (.ZN( u2_out5_23 ) , .A3( u2_u5_u0_n137 ) , .A1( u2_u5_u0_n168 ) , .A2( u2_u5_u0_n171 ) );
  NAND3_X1 u2_u5_u0_U89 (.A3( u2_u5_u0_n127 ) , .A2( u2_u5_u0_n128 ) , .ZN( u2_u5_u0_n135 ) , .A1( u2_u5_u0_n150 ) );
  AND2_X1 u2_u5_u0_U9 (.A1( u2_u5_u0_n131 ) , .ZN( u2_u5_u0_n141 ) , .A2( u2_u5_u0_n150 ) );
  NAND3_X1 u2_u5_u0_U90 (.ZN( u2_u5_u0_n117 ) , .A3( u2_u5_u0_n132 ) , .A2( u2_u5_u0_n139 ) , .A1( u2_u5_u0_n148 ) );
  NAND3_X1 u2_u5_u0_U91 (.ZN( u2_u5_u0_n109 ) , .A2( u2_u5_u0_n114 ) , .A3( u2_u5_u0_n140 ) , .A1( u2_u5_u0_n149 ) );
  NAND3_X1 u2_u5_u0_U92 (.ZN( u2_out5_9 ) , .A3( u2_u5_u0_n106 ) , .A2( u2_u5_u0_n171 ) , .A1( u2_u5_u0_n174 ) );
  NAND3_X1 u2_u5_u0_U93 (.A2( u2_u5_u0_n128 ) , .A1( u2_u5_u0_n132 ) , .A3( u2_u5_u0_n146 ) , .ZN( u2_u5_u0_n97 ) );
  NOR2_X1 u2_u5_u1_U10 (.A1( u2_u5_u1_n112 ) , .A2( u2_u5_u1_n116 ) , .ZN( u2_u5_u1_n118 ) );
  NAND3_X1 u2_u5_u1_U100 (.ZN( u2_u5_u1_n113 ) , .A1( u2_u5_u1_n120 ) , .A3( u2_u5_u1_n133 ) , .A2( u2_u5_u1_n155 ) );
  OAI21_X1 u2_u5_u1_U11 (.ZN( u2_u5_u1_n101 ) , .B1( u2_u5_u1_n141 ) , .A( u2_u5_u1_n146 ) , .B2( u2_u5_u1_n183 ) );
  AOI21_X1 u2_u5_u1_U12 (.B2( u2_u5_u1_n155 ) , .B1( u2_u5_u1_n156 ) , .ZN( u2_u5_u1_n157 ) , .A( u2_u5_u1_n174 ) );
  NAND2_X1 u2_u5_u1_U13 (.ZN( u2_u5_u1_n140 ) , .A2( u2_u5_u1_n150 ) , .A1( u2_u5_u1_n155 ) );
  NAND2_X1 u2_u5_u1_U14 (.A1( u2_u5_u1_n131 ) , .ZN( u2_u5_u1_n147 ) , .A2( u2_u5_u1_n153 ) );
  INV_X1 u2_u5_u1_U15 (.A( u2_u5_u1_n139 ) , .ZN( u2_u5_u1_n174 ) );
  OR4_X1 u2_u5_u1_U16 (.A4( u2_u5_u1_n106 ) , .A3( u2_u5_u1_n107 ) , .ZN( u2_u5_u1_n108 ) , .A1( u2_u5_u1_n117 ) , .A2( u2_u5_u1_n184 ) );
  AOI21_X1 u2_u5_u1_U17 (.ZN( u2_u5_u1_n106 ) , .A( u2_u5_u1_n112 ) , .B1( u2_u5_u1_n154 ) , .B2( u2_u5_u1_n156 ) );
  INV_X1 u2_u5_u1_U18 (.A( u2_u5_u1_n101 ) , .ZN( u2_u5_u1_n184 ) );
  AOI21_X1 u2_u5_u1_U19 (.ZN( u2_u5_u1_n107 ) , .B1( u2_u5_u1_n134 ) , .B2( u2_u5_u1_n149 ) , .A( u2_u5_u1_n174 ) );
  INV_X1 u2_u5_u1_U20 (.A( u2_u5_u1_n112 ) , .ZN( u2_u5_u1_n171 ) );
  NAND2_X1 u2_u5_u1_U21 (.ZN( u2_u5_u1_n141 ) , .A1( u2_u5_u1_n153 ) , .A2( u2_u5_u1_n156 ) );
  AND2_X1 u2_u5_u1_U22 (.A1( u2_u5_u1_n123 ) , .ZN( u2_u5_u1_n134 ) , .A2( u2_u5_u1_n161 ) );
  NAND2_X1 u2_u5_u1_U23 (.A2( u2_u5_u1_n115 ) , .A1( u2_u5_u1_n116 ) , .ZN( u2_u5_u1_n148 ) );
  NAND2_X1 u2_u5_u1_U24 (.A2( u2_u5_u1_n133 ) , .A1( u2_u5_u1_n135 ) , .ZN( u2_u5_u1_n159 ) );
  NAND2_X1 u2_u5_u1_U25 (.A2( u2_u5_u1_n115 ) , .A1( u2_u5_u1_n120 ) , .ZN( u2_u5_u1_n132 ) );
  INV_X1 u2_u5_u1_U26 (.A( u2_u5_u1_n154 ) , .ZN( u2_u5_u1_n178 ) );
  INV_X1 u2_u5_u1_U27 (.A( u2_u5_u1_n151 ) , .ZN( u2_u5_u1_n183 ) );
  AND2_X1 u2_u5_u1_U28 (.A1( u2_u5_u1_n129 ) , .A2( u2_u5_u1_n133 ) , .ZN( u2_u5_u1_n149 ) );
  INV_X1 u2_u5_u1_U29 (.A( u2_u5_u1_n131 ) , .ZN( u2_u5_u1_n180 ) );
  INV_X1 u2_u5_u1_U3 (.A( u2_u5_u1_n159 ) , .ZN( u2_u5_u1_n182 ) );
  OAI221_X1 u2_u5_u1_U30 (.A( u2_u5_u1_n119 ) , .C2( u2_u5_u1_n129 ) , .ZN( u2_u5_u1_n138 ) , .B2( u2_u5_u1_n152 ) , .C1( u2_u5_u1_n174 ) , .B1( u2_u5_u1_n187 ) );
  INV_X1 u2_u5_u1_U31 (.A( u2_u5_u1_n148 ) , .ZN( u2_u5_u1_n187 ) );
  AOI211_X1 u2_u5_u1_U32 (.B( u2_u5_u1_n117 ) , .A( u2_u5_u1_n118 ) , .ZN( u2_u5_u1_n119 ) , .C2( u2_u5_u1_n146 ) , .C1( u2_u5_u1_n159 ) );
  NOR2_X1 u2_u5_u1_U33 (.A1( u2_u5_u1_n168 ) , .A2( u2_u5_u1_n176 ) , .ZN( u2_u5_u1_n98 ) );
  OAI21_X1 u2_u5_u1_U34 (.B2( u2_u5_u1_n123 ) , .ZN( u2_u5_u1_n145 ) , .B1( u2_u5_u1_n160 ) , .A( u2_u5_u1_n185 ) );
  INV_X1 u2_u5_u1_U35 (.A( u2_u5_u1_n122 ) , .ZN( u2_u5_u1_n185 ) );
  AOI21_X1 u2_u5_u1_U36 (.B2( u2_u5_u1_n120 ) , .B1( u2_u5_u1_n121 ) , .ZN( u2_u5_u1_n122 ) , .A( u2_u5_u1_n128 ) );
  NAND2_X1 u2_u5_u1_U37 (.A1( u2_u5_u1_n128 ) , .ZN( u2_u5_u1_n146 ) , .A2( u2_u5_u1_n160 ) );
  NAND2_X1 u2_u5_u1_U38 (.A2( u2_u5_u1_n112 ) , .ZN( u2_u5_u1_n139 ) , .A1( u2_u5_u1_n152 ) );
  NAND2_X1 u2_u5_u1_U39 (.A1( u2_u5_u1_n105 ) , .ZN( u2_u5_u1_n156 ) , .A2( u2_u5_u1_n99 ) );
  AOI221_X1 u2_u5_u1_U4 (.A( u2_u5_u1_n138 ) , .C2( u2_u5_u1_n139 ) , .C1( u2_u5_u1_n140 ) , .B2( u2_u5_u1_n141 ) , .ZN( u2_u5_u1_n142 ) , .B1( u2_u5_u1_n175 ) );
  AOI221_X1 u2_u5_u1_U40 (.B1( u2_u5_u1_n140 ) , .ZN( u2_u5_u1_n167 ) , .B2( u2_u5_u1_n172 ) , .C2( u2_u5_u1_n175 ) , .C1( u2_u5_u1_n178 ) , .A( u2_u5_u1_n188 ) );
  INV_X1 u2_u5_u1_U41 (.ZN( u2_u5_u1_n188 ) , .A( u2_u5_u1_n97 ) );
  AOI211_X1 u2_u5_u1_U42 (.A( u2_u5_u1_n118 ) , .C1( u2_u5_u1_n132 ) , .C2( u2_u5_u1_n139 ) , .B( u2_u5_u1_n96 ) , .ZN( u2_u5_u1_n97 ) );
  AOI21_X1 u2_u5_u1_U43 (.B2( u2_u5_u1_n121 ) , .B1( u2_u5_u1_n135 ) , .A( u2_u5_u1_n152 ) , .ZN( u2_u5_u1_n96 ) );
  NOR2_X1 u2_u5_u1_U44 (.ZN( u2_u5_u1_n117 ) , .A1( u2_u5_u1_n121 ) , .A2( u2_u5_u1_n160 ) );
  AOI21_X1 u2_u5_u1_U45 (.A( u2_u5_u1_n128 ) , .B2( u2_u5_u1_n129 ) , .ZN( u2_u5_u1_n130 ) , .B1( u2_u5_u1_n150 ) );
  NAND2_X1 u2_u5_u1_U46 (.ZN( u2_u5_u1_n112 ) , .A1( u2_u5_u1_n169 ) , .A2( u2_u5_u1_n170 ) );
  NAND2_X1 u2_u5_u1_U47 (.ZN( u2_u5_u1_n129 ) , .A2( u2_u5_u1_n95 ) , .A1( u2_u5_u1_n98 ) );
  NAND2_X1 u2_u5_u1_U48 (.A1( u2_u5_u1_n102 ) , .ZN( u2_u5_u1_n154 ) , .A2( u2_u5_u1_n99 ) );
  NAND2_X1 u2_u5_u1_U49 (.A2( u2_u5_u1_n100 ) , .ZN( u2_u5_u1_n135 ) , .A1( u2_u5_u1_n99 ) );
  AOI211_X1 u2_u5_u1_U5 (.ZN( u2_u5_u1_n124 ) , .A( u2_u5_u1_n138 ) , .C2( u2_u5_u1_n139 ) , .B( u2_u5_u1_n145 ) , .C1( u2_u5_u1_n147 ) );
  AOI21_X1 u2_u5_u1_U50 (.A( u2_u5_u1_n152 ) , .B2( u2_u5_u1_n153 ) , .B1( u2_u5_u1_n154 ) , .ZN( u2_u5_u1_n158 ) );
  INV_X1 u2_u5_u1_U51 (.A( u2_u5_u1_n160 ) , .ZN( u2_u5_u1_n175 ) );
  NAND2_X1 u2_u5_u1_U52 (.A1( u2_u5_u1_n100 ) , .ZN( u2_u5_u1_n116 ) , .A2( u2_u5_u1_n95 ) );
  NAND2_X1 u2_u5_u1_U53 (.A1( u2_u5_u1_n102 ) , .ZN( u2_u5_u1_n131 ) , .A2( u2_u5_u1_n95 ) );
  NAND2_X1 u2_u5_u1_U54 (.A2( u2_u5_u1_n104 ) , .ZN( u2_u5_u1_n121 ) , .A1( u2_u5_u1_n98 ) );
  NAND2_X1 u2_u5_u1_U55 (.A1( u2_u5_u1_n103 ) , .ZN( u2_u5_u1_n153 ) , .A2( u2_u5_u1_n98 ) );
  NAND2_X1 u2_u5_u1_U56 (.A2( u2_u5_u1_n104 ) , .A1( u2_u5_u1_n105 ) , .ZN( u2_u5_u1_n133 ) );
  NAND2_X1 u2_u5_u1_U57 (.ZN( u2_u5_u1_n150 ) , .A2( u2_u5_u1_n98 ) , .A1( u2_u5_u1_n99 ) );
  NAND2_X1 u2_u5_u1_U58 (.A1( u2_u5_u1_n105 ) , .ZN( u2_u5_u1_n155 ) , .A2( u2_u5_u1_n95 ) );
  OAI21_X1 u2_u5_u1_U59 (.ZN( u2_u5_u1_n109 ) , .B1( u2_u5_u1_n129 ) , .B2( u2_u5_u1_n160 ) , .A( u2_u5_u1_n167 ) );
  AOI22_X1 u2_u5_u1_U6 (.B2( u2_u5_u1_n136 ) , .A2( u2_u5_u1_n137 ) , .ZN( u2_u5_u1_n143 ) , .A1( u2_u5_u1_n171 ) , .B1( u2_u5_u1_n173 ) );
  NAND2_X1 u2_u5_u1_U60 (.A2( u2_u5_u1_n100 ) , .A1( u2_u5_u1_n103 ) , .ZN( u2_u5_u1_n120 ) );
  NAND2_X1 u2_u5_u1_U61 (.A1( u2_u5_u1_n102 ) , .A2( u2_u5_u1_n104 ) , .ZN( u2_u5_u1_n115 ) );
  NAND2_X1 u2_u5_u1_U62 (.A2( u2_u5_u1_n100 ) , .A1( u2_u5_u1_n104 ) , .ZN( u2_u5_u1_n151 ) );
  NAND2_X1 u2_u5_u1_U63 (.A2( u2_u5_u1_n103 ) , .A1( u2_u5_u1_n105 ) , .ZN( u2_u5_u1_n161 ) );
  INV_X1 u2_u5_u1_U64 (.A( u2_u5_u1_n152 ) , .ZN( u2_u5_u1_n173 ) );
  INV_X1 u2_u5_u1_U65 (.A( u2_u5_u1_n128 ) , .ZN( u2_u5_u1_n172 ) );
  NAND2_X1 u2_u5_u1_U66 (.A2( u2_u5_u1_n102 ) , .A1( u2_u5_u1_n103 ) , .ZN( u2_u5_u1_n123 ) );
  AOI211_X1 u2_u5_u1_U67 (.B( u2_u5_u1_n162 ) , .A( u2_u5_u1_n163 ) , .C2( u2_u5_u1_n164 ) , .ZN( u2_u5_u1_n165 ) , .C1( u2_u5_u1_n171 ) );
  AOI21_X1 u2_u5_u1_U68 (.A( u2_u5_u1_n160 ) , .B2( u2_u5_u1_n161 ) , .ZN( u2_u5_u1_n162 ) , .B1( u2_u5_u1_n182 ) );
  OR2_X1 u2_u5_u1_U69 (.A2( u2_u5_u1_n157 ) , .A1( u2_u5_u1_n158 ) , .ZN( u2_u5_u1_n163 ) );
  INV_X1 u2_u5_u1_U7 (.A( u2_u5_u1_n147 ) , .ZN( u2_u5_u1_n181 ) );
  NOR2_X1 u2_u5_u1_U70 (.A2( u2_u5_X_7 ) , .A1( u2_u5_X_8 ) , .ZN( u2_u5_u1_n95 ) );
  NOR2_X1 u2_u5_u1_U71 (.A1( u2_u5_X_12 ) , .A2( u2_u5_X_9 ) , .ZN( u2_u5_u1_n100 ) );
  NOR2_X1 u2_u5_u1_U72 (.A2( u2_u5_X_8 ) , .A1( u2_u5_u1_n177 ) , .ZN( u2_u5_u1_n99 ) );
  NOR2_X1 u2_u5_u1_U73 (.A2( u2_u5_X_12 ) , .ZN( u2_u5_u1_n102 ) , .A1( u2_u5_u1_n176 ) );
  NOR2_X1 u2_u5_u1_U74 (.A2( u2_u5_X_9 ) , .ZN( u2_u5_u1_n105 ) , .A1( u2_u5_u1_n168 ) );
  NAND2_X1 u2_u5_u1_U75 (.A1( u2_u5_X_10 ) , .ZN( u2_u5_u1_n160 ) , .A2( u2_u5_u1_n169 ) );
  NAND2_X1 u2_u5_u1_U76 (.A2( u2_u5_X_10 ) , .A1( u2_u5_X_11 ) , .ZN( u2_u5_u1_n152 ) );
  NAND2_X1 u2_u5_u1_U77 (.A1( u2_u5_X_11 ) , .ZN( u2_u5_u1_n128 ) , .A2( u2_u5_u1_n170 ) );
  AND2_X1 u2_u5_u1_U78 (.A2( u2_u5_X_7 ) , .A1( u2_u5_X_8 ) , .ZN( u2_u5_u1_n104 ) );
  AND2_X1 u2_u5_u1_U79 (.A1( u2_u5_X_8 ) , .ZN( u2_u5_u1_n103 ) , .A2( u2_u5_u1_n177 ) );
  AOI22_X1 u2_u5_u1_U8 (.B2( u2_u5_u1_n113 ) , .A2( u2_u5_u1_n114 ) , .ZN( u2_u5_u1_n125 ) , .A1( u2_u5_u1_n171 ) , .B1( u2_u5_u1_n173 ) );
  INV_X1 u2_u5_u1_U80 (.A( u2_u5_X_10 ) , .ZN( u2_u5_u1_n170 ) );
  INV_X1 u2_u5_u1_U81 (.A( u2_u5_X_9 ) , .ZN( u2_u5_u1_n176 ) );
  INV_X1 u2_u5_u1_U82 (.A( u2_u5_X_11 ) , .ZN( u2_u5_u1_n169 ) );
  INV_X1 u2_u5_u1_U83 (.A( u2_u5_X_12 ) , .ZN( u2_u5_u1_n168 ) );
  INV_X1 u2_u5_u1_U84 (.A( u2_u5_X_7 ) , .ZN( u2_u5_u1_n177 ) );
  NAND4_X1 u2_u5_u1_U85 (.ZN( u2_out5_28 ) , .A4( u2_u5_u1_n124 ) , .A3( u2_u5_u1_n125 ) , .A2( u2_u5_u1_n126 ) , .A1( u2_u5_u1_n127 ) );
  OAI21_X1 u2_u5_u1_U86 (.ZN( u2_u5_u1_n127 ) , .B2( u2_u5_u1_n139 ) , .B1( u2_u5_u1_n175 ) , .A( u2_u5_u1_n183 ) );
  OAI21_X1 u2_u5_u1_U87 (.ZN( u2_u5_u1_n126 ) , .B2( u2_u5_u1_n140 ) , .A( u2_u5_u1_n146 ) , .B1( u2_u5_u1_n178 ) );
  NAND4_X1 u2_u5_u1_U88 (.ZN( u2_out5_18 ) , .A4( u2_u5_u1_n165 ) , .A3( u2_u5_u1_n166 ) , .A1( u2_u5_u1_n167 ) , .A2( u2_u5_u1_n186 ) );
  AOI22_X1 u2_u5_u1_U89 (.B2( u2_u5_u1_n146 ) , .B1( u2_u5_u1_n147 ) , .A2( u2_u5_u1_n148 ) , .ZN( u2_u5_u1_n166 ) , .A1( u2_u5_u1_n172 ) );
  NAND2_X1 u2_u5_u1_U9 (.ZN( u2_u5_u1_n114 ) , .A1( u2_u5_u1_n134 ) , .A2( u2_u5_u1_n156 ) );
  INV_X1 u2_u5_u1_U90 (.A( u2_u5_u1_n145 ) , .ZN( u2_u5_u1_n186 ) );
  NAND4_X1 u2_u5_u1_U91 (.ZN( u2_out5_2 ) , .A4( u2_u5_u1_n142 ) , .A3( u2_u5_u1_n143 ) , .A2( u2_u5_u1_n144 ) , .A1( u2_u5_u1_n179 ) );
  OAI21_X1 u2_u5_u1_U92 (.B2( u2_u5_u1_n132 ) , .ZN( u2_u5_u1_n144 ) , .A( u2_u5_u1_n146 ) , .B1( u2_u5_u1_n180 ) );
  INV_X1 u2_u5_u1_U93 (.A( u2_u5_u1_n130 ) , .ZN( u2_u5_u1_n179 ) );
  OR4_X1 u2_u5_u1_U94 (.ZN( u2_out5_13 ) , .A4( u2_u5_u1_n108 ) , .A3( u2_u5_u1_n109 ) , .A2( u2_u5_u1_n110 ) , .A1( u2_u5_u1_n111 ) );
  AOI21_X1 u2_u5_u1_U95 (.ZN( u2_u5_u1_n110 ) , .A( u2_u5_u1_n116 ) , .B1( u2_u5_u1_n152 ) , .B2( u2_u5_u1_n160 ) );
  AOI21_X1 u2_u5_u1_U96 (.ZN( u2_u5_u1_n111 ) , .A( u2_u5_u1_n128 ) , .B2( u2_u5_u1_n131 ) , .B1( u2_u5_u1_n135 ) );
  NAND3_X1 u2_u5_u1_U97 (.A3( u2_u5_u1_n149 ) , .A2( u2_u5_u1_n150 ) , .A1( u2_u5_u1_n151 ) , .ZN( u2_u5_u1_n164 ) );
  NAND3_X1 u2_u5_u1_U98 (.A3( u2_u5_u1_n134 ) , .A2( u2_u5_u1_n135 ) , .ZN( u2_u5_u1_n136 ) , .A1( u2_u5_u1_n151 ) );
  NAND3_X1 u2_u5_u1_U99 (.A1( u2_u5_u1_n133 ) , .ZN( u2_u5_u1_n137 ) , .A2( u2_u5_u1_n154 ) , .A3( u2_u5_u1_n181 ) );
  OAI22_X1 u2_u5_u2_U10 (.ZN( u2_u5_u2_n109 ) , .A2( u2_u5_u2_n113 ) , .B2( u2_u5_u2_n133 ) , .B1( u2_u5_u2_n167 ) , .A1( u2_u5_u2_n168 ) );
  NAND3_X1 u2_u5_u2_U100 (.A2( u2_u5_u2_n100 ) , .A1( u2_u5_u2_n104 ) , .A3( u2_u5_u2_n138 ) , .ZN( u2_u5_u2_n98 ) );
  OAI22_X1 u2_u5_u2_U11 (.B1( u2_u5_u2_n151 ) , .A2( u2_u5_u2_n152 ) , .A1( u2_u5_u2_n153 ) , .ZN( u2_u5_u2_n160 ) , .B2( u2_u5_u2_n168 ) );
  NOR3_X1 u2_u5_u2_U12 (.A1( u2_u5_u2_n150 ) , .ZN( u2_u5_u2_n151 ) , .A3( u2_u5_u2_n175 ) , .A2( u2_u5_u2_n188 ) );
  AOI21_X1 u2_u5_u2_U13 (.ZN( u2_u5_u2_n144 ) , .B2( u2_u5_u2_n155 ) , .A( u2_u5_u2_n172 ) , .B1( u2_u5_u2_n185 ) );
  AOI21_X1 u2_u5_u2_U14 (.B2( u2_u5_u2_n143 ) , .ZN( u2_u5_u2_n145 ) , .B1( u2_u5_u2_n152 ) , .A( u2_u5_u2_n171 ) );
  AOI21_X1 u2_u5_u2_U15 (.B2( u2_u5_u2_n120 ) , .B1( u2_u5_u2_n121 ) , .ZN( u2_u5_u2_n126 ) , .A( u2_u5_u2_n167 ) );
  INV_X1 u2_u5_u2_U16 (.A( u2_u5_u2_n156 ) , .ZN( u2_u5_u2_n171 ) );
  INV_X1 u2_u5_u2_U17 (.A( u2_u5_u2_n120 ) , .ZN( u2_u5_u2_n188 ) );
  NAND2_X1 u2_u5_u2_U18 (.A2( u2_u5_u2_n122 ) , .ZN( u2_u5_u2_n150 ) , .A1( u2_u5_u2_n152 ) );
  INV_X1 u2_u5_u2_U19 (.A( u2_u5_u2_n153 ) , .ZN( u2_u5_u2_n170 ) );
  INV_X1 u2_u5_u2_U20 (.A( u2_u5_u2_n137 ) , .ZN( u2_u5_u2_n173 ) );
  NAND2_X1 u2_u5_u2_U21 (.A1( u2_u5_u2_n132 ) , .A2( u2_u5_u2_n139 ) , .ZN( u2_u5_u2_n157 ) );
  INV_X1 u2_u5_u2_U22 (.A( u2_u5_u2_n113 ) , .ZN( u2_u5_u2_n178 ) );
  INV_X1 u2_u5_u2_U23 (.A( u2_u5_u2_n139 ) , .ZN( u2_u5_u2_n175 ) );
  INV_X1 u2_u5_u2_U24 (.A( u2_u5_u2_n155 ) , .ZN( u2_u5_u2_n181 ) );
  INV_X1 u2_u5_u2_U25 (.A( u2_u5_u2_n119 ) , .ZN( u2_u5_u2_n177 ) );
  INV_X1 u2_u5_u2_U26 (.A( u2_u5_u2_n116 ) , .ZN( u2_u5_u2_n180 ) );
  INV_X1 u2_u5_u2_U27 (.A( u2_u5_u2_n131 ) , .ZN( u2_u5_u2_n179 ) );
  INV_X1 u2_u5_u2_U28 (.A( u2_u5_u2_n154 ) , .ZN( u2_u5_u2_n176 ) );
  NAND2_X1 u2_u5_u2_U29 (.A2( u2_u5_u2_n116 ) , .A1( u2_u5_u2_n117 ) , .ZN( u2_u5_u2_n118 ) );
  NOR2_X1 u2_u5_u2_U3 (.ZN( u2_u5_u2_n121 ) , .A2( u2_u5_u2_n177 ) , .A1( u2_u5_u2_n180 ) );
  INV_X1 u2_u5_u2_U30 (.A( u2_u5_u2_n132 ) , .ZN( u2_u5_u2_n182 ) );
  INV_X1 u2_u5_u2_U31 (.A( u2_u5_u2_n158 ) , .ZN( u2_u5_u2_n183 ) );
  OAI21_X1 u2_u5_u2_U32 (.A( u2_u5_u2_n156 ) , .B1( u2_u5_u2_n157 ) , .ZN( u2_u5_u2_n158 ) , .B2( u2_u5_u2_n179 ) );
  NOR2_X1 u2_u5_u2_U33 (.ZN( u2_u5_u2_n156 ) , .A1( u2_u5_u2_n166 ) , .A2( u2_u5_u2_n169 ) );
  NOR2_X1 u2_u5_u2_U34 (.A2( u2_u5_u2_n114 ) , .ZN( u2_u5_u2_n137 ) , .A1( u2_u5_u2_n140 ) );
  NOR2_X1 u2_u5_u2_U35 (.A2( u2_u5_u2_n138 ) , .ZN( u2_u5_u2_n153 ) , .A1( u2_u5_u2_n156 ) );
  AOI211_X1 u2_u5_u2_U36 (.ZN( u2_u5_u2_n130 ) , .C1( u2_u5_u2_n138 ) , .C2( u2_u5_u2_n179 ) , .B( u2_u5_u2_n96 ) , .A( u2_u5_u2_n97 ) );
  OAI22_X1 u2_u5_u2_U37 (.B1( u2_u5_u2_n133 ) , .A2( u2_u5_u2_n137 ) , .A1( u2_u5_u2_n152 ) , .B2( u2_u5_u2_n168 ) , .ZN( u2_u5_u2_n97 ) );
  OAI221_X1 u2_u5_u2_U38 (.B1( u2_u5_u2_n113 ) , .C1( u2_u5_u2_n132 ) , .A( u2_u5_u2_n149 ) , .B2( u2_u5_u2_n171 ) , .C2( u2_u5_u2_n172 ) , .ZN( u2_u5_u2_n96 ) );
  OAI221_X1 u2_u5_u2_U39 (.A( u2_u5_u2_n115 ) , .C2( u2_u5_u2_n123 ) , .B2( u2_u5_u2_n143 ) , .B1( u2_u5_u2_n153 ) , .ZN( u2_u5_u2_n163 ) , .C1( u2_u5_u2_n168 ) );
  INV_X1 u2_u5_u2_U4 (.A( u2_u5_u2_n134 ) , .ZN( u2_u5_u2_n185 ) );
  OAI21_X1 u2_u5_u2_U40 (.A( u2_u5_u2_n114 ) , .ZN( u2_u5_u2_n115 ) , .B1( u2_u5_u2_n176 ) , .B2( u2_u5_u2_n178 ) );
  OAI221_X1 u2_u5_u2_U41 (.A( u2_u5_u2_n135 ) , .B2( u2_u5_u2_n136 ) , .B1( u2_u5_u2_n137 ) , .ZN( u2_u5_u2_n162 ) , .C2( u2_u5_u2_n167 ) , .C1( u2_u5_u2_n185 ) );
  AND3_X1 u2_u5_u2_U42 (.A3( u2_u5_u2_n131 ) , .A2( u2_u5_u2_n132 ) , .A1( u2_u5_u2_n133 ) , .ZN( u2_u5_u2_n136 ) );
  AOI22_X1 u2_u5_u2_U43 (.ZN( u2_u5_u2_n135 ) , .B1( u2_u5_u2_n140 ) , .A1( u2_u5_u2_n156 ) , .B2( u2_u5_u2_n180 ) , .A2( u2_u5_u2_n188 ) );
  AOI21_X1 u2_u5_u2_U44 (.ZN( u2_u5_u2_n149 ) , .B1( u2_u5_u2_n173 ) , .B2( u2_u5_u2_n188 ) , .A( u2_u5_u2_n95 ) );
  AND3_X1 u2_u5_u2_U45 (.A2( u2_u5_u2_n100 ) , .A1( u2_u5_u2_n104 ) , .A3( u2_u5_u2_n156 ) , .ZN( u2_u5_u2_n95 ) );
  OAI21_X1 u2_u5_u2_U46 (.A( u2_u5_u2_n141 ) , .B2( u2_u5_u2_n142 ) , .ZN( u2_u5_u2_n146 ) , .B1( u2_u5_u2_n153 ) );
  OAI21_X1 u2_u5_u2_U47 (.A( u2_u5_u2_n140 ) , .ZN( u2_u5_u2_n141 ) , .B1( u2_u5_u2_n176 ) , .B2( u2_u5_u2_n177 ) );
  NOR3_X1 u2_u5_u2_U48 (.ZN( u2_u5_u2_n142 ) , .A3( u2_u5_u2_n175 ) , .A2( u2_u5_u2_n178 ) , .A1( u2_u5_u2_n181 ) );
  OAI21_X1 u2_u5_u2_U49 (.A( u2_u5_u2_n101 ) , .B2( u2_u5_u2_n121 ) , .B1( u2_u5_u2_n153 ) , .ZN( u2_u5_u2_n164 ) );
  INV_X1 u2_u5_u2_U5 (.A( u2_u5_u2_n150 ) , .ZN( u2_u5_u2_n184 ) );
  NAND2_X1 u2_u5_u2_U50 (.A2( u2_u5_u2_n100 ) , .A1( u2_u5_u2_n107 ) , .ZN( u2_u5_u2_n155 ) );
  NAND2_X1 u2_u5_u2_U51 (.A2( u2_u5_u2_n105 ) , .A1( u2_u5_u2_n108 ) , .ZN( u2_u5_u2_n143 ) );
  NAND2_X1 u2_u5_u2_U52 (.A1( u2_u5_u2_n104 ) , .A2( u2_u5_u2_n106 ) , .ZN( u2_u5_u2_n152 ) );
  NAND2_X1 u2_u5_u2_U53 (.A1( u2_u5_u2_n100 ) , .A2( u2_u5_u2_n105 ) , .ZN( u2_u5_u2_n132 ) );
  INV_X1 u2_u5_u2_U54 (.A( u2_u5_u2_n140 ) , .ZN( u2_u5_u2_n168 ) );
  INV_X1 u2_u5_u2_U55 (.A( u2_u5_u2_n138 ) , .ZN( u2_u5_u2_n167 ) );
  NAND2_X1 u2_u5_u2_U56 (.A1( u2_u5_u2_n102 ) , .A2( u2_u5_u2_n106 ) , .ZN( u2_u5_u2_n113 ) );
  NAND2_X1 u2_u5_u2_U57 (.A1( u2_u5_u2_n106 ) , .A2( u2_u5_u2_n107 ) , .ZN( u2_u5_u2_n131 ) );
  NAND2_X1 u2_u5_u2_U58 (.A1( u2_u5_u2_n103 ) , .A2( u2_u5_u2_n107 ) , .ZN( u2_u5_u2_n139 ) );
  NAND2_X1 u2_u5_u2_U59 (.A1( u2_u5_u2_n103 ) , .A2( u2_u5_u2_n105 ) , .ZN( u2_u5_u2_n133 ) );
  NOR4_X1 u2_u5_u2_U6 (.A4( u2_u5_u2_n124 ) , .A3( u2_u5_u2_n125 ) , .A2( u2_u5_u2_n126 ) , .A1( u2_u5_u2_n127 ) , .ZN( u2_u5_u2_n128 ) );
  NAND2_X1 u2_u5_u2_U60 (.A1( u2_u5_u2_n102 ) , .A2( u2_u5_u2_n103 ) , .ZN( u2_u5_u2_n154 ) );
  NAND2_X1 u2_u5_u2_U61 (.A2( u2_u5_u2_n103 ) , .A1( u2_u5_u2_n104 ) , .ZN( u2_u5_u2_n119 ) );
  NAND2_X1 u2_u5_u2_U62 (.A2( u2_u5_u2_n107 ) , .A1( u2_u5_u2_n108 ) , .ZN( u2_u5_u2_n123 ) );
  NAND2_X1 u2_u5_u2_U63 (.A1( u2_u5_u2_n104 ) , .A2( u2_u5_u2_n108 ) , .ZN( u2_u5_u2_n122 ) );
  INV_X1 u2_u5_u2_U64 (.A( u2_u5_u2_n114 ) , .ZN( u2_u5_u2_n172 ) );
  NAND2_X1 u2_u5_u2_U65 (.A2( u2_u5_u2_n100 ) , .A1( u2_u5_u2_n102 ) , .ZN( u2_u5_u2_n116 ) );
  NAND2_X1 u2_u5_u2_U66 (.A1( u2_u5_u2_n102 ) , .A2( u2_u5_u2_n108 ) , .ZN( u2_u5_u2_n120 ) );
  NAND2_X1 u2_u5_u2_U67 (.A2( u2_u5_u2_n105 ) , .A1( u2_u5_u2_n106 ) , .ZN( u2_u5_u2_n117 ) );
  INV_X1 u2_u5_u2_U68 (.ZN( u2_u5_u2_n187 ) , .A( u2_u5_u2_n99 ) );
  OAI21_X1 u2_u5_u2_U69 (.B1( u2_u5_u2_n137 ) , .B2( u2_u5_u2_n143 ) , .A( u2_u5_u2_n98 ) , .ZN( u2_u5_u2_n99 ) );
  AOI21_X1 u2_u5_u2_U7 (.B2( u2_u5_u2_n119 ) , .ZN( u2_u5_u2_n127 ) , .A( u2_u5_u2_n137 ) , .B1( u2_u5_u2_n155 ) );
  NOR2_X1 u2_u5_u2_U70 (.A2( u2_u5_X_16 ) , .ZN( u2_u5_u2_n140 ) , .A1( u2_u5_u2_n166 ) );
  NOR2_X1 u2_u5_u2_U71 (.A2( u2_u5_X_13 ) , .A1( u2_u5_X_14 ) , .ZN( u2_u5_u2_n100 ) );
  NOR2_X1 u2_u5_u2_U72 (.A2( u2_u5_X_16 ) , .A1( u2_u5_X_17 ) , .ZN( u2_u5_u2_n138 ) );
  NOR2_X1 u2_u5_u2_U73 (.A2( u2_u5_X_15 ) , .A1( u2_u5_X_18 ) , .ZN( u2_u5_u2_n104 ) );
  NOR2_X1 u2_u5_u2_U74 (.A2( u2_u5_X_14 ) , .ZN( u2_u5_u2_n103 ) , .A1( u2_u5_u2_n174 ) );
  NOR2_X1 u2_u5_u2_U75 (.A2( u2_u5_X_15 ) , .ZN( u2_u5_u2_n102 ) , .A1( u2_u5_u2_n165 ) );
  NOR2_X1 u2_u5_u2_U76 (.A2( u2_u5_X_17 ) , .ZN( u2_u5_u2_n114 ) , .A1( u2_u5_u2_n169 ) );
  AND2_X1 u2_u5_u2_U77 (.A1( u2_u5_X_15 ) , .ZN( u2_u5_u2_n105 ) , .A2( u2_u5_u2_n165 ) );
  AND2_X1 u2_u5_u2_U78 (.A2( u2_u5_X_15 ) , .A1( u2_u5_X_18 ) , .ZN( u2_u5_u2_n107 ) );
  AND2_X1 u2_u5_u2_U79 (.A1( u2_u5_X_14 ) , .ZN( u2_u5_u2_n106 ) , .A2( u2_u5_u2_n174 ) );
  AOI21_X1 u2_u5_u2_U8 (.ZN( u2_u5_u2_n124 ) , .B1( u2_u5_u2_n131 ) , .B2( u2_u5_u2_n143 ) , .A( u2_u5_u2_n172 ) );
  AND2_X1 u2_u5_u2_U80 (.A1( u2_u5_X_13 ) , .A2( u2_u5_X_14 ) , .ZN( u2_u5_u2_n108 ) );
  INV_X1 u2_u5_u2_U81 (.A( u2_u5_X_16 ) , .ZN( u2_u5_u2_n169 ) );
  INV_X1 u2_u5_u2_U82 (.A( u2_u5_X_17 ) , .ZN( u2_u5_u2_n166 ) );
  INV_X1 u2_u5_u2_U83 (.A( u2_u5_X_13 ) , .ZN( u2_u5_u2_n174 ) );
  INV_X1 u2_u5_u2_U84 (.A( u2_u5_X_18 ) , .ZN( u2_u5_u2_n165 ) );
  NAND4_X1 u2_u5_u2_U85 (.ZN( u2_out5_24 ) , .A4( u2_u5_u2_n111 ) , .A3( u2_u5_u2_n112 ) , .A1( u2_u5_u2_n130 ) , .A2( u2_u5_u2_n187 ) );
  AOI221_X1 u2_u5_u2_U86 (.A( u2_u5_u2_n109 ) , .B1( u2_u5_u2_n110 ) , .ZN( u2_u5_u2_n111 ) , .C1( u2_u5_u2_n134 ) , .C2( u2_u5_u2_n170 ) , .B2( u2_u5_u2_n173 ) );
  AOI21_X1 u2_u5_u2_U87 (.ZN( u2_u5_u2_n112 ) , .B2( u2_u5_u2_n156 ) , .A( u2_u5_u2_n164 ) , .B1( u2_u5_u2_n181 ) );
  NAND4_X1 u2_u5_u2_U88 (.ZN( u2_out5_16 ) , .A4( u2_u5_u2_n128 ) , .A3( u2_u5_u2_n129 ) , .A1( u2_u5_u2_n130 ) , .A2( u2_u5_u2_n186 ) );
  AOI22_X1 u2_u5_u2_U89 (.A2( u2_u5_u2_n118 ) , .ZN( u2_u5_u2_n129 ) , .A1( u2_u5_u2_n140 ) , .B1( u2_u5_u2_n157 ) , .B2( u2_u5_u2_n170 ) );
  AOI21_X1 u2_u5_u2_U9 (.B2( u2_u5_u2_n123 ) , .ZN( u2_u5_u2_n125 ) , .A( u2_u5_u2_n171 ) , .B1( u2_u5_u2_n184 ) );
  INV_X1 u2_u5_u2_U90 (.A( u2_u5_u2_n163 ) , .ZN( u2_u5_u2_n186 ) );
  NAND4_X1 u2_u5_u2_U91 (.ZN( u2_out5_30 ) , .A4( u2_u5_u2_n147 ) , .A3( u2_u5_u2_n148 ) , .A2( u2_u5_u2_n149 ) , .A1( u2_u5_u2_n187 ) );
  NOR3_X1 u2_u5_u2_U92 (.A3( u2_u5_u2_n144 ) , .A2( u2_u5_u2_n145 ) , .A1( u2_u5_u2_n146 ) , .ZN( u2_u5_u2_n147 ) );
  AOI21_X1 u2_u5_u2_U93 (.B2( u2_u5_u2_n138 ) , .ZN( u2_u5_u2_n148 ) , .A( u2_u5_u2_n162 ) , .B1( u2_u5_u2_n182 ) );
  OR4_X1 u2_u5_u2_U94 (.ZN( u2_out5_6 ) , .A4( u2_u5_u2_n161 ) , .A3( u2_u5_u2_n162 ) , .A2( u2_u5_u2_n163 ) , .A1( u2_u5_u2_n164 ) );
  OR3_X1 u2_u5_u2_U95 (.A2( u2_u5_u2_n159 ) , .A1( u2_u5_u2_n160 ) , .ZN( u2_u5_u2_n161 ) , .A3( u2_u5_u2_n183 ) );
  AOI21_X1 u2_u5_u2_U96 (.B2( u2_u5_u2_n154 ) , .B1( u2_u5_u2_n155 ) , .ZN( u2_u5_u2_n159 ) , .A( u2_u5_u2_n167 ) );
  NAND3_X1 u2_u5_u2_U97 (.A2( u2_u5_u2_n117 ) , .A1( u2_u5_u2_n122 ) , .A3( u2_u5_u2_n123 ) , .ZN( u2_u5_u2_n134 ) );
  NAND3_X1 u2_u5_u2_U98 (.ZN( u2_u5_u2_n110 ) , .A2( u2_u5_u2_n131 ) , .A3( u2_u5_u2_n139 ) , .A1( u2_u5_u2_n154 ) );
  NAND3_X1 u2_u5_u2_U99 (.A2( u2_u5_u2_n100 ) , .ZN( u2_u5_u2_n101 ) , .A1( u2_u5_u2_n104 ) , .A3( u2_u5_u2_n114 ) );
  OAI22_X1 u2_u5_u3_U10 (.B1( u2_u5_u3_n113 ) , .A2( u2_u5_u3_n135 ) , .A1( u2_u5_u3_n150 ) , .B2( u2_u5_u3_n164 ) , .ZN( u2_u5_u3_n98 ) );
  OAI211_X1 u2_u5_u3_U11 (.B( u2_u5_u3_n106 ) , .ZN( u2_u5_u3_n119 ) , .C2( u2_u5_u3_n128 ) , .C1( u2_u5_u3_n167 ) , .A( u2_u5_u3_n181 ) );
  AOI221_X1 u2_u5_u3_U12 (.C1( u2_u5_u3_n105 ) , .ZN( u2_u5_u3_n106 ) , .A( u2_u5_u3_n131 ) , .B2( u2_u5_u3_n132 ) , .C2( u2_u5_u3_n133 ) , .B1( u2_u5_u3_n169 ) );
  INV_X1 u2_u5_u3_U13 (.ZN( u2_u5_u3_n181 ) , .A( u2_u5_u3_n98 ) );
  NAND2_X1 u2_u5_u3_U14 (.ZN( u2_u5_u3_n105 ) , .A2( u2_u5_u3_n130 ) , .A1( u2_u5_u3_n155 ) );
  AOI22_X1 u2_u5_u3_U15 (.B1( u2_u5_u3_n115 ) , .A2( u2_u5_u3_n116 ) , .ZN( u2_u5_u3_n123 ) , .B2( u2_u5_u3_n133 ) , .A1( u2_u5_u3_n169 ) );
  NAND2_X1 u2_u5_u3_U16 (.ZN( u2_u5_u3_n116 ) , .A2( u2_u5_u3_n151 ) , .A1( u2_u5_u3_n182 ) );
  NOR2_X1 u2_u5_u3_U17 (.ZN( u2_u5_u3_n126 ) , .A2( u2_u5_u3_n150 ) , .A1( u2_u5_u3_n164 ) );
  AOI21_X1 u2_u5_u3_U18 (.ZN( u2_u5_u3_n112 ) , .B2( u2_u5_u3_n146 ) , .B1( u2_u5_u3_n155 ) , .A( u2_u5_u3_n167 ) );
  NAND2_X1 u2_u5_u3_U19 (.A1( u2_u5_u3_n135 ) , .ZN( u2_u5_u3_n142 ) , .A2( u2_u5_u3_n164 ) );
  NAND2_X1 u2_u5_u3_U20 (.ZN( u2_u5_u3_n132 ) , .A2( u2_u5_u3_n152 ) , .A1( u2_u5_u3_n156 ) );
  AND2_X1 u2_u5_u3_U21 (.A2( u2_u5_u3_n113 ) , .A1( u2_u5_u3_n114 ) , .ZN( u2_u5_u3_n151 ) );
  INV_X1 u2_u5_u3_U22 (.A( u2_u5_u3_n133 ) , .ZN( u2_u5_u3_n165 ) );
  INV_X1 u2_u5_u3_U23 (.A( u2_u5_u3_n135 ) , .ZN( u2_u5_u3_n170 ) );
  NAND2_X1 u2_u5_u3_U24 (.A1( u2_u5_u3_n107 ) , .A2( u2_u5_u3_n108 ) , .ZN( u2_u5_u3_n140 ) );
  NAND2_X1 u2_u5_u3_U25 (.ZN( u2_u5_u3_n117 ) , .A1( u2_u5_u3_n124 ) , .A2( u2_u5_u3_n148 ) );
  NAND2_X1 u2_u5_u3_U26 (.ZN( u2_u5_u3_n143 ) , .A1( u2_u5_u3_n165 ) , .A2( u2_u5_u3_n167 ) );
  INV_X1 u2_u5_u3_U27 (.A( u2_u5_u3_n130 ) , .ZN( u2_u5_u3_n177 ) );
  INV_X1 u2_u5_u3_U28 (.A( u2_u5_u3_n128 ) , .ZN( u2_u5_u3_n176 ) );
  INV_X1 u2_u5_u3_U29 (.A( u2_u5_u3_n155 ) , .ZN( u2_u5_u3_n174 ) );
  INV_X1 u2_u5_u3_U3 (.A( u2_u5_u3_n129 ) , .ZN( u2_u5_u3_n183 ) );
  INV_X1 u2_u5_u3_U30 (.A( u2_u5_u3_n139 ) , .ZN( u2_u5_u3_n185 ) );
  NOR2_X1 u2_u5_u3_U31 (.ZN( u2_u5_u3_n135 ) , .A2( u2_u5_u3_n141 ) , .A1( u2_u5_u3_n169 ) );
  OAI222_X1 u2_u5_u3_U32 (.C2( u2_u5_u3_n107 ) , .A2( u2_u5_u3_n108 ) , .B1( u2_u5_u3_n135 ) , .ZN( u2_u5_u3_n138 ) , .B2( u2_u5_u3_n146 ) , .C1( u2_u5_u3_n154 ) , .A1( u2_u5_u3_n164 ) );
  NOR4_X1 u2_u5_u3_U33 (.A4( u2_u5_u3_n157 ) , .A3( u2_u5_u3_n158 ) , .A2( u2_u5_u3_n159 ) , .A1( u2_u5_u3_n160 ) , .ZN( u2_u5_u3_n161 ) );
  AOI21_X1 u2_u5_u3_U34 (.B2( u2_u5_u3_n152 ) , .B1( u2_u5_u3_n153 ) , .ZN( u2_u5_u3_n158 ) , .A( u2_u5_u3_n164 ) );
  AOI21_X1 u2_u5_u3_U35 (.A( u2_u5_u3_n154 ) , .B2( u2_u5_u3_n155 ) , .B1( u2_u5_u3_n156 ) , .ZN( u2_u5_u3_n157 ) );
  AOI21_X1 u2_u5_u3_U36 (.A( u2_u5_u3_n149 ) , .B2( u2_u5_u3_n150 ) , .B1( u2_u5_u3_n151 ) , .ZN( u2_u5_u3_n159 ) );
  AOI211_X1 u2_u5_u3_U37 (.ZN( u2_u5_u3_n109 ) , .A( u2_u5_u3_n119 ) , .C2( u2_u5_u3_n129 ) , .B( u2_u5_u3_n138 ) , .C1( u2_u5_u3_n141 ) );
  AOI211_X1 u2_u5_u3_U38 (.B( u2_u5_u3_n119 ) , .A( u2_u5_u3_n120 ) , .C2( u2_u5_u3_n121 ) , .ZN( u2_u5_u3_n122 ) , .C1( u2_u5_u3_n179 ) );
  INV_X1 u2_u5_u3_U39 (.A( u2_u5_u3_n156 ) , .ZN( u2_u5_u3_n179 ) );
  INV_X1 u2_u5_u3_U4 (.A( u2_u5_u3_n140 ) , .ZN( u2_u5_u3_n182 ) );
  OAI22_X1 u2_u5_u3_U40 (.B1( u2_u5_u3_n118 ) , .ZN( u2_u5_u3_n120 ) , .A1( u2_u5_u3_n135 ) , .B2( u2_u5_u3_n154 ) , .A2( u2_u5_u3_n178 ) );
  AND3_X1 u2_u5_u3_U41 (.ZN( u2_u5_u3_n118 ) , .A2( u2_u5_u3_n124 ) , .A1( u2_u5_u3_n144 ) , .A3( u2_u5_u3_n152 ) );
  INV_X1 u2_u5_u3_U42 (.A( u2_u5_u3_n121 ) , .ZN( u2_u5_u3_n164 ) );
  NAND2_X1 u2_u5_u3_U43 (.ZN( u2_u5_u3_n133 ) , .A1( u2_u5_u3_n154 ) , .A2( u2_u5_u3_n164 ) );
  OAI211_X1 u2_u5_u3_U44 (.B( u2_u5_u3_n127 ) , .ZN( u2_u5_u3_n139 ) , .C1( u2_u5_u3_n150 ) , .C2( u2_u5_u3_n154 ) , .A( u2_u5_u3_n184 ) );
  INV_X1 u2_u5_u3_U45 (.A( u2_u5_u3_n125 ) , .ZN( u2_u5_u3_n184 ) );
  AOI221_X1 u2_u5_u3_U46 (.A( u2_u5_u3_n126 ) , .ZN( u2_u5_u3_n127 ) , .C2( u2_u5_u3_n132 ) , .C1( u2_u5_u3_n169 ) , .B2( u2_u5_u3_n170 ) , .B1( u2_u5_u3_n174 ) );
  OAI22_X1 u2_u5_u3_U47 (.A1( u2_u5_u3_n124 ) , .ZN( u2_u5_u3_n125 ) , .B2( u2_u5_u3_n145 ) , .A2( u2_u5_u3_n165 ) , .B1( u2_u5_u3_n167 ) );
  NOR2_X1 u2_u5_u3_U48 (.A1( u2_u5_u3_n113 ) , .ZN( u2_u5_u3_n131 ) , .A2( u2_u5_u3_n154 ) );
  NAND2_X1 u2_u5_u3_U49 (.A1( u2_u5_u3_n103 ) , .ZN( u2_u5_u3_n150 ) , .A2( u2_u5_u3_n99 ) );
  INV_X1 u2_u5_u3_U5 (.A( u2_u5_u3_n117 ) , .ZN( u2_u5_u3_n178 ) );
  NAND2_X1 u2_u5_u3_U50 (.A2( u2_u5_u3_n102 ) , .ZN( u2_u5_u3_n155 ) , .A1( u2_u5_u3_n97 ) );
  INV_X1 u2_u5_u3_U51 (.A( u2_u5_u3_n141 ) , .ZN( u2_u5_u3_n167 ) );
  AOI21_X1 u2_u5_u3_U52 (.B2( u2_u5_u3_n114 ) , .B1( u2_u5_u3_n146 ) , .A( u2_u5_u3_n154 ) , .ZN( u2_u5_u3_n94 ) );
  AOI21_X1 u2_u5_u3_U53 (.ZN( u2_u5_u3_n110 ) , .B2( u2_u5_u3_n142 ) , .B1( u2_u5_u3_n186 ) , .A( u2_u5_u3_n95 ) );
  INV_X1 u2_u5_u3_U54 (.A( u2_u5_u3_n145 ) , .ZN( u2_u5_u3_n186 ) );
  AOI21_X1 u2_u5_u3_U55 (.B1( u2_u5_u3_n124 ) , .A( u2_u5_u3_n149 ) , .B2( u2_u5_u3_n155 ) , .ZN( u2_u5_u3_n95 ) );
  INV_X1 u2_u5_u3_U56 (.A( u2_u5_u3_n149 ) , .ZN( u2_u5_u3_n169 ) );
  NAND2_X1 u2_u5_u3_U57 (.ZN( u2_u5_u3_n124 ) , .A1( u2_u5_u3_n96 ) , .A2( u2_u5_u3_n97 ) );
  NAND2_X1 u2_u5_u3_U58 (.A2( u2_u5_u3_n100 ) , .ZN( u2_u5_u3_n146 ) , .A1( u2_u5_u3_n96 ) );
  NAND2_X1 u2_u5_u3_U59 (.A1( u2_u5_u3_n101 ) , .ZN( u2_u5_u3_n145 ) , .A2( u2_u5_u3_n99 ) );
  AOI221_X1 u2_u5_u3_U6 (.A( u2_u5_u3_n131 ) , .C2( u2_u5_u3_n132 ) , .C1( u2_u5_u3_n133 ) , .ZN( u2_u5_u3_n134 ) , .B1( u2_u5_u3_n143 ) , .B2( u2_u5_u3_n177 ) );
  NAND2_X1 u2_u5_u3_U60 (.A1( u2_u5_u3_n100 ) , .ZN( u2_u5_u3_n156 ) , .A2( u2_u5_u3_n99 ) );
  NAND2_X1 u2_u5_u3_U61 (.A2( u2_u5_u3_n101 ) , .A1( u2_u5_u3_n104 ) , .ZN( u2_u5_u3_n148 ) );
  NAND2_X1 u2_u5_u3_U62 (.A1( u2_u5_u3_n100 ) , .A2( u2_u5_u3_n102 ) , .ZN( u2_u5_u3_n128 ) );
  NAND2_X1 u2_u5_u3_U63 (.A2( u2_u5_u3_n101 ) , .A1( u2_u5_u3_n102 ) , .ZN( u2_u5_u3_n152 ) );
  NAND2_X1 u2_u5_u3_U64 (.A2( u2_u5_u3_n101 ) , .ZN( u2_u5_u3_n114 ) , .A1( u2_u5_u3_n96 ) );
  NAND2_X1 u2_u5_u3_U65 (.ZN( u2_u5_u3_n107 ) , .A1( u2_u5_u3_n97 ) , .A2( u2_u5_u3_n99 ) );
  NAND2_X1 u2_u5_u3_U66 (.A2( u2_u5_u3_n100 ) , .A1( u2_u5_u3_n104 ) , .ZN( u2_u5_u3_n113 ) );
  NAND2_X1 u2_u5_u3_U67 (.A1( u2_u5_u3_n104 ) , .ZN( u2_u5_u3_n153 ) , .A2( u2_u5_u3_n97 ) );
  NAND2_X1 u2_u5_u3_U68 (.A2( u2_u5_u3_n103 ) , .A1( u2_u5_u3_n104 ) , .ZN( u2_u5_u3_n130 ) );
  NAND2_X1 u2_u5_u3_U69 (.A2( u2_u5_u3_n103 ) , .ZN( u2_u5_u3_n144 ) , .A1( u2_u5_u3_n96 ) );
  OAI22_X1 u2_u5_u3_U7 (.B2( u2_u5_u3_n147 ) , .A2( u2_u5_u3_n148 ) , .ZN( u2_u5_u3_n160 ) , .B1( u2_u5_u3_n165 ) , .A1( u2_u5_u3_n168 ) );
  NAND2_X1 u2_u5_u3_U70 (.A1( u2_u5_u3_n102 ) , .A2( u2_u5_u3_n103 ) , .ZN( u2_u5_u3_n108 ) );
  NOR2_X1 u2_u5_u3_U71 (.A2( u2_u5_X_19 ) , .A1( u2_u5_X_20 ) , .ZN( u2_u5_u3_n99 ) );
  NOR2_X1 u2_u5_u3_U72 (.A2( u2_u5_X_21 ) , .A1( u2_u5_X_24 ) , .ZN( u2_u5_u3_n103 ) );
  NOR2_X1 u2_u5_u3_U73 (.A2( u2_u5_X_24 ) , .A1( u2_u5_u3_n171 ) , .ZN( u2_u5_u3_n97 ) );
  NOR2_X1 u2_u5_u3_U74 (.A2( u2_u5_X_23 ) , .ZN( u2_u5_u3_n141 ) , .A1( u2_u5_u3_n166 ) );
  NOR2_X1 u2_u5_u3_U75 (.A2( u2_u5_X_19 ) , .A1( u2_u5_u3_n172 ) , .ZN( u2_u5_u3_n96 ) );
  NAND2_X1 u2_u5_u3_U76 (.A1( u2_u5_X_22 ) , .A2( u2_u5_X_23 ) , .ZN( u2_u5_u3_n154 ) );
  NAND2_X1 u2_u5_u3_U77 (.A1( u2_u5_X_23 ) , .ZN( u2_u5_u3_n149 ) , .A2( u2_u5_u3_n166 ) );
  NOR2_X1 u2_u5_u3_U78 (.A2( u2_u5_X_22 ) , .A1( u2_u5_X_23 ) , .ZN( u2_u5_u3_n121 ) );
  AND2_X1 u2_u5_u3_U79 (.A1( u2_u5_X_24 ) , .ZN( u2_u5_u3_n101 ) , .A2( u2_u5_u3_n171 ) );
  AND3_X1 u2_u5_u3_U8 (.A3( u2_u5_u3_n144 ) , .A2( u2_u5_u3_n145 ) , .A1( u2_u5_u3_n146 ) , .ZN( u2_u5_u3_n147 ) );
  AND2_X1 u2_u5_u3_U80 (.A1( u2_u5_X_19 ) , .ZN( u2_u5_u3_n102 ) , .A2( u2_u5_u3_n172 ) );
  AND2_X1 u2_u5_u3_U81 (.A1( u2_u5_X_21 ) , .A2( u2_u5_X_24 ) , .ZN( u2_u5_u3_n100 ) );
  AND2_X1 u2_u5_u3_U82 (.A2( u2_u5_X_19 ) , .A1( u2_u5_X_20 ) , .ZN( u2_u5_u3_n104 ) );
  INV_X1 u2_u5_u3_U83 (.A( u2_u5_X_22 ) , .ZN( u2_u5_u3_n166 ) );
  INV_X1 u2_u5_u3_U84 (.A( u2_u5_X_21 ) , .ZN( u2_u5_u3_n171 ) );
  INV_X1 u2_u5_u3_U85 (.A( u2_u5_X_20 ) , .ZN( u2_u5_u3_n172 ) );
  NAND4_X1 u2_u5_u3_U86 (.ZN( u2_out5_26 ) , .A4( u2_u5_u3_n109 ) , .A3( u2_u5_u3_n110 ) , .A2( u2_u5_u3_n111 ) , .A1( u2_u5_u3_n173 ) );
  INV_X1 u2_u5_u3_U87 (.ZN( u2_u5_u3_n173 ) , .A( u2_u5_u3_n94 ) );
  OAI21_X1 u2_u5_u3_U88 (.ZN( u2_u5_u3_n111 ) , .B2( u2_u5_u3_n117 ) , .A( u2_u5_u3_n133 ) , .B1( u2_u5_u3_n176 ) );
  NAND4_X1 u2_u5_u3_U89 (.ZN( u2_out5_20 ) , .A4( u2_u5_u3_n122 ) , .A3( u2_u5_u3_n123 ) , .A1( u2_u5_u3_n175 ) , .A2( u2_u5_u3_n180 ) );
  INV_X1 u2_u5_u3_U9 (.A( u2_u5_u3_n143 ) , .ZN( u2_u5_u3_n168 ) );
  INV_X1 u2_u5_u3_U90 (.A( u2_u5_u3_n126 ) , .ZN( u2_u5_u3_n180 ) );
  INV_X1 u2_u5_u3_U91 (.A( u2_u5_u3_n112 ) , .ZN( u2_u5_u3_n175 ) );
  NAND4_X1 u2_u5_u3_U92 (.ZN( u2_out5_1 ) , .A4( u2_u5_u3_n161 ) , .A3( u2_u5_u3_n162 ) , .A2( u2_u5_u3_n163 ) , .A1( u2_u5_u3_n185 ) );
  NAND2_X1 u2_u5_u3_U93 (.ZN( u2_u5_u3_n163 ) , .A2( u2_u5_u3_n170 ) , .A1( u2_u5_u3_n176 ) );
  AOI22_X1 u2_u5_u3_U94 (.B2( u2_u5_u3_n140 ) , .B1( u2_u5_u3_n141 ) , .A2( u2_u5_u3_n142 ) , .ZN( u2_u5_u3_n162 ) , .A1( u2_u5_u3_n177 ) );
  OR4_X1 u2_u5_u3_U95 (.ZN( u2_out5_10 ) , .A4( u2_u5_u3_n136 ) , .A3( u2_u5_u3_n137 ) , .A1( u2_u5_u3_n138 ) , .A2( u2_u5_u3_n139 ) );
  OAI222_X1 u2_u5_u3_U96 (.C1( u2_u5_u3_n128 ) , .ZN( u2_u5_u3_n137 ) , .B1( u2_u5_u3_n148 ) , .A2( u2_u5_u3_n150 ) , .B2( u2_u5_u3_n154 ) , .C2( u2_u5_u3_n164 ) , .A1( u2_u5_u3_n167 ) );
  OAI221_X1 u2_u5_u3_U97 (.A( u2_u5_u3_n134 ) , .B2( u2_u5_u3_n135 ) , .ZN( u2_u5_u3_n136 ) , .C1( u2_u5_u3_n149 ) , .B1( u2_u5_u3_n151 ) , .C2( u2_u5_u3_n183 ) );
  NAND3_X1 u2_u5_u3_U98 (.A1( u2_u5_u3_n114 ) , .ZN( u2_u5_u3_n115 ) , .A2( u2_u5_u3_n145 ) , .A3( u2_u5_u3_n153 ) );
  NAND3_X1 u2_u5_u3_U99 (.ZN( u2_u5_u3_n129 ) , .A2( u2_u5_u3_n144 ) , .A1( u2_u5_u3_n153 ) , .A3( u2_u5_u3_n182 ) );
  OAI22_X1 u2_u5_u4_U10 (.B2( u2_u5_u4_n135 ) , .ZN( u2_u5_u4_n137 ) , .B1( u2_u5_u4_n153 ) , .A1( u2_u5_u4_n155 ) , .A2( u2_u5_u4_n171 ) );
  AND3_X1 u2_u5_u4_U11 (.A2( u2_u5_u4_n134 ) , .ZN( u2_u5_u4_n135 ) , .A3( u2_u5_u4_n145 ) , .A1( u2_u5_u4_n157 ) );
  NAND2_X1 u2_u5_u4_U12 (.ZN( u2_u5_u4_n132 ) , .A2( u2_u5_u4_n170 ) , .A1( u2_u5_u4_n173 ) );
  AOI21_X1 u2_u5_u4_U13 (.B2( u2_u5_u4_n160 ) , .B1( u2_u5_u4_n161 ) , .ZN( u2_u5_u4_n162 ) , .A( u2_u5_u4_n170 ) );
  AOI21_X1 u2_u5_u4_U14 (.ZN( u2_u5_u4_n107 ) , .B2( u2_u5_u4_n143 ) , .A( u2_u5_u4_n174 ) , .B1( u2_u5_u4_n184 ) );
  AOI21_X1 u2_u5_u4_U15 (.B2( u2_u5_u4_n158 ) , .B1( u2_u5_u4_n159 ) , .ZN( u2_u5_u4_n163 ) , .A( u2_u5_u4_n174 ) );
  AOI21_X1 u2_u5_u4_U16 (.A( u2_u5_u4_n153 ) , .B2( u2_u5_u4_n154 ) , .B1( u2_u5_u4_n155 ) , .ZN( u2_u5_u4_n165 ) );
  AOI21_X1 u2_u5_u4_U17 (.A( u2_u5_u4_n156 ) , .B2( u2_u5_u4_n157 ) , .ZN( u2_u5_u4_n164 ) , .B1( u2_u5_u4_n184 ) );
  INV_X1 u2_u5_u4_U18 (.A( u2_u5_u4_n138 ) , .ZN( u2_u5_u4_n170 ) );
  AND2_X1 u2_u5_u4_U19 (.A2( u2_u5_u4_n120 ) , .ZN( u2_u5_u4_n155 ) , .A1( u2_u5_u4_n160 ) );
  INV_X1 u2_u5_u4_U20 (.A( u2_u5_u4_n156 ) , .ZN( u2_u5_u4_n175 ) );
  NAND2_X1 u2_u5_u4_U21 (.A2( u2_u5_u4_n118 ) , .ZN( u2_u5_u4_n131 ) , .A1( u2_u5_u4_n147 ) );
  NAND2_X1 u2_u5_u4_U22 (.A1( u2_u5_u4_n119 ) , .A2( u2_u5_u4_n120 ) , .ZN( u2_u5_u4_n130 ) );
  NAND2_X1 u2_u5_u4_U23 (.ZN( u2_u5_u4_n117 ) , .A2( u2_u5_u4_n118 ) , .A1( u2_u5_u4_n148 ) );
  NAND2_X1 u2_u5_u4_U24 (.ZN( u2_u5_u4_n129 ) , .A1( u2_u5_u4_n134 ) , .A2( u2_u5_u4_n148 ) );
  AND3_X1 u2_u5_u4_U25 (.A1( u2_u5_u4_n119 ) , .A2( u2_u5_u4_n143 ) , .A3( u2_u5_u4_n154 ) , .ZN( u2_u5_u4_n161 ) );
  AND2_X1 u2_u5_u4_U26 (.A1( u2_u5_u4_n145 ) , .A2( u2_u5_u4_n147 ) , .ZN( u2_u5_u4_n159 ) );
  OR3_X1 u2_u5_u4_U27 (.A3( u2_u5_u4_n114 ) , .A2( u2_u5_u4_n115 ) , .A1( u2_u5_u4_n116 ) , .ZN( u2_u5_u4_n136 ) );
  AOI21_X1 u2_u5_u4_U28 (.A( u2_u5_u4_n113 ) , .ZN( u2_u5_u4_n116 ) , .B2( u2_u5_u4_n173 ) , .B1( u2_u5_u4_n174 ) );
  AOI21_X1 u2_u5_u4_U29 (.ZN( u2_u5_u4_n115 ) , .B2( u2_u5_u4_n145 ) , .B1( u2_u5_u4_n146 ) , .A( u2_u5_u4_n156 ) );
  NOR2_X1 u2_u5_u4_U3 (.ZN( u2_u5_u4_n121 ) , .A1( u2_u5_u4_n181 ) , .A2( u2_u5_u4_n182 ) );
  OAI22_X1 u2_u5_u4_U30 (.ZN( u2_u5_u4_n114 ) , .A2( u2_u5_u4_n121 ) , .B1( u2_u5_u4_n160 ) , .B2( u2_u5_u4_n170 ) , .A1( u2_u5_u4_n171 ) );
  INV_X1 u2_u5_u4_U31 (.A( u2_u5_u4_n158 ) , .ZN( u2_u5_u4_n182 ) );
  INV_X1 u2_u5_u4_U32 (.ZN( u2_u5_u4_n181 ) , .A( u2_u5_u4_n96 ) );
  INV_X1 u2_u5_u4_U33 (.A( u2_u5_u4_n144 ) , .ZN( u2_u5_u4_n179 ) );
  INV_X1 u2_u5_u4_U34 (.A( u2_u5_u4_n157 ) , .ZN( u2_u5_u4_n178 ) );
  NAND2_X1 u2_u5_u4_U35 (.A2( u2_u5_u4_n154 ) , .A1( u2_u5_u4_n96 ) , .ZN( u2_u5_u4_n97 ) );
  INV_X1 u2_u5_u4_U36 (.ZN( u2_u5_u4_n186 ) , .A( u2_u5_u4_n95 ) );
  OAI221_X1 u2_u5_u4_U37 (.C1( u2_u5_u4_n134 ) , .B1( u2_u5_u4_n158 ) , .B2( u2_u5_u4_n171 ) , .C2( u2_u5_u4_n173 ) , .A( u2_u5_u4_n94 ) , .ZN( u2_u5_u4_n95 ) );
  AOI222_X1 u2_u5_u4_U38 (.B2( u2_u5_u4_n132 ) , .A1( u2_u5_u4_n138 ) , .C2( u2_u5_u4_n175 ) , .A2( u2_u5_u4_n179 ) , .C1( u2_u5_u4_n181 ) , .B1( u2_u5_u4_n185 ) , .ZN( u2_u5_u4_n94 ) );
  INV_X1 u2_u5_u4_U39 (.A( u2_u5_u4_n113 ) , .ZN( u2_u5_u4_n185 ) );
  INV_X1 u2_u5_u4_U4 (.A( u2_u5_u4_n117 ) , .ZN( u2_u5_u4_n184 ) );
  INV_X1 u2_u5_u4_U40 (.A( u2_u5_u4_n143 ) , .ZN( u2_u5_u4_n183 ) );
  NOR2_X1 u2_u5_u4_U41 (.ZN( u2_u5_u4_n138 ) , .A1( u2_u5_u4_n168 ) , .A2( u2_u5_u4_n169 ) );
  NOR2_X1 u2_u5_u4_U42 (.A1( u2_u5_u4_n150 ) , .A2( u2_u5_u4_n152 ) , .ZN( u2_u5_u4_n153 ) );
  NOR2_X1 u2_u5_u4_U43 (.A2( u2_u5_u4_n128 ) , .A1( u2_u5_u4_n138 ) , .ZN( u2_u5_u4_n156 ) );
  AOI22_X1 u2_u5_u4_U44 (.B2( u2_u5_u4_n122 ) , .A1( u2_u5_u4_n123 ) , .ZN( u2_u5_u4_n124 ) , .B1( u2_u5_u4_n128 ) , .A2( u2_u5_u4_n172 ) );
  INV_X1 u2_u5_u4_U45 (.A( u2_u5_u4_n153 ) , .ZN( u2_u5_u4_n172 ) );
  NAND2_X1 u2_u5_u4_U46 (.A2( u2_u5_u4_n120 ) , .ZN( u2_u5_u4_n123 ) , .A1( u2_u5_u4_n161 ) );
  AOI22_X1 u2_u5_u4_U47 (.B2( u2_u5_u4_n132 ) , .A2( u2_u5_u4_n133 ) , .ZN( u2_u5_u4_n140 ) , .A1( u2_u5_u4_n150 ) , .B1( u2_u5_u4_n179 ) );
  NAND2_X1 u2_u5_u4_U48 (.ZN( u2_u5_u4_n133 ) , .A2( u2_u5_u4_n146 ) , .A1( u2_u5_u4_n154 ) );
  NAND2_X1 u2_u5_u4_U49 (.A1( u2_u5_u4_n103 ) , .ZN( u2_u5_u4_n154 ) , .A2( u2_u5_u4_n98 ) );
  NOR4_X1 u2_u5_u4_U5 (.A4( u2_u5_u4_n106 ) , .A3( u2_u5_u4_n107 ) , .A2( u2_u5_u4_n108 ) , .A1( u2_u5_u4_n109 ) , .ZN( u2_u5_u4_n110 ) );
  NAND2_X1 u2_u5_u4_U50 (.A1( u2_u5_u4_n101 ) , .ZN( u2_u5_u4_n158 ) , .A2( u2_u5_u4_n99 ) );
  AOI21_X1 u2_u5_u4_U51 (.ZN( u2_u5_u4_n127 ) , .A( u2_u5_u4_n136 ) , .B2( u2_u5_u4_n150 ) , .B1( u2_u5_u4_n180 ) );
  INV_X1 u2_u5_u4_U52 (.A( u2_u5_u4_n160 ) , .ZN( u2_u5_u4_n180 ) );
  NAND2_X1 u2_u5_u4_U53 (.A2( u2_u5_u4_n104 ) , .A1( u2_u5_u4_n105 ) , .ZN( u2_u5_u4_n146 ) );
  NAND2_X1 u2_u5_u4_U54 (.A2( u2_u5_u4_n101 ) , .A1( u2_u5_u4_n102 ) , .ZN( u2_u5_u4_n160 ) );
  NAND2_X1 u2_u5_u4_U55 (.ZN( u2_u5_u4_n134 ) , .A1( u2_u5_u4_n98 ) , .A2( u2_u5_u4_n99 ) );
  NAND2_X1 u2_u5_u4_U56 (.A1( u2_u5_u4_n103 ) , .A2( u2_u5_u4_n104 ) , .ZN( u2_u5_u4_n143 ) );
  NAND2_X1 u2_u5_u4_U57 (.A2( u2_u5_u4_n105 ) , .ZN( u2_u5_u4_n145 ) , .A1( u2_u5_u4_n98 ) );
  NAND2_X1 u2_u5_u4_U58 (.A1( u2_u5_u4_n100 ) , .A2( u2_u5_u4_n105 ) , .ZN( u2_u5_u4_n120 ) );
  NAND2_X1 u2_u5_u4_U59 (.A1( u2_u5_u4_n102 ) , .A2( u2_u5_u4_n104 ) , .ZN( u2_u5_u4_n148 ) );
  AOI21_X1 u2_u5_u4_U6 (.ZN( u2_u5_u4_n106 ) , .B2( u2_u5_u4_n146 ) , .B1( u2_u5_u4_n158 ) , .A( u2_u5_u4_n170 ) );
  NAND2_X1 u2_u5_u4_U60 (.A2( u2_u5_u4_n100 ) , .A1( u2_u5_u4_n103 ) , .ZN( u2_u5_u4_n157 ) );
  INV_X1 u2_u5_u4_U61 (.A( u2_u5_u4_n150 ) , .ZN( u2_u5_u4_n173 ) );
  INV_X1 u2_u5_u4_U62 (.A( u2_u5_u4_n152 ) , .ZN( u2_u5_u4_n171 ) );
  NAND2_X1 u2_u5_u4_U63 (.A1( u2_u5_u4_n100 ) , .ZN( u2_u5_u4_n118 ) , .A2( u2_u5_u4_n99 ) );
  NAND2_X1 u2_u5_u4_U64 (.A2( u2_u5_u4_n100 ) , .A1( u2_u5_u4_n102 ) , .ZN( u2_u5_u4_n144 ) );
  NAND2_X1 u2_u5_u4_U65 (.A2( u2_u5_u4_n101 ) , .A1( u2_u5_u4_n105 ) , .ZN( u2_u5_u4_n96 ) );
  INV_X1 u2_u5_u4_U66 (.A( u2_u5_u4_n128 ) , .ZN( u2_u5_u4_n174 ) );
  NAND2_X1 u2_u5_u4_U67 (.A2( u2_u5_u4_n102 ) , .ZN( u2_u5_u4_n119 ) , .A1( u2_u5_u4_n98 ) );
  NAND2_X1 u2_u5_u4_U68 (.A2( u2_u5_u4_n101 ) , .A1( u2_u5_u4_n103 ) , .ZN( u2_u5_u4_n147 ) );
  NAND2_X1 u2_u5_u4_U69 (.A2( u2_u5_u4_n104 ) , .ZN( u2_u5_u4_n113 ) , .A1( u2_u5_u4_n99 ) );
  AOI21_X1 u2_u5_u4_U7 (.ZN( u2_u5_u4_n108 ) , .B2( u2_u5_u4_n134 ) , .B1( u2_u5_u4_n155 ) , .A( u2_u5_u4_n156 ) );
  NOR2_X1 u2_u5_u4_U70 (.A2( u2_u5_X_28 ) , .ZN( u2_u5_u4_n150 ) , .A1( u2_u5_u4_n168 ) );
  NOR2_X1 u2_u5_u4_U71 (.A2( u2_u5_X_29 ) , .ZN( u2_u5_u4_n152 ) , .A1( u2_u5_u4_n169 ) );
  NOR2_X1 u2_u5_u4_U72 (.A2( u2_u5_X_30 ) , .ZN( u2_u5_u4_n105 ) , .A1( u2_u5_u4_n176 ) );
  NOR2_X1 u2_u5_u4_U73 (.A2( u2_u5_X_26 ) , .ZN( u2_u5_u4_n100 ) , .A1( u2_u5_u4_n177 ) );
  NOR2_X1 u2_u5_u4_U74 (.A2( u2_u5_X_28 ) , .A1( u2_u5_X_29 ) , .ZN( u2_u5_u4_n128 ) );
  NOR2_X1 u2_u5_u4_U75 (.A2( u2_u5_X_27 ) , .A1( u2_u5_X_30 ) , .ZN( u2_u5_u4_n102 ) );
  NOR2_X1 u2_u5_u4_U76 (.A2( u2_u5_X_25 ) , .A1( u2_u5_X_26 ) , .ZN( u2_u5_u4_n98 ) );
  AND2_X1 u2_u5_u4_U77 (.A2( u2_u5_X_25 ) , .A1( u2_u5_X_26 ) , .ZN( u2_u5_u4_n104 ) );
  AND2_X1 u2_u5_u4_U78 (.A1( u2_u5_X_30 ) , .A2( u2_u5_u4_n176 ) , .ZN( u2_u5_u4_n99 ) );
  AND2_X1 u2_u5_u4_U79 (.A1( u2_u5_X_26 ) , .ZN( u2_u5_u4_n101 ) , .A2( u2_u5_u4_n177 ) );
  AOI21_X1 u2_u5_u4_U8 (.ZN( u2_u5_u4_n109 ) , .A( u2_u5_u4_n153 ) , .B1( u2_u5_u4_n159 ) , .B2( u2_u5_u4_n184 ) );
  AND2_X1 u2_u5_u4_U80 (.A1( u2_u5_X_27 ) , .A2( u2_u5_X_30 ) , .ZN( u2_u5_u4_n103 ) );
  INV_X1 u2_u5_u4_U81 (.A( u2_u5_X_28 ) , .ZN( u2_u5_u4_n169 ) );
  INV_X1 u2_u5_u4_U82 (.A( u2_u5_X_29 ) , .ZN( u2_u5_u4_n168 ) );
  INV_X1 u2_u5_u4_U83 (.A( u2_u5_X_25 ) , .ZN( u2_u5_u4_n177 ) );
  INV_X1 u2_u5_u4_U84 (.A( u2_u5_X_27 ) , .ZN( u2_u5_u4_n176 ) );
  NAND4_X1 u2_u5_u4_U85 (.ZN( u2_out5_25 ) , .A4( u2_u5_u4_n139 ) , .A3( u2_u5_u4_n140 ) , .A2( u2_u5_u4_n141 ) , .A1( u2_u5_u4_n142 ) );
  OAI21_X1 u2_u5_u4_U86 (.A( u2_u5_u4_n128 ) , .B2( u2_u5_u4_n129 ) , .B1( u2_u5_u4_n130 ) , .ZN( u2_u5_u4_n142 ) );
  OAI21_X1 u2_u5_u4_U87 (.B2( u2_u5_u4_n131 ) , .ZN( u2_u5_u4_n141 ) , .A( u2_u5_u4_n175 ) , .B1( u2_u5_u4_n183 ) );
  NAND4_X1 u2_u5_u4_U88 (.ZN( u2_out5_14 ) , .A4( u2_u5_u4_n124 ) , .A3( u2_u5_u4_n125 ) , .A2( u2_u5_u4_n126 ) , .A1( u2_u5_u4_n127 ) );
  AOI22_X1 u2_u5_u4_U89 (.B2( u2_u5_u4_n117 ) , .ZN( u2_u5_u4_n126 ) , .A1( u2_u5_u4_n129 ) , .B1( u2_u5_u4_n152 ) , .A2( u2_u5_u4_n175 ) );
  AOI211_X1 u2_u5_u4_U9 (.B( u2_u5_u4_n136 ) , .A( u2_u5_u4_n137 ) , .C2( u2_u5_u4_n138 ) , .ZN( u2_u5_u4_n139 ) , .C1( u2_u5_u4_n182 ) );
  AOI22_X1 u2_u5_u4_U90 (.ZN( u2_u5_u4_n125 ) , .B2( u2_u5_u4_n131 ) , .A2( u2_u5_u4_n132 ) , .B1( u2_u5_u4_n138 ) , .A1( u2_u5_u4_n178 ) );
  NAND4_X1 u2_u5_u4_U91 (.ZN( u2_out5_8 ) , .A4( u2_u5_u4_n110 ) , .A3( u2_u5_u4_n111 ) , .A2( u2_u5_u4_n112 ) , .A1( u2_u5_u4_n186 ) );
  NAND2_X1 u2_u5_u4_U92 (.ZN( u2_u5_u4_n112 ) , .A2( u2_u5_u4_n130 ) , .A1( u2_u5_u4_n150 ) );
  AOI22_X1 u2_u5_u4_U93 (.ZN( u2_u5_u4_n111 ) , .B2( u2_u5_u4_n132 ) , .A1( u2_u5_u4_n152 ) , .B1( u2_u5_u4_n178 ) , .A2( u2_u5_u4_n97 ) );
  AOI22_X1 u2_u5_u4_U94 (.B2( u2_u5_u4_n149 ) , .B1( u2_u5_u4_n150 ) , .A2( u2_u5_u4_n151 ) , .A1( u2_u5_u4_n152 ) , .ZN( u2_u5_u4_n167 ) );
  NOR4_X1 u2_u5_u4_U95 (.A4( u2_u5_u4_n162 ) , .A3( u2_u5_u4_n163 ) , .A2( u2_u5_u4_n164 ) , .A1( u2_u5_u4_n165 ) , .ZN( u2_u5_u4_n166 ) );
  NAND3_X1 u2_u5_u4_U96 (.ZN( u2_out5_3 ) , .A3( u2_u5_u4_n166 ) , .A1( u2_u5_u4_n167 ) , .A2( u2_u5_u4_n186 ) );
  NAND3_X1 u2_u5_u4_U97 (.A3( u2_u5_u4_n146 ) , .A2( u2_u5_u4_n147 ) , .A1( u2_u5_u4_n148 ) , .ZN( u2_u5_u4_n149 ) );
  NAND3_X1 u2_u5_u4_U98 (.A3( u2_u5_u4_n143 ) , .A2( u2_u5_u4_n144 ) , .A1( u2_u5_u4_n145 ) , .ZN( u2_u5_u4_n151 ) );
  NAND3_X1 u2_u5_u4_U99 (.A3( u2_u5_u4_n121 ) , .ZN( u2_u5_u4_n122 ) , .A2( u2_u5_u4_n144 ) , .A1( u2_u5_u4_n154 ) );
  INV_X1 u2_u5_u5_U10 (.A( u2_u5_u5_n121 ) , .ZN( u2_u5_u5_n177 ) );
  NOR3_X1 u2_u5_u5_U100 (.A3( u2_u5_u5_n141 ) , .A1( u2_u5_u5_n142 ) , .ZN( u2_u5_u5_n143 ) , .A2( u2_u5_u5_n191 ) );
  NAND4_X1 u2_u5_u5_U101 (.ZN( u2_out5_4 ) , .A4( u2_u5_u5_n112 ) , .A2( u2_u5_u5_n113 ) , .A1( u2_u5_u5_n114 ) , .A3( u2_u5_u5_n195 ) );
  AOI211_X1 u2_u5_u5_U102 (.A( u2_u5_u5_n110 ) , .C1( u2_u5_u5_n111 ) , .ZN( u2_u5_u5_n112 ) , .B( u2_u5_u5_n118 ) , .C2( u2_u5_u5_n177 ) );
  AOI222_X1 u2_u5_u5_U103 (.ZN( u2_u5_u5_n113 ) , .A1( u2_u5_u5_n131 ) , .C1( u2_u5_u5_n148 ) , .B2( u2_u5_u5_n174 ) , .C2( u2_u5_u5_n178 ) , .A2( u2_u5_u5_n179 ) , .B1( u2_u5_u5_n99 ) );
  NAND3_X1 u2_u5_u5_U104 (.A2( u2_u5_u5_n154 ) , .A3( u2_u5_u5_n158 ) , .A1( u2_u5_u5_n161 ) , .ZN( u2_u5_u5_n99 ) );
  NOR2_X1 u2_u5_u5_U11 (.ZN( u2_u5_u5_n160 ) , .A2( u2_u5_u5_n173 ) , .A1( u2_u5_u5_n177 ) );
  INV_X1 u2_u5_u5_U12 (.A( u2_u5_u5_n150 ) , .ZN( u2_u5_u5_n174 ) );
  AOI21_X1 u2_u5_u5_U13 (.A( u2_u5_u5_n160 ) , .B2( u2_u5_u5_n161 ) , .ZN( u2_u5_u5_n162 ) , .B1( u2_u5_u5_n192 ) );
  INV_X1 u2_u5_u5_U14 (.A( u2_u5_u5_n159 ) , .ZN( u2_u5_u5_n192 ) );
  AOI21_X1 u2_u5_u5_U15 (.A( u2_u5_u5_n156 ) , .B2( u2_u5_u5_n157 ) , .B1( u2_u5_u5_n158 ) , .ZN( u2_u5_u5_n163 ) );
  AOI21_X1 u2_u5_u5_U16 (.B2( u2_u5_u5_n139 ) , .B1( u2_u5_u5_n140 ) , .ZN( u2_u5_u5_n141 ) , .A( u2_u5_u5_n150 ) );
  OAI21_X1 u2_u5_u5_U17 (.A( u2_u5_u5_n133 ) , .B2( u2_u5_u5_n134 ) , .B1( u2_u5_u5_n135 ) , .ZN( u2_u5_u5_n142 ) );
  OAI21_X1 u2_u5_u5_U18 (.ZN( u2_u5_u5_n133 ) , .B2( u2_u5_u5_n147 ) , .A( u2_u5_u5_n173 ) , .B1( u2_u5_u5_n188 ) );
  NAND2_X1 u2_u5_u5_U19 (.A2( u2_u5_u5_n119 ) , .A1( u2_u5_u5_n123 ) , .ZN( u2_u5_u5_n137 ) );
  INV_X1 u2_u5_u5_U20 (.A( u2_u5_u5_n155 ) , .ZN( u2_u5_u5_n194 ) );
  NAND2_X1 u2_u5_u5_U21 (.A1( u2_u5_u5_n121 ) , .ZN( u2_u5_u5_n132 ) , .A2( u2_u5_u5_n172 ) );
  NAND2_X1 u2_u5_u5_U22 (.A2( u2_u5_u5_n122 ) , .ZN( u2_u5_u5_n136 ) , .A1( u2_u5_u5_n154 ) );
  NAND2_X1 u2_u5_u5_U23 (.A2( u2_u5_u5_n119 ) , .A1( u2_u5_u5_n120 ) , .ZN( u2_u5_u5_n159 ) );
  INV_X1 u2_u5_u5_U24 (.A( u2_u5_u5_n156 ) , .ZN( u2_u5_u5_n175 ) );
  INV_X1 u2_u5_u5_U25 (.A( u2_u5_u5_n158 ) , .ZN( u2_u5_u5_n188 ) );
  INV_X1 u2_u5_u5_U26 (.A( u2_u5_u5_n152 ) , .ZN( u2_u5_u5_n179 ) );
  INV_X1 u2_u5_u5_U27 (.A( u2_u5_u5_n140 ) , .ZN( u2_u5_u5_n182 ) );
  INV_X1 u2_u5_u5_U28 (.A( u2_u5_u5_n151 ) , .ZN( u2_u5_u5_n183 ) );
  INV_X1 u2_u5_u5_U29 (.A( u2_u5_u5_n123 ) , .ZN( u2_u5_u5_n185 ) );
  NOR2_X1 u2_u5_u5_U3 (.ZN( u2_u5_u5_n134 ) , .A1( u2_u5_u5_n183 ) , .A2( u2_u5_u5_n190 ) );
  INV_X1 u2_u5_u5_U30 (.A( u2_u5_u5_n161 ) , .ZN( u2_u5_u5_n184 ) );
  INV_X1 u2_u5_u5_U31 (.A( u2_u5_u5_n139 ) , .ZN( u2_u5_u5_n189 ) );
  INV_X1 u2_u5_u5_U32 (.A( u2_u5_u5_n157 ) , .ZN( u2_u5_u5_n190 ) );
  INV_X1 u2_u5_u5_U33 (.A( u2_u5_u5_n120 ) , .ZN( u2_u5_u5_n193 ) );
  NAND2_X1 u2_u5_u5_U34 (.ZN( u2_u5_u5_n111 ) , .A1( u2_u5_u5_n140 ) , .A2( u2_u5_u5_n155 ) );
  NOR2_X1 u2_u5_u5_U35 (.ZN( u2_u5_u5_n100 ) , .A1( u2_u5_u5_n170 ) , .A2( u2_u5_u5_n180 ) );
  INV_X1 u2_u5_u5_U36 (.A( u2_u5_u5_n117 ) , .ZN( u2_u5_u5_n196 ) );
  OAI221_X1 u2_u5_u5_U37 (.A( u2_u5_u5_n116 ) , .ZN( u2_u5_u5_n117 ) , .B2( u2_u5_u5_n119 ) , .C1( u2_u5_u5_n153 ) , .C2( u2_u5_u5_n158 ) , .B1( u2_u5_u5_n172 ) );
  AOI222_X1 u2_u5_u5_U38 (.ZN( u2_u5_u5_n116 ) , .B2( u2_u5_u5_n145 ) , .C1( u2_u5_u5_n148 ) , .A2( u2_u5_u5_n174 ) , .C2( u2_u5_u5_n177 ) , .B1( u2_u5_u5_n187 ) , .A1( u2_u5_u5_n193 ) );
  INV_X1 u2_u5_u5_U39 (.A( u2_u5_u5_n115 ) , .ZN( u2_u5_u5_n187 ) );
  INV_X1 u2_u5_u5_U4 (.A( u2_u5_u5_n138 ) , .ZN( u2_u5_u5_n191 ) );
  AOI22_X1 u2_u5_u5_U40 (.B2( u2_u5_u5_n131 ) , .A2( u2_u5_u5_n146 ) , .ZN( u2_u5_u5_n169 ) , .B1( u2_u5_u5_n174 ) , .A1( u2_u5_u5_n185 ) );
  NOR2_X1 u2_u5_u5_U41 (.A1( u2_u5_u5_n146 ) , .ZN( u2_u5_u5_n150 ) , .A2( u2_u5_u5_n173 ) );
  AOI21_X1 u2_u5_u5_U42 (.A( u2_u5_u5_n118 ) , .B2( u2_u5_u5_n145 ) , .ZN( u2_u5_u5_n168 ) , .B1( u2_u5_u5_n186 ) );
  INV_X1 u2_u5_u5_U43 (.A( u2_u5_u5_n122 ) , .ZN( u2_u5_u5_n186 ) );
  NOR2_X1 u2_u5_u5_U44 (.A1( u2_u5_u5_n146 ) , .ZN( u2_u5_u5_n152 ) , .A2( u2_u5_u5_n176 ) );
  NOR2_X1 u2_u5_u5_U45 (.A1( u2_u5_u5_n115 ) , .ZN( u2_u5_u5_n118 ) , .A2( u2_u5_u5_n153 ) );
  NOR2_X1 u2_u5_u5_U46 (.A2( u2_u5_u5_n145 ) , .ZN( u2_u5_u5_n156 ) , .A1( u2_u5_u5_n174 ) );
  NOR2_X1 u2_u5_u5_U47 (.ZN( u2_u5_u5_n121 ) , .A2( u2_u5_u5_n145 ) , .A1( u2_u5_u5_n176 ) );
  AOI22_X1 u2_u5_u5_U48 (.ZN( u2_u5_u5_n114 ) , .A2( u2_u5_u5_n137 ) , .A1( u2_u5_u5_n145 ) , .B2( u2_u5_u5_n175 ) , .B1( u2_u5_u5_n193 ) );
  OAI211_X1 u2_u5_u5_U49 (.B( u2_u5_u5_n124 ) , .A( u2_u5_u5_n125 ) , .C2( u2_u5_u5_n126 ) , .C1( u2_u5_u5_n127 ) , .ZN( u2_u5_u5_n128 ) );
  OAI21_X1 u2_u5_u5_U5 (.B2( u2_u5_u5_n136 ) , .B1( u2_u5_u5_n137 ) , .ZN( u2_u5_u5_n138 ) , .A( u2_u5_u5_n177 ) );
  NOR3_X1 u2_u5_u5_U50 (.ZN( u2_u5_u5_n127 ) , .A1( u2_u5_u5_n136 ) , .A3( u2_u5_u5_n148 ) , .A2( u2_u5_u5_n182 ) );
  OAI21_X1 u2_u5_u5_U51 (.ZN( u2_u5_u5_n124 ) , .A( u2_u5_u5_n177 ) , .B2( u2_u5_u5_n183 ) , .B1( u2_u5_u5_n189 ) );
  OAI21_X1 u2_u5_u5_U52 (.ZN( u2_u5_u5_n125 ) , .A( u2_u5_u5_n174 ) , .B2( u2_u5_u5_n185 ) , .B1( u2_u5_u5_n190 ) );
  AOI21_X1 u2_u5_u5_U53 (.A( u2_u5_u5_n153 ) , .B2( u2_u5_u5_n154 ) , .B1( u2_u5_u5_n155 ) , .ZN( u2_u5_u5_n164 ) );
  AOI21_X1 u2_u5_u5_U54 (.ZN( u2_u5_u5_n110 ) , .B1( u2_u5_u5_n122 ) , .B2( u2_u5_u5_n139 ) , .A( u2_u5_u5_n153 ) );
  INV_X1 u2_u5_u5_U55 (.A( u2_u5_u5_n153 ) , .ZN( u2_u5_u5_n176 ) );
  INV_X1 u2_u5_u5_U56 (.A( u2_u5_u5_n126 ) , .ZN( u2_u5_u5_n173 ) );
  AND2_X1 u2_u5_u5_U57 (.A2( u2_u5_u5_n104 ) , .A1( u2_u5_u5_n107 ) , .ZN( u2_u5_u5_n147 ) );
  AND2_X1 u2_u5_u5_U58 (.A2( u2_u5_u5_n104 ) , .A1( u2_u5_u5_n108 ) , .ZN( u2_u5_u5_n148 ) );
  NAND2_X1 u2_u5_u5_U59 (.A1( u2_u5_u5_n105 ) , .A2( u2_u5_u5_n106 ) , .ZN( u2_u5_u5_n158 ) );
  INV_X1 u2_u5_u5_U6 (.A( u2_u5_u5_n135 ) , .ZN( u2_u5_u5_n178 ) );
  NAND2_X1 u2_u5_u5_U60 (.A2( u2_u5_u5_n108 ) , .A1( u2_u5_u5_n109 ) , .ZN( u2_u5_u5_n139 ) );
  NAND2_X1 u2_u5_u5_U61 (.A1( u2_u5_u5_n106 ) , .A2( u2_u5_u5_n108 ) , .ZN( u2_u5_u5_n119 ) );
  NAND2_X1 u2_u5_u5_U62 (.A2( u2_u5_u5_n103 ) , .A1( u2_u5_u5_n105 ) , .ZN( u2_u5_u5_n140 ) );
  NAND2_X1 u2_u5_u5_U63 (.A2( u2_u5_u5_n104 ) , .A1( u2_u5_u5_n105 ) , .ZN( u2_u5_u5_n155 ) );
  NAND2_X1 u2_u5_u5_U64 (.A2( u2_u5_u5_n106 ) , .A1( u2_u5_u5_n107 ) , .ZN( u2_u5_u5_n122 ) );
  NAND2_X1 u2_u5_u5_U65 (.A2( u2_u5_u5_n100 ) , .A1( u2_u5_u5_n106 ) , .ZN( u2_u5_u5_n115 ) );
  NAND2_X1 u2_u5_u5_U66 (.A2( u2_u5_u5_n100 ) , .A1( u2_u5_u5_n103 ) , .ZN( u2_u5_u5_n161 ) );
  NAND2_X1 u2_u5_u5_U67 (.A1( u2_u5_u5_n105 ) , .A2( u2_u5_u5_n109 ) , .ZN( u2_u5_u5_n154 ) );
  INV_X1 u2_u5_u5_U68 (.A( u2_u5_u5_n146 ) , .ZN( u2_u5_u5_n172 ) );
  NAND2_X1 u2_u5_u5_U69 (.A1( u2_u5_u5_n103 ) , .A2( u2_u5_u5_n108 ) , .ZN( u2_u5_u5_n123 ) );
  OAI22_X1 u2_u5_u5_U7 (.B2( u2_u5_u5_n149 ) , .B1( u2_u5_u5_n150 ) , .A2( u2_u5_u5_n151 ) , .A1( u2_u5_u5_n152 ) , .ZN( u2_u5_u5_n165 ) );
  NAND2_X1 u2_u5_u5_U70 (.A2( u2_u5_u5_n103 ) , .A1( u2_u5_u5_n107 ) , .ZN( u2_u5_u5_n151 ) );
  NAND2_X1 u2_u5_u5_U71 (.A2( u2_u5_u5_n107 ) , .A1( u2_u5_u5_n109 ) , .ZN( u2_u5_u5_n120 ) );
  NAND2_X1 u2_u5_u5_U72 (.A2( u2_u5_u5_n100 ) , .A1( u2_u5_u5_n109 ) , .ZN( u2_u5_u5_n157 ) );
  AND2_X1 u2_u5_u5_U73 (.A2( u2_u5_u5_n100 ) , .A1( u2_u5_u5_n104 ) , .ZN( u2_u5_u5_n131 ) );
  INV_X1 u2_u5_u5_U74 (.A( u2_u5_u5_n102 ) , .ZN( u2_u5_u5_n195 ) );
  OAI221_X1 u2_u5_u5_U75 (.A( u2_u5_u5_n101 ) , .ZN( u2_u5_u5_n102 ) , .C2( u2_u5_u5_n115 ) , .C1( u2_u5_u5_n126 ) , .B1( u2_u5_u5_n134 ) , .B2( u2_u5_u5_n160 ) );
  OAI21_X1 u2_u5_u5_U76 (.ZN( u2_u5_u5_n101 ) , .B1( u2_u5_u5_n137 ) , .A( u2_u5_u5_n146 ) , .B2( u2_u5_u5_n147 ) );
  NOR2_X1 u2_u5_u5_U77 (.A2( u2_u5_X_34 ) , .A1( u2_u5_X_35 ) , .ZN( u2_u5_u5_n145 ) );
  NOR2_X1 u2_u5_u5_U78 (.A2( u2_u5_X_34 ) , .ZN( u2_u5_u5_n146 ) , .A1( u2_u5_u5_n171 ) );
  NOR2_X1 u2_u5_u5_U79 (.A2( u2_u5_X_31 ) , .A1( u2_u5_X_32 ) , .ZN( u2_u5_u5_n103 ) );
  NOR3_X1 u2_u5_u5_U8 (.A2( u2_u5_u5_n147 ) , .A1( u2_u5_u5_n148 ) , .ZN( u2_u5_u5_n149 ) , .A3( u2_u5_u5_n194 ) );
  NOR2_X1 u2_u5_u5_U80 (.A2( u2_u5_X_36 ) , .ZN( u2_u5_u5_n105 ) , .A1( u2_u5_u5_n180 ) );
  NOR2_X1 u2_u5_u5_U81 (.A2( u2_u5_X_33 ) , .ZN( u2_u5_u5_n108 ) , .A1( u2_u5_u5_n170 ) );
  NOR2_X1 u2_u5_u5_U82 (.A2( u2_u5_X_33 ) , .A1( u2_u5_X_36 ) , .ZN( u2_u5_u5_n107 ) );
  NOR2_X1 u2_u5_u5_U83 (.A2( u2_u5_X_31 ) , .ZN( u2_u5_u5_n104 ) , .A1( u2_u5_u5_n181 ) );
  NAND2_X1 u2_u5_u5_U84 (.A2( u2_u5_X_34 ) , .A1( u2_u5_X_35 ) , .ZN( u2_u5_u5_n153 ) );
  NAND2_X1 u2_u5_u5_U85 (.A1( u2_u5_X_34 ) , .ZN( u2_u5_u5_n126 ) , .A2( u2_u5_u5_n171 ) );
  AND2_X1 u2_u5_u5_U86 (.A1( u2_u5_X_31 ) , .A2( u2_u5_X_32 ) , .ZN( u2_u5_u5_n106 ) );
  AND2_X1 u2_u5_u5_U87 (.A1( u2_u5_X_31 ) , .ZN( u2_u5_u5_n109 ) , .A2( u2_u5_u5_n181 ) );
  INV_X1 u2_u5_u5_U88 (.A( u2_u5_X_33 ) , .ZN( u2_u5_u5_n180 ) );
  INV_X1 u2_u5_u5_U89 (.A( u2_u5_X_35 ) , .ZN( u2_u5_u5_n171 ) );
  NOR2_X1 u2_u5_u5_U9 (.ZN( u2_u5_u5_n135 ) , .A1( u2_u5_u5_n173 ) , .A2( u2_u5_u5_n176 ) );
  INV_X1 u2_u5_u5_U90 (.A( u2_u5_X_36 ) , .ZN( u2_u5_u5_n170 ) );
  INV_X1 u2_u5_u5_U91 (.A( u2_u5_X_32 ) , .ZN( u2_u5_u5_n181 ) );
  NAND4_X1 u2_u5_u5_U92 (.ZN( u2_out5_29 ) , .A4( u2_u5_u5_n129 ) , .A3( u2_u5_u5_n130 ) , .A2( u2_u5_u5_n168 ) , .A1( u2_u5_u5_n196 ) );
  AOI221_X1 u2_u5_u5_U93 (.A( u2_u5_u5_n128 ) , .ZN( u2_u5_u5_n129 ) , .C2( u2_u5_u5_n132 ) , .B2( u2_u5_u5_n159 ) , .B1( u2_u5_u5_n176 ) , .C1( u2_u5_u5_n184 ) );
  AOI222_X1 u2_u5_u5_U94 (.ZN( u2_u5_u5_n130 ) , .A2( u2_u5_u5_n146 ) , .B1( u2_u5_u5_n147 ) , .C2( u2_u5_u5_n175 ) , .B2( u2_u5_u5_n179 ) , .A1( u2_u5_u5_n188 ) , .C1( u2_u5_u5_n194 ) );
  NAND4_X1 u2_u5_u5_U95 (.ZN( u2_out5_19 ) , .A4( u2_u5_u5_n166 ) , .A3( u2_u5_u5_n167 ) , .A2( u2_u5_u5_n168 ) , .A1( u2_u5_u5_n169 ) );
  AOI22_X1 u2_u5_u5_U96 (.B2( u2_u5_u5_n145 ) , .A2( u2_u5_u5_n146 ) , .ZN( u2_u5_u5_n167 ) , .B1( u2_u5_u5_n182 ) , .A1( u2_u5_u5_n189 ) );
  NOR4_X1 u2_u5_u5_U97 (.A4( u2_u5_u5_n162 ) , .A3( u2_u5_u5_n163 ) , .A2( u2_u5_u5_n164 ) , .A1( u2_u5_u5_n165 ) , .ZN( u2_u5_u5_n166 ) );
  NAND4_X1 u2_u5_u5_U98 (.ZN( u2_out5_11 ) , .A4( u2_u5_u5_n143 ) , .A3( u2_u5_u5_n144 ) , .A2( u2_u5_u5_n169 ) , .A1( u2_u5_u5_n196 ) );
  AOI22_X1 u2_u5_u5_U99 (.A2( u2_u5_u5_n132 ) , .ZN( u2_u5_u5_n144 ) , .B2( u2_u5_u5_n145 ) , .B1( u2_u5_u5_n184 ) , .A1( u2_u5_u5_n194 ) );
  OAI21_X1 u2_u5_u6_U10 (.A( u2_u5_u6_n159 ) , .B1( u2_u5_u6_n169 ) , .B2( u2_u5_u6_n173 ) , .ZN( u2_u5_u6_n90 ) );
  INV_X1 u2_u5_u6_U11 (.ZN( u2_u5_u6_n172 ) , .A( u2_u5_u6_n88 ) );
  AOI22_X1 u2_u5_u6_U12 (.A2( u2_u5_u6_n151 ) , .B2( u2_u5_u6_n161 ) , .A1( u2_u5_u6_n167 ) , .B1( u2_u5_u6_n170 ) , .ZN( u2_u5_u6_n89 ) );
  AOI21_X1 u2_u5_u6_U13 (.ZN( u2_u5_u6_n106 ) , .A( u2_u5_u6_n142 ) , .B2( u2_u5_u6_n159 ) , .B1( u2_u5_u6_n164 ) );
  INV_X1 u2_u5_u6_U14 (.A( u2_u5_u6_n155 ) , .ZN( u2_u5_u6_n161 ) );
  INV_X1 u2_u5_u6_U15 (.A( u2_u5_u6_n128 ) , .ZN( u2_u5_u6_n164 ) );
  NAND2_X1 u2_u5_u6_U16 (.ZN( u2_u5_u6_n110 ) , .A1( u2_u5_u6_n122 ) , .A2( u2_u5_u6_n129 ) );
  NAND2_X1 u2_u5_u6_U17 (.ZN( u2_u5_u6_n124 ) , .A2( u2_u5_u6_n146 ) , .A1( u2_u5_u6_n148 ) );
  INV_X1 u2_u5_u6_U18 (.A( u2_u5_u6_n132 ) , .ZN( u2_u5_u6_n171 ) );
  AND2_X1 u2_u5_u6_U19 (.A1( u2_u5_u6_n100 ) , .ZN( u2_u5_u6_n130 ) , .A2( u2_u5_u6_n147 ) );
  INV_X1 u2_u5_u6_U20 (.A( u2_u5_u6_n127 ) , .ZN( u2_u5_u6_n173 ) );
  INV_X1 u2_u5_u6_U21 (.A( u2_u5_u6_n121 ) , .ZN( u2_u5_u6_n167 ) );
  INV_X1 u2_u5_u6_U22 (.A( u2_u5_u6_n100 ) , .ZN( u2_u5_u6_n169 ) );
  INV_X1 u2_u5_u6_U23 (.A( u2_u5_u6_n123 ) , .ZN( u2_u5_u6_n170 ) );
  INV_X1 u2_u5_u6_U24 (.A( u2_u5_u6_n113 ) , .ZN( u2_u5_u6_n168 ) );
  AND2_X1 u2_u5_u6_U25 (.A1( u2_u5_u6_n107 ) , .A2( u2_u5_u6_n119 ) , .ZN( u2_u5_u6_n133 ) );
  AND2_X1 u2_u5_u6_U26 (.A2( u2_u5_u6_n121 ) , .A1( u2_u5_u6_n122 ) , .ZN( u2_u5_u6_n131 ) );
  AND3_X1 u2_u5_u6_U27 (.ZN( u2_u5_u6_n120 ) , .A2( u2_u5_u6_n127 ) , .A1( u2_u5_u6_n132 ) , .A3( u2_u5_u6_n145 ) );
  INV_X1 u2_u5_u6_U28 (.A( u2_u5_u6_n146 ) , .ZN( u2_u5_u6_n163 ) );
  AOI222_X1 u2_u5_u6_U29 (.ZN( u2_u5_u6_n114 ) , .A1( u2_u5_u6_n118 ) , .A2( u2_u5_u6_n126 ) , .B2( u2_u5_u6_n151 ) , .C2( u2_u5_u6_n159 ) , .C1( u2_u5_u6_n168 ) , .B1( u2_u5_u6_n169 ) );
  INV_X1 u2_u5_u6_U3 (.A( u2_u5_u6_n110 ) , .ZN( u2_u5_u6_n166 ) );
  NOR2_X1 u2_u5_u6_U30 (.A1( u2_u5_u6_n162 ) , .A2( u2_u5_u6_n165 ) , .ZN( u2_u5_u6_n98 ) );
  NAND2_X1 u2_u5_u6_U31 (.A1( u2_u5_u6_n144 ) , .ZN( u2_u5_u6_n151 ) , .A2( u2_u5_u6_n158 ) );
  NAND2_X1 u2_u5_u6_U32 (.ZN( u2_u5_u6_n132 ) , .A1( u2_u5_u6_n91 ) , .A2( u2_u5_u6_n97 ) );
  NOR2_X1 u2_u5_u6_U33 (.A2( u2_u5_u6_n126 ) , .ZN( u2_u5_u6_n155 ) , .A1( u2_u5_u6_n160 ) );
  NAND2_X1 u2_u5_u6_U34 (.ZN( u2_u5_u6_n146 ) , .A2( u2_u5_u6_n94 ) , .A1( u2_u5_u6_n99 ) );
  AOI21_X1 u2_u5_u6_U35 (.A( u2_u5_u6_n144 ) , .B2( u2_u5_u6_n145 ) , .B1( u2_u5_u6_n146 ) , .ZN( u2_u5_u6_n150 ) );
  INV_X1 u2_u5_u6_U36 (.A( u2_u5_u6_n111 ) , .ZN( u2_u5_u6_n158 ) );
  NAND2_X1 u2_u5_u6_U37 (.ZN( u2_u5_u6_n127 ) , .A1( u2_u5_u6_n91 ) , .A2( u2_u5_u6_n92 ) );
  NAND2_X1 u2_u5_u6_U38 (.ZN( u2_u5_u6_n129 ) , .A2( u2_u5_u6_n95 ) , .A1( u2_u5_u6_n96 ) );
  INV_X1 u2_u5_u6_U39 (.A( u2_u5_u6_n144 ) , .ZN( u2_u5_u6_n159 ) );
  INV_X1 u2_u5_u6_U4 (.A( u2_u5_u6_n142 ) , .ZN( u2_u5_u6_n174 ) );
  NAND2_X1 u2_u5_u6_U40 (.ZN( u2_u5_u6_n145 ) , .A2( u2_u5_u6_n97 ) , .A1( u2_u5_u6_n98 ) );
  NAND2_X1 u2_u5_u6_U41 (.ZN( u2_u5_u6_n148 ) , .A2( u2_u5_u6_n92 ) , .A1( u2_u5_u6_n94 ) );
  NAND2_X1 u2_u5_u6_U42 (.ZN( u2_u5_u6_n108 ) , .A2( u2_u5_u6_n139 ) , .A1( u2_u5_u6_n144 ) );
  NAND2_X1 u2_u5_u6_U43 (.ZN( u2_u5_u6_n121 ) , .A2( u2_u5_u6_n95 ) , .A1( u2_u5_u6_n97 ) );
  NAND2_X1 u2_u5_u6_U44 (.ZN( u2_u5_u6_n107 ) , .A2( u2_u5_u6_n92 ) , .A1( u2_u5_u6_n95 ) );
  AND2_X1 u2_u5_u6_U45 (.ZN( u2_u5_u6_n118 ) , .A2( u2_u5_u6_n91 ) , .A1( u2_u5_u6_n99 ) );
  AOI22_X1 u2_u5_u6_U46 (.B2( u2_u5_u6_n110 ) , .B1( u2_u5_u6_n111 ) , .A1( u2_u5_u6_n112 ) , .ZN( u2_u5_u6_n115 ) , .A2( u2_u5_u6_n161 ) );
  NAND4_X1 u2_u5_u6_U47 (.A3( u2_u5_u6_n109 ) , .ZN( u2_u5_u6_n112 ) , .A4( u2_u5_u6_n132 ) , .A2( u2_u5_u6_n147 ) , .A1( u2_u5_u6_n166 ) );
  NOR2_X1 u2_u5_u6_U48 (.ZN( u2_u5_u6_n109 ) , .A1( u2_u5_u6_n170 ) , .A2( u2_u5_u6_n173 ) );
  NAND2_X1 u2_u5_u6_U49 (.ZN( u2_u5_u6_n147 ) , .A2( u2_u5_u6_n98 ) , .A1( u2_u5_u6_n99 ) );
  NAND2_X1 u2_u5_u6_U5 (.A2( u2_u5_u6_n143 ) , .ZN( u2_u5_u6_n152 ) , .A1( u2_u5_u6_n166 ) );
  NAND2_X1 u2_u5_u6_U50 (.ZN( u2_u5_u6_n128 ) , .A1( u2_u5_u6_n94 ) , .A2( u2_u5_u6_n96 ) );
  AOI211_X1 u2_u5_u6_U51 (.B( u2_u5_u6_n134 ) , .A( u2_u5_u6_n135 ) , .C1( u2_u5_u6_n136 ) , .ZN( u2_u5_u6_n137 ) , .C2( u2_u5_u6_n151 ) );
  AOI21_X1 u2_u5_u6_U52 (.B2( u2_u5_u6_n132 ) , .B1( u2_u5_u6_n133 ) , .ZN( u2_u5_u6_n134 ) , .A( u2_u5_u6_n158 ) );
  AOI21_X1 u2_u5_u6_U53 (.B1( u2_u5_u6_n131 ) , .ZN( u2_u5_u6_n135 ) , .A( u2_u5_u6_n144 ) , .B2( u2_u5_u6_n146 ) );
  NAND4_X1 u2_u5_u6_U54 (.A4( u2_u5_u6_n127 ) , .A3( u2_u5_u6_n128 ) , .A2( u2_u5_u6_n129 ) , .A1( u2_u5_u6_n130 ) , .ZN( u2_u5_u6_n136 ) );
  NAND2_X1 u2_u5_u6_U55 (.ZN( u2_u5_u6_n119 ) , .A2( u2_u5_u6_n95 ) , .A1( u2_u5_u6_n99 ) );
  NAND2_X1 u2_u5_u6_U56 (.ZN( u2_u5_u6_n123 ) , .A2( u2_u5_u6_n91 ) , .A1( u2_u5_u6_n96 ) );
  NAND2_X1 u2_u5_u6_U57 (.ZN( u2_u5_u6_n100 ) , .A2( u2_u5_u6_n92 ) , .A1( u2_u5_u6_n98 ) );
  NAND2_X1 u2_u5_u6_U58 (.ZN( u2_u5_u6_n122 ) , .A1( u2_u5_u6_n94 ) , .A2( u2_u5_u6_n97 ) );
  INV_X1 u2_u5_u6_U59 (.A( u2_u5_u6_n139 ) , .ZN( u2_u5_u6_n160 ) );
  AOI22_X1 u2_u5_u6_U6 (.B2( u2_u5_u6_n101 ) , .A1( u2_u5_u6_n102 ) , .ZN( u2_u5_u6_n103 ) , .B1( u2_u5_u6_n160 ) , .A2( u2_u5_u6_n161 ) );
  NAND2_X1 u2_u5_u6_U60 (.ZN( u2_u5_u6_n113 ) , .A1( u2_u5_u6_n96 ) , .A2( u2_u5_u6_n98 ) );
  NOR2_X1 u2_u5_u6_U61 (.A2( u2_u5_X_40 ) , .A1( u2_u5_X_41 ) , .ZN( u2_u5_u6_n126 ) );
  NOR2_X1 u2_u5_u6_U62 (.A2( u2_u5_X_39 ) , .A1( u2_u5_X_42 ) , .ZN( u2_u5_u6_n92 ) );
  NOR2_X1 u2_u5_u6_U63 (.A2( u2_u5_X_39 ) , .A1( u2_u5_u6_n156 ) , .ZN( u2_u5_u6_n97 ) );
  NOR2_X1 u2_u5_u6_U64 (.A2( u2_u5_X_38 ) , .A1( u2_u5_u6_n165 ) , .ZN( u2_u5_u6_n95 ) );
  NOR2_X1 u2_u5_u6_U65 (.A2( u2_u5_X_41 ) , .ZN( u2_u5_u6_n111 ) , .A1( u2_u5_u6_n157 ) );
  NOR2_X1 u2_u5_u6_U66 (.A2( u2_u5_X_37 ) , .A1( u2_u5_u6_n162 ) , .ZN( u2_u5_u6_n94 ) );
  NOR2_X1 u2_u5_u6_U67 (.A2( u2_u5_X_37 ) , .A1( u2_u5_X_38 ) , .ZN( u2_u5_u6_n91 ) );
  NAND2_X1 u2_u5_u6_U68 (.A1( u2_u5_X_41 ) , .ZN( u2_u5_u6_n144 ) , .A2( u2_u5_u6_n157 ) );
  NAND2_X1 u2_u5_u6_U69 (.A2( u2_u5_X_40 ) , .A1( u2_u5_X_41 ) , .ZN( u2_u5_u6_n139 ) );
  NOR2_X1 u2_u5_u6_U7 (.A1( u2_u5_u6_n118 ) , .ZN( u2_u5_u6_n143 ) , .A2( u2_u5_u6_n168 ) );
  AND2_X1 u2_u5_u6_U70 (.A1( u2_u5_X_39 ) , .A2( u2_u5_u6_n156 ) , .ZN( u2_u5_u6_n96 ) );
  AND2_X1 u2_u5_u6_U71 (.A1( u2_u5_X_39 ) , .A2( u2_u5_X_42 ) , .ZN( u2_u5_u6_n99 ) );
  INV_X1 u2_u5_u6_U72 (.A( u2_u5_X_40 ) , .ZN( u2_u5_u6_n157 ) );
  INV_X1 u2_u5_u6_U73 (.A( u2_u5_X_37 ) , .ZN( u2_u5_u6_n165 ) );
  INV_X1 u2_u5_u6_U74 (.A( u2_u5_X_38 ) , .ZN( u2_u5_u6_n162 ) );
  INV_X1 u2_u5_u6_U75 (.A( u2_u5_X_42 ) , .ZN( u2_u5_u6_n156 ) );
  NAND4_X1 u2_u5_u6_U76 (.ZN( u2_out5_32 ) , .A4( u2_u5_u6_n103 ) , .A3( u2_u5_u6_n104 ) , .A2( u2_u5_u6_n105 ) , .A1( u2_u5_u6_n106 ) );
  AOI22_X1 u2_u5_u6_U77 (.ZN( u2_u5_u6_n105 ) , .A2( u2_u5_u6_n108 ) , .A1( u2_u5_u6_n118 ) , .B2( u2_u5_u6_n126 ) , .B1( u2_u5_u6_n171 ) );
  AOI22_X1 u2_u5_u6_U78 (.ZN( u2_u5_u6_n104 ) , .A1( u2_u5_u6_n111 ) , .B1( u2_u5_u6_n124 ) , .B2( u2_u5_u6_n151 ) , .A2( u2_u5_u6_n93 ) );
  NAND4_X1 u2_u5_u6_U79 (.ZN( u2_out5_12 ) , .A4( u2_u5_u6_n114 ) , .A3( u2_u5_u6_n115 ) , .A2( u2_u5_u6_n116 ) , .A1( u2_u5_u6_n117 ) );
  AOI21_X1 u2_u5_u6_U8 (.B1( u2_u5_u6_n107 ) , .B2( u2_u5_u6_n132 ) , .A( u2_u5_u6_n158 ) , .ZN( u2_u5_u6_n88 ) );
  OAI22_X1 u2_u5_u6_U80 (.B2( u2_u5_u6_n111 ) , .ZN( u2_u5_u6_n116 ) , .B1( u2_u5_u6_n126 ) , .A2( u2_u5_u6_n164 ) , .A1( u2_u5_u6_n167 ) );
  OAI21_X1 u2_u5_u6_U81 (.A( u2_u5_u6_n108 ) , .ZN( u2_u5_u6_n117 ) , .B2( u2_u5_u6_n141 ) , .B1( u2_u5_u6_n163 ) );
  OAI211_X1 u2_u5_u6_U82 (.ZN( u2_out5_22 ) , .B( u2_u5_u6_n137 ) , .A( u2_u5_u6_n138 ) , .C2( u2_u5_u6_n139 ) , .C1( u2_u5_u6_n140 ) );
  AOI22_X1 u2_u5_u6_U83 (.B1( u2_u5_u6_n124 ) , .A2( u2_u5_u6_n125 ) , .A1( u2_u5_u6_n126 ) , .ZN( u2_u5_u6_n138 ) , .B2( u2_u5_u6_n161 ) );
  AND4_X1 u2_u5_u6_U84 (.A3( u2_u5_u6_n119 ) , .A1( u2_u5_u6_n120 ) , .A4( u2_u5_u6_n129 ) , .ZN( u2_u5_u6_n140 ) , .A2( u2_u5_u6_n143 ) );
  OAI211_X1 u2_u5_u6_U85 (.ZN( u2_out5_7 ) , .B( u2_u5_u6_n153 ) , .C2( u2_u5_u6_n154 ) , .C1( u2_u5_u6_n155 ) , .A( u2_u5_u6_n174 ) );
  NOR3_X1 u2_u5_u6_U86 (.A1( u2_u5_u6_n141 ) , .ZN( u2_u5_u6_n154 ) , .A3( u2_u5_u6_n164 ) , .A2( u2_u5_u6_n171 ) );
  AOI211_X1 u2_u5_u6_U87 (.B( u2_u5_u6_n149 ) , .A( u2_u5_u6_n150 ) , .C2( u2_u5_u6_n151 ) , .C1( u2_u5_u6_n152 ) , .ZN( u2_u5_u6_n153 ) );
  NAND3_X1 u2_u5_u6_U88 (.A2( u2_u5_u6_n123 ) , .ZN( u2_u5_u6_n125 ) , .A1( u2_u5_u6_n130 ) , .A3( u2_u5_u6_n131 ) );
  NAND3_X1 u2_u5_u6_U89 (.A3( u2_u5_u6_n133 ) , .ZN( u2_u5_u6_n141 ) , .A1( u2_u5_u6_n145 ) , .A2( u2_u5_u6_n148 ) );
  AOI21_X1 u2_u5_u6_U9 (.B2( u2_u5_u6_n147 ) , .B1( u2_u5_u6_n148 ) , .ZN( u2_u5_u6_n149 ) , .A( u2_u5_u6_n158 ) );
  NAND3_X1 u2_u5_u6_U90 (.ZN( u2_u5_u6_n101 ) , .A3( u2_u5_u6_n107 ) , .A2( u2_u5_u6_n121 ) , .A1( u2_u5_u6_n127 ) );
  NAND3_X1 u2_u5_u6_U91 (.ZN( u2_u5_u6_n102 ) , .A3( u2_u5_u6_n130 ) , .A2( u2_u5_u6_n145 ) , .A1( u2_u5_u6_n166 ) );
  NAND3_X1 u2_u5_u6_U92 (.A3( u2_u5_u6_n113 ) , .A1( u2_u5_u6_n119 ) , .A2( u2_u5_u6_n123 ) , .ZN( u2_u5_u6_n93 ) );
  NAND3_X1 u2_u5_u6_U93 (.ZN( u2_u5_u6_n142 ) , .A2( u2_u5_u6_n172 ) , .A3( u2_u5_u6_n89 ) , .A1( u2_u5_u6_n90 ) );
  AND3_X1 u2_u5_u7_U10 (.A3( u2_u5_u7_n110 ) , .A2( u2_u5_u7_n127 ) , .A1( u2_u5_u7_n132 ) , .ZN( u2_u5_u7_n92 ) );
  OAI21_X1 u2_u5_u7_U11 (.A( u2_u5_u7_n161 ) , .B1( u2_u5_u7_n168 ) , .B2( u2_u5_u7_n173 ) , .ZN( u2_u5_u7_n91 ) );
  AOI211_X1 u2_u5_u7_U12 (.A( u2_u5_u7_n117 ) , .ZN( u2_u5_u7_n118 ) , .C2( u2_u5_u7_n126 ) , .C1( u2_u5_u7_n177 ) , .B( u2_u5_u7_n180 ) );
  OAI22_X1 u2_u5_u7_U13 (.B1( u2_u5_u7_n115 ) , .ZN( u2_u5_u7_n117 ) , .A2( u2_u5_u7_n133 ) , .A1( u2_u5_u7_n137 ) , .B2( u2_u5_u7_n162 ) );
  INV_X1 u2_u5_u7_U14 (.A( u2_u5_u7_n116 ) , .ZN( u2_u5_u7_n180 ) );
  NOR3_X1 u2_u5_u7_U15 (.ZN( u2_u5_u7_n115 ) , .A3( u2_u5_u7_n145 ) , .A2( u2_u5_u7_n168 ) , .A1( u2_u5_u7_n169 ) );
  OAI211_X1 u2_u5_u7_U16 (.B( u2_u5_u7_n122 ) , .A( u2_u5_u7_n123 ) , .C2( u2_u5_u7_n124 ) , .ZN( u2_u5_u7_n154 ) , .C1( u2_u5_u7_n162 ) );
  AOI222_X1 u2_u5_u7_U17 (.ZN( u2_u5_u7_n122 ) , .C2( u2_u5_u7_n126 ) , .C1( u2_u5_u7_n145 ) , .B1( u2_u5_u7_n161 ) , .A2( u2_u5_u7_n165 ) , .B2( u2_u5_u7_n170 ) , .A1( u2_u5_u7_n176 ) );
  INV_X1 u2_u5_u7_U18 (.A( u2_u5_u7_n133 ) , .ZN( u2_u5_u7_n176 ) );
  NOR3_X1 u2_u5_u7_U19 (.A2( u2_u5_u7_n134 ) , .A1( u2_u5_u7_n135 ) , .ZN( u2_u5_u7_n136 ) , .A3( u2_u5_u7_n171 ) );
  NOR2_X1 u2_u5_u7_U20 (.A1( u2_u5_u7_n130 ) , .A2( u2_u5_u7_n134 ) , .ZN( u2_u5_u7_n153 ) );
  INV_X1 u2_u5_u7_U21 (.A( u2_u5_u7_n101 ) , .ZN( u2_u5_u7_n165 ) );
  NOR2_X1 u2_u5_u7_U22 (.ZN( u2_u5_u7_n111 ) , .A2( u2_u5_u7_n134 ) , .A1( u2_u5_u7_n169 ) );
  AOI21_X1 u2_u5_u7_U23 (.ZN( u2_u5_u7_n104 ) , .B2( u2_u5_u7_n112 ) , .B1( u2_u5_u7_n127 ) , .A( u2_u5_u7_n164 ) );
  AOI21_X1 u2_u5_u7_U24 (.ZN( u2_u5_u7_n106 ) , .B1( u2_u5_u7_n133 ) , .B2( u2_u5_u7_n146 ) , .A( u2_u5_u7_n162 ) );
  AOI21_X1 u2_u5_u7_U25 (.A( u2_u5_u7_n101 ) , .ZN( u2_u5_u7_n107 ) , .B2( u2_u5_u7_n128 ) , .B1( u2_u5_u7_n175 ) );
  INV_X1 u2_u5_u7_U26 (.A( u2_u5_u7_n138 ) , .ZN( u2_u5_u7_n171 ) );
  INV_X1 u2_u5_u7_U27 (.A( u2_u5_u7_n131 ) , .ZN( u2_u5_u7_n177 ) );
  INV_X1 u2_u5_u7_U28 (.A( u2_u5_u7_n110 ) , .ZN( u2_u5_u7_n174 ) );
  NAND2_X1 u2_u5_u7_U29 (.A1( u2_u5_u7_n129 ) , .A2( u2_u5_u7_n132 ) , .ZN( u2_u5_u7_n149 ) );
  OAI21_X1 u2_u5_u7_U3 (.ZN( u2_u5_u7_n159 ) , .A( u2_u5_u7_n165 ) , .B2( u2_u5_u7_n171 ) , .B1( u2_u5_u7_n174 ) );
  NAND2_X1 u2_u5_u7_U30 (.A1( u2_u5_u7_n113 ) , .A2( u2_u5_u7_n124 ) , .ZN( u2_u5_u7_n130 ) );
  INV_X1 u2_u5_u7_U31 (.A( u2_u5_u7_n112 ) , .ZN( u2_u5_u7_n173 ) );
  INV_X1 u2_u5_u7_U32 (.A( u2_u5_u7_n128 ) , .ZN( u2_u5_u7_n168 ) );
  INV_X1 u2_u5_u7_U33 (.A( u2_u5_u7_n148 ) , .ZN( u2_u5_u7_n169 ) );
  INV_X1 u2_u5_u7_U34 (.A( u2_u5_u7_n127 ) , .ZN( u2_u5_u7_n179 ) );
  NOR2_X1 u2_u5_u7_U35 (.ZN( u2_u5_u7_n101 ) , .A2( u2_u5_u7_n150 ) , .A1( u2_u5_u7_n156 ) );
  AOI211_X1 u2_u5_u7_U36 (.B( u2_u5_u7_n154 ) , .A( u2_u5_u7_n155 ) , .C1( u2_u5_u7_n156 ) , .ZN( u2_u5_u7_n157 ) , .C2( u2_u5_u7_n172 ) );
  INV_X1 u2_u5_u7_U37 (.A( u2_u5_u7_n153 ) , .ZN( u2_u5_u7_n172 ) );
  AOI211_X1 u2_u5_u7_U38 (.B( u2_u5_u7_n139 ) , .A( u2_u5_u7_n140 ) , .C2( u2_u5_u7_n141 ) , .ZN( u2_u5_u7_n142 ) , .C1( u2_u5_u7_n156 ) );
  NAND4_X1 u2_u5_u7_U39 (.A3( u2_u5_u7_n127 ) , .A2( u2_u5_u7_n128 ) , .A1( u2_u5_u7_n129 ) , .ZN( u2_u5_u7_n141 ) , .A4( u2_u5_u7_n147 ) );
  INV_X1 u2_u5_u7_U4 (.A( u2_u5_u7_n111 ) , .ZN( u2_u5_u7_n170 ) );
  AOI21_X1 u2_u5_u7_U40 (.A( u2_u5_u7_n137 ) , .B1( u2_u5_u7_n138 ) , .ZN( u2_u5_u7_n139 ) , .B2( u2_u5_u7_n146 ) );
  OAI22_X1 u2_u5_u7_U41 (.B1( u2_u5_u7_n136 ) , .ZN( u2_u5_u7_n140 ) , .A1( u2_u5_u7_n153 ) , .B2( u2_u5_u7_n162 ) , .A2( u2_u5_u7_n164 ) );
  AOI21_X1 u2_u5_u7_U42 (.ZN( u2_u5_u7_n123 ) , .B1( u2_u5_u7_n165 ) , .B2( u2_u5_u7_n177 ) , .A( u2_u5_u7_n97 ) );
  AOI21_X1 u2_u5_u7_U43 (.B2( u2_u5_u7_n113 ) , .B1( u2_u5_u7_n124 ) , .A( u2_u5_u7_n125 ) , .ZN( u2_u5_u7_n97 ) );
  INV_X1 u2_u5_u7_U44 (.A( u2_u5_u7_n125 ) , .ZN( u2_u5_u7_n161 ) );
  INV_X1 u2_u5_u7_U45 (.A( u2_u5_u7_n152 ) , .ZN( u2_u5_u7_n162 ) );
  AOI22_X1 u2_u5_u7_U46 (.A2( u2_u5_u7_n114 ) , .ZN( u2_u5_u7_n119 ) , .B1( u2_u5_u7_n130 ) , .A1( u2_u5_u7_n156 ) , .B2( u2_u5_u7_n165 ) );
  NAND2_X1 u2_u5_u7_U47 (.A2( u2_u5_u7_n112 ) , .ZN( u2_u5_u7_n114 ) , .A1( u2_u5_u7_n175 ) );
  AND2_X1 u2_u5_u7_U48 (.ZN( u2_u5_u7_n145 ) , .A2( u2_u5_u7_n98 ) , .A1( u2_u5_u7_n99 ) );
  NOR2_X1 u2_u5_u7_U49 (.ZN( u2_u5_u7_n137 ) , .A1( u2_u5_u7_n150 ) , .A2( u2_u5_u7_n161 ) );
  INV_X1 u2_u5_u7_U5 (.A( u2_u5_u7_n149 ) , .ZN( u2_u5_u7_n175 ) );
  AOI21_X1 u2_u5_u7_U50 (.ZN( u2_u5_u7_n105 ) , .B2( u2_u5_u7_n110 ) , .A( u2_u5_u7_n125 ) , .B1( u2_u5_u7_n147 ) );
  NAND2_X1 u2_u5_u7_U51 (.ZN( u2_u5_u7_n146 ) , .A1( u2_u5_u7_n95 ) , .A2( u2_u5_u7_n98 ) );
  NAND2_X1 u2_u5_u7_U52 (.A2( u2_u5_u7_n103 ) , .ZN( u2_u5_u7_n147 ) , .A1( u2_u5_u7_n93 ) );
  NAND2_X1 u2_u5_u7_U53 (.A1( u2_u5_u7_n103 ) , .ZN( u2_u5_u7_n127 ) , .A2( u2_u5_u7_n99 ) );
  OR2_X1 u2_u5_u7_U54 (.ZN( u2_u5_u7_n126 ) , .A2( u2_u5_u7_n152 ) , .A1( u2_u5_u7_n156 ) );
  NAND2_X1 u2_u5_u7_U55 (.A2( u2_u5_u7_n102 ) , .A1( u2_u5_u7_n103 ) , .ZN( u2_u5_u7_n133 ) );
  NAND2_X1 u2_u5_u7_U56 (.ZN( u2_u5_u7_n112 ) , .A2( u2_u5_u7_n96 ) , .A1( u2_u5_u7_n99 ) );
  NAND2_X1 u2_u5_u7_U57 (.A2( u2_u5_u7_n102 ) , .ZN( u2_u5_u7_n128 ) , .A1( u2_u5_u7_n98 ) );
  NAND2_X1 u2_u5_u7_U58 (.A1( u2_u5_u7_n100 ) , .ZN( u2_u5_u7_n113 ) , .A2( u2_u5_u7_n93 ) );
  NAND2_X1 u2_u5_u7_U59 (.A2( u2_u5_u7_n102 ) , .ZN( u2_u5_u7_n124 ) , .A1( u2_u5_u7_n96 ) );
  INV_X1 u2_u5_u7_U6 (.A( u2_u5_u7_n154 ) , .ZN( u2_u5_u7_n178 ) );
  NAND2_X1 u2_u5_u7_U60 (.ZN( u2_u5_u7_n110 ) , .A1( u2_u5_u7_n95 ) , .A2( u2_u5_u7_n96 ) );
  INV_X1 u2_u5_u7_U61 (.A( u2_u5_u7_n150 ) , .ZN( u2_u5_u7_n164 ) );
  AND2_X1 u2_u5_u7_U62 (.ZN( u2_u5_u7_n134 ) , .A1( u2_u5_u7_n93 ) , .A2( u2_u5_u7_n98 ) );
  NAND2_X1 u2_u5_u7_U63 (.A1( u2_u5_u7_n100 ) , .A2( u2_u5_u7_n102 ) , .ZN( u2_u5_u7_n129 ) );
  NAND2_X1 u2_u5_u7_U64 (.A2( u2_u5_u7_n103 ) , .ZN( u2_u5_u7_n131 ) , .A1( u2_u5_u7_n95 ) );
  NAND2_X1 u2_u5_u7_U65 (.A1( u2_u5_u7_n100 ) , .ZN( u2_u5_u7_n138 ) , .A2( u2_u5_u7_n99 ) );
  NAND2_X1 u2_u5_u7_U66 (.ZN( u2_u5_u7_n132 ) , .A1( u2_u5_u7_n93 ) , .A2( u2_u5_u7_n96 ) );
  NAND2_X1 u2_u5_u7_U67 (.A1( u2_u5_u7_n100 ) , .ZN( u2_u5_u7_n148 ) , .A2( u2_u5_u7_n95 ) );
  NOR2_X1 u2_u5_u7_U68 (.A2( u2_u5_X_47 ) , .ZN( u2_u5_u7_n150 ) , .A1( u2_u5_u7_n163 ) );
  NOR2_X1 u2_u5_u7_U69 (.A2( u2_u5_X_43 ) , .A1( u2_u5_X_44 ) , .ZN( u2_u5_u7_n103 ) );
  AOI211_X1 u2_u5_u7_U7 (.ZN( u2_u5_u7_n116 ) , .A( u2_u5_u7_n155 ) , .C1( u2_u5_u7_n161 ) , .C2( u2_u5_u7_n171 ) , .B( u2_u5_u7_n94 ) );
  NOR2_X1 u2_u5_u7_U70 (.A2( u2_u5_X_48 ) , .A1( u2_u5_u7_n166 ) , .ZN( u2_u5_u7_n95 ) );
  NOR2_X1 u2_u5_u7_U71 (.A2( u2_u5_X_45 ) , .A1( u2_u5_X_48 ) , .ZN( u2_u5_u7_n99 ) );
  NOR2_X1 u2_u5_u7_U72 (.A2( u2_u5_X_44 ) , .A1( u2_u5_u7_n167 ) , .ZN( u2_u5_u7_n98 ) );
  NOR2_X1 u2_u5_u7_U73 (.A2( u2_u5_X_46 ) , .A1( u2_u5_X_47 ) , .ZN( u2_u5_u7_n152 ) );
  AND2_X1 u2_u5_u7_U74 (.A1( u2_u5_X_47 ) , .ZN( u2_u5_u7_n156 ) , .A2( u2_u5_u7_n163 ) );
  NAND2_X1 u2_u5_u7_U75 (.A2( u2_u5_X_46 ) , .A1( u2_u5_X_47 ) , .ZN( u2_u5_u7_n125 ) );
  AND2_X1 u2_u5_u7_U76 (.A2( u2_u5_X_45 ) , .A1( u2_u5_X_48 ) , .ZN( u2_u5_u7_n102 ) );
  AND2_X1 u2_u5_u7_U77 (.A2( u2_u5_X_43 ) , .A1( u2_u5_X_44 ) , .ZN( u2_u5_u7_n96 ) );
  AND2_X1 u2_u5_u7_U78 (.A1( u2_u5_X_44 ) , .ZN( u2_u5_u7_n100 ) , .A2( u2_u5_u7_n167 ) );
  AND2_X1 u2_u5_u7_U79 (.A1( u2_u5_X_48 ) , .A2( u2_u5_u7_n166 ) , .ZN( u2_u5_u7_n93 ) );
  OAI222_X1 u2_u5_u7_U8 (.C2( u2_u5_u7_n101 ) , .B2( u2_u5_u7_n111 ) , .A1( u2_u5_u7_n113 ) , .C1( u2_u5_u7_n146 ) , .A2( u2_u5_u7_n162 ) , .B1( u2_u5_u7_n164 ) , .ZN( u2_u5_u7_n94 ) );
  INV_X1 u2_u5_u7_U80 (.A( u2_u5_X_46 ) , .ZN( u2_u5_u7_n163 ) );
  INV_X1 u2_u5_u7_U81 (.A( u2_u5_X_43 ) , .ZN( u2_u5_u7_n167 ) );
  INV_X1 u2_u5_u7_U82 (.A( u2_u5_X_45 ) , .ZN( u2_u5_u7_n166 ) );
  NAND4_X1 u2_u5_u7_U83 (.ZN( u2_out5_27 ) , .A4( u2_u5_u7_n118 ) , .A3( u2_u5_u7_n119 ) , .A2( u2_u5_u7_n120 ) , .A1( u2_u5_u7_n121 ) );
  OAI21_X1 u2_u5_u7_U84 (.ZN( u2_u5_u7_n121 ) , .B2( u2_u5_u7_n145 ) , .A( u2_u5_u7_n150 ) , .B1( u2_u5_u7_n174 ) );
  OAI21_X1 u2_u5_u7_U85 (.ZN( u2_u5_u7_n120 ) , .A( u2_u5_u7_n161 ) , .B2( u2_u5_u7_n170 ) , .B1( u2_u5_u7_n179 ) );
  NAND4_X1 u2_u5_u7_U86 (.ZN( u2_out5_21 ) , .A4( u2_u5_u7_n157 ) , .A3( u2_u5_u7_n158 ) , .A2( u2_u5_u7_n159 ) , .A1( u2_u5_u7_n160 ) );
  OAI21_X1 u2_u5_u7_U87 (.B1( u2_u5_u7_n145 ) , .ZN( u2_u5_u7_n160 ) , .A( u2_u5_u7_n161 ) , .B2( u2_u5_u7_n177 ) );
  AOI22_X1 u2_u5_u7_U88 (.B2( u2_u5_u7_n149 ) , .B1( u2_u5_u7_n150 ) , .A2( u2_u5_u7_n151 ) , .A1( u2_u5_u7_n152 ) , .ZN( u2_u5_u7_n158 ) );
  NAND4_X1 u2_u5_u7_U89 (.ZN( u2_out5_15 ) , .A4( u2_u5_u7_n142 ) , .A3( u2_u5_u7_n143 ) , .A2( u2_u5_u7_n144 ) , .A1( u2_u5_u7_n178 ) );
  OAI221_X1 u2_u5_u7_U9 (.C1( u2_u5_u7_n101 ) , .C2( u2_u5_u7_n147 ) , .ZN( u2_u5_u7_n155 ) , .B2( u2_u5_u7_n162 ) , .A( u2_u5_u7_n91 ) , .B1( u2_u5_u7_n92 ) );
  OR2_X1 u2_u5_u7_U90 (.A2( u2_u5_u7_n125 ) , .A1( u2_u5_u7_n129 ) , .ZN( u2_u5_u7_n144 ) );
  AOI22_X1 u2_u5_u7_U91 (.A2( u2_u5_u7_n126 ) , .ZN( u2_u5_u7_n143 ) , .B2( u2_u5_u7_n165 ) , .B1( u2_u5_u7_n173 ) , .A1( u2_u5_u7_n174 ) );
  NAND4_X1 u2_u5_u7_U92 (.ZN( u2_out5_5 ) , .A4( u2_u5_u7_n108 ) , .A3( u2_u5_u7_n109 ) , .A1( u2_u5_u7_n116 ) , .A2( u2_u5_u7_n123 ) );
  AOI22_X1 u2_u5_u7_U93 (.ZN( u2_u5_u7_n109 ) , .A2( u2_u5_u7_n126 ) , .B2( u2_u5_u7_n145 ) , .B1( u2_u5_u7_n156 ) , .A1( u2_u5_u7_n171 ) );
  NOR4_X1 u2_u5_u7_U94 (.A4( u2_u5_u7_n104 ) , .A3( u2_u5_u7_n105 ) , .A2( u2_u5_u7_n106 ) , .A1( u2_u5_u7_n107 ) , .ZN( u2_u5_u7_n108 ) );
  NAND3_X1 u2_u5_u7_U95 (.A3( u2_u5_u7_n146 ) , .A2( u2_u5_u7_n147 ) , .A1( u2_u5_u7_n148 ) , .ZN( u2_u5_u7_n151 ) );
  NAND3_X1 u2_u5_u7_U96 (.A3( u2_u5_u7_n131 ) , .A2( u2_u5_u7_n132 ) , .A1( u2_u5_u7_n133 ) , .ZN( u2_u5_u7_n135 ) );
  XOR2_X1 u2_u6_U11 (.B( u2_K7_44 ) , .A( u2_R5_29 ) , .Z( u2_u6_X_44 ) );
  XOR2_X1 u2_u6_U12 (.B( u2_K7_43 ) , .A( u2_R5_28 ) , .Z( u2_u6_X_43 ) );
  XOR2_X1 u2_u6_U13 (.B( u2_K7_42 ) , .A( u2_R5_29 ) , .Z( u2_u6_X_42 ) );
  XOR2_X1 u2_u6_U14 (.B( u2_K7_41 ) , .A( u2_R5_28 ) , .Z( u2_u6_X_41 ) );
  XOR2_X1 u2_u6_U17 (.B( u2_K7_39 ) , .A( u2_R5_26 ) , .Z( u2_u6_X_39 ) );
  XOR2_X1 u2_u6_U18 (.B( u2_K7_38 ) , .A( u2_R5_25 ) , .Z( u2_u6_X_38 ) );
  XOR2_X1 u2_u6_U19 (.B( u2_K7_37 ) , .A( u2_R5_24 ) , .Z( u2_u6_X_37 ) );
  XOR2_X1 u2_u6_U2 (.B( u2_K7_8 ) , .A( u2_R5_5 ) , .Z( u2_u6_X_8 ) );
  XOR2_X1 u2_u6_U20 (.B( u2_K7_36 ) , .A( u2_R5_25 ) , .Z( u2_u6_X_36 ) );
  XOR2_X1 u2_u6_U21 (.B( u2_K7_35 ) , .A( u2_R5_24 ) , .Z( u2_u6_X_35 ) );
  XOR2_X1 u2_u6_U22 (.B( u2_K7_34 ) , .A( u2_R5_23 ) , .Z( u2_u6_X_34 ) );
  XOR2_X1 u2_u6_U24 (.B( u2_K7_32 ) , .A( u2_R5_21 ) , .Z( u2_u6_X_32 ) );
  XOR2_X1 u2_u6_U25 (.B( u2_K7_31 ) , .A( u2_R5_20 ) , .Z( u2_u6_X_31 ) );
  XOR2_X1 u2_u6_U26 (.B( u2_K7_30 ) , .A( u2_R5_21 ) , .Z( u2_u6_X_30 ) );
  XOR2_X1 u2_u6_U27 (.B( u2_K7_2 ) , .A( u2_R5_1 ) , .Z( u2_u6_X_2 ) );
  XOR2_X1 u2_u6_U28 (.B( u2_K7_29 ) , .A( u2_R5_20 ) , .Z( u2_u6_X_29 ) );
  XOR2_X1 u2_u6_U3 (.B( u2_K7_7 ) , .A( u2_R5_4 ) , .Z( u2_u6_X_7 ) );
  XOR2_X1 u2_u6_U31 (.B( u2_K7_26 ) , .A( u2_R5_17 ) , .Z( u2_u6_X_26 ) );
  XOR2_X1 u2_u6_U32 (.B( u2_K7_25 ) , .A( u2_R5_16 ) , .Z( u2_u6_X_25 ) );
  XOR2_X1 u2_u6_U33 (.B( u2_K7_24 ) , .A( u2_R5_17 ) , .Z( u2_u6_X_24 ) );
  XOR2_X1 u2_u6_U34 (.B( u2_K7_23 ) , .A( u2_R5_16 ) , .Z( u2_u6_X_23 ) );
  XOR2_X1 u2_u6_U36 (.B( u2_K7_21 ) , .A( u2_R5_14 ) , .Z( u2_u6_X_21 ) );
  XOR2_X1 u2_u6_U37 (.B( u2_K7_20 ) , .A( u2_R5_13 ) , .Z( u2_u6_X_20 ) );
  XOR2_X1 u2_u6_U38 (.B( u2_K7_1 ) , .A( u2_R5_32 ) , .Z( u2_u6_X_1 ) );
  XOR2_X1 u2_u6_U39 (.B( u2_K7_19 ) , .A( u2_R5_12 ) , .Z( u2_u6_X_19 ) );
  XOR2_X1 u2_u6_U4 (.B( u2_K7_6 ) , .A( u2_R5_5 ) , .Z( u2_u6_X_6 ) );
  XOR2_X1 u2_u6_U40 (.B( u2_K7_18 ) , .A( u2_R5_13 ) , .Z( u2_u6_X_18 ) );
  XOR2_X1 u2_u6_U41 (.B( u2_K7_17 ) , .A( u2_R5_12 ) , .Z( u2_u6_X_17 ) );
  XOR2_X1 u2_u6_U42 (.B( u2_K7_16 ) , .A( u2_R5_11 ) , .Z( u2_u6_X_16 ) );
  XOR2_X1 u2_u6_U43 (.B( u2_K7_15 ) , .A( u2_R5_10 ) , .Z( u2_u6_X_15 ) );
  XOR2_X1 u2_u6_U44 (.B( u2_K7_14 ) , .A( u2_R5_9 ) , .Z( u2_u6_X_14 ) );
  XOR2_X1 u2_u6_U45 (.B( u2_K7_13 ) , .A( u2_R5_8 ) , .Z( u2_u6_X_13 ) );
  XOR2_X1 u2_u6_U46 (.B( u2_K7_12 ) , .A( u2_R5_9 ) , .Z( u2_u6_X_12 ) );
  XOR2_X1 u2_u6_U47 (.B( u2_K7_11 ) , .A( u2_R5_8 ) , .Z( u2_u6_X_11 ) );
  XOR2_X1 u2_u6_U5 (.B( u2_K7_5 ) , .A( u2_R5_4 ) , .Z( u2_u6_X_5 ) );
  XOR2_X1 u2_u6_U7 (.B( u2_K7_48 ) , .A( u2_R5_1 ) , .Z( u2_u6_X_48 ) );
  XOR2_X1 u2_u6_U8 (.B( u2_K7_47 ) , .A( u2_R5_32 ) , .Z( u2_u6_X_47 ) );
  AND3_X1 u2_u6_u0_U10 (.A2( u2_u6_u0_n112 ) , .ZN( u2_u6_u0_n127 ) , .A3( u2_u6_u0_n130 ) , .A1( u2_u6_u0_n148 ) );
  NAND2_X1 u2_u6_u0_U11 (.ZN( u2_u6_u0_n113 ) , .A1( u2_u6_u0_n139 ) , .A2( u2_u6_u0_n149 ) );
  AND2_X1 u2_u6_u0_U12 (.ZN( u2_u6_u0_n107 ) , .A1( u2_u6_u0_n130 ) , .A2( u2_u6_u0_n140 ) );
  AND2_X1 u2_u6_u0_U13 (.A2( u2_u6_u0_n129 ) , .A1( u2_u6_u0_n130 ) , .ZN( u2_u6_u0_n151 ) );
  AND2_X1 u2_u6_u0_U14 (.A1( u2_u6_u0_n108 ) , .A2( u2_u6_u0_n125 ) , .ZN( u2_u6_u0_n145 ) );
  INV_X1 u2_u6_u0_U15 (.A( u2_u6_u0_n143 ) , .ZN( u2_u6_u0_n173 ) );
  NOR2_X1 u2_u6_u0_U16 (.A2( u2_u6_u0_n136 ) , .ZN( u2_u6_u0_n147 ) , .A1( u2_u6_u0_n160 ) );
  NOR2_X1 u2_u6_u0_U17 (.A1( u2_u6_u0_n163 ) , .A2( u2_u6_u0_n164 ) , .ZN( u2_u6_u0_n95 ) );
  AOI21_X1 u2_u6_u0_U18 (.B1( u2_u6_u0_n103 ) , .ZN( u2_u6_u0_n132 ) , .A( u2_u6_u0_n165 ) , .B2( u2_u6_u0_n93 ) );
  INV_X1 u2_u6_u0_U19 (.A( u2_u6_u0_n142 ) , .ZN( u2_u6_u0_n165 ) );
  OAI22_X1 u2_u6_u0_U20 (.B1( u2_u6_u0_n125 ) , .ZN( u2_u6_u0_n126 ) , .A1( u2_u6_u0_n138 ) , .A2( u2_u6_u0_n146 ) , .B2( u2_u6_u0_n147 ) );
  OAI22_X1 u2_u6_u0_U21 (.B1( u2_u6_u0_n131 ) , .A1( u2_u6_u0_n144 ) , .B2( u2_u6_u0_n147 ) , .A2( u2_u6_u0_n90 ) , .ZN( u2_u6_u0_n91 ) );
  AND3_X1 u2_u6_u0_U22 (.A3( u2_u6_u0_n121 ) , .A2( u2_u6_u0_n125 ) , .A1( u2_u6_u0_n148 ) , .ZN( u2_u6_u0_n90 ) );
  NAND2_X1 u2_u6_u0_U23 (.A1( u2_u6_u0_n100 ) , .A2( u2_u6_u0_n103 ) , .ZN( u2_u6_u0_n125 ) );
  INV_X1 u2_u6_u0_U24 (.A( u2_u6_u0_n136 ) , .ZN( u2_u6_u0_n161 ) );
  AOI22_X1 u2_u6_u0_U25 (.B2( u2_u6_u0_n109 ) , .A2( u2_u6_u0_n110 ) , .ZN( u2_u6_u0_n111 ) , .B1( u2_u6_u0_n118 ) , .A1( u2_u6_u0_n160 ) );
  NAND2_X1 u2_u6_u0_U26 (.A1( u2_u6_u0_n100 ) , .ZN( u2_u6_u0_n129 ) , .A2( u2_u6_u0_n95 ) );
  INV_X1 u2_u6_u0_U27 (.A( u2_u6_u0_n118 ) , .ZN( u2_u6_u0_n158 ) );
  AOI21_X1 u2_u6_u0_U28 (.ZN( u2_u6_u0_n104 ) , .B1( u2_u6_u0_n107 ) , .B2( u2_u6_u0_n141 ) , .A( u2_u6_u0_n144 ) );
  AOI21_X1 u2_u6_u0_U29 (.B1( u2_u6_u0_n127 ) , .B2( u2_u6_u0_n129 ) , .A( u2_u6_u0_n138 ) , .ZN( u2_u6_u0_n96 ) );
  INV_X1 u2_u6_u0_U3 (.A( u2_u6_u0_n113 ) , .ZN( u2_u6_u0_n166 ) );
  AOI21_X1 u2_u6_u0_U30 (.ZN( u2_u6_u0_n116 ) , .B2( u2_u6_u0_n142 ) , .A( u2_u6_u0_n144 ) , .B1( u2_u6_u0_n166 ) );
  NOR2_X1 u2_u6_u0_U31 (.A1( u2_u6_u0_n120 ) , .ZN( u2_u6_u0_n143 ) , .A2( u2_u6_u0_n167 ) );
  OAI221_X1 u2_u6_u0_U32 (.C1( u2_u6_u0_n112 ) , .ZN( u2_u6_u0_n120 ) , .B1( u2_u6_u0_n138 ) , .B2( u2_u6_u0_n141 ) , .C2( u2_u6_u0_n147 ) , .A( u2_u6_u0_n172 ) );
  AOI211_X1 u2_u6_u0_U33 (.B( u2_u6_u0_n115 ) , .A( u2_u6_u0_n116 ) , .C2( u2_u6_u0_n117 ) , .C1( u2_u6_u0_n118 ) , .ZN( u2_u6_u0_n119 ) );
  NAND2_X1 u2_u6_u0_U34 (.A2( u2_u6_u0_n100 ) , .A1( u2_u6_u0_n101 ) , .ZN( u2_u6_u0_n139 ) );
  NAND2_X1 u2_u6_u0_U35 (.A2( u2_u6_u0_n100 ) , .ZN( u2_u6_u0_n131 ) , .A1( u2_u6_u0_n92 ) );
  NAND2_X1 u2_u6_u0_U36 (.A1( u2_u6_u0_n101 ) , .A2( u2_u6_u0_n102 ) , .ZN( u2_u6_u0_n150 ) );
  INV_X1 u2_u6_u0_U37 (.A( u2_u6_u0_n138 ) , .ZN( u2_u6_u0_n160 ) );
  NAND2_X1 u2_u6_u0_U38 (.A1( u2_u6_u0_n102 ) , .ZN( u2_u6_u0_n128 ) , .A2( u2_u6_u0_n95 ) );
  NAND2_X1 u2_u6_u0_U39 (.ZN( u2_u6_u0_n148 ) , .A1( u2_u6_u0_n93 ) , .A2( u2_u6_u0_n95 ) );
  AOI21_X1 u2_u6_u0_U4 (.B1( u2_u6_u0_n114 ) , .ZN( u2_u6_u0_n115 ) , .B2( u2_u6_u0_n129 ) , .A( u2_u6_u0_n161 ) );
  NAND2_X1 u2_u6_u0_U40 (.A2( u2_u6_u0_n102 ) , .A1( u2_u6_u0_n103 ) , .ZN( u2_u6_u0_n149 ) );
  NAND2_X1 u2_u6_u0_U41 (.A2( u2_u6_u0_n102 ) , .ZN( u2_u6_u0_n114 ) , .A1( u2_u6_u0_n92 ) );
  NAND2_X1 u2_u6_u0_U42 (.A2( u2_u6_u0_n101 ) , .ZN( u2_u6_u0_n121 ) , .A1( u2_u6_u0_n93 ) );
  NAND2_X1 u2_u6_u0_U43 (.ZN( u2_u6_u0_n112 ) , .A2( u2_u6_u0_n92 ) , .A1( u2_u6_u0_n93 ) );
  INV_X1 u2_u6_u0_U44 (.ZN( u2_u6_u0_n172 ) , .A( u2_u6_u0_n88 ) );
  OAI222_X1 u2_u6_u0_U45 (.C1( u2_u6_u0_n108 ) , .A1( u2_u6_u0_n125 ) , .B2( u2_u6_u0_n128 ) , .B1( u2_u6_u0_n144 ) , .A2( u2_u6_u0_n158 ) , .C2( u2_u6_u0_n161 ) , .ZN( u2_u6_u0_n88 ) );
  OR3_X1 u2_u6_u0_U46 (.A3( u2_u6_u0_n152 ) , .A2( u2_u6_u0_n153 ) , .A1( u2_u6_u0_n154 ) , .ZN( u2_u6_u0_n155 ) );
  AOI21_X1 u2_u6_u0_U47 (.A( u2_u6_u0_n144 ) , .B2( u2_u6_u0_n145 ) , .B1( u2_u6_u0_n146 ) , .ZN( u2_u6_u0_n154 ) );
  AOI21_X1 u2_u6_u0_U48 (.B2( u2_u6_u0_n150 ) , .B1( u2_u6_u0_n151 ) , .ZN( u2_u6_u0_n152 ) , .A( u2_u6_u0_n158 ) );
  AOI21_X1 u2_u6_u0_U49 (.A( u2_u6_u0_n147 ) , .B2( u2_u6_u0_n148 ) , .B1( u2_u6_u0_n149 ) , .ZN( u2_u6_u0_n153 ) );
  AOI21_X1 u2_u6_u0_U5 (.B2( u2_u6_u0_n131 ) , .ZN( u2_u6_u0_n134 ) , .B1( u2_u6_u0_n151 ) , .A( u2_u6_u0_n158 ) );
  INV_X1 u2_u6_u0_U50 (.ZN( u2_u6_u0_n171 ) , .A( u2_u6_u0_n99 ) );
  OAI211_X1 u2_u6_u0_U51 (.C2( u2_u6_u0_n140 ) , .C1( u2_u6_u0_n161 ) , .A( u2_u6_u0_n169 ) , .B( u2_u6_u0_n98 ) , .ZN( u2_u6_u0_n99 ) );
  INV_X1 u2_u6_u0_U52 (.ZN( u2_u6_u0_n169 ) , .A( u2_u6_u0_n91 ) );
  AOI211_X1 u2_u6_u0_U53 (.C1( u2_u6_u0_n118 ) , .A( u2_u6_u0_n123 ) , .B( u2_u6_u0_n96 ) , .C2( u2_u6_u0_n97 ) , .ZN( u2_u6_u0_n98 ) );
  NOR2_X1 u2_u6_u0_U54 (.A2( u2_u6_X_4 ) , .A1( u2_u6_X_5 ) , .ZN( u2_u6_u0_n118 ) );
  NOR2_X1 u2_u6_u0_U55 (.A2( u2_u6_X_2 ) , .ZN( u2_u6_u0_n103 ) , .A1( u2_u6_u0_n164 ) );
  NOR2_X1 u2_u6_u0_U56 (.A2( u2_u6_X_1 ) , .A1( u2_u6_X_2 ) , .ZN( u2_u6_u0_n92 ) );
  NOR2_X1 u2_u6_u0_U57 (.A2( u2_u6_X_1 ) , .ZN( u2_u6_u0_n101 ) , .A1( u2_u6_u0_n163 ) );
  NAND2_X1 u2_u6_u0_U58 (.A2( u2_u6_X_4 ) , .A1( u2_u6_X_5 ) , .ZN( u2_u6_u0_n144 ) );
  NOR2_X1 u2_u6_u0_U59 (.A2( u2_u6_X_5 ) , .ZN( u2_u6_u0_n136 ) , .A1( u2_u6_u0_n159 ) );
  NOR2_X1 u2_u6_u0_U6 (.A1( u2_u6_u0_n108 ) , .ZN( u2_u6_u0_n123 ) , .A2( u2_u6_u0_n158 ) );
  NAND2_X1 u2_u6_u0_U60 (.A1( u2_u6_X_5 ) , .ZN( u2_u6_u0_n138 ) , .A2( u2_u6_u0_n159 ) );
  INV_X1 u2_u6_u0_U61 (.A( u2_u6_X_4 ) , .ZN( u2_u6_u0_n159 ) );
  INV_X1 u2_u6_u0_U62 (.A( u2_u6_X_1 ) , .ZN( u2_u6_u0_n164 ) );
  INV_X1 u2_u6_u0_U63 (.A( u2_u6_X_2 ) , .ZN( u2_u6_u0_n163 ) );
  INV_X1 u2_u6_u0_U64 (.A( u2_u6_X_3 ) , .ZN( u2_u6_u0_n162 ) );
  INV_X1 u2_u6_u0_U65 (.A( u2_u6_u0_n126 ) , .ZN( u2_u6_u0_n168 ) );
  AOI211_X1 u2_u6_u0_U66 (.B( u2_u6_u0_n133 ) , .A( u2_u6_u0_n134 ) , .C2( u2_u6_u0_n135 ) , .C1( u2_u6_u0_n136 ) , .ZN( u2_u6_u0_n137 ) );
  OR4_X1 u2_u6_u0_U67 (.ZN( u2_out6_17 ) , .A4( u2_u6_u0_n122 ) , .A2( u2_u6_u0_n123 ) , .A1( u2_u6_u0_n124 ) , .A3( u2_u6_u0_n170 ) );
  AOI21_X1 u2_u6_u0_U68 (.B2( u2_u6_u0_n107 ) , .ZN( u2_u6_u0_n124 ) , .B1( u2_u6_u0_n128 ) , .A( u2_u6_u0_n161 ) );
  INV_X1 u2_u6_u0_U69 (.A( u2_u6_u0_n111 ) , .ZN( u2_u6_u0_n170 ) );
  OAI21_X1 u2_u6_u0_U7 (.B1( u2_u6_u0_n150 ) , .B2( u2_u6_u0_n158 ) , .A( u2_u6_u0_n172 ) , .ZN( u2_u6_u0_n89 ) );
  OR4_X1 u2_u6_u0_U70 (.ZN( u2_out6_31 ) , .A4( u2_u6_u0_n155 ) , .A2( u2_u6_u0_n156 ) , .A1( u2_u6_u0_n157 ) , .A3( u2_u6_u0_n173 ) );
  AOI21_X1 u2_u6_u0_U71 (.A( u2_u6_u0_n138 ) , .B2( u2_u6_u0_n139 ) , .B1( u2_u6_u0_n140 ) , .ZN( u2_u6_u0_n157 ) );
  AOI21_X1 u2_u6_u0_U72 (.B2( u2_u6_u0_n141 ) , .B1( u2_u6_u0_n142 ) , .ZN( u2_u6_u0_n156 ) , .A( u2_u6_u0_n161 ) );
  INV_X1 u2_u6_u0_U73 (.ZN( u2_u6_u0_n174 ) , .A( u2_u6_u0_n89 ) );
  AOI211_X1 u2_u6_u0_U74 (.B( u2_u6_u0_n104 ) , .A( u2_u6_u0_n105 ) , .ZN( u2_u6_u0_n106 ) , .C2( u2_u6_u0_n113 ) , .C1( u2_u6_u0_n160 ) );
  AND2_X1 u2_u6_u0_U75 (.A1( u2_u6_X_6 ) , .A2( u2_u6_u0_n162 ) , .ZN( u2_u6_u0_n93 ) );
  NOR2_X1 u2_u6_u0_U76 (.A2( u2_u6_X_3 ) , .A1( u2_u6_X_6 ) , .ZN( u2_u6_u0_n94 ) );
  NOR2_X1 u2_u6_u0_U77 (.A2( u2_u6_X_6 ) , .ZN( u2_u6_u0_n100 ) , .A1( u2_u6_u0_n162 ) );
  AND2_X1 u2_u6_u0_U78 (.A2( u2_u6_X_3 ) , .A1( u2_u6_X_6 ) , .ZN( u2_u6_u0_n102 ) );
  OAI221_X1 u2_u6_u0_U79 (.C1( u2_u6_u0_n121 ) , .ZN( u2_u6_u0_n122 ) , .B2( u2_u6_u0_n127 ) , .A( u2_u6_u0_n143 ) , .B1( u2_u6_u0_n144 ) , .C2( u2_u6_u0_n147 ) );
  AND2_X1 u2_u6_u0_U8 (.A1( u2_u6_u0_n114 ) , .A2( u2_u6_u0_n121 ) , .ZN( u2_u6_u0_n146 ) );
  AOI21_X1 u2_u6_u0_U80 (.B1( u2_u6_u0_n132 ) , .ZN( u2_u6_u0_n133 ) , .A( u2_u6_u0_n144 ) , .B2( u2_u6_u0_n166 ) );
  OAI22_X1 u2_u6_u0_U81 (.ZN( u2_u6_u0_n105 ) , .A2( u2_u6_u0_n132 ) , .B1( u2_u6_u0_n146 ) , .A1( u2_u6_u0_n147 ) , .B2( u2_u6_u0_n161 ) );
  NAND2_X1 u2_u6_u0_U82 (.ZN( u2_u6_u0_n110 ) , .A2( u2_u6_u0_n132 ) , .A1( u2_u6_u0_n145 ) );
  INV_X1 u2_u6_u0_U83 (.A( u2_u6_u0_n119 ) , .ZN( u2_u6_u0_n167 ) );
  NAND2_X1 u2_u6_u0_U84 (.A2( u2_u6_u0_n103 ) , .ZN( u2_u6_u0_n140 ) , .A1( u2_u6_u0_n94 ) );
  NAND2_X1 u2_u6_u0_U85 (.A1( u2_u6_u0_n101 ) , .ZN( u2_u6_u0_n130 ) , .A2( u2_u6_u0_n94 ) );
  NAND2_X1 u2_u6_u0_U86 (.ZN( u2_u6_u0_n108 ) , .A1( u2_u6_u0_n92 ) , .A2( u2_u6_u0_n94 ) );
  NAND2_X1 u2_u6_u0_U87 (.ZN( u2_u6_u0_n142 ) , .A1( u2_u6_u0_n94 ) , .A2( u2_u6_u0_n95 ) );
  NAND3_X1 u2_u6_u0_U88 (.ZN( u2_out6_23 ) , .A3( u2_u6_u0_n137 ) , .A1( u2_u6_u0_n168 ) , .A2( u2_u6_u0_n171 ) );
  NAND3_X1 u2_u6_u0_U89 (.A3( u2_u6_u0_n127 ) , .A2( u2_u6_u0_n128 ) , .ZN( u2_u6_u0_n135 ) , .A1( u2_u6_u0_n150 ) );
  AND2_X1 u2_u6_u0_U9 (.A1( u2_u6_u0_n131 ) , .ZN( u2_u6_u0_n141 ) , .A2( u2_u6_u0_n150 ) );
  NAND3_X1 u2_u6_u0_U90 (.ZN( u2_u6_u0_n117 ) , .A3( u2_u6_u0_n132 ) , .A2( u2_u6_u0_n139 ) , .A1( u2_u6_u0_n148 ) );
  NAND3_X1 u2_u6_u0_U91 (.ZN( u2_u6_u0_n109 ) , .A2( u2_u6_u0_n114 ) , .A3( u2_u6_u0_n140 ) , .A1( u2_u6_u0_n149 ) );
  NAND3_X1 u2_u6_u0_U92 (.ZN( u2_out6_9 ) , .A3( u2_u6_u0_n106 ) , .A2( u2_u6_u0_n171 ) , .A1( u2_u6_u0_n174 ) );
  NAND3_X1 u2_u6_u0_U93 (.A2( u2_u6_u0_n128 ) , .A1( u2_u6_u0_n132 ) , .A3( u2_u6_u0_n146 ) , .ZN( u2_u6_u0_n97 ) );
  AOI21_X1 u2_u6_u1_U10 (.B2( u2_u6_u1_n155 ) , .B1( u2_u6_u1_n156 ) , .ZN( u2_u6_u1_n157 ) , .A( u2_u6_u1_n174 ) );
  NAND3_X1 u2_u6_u1_U100 (.ZN( u2_u6_u1_n113 ) , .A1( u2_u6_u1_n120 ) , .A3( u2_u6_u1_n133 ) , .A2( u2_u6_u1_n155 ) );
  NAND2_X1 u2_u6_u1_U11 (.ZN( u2_u6_u1_n140 ) , .A2( u2_u6_u1_n150 ) , .A1( u2_u6_u1_n155 ) );
  NAND2_X1 u2_u6_u1_U12 (.A1( u2_u6_u1_n131 ) , .ZN( u2_u6_u1_n147 ) , .A2( u2_u6_u1_n153 ) );
  INV_X1 u2_u6_u1_U13 (.A( u2_u6_u1_n139 ) , .ZN( u2_u6_u1_n174 ) );
  OR4_X1 u2_u6_u1_U14 (.A4( u2_u6_u1_n106 ) , .A3( u2_u6_u1_n107 ) , .ZN( u2_u6_u1_n108 ) , .A1( u2_u6_u1_n117 ) , .A2( u2_u6_u1_n184 ) );
  AOI21_X1 u2_u6_u1_U15 (.ZN( u2_u6_u1_n106 ) , .A( u2_u6_u1_n112 ) , .B1( u2_u6_u1_n154 ) , .B2( u2_u6_u1_n156 ) );
  AOI21_X1 u2_u6_u1_U16 (.ZN( u2_u6_u1_n107 ) , .B1( u2_u6_u1_n134 ) , .B2( u2_u6_u1_n149 ) , .A( u2_u6_u1_n174 ) );
  INV_X1 u2_u6_u1_U17 (.A( u2_u6_u1_n101 ) , .ZN( u2_u6_u1_n184 ) );
  INV_X1 u2_u6_u1_U18 (.A( u2_u6_u1_n112 ) , .ZN( u2_u6_u1_n171 ) );
  NAND2_X1 u2_u6_u1_U19 (.ZN( u2_u6_u1_n141 ) , .A1( u2_u6_u1_n153 ) , .A2( u2_u6_u1_n156 ) );
  AND2_X1 u2_u6_u1_U20 (.A1( u2_u6_u1_n123 ) , .ZN( u2_u6_u1_n134 ) , .A2( u2_u6_u1_n161 ) );
  NAND2_X1 u2_u6_u1_U21 (.A2( u2_u6_u1_n115 ) , .A1( u2_u6_u1_n116 ) , .ZN( u2_u6_u1_n148 ) );
  NAND2_X1 u2_u6_u1_U22 (.A2( u2_u6_u1_n133 ) , .A1( u2_u6_u1_n135 ) , .ZN( u2_u6_u1_n159 ) );
  NAND2_X1 u2_u6_u1_U23 (.A2( u2_u6_u1_n115 ) , .A1( u2_u6_u1_n120 ) , .ZN( u2_u6_u1_n132 ) );
  INV_X1 u2_u6_u1_U24 (.A( u2_u6_u1_n154 ) , .ZN( u2_u6_u1_n178 ) );
  AOI22_X1 u2_u6_u1_U25 (.B2( u2_u6_u1_n113 ) , .A2( u2_u6_u1_n114 ) , .ZN( u2_u6_u1_n125 ) , .A1( u2_u6_u1_n171 ) , .B1( u2_u6_u1_n173 ) );
  NAND2_X1 u2_u6_u1_U26 (.ZN( u2_u6_u1_n114 ) , .A1( u2_u6_u1_n134 ) , .A2( u2_u6_u1_n156 ) );
  INV_X1 u2_u6_u1_U27 (.A( u2_u6_u1_n151 ) , .ZN( u2_u6_u1_n183 ) );
  AND2_X1 u2_u6_u1_U28 (.A1( u2_u6_u1_n129 ) , .A2( u2_u6_u1_n133 ) , .ZN( u2_u6_u1_n149 ) );
  INV_X1 u2_u6_u1_U29 (.A( u2_u6_u1_n131 ) , .ZN( u2_u6_u1_n180 ) );
  INV_X1 u2_u6_u1_U3 (.A( u2_u6_u1_n159 ) , .ZN( u2_u6_u1_n182 ) );
  AOI221_X1 u2_u6_u1_U30 (.B1( u2_u6_u1_n140 ) , .ZN( u2_u6_u1_n167 ) , .B2( u2_u6_u1_n172 ) , .C2( u2_u6_u1_n175 ) , .C1( u2_u6_u1_n178 ) , .A( u2_u6_u1_n188 ) );
  INV_X1 u2_u6_u1_U31 (.ZN( u2_u6_u1_n188 ) , .A( u2_u6_u1_n97 ) );
  AOI211_X1 u2_u6_u1_U32 (.A( u2_u6_u1_n118 ) , .C1( u2_u6_u1_n132 ) , .C2( u2_u6_u1_n139 ) , .B( u2_u6_u1_n96 ) , .ZN( u2_u6_u1_n97 ) );
  AOI21_X1 u2_u6_u1_U33 (.B2( u2_u6_u1_n121 ) , .B1( u2_u6_u1_n135 ) , .A( u2_u6_u1_n152 ) , .ZN( u2_u6_u1_n96 ) );
  OAI221_X1 u2_u6_u1_U34 (.A( u2_u6_u1_n119 ) , .C2( u2_u6_u1_n129 ) , .ZN( u2_u6_u1_n138 ) , .B2( u2_u6_u1_n152 ) , .C1( u2_u6_u1_n174 ) , .B1( u2_u6_u1_n187 ) );
  INV_X1 u2_u6_u1_U35 (.A( u2_u6_u1_n148 ) , .ZN( u2_u6_u1_n187 ) );
  AOI211_X1 u2_u6_u1_U36 (.B( u2_u6_u1_n117 ) , .A( u2_u6_u1_n118 ) , .ZN( u2_u6_u1_n119 ) , .C2( u2_u6_u1_n146 ) , .C1( u2_u6_u1_n159 ) );
  NOR2_X1 u2_u6_u1_U37 (.A1( u2_u6_u1_n168 ) , .A2( u2_u6_u1_n176 ) , .ZN( u2_u6_u1_n98 ) );
  AOI211_X1 u2_u6_u1_U38 (.B( u2_u6_u1_n162 ) , .A( u2_u6_u1_n163 ) , .C2( u2_u6_u1_n164 ) , .ZN( u2_u6_u1_n165 ) , .C1( u2_u6_u1_n171 ) );
  AOI21_X1 u2_u6_u1_U39 (.A( u2_u6_u1_n160 ) , .B2( u2_u6_u1_n161 ) , .ZN( u2_u6_u1_n162 ) , .B1( u2_u6_u1_n182 ) );
  AOI221_X1 u2_u6_u1_U4 (.A( u2_u6_u1_n138 ) , .C2( u2_u6_u1_n139 ) , .C1( u2_u6_u1_n140 ) , .B2( u2_u6_u1_n141 ) , .ZN( u2_u6_u1_n142 ) , .B1( u2_u6_u1_n175 ) );
  OR2_X1 u2_u6_u1_U40 (.A2( u2_u6_u1_n157 ) , .A1( u2_u6_u1_n158 ) , .ZN( u2_u6_u1_n163 ) );
  NAND2_X1 u2_u6_u1_U41 (.A1( u2_u6_u1_n128 ) , .ZN( u2_u6_u1_n146 ) , .A2( u2_u6_u1_n160 ) );
  NAND2_X1 u2_u6_u1_U42 (.A2( u2_u6_u1_n112 ) , .ZN( u2_u6_u1_n139 ) , .A1( u2_u6_u1_n152 ) );
  NAND2_X1 u2_u6_u1_U43 (.A1( u2_u6_u1_n105 ) , .ZN( u2_u6_u1_n156 ) , .A2( u2_u6_u1_n99 ) );
  NOR2_X1 u2_u6_u1_U44 (.ZN( u2_u6_u1_n117 ) , .A1( u2_u6_u1_n121 ) , .A2( u2_u6_u1_n160 ) );
  OAI21_X1 u2_u6_u1_U45 (.B2( u2_u6_u1_n123 ) , .ZN( u2_u6_u1_n145 ) , .B1( u2_u6_u1_n160 ) , .A( u2_u6_u1_n185 ) );
  INV_X1 u2_u6_u1_U46 (.A( u2_u6_u1_n122 ) , .ZN( u2_u6_u1_n185 ) );
  AOI21_X1 u2_u6_u1_U47 (.B2( u2_u6_u1_n120 ) , .B1( u2_u6_u1_n121 ) , .ZN( u2_u6_u1_n122 ) , .A( u2_u6_u1_n128 ) );
  AOI21_X1 u2_u6_u1_U48 (.A( u2_u6_u1_n128 ) , .B2( u2_u6_u1_n129 ) , .ZN( u2_u6_u1_n130 ) , .B1( u2_u6_u1_n150 ) );
  NAND2_X1 u2_u6_u1_U49 (.ZN( u2_u6_u1_n112 ) , .A1( u2_u6_u1_n169 ) , .A2( u2_u6_u1_n170 ) );
  AOI211_X1 u2_u6_u1_U5 (.ZN( u2_u6_u1_n124 ) , .A( u2_u6_u1_n138 ) , .C2( u2_u6_u1_n139 ) , .B( u2_u6_u1_n145 ) , .C1( u2_u6_u1_n147 ) );
  NAND2_X1 u2_u6_u1_U50 (.ZN( u2_u6_u1_n129 ) , .A2( u2_u6_u1_n95 ) , .A1( u2_u6_u1_n98 ) );
  NAND2_X1 u2_u6_u1_U51 (.A1( u2_u6_u1_n102 ) , .ZN( u2_u6_u1_n154 ) , .A2( u2_u6_u1_n99 ) );
  NAND2_X1 u2_u6_u1_U52 (.A2( u2_u6_u1_n100 ) , .ZN( u2_u6_u1_n135 ) , .A1( u2_u6_u1_n99 ) );
  AOI21_X1 u2_u6_u1_U53 (.A( u2_u6_u1_n152 ) , .B2( u2_u6_u1_n153 ) , .B1( u2_u6_u1_n154 ) , .ZN( u2_u6_u1_n158 ) );
  INV_X1 u2_u6_u1_U54 (.A( u2_u6_u1_n160 ) , .ZN( u2_u6_u1_n175 ) );
  NAND2_X1 u2_u6_u1_U55 (.A1( u2_u6_u1_n100 ) , .ZN( u2_u6_u1_n116 ) , .A2( u2_u6_u1_n95 ) );
  NAND2_X1 u2_u6_u1_U56 (.A1( u2_u6_u1_n102 ) , .ZN( u2_u6_u1_n131 ) , .A2( u2_u6_u1_n95 ) );
  NAND2_X1 u2_u6_u1_U57 (.A2( u2_u6_u1_n104 ) , .ZN( u2_u6_u1_n121 ) , .A1( u2_u6_u1_n98 ) );
  NAND2_X1 u2_u6_u1_U58 (.A1( u2_u6_u1_n103 ) , .ZN( u2_u6_u1_n153 ) , .A2( u2_u6_u1_n98 ) );
  NAND2_X1 u2_u6_u1_U59 (.A2( u2_u6_u1_n104 ) , .A1( u2_u6_u1_n105 ) , .ZN( u2_u6_u1_n133 ) );
  AOI22_X1 u2_u6_u1_U6 (.B2( u2_u6_u1_n136 ) , .A2( u2_u6_u1_n137 ) , .ZN( u2_u6_u1_n143 ) , .A1( u2_u6_u1_n171 ) , .B1( u2_u6_u1_n173 ) );
  NAND2_X1 u2_u6_u1_U60 (.ZN( u2_u6_u1_n150 ) , .A2( u2_u6_u1_n98 ) , .A1( u2_u6_u1_n99 ) );
  NAND2_X1 u2_u6_u1_U61 (.A1( u2_u6_u1_n105 ) , .ZN( u2_u6_u1_n155 ) , .A2( u2_u6_u1_n95 ) );
  OAI21_X1 u2_u6_u1_U62 (.ZN( u2_u6_u1_n109 ) , .B1( u2_u6_u1_n129 ) , .B2( u2_u6_u1_n160 ) , .A( u2_u6_u1_n167 ) );
  NAND2_X1 u2_u6_u1_U63 (.A2( u2_u6_u1_n100 ) , .A1( u2_u6_u1_n103 ) , .ZN( u2_u6_u1_n120 ) );
  NAND2_X1 u2_u6_u1_U64 (.A1( u2_u6_u1_n102 ) , .A2( u2_u6_u1_n104 ) , .ZN( u2_u6_u1_n115 ) );
  NAND2_X1 u2_u6_u1_U65 (.A2( u2_u6_u1_n100 ) , .A1( u2_u6_u1_n104 ) , .ZN( u2_u6_u1_n151 ) );
  NAND2_X1 u2_u6_u1_U66 (.A2( u2_u6_u1_n103 ) , .A1( u2_u6_u1_n105 ) , .ZN( u2_u6_u1_n161 ) );
  INV_X1 u2_u6_u1_U67 (.A( u2_u6_u1_n152 ) , .ZN( u2_u6_u1_n173 ) );
  INV_X1 u2_u6_u1_U68 (.A( u2_u6_u1_n128 ) , .ZN( u2_u6_u1_n172 ) );
  NAND2_X1 u2_u6_u1_U69 (.A2( u2_u6_u1_n102 ) , .A1( u2_u6_u1_n103 ) , .ZN( u2_u6_u1_n123 ) );
  INV_X1 u2_u6_u1_U7 (.A( u2_u6_u1_n147 ) , .ZN( u2_u6_u1_n181 ) );
  NOR2_X1 u2_u6_u1_U70 (.A2( u2_u6_X_7 ) , .A1( u2_u6_X_8 ) , .ZN( u2_u6_u1_n95 ) );
  NOR2_X1 u2_u6_u1_U71 (.A1( u2_u6_X_12 ) , .A2( u2_u6_X_9 ) , .ZN( u2_u6_u1_n100 ) );
  NOR2_X1 u2_u6_u1_U72 (.A2( u2_u6_X_8 ) , .A1( u2_u6_u1_n177 ) , .ZN( u2_u6_u1_n99 ) );
  NOR2_X1 u2_u6_u1_U73 (.A2( u2_u6_X_12 ) , .ZN( u2_u6_u1_n102 ) , .A1( u2_u6_u1_n176 ) );
  NOR2_X1 u2_u6_u1_U74 (.A2( u2_u6_X_9 ) , .ZN( u2_u6_u1_n105 ) , .A1( u2_u6_u1_n168 ) );
  NAND2_X1 u2_u6_u1_U75 (.A1( u2_u6_X_10 ) , .ZN( u2_u6_u1_n160 ) , .A2( u2_u6_u1_n169 ) );
  NAND2_X1 u2_u6_u1_U76 (.A2( u2_u6_X_10 ) , .A1( u2_u6_X_11 ) , .ZN( u2_u6_u1_n152 ) );
  NAND2_X1 u2_u6_u1_U77 (.A1( u2_u6_X_11 ) , .ZN( u2_u6_u1_n128 ) , .A2( u2_u6_u1_n170 ) );
  AND2_X1 u2_u6_u1_U78 (.A2( u2_u6_X_7 ) , .A1( u2_u6_X_8 ) , .ZN( u2_u6_u1_n104 ) );
  AND2_X1 u2_u6_u1_U79 (.A1( u2_u6_X_8 ) , .ZN( u2_u6_u1_n103 ) , .A2( u2_u6_u1_n177 ) );
  NOR2_X1 u2_u6_u1_U8 (.A1( u2_u6_u1_n112 ) , .A2( u2_u6_u1_n116 ) , .ZN( u2_u6_u1_n118 ) );
  INV_X1 u2_u6_u1_U80 (.A( u2_u6_X_10 ) , .ZN( u2_u6_u1_n170 ) );
  INV_X1 u2_u6_u1_U81 (.A( u2_u6_X_9 ) , .ZN( u2_u6_u1_n176 ) );
  INV_X1 u2_u6_u1_U82 (.A( u2_u6_X_11 ) , .ZN( u2_u6_u1_n169 ) );
  INV_X1 u2_u6_u1_U83 (.A( u2_u6_X_12 ) , .ZN( u2_u6_u1_n168 ) );
  INV_X1 u2_u6_u1_U84 (.A( u2_u6_X_7 ) , .ZN( u2_u6_u1_n177 ) );
  NAND4_X1 u2_u6_u1_U85 (.ZN( u2_out6_28 ) , .A4( u2_u6_u1_n124 ) , .A3( u2_u6_u1_n125 ) , .A2( u2_u6_u1_n126 ) , .A1( u2_u6_u1_n127 ) );
  OAI21_X1 u2_u6_u1_U86 (.ZN( u2_u6_u1_n127 ) , .B2( u2_u6_u1_n139 ) , .B1( u2_u6_u1_n175 ) , .A( u2_u6_u1_n183 ) );
  OAI21_X1 u2_u6_u1_U87 (.ZN( u2_u6_u1_n126 ) , .B2( u2_u6_u1_n140 ) , .A( u2_u6_u1_n146 ) , .B1( u2_u6_u1_n178 ) );
  NAND4_X1 u2_u6_u1_U88 (.ZN( u2_out6_18 ) , .A4( u2_u6_u1_n165 ) , .A3( u2_u6_u1_n166 ) , .A1( u2_u6_u1_n167 ) , .A2( u2_u6_u1_n186 ) );
  AOI22_X1 u2_u6_u1_U89 (.B2( u2_u6_u1_n146 ) , .B1( u2_u6_u1_n147 ) , .A2( u2_u6_u1_n148 ) , .ZN( u2_u6_u1_n166 ) , .A1( u2_u6_u1_n172 ) );
  OAI21_X1 u2_u6_u1_U9 (.ZN( u2_u6_u1_n101 ) , .B1( u2_u6_u1_n141 ) , .A( u2_u6_u1_n146 ) , .B2( u2_u6_u1_n183 ) );
  INV_X1 u2_u6_u1_U90 (.A( u2_u6_u1_n145 ) , .ZN( u2_u6_u1_n186 ) );
  NAND4_X1 u2_u6_u1_U91 (.ZN( u2_out6_2 ) , .A4( u2_u6_u1_n142 ) , .A3( u2_u6_u1_n143 ) , .A2( u2_u6_u1_n144 ) , .A1( u2_u6_u1_n179 ) );
  OAI21_X1 u2_u6_u1_U92 (.B2( u2_u6_u1_n132 ) , .ZN( u2_u6_u1_n144 ) , .A( u2_u6_u1_n146 ) , .B1( u2_u6_u1_n180 ) );
  INV_X1 u2_u6_u1_U93 (.A( u2_u6_u1_n130 ) , .ZN( u2_u6_u1_n179 ) );
  OR4_X1 u2_u6_u1_U94 (.ZN( u2_out6_13 ) , .A4( u2_u6_u1_n108 ) , .A3( u2_u6_u1_n109 ) , .A2( u2_u6_u1_n110 ) , .A1( u2_u6_u1_n111 ) );
  AOI21_X1 u2_u6_u1_U95 (.ZN( u2_u6_u1_n111 ) , .A( u2_u6_u1_n128 ) , .B2( u2_u6_u1_n131 ) , .B1( u2_u6_u1_n135 ) );
  AOI21_X1 u2_u6_u1_U96 (.ZN( u2_u6_u1_n110 ) , .A( u2_u6_u1_n116 ) , .B1( u2_u6_u1_n152 ) , .B2( u2_u6_u1_n160 ) );
  NAND3_X1 u2_u6_u1_U97 (.A3( u2_u6_u1_n149 ) , .A2( u2_u6_u1_n150 ) , .A1( u2_u6_u1_n151 ) , .ZN( u2_u6_u1_n164 ) );
  NAND3_X1 u2_u6_u1_U98 (.A3( u2_u6_u1_n134 ) , .A2( u2_u6_u1_n135 ) , .ZN( u2_u6_u1_n136 ) , .A1( u2_u6_u1_n151 ) );
  NAND3_X1 u2_u6_u1_U99 (.A1( u2_u6_u1_n133 ) , .ZN( u2_u6_u1_n137 ) , .A2( u2_u6_u1_n154 ) , .A3( u2_u6_u1_n181 ) );
  OAI22_X1 u2_u6_u2_U10 (.B1( u2_u6_u2_n151 ) , .A2( u2_u6_u2_n152 ) , .A1( u2_u6_u2_n153 ) , .ZN( u2_u6_u2_n160 ) , .B2( u2_u6_u2_n168 ) );
  NAND3_X1 u2_u6_u2_U100 (.A2( u2_u6_u2_n100 ) , .A1( u2_u6_u2_n104 ) , .A3( u2_u6_u2_n138 ) , .ZN( u2_u6_u2_n98 ) );
  NOR3_X1 u2_u6_u2_U11 (.A1( u2_u6_u2_n150 ) , .ZN( u2_u6_u2_n151 ) , .A3( u2_u6_u2_n175 ) , .A2( u2_u6_u2_n188 ) );
  AOI21_X1 u2_u6_u2_U12 (.B2( u2_u6_u2_n123 ) , .ZN( u2_u6_u2_n125 ) , .A( u2_u6_u2_n171 ) , .B1( u2_u6_u2_n184 ) );
  INV_X1 u2_u6_u2_U13 (.A( u2_u6_u2_n150 ) , .ZN( u2_u6_u2_n184 ) );
  AOI21_X1 u2_u6_u2_U14 (.ZN( u2_u6_u2_n144 ) , .B2( u2_u6_u2_n155 ) , .A( u2_u6_u2_n172 ) , .B1( u2_u6_u2_n185 ) );
  AOI21_X1 u2_u6_u2_U15 (.B2( u2_u6_u2_n143 ) , .ZN( u2_u6_u2_n145 ) , .B1( u2_u6_u2_n152 ) , .A( u2_u6_u2_n171 ) );
  INV_X1 u2_u6_u2_U16 (.A( u2_u6_u2_n156 ) , .ZN( u2_u6_u2_n171 ) );
  INV_X1 u2_u6_u2_U17 (.A( u2_u6_u2_n120 ) , .ZN( u2_u6_u2_n188 ) );
  NAND2_X1 u2_u6_u2_U18 (.A2( u2_u6_u2_n122 ) , .ZN( u2_u6_u2_n150 ) , .A1( u2_u6_u2_n152 ) );
  INV_X1 u2_u6_u2_U19 (.A( u2_u6_u2_n153 ) , .ZN( u2_u6_u2_n170 ) );
  INV_X1 u2_u6_u2_U20 (.A( u2_u6_u2_n137 ) , .ZN( u2_u6_u2_n173 ) );
  NAND2_X1 u2_u6_u2_U21 (.A1( u2_u6_u2_n132 ) , .A2( u2_u6_u2_n139 ) , .ZN( u2_u6_u2_n157 ) );
  INV_X1 u2_u6_u2_U22 (.A( u2_u6_u2_n113 ) , .ZN( u2_u6_u2_n178 ) );
  INV_X1 u2_u6_u2_U23 (.A( u2_u6_u2_n139 ) , .ZN( u2_u6_u2_n175 ) );
  INV_X1 u2_u6_u2_U24 (.A( u2_u6_u2_n155 ) , .ZN( u2_u6_u2_n181 ) );
  INV_X1 u2_u6_u2_U25 (.A( u2_u6_u2_n119 ) , .ZN( u2_u6_u2_n177 ) );
  INV_X1 u2_u6_u2_U26 (.A( u2_u6_u2_n116 ) , .ZN( u2_u6_u2_n180 ) );
  INV_X1 u2_u6_u2_U27 (.A( u2_u6_u2_n131 ) , .ZN( u2_u6_u2_n179 ) );
  INV_X1 u2_u6_u2_U28 (.A( u2_u6_u2_n154 ) , .ZN( u2_u6_u2_n176 ) );
  NAND2_X1 u2_u6_u2_U29 (.A2( u2_u6_u2_n116 ) , .A1( u2_u6_u2_n117 ) , .ZN( u2_u6_u2_n118 ) );
  NOR2_X1 u2_u6_u2_U3 (.ZN( u2_u6_u2_n121 ) , .A2( u2_u6_u2_n177 ) , .A1( u2_u6_u2_n180 ) );
  INV_X1 u2_u6_u2_U30 (.A( u2_u6_u2_n132 ) , .ZN( u2_u6_u2_n182 ) );
  INV_X1 u2_u6_u2_U31 (.A( u2_u6_u2_n158 ) , .ZN( u2_u6_u2_n183 ) );
  OAI21_X1 u2_u6_u2_U32 (.A( u2_u6_u2_n156 ) , .B1( u2_u6_u2_n157 ) , .ZN( u2_u6_u2_n158 ) , .B2( u2_u6_u2_n179 ) );
  NOR2_X1 u2_u6_u2_U33 (.ZN( u2_u6_u2_n156 ) , .A1( u2_u6_u2_n166 ) , .A2( u2_u6_u2_n169 ) );
  NOR2_X1 u2_u6_u2_U34 (.A2( u2_u6_u2_n114 ) , .ZN( u2_u6_u2_n137 ) , .A1( u2_u6_u2_n140 ) );
  NOR2_X1 u2_u6_u2_U35 (.A2( u2_u6_u2_n138 ) , .ZN( u2_u6_u2_n153 ) , .A1( u2_u6_u2_n156 ) );
  AOI211_X1 u2_u6_u2_U36 (.ZN( u2_u6_u2_n130 ) , .C1( u2_u6_u2_n138 ) , .C2( u2_u6_u2_n179 ) , .B( u2_u6_u2_n96 ) , .A( u2_u6_u2_n97 ) );
  OAI22_X1 u2_u6_u2_U37 (.B1( u2_u6_u2_n133 ) , .A2( u2_u6_u2_n137 ) , .A1( u2_u6_u2_n152 ) , .B2( u2_u6_u2_n168 ) , .ZN( u2_u6_u2_n97 ) );
  OAI221_X1 u2_u6_u2_U38 (.B1( u2_u6_u2_n113 ) , .C1( u2_u6_u2_n132 ) , .A( u2_u6_u2_n149 ) , .B2( u2_u6_u2_n171 ) , .C2( u2_u6_u2_n172 ) , .ZN( u2_u6_u2_n96 ) );
  OAI221_X1 u2_u6_u2_U39 (.A( u2_u6_u2_n115 ) , .C2( u2_u6_u2_n123 ) , .B2( u2_u6_u2_n143 ) , .B1( u2_u6_u2_n153 ) , .ZN( u2_u6_u2_n163 ) , .C1( u2_u6_u2_n168 ) );
  INV_X1 u2_u6_u2_U4 (.A( u2_u6_u2_n134 ) , .ZN( u2_u6_u2_n185 ) );
  OAI21_X1 u2_u6_u2_U40 (.A( u2_u6_u2_n114 ) , .ZN( u2_u6_u2_n115 ) , .B1( u2_u6_u2_n176 ) , .B2( u2_u6_u2_n178 ) );
  OAI221_X1 u2_u6_u2_U41 (.A( u2_u6_u2_n135 ) , .B2( u2_u6_u2_n136 ) , .B1( u2_u6_u2_n137 ) , .ZN( u2_u6_u2_n162 ) , .C2( u2_u6_u2_n167 ) , .C1( u2_u6_u2_n185 ) );
  AND3_X1 u2_u6_u2_U42 (.A3( u2_u6_u2_n131 ) , .A2( u2_u6_u2_n132 ) , .A1( u2_u6_u2_n133 ) , .ZN( u2_u6_u2_n136 ) );
  AOI22_X1 u2_u6_u2_U43 (.ZN( u2_u6_u2_n135 ) , .B1( u2_u6_u2_n140 ) , .A1( u2_u6_u2_n156 ) , .B2( u2_u6_u2_n180 ) , .A2( u2_u6_u2_n188 ) );
  AOI21_X1 u2_u6_u2_U44 (.ZN( u2_u6_u2_n149 ) , .B1( u2_u6_u2_n173 ) , .B2( u2_u6_u2_n188 ) , .A( u2_u6_u2_n95 ) );
  AND3_X1 u2_u6_u2_U45 (.A2( u2_u6_u2_n100 ) , .A1( u2_u6_u2_n104 ) , .A3( u2_u6_u2_n156 ) , .ZN( u2_u6_u2_n95 ) );
  OAI21_X1 u2_u6_u2_U46 (.A( u2_u6_u2_n141 ) , .B2( u2_u6_u2_n142 ) , .ZN( u2_u6_u2_n146 ) , .B1( u2_u6_u2_n153 ) );
  OAI21_X1 u2_u6_u2_U47 (.A( u2_u6_u2_n140 ) , .ZN( u2_u6_u2_n141 ) , .B1( u2_u6_u2_n176 ) , .B2( u2_u6_u2_n177 ) );
  NOR3_X1 u2_u6_u2_U48 (.ZN( u2_u6_u2_n142 ) , .A3( u2_u6_u2_n175 ) , .A2( u2_u6_u2_n178 ) , .A1( u2_u6_u2_n181 ) );
  OAI21_X1 u2_u6_u2_U49 (.A( u2_u6_u2_n101 ) , .B2( u2_u6_u2_n121 ) , .B1( u2_u6_u2_n153 ) , .ZN( u2_u6_u2_n164 ) );
  NOR4_X1 u2_u6_u2_U5 (.A4( u2_u6_u2_n124 ) , .A3( u2_u6_u2_n125 ) , .A2( u2_u6_u2_n126 ) , .A1( u2_u6_u2_n127 ) , .ZN( u2_u6_u2_n128 ) );
  NAND2_X1 u2_u6_u2_U50 (.A2( u2_u6_u2_n100 ) , .A1( u2_u6_u2_n107 ) , .ZN( u2_u6_u2_n155 ) );
  NAND2_X1 u2_u6_u2_U51 (.A2( u2_u6_u2_n105 ) , .A1( u2_u6_u2_n108 ) , .ZN( u2_u6_u2_n143 ) );
  NAND2_X1 u2_u6_u2_U52 (.A1( u2_u6_u2_n104 ) , .A2( u2_u6_u2_n106 ) , .ZN( u2_u6_u2_n152 ) );
  NAND2_X1 u2_u6_u2_U53 (.A1( u2_u6_u2_n100 ) , .A2( u2_u6_u2_n105 ) , .ZN( u2_u6_u2_n132 ) );
  INV_X1 u2_u6_u2_U54 (.A( u2_u6_u2_n140 ) , .ZN( u2_u6_u2_n168 ) );
  INV_X1 u2_u6_u2_U55 (.A( u2_u6_u2_n138 ) , .ZN( u2_u6_u2_n167 ) );
  INV_X1 u2_u6_u2_U56 (.ZN( u2_u6_u2_n187 ) , .A( u2_u6_u2_n99 ) );
  OAI21_X1 u2_u6_u2_U57 (.B1( u2_u6_u2_n137 ) , .B2( u2_u6_u2_n143 ) , .A( u2_u6_u2_n98 ) , .ZN( u2_u6_u2_n99 ) );
  NAND2_X1 u2_u6_u2_U58 (.A1( u2_u6_u2_n102 ) , .A2( u2_u6_u2_n106 ) , .ZN( u2_u6_u2_n113 ) );
  NAND2_X1 u2_u6_u2_U59 (.A1( u2_u6_u2_n106 ) , .A2( u2_u6_u2_n107 ) , .ZN( u2_u6_u2_n131 ) );
  AOI21_X1 u2_u6_u2_U6 (.B2( u2_u6_u2_n119 ) , .ZN( u2_u6_u2_n127 ) , .A( u2_u6_u2_n137 ) , .B1( u2_u6_u2_n155 ) );
  NAND2_X1 u2_u6_u2_U60 (.A1( u2_u6_u2_n103 ) , .A2( u2_u6_u2_n107 ) , .ZN( u2_u6_u2_n139 ) );
  NAND2_X1 u2_u6_u2_U61 (.A1( u2_u6_u2_n103 ) , .A2( u2_u6_u2_n105 ) , .ZN( u2_u6_u2_n133 ) );
  NAND2_X1 u2_u6_u2_U62 (.A1( u2_u6_u2_n102 ) , .A2( u2_u6_u2_n103 ) , .ZN( u2_u6_u2_n154 ) );
  NAND2_X1 u2_u6_u2_U63 (.A2( u2_u6_u2_n103 ) , .A1( u2_u6_u2_n104 ) , .ZN( u2_u6_u2_n119 ) );
  NAND2_X1 u2_u6_u2_U64 (.A2( u2_u6_u2_n107 ) , .A1( u2_u6_u2_n108 ) , .ZN( u2_u6_u2_n123 ) );
  NAND2_X1 u2_u6_u2_U65 (.A1( u2_u6_u2_n104 ) , .A2( u2_u6_u2_n108 ) , .ZN( u2_u6_u2_n122 ) );
  INV_X1 u2_u6_u2_U66 (.A( u2_u6_u2_n114 ) , .ZN( u2_u6_u2_n172 ) );
  NAND2_X1 u2_u6_u2_U67 (.A2( u2_u6_u2_n100 ) , .A1( u2_u6_u2_n102 ) , .ZN( u2_u6_u2_n116 ) );
  NAND2_X1 u2_u6_u2_U68 (.A1( u2_u6_u2_n102 ) , .A2( u2_u6_u2_n108 ) , .ZN( u2_u6_u2_n120 ) );
  NAND2_X1 u2_u6_u2_U69 (.A2( u2_u6_u2_n105 ) , .A1( u2_u6_u2_n106 ) , .ZN( u2_u6_u2_n117 ) );
  AOI21_X1 u2_u6_u2_U7 (.ZN( u2_u6_u2_n124 ) , .B1( u2_u6_u2_n131 ) , .B2( u2_u6_u2_n143 ) , .A( u2_u6_u2_n172 ) );
  NOR2_X1 u2_u6_u2_U70 (.A2( u2_u6_X_16 ) , .ZN( u2_u6_u2_n140 ) , .A1( u2_u6_u2_n166 ) );
  NOR2_X1 u2_u6_u2_U71 (.A2( u2_u6_X_13 ) , .A1( u2_u6_X_14 ) , .ZN( u2_u6_u2_n100 ) );
  NOR2_X1 u2_u6_u2_U72 (.A2( u2_u6_X_16 ) , .A1( u2_u6_X_17 ) , .ZN( u2_u6_u2_n138 ) );
  NOR2_X1 u2_u6_u2_U73 (.A2( u2_u6_X_15 ) , .A1( u2_u6_X_18 ) , .ZN( u2_u6_u2_n104 ) );
  NOR2_X1 u2_u6_u2_U74 (.A2( u2_u6_X_14 ) , .ZN( u2_u6_u2_n103 ) , .A1( u2_u6_u2_n174 ) );
  NOR2_X1 u2_u6_u2_U75 (.A2( u2_u6_X_15 ) , .ZN( u2_u6_u2_n102 ) , .A1( u2_u6_u2_n165 ) );
  NOR2_X1 u2_u6_u2_U76 (.A2( u2_u6_X_17 ) , .ZN( u2_u6_u2_n114 ) , .A1( u2_u6_u2_n169 ) );
  AND2_X1 u2_u6_u2_U77 (.A1( u2_u6_X_15 ) , .ZN( u2_u6_u2_n105 ) , .A2( u2_u6_u2_n165 ) );
  AND2_X1 u2_u6_u2_U78 (.A2( u2_u6_X_15 ) , .A1( u2_u6_X_18 ) , .ZN( u2_u6_u2_n107 ) );
  AND2_X1 u2_u6_u2_U79 (.A1( u2_u6_X_14 ) , .ZN( u2_u6_u2_n106 ) , .A2( u2_u6_u2_n174 ) );
  AOI21_X1 u2_u6_u2_U8 (.B2( u2_u6_u2_n120 ) , .B1( u2_u6_u2_n121 ) , .ZN( u2_u6_u2_n126 ) , .A( u2_u6_u2_n167 ) );
  AND2_X1 u2_u6_u2_U80 (.A1( u2_u6_X_13 ) , .A2( u2_u6_X_14 ) , .ZN( u2_u6_u2_n108 ) );
  INV_X1 u2_u6_u2_U81 (.A( u2_u6_X_16 ) , .ZN( u2_u6_u2_n169 ) );
  INV_X1 u2_u6_u2_U82 (.A( u2_u6_X_17 ) , .ZN( u2_u6_u2_n166 ) );
  INV_X1 u2_u6_u2_U83 (.A( u2_u6_X_13 ) , .ZN( u2_u6_u2_n174 ) );
  INV_X1 u2_u6_u2_U84 (.A( u2_u6_X_18 ) , .ZN( u2_u6_u2_n165 ) );
  NAND4_X1 u2_u6_u2_U85 (.ZN( u2_out6_30 ) , .A4( u2_u6_u2_n147 ) , .A3( u2_u6_u2_n148 ) , .A2( u2_u6_u2_n149 ) , .A1( u2_u6_u2_n187 ) );
  AOI21_X1 u2_u6_u2_U86 (.B2( u2_u6_u2_n138 ) , .ZN( u2_u6_u2_n148 ) , .A( u2_u6_u2_n162 ) , .B1( u2_u6_u2_n182 ) );
  NOR3_X1 u2_u6_u2_U87 (.A3( u2_u6_u2_n144 ) , .A2( u2_u6_u2_n145 ) , .A1( u2_u6_u2_n146 ) , .ZN( u2_u6_u2_n147 ) );
  NAND4_X1 u2_u6_u2_U88 (.ZN( u2_out6_24 ) , .A4( u2_u6_u2_n111 ) , .A3( u2_u6_u2_n112 ) , .A1( u2_u6_u2_n130 ) , .A2( u2_u6_u2_n187 ) );
  AOI221_X1 u2_u6_u2_U89 (.A( u2_u6_u2_n109 ) , .B1( u2_u6_u2_n110 ) , .ZN( u2_u6_u2_n111 ) , .C1( u2_u6_u2_n134 ) , .C2( u2_u6_u2_n170 ) , .B2( u2_u6_u2_n173 ) );
  OAI22_X1 u2_u6_u2_U9 (.ZN( u2_u6_u2_n109 ) , .A2( u2_u6_u2_n113 ) , .B2( u2_u6_u2_n133 ) , .B1( u2_u6_u2_n167 ) , .A1( u2_u6_u2_n168 ) );
  AOI21_X1 u2_u6_u2_U90 (.ZN( u2_u6_u2_n112 ) , .B2( u2_u6_u2_n156 ) , .A( u2_u6_u2_n164 ) , .B1( u2_u6_u2_n181 ) );
  NAND4_X1 u2_u6_u2_U91 (.ZN( u2_out6_16 ) , .A4( u2_u6_u2_n128 ) , .A3( u2_u6_u2_n129 ) , .A1( u2_u6_u2_n130 ) , .A2( u2_u6_u2_n186 ) );
  AOI22_X1 u2_u6_u2_U92 (.A2( u2_u6_u2_n118 ) , .ZN( u2_u6_u2_n129 ) , .A1( u2_u6_u2_n140 ) , .B1( u2_u6_u2_n157 ) , .B2( u2_u6_u2_n170 ) );
  INV_X1 u2_u6_u2_U93 (.A( u2_u6_u2_n163 ) , .ZN( u2_u6_u2_n186 ) );
  OR4_X1 u2_u6_u2_U94 (.ZN( u2_out6_6 ) , .A4( u2_u6_u2_n161 ) , .A3( u2_u6_u2_n162 ) , .A2( u2_u6_u2_n163 ) , .A1( u2_u6_u2_n164 ) );
  OR3_X1 u2_u6_u2_U95 (.A2( u2_u6_u2_n159 ) , .A1( u2_u6_u2_n160 ) , .ZN( u2_u6_u2_n161 ) , .A3( u2_u6_u2_n183 ) );
  AOI21_X1 u2_u6_u2_U96 (.B2( u2_u6_u2_n154 ) , .B1( u2_u6_u2_n155 ) , .ZN( u2_u6_u2_n159 ) , .A( u2_u6_u2_n167 ) );
  NAND3_X1 u2_u6_u2_U97 (.A2( u2_u6_u2_n117 ) , .A1( u2_u6_u2_n122 ) , .A3( u2_u6_u2_n123 ) , .ZN( u2_u6_u2_n134 ) );
  NAND3_X1 u2_u6_u2_U98 (.ZN( u2_u6_u2_n110 ) , .A2( u2_u6_u2_n131 ) , .A3( u2_u6_u2_n139 ) , .A1( u2_u6_u2_n154 ) );
  NAND3_X1 u2_u6_u2_U99 (.A2( u2_u6_u2_n100 ) , .ZN( u2_u6_u2_n101 ) , .A1( u2_u6_u2_n104 ) , .A3( u2_u6_u2_n114 ) );
  OAI22_X1 u2_u6_u3_U10 (.B1( u2_u6_u3_n113 ) , .A2( u2_u6_u3_n135 ) , .A1( u2_u6_u3_n150 ) , .B2( u2_u6_u3_n164 ) , .ZN( u2_u6_u3_n98 ) );
  OAI211_X1 u2_u6_u3_U11 (.B( u2_u6_u3_n106 ) , .ZN( u2_u6_u3_n119 ) , .C2( u2_u6_u3_n128 ) , .C1( u2_u6_u3_n167 ) , .A( u2_u6_u3_n181 ) );
  AOI221_X1 u2_u6_u3_U12 (.C1( u2_u6_u3_n105 ) , .ZN( u2_u6_u3_n106 ) , .A( u2_u6_u3_n131 ) , .B2( u2_u6_u3_n132 ) , .C2( u2_u6_u3_n133 ) , .B1( u2_u6_u3_n169 ) );
  INV_X1 u2_u6_u3_U13 (.ZN( u2_u6_u3_n181 ) , .A( u2_u6_u3_n98 ) );
  NAND2_X1 u2_u6_u3_U14 (.ZN( u2_u6_u3_n105 ) , .A2( u2_u6_u3_n130 ) , .A1( u2_u6_u3_n155 ) );
  NOR2_X1 u2_u6_u3_U15 (.ZN( u2_u6_u3_n126 ) , .A2( u2_u6_u3_n150 ) , .A1( u2_u6_u3_n164 ) );
  AOI21_X1 u2_u6_u3_U16 (.ZN( u2_u6_u3_n112 ) , .B2( u2_u6_u3_n146 ) , .B1( u2_u6_u3_n155 ) , .A( u2_u6_u3_n167 ) );
  NAND2_X1 u2_u6_u3_U17 (.A1( u2_u6_u3_n135 ) , .ZN( u2_u6_u3_n142 ) , .A2( u2_u6_u3_n164 ) );
  NAND2_X1 u2_u6_u3_U18 (.ZN( u2_u6_u3_n132 ) , .A2( u2_u6_u3_n152 ) , .A1( u2_u6_u3_n156 ) );
  AND2_X1 u2_u6_u3_U19 (.A2( u2_u6_u3_n113 ) , .A1( u2_u6_u3_n114 ) , .ZN( u2_u6_u3_n151 ) );
  INV_X1 u2_u6_u3_U20 (.A( u2_u6_u3_n133 ) , .ZN( u2_u6_u3_n165 ) );
  INV_X1 u2_u6_u3_U21 (.A( u2_u6_u3_n135 ) , .ZN( u2_u6_u3_n170 ) );
  NAND2_X1 u2_u6_u3_U22 (.A1( u2_u6_u3_n107 ) , .A2( u2_u6_u3_n108 ) , .ZN( u2_u6_u3_n140 ) );
  NAND2_X1 u2_u6_u3_U23 (.ZN( u2_u6_u3_n117 ) , .A1( u2_u6_u3_n124 ) , .A2( u2_u6_u3_n148 ) );
  NAND2_X1 u2_u6_u3_U24 (.ZN( u2_u6_u3_n143 ) , .A1( u2_u6_u3_n165 ) , .A2( u2_u6_u3_n167 ) );
  INV_X1 u2_u6_u3_U25 (.A( u2_u6_u3_n130 ) , .ZN( u2_u6_u3_n177 ) );
  INV_X1 u2_u6_u3_U26 (.A( u2_u6_u3_n128 ) , .ZN( u2_u6_u3_n176 ) );
  INV_X1 u2_u6_u3_U27 (.A( u2_u6_u3_n155 ) , .ZN( u2_u6_u3_n174 ) );
  AOI22_X1 u2_u6_u3_U28 (.B1( u2_u6_u3_n115 ) , .A2( u2_u6_u3_n116 ) , .ZN( u2_u6_u3_n123 ) , .B2( u2_u6_u3_n133 ) , .A1( u2_u6_u3_n169 ) );
  NAND2_X1 u2_u6_u3_U29 (.ZN( u2_u6_u3_n116 ) , .A2( u2_u6_u3_n151 ) , .A1( u2_u6_u3_n182 ) );
  INV_X1 u2_u6_u3_U3 (.A( u2_u6_u3_n129 ) , .ZN( u2_u6_u3_n183 ) );
  INV_X1 u2_u6_u3_U30 (.A( u2_u6_u3_n139 ) , .ZN( u2_u6_u3_n185 ) );
  NOR2_X1 u2_u6_u3_U31 (.ZN( u2_u6_u3_n135 ) , .A2( u2_u6_u3_n141 ) , .A1( u2_u6_u3_n169 ) );
  OAI222_X1 u2_u6_u3_U32 (.C2( u2_u6_u3_n107 ) , .A2( u2_u6_u3_n108 ) , .B1( u2_u6_u3_n135 ) , .ZN( u2_u6_u3_n138 ) , .B2( u2_u6_u3_n146 ) , .C1( u2_u6_u3_n154 ) , .A1( u2_u6_u3_n164 ) );
  NOR4_X1 u2_u6_u3_U33 (.A4( u2_u6_u3_n157 ) , .A3( u2_u6_u3_n158 ) , .A2( u2_u6_u3_n159 ) , .A1( u2_u6_u3_n160 ) , .ZN( u2_u6_u3_n161 ) );
  AOI21_X1 u2_u6_u3_U34 (.B2( u2_u6_u3_n152 ) , .B1( u2_u6_u3_n153 ) , .ZN( u2_u6_u3_n158 ) , .A( u2_u6_u3_n164 ) );
  AOI21_X1 u2_u6_u3_U35 (.A( u2_u6_u3_n154 ) , .B2( u2_u6_u3_n155 ) , .B1( u2_u6_u3_n156 ) , .ZN( u2_u6_u3_n157 ) );
  AOI21_X1 u2_u6_u3_U36 (.A( u2_u6_u3_n149 ) , .B2( u2_u6_u3_n150 ) , .B1( u2_u6_u3_n151 ) , .ZN( u2_u6_u3_n159 ) );
  AOI211_X1 u2_u6_u3_U37 (.ZN( u2_u6_u3_n109 ) , .A( u2_u6_u3_n119 ) , .C2( u2_u6_u3_n129 ) , .B( u2_u6_u3_n138 ) , .C1( u2_u6_u3_n141 ) );
  AOI211_X1 u2_u6_u3_U38 (.B( u2_u6_u3_n119 ) , .A( u2_u6_u3_n120 ) , .C2( u2_u6_u3_n121 ) , .ZN( u2_u6_u3_n122 ) , .C1( u2_u6_u3_n179 ) );
  INV_X1 u2_u6_u3_U39 (.A( u2_u6_u3_n156 ) , .ZN( u2_u6_u3_n179 ) );
  INV_X1 u2_u6_u3_U4 (.A( u2_u6_u3_n140 ) , .ZN( u2_u6_u3_n182 ) );
  OAI22_X1 u2_u6_u3_U40 (.B1( u2_u6_u3_n118 ) , .ZN( u2_u6_u3_n120 ) , .A1( u2_u6_u3_n135 ) , .B2( u2_u6_u3_n154 ) , .A2( u2_u6_u3_n178 ) );
  AND3_X1 u2_u6_u3_U41 (.ZN( u2_u6_u3_n118 ) , .A2( u2_u6_u3_n124 ) , .A1( u2_u6_u3_n144 ) , .A3( u2_u6_u3_n152 ) );
  INV_X1 u2_u6_u3_U42 (.A( u2_u6_u3_n121 ) , .ZN( u2_u6_u3_n164 ) );
  NAND2_X1 u2_u6_u3_U43 (.ZN( u2_u6_u3_n133 ) , .A1( u2_u6_u3_n154 ) , .A2( u2_u6_u3_n164 ) );
  OAI211_X1 u2_u6_u3_U44 (.B( u2_u6_u3_n127 ) , .ZN( u2_u6_u3_n139 ) , .C1( u2_u6_u3_n150 ) , .C2( u2_u6_u3_n154 ) , .A( u2_u6_u3_n184 ) );
  INV_X1 u2_u6_u3_U45 (.A( u2_u6_u3_n125 ) , .ZN( u2_u6_u3_n184 ) );
  AOI221_X1 u2_u6_u3_U46 (.A( u2_u6_u3_n126 ) , .ZN( u2_u6_u3_n127 ) , .C2( u2_u6_u3_n132 ) , .C1( u2_u6_u3_n169 ) , .B2( u2_u6_u3_n170 ) , .B1( u2_u6_u3_n174 ) );
  OAI22_X1 u2_u6_u3_U47 (.A1( u2_u6_u3_n124 ) , .ZN( u2_u6_u3_n125 ) , .B2( u2_u6_u3_n145 ) , .A2( u2_u6_u3_n165 ) , .B1( u2_u6_u3_n167 ) );
  NOR2_X1 u2_u6_u3_U48 (.A1( u2_u6_u3_n113 ) , .ZN( u2_u6_u3_n131 ) , .A2( u2_u6_u3_n154 ) );
  NAND2_X1 u2_u6_u3_U49 (.A1( u2_u6_u3_n103 ) , .ZN( u2_u6_u3_n150 ) , .A2( u2_u6_u3_n99 ) );
  INV_X1 u2_u6_u3_U5 (.A( u2_u6_u3_n117 ) , .ZN( u2_u6_u3_n178 ) );
  NAND2_X1 u2_u6_u3_U50 (.A2( u2_u6_u3_n102 ) , .ZN( u2_u6_u3_n155 ) , .A1( u2_u6_u3_n97 ) );
  INV_X1 u2_u6_u3_U51 (.A( u2_u6_u3_n141 ) , .ZN( u2_u6_u3_n167 ) );
  AOI21_X1 u2_u6_u3_U52 (.B2( u2_u6_u3_n114 ) , .B1( u2_u6_u3_n146 ) , .A( u2_u6_u3_n154 ) , .ZN( u2_u6_u3_n94 ) );
  AOI21_X1 u2_u6_u3_U53 (.ZN( u2_u6_u3_n110 ) , .B2( u2_u6_u3_n142 ) , .B1( u2_u6_u3_n186 ) , .A( u2_u6_u3_n95 ) );
  INV_X1 u2_u6_u3_U54 (.A( u2_u6_u3_n145 ) , .ZN( u2_u6_u3_n186 ) );
  AOI21_X1 u2_u6_u3_U55 (.B1( u2_u6_u3_n124 ) , .A( u2_u6_u3_n149 ) , .B2( u2_u6_u3_n155 ) , .ZN( u2_u6_u3_n95 ) );
  INV_X1 u2_u6_u3_U56 (.A( u2_u6_u3_n149 ) , .ZN( u2_u6_u3_n169 ) );
  NAND2_X1 u2_u6_u3_U57 (.ZN( u2_u6_u3_n124 ) , .A1( u2_u6_u3_n96 ) , .A2( u2_u6_u3_n97 ) );
  NAND2_X1 u2_u6_u3_U58 (.A2( u2_u6_u3_n100 ) , .ZN( u2_u6_u3_n146 ) , .A1( u2_u6_u3_n96 ) );
  NAND2_X1 u2_u6_u3_U59 (.A1( u2_u6_u3_n101 ) , .ZN( u2_u6_u3_n145 ) , .A2( u2_u6_u3_n99 ) );
  AOI221_X1 u2_u6_u3_U6 (.A( u2_u6_u3_n131 ) , .C2( u2_u6_u3_n132 ) , .C1( u2_u6_u3_n133 ) , .ZN( u2_u6_u3_n134 ) , .B1( u2_u6_u3_n143 ) , .B2( u2_u6_u3_n177 ) );
  NAND2_X1 u2_u6_u3_U60 (.A1( u2_u6_u3_n100 ) , .ZN( u2_u6_u3_n156 ) , .A2( u2_u6_u3_n99 ) );
  NAND2_X1 u2_u6_u3_U61 (.A2( u2_u6_u3_n101 ) , .A1( u2_u6_u3_n104 ) , .ZN( u2_u6_u3_n148 ) );
  NAND2_X1 u2_u6_u3_U62 (.A1( u2_u6_u3_n100 ) , .A2( u2_u6_u3_n102 ) , .ZN( u2_u6_u3_n128 ) );
  NAND2_X1 u2_u6_u3_U63 (.A2( u2_u6_u3_n101 ) , .A1( u2_u6_u3_n102 ) , .ZN( u2_u6_u3_n152 ) );
  NAND2_X1 u2_u6_u3_U64 (.A2( u2_u6_u3_n101 ) , .ZN( u2_u6_u3_n114 ) , .A1( u2_u6_u3_n96 ) );
  NAND2_X1 u2_u6_u3_U65 (.ZN( u2_u6_u3_n107 ) , .A1( u2_u6_u3_n97 ) , .A2( u2_u6_u3_n99 ) );
  NAND2_X1 u2_u6_u3_U66 (.A2( u2_u6_u3_n100 ) , .A1( u2_u6_u3_n104 ) , .ZN( u2_u6_u3_n113 ) );
  NAND2_X1 u2_u6_u3_U67 (.A1( u2_u6_u3_n104 ) , .ZN( u2_u6_u3_n153 ) , .A2( u2_u6_u3_n97 ) );
  NAND2_X1 u2_u6_u3_U68 (.A2( u2_u6_u3_n103 ) , .A1( u2_u6_u3_n104 ) , .ZN( u2_u6_u3_n130 ) );
  NAND2_X1 u2_u6_u3_U69 (.A2( u2_u6_u3_n103 ) , .ZN( u2_u6_u3_n144 ) , .A1( u2_u6_u3_n96 ) );
  OAI22_X1 u2_u6_u3_U7 (.B2( u2_u6_u3_n147 ) , .A2( u2_u6_u3_n148 ) , .ZN( u2_u6_u3_n160 ) , .B1( u2_u6_u3_n165 ) , .A1( u2_u6_u3_n168 ) );
  NAND2_X1 u2_u6_u3_U70 (.A1( u2_u6_u3_n102 ) , .A2( u2_u6_u3_n103 ) , .ZN( u2_u6_u3_n108 ) );
  NOR2_X1 u2_u6_u3_U71 (.A2( u2_u6_X_19 ) , .A1( u2_u6_X_20 ) , .ZN( u2_u6_u3_n99 ) );
  NOR2_X1 u2_u6_u3_U72 (.A2( u2_u6_X_21 ) , .A1( u2_u6_X_24 ) , .ZN( u2_u6_u3_n103 ) );
  NOR2_X1 u2_u6_u3_U73 (.A2( u2_u6_X_24 ) , .A1( u2_u6_u3_n171 ) , .ZN( u2_u6_u3_n97 ) );
  NOR2_X1 u2_u6_u3_U74 (.A2( u2_u6_X_23 ) , .ZN( u2_u6_u3_n141 ) , .A1( u2_u6_u3_n166 ) );
  NOR2_X1 u2_u6_u3_U75 (.A2( u2_u6_X_19 ) , .A1( u2_u6_u3_n172 ) , .ZN( u2_u6_u3_n96 ) );
  NAND2_X1 u2_u6_u3_U76 (.A1( u2_u6_X_22 ) , .A2( u2_u6_X_23 ) , .ZN( u2_u6_u3_n154 ) );
  NAND2_X1 u2_u6_u3_U77 (.A1( u2_u6_X_23 ) , .ZN( u2_u6_u3_n149 ) , .A2( u2_u6_u3_n166 ) );
  NOR2_X1 u2_u6_u3_U78 (.A2( u2_u6_X_22 ) , .A1( u2_u6_X_23 ) , .ZN( u2_u6_u3_n121 ) );
  AND2_X1 u2_u6_u3_U79 (.A1( u2_u6_X_24 ) , .ZN( u2_u6_u3_n101 ) , .A2( u2_u6_u3_n171 ) );
  AND3_X1 u2_u6_u3_U8 (.A3( u2_u6_u3_n144 ) , .A2( u2_u6_u3_n145 ) , .A1( u2_u6_u3_n146 ) , .ZN( u2_u6_u3_n147 ) );
  AND2_X1 u2_u6_u3_U80 (.A1( u2_u6_X_19 ) , .ZN( u2_u6_u3_n102 ) , .A2( u2_u6_u3_n172 ) );
  AND2_X1 u2_u6_u3_U81 (.A1( u2_u6_X_21 ) , .A2( u2_u6_X_24 ) , .ZN( u2_u6_u3_n100 ) );
  AND2_X1 u2_u6_u3_U82 (.A2( u2_u6_X_19 ) , .A1( u2_u6_X_20 ) , .ZN( u2_u6_u3_n104 ) );
  INV_X1 u2_u6_u3_U83 (.A( u2_u6_X_22 ) , .ZN( u2_u6_u3_n166 ) );
  INV_X1 u2_u6_u3_U84 (.A( u2_u6_X_21 ) , .ZN( u2_u6_u3_n171 ) );
  INV_X1 u2_u6_u3_U85 (.A( u2_u6_X_20 ) , .ZN( u2_u6_u3_n172 ) );
  NAND4_X1 u2_u6_u3_U86 (.ZN( u2_out6_26 ) , .A4( u2_u6_u3_n109 ) , .A3( u2_u6_u3_n110 ) , .A2( u2_u6_u3_n111 ) , .A1( u2_u6_u3_n173 ) );
  INV_X1 u2_u6_u3_U87 (.ZN( u2_u6_u3_n173 ) , .A( u2_u6_u3_n94 ) );
  OAI21_X1 u2_u6_u3_U88 (.ZN( u2_u6_u3_n111 ) , .B2( u2_u6_u3_n117 ) , .A( u2_u6_u3_n133 ) , .B1( u2_u6_u3_n176 ) );
  NAND4_X1 u2_u6_u3_U89 (.ZN( u2_out6_20 ) , .A4( u2_u6_u3_n122 ) , .A3( u2_u6_u3_n123 ) , .A1( u2_u6_u3_n175 ) , .A2( u2_u6_u3_n180 ) );
  INV_X1 u2_u6_u3_U9 (.A( u2_u6_u3_n143 ) , .ZN( u2_u6_u3_n168 ) );
  INV_X1 u2_u6_u3_U90 (.A( u2_u6_u3_n126 ) , .ZN( u2_u6_u3_n180 ) );
  INV_X1 u2_u6_u3_U91 (.A( u2_u6_u3_n112 ) , .ZN( u2_u6_u3_n175 ) );
  NAND4_X1 u2_u6_u3_U92 (.ZN( u2_out6_1 ) , .A4( u2_u6_u3_n161 ) , .A3( u2_u6_u3_n162 ) , .A2( u2_u6_u3_n163 ) , .A1( u2_u6_u3_n185 ) );
  NAND2_X1 u2_u6_u3_U93 (.ZN( u2_u6_u3_n163 ) , .A2( u2_u6_u3_n170 ) , .A1( u2_u6_u3_n176 ) );
  AOI22_X1 u2_u6_u3_U94 (.B2( u2_u6_u3_n140 ) , .B1( u2_u6_u3_n141 ) , .A2( u2_u6_u3_n142 ) , .ZN( u2_u6_u3_n162 ) , .A1( u2_u6_u3_n177 ) );
  OR4_X1 u2_u6_u3_U95 (.ZN( u2_out6_10 ) , .A4( u2_u6_u3_n136 ) , .A3( u2_u6_u3_n137 ) , .A1( u2_u6_u3_n138 ) , .A2( u2_u6_u3_n139 ) );
  OAI222_X1 u2_u6_u3_U96 (.C1( u2_u6_u3_n128 ) , .ZN( u2_u6_u3_n137 ) , .B1( u2_u6_u3_n148 ) , .A2( u2_u6_u3_n150 ) , .B2( u2_u6_u3_n154 ) , .C2( u2_u6_u3_n164 ) , .A1( u2_u6_u3_n167 ) );
  OAI221_X1 u2_u6_u3_U97 (.A( u2_u6_u3_n134 ) , .B2( u2_u6_u3_n135 ) , .ZN( u2_u6_u3_n136 ) , .C1( u2_u6_u3_n149 ) , .B1( u2_u6_u3_n151 ) , .C2( u2_u6_u3_n183 ) );
  NAND3_X1 u2_u6_u3_U98 (.A1( u2_u6_u3_n114 ) , .ZN( u2_u6_u3_n115 ) , .A2( u2_u6_u3_n145 ) , .A3( u2_u6_u3_n153 ) );
  NAND3_X1 u2_u6_u3_U99 (.ZN( u2_u6_u3_n129 ) , .A2( u2_u6_u3_n144 ) , .A1( u2_u6_u3_n153 ) , .A3( u2_u6_u3_n182 ) );
  OAI22_X1 u2_u6_u4_U10 (.B2( u2_u6_u4_n135 ) , .ZN( u2_u6_u4_n137 ) , .B1( u2_u6_u4_n153 ) , .A1( u2_u6_u4_n155 ) , .A2( u2_u6_u4_n171 ) );
  AND3_X1 u2_u6_u4_U11 (.A2( u2_u6_u4_n134 ) , .ZN( u2_u6_u4_n135 ) , .A3( u2_u6_u4_n145 ) , .A1( u2_u6_u4_n157 ) );
  NAND2_X1 u2_u6_u4_U12 (.ZN( u2_u6_u4_n132 ) , .A2( u2_u6_u4_n170 ) , .A1( u2_u6_u4_n173 ) );
  AOI21_X1 u2_u6_u4_U13 (.B2( u2_u6_u4_n160 ) , .B1( u2_u6_u4_n161 ) , .ZN( u2_u6_u4_n162 ) , .A( u2_u6_u4_n170 ) );
  AOI21_X1 u2_u6_u4_U14 (.ZN( u2_u6_u4_n107 ) , .B2( u2_u6_u4_n143 ) , .A( u2_u6_u4_n174 ) , .B1( u2_u6_u4_n184 ) );
  AOI21_X1 u2_u6_u4_U15 (.B2( u2_u6_u4_n158 ) , .B1( u2_u6_u4_n159 ) , .ZN( u2_u6_u4_n163 ) , .A( u2_u6_u4_n174 ) );
  AOI21_X1 u2_u6_u4_U16 (.A( u2_u6_u4_n153 ) , .B2( u2_u6_u4_n154 ) , .B1( u2_u6_u4_n155 ) , .ZN( u2_u6_u4_n165 ) );
  AOI21_X1 u2_u6_u4_U17 (.A( u2_u6_u4_n156 ) , .B2( u2_u6_u4_n157 ) , .ZN( u2_u6_u4_n164 ) , .B1( u2_u6_u4_n184 ) );
  INV_X1 u2_u6_u4_U18 (.A( u2_u6_u4_n138 ) , .ZN( u2_u6_u4_n170 ) );
  AND2_X1 u2_u6_u4_U19 (.A2( u2_u6_u4_n120 ) , .ZN( u2_u6_u4_n155 ) , .A1( u2_u6_u4_n160 ) );
  INV_X1 u2_u6_u4_U20 (.A( u2_u6_u4_n156 ) , .ZN( u2_u6_u4_n175 ) );
  NAND2_X1 u2_u6_u4_U21 (.A2( u2_u6_u4_n118 ) , .ZN( u2_u6_u4_n131 ) , .A1( u2_u6_u4_n147 ) );
  NAND2_X1 u2_u6_u4_U22 (.A1( u2_u6_u4_n119 ) , .A2( u2_u6_u4_n120 ) , .ZN( u2_u6_u4_n130 ) );
  NAND2_X1 u2_u6_u4_U23 (.ZN( u2_u6_u4_n117 ) , .A2( u2_u6_u4_n118 ) , .A1( u2_u6_u4_n148 ) );
  NAND2_X1 u2_u6_u4_U24 (.ZN( u2_u6_u4_n129 ) , .A1( u2_u6_u4_n134 ) , .A2( u2_u6_u4_n148 ) );
  AND3_X1 u2_u6_u4_U25 (.A1( u2_u6_u4_n119 ) , .A2( u2_u6_u4_n143 ) , .A3( u2_u6_u4_n154 ) , .ZN( u2_u6_u4_n161 ) );
  AND2_X1 u2_u6_u4_U26 (.A1( u2_u6_u4_n145 ) , .A2( u2_u6_u4_n147 ) , .ZN( u2_u6_u4_n159 ) );
  OR3_X1 u2_u6_u4_U27 (.A3( u2_u6_u4_n114 ) , .A2( u2_u6_u4_n115 ) , .A1( u2_u6_u4_n116 ) , .ZN( u2_u6_u4_n136 ) );
  AOI21_X1 u2_u6_u4_U28 (.A( u2_u6_u4_n113 ) , .ZN( u2_u6_u4_n116 ) , .B2( u2_u6_u4_n173 ) , .B1( u2_u6_u4_n174 ) );
  AOI21_X1 u2_u6_u4_U29 (.ZN( u2_u6_u4_n115 ) , .B2( u2_u6_u4_n145 ) , .B1( u2_u6_u4_n146 ) , .A( u2_u6_u4_n156 ) );
  NOR2_X1 u2_u6_u4_U3 (.ZN( u2_u6_u4_n121 ) , .A1( u2_u6_u4_n181 ) , .A2( u2_u6_u4_n182 ) );
  OAI22_X1 u2_u6_u4_U30 (.ZN( u2_u6_u4_n114 ) , .A2( u2_u6_u4_n121 ) , .B1( u2_u6_u4_n160 ) , .B2( u2_u6_u4_n170 ) , .A1( u2_u6_u4_n171 ) );
  INV_X1 u2_u6_u4_U31 (.A( u2_u6_u4_n158 ) , .ZN( u2_u6_u4_n182 ) );
  INV_X1 u2_u6_u4_U32 (.ZN( u2_u6_u4_n181 ) , .A( u2_u6_u4_n96 ) );
  INV_X1 u2_u6_u4_U33 (.A( u2_u6_u4_n144 ) , .ZN( u2_u6_u4_n179 ) );
  INV_X1 u2_u6_u4_U34 (.A( u2_u6_u4_n157 ) , .ZN( u2_u6_u4_n178 ) );
  NAND2_X1 u2_u6_u4_U35 (.A2( u2_u6_u4_n154 ) , .A1( u2_u6_u4_n96 ) , .ZN( u2_u6_u4_n97 ) );
  INV_X1 u2_u6_u4_U36 (.ZN( u2_u6_u4_n186 ) , .A( u2_u6_u4_n95 ) );
  OAI221_X1 u2_u6_u4_U37 (.C1( u2_u6_u4_n134 ) , .B1( u2_u6_u4_n158 ) , .B2( u2_u6_u4_n171 ) , .C2( u2_u6_u4_n173 ) , .A( u2_u6_u4_n94 ) , .ZN( u2_u6_u4_n95 ) );
  AOI222_X1 u2_u6_u4_U38 (.B2( u2_u6_u4_n132 ) , .A1( u2_u6_u4_n138 ) , .C2( u2_u6_u4_n175 ) , .A2( u2_u6_u4_n179 ) , .C1( u2_u6_u4_n181 ) , .B1( u2_u6_u4_n185 ) , .ZN( u2_u6_u4_n94 ) );
  INV_X1 u2_u6_u4_U39 (.A( u2_u6_u4_n113 ) , .ZN( u2_u6_u4_n185 ) );
  INV_X1 u2_u6_u4_U4 (.A( u2_u6_u4_n117 ) , .ZN( u2_u6_u4_n184 ) );
  INV_X1 u2_u6_u4_U40 (.A( u2_u6_u4_n143 ) , .ZN( u2_u6_u4_n183 ) );
  NOR2_X1 u2_u6_u4_U41 (.ZN( u2_u6_u4_n138 ) , .A1( u2_u6_u4_n168 ) , .A2( u2_u6_u4_n169 ) );
  NOR2_X1 u2_u6_u4_U42 (.A1( u2_u6_u4_n150 ) , .A2( u2_u6_u4_n152 ) , .ZN( u2_u6_u4_n153 ) );
  NOR2_X1 u2_u6_u4_U43 (.A2( u2_u6_u4_n128 ) , .A1( u2_u6_u4_n138 ) , .ZN( u2_u6_u4_n156 ) );
  AOI22_X1 u2_u6_u4_U44 (.B2( u2_u6_u4_n122 ) , .A1( u2_u6_u4_n123 ) , .ZN( u2_u6_u4_n124 ) , .B1( u2_u6_u4_n128 ) , .A2( u2_u6_u4_n172 ) );
  INV_X1 u2_u6_u4_U45 (.A( u2_u6_u4_n153 ) , .ZN( u2_u6_u4_n172 ) );
  NAND2_X1 u2_u6_u4_U46 (.A2( u2_u6_u4_n120 ) , .ZN( u2_u6_u4_n123 ) , .A1( u2_u6_u4_n161 ) );
  AOI22_X1 u2_u6_u4_U47 (.B2( u2_u6_u4_n132 ) , .A2( u2_u6_u4_n133 ) , .ZN( u2_u6_u4_n140 ) , .A1( u2_u6_u4_n150 ) , .B1( u2_u6_u4_n179 ) );
  NAND2_X1 u2_u6_u4_U48 (.ZN( u2_u6_u4_n133 ) , .A2( u2_u6_u4_n146 ) , .A1( u2_u6_u4_n154 ) );
  NAND2_X1 u2_u6_u4_U49 (.A1( u2_u6_u4_n103 ) , .ZN( u2_u6_u4_n154 ) , .A2( u2_u6_u4_n98 ) );
  NOR4_X1 u2_u6_u4_U5 (.A4( u2_u6_u4_n106 ) , .A3( u2_u6_u4_n107 ) , .A2( u2_u6_u4_n108 ) , .A1( u2_u6_u4_n109 ) , .ZN( u2_u6_u4_n110 ) );
  NAND2_X1 u2_u6_u4_U50 (.A1( u2_u6_u4_n101 ) , .ZN( u2_u6_u4_n158 ) , .A2( u2_u6_u4_n99 ) );
  AOI21_X1 u2_u6_u4_U51 (.ZN( u2_u6_u4_n127 ) , .A( u2_u6_u4_n136 ) , .B2( u2_u6_u4_n150 ) , .B1( u2_u6_u4_n180 ) );
  INV_X1 u2_u6_u4_U52 (.A( u2_u6_u4_n160 ) , .ZN( u2_u6_u4_n180 ) );
  NAND2_X1 u2_u6_u4_U53 (.A2( u2_u6_u4_n104 ) , .A1( u2_u6_u4_n105 ) , .ZN( u2_u6_u4_n146 ) );
  NAND2_X1 u2_u6_u4_U54 (.A2( u2_u6_u4_n101 ) , .A1( u2_u6_u4_n102 ) , .ZN( u2_u6_u4_n160 ) );
  NAND2_X1 u2_u6_u4_U55 (.ZN( u2_u6_u4_n134 ) , .A1( u2_u6_u4_n98 ) , .A2( u2_u6_u4_n99 ) );
  NAND2_X1 u2_u6_u4_U56 (.A1( u2_u6_u4_n103 ) , .A2( u2_u6_u4_n104 ) , .ZN( u2_u6_u4_n143 ) );
  NAND2_X1 u2_u6_u4_U57 (.A2( u2_u6_u4_n105 ) , .ZN( u2_u6_u4_n145 ) , .A1( u2_u6_u4_n98 ) );
  NAND2_X1 u2_u6_u4_U58 (.A1( u2_u6_u4_n100 ) , .A2( u2_u6_u4_n105 ) , .ZN( u2_u6_u4_n120 ) );
  NAND2_X1 u2_u6_u4_U59 (.A1( u2_u6_u4_n102 ) , .A2( u2_u6_u4_n104 ) , .ZN( u2_u6_u4_n148 ) );
  AOI21_X1 u2_u6_u4_U6 (.ZN( u2_u6_u4_n106 ) , .B2( u2_u6_u4_n146 ) , .B1( u2_u6_u4_n158 ) , .A( u2_u6_u4_n170 ) );
  NAND2_X1 u2_u6_u4_U60 (.A2( u2_u6_u4_n100 ) , .A1( u2_u6_u4_n103 ) , .ZN( u2_u6_u4_n157 ) );
  INV_X1 u2_u6_u4_U61 (.A( u2_u6_u4_n150 ) , .ZN( u2_u6_u4_n173 ) );
  INV_X1 u2_u6_u4_U62 (.A( u2_u6_u4_n152 ) , .ZN( u2_u6_u4_n171 ) );
  NAND2_X1 u2_u6_u4_U63 (.A1( u2_u6_u4_n100 ) , .ZN( u2_u6_u4_n118 ) , .A2( u2_u6_u4_n99 ) );
  NAND2_X1 u2_u6_u4_U64 (.A2( u2_u6_u4_n100 ) , .A1( u2_u6_u4_n102 ) , .ZN( u2_u6_u4_n144 ) );
  NAND2_X1 u2_u6_u4_U65 (.A2( u2_u6_u4_n101 ) , .A1( u2_u6_u4_n105 ) , .ZN( u2_u6_u4_n96 ) );
  INV_X1 u2_u6_u4_U66 (.A( u2_u6_u4_n128 ) , .ZN( u2_u6_u4_n174 ) );
  NAND2_X1 u2_u6_u4_U67 (.A2( u2_u6_u4_n102 ) , .ZN( u2_u6_u4_n119 ) , .A1( u2_u6_u4_n98 ) );
  NAND2_X1 u2_u6_u4_U68 (.A2( u2_u6_u4_n101 ) , .A1( u2_u6_u4_n103 ) , .ZN( u2_u6_u4_n147 ) );
  NAND2_X1 u2_u6_u4_U69 (.A2( u2_u6_u4_n104 ) , .ZN( u2_u6_u4_n113 ) , .A1( u2_u6_u4_n99 ) );
  AOI21_X1 u2_u6_u4_U7 (.ZN( u2_u6_u4_n108 ) , .B2( u2_u6_u4_n134 ) , .B1( u2_u6_u4_n155 ) , .A( u2_u6_u4_n156 ) );
  NOR2_X1 u2_u6_u4_U70 (.A2( u2_u6_X_28 ) , .ZN( u2_u6_u4_n150 ) , .A1( u2_u6_u4_n168 ) );
  NOR2_X1 u2_u6_u4_U71 (.A2( u2_u6_X_29 ) , .ZN( u2_u6_u4_n152 ) , .A1( u2_u6_u4_n169 ) );
  NOR2_X1 u2_u6_u4_U72 (.A2( u2_u6_X_30 ) , .ZN( u2_u6_u4_n105 ) , .A1( u2_u6_u4_n176 ) );
  NOR2_X1 u2_u6_u4_U73 (.A2( u2_u6_X_26 ) , .ZN( u2_u6_u4_n100 ) , .A1( u2_u6_u4_n177 ) );
  NOR2_X1 u2_u6_u4_U74 (.A2( u2_u6_X_28 ) , .A1( u2_u6_X_29 ) , .ZN( u2_u6_u4_n128 ) );
  NOR2_X1 u2_u6_u4_U75 (.A2( u2_u6_X_27 ) , .A1( u2_u6_X_30 ) , .ZN( u2_u6_u4_n102 ) );
  NOR2_X1 u2_u6_u4_U76 (.A2( u2_u6_X_25 ) , .A1( u2_u6_X_26 ) , .ZN( u2_u6_u4_n98 ) );
  AND2_X1 u2_u6_u4_U77 (.A2( u2_u6_X_25 ) , .A1( u2_u6_X_26 ) , .ZN( u2_u6_u4_n104 ) );
  AND2_X1 u2_u6_u4_U78 (.A1( u2_u6_X_30 ) , .A2( u2_u6_u4_n176 ) , .ZN( u2_u6_u4_n99 ) );
  AND2_X1 u2_u6_u4_U79 (.A1( u2_u6_X_26 ) , .ZN( u2_u6_u4_n101 ) , .A2( u2_u6_u4_n177 ) );
  AOI21_X1 u2_u6_u4_U8 (.ZN( u2_u6_u4_n109 ) , .A( u2_u6_u4_n153 ) , .B1( u2_u6_u4_n159 ) , .B2( u2_u6_u4_n184 ) );
  AND2_X1 u2_u6_u4_U80 (.A1( u2_u6_X_27 ) , .A2( u2_u6_X_30 ) , .ZN( u2_u6_u4_n103 ) );
  INV_X1 u2_u6_u4_U81 (.A( u2_u6_X_28 ) , .ZN( u2_u6_u4_n169 ) );
  INV_X1 u2_u6_u4_U82 (.A( u2_u6_X_29 ) , .ZN( u2_u6_u4_n168 ) );
  INV_X1 u2_u6_u4_U83 (.A( u2_u6_X_25 ) , .ZN( u2_u6_u4_n177 ) );
  INV_X1 u2_u6_u4_U84 (.A( u2_u6_X_27 ) , .ZN( u2_u6_u4_n176 ) );
  NAND4_X1 u2_u6_u4_U85 (.ZN( u2_out6_25 ) , .A4( u2_u6_u4_n139 ) , .A3( u2_u6_u4_n140 ) , .A2( u2_u6_u4_n141 ) , .A1( u2_u6_u4_n142 ) );
  OAI21_X1 u2_u6_u4_U86 (.B2( u2_u6_u4_n131 ) , .ZN( u2_u6_u4_n141 ) , .A( u2_u6_u4_n175 ) , .B1( u2_u6_u4_n183 ) );
  OAI21_X1 u2_u6_u4_U87 (.A( u2_u6_u4_n128 ) , .B2( u2_u6_u4_n129 ) , .B1( u2_u6_u4_n130 ) , .ZN( u2_u6_u4_n142 ) );
  NAND4_X1 u2_u6_u4_U88 (.ZN( u2_out6_14 ) , .A4( u2_u6_u4_n124 ) , .A3( u2_u6_u4_n125 ) , .A2( u2_u6_u4_n126 ) , .A1( u2_u6_u4_n127 ) );
  AOI22_X1 u2_u6_u4_U89 (.B2( u2_u6_u4_n117 ) , .ZN( u2_u6_u4_n126 ) , .A1( u2_u6_u4_n129 ) , .B1( u2_u6_u4_n152 ) , .A2( u2_u6_u4_n175 ) );
  AOI211_X1 u2_u6_u4_U9 (.B( u2_u6_u4_n136 ) , .A( u2_u6_u4_n137 ) , .C2( u2_u6_u4_n138 ) , .ZN( u2_u6_u4_n139 ) , .C1( u2_u6_u4_n182 ) );
  AOI22_X1 u2_u6_u4_U90 (.ZN( u2_u6_u4_n125 ) , .B2( u2_u6_u4_n131 ) , .A2( u2_u6_u4_n132 ) , .B1( u2_u6_u4_n138 ) , .A1( u2_u6_u4_n178 ) );
  NAND4_X1 u2_u6_u4_U91 (.ZN( u2_out6_8 ) , .A4( u2_u6_u4_n110 ) , .A3( u2_u6_u4_n111 ) , .A2( u2_u6_u4_n112 ) , .A1( u2_u6_u4_n186 ) );
  NAND2_X1 u2_u6_u4_U92 (.ZN( u2_u6_u4_n112 ) , .A2( u2_u6_u4_n130 ) , .A1( u2_u6_u4_n150 ) );
  AOI22_X1 u2_u6_u4_U93 (.ZN( u2_u6_u4_n111 ) , .B2( u2_u6_u4_n132 ) , .A1( u2_u6_u4_n152 ) , .B1( u2_u6_u4_n178 ) , .A2( u2_u6_u4_n97 ) );
  AOI22_X1 u2_u6_u4_U94 (.B2( u2_u6_u4_n149 ) , .B1( u2_u6_u4_n150 ) , .A2( u2_u6_u4_n151 ) , .A1( u2_u6_u4_n152 ) , .ZN( u2_u6_u4_n167 ) );
  NOR4_X1 u2_u6_u4_U95 (.A4( u2_u6_u4_n162 ) , .A3( u2_u6_u4_n163 ) , .A2( u2_u6_u4_n164 ) , .A1( u2_u6_u4_n165 ) , .ZN( u2_u6_u4_n166 ) );
  NAND3_X1 u2_u6_u4_U96 (.ZN( u2_out6_3 ) , .A3( u2_u6_u4_n166 ) , .A1( u2_u6_u4_n167 ) , .A2( u2_u6_u4_n186 ) );
  NAND3_X1 u2_u6_u4_U97 (.A3( u2_u6_u4_n146 ) , .A2( u2_u6_u4_n147 ) , .A1( u2_u6_u4_n148 ) , .ZN( u2_u6_u4_n149 ) );
  NAND3_X1 u2_u6_u4_U98 (.A3( u2_u6_u4_n143 ) , .A2( u2_u6_u4_n144 ) , .A1( u2_u6_u4_n145 ) , .ZN( u2_u6_u4_n151 ) );
  NAND3_X1 u2_u6_u4_U99 (.A3( u2_u6_u4_n121 ) , .ZN( u2_u6_u4_n122 ) , .A2( u2_u6_u4_n144 ) , .A1( u2_u6_u4_n154 ) );
  INV_X1 u2_u6_u5_U10 (.A( u2_u6_u5_n121 ) , .ZN( u2_u6_u5_n177 ) );
  NOR3_X1 u2_u6_u5_U100 (.A3( u2_u6_u5_n141 ) , .A1( u2_u6_u5_n142 ) , .ZN( u2_u6_u5_n143 ) , .A2( u2_u6_u5_n191 ) );
  NAND4_X1 u2_u6_u5_U101 (.ZN( u2_out6_4 ) , .A4( u2_u6_u5_n112 ) , .A2( u2_u6_u5_n113 ) , .A1( u2_u6_u5_n114 ) , .A3( u2_u6_u5_n195 ) );
  AOI211_X1 u2_u6_u5_U102 (.A( u2_u6_u5_n110 ) , .C1( u2_u6_u5_n111 ) , .ZN( u2_u6_u5_n112 ) , .B( u2_u6_u5_n118 ) , .C2( u2_u6_u5_n177 ) );
  AOI222_X1 u2_u6_u5_U103 (.ZN( u2_u6_u5_n113 ) , .A1( u2_u6_u5_n131 ) , .C1( u2_u6_u5_n148 ) , .B2( u2_u6_u5_n174 ) , .C2( u2_u6_u5_n178 ) , .A2( u2_u6_u5_n179 ) , .B1( u2_u6_u5_n99 ) );
  NAND3_X1 u2_u6_u5_U104 (.A2( u2_u6_u5_n154 ) , .A3( u2_u6_u5_n158 ) , .A1( u2_u6_u5_n161 ) , .ZN( u2_u6_u5_n99 ) );
  NOR2_X1 u2_u6_u5_U11 (.ZN( u2_u6_u5_n160 ) , .A2( u2_u6_u5_n173 ) , .A1( u2_u6_u5_n177 ) );
  INV_X1 u2_u6_u5_U12 (.A( u2_u6_u5_n150 ) , .ZN( u2_u6_u5_n174 ) );
  AOI21_X1 u2_u6_u5_U13 (.A( u2_u6_u5_n160 ) , .B2( u2_u6_u5_n161 ) , .ZN( u2_u6_u5_n162 ) , .B1( u2_u6_u5_n192 ) );
  INV_X1 u2_u6_u5_U14 (.A( u2_u6_u5_n159 ) , .ZN( u2_u6_u5_n192 ) );
  AOI21_X1 u2_u6_u5_U15 (.A( u2_u6_u5_n156 ) , .B2( u2_u6_u5_n157 ) , .B1( u2_u6_u5_n158 ) , .ZN( u2_u6_u5_n163 ) );
  AOI21_X1 u2_u6_u5_U16 (.B2( u2_u6_u5_n139 ) , .B1( u2_u6_u5_n140 ) , .ZN( u2_u6_u5_n141 ) , .A( u2_u6_u5_n150 ) );
  OAI21_X1 u2_u6_u5_U17 (.A( u2_u6_u5_n133 ) , .B2( u2_u6_u5_n134 ) , .B1( u2_u6_u5_n135 ) , .ZN( u2_u6_u5_n142 ) );
  OAI21_X1 u2_u6_u5_U18 (.ZN( u2_u6_u5_n133 ) , .B2( u2_u6_u5_n147 ) , .A( u2_u6_u5_n173 ) , .B1( u2_u6_u5_n188 ) );
  NAND2_X1 u2_u6_u5_U19 (.A2( u2_u6_u5_n119 ) , .A1( u2_u6_u5_n123 ) , .ZN( u2_u6_u5_n137 ) );
  INV_X1 u2_u6_u5_U20 (.A( u2_u6_u5_n155 ) , .ZN( u2_u6_u5_n194 ) );
  NAND2_X1 u2_u6_u5_U21 (.A1( u2_u6_u5_n121 ) , .ZN( u2_u6_u5_n132 ) , .A2( u2_u6_u5_n172 ) );
  NAND2_X1 u2_u6_u5_U22 (.A2( u2_u6_u5_n122 ) , .ZN( u2_u6_u5_n136 ) , .A1( u2_u6_u5_n154 ) );
  NAND2_X1 u2_u6_u5_U23 (.A2( u2_u6_u5_n119 ) , .A1( u2_u6_u5_n120 ) , .ZN( u2_u6_u5_n159 ) );
  INV_X1 u2_u6_u5_U24 (.A( u2_u6_u5_n156 ) , .ZN( u2_u6_u5_n175 ) );
  INV_X1 u2_u6_u5_U25 (.A( u2_u6_u5_n158 ) , .ZN( u2_u6_u5_n188 ) );
  INV_X1 u2_u6_u5_U26 (.A( u2_u6_u5_n152 ) , .ZN( u2_u6_u5_n179 ) );
  INV_X1 u2_u6_u5_U27 (.A( u2_u6_u5_n140 ) , .ZN( u2_u6_u5_n182 ) );
  INV_X1 u2_u6_u5_U28 (.A( u2_u6_u5_n151 ) , .ZN( u2_u6_u5_n183 ) );
  INV_X1 u2_u6_u5_U29 (.A( u2_u6_u5_n123 ) , .ZN( u2_u6_u5_n185 ) );
  NOR2_X1 u2_u6_u5_U3 (.ZN( u2_u6_u5_n134 ) , .A1( u2_u6_u5_n183 ) , .A2( u2_u6_u5_n190 ) );
  INV_X1 u2_u6_u5_U30 (.A( u2_u6_u5_n161 ) , .ZN( u2_u6_u5_n184 ) );
  INV_X1 u2_u6_u5_U31 (.A( u2_u6_u5_n139 ) , .ZN( u2_u6_u5_n189 ) );
  INV_X1 u2_u6_u5_U32 (.A( u2_u6_u5_n157 ) , .ZN( u2_u6_u5_n190 ) );
  INV_X1 u2_u6_u5_U33 (.A( u2_u6_u5_n120 ) , .ZN( u2_u6_u5_n193 ) );
  NAND2_X1 u2_u6_u5_U34 (.ZN( u2_u6_u5_n111 ) , .A1( u2_u6_u5_n140 ) , .A2( u2_u6_u5_n155 ) );
  INV_X1 u2_u6_u5_U35 (.A( u2_u6_u5_n117 ) , .ZN( u2_u6_u5_n196 ) );
  OAI221_X1 u2_u6_u5_U36 (.A( u2_u6_u5_n116 ) , .ZN( u2_u6_u5_n117 ) , .B2( u2_u6_u5_n119 ) , .C1( u2_u6_u5_n153 ) , .C2( u2_u6_u5_n158 ) , .B1( u2_u6_u5_n172 ) );
  AOI222_X1 u2_u6_u5_U37 (.ZN( u2_u6_u5_n116 ) , .B2( u2_u6_u5_n145 ) , .C1( u2_u6_u5_n148 ) , .A2( u2_u6_u5_n174 ) , .C2( u2_u6_u5_n177 ) , .B1( u2_u6_u5_n187 ) , .A1( u2_u6_u5_n193 ) );
  INV_X1 u2_u6_u5_U38 (.A( u2_u6_u5_n115 ) , .ZN( u2_u6_u5_n187 ) );
  NOR2_X1 u2_u6_u5_U39 (.ZN( u2_u6_u5_n100 ) , .A1( u2_u6_u5_n170 ) , .A2( u2_u6_u5_n180 ) );
  INV_X1 u2_u6_u5_U4 (.A( u2_u6_u5_n138 ) , .ZN( u2_u6_u5_n191 ) );
  AOI22_X1 u2_u6_u5_U40 (.B2( u2_u6_u5_n131 ) , .A2( u2_u6_u5_n146 ) , .ZN( u2_u6_u5_n169 ) , .B1( u2_u6_u5_n174 ) , .A1( u2_u6_u5_n185 ) );
  NOR2_X1 u2_u6_u5_U41 (.A1( u2_u6_u5_n146 ) , .ZN( u2_u6_u5_n150 ) , .A2( u2_u6_u5_n173 ) );
  AOI21_X1 u2_u6_u5_U42 (.A( u2_u6_u5_n118 ) , .B2( u2_u6_u5_n145 ) , .ZN( u2_u6_u5_n168 ) , .B1( u2_u6_u5_n186 ) );
  INV_X1 u2_u6_u5_U43 (.A( u2_u6_u5_n122 ) , .ZN( u2_u6_u5_n186 ) );
  NOR2_X1 u2_u6_u5_U44 (.A1( u2_u6_u5_n146 ) , .ZN( u2_u6_u5_n152 ) , .A2( u2_u6_u5_n176 ) );
  NOR2_X1 u2_u6_u5_U45 (.A1( u2_u6_u5_n115 ) , .ZN( u2_u6_u5_n118 ) , .A2( u2_u6_u5_n153 ) );
  NOR2_X1 u2_u6_u5_U46 (.A2( u2_u6_u5_n145 ) , .ZN( u2_u6_u5_n156 ) , .A1( u2_u6_u5_n174 ) );
  NOR2_X1 u2_u6_u5_U47 (.ZN( u2_u6_u5_n121 ) , .A2( u2_u6_u5_n145 ) , .A1( u2_u6_u5_n176 ) );
  AOI22_X1 u2_u6_u5_U48 (.ZN( u2_u6_u5_n114 ) , .A2( u2_u6_u5_n137 ) , .A1( u2_u6_u5_n145 ) , .B2( u2_u6_u5_n175 ) , .B1( u2_u6_u5_n193 ) );
  OAI211_X1 u2_u6_u5_U49 (.B( u2_u6_u5_n124 ) , .A( u2_u6_u5_n125 ) , .C2( u2_u6_u5_n126 ) , .C1( u2_u6_u5_n127 ) , .ZN( u2_u6_u5_n128 ) );
  OAI21_X1 u2_u6_u5_U5 (.B2( u2_u6_u5_n136 ) , .B1( u2_u6_u5_n137 ) , .ZN( u2_u6_u5_n138 ) , .A( u2_u6_u5_n177 ) );
  NOR3_X1 u2_u6_u5_U50 (.ZN( u2_u6_u5_n127 ) , .A1( u2_u6_u5_n136 ) , .A3( u2_u6_u5_n148 ) , .A2( u2_u6_u5_n182 ) );
  OAI21_X1 u2_u6_u5_U51 (.ZN( u2_u6_u5_n124 ) , .A( u2_u6_u5_n177 ) , .B2( u2_u6_u5_n183 ) , .B1( u2_u6_u5_n189 ) );
  OAI21_X1 u2_u6_u5_U52 (.ZN( u2_u6_u5_n125 ) , .A( u2_u6_u5_n174 ) , .B2( u2_u6_u5_n185 ) , .B1( u2_u6_u5_n190 ) );
  AOI21_X1 u2_u6_u5_U53 (.A( u2_u6_u5_n153 ) , .B2( u2_u6_u5_n154 ) , .B1( u2_u6_u5_n155 ) , .ZN( u2_u6_u5_n164 ) );
  AOI21_X1 u2_u6_u5_U54 (.ZN( u2_u6_u5_n110 ) , .B1( u2_u6_u5_n122 ) , .B2( u2_u6_u5_n139 ) , .A( u2_u6_u5_n153 ) );
  INV_X1 u2_u6_u5_U55 (.A( u2_u6_u5_n153 ) , .ZN( u2_u6_u5_n176 ) );
  INV_X1 u2_u6_u5_U56 (.A( u2_u6_u5_n126 ) , .ZN( u2_u6_u5_n173 ) );
  AND2_X1 u2_u6_u5_U57 (.A2( u2_u6_u5_n104 ) , .A1( u2_u6_u5_n107 ) , .ZN( u2_u6_u5_n147 ) );
  AND2_X1 u2_u6_u5_U58 (.A2( u2_u6_u5_n104 ) , .A1( u2_u6_u5_n108 ) , .ZN( u2_u6_u5_n148 ) );
  NAND2_X1 u2_u6_u5_U59 (.A1( u2_u6_u5_n105 ) , .A2( u2_u6_u5_n106 ) , .ZN( u2_u6_u5_n158 ) );
  INV_X1 u2_u6_u5_U6 (.A( u2_u6_u5_n135 ) , .ZN( u2_u6_u5_n178 ) );
  NAND2_X1 u2_u6_u5_U60 (.A2( u2_u6_u5_n108 ) , .A1( u2_u6_u5_n109 ) , .ZN( u2_u6_u5_n139 ) );
  NAND2_X1 u2_u6_u5_U61 (.A1( u2_u6_u5_n106 ) , .A2( u2_u6_u5_n108 ) , .ZN( u2_u6_u5_n119 ) );
  NAND2_X1 u2_u6_u5_U62 (.A2( u2_u6_u5_n103 ) , .A1( u2_u6_u5_n105 ) , .ZN( u2_u6_u5_n140 ) );
  NAND2_X1 u2_u6_u5_U63 (.A2( u2_u6_u5_n104 ) , .A1( u2_u6_u5_n105 ) , .ZN( u2_u6_u5_n155 ) );
  NAND2_X1 u2_u6_u5_U64 (.A2( u2_u6_u5_n106 ) , .A1( u2_u6_u5_n107 ) , .ZN( u2_u6_u5_n122 ) );
  NAND2_X1 u2_u6_u5_U65 (.A2( u2_u6_u5_n100 ) , .A1( u2_u6_u5_n106 ) , .ZN( u2_u6_u5_n115 ) );
  NAND2_X1 u2_u6_u5_U66 (.A2( u2_u6_u5_n100 ) , .A1( u2_u6_u5_n103 ) , .ZN( u2_u6_u5_n161 ) );
  NAND2_X1 u2_u6_u5_U67 (.A1( u2_u6_u5_n105 ) , .A2( u2_u6_u5_n109 ) , .ZN( u2_u6_u5_n154 ) );
  INV_X1 u2_u6_u5_U68 (.A( u2_u6_u5_n146 ) , .ZN( u2_u6_u5_n172 ) );
  NAND2_X1 u2_u6_u5_U69 (.A1( u2_u6_u5_n103 ) , .A2( u2_u6_u5_n108 ) , .ZN( u2_u6_u5_n123 ) );
  OAI22_X1 u2_u6_u5_U7 (.B2( u2_u6_u5_n149 ) , .B1( u2_u6_u5_n150 ) , .A2( u2_u6_u5_n151 ) , .A1( u2_u6_u5_n152 ) , .ZN( u2_u6_u5_n165 ) );
  NAND2_X1 u2_u6_u5_U70 (.A2( u2_u6_u5_n103 ) , .A1( u2_u6_u5_n107 ) , .ZN( u2_u6_u5_n151 ) );
  NAND2_X1 u2_u6_u5_U71 (.A2( u2_u6_u5_n107 ) , .A1( u2_u6_u5_n109 ) , .ZN( u2_u6_u5_n120 ) );
  NAND2_X1 u2_u6_u5_U72 (.A2( u2_u6_u5_n100 ) , .A1( u2_u6_u5_n109 ) , .ZN( u2_u6_u5_n157 ) );
  AND2_X1 u2_u6_u5_U73 (.A2( u2_u6_u5_n100 ) , .A1( u2_u6_u5_n104 ) , .ZN( u2_u6_u5_n131 ) );
  INV_X1 u2_u6_u5_U74 (.A( u2_u6_u5_n102 ) , .ZN( u2_u6_u5_n195 ) );
  OAI221_X1 u2_u6_u5_U75 (.A( u2_u6_u5_n101 ) , .ZN( u2_u6_u5_n102 ) , .C2( u2_u6_u5_n115 ) , .C1( u2_u6_u5_n126 ) , .B1( u2_u6_u5_n134 ) , .B2( u2_u6_u5_n160 ) );
  OAI21_X1 u2_u6_u5_U76 (.ZN( u2_u6_u5_n101 ) , .B1( u2_u6_u5_n137 ) , .A( u2_u6_u5_n146 ) , .B2( u2_u6_u5_n147 ) );
  NOR2_X1 u2_u6_u5_U77 (.A2( u2_u6_X_34 ) , .A1( u2_u6_X_35 ) , .ZN( u2_u6_u5_n145 ) );
  NOR2_X1 u2_u6_u5_U78 (.A2( u2_u6_X_34 ) , .ZN( u2_u6_u5_n146 ) , .A1( u2_u6_u5_n171 ) );
  NOR2_X1 u2_u6_u5_U79 (.A2( u2_u6_X_31 ) , .A1( u2_u6_X_32 ) , .ZN( u2_u6_u5_n103 ) );
  NOR3_X1 u2_u6_u5_U8 (.A2( u2_u6_u5_n147 ) , .A1( u2_u6_u5_n148 ) , .ZN( u2_u6_u5_n149 ) , .A3( u2_u6_u5_n194 ) );
  NOR2_X1 u2_u6_u5_U80 (.A2( u2_u6_X_36 ) , .ZN( u2_u6_u5_n105 ) , .A1( u2_u6_u5_n180 ) );
  NOR2_X1 u2_u6_u5_U81 (.A2( u2_u6_X_33 ) , .ZN( u2_u6_u5_n108 ) , .A1( u2_u6_u5_n170 ) );
  NOR2_X1 u2_u6_u5_U82 (.A2( u2_u6_X_33 ) , .A1( u2_u6_X_36 ) , .ZN( u2_u6_u5_n107 ) );
  NOR2_X1 u2_u6_u5_U83 (.A2( u2_u6_X_31 ) , .ZN( u2_u6_u5_n104 ) , .A1( u2_u6_u5_n181 ) );
  NAND2_X1 u2_u6_u5_U84 (.A2( u2_u6_X_34 ) , .A1( u2_u6_X_35 ) , .ZN( u2_u6_u5_n153 ) );
  NAND2_X1 u2_u6_u5_U85 (.A1( u2_u6_X_34 ) , .ZN( u2_u6_u5_n126 ) , .A2( u2_u6_u5_n171 ) );
  AND2_X1 u2_u6_u5_U86 (.A1( u2_u6_X_31 ) , .A2( u2_u6_X_32 ) , .ZN( u2_u6_u5_n106 ) );
  AND2_X1 u2_u6_u5_U87 (.A1( u2_u6_X_31 ) , .ZN( u2_u6_u5_n109 ) , .A2( u2_u6_u5_n181 ) );
  INV_X1 u2_u6_u5_U88 (.A( u2_u6_X_33 ) , .ZN( u2_u6_u5_n180 ) );
  INV_X1 u2_u6_u5_U89 (.A( u2_u6_X_35 ) , .ZN( u2_u6_u5_n171 ) );
  NOR2_X1 u2_u6_u5_U9 (.ZN( u2_u6_u5_n135 ) , .A1( u2_u6_u5_n173 ) , .A2( u2_u6_u5_n176 ) );
  INV_X1 u2_u6_u5_U90 (.A( u2_u6_X_36 ) , .ZN( u2_u6_u5_n170 ) );
  INV_X1 u2_u6_u5_U91 (.A( u2_u6_X_32 ) , .ZN( u2_u6_u5_n181 ) );
  NAND4_X1 u2_u6_u5_U92 (.ZN( u2_out6_29 ) , .A4( u2_u6_u5_n129 ) , .A3( u2_u6_u5_n130 ) , .A2( u2_u6_u5_n168 ) , .A1( u2_u6_u5_n196 ) );
  AOI221_X1 u2_u6_u5_U93 (.A( u2_u6_u5_n128 ) , .ZN( u2_u6_u5_n129 ) , .C2( u2_u6_u5_n132 ) , .B2( u2_u6_u5_n159 ) , .B1( u2_u6_u5_n176 ) , .C1( u2_u6_u5_n184 ) );
  AOI222_X1 u2_u6_u5_U94 (.ZN( u2_u6_u5_n130 ) , .A2( u2_u6_u5_n146 ) , .B1( u2_u6_u5_n147 ) , .C2( u2_u6_u5_n175 ) , .B2( u2_u6_u5_n179 ) , .A1( u2_u6_u5_n188 ) , .C1( u2_u6_u5_n194 ) );
  NAND4_X1 u2_u6_u5_U95 (.ZN( u2_out6_19 ) , .A4( u2_u6_u5_n166 ) , .A3( u2_u6_u5_n167 ) , .A2( u2_u6_u5_n168 ) , .A1( u2_u6_u5_n169 ) );
  AOI22_X1 u2_u6_u5_U96 (.B2( u2_u6_u5_n145 ) , .A2( u2_u6_u5_n146 ) , .ZN( u2_u6_u5_n167 ) , .B1( u2_u6_u5_n182 ) , .A1( u2_u6_u5_n189 ) );
  NOR4_X1 u2_u6_u5_U97 (.A4( u2_u6_u5_n162 ) , .A3( u2_u6_u5_n163 ) , .A2( u2_u6_u5_n164 ) , .A1( u2_u6_u5_n165 ) , .ZN( u2_u6_u5_n166 ) );
  NAND4_X1 u2_u6_u5_U98 (.ZN( u2_out6_11 ) , .A4( u2_u6_u5_n143 ) , .A3( u2_u6_u5_n144 ) , .A2( u2_u6_u5_n169 ) , .A1( u2_u6_u5_n196 ) );
  AOI22_X1 u2_u6_u5_U99 (.A2( u2_u6_u5_n132 ) , .ZN( u2_u6_u5_n144 ) , .B2( u2_u6_u5_n145 ) , .B1( u2_u6_u5_n184 ) , .A1( u2_u6_u5_n194 ) );
  AOI21_X1 u2_u6_u6_U10 (.ZN( u2_u6_u6_n106 ) , .A( u2_u6_u6_n142 ) , .B2( u2_u6_u6_n159 ) , .B1( u2_u6_u6_n164 ) );
  INV_X1 u2_u6_u6_U11 (.A( u2_u6_u6_n155 ) , .ZN( u2_u6_u6_n161 ) );
  INV_X1 u2_u6_u6_U12 (.A( u2_u6_u6_n128 ) , .ZN( u2_u6_u6_n164 ) );
  NAND2_X1 u2_u6_u6_U13 (.ZN( u2_u6_u6_n110 ) , .A1( u2_u6_u6_n122 ) , .A2( u2_u6_u6_n129 ) );
  NAND2_X1 u2_u6_u6_U14 (.ZN( u2_u6_u6_n124 ) , .A2( u2_u6_u6_n146 ) , .A1( u2_u6_u6_n148 ) );
  INV_X1 u2_u6_u6_U15 (.A( u2_u6_u6_n132 ) , .ZN( u2_u6_u6_n171 ) );
  AND2_X1 u2_u6_u6_U16 (.A1( u2_u6_u6_n100 ) , .ZN( u2_u6_u6_n130 ) , .A2( u2_u6_u6_n147 ) );
  INV_X1 u2_u6_u6_U17 (.A( u2_u6_u6_n127 ) , .ZN( u2_u6_u6_n173 ) );
  INV_X1 u2_u6_u6_U18 (.A( u2_u6_u6_n121 ) , .ZN( u2_u6_u6_n167 ) );
  INV_X1 u2_u6_u6_U19 (.A( u2_u6_u6_n100 ) , .ZN( u2_u6_u6_n169 ) );
  INV_X1 u2_u6_u6_U20 (.A( u2_u6_u6_n123 ) , .ZN( u2_u6_u6_n170 ) );
  INV_X1 u2_u6_u6_U21 (.A( u2_u6_u6_n113 ) , .ZN( u2_u6_u6_n168 ) );
  AND2_X1 u2_u6_u6_U22 (.A1( u2_u6_u6_n107 ) , .A2( u2_u6_u6_n119 ) , .ZN( u2_u6_u6_n133 ) );
  AND2_X1 u2_u6_u6_U23 (.A2( u2_u6_u6_n121 ) , .A1( u2_u6_u6_n122 ) , .ZN( u2_u6_u6_n131 ) );
  AND3_X1 u2_u6_u6_U24 (.ZN( u2_u6_u6_n120 ) , .A2( u2_u6_u6_n127 ) , .A1( u2_u6_u6_n132 ) , .A3( u2_u6_u6_n145 ) );
  INV_X1 u2_u6_u6_U25 (.A( u2_u6_u6_n146 ) , .ZN( u2_u6_u6_n163 ) );
  AOI222_X1 u2_u6_u6_U26 (.ZN( u2_u6_u6_n114 ) , .A1( u2_u6_u6_n118 ) , .A2( u2_u6_u6_n126 ) , .B2( u2_u6_u6_n151 ) , .C2( u2_u6_u6_n159 ) , .C1( u2_u6_u6_n168 ) , .B1( u2_u6_u6_n169 ) );
  NOR2_X1 u2_u6_u6_U27 (.A1( u2_u6_u6_n162 ) , .A2( u2_u6_u6_n165 ) , .ZN( u2_u6_u6_n98 ) );
  AOI211_X1 u2_u6_u6_U28 (.B( u2_u6_u6_n149 ) , .A( u2_u6_u6_n150 ) , .C2( u2_u6_u6_n151 ) , .C1( u2_u6_u6_n152 ) , .ZN( u2_u6_u6_n153 ) );
  AOI21_X1 u2_u6_u6_U29 (.B2( u2_u6_u6_n147 ) , .B1( u2_u6_u6_n148 ) , .ZN( u2_u6_u6_n149 ) , .A( u2_u6_u6_n158 ) );
  INV_X1 u2_u6_u6_U3 (.A( u2_u6_u6_n110 ) , .ZN( u2_u6_u6_n166 ) );
  AOI21_X1 u2_u6_u6_U30 (.A( u2_u6_u6_n144 ) , .B2( u2_u6_u6_n145 ) , .B1( u2_u6_u6_n146 ) , .ZN( u2_u6_u6_n150 ) );
  NAND2_X1 u2_u6_u6_U31 (.A2( u2_u6_u6_n143 ) , .ZN( u2_u6_u6_n152 ) , .A1( u2_u6_u6_n166 ) );
  NAND2_X1 u2_u6_u6_U32 (.A1( u2_u6_u6_n144 ) , .ZN( u2_u6_u6_n151 ) , .A2( u2_u6_u6_n158 ) );
  NAND2_X1 u2_u6_u6_U33 (.ZN( u2_u6_u6_n132 ) , .A1( u2_u6_u6_n91 ) , .A2( u2_u6_u6_n97 ) );
  AOI22_X1 u2_u6_u6_U34 (.B2( u2_u6_u6_n110 ) , .B1( u2_u6_u6_n111 ) , .A1( u2_u6_u6_n112 ) , .ZN( u2_u6_u6_n115 ) , .A2( u2_u6_u6_n161 ) );
  NAND4_X1 u2_u6_u6_U35 (.A3( u2_u6_u6_n109 ) , .ZN( u2_u6_u6_n112 ) , .A4( u2_u6_u6_n132 ) , .A2( u2_u6_u6_n147 ) , .A1( u2_u6_u6_n166 ) );
  NOR2_X1 u2_u6_u6_U36 (.ZN( u2_u6_u6_n109 ) , .A1( u2_u6_u6_n170 ) , .A2( u2_u6_u6_n173 ) );
  NOR2_X1 u2_u6_u6_U37 (.A2( u2_u6_u6_n126 ) , .ZN( u2_u6_u6_n155 ) , .A1( u2_u6_u6_n160 ) );
  NAND2_X1 u2_u6_u6_U38 (.ZN( u2_u6_u6_n146 ) , .A2( u2_u6_u6_n94 ) , .A1( u2_u6_u6_n99 ) );
  AOI211_X1 u2_u6_u6_U39 (.B( u2_u6_u6_n134 ) , .A( u2_u6_u6_n135 ) , .C1( u2_u6_u6_n136 ) , .ZN( u2_u6_u6_n137 ) , .C2( u2_u6_u6_n151 ) );
  AOI22_X1 u2_u6_u6_U4 (.B2( u2_u6_u6_n101 ) , .A1( u2_u6_u6_n102 ) , .ZN( u2_u6_u6_n103 ) , .B1( u2_u6_u6_n160 ) , .A2( u2_u6_u6_n161 ) );
  NAND4_X1 u2_u6_u6_U40 (.A4( u2_u6_u6_n127 ) , .A3( u2_u6_u6_n128 ) , .A2( u2_u6_u6_n129 ) , .A1( u2_u6_u6_n130 ) , .ZN( u2_u6_u6_n136 ) );
  AOI21_X1 u2_u6_u6_U41 (.B2( u2_u6_u6_n132 ) , .B1( u2_u6_u6_n133 ) , .ZN( u2_u6_u6_n134 ) , .A( u2_u6_u6_n158 ) );
  AOI21_X1 u2_u6_u6_U42 (.B1( u2_u6_u6_n131 ) , .ZN( u2_u6_u6_n135 ) , .A( u2_u6_u6_n144 ) , .B2( u2_u6_u6_n146 ) );
  INV_X1 u2_u6_u6_U43 (.A( u2_u6_u6_n111 ) , .ZN( u2_u6_u6_n158 ) );
  NAND2_X1 u2_u6_u6_U44 (.ZN( u2_u6_u6_n127 ) , .A1( u2_u6_u6_n91 ) , .A2( u2_u6_u6_n92 ) );
  NAND2_X1 u2_u6_u6_U45 (.ZN( u2_u6_u6_n129 ) , .A2( u2_u6_u6_n95 ) , .A1( u2_u6_u6_n96 ) );
  INV_X1 u2_u6_u6_U46 (.A( u2_u6_u6_n144 ) , .ZN( u2_u6_u6_n159 ) );
  NAND2_X1 u2_u6_u6_U47 (.ZN( u2_u6_u6_n145 ) , .A2( u2_u6_u6_n97 ) , .A1( u2_u6_u6_n98 ) );
  NAND2_X1 u2_u6_u6_U48 (.ZN( u2_u6_u6_n148 ) , .A2( u2_u6_u6_n92 ) , .A1( u2_u6_u6_n94 ) );
  NAND2_X1 u2_u6_u6_U49 (.ZN( u2_u6_u6_n108 ) , .A2( u2_u6_u6_n139 ) , .A1( u2_u6_u6_n144 ) );
  NOR2_X1 u2_u6_u6_U5 (.A1( u2_u6_u6_n118 ) , .ZN( u2_u6_u6_n143 ) , .A2( u2_u6_u6_n168 ) );
  NAND2_X1 u2_u6_u6_U50 (.ZN( u2_u6_u6_n121 ) , .A2( u2_u6_u6_n95 ) , .A1( u2_u6_u6_n97 ) );
  NAND2_X1 u2_u6_u6_U51 (.ZN( u2_u6_u6_n107 ) , .A2( u2_u6_u6_n92 ) , .A1( u2_u6_u6_n95 ) );
  AND2_X1 u2_u6_u6_U52 (.ZN( u2_u6_u6_n118 ) , .A2( u2_u6_u6_n91 ) , .A1( u2_u6_u6_n99 ) );
  NAND2_X1 u2_u6_u6_U53 (.ZN( u2_u6_u6_n147 ) , .A2( u2_u6_u6_n98 ) , .A1( u2_u6_u6_n99 ) );
  NAND2_X1 u2_u6_u6_U54 (.ZN( u2_u6_u6_n128 ) , .A1( u2_u6_u6_n94 ) , .A2( u2_u6_u6_n96 ) );
  NAND2_X1 u2_u6_u6_U55 (.ZN( u2_u6_u6_n119 ) , .A2( u2_u6_u6_n95 ) , .A1( u2_u6_u6_n99 ) );
  NAND2_X1 u2_u6_u6_U56 (.ZN( u2_u6_u6_n123 ) , .A2( u2_u6_u6_n91 ) , .A1( u2_u6_u6_n96 ) );
  NAND2_X1 u2_u6_u6_U57 (.ZN( u2_u6_u6_n100 ) , .A2( u2_u6_u6_n92 ) , .A1( u2_u6_u6_n98 ) );
  NAND2_X1 u2_u6_u6_U58 (.ZN( u2_u6_u6_n122 ) , .A1( u2_u6_u6_n94 ) , .A2( u2_u6_u6_n97 ) );
  INV_X1 u2_u6_u6_U59 (.A( u2_u6_u6_n139 ) , .ZN( u2_u6_u6_n160 ) );
  AOI21_X1 u2_u6_u6_U6 (.B1( u2_u6_u6_n107 ) , .B2( u2_u6_u6_n132 ) , .A( u2_u6_u6_n158 ) , .ZN( u2_u6_u6_n88 ) );
  NAND2_X1 u2_u6_u6_U60 (.ZN( u2_u6_u6_n113 ) , .A1( u2_u6_u6_n96 ) , .A2( u2_u6_u6_n98 ) );
  NOR2_X1 u2_u6_u6_U61 (.A2( u2_u6_X_40 ) , .A1( u2_u6_X_41 ) , .ZN( u2_u6_u6_n126 ) );
  NOR2_X1 u2_u6_u6_U62 (.A2( u2_u6_X_39 ) , .A1( u2_u6_X_42 ) , .ZN( u2_u6_u6_n92 ) );
  NOR2_X1 u2_u6_u6_U63 (.A2( u2_u6_X_39 ) , .A1( u2_u6_u6_n156 ) , .ZN( u2_u6_u6_n97 ) );
  NOR2_X1 u2_u6_u6_U64 (.A2( u2_u6_X_38 ) , .A1( u2_u6_u6_n165 ) , .ZN( u2_u6_u6_n95 ) );
  NOR2_X1 u2_u6_u6_U65 (.A2( u2_u6_X_41 ) , .ZN( u2_u6_u6_n111 ) , .A1( u2_u6_u6_n157 ) );
  NOR2_X1 u2_u6_u6_U66 (.A2( u2_u6_X_37 ) , .A1( u2_u6_u6_n162 ) , .ZN( u2_u6_u6_n94 ) );
  NOR2_X1 u2_u6_u6_U67 (.A2( u2_u6_X_37 ) , .A1( u2_u6_X_38 ) , .ZN( u2_u6_u6_n91 ) );
  NAND2_X1 u2_u6_u6_U68 (.A1( u2_u6_X_41 ) , .ZN( u2_u6_u6_n144 ) , .A2( u2_u6_u6_n157 ) );
  NAND2_X1 u2_u6_u6_U69 (.A2( u2_u6_X_40 ) , .A1( u2_u6_X_41 ) , .ZN( u2_u6_u6_n139 ) );
  OAI21_X1 u2_u6_u6_U7 (.A( u2_u6_u6_n159 ) , .B1( u2_u6_u6_n169 ) , .B2( u2_u6_u6_n173 ) , .ZN( u2_u6_u6_n90 ) );
  AND2_X1 u2_u6_u6_U70 (.A1( u2_u6_X_39 ) , .A2( u2_u6_u6_n156 ) , .ZN( u2_u6_u6_n96 ) );
  AND2_X1 u2_u6_u6_U71 (.A1( u2_u6_X_39 ) , .A2( u2_u6_X_42 ) , .ZN( u2_u6_u6_n99 ) );
  INV_X1 u2_u6_u6_U72 (.A( u2_u6_X_40 ) , .ZN( u2_u6_u6_n157 ) );
  INV_X1 u2_u6_u6_U73 (.A( u2_u6_X_37 ) , .ZN( u2_u6_u6_n165 ) );
  INV_X1 u2_u6_u6_U74 (.A( u2_u6_X_38 ) , .ZN( u2_u6_u6_n162 ) );
  INV_X1 u2_u6_u6_U75 (.A( u2_u6_X_42 ) , .ZN( u2_u6_u6_n156 ) );
  NAND4_X1 u2_u6_u6_U76 (.ZN( u2_out6_32 ) , .A4( u2_u6_u6_n103 ) , .A3( u2_u6_u6_n104 ) , .A2( u2_u6_u6_n105 ) , .A1( u2_u6_u6_n106 ) );
  AOI22_X1 u2_u6_u6_U77 (.ZN( u2_u6_u6_n104 ) , .A1( u2_u6_u6_n111 ) , .B1( u2_u6_u6_n124 ) , .B2( u2_u6_u6_n151 ) , .A2( u2_u6_u6_n93 ) );
  AOI22_X1 u2_u6_u6_U78 (.ZN( u2_u6_u6_n105 ) , .A2( u2_u6_u6_n108 ) , .A1( u2_u6_u6_n118 ) , .B2( u2_u6_u6_n126 ) , .B1( u2_u6_u6_n171 ) );
  NAND4_X1 u2_u6_u6_U79 (.ZN( u2_out6_12 ) , .A4( u2_u6_u6_n114 ) , .A3( u2_u6_u6_n115 ) , .A2( u2_u6_u6_n116 ) , .A1( u2_u6_u6_n117 ) );
  INV_X1 u2_u6_u6_U8 (.ZN( u2_u6_u6_n172 ) , .A( u2_u6_u6_n88 ) );
  OAI22_X1 u2_u6_u6_U80 (.B2( u2_u6_u6_n111 ) , .ZN( u2_u6_u6_n116 ) , .B1( u2_u6_u6_n126 ) , .A2( u2_u6_u6_n164 ) , .A1( u2_u6_u6_n167 ) );
  OAI21_X1 u2_u6_u6_U81 (.A( u2_u6_u6_n108 ) , .ZN( u2_u6_u6_n117 ) , .B2( u2_u6_u6_n141 ) , .B1( u2_u6_u6_n163 ) );
  OAI211_X1 u2_u6_u6_U82 (.ZN( u2_out6_22 ) , .B( u2_u6_u6_n137 ) , .A( u2_u6_u6_n138 ) , .C2( u2_u6_u6_n139 ) , .C1( u2_u6_u6_n140 ) );
  AOI22_X1 u2_u6_u6_U83 (.B1( u2_u6_u6_n124 ) , .A2( u2_u6_u6_n125 ) , .A1( u2_u6_u6_n126 ) , .ZN( u2_u6_u6_n138 ) , .B2( u2_u6_u6_n161 ) );
  AND4_X1 u2_u6_u6_U84 (.A3( u2_u6_u6_n119 ) , .A1( u2_u6_u6_n120 ) , .A4( u2_u6_u6_n129 ) , .ZN( u2_u6_u6_n140 ) , .A2( u2_u6_u6_n143 ) );
  OAI211_X1 u2_u6_u6_U85 (.ZN( u2_out6_7 ) , .B( u2_u6_u6_n153 ) , .C2( u2_u6_u6_n154 ) , .C1( u2_u6_u6_n155 ) , .A( u2_u6_u6_n174 ) );
  NOR3_X1 u2_u6_u6_U86 (.A1( u2_u6_u6_n141 ) , .ZN( u2_u6_u6_n154 ) , .A3( u2_u6_u6_n164 ) , .A2( u2_u6_u6_n171 ) );
  INV_X1 u2_u6_u6_U87 (.A( u2_u6_u6_n142 ) , .ZN( u2_u6_u6_n174 ) );
  NAND3_X1 u2_u6_u6_U88 (.A2( u2_u6_u6_n123 ) , .ZN( u2_u6_u6_n125 ) , .A1( u2_u6_u6_n130 ) , .A3( u2_u6_u6_n131 ) );
  NAND3_X1 u2_u6_u6_U89 (.A3( u2_u6_u6_n133 ) , .ZN( u2_u6_u6_n141 ) , .A1( u2_u6_u6_n145 ) , .A2( u2_u6_u6_n148 ) );
  AOI22_X1 u2_u6_u6_U9 (.A2( u2_u6_u6_n151 ) , .B2( u2_u6_u6_n161 ) , .A1( u2_u6_u6_n167 ) , .B1( u2_u6_u6_n170 ) , .ZN( u2_u6_u6_n89 ) );
  NAND3_X1 u2_u6_u6_U90 (.ZN( u2_u6_u6_n101 ) , .A3( u2_u6_u6_n107 ) , .A2( u2_u6_u6_n121 ) , .A1( u2_u6_u6_n127 ) );
  NAND3_X1 u2_u6_u6_U91 (.ZN( u2_u6_u6_n102 ) , .A3( u2_u6_u6_n130 ) , .A2( u2_u6_u6_n145 ) , .A1( u2_u6_u6_n166 ) );
  NAND3_X1 u2_u6_u6_U92 (.A3( u2_u6_u6_n113 ) , .A1( u2_u6_u6_n119 ) , .A2( u2_u6_u6_n123 ) , .ZN( u2_u6_u6_n93 ) );
  NAND3_X1 u2_u6_u6_U93 (.ZN( u2_u6_u6_n142 ) , .A2( u2_u6_u6_n172 ) , .A3( u2_u6_u6_n89 ) , .A1( u2_u6_u6_n90 ) );
  AND3_X1 u2_u6_u7_U10 (.A3( u2_u6_u7_n110 ) , .A2( u2_u6_u7_n127 ) , .A1( u2_u6_u7_n132 ) , .ZN( u2_u6_u7_n92 ) );
  OAI21_X1 u2_u6_u7_U11 (.A( u2_u6_u7_n161 ) , .B1( u2_u6_u7_n168 ) , .B2( u2_u6_u7_n173 ) , .ZN( u2_u6_u7_n91 ) );
  AOI211_X1 u2_u6_u7_U12 (.A( u2_u6_u7_n117 ) , .ZN( u2_u6_u7_n118 ) , .C2( u2_u6_u7_n126 ) , .C1( u2_u6_u7_n177 ) , .B( u2_u6_u7_n180 ) );
  OAI22_X1 u2_u6_u7_U13 (.B1( u2_u6_u7_n115 ) , .ZN( u2_u6_u7_n117 ) , .A2( u2_u6_u7_n133 ) , .A1( u2_u6_u7_n137 ) , .B2( u2_u6_u7_n162 ) );
  INV_X1 u2_u6_u7_U14 (.A( u2_u6_u7_n116 ) , .ZN( u2_u6_u7_n180 ) );
  NOR3_X1 u2_u6_u7_U15 (.ZN( u2_u6_u7_n115 ) , .A3( u2_u6_u7_n145 ) , .A2( u2_u6_u7_n168 ) , .A1( u2_u6_u7_n169 ) );
  OAI211_X1 u2_u6_u7_U16 (.B( u2_u6_u7_n122 ) , .A( u2_u6_u7_n123 ) , .C2( u2_u6_u7_n124 ) , .ZN( u2_u6_u7_n154 ) , .C1( u2_u6_u7_n162 ) );
  AOI222_X1 u2_u6_u7_U17 (.ZN( u2_u6_u7_n122 ) , .C2( u2_u6_u7_n126 ) , .C1( u2_u6_u7_n145 ) , .B1( u2_u6_u7_n161 ) , .A2( u2_u6_u7_n165 ) , .B2( u2_u6_u7_n170 ) , .A1( u2_u6_u7_n176 ) );
  INV_X1 u2_u6_u7_U18 (.A( u2_u6_u7_n133 ) , .ZN( u2_u6_u7_n176 ) );
  NOR3_X1 u2_u6_u7_U19 (.A2( u2_u6_u7_n134 ) , .A1( u2_u6_u7_n135 ) , .ZN( u2_u6_u7_n136 ) , .A3( u2_u6_u7_n171 ) );
  NOR2_X1 u2_u6_u7_U20 (.A1( u2_u6_u7_n130 ) , .A2( u2_u6_u7_n134 ) , .ZN( u2_u6_u7_n153 ) );
  INV_X1 u2_u6_u7_U21 (.A( u2_u6_u7_n101 ) , .ZN( u2_u6_u7_n165 ) );
  NOR2_X1 u2_u6_u7_U22 (.ZN( u2_u6_u7_n111 ) , .A2( u2_u6_u7_n134 ) , .A1( u2_u6_u7_n169 ) );
  AOI21_X1 u2_u6_u7_U23 (.ZN( u2_u6_u7_n104 ) , .B2( u2_u6_u7_n112 ) , .B1( u2_u6_u7_n127 ) , .A( u2_u6_u7_n164 ) );
  AOI21_X1 u2_u6_u7_U24 (.ZN( u2_u6_u7_n106 ) , .B1( u2_u6_u7_n133 ) , .B2( u2_u6_u7_n146 ) , .A( u2_u6_u7_n162 ) );
  AOI21_X1 u2_u6_u7_U25 (.A( u2_u6_u7_n101 ) , .ZN( u2_u6_u7_n107 ) , .B2( u2_u6_u7_n128 ) , .B1( u2_u6_u7_n175 ) );
  INV_X1 u2_u6_u7_U26 (.A( u2_u6_u7_n138 ) , .ZN( u2_u6_u7_n171 ) );
  INV_X1 u2_u6_u7_U27 (.A( u2_u6_u7_n131 ) , .ZN( u2_u6_u7_n177 ) );
  INV_X1 u2_u6_u7_U28 (.A( u2_u6_u7_n110 ) , .ZN( u2_u6_u7_n174 ) );
  NAND2_X1 u2_u6_u7_U29 (.A1( u2_u6_u7_n129 ) , .A2( u2_u6_u7_n132 ) , .ZN( u2_u6_u7_n149 ) );
  OAI21_X1 u2_u6_u7_U3 (.ZN( u2_u6_u7_n159 ) , .A( u2_u6_u7_n165 ) , .B2( u2_u6_u7_n171 ) , .B1( u2_u6_u7_n174 ) );
  NAND2_X1 u2_u6_u7_U30 (.A1( u2_u6_u7_n113 ) , .A2( u2_u6_u7_n124 ) , .ZN( u2_u6_u7_n130 ) );
  INV_X1 u2_u6_u7_U31 (.A( u2_u6_u7_n112 ) , .ZN( u2_u6_u7_n173 ) );
  INV_X1 u2_u6_u7_U32 (.A( u2_u6_u7_n128 ) , .ZN( u2_u6_u7_n168 ) );
  INV_X1 u2_u6_u7_U33 (.A( u2_u6_u7_n148 ) , .ZN( u2_u6_u7_n169 ) );
  INV_X1 u2_u6_u7_U34 (.A( u2_u6_u7_n127 ) , .ZN( u2_u6_u7_n179 ) );
  NOR2_X1 u2_u6_u7_U35 (.ZN( u2_u6_u7_n101 ) , .A2( u2_u6_u7_n150 ) , .A1( u2_u6_u7_n156 ) );
  AOI211_X1 u2_u6_u7_U36 (.B( u2_u6_u7_n154 ) , .A( u2_u6_u7_n155 ) , .C1( u2_u6_u7_n156 ) , .ZN( u2_u6_u7_n157 ) , .C2( u2_u6_u7_n172 ) );
  INV_X1 u2_u6_u7_U37 (.A( u2_u6_u7_n153 ) , .ZN( u2_u6_u7_n172 ) );
  AOI211_X1 u2_u6_u7_U38 (.B( u2_u6_u7_n139 ) , .A( u2_u6_u7_n140 ) , .C2( u2_u6_u7_n141 ) , .ZN( u2_u6_u7_n142 ) , .C1( u2_u6_u7_n156 ) );
  NAND4_X1 u2_u6_u7_U39 (.A3( u2_u6_u7_n127 ) , .A2( u2_u6_u7_n128 ) , .A1( u2_u6_u7_n129 ) , .ZN( u2_u6_u7_n141 ) , .A4( u2_u6_u7_n147 ) );
  INV_X1 u2_u6_u7_U4 (.A( u2_u6_u7_n111 ) , .ZN( u2_u6_u7_n170 ) );
  AOI21_X1 u2_u6_u7_U40 (.A( u2_u6_u7_n137 ) , .B1( u2_u6_u7_n138 ) , .ZN( u2_u6_u7_n139 ) , .B2( u2_u6_u7_n146 ) );
  OAI22_X1 u2_u6_u7_U41 (.B1( u2_u6_u7_n136 ) , .ZN( u2_u6_u7_n140 ) , .A1( u2_u6_u7_n153 ) , .B2( u2_u6_u7_n162 ) , .A2( u2_u6_u7_n164 ) );
  AOI21_X1 u2_u6_u7_U42 (.ZN( u2_u6_u7_n123 ) , .B1( u2_u6_u7_n165 ) , .B2( u2_u6_u7_n177 ) , .A( u2_u6_u7_n97 ) );
  AOI21_X1 u2_u6_u7_U43 (.B2( u2_u6_u7_n113 ) , .B1( u2_u6_u7_n124 ) , .A( u2_u6_u7_n125 ) , .ZN( u2_u6_u7_n97 ) );
  INV_X1 u2_u6_u7_U44 (.A( u2_u6_u7_n125 ) , .ZN( u2_u6_u7_n161 ) );
  INV_X1 u2_u6_u7_U45 (.A( u2_u6_u7_n152 ) , .ZN( u2_u6_u7_n162 ) );
  AOI22_X1 u2_u6_u7_U46 (.A2( u2_u6_u7_n114 ) , .ZN( u2_u6_u7_n119 ) , .B1( u2_u6_u7_n130 ) , .A1( u2_u6_u7_n156 ) , .B2( u2_u6_u7_n165 ) );
  NAND2_X1 u2_u6_u7_U47 (.A2( u2_u6_u7_n112 ) , .ZN( u2_u6_u7_n114 ) , .A1( u2_u6_u7_n175 ) );
  AND2_X1 u2_u6_u7_U48 (.ZN( u2_u6_u7_n145 ) , .A2( u2_u6_u7_n98 ) , .A1( u2_u6_u7_n99 ) );
  NOR2_X1 u2_u6_u7_U49 (.ZN( u2_u6_u7_n137 ) , .A1( u2_u6_u7_n150 ) , .A2( u2_u6_u7_n161 ) );
  INV_X1 u2_u6_u7_U5 (.A( u2_u6_u7_n149 ) , .ZN( u2_u6_u7_n175 ) );
  AOI21_X1 u2_u6_u7_U50 (.ZN( u2_u6_u7_n105 ) , .B2( u2_u6_u7_n110 ) , .A( u2_u6_u7_n125 ) , .B1( u2_u6_u7_n147 ) );
  NAND2_X1 u2_u6_u7_U51 (.ZN( u2_u6_u7_n146 ) , .A1( u2_u6_u7_n95 ) , .A2( u2_u6_u7_n98 ) );
  NAND2_X1 u2_u6_u7_U52 (.A2( u2_u6_u7_n103 ) , .ZN( u2_u6_u7_n147 ) , .A1( u2_u6_u7_n93 ) );
  NAND2_X1 u2_u6_u7_U53 (.A1( u2_u6_u7_n103 ) , .ZN( u2_u6_u7_n127 ) , .A2( u2_u6_u7_n99 ) );
  OR2_X1 u2_u6_u7_U54 (.ZN( u2_u6_u7_n126 ) , .A2( u2_u6_u7_n152 ) , .A1( u2_u6_u7_n156 ) );
  NAND2_X1 u2_u6_u7_U55 (.A2( u2_u6_u7_n102 ) , .A1( u2_u6_u7_n103 ) , .ZN( u2_u6_u7_n133 ) );
  NAND2_X1 u2_u6_u7_U56 (.ZN( u2_u6_u7_n112 ) , .A2( u2_u6_u7_n96 ) , .A1( u2_u6_u7_n99 ) );
  NAND2_X1 u2_u6_u7_U57 (.A2( u2_u6_u7_n102 ) , .ZN( u2_u6_u7_n128 ) , .A1( u2_u6_u7_n98 ) );
  NAND2_X1 u2_u6_u7_U58 (.A1( u2_u6_u7_n100 ) , .ZN( u2_u6_u7_n113 ) , .A2( u2_u6_u7_n93 ) );
  NAND2_X1 u2_u6_u7_U59 (.A2( u2_u6_u7_n102 ) , .ZN( u2_u6_u7_n124 ) , .A1( u2_u6_u7_n96 ) );
  INV_X1 u2_u6_u7_U6 (.A( u2_u6_u7_n154 ) , .ZN( u2_u6_u7_n178 ) );
  NAND2_X1 u2_u6_u7_U60 (.ZN( u2_u6_u7_n110 ) , .A1( u2_u6_u7_n95 ) , .A2( u2_u6_u7_n96 ) );
  INV_X1 u2_u6_u7_U61 (.A( u2_u6_u7_n150 ) , .ZN( u2_u6_u7_n164 ) );
  AND2_X1 u2_u6_u7_U62 (.ZN( u2_u6_u7_n134 ) , .A1( u2_u6_u7_n93 ) , .A2( u2_u6_u7_n98 ) );
  NAND2_X1 u2_u6_u7_U63 (.A1( u2_u6_u7_n100 ) , .A2( u2_u6_u7_n102 ) , .ZN( u2_u6_u7_n129 ) );
  NAND2_X1 u2_u6_u7_U64 (.A2( u2_u6_u7_n103 ) , .ZN( u2_u6_u7_n131 ) , .A1( u2_u6_u7_n95 ) );
  NAND2_X1 u2_u6_u7_U65 (.A1( u2_u6_u7_n100 ) , .ZN( u2_u6_u7_n138 ) , .A2( u2_u6_u7_n99 ) );
  NAND2_X1 u2_u6_u7_U66 (.ZN( u2_u6_u7_n132 ) , .A1( u2_u6_u7_n93 ) , .A2( u2_u6_u7_n96 ) );
  NAND2_X1 u2_u6_u7_U67 (.A1( u2_u6_u7_n100 ) , .ZN( u2_u6_u7_n148 ) , .A2( u2_u6_u7_n95 ) );
  NOR2_X1 u2_u6_u7_U68 (.A2( u2_u6_X_47 ) , .ZN( u2_u6_u7_n150 ) , .A1( u2_u6_u7_n163 ) );
  NOR2_X1 u2_u6_u7_U69 (.A2( u2_u6_X_43 ) , .A1( u2_u6_X_44 ) , .ZN( u2_u6_u7_n103 ) );
  AOI211_X1 u2_u6_u7_U7 (.ZN( u2_u6_u7_n116 ) , .A( u2_u6_u7_n155 ) , .C1( u2_u6_u7_n161 ) , .C2( u2_u6_u7_n171 ) , .B( u2_u6_u7_n94 ) );
  NOR2_X1 u2_u6_u7_U70 (.A2( u2_u6_X_48 ) , .A1( u2_u6_u7_n166 ) , .ZN( u2_u6_u7_n95 ) );
  NOR2_X1 u2_u6_u7_U71 (.A2( u2_u6_X_45 ) , .A1( u2_u6_X_48 ) , .ZN( u2_u6_u7_n99 ) );
  NOR2_X1 u2_u6_u7_U72 (.A2( u2_u6_X_44 ) , .A1( u2_u6_u7_n167 ) , .ZN( u2_u6_u7_n98 ) );
  NOR2_X1 u2_u6_u7_U73 (.A2( u2_u6_X_46 ) , .A1( u2_u6_X_47 ) , .ZN( u2_u6_u7_n152 ) );
  AND2_X1 u2_u6_u7_U74 (.A1( u2_u6_X_47 ) , .ZN( u2_u6_u7_n156 ) , .A2( u2_u6_u7_n163 ) );
  NAND2_X1 u2_u6_u7_U75 (.A2( u2_u6_X_46 ) , .A1( u2_u6_X_47 ) , .ZN( u2_u6_u7_n125 ) );
  AND2_X1 u2_u6_u7_U76 (.A2( u2_u6_X_45 ) , .A1( u2_u6_X_48 ) , .ZN( u2_u6_u7_n102 ) );
  AND2_X1 u2_u6_u7_U77 (.A2( u2_u6_X_43 ) , .A1( u2_u6_X_44 ) , .ZN( u2_u6_u7_n96 ) );
  AND2_X1 u2_u6_u7_U78 (.A1( u2_u6_X_44 ) , .ZN( u2_u6_u7_n100 ) , .A2( u2_u6_u7_n167 ) );
  AND2_X1 u2_u6_u7_U79 (.A1( u2_u6_X_48 ) , .A2( u2_u6_u7_n166 ) , .ZN( u2_u6_u7_n93 ) );
  OAI222_X1 u2_u6_u7_U8 (.C2( u2_u6_u7_n101 ) , .B2( u2_u6_u7_n111 ) , .A1( u2_u6_u7_n113 ) , .C1( u2_u6_u7_n146 ) , .A2( u2_u6_u7_n162 ) , .B1( u2_u6_u7_n164 ) , .ZN( u2_u6_u7_n94 ) );
  INV_X1 u2_u6_u7_U80 (.A( u2_u6_X_46 ) , .ZN( u2_u6_u7_n163 ) );
  INV_X1 u2_u6_u7_U81 (.A( u2_u6_X_43 ) , .ZN( u2_u6_u7_n167 ) );
  INV_X1 u2_u6_u7_U82 (.A( u2_u6_X_45 ) , .ZN( u2_u6_u7_n166 ) );
  NAND4_X1 u2_u6_u7_U83 (.ZN( u2_out6_5 ) , .A4( u2_u6_u7_n108 ) , .A3( u2_u6_u7_n109 ) , .A1( u2_u6_u7_n116 ) , .A2( u2_u6_u7_n123 ) );
  AOI22_X1 u2_u6_u7_U84 (.ZN( u2_u6_u7_n109 ) , .A2( u2_u6_u7_n126 ) , .B2( u2_u6_u7_n145 ) , .B1( u2_u6_u7_n156 ) , .A1( u2_u6_u7_n171 ) );
  NOR4_X1 u2_u6_u7_U85 (.A4( u2_u6_u7_n104 ) , .A3( u2_u6_u7_n105 ) , .A2( u2_u6_u7_n106 ) , .A1( u2_u6_u7_n107 ) , .ZN( u2_u6_u7_n108 ) );
  NAND4_X1 u2_u6_u7_U86 (.ZN( u2_out6_27 ) , .A4( u2_u6_u7_n118 ) , .A3( u2_u6_u7_n119 ) , .A2( u2_u6_u7_n120 ) , .A1( u2_u6_u7_n121 ) );
  OAI21_X1 u2_u6_u7_U87 (.ZN( u2_u6_u7_n121 ) , .B2( u2_u6_u7_n145 ) , .A( u2_u6_u7_n150 ) , .B1( u2_u6_u7_n174 ) );
  OAI21_X1 u2_u6_u7_U88 (.ZN( u2_u6_u7_n120 ) , .A( u2_u6_u7_n161 ) , .B2( u2_u6_u7_n170 ) , .B1( u2_u6_u7_n179 ) );
  NAND4_X1 u2_u6_u7_U89 (.ZN( u2_out6_21 ) , .A4( u2_u6_u7_n157 ) , .A3( u2_u6_u7_n158 ) , .A2( u2_u6_u7_n159 ) , .A1( u2_u6_u7_n160 ) );
  OAI221_X1 u2_u6_u7_U9 (.C1( u2_u6_u7_n101 ) , .C2( u2_u6_u7_n147 ) , .ZN( u2_u6_u7_n155 ) , .B2( u2_u6_u7_n162 ) , .A( u2_u6_u7_n91 ) , .B1( u2_u6_u7_n92 ) );
  OAI21_X1 u2_u6_u7_U90 (.B1( u2_u6_u7_n145 ) , .ZN( u2_u6_u7_n160 ) , .A( u2_u6_u7_n161 ) , .B2( u2_u6_u7_n177 ) );
  AOI22_X1 u2_u6_u7_U91 (.B2( u2_u6_u7_n149 ) , .B1( u2_u6_u7_n150 ) , .A2( u2_u6_u7_n151 ) , .A1( u2_u6_u7_n152 ) , .ZN( u2_u6_u7_n158 ) );
  NAND4_X1 u2_u6_u7_U92 (.ZN( u2_out6_15 ) , .A4( u2_u6_u7_n142 ) , .A3( u2_u6_u7_n143 ) , .A2( u2_u6_u7_n144 ) , .A1( u2_u6_u7_n178 ) );
  OR2_X1 u2_u6_u7_U93 (.A2( u2_u6_u7_n125 ) , .A1( u2_u6_u7_n129 ) , .ZN( u2_u6_u7_n144 ) );
  AOI22_X1 u2_u6_u7_U94 (.A2( u2_u6_u7_n126 ) , .ZN( u2_u6_u7_n143 ) , .B2( u2_u6_u7_n165 ) , .B1( u2_u6_u7_n173 ) , .A1( u2_u6_u7_n174 ) );
  NAND3_X1 u2_u6_u7_U95 (.A3( u2_u6_u7_n146 ) , .A2( u2_u6_u7_n147 ) , .A1( u2_u6_u7_n148 ) , .ZN( u2_u6_u7_n151 ) );
  NAND3_X1 u2_u6_u7_U96 (.A3( u2_u6_u7_n131 ) , .A2( u2_u6_u7_n132 ) , .A1( u2_u6_u7_n133 ) , .ZN( u2_u6_u7_n135 ) );
  XOR2_X1 u2_u8_U1 (.B( u2_K9_9 ) , .A( u2_R7_6 ) , .Z( u2_u8_X_9 ) );
  XOR2_X1 u2_u8_U2 (.B( u2_K9_8 ) , .A( u2_R7_5 ) , .Z( u2_u8_X_8 ) );
  XOR2_X1 u2_u8_U27 (.B( u2_K9_2 ) , .A( u2_R7_1 ) , .Z( u2_u8_X_2 ) );
  XOR2_X1 u2_u8_U3 (.B( u2_K9_7 ) , .A( u2_R7_4 ) , .Z( u2_u8_X_7 ) );
  XOR2_X1 u2_u8_U31 (.B( u2_K9_26 ) , .A( u2_R7_17 ) , .Z( u2_u8_X_26 ) );
  XOR2_X1 u2_u8_U32 (.B( u2_K9_25 ) , .A( u2_R7_16 ) , .Z( u2_u8_X_25 ) );
  XOR2_X1 u2_u8_U33 (.B( u2_K9_24 ) , .A( u2_R7_17 ) , .Z( u2_u8_X_24 ) );
  XOR2_X1 u2_u8_U34 (.B( u2_K9_23 ) , .A( u2_R7_16 ) , .Z( u2_u8_X_23 ) );
  XOR2_X1 u2_u8_U35 (.B( u2_K9_22 ) , .A( u2_R7_15 ) , .Z( u2_u8_X_22 ) );
  XOR2_X1 u2_u8_U36 (.B( u2_K9_21 ) , .A( u2_R7_14 ) , .Z( u2_u8_X_21 ) );
  XOR2_X1 u2_u8_U37 (.B( u2_K9_20 ) , .A( u2_R7_13 ) , .Z( u2_u8_X_20 ) );
  XOR2_X1 u2_u8_U39 (.B( u2_K9_19 ) , .A( u2_R7_12 ) , .Z( u2_u8_X_19 ) );
  XOR2_X1 u2_u8_U4 (.B( u2_K9_6 ) , .A( u2_R7_5 ) , .Z( u2_u8_X_6 ) );
  XOR2_X1 u2_u8_U40 (.B( u2_K9_18 ) , .A( u2_R7_13 ) , .Z( u2_u8_X_18 ) );
  XOR2_X1 u2_u8_U41 (.B( u2_K9_17 ) , .A( u2_R7_12 ) , .Z( u2_u8_X_17 ) );
  XOR2_X1 u2_u8_U42 (.B( u2_K9_16 ) , .A( u2_R7_11 ) , .Z( u2_u8_X_16 ) );
  XOR2_X1 u2_u8_U44 (.B( u2_K9_14 ) , .A( u2_R7_9 ) , .Z( u2_u8_X_14 ) );
  XOR2_X1 u2_u8_U45 (.B( u2_K9_13 ) , .A( u2_R7_8 ) , .Z( u2_u8_X_13 ) );
  XOR2_X1 u2_u8_U46 (.B( u2_K9_12 ) , .A( u2_R7_9 ) , .Z( u2_u8_X_12 ) );
  XOR2_X1 u2_u8_U47 (.B( u2_K9_11 ) , .A( u2_R7_8 ) , .Z( u2_u8_X_11 ) );
  XOR2_X1 u2_u8_U48 (.B( u2_K9_10 ) , .A( u2_R7_7 ) , .Z( u2_u8_X_10 ) );
  XOR2_X1 u2_u8_U5 (.B( u2_K9_5 ) , .A( u2_R7_4 ) , .Z( u2_u8_X_5 ) );
  XOR2_X1 u2_u8_U6 (.B( u2_K9_4 ) , .A( u2_R7_3 ) , .Z( u2_u8_X_4 ) );
  AND2_X1 u2_u8_u0_U10 (.A1( u2_u8_u0_n131 ) , .ZN( u2_u8_u0_n141 ) , .A2( u2_u8_u0_n150 ) );
  AND3_X1 u2_u8_u0_U11 (.A2( u2_u8_u0_n112 ) , .ZN( u2_u8_u0_n127 ) , .A3( u2_u8_u0_n130 ) , .A1( u2_u8_u0_n148 ) );
  AND2_X1 u2_u8_u0_U12 (.ZN( u2_u8_u0_n107 ) , .A1( u2_u8_u0_n130 ) , .A2( u2_u8_u0_n140 ) );
  AND2_X1 u2_u8_u0_U13 (.A2( u2_u8_u0_n129 ) , .A1( u2_u8_u0_n130 ) , .ZN( u2_u8_u0_n151 ) );
  AND2_X1 u2_u8_u0_U14 (.A1( u2_u8_u0_n108 ) , .A2( u2_u8_u0_n125 ) , .ZN( u2_u8_u0_n145 ) );
  INV_X1 u2_u8_u0_U15 (.A( u2_u8_u0_n143 ) , .ZN( u2_u8_u0_n173 ) );
  NOR2_X1 u2_u8_u0_U16 (.A2( u2_u8_u0_n136 ) , .ZN( u2_u8_u0_n147 ) , .A1( u2_u8_u0_n160 ) );
  AOI21_X1 u2_u8_u0_U17 (.B1( u2_u8_u0_n103 ) , .ZN( u2_u8_u0_n132 ) , .A( u2_u8_u0_n165 ) , .B2( u2_u8_u0_n93 ) );
  OAI22_X1 u2_u8_u0_U18 (.B1( u2_u8_u0_n131 ) , .A1( u2_u8_u0_n144 ) , .B2( u2_u8_u0_n147 ) , .A2( u2_u8_u0_n90 ) , .ZN( u2_u8_u0_n91 ) );
  AND3_X1 u2_u8_u0_U19 (.A3( u2_u8_u0_n121 ) , .A2( u2_u8_u0_n125 ) , .A1( u2_u8_u0_n148 ) , .ZN( u2_u8_u0_n90 ) );
  OAI22_X1 u2_u8_u0_U20 (.B1( u2_u8_u0_n125 ) , .ZN( u2_u8_u0_n126 ) , .A1( u2_u8_u0_n138 ) , .A2( u2_u8_u0_n146 ) , .B2( u2_u8_u0_n147 ) );
  NOR2_X1 u2_u8_u0_U21 (.A1( u2_u8_u0_n163 ) , .A2( u2_u8_u0_n164 ) , .ZN( u2_u8_u0_n95 ) );
  AOI22_X1 u2_u8_u0_U22 (.B2( u2_u8_u0_n109 ) , .A2( u2_u8_u0_n110 ) , .ZN( u2_u8_u0_n111 ) , .B1( u2_u8_u0_n118 ) , .A1( u2_u8_u0_n160 ) );
  NAND2_X1 u2_u8_u0_U23 (.A2( u2_u8_u0_n102 ) , .A1( u2_u8_u0_n103 ) , .ZN( u2_u8_u0_n149 ) );
  INV_X1 u2_u8_u0_U24 (.A( u2_u8_u0_n136 ) , .ZN( u2_u8_u0_n161 ) );
  INV_X1 u2_u8_u0_U25 (.A( u2_u8_u0_n118 ) , .ZN( u2_u8_u0_n158 ) );
  NAND2_X1 u2_u8_u0_U26 (.A2( u2_u8_u0_n100 ) , .ZN( u2_u8_u0_n131 ) , .A1( u2_u8_u0_n92 ) );
  NAND2_X1 u2_u8_u0_U27 (.ZN( u2_u8_u0_n108 ) , .A1( u2_u8_u0_n92 ) , .A2( u2_u8_u0_n94 ) );
  AOI21_X1 u2_u8_u0_U28 (.ZN( u2_u8_u0_n104 ) , .B1( u2_u8_u0_n107 ) , .B2( u2_u8_u0_n141 ) , .A( u2_u8_u0_n144 ) );
  AOI21_X1 u2_u8_u0_U29 (.B1( u2_u8_u0_n127 ) , .B2( u2_u8_u0_n129 ) , .A( u2_u8_u0_n138 ) , .ZN( u2_u8_u0_n96 ) );
  INV_X1 u2_u8_u0_U3 (.A( u2_u8_u0_n113 ) , .ZN( u2_u8_u0_n166 ) );
  NAND2_X1 u2_u8_u0_U30 (.A2( u2_u8_u0_n102 ) , .ZN( u2_u8_u0_n114 ) , .A1( u2_u8_u0_n92 ) );
  NOR2_X1 u2_u8_u0_U31 (.A1( u2_u8_u0_n120 ) , .ZN( u2_u8_u0_n143 ) , .A2( u2_u8_u0_n167 ) );
  OAI221_X1 u2_u8_u0_U32 (.C1( u2_u8_u0_n112 ) , .ZN( u2_u8_u0_n120 ) , .B1( u2_u8_u0_n138 ) , .B2( u2_u8_u0_n141 ) , .C2( u2_u8_u0_n147 ) , .A( u2_u8_u0_n172 ) );
  AOI211_X1 u2_u8_u0_U33 (.B( u2_u8_u0_n115 ) , .A( u2_u8_u0_n116 ) , .C2( u2_u8_u0_n117 ) , .C1( u2_u8_u0_n118 ) , .ZN( u2_u8_u0_n119 ) );
  NAND2_X1 u2_u8_u0_U34 (.A2( u2_u8_u0_n103 ) , .ZN( u2_u8_u0_n140 ) , .A1( u2_u8_u0_n94 ) );
  NAND2_X1 u2_u8_u0_U35 (.A1( u2_u8_u0_n100 ) , .A2( u2_u8_u0_n103 ) , .ZN( u2_u8_u0_n125 ) );
  NAND2_X1 u2_u8_u0_U36 (.A1( u2_u8_u0_n101 ) , .A2( u2_u8_u0_n102 ) , .ZN( u2_u8_u0_n150 ) );
  INV_X1 u2_u8_u0_U37 (.A( u2_u8_u0_n138 ) , .ZN( u2_u8_u0_n160 ) );
  NAND2_X1 u2_u8_u0_U38 (.A2( u2_u8_u0_n100 ) , .A1( u2_u8_u0_n101 ) , .ZN( u2_u8_u0_n139 ) );
  NAND2_X1 u2_u8_u0_U39 (.ZN( u2_u8_u0_n112 ) , .A2( u2_u8_u0_n92 ) , .A1( u2_u8_u0_n93 ) );
  AOI21_X1 u2_u8_u0_U4 (.B1( u2_u8_u0_n114 ) , .ZN( u2_u8_u0_n115 ) , .B2( u2_u8_u0_n129 ) , .A( u2_u8_u0_n161 ) );
  NAND2_X1 u2_u8_u0_U40 (.A1( u2_u8_u0_n101 ) , .ZN( u2_u8_u0_n130 ) , .A2( u2_u8_u0_n94 ) );
  INV_X1 u2_u8_u0_U41 (.ZN( u2_u8_u0_n172 ) , .A( u2_u8_u0_n88 ) );
  OAI222_X1 u2_u8_u0_U42 (.C1( u2_u8_u0_n108 ) , .A1( u2_u8_u0_n125 ) , .B2( u2_u8_u0_n128 ) , .B1( u2_u8_u0_n144 ) , .A2( u2_u8_u0_n158 ) , .C2( u2_u8_u0_n161 ) , .ZN( u2_u8_u0_n88 ) );
  NAND2_X1 u2_u8_u0_U43 (.A2( u2_u8_u0_n101 ) , .ZN( u2_u8_u0_n121 ) , .A1( u2_u8_u0_n93 ) );
  OR3_X1 u2_u8_u0_U44 (.A3( u2_u8_u0_n152 ) , .A2( u2_u8_u0_n153 ) , .A1( u2_u8_u0_n154 ) , .ZN( u2_u8_u0_n155 ) );
  AOI21_X1 u2_u8_u0_U45 (.A( u2_u8_u0_n144 ) , .B2( u2_u8_u0_n145 ) , .B1( u2_u8_u0_n146 ) , .ZN( u2_u8_u0_n154 ) );
  AOI21_X1 u2_u8_u0_U46 (.B2( u2_u8_u0_n150 ) , .B1( u2_u8_u0_n151 ) , .ZN( u2_u8_u0_n152 ) , .A( u2_u8_u0_n158 ) );
  AOI21_X1 u2_u8_u0_U47 (.A( u2_u8_u0_n147 ) , .B2( u2_u8_u0_n148 ) , .B1( u2_u8_u0_n149 ) , .ZN( u2_u8_u0_n153 ) );
  INV_X1 u2_u8_u0_U48 (.ZN( u2_u8_u0_n171 ) , .A( u2_u8_u0_n99 ) );
  OAI211_X1 u2_u8_u0_U49 (.C2( u2_u8_u0_n140 ) , .C1( u2_u8_u0_n161 ) , .A( u2_u8_u0_n169 ) , .B( u2_u8_u0_n98 ) , .ZN( u2_u8_u0_n99 ) );
  AOI21_X1 u2_u8_u0_U5 (.B2( u2_u8_u0_n131 ) , .ZN( u2_u8_u0_n134 ) , .B1( u2_u8_u0_n151 ) , .A( u2_u8_u0_n158 ) );
  INV_X1 u2_u8_u0_U50 (.ZN( u2_u8_u0_n169 ) , .A( u2_u8_u0_n91 ) );
  AOI211_X1 u2_u8_u0_U51 (.C1( u2_u8_u0_n118 ) , .A( u2_u8_u0_n123 ) , .B( u2_u8_u0_n96 ) , .C2( u2_u8_u0_n97 ) , .ZN( u2_u8_u0_n98 ) );
  NOR2_X1 u2_u8_u0_U52 (.A2( u2_u8_X_4 ) , .A1( u2_u8_X_5 ) , .ZN( u2_u8_u0_n118 ) );
  NOR2_X1 u2_u8_u0_U53 (.A2( u2_u8_X_1 ) , .ZN( u2_u8_u0_n101 ) , .A1( u2_u8_u0_n163 ) );
  NOR2_X1 u2_u8_u0_U54 (.A2( u2_u8_X_3 ) , .A1( u2_u8_X_6 ) , .ZN( u2_u8_u0_n94 ) );
  NOR2_X1 u2_u8_u0_U55 (.A2( u2_u8_X_6 ) , .ZN( u2_u8_u0_n100 ) , .A1( u2_u8_u0_n162 ) );
  NAND2_X1 u2_u8_u0_U56 (.A2( u2_u8_X_4 ) , .A1( u2_u8_X_5 ) , .ZN( u2_u8_u0_n144 ) );
  NOR2_X1 u2_u8_u0_U57 (.A2( u2_u8_X_5 ) , .ZN( u2_u8_u0_n136 ) , .A1( u2_u8_u0_n159 ) );
  NAND2_X1 u2_u8_u0_U58 (.A1( u2_u8_X_5 ) , .ZN( u2_u8_u0_n138 ) , .A2( u2_u8_u0_n159 ) );
  AND2_X1 u2_u8_u0_U59 (.A2( u2_u8_X_3 ) , .A1( u2_u8_X_6 ) , .ZN( u2_u8_u0_n102 ) );
  NOR2_X1 u2_u8_u0_U6 (.A1( u2_u8_u0_n108 ) , .ZN( u2_u8_u0_n123 ) , .A2( u2_u8_u0_n158 ) );
  AND2_X1 u2_u8_u0_U60 (.A1( u2_u8_X_6 ) , .A2( u2_u8_u0_n162 ) , .ZN( u2_u8_u0_n93 ) );
  INV_X1 u2_u8_u0_U61 (.A( u2_u8_X_4 ) , .ZN( u2_u8_u0_n159 ) );
  INV_X1 u2_u8_u0_U62 (.A( u2_u8_X_1 ) , .ZN( u2_u8_u0_n164 ) );
  INV_X1 u2_u8_u0_U63 (.A( u2_u8_X_3 ) , .ZN( u2_u8_u0_n162 ) );
  INV_X1 u2_u8_u0_U64 (.A( u2_u8_u0_n126 ) , .ZN( u2_u8_u0_n168 ) );
  AOI211_X1 u2_u8_u0_U65 (.B( u2_u8_u0_n133 ) , .A( u2_u8_u0_n134 ) , .C2( u2_u8_u0_n135 ) , .C1( u2_u8_u0_n136 ) , .ZN( u2_u8_u0_n137 ) );
  OR4_X1 u2_u8_u0_U66 (.ZN( u2_out8_17 ) , .A4( u2_u8_u0_n122 ) , .A2( u2_u8_u0_n123 ) , .A1( u2_u8_u0_n124 ) , .A3( u2_u8_u0_n170 ) );
  AOI21_X1 u2_u8_u0_U67 (.B2( u2_u8_u0_n107 ) , .ZN( u2_u8_u0_n124 ) , .B1( u2_u8_u0_n128 ) , .A( u2_u8_u0_n161 ) );
  INV_X1 u2_u8_u0_U68 (.A( u2_u8_u0_n111 ) , .ZN( u2_u8_u0_n170 ) );
  OR4_X1 u2_u8_u0_U69 (.ZN( u2_out8_31 ) , .A4( u2_u8_u0_n155 ) , .A2( u2_u8_u0_n156 ) , .A1( u2_u8_u0_n157 ) , .A3( u2_u8_u0_n173 ) );
  OAI21_X1 u2_u8_u0_U7 (.B1( u2_u8_u0_n150 ) , .B2( u2_u8_u0_n158 ) , .A( u2_u8_u0_n172 ) , .ZN( u2_u8_u0_n89 ) );
  AOI21_X1 u2_u8_u0_U70 (.A( u2_u8_u0_n138 ) , .B2( u2_u8_u0_n139 ) , .B1( u2_u8_u0_n140 ) , .ZN( u2_u8_u0_n157 ) );
  AOI211_X1 u2_u8_u0_U71 (.B( u2_u8_u0_n104 ) , .A( u2_u8_u0_n105 ) , .ZN( u2_u8_u0_n106 ) , .C2( u2_u8_u0_n113 ) , .C1( u2_u8_u0_n160 ) );
  INV_X1 u2_u8_u0_U72 (.ZN( u2_u8_u0_n174 ) , .A( u2_u8_u0_n89 ) );
  INV_X1 u2_u8_u0_U73 (.A( u2_u8_u0_n142 ) , .ZN( u2_u8_u0_n165 ) );
  AOI21_X1 u2_u8_u0_U74 (.ZN( u2_u8_u0_n116 ) , .B2( u2_u8_u0_n142 ) , .A( u2_u8_u0_n144 ) , .B1( u2_u8_u0_n166 ) );
  AOI21_X1 u2_u8_u0_U75 (.B2( u2_u8_u0_n141 ) , .B1( u2_u8_u0_n142 ) , .ZN( u2_u8_u0_n156 ) , .A( u2_u8_u0_n161 ) );
  OAI221_X1 u2_u8_u0_U76 (.C1( u2_u8_u0_n121 ) , .ZN( u2_u8_u0_n122 ) , .B2( u2_u8_u0_n127 ) , .A( u2_u8_u0_n143 ) , .B1( u2_u8_u0_n144 ) , .C2( u2_u8_u0_n147 ) );
  AOI21_X1 u2_u8_u0_U77 (.B1( u2_u8_u0_n132 ) , .ZN( u2_u8_u0_n133 ) , .A( u2_u8_u0_n144 ) , .B2( u2_u8_u0_n166 ) );
  OAI22_X1 u2_u8_u0_U78 (.ZN( u2_u8_u0_n105 ) , .A2( u2_u8_u0_n132 ) , .B1( u2_u8_u0_n146 ) , .A1( u2_u8_u0_n147 ) , .B2( u2_u8_u0_n161 ) );
  NAND2_X1 u2_u8_u0_U79 (.ZN( u2_u8_u0_n110 ) , .A2( u2_u8_u0_n132 ) , .A1( u2_u8_u0_n145 ) );
  AND2_X1 u2_u8_u0_U8 (.A1( u2_u8_u0_n114 ) , .A2( u2_u8_u0_n121 ) , .ZN( u2_u8_u0_n146 ) );
  INV_X1 u2_u8_u0_U80 (.A( u2_u8_u0_n119 ) , .ZN( u2_u8_u0_n167 ) );
  NAND2_X1 u2_u8_u0_U81 (.ZN( u2_u8_u0_n148 ) , .A1( u2_u8_u0_n93 ) , .A2( u2_u8_u0_n95 ) );
  NAND2_X1 u2_u8_u0_U82 (.A1( u2_u8_u0_n100 ) , .ZN( u2_u8_u0_n129 ) , .A2( u2_u8_u0_n95 ) );
  NAND2_X1 u2_u8_u0_U83 (.A1( u2_u8_u0_n102 ) , .ZN( u2_u8_u0_n128 ) , .A2( u2_u8_u0_n95 ) );
  NOR2_X1 u2_u8_u0_U84 (.A2( u2_u8_X_1 ) , .A1( u2_u8_X_2 ) , .ZN( u2_u8_u0_n92 ) );
  NAND2_X1 u2_u8_u0_U85 (.ZN( u2_u8_u0_n142 ) , .A1( u2_u8_u0_n94 ) , .A2( u2_u8_u0_n95 ) );
  NOR2_X1 u2_u8_u0_U86 (.A2( u2_u8_X_2 ) , .ZN( u2_u8_u0_n103 ) , .A1( u2_u8_u0_n164 ) );
  INV_X1 u2_u8_u0_U87 (.A( u2_u8_X_2 ) , .ZN( u2_u8_u0_n163 ) );
  NAND3_X1 u2_u8_u0_U88 (.ZN( u2_out8_23 ) , .A3( u2_u8_u0_n137 ) , .A1( u2_u8_u0_n168 ) , .A2( u2_u8_u0_n171 ) );
  NAND3_X1 u2_u8_u0_U89 (.A3( u2_u8_u0_n127 ) , .A2( u2_u8_u0_n128 ) , .ZN( u2_u8_u0_n135 ) , .A1( u2_u8_u0_n150 ) );
  NAND2_X1 u2_u8_u0_U9 (.ZN( u2_u8_u0_n113 ) , .A1( u2_u8_u0_n139 ) , .A2( u2_u8_u0_n149 ) );
  NAND3_X1 u2_u8_u0_U90 (.ZN( u2_u8_u0_n117 ) , .A3( u2_u8_u0_n132 ) , .A2( u2_u8_u0_n139 ) , .A1( u2_u8_u0_n148 ) );
  NAND3_X1 u2_u8_u0_U91 (.ZN( u2_u8_u0_n109 ) , .A2( u2_u8_u0_n114 ) , .A3( u2_u8_u0_n140 ) , .A1( u2_u8_u0_n149 ) );
  NAND3_X1 u2_u8_u0_U92 (.ZN( u2_out8_9 ) , .A3( u2_u8_u0_n106 ) , .A2( u2_u8_u0_n171 ) , .A1( u2_u8_u0_n174 ) );
  NAND3_X1 u2_u8_u0_U93 (.A2( u2_u8_u0_n128 ) , .A1( u2_u8_u0_n132 ) , .A3( u2_u8_u0_n146 ) , .ZN( u2_u8_u0_n97 ) );
  AOI21_X1 u2_u8_u1_U10 (.B2( u2_u8_u1_n155 ) , .B1( u2_u8_u1_n156 ) , .ZN( u2_u8_u1_n157 ) , .A( u2_u8_u1_n174 ) );
  NAND3_X1 u2_u8_u1_U100 (.ZN( u2_u8_u1_n113 ) , .A1( u2_u8_u1_n120 ) , .A3( u2_u8_u1_n133 ) , .A2( u2_u8_u1_n155 ) );
  NAND2_X1 u2_u8_u1_U11 (.ZN( u2_u8_u1_n140 ) , .A2( u2_u8_u1_n150 ) , .A1( u2_u8_u1_n155 ) );
  NAND2_X1 u2_u8_u1_U12 (.A1( u2_u8_u1_n131 ) , .ZN( u2_u8_u1_n147 ) , .A2( u2_u8_u1_n153 ) );
  AOI22_X1 u2_u8_u1_U13 (.B2( u2_u8_u1_n136 ) , .A2( u2_u8_u1_n137 ) , .ZN( u2_u8_u1_n143 ) , .A1( u2_u8_u1_n171 ) , .B1( u2_u8_u1_n173 ) );
  INV_X1 u2_u8_u1_U14 (.A( u2_u8_u1_n147 ) , .ZN( u2_u8_u1_n181 ) );
  INV_X1 u2_u8_u1_U15 (.A( u2_u8_u1_n139 ) , .ZN( u2_u8_u1_n174 ) );
  OR4_X1 u2_u8_u1_U16 (.A4( u2_u8_u1_n106 ) , .A3( u2_u8_u1_n107 ) , .ZN( u2_u8_u1_n108 ) , .A1( u2_u8_u1_n117 ) , .A2( u2_u8_u1_n184 ) );
  AOI21_X1 u2_u8_u1_U17 (.ZN( u2_u8_u1_n106 ) , .A( u2_u8_u1_n112 ) , .B1( u2_u8_u1_n154 ) , .B2( u2_u8_u1_n156 ) );
  AOI21_X1 u2_u8_u1_U18 (.ZN( u2_u8_u1_n107 ) , .B1( u2_u8_u1_n134 ) , .B2( u2_u8_u1_n149 ) , .A( u2_u8_u1_n174 ) );
  INV_X1 u2_u8_u1_U19 (.A( u2_u8_u1_n101 ) , .ZN( u2_u8_u1_n184 ) );
  INV_X1 u2_u8_u1_U20 (.A( u2_u8_u1_n112 ) , .ZN( u2_u8_u1_n171 ) );
  NAND2_X1 u2_u8_u1_U21 (.ZN( u2_u8_u1_n141 ) , .A1( u2_u8_u1_n153 ) , .A2( u2_u8_u1_n156 ) );
  AND2_X1 u2_u8_u1_U22 (.A1( u2_u8_u1_n123 ) , .ZN( u2_u8_u1_n134 ) , .A2( u2_u8_u1_n161 ) );
  NAND2_X1 u2_u8_u1_U23 (.A2( u2_u8_u1_n115 ) , .A1( u2_u8_u1_n116 ) , .ZN( u2_u8_u1_n148 ) );
  NAND2_X1 u2_u8_u1_U24 (.A2( u2_u8_u1_n133 ) , .A1( u2_u8_u1_n135 ) , .ZN( u2_u8_u1_n159 ) );
  NAND2_X1 u2_u8_u1_U25 (.A2( u2_u8_u1_n115 ) , .A1( u2_u8_u1_n120 ) , .ZN( u2_u8_u1_n132 ) );
  INV_X1 u2_u8_u1_U26 (.A( u2_u8_u1_n154 ) , .ZN( u2_u8_u1_n178 ) );
  INV_X1 u2_u8_u1_U27 (.A( u2_u8_u1_n151 ) , .ZN( u2_u8_u1_n183 ) );
  AND2_X1 u2_u8_u1_U28 (.A1( u2_u8_u1_n129 ) , .A2( u2_u8_u1_n133 ) , .ZN( u2_u8_u1_n149 ) );
  INV_X1 u2_u8_u1_U29 (.A( u2_u8_u1_n131 ) , .ZN( u2_u8_u1_n180 ) );
  INV_X1 u2_u8_u1_U3 (.A( u2_u8_u1_n159 ) , .ZN( u2_u8_u1_n182 ) );
  AOI221_X1 u2_u8_u1_U30 (.B1( u2_u8_u1_n140 ) , .ZN( u2_u8_u1_n167 ) , .B2( u2_u8_u1_n172 ) , .C2( u2_u8_u1_n175 ) , .C1( u2_u8_u1_n178 ) , .A( u2_u8_u1_n188 ) );
  INV_X1 u2_u8_u1_U31 (.ZN( u2_u8_u1_n188 ) , .A( u2_u8_u1_n97 ) );
  AOI211_X1 u2_u8_u1_U32 (.A( u2_u8_u1_n118 ) , .C1( u2_u8_u1_n132 ) , .C2( u2_u8_u1_n139 ) , .B( u2_u8_u1_n96 ) , .ZN( u2_u8_u1_n97 ) );
  AOI21_X1 u2_u8_u1_U33 (.B2( u2_u8_u1_n121 ) , .B1( u2_u8_u1_n135 ) , .A( u2_u8_u1_n152 ) , .ZN( u2_u8_u1_n96 ) );
  OAI221_X1 u2_u8_u1_U34 (.A( u2_u8_u1_n119 ) , .C2( u2_u8_u1_n129 ) , .ZN( u2_u8_u1_n138 ) , .B2( u2_u8_u1_n152 ) , .C1( u2_u8_u1_n174 ) , .B1( u2_u8_u1_n187 ) );
  INV_X1 u2_u8_u1_U35 (.A( u2_u8_u1_n148 ) , .ZN( u2_u8_u1_n187 ) );
  AOI211_X1 u2_u8_u1_U36 (.B( u2_u8_u1_n117 ) , .A( u2_u8_u1_n118 ) , .ZN( u2_u8_u1_n119 ) , .C2( u2_u8_u1_n146 ) , .C1( u2_u8_u1_n159 ) );
  NOR2_X1 u2_u8_u1_U37 (.A1( u2_u8_u1_n168 ) , .A2( u2_u8_u1_n176 ) , .ZN( u2_u8_u1_n98 ) );
  AOI211_X1 u2_u8_u1_U38 (.B( u2_u8_u1_n162 ) , .A( u2_u8_u1_n163 ) , .C2( u2_u8_u1_n164 ) , .ZN( u2_u8_u1_n165 ) , .C1( u2_u8_u1_n171 ) );
  AOI21_X1 u2_u8_u1_U39 (.A( u2_u8_u1_n160 ) , .B2( u2_u8_u1_n161 ) , .ZN( u2_u8_u1_n162 ) , .B1( u2_u8_u1_n182 ) );
  AOI221_X1 u2_u8_u1_U4 (.A( u2_u8_u1_n138 ) , .C2( u2_u8_u1_n139 ) , .C1( u2_u8_u1_n140 ) , .B2( u2_u8_u1_n141 ) , .ZN( u2_u8_u1_n142 ) , .B1( u2_u8_u1_n175 ) );
  OR2_X1 u2_u8_u1_U40 (.A2( u2_u8_u1_n157 ) , .A1( u2_u8_u1_n158 ) , .ZN( u2_u8_u1_n163 ) );
  NAND2_X1 u2_u8_u1_U41 (.A1( u2_u8_u1_n128 ) , .ZN( u2_u8_u1_n146 ) , .A2( u2_u8_u1_n160 ) );
  NAND2_X1 u2_u8_u1_U42 (.A2( u2_u8_u1_n112 ) , .ZN( u2_u8_u1_n139 ) , .A1( u2_u8_u1_n152 ) );
  NAND2_X1 u2_u8_u1_U43 (.A1( u2_u8_u1_n105 ) , .ZN( u2_u8_u1_n156 ) , .A2( u2_u8_u1_n99 ) );
  NOR2_X1 u2_u8_u1_U44 (.ZN( u2_u8_u1_n117 ) , .A1( u2_u8_u1_n121 ) , .A2( u2_u8_u1_n160 ) );
  OAI21_X1 u2_u8_u1_U45 (.B2( u2_u8_u1_n123 ) , .ZN( u2_u8_u1_n145 ) , .B1( u2_u8_u1_n160 ) , .A( u2_u8_u1_n185 ) );
  INV_X1 u2_u8_u1_U46 (.A( u2_u8_u1_n122 ) , .ZN( u2_u8_u1_n185 ) );
  AOI21_X1 u2_u8_u1_U47 (.B2( u2_u8_u1_n120 ) , .B1( u2_u8_u1_n121 ) , .ZN( u2_u8_u1_n122 ) , .A( u2_u8_u1_n128 ) );
  AOI21_X1 u2_u8_u1_U48 (.A( u2_u8_u1_n128 ) , .B2( u2_u8_u1_n129 ) , .ZN( u2_u8_u1_n130 ) , .B1( u2_u8_u1_n150 ) );
  NAND2_X1 u2_u8_u1_U49 (.ZN( u2_u8_u1_n112 ) , .A1( u2_u8_u1_n169 ) , .A2( u2_u8_u1_n170 ) );
  AOI211_X1 u2_u8_u1_U5 (.ZN( u2_u8_u1_n124 ) , .A( u2_u8_u1_n138 ) , .C2( u2_u8_u1_n139 ) , .B( u2_u8_u1_n145 ) , .C1( u2_u8_u1_n147 ) );
  NAND2_X1 u2_u8_u1_U50 (.ZN( u2_u8_u1_n129 ) , .A2( u2_u8_u1_n95 ) , .A1( u2_u8_u1_n98 ) );
  NAND2_X1 u2_u8_u1_U51 (.A1( u2_u8_u1_n102 ) , .ZN( u2_u8_u1_n154 ) , .A2( u2_u8_u1_n99 ) );
  NAND2_X1 u2_u8_u1_U52 (.A2( u2_u8_u1_n100 ) , .ZN( u2_u8_u1_n135 ) , .A1( u2_u8_u1_n99 ) );
  AOI21_X1 u2_u8_u1_U53 (.A( u2_u8_u1_n152 ) , .B2( u2_u8_u1_n153 ) , .B1( u2_u8_u1_n154 ) , .ZN( u2_u8_u1_n158 ) );
  INV_X1 u2_u8_u1_U54 (.A( u2_u8_u1_n160 ) , .ZN( u2_u8_u1_n175 ) );
  NAND2_X1 u2_u8_u1_U55 (.A1( u2_u8_u1_n100 ) , .ZN( u2_u8_u1_n116 ) , .A2( u2_u8_u1_n95 ) );
  NAND2_X1 u2_u8_u1_U56 (.A1( u2_u8_u1_n102 ) , .ZN( u2_u8_u1_n131 ) , .A2( u2_u8_u1_n95 ) );
  NAND2_X1 u2_u8_u1_U57 (.A2( u2_u8_u1_n104 ) , .ZN( u2_u8_u1_n121 ) , .A1( u2_u8_u1_n98 ) );
  NAND2_X1 u2_u8_u1_U58 (.A1( u2_u8_u1_n103 ) , .ZN( u2_u8_u1_n153 ) , .A2( u2_u8_u1_n98 ) );
  NAND2_X1 u2_u8_u1_U59 (.A2( u2_u8_u1_n104 ) , .A1( u2_u8_u1_n105 ) , .ZN( u2_u8_u1_n133 ) );
  AOI22_X1 u2_u8_u1_U6 (.B2( u2_u8_u1_n113 ) , .A2( u2_u8_u1_n114 ) , .ZN( u2_u8_u1_n125 ) , .A1( u2_u8_u1_n171 ) , .B1( u2_u8_u1_n173 ) );
  NAND2_X1 u2_u8_u1_U60 (.ZN( u2_u8_u1_n150 ) , .A2( u2_u8_u1_n98 ) , .A1( u2_u8_u1_n99 ) );
  NAND2_X1 u2_u8_u1_U61 (.A1( u2_u8_u1_n105 ) , .ZN( u2_u8_u1_n155 ) , .A2( u2_u8_u1_n95 ) );
  OAI21_X1 u2_u8_u1_U62 (.ZN( u2_u8_u1_n109 ) , .B1( u2_u8_u1_n129 ) , .B2( u2_u8_u1_n160 ) , .A( u2_u8_u1_n167 ) );
  NAND2_X1 u2_u8_u1_U63 (.A2( u2_u8_u1_n100 ) , .A1( u2_u8_u1_n103 ) , .ZN( u2_u8_u1_n120 ) );
  NAND2_X1 u2_u8_u1_U64 (.A1( u2_u8_u1_n102 ) , .A2( u2_u8_u1_n104 ) , .ZN( u2_u8_u1_n115 ) );
  NAND2_X1 u2_u8_u1_U65 (.A2( u2_u8_u1_n100 ) , .A1( u2_u8_u1_n104 ) , .ZN( u2_u8_u1_n151 ) );
  NAND2_X1 u2_u8_u1_U66 (.A2( u2_u8_u1_n103 ) , .A1( u2_u8_u1_n105 ) , .ZN( u2_u8_u1_n161 ) );
  INV_X1 u2_u8_u1_U67 (.A( u2_u8_u1_n152 ) , .ZN( u2_u8_u1_n173 ) );
  INV_X1 u2_u8_u1_U68 (.A( u2_u8_u1_n128 ) , .ZN( u2_u8_u1_n172 ) );
  NAND2_X1 u2_u8_u1_U69 (.A2( u2_u8_u1_n102 ) , .A1( u2_u8_u1_n103 ) , .ZN( u2_u8_u1_n123 ) );
  NAND2_X1 u2_u8_u1_U7 (.ZN( u2_u8_u1_n114 ) , .A1( u2_u8_u1_n134 ) , .A2( u2_u8_u1_n156 ) );
  NOR2_X1 u2_u8_u1_U70 (.A2( u2_u8_X_7 ) , .A1( u2_u8_X_8 ) , .ZN( u2_u8_u1_n95 ) );
  NOR2_X1 u2_u8_u1_U71 (.A1( u2_u8_X_12 ) , .A2( u2_u8_X_9 ) , .ZN( u2_u8_u1_n100 ) );
  NOR2_X1 u2_u8_u1_U72 (.A2( u2_u8_X_8 ) , .A1( u2_u8_u1_n177 ) , .ZN( u2_u8_u1_n99 ) );
  NOR2_X1 u2_u8_u1_U73 (.A2( u2_u8_X_12 ) , .ZN( u2_u8_u1_n102 ) , .A1( u2_u8_u1_n176 ) );
  NOR2_X1 u2_u8_u1_U74 (.A2( u2_u8_X_9 ) , .ZN( u2_u8_u1_n105 ) , .A1( u2_u8_u1_n168 ) );
  NAND2_X1 u2_u8_u1_U75 (.A1( u2_u8_X_10 ) , .ZN( u2_u8_u1_n160 ) , .A2( u2_u8_u1_n169 ) );
  NAND2_X1 u2_u8_u1_U76 (.A2( u2_u8_X_10 ) , .A1( u2_u8_X_11 ) , .ZN( u2_u8_u1_n152 ) );
  NAND2_X1 u2_u8_u1_U77 (.A1( u2_u8_X_11 ) , .ZN( u2_u8_u1_n128 ) , .A2( u2_u8_u1_n170 ) );
  AND2_X1 u2_u8_u1_U78 (.A2( u2_u8_X_7 ) , .A1( u2_u8_X_8 ) , .ZN( u2_u8_u1_n104 ) );
  AND2_X1 u2_u8_u1_U79 (.A1( u2_u8_X_8 ) , .ZN( u2_u8_u1_n103 ) , .A2( u2_u8_u1_n177 ) );
  NOR2_X1 u2_u8_u1_U8 (.A1( u2_u8_u1_n112 ) , .A2( u2_u8_u1_n116 ) , .ZN( u2_u8_u1_n118 ) );
  INV_X1 u2_u8_u1_U80 (.A( u2_u8_X_10 ) , .ZN( u2_u8_u1_n170 ) );
  INV_X1 u2_u8_u1_U81 (.A( u2_u8_X_9 ) , .ZN( u2_u8_u1_n176 ) );
  INV_X1 u2_u8_u1_U82 (.A( u2_u8_X_11 ) , .ZN( u2_u8_u1_n169 ) );
  INV_X1 u2_u8_u1_U83 (.A( u2_u8_X_12 ) , .ZN( u2_u8_u1_n168 ) );
  INV_X1 u2_u8_u1_U84 (.A( u2_u8_X_7 ) , .ZN( u2_u8_u1_n177 ) );
  NAND4_X1 u2_u8_u1_U85 (.ZN( u2_out8_28 ) , .A4( u2_u8_u1_n124 ) , .A3( u2_u8_u1_n125 ) , .A2( u2_u8_u1_n126 ) , .A1( u2_u8_u1_n127 ) );
  OAI21_X1 u2_u8_u1_U86 (.ZN( u2_u8_u1_n127 ) , .B2( u2_u8_u1_n139 ) , .B1( u2_u8_u1_n175 ) , .A( u2_u8_u1_n183 ) );
  OAI21_X1 u2_u8_u1_U87 (.ZN( u2_u8_u1_n126 ) , .B2( u2_u8_u1_n140 ) , .A( u2_u8_u1_n146 ) , .B1( u2_u8_u1_n178 ) );
  NAND4_X1 u2_u8_u1_U88 (.ZN( u2_out8_18 ) , .A4( u2_u8_u1_n165 ) , .A3( u2_u8_u1_n166 ) , .A1( u2_u8_u1_n167 ) , .A2( u2_u8_u1_n186 ) );
  AOI22_X1 u2_u8_u1_U89 (.B2( u2_u8_u1_n146 ) , .B1( u2_u8_u1_n147 ) , .A2( u2_u8_u1_n148 ) , .ZN( u2_u8_u1_n166 ) , .A1( u2_u8_u1_n172 ) );
  OAI21_X1 u2_u8_u1_U9 (.ZN( u2_u8_u1_n101 ) , .B1( u2_u8_u1_n141 ) , .A( u2_u8_u1_n146 ) , .B2( u2_u8_u1_n183 ) );
  INV_X1 u2_u8_u1_U90 (.A( u2_u8_u1_n145 ) , .ZN( u2_u8_u1_n186 ) );
  NAND4_X1 u2_u8_u1_U91 (.ZN( u2_out8_2 ) , .A4( u2_u8_u1_n142 ) , .A3( u2_u8_u1_n143 ) , .A2( u2_u8_u1_n144 ) , .A1( u2_u8_u1_n179 ) );
  OAI21_X1 u2_u8_u1_U92 (.B2( u2_u8_u1_n132 ) , .ZN( u2_u8_u1_n144 ) , .A( u2_u8_u1_n146 ) , .B1( u2_u8_u1_n180 ) );
  INV_X1 u2_u8_u1_U93 (.A( u2_u8_u1_n130 ) , .ZN( u2_u8_u1_n179 ) );
  OR4_X1 u2_u8_u1_U94 (.ZN( u2_out8_13 ) , .A4( u2_u8_u1_n108 ) , .A3( u2_u8_u1_n109 ) , .A2( u2_u8_u1_n110 ) , .A1( u2_u8_u1_n111 ) );
  AOI21_X1 u2_u8_u1_U95 (.ZN( u2_u8_u1_n111 ) , .A( u2_u8_u1_n128 ) , .B2( u2_u8_u1_n131 ) , .B1( u2_u8_u1_n135 ) );
  AOI21_X1 u2_u8_u1_U96 (.ZN( u2_u8_u1_n110 ) , .A( u2_u8_u1_n116 ) , .B1( u2_u8_u1_n152 ) , .B2( u2_u8_u1_n160 ) );
  NAND3_X1 u2_u8_u1_U97 (.A3( u2_u8_u1_n149 ) , .A2( u2_u8_u1_n150 ) , .A1( u2_u8_u1_n151 ) , .ZN( u2_u8_u1_n164 ) );
  NAND3_X1 u2_u8_u1_U98 (.A3( u2_u8_u1_n134 ) , .A2( u2_u8_u1_n135 ) , .ZN( u2_u8_u1_n136 ) , .A1( u2_u8_u1_n151 ) );
  NAND3_X1 u2_u8_u1_U99 (.A1( u2_u8_u1_n133 ) , .ZN( u2_u8_u1_n137 ) , .A2( u2_u8_u1_n154 ) , .A3( u2_u8_u1_n181 ) );
  OAI22_X1 u2_u8_u2_U10 (.B1( u2_u8_u2_n151 ) , .A2( u2_u8_u2_n152 ) , .A1( u2_u8_u2_n153 ) , .ZN( u2_u8_u2_n160 ) , .B2( u2_u8_u2_n168 ) );
  NAND3_X1 u2_u8_u2_U100 (.A2( u2_u8_u2_n100 ) , .A1( u2_u8_u2_n104 ) , .A3( u2_u8_u2_n138 ) , .ZN( u2_u8_u2_n98 ) );
  NOR3_X1 u2_u8_u2_U11 (.A1( u2_u8_u2_n150 ) , .ZN( u2_u8_u2_n151 ) , .A3( u2_u8_u2_n175 ) , .A2( u2_u8_u2_n188 ) );
  AOI21_X1 u2_u8_u2_U12 (.B2( u2_u8_u2_n123 ) , .ZN( u2_u8_u2_n125 ) , .A( u2_u8_u2_n171 ) , .B1( u2_u8_u2_n184 ) );
  INV_X1 u2_u8_u2_U13 (.A( u2_u8_u2_n150 ) , .ZN( u2_u8_u2_n184 ) );
  AOI21_X1 u2_u8_u2_U14 (.ZN( u2_u8_u2_n144 ) , .B2( u2_u8_u2_n155 ) , .A( u2_u8_u2_n172 ) , .B1( u2_u8_u2_n185 ) );
  AOI21_X1 u2_u8_u2_U15 (.B2( u2_u8_u2_n143 ) , .ZN( u2_u8_u2_n145 ) , .B1( u2_u8_u2_n152 ) , .A( u2_u8_u2_n171 ) );
  INV_X1 u2_u8_u2_U16 (.A( u2_u8_u2_n156 ) , .ZN( u2_u8_u2_n171 ) );
  INV_X1 u2_u8_u2_U17 (.A( u2_u8_u2_n120 ) , .ZN( u2_u8_u2_n188 ) );
  NAND2_X1 u2_u8_u2_U18 (.A2( u2_u8_u2_n122 ) , .ZN( u2_u8_u2_n150 ) , .A1( u2_u8_u2_n152 ) );
  INV_X1 u2_u8_u2_U19 (.A( u2_u8_u2_n153 ) , .ZN( u2_u8_u2_n170 ) );
  INV_X1 u2_u8_u2_U20 (.A( u2_u8_u2_n137 ) , .ZN( u2_u8_u2_n173 ) );
  NAND2_X1 u2_u8_u2_U21 (.A1( u2_u8_u2_n132 ) , .A2( u2_u8_u2_n139 ) , .ZN( u2_u8_u2_n157 ) );
  INV_X1 u2_u8_u2_U22 (.A( u2_u8_u2_n113 ) , .ZN( u2_u8_u2_n178 ) );
  INV_X1 u2_u8_u2_U23 (.A( u2_u8_u2_n139 ) , .ZN( u2_u8_u2_n175 ) );
  INV_X1 u2_u8_u2_U24 (.A( u2_u8_u2_n155 ) , .ZN( u2_u8_u2_n181 ) );
  INV_X1 u2_u8_u2_U25 (.A( u2_u8_u2_n119 ) , .ZN( u2_u8_u2_n177 ) );
  INV_X1 u2_u8_u2_U26 (.A( u2_u8_u2_n116 ) , .ZN( u2_u8_u2_n180 ) );
  INV_X1 u2_u8_u2_U27 (.A( u2_u8_u2_n131 ) , .ZN( u2_u8_u2_n179 ) );
  INV_X1 u2_u8_u2_U28 (.A( u2_u8_u2_n154 ) , .ZN( u2_u8_u2_n176 ) );
  NAND2_X1 u2_u8_u2_U29 (.A2( u2_u8_u2_n116 ) , .A1( u2_u8_u2_n117 ) , .ZN( u2_u8_u2_n118 ) );
  NOR2_X1 u2_u8_u2_U3 (.ZN( u2_u8_u2_n121 ) , .A2( u2_u8_u2_n177 ) , .A1( u2_u8_u2_n180 ) );
  INV_X1 u2_u8_u2_U30 (.A( u2_u8_u2_n132 ) , .ZN( u2_u8_u2_n182 ) );
  INV_X1 u2_u8_u2_U31 (.A( u2_u8_u2_n158 ) , .ZN( u2_u8_u2_n183 ) );
  OAI21_X1 u2_u8_u2_U32 (.A( u2_u8_u2_n156 ) , .B1( u2_u8_u2_n157 ) , .ZN( u2_u8_u2_n158 ) , .B2( u2_u8_u2_n179 ) );
  NOR2_X1 u2_u8_u2_U33 (.ZN( u2_u8_u2_n156 ) , .A1( u2_u8_u2_n166 ) , .A2( u2_u8_u2_n169 ) );
  NOR2_X1 u2_u8_u2_U34 (.A2( u2_u8_u2_n114 ) , .ZN( u2_u8_u2_n137 ) , .A1( u2_u8_u2_n140 ) );
  NOR2_X1 u2_u8_u2_U35 (.A2( u2_u8_u2_n138 ) , .ZN( u2_u8_u2_n153 ) , .A1( u2_u8_u2_n156 ) );
  AOI211_X1 u2_u8_u2_U36 (.ZN( u2_u8_u2_n130 ) , .C1( u2_u8_u2_n138 ) , .C2( u2_u8_u2_n179 ) , .B( u2_u8_u2_n96 ) , .A( u2_u8_u2_n97 ) );
  OAI22_X1 u2_u8_u2_U37 (.B1( u2_u8_u2_n133 ) , .A2( u2_u8_u2_n137 ) , .A1( u2_u8_u2_n152 ) , .B2( u2_u8_u2_n168 ) , .ZN( u2_u8_u2_n97 ) );
  OAI221_X1 u2_u8_u2_U38 (.B1( u2_u8_u2_n113 ) , .C1( u2_u8_u2_n132 ) , .A( u2_u8_u2_n149 ) , .B2( u2_u8_u2_n171 ) , .C2( u2_u8_u2_n172 ) , .ZN( u2_u8_u2_n96 ) );
  OAI221_X1 u2_u8_u2_U39 (.A( u2_u8_u2_n115 ) , .C2( u2_u8_u2_n123 ) , .B2( u2_u8_u2_n143 ) , .B1( u2_u8_u2_n153 ) , .ZN( u2_u8_u2_n163 ) , .C1( u2_u8_u2_n168 ) );
  INV_X1 u2_u8_u2_U4 (.A( u2_u8_u2_n134 ) , .ZN( u2_u8_u2_n185 ) );
  OAI21_X1 u2_u8_u2_U40 (.A( u2_u8_u2_n114 ) , .ZN( u2_u8_u2_n115 ) , .B1( u2_u8_u2_n176 ) , .B2( u2_u8_u2_n178 ) );
  OAI221_X1 u2_u8_u2_U41 (.A( u2_u8_u2_n135 ) , .B2( u2_u8_u2_n136 ) , .B1( u2_u8_u2_n137 ) , .ZN( u2_u8_u2_n162 ) , .C2( u2_u8_u2_n167 ) , .C1( u2_u8_u2_n185 ) );
  AND3_X1 u2_u8_u2_U42 (.A3( u2_u8_u2_n131 ) , .A2( u2_u8_u2_n132 ) , .A1( u2_u8_u2_n133 ) , .ZN( u2_u8_u2_n136 ) );
  AOI22_X1 u2_u8_u2_U43 (.ZN( u2_u8_u2_n135 ) , .B1( u2_u8_u2_n140 ) , .A1( u2_u8_u2_n156 ) , .B2( u2_u8_u2_n180 ) , .A2( u2_u8_u2_n188 ) );
  AOI21_X1 u2_u8_u2_U44 (.ZN( u2_u8_u2_n149 ) , .B1( u2_u8_u2_n173 ) , .B2( u2_u8_u2_n188 ) , .A( u2_u8_u2_n95 ) );
  AND3_X1 u2_u8_u2_U45 (.A2( u2_u8_u2_n100 ) , .A1( u2_u8_u2_n104 ) , .A3( u2_u8_u2_n156 ) , .ZN( u2_u8_u2_n95 ) );
  OAI21_X1 u2_u8_u2_U46 (.A( u2_u8_u2_n141 ) , .B2( u2_u8_u2_n142 ) , .ZN( u2_u8_u2_n146 ) , .B1( u2_u8_u2_n153 ) );
  OAI21_X1 u2_u8_u2_U47 (.A( u2_u8_u2_n140 ) , .ZN( u2_u8_u2_n141 ) , .B1( u2_u8_u2_n176 ) , .B2( u2_u8_u2_n177 ) );
  NOR3_X1 u2_u8_u2_U48 (.ZN( u2_u8_u2_n142 ) , .A3( u2_u8_u2_n175 ) , .A2( u2_u8_u2_n178 ) , .A1( u2_u8_u2_n181 ) );
  OAI21_X1 u2_u8_u2_U49 (.A( u2_u8_u2_n101 ) , .B2( u2_u8_u2_n121 ) , .B1( u2_u8_u2_n153 ) , .ZN( u2_u8_u2_n164 ) );
  NOR4_X1 u2_u8_u2_U5 (.A4( u2_u8_u2_n124 ) , .A3( u2_u8_u2_n125 ) , .A2( u2_u8_u2_n126 ) , .A1( u2_u8_u2_n127 ) , .ZN( u2_u8_u2_n128 ) );
  NAND2_X1 u2_u8_u2_U50 (.A2( u2_u8_u2_n100 ) , .A1( u2_u8_u2_n107 ) , .ZN( u2_u8_u2_n155 ) );
  NAND2_X1 u2_u8_u2_U51 (.A2( u2_u8_u2_n105 ) , .A1( u2_u8_u2_n108 ) , .ZN( u2_u8_u2_n143 ) );
  NAND2_X1 u2_u8_u2_U52 (.A1( u2_u8_u2_n104 ) , .A2( u2_u8_u2_n106 ) , .ZN( u2_u8_u2_n152 ) );
  NAND2_X1 u2_u8_u2_U53 (.A1( u2_u8_u2_n100 ) , .A2( u2_u8_u2_n105 ) , .ZN( u2_u8_u2_n132 ) );
  INV_X1 u2_u8_u2_U54 (.A( u2_u8_u2_n140 ) , .ZN( u2_u8_u2_n168 ) );
  INV_X1 u2_u8_u2_U55 (.A( u2_u8_u2_n138 ) , .ZN( u2_u8_u2_n167 ) );
  NAND2_X1 u2_u8_u2_U56 (.A1( u2_u8_u2_n102 ) , .A2( u2_u8_u2_n106 ) , .ZN( u2_u8_u2_n113 ) );
  NAND2_X1 u2_u8_u2_U57 (.A1( u2_u8_u2_n106 ) , .A2( u2_u8_u2_n107 ) , .ZN( u2_u8_u2_n131 ) );
  NAND2_X1 u2_u8_u2_U58 (.A1( u2_u8_u2_n103 ) , .A2( u2_u8_u2_n107 ) , .ZN( u2_u8_u2_n139 ) );
  NAND2_X1 u2_u8_u2_U59 (.A1( u2_u8_u2_n103 ) , .A2( u2_u8_u2_n105 ) , .ZN( u2_u8_u2_n133 ) );
  AOI21_X1 u2_u8_u2_U6 (.B2( u2_u8_u2_n119 ) , .ZN( u2_u8_u2_n127 ) , .A( u2_u8_u2_n137 ) , .B1( u2_u8_u2_n155 ) );
  NAND2_X1 u2_u8_u2_U60 (.A1( u2_u8_u2_n102 ) , .A2( u2_u8_u2_n103 ) , .ZN( u2_u8_u2_n154 ) );
  NAND2_X1 u2_u8_u2_U61 (.A2( u2_u8_u2_n103 ) , .A1( u2_u8_u2_n104 ) , .ZN( u2_u8_u2_n119 ) );
  NAND2_X1 u2_u8_u2_U62 (.A2( u2_u8_u2_n107 ) , .A1( u2_u8_u2_n108 ) , .ZN( u2_u8_u2_n123 ) );
  NAND2_X1 u2_u8_u2_U63 (.A1( u2_u8_u2_n104 ) , .A2( u2_u8_u2_n108 ) , .ZN( u2_u8_u2_n122 ) );
  INV_X1 u2_u8_u2_U64 (.A( u2_u8_u2_n114 ) , .ZN( u2_u8_u2_n172 ) );
  NAND2_X1 u2_u8_u2_U65 (.A2( u2_u8_u2_n100 ) , .A1( u2_u8_u2_n102 ) , .ZN( u2_u8_u2_n116 ) );
  NAND2_X1 u2_u8_u2_U66 (.A1( u2_u8_u2_n102 ) , .A2( u2_u8_u2_n108 ) , .ZN( u2_u8_u2_n120 ) );
  NAND2_X1 u2_u8_u2_U67 (.A2( u2_u8_u2_n105 ) , .A1( u2_u8_u2_n106 ) , .ZN( u2_u8_u2_n117 ) );
  INV_X1 u2_u8_u2_U68 (.ZN( u2_u8_u2_n187 ) , .A( u2_u8_u2_n99 ) );
  OAI21_X1 u2_u8_u2_U69 (.B1( u2_u8_u2_n137 ) , .B2( u2_u8_u2_n143 ) , .A( u2_u8_u2_n98 ) , .ZN( u2_u8_u2_n99 ) );
  AOI21_X1 u2_u8_u2_U7 (.ZN( u2_u8_u2_n124 ) , .B1( u2_u8_u2_n131 ) , .B2( u2_u8_u2_n143 ) , .A( u2_u8_u2_n172 ) );
  NOR2_X1 u2_u8_u2_U70 (.A2( u2_u8_X_16 ) , .ZN( u2_u8_u2_n140 ) , .A1( u2_u8_u2_n166 ) );
  NOR2_X1 u2_u8_u2_U71 (.A2( u2_u8_X_13 ) , .A1( u2_u8_X_14 ) , .ZN( u2_u8_u2_n100 ) );
  NOR2_X1 u2_u8_u2_U72 (.A2( u2_u8_X_16 ) , .A1( u2_u8_X_17 ) , .ZN( u2_u8_u2_n138 ) );
  NOR2_X1 u2_u8_u2_U73 (.A2( u2_u8_X_15 ) , .A1( u2_u8_X_18 ) , .ZN( u2_u8_u2_n104 ) );
  NOR2_X1 u2_u8_u2_U74 (.A2( u2_u8_X_14 ) , .ZN( u2_u8_u2_n103 ) , .A1( u2_u8_u2_n174 ) );
  NOR2_X1 u2_u8_u2_U75 (.A2( u2_u8_X_15 ) , .ZN( u2_u8_u2_n102 ) , .A1( u2_u8_u2_n165 ) );
  NOR2_X1 u2_u8_u2_U76 (.A2( u2_u8_X_17 ) , .ZN( u2_u8_u2_n114 ) , .A1( u2_u8_u2_n169 ) );
  AND2_X1 u2_u8_u2_U77 (.A1( u2_u8_X_15 ) , .ZN( u2_u8_u2_n105 ) , .A2( u2_u8_u2_n165 ) );
  AND2_X1 u2_u8_u2_U78 (.A2( u2_u8_X_15 ) , .A1( u2_u8_X_18 ) , .ZN( u2_u8_u2_n107 ) );
  AND2_X1 u2_u8_u2_U79 (.A1( u2_u8_X_14 ) , .ZN( u2_u8_u2_n106 ) , .A2( u2_u8_u2_n174 ) );
  AOI21_X1 u2_u8_u2_U8 (.B2( u2_u8_u2_n120 ) , .B1( u2_u8_u2_n121 ) , .ZN( u2_u8_u2_n126 ) , .A( u2_u8_u2_n167 ) );
  AND2_X1 u2_u8_u2_U80 (.A1( u2_u8_X_13 ) , .A2( u2_u8_X_14 ) , .ZN( u2_u8_u2_n108 ) );
  INV_X1 u2_u8_u2_U81 (.A( u2_u8_X_16 ) , .ZN( u2_u8_u2_n169 ) );
  INV_X1 u2_u8_u2_U82 (.A( u2_u8_X_17 ) , .ZN( u2_u8_u2_n166 ) );
  INV_X1 u2_u8_u2_U83 (.A( u2_u8_X_13 ) , .ZN( u2_u8_u2_n174 ) );
  INV_X1 u2_u8_u2_U84 (.A( u2_u8_X_18 ) , .ZN( u2_u8_u2_n165 ) );
  NAND4_X1 u2_u8_u2_U85 (.ZN( u2_out8_30 ) , .A4( u2_u8_u2_n147 ) , .A3( u2_u8_u2_n148 ) , .A2( u2_u8_u2_n149 ) , .A1( u2_u8_u2_n187 ) );
  NOR3_X1 u2_u8_u2_U86 (.A3( u2_u8_u2_n144 ) , .A2( u2_u8_u2_n145 ) , .A1( u2_u8_u2_n146 ) , .ZN( u2_u8_u2_n147 ) );
  AOI21_X1 u2_u8_u2_U87 (.B2( u2_u8_u2_n138 ) , .ZN( u2_u8_u2_n148 ) , .A( u2_u8_u2_n162 ) , .B1( u2_u8_u2_n182 ) );
  NAND4_X1 u2_u8_u2_U88 (.ZN( u2_out8_24 ) , .A4( u2_u8_u2_n111 ) , .A3( u2_u8_u2_n112 ) , .A1( u2_u8_u2_n130 ) , .A2( u2_u8_u2_n187 ) );
  AOI221_X1 u2_u8_u2_U89 (.A( u2_u8_u2_n109 ) , .B1( u2_u8_u2_n110 ) , .ZN( u2_u8_u2_n111 ) , .C1( u2_u8_u2_n134 ) , .C2( u2_u8_u2_n170 ) , .B2( u2_u8_u2_n173 ) );
  OAI22_X1 u2_u8_u2_U9 (.ZN( u2_u8_u2_n109 ) , .A2( u2_u8_u2_n113 ) , .B2( u2_u8_u2_n133 ) , .B1( u2_u8_u2_n167 ) , .A1( u2_u8_u2_n168 ) );
  AOI21_X1 u2_u8_u2_U90 (.ZN( u2_u8_u2_n112 ) , .B2( u2_u8_u2_n156 ) , .A( u2_u8_u2_n164 ) , .B1( u2_u8_u2_n181 ) );
  NAND4_X1 u2_u8_u2_U91 (.ZN( u2_out8_16 ) , .A4( u2_u8_u2_n128 ) , .A3( u2_u8_u2_n129 ) , .A1( u2_u8_u2_n130 ) , .A2( u2_u8_u2_n186 ) );
  AOI22_X1 u2_u8_u2_U92 (.A2( u2_u8_u2_n118 ) , .ZN( u2_u8_u2_n129 ) , .A1( u2_u8_u2_n140 ) , .B1( u2_u8_u2_n157 ) , .B2( u2_u8_u2_n170 ) );
  INV_X1 u2_u8_u2_U93 (.A( u2_u8_u2_n163 ) , .ZN( u2_u8_u2_n186 ) );
  OR4_X1 u2_u8_u2_U94 (.ZN( u2_out8_6 ) , .A4( u2_u8_u2_n161 ) , .A3( u2_u8_u2_n162 ) , .A2( u2_u8_u2_n163 ) , .A1( u2_u8_u2_n164 ) );
  OR3_X1 u2_u8_u2_U95 (.A2( u2_u8_u2_n159 ) , .A1( u2_u8_u2_n160 ) , .ZN( u2_u8_u2_n161 ) , .A3( u2_u8_u2_n183 ) );
  AOI21_X1 u2_u8_u2_U96 (.B2( u2_u8_u2_n154 ) , .B1( u2_u8_u2_n155 ) , .ZN( u2_u8_u2_n159 ) , .A( u2_u8_u2_n167 ) );
  NAND3_X1 u2_u8_u2_U97 (.A2( u2_u8_u2_n117 ) , .A1( u2_u8_u2_n122 ) , .A3( u2_u8_u2_n123 ) , .ZN( u2_u8_u2_n134 ) );
  NAND3_X1 u2_u8_u2_U98 (.ZN( u2_u8_u2_n110 ) , .A2( u2_u8_u2_n131 ) , .A3( u2_u8_u2_n139 ) , .A1( u2_u8_u2_n154 ) );
  NAND3_X1 u2_u8_u2_U99 (.A2( u2_u8_u2_n100 ) , .ZN( u2_u8_u2_n101 ) , .A1( u2_u8_u2_n104 ) , .A3( u2_u8_u2_n114 ) );
  OAI22_X1 u2_u8_u3_U10 (.B1( u2_u8_u3_n113 ) , .A2( u2_u8_u3_n135 ) , .A1( u2_u8_u3_n150 ) , .B2( u2_u8_u3_n164 ) , .ZN( u2_u8_u3_n98 ) );
  OAI211_X1 u2_u8_u3_U11 (.B( u2_u8_u3_n106 ) , .ZN( u2_u8_u3_n119 ) , .C2( u2_u8_u3_n128 ) , .C1( u2_u8_u3_n167 ) , .A( u2_u8_u3_n181 ) );
  AOI221_X1 u2_u8_u3_U12 (.C1( u2_u8_u3_n105 ) , .ZN( u2_u8_u3_n106 ) , .A( u2_u8_u3_n131 ) , .B2( u2_u8_u3_n132 ) , .C2( u2_u8_u3_n133 ) , .B1( u2_u8_u3_n169 ) );
  INV_X1 u2_u8_u3_U13 (.ZN( u2_u8_u3_n181 ) , .A( u2_u8_u3_n98 ) );
  NAND2_X1 u2_u8_u3_U14 (.ZN( u2_u8_u3_n105 ) , .A2( u2_u8_u3_n130 ) , .A1( u2_u8_u3_n155 ) );
  AOI22_X1 u2_u8_u3_U15 (.B1( u2_u8_u3_n115 ) , .A2( u2_u8_u3_n116 ) , .ZN( u2_u8_u3_n123 ) , .B2( u2_u8_u3_n133 ) , .A1( u2_u8_u3_n169 ) );
  NAND2_X1 u2_u8_u3_U16 (.ZN( u2_u8_u3_n116 ) , .A2( u2_u8_u3_n151 ) , .A1( u2_u8_u3_n182 ) );
  NOR2_X1 u2_u8_u3_U17 (.ZN( u2_u8_u3_n126 ) , .A2( u2_u8_u3_n150 ) , .A1( u2_u8_u3_n164 ) );
  AOI21_X1 u2_u8_u3_U18 (.ZN( u2_u8_u3_n112 ) , .B2( u2_u8_u3_n146 ) , .B1( u2_u8_u3_n155 ) , .A( u2_u8_u3_n167 ) );
  NAND2_X1 u2_u8_u3_U19 (.A1( u2_u8_u3_n135 ) , .ZN( u2_u8_u3_n142 ) , .A2( u2_u8_u3_n164 ) );
  NAND2_X1 u2_u8_u3_U20 (.ZN( u2_u8_u3_n132 ) , .A2( u2_u8_u3_n152 ) , .A1( u2_u8_u3_n156 ) );
  AND2_X1 u2_u8_u3_U21 (.A2( u2_u8_u3_n113 ) , .A1( u2_u8_u3_n114 ) , .ZN( u2_u8_u3_n151 ) );
  INV_X1 u2_u8_u3_U22 (.A( u2_u8_u3_n133 ) , .ZN( u2_u8_u3_n165 ) );
  INV_X1 u2_u8_u3_U23 (.A( u2_u8_u3_n135 ) , .ZN( u2_u8_u3_n170 ) );
  NAND2_X1 u2_u8_u3_U24 (.A1( u2_u8_u3_n107 ) , .A2( u2_u8_u3_n108 ) , .ZN( u2_u8_u3_n140 ) );
  NAND2_X1 u2_u8_u3_U25 (.ZN( u2_u8_u3_n117 ) , .A1( u2_u8_u3_n124 ) , .A2( u2_u8_u3_n148 ) );
  NAND2_X1 u2_u8_u3_U26 (.ZN( u2_u8_u3_n143 ) , .A1( u2_u8_u3_n165 ) , .A2( u2_u8_u3_n167 ) );
  INV_X1 u2_u8_u3_U27 (.A( u2_u8_u3_n130 ) , .ZN( u2_u8_u3_n177 ) );
  INV_X1 u2_u8_u3_U28 (.A( u2_u8_u3_n128 ) , .ZN( u2_u8_u3_n176 ) );
  INV_X1 u2_u8_u3_U29 (.A( u2_u8_u3_n155 ) , .ZN( u2_u8_u3_n174 ) );
  INV_X1 u2_u8_u3_U3 (.A( u2_u8_u3_n129 ) , .ZN( u2_u8_u3_n183 ) );
  INV_X1 u2_u8_u3_U30 (.A( u2_u8_u3_n139 ) , .ZN( u2_u8_u3_n185 ) );
  NOR2_X1 u2_u8_u3_U31 (.ZN( u2_u8_u3_n135 ) , .A2( u2_u8_u3_n141 ) , .A1( u2_u8_u3_n169 ) );
  OAI222_X1 u2_u8_u3_U32 (.C2( u2_u8_u3_n107 ) , .A2( u2_u8_u3_n108 ) , .B1( u2_u8_u3_n135 ) , .ZN( u2_u8_u3_n138 ) , .B2( u2_u8_u3_n146 ) , .C1( u2_u8_u3_n154 ) , .A1( u2_u8_u3_n164 ) );
  NOR4_X1 u2_u8_u3_U33 (.A4( u2_u8_u3_n157 ) , .A3( u2_u8_u3_n158 ) , .A2( u2_u8_u3_n159 ) , .A1( u2_u8_u3_n160 ) , .ZN( u2_u8_u3_n161 ) );
  AOI21_X1 u2_u8_u3_U34 (.B2( u2_u8_u3_n152 ) , .B1( u2_u8_u3_n153 ) , .ZN( u2_u8_u3_n158 ) , .A( u2_u8_u3_n164 ) );
  AOI21_X1 u2_u8_u3_U35 (.A( u2_u8_u3_n149 ) , .B2( u2_u8_u3_n150 ) , .B1( u2_u8_u3_n151 ) , .ZN( u2_u8_u3_n159 ) );
  AOI21_X1 u2_u8_u3_U36 (.A( u2_u8_u3_n154 ) , .B2( u2_u8_u3_n155 ) , .B1( u2_u8_u3_n156 ) , .ZN( u2_u8_u3_n157 ) );
  AOI211_X1 u2_u8_u3_U37 (.ZN( u2_u8_u3_n109 ) , .A( u2_u8_u3_n119 ) , .C2( u2_u8_u3_n129 ) , .B( u2_u8_u3_n138 ) , .C1( u2_u8_u3_n141 ) );
  AOI211_X1 u2_u8_u3_U38 (.B( u2_u8_u3_n119 ) , .A( u2_u8_u3_n120 ) , .C2( u2_u8_u3_n121 ) , .ZN( u2_u8_u3_n122 ) , .C1( u2_u8_u3_n179 ) );
  INV_X1 u2_u8_u3_U39 (.A( u2_u8_u3_n156 ) , .ZN( u2_u8_u3_n179 ) );
  INV_X1 u2_u8_u3_U4 (.A( u2_u8_u3_n140 ) , .ZN( u2_u8_u3_n182 ) );
  OAI22_X1 u2_u8_u3_U40 (.B1( u2_u8_u3_n118 ) , .ZN( u2_u8_u3_n120 ) , .A1( u2_u8_u3_n135 ) , .B2( u2_u8_u3_n154 ) , .A2( u2_u8_u3_n178 ) );
  AND3_X1 u2_u8_u3_U41 (.ZN( u2_u8_u3_n118 ) , .A2( u2_u8_u3_n124 ) , .A1( u2_u8_u3_n144 ) , .A3( u2_u8_u3_n152 ) );
  INV_X1 u2_u8_u3_U42 (.A( u2_u8_u3_n121 ) , .ZN( u2_u8_u3_n164 ) );
  NAND2_X1 u2_u8_u3_U43 (.ZN( u2_u8_u3_n133 ) , .A1( u2_u8_u3_n154 ) , .A2( u2_u8_u3_n164 ) );
  OAI211_X1 u2_u8_u3_U44 (.B( u2_u8_u3_n127 ) , .ZN( u2_u8_u3_n139 ) , .C1( u2_u8_u3_n150 ) , .C2( u2_u8_u3_n154 ) , .A( u2_u8_u3_n184 ) );
  INV_X1 u2_u8_u3_U45 (.A( u2_u8_u3_n125 ) , .ZN( u2_u8_u3_n184 ) );
  AOI221_X1 u2_u8_u3_U46 (.A( u2_u8_u3_n126 ) , .ZN( u2_u8_u3_n127 ) , .C2( u2_u8_u3_n132 ) , .C1( u2_u8_u3_n169 ) , .B2( u2_u8_u3_n170 ) , .B1( u2_u8_u3_n174 ) );
  OAI22_X1 u2_u8_u3_U47 (.A1( u2_u8_u3_n124 ) , .ZN( u2_u8_u3_n125 ) , .B2( u2_u8_u3_n145 ) , .A2( u2_u8_u3_n165 ) , .B1( u2_u8_u3_n167 ) );
  NOR2_X1 u2_u8_u3_U48 (.A1( u2_u8_u3_n113 ) , .ZN( u2_u8_u3_n131 ) , .A2( u2_u8_u3_n154 ) );
  NAND2_X1 u2_u8_u3_U49 (.A1( u2_u8_u3_n103 ) , .ZN( u2_u8_u3_n150 ) , .A2( u2_u8_u3_n99 ) );
  INV_X1 u2_u8_u3_U5 (.A( u2_u8_u3_n117 ) , .ZN( u2_u8_u3_n178 ) );
  NAND2_X1 u2_u8_u3_U50 (.A2( u2_u8_u3_n102 ) , .ZN( u2_u8_u3_n155 ) , .A1( u2_u8_u3_n97 ) );
  INV_X1 u2_u8_u3_U51 (.A( u2_u8_u3_n141 ) , .ZN( u2_u8_u3_n167 ) );
  AOI21_X1 u2_u8_u3_U52 (.B2( u2_u8_u3_n114 ) , .B1( u2_u8_u3_n146 ) , .A( u2_u8_u3_n154 ) , .ZN( u2_u8_u3_n94 ) );
  AOI21_X1 u2_u8_u3_U53 (.ZN( u2_u8_u3_n110 ) , .B2( u2_u8_u3_n142 ) , .B1( u2_u8_u3_n186 ) , .A( u2_u8_u3_n95 ) );
  INV_X1 u2_u8_u3_U54 (.A( u2_u8_u3_n145 ) , .ZN( u2_u8_u3_n186 ) );
  AOI21_X1 u2_u8_u3_U55 (.B1( u2_u8_u3_n124 ) , .A( u2_u8_u3_n149 ) , .B2( u2_u8_u3_n155 ) , .ZN( u2_u8_u3_n95 ) );
  INV_X1 u2_u8_u3_U56 (.A( u2_u8_u3_n149 ) , .ZN( u2_u8_u3_n169 ) );
  NAND2_X1 u2_u8_u3_U57 (.ZN( u2_u8_u3_n124 ) , .A1( u2_u8_u3_n96 ) , .A2( u2_u8_u3_n97 ) );
  NAND2_X1 u2_u8_u3_U58 (.A2( u2_u8_u3_n100 ) , .ZN( u2_u8_u3_n146 ) , .A1( u2_u8_u3_n96 ) );
  NAND2_X1 u2_u8_u3_U59 (.A1( u2_u8_u3_n101 ) , .ZN( u2_u8_u3_n145 ) , .A2( u2_u8_u3_n99 ) );
  AOI221_X1 u2_u8_u3_U6 (.A( u2_u8_u3_n131 ) , .C2( u2_u8_u3_n132 ) , .C1( u2_u8_u3_n133 ) , .ZN( u2_u8_u3_n134 ) , .B1( u2_u8_u3_n143 ) , .B2( u2_u8_u3_n177 ) );
  NAND2_X1 u2_u8_u3_U60 (.A1( u2_u8_u3_n100 ) , .ZN( u2_u8_u3_n156 ) , .A2( u2_u8_u3_n99 ) );
  NAND2_X1 u2_u8_u3_U61 (.A2( u2_u8_u3_n101 ) , .A1( u2_u8_u3_n104 ) , .ZN( u2_u8_u3_n148 ) );
  NAND2_X1 u2_u8_u3_U62 (.A1( u2_u8_u3_n100 ) , .A2( u2_u8_u3_n102 ) , .ZN( u2_u8_u3_n128 ) );
  NAND2_X1 u2_u8_u3_U63 (.A2( u2_u8_u3_n101 ) , .A1( u2_u8_u3_n102 ) , .ZN( u2_u8_u3_n152 ) );
  NAND2_X1 u2_u8_u3_U64 (.A2( u2_u8_u3_n101 ) , .ZN( u2_u8_u3_n114 ) , .A1( u2_u8_u3_n96 ) );
  NAND2_X1 u2_u8_u3_U65 (.ZN( u2_u8_u3_n107 ) , .A1( u2_u8_u3_n97 ) , .A2( u2_u8_u3_n99 ) );
  NAND2_X1 u2_u8_u3_U66 (.A2( u2_u8_u3_n100 ) , .A1( u2_u8_u3_n104 ) , .ZN( u2_u8_u3_n113 ) );
  NAND2_X1 u2_u8_u3_U67 (.A1( u2_u8_u3_n104 ) , .ZN( u2_u8_u3_n153 ) , .A2( u2_u8_u3_n97 ) );
  NAND2_X1 u2_u8_u3_U68 (.A2( u2_u8_u3_n103 ) , .A1( u2_u8_u3_n104 ) , .ZN( u2_u8_u3_n130 ) );
  NAND2_X1 u2_u8_u3_U69 (.A2( u2_u8_u3_n103 ) , .ZN( u2_u8_u3_n144 ) , .A1( u2_u8_u3_n96 ) );
  OAI22_X1 u2_u8_u3_U7 (.B2( u2_u8_u3_n147 ) , .A2( u2_u8_u3_n148 ) , .ZN( u2_u8_u3_n160 ) , .B1( u2_u8_u3_n165 ) , .A1( u2_u8_u3_n168 ) );
  NAND2_X1 u2_u8_u3_U70 (.A1( u2_u8_u3_n102 ) , .A2( u2_u8_u3_n103 ) , .ZN( u2_u8_u3_n108 ) );
  NOR2_X1 u2_u8_u3_U71 (.A2( u2_u8_X_19 ) , .A1( u2_u8_X_20 ) , .ZN( u2_u8_u3_n99 ) );
  NOR2_X1 u2_u8_u3_U72 (.A2( u2_u8_X_21 ) , .A1( u2_u8_X_24 ) , .ZN( u2_u8_u3_n103 ) );
  NOR2_X1 u2_u8_u3_U73 (.A2( u2_u8_X_24 ) , .A1( u2_u8_u3_n171 ) , .ZN( u2_u8_u3_n97 ) );
  NOR2_X1 u2_u8_u3_U74 (.A2( u2_u8_X_23 ) , .ZN( u2_u8_u3_n141 ) , .A1( u2_u8_u3_n166 ) );
  NOR2_X1 u2_u8_u3_U75 (.A2( u2_u8_X_19 ) , .A1( u2_u8_u3_n172 ) , .ZN( u2_u8_u3_n96 ) );
  NAND2_X1 u2_u8_u3_U76 (.A1( u2_u8_X_22 ) , .A2( u2_u8_X_23 ) , .ZN( u2_u8_u3_n154 ) );
  NAND2_X1 u2_u8_u3_U77 (.A1( u2_u8_X_23 ) , .ZN( u2_u8_u3_n149 ) , .A2( u2_u8_u3_n166 ) );
  NOR2_X1 u2_u8_u3_U78 (.A2( u2_u8_X_22 ) , .A1( u2_u8_X_23 ) , .ZN( u2_u8_u3_n121 ) );
  AND2_X1 u2_u8_u3_U79 (.A1( u2_u8_X_24 ) , .ZN( u2_u8_u3_n101 ) , .A2( u2_u8_u3_n171 ) );
  AND3_X1 u2_u8_u3_U8 (.A3( u2_u8_u3_n144 ) , .A2( u2_u8_u3_n145 ) , .A1( u2_u8_u3_n146 ) , .ZN( u2_u8_u3_n147 ) );
  AND2_X1 u2_u8_u3_U80 (.A1( u2_u8_X_19 ) , .ZN( u2_u8_u3_n102 ) , .A2( u2_u8_u3_n172 ) );
  AND2_X1 u2_u8_u3_U81 (.A1( u2_u8_X_21 ) , .A2( u2_u8_X_24 ) , .ZN( u2_u8_u3_n100 ) );
  AND2_X1 u2_u8_u3_U82 (.A2( u2_u8_X_19 ) , .A1( u2_u8_X_20 ) , .ZN( u2_u8_u3_n104 ) );
  INV_X1 u2_u8_u3_U83 (.A( u2_u8_X_22 ) , .ZN( u2_u8_u3_n166 ) );
  INV_X1 u2_u8_u3_U84 (.A( u2_u8_X_21 ) , .ZN( u2_u8_u3_n171 ) );
  INV_X1 u2_u8_u3_U85 (.A( u2_u8_X_20 ) , .ZN( u2_u8_u3_n172 ) );
  OR4_X1 u2_u8_u3_U86 (.ZN( u2_out8_10 ) , .A4( u2_u8_u3_n136 ) , .A3( u2_u8_u3_n137 ) , .A1( u2_u8_u3_n138 ) , .A2( u2_u8_u3_n139 ) );
  OAI222_X1 u2_u8_u3_U87 (.C1( u2_u8_u3_n128 ) , .ZN( u2_u8_u3_n137 ) , .B1( u2_u8_u3_n148 ) , .A2( u2_u8_u3_n150 ) , .B2( u2_u8_u3_n154 ) , .C2( u2_u8_u3_n164 ) , .A1( u2_u8_u3_n167 ) );
  OAI221_X1 u2_u8_u3_U88 (.A( u2_u8_u3_n134 ) , .B2( u2_u8_u3_n135 ) , .ZN( u2_u8_u3_n136 ) , .C1( u2_u8_u3_n149 ) , .B1( u2_u8_u3_n151 ) , .C2( u2_u8_u3_n183 ) );
  NAND4_X1 u2_u8_u3_U89 (.ZN( u2_out8_26 ) , .A4( u2_u8_u3_n109 ) , .A3( u2_u8_u3_n110 ) , .A2( u2_u8_u3_n111 ) , .A1( u2_u8_u3_n173 ) );
  INV_X1 u2_u8_u3_U9 (.A( u2_u8_u3_n143 ) , .ZN( u2_u8_u3_n168 ) );
  INV_X1 u2_u8_u3_U90 (.ZN( u2_u8_u3_n173 ) , .A( u2_u8_u3_n94 ) );
  OAI21_X1 u2_u8_u3_U91 (.ZN( u2_u8_u3_n111 ) , .B2( u2_u8_u3_n117 ) , .A( u2_u8_u3_n133 ) , .B1( u2_u8_u3_n176 ) );
  NAND4_X1 u2_u8_u3_U92 (.ZN( u2_out8_20 ) , .A4( u2_u8_u3_n122 ) , .A3( u2_u8_u3_n123 ) , .A1( u2_u8_u3_n175 ) , .A2( u2_u8_u3_n180 ) );
  INV_X1 u2_u8_u3_U93 (.A( u2_u8_u3_n126 ) , .ZN( u2_u8_u3_n180 ) );
  INV_X1 u2_u8_u3_U94 (.A( u2_u8_u3_n112 ) , .ZN( u2_u8_u3_n175 ) );
  NAND4_X1 u2_u8_u3_U95 (.ZN( u2_out8_1 ) , .A4( u2_u8_u3_n161 ) , .A3( u2_u8_u3_n162 ) , .A2( u2_u8_u3_n163 ) , .A1( u2_u8_u3_n185 ) );
  NAND2_X1 u2_u8_u3_U96 (.ZN( u2_u8_u3_n163 ) , .A2( u2_u8_u3_n170 ) , .A1( u2_u8_u3_n176 ) );
  AOI22_X1 u2_u8_u3_U97 (.B2( u2_u8_u3_n140 ) , .B1( u2_u8_u3_n141 ) , .A2( u2_u8_u3_n142 ) , .ZN( u2_u8_u3_n162 ) , .A1( u2_u8_u3_n177 ) );
  NAND3_X1 u2_u8_u3_U98 (.A1( u2_u8_u3_n114 ) , .ZN( u2_u8_u3_n115 ) , .A2( u2_u8_u3_n145 ) , .A3( u2_u8_u3_n153 ) );
  NAND3_X1 u2_u8_u3_U99 (.ZN( u2_u8_u3_n129 ) , .A2( u2_u8_u3_n144 ) , .A1( u2_u8_u3_n153 ) , .A3( u2_u8_u3_n182 ) );
  OAI22_X1 u2_u8_u4_U10 (.B2( u2_u8_u4_n135 ) , .ZN( u2_u8_u4_n137 ) , .B1( u2_u8_u4_n153 ) , .A1( u2_u8_u4_n155 ) , .A2( u2_u8_u4_n171 ) );
  AND3_X1 u2_u8_u4_U11 (.A2( u2_u8_u4_n134 ) , .ZN( u2_u8_u4_n135 ) , .A3( u2_u8_u4_n145 ) , .A1( u2_u8_u4_n157 ) );
  NAND2_X1 u2_u8_u4_U12 (.ZN( u2_u8_u4_n132 ) , .A2( u2_u8_u4_n170 ) , .A1( u2_u8_u4_n173 ) );
  AOI21_X1 u2_u8_u4_U13 (.B2( u2_u8_u4_n160 ) , .B1( u2_u8_u4_n161 ) , .ZN( u2_u8_u4_n162 ) , .A( u2_u8_u4_n170 ) );
  AOI21_X1 u2_u8_u4_U14 (.ZN( u2_u8_u4_n107 ) , .B2( u2_u8_u4_n143 ) , .A( u2_u8_u4_n174 ) , .B1( u2_u8_u4_n184 ) );
  AOI21_X1 u2_u8_u4_U15 (.B2( u2_u8_u4_n158 ) , .B1( u2_u8_u4_n159 ) , .ZN( u2_u8_u4_n163 ) , .A( u2_u8_u4_n174 ) );
  AOI21_X1 u2_u8_u4_U16 (.A( u2_u8_u4_n153 ) , .B2( u2_u8_u4_n154 ) , .B1( u2_u8_u4_n155 ) , .ZN( u2_u8_u4_n165 ) );
  AOI21_X1 u2_u8_u4_U17 (.A( u2_u8_u4_n156 ) , .B2( u2_u8_u4_n157 ) , .ZN( u2_u8_u4_n164 ) , .B1( u2_u8_u4_n184 ) );
  INV_X1 u2_u8_u4_U18 (.A( u2_u8_u4_n138 ) , .ZN( u2_u8_u4_n170 ) );
  AND2_X1 u2_u8_u4_U19 (.A2( u2_u8_u4_n120 ) , .ZN( u2_u8_u4_n155 ) , .A1( u2_u8_u4_n160 ) );
  INV_X1 u2_u8_u4_U20 (.A( u2_u8_u4_n156 ) , .ZN( u2_u8_u4_n175 ) );
  NAND2_X1 u2_u8_u4_U21 (.A2( u2_u8_u4_n118 ) , .ZN( u2_u8_u4_n131 ) , .A1( u2_u8_u4_n147 ) );
  NAND2_X1 u2_u8_u4_U22 (.A1( u2_u8_u4_n119 ) , .A2( u2_u8_u4_n120 ) , .ZN( u2_u8_u4_n130 ) );
  NAND2_X1 u2_u8_u4_U23 (.ZN( u2_u8_u4_n117 ) , .A2( u2_u8_u4_n118 ) , .A1( u2_u8_u4_n148 ) );
  NAND2_X1 u2_u8_u4_U24 (.ZN( u2_u8_u4_n129 ) , .A1( u2_u8_u4_n134 ) , .A2( u2_u8_u4_n148 ) );
  AND3_X1 u2_u8_u4_U25 (.A1( u2_u8_u4_n119 ) , .A2( u2_u8_u4_n143 ) , .A3( u2_u8_u4_n154 ) , .ZN( u2_u8_u4_n161 ) );
  AND2_X1 u2_u8_u4_U26 (.A1( u2_u8_u4_n145 ) , .A2( u2_u8_u4_n147 ) , .ZN( u2_u8_u4_n159 ) );
  OR3_X1 u2_u8_u4_U27 (.A3( u2_u8_u4_n114 ) , .A2( u2_u8_u4_n115 ) , .A1( u2_u8_u4_n116 ) , .ZN( u2_u8_u4_n136 ) );
  AOI21_X1 u2_u8_u4_U28 (.A( u2_u8_u4_n113 ) , .ZN( u2_u8_u4_n116 ) , .B2( u2_u8_u4_n173 ) , .B1( u2_u8_u4_n174 ) );
  AOI21_X1 u2_u8_u4_U29 (.ZN( u2_u8_u4_n115 ) , .B2( u2_u8_u4_n145 ) , .B1( u2_u8_u4_n146 ) , .A( u2_u8_u4_n156 ) );
  NOR2_X1 u2_u8_u4_U3 (.ZN( u2_u8_u4_n121 ) , .A1( u2_u8_u4_n181 ) , .A2( u2_u8_u4_n182 ) );
  OAI22_X1 u2_u8_u4_U30 (.ZN( u2_u8_u4_n114 ) , .A2( u2_u8_u4_n121 ) , .B1( u2_u8_u4_n160 ) , .B2( u2_u8_u4_n170 ) , .A1( u2_u8_u4_n171 ) );
  INV_X1 u2_u8_u4_U31 (.A( u2_u8_u4_n158 ) , .ZN( u2_u8_u4_n182 ) );
  INV_X1 u2_u8_u4_U32 (.ZN( u2_u8_u4_n181 ) , .A( u2_u8_u4_n96 ) );
  INV_X1 u2_u8_u4_U33 (.A( u2_u8_u4_n144 ) , .ZN( u2_u8_u4_n179 ) );
  INV_X1 u2_u8_u4_U34 (.A( u2_u8_u4_n157 ) , .ZN( u2_u8_u4_n178 ) );
  NAND2_X1 u2_u8_u4_U35 (.A2( u2_u8_u4_n154 ) , .A1( u2_u8_u4_n96 ) , .ZN( u2_u8_u4_n97 ) );
  INV_X1 u2_u8_u4_U36 (.ZN( u2_u8_u4_n186 ) , .A( u2_u8_u4_n95 ) );
  OAI221_X1 u2_u8_u4_U37 (.C1( u2_u8_u4_n134 ) , .B1( u2_u8_u4_n158 ) , .B2( u2_u8_u4_n171 ) , .C2( u2_u8_u4_n173 ) , .A( u2_u8_u4_n94 ) , .ZN( u2_u8_u4_n95 ) );
  AOI222_X1 u2_u8_u4_U38 (.B2( u2_u8_u4_n132 ) , .A1( u2_u8_u4_n138 ) , .C2( u2_u8_u4_n175 ) , .A2( u2_u8_u4_n179 ) , .C1( u2_u8_u4_n181 ) , .B1( u2_u8_u4_n185 ) , .ZN( u2_u8_u4_n94 ) );
  INV_X1 u2_u8_u4_U39 (.A( u2_u8_u4_n113 ) , .ZN( u2_u8_u4_n185 ) );
  INV_X1 u2_u8_u4_U4 (.A( u2_u8_u4_n117 ) , .ZN( u2_u8_u4_n184 ) );
  INV_X1 u2_u8_u4_U40 (.A( u2_u8_u4_n143 ) , .ZN( u2_u8_u4_n183 ) );
  NOR2_X1 u2_u8_u4_U41 (.ZN( u2_u8_u4_n138 ) , .A1( u2_u8_u4_n168 ) , .A2( u2_u8_u4_n169 ) );
  NOR2_X1 u2_u8_u4_U42 (.A1( u2_u8_u4_n150 ) , .A2( u2_u8_u4_n152 ) , .ZN( u2_u8_u4_n153 ) );
  NOR2_X1 u2_u8_u4_U43 (.A2( u2_u8_u4_n128 ) , .A1( u2_u8_u4_n138 ) , .ZN( u2_u8_u4_n156 ) );
  AOI22_X1 u2_u8_u4_U44 (.B2( u2_u8_u4_n122 ) , .A1( u2_u8_u4_n123 ) , .ZN( u2_u8_u4_n124 ) , .B1( u2_u8_u4_n128 ) , .A2( u2_u8_u4_n172 ) );
  INV_X1 u2_u8_u4_U45 (.A( u2_u8_u4_n153 ) , .ZN( u2_u8_u4_n172 ) );
  NAND2_X1 u2_u8_u4_U46 (.A2( u2_u8_u4_n120 ) , .ZN( u2_u8_u4_n123 ) , .A1( u2_u8_u4_n161 ) );
  AOI22_X1 u2_u8_u4_U47 (.B2( u2_u8_u4_n132 ) , .A2( u2_u8_u4_n133 ) , .ZN( u2_u8_u4_n140 ) , .A1( u2_u8_u4_n150 ) , .B1( u2_u8_u4_n179 ) );
  NAND2_X1 u2_u8_u4_U48 (.ZN( u2_u8_u4_n133 ) , .A2( u2_u8_u4_n146 ) , .A1( u2_u8_u4_n154 ) );
  NAND2_X1 u2_u8_u4_U49 (.A1( u2_u8_u4_n103 ) , .ZN( u2_u8_u4_n154 ) , .A2( u2_u8_u4_n98 ) );
  NOR4_X1 u2_u8_u4_U5 (.A4( u2_u8_u4_n106 ) , .A3( u2_u8_u4_n107 ) , .A2( u2_u8_u4_n108 ) , .A1( u2_u8_u4_n109 ) , .ZN( u2_u8_u4_n110 ) );
  NAND2_X1 u2_u8_u4_U50 (.A1( u2_u8_u4_n101 ) , .ZN( u2_u8_u4_n158 ) , .A2( u2_u8_u4_n99 ) );
  AOI21_X1 u2_u8_u4_U51 (.ZN( u2_u8_u4_n127 ) , .A( u2_u8_u4_n136 ) , .B2( u2_u8_u4_n150 ) , .B1( u2_u8_u4_n180 ) );
  INV_X1 u2_u8_u4_U52 (.A( u2_u8_u4_n160 ) , .ZN( u2_u8_u4_n180 ) );
  NAND2_X1 u2_u8_u4_U53 (.A2( u2_u8_u4_n104 ) , .A1( u2_u8_u4_n105 ) , .ZN( u2_u8_u4_n146 ) );
  NAND2_X1 u2_u8_u4_U54 (.A2( u2_u8_u4_n101 ) , .A1( u2_u8_u4_n102 ) , .ZN( u2_u8_u4_n160 ) );
  NAND2_X1 u2_u8_u4_U55 (.ZN( u2_u8_u4_n134 ) , .A1( u2_u8_u4_n98 ) , .A2( u2_u8_u4_n99 ) );
  NAND2_X1 u2_u8_u4_U56 (.A1( u2_u8_u4_n103 ) , .A2( u2_u8_u4_n104 ) , .ZN( u2_u8_u4_n143 ) );
  NAND2_X1 u2_u8_u4_U57 (.A2( u2_u8_u4_n105 ) , .ZN( u2_u8_u4_n145 ) , .A1( u2_u8_u4_n98 ) );
  NAND2_X1 u2_u8_u4_U58 (.A1( u2_u8_u4_n100 ) , .A2( u2_u8_u4_n105 ) , .ZN( u2_u8_u4_n120 ) );
  NAND2_X1 u2_u8_u4_U59 (.A1( u2_u8_u4_n102 ) , .A2( u2_u8_u4_n104 ) , .ZN( u2_u8_u4_n148 ) );
  AOI21_X1 u2_u8_u4_U6 (.ZN( u2_u8_u4_n106 ) , .B2( u2_u8_u4_n146 ) , .B1( u2_u8_u4_n158 ) , .A( u2_u8_u4_n170 ) );
  NAND2_X1 u2_u8_u4_U60 (.A2( u2_u8_u4_n100 ) , .A1( u2_u8_u4_n103 ) , .ZN( u2_u8_u4_n157 ) );
  INV_X1 u2_u8_u4_U61 (.A( u2_u8_u4_n150 ) , .ZN( u2_u8_u4_n173 ) );
  INV_X1 u2_u8_u4_U62 (.A( u2_u8_u4_n152 ) , .ZN( u2_u8_u4_n171 ) );
  NAND2_X1 u2_u8_u4_U63 (.A1( u2_u8_u4_n100 ) , .ZN( u2_u8_u4_n118 ) , .A2( u2_u8_u4_n99 ) );
  NAND2_X1 u2_u8_u4_U64 (.A2( u2_u8_u4_n100 ) , .A1( u2_u8_u4_n102 ) , .ZN( u2_u8_u4_n144 ) );
  NAND2_X1 u2_u8_u4_U65 (.A2( u2_u8_u4_n101 ) , .A1( u2_u8_u4_n105 ) , .ZN( u2_u8_u4_n96 ) );
  INV_X1 u2_u8_u4_U66 (.A( u2_u8_u4_n128 ) , .ZN( u2_u8_u4_n174 ) );
  NAND2_X1 u2_u8_u4_U67 (.A2( u2_u8_u4_n102 ) , .ZN( u2_u8_u4_n119 ) , .A1( u2_u8_u4_n98 ) );
  NAND2_X1 u2_u8_u4_U68 (.A2( u2_u8_u4_n101 ) , .A1( u2_u8_u4_n103 ) , .ZN( u2_u8_u4_n147 ) );
  NAND2_X1 u2_u8_u4_U69 (.A2( u2_u8_u4_n104 ) , .ZN( u2_u8_u4_n113 ) , .A1( u2_u8_u4_n99 ) );
  AOI21_X1 u2_u8_u4_U7 (.ZN( u2_u8_u4_n108 ) , .B2( u2_u8_u4_n134 ) , .B1( u2_u8_u4_n155 ) , .A( u2_u8_u4_n156 ) );
  NOR2_X1 u2_u8_u4_U70 (.A2( u2_u8_X_28 ) , .ZN( u2_u8_u4_n150 ) , .A1( u2_u8_u4_n168 ) );
  NOR2_X1 u2_u8_u4_U71 (.A2( u2_u8_X_29 ) , .ZN( u2_u8_u4_n152 ) , .A1( u2_u8_u4_n169 ) );
  NOR2_X1 u2_u8_u4_U72 (.A2( u2_u8_X_30 ) , .ZN( u2_u8_u4_n105 ) , .A1( u2_u8_u4_n176 ) );
  NOR2_X1 u2_u8_u4_U73 (.A2( u2_u8_X_26 ) , .ZN( u2_u8_u4_n100 ) , .A1( u2_u8_u4_n177 ) );
  NOR2_X1 u2_u8_u4_U74 (.A2( u2_u8_X_28 ) , .A1( u2_u8_X_29 ) , .ZN( u2_u8_u4_n128 ) );
  NOR2_X1 u2_u8_u4_U75 (.A2( u2_u8_X_27 ) , .A1( u2_u8_X_30 ) , .ZN( u2_u8_u4_n102 ) );
  NOR2_X1 u2_u8_u4_U76 (.A2( u2_u8_X_25 ) , .A1( u2_u8_X_26 ) , .ZN( u2_u8_u4_n98 ) );
  AND2_X1 u2_u8_u4_U77 (.A2( u2_u8_X_25 ) , .A1( u2_u8_X_26 ) , .ZN( u2_u8_u4_n104 ) );
  AND2_X1 u2_u8_u4_U78 (.A1( u2_u8_X_30 ) , .A2( u2_u8_u4_n176 ) , .ZN( u2_u8_u4_n99 ) );
  AND2_X1 u2_u8_u4_U79 (.A1( u2_u8_X_26 ) , .ZN( u2_u8_u4_n101 ) , .A2( u2_u8_u4_n177 ) );
  AOI21_X1 u2_u8_u4_U8 (.ZN( u2_u8_u4_n109 ) , .A( u2_u8_u4_n153 ) , .B1( u2_u8_u4_n159 ) , .B2( u2_u8_u4_n184 ) );
  AND2_X1 u2_u8_u4_U80 (.A1( u2_u8_X_27 ) , .A2( u2_u8_X_30 ) , .ZN( u2_u8_u4_n103 ) );
  INV_X1 u2_u8_u4_U81 (.A( u2_u8_X_28 ) , .ZN( u2_u8_u4_n169 ) );
  INV_X1 u2_u8_u4_U82 (.A( u2_u8_X_29 ) , .ZN( u2_u8_u4_n168 ) );
  INV_X1 u2_u8_u4_U83 (.A( u2_u8_X_25 ) , .ZN( u2_u8_u4_n177 ) );
  INV_X1 u2_u8_u4_U84 (.A( u2_u8_X_27 ) , .ZN( u2_u8_u4_n176 ) );
  NAND4_X1 u2_u8_u4_U85 (.ZN( u2_out8_25 ) , .A4( u2_u8_u4_n139 ) , .A3( u2_u8_u4_n140 ) , .A2( u2_u8_u4_n141 ) , .A1( u2_u8_u4_n142 ) );
  OAI21_X1 u2_u8_u4_U86 (.B2( u2_u8_u4_n131 ) , .ZN( u2_u8_u4_n141 ) , .A( u2_u8_u4_n175 ) , .B1( u2_u8_u4_n183 ) );
  OAI21_X1 u2_u8_u4_U87 (.A( u2_u8_u4_n128 ) , .B2( u2_u8_u4_n129 ) , .B1( u2_u8_u4_n130 ) , .ZN( u2_u8_u4_n142 ) );
  NAND4_X1 u2_u8_u4_U88 (.ZN( u2_out8_14 ) , .A4( u2_u8_u4_n124 ) , .A3( u2_u8_u4_n125 ) , .A2( u2_u8_u4_n126 ) , .A1( u2_u8_u4_n127 ) );
  AOI22_X1 u2_u8_u4_U89 (.B2( u2_u8_u4_n117 ) , .ZN( u2_u8_u4_n126 ) , .A1( u2_u8_u4_n129 ) , .B1( u2_u8_u4_n152 ) , .A2( u2_u8_u4_n175 ) );
  AOI211_X1 u2_u8_u4_U9 (.B( u2_u8_u4_n136 ) , .A( u2_u8_u4_n137 ) , .C2( u2_u8_u4_n138 ) , .ZN( u2_u8_u4_n139 ) , .C1( u2_u8_u4_n182 ) );
  AOI22_X1 u2_u8_u4_U90 (.ZN( u2_u8_u4_n125 ) , .B2( u2_u8_u4_n131 ) , .A2( u2_u8_u4_n132 ) , .B1( u2_u8_u4_n138 ) , .A1( u2_u8_u4_n178 ) );
  NAND4_X1 u2_u8_u4_U91 (.ZN( u2_out8_8 ) , .A4( u2_u8_u4_n110 ) , .A3( u2_u8_u4_n111 ) , .A2( u2_u8_u4_n112 ) , .A1( u2_u8_u4_n186 ) );
  NAND2_X1 u2_u8_u4_U92 (.ZN( u2_u8_u4_n112 ) , .A2( u2_u8_u4_n130 ) , .A1( u2_u8_u4_n150 ) );
  AOI22_X1 u2_u8_u4_U93 (.ZN( u2_u8_u4_n111 ) , .B2( u2_u8_u4_n132 ) , .A1( u2_u8_u4_n152 ) , .B1( u2_u8_u4_n178 ) , .A2( u2_u8_u4_n97 ) );
  AOI22_X1 u2_u8_u4_U94 (.B2( u2_u8_u4_n149 ) , .B1( u2_u8_u4_n150 ) , .A2( u2_u8_u4_n151 ) , .A1( u2_u8_u4_n152 ) , .ZN( u2_u8_u4_n167 ) );
  NOR4_X1 u2_u8_u4_U95 (.A4( u2_u8_u4_n162 ) , .A3( u2_u8_u4_n163 ) , .A2( u2_u8_u4_n164 ) , .A1( u2_u8_u4_n165 ) , .ZN( u2_u8_u4_n166 ) );
  NAND3_X1 u2_u8_u4_U96 (.ZN( u2_out8_3 ) , .A3( u2_u8_u4_n166 ) , .A1( u2_u8_u4_n167 ) , .A2( u2_u8_u4_n186 ) );
  NAND3_X1 u2_u8_u4_U97 (.A3( u2_u8_u4_n146 ) , .A2( u2_u8_u4_n147 ) , .A1( u2_u8_u4_n148 ) , .ZN( u2_u8_u4_n149 ) );
  NAND3_X1 u2_u8_u4_U98 (.A3( u2_u8_u4_n143 ) , .A2( u2_u8_u4_n144 ) , .A1( u2_u8_u4_n145 ) , .ZN( u2_u8_u4_n151 ) );
  NAND3_X1 u2_u8_u4_U99 (.A3( u2_u8_u4_n121 ) , .ZN( u2_u8_u4_n122 ) , .A2( u2_u8_u4_n144 ) , .A1( u2_u8_u4_n154 ) );
  XOR2_X1 u2_u9_U11 (.B( u2_K10_44 ) , .A( u2_R8_29 ) , .Z( u2_u9_X_44 ) );
  XOR2_X1 u2_u9_U12 (.B( u2_K10_43 ) , .A( u2_R8_28 ) , .Z( u2_u9_X_43 ) );
  XOR2_X1 u2_u9_U13 (.B( u2_K10_42 ) , .A( u2_R8_29 ) , .Z( u2_u9_X_42 ) );
  XOR2_X1 u2_u9_U14 (.B( u2_K10_41 ) , .A( u2_R8_28 ) , .Z( u2_u9_X_41 ) );
  XOR2_X1 u2_u9_U15 (.B( u2_K10_40 ) , .A( u2_R8_27 ) , .Z( u2_u9_X_40 ) );
  XOR2_X1 u2_u9_U17 (.B( u2_K10_39 ) , .A( u2_R8_26 ) , .Z( u2_u9_X_39 ) );
  XOR2_X1 u2_u9_U18 (.B( u2_K10_38 ) , .A( u2_R8_25 ) , .Z( u2_u9_X_38 ) );
  XOR2_X1 u2_u9_U19 (.B( u2_K10_37 ) , .A( u2_R8_24 ) , .Z( u2_u9_X_37 ) );
  XOR2_X1 u2_u9_U20 (.B( u2_K10_36 ) , .A( u2_R8_25 ) , .Z( u2_u9_X_36 ) );
  XOR2_X1 u2_u9_U21 (.B( u2_K10_35 ) , .A( u2_R8_24 ) , .Z( u2_u9_X_35 ) );
  XOR2_X1 u2_u9_U23 (.B( u2_K10_33 ) , .A( u2_R8_22 ) , .Z( u2_u9_X_33 ) );
  XOR2_X1 u2_u9_U25 (.B( u2_K10_31 ) , .A( u2_R8_20 ) , .Z( u2_u9_X_31 ) );
  XOR2_X1 u2_u9_U27 (.B( u2_K10_2 ) , .A( u2_R8_1 ) , .Z( u2_u9_X_2 ) );
  XOR2_X1 u2_u9_U38 (.B( u2_K10_1 ) , .A( u2_R8_32 ) , .Z( u2_u9_X_1 ) );
  XOR2_X1 u2_u9_U5 (.B( u2_K10_5 ) , .A( u2_R8_4 ) , .Z( u2_u9_X_5 ) );
  XOR2_X1 u2_u9_U7 (.B( u2_K10_48 ) , .A( u2_R8_1 ) , .Z( u2_u9_X_48 ) );
  XOR2_X1 u2_u9_U8 (.B( u2_K10_47 ) , .A( u2_R8_32 ) , .Z( u2_u9_X_47 ) );
  AND3_X1 u2_u9_u0_U10 (.A2( u2_u9_u0_n112 ) , .ZN( u2_u9_u0_n127 ) , .A3( u2_u9_u0_n130 ) , .A1( u2_u9_u0_n148 ) );
  NAND2_X1 u2_u9_u0_U11 (.ZN( u2_u9_u0_n113 ) , .A1( u2_u9_u0_n139 ) , .A2( u2_u9_u0_n149 ) );
  AND2_X1 u2_u9_u0_U12 (.ZN( u2_u9_u0_n107 ) , .A1( u2_u9_u0_n130 ) , .A2( u2_u9_u0_n140 ) );
  AND2_X1 u2_u9_u0_U13 (.A2( u2_u9_u0_n129 ) , .A1( u2_u9_u0_n130 ) , .ZN( u2_u9_u0_n151 ) );
  AND2_X1 u2_u9_u0_U14 (.A1( u2_u9_u0_n108 ) , .A2( u2_u9_u0_n125 ) , .ZN( u2_u9_u0_n145 ) );
  INV_X1 u2_u9_u0_U15 (.A( u2_u9_u0_n143 ) , .ZN( u2_u9_u0_n173 ) );
  NOR2_X1 u2_u9_u0_U16 (.A2( u2_u9_u0_n136 ) , .ZN( u2_u9_u0_n147 ) , .A1( u2_u9_u0_n160 ) );
  OAI221_X1 u2_u9_u0_U17 (.C1( u2_u9_u0_n112 ) , .ZN( u2_u9_u0_n120 ) , .B1( u2_u9_u0_n138 ) , .B2( u2_u9_u0_n141 ) , .C2( u2_u9_u0_n147 ) , .A( u2_u9_u0_n172 ) );
  AOI211_X1 u2_u9_u0_U18 (.B( u2_u9_u0_n115 ) , .A( u2_u9_u0_n116 ) , .C2( u2_u9_u0_n117 ) , .C1( u2_u9_u0_n118 ) , .ZN( u2_u9_u0_n119 ) );
  OAI22_X1 u2_u9_u0_U19 (.B1( u2_u9_u0_n125 ) , .ZN( u2_u9_u0_n126 ) , .A1( u2_u9_u0_n138 ) , .A2( u2_u9_u0_n146 ) , .B2( u2_u9_u0_n147 ) );
  OAI22_X1 u2_u9_u0_U20 (.B1( u2_u9_u0_n131 ) , .A1( u2_u9_u0_n144 ) , .B2( u2_u9_u0_n147 ) , .A2( u2_u9_u0_n90 ) , .ZN( u2_u9_u0_n91 ) );
  AND3_X1 u2_u9_u0_U21 (.A3( u2_u9_u0_n121 ) , .A2( u2_u9_u0_n125 ) , .A1( u2_u9_u0_n148 ) , .ZN( u2_u9_u0_n90 ) );
  NOR2_X1 u2_u9_u0_U22 (.A1( u2_u9_u0_n163 ) , .A2( u2_u9_u0_n164 ) , .ZN( u2_u9_u0_n95 ) );
  INV_X1 u2_u9_u0_U23 (.A( u2_u9_u0_n136 ) , .ZN( u2_u9_u0_n161 ) );
  AOI22_X1 u2_u9_u0_U24 (.B2( u2_u9_u0_n109 ) , .A2( u2_u9_u0_n110 ) , .ZN( u2_u9_u0_n111 ) , .B1( u2_u9_u0_n118 ) , .A1( u2_u9_u0_n160 ) );
  INV_X1 u2_u9_u0_U25 (.A( u2_u9_u0_n118 ) , .ZN( u2_u9_u0_n158 ) );
  AOI21_X1 u2_u9_u0_U26 (.ZN( u2_u9_u0_n104 ) , .B1( u2_u9_u0_n107 ) , .B2( u2_u9_u0_n141 ) , .A( u2_u9_u0_n144 ) );
  AOI21_X1 u2_u9_u0_U27 (.B1( u2_u9_u0_n127 ) , .B2( u2_u9_u0_n129 ) , .A( u2_u9_u0_n138 ) , .ZN( u2_u9_u0_n96 ) );
  AOI21_X1 u2_u9_u0_U28 (.ZN( u2_u9_u0_n116 ) , .B2( u2_u9_u0_n142 ) , .A( u2_u9_u0_n144 ) , .B1( u2_u9_u0_n166 ) );
  NAND2_X1 u2_u9_u0_U29 (.A1( u2_u9_u0_n100 ) , .A2( u2_u9_u0_n103 ) , .ZN( u2_u9_u0_n125 ) );
  INV_X1 u2_u9_u0_U3 (.A( u2_u9_u0_n113 ) , .ZN( u2_u9_u0_n166 ) );
  NAND2_X1 u2_u9_u0_U30 (.A2( u2_u9_u0_n103 ) , .ZN( u2_u9_u0_n140 ) , .A1( u2_u9_u0_n94 ) );
  NAND2_X1 u2_u9_u0_U31 (.A1( u2_u9_u0_n101 ) , .A2( u2_u9_u0_n102 ) , .ZN( u2_u9_u0_n150 ) );
  INV_X1 u2_u9_u0_U32 (.A( u2_u9_u0_n138 ) , .ZN( u2_u9_u0_n160 ) );
  NAND2_X1 u2_u9_u0_U33 (.A2( u2_u9_u0_n102 ) , .A1( u2_u9_u0_n103 ) , .ZN( u2_u9_u0_n149 ) );
  NAND2_X1 u2_u9_u0_U34 (.A2( u2_u9_u0_n100 ) , .A1( u2_u9_u0_n101 ) , .ZN( u2_u9_u0_n139 ) );
  NAND2_X1 u2_u9_u0_U35 (.A2( u2_u9_u0_n100 ) , .ZN( u2_u9_u0_n131 ) , .A1( u2_u9_u0_n92 ) );
  NAND2_X1 u2_u9_u0_U36 (.ZN( u2_u9_u0_n108 ) , .A1( u2_u9_u0_n92 ) , .A2( u2_u9_u0_n94 ) );
  NAND2_X1 u2_u9_u0_U37 (.A2( u2_u9_u0_n102 ) , .ZN( u2_u9_u0_n114 ) , .A1( u2_u9_u0_n92 ) );
  NAND2_X1 u2_u9_u0_U38 (.A1( u2_u9_u0_n101 ) , .ZN( u2_u9_u0_n130 ) , .A2( u2_u9_u0_n94 ) );
  NAND2_X1 u2_u9_u0_U39 (.A2( u2_u9_u0_n101 ) , .ZN( u2_u9_u0_n121 ) , .A1( u2_u9_u0_n93 ) );
  AOI21_X1 u2_u9_u0_U4 (.B1( u2_u9_u0_n114 ) , .ZN( u2_u9_u0_n115 ) , .B2( u2_u9_u0_n129 ) , .A( u2_u9_u0_n161 ) );
  INV_X1 u2_u9_u0_U40 (.ZN( u2_u9_u0_n172 ) , .A( u2_u9_u0_n88 ) );
  OAI222_X1 u2_u9_u0_U41 (.C1( u2_u9_u0_n108 ) , .A1( u2_u9_u0_n125 ) , .B2( u2_u9_u0_n128 ) , .B1( u2_u9_u0_n144 ) , .A2( u2_u9_u0_n158 ) , .C2( u2_u9_u0_n161 ) , .ZN( u2_u9_u0_n88 ) );
  NAND2_X1 u2_u9_u0_U42 (.ZN( u2_u9_u0_n112 ) , .A2( u2_u9_u0_n92 ) , .A1( u2_u9_u0_n93 ) );
  OR3_X1 u2_u9_u0_U43 (.A3( u2_u9_u0_n152 ) , .A2( u2_u9_u0_n153 ) , .A1( u2_u9_u0_n154 ) , .ZN( u2_u9_u0_n155 ) );
  AOI21_X1 u2_u9_u0_U44 (.A( u2_u9_u0_n144 ) , .B2( u2_u9_u0_n145 ) , .B1( u2_u9_u0_n146 ) , .ZN( u2_u9_u0_n154 ) );
  AOI21_X1 u2_u9_u0_U45 (.B2( u2_u9_u0_n150 ) , .B1( u2_u9_u0_n151 ) , .ZN( u2_u9_u0_n152 ) , .A( u2_u9_u0_n158 ) );
  AOI21_X1 u2_u9_u0_U46 (.A( u2_u9_u0_n147 ) , .B2( u2_u9_u0_n148 ) , .B1( u2_u9_u0_n149 ) , .ZN( u2_u9_u0_n153 ) );
  AOI21_X1 u2_u9_u0_U47 (.B1( u2_u9_u0_n103 ) , .ZN( u2_u9_u0_n132 ) , .A( u2_u9_u0_n165 ) , .B2( u2_u9_u0_n93 ) );
  INV_X1 u2_u9_u0_U48 (.A( u2_u9_u0_n142 ) , .ZN( u2_u9_u0_n165 ) );
  INV_X1 u2_u9_u0_U49 (.ZN( u2_u9_u0_n171 ) , .A( u2_u9_u0_n99 ) );
  AOI21_X1 u2_u9_u0_U5 (.B2( u2_u9_u0_n131 ) , .ZN( u2_u9_u0_n134 ) , .B1( u2_u9_u0_n151 ) , .A( u2_u9_u0_n158 ) );
  OAI211_X1 u2_u9_u0_U50 (.C2( u2_u9_u0_n140 ) , .C1( u2_u9_u0_n161 ) , .A( u2_u9_u0_n169 ) , .B( u2_u9_u0_n98 ) , .ZN( u2_u9_u0_n99 ) );
  INV_X1 u2_u9_u0_U51 (.ZN( u2_u9_u0_n169 ) , .A( u2_u9_u0_n91 ) );
  AOI211_X1 u2_u9_u0_U52 (.C1( u2_u9_u0_n118 ) , .A( u2_u9_u0_n123 ) , .B( u2_u9_u0_n96 ) , .C2( u2_u9_u0_n97 ) , .ZN( u2_u9_u0_n98 ) );
  NOR2_X1 u2_u9_u0_U53 (.A2( u2_u9_X_2 ) , .ZN( u2_u9_u0_n103 ) , .A1( u2_u9_u0_n164 ) );
  NOR2_X1 u2_u9_u0_U54 (.A2( u2_u9_X_4 ) , .A1( u2_u9_X_5 ) , .ZN( u2_u9_u0_n118 ) );
  NOR2_X1 u2_u9_u0_U55 (.A2( u2_u9_X_1 ) , .A1( u2_u9_X_2 ) , .ZN( u2_u9_u0_n92 ) );
  NOR2_X1 u2_u9_u0_U56 (.A2( u2_u9_X_1 ) , .ZN( u2_u9_u0_n101 ) , .A1( u2_u9_u0_n163 ) );
  NOR2_X1 u2_u9_u0_U57 (.A2( u2_u9_X_3 ) , .A1( u2_u9_X_6 ) , .ZN( u2_u9_u0_n94 ) );
  NOR2_X1 u2_u9_u0_U58 (.A2( u2_u9_X_6 ) , .ZN( u2_u9_u0_n100 ) , .A1( u2_u9_u0_n162 ) );
  NAND2_X1 u2_u9_u0_U59 (.A2( u2_u9_X_4 ) , .A1( u2_u9_X_5 ) , .ZN( u2_u9_u0_n144 ) );
  NOR2_X1 u2_u9_u0_U6 (.A1( u2_u9_u0_n108 ) , .ZN( u2_u9_u0_n123 ) , .A2( u2_u9_u0_n158 ) );
  NOR2_X1 u2_u9_u0_U60 (.A2( u2_u9_X_5 ) , .ZN( u2_u9_u0_n136 ) , .A1( u2_u9_u0_n159 ) );
  NAND2_X1 u2_u9_u0_U61 (.A1( u2_u9_X_5 ) , .ZN( u2_u9_u0_n138 ) , .A2( u2_u9_u0_n159 ) );
  AND2_X1 u2_u9_u0_U62 (.A2( u2_u9_X_3 ) , .A1( u2_u9_X_6 ) , .ZN( u2_u9_u0_n102 ) );
  AND2_X1 u2_u9_u0_U63 (.A1( u2_u9_X_6 ) , .A2( u2_u9_u0_n162 ) , .ZN( u2_u9_u0_n93 ) );
  INV_X1 u2_u9_u0_U64 (.A( u2_u9_X_4 ) , .ZN( u2_u9_u0_n159 ) );
  INV_X1 u2_u9_u0_U65 (.A( u2_u9_X_1 ) , .ZN( u2_u9_u0_n164 ) );
  INV_X1 u2_u9_u0_U66 (.A( u2_u9_X_2 ) , .ZN( u2_u9_u0_n163 ) );
  INV_X1 u2_u9_u0_U67 (.A( u2_u9_X_3 ) , .ZN( u2_u9_u0_n162 ) );
  INV_X1 u2_u9_u0_U68 (.A( u2_u9_u0_n126 ) , .ZN( u2_u9_u0_n168 ) );
  AOI211_X1 u2_u9_u0_U69 (.B( u2_u9_u0_n133 ) , .A( u2_u9_u0_n134 ) , .C2( u2_u9_u0_n135 ) , .C1( u2_u9_u0_n136 ) , .ZN( u2_u9_u0_n137 ) );
  OAI21_X1 u2_u9_u0_U7 (.B1( u2_u9_u0_n150 ) , .B2( u2_u9_u0_n158 ) , .A( u2_u9_u0_n172 ) , .ZN( u2_u9_u0_n89 ) );
  OR4_X1 u2_u9_u0_U70 (.ZN( u2_out9_17 ) , .A4( u2_u9_u0_n122 ) , .A2( u2_u9_u0_n123 ) , .A1( u2_u9_u0_n124 ) , .A3( u2_u9_u0_n170 ) );
  AOI21_X1 u2_u9_u0_U71 (.B2( u2_u9_u0_n107 ) , .ZN( u2_u9_u0_n124 ) , .B1( u2_u9_u0_n128 ) , .A( u2_u9_u0_n161 ) );
  INV_X1 u2_u9_u0_U72 (.A( u2_u9_u0_n111 ) , .ZN( u2_u9_u0_n170 ) );
  OR4_X1 u2_u9_u0_U73 (.ZN( u2_out9_31 ) , .A4( u2_u9_u0_n155 ) , .A2( u2_u9_u0_n156 ) , .A1( u2_u9_u0_n157 ) , .A3( u2_u9_u0_n173 ) );
  AOI21_X1 u2_u9_u0_U74 (.A( u2_u9_u0_n138 ) , .B2( u2_u9_u0_n139 ) , .B1( u2_u9_u0_n140 ) , .ZN( u2_u9_u0_n157 ) );
  AOI21_X1 u2_u9_u0_U75 (.B2( u2_u9_u0_n141 ) , .B1( u2_u9_u0_n142 ) , .ZN( u2_u9_u0_n156 ) , .A( u2_u9_u0_n161 ) );
  INV_X1 u2_u9_u0_U76 (.ZN( u2_u9_u0_n174 ) , .A( u2_u9_u0_n89 ) );
  AOI211_X1 u2_u9_u0_U77 (.B( u2_u9_u0_n104 ) , .A( u2_u9_u0_n105 ) , .ZN( u2_u9_u0_n106 ) , .C2( u2_u9_u0_n113 ) , .C1( u2_u9_u0_n160 ) );
  OAI221_X1 u2_u9_u0_U78 (.C1( u2_u9_u0_n121 ) , .ZN( u2_u9_u0_n122 ) , .B2( u2_u9_u0_n127 ) , .A( u2_u9_u0_n143 ) , .B1( u2_u9_u0_n144 ) , .C2( u2_u9_u0_n147 ) );
  NOR2_X1 u2_u9_u0_U79 (.A1( u2_u9_u0_n120 ) , .ZN( u2_u9_u0_n143 ) , .A2( u2_u9_u0_n167 ) );
  AND2_X1 u2_u9_u0_U8 (.A1( u2_u9_u0_n114 ) , .A2( u2_u9_u0_n121 ) , .ZN( u2_u9_u0_n146 ) );
  AOI21_X1 u2_u9_u0_U80 (.B1( u2_u9_u0_n132 ) , .ZN( u2_u9_u0_n133 ) , .A( u2_u9_u0_n144 ) , .B2( u2_u9_u0_n166 ) );
  OAI22_X1 u2_u9_u0_U81 (.ZN( u2_u9_u0_n105 ) , .A2( u2_u9_u0_n132 ) , .B1( u2_u9_u0_n146 ) , .A1( u2_u9_u0_n147 ) , .B2( u2_u9_u0_n161 ) );
  NAND2_X1 u2_u9_u0_U82 (.ZN( u2_u9_u0_n110 ) , .A2( u2_u9_u0_n132 ) , .A1( u2_u9_u0_n145 ) );
  INV_X1 u2_u9_u0_U83 (.A( u2_u9_u0_n119 ) , .ZN( u2_u9_u0_n167 ) );
  NAND2_X1 u2_u9_u0_U84 (.ZN( u2_u9_u0_n148 ) , .A1( u2_u9_u0_n93 ) , .A2( u2_u9_u0_n95 ) );
  NAND2_X1 u2_u9_u0_U85 (.A1( u2_u9_u0_n100 ) , .ZN( u2_u9_u0_n129 ) , .A2( u2_u9_u0_n95 ) );
  NAND2_X1 u2_u9_u0_U86 (.A1( u2_u9_u0_n102 ) , .ZN( u2_u9_u0_n128 ) , .A2( u2_u9_u0_n95 ) );
  NAND2_X1 u2_u9_u0_U87 (.ZN( u2_u9_u0_n142 ) , .A1( u2_u9_u0_n94 ) , .A2( u2_u9_u0_n95 ) );
  NAND3_X1 u2_u9_u0_U88 (.ZN( u2_out9_23 ) , .A3( u2_u9_u0_n137 ) , .A1( u2_u9_u0_n168 ) , .A2( u2_u9_u0_n171 ) );
  NAND3_X1 u2_u9_u0_U89 (.A3( u2_u9_u0_n127 ) , .A2( u2_u9_u0_n128 ) , .ZN( u2_u9_u0_n135 ) , .A1( u2_u9_u0_n150 ) );
  AND2_X1 u2_u9_u0_U9 (.A1( u2_u9_u0_n131 ) , .ZN( u2_u9_u0_n141 ) , .A2( u2_u9_u0_n150 ) );
  NAND3_X1 u2_u9_u0_U90 (.ZN( u2_u9_u0_n117 ) , .A3( u2_u9_u0_n132 ) , .A2( u2_u9_u0_n139 ) , .A1( u2_u9_u0_n148 ) );
  NAND3_X1 u2_u9_u0_U91 (.ZN( u2_u9_u0_n109 ) , .A2( u2_u9_u0_n114 ) , .A3( u2_u9_u0_n140 ) , .A1( u2_u9_u0_n149 ) );
  NAND3_X1 u2_u9_u0_U92 (.ZN( u2_out9_9 ) , .A3( u2_u9_u0_n106 ) , .A2( u2_u9_u0_n171 ) , .A1( u2_u9_u0_n174 ) );
  NAND3_X1 u2_u9_u0_U93 (.A2( u2_u9_u0_n128 ) , .A1( u2_u9_u0_n132 ) , .A3( u2_u9_u0_n146 ) , .ZN( u2_u9_u0_n97 ) );
  NOR2_X1 u2_u9_u5_U10 (.ZN( u2_u9_u5_n135 ) , .A1( u2_u9_u5_n173 ) , .A2( u2_u9_u5_n176 ) );
  NOR3_X1 u2_u9_u5_U100 (.A3( u2_u9_u5_n141 ) , .A1( u2_u9_u5_n142 ) , .ZN( u2_u9_u5_n143 ) , .A2( u2_u9_u5_n191 ) );
  NAND4_X1 u2_u9_u5_U101 (.ZN( u2_out9_4 ) , .A4( u2_u9_u5_n112 ) , .A2( u2_u9_u5_n113 ) , .A1( u2_u9_u5_n114 ) , .A3( u2_u9_u5_n195 ) );
  AOI211_X1 u2_u9_u5_U102 (.A( u2_u9_u5_n110 ) , .C1( u2_u9_u5_n111 ) , .ZN( u2_u9_u5_n112 ) , .B( u2_u9_u5_n118 ) , .C2( u2_u9_u5_n177 ) );
  INV_X1 u2_u9_u5_U103 (.A( u2_u9_u5_n102 ) , .ZN( u2_u9_u5_n195 ) );
  NAND3_X1 u2_u9_u5_U104 (.A2( u2_u9_u5_n154 ) , .A3( u2_u9_u5_n158 ) , .A1( u2_u9_u5_n161 ) , .ZN( u2_u9_u5_n99 ) );
  INV_X1 u2_u9_u5_U11 (.A( u2_u9_u5_n121 ) , .ZN( u2_u9_u5_n177 ) );
  NOR2_X1 u2_u9_u5_U12 (.ZN( u2_u9_u5_n160 ) , .A2( u2_u9_u5_n173 ) , .A1( u2_u9_u5_n177 ) );
  INV_X1 u2_u9_u5_U13 (.A( u2_u9_u5_n150 ) , .ZN( u2_u9_u5_n174 ) );
  AOI21_X1 u2_u9_u5_U14 (.A( u2_u9_u5_n160 ) , .B2( u2_u9_u5_n161 ) , .ZN( u2_u9_u5_n162 ) , .B1( u2_u9_u5_n192 ) );
  INV_X1 u2_u9_u5_U15 (.A( u2_u9_u5_n159 ) , .ZN( u2_u9_u5_n192 ) );
  AOI21_X1 u2_u9_u5_U16 (.A( u2_u9_u5_n156 ) , .B2( u2_u9_u5_n157 ) , .B1( u2_u9_u5_n158 ) , .ZN( u2_u9_u5_n163 ) );
  AOI21_X1 u2_u9_u5_U17 (.B2( u2_u9_u5_n139 ) , .B1( u2_u9_u5_n140 ) , .ZN( u2_u9_u5_n141 ) , .A( u2_u9_u5_n150 ) );
  OAI21_X1 u2_u9_u5_U18 (.A( u2_u9_u5_n133 ) , .B2( u2_u9_u5_n134 ) , .B1( u2_u9_u5_n135 ) , .ZN( u2_u9_u5_n142 ) );
  OAI21_X1 u2_u9_u5_U19 (.ZN( u2_u9_u5_n133 ) , .B2( u2_u9_u5_n147 ) , .A( u2_u9_u5_n173 ) , .B1( u2_u9_u5_n188 ) );
  NAND2_X1 u2_u9_u5_U20 (.A2( u2_u9_u5_n119 ) , .A1( u2_u9_u5_n123 ) , .ZN( u2_u9_u5_n137 ) );
  INV_X1 u2_u9_u5_U21 (.A( u2_u9_u5_n155 ) , .ZN( u2_u9_u5_n194 ) );
  NAND2_X1 u2_u9_u5_U22 (.A1( u2_u9_u5_n121 ) , .ZN( u2_u9_u5_n132 ) , .A2( u2_u9_u5_n172 ) );
  NAND2_X1 u2_u9_u5_U23 (.A2( u2_u9_u5_n122 ) , .ZN( u2_u9_u5_n136 ) , .A1( u2_u9_u5_n154 ) );
  NAND2_X1 u2_u9_u5_U24 (.A2( u2_u9_u5_n119 ) , .A1( u2_u9_u5_n120 ) , .ZN( u2_u9_u5_n159 ) );
  INV_X1 u2_u9_u5_U25 (.A( u2_u9_u5_n156 ) , .ZN( u2_u9_u5_n175 ) );
  INV_X1 u2_u9_u5_U26 (.A( u2_u9_u5_n158 ) , .ZN( u2_u9_u5_n188 ) );
  INV_X1 u2_u9_u5_U27 (.A( u2_u9_u5_n152 ) , .ZN( u2_u9_u5_n179 ) );
  INV_X1 u2_u9_u5_U28 (.A( u2_u9_u5_n140 ) , .ZN( u2_u9_u5_n182 ) );
  INV_X1 u2_u9_u5_U29 (.A( u2_u9_u5_n151 ) , .ZN( u2_u9_u5_n183 ) );
  NOR2_X1 u2_u9_u5_U3 (.ZN( u2_u9_u5_n134 ) , .A1( u2_u9_u5_n183 ) , .A2( u2_u9_u5_n190 ) );
  INV_X1 u2_u9_u5_U30 (.A( u2_u9_u5_n123 ) , .ZN( u2_u9_u5_n185 ) );
  INV_X1 u2_u9_u5_U31 (.A( u2_u9_u5_n161 ) , .ZN( u2_u9_u5_n184 ) );
  INV_X1 u2_u9_u5_U32 (.A( u2_u9_u5_n139 ) , .ZN( u2_u9_u5_n189 ) );
  INV_X1 u2_u9_u5_U33 (.A( u2_u9_u5_n157 ) , .ZN( u2_u9_u5_n190 ) );
  INV_X1 u2_u9_u5_U34 (.A( u2_u9_u5_n120 ) , .ZN( u2_u9_u5_n193 ) );
  NAND2_X1 u2_u9_u5_U35 (.ZN( u2_u9_u5_n111 ) , .A1( u2_u9_u5_n140 ) , .A2( u2_u9_u5_n155 ) );
  NOR2_X1 u2_u9_u5_U36 (.ZN( u2_u9_u5_n100 ) , .A1( u2_u9_u5_n170 ) , .A2( u2_u9_u5_n180 ) );
  INV_X1 u2_u9_u5_U37 (.A( u2_u9_u5_n117 ) , .ZN( u2_u9_u5_n196 ) );
  OAI221_X1 u2_u9_u5_U38 (.A( u2_u9_u5_n116 ) , .ZN( u2_u9_u5_n117 ) , .B2( u2_u9_u5_n119 ) , .C1( u2_u9_u5_n153 ) , .C2( u2_u9_u5_n158 ) , .B1( u2_u9_u5_n172 ) );
  AOI222_X1 u2_u9_u5_U39 (.ZN( u2_u9_u5_n116 ) , .B2( u2_u9_u5_n145 ) , .C1( u2_u9_u5_n148 ) , .A2( u2_u9_u5_n174 ) , .C2( u2_u9_u5_n177 ) , .B1( u2_u9_u5_n187 ) , .A1( u2_u9_u5_n193 ) );
  INV_X1 u2_u9_u5_U4 (.A( u2_u9_u5_n138 ) , .ZN( u2_u9_u5_n191 ) );
  INV_X1 u2_u9_u5_U40 (.A( u2_u9_u5_n115 ) , .ZN( u2_u9_u5_n187 ) );
  OAI221_X1 u2_u9_u5_U41 (.A( u2_u9_u5_n101 ) , .ZN( u2_u9_u5_n102 ) , .C2( u2_u9_u5_n115 ) , .C1( u2_u9_u5_n126 ) , .B1( u2_u9_u5_n134 ) , .B2( u2_u9_u5_n160 ) );
  OAI21_X1 u2_u9_u5_U42 (.ZN( u2_u9_u5_n101 ) , .B1( u2_u9_u5_n137 ) , .A( u2_u9_u5_n146 ) , .B2( u2_u9_u5_n147 ) );
  AOI22_X1 u2_u9_u5_U43 (.B2( u2_u9_u5_n131 ) , .A2( u2_u9_u5_n146 ) , .ZN( u2_u9_u5_n169 ) , .B1( u2_u9_u5_n174 ) , .A1( u2_u9_u5_n185 ) );
  NOR2_X1 u2_u9_u5_U44 (.A1( u2_u9_u5_n146 ) , .ZN( u2_u9_u5_n150 ) , .A2( u2_u9_u5_n173 ) );
  AOI21_X1 u2_u9_u5_U45 (.A( u2_u9_u5_n118 ) , .B2( u2_u9_u5_n145 ) , .ZN( u2_u9_u5_n168 ) , .B1( u2_u9_u5_n186 ) );
  INV_X1 u2_u9_u5_U46 (.A( u2_u9_u5_n122 ) , .ZN( u2_u9_u5_n186 ) );
  NOR2_X1 u2_u9_u5_U47 (.A1( u2_u9_u5_n146 ) , .ZN( u2_u9_u5_n152 ) , .A2( u2_u9_u5_n176 ) );
  NOR2_X1 u2_u9_u5_U48 (.A1( u2_u9_u5_n115 ) , .ZN( u2_u9_u5_n118 ) , .A2( u2_u9_u5_n153 ) );
  NOR2_X1 u2_u9_u5_U49 (.A2( u2_u9_u5_n145 ) , .ZN( u2_u9_u5_n156 ) , .A1( u2_u9_u5_n174 ) );
  OAI21_X1 u2_u9_u5_U5 (.B2( u2_u9_u5_n136 ) , .B1( u2_u9_u5_n137 ) , .ZN( u2_u9_u5_n138 ) , .A( u2_u9_u5_n177 ) );
  NOR2_X1 u2_u9_u5_U50 (.ZN( u2_u9_u5_n121 ) , .A2( u2_u9_u5_n145 ) , .A1( u2_u9_u5_n176 ) );
  AOI22_X1 u2_u9_u5_U51 (.ZN( u2_u9_u5_n114 ) , .A2( u2_u9_u5_n137 ) , .A1( u2_u9_u5_n145 ) , .B2( u2_u9_u5_n175 ) , .B1( u2_u9_u5_n193 ) );
  OAI211_X1 u2_u9_u5_U52 (.B( u2_u9_u5_n124 ) , .A( u2_u9_u5_n125 ) , .C2( u2_u9_u5_n126 ) , .C1( u2_u9_u5_n127 ) , .ZN( u2_u9_u5_n128 ) );
  NOR3_X1 u2_u9_u5_U53 (.ZN( u2_u9_u5_n127 ) , .A1( u2_u9_u5_n136 ) , .A3( u2_u9_u5_n148 ) , .A2( u2_u9_u5_n182 ) );
  OAI21_X1 u2_u9_u5_U54 (.ZN( u2_u9_u5_n124 ) , .A( u2_u9_u5_n177 ) , .B2( u2_u9_u5_n183 ) , .B1( u2_u9_u5_n189 ) );
  OAI21_X1 u2_u9_u5_U55 (.ZN( u2_u9_u5_n125 ) , .A( u2_u9_u5_n174 ) , .B2( u2_u9_u5_n185 ) , .B1( u2_u9_u5_n190 ) );
  AOI21_X1 u2_u9_u5_U56 (.A( u2_u9_u5_n153 ) , .B2( u2_u9_u5_n154 ) , .B1( u2_u9_u5_n155 ) , .ZN( u2_u9_u5_n164 ) );
  AOI21_X1 u2_u9_u5_U57 (.ZN( u2_u9_u5_n110 ) , .B1( u2_u9_u5_n122 ) , .B2( u2_u9_u5_n139 ) , .A( u2_u9_u5_n153 ) );
  INV_X1 u2_u9_u5_U58 (.A( u2_u9_u5_n153 ) , .ZN( u2_u9_u5_n176 ) );
  INV_X1 u2_u9_u5_U59 (.A( u2_u9_u5_n126 ) , .ZN( u2_u9_u5_n173 ) );
  AOI222_X1 u2_u9_u5_U6 (.ZN( u2_u9_u5_n113 ) , .A1( u2_u9_u5_n131 ) , .C1( u2_u9_u5_n148 ) , .B2( u2_u9_u5_n174 ) , .C2( u2_u9_u5_n178 ) , .A2( u2_u9_u5_n179 ) , .B1( u2_u9_u5_n99 ) );
  AND2_X1 u2_u9_u5_U60 (.A2( u2_u9_u5_n104 ) , .A1( u2_u9_u5_n107 ) , .ZN( u2_u9_u5_n147 ) );
  AND2_X1 u2_u9_u5_U61 (.A2( u2_u9_u5_n104 ) , .A1( u2_u9_u5_n108 ) , .ZN( u2_u9_u5_n148 ) );
  NAND2_X1 u2_u9_u5_U62 (.A1( u2_u9_u5_n105 ) , .A2( u2_u9_u5_n106 ) , .ZN( u2_u9_u5_n158 ) );
  NAND2_X1 u2_u9_u5_U63 (.A2( u2_u9_u5_n108 ) , .A1( u2_u9_u5_n109 ) , .ZN( u2_u9_u5_n139 ) );
  NAND2_X1 u2_u9_u5_U64 (.A1( u2_u9_u5_n106 ) , .A2( u2_u9_u5_n108 ) , .ZN( u2_u9_u5_n119 ) );
  NAND2_X1 u2_u9_u5_U65 (.A2( u2_u9_u5_n103 ) , .A1( u2_u9_u5_n105 ) , .ZN( u2_u9_u5_n140 ) );
  NAND2_X1 u2_u9_u5_U66 (.A2( u2_u9_u5_n104 ) , .A1( u2_u9_u5_n105 ) , .ZN( u2_u9_u5_n155 ) );
  NAND2_X1 u2_u9_u5_U67 (.A2( u2_u9_u5_n106 ) , .A1( u2_u9_u5_n107 ) , .ZN( u2_u9_u5_n122 ) );
  NAND2_X1 u2_u9_u5_U68 (.A2( u2_u9_u5_n100 ) , .A1( u2_u9_u5_n106 ) , .ZN( u2_u9_u5_n115 ) );
  NAND2_X1 u2_u9_u5_U69 (.A2( u2_u9_u5_n100 ) , .A1( u2_u9_u5_n103 ) , .ZN( u2_u9_u5_n161 ) );
  INV_X1 u2_u9_u5_U7 (.A( u2_u9_u5_n135 ) , .ZN( u2_u9_u5_n178 ) );
  NAND2_X1 u2_u9_u5_U70 (.A1( u2_u9_u5_n105 ) , .A2( u2_u9_u5_n109 ) , .ZN( u2_u9_u5_n154 ) );
  INV_X1 u2_u9_u5_U71 (.A( u2_u9_u5_n146 ) , .ZN( u2_u9_u5_n172 ) );
  NAND2_X1 u2_u9_u5_U72 (.A1( u2_u9_u5_n103 ) , .A2( u2_u9_u5_n108 ) , .ZN( u2_u9_u5_n123 ) );
  NAND2_X1 u2_u9_u5_U73 (.A2( u2_u9_u5_n103 ) , .A1( u2_u9_u5_n107 ) , .ZN( u2_u9_u5_n151 ) );
  NAND2_X1 u2_u9_u5_U74 (.A2( u2_u9_u5_n107 ) , .A1( u2_u9_u5_n109 ) , .ZN( u2_u9_u5_n120 ) );
  NAND2_X1 u2_u9_u5_U75 (.A2( u2_u9_u5_n100 ) , .A1( u2_u9_u5_n109 ) , .ZN( u2_u9_u5_n157 ) );
  AND2_X1 u2_u9_u5_U76 (.A2( u2_u9_u5_n100 ) , .A1( u2_u9_u5_n104 ) , .ZN( u2_u9_u5_n131 ) );
  NOR2_X1 u2_u9_u5_U77 (.A2( u2_u9_X_34 ) , .A1( u2_u9_X_35 ) , .ZN( u2_u9_u5_n145 ) );
  NOR2_X1 u2_u9_u5_U78 (.A2( u2_u9_X_34 ) , .ZN( u2_u9_u5_n146 ) , .A1( u2_u9_u5_n171 ) );
  NOR2_X1 u2_u9_u5_U79 (.A2( u2_u9_X_31 ) , .A1( u2_u9_X_32 ) , .ZN( u2_u9_u5_n103 ) );
  OAI22_X1 u2_u9_u5_U8 (.B2( u2_u9_u5_n149 ) , .B1( u2_u9_u5_n150 ) , .A2( u2_u9_u5_n151 ) , .A1( u2_u9_u5_n152 ) , .ZN( u2_u9_u5_n165 ) );
  NOR2_X1 u2_u9_u5_U80 (.A2( u2_u9_X_36 ) , .ZN( u2_u9_u5_n105 ) , .A1( u2_u9_u5_n180 ) );
  NOR2_X1 u2_u9_u5_U81 (.A2( u2_u9_X_33 ) , .ZN( u2_u9_u5_n108 ) , .A1( u2_u9_u5_n170 ) );
  NOR2_X1 u2_u9_u5_U82 (.A2( u2_u9_X_33 ) , .A1( u2_u9_X_36 ) , .ZN( u2_u9_u5_n107 ) );
  NOR2_X1 u2_u9_u5_U83 (.A2( u2_u9_X_31 ) , .ZN( u2_u9_u5_n104 ) , .A1( u2_u9_u5_n181 ) );
  NAND2_X1 u2_u9_u5_U84 (.A2( u2_u9_X_34 ) , .A1( u2_u9_X_35 ) , .ZN( u2_u9_u5_n153 ) );
  NAND2_X1 u2_u9_u5_U85 (.A1( u2_u9_X_34 ) , .ZN( u2_u9_u5_n126 ) , .A2( u2_u9_u5_n171 ) );
  AND2_X1 u2_u9_u5_U86 (.A1( u2_u9_X_31 ) , .A2( u2_u9_X_32 ) , .ZN( u2_u9_u5_n106 ) );
  AND2_X1 u2_u9_u5_U87 (.A1( u2_u9_X_31 ) , .ZN( u2_u9_u5_n109 ) , .A2( u2_u9_u5_n181 ) );
  INV_X1 u2_u9_u5_U88 (.A( u2_u9_X_33 ) , .ZN( u2_u9_u5_n180 ) );
  INV_X1 u2_u9_u5_U89 (.A( u2_u9_X_35 ) , .ZN( u2_u9_u5_n171 ) );
  NOR3_X1 u2_u9_u5_U9 (.A2( u2_u9_u5_n147 ) , .A1( u2_u9_u5_n148 ) , .ZN( u2_u9_u5_n149 ) , .A3( u2_u9_u5_n194 ) );
  INV_X1 u2_u9_u5_U90 (.A( u2_u9_X_36 ) , .ZN( u2_u9_u5_n170 ) );
  INV_X1 u2_u9_u5_U91 (.A( u2_u9_X_32 ) , .ZN( u2_u9_u5_n181 ) );
  NAND4_X1 u2_u9_u5_U92 (.ZN( u2_out9_29 ) , .A4( u2_u9_u5_n129 ) , .A3( u2_u9_u5_n130 ) , .A2( u2_u9_u5_n168 ) , .A1( u2_u9_u5_n196 ) );
  AOI221_X1 u2_u9_u5_U93 (.A( u2_u9_u5_n128 ) , .ZN( u2_u9_u5_n129 ) , .C2( u2_u9_u5_n132 ) , .B2( u2_u9_u5_n159 ) , .B1( u2_u9_u5_n176 ) , .C1( u2_u9_u5_n184 ) );
  AOI222_X1 u2_u9_u5_U94 (.ZN( u2_u9_u5_n130 ) , .A2( u2_u9_u5_n146 ) , .B1( u2_u9_u5_n147 ) , .C2( u2_u9_u5_n175 ) , .B2( u2_u9_u5_n179 ) , .A1( u2_u9_u5_n188 ) , .C1( u2_u9_u5_n194 ) );
  NAND4_X1 u2_u9_u5_U95 (.ZN( u2_out9_19 ) , .A4( u2_u9_u5_n166 ) , .A3( u2_u9_u5_n167 ) , .A2( u2_u9_u5_n168 ) , .A1( u2_u9_u5_n169 ) );
  AOI22_X1 u2_u9_u5_U96 (.B2( u2_u9_u5_n145 ) , .A2( u2_u9_u5_n146 ) , .ZN( u2_u9_u5_n167 ) , .B1( u2_u9_u5_n182 ) , .A1( u2_u9_u5_n189 ) );
  NOR4_X1 u2_u9_u5_U97 (.A4( u2_u9_u5_n162 ) , .A3( u2_u9_u5_n163 ) , .A2( u2_u9_u5_n164 ) , .A1( u2_u9_u5_n165 ) , .ZN( u2_u9_u5_n166 ) );
  NAND4_X1 u2_u9_u5_U98 (.ZN( u2_out9_11 ) , .A4( u2_u9_u5_n143 ) , .A3( u2_u9_u5_n144 ) , .A2( u2_u9_u5_n169 ) , .A1( u2_u9_u5_n196 ) );
  AOI22_X1 u2_u9_u5_U99 (.A2( u2_u9_u5_n132 ) , .ZN( u2_u9_u5_n144 ) , .B2( u2_u9_u5_n145 ) , .B1( u2_u9_u5_n184 ) , .A1( u2_u9_u5_n194 ) );
  AOI22_X1 u2_u9_u6_U10 (.A2( u2_u9_u6_n151 ) , .B2( u2_u9_u6_n161 ) , .A1( u2_u9_u6_n167 ) , .B1( u2_u9_u6_n170 ) , .ZN( u2_u9_u6_n89 ) );
  AOI21_X1 u2_u9_u6_U11 (.B1( u2_u9_u6_n107 ) , .B2( u2_u9_u6_n132 ) , .A( u2_u9_u6_n158 ) , .ZN( u2_u9_u6_n88 ) );
  AOI21_X1 u2_u9_u6_U12 (.B2( u2_u9_u6_n147 ) , .B1( u2_u9_u6_n148 ) , .ZN( u2_u9_u6_n149 ) , .A( u2_u9_u6_n158 ) );
  AOI21_X1 u2_u9_u6_U13 (.ZN( u2_u9_u6_n106 ) , .A( u2_u9_u6_n142 ) , .B2( u2_u9_u6_n159 ) , .B1( u2_u9_u6_n164 ) );
  INV_X1 u2_u9_u6_U14 (.A( u2_u9_u6_n155 ) , .ZN( u2_u9_u6_n161 ) );
  INV_X1 u2_u9_u6_U15 (.A( u2_u9_u6_n128 ) , .ZN( u2_u9_u6_n164 ) );
  NAND2_X1 u2_u9_u6_U16 (.ZN( u2_u9_u6_n110 ) , .A1( u2_u9_u6_n122 ) , .A2( u2_u9_u6_n129 ) );
  NAND2_X1 u2_u9_u6_U17 (.ZN( u2_u9_u6_n124 ) , .A2( u2_u9_u6_n146 ) , .A1( u2_u9_u6_n148 ) );
  INV_X1 u2_u9_u6_U18 (.A( u2_u9_u6_n132 ) , .ZN( u2_u9_u6_n171 ) );
  AND2_X1 u2_u9_u6_U19 (.A1( u2_u9_u6_n100 ) , .ZN( u2_u9_u6_n130 ) , .A2( u2_u9_u6_n147 ) );
  INV_X1 u2_u9_u6_U20 (.A( u2_u9_u6_n127 ) , .ZN( u2_u9_u6_n173 ) );
  INV_X1 u2_u9_u6_U21 (.A( u2_u9_u6_n121 ) , .ZN( u2_u9_u6_n167 ) );
  INV_X1 u2_u9_u6_U22 (.A( u2_u9_u6_n100 ) , .ZN( u2_u9_u6_n169 ) );
  INV_X1 u2_u9_u6_U23 (.A( u2_u9_u6_n123 ) , .ZN( u2_u9_u6_n170 ) );
  INV_X1 u2_u9_u6_U24 (.A( u2_u9_u6_n113 ) , .ZN( u2_u9_u6_n168 ) );
  AND2_X1 u2_u9_u6_U25 (.A1( u2_u9_u6_n107 ) , .A2( u2_u9_u6_n119 ) , .ZN( u2_u9_u6_n133 ) );
  AND2_X1 u2_u9_u6_U26 (.A2( u2_u9_u6_n121 ) , .A1( u2_u9_u6_n122 ) , .ZN( u2_u9_u6_n131 ) );
  AND3_X1 u2_u9_u6_U27 (.ZN( u2_u9_u6_n120 ) , .A2( u2_u9_u6_n127 ) , .A1( u2_u9_u6_n132 ) , .A3( u2_u9_u6_n145 ) );
  INV_X1 u2_u9_u6_U28 (.A( u2_u9_u6_n146 ) , .ZN( u2_u9_u6_n163 ) );
  AOI222_X1 u2_u9_u6_U29 (.ZN( u2_u9_u6_n114 ) , .A1( u2_u9_u6_n118 ) , .A2( u2_u9_u6_n126 ) , .B2( u2_u9_u6_n151 ) , .C2( u2_u9_u6_n159 ) , .C1( u2_u9_u6_n168 ) , .B1( u2_u9_u6_n169 ) );
  INV_X1 u2_u9_u6_U3 (.A( u2_u9_u6_n110 ) , .ZN( u2_u9_u6_n166 ) );
  NOR2_X1 u2_u9_u6_U30 (.A1( u2_u9_u6_n162 ) , .A2( u2_u9_u6_n165 ) , .ZN( u2_u9_u6_n98 ) );
  NAND2_X1 u2_u9_u6_U31 (.A1( u2_u9_u6_n144 ) , .ZN( u2_u9_u6_n151 ) , .A2( u2_u9_u6_n158 ) );
  NAND2_X1 u2_u9_u6_U32 (.ZN( u2_u9_u6_n132 ) , .A1( u2_u9_u6_n91 ) , .A2( u2_u9_u6_n97 ) );
  AOI22_X1 u2_u9_u6_U33 (.B2( u2_u9_u6_n110 ) , .B1( u2_u9_u6_n111 ) , .A1( u2_u9_u6_n112 ) , .ZN( u2_u9_u6_n115 ) , .A2( u2_u9_u6_n161 ) );
  NAND4_X1 u2_u9_u6_U34 (.A3( u2_u9_u6_n109 ) , .ZN( u2_u9_u6_n112 ) , .A4( u2_u9_u6_n132 ) , .A2( u2_u9_u6_n147 ) , .A1( u2_u9_u6_n166 ) );
  NOR2_X1 u2_u9_u6_U35 (.ZN( u2_u9_u6_n109 ) , .A1( u2_u9_u6_n170 ) , .A2( u2_u9_u6_n173 ) );
  NOR2_X1 u2_u9_u6_U36 (.A2( u2_u9_u6_n126 ) , .ZN( u2_u9_u6_n155 ) , .A1( u2_u9_u6_n160 ) );
  NAND2_X1 u2_u9_u6_U37 (.ZN( u2_u9_u6_n146 ) , .A2( u2_u9_u6_n94 ) , .A1( u2_u9_u6_n99 ) );
  AOI21_X1 u2_u9_u6_U38 (.A( u2_u9_u6_n144 ) , .B2( u2_u9_u6_n145 ) , .B1( u2_u9_u6_n146 ) , .ZN( u2_u9_u6_n150 ) );
  AOI211_X1 u2_u9_u6_U39 (.B( u2_u9_u6_n134 ) , .A( u2_u9_u6_n135 ) , .C1( u2_u9_u6_n136 ) , .ZN( u2_u9_u6_n137 ) , .C2( u2_u9_u6_n151 ) );
  INV_X1 u2_u9_u6_U4 (.A( u2_u9_u6_n142 ) , .ZN( u2_u9_u6_n174 ) );
  NAND4_X1 u2_u9_u6_U40 (.A4( u2_u9_u6_n127 ) , .A3( u2_u9_u6_n128 ) , .A2( u2_u9_u6_n129 ) , .A1( u2_u9_u6_n130 ) , .ZN( u2_u9_u6_n136 ) );
  AOI21_X1 u2_u9_u6_U41 (.B2( u2_u9_u6_n132 ) , .B1( u2_u9_u6_n133 ) , .ZN( u2_u9_u6_n134 ) , .A( u2_u9_u6_n158 ) );
  AOI21_X1 u2_u9_u6_U42 (.B1( u2_u9_u6_n131 ) , .ZN( u2_u9_u6_n135 ) , .A( u2_u9_u6_n144 ) , .B2( u2_u9_u6_n146 ) );
  INV_X1 u2_u9_u6_U43 (.A( u2_u9_u6_n111 ) , .ZN( u2_u9_u6_n158 ) );
  NAND2_X1 u2_u9_u6_U44 (.ZN( u2_u9_u6_n127 ) , .A1( u2_u9_u6_n91 ) , .A2( u2_u9_u6_n92 ) );
  NAND2_X1 u2_u9_u6_U45 (.ZN( u2_u9_u6_n129 ) , .A2( u2_u9_u6_n95 ) , .A1( u2_u9_u6_n96 ) );
  INV_X1 u2_u9_u6_U46 (.A( u2_u9_u6_n144 ) , .ZN( u2_u9_u6_n159 ) );
  NAND2_X1 u2_u9_u6_U47 (.ZN( u2_u9_u6_n145 ) , .A2( u2_u9_u6_n97 ) , .A1( u2_u9_u6_n98 ) );
  NAND2_X1 u2_u9_u6_U48 (.ZN( u2_u9_u6_n148 ) , .A2( u2_u9_u6_n92 ) , .A1( u2_u9_u6_n94 ) );
  NAND2_X1 u2_u9_u6_U49 (.ZN( u2_u9_u6_n108 ) , .A2( u2_u9_u6_n139 ) , .A1( u2_u9_u6_n144 ) );
  NAND2_X1 u2_u9_u6_U5 (.A2( u2_u9_u6_n143 ) , .ZN( u2_u9_u6_n152 ) , .A1( u2_u9_u6_n166 ) );
  NAND2_X1 u2_u9_u6_U50 (.ZN( u2_u9_u6_n121 ) , .A2( u2_u9_u6_n95 ) , .A1( u2_u9_u6_n97 ) );
  NAND2_X1 u2_u9_u6_U51 (.ZN( u2_u9_u6_n107 ) , .A2( u2_u9_u6_n92 ) , .A1( u2_u9_u6_n95 ) );
  AND2_X1 u2_u9_u6_U52 (.ZN( u2_u9_u6_n118 ) , .A2( u2_u9_u6_n91 ) , .A1( u2_u9_u6_n99 ) );
  NAND2_X1 u2_u9_u6_U53 (.ZN( u2_u9_u6_n147 ) , .A2( u2_u9_u6_n98 ) , .A1( u2_u9_u6_n99 ) );
  NAND2_X1 u2_u9_u6_U54 (.ZN( u2_u9_u6_n128 ) , .A1( u2_u9_u6_n94 ) , .A2( u2_u9_u6_n96 ) );
  NAND2_X1 u2_u9_u6_U55 (.ZN( u2_u9_u6_n119 ) , .A2( u2_u9_u6_n95 ) , .A1( u2_u9_u6_n99 ) );
  NAND2_X1 u2_u9_u6_U56 (.ZN( u2_u9_u6_n123 ) , .A2( u2_u9_u6_n91 ) , .A1( u2_u9_u6_n96 ) );
  NAND2_X1 u2_u9_u6_U57 (.ZN( u2_u9_u6_n100 ) , .A2( u2_u9_u6_n92 ) , .A1( u2_u9_u6_n98 ) );
  NAND2_X1 u2_u9_u6_U58 (.ZN( u2_u9_u6_n122 ) , .A1( u2_u9_u6_n94 ) , .A2( u2_u9_u6_n97 ) );
  INV_X1 u2_u9_u6_U59 (.A( u2_u9_u6_n139 ) , .ZN( u2_u9_u6_n160 ) );
  AOI22_X1 u2_u9_u6_U6 (.B2( u2_u9_u6_n101 ) , .A1( u2_u9_u6_n102 ) , .ZN( u2_u9_u6_n103 ) , .B1( u2_u9_u6_n160 ) , .A2( u2_u9_u6_n161 ) );
  NAND2_X1 u2_u9_u6_U60 (.ZN( u2_u9_u6_n113 ) , .A1( u2_u9_u6_n96 ) , .A2( u2_u9_u6_n98 ) );
  NOR2_X1 u2_u9_u6_U61 (.A2( u2_u9_X_40 ) , .A1( u2_u9_X_41 ) , .ZN( u2_u9_u6_n126 ) );
  NOR2_X1 u2_u9_u6_U62 (.A2( u2_u9_X_39 ) , .A1( u2_u9_X_42 ) , .ZN( u2_u9_u6_n92 ) );
  NOR2_X1 u2_u9_u6_U63 (.A2( u2_u9_X_39 ) , .A1( u2_u9_u6_n156 ) , .ZN( u2_u9_u6_n97 ) );
  NOR2_X1 u2_u9_u6_U64 (.A2( u2_u9_X_38 ) , .A1( u2_u9_u6_n165 ) , .ZN( u2_u9_u6_n95 ) );
  NOR2_X1 u2_u9_u6_U65 (.A2( u2_u9_X_41 ) , .ZN( u2_u9_u6_n111 ) , .A1( u2_u9_u6_n157 ) );
  NOR2_X1 u2_u9_u6_U66 (.A2( u2_u9_X_37 ) , .A1( u2_u9_u6_n162 ) , .ZN( u2_u9_u6_n94 ) );
  NOR2_X1 u2_u9_u6_U67 (.A2( u2_u9_X_37 ) , .A1( u2_u9_X_38 ) , .ZN( u2_u9_u6_n91 ) );
  NAND2_X1 u2_u9_u6_U68 (.A1( u2_u9_X_41 ) , .ZN( u2_u9_u6_n144 ) , .A2( u2_u9_u6_n157 ) );
  NAND2_X1 u2_u9_u6_U69 (.A2( u2_u9_X_40 ) , .A1( u2_u9_X_41 ) , .ZN( u2_u9_u6_n139 ) );
  NOR2_X1 u2_u9_u6_U7 (.A1( u2_u9_u6_n118 ) , .ZN( u2_u9_u6_n143 ) , .A2( u2_u9_u6_n168 ) );
  AND2_X1 u2_u9_u6_U70 (.A1( u2_u9_X_39 ) , .A2( u2_u9_u6_n156 ) , .ZN( u2_u9_u6_n96 ) );
  AND2_X1 u2_u9_u6_U71 (.A1( u2_u9_X_39 ) , .A2( u2_u9_X_42 ) , .ZN( u2_u9_u6_n99 ) );
  INV_X1 u2_u9_u6_U72 (.A( u2_u9_X_40 ) , .ZN( u2_u9_u6_n157 ) );
  INV_X1 u2_u9_u6_U73 (.A( u2_u9_X_37 ) , .ZN( u2_u9_u6_n165 ) );
  INV_X1 u2_u9_u6_U74 (.A( u2_u9_X_38 ) , .ZN( u2_u9_u6_n162 ) );
  INV_X1 u2_u9_u6_U75 (.A( u2_u9_X_42 ) , .ZN( u2_u9_u6_n156 ) );
  NAND4_X1 u2_u9_u6_U76 (.ZN( u2_out9_32 ) , .A4( u2_u9_u6_n103 ) , .A3( u2_u9_u6_n104 ) , .A2( u2_u9_u6_n105 ) , .A1( u2_u9_u6_n106 ) );
  AOI22_X1 u2_u9_u6_U77 (.ZN( u2_u9_u6_n105 ) , .A2( u2_u9_u6_n108 ) , .A1( u2_u9_u6_n118 ) , .B2( u2_u9_u6_n126 ) , .B1( u2_u9_u6_n171 ) );
  AOI22_X1 u2_u9_u6_U78 (.ZN( u2_u9_u6_n104 ) , .A1( u2_u9_u6_n111 ) , .B1( u2_u9_u6_n124 ) , .B2( u2_u9_u6_n151 ) , .A2( u2_u9_u6_n93 ) );
  NAND4_X1 u2_u9_u6_U79 (.ZN( u2_out9_12 ) , .A4( u2_u9_u6_n114 ) , .A3( u2_u9_u6_n115 ) , .A2( u2_u9_u6_n116 ) , .A1( u2_u9_u6_n117 ) );
  OAI21_X1 u2_u9_u6_U8 (.A( u2_u9_u6_n159 ) , .B1( u2_u9_u6_n169 ) , .B2( u2_u9_u6_n173 ) , .ZN( u2_u9_u6_n90 ) );
  OAI22_X1 u2_u9_u6_U80 (.B2( u2_u9_u6_n111 ) , .ZN( u2_u9_u6_n116 ) , .B1( u2_u9_u6_n126 ) , .A2( u2_u9_u6_n164 ) , .A1( u2_u9_u6_n167 ) );
  OAI21_X1 u2_u9_u6_U81 (.A( u2_u9_u6_n108 ) , .ZN( u2_u9_u6_n117 ) , .B2( u2_u9_u6_n141 ) , .B1( u2_u9_u6_n163 ) );
  OAI211_X1 u2_u9_u6_U82 (.ZN( u2_out9_7 ) , .B( u2_u9_u6_n153 ) , .C2( u2_u9_u6_n154 ) , .C1( u2_u9_u6_n155 ) , .A( u2_u9_u6_n174 ) );
  NOR3_X1 u2_u9_u6_U83 (.A1( u2_u9_u6_n141 ) , .ZN( u2_u9_u6_n154 ) , .A3( u2_u9_u6_n164 ) , .A2( u2_u9_u6_n171 ) );
  AOI211_X1 u2_u9_u6_U84 (.B( u2_u9_u6_n149 ) , .A( u2_u9_u6_n150 ) , .C2( u2_u9_u6_n151 ) , .C1( u2_u9_u6_n152 ) , .ZN( u2_u9_u6_n153 ) );
  OAI211_X1 u2_u9_u6_U85 (.ZN( u2_out9_22 ) , .B( u2_u9_u6_n137 ) , .A( u2_u9_u6_n138 ) , .C2( u2_u9_u6_n139 ) , .C1( u2_u9_u6_n140 ) );
  AOI22_X1 u2_u9_u6_U86 (.B1( u2_u9_u6_n124 ) , .A2( u2_u9_u6_n125 ) , .A1( u2_u9_u6_n126 ) , .ZN( u2_u9_u6_n138 ) , .B2( u2_u9_u6_n161 ) );
  AND4_X1 u2_u9_u6_U87 (.A3( u2_u9_u6_n119 ) , .A1( u2_u9_u6_n120 ) , .A4( u2_u9_u6_n129 ) , .ZN( u2_u9_u6_n140 ) , .A2( u2_u9_u6_n143 ) );
  NAND3_X1 u2_u9_u6_U88 (.A2( u2_u9_u6_n123 ) , .ZN( u2_u9_u6_n125 ) , .A1( u2_u9_u6_n130 ) , .A3( u2_u9_u6_n131 ) );
  NAND3_X1 u2_u9_u6_U89 (.A3( u2_u9_u6_n133 ) , .ZN( u2_u9_u6_n141 ) , .A1( u2_u9_u6_n145 ) , .A2( u2_u9_u6_n148 ) );
  INV_X1 u2_u9_u6_U9 (.ZN( u2_u9_u6_n172 ) , .A( u2_u9_u6_n88 ) );
  NAND3_X1 u2_u9_u6_U90 (.ZN( u2_u9_u6_n101 ) , .A3( u2_u9_u6_n107 ) , .A2( u2_u9_u6_n121 ) , .A1( u2_u9_u6_n127 ) );
  NAND3_X1 u2_u9_u6_U91 (.ZN( u2_u9_u6_n102 ) , .A3( u2_u9_u6_n130 ) , .A2( u2_u9_u6_n145 ) , .A1( u2_u9_u6_n166 ) );
  NAND3_X1 u2_u9_u6_U92 (.A3( u2_u9_u6_n113 ) , .A1( u2_u9_u6_n119 ) , .A2( u2_u9_u6_n123 ) , .ZN( u2_u9_u6_n93 ) );
  NAND3_X1 u2_u9_u6_U93 (.ZN( u2_u9_u6_n142 ) , .A2( u2_u9_u6_n172 ) , .A3( u2_u9_u6_n89 ) , .A1( u2_u9_u6_n90 ) );
  AND3_X1 u2_u9_u7_U10 (.A3( u2_u9_u7_n110 ) , .A2( u2_u9_u7_n127 ) , .A1( u2_u9_u7_n132 ) , .ZN( u2_u9_u7_n92 ) );
  OAI21_X1 u2_u9_u7_U11 (.A( u2_u9_u7_n161 ) , .B1( u2_u9_u7_n168 ) , .B2( u2_u9_u7_n173 ) , .ZN( u2_u9_u7_n91 ) );
  AOI211_X1 u2_u9_u7_U12 (.A( u2_u9_u7_n117 ) , .ZN( u2_u9_u7_n118 ) , .C2( u2_u9_u7_n126 ) , .C1( u2_u9_u7_n177 ) , .B( u2_u9_u7_n180 ) );
  OAI22_X1 u2_u9_u7_U13 (.B1( u2_u9_u7_n115 ) , .ZN( u2_u9_u7_n117 ) , .A2( u2_u9_u7_n133 ) , .A1( u2_u9_u7_n137 ) , .B2( u2_u9_u7_n162 ) );
  INV_X1 u2_u9_u7_U14 (.A( u2_u9_u7_n116 ) , .ZN( u2_u9_u7_n180 ) );
  NOR3_X1 u2_u9_u7_U15 (.ZN( u2_u9_u7_n115 ) , .A3( u2_u9_u7_n145 ) , .A2( u2_u9_u7_n168 ) , .A1( u2_u9_u7_n169 ) );
  OAI211_X1 u2_u9_u7_U16 (.B( u2_u9_u7_n122 ) , .A( u2_u9_u7_n123 ) , .C2( u2_u9_u7_n124 ) , .ZN( u2_u9_u7_n154 ) , .C1( u2_u9_u7_n162 ) );
  AOI222_X1 u2_u9_u7_U17 (.ZN( u2_u9_u7_n122 ) , .C2( u2_u9_u7_n126 ) , .C1( u2_u9_u7_n145 ) , .B1( u2_u9_u7_n161 ) , .A2( u2_u9_u7_n165 ) , .B2( u2_u9_u7_n170 ) , .A1( u2_u9_u7_n176 ) );
  INV_X1 u2_u9_u7_U18 (.A( u2_u9_u7_n133 ) , .ZN( u2_u9_u7_n176 ) );
  NOR3_X1 u2_u9_u7_U19 (.A2( u2_u9_u7_n134 ) , .A1( u2_u9_u7_n135 ) , .ZN( u2_u9_u7_n136 ) , .A3( u2_u9_u7_n171 ) );
  NOR2_X1 u2_u9_u7_U20 (.A1( u2_u9_u7_n130 ) , .A2( u2_u9_u7_n134 ) , .ZN( u2_u9_u7_n153 ) );
  INV_X1 u2_u9_u7_U21 (.A( u2_u9_u7_n101 ) , .ZN( u2_u9_u7_n165 ) );
  NOR2_X1 u2_u9_u7_U22 (.ZN( u2_u9_u7_n111 ) , .A2( u2_u9_u7_n134 ) , .A1( u2_u9_u7_n169 ) );
  AOI21_X1 u2_u9_u7_U23 (.ZN( u2_u9_u7_n104 ) , .B2( u2_u9_u7_n112 ) , .B1( u2_u9_u7_n127 ) , .A( u2_u9_u7_n164 ) );
  AOI21_X1 u2_u9_u7_U24 (.ZN( u2_u9_u7_n106 ) , .B1( u2_u9_u7_n133 ) , .B2( u2_u9_u7_n146 ) , .A( u2_u9_u7_n162 ) );
  AOI21_X1 u2_u9_u7_U25 (.A( u2_u9_u7_n101 ) , .ZN( u2_u9_u7_n107 ) , .B2( u2_u9_u7_n128 ) , .B1( u2_u9_u7_n175 ) );
  INV_X1 u2_u9_u7_U26 (.A( u2_u9_u7_n138 ) , .ZN( u2_u9_u7_n171 ) );
  INV_X1 u2_u9_u7_U27 (.A( u2_u9_u7_n131 ) , .ZN( u2_u9_u7_n177 ) );
  INV_X1 u2_u9_u7_U28 (.A( u2_u9_u7_n110 ) , .ZN( u2_u9_u7_n174 ) );
  NAND2_X1 u2_u9_u7_U29 (.A1( u2_u9_u7_n129 ) , .A2( u2_u9_u7_n132 ) , .ZN( u2_u9_u7_n149 ) );
  OAI21_X1 u2_u9_u7_U3 (.ZN( u2_u9_u7_n159 ) , .A( u2_u9_u7_n165 ) , .B2( u2_u9_u7_n171 ) , .B1( u2_u9_u7_n174 ) );
  NAND2_X1 u2_u9_u7_U30 (.A1( u2_u9_u7_n113 ) , .A2( u2_u9_u7_n124 ) , .ZN( u2_u9_u7_n130 ) );
  INV_X1 u2_u9_u7_U31 (.A( u2_u9_u7_n112 ) , .ZN( u2_u9_u7_n173 ) );
  INV_X1 u2_u9_u7_U32 (.A( u2_u9_u7_n128 ) , .ZN( u2_u9_u7_n168 ) );
  INV_X1 u2_u9_u7_U33 (.A( u2_u9_u7_n148 ) , .ZN( u2_u9_u7_n169 ) );
  INV_X1 u2_u9_u7_U34 (.A( u2_u9_u7_n127 ) , .ZN( u2_u9_u7_n179 ) );
  NOR2_X1 u2_u9_u7_U35 (.ZN( u2_u9_u7_n101 ) , .A2( u2_u9_u7_n150 ) , .A1( u2_u9_u7_n156 ) );
  AOI211_X1 u2_u9_u7_U36 (.B( u2_u9_u7_n154 ) , .A( u2_u9_u7_n155 ) , .C1( u2_u9_u7_n156 ) , .ZN( u2_u9_u7_n157 ) , .C2( u2_u9_u7_n172 ) );
  INV_X1 u2_u9_u7_U37 (.A( u2_u9_u7_n153 ) , .ZN( u2_u9_u7_n172 ) );
  AOI211_X1 u2_u9_u7_U38 (.B( u2_u9_u7_n139 ) , .A( u2_u9_u7_n140 ) , .C2( u2_u9_u7_n141 ) , .ZN( u2_u9_u7_n142 ) , .C1( u2_u9_u7_n156 ) );
  NAND4_X1 u2_u9_u7_U39 (.A3( u2_u9_u7_n127 ) , .A2( u2_u9_u7_n128 ) , .A1( u2_u9_u7_n129 ) , .ZN( u2_u9_u7_n141 ) , .A4( u2_u9_u7_n147 ) );
  INV_X1 u2_u9_u7_U4 (.A( u2_u9_u7_n111 ) , .ZN( u2_u9_u7_n170 ) );
  AOI21_X1 u2_u9_u7_U40 (.A( u2_u9_u7_n137 ) , .B1( u2_u9_u7_n138 ) , .ZN( u2_u9_u7_n139 ) , .B2( u2_u9_u7_n146 ) );
  OAI22_X1 u2_u9_u7_U41 (.B1( u2_u9_u7_n136 ) , .ZN( u2_u9_u7_n140 ) , .A1( u2_u9_u7_n153 ) , .B2( u2_u9_u7_n162 ) , .A2( u2_u9_u7_n164 ) );
  AOI21_X1 u2_u9_u7_U42 (.ZN( u2_u9_u7_n123 ) , .B1( u2_u9_u7_n165 ) , .B2( u2_u9_u7_n177 ) , .A( u2_u9_u7_n97 ) );
  AOI21_X1 u2_u9_u7_U43 (.B2( u2_u9_u7_n113 ) , .B1( u2_u9_u7_n124 ) , .A( u2_u9_u7_n125 ) , .ZN( u2_u9_u7_n97 ) );
  INV_X1 u2_u9_u7_U44 (.A( u2_u9_u7_n125 ) , .ZN( u2_u9_u7_n161 ) );
  INV_X1 u2_u9_u7_U45 (.A( u2_u9_u7_n152 ) , .ZN( u2_u9_u7_n162 ) );
  AOI22_X1 u2_u9_u7_U46 (.A2( u2_u9_u7_n114 ) , .ZN( u2_u9_u7_n119 ) , .B1( u2_u9_u7_n130 ) , .A1( u2_u9_u7_n156 ) , .B2( u2_u9_u7_n165 ) );
  NAND2_X1 u2_u9_u7_U47 (.A2( u2_u9_u7_n112 ) , .ZN( u2_u9_u7_n114 ) , .A1( u2_u9_u7_n175 ) );
  AND2_X1 u2_u9_u7_U48 (.ZN( u2_u9_u7_n145 ) , .A2( u2_u9_u7_n98 ) , .A1( u2_u9_u7_n99 ) );
  NOR2_X1 u2_u9_u7_U49 (.ZN( u2_u9_u7_n137 ) , .A1( u2_u9_u7_n150 ) , .A2( u2_u9_u7_n161 ) );
  INV_X1 u2_u9_u7_U5 (.A( u2_u9_u7_n149 ) , .ZN( u2_u9_u7_n175 ) );
  AOI21_X1 u2_u9_u7_U50 (.ZN( u2_u9_u7_n105 ) , .B2( u2_u9_u7_n110 ) , .A( u2_u9_u7_n125 ) , .B1( u2_u9_u7_n147 ) );
  NAND2_X1 u2_u9_u7_U51 (.ZN( u2_u9_u7_n146 ) , .A1( u2_u9_u7_n95 ) , .A2( u2_u9_u7_n98 ) );
  NAND2_X1 u2_u9_u7_U52 (.A2( u2_u9_u7_n103 ) , .ZN( u2_u9_u7_n147 ) , .A1( u2_u9_u7_n93 ) );
  NAND2_X1 u2_u9_u7_U53 (.A1( u2_u9_u7_n103 ) , .ZN( u2_u9_u7_n127 ) , .A2( u2_u9_u7_n99 ) );
  OR2_X1 u2_u9_u7_U54 (.ZN( u2_u9_u7_n126 ) , .A2( u2_u9_u7_n152 ) , .A1( u2_u9_u7_n156 ) );
  NAND2_X1 u2_u9_u7_U55 (.A2( u2_u9_u7_n102 ) , .A1( u2_u9_u7_n103 ) , .ZN( u2_u9_u7_n133 ) );
  NAND2_X1 u2_u9_u7_U56 (.ZN( u2_u9_u7_n112 ) , .A2( u2_u9_u7_n96 ) , .A1( u2_u9_u7_n99 ) );
  NAND2_X1 u2_u9_u7_U57 (.A2( u2_u9_u7_n102 ) , .ZN( u2_u9_u7_n128 ) , .A1( u2_u9_u7_n98 ) );
  NAND2_X1 u2_u9_u7_U58 (.A1( u2_u9_u7_n100 ) , .ZN( u2_u9_u7_n113 ) , .A2( u2_u9_u7_n93 ) );
  NAND2_X1 u2_u9_u7_U59 (.A2( u2_u9_u7_n102 ) , .ZN( u2_u9_u7_n124 ) , .A1( u2_u9_u7_n96 ) );
  INV_X1 u2_u9_u7_U6 (.A( u2_u9_u7_n154 ) , .ZN( u2_u9_u7_n178 ) );
  NAND2_X1 u2_u9_u7_U60 (.ZN( u2_u9_u7_n110 ) , .A1( u2_u9_u7_n95 ) , .A2( u2_u9_u7_n96 ) );
  INV_X1 u2_u9_u7_U61 (.A( u2_u9_u7_n150 ) , .ZN( u2_u9_u7_n164 ) );
  AND2_X1 u2_u9_u7_U62 (.ZN( u2_u9_u7_n134 ) , .A1( u2_u9_u7_n93 ) , .A2( u2_u9_u7_n98 ) );
  NAND2_X1 u2_u9_u7_U63 (.A1( u2_u9_u7_n100 ) , .A2( u2_u9_u7_n102 ) , .ZN( u2_u9_u7_n129 ) );
  NAND2_X1 u2_u9_u7_U64 (.A2( u2_u9_u7_n103 ) , .ZN( u2_u9_u7_n131 ) , .A1( u2_u9_u7_n95 ) );
  NAND2_X1 u2_u9_u7_U65 (.A1( u2_u9_u7_n100 ) , .ZN( u2_u9_u7_n138 ) , .A2( u2_u9_u7_n99 ) );
  NAND2_X1 u2_u9_u7_U66 (.ZN( u2_u9_u7_n132 ) , .A1( u2_u9_u7_n93 ) , .A2( u2_u9_u7_n96 ) );
  NAND2_X1 u2_u9_u7_U67 (.A1( u2_u9_u7_n100 ) , .ZN( u2_u9_u7_n148 ) , .A2( u2_u9_u7_n95 ) );
  NOR2_X1 u2_u9_u7_U68 (.A2( u2_u9_X_47 ) , .ZN( u2_u9_u7_n150 ) , .A1( u2_u9_u7_n163 ) );
  NOR2_X1 u2_u9_u7_U69 (.A2( u2_u9_X_43 ) , .A1( u2_u9_X_44 ) , .ZN( u2_u9_u7_n103 ) );
  AOI211_X1 u2_u9_u7_U7 (.ZN( u2_u9_u7_n116 ) , .A( u2_u9_u7_n155 ) , .C1( u2_u9_u7_n161 ) , .C2( u2_u9_u7_n171 ) , .B( u2_u9_u7_n94 ) );
  NOR2_X1 u2_u9_u7_U70 (.A2( u2_u9_X_48 ) , .A1( u2_u9_u7_n166 ) , .ZN( u2_u9_u7_n95 ) );
  NOR2_X1 u2_u9_u7_U71 (.A2( u2_u9_X_45 ) , .A1( u2_u9_X_48 ) , .ZN( u2_u9_u7_n99 ) );
  NOR2_X1 u2_u9_u7_U72 (.A2( u2_u9_X_44 ) , .A1( u2_u9_u7_n167 ) , .ZN( u2_u9_u7_n98 ) );
  NOR2_X1 u2_u9_u7_U73 (.A2( u2_u9_X_46 ) , .A1( u2_u9_X_47 ) , .ZN( u2_u9_u7_n152 ) );
  AND2_X1 u2_u9_u7_U74 (.A1( u2_u9_X_47 ) , .ZN( u2_u9_u7_n156 ) , .A2( u2_u9_u7_n163 ) );
  NAND2_X1 u2_u9_u7_U75 (.A2( u2_u9_X_46 ) , .A1( u2_u9_X_47 ) , .ZN( u2_u9_u7_n125 ) );
  AND2_X1 u2_u9_u7_U76 (.A2( u2_u9_X_45 ) , .A1( u2_u9_X_48 ) , .ZN( u2_u9_u7_n102 ) );
  AND2_X1 u2_u9_u7_U77 (.A2( u2_u9_X_43 ) , .A1( u2_u9_X_44 ) , .ZN( u2_u9_u7_n96 ) );
  AND2_X1 u2_u9_u7_U78 (.A1( u2_u9_X_44 ) , .ZN( u2_u9_u7_n100 ) , .A2( u2_u9_u7_n167 ) );
  AND2_X1 u2_u9_u7_U79 (.A1( u2_u9_X_48 ) , .A2( u2_u9_u7_n166 ) , .ZN( u2_u9_u7_n93 ) );
  OAI222_X1 u2_u9_u7_U8 (.C2( u2_u9_u7_n101 ) , .B2( u2_u9_u7_n111 ) , .A1( u2_u9_u7_n113 ) , .C1( u2_u9_u7_n146 ) , .A2( u2_u9_u7_n162 ) , .B1( u2_u9_u7_n164 ) , .ZN( u2_u9_u7_n94 ) );
  INV_X1 u2_u9_u7_U80 (.A( u2_u9_X_46 ) , .ZN( u2_u9_u7_n163 ) );
  INV_X1 u2_u9_u7_U81 (.A( u2_u9_X_43 ) , .ZN( u2_u9_u7_n167 ) );
  INV_X1 u2_u9_u7_U82 (.A( u2_u9_X_45 ) , .ZN( u2_u9_u7_n166 ) );
  NAND4_X1 u2_u9_u7_U83 (.ZN( u2_out9_27 ) , .A4( u2_u9_u7_n118 ) , .A3( u2_u9_u7_n119 ) , .A2( u2_u9_u7_n120 ) , .A1( u2_u9_u7_n121 ) );
  OAI21_X1 u2_u9_u7_U84 (.ZN( u2_u9_u7_n121 ) , .B2( u2_u9_u7_n145 ) , .A( u2_u9_u7_n150 ) , .B1( u2_u9_u7_n174 ) );
  OAI21_X1 u2_u9_u7_U85 (.ZN( u2_u9_u7_n120 ) , .A( u2_u9_u7_n161 ) , .B2( u2_u9_u7_n170 ) , .B1( u2_u9_u7_n179 ) );
  NAND4_X1 u2_u9_u7_U86 (.ZN( u2_out9_21 ) , .A4( u2_u9_u7_n157 ) , .A3( u2_u9_u7_n158 ) , .A2( u2_u9_u7_n159 ) , .A1( u2_u9_u7_n160 ) );
  OAI21_X1 u2_u9_u7_U87 (.B1( u2_u9_u7_n145 ) , .ZN( u2_u9_u7_n160 ) , .A( u2_u9_u7_n161 ) , .B2( u2_u9_u7_n177 ) );
  AOI22_X1 u2_u9_u7_U88 (.B2( u2_u9_u7_n149 ) , .B1( u2_u9_u7_n150 ) , .A2( u2_u9_u7_n151 ) , .A1( u2_u9_u7_n152 ) , .ZN( u2_u9_u7_n158 ) );
  NAND4_X1 u2_u9_u7_U89 (.ZN( u2_out9_15 ) , .A4( u2_u9_u7_n142 ) , .A3( u2_u9_u7_n143 ) , .A2( u2_u9_u7_n144 ) , .A1( u2_u9_u7_n178 ) );
  OAI221_X1 u2_u9_u7_U9 (.C1( u2_u9_u7_n101 ) , .C2( u2_u9_u7_n147 ) , .ZN( u2_u9_u7_n155 ) , .B2( u2_u9_u7_n162 ) , .A( u2_u9_u7_n91 ) , .B1( u2_u9_u7_n92 ) );
  OR2_X1 u2_u9_u7_U90 (.A2( u2_u9_u7_n125 ) , .A1( u2_u9_u7_n129 ) , .ZN( u2_u9_u7_n144 ) );
  AOI22_X1 u2_u9_u7_U91 (.A2( u2_u9_u7_n126 ) , .ZN( u2_u9_u7_n143 ) , .B2( u2_u9_u7_n165 ) , .B1( u2_u9_u7_n173 ) , .A1( u2_u9_u7_n174 ) );
  NAND4_X1 u2_u9_u7_U92 (.ZN( u2_out9_5 ) , .A4( u2_u9_u7_n108 ) , .A3( u2_u9_u7_n109 ) , .A1( u2_u9_u7_n116 ) , .A2( u2_u9_u7_n123 ) );
  AOI22_X1 u2_u9_u7_U93 (.ZN( u2_u9_u7_n109 ) , .A2( u2_u9_u7_n126 ) , .B2( u2_u9_u7_n145 ) , .B1( u2_u9_u7_n156 ) , .A1( u2_u9_u7_n171 ) );
  NOR4_X1 u2_u9_u7_U94 (.A4( u2_u9_u7_n104 ) , .A3( u2_u9_u7_n105 ) , .A2( u2_u9_u7_n106 ) , .A1( u2_u9_u7_n107 ) , .ZN( u2_u9_u7_n108 ) );
  NAND3_X1 u2_u9_u7_U95 (.A3( u2_u9_u7_n146 ) , .A2( u2_u9_u7_n147 ) , .A1( u2_u9_u7_n148 ) , .ZN( u2_u9_u7_n151 ) );
  NAND3_X1 u2_u9_u7_U96 (.A3( u2_u9_u7_n131 ) , .A2( u2_u9_u7_n132 ) , .A1( u2_u9_u7_n133 ) , .ZN( u2_u9_u7_n135 ) );
  INV_X1 u2_uk_U10 (.A( u2_uk_n188 ) , .ZN( u2_uk_n27 ) );
  OAI21_X1 u2_uk_U1003 (.ZN( u2_K12_7 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1720 ) , .A( u2_uk_n520 ) );
  OAI21_X1 u2_uk_U1021 (.ZN( u2_K6_41 ) , .A( u2_uk_n1069 ) , .B1( u2_uk_n110 ) , .B2( u2_uk_n1445 ) );
  OAI21_X1 u2_uk_U1025 (.ZN( u2_K4_28 ) , .A( u2_uk_n1029 ) , .B2( u2_uk_n1351 ) , .B1( u2_uk_n17 ) );
  NAND2_X1 u2_uk_U1026 (.A1( u2_uk_K_r2_21 ) , .ZN( u2_uk_n1029 ) , .A2( u2_uk_n99 ) );
  OAI21_X1 u2_uk_U1031 (.ZN( u2_K15_14 ) , .B1( u2_uk_n109 ) , .B2( u2_uk_n1821 ) , .A( u2_uk_n936 ) );
  NAND2_X1 u2_uk_U1032 (.A1( u2_uk_K_r13_32 ) , .A2( u2_uk_n83 ) , .ZN( u2_uk_n936 ) );
  OAI21_X1 u2_uk_U1037 (.ZN( u2_K5_42 ) , .A( u2_uk_n1052 ) , .B2( u2_uk_n1382 ) , .B1( u2_uk_n17 ) );
  NAND2_X1 u2_uk_U1038 (.A1( u2_uk_K_r3_9 ) , .ZN( u2_uk_n1052 ) , .A2( u2_uk_n60 ) );
  INV_X1 u2_uk_U1044 (.A( u2_key_r_7 ) , .ZN( u2_uk_n1147 ) );
  INV_X1 u2_uk_U1047 (.A( u2_key_r_23 ) , .ZN( u2_uk_n1158 ) );
  INV_X1 u2_uk_U1049 (.A( u2_key_r_30 ) , .ZN( u2_uk_n1165 ) );
  OAI22_X1 u2_uk_U106 (.ZN( u2_K10_41 ) , .A2( u2_uk_n1594 ) , .B2( u2_uk_n1622 ) , .B1( u2_uk_n17 ) , .A1( u2_uk_n231 ) );
  OAI21_X1 u2_uk_U1072 (.ZN( u2_K3_40 ) , .A( u2_uk_n1014 ) , .B2( u2_uk_n1300 ) , .B1( u2_uk_n230 ) );
  NAND2_X1 u2_uk_U1073 (.A1( u2_uk_K_r1_21 ) , .ZN( u2_uk_n1014 ) , .A2( u2_uk_n148 ) );
  OAI22_X1 u2_uk_U109 (.ZN( u2_K3_41 ) , .A2( u2_uk_n1283 ) , .B2( u2_uk_n1288 ) , .B1( u2_uk_n141 ) , .A1( u2_uk_n83 ) );
  INV_X1 u2_uk_U1090 (.ZN( u2_K7_6 ) , .A( u2_uk_n1095 ) );
  AOI22_X1 u2_uk_U1091 (.B2( u2_uk_K_r5_39 ) , .A2( u2_uk_K_r5_4 ) , .ZN( u2_uk_n1095 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n182 ) );
  INV_X1 u2_uk_U1092 (.ZN( u2_K1_41 ) , .A( u2_uk_n985 ) );
  INV_X1 u2_uk_U11 (.A( u2_uk_n163 ) , .ZN( u2_uk_n60 ) );
  INV_X1 u2_uk_U1104 (.ZN( u2_K4_3 ) , .A( u2_uk_n1035 ) );
  INV_X1 u2_uk_U1106 (.ZN( u2_K12_23 ) , .A( u2_uk_n454 ) );
  INV_X1 u2_uk_U1110 (.ZN( u2_K12_32 ) , .A( u2_uk_n467 ) );
  INV_X1 u2_uk_U1112 (.ZN( u2_K9_20 ) , .A( u2_uk_n1126 ) );
  AOI22_X1 u2_uk_U1113 (.B2( u2_uk_K_r7_32 ) , .A2( u2_uk_K_r7_39 ) , .ZN( u2_uk_n1126 ) , .A1( u2_uk_n162 ) , .B1( u2_uk_n63 ) );
  INV_X1 u2_uk_U1114 (.ZN( u2_K5_20 ) , .A( u2_uk_n1043 ) );
  INV_X1 u2_uk_U1116 (.ZN( u2_K7_13 ) , .A( u2_uk_n1076 ) );
  INV_X1 u2_uk_U1120 (.ZN( u2_K7_32 ) , .A( u2_uk_n1088 ) );
  INV_X1 u2_uk_U1122 (.ZN( u2_K4_20 ) , .A( u2_uk_n1024 ) );
  INV_X1 u2_uk_U1124 (.ZN( u2_K4_4 ) , .A( u2_uk_n1037 ) );
  AOI22_X1 u2_uk_U1125 (.B2( u2_uk_K_r2_13 ) , .A2( u2_uk_K_r2_18 ) , .ZN( u2_uk_n1037 ) , .B1( u2_uk_n147 ) , .A1( u2_uk_n83 ) );
  INV_X1 u2_uk_U1126 (.ZN( u2_K5_35 ) , .A( u2_uk_n1049 ) );
  INV_X1 u2_uk_U113 (.ZN( u2_K11_47 ) , .A( u2_uk_n386 ) );
  INV_X1 u2_uk_U1130 (.ZN( u2_K4_10 ) , .A( u2_uk_n1020 ) );
  INV_X1 u2_uk_U1145 (.ZN( u2_K12_1 ) , .A( u2_uk_n421 ) );
  INV_X1 u2_uk_U1146 (.ZN( u2_K13_2 ) , .A( u2_uk_n665 ) );
  OAI22_X1 u2_uk_U115 (.ZN( u2_K10_47 ) , .A2( u2_uk_n1594 ) , .B2( u2_uk_n1609 ) , .B1( u2_uk_n164 ) , .A1( u2_uk_n93 ) );
  INV_X1 u2_uk_U1153 (.ZN( u2_K9_2 ) , .A( u2_uk_n1130 ) );
  AOI22_X1 u2_uk_U1154 (.B2( u2_uk_K_r4_17 ) , .A2( u2_uk_K_r4_55 ) , .ZN( u2_uk_n1066 ) , .B1( u2_uk_n148 ) , .A1( u2_uk_n63 ) );
  INV_X1 u2_uk_U1155 (.ZN( u2_K6_2 ) , .A( u2_uk_n1066 ) );
  INV_X1 u2_uk_U1157 (.ZN( u2_K4_2 ) , .A( u2_uk_n1031 ) );
  OAI22_X1 u2_uk_U117 (.ZN( u2_K7_47 ) , .A2( u2_uk_n1456 ) , .B2( u2_uk_n1470 ) , .A1( u2_uk_n164 ) , .B1( u2_uk_n31 ) );
  INV_X1 u2_uk_U12 (.A( u2_uk_n145 ) , .ZN( u2_uk_n83 ) );
  OAI22_X1 u2_uk_U121 (.ZN( u2_K4_47 ) , .B2( u2_uk_n1350 ) , .A2( u2_uk_n1359 ) , .A1( u2_uk_n187 ) , .B1( u2_uk_n63 ) );
  OAI22_X1 u2_uk_U125 (.ZN( u2_K4_15 ) , .B2( u2_uk_n1328 ) , .A2( u2_uk_n1356 ) , .A1( u2_uk_n182 ) , .B1( u2_uk_n63 ) );
  INV_X1 u2_uk_U13 (.A( u2_uk_n182 ) , .ZN( u2_uk_n92 ) );
  OAI22_X1 u2_uk_U130 (.ZN( u2_K7_15 ) , .A2( u2_uk_n1454 ) , .A1( u2_uk_n148 ) , .B2( u2_uk_n1494 ) , .B1( u2_uk_n31 ) );
  INV_X1 u2_uk_U14 (.A( u2_uk_n145 ) , .ZN( u2_uk_n94 ) );
  INV_X1 u2_uk_U149 (.ZN( u2_K11_19 ) , .A( u2_uk_n338 ) );
  INV_X1 u2_uk_U15 (.A( u2_uk_n164 ) , .ZN( u2_uk_n93 ) );
  AOI22_X1 u2_uk_U150 (.B2( u2_uk_K_r9_10 ) , .A2( u2_uk_K_r9_48 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n163 ) , .ZN( u2_uk_n338 ) );
  INV_X1 u2_uk_U151 (.ZN( u2_K9_19 ) , .A( u2_uk_n1124 ) );
  OAI22_X1 u2_uk_U153 (.ZN( u2_K7_19 ) , .B2( u2_uk_n1465 ) , .A2( u2_uk_n1475 ) , .A1( u2_uk_n209 ) , .B1( u2_uk_n31 ) );
  INV_X1 u2_uk_U16 (.A( u2_uk_n146 ) , .ZN( u2_uk_n99 ) );
  OAI22_X1 u2_uk_U163 (.ZN( u2_K14_30 ) , .B1( u2_uk_n142 ) , .B2( u2_uk_n1781 ) , .A2( u2_uk_n1808 ) , .A1( u2_uk_n94 ) );
  INV_X1 u2_uk_U164 (.ZN( u2_K12_30 ) , .A( u2_uk_n456 ) );
  INV_X1 u2_uk_U17 (.ZN( u2_uk_n109 ) , .A( u2_uk_n146 ) );
  OAI22_X1 u2_uk_U176 (.ZN( u2_K12_14 ) , .B2( u2_uk_n1688 ) , .A2( u2_uk_n1693 ) , .B1( u2_uk_n214 ) , .A1( u2_uk_n92 ) );
  INV_X1 u2_uk_U18 (.ZN( u2_uk_n110 ) , .A( u2_uk_n209 ) );
  INV_X1 u2_uk_U19 (.ZN( u2_uk_n100 ) , .A( u2_uk_n146 ) );
  OAI21_X1 u2_uk_U190 (.ZN( u2_K13_30 ) , .B1( u2_uk_n110 ) , .B2( u2_uk_n1746 ) , .A( u2_uk_n671 ) );
  NAND2_X1 u2_uk_U191 (.A1( u2_uk_K_r11_28 ) , .A2( u2_uk_n17 ) , .ZN( u2_uk_n671 ) );
  INV_X1 u2_uk_U194 (.ZN( u2_K7_24 ) , .A( u2_uk_n1083 ) );
  INV_X1 u2_uk_U197 (.ZN( u2_K3_24 ) , .A( u2_uk_n1008 ) );
  OAI22_X1 u2_uk_U199 (.ZN( u2_K15_24 ) , .A2( u2_uk_n1816 ) , .B2( u2_uk_n1834 ) , .B1( u2_uk_n222 ) , .A1( u2_uk_n93 ) );
  INV_X1 u2_uk_U20 (.ZN( u2_uk_n102 ) , .A( u2_uk_n146 ) );
  OAI21_X1 u2_uk_U204 (.ZN( u2_K4_30 ) , .A( u2_uk_n1032 ) , .B2( u2_uk_n1345 ) , .B1( u2_uk_n187 ) );
  NAND2_X1 u2_uk_U205 (.A1( u2_uk_K_r2_28 ) , .ZN( u2_uk_n1032 ) , .A2( u2_uk_n148 ) );
  OAI22_X1 u2_uk_U208 (.ZN( u2_K3_14 ) , .B1( u2_uk_n10 ) , .B2( u2_uk_n1310 ) , .A2( u2_uk_n1317 ) , .A1( u2_uk_n202 ) );
  INV_X1 u2_uk_U209 (.ZN( u2_K4_31 ) , .A( u2_uk_n1033 ) );
  INV_X1 u2_uk_U21 (.ZN( u2_uk_n128 ) , .A( u2_uk_n223 ) );
  AOI22_X1 u2_uk_U210 (.B2( u2_uk_K_r2_31 ) , .A2( u2_uk_K_r2_49 ) , .B1( u2_uk_n10 ) , .ZN( u2_uk_n1033 ) , .A1( u2_uk_n188 ) );
  OAI22_X1 u2_uk_U211 (.ZN( u2_K1_31 ) , .A2( u2_uk_n1147 ) , .B2( u2_uk_n1151 ) , .A1( u2_uk_n208 ) , .B1( u2_uk_n31 ) );
  INV_X1 u2_uk_U212 (.A( u2_key_r_14 ) , .ZN( u2_uk_n1151 ) );
  INV_X1 u2_uk_U217 (.ZN( u2_K11_31 ) , .A( u2_uk_n373 ) );
  BUF_X1 u2_uk_U22 (.Z( u2_uk_n141 ) , .A( u2_uk_n223 ) );
  INV_X1 u2_uk_U222 (.ZN( u2_K10_39 ) , .A( u2_uk_n305 ) );
  OAI21_X1 u2_uk_U225 (.ZN( u2_K10_31 ) , .B2( u2_uk_n1615 ) , .B1( u2_uk_n164 ) , .A( u2_uk_n291 ) );
  NAND2_X1 u2_uk_U226 (.A1( u2_uk_K_r8_16 ) , .A2( u2_uk_n155 ) , .ZN( u2_uk_n291 ) );
  BUF_X1 u2_uk_U23 (.Z( u2_uk_n155 ) , .A( u2_uk_n214 ) );
  OAI22_X1 u2_uk_U235 (.ZN( u2_K14_31 ) , .B1( u2_uk_n142 ) , .B2( u2_uk_n1797 ) , .A2( u2_uk_n1803 ) , .A1( u2_uk_n94 ) );
  BUF_X1 u2_uk_U24 (.Z( u2_uk_n145 ) , .A( u2_uk_n222 ) );
  BUF_X1 u2_uk_U25 (.Z( u2_uk_n142 ) , .A( u2_uk_n222 ) );
  OAI21_X1 u2_uk_U250 (.ZN( u2_K15_48 ) , .B1( u2_uk_n109 ) , .B2( u2_uk_n1824 ) , .A( u2_uk_n945 ) );
  INV_X1 u2_uk_U256 (.ZN( u2_K12_44 ) , .A( u2_uk_n504 ) );
  BUF_X1 u2_uk_U26 (.Z( u2_uk_n148 ) , .A( u2_uk_n217 ) );
  OAI22_X1 u2_uk_U267 (.ZN( u2_K7_44 ) , .A1( u2_uk_n118 ) , .B1( u2_uk_n142 ) , .B2( u2_uk_n1459 ) , .A2( u2_uk_n1480 ) );
  OAI22_X1 u2_uk_U269 (.ZN( u2_K6_44 ) , .B2( u2_uk_n1428 ) , .A2( u2_uk_n1446 ) , .B1( u2_uk_n182 ) , .A1( u2_uk_n93 ) );
  BUF_X1 u2_uk_U27 (.Z( u2_uk_n129 ) , .A( u2_uk_n220 ) );
  OAI22_X1 u2_uk_U270 (.ZN( u2_K6_48 ) , .B2( u2_uk_n1433 ) , .A2( u2_uk_n1440 ) , .A1( u2_uk_n222 ) , .B1( u2_uk_n60 ) );
  OAI21_X1 u2_uk_U272 (.ZN( u2_K3_44 ) , .A( u2_uk_n1015 ) , .B1( u2_uk_n109 ) , .B2( u2_uk_n1284 ) );
  NAND2_X1 u2_uk_U273 (.A1( u2_uk_K_r1_15 ) , .ZN( u2_uk_n1015 ) , .A2( u2_uk_n60 ) );
  OAI22_X1 u2_uk_U277 (.ZN( u2_K15_6 ) , .B1( u2_uk_n17 ) , .B2( u2_uk_n1834 ) , .A2( u2_uk_n1852 ) , .A1( u2_uk_n217 ) );
  BUF_X1 u2_uk_U28 (.Z( u2_uk_n146 ) , .A( u2_uk_n182 ) );
  OAI22_X1 u2_uk_U283 (.ZN( u2_K3_6 ) , .A2( u2_uk_n1282 ) , .B2( u2_uk_n1287 ) , .B1( u2_uk_n222 ) , .A1( u2_uk_n92 ) );
  INV_X1 u2_uk_U285 (.ZN( u2_K15_8 ) , .A( u2_uk_n946 ) );
  INV_X1 u2_uk_U289 (.ZN( u2_K7_8 ) , .A( u2_uk_n1096 ) );
  BUF_X1 u2_uk_U29 (.Z( u2_uk_n147 ) , .A( u2_uk_n217 ) );
  INV_X1 u2_uk_U292 (.ZN( u2_K4_8 ) , .A( u2_uk_n1040 ) );
  OAI22_X1 u2_uk_U294 (.ZN( u2_K3_8 ) , .A2( u2_uk_n1280 ) , .B2( u2_uk_n1296 ) , .A1( u2_uk_n164 ) , .B1( u2_uk_n94 ) );
  INV_X1 u2_uk_U3 (.ZN( u2_uk_n10 ) , .A( u2_uk_n141 ) );
  BUF_X1 u2_uk_U30 (.Z( u2_uk_n161 ) , .A( u2_uk_n213 ) );
  INV_X1 u2_uk_U301 (.ZN( u2_K9_26 ) , .A( u2_uk_n1128 ) );
  INV_X1 u2_uk_U303 (.ZN( u2_K4_26 ) , .A( u2_uk_n1028 ) );
  INV_X1 u2_uk_U305 (.ZN( u2_K15_26 ) , .A( u2_uk_n939 ) );
  OAI21_X1 u2_uk_U307 (.ZN( u2_K6_26 ) , .A( u2_uk_n1064 ) , .B2( u2_uk_n1439 ) , .B1( u2_uk_n188 ) );
  NAND2_X1 u2_uk_U308 (.A1( u2_uk_K_r4_35 ) , .ZN( u2_uk_n1064 ) , .A2( u2_uk_n191 ) );
  BUF_X1 u2_uk_U31 (.Z( u2_uk_n163 ) , .A( u2_uk_n209 ) );
  BUF_X1 u2_uk_U32 (.Z( u2_uk_n162 ) , .A( u2_uk_n223 ) );
  OAI21_X1 u2_uk_U326 (.ZN( u2_K3_46 ) , .A( u2_uk_n1017 ) , .B2( u2_uk_n1297 ) , .B1( u2_uk_n202 ) );
  NAND2_X1 u2_uk_U327 (.A1( u2_uk_K_r1_22 ) , .ZN( u2_uk_n1017 ) , .A2( u2_uk_n148 ) );
  BUF_X1 u2_uk_U33 (.Z( u2_uk_n182 ) , .A( u2_uk_n208 ) );
  INV_X1 u2_uk_U338 (.ZN( u2_K12_4 ) , .A( u2_uk_n515 ) );
  BUF_X1 u2_uk_U34 (.Z( u2_uk_n164 ) , .A( u2_uk_n208 ) );
  OAI22_X1 u2_uk_U342 (.ZN( u2_K3_4 ) , .B2( u2_uk_n1293 ) , .A2( u2_uk_n1301 ) , .A1( u2_uk_n213 ) , .B1( u2_uk_n93 ) );
  BUF_X1 u2_uk_U35 (.A( u2_uk_n164 ) , .Z( u2_uk_n187 ) );
  INV_X1 u2_uk_U350 (.ZN( u2_K10_40 ) , .A( u2_uk_n306 ) );
  AOI22_X1 u2_uk_U351 (.A2( u2_uk_K_r8_2 ) , .B2( u2_uk_K_r8_22 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n203 ) , .ZN( u2_uk_n306 ) );
  OAI22_X1 u2_uk_U355 (.ZN( u2_K15_40 ) , .A1( u2_uk_n162 ) , .B1( u2_uk_n17 ) , .A2( u2_uk_n1817 ) , .B2( u2_uk_n1849 ) );
  BUF_X1 u2_uk_U36 (.Z( u2_uk_n188 ) , .A( u2_uk_n209 ) );
  OAI21_X1 u2_uk_U362 (.ZN( u2_K15_33 ) , .B1( u2_uk_n109 ) , .B2( u2_uk_n1840 ) , .A( u2_uk_n942 ) );
  BUF_X1 u2_uk_U37 (.Z( u2_uk_n213 ) , .A( u2_uk_n231 ) );
  OAI21_X1 u2_uk_U374 (.ZN( u2_K5_33 ) , .A( u2_uk_n1048 ) , .B2( u2_uk_n1401 ) , .B1( u2_uk_n202 ) );
  NAND2_X1 u2_uk_U375 (.A1( u2_uk_K_r3_14 ) , .ZN( u2_uk_n1048 ) , .A2( u2_uk_n203 ) );
  BUF_X1 u2_uk_U38 (.Z( u2_uk_n208 ) , .A( u2_uk_n231 ) );
  OAI21_X1 u2_uk_U388 (.ZN( u2_K4_1 ) , .A( u2_uk_n1023 ) , .B2( u2_uk_n1323 ) , .B1( u2_uk_n208 ) );
  NAND2_X1 u2_uk_U389 (.A1( u2_uk_K_r2_25 ) , .ZN( u2_uk_n1023 ) , .A2( u2_uk_n214 ) );
  BUF_X1 u2_uk_U39 (.Z( u2_uk_n214 ) , .A( u2_uk_n231 ) );
  OAI22_X1 u2_uk_U390 (.ZN( u2_K3_1 ) , .B2( u2_uk_n1285 ) , .A1( u2_uk_n129 ) , .A2( u2_uk_n1290 ) , .B1( u2_uk_n27 ) );
  OAI21_X1 u2_uk_U392 (.ZN( u2_K7_1 ) , .A( u2_uk_n1078 ) , .B2( u2_uk_n1462 ) , .B1( u2_uk_n208 ) );
  NAND2_X1 u2_uk_U393 (.A1( u2_uk_K_r5_10 ) , .ZN( u2_uk_n1078 ) , .A2( u2_uk_n129 ) );
  OAI22_X1 u2_uk_U398 (.ZN( u2_K9_16 ) , .B2( u2_uk_n1548 ) , .A2( u2_uk_n1555 ) , .B1( u2_uk_n220 ) , .A1( u2_uk_n99 ) );
  INV_X1 u2_uk_U4 (.ZN( u2_uk_n118 ) , .A( u2_uk_n187 ) );
  BUF_X1 u2_uk_U40 (.Z( u2_uk_n209 ) , .A( u2_uk_n231 ) );
  OAI21_X1 u2_uk_U400 (.ZN( u2_K7_16 ) , .A( u2_uk_n1077 ) , .B1( u2_uk_n110 ) , .B2( u2_uk_n1496 ) );
  OAI22_X1 u2_uk_U403 (.ZN( u2_K4_16 ) , .B2( u2_uk_n1329 ) , .A2( u2_uk_n1333 ) , .A1( u2_uk_n207 ) , .B1( u2_uk_n99 ) );
  BUF_X1 u2_uk_U41 (.Z( u2_uk_n203 ) , .A( u2_uk_n222 ) );
  OAI22_X1 u2_uk_U415 (.ZN( u2_K4_9 ) , .A1( u2_uk_n118 ) , .B2( u2_uk_n1329 ) , .A2( u2_uk_n1339 ) , .B1( u2_uk_n238 ) );
  INV_X1 u2_uk_U416 (.ZN( u2_K10_37 ) , .A( u2_uk_n299 ) );
  BUF_X1 u2_uk_U42 (.A( u2_uk_n182 ) , .Z( u2_uk_n202 ) );
  INV_X1 u2_uk_U422 (.ZN( u2_K9_9 ) , .A( u2_uk_n1141 ) );
  INV_X1 u2_uk_U424 (.ZN( u2_K6_9 ) , .A( u2_uk_n1074 ) );
  OAI21_X1 u2_uk_U428 (.ZN( u2_K3_9 ) , .A( u2_uk_n1019 ) , .B2( u2_uk_n1295 ) , .B1( u2_uk_n202 ) );
  NAND2_X1 u2_uk_U429 (.A1( u2_uk_K_r1_18 ) , .ZN( u2_uk_n1019 ) , .A2( u2_uk_n217 ) );
  BUF_X1 u2_uk_U43 (.A( u2_uk_n141 ) , .Z( u2_uk_n222 ) );
  BUF_X1 u2_uk_U44 (.A( u2_uk_n182 ) , .Z( u2_uk_n220 ) );
  INV_X1 u2_uk_U446 (.ZN( u2_K10_33 ) , .A( u2_uk_n294 ) );
  AOI22_X1 u2_uk_U447 (.B2( u2_uk_K_r8_22 ) , .A2( u2_uk_K_r8_42 ) , .A1( u2_uk_n117 ) , .B1( u2_uk_n217 ) , .ZN( u2_uk_n294 ) );
  BUF_X1 u2_uk_U45 (.A( u2_uk_n203 ) , .Z( u2_uk_n207 ) );
  OAI22_X1 u2_uk_U453 (.ZN( u2_K14_33 ) , .A1( u2_uk_n155 ) , .B2( u2_uk_n1785 ) , .A2( u2_uk_n1803 ) , .B1( u2_uk_n83 ) );
  OAI22_X1 u2_uk_U457 (.ZN( u2_K6_33 ) , .B2( u2_uk_n1428 ) , .A2( u2_uk_n1433 ) , .A1( u2_uk_n188 ) , .B1( u2_uk_n60 ) );
  BUF_X1 u2_uk_U46 (.A( u2_uk_n155 ) , .Z( u2_uk_n217 ) );
  OAI22_X1 u2_uk_U460 (.ZN( u2_K15_37 ) , .A2( u2_uk_n1819 ) , .B2( u2_uk_n1846 ) , .A1( u2_uk_n223 ) , .B1( u2_uk_n99 ) );
  OAI21_X1 u2_uk_U468 (.ZN( u2_K6_37 ) , .A( u2_uk_n1068 ) , .B2( u2_uk_n1438 ) , .B1( u2_uk_n187 ) );
  NAND2_X1 u2_uk_U469 (.A1( u2_uk_K_r4_38 ) , .ZN( u2_uk_n1068 ) , .A2( u2_uk_n217 ) );
  BUF_X1 u2_uk_U47 (.Z( u2_uk_n223 ) , .A( u2_uk_n230 ) );
  OAI22_X1 u2_uk_U472 (.ZN( u2_K1_29 ) , .B2( u2_uk_n1152 ) , .A2( u2_uk_n1158 ) , .B1( u2_uk_n182 ) , .A1( u2_uk_n94 ) );
  OAI21_X1 u2_uk_U475 (.ZN( u2_K14_29 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1807 ) , .A( u2_uk_n689 ) );
  BUF_X1 u2_uk_U48 (.Z( u2_uk_n191 ) , .A( u2_uk_n217 ) );
  INV_X1 u2_uk_U483 (.ZN( u2_K4_29 ) , .A( u2_uk_n1030 ) );
  AOI22_X1 u2_uk_U484 (.B2( u2_uk_K_r2_31 ) , .A2( u2_uk_K_r2_36 ) , .ZN( u2_uk_n1030 ) , .B1( u2_uk_n191 ) , .A1( u2_uk_n83 ) );
  BUF_X1 u2_uk_U49 (.Z( u2_uk_n231 ) , .A( u2_uk_n238 ) );
  OAI22_X1 u2_uk_U493 (.ZN( u2_K7_29 ) , .B2( u2_uk_n1459 ) , .A2( u2_uk_n1490 ) , .A1( u2_uk_n238 ) , .B1( u2_uk_n31 ) );
  OAI21_X1 u2_uk_U497 (.ZN( u2_K10_2 ) , .B2( u2_uk_n1592 ) , .B1( u2_uk_n220 ) , .A( u2_uk_n286 ) );
  NAND2_X1 u2_uk_U498 (.A1( u2_uk_K_r8_41 ) , .A2( u2_uk_n230 ) , .ZN( u2_uk_n286 ) );
  INV_X1 u2_uk_U5 (.ZN( u2_uk_n117 ) , .A( u2_uk_n161 ) );
  BUF_X1 u2_uk_U50 (.Z( u2_uk_n230 ) , .A( u2_uk_n238 ) );
  OAI22_X1 u2_uk_U502 (.ZN( u2_K3_2 ) , .B2( u2_uk_n1301 ) , .A2( u2_uk_n1306 ) , .A1( u2_uk_n220 ) , .B1( u2_uk_n83 ) );
  OAI21_X1 u2_uk_U503 (.ZN( u2_K7_2 ) , .B1( u2_uk_n100 ) , .A( u2_uk_n1086 ) , .B2( u2_uk_n1454 ) );
  NAND2_X1 u2_uk_U504 (.A1( u2_uk_K_r5_41 ) , .ZN( u2_uk_n1086 ) , .A2( u2_uk_n63 ) );
  OAI21_X1 u2_uk_U512 (.ZN( u2_K9_17 ) , .B1( u2_uk_n102 ) , .A( u2_uk_n1122 ) , .B2( u2_uk_n1568 ) );
  NAND2_X1 u2_uk_U513 (.A1( u2_uk_K_r7_26 ) , .ZN( u2_uk_n1122 ) , .A2( u2_uk_n99 ) );
  OAI22_X1 u2_uk_U516 (.ZN( u2_K7_17 ) , .B2( u2_uk_n1458 ) , .A2( u2_uk_n1488 ) , .A1( u2_uk_n230 ) , .B1( u2_uk_n31 ) );
  OAI21_X1 u2_uk_U517 (.ZN( u2_K4_17 ) , .A( u2_uk_n1021 ) , .B2( u2_uk_n1339 ) , .B1( u2_uk_n187 ) );
  NAND2_X1 u2_uk_U518 (.A1( u2_uk_K_r2_27 ) , .ZN( u2_uk_n1021 ) , .A2( u2_uk_n155 ) );
  OAI22_X1 u2_uk_U519 (.ZN( u2_K3_17 ) , .B1( u2_uk_n10 ) , .B2( u2_uk_n1287 ) , .A2( u2_uk_n1310 ) , .A1( u2_uk_n202 ) );
  OAI21_X1 u2_uk_U523 (.ZN( u2_K12_12 ) , .B2( u2_uk_n1689 ) , .B1( u2_uk_n31 ) , .A( u2_uk_n408 ) );
  INV_X1 u2_uk_U525 (.ZN( u2_K7_12 ) , .A( u2_uk_n1075 ) );
  AOI22_X1 u2_uk_U526 (.B2( u2_uk_K_r5_17 ) , .A2( u2_uk_K_r5_39 ) , .ZN( u2_uk_n1075 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n230 ) );
  OAI21_X1 u2_uk_U527 (.ZN( u2_K5_12 ) , .A( u2_uk_n1041 ) , .B2( u2_uk_n1375 ) , .B1( u2_uk_n163 ) );
  NAND2_X1 u2_uk_U528 (.A1( u2_uk_K_r3_11 ) , .ZN( u2_uk_n1041 ) , .A2( u2_uk_n155 ) );
  OAI22_X1 u2_uk_U529 (.ZN( u2_K4_12 ) , .A1( u2_uk_n109 ) , .B2( u2_uk_n1341 ) , .A2( u2_uk_n1361 ) , .B1( u2_uk_n230 ) );
  OAI22_X1 u2_uk_U530 (.ZN( u2_K3_12 ) , .B1( u2_uk_n10 ) , .B2( u2_uk_n1306 ) , .A2( u2_uk_n1311 ) , .A1( u2_uk_n203 ) );
  OAI22_X1 u2_uk_U533 (.ZN( u2_K1_36 ) , .B2( u2_uk_n1158 ) , .A2( u2_uk_n1165 ) , .B1( u2_uk_n222 ) , .A1( u2_uk_n94 ) );
  INV_X1 u2_uk_U542 (.ZN( u2_K12_17 ) , .A( u2_uk_n415 ) );
  INV_X1 u2_uk_U546 (.ZN( u2_K6_17 ) , .A( u2_uk_n1059 ) );
  AOI22_X1 u2_uk_U547 (.B2( u2_uk_K_r4_4 ) , .A2( u2_uk_K_r4_55 ) , .ZN( u2_uk_n1059 ) , .B1( u2_uk_n118 ) , .A1( u2_uk_n147 ) );
  OAI22_X1 u2_uk_U548 (.ZN( u2_K15_36 ) , .B2( u2_uk_n1826 ) , .A2( u2_uk_n1840 ) , .A1( u2_uk_n222 ) , .B1( u2_uk_n92 ) );
  OAI22_X1 u2_uk_U549 (.ZN( u2_K14_36 ) , .A1( u2_uk_n141 ) , .B2( u2_uk_n1770 ) , .A2( u2_uk_n1808 ) , .B1( u2_uk_n63 ) );
  OAI22_X1 u2_uk_U551 (.ZN( u2_K3_36 ) , .B2( u2_uk_n1279 ) , .A1( u2_uk_n128 ) , .A2( u2_uk_n1314 ) , .B1( u2_uk_n145 ) );
  OAI22_X1 u2_uk_U553 (.ZN( u2_K1_38 ) , .A1( u2_uk_n10 ) , .B2( u2_uk_n1165 ) , .A2( u2_uk_n1171 ) , .B1( u2_uk_n203 ) );
  INV_X1 u2_uk_U557 (.ZN( u2_K7_36 ) , .A( u2_uk_n1091 ) );
  INV_X1 u2_uk_U561 (.ZN( u2_K5_36 ) , .A( u2_uk_n1050 ) );
  INV_X1 u2_uk_U564 (.ZN( u2_K15_38 ) , .A( u2_uk_n943 ) );
  INV_X1 u2_uk_U566 (.ZN( u2_K10_38 ) , .A( u2_uk_n301 ) );
  INV_X1 u2_uk_U579 (.ZN( u2_K9_10 ) , .A( u2_uk_n1117 ) );
  INV_X1 u2_uk_U58 (.ZN( u2_K7_34 ) , .A( u2_uk_n1089 ) );
  AOI22_X1 u2_uk_U580 (.B2( u2_uk_K_r7_25 ) , .A2( u2_uk_K_r7_32 ) , .B1( u2_uk_n110 ) , .ZN( u2_uk_n1117 ) , .A1( u2_uk_n163 ) );
  OAI22_X1 u2_uk_U587 (.ZN( u2_K3_22 ) , .B2( u2_uk_n1281 ) , .A2( u2_uk_n1316 ) , .B1( u2_uk_n141 ) , .A1( u2_uk_n94 ) );
  INV_X1 u2_uk_U595 (.ZN( u2_K9_22 ) , .A( u2_uk_n1127 ) );
  AOI22_X1 u2_uk_U596 (.B2( u2_uk_K_r7_41 ) , .A2( u2_uk_K_r7_48 ) , .B1( u2_uk_n109 ) , .ZN( u2_uk_n1127 ) , .A1( u2_uk_n213 ) );
  INV_X1 u2_uk_U6 (.A( u2_uk_n146 ) , .ZN( u2_uk_n17 ) );
  INV_X1 u2_uk_U614 (.ZN( u2_K10_35 ) , .A( u2_uk_n297 ) );
  AOI22_X1 u2_uk_U615 (.B2( u2_uk_K_r8_2 ) , .A2( u2_uk_K_r8_37 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n238 ) , .ZN( u2_uk_n297 ) );
  OAI22_X1 u2_uk_U618 (.ZN( u2_K6_35 ) , .B2( u2_uk_n1439 ) , .A2( u2_uk_n1446 ) , .A1( u2_uk_n217 ) , .B1( u2_uk_n60 ) );
  OAI22_X1 u2_uk_U625 (.ZN( u2_K7_11 ) , .B2( u2_uk_n1458 ) , .A2( u2_uk_n1475 ) , .B1( u2_uk_n208 ) , .A1( u2_uk_n93 ) );
  INV_X1 u2_uk_U635 (.ZN( u2_K9_11 ) , .A( u2_uk_n1118 ) );
  AOI22_X1 u2_uk_U636 (.B2( u2_uk_K_r7_48 ) , .A2( u2_uk_K_r7_55 ) , .B1( u2_uk_n100 ) , .ZN( u2_uk_n1118 ) , .A1( u2_uk_n223 ) );
  OAI22_X1 u2_uk_U639 (.ZN( u2_K3_11 ) , .A2( u2_uk_n1280 ) , .B2( u2_uk_n1285 ) , .B1( u2_uk_n141 ) , .A1( u2_uk_n99 ) );
  INV_X1 u2_uk_U644 (.ZN( u2_K1_44 ) , .A( u2_uk_n987 ) );
  INV_X1 u2_uk_U663 (.ZN( u2_K5_43 ) , .A( u2_uk_n1053 ) );
  OAI21_X1 u2_uk_U680 (.ZN( u2_K6_7 ) , .A( u2_uk_n1072 ) , .B2( u2_uk_n1435 ) , .B1( u2_uk_n238 ) );
  NAND2_X1 u2_uk_U681 (.A1( u2_uk_K_r4_33 ) , .ZN( u2_uk_n1072 ) , .A2( u2_uk_n217 ) );
  OAI21_X1 u2_uk_U682 (.ZN( u2_K3_3 ) , .A( u2_uk_n1013 ) , .B2( u2_uk_n1318 ) , .B1( u2_uk_n231 ) );
  NAND2_X1 u2_uk_U683 (.A1( u2_uk_K_r1_47 ) , .ZN( u2_uk_n1013 ) , .A2( u2_uk_n214 ) );
  INV_X1 u2_uk_U697 (.ZN( u2_K13_7 ) , .A( u2_uk_n682 ) );
  OAI21_X1 u2_uk_U699 (.ZN( u2_K5_7 ) , .A( u2_uk_n1057 ) , .B2( u2_uk_n1405 ) , .B1( u2_uk_n214 ) );
  INV_X1 u2_uk_U7 (.ZN( u2_uk_n11 ) , .A( u2_uk_n141 ) );
  NAND2_X1 u2_uk_U700 (.A1( u2_uk_K_r3_19 ) , .ZN( u2_uk_n1057 ) , .A2( u2_uk_n217 ) );
  INV_X1 u2_uk_U701 (.ZN( u2_K7_25 ) , .A( u2_uk_n1084 ) );
  INV_X1 u2_uk_U705 (.ZN( u2_K4_25 ) , .A( u2_uk_n1027 ) );
  OAI21_X1 u2_uk_U707 (.ZN( u2_K15_25 ) , .B1( u2_uk_n146 ) , .B2( u2_uk_n1846 ) , .A( u2_uk_n938 ) );
  NAND2_X1 u2_uk_U708 (.A1( u2_uk_K_r13_22 ) , .A2( u2_uk_n214 ) , .ZN( u2_uk_n938 ) );
  OAI22_X1 u2_uk_U713 (.ZN( u2_K4_32 ) , .A1( u2_uk_n109 ) , .A2( u2_uk_n1326 ) , .B2( u2_uk_n1350 ) , .B1( u2_uk_n209 ) );
  OAI22_X1 u2_uk_U723 (.ZN( u2_K14_32 ) , .A1( u2_uk_n155 ) , .B2( u2_uk_n1769 ) , .A2( u2_uk_n1807 ) , .B1( u2_uk_n83 ) );
  OAI22_X1 u2_uk_U727 (.ZN( u2_K15_42 ) , .B1( u2_uk_n161 ) , .B2( u2_uk_n1849 ) , .A2( u2_uk_n1855 ) , .A1( u2_uk_n31 ) );
  INV_X1 u2_uk_U737 (.ZN( u2_K7_42 ) , .A( u2_uk_n1093 ) );
  INV_X1 u2_uk_U739 (.ZN( u2_K1_42 ) , .A( u2_uk_n986 ) );
  OAI22_X1 u2_uk_U748 (.ZN( u2_K12_13 ) , .B2( u2_uk_n1689 ) , .A2( u2_uk_n1721 ) , .B1( u2_uk_n209 ) , .A1( u2_uk_n92 ) );
  OAI21_X1 u2_uk_U754 (.ZN( u2_K9_13 ) , .B1( u2_uk_n102 ) , .A( u2_uk_n1120 ) , .B2( u2_uk_n1549 ) );
  INV_X1 u2_uk_U76 (.ZN( u2_K4_23 ) , .A( u2_uk_n1026 ) );
  OAI22_X1 u2_uk_U761 (.ZN( u2_K9_21 ) , .A1( u2_uk_n117 ) , .B2( u2_uk_n1568 ) , .A2( u2_uk_n1573 ) , .B1( u2_uk_n208 ) );
  AOI22_X1 u2_uk_U77 (.B2( u2_uk_K_r2_18 ) , .A2( u2_uk_K_r2_55 ) , .ZN( u2_uk_n1026 ) , .B1( u2_uk_n191 ) , .A1( u2_uk_n83 ) );
  OAI22_X1 u2_uk_U775 (.ZN( u2_K4_13 ) , .A1( u2_uk_n102 ) , .A2( u2_uk_n1324 ) , .B2( u2_uk_n1328 ) , .B1( u2_uk_n230 ) );
  INV_X1 u2_uk_U778 (.ZN( u2_K6_21 ) , .A( u2_uk_n1062 ) );
  AOI22_X1 u2_uk_U779 (.B2( u2_uk_K_r4_11 ) , .A2( u2_uk_K_r4_5 ) , .ZN( u2_uk_n1062 ) , .B1( u2_uk_n118 ) , .A1( u2_uk_n217 ) );
  OAI21_X1 u2_uk_U782 (.ZN( u2_K7_21 ) , .A( u2_uk_n1080 ) , .B2( u2_uk_n1496 ) , .B1( u2_uk_n231 ) );
  NAND2_X1 u2_uk_U783 (.A1( u2_uk_K_r5_19 ) , .ZN( u2_uk_n1080 ) , .A2( u2_uk_n129 ) );
  INV_X1 u2_uk_U785 (.ZN( u2_K5_27 ) , .A( u2_uk_n1046 ) );
  INV_X1 u2_uk_U8 (.A( u2_uk_n145 ) , .ZN( u2_uk_n63 ) );
  OAI22_X1 u2_uk_U802 (.ZN( u2_K7_18 ) , .A2( u2_uk_n1453 ) , .B2( u2_uk_n1466 ) , .A1( u2_uk_n223 ) , .B1( u2_uk_n31 ) );
  INV_X1 u2_uk_U820 (.ZN( u2_K9_18 ) , .A( u2_uk_n1123 ) );
  INV_X1 u2_uk_U822 (.ZN( u2_K6_18 ) , .A( u2_uk_n1060 ) );
  AOI22_X1 u2_uk_U823 (.B2( u2_uk_K_r4_11 ) , .A2( u2_uk_K_r4_17 ) , .A1( u2_uk_n100 ) , .ZN( u2_uk_n1060 ) , .B1( u2_uk_n155 ) );
  INV_X1 u2_uk_U824 (.ZN( u2_K11_20 ) , .A( u2_uk_n342 ) );
  AOI22_X1 u2_uk_U825 (.B2( u2_uk_K_r9_10 ) , .A2( u2_uk_K_r9_4 ) , .A1( u2_uk_n110 ) , .B1( u2_uk_n162 ) , .ZN( u2_uk_n342 ) );
  INV_X1 u2_uk_U826 (.ZN( u2_K7_20 ) , .A( u2_uk_n1079 ) );
  OAI22_X1 u2_uk_U845 (.ZN( u2_K3_18 ) , .B1( u2_uk_n10 ) , .B2( u2_uk_n1295 ) , .A2( u2_uk_n1302 ) , .A1( u2_uk_n220 ) );
  OAI22_X1 u2_uk_U858 (.ZN( u2_K6_5 ) , .B2( u2_uk_n1422 ) , .A2( u2_uk_n1426 ) , .A1( u2_uk_n230 ) , .B1( u2_uk_n60 ) );
  OAI22_X1 u2_uk_U859 (.ZN( u2_K12_10 ) , .B1( u2_uk_n10 ) , .B2( u2_uk_n1688 ) , .A2( u2_uk_n1709 ) , .A1( u2_uk_n207 ) );
  OAI22_X1 u2_uk_U860 (.ZN( u2_K12_11 ) , .A1( u2_uk_n146 ) , .A2( u2_uk_n1683 ) , .B2( u2_uk_n1709 ) , .B1( u2_uk_n63 ) );
  OAI22_X1 u2_uk_U862 (.ZN( u2_K4_11 ) , .B2( u2_uk_n1333 ) , .A2( u2_uk_n1361 ) , .A1( u2_uk_n164 ) , .B1( u2_uk_n94 ) );
  OAI22_X1 u2_uk_U863 (.ZN( u2_K3_10 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1286 ) , .A1( u2_uk_n129 ) , .A2( u2_uk_n1291 ) );
  OAI22_X1 u2_uk_U873 (.ZN( u2_K9_7 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n146 ) , .A2( u2_uk_n1544 ) , .B2( u2_uk_n1548 ) );
  OAI22_X1 u2_uk_U874 (.ZN( u2_K6_12 ) , .A2( u2_uk_n1410 ) , .B2( u2_uk_n1426 ) , .A1( u2_uk_n207 ) , .B1( u2_uk_n93 ) );
  OAI22_X1 u2_uk_U875 (.ZN( u2_K7_14 ) , .B2( u2_uk_n1462 ) , .A2( u2_uk_n1497 ) , .A1( u2_uk_n222 ) , .B1( u2_uk_n31 ) );
  OAI22_X1 u2_uk_U880 (.ZN( u2_K3_21 ) , .B1( u2_uk_n109 ) , .B2( u2_uk_n1291 ) , .A2( u2_uk_n1316 ) , .A1( u2_uk_n161 ) );
  OAI22_X1 u2_uk_U881 (.ZN( u2_K9_24 ) , .B1( u2_uk_n128 ) , .B2( u2_uk_n1544 ) , .A2( u2_uk_n1586 ) , .A1( u2_uk_n220 ) );
  OAI22_X1 u2_uk_U893 (.ZN( u2_K4_36 ) , .B1( u2_uk_n109 ) , .B2( u2_uk_n1346 ) , .A2( u2_uk_n1351 ) , .A1( u2_uk_n161 ) );
  OAI22_X1 u2_uk_U895 (.ZN( u2_K6_30 ) , .B2( u2_uk_n1408 ) , .A2( u2_uk_n1413 ) , .A1( u2_uk_n164 ) , .B1( u2_uk_n60 ) );
  OAI22_X1 u2_uk_U896 (.ZN( u2_K3_25 ) , .B1( u2_uk_n117 ) , .B2( u2_uk_n1279 ) , .A2( u2_uk_n1283 ) , .A1( u2_uk_n207 ) );
  OAI22_X1 u2_uk_U899 (.ZN( u2_K7_39 ) , .B2( u2_uk_n1486 ) , .A2( u2_uk_n1493 ) , .A1( u2_uk_n161 ) , .B1( u2_uk_n31 ) );
  INV_X1 u2_uk_U9 (.A( u2_uk_n129 ) , .ZN( u2_uk_n31 ) );
  OAI22_X1 u2_uk_U90 (.ZN( u2_K7_41 ) , .A1( u2_uk_n118 ) , .A2( u2_uk_n1456 ) , .B2( u2_uk_n1486 ) , .B1( u2_uk_n208 ) );
  OAI22_X1 u2_uk_U900 (.ZN( u2_K6_42 ) , .B2( u2_uk_n1438 ) , .A2( u2_uk_n1445 ) , .A1( u2_uk_n163 ) , .B1( u2_uk_n60 ) );
  OAI22_X1 u2_uk_U903 (.ZN( u2_K3_38 ) , .B1( u2_uk_n128 ) , .A2( u2_uk_n1284 ) , .A1( u2_uk_n129 ) , .B2( u2_uk_n1300 ) );
  OAI22_X1 u2_uk_U913 (.ZN( u2_K9_6 ) , .A1( u2_uk_n100 ) , .B2( u2_uk_n1555 ) , .A2( u2_uk_n1563 ) , .B1( u2_uk_n217 ) );
  OAI22_X1 u2_uk_U914 (.ZN( u2_K9_8 ) , .B1( u2_uk_n129 ) , .B2( u2_uk_n1573 ) , .A2( u2_uk_n1580 ) , .A1( u2_uk_n92 ) );
  OAI22_X1 u2_uk_U916 (.ZN( u2_K12_18 ) , .A2( u2_uk_n1683 ) , .B2( u2_uk_n1721 ) , .B1( u2_uk_n231 ) , .A1( u2_uk_n92 ) );
  OAI22_X1 u2_uk_U923 (.ZN( u2_K15_47 ) , .A1( u2_uk_n117 ) , .B2( u2_uk_n1824 ) , .A2( u2_uk_n1856 ) , .B1( u2_uk_n220 ) );
  OAI22_X1 u2_uk_U928 (.ZN( u2_K6_46 ) , .A2( u2_uk_n1413 ) , .B2( u2_uk_n1441 ) , .B1( u2_uk_n208 ) , .A1( u2_uk_n93 ) );
  OAI22_X1 u2_uk_U930 (.ZN( u2_K9_4 ) , .A1( u2_uk_n110 ) , .B2( u2_uk_n1549 ) , .A2( u2_uk_n1556 ) , .B1( u2_uk_n231 ) );
  OAI22_X1 u2_uk_U938 (.ZN( u2_K12_19 ) , .A1( u2_uk_n128 ) , .A2( u2_uk_n1682 ) , .B2( u2_uk_n1720 ) , .B1( u2_uk_n231 ) );
  OAI22_X1 u2_uk_U939 (.ZN( u2_K15_19 ) , .A1( u2_uk_n118 ) , .B2( u2_uk_n1821 ) , .A2( u2_uk_n1851 ) , .B1( u2_uk_n207 ) );
  OAI22_X1 u2_uk_U954 (.ZN( u2_K6_43 ) , .B2( u2_uk_n1408 ) , .A2( u2_uk_n1447 ) , .B1( u2_uk_n182 ) , .A1( u2_uk_n93 ) );
  INV_X1 u2_uk_U96 (.ZN( u2_K13_5 ) , .A( u2_uk_n678 ) );
  OAI22_X1 u2_uk_U966 (.ZN( u2_K1_47 ) , .B2( u2_uk_n1142 ) , .A2( u2_uk_n1147 ) , .B1( u2_uk_n142 ) , .A1( u2_uk_n99 ) );
  AOI22_X1 u2_uk_U97 (.B2( u2_uk_K_r11_48 ) , .A2( u2_uk_K_r11_53 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n203 ) , .ZN( u2_uk_n678 ) );
  INV_X1 u2_uk_U970 (.ZN( u2_K12_42 ) , .A( u2_uk_n503 ) );
  OAI21_X1 u2_uk_U977 (.ZN( u2_K7_23 ) , .B1( u2_uk_n100 ) , .A( u2_uk_n1082 ) , .B2( u2_uk_n1453 ) );
  OAI22_X1 u2_uk_U98 (.ZN( u2_K12_5 ) , .A2( u2_uk_n1682 ) , .B2( u2_uk_n1708 ) , .A1( u2_uk_n202 ) , .B1( u2_uk_n94 ) );
  OAI21_X1 u2_uk_U985 (.ZN( u2_K4_5 ) , .A( u2_uk_n1038 ) , .B2( u2_uk_n1356 ) , .B1( u2_uk_n27 ) );
  OAI21_X1 u2_uk_U995 (.ZN( u2_K5_45 ) , .A( u2_uk_n1054 ) , .B2( u2_uk_n1370 ) , .B1( u2_uk_n27 ) );
  NAND2_X1 u2_uk_U996 (.A1( u2_uk_K_r3_43 ) , .ZN( u2_uk_n1054 ) , .A2( u2_uk_n17 ) );
  OAI21_X1 u2_uk_U997 (.ZN( u2_K3_45 ) , .A( u2_uk_n1016 ) , .B1( u2_uk_n102 ) , .B2( u2_uk_n1305 ) );
  NAND2_X1 u2_uk_U998 (.A1( u2_uk_K_r1_16 ) , .ZN( u2_uk_n1016 ) , .A2( u2_uk_n27 ) );
endmodule

