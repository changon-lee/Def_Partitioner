module des_des_die_12 ( u0_FP_33, u0_FP_40, u0_FP_41, u0_FP_42, u0_FP_43, u0_FP_44, u0_FP_45, u0_FP_46, u0_FP_47, 
       u0_FP_48, u0_FP_49, u0_FP_60, u0_FP_61, u0_FP_62, u0_FP_63, u0_FP_64, u0_K12_19, u0_K12_22, 
       u0_K12_7, u0_K12_9, u0_K16_18, u0_K16_19, u0_K16_22, u0_K16_24, u0_K1_30, u0_K1_31, u0_K1_45, 
       u0_K1_46, u0_K5_26, u0_K5_28, u0_K5_31, u0_K5_32, u0_K5_34, u0_K5_38, u0_K5_41, u0_L10_1, 
       u0_L10_10, u0_L10_13, u0_L10_16, u0_L10_17, u0_L10_18, u0_L10_2, u0_L10_20, u0_L10_23, u0_L10_24, 
       u0_L10_26, u0_L10_28, u0_L10_30, u0_L10_31, u0_L10_6, u0_L10_9, u0_L14_1, u0_L14_10, u0_L14_15, 
       u0_L14_16, u0_L14_20, u0_L14_21, u0_L14_24, u0_L14_26, u0_L14_27, u0_L14_30, u0_L14_5, u0_L14_6, 
       u0_L3_11, u0_L3_12, u0_L3_14, u0_L3_19, u0_L3_22, u0_L3_25, u0_L3_29, u0_L3_3, u0_L3_32, 
       u0_L3_4, u0_L3_7, u0_L3_8, u0_R10_1, u0_R10_10, u0_R10_11, u0_R10_12, u0_R10_13, u0_R10_14, 
       u0_R10_15, u0_R10_16, u0_R10_17, u0_R10_2, u0_R10_3, u0_R10_32, u0_R10_4, u0_R10_5, u0_R10_6, 
       u0_R10_7, u0_R10_8, u0_R10_9, u0_R3_16, u0_R3_17, u0_R3_18, u0_R3_19, u0_R3_20, u0_R3_21, 
       u0_R3_22, u0_R3_23, u0_R3_24, u0_R3_25, u0_R3_26, u0_R3_27, u0_R3_28, u0_R3_29, u0_desIn_r_0, 
       u0_desIn_r_1, u0_desIn_r_11, u0_desIn_r_16, u0_desIn_r_17, u0_desIn_r_18, u0_desIn_r_19, u0_desIn_r_20, u0_desIn_r_22, u0_desIn_r_25, 
       u0_desIn_r_27, u0_desIn_r_28, u0_desIn_r_3, u0_desIn_r_30, u0_desIn_r_32, u0_desIn_r_33, u0_desIn_r_34, u0_desIn_r_35, u0_desIn_r_38, 
       u0_desIn_r_41, u0_desIn_r_42, u0_desIn_r_43, u0_desIn_r_44, u0_desIn_r_49, u0_desIn_r_51, u0_desIn_r_52, u0_desIn_r_54, u0_desIn_r_56, 
       u0_desIn_r_57, u0_desIn_r_59, u0_desIn_r_61, u0_desIn_r_62, u0_desIn_r_7, u0_desIn_r_9, u0_key_r_0, u0_key_r_1, u0_key_r_14, 
       u0_key_r_16, u0_key_r_2, u0_key_r_21, u0_key_r_22, u0_key_r_23, u0_key_r_28, u0_key_r_29, u0_key_r_30, u0_key_r_31, 
       u0_key_r_35, u0_key_r_36, u0_key_r_37, u0_key_r_38, u0_key_r_42, u0_key_r_43, u0_key_r_50, u0_key_r_51, u0_key_r_52, 
       u0_key_r_7, u0_key_r_8, u0_key_r_9, u0_uk_K_r10_10, u0_uk_K_r10_18, u0_uk_K_r10_25, u0_uk_K_r10_27, u0_uk_K_r10_32, u0_uk_K_r10_34, 
       u0_uk_K_r10_39, u0_uk_K_r10_41, u0_uk_K_r10_47, u0_uk_K_r10_48, u0_uk_K_r14_10, u0_uk_K_r14_16, u0_uk_K_r14_18, u0_uk_K_r14_43, u0_uk_K_r14_46, 
       u0_uk_K_r14_9, u0_uk_K_r1_10, u0_uk_K_r2_29, u0_uk_K_r3_14, u0_uk_K_r3_16, u0_uk_K_r3_29, u0_uk_K_r3_35, u0_uk_K_r3_52, u0_uk_K_r3_9, 
       u0_uk_K_r9_38, u0_uk_n10, u0_uk_n100, u0_uk_n102, u0_uk_n109, u0_uk_n11, u0_uk_n110, u0_uk_n117, u0_uk_n118, 
       u0_uk_n128, u0_uk_n129, u0_uk_n136, u0_uk_n137, u0_uk_n141, u0_uk_n142, u0_uk_n143, u0_uk_n145, u0_uk_n146, 
       u0_uk_n147, u0_uk_n148, u0_uk_n149, u0_uk_n150, u0_uk_n155, u0_uk_n156, u0_uk_n157, u0_uk_n161, u0_uk_n163, 
       u0_uk_n164, u0_uk_n165, u0_uk_n166, u0_uk_n169, u0_uk_n170, u0_uk_n172, u0_uk_n175, u0_uk_n176, u0_uk_n177, 
       u0_uk_n182, u0_uk_n187, u0_uk_n188, u0_uk_n191, u0_uk_n202, u0_uk_n207, u0_uk_n209, u0_uk_n213, u0_uk_n220, 
       u0_uk_n222, u0_uk_n223, u0_uk_n230, u0_uk_n238, u0_uk_n240, u0_uk_n242, u0_uk_n250, u0_uk_n251, u0_uk_n252, 
       u0_uk_n257, u0_uk_n27, u0_uk_n31, u0_uk_n455, u0_uk_n457, u0_uk_n458, u0_uk_n462, u0_uk_n463, u0_uk_n475, 
       u0_uk_n476, u0_uk_n480, u0_uk_n481, u0_uk_n482, u0_uk_n493, u0_uk_n629, u0_uk_n631, u0_uk_n635, u0_uk_n636, 
       u0_uk_n638, u0_uk_n640, u0_uk_n641, u0_uk_n642, u0_uk_n644, u0_uk_n645, u0_uk_n650, u0_uk_n651, u0_uk_n652, 
       u0_uk_n653, u0_uk_n654, u0_uk_n658, u0_uk_n661, u0_uk_n666, u0_uk_n669, u0_uk_n670, u0_uk_n810, u0_uk_n813, 
       u0_uk_n83, u0_uk_n875, u0_uk_n878, u0_uk_n93, u0_uk_n94, u0_uk_n963, u0_uk_n981, u0_uk_n99, u2_K11_29, 
       u2_K13_14, u2_K13_3, u2_K13_37, u2_K13_40, u2_K13_42, u2_K13_44, u2_K13_45, u2_K13_46, u2_K13_47, 
       u2_K13_8, u2_K4_6, u2_K4_7, u2_K6_25, u2_K6_27, u2_K8_24, u2_K8_26, u2_K8_31, u2_K8_41, 
       u2_L11_12, u2_L11_13, u2_L11_15, u2_L11_16, u2_L11_17, u2_L11_18, u2_L11_2, u2_L11_21, u2_L11_22, 
       u2_L11_23, u2_L11_24, u2_L11_27, u2_L11_28, u2_L11_30, u2_L11_31, u2_L11_32, u2_L11_5, u2_L11_6, 
       u2_L11_7, u2_L11_9, u2_L2_13, u2_L2_15, u2_L2_17, u2_L2_18, u2_L2_2, u2_L2_21, u2_L2_23, 
       u2_L2_27, u2_L2_28, u2_L2_31, u2_L2_5, u2_L2_9, u2_L4_14, u2_L4_25, u2_L4_3, u2_L4_8, 
       u2_L6_1, u2_L6_10, u2_L6_11, u2_L6_12, u2_L6_14, u2_L6_19, u2_L6_20, u2_L6_22, u2_L6_25, 
       u2_L6_26, u2_L6_29, u2_L6_3, u2_L6_32, u2_L6_4, u2_L6_7, u2_L6_8, u2_L9_14, u2_L9_25, 
       u2_L9_3, u2_L9_8, u2_R11_1, u2_R11_10, u2_R11_11, u2_R11_12, u2_R11_13, u2_R11_2, u2_R11_24, 
       u2_R11_25, u2_R11_26, u2_R11_27, u2_R11_28, u2_R11_29, u2_R11_3, u2_R11_30, u2_R11_31, u2_R11_32, 
       u2_R11_4, u2_R11_5, u2_R11_6, u2_R11_7, u2_R11_8, u2_R11_9, u2_R2_1, u2_R2_2, u2_R2_28, 
       u2_R2_29, u2_R2_3, u2_R2_30, u2_R2_31, u2_R2_32, u2_R2_4, u2_R2_5, u2_R2_6, u2_R2_7, 
       u2_R2_8, u2_R2_9, u2_R4_16, u2_R4_17, u2_R4_18, u2_R4_19, u2_R4_20, u2_R4_21, u2_R6_12, 
       u2_R6_13, u2_R6_14, u2_R6_15, u2_R6_16, u2_R6_17, u2_R6_18, u2_R6_19, u2_R6_20, u2_R6_21, 
       u2_R6_22, u2_R6_23, u2_R6_24, u2_R6_25, u2_R6_26, u2_R6_27, u2_R6_28, u2_R6_29, u2_R9_16, 
       u2_R9_17, u2_R9_18, u2_R9_19, u2_R9_20, u2_R9_21, u2_uk_K_r11_11, u2_uk_K_r11_19, u2_uk_K_r11_20, u2_uk_K_r11_24, 
       u2_uk_K_r11_25, u2_uk_K_r11_26, u2_uk_K_r11_27, u2_uk_K_r11_29, u2_uk_K_r11_48, u2_uk_K_r11_53, u2_uk_K_r11_6, u2_uk_K_r2_13, u2_uk_K_r2_18, 
       u2_uk_K_r2_25, u2_uk_K_r2_26, u2_uk_K_r2_6, u2_uk_K_r4_0, u2_uk_K_r4_35, u2_uk_K_r6_14, u2_uk_K_r6_29, u2_uk_K_r6_31, u2_uk_K_r6_51, 
       u2_uk_K_r6_7, u2_uk_K_r9_1, u2_uk_K_r9_33, u2_uk_K_r9_5, u2_uk_K_r9_9, u2_uk_n102, u2_uk_n1031, u2_uk_n1035, u2_uk_n1036, 
       u2_uk_n1038, u2_uk_n1040, u2_uk_n109, u2_uk_n110, u2_uk_n1104, u2_uk_n1107, u2_uk_n1112, u2_uk_n117, u2_uk_n128, 
       u2_uk_n129, u2_uk_n1320, u2_uk_n1321, u2_uk_n1323, u2_uk_n1325, u2_uk_n1329, u2_uk_n1330, u2_uk_n1333, u2_uk_n1337, 
       u2_uk_n1339, u2_uk_n1341, u2_uk_n1344, u2_uk_n1350, u2_uk_n1353, u2_uk_n1356, u2_uk_n1359, u2_uk_n1360, u2_uk_n1361, 
       u2_uk_n1408, u2_uk_n1412, u2_uk_n1413, u2_uk_n1420, u2_uk_n1439, u2_uk_n1447, u2_uk_n145, u2_uk_n146, u2_uk_n147, 
       u2_uk_n148, u2_uk_n1498, u2_uk_n1499, u2_uk_n1503, u2_uk_n1504, u2_uk_n1508, u2_uk_n1510, u2_uk_n1511, u2_uk_n1513, 
       u2_uk_n1515, u2_uk_n1517, u2_uk_n1518, u2_uk_n1521, u2_uk_n1522, u2_uk_n1524, u2_uk_n1525, u2_uk_n1526, u2_uk_n1527, 
       u2_uk_n1528, u2_uk_n1529, u2_uk_n1530, u2_uk_n1531, u2_uk_n1532, u2_uk_n1533, u2_uk_n1535, u2_uk_n1536, u2_uk_n1538, 
       u2_uk_n155, u2_uk_n161, u2_uk_n162, u2_uk_n163, u2_uk_n164, u2_uk_n1642, u2_uk_n1647, u2_uk_n1654, u2_uk_n1660, 
       u2_uk_n1665, u2_uk_n1666, u2_uk_n1674, u2_uk_n17, u2_uk_n1723, u2_uk_n1725, u2_uk_n1727, u2_uk_n1731, u2_uk_n1732, 
       u2_uk_n1736, u2_uk_n1737, u2_uk_n1738, u2_uk_n1743, u2_uk_n1744, u2_uk_n1750, u2_uk_n1755, u2_uk_n1761, u2_uk_n1762, 
       u2_uk_n182, u2_uk_n188, u2_uk_n191, u2_uk_n202, u2_uk_n203, u2_uk_n208, u2_uk_n213, u2_uk_n214, u2_uk_n220, 
       u2_uk_n222, u2_uk_n223, u2_uk_n230, u2_uk_n231, u2_uk_n238, u2_uk_n363, u2_uk_n526, u2_uk_n551, u2_uk_n586, 
       u2_uk_n60, u2_uk_n63, u2_uk_n665, u2_uk_n677, u2_uk_n682, u2_uk_n83, u2_uk_n94, u2_uk_n99, u0_FP_1, u0_FP_10, u0_FP_15, u0_FP_16, u0_FP_20, u0_FP_21, u0_FP_24, u0_FP_26, u0_FP_27, 
        u0_FP_30, u0_FP_5, u0_FP_6, u0_N10, u0_N11, u0_N13, u0_N130, u0_N131, u0_N134, 
        u0_N135, u0_N138, u0_N139, u0_N14, u0_N141, u0_N146, u0_N149, u0_N152, u0_N156, 
        u0_N159, u0_N18, u0_N2, u0_N20, u0_N21, u0_N24, u0_N26, u0_N28, u0_N3, 
        u0_N31, u0_N352, u0_N353, u0_N357, u0_N360, u0_N361, u0_N364, u0_N367, u0_N368, 
        u0_N369, u0_N371, u0_N374, u0_N375, u0_N377, u0_N379, u0_N381, u0_N382, u0_N4, 
        u0_N6, u0_N7, u0_uk_n17, u0_uk_n208, u0_uk_n675, u0_uk_n687, u0_uk_n707, u0_uk_n711, u0_uk_n715, 
        u0_uk_n823, u0_uk_n841, u0_uk_n92, u0_uk_n989, u2_N100, u2_N104, u2_N108, u2_N110, u2_N112, 
        u2_N113, u2_N116, u2_N118, u2_N122, u2_N123, u2_N126, u2_N162, u2_N167, u2_N173, 
        u2_N184, u2_N224, u2_N226, u2_N227, u2_N230, u2_N231, u2_N233, u2_N234, u2_N235, 
        u2_N237, u2_N242, u2_N243, u2_N245, u2_N248, u2_N249, u2_N252, u2_N255, u2_N322, 
        u2_N327, u2_N333, u2_N344, u2_N385, u2_N388, u2_N389, u2_N390, u2_N392, u2_N395, 
        u2_N396, u2_N398, u2_N399, u2_N400, u2_N401, u2_N404, u2_N405, u2_N406, u2_N407, 
        u2_N410, u2_N411, u2_N413, u2_N414, u2_N415, u2_N97, u2_uk_n118, u2_uk_n187, u2_uk_n27, 
        u2_uk_n346, u2_uk_n395, u2_uk_n93 );
  input u0_FP_33, u0_FP_40, u0_FP_41, u0_FP_42, u0_FP_43, u0_FP_44, u0_FP_45, u0_FP_46, u0_FP_47, 
        u0_FP_48, u0_FP_49, u0_FP_60, u0_FP_61, u0_FP_62, u0_FP_63, u0_FP_64, u0_K12_19, u0_K12_22, 
        u0_K12_7, u0_K12_9, u0_K16_18, u0_K16_19, u0_K16_22, u0_K16_24, u0_K1_30, u0_K1_31, u0_K1_45, 
        u0_K1_46, u0_K5_26, u0_K5_28, u0_K5_31, u0_K5_32, u0_K5_34, u0_K5_38, u0_K5_41, u0_L10_1, 
        u0_L10_10, u0_L10_13, u0_L10_16, u0_L10_17, u0_L10_18, u0_L10_2, u0_L10_20, u0_L10_23, u0_L10_24, 
        u0_L10_26, u0_L10_28, u0_L10_30, u0_L10_31, u0_L10_6, u0_L10_9, u0_L14_1, u0_L14_10, u0_L14_15, 
        u0_L14_16, u0_L14_20, u0_L14_21, u0_L14_24, u0_L14_26, u0_L14_27, u0_L14_30, u0_L14_5, u0_L14_6, 
        u0_L3_11, u0_L3_12, u0_L3_14, u0_L3_19, u0_L3_22, u0_L3_25, u0_L3_29, u0_L3_3, u0_L3_32, 
        u0_L3_4, u0_L3_7, u0_L3_8, u0_R10_1, u0_R10_10, u0_R10_11, u0_R10_12, u0_R10_13, u0_R10_14, 
        u0_R10_15, u0_R10_16, u0_R10_17, u0_R10_2, u0_R10_3, u0_R10_32, u0_R10_4, u0_R10_5, u0_R10_6, 
        u0_R10_7, u0_R10_8, u0_R10_9, u0_R3_16, u0_R3_17, u0_R3_18, u0_R3_19, u0_R3_20, u0_R3_21, 
        u0_R3_22, u0_R3_23, u0_R3_24, u0_R3_25, u0_R3_26, u0_R3_27, u0_R3_28, u0_R3_29, u0_desIn_r_0, 
        u0_desIn_r_1, u0_desIn_r_11, u0_desIn_r_16, u0_desIn_r_17, u0_desIn_r_18, u0_desIn_r_19, u0_desIn_r_20, u0_desIn_r_22, u0_desIn_r_25, 
        u0_desIn_r_27, u0_desIn_r_28, u0_desIn_r_3, u0_desIn_r_30, u0_desIn_r_32, u0_desIn_r_33, u0_desIn_r_34, u0_desIn_r_35, u0_desIn_r_38, 
        u0_desIn_r_41, u0_desIn_r_42, u0_desIn_r_43, u0_desIn_r_44, u0_desIn_r_49, u0_desIn_r_51, u0_desIn_r_52, u0_desIn_r_54, u0_desIn_r_56, 
        u0_desIn_r_57, u0_desIn_r_59, u0_desIn_r_61, u0_desIn_r_62, u0_desIn_r_7, u0_desIn_r_9, u0_key_r_0, u0_key_r_1, u0_key_r_14, 
        u0_key_r_16, u0_key_r_2, u0_key_r_21, u0_key_r_22, u0_key_r_23, u0_key_r_28, u0_key_r_29, u0_key_r_30, u0_key_r_31, 
        u0_key_r_35, u0_key_r_36, u0_key_r_37, u0_key_r_38, u0_key_r_42, u0_key_r_43, u0_key_r_50, u0_key_r_51, u0_key_r_52, 
        u0_key_r_7, u0_key_r_8, u0_key_r_9, u0_uk_K_r10_10, u0_uk_K_r10_18, u0_uk_K_r10_25, u0_uk_K_r10_27, u0_uk_K_r10_32, u0_uk_K_r10_34, 
        u0_uk_K_r10_39, u0_uk_K_r10_41, u0_uk_K_r10_47, u0_uk_K_r10_48, u0_uk_K_r14_10, u0_uk_K_r14_16, u0_uk_K_r14_18, u0_uk_K_r14_43, u0_uk_K_r14_46, 
        u0_uk_K_r14_9, u0_uk_K_r1_10, u0_uk_K_r2_29, u0_uk_K_r3_14, u0_uk_K_r3_16, u0_uk_K_r3_29, u0_uk_K_r3_35, u0_uk_K_r3_52, u0_uk_K_r3_9, 
        u0_uk_K_r9_38, u0_uk_n10, u0_uk_n100, u0_uk_n102, u0_uk_n109, u0_uk_n11, u0_uk_n110, u0_uk_n117, u0_uk_n118, 
        u0_uk_n128, u0_uk_n129, u0_uk_n136, u0_uk_n137, u0_uk_n141, u0_uk_n142, u0_uk_n143, u0_uk_n145, u0_uk_n146, 
        u0_uk_n147, u0_uk_n148, u0_uk_n149, u0_uk_n150, u0_uk_n155, u0_uk_n156, u0_uk_n157, u0_uk_n161, u0_uk_n163, 
        u0_uk_n164, u0_uk_n165, u0_uk_n166, u0_uk_n169, u0_uk_n170, u0_uk_n172, u0_uk_n175, u0_uk_n176, u0_uk_n177, 
        u0_uk_n182, u0_uk_n187, u0_uk_n188, u0_uk_n191, u0_uk_n202, u0_uk_n207, u0_uk_n209, u0_uk_n213, u0_uk_n220, 
        u0_uk_n222, u0_uk_n223, u0_uk_n230, u0_uk_n238, u0_uk_n240, u0_uk_n242, u0_uk_n250, u0_uk_n251, u0_uk_n252, 
        u0_uk_n257, u0_uk_n27, u0_uk_n31, u0_uk_n455, u0_uk_n457, u0_uk_n458, u0_uk_n462, u0_uk_n463, u0_uk_n475, 
        u0_uk_n476, u0_uk_n480, u0_uk_n481, u0_uk_n482, u0_uk_n493, u0_uk_n629, u0_uk_n631, u0_uk_n635, u0_uk_n636, 
        u0_uk_n638, u0_uk_n640, u0_uk_n641, u0_uk_n642, u0_uk_n644, u0_uk_n645, u0_uk_n650, u0_uk_n651, u0_uk_n652, 
        u0_uk_n653, u0_uk_n654, u0_uk_n658, u0_uk_n661, u0_uk_n666, u0_uk_n669, u0_uk_n670, u0_uk_n810, u0_uk_n813, 
        u0_uk_n83, u0_uk_n875, u0_uk_n878, u0_uk_n93, u0_uk_n94, u0_uk_n963, u0_uk_n981, u0_uk_n99, u2_K11_29, 
        u2_K13_14, u2_K13_3, u2_K13_37, u2_K13_40, u2_K13_42, u2_K13_44, u2_K13_45, u2_K13_46, u2_K13_47, 
        u2_K13_8, u2_K4_6, u2_K4_7, u2_K6_25, u2_K6_27, u2_K8_24, u2_K8_26, u2_K8_31, u2_K8_41, 
        u2_L11_12, u2_L11_13, u2_L11_15, u2_L11_16, u2_L11_17, u2_L11_18, u2_L11_2, u2_L11_21, u2_L11_22, 
        u2_L11_23, u2_L11_24, u2_L11_27, u2_L11_28, u2_L11_30, u2_L11_31, u2_L11_32, u2_L11_5, u2_L11_6, 
        u2_L11_7, u2_L11_9, u2_L2_13, u2_L2_15, u2_L2_17, u2_L2_18, u2_L2_2, u2_L2_21, u2_L2_23, 
        u2_L2_27, u2_L2_28, u2_L2_31, u2_L2_5, u2_L2_9, u2_L4_14, u2_L4_25, u2_L4_3, u2_L4_8, 
        u2_L6_1, u2_L6_10, u2_L6_11, u2_L6_12, u2_L6_14, u2_L6_19, u2_L6_20, u2_L6_22, u2_L6_25, 
        u2_L6_26, u2_L6_29, u2_L6_3, u2_L6_32, u2_L6_4, u2_L6_7, u2_L6_8, u2_L9_14, u2_L9_25, 
        u2_L9_3, u2_L9_8, u2_R11_1, u2_R11_10, u2_R11_11, u2_R11_12, u2_R11_13, u2_R11_2, u2_R11_24, 
        u2_R11_25, u2_R11_26, u2_R11_27, u2_R11_28, u2_R11_29, u2_R11_3, u2_R11_30, u2_R11_31, u2_R11_32, 
        u2_R11_4, u2_R11_5, u2_R11_6, u2_R11_7, u2_R11_8, u2_R11_9, u2_R2_1, u2_R2_2, u2_R2_28, 
        u2_R2_29, u2_R2_3, u2_R2_30, u2_R2_31, u2_R2_32, u2_R2_4, u2_R2_5, u2_R2_6, u2_R2_7, 
        u2_R2_8, u2_R2_9, u2_R4_16, u2_R4_17, u2_R4_18, u2_R4_19, u2_R4_20, u2_R4_21, u2_R6_12, 
        u2_R6_13, u2_R6_14, u2_R6_15, u2_R6_16, u2_R6_17, u2_R6_18, u2_R6_19, u2_R6_20, u2_R6_21, 
        u2_R6_22, u2_R6_23, u2_R6_24, u2_R6_25, u2_R6_26, u2_R6_27, u2_R6_28, u2_R6_29, u2_R9_16, 
        u2_R9_17, u2_R9_18, u2_R9_19, u2_R9_20, u2_R9_21, u2_uk_K_r11_11, u2_uk_K_r11_19, u2_uk_K_r11_20, u2_uk_K_r11_24, 
        u2_uk_K_r11_25, u2_uk_K_r11_26, u2_uk_K_r11_27, u2_uk_K_r11_29, u2_uk_K_r11_48, u2_uk_K_r11_53, u2_uk_K_r11_6, u2_uk_K_r2_13, u2_uk_K_r2_18, 
        u2_uk_K_r2_25, u2_uk_K_r2_26, u2_uk_K_r2_6, u2_uk_K_r4_0, u2_uk_K_r4_35, u2_uk_K_r6_14, u2_uk_K_r6_29, u2_uk_K_r6_31, u2_uk_K_r6_51, 
        u2_uk_K_r6_7, u2_uk_K_r9_1, u2_uk_K_r9_33, u2_uk_K_r9_5, u2_uk_K_r9_9, u2_uk_n102, u2_uk_n1031, u2_uk_n1035, u2_uk_n1036, 
        u2_uk_n1038, u2_uk_n1040, u2_uk_n109, u2_uk_n110, u2_uk_n1104, u2_uk_n1107, u2_uk_n1112, u2_uk_n117, u2_uk_n128, 
        u2_uk_n129, u2_uk_n1320, u2_uk_n1321, u2_uk_n1323, u2_uk_n1325, u2_uk_n1329, u2_uk_n1330, u2_uk_n1333, u2_uk_n1337, 
        u2_uk_n1339, u2_uk_n1341, u2_uk_n1344, u2_uk_n1350, u2_uk_n1353, u2_uk_n1356, u2_uk_n1359, u2_uk_n1360, u2_uk_n1361, 
        u2_uk_n1408, u2_uk_n1412, u2_uk_n1413, u2_uk_n1420, u2_uk_n1439, u2_uk_n1447, u2_uk_n145, u2_uk_n146, u2_uk_n147, 
        u2_uk_n148, u2_uk_n1498, u2_uk_n1499, u2_uk_n1503, u2_uk_n1504, u2_uk_n1508, u2_uk_n1510, u2_uk_n1511, u2_uk_n1513, 
        u2_uk_n1515, u2_uk_n1517, u2_uk_n1518, u2_uk_n1521, u2_uk_n1522, u2_uk_n1524, u2_uk_n1525, u2_uk_n1526, u2_uk_n1527, 
        u2_uk_n1528, u2_uk_n1529, u2_uk_n1530, u2_uk_n1531, u2_uk_n1532, u2_uk_n1533, u2_uk_n1535, u2_uk_n1536, u2_uk_n1538, 
        u2_uk_n155, u2_uk_n161, u2_uk_n162, u2_uk_n163, u2_uk_n164, u2_uk_n1642, u2_uk_n1647, u2_uk_n1654, u2_uk_n1660, 
        u2_uk_n1665, u2_uk_n1666, u2_uk_n1674, u2_uk_n17, u2_uk_n1723, u2_uk_n1725, u2_uk_n1727, u2_uk_n1731, u2_uk_n1732, 
        u2_uk_n1736, u2_uk_n1737, u2_uk_n1738, u2_uk_n1743, u2_uk_n1744, u2_uk_n1750, u2_uk_n1755, u2_uk_n1761, u2_uk_n1762, 
        u2_uk_n182, u2_uk_n188, u2_uk_n191, u2_uk_n202, u2_uk_n203, u2_uk_n208, u2_uk_n213, u2_uk_n214, u2_uk_n220, 
        u2_uk_n222, u2_uk_n223, u2_uk_n230, u2_uk_n231, u2_uk_n238, u2_uk_n363, u2_uk_n526, u2_uk_n551, u2_uk_n586, 
        u2_uk_n60, u2_uk_n63, u2_uk_n665, u2_uk_n677, u2_uk_n682, u2_uk_n83, u2_uk_n94, u2_uk_n99;
  output u0_FP_1, u0_FP_10, u0_FP_15, u0_FP_16, u0_FP_20, u0_FP_21, u0_FP_24, u0_FP_26, u0_FP_27, 
        u0_FP_30, u0_FP_5, u0_FP_6, u0_N10, u0_N11, u0_N13, u0_N130, u0_N131, u0_N134, 
        u0_N135, u0_N138, u0_N139, u0_N14, u0_N141, u0_N146, u0_N149, u0_N152, u0_N156, 
        u0_N159, u0_N18, u0_N2, u0_N20, u0_N21, u0_N24, u0_N26, u0_N28, u0_N3, 
        u0_N31, u0_N352, u0_N353, u0_N357, u0_N360, u0_N361, u0_N364, u0_N367, u0_N368, 
        u0_N369, u0_N371, u0_N374, u0_N375, u0_N377, u0_N379, u0_N381, u0_N382, u0_N4, 
        u0_N6, u0_N7, u0_uk_n17, u0_uk_n208, u0_uk_n675, u0_uk_n687, u0_uk_n707, u0_uk_n711, u0_uk_n715, 
        u0_uk_n823, u0_uk_n841, u0_uk_n92, u0_uk_n989, u2_N100, u2_N104, u2_N108, u2_N110, u2_N112, 
        u2_N113, u2_N116, u2_N118, u2_N122, u2_N123, u2_N126, u2_N162, u2_N167, u2_N173, 
        u2_N184, u2_N224, u2_N226, u2_N227, u2_N230, u2_N231, u2_N233, u2_N234, u2_N235, 
        u2_N237, u2_N242, u2_N243, u2_N245, u2_N248, u2_N249, u2_N252, u2_N255, u2_N322, 
        u2_N327, u2_N333, u2_N344, u2_N385, u2_N388, u2_N389, u2_N390, u2_N392, u2_N395, 
        u2_N396, u2_N398, u2_N399, u2_N400, u2_N401, u2_N404, u2_N405, u2_N406, u2_N407, 
        u2_N410, u2_N411, u2_N413, u2_N414, u2_N415, u2_N97, u2_uk_n118, u2_uk_n187, u2_uk_n27, 
        u2_uk_n346, u2_uk_n395, u2_uk_n93;
  wire u0_K12_1, u0_K12_10, u0_K12_11, u0_K12_12, u0_K12_13, u0_K12_14, u0_K12_15, u0_K12_16, u0_K12_17, 
       u0_K12_18, u0_K12_2, u0_K12_20, u0_K12_21, u0_K12_23, u0_K12_24, u0_K12_3, u0_K12_4, u0_K12_5, 
       u0_K12_6, u0_K12_8, u0_K16_13, u0_K16_14, u0_K16_15, u0_K16_16, u0_K16_17, u0_K16_20, u0_K16_21, 
       u0_K16_23, u0_K16_43, u0_K16_44, u0_K16_45, u0_K16_46, u0_K16_47, u0_K16_48, u0_K1_25, u0_K1_26, 
       u0_K1_27, u0_K1_28, u0_K1_29, u0_K1_32, u0_K1_33, u0_K1_34, u0_K1_35, u0_K1_36, u0_K1_37, 
       u0_K1_38, u0_K1_39, u0_K1_40, u0_K1_41, u0_K1_42, u0_K1_43, u0_K1_44, u0_K1_47, u0_K1_48, 
       u0_K5_25, u0_K5_27, u0_K5_29, u0_K5_30, u0_K5_33, u0_K5_35, u0_K5_36, u0_K5_37, u0_K5_39, 
       u0_K5_40, u0_K5_42, u0_out0_11, u0_out0_12, u0_out0_14, u0_out0_15, u0_out0_19, u0_out0_21, u0_out0_22, 
       u0_out0_25, u0_out0_27, u0_out0_29, u0_out0_3, u0_out0_32, u0_out0_4, u0_out0_5, u0_out0_7, u0_out0_8, 
       u0_out11_1, u0_out11_10, u0_out11_13, u0_out11_16, u0_out11_17, u0_out11_18, u0_out11_2, u0_out11_20, u0_out11_23, 
       u0_out11_24, u0_out11_26, u0_out11_28, u0_out11_30, u0_out11_31, u0_out11_6, u0_out11_9, u0_out15_1, u0_out15_10, 
       u0_out15_15, u0_out15_16, u0_out15_20, u0_out15_21, u0_out15_24, u0_out15_26, u0_out15_27, u0_out15_30, u0_out15_5, 
       u0_out15_6, u0_out4_11, u0_out4_12, u0_out4_14, u0_out4_19, u0_out4_22, u0_out4_25, u0_out4_29, u0_out4_3, 
       u0_out4_32, u0_out4_4, u0_out4_7, u0_out4_8, u0_u0_X_25, u0_u0_X_26, u0_u0_X_27, u0_u0_X_28, u0_u0_X_29, 
       u0_u0_X_30, u0_u0_X_31, u0_u0_X_32, u0_u0_X_33, u0_u0_X_34, u0_u0_X_35, u0_u0_X_36, u0_u0_X_37, u0_u0_X_38, 
       u0_u0_X_39, u0_u0_X_40, u0_u0_X_41, u0_u0_X_42, u0_u0_X_43, u0_u0_X_44, u0_u0_X_45, u0_u0_X_46, u0_u0_X_47, 
       u0_u0_X_48, u0_u0_u4_n1, u0_u0_u4_n10, u0_u0_u4_n11, u0_u0_u4_n12, u0_u0_u4_n13, u0_u0_u4_n14, u0_u0_u4_n15, u0_u0_u4_n16, 
       u0_u0_u4_n17, u0_u0_u4_n18, u0_u0_u4_n19, u0_u0_u4_n2, u0_u0_u4_n20, u0_u0_u4_n21, u0_u0_u4_n22, u0_u0_u4_n23, u0_u0_u4_n24, 
       u0_u0_u4_n25, u0_u0_u4_n26, u0_u0_u4_n27, u0_u0_u4_n28, u0_u0_u4_n29, u0_u0_u4_n3, u0_u0_u4_n30, u0_u0_u4_n31, u0_u0_u4_n32, 
       u0_u0_u4_n33, u0_u0_u4_n34, u0_u0_u4_n35, u0_u0_u4_n36, u0_u0_u4_n37, u0_u0_u4_n38, u0_u0_u4_n39, u0_u0_u4_n4, u0_u0_u4_n40, 
       u0_u0_u4_n41, u0_u0_u4_n42, u0_u0_u4_n43, u0_u0_u4_n44, u0_u0_u4_n45, u0_u0_u4_n46, u0_u0_u4_n47, u0_u0_u4_n48, u0_u0_u4_n49, 
       u0_u0_u4_n5, u0_u0_u4_n50, u0_u0_u4_n51, u0_u0_u4_n52, u0_u0_u4_n53, u0_u0_u4_n54, u0_u0_u4_n55, u0_u0_u4_n56, u0_u0_u4_n57, 
       u0_u0_u4_n58, u0_u0_u4_n59, u0_u0_u4_n6, u0_u0_u4_n60, u0_u0_u4_n61, u0_u0_u4_n62, u0_u0_u4_n63, u0_u0_u4_n64, u0_u0_u4_n65, 
       u0_u0_u4_n66, u0_u0_u4_n67, u0_u0_u4_n68, u0_u0_u4_n69, u0_u0_u4_n7, u0_u0_u4_n70, u0_u0_u4_n71, u0_u0_u4_n72, u0_u0_u4_n73, 
       u0_u0_u4_n74, u0_u0_u4_n75, u0_u0_u4_n76, u0_u0_u4_n77, u0_u0_u4_n78, u0_u0_u4_n79, u0_u0_u4_n8, u0_u0_u4_n80, u0_u0_u4_n81, 
       u0_u0_u4_n82, u0_u0_u4_n83, u0_u0_u4_n84, u0_u0_u4_n85, u0_u0_u4_n86, u0_u0_u4_n87, u0_u0_u4_n88, u0_u0_u4_n89, u0_u0_u4_n9, 
       u0_u0_u4_n90, u0_u0_u4_n91, u0_u0_u4_n92, u0_u0_u4_n93, u0_u0_u5_n1, u0_u0_u5_n10, u0_u0_u5_n11, u0_u0_u5_n12, u0_u0_u5_n13, 
       u0_u0_u5_n14, u0_u0_u5_n15, u0_u0_u5_n16, u0_u0_u5_n17, u0_u0_u5_n18, u0_u0_u5_n19, u0_u0_u5_n2, u0_u0_u5_n20, u0_u0_u5_n21, 
       u0_u0_u5_n22, u0_u0_u5_n23, u0_u0_u5_n24, u0_u0_u5_n25, u0_u0_u5_n26, u0_u0_u5_n27, u0_u0_u5_n28, u0_u0_u5_n29, u0_u0_u5_n3, 
       u0_u0_u5_n30, u0_u0_u5_n31, u0_u0_u5_n32, u0_u0_u5_n33, u0_u0_u5_n34, u0_u0_u5_n35, u0_u0_u5_n36, u0_u0_u5_n37, u0_u0_u5_n38, 
       u0_u0_u5_n39, u0_u0_u5_n4, u0_u0_u5_n40, u0_u0_u5_n41, u0_u0_u5_n42, u0_u0_u5_n43, u0_u0_u5_n44, u0_u0_u5_n45, u0_u0_u5_n46, 
       u0_u0_u5_n47, u0_u0_u5_n48, u0_u0_u5_n49, u0_u0_u5_n5, u0_u0_u5_n50, u0_u0_u5_n51, u0_u0_u5_n52, u0_u0_u5_n53, u0_u0_u5_n54, 
       u0_u0_u5_n55, u0_u0_u5_n56, u0_u0_u5_n57, u0_u0_u5_n58, u0_u0_u5_n59, u0_u0_u5_n6, u0_u0_u5_n60, u0_u0_u5_n61, u0_u0_u5_n62, 
       u0_u0_u5_n63, u0_u0_u5_n64, u0_u0_u5_n65, u0_u0_u5_n66, u0_u0_u5_n67, u0_u0_u5_n68, u0_u0_u5_n69, u0_u0_u5_n7, u0_u0_u5_n70, 
       u0_u0_u5_n71, u0_u0_u5_n72, u0_u0_u5_n73, u0_u0_u5_n74, u0_u0_u5_n75, u0_u0_u5_n76, u0_u0_u5_n77, u0_u0_u5_n78, u0_u0_u5_n79, 
       u0_u0_u5_n8, u0_u0_u5_n80, u0_u0_u5_n81, u0_u0_u5_n82, u0_u0_u5_n83, u0_u0_u5_n84, u0_u0_u5_n85, u0_u0_u5_n86, u0_u0_u5_n87, 
       u0_u0_u5_n88, u0_u0_u5_n89, u0_u0_u5_n9, u0_u0_u5_n90, u0_u0_u5_n91, u0_u0_u5_n92, u0_u0_u5_n93, u0_u0_u5_n94, u0_u0_u5_n95, 
       u0_u0_u5_n96, u0_u0_u5_n97, u0_u0_u5_n98, u0_u0_u6_n1, u0_u0_u6_n10, u0_u0_u6_n11, u0_u0_u6_n12, u0_u0_u6_n13, u0_u0_u6_n14, 
       u0_u0_u6_n15, u0_u0_u6_n16, u0_u0_u6_n17, u0_u0_u6_n18, u0_u0_u6_n19, u0_u0_u6_n2, u0_u0_u6_n20, u0_u0_u6_n21, u0_u0_u6_n22, 
       u0_u0_u6_n23, u0_u0_u6_n24, u0_u0_u6_n25, u0_u0_u6_n26, u0_u0_u6_n27, u0_u0_u6_n28, u0_u0_u6_n29, u0_u0_u6_n3, u0_u0_u6_n30, 
       u0_u0_u6_n31, u0_u0_u6_n32, u0_u0_u6_n33, u0_u0_u6_n34, u0_u0_u6_n35, u0_u0_u6_n36, u0_u0_u6_n37, u0_u0_u6_n38, u0_u0_u6_n39, 
       u0_u0_u6_n4, u0_u0_u6_n40, u0_u0_u6_n41, u0_u0_u6_n42, u0_u0_u6_n43, u0_u0_u6_n44, u0_u0_u6_n45, u0_u0_u6_n46, u0_u0_u6_n47, 
       u0_u0_u6_n48, u0_u0_u6_n49, u0_u0_u6_n5, u0_u0_u6_n50, u0_u0_u6_n51, u0_u0_u6_n52, u0_u0_u6_n53, u0_u0_u6_n54, u0_u0_u6_n55, 
       u0_u0_u6_n56, u0_u0_u6_n57, u0_u0_u6_n58, u0_u0_u6_n59, u0_u0_u6_n6, u0_u0_u6_n60, u0_u0_u6_n61, u0_u0_u6_n62, u0_u0_u6_n63, 
       u0_u0_u6_n64, u0_u0_u6_n65, u0_u0_u6_n66, u0_u0_u6_n67, u0_u0_u6_n68, u0_u0_u6_n69, u0_u0_u6_n7, u0_u0_u6_n70, u0_u0_u6_n71, 
       u0_u0_u6_n72, u0_u0_u6_n73, u0_u0_u6_n74, u0_u0_u6_n75, u0_u0_u6_n76, u0_u0_u6_n77, u0_u0_u6_n78, u0_u0_u6_n79, u0_u0_u6_n8, 
       u0_u0_u6_n80, u0_u0_u6_n81, u0_u0_u6_n82, u0_u0_u6_n83, u0_u0_u6_n84, u0_u0_u6_n85, u0_u0_u6_n86, u0_u0_u6_n87, u0_u0_u6_n9, 
       u0_u0_u7_n1, u0_u0_u7_n10, u0_u0_u7_n11, u0_u0_u7_n12, u0_u0_u7_n13, u0_u0_u7_n14, u0_u0_u7_n15, u0_u0_u7_n16, u0_u0_u7_n17, 
       u0_u0_u7_n18, u0_u0_u7_n19, u0_u0_u7_n2, u0_u0_u7_n20, u0_u0_u7_n21, u0_u0_u7_n22, u0_u0_u7_n23, u0_u0_u7_n24, u0_u0_u7_n25, 
       u0_u0_u7_n26, u0_u0_u7_n27, u0_u0_u7_n28, u0_u0_u7_n29, u0_u0_u7_n3, u0_u0_u7_n30, u0_u0_u7_n31, u0_u0_u7_n32, u0_u0_u7_n33, 
       u0_u0_u7_n34, u0_u0_u7_n35, u0_u0_u7_n36, u0_u0_u7_n37, u0_u0_u7_n38, u0_u0_u7_n39, u0_u0_u7_n4, u0_u0_u7_n40, u0_u0_u7_n41, 
       u0_u0_u7_n42, u0_u0_u7_n43, u0_u0_u7_n44, u0_u0_u7_n45, u0_u0_u7_n46, u0_u0_u7_n47, u0_u0_u7_n48, u0_u0_u7_n49, u0_u0_u7_n5, 
       u0_u0_u7_n50, u0_u0_u7_n51, u0_u0_u7_n52, u0_u0_u7_n53, u0_u0_u7_n54, u0_u0_u7_n55, u0_u0_u7_n56, u0_u0_u7_n57, u0_u0_u7_n58, 
       u0_u0_u7_n59, u0_u0_u7_n6, u0_u0_u7_n60, u0_u0_u7_n61, u0_u0_u7_n62, u0_u0_u7_n63, u0_u0_u7_n64, u0_u0_u7_n65, u0_u0_u7_n66, 
       u0_u0_u7_n67, u0_u0_u7_n68, u0_u0_u7_n69, u0_u0_u7_n7, u0_u0_u7_n70, u0_u0_u7_n71, u0_u0_u7_n72, u0_u0_u7_n73, u0_u0_u7_n74, 
       u0_u0_u7_n75, u0_u0_u7_n76, u0_u0_u7_n77, u0_u0_u7_n78, u0_u0_u7_n79, u0_u0_u7_n8, u0_u0_u7_n80, u0_u0_u7_n81, u0_u0_u7_n82, 
       u0_u0_u7_n83, u0_u0_u7_n84, u0_u0_u7_n85, u0_u0_u7_n86, u0_u0_u7_n87, u0_u0_u7_n88, u0_u0_u7_n89, u0_u0_u7_n9, u0_u0_u7_n90, 
       u0_u11_X_1, u0_u11_X_10, u0_u11_X_11, u0_u11_X_12, u0_u11_X_13, u0_u11_X_14, u0_u11_X_15, u0_u11_X_16, u0_u11_X_17, 
       u0_u11_X_18, u0_u11_X_19, u0_u11_X_2, u0_u11_X_20, u0_u11_X_21, u0_u11_X_22, u0_u11_X_23, u0_u11_X_24, u0_u11_X_3, 
       u0_u11_X_4, u0_u11_X_5, u0_u11_X_6, u0_u11_X_7, u0_u11_X_8, u0_u11_X_9, u0_u11_u0_n100, u0_u11_u0_n101, u0_u11_u0_n102, 
       u0_u11_u0_n103, u0_u11_u0_n104, u0_u11_u0_n105, u0_u11_u0_n106, u0_u11_u0_n107, u0_u11_u0_n108, u0_u11_u0_n109, u0_u11_u0_n110, u0_u11_u0_n111, 
       u0_u11_u0_n112, u0_u11_u0_n113, u0_u11_u0_n114, u0_u11_u0_n115, u0_u11_u0_n116, u0_u11_u0_n117, u0_u11_u0_n118, u0_u11_u0_n119, u0_u11_u0_n120, 
       u0_u11_u0_n121, u0_u11_u0_n122, u0_u11_u0_n123, u0_u11_u0_n124, u0_u11_u0_n125, u0_u11_u0_n126, u0_u11_u0_n127, u0_u11_u0_n128, u0_u11_u0_n129, 
       u0_u11_u0_n130, u0_u11_u0_n131, u0_u11_u0_n132, u0_u11_u0_n133, u0_u11_u0_n134, u0_u11_u0_n135, u0_u11_u0_n136, u0_u11_u0_n137, u0_u11_u0_n138, 
       u0_u11_u0_n139, u0_u11_u0_n140, u0_u11_u0_n141, u0_u11_u0_n142, u0_u11_u0_n143, u0_u11_u0_n144, u0_u11_u0_n145, u0_u11_u0_n146, u0_u11_u0_n147, 
       u0_u11_u0_n148, u0_u11_u0_n149, u0_u11_u0_n150, u0_u11_u0_n151, u0_u11_u0_n152, u0_u11_u0_n153, u0_u11_u0_n154, u0_u11_u0_n155, u0_u11_u0_n156, 
       u0_u11_u0_n157, u0_u11_u0_n158, u0_u11_u0_n159, u0_u11_u0_n160, u0_u11_u0_n161, u0_u11_u0_n162, u0_u11_u0_n163, u0_u11_u0_n164, u0_u11_u0_n165, 
       u0_u11_u0_n166, u0_u11_u0_n167, u0_u11_u0_n168, u0_u11_u0_n169, u0_u11_u0_n170, u0_u11_u0_n171, u0_u11_u0_n172, u0_u11_u0_n173, u0_u11_u0_n174, 
       u0_u11_u0_n88, u0_u11_u0_n89, u0_u11_u0_n90, u0_u11_u0_n91, u0_u11_u0_n92, u0_u11_u0_n93, u0_u11_u0_n94, u0_u11_u0_n95, u0_u11_u0_n96, 
       u0_u11_u0_n97, u0_u11_u0_n98, u0_u11_u0_n99, u0_u11_u1_n100, u0_u11_u1_n101, u0_u11_u1_n102, u0_u11_u1_n103, u0_u11_u1_n104, u0_u11_u1_n105, 
       u0_u11_u1_n106, u0_u11_u1_n107, u0_u11_u1_n108, u0_u11_u1_n109, u0_u11_u1_n110, u0_u11_u1_n111, u0_u11_u1_n112, u0_u11_u1_n113, u0_u11_u1_n114, 
       u0_u11_u1_n115, u0_u11_u1_n116, u0_u11_u1_n117, u0_u11_u1_n118, u0_u11_u1_n119, u0_u11_u1_n120, u0_u11_u1_n121, u0_u11_u1_n122, u0_u11_u1_n123, 
       u0_u11_u1_n124, u0_u11_u1_n125, u0_u11_u1_n126, u0_u11_u1_n127, u0_u11_u1_n128, u0_u11_u1_n129, u0_u11_u1_n130, u0_u11_u1_n131, u0_u11_u1_n132, 
       u0_u11_u1_n133, u0_u11_u1_n134, u0_u11_u1_n135, u0_u11_u1_n136, u0_u11_u1_n137, u0_u11_u1_n138, u0_u11_u1_n139, u0_u11_u1_n140, u0_u11_u1_n141, 
       u0_u11_u1_n142, u0_u11_u1_n143, u0_u11_u1_n144, u0_u11_u1_n145, u0_u11_u1_n146, u0_u11_u1_n147, u0_u11_u1_n148, u0_u11_u1_n149, u0_u11_u1_n150, 
       u0_u11_u1_n151, u0_u11_u1_n152, u0_u11_u1_n153, u0_u11_u1_n154, u0_u11_u1_n155, u0_u11_u1_n156, u0_u11_u1_n157, u0_u11_u1_n158, u0_u11_u1_n159, 
       u0_u11_u1_n160, u0_u11_u1_n161, u0_u11_u1_n162, u0_u11_u1_n163, u0_u11_u1_n164, u0_u11_u1_n165, u0_u11_u1_n166, u0_u11_u1_n167, u0_u11_u1_n168, 
       u0_u11_u1_n169, u0_u11_u1_n170, u0_u11_u1_n171, u0_u11_u1_n172, u0_u11_u1_n173, u0_u11_u1_n174, u0_u11_u1_n175, u0_u11_u1_n176, u0_u11_u1_n177, 
       u0_u11_u1_n178, u0_u11_u1_n179, u0_u11_u1_n180, u0_u11_u1_n181, u0_u11_u1_n182, u0_u11_u1_n183, u0_u11_u1_n184, u0_u11_u1_n185, u0_u11_u1_n186, 
       u0_u11_u1_n187, u0_u11_u1_n188, u0_u11_u1_n95, u0_u11_u1_n96, u0_u11_u1_n97, u0_u11_u1_n98, u0_u11_u1_n99, u0_u11_u2_n100, u0_u11_u2_n101, 
       u0_u11_u2_n102, u0_u11_u2_n103, u0_u11_u2_n104, u0_u11_u2_n105, u0_u11_u2_n106, u0_u11_u2_n107, u0_u11_u2_n108, u0_u11_u2_n109, u0_u11_u2_n110, 
       u0_u11_u2_n111, u0_u11_u2_n112, u0_u11_u2_n113, u0_u11_u2_n114, u0_u11_u2_n115, u0_u11_u2_n116, u0_u11_u2_n117, u0_u11_u2_n118, u0_u11_u2_n119, 
       u0_u11_u2_n120, u0_u11_u2_n121, u0_u11_u2_n122, u0_u11_u2_n123, u0_u11_u2_n124, u0_u11_u2_n125, u0_u11_u2_n126, u0_u11_u2_n127, u0_u11_u2_n128, 
       u0_u11_u2_n129, u0_u11_u2_n130, u0_u11_u2_n131, u0_u11_u2_n132, u0_u11_u2_n133, u0_u11_u2_n134, u0_u11_u2_n135, u0_u11_u2_n136, u0_u11_u2_n137, 
       u0_u11_u2_n138, u0_u11_u2_n139, u0_u11_u2_n140, u0_u11_u2_n141, u0_u11_u2_n142, u0_u11_u2_n143, u0_u11_u2_n144, u0_u11_u2_n145, u0_u11_u2_n146, 
       u0_u11_u2_n147, u0_u11_u2_n148, u0_u11_u2_n149, u0_u11_u2_n150, u0_u11_u2_n151, u0_u11_u2_n152, u0_u11_u2_n153, u0_u11_u2_n154, u0_u11_u2_n155, 
       u0_u11_u2_n156, u0_u11_u2_n157, u0_u11_u2_n158, u0_u11_u2_n159, u0_u11_u2_n160, u0_u11_u2_n161, u0_u11_u2_n162, u0_u11_u2_n163, u0_u11_u2_n164, 
       u0_u11_u2_n165, u0_u11_u2_n166, u0_u11_u2_n167, u0_u11_u2_n168, u0_u11_u2_n169, u0_u11_u2_n170, u0_u11_u2_n171, u0_u11_u2_n172, u0_u11_u2_n173, 
       u0_u11_u2_n174, u0_u11_u2_n175, u0_u11_u2_n176, u0_u11_u2_n177, u0_u11_u2_n178, u0_u11_u2_n179, u0_u11_u2_n180, u0_u11_u2_n181, u0_u11_u2_n182, 
       u0_u11_u2_n183, u0_u11_u2_n184, u0_u11_u2_n185, u0_u11_u2_n186, u0_u11_u2_n187, u0_u11_u2_n188, u0_u11_u2_n95, u0_u11_u2_n96, u0_u11_u2_n97, 
       u0_u11_u2_n98, u0_u11_u2_n99, u0_u11_u3_n100, u0_u11_u3_n101, u0_u11_u3_n102, u0_u11_u3_n103, u0_u11_u3_n104, u0_u11_u3_n105, u0_u11_u3_n106, 
       u0_u11_u3_n107, u0_u11_u3_n108, u0_u11_u3_n109, u0_u11_u3_n110, u0_u11_u3_n111, u0_u11_u3_n112, u0_u11_u3_n113, u0_u11_u3_n114, u0_u11_u3_n115, 
       u0_u11_u3_n116, u0_u11_u3_n117, u0_u11_u3_n118, u0_u11_u3_n119, u0_u11_u3_n120, u0_u11_u3_n121, u0_u11_u3_n122, u0_u11_u3_n123, u0_u11_u3_n124, 
       u0_u11_u3_n125, u0_u11_u3_n126, u0_u11_u3_n127, u0_u11_u3_n128, u0_u11_u3_n129, u0_u11_u3_n130, u0_u11_u3_n131, u0_u11_u3_n132, u0_u11_u3_n133, 
       u0_u11_u3_n134, u0_u11_u3_n135, u0_u11_u3_n136, u0_u11_u3_n137, u0_u11_u3_n138, u0_u11_u3_n139, u0_u11_u3_n140, u0_u11_u3_n141, u0_u11_u3_n142, 
       u0_u11_u3_n143, u0_u11_u3_n144, u0_u11_u3_n145, u0_u11_u3_n146, u0_u11_u3_n147, u0_u11_u3_n148, u0_u11_u3_n149, u0_u11_u3_n150, u0_u11_u3_n151, 
       u0_u11_u3_n152, u0_u11_u3_n153, u0_u11_u3_n154, u0_u11_u3_n155, u0_u11_u3_n156, u0_u11_u3_n157, u0_u11_u3_n158, u0_u11_u3_n159, u0_u11_u3_n160, 
       u0_u11_u3_n161, u0_u11_u3_n162, u0_u11_u3_n163, u0_u11_u3_n164, u0_u11_u3_n165, u0_u11_u3_n166, u0_u11_u3_n167, u0_u11_u3_n168, u0_u11_u3_n169, 
       u0_u11_u3_n170, u0_u11_u3_n171, u0_u11_u3_n172, u0_u11_u3_n173, u0_u11_u3_n174, u0_u11_u3_n175, u0_u11_u3_n176, u0_u11_u3_n177, u0_u11_u3_n178, 
       u0_u11_u3_n179, u0_u11_u3_n180, u0_u11_u3_n181, u0_u11_u3_n182, u0_u11_u3_n183, u0_u11_u3_n184, u0_u11_u3_n185, u0_u11_u3_n186, u0_u11_u3_n94, 
       u0_u11_u3_n95, u0_u11_u3_n96, u0_u11_u3_n97, u0_u11_u3_n98, u0_u11_u3_n99, u0_u15_X_13, u0_u15_X_14, u0_u15_X_15, u0_u15_X_16, 
       u0_u15_X_17, u0_u15_X_18, u0_u15_X_19, u0_u15_X_20, u0_u15_X_21, u0_u15_X_22, u0_u15_X_23, u0_u15_X_24, u0_u15_X_43, 
       u0_u15_X_44, u0_u15_X_45, u0_u15_X_46, u0_u15_X_47, u0_u15_X_48, u0_u15_u2_n100, u0_u15_u2_n101, u0_u15_u2_n102, u0_u15_u2_n103, 
       u0_u15_u2_n104, u0_u15_u2_n105, u0_u15_u2_n106, u0_u15_u2_n107, u0_u15_u2_n108, u0_u15_u2_n109, u0_u15_u2_n110, u0_u15_u2_n111, u0_u15_u2_n112, 
       u0_u15_u2_n113, u0_u15_u2_n114, u0_u15_u2_n115, u0_u15_u2_n116, u0_u15_u2_n117, u0_u15_u2_n118, u0_u15_u2_n119, u0_u15_u2_n120, u0_u15_u2_n121, 
       u0_u15_u2_n122, u0_u15_u2_n123, u0_u15_u2_n124, u0_u15_u2_n125, u0_u15_u2_n126, u0_u15_u2_n127, u0_u15_u2_n128, u0_u15_u2_n129, u0_u15_u2_n130, 
       u0_u15_u2_n131, u0_u15_u2_n132, u0_u15_u2_n133, u0_u15_u2_n134, u0_u15_u2_n135, u0_u15_u2_n136, u0_u15_u2_n137, u0_u15_u2_n138, u0_u15_u2_n139, 
       u0_u15_u2_n140, u0_u15_u2_n141, u0_u15_u2_n142, u0_u15_u2_n143, u0_u15_u2_n144, u0_u15_u2_n145, u0_u15_u2_n146, u0_u15_u2_n147, u0_u15_u2_n148, 
       u0_u15_u2_n149, u0_u15_u2_n150, u0_u15_u2_n151, u0_u15_u2_n152, u0_u15_u2_n153, u0_u15_u2_n154, u0_u15_u2_n155, u0_u15_u2_n156, u0_u15_u2_n157, 
       u0_u15_u2_n158, u0_u15_u2_n159, u0_u15_u2_n160, u0_u15_u2_n161, u0_u15_u2_n162, u0_u15_u2_n163, u0_u15_u2_n164, u0_u15_u2_n165, u0_u15_u2_n166, 
       u0_u15_u2_n167, u0_u15_u2_n168, u0_u15_u2_n169, u0_u15_u2_n170, u0_u15_u2_n171, u0_u15_u2_n172, u0_u15_u2_n173, u0_u15_u2_n174, u0_u15_u2_n175, 
       u0_u15_u2_n176, u0_u15_u2_n177, u0_u15_u2_n178, u0_u15_u2_n179, u0_u15_u2_n180, u0_u15_u2_n181, u0_u15_u2_n182, u0_u15_u2_n183, u0_u15_u2_n184, 
       u0_u15_u2_n185, u0_u15_u2_n186, u0_u15_u2_n187, u0_u15_u2_n188, u0_u15_u2_n95, u0_u15_u2_n96, u0_u15_u2_n97, u0_u15_u2_n98, u0_u15_u2_n99, 
       u0_u15_u3_n100, u0_u15_u3_n101, u0_u15_u3_n102, u0_u15_u3_n103, u0_u15_u3_n104, u0_u15_u3_n105, u0_u15_u3_n106, u0_u15_u3_n107, u0_u15_u3_n108, 
       u0_u15_u3_n109, u0_u15_u3_n110, u0_u15_u3_n111, u0_u15_u3_n112, u0_u15_u3_n113, u0_u15_u3_n114, u0_u15_u3_n115, u0_u15_u3_n116, u0_u15_u3_n117, 
       u0_u15_u3_n118, u0_u15_u3_n119, u0_u15_u3_n120, u0_u15_u3_n121, u0_u15_u3_n122, u0_u15_u3_n123, u0_u15_u3_n124, u0_u15_u3_n125, u0_u15_u3_n126, 
       u0_u15_u3_n127, u0_u15_u3_n128, u0_u15_u3_n129, u0_u15_u3_n130, u0_u15_u3_n131, u0_u15_u3_n132, u0_u15_u3_n133, u0_u15_u3_n134, u0_u15_u3_n135, 
       u0_u15_u3_n136, u0_u15_u3_n137, u0_u15_u3_n138, u0_u15_u3_n139, u0_u15_u3_n140, u0_u15_u3_n141, u0_u15_u3_n142, u0_u15_u3_n143, u0_u15_u3_n144, 
       u0_u15_u3_n145, u0_u15_u3_n146, u0_u15_u3_n147, u0_u15_u3_n148, u0_u15_u3_n149, u0_u15_u3_n150, u0_u15_u3_n151, u0_u15_u3_n152, u0_u15_u3_n153, 
       u0_u15_u3_n154, u0_u15_u3_n155, u0_u15_u3_n156, u0_u15_u3_n157, u0_u15_u3_n158, u0_u15_u3_n159, u0_u15_u3_n160, u0_u15_u3_n161, u0_u15_u3_n162, 
       u0_u15_u3_n163, u0_u15_u3_n164, u0_u15_u3_n165, u0_u15_u3_n166, u0_u15_u3_n167, u0_u15_u3_n168, u0_u15_u3_n169, u0_u15_u3_n170, u0_u15_u3_n171, 
       u0_u15_u3_n172, u0_u15_u3_n173, u0_u15_u3_n174, u0_u15_u3_n175, u0_u15_u3_n176, u0_u15_u3_n177, u0_u15_u3_n178, u0_u15_u3_n179, u0_u15_u3_n180, 
       u0_u15_u3_n181, u0_u15_u3_n182, u0_u15_u3_n183, u0_u15_u3_n184, u0_u15_u3_n185, u0_u15_u3_n186, u0_u15_u3_n94, u0_u15_u3_n95, u0_u15_u3_n96, 
       u0_u15_u3_n97, u0_u15_u3_n98, u0_u15_u3_n99, u0_u15_u7_n100, u0_u15_u7_n101, u0_u15_u7_n102, u0_u15_u7_n103, u0_u15_u7_n104, u0_u15_u7_n105, 
       u0_u15_u7_n106, u0_u15_u7_n107, u0_u15_u7_n108, u0_u15_u7_n109, u0_u15_u7_n110, u0_u15_u7_n111, u0_u15_u7_n112, u0_u15_u7_n113, u0_u15_u7_n114, 
       u0_u15_u7_n115, u0_u15_u7_n116, u0_u15_u7_n117, u0_u15_u7_n118, u0_u15_u7_n119, u0_u15_u7_n120, u0_u15_u7_n121, u0_u15_u7_n122, u0_u15_u7_n123, 
       u0_u15_u7_n124, u0_u15_u7_n125, u0_u15_u7_n126, u0_u15_u7_n127, u0_u15_u7_n128, u0_u15_u7_n129, u0_u15_u7_n130, u0_u15_u7_n131, u0_u15_u7_n132, 
       u0_u15_u7_n133, u0_u15_u7_n134, u0_u15_u7_n135, u0_u15_u7_n136, u0_u15_u7_n137, u0_u15_u7_n138, u0_u15_u7_n139, u0_u15_u7_n140, u0_u15_u7_n141, 
       u0_u15_u7_n142, u0_u15_u7_n143, u0_u15_u7_n144, u0_u15_u7_n145, u0_u15_u7_n146, u0_u15_u7_n147, u0_u15_u7_n148, u0_u15_u7_n149, u0_u15_u7_n150, 
       u0_u15_u7_n151, u0_u15_u7_n152, u0_u15_u7_n153, u0_u15_u7_n154, u0_u15_u7_n155, u0_u15_u7_n156, u0_u15_u7_n157, u0_u15_u7_n158, u0_u15_u7_n159, 
       u0_u15_u7_n160, u0_u15_u7_n161, u0_u15_u7_n162, u0_u15_u7_n163, u0_u15_u7_n164, u0_u15_u7_n165, u0_u15_u7_n166, u0_u15_u7_n167, u0_u15_u7_n168, 
       u0_u15_u7_n169, u0_u15_u7_n170, u0_u15_u7_n171, u0_u15_u7_n172, u0_u15_u7_n173, u0_u15_u7_n174, u0_u15_u7_n175, u0_u15_u7_n176, u0_u15_u7_n177, 
       u0_u15_u7_n178, u0_u15_u7_n179, u0_u15_u7_n180, u0_u15_u7_n91, u0_u15_u7_n92, u0_u15_u7_n93, u0_u15_u7_n94, u0_u15_u7_n95, u0_u15_u7_n96, 
       u0_u15_u7_n97, u0_u15_u7_n98, u0_u15_u7_n99, u0_u4_X_25, u0_u4_X_26, u0_u4_X_27, u0_u4_X_28, u0_u4_X_29, u0_u4_X_30, 
       u0_u4_X_31, u0_u4_X_32, u0_u4_X_33, u0_u4_X_34, u0_u4_X_35, u0_u4_X_36, u0_u4_X_37, u0_u4_X_38, u0_u4_X_39, 
       u0_u4_X_40, u0_u4_X_41, u0_u4_X_42, u0_u4_u4_n100, u0_u4_u4_n101, u0_u4_u4_n102, u0_u4_u4_n103, u0_u4_u4_n104, u0_u4_u4_n105, 
       u0_u4_u4_n106, u0_u4_u4_n107, u0_u4_u4_n108, u0_u4_u4_n109, u0_u4_u4_n110, u0_u4_u4_n111, u0_u4_u4_n112, u0_u4_u4_n113, u0_u4_u4_n114, 
       u0_u4_u4_n115, u0_u4_u4_n116, u0_u4_u4_n117, u0_u4_u4_n118, u0_u4_u4_n119, u0_u4_u4_n120, u0_u4_u4_n121, u0_u4_u4_n122, u0_u4_u4_n123, 
       u0_u4_u4_n124, u0_u4_u4_n125, u0_u4_u4_n126, u0_u4_u4_n127, u0_u4_u4_n128, u0_u4_u4_n129, u0_u4_u4_n130, u0_u4_u4_n131, u0_u4_u4_n132, 
       u0_u4_u4_n133, u0_u4_u4_n134, u0_u4_u4_n135, u0_u4_u4_n136, u0_u4_u4_n137, u0_u4_u4_n138, u0_u4_u4_n139, u0_u4_u4_n140, u0_u4_u4_n141, 
       u0_u4_u4_n142, u0_u4_u4_n143, u0_u4_u4_n144, u0_u4_u4_n145, u0_u4_u4_n146, u0_u4_u4_n147, u0_u4_u4_n148, u0_u4_u4_n149, u0_u4_u4_n150, 
       u0_u4_u4_n151, u0_u4_u4_n152, u0_u4_u4_n153, u0_u4_u4_n154, u0_u4_u4_n155, u0_u4_u4_n156, u0_u4_u4_n157, u0_u4_u4_n158, u0_u4_u4_n159, 
       u0_u4_u4_n160, u0_u4_u4_n161, u0_u4_u4_n162, u0_u4_u4_n163, u0_u4_u4_n164, u0_u4_u4_n165, u0_u4_u4_n166, u0_u4_u4_n167, u0_u4_u4_n168, 
       u0_u4_u4_n169, u0_u4_u4_n170, u0_u4_u4_n171, u0_u4_u4_n172, u0_u4_u4_n173, u0_u4_u4_n174, u0_u4_u4_n175, u0_u4_u4_n176, u0_u4_u4_n177, 
       u0_u4_u4_n178, u0_u4_u4_n179, u0_u4_u4_n180, u0_u4_u4_n181, u0_u4_u4_n182, u0_u4_u4_n183, u0_u4_u4_n184, u0_u4_u4_n185, u0_u4_u4_n186, 
       u0_u4_u4_n94, u0_u4_u4_n95, u0_u4_u4_n96, u0_u4_u4_n97, u0_u4_u4_n98, u0_u4_u4_n99, u0_u4_u5_n100, u0_u4_u5_n101, u0_u4_u5_n102, 
       u0_u4_u5_n103, u0_u4_u5_n104, u0_u4_u5_n105, u0_u4_u5_n106, u0_u4_u5_n107, u0_u4_u5_n108, u0_u4_u5_n109, u0_u4_u5_n110, u0_u4_u5_n111, 
       u0_u4_u5_n112, u0_u4_u5_n113, u0_u4_u5_n114, u0_u4_u5_n115, u0_u4_u5_n116, u0_u4_u5_n117, u0_u4_u5_n118, u0_u4_u5_n119, u0_u4_u5_n120, 
       u0_u4_u5_n121, u0_u4_u5_n122, u0_u4_u5_n123, u0_u4_u5_n124, u0_u4_u5_n125, u0_u4_u5_n126, u0_u4_u5_n127, u0_u4_u5_n128, u0_u4_u5_n129, 
       u0_u4_u5_n130, u0_u4_u5_n131, u0_u4_u5_n132, u0_u4_u5_n133, u0_u4_u5_n134, u0_u4_u5_n135, u0_u4_u5_n136, u0_u4_u5_n137, u0_u4_u5_n138, 
       u0_u4_u5_n139, u0_u4_u5_n140, u0_u4_u5_n141, u0_u4_u5_n142, u0_u4_u5_n143, u0_u4_u5_n144, u0_u4_u5_n145, u0_u4_u5_n146, u0_u4_u5_n147, 
       u0_u4_u5_n148, u0_u4_u5_n149, u0_u4_u5_n150, u0_u4_u5_n151, u0_u4_u5_n152, u0_u4_u5_n153, u0_u4_u5_n154, u0_u4_u5_n155, u0_u4_u5_n156, 
       u0_u4_u5_n157, u0_u4_u5_n158, u0_u4_u5_n159, u0_u4_u5_n160, u0_u4_u5_n161, u0_u4_u5_n162, u0_u4_u5_n163, u0_u4_u5_n164, u0_u4_u5_n165, 
       u0_u4_u5_n166, u0_u4_u5_n167, u0_u4_u5_n168, u0_u4_u5_n169, u0_u4_u5_n170, u0_u4_u5_n171, u0_u4_u5_n172, u0_u4_u5_n173, u0_u4_u5_n174, 
       u0_u4_u5_n175, u0_u4_u5_n176, u0_u4_u5_n177, u0_u4_u5_n178, u0_u4_u5_n179, u0_u4_u5_n180, u0_u4_u5_n181, u0_u4_u5_n182, u0_u4_u5_n183, 
       u0_u4_u5_n184, u0_u4_u5_n185, u0_u4_u5_n186, u0_u4_u5_n187, u0_u4_u5_n188, u0_u4_u5_n189, u0_u4_u5_n190, u0_u4_u5_n191, u0_u4_u5_n192, 
       u0_u4_u5_n193, u0_u4_u5_n194, u0_u4_u5_n195, u0_u4_u5_n196, u0_u4_u5_n99, u0_u4_u6_n100, u0_u4_u6_n101, u0_u4_u6_n102, u0_u4_u6_n103, 
       u0_u4_u6_n104, u0_u4_u6_n105, u0_u4_u6_n106, u0_u4_u6_n107, u0_u4_u6_n108, u0_u4_u6_n109, u0_u4_u6_n110, u0_u4_u6_n111, u0_u4_u6_n112, 
       u0_u4_u6_n113, u0_u4_u6_n114, u0_u4_u6_n115, u0_u4_u6_n116, u0_u4_u6_n117, u0_u4_u6_n118, u0_u4_u6_n119, u0_u4_u6_n120, u0_u4_u6_n121, 
       u0_u4_u6_n122, u0_u4_u6_n123, u0_u4_u6_n124, u0_u4_u6_n125, u0_u4_u6_n126, u0_u4_u6_n127, u0_u4_u6_n128, u0_u4_u6_n129, u0_u4_u6_n130, 
       u0_u4_u6_n131, u0_u4_u6_n132, u0_u4_u6_n133, u0_u4_u6_n134, u0_u4_u6_n135, u0_u4_u6_n136, u0_u4_u6_n137, u0_u4_u6_n138, u0_u4_u6_n139, 
       u0_u4_u6_n140, u0_u4_u6_n141, u0_u4_u6_n142, u0_u4_u6_n143, u0_u4_u6_n144, u0_u4_u6_n145, u0_u4_u6_n146, u0_u4_u6_n147, u0_u4_u6_n148, 
       u0_u4_u6_n149, u0_u4_u6_n150, u0_u4_u6_n151, u0_u4_u6_n152, u0_u4_u6_n153, u0_u4_u6_n154, u0_u4_u6_n155, u0_u4_u6_n156, u0_u4_u6_n157, 
       u0_u4_u6_n158, u0_u4_u6_n159, u0_u4_u6_n160, u0_u4_u6_n161, u0_u4_u6_n162, u0_u4_u6_n163, u0_u4_u6_n164, u0_u4_u6_n165, u0_u4_u6_n166, 
       u0_u4_u6_n167, u0_u4_u6_n168, u0_u4_u6_n169, u0_u4_u6_n170, u0_u4_u6_n171, u0_u4_u6_n172, u0_u4_u6_n173, u0_u4_u6_n174, u0_u4_u6_n88, 
       u0_u4_u6_n89, u0_u4_u6_n90, u0_u4_u6_n91, u0_u4_u6_n92, u0_u4_u6_n93, u0_u4_u6_n94, u0_u4_u6_n95, u0_u4_u6_n96, u0_u4_u6_n97, 
       u0_u4_u6_n98, u0_u4_u6_n99, u0_uk_n693, u0_uk_n700, u0_uk_n701, u0_uk_n706, u0_uk_n709, u0_uk_n710, u0_uk_n714, 
       u0_uk_n716, u0_uk_n807, u0_uk_n808, u0_uk_n809, u0_uk_n811, u0_uk_n814, u0_uk_n870, u0_uk_n872, u0_uk_n873, 
       u0_uk_n874, u0_uk_n876, u0_uk_n877, u0_uk_n879, u0_uk_n882, u0_uk_n883, u0_uk_n884, u0_uk_n895, u0_uk_n896, 
       u0_uk_n907, u0_uk_n908, u0_uk_n909, u0_uk_n962, u0_uk_n968, u0_uk_n975, u0_uk_n976, u0_uk_n977, u0_uk_n978, 
       u0_uk_n979, u0_uk_n980, u2_K11_25, u2_K11_26, u2_K11_27, u2_K11_28, u2_K11_30, u2_K13_1, u2_K13_10, 
       u2_K13_11, u2_K13_12, u2_K13_13, u2_K13_15, u2_K13_16, u2_K13_17, u2_K13_18, u2_K13_2, u2_K13_38, 
       u2_K13_39, u2_K13_4, u2_K13_41, u2_K13_43, u2_K13_48, u2_K13_5, u2_K13_6, u2_K13_7, u2_K13_9, 
       u2_K4_1, u2_K4_10, u2_K4_11, u2_K4_12, u2_K4_2, u2_K4_3, u2_K4_4, u2_K4_43, u2_K4_44, 
       u2_K4_45, u2_K4_46, u2_K4_47, u2_K4_48, u2_K4_5, u2_K4_8, u2_K4_9, u2_K6_26, u2_K6_28, 
       u2_K6_29, u2_K6_30, u2_K8_19, u2_K8_20, u2_K8_21, u2_K8_22, u2_K8_23, u2_K8_25, u2_K8_27, 
       u2_K8_28, u2_K8_29, u2_K8_30, u2_K8_32, u2_K8_33, u2_K8_34, u2_K8_35, u2_K8_36, u2_K8_37, 
       u2_K8_38, u2_K8_39, u2_K8_40, u2_K8_42, u2_out10_14, u2_out10_25, u2_out10_3, u2_out10_8, u2_out12_12, 
       u2_out12_13, u2_out12_15, u2_out12_16, u2_out12_17, u2_out12_18, u2_out12_2, u2_out12_21, u2_out12_22, u2_out12_23, 
       u2_out12_24, u2_out12_27, u2_out12_28, u2_out12_30, u2_out12_31, u2_out12_32, u2_out12_5, u2_out12_6, u2_out12_7, 
       u2_out12_9, u2_out3_13, u2_out3_15, u2_out3_17, u2_out3_18, u2_out3_2, u2_out3_21, u2_out3_23, u2_out3_27, 
       u2_out3_28, u2_out3_31, u2_out3_5, u2_out3_9, u2_out5_14, u2_out5_25, u2_out5_3, u2_out5_8, u2_out7_1, 
       u2_out7_10, u2_out7_11, u2_out7_12, u2_out7_14, u2_out7_19, u2_out7_20, u2_out7_22, u2_out7_25, u2_out7_26, 
       u2_out7_29, u2_out7_3, u2_out7_32, u2_out7_4, u2_out7_7, u2_out7_8, u2_u10_X_25, u2_u10_X_26, u2_u10_X_27, 
       u2_u10_X_28, u2_u10_X_29, u2_u10_X_30, u2_u10_u4_n100, u2_u10_u4_n101, u2_u10_u4_n102, u2_u10_u4_n103, u2_u10_u4_n104, u2_u10_u4_n105, 
       u2_u10_u4_n106, u2_u10_u4_n107, u2_u10_u4_n108, u2_u10_u4_n109, u2_u10_u4_n110, u2_u10_u4_n111, u2_u10_u4_n112, u2_u10_u4_n113, u2_u10_u4_n114, 
       u2_u10_u4_n115, u2_u10_u4_n116, u2_u10_u4_n117, u2_u10_u4_n118, u2_u10_u4_n119, u2_u10_u4_n120, u2_u10_u4_n121, u2_u10_u4_n122, u2_u10_u4_n123, 
       u2_u10_u4_n124, u2_u10_u4_n125, u2_u10_u4_n126, u2_u10_u4_n127, u2_u10_u4_n128, u2_u10_u4_n129, u2_u10_u4_n130, u2_u10_u4_n131, u2_u10_u4_n132, 
       u2_u10_u4_n133, u2_u10_u4_n134, u2_u10_u4_n135, u2_u10_u4_n136, u2_u10_u4_n137, u2_u10_u4_n138, u2_u10_u4_n139, u2_u10_u4_n140, u2_u10_u4_n141, 
       u2_u10_u4_n142, u2_u10_u4_n143, u2_u10_u4_n144, u2_u10_u4_n145, u2_u10_u4_n146, u2_u10_u4_n147, u2_u10_u4_n148, u2_u10_u4_n149, u2_u10_u4_n150, 
       u2_u10_u4_n151, u2_u10_u4_n152, u2_u10_u4_n153, u2_u10_u4_n154, u2_u10_u4_n155, u2_u10_u4_n156, u2_u10_u4_n157, u2_u10_u4_n158, u2_u10_u4_n159, 
       u2_u10_u4_n160, u2_u10_u4_n161, u2_u10_u4_n162, u2_u10_u4_n163, u2_u10_u4_n164, u2_u10_u4_n165, u2_u10_u4_n166, u2_u10_u4_n167, u2_u10_u4_n168, 
       u2_u10_u4_n169, u2_u10_u4_n170, u2_u10_u4_n171, u2_u10_u4_n172, u2_u10_u4_n173, u2_u10_u4_n174, u2_u10_u4_n175, u2_u10_u4_n176, u2_u10_u4_n177, 
       u2_u10_u4_n178, u2_u10_u4_n179, u2_u10_u4_n180, u2_u10_u4_n181, u2_u10_u4_n182, u2_u10_u4_n183, u2_u10_u4_n184, u2_u10_u4_n185, u2_u10_u4_n186, 
       u2_u10_u4_n94, u2_u10_u4_n95, u2_u10_u4_n96, u2_u10_u4_n97, u2_u10_u4_n98, u2_u10_u4_n99, u2_u12_X_1, u2_u12_X_10, u2_u12_X_11, 
       u2_u12_X_12, u2_u12_X_13, u2_u12_X_14, u2_u12_X_15, u2_u12_X_16, u2_u12_X_17, u2_u12_X_18, u2_u12_X_2, u2_u12_X_3, 
       u2_u12_X_37, u2_u12_X_38, u2_u12_X_39, u2_u12_X_4, u2_u12_X_40, u2_u12_X_41, u2_u12_X_42, u2_u12_X_43, u2_u12_X_44, 
       u2_u12_X_45, u2_u12_X_46, u2_u12_X_47, u2_u12_X_48, u2_u12_X_5, u2_u12_X_6, u2_u12_X_7, u2_u12_X_8, u2_u12_X_9, 
       u2_u12_u0_n100, u2_u12_u0_n101, u2_u12_u0_n102, u2_u12_u0_n103, u2_u12_u0_n104, u2_u12_u0_n105, u2_u12_u0_n106, u2_u12_u0_n107, u2_u12_u0_n108, 
       u2_u12_u0_n109, u2_u12_u0_n110, u2_u12_u0_n111, u2_u12_u0_n112, u2_u12_u0_n113, u2_u12_u0_n114, u2_u12_u0_n115, u2_u12_u0_n116, u2_u12_u0_n117, 
       u2_u12_u0_n118, u2_u12_u0_n119, u2_u12_u0_n120, u2_u12_u0_n121, u2_u12_u0_n122, u2_u12_u0_n123, u2_u12_u0_n124, u2_u12_u0_n125, u2_u12_u0_n126, 
       u2_u12_u0_n127, u2_u12_u0_n128, u2_u12_u0_n129, u2_u12_u0_n130, u2_u12_u0_n131, u2_u12_u0_n132, u2_u12_u0_n133, u2_u12_u0_n134, u2_u12_u0_n135, 
       u2_u12_u0_n136, u2_u12_u0_n137, u2_u12_u0_n138, u2_u12_u0_n139, u2_u12_u0_n140, u2_u12_u0_n141, u2_u12_u0_n142, u2_u12_u0_n143, u2_u12_u0_n144, 
       u2_u12_u0_n145, u2_u12_u0_n146, u2_u12_u0_n147, u2_u12_u0_n148, u2_u12_u0_n149, u2_u12_u0_n150, u2_u12_u0_n151, u2_u12_u0_n152, u2_u12_u0_n153, 
       u2_u12_u0_n154, u2_u12_u0_n155, u2_u12_u0_n156, u2_u12_u0_n157, u2_u12_u0_n158, u2_u12_u0_n159, u2_u12_u0_n160, u2_u12_u0_n161, u2_u12_u0_n162, 
       u2_u12_u0_n163, u2_u12_u0_n164, u2_u12_u0_n165, u2_u12_u0_n166, u2_u12_u0_n167, u2_u12_u0_n168, u2_u12_u0_n169, u2_u12_u0_n170, u2_u12_u0_n171, 
       u2_u12_u0_n172, u2_u12_u0_n173, u2_u12_u0_n174, u2_u12_u0_n88, u2_u12_u0_n89, u2_u12_u0_n90, u2_u12_u0_n91, u2_u12_u0_n92, u2_u12_u0_n93, 
       u2_u12_u0_n94, u2_u12_u0_n95, u2_u12_u0_n96, u2_u12_u0_n97, u2_u12_u0_n98, u2_u12_u0_n99, u2_u12_u1_n100, u2_u12_u1_n101, u2_u12_u1_n102, 
       u2_u12_u1_n103, u2_u12_u1_n104, u2_u12_u1_n105, u2_u12_u1_n106, u2_u12_u1_n107, u2_u12_u1_n108, u2_u12_u1_n109, u2_u12_u1_n110, u2_u12_u1_n111, 
       u2_u12_u1_n112, u2_u12_u1_n113, u2_u12_u1_n114, u2_u12_u1_n115, u2_u12_u1_n116, u2_u12_u1_n117, u2_u12_u1_n118, u2_u12_u1_n119, u2_u12_u1_n120, 
       u2_u12_u1_n121, u2_u12_u1_n122, u2_u12_u1_n123, u2_u12_u1_n124, u2_u12_u1_n125, u2_u12_u1_n126, u2_u12_u1_n127, u2_u12_u1_n128, u2_u12_u1_n129, 
       u2_u12_u1_n130, u2_u12_u1_n131, u2_u12_u1_n132, u2_u12_u1_n133, u2_u12_u1_n134, u2_u12_u1_n135, u2_u12_u1_n136, u2_u12_u1_n137, u2_u12_u1_n138, 
       u2_u12_u1_n139, u2_u12_u1_n140, u2_u12_u1_n141, u2_u12_u1_n142, u2_u12_u1_n143, u2_u12_u1_n144, u2_u12_u1_n145, u2_u12_u1_n146, u2_u12_u1_n147, 
       u2_u12_u1_n148, u2_u12_u1_n149, u2_u12_u1_n150, u2_u12_u1_n151, u2_u12_u1_n152, u2_u12_u1_n153, u2_u12_u1_n154, u2_u12_u1_n155, u2_u12_u1_n156, 
       u2_u12_u1_n157, u2_u12_u1_n158, u2_u12_u1_n159, u2_u12_u1_n160, u2_u12_u1_n161, u2_u12_u1_n162, u2_u12_u1_n163, u2_u12_u1_n164, u2_u12_u1_n165, 
       u2_u12_u1_n166, u2_u12_u1_n167, u2_u12_u1_n168, u2_u12_u1_n169, u2_u12_u1_n170, u2_u12_u1_n171, u2_u12_u1_n172, u2_u12_u1_n173, u2_u12_u1_n174, 
       u2_u12_u1_n175, u2_u12_u1_n176, u2_u12_u1_n177, u2_u12_u1_n178, u2_u12_u1_n179, u2_u12_u1_n180, u2_u12_u1_n181, u2_u12_u1_n182, u2_u12_u1_n183, 
       u2_u12_u1_n184, u2_u12_u1_n185, u2_u12_u1_n186, u2_u12_u1_n187, u2_u12_u1_n188, u2_u12_u1_n95, u2_u12_u1_n96, u2_u12_u1_n97, u2_u12_u1_n98, 
       u2_u12_u1_n99, u2_u12_u2_n100, u2_u12_u2_n101, u2_u12_u2_n102, u2_u12_u2_n103, u2_u12_u2_n104, u2_u12_u2_n105, u2_u12_u2_n106, u2_u12_u2_n107, 
       u2_u12_u2_n108, u2_u12_u2_n109, u2_u12_u2_n110, u2_u12_u2_n111, u2_u12_u2_n112, u2_u12_u2_n113, u2_u12_u2_n114, u2_u12_u2_n115, u2_u12_u2_n116, 
       u2_u12_u2_n117, u2_u12_u2_n118, u2_u12_u2_n119, u2_u12_u2_n120, u2_u12_u2_n121, u2_u12_u2_n122, u2_u12_u2_n123, u2_u12_u2_n124, u2_u12_u2_n125, 
       u2_u12_u2_n126, u2_u12_u2_n127, u2_u12_u2_n128, u2_u12_u2_n129, u2_u12_u2_n130, u2_u12_u2_n131, u2_u12_u2_n132, u2_u12_u2_n133, u2_u12_u2_n134, 
       u2_u12_u2_n135, u2_u12_u2_n136, u2_u12_u2_n137, u2_u12_u2_n138, u2_u12_u2_n139, u2_u12_u2_n140, u2_u12_u2_n141, u2_u12_u2_n142, u2_u12_u2_n143, 
       u2_u12_u2_n144, u2_u12_u2_n145, u2_u12_u2_n146, u2_u12_u2_n147, u2_u12_u2_n148, u2_u12_u2_n149, u2_u12_u2_n150, u2_u12_u2_n151, u2_u12_u2_n152, 
       u2_u12_u2_n153, u2_u12_u2_n154, u2_u12_u2_n155, u2_u12_u2_n156, u2_u12_u2_n157, u2_u12_u2_n158, u2_u12_u2_n159, u2_u12_u2_n160, u2_u12_u2_n161, 
       u2_u12_u2_n162, u2_u12_u2_n163, u2_u12_u2_n164, u2_u12_u2_n165, u2_u12_u2_n166, u2_u12_u2_n167, u2_u12_u2_n168, u2_u12_u2_n169, u2_u12_u2_n170, 
       u2_u12_u2_n171, u2_u12_u2_n172, u2_u12_u2_n173, u2_u12_u2_n174, u2_u12_u2_n175, u2_u12_u2_n176, u2_u12_u2_n177, u2_u12_u2_n178, u2_u12_u2_n179, 
       u2_u12_u2_n180, u2_u12_u2_n181, u2_u12_u2_n182, u2_u12_u2_n183, u2_u12_u2_n184, u2_u12_u2_n185, u2_u12_u2_n186, u2_u12_u2_n187, u2_u12_u2_n188, 
       u2_u12_u2_n95, u2_u12_u2_n96, u2_u12_u2_n97, u2_u12_u2_n98, u2_u12_u2_n99, u2_u12_u6_n100, u2_u12_u6_n101, u2_u12_u6_n102, u2_u12_u6_n103, 
       u2_u12_u6_n104, u2_u12_u6_n105, u2_u12_u6_n106, u2_u12_u6_n107, u2_u12_u6_n108, u2_u12_u6_n109, u2_u12_u6_n110, u2_u12_u6_n111, u2_u12_u6_n112, 
       u2_u12_u6_n113, u2_u12_u6_n114, u2_u12_u6_n115, u2_u12_u6_n116, u2_u12_u6_n117, u2_u12_u6_n118, u2_u12_u6_n119, u2_u12_u6_n120, u2_u12_u6_n121, 
       u2_u12_u6_n122, u2_u12_u6_n123, u2_u12_u6_n124, u2_u12_u6_n125, u2_u12_u6_n126, u2_u12_u6_n127, u2_u12_u6_n128, u2_u12_u6_n129, u2_u12_u6_n130, 
       u2_u12_u6_n131, u2_u12_u6_n132, u2_u12_u6_n133, u2_u12_u6_n134, u2_u12_u6_n135, u2_u12_u6_n136, u2_u12_u6_n137, u2_u12_u6_n138, u2_u12_u6_n139, 
       u2_u12_u6_n140, u2_u12_u6_n141, u2_u12_u6_n142, u2_u12_u6_n143, u2_u12_u6_n144, u2_u12_u6_n145, u2_u12_u6_n146, u2_u12_u6_n147, u2_u12_u6_n148, 
       u2_u12_u6_n149, u2_u12_u6_n150, u2_u12_u6_n151, u2_u12_u6_n152, u2_u12_u6_n153, u2_u12_u6_n154, u2_u12_u6_n155, u2_u12_u6_n156, u2_u12_u6_n157, 
       u2_u12_u6_n158, u2_u12_u6_n159, u2_u12_u6_n160, u2_u12_u6_n161, u2_u12_u6_n162, u2_u12_u6_n163, u2_u12_u6_n164, u2_u12_u6_n165, u2_u12_u6_n166, 
       u2_u12_u6_n167, u2_u12_u6_n168, u2_u12_u6_n169, u2_u12_u6_n170, u2_u12_u6_n171, u2_u12_u6_n172, u2_u12_u6_n173, u2_u12_u6_n174, u2_u12_u6_n88, 
       u2_u12_u6_n89, u2_u12_u6_n90, u2_u12_u6_n91, u2_u12_u6_n92, u2_u12_u6_n93, u2_u12_u6_n94, u2_u12_u6_n95, u2_u12_u6_n96, u2_u12_u6_n97, 
       u2_u12_u6_n98, u2_u12_u6_n99, u2_u12_u7_n100, u2_u12_u7_n101, u2_u12_u7_n102, u2_u12_u7_n103, u2_u12_u7_n104, u2_u12_u7_n105, u2_u12_u7_n106, 
       u2_u12_u7_n107, u2_u12_u7_n108, u2_u12_u7_n109, u2_u12_u7_n110, u2_u12_u7_n111, u2_u12_u7_n112, u2_u12_u7_n113, u2_u12_u7_n114, u2_u12_u7_n115, 
       u2_u12_u7_n116, u2_u12_u7_n117, u2_u12_u7_n118, u2_u12_u7_n119, u2_u12_u7_n120, u2_u12_u7_n121, u2_u12_u7_n122, u2_u12_u7_n123, u2_u12_u7_n124, 
       u2_u12_u7_n125, u2_u12_u7_n126, u2_u12_u7_n127, u2_u12_u7_n128, u2_u12_u7_n129, u2_u12_u7_n130, u2_u12_u7_n131, u2_u12_u7_n132, u2_u12_u7_n133, 
       u2_u12_u7_n134, u2_u12_u7_n135, u2_u12_u7_n136, u2_u12_u7_n137, u2_u12_u7_n138, u2_u12_u7_n139, u2_u12_u7_n140, u2_u12_u7_n141, u2_u12_u7_n142, 
       u2_u12_u7_n143, u2_u12_u7_n144, u2_u12_u7_n145, u2_u12_u7_n146, u2_u12_u7_n147, u2_u12_u7_n148, u2_u12_u7_n149, u2_u12_u7_n150, u2_u12_u7_n151, 
       u2_u12_u7_n152, u2_u12_u7_n153, u2_u12_u7_n154, u2_u12_u7_n155, u2_u12_u7_n156, u2_u12_u7_n157, u2_u12_u7_n158, u2_u12_u7_n159, u2_u12_u7_n160, 
       u2_u12_u7_n161, u2_u12_u7_n162, u2_u12_u7_n163, u2_u12_u7_n164, u2_u12_u7_n165, u2_u12_u7_n166, u2_u12_u7_n167, u2_u12_u7_n168, u2_u12_u7_n169, 
       u2_u12_u7_n170, u2_u12_u7_n171, u2_u12_u7_n172, u2_u12_u7_n173, u2_u12_u7_n174, u2_u12_u7_n175, u2_u12_u7_n176, u2_u12_u7_n177, u2_u12_u7_n178, 
       u2_u12_u7_n179, u2_u12_u7_n180, u2_u12_u7_n91, u2_u12_u7_n92, u2_u12_u7_n93, u2_u12_u7_n94, u2_u12_u7_n95, u2_u12_u7_n96, u2_u12_u7_n97, 
       u2_u12_u7_n98, u2_u12_u7_n99, u2_u3_X_1, u2_u3_X_10, u2_u3_X_11, u2_u3_X_12, u2_u3_X_2, u2_u3_X_3, u2_u3_X_4, 
       u2_u3_X_43, u2_u3_X_44, u2_u3_X_45, u2_u3_X_46, u2_u3_X_47, u2_u3_X_48, u2_u3_X_5, u2_u3_X_6, u2_u3_X_7, 
       u2_u3_X_8, u2_u3_X_9, u2_u3_u0_n100, u2_u3_u0_n101, u2_u3_u0_n102, u2_u3_u0_n103, u2_u3_u0_n104, u2_u3_u0_n105, u2_u3_u0_n106, 
       u2_u3_u0_n107, u2_u3_u0_n108, u2_u3_u0_n109, u2_u3_u0_n110, u2_u3_u0_n111, u2_u3_u0_n112, u2_u3_u0_n113, u2_u3_u0_n114, u2_u3_u0_n115, 
       u2_u3_u0_n116, u2_u3_u0_n117, u2_u3_u0_n118, u2_u3_u0_n119, u2_u3_u0_n120, u2_u3_u0_n121, u2_u3_u0_n122, u2_u3_u0_n123, u2_u3_u0_n124, 
       u2_u3_u0_n125, u2_u3_u0_n126, u2_u3_u0_n127, u2_u3_u0_n128, u2_u3_u0_n129, u2_u3_u0_n130, u2_u3_u0_n131, u2_u3_u0_n132, u2_u3_u0_n133, 
       u2_u3_u0_n134, u2_u3_u0_n135, u2_u3_u0_n136, u2_u3_u0_n137, u2_u3_u0_n138, u2_u3_u0_n139, u2_u3_u0_n140, u2_u3_u0_n141, u2_u3_u0_n142, 
       u2_u3_u0_n143, u2_u3_u0_n144, u2_u3_u0_n145, u2_u3_u0_n146, u2_u3_u0_n147, u2_u3_u0_n148, u2_u3_u0_n149, u2_u3_u0_n150, u2_u3_u0_n151, 
       u2_u3_u0_n152, u2_u3_u0_n153, u2_u3_u0_n154, u2_u3_u0_n155, u2_u3_u0_n156, u2_u3_u0_n157, u2_u3_u0_n158, u2_u3_u0_n159, u2_u3_u0_n160, 
       u2_u3_u0_n161, u2_u3_u0_n162, u2_u3_u0_n163, u2_u3_u0_n164, u2_u3_u0_n165, u2_u3_u0_n166, u2_u3_u0_n167, u2_u3_u0_n168, u2_u3_u0_n169, 
       u2_u3_u0_n170, u2_u3_u0_n171, u2_u3_u0_n172, u2_u3_u0_n173, u2_u3_u0_n174, u2_u3_u0_n88, u2_u3_u0_n89, u2_u3_u0_n90, u2_u3_u0_n91, 
       u2_u3_u0_n92, u2_u3_u0_n93, u2_u3_u0_n94, u2_u3_u0_n95, u2_u3_u0_n96, u2_u3_u0_n97, u2_u3_u0_n98, u2_u3_u0_n99, u2_u3_u1_n100, 
       u2_u3_u1_n101, u2_u3_u1_n102, u2_u3_u1_n103, u2_u3_u1_n104, u2_u3_u1_n105, u2_u3_u1_n106, u2_u3_u1_n107, u2_u3_u1_n108, u2_u3_u1_n109, 
       u2_u3_u1_n110, u2_u3_u1_n111, u2_u3_u1_n112, u2_u3_u1_n113, u2_u3_u1_n114, u2_u3_u1_n115, u2_u3_u1_n116, u2_u3_u1_n117, u2_u3_u1_n118, 
       u2_u3_u1_n119, u2_u3_u1_n120, u2_u3_u1_n121, u2_u3_u1_n122, u2_u3_u1_n123, u2_u3_u1_n124, u2_u3_u1_n125, u2_u3_u1_n126, u2_u3_u1_n127, 
       u2_u3_u1_n128, u2_u3_u1_n129, u2_u3_u1_n130, u2_u3_u1_n131, u2_u3_u1_n132, u2_u3_u1_n133, u2_u3_u1_n134, u2_u3_u1_n135, u2_u3_u1_n136, 
       u2_u3_u1_n137, u2_u3_u1_n138, u2_u3_u1_n139, u2_u3_u1_n140, u2_u3_u1_n141, u2_u3_u1_n142, u2_u3_u1_n143, u2_u3_u1_n144, u2_u3_u1_n145, 
       u2_u3_u1_n146, u2_u3_u1_n147, u2_u3_u1_n148, u2_u3_u1_n149, u2_u3_u1_n150, u2_u3_u1_n151, u2_u3_u1_n152, u2_u3_u1_n153, u2_u3_u1_n154, 
       u2_u3_u1_n155, u2_u3_u1_n156, u2_u3_u1_n157, u2_u3_u1_n158, u2_u3_u1_n159, u2_u3_u1_n160, u2_u3_u1_n161, u2_u3_u1_n162, u2_u3_u1_n163, 
       u2_u3_u1_n164, u2_u3_u1_n165, u2_u3_u1_n166, u2_u3_u1_n167, u2_u3_u1_n168, u2_u3_u1_n169, u2_u3_u1_n170, u2_u3_u1_n171, u2_u3_u1_n172, 
       u2_u3_u1_n173, u2_u3_u1_n174, u2_u3_u1_n175, u2_u3_u1_n176, u2_u3_u1_n177, u2_u3_u1_n178, u2_u3_u1_n179, u2_u3_u1_n180, u2_u3_u1_n181, 
       u2_u3_u1_n182, u2_u3_u1_n183, u2_u3_u1_n184, u2_u3_u1_n185, u2_u3_u1_n186, u2_u3_u1_n187, u2_u3_u1_n188, u2_u3_u1_n95, u2_u3_u1_n96, 
       u2_u3_u1_n97, u2_u3_u1_n98, u2_u3_u1_n99, u2_u3_u7_n100, u2_u3_u7_n101, u2_u3_u7_n102, u2_u3_u7_n103, u2_u3_u7_n104, u2_u3_u7_n105, 
       u2_u3_u7_n106, u2_u3_u7_n107, u2_u3_u7_n108, u2_u3_u7_n109, u2_u3_u7_n110, u2_u3_u7_n111, u2_u3_u7_n112, u2_u3_u7_n113, u2_u3_u7_n114, 
       u2_u3_u7_n115, u2_u3_u7_n116, u2_u3_u7_n117, u2_u3_u7_n118, u2_u3_u7_n119, u2_u3_u7_n120, u2_u3_u7_n121, u2_u3_u7_n122, u2_u3_u7_n123, 
       u2_u3_u7_n124, u2_u3_u7_n125, u2_u3_u7_n126, u2_u3_u7_n127, u2_u3_u7_n128, u2_u3_u7_n129, u2_u3_u7_n130, u2_u3_u7_n131, u2_u3_u7_n132, 
       u2_u3_u7_n133, u2_u3_u7_n134, u2_u3_u7_n135, u2_u3_u7_n136, u2_u3_u7_n137, u2_u3_u7_n138, u2_u3_u7_n139, u2_u3_u7_n140, u2_u3_u7_n141, 
       u2_u3_u7_n142, u2_u3_u7_n143, u2_u3_u7_n144, u2_u3_u7_n145, u2_u3_u7_n146, u2_u3_u7_n147, u2_u3_u7_n148, u2_u3_u7_n149, u2_u3_u7_n150, 
       u2_u3_u7_n151, u2_u3_u7_n152, u2_u3_u7_n153, u2_u3_u7_n154, u2_u3_u7_n155, u2_u3_u7_n156, u2_u3_u7_n157, u2_u3_u7_n158, u2_u3_u7_n159, 
       u2_u3_u7_n160, u2_u3_u7_n161, u2_u3_u7_n162, u2_u3_u7_n163, u2_u3_u7_n164, u2_u3_u7_n165, u2_u3_u7_n166, u2_u3_u7_n167, u2_u3_u7_n168, 
       u2_u3_u7_n169, u2_u3_u7_n170, u2_u3_u7_n171, u2_u3_u7_n172, u2_u3_u7_n173, u2_u3_u7_n174, u2_u3_u7_n175, u2_u3_u7_n176, u2_u3_u7_n177, 
       u2_u3_u7_n178, u2_u3_u7_n179, u2_u3_u7_n180, u2_u3_u7_n91, u2_u3_u7_n92, u2_u3_u7_n93, u2_u3_u7_n94, u2_u3_u7_n95, u2_u3_u7_n96, 
       u2_u3_u7_n97, u2_u3_u7_n98, u2_u3_u7_n99, u2_u5_X_25, u2_u5_X_26, u2_u5_X_27, u2_u5_X_28, u2_u5_X_29, u2_u5_X_30, 
       u2_u5_u4_n100, u2_u5_u4_n101, u2_u5_u4_n102, u2_u5_u4_n103, u2_u5_u4_n104, u2_u5_u4_n105, u2_u5_u4_n106, u2_u5_u4_n107, u2_u5_u4_n108, 
       u2_u5_u4_n109, u2_u5_u4_n110, u2_u5_u4_n111, u2_u5_u4_n112, u2_u5_u4_n113, u2_u5_u4_n114, u2_u5_u4_n115, u2_u5_u4_n116, u2_u5_u4_n117, 
       u2_u5_u4_n118, u2_u5_u4_n119, u2_u5_u4_n120, u2_u5_u4_n121, u2_u5_u4_n122, u2_u5_u4_n123, u2_u5_u4_n124, u2_u5_u4_n125, u2_u5_u4_n126, 
       u2_u5_u4_n127, u2_u5_u4_n128, u2_u5_u4_n129, u2_u5_u4_n130, u2_u5_u4_n131, u2_u5_u4_n132, u2_u5_u4_n133, u2_u5_u4_n134, u2_u5_u4_n135, 
       u2_u5_u4_n136, u2_u5_u4_n137, u2_u5_u4_n138, u2_u5_u4_n139, u2_u5_u4_n140, u2_u5_u4_n141, u2_u5_u4_n142, u2_u5_u4_n143, u2_u5_u4_n144, 
       u2_u5_u4_n145, u2_u5_u4_n146, u2_u5_u4_n147, u2_u5_u4_n148, u2_u5_u4_n149, u2_u5_u4_n150, u2_u5_u4_n151, u2_u5_u4_n152, u2_u5_u4_n153, 
       u2_u5_u4_n154, u2_u5_u4_n155, u2_u5_u4_n156, u2_u5_u4_n157, u2_u5_u4_n158, u2_u5_u4_n159, u2_u5_u4_n160, u2_u5_u4_n161, u2_u5_u4_n162, 
       u2_u5_u4_n163, u2_u5_u4_n164, u2_u5_u4_n165, u2_u5_u4_n166, u2_u5_u4_n167, u2_u5_u4_n168, u2_u5_u4_n169, u2_u5_u4_n170, u2_u5_u4_n171, 
       u2_u5_u4_n172, u2_u5_u4_n173, u2_u5_u4_n174, u2_u5_u4_n175, u2_u5_u4_n176, u2_u5_u4_n177, u2_u5_u4_n178, u2_u5_u4_n179, u2_u5_u4_n180, 
       u2_u5_u4_n181, u2_u5_u4_n182, u2_u5_u4_n183, u2_u5_u4_n184, u2_u5_u4_n185, u2_u5_u4_n186, u2_u5_u4_n94, u2_u5_u4_n95, u2_u5_u4_n96, 
       u2_u5_u4_n97, u2_u5_u4_n98, u2_u5_u4_n99, u2_u7_X_19, u2_u7_X_20, u2_u7_X_21, u2_u7_X_22, u2_u7_X_23, u2_u7_X_24, 
       u2_u7_X_25, u2_u7_X_26, u2_u7_X_27, u2_u7_X_28, u2_u7_X_29, u2_u7_X_30, u2_u7_X_31, u2_u7_X_32, u2_u7_X_33, 
       u2_u7_X_34, u2_u7_X_35, u2_u7_X_36, u2_u7_X_37, u2_u7_X_38, u2_u7_X_39, u2_u7_X_40, u2_u7_X_41, u2_u7_X_42, 
       u2_u7_u3_n100, u2_u7_u3_n101, u2_u7_u3_n102, u2_u7_u3_n103, u2_u7_u3_n104, u2_u7_u3_n105, u2_u7_u3_n106, u2_u7_u3_n107, u2_u7_u3_n108, 
       u2_u7_u3_n109, u2_u7_u3_n110, u2_u7_u3_n111, u2_u7_u3_n112, u2_u7_u3_n113, u2_u7_u3_n114, u2_u7_u3_n115, u2_u7_u3_n116, u2_u7_u3_n117, 
       u2_u7_u3_n118, u2_u7_u3_n119, u2_u7_u3_n120, u2_u7_u3_n121, u2_u7_u3_n122, u2_u7_u3_n123, u2_u7_u3_n124, u2_u7_u3_n125, u2_u7_u3_n126, 
       u2_u7_u3_n127, u2_u7_u3_n128, u2_u7_u3_n129, u2_u7_u3_n130, u2_u7_u3_n131, u2_u7_u3_n132, u2_u7_u3_n133, u2_u7_u3_n134, u2_u7_u3_n135, 
       u2_u7_u3_n136, u2_u7_u3_n137, u2_u7_u3_n138, u2_u7_u3_n139, u2_u7_u3_n140, u2_u7_u3_n141, u2_u7_u3_n142, u2_u7_u3_n143, u2_u7_u3_n144, 
       u2_u7_u3_n145, u2_u7_u3_n146, u2_u7_u3_n147, u2_u7_u3_n148, u2_u7_u3_n149, u2_u7_u3_n150, u2_u7_u3_n151, u2_u7_u3_n152, u2_u7_u3_n153, 
       u2_u7_u3_n154, u2_u7_u3_n155, u2_u7_u3_n156, u2_u7_u3_n157, u2_u7_u3_n158, u2_u7_u3_n159, u2_u7_u3_n160, u2_u7_u3_n161, u2_u7_u3_n162, 
       u2_u7_u3_n163, u2_u7_u3_n164, u2_u7_u3_n165, u2_u7_u3_n166, u2_u7_u3_n167, u2_u7_u3_n168, u2_u7_u3_n169, u2_u7_u3_n170, u2_u7_u3_n171, 
       u2_u7_u3_n172, u2_u7_u3_n173, u2_u7_u3_n174, u2_u7_u3_n175, u2_u7_u3_n176, u2_u7_u3_n177, u2_u7_u3_n178, u2_u7_u3_n179, u2_u7_u3_n180, 
       u2_u7_u3_n181, u2_u7_u3_n182, u2_u7_u3_n183, u2_u7_u3_n184, u2_u7_u3_n185, u2_u7_u3_n186, u2_u7_u3_n94, u2_u7_u3_n95, u2_u7_u3_n96, 
       u2_u7_u3_n97, u2_u7_u3_n98, u2_u7_u3_n99, u2_u7_u4_n100, u2_u7_u4_n101, u2_u7_u4_n102, u2_u7_u4_n103, u2_u7_u4_n104, u2_u7_u4_n105, 
       u2_u7_u4_n106, u2_u7_u4_n107, u2_u7_u4_n108, u2_u7_u4_n109, u2_u7_u4_n110, u2_u7_u4_n111, u2_u7_u4_n112, u2_u7_u4_n113, u2_u7_u4_n114, 
       u2_u7_u4_n115, u2_u7_u4_n116, u2_u7_u4_n117, u2_u7_u4_n118, u2_u7_u4_n119, u2_u7_u4_n120, u2_u7_u4_n121, u2_u7_u4_n122, u2_u7_u4_n123, 
       u2_u7_u4_n124, u2_u7_u4_n125, u2_u7_u4_n126, u2_u7_u4_n127, u2_u7_u4_n128, u2_u7_u4_n129, u2_u7_u4_n130, u2_u7_u4_n131, u2_u7_u4_n132, 
       u2_u7_u4_n133, u2_u7_u4_n134, u2_u7_u4_n135, u2_u7_u4_n136, u2_u7_u4_n137, u2_u7_u4_n138, u2_u7_u4_n139, u2_u7_u4_n140, u2_u7_u4_n141, 
       u2_u7_u4_n142, u2_u7_u4_n143, u2_u7_u4_n144, u2_u7_u4_n145, u2_u7_u4_n146, u2_u7_u4_n147, u2_u7_u4_n148, u2_u7_u4_n149, u2_u7_u4_n150, 
       u2_u7_u4_n151, u2_u7_u4_n152, u2_u7_u4_n153, u2_u7_u4_n154, u2_u7_u4_n155, u2_u7_u4_n156, u2_u7_u4_n157, u2_u7_u4_n158, u2_u7_u4_n159, 
       u2_u7_u4_n160, u2_u7_u4_n161, u2_u7_u4_n162, u2_u7_u4_n163, u2_u7_u4_n164, u2_u7_u4_n165, u2_u7_u4_n166, u2_u7_u4_n167, u2_u7_u4_n168, 
       u2_u7_u4_n169, u2_u7_u4_n170, u2_u7_u4_n171, u2_u7_u4_n172, u2_u7_u4_n173, u2_u7_u4_n174, u2_u7_u4_n175, u2_u7_u4_n176, u2_u7_u4_n177, 
       u2_u7_u4_n178, u2_u7_u4_n179, u2_u7_u4_n180, u2_u7_u4_n181, u2_u7_u4_n182, u2_u7_u4_n183, u2_u7_u4_n184, u2_u7_u4_n185, u2_u7_u4_n186, 
       u2_u7_u4_n94, u2_u7_u4_n95, u2_u7_u4_n96, u2_u7_u4_n97, u2_u7_u4_n98, u2_u7_u4_n99, u2_u7_u5_n100, u2_u7_u5_n101, u2_u7_u5_n102, 
       u2_u7_u5_n103, u2_u7_u5_n104, u2_u7_u5_n105, u2_u7_u5_n106, u2_u7_u5_n107, u2_u7_u5_n108, u2_u7_u5_n109, u2_u7_u5_n110, u2_u7_u5_n111, 
       u2_u7_u5_n112, u2_u7_u5_n113, u2_u7_u5_n114, u2_u7_u5_n115, u2_u7_u5_n116, u2_u7_u5_n117, u2_u7_u5_n118, u2_u7_u5_n119, u2_u7_u5_n120, 
       u2_u7_u5_n121, u2_u7_u5_n122, u2_u7_u5_n123, u2_u7_u5_n124, u2_u7_u5_n125, u2_u7_u5_n126, u2_u7_u5_n127, u2_u7_u5_n128, u2_u7_u5_n129, 
       u2_u7_u5_n130, u2_u7_u5_n131, u2_u7_u5_n132, u2_u7_u5_n133, u2_u7_u5_n134, u2_u7_u5_n135, u2_u7_u5_n136, u2_u7_u5_n137, u2_u7_u5_n138, 
       u2_u7_u5_n139, u2_u7_u5_n140, u2_u7_u5_n141, u2_u7_u5_n142, u2_u7_u5_n143, u2_u7_u5_n144, u2_u7_u5_n145, u2_u7_u5_n146, u2_u7_u5_n147, 
       u2_u7_u5_n148, u2_u7_u5_n149, u2_u7_u5_n150, u2_u7_u5_n151, u2_u7_u5_n152, u2_u7_u5_n153, u2_u7_u5_n154, u2_u7_u5_n155, u2_u7_u5_n156, 
       u2_u7_u5_n157, u2_u7_u5_n158, u2_u7_u5_n159, u2_u7_u5_n160, u2_u7_u5_n161, u2_u7_u5_n162, u2_u7_u5_n163, u2_u7_u5_n164, u2_u7_u5_n165, 
       u2_u7_u5_n166, u2_u7_u5_n167, u2_u7_u5_n168, u2_u7_u5_n169, u2_u7_u5_n170, u2_u7_u5_n171, u2_u7_u5_n172, u2_u7_u5_n173, u2_u7_u5_n174, 
       u2_u7_u5_n175, u2_u7_u5_n176, u2_u7_u5_n177, u2_u7_u5_n178, u2_u7_u5_n179, u2_u7_u5_n180, u2_u7_u5_n181, u2_u7_u5_n182, u2_u7_u5_n183, 
       u2_u7_u5_n184, u2_u7_u5_n185, u2_u7_u5_n186, u2_u7_u5_n187, u2_u7_u5_n188, u2_u7_u5_n189, u2_u7_u5_n190, u2_u7_u5_n191, u2_u7_u5_n192, 
       u2_u7_u5_n193, u2_u7_u5_n194, u2_u7_u5_n195, u2_u7_u5_n196, u2_u7_u5_n99, u2_u7_u6_n100, u2_u7_u6_n101, u2_u7_u6_n102, u2_u7_u6_n103, 
       u2_u7_u6_n104, u2_u7_u6_n105, u2_u7_u6_n106, u2_u7_u6_n107, u2_u7_u6_n108, u2_u7_u6_n109, u2_u7_u6_n110, u2_u7_u6_n111, u2_u7_u6_n112, 
       u2_u7_u6_n113, u2_u7_u6_n114, u2_u7_u6_n115, u2_u7_u6_n116, u2_u7_u6_n117, u2_u7_u6_n118, u2_u7_u6_n119, u2_u7_u6_n120, u2_u7_u6_n121, 
       u2_u7_u6_n122, u2_u7_u6_n123, u2_u7_u6_n124, u2_u7_u6_n125, u2_u7_u6_n126, u2_u7_u6_n127, u2_u7_u6_n128, u2_u7_u6_n129, u2_u7_u6_n130, 
       u2_u7_u6_n131, u2_u7_u6_n132, u2_u7_u6_n133, u2_u7_u6_n134, u2_u7_u6_n135, u2_u7_u6_n136, u2_u7_u6_n137, u2_u7_u6_n138, u2_u7_u6_n139, 
       u2_u7_u6_n140, u2_u7_u6_n141, u2_u7_u6_n142, u2_u7_u6_n143, u2_u7_u6_n144, u2_u7_u6_n145, u2_u7_u6_n146, u2_u7_u6_n147, u2_u7_u6_n148, 
       u2_u7_u6_n149, u2_u7_u6_n150, u2_u7_u6_n151, u2_u7_u6_n152, u2_u7_u6_n153, u2_u7_u6_n154, u2_u7_u6_n155, u2_u7_u6_n156, u2_u7_u6_n157, 
       u2_u7_u6_n158, u2_u7_u6_n159, u2_u7_u6_n160, u2_u7_u6_n161, u2_u7_u6_n162, u2_u7_u6_n163, u2_u7_u6_n164, u2_u7_u6_n165, u2_u7_u6_n166, 
       u2_u7_u6_n167, u2_u7_u6_n168, u2_u7_u6_n169, u2_u7_u6_n170, u2_u7_u6_n171, u2_u7_u6_n172, u2_u7_u6_n173, u2_u7_u6_n174, u2_u7_u6_n88, 
       u2_u7_u6_n89, u2_u7_u6_n90, u2_u7_u6_n91, u2_u7_u6_n92, u2_u7_u6_n93, u2_u7_u6_n94, u2_u7_u6_n95, u2_u7_u6_n96, u2_u7_u6_n97, 
       u2_u7_u6_n98, u2_u7_u6_n99, u2_uk_n1020, u2_uk_n1023, u2_uk_n1037, u2_uk_n1064, u2_uk_n1065, u2_uk_n1103, u2_uk_n1106, 
       u2_uk_n1108, u2_uk_n1109, u2_uk_n369, u2_uk_n524, u2_uk_n582, u2_uk_n587, u2_uk_n590, u2_uk_n603, u2_uk_n676, 
       u2_uk_n678,  u2_uk_n681;
  XOR2_X1 u0_U148 (.Z( u0_N4 ) , .B( u0_desIn_r_38 ) , .A( u0_out0_5 ) );
  XOR2_X1 u0_U167 (.B( u0_L10_31 ) , .Z( u0_N382 ) , .A( u0_out11_31 ) );
  XOR2_X1 u0_U168 (.B( u0_L10_30 ) , .Z( u0_N381 ) , .A( u0_out11_30 ) );
  XOR2_X1 u0_U171 (.B( u0_L10_28 ) , .Z( u0_N379 ) , .A( u0_out11_28 ) );
  XOR2_X1 u0_U173 (.B( u0_L10_26 ) , .Z( u0_N377 ) , .A( u0_out11_26 ) );
  XOR2_X1 u0_U175 (.B( u0_L10_24 ) , .Z( u0_N375 ) , .A( u0_out11_24 ) );
  XOR2_X1 u0_U176 (.B( u0_L10_23 ) , .Z( u0_N374 ) , .A( u0_out11_23 ) );
  XOR2_X1 u0_U179 (.B( u0_L10_20 ) , .Z( u0_N371 ) , .A( u0_out11_20 ) );
  XOR2_X1 u0_U182 (.B( u0_L10_18 ) , .Z( u0_N369 ) , .A( u0_out11_18 ) );
  XOR2_X1 u0_U183 (.B( u0_L10_17 ) , .Z( u0_N368 ) , .A( u0_out11_17 ) );
  XOR2_X1 u0_U184 (.B( u0_L10_16 ) , .Z( u0_N367 ) , .A( u0_out11_16 ) );
  XOR2_X1 u0_U187 (.B( u0_L10_13 ) , .Z( u0_N364 ) , .A( u0_out11_13 ) );
  XOR2_X1 u0_U190 (.B( u0_L10_10 ) , .Z( u0_N361 ) , .A( u0_out11_10 ) );
  XOR2_X1 u0_U191 (.B( u0_L10_9 ) , .Z( u0_N360 ) , .A( u0_out11_9 ) );
  XOR2_X1 u0_U195 (.B( u0_L10_6 ) , .Z( u0_N357 ) , .A( u0_out11_6 ) );
  XOR2_X1 u0_U199 (.B( u0_L10_2 ) , .Z( u0_N353 ) , .A( u0_out11_2 ) );
  XOR2_X1 u0_U200 (.B( u0_L10_1 ) , .Z( u0_N352 ) , .A( u0_out11_1 ) );
  XOR2_X1 u0_U247 (.Z( u0_N31 ) , .B( u0_desIn_r_56 ) , .A( u0_out0_32 ) );
  XOR2_X1 u0_U259 (.Z( u0_N3 ) , .B( u0_desIn_r_30 ) , .A( u0_out0_4 ) );
  XOR2_X1 u0_U281 (.Z( u0_N28 ) , .B( u0_desIn_r_32 ) , .A( u0_out0_29 ) );
  XOR2_X1 u0_U303 (.Z( u0_N26 ) , .B( u0_desIn_r_16 ) , .A( u0_out0_27 ) );
  XOR2_X1 u0_U325 (.Z( u0_N24 ) , .B( u0_desIn_r_0 ) , .A( u0_out0_25 ) );
  XOR2_X1 u0_U35 (.Z( u0_N7 ) , .B( u0_desIn_r_62 ) , .A( u0_out0_8 ) );
  XOR2_X1 u0_U358 (.Z( u0_N21 ) , .B( u0_desIn_r_42 ) , .A( u0_out0_22 ) );
  XOR2_X1 u0_U369 (.Z( u0_N20 ) , .B( u0_desIn_r_34 ) , .A( u0_out0_21 ) );
  XOR2_X1 u0_U370 (.Z( u0_N2 ) , .B( u0_desIn_r_22 ) , .A( u0_out0_3 ) );
  XOR2_X1 u0_U392 (.Z( u0_N18 ) , .B( u0_desIn_r_18 ) , .A( u0_out0_19 ) );
  XOR2_X1 u0_U415 (.B( u0_L3_32 ) , .Z( u0_N159 ) , .A( u0_out4_32 ) );
  XOR2_X1 u0_U418 (.B( u0_L3_29 ) , .Z( u0_N156 ) , .A( u0_out4_29 ) );
  XOR2_X1 u0_U422 (.B( u0_L3_25 ) , .Z( u0_N152 ) , .A( u0_out4_25 ) );
  XOR2_X1 u0_U426 (.B( u0_L3_22 ) , .Z( u0_N149 ) , .A( u0_out4_22 ) );
  XOR2_X1 u0_U429 (.B( u0_L3_19 ) , .Z( u0_N146 ) , .A( u0_out4_19 ) );
  XOR2_X1 u0_U434 (.B( u0_L3_14 ) , .Z( u0_N141 ) , .A( u0_out4_14 ) );
  XOR2_X1 u0_U436 (.Z( u0_N14 ) , .B( u0_desIn_r_52 ) , .A( u0_out0_15 ) );
  XOR2_X1 u0_U437 (.B( u0_L3_12 ) , .Z( u0_N139 ) , .A( u0_out4_12 ) );
  XOR2_X1 u0_U438 (.B( u0_L3_11 ) , .Z( u0_N138 ) , .A( u0_out4_11 ) );
  XOR2_X1 u0_U441 (.B( u0_L3_8 ) , .Z( u0_N135 ) , .A( u0_out4_8 ) );
  XOR2_X1 u0_U442 (.B( u0_L3_7 ) , .Z( u0_N134 ) , .A( u0_out4_7 ) );
  XOR2_X1 u0_U445 (.B( u0_L3_4 ) , .Z( u0_N131 ) , .A( u0_out4_4 ) );
  XOR2_X1 u0_U446 (.B( u0_L3_3 ) , .Z( u0_N130 ) , .A( u0_out4_3 ) );
  XOR2_X1 u0_U447 (.Z( u0_N13 ) , .B( u0_desIn_r_44 ) , .A( u0_out0_14 ) );
  XOR2_X1 u0_U46 (.Z( u0_N6 ) , .B( u0_desIn_r_54 ) , .A( u0_out0_7 ) );
  XOR2_X1 u0_U469 (.Z( u0_N11 ) , .B( u0_desIn_r_28 ) , .A( u0_out0_12 ) );
  XOR2_X1 u0_U480 (.Z( u0_N10 ) , .B( u0_desIn_r_20 ) , .A( u0_out0_11 ) );
  XOR2_X1 u0_U486 (.Z( u0_FP_6 ) , .B( u0_L14_6 ) , .A( u0_out15_6 ) );
  XOR2_X1 u0_U487 (.Z( u0_FP_5 ) , .B( u0_L14_5 ) , .A( u0_out15_5 ) );
  XOR2_X1 u0_U492 (.Z( u0_FP_30 ) , .B( u0_L14_30 ) , .A( u0_out15_30 ) );
  XOR2_X1 u0_U496 (.Z( u0_FP_27 ) , .B( u0_L14_27 ) , .A( u0_out15_27 ) );
  XOR2_X1 u0_U497 (.Z( u0_FP_26 ) , .B( u0_L14_26 ) , .A( u0_out15_26 ) );
  XOR2_X1 u0_U499 (.Z( u0_FP_24 ) , .B( u0_L14_24 ) , .A( u0_out15_24 ) );
  XOR2_X1 u0_U502 (.Z( u0_FP_21 ) , .B( u0_L14_21 ) , .A( u0_out15_21 ) );
  XOR2_X1 u0_U503 (.Z( u0_FP_20 ) , .B( u0_L14_20 ) , .A( u0_out15_20 ) );
  XOR2_X1 u0_U504 (.Z( u0_FP_1 ) , .B( u0_L14_1 ) , .A( u0_out15_1 ) );
  XOR2_X1 u0_U508 (.Z( u0_FP_16 ) , .B( u0_L14_16 ) , .A( u0_out15_16 ) );
  XOR2_X1 u0_U509 (.Z( u0_FP_15 ) , .B( u0_L14_15 ) , .A( u0_out15_15 ) );
  XOR2_X1 u0_U514 (.Z( u0_FP_10 ) , .B( u0_L14_10 ) , .A( u0_out15_10 ) );
  XOR2_X1 u0_u0_U10 (.B( u0_K1_45 ) , .A( u0_desIn_r_41 ) , .Z( u0_u0_X_45 ) );
  XOR2_X1 u0_u0_U11 (.B( u0_K1_44 ) , .A( u0_desIn_r_33 ) , .Z( u0_u0_X_44 ) );
  XOR2_X1 u0_u0_U12 (.B( u0_K1_43 ) , .A( u0_desIn_r_25 ) , .Z( u0_u0_X_43 ) );
  XOR2_X1 u0_u0_U13 (.B( u0_K1_42 ) , .A( u0_desIn_r_33 ) , .Z( u0_u0_X_42 ) );
  XOR2_X1 u0_u0_U14 (.B( u0_K1_41 ) , .A( u0_desIn_r_25 ) , .Z( u0_u0_X_41 ) );
  XOR2_X1 u0_u0_U15 (.B( u0_K1_40 ) , .A( u0_desIn_r_17 ) , .Z( u0_u0_X_40 ) );
  XOR2_X1 u0_u0_U17 (.B( u0_K1_39 ) , .A( u0_desIn_r_9 ) , .Z( u0_u0_X_39 ) );
  XOR2_X1 u0_u0_U18 (.B( u0_K1_38 ) , .A( u0_desIn_r_1 ) , .Z( u0_u0_X_38 ) );
  XOR2_X1 u0_u0_U19 (.B( u0_K1_37 ) , .A( u0_desIn_r_59 ) , .Z( u0_u0_X_37 ) );
  XOR2_X1 u0_u0_U20 (.B( u0_K1_36 ) , .A( u0_desIn_r_1 ) , .Z( u0_u0_X_36 ) );
  XOR2_X1 u0_u0_U21 (.B( u0_K1_35 ) , .A( u0_desIn_r_59 ) , .Z( u0_u0_X_35 ) );
  XOR2_X1 u0_u0_U22 (.B( u0_K1_34 ) , .A( u0_desIn_r_51 ) , .Z( u0_u0_X_34 ) );
  XOR2_X1 u0_u0_U23 (.B( u0_K1_33 ) , .A( u0_desIn_r_43 ) , .Z( u0_u0_X_33 ) );
  XOR2_X1 u0_u0_U24 (.B( u0_K1_32 ) , .A( u0_desIn_r_35 ) , .Z( u0_u0_X_32 ) );
  XOR2_X1 u0_u0_U25 (.B( u0_K1_31 ) , .A( u0_desIn_r_27 ) , .Z( u0_u0_X_31 ) );
  XOR2_X1 u0_u0_U26 (.B( u0_K1_30 ) , .A( u0_desIn_r_35 ) , .Z( u0_u0_X_30 ) );
  XOR2_X1 u0_u0_U28 (.B( u0_K1_29 ) , .A( u0_desIn_r_27 ) , .Z( u0_u0_X_29 ) );
  XOR2_X1 u0_u0_U29 (.B( u0_K1_28 ) , .A( u0_desIn_r_19 ) , .Z( u0_u0_X_28 ) );
  XOR2_X1 u0_u0_U30 (.B( u0_K1_27 ) , .A( u0_desIn_r_11 ) , .Z( u0_u0_X_27 ) );
  XOR2_X1 u0_u0_U31 (.B( u0_K1_26 ) , .A( u0_desIn_r_3 ) , .Z( u0_u0_X_26 ) );
  XOR2_X1 u0_u0_U32 (.B( u0_K1_25 ) , .A( u0_desIn_r_61 ) , .Z( u0_u0_X_25 ) );
  XOR2_X1 u0_u0_U7 (.B( u0_K1_48 ) , .A( u0_desIn_r_7 ) , .Z( u0_u0_X_48 ) );
  XOR2_X1 u0_u0_U8 (.B( u0_K1_47 ) , .A( u0_desIn_r_57 ) , .Z( u0_u0_X_47 ) );
  XOR2_X1 u0_u0_U9 (.B( u0_K1_46 ) , .A( u0_desIn_r_49 ) , .Z( u0_u0_X_46 ) );
  OAI22_X1 u0_u0_u4_U10 (.A2( u0_u0_u4_n16 ) , .A1( u0_u0_u4_n32 ) , .B1( u0_u0_u4_n34 ) , .ZN( u0_u0_u4_n50 ) , .B2( u0_u0_u4_n52 ) );
  AND3_X1 u0_u0_u4_U11 (.A1( u0_u0_u4_n30 ) , .A3( u0_u0_u4_n42 ) , .ZN( u0_u0_u4_n52 ) , .A2( u0_u0_u4_n53 ) );
  NAND2_X1 u0_u0_u4_U12 (.A1( u0_u0_u4_n14 ) , .A2( u0_u0_u4_n17 ) , .ZN( u0_u0_u4_n55 ) );
  AOI21_X1 u0_u0_u4_U13 (.A( u0_u0_u4_n17 ) , .ZN( u0_u0_u4_n25 ) , .B1( u0_u0_u4_n26 ) , .B2( u0_u0_u4_n27 ) );
  AOI21_X1 u0_u0_u4_U14 (.A( u0_u0_u4_n13 ) , .B1( u0_u0_u4_n3 ) , .B2( u0_u0_u4_n44 ) , .ZN( u0_u0_u4_n80 ) );
  AOI21_X1 u0_u0_u4_U15 (.A( u0_u0_u4_n13 ) , .ZN( u0_u0_u4_n24 ) , .B1( u0_u0_u4_n28 ) , .B2( u0_u0_u4_n29 ) );
  AOI21_X1 u0_u0_u4_U16 (.ZN( u0_u0_u4_n22 ) , .B1( u0_u0_u4_n32 ) , .B2( u0_u0_u4_n33 ) , .A( u0_u0_u4_n34 ) );
  AOI21_X1 u0_u0_u4_U17 (.ZN( u0_u0_u4_n23 ) , .B1( u0_u0_u4_n3 ) , .B2( u0_u0_u4_n30 ) , .A( u0_u0_u4_n31 ) );
  INV_X1 u0_u0_u4_U18 (.ZN( u0_u0_u4_n17 ) , .A( u0_u0_u4_n49 ) );
  AND2_X1 u0_u0_u4_U19 (.A1( u0_u0_u4_n27 ) , .ZN( u0_u0_u4_n32 ) , .A2( u0_u0_u4_n67 ) );
  INV_X1 u0_u0_u4_U20 (.ZN( u0_u0_u4_n12 ) , .A( u0_u0_u4_n31 ) );
  NAND2_X1 u0_u0_u4_U21 (.A1( u0_u0_u4_n40 ) , .ZN( u0_u0_u4_n56 ) , .A2( u0_u0_u4_n69 ) );
  NAND2_X1 u0_u0_u4_U22 (.ZN( u0_u0_u4_n57 ) , .A2( u0_u0_u4_n67 ) , .A1( u0_u0_u4_n68 ) );
  NAND2_X1 u0_u0_u4_U23 (.A1( u0_u0_u4_n39 ) , .A2( u0_u0_u4_n69 ) , .ZN( u0_u0_u4_n70 ) );
  NAND2_X1 u0_u0_u4_U24 (.A2( u0_u0_u4_n39 ) , .A1( u0_u0_u4_n53 ) , .ZN( u0_u0_u4_n58 ) );
  AND3_X1 u0_u0_u4_U25 (.ZN( u0_u0_u4_n26 ) , .A3( u0_u0_u4_n33 ) , .A2( u0_u0_u4_n44 ) , .A1( u0_u0_u4_n68 ) );
  AND2_X1 u0_u0_u4_U26 (.ZN( u0_u0_u4_n28 ) , .A2( u0_u0_u4_n40 ) , .A1( u0_u0_u4_n42 ) );
  OR3_X1 u0_u0_u4_U27 (.ZN( u0_u0_u4_n51 ) , .A1( u0_u0_u4_n71 ) , .A2( u0_u0_u4_n72 ) , .A3( u0_u0_u4_n73 ) );
  AOI21_X1 u0_u0_u4_U28 (.B1( u0_u0_u4_n13 ) , .B2( u0_u0_u4_n14 ) , .ZN( u0_u0_u4_n71 ) , .A( u0_u0_u4_n74 ) );
  AOI21_X1 u0_u0_u4_U29 (.A( u0_u0_u4_n31 ) , .B1( u0_u0_u4_n41 ) , .B2( u0_u0_u4_n42 ) , .ZN( u0_u0_u4_n72 ) );
  NOR2_X1 u0_u0_u4_U3 (.A2( u0_u0_u4_n5 ) , .A1( u0_u0_u4_n6 ) , .ZN( u0_u0_u4_n66 ) );
  OAI22_X1 u0_u0_u4_U30 (.A1( u0_u0_u4_n16 ) , .B2( u0_u0_u4_n17 ) , .B1( u0_u0_u4_n27 ) , .A2( u0_u0_u4_n66 ) , .ZN( u0_u0_u4_n73 ) );
  INV_X1 u0_u0_u4_U31 (.A( u0_u0_u4_n29 ) , .ZN( u0_u0_u4_n5 ) );
  INV_X1 u0_u0_u4_U32 (.ZN( u0_u0_u4_n6 ) , .A( u0_u0_u4_n91 ) );
  INV_X1 u0_u0_u4_U33 (.A( u0_u0_u4_n43 ) , .ZN( u0_u0_u4_n8 ) );
  INV_X1 u0_u0_u4_U34 (.A( u0_u0_u4_n30 ) , .ZN( u0_u0_u4_n9 ) );
  NAND2_X1 u0_u0_u4_U35 (.A2( u0_u0_u4_n33 ) , .ZN( u0_u0_u4_n90 ) , .A1( u0_u0_u4_n91 ) );
  INV_X1 u0_u0_u4_U36 (.ZN( u0_u0_u4_n1 ) , .A( u0_u0_u4_n92 ) );
  OAI221_X1 u0_u0_u4_U37 (.C2( u0_u0_u4_n14 ) , .B2( u0_u0_u4_n16 ) , .B1( u0_u0_u4_n29 ) , .C1( u0_u0_u4_n53 ) , .ZN( u0_u0_u4_n92 ) , .A( u0_u0_u4_n93 ) );
  AOI222_X1 u0_u0_u4_U38 (.C2( u0_u0_u4_n12 ) , .B1( u0_u0_u4_n2 ) , .A1( u0_u0_u4_n49 ) , .B2( u0_u0_u4_n55 ) , .C1( u0_u0_u4_n6 ) , .A2( u0_u0_u4_n8 ) , .ZN( u0_u0_u4_n93 ) );
  INV_X1 u0_u0_u4_U39 (.ZN( u0_u0_u4_n2 ) , .A( u0_u0_u4_n74 ) );
  INV_X1 u0_u0_u4_U4 (.ZN( u0_u0_u4_n3 ) , .A( u0_u0_u4_n70 ) );
  INV_X1 u0_u0_u4_U40 (.ZN( u0_u0_u4_n4 ) , .A( u0_u0_u4_n44 ) );
  NOR2_X1 u0_u0_u4_U41 (.A2( u0_u0_u4_n18 ) , .A1( u0_u0_u4_n19 ) , .ZN( u0_u0_u4_n49 ) );
  NOR2_X1 u0_u0_u4_U42 (.ZN( u0_u0_u4_n34 ) , .A2( u0_u0_u4_n35 ) , .A1( u0_u0_u4_n37 ) );
  NOR2_X1 u0_u0_u4_U43 (.ZN( u0_u0_u4_n31 ) , .A1( u0_u0_u4_n49 ) , .A2( u0_u0_u4_n59 ) );
  AOI22_X1 u0_u0_u4_U44 (.A2( u0_u0_u4_n15 ) , .B1( u0_u0_u4_n59 ) , .ZN( u0_u0_u4_n63 ) , .A1( u0_u0_u4_n64 ) , .B2( u0_u0_u4_n65 ) );
  INV_X1 u0_u0_u4_U45 (.ZN( u0_u0_u4_n15 ) , .A( u0_u0_u4_n34 ) );
  NAND2_X1 u0_u0_u4_U46 (.A1( u0_u0_u4_n26 ) , .ZN( u0_u0_u4_n64 ) , .A2( u0_u0_u4_n67 ) );
  AOI22_X1 u0_u0_u4_U47 (.A1( u0_u0_u4_n37 ) , .ZN( u0_u0_u4_n47 ) , .A2( u0_u0_u4_n54 ) , .B2( u0_u0_u4_n55 ) , .B1( u0_u0_u4_n8 ) );
  NAND2_X1 u0_u0_u4_U48 (.A1( u0_u0_u4_n33 ) , .A2( u0_u0_u4_n41 ) , .ZN( u0_u0_u4_n54 ) );
  NAND2_X1 u0_u0_u4_U49 (.ZN( u0_u0_u4_n33 ) , .A1( u0_u0_u4_n84 ) , .A2( u0_u0_u4_n89 ) );
  NOR4_X1 u0_u0_u4_U5 (.ZN( u0_u0_u4_n77 ) , .A1( u0_u0_u4_n78 ) , .A2( u0_u0_u4_n79 ) , .A3( u0_u0_u4_n80 ) , .A4( u0_u0_u4_n81 ) );
  NAND2_X1 u0_u0_u4_U50 (.ZN( u0_u0_u4_n29 ) , .A1( u0_u0_u4_n86 ) , .A2( u0_u0_u4_n88 ) );
  AOI21_X1 u0_u0_u4_U51 (.B2( u0_u0_u4_n37 ) , .A( u0_u0_u4_n51 ) , .ZN( u0_u0_u4_n60 ) , .B1( u0_u0_u4_n7 ) );
  INV_X1 u0_u0_u4_U52 (.A( u0_u0_u4_n27 ) , .ZN( u0_u0_u4_n7 ) );
  NAND2_X1 u0_u0_u4_U53 (.ZN( u0_u0_u4_n41 ) , .A1( u0_u0_u4_n82 ) , .A2( u0_u0_u4_n83 ) );
  NAND2_X1 u0_u0_u4_U54 (.ZN( u0_u0_u4_n27 ) , .A1( u0_u0_u4_n85 ) , .A2( u0_u0_u4_n86 ) );
  NAND2_X1 u0_u0_u4_U55 (.ZN( u0_u0_u4_n53 ) , .A2( u0_u0_u4_n88 ) , .A1( u0_u0_u4_n89 ) );
  NAND2_X1 u0_u0_u4_U56 (.ZN( u0_u0_u4_n44 ) , .A2( u0_u0_u4_n83 ) , .A1( u0_u0_u4_n84 ) );
  NAND2_X1 u0_u0_u4_U57 (.ZN( u0_u0_u4_n42 ) , .A2( u0_u0_u4_n82 ) , .A1( u0_u0_u4_n89 ) );
  NAND2_X1 u0_u0_u4_U58 (.ZN( u0_u0_u4_n67 ) , .A2( u0_u0_u4_n82 ) , .A1( u0_u0_u4_n87 ) );
  NAND2_X1 u0_u0_u4_U59 (.ZN( u0_u0_u4_n39 ) , .A2( u0_u0_u4_n83 ) , .A1( u0_u0_u4_n85 ) );
  AOI21_X1 u0_u0_u4_U6 (.A( u0_u0_u4_n17 ) , .B1( u0_u0_u4_n29 ) , .B2( u0_u0_u4_n41 ) , .ZN( u0_u0_u4_n81 ) );
  NAND2_X1 u0_u0_u4_U60 (.ZN( u0_u0_u4_n30 ) , .A1( u0_u0_u4_n84 ) , .A2( u0_u0_u4_n87 ) );
  INV_X1 u0_u0_u4_U61 (.ZN( u0_u0_u4_n14 ) , .A( u0_u0_u4_n37 ) );
  INV_X1 u0_u0_u4_U62 (.ZN( u0_u0_u4_n16 ) , .A( u0_u0_u4_n35 ) );
  NAND2_X1 u0_u0_u4_U63 (.ZN( u0_u0_u4_n69 ) , .A1( u0_u0_u4_n87 ) , .A2( u0_u0_u4_n88 ) );
  NAND2_X1 u0_u0_u4_U64 (.ZN( u0_u0_u4_n43 ) , .A1( u0_u0_u4_n85 ) , .A2( u0_u0_u4_n87 ) );
  NAND2_X1 u0_u0_u4_U65 (.A1( u0_u0_u4_n82 ) , .A2( u0_u0_u4_n86 ) , .ZN( u0_u0_u4_n91 ) );
  INV_X1 u0_u0_u4_U66 (.ZN( u0_u0_u4_n13 ) , .A( u0_u0_u4_n59 ) );
  NAND2_X1 u0_u0_u4_U67 (.ZN( u0_u0_u4_n68 ) , .A2( u0_u0_u4_n85 ) , .A1( u0_u0_u4_n89 ) );
  NAND2_X1 u0_u0_u4_U68 (.ZN( u0_u0_u4_n40 ) , .A1( u0_u0_u4_n84 ) , .A2( u0_u0_u4_n86 ) );
  NAND2_X1 u0_u0_u4_U69 (.ZN( u0_u0_u4_n74 ) , .A2( u0_u0_u4_n83 ) , .A1( u0_u0_u4_n88 ) );
  AOI21_X1 u0_u0_u4_U7 (.A( u0_u0_u4_n31 ) , .B1( u0_u0_u4_n32 ) , .B2( u0_u0_u4_n53 ) , .ZN( u0_u0_u4_n79 ) );
  NOR2_X1 u0_u0_u4_U70 (.A2( u0_u0_X_28 ) , .A1( u0_u0_u4_n19 ) , .ZN( u0_u0_u4_n37 ) );
  NOR2_X1 u0_u0_u4_U71 (.A2( u0_u0_X_29 ) , .A1( u0_u0_u4_n18 ) , .ZN( u0_u0_u4_n35 ) );
  NOR2_X1 u0_u0_u4_U72 (.A2( u0_u0_X_30 ) , .A1( u0_u0_u4_n11 ) , .ZN( u0_u0_u4_n82 ) );
  NOR2_X1 u0_u0_u4_U73 (.A2( u0_u0_X_26 ) , .A1( u0_u0_u4_n10 ) , .ZN( u0_u0_u4_n87 ) );
  NOR2_X1 u0_u0_u4_U74 (.A2( u0_u0_X_28 ) , .A1( u0_u0_X_29 ) , .ZN( u0_u0_u4_n59 ) );
  NOR2_X1 u0_u0_u4_U75 (.A2( u0_u0_X_27 ) , .A1( u0_u0_X_30 ) , .ZN( u0_u0_u4_n85 ) );
  NOR2_X1 u0_u0_u4_U76 (.A2( u0_u0_X_25 ) , .A1( u0_u0_X_26 ) , .ZN( u0_u0_u4_n89 ) );
  AND2_X1 u0_u0_u4_U77 (.A2( u0_u0_X_25 ) , .A1( u0_u0_X_26 ) , .ZN( u0_u0_u4_n83 ) );
  AND2_X1 u0_u0_u4_U78 (.A1( u0_u0_X_30 ) , .A2( u0_u0_u4_n11 ) , .ZN( u0_u0_u4_n88 ) );
  AND2_X1 u0_u0_u4_U79 (.A1( u0_u0_X_26 ) , .A2( u0_u0_u4_n10 ) , .ZN( u0_u0_u4_n86 ) );
  AOI21_X1 u0_u0_u4_U8 (.B1( u0_u0_u4_n28 ) , .B2( u0_u0_u4_n3 ) , .A( u0_u0_u4_n34 ) , .ZN( u0_u0_u4_n78 ) );
  AND2_X1 u0_u0_u4_U80 (.A1( u0_u0_X_27 ) , .A2( u0_u0_X_30 ) , .ZN( u0_u0_u4_n84 ) );
  INV_X1 u0_u0_u4_U81 (.A( u0_u0_X_28 ) , .ZN( u0_u0_u4_n18 ) );
  INV_X1 u0_u0_u4_U82 (.A( u0_u0_X_29 ) , .ZN( u0_u0_u4_n19 ) );
  INV_X1 u0_u0_u4_U83 (.A( u0_u0_X_25 ) , .ZN( u0_u0_u4_n10 ) );
  INV_X1 u0_u0_u4_U84 (.A( u0_u0_X_27 ) , .ZN( u0_u0_u4_n11 ) );
  NAND4_X1 u0_u0_u4_U85 (.ZN( u0_out0_25 ) , .A1( u0_u0_u4_n45 ) , .A2( u0_u0_u4_n46 ) , .A3( u0_u0_u4_n47 ) , .A4( u0_u0_u4_n48 ) );
  OAI21_X1 u0_u0_u4_U86 (.ZN( u0_u0_u4_n45 ) , .B1( u0_u0_u4_n57 ) , .B2( u0_u0_u4_n58 ) , .A( u0_u0_u4_n59 ) );
  OAI21_X1 u0_u0_u4_U87 (.A( u0_u0_u4_n12 ) , .B1( u0_u0_u4_n4 ) , .ZN( u0_u0_u4_n46 ) , .B2( u0_u0_u4_n56 ) );
  NAND4_X1 u0_u0_u4_U88 (.ZN( u0_out0_14 ) , .A1( u0_u0_u4_n60 ) , .A2( u0_u0_u4_n61 ) , .A3( u0_u0_u4_n62 ) , .A4( u0_u0_u4_n63 ) );
  AOI22_X1 u0_u0_u4_U89 (.A2( u0_u0_u4_n12 ) , .B1( u0_u0_u4_n35 ) , .A1( u0_u0_u4_n58 ) , .ZN( u0_u0_u4_n61 ) , .B2( u0_u0_u4_n70 ) );
  AOI211_X1 u0_u0_u4_U9 (.ZN( u0_u0_u4_n48 ) , .C2( u0_u0_u4_n49 ) , .C1( u0_u0_u4_n5 ) , .A( u0_u0_u4_n50 ) , .B( u0_u0_u4_n51 ) );
  AOI22_X1 u0_u0_u4_U90 (.B1( u0_u0_u4_n49 ) , .A2( u0_u0_u4_n55 ) , .B2( u0_u0_u4_n56 ) , .ZN( u0_u0_u4_n62 ) , .A1( u0_u0_u4_n9 ) );
  NAND4_X1 u0_u0_u4_U91 (.ZN( u0_out0_8 ) , .A1( u0_u0_u4_n1 ) , .A2( u0_u0_u4_n75 ) , .A3( u0_u0_u4_n76 ) , .A4( u0_u0_u4_n77 ) );
  NAND2_X1 u0_u0_u4_U92 (.A1( u0_u0_u4_n37 ) , .A2( u0_u0_u4_n57 ) , .ZN( u0_u0_u4_n75 ) );
  AOI22_X1 u0_u0_u4_U93 (.A1( u0_u0_u4_n35 ) , .B2( u0_u0_u4_n55 ) , .ZN( u0_u0_u4_n76 ) , .B1( u0_u0_u4_n9 ) , .A2( u0_u0_u4_n90 ) );
  AOI22_X1 u0_u0_u4_U94 (.ZN( u0_u0_u4_n20 ) , .A1( u0_u0_u4_n35 ) , .A2( u0_u0_u4_n36 ) , .B1( u0_u0_u4_n37 ) , .B2( u0_u0_u4_n38 ) );
  NOR4_X1 u0_u0_u4_U95 (.ZN( u0_u0_u4_n21 ) , .A1( u0_u0_u4_n22 ) , .A2( u0_u0_u4_n23 ) , .A3( u0_u0_u4_n24 ) , .A4( u0_u0_u4_n25 ) );
  NAND3_X1 u0_u0_u4_U96 (.ZN( u0_out0_3 ) , .A2( u0_u0_u4_n1 ) , .A1( u0_u0_u4_n20 ) , .A3( u0_u0_u4_n21 ) );
  NAND3_X1 u0_u0_u4_U97 (.ZN( u0_u0_u4_n38 ) , .A1( u0_u0_u4_n39 ) , .A2( u0_u0_u4_n40 ) , .A3( u0_u0_u4_n41 ) );
  NAND3_X1 u0_u0_u4_U98 (.ZN( u0_u0_u4_n36 ) , .A1( u0_u0_u4_n42 ) , .A2( u0_u0_u4_n43 ) , .A3( u0_u0_u4_n44 ) );
  NAND3_X1 u0_u0_u4_U99 (.A1( u0_u0_u4_n33 ) , .A2( u0_u0_u4_n43 ) , .ZN( u0_u0_u4_n65 ) , .A3( u0_u0_u4_n66 ) );
  INV_X1 u0_u0_u5_U10 (.ZN( u0_u0_u5_n20 ) , .A( u0_u0_u5_n76 ) );
  AOI222_X1 u0_u0_u5_U100 (.A2( u0_u0_u5_n18 ) , .C2( u0_u0_u5_n19 ) , .B2( u0_u0_u5_n23 ) , .C1( u0_u0_u5_n49 ) , .A1( u0_u0_u5_n66 ) , .ZN( u0_u0_u5_n84 ) , .B1( u0_u0_u5_n98 ) );
  NAND4_X1 u0_u0_u5_U101 (.ZN( u0_out0_29 ) , .A1( u0_u0_u5_n1 ) , .A2( u0_u0_u5_n29 ) , .A3( u0_u0_u5_n67 ) , .A4( u0_u0_u5_n68 ) );
  AOI221_X1 u0_u0_u5_U102 (.C1( u0_u0_u5_n13 ) , .B1( u0_u0_u5_n21 ) , .B2( u0_u0_u5_n38 ) , .C2( u0_u0_u5_n65 ) , .ZN( u0_u0_u5_n68 ) , .A( u0_u0_u5_n69 ) );
  AOI222_X1 u0_u0_u5_U103 (.B2( u0_u0_u5_n18 ) , .C2( u0_u0_u5_n22 ) , .C1( u0_u0_u5_n3 ) , .B1( u0_u0_u5_n50 ) , .A2( u0_u0_u5_n51 ) , .ZN( u0_u0_u5_n67 ) , .A1( u0_u0_u5_n9 ) );
  NAND3_X1 u0_u0_u5_U104 (.A1( u0_u0_u5_n36 ) , .A3( u0_u0_u5_n39 ) , .A2( u0_u0_u5_n43 ) , .ZN( u0_u0_u5_n98 ) );
  NOR2_X1 u0_u0_u5_U11 (.A1( u0_u0_u5_n20 ) , .A2( u0_u0_u5_n24 ) , .ZN( u0_u0_u5_n37 ) );
  INV_X1 u0_u0_u5_U12 (.ZN( u0_u0_u5_n23 ) , .A( u0_u0_u5_n47 ) );
  AOI21_X1 u0_u0_u5_U13 (.ZN( u0_u0_u5_n35 ) , .B2( u0_u0_u5_n36 ) , .A( u0_u0_u5_n37 ) , .B1( u0_u0_u5_n5 ) );
  INV_X1 u0_u0_u5_U14 (.A( u0_u0_u5_n38 ) , .ZN( u0_u0_u5_n5 ) );
  AOI21_X1 u0_u0_u5_U15 (.ZN( u0_u0_u5_n34 ) , .B1( u0_u0_u5_n39 ) , .B2( u0_u0_u5_n40 ) , .A( u0_u0_u5_n41 ) );
  AOI21_X1 u0_u0_u5_U16 (.A( u0_u0_u5_n47 ) , .ZN( u0_u0_u5_n56 ) , .B1( u0_u0_u5_n57 ) , .B2( u0_u0_u5_n58 ) );
  OAI21_X1 u0_u0_u5_U17 (.ZN( u0_u0_u5_n55 ) , .B1( u0_u0_u5_n62 ) , .B2( u0_u0_u5_n63 ) , .A( u0_u0_u5_n64 ) );
  OAI21_X1 u0_u0_u5_U18 (.A( u0_u0_u5_n24 ) , .B2( u0_u0_u5_n50 ) , .ZN( u0_u0_u5_n64 ) , .B1( u0_u0_u5_n9 ) );
  NAND2_X1 u0_u0_u5_U19 (.ZN( u0_u0_u5_n60 ) , .A1( u0_u0_u5_n74 ) , .A2( u0_u0_u5_n78 ) );
  INV_X1 u0_u0_u5_U20 (.ZN( u0_u0_u5_n3 ) , .A( u0_u0_u5_n42 ) );
  NAND2_X1 u0_u0_u5_U21 (.A2( u0_u0_u5_n25 ) , .ZN( u0_u0_u5_n65 ) , .A1( u0_u0_u5_n76 ) );
  NAND2_X1 u0_u0_u5_U22 (.A1( u0_u0_u5_n43 ) , .ZN( u0_u0_u5_n61 ) , .A2( u0_u0_u5_n75 ) );
  NAND2_X1 u0_u0_u5_U23 (.ZN( u0_u0_u5_n38 ) , .A1( u0_u0_u5_n77 ) , .A2( u0_u0_u5_n78 ) );
  INV_X1 u0_u0_u5_U24 (.ZN( u0_u0_u5_n22 ) , .A( u0_u0_u5_n41 ) );
  INV_X1 u0_u0_u5_U25 (.A( u0_u0_u5_n39 ) , .ZN( u0_u0_u5_n9 ) );
  INV_X1 u0_u0_u5_U26 (.ZN( u0_u0_u5_n18 ) , .A( u0_u0_u5_n45 ) );
  INV_X1 u0_u0_u5_U27 (.ZN( u0_u0_u5_n15 ) , .A( u0_u0_u5_n57 ) );
  INV_X1 u0_u0_u5_U28 (.ZN( u0_u0_u5_n14 ) , .A( u0_u0_u5_n46 ) );
  INV_X1 u0_u0_u5_U29 (.ZN( u0_u0_u5_n12 ) , .A( u0_u0_u5_n74 ) );
  NOR2_X1 u0_u0_u5_U3 (.A1( u0_u0_u5_n14 ) , .ZN( u0_u0_u5_n63 ) , .A2( u0_u0_u5_n7 ) );
  INV_X1 u0_u0_u5_U30 (.ZN( u0_u0_u5_n13 ) , .A( u0_u0_u5_n36 ) );
  INV_X1 u0_u0_u5_U31 (.A( u0_u0_u5_n58 ) , .ZN( u0_u0_u5_n8 ) );
  INV_X1 u0_u0_u5_U32 (.A( u0_u0_u5_n40 ) , .ZN( u0_u0_u5_n7 ) );
  INV_X1 u0_u0_u5_U33 (.ZN( u0_u0_u5_n4 ) , .A( u0_u0_u5_n77 ) );
  NAND2_X1 u0_u0_u5_U34 (.A2( u0_u0_u5_n42 ) , .A1( u0_u0_u5_n57 ) , .ZN( u0_u0_u5_n86 ) );
  NOR2_X1 u0_u0_u5_U35 (.A2( u0_u0_u5_n17 ) , .A1( u0_u0_u5_n27 ) , .ZN( u0_u0_u5_n97 ) );
  INV_X1 u0_u0_u5_U36 (.ZN( u0_u0_u5_n1 ) , .A( u0_u0_u5_n80 ) );
  OAI221_X1 u0_u0_u5_U37 (.B1( u0_u0_u5_n25 ) , .C2( u0_u0_u5_n39 ) , .C1( u0_u0_u5_n44 ) , .B2( u0_u0_u5_n78 ) , .ZN( u0_u0_u5_n80 ) , .A( u0_u0_u5_n81 ) );
  AOI222_X1 u0_u0_u5_U38 (.B1( u0_u0_u5_n10 ) , .C2( u0_u0_u5_n20 ) , .A2( u0_u0_u5_n23 ) , .A1( u0_u0_u5_n4 ) , .C1( u0_u0_u5_n49 ) , .B2( u0_u0_u5_n52 ) , .ZN( u0_u0_u5_n81 ) );
  INV_X1 u0_u0_u5_U39 (.ZN( u0_u0_u5_n10 ) , .A( u0_u0_u5_n82 ) );
  INV_X1 u0_u0_u5_U4 (.A( u0_u0_u5_n59 ) , .ZN( u0_u0_u5_n6 ) );
  AOI22_X1 u0_u0_u5_U40 (.A1( u0_u0_u5_n12 ) , .B1( u0_u0_u5_n23 ) , .ZN( u0_u0_u5_n28 ) , .A2( u0_u0_u5_n51 ) , .B2( u0_u0_u5_n66 ) );
  NOR2_X1 u0_u0_u5_U41 (.A2( u0_u0_u5_n24 ) , .ZN( u0_u0_u5_n47 ) , .A1( u0_u0_u5_n51 ) );
  AOI21_X1 u0_u0_u5_U42 (.B1( u0_u0_u5_n11 ) , .ZN( u0_u0_u5_n29 ) , .B2( u0_u0_u5_n52 ) , .A( u0_u0_u5_n79 ) );
  INV_X1 u0_u0_u5_U43 (.ZN( u0_u0_u5_n11 ) , .A( u0_u0_u5_n75 ) );
  NOR2_X1 u0_u0_u5_U44 (.A2( u0_u0_u5_n21 ) , .ZN( u0_u0_u5_n45 ) , .A1( u0_u0_u5_n51 ) );
  NOR2_X1 u0_u0_u5_U45 (.A2( u0_u0_u5_n44 ) , .ZN( u0_u0_u5_n79 ) , .A1( u0_u0_u5_n82 ) );
  NOR2_X1 u0_u0_u5_U46 (.A1( u0_u0_u5_n23 ) , .ZN( u0_u0_u5_n41 ) , .A2( u0_u0_u5_n52 ) );
  NOR2_X1 u0_u0_u5_U47 (.A1( u0_u0_u5_n21 ) , .A2( u0_u0_u5_n52 ) , .ZN( u0_u0_u5_n76 ) );
  AOI22_X1 u0_u0_u5_U48 (.B2( u0_u0_u5_n22 ) , .B1( u0_u0_u5_n4 ) , .A1( u0_u0_u5_n52 ) , .A2( u0_u0_u5_n60 ) , .ZN( u0_u0_u5_n83 ) );
  OAI211_X1 u0_u0_u5_U49 (.ZN( u0_u0_u5_n69 ) , .C1( u0_u0_u5_n70 ) , .C2( u0_u0_u5_n71 ) , .A( u0_u0_u5_n72 ) , .B( u0_u0_u5_n73 ) );
  OAI21_X1 u0_u0_u5_U5 (.A( u0_u0_u5_n20 ) , .ZN( u0_u0_u5_n59 ) , .B1( u0_u0_u5_n60 ) , .B2( u0_u0_u5_n61 ) );
  NOR3_X1 u0_u0_u5_U50 (.A2( u0_u0_u5_n15 ) , .A3( u0_u0_u5_n49 ) , .A1( u0_u0_u5_n61 ) , .ZN( u0_u0_u5_n70 ) );
  OAI21_X1 u0_u0_u5_U51 (.B2( u0_u0_u5_n14 ) , .A( u0_u0_u5_n20 ) , .ZN( u0_u0_u5_n73 ) , .B1( u0_u0_u5_n8 ) );
  OAI21_X1 u0_u0_u5_U52 (.B2( u0_u0_u5_n12 ) , .A( u0_u0_u5_n23 ) , .B1( u0_u0_u5_n7 ) , .ZN( u0_u0_u5_n72 ) );
  AOI21_X1 u0_u0_u5_U53 (.ZN( u0_u0_u5_n33 ) , .B1( u0_u0_u5_n42 ) , .B2( u0_u0_u5_n43 ) , .A( u0_u0_u5_n44 ) );
  AOI21_X1 u0_u0_u5_U54 (.A( u0_u0_u5_n44 ) , .B2( u0_u0_u5_n58 ) , .B1( u0_u0_u5_n75 ) , .ZN( u0_u0_u5_n87 ) );
  INV_X1 u0_u0_u5_U55 (.ZN( u0_u0_u5_n21 ) , .A( u0_u0_u5_n44 ) );
  INV_X1 u0_u0_u5_U56 (.ZN( u0_u0_u5_n24 ) , .A( u0_u0_u5_n71 ) );
  AND2_X1 u0_u0_u5_U57 (.ZN( u0_u0_u5_n50 ) , .A1( u0_u0_u5_n90 ) , .A2( u0_u0_u5_n93 ) );
  AND2_X1 u0_u0_u5_U58 (.ZN( u0_u0_u5_n49 ) , .A1( u0_u0_u5_n89 ) , .A2( u0_u0_u5_n93 ) );
  NAND2_X1 u0_u0_u5_U59 (.ZN( u0_u0_u5_n39 ) , .A2( u0_u0_u5_n91 ) , .A1( u0_u0_u5_n92 ) );
  INV_X1 u0_u0_u5_U6 (.ZN( u0_u0_u5_n19 ) , .A( u0_u0_u5_n62 ) );
  NAND2_X1 u0_u0_u5_U60 (.ZN( u0_u0_u5_n58 ) , .A1( u0_u0_u5_n88 ) , .A2( u0_u0_u5_n89 ) );
  NAND2_X1 u0_u0_u5_U61 (.ZN( u0_u0_u5_n78 ) , .A2( u0_u0_u5_n89 ) , .A1( u0_u0_u5_n91 ) );
  NAND2_X1 u0_u0_u5_U62 (.ZN( u0_u0_u5_n57 ) , .A1( u0_u0_u5_n92 ) , .A2( u0_u0_u5_n94 ) );
  NAND2_X1 u0_u0_u5_U63 (.ZN( u0_u0_u5_n42 ) , .A1( u0_u0_u5_n92 ) , .A2( u0_u0_u5_n93 ) );
  NAND2_X1 u0_u0_u5_U64 (.ZN( u0_u0_u5_n75 ) , .A1( u0_u0_u5_n90 ) , .A2( u0_u0_u5_n91 ) );
  NAND2_X1 u0_u0_u5_U65 (.ZN( u0_u0_u5_n82 ) , .A1( u0_u0_u5_n91 ) , .A2( u0_u0_u5_n97 ) );
  NAND2_X1 u0_u0_u5_U66 (.ZN( u0_u0_u5_n36 ) , .A1( u0_u0_u5_n94 ) , .A2( u0_u0_u5_n97 ) );
  NAND2_X1 u0_u0_u5_U67 (.ZN( u0_u0_u5_n43 ) , .A2( u0_u0_u5_n88 ) , .A1( u0_u0_u5_n92 ) );
  INV_X1 u0_u0_u5_U68 (.ZN( u0_u0_u5_n25 ) , .A( u0_u0_u5_n51 ) );
  NAND2_X1 u0_u0_u5_U69 (.ZN( u0_u0_u5_n74 ) , .A2( u0_u0_u5_n89 ) , .A1( u0_u0_u5_n94 ) );
  OAI22_X1 u0_u0_u5_U7 (.ZN( u0_u0_u5_n32 ) , .A1( u0_u0_u5_n45 ) , .A2( u0_u0_u5_n46 ) , .B1( u0_u0_u5_n47 ) , .B2( u0_u0_u5_n48 ) );
  NAND2_X1 u0_u0_u5_U70 (.ZN( u0_u0_u5_n46 ) , .A1( u0_u0_u5_n90 ) , .A2( u0_u0_u5_n94 ) );
  NAND2_X1 u0_u0_u5_U71 (.ZN( u0_u0_u5_n77 ) , .A1( u0_u0_u5_n88 ) , .A2( u0_u0_u5_n90 ) );
  NAND2_X1 u0_u0_u5_U72 (.ZN( u0_u0_u5_n40 ) , .A1( u0_u0_u5_n88 ) , .A2( u0_u0_u5_n97 ) );
  AND2_X1 u0_u0_u5_U73 (.ZN( u0_u0_u5_n66 ) , .A1( u0_u0_u5_n93 ) , .A2( u0_u0_u5_n97 ) );
  INV_X1 u0_u0_u5_U74 (.ZN( u0_u0_u5_n2 ) , .A( u0_u0_u5_n95 ) );
  OAI221_X1 u0_u0_u5_U75 (.B2( u0_u0_u5_n37 ) , .B1( u0_u0_u5_n63 ) , .C1( u0_u0_u5_n71 ) , .C2( u0_u0_u5_n82 ) , .ZN( u0_u0_u5_n95 ) , .A( u0_u0_u5_n96 ) );
  OAI21_X1 u0_u0_u5_U76 (.B2( u0_u0_u5_n50 ) , .A( u0_u0_u5_n51 ) , .B1( u0_u0_u5_n60 ) , .ZN( u0_u0_u5_n96 ) );
  NOR2_X1 u0_u0_u5_U77 (.A2( u0_u0_X_34 ) , .A1( u0_u0_X_35 ) , .ZN( u0_u0_u5_n52 ) );
  NOR2_X1 u0_u0_u5_U78 (.A2( u0_u0_X_34 ) , .A1( u0_u0_u5_n26 ) , .ZN( u0_u0_u5_n51 ) );
  NOR2_X1 u0_u0_u5_U79 (.A2( u0_u0_X_31 ) , .A1( u0_u0_X_32 ) , .ZN( u0_u0_u5_n94 ) );
  NOR3_X1 u0_u0_u5_U8 (.A3( u0_u0_u5_n3 ) , .ZN( u0_u0_u5_n48 ) , .A1( u0_u0_u5_n49 ) , .A2( u0_u0_u5_n50 ) );
  NOR2_X1 u0_u0_u5_U80 (.A2( u0_u0_X_36 ) , .A1( u0_u0_u5_n17 ) , .ZN( u0_u0_u5_n92 ) );
  NOR2_X1 u0_u0_u5_U81 (.A2( u0_u0_X_33 ) , .A1( u0_u0_u5_n27 ) , .ZN( u0_u0_u5_n89 ) );
  NOR2_X1 u0_u0_u5_U82 (.A2( u0_u0_X_33 ) , .A1( u0_u0_X_36 ) , .ZN( u0_u0_u5_n90 ) );
  NOR2_X1 u0_u0_u5_U83 (.A2( u0_u0_X_31 ) , .A1( u0_u0_u5_n16 ) , .ZN( u0_u0_u5_n93 ) );
  NAND2_X1 u0_u0_u5_U84 (.A2( u0_u0_X_34 ) , .A1( u0_u0_X_35 ) , .ZN( u0_u0_u5_n44 ) );
  NAND2_X1 u0_u0_u5_U85 (.A1( u0_u0_X_34 ) , .A2( u0_u0_u5_n26 ) , .ZN( u0_u0_u5_n71 ) );
  AND2_X1 u0_u0_u5_U86 (.A1( u0_u0_X_31 ) , .A2( u0_u0_X_32 ) , .ZN( u0_u0_u5_n91 ) );
  AND2_X1 u0_u0_u5_U87 (.A1( u0_u0_X_31 ) , .A2( u0_u0_u5_n16 ) , .ZN( u0_u0_u5_n88 ) );
  INV_X1 u0_u0_u5_U88 (.A( u0_u0_X_33 ) , .ZN( u0_u0_u5_n17 ) );
  INV_X1 u0_u0_u5_U89 (.A( u0_u0_X_35 ) , .ZN( u0_u0_u5_n26 ) );
  NOR2_X1 u0_u0_u5_U9 (.A2( u0_u0_u5_n21 ) , .A1( u0_u0_u5_n24 ) , .ZN( u0_u0_u5_n62 ) );
  INV_X1 u0_u0_u5_U90 (.A( u0_u0_X_36 ) , .ZN( u0_u0_u5_n27 ) );
  INV_X1 u0_u0_u5_U91 (.A( u0_u0_X_32 ) , .ZN( u0_u0_u5_n16 ) );
  NAND4_X1 u0_u0_u5_U92 (.ZN( u0_out0_19 ) , .A1( u0_u0_u5_n28 ) , .A2( u0_u0_u5_n29 ) , .A3( u0_u0_u5_n30 ) , .A4( u0_u0_u5_n31 ) );
  AOI22_X1 u0_u0_u5_U93 (.B1( u0_u0_u5_n15 ) , .ZN( u0_u0_u5_n30 ) , .A2( u0_u0_u5_n51 ) , .B2( u0_u0_u5_n52 ) , .A1( u0_u0_u5_n8 ) );
  NOR4_X1 u0_u0_u5_U94 (.ZN( u0_u0_u5_n31 ) , .A1( u0_u0_u5_n32 ) , .A2( u0_u0_u5_n33 ) , .A3( u0_u0_u5_n34 ) , .A4( u0_u0_u5_n35 ) );
  NAND4_X1 u0_u0_u5_U95 (.ZN( u0_out0_11 ) , .A1( u0_u0_u5_n1 ) , .A2( u0_u0_u5_n28 ) , .A3( u0_u0_u5_n53 ) , .A4( u0_u0_u5_n54 ) );
  AOI22_X1 u0_u0_u5_U96 (.B1( u0_u0_u5_n13 ) , .A1( u0_u0_u5_n3 ) , .B2( u0_u0_u5_n52 ) , .ZN( u0_u0_u5_n53 ) , .A2( u0_u0_u5_n65 ) );
  NOR3_X1 u0_u0_u5_U97 (.ZN( u0_u0_u5_n54 ) , .A1( u0_u0_u5_n55 ) , .A3( u0_u0_u5_n56 ) , .A2( u0_u0_u5_n6 ) );
  NAND4_X1 u0_u0_u5_U98 (.ZN( u0_out0_4 ) , .A3( u0_u0_u5_n2 ) , .A1( u0_u0_u5_n83 ) , .A2( u0_u0_u5_n84 ) , .A4( u0_u0_u5_n85 ) );
  AOI211_X1 u0_u0_u5_U99 (.C2( u0_u0_u5_n20 ) , .B( u0_u0_u5_n79 ) , .ZN( u0_u0_u5_n85 ) , .C1( u0_u0_u5_n86 ) , .A( u0_u0_u5_n87 ) );
  AOI22_X1 u0_u0_u6_U10 (.B2( u0_u0_u6_n14 ) , .A2( u0_u0_u6_n24 ) , .B1( u0_u0_u6_n5 ) , .A1( u0_u0_u6_n8 ) , .ZN( u0_u0_u6_n86 ) );
  AOI21_X1 u0_u0_u6_U11 (.A( u0_u0_u6_n17 ) , .B2( u0_u0_u6_n43 ) , .B1( u0_u0_u6_n68 ) , .ZN( u0_u0_u6_n87 ) );
  AOI21_X1 u0_u0_u6_U12 (.A( u0_u0_u6_n17 ) , .ZN( u0_u0_u6_n26 ) , .B1( u0_u0_u6_n27 ) , .B2( u0_u0_u6_n28 ) );
  AOI21_X1 u0_u0_u6_U13 (.B1( u0_u0_u6_n11 ) , .B2( u0_u0_u6_n16 ) , .A( u0_u0_u6_n33 ) , .ZN( u0_u0_u6_n69 ) );
  INV_X1 u0_u0_u6_U14 (.ZN( u0_u0_u6_n14 ) , .A( u0_u0_u6_n20 ) );
  INV_X1 u0_u0_u6_U15 (.ZN( u0_u0_u6_n11 ) , .A( u0_u0_u6_n47 ) );
  NAND2_X1 u0_u0_u6_U16 (.A2( u0_u0_u6_n46 ) , .A1( u0_u0_u6_n53 ) , .ZN( u0_u0_u6_n65 ) );
  NAND2_X1 u0_u0_u6_U17 (.A1( u0_u0_u6_n27 ) , .A2( u0_u0_u6_n29 ) , .ZN( u0_u0_u6_n51 ) );
  INV_X1 u0_u0_u6_U18 (.ZN( u0_u0_u6_n4 ) , .A( u0_u0_u6_n43 ) );
  AND2_X1 u0_u0_u6_U19 (.A2( u0_u0_u6_n28 ) , .ZN( u0_u0_u6_n45 ) , .A1( u0_u0_u6_n75 ) );
  INV_X1 u0_u0_u6_U20 (.ZN( u0_u0_u6_n2 ) , .A( u0_u0_u6_n48 ) );
  INV_X1 u0_u0_u6_U21 (.A( u0_u0_u6_n54 ) , .ZN( u0_u0_u6_n8 ) );
  INV_X1 u0_u0_u6_U22 (.ZN( u0_u0_u6_n6 ) , .A( u0_u0_u6_n75 ) );
  INV_X1 u0_u0_u6_U23 (.ZN( u0_u0_u6_n5 ) , .A( u0_u0_u6_n52 ) );
  INV_X1 u0_u0_u6_U24 (.A( u0_u0_u6_n62 ) , .ZN( u0_u0_u6_n7 ) );
  AND2_X1 u0_u0_u6_U25 (.ZN( u0_u0_u6_n42 ) , .A2( u0_u0_u6_n56 ) , .A1( u0_u0_u6_n68 ) );
  AND2_X1 u0_u0_u6_U26 (.ZN( u0_u0_u6_n44 ) , .A1( u0_u0_u6_n53 ) , .A2( u0_u0_u6_n54 ) );
  AND3_X1 u0_u0_u6_U27 (.A3( u0_u0_u6_n30 ) , .A1( u0_u0_u6_n43 ) , .A2( u0_u0_u6_n48 ) , .ZN( u0_u0_u6_n55 ) );
  INV_X1 u0_u0_u6_U28 (.ZN( u0_u0_u6_n12 ) , .A( u0_u0_u6_n29 ) );
  AOI222_X1 u0_u0_u6_U29 (.C2( u0_u0_u6_n16 ) , .B2( u0_u0_u6_n24 ) , .A2( u0_u0_u6_n49 ) , .A1( u0_u0_u6_n57 ) , .B1( u0_u0_u6_n6 ) , .ZN( u0_u0_u6_n61 ) , .C1( u0_u0_u6_n7 ) );
  INV_X1 u0_u0_u6_U3 (.A( u0_u0_u6_n65 ) , .ZN( u0_u0_u6_n9 ) );
  NOR2_X1 u0_u0_u6_U30 (.A2( u0_u0_u6_n10 ) , .A1( u0_u0_u6_n13 ) , .ZN( u0_u0_u6_n77 ) );
  AOI211_X1 u0_u0_u6_U31 (.C2( u0_u0_u6_n24 ) , .ZN( u0_u0_u6_n38 ) , .C1( u0_u0_u6_n39 ) , .A( u0_u0_u6_n40 ) , .B( u0_u0_u6_n41 ) );
  AOI21_X1 u0_u0_u6_U32 (.A( u0_u0_u6_n17 ) , .ZN( u0_u0_u6_n41 ) , .B1( u0_u0_u6_n42 ) , .B2( u0_u0_u6_n43 ) );
  NAND4_X1 u0_u0_u6_U33 (.ZN( u0_u0_u6_n39 ) , .A1( u0_u0_u6_n45 ) , .A2( u0_u0_u6_n46 ) , .A3( u0_u0_u6_n47 ) , .A4( u0_u0_u6_n48 ) );
  AOI21_X1 u0_u0_u6_U34 (.B2( u0_u0_u6_n29 ) , .A( u0_u0_u6_n31 ) , .ZN( u0_u0_u6_n40 ) , .B1( u0_u0_u6_n44 ) );
  NAND2_X1 u0_u0_u6_U35 (.A2( u0_u0_u6_n17 ) , .ZN( u0_u0_u6_n24 ) , .A1( u0_u0_u6_n31 ) );
  NAND2_X1 u0_u0_u6_U36 (.ZN( u0_u0_u6_n43 ) , .A2( u0_u0_u6_n78 ) , .A1( u0_u0_u6_n84 ) );
  AOI22_X1 u0_u0_u6_U37 (.A2( u0_u0_u6_n14 ) , .ZN( u0_u0_u6_n60 ) , .A1( u0_u0_u6_n63 ) , .B1( u0_u0_u6_n64 ) , .B2( u0_u0_u6_n65 ) );
  NAND4_X1 u0_u0_u6_U38 (.A2( u0_u0_u6_n28 ) , .A4( u0_u0_u6_n43 ) , .ZN( u0_u0_u6_n63 ) , .A3( u0_u0_u6_n66 ) , .A1( u0_u0_u6_n9 ) );
  NOR2_X1 u0_u0_u6_U39 (.A2( u0_u0_u6_n2 ) , .A1( u0_u0_u6_n5 ) , .ZN( u0_u0_u6_n66 ) );
  INV_X1 u0_u0_u6_U4 (.ZN( u0_u0_u6_n1 ) , .A( u0_u0_u6_n33 ) );
  NOR2_X1 u0_u0_u6_U40 (.A1( u0_u0_u6_n15 ) , .ZN( u0_u0_u6_n20 ) , .A2( u0_u0_u6_n49 ) );
  NAND2_X1 u0_u0_u6_U41 (.ZN( u0_u0_u6_n29 ) , .A1( u0_u0_u6_n76 ) , .A2( u0_u0_u6_n81 ) );
  AOI21_X1 u0_u0_u6_U42 (.ZN( u0_u0_u6_n25 ) , .B1( u0_u0_u6_n29 ) , .B2( u0_u0_u6_n30 ) , .A( u0_u0_u6_n31 ) );
  INV_X1 u0_u0_u6_U43 (.ZN( u0_u0_u6_n17 ) , .A( u0_u0_u6_n64 ) );
  NAND2_X1 u0_u0_u6_U44 (.ZN( u0_u0_u6_n48 ) , .A2( u0_u0_u6_n83 ) , .A1( u0_u0_u6_n84 ) );
  NAND2_X1 u0_u0_u6_U45 (.ZN( u0_u0_u6_n46 ) , .A1( u0_u0_u6_n79 ) , .A2( u0_u0_u6_n80 ) );
  INV_X1 u0_u0_u6_U46 (.ZN( u0_u0_u6_n16 ) , .A( u0_u0_u6_n31 ) );
  NAND2_X1 u0_u0_u6_U47 (.ZN( u0_u0_u6_n30 ) , .A1( u0_u0_u6_n77 ) , .A2( u0_u0_u6_n78 ) );
  NAND2_X1 u0_u0_u6_U48 (.ZN( u0_u0_u6_n27 ) , .A1( u0_u0_u6_n81 ) , .A2( u0_u0_u6_n83 ) );
  NAND2_X1 u0_u0_u6_U49 (.A1( u0_u0_u6_n31 ) , .A2( u0_u0_u6_n36 ) , .ZN( u0_u0_u6_n67 ) );
  NAND2_X1 u0_u0_u6_U5 (.ZN( u0_u0_u6_n23 ) , .A2( u0_u0_u6_n32 ) , .A1( u0_u0_u6_n9 ) );
  NAND2_X1 u0_u0_u6_U50 (.ZN( u0_u0_u6_n54 ) , .A1( u0_u0_u6_n78 ) , .A2( u0_u0_u6_n80 ) );
  NAND2_X1 u0_u0_u6_U51 (.ZN( u0_u0_u6_n68 ) , .A1( u0_u0_u6_n80 ) , .A2( u0_u0_u6_n83 ) );
  AND2_X1 u0_u0_u6_U52 (.ZN( u0_u0_u6_n57 ) , .A1( u0_u0_u6_n76 ) , .A2( u0_u0_u6_n84 ) );
  NAND2_X1 u0_u0_u6_U53 (.ZN( u0_u0_u6_n28 ) , .A1( u0_u0_u6_n76 ) , .A2( u0_u0_u6_n77 ) );
  NAND2_X1 u0_u0_u6_U54 (.ZN( u0_u0_u6_n47 ) , .A2( u0_u0_u6_n79 ) , .A1( u0_u0_u6_n81 ) );
  NAND2_X1 u0_u0_u6_U55 (.ZN( u0_u0_u6_n56 ) , .A1( u0_u0_u6_n76 ) , .A2( u0_u0_u6_n80 ) );
  NAND2_X1 u0_u0_u6_U56 (.ZN( u0_u0_u6_n52 ) , .A1( u0_u0_u6_n79 ) , .A2( u0_u0_u6_n84 ) );
  NAND2_X1 u0_u0_u6_U57 (.ZN( u0_u0_u6_n75 ) , .A1( u0_u0_u6_n77 ) , .A2( u0_u0_u6_n83 ) );
  NAND2_X1 u0_u0_u6_U58 (.ZN( u0_u0_u6_n53 ) , .A2( u0_u0_u6_n78 ) , .A1( u0_u0_u6_n81 ) );
  INV_X1 u0_u0_u6_U59 (.ZN( u0_u0_u6_n15 ) , .A( u0_u0_u6_n36 ) );
  AOI22_X1 u0_u0_u6_U6 (.A2( u0_u0_u6_n14 ) , .B1( u0_u0_u6_n15 ) , .ZN( u0_u0_u6_n72 ) , .A1( u0_u0_u6_n73 ) , .B2( u0_u0_u6_n74 ) );
  NAND2_X1 u0_u0_u6_U60 (.ZN( u0_u0_u6_n62 ) , .A2( u0_u0_u6_n77 ) , .A1( u0_u0_u6_n79 ) );
  NOR2_X1 u0_u0_u6_U61 (.A2( u0_u0_X_40 ) , .A1( u0_u0_X_41 ) , .ZN( u0_u0_u6_n49 ) );
  NOR2_X1 u0_u0_u6_U62 (.A2( u0_u0_X_39 ) , .A1( u0_u0_X_42 ) , .ZN( u0_u0_u6_n83 ) );
  NOR2_X1 u0_u0_u6_U63 (.A2( u0_u0_X_39 ) , .A1( u0_u0_u6_n19 ) , .ZN( u0_u0_u6_n78 ) );
  NOR2_X1 u0_u0_u6_U64 (.A2( u0_u0_X_38 ) , .A1( u0_u0_u6_n10 ) , .ZN( u0_u0_u6_n80 ) );
  NOR2_X1 u0_u0_u6_U65 (.A2( u0_u0_X_41 ) , .A1( u0_u0_u6_n18 ) , .ZN( u0_u0_u6_n64 ) );
  NOR2_X1 u0_u0_u6_U66 (.A2( u0_u0_X_37 ) , .A1( u0_u0_u6_n13 ) , .ZN( u0_u0_u6_n81 ) );
  NOR2_X1 u0_u0_u6_U67 (.A2( u0_u0_X_37 ) , .A1( u0_u0_X_38 ) , .ZN( u0_u0_u6_n84 ) );
  NAND2_X1 u0_u0_u6_U68 (.A1( u0_u0_X_41 ) , .A2( u0_u0_u6_n18 ) , .ZN( u0_u0_u6_n31 ) );
  NAND2_X1 u0_u0_u6_U69 (.A2( u0_u0_X_40 ) , .A1( u0_u0_X_41 ) , .ZN( u0_u0_u6_n36 ) );
  NOR2_X1 u0_u0_u6_U7 (.ZN( u0_u0_u6_n32 ) , .A1( u0_u0_u6_n57 ) , .A2( u0_u0_u6_n7 ) );
  AND2_X1 u0_u0_u6_U70 (.A1( u0_u0_X_39 ) , .A2( u0_u0_u6_n19 ) , .ZN( u0_u0_u6_n79 ) );
  AND2_X1 u0_u0_u6_U71 (.A1( u0_u0_X_39 ) , .A2( u0_u0_X_42 ) , .ZN( u0_u0_u6_n76 ) );
  INV_X1 u0_u0_u6_U72 (.A( u0_u0_X_40 ) , .ZN( u0_u0_u6_n18 ) );
  INV_X1 u0_u0_u6_U73 (.A( u0_u0_X_37 ) , .ZN( u0_u0_u6_n10 ) );
  INV_X1 u0_u0_u6_U74 (.A( u0_u0_X_38 ) , .ZN( u0_u0_u6_n13 ) );
  INV_X1 u0_u0_u6_U75 (.A( u0_u0_X_42 ) , .ZN( u0_u0_u6_n19 ) );
  NAND4_X1 u0_u0_u6_U76 (.ZN( u0_out0_12 ) , .A1( u0_u0_u6_n58 ) , .A2( u0_u0_u6_n59 ) , .A3( u0_u0_u6_n60 ) , .A4( u0_u0_u6_n61 ) );
  OAI22_X1 u0_u0_u6_U77 (.A2( u0_u0_u6_n11 ) , .B1( u0_u0_u6_n49 ) , .ZN( u0_u0_u6_n59 ) , .B2( u0_u0_u6_n64 ) , .A1( u0_u0_u6_n8 ) );
  OAI21_X1 u0_u0_u6_U78 (.B1( u0_u0_u6_n12 ) , .B2( u0_u0_u6_n34 ) , .ZN( u0_u0_u6_n58 ) , .A( u0_u0_u6_n67 ) );
  NAND4_X1 u0_u0_u6_U79 (.ZN( u0_out0_32 ) , .A1( u0_u0_u6_n69 ) , .A2( u0_u0_u6_n70 ) , .A3( u0_u0_u6_n71 ) , .A4( u0_u0_u6_n72 ) );
  OAI21_X1 u0_u0_u6_U8 (.A( u0_u0_u6_n16 ) , .B2( u0_u0_u6_n2 ) , .B1( u0_u0_u6_n6 ) , .ZN( u0_u0_u6_n85 ) );
  AOI22_X1 u0_u0_u6_U80 (.B1( u0_u0_u6_n4 ) , .B2( u0_u0_u6_n49 ) , .A1( u0_u0_u6_n57 ) , .A2( u0_u0_u6_n67 ) , .ZN( u0_u0_u6_n70 ) );
  AOI22_X1 u0_u0_u6_U81 (.B2( u0_u0_u6_n24 ) , .B1( u0_u0_u6_n51 ) , .A1( u0_u0_u6_n64 ) , .ZN( u0_u0_u6_n71 ) , .A2( u0_u0_u6_n82 ) );
  OAI211_X1 u0_u0_u6_U82 (.ZN( u0_out0_7 ) , .A( u0_u0_u6_n1 ) , .C1( u0_u0_u6_n20 ) , .C2( u0_u0_u6_n21 ) , .B( u0_u0_u6_n22 ) );
  NOR3_X1 u0_u0_u6_U83 (.A3( u0_u0_u6_n11 ) , .ZN( u0_u0_u6_n21 ) , .A1( u0_u0_u6_n34 ) , .A2( u0_u0_u6_n4 ) );
  AOI211_X1 u0_u0_u6_U84 (.ZN( u0_u0_u6_n22 ) , .C1( u0_u0_u6_n23 ) , .C2( u0_u0_u6_n24 ) , .A( u0_u0_u6_n25 ) , .B( u0_u0_u6_n26 ) );
  OAI211_X1 u0_u0_u6_U85 (.ZN( u0_out0_22 ) , .C1( u0_u0_u6_n35 ) , .C2( u0_u0_u6_n36 ) , .A( u0_u0_u6_n37 ) , .B( u0_u0_u6_n38 ) );
  AOI22_X1 u0_u0_u6_U86 (.B2( u0_u0_u6_n14 ) , .ZN( u0_u0_u6_n37 ) , .A1( u0_u0_u6_n49 ) , .A2( u0_u0_u6_n50 ) , .B1( u0_u0_u6_n51 ) );
  AND4_X1 u0_u0_u6_U87 (.A2( u0_u0_u6_n32 ) , .ZN( u0_u0_u6_n35 ) , .A4( u0_u0_u6_n46 ) , .A1( u0_u0_u6_n55 ) , .A3( u0_u0_u6_n56 ) );
  NAND3_X1 u0_u0_u6_U88 (.A3( u0_u0_u6_n44 ) , .A1( u0_u0_u6_n45 ) , .ZN( u0_u0_u6_n50 ) , .A2( u0_u0_u6_n52 ) );
  NAND3_X1 u0_u0_u6_U89 (.A2( u0_u0_u6_n27 ) , .A1( u0_u0_u6_n30 ) , .ZN( u0_u0_u6_n34 ) , .A3( u0_u0_u6_n42 ) );
  INV_X1 u0_u0_u6_U9 (.ZN( u0_u0_u6_n3 ) , .A( u0_u0_u6_n87 ) );
  NAND3_X1 u0_u0_u6_U90 (.A1( u0_u0_u6_n48 ) , .A2( u0_u0_u6_n54 ) , .A3( u0_u0_u6_n68 ) , .ZN( u0_u0_u6_n74 ) );
  NAND3_X1 u0_u0_u6_U91 (.A2( u0_u0_u6_n30 ) , .A3( u0_u0_u6_n45 ) , .ZN( u0_u0_u6_n73 ) , .A1( u0_u0_u6_n9 ) );
  NAND3_X1 u0_u0_u6_U92 (.A2( u0_u0_u6_n52 ) , .A1( u0_u0_u6_n56 ) , .A3( u0_u0_u6_n62 ) , .ZN( u0_u0_u6_n82 ) );
  NAND3_X1 u0_u0_u6_U93 (.A2( u0_u0_u6_n3 ) , .ZN( u0_u0_u6_n33 ) , .A1( u0_u0_u6_n85 ) , .A3( u0_u0_u6_n86 ) );
  OAI21_X1 u0_u0_u7_U10 (.B1( u0_u0_u7_n13 ) , .A( u0_u0_u7_n20 ) , .B2( u0_u0_u7_n8 ) , .ZN( u0_u0_u7_n90 ) );
  AOI211_X1 u0_u0_u7_U11 (.B( u0_u0_u7_n1 ) , .C1( u0_u0_u7_n4 ) , .C2( u0_u0_u7_n55 ) , .ZN( u0_u0_u7_n63 ) , .A( u0_u0_u7_n64 ) );
  OAI22_X1 u0_u0_u7_U12 (.B2( u0_u0_u7_n19 ) , .A1( u0_u0_u7_n44 ) , .A2( u0_u0_u7_n48 ) , .ZN( u0_u0_u7_n64 ) , .B1( u0_u0_u7_n66 ) );
  INV_X1 u0_u0_u7_U13 (.ZN( u0_u0_u7_n1 ) , .A( u0_u0_u7_n65 ) );
  NOR3_X1 u0_u0_u7_U14 (.A1( u0_u0_u7_n12 ) , .A2( u0_u0_u7_n13 ) , .A3( u0_u0_u7_n36 ) , .ZN( u0_u0_u7_n66 ) );
  INV_X1 u0_u0_u7_U15 (.A( u0_u0_u7_n48 ) , .ZN( u0_u0_u7_n5 ) );
  NOR3_X1 u0_u0_u7_U16 (.A3( u0_u0_u7_n10 ) , .ZN( u0_u0_u7_n45 ) , .A1( u0_u0_u7_n46 ) , .A2( u0_u0_u7_n47 ) );
  NOR2_X1 u0_u0_u7_U17 (.ZN( u0_u0_u7_n28 ) , .A2( u0_u0_u7_n47 ) , .A1( u0_u0_u7_n51 ) );
  AOI21_X1 u0_u0_u7_U18 (.A( u0_u0_u7_n17 ) , .B1( u0_u0_u7_n54 ) , .B2( u0_u0_u7_n69 ) , .ZN( u0_u0_u7_n77 ) );
  AOI21_X1 u0_u0_u7_U19 (.A( u0_u0_u7_n19 ) , .B2( u0_u0_u7_n35 ) , .B1( u0_u0_u7_n48 ) , .ZN( u0_u0_u7_n75 ) );
  AOI21_X1 u0_u0_u7_U20 (.B2( u0_u0_u7_n53 ) , .B1( u0_u0_u7_n6 ) , .ZN( u0_u0_u7_n74 ) , .A( u0_u0_u7_n80 ) );
  INV_X1 u0_u0_u7_U21 (.ZN( u0_u0_u7_n16 ) , .A( u0_u0_u7_n80 ) );
  NOR2_X1 u0_u0_u7_U22 (.A1( u0_u0_u7_n12 ) , .A2( u0_u0_u7_n47 ) , .ZN( u0_u0_u7_n70 ) );
  INV_X1 u0_u0_u7_U23 (.ZN( u0_u0_u7_n10 ) , .A( u0_u0_u7_n43 ) );
  INV_X1 u0_u0_u7_U24 (.ZN( u0_u0_u7_n4 ) , .A( u0_u0_u7_n50 ) );
  INV_X1 u0_u0_u7_U25 (.ZN( u0_u0_u7_n7 ) , .A( u0_u0_u7_n71 ) );
  NAND2_X1 u0_u0_u7_U26 (.ZN( u0_u0_u7_n32 ) , .A2( u0_u0_u7_n49 ) , .A1( u0_u0_u7_n52 ) );
  NAND2_X1 u0_u0_u7_U27 (.ZN( u0_u0_u7_n51 ) , .A2( u0_u0_u7_n57 ) , .A1( u0_u0_u7_n68 ) );
  INV_X1 u0_u0_u7_U28 (.A( u0_u0_u7_n69 ) , .ZN( u0_u0_u7_n8 ) );
  INV_X1 u0_u0_u7_U29 (.ZN( u0_u0_u7_n13 ) , .A( u0_u0_u7_n53 ) );
  OAI21_X1 u0_u0_u7_U3 (.B2( u0_u0_u7_n10 ) , .A( u0_u0_u7_n16 ) , .ZN( u0_u0_u7_n22 ) , .B1( u0_u0_u7_n7 ) );
  INV_X1 u0_u0_u7_U30 (.ZN( u0_u0_u7_n12 ) , .A( u0_u0_u7_n33 ) );
  INV_X1 u0_u0_u7_U31 (.ZN( u0_u0_u7_n2 ) , .A( u0_u0_u7_n54 ) );
  INV_X1 u0_u0_u7_U32 (.A( u0_u0_u7_n28 ) , .ZN( u0_u0_u7_n9 ) );
  NOR2_X1 u0_u0_u7_U33 (.A1( u0_u0_u7_n25 ) , .A2( u0_u0_u7_n31 ) , .ZN( u0_u0_u7_n80 ) );
  AOI211_X1 u0_u0_u7_U34 (.C1( u0_u0_u7_n25 ) , .ZN( u0_u0_u7_n39 ) , .C2( u0_u0_u7_n40 ) , .A( u0_u0_u7_n41 ) , .B( u0_u0_u7_n42 ) );
  NAND4_X1 u0_u0_u7_U35 (.A4( u0_u0_u7_n34 ) , .ZN( u0_u0_u7_n40 ) , .A1( u0_u0_u7_n52 ) , .A2( u0_u0_u7_n53 ) , .A3( u0_u0_u7_n54 ) );
  AOI21_X1 u0_u0_u7_U36 (.B2( u0_u0_u7_n35 ) , .ZN( u0_u0_u7_n42 ) , .B1( u0_u0_u7_n43 ) , .A( u0_u0_u7_n44 ) );
  OAI22_X1 u0_u0_u7_U37 (.A2( u0_u0_u7_n17 ) , .B2( u0_u0_u7_n19 ) , .A1( u0_u0_u7_n28 ) , .ZN( u0_u0_u7_n41 ) , .B1( u0_u0_u7_n45 ) );
  INV_X1 u0_u0_u7_U38 (.ZN( u0_u0_u7_n20 ) , .A( u0_u0_u7_n56 ) );
  AOI21_X1 u0_u0_u7_U39 (.B1( u0_u0_u7_n16 ) , .B2( u0_u0_u7_n4 ) , .ZN( u0_u0_u7_n58 ) , .A( u0_u0_u7_n84 ) );
  INV_X1 u0_u0_u7_U4 (.A( u0_u0_u7_n32 ) , .ZN( u0_u0_u7_n6 ) );
  AOI21_X1 u0_u0_u7_U40 (.A( u0_u0_u7_n56 ) , .B1( u0_u0_u7_n57 ) , .B2( u0_u0_u7_n68 ) , .ZN( u0_u0_u7_n84 ) );
  INV_X1 u0_u0_u7_U41 (.ZN( u0_u0_u7_n19 ) , .A( u0_u0_u7_n29 ) );
  AOI22_X1 u0_u0_u7_U42 (.B2( u0_u0_u7_n16 ) , .A1( u0_u0_u7_n25 ) , .B1( u0_u0_u7_n51 ) , .ZN( u0_u0_u7_n62 ) , .A2( u0_u0_u7_n67 ) );
  NAND2_X1 u0_u0_u7_U43 (.A1( u0_u0_u7_n6 ) , .ZN( u0_u0_u7_n67 ) , .A2( u0_u0_u7_n69 ) );
  NOR2_X1 u0_u0_u7_U44 (.A2( u0_u0_u7_n20 ) , .A1( u0_u0_u7_n31 ) , .ZN( u0_u0_u7_n44 ) );
  AND2_X1 u0_u0_u7_U45 (.ZN( u0_u0_u7_n36 ) , .A1( u0_u0_u7_n82 ) , .A2( u0_u0_u7_n83 ) );
  AOI21_X1 u0_u0_u7_U46 (.B1( u0_u0_u7_n34 ) , .A( u0_u0_u7_n56 ) , .B2( u0_u0_u7_n71 ) , .ZN( u0_u0_u7_n76 ) );
  NAND2_X1 u0_u0_u7_U47 (.ZN( u0_u0_u7_n35 ) , .A2( u0_u0_u7_n83 ) , .A1( u0_u0_u7_n86 ) );
  NAND2_X1 u0_u0_u7_U48 (.ZN( u0_u0_u7_n34 ) , .A2( u0_u0_u7_n78 ) , .A1( u0_u0_u7_n88 ) );
  NAND2_X1 u0_u0_u7_U49 (.ZN( u0_u0_u7_n54 ) , .A1( u0_u0_u7_n78 ) , .A2( u0_u0_u7_n82 ) );
  INV_X1 u0_u0_u7_U5 (.A( u0_u0_u7_n27 ) , .ZN( u0_u0_u7_n3 ) );
  NAND2_X1 u0_u0_u7_U50 (.ZN( u0_u0_u7_n48 ) , .A1( u0_u0_u7_n78 ) , .A2( u0_u0_u7_n79 ) );
  OR2_X1 u0_u0_u7_U51 (.A1( u0_u0_u7_n25 ) , .A2( u0_u0_u7_n29 ) , .ZN( u0_u0_u7_n55 ) );
  NAND2_X1 u0_u0_u7_U52 (.ZN( u0_u0_u7_n69 ) , .A1( u0_u0_u7_n82 ) , .A2( u0_u0_u7_n85 ) );
  NAND2_X1 u0_u0_u7_U53 (.ZN( u0_u0_u7_n53 ) , .A2( u0_u0_u7_n79 ) , .A1( u0_u0_u7_n83 ) );
  NAND2_X1 u0_u0_u7_U54 (.ZN( u0_u0_u7_n68 ) , .A1( u0_u0_u7_n81 ) , .A2( u0_u0_u7_n88 ) );
  NAND2_X1 u0_u0_u7_U55 (.ZN( u0_u0_u7_n71 ) , .A2( u0_u0_u7_n85 ) , .A1( u0_u0_u7_n86 ) );
  INV_X1 u0_u0_u7_U56 (.ZN( u0_u0_u7_n17 ) , .A( u0_u0_u7_n31 ) );
  AND2_X1 u0_u0_u7_U57 (.ZN( u0_u0_u7_n47 ) , .A2( u0_u0_u7_n83 ) , .A1( u0_u0_u7_n88 ) );
  NAND2_X1 u0_u0_u7_U58 (.ZN( u0_u0_u7_n57 ) , .A2( u0_u0_u7_n79 ) , .A1( u0_u0_u7_n85 ) );
  NAND2_X1 u0_u0_u7_U59 (.ZN( u0_u0_u7_n52 ) , .A2( u0_u0_u7_n79 ) , .A1( u0_u0_u7_n81 ) );
  AOI211_X1 u0_u0_u7_U6 (.C2( u0_u0_u7_n10 ) , .C1( u0_u0_u7_n20 ) , .A( u0_u0_u7_n26 ) , .ZN( u0_u0_u7_n65 ) , .B( u0_u0_u7_n87 ) );
  NAND2_X1 u0_u0_u7_U60 (.ZN( u0_u0_u7_n50 ) , .A2( u0_u0_u7_n78 ) , .A1( u0_u0_u7_n86 ) );
  NAND2_X1 u0_u0_u7_U61 (.ZN( u0_u0_u7_n43 ) , .A1( u0_u0_u7_n81 ) , .A2( u0_u0_u7_n82 ) );
  NAND2_X1 u0_u0_u7_U62 (.ZN( u0_u0_u7_n49 ) , .A2( u0_u0_u7_n85 ) , .A1( u0_u0_u7_n88 ) );
  NAND2_X1 u0_u0_u7_U63 (.ZN( u0_u0_u7_n33 ) , .A1( u0_u0_u7_n81 ) , .A2( u0_u0_u7_n86 ) );
  NOR2_X1 u0_u0_u7_U64 (.A2( u0_u0_X_47 ) , .A1( u0_u0_u7_n18 ) , .ZN( u0_u0_u7_n31 ) );
  NOR2_X1 u0_u0_u7_U65 (.A2( u0_u0_X_43 ) , .A1( u0_u0_X_44 ) , .ZN( u0_u0_u7_n78 ) );
  NOR2_X1 u0_u0_u7_U66 (.A2( u0_u0_X_48 ) , .A1( u0_u0_u7_n15 ) , .ZN( u0_u0_u7_n86 ) );
  NOR2_X1 u0_u0_u7_U67 (.A2( u0_u0_X_45 ) , .A1( u0_u0_X_48 ) , .ZN( u0_u0_u7_n82 ) );
  NOR2_X1 u0_u0_u7_U68 (.A2( u0_u0_X_44 ) , .A1( u0_u0_u7_n14 ) , .ZN( u0_u0_u7_n83 ) );
  NOR2_X1 u0_u0_u7_U69 (.A2( u0_u0_X_46 ) , .A1( u0_u0_X_47 ) , .ZN( u0_u0_u7_n29 ) );
  OAI222_X1 u0_u0_u7_U7 (.B1( u0_u0_u7_n17 ) , .A2( u0_u0_u7_n19 ) , .C1( u0_u0_u7_n35 ) , .A1( u0_u0_u7_n68 ) , .B2( u0_u0_u7_n70 ) , .C2( u0_u0_u7_n80 ) , .ZN( u0_u0_u7_n87 ) );
  NAND2_X1 u0_u0_u7_U70 (.A2( u0_u0_X_46 ) , .A1( u0_u0_X_47 ) , .ZN( u0_u0_u7_n56 ) );
  AND2_X1 u0_u0_u7_U71 (.A1( u0_u0_X_47 ) , .A2( u0_u0_u7_n18 ) , .ZN( u0_u0_u7_n25 ) );
  AND2_X1 u0_u0_u7_U72 (.A2( u0_u0_X_45 ) , .A1( u0_u0_X_48 ) , .ZN( u0_u0_u7_n79 ) );
  AND2_X1 u0_u0_u7_U73 (.A2( u0_u0_X_43 ) , .A1( u0_u0_X_44 ) , .ZN( u0_u0_u7_n85 ) );
  AND2_X1 u0_u0_u7_U74 (.A1( u0_u0_X_44 ) , .A2( u0_u0_u7_n14 ) , .ZN( u0_u0_u7_n81 ) );
  AND2_X1 u0_u0_u7_U75 (.A1( u0_u0_X_48 ) , .A2( u0_u0_u7_n15 ) , .ZN( u0_u0_u7_n88 ) );
  INV_X1 u0_u0_u7_U76 (.A( u0_u0_X_46 ) , .ZN( u0_u0_u7_n18 ) );
  INV_X1 u0_u0_u7_U77 (.A( u0_u0_X_45 ) , .ZN( u0_u0_u7_n15 ) );
  NAND4_X1 u0_u0_u7_U78 (.ZN( u0_out0_27 ) , .A1( u0_u0_u7_n60 ) , .A2( u0_u0_u7_n61 ) , .A3( u0_u0_u7_n62 ) , .A4( u0_u0_u7_n63 ) );
  OAI21_X1 u0_u0_u7_U79 (.A( u0_u0_u7_n31 ) , .B2( u0_u0_u7_n36 ) , .ZN( u0_u0_u7_n60 ) , .B1( u0_u0_u7_n7 ) );
  OAI221_X1 u0_u0_u7_U8 (.B2( u0_u0_u7_n19 ) , .ZN( u0_u0_u7_n26 ) , .C2( u0_u0_u7_n34 ) , .C1( u0_u0_u7_n80 ) , .B1( u0_u0_u7_n89 ) , .A( u0_u0_u7_n90 ) );
  OAI21_X1 u0_u0_u7_U80 (.B2( u0_u0_u7_n11 ) , .B1( u0_u0_u7_n2 ) , .A( u0_u0_u7_n20 ) , .ZN( u0_u0_u7_n61 ) );
  NAND4_X1 u0_u0_u7_U81 (.ZN( u0_out0_21 ) , .A1( u0_u0_u7_n21 ) , .A2( u0_u0_u7_n22 ) , .A3( u0_u0_u7_n23 ) , .A4( u0_u0_u7_n24 ) );
  OAI21_X1 u0_u0_u7_U82 (.A( u0_u0_u7_n20 ) , .ZN( u0_u0_u7_n21 ) , .B1( u0_u0_u7_n36 ) , .B2( u0_u0_u7_n4 ) );
  AOI22_X1 u0_u0_u7_U83 (.ZN( u0_u0_u7_n23 ) , .A1( u0_u0_u7_n29 ) , .A2( u0_u0_u7_n30 ) , .B1( u0_u0_u7_n31 ) , .B2( u0_u0_u7_n32 ) );
  NAND4_X1 u0_u0_u7_U84 (.ZN( u0_out0_5 ) , .A2( u0_u0_u7_n58 ) , .A1( u0_u0_u7_n65 ) , .A3( u0_u0_u7_n72 ) , .A4( u0_u0_u7_n73 ) );
  AOI22_X1 u0_u0_u7_U85 (.A1( u0_u0_u7_n10 ) , .B1( u0_u0_u7_n25 ) , .B2( u0_u0_u7_n36 ) , .A2( u0_u0_u7_n55 ) , .ZN( u0_u0_u7_n72 ) );
  NOR4_X1 u0_u0_u7_U86 (.ZN( u0_u0_u7_n73 ) , .A1( u0_u0_u7_n74 ) , .A2( u0_u0_u7_n75 ) , .A3( u0_u0_u7_n76 ) , .A4( u0_u0_u7_n77 ) );
  NAND4_X1 u0_u0_u7_U87 (.ZN( u0_out0_15 ) , .A1( u0_u0_u7_n3 ) , .A2( u0_u0_u7_n37 ) , .A3( u0_u0_u7_n38 ) , .A4( u0_u0_u7_n39 ) );
  OR2_X1 u0_u0_u7_U88 (.ZN( u0_u0_u7_n37 ) , .A1( u0_u0_u7_n52 ) , .A2( u0_u0_u7_n56 ) );
  AOI22_X1 u0_u0_u7_U89 (.B2( u0_u0_u7_n16 ) , .ZN( u0_u0_u7_n38 ) , .A2( u0_u0_u7_n55 ) , .A1( u0_u0_u7_n7 ) , .B1( u0_u0_u7_n8 ) );
  AND3_X1 u0_u0_u7_U9 (.A1( u0_u0_u7_n49 ) , .A2( u0_u0_u7_n54 ) , .A3( u0_u0_u7_n71 ) , .ZN( u0_u0_u7_n89 ) );
  INV_X1 u0_u0_u7_U90 (.A( u0_u0_X_43 ) , .ZN( u0_u0_u7_n14 ) );
  AOI211_X1 u0_u0_u7_U91 (.ZN( u0_u0_u7_n24 ) , .C1( u0_u0_u7_n25 ) , .A( u0_u0_u7_n26 ) , .B( u0_u0_u7_n27 ) , .C2( u0_u0_u7_n9 ) );
  OAI211_X1 u0_u0_u7_U92 (.C1( u0_u0_u7_n19 ) , .ZN( u0_u0_u7_n27 ) , .C2( u0_u0_u7_n57 ) , .A( u0_u0_u7_n58 ) , .B( u0_u0_u7_n59 ) );
  AOI222_X1 u0_u0_u7_U93 (.B2( u0_u0_u7_n11 ) , .A2( u0_u0_u7_n16 ) , .B1( u0_u0_u7_n20 ) , .C1( u0_u0_u7_n36 ) , .A1( u0_u0_u7_n5 ) , .C2( u0_u0_u7_n55 ) , .ZN( u0_u0_u7_n59 ) );
  INV_X1 u0_u0_u7_U94 (.ZN( u0_u0_u7_n11 ) , .A( u0_u0_u7_n70 ) );
  NAND3_X1 u0_u0_u7_U95 (.ZN( u0_u0_u7_n30 ) , .A1( u0_u0_u7_n33 ) , .A2( u0_u0_u7_n34 ) , .A3( u0_u0_u7_n35 ) );
  NAND3_X1 u0_u0_u7_U96 (.ZN( u0_u0_u7_n46 ) , .A1( u0_u0_u7_n48 ) , .A2( u0_u0_u7_n49 ) , .A3( u0_u0_u7_n50 ) );
  XOR2_X1 u0_u11_U1 (.B( u0_K12_9 ) , .A( u0_R10_6 ) , .Z( u0_u11_X_9 ) );
  XOR2_X1 u0_u11_U16 (.B( u0_K12_3 ) , .A( u0_R10_2 ) , .Z( u0_u11_X_3 ) );
  XOR2_X1 u0_u11_U2 (.B( u0_K12_8 ) , .A( u0_R10_5 ) , .Z( u0_u11_X_8 ) );
  XOR2_X1 u0_u11_U27 (.B( u0_K12_2 ) , .A( u0_R10_1 ) , .Z( u0_u11_X_2 ) );
  XOR2_X1 u0_u11_U3 (.B( u0_K12_7 ) , .A( u0_R10_4 ) , .Z( u0_u11_X_7 ) );
  XOR2_X1 u0_u11_U33 (.B( u0_K12_24 ) , .A( u0_R10_17 ) , .Z( u0_u11_X_24 ) );
  XOR2_X1 u0_u11_U34 (.B( u0_K12_23 ) , .A( u0_R10_16 ) , .Z( u0_u11_X_23 ) );
  XOR2_X1 u0_u11_U35 (.B( u0_K12_22 ) , .A( u0_R10_15 ) , .Z( u0_u11_X_22 ) );
  XOR2_X1 u0_u11_U36 (.B( u0_K12_21 ) , .A( u0_R10_14 ) , .Z( u0_u11_X_21 ) );
  XOR2_X1 u0_u11_U37 (.B( u0_K12_20 ) , .A( u0_R10_13 ) , .Z( u0_u11_X_20 ) );
  XOR2_X1 u0_u11_U38 (.B( u0_K12_1 ) , .A( u0_R10_32 ) , .Z( u0_u11_X_1 ) );
  XOR2_X1 u0_u11_U39 (.B( u0_K12_19 ) , .A( u0_R10_12 ) , .Z( u0_u11_X_19 ) );
  XOR2_X1 u0_u11_U4 (.B( u0_K12_6 ) , .A( u0_R10_5 ) , .Z( u0_u11_X_6 ) );
  XOR2_X1 u0_u11_U40 (.B( u0_K12_18 ) , .A( u0_R10_13 ) , .Z( u0_u11_X_18 ) );
  XOR2_X1 u0_u11_U41 (.B( u0_K12_17 ) , .A( u0_R10_12 ) , .Z( u0_u11_X_17 ) );
  XOR2_X1 u0_u11_U42 (.B( u0_K12_16 ) , .A( u0_R10_11 ) , .Z( u0_u11_X_16 ) );
  XOR2_X1 u0_u11_U43 (.B( u0_K12_15 ) , .A( u0_R10_10 ) , .Z( u0_u11_X_15 ) );
  XOR2_X1 u0_u11_U44 (.B( u0_K12_14 ) , .A( u0_R10_9 ) , .Z( u0_u11_X_14 ) );
  XOR2_X1 u0_u11_U45 (.B( u0_K12_13 ) , .A( u0_R10_8 ) , .Z( u0_u11_X_13 ) );
  XOR2_X1 u0_u11_U46 (.B( u0_K12_12 ) , .A( u0_R10_9 ) , .Z( u0_u11_X_12 ) );
  XOR2_X1 u0_u11_U47 (.B( u0_K12_11 ) , .A( u0_R10_8 ) , .Z( u0_u11_X_11 ) );
  XOR2_X1 u0_u11_U48 (.B( u0_K12_10 ) , .A( u0_R10_7 ) , .Z( u0_u11_X_10 ) );
  XOR2_X1 u0_u11_U5 (.B( u0_K12_5 ) , .A( u0_R10_4 ) , .Z( u0_u11_X_5 ) );
  XOR2_X1 u0_u11_U6 (.B( u0_K12_4 ) , .A( u0_R10_3 ) , .Z( u0_u11_X_4 ) );
  AND3_X1 u0_u11_u0_U10 (.A2( u0_u11_u0_n112 ) , .ZN( u0_u11_u0_n127 ) , .A3( u0_u11_u0_n130 ) , .A1( u0_u11_u0_n148 ) );
  NAND2_X1 u0_u11_u0_U11 (.ZN( u0_u11_u0_n113 ) , .A1( u0_u11_u0_n139 ) , .A2( u0_u11_u0_n149 ) );
  AND2_X1 u0_u11_u0_U12 (.ZN( u0_u11_u0_n107 ) , .A1( u0_u11_u0_n130 ) , .A2( u0_u11_u0_n140 ) );
  AND2_X1 u0_u11_u0_U13 (.A2( u0_u11_u0_n129 ) , .A1( u0_u11_u0_n130 ) , .ZN( u0_u11_u0_n151 ) );
  AND2_X1 u0_u11_u0_U14 (.A1( u0_u11_u0_n108 ) , .A2( u0_u11_u0_n125 ) , .ZN( u0_u11_u0_n145 ) );
  INV_X1 u0_u11_u0_U15 (.A( u0_u11_u0_n143 ) , .ZN( u0_u11_u0_n173 ) );
  NOR2_X1 u0_u11_u0_U16 (.A2( u0_u11_u0_n136 ) , .ZN( u0_u11_u0_n147 ) , .A1( u0_u11_u0_n160 ) );
  AOI21_X1 u0_u11_u0_U17 (.B1( u0_u11_u0_n103 ) , .ZN( u0_u11_u0_n132 ) , .A( u0_u11_u0_n165 ) , .B2( u0_u11_u0_n93 ) );
  INV_X1 u0_u11_u0_U18 (.A( u0_u11_u0_n142 ) , .ZN( u0_u11_u0_n165 ) );
  OAI22_X1 u0_u11_u0_U19 (.B1( u0_u11_u0_n125 ) , .ZN( u0_u11_u0_n126 ) , .A1( u0_u11_u0_n138 ) , .A2( u0_u11_u0_n146 ) , .B2( u0_u11_u0_n147 ) );
  OAI22_X1 u0_u11_u0_U20 (.B1( u0_u11_u0_n131 ) , .A1( u0_u11_u0_n144 ) , .B2( u0_u11_u0_n147 ) , .A2( u0_u11_u0_n90 ) , .ZN( u0_u11_u0_n91 ) );
  AND3_X1 u0_u11_u0_U21 (.A3( u0_u11_u0_n121 ) , .A2( u0_u11_u0_n125 ) , .A1( u0_u11_u0_n148 ) , .ZN( u0_u11_u0_n90 ) );
  INV_X1 u0_u11_u0_U22 (.A( u0_u11_u0_n136 ) , .ZN( u0_u11_u0_n161 ) );
  AOI22_X1 u0_u11_u0_U23 (.B2( u0_u11_u0_n109 ) , .A2( u0_u11_u0_n110 ) , .ZN( u0_u11_u0_n111 ) , .B1( u0_u11_u0_n118 ) , .A1( u0_u11_u0_n160 ) );
  NAND2_X1 u0_u11_u0_U24 (.A1( u0_u11_u0_n100 ) , .A2( u0_u11_u0_n103 ) , .ZN( u0_u11_u0_n125 ) );
  INV_X1 u0_u11_u0_U25 (.A( u0_u11_u0_n118 ) , .ZN( u0_u11_u0_n158 ) );
  AOI21_X1 u0_u11_u0_U26 (.B1( u0_u11_u0_n127 ) , .B2( u0_u11_u0_n129 ) , .A( u0_u11_u0_n138 ) , .ZN( u0_u11_u0_n96 ) );
  AOI21_X1 u0_u11_u0_U27 (.ZN( u0_u11_u0_n104 ) , .B1( u0_u11_u0_n107 ) , .B2( u0_u11_u0_n141 ) , .A( u0_u11_u0_n144 ) );
  AOI21_X1 u0_u11_u0_U28 (.ZN( u0_u11_u0_n116 ) , .B2( u0_u11_u0_n142 ) , .A( u0_u11_u0_n144 ) , .B1( u0_u11_u0_n166 ) );
  NOR2_X1 u0_u11_u0_U29 (.A1( u0_u11_u0_n120 ) , .ZN( u0_u11_u0_n143 ) , .A2( u0_u11_u0_n167 ) );
  INV_X1 u0_u11_u0_U3 (.A( u0_u11_u0_n113 ) , .ZN( u0_u11_u0_n166 ) );
  OAI221_X1 u0_u11_u0_U30 (.C1( u0_u11_u0_n112 ) , .ZN( u0_u11_u0_n120 ) , .B1( u0_u11_u0_n138 ) , .B2( u0_u11_u0_n141 ) , .C2( u0_u11_u0_n147 ) , .A( u0_u11_u0_n172 ) );
  AOI211_X1 u0_u11_u0_U31 (.B( u0_u11_u0_n115 ) , .A( u0_u11_u0_n116 ) , .C2( u0_u11_u0_n117 ) , .C1( u0_u11_u0_n118 ) , .ZN( u0_u11_u0_n119 ) );
  NAND2_X1 u0_u11_u0_U32 (.A2( u0_u11_u0_n103 ) , .ZN( u0_u11_u0_n140 ) , .A1( u0_u11_u0_n94 ) );
  NAND2_X1 u0_u11_u0_U33 (.A1( u0_u11_u0_n101 ) , .A2( u0_u11_u0_n102 ) , .ZN( u0_u11_u0_n150 ) );
  INV_X1 u0_u11_u0_U34 (.A( u0_u11_u0_n138 ) , .ZN( u0_u11_u0_n160 ) );
  NAND2_X1 u0_u11_u0_U35 (.A2( u0_u11_u0_n100 ) , .A1( u0_u11_u0_n101 ) , .ZN( u0_u11_u0_n139 ) );
  NAND2_X1 u0_u11_u0_U36 (.A2( u0_u11_u0_n100 ) , .ZN( u0_u11_u0_n131 ) , .A1( u0_u11_u0_n92 ) );
  NAND2_X1 u0_u11_u0_U37 (.A2( u0_u11_u0_n102 ) , .A1( u0_u11_u0_n103 ) , .ZN( u0_u11_u0_n149 ) );
  NAND2_X1 u0_u11_u0_U38 (.ZN( u0_u11_u0_n108 ) , .A1( u0_u11_u0_n92 ) , .A2( u0_u11_u0_n94 ) );
  NAND2_X1 u0_u11_u0_U39 (.A2( u0_u11_u0_n102 ) , .ZN( u0_u11_u0_n114 ) , .A1( u0_u11_u0_n92 ) );
  AOI21_X1 u0_u11_u0_U4 (.B1( u0_u11_u0_n114 ) , .ZN( u0_u11_u0_n115 ) , .B2( u0_u11_u0_n129 ) , .A( u0_u11_u0_n161 ) );
  NAND2_X1 u0_u11_u0_U40 (.A1( u0_u11_u0_n101 ) , .ZN( u0_u11_u0_n130 ) , .A2( u0_u11_u0_n94 ) );
  INV_X1 u0_u11_u0_U41 (.ZN( u0_u11_u0_n172 ) , .A( u0_u11_u0_n88 ) );
  OAI222_X1 u0_u11_u0_U42 (.C1( u0_u11_u0_n108 ) , .A1( u0_u11_u0_n125 ) , .B2( u0_u11_u0_n128 ) , .B1( u0_u11_u0_n144 ) , .A2( u0_u11_u0_n158 ) , .C2( u0_u11_u0_n161 ) , .ZN( u0_u11_u0_n88 ) );
  NAND2_X1 u0_u11_u0_U43 (.ZN( u0_u11_u0_n112 ) , .A2( u0_u11_u0_n92 ) , .A1( u0_u11_u0_n93 ) );
  NAND2_X1 u0_u11_u0_U44 (.A2( u0_u11_u0_n101 ) , .ZN( u0_u11_u0_n121 ) , .A1( u0_u11_u0_n93 ) );
  OR3_X1 u0_u11_u0_U45 (.A3( u0_u11_u0_n152 ) , .A2( u0_u11_u0_n153 ) , .A1( u0_u11_u0_n154 ) , .ZN( u0_u11_u0_n155 ) );
  AOI21_X1 u0_u11_u0_U46 (.A( u0_u11_u0_n144 ) , .B2( u0_u11_u0_n145 ) , .B1( u0_u11_u0_n146 ) , .ZN( u0_u11_u0_n154 ) );
  AOI21_X1 u0_u11_u0_U47 (.B2( u0_u11_u0_n150 ) , .B1( u0_u11_u0_n151 ) , .ZN( u0_u11_u0_n152 ) , .A( u0_u11_u0_n158 ) );
  AOI21_X1 u0_u11_u0_U48 (.A( u0_u11_u0_n147 ) , .B2( u0_u11_u0_n148 ) , .B1( u0_u11_u0_n149 ) , .ZN( u0_u11_u0_n153 ) );
  INV_X1 u0_u11_u0_U49 (.ZN( u0_u11_u0_n171 ) , .A( u0_u11_u0_n99 ) );
  AOI21_X1 u0_u11_u0_U5 (.B2( u0_u11_u0_n131 ) , .ZN( u0_u11_u0_n134 ) , .B1( u0_u11_u0_n151 ) , .A( u0_u11_u0_n158 ) );
  OAI211_X1 u0_u11_u0_U50 (.C2( u0_u11_u0_n140 ) , .C1( u0_u11_u0_n161 ) , .A( u0_u11_u0_n169 ) , .B( u0_u11_u0_n98 ) , .ZN( u0_u11_u0_n99 ) );
  AOI211_X1 u0_u11_u0_U51 (.C1( u0_u11_u0_n118 ) , .A( u0_u11_u0_n123 ) , .B( u0_u11_u0_n96 ) , .C2( u0_u11_u0_n97 ) , .ZN( u0_u11_u0_n98 ) );
  INV_X1 u0_u11_u0_U52 (.ZN( u0_u11_u0_n169 ) , .A( u0_u11_u0_n91 ) );
  NOR2_X1 u0_u11_u0_U53 (.A2( u0_u11_X_2 ) , .ZN( u0_u11_u0_n103 ) , .A1( u0_u11_u0_n164 ) );
  NOR2_X1 u0_u11_u0_U54 (.A2( u0_u11_X_4 ) , .A1( u0_u11_X_5 ) , .ZN( u0_u11_u0_n118 ) );
  NOR2_X1 u0_u11_u0_U55 (.A2( u0_u11_X_1 ) , .A1( u0_u11_X_2 ) , .ZN( u0_u11_u0_n92 ) );
  NOR2_X1 u0_u11_u0_U56 (.A2( u0_u11_X_1 ) , .ZN( u0_u11_u0_n101 ) , .A1( u0_u11_u0_n163 ) );
  NOR2_X1 u0_u11_u0_U57 (.A2( u0_u11_X_3 ) , .A1( u0_u11_X_6 ) , .ZN( u0_u11_u0_n94 ) );
  NAND2_X1 u0_u11_u0_U58 (.A2( u0_u11_X_4 ) , .A1( u0_u11_X_5 ) , .ZN( u0_u11_u0_n144 ) );
  NOR2_X1 u0_u11_u0_U59 (.A2( u0_u11_X_5 ) , .ZN( u0_u11_u0_n136 ) , .A1( u0_u11_u0_n159 ) );
  NOR2_X1 u0_u11_u0_U6 (.A1( u0_u11_u0_n108 ) , .ZN( u0_u11_u0_n123 ) , .A2( u0_u11_u0_n158 ) );
  NAND2_X1 u0_u11_u0_U60 (.A1( u0_u11_X_5 ) , .ZN( u0_u11_u0_n138 ) , .A2( u0_u11_u0_n159 ) );
  AND2_X1 u0_u11_u0_U61 (.A2( u0_u11_X_3 ) , .A1( u0_u11_X_6 ) , .ZN( u0_u11_u0_n102 ) );
  AND2_X1 u0_u11_u0_U62 (.A1( u0_u11_X_6 ) , .A2( u0_u11_u0_n162 ) , .ZN( u0_u11_u0_n93 ) );
  INV_X1 u0_u11_u0_U63 (.A( u0_u11_X_4 ) , .ZN( u0_u11_u0_n159 ) );
  INV_X1 u0_u11_u0_U64 (.A( u0_u11_X_2 ) , .ZN( u0_u11_u0_n163 ) );
  INV_X1 u0_u11_u0_U65 (.A( u0_u11_X_1 ) , .ZN( u0_u11_u0_n164 ) );
  INV_X1 u0_u11_u0_U66 (.A( u0_u11_u0_n126 ) , .ZN( u0_u11_u0_n168 ) );
  AOI211_X1 u0_u11_u0_U67 (.B( u0_u11_u0_n133 ) , .A( u0_u11_u0_n134 ) , .C2( u0_u11_u0_n135 ) , .C1( u0_u11_u0_n136 ) , .ZN( u0_u11_u0_n137 ) );
  OR4_X1 u0_u11_u0_U68 (.ZN( u0_out11_17 ) , .A4( u0_u11_u0_n122 ) , .A2( u0_u11_u0_n123 ) , .A1( u0_u11_u0_n124 ) , .A3( u0_u11_u0_n170 ) );
  AOI21_X1 u0_u11_u0_U69 (.B2( u0_u11_u0_n107 ) , .ZN( u0_u11_u0_n124 ) , .B1( u0_u11_u0_n128 ) , .A( u0_u11_u0_n161 ) );
  OAI21_X1 u0_u11_u0_U7 (.B1( u0_u11_u0_n150 ) , .B2( u0_u11_u0_n158 ) , .A( u0_u11_u0_n172 ) , .ZN( u0_u11_u0_n89 ) );
  INV_X1 u0_u11_u0_U70 (.A( u0_u11_u0_n111 ) , .ZN( u0_u11_u0_n170 ) );
  OR4_X1 u0_u11_u0_U71 (.ZN( u0_out11_31 ) , .A4( u0_u11_u0_n155 ) , .A2( u0_u11_u0_n156 ) , .A1( u0_u11_u0_n157 ) , .A3( u0_u11_u0_n173 ) );
  AOI21_X1 u0_u11_u0_U72 (.A( u0_u11_u0_n138 ) , .B2( u0_u11_u0_n139 ) , .B1( u0_u11_u0_n140 ) , .ZN( u0_u11_u0_n157 ) );
  AOI21_X1 u0_u11_u0_U73 (.B2( u0_u11_u0_n141 ) , .B1( u0_u11_u0_n142 ) , .ZN( u0_u11_u0_n156 ) , .A( u0_u11_u0_n161 ) );
  INV_X1 u0_u11_u0_U74 (.ZN( u0_u11_u0_n174 ) , .A( u0_u11_u0_n89 ) );
  AOI211_X1 u0_u11_u0_U75 (.B( u0_u11_u0_n104 ) , .A( u0_u11_u0_n105 ) , .ZN( u0_u11_u0_n106 ) , .C2( u0_u11_u0_n113 ) , .C1( u0_u11_u0_n160 ) );
  NOR2_X1 u0_u11_u0_U76 (.A2( u0_u11_X_6 ) , .ZN( u0_u11_u0_n100 ) , .A1( u0_u11_u0_n162 ) );
  INV_X1 u0_u11_u0_U77 (.A( u0_u11_X_3 ) , .ZN( u0_u11_u0_n162 ) );
  NOR2_X1 u0_u11_u0_U78 (.A1( u0_u11_u0_n163 ) , .A2( u0_u11_u0_n164 ) , .ZN( u0_u11_u0_n95 ) );
  OAI221_X1 u0_u11_u0_U79 (.C1( u0_u11_u0_n121 ) , .ZN( u0_u11_u0_n122 ) , .B2( u0_u11_u0_n127 ) , .A( u0_u11_u0_n143 ) , .B1( u0_u11_u0_n144 ) , .C2( u0_u11_u0_n147 ) );
  AND2_X1 u0_u11_u0_U8 (.A1( u0_u11_u0_n114 ) , .A2( u0_u11_u0_n121 ) , .ZN( u0_u11_u0_n146 ) );
  AOI21_X1 u0_u11_u0_U80 (.B1( u0_u11_u0_n132 ) , .ZN( u0_u11_u0_n133 ) , .A( u0_u11_u0_n144 ) , .B2( u0_u11_u0_n166 ) );
  OAI22_X1 u0_u11_u0_U81 (.ZN( u0_u11_u0_n105 ) , .A2( u0_u11_u0_n132 ) , .B1( u0_u11_u0_n146 ) , .A1( u0_u11_u0_n147 ) , .B2( u0_u11_u0_n161 ) );
  NAND2_X1 u0_u11_u0_U82 (.ZN( u0_u11_u0_n110 ) , .A2( u0_u11_u0_n132 ) , .A1( u0_u11_u0_n145 ) );
  INV_X1 u0_u11_u0_U83 (.A( u0_u11_u0_n119 ) , .ZN( u0_u11_u0_n167 ) );
  NAND2_X1 u0_u11_u0_U84 (.ZN( u0_u11_u0_n148 ) , .A1( u0_u11_u0_n93 ) , .A2( u0_u11_u0_n95 ) );
  NAND2_X1 u0_u11_u0_U85 (.A1( u0_u11_u0_n100 ) , .ZN( u0_u11_u0_n129 ) , .A2( u0_u11_u0_n95 ) );
  NAND2_X1 u0_u11_u0_U86 (.A1( u0_u11_u0_n102 ) , .ZN( u0_u11_u0_n128 ) , .A2( u0_u11_u0_n95 ) );
  NAND2_X1 u0_u11_u0_U87 (.ZN( u0_u11_u0_n142 ) , .A1( u0_u11_u0_n94 ) , .A2( u0_u11_u0_n95 ) );
  NAND3_X1 u0_u11_u0_U88 (.ZN( u0_out11_23 ) , .A3( u0_u11_u0_n137 ) , .A1( u0_u11_u0_n168 ) , .A2( u0_u11_u0_n171 ) );
  NAND3_X1 u0_u11_u0_U89 (.A3( u0_u11_u0_n127 ) , .A2( u0_u11_u0_n128 ) , .ZN( u0_u11_u0_n135 ) , .A1( u0_u11_u0_n150 ) );
  AND2_X1 u0_u11_u0_U9 (.A1( u0_u11_u0_n131 ) , .ZN( u0_u11_u0_n141 ) , .A2( u0_u11_u0_n150 ) );
  NAND3_X1 u0_u11_u0_U90 (.ZN( u0_u11_u0_n117 ) , .A3( u0_u11_u0_n132 ) , .A2( u0_u11_u0_n139 ) , .A1( u0_u11_u0_n148 ) );
  NAND3_X1 u0_u11_u0_U91 (.ZN( u0_u11_u0_n109 ) , .A2( u0_u11_u0_n114 ) , .A3( u0_u11_u0_n140 ) , .A1( u0_u11_u0_n149 ) );
  NAND3_X1 u0_u11_u0_U92 (.ZN( u0_out11_9 ) , .A3( u0_u11_u0_n106 ) , .A2( u0_u11_u0_n171 ) , .A1( u0_u11_u0_n174 ) );
  NAND3_X1 u0_u11_u0_U93 (.A2( u0_u11_u0_n128 ) , .A1( u0_u11_u0_n132 ) , .A3( u0_u11_u0_n146 ) , .ZN( u0_u11_u0_n97 ) );
  NOR2_X1 u0_u11_u1_U10 (.A1( u0_u11_u1_n112 ) , .A2( u0_u11_u1_n116 ) , .ZN( u0_u11_u1_n118 ) );
  NAND3_X1 u0_u11_u1_U100 (.ZN( u0_u11_u1_n113 ) , .A1( u0_u11_u1_n120 ) , .A3( u0_u11_u1_n133 ) , .A2( u0_u11_u1_n155 ) );
  OAI21_X1 u0_u11_u1_U11 (.ZN( u0_u11_u1_n101 ) , .B1( u0_u11_u1_n141 ) , .A( u0_u11_u1_n146 ) , .B2( u0_u11_u1_n183 ) );
  AOI21_X1 u0_u11_u1_U12 (.B2( u0_u11_u1_n155 ) , .B1( u0_u11_u1_n156 ) , .ZN( u0_u11_u1_n157 ) , .A( u0_u11_u1_n174 ) );
  NAND2_X1 u0_u11_u1_U13 (.ZN( u0_u11_u1_n140 ) , .A2( u0_u11_u1_n150 ) , .A1( u0_u11_u1_n155 ) );
  NAND2_X1 u0_u11_u1_U14 (.A1( u0_u11_u1_n131 ) , .ZN( u0_u11_u1_n147 ) , .A2( u0_u11_u1_n153 ) );
  INV_X1 u0_u11_u1_U15 (.A( u0_u11_u1_n139 ) , .ZN( u0_u11_u1_n174 ) );
  OR4_X1 u0_u11_u1_U16 (.A4( u0_u11_u1_n106 ) , .A3( u0_u11_u1_n107 ) , .ZN( u0_u11_u1_n108 ) , .A1( u0_u11_u1_n117 ) , .A2( u0_u11_u1_n184 ) );
  AOI21_X1 u0_u11_u1_U17 (.ZN( u0_u11_u1_n106 ) , .A( u0_u11_u1_n112 ) , .B1( u0_u11_u1_n154 ) , .B2( u0_u11_u1_n156 ) );
  AOI21_X1 u0_u11_u1_U18 (.ZN( u0_u11_u1_n107 ) , .B1( u0_u11_u1_n134 ) , .B2( u0_u11_u1_n149 ) , .A( u0_u11_u1_n174 ) );
  INV_X1 u0_u11_u1_U19 (.A( u0_u11_u1_n101 ) , .ZN( u0_u11_u1_n184 ) );
  INV_X1 u0_u11_u1_U20 (.A( u0_u11_u1_n112 ) , .ZN( u0_u11_u1_n171 ) );
  NAND2_X1 u0_u11_u1_U21 (.ZN( u0_u11_u1_n141 ) , .A1( u0_u11_u1_n153 ) , .A2( u0_u11_u1_n156 ) );
  AND2_X1 u0_u11_u1_U22 (.A1( u0_u11_u1_n123 ) , .ZN( u0_u11_u1_n134 ) , .A2( u0_u11_u1_n161 ) );
  NAND2_X1 u0_u11_u1_U23 (.A2( u0_u11_u1_n115 ) , .A1( u0_u11_u1_n116 ) , .ZN( u0_u11_u1_n148 ) );
  NAND2_X1 u0_u11_u1_U24 (.A2( u0_u11_u1_n133 ) , .A1( u0_u11_u1_n135 ) , .ZN( u0_u11_u1_n159 ) );
  NAND2_X1 u0_u11_u1_U25 (.A2( u0_u11_u1_n115 ) , .A1( u0_u11_u1_n120 ) , .ZN( u0_u11_u1_n132 ) );
  INV_X1 u0_u11_u1_U26 (.A( u0_u11_u1_n154 ) , .ZN( u0_u11_u1_n178 ) );
  INV_X1 u0_u11_u1_U27 (.A( u0_u11_u1_n151 ) , .ZN( u0_u11_u1_n183 ) );
  AND2_X1 u0_u11_u1_U28 (.A1( u0_u11_u1_n129 ) , .A2( u0_u11_u1_n133 ) , .ZN( u0_u11_u1_n149 ) );
  INV_X1 u0_u11_u1_U29 (.A( u0_u11_u1_n131 ) , .ZN( u0_u11_u1_n180 ) );
  INV_X1 u0_u11_u1_U3 (.A( u0_u11_u1_n159 ) , .ZN( u0_u11_u1_n182 ) );
  OAI221_X1 u0_u11_u1_U30 (.A( u0_u11_u1_n119 ) , .C2( u0_u11_u1_n129 ) , .ZN( u0_u11_u1_n138 ) , .B2( u0_u11_u1_n152 ) , .C1( u0_u11_u1_n174 ) , .B1( u0_u11_u1_n187 ) );
  INV_X1 u0_u11_u1_U31 (.A( u0_u11_u1_n148 ) , .ZN( u0_u11_u1_n187 ) );
  AOI211_X1 u0_u11_u1_U32 (.B( u0_u11_u1_n117 ) , .A( u0_u11_u1_n118 ) , .ZN( u0_u11_u1_n119 ) , .C2( u0_u11_u1_n146 ) , .C1( u0_u11_u1_n159 ) );
  NOR2_X1 u0_u11_u1_U33 (.A1( u0_u11_u1_n168 ) , .A2( u0_u11_u1_n176 ) , .ZN( u0_u11_u1_n98 ) );
  AOI211_X1 u0_u11_u1_U34 (.B( u0_u11_u1_n162 ) , .A( u0_u11_u1_n163 ) , .C2( u0_u11_u1_n164 ) , .ZN( u0_u11_u1_n165 ) , .C1( u0_u11_u1_n171 ) );
  AOI21_X1 u0_u11_u1_U35 (.A( u0_u11_u1_n160 ) , .B2( u0_u11_u1_n161 ) , .ZN( u0_u11_u1_n162 ) , .B1( u0_u11_u1_n182 ) );
  OR2_X1 u0_u11_u1_U36 (.A2( u0_u11_u1_n157 ) , .A1( u0_u11_u1_n158 ) , .ZN( u0_u11_u1_n163 ) );
  NAND2_X1 u0_u11_u1_U37 (.A1( u0_u11_u1_n128 ) , .ZN( u0_u11_u1_n146 ) , .A2( u0_u11_u1_n160 ) );
  NAND2_X1 u0_u11_u1_U38 (.A2( u0_u11_u1_n112 ) , .ZN( u0_u11_u1_n139 ) , .A1( u0_u11_u1_n152 ) );
  NAND2_X1 u0_u11_u1_U39 (.A1( u0_u11_u1_n105 ) , .ZN( u0_u11_u1_n156 ) , .A2( u0_u11_u1_n99 ) );
  AOI221_X1 u0_u11_u1_U4 (.A( u0_u11_u1_n138 ) , .C2( u0_u11_u1_n139 ) , .C1( u0_u11_u1_n140 ) , .B2( u0_u11_u1_n141 ) , .ZN( u0_u11_u1_n142 ) , .B1( u0_u11_u1_n175 ) );
  AOI221_X1 u0_u11_u1_U40 (.B1( u0_u11_u1_n140 ) , .ZN( u0_u11_u1_n167 ) , .B2( u0_u11_u1_n172 ) , .C2( u0_u11_u1_n175 ) , .C1( u0_u11_u1_n178 ) , .A( u0_u11_u1_n188 ) );
  INV_X1 u0_u11_u1_U41 (.ZN( u0_u11_u1_n188 ) , .A( u0_u11_u1_n97 ) );
  AOI211_X1 u0_u11_u1_U42 (.A( u0_u11_u1_n118 ) , .C1( u0_u11_u1_n132 ) , .C2( u0_u11_u1_n139 ) , .B( u0_u11_u1_n96 ) , .ZN( u0_u11_u1_n97 ) );
  AOI21_X1 u0_u11_u1_U43 (.B2( u0_u11_u1_n121 ) , .B1( u0_u11_u1_n135 ) , .A( u0_u11_u1_n152 ) , .ZN( u0_u11_u1_n96 ) );
  NOR2_X1 u0_u11_u1_U44 (.ZN( u0_u11_u1_n117 ) , .A1( u0_u11_u1_n121 ) , .A2( u0_u11_u1_n160 ) );
  OAI21_X1 u0_u11_u1_U45 (.B2( u0_u11_u1_n123 ) , .ZN( u0_u11_u1_n145 ) , .B1( u0_u11_u1_n160 ) , .A( u0_u11_u1_n185 ) );
  INV_X1 u0_u11_u1_U46 (.A( u0_u11_u1_n122 ) , .ZN( u0_u11_u1_n185 ) );
  AOI21_X1 u0_u11_u1_U47 (.B2( u0_u11_u1_n120 ) , .B1( u0_u11_u1_n121 ) , .ZN( u0_u11_u1_n122 ) , .A( u0_u11_u1_n128 ) );
  AOI21_X1 u0_u11_u1_U48 (.A( u0_u11_u1_n128 ) , .B2( u0_u11_u1_n129 ) , .ZN( u0_u11_u1_n130 ) , .B1( u0_u11_u1_n150 ) );
  NAND2_X1 u0_u11_u1_U49 (.ZN( u0_u11_u1_n112 ) , .A1( u0_u11_u1_n169 ) , .A2( u0_u11_u1_n170 ) );
  AOI211_X1 u0_u11_u1_U5 (.ZN( u0_u11_u1_n124 ) , .A( u0_u11_u1_n138 ) , .C2( u0_u11_u1_n139 ) , .B( u0_u11_u1_n145 ) , .C1( u0_u11_u1_n147 ) );
  NAND2_X1 u0_u11_u1_U50 (.ZN( u0_u11_u1_n129 ) , .A2( u0_u11_u1_n95 ) , .A1( u0_u11_u1_n98 ) );
  NAND2_X1 u0_u11_u1_U51 (.A1( u0_u11_u1_n102 ) , .ZN( u0_u11_u1_n154 ) , .A2( u0_u11_u1_n99 ) );
  NAND2_X1 u0_u11_u1_U52 (.A2( u0_u11_u1_n100 ) , .ZN( u0_u11_u1_n135 ) , .A1( u0_u11_u1_n99 ) );
  AOI21_X1 u0_u11_u1_U53 (.A( u0_u11_u1_n152 ) , .B2( u0_u11_u1_n153 ) , .B1( u0_u11_u1_n154 ) , .ZN( u0_u11_u1_n158 ) );
  INV_X1 u0_u11_u1_U54 (.A( u0_u11_u1_n160 ) , .ZN( u0_u11_u1_n175 ) );
  NAND2_X1 u0_u11_u1_U55 (.A1( u0_u11_u1_n100 ) , .ZN( u0_u11_u1_n116 ) , .A2( u0_u11_u1_n95 ) );
  NAND2_X1 u0_u11_u1_U56 (.A1( u0_u11_u1_n102 ) , .ZN( u0_u11_u1_n131 ) , .A2( u0_u11_u1_n95 ) );
  NAND2_X1 u0_u11_u1_U57 (.A2( u0_u11_u1_n104 ) , .ZN( u0_u11_u1_n121 ) , .A1( u0_u11_u1_n98 ) );
  NAND2_X1 u0_u11_u1_U58 (.A1( u0_u11_u1_n103 ) , .ZN( u0_u11_u1_n153 ) , .A2( u0_u11_u1_n98 ) );
  NAND2_X1 u0_u11_u1_U59 (.A2( u0_u11_u1_n104 ) , .A1( u0_u11_u1_n105 ) , .ZN( u0_u11_u1_n133 ) );
  AOI22_X1 u0_u11_u1_U6 (.B2( u0_u11_u1_n113 ) , .A2( u0_u11_u1_n114 ) , .ZN( u0_u11_u1_n125 ) , .A1( u0_u11_u1_n171 ) , .B1( u0_u11_u1_n173 ) );
  NAND2_X1 u0_u11_u1_U60 (.ZN( u0_u11_u1_n150 ) , .A2( u0_u11_u1_n98 ) , .A1( u0_u11_u1_n99 ) );
  NAND2_X1 u0_u11_u1_U61 (.A1( u0_u11_u1_n105 ) , .ZN( u0_u11_u1_n155 ) , .A2( u0_u11_u1_n95 ) );
  OAI21_X1 u0_u11_u1_U62 (.ZN( u0_u11_u1_n109 ) , .B1( u0_u11_u1_n129 ) , .B2( u0_u11_u1_n160 ) , .A( u0_u11_u1_n167 ) );
  NAND2_X1 u0_u11_u1_U63 (.A2( u0_u11_u1_n100 ) , .A1( u0_u11_u1_n103 ) , .ZN( u0_u11_u1_n120 ) );
  NAND2_X1 u0_u11_u1_U64 (.A1( u0_u11_u1_n102 ) , .A2( u0_u11_u1_n104 ) , .ZN( u0_u11_u1_n115 ) );
  NAND2_X1 u0_u11_u1_U65 (.A2( u0_u11_u1_n100 ) , .A1( u0_u11_u1_n104 ) , .ZN( u0_u11_u1_n151 ) );
  NAND2_X1 u0_u11_u1_U66 (.A2( u0_u11_u1_n103 ) , .A1( u0_u11_u1_n105 ) , .ZN( u0_u11_u1_n161 ) );
  INV_X1 u0_u11_u1_U67 (.A( u0_u11_u1_n152 ) , .ZN( u0_u11_u1_n173 ) );
  INV_X1 u0_u11_u1_U68 (.A( u0_u11_u1_n128 ) , .ZN( u0_u11_u1_n172 ) );
  NAND2_X1 u0_u11_u1_U69 (.A2( u0_u11_u1_n102 ) , .A1( u0_u11_u1_n103 ) , .ZN( u0_u11_u1_n123 ) );
  NAND2_X1 u0_u11_u1_U7 (.ZN( u0_u11_u1_n114 ) , .A1( u0_u11_u1_n134 ) , .A2( u0_u11_u1_n156 ) );
  NOR2_X1 u0_u11_u1_U70 (.A2( u0_u11_X_7 ) , .A1( u0_u11_X_8 ) , .ZN( u0_u11_u1_n95 ) );
  NOR2_X1 u0_u11_u1_U71 (.A1( u0_u11_X_12 ) , .A2( u0_u11_X_9 ) , .ZN( u0_u11_u1_n100 ) );
  NOR2_X1 u0_u11_u1_U72 (.A2( u0_u11_X_8 ) , .A1( u0_u11_u1_n177 ) , .ZN( u0_u11_u1_n99 ) );
  NOR2_X1 u0_u11_u1_U73 (.A2( u0_u11_X_12 ) , .ZN( u0_u11_u1_n102 ) , .A1( u0_u11_u1_n176 ) );
  NOR2_X1 u0_u11_u1_U74 (.A2( u0_u11_X_9 ) , .ZN( u0_u11_u1_n105 ) , .A1( u0_u11_u1_n168 ) );
  NAND2_X1 u0_u11_u1_U75 (.A1( u0_u11_X_10 ) , .ZN( u0_u11_u1_n160 ) , .A2( u0_u11_u1_n169 ) );
  NAND2_X1 u0_u11_u1_U76 (.A2( u0_u11_X_10 ) , .A1( u0_u11_X_11 ) , .ZN( u0_u11_u1_n152 ) );
  NAND2_X1 u0_u11_u1_U77 (.A1( u0_u11_X_11 ) , .ZN( u0_u11_u1_n128 ) , .A2( u0_u11_u1_n170 ) );
  AND2_X1 u0_u11_u1_U78 (.A2( u0_u11_X_7 ) , .A1( u0_u11_X_8 ) , .ZN( u0_u11_u1_n104 ) );
  AND2_X1 u0_u11_u1_U79 (.A1( u0_u11_X_8 ) , .ZN( u0_u11_u1_n103 ) , .A2( u0_u11_u1_n177 ) );
  AOI22_X1 u0_u11_u1_U8 (.B2( u0_u11_u1_n136 ) , .A2( u0_u11_u1_n137 ) , .ZN( u0_u11_u1_n143 ) , .A1( u0_u11_u1_n171 ) , .B1( u0_u11_u1_n173 ) );
  INV_X1 u0_u11_u1_U80 (.A( u0_u11_X_10 ) , .ZN( u0_u11_u1_n170 ) );
  INV_X1 u0_u11_u1_U81 (.A( u0_u11_X_9 ) , .ZN( u0_u11_u1_n176 ) );
  INV_X1 u0_u11_u1_U82 (.A( u0_u11_X_11 ) , .ZN( u0_u11_u1_n169 ) );
  INV_X1 u0_u11_u1_U83 (.A( u0_u11_X_12 ) , .ZN( u0_u11_u1_n168 ) );
  INV_X1 u0_u11_u1_U84 (.A( u0_u11_X_7 ) , .ZN( u0_u11_u1_n177 ) );
  NAND4_X1 u0_u11_u1_U85 (.ZN( u0_out11_28 ) , .A4( u0_u11_u1_n124 ) , .A3( u0_u11_u1_n125 ) , .A2( u0_u11_u1_n126 ) , .A1( u0_u11_u1_n127 ) );
  OAI21_X1 u0_u11_u1_U86 (.ZN( u0_u11_u1_n127 ) , .B2( u0_u11_u1_n139 ) , .B1( u0_u11_u1_n175 ) , .A( u0_u11_u1_n183 ) );
  OAI21_X1 u0_u11_u1_U87 (.ZN( u0_u11_u1_n126 ) , .B2( u0_u11_u1_n140 ) , .A( u0_u11_u1_n146 ) , .B1( u0_u11_u1_n178 ) );
  NAND4_X1 u0_u11_u1_U88 (.ZN( u0_out11_18 ) , .A4( u0_u11_u1_n165 ) , .A3( u0_u11_u1_n166 ) , .A1( u0_u11_u1_n167 ) , .A2( u0_u11_u1_n186 ) );
  AOI22_X1 u0_u11_u1_U89 (.B2( u0_u11_u1_n146 ) , .B1( u0_u11_u1_n147 ) , .A2( u0_u11_u1_n148 ) , .ZN( u0_u11_u1_n166 ) , .A1( u0_u11_u1_n172 ) );
  INV_X1 u0_u11_u1_U9 (.A( u0_u11_u1_n147 ) , .ZN( u0_u11_u1_n181 ) );
  INV_X1 u0_u11_u1_U90 (.A( u0_u11_u1_n145 ) , .ZN( u0_u11_u1_n186 ) );
  NAND4_X1 u0_u11_u1_U91 (.ZN( u0_out11_2 ) , .A4( u0_u11_u1_n142 ) , .A3( u0_u11_u1_n143 ) , .A2( u0_u11_u1_n144 ) , .A1( u0_u11_u1_n179 ) );
  OAI21_X1 u0_u11_u1_U92 (.B2( u0_u11_u1_n132 ) , .ZN( u0_u11_u1_n144 ) , .A( u0_u11_u1_n146 ) , .B1( u0_u11_u1_n180 ) );
  INV_X1 u0_u11_u1_U93 (.A( u0_u11_u1_n130 ) , .ZN( u0_u11_u1_n179 ) );
  OR4_X1 u0_u11_u1_U94 (.ZN( u0_out11_13 ) , .A4( u0_u11_u1_n108 ) , .A3( u0_u11_u1_n109 ) , .A2( u0_u11_u1_n110 ) , .A1( u0_u11_u1_n111 ) );
  AOI21_X1 u0_u11_u1_U95 (.ZN( u0_u11_u1_n111 ) , .A( u0_u11_u1_n128 ) , .B2( u0_u11_u1_n131 ) , .B1( u0_u11_u1_n135 ) );
  AOI21_X1 u0_u11_u1_U96 (.ZN( u0_u11_u1_n110 ) , .A( u0_u11_u1_n116 ) , .B1( u0_u11_u1_n152 ) , .B2( u0_u11_u1_n160 ) );
  NAND3_X1 u0_u11_u1_U97 (.A3( u0_u11_u1_n149 ) , .A2( u0_u11_u1_n150 ) , .A1( u0_u11_u1_n151 ) , .ZN( u0_u11_u1_n164 ) );
  NAND3_X1 u0_u11_u1_U98 (.A3( u0_u11_u1_n134 ) , .A2( u0_u11_u1_n135 ) , .ZN( u0_u11_u1_n136 ) , .A1( u0_u11_u1_n151 ) );
  NAND3_X1 u0_u11_u1_U99 (.A1( u0_u11_u1_n133 ) , .ZN( u0_u11_u1_n137 ) , .A2( u0_u11_u1_n154 ) , .A3( u0_u11_u1_n181 ) );
  OAI22_X1 u0_u11_u2_U10 (.ZN( u0_u11_u2_n109 ) , .A2( u0_u11_u2_n113 ) , .B2( u0_u11_u2_n133 ) , .B1( u0_u11_u2_n167 ) , .A1( u0_u11_u2_n168 ) );
  NAND3_X1 u0_u11_u2_U100 (.A2( u0_u11_u2_n100 ) , .A1( u0_u11_u2_n104 ) , .A3( u0_u11_u2_n138 ) , .ZN( u0_u11_u2_n98 ) );
  OAI22_X1 u0_u11_u2_U11 (.B1( u0_u11_u2_n151 ) , .A2( u0_u11_u2_n152 ) , .A1( u0_u11_u2_n153 ) , .ZN( u0_u11_u2_n160 ) , .B2( u0_u11_u2_n168 ) );
  NOR3_X1 u0_u11_u2_U12 (.A1( u0_u11_u2_n150 ) , .ZN( u0_u11_u2_n151 ) , .A3( u0_u11_u2_n175 ) , .A2( u0_u11_u2_n188 ) );
  AOI21_X1 u0_u11_u2_U13 (.ZN( u0_u11_u2_n144 ) , .B2( u0_u11_u2_n155 ) , .A( u0_u11_u2_n172 ) , .B1( u0_u11_u2_n185 ) );
  AOI21_X1 u0_u11_u2_U14 (.B2( u0_u11_u2_n143 ) , .ZN( u0_u11_u2_n145 ) , .B1( u0_u11_u2_n152 ) , .A( u0_u11_u2_n171 ) );
  AOI21_X1 u0_u11_u2_U15 (.B2( u0_u11_u2_n120 ) , .B1( u0_u11_u2_n121 ) , .ZN( u0_u11_u2_n126 ) , .A( u0_u11_u2_n167 ) );
  INV_X1 u0_u11_u2_U16 (.A( u0_u11_u2_n156 ) , .ZN( u0_u11_u2_n171 ) );
  INV_X1 u0_u11_u2_U17 (.A( u0_u11_u2_n120 ) , .ZN( u0_u11_u2_n188 ) );
  NAND2_X1 u0_u11_u2_U18 (.A2( u0_u11_u2_n122 ) , .ZN( u0_u11_u2_n150 ) , .A1( u0_u11_u2_n152 ) );
  INV_X1 u0_u11_u2_U19 (.A( u0_u11_u2_n153 ) , .ZN( u0_u11_u2_n170 ) );
  INV_X1 u0_u11_u2_U20 (.A( u0_u11_u2_n137 ) , .ZN( u0_u11_u2_n173 ) );
  NAND2_X1 u0_u11_u2_U21 (.A1( u0_u11_u2_n132 ) , .A2( u0_u11_u2_n139 ) , .ZN( u0_u11_u2_n157 ) );
  INV_X1 u0_u11_u2_U22 (.A( u0_u11_u2_n113 ) , .ZN( u0_u11_u2_n178 ) );
  INV_X1 u0_u11_u2_U23 (.A( u0_u11_u2_n139 ) , .ZN( u0_u11_u2_n175 ) );
  INV_X1 u0_u11_u2_U24 (.A( u0_u11_u2_n155 ) , .ZN( u0_u11_u2_n181 ) );
  INV_X1 u0_u11_u2_U25 (.A( u0_u11_u2_n119 ) , .ZN( u0_u11_u2_n177 ) );
  INV_X1 u0_u11_u2_U26 (.A( u0_u11_u2_n116 ) , .ZN( u0_u11_u2_n180 ) );
  INV_X1 u0_u11_u2_U27 (.A( u0_u11_u2_n131 ) , .ZN( u0_u11_u2_n179 ) );
  INV_X1 u0_u11_u2_U28 (.A( u0_u11_u2_n154 ) , .ZN( u0_u11_u2_n176 ) );
  NAND2_X1 u0_u11_u2_U29 (.A2( u0_u11_u2_n116 ) , .A1( u0_u11_u2_n117 ) , .ZN( u0_u11_u2_n118 ) );
  NOR2_X1 u0_u11_u2_U3 (.ZN( u0_u11_u2_n121 ) , .A2( u0_u11_u2_n177 ) , .A1( u0_u11_u2_n180 ) );
  INV_X1 u0_u11_u2_U30 (.A( u0_u11_u2_n132 ) , .ZN( u0_u11_u2_n182 ) );
  INV_X1 u0_u11_u2_U31 (.A( u0_u11_u2_n158 ) , .ZN( u0_u11_u2_n183 ) );
  OAI21_X1 u0_u11_u2_U32 (.A( u0_u11_u2_n156 ) , .B1( u0_u11_u2_n157 ) , .ZN( u0_u11_u2_n158 ) , .B2( u0_u11_u2_n179 ) );
  NOR2_X1 u0_u11_u2_U33 (.ZN( u0_u11_u2_n156 ) , .A1( u0_u11_u2_n166 ) , .A2( u0_u11_u2_n169 ) );
  NOR2_X1 u0_u11_u2_U34 (.A2( u0_u11_u2_n114 ) , .ZN( u0_u11_u2_n137 ) , .A1( u0_u11_u2_n140 ) );
  NOR2_X1 u0_u11_u2_U35 (.A2( u0_u11_u2_n138 ) , .ZN( u0_u11_u2_n153 ) , .A1( u0_u11_u2_n156 ) );
  AOI211_X1 u0_u11_u2_U36 (.ZN( u0_u11_u2_n130 ) , .C1( u0_u11_u2_n138 ) , .C2( u0_u11_u2_n179 ) , .B( u0_u11_u2_n96 ) , .A( u0_u11_u2_n97 ) );
  OAI22_X1 u0_u11_u2_U37 (.B1( u0_u11_u2_n133 ) , .A2( u0_u11_u2_n137 ) , .A1( u0_u11_u2_n152 ) , .B2( u0_u11_u2_n168 ) , .ZN( u0_u11_u2_n97 ) );
  OAI221_X1 u0_u11_u2_U38 (.B1( u0_u11_u2_n113 ) , .C1( u0_u11_u2_n132 ) , .A( u0_u11_u2_n149 ) , .B2( u0_u11_u2_n171 ) , .C2( u0_u11_u2_n172 ) , .ZN( u0_u11_u2_n96 ) );
  OAI221_X1 u0_u11_u2_U39 (.A( u0_u11_u2_n115 ) , .C2( u0_u11_u2_n123 ) , .B2( u0_u11_u2_n143 ) , .B1( u0_u11_u2_n153 ) , .ZN( u0_u11_u2_n163 ) , .C1( u0_u11_u2_n168 ) );
  INV_X1 u0_u11_u2_U4 (.A( u0_u11_u2_n134 ) , .ZN( u0_u11_u2_n185 ) );
  OAI21_X1 u0_u11_u2_U40 (.A( u0_u11_u2_n114 ) , .ZN( u0_u11_u2_n115 ) , .B1( u0_u11_u2_n176 ) , .B2( u0_u11_u2_n178 ) );
  OAI221_X1 u0_u11_u2_U41 (.A( u0_u11_u2_n135 ) , .B2( u0_u11_u2_n136 ) , .B1( u0_u11_u2_n137 ) , .ZN( u0_u11_u2_n162 ) , .C2( u0_u11_u2_n167 ) , .C1( u0_u11_u2_n185 ) );
  AND3_X1 u0_u11_u2_U42 (.A3( u0_u11_u2_n131 ) , .A2( u0_u11_u2_n132 ) , .A1( u0_u11_u2_n133 ) , .ZN( u0_u11_u2_n136 ) );
  AOI22_X1 u0_u11_u2_U43 (.ZN( u0_u11_u2_n135 ) , .B1( u0_u11_u2_n140 ) , .A1( u0_u11_u2_n156 ) , .B2( u0_u11_u2_n180 ) , .A2( u0_u11_u2_n188 ) );
  AOI21_X1 u0_u11_u2_U44 (.ZN( u0_u11_u2_n149 ) , .B1( u0_u11_u2_n173 ) , .B2( u0_u11_u2_n188 ) , .A( u0_u11_u2_n95 ) );
  AND3_X1 u0_u11_u2_U45 (.A2( u0_u11_u2_n100 ) , .A1( u0_u11_u2_n104 ) , .A3( u0_u11_u2_n156 ) , .ZN( u0_u11_u2_n95 ) );
  OAI21_X1 u0_u11_u2_U46 (.A( u0_u11_u2_n101 ) , .B2( u0_u11_u2_n121 ) , .B1( u0_u11_u2_n153 ) , .ZN( u0_u11_u2_n164 ) );
  NAND2_X1 u0_u11_u2_U47 (.A2( u0_u11_u2_n100 ) , .A1( u0_u11_u2_n107 ) , .ZN( u0_u11_u2_n155 ) );
  NAND2_X1 u0_u11_u2_U48 (.A2( u0_u11_u2_n105 ) , .A1( u0_u11_u2_n108 ) , .ZN( u0_u11_u2_n143 ) );
  NAND2_X1 u0_u11_u2_U49 (.A1( u0_u11_u2_n104 ) , .A2( u0_u11_u2_n106 ) , .ZN( u0_u11_u2_n152 ) );
  INV_X1 u0_u11_u2_U5 (.A( u0_u11_u2_n150 ) , .ZN( u0_u11_u2_n184 ) );
  NAND2_X1 u0_u11_u2_U50 (.A1( u0_u11_u2_n100 ) , .A2( u0_u11_u2_n105 ) , .ZN( u0_u11_u2_n132 ) );
  INV_X1 u0_u11_u2_U51 (.A( u0_u11_u2_n140 ) , .ZN( u0_u11_u2_n168 ) );
  INV_X1 u0_u11_u2_U52 (.A( u0_u11_u2_n138 ) , .ZN( u0_u11_u2_n167 ) );
  OAI21_X1 u0_u11_u2_U53 (.A( u0_u11_u2_n141 ) , .B2( u0_u11_u2_n142 ) , .ZN( u0_u11_u2_n146 ) , .B1( u0_u11_u2_n153 ) );
  OAI21_X1 u0_u11_u2_U54 (.A( u0_u11_u2_n140 ) , .ZN( u0_u11_u2_n141 ) , .B1( u0_u11_u2_n176 ) , .B2( u0_u11_u2_n177 ) );
  NOR3_X1 u0_u11_u2_U55 (.ZN( u0_u11_u2_n142 ) , .A3( u0_u11_u2_n175 ) , .A2( u0_u11_u2_n178 ) , .A1( u0_u11_u2_n181 ) );
  NAND2_X1 u0_u11_u2_U56 (.A1( u0_u11_u2_n102 ) , .A2( u0_u11_u2_n106 ) , .ZN( u0_u11_u2_n113 ) );
  NAND2_X1 u0_u11_u2_U57 (.A1( u0_u11_u2_n106 ) , .A2( u0_u11_u2_n107 ) , .ZN( u0_u11_u2_n131 ) );
  NAND2_X1 u0_u11_u2_U58 (.A1( u0_u11_u2_n103 ) , .A2( u0_u11_u2_n107 ) , .ZN( u0_u11_u2_n139 ) );
  NAND2_X1 u0_u11_u2_U59 (.A1( u0_u11_u2_n103 ) , .A2( u0_u11_u2_n105 ) , .ZN( u0_u11_u2_n133 ) );
  NOR4_X1 u0_u11_u2_U6 (.A4( u0_u11_u2_n124 ) , .A3( u0_u11_u2_n125 ) , .A2( u0_u11_u2_n126 ) , .A1( u0_u11_u2_n127 ) , .ZN( u0_u11_u2_n128 ) );
  NAND2_X1 u0_u11_u2_U60 (.A1( u0_u11_u2_n102 ) , .A2( u0_u11_u2_n103 ) , .ZN( u0_u11_u2_n154 ) );
  NAND2_X1 u0_u11_u2_U61 (.A2( u0_u11_u2_n103 ) , .A1( u0_u11_u2_n104 ) , .ZN( u0_u11_u2_n119 ) );
  NAND2_X1 u0_u11_u2_U62 (.A2( u0_u11_u2_n107 ) , .A1( u0_u11_u2_n108 ) , .ZN( u0_u11_u2_n123 ) );
  NAND2_X1 u0_u11_u2_U63 (.A1( u0_u11_u2_n104 ) , .A2( u0_u11_u2_n108 ) , .ZN( u0_u11_u2_n122 ) );
  INV_X1 u0_u11_u2_U64 (.A( u0_u11_u2_n114 ) , .ZN( u0_u11_u2_n172 ) );
  NAND2_X1 u0_u11_u2_U65 (.A2( u0_u11_u2_n100 ) , .A1( u0_u11_u2_n102 ) , .ZN( u0_u11_u2_n116 ) );
  NAND2_X1 u0_u11_u2_U66 (.A1( u0_u11_u2_n102 ) , .A2( u0_u11_u2_n108 ) , .ZN( u0_u11_u2_n120 ) );
  NAND2_X1 u0_u11_u2_U67 (.A2( u0_u11_u2_n105 ) , .A1( u0_u11_u2_n106 ) , .ZN( u0_u11_u2_n117 ) );
  INV_X1 u0_u11_u2_U68 (.ZN( u0_u11_u2_n187 ) , .A( u0_u11_u2_n99 ) );
  OAI21_X1 u0_u11_u2_U69 (.B1( u0_u11_u2_n137 ) , .B2( u0_u11_u2_n143 ) , .A( u0_u11_u2_n98 ) , .ZN( u0_u11_u2_n99 ) );
  AOI21_X1 u0_u11_u2_U7 (.ZN( u0_u11_u2_n124 ) , .B1( u0_u11_u2_n131 ) , .B2( u0_u11_u2_n143 ) , .A( u0_u11_u2_n172 ) );
  NOR2_X1 u0_u11_u2_U70 (.A2( u0_u11_X_16 ) , .ZN( u0_u11_u2_n140 ) , .A1( u0_u11_u2_n166 ) );
  NOR2_X1 u0_u11_u2_U71 (.A2( u0_u11_X_13 ) , .A1( u0_u11_X_14 ) , .ZN( u0_u11_u2_n100 ) );
  NOR2_X1 u0_u11_u2_U72 (.A2( u0_u11_X_16 ) , .A1( u0_u11_X_17 ) , .ZN( u0_u11_u2_n138 ) );
  NOR2_X1 u0_u11_u2_U73 (.A2( u0_u11_X_15 ) , .A1( u0_u11_X_18 ) , .ZN( u0_u11_u2_n104 ) );
  NOR2_X1 u0_u11_u2_U74 (.A2( u0_u11_X_14 ) , .ZN( u0_u11_u2_n103 ) , .A1( u0_u11_u2_n174 ) );
  NOR2_X1 u0_u11_u2_U75 (.A2( u0_u11_X_15 ) , .ZN( u0_u11_u2_n102 ) , .A1( u0_u11_u2_n165 ) );
  NOR2_X1 u0_u11_u2_U76 (.A2( u0_u11_X_17 ) , .ZN( u0_u11_u2_n114 ) , .A1( u0_u11_u2_n169 ) );
  AND2_X1 u0_u11_u2_U77 (.A1( u0_u11_X_15 ) , .ZN( u0_u11_u2_n105 ) , .A2( u0_u11_u2_n165 ) );
  AND2_X1 u0_u11_u2_U78 (.A2( u0_u11_X_15 ) , .A1( u0_u11_X_18 ) , .ZN( u0_u11_u2_n107 ) );
  AND2_X1 u0_u11_u2_U79 (.A1( u0_u11_X_14 ) , .ZN( u0_u11_u2_n106 ) , .A2( u0_u11_u2_n174 ) );
  AOI21_X1 u0_u11_u2_U8 (.B2( u0_u11_u2_n119 ) , .ZN( u0_u11_u2_n127 ) , .A( u0_u11_u2_n137 ) , .B1( u0_u11_u2_n155 ) );
  AND2_X1 u0_u11_u2_U80 (.A1( u0_u11_X_13 ) , .A2( u0_u11_X_14 ) , .ZN( u0_u11_u2_n108 ) );
  INV_X1 u0_u11_u2_U81 (.A( u0_u11_X_16 ) , .ZN( u0_u11_u2_n169 ) );
  INV_X1 u0_u11_u2_U82 (.A( u0_u11_X_17 ) , .ZN( u0_u11_u2_n166 ) );
  INV_X1 u0_u11_u2_U83 (.A( u0_u11_X_13 ) , .ZN( u0_u11_u2_n174 ) );
  INV_X1 u0_u11_u2_U84 (.A( u0_u11_X_18 ) , .ZN( u0_u11_u2_n165 ) );
  NAND4_X1 u0_u11_u2_U85 (.ZN( u0_out11_30 ) , .A4( u0_u11_u2_n147 ) , .A3( u0_u11_u2_n148 ) , .A2( u0_u11_u2_n149 ) , .A1( u0_u11_u2_n187 ) );
  NOR3_X1 u0_u11_u2_U86 (.A3( u0_u11_u2_n144 ) , .A2( u0_u11_u2_n145 ) , .A1( u0_u11_u2_n146 ) , .ZN( u0_u11_u2_n147 ) );
  AOI21_X1 u0_u11_u2_U87 (.B2( u0_u11_u2_n138 ) , .ZN( u0_u11_u2_n148 ) , .A( u0_u11_u2_n162 ) , .B1( u0_u11_u2_n182 ) );
  NAND4_X1 u0_u11_u2_U88 (.ZN( u0_out11_24 ) , .A4( u0_u11_u2_n111 ) , .A3( u0_u11_u2_n112 ) , .A1( u0_u11_u2_n130 ) , .A2( u0_u11_u2_n187 ) );
  AOI221_X1 u0_u11_u2_U89 (.A( u0_u11_u2_n109 ) , .B1( u0_u11_u2_n110 ) , .ZN( u0_u11_u2_n111 ) , .C1( u0_u11_u2_n134 ) , .C2( u0_u11_u2_n170 ) , .B2( u0_u11_u2_n173 ) );
  AOI21_X1 u0_u11_u2_U9 (.B2( u0_u11_u2_n123 ) , .ZN( u0_u11_u2_n125 ) , .A( u0_u11_u2_n171 ) , .B1( u0_u11_u2_n184 ) );
  AOI21_X1 u0_u11_u2_U90 (.ZN( u0_u11_u2_n112 ) , .B2( u0_u11_u2_n156 ) , .A( u0_u11_u2_n164 ) , .B1( u0_u11_u2_n181 ) );
  NAND4_X1 u0_u11_u2_U91 (.ZN( u0_out11_16 ) , .A4( u0_u11_u2_n128 ) , .A3( u0_u11_u2_n129 ) , .A1( u0_u11_u2_n130 ) , .A2( u0_u11_u2_n186 ) );
  AOI22_X1 u0_u11_u2_U92 (.A2( u0_u11_u2_n118 ) , .ZN( u0_u11_u2_n129 ) , .A1( u0_u11_u2_n140 ) , .B1( u0_u11_u2_n157 ) , .B2( u0_u11_u2_n170 ) );
  INV_X1 u0_u11_u2_U93 (.A( u0_u11_u2_n163 ) , .ZN( u0_u11_u2_n186 ) );
  OR4_X1 u0_u11_u2_U94 (.ZN( u0_out11_6 ) , .A4( u0_u11_u2_n161 ) , .A3( u0_u11_u2_n162 ) , .A2( u0_u11_u2_n163 ) , .A1( u0_u11_u2_n164 ) );
  OR3_X1 u0_u11_u2_U95 (.A2( u0_u11_u2_n159 ) , .A1( u0_u11_u2_n160 ) , .ZN( u0_u11_u2_n161 ) , .A3( u0_u11_u2_n183 ) );
  AOI21_X1 u0_u11_u2_U96 (.B2( u0_u11_u2_n154 ) , .B1( u0_u11_u2_n155 ) , .ZN( u0_u11_u2_n159 ) , .A( u0_u11_u2_n167 ) );
  NAND3_X1 u0_u11_u2_U97 (.A2( u0_u11_u2_n117 ) , .A1( u0_u11_u2_n122 ) , .A3( u0_u11_u2_n123 ) , .ZN( u0_u11_u2_n134 ) );
  NAND3_X1 u0_u11_u2_U98 (.ZN( u0_u11_u2_n110 ) , .A2( u0_u11_u2_n131 ) , .A3( u0_u11_u2_n139 ) , .A1( u0_u11_u2_n154 ) );
  NAND3_X1 u0_u11_u2_U99 (.A2( u0_u11_u2_n100 ) , .ZN( u0_u11_u2_n101 ) , .A1( u0_u11_u2_n104 ) , .A3( u0_u11_u2_n114 ) );
  OAI211_X1 u0_u11_u3_U10 (.B( u0_u11_u3_n106 ) , .ZN( u0_u11_u3_n119 ) , .C2( u0_u11_u3_n128 ) , .C1( u0_u11_u3_n167 ) , .A( u0_u11_u3_n181 ) );
  INV_X1 u0_u11_u3_U11 (.ZN( u0_u11_u3_n181 ) , .A( u0_u11_u3_n98 ) );
  AOI221_X1 u0_u11_u3_U12 (.C1( u0_u11_u3_n105 ) , .ZN( u0_u11_u3_n106 ) , .A( u0_u11_u3_n131 ) , .B2( u0_u11_u3_n132 ) , .C2( u0_u11_u3_n133 ) , .B1( u0_u11_u3_n169 ) );
  OAI22_X1 u0_u11_u3_U13 (.B1( u0_u11_u3_n113 ) , .A2( u0_u11_u3_n135 ) , .A1( u0_u11_u3_n150 ) , .B2( u0_u11_u3_n164 ) , .ZN( u0_u11_u3_n98 ) );
  AOI22_X1 u0_u11_u3_U14 (.B1( u0_u11_u3_n115 ) , .A2( u0_u11_u3_n116 ) , .ZN( u0_u11_u3_n123 ) , .B2( u0_u11_u3_n133 ) , .A1( u0_u11_u3_n169 ) );
  NAND2_X1 u0_u11_u3_U15 (.ZN( u0_u11_u3_n116 ) , .A2( u0_u11_u3_n151 ) , .A1( u0_u11_u3_n182 ) );
  NOR2_X1 u0_u11_u3_U16 (.ZN( u0_u11_u3_n126 ) , .A2( u0_u11_u3_n150 ) , .A1( u0_u11_u3_n164 ) );
  AOI21_X1 u0_u11_u3_U17 (.ZN( u0_u11_u3_n112 ) , .B2( u0_u11_u3_n146 ) , .B1( u0_u11_u3_n155 ) , .A( u0_u11_u3_n167 ) );
  NAND2_X1 u0_u11_u3_U18 (.A1( u0_u11_u3_n135 ) , .ZN( u0_u11_u3_n142 ) , .A2( u0_u11_u3_n164 ) );
  NAND2_X1 u0_u11_u3_U19 (.ZN( u0_u11_u3_n132 ) , .A2( u0_u11_u3_n152 ) , .A1( u0_u11_u3_n156 ) );
  INV_X1 u0_u11_u3_U20 (.A( u0_u11_u3_n133 ) , .ZN( u0_u11_u3_n165 ) );
  NAND2_X1 u0_u11_u3_U21 (.ZN( u0_u11_u3_n143 ) , .A1( u0_u11_u3_n165 ) , .A2( u0_u11_u3_n167 ) );
  AND2_X1 u0_u11_u3_U22 (.A2( u0_u11_u3_n113 ) , .A1( u0_u11_u3_n114 ) , .ZN( u0_u11_u3_n151 ) );
  INV_X1 u0_u11_u3_U23 (.A( u0_u11_u3_n135 ) , .ZN( u0_u11_u3_n170 ) );
  NAND2_X1 u0_u11_u3_U24 (.A1( u0_u11_u3_n107 ) , .A2( u0_u11_u3_n108 ) , .ZN( u0_u11_u3_n140 ) );
  NAND2_X1 u0_u11_u3_U25 (.ZN( u0_u11_u3_n117 ) , .A1( u0_u11_u3_n124 ) , .A2( u0_u11_u3_n148 ) );
  INV_X1 u0_u11_u3_U26 (.A( u0_u11_u3_n130 ) , .ZN( u0_u11_u3_n177 ) );
  INV_X1 u0_u11_u3_U27 (.A( u0_u11_u3_n128 ) , .ZN( u0_u11_u3_n176 ) );
  NAND2_X1 u0_u11_u3_U28 (.ZN( u0_u11_u3_n105 ) , .A2( u0_u11_u3_n130 ) , .A1( u0_u11_u3_n155 ) );
  INV_X1 u0_u11_u3_U29 (.A( u0_u11_u3_n155 ) , .ZN( u0_u11_u3_n174 ) );
  INV_X1 u0_u11_u3_U3 (.A( u0_u11_u3_n140 ) , .ZN( u0_u11_u3_n182 ) );
  INV_X1 u0_u11_u3_U30 (.A( u0_u11_u3_n139 ) , .ZN( u0_u11_u3_n185 ) );
  NOR2_X1 u0_u11_u3_U31 (.ZN( u0_u11_u3_n135 ) , .A2( u0_u11_u3_n141 ) , .A1( u0_u11_u3_n169 ) );
  INV_X1 u0_u11_u3_U32 (.A( u0_u11_u3_n156 ) , .ZN( u0_u11_u3_n179 ) );
  OAI22_X1 u0_u11_u3_U33 (.B1( u0_u11_u3_n118 ) , .ZN( u0_u11_u3_n120 ) , .A1( u0_u11_u3_n135 ) , .B2( u0_u11_u3_n154 ) , .A2( u0_u11_u3_n178 ) );
  AND3_X1 u0_u11_u3_U34 (.ZN( u0_u11_u3_n118 ) , .A2( u0_u11_u3_n124 ) , .A1( u0_u11_u3_n144 ) , .A3( u0_u11_u3_n152 ) );
  OAI222_X1 u0_u11_u3_U35 (.C2( u0_u11_u3_n107 ) , .A2( u0_u11_u3_n108 ) , .B1( u0_u11_u3_n135 ) , .ZN( u0_u11_u3_n138 ) , .B2( u0_u11_u3_n146 ) , .C1( u0_u11_u3_n154 ) , .A1( u0_u11_u3_n164 ) );
  NOR4_X1 u0_u11_u3_U36 (.A4( u0_u11_u3_n157 ) , .A3( u0_u11_u3_n158 ) , .A2( u0_u11_u3_n159 ) , .A1( u0_u11_u3_n160 ) , .ZN( u0_u11_u3_n161 ) );
  AOI21_X1 u0_u11_u3_U37 (.B2( u0_u11_u3_n152 ) , .B1( u0_u11_u3_n153 ) , .ZN( u0_u11_u3_n158 ) , .A( u0_u11_u3_n164 ) );
  AOI21_X1 u0_u11_u3_U38 (.A( u0_u11_u3_n154 ) , .B2( u0_u11_u3_n155 ) , .B1( u0_u11_u3_n156 ) , .ZN( u0_u11_u3_n157 ) );
  AOI21_X1 u0_u11_u3_U39 (.A( u0_u11_u3_n149 ) , .B2( u0_u11_u3_n150 ) , .B1( u0_u11_u3_n151 ) , .ZN( u0_u11_u3_n159 ) );
  INV_X1 u0_u11_u3_U4 (.A( u0_u11_u3_n129 ) , .ZN( u0_u11_u3_n183 ) );
  AOI211_X1 u0_u11_u3_U40 (.ZN( u0_u11_u3_n109 ) , .A( u0_u11_u3_n119 ) , .C2( u0_u11_u3_n129 ) , .B( u0_u11_u3_n138 ) , .C1( u0_u11_u3_n141 ) );
  INV_X1 u0_u11_u3_U41 (.A( u0_u11_u3_n121 ) , .ZN( u0_u11_u3_n164 ) );
  NAND2_X1 u0_u11_u3_U42 (.ZN( u0_u11_u3_n133 ) , .A1( u0_u11_u3_n154 ) , .A2( u0_u11_u3_n164 ) );
  OAI211_X1 u0_u11_u3_U43 (.B( u0_u11_u3_n127 ) , .ZN( u0_u11_u3_n139 ) , .C1( u0_u11_u3_n150 ) , .C2( u0_u11_u3_n154 ) , .A( u0_u11_u3_n184 ) );
  INV_X1 u0_u11_u3_U44 (.A( u0_u11_u3_n125 ) , .ZN( u0_u11_u3_n184 ) );
  AOI221_X1 u0_u11_u3_U45 (.A( u0_u11_u3_n126 ) , .ZN( u0_u11_u3_n127 ) , .C2( u0_u11_u3_n132 ) , .C1( u0_u11_u3_n169 ) , .B2( u0_u11_u3_n170 ) , .B1( u0_u11_u3_n174 ) );
  OAI22_X1 u0_u11_u3_U46 (.A1( u0_u11_u3_n124 ) , .ZN( u0_u11_u3_n125 ) , .B2( u0_u11_u3_n145 ) , .A2( u0_u11_u3_n165 ) , .B1( u0_u11_u3_n167 ) );
  NOR2_X1 u0_u11_u3_U47 (.A1( u0_u11_u3_n113 ) , .ZN( u0_u11_u3_n131 ) , .A2( u0_u11_u3_n154 ) );
  NAND2_X1 u0_u11_u3_U48 (.A1( u0_u11_u3_n103 ) , .ZN( u0_u11_u3_n150 ) , .A2( u0_u11_u3_n99 ) );
  NAND2_X1 u0_u11_u3_U49 (.A2( u0_u11_u3_n102 ) , .ZN( u0_u11_u3_n155 ) , .A1( u0_u11_u3_n97 ) );
  INV_X1 u0_u11_u3_U5 (.A( u0_u11_u3_n117 ) , .ZN( u0_u11_u3_n178 ) );
  INV_X1 u0_u11_u3_U50 (.A( u0_u11_u3_n141 ) , .ZN( u0_u11_u3_n167 ) );
  AOI21_X1 u0_u11_u3_U51 (.B2( u0_u11_u3_n114 ) , .B1( u0_u11_u3_n146 ) , .A( u0_u11_u3_n154 ) , .ZN( u0_u11_u3_n94 ) );
  AOI21_X1 u0_u11_u3_U52 (.ZN( u0_u11_u3_n110 ) , .B2( u0_u11_u3_n142 ) , .B1( u0_u11_u3_n186 ) , .A( u0_u11_u3_n95 ) );
  INV_X1 u0_u11_u3_U53 (.A( u0_u11_u3_n145 ) , .ZN( u0_u11_u3_n186 ) );
  AOI21_X1 u0_u11_u3_U54 (.B1( u0_u11_u3_n124 ) , .A( u0_u11_u3_n149 ) , .B2( u0_u11_u3_n155 ) , .ZN( u0_u11_u3_n95 ) );
  INV_X1 u0_u11_u3_U55 (.A( u0_u11_u3_n149 ) , .ZN( u0_u11_u3_n169 ) );
  NAND2_X1 u0_u11_u3_U56 (.ZN( u0_u11_u3_n124 ) , .A1( u0_u11_u3_n96 ) , .A2( u0_u11_u3_n97 ) );
  NAND2_X1 u0_u11_u3_U57 (.A2( u0_u11_u3_n100 ) , .ZN( u0_u11_u3_n146 ) , .A1( u0_u11_u3_n96 ) );
  NAND2_X1 u0_u11_u3_U58 (.A1( u0_u11_u3_n101 ) , .ZN( u0_u11_u3_n145 ) , .A2( u0_u11_u3_n99 ) );
  NAND2_X1 u0_u11_u3_U59 (.A1( u0_u11_u3_n100 ) , .ZN( u0_u11_u3_n156 ) , .A2( u0_u11_u3_n99 ) );
  AOI221_X1 u0_u11_u3_U6 (.A( u0_u11_u3_n131 ) , .C2( u0_u11_u3_n132 ) , .C1( u0_u11_u3_n133 ) , .ZN( u0_u11_u3_n134 ) , .B1( u0_u11_u3_n143 ) , .B2( u0_u11_u3_n177 ) );
  NAND2_X1 u0_u11_u3_U60 (.A2( u0_u11_u3_n101 ) , .A1( u0_u11_u3_n104 ) , .ZN( u0_u11_u3_n148 ) );
  NAND2_X1 u0_u11_u3_U61 (.A1( u0_u11_u3_n100 ) , .A2( u0_u11_u3_n102 ) , .ZN( u0_u11_u3_n128 ) );
  NAND2_X1 u0_u11_u3_U62 (.A2( u0_u11_u3_n101 ) , .A1( u0_u11_u3_n102 ) , .ZN( u0_u11_u3_n152 ) );
  NAND2_X1 u0_u11_u3_U63 (.A2( u0_u11_u3_n101 ) , .ZN( u0_u11_u3_n114 ) , .A1( u0_u11_u3_n96 ) );
  NAND2_X1 u0_u11_u3_U64 (.ZN( u0_u11_u3_n107 ) , .A1( u0_u11_u3_n97 ) , .A2( u0_u11_u3_n99 ) );
  NAND2_X1 u0_u11_u3_U65 (.A2( u0_u11_u3_n100 ) , .A1( u0_u11_u3_n104 ) , .ZN( u0_u11_u3_n113 ) );
  NAND2_X1 u0_u11_u3_U66 (.A1( u0_u11_u3_n104 ) , .ZN( u0_u11_u3_n153 ) , .A2( u0_u11_u3_n97 ) );
  NAND2_X1 u0_u11_u3_U67 (.A2( u0_u11_u3_n103 ) , .A1( u0_u11_u3_n104 ) , .ZN( u0_u11_u3_n130 ) );
  NAND2_X1 u0_u11_u3_U68 (.A2( u0_u11_u3_n103 ) , .ZN( u0_u11_u3_n144 ) , .A1( u0_u11_u3_n96 ) );
  NAND2_X1 u0_u11_u3_U69 (.A1( u0_u11_u3_n102 ) , .A2( u0_u11_u3_n103 ) , .ZN( u0_u11_u3_n108 ) );
  OAI22_X1 u0_u11_u3_U7 (.B2( u0_u11_u3_n147 ) , .A2( u0_u11_u3_n148 ) , .ZN( u0_u11_u3_n160 ) , .B1( u0_u11_u3_n165 ) , .A1( u0_u11_u3_n168 ) );
  NOR2_X1 u0_u11_u3_U70 (.A2( u0_u11_X_19 ) , .A1( u0_u11_X_20 ) , .ZN( u0_u11_u3_n99 ) );
  NOR2_X1 u0_u11_u3_U71 (.A2( u0_u11_X_21 ) , .A1( u0_u11_X_24 ) , .ZN( u0_u11_u3_n103 ) );
  NOR2_X1 u0_u11_u3_U72 (.A2( u0_u11_X_24 ) , .A1( u0_u11_u3_n171 ) , .ZN( u0_u11_u3_n97 ) );
  NOR2_X1 u0_u11_u3_U73 (.A2( u0_u11_X_19 ) , .A1( u0_u11_u3_n172 ) , .ZN( u0_u11_u3_n96 ) );
  NAND2_X1 u0_u11_u3_U74 (.A1( u0_u11_X_22 ) , .A2( u0_u11_X_23 ) , .ZN( u0_u11_u3_n154 ) );
  AND2_X1 u0_u11_u3_U75 (.A1( u0_u11_X_24 ) , .ZN( u0_u11_u3_n101 ) , .A2( u0_u11_u3_n171 ) );
  AND2_X1 u0_u11_u3_U76 (.A1( u0_u11_X_19 ) , .ZN( u0_u11_u3_n102 ) , .A2( u0_u11_u3_n172 ) );
  AND2_X1 u0_u11_u3_U77 (.A1( u0_u11_X_21 ) , .A2( u0_u11_X_24 ) , .ZN( u0_u11_u3_n100 ) );
  AND2_X1 u0_u11_u3_U78 (.A2( u0_u11_X_19 ) , .A1( u0_u11_X_20 ) , .ZN( u0_u11_u3_n104 ) );
  INV_X1 u0_u11_u3_U79 (.A( u0_u11_X_21 ) , .ZN( u0_u11_u3_n171 ) );
  AND3_X1 u0_u11_u3_U8 (.A3( u0_u11_u3_n144 ) , .A2( u0_u11_u3_n145 ) , .A1( u0_u11_u3_n146 ) , .ZN( u0_u11_u3_n147 ) );
  INV_X1 u0_u11_u3_U80 (.A( u0_u11_X_20 ) , .ZN( u0_u11_u3_n172 ) );
  INV_X1 u0_u11_u3_U81 (.A( u0_u11_X_22 ) , .ZN( u0_u11_u3_n166 ) );
  NAND4_X1 u0_u11_u3_U82 (.ZN( u0_out11_26 ) , .A4( u0_u11_u3_n109 ) , .A3( u0_u11_u3_n110 ) , .A2( u0_u11_u3_n111 ) , .A1( u0_u11_u3_n173 ) );
  INV_X1 u0_u11_u3_U83 (.ZN( u0_u11_u3_n173 ) , .A( u0_u11_u3_n94 ) );
  OAI21_X1 u0_u11_u3_U84 (.ZN( u0_u11_u3_n111 ) , .B2( u0_u11_u3_n117 ) , .A( u0_u11_u3_n133 ) , .B1( u0_u11_u3_n176 ) );
  NAND4_X1 u0_u11_u3_U85 (.ZN( u0_out11_1 ) , .A4( u0_u11_u3_n161 ) , .A3( u0_u11_u3_n162 ) , .A2( u0_u11_u3_n163 ) , .A1( u0_u11_u3_n185 ) );
  NAND2_X1 u0_u11_u3_U86 (.ZN( u0_u11_u3_n163 ) , .A2( u0_u11_u3_n170 ) , .A1( u0_u11_u3_n176 ) );
  AOI22_X1 u0_u11_u3_U87 (.B2( u0_u11_u3_n140 ) , .B1( u0_u11_u3_n141 ) , .A2( u0_u11_u3_n142 ) , .ZN( u0_u11_u3_n162 ) , .A1( u0_u11_u3_n177 ) );
  NAND4_X1 u0_u11_u3_U88 (.ZN( u0_out11_20 ) , .A4( u0_u11_u3_n122 ) , .A3( u0_u11_u3_n123 ) , .A1( u0_u11_u3_n175 ) , .A2( u0_u11_u3_n180 ) );
  INV_X1 u0_u11_u3_U89 (.A( u0_u11_u3_n126 ) , .ZN( u0_u11_u3_n180 ) );
  INV_X1 u0_u11_u3_U9 (.A( u0_u11_u3_n143 ) , .ZN( u0_u11_u3_n168 ) );
  INV_X1 u0_u11_u3_U90 (.A( u0_u11_u3_n112 ) , .ZN( u0_u11_u3_n175 ) );
  OR4_X1 u0_u11_u3_U91 (.ZN( u0_out11_10 ) , .A4( u0_u11_u3_n136 ) , .A3( u0_u11_u3_n137 ) , .A1( u0_u11_u3_n138 ) , .A2( u0_u11_u3_n139 ) );
  OAI222_X1 u0_u11_u3_U92 (.C1( u0_u11_u3_n128 ) , .ZN( u0_u11_u3_n137 ) , .B1( u0_u11_u3_n148 ) , .A2( u0_u11_u3_n150 ) , .B2( u0_u11_u3_n154 ) , .C2( u0_u11_u3_n164 ) , .A1( u0_u11_u3_n167 ) );
  AOI211_X1 u0_u11_u3_U93 (.B( u0_u11_u3_n119 ) , .A( u0_u11_u3_n120 ) , .C2( u0_u11_u3_n121 ) , .ZN( u0_u11_u3_n122 ) , .C1( u0_u11_u3_n179 ) );
  OAI221_X1 u0_u11_u3_U94 (.A( u0_u11_u3_n134 ) , .B2( u0_u11_u3_n135 ) , .ZN( u0_u11_u3_n136 ) , .C1( u0_u11_u3_n149 ) , .B1( u0_u11_u3_n151 ) , .C2( u0_u11_u3_n183 ) );
  NOR2_X1 u0_u11_u3_U95 (.A2( u0_u11_X_23 ) , .ZN( u0_u11_u3_n141 ) , .A1( u0_u11_u3_n166 ) );
  NAND2_X1 u0_u11_u3_U96 (.A1( u0_u11_X_23 ) , .ZN( u0_u11_u3_n149 ) , .A2( u0_u11_u3_n166 ) );
  NOR2_X1 u0_u11_u3_U97 (.A2( u0_u11_X_22 ) , .A1( u0_u11_X_23 ) , .ZN( u0_u11_u3_n121 ) );
  NAND3_X1 u0_u11_u3_U98 (.A1( u0_u11_u3_n114 ) , .ZN( u0_u11_u3_n115 ) , .A2( u0_u11_u3_n145 ) , .A3( u0_u11_u3_n153 ) );
  NAND3_X1 u0_u11_u3_U99 (.ZN( u0_u11_u3_n129 ) , .A2( u0_u11_u3_n144 ) , .A1( u0_u11_u3_n153 ) , .A3( u0_u11_u3_n182 ) );
  XOR2_X1 u0_u15_U10 (.A( u0_FP_62 ) , .B( u0_K16_45 ) , .Z( u0_u15_X_45 ) );
  XOR2_X1 u0_u15_U11 (.A( u0_FP_61 ) , .B( u0_K16_44 ) , .Z( u0_u15_X_44 ) );
  XOR2_X1 u0_u15_U12 (.A( u0_FP_60 ) , .B( u0_K16_43 ) , .Z( u0_u15_X_43 ) );
  XOR2_X1 u0_u15_U33 (.A( u0_FP_49 ) , .B( u0_K16_24 ) , .Z( u0_u15_X_24 ) );
  XOR2_X1 u0_u15_U34 (.A( u0_FP_48 ) , .B( u0_K16_23 ) , .Z( u0_u15_X_23 ) );
  XOR2_X1 u0_u15_U35 (.A( u0_FP_47 ) , .B( u0_K16_22 ) , .Z( u0_u15_X_22 ) );
  XOR2_X1 u0_u15_U36 (.A( u0_FP_46 ) , .B( u0_K16_21 ) , .Z( u0_u15_X_21 ) );
  XOR2_X1 u0_u15_U37 (.A( u0_FP_45 ) , .B( u0_K16_20 ) , .Z( u0_u15_X_20 ) );
  XOR2_X1 u0_u15_U39 (.A( u0_FP_44 ) , .B( u0_K16_19 ) , .Z( u0_u15_X_19 ) );
  XOR2_X1 u0_u15_U40 (.A( u0_FP_45 ) , .B( u0_K16_18 ) , .Z( u0_u15_X_18 ) );
  XOR2_X1 u0_u15_U41 (.A( u0_FP_44 ) , .B( u0_K16_17 ) , .Z( u0_u15_X_17 ) );
  XOR2_X1 u0_u15_U42 (.A( u0_FP_43 ) , .B( u0_K16_16 ) , .Z( u0_u15_X_16 ) );
  XOR2_X1 u0_u15_U43 (.A( u0_FP_42 ) , .B( u0_K16_15 ) , .Z( u0_u15_X_15 ) );
  XOR2_X1 u0_u15_U44 (.A( u0_FP_41 ) , .B( u0_K16_14 ) , .Z( u0_u15_X_14 ) );
  XOR2_X1 u0_u15_U45 (.A( u0_FP_40 ) , .B( u0_K16_13 ) , .Z( u0_u15_X_13 ) );
  XOR2_X1 u0_u15_U7 (.A( u0_FP_33 ) , .B( u0_K16_48 ) , .Z( u0_u15_X_48 ) );
  XOR2_X1 u0_u15_U8 (.A( u0_FP_64 ) , .B( u0_K16_47 ) , .Z( u0_u15_X_47 ) );
  XOR2_X1 u0_u15_U9 (.A( u0_FP_63 ) , .B( u0_K16_46 ) , .Z( u0_u15_X_46 ) );
  OAI22_X1 u0_u15_u2_U10 (.B1( u0_u15_u2_n151 ) , .A2( u0_u15_u2_n152 ) , .A1( u0_u15_u2_n153 ) , .ZN( u0_u15_u2_n160 ) , .B2( u0_u15_u2_n168 ) );
  NAND3_X1 u0_u15_u2_U100 (.A2( u0_u15_u2_n100 ) , .A1( u0_u15_u2_n104 ) , .A3( u0_u15_u2_n138 ) , .ZN( u0_u15_u2_n98 ) );
  NOR3_X1 u0_u15_u2_U11 (.A1( u0_u15_u2_n150 ) , .ZN( u0_u15_u2_n151 ) , .A3( u0_u15_u2_n175 ) , .A2( u0_u15_u2_n188 ) );
  AOI21_X1 u0_u15_u2_U12 (.B2( u0_u15_u2_n123 ) , .ZN( u0_u15_u2_n125 ) , .A( u0_u15_u2_n171 ) , .B1( u0_u15_u2_n184 ) );
  INV_X1 u0_u15_u2_U13 (.A( u0_u15_u2_n150 ) , .ZN( u0_u15_u2_n184 ) );
  AOI21_X1 u0_u15_u2_U14 (.ZN( u0_u15_u2_n144 ) , .B2( u0_u15_u2_n155 ) , .A( u0_u15_u2_n172 ) , .B1( u0_u15_u2_n185 ) );
  AOI21_X1 u0_u15_u2_U15 (.B2( u0_u15_u2_n143 ) , .ZN( u0_u15_u2_n145 ) , .B1( u0_u15_u2_n152 ) , .A( u0_u15_u2_n171 ) );
  INV_X1 u0_u15_u2_U16 (.A( u0_u15_u2_n156 ) , .ZN( u0_u15_u2_n171 ) );
  INV_X1 u0_u15_u2_U17 (.A( u0_u15_u2_n120 ) , .ZN( u0_u15_u2_n188 ) );
  NAND2_X1 u0_u15_u2_U18 (.A2( u0_u15_u2_n122 ) , .ZN( u0_u15_u2_n150 ) , .A1( u0_u15_u2_n152 ) );
  INV_X1 u0_u15_u2_U19 (.A( u0_u15_u2_n153 ) , .ZN( u0_u15_u2_n170 ) );
  INV_X1 u0_u15_u2_U20 (.A( u0_u15_u2_n137 ) , .ZN( u0_u15_u2_n173 ) );
  NAND2_X1 u0_u15_u2_U21 (.A1( u0_u15_u2_n132 ) , .A2( u0_u15_u2_n139 ) , .ZN( u0_u15_u2_n157 ) );
  INV_X1 u0_u15_u2_U22 (.A( u0_u15_u2_n113 ) , .ZN( u0_u15_u2_n178 ) );
  INV_X1 u0_u15_u2_U23 (.A( u0_u15_u2_n139 ) , .ZN( u0_u15_u2_n175 ) );
  INV_X1 u0_u15_u2_U24 (.A( u0_u15_u2_n155 ) , .ZN( u0_u15_u2_n181 ) );
  INV_X1 u0_u15_u2_U25 (.A( u0_u15_u2_n119 ) , .ZN( u0_u15_u2_n177 ) );
  INV_X1 u0_u15_u2_U26 (.A( u0_u15_u2_n116 ) , .ZN( u0_u15_u2_n180 ) );
  INV_X1 u0_u15_u2_U27 (.A( u0_u15_u2_n131 ) , .ZN( u0_u15_u2_n179 ) );
  INV_X1 u0_u15_u2_U28 (.A( u0_u15_u2_n154 ) , .ZN( u0_u15_u2_n176 ) );
  NAND2_X1 u0_u15_u2_U29 (.A2( u0_u15_u2_n116 ) , .A1( u0_u15_u2_n117 ) , .ZN( u0_u15_u2_n118 ) );
  NOR2_X1 u0_u15_u2_U3 (.ZN( u0_u15_u2_n121 ) , .A2( u0_u15_u2_n177 ) , .A1( u0_u15_u2_n180 ) );
  INV_X1 u0_u15_u2_U30 (.A( u0_u15_u2_n132 ) , .ZN( u0_u15_u2_n182 ) );
  INV_X1 u0_u15_u2_U31 (.A( u0_u15_u2_n158 ) , .ZN( u0_u15_u2_n183 ) );
  OAI21_X1 u0_u15_u2_U32 (.A( u0_u15_u2_n156 ) , .B1( u0_u15_u2_n157 ) , .ZN( u0_u15_u2_n158 ) , .B2( u0_u15_u2_n179 ) );
  NOR2_X1 u0_u15_u2_U33 (.ZN( u0_u15_u2_n156 ) , .A1( u0_u15_u2_n166 ) , .A2( u0_u15_u2_n169 ) );
  NOR2_X1 u0_u15_u2_U34 (.A2( u0_u15_u2_n114 ) , .ZN( u0_u15_u2_n137 ) , .A1( u0_u15_u2_n140 ) );
  NOR2_X1 u0_u15_u2_U35 (.A2( u0_u15_u2_n138 ) , .ZN( u0_u15_u2_n153 ) , .A1( u0_u15_u2_n156 ) );
  AOI211_X1 u0_u15_u2_U36 (.ZN( u0_u15_u2_n130 ) , .C1( u0_u15_u2_n138 ) , .C2( u0_u15_u2_n179 ) , .B( u0_u15_u2_n96 ) , .A( u0_u15_u2_n97 ) );
  OAI22_X1 u0_u15_u2_U37 (.B1( u0_u15_u2_n133 ) , .A2( u0_u15_u2_n137 ) , .A1( u0_u15_u2_n152 ) , .B2( u0_u15_u2_n168 ) , .ZN( u0_u15_u2_n97 ) );
  OAI221_X1 u0_u15_u2_U38 (.B1( u0_u15_u2_n113 ) , .C1( u0_u15_u2_n132 ) , .A( u0_u15_u2_n149 ) , .B2( u0_u15_u2_n171 ) , .C2( u0_u15_u2_n172 ) , .ZN( u0_u15_u2_n96 ) );
  OAI221_X1 u0_u15_u2_U39 (.A( u0_u15_u2_n115 ) , .C2( u0_u15_u2_n123 ) , .B2( u0_u15_u2_n143 ) , .B1( u0_u15_u2_n153 ) , .ZN( u0_u15_u2_n163 ) , .C1( u0_u15_u2_n168 ) );
  INV_X1 u0_u15_u2_U4 (.A( u0_u15_u2_n134 ) , .ZN( u0_u15_u2_n185 ) );
  OAI21_X1 u0_u15_u2_U40 (.A( u0_u15_u2_n114 ) , .ZN( u0_u15_u2_n115 ) , .B1( u0_u15_u2_n176 ) , .B2( u0_u15_u2_n178 ) );
  OAI221_X1 u0_u15_u2_U41 (.A( u0_u15_u2_n135 ) , .B2( u0_u15_u2_n136 ) , .B1( u0_u15_u2_n137 ) , .ZN( u0_u15_u2_n162 ) , .C2( u0_u15_u2_n167 ) , .C1( u0_u15_u2_n185 ) );
  AND3_X1 u0_u15_u2_U42 (.A3( u0_u15_u2_n131 ) , .A2( u0_u15_u2_n132 ) , .A1( u0_u15_u2_n133 ) , .ZN( u0_u15_u2_n136 ) );
  AOI22_X1 u0_u15_u2_U43 (.ZN( u0_u15_u2_n135 ) , .B1( u0_u15_u2_n140 ) , .A1( u0_u15_u2_n156 ) , .B2( u0_u15_u2_n180 ) , .A2( u0_u15_u2_n188 ) );
  AOI21_X1 u0_u15_u2_U44 (.ZN( u0_u15_u2_n149 ) , .B1( u0_u15_u2_n173 ) , .B2( u0_u15_u2_n188 ) , .A( u0_u15_u2_n95 ) );
  AND3_X1 u0_u15_u2_U45 (.A2( u0_u15_u2_n100 ) , .A1( u0_u15_u2_n104 ) , .A3( u0_u15_u2_n156 ) , .ZN( u0_u15_u2_n95 ) );
  OAI21_X1 u0_u15_u2_U46 (.A( u0_u15_u2_n141 ) , .B2( u0_u15_u2_n142 ) , .ZN( u0_u15_u2_n146 ) , .B1( u0_u15_u2_n153 ) );
  OAI21_X1 u0_u15_u2_U47 (.A( u0_u15_u2_n140 ) , .ZN( u0_u15_u2_n141 ) , .B1( u0_u15_u2_n176 ) , .B2( u0_u15_u2_n177 ) );
  NOR3_X1 u0_u15_u2_U48 (.ZN( u0_u15_u2_n142 ) , .A3( u0_u15_u2_n175 ) , .A2( u0_u15_u2_n178 ) , .A1( u0_u15_u2_n181 ) );
  OAI21_X1 u0_u15_u2_U49 (.A( u0_u15_u2_n101 ) , .B2( u0_u15_u2_n121 ) , .B1( u0_u15_u2_n153 ) , .ZN( u0_u15_u2_n164 ) );
  NOR4_X1 u0_u15_u2_U5 (.A4( u0_u15_u2_n124 ) , .A3( u0_u15_u2_n125 ) , .A2( u0_u15_u2_n126 ) , .A1( u0_u15_u2_n127 ) , .ZN( u0_u15_u2_n128 ) );
  NAND2_X1 u0_u15_u2_U50 (.A2( u0_u15_u2_n100 ) , .A1( u0_u15_u2_n107 ) , .ZN( u0_u15_u2_n155 ) );
  NAND2_X1 u0_u15_u2_U51 (.A2( u0_u15_u2_n105 ) , .A1( u0_u15_u2_n108 ) , .ZN( u0_u15_u2_n143 ) );
  NAND2_X1 u0_u15_u2_U52 (.A1( u0_u15_u2_n104 ) , .A2( u0_u15_u2_n106 ) , .ZN( u0_u15_u2_n152 ) );
  NAND2_X1 u0_u15_u2_U53 (.A1( u0_u15_u2_n100 ) , .A2( u0_u15_u2_n105 ) , .ZN( u0_u15_u2_n132 ) );
  INV_X1 u0_u15_u2_U54 (.A( u0_u15_u2_n140 ) , .ZN( u0_u15_u2_n168 ) );
  INV_X1 u0_u15_u2_U55 (.A( u0_u15_u2_n138 ) , .ZN( u0_u15_u2_n167 ) );
  INV_X1 u0_u15_u2_U56 (.ZN( u0_u15_u2_n187 ) , .A( u0_u15_u2_n99 ) );
  OAI21_X1 u0_u15_u2_U57 (.B1( u0_u15_u2_n137 ) , .B2( u0_u15_u2_n143 ) , .A( u0_u15_u2_n98 ) , .ZN( u0_u15_u2_n99 ) );
  NAND2_X1 u0_u15_u2_U58 (.A1( u0_u15_u2_n102 ) , .A2( u0_u15_u2_n106 ) , .ZN( u0_u15_u2_n113 ) );
  NAND2_X1 u0_u15_u2_U59 (.A1( u0_u15_u2_n106 ) , .A2( u0_u15_u2_n107 ) , .ZN( u0_u15_u2_n131 ) );
  AOI21_X1 u0_u15_u2_U6 (.B2( u0_u15_u2_n119 ) , .ZN( u0_u15_u2_n127 ) , .A( u0_u15_u2_n137 ) , .B1( u0_u15_u2_n155 ) );
  NAND2_X1 u0_u15_u2_U60 (.A1( u0_u15_u2_n103 ) , .A2( u0_u15_u2_n107 ) , .ZN( u0_u15_u2_n139 ) );
  NAND2_X1 u0_u15_u2_U61 (.A1( u0_u15_u2_n103 ) , .A2( u0_u15_u2_n105 ) , .ZN( u0_u15_u2_n133 ) );
  NAND2_X1 u0_u15_u2_U62 (.A1( u0_u15_u2_n102 ) , .A2( u0_u15_u2_n103 ) , .ZN( u0_u15_u2_n154 ) );
  NAND2_X1 u0_u15_u2_U63 (.A2( u0_u15_u2_n103 ) , .A1( u0_u15_u2_n104 ) , .ZN( u0_u15_u2_n119 ) );
  NAND2_X1 u0_u15_u2_U64 (.A2( u0_u15_u2_n107 ) , .A1( u0_u15_u2_n108 ) , .ZN( u0_u15_u2_n123 ) );
  NAND2_X1 u0_u15_u2_U65 (.A1( u0_u15_u2_n104 ) , .A2( u0_u15_u2_n108 ) , .ZN( u0_u15_u2_n122 ) );
  INV_X1 u0_u15_u2_U66 (.A( u0_u15_u2_n114 ) , .ZN( u0_u15_u2_n172 ) );
  NAND2_X1 u0_u15_u2_U67 (.A2( u0_u15_u2_n100 ) , .A1( u0_u15_u2_n102 ) , .ZN( u0_u15_u2_n116 ) );
  NAND2_X1 u0_u15_u2_U68 (.A1( u0_u15_u2_n102 ) , .A2( u0_u15_u2_n108 ) , .ZN( u0_u15_u2_n120 ) );
  NAND2_X1 u0_u15_u2_U69 (.A2( u0_u15_u2_n105 ) , .A1( u0_u15_u2_n106 ) , .ZN( u0_u15_u2_n117 ) );
  AOI21_X1 u0_u15_u2_U7 (.ZN( u0_u15_u2_n124 ) , .B1( u0_u15_u2_n131 ) , .B2( u0_u15_u2_n143 ) , .A( u0_u15_u2_n172 ) );
  NOR2_X1 u0_u15_u2_U70 (.A2( u0_u15_X_16 ) , .ZN( u0_u15_u2_n140 ) , .A1( u0_u15_u2_n166 ) );
  NOR2_X1 u0_u15_u2_U71 (.A2( u0_u15_X_13 ) , .A1( u0_u15_X_14 ) , .ZN( u0_u15_u2_n100 ) );
  NOR2_X1 u0_u15_u2_U72 (.A2( u0_u15_X_16 ) , .A1( u0_u15_X_17 ) , .ZN( u0_u15_u2_n138 ) );
  NOR2_X1 u0_u15_u2_U73 (.A2( u0_u15_X_15 ) , .A1( u0_u15_X_18 ) , .ZN( u0_u15_u2_n104 ) );
  NOR2_X1 u0_u15_u2_U74 (.A2( u0_u15_X_14 ) , .ZN( u0_u15_u2_n103 ) , .A1( u0_u15_u2_n174 ) );
  NOR2_X1 u0_u15_u2_U75 (.A2( u0_u15_X_15 ) , .ZN( u0_u15_u2_n102 ) , .A1( u0_u15_u2_n165 ) );
  NOR2_X1 u0_u15_u2_U76 (.A2( u0_u15_X_17 ) , .ZN( u0_u15_u2_n114 ) , .A1( u0_u15_u2_n169 ) );
  AND2_X1 u0_u15_u2_U77 (.A1( u0_u15_X_15 ) , .ZN( u0_u15_u2_n105 ) , .A2( u0_u15_u2_n165 ) );
  AND2_X1 u0_u15_u2_U78 (.A2( u0_u15_X_15 ) , .A1( u0_u15_X_18 ) , .ZN( u0_u15_u2_n107 ) );
  AND2_X1 u0_u15_u2_U79 (.A1( u0_u15_X_14 ) , .ZN( u0_u15_u2_n106 ) , .A2( u0_u15_u2_n174 ) );
  AOI21_X1 u0_u15_u2_U8 (.B2( u0_u15_u2_n120 ) , .B1( u0_u15_u2_n121 ) , .ZN( u0_u15_u2_n126 ) , .A( u0_u15_u2_n167 ) );
  AND2_X1 u0_u15_u2_U80 (.A1( u0_u15_X_13 ) , .A2( u0_u15_X_14 ) , .ZN( u0_u15_u2_n108 ) );
  INV_X1 u0_u15_u2_U81 (.A( u0_u15_X_16 ) , .ZN( u0_u15_u2_n169 ) );
  INV_X1 u0_u15_u2_U82 (.A( u0_u15_X_17 ) , .ZN( u0_u15_u2_n166 ) );
  INV_X1 u0_u15_u2_U83 (.A( u0_u15_X_13 ) , .ZN( u0_u15_u2_n174 ) );
  INV_X1 u0_u15_u2_U84 (.A( u0_u15_X_18 ) , .ZN( u0_u15_u2_n165 ) );
  NAND4_X1 u0_u15_u2_U85 (.ZN( u0_out15_30 ) , .A4( u0_u15_u2_n147 ) , .A3( u0_u15_u2_n148 ) , .A2( u0_u15_u2_n149 ) , .A1( u0_u15_u2_n187 ) );
  NOR3_X1 u0_u15_u2_U86 (.A3( u0_u15_u2_n144 ) , .A2( u0_u15_u2_n145 ) , .A1( u0_u15_u2_n146 ) , .ZN( u0_u15_u2_n147 ) );
  AOI21_X1 u0_u15_u2_U87 (.B2( u0_u15_u2_n138 ) , .ZN( u0_u15_u2_n148 ) , .A( u0_u15_u2_n162 ) , .B1( u0_u15_u2_n182 ) );
  NAND4_X1 u0_u15_u2_U88 (.ZN( u0_out15_24 ) , .A4( u0_u15_u2_n111 ) , .A3( u0_u15_u2_n112 ) , .A1( u0_u15_u2_n130 ) , .A2( u0_u15_u2_n187 ) );
  AOI221_X1 u0_u15_u2_U89 (.A( u0_u15_u2_n109 ) , .B1( u0_u15_u2_n110 ) , .ZN( u0_u15_u2_n111 ) , .C1( u0_u15_u2_n134 ) , .C2( u0_u15_u2_n170 ) , .B2( u0_u15_u2_n173 ) );
  OAI22_X1 u0_u15_u2_U9 (.ZN( u0_u15_u2_n109 ) , .A2( u0_u15_u2_n113 ) , .B2( u0_u15_u2_n133 ) , .B1( u0_u15_u2_n167 ) , .A1( u0_u15_u2_n168 ) );
  AOI21_X1 u0_u15_u2_U90 (.ZN( u0_u15_u2_n112 ) , .B2( u0_u15_u2_n156 ) , .A( u0_u15_u2_n164 ) , .B1( u0_u15_u2_n181 ) );
  NAND4_X1 u0_u15_u2_U91 (.ZN( u0_out15_16 ) , .A4( u0_u15_u2_n128 ) , .A3( u0_u15_u2_n129 ) , .A1( u0_u15_u2_n130 ) , .A2( u0_u15_u2_n186 ) );
  AOI22_X1 u0_u15_u2_U92 (.A2( u0_u15_u2_n118 ) , .ZN( u0_u15_u2_n129 ) , .A1( u0_u15_u2_n140 ) , .B1( u0_u15_u2_n157 ) , .B2( u0_u15_u2_n170 ) );
  INV_X1 u0_u15_u2_U93 (.A( u0_u15_u2_n163 ) , .ZN( u0_u15_u2_n186 ) );
  OR4_X1 u0_u15_u2_U94 (.ZN( u0_out15_6 ) , .A4( u0_u15_u2_n161 ) , .A3( u0_u15_u2_n162 ) , .A2( u0_u15_u2_n163 ) , .A1( u0_u15_u2_n164 ) );
  OR3_X1 u0_u15_u2_U95 (.A2( u0_u15_u2_n159 ) , .A1( u0_u15_u2_n160 ) , .ZN( u0_u15_u2_n161 ) , .A3( u0_u15_u2_n183 ) );
  AOI21_X1 u0_u15_u2_U96 (.B2( u0_u15_u2_n154 ) , .B1( u0_u15_u2_n155 ) , .ZN( u0_u15_u2_n159 ) , .A( u0_u15_u2_n167 ) );
  NAND3_X1 u0_u15_u2_U97 (.A2( u0_u15_u2_n117 ) , .A1( u0_u15_u2_n122 ) , .A3( u0_u15_u2_n123 ) , .ZN( u0_u15_u2_n134 ) );
  NAND3_X1 u0_u15_u2_U98 (.ZN( u0_u15_u2_n110 ) , .A2( u0_u15_u2_n131 ) , .A3( u0_u15_u2_n139 ) , .A1( u0_u15_u2_n154 ) );
  NAND3_X1 u0_u15_u2_U99 (.A2( u0_u15_u2_n100 ) , .ZN( u0_u15_u2_n101 ) , .A1( u0_u15_u2_n104 ) , .A3( u0_u15_u2_n114 ) );
  OAI22_X1 u0_u15_u3_U10 (.B1( u0_u15_u3_n113 ) , .A2( u0_u15_u3_n135 ) , .A1( u0_u15_u3_n150 ) , .B2( u0_u15_u3_n164 ) , .ZN( u0_u15_u3_n98 ) );
  OAI211_X1 u0_u15_u3_U11 (.B( u0_u15_u3_n106 ) , .ZN( u0_u15_u3_n119 ) , .C2( u0_u15_u3_n128 ) , .C1( u0_u15_u3_n167 ) , .A( u0_u15_u3_n181 ) );
  AOI221_X1 u0_u15_u3_U12 (.C1( u0_u15_u3_n105 ) , .ZN( u0_u15_u3_n106 ) , .A( u0_u15_u3_n131 ) , .B2( u0_u15_u3_n132 ) , .C2( u0_u15_u3_n133 ) , .B1( u0_u15_u3_n169 ) );
  INV_X1 u0_u15_u3_U13 (.ZN( u0_u15_u3_n181 ) , .A( u0_u15_u3_n98 ) );
  NAND2_X1 u0_u15_u3_U14 (.ZN( u0_u15_u3_n105 ) , .A2( u0_u15_u3_n130 ) , .A1( u0_u15_u3_n155 ) );
  AOI22_X1 u0_u15_u3_U15 (.B1( u0_u15_u3_n115 ) , .A2( u0_u15_u3_n116 ) , .ZN( u0_u15_u3_n123 ) , .B2( u0_u15_u3_n133 ) , .A1( u0_u15_u3_n169 ) );
  NAND2_X1 u0_u15_u3_U16 (.ZN( u0_u15_u3_n116 ) , .A2( u0_u15_u3_n151 ) , .A1( u0_u15_u3_n182 ) );
  NOR2_X1 u0_u15_u3_U17 (.ZN( u0_u15_u3_n126 ) , .A2( u0_u15_u3_n150 ) , .A1( u0_u15_u3_n164 ) );
  AOI21_X1 u0_u15_u3_U18 (.ZN( u0_u15_u3_n112 ) , .B2( u0_u15_u3_n146 ) , .B1( u0_u15_u3_n155 ) , .A( u0_u15_u3_n167 ) );
  NAND2_X1 u0_u15_u3_U19 (.A1( u0_u15_u3_n135 ) , .ZN( u0_u15_u3_n142 ) , .A2( u0_u15_u3_n164 ) );
  NAND2_X1 u0_u15_u3_U20 (.ZN( u0_u15_u3_n132 ) , .A2( u0_u15_u3_n152 ) , .A1( u0_u15_u3_n156 ) );
  AND2_X1 u0_u15_u3_U21 (.A2( u0_u15_u3_n113 ) , .A1( u0_u15_u3_n114 ) , .ZN( u0_u15_u3_n151 ) );
  INV_X1 u0_u15_u3_U22 (.A( u0_u15_u3_n133 ) , .ZN( u0_u15_u3_n165 ) );
  INV_X1 u0_u15_u3_U23 (.A( u0_u15_u3_n135 ) , .ZN( u0_u15_u3_n170 ) );
  NAND2_X1 u0_u15_u3_U24 (.A1( u0_u15_u3_n107 ) , .A2( u0_u15_u3_n108 ) , .ZN( u0_u15_u3_n140 ) );
  NAND2_X1 u0_u15_u3_U25 (.ZN( u0_u15_u3_n117 ) , .A1( u0_u15_u3_n124 ) , .A2( u0_u15_u3_n148 ) );
  NAND2_X1 u0_u15_u3_U26 (.ZN( u0_u15_u3_n143 ) , .A1( u0_u15_u3_n165 ) , .A2( u0_u15_u3_n167 ) );
  INV_X1 u0_u15_u3_U27 (.A( u0_u15_u3_n130 ) , .ZN( u0_u15_u3_n177 ) );
  INV_X1 u0_u15_u3_U28 (.A( u0_u15_u3_n128 ) , .ZN( u0_u15_u3_n176 ) );
  INV_X1 u0_u15_u3_U29 (.A( u0_u15_u3_n155 ) , .ZN( u0_u15_u3_n174 ) );
  INV_X1 u0_u15_u3_U3 (.A( u0_u15_u3_n129 ) , .ZN( u0_u15_u3_n183 ) );
  INV_X1 u0_u15_u3_U30 (.A( u0_u15_u3_n139 ) , .ZN( u0_u15_u3_n185 ) );
  NOR2_X1 u0_u15_u3_U31 (.ZN( u0_u15_u3_n135 ) , .A2( u0_u15_u3_n141 ) , .A1( u0_u15_u3_n169 ) );
  OAI222_X1 u0_u15_u3_U32 (.C2( u0_u15_u3_n107 ) , .A2( u0_u15_u3_n108 ) , .B1( u0_u15_u3_n135 ) , .ZN( u0_u15_u3_n138 ) , .B2( u0_u15_u3_n146 ) , .C1( u0_u15_u3_n154 ) , .A1( u0_u15_u3_n164 ) );
  NOR4_X1 u0_u15_u3_U33 (.A4( u0_u15_u3_n157 ) , .A3( u0_u15_u3_n158 ) , .A2( u0_u15_u3_n159 ) , .A1( u0_u15_u3_n160 ) , .ZN( u0_u15_u3_n161 ) );
  AOI21_X1 u0_u15_u3_U34 (.B2( u0_u15_u3_n152 ) , .B1( u0_u15_u3_n153 ) , .ZN( u0_u15_u3_n158 ) , .A( u0_u15_u3_n164 ) );
  AOI21_X1 u0_u15_u3_U35 (.A( u0_u15_u3_n154 ) , .B2( u0_u15_u3_n155 ) , .B1( u0_u15_u3_n156 ) , .ZN( u0_u15_u3_n157 ) );
  AOI21_X1 u0_u15_u3_U36 (.A( u0_u15_u3_n149 ) , .B2( u0_u15_u3_n150 ) , .B1( u0_u15_u3_n151 ) , .ZN( u0_u15_u3_n159 ) );
  AOI211_X1 u0_u15_u3_U37 (.ZN( u0_u15_u3_n109 ) , .A( u0_u15_u3_n119 ) , .C2( u0_u15_u3_n129 ) , .B( u0_u15_u3_n138 ) , .C1( u0_u15_u3_n141 ) );
  AOI211_X1 u0_u15_u3_U38 (.B( u0_u15_u3_n119 ) , .A( u0_u15_u3_n120 ) , .C2( u0_u15_u3_n121 ) , .ZN( u0_u15_u3_n122 ) , .C1( u0_u15_u3_n179 ) );
  INV_X1 u0_u15_u3_U39 (.A( u0_u15_u3_n156 ) , .ZN( u0_u15_u3_n179 ) );
  INV_X1 u0_u15_u3_U4 (.A( u0_u15_u3_n140 ) , .ZN( u0_u15_u3_n182 ) );
  OAI22_X1 u0_u15_u3_U40 (.B1( u0_u15_u3_n118 ) , .ZN( u0_u15_u3_n120 ) , .A1( u0_u15_u3_n135 ) , .B2( u0_u15_u3_n154 ) , .A2( u0_u15_u3_n178 ) );
  AND3_X1 u0_u15_u3_U41 (.ZN( u0_u15_u3_n118 ) , .A2( u0_u15_u3_n124 ) , .A1( u0_u15_u3_n144 ) , .A3( u0_u15_u3_n152 ) );
  INV_X1 u0_u15_u3_U42 (.A( u0_u15_u3_n121 ) , .ZN( u0_u15_u3_n164 ) );
  NAND2_X1 u0_u15_u3_U43 (.ZN( u0_u15_u3_n133 ) , .A1( u0_u15_u3_n154 ) , .A2( u0_u15_u3_n164 ) );
  OAI211_X1 u0_u15_u3_U44 (.B( u0_u15_u3_n127 ) , .ZN( u0_u15_u3_n139 ) , .C1( u0_u15_u3_n150 ) , .C2( u0_u15_u3_n154 ) , .A( u0_u15_u3_n184 ) );
  INV_X1 u0_u15_u3_U45 (.A( u0_u15_u3_n125 ) , .ZN( u0_u15_u3_n184 ) );
  AOI221_X1 u0_u15_u3_U46 (.A( u0_u15_u3_n126 ) , .ZN( u0_u15_u3_n127 ) , .C2( u0_u15_u3_n132 ) , .C1( u0_u15_u3_n169 ) , .B2( u0_u15_u3_n170 ) , .B1( u0_u15_u3_n174 ) );
  OAI22_X1 u0_u15_u3_U47 (.A1( u0_u15_u3_n124 ) , .ZN( u0_u15_u3_n125 ) , .B2( u0_u15_u3_n145 ) , .A2( u0_u15_u3_n165 ) , .B1( u0_u15_u3_n167 ) );
  NOR2_X1 u0_u15_u3_U48 (.A1( u0_u15_u3_n113 ) , .ZN( u0_u15_u3_n131 ) , .A2( u0_u15_u3_n154 ) );
  NAND2_X1 u0_u15_u3_U49 (.A1( u0_u15_u3_n103 ) , .ZN( u0_u15_u3_n150 ) , .A2( u0_u15_u3_n99 ) );
  INV_X1 u0_u15_u3_U5 (.A( u0_u15_u3_n117 ) , .ZN( u0_u15_u3_n178 ) );
  NAND2_X1 u0_u15_u3_U50 (.A2( u0_u15_u3_n102 ) , .ZN( u0_u15_u3_n155 ) , .A1( u0_u15_u3_n97 ) );
  INV_X1 u0_u15_u3_U51 (.A( u0_u15_u3_n141 ) , .ZN( u0_u15_u3_n167 ) );
  AOI21_X1 u0_u15_u3_U52 (.B2( u0_u15_u3_n114 ) , .B1( u0_u15_u3_n146 ) , .A( u0_u15_u3_n154 ) , .ZN( u0_u15_u3_n94 ) );
  AOI21_X1 u0_u15_u3_U53 (.ZN( u0_u15_u3_n110 ) , .B2( u0_u15_u3_n142 ) , .B1( u0_u15_u3_n186 ) , .A( u0_u15_u3_n95 ) );
  INV_X1 u0_u15_u3_U54 (.A( u0_u15_u3_n145 ) , .ZN( u0_u15_u3_n186 ) );
  AOI21_X1 u0_u15_u3_U55 (.B1( u0_u15_u3_n124 ) , .A( u0_u15_u3_n149 ) , .B2( u0_u15_u3_n155 ) , .ZN( u0_u15_u3_n95 ) );
  INV_X1 u0_u15_u3_U56 (.A( u0_u15_u3_n149 ) , .ZN( u0_u15_u3_n169 ) );
  NAND2_X1 u0_u15_u3_U57 (.ZN( u0_u15_u3_n124 ) , .A1( u0_u15_u3_n96 ) , .A2( u0_u15_u3_n97 ) );
  NAND2_X1 u0_u15_u3_U58 (.A2( u0_u15_u3_n100 ) , .ZN( u0_u15_u3_n146 ) , .A1( u0_u15_u3_n96 ) );
  NAND2_X1 u0_u15_u3_U59 (.A1( u0_u15_u3_n101 ) , .ZN( u0_u15_u3_n145 ) , .A2( u0_u15_u3_n99 ) );
  AOI221_X1 u0_u15_u3_U6 (.A( u0_u15_u3_n131 ) , .C2( u0_u15_u3_n132 ) , .C1( u0_u15_u3_n133 ) , .ZN( u0_u15_u3_n134 ) , .B1( u0_u15_u3_n143 ) , .B2( u0_u15_u3_n177 ) );
  NAND2_X1 u0_u15_u3_U60 (.A1( u0_u15_u3_n100 ) , .ZN( u0_u15_u3_n156 ) , .A2( u0_u15_u3_n99 ) );
  NAND2_X1 u0_u15_u3_U61 (.A2( u0_u15_u3_n101 ) , .A1( u0_u15_u3_n104 ) , .ZN( u0_u15_u3_n148 ) );
  NAND2_X1 u0_u15_u3_U62 (.A1( u0_u15_u3_n100 ) , .A2( u0_u15_u3_n102 ) , .ZN( u0_u15_u3_n128 ) );
  NAND2_X1 u0_u15_u3_U63 (.A2( u0_u15_u3_n101 ) , .A1( u0_u15_u3_n102 ) , .ZN( u0_u15_u3_n152 ) );
  NAND2_X1 u0_u15_u3_U64 (.A2( u0_u15_u3_n101 ) , .ZN( u0_u15_u3_n114 ) , .A1( u0_u15_u3_n96 ) );
  NAND2_X1 u0_u15_u3_U65 (.ZN( u0_u15_u3_n107 ) , .A1( u0_u15_u3_n97 ) , .A2( u0_u15_u3_n99 ) );
  NAND2_X1 u0_u15_u3_U66 (.A2( u0_u15_u3_n100 ) , .A1( u0_u15_u3_n104 ) , .ZN( u0_u15_u3_n113 ) );
  NAND2_X1 u0_u15_u3_U67 (.A1( u0_u15_u3_n104 ) , .ZN( u0_u15_u3_n153 ) , .A2( u0_u15_u3_n97 ) );
  NAND2_X1 u0_u15_u3_U68 (.A2( u0_u15_u3_n103 ) , .A1( u0_u15_u3_n104 ) , .ZN( u0_u15_u3_n130 ) );
  NAND2_X1 u0_u15_u3_U69 (.A2( u0_u15_u3_n103 ) , .ZN( u0_u15_u3_n144 ) , .A1( u0_u15_u3_n96 ) );
  OAI22_X1 u0_u15_u3_U7 (.B2( u0_u15_u3_n147 ) , .A2( u0_u15_u3_n148 ) , .ZN( u0_u15_u3_n160 ) , .B1( u0_u15_u3_n165 ) , .A1( u0_u15_u3_n168 ) );
  NAND2_X1 u0_u15_u3_U70 (.A1( u0_u15_u3_n102 ) , .A2( u0_u15_u3_n103 ) , .ZN( u0_u15_u3_n108 ) );
  NOR2_X1 u0_u15_u3_U71 (.A2( u0_u15_X_19 ) , .A1( u0_u15_X_20 ) , .ZN( u0_u15_u3_n99 ) );
  NOR2_X1 u0_u15_u3_U72 (.A2( u0_u15_X_21 ) , .A1( u0_u15_X_24 ) , .ZN( u0_u15_u3_n103 ) );
  NOR2_X1 u0_u15_u3_U73 (.A2( u0_u15_X_24 ) , .A1( u0_u15_u3_n171 ) , .ZN( u0_u15_u3_n97 ) );
  NOR2_X1 u0_u15_u3_U74 (.A2( u0_u15_X_23 ) , .ZN( u0_u15_u3_n141 ) , .A1( u0_u15_u3_n166 ) );
  NOR2_X1 u0_u15_u3_U75 (.A2( u0_u15_X_19 ) , .A1( u0_u15_u3_n172 ) , .ZN( u0_u15_u3_n96 ) );
  NAND2_X1 u0_u15_u3_U76 (.A1( u0_u15_X_22 ) , .A2( u0_u15_X_23 ) , .ZN( u0_u15_u3_n154 ) );
  NAND2_X1 u0_u15_u3_U77 (.A1( u0_u15_X_23 ) , .ZN( u0_u15_u3_n149 ) , .A2( u0_u15_u3_n166 ) );
  NOR2_X1 u0_u15_u3_U78 (.A2( u0_u15_X_22 ) , .A1( u0_u15_X_23 ) , .ZN( u0_u15_u3_n121 ) );
  AND2_X1 u0_u15_u3_U79 (.A1( u0_u15_X_24 ) , .ZN( u0_u15_u3_n101 ) , .A2( u0_u15_u3_n171 ) );
  AND3_X1 u0_u15_u3_U8 (.A3( u0_u15_u3_n144 ) , .A2( u0_u15_u3_n145 ) , .A1( u0_u15_u3_n146 ) , .ZN( u0_u15_u3_n147 ) );
  AND2_X1 u0_u15_u3_U80 (.A1( u0_u15_X_19 ) , .ZN( u0_u15_u3_n102 ) , .A2( u0_u15_u3_n172 ) );
  AND2_X1 u0_u15_u3_U81 (.A1( u0_u15_X_21 ) , .A2( u0_u15_X_24 ) , .ZN( u0_u15_u3_n100 ) );
  AND2_X1 u0_u15_u3_U82 (.A2( u0_u15_X_19 ) , .A1( u0_u15_X_20 ) , .ZN( u0_u15_u3_n104 ) );
  INV_X1 u0_u15_u3_U83 (.A( u0_u15_X_22 ) , .ZN( u0_u15_u3_n166 ) );
  INV_X1 u0_u15_u3_U84 (.A( u0_u15_X_21 ) , .ZN( u0_u15_u3_n171 ) );
  INV_X1 u0_u15_u3_U85 (.A( u0_u15_X_20 ) , .ZN( u0_u15_u3_n172 ) );
  OR4_X1 u0_u15_u3_U86 (.ZN( u0_out15_10 ) , .A4( u0_u15_u3_n136 ) , .A3( u0_u15_u3_n137 ) , .A1( u0_u15_u3_n138 ) , .A2( u0_u15_u3_n139 ) );
  OAI222_X1 u0_u15_u3_U87 (.C1( u0_u15_u3_n128 ) , .ZN( u0_u15_u3_n137 ) , .B1( u0_u15_u3_n148 ) , .A2( u0_u15_u3_n150 ) , .B2( u0_u15_u3_n154 ) , .C2( u0_u15_u3_n164 ) , .A1( u0_u15_u3_n167 ) );
  OAI221_X1 u0_u15_u3_U88 (.A( u0_u15_u3_n134 ) , .B2( u0_u15_u3_n135 ) , .ZN( u0_u15_u3_n136 ) , .C1( u0_u15_u3_n149 ) , .B1( u0_u15_u3_n151 ) , .C2( u0_u15_u3_n183 ) );
  NAND4_X1 u0_u15_u3_U89 (.ZN( u0_out15_26 ) , .A4( u0_u15_u3_n109 ) , .A3( u0_u15_u3_n110 ) , .A2( u0_u15_u3_n111 ) , .A1( u0_u15_u3_n173 ) );
  INV_X1 u0_u15_u3_U9 (.A( u0_u15_u3_n143 ) , .ZN( u0_u15_u3_n168 ) );
  INV_X1 u0_u15_u3_U90 (.ZN( u0_u15_u3_n173 ) , .A( u0_u15_u3_n94 ) );
  OAI21_X1 u0_u15_u3_U91 (.ZN( u0_u15_u3_n111 ) , .B2( u0_u15_u3_n117 ) , .A( u0_u15_u3_n133 ) , .B1( u0_u15_u3_n176 ) );
  NAND4_X1 u0_u15_u3_U92 (.ZN( u0_out15_20 ) , .A4( u0_u15_u3_n122 ) , .A3( u0_u15_u3_n123 ) , .A1( u0_u15_u3_n175 ) , .A2( u0_u15_u3_n180 ) );
  INV_X1 u0_u15_u3_U93 (.A( u0_u15_u3_n126 ) , .ZN( u0_u15_u3_n180 ) );
  INV_X1 u0_u15_u3_U94 (.A( u0_u15_u3_n112 ) , .ZN( u0_u15_u3_n175 ) );
  NAND4_X1 u0_u15_u3_U95 (.ZN( u0_out15_1 ) , .A4( u0_u15_u3_n161 ) , .A3( u0_u15_u3_n162 ) , .A2( u0_u15_u3_n163 ) , .A1( u0_u15_u3_n185 ) );
  NAND2_X1 u0_u15_u3_U96 (.ZN( u0_u15_u3_n163 ) , .A2( u0_u15_u3_n170 ) , .A1( u0_u15_u3_n176 ) );
  AOI22_X1 u0_u15_u3_U97 (.B2( u0_u15_u3_n140 ) , .B1( u0_u15_u3_n141 ) , .A2( u0_u15_u3_n142 ) , .ZN( u0_u15_u3_n162 ) , .A1( u0_u15_u3_n177 ) );
  NAND3_X1 u0_u15_u3_U98 (.A1( u0_u15_u3_n114 ) , .ZN( u0_u15_u3_n115 ) , .A2( u0_u15_u3_n145 ) , .A3( u0_u15_u3_n153 ) );
  NAND3_X1 u0_u15_u3_U99 (.ZN( u0_u15_u3_n129 ) , .A2( u0_u15_u3_n144 ) , .A1( u0_u15_u3_n153 ) , .A3( u0_u15_u3_n182 ) );
  OAI21_X1 u0_u15_u7_U10 (.A( u0_u15_u7_n161 ) , .B1( u0_u15_u7_n168 ) , .B2( u0_u15_u7_n173 ) , .ZN( u0_u15_u7_n91 ) );
  AOI211_X1 u0_u15_u7_U11 (.A( u0_u15_u7_n117 ) , .ZN( u0_u15_u7_n118 ) , .C2( u0_u15_u7_n126 ) , .C1( u0_u15_u7_n177 ) , .B( u0_u15_u7_n180 ) );
  OAI22_X1 u0_u15_u7_U12 (.B1( u0_u15_u7_n115 ) , .ZN( u0_u15_u7_n117 ) , .A2( u0_u15_u7_n133 ) , .A1( u0_u15_u7_n137 ) , .B2( u0_u15_u7_n162 ) );
  INV_X1 u0_u15_u7_U13 (.A( u0_u15_u7_n116 ) , .ZN( u0_u15_u7_n180 ) );
  NOR3_X1 u0_u15_u7_U14 (.ZN( u0_u15_u7_n115 ) , .A3( u0_u15_u7_n145 ) , .A2( u0_u15_u7_n168 ) , .A1( u0_u15_u7_n169 ) );
  OAI211_X1 u0_u15_u7_U15 (.B( u0_u15_u7_n122 ) , .A( u0_u15_u7_n123 ) , .C2( u0_u15_u7_n124 ) , .ZN( u0_u15_u7_n154 ) , .C1( u0_u15_u7_n162 ) );
  AOI222_X1 u0_u15_u7_U16 (.ZN( u0_u15_u7_n122 ) , .C2( u0_u15_u7_n126 ) , .C1( u0_u15_u7_n145 ) , .B1( u0_u15_u7_n161 ) , .A2( u0_u15_u7_n165 ) , .B2( u0_u15_u7_n170 ) , .A1( u0_u15_u7_n176 ) );
  INV_X1 u0_u15_u7_U17 (.A( u0_u15_u7_n133 ) , .ZN( u0_u15_u7_n176 ) );
  NOR3_X1 u0_u15_u7_U18 (.A2( u0_u15_u7_n134 ) , .A1( u0_u15_u7_n135 ) , .ZN( u0_u15_u7_n136 ) , .A3( u0_u15_u7_n171 ) );
  NOR2_X1 u0_u15_u7_U19 (.A1( u0_u15_u7_n130 ) , .A2( u0_u15_u7_n134 ) , .ZN( u0_u15_u7_n153 ) );
  INV_X1 u0_u15_u7_U20 (.A( u0_u15_u7_n101 ) , .ZN( u0_u15_u7_n165 ) );
  NOR2_X1 u0_u15_u7_U21 (.ZN( u0_u15_u7_n111 ) , .A2( u0_u15_u7_n134 ) , .A1( u0_u15_u7_n169 ) );
  AOI21_X1 u0_u15_u7_U22 (.ZN( u0_u15_u7_n104 ) , .B2( u0_u15_u7_n112 ) , .B1( u0_u15_u7_n127 ) , .A( u0_u15_u7_n164 ) );
  AOI21_X1 u0_u15_u7_U23 (.ZN( u0_u15_u7_n106 ) , .B1( u0_u15_u7_n133 ) , .B2( u0_u15_u7_n146 ) , .A( u0_u15_u7_n162 ) );
  AOI21_X1 u0_u15_u7_U24 (.A( u0_u15_u7_n101 ) , .ZN( u0_u15_u7_n107 ) , .B2( u0_u15_u7_n128 ) , .B1( u0_u15_u7_n175 ) );
  INV_X1 u0_u15_u7_U25 (.A( u0_u15_u7_n138 ) , .ZN( u0_u15_u7_n171 ) );
  INV_X1 u0_u15_u7_U26 (.A( u0_u15_u7_n131 ) , .ZN( u0_u15_u7_n177 ) );
  INV_X1 u0_u15_u7_U27 (.A( u0_u15_u7_n110 ) , .ZN( u0_u15_u7_n174 ) );
  NAND2_X1 u0_u15_u7_U28 (.A1( u0_u15_u7_n129 ) , .A2( u0_u15_u7_n132 ) , .ZN( u0_u15_u7_n149 ) );
  NAND2_X1 u0_u15_u7_U29 (.A1( u0_u15_u7_n113 ) , .A2( u0_u15_u7_n124 ) , .ZN( u0_u15_u7_n130 ) );
  INV_X1 u0_u15_u7_U3 (.A( u0_u15_u7_n111 ) , .ZN( u0_u15_u7_n170 ) );
  INV_X1 u0_u15_u7_U30 (.A( u0_u15_u7_n112 ) , .ZN( u0_u15_u7_n173 ) );
  INV_X1 u0_u15_u7_U31 (.A( u0_u15_u7_n128 ) , .ZN( u0_u15_u7_n168 ) );
  INV_X1 u0_u15_u7_U32 (.A( u0_u15_u7_n148 ) , .ZN( u0_u15_u7_n169 ) );
  INV_X1 u0_u15_u7_U33 (.A( u0_u15_u7_n127 ) , .ZN( u0_u15_u7_n179 ) );
  NOR2_X1 u0_u15_u7_U34 (.ZN( u0_u15_u7_n101 ) , .A2( u0_u15_u7_n150 ) , .A1( u0_u15_u7_n156 ) );
  AOI211_X1 u0_u15_u7_U35 (.B( u0_u15_u7_n154 ) , .A( u0_u15_u7_n155 ) , .C1( u0_u15_u7_n156 ) , .ZN( u0_u15_u7_n157 ) , .C2( u0_u15_u7_n172 ) );
  INV_X1 u0_u15_u7_U36 (.A( u0_u15_u7_n153 ) , .ZN( u0_u15_u7_n172 ) );
  AOI211_X1 u0_u15_u7_U37 (.B( u0_u15_u7_n139 ) , .A( u0_u15_u7_n140 ) , .C2( u0_u15_u7_n141 ) , .ZN( u0_u15_u7_n142 ) , .C1( u0_u15_u7_n156 ) );
  NAND4_X1 u0_u15_u7_U38 (.A3( u0_u15_u7_n127 ) , .A2( u0_u15_u7_n128 ) , .A1( u0_u15_u7_n129 ) , .ZN( u0_u15_u7_n141 ) , .A4( u0_u15_u7_n147 ) );
  AOI21_X1 u0_u15_u7_U39 (.A( u0_u15_u7_n137 ) , .B1( u0_u15_u7_n138 ) , .ZN( u0_u15_u7_n139 ) , .B2( u0_u15_u7_n146 ) );
  INV_X1 u0_u15_u7_U4 (.A( u0_u15_u7_n149 ) , .ZN( u0_u15_u7_n175 ) );
  OAI22_X1 u0_u15_u7_U40 (.B1( u0_u15_u7_n136 ) , .ZN( u0_u15_u7_n140 ) , .A1( u0_u15_u7_n153 ) , .B2( u0_u15_u7_n162 ) , .A2( u0_u15_u7_n164 ) );
  AOI21_X1 u0_u15_u7_U41 (.ZN( u0_u15_u7_n123 ) , .B1( u0_u15_u7_n165 ) , .B2( u0_u15_u7_n177 ) , .A( u0_u15_u7_n97 ) );
  AOI21_X1 u0_u15_u7_U42 (.B2( u0_u15_u7_n113 ) , .B1( u0_u15_u7_n124 ) , .A( u0_u15_u7_n125 ) , .ZN( u0_u15_u7_n97 ) );
  INV_X1 u0_u15_u7_U43 (.A( u0_u15_u7_n125 ) , .ZN( u0_u15_u7_n161 ) );
  INV_X1 u0_u15_u7_U44 (.A( u0_u15_u7_n152 ) , .ZN( u0_u15_u7_n162 ) );
  AOI22_X1 u0_u15_u7_U45 (.A2( u0_u15_u7_n114 ) , .ZN( u0_u15_u7_n119 ) , .B1( u0_u15_u7_n130 ) , .A1( u0_u15_u7_n156 ) , .B2( u0_u15_u7_n165 ) );
  NAND2_X1 u0_u15_u7_U46 (.A2( u0_u15_u7_n112 ) , .ZN( u0_u15_u7_n114 ) , .A1( u0_u15_u7_n175 ) );
  AOI22_X1 u0_u15_u7_U47 (.B2( u0_u15_u7_n149 ) , .B1( u0_u15_u7_n150 ) , .A2( u0_u15_u7_n151 ) , .A1( u0_u15_u7_n152 ) , .ZN( u0_u15_u7_n158 ) );
  AND2_X1 u0_u15_u7_U48 (.ZN( u0_u15_u7_n145 ) , .A2( u0_u15_u7_n98 ) , .A1( u0_u15_u7_n99 ) );
  NOR2_X1 u0_u15_u7_U49 (.ZN( u0_u15_u7_n137 ) , .A1( u0_u15_u7_n150 ) , .A2( u0_u15_u7_n161 ) );
  INV_X1 u0_u15_u7_U5 (.A( u0_u15_u7_n154 ) , .ZN( u0_u15_u7_n178 ) );
  AOI21_X1 u0_u15_u7_U50 (.ZN( u0_u15_u7_n105 ) , .B2( u0_u15_u7_n110 ) , .A( u0_u15_u7_n125 ) , .B1( u0_u15_u7_n147 ) );
  NAND2_X1 u0_u15_u7_U51 (.ZN( u0_u15_u7_n146 ) , .A1( u0_u15_u7_n95 ) , .A2( u0_u15_u7_n98 ) );
  NAND2_X1 u0_u15_u7_U52 (.A2( u0_u15_u7_n103 ) , .ZN( u0_u15_u7_n147 ) , .A1( u0_u15_u7_n93 ) );
  NAND2_X1 u0_u15_u7_U53 (.A1( u0_u15_u7_n103 ) , .ZN( u0_u15_u7_n127 ) , .A2( u0_u15_u7_n99 ) );
  OR2_X1 u0_u15_u7_U54 (.ZN( u0_u15_u7_n126 ) , .A2( u0_u15_u7_n152 ) , .A1( u0_u15_u7_n156 ) );
  NAND2_X1 u0_u15_u7_U55 (.A2( u0_u15_u7_n102 ) , .A1( u0_u15_u7_n103 ) , .ZN( u0_u15_u7_n133 ) );
  NAND2_X1 u0_u15_u7_U56 (.ZN( u0_u15_u7_n112 ) , .A2( u0_u15_u7_n96 ) , .A1( u0_u15_u7_n99 ) );
  NAND2_X1 u0_u15_u7_U57 (.A2( u0_u15_u7_n102 ) , .ZN( u0_u15_u7_n128 ) , .A1( u0_u15_u7_n98 ) );
  NAND2_X1 u0_u15_u7_U58 (.A1( u0_u15_u7_n100 ) , .ZN( u0_u15_u7_n113 ) , .A2( u0_u15_u7_n93 ) );
  NAND2_X1 u0_u15_u7_U59 (.A2( u0_u15_u7_n102 ) , .ZN( u0_u15_u7_n124 ) , .A1( u0_u15_u7_n96 ) );
  AOI211_X1 u0_u15_u7_U6 (.ZN( u0_u15_u7_n116 ) , .A( u0_u15_u7_n155 ) , .C1( u0_u15_u7_n161 ) , .C2( u0_u15_u7_n171 ) , .B( u0_u15_u7_n94 ) );
  NAND2_X1 u0_u15_u7_U60 (.ZN( u0_u15_u7_n110 ) , .A1( u0_u15_u7_n95 ) , .A2( u0_u15_u7_n96 ) );
  INV_X1 u0_u15_u7_U61 (.A( u0_u15_u7_n150 ) , .ZN( u0_u15_u7_n164 ) );
  AND2_X1 u0_u15_u7_U62 (.ZN( u0_u15_u7_n134 ) , .A1( u0_u15_u7_n93 ) , .A2( u0_u15_u7_n98 ) );
  NAND2_X1 u0_u15_u7_U63 (.A1( u0_u15_u7_n100 ) , .A2( u0_u15_u7_n102 ) , .ZN( u0_u15_u7_n129 ) );
  NAND2_X1 u0_u15_u7_U64 (.A2( u0_u15_u7_n103 ) , .ZN( u0_u15_u7_n131 ) , .A1( u0_u15_u7_n95 ) );
  NAND2_X1 u0_u15_u7_U65 (.A1( u0_u15_u7_n100 ) , .ZN( u0_u15_u7_n138 ) , .A2( u0_u15_u7_n99 ) );
  NAND2_X1 u0_u15_u7_U66 (.ZN( u0_u15_u7_n132 ) , .A1( u0_u15_u7_n93 ) , .A2( u0_u15_u7_n96 ) );
  NAND2_X1 u0_u15_u7_U67 (.A1( u0_u15_u7_n100 ) , .ZN( u0_u15_u7_n148 ) , .A2( u0_u15_u7_n95 ) );
  NOR2_X1 u0_u15_u7_U68 (.A2( u0_u15_X_47 ) , .ZN( u0_u15_u7_n150 ) , .A1( u0_u15_u7_n163 ) );
  NOR2_X1 u0_u15_u7_U69 (.A2( u0_u15_X_43 ) , .A1( u0_u15_X_44 ) , .ZN( u0_u15_u7_n103 ) );
  OAI222_X1 u0_u15_u7_U7 (.C2( u0_u15_u7_n101 ) , .B2( u0_u15_u7_n111 ) , .A1( u0_u15_u7_n113 ) , .C1( u0_u15_u7_n146 ) , .A2( u0_u15_u7_n162 ) , .B1( u0_u15_u7_n164 ) , .ZN( u0_u15_u7_n94 ) );
  NOR2_X1 u0_u15_u7_U70 (.A2( u0_u15_X_48 ) , .A1( u0_u15_u7_n166 ) , .ZN( u0_u15_u7_n95 ) );
  NOR2_X1 u0_u15_u7_U71 (.A2( u0_u15_X_45 ) , .A1( u0_u15_X_48 ) , .ZN( u0_u15_u7_n99 ) );
  NOR2_X1 u0_u15_u7_U72 (.A2( u0_u15_X_44 ) , .A1( u0_u15_u7_n167 ) , .ZN( u0_u15_u7_n98 ) );
  NOR2_X1 u0_u15_u7_U73 (.A2( u0_u15_X_46 ) , .A1( u0_u15_X_47 ) , .ZN( u0_u15_u7_n152 ) );
  AND2_X1 u0_u15_u7_U74 (.A1( u0_u15_X_47 ) , .ZN( u0_u15_u7_n156 ) , .A2( u0_u15_u7_n163 ) );
  NAND2_X1 u0_u15_u7_U75 (.A2( u0_u15_X_46 ) , .A1( u0_u15_X_47 ) , .ZN( u0_u15_u7_n125 ) );
  AND2_X1 u0_u15_u7_U76 (.A2( u0_u15_X_45 ) , .A1( u0_u15_X_48 ) , .ZN( u0_u15_u7_n102 ) );
  AND2_X1 u0_u15_u7_U77 (.A2( u0_u15_X_43 ) , .A1( u0_u15_X_44 ) , .ZN( u0_u15_u7_n96 ) );
  AND2_X1 u0_u15_u7_U78 (.A1( u0_u15_X_44 ) , .ZN( u0_u15_u7_n100 ) , .A2( u0_u15_u7_n167 ) );
  AND2_X1 u0_u15_u7_U79 (.A1( u0_u15_X_48 ) , .A2( u0_u15_u7_n166 ) , .ZN( u0_u15_u7_n93 ) );
  OAI221_X1 u0_u15_u7_U8 (.C1( u0_u15_u7_n101 ) , .C2( u0_u15_u7_n147 ) , .ZN( u0_u15_u7_n155 ) , .B2( u0_u15_u7_n162 ) , .A( u0_u15_u7_n91 ) , .B1( u0_u15_u7_n92 ) );
  INV_X1 u0_u15_u7_U80 (.A( u0_u15_X_46 ) , .ZN( u0_u15_u7_n163 ) );
  INV_X1 u0_u15_u7_U81 (.A( u0_u15_X_45 ) , .ZN( u0_u15_u7_n166 ) );
  INV_X1 u0_u15_u7_U82 (.A( u0_u15_X_43 ) , .ZN( u0_u15_u7_n167 ) );
  NAND4_X1 u0_u15_u7_U83 (.ZN( u0_out15_5 ) , .A4( u0_u15_u7_n108 ) , .A3( u0_u15_u7_n109 ) , .A1( u0_u15_u7_n116 ) , .A2( u0_u15_u7_n123 ) );
  AOI22_X1 u0_u15_u7_U84 (.ZN( u0_u15_u7_n109 ) , .A2( u0_u15_u7_n126 ) , .B2( u0_u15_u7_n145 ) , .B1( u0_u15_u7_n156 ) , .A1( u0_u15_u7_n171 ) );
  NOR4_X1 u0_u15_u7_U85 (.A4( u0_u15_u7_n104 ) , .A3( u0_u15_u7_n105 ) , .A2( u0_u15_u7_n106 ) , .A1( u0_u15_u7_n107 ) , .ZN( u0_u15_u7_n108 ) );
  NAND4_X1 u0_u15_u7_U86 (.ZN( u0_out15_21 ) , .A4( u0_u15_u7_n157 ) , .A3( u0_u15_u7_n158 ) , .A2( u0_u15_u7_n159 ) , .A1( u0_u15_u7_n160 ) );
  OAI21_X1 u0_u15_u7_U87 (.B1( u0_u15_u7_n145 ) , .ZN( u0_u15_u7_n160 ) , .A( u0_u15_u7_n161 ) , .B2( u0_u15_u7_n177 ) );
  OAI21_X1 u0_u15_u7_U88 (.ZN( u0_u15_u7_n159 ) , .A( u0_u15_u7_n165 ) , .B2( u0_u15_u7_n171 ) , .B1( u0_u15_u7_n174 ) );
  NAND4_X1 u0_u15_u7_U89 (.ZN( u0_out15_15 ) , .A4( u0_u15_u7_n142 ) , .A3( u0_u15_u7_n143 ) , .A2( u0_u15_u7_n144 ) , .A1( u0_u15_u7_n178 ) );
  AND3_X1 u0_u15_u7_U9 (.A3( u0_u15_u7_n110 ) , .A2( u0_u15_u7_n127 ) , .A1( u0_u15_u7_n132 ) , .ZN( u0_u15_u7_n92 ) );
  OR2_X1 u0_u15_u7_U90 (.A2( u0_u15_u7_n125 ) , .A1( u0_u15_u7_n129 ) , .ZN( u0_u15_u7_n144 ) );
  AOI22_X1 u0_u15_u7_U91 (.A2( u0_u15_u7_n126 ) , .ZN( u0_u15_u7_n143 ) , .B2( u0_u15_u7_n165 ) , .B1( u0_u15_u7_n173 ) , .A1( u0_u15_u7_n174 ) );
  NAND4_X1 u0_u15_u7_U92 (.ZN( u0_out15_27 ) , .A4( u0_u15_u7_n118 ) , .A3( u0_u15_u7_n119 ) , .A2( u0_u15_u7_n120 ) , .A1( u0_u15_u7_n121 ) );
  OAI21_X1 u0_u15_u7_U93 (.ZN( u0_u15_u7_n121 ) , .B2( u0_u15_u7_n145 ) , .A( u0_u15_u7_n150 ) , .B1( u0_u15_u7_n174 ) );
  OAI21_X1 u0_u15_u7_U94 (.ZN( u0_u15_u7_n120 ) , .A( u0_u15_u7_n161 ) , .B2( u0_u15_u7_n170 ) , .B1( u0_u15_u7_n179 ) );
  NAND3_X1 u0_u15_u7_U95 (.A3( u0_u15_u7_n146 ) , .A2( u0_u15_u7_n147 ) , .A1( u0_u15_u7_n148 ) , .ZN( u0_u15_u7_n151 ) );
  NAND3_X1 u0_u15_u7_U96 (.A3( u0_u15_u7_n131 ) , .A2( u0_u15_u7_n132 ) , .A1( u0_u15_u7_n133 ) , .ZN( u0_u15_u7_n135 ) );
  XOR2_X1 u0_u4_U13 (.B( u0_K5_42 ) , .A( u0_R3_29 ) , .Z( u0_u4_X_42 ) );
  XOR2_X1 u0_u4_U14 (.B( u0_K5_41 ) , .A( u0_R3_28 ) , .Z( u0_u4_X_41 ) );
  XOR2_X1 u0_u4_U15 (.B( u0_K5_40 ) , .A( u0_R3_27 ) , .Z( u0_u4_X_40 ) );
  XOR2_X1 u0_u4_U17 (.B( u0_K5_39 ) , .A( u0_R3_26 ) , .Z( u0_u4_X_39 ) );
  XOR2_X1 u0_u4_U18 (.B( u0_K5_38 ) , .A( u0_R3_25 ) , .Z( u0_u4_X_38 ) );
  XOR2_X1 u0_u4_U19 (.B( u0_K5_37 ) , .A( u0_R3_24 ) , .Z( u0_u4_X_37 ) );
  XOR2_X1 u0_u4_U20 (.B( u0_K5_36 ) , .A( u0_R3_25 ) , .Z( u0_u4_X_36 ) );
  XOR2_X1 u0_u4_U21 (.B( u0_K5_35 ) , .A( u0_R3_24 ) , .Z( u0_u4_X_35 ) );
  XOR2_X1 u0_u4_U22 (.B( u0_K5_34 ) , .A( u0_R3_23 ) , .Z( u0_u4_X_34 ) );
  XOR2_X1 u0_u4_U23 (.B( u0_K5_33 ) , .A( u0_R3_22 ) , .Z( u0_u4_X_33 ) );
  XOR2_X1 u0_u4_U24 (.B( u0_K5_32 ) , .A( u0_R3_21 ) , .Z( u0_u4_X_32 ) );
  XOR2_X1 u0_u4_U25 (.B( u0_K5_31 ) , .A( u0_R3_20 ) , .Z( u0_u4_X_31 ) );
  XOR2_X1 u0_u4_U26 (.B( u0_K5_30 ) , .A( u0_R3_21 ) , .Z( u0_u4_X_30 ) );
  XOR2_X1 u0_u4_U28 (.B( u0_K5_29 ) , .A( u0_R3_20 ) , .Z( u0_u4_X_29 ) );
  XOR2_X1 u0_u4_U29 (.B( u0_K5_28 ) , .A( u0_R3_19 ) , .Z( u0_u4_X_28 ) );
  XOR2_X1 u0_u4_U30 (.B( u0_K5_27 ) , .A( u0_R3_18 ) , .Z( u0_u4_X_27 ) );
  XOR2_X1 u0_u4_U31 (.B( u0_K5_26 ) , .A( u0_R3_17 ) , .Z( u0_u4_X_26 ) );
  XOR2_X1 u0_u4_U32 (.B( u0_K5_25 ) , .A( u0_R3_16 ) , .Z( u0_u4_X_25 ) );
  OAI22_X1 u0_u4_u4_U10 (.B2( u0_u4_u4_n135 ) , .ZN( u0_u4_u4_n137 ) , .B1( u0_u4_u4_n153 ) , .A1( u0_u4_u4_n155 ) , .A2( u0_u4_u4_n171 ) );
  AND3_X1 u0_u4_u4_U11 (.A2( u0_u4_u4_n134 ) , .ZN( u0_u4_u4_n135 ) , .A3( u0_u4_u4_n145 ) , .A1( u0_u4_u4_n157 ) );
  NAND2_X1 u0_u4_u4_U12 (.ZN( u0_u4_u4_n132 ) , .A2( u0_u4_u4_n170 ) , .A1( u0_u4_u4_n173 ) );
  AOI21_X1 u0_u4_u4_U13 (.B2( u0_u4_u4_n160 ) , .B1( u0_u4_u4_n161 ) , .ZN( u0_u4_u4_n162 ) , .A( u0_u4_u4_n170 ) );
  AOI21_X1 u0_u4_u4_U14 (.ZN( u0_u4_u4_n107 ) , .B2( u0_u4_u4_n143 ) , .A( u0_u4_u4_n174 ) , .B1( u0_u4_u4_n184 ) );
  AOI21_X1 u0_u4_u4_U15 (.B2( u0_u4_u4_n158 ) , .B1( u0_u4_u4_n159 ) , .ZN( u0_u4_u4_n163 ) , .A( u0_u4_u4_n174 ) );
  AOI21_X1 u0_u4_u4_U16 (.A( u0_u4_u4_n153 ) , .B2( u0_u4_u4_n154 ) , .B1( u0_u4_u4_n155 ) , .ZN( u0_u4_u4_n165 ) );
  AOI21_X1 u0_u4_u4_U17 (.A( u0_u4_u4_n156 ) , .B2( u0_u4_u4_n157 ) , .ZN( u0_u4_u4_n164 ) , .B1( u0_u4_u4_n184 ) );
  INV_X1 u0_u4_u4_U18 (.A( u0_u4_u4_n138 ) , .ZN( u0_u4_u4_n170 ) );
  AND2_X1 u0_u4_u4_U19 (.A2( u0_u4_u4_n120 ) , .ZN( u0_u4_u4_n155 ) , .A1( u0_u4_u4_n160 ) );
  INV_X1 u0_u4_u4_U20 (.A( u0_u4_u4_n156 ) , .ZN( u0_u4_u4_n175 ) );
  NAND2_X1 u0_u4_u4_U21 (.A2( u0_u4_u4_n118 ) , .ZN( u0_u4_u4_n131 ) , .A1( u0_u4_u4_n147 ) );
  NAND2_X1 u0_u4_u4_U22 (.A1( u0_u4_u4_n119 ) , .A2( u0_u4_u4_n120 ) , .ZN( u0_u4_u4_n130 ) );
  NAND2_X1 u0_u4_u4_U23 (.ZN( u0_u4_u4_n117 ) , .A2( u0_u4_u4_n118 ) , .A1( u0_u4_u4_n148 ) );
  NAND2_X1 u0_u4_u4_U24 (.ZN( u0_u4_u4_n129 ) , .A1( u0_u4_u4_n134 ) , .A2( u0_u4_u4_n148 ) );
  AND3_X1 u0_u4_u4_U25 (.A1( u0_u4_u4_n119 ) , .A2( u0_u4_u4_n143 ) , .A3( u0_u4_u4_n154 ) , .ZN( u0_u4_u4_n161 ) );
  AND2_X1 u0_u4_u4_U26 (.A1( u0_u4_u4_n145 ) , .A2( u0_u4_u4_n147 ) , .ZN( u0_u4_u4_n159 ) );
  OR3_X1 u0_u4_u4_U27 (.A3( u0_u4_u4_n114 ) , .A2( u0_u4_u4_n115 ) , .A1( u0_u4_u4_n116 ) , .ZN( u0_u4_u4_n136 ) );
  AOI21_X1 u0_u4_u4_U28 (.A( u0_u4_u4_n113 ) , .ZN( u0_u4_u4_n116 ) , .B2( u0_u4_u4_n173 ) , .B1( u0_u4_u4_n174 ) );
  AOI21_X1 u0_u4_u4_U29 (.ZN( u0_u4_u4_n115 ) , .B2( u0_u4_u4_n145 ) , .B1( u0_u4_u4_n146 ) , .A( u0_u4_u4_n156 ) );
  NOR2_X1 u0_u4_u4_U3 (.ZN( u0_u4_u4_n121 ) , .A1( u0_u4_u4_n181 ) , .A2( u0_u4_u4_n182 ) );
  OAI22_X1 u0_u4_u4_U30 (.ZN( u0_u4_u4_n114 ) , .A2( u0_u4_u4_n121 ) , .B1( u0_u4_u4_n160 ) , .B2( u0_u4_u4_n170 ) , .A1( u0_u4_u4_n171 ) );
  INV_X1 u0_u4_u4_U31 (.A( u0_u4_u4_n158 ) , .ZN( u0_u4_u4_n182 ) );
  INV_X1 u0_u4_u4_U32 (.ZN( u0_u4_u4_n181 ) , .A( u0_u4_u4_n96 ) );
  INV_X1 u0_u4_u4_U33 (.A( u0_u4_u4_n144 ) , .ZN( u0_u4_u4_n179 ) );
  INV_X1 u0_u4_u4_U34 (.A( u0_u4_u4_n157 ) , .ZN( u0_u4_u4_n178 ) );
  NAND2_X1 u0_u4_u4_U35 (.A2( u0_u4_u4_n154 ) , .A1( u0_u4_u4_n96 ) , .ZN( u0_u4_u4_n97 ) );
  INV_X1 u0_u4_u4_U36 (.ZN( u0_u4_u4_n186 ) , .A( u0_u4_u4_n95 ) );
  OAI221_X1 u0_u4_u4_U37 (.C1( u0_u4_u4_n134 ) , .B1( u0_u4_u4_n158 ) , .B2( u0_u4_u4_n171 ) , .C2( u0_u4_u4_n173 ) , .A( u0_u4_u4_n94 ) , .ZN( u0_u4_u4_n95 ) );
  AOI222_X1 u0_u4_u4_U38 (.B2( u0_u4_u4_n132 ) , .A1( u0_u4_u4_n138 ) , .C2( u0_u4_u4_n175 ) , .A2( u0_u4_u4_n179 ) , .C1( u0_u4_u4_n181 ) , .B1( u0_u4_u4_n185 ) , .ZN( u0_u4_u4_n94 ) );
  INV_X1 u0_u4_u4_U39 (.A( u0_u4_u4_n113 ) , .ZN( u0_u4_u4_n185 ) );
  INV_X1 u0_u4_u4_U4 (.A( u0_u4_u4_n117 ) , .ZN( u0_u4_u4_n184 ) );
  INV_X1 u0_u4_u4_U40 (.A( u0_u4_u4_n143 ) , .ZN( u0_u4_u4_n183 ) );
  NOR2_X1 u0_u4_u4_U41 (.ZN( u0_u4_u4_n138 ) , .A1( u0_u4_u4_n168 ) , .A2( u0_u4_u4_n169 ) );
  NOR2_X1 u0_u4_u4_U42 (.A1( u0_u4_u4_n150 ) , .A2( u0_u4_u4_n152 ) , .ZN( u0_u4_u4_n153 ) );
  NOR2_X1 u0_u4_u4_U43 (.A2( u0_u4_u4_n128 ) , .A1( u0_u4_u4_n138 ) , .ZN( u0_u4_u4_n156 ) );
  AOI22_X1 u0_u4_u4_U44 (.B2( u0_u4_u4_n122 ) , .A1( u0_u4_u4_n123 ) , .ZN( u0_u4_u4_n124 ) , .B1( u0_u4_u4_n128 ) , .A2( u0_u4_u4_n172 ) );
  INV_X1 u0_u4_u4_U45 (.A( u0_u4_u4_n153 ) , .ZN( u0_u4_u4_n172 ) );
  NAND2_X1 u0_u4_u4_U46 (.A2( u0_u4_u4_n120 ) , .ZN( u0_u4_u4_n123 ) , .A1( u0_u4_u4_n161 ) );
  AOI22_X1 u0_u4_u4_U47 (.B2( u0_u4_u4_n132 ) , .A2( u0_u4_u4_n133 ) , .ZN( u0_u4_u4_n140 ) , .A1( u0_u4_u4_n150 ) , .B1( u0_u4_u4_n179 ) );
  NAND2_X1 u0_u4_u4_U48 (.ZN( u0_u4_u4_n133 ) , .A2( u0_u4_u4_n146 ) , .A1( u0_u4_u4_n154 ) );
  NAND2_X1 u0_u4_u4_U49 (.A1( u0_u4_u4_n103 ) , .ZN( u0_u4_u4_n154 ) , .A2( u0_u4_u4_n98 ) );
  NOR4_X1 u0_u4_u4_U5 (.A4( u0_u4_u4_n106 ) , .A3( u0_u4_u4_n107 ) , .A2( u0_u4_u4_n108 ) , .A1( u0_u4_u4_n109 ) , .ZN( u0_u4_u4_n110 ) );
  NAND2_X1 u0_u4_u4_U50 (.A1( u0_u4_u4_n101 ) , .ZN( u0_u4_u4_n158 ) , .A2( u0_u4_u4_n99 ) );
  AOI21_X1 u0_u4_u4_U51 (.ZN( u0_u4_u4_n127 ) , .A( u0_u4_u4_n136 ) , .B2( u0_u4_u4_n150 ) , .B1( u0_u4_u4_n180 ) );
  INV_X1 u0_u4_u4_U52 (.A( u0_u4_u4_n160 ) , .ZN( u0_u4_u4_n180 ) );
  NAND2_X1 u0_u4_u4_U53 (.A2( u0_u4_u4_n104 ) , .A1( u0_u4_u4_n105 ) , .ZN( u0_u4_u4_n146 ) );
  NAND2_X1 u0_u4_u4_U54 (.A2( u0_u4_u4_n101 ) , .A1( u0_u4_u4_n102 ) , .ZN( u0_u4_u4_n160 ) );
  NAND2_X1 u0_u4_u4_U55 (.ZN( u0_u4_u4_n134 ) , .A1( u0_u4_u4_n98 ) , .A2( u0_u4_u4_n99 ) );
  NAND2_X1 u0_u4_u4_U56 (.A1( u0_u4_u4_n103 ) , .A2( u0_u4_u4_n104 ) , .ZN( u0_u4_u4_n143 ) );
  NAND2_X1 u0_u4_u4_U57 (.A2( u0_u4_u4_n105 ) , .ZN( u0_u4_u4_n145 ) , .A1( u0_u4_u4_n98 ) );
  NAND2_X1 u0_u4_u4_U58 (.A1( u0_u4_u4_n100 ) , .A2( u0_u4_u4_n105 ) , .ZN( u0_u4_u4_n120 ) );
  NAND2_X1 u0_u4_u4_U59 (.A1( u0_u4_u4_n102 ) , .A2( u0_u4_u4_n104 ) , .ZN( u0_u4_u4_n148 ) );
  AOI21_X1 u0_u4_u4_U6 (.ZN( u0_u4_u4_n106 ) , .B2( u0_u4_u4_n146 ) , .B1( u0_u4_u4_n158 ) , .A( u0_u4_u4_n170 ) );
  NAND2_X1 u0_u4_u4_U60 (.A2( u0_u4_u4_n100 ) , .A1( u0_u4_u4_n103 ) , .ZN( u0_u4_u4_n157 ) );
  INV_X1 u0_u4_u4_U61 (.A( u0_u4_u4_n150 ) , .ZN( u0_u4_u4_n173 ) );
  INV_X1 u0_u4_u4_U62 (.A( u0_u4_u4_n152 ) , .ZN( u0_u4_u4_n171 ) );
  NAND2_X1 u0_u4_u4_U63 (.A1( u0_u4_u4_n100 ) , .ZN( u0_u4_u4_n118 ) , .A2( u0_u4_u4_n99 ) );
  NAND2_X1 u0_u4_u4_U64 (.A2( u0_u4_u4_n100 ) , .A1( u0_u4_u4_n102 ) , .ZN( u0_u4_u4_n144 ) );
  NAND2_X1 u0_u4_u4_U65 (.A2( u0_u4_u4_n101 ) , .A1( u0_u4_u4_n105 ) , .ZN( u0_u4_u4_n96 ) );
  INV_X1 u0_u4_u4_U66 (.A( u0_u4_u4_n128 ) , .ZN( u0_u4_u4_n174 ) );
  NAND2_X1 u0_u4_u4_U67 (.A2( u0_u4_u4_n102 ) , .ZN( u0_u4_u4_n119 ) , .A1( u0_u4_u4_n98 ) );
  NAND2_X1 u0_u4_u4_U68 (.A2( u0_u4_u4_n101 ) , .A1( u0_u4_u4_n103 ) , .ZN( u0_u4_u4_n147 ) );
  NAND2_X1 u0_u4_u4_U69 (.A2( u0_u4_u4_n104 ) , .ZN( u0_u4_u4_n113 ) , .A1( u0_u4_u4_n99 ) );
  AOI21_X1 u0_u4_u4_U7 (.ZN( u0_u4_u4_n108 ) , .B2( u0_u4_u4_n134 ) , .B1( u0_u4_u4_n155 ) , .A( u0_u4_u4_n156 ) );
  NOR2_X1 u0_u4_u4_U70 (.A2( u0_u4_X_28 ) , .ZN( u0_u4_u4_n150 ) , .A1( u0_u4_u4_n168 ) );
  NOR2_X1 u0_u4_u4_U71 (.A2( u0_u4_X_29 ) , .ZN( u0_u4_u4_n152 ) , .A1( u0_u4_u4_n169 ) );
  NOR2_X1 u0_u4_u4_U72 (.A2( u0_u4_X_30 ) , .ZN( u0_u4_u4_n105 ) , .A1( u0_u4_u4_n176 ) );
  NOR2_X1 u0_u4_u4_U73 (.A2( u0_u4_X_26 ) , .ZN( u0_u4_u4_n100 ) , .A1( u0_u4_u4_n177 ) );
  NOR2_X1 u0_u4_u4_U74 (.A2( u0_u4_X_28 ) , .A1( u0_u4_X_29 ) , .ZN( u0_u4_u4_n128 ) );
  NOR2_X1 u0_u4_u4_U75 (.A2( u0_u4_X_27 ) , .A1( u0_u4_X_30 ) , .ZN( u0_u4_u4_n102 ) );
  NOR2_X1 u0_u4_u4_U76 (.A2( u0_u4_X_25 ) , .A1( u0_u4_X_26 ) , .ZN( u0_u4_u4_n98 ) );
  AND2_X1 u0_u4_u4_U77 (.A2( u0_u4_X_25 ) , .A1( u0_u4_X_26 ) , .ZN( u0_u4_u4_n104 ) );
  AND2_X1 u0_u4_u4_U78 (.A1( u0_u4_X_30 ) , .A2( u0_u4_u4_n176 ) , .ZN( u0_u4_u4_n99 ) );
  AND2_X1 u0_u4_u4_U79 (.A1( u0_u4_X_26 ) , .ZN( u0_u4_u4_n101 ) , .A2( u0_u4_u4_n177 ) );
  AOI21_X1 u0_u4_u4_U8 (.ZN( u0_u4_u4_n109 ) , .A( u0_u4_u4_n153 ) , .B1( u0_u4_u4_n159 ) , .B2( u0_u4_u4_n184 ) );
  AND2_X1 u0_u4_u4_U80 (.A1( u0_u4_X_27 ) , .A2( u0_u4_X_30 ) , .ZN( u0_u4_u4_n103 ) );
  INV_X1 u0_u4_u4_U81 (.A( u0_u4_X_28 ) , .ZN( u0_u4_u4_n169 ) );
  INV_X1 u0_u4_u4_U82 (.A( u0_u4_X_29 ) , .ZN( u0_u4_u4_n168 ) );
  INV_X1 u0_u4_u4_U83 (.A( u0_u4_X_25 ) , .ZN( u0_u4_u4_n177 ) );
  INV_X1 u0_u4_u4_U84 (.A( u0_u4_X_27 ) , .ZN( u0_u4_u4_n176 ) );
  NAND4_X1 u0_u4_u4_U85 (.ZN( u0_out4_25 ) , .A4( u0_u4_u4_n139 ) , .A3( u0_u4_u4_n140 ) , .A2( u0_u4_u4_n141 ) , .A1( u0_u4_u4_n142 ) );
  OAI21_X1 u0_u4_u4_U86 (.B2( u0_u4_u4_n131 ) , .ZN( u0_u4_u4_n141 ) , .A( u0_u4_u4_n175 ) , .B1( u0_u4_u4_n183 ) );
  OAI21_X1 u0_u4_u4_U87 (.A( u0_u4_u4_n128 ) , .B2( u0_u4_u4_n129 ) , .B1( u0_u4_u4_n130 ) , .ZN( u0_u4_u4_n142 ) );
  NAND4_X1 u0_u4_u4_U88 (.ZN( u0_out4_14 ) , .A4( u0_u4_u4_n124 ) , .A3( u0_u4_u4_n125 ) , .A2( u0_u4_u4_n126 ) , .A1( u0_u4_u4_n127 ) );
  AOI22_X1 u0_u4_u4_U89 (.B2( u0_u4_u4_n117 ) , .ZN( u0_u4_u4_n126 ) , .A1( u0_u4_u4_n129 ) , .B1( u0_u4_u4_n152 ) , .A2( u0_u4_u4_n175 ) );
  AOI211_X1 u0_u4_u4_U9 (.B( u0_u4_u4_n136 ) , .A( u0_u4_u4_n137 ) , .C2( u0_u4_u4_n138 ) , .ZN( u0_u4_u4_n139 ) , .C1( u0_u4_u4_n182 ) );
  AOI22_X1 u0_u4_u4_U90 (.ZN( u0_u4_u4_n125 ) , .B2( u0_u4_u4_n131 ) , .A2( u0_u4_u4_n132 ) , .B1( u0_u4_u4_n138 ) , .A1( u0_u4_u4_n178 ) );
  NAND4_X1 u0_u4_u4_U91 (.ZN( u0_out4_8 ) , .A4( u0_u4_u4_n110 ) , .A3( u0_u4_u4_n111 ) , .A2( u0_u4_u4_n112 ) , .A1( u0_u4_u4_n186 ) );
  NAND2_X1 u0_u4_u4_U92 (.ZN( u0_u4_u4_n112 ) , .A2( u0_u4_u4_n130 ) , .A1( u0_u4_u4_n150 ) );
  AOI22_X1 u0_u4_u4_U93 (.ZN( u0_u4_u4_n111 ) , .B2( u0_u4_u4_n132 ) , .A1( u0_u4_u4_n152 ) , .B1( u0_u4_u4_n178 ) , .A2( u0_u4_u4_n97 ) );
  AOI22_X1 u0_u4_u4_U94 (.B2( u0_u4_u4_n149 ) , .B1( u0_u4_u4_n150 ) , .A2( u0_u4_u4_n151 ) , .A1( u0_u4_u4_n152 ) , .ZN( u0_u4_u4_n167 ) );
  NOR4_X1 u0_u4_u4_U95 (.A4( u0_u4_u4_n162 ) , .A3( u0_u4_u4_n163 ) , .A2( u0_u4_u4_n164 ) , .A1( u0_u4_u4_n165 ) , .ZN( u0_u4_u4_n166 ) );
  NAND3_X1 u0_u4_u4_U96 (.ZN( u0_out4_3 ) , .A3( u0_u4_u4_n166 ) , .A1( u0_u4_u4_n167 ) , .A2( u0_u4_u4_n186 ) );
  NAND3_X1 u0_u4_u4_U97 (.A3( u0_u4_u4_n146 ) , .A2( u0_u4_u4_n147 ) , .A1( u0_u4_u4_n148 ) , .ZN( u0_u4_u4_n149 ) );
  NAND3_X1 u0_u4_u4_U98 (.A3( u0_u4_u4_n143 ) , .A2( u0_u4_u4_n144 ) , .A1( u0_u4_u4_n145 ) , .ZN( u0_u4_u4_n151 ) );
  NAND3_X1 u0_u4_u4_U99 (.A3( u0_u4_u4_n121 ) , .ZN( u0_u4_u4_n122 ) , .A2( u0_u4_u4_n144 ) , .A1( u0_u4_u4_n154 ) );
  NOR2_X1 u0_u4_u5_U10 (.ZN( u0_u4_u5_n135 ) , .A1( u0_u4_u5_n173 ) , .A2( u0_u4_u5_n176 ) );
  NOR3_X1 u0_u4_u5_U100 (.A3( u0_u4_u5_n141 ) , .A1( u0_u4_u5_n142 ) , .ZN( u0_u4_u5_n143 ) , .A2( u0_u4_u5_n191 ) );
  NAND4_X1 u0_u4_u5_U101 (.ZN( u0_out4_4 ) , .A4( u0_u4_u5_n112 ) , .A2( u0_u4_u5_n113 ) , .A1( u0_u4_u5_n114 ) , .A3( u0_u4_u5_n195 ) );
  AOI211_X1 u0_u4_u5_U102 (.A( u0_u4_u5_n110 ) , .C1( u0_u4_u5_n111 ) , .ZN( u0_u4_u5_n112 ) , .B( u0_u4_u5_n118 ) , .C2( u0_u4_u5_n177 ) );
  INV_X1 u0_u4_u5_U103 (.A( u0_u4_u5_n102 ) , .ZN( u0_u4_u5_n195 ) );
  NAND3_X1 u0_u4_u5_U104 (.A2( u0_u4_u5_n154 ) , .A3( u0_u4_u5_n158 ) , .A1( u0_u4_u5_n161 ) , .ZN( u0_u4_u5_n99 ) );
  INV_X1 u0_u4_u5_U11 (.A( u0_u4_u5_n121 ) , .ZN( u0_u4_u5_n177 ) );
  NOR2_X1 u0_u4_u5_U12 (.ZN( u0_u4_u5_n160 ) , .A2( u0_u4_u5_n173 ) , .A1( u0_u4_u5_n177 ) );
  INV_X1 u0_u4_u5_U13 (.A( u0_u4_u5_n150 ) , .ZN( u0_u4_u5_n174 ) );
  AOI21_X1 u0_u4_u5_U14 (.A( u0_u4_u5_n160 ) , .B2( u0_u4_u5_n161 ) , .ZN( u0_u4_u5_n162 ) , .B1( u0_u4_u5_n192 ) );
  INV_X1 u0_u4_u5_U15 (.A( u0_u4_u5_n159 ) , .ZN( u0_u4_u5_n192 ) );
  AOI21_X1 u0_u4_u5_U16 (.A( u0_u4_u5_n156 ) , .B2( u0_u4_u5_n157 ) , .B1( u0_u4_u5_n158 ) , .ZN( u0_u4_u5_n163 ) );
  AOI21_X1 u0_u4_u5_U17 (.B2( u0_u4_u5_n139 ) , .B1( u0_u4_u5_n140 ) , .ZN( u0_u4_u5_n141 ) , .A( u0_u4_u5_n150 ) );
  OAI21_X1 u0_u4_u5_U18 (.A( u0_u4_u5_n133 ) , .B2( u0_u4_u5_n134 ) , .B1( u0_u4_u5_n135 ) , .ZN( u0_u4_u5_n142 ) );
  OAI21_X1 u0_u4_u5_U19 (.ZN( u0_u4_u5_n133 ) , .B2( u0_u4_u5_n147 ) , .A( u0_u4_u5_n173 ) , .B1( u0_u4_u5_n188 ) );
  NAND2_X1 u0_u4_u5_U20 (.A2( u0_u4_u5_n119 ) , .A1( u0_u4_u5_n123 ) , .ZN( u0_u4_u5_n137 ) );
  INV_X1 u0_u4_u5_U21 (.A( u0_u4_u5_n155 ) , .ZN( u0_u4_u5_n194 ) );
  NAND2_X1 u0_u4_u5_U22 (.A1( u0_u4_u5_n121 ) , .ZN( u0_u4_u5_n132 ) , .A2( u0_u4_u5_n172 ) );
  NAND2_X1 u0_u4_u5_U23 (.A2( u0_u4_u5_n122 ) , .ZN( u0_u4_u5_n136 ) , .A1( u0_u4_u5_n154 ) );
  NAND2_X1 u0_u4_u5_U24 (.A2( u0_u4_u5_n119 ) , .A1( u0_u4_u5_n120 ) , .ZN( u0_u4_u5_n159 ) );
  INV_X1 u0_u4_u5_U25 (.A( u0_u4_u5_n156 ) , .ZN( u0_u4_u5_n175 ) );
  INV_X1 u0_u4_u5_U26 (.A( u0_u4_u5_n158 ) , .ZN( u0_u4_u5_n188 ) );
  INV_X1 u0_u4_u5_U27 (.A( u0_u4_u5_n152 ) , .ZN( u0_u4_u5_n179 ) );
  INV_X1 u0_u4_u5_U28 (.A( u0_u4_u5_n140 ) , .ZN( u0_u4_u5_n182 ) );
  INV_X1 u0_u4_u5_U29 (.A( u0_u4_u5_n151 ) , .ZN( u0_u4_u5_n183 ) );
  NOR2_X1 u0_u4_u5_U3 (.ZN( u0_u4_u5_n134 ) , .A1( u0_u4_u5_n183 ) , .A2( u0_u4_u5_n190 ) );
  INV_X1 u0_u4_u5_U30 (.A( u0_u4_u5_n123 ) , .ZN( u0_u4_u5_n185 ) );
  INV_X1 u0_u4_u5_U31 (.A( u0_u4_u5_n161 ) , .ZN( u0_u4_u5_n184 ) );
  INV_X1 u0_u4_u5_U32 (.A( u0_u4_u5_n139 ) , .ZN( u0_u4_u5_n189 ) );
  INV_X1 u0_u4_u5_U33 (.A( u0_u4_u5_n157 ) , .ZN( u0_u4_u5_n190 ) );
  INV_X1 u0_u4_u5_U34 (.A( u0_u4_u5_n120 ) , .ZN( u0_u4_u5_n193 ) );
  NAND2_X1 u0_u4_u5_U35 (.ZN( u0_u4_u5_n111 ) , .A1( u0_u4_u5_n140 ) , .A2( u0_u4_u5_n155 ) );
  INV_X1 u0_u4_u5_U36 (.A( u0_u4_u5_n117 ) , .ZN( u0_u4_u5_n196 ) );
  OAI221_X1 u0_u4_u5_U37 (.A( u0_u4_u5_n116 ) , .ZN( u0_u4_u5_n117 ) , .B2( u0_u4_u5_n119 ) , .C1( u0_u4_u5_n153 ) , .C2( u0_u4_u5_n158 ) , .B1( u0_u4_u5_n172 ) );
  AOI222_X1 u0_u4_u5_U38 (.ZN( u0_u4_u5_n116 ) , .B2( u0_u4_u5_n145 ) , .C1( u0_u4_u5_n148 ) , .A2( u0_u4_u5_n174 ) , .C2( u0_u4_u5_n177 ) , .B1( u0_u4_u5_n187 ) , .A1( u0_u4_u5_n193 ) );
  INV_X1 u0_u4_u5_U39 (.A( u0_u4_u5_n115 ) , .ZN( u0_u4_u5_n187 ) );
  INV_X1 u0_u4_u5_U4 (.A( u0_u4_u5_n138 ) , .ZN( u0_u4_u5_n191 ) );
  NOR2_X1 u0_u4_u5_U40 (.ZN( u0_u4_u5_n100 ) , .A1( u0_u4_u5_n170 ) , .A2( u0_u4_u5_n180 ) );
  OAI221_X1 u0_u4_u5_U41 (.A( u0_u4_u5_n101 ) , .ZN( u0_u4_u5_n102 ) , .C2( u0_u4_u5_n115 ) , .C1( u0_u4_u5_n126 ) , .B1( u0_u4_u5_n134 ) , .B2( u0_u4_u5_n160 ) );
  OAI21_X1 u0_u4_u5_U42 (.ZN( u0_u4_u5_n101 ) , .B1( u0_u4_u5_n137 ) , .A( u0_u4_u5_n146 ) , .B2( u0_u4_u5_n147 ) );
  AOI22_X1 u0_u4_u5_U43 (.B2( u0_u4_u5_n131 ) , .A2( u0_u4_u5_n146 ) , .ZN( u0_u4_u5_n169 ) , .B1( u0_u4_u5_n174 ) , .A1( u0_u4_u5_n185 ) );
  NOR2_X1 u0_u4_u5_U44 (.A1( u0_u4_u5_n146 ) , .ZN( u0_u4_u5_n150 ) , .A2( u0_u4_u5_n173 ) );
  AOI21_X1 u0_u4_u5_U45 (.A( u0_u4_u5_n118 ) , .B2( u0_u4_u5_n145 ) , .ZN( u0_u4_u5_n168 ) , .B1( u0_u4_u5_n186 ) );
  INV_X1 u0_u4_u5_U46 (.A( u0_u4_u5_n122 ) , .ZN( u0_u4_u5_n186 ) );
  NOR2_X1 u0_u4_u5_U47 (.A1( u0_u4_u5_n146 ) , .ZN( u0_u4_u5_n152 ) , .A2( u0_u4_u5_n176 ) );
  NOR2_X1 u0_u4_u5_U48 (.A1( u0_u4_u5_n115 ) , .ZN( u0_u4_u5_n118 ) , .A2( u0_u4_u5_n153 ) );
  NOR2_X1 u0_u4_u5_U49 (.A2( u0_u4_u5_n145 ) , .ZN( u0_u4_u5_n156 ) , .A1( u0_u4_u5_n174 ) );
  OAI21_X1 u0_u4_u5_U5 (.B2( u0_u4_u5_n136 ) , .B1( u0_u4_u5_n137 ) , .ZN( u0_u4_u5_n138 ) , .A( u0_u4_u5_n177 ) );
  NOR2_X1 u0_u4_u5_U50 (.ZN( u0_u4_u5_n121 ) , .A2( u0_u4_u5_n145 ) , .A1( u0_u4_u5_n176 ) );
  AOI22_X1 u0_u4_u5_U51 (.ZN( u0_u4_u5_n114 ) , .A2( u0_u4_u5_n137 ) , .A1( u0_u4_u5_n145 ) , .B2( u0_u4_u5_n175 ) , .B1( u0_u4_u5_n193 ) );
  OAI211_X1 u0_u4_u5_U52 (.B( u0_u4_u5_n124 ) , .A( u0_u4_u5_n125 ) , .C2( u0_u4_u5_n126 ) , .C1( u0_u4_u5_n127 ) , .ZN( u0_u4_u5_n128 ) );
  NOR3_X1 u0_u4_u5_U53 (.ZN( u0_u4_u5_n127 ) , .A1( u0_u4_u5_n136 ) , .A3( u0_u4_u5_n148 ) , .A2( u0_u4_u5_n182 ) );
  OAI21_X1 u0_u4_u5_U54 (.ZN( u0_u4_u5_n124 ) , .A( u0_u4_u5_n177 ) , .B2( u0_u4_u5_n183 ) , .B1( u0_u4_u5_n189 ) );
  OAI21_X1 u0_u4_u5_U55 (.ZN( u0_u4_u5_n125 ) , .A( u0_u4_u5_n174 ) , .B2( u0_u4_u5_n185 ) , .B1( u0_u4_u5_n190 ) );
  AOI21_X1 u0_u4_u5_U56 (.A( u0_u4_u5_n153 ) , .B2( u0_u4_u5_n154 ) , .B1( u0_u4_u5_n155 ) , .ZN( u0_u4_u5_n164 ) );
  AOI21_X1 u0_u4_u5_U57 (.ZN( u0_u4_u5_n110 ) , .B1( u0_u4_u5_n122 ) , .B2( u0_u4_u5_n139 ) , .A( u0_u4_u5_n153 ) );
  INV_X1 u0_u4_u5_U58 (.A( u0_u4_u5_n153 ) , .ZN( u0_u4_u5_n176 ) );
  INV_X1 u0_u4_u5_U59 (.A( u0_u4_u5_n126 ) , .ZN( u0_u4_u5_n173 ) );
  AOI222_X1 u0_u4_u5_U6 (.ZN( u0_u4_u5_n113 ) , .A1( u0_u4_u5_n131 ) , .C1( u0_u4_u5_n148 ) , .B2( u0_u4_u5_n174 ) , .C2( u0_u4_u5_n178 ) , .A2( u0_u4_u5_n179 ) , .B1( u0_u4_u5_n99 ) );
  AND2_X1 u0_u4_u5_U60 (.A2( u0_u4_u5_n104 ) , .A1( u0_u4_u5_n107 ) , .ZN( u0_u4_u5_n147 ) );
  AND2_X1 u0_u4_u5_U61 (.A2( u0_u4_u5_n104 ) , .A1( u0_u4_u5_n108 ) , .ZN( u0_u4_u5_n148 ) );
  NAND2_X1 u0_u4_u5_U62 (.A1( u0_u4_u5_n105 ) , .A2( u0_u4_u5_n106 ) , .ZN( u0_u4_u5_n158 ) );
  NAND2_X1 u0_u4_u5_U63 (.A2( u0_u4_u5_n108 ) , .A1( u0_u4_u5_n109 ) , .ZN( u0_u4_u5_n139 ) );
  NAND2_X1 u0_u4_u5_U64 (.A1( u0_u4_u5_n106 ) , .A2( u0_u4_u5_n108 ) , .ZN( u0_u4_u5_n119 ) );
  NAND2_X1 u0_u4_u5_U65 (.A2( u0_u4_u5_n103 ) , .A1( u0_u4_u5_n105 ) , .ZN( u0_u4_u5_n140 ) );
  NAND2_X1 u0_u4_u5_U66 (.A2( u0_u4_u5_n104 ) , .A1( u0_u4_u5_n105 ) , .ZN( u0_u4_u5_n155 ) );
  NAND2_X1 u0_u4_u5_U67 (.A2( u0_u4_u5_n106 ) , .A1( u0_u4_u5_n107 ) , .ZN( u0_u4_u5_n122 ) );
  NAND2_X1 u0_u4_u5_U68 (.A2( u0_u4_u5_n100 ) , .A1( u0_u4_u5_n106 ) , .ZN( u0_u4_u5_n115 ) );
  NAND2_X1 u0_u4_u5_U69 (.A2( u0_u4_u5_n100 ) , .A1( u0_u4_u5_n103 ) , .ZN( u0_u4_u5_n161 ) );
  INV_X1 u0_u4_u5_U7 (.A( u0_u4_u5_n135 ) , .ZN( u0_u4_u5_n178 ) );
  NAND2_X1 u0_u4_u5_U70 (.A1( u0_u4_u5_n105 ) , .A2( u0_u4_u5_n109 ) , .ZN( u0_u4_u5_n154 ) );
  INV_X1 u0_u4_u5_U71 (.A( u0_u4_u5_n146 ) , .ZN( u0_u4_u5_n172 ) );
  NAND2_X1 u0_u4_u5_U72 (.A1( u0_u4_u5_n103 ) , .A2( u0_u4_u5_n108 ) , .ZN( u0_u4_u5_n123 ) );
  NAND2_X1 u0_u4_u5_U73 (.A2( u0_u4_u5_n103 ) , .A1( u0_u4_u5_n107 ) , .ZN( u0_u4_u5_n151 ) );
  NAND2_X1 u0_u4_u5_U74 (.A2( u0_u4_u5_n107 ) , .A1( u0_u4_u5_n109 ) , .ZN( u0_u4_u5_n120 ) );
  NAND2_X1 u0_u4_u5_U75 (.A2( u0_u4_u5_n100 ) , .A1( u0_u4_u5_n109 ) , .ZN( u0_u4_u5_n157 ) );
  AND2_X1 u0_u4_u5_U76 (.A2( u0_u4_u5_n100 ) , .A1( u0_u4_u5_n104 ) , .ZN( u0_u4_u5_n131 ) );
  NOR2_X1 u0_u4_u5_U77 (.A2( u0_u4_X_34 ) , .A1( u0_u4_X_35 ) , .ZN( u0_u4_u5_n145 ) );
  NOR2_X1 u0_u4_u5_U78 (.A2( u0_u4_X_34 ) , .ZN( u0_u4_u5_n146 ) , .A1( u0_u4_u5_n171 ) );
  NOR2_X1 u0_u4_u5_U79 (.A2( u0_u4_X_31 ) , .A1( u0_u4_X_32 ) , .ZN( u0_u4_u5_n103 ) );
  OAI22_X1 u0_u4_u5_U8 (.B2( u0_u4_u5_n149 ) , .B1( u0_u4_u5_n150 ) , .A2( u0_u4_u5_n151 ) , .A1( u0_u4_u5_n152 ) , .ZN( u0_u4_u5_n165 ) );
  NOR2_X1 u0_u4_u5_U80 (.A2( u0_u4_X_36 ) , .ZN( u0_u4_u5_n105 ) , .A1( u0_u4_u5_n180 ) );
  NOR2_X1 u0_u4_u5_U81 (.A2( u0_u4_X_33 ) , .ZN( u0_u4_u5_n108 ) , .A1( u0_u4_u5_n170 ) );
  NOR2_X1 u0_u4_u5_U82 (.A2( u0_u4_X_33 ) , .A1( u0_u4_X_36 ) , .ZN( u0_u4_u5_n107 ) );
  NOR2_X1 u0_u4_u5_U83 (.A2( u0_u4_X_31 ) , .ZN( u0_u4_u5_n104 ) , .A1( u0_u4_u5_n181 ) );
  NAND2_X1 u0_u4_u5_U84 (.A2( u0_u4_X_34 ) , .A1( u0_u4_X_35 ) , .ZN( u0_u4_u5_n153 ) );
  NAND2_X1 u0_u4_u5_U85 (.A1( u0_u4_X_34 ) , .ZN( u0_u4_u5_n126 ) , .A2( u0_u4_u5_n171 ) );
  AND2_X1 u0_u4_u5_U86 (.A1( u0_u4_X_31 ) , .A2( u0_u4_X_32 ) , .ZN( u0_u4_u5_n106 ) );
  AND2_X1 u0_u4_u5_U87 (.A1( u0_u4_X_31 ) , .ZN( u0_u4_u5_n109 ) , .A2( u0_u4_u5_n181 ) );
  INV_X1 u0_u4_u5_U88 (.A( u0_u4_X_33 ) , .ZN( u0_u4_u5_n180 ) );
  INV_X1 u0_u4_u5_U89 (.A( u0_u4_X_35 ) , .ZN( u0_u4_u5_n171 ) );
  NOR3_X1 u0_u4_u5_U9 (.A2( u0_u4_u5_n147 ) , .A1( u0_u4_u5_n148 ) , .ZN( u0_u4_u5_n149 ) , .A3( u0_u4_u5_n194 ) );
  INV_X1 u0_u4_u5_U90 (.A( u0_u4_X_36 ) , .ZN( u0_u4_u5_n170 ) );
  INV_X1 u0_u4_u5_U91 (.A( u0_u4_X_32 ) , .ZN( u0_u4_u5_n181 ) );
  NAND4_X1 u0_u4_u5_U92 (.ZN( u0_out4_29 ) , .A4( u0_u4_u5_n129 ) , .A3( u0_u4_u5_n130 ) , .A2( u0_u4_u5_n168 ) , .A1( u0_u4_u5_n196 ) );
  AOI221_X1 u0_u4_u5_U93 (.A( u0_u4_u5_n128 ) , .ZN( u0_u4_u5_n129 ) , .C2( u0_u4_u5_n132 ) , .B2( u0_u4_u5_n159 ) , .B1( u0_u4_u5_n176 ) , .C1( u0_u4_u5_n184 ) );
  AOI222_X1 u0_u4_u5_U94 (.ZN( u0_u4_u5_n130 ) , .A2( u0_u4_u5_n146 ) , .B1( u0_u4_u5_n147 ) , .C2( u0_u4_u5_n175 ) , .B2( u0_u4_u5_n179 ) , .A1( u0_u4_u5_n188 ) , .C1( u0_u4_u5_n194 ) );
  NAND4_X1 u0_u4_u5_U95 (.ZN( u0_out4_19 ) , .A4( u0_u4_u5_n166 ) , .A3( u0_u4_u5_n167 ) , .A2( u0_u4_u5_n168 ) , .A1( u0_u4_u5_n169 ) );
  AOI22_X1 u0_u4_u5_U96 (.B2( u0_u4_u5_n145 ) , .A2( u0_u4_u5_n146 ) , .ZN( u0_u4_u5_n167 ) , .B1( u0_u4_u5_n182 ) , .A1( u0_u4_u5_n189 ) );
  NOR4_X1 u0_u4_u5_U97 (.A4( u0_u4_u5_n162 ) , .A3( u0_u4_u5_n163 ) , .A2( u0_u4_u5_n164 ) , .A1( u0_u4_u5_n165 ) , .ZN( u0_u4_u5_n166 ) );
  NAND4_X1 u0_u4_u5_U98 (.ZN( u0_out4_11 ) , .A4( u0_u4_u5_n143 ) , .A3( u0_u4_u5_n144 ) , .A2( u0_u4_u5_n169 ) , .A1( u0_u4_u5_n196 ) );
  AOI22_X1 u0_u4_u5_U99 (.A2( u0_u4_u5_n132 ) , .ZN( u0_u4_u5_n144 ) , .B2( u0_u4_u5_n145 ) , .B1( u0_u4_u5_n184 ) , .A1( u0_u4_u5_n194 ) );
  AOI22_X1 u0_u4_u6_U10 (.A2( u0_u4_u6_n151 ) , .B2( u0_u4_u6_n161 ) , .A1( u0_u4_u6_n167 ) , .B1( u0_u4_u6_n170 ) , .ZN( u0_u4_u6_n89 ) );
  AOI21_X1 u0_u4_u6_U11 (.B1( u0_u4_u6_n107 ) , .B2( u0_u4_u6_n132 ) , .A( u0_u4_u6_n158 ) , .ZN( u0_u4_u6_n88 ) );
  AOI21_X1 u0_u4_u6_U12 (.B2( u0_u4_u6_n147 ) , .B1( u0_u4_u6_n148 ) , .ZN( u0_u4_u6_n149 ) , .A( u0_u4_u6_n158 ) );
  AOI21_X1 u0_u4_u6_U13 (.ZN( u0_u4_u6_n106 ) , .A( u0_u4_u6_n142 ) , .B2( u0_u4_u6_n159 ) , .B1( u0_u4_u6_n164 ) );
  INV_X1 u0_u4_u6_U14 (.A( u0_u4_u6_n155 ) , .ZN( u0_u4_u6_n161 ) );
  INV_X1 u0_u4_u6_U15 (.A( u0_u4_u6_n128 ) , .ZN( u0_u4_u6_n164 ) );
  NAND2_X1 u0_u4_u6_U16 (.ZN( u0_u4_u6_n110 ) , .A1( u0_u4_u6_n122 ) , .A2( u0_u4_u6_n129 ) );
  NAND2_X1 u0_u4_u6_U17 (.ZN( u0_u4_u6_n124 ) , .A2( u0_u4_u6_n146 ) , .A1( u0_u4_u6_n148 ) );
  INV_X1 u0_u4_u6_U18 (.A( u0_u4_u6_n132 ) , .ZN( u0_u4_u6_n171 ) );
  AND2_X1 u0_u4_u6_U19 (.A1( u0_u4_u6_n100 ) , .ZN( u0_u4_u6_n130 ) , .A2( u0_u4_u6_n147 ) );
  INV_X1 u0_u4_u6_U20 (.A( u0_u4_u6_n127 ) , .ZN( u0_u4_u6_n173 ) );
  INV_X1 u0_u4_u6_U21 (.A( u0_u4_u6_n121 ) , .ZN( u0_u4_u6_n167 ) );
  INV_X1 u0_u4_u6_U22 (.A( u0_u4_u6_n100 ) , .ZN( u0_u4_u6_n169 ) );
  INV_X1 u0_u4_u6_U23 (.A( u0_u4_u6_n123 ) , .ZN( u0_u4_u6_n170 ) );
  INV_X1 u0_u4_u6_U24 (.A( u0_u4_u6_n113 ) , .ZN( u0_u4_u6_n168 ) );
  AND2_X1 u0_u4_u6_U25 (.A1( u0_u4_u6_n107 ) , .A2( u0_u4_u6_n119 ) , .ZN( u0_u4_u6_n133 ) );
  AND2_X1 u0_u4_u6_U26 (.A2( u0_u4_u6_n121 ) , .A1( u0_u4_u6_n122 ) , .ZN( u0_u4_u6_n131 ) );
  AND3_X1 u0_u4_u6_U27 (.ZN( u0_u4_u6_n120 ) , .A2( u0_u4_u6_n127 ) , .A1( u0_u4_u6_n132 ) , .A3( u0_u4_u6_n145 ) );
  INV_X1 u0_u4_u6_U28 (.A( u0_u4_u6_n146 ) , .ZN( u0_u4_u6_n163 ) );
  AOI222_X1 u0_u4_u6_U29 (.ZN( u0_u4_u6_n114 ) , .A1( u0_u4_u6_n118 ) , .A2( u0_u4_u6_n126 ) , .B2( u0_u4_u6_n151 ) , .C2( u0_u4_u6_n159 ) , .C1( u0_u4_u6_n168 ) , .B1( u0_u4_u6_n169 ) );
  INV_X1 u0_u4_u6_U3 (.A( u0_u4_u6_n110 ) , .ZN( u0_u4_u6_n166 ) );
  NOR2_X1 u0_u4_u6_U30 (.A1( u0_u4_u6_n162 ) , .A2( u0_u4_u6_n165 ) , .ZN( u0_u4_u6_n98 ) );
  NAND2_X1 u0_u4_u6_U31 (.A1( u0_u4_u6_n144 ) , .ZN( u0_u4_u6_n151 ) , .A2( u0_u4_u6_n158 ) );
  NAND2_X1 u0_u4_u6_U32 (.ZN( u0_u4_u6_n132 ) , .A1( u0_u4_u6_n91 ) , .A2( u0_u4_u6_n97 ) );
  AOI22_X1 u0_u4_u6_U33 (.B2( u0_u4_u6_n110 ) , .B1( u0_u4_u6_n111 ) , .A1( u0_u4_u6_n112 ) , .ZN( u0_u4_u6_n115 ) , .A2( u0_u4_u6_n161 ) );
  NAND4_X1 u0_u4_u6_U34 (.A3( u0_u4_u6_n109 ) , .ZN( u0_u4_u6_n112 ) , .A4( u0_u4_u6_n132 ) , .A2( u0_u4_u6_n147 ) , .A1( u0_u4_u6_n166 ) );
  NOR2_X1 u0_u4_u6_U35 (.ZN( u0_u4_u6_n109 ) , .A1( u0_u4_u6_n170 ) , .A2( u0_u4_u6_n173 ) );
  NOR2_X1 u0_u4_u6_U36 (.A2( u0_u4_u6_n126 ) , .ZN( u0_u4_u6_n155 ) , .A1( u0_u4_u6_n160 ) );
  NAND2_X1 u0_u4_u6_U37 (.ZN( u0_u4_u6_n146 ) , .A2( u0_u4_u6_n94 ) , .A1( u0_u4_u6_n99 ) );
  AOI21_X1 u0_u4_u6_U38 (.A( u0_u4_u6_n144 ) , .B2( u0_u4_u6_n145 ) , .B1( u0_u4_u6_n146 ) , .ZN( u0_u4_u6_n150 ) );
  AOI211_X1 u0_u4_u6_U39 (.B( u0_u4_u6_n134 ) , .A( u0_u4_u6_n135 ) , .C1( u0_u4_u6_n136 ) , .ZN( u0_u4_u6_n137 ) , .C2( u0_u4_u6_n151 ) );
  INV_X1 u0_u4_u6_U4 (.A( u0_u4_u6_n142 ) , .ZN( u0_u4_u6_n174 ) );
  NAND4_X1 u0_u4_u6_U40 (.A4( u0_u4_u6_n127 ) , .A3( u0_u4_u6_n128 ) , .A2( u0_u4_u6_n129 ) , .A1( u0_u4_u6_n130 ) , .ZN( u0_u4_u6_n136 ) );
  AOI21_X1 u0_u4_u6_U41 (.B2( u0_u4_u6_n132 ) , .B1( u0_u4_u6_n133 ) , .ZN( u0_u4_u6_n134 ) , .A( u0_u4_u6_n158 ) );
  AOI21_X1 u0_u4_u6_U42 (.B1( u0_u4_u6_n131 ) , .ZN( u0_u4_u6_n135 ) , .A( u0_u4_u6_n144 ) , .B2( u0_u4_u6_n146 ) );
  INV_X1 u0_u4_u6_U43 (.A( u0_u4_u6_n111 ) , .ZN( u0_u4_u6_n158 ) );
  NAND2_X1 u0_u4_u6_U44 (.ZN( u0_u4_u6_n127 ) , .A1( u0_u4_u6_n91 ) , .A2( u0_u4_u6_n92 ) );
  NAND2_X1 u0_u4_u6_U45 (.ZN( u0_u4_u6_n129 ) , .A2( u0_u4_u6_n95 ) , .A1( u0_u4_u6_n96 ) );
  INV_X1 u0_u4_u6_U46 (.A( u0_u4_u6_n144 ) , .ZN( u0_u4_u6_n159 ) );
  NAND2_X1 u0_u4_u6_U47 (.ZN( u0_u4_u6_n145 ) , .A2( u0_u4_u6_n97 ) , .A1( u0_u4_u6_n98 ) );
  NAND2_X1 u0_u4_u6_U48 (.ZN( u0_u4_u6_n148 ) , .A2( u0_u4_u6_n92 ) , .A1( u0_u4_u6_n94 ) );
  NAND2_X1 u0_u4_u6_U49 (.ZN( u0_u4_u6_n108 ) , .A2( u0_u4_u6_n139 ) , .A1( u0_u4_u6_n144 ) );
  NAND2_X1 u0_u4_u6_U5 (.A2( u0_u4_u6_n143 ) , .ZN( u0_u4_u6_n152 ) , .A1( u0_u4_u6_n166 ) );
  NAND2_X1 u0_u4_u6_U50 (.ZN( u0_u4_u6_n121 ) , .A2( u0_u4_u6_n95 ) , .A1( u0_u4_u6_n97 ) );
  NAND2_X1 u0_u4_u6_U51 (.ZN( u0_u4_u6_n107 ) , .A2( u0_u4_u6_n92 ) , .A1( u0_u4_u6_n95 ) );
  AND2_X1 u0_u4_u6_U52 (.ZN( u0_u4_u6_n118 ) , .A2( u0_u4_u6_n91 ) , .A1( u0_u4_u6_n99 ) );
  NAND2_X1 u0_u4_u6_U53 (.ZN( u0_u4_u6_n147 ) , .A2( u0_u4_u6_n98 ) , .A1( u0_u4_u6_n99 ) );
  NAND2_X1 u0_u4_u6_U54 (.ZN( u0_u4_u6_n128 ) , .A1( u0_u4_u6_n94 ) , .A2( u0_u4_u6_n96 ) );
  NAND2_X1 u0_u4_u6_U55 (.ZN( u0_u4_u6_n119 ) , .A2( u0_u4_u6_n95 ) , .A1( u0_u4_u6_n99 ) );
  NAND2_X1 u0_u4_u6_U56 (.ZN( u0_u4_u6_n123 ) , .A2( u0_u4_u6_n91 ) , .A1( u0_u4_u6_n96 ) );
  NAND2_X1 u0_u4_u6_U57 (.ZN( u0_u4_u6_n100 ) , .A2( u0_u4_u6_n92 ) , .A1( u0_u4_u6_n98 ) );
  NAND2_X1 u0_u4_u6_U58 (.ZN( u0_u4_u6_n122 ) , .A1( u0_u4_u6_n94 ) , .A2( u0_u4_u6_n97 ) );
  INV_X1 u0_u4_u6_U59 (.A( u0_u4_u6_n139 ) , .ZN( u0_u4_u6_n160 ) );
  AOI22_X1 u0_u4_u6_U6 (.B2( u0_u4_u6_n101 ) , .A1( u0_u4_u6_n102 ) , .ZN( u0_u4_u6_n103 ) , .B1( u0_u4_u6_n160 ) , .A2( u0_u4_u6_n161 ) );
  NAND2_X1 u0_u4_u6_U60 (.ZN( u0_u4_u6_n113 ) , .A1( u0_u4_u6_n96 ) , .A2( u0_u4_u6_n98 ) );
  NOR2_X1 u0_u4_u6_U61 (.A2( u0_u4_X_40 ) , .A1( u0_u4_X_41 ) , .ZN( u0_u4_u6_n126 ) );
  NOR2_X1 u0_u4_u6_U62 (.A2( u0_u4_X_39 ) , .A1( u0_u4_X_42 ) , .ZN( u0_u4_u6_n92 ) );
  NOR2_X1 u0_u4_u6_U63 (.A2( u0_u4_X_39 ) , .A1( u0_u4_u6_n156 ) , .ZN( u0_u4_u6_n97 ) );
  NOR2_X1 u0_u4_u6_U64 (.A2( u0_u4_X_38 ) , .A1( u0_u4_u6_n165 ) , .ZN( u0_u4_u6_n95 ) );
  NOR2_X1 u0_u4_u6_U65 (.A2( u0_u4_X_41 ) , .ZN( u0_u4_u6_n111 ) , .A1( u0_u4_u6_n157 ) );
  NOR2_X1 u0_u4_u6_U66 (.A2( u0_u4_X_37 ) , .A1( u0_u4_u6_n162 ) , .ZN( u0_u4_u6_n94 ) );
  NOR2_X1 u0_u4_u6_U67 (.A2( u0_u4_X_37 ) , .A1( u0_u4_X_38 ) , .ZN( u0_u4_u6_n91 ) );
  NAND2_X1 u0_u4_u6_U68 (.A1( u0_u4_X_41 ) , .ZN( u0_u4_u6_n144 ) , .A2( u0_u4_u6_n157 ) );
  NAND2_X1 u0_u4_u6_U69 (.A2( u0_u4_X_40 ) , .A1( u0_u4_X_41 ) , .ZN( u0_u4_u6_n139 ) );
  NOR2_X1 u0_u4_u6_U7 (.A1( u0_u4_u6_n118 ) , .ZN( u0_u4_u6_n143 ) , .A2( u0_u4_u6_n168 ) );
  AND2_X1 u0_u4_u6_U70 (.A1( u0_u4_X_39 ) , .A2( u0_u4_u6_n156 ) , .ZN( u0_u4_u6_n96 ) );
  AND2_X1 u0_u4_u6_U71 (.A1( u0_u4_X_39 ) , .A2( u0_u4_X_42 ) , .ZN( u0_u4_u6_n99 ) );
  INV_X1 u0_u4_u6_U72 (.A( u0_u4_X_40 ) , .ZN( u0_u4_u6_n157 ) );
  INV_X1 u0_u4_u6_U73 (.A( u0_u4_X_37 ) , .ZN( u0_u4_u6_n165 ) );
  INV_X1 u0_u4_u6_U74 (.A( u0_u4_X_38 ) , .ZN( u0_u4_u6_n162 ) );
  INV_X1 u0_u4_u6_U75 (.A( u0_u4_X_42 ) , .ZN( u0_u4_u6_n156 ) );
  NAND4_X1 u0_u4_u6_U76 (.ZN( u0_out4_32 ) , .A4( u0_u4_u6_n103 ) , .A3( u0_u4_u6_n104 ) , .A2( u0_u4_u6_n105 ) , .A1( u0_u4_u6_n106 ) );
  AOI22_X1 u0_u4_u6_U77 (.ZN( u0_u4_u6_n105 ) , .A2( u0_u4_u6_n108 ) , .A1( u0_u4_u6_n118 ) , .B2( u0_u4_u6_n126 ) , .B1( u0_u4_u6_n171 ) );
  AOI22_X1 u0_u4_u6_U78 (.ZN( u0_u4_u6_n104 ) , .A1( u0_u4_u6_n111 ) , .B1( u0_u4_u6_n124 ) , .B2( u0_u4_u6_n151 ) , .A2( u0_u4_u6_n93 ) );
  NAND4_X1 u0_u4_u6_U79 (.ZN( u0_out4_12 ) , .A4( u0_u4_u6_n114 ) , .A3( u0_u4_u6_n115 ) , .A2( u0_u4_u6_n116 ) , .A1( u0_u4_u6_n117 ) );
  INV_X1 u0_u4_u6_U8 (.ZN( u0_u4_u6_n172 ) , .A( u0_u4_u6_n88 ) );
  OAI22_X1 u0_u4_u6_U80 (.B2( u0_u4_u6_n111 ) , .ZN( u0_u4_u6_n116 ) , .B1( u0_u4_u6_n126 ) , .A2( u0_u4_u6_n164 ) , .A1( u0_u4_u6_n167 ) );
  OAI21_X1 u0_u4_u6_U81 (.A( u0_u4_u6_n108 ) , .ZN( u0_u4_u6_n117 ) , .B2( u0_u4_u6_n141 ) , .B1( u0_u4_u6_n163 ) );
  OAI211_X1 u0_u4_u6_U82 (.ZN( u0_out4_22 ) , .B( u0_u4_u6_n137 ) , .A( u0_u4_u6_n138 ) , .C2( u0_u4_u6_n139 ) , .C1( u0_u4_u6_n140 ) );
  AOI22_X1 u0_u4_u6_U83 (.B1( u0_u4_u6_n124 ) , .A2( u0_u4_u6_n125 ) , .A1( u0_u4_u6_n126 ) , .ZN( u0_u4_u6_n138 ) , .B2( u0_u4_u6_n161 ) );
  AND4_X1 u0_u4_u6_U84 (.A3( u0_u4_u6_n119 ) , .A1( u0_u4_u6_n120 ) , .A4( u0_u4_u6_n129 ) , .ZN( u0_u4_u6_n140 ) , .A2( u0_u4_u6_n143 ) );
  OAI211_X1 u0_u4_u6_U85 (.ZN( u0_out4_7 ) , .B( u0_u4_u6_n153 ) , .C2( u0_u4_u6_n154 ) , .C1( u0_u4_u6_n155 ) , .A( u0_u4_u6_n174 ) );
  NOR3_X1 u0_u4_u6_U86 (.A1( u0_u4_u6_n141 ) , .ZN( u0_u4_u6_n154 ) , .A3( u0_u4_u6_n164 ) , .A2( u0_u4_u6_n171 ) );
  AOI211_X1 u0_u4_u6_U87 (.B( u0_u4_u6_n149 ) , .A( u0_u4_u6_n150 ) , .C2( u0_u4_u6_n151 ) , .C1( u0_u4_u6_n152 ) , .ZN( u0_u4_u6_n153 ) );
  NAND3_X1 u0_u4_u6_U88 (.A2( u0_u4_u6_n123 ) , .ZN( u0_u4_u6_n125 ) , .A1( u0_u4_u6_n130 ) , .A3( u0_u4_u6_n131 ) );
  NAND3_X1 u0_u4_u6_U89 (.A3( u0_u4_u6_n133 ) , .ZN( u0_u4_u6_n141 ) , .A1( u0_u4_u6_n145 ) , .A2( u0_u4_u6_n148 ) );
  OAI21_X1 u0_u4_u6_U9 (.A( u0_u4_u6_n159 ) , .B1( u0_u4_u6_n169 ) , .B2( u0_u4_u6_n173 ) , .ZN( u0_u4_u6_n90 ) );
  NAND3_X1 u0_u4_u6_U90 (.ZN( u0_u4_u6_n101 ) , .A3( u0_u4_u6_n107 ) , .A2( u0_u4_u6_n121 ) , .A1( u0_u4_u6_n127 ) );
  NAND3_X1 u0_u4_u6_U91 (.ZN( u0_u4_u6_n102 ) , .A3( u0_u4_u6_n130 ) , .A2( u0_u4_u6_n145 ) , .A1( u0_u4_u6_n166 ) );
  NAND3_X1 u0_u4_u6_U92 (.A3( u0_u4_u6_n113 ) , .A1( u0_u4_u6_n119 ) , .A2( u0_u4_u6_n123 ) , .ZN( u0_u4_u6_n93 ) );
  NAND3_X1 u0_u4_u6_U93 (.ZN( u0_u4_u6_n142 ) , .A2( u0_u4_u6_n172 ) , .A3( u0_u4_u6_n89 ) , .A1( u0_u4_u6_n90 ) );
  OAI22_X1 u0_uk_U100 (.ZN( u0_K12_5 ) , .B2( u0_uk_n150 ) , .A2( u0_uk_n176 ) , .A1( u0_uk_n209 ) , .B1( u0_uk_n83 ) );
  NAND2_X1 u0_uk_U1005 (.A1( u0_uk_K_r1_10 ) , .A2( u0_uk_n100 ) , .ZN( u0_uk_n841 ) );
  OAI21_X1 u0_uk_U1014 (.ZN( u0_K1_37 ) , .B1( u0_uk_n129 ) , .B2( u0_uk_n714 ) , .A( u0_uk_n876 ) );
  NAND2_X1 u0_uk_U1015 (.A1( u0_key_r_50 ) , .A2( u0_uk_n17 ) , .ZN( u0_uk_n876 ) );
  INV_X1 u0_uk_U1062 (.A( u0_key_r_9 ) , .ZN( u0_uk_n709 ) );
  INV_X1 u0_uk_U1063 (.A( u0_key_r_7 ) , .ZN( u0_uk_n711 ) );
  INV_X1 u0_uk_U1067 (.A( u0_key_r_23 ) , .ZN( u0_uk_n700 ) );
  INV_X1 u0_uk_U1069 (.A( u0_key_r_30 ) , .ZN( u0_uk_n693 ) );
  INV_X1 u0_uk_U1074 (.A( u0_key_r_37 ) , .ZN( u0_uk_n687 ) );
  INV_X1 u0_uk_U1075 (.A( u0_key_r_52 ) , .ZN( u0_uk_n675 ) );
  INV_X1 u0_uk_U1076 (.A( u0_key_r_0 ) , .ZN( u0_uk_n716 ) );
  INV_X1 u0_uk_U1077 (.A( u0_key_r_16 ) , .ZN( u0_uk_n706 ) );
  INV_X1 u0_uk_U1079 (.A( u0_key_r_1 ) , .ZN( u0_uk_n715 ) );
  INV_X1 u0_uk_U1080 (.A( u0_key_r_2 ) , .ZN( u0_uk_n714 ) );
  OAI21_X1 u0_uk_U1089 (.ZN( u0_K16_14 ) , .B1( u0_uk_n252 ) , .B2( u0_uk_n653 ) , .A( u0_uk_n908 ) );
  NAND2_X1 u0_uk_U1090 (.A1( u0_uk_K_r14_18 ) , .A2( u0_uk_n207 ) , .ZN( u0_uk_n908 ) );
  OAI21_X1 u0_uk_U1097 (.ZN( u0_K5_39 ) , .B1( u0_uk_n208 ) , .B2( u0_uk_n482 ) , .A( u0_uk_n808 ) );
  NAND2_X1 u0_uk_U1098 (.A1( u0_uk_K_r3_16 ) , .A2( u0_uk_n208 ) , .ZN( u0_uk_n808 ) );
  INV_X1 u0_uk_U1107 (.ZN( u0_K1_41 ) , .A( u0_uk_n874 ) );
  AOI22_X1 u0_uk_U1108 (.B2( u0_key_r_35 ) , .A2( u0_key_r_42 ) , .B1( u0_uk_n145 ) , .A1( u0_uk_n251 ) , .ZN( u0_uk_n874 ) );
  INV_X1 u0_uk_U1117 (.ZN( u0_K12_4 ) , .A( u0_uk_n963 ) );
  OAI22_X1 u0_uk_U112 (.ZN( u0_K16_47 ) , .B1( u0_uk_n128 ) , .A1( u0_uk_n187 ) , .A2( u0_uk_n666 ) , .B2( u0_uk_n670 ) );
  INV_X1 u0_uk_U1125 (.ZN( u0_K1_32 ) , .A( u0_uk_n879 ) );
  AOI22_X1 u0_uk_U1126 (.B2( u0_key_r_22 ) , .A2( u0_key_r_29 ) , .B1( u0_uk_n146 ) , .A1( u0_uk_n242 ) , .ZN( u0_uk_n879 ) );
  INV_X1 u0_uk_U1147 (.ZN( u0_K5_35 ) , .A( u0_uk_n810 ) );
  AOI22_X1 u0_uk_U1160 (.B2( u0_uk_K_r10_39 ) , .A2( u0_uk_K_r10_48 ) , .B1( u0_uk_n11 ) , .A1( u0_uk_n213 ) , .ZN( u0_uk_n978 ) );
  INV_X1 u0_uk_U1161 (.ZN( u0_K12_1 ) , .A( u0_uk_n978 ) );
  INV_X1 u0_uk_U12 (.A( u0_uk_n187 ) , .ZN( u0_uk_n92 ) );
  INV_X1 u0_uk_U133 (.ZN( u0_K12_15 ) , .A( u0_uk_n980 ) );
  AOI22_X1 u0_uk_U134 (.B2( u0_uk_K_r10_25 ) , .A2( u0_uk_K_r10_34 ) , .B1( u0_uk_n141 ) , .A1( u0_uk_n257 ) , .ZN( u0_uk_n980 ) );
  OAI22_X1 u0_uk_U145 (.ZN( u0_K16_15 ) , .B1( u0_uk_n17 ) , .A1( u0_uk_n187 ) , .A2( u0_uk_n645 ) , .B2( u0_uk_n652 ) );
  OAI22_X1 u0_uk_U164 (.ZN( u0_K5_30 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n222 ) , .A2( u0_uk_n463 ) , .B2( u0_uk_n480 ) );
  OAI22_X1 u0_uk_U178 (.ZN( u0_K12_14 ) , .A1( u0_uk_n100 ) , .A2( u0_uk_n165 ) , .B2( u0_uk_n170 ) , .B1( u0_uk_n202 ) );
  OAI22_X1 u0_uk_U179 (.ZN( u0_K12_24 ) , .A1( u0_uk_n102 ) , .A2( u0_uk_n143 ) , .B1( u0_uk_n163 ) , .B2( u0_uk_n172 ) );
  INV_X1 u0_uk_U213 (.A( u0_key_r_14 ) , .ZN( u0_uk_n707 ) );
  OAI21_X1 u0_uk_U231 (.ZN( u0_K1_39 ) , .B1( u0_uk_n118 ) , .B2( u0_uk_n701 ) , .A( u0_uk_n875 ) );
  INV_X1 u0_uk_U233 (.A( u0_key_r_22 ) , .ZN( u0_uk_n701 ) );
  OAI22_X1 u0_uk_U241 (.ZN( u0_K16_48 ) , .B1( u0_uk_n102 ) , .A1( u0_uk_n187 ) , .A2( u0_uk_n650 ) , .B2( u0_uk_n658 ) );
  OAI21_X1 u0_uk_U242 (.ZN( u0_K16_44 ) , .B1( u0_uk_n110 ) , .B2( u0_uk_n642 ) , .A( u0_uk_n895 ) );
  NAND2_X1 u0_uk_U243 (.A1( u0_uk_K_r14_43 ) , .ZN( u0_uk_n895 ) , .A2( u0_uk_n99 ) );
  INV_X1 u0_uk_U250 (.ZN( u0_K1_48 ) , .A( u0_uk_n870 ) );
  AOI22_X1 u0_uk_U251 (.B2( u0_key_r_21 ) , .A2( u0_key_r_28 ) , .B1( u0_uk_n145 ) , .A1( u0_uk_n213 ) , .ZN( u0_uk_n870 ) );
  INV_X1 u0_uk_U252 (.ZN( u0_K1_44 ) , .A( u0_uk_n872 ) );
  AOI22_X1 u0_uk_U253 (.B2( u0_key_r_36 ) , .A2( u0_key_r_43 ) , .B1( u0_uk_n145 ) , .A1( u0_uk_n223 ) , .ZN( u0_uk_n872 ) );
  OAI22_X1 u0_uk_U286 (.ZN( u0_K12_8 ) , .A2( u0_uk_n136 ) , .B2( u0_uk_n157 ) , .A1( u0_uk_n191 ) , .B1( u0_uk_n83 ) );
  INV_X1 u0_uk_U297 (.ZN( u0_K1_26 ) , .A( u0_uk_n883 ) );
  AOI22_X1 u0_uk_U298 (.B2( u0_key_r_31 ) , .A2( u0_key_r_51 ) , .A1( u0_uk_n146 ) , .B1( u0_uk_n207 ) , .ZN( u0_uk_n883 ) );
  OAI22_X1 u0_uk_U357 (.ZN( u0_K1_40 ) , .A1( u0_uk_n230 ) , .A2( u0_uk_n675 ) , .B2( u0_uk_n716 ) , .B1( u0_uk_n99 ) );
  OAI22_X1 u0_uk_U371 (.ZN( u0_K1_28 ) , .A1( u0_uk_n118 ) , .B1( u0_uk_n220 ) , .A2( u0_uk_n710 ) , .B2( u0_uk_n715 ) );
  INV_X1 u0_uk_U372 (.A( u0_key_r_8 ) , .ZN( u0_uk_n710 ) );
  OAI21_X1 u0_uk_U379 (.ZN( u0_K5_33 ) , .B1( u0_uk_n250 ) , .B2( u0_uk_n457 ) , .A( u0_uk_n811 ) );
  NAND2_X1 u0_uk_U380 (.A1( u0_uk_K_r3_14 ) , .A2( u0_uk_n220 ) , .ZN( u0_uk_n811 ) );
  INV_X1 u0_uk_U426 (.ZN( u0_K1_33 ) , .A( u0_uk_n878 ) );
  OAI22_X1 u0_uk_U430 (.ZN( u0_K16_16 ) , .B1( u0_uk_n17 ) , .A1( u0_uk_n187 ) , .A2( u0_uk_n644 ) , .B2( u0_uk_n651 ) );
  NAND2_X1 u0_uk_U458 (.A1( u0_uk_K_r9_38 ) , .A2( u0_uk_n128 ) , .ZN( u0_uk_n989 ) );
  OAI22_X1 u0_uk_U467 (.ZN( u0_K5_37 ) , .A1( u0_uk_n100 ) , .B1( u0_uk_n222 ) , .A2( u0_uk_n455 ) , .B2( u0_uk_n493 ) );
  OAI22_X1 u0_uk_U469 (.ZN( u0_K1_29 ) , .A1( u0_uk_n142 ) , .B1( u0_uk_n188 ) , .A2( u0_uk_n700 ) , .B2( u0_uk_n706 ) );
  OAI22_X1 u0_uk_U487 (.ZN( u0_K5_29 ) , .A1( u0_uk_n118 ) , .B1( u0_uk_n222 ) , .A2( u0_uk_n462 ) , .B2( u0_uk_n481 ) );
  OAI22_X1 u0_uk_U489 (.ZN( u0_K12_2 ) , .A1( u0_uk_n148 ) , .B2( u0_uk_n172 ) , .A2( u0_uk_n177 ) , .B1( u0_uk_n92 ) );
  OAI21_X1 u0_uk_U520 (.ZN( u0_K12_12 ) , .B1( u0_uk_n109 ) , .B2( u0_uk_n169 ) , .A( u0_uk_n981 ) );
  BUF_X1 u0_uk_U53 (.A( u0_uk_n163 ) , .Z( u0_uk_n208 ) );
  OAI22_X1 u0_uk_U531 (.ZN( u0_K1_36 ) , .A1( u0_uk_n128 ) , .B1( u0_uk_n188 ) , .A2( u0_uk_n693 ) , .B2( u0_uk_n700 ) );
  OAI21_X1 u0_uk_U534 (.ZN( u0_K16_17 ) , .B1( u0_uk_n252 ) , .B2( u0_uk_n661 ) , .A( u0_uk_n907 ) );
  NAND2_X1 u0_uk_U535 (.A1( u0_uk_K_r14_10 ) , .A2( u0_uk_n202 ) , .ZN( u0_uk_n907 ) );
  INV_X1 u0_uk_U540 (.ZN( u0_K12_17 ) , .A( u0_uk_n979 ) );
  AOI22_X1 u0_uk_U541 (.B2( u0_uk_K_r10_18 ) , .A2( u0_uk_K_r10_41 ) , .A1( u0_uk_n129 ) , .B1( u0_uk_n207 ) , .ZN( u0_uk_n979 ) );
  OAI22_X1 u0_uk_U549 (.ZN( u0_K1_38 ) , .A1( u0_uk_n118 ) , .B1( u0_uk_n188 ) , .A2( u0_uk_n687 ) , .B2( u0_uk_n693 ) );
  INV_X1 u0_uk_U550 (.ZN( u0_K5_36 ) , .A( u0_uk_n809 ) );
  AOI22_X1 u0_uk_U551 (.B2( u0_uk_K_r3_29 ) , .A2( u0_uk_K_r3_52 ) , .B1( u0_uk_n141 ) , .A1( u0_uk_n223 ) , .ZN( u0_uk_n809 ) );
  INV_X1 u0_uk_U620 (.ZN( u0_K1_35 ) , .A( u0_uk_n877 ) );
  AOI22_X1 u0_uk_U621 (.B2( u0_key_r_28 ) , .A2( u0_key_r_35 ) , .B1( u0_uk_n146 ) , .A1( u0_uk_n161 ) , .ZN( u0_uk_n877 ) );
  INV_X1 u0_uk_U641 (.ZN( u0_K12_23 ) , .A( u0_uk_n975 ) );
  AOI22_X1 u0_uk_U642 (.B2( u0_uk_K_r10_32 ) , .A2( u0_uk_K_r10_41 ) , .A1( u0_uk_n220 ) , .B1( u0_uk_n83 ) , .ZN( u0_uk_n975 ) );
  OAI21_X1 u0_uk_U645 (.ZN( u0_K12_6 ) , .B1( u0_uk_n147 ) , .B2( u0_uk_n156 ) , .A( u0_uk_n962 ) );
  NAND2_X1 u0_uk_U646 (.A1( u0_uk_K_r10_10 ) , .A2( u0_uk_n163 ) , .ZN( u0_uk_n962 ) );
  OAI22_X1 u0_uk_U647 (.ZN( u0_K16_45 ) , .B1( u0_uk_n110 ) , .A1( u0_uk_n155 ) , .A2( u0_uk_n638 ) , .B2( u0_uk_n641 ) );
  INV_X1 u0_uk_U658 (.ZN( u0_K16_43 ) , .A( u0_uk_n896 ) );
  AOI22_X1 u0_uk_U659 (.B2( u0_uk_K_r14_16 ) , .A2( u0_uk_K_r14_9 ) , .B1( u0_uk_n142 ) , .A1( u0_uk_n191 ) , .ZN( u0_uk_n896 ) );
  NAND2_X1 u0_uk_U676 (.A1( u0_uk_K_r2_29 ) , .A2( u0_uk_n100 ) , .ZN( u0_uk_n823 ) );
  OAI21_X1 u0_uk_U690 (.ZN( u0_K5_25 ) , .B1( u0_uk_n129 ) , .B2( u0_uk_n475 ) , .A( u0_uk_n814 ) );
  NAND2_X1 u0_uk_U691 (.A1( u0_uk_K_r3_35 ) , .A2( u0_uk_n128 ) , .ZN( u0_uk_n814 ) );
  INV_X1 u0_uk_U710 (.ZN( u0_K1_25 ) , .A( u0_uk_n884 ) );
  AOI22_X1 u0_uk_U711 (.B2( u0_key_r_29 ) , .A2( u0_key_r_36 ) , .B1( u0_uk_n146 ) , .A1( u0_uk_n242 ) , .ZN( u0_uk_n884 ) );
  OAI21_X1 u0_uk_U731 (.ZN( u0_K5_42 ) , .B1( u0_uk_n128 ) , .B2( u0_uk_n476 ) , .A( u0_uk_n807 ) );
  NAND2_X1 u0_uk_U732 (.A1( u0_uk_K_r3_9 ) , .ZN( u0_uk_n807 ) , .A2( u0_uk_n92 ) );
  OAI22_X1 u0_uk_U74 (.ZN( u0_K16_23 ) , .A1( u0_uk_n164 ) , .A2( u0_uk_n640 ) , .B2( u0_uk_n645 ) , .B1( u0_uk_n92 ) );
  INV_X1 u0_uk_U742 (.ZN( u0_K1_42 ) , .A( u0_uk_n873 ) );
  AOI22_X1 u0_uk_U743 (.B2( u0_key_r_31 ) , .A2( u0_key_r_38 ) , .B1( u0_uk_n145 ) , .A1( u0_uk_n251 ) , .ZN( u0_uk_n873 ) );
  OAI22_X1 u0_uk_U751 (.ZN( u0_K12_13 ) , .A1( u0_uk_n100 ) , .A2( u0_uk_n137 ) , .B2( u0_uk_n169 ) , .B1( u0_uk_n238 ) );
  INV_X1 u0_uk_U774 (.ZN( u0_K5_27 ) , .A( u0_uk_n813 ) );
  INV_X1 u0_uk_U784 (.ZN( u0_K12_21 ) , .A( u0_uk_n976 ) );
  AOI22_X1 u0_uk_U785 (.B2( u0_uk_K_r10_25 ) , .A2( u0_uk_K_r10_48 ) , .A1( u0_uk_n10 ) , .B1( u0_uk_n207 ) , .ZN( u0_uk_n976 ) );
  OAI21_X1 u0_uk_U788 (.ZN( u0_K16_13 ) , .B1( u0_uk_n147 ) , .B2( u0_uk_n631 ) , .A( u0_uk_n909 ) );
  NAND2_X1 u0_uk_U789 (.A1( u0_uk_K_r14_46 ) , .A2( u0_uk_n208 ) , .ZN( u0_uk_n909 ) );
  INV_X1 u0_uk_U794 (.ZN( u0_K1_27 ) , .A( u0_uk_n882 ) );
  AOI22_X1 u0_uk_U795 (.B2( u0_key_r_14 ) , .A2( u0_key_r_21 ) , .B1( u0_uk_n146 ) , .A1( u0_uk_n238 ) , .ZN( u0_uk_n882 ) );
  OAI21_X1 u0_uk_U810 (.ZN( u0_K12_20 ) , .B1( u0_uk_n129 ) , .B2( u0_uk_n166 ) , .A( u0_uk_n977 ) );
  NAND2_X1 u0_uk_U811 (.A1( u0_uk_K_r10_47 ) , .A2( u0_uk_n31 ) , .ZN( u0_uk_n977 ) );
  OAI22_X1 u0_uk_U822 (.ZN( u0_K16_20 ) , .A1( u0_uk_n155 ) , .B1( u0_uk_n17 ) , .A2( u0_uk_n629 ) , .B2( u0_uk_n636 ) );
  OAI22_X1 u0_uk_U843 (.ZN( u0_K1_43 ) , .B1( u0_uk_n109 ) , .A1( u0_uk_n164 ) , .B2( u0_uk_n706 ) , .A2( u0_uk_n709 ) );
  INV_X1 u0_uk_U844 (.ZN( u0_K12_3 ) , .A( u0_uk_n968 ) );
  AOI22_X1 u0_uk_U845 (.B2( u0_uk_K_r10_18 ) , .A2( u0_uk_K_r10_27 ) , .A1( u0_uk_n188 ) , .B1( u0_uk_n27 ) , .ZN( u0_uk_n968 ) );
  OAI22_X1 u0_uk_U881 (.ZN( u0_K12_10 ) , .B1( u0_uk_n142 ) , .A2( u0_uk_n149 ) , .B2( u0_uk_n170 ) , .A1( u0_uk_n191 ) );
  OAI22_X1 u0_uk_U882 (.ZN( u0_K12_11 ) , .B2( u0_uk_n149 ) , .A2( u0_uk_n175 ) , .A1( u0_uk_n182 ) , .B1( u0_uk_n93 ) );
  INV_X1 u0_uk_U9 (.A( u0_uk_n147 ) , .ZN( u0_uk_n17 ) );
  OAI22_X1 u0_uk_U908 (.ZN( u0_K16_21 ) , .A1( u0_uk_n187 ) , .A2( u0_uk_n654 ) , .B2( u0_uk_n661 ) , .B1( u0_uk_n94 ) );
  OAI22_X1 u0_uk_U932 (.ZN( u0_K12_16 ) , .A1( u0_uk_n100 ) , .B1( u0_uk_n163 ) , .B2( u0_uk_n165 ) , .A2( u0_uk_n177 ) );
  OAI22_X1 u0_uk_U939 (.ZN( u0_K12_18 ) , .A1( u0_uk_n100 ) , .B2( u0_uk_n137 ) , .B1( u0_uk_n163 ) , .A2( u0_uk_n175 ) );
  OAI22_X1 u0_uk_U945 (.ZN( u0_K16_46 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n223 ) , .A2( u0_uk_n635 ) , .B2( u0_uk_n669 ) );
  OAI22_X1 u0_uk_U972 (.ZN( u0_K5_40 ) , .A1( u0_uk_n100 ) , .B1( u0_uk_n182 ) , .A2( u0_uk_n458 ) , .B2( u0_uk_n475 ) );
  OAI22_X1 u0_uk_U991 (.ZN( u0_K1_34 ) , .A1( u0_uk_n118 ) , .B1( u0_uk_n188 ) , .A2( u0_uk_n709 ) , .B2( u0_uk_n714 ) );
  OAI22_X1 u0_uk_U992 (.ZN( u0_K1_47 ) , .A1( u0_uk_n146 ) , .B1( u0_uk_n240 ) , .A2( u0_uk_n711 ) , .B2( u0_uk_n716 ) );
  XOR2_X1 u2_U130 (.B( u2_L11_32 ) , .Z( u2_N415 ) , .A( u2_out12_32 ) );
  XOR2_X1 u2_U131 (.B( u2_L11_31 ) , .Z( u2_N414 ) , .A( u2_out12_31 ) );
  XOR2_X1 u2_U132 (.B( u2_L11_30 ) , .Z( u2_N413 ) , .A( u2_out12_30 ) );
  XOR2_X1 u2_U134 (.B( u2_L11_28 ) , .Z( u2_N411 ) , .A( u2_out12_28 ) );
  XOR2_X1 u2_U135 (.B( u2_L11_27 ) , .Z( u2_N410 ) , .A( u2_out12_27 ) );
  XOR2_X1 u2_U139 (.B( u2_L11_24 ) , .Z( u2_N407 ) , .A( u2_out12_24 ) );
  XOR2_X1 u2_U140 (.B( u2_L11_23 ) , .Z( u2_N406 ) , .A( u2_out12_23 ) );
  XOR2_X1 u2_U141 (.B( u2_L11_22 ) , .Z( u2_N405 ) , .A( u2_out12_22 ) );
  XOR2_X1 u2_U142 (.B( u2_L11_21 ) , .Z( u2_N404 ) , .A( u2_out12_21 ) );
  XOR2_X1 u2_U145 (.B( u2_L11_18 ) , .Z( u2_N401 ) , .A( u2_out12_18 ) );
  XOR2_X1 u2_U146 (.B( u2_L11_17 ) , .Z( u2_N400 ) , .A( u2_out12_17 ) );
  XOR2_X1 u2_U149 (.B( u2_L11_16 ) , .Z( u2_N399 ) , .A( u2_out12_16 ) );
  XOR2_X1 u2_U150 (.B( u2_L11_15 ) , .Z( u2_N398 ) , .A( u2_out12_15 ) );
  XOR2_X1 u2_U152 (.B( u2_L11_13 ) , .Z( u2_N396 ) , .A( u2_out12_13 ) );
  XOR2_X1 u2_U153 (.B( u2_L11_12 ) , .Z( u2_N395 ) , .A( u2_out12_12 ) );
  XOR2_X1 u2_U156 (.B( u2_L11_9 ) , .Z( u2_N392 ) , .A( u2_out12_9 ) );
  XOR2_X1 u2_U158 (.B( u2_L11_7 ) , .Z( u2_N390 ) , .A( u2_out12_7 ) );
  XOR2_X1 u2_U160 (.B( u2_L11_6 ) , .Z( u2_N389 ) , .A( u2_out12_6 ) );
  XOR2_X1 u2_U161 (.B( u2_L11_5 ) , .Z( u2_N388 ) , .A( u2_out12_5 ) );
  XOR2_X1 u2_U164 (.B( u2_L11_2 ) , .Z( u2_N385 ) , .A( u2_out12_2 ) );
  XOR2_X1 u2_U209 (.B( u2_L9_25 ) , .Z( u2_N344 ) , .A( u2_out10_25 ) );
  XOR2_X1 u2_U221 (.B( u2_L9_14 ) , .Z( u2_N333 ) , .A( u2_out10_14 ) );
  XOR2_X1 u2_U228 (.B( u2_L9_8 ) , .Z( u2_N327 ) , .A( u2_out10_8 ) );
  XOR2_X1 u2_U233 (.B( u2_L9_3 ) , .Z( u2_N322 ) , .A( u2_out10_3 ) );
  XOR2_X1 u2_U308 (.B( u2_L6_32 ) , .Z( u2_N255 ) , .A( u2_out7_32 ) );
  XOR2_X1 u2_U311 (.B( u2_L6_29 ) , .Z( u2_N252 ) , .A( u2_out7_29 ) );
  XOR2_X1 u2_U315 (.B( u2_L6_26 ) , .Z( u2_N249 ) , .A( u2_out7_26 ) );
  XOR2_X1 u2_U316 (.B( u2_L6_25 ) , .Z( u2_N248 ) , .A( u2_out7_25 ) );
  XOR2_X1 u2_U319 (.B( u2_L6_22 ) , .Z( u2_N245 ) , .A( u2_out7_22 ) );
  XOR2_X1 u2_U321 (.B( u2_L6_20 ) , .Z( u2_N243 ) , .A( u2_out7_20 ) );
  XOR2_X1 u2_U322 (.B( u2_L6_19 ) , .Z( u2_N242 ) , .A( u2_out7_19 ) );
  XOR2_X1 u2_U328 (.B( u2_L6_14 ) , .Z( u2_N237 ) , .A( u2_out7_14 ) );
  XOR2_X1 u2_U330 (.B( u2_L6_12 ) , .Z( u2_N235 ) , .A( u2_out7_12 ) );
  XOR2_X1 u2_U331 (.B( u2_L6_11 ) , .Z( u2_N234 ) , .A( u2_out7_11 ) );
  XOR2_X1 u2_U332 (.B( u2_L6_10 ) , .Z( u2_N233 ) , .A( u2_out7_10 ) );
  XOR2_X1 u2_U334 (.B( u2_L6_8 ) , .Z( u2_N231 ) , .A( u2_out7_8 ) );
  XOR2_X1 u2_U335 (.B( u2_L6_7 ) , .Z( u2_N230 ) , .A( u2_out7_7 ) );
  XOR2_X1 u2_U339 (.B( u2_L6_4 ) , .Z( u2_N227 ) , .A( u2_out7_4 ) );
  XOR2_X1 u2_U340 (.B( u2_L6_3 ) , .Z( u2_N226 ) , .A( u2_out7_3 ) );
  XOR2_X1 u2_U342 (.B( u2_L6_1 ) , .Z( u2_N224 ) , .A( u2_out7_1 ) );
  XOR2_X1 u2_U387 (.B( u2_L4_25 ) , .Z( u2_N184 ) , .A( u2_out5_25 ) );
  XOR2_X1 u2_U399 (.B( u2_L4_14 ) , .Z( u2_N173 ) , .A( u2_out5_14 ) );
  XOR2_X1 u2_U406 (.B( u2_L4_8 ) , .Z( u2_N167 ) , .A( u2_out5_8 ) );
  XOR2_X1 u2_U411 (.B( u2_L4_3 ) , .Z( u2_N162 ) , .A( u2_out5_3 ) );
  XOR2_X1 u2_U451 (.B( u2_L2_31 ) , .Z( u2_N126 ) , .A( u2_out3_31 ) );
  XOR2_X1 u2_U454 (.B( u2_L2_28 ) , .Z( u2_N123 ) , .A( u2_out3_28 ) );
  XOR2_X1 u2_U455 (.B( u2_L2_27 ) , .Z( u2_N122 ) , .A( u2_out3_27 ) );
  XOR2_X1 u2_U460 (.B( u2_L2_23 ) , .Z( u2_N118 ) , .A( u2_out3_23 ) );
  XOR2_X1 u2_U462 (.B( u2_L2_21 ) , .Z( u2_N116 ) , .A( u2_out3_21 ) );
  XOR2_X1 u2_U465 (.B( u2_L2_18 ) , .Z( u2_N113 ) , .A( u2_out3_18 ) );
  XOR2_X1 u2_U466 (.B( u2_L2_17 ) , .Z( u2_N112 ) , .A( u2_out3_17 ) );
  XOR2_X1 u2_U468 (.B( u2_L2_15 ) , .Z( u2_N110 ) , .A( u2_out3_15 ) );
  XOR2_X1 u2_U471 (.B( u2_L2_13 ) , .Z( u2_N108 ) , .A( u2_out3_13 ) );
  XOR2_X1 u2_U475 (.B( u2_L2_9 ) , .Z( u2_N104 ) , .A( u2_out3_9 ) );
  XOR2_X1 u2_U479 (.B( u2_L2_5 ) , .Z( u2_N100 ) , .A( u2_out3_5 ) );
  XOR2_X1 u2_U5 (.B( u2_L2_2 ) , .Z( u2_N97 ) , .A( u2_out3_2 ) );
  XOR2_X1 u2_u10_U26 (.B( u2_K11_30 ) , .A( u2_R9_21 ) , .Z( u2_u10_X_30 ) );
  XOR2_X1 u2_u10_U28 (.B( u2_K11_29 ) , .A( u2_R9_20 ) , .Z( u2_u10_X_29 ) );
  XOR2_X1 u2_u10_U29 (.B( u2_K11_28 ) , .A( u2_R9_19 ) , .Z( u2_u10_X_28 ) );
  XOR2_X1 u2_u10_U30 (.B( u2_K11_27 ) , .A( u2_R9_18 ) , .Z( u2_u10_X_27 ) );
  XOR2_X1 u2_u10_U31 (.B( u2_K11_26 ) , .A( u2_R9_17 ) , .Z( u2_u10_X_26 ) );
  XOR2_X1 u2_u10_U32 (.B( u2_K11_25 ) , .A( u2_R9_16 ) , .Z( u2_u10_X_25 ) );
  AOI21_X1 u2_u10_u4_U10 (.ZN( u2_u10_u4_n106 ) , .B2( u2_u10_u4_n146 ) , .B1( u2_u10_u4_n158 ) , .A( u2_u10_u4_n170 ) );
  AOI21_X1 u2_u10_u4_U11 (.ZN( u2_u10_u4_n108 ) , .B2( u2_u10_u4_n134 ) , .B1( u2_u10_u4_n155 ) , .A( u2_u10_u4_n156 ) );
  AOI21_X1 u2_u10_u4_U12 (.ZN( u2_u10_u4_n109 ) , .A( u2_u10_u4_n153 ) , .B1( u2_u10_u4_n159 ) , .B2( u2_u10_u4_n184 ) );
  AOI211_X1 u2_u10_u4_U13 (.B( u2_u10_u4_n136 ) , .A( u2_u10_u4_n137 ) , .C2( u2_u10_u4_n138 ) , .ZN( u2_u10_u4_n139 ) , .C1( u2_u10_u4_n182 ) );
  OAI22_X1 u2_u10_u4_U14 (.B2( u2_u10_u4_n135 ) , .ZN( u2_u10_u4_n137 ) , .B1( u2_u10_u4_n153 ) , .A1( u2_u10_u4_n155 ) , .A2( u2_u10_u4_n171 ) );
  AND3_X1 u2_u10_u4_U15 (.A2( u2_u10_u4_n134 ) , .ZN( u2_u10_u4_n135 ) , .A3( u2_u10_u4_n145 ) , .A1( u2_u10_u4_n157 ) );
  NAND2_X1 u2_u10_u4_U16 (.ZN( u2_u10_u4_n132 ) , .A2( u2_u10_u4_n170 ) , .A1( u2_u10_u4_n173 ) );
  AOI21_X1 u2_u10_u4_U17 (.B2( u2_u10_u4_n160 ) , .B1( u2_u10_u4_n161 ) , .ZN( u2_u10_u4_n162 ) , .A( u2_u10_u4_n170 ) );
  AOI21_X1 u2_u10_u4_U18 (.ZN( u2_u10_u4_n107 ) , .B2( u2_u10_u4_n143 ) , .A( u2_u10_u4_n174 ) , .B1( u2_u10_u4_n184 ) );
  AOI21_X1 u2_u10_u4_U19 (.B2( u2_u10_u4_n158 ) , .B1( u2_u10_u4_n159 ) , .ZN( u2_u10_u4_n163 ) , .A( u2_u10_u4_n174 ) );
  AOI21_X1 u2_u10_u4_U20 (.A( u2_u10_u4_n153 ) , .B2( u2_u10_u4_n154 ) , .B1( u2_u10_u4_n155 ) , .ZN( u2_u10_u4_n165 ) );
  AOI21_X1 u2_u10_u4_U21 (.A( u2_u10_u4_n156 ) , .B2( u2_u10_u4_n157 ) , .ZN( u2_u10_u4_n164 ) , .B1( u2_u10_u4_n184 ) );
  INV_X1 u2_u10_u4_U22 (.A( u2_u10_u4_n138 ) , .ZN( u2_u10_u4_n170 ) );
  AND2_X1 u2_u10_u4_U23 (.A2( u2_u10_u4_n120 ) , .ZN( u2_u10_u4_n155 ) , .A1( u2_u10_u4_n160 ) );
  INV_X1 u2_u10_u4_U24 (.A( u2_u10_u4_n156 ) , .ZN( u2_u10_u4_n175 ) );
  NAND2_X1 u2_u10_u4_U25 (.A2( u2_u10_u4_n118 ) , .ZN( u2_u10_u4_n131 ) , .A1( u2_u10_u4_n147 ) );
  NAND2_X1 u2_u10_u4_U26 (.A1( u2_u10_u4_n119 ) , .A2( u2_u10_u4_n120 ) , .ZN( u2_u10_u4_n130 ) );
  NAND2_X1 u2_u10_u4_U27 (.ZN( u2_u10_u4_n117 ) , .A2( u2_u10_u4_n118 ) , .A1( u2_u10_u4_n148 ) );
  NAND2_X1 u2_u10_u4_U28 (.ZN( u2_u10_u4_n129 ) , .A1( u2_u10_u4_n134 ) , .A2( u2_u10_u4_n148 ) );
  AND3_X1 u2_u10_u4_U29 (.A1( u2_u10_u4_n119 ) , .A2( u2_u10_u4_n143 ) , .A3( u2_u10_u4_n154 ) , .ZN( u2_u10_u4_n161 ) );
  NOR2_X1 u2_u10_u4_U3 (.ZN( u2_u10_u4_n121 ) , .A1( u2_u10_u4_n181 ) , .A2( u2_u10_u4_n182 ) );
  AND2_X1 u2_u10_u4_U30 (.A1( u2_u10_u4_n145 ) , .A2( u2_u10_u4_n147 ) , .ZN( u2_u10_u4_n159 ) );
  OR3_X1 u2_u10_u4_U31 (.A3( u2_u10_u4_n114 ) , .A2( u2_u10_u4_n115 ) , .A1( u2_u10_u4_n116 ) , .ZN( u2_u10_u4_n136 ) );
  AOI21_X1 u2_u10_u4_U32 (.A( u2_u10_u4_n113 ) , .ZN( u2_u10_u4_n116 ) , .B2( u2_u10_u4_n173 ) , .B1( u2_u10_u4_n174 ) );
  AOI21_X1 u2_u10_u4_U33 (.ZN( u2_u10_u4_n115 ) , .B2( u2_u10_u4_n145 ) , .B1( u2_u10_u4_n146 ) , .A( u2_u10_u4_n156 ) );
  OAI22_X1 u2_u10_u4_U34 (.ZN( u2_u10_u4_n114 ) , .A2( u2_u10_u4_n121 ) , .B1( u2_u10_u4_n160 ) , .B2( u2_u10_u4_n170 ) , .A1( u2_u10_u4_n171 ) );
  INV_X1 u2_u10_u4_U35 (.A( u2_u10_u4_n158 ) , .ZN( u2_u10_u4_n182 ) );
  INV_X1 u2_u10_u4_U36 (.ZN( u2_u10_u4_n181 ) , .A( u2_u10_u4_n96 ) );
  INV_X1 u2_u10_u4_U37 (.A( u2_u10_u4_n144 ) , .ZN( u2_u10_u4_n179 ) );
  INV_X1 u2_u10_u4_U38 (.A( u2_u10_u4_n157 ) , .ZN( u2_u10_u4_n178 ) );
  NAND2_X1 u2_u10_u4_U39 (.A2( u2_u10_u4_n154 ) , .A1( u2_u10_u4_n96 ) , .ZN( u2_u10_u4_n97 ) );
  INV_X1 u2_u10_u4_U4 (.A( u2_u10_u4_n117 ) , .ZN( u2_u10_u4_n184 ) );
  INV_X1 u2_u10_u4_U40 (.A( u2_u10_u4_n143 ) , .ZN( u2_u10_u4_n183 ) );
  NOR2_X1 u2_u10_u4_U41 (.ZN( u2_u10_u4_n138 ) , .A1( u2_u10_u4_n168 ) , .A2( u2_u10_u4_n169 ) );
  NOR2_X1 u2_u10_u4_U42 (.A1( u2_u10_u4_n150 ) , .A2( u2_u10_u4_n152 ) , .ZN( u2_u10_u4_n153 ) );
  NOR2_X1 u2_u10_u4_U43 (.A2( u2_u10_u4_n128 ) , .A1( u2_u10_u4_n138 ) , .ZN( u2_u10_u4_n156 ) );
  AOI22_X1 u2_u10_u4_U44 (.B2( u2_u10_u4_n122 ) , .A1( u2_u10_u4_n123 ) , .ZN( u2_u10_u4_n124 ) , .B1( u2_u10_u4_n128 ) , .A2( u2_u10_u4_n172 ) );
  INV_X1 u2_u10_u4_U45 (.A( u2_u10_u4_n153 ) , .ZN( u2_u10_u4_n172 ) );
  NAND2_X1 u2_u10_u4_U46 (.A2( u2_u10_u4_n120 ) , .ZN( u2_u10_u4_n123 ) , .A1( u2_u10_u4_n161 ) );
  AOI22_X1 u2_u10_u4_U47 (.B2( u2_u10_u4_n132 ) , .A2( u2_u10_u4_n133 ) , .ZN( u2_u10_u4_n140 ) , .A1( u2_u10_u4_n150 ) , .B1( u2_u10_u4_n179 ) );
  NAND2_X1 u2_u10_u4_U48 (.ZN( u2_u10_u4_n133 ) , .A2( u2_u10_u4_n146 ) , .A1( u2_u10_u4_n154 ) );
  NAND2_X1 u2_u10_u4_U49 (.A1( u2_u10_u4_n103 ) , .ZN( u2_u10_u4_n154 ) , .A2( u2_u10_u4_n98 ) );
  INV_X1 u2_u10_u4_U5 (.ZN( u2_u10_u4_n186 ) , .A( u2_u10_u4_n95 ) );
  NAND2_X1 u2_u10_u4_U50 (.A1( u2_u10_u4_n101 ) , .ZN( u2_u10_u4_n158 ) , .A2( u2_u10_u4_n99 ) );
  AOI21_X1 u2_u10_u4_U51 (.ZN( u2_u10_u4_n127 ) , .A( u2_u10_u4_n136 ) , .B2( u2_u10_u4_n150 ) , .B1( u2_u10_u4_n180 ) );
  INV_X1 u2_u10_u4_U52 (.A( u2_u10_u4_n160 ) , .ZN( u2_u10_u4_n180 ) );
  NAND2_X1 u2_u10_u4_U53 (.A2( u2_u10_u4_n104 ) , .A1( u2_u10_u4_n105 ) , .ZN( u2_u10_u4_n146 ) );
  NAND2_X1 u2_u10_u4_U54 (.A2( u2_u10_u4_n101 ) , .A1( u2_u10_u4_n102 ) , .ZN( u2_u10_u4_n160 ) );
  NAND2_X1 u2_u10_u4_U55 (.ZN( u2_u10_u4_n134 ) , .A1( u2_u10_u4_n98 ) , .A2( u2_u10_u4_n99 ) );
  NAND2_X1 u2_u10_u4_U56 (.A1( u2_u10_u4_n103 ) , .A2( u2_u10_u4_n104 ) , .ZN( u2_u10_u4_n143 ) );
  NAND2_X1 u2_u10_u4_U57 (.A2( u2_u10_u4_n105 ) , .ZN( u2_u10_u4_n145 ) , .A1( u2_u10_u4_n98 ) );
  NAND2_X1 u2_u10_u4_U58 (.A1( u2_u10_u4_n100 ) , .A2( u2_u10_u4_n105 ) , .ZN( u2_u10_u4_n120 ) );
  NAND2_X1 u2_u10_u4_U59 (.A1( u2_u10_u4_n102 ) , .A2( u2_u10_u4_n104 ) , .ZN( u2_u10_u4_n148 ) );
  OAI221_X1 u2_u10_u4_U6 (.C1( u2_u10_u4_n134 ) , .B1( u2_u10_u4_n158 ) , .B2( u2_u10_u4_n171 ) , .C2( u2_u10_u4_n173 ) , .A( u2_u10_u4_n94 ) , .ZN( u2_u10_u4_n95 ) );
  NAND2_X1 u2_u10_u4_U60 (.A2( u2_u10_u4_n100 ) , .A1( u2_u10_u4_n103 ) , .ZN( u2_u10_u4_n157 ) );
  INV_X1 u2_u10_u4_U61 (.A( u2_u10_u4_n150 ) , .ZN( u2_u10_u4_n173 ) );
  INV_X1 u2_u10_u4_U62 (.A( u2_u10_u4_n152 ) , .ZN( u2_u10_u4_n171 ) );
  NAND2_X1 u2_u10_u4_U63 (.A1( u2_u10_u4_n100 ) , .ZN( u2_u10_u4_n118 ) , .A2( u2_u10_u4_n99 ) );
  NAND2_X1 u2_u10_u4_U64 (.A2( u2_u10_u4_n100 ) , .A1( u2_u10_u4_n102 ) , .ZN( u2_u10_u4_n144 ) );
  NAND2_X1 u2_u10_u4_U65 (.A2( u2_u10_u4_n101 ) , .A1( u2_u10_u4_n105 ) , .ZN( u2_u10_u4_n96 ) );
  INV_X1 u2_u10_u4_U66 (.A( u2_u10_u4_n128 ) , .ZN( u2_u10_u4_n174 ) );
  NAND2_X1 u2_u10_u4_U67 (.A2( u2_u10_u4_n102 ) , .ZN( u2_u10_u4_n119 ) , .A1( u2_u10_u4_n98 ) );
  NAND2_X1 u2_u10_u4_U68 (.A2( u2_u10_u4_n101 ) , .A1( u2_u10_u4_n103 ) , .ZN( u2_u10_u4_n147 ) );
  NAND2_X1 u2_u10_u4_U69 (.A2( u2_u10_u4_n104 ) , .ZN( u2_u10_u4_n113 ) , .A1( u2_u10_u4_n99 ) );
  AOI222_X1 u2_u10_u4_U7 (.B2( u2_u10_u4_n132 ) , .A1( u2_u10_u4_n138 ) , .C2( u2_u10_u4_n175 ) , .A2( u2_u10_u4_n179 ) , .C1( u2_u10_u4_n181 ) , .B1( u2_u10_u4_n185 ) , .ZN( u2_u10_u4_n94 ) );
  NOR2_X1 u2_u10_u4_U70 (.A2( u2_u10_X_28 ) , .ZN( u2_u10_u4_n150 ) , .A1( u2_u10_u4_n168 ) );
  NOR2_X1 u2_u10_u4_U71 (.A2( u2_u10_X_29 ) , .ZN( u2_u10_u4_n152 ) , .A1( u2_u10_u4_n169 ) );
  NOR2_X1 u2_u10_u4_U72 (.A2( u2_u10_X_30 ) , .ZN( u2_u10_u4_n105 ) , .A1( u2_u10_u4_n176 ) );
  NOR2_X1 u2_u10_u4_U73 (.A2( u2_u10_X_26 ) , .ZN( u2_u10_u4_n100 ) , .A1( u2_u10_u4_n177 ) );
  NOR2_X1 u2_u10_u4_U74 (.A2( u2_u10_X_28 ) , .A1( u2_u10_X_29 ) , .ZN( u2_u10_u4_n128 ) );
  NOR2_X1 u2_u10_u4_U75 (.A2( u2_u10_X_27 ) , .A1( u2_u10_X_30 ) , .ZN( u2_u10_u4_n102 ) );
  NOR2_X1 u2_u10_u4_U76 (.A2( u2_u10_X_25 ) , .A1( u2_u10_X_26 ) , .ZN( u2_u10_u4_n98 ) );
  AND2_X1 u2_u10_u4_U77 (.A2( u2_u10_X_25 ) , .A1( u2_u10_X_26 ) , .ZN( u2_u10_u4_n104 ) );
  AND2_X1 u2_u10_u4_U78 (.A1( u2_u10_X_30 ) , .A2( u2_u10_u4_n176 ) , .ZN( u2_u10_u4_n99 ) );
  AND2_X1 u2_u10_u4_U79 (.A1( u2_u10_X_26 ) , .ZN( u2_u10_u4_n101 ) , .A2( u2_u10_u4_n177 ) );
  INV_X1 u2_u10_u4_U8 (.A( u2_u10_u4_n113 ) , .ZN( u2_u10_u4_n185 ) );
  AND2_X1 u2_u10_u4_U80 (.A1( u2_u10_X_27 ) , .A2( u2_u10_X_30 ) , .ZN( u2_u10_u4_n103 ) );
  INV_X1 u2_u10_u4_U81 (.A( u2_u10_X_28 ) , .ZN( u2_u10_u4_n169 ) );
  INV_X1 u2_u10_u4_U82 (.A( u2_u10_X_29 ) , .ZN( u2_u10_u4_n168 ) );
  INV_X1 u2_u10_u4_U83 (.A( u2_u10_X_25 ) , .ZN( u2_u10_u4_n177 ) );
  INV_X1 u2_u10_u4_U84 (.A( u2_u10_X_27 ) , .ZN( u2_u10_u4_n176 ) );
  NAND4_X1 u2_u10_u4_U85 (.ZN( u2_out10_25 ) , .A4( u2_u10_u4_n139 ) , .A3( u2_u10_u4_n140 ) , .A2( u2_u10_u4_n141 ) , .A1( u2_u10_u4_n142 ) );
  OAI21_X1 u2_u10_u4_U86 (.A( u2_u10_u4_n128 ) , .B2( u2_u10_u4_n129 ) , .B1( u2_u10_u4_n130 ) , .ZN( u2_u10_u4_n142 ) );
  OAI21_X1 u2_u10_u4_U87 (.B2( u2_u10_u4_n131 ) , .ZN( u2_u10_u4_n141 ) , .A( u2_u10_u4_n175 ) , .B1( u2_u10_u4_n183 ) );
  NAND4_X1 u2_u10_u4_U88 (.ZN( u2_out10_14 ) , .A4( u2_u10_u4_n124 ) , .A3( u2_u10_u4_n125 ) , .A2( u2_u10_u4_n126 ) , .A1( u2_u10_u4_n127 ) );
  AOI22_X1 u2_u10_u4_U89 (.B2( u2_u10_u4_n117 ) , .ZN( u2_u10_u4_n126 ) , .A1( u2_u10_u4_n129 ) , .B1( u2_u10_u4_n152 ) , .A2( u2_u10_u4_n175 ) );
  NOR4_X1 u2_u10_u4_U9 (.A4( u2_u10_u4_n106 ) , .A3( u2_u10_u4_n107 ) , .A2( u2_u10_u4_n108 ) , .A1( u2_u10_u4_n109 ) , .ZN( u2_u10_u4_n110 ) );
  AOI22_X1 u2_u10_u4_U90 (.ZN( u2_u10_u4_n125 ) , .B2( u2_u10_u4_n131 ) , .A2( u2_u10_u4_n132 ) , .B1( u2_u10_u4_n138 ) , .A1( u2_u10_u4_n178 ) );
  NAND4_X1 u2_u10_u4_U91 (.ZN( u2_out10_8 ) , .A4( u2_u10_u4_n110 ) , .A3( u2_u10_u4_n111 ) , .A2( u2_u10_u4_n112 ) , .A1( u2_u10_u4_n186 ) );
  NAND2_X1 u2_u10_u4_U92 (.ZN( u2_u10_u4_n112 ) , .A2( u2_u10_u4_n130 ) , .A1( u2_u10_u4_n150 ) );
  AOI22_X1 u2_u10_u4_U93 (.ZN( u2_u10_u4_n111 ) , .B2( u2_u10_u4_n132 ) , .A1( u2_u10_u4_n152 ) , .B1( u2_u10_u4_n178 ) , .A2( u2_u10_u4_n97 ) );
  AOI22_X1 u2_u10_u4_U94 (.B2( u2_u10_u4_n149 ) , .B1( u2_u10_u4_n150 ) , .A2( u2_u10_u4_n151 ) , .A1( u2_u10_u4_n152 ) , .ZN( u2_u10_u4_n167 ) );
  NOR4_X1 u2_u10_u4_U95 (.A4( u2_u10_u4_n162 ) , .A3( u2_u10_u4_n163 ) , .A2( u2_u10_u4_n164 ) , .A1( u2_u10_u4_n165 ) , .ZN( u2_u10_u4_n166 ) );
  NAND3_X1 u2_u10_u4_U96 (.ZN( u2_out10_3 ) , .A3( u2_u10_u4_n166 ) , .A1( u2_u10_u4_n167 ) , .A2( u2_u10_u4_n186 ) );
  NAND3_X1 u2_u10_u4_U97 (.A3( u2_u10_u4_n146 ) , .A2( u2_u10_u4_n147 ) , .A1( u2_u10_u4_n148 ) , .ZN( u2_u10_u4_n149 ) );
  NAND3_X1 u2_u10_u4_U98 (.A3( u2_u10_u4_n143 ) , .A2( u2_u10_u4_n144 ) , .A1( u2_u10_u4_n145 ) , .ZN( u2_u10_u4_n151 ) );
  NAND3_X1 u2_u10_u4_U99 (.A3( u2_u10_u4_n121 ) , .ZN( u2_u10_u4_n122 ) , .A2( u2_u10_u4_n144 ) , .A1( u2_u10_u4_n154 ) );
  XOR2_X1 u2_u12_U1 (.B( u2_K13_9 ) , .A( u2_R11_6 ) , .Z( u2_u12_X_9 ) );
  XOR2_X1 u2_u12_U10 (.B( u2_K13_45 ) , .A( u2_R11_30 ) , .Z( u2_u12_X_45 ) );
  XOR2_X1 u2_u12_U11 (.B( u2_K13_44 ) , .A( u2_R11_29 ) , .Z( u2_u12_X_44 ) );
  XOR2_X1 u2_u12_U12 (.B( u2_K13_43 ) , .A( u2_R11_28 ) , .Z( u2_u12_X_43 ) );
  XOR2_X1 u2_u12_U13 (.B( u2_K13_42 ) , .A( u2_R11_29 ) , .Z( u2_u12_X_42 ) );
  XOR2_X1 u2_u12_U14 (.B( u2_K13_41 ) , .A( u2_R11_28 ) , .Z( u2_u12_X_41 ) );
  XOR2_X1 u2_u12_U15 (.B( u2_K13_40 ) , .A( u2_R11_27 ) , .Z( u2_u12_X_40 ) );
  XOR2_X1 u2_u12_U16 (.B( u2_K13_3 ) , .A( u2_R11_2 ) , .Z( u2_u12_X_3 ) );
  XOR2_X1 u2_u12_U17 (.B( u2_K13_39 ) , .A( u2_R11_26 ) , .Z( u2_u12_X_39 ) );
  XOR2_X1 u2_u12_U18 (.B( u2_K13_38 ) , .A( u2_R11_25 ) , .Z( u2_u12_X_38 ) );
  XOR2_X1 u2_u12_U19 (.B( u2_K13_37 ) , .A( u2_R11_24 ) , .Z( u2_u12_X_37 ) );
  XOR2_X1 u2_u12_U2 (.B( u2_K13_8 ) , .A( u2_R11_5 ) , .Z( u2_u12_X_8 ) );
  XOR2_X1 u2_u12_U27 (.B( u2_K13_2 ) , .A( u2_R11_1 ) , .Z( u2_u12_X_2 ) );
  XOR2_X1 u2_u12_U3 (.B( u2_K13_7 ) , .A( u2_R11_4 ) , .Z( u2_u12_X_7 ) );
  XOR2_X1 u2_u12_U38 (.B( u2_K13_1 ) , .A( u2_R11_32 ) , .Z( u2_u12_X_1 ) );
  XOR2_X1 u2_u12_U4 (.B( u2_K13_6 ) , .A( u2_R11_5 ) , .Z( u2_u12_X_6 ) );
  XOR2_X1 u2_u12_U40 (.B( u2_K13_18 ) , .A( u2_R11_13 ) , .Z( u2_u12_X_18 ) );
  XOR2_X1 u2_u12_U41 (.B( u2_K13_17 ) , .A( u2_R11_12 ) , .Z( u2_u12_X_17 ) );
  XOR2_X1 u2_u12_U42 (.B( u2_K13_16 ) , .A( u2_R11_11 ) , .Z( u2_u12_X_16 ) );
  XOR2_X1 u2_u12_U43 (.B( u2_K13_15 ) , .A( u2_R11_10 ) , .Z( u2_u12_X_15 ) );
  XOR2_X1 u2_u12_U44 (.B( u2_K13_14 ) , .A( u2_R11_9 ) , .Z( u2_u12_X_14 ) );
  XOR2_X1 u2_u12_U45 (.B( u2_K13_13 ) , .A( u2_R11_8 ) , .Z( u2_u12_X_13 ) );
  XOR2_X1 u2_u12_U46 (.B( u2_K13_12 ) , .A( u2_R11_9 ) , .Z( u2_u12_X_12 ) );
  XOR2_X1 u2_u12_U47 (.B( u2_K13_11 ) , .A( u2_R11_8 ) , .Z( u2_u12_X_11 ) );
  XOR2_X1 u2_u12_U48 (.B( u2_K13_10 ) , .A( u2_R11_7 ) , .Z( u2_u12_X_10 ) );
  XOR2_X1 u2_u12_U5 (.B( u2_K13_5 ) , .A( u2_R11_4 ) , .Z( u2_u12_X_5 ) );
  XOR2_X1 u2_u12_U6 (.B( u2_K13_4 ) , .A( u2_R11_3 ) , .Z( u2_u12_X_4 ) );
  XOR2_X1 u2_u12_U7 (.B( u2_K13_48 ) , .A( u2_R11_1 ) , .Z( u2_u12_X_48 ) );
  XOR2_X1 u2_u12_U8 (.B( u2_K13_47 ) , .A( u2_R11_32 ) , .Z( u2_u12_X_47 ) );
  XOR2_X1 u2_u12_U9 (.B( u2_K13_46 ) , .A( u2_R11_31 ) , .Z( u2_u12_X_46 ) );
  AND2_X1 u2_u12_u0_U10 (.A1( u2_u12_u0_n131 ) , .ZN( u2_u12_u0_n141 ) , .A2( u2_u12_u0_n150 ) );
  AND3_X1 u2_u12_u0_U11 (.A2( u2_u12_u0_n112 ) , .ZN( u2_u12_u0_n127 ) , .A3( u2_u12_u0_n130 ) , .A1( u2_u12_u0_n148 ) );
  AND2_X1 u2_u12_u0_U12 (.ZN( u2_u12_u0_n107 ) , .A1( u2_u12_u0_n130 ) , .A2( u2_u12_u0_n140 ) );
  AND2_X1 u2_u12_u0_U13 (.A2( u2_u12_u0_n129 ) , .A1( u2_u12_u0_n130 ) , .ZN( u2_u12_u0_n151 ) );
  AND2_X1 u2_u12_u0_U14 (.A1( u2_u12_u0_n108 ) , .A2( u2_u12_u0_n125 ) , .ZN( u2_u12_u0_n145 ) );
  INV_X1 u2_u12_u0_U15 (.A( u2_u12_u0_n143 ) , .ZN( u2_u12_u0_n173 ) );
  NOR2_X1 u2_u12_u0_U16 (.A2( u2_u12_u0_n136 ) , .ZN( u2_u12_u0_n147 ) , .A1( u2_u12_u0_n160 ) );
  AOI21_X1 u2_u12_u0_U17 (.B1( u2_u12_u0_n103 ) , .ZN( u2_u12_u0_n132 ) , .A( u2_u12_u0_n165 ) , .B2( u2_u12_u0_n93 ) );
  OAI22_X1 u2_u12_u0_U18 (.B1( u2_u12_u0_n125 ) , .ZN( u2_u12_u0_n126 ) , .A1( u2_u12_u0_n138 ) , .A2( u2_u12_u0_n146 ) , .B2( u2_u12_u0_n147 ) );
  OAI22_X1 u2_u12_u0_U19 (.B1( u2_u12_u0_n131 ) , .A1( u2_u12_u0_n144 ) , .B2( u2_u12_u0_n147 ) , .A2( u2_u12_u0_n90 ) , .ZN( u2_u12_u0_n91 ) );
  AND3_X1 u2_u12_u0_U20 (.A3( u2_u12_u0_n121 ) , .A2( u2_u12_u0_n125 ) , .A1( u2_u12_u0_n148 ) , .ZN( u2_u12_u0_n90 ) );
  NOR2_X1 u2_u12_u0_U21 (.A1( u2_u12_u0_n163 ) , .A2( u2_u12_u0_n164 ) , .ZN( u2_u12_u0_n95 ) );
  AOI22_X1 u2_u12_u0_U22 (.B2( u2_u12_u0_n109 ) , .A2( u2_u12_u0_n110 ) , .ZN( u2_u12_u0_n111 ) , .B1( u2_u12_u0_n118 ) , .A1( u2_u12_u0_n160 ) );
  NAND2_X1 u2_u12_u0_U23 (.A1( u2_u12_u0_n100 ) , .A2( u2_u12_u0_n103 ) , .ZN( u2_u12_u0_n125 ) );
  INV_X1 u2_u12_u0_U24 (.A( u2_u12_u0_n136 ) , .ZN( u2_u12_u0_n161 ) );
  INV_X1 u2_u12_u0_U25 (.A( u2_u12_u0_n118 ) , .ZN( u2_u12_u0_n158 ) );
  AOI21_X1 u2_u12_u0_U26 (.B1( u2_u12_u0_n127 ) , .B2( u2_u12_u0_n129 ) , .A( u2_u12_u0_n138 ) , .ZN( u2_u12_u0_n96 ) );
  AOI21_X1 u2_u12_u0_U27 (.ZN( u2_u12_u0_n104 ) , .B1( u2_u12_u0_n107 ) , .B2( u2_u12_u0_n141 ) , .A( u2_u12_u0_n144 ) );
  NAND2_X1 u2_u12_u0_U28 (.A2( u2_u12_u0_n102 ) , .A1( u2_u12_u0_n103 ) , .ZN( u2_u12_u0_n149 ) );
  NAND2_X1 u2_u12_u0_U29 (.A2( u2_u12_u0_n100 ) , .ZN( u2_u12_u0_n131 ) , .A1( u2_u12_u0_n92 ) );
  INV_X1 u2_u12_u0_U3 (.A( u2_u12_u0_n113 ) , .ZN( u2_u12_u0_n166 ) );
  NAND2_X1 u2_u12_u0_U30 (.A2( u2_u12_u0_n102 ) , .ZN( u2_u12_u0_n114 ) , .A1( u2_u12_u0_n92 ) );
  NOR2_X1 u2_u12_u0_U31 (.A1( u2_u12_u0_n120 ) , .ZN( u2_u12_u0_n143 ) , .A2( u2_u12_u0_n167 ) );
  OAI221_X1 u2_u12_u0_U32 (.C1( u2_u12_u0_n112 ) , .ZN( u2_u12_u0_n120 ) , .B1( u2_u12_u0_n138 ) , .B2( u2_u12_u0_n141 ) , .C2( u2_u12_u0_n147 ) , .A( u2_u12_u0_n172 ) );
  AOI211_X1 u2_u12_u0_U33 (.B( u2_u12_u0_n115 ) , .A( u2_u12_u0_n116 ) , .C2( u2_u12_u0_n117 ) , .C1( u2_u12_u0_n118 ) , .ZN( u2_u12_u0_n119 ) );
  NAND2_X1 u2_u12_u0_U34 (.A1( u2_u12_u0_n101 ) , .A2( u2_u12_u0_n102 ) , .ZN( u2_u12_u0_n150 ) );
  INV_X1 u2_u12_u0_U35 (.A( u2_u12_u0_n138 ) , .ZN( u2_u12_u0_n160 ) );
  NAND2_X1 u2_u12_u0_U36 (.A2( u2_u12_u0_n100 ) , .A1( u2_u12_u0_n101 ) , .ZN( u2_u12_u0_n139 ) );
  NAND2_X1 u2_u12_u0_U37 (.ZN( u2_u12_u0_n112 ) , .A2( u2_u12_u0_n92 ) , .A1( u2_u12_u0_n93 ) );
  INV_X1 u2_u12_u0_U38 (.ZN( u2_u12_u0_n172 ) , .A( u2_u12_u0_n88 ) );
  OAI222_X1 u2_u12_u0_U39 (.C1( u2_u12_u0_n108 ) , .A1( u2_u12_u0_n125 ) , .B2( u2_u12_u0_n128 ) , .B1( u2_u12_u0_n144 ) , .A2( u2_u12_u0_n158 ) , .C2( u2_u12_u0_n161 ) , .ZN( u2_u12_u0_n88 ) );
  AOI21_X1 u2_u12_u0_U4 (.B1( u2_u12_u0_n114 ) , .ZN( u2_u12_u0_n115 ) , .B2( u2_u12_u0_n129 ) , .A( u2_u12_u0_n161 ) );
  NAND2_X1 u2_u12_u0_U40 (.A2( u2_u12_u0_n101 ) , .ZN( u2_u12_u0_n121 ) , .A1( u2_u12_u0_n93 ) );
  OR3_X1 u2_u12_u0_U41 (.A3( u2_u12_u0_n152 ) , .A2( u2_u12_u0_n153 ) , .A1( u2_u12_u0_n154 ) , .ZN( u2_u12_u0_n155 ) );
  AOI21_X1 u2_u12_u0_U42 (.B2( u2_u12_u0_n150 ) , .B1( u2_u12_u0_n151 ) , .ZN( u2_u12_u0_n152 ) , .A( u2_u12_u0_n158 ) );
  AOI21_X1 u2_u12_u0_U43 (.A( u2_u12_u0_n144 ) , .B2( u2_u12_u0_n145 ) , .B1( u2_u12_u0_n146 ) , .ZN( u2_u12_u0_n154 ) );
  AOI21_X1 u2_u12_u0_U44 (.A( u2_u12_u0_n147 ) , .B2( u2_u12_u0_n148 ) , .B1( u2_u12_u0_n149 ) , .ZN( u2_u12_u0_n153 ) );
  INV_X1 u2_u12_u0_U45 (.ZN( u2_u12_u0_n171 ) , .A( u2_u12_u0_n99 ) );
  OAI211_X1 u2_u12_u0_U46 (.C2( u2_u12_u0_n140 ) , .C1( u2_u12_u0_n161 ) , .A( u2_u12_u0_n169 ) , .B( u2_u12_u0_n98 ) , .ZN( u2_u12_u0_n99 ) );
  INV_X1 u2_u12_u0_U47 (.ZN( u2_u12_u0_n169 ) , .A( u2_u12_u0_n91 ) );
  AOI211_X1 u2_u12_u0_U48 (.C1( u2_u12_u0_n118 ) , .A( u2_u12_u0_n123 ) , .B( u2_u12_u0_n96 ) , .C2( u2_u12_u0_n97 ) , .ZN( u2_u12_u0_n98 ) );
  NOR2_X1 u2_u12_u0_U49 (.A2( u2_u12_X_4 ) , .A1( u2_u12_X_5 ) , .ZN( u2_u12_u0_n118 ) );
  NOR2_X1 u2_u12_u0_U5 (.A1( u2_u12_u0_n108 ) , .ZN( u2_u12_u0_n123 ) , .A2( u2_u12_u0_n158 ) );
  NOR2_X1 u2_u12_u0_U50 (.A2( u2_u12_X_1 ) , .ZN( u2_u12_u0_n101 ) , .A1( u2_u12_u0_n163 ) );
  NAND2_X1 u2_u12_u0_U51 (.A2( u2_u12_X_4 ) , .A1( u2_u12_X_5 ) , .ZN( u2_u12_u0_n144 ) );
  NOR2_X1 u2_u12_u0_U52 (.A2( u2_u12_X_5 ) , .ZN( u2_u12_u0_n136 ) , .A1( u2_u12_u0_n159 ) );
  NAND2_X1 u2_u12_u0_U53 (.A1( u2_u12_X_5 ) , .ZN( u2_u12_u0_n138 ) , .A2( u2_u12_u0_n159 ) );
  AND2_X1 u2_u12_u0_U54 (.A2( u2_u12_X_3 ) , .A1( u2_u12_X_6 ) , .ZN( u2_u12_u0_n102 ) );
  INV_X1 u2_u12_u0_U55 (.A( u2_u12_X_4 ) , .ZN( u2_u12_u0_n159 ) );
  INV_X1 u2_u12_u0_U56 (.A( u2_u12_X_1 ) , .ZN( u2_u12_u0_n164 ) );
  INV_X1 u2_u12_u0_U57 (.A( u2_u12_X_3 ) , .ZN( u2_u12_u0_n162 ) );
  INV_X1 u2_u12_u0_U58 (.A( u2_u12_u0_n126 ) , .ZN( u2_u12_u0_n168 ) );
  AOI211_X1 u2_u12_u0_U59 (.B( u2_u12_u0_n133 ) , .A( u2_u12_u0_n134 ) , .C2( u2_u12_u0_n135 ) , .C1( u2_u12_u0_n136 ) , .ZN( u2_u12_u0_n137 ) );
  AOI21_X1 u2_u12_u0_U6 (.B2( u2_u12_u0_n131 ) , .ZN( u2_u12_u0_n134 ) , .B1( u2_u12_u0_n151 ) , .A( u2_u12_u0_n158 ) );
  OR4_X1 u2_u12_u0_U60 (.ZN( u2_out12_17 ) , .A4( u2_u12_u0_n122 ) , .A2( u2_u12_u0_n123 ) , .A1( u2_u12_u0_n124 ) , .A3( u2_u12_u0_n170 ) );
  AOI21_X1 u2_u12_u0_U61 (.B2( u2_u12_u0_n107 ) , .ZN( u2_u12_u0_n124 ) , .B1( u2_u12_u0_n128 ) , .A( u2_u12_u0_n161 ) );
  INV_X1 u2_u12_u0_U62 (.A( u2_u12_u0_n111 ) , .ZN( u2_u12_u0_n170 ) );
  OR4_X1 u2_u12_u0_U63 (.ZN( u2_out12_31 ) , .A4( u2_u12_u0_n155 ) , .A2( u2_u12_u0_n156 ) , .A1( u2_u12_u0_n157 ) , .A3( u2_u12_u0_n173 ) );
  AOI21_X1 u2_u12_u0_U64 (.A( u2_u12_u0_n138 ) , .B2( u2_u12_u0_n139 ) , .B1( u2_u12_u0_n140 ) , .ZN( u2_u12_u0_n157 ) );
  INV_X1 u2_u12_u0_U65 (.ZN( u2_u12_u0_n174 ) , .A( u2_u12_u0_n89 ) );
  AOI211_X1 u2_u12_u0_U66 (.B( u2_u12_u0_n104 ) , .A( u2_u12_u0_n105 ) , .ZN( u2_u12_u0_n106 ) , .C2( u2_u12_u0_n113 ) , .C1( u2_u12_u0_n160 ) );
  AOI21_X1 u2_u12_u0_U67 (.B2( u2_u12_u0_n141 ) , .B1( u2_u12_u0_n142 ) , .ZN( u2_u12_u0_n156 ) , .A( u2_u12_u0_n161 ) );
  AOI21_X1 u2_u12_u0_U68 (.ZN( u2_u12_u0_n116 ) , .B2( u2_u12_u0_n142 ) , .A( u2_u12_u0_n144 ) , .B1( u2_u12_u0_n166 ) );
  INV_X1 u2_u12_u0_U69 (.A( u2_u12_u0_n142 ) , .ZN( u2_u12_u0_n165 ) );
  OAI21_X1 u2_u12_u0_U7 (.B1( u2_u12_u0_n150 ) , .B2( u2_u12_u0_n158 ) , .A( u2_u12_u0_n172 ) , .ZN( u2_u12_u0_n89 ) );
  NAND2_X1 u2_u12_u0_U70 (.A2( u2_u12_u0_n103 ) , .ZN( u2_u12_u0_n140 ) , .A1( u2_u12_u0_n94 ) );
  NAND2_X1 u2_u12_u0_U71 (.A1( u2_u12_u0_n101 ) , .ZN( u2_u12_u0_n130 ) , .A2( u2_u12_u0_n94 ) );
  NAND2_X1 u2_u12_u0_U72 (.ZN( u2_u12_u0_n108 ) , .A1( u2_u12_u0_n92 ) , .A2( u2_u12_u0_n94 ) );
  AND2_X1 u2_u12_u0_U73 (.A1( u2_u12_X_6 ) , .A2( u2_u12_u0_n162 ) , .ZN( u2_u12_u0_n93 ) );
  NOR2_X1 u2_u12_u0_U74 (.A2( u2_u12_X_6 ) , .ZN( u2_u12_u0_n100 ) , .A1( u2_u12_u0_n162 ) );
  NOR2_X1 u2_u12_u0_U75 (.A2( u2_u12_X_3 ) , .A1( u2_u12_X_6 ) , .ZN( u2_u12_u0_n94 ) );
  OAI221_X1 u2_u12_u0_U76 (.C1( u2_u12_u0_n121 ) , .ZN( u2_u12_u0_n122 ) , .B2( u2_u12_u0_n127 ) , .A( u2_u12_u0_n143 ) , .B1( u2_u12_u0_n144 ) , .C2( u2_u12_u0_n147 ) );
  AOI21_X1 u2_u12_u0_U77 (.B1( u2_u12_u0_n132 ) , .ZN( u2_u12_u0_n133 ) , .A( u2_u12_u0_n144 ) , .B2( u2_u12_u0_n166 ) );
  OAI22_X1 u2_u12_u0_U78 (.ZN( u2_u12_u0_n105 ) , .A2( u2_u12_u0_n132 ) , .B1( u2_u12_u0_n146 ) , .A1( u2_u12_u0_n147 ) , .B2( u2_u12_u0_n161 ) );
  NAND2_X1 u2_u12_u0_U79 (.ZN( u2_u12_u0_n110 ) , .A2( u2_u12_u0_n132 ) , .A1( u2_u12_u0_n145 ) );
  AND2_X1 u2_u12_u0_U8 (.A1( u2_u12_u0_n114 ) , .A2( u2_u12_u0_n121 ) , .ZN( u2_u12_u0_n146 ) );
  INV_X1 u2_u12_u0_U80 (.A( u2_u12_u0_n119 ) , .ZN( u2_u12_u0_n167 ) );
  NAND2_X1 u2_u12_u0_U81 (.ZN( u2_u12_u0_n148 ) , .A1( u2_u12_u0_n93 ) , .A2( u2_u12_u0_n95 ) );
  NAND2_X1 u2_u12_u0_U82 (.A1( u2_u12_u0_n100 ) , .ZN( u2_u12_u0_n129 ) , .A2( u2_u12_u0_n95 ) );
  NAND2_X1 u2_u12_u0_U83 (.A1( u2_u12_u0_n102 ) , .ZN( u2_u12_u0_n128 ) , .A2( u2_u12_u0_n95 ) );
  NOR2_X1 u2_u12_u0_U84 (.A2( u2_u12_X_1 ) , .A1( u2_u12_X_2 ) , .ZN( u2_u12_u0_n92 ) );
  NAND2_X1 u2_u12_u0_U85 (.ZN( u2_u12_u0_n142 ) , .A1( u2_u12_u0_n94 ) , .A2( u2_u12_u0_n95 ) );
  NOR2_X1 u2_u12_u0_U86 (.A2( u2_u12_X_2 ) , .ZN( u2_u12_u0_n103 ) , .A1( u2_u12_u0_n164 ) );
  INV_X1 u2_u12_u0_U87 (.A( u2_u12_X_2 ) , .ZN( u2_u12_u0_n163 ) );
  NAND3_X1 u2_u12_u0_U88 (.ZN( u2_out12_23 ) , .A3( u2_u12_u0_n137 ) , .A1( u2_u12_u0_n168 ) , .A2( u2_u12_u0_n171 ) );
  NAND3_X1 u2_u12_u0_U89 (.A3( u2_u12_u0_n127 ) , .A2( u2_u12_u0_n128 ) , .ZN( u2_u12_u0_n135 ) , .A1( u2_u12_u0_n150 ) );
  NAND2_X1 u2_u12_u0_U9 (.ZN( u2_u12_u0_n113 ) , .A1( u2_u12_u0_n139 ) , .A2( u2_u12_u0_n149 ) );
  NAND3_X1 u2_u12_u0_U90 (.ZN( u2_u12_u0_n117 ) , .A3( u2_u12_u0_n132 ) , .A2( u2_u12_u0_n139 ) , .A1( u2_u12_u0_n148 ) );
  NAND3_X1 u2_u12_u0_U91 (.ZN( u2_u12_u0_n109 ) , .A2( u2_u12_u0_n114 ) , .A3( u2_u12_u0_n140 ) , .A1( u2_u12_u0_n149 ) );
  NAND3_X1 u2_u12_u0_U92 (.ZN( u2_out12_9 ) , .A3( u2_u12_u0_n106 ) , .A2( u2_u12_u0_n171 ) , .A1( u2_u12_u0_n174 ) );
  NAND3_X1 u2_u12_u0_U93 (.A2( u2_u12_u0_n128 ) , .A1( u2_u12_u0_n132 ) , .A3( u2_u12_u0_n146 ) , .ZN( u2_u12_u0_n97 ) );
  NOR2_X1 u2_u12_u1_U10 (.A1( u2_u12_u1_n112 ) , .A2( u2_u12_u1_n116 ) , .ZN( u2_u12_u1_n118 ) );
  NAND3_X1 u2_u12_u1_U100 (.ZN( u2_u12_u1_n113 ) , .A1( u2_u12_u1_n120 ) , .A3( u2_u12_u1_n133 ) , .A2( u2_u12_u1_n155 ) );
  OAI21_X1 u2_u12_u1_U11 (.ZN( u2_u12_u1_n101 ) , .B1( u2_u12_u1_n141 ) , .A( u2_u12_u1_n146 ) , .B2( u2_u12_u1_n183 ) );
  AOI21_X1 u2_u12_u1_U12 (.B2( u2_u12_u1_n155 ) , .B1( u2_u12_u1_n156 ) , .ZN( u2_u12_u1_n157 ) , .A( u2_u12_u1_n174 ) );
  NAND2_X1 u2_u12_u1_U13 (.ZN( u2_u12_u1_n140 ) , .A2( u2_u12_u1_n150 ) , .A1( u2_u12_u1_n155 ) );
  NAND2_X1 u2_u12_u1_U14 (.A1( u2_u12_u1_n131 ) , .ZN( u2_u12_u1_n147 ) , .A2( u2_u12_u1_n153 ) );
  INV_X1 u2_u12_u1_U15 (.A( u2_u12_u1_n139 ) , .ZN( u2_u12_u1_n174 ) );
  INV_X1 u2_u12_u1_U16 (.A( u2_u12_u1_n112 ) , .ZN( u2_u12_u1_n171 ) );
  NAND2_X1 u2_u12_u1_U17 (.ZN( u2_u12_u1_n141 ) , .A1( u2_u12_u1_n153 ) , .A2( u2_u12_u1_n156 ) );
  AND2_X1 u2_u12_u1_U18 (.A1( u2_u12_u1_n123 ) , .ZN( u2_u12_u1_n134 ) , .A2( u2_u12_u1_n161 ) );
  NAND2_X1 u2_u12_u1_U19 (.A2( u2_u12_u1_n115 ) , .A1( u2_u12_u1_n116 ) , .ZN( u2_u12_u1_n148 ) );
  NAND2_X1 u2_u12_u1_U20 (.A2( u2_u12_u1_n133 ) , .A1( u2_u12_u1_n135 ) , .ZN( u2_u12_u1_n159 ) );
  NAND2_X1 u2_u12_u1_U21 (.A2( u2_u12_u1_n115 ) , .A1( u2_u12_u1_n120 ) , .ZN( u2_u12_u1_n132 ) );
  INV_X1 u2_u12_u1_U22 (.A( u2_u12_u1_n154 ) , .ZN( u2_u12_u1_n178 ) );
  INV_X1 u2_u12_u1_U23 (.A( u2_u12_u1_n151 ) , .ZN( u2_u12_u1_n183 ) );
  AND2_X1 u2_u12_u1_U24 (.A1( u2_u12_u1_n129 ) , .A2( u2_u12_u1_n133 ) , .ZN( u2_u12_u1_n149 ) );
  INV_X1 u2_u12_u1_U25 (.A( u2_u12_u1_n131 ) , .ZN( u2_u12_u1_n180 ) );
  OR4_X1 u2_u12_u1_U26 (.A4( u2_u12_u1_n106 ) , .A3( u2_u12_u1_n107 ) , .ZN( u2_u12_u1_n108 ) , .A1( u2_u12_u1_n117 ) , .A2( u2_u12_u1_n184 ) );
  AOI21_X1 u2_u12_u1_U27 (.ZN( u2_u12_u1_n106 ) , .A( u2_u12_u1_n112 ) , .B1( u2_u12_u1_n154 ) , .B2( u2_u12_u1_n156 ) );
  AOI21_X1 u2_u12_u1_U28 (.ZN( u2_u12_u1_n107 ) , .B1( u2_u12_u1_n134 ) , .B2( u2_u12_u1_n149 ) , .A( u2_u12_u1_n174 ) );
  INV_X1 u2_u12_u1_U29 (.A( u2_u12_u1_n101 ) , .ZN( u2_u12_u1_n184 ) );
  INV_X1 u2_u12_u1_U3 (.A( u2_u12_u1_n159 ) , .ZN( u2_u12_u1_n182 ) );
  AOI221_X1 u2_u12_u1_U30 (.B1( u2_u12_u1_n140 ) , .ZN( u2_u12_u1_n167 ) , .B2( u2_u12_u1_n172 ) , .C2( u2_u12_u1_n175 ) , .C1( u2_u12_u1_n178 ) , .A( u2_u12_u1_n188 ) );
  INV_X1 u2_u12_u1_U31 (.ZN( u2_u12_u1_n188 ) , .A( u2_u12_u1_n97 ) );
  AOI211_X1 u2_u12_u1_U32 (.A( u2_u12_u1_n118 ) , .C1( u2_u12_u1_n132 ) , .C2( u2_u12_u1_n139 ) , .B( u2_u12_u1_n96 ) , .ZN( u2_u12_u1_n97 ) );
  AOI21_X1 u2_u12_u1_U33 (.B2( u2_u12_u1_n121 ) , .B1( u2_u12_u1_n135 ) , .A( u2_u12_u1_n152 ) , .ZN( u2_u12_u1_n96 ) );
  OAI221_X1 u2_u12_u1_U34 (.A( u2_u12_u1_n119 ) , .C2( u2_u12_u1_n129 ) , .ZN( u2_u12_u1_n138 ) , .B2( u2_u12_u1_n152 ) , .C1( u2_u12_u1_n174 ) , .B1( u2_u12_u1_n187 ) );
  INV_X1 u2_u12_u1_U35 (.A( u2_u12_u1_n148 ) , .ZN( u2_u12_u1_n187 ) );
  AOI211_X1 u2_u12_u1_U36 (.B( u2_u12_u1_n117 ) , .A( u2_u12_u1_n118 ) , .ZN( u2_u12_u1_n119 ) , .C2( u2_u12_u1_n146 ) , .C1( u2_u12_u1_n159 ) );
  NOR2_X1 u2_u12_u1_U37 (.A1( u2_u12_u1_n168 ) , .A2( u2_u12_u1_n176 ) , .ZN( u2_u12_u1_n98 ) );
  AOI211_X1 u2_u12_u1_U38 (.B( u2_u12_u1_n162 ) , .A( u2_u12_u1_n163 ) , .C2( u2_u12_u1_n164 ) , .ZN( u2_u12_u1_n165 ) , .C1( u2_u12_u1_n171 ) );
  AOI21_X1 u2_u12_u1_U39 (.A( u2_u12_u1_n160 ) , .B2( u2_u12_u1_n161 ) , .ZN( u2_u12_u1_n162 ) , .B1( u2_u12_u1_n182 ) );
  AOI221_X1 u2_u12_u1_U4 (.A( u2_u12_u1_n138 ) , .C2( u2_u12_u1_n139 ) , .C1( u2_u12_u1_n140 ) , .B2( u2_u12_u1_n141 ) , .ZN( u2_u12_u1_n142 ) , .B1( u2_u12_u1_n175 ) );
  OR2_X1 u2_u12_u1_U40 (.A2( u2_u12_u1_n157 ) , .A1( u2_u12_u1_n158 ) , .ZN( u2_u12_u1_n163 ) );
  NAND2_X1 u2_u12_u1_U41 (.A1( u2_u12_u1_n128 ) , .ZN( u2_u12_u1_n146 ) , .A2( u2_u12_u1_n160 ) );
  NAND2_X1 u2_u12_u1_U42 (.A2( u2_u12_u1_n112 ) , .ZN( u2_u12_u1_n139 ) , .A1( u2_u12_u1_n152 ) );
  NAND2_X1 u2_u12_u1_U43 (.A1( u2_u12_u1_n105 ) , .ZN( u2_u12_u1_n156 ) , .A2( u2_u12_u1_n99 ) );
  NOR2_X1 u2_u12_u1_U44 (.ZN( u2_u12_u1_n117 ) , .A1( u2_u12_u1_n121 ) , .A2( u2_u12_u1_n160 ) );
  OAI21_X1 u2_u12_u1_U45 (.B2( u2_u12_u1_n123 ) , .ZN( u2_u12_u1_n145 ) , .B1( u2_u12_u1_n160 ) , .A( u2_u12_u1_n185 ) );
  INV_X1 u2_u12_u1_U46 (.A( u2_u12_u1_n122 ) , .ZN( u2_u12_u1_n185 ) );
  AOI21_X1 u2_u12_u1_U47 (.B2( u2_u12_u1_n120 ) , .B1( u2_u12_u1_n121 ) , .ZN( u2_u12_u1_n122 ) , .A( u2_u12_u1_n128 ) );
  AOI21_X1 u2_u12_u1_U48 (.A( u2_u12_u1_n128 ) , .B2( u2_u12_u1_n129 ) , .ZN( u2_u12_u1_n130 ) , .B1( u2_u12_u1_n150 ) );
  NAND2_X1 u2_u12_u1_U49 (.ZN( u2_u12_u1_n112 ) , .A1( u2_u12_u1_n169 ) , .A2( u2_u12_u1_n170 ) );
  AOI211_X1 u2_u12_u1_U5 (.ZN( u2_u12_u1_n124 ) , .A( u2_u12_u1_n138 ) , .C2( u2_u12_u1_n139 ) , .B( u2_u12_u1_n145 ) , .C1( u2_u12_u1_n147 ) );
  NAND2_X1 u2_u12_u1_U50 (.ZN( u2_u12_u1_n129 ) , .A2( u2_u12_u1_n95 ) , .A1( u2_u12_u1_n98 ) );
  NAND2_X1 u2_u12_u1_U51 (.A1( u2_u12_u1_n102 ) , .ZN( u2_u12_u1_n154 ) , .A2( u2_u12_u1_n99 ) );
  NAND2_X1 u2_u12_u1_U52 (.A2( u2_u12_u1_n100 ) , .ZN( u2_u12_u1_n135 ) , .A1( u2_u12_u1_n99 ) );
  AOI21_X1 u2_u12_u1_U53 (.A( u2_u12_u1_n152 ) , .B2( u2_u12_u1_n153 ) , .B1( u2_u12_u1_n154 ) , .ZN( u2_u12_u1_n158 ) );
  INV_X1 u2_u12_u1_U54 (.A( u2_u12_u1_n160 ) , .ZN( u2_u12_u1_n175 ) );
  NAND2_X1 u2_u12_u1_U55 (.A1( u2_u12_u1_n100 ) , .ZN( u2_u12_u1_n116 ) , .A2( u2_u12_u1_n95 ) );
  NAND2_X1 u2_u12_u1_U56 (.A1( u2_u12_u1_n102 ) , .ZN( u2_u12_u1_n131 ) , .A2( u2_u12_u1_n95 ) );
  NAND2_X1 u2_u12_u1_U57 (.A2( u2_u12_u1_n104 ) , .ZN( u2_u12_u1_n121 ) , .A1( u2_u12_u1_n98 ) );
  NAND2_X1 u2_u12_u1_U58 (.A1( u2_u12_u1_n103 ) , .ZN( u2_u12_u1_n153 ) , .A2( u2_u12_u1_n98 ) );
  NAND2_X1 u2_u12_u1_U59 (.A2( u2_u12_u1_n104 ) , .A1( u2_u12_u1_n105 ) , .ZN( u2_u12_u1_n133 ) );
  AOI22_X1 u2_u12_u1_U6 (.B2( u2_u12_u1_n113 ) , .A2( u2_u12_u1_n114 ) , .ZN( u2_u12_u1_n125 ) , .A1( u2_u12_u1_n171 ) , .B1( u2_u12_u1_n173 ) );
  NAND2_X1 u2_u12_u1_U60 (.ZN( u2_u12_u1_n150 ) , .A2( u2_u12_u1_n98 ) , .A1( u2_u12_u1_n99 ) );
  NAND2_X1 u2_u12_u1_U61 (.A1( u2_u12_u1_n105 ) , .ZN( u2_u12_u1_n155 ) , .A2( u2_u12_u1_n95 ) );
  OAI21_X1 u2_u12_u1_U62 (.ZN( u2_u12_u1_n109 ) , .B1( u2_u12_u1_n129 ) , .B2( u2_u12_u1_n160 ) , .A( u2_u12_u1_n167 ) );
  NAND2_X1 u2_u12_u1_U63 (.A2( u2_u12_u1_n100 ) , .A1( u2_u12_u1_n103 ) , .ZN( u2_u12_u1_n120 ) );
  NAND2_X1 u2_u12_u1_U64 (.A1( u2_u12_u1_n102 ) , .A2( u2_u12_u1_n104 ) , .ZN( u2_u12_u1_n115 ) );
  NAND2_X1 u2_u12_u1_U65 (.A2( u2_u12_u1_n100 ) , .A1( u2_u12_u1_n104 ) , .ZN( u2_u12_u1_n151 ) );
  NAND2_X1 u2_u12_u1_U66 (.A2( u2_u12_u1_n103 ) , .A1( u2_u12_u1_n105 ) , .ZN( u2_u12_u1_n161 ) );
  INV_X1 u2_u12_u1_U67 (.A( u2_u12_u1_n152 ) , .ZN( u2_u12_u1_n173 ) );
  INV_X1 u2_u12_u1_U68 (.A( u2_u12_u1_n128 ) , .ZN( u2_u12_u1_n172 ) );
  NAND2_X1 u2_u12_u1_U69 (.A2( u2_u12_u1_n102 ) , .A1( u2_u12_u1_n103 ) , .ZN( u2_u12_u1_n123 ) );
  NAND2_X1 u2_u12_u1_U7 (.ZN( u2_u12_u1_n114 ) , .A1( u2_u12_u1_n134 ) , .A2( u2_u12_u1_n156 ) );
  NOR2_X1 u2_u12_u1_U70 (.A2( u2_u12_X_7 ) , .A1( u2_u12_X_8 ) , .ZN( u2_u12_u1_n95 ) );
  NOR2_X1 u2_u12_u1_U71 (.A1( u2_u12_X_12 ) , .A2( u2_u12_X_9 ) , .ZN( u2_u12_u1_n100 ) );
  NOR2_X1 u2_u12_u1_U72 (.A2( u2_u12_X_8 ) , .A1( u2_u12_u1_n177 ) , .ZN( u2_u12_u1_n99 ) );
  NOR2_X1 u2_u12_u1_U73 (.A2( u2_u12_X_12 ) , .ZN( u2_u12_u1_n102 ) , .A1( u2_u12_u1_n176 ) );
  NOR2_X1 u2_u12_u1_U74 (.A2( u2_u12_X_9 ) , .ZN( u2_u12_u1_n105 ) , .A1( u2_u12_u1_n168 ) );
  NAND2_X1 u2_u12_u1_U75 (.A1( u2_u12_X_10 ) , .ZN( u2_u12_u1_n160 ) , .A2( u2_u12_u1_n169 ) );
  NAND2_X1 u2_u12_u1_U76 (.A2( u2_u12_X_10 ) , .A1( u2_u12_X_11 ) , .ZN( u2_u12_u1_n152 ) );
  NAND2_X1 u2_u12_u1_U77 (.A1( u2_u12_X_11 ) , .ZN( u2_u12_u1_n128 ) , .A2( u2_u12_u1_n170 ) );
  AND2_X1 u2_u12_u1_U78 (.A2( u2_u12_X_7 ) , .A1( u2_u12_X_8 ) , .ZN( u2_u12_u1_n104 ) );
  AND2_X1 u2_u12_u1_U79 (.A1( u2_u12_X_8 ) , .ZN( u2_u12_u1_n103 ) , .A2( u2_u12_u1_n177 ) );
  AOI22_X1 u2_u12_u1_U8 (.B2( u2_u12_u1_n136 ) , .A2( u2_u12_u1_n137 ) , .ZN( u2_u12_u1_n143 ) , .A1( u2_u12_u1_n171 ) , .B1( u2_u12_u1_n173 ) );
  INV_X1 u2_u12_u1_U80 (.A( u2_u12_X_10 ) , .ZN( u2_u12_u1_n170 ) );
  INV_X1 u2_u12_u1_U81 (.A( u2_u12_X_9 ) , .ZN( u2_u12_u1_n176 ) );
  INV_X1 u2_u12_u1_U82 (.A( u2_u12_X_11 ) , .ZN( u2_u12_u1_n169 ) );
  INV_X1 u2_u12_u1_U83 (.A( u2_u12_X_12 ) , .ZN( u2_u12_u1_n168 ) );
  INV_X1 u2_u12_u1_U84 (.A( u2_u12_X_7 ) , .ZN( u2_u12_u1_n177 ) );
  NAND4_X1 u2_u12_u1_U85 (.ZN( u2_out12_28 ) , .A4( u2_u12_u1_n124 ) , .A3( u2_u12_u1_n125 ) , .A2( u2_u12_u1_n126 ) , .A1( u2_u12_u1_n127 ) );
  OAI21_X1 u2_u12_u1_U86 (.ZN( u2_u12_u1_n127 ) , .B2( u2_u12_u1_n139 ) , .B1( u2_u12_u1_n175 ) , .A( u2_u12_u1_n183 ) );
  OAI21_X1 u2_u12_u1_U87 (.ZN( u2_u12_u1_n126 ) , .B2( u2_u12_u1_n140 ) , .A( u2_u12_u1_n146 ) , .B1( u2_u12_u1_n178 ) );
  NAND4_X1 u2_u12_u1_U88 (.ZN( u2_out12_18 ) , .A4( u2_u12_u1_n165 ) , .A3( u2_u12_u1_n166 ) , .A1( u2_u12_u1_n167 ) , .A2( u2_u12_u1_n186 ) );
  AOI22_X1 u2_u12_u1_U89 (.B2( u2_u12_u1_n146 ) , .B1( u2_u12_u1_n147 ) , .A2( u2_u12_u1_n148 ) , .ZN( u2_u12_u1_n166 ) , .A1( u2_u12_u1_n172 ) );
  INV_X1 u2_u12_u1_U9 (.A( u2_u12_u1_n147 ) , .ZN( u2_u12_u1_n181 ) );
  INV_X1 u2_u12_u1_U90 (.A( u2_u12_u1_n145 ) , .ZN( u2_u12_u1_n186 ) );
  NAND4_X1 u2_u12_u1_U91 (.ZN( u2_out12_2 ) , .A4( u2_u12_u1_n142 ) , .A3( u2_u12_u1_n143 ) , .A2( u2_u12_u1_n144 ) , .A1( u2_u12_u1_n179 ) );
  OAI21_X1 u2_u12_u1_U92 (.B2( u2_u12_u1_n132 ) , .ZN( u2_u12_u1_n144 ) , .A( u2_u12_u1_n146 ) , .B1( u2_u12_u1_n180 ) );
  INV_X1 u2_u12_u1_U93 (.A( u2_u12_u1_n130 ) , .ZN( u2_u12_u1_n179 ) );
  OR4_X1 u2_u12_u1_U94 (.ZN( u2_out12_13 ) , .A4( u2_u12_u1_n108 ) , .A3( u2_u12_u1_n109 ) , .A2( u2_u12_u1_n110 ) , .A1( u2_u12_u1_n111 ) );
  AOI21_X1 u2_u12_u1_U95 (.ZN( u2_u12_u1_n111 ) , .A( u2_u12_u1_n128 ) , .B2( u2_u12_u1_n131 ) , .B1( u2_u12_u1_n135 ) );
  AOI21_X1 u2_u12_u1_U96 (.ZN( u2_u12_u1_n110 ) , .A( u2_u12_u1_n116 ) , .B1( u2_u12_u1_n152 ) , .B2( u2_u12_u1_n160 ) );
  NAND3_X1 u2_u12_u1_U97 (.A3( u2_u12_u1_n149 ) , .A2( u2_u12_u1_n150 ) , .A1( u2_u12_u1_n151 ) , .ZN( u2_u12_u1_n164 ) );
  NAND3_X1 u2_u12_u1_U98 (.A3( u2_u12_u1_n134 ) , .A2( u2_u12_u1_n135 ) , .ZN( u2_u12_u1_n136 ) , .A1( u2_u12_u1_n151 ) );
  NAND3_X1 u2_u12_u1_U99 (.A1( u2_u12_u1_n133 ) , .ZN( u2_u12_u1_n137 ) , .A2( u2_u12_u1_n154 ) , .A3( u2_u12_u1_n181 ) );
  OAI22_X1 u2_u12_u2_U10 (.B1( u2_u12_u2_n151 ) , .A2( u2_u12_u2_n152 ) , .A1( u2_u12_u2_n153 ) , .ZN( u2_u12_u2_n160 ) , .B2( u2_u12_u2_n168 ) );
  NAND3_X1 u2_u12_u2_U100 (.A2( u2_u12_u2_n100 ) , .A1( u2_u12_u2_n104 ) , .A3( u2_u12_u2_n138 ) , .ZN( u2_u12_u2_n98 ) );
  NOR3_X1 u2_u12_u2_U11 (.A1( u2_u12_u2_n150 ) , .ZN( u2_u12_u2_n151 ) , .A3( u2_u12_u2_n175 ) , .A2( u2_u12_u2_n188 ) );
  AOI21_X1 u2_u12_u2_U12 (.B2( u2_u12_u2_n123 ) , .ZN( u2_u12_u2_n125 ) , .A( u2_u12_u2_n171 ) , .B1( u2_u12_u2_n184 ) );
  INV_X1 u2_u12_u2_U13 (.A( u2_u12_u2_n150 ) , .ZN( u2_u12_u2_n184 ) );
  AOI21_X1 u2_u12_u2_U14 (.ZN( u2_u12_u2_n144 ) , .B2( u2_u12_u2_n155 ) , .A( u2_u12_u2_n172 ) , .B1( u2_u12_u2_n185 ) );
  AOI21_X1 u2_u12_u2_U15 (.B2( u2_u12_u2_n143 ) , .ZN( u2_u12_u2_n145 ) , .B1( u2_u12_u2_n152 ) , .A( u2_u12_u2_n171 ) );
  INV_X1 u2_u12_u2_U16 (.A( u2_u12_u2_n156 ) , .ZN( u2_u12_u2_n171 ) );
  INV_X1 u2_u12_u2_U17 (.A( u2_u12_u2_n120 ) , .ZN( u2_u12_u2_n188 ) );
  NAND2_X1 u2_u12_u2_U18 (.A2( u2_u12_u2_n122 ) , .ZN( u2_u12_u2_n150 ) , .A1( u2_u12_u2_n152 ) );
  INV_X1 u2_u12_u2_U19 (.A( u2_u12_u2_n153 ) , .ZN( u2_u12_u2_n170 ) );
  INV_X1 u2_u12_u2_U20 (.A( u2_u12_u2_n137 ) , .ZN( u2_u12_u2_n173 ) );
  NAND2_X1 u2_u12_u2_U21 (.A1( u2_u12_u2_n132 ) , .A2( u2_u12_u2_n139 ) , .ZN( u2_u12_u2_n157 ) );
  INV_X1 u2_u12_u2_U22 (.A( u2_u12_u2_n113 ) , .ZN( u2_u12_u2_n178 ) );
  INV_X1 u2_u12_u2_U23 (.A( u2_u12_u2_n139 ) , .ZN( u2_u12_u2_n175 ) );
  INV_X1 u2_u12_u2_U24 (.A( u2_u12_u2_n155 ) , .ZN( u2_u12_u2_n181 ) );
  INV_X1 u2_u12_u2_U25 (.A( u2_u12_u2_n119 ) , .ZN( u2_u12_u2_n177 ) );
  INV_X1 u2_u12_u2_U26 (.A( u2_u12_u2_n116 ) , .ZN( u2_u12_u2_n180 ) );
  INV_X1 u2_u12_u2_U27 (.A( u2_u12_u2_n131 ) , .ZN( u2_u12_u2_n179 ) );
  INV_X1 u2_u12_u2_U28 (.A( u2_u12_u2_n154 ) , .ZN( u2_u12_u2_n176 ) );
  NAND2_X1 u2_u12_u2_U29 (.A2( u2_u12_u2_n116 ) , .A1( u2_u12_u2_n117 ) , .ZN( u2_u12_u2_n118 ) );
  NOR2_X1 u2_u12_u2_U3 (.ZN( u2_u12_u2_n121 ) , .A2( u2_u12_u2_n177 ) , .A1( u2_u12_u2_n180 ) );
  INV_X1 u2_u12_u2_U30 (.A( u2_u12_u2_n132 ) , .ZN( u2_u12_u2_n182 ) );
  INV_X1 u2_u12_u2_U31 (.A( u2_u12_u2_n158 ) , .ZN( u2_u12_u2_n183 ) );
  OAI21_X1 u2_u12_u2_U32 (.A( u2_u12_u2_n156 ) , .B1( u2_u12_u2_n157 ) , .ZN( u2_u12_u2_n158 ) , .B2( u2_u12_u2_n179 ) );
  NOR2_X1 u2_u12_u2_U33 (.ZN( u2_u12_u2_n156 ) , .A1( u2_u12_u2_n166 ) , .A2( u2_u12_u2_n169 ) );
  NOR2_X1 u2_u12_u2_U34 (.A2( u2_u12_u2_n114 ) , .ZN( u2_u12_u2_n137 ) , .A1( u2_u12_u2_n140 ) );
  NOR2_X1 u2_u12_u2_U35 (.A2( u2_u12_u2_n138 ) , .ZN( u2_u12_u2_n153 ) , .A1( u2_u12_u2_n156 ) );
  AOI211_X1 u2_u12_u2_U36 (.ZN( u2_u12_u2_n130 ) , .C1( u2_u12_u2_n138 ) , .C2( u2_u12_u2_n179 ) , .B( u2_u12_u2_n96 ) , .A( u2_u12_u2_n97 ) );
  OAI22_X1 u2_u12_u2_U37 (.B1( u2_u12_u2_n133 ) , .A2( u2_u12_u2_n137 ) , .A1( u2_u12_u2_n152 ) , .B2( u2_u12_u2_n168 ) , .ZN( u2_u12_u2_n97 ) );
  OAI221_X1 u2_u12_u2_U38 (.B1( u2_u12_u2_n113 ) , .C1( u2_u12_u2_n132 ) , .A( u2_u12_u2_n149 ) , .B2( u2_u12_u2_n171 ) , .C2( u2_u12_u2_n172 ) , .ZN( u2_u12_u2_n96 ) );
  OAI221_X1 u2_u12_u2_U39 (.A( u2_u12_u2_n115 ) , .C2( u2_u12_u2_n123 ) , .B2( u2_u12_u2_n143 ) , .B1( u2_u12_u2_n153 ) , .ZN( u2_u12_u2_n163 ) , .C1( u2_u12_u2_n168 ) );
  INV_X1 u2_u12_u2_U4 (.A( u2_u12_u2_n134 ) , .ZN( u2_u12_u2_n185 ) );
  OAI21_X1 u2_u12_u2_U40 (.A( u2_u12_u2_n114 ) , .ZN( u2_u12_u2_n115 ) , .B1( u2_u12_u2_n176 ) , .B2( u2_u12_u2_n178 ) );
  OAI221_X1 u2_u12_u2_U41 (.A( u2_u12_u2_n135 ) , .B2( u2_u12_u2_n136 ) , .B1( u2_u12_u2_n137 ) , .ZN( u2_u12_u2_n162 ) , .C2( u2_u12_u2_n167 ) , .C1( u2_u12_u2_n185 ) );
  AND3_X1 u2_u12_u2_U42 (.A3( u2_u12_u2_n131 ) , .A2( u2_u12_u2_n132 ) , .A1( u2_u12_u2_n133 ) , .ZN( u2_u12_u2_n136 ) );
  AOI22_X1 u2_u12_u2_U43 (.ZN( u2_u12_u2_n135 ) , .B1( u2_u12_u2_n140 ) , .A1( u2_u12_u2_n156 ) , .B2( u2_u12_u2_n180 ) , .A2( u2_u12_u2_n188 ) );
  AOI21_X1 u2_u12_u2_U44 (.ZN( u2_u12_u2_n149 ) , .B1( u2_u12_u2_n173 ) , .B2( u2_u12_u2_n188 ) , .A( u2_u12_u2_n95 ) );
  AND3_X1 u2_u12_u2_U45 (.A2( u2_u12_u2_n100 ) , .A1( u2_u12_u2_n104 ) , .A3( u2_u12_u2_n156 ) , .ZN( u2_u12_u2_n95 ) );
  OAI21_X1 u2_u12_u2_U46 (.A( u2_u12_u2_n101 ) , .B2( u2_u12_u2_n121 ) , .B1( u2_u12_u2_n153 ) , .ZN( u2_u12_u2_n164 ) );
  NAND2_X1 u2_u12_u2_U47 (.A2( u2_u12_u2_n100 ) , .A1( u2_u12_u2_n107 ) , .ZN( u2_u12_u2_n155 ) );
  NAND2_X1 u2_u12_u2_U48 (.A2( u2_u12_u2_n105 ) , .A1( u2_u12_u2_n108 ) , .ZN( u2_u12_u2_n143 ) );
  NAND2_X1 u2_u12_u2_U49 (.A1( u2_u12_u2_n104 ) , .A2( u2_u12_u2_n106 ) , .ZN( u2_u12_u2_n152 ) );
  NOR4_X1 u2_u12_u2_U5 (.A4( u2_u12_u2_n124 ) , .A3( u2_u12_u2_n125 ) , .A2( u2_u12_u2_n126 ) , .A1( u2_u12_u2_n127 ) , .ZN( u2_u12_u2_n128 ) );
  NAND2_X1 u2_u12_u2_U50 (.A1( u2_u12_u2_n100 ) , .A2( u2_u12_u2_n105 ) , .ZN( u2_u12_u2_n132 ) );
  INV_X1 u2_u12_u2_U51 (.A( u2_u12_u2_n140 ) , .ZN( u2_u12_u2_n168 ) );
  INV_X1 u2_u12_u2_U52 (.A( u2_u12_u2_n138 ) , .ZN( u2_u12_u2_n167 ) );
  OAI21_X1 u2_u12_u2_U53 (.A( u2_u12_u2_n141 ) , .B2( u2_u12_u2_n142 ) , .ZN( u2_u12_u2_n146 ) , .B1( u2_u12_u2_n153 ) );
  OAI21_X1 u2_u12_u2_U54 (.A( u2_u12_u2_n140 ) , .ZN( u2_u12_u2_n141 ) , .B1( u2_u12_u2_n176 ) , .B2( u2_u12_u2_n177 ) );
  NOR3_X1 u2_u12_u2_U55 (.ZN( u2_u12_u2_n142 ) , .A3( u2_u12_u2_n175 ) , .A2( u2_u12_u2_n178 ) , .A1( u2_u12_u2_n181 ) );
  NAND2_X1 u2_u12_u2_U56 (.A1( u2_u12_u2_n102 ) , .A2( u2_u12_u2_n106 ) , .ZN( u2_u12_u2_n113 ) );
  NAND2_X1 u2_u12_u2_U57 (.A1( u2_u12_u2_n106 ) , .A2( u2_u12_u2_n107 ) , .ZN( u2_u12_u2_n131 ) );
  NAND2_X1 u2_u12_u2_U58 (.A1( u2_u12_u2_n103 ) , .A2( u2_u12_u2_n107 ) , .ZN( u2_u12_u2_n139 ) );
  NAND2_X1 u2_u12_u2_U59 (.A1( u2_u12_u2_n103 ) , .A2( u2_u12_u2_n105 ) , .ZN( u2_u12_u2_n133 ) );
  AOI21_X1 u2_u12_u2_U6 (.B2( u2_u12_u2_n119 ) , .ZN( u2_u12_u2_n127 ) , .A( u2_u12_u2_n137 ) , .B1( u2_u12_u2_n155 ) );
  NAND2_X1 u2_u12_u2_U60 (.A1( u2_u12_u2_n102 ) , .A2( u2_u12_u2_n103 ) , .ZN( u2_u12_u2_n154 ) );
  NAND2_X1 u2_u12_u2_U61 (.A2( u2_u12_u2_n103 ) , .A1( u2_u12_u2_n104 ) , .ZN( u2_u12_u2_n119 ) );
  NAND2_X1 u2_u12_u2_U62 (.A2( u2_u12_u2_n107 ) , .A1( u2_u12_u2_n108 ) , .ZN( u2_u12_u2_n123 ) );
  NAND2_X1 u2_u12_u2_U63 (.A1( u2_u12_u2_n104 ) , .A2( u2_u12_u2_n108 ) , .ZN( u2_u12_u2_n122 ) );
  INV_X1 u2_u12_u2_U64 (.A( u2_u12_u2_n114 ) , .ZN( u2_u12_u2_n172 ) );
  NAND2_X1 u2_u12_u2_U65 (.A2( u2_u12_u2_n100 ) , .A1( u2_u12_u2_n102 ) , .ZN( u2_u12_u2_n116 ) );
  NAND2_X1 u2_u12_u2_U66 (.A1( u2_u12_u2_n102 ) , .A2( u2_u12_u2_n108 ) , .ZN( u2_u12_u2_n120 ) );
  NAND2_X1 u2_u12_u2_U67 (.A2( u2_u12_u2_n105 ) , .A1( u2_u12_u2_n106 ) , .ZN( u2_u12_u2_n117 ) );
  INV_X1 u2_u12_u2_U68 (.ZN( u2_u12_u2_n187 ) , .A( u2_u12_u2_n99 ) );
  OAI21_X1 u2_u12_u2_U69 (.B1( u2_u12_u2_n137 ) , .B2( u2_u12_u2_n143 ) , .A( u2_u12_u2_n98 ) , .ZN( u2_u12_u2_n99 ) );
  AOI21_X1 u2_u12_u2_U7 (.ZN( u2_u12_u2_n124 ) , .B1( u2_u12_u2_n131 ) , .B2( u2_u12_u2_n143 ) , .A( u2_u12_u2_n172 ) );
  NOR2_X1 u2_u12_u2_U70 (.A2( u2_u12_X_16 ) , .ZN( u2_u12_u2_n140 ) , .A1( u2_u12_u2_n166 ) );
  NOR2_X1 u2_u12_u2_U71 (.A2( u2_u12_X_13 ) , .A1( u2_u12_X_14 ) , .ZN( u2_u12_u2_n100 ) );
  NOR2_X1 u2_u12_u2_U72 (.A2( u2_u12_X_16 ) , .A1( u2_u12_X_17 ) , .ZN( u2_u12_u2_n138 ) );
  NOR2_X1 u2_u12_u2_U73 (.A2( u2_u12_X_15 ) , .A1( u2_u12_X_18 ) , .ZN( u2_u12_u2_n104 ) );
  NOR2_X1 u2_u12_u2_U74 (.A2( u2_u12_X_14 ) , .ZN( u2_u12_u2_n103 ) , .A1( u2_u12_u2_n174 ) );
  NOR2_X1 u2_u12_u2_U75 (.A2( u2_u12_X_15 ) , .ZN( u2_u12_u2_n102 ) , .A1( u2_u12_u2_n165 ) );
  NOR2_X1 u2_u12_u2_U76 (.A2( u2_u12_X_17 ) , .ZN( u2_u12_u2_n114 ) , .A1( u2_u12_u2_n169 ) );
  AND2_X1 u2_u12_u2_U77 (.A1( u2_u12_X_15 ) , .ZN( u2_u12_u2_n105 ) , .A2( u2_u12_u2_n165 ) );
  AND2_X1 u2_u12_u2_U78 (.A2( u2_u12_X_15 ) , .A1( u2_u12_X_18 ) , .ZN( u2_u12_u2_n107 ) );
  AND2_X1 u2_u12_u2_U79 (.A1( u2_u12_X_14 ) , .ZN( u2_u12_u2_n106 ) , .A2( u2_u12_u2_n174 ) );
  AOI21_X1 u2_u12_u2_U8 (.B2( u2_u12_u2_n120 ) , .B1( u2_u12_u2_n121 ) , .ZN( u2_u12_u2_n126 ) , .A( u2_u12_u2_n167 ) );
  AND2_X1 u2_u12_u2_U80 (.A1( u2_u12_X_13 ) , .A2( u2_u12_X_14 ) , .ZN( u2_u12_u2_n108 ) );
  INV_X1 u2_u12_u2_U81 (.A( u2_u12_X_16 ) , .ZN( u2_u12_u2_n169 ) );
  INV_X1 u2_u12_u2_U82 (.A( u2_u12_X_17 ) , .ZN( u2_u12_u2_n166 ) );
  INV_X1 u2_u12_u2_U83 (.A( u2_u12_X_13 ) , .ZN( u2_u12_u2_n174 ) );
  INV_X1 u2_u12_u2_U84 (.A( u2_u12_X_18 ) , .ZN( u2_u12_u2_n165 ) );
  NAND4_X1 u2_u12_u2_U85 (.ZN( u2_out12_30 ) , .A4( u2_u12_u2_n147 ) , .A3( u2_u12_u2_n148 ) , .A2( u2_u12_u2_n149 ) , .A1( u2_u12_u2_n187 ) );
  AOI21_X1 u2_u12_u2_U86 (.B2( u2_u12_u2_n138 ) , .ZN( u2_u12_u2_n148 ) , .A( u2_u12_u2_n162 ) , .B1( u2_u12_u2_n182 ) );
  NOR3_X1 u2_u12_u2_U87 (.A3( u2_u12_u2_n144 ) , .A2( u2_u12_u2_n145 ) , .A1( u2_u12_u2_n146 ) , .ZN( u2_u12_u2_n147 ) );
  NAND4_X1 u2_u12_u2_U88 (.ZN( u2_out12_24 ) , .A4( u2_u12_u2_n111 ) , .A3( u2_u12_u2_n112 ) , .A1( u2_u12_u2_n130 ) , .A2( u2_u12_u2_n187 ) );
  AOI221_X1 u2_u12_u2_U89 (.A( u2_u12_u2_n109 ) , .B1( u2_u12_u2_n110 ) , .ZN( u2_u12_u2_n111 ) , .C1( u2_u12_u2_n134 ) , .C2( u2_u12_u2_n170 ) , .B2( u2_u12_u2_n173 ) );
  OAI22_X1 u2_u12_u2_U9 (.ZN( u2_u12_u2_n109 ) , .A2( u2_u12_u2_n113 ) , .B2( u2_u12_u2_n133 ) , .B1( u2_u12_u2_n167 ) , .A1( u2_u12_u2_n168 ) );
  AOI21_X1 u2_u12_u2_U90 (.ZN( u2_u12_u2_n112 ) , .B2( u2_u12_u2_n156 ) , .A( u2_u12_u2_n164 ) , .B1( u2_u12_u2_n181 ) );
  NAND4_X1 u2_u12_u2_U91 (.ZN( u2_out12_16 ) , .A4( u2_u12_u2_n128 ) , .A3( u2_u12_u2_n129 ) , .A1( u2_u12_u2_n130 ) , .A2( u2_u12_u2_n186 ) );
  AOI22_X1 u2_u12_u2_U92 (.A2( u2_u12_u2_n118 ) , .ZN( u2_u12_u2_n129 ) , .A1( u2_u12_u2_n140 ) , .B1( u2_u12_u2_n157 ) , .B2( u2_u12_u2_n170 ) );
  INV_X1 u2_u12_u2_U93 (.A( u2_u12_u2_n163 ) , .ZN( u2_u12_u2_n186 ) );
  OR4_X1 u2_u12_u2_U94 (.ZN( u2_out12_6 ) , .A4( u2_u12_u2_n161 ) , .A3( u2_u12_u2_n162 ) , .A2( u2_u12_u2_n163 ) , .A1( u2_u12_u2_n164 ) );
  OR3_X1 u2_u12_u2_U95 (.A2( u2_u12_u2_n159 ) , .A1( u2_u12_u2_n160 ) , .ZN( u2_u12_u2_n161 ) , .A3( u2_u12_u2_n183 ) );
  AOI21_X1 u2_u12_u2_U96 (.B2( u2_u12_u2_n154 ) , .B1( u2_u12_u2_n155 ) , .ZN( u2_u12_u2_n159 ) , .A( u2_u12_u2_n167 ) );
  NAND3_X1 u2_u12_u2_U97 (.A2( u2_u12_u2_n117 ) , .A1( u2_u12_u2_n122 ) , .A3( u2_u12_u2_n123 ) , .ZN( u2_u12_u2_n134 ) );
  NAND3_X1 u2_u12_u2_U98 (.ZN( u2_u12_u2_n110 ) , .A2( u2_u12_u2_n131 ) , .A3( u2_u12_u2_n139 ) , .A1( u2_u12_u2_n154 ) );
  NAND3_X1 u2_u12_u2_U99 (.A2( u2_u12_u2_n100 ) , .ZN( u2_u12_u2_n101 ) , .A1( u2_u12_u2_n104 ) , .A3( u2_u12_u2_n114 ) );
  AOI22_X1 u2_u12_u6_U10 (.A2( u2_u12_u6_n151 ) , .B2( u2_u12_u6_n161 ) , .A1( u2_u12_u6_n167 ) , .B1( u2_u12_u6_n170 ) , .ZN( u2_u12_u6_n89 ) );
  AOI21_X1 u2_u12_u6_U11 (.B1( u2_u12_u6_n107 ) , .B2( u2_u12_u6_n132 ) , .A( u2_u12_u6_n158 ) , .ZN( u2_u12_u6_n88 ) );
  AOI21_X1 u2_u12_u6_U12 (.B2( u2_u12_u6_n147 ) , .B1( u2_u12_u6_n148 ) , .ZN( u2_u12_u6_n149 ) , .A( u2_u12_u6_n158 ) );
  AOI21_X1 u2_u12_u6_U13 (.ZN( u2_u12_u6_n106 ) , .A( u2_u12_u6_n142 ) , .B2( u2_u12_u6_n159 ) , .B1( u2_u12_u6_n164 ) );
  INV_X1 u2_u12_u6_U14 (.A( u2_u12_u6_n155 ) , .ZN( u2_u12_u6_n161 ) );
  INV_X1 u2_u12_u6_U15 (.A( u2_u12_u6_n128 ) , .ZN( u2_u12_u6_n164 ) );
  NAND2_X1 u2_u12_u6_U16 (.ZN( u2_u12_u6_n110 ) , .A1( u2_u12_u6_n122 ) , .A2( u2_u12_u6_n129 ) );
  NAND2_X1 u2_u12_u6_U17 (.ZN( u2_u12_u6_n124 ) , .A2( u2_u12_u6_n146 ) , .A1( u2_u12_u6_n148 ) );
  INV_X1 u2_u12_u6_U18 (.A( u2_u12_u6_n132 ) , .ZN( u2_u12_u6_n171 ) );
  AND2_X1 u2_u12_u6_U19 (.A1( u2_u12_u6_n100 ) , .ZN( u2_u12_u6_n130 ) , .A2( u2_u12_u6_n147 ) );
  INV_X1 u2_u12_u6_U20 (.A( u2_u12_u6_n127 ) , .ZN( u2_u12_u6_n173 ) );
  INV_X1 u2_u12_u6_U21 (.A( u2_u12_u6_n121 ) , .ZN( u2_u12_u6_n167 ) );
  INV_X1 u2_u12_u6_U22 (.A( u2_u12_u6_n100 ) , .ZN( u2_u12_u6_n169 ) );
  INV_X1 u2_u12_u6_U23 (.A( u2_u12_u6_n123 ) , .ZN( u2_u12_u6_n170 ) );
  INV_X1 u2_u12_u6_U24 (.A( u2_u12_u6_n113 ) , .ZN( u2_u12_u6_n168 ) );
  AND2_X1 u2_u12_u6_U25 (.A1( u2_u12_u6_n107 ) , .A2( u2_u12_u6_n119 ) , .ZN( u2_u12_u6_n133 ) );
  AND2_X1 u2_u12_u6_U26 (.A2( u2_u12_u6_n121 ) , .A1( u2_u12_u6_n122 ) , .ZN( u2_u12_u6_n131 ) );
  AND3_X1 u2_u12_u6_U27 (.ZN( u2_u12_u6_n120 ) , .A2( u2_u12_u6_n127 ) , .A1( u2_u12_u6_n132 ) , .A3( u2_u12_u6_n145 ) );
  INV_X1 u2_u12_u6_U28 (.A( u2_u12_u6_n146 ) , .ZN( u2_u12_u6_n163 ) );
  AOI222_X1 u2_u12_u6_U29 (.ZN( u2_u12_u6_n114 ) , .A1( u2_u12_u6_n118 ) , .A2( u2_u12_u6_n126 ) , .B2( u2_u12_u6_n151 ) , .C2( u2_u12_u6_n159 ) , .C1( u2_u12_u6_n168 ) , .B1( u2_u12_u6_n169 ) );
  INV_X1 u2_u12_u6_U3 (.A( u2_u12_u6_n110 ) , .ZN( u2_u12_u6_n166 ) );
  NOR2_X1 u2_u12_u6_U30 (.A1( u2_u12_u6_n162 ) , .A2( u2_u12_u6_n165 ) , .ZN( u2_u12_u6_n98 ) );
  AOI211_X1 u2_u12_u6_U31 (.B( u2_u12_u6_n134 ) , .A( u2_u12_u6_n135 ) , .C1( u2_u12_u6_n136 ) , .ZN( u2_u12_u6_n137 ) , .C2( u2_u12_u6_n151 ) );
  AOI21_X1 u2_u12_u6_U32 (.B2( u2_u12_u6_n132 ) , .B1( u2_u12_u6_n133 ) , .ZN( u2_u12_u6_n134 ) , .A( u2_u12_u6_n158 ) );
  AOI21_X1 u2_u12_u6_U33 (.B1( u2_u12_u6_n131 ) , .ZN( u2_u12_u6_n135 ) , .A( u2_u12_u6_n144 ) , .B2( u2_u12_u6_n146 ) );
  NAND4_X1 u2_u12_u6_U34 (.A4( u2_u12_u6_n127 ) , .A3( u2_u12_u6_n128 ) , .A2( u2_u12_u6_n129 ) , .A1( u2_u12_u6_n130 ) , .ZN( u2_u12_u6_n136 ) );
  NAND2_X1 u2_u12_u6_U35 (.A1( u2_u12_u6_n144 ) , .ZN( u2_u12_u6_n151 ) , .A2( u2_u12_u6_n158 ) );
  NAND2_X1 u2_u12_u6_U36 (.ZN( u2_u12_u6_n132 ) , .A1( u2_u12_u6_n91 ) , .A2( u2_u12_u6_n97 ) );
  AOI22_X1 u2_u12_u6_U37 (.B2( u2_u12_u6_n110 ) , .B1( u2_u12_u6_n111 ) , .A1( u2_u12_u6_n112 ) , .ZN( u2_u12_u6_n115 ) , .A2( u2_u12_u6_n161 ) );
  NAND4_X1 u2_u12_u6_U38 (.A3( u2_u12_u6_n109 ) , .ZN( u2_u12_u6_n112 ) , .A4( u2_u12_u6_n132 ) , .A2( u2_u12_u6_n147 ) , .A1( u2_u12_u6_n166 ) );
  NOR2_X1 u2_u12_u6_U39 (.ZN( u2_u12_u6_n109 ) , .A1( u2_u12_u6_n170 ) , .A2( u2_u12_u6_n173 ) );
  INV_X1 u2_u12_u6_U4 (.A( u2_u12_u6_n142 ) , .ZN( u2_u12_u6_n174 ) );
  NOR2_X1 u2_u12_u6_U40 (.A2( u2_u12_u6_n126 ) , .ZN( u2_u12_u6_n155 ) , .A1( u2_u12_u6_n160 ) );
  NAND2_X1 u2_u12_u6_U41 (.ZN( u2_u12_u6_n146 ) , .A2( u2_u12_u6_n94 ) , .A1( u2_u12_u6_n99 ) );
  AOI21_X1 u2_u12_u6_U42 (.A( u2_u12_u6_n144 ) , .B2( u2_u12_u6_n145 ) , .B1( u2_u12_u6_n146 ) , .ZN( u2_u12_u6_n150 ) );
  INV_X1 u2_u12_u6_U43 (.A( u2_u12_u6_n111 ) , .ZN( u2_u12_u6_n158 ) );
  NAND2_X1 u2_u12_u6_U44 (.ZN( u2_u12_u6_n127 ) , .A1( u2_u12_u6_n91 ) , .A2( u2_u12_u6_n92 ) );
  NAND2_X1 u2_u12_u6_U45 (.ZN( u2_u12_u6_n129 ) , .A2( u2_u12_u6_n95 ) , .A1( u2_u12_u6_n96 ) );
  INV_X1 u2_u12_u6_U46 (.A( u2_u12_u6_n144 ) , .ZN( u2_u12_u6_n159 ) );
  NAND2_X1 u2_u12_u6_U47 (.ZN( u2_u12_u6_n145 ) , .A2( u2_u12_u6_n97 ) , .A1( u2_u12_u6_n98 ) );
  NAND2_X1 u2_u12_u6_U48 (.ZN( u2_u12_u6_n148 ) , .A2( u2_u12_u6_n92 ) , .A1( u2_u12_u6_n94 ) );
  NAND2_X1 u2_u12_u6_U49 (.ZN( u2_u12_u6_n108 ) , .A2( u2_u12_u6_n139 ) , .A1( u2_u12_u6_n144 ) );
  NAND2_X1 u2_u12_u6_U5 (.A2( u2_u12_u6_n143 ) , .ZN( u2_u12_u6_n152 ) , .A1( u2_u12_u6_n166 ) );
  NAND2_X1 u2_u12_u6_U50 (.ZN( u2_u12_u6_n121 ) , .A2( u2_u12_u6_n95 ) , .A1( u2_u12_u6_n97 ) );
  NAND2_X1 u2_u12_u6_U51 (.ZN( u2_u12_u6_n107 ) , .A2( u2_u12_u6_n92 ) , .A1( u2_u12_u6_n95 ) );
  AND2_X1 u2_u12_u6_U52 (.ZN( u2_u12_u6_n118 ) , .A2( u2_u12_u6_n91 ) , .A1( u2_u12_u6_n99 ) );
  NAND2_X1 u2_u12_u6_U53 (.ZN( u2_u12_u6_n147 ) , .A2( u2_u12_u6_n98 ) , .A1( u2_u12_u6_n99 ) );
  NAND2_X1 u2_u12_u6_U54 (.ZN( u2_u12_u6_n128 ) , .A1( u2_u12_u6_n94 ) , .A2( u2_u12_u6_n96 ) );
  NAND2_X1 u2_u12_u6_U55 (.ZN( u2_u12_u6_n119 ) , .A2( u2_u12_u6_n95 ) , .A1( u2_u12_u6_n99 ) );
  NAND2_X1 u2_u12_u6_U56 (.ZN( u2_u12_u6_n123 ) , .A2( u2_u12_u6_n91 ) , .A1( u2_u12_u6_n96 ) );
  NAND2_X1 u2_u12_u6_U57 (.ZN( u2_u12_u6_n100 ) , .A2( u2_u12_u6_n92 ) , .A1( u2_u12_u6_n98 ) );
  NAND2_X1 u2_u12_u6_U58 (.ZN( u2_u12_u6_n122 ) , .A1( u2_u12_u6_n94 ) , .A2( u2_u12_u6_n97 ) );
  INV_X1 u2_u12_u6_U59 (.A( u2_u12_u6_n139 ) , .ZN( u2_u12_u6_n160 ) );
  AOI22_X1 u2_u12_u6_U6 (.B2( u2_u12_u6_n101 ) , .A1( u2_u12_u6_n102 ) , .ZN( u2_u12_u6_n103 ) , .B1( u2_u12_u6_n160 ) , .A2( u2_u12_u6_n161 ) );
  NAND2_X1 u2_u12_u6_U60 (.ZN( u2_u12_u6_n113 ) , .A1( u2_u12_u6_n96 ) , .A2( u2_u12_u6_n98 ) );
  NOR2_X1 u2_u12_u6_U61 (.A2( u2_u12_X_40 ) , .A1( u2_u12_X_41 ) , .ZN( u2_u12_u6_n126 ) );
  NOR2_X1 u2_u12_u6_U62 (.A2( u2_u12_X_39 ) , .A1( u2_u12_X_42 ) , .ZN( u2_u12_u6_n92 ) );
  NOR2_X1 u2_u12_u6_U63 (.A2( u2_u12_X_39 ) , .A1( u2_u12_u6_n156 ) , .ZN( u2_u12_u6_n97 ) );
  NOR2_X1 u2_u12_u6_U64 (.A2( u2_u12_X_38 ) , .A1( u2_u12_u6_n165 ) , .ZN( u2_u12_u6_n95 ) );
  NOR2_X1 u2_u12_u6_U65 (.A2( u2_u12_X_41 ) , .ZN( u2_u12_u6_n111 ) , .A1( u2_u12_u6_n157 ) );
  NOR2_X1 u2_u12_u6_U66 (.A2( u2_u12_X_37 ) , .A1( u2_u12_u6_n162 ) , .ZN( u2_u12_u6_n94 ) );
  NOR2_X1 u2_u12_u6_U67 (.A2( u2_u12_X_37 ) , .A1( u2_u12_X_38 ) , .ZN( u2_u12_u6_n91 ) );
  NAND2_X1 u2_u12_u6_U68 (.A1( u2_u12_X_41 ) , .ZN( u2_u12_u6_n144 ) , .A2( u2_u12_u6_n157 ) );
  NAND2_X1 u2_u12_u6_U69 (.A2( u2_u12_X_40 ) , .A1( u2_u12_X_41 ) , .ZN( u2_u12_u6_n139 ) );
  NOR2_X1 u2_u12_u6_U7 (.A1( u2_u12_u6_n118 ) , .ZN( u2_u12_u6_n143 ) , .A2( u2_u12_u6_n168 ) );
  AND2_X1 u2_u12_u6_U70 (.A1( u2_u12_X_39 ) , .A2( u2_u12_u6_n156 ) , .ZN( u2_u12_u6_n96 ) );
  AND2_X1 u2_u12_u6_U71 (.A1( u2_u12_X_39 ) , .A2( u2_u12_X_42 ) , .ZN( u2_u12_u6_n99 ) );
  INV_X1 u2_u12_u6_U72 (.A( u2_u12_X_40 ) , .ZN( u2_u12_u6_n157 ) );
  INV_X1 u2_u12_u6_U73 (.A( u2_u12_X_37 ) , .ZN( u2_u12_u6_n165 ) );
  INV_X1 u2_u12_u6_U74 (.A( u2_u12_X_38 ) , .ZN( u2_u12_u6_n162 ) );
  INV_X1 u2_u12_u6_U75 (.A( u2_u12_X_42 ) , .ZN( u2_u12_u6_n156 ) );
  NAND4_X1 u2_u12_u6_U76 (.ZN( u2_out12_32 ) , .A4( u2_u12_u6_n103 ) , .A3( u2_u12_u6_n104 ) , .A2( u2_u12_u6_n105 ) , .A1( u2_u12_u6_n106 ) );
  AOI22_X1 u2_u12_u6_U77 (.ZN( u2_u12_u6_n105 ) , .A2( u2_u12_u6_n108 ) , .A1( u2_u12_u6_n118 ) , .B2( u2_u12_u6_n126 ) , .B1( u2_u12_u6_n171 ) );
  AOI22_X1 u2_u12_u6_U78 (.ZN( u2_u12_u6_n104 ) , .A1( u2_u12_u6_n111 ) , .B1( u2_u12_u6_n124 ) , .B2( u2_u12_u6_n151 ) , .A2( u2_u12_u6_n93 ) );
  NAND4_X1 u2_u12_u6_U79 (.ZN( u2_out12_12 ) , .A4( u2_u12_u6_n114 ) , .A3( u2_u12_u6_n115 ) , .A2( u2_u12_u6_n116 ) , .A1( u2_u12_u6_n117 ) );
  INV_X1 u2_u12_u6_U8 (.ZN( u2_u12_u6_n172 ) , .A( u2_u12_u6_n88 ) );
  OAI22_X1 u2_u12_u6_U80 (.B2( u2_u12_u6_n111 ) , .ZN( u2_u12_u6_n116 ) , .B1( u2_u12_u6_n126 ) , .A2( u2_u12_u6_n164 ) , .A1( u2_u12_u6_n167 ) );
  OAI21_X1 u2_u12_u6_U81 (.A( u2_u12_u6_n108 ) , .ZN( u2_u12_u6_n117 ) , .B2( u2_u12_u6_n141 ) , .B1( u2_u12_u6_n163 ) );
  OAI211_X1 u2_u12_u6_U82 (.ZN( u2_out12_22 ) , .B( u2_u12_u6_n137 ) , .A( u2_u12_u6_n138 ) , .C2( u2_u12_u6_n139 ) , .C1( u2_u12_u6_n140 ) );
  AOI22_X1 u2_u12_u6_U83 (.B1( u2_u12_u6_n124 ) , .A2( u2_u12_u6_n125 ) , .A1( u2_u12_u6_n126 ) , .ZN( u2_u12_u6_n138 ) , .B2( u2_u12_u6_n161 ) );
  AND4_X1 u2_u12_u6_U84 (.A3( u2_u12_u6_n119 ) , .A1( u2_u12_u6_n120 ) , .A4( u2_u12_u6_n129 ) , .ZN( u2_u12_u6_n140 ) , .A2( u2_u12_u6_n143 ) );
  OAI211_X1 u2_u12_u6_U85 (.ZN( u2_out12_7 ) , .B( u2_u12_u6_n153 ) , .C2( u2_u12_u6_n154 ) , .C1( u2_u12_u6_n155 ) , .A( u2_u12_u6_n174 ) );
  NOR3_X1 u2_u12_u6_U86 (.A1( u2_u12_u6_n141 ) , .ZN( u2_u12_u6_n154 ) , .A3( u2_u12_u6_n164 ) , .A2( u2_u12_u6_n171 ) );
  AOI211_X1 u2_u12_u6_U87 (.B( u2_u12_u6_n149 ) , .A( u2_u12_u6_n150 ) , .C2( u2_u12_u6_n151 ) , .C1( u2_u12_u6_n152 ) , .ZN( u2_u12_u6_n153 ) );
  NAND3_X1 u2_u12_u6_U88 (.A2( u2_u12_u6_n123 ) , .ZN( u2_u12_u6_n125 ) , .A1( u2_u12_u6_n130 ) , .A3( u2_u12_u6_n131 ) );
  NAND3_X1 u2_u12_u6_U89 (.A3( u2_u12_u6_n133 ) , .ZN( u2_u12_u6_n141 ) , .A1( u2_u12_u6_n145 ) , .A2( u2_u12_u6_n148 ) );
  OAI21_X1 u2_u12_u6_U9 (.A( u2_u12_u6_n159 ) , .B1( u2_u12_u6_n169 ) , .B2( u2_u12_u6_n173 ) , .ZN( u2_u12_u6_n90 ) );
  NAND3_X1 u2_u12_u6_U90 (.ZN( u2_u12_u6_n101 ) , .A3( u2_u12_u6_n107 ) , .A2( u2_u12_u6_n121 ) , .A1( u2_u12_u6_n127 ) );
  NAND3_X1 u2_u12_u6_U91 (.ZN( u2_u12_u6_n102 ) , .A3( u2_u12_u6_n130 ) , .A2( u2_u12_u6_n145 ) , .A1( u2_u12_u6_n166 ) );
  NAND3_X1 u2_u12_u6_U92 (.A3( u2_u12_u6_n113 ) , .A1( u2_u12_u6_n119 ) , .A2( u2_u12_u6_n123 ) , .ZN( u2_u12_u6_n93 ) );
  NAND3_X1 u2_u12_u6_U93 (.ZN( u2_u12_u6_n142 ) , .A2( u2_u12_u6_n172 ) , .A3( u2_u12_u6_n89 ) , .A1( u2_u12_u6_n90 ) );
  AND3_X1 u2_u12_u7_U10 (.A3( u2_u12_u7_n110 ) , .A2( u2_u12_u7_n127 ) , .A1( u2_u12_u7_n132 ) , .ZN( u2_u12_u7_n92 ) );
  OAI21_X1 u2_u12_u7_U11 (.A( u2_u12_u7_n161 ) , .B1( u2_u12_u7_n168 ) , .B2( u2_u12_u7_n173 ) , .ZN( u2_u12_u7_n91 ) );
  AOI211_X1 u2_u12_u7_U12 (.A( u2_u12_u7_n117 ) , .ZN( u2_u12_u7_n118 ) , .C2( u2_u12_u7_n126 ) , .C1( u2_u12_u7_n177 ) , .B( u2_u12_u7_n180 ) );
  OAI22_X1 u2_u12_u7_U13 (.B1( u2_u12_u7_n115 ) , .ZN( u2_u12_u7_n117 ) , .A2( u2_u12_u7_n133 ) , .A1( u2_u12_u7_n137 ) , .B2( u2_u12_u7_n162 ) );
  INV_X1 u2_u12_u7_U14 (.A( u2_u12_u7_n116 ) , .ZN( u2_u12_u7_n180 ) );
  NOR3_X1 u2_u12_u7_U15 (.ZN( u2_u12_u7_n115 ) , .A3( u2_u12_u7_n145 ) , .A2( u2_u12_u7_n168 ) , .A1( u2_u12_u7_n169 ) );
  OAI211_X1 u2_u12_u7_U16 (.B( u2_u12_u7_n122 ) , .A( u2_u12_u7_n123 ) , .C2( u2_u12_u7_n124 ) , .ZN( u2_u12_u7_n154 ) , .C1( u2_u12_u7_n162 ) );
  AOI222_X1 u2_u12_u7_U17 (.ZN( u2_u12_u7_n122 ) , .C2( u2_u12_u7_n126 ) , .C1( u2_u12_u7_n145 ) , .B1( u2_u12_u7_n161 ) , .A2( u2_u12_u7_n165 ) , .B2( u2_u12_u7_n170 ) , .A1( u2_u12_u7_n176 ) );
  INV_X1 u2_u12_u7_U18 (.A( u2_u12_u7_n133 ) , .ZN( u2_u12_u7_n176 ) );
  NOR3_X1 u2_u12_u7_U19 (.A2( u2_u12_u7_n134 ) , .A1( u2_u12_u7_n135 ) , .ZN( u2_u12_u7_n136 ) , .A3( u2_u12_u7_n171 ) );
  NOR2_X1 u2_u12_u7_U20 (.A1( u2_u12_u7_n130 ) , .A2( u2_u12_u7_n134 ) , .ZN( u2_u12_u7_n153 ) );
  INV_X1 u2_u12_u7_U21 (.A( u2_u12_u7_n101 ) , .ZN( u2_u12_u7_n165 ) );
  NOR2_X1 u2_u12_u7_U22 (.ZN( u2_u12_u7_n111 ) , .A2( u2_u12_u7_n134 ) , .A1( u2_u12_u7_n169 ) );
  AOI21_X1 u2_u12_u7_U23 (.ZN( u2_u12_u7_n104 ) , .B2( u2_u12_u7_n112 ) , .B1( u2_u12_u7_n127 ) , .A( u2_u12_u7_n164 ) );
  AOI21_X1 u2_u12_u7_U24 (.ZN( u2_u12_u7_n106 ) , .B1( u2_u12_u7_n133 ) , .B2( u2_u12_u7_n146 ) , .A( u2_u12_u7_n162 ) );
  AOI21_X1 u2_u12_u7_U25 (.A( u2_u12_u7_n101 ) , .ZN( u2_u12_u7_n107 ) , .B2( u2_u12_u7_n128 ) , .B1( u2_u12_u7_n175 ) );
  INV_X1 u2_u12_u7_U26 (.A( u2_u12_u7_n138 ) , .ZN( u2_u12_u7_n171 ) );
  INV_X1 u2_u12_u7_U27 (.A( u2_u12_u7_n131 ) , .ZN( u2_u12_u7_n177 ) );
  INV_X1 u2_u12_u7_U28 (.A( u2_u12_u7_n110 ) , .ZN( u2_u12_u7_n174 ) );
  NAND2_X1 u2_u12_u7_U29 (.A1( u2_u12_u7_n129 ) , .A2( u2_u12_u7_n132 ) , .ZN( u2_u12_u7_n149 ) );
  OAI21_X1 u2_u12_u7_U3 (.ZN( u2_u12_u7_n159 ) , .A( u2_u12_u7_n165 ) , .B2( u2_u12_u7_n171 ) , .B1( u2_u12_u7_n174 ) );
  NAND2_X1 u2_u12_u7_U30 (.A1( u2_u12_u7_n113 ) , .A2( u2_u12_u7_n124 ) , .ZN( u2_u12_u7_n130 ) );
  INV_X1 u2_u12_u7_U31 (.A( u2_u12_u7_n112 ) , .ZN( u2_u12_u7_n173 ) );
  INV_X1 u2_u12_u7_U32 (.A( u2_u12_u7_n128 ) , .ZN( u2_u12_u7_n168 ) );
  INV_X1 u2_u12_u7_U33 (.A( u2_u12_u7_n148 ) , .ZN( u2_u12_u7_n169 ) );
  INV_X1 u2_u12_u7_U34 (.A( u2_u12_u7_n127 ) , .ZN( u2_u12_u7_n179 ) );
  NOR2_X1 u2_u12_u7_U35 (.ZN( u2_u12_u7_n101 ) , .A2( u2_u12_u7_n150 ) , .A1( u2_u12_u7_n156 ) );
  AOI211_X1 u2_u12_u7_U36 (.B( u2_u12_u7_n154 ) , .A( u2_u12_u7_n155 ) , .C1( u2_u12_u7_n156 ) , .ZN( u2_u12_u7_n157 ) , .C2( u2_u12_u7_n172 ) );
  INV_X1 u2_u12_u7_U37 (.A( u2_u12_u7_n153 ) , .ZN( u2_u12_u7_n172 ) );
  AOI211_X1 u2_u12_u7_U38 (.B( u2_u12_u7_n139 ) , .A( u2_u12_u7_n140 ) , .C2( u2_u12_u7_n141 ) , .ZN( u2_u12_u7_n142 ) , .C1( u2_u12_u7_n156 ) );
  NAND4_X1 u2_u12_u7_U39 (.A3( u2_u12_u7_n127 ) , .A2( u2_u12_u7_n128 ) , .A1( u2_u12_u7_n129 ) , .ZN( u2_u12_u7_n141 ) , .A4( u2_u12_u7_n147 ) );
  INV_X1 u2_u12_u7_U4 (.A( u2_u12_u7_n111 ) , .ZN( u2_u12_u7_n170 ) );
  AOI21_X1 u2_u12_u7_U40 (.A( u2_u12_u7_n137 ) , .B1( u2_u12_u7_n138 ) , .ZN( u2_u12_u7_n139 ) , .B2( u2_u12_u7_n146 ) );
  OAI22_X1 u2_u12_u7_U41 (.B1( u2_u12_u7_n136 ) , .ZN( u2_u12_u7_n140 ) , .A1( u2_u12_u7_n153 ) , .B2( u2_u12_u7_n162 ) , .A2( u2_u12_u7_n164 ) );
  AOI21_X1 u2_u12_u7_U42 (.ZN( u2_u12_u7_n123 ) , .B1( u2_u12_u7_n165 ) , .B2( u2_u12_u7_n177 ) , .A( u2_u12_u7_n97 ) );
  AOI21_X1 u2_u12_u7_U43 (.B2( u2_u12_u7_n113 ) , .B1( u2_u12_u7_n124 ) , .A( u2_u12_u7_n125 ) , .ZN( u2_u12_u7_n97 ) );
  INV_X1 u2_u12_u7_U44 (.A( u2_u12_u7_n125 ) , .ZN( u2_u12_u7_n161 ) );
  INV_X1 u2_u12_u7_U45 (.A( u2_u12_u7_n152 ) , .ZN( u2_u12_u7_n162 ) );
  AOI22_X1 u2_u12_u7_U46 (.A2( u2_u12_u7_n114 ) , .ZN( u2_u12_u7_n119 ) , .B1( u2_u12_u7_n130 ) , .A1( u2_u12_u7_n156 ) , .B2( u2_u12_u7_n165 ) );
  NAND2_X1 u2_u12_u7_U47 (.A2( u2_u12_u7_n112 ) , .ZN( u2_u12_u7_n114 ) , .A1( u2_u12_u7_n175 ) );
  AND2_X1 u2_u12_u7_U48 (.ZN( u2_u12_u7_n145 ) , .A2( u2_u12_u7_n98 ) , .A1( u2_u12_u7_n99 ) );
  NOR2_X1 u2_u12_u7_U49 (.ZN( u2_u12_u7_n137 ) , .A1( u2_u12_u7_n150 ) , .A2( u2_u12_u7_n161 ) );
  INV_X1 u2_u12_u7_U5 (.A( u2_u12_u7_n149 ) , .ZN( u2_u12_u7_n175 ) );
  AOI21_X1 u2_u12_u7_U50 (.ZN( u2_u12_u7_n105 ) , .B2( u2_u12_u7_n110 ) , .A( u2_u12_u7_n125 ) , .B1( u2_u12_u7_n147 ) );
  NAND2_X1 u2_u12_u7_U51 (.ZN( u2_u12_u7_n146 ) , .A1( u2_u12_u7_n95 ) , .A2( u2_u12_u7_n98 ) );
  NAND2_X1 u2_u12_u7_U52 (.A2( u2_u12_u7_n103 ) , .ZN( u2_u12_u7_n147 ) , .A1( u2_u12_u7_n93 ) );
  NAND2_X1 u2_u12_u7_U53 (.A1( u2_u12_u7_n103 ) , .ZN( u2_u12_u7_n127 ) , .A2( u2_u12_u7_n99 ) );
  OR2_X1 u2_u12_u7_U54 (.ZN( u2_u12_u7_n126 ) , .A2( u2_u12_u7_n152 ) , .A1( u2_u12_u7_n156 ) );
  NAND2_X1 u2_u12_u7_U55 (.A2( u2_u12_u7_n102 ) , .A1( u2_u12_u7_n103 ) , .ZN( u2_u12_u7_n133 ) );
  NAND2_X1 u2_u12_u7_U56 (.ZN( u2_u12_u7_n112 ) , .A2( u2_u12_u7_n96 ) , .A1( u2_u12_u7_n99 ) );
  NAND2_X1 u2_u12_u7_U57 (.A2( u2_u12_u7_n102 ) , .ZN( u2_u12_u7_n128 ) , .A1( u2_u12_u7_n98 ) );
  NAND2_X1 u2_u12_u7_U58 (.A1( u2_u12_u7_n100 ) , .ZN( u2_u12_u7_n113 ) , .A2( u2_u12_u7_n93 ) );
  NAND2_X1 u2_u12_u7_U59 (.A2( u2_u12_u7_n102 ) , .ZN( u2_u12_u7_n124 ) , .A1( u2_u12_u7_n96 ) );
  INV_X1 u2_u12_u7_U6 (.A( u2_u12_u7_n154 ) , .ZN( u2_u12_u7_n178 ) );
  NAND2_X1 u2_u12_u7_U60 (.ZN( u2_u12_u7_n110 ) , .A1( u2_u12_u7_n95 ) , .A2( u2_u12_u7_n96 ) );
  INV_X1 u2_u12_u7_U61 (.A( u2_u12_u7_n150 ) , .ZN( u2_u12_u7_n164 ) );
  AND2_X1 u2_u12_u7_U62 (.ZN( u2_u12_u7_n134 ) , .A1( u2_u12_u7_n93 ) , .A2( u2_u12_u7_n98 ) );
  NAND2_X1 u2_u12_u7_U63 (.A1( u2_u12_u7_n100 ) , .A2( u2_u12_u7_n102 ) , .ZN( u2_u12_u7_n129 ) );
  NAND2_X1 u2_u12_u7_U64 (.A2( u2_u12_u7_n103 ) , .ZN( u2_u12_u7_n131 ) , .A1( u2_u12_u7_n95 ) );
  NAND2_X1 u2_u12_u7_U65 (.A1( u2_u12_u7_n100 ) , .ZN( u2_u12_u7_n138 ) , .A2( u2_u12_u7_n99 ) );
  NAND2_X1 u2_u12_u7_U66 (.ZN( u2_u12_u7_n132 ) , .A1( u2_u12_u7_n93 ) , .A2( u2_u12_u7_n96 ) );
  NAND2_X1 u2_u12_u7_U67 (.A1( u2_u12_u7_n100 ) , .ZN( u2_u12_u7_n148 ) , .A2( u2_u12_u7_n95 ) );
  NOR2_X1 u2_u12_u7_U68 (.A2( u2_u12_X_47 ) , .ZN( u2_u12_u7_n150 ) , .A1( u2_u12_u7_n163 ) );
  NOR2_X1 u2_u12_u7_U69 (.A2( u2_u12_X_43 ) , .A1( u2_u12_X_44 ) , .ZN( u2_u12_u7_n103 ) );
  AOI211_X1 u2_u12_u7_U7 (.ZN( u2_u12_u7_n116 ) , .A( u2_u12_u7_n155 ) , .C1( u2_u12_u7_n161 ) , .C2( u2_u12_u7_n171 ) , .B( u2_u12_u7_n94 ) );
  NOR2_X1 u2_u12_u7_U70 (.A2( u2_u12_X_48 ) , .A1( u2_u12_u7_n166 ) , .ZN( u2_u12_u7_n95 ) );
  NOR2_X1 u2_u12_u7_U71 (.A2( u2_u12_X_45 ) , .A1( u2_u12_X_48 ) , .ZN( u2_u12_u7_n99 ) );
  NOR2_X1 u2_u12_u7_U72 (.A2( u2_u12_X_44 ) , .A1( u2_u12_u7_n167 ) , .ZN( u2_u12_u7_n98 ) );
  NOR2_X1 u2_u12_u7_U73 (.A2( u2_u12_X_46 ) , .A1( u2_u12_X_47 ) , .ZN( u2_u12_u7_n152 ) );
  AND2_X1 u2_u12_u7_U74 (.A1( u2_u12_X_47 ) , .ZN( u2_u12_u7_n156 ) , .A2( u2_u12_u7_n163 ) );
  NAND2_X1 u2_u12_u7_U75 (.A2( u2_u12_X_46 ) , .A1( u2_u12_X_47 ) , .ZN( u2_u12_u7_n125 ) );
  AND2_X1 u2_u12_u7_U76 (.A2( u2_u12_X_45 ) , .A1( u2_u12_X_48 ) , .ZN( u2_u12_u7_n102 ) );
  AND2_X1 u2_u12_u7_U77 (.A2( u2_u12_X_43 ) , .A1( u2_u12_X_44 ) , .ZN( u2_u12_u7_n96 ) );
  AND2_X1 u2_u12_u7_U78 (.A1( u2_u12_X_44 ) , .ZN( u2_u12_u7_n100 ) , .A2( u2_u12_u7_n167 ) );
  AND2_X1 u2_u12_u7_U79 (.A1( u2_u12_X_48 ) , .A2( u2_u12_u7_n166 ) , .ZN( u2_u12_u7_n93 ) );
  OAI222_X1 u2_u12_u7_U8 (.C2( u2_u12_u7_n101 ) , .B2( u2_u12_u7_n111 ) , .A1( u2_u12_u7_n113 ) , .C1( u2_u12_u7_n146 ) , .A2( u2_u12_u7_n162 ) , .B1( u2_u12_u7_n164 ) , .ZN( u2_u12_u7_n94 ) );
  INV_X1 u2_u12_u7_U80 (.A( u2_u12_X_46 ) , .ZN( u2_u12_u7_n163 ) );
  INV_X1 u2_u12_u7_U81 (.A( u2_u12_X_43 ) , .ZN( u2_u12_u7_n167 ) );
  INV_X1 u2_u12_u7_U82 (.A( u2_u12_X_45 ) , .ZN( u2_u12_u7_n166 ) );
  NAND4_X1 u2_u12_u7_U83 (.ZN( u2_out12_27 ) , .A4( u2_u12_u7_n118 ) , .A3( u2_u12_u7_n119 ) , .A2( u2_u12_u7_n120 ) , .A1( u2_u12_u7_n121 ) );
  OAI21_X1 u2_u12_u7_U84 (.ZN( u2_u12_u7_n121 ) , .B2( u2_u12_u7_n145 ) , .A( u2_u12_u7_n150 ) , .B1( u2_u12_u7_n174 ) );
  OAI21_X1 u2_u12_u7_U85 (.ZN( u2_u12_u7_n120 ) , .A( u2_u12_u7_n161 ) , .B2( u2_u12_u7_n170 ) , .B1( u2_u12_u7_n179 ) );
  NAND4_X1 u2_u12_u7_U86 (.ZN( u2_out12_21 ) , .A4( u2_u12_u7_n157 ) , .A3( u2_u12_u7_n158 ) , .A2( u2_u12_u7_n159 ) , .A1( u2_u12_u7_n160 ) );
  OAI21_X1 u2_u12_u7_U87 (.B1( u2_u12_u7_n145 ) , .ZN( u2_u12_u7_n160 ) , .A( u2_u12_u7_n161 ) , .B2( u2_u12_u7_n177 ) );
  AOI22_X1 u2_u12_u7_U88 (.B2( u2_u12_u7_n149 ) , .B1( u2_u12_u7_n150 ) , .A2( u2_u12_u7_n151 ) , .A1( u2_u12_u7_n152 ) , .ZN( u2_u12_u7_n158 ) );
  NAND4_X1 u2_u12_u7_U89 (.ZN( u2_out12_15 ) , .A4( u2_u12_u7_n142 ) , .A3( u2_u12_u7_n143 ) , .A2( u2_u12_u7_n144 ) , .A1( u2_u12_u7_n178 ) );
  OAI221_X1 u2_u12_u7_U9 (.C1( u2_u12_u7_n101 ) , .C2( u2_u12_u7_n147 ) , .ZN( u2_u12_u7_n155 ) , .B2( u2_u12_u7_n162 ) , .A( u2_u12_u7_n91 ) , .B1( u2_u12_u7_n92 ) );
  OR2_X1 u2_u12_u7_U90 (.A2( u2_u12_u7_n125 ) , .A1( u2_u12_u7_n129 ) , .ZN( u2_u12_u7_n144 ) );
  AOI22_X1 u2_u12_u7_U91 (.A2( u2_u12_u7_n126 ) , .ZN( u2_u12_u7_n143 ) , .B2( u2_u12_u7_n165 ) , .B1( u2_u12_u7_n173 ) , .A1( u2_u12_u7_n174 ) );
  NAND4_X1 u2_u12_u7_U92 (.ZN( u2_out12_5 ) , .A4( u2_u12_u7_n108 ) , .A3( u2_u12_u7_n109 ) , .A1( u2_u12_u7_n116 ) , .A2( u2_u12_u7_n123 ) );
  AOI22_X1 u2_u12_u7_U93 (.ZN( u2_u12_u7_n109 ) , .A2( u2_u12_u7_n126 ) , .B2( u2_u12_u7_n145 ) , .B1( u2_u12_u7_n156 ) , .A1( u2_u12_u7_n171 ) );
  NOR4_X1 u2_u12_u7_U94 (.A4( u2_u12_u7_n104 ) , .A3( u2_u12_u7_n105 ) , .A2( u2_u12_u7_n106 ) , .A1( u2_u12_u7_n107 ) , .ZN( u2_u12_u7_n108 ) );
  NAND3_X1 u2_u12_u7_U95 (.A3( u2_u12_u7_n146 ) , .A2( u2_u12_u7_n147 ) , .A1( u2_u12_u7_n148 ) , .ZN( u2_u12_u7_n151 ) );
  NAND3_X1 u2_u12_u7_U96 (.A3( u2_u12_u7_n131 ) , .A2( u2_u12_u7_n132 ) , .A1( u2_u12_u7_n133 ) , .ZN( u2_u12_u7_n135 ) );
  XOR2_X1 u2_u3_U1 (.B( u2_K4_9 ) , .A( u2_R2_6 ) , .Z( u2_u3_X_9 ) );
  XOR2_X1 u2_u3_U10 (.B( u2_K4_45 ) , .A( u2_R2_30 ) , .Z( u2_u3_X_45 ) );
  XOR2_X1 u2_u3_U11 (.B( u2_K4_44 ) , .A( u2_R2_29 ) , .Z( u2_u3_X_44 ) );
  XOR2_X1 u2_u3_U12 (.B( u2_K4_43 ) , .A( u2_R2_28 ) , .Z( u2_u3_X_43 ) );
  XOR2_X1 u2_u3_U16 (.B( u2_K4_3 ) , .A( u2_R2_2 ) , .Z( u2_u3_X_3 ) );
  XOR2_X1 u2_u3_U2 (.B( u2_K4_8 ) , .A( u2_R2_5 ) , .Z( u2_u3_X_8 ) );
  XOR2_X1 u2_u3_U27 (.B( u2_K4_2 ) , .A( u2_R2_1 ) , .Z( u2_u3_X_2 ) );
  XOR2_X1 u2_u3_U3 (.B( u2_K4_7 ) , .A( u2_R2_4 ) , .Z( u2_u3_X_7 ) );
  XOR2_X1 u2_u3_U38 (.B( u2_K4_1 ) , .A( u2_R2_32 ) , .Z( u2_u3_X_1 ) );
  XOR2_X1 u2_u3_U4 (.B( u2_K4_6 ) , .A( u2_R2_5 ) , .Z( u2_u3_X_6 ) );
  XOR2_X1 u2_u3_U46 (.B( u2_K4_12 ) , .A( u2_R2_9 ) , .Z( u2_u3_X_12 ) );
  XOR2_X1 u2_u3_U47 (.B( u2_K4_11 ) , .A( u2_R2_8 ) , .Z( u2_u3_X_11 ) );
  XOR2_X1 u2_u3_U48 (.B( u2_K4_10 ) , .A( u2_R2_7 ) , .Z( u2_u3_X_10 ) );
  XOR2_X1 u2_u3_U5 (.B( u2_K4_5 ) , .A( u2_R2_4 ) , .Z( u2_u3_X_5 ) );
  XOR2_X1 u2_u3_U6 (.B( u2_K4_4 ) , .A( u2_R2_3 ) , .Z( u2_u3_X_4 ) );
  XOR2_X1 u2_u3_U7 (.B( u2_K4_48 ) , .A( u2_R2_1 ) , .Z( u2_u3_X_48 ) );
  XOR2_X1 u2_u3_U8 (.B( u2_K4_47 ) , .A( u2_R2_32 ) , .Z( u2_u3_X_47 ) );
  XOR2_X1 u2_u3_U9 (.B( u2_K4_46 ) , .A( u2_R2_31 ) , .Z( u2_u3_X_46 ) );
  AND3_X1 u2_u3_u0_U10 (.A2( u2_u3_u0_n112 ) , .ZN( u2_u3_u0_n127 ) , .A3( u2_u3_u0_n130 ) , .A1( u2_u3_u0_n148 ) );
  NAND2_X1 u2_u3_u0_U11 (.ZN( u2_u3_u0_n113 ) , .A1( u2_u3_u0_n139 ) , .A2( u2_u3_u0_n149 ) );
  AND2_X1 u2_u3_u0_U12 (.ZN( u2_u3_u0_n107 ) , .A1( u2_u3_u0_n130 ) , .A2( u2_u3_u0_n140 ) );
  AND2_X1 u2_u3_u0_U13 (.A2( u2_u3_u0_n129 ) , .A1( u2_u3_u0_n130 ) , .ZN( u2_u3_u0_n151 ) );
  AND2_X1 u2_u3_u0_U14 (.A1( u2_u3_u0_n108 ) , .A2( u2_u3_u0_n125 ) , .ZN( u2_u3_u0_n145 ) );
  INV_X1 u2_u3_u0_U15 (.A( u2_u3_u0_n143 ) , .ZN( u2_u3_u0_n173 ) );
  NOR2_X1 u2_u3_u0_U16 (.A2( u2_u3_u0_n136 ) , .ZN( u2_u3_u0_n147 ) , .A1( u2_u3_u0_n160 ) );
  INV_X1 u2_u3_u0_U17 (.ZN( u2_u3_u0_n172 ) , .A( u2_u3_u0_n88 ) );
  OAI222_X1 u2_u3_u0_U18 (.C1( u2_u3_u0_n108 ) , .A1( u2_u3_u0_n125 ) , .B2( u2_u3_u0_n128 ) , .B1( u2_u3_u0_n144 ) , .A2( u2_u3_u0_n158 ) , .C2( u2_u3_u0_n161 ) , .ZN( u2_u3_u0_n88 ) );
  AOI21_X1 u2_u3_u0_U19 (.B1( u2_u3_u0_n103 ) , .ZN( u2_u3_u0_n132 ) , .A( u2_u3_u0_n165 ) , .B2( u2_u3_u0_n93 ) );
  INV_X1 u2_u3_u0_U20 (.A( u2_u3_u0_n142 ) , .ZN( u2_u3_u0_n165 ) );
  OAI22_X1 u2_u3_u0_U21 (.B1( u2_u3_u0_n125 ) , .ZN( u2_u3_u0_n126 ) , .A1( u2_u3_u0_n138 ) , .A2( u2_u3_u0_n146 ) , .B2( u2_u3_u0_n147 ) );
  OAI22_X1 u2_u3_u0_U22 (.B1( u2_u3_u0_n131 ) , .A1( u2_u3_u0_n144 ) , .B2( u2_u3_u0_n147 ) , .A2( u2_u3_u0_n90 ) , .ZN( u2_u3_u0_n91 ) );
  AND3_X1 u2_u3_u0_U23 (.A3( u2_u3_u0_n121 ) , .A2( u2_u3_u0_n125 ) , .A1( u2_u3_u0_n148 ) , .ZN( u2_u3_u0_n90 ) );
  INV_X1 u2_u3_u0_U24 (.A( u2_u3_u0_n136 ) , .ZN( u2_u3_u0_n161 ) );
  AOI22_X1 u2_u3_u0_U25 (.B2( u2_u3_u0_n109 ) , .A2( u2_u3_u0_n110 ) , .ZN( u2_u3_u0_n111 ) , .B1( u2_u3_u0_n118 ) , .A1( u2_u3_u0_n160 ) );
  NAND2_X1 u2_u3_u0_U26 (.A2( u2_u3_u0_n103 ) , .ZN( u2_u3_u0_n140 ) , .A1( u2_u3_u0_n94 ) );
  INV_X1 u2_u3_u0_U27 (.A( u2_u3_u0_n118 ) , .ZN( u2_u3_u0_n158 ) );
  AOI21_X1 u2_u3_u0_U28 (.ZN( u2_u3_u0_n104 ) , .B1( u2_u3_u0_n107 ) , .B2( u2_u3_u0_n141 ) , .A( u2_u3_u0_n144 ) );
  AOI21_X1 u2_u3_u0_U29 (.B1( u2_u3_u0_n127 ) , .B2( u2_u3_u0_n129 ) , .A( u2_u3_u0_n138 ) , .ZN( u2_u3_u0_n96 ) );
  INV_X1 u2_u3_u0_U3 (.A( u2_u3_u0_n113 ) , .ZN( u2_u3_u0_n166 ) );
  NOR2_X1 u2_u3_u0_U30 (.A1( u2_u3_u0_n120 ) , .ZN( u2_u3_u0_n143 ) , .A2( u2_u3_u0_n167 ) );
  OAI221_X1 u2_u3_u0_U31 (.C1( u2_u3_u0_n112 ) , .ZN( u2_u3_u0_n120 ) , .B1( u2_u3_u0_n138 ) , .B2( u2_u3_u0_n141 ) , .C2( u2_u3_u0_n147 ) , .A( u2_u3_u0_n172 ) );
  AOI21_X1 u2_u3_u0_U32 (.ZN( u2_u3_u0_n116 ) , .B2( u2_u3_u0_n142 ) , .A( u2_u3_u0_n144 ) , .B1( u2_u3_u0_n166 ) );
  NAND2_X1 u2_u3_u0_U33 (.A1( u2_u3_u0_n101 ) , .A2( u2_u3_u0_n102 ) , .ZN( u2_u3_u0_n150 ) );
  INV_X1 u2_u3_u0_U34 (.A( u2_u3_u0_n138 ) , .ZN( u2_u3_u0_n160 ) );
  NAND2_X1 u2_u3_u0_U35 (.ZN( u2_u3_u0_n108 ) , .A1( u2_u3_u0_n92 ) , .A2( u2_u3_u0_n94 ) );
  NAND2_X1 u2_u3_u0_U36 (.A2( u2_u3_u0_n102 ) , .A1( u2_u3_u0_n103 ) , .ZN( u2_u3_u0_n149 ) );
  NAND2_X1 u2_u3_u0_U37 (.A1( u2_u3_u0_n101 ) , .ZN( u2_u3_u0_n130 ) , .A2( u2_u3_u0_n94 ) );
  NAND2_X1 u2_u3_u0_U38 (.A2( u2_u3_u0_n102 ) , .ZN( u2_u3_u0_n114 ) , .A1( u2_u3_u0_n92 ) );
  NAND2_X1 u2_u3_u0_U39 (.A2( u2_u3_u0_n101 ) , .ZN( u2_u3_u0_n121 ) , .A1( u2_u3_u0_n93 ) );
  AOI21_X1 u2_u3_u0_U4 (.B2( u2_u3_u0_n131 ) , .ZN( u2_u3_u0_n134 ) , .B1( u2_u3_u0_n151 ) , .A( u2_u3_u0_n158 ) );
  NAND2_X1 u2_u3_u0_U40 (.ZN( u2_u3_u0_n112 ) , .A2( u2_u3_u0_n92 ) , .A1( u2_u3_u0_n93 ) );
  OR3_X1 u2_u3_u0_U41 (.A3( u2_u3_u0_n152 ) , .A2( u2_u3_u0_n153 ) , .A1( u2_u3_u0_n154 ) , .ZN( u2_u3_u0_n155 ) );
  AOI21_X1 u2_u3_u0_U42 (.A( u2_u3_u0_n144 ) , .B2( u2_u3_u0_n145 ) , .B1( u2_u3_u0_n146 ) , .ZN( u2_u3_u0_n154 ) );
  AOI21_X1 u2_u3_u0_U43 (.B2( u2_u3_u0_n150 ) , .B1( u2_u3_u0_n151 ) , .ZN( u2_u3_u0_n152 ) , .A( u2_u3_u0_n158 ) );
  AOI21_X1 u2_u3_u0_U44 (.A( u2_u3_u0_n147 ) , .B2( u2_u3_u0_n148 ) , .B1( u2_u3_u0_n149 ) , .ZN( u2_u3_u0_n153 ) );
  INV_X1 u2_u3_u0_U45 (.ZN( u2_u3_u0_n171 ) , .A( u2_u3_u0_n99 ) );
  OAI211_X1 u2_u3_u0_U46 (.C2( u2_u3_u0_n140 ) , .C1( u2_u3_u0_n161 ) , .A( u2_u3_u0_n169 ) , .B( u2_u3_u0_n98 ) , .ZN( u2_u3_u0_n99 ) );
  AOI211_X1 u2_u3_u0_U47 (.C1( u2_u3_u0_n118 ) , .A( u2_u3_u0_n123 ) , .B( u2_u3_u0_n96 ) , .C2( u2_u3_u0_n97 ) , .ZN( u2_u3_u0_n98 ) );
  INV_X1 u2_u3_u0_U48 (.ZN( u2_u3_u0_n169 ) , .A( u2_u3_u0_n91 ) );
  NOR2_X1 u2_u3_u0_U49 (.A2( u2_u3_X_2 ) , .ZN( u2_u3_u0_n103 ) , .A1( u2_u3_u0_n164 ) );
  NOR2_X1 u2_u3_u0_U5 (.A1( u2_u3_u0_n108 ) , .ZN( u2_u3_u0_n123 ) , .A2( u2_u3_u0_n158 ) );
  NOR2_X1 u2_u3_u0_U50 (.A2( u2_u3_X_1 ) , .A1( u2_u3_X_2 ) , .ZN( u2_u3_u0_n92 ) );
  NOR2_X1 u2_u3_u0_U51 (.A2( u2_u3_X_4 ) , .A1( u2_u3_X_5 ) , .ZN( u2_u3_u0_n118 ) );
  NOR2_X1 u2_u3_u0_U52 (.A2( u2_u3_X_1 ) , .ZN( u2_u3_u0_n101 ) , .A1( u2_u3_u0_n163 ) );
  NAND2_X1 u2_u3_u0_U53 (.A2( u2_u3_X_4 ) , .A1( u2_u3_X_5 ) , .ZN( u2_u3_u0_n144 ) );
  NOR2_X1 u2_u3_u0_U54 (.A2( u2_u3_X_5 ) , .ZN( u2_u3_u0_n136 ) , .A1( u2_u3_u0_n159 ) );
  NAND2_X1 u2_u3_u0_U55 (.A1( u2_u3_X_5 ) , .ZN( u2_u3_u0_n138 ) , .A2( u2_u3_u0_n159 ) );
  NOR2_X1 u2_u3_u0_U56 (.A2( u2_u3_X_6 ) , .ZN( u2_u3_u0_n100 ) , .A1( u2_u3_u0_n162 ) );
  AND2_X1 u2_u3_u0_U57 (.A2( u2_u3_X_3 ) , .A1( u2_u3_X_6 ) , .ZN( u2_u3_u0_n102 ) );
  AND2_X1 u2_u3_u0_U58 (.A1( u2_u3_X_6 ) , .A2( u2_u3_u0_n162 ) , .ZN( u2_u3_u0_n93 ) );
  INV_X1 u2_u3_u0_U59 (.A( u2_u3_X_4 ) , .ZN( u2_u3_u0_n159 ) );
  OAI21_X1 u2_u3_u0_U6 (.B1( u2_u3_u0_n150 ) , .B2( u2_u3_u0_n158 ) , .A( u2_u3_u0_n172 ) , .ZN( u2_u3_u0_n89 ) );
  INV_X1 u2_u3_u0_U60 (.A( u2_u3_X_1 ) , .ZN( u2_u3_u0_n164 ) );
  INV_X1 u2_u3_u0_U61 (.A( u2_u3_X_2 ) , .ZN( u2_u3_u0_n163 ) );
  INV_X1 u2_u3_u0_U62 (.A( u2_u3_u0_n126 ) , .ZN( u2_u3_u0_n168 ) );
  AOI211_X1 u2_u3_u0_U63 (.B( u2_u3_u0_n133 ) , .A( u2_u3_u0_n134 ) , .C2( u2_u3_u0_n135 ) , .C1( u2_u3_u0_n136 ) , .ZN( u2_u3_u0_n137 ) );
  OR4_X1 u2_u3_u0_U64 (.ZN( u2_out3_17 ) , .A4( u2_u3_u0_n122 ) , .A2( u2_u3_u0_n123 ) , .A1( u2_u3_u0_n124 ) , .A3( u2_u3_u0_n170 ) );
  AOI21_X1 u2_u3_u0_U65 (.B2( u2_u3_u0_n107 ) , .ZN( u2_u3_u0_n124 ) , .B1( u2_u3_u0_n128 ) , .A( u2_u3_u0_n161 ) );
  INV_X1 u2_u3_u0_U66 (.A( u2_u3_u0_n111 ) , .ZN( u2_u3_u0_n170 ) );
  OR4_X1 u2_u3_u0_U67 (.ZN( u2_out3_31 ) , .A4( u2_u3_u0_n155 ) , .A2( u2_u3_u0_n156 ) , .A1( u2_u3_u0_n157 ) , .A3( u2_u3_u0_n173 ) );
  AOI21_X1 u2_u3_u0_U68 (.A( u2_u3_u0_n138 ) , .B2( u2_u3_u0_n139 ) , .B1( u2_u3_u0_n140 ) , .ZN( u2_u3_u0_n157 ) );
  AOI21_X1 u2_u3_u0_U69 (.B2( u2_u3_u0_n141 ) , .B1( u2_u3_u0_n142 ) , .ZN( u2_u3_u0_n156 ) , .A( u2_u3_u0_n161 ) );
  AOI21_X1 u2_u3_u0_U7 (.B1( u2_u3_u0_n114 ) , .ZN( u2_u3_u0_n115 ) , .B2( u2_u3_u0_n129 ) , .A( u2_u3_u0_n161 ) );
  INV_X1 u2_u3_u0_U70 (.ZN( u2_u3_u0_n174 ) , .A( u2_u3_u0_n89 ) );
  AOI211_X1 u2_u3_u0_U71 (.B( u2_u3_u0_n104 ) , .A( u2_u3_u0_n105 ) , .ZN( u2_u3_u0_n106 ) , .C2( u2_u3_u0_n113 ) , .C1( u2_u3_u0_n160 ) );
  AOI211_X1 u2_u3_u0_U72 (.B( u2_u3_u0_n115 ) , .A( u2_u3_u0_n116 ) , .C2( u2_u3_u0_n117 ) , .C1( u2_u3_u0_n118 ) , .ZN( u2_u3_u0_n119 ) );
  NAND2_X1 u2_u3_u0_U73 (.A2( u2_u3_u0_n100 ) , .ZN( u2_u3_u0_n131 ) , .A1( u2_u3_u0_n92 ) );
  NAND2_X1 u2_u3_u0_U74 (.A1( u2_u3_u0_n100 ) , .A2( u2_u3_u0_n103 ) , .ZN( u2_u3_u0_n125 ) );
  NAND2_X1 u2_u3_u0_U75 (.A2( u2_u3_u0_n100 ) , .A1( u2_u3_u0_n101 ) , .ZN( u2_u3_u0_n139 ) );
  NOR2_X1 u2_u3_u0_U76 (.A2( u2_u3_X_3 ) , .A1( u2_u3_X_6 ) , .ZN( u2_u3_u0_n94 ) );
  INV_X1 u2_u3_u0_U77 (.A( u2_u3_X_3 ) , .ZN( u2_u3_u0_n162 ) );
  NOR2_X1 u2_u3_u0_U78 (.A1( u2_u3_u0_n163 ) , .A2( u2_u3_u0_n164 ) , .ZN( u2_u3_u0_n95 ) );
  OAI221_X1 u2_u3_u0_U79 (.C1( u2_u3_u0_n121 ) , .ZN( u2_u3_u0_n122 ) , .B2( u2_u3_u0_n127 ) , .A( u2_u3_u0_n143 ) , .B1( u2_u3_u0_n144 ) , .C2( u2_u3_u0_n147 ) );
  AND2_X1 u2_u3_u0_U8 (.A1( u2_u3_u0_n114 ) , .A2( u2_u3_u0_n121 ) , .ZN( u2_u3_u0_n146 ) );
  AOI21_X1 u2_u3_u0_U80 (.B1( u2_u3_u0_n132 ) , .ZN( u2_u3_u0_n133 ) , .A( u2_u3_u0_n144 ) , .B2( u2_u3_u0_n166 ) );
  OAI22_X1 u2_u3_u0_U81 (.ZN( u2_u3_u0_n105 ) , .A2( u2_u3_u0_n132 ) , .B1( u2_u3_u0_n146 ) , .A1( u2_u3_u0_n147 ) , .B2( u2_u3_u0_n161 ) );
  NAND2_X1 u2_u3_u0_U82 (.ZN( u2_u3_u0_n110 ) , .A2( u2_u3_u0_n132 ) , .A1( u2_u3_u0_n145 ) );
  INV_X1 u2_u3_u0_U83 (.A( u2_u3_u0_n119 ) , .ZN( u2_u3_u0_n167 ) );
  NAND2_X1 u2_u3_u0_U84 (.ZN( u2_u3_u0_n148 ) , .A1( u2_u3_u0_n93 ) , .A2( u2_u3_u0_n95 ) );
  NAND2_X1 u2_u3_u0_U85 (.A1( u2_u3_u0_n100 ) , .ZN( u2_u3_u0_n129 ) , .A2( u2_u3_u0_n95 ) );
  NAND2_X1 u2_u3_u0_U86 (.A1( u2_u3_u0_n102 ) , .ZN( u2_u3_u0_n128 ) , .A2( u2_u3_u0_n95 ) );
  NAND2_X1 u2_u3_u0_U87 (.ZN( u2_u3_u0_n142 ) , .A1( u2_u3_u0_n94 ) , .A2( u2_u3_u0_n95 ) );
  NAND3_X1 u2_u3_u0_U88 (.ZN( u2_out3_23 ) , .A3( u2_u3_u0_n137 ) , .A1( u2_u3_u0_n168 ) , .A2( u2_u3_u0_n171 ) );
  NAND3_X1 u2_u3_u0_U89 (.A3( u2_u3_u0_n127 ) , .A2( u2_u3_u0_n128 ) , .ZN( u2_u3_u0_n135 ) , .A1( u2_u3_u0_n150 ) );
  AND2_X1 u2_u3_u0_U9 (.A1( u2_u3_u0_n131 ) , .ZN( u2_u3_u0_n141 ) , .A2( u2_u3_u0_n150 ) );
  NAND3_X1 u2_u3_u0_U90 (.ZN( u2_u3_u0_n117 ) , .A3( u2_u3_u0_n132 ) , .A2( u2_u3_u0_n139 ) , .A1( u2_u3_u0_n148 ) );
  NAND3_X1 u2_u3_u0_U91 (.ZN( u2_u3_u0_n109 ) , .A2( u2_u3_u0_n114 ) , .A3( u2_u3_u0_n140 ) , .A1( u2_u3_u0_n149 ) );
  NAND3_X1 u2_u3_u0_U92 (.ZN( u2_out3_9 ) , .A3( u2_u3_u0_n106 ) , .A2( u2_u3_u0_n171 ) , .A1( u2_u3_u0_n174 ) );
  NAND3_X1 u2_u3_u0_U93 (.A2( u2_u3_u0_n128 ) , .A1( u2_u3_u0_n132 ) , .A3( u2_u3_u0_n146 ) , .ZN( u2_u3_u0_n97 ) );
  NOR2_X1 u2_u3_u1_U10 (.A1( u2_u3_u1_n112 ) , .A2( u2_u3_u1_n116 ) , .ZN( u2_u3_u1_n118 ) );
  NAND3_X1 u2_u3_u1_U100 (.ZN( u2_u3_u1_n113 ) , .A1( u2_u3_u1_n120 ) , .A3( u2_u3_u1_n133 ) , .A2( u2_u3_u1_n155 ) );
  OAI21_X1 u2_u3_u1_U11 (.ZN( u2_u3_u1_n101 ) , .B1( u2_u3_u1_n141 ) , .A( u2_u3_u1_n146 ) , .B2( u2_u3_u1_n183 ) );
  AOI21_X1 u2_u3_u1_U12 (.B2( u2_u3_u1_n155 ) , .B1( u2_u3_u1_n156 ) , .ZN( u2_u3_u1_n157 ) , .A( u2_u3_u1_n174 ) );
  NAND2_X1 u2_u3_u1_U13 (.ZN( u2_u3_u1_n140 ) , .A2( u2_u3_u1_n150 ) , .A1( u2_u3_u1_n155 ) );
  NAND2_X1 u2_u3_u1_U14 (.A1( u2_u3_u1_n131 ) , .ZN( u2_u3_u1_n147 ) , .A2( u2_u3_u1_n153 ) );
  INV_X1 u2_u3_u1_U15 (.A( u2_u3_u1_n139 ) , .ZN( u2_u3_u1_n174 ) );
  OR4_X1 u2_u3_u1_U16 (.A4( u2_u3_u1_n106 ) , .A3( u2_u3_u1_n107 ) , .ZN( u2_u3_u1_n108 ) , .A1( u2_u3_u1_n117 ) , .A2( u2_u3_u1_n184 ) );
  AOI21_X1 u2_u3_u1_U17 (.ZN( u2_u3_u1_n106 ) , .A( u2_u3_u1_n112 ) , .B1( u2_u3_u1_n154 ) , .B2( u2_u3_u1_n156 ) );
  INV_X1 u2_u3_u1_U18 (.A( u2_u3_u1_n101 ) , .ZN( u2_u3_u1_n184 ) );
  AOI21_X1 u2_u3_u1_U19 (.ZN( u2_u3_u1_n107 ) , .B1( u2_u3_u1_n134 ) , .B2( u2_u3_u1_n149 ) , .A( u2_u3_u1_n174 ) );
  INV_X1 u2_u3_u1_U20 (.A( u2_u3_u1_n112 ) , .ZN( u2_u3_u1_n171 ) );
  NAND2_X1 u2_u3_u1_U21 (.ZN( u2_u3_u1_n141 ) , .A1( u2_u3_u1_n153 ) , .A2( u2_u3_u1_n156 ) );
  AND2_X1 u2_u3_u1_U22 (.A1( u2_u3_u1_n123 ) , .ZN( u2_u3_u1_n134 ) , .A2( u2_u3_u1_n161 ) );
  NAND2_X1 u2_u3_u1_U23 (.A2( u2_u3_u1_n115 ) , .A1( u2_u3_u1_n116 ) , .ZN( u2_u3_u1_n148 ) );
  NAND2_X1 u2_u3_u1_U24 (.A2( u2_u3_u1_n133 ) , .A1( u2_u3_u1_n135 ) , .ZN( u2_u3_u1_n159 ) );
  NAND2_X1 u2_u3_u1_U25 (.A2( u2_u3_u1_n115 ) , .A1( u2_u3_u1_n120 ) , .ZN( u2_u3_u1_n132 ) );
  INV_X1 u2_u3_u1_U26 (.A( u2_u3_u1_n154 ) , .ZN( u2_u3_u1_n178 ) );
  INV_X1 u2_u3_u1_U27 (.A( u2_u3_u1_n151 ) , .ZN( u2_u3_u1_n183 ) );
  AND2_X1 u2_u3_u1_U28 (.A1( u2_u3_u1_n129 ) , .A2( u2_u3_u1_n133 ) , .ZN( u2_u3_u1_n149 ) );
  INV_X1 u2_u3_u1_U29 (.A( u2_u3_u1_n131 ) , .ZN( u2_u3_u1_n180 ) );
  INV_X1 u2_u3_u1_U3 (.A( u2_u3_u1_n159 ) , .ZN( u2_u3_u1_n182 ) );
  AOI221_X1 u2_u3_u1_U30 (.B1( u2_u3_u1_n140 ) , .ZN( u2_u3_u1_n167 ) , .B2( u2_u3_u1_n172 ) , .C2( u2_u3_u1_n175 ) , .C1( u2_u3_u1_n178 ) , .A( u2_u3_u1_n188 ) );
  INV_X1 u2_u3_u1_U31 (.ZN( u2_u3_u1_n188 ) , .A( u2_u3_u1_n97 ) );
  AOI211_X1 u2_u3_u1_U32 (.A( u2_u3_u1_n118 ) , .C1( u2_u3_u1_n132 ) , .C2( u2_u3_u1_n139 ) , .B( u2_u3_u1_n96 ) , .ZN( u2_u3_u1_n97 ) );
  AOI21_X1 u2_u3_u1_U33 (.B2( u2_u3_u1_n121 ) , .B1( u2_u3_u1_n135 ) , .A( u2_u3_u1_n152 ) , .ZN( u2_u3_u1_n96 ) );
  OAI221_X1 u2_u3_u1_U34 (.A( u2_u3_u1_n119 ) , .C2( u2_u3_u1_n129 ) , .ZN( u2_u3_u1_n138 ) , .B2( u2_u3_u1_n152 ) , .C1( u2_u3_u1_n174 ) , .B1( u2_u3_u1_n187 ) );
  INV_X1 u2_u3_u1_U35 (.A( u2_u3_u1_n148 ) , .ZN( u2_u3_u1_n187 ) );
  AOI211_X1 u2_u3_u1_U36 (.B( u2_u3_u1_n117 ) , .A( u2_u3_u1_n118 ) , .ZN( u2_u3_u1_n119 ) , .C2( u2_u3_u1_n146 ) , .C1( u2_u3_u1_n159 ) );
  NOR2_X1 u2_u3_u1_U37 (.A1( u2_u3_u1_n168 ) , .A2( u2_u3_u1_n176 ) , .ZN( u2_u3_u1_n98 ) );
  NAND2_X1 u2_u3_u1_U38 (.A1( u2_u3_u1_n128 ) , .ZN( u2_u3_u1_n146 ) , .A2( u2_u3_u1_n160 ) );
  NAND2_X1 u2_u3_u1_U39 (.A2( u2_u3_u1_n112 ) , .ZN( u2_u3_u1_n139 ) , .A1( u2_u3_u1_n152 ) );
  AOI221_X1 u2_u3_u1_U4 (.A( u2_u3_u1_n138 ) , .C2( u2_u3_u1_n139 ) , .C1( u2_u3_u1_n140 ) , .B2( u2_u3_u1_n141 ) , .ZN( u2_u3_u1_n142 ) , .B1( u2_u3_u1_n175 ) );
  NAND2_X1 u2_u3_u1_U40 (.A1( u2_u3_u1_n105 ) , .ZN( u2_u3_u1_n156 ) , .A2( u2_u3_u1_n99 ) );
  NOR2_X1 u2_u3_u1_U41 (.ZN( u2_u3_u1_n117 ) , .A1( u2_u3_u1_n121 ) , .A2( u2_u3_u1_n160 ) );
  OAI21_X1 u2_u3_u1_U42 (.B2( u2_u3_u1_n123 ) , .ZN( u2_u3_u1_n145 ) , .B1( u2_u3_u1_n160 ) , .A( u2_u3_u1_n185 ) );
  INV_X1 u2_u3_u1_U43 (.A( u2_u3_u1_n122 ) , .ZN( u2_u3_u1_n185 ) );
  AOI21_X1 u2_u3_u1_U44 (.B2( u2_u3_u1_n120 ) , .B1( u2_u3_u1_n121 ) , .ZN( u2_u3_u1_n122 ) , .A( u2_u3_u1_n128 ) );
  AOI21_X1 u2_u3_u1_U45 (.A( u2_u3_u1_n128 ) , .B2( u2_u3_u1_n129 ) , .ZN( u2_u3_u1_n130 ) , .B1( u2_u3_u1_n150 ) );
  NAND2_X1 u2_u3_u1_U46 (.ZN( u2_u3_u1_n112 ) , .A1( u2_u3_u1_n169 ) , .A2( u2_u3_u1_n170 ) );
  NAND2_X1 u2_u3_u1_U47 (.ZN( u2_u3_u1_n129 ) , .A2( u2_u3_u1_n95 ) , .A1( u2_u3_u1_n98 ) );
  NAND2_X1 u2_u3_u1_U48 (.A1( u2_u3_u1_n102 ) , .ZN( u2_u3_u1_n154 ) , .A2( u2_u3_u1_n99 ) );
  NAND2_X1 u2_u3_u1_U49 (.A2( u2_u3_u1_n100 ) , .ZN( u2_u3_u1_n135 ) , .A1( u2_u3_u1_n99 ) );
  AOI211_X1 u2_u3_u1_U5 (.ZN( u2_u3_u1_n124 ) , .A( u2_u3_u1_n138 ) , .C2( u2_u3_u1_n139 ) , .B( u2_u3_u1_n145 ) , .C1( u2_u3_u1_n147 ) );
  AOI21_X1 u2_u3_u1_U50 (.A( u2_u3_u1_n152 ) , .B2( u2_u3_u1_n153 ) , .B1( u2_u3_u1_n154 ) , .ZN( u2_u3_u1_n158 ) );
  INV_X1 u2_u3_u1_U51 (.A( u2_u3_u1_n160 ) , .ZN( u2_u3_u1_n175 ) );
  NAND2_X1 u2_u3_u1_U52 (.A1( u2_u3_u1_n100 ) , .ZN( u2_u3_u1_n116 ) , .A2( u2_u3_u1_n95 ) );
  NAND2_X1 u2_u3_u1_U53 (.A1( u2_u3_u1_n102 ) , .ZN( u2_u3_u1_n131 ) , .A2( u2_u3_u1_n95 ) );
  NAND2_X1 u2_u3_u1_U54 (.A2( u2_u3_u1_n104 ) , .ZN( u2_u3_u1_n121 ) , .A1( u2_u3_u1_n98 ) );
  NAND2_X1 u2_u3_u1_U55 (.A1( u2_u3_u1_n103 ) , .ZN( u2_u3_u1_n153 ) , .A2( u2_u3_u1_n98 ) );
  NAND2_X1 u2_u3_u1_U56 (.A2( u2_u3_u1_n104 ) , .A1( u2_u3_u1_n105 ) , .ZN( u2_u3_u1_n133 ) );
  NAND2_X1 u2_u3_u1_U57 (.ZN( u2_u3_u1_n150 ) , .A2( u2_u3_u1_n98 ) , .A1( u2_u3_u1_n99 ) );
  NAND2_X1 u2_u3_u1_U58 (.A1( u2_u3_u1_n105 ) , .ZN( u2_u3_u1_n155 ) , .A2( u2_u3_u1_n95 ) );
  OAI21_X1 u2_u3_u1_U59 (.ZN( u2_u3_u1_n109 ) , .B1( u2_u3_u1_n129 ) , .B2( u2_u3_u1_n160 ) , .A( u2_u3_u1_n167 ) );
  AOI22_X1 u2_u3_u1_U6 (.B2( u2_u3_u1_n113 ) , .A2( u2_u3_u1_n114 ) , .ZN( u2_u3_u1_n125 ) , .A1( u2_u3_u1_n171 ) , .B1( u2_u3_u1_n173 ) );
  NAND2_X1 u2_u3_u1_U60 (.A2( u2_u3_u1_n100 ) , .A1( u2_u3_u1_n103 ) , .ZN( u2_u3_u1_n120 ) );
  NAND2_X1 u2_u3_u1_U61 (.A1( u2_u3_u1_n102 ) , .A2( u2_u3_u1_n104 ) , .ZN( u2_u3_u1_n115 ) );
  NAND2_X1 u2_u3_u1_U62 (.A2( u2_u3_u1_n100 ) , .A1( u2_u3_u1_n104 ) , .ZN( u2_u3_u1_n151 ) );
  NAND2_X1 u2_u3_u1_U63 (.A2( u2_u3_u1_n103 ) , .A1( u2_u3_u1_n105 ) , .ZN( u2_u3_u1_n161 ) );
  INV_X1 u2_u3_u1_U64 (.A( u2_u3_u1_n152 ) , .ZN( u2_u3_u1_n173 ) );
  INV_X1 u2_u3_u1_U65 (.A( u2_u3_u1_n128 ) , .ZN( u2_u3_u1_n172 ) );
  NAND2_X1 u2_u3_u1_U66 (.A2( u2_u3_u1_n102 ) , .A1( u2_u3_u1_n103 ) , .ZN( u2_u3_u1_n123 ) );
  AOI211_X1 u2_u3_u1_U67 (.B( u2_u3_u1_n162 ) , .A( u2_u3_u1_n163 ) , .C2( u2_u3_u1_n164 ) , .ZN( u2_u3_u1_n165 ) , .C1( u2_u3_u1_n171 ) );
  AOI21_X1 u2_u3_u1_U68 (.A( u2_u3_u1_n160 ) , .B2( u2_u3_u1_n161 ) , .ZN( u2_u3_u1_n162 ) , .B1( u2_u3_u1_n182 ) );
  OR2_X1 u2_u3_u1_U69 (.A2( u2_u3_u1_n157 ) , .A1( u2_u3_u1_n158 ) , .ZN( u2_u3_u1_n163 ) );
  NAND2_X1 u2_u3_u1_U7 (.ZN( u2_u3_u1_n114 ) , .A1( u2_u3_u1_n134 ) , .A2( u2_u3_u1_n156 ) );
  NOR2_X1 u2_u3_u1_U70 (.A2( u2_u3_X_7 ) , .A1( u2_u3_X_8 ) , .ZN( u2_u3_u1_n95 ) );
  NOR2_X1 u2_u3_u1_U71 (.A1( u2_u3_X_12 ) , .A2( u2_u3_X_9 ) , .ZN( u2_u3_u1_n100 ) );
  NOR2_X1 u2_u3_u1_U72 (.A2( u2_u3_X_8 ) , .A1( u2_u3_u1_n177 ) , .ZN( u2_u3_u1_n99 ) );
  NOR2_X1 u2_u3_u1_U73 (.A2( u2_u3_X_12 ) , .ZN( u2_u3_u1_n102 ) , .A1( u2_u3_u1_n176 ) );
  NOR2_X1 u2_u3_u1_U74 (.A2( u2_u3_X_9 ) , .ZN( u2_u3_u1_n105 ) , .A1( u2_u3_u1_n168 ) );
  NAND2_X1 u2_u3_u1_U75 (.A1( u2_u3_X_10 ) , .ZN( u2_u3_u1_n160 ) , .A2( u2_u3_u1_n169 ) );
  NAND2_X1 u2_u3_u1_U76 (.A2( u2_u3_X_10 ) , .A1( u2_u3_X_11 ) , .ZN( u2_u3_u1_n152 ) );
  NAND2_X1 u2_u3_u1_U77 (.A1( u2_u3_X_11 ) , .ZN( u2_u3_u1_n128 ) , .A2( u2_u3_u1_n170 ) );
  AND2_X1 u2_u3_u1_U78 (.A2( u2_u3_X_7 ) , .A1( u2_u3_X_8 ) , .ZN( u2_u3_u1_n104 ) );
  AND2_X1 u2_u3_u1_U79 (.A1( u2_u3_X_8 ) , .ZN( u2_u3_u1_n103 ) , .A2( u2_u3_u1_n177 ) );
  AOI22_X1 u2_u3_u1_U8 (.B2( u2_u3_u1_n136 ) , .A2( u2_u3_u1_n137 ) , .ZN( u2_u3_u1_n143 ) , .A1( u2_u3_u1_n171 ) , .B1( u2_u3_u1_n173 ) );
  INV_X1 u2_u3_u1_U80 (.A( u2_u3_X_10 ) , .ZN( u2_u3_u1_n170 ) );
  INV_X1 u2_u3_u1_U81 (.A( u2_u3_X_9 ) , .ZN( u2_u3_u1_n176 ) );
  INV_X1 u2_u3_u1_U82 (.A( u2_u3_X_11 ) , .ZN( u2_u3_u1_n169 ) );
  INV_X1 u2_u3_u1_U83 (.A( u2_u3_X_12 ) , .ZN( u2_u3_u1_n168 ) );
  INV_X1 u2_u3_u1_U84 (.A( u2_u3_X_7 ) , .ZN( u2_u3_u1_n177 ) );
  NAND4_X1 u2_u3_u1_U85 (.ZN( u2_out3_28 ) , .A4( u2_u3_u1_n124 ) , .A3( u2_u3_u1_n125 ) , .A2( u2_u3_u1_n126 ) , .A1( u2_u3_u1_n127 ) );
  OAI21_X1 u2_u3_u1_U86 (.ZN( u2_u3_u1_n127 ) , .B2( u2_u3_u1_n139 ) , .B1( u2_u3_u1_n175 ) , .A( u2_u3_u1_n183 ) );
  OAI21_X1 u2_u3_u1_U87 (.ZN( u2_u3_u1_n126 ) , .B2( u2_u3_u1_n140 ) , .A( u2_u3_u1_n146 ) , .B1( u2_u3_u1_n178 ) );
  NAND4_X1 u2_u3_u1_U88 (.ZN( u2_out3_18 ) , .A4( u2_u3_u1_n165 ) , .A3( u2_u3_u1_n166 ) , .A1( u2_u3_u1_n167 ) , .A2( u2_u3_u1_n186 ) );
  AOI22_X1 u2_u3_u1_U89 (.B2( u2_u3_u1_n146 ) , .B1( u2_u3_u1_n147 ) , .A2( u2_u3_u1_n148 ) , .ZN( u2_u3_u1_n166 ) , .A1( u2_u3_u1_n172 ) );
  INV_X1 u2_u3_u1_U9 (.A( u2_u3_u1_n147 ) , .ZN( u2_u3_u1_n181 ) );
  INV_X1 u2_u3_u1_U90 (.A( u2_u3_u1_n145 ) , .ZN( u2_u3_u1_n186 ) );
  NAND4_X1 u2_u3_u1_U91 (.ZN( u2_out3_2 ) , .A4( u2_u3_u1_n142 ) , .A3( u2_u3_u1_n143 ) , .A2( u2_u3_u1_n144 ) , .A1( u2_u3_u1_n179 ) );
  OAI21_X1 u2_u3_u1_U92 (.B2( u2_u3_u1_n132 ) , .ZN( u2_u3_u1_n144 ) , .A( u2_u3_u1_n146 ) , .B1( u2_u3_u1_n180 ) );
  INV_X1 u2_u3_u1_U93 (.A( u2_u3_u1_n130 ) , .ZN( u2_u3_u1_n179 ) );
  OR4_X1 u2_u3_u1_U94 (.ZN( u2_out3_13 ) , .A4( u2_u3_u1_n108 ) , .A3( u2_u3_u1_n109 ) , .A2( u2_u3_u1_n110 ) , .A1( u2_u3_u1_n111 ) );
  AOI21_X1 u2_u3_u1_U95 (.ZN( u2_u3_u1_n111 ) , .A( u2_u3_u1_n128 ) , .B2( u2_u3_u1_n131 ) , .B1( u2_u3_u1_n135 ) );
  AOI21_X1 u2_u3_u1_U96 (.ZN( u2_u3_u1_n110 ) , .A( u2_u3_u1_n116 ) , .B1( u2_u3_u1_n152 ) , .B2( u2_u3_u1_n160 ) );
  NAND3_X1 u2_u3_u1_U97 (.A3( u2_u3_u1_n149 ) , .A2( u2_u3_u1_n150 ) , .A1( u2_u3_u1_n151 ) , .ZN( u2_u3_u1_n164 ) );
  NAND3_X1 u2_u3_u1_U98 (.A3( u2_u3_u1_n134 ) , .A2( u2_u3_u1_n135 ) , .ZN( u2_u3_u1_n136 ) , .A1( u2_u3_u1_n151 ) );
  NAND3_X1 u2_u3_u1_U99 (.A1( u2_u3_u1_n133 ) , .ZN( u2_u3_u1_n137 ) , .A2( u2_u3_u1_n154 ) , .A3( u2_u3_u1_n181 ) );
  AND3_X1 u2_u3_u7_U10 (.A3( u2_u3_u7_n110 ) , .A2( u2_u3_u7_n127 ) , .A1( u2_u3_u7_n132 ) , .ZN( u2_u3_u7_n92 ) );
  OAI21_X1 u2_u3_u7_U11 (.A( u2_u3_u7_n161 ) , .B1( u2_u3_u7_n168 ) , .B2( u2_u3_u7_n173 ) , .ZN( u2_u3_u7_n91 ) );
  AOI211_X1 u2_u3_u7_U12 (.A( u2_u3_u7_n117 ) , .ZN( u2_u3_u7_n118 ) , .C2( u2_u3_u7_n126 ) , .C1( u2_u3_u7_n177 ) , .B( u2_u3_u7_n180 ) );
  OAI22_X1 u2_u3_u7_U13 (.B1( u2_u3_u7_n115 ) , .ZN( u2_u3_u7_n117 ) , .A2( u2_u3_u7_n133 ) , .A1( u2_u3_u7_n137 ) , .B2( u2_u3_u7_n162 ) );
  INV_X1 u2_u3_u7_U14 (.A( u2_u3_u7_n116 ) , .ZN( u2_u3_u7_n180 ) );
  NOR3_X1 u2_u3_u7_U15 (.ZN( u2_u3_u7_n115 ) , .A3( u2_u3_u7_n145 ) , .A2( u2_u3_u7_n168 ) , .A1( u2_u3_u7_n169 ) );
  OAI211_X1 u2_u3_u7_U16 (.B( u2_u3_u7_n122 ) , .A( u2_u3_u7_n123 ) , .C2( u2_u3_u7_n124 ) , .ZN( u2_u3_u7_n154 ) , .C1( u2_u3_u7_n162 ) );
  AOI222_X1 u2_u3_u7_U17 (.ZN( u2_u3_u7_n122 ) , .C2( u2_u3_u7_n126 ) , .C1( u2_u3_u7_n145 ) , .B1( u2_u3_u7_n161 ) , .A2( u2_u3_u7_n165 ) , .B2( u2_u3_u7_n170 ) , .A1( u2_u3_u7_n176 ) );
  INV_X1 u2_u3_u7_U18 (.A( u2_u3_u7_n133 ) , .ZN( u2_u3_u7_n176 ) );
  NOR3_X1 u2_u3_u7_U19 (.A2( u2_u3_u7_n134 ) , .A1( u2_u3_u7_n135 ) , .ZN( u2_u3_u7_n136 ) , .A3( u2_u3_u7_n171 ) );
  NOR2_X1 u2_u3_u7_U20 (.A1( u2_u3_u7_n130 ) , .A2( u2_u3_u7_n134 ) , .ZN( u2_u3_u7_n153 ) );
  INV_X1 u2_u3_u7_U21 (.A( u2_u3_u7_n101 ) , .ZN( u2_u3_u7_n165 ) );
  NOR2_X1 u2_u3_u7_U22 (.ZN( u2_u3_u7_n111 ) , .A2( u2_u3_u7_n134 ) , .A1( u2_u3_u7_n169 ) );
  AOI21_X1 u2_u3_u7_U23 (.ZN( u2_u3_u7_n104 ) , .B2( u2_u3_u7_n112 ) , .B1( u2_u3_u7_n127 ) , .A( u2_u3_u7_n164 ) );
  AOI21_X1 u2_u3_u7_U24 (.ZN( u2_u3_u7_n106 ) , .B1( u2_u3_u7_n133 ) , .B2( u2_u3_u7_n146 ) , .A( u2_u3_u7_n162 ) );
  AOI21_X1 u2_u3_u7_U25 (.A( u2_u3_u7_n101 ) , .ZN( u2_u3_u7_n107 ) , .B2( u2_u3_u7_n128 ) , .B1( u2_u3_u7_n175 ) );
  INV_X1 u2_u3_u7_U26 (.A( u2_u3_u7_n138 ) , .ZN( u2_u3_u7_n171 ) );
  INV_X1 u2_u3_u7_U27 (.A( u2_u3_u7_n131 ) , .ZN( u2_u3_u7_n177 ) );
  INV_X1 u2_u3_u7_U28 (.A( u2_u3_u7_n110 ) , .ZN( u2_u3_u7_n174 ) );
  NAND2_X1 u2_u3_u7_U29 (.A1( u2_u3_u7_n129 ) , .A2( u2_u3_u7_n132 ) , .ZN( u2_u3_u7_n149 ) );
  OAI21_X1 u2_u3_u7_U3 (.ZN( u2_u3_u7_n159 ) , .A( u2_u3_u7_n165 ) , .B2( u2_u3_u7_n171 ) , .B1( u2_u3_u7_n174 ) );
  NAND2_X1 u2_u3_u7_U30 (.A1( u2_u3_u7_n113 ) , .A2( u2_u3_u7_n124 ) , .ZN( u2_u3_u7_n130 ) );
  INV_X1 u2_u3_u7_U31 (.A( u2_u3_u7_n112 ) , .ZN( u2_u3_u7_n173 ) );
  INV_X1 u2_u3_u7_U32 (.A( u2_u3_u7_n128 ) , .ZN( u2_u3_u7_n168 ) );
  INV_X1 u2_u3_u7_U33 (.A( u2_u3_u7_n148 ) , .ZN( u2_u3_u7_n169 ) );
  INV_X1 u2_u3_u7_U34 (.A( u2_u3_u7_n127 ) , .ZN( u2_u3_u7_n179 ) );
  NOR2_X1 u2_u3_u7_U35 (.ZN( u2_u3_u7_n101 ) , .A2( u2_u3_u7_n150 ) , .A1( u2_u3_u7_n156 ) );
  AOI211_X1 u2_u3_u7_U36 (.B( u2_u3_u7_n154 ) , .A( u2_u3_u7_n155 ) , .C1( u2_u3_u7_n156 ) , .ZN( u2_u3_u7_n157 ) , .C2( u2_u3_u7_n172 ) );
  INV_X1 u2_u3_u7_U37 (.A( u2_u3_u7_n153 ) , .ZN( u2_u3_u7_n172 ) );
  AOI211_X1 u2_u3_u7_U38 (.B( u2_u3_u7_n139 ) , .A( u2_u3_u7_n140 ) , .C2( u2_u3_u7_n141 ) , .ZN( u2_u3_u7_n142 ) , .C1( u2_u3_u7_n156 ) );
  NAND4_X1 u2_u3_u7_U39 (.A3( u2_u3_u7_n127 ) , .A2( u2_u3_u7_n128 ) , .A1( u2_u3_u7_n129 ) , .ZN( u2_u3_u7_n141 ) , .A4( u2_u3_u7_n147 ) );
  INV_X1 u2_u3_u7_U4 (.A( u2_u3_u7_n111 ) , .ZN( u2_u3_u7_n170 ) );
  AOI21_X1 u2_u3_u7_U40 (.A( u2_u3_u7_n137 ) , .B1( u2_u3_u7_n138 ) , .ZN( u2_u3_u7_n139 ) , .B2( u2_u3_u7_n146 ) );
  OAI22_X1 u2_u3_u7_U41 (.B1( u2_u3_u7_n136 ) , .ZN( u2_u3_u7_n140 ) , .A1( u2_u3_u7_n153 ) , .B2( u2_u3_u7_n162 ) , .A2( u2_u3_u7_n164 ) );
  AOI21_X1 u2_u3_u7_U42 (.ZN( u2_u3_u7_n123 ) , .B1( u2_u3_u7_n165 ) , .B2( u2_u3_u7_n177 ) , .A( u2_u3_u7_n97 ) );
  AOI21_X1 u2_u3_u7_U43 (.B2( u2_u3_u7_n113 ) , .B1( u2_u3_u7_n124 ) , .A( u2_u3_u7_n125 ) , .ZN( u2_u3_u7_n97 ) );
  INV_X1 u2_u3_u7_U44 (.A( u2_u3_u7_n125 ) , .ZN( u2_u3_u7_n161 ) );
  INV_X1 u2_u3_u7_U45 (.A( u2_u3_u7_n152 ) , .ZN( u2_u3_u7_n162 ) );
  AOI22_X1 u2_u3_u7_U46 (.A2( u2_u3_u7_n114 ) , .ZN( u2_u3_u7_n119 ) , .B1( u2_u3_u7_n130 ) , .A1( u2_u3_u7_n156 ) , .B2( u2_u3_u7_n165 ) );
  NAND2_X1 u2_u3_u7_U47 (.A2( u2_u3_u7_n112 ) , .ZN( u2_u3_u7_n114 ) , .A1( u2_u3_u7_n175 ) );
  AND2_X1 u2_u3_u7_U48 (.ZN( u2_u3_u7_n145 ) , .A2( u2_u3_u7_n98 ) , .A1( u2_u3_u7_n99 ) );
  NOR2_X1 u2_u3_u7_U49 (.ZN( u2_u3_u7_n137 ) , .A1( u2_u3_u7_n150 ) , .A2( u2_u3_u7_n161 ) );
  INV_X1 u2_u3_u7_U5 (.A( u2_u3_u7_n149 ) , .ZN( u2_u3_u7_n175 ) );
  AOI21_X1 u2_u3_u7_U50 (.ZN( u2_u3_u7_n105 ) , .B2( u2_u3_u7_n110 ) , .A( u2_u3_u7_n125 ) , .B1( u2_u3_u7_n147 ) );
  NAND2_X1 u2_u3_u7_U51 (.ZN( u2_u3_u7_n146 ) , .A1( u2_u3_u7_n95 ) , .A2( u2_u3_u7_n98 ) );
  NAND2_X1 u2_u3_u7_U52 (.A2( u2_u3_u7_n103 ) , .ZN( u2_u3_u7_n147 ) , .A1( u2_u3_u7_n93 ) );
  NAND2_X1 u2_u3_u7_U53 (.A1( u2_u3_u7_n103 ) , .ZN( u2_u3_u7_n127 ) , .A2( u2_u3_u7_n99 ) );
  OR2_X1 u2_u3_u7_U54 (.ZN( u2_u3_u7_n126 ) , .A2( u2_u3_u7_n152 ) , .A1( u2_u3_u7_n156 ) );
  NAND2_X1 u2_u3_u7_U55 (.A2( u2_u3_u7_n102 ) , .A1( u2_u3_u7_n103 ) , .ZN( u2_u3_u7_n133 ) );
  NAND2_X1 u2_u3_u7_U56 (.ZN( u2_u3_u7_n112 ) , .A2( u2_u3_u7_n96 ) , .A1( u2_u3_u7_n99 ) );
  NAND2_X1 u2_u3_u7_U57 (.A2( u2_u3_u7_n102 ) , .ZN( u2_u3_u7_n128 ) , .A1( u2_u3_u7_n98 ) );
  NAND2_X1 u2_u3_u7_U58 (.A1( u2_u3_u7_n100 ) , .ZN( u2_u3_u7_n113 ) , .A2( u2_u3_u7_n93 ) );
  NAND2_X1 u2_u3_u7_U59 (.A2( u2_u3_u7_n102 ) , .ZN( u2_u3_u7_n124 ) , .A1( u2_u3_u7_n96 ) );
  INV_X1 u2_u3_u7_U6 (.A( u2_u3_u7_n154 ) , .ZN( u2_u3_u7_n178 ) );
  NAND2_X1 u2_u3_u7_U60 (.ZN( u2_u3_u7_n110 ) , .A1( u2_u3_u7_n95 ) , .A2( u2_u3_u7_n96 ) );
  INV_X1 u2_u3_u7_U61 (.A( u2_u3_u7_n150 ) , .ZN( u2_u3_u7_n164 ) );
  AND2_X1 u2_u3_u7_U62 (.ZN( u2_u3_u7_n134 ) , .A1( u2_u3_u7_n93 ) , .A2( u2_u3_u7_n98 ) );
  NAND2_X1 u2_u3_u7_U63 (.A1( u2_u3_u7_n100 ) , .A2( u2_u3_u7_n102 ) , .ZN( u2_u3_u7_n129 ) );
  NAND2_X1 u2_u3_u7_U64 (.A2( u2_u3_u7_n103 ) , .ZN( u2_u3_u7_n131 ) , .A1( u2_u3_u7_n95 ) );
  NAND2_X1 u2_u3_u7_U65 (.A1( u2_u3_u7_n100 ) , .ZN( u2_u3_u7_n138 ) , .A2( u2_u3_u7_n99 ) );
  NAND2_X1 u2_u3_u7_U66 (.ZN( u2_u3_u7_n132 ) , .A1( u2_u3_u7_n93 ) , .A2( u2_u3_u7_n96 ) );
  NAND2_X1 u2_u3_u7_U67 (.A1( u2_u3_u7_n100 ) , .ZN( u2_u3_u7_n148 ) , .A2( u2_u3_u7_n95 ) );
  NOR2_X1 u2_u3_u7_U68 (.A2( u2_u3_X_47 ) , .ZN( u2_u3_u7_n150 ) , .A1( u2_u3_u7_n163 ) );
  NOR2_X1 u2_u3_u7_U69 (.A2( u2_u3_X_43 ) , .A1( u2_u3_X_44 ) , .ZN( u2_u3_u7_n103 ) );
  AOI211_X1 u2_u3_u7_U7 (.ZN( u2_u3_u7_n116 ) , .A( u2_u3_u7_n155 ) , .C1( u2_u3_u7_n161 ) , .C2( u2_u3_u7_n171 ) , .B( u2_u3_u7_n94 ) );
  NOR2_X1 u2_u3_u7_U70 (.A2( u2_u3_X_48 ) , .A1( u2_u3_u7_n166 ) , .ZN( u2_u3_u7_n95 ) );
  NOR2_X1 u2_u3_u7_U71 (.A2( u2_u3_X_45 ) , .A1( u2_u3_X_48 ) , .ZN( u2_u3_u7_n99 ) );
  NOR2_X1 u2_u3_u7_U72 (.A2( u2_u3_X_44 ) , .A1( u2_u3_u7_n167 ) , .ZN( u2_u3_u7_n98 ) );
  NOR2_X1 u2_u3_u7_U73 (.A2( u2_u3_X_46 ) , .A1( u2_u3_X_47 ) , .ZN( u2_u3_u7_n152 ) );
  AND2_X1 u2_u3_u7_U74 (.A1( u2_u3_X_47 ) , .ZN( u2_u3_u7_n156 ) , .A2( u2_u3_u7_n163 ) );
  NAND2_X1 u2_u3_u7_U75 (.A2( u2_u3_X_46 ) , .A1( u2_u3_X_47 ) , .ZN( u2_u3_u7_n125 ) );
  AND2_X1 u2_u3_u7_U76 (.A2( u2_u3_X_45 ) , .A1( u2_u3_X_48 ) , .ZN( u2_u3_u7_n102 ) );
  AND2_X1 u2_u3_u7_U77 (.A2( u2_u3_X_43 ) , .A1( u2_u3_X_44 ) , .ZN( u2_u3_u7_n96 ) );
  AND2_X1 u2_u3_u7_U78 (.A1( u2_u3_X_44 ) , .ZN( u2_u3_u7_n100 ) , .A2( u2_u3_u7_n167 ) );
  AND2_X1 u2_u3_u7_U79 (.A1( u2_u3_X_48 ) , .A2( u2_u3_u7_n166 ) , .ZN( u2_u3_u7_n93 ) );
  OAI222_X1 u2_u3_u7_U8 (.C2( u2_u3_u7_n101 ) , .B2( u2_u3_u7_n111 ) , .A1( u2_u3_u7_n113 ) , .C1( u2_u3_u7_n146 ) , .A2( u2_u3_u7_n162 ) , .B1( u2_u3_u7_n164 ) , .ZN( u2_u3_u7_n94 ) );
  INV_X1 u2_u3_u7_U80 (.A( u2_u3_X_46 ) , .ZN( u2_u3_u7_n163 ) );
  INV_X1 u2_u3_u7_U81 (.A( u2_u3_X_43 ) , .ZN( u2_u3_u7_n167 ) );
  INV_X1 u2_u3_u7_U82 (.A( u2_u3_X_45 ) , .ZN( u2_u3_u7_n166 ) );
  NAND4_X1 u2_u3_u7_U83 (.ZN( u2_out3_5 ) , .A4( u2_u3_u7_n108 ) , .A3( u2_u3_u7_n109 ) , .A1( u2_u3_u7_n116 ) , .A2( u2_u3_u7_n123 ) );
  AOI22_X1 u2_u3_u7_U84 (.ZN( u2_u3_u7_n109 ) , .A2( u2_u3_u7_n126 ) , .B2( u2_u3_u7_n145 ) , .B1( u2_u3_u7_n156 ) , .A1( u2_u3_u7_n171 ) );
  NOR4_X1 u2_u3_u7_U85 (.A4( u2_u3_u7_n104 ) , .A3( u2_u3_u7_n105 ) , .A2( u2_u3_u7_n106 ) , .A1( u2_u3_u7_n107 ) , .ZN( u2_u3_u7_n108 ) );
  NAND4_X1 u2_u3_u7_U86 (.ZN( u2_out3_27 ) , .A4( u2_u3_u7_n118 ) , .A3( u2_u3_u7_n119 ) , .A2( u2_u3_u7_n120 ) , .A1( u2_u3_u7_n121 ) );
  OAI21_X1 u2_u3_u7_U87 (.ZN( u2_u3_u7_n121 ) , .B2( u2_u3_u7_n145 ) , .A( u2_u3_u7_n150 ) , .B1( u2_u3_u7_n174 ) );
  OAI21_X1 u2_u3_u7_U88 (.ZN( u2_u3_u7_n120 ) , .A( u2_u3_u7_n161 ) , .B2( u2_u3_u7_n170 ) , .B1( u2_u3_u7_n179 ) );
  NAND4_X1 u2_u3_u7_U89 (.ZN( u2_out3_21 ) , .A4( u2_u3_u7_n157 ) , .A3( u2_u3_u7_n158 ) , .A2( u2_u3_u7_n159 ) , .A1( u2_u3_u7_n160 ) );
  OAI221_X1 u2_u3_u7_U9 (.C1( u2_u3_u7_n101 ) , .C2( u2_u3_u7_n147 ) , .ZN( u2_u3_u7_n155 ) , .B2( u2_u3_u7_n162 ) , .A( u2_u3_u7_n91 ) , .B1( u2_u3_u7_n92 ) );
  OAI21_X1 u2_u3_u7_U90 (.B1( u2_u3_u7_n145 ) , .ZN( u2_u3_u7_n160 ) , .A( u2_u3_u7_n161 ) , .B2( u2_u3_u7_n177 ) );
  AOI22_X1 u2_u3_u7_U91 (.B2( u2_u3_u7_n149 ) , .B1( u2_u3_u7_n150 ) , .A2( u2_u3_u7_n151 ) , .A1( u2_u3_u7_n152 ) , .ZN( u2_u3_u7_n158 ) );
  NAND4_X1 u2_u3_u7_U92 (.ZN( u2_out3_15 ) , .A4( u2_u3_u7_n142 ) , .A3( u2_u3_u7_n143 ) , .A2( u2_u3_u7_n144 ) , .A1( u2_u3_u7_n178 ) );
  OR2_X1 u2_u3_u7_U93 (.A2( u2_u3_u7_n125 ) , .A1( u2_u3_u7_n129 ) , .ZN( u2_u3_u7_n144 ) );
  AOI22_X1 u2_u3_u7_U94 (.A2( u2_u3_u7_n126 ) , .ZN( u2_u3_u7_n143 ) , .B2( u2_u3_u7_n165 ) , .B1( u2_u3_u7_n173 ) , .A1( u2_u3_u7_n174 ) );
  NAND3_X1 u2_u3_u7_U95 (.A3( u2_u3_u7_n146 ) , .A2( u2_u3_u7_n147 ) , .A1( u2_u3_u7_n148 ) , .ZN( u2_u3_u7_n151 ) );
  NAND3_X1 u2_u3_u7_U96 (.A3( u2_u3_u7_n131 ) , .A2( u2_u3_u7_n132 ) , .A1( u2_u3_u7_n133 ) , .ZN( u2_u3_u7_n135 ) );
  XOR2_X1 u2_u5_U26 (.B( u2_K6_30 ) , .A( u2_R4_21 ) , .Z( u2_u5_X_30 ) );
  XOR2_X1 u2_u5_U28 (.B( u2_K6_29 ) , .A( u2_R4_20 ) , .Z( u2_u5_X_29 ) );
  XOR2_X1 u2_u5_U29 (.B( u2_K6_28 ) , .A( u2_R4_19 ) , .Z( u2_u5_X_28 ) );
  XOR2_X1 u2_u5_U30 (.B( u2_K6_27 ) , .A( u2_R4_18 ) , .Z( u2_u5_X_27 ) );
  XOR2_X1 u2_u5_U31 (.B( u2_K6_26 ) , .A( u2_R4_17 ) , .Z( u2_u5_X_26 ) );
  XOR2_X1 u2_u5_U32 (.B( u2_K6_25 ) , .A( u2_R4_16 ) , .Z( u2_u5_X_25 ) );
  OAI22_X1 u2_u5_u4_U10 (.B2( u2_u5_u4_n135 ) , .ZN( u2_u5_u4_n137 ) , .B1( u2_u5_u4_n153 ) , .A1( u2_u5_u4_n155 ) , .A2( u2_u5_u4_n171 ) );
  AND3_X1 u2_u5_u4_U11 (.A2( u2_u5_u4_n134 ) , .ZN( u2_u5_u4_n135 ) , .A3( u2_u5_u4_n145 ) , .A1( u2_u5_u4_n157 ) );
  NAND2_X1 u2_u5_u4_U12 (.ZN( u2_u5_u4_n132 ) , .A2( u2_u5_u4_n170 ) , .A1( u2_u5_u4_n173 ) );
  AOI21_X1 u2_u5_u4_U13 (.B2( u2_u5_u4_n160 ) , .B1( u2_u5_u4_n161 ) , .ZN( u2_u5_u4_n162 ) , .A( u2_u5_u4_n170 ) );
  AOI21_X1 u2_u5_u4_U14 (.ZN( u2_u5_u4_n107 ) , .B2( u2_u5_u4_n143 ) , .A( u2_u5_u4_n174 ) , .B1( u2_u5_u4_n184 ) );
  AOI21_X1 u2_u5_u4_U15 (.B2( u2_u5_u4_n158 ) , .B1( u2_u5_u4_n159 ) , .ZN( u2_u5_u4_n163 ) , .A( u2_u5_u4_n174 ) );
  AOI21_X1 u2_u5_u4_U16 (.A( u2_u5_u4_n153 ) , .B2( u2_u5_u4_n154 ) , .B1( u2_u5_u4_n155 ) , .ZN( u2_u5_u4_n165 ) );
  AOI21_X1 u2_u5_u4_U17 (.A( u2_u5_u4_n156 ) , .B2( u2_u5_u4_n157 ) , .ZN( u2_u5_u4_n164 ) , .B1( u2_u5_u4_n184 ) );
  INV_X1 u2_u5_u4_U18 (.A( u2_u5_u4_n138 ) , .ZN( u2_u5_u4_n170 ) );
  AND2_X1 u2_u5_u4_U19 (.A2( u2_u5_u4_n120 ) , .ZN( u2_u5_u4_n155 ) , .A1( u2_u5_u4_n160 ) );
  INV_X1 u2_u5_u4_U20 (.A( u2_u5_u4_n156 ) , .ZN( u2_u5_u4_n175 ) );
  NAND2_X1 u2_u5_u4_U21 (.A2( u2_u5_u4_n118 ) , .ZN( u2_u5_u4_n131 ) , .A1( u2_u5_u4_n147 ) );
  NAND2_X1 u2_u5_u4_U22 (.A1( u2_u5_u4_n119 ) , .A2( u2_u5_u4_n120 ) , .ZN( u2_u5_u4_n130 ) );
  NAND2_X1 u2_u5_u4_U23 (.ZN( u2_u5_u4_n117 ) , .A2( u2_u5_u4_n118 ) , .A1( u2_u5_u4_n148 ) );
  NAND2_X1 u2_u5_u4_U24 (.ZN( u2_u5_u4_n129 ) , .A1( u2_u5_u4_n134 ) , .A2( u2_u5_u4_n148 ) );
  AND3_X1 u2_u5_u4_U25 (.A1( u2_u5_u4_n119 ) , .A2( u2_u5_u4_n143 ) , .A3( u2_u5_u4_n154 ) , .ZN( u2_u5_u4_n161 ) );
  AND2_X1 u2_u5_u4_U26 (.A1( u2_u5_u4_n145 ) , .A2( u2_u5_u4_n147 ) , .ZN( u2_u5_u4_n159 ) );
  OR3_X1 u2_u5_u4_U27 (.A3( u2_u5_u4_n114 ) , .A2( u2_u5_u4_n115 ) , .A1( u2_u5_u4_n116 ) , .ZN( u2_u5_u4_n136 ) );
  AOI21_X1 u2_u5_u4_U28 (.A( u2_u5_u4_n113 ) , .ZN( u2_u5_u4_n116 ) , .B2( u2_u5_u4_n173 ) , .B1( u2_u5_u4_n174 ) );
  AOI21_X1 u2_u5_u4_U29 (.ZN( u2_u5_u4_n115 ) , .B2( u2_u5_u4_n145 ) , .B1( u2_u5_u4_n146 ) , .A( u2_u5_u4_n156 ) );
  NOR2_X1 u2_u5_u4_U3 (.ZN( u2_u5_u4_n121 ) , .A1( u2_u5_u4_n181 ) , .A2( u2_u5_u4_n182 ) );
  OAI22_X1 u2_u5_u4_U30 (.ZN( u2_u5_u4_n114 ) , .A2( u2_u5_u4_n121 ) , .B1( u2_u5_u4_n160 ) , .B2( u2_u5_u4_n170 ) , .A1( u2_u5_u4_n171 ) );
  INV_X1 u2_u5_u4_U31 (.A( u2_u5_u4_n158 ) , .ZN( u2_u5_u4_n182 ) );
  INV_X1 u2_u5_u4_U32 (.ZN( u2_u5_u4_n181 ) , .A( u2_u5_u4_n96 ) );
  INV_X1 u2_u5_u4_U33 (.A( u2_u5_u4_n144 ) , .ZN( u2_u5_u4_n179 ) );
  INV_X1 u2_u5_u4_U34 (.A( u2_u5_u4_n157 ) , .ZN( u2_u5_u4_n178 ) );
  NAND2_X1 u2_u5_u4_U35 (.A2( u2_u5_u4_n154 ) , .A1( u2_u5_u4_n96 ) , .ZN( u2_u5_u4_n97 ) );
  INV_X1 u2_u5_u4_U36 (.ZN( u2_u5_u4_n186 ) , .A( u2_u5_u4_n95 ) );
  OAI221_X1 u2_u5_u4_U37 (.C1( u2_u5_u4_n134 ) , .B1( u2_u5_u4_n158 ) , .B2( u2_u5_u4_n171 ) , .C2( u2_u5_u4_n173 ) , .A( u2_u5_u4_n94 ) , .ZN( u2_u5_u4_n95 ) );
  AOI222_X1 u2_u5_u4_U38 (.B2( u2_u5_u4_n132 ) , .A1( u2_u5_u4_n138 ) , .C2( u2_u5_u4_n175 ) , .A2( u2_u5_u4_n179 ) , .C1( u2_u5_u4_n181 ) , .B1( u2_u5_u4_n185 ) , .ZN( u2_u5_u4_n94 ) );
  INV_X1 u2_u5_u4_U39 (.A( u2_u5_u4_n113 ) , .ZN( u2_u5_u4_n185 ) );
  INV_X1 u2_u5_u4_U4 (.A( u2_u5_u4_n117 ) , .ZN( u2_u5_u4_n184 ) );
  INV_X1 u2_u5_u4_U40 (.A( u2_u5_u4_n143 ) , .ZN( u2_u5_u4_n183 ) );
  NOR2_X1 u2_u5_u4_U41 (.ZN( u2_u5_u4_n138 ) , .A1( u2_u5_u4_n168 ) , .A2( u2_u5_u4_n169 ) );
  NOR2_X1 u2_u5_u4_U42 (.A1( u2_u5_u4_n150 ) , .A2( u2_u5_u4_n152 ) , .ZN( u2_u5_u4_n153 ) );
  NOR2_X1 u2_u5_u4_U43 (.A2( u2_u5_u4_n128 ) , .A1( u2_u5_u4_n138 ) , .ZN( u2_u5_u4_n156 ) );
  AOI22_X1 u2_u5_u4_U44 (.B2( u2_u5_u4_n122 ) , .A1( u2_u5_u4_n123 ) , .ZN( u2_u5_u4_n124 ) , .B1( u2_u5_u4_n128 ) , .A2( u2_u5_u4_n172 ) );
  INV_X1 u2_u5_u4_U45 (.A( u2_u5_u4_n153 ) , .ZN( u2_u5_u4_n172 ) );
  NAND2_X1 u2_u5_u4_U46 (.A2( u2_u5_u4_n120 ) , .ZN( u2_u5_u4_n123 ) , .A1( u2_u5_u4_n161 ) );
  AOI22_X1 u2_u5_u4_U47 (.B2( u2_u5_u4_n132 ) , .A2( u2_u5_u4_n133 ) , .ZN( u2_u5_u4_n140 ) , .A1( u2_u5_u4_n150 ) , .B1( u2_u5_u4_n179 ) );
  NAND2_X1 u2_u5_u4_U48 (.ZN( u2_u5_u4_n133 ) , .A2( u2_u5_u4_n146 ) , .A1( u2_u5_u4_n154 ) );
  NAND2_X1 u2_u5_u4_U49 (.A1( u2_u5_u4_n103 ) , .ZN( u2_u5_u4_n154 ) , .A2( u2_u5_u4_n98 ) );
  NOR4_X1 u2_u5_u4_U5 (.A4( u2_u5_u4_n106 ) , .A3( u2_u5_u4_n107 ) , .A2( u2_u5_u4_n108 ) , .A1( u2_u5_u4_n109 ) , .ZN( u2_u5_u4_n110 ) );
  NAND2_X1 u2_u5_u4_U50 (.A1( u2_u5_u4_n101 ) , .ZN( u2_u5_u4_n158 ) , .A2( u2_u5_u4_n99 ) );
  AOI21_X1 u2_u5_u4_U51 (.ZN( u2_u5_u4_n127 ) , .A( u2_u5_u4_n136 ) , .B2( u2_u5_u4_n150 ) , .B1( u2_u5_u4_n180 ) );
  INV_X1 u2_u5_u4_U52 (.A( u2_u5_u4_n160 ) , .ZN( u2_u5_u4_n180 ) );
  NAND2_X1 u2_u5_u4_U53 (.A2( u2_u5_u4_n104 ) , .A1( u2_u5_u4_n105 ) , .ZN( u2_u5_u4_n146 ) );
  NAND2_X1 u2_u5_u4_U54 (.A2( u2_u5_u4_n101 ) , .A1( u2_u5_u4_n102 ) , .ZN( u2_u5_u4_n160 ) );
  NAND2_X1 u2_u5_u4_U55 (.ZN( u2_u5_u4_n134 ) , .A1( u2_u5_u4_n98 ) , .A2( u2_u5_u4_n99 ) );
  NAND2_X1 u2_u5_u4_U56 (.A1( u2_u5_u4_n103 ) , .A2( u2_u5_u4_n104 ) , .ZN( u2_u5_u4_n143 ) );
  NAND2_X1 u2_u5_u4_U57 (.A2( u2_u5_u4_n105 ) , .ZN( u2_u5_u4_n145 ) , .A1( u2_u5_u4_n98 ) );
  NAND2_X1 u2_u5_u4_U58 (.A1( u2_u5_u4_n100 ) , .A2( u2_u5_u4_n105 ) , .ZN( u2_u5_u4_n120 ) );
  NAND2_X1 u2_u5_u4_U59 (.A1( u2_u5_u4_n102 ) , .A2( u2_u5_u4_n104 ) , .ZN( u2_u5_u4_n148 ) );
  AOI21_X1 u2_u5_u4_U6 (.ZN( u2_u5_u4_n106 ) , .B2( u2_u5_u4_n146 ) , .B1( u2_u5_u4_n158 ) , .A( u2_u5_u4_n170 ) );
  NAND2_X1 u2_u5_u4_U60 (.A2( u2_u5_u4_n100 ) , .A1( u2_u5_u4_n103 ) , .ZN( u2_u5_u4_n157 ) );
  INV_X1 u2_u5_u4_U61 (.A( u2_u5_u4_n150 ) , .ZN( u2_u5_u4_n173 ) );
  INV_X1 u2_u5_u4_U62 (.A( u2_u5_u4_n152 ) , .ZN( u2_u5_u4_n171 ) );
  NAND2_X1 u2_u5_u4_U63 (.A1( u2_u5_u4_n100 ) , .ZN( u2_u5_u4_n118 ) , .A2( u2_u5_u4_n99 ) );
  NAND2_X1 u2_u5_u4_U64 (.A2( u2_u5_u4_n100 ) , .A1( u2_u5_u4_n102 ) , .ZN( u2_u5_u4_n144 ) );
  NAND2_X1 u2_u5_u4_U65 (.A2( u2_u5_u4_n101 ) , .A1( u2_u5_u4_n105 ) , .ZN( u2_u5_u4_n96 ) );
  INV_X1 u2_u5_u4_U66 (.A( u2_u5_u4_n128 ) , .ZN( u2_u5_u4_n174 ) );
  NAND2_X1 u2_u5_u4_U67 (.A2( u2_u5_u4_n102 ) , .ZN( u2_u5_u4_n119 ) , .A1( u2_u5_u4_n98 ) );
  NAND2_X1 u2_u5_u4_U68 (.A2( u2_u5_u4_n101 ) , .A1( u2_u5_u4_n103 ) , .ZN( u2_u5_u4_n147 ) );
  NAND2_X1 u2_u5_u4_U69 (.A2( u2_u5_u4_n104 ) , .ZN( u2_u5_u4_n113 ) , .A1( u2_u5_u4_n99 ) );
  AOI21_X1 u2_u5_u4_U7 (.ZN( u2_u5_u4_n108 ) , .B2( u2_u5_u4_n134 ) , .B1( u2_u5_u4_n155 ) , .A( u2_u5_u4_n156 ) );
  NOR2_X1 u2_u5_u4_U70 (.A2( u2_u5_X_28 ) , .ZN( u2_u5_u4_n150 ) , .A1( u2_u5_u4_n168 ) );
  NOR2_X1 u2_u5_u4_U71 (.A2( u2_u5_X_29 ) , .ZN( u2_u5_u4_n152 ) , .A1( u2_u5_u4_n169 ) );
  NOR2_X1 u2_u5_u4_U72 (.A2( u2_u5_X_30 ) , .ZN( u2_u5_u4_n105 ) , .A1( u2_u5_u4_n176 ) );
  NOR2_X1 u2_u5_u4_U73 (.A2( u2_u5_X_26 ) , .ZN( u2_u5_u4_n100 ) , .A1( u2_u5_u4_n177 ) );
  NOR2_X1 u2_u5_u4_U74 (.A2( u2_u5_X_28 ) , .A1( u2_u5_X_29 ) , .ZN( u2_u5_u4_n128 ) );
  NOR2_X1 u2_u5_u4_U75 (.A2( u2_u5_X_27 ) , .A1( u2_u5_X_30 ) , .ZN( u2_u5_u4_n102 ) );
  NOR2_X1 u2_u5_u4_U76 (.A2( u2_u5_X_25 ) , .A1( u2_u5_X_26 ) , .ZN( u2_u5_u4_n98 ) );
  AND2_X1 u2_u5_u4_U77 (.A2( u2_u5_X_25 ) , .A1( u2_u5_X_26 ) , .ZN( u2_u5_u4_n104 ) );
  AND2_X1 u2_u5_u4_U78 (.A1( u2_u5_X_30 ) , .A2( u2_u5_u4_n176 ) , .ZN( u2_u5_u4_n99 ) );
  AND2_X1 u2_u5_u4_U79 (.A1( u2_u5_X_26 ) , .ZN( u2_u5_u4_n101 ) , .A2( u2_u5_u4_n177 ) );
  AOI21_X1 u2_u5_u4_U8 (.ZN( u2_u5_u4_n109 ) , .A( u2_u5_u4_n153 ) , .B1( u2_u5_u4_n159 ) , .B2( u2_u5_u4_n184 ) );
  AND2_X1 u2_u5_u4_U80 (.A1( u2_u5_X_27 ) , .A2( u2_u5_X_30 ) , .ZN( u2_u5_u4_n103 ) );
  INV_X1 u2_u5_u4_U81 (.A( u2_u5_X_28 ) , .ZN( u2_u5_u4_n169 ) );
  INV_X1 u2_u5_u4_U82 (.A( u2_u5_X_29 ) , .ZN( u2_u5_u4_n168 ) );
  INV_X1 u2_u5_u4_U83 (.A( u2_u5_X_25 ) , .ZN( u2_u5_u4_n177 ) );
  INV_X1 u2_u5_u4_U84 (.A( u2_u5_X_27 ) , .ZN( u2_u5_u4_n176 ) );
  NAND4_X1 u2_u5_u4_U85 (.ZN( u2_out5_25 ) , .A4( u2_u5_u4_n139 ) , .A3( u2_u5_u4_n140 ) , .A2( u2_u5_u4_n141 ) , .A1( u2_u5_u4_n142 ) );
  OAI21_X1 u2_u5_u4_U86 (.A( u2_u5_u4_n128 ) , .B2( u2_u5_u4_n129 ) , .B1( u2_u5_u4_n130 ) , .ZN( u2_u5_u4_n142 ) );
  OAI21_X1 u2_u5_u4_U87 (.B2( u2_u5_u4_n131 ) , .ZN( u2_u5_u4_n141 ) , .A( u2_u5_u4_n175 ) , .B1( u2_u5_u4_n183 ) );
  NAND4_X1 u2_u5_u4_U88 (.ZN( u2_out5_14 ) , .A4( u2_u5_u4_n124 ) , .A3( u2_u5_u4_n125 ) , .A2( u2_u5_u4_n126 ) , .A1( u2_u5_u4_n127 ) );
  AOI22_X1 u2_u5_u4_U89 (.B2( u2_u5_u4_n117 ) , .ZN( u2_u5_u4_n126 ) , .A1( u2_u5_u4_n129 ) , .B1( u2_u5_u4_n152 ) , .A2( u2_u5_u4_n175 ) );
  AOI211_X1 u2_u5_u4_U9 (.B( u2_u5_u4_n136 ) , .A( u2_u5_u4_n137 ) , .C2( u2_u5_u4_n138 ) , .ZN( u2_u5_u4_n139 ) , .C1( u2_u5_u4_n182 ) );
  AOI22_X1 u2_u5_u4_U90 (.ZN( u2_u5_u4_n125 ) , .B2( u2_u5_u4_n131 ) , .A2( u2_u5_u4_n132 ) , .B1( u2_u5_u4_n138 ) , .A1( u2_u5_u4_n178 ) );
  NAND4_X1 u2_u5_u4_U91 (.ZN( u2_out5_8 ) , .A4( u2_u5_u4_n110 ) , .A3( u2_u5_u4_n111 ) , .A2( u2_u5_u4_n112 ) , .A1( u2_u5_u4_n186 ) );
  NAND2_X1 u2_u5_u4_U92 (.ZN( u2_u5_u4_n112 ) , .A2( u2_u5_u4_n130 ) , .A1( u2_u5_u4_n150 ) );
  AOI22_X1 u2_u5_u4_U93 (.ZN( u2_u5_u4_n111 ) , .B2( u2_u5_u4_n132 ) , .A1( u2_u5_u4_n152 ) , .B1( u2_u5_u4_n178 ) , .A2( u2_u5_u4_n97 ) );
  AOI22_X1 u2_u5_u4_U94 (.B2( u2_u5_u4_n149 ) , .B1( u2_u5_u4_n150 ) , .A2( u2_u5_u4_n151 ) , .A1( u2_u5_u4_n152 ) , .ZN( u2_u5_u4_n167 ) );
  NOR4_X1 u2_u5_u4_U95 (.A4( u2_u5_u4_n162 ) , .A3( u2_u5_u4_n163 ) , .A2( u2_u5_u4_n164 ) , .A1( u2_u5_u4_n165 ) , .ZN( u2_u5_u4_n166 ) );
  NAND3_X1 u2_u5_u4_U96 (.ZN( u2_out5_3 ) , .A3( u2_u5_u4_n166 ) , .A1( u2_u5_u4_n167 ) , .A2( u2_u5_u4_n186 ) );
  NAND3_X1 u2_u5_u4_U97 (.A3( u2_u5_u4_n146 ) , .A2( u2_u5_u4_n147 ) , .A1( u2_u5_u4_n148 ) , .ZN( u2_u5_u4_n149 ) );
  NAND3_X1 u2_u5_u4_U98 (.A3( u2_u5_u4_n143 ) , .A2( u2_u5_u4_n144 ) , .A1( u2_u5_u4_n145 ) , .ZN( u2_u5_u4_n151 ) );
  NAND3_X1 u2_u5_u4_U99 (.A3( u2_u5_u4_n121 ) , .ZN( u2_u5_u4_n122 ) , .A2( u2_u5_u4_n144 ) , .A1( u2_u5_u4_n154 ) );
  XOR2_X1 u2_u7_U13 (.B( u2_K8_42 ) , .A( u2_R6_29 ) , .Z( u2_u7_X_42 ) );
  XOR2_X1 u2_u7_U14 (.B( u2_K8_41 ) , .A( u2_R6_28 ) , .Z( u2_u7_X_41 ) );
  XOR2_X1 u2_u7_U15 (.B( u2_K8_40 ) , .A( u2_R6_27 ) , .Z( u2_u7_X_40 ) );
  XOR2_X1 u2_u7_U17 (.B( u2_K8_39 ) , .A( u2_R6_26 ) , .Z( u2_u7_X_39 ) );
  XOR2_X1 u2_u7_U18 (.B( u2_K8_38 ) , .A( u2_R6_25 ) , .Z( u2_u7_X_38 ) );
  XOR2_X1 u2_u7_U19 (.B( u2_K8_37 ) , .A( u2_R6_24 ) , .Z( u2_u7_X_37 ) );
  XOR2_X1 u2_u7_U20 (.B( u2_K8_36 ) , .A( u2_R6_25 ) , .Z( u2_u7_X_36 ) );
  XOR2_X1 u2_u7_U21 (.B( u2_K8_35 ) , .A( u2_R6_24 ) , .Z( u2_u7_X_35 ) );
  XOR2_X1 u2_u7_U22 (.B( u2_K8_34 ) , .A( u2_R6_23 ) , .Z( u2_u7_X_34 ) );
  XOR2_X1 u2_u7_U23 (.B( u2_K8_33 ) , .A( u2_R6_22 ) , .Z( u2_u7_X_33 ) );
  XOR2_X1 u2_u7_U24 (.B( u2_K8_32 ) , .A( u2_R6_21 ) , .Z( u2_u7_X_32 ) );
  XOR2_X1 u2_u7_U25 (.B( u2_K8_31 ) , .A( u2_R6_20 ) , .Z( u2_u7_X_31 ) );
  XOR2_X1 u2_u7_U26 (.B( u2_K8_30 ) , .A( u2_R6_21 ) , .Z( u2_u7_X_30 ) );
  XOR2_X1 u2_u7_U28 (.B( u2_K8_29 ) , .A( u2_R6_20 ) , .Z( u2_u7_X_29 ) );
  XOR2_X1 u2_u7_U29 (.B( u2_K8_28 ) , .A( u2_R6_19 ) , .Z( u2_u7_X_28 ) );
  XOR2_X1 u2_u7_U30 (.B( u2_K8_27 ) , .A( u2_R6_18 ) , .Z( u2_u7_X_27 ) );
  XOR2_X1 u2_u7_U31 (.B( u2_K8_26 ) , .A( u2_R6_17 ) , .Z( u2_u7_X_26 ) );
  XOR2_X1 u2_u7_U32 (.B( u2_K8_25 ) , .A( u2_R6_16 ) , .Z( u2_u7_X_25 ) );
  XOR2_X1 u2_u7_U33 (.B( u2_K8_24 ) , .A( u2_R6_17 ) , .Z( u2_u7_X_24 ) );
  XOR2_X1 u2_u7_U34 (.B( u2_K8_23 ) , .A( u2_R6_16 ) , .Z( u2_u7_X_23 ) );
  XOR2_X1 u2_u7_U35 (.B( u2_K8_22 ) , .A( u2_R6_15 ) , .Z( u2_u7_X_22 ) );
  XOR2_X1 u2_u7_U36 (.B( u2_K8_21 ) , .A( u2_R6_14 ) , .Z( u2_u7_X_21 ) );
  XOR2_X1 u2_u7_U37 (.B( u2_K8_20 ) , .A( u2_R6_13 ) , .Z( u2_u7_X_20 ) );
  XOR2_X1 u2_u7_U39 (.B( u2_K8_19 ) , .A( u2_R6_12 ) , .Z( u2_u7_X_19 ) );
  OAI22_X1 u2_u7_u3_U10 (.B1( u2_u7_u3_n113 ) , .A2( u2_u7_u3_n135 ) , .A1( u2_u7_u3_n150 ) , .B2( u2_u7_u3_n164 ) , .ZN( u2_u7_u3_n98 ) );
  OAI211_X1 u2_u7_u3_U11 (.B( u2_u7_u3_n106 ) , .ZN( u2_u7_u3_n119 ) , .C2( u2_u7_u3_n128 ) , .C1( u2_u7_u3_n167 ) , .A( u2_u7_u3_n181 ) );
  AOI221_X1 u2_u7_u3_U12 (.C1( u2_u7_u3_n105 ) , .ZN( u2_u7_u3_n106 ) , .A( u2_u7_u3_n131 ) , .B2( u2_u7_u3_n132 ) , .C2( u2_u7_u3_n133 ) , .B1( u2_u7_u3_n169 ) );
  INV_X1 u2_u7_u3_U13 (.ZN( u2_u7_u3_n181 ) , .A( u2_u7_u3_n98 ) );
  NAND2_X1 u2_u7_u3_U14 (.ZN( u2_u7_u3_n105 ) , .A2( u2_u7_u3_n130 ) , .A1( u2_u7_u3_n155 ) );
  AOI22_X1 u2_u7_u3_U15 (.B1( u2_u7_u3_n115 ) , .A2( u2_u7_u3_n116 ) , .ZN( u2_u7_u3_n123 ) , .B2( u2_u7_u3_n133 ) , .A1( u2_u7_u3_n169 ) );
  NAND2_X1 u2_u7_u3_U16 (.ZN( u2_u7_u3_n116 ) , .A2( u2_u7_u3_n151 ) , .A1( u2_u7_u3_n182 ) );
  NOR2_X1 u2_u7_u3_U17 (.ZN( u2_u7_u3_n126 ) , .A2( u2_u7_u3_n150 ) , .A1( u2_u7_u3_n164 ) );
  AOI21_X1 u2_u7_u3_U18 (.ZN( u2_u7_u3_n112 ) , .B2( u2_u7_u3_n146 ) , .B1( u2_u7_u3_n155 ) , .A( u2_u7_u3_n167 ) );
  NAND2_X1 u2_u7_u3_U19 (.A1( u2_u7_u3_n135 ) , .ZN( u2_u7_u3_n142 ) , .A2( u2_u7_u3_n164 ) );
  NAND2_X1 u2_u7_u3_U20 (.ZN( u2_u7_u3_n132 ) , .A2( u2_u7_u3_n152 ) , .A1( u2_u7_u3_n156 ) );
  AND2_X1 u2_u7_u3_U21 (.A2( u2_u7_u3_n113 ) , .A1( u2_u7_u3_n114 ) , .ZN( u2_u7_u3_n151 ) );
  INV_X1 u2_u7_u3_U22 (.A( u2_u7_u3_n133 ) , .ZN( u2_u7_u3_n165 ) );
  INV_X1 u2_u7_u3_U23 (.A( u2_u7_u3_n135 ) , .ZN( u2_u7_u3_n170 ) );
  NAND2_X1 u2_u7_u3_U24 (.A1( u2_u7_u3_n107 ) , .A2( u2_u7_u3_n108 ) , .ZN( u2_u7_u3_n140 ) );
  NAND2_X1 u2_u7_u3_U25 (.ZN( u2_u7_u3_n117 ) , .A1( u2_u7_u3_n124 ) , .A2( u2_u7_u3_n148 ) );
  NAND2_X1 u2_u7_u3_U26 (.ZN( u2_u7_u3_n143 ) , .A1( u2_u7_u3_n165 ) , .A2( u2_u7_u3_n167 ) );
  INV_X1 u2_u7_u3_U27 (.A( u2_u7_u3_n130 ) , .ZN( u2_u7_u3_n177 ) );
  INV_X1 u2_u7_u3_U28 (.A( u2_u7_u3_n128 ) , .ZN( u2_u7_u3_n176 ) );
  INV_X1 u2_u7_u3_U29 (.A( u2_u7_u3_n155 ) , .ZN( u2_u7_u3_n174 ) );
  INV_X1 u2_u7_u3_U3 (.A( u2_u7_u3_n129 ) , .ZN( u2_u7_u3_n183 ) );
  INV_X1 u2_u7_u3_U30 (.A( u2_u7_u3_n139 ) , .ZN( u2_u7_u3_n185 ) );
  NOR2_X1 u2_u7_u3_U31 (.ZN( u2_u7_u3_n135 ) , .A2( u2_u7_u3_n141 ) , .A1( u2_u7_u3_n169 ) );
  OAI222_X1 u2_u7_u3_U32 (.C2( u2_u7_u3_n107 ) , .A2( u2_u7_u3_n108 ) , .B1( u2_u7_u3_n135 ) , .ZN( u2_u7_u3_n138 ) , .B2( u2_u7_u3_n146 ) , .C1( u2_u7_u3_n154 ) , .A1( u2_u7_u3_n164 ) );
  NOR4_X1 u2_u7_u3_U33 (.A4( u2_u7_u3_n157 ) , .A3( u2_u7_u3_n158 ) , .A2( u2_u7_u3_n159 ) , .A1( u2_u7_u3_n160 ) , .ZN( u2_u7_u3_n161 ) );
  AOI21_X1 u2_u7_u3_U34 (.B2( u2_u7_u3_n152 ) , .B1( u2_u7_u3_n153 ) , .ZN( u2_u7_u3_n158 ) , .A( u2_u7_u3_n164 ) );
  AOI21_X1 u2_u7_u3_U35 (.A( u2_u7_u3_n154 ) , .B2( u2_u7_u3_n155 ) , .B1( u2_u7_u3_n156 ) , .ZN( u2_u7_u3_n157 ) );
  AOI21_X1 u2_u7_u3_U36 (.A( u2_u7_u3_n149 ) , .B2( u2_u7_u3_n150 ) , .B1( u2_u7_u3_n151 ) , .ZN( u2_u7_u3_n159 ) );
  AOI211_X1 u2_u7_u3_U37 (.ZN( u2_u7_u3_n109 ) , .A( u2_u7_u3_n119 ) , .C2( u2_u7_u3_n129 ) , .B( u2_u7_u3_n138 ) , .C1( u2_u7_u3_n141 ) );
  AOI211_X1 u2_u7_u3_U38 (.B( u2_u7_u3_n119 ) , .A( u2_u7_u3_n120 ) , .C2( u2_u7_u3_n121 ) , .ZN( u2_u7_u3_n122 ) , .C1( u2_u7_u3_n179 ) );
  INV_X1 u2_u7_u3_U39 (.A( u2_u7_u3_n156 ) , .ZN( u2_u7_u3_n179 ) );
  INV_X1 u2_u7_u3_U4 (.A( u2_u7_u3_n140 ) , .ZN( u2_u7_u3_n182 ) );
  OAI22_X1 u2_u7_u3_U40 (.B1( u2_u7_u3_n118 ) , .ZN( u2_u7_u3_n120 ) , .A1( u2_u7_u3_n135 ) , .B2( u2_u7_u3_n154 ) , .A2( u2_u7_u3_n178 ) );
  AND3_X1 u2_u7_u3_U41 (.ZN( u2_u7_u3_n118 ) , .A2( u2_u7_u3_n124 ) , .A1( u2_u7_u3_n144 ) , .A3( u2_u7_u3_n152 ) );
  INV_X1 u2_u7_u3_U42 (.A( u2_u7_u3_n121 ) , .ZN( u2_u7_u3_n164 ) );
  NAND2_X1 u2_u7_u3_U43 (.ZN( u2_u7_u3_n133 ) , .A1( u2_u7_u3_n154 ) , .A2( u2_u7_u3_n164 ) );
  OAI211_X1 u2_u7_u3_U44 (.B( u2_u7_u3_n127 ) , .ZN( u2_u7_u3_n139 ) , .C1( u2_u7_u3_n150 ) , .C2( u2_u7_u3_n154 ) , .A( u2_u7_u3_n184 ) );
  INV_X1 u2_u7_u3_U45 (.A( u2_u7_u3_n125 ) , .ZN( u2_u7_u3_n184 ) );
  AOI221_X1 u2_u7_u3_U46 (.A( u2_u7_u3_n126 ) , .ZN( u2_u7_u3_n127 ) , .C2( u2_u7_u3_n132 ) , .C1( u2_u7_u3_n169 ) , .B2( u2_u7_u3_n170 ) , .B1( u2_u7_u3_n174 ) );
  OAI22_X1 u2_u7_u3_U47 (.A1( u2_u7_u3_n124 ) , .ZN( u2_u7_u3_n125 ) , .B2( u2_u7_u3_n145 ) , .A2( u2_u7_u3_n165 ) , .B1( u2_u7_u3_n167 ) );
  NOR2_X1 u2_u7_u3_U48 (.A1( u2_u7_u3_n113 ) , .ZN( u2_u7_u3_n131 ) , .A2( u2_u7_u3_n154 ) );
  NAND2_X1 u2_u7_u3_U49 (.A1( u2_u7_u3_n103 ) , .ZN( u2_u7_u3_n150 ) , .A2( u2_u7_u3_n99 ) );
  INV_X1 u2_u7_u3_U5 (.A( u2_u7_u3_n117 ) , .ZN( u2_u7_u3_n178 ) );
  NAND2_X1 u2_u7_u3_U50 (.A2( u2_u7_u3_n102 ) , .ZN( u2_u7_u3_n155 ) , .A1( u2_u7_u3_n97 ) );
  INV_X1 u2_u7_u3_U51 (.A( u2_u7_u3_n141 ) , .ZN( u2_u7_u3_n167 ) );
  AOI21_X1 u2_u7_u3_U52 (.B2( u2_u7_u3_n114 ) , .B1( u2_u7_u3_n146 ) , .A( u2_u7_u3_n154 ) , .ZN( u2_u7_u3_n94 ) );
  AOI21_X1 u2_u7_u3_U53 (.ZN( u2_u7_u3_n110 ) , .B2( u2_u7_u3_n142 ) , .B1( u2_u7_u3_n186 ) , .A( u2_u7_u3_n95 ) );
  INV_X1 u2_u7_u3_U54 (.A( u2_u7_u3_n145 ) , .ZN( u2_u7_u3_n186 ) );
  AOI21_X1 u2_u7_u3_U55 (.B1( u2_u7_u3_n124 ) , .A( u2_u7_u3_n149 ) , .B2( u2_u7_u3_n155 ) , .ZN( u2_u7_u3_n95 ) );
  INV_X1 u2_u7_u3_U56 (.A( u2_u7_u3_n149 ) , .ZN( u2_u7_u3_n169 ) );
  NAND2_X1 u2_u7_u3_U57 (.ZN( u2_u7_u3_n124 ) , .A1( u2_u7_u3_n96 ) , .A2( u2_u7_u3_n97 ) );
  NAND2_X1 u2_u7_u3_U58 (.A2( u2_u7_u3_n100 ) , .ZN( u2_u7_u3_n146 ) , .A1( u2_u7_u3_n96 ) );
  NAND2_X1 u2_u7_u3_U59 (.A1( u2_u7_u3_n101 ) , .ZN( u2_u7_u3_n145 ) , .A2( u2_u7_u3_n99 ) );
  AOI221_X1 u2_u7_u3_U6 (.A( u2_u7_u3_n131 ) , .C2( u2_u7_u3_n132 ) , .C1( u2_u7_u3_n133 ) , .ZN( u2_u7_u3_n134 ) , .B1( u2_u7_u3_n143 ) , .B2( u2_u7_u3_n177 ) );
  NAND2_X1 u2_u7_u3_U60 (.A1( u2_u7_u3_n100 ) , .ZN( u2_u7_u3_n156 ) , .A2( u2_u7_u3_n99 ) );
  NAND2_X1 u2_u7_u3_U61 (.A2( u2_u7_u3_n101 ) , .A1( u2_u7_u3_n104 ) , .ZN( u2_u7_u3_n148 ) );
  NAND2_X1 u2_u7_u3_U62 (.A1( u2_u7_u3_n100 ) , .A2( u2_u7_u3_n102 ) , .ZN( u2_u7_u3_n128 ) );
  NAND2_X1 u2_u7_u3_U63 (.A2( u2_u7_u3_n101 ) , .A1( u2_u7_u3_n102 ) , .ZN( u2_u7_u3_n152 ) );
  NAND2_X1 u2_u7_u3_U64 (.A2( u2_u7_u3_n101 ) , .ZN( u2_u7_u3_n114 ) , .A1( u2_u7_u3_n96 ) );
  NAND2_X1 u2_u7_u3_U65 (.ZN( u2_u7_u3_n107 ) , .A1( u2_u7_u3_n97 ) , .A2( u2_u7_u3_n99 ) );
  NAND2_X1 u2_u7_u3_U66 (.A2( u2_u7_u3_n100 ) , .A1( u2_u7_u3_n104 ) , .ZN( u2_u7_u3_n113 ) );
  NAND2_X1 u2_u7_u3_U67 (.A1( u2_u7_u3_n104 ) , .ZN( u2_u7_u3_n153 ) , .A2( u2_u7_u3_n97 ) );
  NAND2_X1 u2_u7_u3_U68 (.A2( u2_u7_u3_n103 ) , .A1( u2_u7_u3_n104 ) , .ZN( u2_u7_u3_n130 ) );
  NAND2_X1 u2_u7_u3_U69 (.A2( u2_u7_u3_n103 ) , .ZN( u2_u7_u3_n144 ) , .A1( u2_u7_u3_n96 ) );
  OAI22_X1 u2_u7_u3_U7 (.B2( u2_u7_u3_n147 ) , .A2( u2_u7_u3_n148 ) , .ZN( u2_u7_u3_n160 ) , .B1( u2_u7_u3_n165 ) , .A1( u2_u7_u3_n168 ) );
  NAND2_X1 u2_u7_u3_U70 (.A1( u2_u7_u3_n102 ) , .A2( u2_u7_u3_n103 ) , .ZN( u2_u7_u3_n108 ) );
  NOR2_X1 u2_u7_u3_U71 (.A2( u2_u7_X_19 ) , .A1( u2_u7_X_20 ) , .ZN( u2_u7_u3_n99 ) );
  NOR2_X1 u2_u7_u3_U72 (.A2( u2_u7_X_21 ) , .A1( u2_u7_X_24 ) , .ZN( u2_u7_u3_n103 ) );
  NOR2_X1 u2_u7_u3_U73 (.A2( u2_u7_X_24 ) , .A1( u2_u7_u3_n171 ) , .ZN( u2_u7_u3_n97 ) );
  NOR2_X1 u2_u7_u3_U74 (.A2( u2_u7_X_23 ) , .ZN( u2_u7_u3_n141 ) , .A1( u2_u7_u3_n166 ) );
  NOR2_X1 u2_u7_u3_U75 (.A2( u2_u7_X_19 ) , .A1( u2_u7_u3_n172 ) , .ZN( u2_u7_u3_n96 ) );
  NAND2_X1 u2_u7_u3_U76 (.A1( u2_u7_X_22 ) , .A2( u2_u7_X_23 ) , .ZN( u2_u7_u3_n154 ) );
  NAND2_X1 u2_u7_u3_U77 (.A1( u2_u7_X_23 ) , .ZN( u2_u7_u3_n149 ) , .A2( u2_u7_u3_n166 ) );
  NOR2_X1 u2_u7_u3_U78 (.A2( u2_u7_X_22 ) , .A1( u2_u7_X_23 ) , .ZN( u2_u7_u3_n121 ) );
  AND2_X1 u2_u7_u3_U79 (.A1( u2_u7_X_24 ) , .ZN( u2_u7_u3_n101 ) , .A2( u2_u7_u3_n171 ) );
  AND3_X1 u2_u7_u3_U8 (.A3( u2_u7_u3_n144 ) , .A2( u2_u7_u3_n145 ) , .A1( u2_u7_u3_n146 ) , .ZN( u2_u7_u3_n147 ) );
  AND2_X1 u2_u7_u3_U80 (.A1( u2_u7_X_19 ) , .ZN( u2_u7_u3_n102 ) , .A2( u2_u7_u3_n172 ) );
  AND2_X1 u2_u7_u3_U81 (.A1( u2_u7_X_21 ) , .A2( u2_u7_X_24 ) , .ZN( u2_u7_u3_n100 ) );
  AND2_X1 u2_u7_u3_U82 (.A2( u2_u7_X_19 ) , .A1( u2_u7_X_20 ) , .ZN( u2_u7_u3_n104 ) );
  INV_X1 u2_u7_u3_U83 (.A( u2_u7_X_22 ) , .ZN( u2_u7_u3_n166 ) );
  INV_X1 u2_u7_u3_U84 (.A( u2_u7_X_21 ) , .ZN( u2_u7_u3_n171 ) );
  INV_X1 u2_u7_u3_U85 (.A( u2_u7_X_20 ) , .ZN( u2_u7_u3_n172 ) );
  OR4_X1 u2_u7_u3_U86 (.ZN( u2_out7_10 ) , .A4( u2_u7_u3_n136 ) , .A3( u2_u7_u3_n137 ) , .A1( u2_u7_u3_n138 ) , .A2( u2_u7_u3_n139 ) );
  OAI222_X1 u2_u7_u3_U87 (.C1( u2_u7_u3_n128 ) , .ZN( u2_u7_u3_n137 ) , .B1( u2_u7_u3_n148 ) , .A2( u2_u7_u3_n150 ) , .B2( u2_u7_u3_n154 ) , .C2( u2_u7_u3_n164 ) , .A1( u2_u7_u3_n167 ) );
  OAI221_X1 u2_u7_u3_U88 (.A( u2_u7_u3_n134 ) , .B2( u2_u7_u3_n135 ) , .ZN( u2_u7_u3_n136 ) , .C1( u2_u7_u3_n149 ) , .B1( u2_u7_u3_n151 ) , .C2( u2_u7_u3_n183 ) );
  NAND4_X1 u2_u7_u3_U89 (.ZN( u2_out7_26 ) , .A4( u2_u7_u3_n109 ) , .A3( u2_u7_u3_n110 ) , .A2( u2_u7_u3_n111 ) , .A1( u2_u7_u3_n173 ) );
  INV_X1 u2_u7_u3_U9 (.A( u2_u7_u3_n143 ) , .ZN( u2_u7_u3_n168 ) );
  INV_X1 u2_u7_u3_U90 (.ZN( u2_u7_u3_n173 ) , .A( u2_u7_u3_n94 ) );
  OAI21_X1 u2_u7_u3_U91 (.ZN( u2_u7_u3_n111 ) , .B2( u2_u7_u3_n117 ) , .A( u2_u7_u3_n133 ) , .B1( u2_u7_u3_n176 ) );
  NAND4_X1 u2_u7_u3_U92 (.ZN( u2_out7_20 ) , .A4( u2_u7_u3_n122 ) , .A3( u2_u7_u3_n123 ) , .A1( u2_u7_u3_n175 ) , .A2( u2_u7_u3_n180 ) );
  INV_X1 u2_u7_u3_U93 (.A( u2_u7_u3_n126 ) , .ZN( u2_u7_u3_n180 ) );
  INV_X1 u2_u7_u3_U94 (.A( u2_u7_u3_n112 ) , .ZN( u2_u7_u3_n175 ) );
  NAND4_X1 u2_u7_u3_U95 (.ZN( u2_out7_1 ) , .A4( u2_u7_u3_n161 ) , .A3( u2_u7_u3_n162 ) , .A2( u2_u7_u3_n163 ) , .A1( u2_u7_u3_n185 ) );
  NAND2_X1 u2_u7_u3_U96 (.ZN( u2_u7_u3_n163 ) , .A2( u2_u7_u3_n170 ) , .A1( u2_u7_u3_n176 ) );
  AOI22_X1 u2_u7_u3_U97 (.B2( u2_u7_u3_n140 ) , .B1( u2_u7_u3_n141 ) , .A2( u2_u7_u3_n142 ) , .ZN( u2_u7_u3_n162 ) , .A1( u2_u7_u3_n177 ) );
  NAND3_X1 u2_u7_u3_U98 (.A1( u2_u7_u3_n114 ) , .ZN( u2_u7_u3_n115 ) , .A2( u2_u7_u3_n145 ) , .A3( u2_u7_u3_n153 ) );
  NAND3_X1 u2_u7_u3_U99 (.ZN( u2_u7_u3_n129 ) , .A2( u2_u7_u3_n144 ) , .A1( u2_u7_u3_n153 ) , .A3( u2_u7_u3_n182 ) );
  OAI22_X1 u2_u7_u4_U10 (.B2( u2_u7_u4_n135 ) , .ZN( u2_u7_u4_n137 ) , .B1( u2_u7_u4_n153 ) , .A1( u2_u7_u4_n155 ) , .A2( u2_u7_u4_n171 ) );
  AND3_X1 u2_u7_u4_U11 (.A2( u2_u7_u4_n134 ) , .ZN( u2_u7_u4_n135 ) , .A3( u2_u7_u4_n145 ) , .A1( u2_u7_u4_n157 ) );
  OR3_X1 u2_u7_u4_U12 (.A3( u2_u7_u4_n114 ) , .A2( u2_u7_u4_n115 ) , .A1( u2_u7_u4_n116 ) , .ZN( u2_u7_u4_n136 ) );
  AOI21_X1 u2_u7_u4_U13 (.A( u2_u7_u4_n113 ) , .ZN( u2_u7_u4_n116 ) , .B2( u2_u7_u4_n173 ) , .B1( u2_u7_u4_n174 ) );
  AOI21_X1 u2_u7_u4_U14 (.ZN( u2_u7_u4_n115 ) , .B2( u2_u7_u4_n145 ) , .B1( u2_u7_u4_n146 ) , .A( u2_u7_u4_n156 ) );
  OAI22_X1 u2_u7_u4_U15 (.ZN( u2_u7_u4_n114 ) , .A2( u2_u7_u4_n121 ) , .B1( u2_u7_u4_n160 ) , .B2( u2_u7_u4_n170 ) , .A1( u2_u7_u4_n171 ) );
  NAND2_X1 u2_u7_u4_U16 (.ZN( u2_u7_u4_n132 ) , .A2( u2_u7_u4_n170 ) , .A1( u2_u7_u4_n173 ) );
  AOI21_X1 u2_u7_u4_U17 (.B2( u2_u7_u4_n160 ) , .B1( u2_u7_u4_n161 ) , .ZN( u2_u7_u4_n162 ) , .A( u2_u7_u4_n170 ) );
  AOI21_X1 u2_u7_u4_U18 (.ZN( u2_u7_u4_n107 ) , .B2( u2_u7_u4_n143 ) , .A( u2_u7_u4_n174 ) , .B1( u2_u7_u4_n184 ) );
  AOI21_X1 u2_u7_u4_U19 (.B2( u2_u7_u4_n158 ) , .B1( u2_u7_u4_n159 ) , .ZN( u2_u7_u4_n163 ) , .A( u2_u7_u4_n174 ) );
  AOI21_X1 u2_u7_u4_U20 (.A( u2_u7_u4_n153 ) , .B2( u2_u7_u4_n154 ) , .B1( u2_u7_u4_n155 ) , .ZN( u2_u7_u4_n165 ) );
  AOI21_X1 u2_u7_u4_U21 (.A( u2_u7_u4_n156 ) , .B2( u2_u7_u4_n157 ) , .ZN( u2_u7_u4_n164 ) , .B1( u2_u7_u4_n184 ) );
  INV_X1 u2_u7_u4_U22 (.A( u2_u7_u4_n138 ) , .ZN( u2_u7_u4_n170 ) );
  AND2_X1 u2_u7_u4_U23 (.A2( u2_u7_u4_n120 ) , .ZN( u2_u7_u4_n155 ) , .A1( u2_u7_u4_n160 ) );
  INV_X1 u2_u7_u4_U24 (.A( u2_u7_u4_n156 ) , .ZN( u2_u7_u4_n175 ) );
  NAND2_X1 u2_u7_u4_U25 (.A2( u2_u7_u4_n118 ) , .ZN( u2_u7_u4_n131 ) , .A1( u2_u7_u4_n147 ) );
  NAND2_X1 u2_u7_u4_U26 (.A1( u2_u7_u4_n119 ) , .A2( u2_u7_u4_n120 ) , .ZN( u2_u7_u4_n130 ) );
  NAND2_X1 u2_u7_u4_U27 (.ZN( u2_u7_u4_n117 ) , .A2( u2_u7_u4_n118 ) , .A1( u2_u7_u4_n148 ) );
  NAND2_X1 u2_u7_u4_U28 (.ZN( u2_u7_u4_n129 ) , .A1( u2_u7_u4_n134 ) , .A2( u2_u7_u4_n148 ) );
  AND3_X1 u2_u7_u4_U29 (.A1( u2_u7_u4_n119 ) , .A2( u2_u7_u4_n143 ) , .A3( u2_u7_u4_n154 ) , .ZN( u2_u7_u4_n161 ) );
  NOR2_X1 u2_u7_u4_U3 (.ZN( u2_u7_u4_n121 ) , .A1( u2_u7_u4_n181 ) , .A2( u2_u7_u4_n182 ) );
  AND2_X1 u2_u7_u4_U30 (.A1( u2_u7_u4_n145 ) , .A2( u2_u7_u4_n147 ) , .ZN( u2_u7_u4_n159 ) );
  INV_X1 u2_u7_u4_U31 (.A( u2_u7_u4_n158 ) , .ZN( u2_u7_u4_n182 ) );
  INV_X1 u2_u7_u4_U32 (.ZN( u2_u7_u4_n181 ) , .A( u2_u7_u4_n96 ) );
  INV_X1 u2_u7_u4_U33 (.A( u2_u7_u4_n144 ) , .ZN( u2_u7_u4_n179 ) );
  INV_X1 u2_u7_u4_U34 (.A( u2_u7_u4_n157 ) , .ZN( u2_u7_u4_n178 ) );
  NAND2_X1 u2_u7_u4_U35 (.A2( u2_u7_u4_n154 ) , .A1( u2_u7_u4_n96 ) , .ZN( u2_u7_u4_n97 ) );
  INV_X1 u2_u7_u4_U36 (.ZN( u2_u7_u4_n186 ) , .A( u2_u7_u4_n95 ) );
  OAI221_X1 u2_u7_u4_U37 (.C1( u2_u7_u4_n134 ) , .B1( u2_u7_u4_n158 ) , .B2( u2_u7_u4_n171 ) , .C2( u2_u7_u4_n173 ) , .A( u2_u7_u4_n94 ) , .ZN( u2_u7_u4_n95 ) );
  AOI222_X1 u2_u7_u4_U38 (.B2( u2_u7_u4_n132 ) , .A1( u2_u7_u4_n138 ) , .C2( u2_u7_u4_n175 ) , .A2( u2_u7_u4_n179 ) , .C1( u2_u7_u4_n181 ) , .B1( u2_u7_u4_n185 ) , .ZN( u2_u7_u4_n94 ) );
  INV_X1 u2_u7_u4_U39 (.A( u2_u7_u4_n113 ) , .ZN( u2_u7_u4_n185 ) );
  INV_X1 u2_u7_u4_U4 (.A( u2_u7_u4_n117 ) , .ZN( u2_u7_u4_n184 ) );
  INV_X1 u2_u7_u4_U40 (.A( u2_u7_u4_n143 ) , .ZN( u2_u7_u4_n183 ) );
  NOR2_X1 u2_u7_u4_U41 (.ZN( u2_u7_u4_n138 ) , .A1( u2_u7_u4_n168 ) , .A2( u2_u7_u4_n169 ) );
  NOR2_X1 u2_u7_u4_U42 (.A1( u2_u7_u4_n150 ) , .A2( u2_u7_u4_n152 ) , .ZN( u2_u7_u4_n153 ) );
  NOR2_X1 u2_u7_u4_U43 (.A2( u2_u7_u4_n128 ) , .A1( u2_u7_u4_n138 ) , .ZN( u2_u7_u4_n156 ) );
  AOI22_X1 u2_u7_u4_U44 (.B2( u2_u7_u4_n122 ) , .A1( u2_u7_u4_n123 ) , .ZN( u2_u7_u4_n124 ) , .B1( u2_u7_u4_n128 ) , .A2( u2_u7_u4_n172 ) );
  NAND2_X1 u2_u7_u4_U45 (.A2( u2_u7_u4_n120 ) , .ZN( u2_u7_u4_n123 ) , .A1( u2_u7_u4_n161 ) );
  INV_X1 u2_u7_u4_U46 (.A( u2_u7_u4_n153 ) , .ZN( u2_u7_u4_n172 ) );
  AOI22_X1 u2_u7_u4_U47 (.B2( u2_u7_u4_n132 ) , .A2( u2_u7_u4_n133 ) , .ZN( u2_u7_u4_n140 ) , .A1( u2_u7_u4_n150 ) , .B1( u2_u7_u4_n179 ) );
  NAND2_X1 u2_u7_u4_U48 (.ZN( u2_u7_u4_n133 ) , .A2( u2_u7_u4_n146 ) , .A1( u2_u7_u4_n154 ) );
  NAND2_X1 u2_u7_u4_U49 (.A1( u2_u7_u4_n103 ) , .ZN( u2_u7_u4_n154 ) , .A2( u2_u7_u4_n98 ) );
  NOR4_X1 u2_u7_u4_U5 (.A4( u2_u7_u4_n106 ) , .A3( u2_u7_u4_n107 ) , .A2( u2_u7_u4_n108 ) , .A1( u2_u7_u4_n109 ) , .ZN( u2_u7_u4_n110 ) );
  NAND2_X1 u2_u7_u4_U50 (.A1( u2_u7_u4_n101 ) , .ZN( u2_u7_u4_n158 ) , .A2( u2_u7_u4_n99 ) );
  AOI21_X1 u2_u7_u4_U51 (.ZN( u2_u7_u4_n127 ) , .A( u2_u7_u4_n136 ) , .B2( u2_u7_u4_n150 ) , .B1( u2_u7_u4_n180 ) );
  INV_X1 u2_u7_u4_U52 (.A( u2_u7_u4_n160 ) , .ZN( u2_u7_u4_n180 ) );
  NAND2_X1 u2_u7_u4_U53 (.A2( u2_u7_u4_n104 ) , .A1( u2_u7_u4_n105 ) , .ZN( u2_u7_u4_n146 ) );
  NAND2_X1 u2_u7_u4_U54 (.A2( u2_u7_u4_n101 ) , .A1( u2_u7_u4_n102 ) , .ZN( u2_u7_u4_n160 ) );
  NAND2_X1 u2_u7_u4_U55 (.ZN( u2_u7_u4_n134 ) , .A1( u2_u7_u4_n98 ) , .A2( u2_u7_u4_n99 ) );
  NAND2_X1 u2_u7_u4_U56 (.A1( u2_u7_u4_n103 ) , .A2( u2_u7_u4_n104 ) , .ZN( u2_u7_u4_n143 ) );
  NAND2_X1 u2_u7_u4_U57 (.A2( u2_u7_u4_n105 ) , .ZN( u2_u7_u4_n145 ) , .A1( u2_u7_u4_n98 ) );
  NAND2_X1 u2_u7_u4_U58 (.A1( u2_u7_u4_n100 ) , .A2( u2_u7_u4_n105 ) , .ZN( u2_u7_u4_n120 ) );
  NAND2_X1 u2_u7_u4_U59 (.A1( u2_u7_u4_n102 ) , .A2( u2_u7_u4_n104 ) , .ZN( u2_u7_u4_n148 ) );
  AOI21_X1 u2_u7_u4_U6 (.ZN( u2_u7_u4_n106 ) , .B2( u2_u7_u4_n146 ) , .B1( u2_u7_u4_n158 ) , .A( u2_u7_u4_n170 ) );
  NAND2_X1 u2_u7_u4_U60 (.A2( u2_u7_u4_n100 ) , .A1( u2_u7_u4_n103 ) , .ZN( u2_u7_u4_n157 ) );
  INV_X1 u2_u7_u4_U61 (.A( u2_u7_u4_n150 ) , .ZN( u2_u7_u4_n173 ) );
  INV_X1 u2_u7_u4_U62 (.A( u2_u7_u4_n152 ) , .ZN( u2_u7_u4_n171 ) );
  NAND2_X1 u2_u7_u4_U63 (.A1( u2_u7_u4_n100 ) , .ZN( u2_u7_u4_n118 ) , .A2( u2_u7_u4_n99 ) );
  NAND2_X1 u2_u7_u4_U64 (.A2( u2_u7_u4_n100 ) , .A1( u2_u7_u4_n102 ) , .ZN( u2_u7_u4_n144 ) );
  NAND2_X1 u2_u7_u4_U65 (.A2( u2_u7_u4_n101 ) , .A1( u2_u7_u4_n105 ) , .ZN( u2_u7_u4_n96 ) );
  INV_X1 u2_u7_u4_U66 (.A( u2_u7_u4_n128 ) , .ZN( u2_u7_u4_n174 ) );
  NAND2_X1 u2_u7_u4_U67 (.A2( u2_u7_u4_n102 ) , .ZN( u2_u7_u4_n119 ) , .A1( u2_u7_u4_n98 ) );
  NAND2_X1 u2_u7_u4_U68 (.A2( u2_u7_u4_n101 ) , .A1( u2_u7_u4_n103 ) , .ZN( u2_u7_u4_n147 ) );
  NAND2_X1 u2_u7_u4_U69 (.A2( u2_u7_u4_n104 ) , .ZN( u2_u7_u4_n113 ) , .A1( u2_u7_u4_n99 ) );
  AOI21_X1 u2_u7_u4_U7 (.ZN( u2_u7_u4_n108 ) , .B2( u2_u7_u4_n134 ) , .B1( u2_u7_u4_n155 ) , .A( u2_u7_u4_n156 ) );
  NOR2_X1 u2_u7_u4_U70 (.A2( u2_u7_X_28 ) , .ZN( u2_u7_u4_n150 ) , .A1( u2_u7_u4_n168 ) );
  NOR2_X1 u2_u7_u4_U71 (.A2( u2_u7_X_29 ) , .ZN( u2_u7_u4_n152 ) , .A1( u2_u7_u4_n169 ) );
  NOR2_X1 u2_u7_u4_U72 (.A2( u2_u7_X_26 ) , .ZN( u2_u7_u4_n100 ) , .A1( u2_u7_u4_n177 ) );
  NOR2_X1 u2_u7_u4_U73 (.A2( u2_u7_X_30 ) , .ZN( u2_u7_u4_n105 ) , .A1( u2_u7_u4_n176 ) );
  NOR2_X1 u2_u7_u4_U74 (.A2( u2_u7_X_28 ) , .A1( u2_u7_X_29 ) , .ZN( u2_u7_u4_n128 ) );
  NOR2_X1 u2_u7_u4_U75 (.A2( u2_u7_X_25 ) , .A1( u2_u7_X_26 ) , .ZN( u2_u7_u4_n98 ) );
  NOR2_X1 u2_u7_u4_U76 (.A2( u2_u7_X_27 ) , .A1( u2_u7_X_30 ) , .ZN( u2_u7_u4_n102 ) );
  AND2_X1 u2_u7_u4_U77 (.A2( u2_u7_X_25 ) , .A1( u2_u7_X_26 ) , .ZN( u2_u7_u4_n104 ) );
  AND2_X1 u2_u7_u4_U78 (.A1( u2_u7_X_30 ) , .A2( u2_u7_u4_n176 ) , .ZN( u2_u7_u4_n99 ) );
  AND2_X1 u2_u7_u4_U79 (.A1( u2_u7_X_26 ) , .ZN( u2_u7_u4_n101 ) , .A2( u2_u7_u4_n177 ) );
  AOI21_X1 u2_u7_u4_U8 (.ZN( u2_u7_u4_n109 ) , .A( u2_u7_u4_n153 ) , .B1( u2_u7_u4_n159 ) , .B2( u2_u7_u4_n184 ) );
  AND2_X1 u2_u7_u4_U80 (.A1( u2_u7_X_27 ) , .A2( u2_u7_X_30 ) , .ZN( u2_u7_u4_n103 ) );
  INV_X1 u2_u7_u4_U81 (.A( u2_u7_X_28 ) , .ZN( u2_u7_u4_n169 ) );
  INV_X1 u2_u7_u4_U82 (.A( u2_u7_X_29 ) , .ZN( u2_u7_u4_n168 ) );
  INV_X1 u2_u7_u4_U83 (.A( u2_u7_X_25 ) , .ZN( u2_u7_u4_n177 ) );
  INV_X1 u2_u7_u4_U84 (.A( u2_u7_X_27 ) , .ZN( u2_u7_u4_n176 ) );
  NAND4_X1 u2_u7_u4_U85 (.ZN( u2_out7_25 ) , .A4( u2_u7_u4_n139 ) , .A3( u2_u7_u4_n140 ) , .A2( u2_u7_u4_n141 ) , .A1( u2_u7_u4_n142 ) );
  OAI21_X1 u2_u7_u4_U86 (.A( u2_u7_u4_n128 ) , .B2( u2_u7_u4_n129 ) , .B1( u2_u7_u4_n130 ) , .ZN( u2_u7_u4_n142 ) );
  OAI21_X1 u2_u7_u4_U87 (.B2( u2_u7_u4_n131 ) , .ZN( u2_u7_u4_n141 ) , .A( u2_u7_u4_n175 ) , .B1( u2_u7_u4_n183 ) );
  NAND4_X1 u2_u7_u4_U88 (.ZN( u2_out7_14 ) , .A4( u2_u7_u4_n124 ) , .A3( u2_u7_u4_n125 ) , .A2( u2_u7_u4_n126 ) , .A1( u2_u7_u4_n127 ) );
  AOI22_X1 u2_u7_u4_U89 (.B2( u2_u7_u4_n117 ) , .ZN( u2_u7_u4_n126 ) , .A1( u2_u7_u4_n129 ) , .B1( u2_u7_u4_n152 ) , .A2( u2_u7_u4_n175 ) );
  AOI211_X1 u2_u7_u4_U9 (.B( u2_u7_u4_n136 ) , .A( u2_u7_u4_n137 ) , .C2( u2_u7_u4_n138 ) , .ZN( u2_u7_u4_n139 ) , .C1( u2_u7_u4_n182 ) );
  AOI22_X1 u2_u7_u4_U90 (.ZN( u2_u7_u4_n125 ) , .B2( u2_u7_u4_n131 ) , .A2( u2_u7_u4_n132 ) , .B1( u2_u7_u4_n138 ) , .A1( u2_u7_u4_n178 ) );
  NAND4_X1 u2_u7_u4_U91 (.ZN( u2_out7_8 ) , .A4( u2_u7_u4_n110 ) , .A3( u2_u7_u4_n111 ) , .A2( u2_u7_u4_n112 ) , .A1( u2_u7_u4_n186 ) );
  NAND2_X1 u2_u7_u4_U92 (.ZN( u2_u7_u4_n112 ) , .A2( u2_u7_u4_n130 ) , .A1( u2_u7_u4_n150 ) );
  AOI22_X1 u2_u7_u4_U93 (.ZN( u2_u7_u4_n111 ) , .B2( u2_u7_u4_n132 ) , .A1( u2_u7_u4_n152 ) , .B1( u2_u7_u4_n178 ) , .A2( u2_u7_u4_n97 ) );
  AOI22_X1 u2_u7_u4_U94 (.B2( u2_u7_u4_n149 ) , .B1( u2_u7_u4_n150 ) , .A2( u2_u7_u4_n151 ) , .A1( u2_u7_u4_n152 ) , .ZN( u2_u7_u4_n167 ) );
  NOR4_X1 u2_u7_u4_U95 (.A4( u2_u7_u4_n162 ) , .A3( u2_u7_u4_n163 ) , .A2( u2_u7_u4_n164 ) , .A1( u2_u7_u4_n165 ) , .ZN( u2_u7_u4_n166 ) );
  NAND3_X1 u2_u7_u4_U96 (.ZN( u2_out7_3 ) , .A3( u2_u7_u4_n166 ) , .A1( u2_u7_u4_n167 ) , .A2( u2_u7_u4_n186 ) );
  NAND3_X1 u2_u7_u4_U97 (.A3( u2_u7_u4_n146 ) , .A2( u2_u7_u4_n147 ) , .A1( u2_u7_u4_n148 ) , .ZN( u2_u7_u4_n149 ) );
  NAND3_X1 u2_u7_u4_U98 (.A3( u2_u7_u4_n143 ) , .A2( u2_u7_u4_n144 ) , .A1( u2_u7_u4_n145 ) , .ZN( u2_u7_u4_n151 ) );
  NAND3_X1 u2_u7_u4_U99 (.A3( u2_u7_u4_n121 ) , .ZN( u2_u7_u4_n122 ) , .A2( u2_u7_u4_n144 ) , .A1( u2_u7_u4_n154 ) );
  INV_X1 u2_u7_u5_U10 (.A( u2_u7_u5_n121 ) , .ZN( u2_u7_u5_n177 ) );
  NOR3_X1 u2_u7_u5_U100 (.A3( u2_u7_u5_n141 ) , .A1( u2_u7_u5_n142 ) , .ZN( u2_u7_u5_n143 ) , .A2( u2_u7_u5_n191 ) );
  NAND4_X1 u2_u7_u5_U101 (.ZN( u2_out7_4 ) , .A4( u2_u7_u5_n112 ) , .A2( u2_u7_u5_n113 ) , .A1( u2_u7_u5_n114 ) , .A3( u2_u7_u5_n195 ) );
  AOI211_X1 u2_u7_u5_U102 (.A( u2_u7_u5_n110 ) , .C1( u2_u7_u5_n111 ) , .ZN( u2_u7_u5_n112 ) , .B( u2_u7_u5_n118 ) , .C2( u2_u7_u5_n177 ) );
  AOI222_X1 u2_u7_u5_U103 (.ZN( u2_u7_u5_n113 ) , .A1( u2_u7_u5_n131 ) , .C1( u2_u7_u5_n148 ) , .B2( u2_u7_u5_n174 ) , .C2( u2_u7_u5_n178 ) , .A2( u2_u7_u5_n179 ) , .B1( u2_u7_u5_n99 ) );
  NAND3_X1 u2_u7_u5_U104 (.A2( u2_u7_u5_n154 ) , .A3( u2_u7_u5_n158 ) , .A1( u2_u7_u5_n161 ) , .ZN( u2_u7_u5_n99 ) );
  NOR2_X1 u2_u7_u5_U11 (.ZN( u2_u7_u5_n160 ) , .A2( u2_u7_u5_n173 ) , .A1( u2_u7_u5_n177 ) );
  INV_X1 u2_u7_u5_U12 (.A( u2_u7_u5_n150 ) , .ZN( u2_u7_u5_n174 ) );
  AOI21_X1 u2_u7_u5_U13 (.A( u2_u7_u5_n160 ) , .B2( u2_u7_u5_n161 ) , .ZN( u2_u7_u5_n162 ) , .B1( u2_u7_u5_n192 ) );
  INV_X1 u2_u7_u5_U14 (.A( u2_u7_u5_n159 ) , .ZN( u2_u7_u5_n192 ) );
  AOI21_X1 u2_u7_u5_U15 (.A( u2_u7_u5_n156 ) , .B2( u2_u7_u5_n157 ) , .B1( u2_u7_u5_n158 ) , .ZN( u2_u7_u5_n163 ) );
  AOI21_X1 u2_u7_u5_U16 (.B2( u2_u7_u5_n139 ) , .B1( u2_u7_u5_n140 ) , .ZN( u2_u7_u5_n141 ) , .A( u2_u7_u5_n150 ) );
  OAI21_X1 u2_u7_u5_U17 (.A( u2_u7_u5_n133 ) , .B2( u2_u7_u5_n134 ) , .B1( u2_u7_u5_n135 ) , .ZN( u2_u7_u5_n142 ) );
  OAI21_X1 u2_u7_u5_U18 (.ZN( u2_u7_u5_n133 ) , .B2( u2_u7_u5_n147 ) , .A( u2_u7_u5_n173 ) , .B1( u2_u7_u5_n188 ) );
  NAND2_X1 u2_u7_u5_U19 (.A2( u2_u7_u5_n119 ) , .A1( u2_u7_u5_n123 ) , .ZN( u2_u7_u5_n137 ) );
  INV_X1 u2_u7_u5_U20 (.A( u2_u7_u5_n155 ) , .ZN( u2_u7_u5_n194 ) );
  NAND2_X1 u2_u7_u5_U21 (.A1( u2_u7_u5_n121 ) , .ZN( u2_u7_u5_n132 ) , .A2( u2_u7_u5_n172 ) );
  NAND2_X1 u2_u7_u5_U22 (.A2( u2_u7_u5_n122 ) , .ZN( u2_u7_u5_n136 ) , .A1( u2_u7_u5_n154 ) );
  NAND2_X1 u2_u7_u5_U23 (.A2( u2_u7_u5_n119 ) , .A1( u2_u7_u5_n120 ) , .ZN( u2_u7_u5_n159 ) );
  INV_X1 u2_u7_u5_U24 (.A( u2_u7_u5_n156 ) , .ZN( u2_u7_u5_n175 ) );
  INV_X1 u2_u7_u5_U25 (.A( u2_u7_u5_n158 ) , .ZN( u2_u7_u5_n188 ) );
  INV_X1 u2_u7_u5_U26 (.A( u2_u7_u5_n152 ) , .ZN( u2_u7_u5_n179 ) );
  INV_X1 u2_u7_u5_U27 (.A( u2_u7_u5_n140 ) , .ZN( u2_u7_u5_n182 ) );
  INV_X1 u2_u7_u5_U28 (.A( u2_u7_u5_n151 ) , .ZN( u2_u7_u5_n183 ) );
  INV_X1 u2_u7_u5_U29 (.A( u2_u7_u5_n123 ) , .ZN( u2_u7_u5_n185 ) );
  NOR2_X1 u2_u7_u5_U3 (.ZN( u2_u7_u5_n134 ) , .A1( u2_u7_u5_n183 ) , .A2( u2_u7_u5_n190 ) );
  INV_X1 u2_u7_u5_U30 (.A( u2_u7_u5_n161 ) , .ZN( u2_u7_u5_n184 ) );
  INV_X1 u2_u7_u5_U31 (.A( u2_u7_u5_n139 ) , .ZN( u2_u7_u5_n189 ) );
  INV_X1 u2_u7_u5_U32 (.A( u2_u7_u5_n157 ) , .ZN( u2_u7_u5_n190 ) );
  INV_X1 u2_u7_u5_U33 (.A( u2_u7_u5_n120 ) , .ZN( u2_u7_u5_n193 ) );
  NAND2_X1 u2_u7_u5_U34 (.ZN( u2_u7_u5_n111 ) , .A1( u2_u7_u5_n140 ) , .A2( u2_u7_u5_n155 ) );
  NOR2_X1 u2_u7_u5_U35 (.ZN( u2_u7_u5_n100 ) , .A1( u2_u7_u5_n170 ) , .A2( u2_u7_u5_n180 ) );
  INV_X1 u2_u7_u5_U36 (.A( u2_u7_u5_n117 ) , .ZN( u2_u7_u5_n196 ) );
  OAI221_X1 u2_u7_u5_U37 (.A( u2_u7_u5_n116 ) , .ZN( u2_u7_u5_n117 ) , .B2( u2_u7_u5_n119 ) , .C1( u2_u7_u5_n153 ) , .C2( u2_u7_u5_n158 ) , .B1( u2_u7_u5_n172 ) );
  AOI222_X1 u2_u7_u5_U38 (.ZN( u2_u7_u5_n116 ) , .B2( u2_u7_u5_n145 ) , .C1( u2_u7_u5_n148 ) , .A2( u2_u7_u5_n174 ) , .C2( u2_u7_u5_n177 ) , .B1( u2_u7_u5_n187 ) , .A1( u2_u7_u5_n193 ) );
  INV_X1 u2_u7_u5_U39 (.A( u2_u7_u5_n115 ) , .ZN( u2_u7_u5_n187 ) );
  INV_X1 u2_u7_u5_U4 (.A( u2_u7_u5_n138 ) , .ZN( u2_u7_u5_n191 ) );
  AOI22_X1 u2_u7_u5_U40 (.B2( u2_u7_u5_n131 ) , .A2( u2_u7_u5_n146 ) , .ZN( u2_u7_u5_n169 ) , .B1( u2_u7_u5_n174 ) , .A1( u2_u7_u5_n185 ) );
  NOR2_X1 u2_u7_u5_U41 (.A1( u2_u7_u5_n146 ) , .ZN( u2_u7_u5_n150 ) , .A2( u2_u7_u5_n173 ) );
  AOI21_X1 u2_u7_u5_U42 (.A( u2_u7_u5_n118 ) , .B2( u2_u7_u5_n145 ) , .ZN( u2_u7_u5_n168 ) , .B1( u2_u7_u5_n186 ) );
  INV_X1 u2_u7_u5_U43 (.A( u2_u7_u5_n122 ) , .ZN( u2_u7_u5_n186 ) );
  NOR2_X1 u2_u7_u5_U44 (.A1( u2_u7_u5_n146 ) , .ZN( u2_u7_u5_n152 ) , .A2( u2_u7_u5_n176 ) );
  NOR2_X1 u2_u7_u5_U45 (.A1( u2_u7_u5_n115 ) , .ZN( u2_u7_u5_n118 ) , .A2( u2_u7_u5_n153 ) );
  NOR2_X1 u2_u7_u5_U46 (.A2( u2_u7_u5_n145 ) , .ZN( u2_u7_u5_n156 ) , .A1( u2_u7_u5_n174 ) );
  NOR2_X1 u2_u7_u5_U47 (.ZN( u2_u7_u5_n121 ) , .A2( u2_u7_u5_n145 ) , .A1( u2_u7_u5_n176 ) );
  AOI22_X1 u2_u7_u5_U48 (.ZN( u2_u7_u5_n114 ) , .A2( u2_u7_u5_n137 ) , .A1( u2_u7_u5_n145 ) , .B2( u2_u7_u5_n175 ) , .B1( u2_u7_u5_n193 ) );
  OAI211_X1 u2_u7_u5_U49 (.B( u2_u7_u5_n124 ) , .A( u2_u7_u5_n125 ) , .C2( u2_u7_u5_n126 ) , .C1( u2_u7_u5_n127 ) , .ZN( u2_u7_u5_n128 ) );
  OAI21_X1 u2_u7_u5_U5 (.B2( u2_u7_u5_n136 ) , .B1( u2_u7_u5_n137 ) , .ZN( u2_u7_u5_n138 ) , .A( u2_u7_u5_n177 ) );
  NOR3_X1 u2_u7_u5_U50 (.ZN( u2_u7_u5_n127 ) , .A1( u2_u7_u5_n136 ) , .A3( u2_u7_u5_n148 ) , .A2( u2_u7_u5_n182 ) );
  OAI21_X1 u2_u7_u5_U51 (.ZN( u2_u7_u5_n124 ) , .A( u2_u7_u5_n177 ) , .B2( u2_u7_u5_n183 ) , .B1( u2_u7_u5_n189 ) );
  OAI21_X1 u2_u7_u5_U52 (.ZN( u2_u7_u5_n125 ) , .A( u2_u7_u5_n174 ) , .B2( u2_u7_u5_n185 ) , .B1( u2_u7_u5_n190 ) );
  AOI21_X1 u2_u7_u5_U53 (.A( u2_u7_u5_n153 ) , .B2( u2_u7_u5_n154 ) , .B1( u2_u7_u5_n155 ) , .ZN( u2_u7_u5_n164 ) );
  AOI21_X1 u2_u7_u5_U54 (.ZN( u2_u7_u5_n110 ) , .B1( u2_u7_u5_n122 ) , .B2( u2_u7_u5_n139 ) , .A( u2_u7_u5_n153 ) );
  INV_X1 u2_u7_u5_U55 (.A( u2_u7_u5_n153 ) , .ZN( u2_u7_u5_n176 ) );
  INV_X1 u2_u7_u5_U56 (.A( u2_u7_u5_n126 ) , .ZN( u2_u7_u5_n173 ) );
  AND2_X1 u2_u7_u5_U57 (.A2( u2_u7_u5_n104 ) , .A1( u2_u7_u5_n107 ) , .ZN( u2_u7_u5_n147 ) );
  AND2_X1 u2_u7_u5_U58 (.A2( u2_u7_u5_n104 ) , .A1( u2_u7_u5_n108 ) , .ZN( u2_u7_u5_n148 ) );
  NAND2_X1 u2_u7_u5_U59 (.A1( u2_u7_u5_n105 ) , .A2( u2_u7_u5_n106 ) , .ZN( u2_u7_u5_n158 ) );
  INV_X1 u2_u7_u5_U6 (.A( u2_u7_u5_n135 ) , .ZN( u2_u7_u5_n178 ) );
  NAND2_X1 u2_u7_u5_U60 (.A2( u2_u7_u5_n108 ) , .A1( u2_u7_u5_n109 ) , .ZN( u2_u7_u5_n139 ) );
  NAND2_X1 u2_u7_u5_U61 (.A1( u2_u7_u5_n106 ) , .A2( u2_u7_u5_n108 ) , .ZN( u2_u7_u5_n119 ) );
  NAND2_X1 u2_u7_u5_U62 (.A2( u2_u7_u5_n103 ) , .A1( u2_u7_u5_n105 ) , .ZN( u2_u7_u5_n140 ) );
  NAND2_X1 u2_u7_u5_U63 (.A2( u2_u7_u5_n104 ) , .A1( u2_u7_u5_n105 ) , .ZN( u2_u7_u5_n155 ) );
  NAND2_X1 u2_u7_u5_U64 (.A2( u2_u7_u5_n106 ) , .A1( u2_u7_u5_n107 ) , .ZN( u2_u7_u5_n122 ) );
  NAND2_X1 u2_u7_u5_U65 (.A2( u2_u7_u5_n100 ) , .A1( u2_u7_u5_n106 ) , .ZN( u2_u7_u5_n115 ) );
  NAND2_X1 u2_u7_u5_U66 (.A2( u2_u7_u5_n100 ) , .A1( u2_u7_u5_n103 ) , .ZN( u2_u7_u5_n161 ) );
  NAND2_X1 u2_u7_u5_U67 (.A1( u2_u7_u5_n105 ) , .A2( u2_u7_u5_n109 ) , .ZN( u2_u7_u5_n154 ) );
  INV_X1 u2_u7_u5_U68 (.A( u2_u7_u5_n146 ) , .ZN( u2_u7_u5_n172 ) );
  NAND2_X1 u2_u7_u5_U69 (.A1( u2_u7_u5_n103 ) , .A2( u2_u7_u5_n108 ) , .ZN( u2_u7_u5_n123 ) );
  OAI22_X1 u2_u7_u5_U7 (.B2( u2_u7_u5_n149 ) , .B1( u2_u7_u5_n150 ) , .A2( u2_u7_u5_n151 ) , .A1( u2_u7_u5_n152 ) , .ZN( u2_u7_u5_n165 ) );
  NAND2_X1 u2_u7_u5_U70 (.A2( u2_u7_u5_n103 ) , .A1( u2_u7_u5_n107 ) , .ZN( u2_u7_u5_n151 ) );
  NAND2_X1 u2_u7_u5_U71 (.A2( u2_u7_u5_n107 ) , .A1( u2_u7_u5_n109 ) , .ZN( u2_u7_u5_n120 ) );
  NAND2_X1 u2_u7_u5_U72 (.A2( u2_u7_u5_n100 ) , .A1( u2_u7_u5_n109 ) , .ZN( u2_u7_u5_n157 ) );
  AND2_X1 u2_u7_u5_U73 (.A2( u2_u7_u5_n100 ) , .A1( u2_u7_u5_n104 ) , .ZN( u2_u7_u5_n131 ) );
  INV_X1 u2_u7_u5_U74 (.A( u2_u7_u5_n102 ) , .ZN( u2_u7_u5_n195 ) );
  OAI221_X1 u2_u7_u5_U75 (.A( u2_u7_u5_n101 ) , .ZN( u2_u7_u5_n102 ) , .C2( u2_u7_u5_n115 ) , .C1( u2_u7_u5_n126 ) , .B1( u2_u7_u5_n134 ) , .B2( u2_u7_u5_n160 ) );
  OAI21_X1 u2_u7_u5_U76 (.ZN( u2_u7_u5_n101 ) , .B1( u2_u7_u5_n137 ) , .A( u2_u7_u5_n146 ) , .B2( u2_u7_u5_n147 ) );
  NOR2_X1 u2_u7_u5_U77 (.A2( u2_u7_X_34 ) , .A1( u2_u7_X_35 ) , .ZN( u2_u7_u5_n145 ) );
  NOR2_X1 u2_u7_u5_U78 (.A2( u2_u7_X_34 ) , .ZN( u2_u7_u5_n146 ) , .A1( u2_u7_u5_n171 ) );
  NOR2_X1 u2_u7_u5_U79 (.A2( u2_u7_X_31 ) , .A1( u2_u7_X_32 ) , .ZN( u2_u7_u5_n103 ) );
  NOR3_X1 u2_u7_u5_U8 (.A2( u2_u7_u5_n147 ) , .A1( u2_u7_u5_n148 ) , .ZN( u2_u7_u5_n149 ) , .A3( u2_u7_u5_n194 ) );
  NOR2_X1 u2_u7_u5_U80 (.A2( u2_u7_X_36 ) , .ZN( u2_u7_u5_n105 ) , .A1( u2_u7_u5_n180 ) );
  NOR2_X1 u2_u7_u5_U81 (.A2( u2_u7_X_33 ) , .ZN( u2_u7_u5_n108 ) , .A1( u2_u7_u5_n170 ) );
  NOR2_X1 u2_u7_u5_U82 (.A2( u2_u7_X_33 ) , .A1( u2_u7_X_36 ) , .ZN( u2_u7_u5_n107 ) );
  NOR2_X1 u2_u7_u5_U83 (.A2( u2_u7_X_31 ) , .ZN( u2_u7_u5_n104 ) , .A1( u2_u7_u5_n181 ) );
  NAND2_X1 u2_u7_u5_U84 (.A2( u2_u7_X_34 ) , .A1( u2_u7_X_35 ) , .ZN( u2_u7_u5_n153 ) );
  NAND2_X1 u2_u7_u5_U85 (.A1( u2_u7_X_34 ) , .ZN( u2_u7_u5_n126 ) , .A2( u2_u7_u5_n171 ) );
  AND2_X1 u2_u7_u5_U86 (.A1( u2_u7_X_31 ) , .A2( u2_u7_X_32 ) , .ZN( u2_u7_u5_n106 ) );
  AND2_X1 u2_u7_u5_U87 (.A1( u2_u7_X_31 ) , .ZN( u2_u7_u5_n109 ) , .A2( u2_u7_u5_n181 ) );
  INV_X1 u2_u7_u5_U88 (.A( u2_u7_X_33 ) , .ZN( u2_u7_u5_n180 ) );
  INV_X1 u2_u7_u5_U89 (.A( u2_u7_X_35 ) , .ZN( u2_u7_u5_n171 ) );
  NOR2_X1 u2_u7_u5_U9 (.ZN( u2_u7_u5_n135 ) , .A1( u2_u7_u5_n173 ) , .A2( u2_u7_u5_n176 ) );
  INV_X1 u2_u7_u5_U90 (.A( u2_u7_X_36 ) , .ZN( u2_u7_u5_n170 ) );
  INV_X1 u2_u7_u5_U91 (.A( u2_u7_X_32 ) , .ZN( u2_u7_u5_n181 ) );
  NAND4_X1 u2_u7_u5_U92 (.ZN( u2_out7_29 ) , .A4( u2_u7_u5_n129 ) , .A3( u2_u7_u5_n130 ) , .A2( u2_u7_u5_n168 ) , .A1( u2_u7_u5_n196 ) );
  AOI221_X1 u2_u7_u5_U93 (.A( u2_u7_u5_n128 ) , .ZN( u2_u7_u5_n129 ) , .C2( u2_u7_u5_n132 ) , .B2( u2_u7_u5_n159 ) , .B1( u2_u7_u5_n176 ) , .C1( u2_u7_u5_n184 ) );
  AOI222_X1 u2_u7_u5_U94 (.ZN( u2_u7_u5_n130 ) , .A2( u2_u7_u5_n146 ) , .B1( u2_u7_u5_n147 ) , .C2( u2_u7_u5_n175 ) , .B2( u2_u7_u5_n179 ) , .A1( u2_u7_u5_n188 ) , .C1( u2_u7_u5_n194 ) );
  NAND4_X1 u2_u7_u5_U95 (.ZN( u2_out7_19 ) , .A4( u2_u7_u5_n166 ) , .A3( u2_u7_u5_n167 ) , .A2( u2_u7_u5_n168 ) , .A1( u2_u7_u5_n169 ) );
  AOI22_X1 u2_u7_u5_U96 (.B2( u2_u7_u5_n145 ) , .A2( u2_u7_u5_n146 ) , .ZN( u2_u7_u5_n167 ) , .B1( u2_u7_u5_n182 ) , .A1( u2_u7_u5_n189 ) );
  NOR4_X1 u2_u7_u5_U97 (.A4( u2_u7_u5_n162 ) , .A3( u2_u7_u5_n163 ) , .A2( u2_u7_u5_n164 ) , .A1( u2_u7_u5_n165 ) , .ZN( u2_u7_u5_n166 ) );
  NAND4_X1 u2_u7_u5_U98 (.ZN( u2_out7_11 ) , .A4( u2_u7_u5_n143 ) , .A3( u2_u7_u5_n144 ) , .A2( u2_u7_u5_n169 ) , .A1( u2_u7_u5_n196 ) );
  AOI22_X1 u2_u7_u5_U99 (.A2( u2_u7_u5_n132 ) , .ZN( u2_u7_u5_n144 ) , .B2( u2_u7_u5_n145 ) , .B1( u2_u7_u5_n184 ) , .A1( u2_u7_u5_n194 ) );
  INV_X1 u2_u7_u6_U10 (.ZN( u2_u7_u6_n172 ) , .A( u2_u7_u6_n88 ) );
  OAI21_X1 u2_u7_u6_U11 (.A( u2_u7_u6_n159 ) , .B1( u2_u7_u6_n169 ) , .B2( u2_u7_u6_n173 ) , .ZN( u2_u7_u6_n90 ) );
  AOI22_X1 u2_u7_u6_U12 (.A2( u2_u7_u6_n151 ) , .B2( u2_u7_u6_n161 ) , .A1( u2_u7_u6_n167 ) , .B1( u2_u7_u6_n170 ) , .ZN( u2_u7_u6_n89 ) );
  AOI21_X1 u2_u7_u6_U13 (.ZN( u2_u7_u6_n106 ) , .A( u2_u7_u6_n142 ) , .B2( u2_u7_u6_n159 ) , .B1( u2_u7_u6_n164 ) );
  INV_X1 u2_u7_u6_U14 (.A( u2_u7_u6_n155 ) , .ZN( u2_u7_u6_n161 ) );
  INV_X1 u2_u7_u6_U15 (.A( u2_u7_u6_n128 ) , .ZN( u2_u7_u6_n164 ) );
  NAND2_X1 u2_u7_u6_U16 (.ZN( u2_u7_u6_n110 ) , .A1( u2_u7_u6_n122 ) , .A2( u2_u7_u6_n129 ) );
  NAND2_X1 u2_u7_u6_U17 (.ZN( u2_u7_u6_n124 ) , .A2( u2_u7_u6_n146 ) , .A1( u2_u7_u6_n148 ) );
  INV_X1 u2_u7_u6_U18 (.A( u2_u7_u6_n132 ) , .ZN( u2_u7_u6_n171 ) );
  AND2_X1 u2_u7_u6_U19 (.A1( u2_u7_u6_n100 ) , .ZN( u2_u7_u6_n130 ) , .A2( u2_u7_u6_n147 ) );
  INV_X1 u2_u7_u6_U20 (.A( u2_u7_u6_n127 ) , .ZN( u2_u7_u6_n173 ) );
  INV_X1 u2_u7_u6_U21 (.A( u2_u7_u6_n121 ) , .ZN( u2_u7_u6_n167 ) );
  INV_X1 u2_u7_u6_U22 (.A( u2_u7_u6_n100 ) , .ZN( u2_u7_u6_n169 ) );
  INV_X1 u2_u7_u6_U23 (.A( u2_u7_u6_n123 ) , .ZN( u2_u7_u6_n170 ) );
  INV_X1 u2_u7_u6_U24 (.A( u2_u7_u6_n113 ) , .ZN( u2_u7_u6_n168 ) );
  AND2_X1 u2_u7_u6_U25 (.A1( u2_u7_u6_n107 ) , .A2( u2_u7_u6_n119 ) , .ZN( u2_u7_u6_n133 ) );
  AND2_X1 u2_u7_u6_U26 (.A2( u2_u7_u6_n121 ) , .A1( u2_u7_u6_n122 ) , .ZN( u2_u7_u6_n131 ) );
  AND3_X1 u2_u7_u6_U27 (.ZN( u2_u7_u6_n120 ) , .A2( u2_u7_u6_n127 ) , .A1( u2_u7_u6_n132 ) , .A3( u2_u7_u6_n145 ) );
  INV_X1 u2_u7_u6_U28 (.A( u2_u7_u6_n146 ) , .ZN( u2_u7_u6_n163 ) );
  AOI222_X1 u2_u7_u6_U29 (.ZN( u2_u7_u6_n114 ) , .A1( u2_u7_u6_n118 ) , .A2( u2_u7_u6_n126 ) , .B2( u2_u7_u6_n151 ) , .C2( u2_u7_u6_n159 ) , .C1( u2_u7_u6_n168 ) , .B1( u2_u7_u6_n169 ) );
  INV_X1 u2_u7_u6_U3 (.A( u2_u7_u6_n110 ) , .ZN( u2_u7_u6_n166 ) );
  NOR2_X1 u2_u7_u6_U30 (.A1( u2_u7_u6_n162 ) , .A2( u2_u7_u6_n165 ) , .ZN( u2_u7_u6_n98 ) );
  NAND2_X1 u2_u7_u6_U31 (.A1( u2_u7_u6_n144 ) , .ZN( u2_u7_u6_n151 ) , .A2( u2_u7_u6_n158 ) );
  NAND2_X1 u2_u7_u6_U32 (.ZN( u2_u7_u6_n132 ) , .A1( u2_u7_u6_n91 ) , .A2( u2_u7_u6_n97 ) );
  AOI22_X1 u2_u7_u6_U33 (.B2( u2_u7_u6_n110 ) , .B1( u2_u7_u6_n111 ) , .A1( u2_u7_u6_n112 ) , .ZN( u2_u7_u6_n115 ) , .A2( u2_u7_u6_n161 ) );
  NAND4_X1 u2_u7_u6_U34 (.A3( u2_u7_u6_n109 ) , .ZN( u2_u7_u6_n112 ) , .A4( u2_u7_u6_n132 ) , .A2( u2_u7_u6_n147 ) , .A1( u2_u7_u6_n166 ) );
  NOR2_X1 u2_u7_u6_U35 (.ZN( u2_u7_u6_n109 ) , .A1( u2_u7_u6_n170 ) , .A2( u2_u7_u6_n173 ) );
  NOR2_X1 u2_u7_u6_U36 (.A2( u2_u7_u6_n126 ) , .ZN( u2_u7_u6_n155 ) , .A1( u2_u7_u6_n160 ) );
  NAND2_X1 u2_u7_u6_U37 (.ZN( u2_u7_u6_n146 ) , .A2( u2_u7_u6_n94 ) , .A1( u2_u7_u6_n99 ) );
  AOI21_X1 u2_u7_u6_U38 (.A( u2_u7_u6_n144 ) , .B2( u2_u7_u6_n145 ) , .B1( u2_u7_u6_n146 ) , .ZN( u2_u7_u6_n150 ) );
  AOI211_X1 u2_u7_u6_U39 (.B( u2_u7_u6_n134 ) , .A( u2_u7_u6_n135 ) , .C1( u2_u7_u6_n136 ) , .ZN( u2_u7_u6_n137 ) , .C2( u2_u7_u6_n151 ) );
  INV_X1 u2_u7_u6_U4 (.A( u2_u7_u6_n142 ) , .ZN( u2_u7_u6_n174 ) );
  NAND4_X1 u2_u7_u6_U40 (.A4( u2_u7_u6_n127 ) , .A3( u2_u7_u6_n128 ) , .A2( u2_u7_u6_n129 ) , .A1( u2_u7_u6_n130 ) , .ZN( u2_u7_u6_n136 ) );
  AOI21_X1 u2_u7_u6_U41 (.B2( u2_u7_u6_n132 ) , .B1( u2_u7_u6_n133 ) , .ZN( u2_u7_u6_n134 ) , .A( u2_u7_u6_n158 ) );
  AOI21_X1 u2_u7_u6_U42 (.B1( u2_u7_u6_n131 ) , .ZN( u2_u7_u6_n135 ) , .A( u2_u7_u6_n144 ) , .B2( u2_u7_u6_n146 ) );
  INV_X1 u2_u7_u6_U43 (.A( u2_u7_u6_n111 ) , .ZN( u2_u7_u6_n158 ) );
  NAND2_X1 u2_u7_u6_U44 (.ZN( u2_u7_u6_n127 ) , .A1( u2_u7_u6_n91 ) , .A2( u2_u7_u6_n92 ) );
  NAND2_X1 u2_u7_u6_U45 (.ZN( u2_u7_u6_n129 ) , .A2( u2_u7_u6_n95 ) , .A1( u2_u7_u6_n96 ) );
  INV_X1 u2_u7_u6_U46 (.A( u2_u7_u6_n144 ) , .ZN( u2_u7_u6_n159 ) );
  NAND2_X1 u2_u7_u6_U47 (.ZN( u2_u7_u6_n145 ) , .A2( u2_u7_u6_n97 ) , .A1( u2_u7_u6_n98 ) );
  NAND2_X1 u2_u7_u6_U48 (.ZN( u2_u7_u6_n148 ) , .A2( u2_u7_u6_n92 ) , .A1( u2_u7_u6_n94 ) );
  NAND2_X1 u2_u7_u6_U49 (.ZN( u2_u7_u6_n108 ) , .A2( u2_u7_u6_n139 ) , .A1( u2_u7_u6_n144 ) );
  NAND2_X1 u2_u7_u6_U5 (.A2( u2_u7_u6_n143 ) , .ZN( u2_u7_u6_n152 ) , .A1( u2_u7_u6_n166 ) );
  NAND2_X1 u2_u7_u6_U50 (.ZN( u2_u7_u6_n121 ) , .A2( u2_u7_u6_n95 ) , .A1( u2_u7_u6_n97 ) );
  NAND2_X1 u2_u7_u6_U51 (.ZN( u2_u7_u6_n107 ) , .A2( u2_u7_u6_n92 ) , .A1( u2_u7_u6_n95 ) );
  AND2_X1 u2_u7_u6_U52 (.ZN( u2_u7_u6_n118 ) , .A2( u2_u7_u6_n91 ) , .A1( u2_u7_u6_n99 ) );
  NAND2_X1 u2_u7_u6_U53 (.ZN( u2_u7_u6_n147 ) , .A2( u2_u7_u6_n98 ) , .A1( u2_u7_u6_n99 ) );
  NAND2_X1 u2_u7_u6_U54 (.ZN( u2_u7_u6_n128 ) , .A1( u2_u7_u6_n94 ) , .A2( u2_u7_u6_n96 ) );
  NAND2_X1 u2_u7_u6_U55 (.ZN( u2_u7_u6_n119 ) , .A2( u2_u7_u6_n95 ) , .A1( u2_u7_u6_n99 ) );
  NAND2_X1 u2_u7_u6_U56 (.ZN( u2_u7_u6_n123 ) , .A2( u2_u7_u6_n91 ) , .A1( u2_u7_u6_n96 ) );
  NAND2_X1 u2_u7_u6_U57 (.ZN( u2_u7_u6_n100 ) , .A2( u2_u7_u6_n92 ) , .A1( u2_u7_u6_n98 ) );
  NAND2_X1 u2_u7_u6_U58 (.ZN( u2_u7_u6_n122 ) , .A1( u2_u7_u6_n94 ) , .A2( u2_u7_u6_n97 ) );
  INV_X1 u2_u7_u6_U59 (.A( u2_u7_u6_n139 ) , .ZN( u2_u7_u6_n160 ) );
  AOI22_X1 u2_u7_u6_U6 (.B2( u2_u7_u6_n101 ) , .A1( u2_u7_u6_n102 ) , .ZN( u2_u7_u6_n103 ) , .B1( u2_u7_u6_n160 ) , .A2( u2_u7_u6_n161 ) );
  NAND2_X1 u2_u7_u6_U60 (.ZN( u2_u7_u6_n113 ) , .A1( u2_u7_u6_n96 ) , .A2( u2_u7_u6_n98 ) );
  NOR2_X1 u2_u7_u6_U61 (.A2( u2_u7_X_40 ) , .A1( u2_u7_X_41 ) , .ZN( u2_u7_u6_n126 ) );
  NOR2_X1 u2_u7_u6_U62 (.A2( u2_u7_X_39 ) , .A1( u2_u7_X_42 ) , .ZN( u2_u7_u6_n92 ) );
  NOR2_X1 u2_u7_u6_U63 (.A2( u2_u7_X_39 ) , .A1( u2_u7_u6_n156 ) , .ZN( u2_u7_u6_n97 ) );
  NOR2_X1 u2_u7_u6_U64 (.A2( u2_u7_X_38 ) , .A1( u2_u7_u6_n165 ) , .ZN( u2_u7_u6_n95 ) );
  NOR2_X1 u2_u7_u6_U65 (.A2( u2_u7_X_41 ) , .ZN( u2_u7_u6_n111 ) , .A1( u2_u7_u6_n157 ) );
  NOR2_X1 u2_u7_u6_U66 (.A2( u2_u7_X_37 ) , .A1( u2_u7_u6_n162 ) , .ZN( u2_u7_u6_n94 ) );
  NOR2_X1 u2_u7_u6_U67 (.A2( u2_u7_X_37 ) , .A1( u2_u7_X_38 ) , .ZN( u2_u7_u6_n91 ) );
  NAND2_X1 u2_u7_u6_U68 (.A1( u2_u7_X_41 ) , .ZN( u2_u7_u6_n144 ) , .A2( u2_u7_u6_n157 ) );
  NAND2_X1 u2_u7_u6_U69 (.A2( u2_u7_X_40 ) , .A1( u2_u7_X_41 ) , .ZN( u2_u7_u6_n139 ) );
  NOR2_X1 u2_u7_u6_U7 (.A1( u2_u7_u6_n118 ) , .ZN( u2_u7_u6_n143 ) , .A2( u2_u7_u6_n168 ) );
  AND2_X1 u2_u7_u6_U70 (.A1( u2_u7_X_39 ) , .A2( u2_u7_u6_n156 ) , .ZN( u2_u7_u6_n96 ) );
  AND2_X1 u2_u7_u6_U71 (.A1( u2_u7_X_39 ) , .A2( u2_u7_X_42 ) , .ZN( u2_u7_u6_n99 ) );
  INV_X1 u2_u7_u6_U72 (.A( u2_u7_X_40 ) , .ZN( u2_u7_u6_n157 ) );
  INV_X1 u2_u7_u6_U73 (.A( u2_u7_X_37 ) , .ZN( u2_u7_u6_n165 ) );
  INV_X1 u2_u7_u6_U74 (.A( u2_u7_X_38 ) , .ZN( u2_u7_u6_n162 ) );
  INV_X1 u2_u7_u6_U75 (.A( u2_u7_X_42 ) , .ZN( u2_u7_u6_n156 ) );
  NAND4_X1 u2_u7_u6_U76 (.ZN( u2_out7_12 ) , .A4( u2_u7_u6_n114 ) , .A3( u2_u7_u6_n115 ) , .A2( u2_u7_u6_n116 ) , .A1( u2_u7_u6_n117 ) );
  OAI22_X1 u2_u7_u6_U77 (.B2( u2_u7_u6_n111 ) , .ZN( u2_u7_u6_n116 ) , .B1( u2_u7_u6_n126 ) , .A2( u2_u7_u6_n164 ) , .A1( u2_u7_u6_n167 ) );
  OAI21_X1 u2_u7_u6_U78 (.A( u2_u7_u6_n108 ) , .ZN( u2_u7_u6_n117 ) , .B2( u2_u7_u6_n141 ) , .B1( u2_u7_u6_n163 ) );
  NAND4_X1 u2_u7_u6_U79 (.ZN( u2_out7_32 ) , .A4( u2_u7_u6_n103 ) , .A3( u2_u7_u6_n104 ) , .A2( u2_u7_u6_n105 ) , .A1( u2_u7_u6_n106 ) );
  AOI21_X1 u2_u7_u6_U8 (.B1( u2_u7_u6_n107 ) , .B2( u2_u7_u6_n132 ) , .A( u2_u7_u6_n158 ) , .ZN( u2_u7_u6_n88 ) );
  AOI22_X1 u2_u7_u6_U80 (.ZN( u2_u7_u6_n105 ) , .A2( u2_u7_u6_n108 ) , .A1( u2_u7_u6_n118 ) , .B2( u2_u7_u6_n126 ) , .B1( u2_u7_u6_n171 ) );
  AOI22_X1 u2_u7_u6_U81 (.ZN( u2_u7_u6_n104 ) , .A1( u2_u7_u6_n111 ) , .B1( u2_u7_u6_n124 ) , .B2( u2_u7_u6_n151 ) , .A2( u2_u7_u6_n93 ) );
  OAI211_X1 u2_u7_u6_U82 (.ZN( u2_out7_22 ) , .B( u2_u7_u6_n137 ) , .A( u2_u7_u6_n138 ) , .C2( u2_u7_u6_n139 ) , .C1( u2_u7_u6_n140 ) );
  AOI22_X1 u2_u7_u6_U83 (.B1( u2_u7_u6_n124 ) , .A2( u2_u7_u6_n125 ) , .A1( u2_u7_u6_n126 ) , .ZN( u2_u7_u6_n138 ) , .B2( u2_u7_u6_n161 ) );
  AND4_X1 u2_u7_u6_U84 (.A3( u2_u7_u6_n119 ) , .A1( u2_u7_u6_n120 ) , .A4( u2_u7_u6_n129 ) , .ZN( u2_u7_u6_n140 ) , .A2( u2_u7_u6_n143 ) );
  OAI211_X1 u2_u7_u6_U85 (.ZN( u2_out7_7 ) , .B( u2_u7_u6_n153 ) , .C2( u2_u7_u6_n154 ) , .C1( u2_u7_u6_n155 ) , .A( u2_u7_u6_n174 ) );
  NOR3_X1 u2_u7_u6_U86 (.A1( u2_u7_u6_n141 ) , .ZN( u2_u7_u6_n154 ) , .A3( u2_u7_u6_n164 ) , .A2( u2_u7_u6_n171 ) );
  AOI211_X1 u2_u7_u6_U87 (.B( u2_u7_u6_n149 ) , .A( u2_u7_u6_n150 ) , .C2( u2_u7_u6_n151 ) , .C1( u2_u7_u6_n152 ) , .ZN( u2_u7_u6_n153 ) );
  NAND3_X1 u2_u7_u6_U88 (.A2( u2_u7_u6_n123 ) , .ZN( u2_u7_u6_n125 ) , .A1( u2_u7_u6_n130 ) , .A3( u2_u7_u6_n131 ) );
  NAND3_X1 u2_u7_u6_U89 (.A3( u2_u7_u6_n133 ) , .ZN( u2_u7_u6_n141 ) , .A1( u2_u7_u6_n145 ) , .A2( u2_u7_u6_n148 ) );
  AOI21_X1 u2_u7_u6_U9 (.B2( u2_u7_u6_n147 ) , .B1( u2_u7_u6_n148 ) , .ZN( u2_u7_u6_n149 ) , .A( u2_u7_u6_n158 ) );
  NAND3_X1 u2_u7_u6_U90 (.ZN( u2_u7_u6_n101 ) , .A3( u2_u7_u6_n107 ) , .A2( u2_u7_u6_n121 ) , .A1( u2_u7_u6_n127 ) );
  NAND3_X1 u2_u7_u6_U91 (.ZN( u2_u7_u6_n102 ) , .A3( u2_u7_u6_n130 ) , .A2( u2_u7_u6_n145 ) , .A1( u2_u7_u6_n166 ) );
  NAND3_X1 u2_u7_u6_U92 (.A3( u2_u7_u6_n113 ) , .A1( u2_u7_u6_n119 ) , .A2( u2_u7_u6_n123 ) , .ZN( u2_u7_u6_n93 ) );
  NAND3_X1 u2_u7_u6_U93 (.ZN( u2_u7_u6_n142 ) , .A2( u2_u7_u6_n172 ) , .A3( u2_u7_u6_n89 ) , .A1( u2_u7_u6_n90 ) );
  INV_X1 u2_uk_U10 (.A( u2_uk_n188 ) , .ZN( u2_uk_n27 ) );
  OAI21_X1 u2_uk_U1023 (.ZN( u2_K8_28 ) , .A( u2_uk_n1103 ) , .B2( u2_uk_n1532 ) , .B1( u2_uk_n27 ) );
  NAND2_X1 u2_uk_U1024 (.A1( u2_uk_K_r6_51 ) , .ZN( u2_uk_n1103 ) , .A2( u2_uk_n27 ) );
  OAI21_X1 u2_uk_U1076 (.ZN( u2_K8_39 ) , .A( u2_uk_n1109 ) , .B2( u2_uk_n1526 ) , .B1( u2_uk_n202 ) );
  NAND2_X1 u2_uk_U1077 (.A1( u2_uk_K_r6_31 ) , .ZN( u2_uk_n1109 ) , .A2( u2_uk_n155 ) );
  INV_X1 u2_uk_U1081 (.ZN( u2_K13_10 ) , .A( u2_uk_n524 ) );
  INV_X1 u2_uk_U1104 (.ZN( u2_K4_3 ) , .A( u2_uk_n1035 ) );
  INV_X1 u2_uk_U1124 (.ZN( u2_K4_4 ) , .A( u2_uk_n1037 ) );
  AOI22_X1 u2_uk_U1125 (.B2( u2_uk_K_r2_13 ) , .A2( u2_uk_K_r2_18 ) , .ZN( u2_uk_n1037 ) , .B1( u2_uk_n147 ) , .A1( u2_uk_n83 ) );
  INV_X1 u2_uk_U1130 (.ZN( u2_K4_10 ) , .A( u2_uk_n1020 ) );
  AOI22_X1 u2_uk_U1131 (.B2( u2_uk_K_r2_26 ) , .A2( u2_uk_K_r2_6 ) , .ZN( u2_uk_n1020 ) , .B1( u2_uk_n231 ) , .A1( u2_uk_n60 ) );
  INV_X1 u2_uk_U1134 (.ZN( u2_K13_12 ) , .A( u2_uk_n551 ) );
  INV_X1 u2_uk_U1146 (.ZN( u2_K13_2 ) , .A( u2_uk_n665 ) );
  AOI22_X1 u2_uk_U1147 (.B2( u2_uk_K_r11_26 ) , .A2( u2_uk_K_r11_6 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n203 ) , .ZN( u2_uk_n524 ) );
  INV_X1 u2_uk_U1149 (.ZN( u2_K13_6 ) , .A( u2_uk_n681 ) );
  INV_X1 u2_uk_U1157 (.ZN( u2_K4_2 ) , .A( u2_uk_n1031 ) );
  OAI22_X1 u2_uk_U121 (.ZN( u2_K4_47 ) , .B2( u2_uk_n1350 ) , .A2( u2_uk_n1359 ) , .A1( u2_uk_n187 ) , .B1( u2_uk_n63 ) );
  INV_X1 u2_uk_U128 (.ZN( u2_K13_15 ) , .A( u2_uk_n586 ) );
  INV_X1 u2_uk_U15 (.A( u2_uk_n164 ) , .ZN( u2_uk_n93 ) );
  OAI22_X1 u2_uk_U159 (.ZN( u2_K8_19 ) , .B2( u2_uk_n1508 ) , .A2( u2_uk_n1515 ) , .A1( u2_uk_n202 ) , .B1( u2_uk_n27 ) );
  OAI21_X1 u2_uk_U171 (.ZN( u2_K8_30 ) , .A( u2_uk_n1106 ) , .B2( u2_uk_n1525 ) , .B1( u2_uk_n187 ) );
  NAND2_X1 u2_uk_U172 (.A1( u2_uk_K_r6_29 ) , .ZN( u2_uk_n1106 ) , .A2( u2_uk_n191 ) );
  INV_X1 u2_uk_U187 (.ZN( u2_K11_30 ) , .A( u2_uk_n369 ) );
  AOI22_X1 u2_uk_U188 (.B2( u2_uk_K_r9_1 ) , .A2( u2_uk_K_r9_9 ) , .B1( u2_uk_n110 ) , .A1( u2_uk_n213 ) , .ZN( u2_uk_n369 ) );
  OAI22_X1 u2_uk_U239 (.ZN( u2_K13_39 ) , .B1( u2_uk_n161 ) , .B2( u2_uk_n1725 ) , .A2( u2_uk_n1744 ) , .A1( u2_uk_n99 ) );
  OAI21_X1 u2_uk_U254 (.ZN( u2_K13_48 ) , .B1( u2_uk_n110 ) , .B2( u2_uk_n1755 ) , .A( u2_uk_n677 ) );
  OAI22_X1 u2_uk_U271 (.ZN( u2_K4_44 ) , .A1( u2_uk_n117 ) , .B2( u2_uk_n1320 ) , .A2( u2_uk_n1337 ) , .B1( u2_uk_n147 ) );
  INV_X1 u2_uk_U292 (.ZN( u2_K4_8 ) , .A( u2_uk_n1040 ) );
  OAI21_X1 u2_uk_U307 (.ZN( u2_K6_26 ) , .A( u2_uk_n1064 ) , .B2( u2_uk_n1439 ) , .B1( u2_uk_n188 ) );
  NAND2_X1 u2_uk_U308 (.A1( u2_uk_K_r4_35 ) , .ZN( u2_uk_n1064 ) , .A2( u2_uk_n191 ) );
  OAI21_X1 u2_uk_U309 (.ZN( u2_K11_26 ) , .B1( u2_uk_n102 ) , .B2( u2_uk_n1665 ) , .A( u2_uk_n363 ) );
  OAI22_X1 u2_uk_U325 (.ZN( u2_K4_46 ) , .A1( u2_uk_n128 ) , .B2( u2_uk_n1330 ) , .A2( u2_uk_n1344 ) , .B1( u2_uk_n155 ) );
  BUF_X1 u2_uk_U35 (.A( u2_uk_n164 ) , .Z( u2_uk_n187 ) );
  OAI22_X1 u2_uk_U358 (.ZN( u2_K8_40 ) , .B2( u2_uk_n1525 ) , .A2( u2_uk_n1531 ) , .A1( u2_uk_n182 ) , .B1( u2_uk_n93 ) );
  OAI22_X1 u2_uk_U371 (.ZN( u2_K11_28 ) , .B1( u2_uk_n148 ) , .B2( u2_uk_n1642 ) , .A2( u2_uk_n1674 ) , .A1( u2_uk_n93 ) );
  OAI22_X1 u2_uk_U372 (.ZN( u2_K6_28 ) , .B2( u2_uk_n1420 ) , .A2( u2_uk_n1447 ) , .A1( u2_uk_n220 ) , .B1( u2_uk_n60 ) );
  OAI21_X1 u2_uk_U388 (.ZN( u2_K4_1 ) , .A( u2_uk_n1023 ) , .B2( u2_uk_n1323 ) , .B1( u2_uk_n208 ) );
  NAND2_X1 u2_uk_U389 (.A1( u2_uk_K_r2_25 ) , .ZN( u2_uk_n1023 ) , .A2( u2_uk_n214 ) );
  OAI22_X1 u2_uk_U395 (.ZN( u2_K13_16 ) , .B2( u2_uk_n1731 ) , .A2( u2_uk_n1736 ) , .B1( u2_uk_n223 ) , .A1( u2_uk_n99 ) );
  INV_X1 u2_uk_U4 (.ZN( u2_uk_n118 ) , .A( u2_uk_n187 ) );
  OAI22_X1 u2_uk_U411 (.ZN( u2_K13_9 ) , .A1( u2_uk_n145 ) , .B2( u2_uk_n1731 ) , .A2( u2_uk_n1743 ) , .B1( u2_uk_n63 ) );
  OAI22_X1 u2_uk_U415 (.ZN( u2_K4_9 ) , .A1( u2_uk_n118 ) , .B2( u2_uk_n1329 ) , .A2( u2_uk_n1339 ) , .B1( u2_uk_n238 ) );
  INV_X1 u2_uk_U418 (.ZN( u2_K8_37 ) , .A( u2_uk_n1108 ) );
  AOI22_X1 u2_uk_U419 (.B2( u2_uk_K_r6_14 ) , .A2( u2_uk_K_r6_7 ) , .ZN( u2_uk_n1108 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n162 ) );
  OAI22_X1 u2_uk_U456 (.ZN( u2_K8_33 ) , .B2( u2_uk_n1498 ) , .A2( u2_uk_n1503 ) , .A1( u2_uk_n188 ) , .B1( u2_uk_n27 ) );
  OAI21_X1 u2_uk_U478 (.ZN( u2_K6_29 ) , .A( u2_uk_n1065 ) , .B2( u2_uk_n1412 ) , .B1( u2_uk_n161 ) );
  NAND2_X1 u2_uk_U479 (.A1( u2_uk_K_r4_0 ) , .ZN( u2_uk_n1065 ) , .A2( u2_uk_n191 ) );
  INV_X1 u2_uk_U491 (.ZN( u2_K8_29 ) , .A( u2_uk_n1104 ) );
  OAI21_X1 u2_uk_U509 (.ZN( u2_K13_17 ) , .B2( u2_uk_n1743 ) , .A( u2_uk_n587 ) , .B1( u2_uk_n60 ) );
  NAND2_X1 u2_uk_U510 (.A1( u2_uk_K_r11_27 ) , .ZN( u2_uk_n587 ) , .A2( u2_uk_n60 ) );
  OAI22_X1 u2_uk_U529 (.ZN( u2_K4_12 ) , .A1( u2_uk_n109 ) , .B2( u2_uk_n1341 ) , .A2( u2_uk_n1361 ) , .B1( u2_uk_n230 ) );
  INV_X1 u2_uk_U56 (.ZN( u2_K8_34 ) , .A( u2_uk_n1107 ) );
  OAI22_X1 u2_uk_U568 (.ZN( u2_K8_36 ) , .A1( u2_uk_n146 ) , .B2( u2_uk_n1524 ) , .A2( u2_uk_n1530 ) , .B1( u2_uk_n27 ) );
  OAI22_X1 u2_uk_U597 (.ZN( u2_K8_22 ) , .B2( u2_uk_n1529 ) , .A2( u2_uk_n1535 ) , .A1( u2_uk_n220 ) , .B1( u2_uk_n27 ) );
  OAI22_X1 u2_uk_U606 (.ZN( u2_K8_35 ) , .B2( u2_uk_n1511 ) , .A2( u2_uk_n1517 ) , .A1( u2_uk_n203 ) , .B1( u2_uk_n27 ) );
  INV_X1 u2_uk_U630 (.ZN( u2_K13_11 ) , .A( u2_uk_n526 ) );
  OAI21_X1 u2_uk_U653 (.ZN( u2_K4_43 ) , .A( u2_uk_n1036 ) , .B1( u2_uk_n110 ) , .B2( u2_uk_n1359 ) );
  OAI21_X1 u2_uk_U667 (.ZN( u2_K13_43 ) , .B2( u2_uk_n1762 ) , .B1( u2_uk_n187 ) , .A( u2_uk_n676 ) );
  NAND2_X1 u2_uk_U668 (.A1( u2_uk_K_r11_29 ) , .A2( u2_uk_n147 ) , .ZN( u2_uk_n676 ) );
  NAND2_X1 u2_uk_U686 (.A1( u2_uk_K_r9_33 ) , .A2( u2_uk_n27 ) , .ZN( u2_uk_n395 ) );
  OAI22_X1 u2_uk_U688 (.ZN( u2_K11_25 ) , .A1( u2_uk_n163 ) , .B2( u2_uk_n1647 ) , .A2( u2_uk_n1666 ) , .B1( u2_uk_n83 ) );
  OAI22_X1 u2_uk_U696 (.ZN( u2_K8_25 ) , .B2( u2_uk_n1533 ) , .A2( u2_uk_n1538 ) , .A1( u2_uk_n222 ) , .B1( u2_uk_n27 ) );
  INV_X1 u2_uk_U697 (.ZN( u2_K13_7 ) , .A( u2_uk_n682 ) );
  OAI22_X1 u2_uk_U715 (.ZN( u2_K8_32 ) , .B2( u2_uk_n1526 ) , .A2( u2_uk_n1533 ) , .A1( u2_uk_n238 ) , .B1( u2_uk_n27 ) );
  OAI21_X1 u2_uk_U732 (.ZN( u2_K8_42 ) , .A( u2_uk_n1112 ) , .B2( u2_uk_n1510 ) , .B1( u2_uk_n17 ) );
  OAI22_X1 u2_uk_U746 (.ZN( u2_K8_27 ) , .B2( u2_uk_n1499 ) , .A2( u2_uk_n1504 ) , .A1( u2_uk_n213 ) , .B1( u2_uk_n27 ) );
  OAI22_X1 u2_uk_U75 (.ZN( u2_K8_23 ) , .B2( u2_uk_n1513 ) , .A2( u2_uk_n1518 ) , .A1( u2_uk_n220 ) , .B1( u2_uk_n27 ) );
  OAI22_X1 u2_uk_U756 (.ZN( u2_K11_27 ) , .B1( u2_uk_n146 ) , .B2( u2_uk_n1654 ) , .A2( u2_uk_n1660 ) , .A1( u2_uk_n93 ) );
  NAND2_X1 u2_uk_U760 (.A1( u2_uk_K_r9_5 ) , .A2( u2_uk_n27 ) , .ZN( u2_uk_n346 ) );
  INV_X1 u2_uk_U787 (.ZN( u2_K13_13 ) , .A( u2_uk_n582 ) );
  AOI22_X1 u2_uk_U788 (.B2( u2_uk_K_r11_11 ) , .A2( u2_uk_K_r11_6 ) , .B1( u2_uk_n214 ) , .ZN( u2_uk_n582 ) , .A1( u2_uk_n83 ) );
  OAI21_X1 u2_uk_U795 (.ZN( u2_K13_1 ) , .B1( u2_uk_n109 ) , .B2( u2_uk_n1727 ) , .A( u2_uk_n603 ) );
  NAND2_X1 u2_uk_U796 (.A1( u2_uk_K_r11_25 ) , .ZN( u2_uk_n603 ) , .A2( u2_uk_n93 ) );
  OAI21_X1 u2_uk_U812 (.ZN( u2_K13_18 ) , .B2( u2_uk_n1750 ) , .B1( u2_uk_n187 ) , .A( u2_uk_n590 ) );
  NAND2_X1 u2_uk_U813 (.A1( u2_uk_K_r11_20 ) , .A2( u2_uk_n147 ) , .ZN( u2_uk_n590 ) );
  OAI22_X1 u2_uk_U819 (.ZN( u2_K8_20 ) , .B2( u2_uk_n1521 ) , .A2( u2_uk_n1527 ) , .A1( u2_uk_n220 ) , .B1( u2_uk_n27 ) );
  OAI22_X1 u2_uk_U862 (.ZN( u2_K4_11 ) , .B2( u2_uk_n1333 ) , .A2( u2_uk_n1361 ) , .A1( u2_uk_n164 ) , .B1( u2_uk_n94 ) );
  OAI22_X1 u2_uk_U886 (.ZN( u2_K8_21 ) , .B2( u2_uk_n1522 ) , .A2( u2_uk_n1528 ) , .A1( u2_uk_n213 ) , .B1( u2_uk_n27 ) );
  OAI22_X1 u2_uk_U89 (.ZN( u2_K13_41 ) , .A1( u2_uk_n129 ) , .B2( u2_uk_n1723 ) , .A2( u2_uk_n1738 ) , .B1( u2_uk_n63 ) );
  OAI22_X1 u2_uk_U895 (.ZN( u2_K6_30 ) , .B2( u2_uk_n1408 ) , .A2( u2_uk_n1413 ) , .A1( u2_uk_n164 ) , .B1( u2_uk_n60 ) );
  OAI22_X1 u2_uk_U898 (.ZN( u2_K8_38 ) , .B1( u2_uk_n118 ) , .B2( u2_uk_n1530 ) , .A2( u2_uk_n1536 ) , .A1( u2_uk_n163 ) );
  OAI22_X1 u2_uk_U929 (.ZN( u2_K13_4 ) , .B2( u2_uk_n1732 ) , .A2( u2_uk_n1737 ) , .B1( u2_uk_n187 ) , .A1( u2_uk_n94 ) );
  OAI22_X1 u2_uk_U931 (.ZN( u2_K4_48 ) , .A1( u2_uk_n109 ) , .A2( u2_uk_n1325 ) , .B2( u2_uk_n1353 ) , .B1( u2_uk_n191 ) );
  OAI22_X1 u2_uk_U944 (.ZN( u2_K13_38 ) , .B1( u2_uk_n145 ) , .B2( u2_uk_n1755 ) , .A2( u2_uk_n1761 ) , .A1( u2_uk_n99 ) );
  OAI22_X1 u2_uk_U955 (.ZN( u2_K4_45 ) , .A1( u2_uk_n102 ) , .B2( u2_uk_n1321 ) , .A2( u2_uk_n1360 ) , .B1( u2_uk_n155 ) );
  INV_X1 u2_uk_U96 (.ZN( u2_K13_5 ) , .A( u2_uk_n678 ) );
  AOI22_X1 u2_uk_U97 (.B2( u2_uk_K_r11_48 ) , .A2( u2_uk_K_r11_53 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n203 ) , .ZN( u2_uk_n678 ) );
  AOI22_X1 u2_uk_U974 (.B2( u2_uk_K_r11_19 ) , .A2( u2_uk_K_r11_24 ) , .B1( u2_uk_n118 ) , .A1( u2_uk_n187 ) , .ZN( u2_uk_n681 ) );
  OAI21_X1 u2_uk_U985 (.ZN( u2_K4_5 ) , .A( u2_uk_n1038 ) , .B2( u2_uk_n1356 ) , .B1( u2_uk_n27 ) );
endmodule

