module aes_aes_die_3 ( sa02_0, sa02_1, sa02_2, sa02_3, sa02_4, sa02_5, sa02_6, sa02_7, sa21_0, 
       sa21_1, sa21_2, sa21_3, sa21_4, sa21_5, sa21_6, sa21_7, sa23_0, sa23_1, 
       sa23_2, sa23_3, sa23_4, sa23_5, sa23_6, sa23_7, sa30_0, sa30_1, sa30_2, 
       sa30_3, sa30_4, sa30_5, sa30_6, sa30_7, sa32_0, sa32_1, sa32_2, sa32_3, 
       sa32_4, sa32_5, sa32_6, sa32_7, u0_n268, u0_n270, u0_n272, u0_n274, w3_10, 
       w3_11, w3_8, w3_9, sa02_sr_0, sa02_sr_1, sa02_sr_2, sa02_sr_3, sa02_sr_4, sa02_sr_5, sa02_sr_6, sa02_sr_7, sa21_sr_0, 
        sa21_sr_1, sa21_sr_2, sa21_sr_3, sa21_sr_4, sa21_sr_5, sa21_sr_6, sa21_sr_7, sa23_sr_0, sa23_sr_1, 
        sa23_sr_2, sa23_sr_3, sa23_sr_4, sa23_sr_5, sa23_sr_6, sa23_sr_7, sa31_sr_0, sa31_sr_1, sa31_sr_2, 
        sa31_sr_3, sa31_sr_4, sa31_sr_5, sa31_sr_6, sa31_sr_7, sa33_sr_0, sa33_sr_1, sa33_sr_2, sa33_sr_3, 
        sa33_sr_4, sa33_sr_5, sa33_sr_6, sa33_sr_7, u0_subword_16, u0_subword_17, u0_subword_18, u0_subword_19, u0_subword_20, 
        u0_subword_21, u0_subword_22, u0_subword_23 );
  input sa02_0, sa02_1, sa02_2, sa02_3, sa02_4, sa02_5, sa02_6, sa02_7, sa21_0, 
        sa21_1, sa21_2, sa21_3, sa21_4, sa21_5, sa21_6, sa21_7, sa23_0, sa23_1, 
        sa23_2, sa23_3, sa23_4, sa23_5, sa23_6, sa23_7, sa30_0, sa30_1, sa30_2, 
        sa30_3, sa30_4, sa30_5, sa30_6, sa30_7, sa32_0, sa32_1, sa32_2, sa32_3, 
        sa32_4, sa32_5, sa32_6, sa32_7, u0_n268, u0_n270, u0_n272, u0_n274, w3_10, 
        w3_11, w3_8, w3_9;
  output sa02_sr_0, sa02_sr_1, sa02_sr_2, sa02_sr_3, sa02_sr_4, sa02_sr_5, sa02_sr_6, sa02_sr_7, sa21_sr_0, 
        sa21_sr_1, sa21_sr_2, sa21_sr_3, sa21_sr_4, sa21_sr_5, sa21_sr_6, sa21_sr_7, sa23_sr_0, sa23_sr_1, 
        sa23_sr_2, sa23_sr_3, sa23_sr_4, sa23_sr_5, sa23_sr_6, sa23_sr_7, sa31_sr_0, sa31_sr_1, sa31_sr_2, 
        sa31_sr_3, sa31_sr_4, sa31_sr_5, sa31_sr_6, sa31_sr_7, sa33_sr_0, sa33_sr_1, sa33_sr_2, sa33_sr_3, 
        sa33_sr_4, sa33_sr_5, sa33_sr_6, sa33_sr_7, u0_subword_16, u0_subword_17, u0_subword_18, u0_subword_19, u0_subword_20, 
        u0_subword_21, u0_subword_22, u0_subword_23;
  wire u0_u1_n41, u0_u1_n438, u0_u1_n439, u0_u1_n440, u0_u1_n441, u0_u1_n442, u0_u1_n443, u0_u1_n444, u0_u1_n445, 
       u0_u1_n446, u0_u1_n447, u0_u1_n448, u0_u1_n449, u0_u1_n450, u0_u1_n451, u0_u1_n452, u0_u1_n453, u0_u1_n454, 
       u0_u1_n455, u0_u1_n456, u0_u1_n457, u0_u1_n458, u0_u1_n459, u0_u1_n460, u0_u1_n461, u0_u1_n462, u0_u1_n463, 
       u0_u1_n464, u0_u1_n465, u0_u1_n466, u0_u1_n467, u0_u1_n468, u0_u1_n469, u0_u1_n470, u0_u1_n471, u0_u1_n472, 
       u0_u1_n473, u0_u1_n474, u0_u1_n475, u0_u1_n476, u0_u1_n477, u0_u1_n478, u0_u1_n479, u0_u1_n480, u0_u1_n481, 
       u0_u1_n482, u0_u1_n483, u0_u1_n484, u0_u1_n485, u0_u1_n486, u0_u1_n487, u0_u1_n488, u0_u1_n489, u0_u1_n490, 
       u0_u1_n491, u0_u1_n492, u0_u1_n493, u0_u1_n494, u0_u1_n495, u0_u1_n496, u0_u1_n497, u0_u1_n498, u0_u1_n499, 
       u0_u1_n500, u0_u1_n501, u0_u1_n502, u0_u1_n503, u0_u1_n504, u0_u1_n505, u0_u1_n506, u0_u1_n507, u0_u1_n508, 
       u0_u1_n509, u0_u1_n510, u0_u1_n511, u0_u1_n512, u0_u1_n513, u0_u1_n514, u0_u1_n515, u0_u1_n516, u0_u1_n517, 
       u0_u1_n518, u0_u1_n519, u0_u1_n520, u0_u1_n521, u0_u1_n522, u0_u1_n523, u0_u1_n524, u0_u1_n525, u0_u1_n526, 
       u0_u1_n527, u0_u1_n528, u0_u1_n529, u0_u1_n530, u0_u1_n531, u0_u1_n532, u0_u1_n533, u0_u1_n534, u0_u1_n535, 
       u0_u1_n536, u0_u1_n537, u0_u1_n538, u0_u1_n539, u0_u1_n540, u0_u1_n541, u0_u1_n542, u0_u1_n543, u0_u1_n544, 
       u0_u1_n545, u0_u1_n546, u0_u1_n547, u0_u1_n548, u0_u1_n549, u0_u1_n550, u0_u1_n551, u0_u1_n552, u0_u1_n553, 
       u0_u1_n554, u0_u1_n555, u0_u1_n556, u0_u1_n557, u0_u1_n558, u0_u1_n559, u0_u1_n560, u0_u1_n561, u0_u1_n562, 
       u0_u1_n563, u0_u1_n564, u0_u1_n565, u0_u1_n566, u0_u1_n567, u0_u1_n568, u0_u1_n569, u0_u1_n570, u0_u1_n571, 
       u0_u1_n572, u0_u1_n573, u0_u1_n574, u0_u1_n575, u0_u1_n576, u0_u1_n577, u0_u1_n578, u0_u1_n579, u0_u1_n580, 
       u0_u1_n581, u0_u1_n582, u0_u1_n583, u0_u1_n584, u0_u1_n585, u0_u1_n586, u0_u1_n587, u0_u1_n588, u0_u1_n589, 
       u0_u1_n590, u0_u1_n591, u0_u1_n592, u0_u1_n593, u0_u1_n594, u0_u1_n595, u0_u1_n596, u0_u1_n597, u0_u1_n598, 
       u0_u1_n599, u0_u1_n600, u0_u1_n601, u0_u1_n602, u0_u1_n603, u0_u1_n604, u0_u1_n605, u0_u1_n606, u0_u1_n607, 
       u0_u1_n608, u0_u1_n609, u0_u1_n610, u0_u1_n611, u0_u1_n612, u0_u1_n613, u0_u1_n614, u0_u1_n615, u0_u1_n616, 
       u0_u1_n617, u0_u1_n618, u0_u1_n619, u0_u1_n620, u0_u1_n621, u0_u1_n622, u0_u1_n623, u0_u1_n624, u0_u1_n625, 
       u0_u1_n626, u0_u1_n627, u0_u1_n628, u0_u1_n629, u0_u1_n630, u0_u1_n631, u0_u1_n632, u0_u1_n633, u0_u1_n634, 
       u0_u1_n635, u0_u1_n636, u0_u1_n637, u0_u1_n638, u0_u1_n639, u0_u1_n640, u0_u1_n641, u0_u1_n642, u0_u1_n643, 
       u0_u1_n644, u0_u1_n645, u0_u1_n646, u0_u1_n647, u0_u1_n648, u0_u1_n649, u0_u1_n650, u0_u1_n651, u0_u1_n652, 
       u0_u1_n653, u0_u1_n654, u0_u1_n655, u0_u1_n656, u0_u1_n657, u0_u1_n658, u0_u1_n659, u0_u1_n660, u0_u1_n661, 
       u0_u1_n662, u0_u1_n663, u0_u1_n664, u0_u1_n665, u0_u1_n666, u0_u1_n667, u0_u1_n668, u0_u1_n669, u0_u1_n670, 
       u0_u1_n671, u0_u1_n672, u0_u1_n673, u0_u1_n674, u0_u1_n675, u0_u1_n676, u0_u1_n677, u0_u1_n678, u0_u1_n679, 
       u0_u1_n680, u0_u1_n681, u0_u1_n682, u0_u1_n683, u0_u1_n684, u0_u1_n685, u0_u1_n686, u0_u1_n687, u0_u1_n688, 
       u0_u1_n689, u0_u1_n690, u0_u1_n691, u0_u1_n692, u0_u1_n693, u0_u1_n694, u0_u1_n695, u0_u1_n696, u0_u1_n697, 
       u0_u1_n698, u0_u1_n699, u0_u1_n700, u0_u1_n701, u0_u1_n702, u0_u1_n703, u0_u1_n704, u0_u1_n705, u0_u1_n706, 
       u0_u1_n707, u0_u1_n708, u0_u1_n709, u0_u1_n710, u0_u1_n711, u0_u1_n712, u0_u1_n713, u0_u1_n714, u0_u1_n715, 
       u0_u1_n716, u0_u1_n717, u0_u1_n718, u0_u1_n719, u0_u1_n720, u0_u1_n721, u0_u1_n722, u0_u1_n723, u0_u1_n724, 
       u0_u1_n725, u0_u1_n726, u0_u1_n727, u0_u1_n728, u0_u1_n729, u0_u1_n730, u0_u1_n731, u0_u1_n732, u0_u1_n733, 
       u0_u1_n734, u0_u1_n735, u0_u1_n736, u0_u1_n737, u0_u1_n738, u0_u1_n739, u0_u1_n740, u0_u1_n741, u0_u1_n742, 
       u0_u1_n743, u0_u1_n744, u0_u1_n745, u0_u1_n746, u0_u1_n747, u0_u1_n748, u0_u1_n749, u0_u1_n750, u0_u1_n751, 
       u0_u1_n752, u0_u1_n753, u0_u1_n754, u0_u1_n755, u0_u1_n756, u0_u1_n757, u0_u1_n758, u0_u1_n759, u0_u1_n760, 
       u0_u1_n761, u0_u1_n762, u0_u1_n763, u0_u1_n764, u0_u1_n765, u0_u1_n766, u0_u1_n767, u0_u1_n768, u0_u1_n769, 
       u0_u1_n770, u0_u1_n771, u0_u1_n772, u0_u1_n773, u0_u1_n774, u0_u1_n775, u0_u1_n776, u0_u1_n777, u0_u1_n778, 
       u0_u1_n779, u0_u1_n780, u0_u1_n781, u0_u1_n782, u0_u1_n783, u0_u1_n784, u0_u1_n785, u0_u1_n786, u0_u1_n787, 
       u0_u1_n788, u0_u1_n789, u0_u1_n790, u0_u1_n791, u0_u1_n792, u0_u1_n793, u0_u1_n794, u0_u1_n795, u0_u1_n796, 
       u0_u1_n797, u0_u1_n798, u0_u1_n799, u0_u1_n800, u0_u1_n801, u0_u1_n802, u0_u1_n803, u0_u1_n804, u0_u1_n805, 
       u0_u1_n806, u0_u1_n807, u0_u1_n808, u0_u1_n809, u0_u1_n810, u0_u1_n811, u0_u1_n812, u0_u1_n813, u0_u1_n814, 
       u0_u1_n815, u0_u1_n816, u0_u1_n817, u0_u1_n818, u0_u1_n819, u0_u1_n820, u0_u1_n821, u0_u1_n822, u0_u1_n823, 
       u0_u1_n824, u0_u1_n825, u0_u1_n826, u0_u1_n827, u0_u1_n828, u0_u1_n829, u0_u1_n830, u0_u1_n831, u0_u1_n832, 
       u0_u1_n833, u0_u1_n834, u0_u1_n835, u0_u1_n836, u0_u1_n837, u0_u1_n838, u0_u1_n839, u0_u1_n840, u0_u1_n841, 
       u0_u1_n842, u0_u1_n843, u0_u1_n844, u0_u1_n845, u0_u1_n846, u0_u1_n847, u0_u1_n848, u0_u1_n849, u0_u1_n850, 
       u0_u1_n851, u0_u1_n852, u0_u1_n853, u0_u1_n854, u0_u1_n855, u0_u1_n856, u0_u1_n857, u0_u1_n858, u0_u1_n859, 
       u0_u1_n860, u0_u1_n861, u0_u1_n862, u0_u1_n863, u0_u1_n864, u0_u1_n865, u0_u1_n866, u0_u1_n867, u0_u1_n868, 
       u0_u1_n869, u0_u1_n870, u0_u1_n871, u0_u1_n872, u0_u1_n873, u0_u1_n874, u0_u1_n875, u0_u1_n876, u0_u1_n877, 
       us02_n438, us02_n439, us02_n440, us02_n441, us02_n442, us02_n443, us02_n444, us02_n445, us02_n446, 
       us02_n447, us02_n448, us02_n449, us02_n450, us02_n451, us02_n452, us02_n453, us02_n454, us02_n455, 
       us02_n456, us02_n457, us02_n458, us02_n459, us02_n460, us02_n461, us02_n462, us02_n463, us02_n464, 
       us02_n465, us02_n466, us02_n467, us02_n468, us02_n469, us02_n470, us02_n471, us02_n472, us02_n473, 
       us02_n474, us02_n475, us02_n476, us02_n477, us02_n478, us02_n479, us02_n480, us02_n481, us02_n482, 
       us02_n483, us02_n484, us02_n485, us02_n486, us02_n487, us02_n488, us02_n489, us02_n490, us02_n491, 
       us02_n492, us02_n493, us02_n494, us02_n495, us02_n496, us02_n497, us02_n498, us02_n499, us02_n500, 
       us02_n501, us02_n502, us02_n503, us02_n504, us02_n505, us02_n506, us02_n507, us02_n508, us02_n509, 
       us02_n510, us02_n511, us02_n512, us02_n513, us02_n514, us02_n515, us02_n516, us02_n517, us02_n518, 
       us02_n519, us02_n520, us02_n521, us02_n522, us02_n523, us02_n524, us02_n525, us02_n526, us02_n527, 
       us02_n528, us02_n529, us02_n530, us02_n531, us02_n532, us02_n533, us02_n534, us02_n535, us02_n536, 
       us02_n537, us02_n538, us02_n539, us02_n540, us02_n541, us02_n542, us02_n543, us02_n544, us02_n545, 
       us02_n546, us02_n547, us02_n548, us02_n549, us02_n550, us02_n551, us02_n552, us02_n553, us02_n554, 
       us02_n555, us02_n556, us02_n557, us02_n558, us02_n559, us02_n560, us02_n561, us02_n562, us02_n563, 
       us02_n564, us02_n565, us02_n566, us02_n567, us02_n568, us02_n569, us02_n570, us02_n571, us02_n572, 
       us02_n573, us02_n574, us02_n575, us02_n576, us02_n577, us02_n578, us02_n579, us02_n580, us02_n581, 
       us02_n582, us02_n583, us02_n584, us02_n585, us02_n586, us02_n587, us02_n588, us02_n589, us02_n590, 
       us02_n591, us02_n592, us02_n593, us02_n594, us02_n595, us02_n596, us02_n597, us02_n598, us02_n599, 
       us02_n600, us02_n601, us02_n602, us02_n603, us02_n604, us02_n605, us02_n606, us02_n607, us02_n608, 
       us02_n609, us02_n610, us02_n611, us02_n612, us02_n613, us02_n614, us02_n615, us02_n616, us02_n617, 
       us02_n618, us02_n619, us02_n620, us02_n621, us02_n622, us02_n623, us02_n624, us02_n625, us02_n626, 
       us02_n627, us02_n628, us02_n629, us02_n630, us02_n631, us02_n632, us02_n633, us02_n634, us02_n635, 
       us02_n636, us02_n637, us02_n638, us02_n639, us02_n640, us02_n641, us02_n642, us02_n643, us02_n644, 
       us02_n645, us02_n646, us02_n647, us02_n648, us02_n649, us02_n650, us02_n651, us02_n652, us02_n653, 
       us02_n654, us02_n655, us02_n656, us02_n657, us02_n658, us02_n659, us02_n660, us02_n661, us02_n662, 
       us02_n663, us02_n664, us02_n665, us02_n666, us02_n667, us02_n668, us02_n669, us02_n670, us02_n671, 
       us02_n672, us02_n673, us02_n674, us02_n675, us02_n676, us02_n677, us02_n678, us02_n679, us02_n680, 
       us02_n681, us02_n682, us02_n683, us02_n684, us02_n685, us02_n686, us02_n687, us02_n688, us02_n689, 
       us02_n690, us02_n691, us02_n692, us02_n693, us02_n694, us02_n695, us02_n696, us02_n697, us02_n698, 
       us02_n699, us02_n700, us02_n701, us02_n702, us02_n703, us02_n704, us02_n705, us02_n706, us02_n707, 
       us02_n708, us02_n709, us02_n710, us02_n711, us02_n712, us02_n713, us02_n714, us02_n715, us02_n716, 
       us02_n717, us02_n718, us02_n719, us02_n720, us02_n721, us02_n722, us02_n723, us02_n724, us02_n725, 
       us02_n726, us02_n727, us02_n728, us02_n729, us02_n730, us02_n731, us02_n732, us02_n733, us02_n734, 
       us02_n735, us02_n736, us02_n737, us02_n738, us02_n739, us02_n740, us02_n741, us02_n742, us02_n743, 
       us02_n744, us02_n745, us02_n746, us02_n747, us02_n748, us02_n749, us02_n750, us02_n751, us02_n752, 
       us02_n753, us02_n754, us02_n755, us02_n756, us02_n757, us02_n758, us02_n759, us02_n760, us02_n761, 
       us02_n762, us02_n763, us02_n764, us02_n765, us02_n766, us02_n767, us02_n768, us02_n769, us02_n770, 
       us02_n771, us02_n772, us02_n773, us02_n774, us02_n775, us02_n776, us02_n777, us02_n778, us02_n779, 
       us02_n780, us02_n781, us02_n782, us02_n783, us02_n784, us02_n785, us02_n786, us02_n787, us02_n788, 
       us02_n789, us02_n790, us02_n791, us02_n792, us02_n793, us02_n794, us02_n795, us02_n796, us02_n797, 
       us02_n798, us02_n799, us02_n800, us02_n801, us02_n802, us02_n803, us02_n804, us02_n805, us02_n806, 
       us02_n807, us02_n808, us02_n809, us02_n810, us02_n811, us02_n812, us02_n813, us02_n814, us02_n815, 
       us02_n816, us02_n817, us02_n818, us02_n819, us02_n820, us02_n821, us02_n822, us02_n823, us02_n824, 
       us02_n825, us02_n826, us02_n827, us02_n828, us02_n829, us02_n830, us02_n831, us02_n832, us02_n833, 
       us02_n834, us02_n835, us02_n836, us02_n837, us02_n838, us02_n839, us02_n840, us02_n841, us02_n842, 
       us02_n843, us02_n844, us02_n845, us02_n846, us02_n847, us02_n848, us02_n849, us02_n850, us02_n851, 
       us02_n852, us02_n853, us02_n854, us02_n855, us02_n856, us02_n857, us02_n858, us02_n859, us02_n860, 
       us02_n861, us02_n862, us02_n863, us02_n864, us02_n865, us02_n866, us02_n867, us02_n868, us02_n869, 
       us02_n870, us02_n871, us02_n872, us02_n873, us02_n874, us02_n875, us21_n438, us21_n439, us21_n440, 
       us21_n441, us21_n442, us21_n443, us21_n444, us21_n445, us21_n446, us21_n447, us21_n448, us21_n449, 
       us21_n450, us21_n451, us21_n452, us21_n453, us21_n454, us21_n455, us21_n456, us21_n457, us21_n458, 
       us21_n459, us21_n460, us21_n461, us21_n462, us21_n463, us21_n464, us21_n465, us21_n466, us21_n467, 
       us21_n468, us21_n469, us21_n470, us21_n471, us21_n472, us21_n473, us21_n474, us21_n475, us21_n476, 
       us21_n477, us21_n478, us21_n479, us21_n480, us21_n481, us21_n482, us21_n483, us21_n484, us21_n485, 
       us21_n486, us21_n487, us21_n488, us21_n489, us21_n490, us21_n491, us21_n492, us21_n493, us21_n494, 
       us21_n495, us21_n496, us21_n497, us21_n498, us21_n499, us21_n500, us21_n501, us21_n502, us21_n503, 
       us21_n504, us21_n505, us21_n506, us21_n507, us21_n508, us21_n509, us21_n510, us21_n511, us21_n512, 
       us21_n513, us21_n514, us21_n515, us21_n516, us21_n517, us21_n518, us21_n519, us21_n520, us21_n521, 
       us21_n522, us21_n523, us21_n524, us21_n525, us21_n526, us21_n527, us21_n528, us21_n529, us21_n530, 
       us21_n531, us21_n532, us21_n533, us21_n534, us21_n535, us21_n536, us21_n537, us21_n538, us21_n539, 
       us21_n540, us21_n541, us21_n542, us21_n543, us21_n544, us21_n545, us21_n546, us21_n547, us21_n548, 
       us21_n549, us21_n550, us21_n551, us21_n552, us21_n553, us21_n554, us21_n555, us21_n556, us21_n557, 
       us21_n558, us21_n559, us21_n560, us21_n561, us21_n562, us21_n563, us21_n564, us21_n565, us21_n566, 
       us21_n567, us21_n568, us21_n569, us21_n570, us21_n571, us21_n572, us21_n573, us21_n574, us21_n575, 
       us21_n576, us21_n577, us21_n578, us21_n579, us21_n580, us21_n581, us21_n582, us21_n583, us21_n584, 
       us21_n585, us21_n586, us21_n587, us21_n588, us21_n589, us21_n590, us21_n591, us21_n592, us21_n593, 
       us21_n594, us21_n595, us21_n596, us21_n597, us21_n598, us21_n599, us21_n600, us21_n601, us21_n602, 
       us21_n603, us21_n604, us21_n605, us21_n606, us21_n607, us21_n608, us21_n609, us21_n610, us21_n611, 
       us21_n612, us21_n613, us21_n614, us21_n615, us21_n616, us21_n617, us21_n618, us21_n619, us21_n620, 
       us21_n621, us21_n622, us21_n623, us21_n624, us21_n625, us21_n626, us21_n627, us21_n628, us21_n629, 
       us21_n630, us21_n631, us21_n632, us21_n633, us21_n634, us21_n635, us21_n636, us21_n637, us21_n638, 
       us21_n639, us21_n640, us21_n641, us21_n642, us21_n643, us21_n644, us21_n645, us21_n646, us21_n647, 
       us21_n648, us21_n649, us21_n650, us21_n651, us21_n652, us21_n653, us21_n654, us21_n655, us21_n656, 
       us21_n657, us21_n658, us21_n659, us21_n660, us21_n661, us21_n662, us21_n663, us21_n664, us21_n665, 
       us21_n666, us21_n667, us21_n668, us21_n669, us21_n670, us21_n671, us21_n672, us21_n673, us21_n674, 
       us21_n675, us21_n676, us21_n677, us21_n678, us21_n679, us21_n680, us21_n681, us21_n682, us21_n683, 
       us21_n684, us21_n685, us21_n686, us21_n687, us21_n688, us21_n689, us21_n690, us21_n691, us21_n692, 
       us21_n693, us21_n694, us21_n695, us21_n696, us21_n697, us21_n698, us21_n699, us21_n700, us21_n701, 
       us21_n702, us21_n703, us21_n704, us21_n705, us21_n706, us21_n707, us21_n708, us21_n709, us21_n710, 
       us21_n711, us21_n712, us21_n713, us21_n714, us21_n715, us21_n716, us21_n717, us21_n718, us21_n719, 
       us21_n720, us21_n721, us21_n722, us21_n723, us21_n724, us21_n725, us21_n726, us21_n727, us21_n728, 
       us21_n729, us21_n730, us21_n731, us21_n732, us21_n733, us21_n734, us21_n735, us21_n736, us21_n737, 
       us21_n738, us21_n739, us21_n740, us21_n741, us21_n742, us21_n743, us21_n744, us21_n745, us21_n746, 
       us21_n747, us21_n748, us21_n749, us21_n750, us21_n751, us21_n752, us21_n753, us21_n754, us21_n755, 
       us21_n756, us21_n757, us21_n758, us21_n759, us21_n760, us21_n761, us21_n762, us21_n763, us21_n764, 
       us21_n765, us21_n766, us21_n767, us21_n768, us21_n769, us21_n770, us21_n771, us21_n772, us21_n773, 
       us21_n774, us21_n775, us21_n776, us21_n777, us21_n778, us21_n779, us21_n780, us21_n781, us21_n782, 
       us21_n783, us21_n784, us21_n785, us21_n786, us21_n787, us21_n788, us21_n789, us21_n790, us21_n791, 
       us21_n792, us21_n793, us21_n794, us21_n795, us21_n796, us21_n797, us21_n798, us21_n799, us21_n800, 
       us21_n801, us21_n802, us21_n803, us21_n804, us21_n805, us21_n806, us21_n807, us21_n808, us21_n809, 
       us21_n810, us21_n811, us21_n812, us21_n813, us21_n814, us21_n815, us21_n816, us21_n817, us21_n818, 
       us21_n819, us21_n820, us21_n821, us21_n822, us21_n823, us21_n824, us21_n825, us21_n826, us21_n827, 
       us21_n828, us21_n829, us21_n830, us21_n831, us21_n832, us21_n833, us21_n834, us21_n835, us21_n836, 
       us21_n837, us21_n838, us21_n839, us21_n840, us21_n841, us21_n842, us21_n843, us21_n844, us21_n845, 
       us21_n846, us21_n847, us21_n848, us21_n849, us21_n850, us21_n851, us21_n852, us21_n853, us21_n854, 
       us21_n855, us21_n856, us21_n857, us21_n858, us21_n859, us21_n860, us21_n861, us21_n862, us21_n863, 
       us21_n864, us21_n865, us21_n866, us21_n867, us21_n868, us21_n869, us21_n870, us21_n871, us21_n872, 
       us21_n873, us21_n874, us23_n438, us23_n439, us23_n440, us23_n441, us23_n442, us23_n443, us23_n444, 
       us23_n445, us23_n446, us23_n447, us23_n448, us23_n449, us23_n450, us23_n451, us23_n452, us23_n453, 
       us23_n454, us23_n455, us23_n456, us23_n457, us23_n458, us23_n459, us23_n460, us23_n461, us23_n462, 
       us23_n463, us23_n464, us23_n465, us23_n466, us23_n467, us23_n468, us23_n469, us23_n470, us23_n471, 
       us23_n472, us23_n473, us23_n474, us23_n475, us23_n476, us23_n477, us23_n478, us23_n479, us23_n480, 
       us23_n481, us23_n482, us23_n483, us23_n484, us23_n485, us23_n486, us23_n487, us23_n488, us23_n489, 
       us23_n490, us23_n491, us23_n492, us23_n493, us23_n494, us23_n495, us23_n496, us23_n497, us23_n498, 
       us23_n499, us23_n500, us23_n501, us23_n502, us23_n503, us23_n504, us23_n505, us23_n506, us23_n507, 
       us23_n508, us23_n509, us23_n510, us23_n511, us23_n512, us23_n513, us23_n514, us23_n515, us23_n516, 
       us23_n517, us23_n518, us23_n519, us23_n520, us23_n521, us23_n522, us23_n523, us23_n524, us23_n525, 
       us23_n526, us23_n527, us23_n528, us23_n529, us23_n530, us23_n531, us23_n532, us23_n533, us23_n534, 
       us23_n535, us23_n536, us23_n537, us23_n538, us23_n539, us23_n540, us23_n541, us23_n542, us23_n543, 
       us23_n544, us23_n545, us23_n546, us23_n547, us23_n548, us23_n549, us23_n550, us23_n551, us23_n552, 
       us23_n553, us23_n554, us23_n555, us23_n556, us23_n557, us23_n558, us23_n559, us23_n560, us23_n561, 
       us23_n562, us23_n563, us23_n564, us23_n565, us23_n566, us23_n567, us23_n568, us23_n569, us23_n570, 
       us23_n571, us23_n572, us23_n573, us23_n574, us23_n575, us23_n576, us23_n577, us23_n578, us23_n579, 
       us23_n580, us23_n581, us23_n582, us23_n583, us23_n584, us23_n585, us23_n586, us23_n587, us23_n588, 
       us23_n589, us23_n590, us23_n591, us23_n592, us23_n593, us23_n594, us23_n595, us23_n596, us23_n597, 
       us23_n598, us23_n599, us23_n600, us23_n601, us23_n602, us23_n603, us23_n604, us23_n605, us23_n606, 
       us23_n607, us23_n608, us23_n609, us23_n610, us23_n611, us23_n612, us23_n613, us23_n614, us23_n615, 
       us23_n616, us23_n617, us23_n618, us23_n619, us23_n620, us23_n621, us23_n622, us23_n623, us23_n624, 
       us23_n625, us23_n626, us23_n627, us23_n628, us23_n629, us23_n630, us23_n631, us23_n632, us23_n633, 
       us23_n634, us23_n635, us23_n636, us23_n637, us23_n638, us23_n639, us23_n640, us23_n641, us23_n642, 
       us23_n643, us23_n644, us23_n645, us23_n646, us23_n647, us23_n648, us23_n649, us23_n650, us23_n651, 
       us23_n652, us23_n653, us23_n654, us23_n655, us23_n656, us23_n657, us23_n658, us23_n659, us23_n660, 
       us23_n661, us23_n662, us23_n663, us23_n664, us23_n665, us23_n666, us23_n667, us23_n668, us23_n669, 
       us23_n670, us23_n671, us23_n672, us23_n673, us23_n674, us23_n675, us23_n676, us23_n677, us23_n678, 
       us23_n679, us23_n680, us23_n681, us23_n682, us23_n683, us23_n684, us23_n685, us23_n686, us23_n687, 
       us23_n688, us23_n689, us23_n690, us23_n691, us23_n692, us23_n693, us23_n694, us23_n695, us23_n696, 
       us23_n697, us23_n698, us23_n699, us23_n700, us23_n701, us23_n702, us23_n703, us23_n704, us23_n705, 
       us23_n706, us23_n707, us23_n708, us23_n709, us23_n710, us23_n711, us23_n712, us23_n713, us23_n714, 
       us23_n715, us23_n716, us23_n717, us23_n718, us23_n719, us23_n720, us23_n721, us23_n722, us23_n723, 
       us23_n724, us23_n725, us23_n726, us23_n727, us23_n728, us23_n729, us23_n730, us23_n731, us23_n732, 
       us23_n733, us23_n734, us23_n735, us23_n736, us23_n737, us23_n738, us23_n739, us23_n740, us23_n741, 
       us23_n742, us23_n743, us23_n744, us23_n745, us23_n746, us23_n747, us23_n748, us23_n749, us23_n750, 
       us23_n751, us23_n752, us23_n753, us23_n754, us23_n755, us23_n756, us23_n757, us23_n758, us23_n759, 
       us23_n760, us23_n761, us23_n762, us23_n763, us23_n764, us23_n765, us23_n766, us23_n767, us23_n768, 
       us23_n769, us23_n770, us23_n771, us23_n772, us23_n773, us23_n774, us23_n775, us23_n776, us23_n777, 
       us23_n778, us23_n779, us23_n780, us23_n781, us23_n782, us23_n783, us23_n784, us23_n785, us23_n786, 
       us23_n787, us23_n788, us23_n789, us23_n790, us23_n791, us23_n792, us23_n793, us23_n794, us23_n795, 
       us23_n796, us23_n797, us23_n798, us23_n799, us23_n800, us23_n801, us23_n802, us23_n803, us23_n804, 
       us23_n805, us23_n806, us23_n807, us23_n808, us23_n809, us23_n810, us23_n811, us23_n812, us23_n813, 
       us23_n814, us23_n815, us23_n816, us23_n817, us23_n818, us23_n819, us23_n820, us23_n821, us23_n822, 
       us23_n823, us23_n824, us23_n825, us23_n826, us23_n827, us23_n828, us23_n829, us23_n830, us23_n831, 
       us23_n832, us23_n833, us23_n834, us23_n835, us23_n836, us23_n837, us23_n838, us23_n839, us23_n840, 
       us23_n841, us23_n842, us23_n843, us23_n844, us23_n845, us23_n846, us23_n847, us23_n848, us23_n849, 
       us23_n850, us23_n851, us23_n852, us23_n853, us23_n854, us23_n855, us23_n856, us23_n857, us23_n858, 
       us23_n859, us23_n860, us23_n861, us23_n862, us23_n863, us23_n864, us23_n865, us23_n866, us23_n867, 
       us23_n868, us23_n869, us23_n870, us23_n871, us23_n872, us23_n873, us23_n874, us23_n875, us30_n438, 
       us30_n439, us30_n440, us30_n441, us30_n442, us30_n443, us30_n444, us30_n445, us30_n446, us30_n447, 
       us30_n448, us30_n449, us30_n450, us30_n451, us30_n452, us30_n453, us30_n454, us30_n455, us30_n456, 
       us30_n457, us30_n458, us30_n459, us30_n460, us30_n461, us30_n462, us30_n463, us30_n464, us30_n465, 
       us30_n466, us30_n467, us30_n468, us30_n469, us30_n470, us30_n471, us30_n472, us30_n473, us30_n474, 
       us30_n475, us30_n476, us30_n477, us30_n478, us30_n479, us30_n480, us30_n481, us30_n482, us30_n483, 
       us30_n484, us30_n485, us30_n486, us30_n487, us30_n488, us30_n489, us30_n490, us30_n491, us30_n492, 
       us30_n493, us30_n494, us30_n495, us30_n496, us30_n497, us30_n498, us30_n499, us30_n500, us30_n501, 
       us30_n502, us30_n503, us30_n504, us30_n505, us30_n506, us30_n507, us30_n508, us30_n509, us30_n510, 
       us30_n511, us30_n512, us30_n513, us30_n514, us30_n515, us30_n516, us30_n517, us30_n518, us30_n519, 
       us30_n520, us30_n521, us30_n522, us30_n523, us30_n524, us30_n525, us30_n526, us30_n527, us30_n528, 
       us30_n529, us30_n530, us30_n531, us30_n532, us30_n533, us30_n534, us30_n535, us30_n536, us30_n537, 
       us30_n538, us30_n539, us30_n540, us30_n541, us30_n542, us30_n543, us30_n544, us30_n545, us30_n546, 
       us30_n547, us30_n548, us30_n549, us30_n550, us30_n551, us30_n552, us30_n553, us30_n554, us30_n555, 
       us30_n556, us30_n557, us30_n558, us30_n559, us30_n560, us30_n561, us30_n562, us30_n563, us30_n564, 
       us30_n565, us30_n566, us30_n567, us30_n568, us30_n569, us30_n570, us30_n571, us30_n572, us30_n573, 
       us30_n574, us30_n575, us30_n576, us30_n577, us30_n578, us30_n579, us30_n580, us30_n581, us30_n582, 
       us30_n583, us30_n584, us30_n585, us30_n586, us30_n587, us30_n588, us30_n589, us30_n590, us30_n591, 
       us30_n592, us30_n593, us30_n594, us30_n595, us30_n596, us30_n597, us30_n598, us30_n599, us30_n600, 
       us30_n601, us30_n602, us30_n603, us30_n604, us30_n605, us30_n606, us30_n607, us30_n608, us30_n609, 
       us30_n610, us30_n611, us30_n612, us30_n613, us30_n614, us30_n615, us30_n616, us30_n617, us30_n618, 
       us30_n619, us30_n620, us30_n621, us30_n622, us30_n623, us30_n624, us30_n625, us30_n626, us30_n627, 
       us30_n628, us30_n629, us30_n630, us30_n631, us30_n632, us30_n633, us30_n634, us30_n635, us30_n636, 
       us30_n637, us30_n638, us30_n639, us30_n640, us30_n641, us30_n642, us30_n643, us30_n644, us30_n645, 
       us30_n646, us30_n647, us30_n648, us30_n649, us30_n650, us30_n651, us30_n652, us30_n653, us30_n654, 
       us30_n655, us30_n656, us30_n657, us30_n658, us30_n659, us30_n660, us30_n661, us30_n662, us30_n663, 
       us30_n664, us30_n665, us30_n666, us30_n667, us30_n668, us30_n669, us30_n670, us30_n671, us30_n672, 
       us30_n673, us30_n674, us30_n675, us30_n676, us30_n677, us30_n678, us30_n679, us30_n680, us30_n681, 
       us30_n682, us30_n683, us30_n684, us30_n685, us30_n686, us30_n687, us30_n688, us30_n689, us30_n690, 
       us30_n691, us30_n692, us30_n693, us30_n694, us30_n695, us30_n696, us30_n697, us30_n698, us30_n699, 
       us30_n700, us30_n701, us30_n702, us30_n703, us30_n704, us30_n705, us30_n706, us30_n707, us30_n708, 
       us30_n709, us30_n710, us30_n711, us30_n712, us30_n713, us30_n714, us30_n715, us30_n716, us30_n717, 
       us30_n718, us30_n719, us30_n720, us30_n721, us30_n722, us30_n723, us30_n724, us30_n725, us30_n726, 
       us30_n727, us30_n728, us30_n729, us30_n730, us30_n731, us30_n732, us30_n733, us30_n734, us30_n735, 
       us30_n736, us30_n737, us30_n738, us30_n739, us30_n740, us30_n741, us30_n742, us30_n743, us30_n744, 
       us30_n745, us30_n746, us30_n747, us30_n748, us30_n749, us30_n750, us30_n751, us30_n752, us30_n753, 
       us30_n754, us30_n755, us30_n756, us30_n757, us30_n758, us30_n759, us30_n760, us30_n761, us30_n762, 
       us30_n763, us30_n764, us30_n765, us30_n766, us30_n767, us30_n768, us30_n769, us30_n770, us30_n771, 
       us30_n772, us30_n773, us30_n774, us30_n775, us30_n776, us30_n777, us30_n778, us30_n779, us30_n780, 
       us30_n781, us30_n782, us30_n783, us30_n784, us30_n785, us30_n786, us30_n787, us30_n788, us30_n789, 
       us30_n790, us30_n791, us30_n792, us30_n793, us30_n794, us30_n795, us30_n796, us30_n797, us30_n798, 
       us30_n799, us30_n800, us30_n801, us30_n802, us30_n803, us30_n804, us30_n805, us30_n806, us30_n807, 
       us30_n808, us30_n809, us30_n810, us30_n811, us30_n812, us30_n813, us30_n814, us30_n815, us30_n816, 
       us30_n817, us30_n818, us30_n819, us30_n820, us30_n821, us30_n822, us30_n823, us30_n824, us30_n825, 
       us30_n826, us30_n827, us30_n828, us30_n829, us30_n830, us30_n831, us30_n832, us30_n833, us30_n834, 
       us30_n835, us30_n836, us30_n837, us30_n838, us30_n839, us30_n840, us30_n841, us30_n842, us30_n843, 
       us30_n844, us30_n845, us30_n846, us30_n847, us30_n848, us30_n849, us30_n850, us30_n851, us30_n852, 
       us30_n853, us30_n854, us30_n855, us30_n856, us30_n857, us30_n858, us30_n859, us30_n860, us30_n861, 
       us30_n862, us30_n863, us30_n864, us30_n865, us30_n866, us30_n867, us30_n868, us30_n869, us30_n870, 
       us30_n871, us30_n872, us30_n873, us30_n874, us30_n875, us30_n876, us32_n438, us32_n439, us32_n440, 
       us32_n441, us32_n442, us32_n443, us32_n444, us32_n445, us32_n446, us32_n447, us32_n448, us32_n449, 
       us32_n450, us32_n451, us32_n452, us32_n453, us32_n454, us32_n455, us32_n456, us32_n457, us32_n458, 
       us32_n459, us32_n460, us32_n461, us32_n462, us32_n463, us32_n464, us32_n465, us32_n466, us32_n467, 
       us32_n468, us32_n469, us32_n470, us32_n471, us32_n472, us32_n473, us32_n474, us32_n475, us32_n476, 
       us32_n477, us32_n478, us32_n479, us32_n480, us32_n481, us32_n482, us32_n483, us32_n484, us32_n485, 
       us32_n486, us32_n487, us32_n488, us32_n489, us32_n490, us32_n491, us32_n492, us32_n493, us32_n494, 
       us32_n495, us32_n496, us32_n497, us32_n498, us32_n499, us32_n500, us32_n501, us32_n502, us32_n503, 
       us32_n504, us32_n505, us32_n506, us32_n507, us32_n508, us32_n509, us32_n510, us32_n511, us32_n512, 
       us32_n513, us32_n514, us32_n515, us32_n516, us32_n517, us32_n518, us32_n519, us32_n520, us32_n521, 
       us32_n522, us32_n523, us32_n524, us32_n525, us32_n526, us32_n527, us32_n528, us32_n529, us32_n530, 
       us32_n531, us32_n532, us32_n533, us32_n534, us32_n535, us32_n536, us32_n537, us32_n538, us32_n539, 
       us32_n540, us32_n541, us32_n542, us32_n543, us32_n544, us32_n545, us32_n546, us32_n547, us32_n548, 
       us32_n549, us32_n550, us32_n551, us32_n552, us32_n553, us32_n554, us32_n555, us32_n556, us32_n557, 
       us32_n558, us32_n559, us32_n560, us32_n561, us32_n562, us32_n563, us32_n564, us32_n565, us32_n566, 
       us32_n567, us32_n568, us32_n569, us32_n570, us32_n571, us32_n572, us32_n573, us32_n574, us32_n575, 
       us32_n576, us32_n577, us32_n578, us32_n579, us32_n580, us32_n581, us32_n582, us32_n583, us32_n584, 
       us32_n585, us32_n586, us32_n587, us32_n588, us32_n589, us32_n590, us32_n591, us32_n592, us32_n593, 
       us32_n594, us32_n595, us32_n596, us32_n597, us32_n598, us32_n599, us32_n600, us32_n601, us32_n602, 
       us32_n603, us32_n604, us32_n605, us32_n606, us32_n607, us32_n608, us32_n609, us32_n610, us32_n611, 
       us32_n612, us32_n613, us32_n614, us32_n615, us32_n616, us32_n617, us32_n618, us32_n619, us32_n620, 
       us32_n621, us32_n622, us32_n623, us32_n624, us32_n625, us32_n626, us32_n627, us32_n628, us32_n629, 
       us32_n630, us32_n631, us32_n632, us32_n633, us32_n634, us32_n635, us32_n636, us32_n637, us32_n638, 
       us32_n639, us32_n640, us32_n641, us32_n642, us32_n643, us32_n644, us32_n645, us32_n646, us32_n647, 
       us32_n648, us32_n649, us32_n650, us32_n651, us32_n652, us32_n653, us32_n654, us32_n655, us32_n656, 
       us32_n657, us32_n658, us32_n659, us32_n660, us32_n661, us32_n662, us32_n663, us32_n664, us32_n665, 
       us32_n666, us32_n667, us32_n668, us32_n669, us32_n670, us32_n671, us32_n672, us32_n673, us32_n674, 
       us32_n675, us32_n676, us32_n677, us32_n678, us32_n679, us32_n680, us32_n681, us32_n682, us32_n683, 
       us32_n684, us32_n685, us32_n686, us32_n687, us32_n688, us32_n689, us32_n690, us32_n691, us32_n692, 
       us32_n693, us32_n694, us32_n695, us32_n696, us32_n697, us32_n698, us32_n699, us32_n700, us32_n701, 
       us32_n702, us32_n703, us32_n704, us32_n705, us32_n706, us32_n707, us32_n708, us32_n709, us32_n710, 
       us32_n711, us32_n712, us32_n713, us32_n714, us32_n715, us32_n716, us32_n717, us32_n718, us32_n719, 
       us32_n720, us32_n721, us32_n722, us32_n723, us32_n724, us32_n725, us32_n726, us32_n727, us32_n728, 
       us32_n729, us32_n730, us32_n731, us32_n732, us32_n733, us32_n734, us32_n735, us32_n736, us32_n737, 
       us32_n738, us32_n739, us32_n740, us32_n741, us32_n742, us32_n743, us32_n744, us32_n745, us32_n746, 
       us32_n747, us32_n748, us32_n749, us32_n750, us32_n751, us32_n752, us32_n753, us32_n754, us32_n755, 
       us32_n756, us32_n757, us32_n758, us32_n759, us32_n760, us32_n761, us32_n762, us32_n763, us32_n764, 
       us32_n765, us32_n766, us32_n767, us32_n768, us32_n769, us32_n770, us32_n771, us32_n772, us32_n773, 
       us32_n774, us32_n775, us32_n776, us32_n777, us32_n778, us32_n779, us32_n780, us32_n781, us32_n782, 
       us32_n783, us32_n784, us32_n785, us32_n786, us32_n787, us32_n788, us32_n789, us32_n790, us32_n791, 
       us32_n792, us32_n793, us32_n794, us32_n795, us32_n796, us32_n797, us32_n798, us32_n799, us32_n800, 
       us32_n801, us32_n802, us32_n803, us32_n804, us32_n805, us32_n806, us32_n807, us32_n808, us32_n809, 
       us32_n810, us32_n811, us32_n812, us32_n813, us32_n814, us32_n815, us32_n816, us32_n817, us32_n818, 
       us32_n819, us32_n820, us32_n821, us32_n822, us32_n823, us32_n824, us32_n825, us32_n826, us32_n827, 
       us32_n828, us32_n829, us32_n830, us32_n831, us32_n832, us32_n833, us32_n834, us32_n835, us32_n836, 
       us32_n837, us32_n838, us32_n839, us32_n840, us32_n841, us32_n842, us32_n843, us32_n844, us32_n845, 
       us32_n846, us32_n847, us32_n848, us32_n849, us32_n850, us32_n851, us32_n852, us32_n853, us32_n854, 
       us32_n855, us32_n856, us32_n857, us32_n858, us32_n859, us32_n860, us32_n861, us32_n862, us32_n863, 
       us32_n864, us32_n865, us32_n866, us32_n867, us32_n868, us32_n869, us32_n870, us32_n871, us32_n872, 
       us32_n873, us32_n874, us32_n875,  us32_n876;
  NOR2_X1 u0_u1_U10 (.ZN( u0_u1_n709 ) , .A2( u0_u1_n778 ) , .A1( u0_u1_n802 ) );
  INV_X1 u0_u1_U100 (.A( u0_u1_n819 ) , .ZN( u0_u1_n845 ) );
  INV_X1 u0_u1_U101 (.A( u0_u1_n674 ) , .ZN( u0_u1_n860 ) );
  AOI21_X1 u0_u1_U102 (.A( u0_u1_n672 ) , .B1( u0_u1_n673 ) , .ZN( u0_u1_n674 ) , .B2( u0_u1_n857 ) );
  INV_X1 u0_u1_U103 (.A( u0_u1_n756 ) , .ZN( u0_u1_n870 ) );
  OAI21_X1 u0_u1_U104 (.B1( u0_u1_n755 ) , .ZN( u0_u1_n756 ) , .A( u0_u1_n846 ) , .B2( u0_u1_n869 ) );
  AOI221_X1 u0_u1_U105 (.A( u0_u1_n715 ) , .B2( u0_u1_n716 ) , .ZN( u0_u1_n722 ) , .C1( u0_u1_n834 ) , .B1( u0_u1_n840 ) , .C2( u0_u1_n864 ) );
  OR2_X1 u0_u1_U106 (.A2( u0_u1_n713 ) , .A1( u0_u1_n714 ) , .ZN( u0_u1_n715 ) );
  NAND2_X1 u0_u1_U107 (.A1( u0_u1_n449 ) , .A2( u0_u1_n451 ) , .ZN( u0_u1_n807 ) );
  NOR3_X1 u0_u1_U108 (.ZN( u0_u1_n754 ) , .A2( u0_u1_n854 ) , .A1( u0_u1_n864 ) , .A3( u0_u1_n866 ) );
  NOR2_X1 u0_u1_U109 (.ZN( u0_u1_n753 ) , .A2( u0_u1_n853 ) , .A1( u0_u1_n861 ) );
  NOR2_X1 u0_u1_U11 (.A1( u0_u1_n680 ) , .ZN( u0_u1_n695 ) , .A2( u0_u1_n809 ) );
  INV_X1 u0_u1_U110 (.A( u0_u1_n440 ) , .ZN( u0_u1_n815 ) );
  NAND2_X1 u0_u1_U111 (.A1( u0_u1_n449 ) , .A2( u0_u1_n467 ) , .ZN( u0_u1_n751 ) );
  AOI211_X1 u0_u1_U112 (.B( u0_u1_n809 ) , .A( u0_u1_n810 ) , .ZN( u0_u1_n826 ) , .C1( u0_u1_n843 ) , .C2( u0_u1_n851 ) );
  NOR2_X1 u0_u1_U113 (.ZN( u0_u1_n509 ) , .A1( u0_u1_n814 ) , .A2( u0_u1_n819 ) );
  OAI22_X1 u0_u1_U114 (.B1( u0_u1_n492 ) , .ZN( u0_u1_n493 ) , .A1( u0_u1_n688 ) , .A2( u0_u1_n765 ) , .B2( u0_u1_n819 ) );
  NOR3_X1 u0_u1_U115 (.ZN( u0_u1_n492 ) , .A1( u0_u1_n784 ) , .A2( u0_u1_n851 ) , .A3( u0_u1_n864 ) );
  NOR2_X1 u0_u1_U116 (.ZN( u0_u1_n579 ) , .A2( u0_u1_n701 ) , .A1( u0_u1_n816 ) );
  NOR2_X1 u0_u1_U117 (.ZN( u0_u1_n548 ) , .A2( u0_u1_n782 ) , .A1( u0_u1_n816 ) );
  NOR2_X1 u0_u1_U118 (.ZN( u0_u1_n508 ) , .A2( u0_u1_n730 ) , .A1( u0_u1_n764 ) );
  INV_X1 u0_u1_U119 (.A( u0_u1_n814 ) , .ZN( u0_u1_n855 ) );
  INV_X1 u0_u1_U12 (.A( u0_u1_n609 ) , .ZN( u0_u1_n875 ) );
  NOR2_X1 u0_u1_U120 (.ZN( u0_u1_n534 ) , .A2( u0_u1_n751 ) , .A1( u0_u1_n752 ) );
  NOR2_X1 u0_u1_U121 (.ZN( u0_u1_n603 ) , .A2( u0_u1_n782 ) , .A1( u0_u1_n805 ) );
  NOR2_X1 u0_u1_U122 (.ZN( u0_u1_n530 ) , .A2( u0_u1_n726 ) , .A1( u0_u1_n805 ) );
  INV_X1 u0_u1_U123 (.A( u0_u1_n816 ) , .ZN( u0_u1_n835 ) );
  AOI21_X1 u0_u1_U124 (.B1( u0_u1_n701 ) , .ZN( u0_u1_n702 ) , .A( u0_u1_n734 ) , .B2( u0_u1_n765 ) );
  NOR2_X1 u0_u1_U125 (.ZN( u0_u1_n557 ) , .A1( u0_u1_n752 ) , .A2( u0_u1_n793 ) );
  NOR2_X1 u0_u1_U126 (.ZN( u0_u1_n668 ) , .A1( u0_u1_n730 ) , .A2( u0_u1_n805 ) );
  NOR2_X1 u0_u1_U127 (.ZN( u0_u1_n547 ) , .A1( u0_u1_n751 ) , .A2( u0_u1_n816 ) );
  NOR2_X1 u0_u1_U128 (.ZN( u0_u1_n511 ) , .A1( u0_u1_n731 ) , .A2( u0_u1_n781 ) );
  NOR2_X1 u0_u1_U129 (.A1( u0_u1_n751 ) , .ZN( u0_u1_n769 ) , .A2( u0_u1_n805 ) );
  INV_X1 u0_u1_U13 (.A( u0_u1_n649 ) , .ZN( u0_u1_n871 ) );
  NOR2_X1 u0_u1_U130 (.ZN( u0_u1_n654 ) , .A1( u0_u1_n671 ) , .A2( u0_u1_n816 ) );
  NOR2_X1 u0_u1_U131 (.ZN( u0_u1_n604 ) , .A1( u0_u1_n671 ) , .A2( u0_u1_n805 ) );
  NOR2_X1 u0_u1_U132 (.ZN( u0_u1_n658 ) , .A1( u0_u1_n749 ) , .A2( u0_u1_n782 ) );
  NOR2_X1 u0_u1_U133 (.ZN( u0_u1_n529 ) , .A1( u0_u1_n671 ) , .A2( u0_u1_n781 ) );
  INV_X1 u0_u1_U134 (.A( u0_u1_n701 ) , .ZN( u0_u1_n854 ) );
  NOR2_X1 u0_u1_U135 (.ZN( u0_u1_n611 ) , .A2( u0_u1_n726 ) , .A1( u0_u1_n819 ) );
  AOI21_X1 u0_u1_U136 (.ZN( u0_u1_n571 ) , .B1( u0_u1_n752 ) , .B2( u0_u1_n764 ) , .A( u0_u1_n782 ) );
  AOI21_X1 u0_u1_U137 (.ZN( u0_u1_n500 ) , .A( u0_u1_n726 ) , .B2( u0_u1_n764 ) , .B1( u0_u1_n816 ) );
  NOR2_X1 u0_u1_U138 (.ZN( u0_u1_n685 ) , .A2( u0_u1_n701 ) , .A1( u0_u1_n805 ) );
  NOR2_X1 u0_u1_U139 (.ZN( u0_u1_n713 ) , .A1( u0_u1_n764 ) , .A2( u0_u1_n765 ) );
  NOR4_X1 u0_u1_U14 (.ZN( u0_u1_n458 ) , .A2( u0_u1_n519 ) , .A1( u0_u1_n545 ) , .A3( u0_u1_n581 ) , .A4( u0_u1_n617 ) );
  INV_X1 u0_u1_U140 (.A( u0_u1_n805 ) , .ZN( u0_u1_n844 ) );
  AOI21_X1 u0_u1_U141 (.ZN( u0_u1_n517 ) , .A( u0_u1_n731 ) , .B1( u0_u1_n752 ) , .B2( u0_u1_n805 ) );
  AOI21_X1 u0_u1_U142 (.B1( u0_u1_n627 ) , .ZN( u0_u1_n629 ) , .A( u0_u1_n765 ) , .B2( u0_u1_n816 ) );
  INV_X1 u0_u1_U143 (.A( u0_u1_n792 ) , .ZN( u0_u1_n834 ) );
  NOR2_X1 u0_u1_U144 (.ZN( u0_u1_n616 ) , .A1( u0_u1_n764 ) , .A2( u0_u1_n814 ) );
  NOR2_X1 u0_u1_U145 (.ZN( u0_u1_n561 ) , .A2( u0_u1_n793 ) , .A1( u0_u1_n805 ) );
  NAND2_X1 u0_u1_U146 (.A1( u0_u1_n701 ) , .A2( u0_u1_n731 ) , .ZN( u0_u1_n784 ) );
  INV_X1 u0_u1_U147 (.A( u0_u1_n749 ) , .ZN( u0_u1_n836 ) );
  INV_X1 u0_u1_U148 (.A( u0_u1_n752 ) , .ZN( u0_u1_n843 ) );
  NOR2_X1 u0_u1_U149 (.ZN( u0_u1_n570 ) , .A1( u0_u1_n731 ) , .A2( u0_u1_n764 ) );
  NOR4_X1 u0_u1_U15 (.ZN( u0_u1_n487 ) , .A2( u0_u1_n535 ) , .A1( u0_u1_n560 ) , .A3( u0_u1_n633 ) , .A4( u0_u1_n720 ) );
  INV_X1 u0_u1_U150 (.A( u0_u1_n730 ) , .ZN( u0_u1_n853 ) );
  AOI21_X1 u0_u1_U151 (.ZN( u0_u1_n566 ) , .B1( u0_u1_n726 ) , .A( u0_u1_n781 ) , .B2( u0_u1_n793 ) );
  AOI21_X1 u0_u1_U152 (.B1( u0_u1_n688 ) , .ZN( u0_u1_n689 ) , .A( u0_u1_n730 ) , .B2( u0_u1_n763 ) );
  INV_X1 u0_u1_U153 (.A( u0_u1_n731 ) , .ZN( u0_u1_n869 ) );
  AOI211_X1 u0_u1_U154 (.C2( u0_u1_n440 ) , .B( u0_u1_n625 ) , .A( u0_u1_n626 ) , .ZN( u0_u1_n637 ) , .C1( u0_u1_n864 ) );
  NOR4_X1 u0_u1_U155 (.A4( u0_u1_n631 ) , .A3( u0_u1_n632 ) , .A2( u0_u1_n633 ) , .A1( u0_u1_n634 ) , .ZN( u0_u1_n635 ) );
  NOR4_X1 u0_u1_U156 (.A4( u0_u1_n628 ) , .A3( u0_u1_n629 ) , .A2( u0_u1_n630 ) , .ZN( u0_u1_n636 ) , .A1( u0_u1_n666 ) );
  AOI21_X1 u0_u1_U157 (.ZN( u0_u1_n542 ) , .A( u0_u1_n765 ) , .B2( u0_u1_n781 ) , .B1( u0_u1_n819 ) );
  OAI21_X1 u0_u1_U158 (.A( u0_u1_n700 ) , .ZN( u0_u1_n704 ) , .B2( u0_u1_n752 ) , .B1( u0_u1_n806 ) );
  OAI21_X1 u0_u1_U159 (.ZN( u0_u1_n700 ) , .B2( u0_u1_n835 ) , .B1( u0_u1_n839 ) , .A( u0_u1_n861 ) );
  NOR4_X1 u0_u1_U16 (.A4( u0_u1_n447 ) , .A3( u0_u1_n448 ) , .A2( u0_u1_n518 ) , .A1( u0_u1_n543 ) , .ZN( u0_u1_n708 ) );
  INV_X1 u0_u1_U160 (.A( u0_u1_n765 ) , .ZN( u0_u1_n867 ) );
  NOR2_X1 u0_u1_U161 (.ZN( u0_u1_n528 ) , .A1( u0_u1_n726 ) , .A2( u0_u1_n752 ) );
  AOI21_X1 u0_u1_U162 (.ZN( u0_u1_n445 ) , .B1( u0_u1_n791 ) , .B2( u0_u1_n793 ) , .A( u0_u1_n816 ) );
  NAND4_X1 u0_u1_U163 (.A4( u0_u1_n495 ) , .A3( u0_u1_n496 ) , .A1( u0_u1_n497 ) , .ZN( u0_u1_n804 ) , .A2( u0_u1_n868 ) );
  AOI221_X1 u0_u1_U164 (.B2( u0_u1_n440 ) , .A( u0_u1_n491 ) , .ZN( u0_u1_n496 ) , .C2( u0_u1_n842 ) , .C1( u0_u1_n852 ) , .B1( u0_u1_n861 ) );
  NOR4_X1 u0_u1_U165 (.A3( u0_u1_n439 ) , .A2( u0_u1_n493 ) , .A1( u0_u1_n494 ) , .ZN( u0_u1_n495 ) , .A4( u0_u1_n614 ) );
  INV_X1 u0_u1_U166 (.A( u0_u1_n780 ) , .ZN( u0_u1_n868 ) );
  AOI21_X1 u0_u1_U167 (.ZN( u0_u1_n499 ) , .A( u0_u1_n781 ) , .B2( u0_u1_n793 ) , .B1( u0_u1_n806 ) );
  INV_X1 u0_u1_U168 (.A( u0_u1_n782 ) , .ZN( u0_u1_n851 ) );
  NAND2_X1 u0_u1_U169 (.ZN( u0_u1_n716 ) , .A1( u0_u1_n730 ) , .A2( u0_u1_n782 ) );
  OR3_X1 u0_u1_U17 (.ZN( u0_u1_n448 ) , .A1( u0_u1_n530 ) , .A3( u0_u1_n579 ) , .A2( u0_u1_n876 ) );
  BUF_X2 u0_u1_U170 (.Z( u0_u1_n41 ) , .A( u0_u1_n699 ) );
  OR4_X1 u0_u1_U171 (.A4( u0_u1_n582 ) , .A3( u0_u1_n583 ) , .A2( u0_u1_n584 ) , .A1( u0_u1_n585 ) , .ZN( u0_u1_n586 ) );
  INV_X1 u0_u1_U172 (.A( u0_u1_n726 ) , .ZN( u0_u1_n857 ) );
  OAI222_X1 u0_u1_U173 (.B2( u0_u1_n710 ) , .ZN( u0_u1_n711 ) , .C2( u0_u1_n726 ) , .B1( u0_u1_n749 ) , .A1( u0_u1_n808 ) , .C1( u0_u1_n816 ) , .A2( u0_u1_n817 ) );
  AOI221_X1 u0_u1_U174 (.A( u0_u1_n766 ) , .ZN( u0_u1_n776 ) , .C2( u0_u1_n812 ) , .B2( u0_u1_n837 ) , .C1( u0_u1_n856 ) , .B1( u0_u1_n867 ) );
  INV_X1 u0_u1_U175 (.A( u0_u1_n763 ) , .ZN( u0_u1_n837 ) );
  OAI221_X1 u0_u1_U176 (.A( u0_u1_n729 ) , .C2( u0_u1_n730 ) , .B2( u0_u1_n731 ) , .B1( u0_u1_n732 ) , .ZN( u0_u1_n739 ) , .C1( u0_u1_n819 ) );
  OAI221_X1 u0_u1_U177 (.C2( u0_u1_n441 ) , .A( u0_u1_n785 ) , .B2( u0_u1_n787 ) , .B1( u0_u1_n788 ) , .ZN( u0_u1_n798 ) , .C1( u0_u1_n815 ) );
  AOI22_X1 u0_u1_U178 (.A2( u0_u1_n784 ) , .ZN( u0_u1_n785 ) , .B2( u0_u1_n833 ) , .A1( u0_u1_n836 ) , .B1( u0_u1_n864 ) );
  OAI221_X1 u0_u1_U179 (.C2( u0_u1_n441 ) , .A( u0_u1_n698 ) , .ZN( u0_u1_n705 ) , .C1( u0_u1_n787 ) , .B1( u0_u1_n788 ) , .B2( u0_u1_n808 ) );
  OR4_X1 u0_u1_U18 (.A4( u0_u1_n444 ) , .A2( u0_u1_n445 ) , .A1( u0_u1_n446 ) , .ZN( u0_u1_n447 ) , .A3( u0_u1_n555 ) );
  AOI22_X1 u0_u1_U180 (.ZN( u0_u1_n698 ) , .A1( u0_u1_n832 ) , .B2( u0_u1_n844 ) , .A2( u0_u1_n866 ) , .B1( u0_u1_n869 ) );
  OAI222_X1 u0_u1_U181 (.B1( u0_u1_n41 ) , .ZN( u0_u1_n619 ) , .C1( u0_u1_n726 ) , .C2( u0_u1_n749 ) , .B2( u0_u1_n788 ) , .A2( u0_u1_n794 ) , .A1( u0_u1_n818 ) );
  NAND2_X1 u0_u1_U182 (.A2( u0_u1_n450 ) , .A1( u0_u1_n466 ) , .ZN( u0_u1_n817 ) );
  NAND2_X1 u0_u1_U183 (.A2( u0_u1_n456 ) , .A1( u0_u1_n474 ) , .ZN( u0_u1_n781 ) );
  NAND2_X1 u0_u1_U184 (.A2( u0_u1_n450 ) , .A1( u0_u1_n454 ) , .ZN( u0_u1_n731 ) );
  NAND2_X1 u0_u1_U185 (.A1( u0_u1_n455 ) , .A2( u0_u1_n474 ) , .ZN( u0_u1_n787 ) );
  NAND2_X1 u0_u1_U186 (.A1( u0_u1_n455 ) , .A2( u0_u1_n463 ) , .ZN( u0_u1_n746 ) );
  NAND2_X1 u0_u1_U187 (.A1( u0_u1_n453 ) , .A2( u0_u1_n473 ) , .ZN( u0_u1_n818 ) );
  NAND2_X1 u0_u1_U188 (.A2( u0_u1_n455 ) , .A1( u0_u1_n457 ) , .ZN( u0_u1_n808 ) );
  NOR2_X1 u0_u1_U189 (.ZN( u0_u1_n467 ) , .A2( u0_u1_n848 ) , .A1( u0_u1_n849 ) );
  INV_X1 u0_u1_U19 (.A( u0_u1_n615 ) , .ZN( u0_u1_n876 ) );
  NAND2_X1 u0_u1_U190 (.A1( u0_u1_n449 ) , .A2( u0_u1_n450 ) , .ZN( u0_u1_n788 ) );
  NAND2_X1 u0_u1_U191 (.A2( u0_u1_n463 ) , .A1( u0_u1_n464 ) , .ZN( u0_u1_n749 ) );
  NAND2_X1 u0_u1_U192 (.A1( u0_u1_n464 ) , .A2( u0_u1_n474 ) , .ZN( u0_u1_n790 ) );
  NAND2_X1 u0_u1_U193 (.A1( u0_u1_n453 ) , .A2( u0_u1_n464 ) , .ZN( u0_u1_n792 ) );
  AND2_X1 u0_u1_U194 (.ZN( u0_u1_n440 ) , .A1( u0_u1_n456 ) , .A2( u0_u1_n463 ) );
  NOR2_X1 u0_u1_U195 (.A2( u0_n268 ) , .ZN( u0_u1_n462 ) , .A1( u0_u1_n850 ) );
  AOI222_X1 u0_u1_U196 (.B2( u0_u1_n640 ) , .ZN( u0_u1_n646 ) , .B1( u0_u1_n842 ) , .A1( u0_u1_n843 ) , .C2( u0_u1_n847 ) , .C1( u0_u1_n864 ) , .A2( u0_u1_n866 ) );
  NOR4_X1 u0_u1_U197 (.A4( u0_u1_n641 ) , .A3( u0_u1_n642 ) , .A2( u0_u1_n643 ) , .A1( u0_u1_n644 ) , .ZN( u0_u1_n645 ) );
  NOR4_X1 u0_u1_U198 (.A4( u0_u1_n500 ) , .A3( u0_u1_n501 ) , .A2( u0_u1_n502 ) , .ZN( u0_u1_n503 ) , .A1( u0_u1_n529 ) );
  AOI221_X1 u0_u1_U199 (.A( u0_u1_n499 ) , .ZN( u0_u1_n504 ) , .B2( u0_u1_n844 ) , .C1( u0_u1_n847 ) , .C2( u0_u1_n861 ) , .B1( u0_u1_n863 ) );
  NOR4_X1 u0_u1_U20 (.ZN( u0_u1_n622 ) , .A1( u0_u1_n658 ) , .A3( u0_u1_n668 ) , .A4( u0_u1_n684 ) , .A2( u0_u1_n768 ) );
  AOI221_X1 u0_u1_U200 (.A( u0_u1_n783 ) , .ZN( u0_u1_n800 ) , .C2( u0_u1_n838 ) , .B2( u0_u1_n839 ) , .B1( u0_u1_n866 ) , .C1( u0_u1_n867 ) );
  NOR4_X1 u0_u1_U201 (.A4( u0_u1_n795 ) , .A3( u0_u1_n796 ) , .A2( u0_u1_n797 ) , .A1( u0_u1_n798 ) , .ZN( u0_u1_n799 ) );
  NAND4_X1 u0_u1_U202 (.ZN( u0_subword_23 ) , .A4( u0_u1_n824 ) , .A3( u0_u1_n825 ) , .A2( u0_u1_n826 ) , .A1( u0_u1_n827 ) );
  NOR4_X1 u0_u1_U203 (.A4( u0_u1_n820 ) , .A3( u0_u1_n821 ) , .A2( u0_u1_n822 ) , .A1( u0_u1_n823 ) , .ZN( u0_u1_n824 ) );
  NOR4_X1 u0_u1_U204 (.A4( u0_u1_n736 ) , .A3( u0_u1_n737 ) , .A2( u0_u1_n738 ) , .A1( u0_u1_n739 ) , .ZN( u0_u1_n740 ) );
  NOR4_X1 u0_u1_U205 (.A3( u0_u1_n757 ) , .A2( u0_u1_n758 ) , .A1( u0_u1_n759 ) , .ZN( u0_u1_n760 ) , .A4( u0_u1_n870 ) );
  AOI211_X1 u0_u1_U206 (.B( u0_u1_n747 ) , .A( u0_u1_n748 ) , .ZN( u0_u1_n761 ) , .C1( u0_u1_n834 ) , .C2( u0_u1_n854 ) );
  NOR4_X1 u0_u1_U207 (.A4( u0_u1_n702 ) , .A3( u0_u1_n703 ) , .A2( u0_u1_n704 ) , .A1( u0_u1_n705 ) , .ZN( u0_u1_n706 ) );
  AOI211_X1 u0_u1_U208 (.B( u0_u1_n696 ) , .A( u0_u1_n697 ) , .ZN( u0_u1_n707 ) , .C2( u0_u1_n833 ) , .C1( u0_u1_n852 ) );
  NAND4_X1 u0_u1_U209 (.ZN( u0_subword_17 ) , .A4( u0_u1_n597 ) , .A3( u0_u1_n598 ) , .A2( u0_u1_n599 ) , .A1( u0_u1_n600 ) );
  NOR4_X1 u0_u1_U21 (.A4( u0_u1_n611 ) , .A3( u0_u1_n612 ) , .A2( u0_u1_n613 ) , .A1( u0_u1_n614 ) , .ZN( u0_u1_n621 ) );
  NOR4_X1 u0_u1_U210 (.A4( u0_u1_n593 ) , .A3( u0_u1_n594 ) , .A2( u0_u1_n595 ) , .A1( u0_u1_n596 ) , .ZN( u0_u1_n597 ) );
  AOI211_X1 u0_u1_U211 (.B( u0_u1_n591 ) , .A( u0_u1_n592 ) , .ZN( u0_u1_n598 ) , .C2( u0_u1_n813 ) , .C1( u0_u1_n835 ) );
  NAND2_X1 u0_u1_U212 (.A2( u0_u1_n443 ) , .A1( u0_u1_n454 ) , .ZN( u0_u1_n793 ) );
  AOI21_X1 u0_u1_U213 (.ZN( u0_u1_n642 ) , .B2( u0_u1_n749 ) , .A( u0_u1_n794 ) , .B1( u0_u1_n805 ) );
  AOI21_X1 u0_u1_U214 (.ZN( u0_u1_n516 ) , .A( u0_u1_n781 ) , .B2( u0_u1_n794 ) , .B1( u0_u1_n814 ) );
  INV_X1 u0_u1_U215 (.A( u0_u1_n794 ) , .ZN( u0_u1_n852 ) );
  NOR2_X1 u0_u1_U216 (.ZN( u0_u1_n559 ) , .A1( u0_u1_n794 ) , .A2( u0_u1_n816 ) );
  NOR2_X1 u0_u1_U217 (.ZN( u0_u1_n585 ) , .A1( u0_u1_n794 ) , .A2( u0_u1_n819 ) );
  NAND2_X2 u0_u1_U218 (.A1( u0_u1_n453 ) , .A2( u0_u1_n455 ) , .ZN( u0_u1_n764 ) );
  NAND2_X2 u0_u1_U219 (.A1( u0_u1_n453 ) , .A2( u0_u1_n456 ) , .ZN( u0_u1_n816 ) );
  NOR4_X1 u0_u1_U22 (.ZN( u0_u1_n563 ) , .A1( u0_u1_n655 ) , .A3( u0_u1_n663 ) , .A4( u0_u1_n687 ) , .A2( u0_u1_n770 ) );
  NOR2_X1 u0_u1_U220 (.ZN( u0_u1_n453 ) , .A1( u0_u1_n830 ) , .A2( u0_u1_n831 ) );
  NAND2_X1 u0_u1_U221 (.A1( u0_u1_n454 ) , .A2( u0_u1_n467 ) , .ZN( u0_u1_n671 ) );
  NAND2_X1 u0_u1_U222 (.A1( u0_u1_n443 ) , .A2( u0_u1_n462 ) , .ZN( u0_u1_n701 ) );
  NOR2_X1 u0_u1_U223 (.ZN( u0_u1_n455 ) , .A1( u0_u1_n828 ) , .A2( u0_u1_n829 ) );
  AOI211_X1 u0_u1_U224 (.B( u0_u1_n727 ) , .A( u0_u1_n728 ) , .ZN( u0_u1_n741 ) , .C1( u0_u1_n844 ) , .C2( u0_u1_n856 ) );
  NOR2_X1 u0_u1_U225 (.A2( u0_u1_n710 ) , .A1( u0_u1_n764 ) , .ZN( u0_u1_n796 ) );
  NOR2_X1 u0_u1_U226 (.ZN( u0_u1_n519 ) , .A1( u0_u1_n710 ) , .A2( u0_u1_n805 ) );
  NOR2_X1 u0_u1_U227 (.ZN( u0_u1_n684 ) , .A2( u0_u1_n710 ) , .A1( u0_u1_n819 ) );
  NOR2_X1 u0_u1_U228 (.A2( u0_u1_n710 ) , .A1( u0_u1_n752 ) , .ZN( u0_u1_n773 ) );
  NOR2_X1 u0_u1_U229 (.ZN( u0_u1_n522 ) , .A2( u0_u1_n710 ) , .A1( u0_u1_n816 ) );
  NOR4_X1 u0_u1_U23 (.ZN( u0_u1_n477 ) , .A1( u0_u1_n533 ) , .A3( u0_u1_n570 ) , .A4( u0_u1_n602 ) , .A2( u0_u1_n644 ) );
  NOR2_X1 u0_u1_U230 (.ZN( u0_u1_n531 ) , .A1( u0_u1_n710 ) , .A2( u0_u1_n781 ) );
  INV_X1 u0_u1_U231 (.A( u0_u1_n682 ) , .ZN( u0_u1_n841 ) );
  AOI21_X1 u0_u1_U232 (.ZN( u0_u1_n643 ) , .B1( u0_u1_n682 ) , .A( u0_u1_n793 ) , .B2( u0_u1_n819 ) );
  OAI22_X1 u0_u1_U233 (.B2( u0_u1_n781 ) , .B1( u0_u1_n782 ) , .ZN( u0_u1_n783 ) , .A2( u0_u1_n816 ) , .A1( u0_u1_n817 ) );
  AOI21_X1 u0_u1_U234 (.ZN( u0_u1_n591 ) , .B2( u0_u1_n701 ) , .B1( u0_u1_n817 ) , .A( u0_u1_n819 ) );
  INV_X1 u0_u1_U235 (.A( u0_u1_n817 ) , .ZN( u0_u1_n856 ) );
  NOR2_X1 u0_u1_U236 (.ZN( u0_u1_n669 ) , .A1( u0_u1_n752 ) , .A2( u0_u1_n817 ) );
  AOI21_X1 u0_u1_U237 (.ZN( u0_u1_n541 ) , .B2( u0_u1_n814 ) , .A( u0_u1_n816 ) , .B1( u0_u1_n817 ) );
  AOI21_X1 u0_u1_U238 (.ZN( u0_u1_n452 ) , .B2( u0_u1_n794 ) , .A( u0_u1_n805 ) , .B1( u0_u1_n817 ) );
  NOR2_X1 u0_u1_U239 (.ZN( u0_u1_n472 ) , .A2( u0_u1_n781 ) , .A1( u0_u1_n817 ) );
  NOR4_X1 u0_u1_U24 (.ZN( u0_u1_n483 ) , .A3( u0_u1_n534 ) , .A4( u0_u1_n547 ) , .A2( u0_u1_n569 ) , .A1( u0_u1_n719 ) );
  OAI222_X1 u0_u1_U240 (.A2( u0_u1_n671 ) , .ZN( u0_u1_n676 ) , .B1( u0_u1_n749 ) , .B2( u0_u1_n786 ) , .C2( u0_u1_n790 ) , .C1( u0_u1_n817 ) , .A1( u0_u1_n819 ) );
  NOR2_X1 u0_u1_U241 (.ZN( u0_u1_n632 ) , .A1( u0_u1_n749 ) , .A2( u0_u1_n817 ) );
  NAND2_X1 u0_u1_U242 (.A1( u0_u1_n443 ) , .A2( u0_u1_n466 ) , .ZN( u0_u1_n710 ) );
  NAND2_X1 u0_u1_U243 (.A2( u0_u1_n463 ) , .A1( u0_u1_n473 ) , .ZN( u0_u1_n699 ) );
  INV_X1 u0_u1_U244 (.ZN( u0_u1_n438 ) , .A( u0_u1_n788 ) );
  INV_X1 u0_u1_U245 (.ZN( u0_u1_n828 ) , .A( w3_8 ) );
  NOR2_X1 u0_u1_U246 (.ZN( u0_u1_n456 ) , .A1( u0_u1_n829 ) , .A2( w3_8 ) );
  NOR2_X1 u0_u1_U247 (.A2( u0_n270 ) , .ZN( u0_u1_n454 ) , .A1( u0_u1_n859 ) );
  OAI21_X1 u0_u1_U248 (.A( u0_u1_n789 ) , .B2( u0_u1_n790 ) , .B1( u0_u1_n791 ) , .ZN( u0_u1_n797 ) );
  AOI21_X1 u0_u1_U249 (.ZN( u0_u1_n641 ) , .B2( u0_u1_n751 ) , .A( u0_u1_n790 ) , .B1( u0_u1_n814 ) );
  INV_X1 u0_u1_U25 (.A( u0_u1_n751 ) , .ZN( u0_u1_n864 ) );
  AOI21_X1 u0_u1_U250 (.A( u0_u1_n735 ) , .ZN( u0_u1_n736 ) , .B2( u0_u1_n782 ) , .B1( u0_u1_n794 ) );
  AOI21_X1 u0_u1_U251 (.B2( u0_u1_n765 ) , .ZN( u0_u1_n766 ) , .A( u0_u1_n790 ) , .B1( u0_u1_n794 ) );
  AOI21_X1 u0_u1_U252 (.ZN( u0_u1_n444 ) , .A( u0_u1_n701 ) , .B1( u0_u1_n735 ) , .B2( u0_u1_n752 ) );
  NOR2_X1 u0_u1_U253 (.ZN( u0_u1_n520 ) , .A1( u0_u1_n710 ) , .A2( u0_u1_n790 ) );
  NOR2_X1 u0_u1_U254 (.ZN( u0_u1_n536 ) , .A1( u0_u1_n726 ) , .A2( u0_u1_n790 ) );
  NOR2_X1 u0_u1_U255 (.ZN( u0_u1_n644 ) , .A2( u0_u1_n790 ) , .A1( u0_u1_n793 ) );
  NOR2_X1 u0_u1_U256 (.ZN( u0_u1_n583 ) , .A1( u0_u1_n671 ) , .A2( u0_u1_n790 ) );
  INV_X1 u0_u1_U257 (.A( u0_u1_n790 ) , .ZN( u0_u1_n846 ) );
  AOI222_X1 u0_u1_U258 (.ZN( u0_u1_n527 ) , .A1( u0_u1_n836 ) , .B2( u0_u1_n838 ) , .C1( u0_u1_n845 ) , .C2( u0_u1_n851 ) , .A2( u0_u1_n853 ) , .B1( u0_u1_n867 ) );
  NOR3_X1 u0_u1_U259 (.A2( u0_u1_n440 ) , .ZN( u0_u1_n442 ) , .A3( u0_u1_n838 ) , .A1( u0_u1_n847 ) );
  NOR4_X1 u0_u1_U26 (.A1( u0_u1_n533 ) , .ZN( u0_u1_n538 ) , .A2( u0_u1_n656 ) , .A4( u0_u1_n670 ) , .A3( u0_u1_n767 ) );
  NAND2_X1 u0_u1_U260 (.ZN( u0_u1_n615 ) , .A2( u0_u1_n838 ) , .A1( u0_u1_n874 ) );
  AND2_X1 u0_u1_U261 (.ZN( u0_u1_n627 ) , .A1( u0_u1_n732 ) , .A2( u0_u1_n815 ) );
  NAND2_X1 u0_u1_U262 (.A2( u0_u1_n456 ) , .A1( u0_u1_n457 ) , .ZN( u0_u1_n732 ) );
  NOR2_X1 u0_u1_U263 (.A2( u0_u1_n41 ) , .ZN( u0_u1_n439 ) , .A1( u0_u1_n793 ) );
  AOI21_X1 u0_u1_U264 (.ZN( u0_u1_n593 ) , .B2( u0_u1_n765 ) , .A( u0_u1_n787 ) , .B1( u0_u1_n814 ) );
  AND2_X1 u0_u1_U265 (.ZN( u0_u1_n734 ) , .A1( u0_u1_n781 ) , .A2( u0_u1_n787 ) );
  NAND4_X1 u0_u1_U266 (.A4( u0_u1_n550 ) , .A3( u0_u1_n551 ) , .A2( u0_u1_n552 ) , .A1( u0_u1_n553 ) , .ZN( u0_u1_n747 ) );
  NOR2_X1 u0_u1_U267 (.ZN( u0_u1_n666 ) , .A1( u0_u1_n787 ) , .A2( u0_u1_n793 ) );
  NOR2_X1 u0_u1_U268 (.ZN( u0_u1_n665 ) , .A1( u0_u1_n731 ) , .A2( u0_u1_n787 ) );
  NOR2_X1 u0_u1_U269 (.ZN( u0_u1_n510 ) , .A2( u0_u1_n782 ) , .A1( u0_u1_n787 ) );
  NOR4_X1 u0_u1_U27 (.A4( u0_u1_n543 ) , .A3( u0_u1_n544 ) , .A2( u0_u1_n545 ) , .ZN( u0_u1_n552 ) , .A1( u0_u1_n690 ) );
  NOR2_X1 u0_u1_U270 (.ZN( u0_u1_n630 ) , .A2( u0_u1_n671 ) , .A1( u0_u1_n787 ) );
  NOR2_X1 u0_u1_U271 (.ZN( u0_u1_n617 ) , .A1( u0_u1_n787 ) , .A2( u0_u1_n817 ) );
  INV_X1 u0_u1_U272 (.A( u0_u1_n787 ) , .ZN( u0_u1_n847 ) );
  NOR2_X1 u0_u1_U273 (.ZN( u0_u1_n545 ) , .A2( u0_u1_n710 ) , .A1( u0_u1_n787 ) );
  NOR2_X1 u0_u1_U274 (.ZN( u0_u1_n546 ) , .A2( u0_u1_n787 ) , .A1( u0_u1_n794 ) );
  NAND2_X1 u0_u1_U275 (.A2( u0_u1_n473 ) , .A1( u0_u1_n474 ) , .ZN( u0_u1_n819 ) );
  AOI222_X1 u0_u1_U276 (.C2( u0_u1_n811 ) , .B2( u0_u1_n812 ) , .A2( u0_u1_n813 ) , .ZN( u0_u1_n825 ) , .C1( u0_u1_n834 ) , .A1( u0_u1_n840 ) , .B1( u0_u1_n854 ) );
  AOI22_X1 u0_u1_U277 (.ZN( u0_u1_n729 ) , .B1( u0_u1_n834 ) , .A2( u0_u1_n839 ) , .A1( u0_u1_n864 ) , .B2( u0_u1_n867 ) );
  AOI222_X1 u0_u1_U278 (.ZN( u0_u1_n471 ) , .B1( u0_u1_n834 ) , .A1( u0_u1_n840 ) , .C1( u0_u1_n843 ) , .C2( u0_u1_n852 ) , .A2( u0_u1_n856 ) , .B2( u0_u1_n866 ) );
  NOR2_X1 u0_u1_U279 (.ZN( u0_u1_n688 ) , .A1( u0_u1_n833 ) , .A2( u0_u1_n834 ) );
  NOR2_X1 u0_u1_U28 (.ZN( u0_u1_n544 ) , .A1( u0_u1_n764 ) , .A2( u0_u1_n793 ) );
  NOR2_X1 u0_u1_U280 (.ZN( u0_u1_n735 ) , .A2( u0_u1_n834 ) , .A1( u0_u1_n846 ) );
  NAND4_X1 u0_u1_U281 (.A4( u0_u1_n537 ) , .A3( u0_u1_n538 ) , .A2( u0_u1_n539 ) , .A1( u0_u1_n540 ) , .ZN( u0_u1_n624 ) );
  NAND2_X2 u0_u1_U282 (.A1( u0_u1_n451 ) , .A2( u0_u1_n462 ) , .ZN( u0_u1_n794 ) );
  NAND2_X1 u0_u1_U283 (.A2( u0_u1_n466 ) , .A1( u0_u1_n467 ) , .ZN( u0_u1_n814 ) );
  NOR2_X1 u0_u1_U284 (.ZN( u0_u1_n631 ) , .A2( u0_u1_n730 ) , .A1( u0_u1_n787 ) );
  NAND2_X2 u0_u1_U285 (.A2( u0_u1_n450 ) , .A1( u0_u1_n462 ) , .ZN( u0_u1_n730 ) );
  NOR2_X1 u0_u1_U286 (.A2( u0_n274 ) , .ZN( u0_u1_n451 ) , .A1( u0_u1_n849 ) );
  NOR2_X1 u0_u1_U287 (.A1( u0_n272 ) , .A2( u0_n274 ) , .ZN( u0_u1_n443 ) );
  OAI22_X1 u0_u1_U288 (.ZN( u0_u1_n697 ) , .A2( u0_u1_n732 ) , .A1( u0_u1_n782 ) , .B1( u0_u1_n793 ) , .B2( u0_u1_n819 ) );
  AOI21_X1 u0_u1_U289 (.ZN( u0_u1_n512 ) , .B2( u0_u1_n671 ) , .A( u0_u1_n732 ) , .B1( u0_u1_n817 ) );
  NAND4_X1 u0_u1_U29 (.A4( u0_u1_n605 ) , .A3( u0_u1_n606 ) , .A2( u0_u1_n607 ) , .A1( u0_u1_n608 ) , .ZN( u0_u1_n724 ) );
  OAI22_X1 u0_u1_U290 (.ZN( u0_u1_n491 ) , .A1( u0_u1_n726 ) , .B2( u0_u1_n730 ) , .B1( u0_u1_n732 ) , .A2( u0_u1_n781 ) );
  NOR2_X1 u0_u1_U291 (.ZN( u0_u1_n581 ) , .A2( u0_u1_n710 ) , .A1( u0_u1_n732 ) );
  NOR2_X1 u0_u1_U292 (.ZN( u0_u1_n535 ) , .A2( u0_u1_n726 ) , .A1( u0_u1_n732 ) );
  INV_X1 u0_u1_U293 (.A( u0_u1_n732 ) , .ZN( u0_u1_n840 ) );
  AOI211_X1 u0_u1_U294 (.A( u0_u1_n498 ) , .ZN( u0_u1_n505 ) , .B( u0_u1_n804 ) , .C2( u0_u1_n840 ) , .C1( u0_u1_n852 ) );
  OAI21_X1 u0_u1_U295 (.ZN( u0_u1_n789 ) , .A( u0_u1_n840 ) , .B1( u0_u1_n864 ) , .B2( u0_u1_n874 ) );
  AOI222_X1 u0_u1_U296 (.ZN( u0_u1_n662 ) , .A2( u0_u1_n840 ) , .B1( u0_u1_n842 ) , .C2( u0_u1_n846 ) , .A1( u0_u1_n861 ) , .C1( u0_u1_n864 ) , .B2( u0_u1_n871 ) );
  AOI211_X1 u0_u1_U297 (.B( u0_u1_n541 ) , .A( u0_u1_n542 ) , .ZN( u0_u1_n553 ) , .C2( u0_u1_n840 ) , .C1( u0_u1_n852 ) );
  NOR2_X1 u0_u1_U298 (.ZN( u0_u1_n682 ) , .A2( u0_u1_n836 ) , .A1( u0_u1_n840 ) );
  NAND4_X1 u0_u1_U299 (.ZN( u0_subword_16 ) , .A4( u0_u1_n503 ) , .A3( u0_u1_n504 ) , .A2( u0_u1_n505 ) , .A1( u0_u1_n506 ) );
  NAND2_X1 u0_u1_U3 (.A1( u0_u1_n451 ) , .A2( u0_u1_n466 ) , .ZN( u0_u1_n726 ) );
  NOR4_X1 u0_u1_U30 (.A3( u0_u1_n602 ) , .A2( u0_u1_n603 ) , .A1( u0_u1_n604 ) , .ZN( u0_u1_n605 ) , .A4( u0_u1_n657 ) );
  AOI21_X1 u0_u1_U300 (.A( u0_u1_n792 ) , .B2( u0_u1_n793 ) , .B1( u0_u1_n794 ) , .ZN( u0_u1_n795 ) );
  AOI21_X1 u0_u1_U301 (.ZN( u0_u1_n628 ) , .B2( u0_u1_n671 ) , .A( u0_u1_n792 ) , .B1( u0_u1_n793 ) );
  NOR2_X1 u0_u1_U302 (.ZN( u0_u1_n657 ) , .A1( u0_u1_n792 ) , .A2( u0_u1_n817 ) );
  NOR2_X1 u0_u1_U303 (.ZN( u0_u1_n714 ) , .A2( u0_u1_n726 ) , .A1( u0_u1_n792 ) );
  NOR2_X1 u0_u1_U304 (.ZN( u0_u1_n523 ) , .A1( u0_u1_n792 ) , .A2( u0_u1_n814 ) );
  NOR2_X1 u0_u1_U305 (.ZN( u0_u1_n663 ) , .A1( u0_u1_n731 ) , .A2( u0_u1_n792 ) );
  NOR2_X1 u0_u1_U306 (.ZN( u0_u1_n670 ) , .A2( u0_u1_n710 ) , .A1( u0_u1_n792 ) );
  NOR3_X1 u0_u1_U307 (.A3( u0_u1_n743 ) , .A2( u0_u1_n744 ) , .A1( u0_u1_n745 ) , .ZN( u0_u1_n762 ) );
  NAND2_X2 u0_u1_U308 (.A2( u0_u1_n451 ) , .A1( u0_u1_n454 ) , .ZN( u0_u1_n765 ) );
  OAI22_X1 u0_u1_U309 (.ZN( u0_u1_n639 ) , .A1( u0_u1_n701 ) , .B2( u0_u1_n730 ) , .A2( u0_u1_n764 ) , .B1( u0_u1_n818 ) );
  NOR3_X1 u0_u1_U31 (.A1( u0_u1_n601 ) , .ZN( u0_u1_n606 ) , .A3( u0_u1_n665 ) , .A2( u0_u1_n772 ) );
  AOI21_X1 u0_u1_U310 (.ZN( u0_u1_n501 ) , .B1( u0_u1_n682 ) , .A( u0_u1_n814 ) , .B2( u0_u1_n818 ) );
  OAI22_X1 u0_u1_U311 (.A1( u0_u1_n726 ) , .ZN( u0_u1_n728 ) , .B2( u0_u1_n752 ) , .B1( u0_u1_n814 ) , .A2( u0_u1_n818 ) );
  AOI21_X1 u0_u1_U312 (.A( u0_u1_n817 ) , .B2( u0_u1_n818 ) , .B1( u0_u1_n819 ) , .ZN( u0_u1_n820 ) );
  OAI22_X1 u0_u1_U313 (.ZN( u0_u1_n626 ) , .B1( u0_u1_n671 ) , .B2( u0_u1_n749 ) , .A1( u0_u1_n817 ) , .A2( u0_u1_n818 ) );
  NOR2_X1 u0_u1_U314 (.ZN( u0_u1_n601 ) , .A2( u0_u1_n793 ) , .A1( u0_u1_n818 ) );
  NOR2_X1 u0_u1_U315 (.ZN( u0_u1_n533 ) , .A2( u0_u1_n782 ) , .A1( u0_u1_n818 ) );
  NOR2_X1 u0_u1_U316 (.A1( u0_u1_n671 ) , .ZN( u0_u1_n690 ) , .A2( u0_u1_n818 ) );
  NOR2_X1 u0_u1_U317 (.ZN( u0_u1_n521 ) , .A2( u0_u1_n701 ) , .A1( u0_u1_n818 ) );
  NOR2_X1 u0_u1_U318 (.ZN( u0_u1_n560 ) , .A1( u0_u1_n710 ) , .A2( u0_u1_n818 ) );
  NOR2_X1 u0_u1_U319 (.ZN( u0_u1_n687 ) , .A1( u0_u1_n731 ) , .A2( u0_u1_n818 ) );
  NOR3_X1 u0_u1_U32 (.ZN( u0_u1_n551 ) , .A2( u0_u1_n653 ) , .A1( u0_u1_n669 ) , .A3( u0_u1_n773 ) );
  INV_X1 u0_u1_U320 (.A( u0_u1_n818 ) , .ZN( u0_u1_n833 ) );
  BUF_X2 u0_u1_U321 (.Z( u0_u1_n441 ) , .A( u0_u1_n786 ) );
  NAND2_X1 u0_u1_U322 (.A2( u0_u1_n443 ) , .A1( u0_u1_n449 ) , .ZN( u0_u1_n786 ) );
  AOI222_X1 u0_u1_U323 (.ZN( u0_u1_n777 ) , .A1( u0_u1_n832 ) , .C1( u0_u1_n836 ) , .B2( u0_u1_n842 ) , .A2( u0_u1_n851 ) , .B1( u0_u1_n862 ) , .C2( u0_u1_n874 ) );
  INV_X1 u0_u1_U324 (.A( u0_n268 ) , .ZN( u0_u1_n859 ) );
  INV_X1 u0_u1_U325 (.A( u0_n274 ) , .ZN( u0_u1_n848 ) );
  INV_X1 u0_u1_U326 (.A( u0_u1_n786 ) , .ZN( u0_u1_n862 ) );
  OAI22_X1 u0_u1_U327 (.B2( u0_u1_n752 ) , .B1( u0_u1_n753 ) , .A1( u0_u1_n754 ) , .ZN( u0_u1_n758 ) , .A2( u0_u1_n808 ) );
  OAI222_X1 u0_u1_U328 (.ZN( u0_u1_n507 ) , .C2( u0_u1_n627 ) , .B2( u0_u1_n649 ) , .B1( u0_u1_n749 ) , .A2( u0_u1_n750 ) , .C1( u0_u1_n807 ) , .A1( u0_u1_n808 ) );
  AOI21_X1 u0_u1_U329 (.ZN( u0_u1_n691 ) , .B2( u0_u1_n751 ) , .B1( u0_u1_n765 ) , .A( u0_u1_n808 ) );
  NOR4_X1 u0_u1_U33 (.A4( u0_u1_n546 ) , .A3( u0_u1_n547 ) , .A2( u0_u1_n548 ) , .A1( u0_u1_n549 ) , .ZN( u0_u1_n550 ) );
  NAND2_X1 u0_u1_U330 (.A2( u0_u1_n764 ) , .A1( u0_u1_n808 ) , .ZN( u0_u1_n812 ) );
  NOR2_X1 u0_u1_U331 (.ZN( u0_u1_n572 ) , .A1( u0_u1_n730 ) , .A2( u0_u1_n808 ) );
  AOI21_X1 u0_u1_U332 (.ZN( u0_u1_n479 ) , .A( u0_u1_n671 ) , .B1( u0_u1_n752 ) , .B2( u0_u1_n808 ) );
  OAI22_X1 u0_u1_U333 (.ZN( u0_u1_n485 ) , .A1( u0_u1_n710 ) , .B2( u0_u1_n787 ) , .A2( u0_u1_n808 ) , .B1( u0_u1_n814 ) );
  NOR2_X1 u0_u1_U334 (.ZN( u0_u1_n613 ) , .A2( u0_u1_n782 ) , .A1( u0_u1_n808 ) );
  INV_X1 u0_u1_U335 (.A( u0_u1_n808 ) , .ZN( u0_u1_n842 ) );
  NAND2_X1 u0_u1_U336 (.ZN( u0_u1_n673 ) , .A1( u0_u1_n808 ) , .A2( u0_u1_n818 ) );
  NOR2_X1 u0_u1_U337 (.ZN( u0_u1_n464 ) , .A2( w3_8 ) , .A1( w3_9 ) );
  NOR2_X1 u0_u1_U338 (.ZN( u0_u1_n473 ) , .A1( u0_u1_n828 ) , .A2( w3_9 ) );
  INV_X1 u0_u1_U339 (.ZN( u0_u1_n829 ) , .A( w3_9 ) );
  NOR2_X1 u0_u1_U34 (.ZN( u0_u1_n806 ) , .A1( u0_u1_n855 ) , .A2( u0_u1_n862 ) );
  NAND2_X2 u0_u1_U340 (.A1( u0_u1_n457 ) , .A2( u0_u1_n464 ) , .ZN( u0_u1_n752 ) );
  NOR2_X1 u0_u1_U341 (.ZN( u0_u1_n463 ) , .A1( u0_u1_n831 ) , .A2( w3_10 ) );
  INV_X1 u0_u1_U342 (.ZN( u0_u1_n830 ) , .A( w3_10 ) );
  AOI211_X1 u0_u1_U343 (.A( u0_u1_n590 ) , .ZN( u0_u1_n599 ) , .B( u0_u1_n623 ) , .C1( u0_u1_n846 ) , .C2( u0_u1_n856 ) );
  NOR3_X1 u0_u1_U344 (.A3( u0_u1_n623 ) , .A2( u0_u1_n624 ) , .ZN( u0_u1_n638 ) , .A1( u0_u1_n727 ) );
  AOI211_X1 u0_u1_U345 (.B( u0_u1_n479 ) , .A( u0_u1_n480 ) , .ZN( u0_u1_n484 ) , .C2( u0_u1_n835 ) , .C1( u0_u1_n862 ) );
  AOI222_X1 u0_u1_U346 (.ZN( u0_u1_n608 ) , .A1( u0_u1_n832 ) , .C2( u0_u1_n838 ) , .B1( u0_u1_n843 ) , .A2( u0_u1_n857 ) , .B2( u0_u1_n862 ) , .C1( u0_u1_n869 ) );
  AOI21_X1 u0_u1_U347 (.ZN( u0_u1_n595 ) , .B1( u0_u1_n752 ) , .A( u0_u1_n794 ) , .B2( u0_u1_n815 ) );
  AOI21_X1 u0_u1_U348 (.A( u0_u1_n814 ) , .B2( u0_u1_n815 ) , .B1( u0_u1_n816 ) , .ZN( u0_u1_n821 ) );
  AOI21_X1 u0_u1_U349 (.ZN( u0_u1_n651 ) , .B1( u0_u1_n731 ) , .B2( u0_u1_n765 ) , .A( u0_u1_n815 ) );
  NAND4_X1 u0_u1_U35 (.A4( u0_u1_n659 ) , .A3( u0_u1_n660 ) , .A2( u0_u1_n661 ) , .A1( u0_u1_n662 ) , .ZN( u0_u1_n802 ) );
  NOR4_X1 u0_u1_U350 (.A4( u0_u1_n616 ) , .A3( u0_u1_n617 ) , .A2( u0_u1_n618 ) , .A1( u0_u1_n619 ) , .ZN( u0_u1_n620 ) );
  NOR2_X1 u0_u1_U351 (.A1( u0_u1_n671 ) , .ZN( u0_u1_n768 ) , .A2( u0_u1_n815 ) );
  NOR2_X1 u0_u1_U352 (.A2( u0_u1_n815 ) , .A1( u0_u1_n817 ) , .ZN( u0_u1_n823 ) );
  NOR2_X1 u0_u1_U353 (.ZN( u0_u1_n580 ) , .A1( u0_u1_n710 ) , .A2( u0_u1_n815 ) );
  NOR2_X1 u0_u1_U354 (.ZN( u0_u1_n667 ) , .A1( u0_u1_n782 ) , .A2( u0_u1_n815 ) );
  NOR2_X1 u0_u1_U355 (.ZN( u0_u1_n686 ) , .A1( u0_u1_n793 ) , .A2( u0_u1_n815 ) );
  NOR2_X1 u0_u1_U356 (.A1( u0_u1_n701 ) , .ZN( u0_u1_n770 ) , .A2( u0_u1_n815 ) );
  NOR2_X1 u0_u1_U357 (.ZN( u0_u1_n656 ) , .A1( u0_u1_n730 ) , .A2( u0_u1_n815 ) );
  NOR2_X1 u0_u1_U358 (.ZN( u0_u1_n633 ) , .A1( u0_u1_n726 ) , .A2( u0_u1_n815 ) );
  NOR2_X1 u0_u1_U359 (.ZN( u0_u1_n457 ) , .A1( u0_u1_n830 ) , .A2( w3_11 ) );
  NOR3_X1 u0_u1_U36 (.A3( u0_u1_n650 ) , .A2( u0_u1_n651 ) , .A1( u0_u1_n652 ) , .ZN( u0_u1_n661 ) );
  NOR2_X1 u0_u1_U360 (.ZN( u0_u1_n474 ) , .A2( w3_10 ) , .A1( w3_11 ) );
  INV_X1 u0_u1_U361 (.ZN( u0_u1_n831 ) , .A( w3_11 ) );
  INV_X1 u0_u1_U362 (.A( u0_n270 ) , .ZN( u0_u1_n850 ) );
  NOR2_X1 u0_u1_U363 (.A1( u0_n268 ) , .A2( u0_n270 ) , .ZN( u0_u1_n466 ) );
  NOR2_X1 u0_u1_U364 (.ZN( u0_u1_n449 ) , .A2( u0_u1_n850 ) , .A1( u0_u1_n859 ) );
  INV_X1 u0_u1_U365 (.A( u0_n272 ) , .ZN( u0_u1_n849 ) );
  NOR2_X1 u0_u1_U366 (.A2( u0_n272 ) , .ZN( u0_u1_n450 ) , .A1( u0_u1_n848 ) );
  NOR2_X1 u0_u1_U367 (.A2( u0_u1_n438 ) , .ZN( u0_u1_n750 ) , .A1( u0_u1_n862 ) );
  NOR4_X1 u0_u1_U368 (.A4( u0_u1_n778 ) , .A3( u0_u1_n779 ) , .A1( u0_u1_n780 ) , .ZN( u0_u1_n801 ) , .A2( u0_u1_n803 ) );
  NAND4_X1 u0_u1_U369 (.A4( u0_u1_n693 ) , .A3( u0_u1_n694 ) , .A1( u0_u1_n695 ) , .ZN( u0_u1_n778 ) , .A2( u0_u1_n873 ) );
  NOR3_X1 u0_u1_U37 (.A3( u0_u1_n653 ) , .A2( u0_u1_n654 ) , .A1( u0_u1_n655 ) , .ZN( u0_u1_n660 ) );
  INV_X1 u0_u1_U370 (.A( u0_u1_n41 ) , .ZN( u0_u1_n839 ) );
  NOR2_X1 u0_u1_U371 (.A1( u0_u1_n41 ) , .ZN( u0_u1_n772 ) , .A2( u0_u1_n817 ) );
  NAND2_X2 u0_u1_U372 (.A1( u0_u1_n457 ) , .A2( u0_u1_n473 ) , .ZN( u0_u1_n805 ) );
  AOI21_X1 u0_u1_U373 (.B2( u0_u1_n41 ) , .ZN( u0_u1_n573 ) , .B1( u0_u1_n808 ) , .A( u0_u1_n814 ) );
  NOR2_X1 u0_u1_U374 (.A2( u0_u1_n41 ) , .A1( u0_u1_n782 ) , .ZN( u0_u1_n822 ) );
  NOR2_X1 u0_u1_U375 (.A2( u0_u1_n41 ) , .ZN( u0_u1_n634 ) , .A1( u0_u1_n726 ) );
  NOR2_X1 u0_u1_U376 (.A2( u0_u1_n41 ) , .ZN( u0_u1_n568 ) , .A1( u0_u1_n765 ) );
  NOR2_X1 u0_u1_U377 (.A2( u0_u1_n41 ) , .ZN( u0_u1_n664 ) , .A1( u0_u1_n731 ) );
  AOI21_X1 u0_u1_U378 (.B2( u0_u1_n41 ) , .ZN( u0_u1_n480 ) , .A( u0_u1_n751 ) , .B1( u0_u1_n781 ) );
  NOR2_X1 u0_u1_U379 (.A2( u0_u1_n41 ) , .ZN( u0_u1_n718 ) , .A1( u0_u1_n794 ) );
  NOR3_X1 u0_u1_U38 (.A3( u0_u1_n656 ) , .A2( u0_u1_n657 ) , .A1( u0_u1_n658 ) , .ZN( u0_u1_n659 ) );
  NOR2_X1 u0_u1_U380 (.A2( u0_u1_n41 ) , .ZN( u0_u1_n596 ) , .A1( u0_u1_n730 ) );
  NOR2_X1 u0_u1_U381 (.A2( u0_u1_n41 ) , .ZN( u0_u1_n543 ) , .A1( u0_u1_n701 ) );
  NOR2_X1 u0_u1_U382 (.ZN( u0_u1_n582 ) , .A2( u0_u1_n699 ) , .A1( u0_u1_n793 ) );
  NAND4_X1 u0_u1_U383 (.ZN( u0_subword_18 ) , .A4( u0_u1_n645 ) , .A3( u0_u1_n646 ) , .A2( u0_u1_n647 ) , .A1( u0_u1_n648 ) );
  OAI21_X1 u0_u1_U384 (.A( u0_u1_n733 ) , .B1( u0_u1_n734 ) , .ZN( u0_u1_n738 ) , .B2( u0_u1_n807 ) );
  OAI222_X1 u0_u1_U385 (.B2( u0_u1_n749 ) , .B1( u0_u1_n750 ) , .A2( u0_u1_n751 ) , .ZN( u0_u1_n759 ) , .C2( u0_u1_n807 ) , .C1( u0_u1_n816 ) , .A1( u0_u1_n819 ) );
  OAI22_X1 u0_u1_U386 (.B2( u0_u1_n805 ) , .B1( u0_u1_n806 ) , .A2( u0_u1_n807 ) , .A1( u0_u1_n808 ) , .ZN( u0_u1_n810 ) );
  AOI21_X1 u0_u1_U387 (.ZN( u0_u1_n652 ) , .A( u0_u1_n781 ) , .B1( u0_u1_n794 ) , .B2( u0_u1_n807 ) );
  INV_X1 u0_u1_U388 (.A( u0_u1_n807 ) , .ZN( u0_u1_n861 ) );
  NOR2_X1 u0_u1_U389 (.ZN( u0_u1_n737 ) , .A2( u0_u1_n805 ) , .A1( u0_u1_n807 ) );
  OAI21_X1 u0_u1_U39 (.ZN( u0_u1_n733 ) , .A( u0_u1_n835 ) , .B2( u0_u1_n853 ) , .B1( u0_u1_n874 ) );
  NOR2_X1 u0_u1_U390 (.ZN( u0_u1_n486 ) , .A1( u0_u1_n790 ) , .A2( u0_u1_n807 ) );
  NOR2_X1 u0_u1_U391 (.ZN( u0_u1_n569 ) , .A1( u0_u1_n749 ) , .A2( u0_u1_n807 ) );
  AOI21_X1 u0_u1_U392 (.A( u0_u1_n41 ) , .ZN( u0_u1_n554 ) , .B1( u0_u1_n671 ) , .B2( u0_u1_n807 ) );
  NAND2_X1 u0_u1_U393 (.ZN( u0_u1_n755 ) , .A1( u0_u1_n765 ) , .A2( u0_u1_n807 ) );
  NOR2_X1 u0_u1_U394 (.ZN( u0_u1_n717 ) , .A1( u0_u1_n807 ) , .A2( u0_u1_n819 ) );
  NOR2_X1 u0_u1_U395 (.ZN( u0_u1_n558 ) , .A1( u0_u1_n764 ) , .A2( u0_u1_n807 ) );
  NOR2_X1 u0_u1_U396 (.ZN( u0_u1_n672 ) , .A1( u0_u1_n792 ) , .A2( u0_u1_n807 ) );
  NAND4_X1 u0_u1_U397 (.ZN( u0_subword_19 ) , .A4( u0_u1_n706 ) , .A3( u0_u1_n707 ) , .A2( u0_u1_n708 ) , .A1( u0_u1_n709 ) );
  INV_X1 u0_u1_U398 (.A( u0_u1_n708 ) , .ZN( u0_u1_n877 ) );
  OAI22_X1 u0_u1_U399 (.B2( u0_u1_n746 ) , .ZN( u0_u1_n748 ) , .A2( u0_u1_n764 ) , .B1( u0_u1_n782 ) , .A1( u0_u1_n794 ) );
  NAND2_X1 u0_u1_U4 (.A2( u0_u1_n462 ) , .A1( u0_u1_n467 ) , .ZN( u0_u1_n782 ) );
  INV_X1 u0_u1_U40 (.A( u0_u1_n681 ) , .ZN( u0_u1_n873 ) );
  OAI22_X1 u0_u1_U400 (.ZN( u0_u1_n498 ) , .A2( u0_u1_n746 ) , .A1( u0_u1_n782 ) , .B1( u0_u1_n793 ) , .B2( u0_u1_n808 ) );
  NOR2_X1 u0_u1_U401 (.ZN( u0_u1_n518 ) , .A1( u0_u1_n710 ) , .A2( u0_u1_n746 ) );
  OAI22_X1 u0_u1_U402 (.ZN( u0_u1_n712 ) , .A2( u0_u1_n730 ) , .B2( u0_u1_n731 ) , .A1( u0_u1_n746 ) , .B1( u0_u1_n815 ) );
  NOR2_X1 u0_u1_U403 (.A2( u0_u1_n746 ) , .ZN( u0_u1_n771 ) , .A1( u0_u1_n814 ) );
  OAI22_X1 u0_u1_U404 (.B1( u0_u1_n442 ) , .ZN( u0_u1_n446 ) , .A2( u0_u1_n730 ) , .A1( u0_u1_n746 ) , .B2( u0_u1_n751 ) );
  NOR2_X1 u0_u1_U405 (.ZN( u0_u1_n549 ) , .A1( u0_u1_n701 ) , .A2( u0_u1_n746 ) );
  NOR2_X1 u0_u1_U406 (.ZN( u0_u1_n532 ) , .A2( u0_u1_n746 ) , .A1( u0_u1_n794 ) );
  NOR2_X1 u0_u1_U407 (.A2( u0_u1_n746 ) , .ZN( u0_u1_n757 ) , .A1( u0_u1_n807 ) );
  NOR2_X1 u0_u1_U408 (.A1( u0_u1_n671 ) , .ZN( u0_u1_n675 ) , .A2( u0_u1_n746 ) );
  NOR2_X1 u0_u1_U409 (.ZN( u0_u1_n720 ) , .A2( u0_u1_n726 ) , .A1( u0_u1_n746 ) );
  NOR4_X1 u0_u1_U41 (.A4( u0_u1_n689 ) , .A3( u0_u1_n690 ) , .A2( u0_u1_n691 ) , .A1( u0_u1_n692 ) , .ZN( u0_u1_n693 ) );
  NOR2_X1 u0_u1_U410 (.ZN( u0_u1_n584 ) , .A1( u0_u1_n746 ) , .A2( u0_u1_n817 ) );
  INV_X1 u0_u1_U411 (.A( u0_u1_n746 ) , .ZN( u0_u1_n838 ) );
  AOI221_X1 u0_u1_U412 (.A( u0_u1_n578 ) , .ZN( u0_u1_n589 ) , .B2( u0_u1_n833 ) , .C2( u0_u1_n844 ) , .B1( u0_u1_n855 ) , .C1( u0_u1_n862 ) );
  AOI21_X1 u0_u1_U413 (.ZN( u0_u1_n578 ) , .B2( u0_u1_n726 ) , .B1( u0_u1_n750 ) , .A( u0_u1_n787 ) );
  AOI211_X1 u0_u1_U414 (.A( u0_u1_n639 ) , .ZN( u0_u1_n647 ) , .B( u0_u1_n745 ) , .C2( u0_u1_n840 ) , .C1( u0_u1_n855 ) );
  NAND4_X1 u0_u1_U415 (.A4( u0_u1_n635 ) , .A3( u0_u1_n636 ) , .A2( u0_u1_n637 ) , .A1( u0_u1_n638 ) , .ZN( u0_u1_n745 ) );
  OAI22_X1 u0_u1_U416 (.B1( u0_u1_n441 ) , .ZN( u0_u1_n590 ) , .A2( u0_u1_n749 ) , .B2( u0_u1_n764 ) , .A1( u0_u1_n765 ) );
  NAND2_X1 u0_u1_U417 (.A2( u0_u1_n441 ) , .A1( u0_u1_n731 ) , .ZN( u0_u1_n813 ) );
  AOI21_X1 u0_u1_U418 (.B2( u0_u1_n441 ) , .ZN( u0_u1_n594 ) , .B1( u0_u1_n730 ) , .A( u0_u1_n792 ) );
  AOI21_X1 u0_u1_U419 (.B2( u0_u1_n441 ) , .ZN( u0_u1_n650 ) , .A( u0_u1_n764 ) , .B1( u0_u1_n794 ) );
  AOI221_X1 u0_u1_U42 (.A( u0_u1_n683 ) , .ZN( u0_u1_n694 ) , .B2( u0_u1_n841 ) , .C1( u0_u1_n843 ) , .C2( u0_u1_n863 ) , .B1( u0_u1_n866 ) );
  AOI21_X1 u0_u1_U420 (.B2( u0_u1_n441 ) , .ZN( u0_u1_n625 ) , .B1( u0_u1_n701 ) , .A( u0_u1_n781 ) );
  OAI22_X1 u0_u1_U421 (.B2( u0_u1_n441 ) , .ZN( u0_u1_n683 ) , .A1( u0_u1_n701 ) , .A2( u0_u1_n732 ) , .B1( u0_u1_n819 ) );
  NOR2_X1 u0_u1_U422 (.ZN( u0_u1_n653 ) , .A1( u0_u1_n786 ) , .A2( u0_u1_n790 ) );
  OAI21_X1 u0_u1_U423 (.B2( u0_u1_n441 ) , .A( u0_u1_n615 ) , .ZN( u0_u1_n618 ) , .B1( u0_u1_n627 ) );
  NOR2_X1 u0_u1_U424 (.A1( u0_u1_n441 ) , .ZN( u0_u1_n612 ) , .A2( u0_u1_n818 ) );
  NOR2_X1 u0_u1_U425 (.ZN( u0_u1_n555 ) , .A2( u0_u1_n746 ) , .A1( u0_u1_n786 ) );
  NOR2_X1 u0_u1_U426 (.A2( u0_u1_n41 ) , .ZN( u0_u1_n602 ) , .A1( u0_u1_n786 ) );
  AOI21_X1 u0_u1_U427 (.A( u0_u1_n41 ) , .ZN( u0_u1_n502 ) , .B1( u0_u1_n710 ) , .B2( u0_u1_n788 ) );
  OAI22_X1 u0_u1_U428 (.ZN( u0_u1_n592 ) , .B1( u0_u1_n732 ) , .B2( u0_u1_n751 ) , .A2( u0_u1_n788 ) , .A1( u0_u1_n805 ) );
  AOI222_X1 u0_u1_U429 (.ZN( u0_u1_n515 ) , .C1( u0_u1_n834 ) , .B2( u0_u1_n838 ) , .A2( u0_u1_n844 ) , .C2( u0_u1_n863 ) , .B1( u0_u1_n864 ) , .A1( u0_u1_n867 ) );
  NOR4_X1 u0_u1_U43 (.A4( u0_u1_n528 ) , .A2( u0_u1_n529 ) , .A1( u0_u1_n530 ) , .ZN( u0_u1_n540 ) , .A3( u0_u1_n703 ) );
  AOI222_X1 u0_u1_U430 (.ZN( u0_u1_n607 ) , .B2( u0_u1_n673 ) , .B1( u0_u1_n755 ) , .C2( u0_u1_n833 ) , .A1( u0_u1_n835 ) , .A2( u0_u1_n863 ) , .C1( u0_u1_n864 ) );
  AOI221_X1 u0_u1_U431 (.A( u0_u1_n485 ) , .ZN( u0_u1_n490 ) , .B1( u0_u1_n833 ) , .C2( u0_u1_n845 ) , .C1( u0_u1_n853 ) , .B2( u0_u1_n863 ) );
  NOR2_X1 u0_u1_U432 (.ZN( u0_u1_n655 ) , .A1( u0_u1_n764 ) , .A2( u0_u1_n788 ) );
  NAND2_X1 u0_u1_U433 (.A2( u0_u1_n751 ) , .A1( u0_u1_n788 ) , .ZN( u0_u1_n811 ) );
  NOR2_X1 u0_u1_U434 (.ZN( u0_u1_n556 ) , .A1( u0_u1_n788 ) , .A2( u0_u1_n815 ) );
  NOR2_X1 u0_u1_U435 (.ZN( u0_u1_n614 ) , .A1( u0_u1_n781 ) , .A2( u0_u1_n788 ) );
  NOR2_X1 u0_u1_U436 (.ZN( u0_u1_n719 ) , .A2( u0_u1_n746 ) , .A1( u0_u1_n788 ) );
  NAND3_X1 u0_u1_U437 (.ZN( u0_subword_22 ) , .A3( u0_u1_n799 ) , .A2( u0_u1_n800 ) , .A1( u0_u1_n801 ) );
  NAND3_X1 u0_u1_U438 (.ZN( u0_subword_21 ) , .A3( u0_u1_n760 ) , .A2( u0_u1_n761 ) , .A1( u0_u1_n762 ) );
  NAND3_X1 u0_u1_U439 (.ZN( u0_subword_20 ) , .A3( u0_u1_n740 ) , .A2( u0_u1_n741 ) , .A1( u0_u1_n742 ) );
  NOR4_X1 u0_u1_U44 (.A4( u0_u1_n534 ) , .A3( u0_u1_n535 ) , .A2( u0_u1_n536 ) , .ZN( u0_u1_n537 ) , .A1( u0_u1_n822 ) );
  NAND3_X1 u0_u1_U440 (.A3( u0_u1_n677 ) , .A2( u0_u1_n678 ) , .A1( u0_u1_n679 ) , .ZN( u0_u1_n809 ) );
  NAND3_X1 u0_u1_U441 (.ZN( u0_u1_n640 ) , .A3( u0_u1_n710 ) , .A2( u0_u1_n726 ) , .A1( u0_u1_n794 ) );
  NAND3_X1 u0_u1_U442 (.A3( u0_u1_n620 ) , .A2( u0_u1_n621 ) , .A1( u0_u1_n622 ) , .ZN( u0_u1_n727 ) );
  NAND3_X1 u0_u1_U443 (.A3( u0_u1_n587 ) , .A2( u0_u1_n588 ) , .A1( u0_u1_n589 ) , .ZN( u0_u1_n623 ) );
  NAND3_X1 u0_u1_U444 (.ZN( u0_u1_n567 ) , .A3( u0_u1_n682 ) , .A2( u0_u1_n752 ) , .A1( u0_u1_n787 ) );
  NAND3_X1 u0_u1_U445 (.A3( u0_u1_n525 ) , .A2( u0_u1_n526 ) , .A1( u0_u1_n527 ) , .ZN( u0_u1_n744 ) );
  NAND3_X1 u0_u1_U446 (.A3( u0_u1_n514 ) , .A1( u0_u1_n515 ) , .ZN( u0_u1_n610 ) , .A2( u0_u1_n872 ) );
  NAND3_X1 u0_u1_U447 (.A3( u0_u1_n469 ) , .A2( u0_u1_n470 ) , .A1( u0_u1_n471 ) , .ZN( u0_u1_n779 ) );
  NOR2_X1 u0_u1_U448 (.ZN( u0_u1_n791 ) , .A2( u0_u1_n863 ) , .A1( u0_u1_n869 ) );
  NOR2_X1 u0_u1_U449 (.ZN( u0_u1_n703 ) , .A2( u0_u1_n788 ) , .A1( u0_u1_n819 ) );
  NOR4_X1 u0_u1_U45 (.A4( u0_u1_n531 ) , .A3( u0_u1_n532 ) , .ZN( u0_u1_n539 ) , .A2( u0_u1_n686 ) , .A1( u0_u1_n796 ) );
  NOR2_X1 u0_u1_U450 (.A1( u0_u1_n732 ) , .ZN( u0_u1_n767 ) , .A2( u0_u1_n788 ) );
  INV_X1 u0_u1_U451 (.A( u0_u1_n788 ) , .ZN( u0_u1_n863 ) );
  NOR3_X1 u0_u1_U46 (.A3( u0_u1_n802 ) , .A2( u0_u1_n803 ) , .A1( u0_u1_n804 ) , .ZN( u0_u1_n827 ) );
  NAND4_X1 u0_u1_U47 (.A4( u0_u1_n481 ) , .A3( u0_u1_n482 ) , .A2( u0_u1_n483 ) , .A1( u0_u1_n484 ) , .ZN( u0_u1_n696 ) );
  NOR3_X1 u0_u1_U48 (.ZN( u0_u1_n482 ) , .A2( u0_u1_n510 ) , .A3( u0_u1_n603 ) , .A1( u0_u1_n612 ) );
  NOR4_X1 u0_u1_U49 (.ZN( u0_u1_n481 ) , .A1( u0_u1_n522 ) , .A4( u0_u1_n559 ) , .A3( u0_u1_n584 ) , .A2( u0_u1_n632 ) );
  NOR3_X1 u0_u1_U5 (.ZN( u0_u1_n600 ) , .A1( u0_u1_n610 ) , .A3( u0_u1_n725 ) , .A2( u0_u1_n744 ) );
  NAND4_X1 u0_u1_U50 (.A4( u0_u1_n774 ) , .A3( u0_u1_n775 ) , .A2( u0_u1_n776 ) , .A1( u0_u1_n777 ) , .ZN( u0_u1_n803 ) );
  NOR3_X1 u0_u1_U51 (.A3( u0_u1_n767 ) , .A2( u0_u1_n768 ) , .A1( u0_u1_n769 ) , .ZN( u0_u1_n775 ) );
  NOR4_X1 u0_u1_U52 (.A4( u0_u1_n770 ) , .A3( u0_u1_n771 ) , .A2( u0_u1_n772 ) , .A1( u0_u1_n773 ) , .ZN( u0_u1_n774 ) );
  NAND4_X1 u0_u1_U53 (.A4( u0_u1_n562 ) , .A3( u0_u1_n563 ) , .A2( u0_u1_n564 ) , .A1( u0_u1_n565 ) , .ZN( u0_u1_n609 ) );
  NOR4_X1 u0_u1_U54 (.A4( u0_u1_n554 ) , .A3( u0_u1_n555 ) , .A2( u0_u1_n556 ) , .A1( u0_u1_n557 ) , .ZN( u0_u1_n564 ) );
  AOI222_X1 u0_u1_U55 (.ZN( u0_u1_n565 ) , .B1( u0_u1_n832 ) , .C1( u0_u1_n842 ) , .A2( u0_u1_n844 ) , .A1( u0_u1_n855 ) , .B2( u0_u1_n864 ) , .C2( u0_u1_n874 ) );
  NOR4_X1 u0_u1_U56 (.A4( u0_u1_n558 ) , .A3( u0_u1_n559 ) , .A2( u0_u1_n560 ) , .A1( u0_u1_n561 ) , .ZN( u0_u1_n562 ) );
  INV_X1 u0_u1_U57 (.A( u0_u1_n507 ) , .ZN( u0_u1_n872 ) );
  NOR4_X1 u0_u1_U58 (.A4( u0_u1_n511 ) , .A2( u0_u1_n512 ) , .A1( u0_u1_n513 ) , .ZN( u0_u1_n514 ) , .A3( u0_u1_n672 ) );
  NOR4_X1 u0_u1_U59 (.A4( u0_u1_n663 ) , .A3( u0_u1_n664 ) , .A2( u0_u1_n665 ) , .A1( u0_u1_n666 ) , .ZN( u0_u1_n679 ) );
  NOR3_X1 u0_u1_U6 (.A2( u0_u1_n609 ) , .A1( u0_u1_n610 ) , .ZN( u0_u1_n648 ) , .A3( u0_u1_n724 ) );
  NOR4_X1 u0_u1_U60 (.A4( u0_u1_n667 ) , .A3( u0_u1_n668 ) , .A2( u0_u1_n669 ) , .A1( u0_u1_n670 ) , .ZN( u0_u1_n678 ) );
  NOR4_X1 u0_u1_U61 (.A3( u0_u1_n675 ) , .A1( u0_u1_n676 ) , .ZN( u0_u1_n677 ) , .A4( u0_u1_n717 ) , .A2( u0_u1_n860 ) );
  AOI221_X1 u0_u1_U62 (.ZN( u0_u1_n470 ) , .C2( u0_u1_n716 ) , .B2( u0_u1_n833 ) , .C1( u0_u1_n846 ) , .B1( u0_u1_n861 ) , .A( u0_u1_n865 ) );
  NOR4_X1 u0_u1_U63 (.A1( u0_u1_n468 ) , .ZN( u0_u1_n469 ) , .A4( u0_u1_n544 ) , .A2( u0_u1_n556 ) , .A3( u0_u1_n616 ) );
  NAND4_X1 u0_u1_U64 (.A4( u0_u1_n487 ) , .A3( u0_u1_n488 ) , .A2( u0_u1_n489 ) , .A1( u0_u1_n490 ) , .ZN( u0_u1_n780 ) );
  NOR4_X1 u0_u1_U65 (.A4( u0_u1_n486 ) , .ZN( u0_u1_n489 ) , .A1( u0_u1_n568 ) , .A2( u0_u1_n583 ) , .A3( u0_u1_n604 ) );
  NOR4_X1 u0_u1_U66 (.ZN( u0_u1_n488 ) , .A1( u0_u1_n509 ) , .A2( u0_u1_n521 ) , .A4( u0_u1_n548 ) , .A3( u0_u1_n613 ) );
  NOR2_X1 u0_u1_U67 (.ZN( u0_u1_n763 ) , .A1( u0_u1_n835 ) , .A2( u0_u1_n836 ) );
  NOR4_X1 u0_u1_U68 (.A4( u0_u1_n516 ) , .A3( u0_u1_n517 ) , .A2( u0_u1_n518 ) , .A1( u0_u1_n519 ) , .ZN( u0_u1_n526 ) );
  NOR4_X1 u0_u1_U69 (.A3( u0_u1_n523 ) , .A1( u0_u1_n524 ) , .ZN( u0_u1_n525 ) , .A2( u0_u1_n675 ) , .A4( u0_u1_n771 ) );
  NOR3_X1 u0_u1_U7 (.A3( u0_u1_n724 ) , .A1( u0_u1_n725 ) , .ZN( u0_u1_n742 ) , .A2( u0_u1_n743 ) );
  NAND4_X1 u0_u1_U70 (.A4( u0_u1_n475 ) , .A3( u0_u1_n476 ) , .A2( u0_u1_n477 ) , .A1( u0_u1_n478 ) , .ZN( u0_u1_n680 ) );
  NOR4_X1 u0_u1_U71 (.ZN( u0_u1_n476 ) , .A1( u0_u1_n508 ) , .A3( u0_u1_n546 ) , .A2( u0_u1_n585 ) , .A4( u0_u1_n718 ) );
  NOR4_X1 u0_u1_U72 (.ZN( u0_u1_n475 ) , .A2( u0_u1_n523 ) , .A4( u0_u1_n596 ) , .A1( u0_u1_n611 ) , .A3( u0_u1_n631 ) );
  NOR4_X1 u0_u1_U73 (.A4( u0_u1_n472 ) , .ZN( u0_u1_n478 ) , .A3( u0_u1_n558 ) , .A1( u0_u1_n737 ) , .A2( u0_u1_n757 ) );
  NAND4_X1 u0_u1_U74 (.A4( u0_u1_n458 ) , .A3( u0_u1_n459 ) , .A2( u0_u1_n460 ) , .A1( u0_u1_n461 ) , .ZN( u0_u1_n681 ) );
  NOR3_X1 u0_u1_U75 (.ZN( u0_u1_n459 ) , .A3( u0_u1_n532 ) , .A1( u0_u1_n557 ) , .A2( u0_u1_n572 ) );
  AOI221_X1 u0_u1_U76 (.A( u0_u1_n452 ) , .ZN( u0_u1_n461 ) , .C2( u0_u1_n755 ) , .B1( u0_u1_n834 ) , .C1( u0_u1_n843 ) , .B2( u0_u1_n862 ) );
  NOR4_X1 u0_u1_U77 (.ZN( u0_u1_n460 ) , .A2( u0_u1_n511 ) , .A1( u0_u1_n601 ) , .A4( u0_u1_n630 ) , .A3( u0_u1_n713 ) );
  INV_X1 u0_u1_U78 (.A( u0_u1_n671 ) , .ZN( u0_u1_n866 ) );
  NAND4_X1 u0_u1_U79 (.A4( u0_u1_n575 ) , .A3( u0_u1_n576 ) , .A1( u0_u1_n577 ) , .ZN( u0_u1_n725 ) , .A2( u0_u1_n875 ) );
  NOR3_X1 u0_u1_U8 (.ZN( u0_u1_n506 ) , .A2( u0_u1_n681 ) , .A3( u0_u1_n779 ) , .A1( u0_u1_n877 ) );
  NOR4_X1 u0_u1_U80 (.A4( u0_u1_n571 ) , .A3( u0_u1_n572 ) , .A2( u0_u1_n573 ) , .A1( u0_u1_n574 ) , .ZN( u0_u1_n575 ) );
  AOI221_X1 u0_u1_U81 (.A( u0_u1_n566 ) , .C2( u0_u1_n567 ) , .ZN( u0_u1_n576 ) , .B2( u0_u1_n846 ) , .B1( u0_u1_n853 ) , .C1( u0_u1_n854 ) );
  NOR2_X1 u0_u1_U82 (.ZN( u0_u1_n577 ) , .A1( u0_u1_n624 ) , .A2( u0_u1_n747 ) );
  INV_X1 u0_u1_U83 (.A( u0_u1_n764 ) , .ZN( u0_u1_n832 ) );
  NOR2_X1 u0_u1_U84 (.ZN( u0_u1_n649 ) , .A1( u0_u1_n855 ) , .A2( u0_u1_n869 ) );
  NOR4_X1 u0_u1_U85 (.A4( u0_u1_n579 ) , .A3( u0_u1_n580 ) , .A2( u0_u1_n581 ) , .ZN( u0_u1_n588 ) , .A1( u0_u1_n685 ) );
  NOR4_X1 u0_u1_U86 (.A1( u0_u1_n586 ) , .ZN( u0_u1_n587 ) , .A3( u0_u1_n654 ) , .A2( u0_u1_n664 ) , .A4( u0_u1_n769 ) );
  NAND4_X1 u0_u1_U87 (.A4( u0_u1_n721 ) , .A3( u0_u1_n722 ) , .A2( u0_u1_n723 ) , .ZN( u0_u1_n743 ) , .A1( u0_u1_n858 ) );
  NOR4_X1 u0_u1_U88 (.A4( u0_u1_n717 ) , .A3( u0_u1_n718 ) , .A2( u0_u1_n719 ) , .A1( u0_u1_n720 ) , .ZN( u0_u1_n721 ) );
  INV_X1 u0_u1_U89 (.A( u0_u1_n711 ) , .ZN( u0_u1_n858 ) );
  NOR2_X1 u0_u1_U9 (.ZN( u0_u1_n497 ) , .A1( u0_u1_n680 ) , .A2( u0_u1_n696 ) );
  AOI221_X1 u0_u1_U90 (.A( u0_u1_n712 ) , .ZN( u0_u1_n723 ) , .C2( u0_u1_n845 ) , .B2( u0_u1_n846 ) , .C1( u0_u1_n862 ) , .B1( u0_u1_n863 ) );
  INV_X1 u0_u1_U91 (.A( u0_u1_n465 ) , .ZN( u0_u1_n865 ) );
  OAI21_X1 u0_u1_U92 (.ZN( u0_u1_n465 ) , .B1( u0_u1_n811 ) , .A( u0_u1_n836 ) , .B2( u0_u1_n852 ) );
  INV_X1 u0_u1_U93 (.A( u0_u1_n793 ) , .ZN( u0_u1_n874 ) );
  OR4_X1 u0_u1_U94 (.A4( u0_u1_n568 ) , .A3( u0_u1_n569 ) , .A2( u0_u1_n570 ) , .ZN( u0_u1_n574 ) , .A1( u0_u1_n667 ) );
  OR4_X1 u0_u1_U95 (.A4( u0_u1_n520 ) , .A2( u0_u1_n521 ) , .A1( u0_u1_n522 ) , .ZN( u0_u1_n524 ) , .A3( u0_u1_n823 ) );
  OR4_X1 u0_u1_U96 (.ZN( u0_u1_n494 ) , .A4( u0_u1_n536 ) , .A2( u0_u1_n549 ) , .A1( u0_u1_n561 ) , .A3( u0_u1_n634 ) );
  OR4_X1 u0_u1_U97 (.ZN( u0_u1_n468 ) , .A4( u0_u1_n520 ) , .A3( u0_u1_n531 ) , .A2( u0_u1_n580 ) , .A1( u0_u1_n714 ) );
  OR4_X1 u0_u1_U98 (.A4( u0_u1_n684 ) , .A3( u0_u1_n685 ) , .A2( u0_u1_n686 ) , .A1( u0_u1_n687 ) , .ZN( u0_u1_n692 ) );
  OR3_X1 u0_u1_U99 (.A3( u0_u1_n508 ) , .A2( u0_u1_n509 ) , .A1( u0_u1_n510 ) , .ZN( u0_u1_n513 ) );
  NOR2_X1 us02_U10 (.ZN( us02_n574 ) , .A1( us02_n621 ) , .A2( us02_n744 ) );
  NOR2_X1 us02_U100 (.ZN( us02_n685 ) , .A1( us02_n830 ) , .A2( us02_n831 ) );
  NOR4_X1 us02_U101 (.ZN( us02_n619 ) , .A1( us02_n655 ) , .A3( us02_n665 ) , .A4( us02_n681 ) , .A2( us02_n765 ) );
  NOR4_X1 us02_U102 (.A4( us02_n608 ) , .A3( us02_n609 ) , .A2( us02_n610 ) , .A1( us02_n611 ) , .ZN( us02_n618 ) );
  NOR4_X1 us02_U103 (.A4( us02_n613 ) , .A3( us02_n614 ) , .A2( us02_n615 ) , .A1( us02_n616 ) , .ZN( us02_n617 ) );
  NAND4_X1 us02_U104 (.A4( us02_n484 ) , .A3( us02_n485 ) , .A2( us02_n486 ) , .A1( us02_n487 ) , .ZN( us02_n777 ) );
  NOR4_X1 us02_U105 (.A4( us02_n483 ) , .ZN( us02_n486 ) , .A1( us02_n565 ) , .A2( us02_n580 ) , .A3( us02_n601 ) );
  NOR4_X1 us02_U106 (.ZN( us02_n485 ) , .A1( us02_n506 ) , .A2( us02_n518 ) , .A4( us02_n545 ) , .A3( us02_n610 ) );
  NOR4_X1 us02_U107 (.ZN( us02_n484 ) , .A2( us02_n532 ) , .A1( us02_n557 ) , .A3( us02_n630 ) , .A4( us02_n717 ) );
  NAND4_X1 us02_U108 (.A4( us02_n690 ) , .A3( us02_n691 ) , .A1( us02_n692 ) , .ZN( us02_n775 ) , .A2( us02_n871 ) );
  AOI221_X1 us02_U109 (.A( us02_n680 ) , .ZN( us02_n691 ) , .B2( us02_n839 ) , .C1( us02_n841 ) , .C2( us02_n861 ) , .B1( us02_n864 ) );
  NOR2_X1 us02_U11 (.A1( us02_n677 ) , .ZN( us02_n692 ) , .A2( us02_n806 ) );
  INV_X1 us02_U110 (.A( us02_n678 ) , .ZN( us02_n871 ) );
  NOR4_X1 us02_U111 (.A4( us02_n686 ) , .A3( us02_n687 ) , .A2( us02_n688 ) , .A1( us02_n689 ) , .ZN( us02_n690 ) );
  NAND4_X1 us02_U112 (.A4( us02_n559 ) , .A3( us02_n560 ) , .A2( us02_n561 ) , .A1( us02_n562 ) , .ZN( us02_n606 ) );
  NOR4_X1 us02_U113 (.ZN( us02_n560 ) , .A1( us02_n652 ) , .A3( us02_n660 ) , .A4( us02_n684 ) , .A2( us02_n767 ) );
  NOR4_X1 us02_U114 (.A4( us02_n551 ) , .A3( us02_n552 ) , .A2( us02_n553 ) , .A1( us02_n554 ) , .ZN( us02_n561 ) );
  NOR4_X1 us02_U115 (.A4( us02_n555 ) , .A3( us02_n556 ) , .A2( us02_n557 ) , .A1( us02_n558 ) , .ZN( us02_n559 ) );
  NAND4_X1 us02_U116 (.A4( us02_n718 ) , .A3( us02_n719 ) , .A2( us02_n720 ) , .ZN( us02_n740 ) , .A1( us02_n856 ) );
  INV_X1 us02_U117 (.A( us02_n708 ) , .ZN( us02_n856 ) );
  AOI221_X1 us02_U118 (.A( us02_n709 ) , .ZN( us02_n720 ) , .C2( us02_n843 ) , .B2( us02_n844 ) , .C1( us02_n860 ) , .B1( us02_n861 ) );
  NOR4_X1 us02_U119 (.A4( us02_n714 ) , .A3( us02_n715 ) , .A2( us02_n716 ) , .A1( us02_n717 ) , .ZN( us02_n718 ) );
  INV_X1 us02_U12 (.A( us02_n679 ) , .ZN( us02_n839 ) );
  NAND4_X1 us02_U120 (.A4( us02_n472 ) , .A3( us02_n473 ) , .A2( us02_n474 ) , .A1( us02_n475 ) , .ZN( us02_n677 ) );
  NOR4_X1 us02_U121 (.A4( us02_n469 ) , .ZN( us02_n475 ) , .A3( us02_n555 ) , .A1( us02_n734 ) , .A2( us02_n754 ) );
  NOR4_X1 us02_U122 (.ZN( us02_n474 ) , .A1( us02_n530 ) , .A3( us02_n567 ) , .A4( us02_n599 ) , .A2( us02_n641 ) );
  NOR4_X1 us02_U123 (.ZN( us02_n473 ) , .A1( us02_n505 ) , .A3( us02_n543 ) , .A2( us02_n582 ) , .A4( us02_n715 ) );
  NOR2_X1 us02_U124 (.ZN( us02_n732 ) , .A2( us02_n831 ) , .A1( us02_n844 ) );
  NOR2_X1 us02_U125 (.ZN( us02_n788 ) , .A2( us02_n861 ) , .A1( us02_n867 ) );
  NOR2_X1 us02_U126 (.ZN( us02_n646 ) , .A1( us02_n853 ) , .A2( us02_n867 ) );
  NAND4_X1 us02_U127 (.A4( us02_n572 ) , .A3( us02_n573 ) , .A1( us02_n574 ) , .ZN( us02_n722 ) , .A2( us02_n873 ) );
  NOR4_X1 us02_U128 (.A4( us02_n568 ) , .A3( us02_n569 ) , .A2( us02_n570 ) , .A1( us02_n571 ) , .ZN( us02_n572 ) );
  AOI221_X1 us02_U129 (.A( us02_n563 ) , .C2( us02_n564 ) , .ZN( us02_n573 ) , .B2( us02_n844 ) , .B1( us02_n851 ) , .C1( us02_n852 ) );
  NOR4_X1 us02_U13 (.A4( us02_n444 ) , .A3( us02_n445 ) , .A2( us02_n515 ) , .A1( us02_n540 ) , .ZN( us02_n705 ) );
  INV_X1 us02_U130 (.A( us02_n606 ) , .ZN( us02_n873 ) );
  NAND4_X1 us02_U131 (.A4( us02_n492 ) , .A3( us02_n493 ) , .A1( us02_n494 ) , .ZN( us02_n801 ) , .A2( us02_n866 ) );
  AOI221_X1 us02_U132 (.A( us02_n488 ) , .ZN( us02_n493 ) , .B2( us02_n835 ) , .C2( us02_n840 ) , .C1( us02_n850 ) , .B1( us02_n859 ) );
  INV_X1 us02_U133 (.A( us02_n777 ) , .ZN( us02_n866 ) );
  NOR2_X1 us02_U134 (.ZN( us02_n494 ) , .A1( us02_n677 ) , .A2( us02_n693 ) );
  AOI222_X1 us02_U135 (.ZN( us02_n512 ) , .C1( us02_n831 ) , .B2( us02_n836 ) , .A2( us02_n842 ) , .C2( us02_n861 ) , .B1( us02_n862 ) , .A1( us02_n865 ) );
  NOR4_X1 us02_U136 (.A4( us02_n508 ) , .A2( us02_n509 ) , .A1( us02_n510 ) , .ZN( us02_n511 ) , .A3( us02_n669 ) );
  INV_X1 us02_U137 (.A( us02_n504 ) , .ZN( us02_n870 ) );
  INV_X1 us02_U138 (.A( us02_n761 ) , .ZN( us02_n829 ) );
  INV_X1 us02_U139 (.A( us02_n462 ) , .ZN( us02_n863 ) );
  OR3_X1 us02_U14 (.ZN( us02_n445 ) , .A1( us02_n527 ) , .A3( us02_n576 ) , .A2( us02_n874 ) );
  OAI21_X1 us02_U140 (.ZN( us02_n462 ) , .B1( us02_n808 ) , .A( us02_n833 ) , .B2( us02_n850 ) );
  OR4_X1 us02_U141 (.A4( us02_n565 ) , .A3( us02_n566 ) , .A2( us02_n567 ) , .ZN( us02_n571 ) , .A1( us02_n664 ) );
  OR4_X1 us02_U142 (.A4( us02_n517 ) , .A2( us02_n518 ) , .A1( us02_n519 ) , .ZN( us02_n521 ) , .A3( us02_n820 ) );
  OR4_X1 us02_U143 (.ZN( us02_n465 ) , .A4( us02_n517 ) , .A3( us02_n528 ) , .A2( us02_n577 ) , .A1( us02_n711 ) );
  OR4_X1 us02_U144 (.A4( us02_n681 ) , .A3( us02_n682 ) , .A2( us02_n683 ) , .A1( us02_n684 ) , .ZN( us02_n689 ) );
  OR4_X1 us02_U145 (.A4( us02_n579 ) , .A3( us02_n580 ) , .A2( us02_n581 ) , .A1( us02_n582 ) , .ZN( us02_n583 ) );
  NAND2_X1 us02_U146 (.ZN( us02_n612 ) , .A2( us02_n836 ) , .A1( us02_n872 ) );
  OR3_X1 us02_U147 (.A3( us02_n505 ) , .A2( us02_n506 ) , .A1( us02_n507 ) , .ZN( us02_n510 ) );
  AOI221_X1 us02_U148 (.A( us02_n712 ) , .B2( us02_n713 ) , .ZN( us02_n719 ) , .C1( us02_n831 ) , .B1( us02_n838 ) , .C2( us02_n862 ) );
  OR2_X1 us02_U149 (.A2( us02_n710 ) , .A1( us02_n711 ) , .ZN( us02_n712 ) );
  OR4_X1 us02_U15 (.A4( us02_n441 ) , .A2( us02_n442 ) , .A1( us02_n443 ) , .ZN( us02_n444 ) , .A3( us02_n552 ) );
  INV_X1 us02_U150 (.A( us02_n753 ) , .ZN( us02_n868 ) );
  OAI21_X1 us02_U151 (.B1( us02_n752 ) , .ZN( us02_n753 ) , .A( us02_n844 ) , .B2( us02_n867 ) );
  INV_X1 us02_U152 (.A( us02_n671 ) , .ZN( us02_n858 ) );
  AOI21_X1 us02_U153 (.A( us02_n669 ) , .B1( us02_n670 ) , .ZN( us02_n671 ) , .B2( us02_n855 ) );
  NAND2_X1 us02_U154 (.A1( us02_n446 ) , .A2( us02_n464 ) , .ZN( us02_n748 ) );
  OAI222_X1 us02_U155 (.B2( us02_n746 ) , .B1( us02_n747 ) , .A2( us02_n748 ) , .ZN( us02_n756 ) , .C2( us02_n804 ) , .C1( us02_n813 ) , .A1( us02_n816 ) );
  OAI222_X1 us02_U156 (.ZN( us02_n504 ) , .C2( us02_n624 ) , .B2( us02_n646 ) , .B1( us02_n746 ) , .A2( us02_n747 ) , .C1( us02_n804 ) , .A1( us02_n805 ) );
  OAI222_X1 us02_U157 (.B2( us02_n707 ) , .ZN( us02_n708 ) , .C2( us02_n723 ) , .B1( us02_n746 ) , .A1( us02_n805 ) , .C1( us02_n813 ) , .A2( us02_n814 ) );
  OAI222_X1 us02_U158 (.ZN( us02_n616 ) , .B1( us02_n696 ) , .C1( us02_n723 ) , .C2( us02_n746 ) , .B2( us02_n785 ) , .A2( us02_n791 ) , .A1( us02_n815 ) );
  NOR4_X1 us02_U159 (.A2( us02_n490 ) , .A1( us02_n491 ) , .ZN( us02_n492 ) , .A3( us02_n579 ) , .A4( us02_n611 ) );
  INV_X1 us02_U16 (.A( us02_n612 ) , .ZN( us02_n874 ) );
  OR4_X1 us02_U160 (.ZN( us02_n491 ) , .A4( us02_n533 ) , .A2( us02_n546 ) , .A1( us02_n558 ) , .A3( us02_n631 ) );
  OAI22_X1 us02_U161 (.B1( us02_n489 ) , .ZN( us02_n490 ) , .A1( us02_n685 ) , .A2( us02_n762 ) , .B2( us02_n816 ) );
  NOR3_X1 us02_U162 (.ZN( us02_n489 ) , .A1( us02_n781 ) , .A2( us02_n849 ) , .A3( us02_n862 ) );
  AOI22_X1 us02_U163 (.ZN( us02_n695 ) , .A1( us02_n829 ) , .B2( us02_n842 ) , .A2( us02_n864 ) , .B1( us02_n867 ) );
  INV_X1 us02_U164 (.A( us02_n729 ) , .ZN( us02_n838 ) );
  AOI221_X1 us02_U165 (.A( us02_n763 ) , .ZN( us02_n773 ) , .C2( us02_n809 ) , .B2( us02_n834 ) , .C1( us02_n854 ) , .B1( us02_n865 ) );
  AOI21_X1 us02_U166 (.B2( us02_n762 ) , .ZN( us02_n763 ) , .A( us02_n787 ) , .B1( us02_n791 ) );
  INV_X1 us02_U167 (.A( us02_n760 ) , .ZN( us02_n834 ) );
  AOI221_X1 us02_U168 (.A( us02_n482 ) , .ZN( us02_n487 ) , .B1( us02_n830 ) , .C2( us02_n843 ) , .C1( us02_n851 ) , .B2( us02_n861 ) );
  OAI22_X1 us02_U169 (.ZN( us02_n482 ) , .A1( us02_n707 ) , .B2( us02_n784 ) , .A2( us02_n805 ) , .B1( us02_n811 ) );
  INV_X1 us02_U17 (.A( us02_n748 ) , .ZN( us02_n862 ) );
  INV_X1 us02_U170 (.A( us02_n789 ) , .ZN( us02_n831 ) );
  NAND2_X1 us02_U171 (.A1( us02_n450 ) , .A2( us02_n452 ) , .ZN( us02_n761 ) );
  OAI221_X1 us02_U172 (.A( us02_n726 ) , .C2( us02_n727 ) , .B2( us02_n728 ) , .B1( us02_n729 ) , .ZN( us02_n736 ) , .C1( us02_n816 ) );
  AOI22_X1 us02_U173 (.ZN( us02_n726 ) , .B1( us02_n831 ) , .A2( us02_n837 ) , .A1( us02_n862 ) , .B2( us02_n865 ) );
  INV_X1 us02_U174 (.A( us02_n785 ) , .ZN( us02_n861 ) );
  OAI22_X1 us02_U175 (.ZN( us02_n709 ) , .A2( us02_n727 ) , .B2( us02_n728 ) , .A1( us02_n743 ) , .B1( us02_n812 ) );
  INV_X1 us02_U176 (.A( us02_n815 ) , .ZN( us02_n830 ) );
  OAI22_X1 us02_U177 (.ZN( us02_n488 ) , .A1( us02_n723 ) , .B2( us02_n727 ) , .B1( us02_n729 ) , .A2( us02_n778 ) );
  OAI22_X1 us02_U178 (.ZN( us02_n623 ) , .B1( us02_n668 ) , .B2( us02_n746 ) , .A1( us02_n814 ) , .A2( us02_n815 ) );
  INV_X1 us02_U179 (.A( us02_n743 ) , .ZN( us02_n836 ) );
  AOI222_X1 us02_U18 (.ZN( us02_n604 ) , .B2( us02_n670 ) , .B1( us02_n752 ) , .C2( us02_n830 ) , .A1( us02_n832 ) , .A2( us02_n861 ) , .C1( us02_n862 ) );
  OAI22_X1 us02_U180 (.A1( us02_n723 ) , .ZN( us02_n725 ) , .B2( us02_n749 ) , .B1( us02_n811 ) , .A2( us02_n815 ) );
  OAI22_X1 us02_U181 (.B2( us02_n778 ) , .B1( us02_n779 ) , .ZN( us02_n780 ) , .A2( us02_n813 ) , .A1( us02_n814 ) );
  INV_X1 us02_U182 (.A( us02_n787 ) , .ZN( us02_n844 ) );
  INV_X1 us02_U183 (.A( us02_n804 ) , .ZN( us02_n859 ) );
  INV_X1 us02_U184 (.A( us02_n813 ) , .ZN( us02_n832 ) );
  OAI22_X1 us02_U185 (.B2( us02_n743 ) , .ZN( us02_n745 ) , .A2( us02_n761 ) , .B1( us02_n779 ) , .A1( us02_n791 ) );
  OAI22_X1 us02_U186 (.B2( us02_n802 ) , .B1( us02_n803 ) , .A2( us02_n804 ) , .A1( us02_n805 ) , .ZN( us02_n807 ) );
  OAI22_X1 us02_U187 (.ZN( us02_n495 ) , .A2( us02_n743 ) , .A1( us02_n779 ) , .B1( us02_n790 ) , .B2( us02_n805 ) );
  OAI22_X1 us02_U188 (.ZN( us02_n589 ) , .B1( us02_n729 ) , .B2( us02_n748 ) , .A2( us02_n785 ) , .A1( us02_n802 ) );
  OAI22_X1 us02_U189 (.ZN( us02_n694 ) , .A2( us02_n729 ) , .A1( us02_n779 ) , .B1( us02_n790 ) , .B2( us02_n816 ) );
  AOI222_X1 us02_U19 (.ZN( us02_n562 ) , .B1( us02_n829 ) , .C1( us02_n840 ) , .A2( us02_n842 ) , .A1( us02_n853 ) , .B2( us02_n862 ) , .C2( us02_n872 ) );
  INV_X1 us02_U190 (.A( us02_n802 ) , .ZN( us02_n842 ) );
  INV_X1 us02_U191 (.A( us02_n668 ) , .ZN( us02_n864 ) );
  OAI22_X1 us02_U192 (.ZN( us02_n636 ) , .A1( us02_n698 ) , .B2( us02_n727 ) , .A2( us02_n761 ) , .B1( us02_n815 ) );
  NOR2_X1 us02_U193 (.ZN( us02_n714 ) , .A1( us02_n804 ) , .A2( us02_n816 ) );
  NOR2_X1 us02_U194 (.A1( us02_n696 ) , .ZN( us02_n769 ) , .A2( us02_n814 ) );
  NOR2_X1 us02_U195 (.ZN( us02_n665 ) , .A1( us02_n727 ) , .A2( us02_n802 ) );
  NOR2_X1 us02_U196 (.ZN( us02_n593 ) , .A2( us02_n696 ) , .A1( us02_n727 ) );
  NOR2_X1 us02_U197 (.ZN( us02_n569 ) , .A1( us02_n727 ) , .A2( us02_n805 ) );
  NOR2_X1 us02_U198 (.A2( us02_n743 ) , .ZN( us02_n754 ) , .A1( us02_n804 ) );
  NOR2_X1 us02_U199 (.ZN( us02_n717 ) , .A2( us02_n723 ) , .A1( us02_n743 ) );
  AOI222_X1 us02_U20 (.ZN( us02_n659 ) , .A2( us02_n838 ) , .B1( us02_n840 ) , .C2( us02_n844 ) , .A1( us02_n859 ) , .C1( us02_n862 ) , .B2( us02_n869 ) );
  NOR2_X1 us02_U200 (.ZN( us02_n734 ) , .A2( us02_n802 ) , .A1( us02_n804 ) );
  NOR2_X1 us02_U201 (.ZN( us02_n545 ) , .A2( us02_n779 ) , .A1( us02_n813 ) );
  NOR2_X1 us02_U202 (.ZN( us02_n576 ) , .A2( us02_n698 ) , .A1( us02_n813 ) );
  NOR2_X1 us02_U203 (.ZN( us02_n653 ) , .A1( us02_n727 ) , .A2( us02_n812 ) );
  NOR2_X1 us02_U204 (.ZN( us02_n611 ) , .A1( us02_n778 ) , .A2( us02_n785 ) );
  INV_X1 us02_U205 (.A( us02_n749 ) , .ZN( us02_n841 ) );
  NOR2_X1 us02_U206 (.ZN( us02_n531 ) , .A2( us02_n748 ) , .A1( us02_n749 ) );
  NOR2_X1 us02_U207 (.ZN( us02_n628 ) , .A2( us02_n727 ) , .A1( us02_n784 ) );
  NOR2_X1 us02_U208 (.ZN( us02_n614 ) , .A1( us02_n784 ) , .A2( us02_n814 ) );
  NOR2_X1 us02_U209 (.ZN( us02_n600 ) , .A2( us02_n779 ) , .A1( us02_n802 ) );
  INV_X1 us02_U21 (.A( us02_n646 ) , .ZN( us02_n869 ) );
  NOR2_X1 us02_U210 (.ZN( us02_n610 ) , .A2( us02_n779 ) , .A1( us02_n805 ) );
  INV_X1 us02_U211 (.A( us02_n746 ) , .ZN( us02_n833 ) );
  NOR2_X1 us02_U212 (.A2( us02_n743 ) , .ZN( us02_n768 ) , .A1( us02_n811 ) );
  NOR2_X1 us02_U213 (.ZN( us02_n527 ) , .A2( us02_n723 ) , .A1( us02_n802 ) );
  NOR2_X1 us02_U214 (.ZN( us02_n530 ) , .A2( us02_n779 ) , .A1( us02_n815 ) );
  NOR2_X1 us02_U215 (.ZN( us02_n627 ) , .A2( us02_n668 ) , .A1( us02_n784 ) );
  NOR2_X1 us02_U216 (.ZN( us02_n598 ) , .A2( us02_n790 ) , .A1( us02_n815 ) );
  INV_X1 us02_U217 (.A( us02_n727 ) , .ZN( us02_n851 ) );
  NOR2_X1 us02_U218 (.ZN( us02_n651 ) , .A1( us02_n668 ) , .A2( us02_n813 ) );
  NOR2_X1 us02_U219 (.A1( us02_n668 ) , .ZN( us02_n672 ) , .A2( us02_n743 ) );
  NOR4_X1 us02_U22 (.ZN( us02_n472 ) , .A2( us02_n520 ) , .A4( us02_n593 ) , .A1( us02_n608 ) , .A3( us02_n628 ) );
  NOR2_X1 us02_U220 (.ZN( us02_n601 ) , .A1( us02_n668 ) , .A2( us02_n802 ) );
  NOR2_X1 us02_U221 (.A1( us02_n668 ) , .ZN( us02_n687 ) , .A2( us02_n815 ) );
  INV_X1 us02_U222 (.A( us02_n791 ) , .ZN( us02_n850 ) );
  NOR2_X1 us02_U223 (.A2( us02_n707 ) , .A1( us02_n749 ) , .ZN( us02_n770 ) );
  NOR2_X1 us02_U224 (.A1( us02_n668 ) , .ZN( us02_n765 ) , .A2( us02_n812 ) );
  NOR2_X1 us02_U225 (.A1( us02_n698 ) , .ZN( us02_n767 ) , .A2( us02_n812 ) );
  NOR2_X1 us02_U226 (.ZN( us02_n540 ) , .A2( us02_n696 ) , .A1( us02_n698 ) );
  NOR2_X1 us02_U227 (.ZN( us02_n526 ) , .A1( us02_n668 ) , .A2( us02_n778 ) );
  NOR2_X1 us02_U228 (.ZN( us02_n666 ) , .A1( us02_n749 ) , .A2( us02_n814 ) );
  NOR2_X1 us02_U229 (.ZN( us02_n554 ) , .A1( us02_n749 ) , .A2( us02_n790 ) );
  NOR4_X1 us02_U23 (.ZN( us02_n478 ) , .A1( us02_n519 ) , .A4( us02_n556 ) , .A3( us02_n581 ) , .A2( us02_n629 ) );
  NOR2_X1 us02_U230 (.ZN( us02_n507 ) , .A2( us02_n779 ) , .A1( us02_n784 ) );
  NOR2_X1 us02_U231 (.ZN( us02_n542 ) , .A2( us02_n707 ) , .A1( us02_n784 ) );
  NOR2_X1 us02_U232 (.ZN( us02_n663 ) , .A1( us02_n784 ) , .A2( us02_n790 ) );
  NOR2_X1 us02_U233 (.A2( us02_n696 ) , .ZN( us02_n715 ) , .A1( us02_n791 ) );
  NOR2_X1 us02_U234 (.ZN( us02_n506 ) , .A1( us02_n811 ) , .A2( us02_n816 ) );
  NOR2_X1 us02_U235 (.ZN( us02_n555 ) , .A1( us02_n761 ) , .A2( us02_n804 ) );
  NOR2_X1 us02_U236 (.ZN( us02_n660 ) , .A1( us02_n728 ) , .A2( us02_n789 ) );
  NOR2_X1 us02_U237 (.ZN( us02_n661 ) , .A2( us02_n696 ) , .A1( us02_n728 ) );
  NOR2_X1 us02_U238 (.ZN( us02_n556 ) , .A1( us02_n791 ) , .A2( us02_n813 ) );
  NOR2_X1 us02_U239 (.ZN( us02_n544 ) , .A1( us02_n748 ) , .A2( us02_n813 ) );
  NOR4_X1 us02_U24 (.A4( us02_n531 ) , .A3( us02_n532 ) , .A2( us02_n533 ) , .ZN( us02_n534 ) , .A1( us02_n819 ) );
  NOR2_X1 us02_U240 (.ZN( us02_n508 ) , .A1( us02_n728 ) , .A2( us02_n778 ) );
  NOR2_X1 us02_U241 (.A2( us02_n696 ) , .A1( us02_n779 ) , .ZN( us02_n819 ) );
  OAI22_X1 us02_U242 (.B2( us02_n749 ) , .B1( us02_n750 ) , .A1( us02_n751 ) , .ZN( us02_n755 ) , .A2( us02_n805 ) );
  NOR2_X1 us02_U243 (.ZN( us02_n750 ) , .A2( us02_n851 ) , .A1( us02_n859 ) );
  NOR3_X1 us02_U244 (.ZN( us02_n751 ) , .A2( us02_n852 ) , .A1( us02_n862 ) , .A3( us02_n864 ) );
  NOR2_X1 us02_U245 (.ZN( us02_n529 ) , .A2( us02_n743 ) , .A1( us02_n791 ) );
  NOR2_X1 us02_U246 (.A1( us02_n748 ) , .ZN( us02_n766 ) , .A2( us02_n802 ) );
  NOR2_X1 us02_U247 (.ZN( us02_n543 ) , .A2( us02_n784 ) , .A1( us02_n791 ) );
  NOR2_X1 us02_U248 (.ZN( us02_n662 ) , .A1( us02_n728 ) , .A2( us02_n784 ) );
  NOR2_X1 us02_U249 (.ZN( us02_n630 ) , .A1( us02_n723 ) , .A2( us02_n812 ) );
  NOR4_X1 us02_U25 (.ZN( us02_n455 ) , .A2( us02_n516 ) , .A1( us02_n542 ) , .A3( us02_n578 ) , .A4( us02_n614 ) );
  NOR2_X1 us02_U250 (.ZN( us02_n613 ) , .A1( us02_n761 ) , .A2( us02_n811 ) );
  OAI22_X1 us02_U251 (.B1( us02_n439 ) , .ZN( us02_n443 ) , .A2( us02_n727 ) , .A1( us02_n743 ) , .B2( us02_n748 ) );
  NOR3_X1 us02_U252 (.ZN( us02_n439 ) , .A2( us02_n835 ) , .A3( us02_n836 ) , .A1( us02_n845 ) );
  NOR2_X1 us02_U253 (.ZN( us02_n505 ) , .A2( us02_n727 ) , .A1( us02_n761 ) );
  NOR2_X1 us02_U254 (.ZN( us02_n515 ) , .A1( us02_n707 ) , .A2( us02_n743 ) );
  NOR2_X1 us02_U255 (.ZN( us02_n716 ) , .A2( us02_n743 ) , .A1( us02_n785 ) );
  NOR2_X1 us02_U256 (.ZN( us02_n553 ) , .A1( us02_n785 ) , .A2( us02_n812 ) );
  NOR2_X1 us02_U257 (.ZN( us02_n516 ) , .A1( us02_n707 ) , .A2( us02_n802 ) );
  NOR2_X1 us02_U258 (.ZN( us02_n557 ) , .A1( us02_n707 ) , .A2( us02_n815 ) );
  NOR2_X1 us02_U259 (.ZN( us02_n669 ) , .A1( us02_n789 ) , .A2( us02_n804 ) );
  NOR4_X1 us02_U26 (.A4( us02_n540 ) , .A3( us02_n541 ) , .A2( us02_n542 ) , .ZN( us02_n549 ) , .A1( us02_n687 ) );
  NOR2_X1 us02_U260 (.ZN( us02_n520 ) , .A1( us02_n789 ) , .A2( us02_n811 ) );
  NOR2_X1 us02_U261 (.ZN( us02_n629 ) , .A1( us02_n746 ) , .A2( us02_n814 ) );
  INV_X1 us02_U262 (.A( us02_n805 ) , .ZN( us02_n840 ) );
  AOI21_X1 us02_U263 (.ZN( us02_n570 ) , .B2( us02_n696 ) , .B1( us02_n805 ) , .A( us02_n811 ) );
  NOR2_X1 us02_U264 (.ZN( us02_n654 ) , .A1( us02_n789 ) , .A2( us02_n814 ) );
  INV_X1 us02_U265 (.A( us02_n762 ) , .ZN( us02_n865 ) );
  AOI21_X1 us02_U266 (.ZN( us02_n551 ) , .B1( us02_n668 ) , .A( us02_n696 ) , .B2( us02_n804 ) );
  NOR2_X1 us02_U267 (.ZN( us02_n667 ) , .A2( us02_n707 ) , .A1( us02_n789 ) );
  NOR2_X1 us02_U268 (.ZN( us02_n655 ) , .A1( us02_n746 ) , .A2( us02_n779 ) );
  NOR2_X1 us02_U269 (.ZN( us02_n541 ) , .A1( us02_n761 ) , .A2( us02_n790 ) );
  NOR2_X1 us02_U27 (.ZN( us02_n679 ) , .A2( us02_n833 ) , .A1( us02_n838 ) );
  NOR2_X1 us02_U270 (.ZN( us02_n700 ) , .A2( us02_n785 ) , .A1( us02_n816 ) );
  NOR2_X1 us02_U271 (.ZN( us02_n608 ) , .A2( us02_n723 ) , .A1( us02_n816 ) );
  NOR2_X1 us02_U272 (.A1( us02_n729 ) , .ZN( us02_n764 ) , .A2( us02_n785 ) );
  AOI21_X1 us02_U273 (.A( us02_n814 ) , .B2( us02_n815 ) , .B1( us02_n816 ) , .ZN( us02_n817 ) );
  INV_X1 us02_U274 (.A( us02_n728 ) , .ZN( us02_n867 ) );
  NOR2_X1 us02_U275 (.ZN( us02_n578 ) , .A2( us02_n707 ) , .A1( us02_n729 ) );
  NOR2_X1 us02_U276 (.ZN( us02_n532 ) , .A2( us02_n723 ) , .A1( us02_n729 ) );
  AOI21_X1 us02_U277 (.B1( us02_n624 ) , .ZN( us02_n626 ) , .A( us02_n762 ) , .B2( us02_n813 ) );
  AOI21_X1 us02_U278 (.A( us02_n811 ) , .B2( us02_n812 ) , .B1( us02_n813 ) , .ZN( us02_n818 ) );
  AOI21_X1 us02_U279 (.ZN( us02_n514 ) , .A( us02_n728 ) , .B1( us02_n749 ) , .B2( us02_n802 ) );
  AOI222_X1 us02_U28 (.ZN( us02_n468 ) , .B1( us02_n831 ) , .A1( us02_n838 ) , .C1( us02_n841 ) , .C2( us02_n850 ) , .A2( us02_n854 ) , .B2( us02_n864 ) );
  AOI21_X1 us02_U280 (.ZN( us02_n498 ) , .B1( us02_n679 ) , .A( us02_n811 ) , .B2( us02_n815 ) );
  AOI21_X1 us02_U281 (.ZN( us02_n649 ) , .A( us02_n778 ) , .B1( us02_n791 ) , .B2( us02_n804 ) );
  AOI21_X1 us02_U282 (.ZN( us02_n477 ) , .B2( us02_n696 ) , .A( us02_n748 ) , .B1( us02_n778 ) );
  NOR2_X1 us02_U283 (.ZN( us02_n581 ) , .A1( us02_n743 ) , .A2( us02_n814 ) );
  AOI21_X1 us02_U284 (.ZN( us02_n592 ) , .B1( us02_n749 ) , .A( us02_n791 ) , .B2( us02_n812 ) );
  NOR2_X1 us02_U285 (.A2( us02_n707 ) , .A1( us02_n761 ) , .ZN( us02_n793 ) );
  AOI21_X1 us02_U286 (.ZN( us02_n625 ) , .B2( us02_n668 ) , .A( us02_n789 ) , .B1( us02_n790 ) );
  NOR2_X1 us02_U287 (.ZN( us02_n519 ) , .A2( us02_n707 ) , .A1( us02_n813 ) );
  AOI21_X1 us02_U288 (.ZN( us02_n476 ) , .A( us02_n668 ) , .B1( us02_n749 ) , .B2( us02_n805 ) );
  NOR2_X1 us02_U289 (.ZN( us02_n558 ) , .A2( us02_n790 ) , .A1( us02_n802 ) );
  NOR4_X1 us02_U29 (.A1( us02_n465 ) , .ZN( us02_n466 ) , .A4( us02_n541 ) , .A2( us02_n553 ) , .A3( us02_n613 ) );
  NOR2_X1 us02_U290 (.ZN( us02_n518 ) , .A2( us02_n698 ) , .A1( us02_n815 ) );
  NOR2_X1 us02_U291 (.ZN( us02_n682 ) , .A2( us02_n698 ) , .A1( us02_n802 ) );
  NOR2_X1 us02_U292 (.ZN( us02_n652 ) , .A1( us02_n761 ) , .A2( us02_n785 ) );
  INV_X1 us02_U293 (.A( us02_n812 ) , .ZN( us02_n835 ) );
  AOI21_X1 us02_U294 (.ZN( us02_n509 ) , .B2( us02_n668 ) , .A( us02_n729 ) , .B1( us02_n814 ) );
  AOI21_X1 us02_U295 (.ZN( us02_n538 ) , .B2( us02_n811 ) , .A( us02_n813 ) , .B1( us02_n814 ) );
  AOI21_X1 us02_U296 (.ZN( us02_n539 ) , .A( us02_n762 ) , .B2( us02_n778 ) , .B1( us02_n816 ) );
  NOR2_X1 us02_U297 (.ZN( us02_n580 ) , .A1( us02_n668 ) , .A2( us02_n787 ) );
  AOI21_X1 us02_U298 (.ZN( us02_n588 ) , .B2( us02_n698 ) , .B1( us02_n814 ) , .A( us02_n816 ) );
  AOI21_X1 us02_U299 (.B1( us02_n698 ) , .ZN( us02_n699 ) , .A( us02_n731 ) , .B2( us02_n762 ) );
  NAND2_X1 us02_U3 (.A1( us02_n440 ) , .A2( us02_n463 ) , .ZN( us02_n707 ) );
  AOI221_X1 us02_U30 (.ZN( us02_n467 ) , .C2( us02_n713 ) , .B2( us02_n830 ) , .C1( us02_n844 ) , .B1( us02_n859 ) , .A( us02_n863 ) );
  AOI21_X1 us02_U300 (.ZN( us02_n590 ) , .B2( us02_n762 ) , .A( us02_n784 ) , .B1( us02_n811 ) );
  AOI21_X1 us02_U301 (.ZN( us02_n497 ) , .A( us02_n723 ) , .B2( us02_n761 ) , .B1( us02_n813 ) );
  NOR2_X1 us02_U302 (.ZN( us02_n546 ) , .A1( us02_n698 ) , .A2( us02_n743 ) );
  INV_X1 us02_U303 (.A( us02_n790 ) , .ZN( us02_n872 ) );
  INV_X1 us02_U304 (.A( us02_n811 ) , .ZN( us02_n853 ) );
  AOI21_X1 us02_U305 (.ZN( us02_n648 ) , .B1( us02_n728 ) , .B2( us02_n762 ) , .A( us02_n812 ) );
  NOR2_X1 us02_U306 (.ZN( us02_n684 ) , .A1( us02_n728 ) , .A2( us02_n815 ) );
  AOI21_X1 us02_U307 (.B1( us02_n685 ) , .ZN( us02_n686 ) , .A( us02_n727 ) , .B2( us02_n760 ) );
  AOI21_X1 us02_U308 (.ZN( us02_n568 ) , .B1( us02_n749 ) , .B2( us02_n761 ) , .A( us02_n779 ) );
  AOI21_X1 us02_U309 (.ZN( us02_n499 ) , .A( us02_n696 ) , .B1( us02_n707 ) , .B2( us02_n785 ) );
  NOR4_X1 us02_U31 (.A4( us02_n513 ) , .A3( us02_n514 ) , .A2( us02_n515 ) , .A1( us02_n516 ) , .ZN( us02_n523 ) );
  NOR2_X1 us02_U310 (.ZN( us02_n567 ) , .A1( us02_n728 ) , .A2( us02_n761 ) );
  NOR2_X1 us02_U311 (.ZN( us02_n579 ) , .A2( us02_n696 ) , .A1( us02_n790 ) );
  NOR2_X1 us02_U312 (.ZN( us02_n565 ) , .A2( us02_n696 ) , .A1( us02_n762 ) );
  AOI21_X1 us02_U313 (.ZN( us02_n513 ) , .A( us02_n778 ) , .B2( us02_n791 ) , .B1( us02_n811 ) );
  INV_X1 us02_U314 (.A( us02_n698 ) , .ZN( us02_n852 ) );
  NOR2_X1 us02_U315 (.ZN( us02_n664 ) , .A1( us02_n779 ) , .A2( us02_n812 ) );
  AOI21_X1 us02_U316 (.ZN( us02_n449 ) , .B2( us02_n791 ) , .A( us02_n802 ) , .B1( us02_n814 ) );
  NOR2_X1 us02_U317 (.ZN( us02_n631 ) , .A2( us02_n696 ) , .A1( us02_n723 ) );
  AOI21_X1 us02_U318 (.ZN( us02_n563 ) , .B1( us02_n723 ) , .A( us02_n778 ) , .B2( us02_n790 ) );
  AOI21_X1 us02_U319 (.ZN( us02_n496 ) , .A( us02_n778 ) , .B2( us02_n790 ) , .B1( us02_n803 ) );
  AOI222_X1 us02_U32 (.ZN( us02_n524 ) , .A1( us02_n833 ) , .B2( us02_n836 ) , .C1( us02_n843 ) , .C2( us02_n849 ) , .A2( us02_n851 ) , .B1( us02_n865 ) );
  NAND2_X1 us02_U320 (.ZN( us02_n752 ) , .A1( us02_n762 ) , .A2( us02_n804 ) );
  NOR2_X1 us02_U321 (.ZN( us02_n528 ) , .A1( us02_n707 ) , .A2( us02_n778 ) );
  NOR2_X1 us02_U322 (.ZN( us02_n577 ) , .A1( us02_n707 ) , .A2( us02_n812 ) );
  AOI21_X1 us02_U323 (.ZN( us02_n688 ) , .B2( us02_n748 ) , .B1( us02_n762 ) , .A( us02_n805 ) );
  NOR2_X1 us02_U324 (.ZN( us02_n566 ) , .A1( us02_n746 ) , .A2( us02_n804 ) );
  NOR2_X1 us02_U325 (.ZN( us02_n683 ) , .A1( us02_n790 ) , .A2( us02_n812 ) );
  NOR2_X1 us02_U326 (.A2( us02_n812 ) , .A1( us02_n814 ) , .ZN( us02_n820 ) );
  AOI21_X1 us02_U327 (.A( us02_n789 ) , .B2( us02_n790 ) , .B1( us02_n791 ) , .ZN( us02_n792 ) );
  AOI21_X1 us02_U328 (.A( us02_n732 ) , .ZN( us02_n733 ) , .B2( us02_n779 ) , .B1( us02_n791 ) );
  NOR2_X1 us02_U329 (.ZN( us02_n710 ) , .A1( us02_n761 ) , .A2( us02_n762 ) );
  NOR4_X1 us02_U33 (.A3( us02_n520 ) , .A1( us02_n521 ) , .ZN( us02_n522 ) , .A2( us02_n672 ) , .A4( us02_n768 ) );
  NOR2_X1 us02_U330 (.ZN( us02_n582 ) , .A1( us02_n791 ) , .A2( us02_n816 ) );
  NOR2_X1 us02_U331 (.ZN( us02_n533 ) , .A1( us02_n723 ) , .A2( us02_n787 ) );
  NOR2_X1 us02_U332 (.ZN( us02_n681 ) , .A2( us02_n707 ) , .A1( us02_n816 ) );
  INV_X1 us02_U333 (.A( us02_n696 ) , .ZN( us02_n837 ) );
  NOR2_X1 us02_U334 (.ZN( us02_n641 ) , .A2( us02_n787 ) , .A1( us02_n790 ) );
  INV_X1 us02_U335 (.A( us02_n814 ) , .ZN( us02_n854 ) );
  AOI21_X1 us02_U336 (.ZN( us02_n441 ) , .A( us02_n698 ) , .B1( us02_n732 ) , .B2( us02_n749 ) );
  INV_X1 us02_U337 (.A( us02_n779 ) , .ZN( us02_n849 ) );
  AOI22_X1 us02_U338 (.A2( us02_n781 ) , .ZN( us02_n782 ) , .B2( us02_n830 ) , .A1( us02_n833 ) , .B1( us02_n862 ) );
  NAND2_X1 us02_U339 (.ZN( us02_n670 ) , .A1( us02_n805 ) , .A2( us02_n815 ) );
  NOR4_X1 us02_U34 (.A3( us02_n754 ) , .A2( us02_n755 ) , .A1( us02_n756 ) , .ZN( us02_n757 ) , .A4( us02_n868 ) );
  NAND2_X1 us02_U340 (.ZN( us02_n713 ) , .A1( us02_n727 ) , .A2( us02_n779 ) );
  NAND2_X1 us02_U341 (.A2( us02_n761 ) , .A1( us02_n805 ) , .ZN( us02_n809 ) );
  AOI21_X1 us02_U342 (.ZN( us02_n442 ) , .B1( us02_n788 ) , .B2( us02_n790 ) , .A( us02_n813 ) );
  NOR2_X1 us02_U343 (.ZN( us02_n483 ) , .A1( us02_n787 ) , .A2( us02_n804 ) );
  NOR2_X1 us02_U344 (.ZN( us02_n469 ) , .A2( us02_n778 ) , .A1( us02_n814 ) );
  INV_X1 us02_U345 (.A( us02_n784 ) , .ZN( us02_n845 ) );
  OAI21_X1 us02_U346 (.A( us02_n786 ) , .B2( us02_n787 ) , .B1( us02_n788 ) , .ZN( us02_n794 ) );
  OAI21_X1 us02_U347 (.ZN( us02_n786 ) , .A( us02_n838 ) , .B1( us02_n862 ) , .B2( us02_n872 ) );
  NOR2_X1 us02_U348 (.ZN( us02_n711 ) , .A2( us02_n723 ) , .A1( us02_n789 ) );
  NOR2_X1 us02_U349 (.ZN( us02_n525 ) , .A1( us02_n723 ) , .A2( us02_n749 ) );
  AOI211_X1 us02_U35 (.B( us02_n744 ) , .A( us02_n745 ) , .ZN( us02_n758 ) , .C1( us02_n831 ) , .C2( us02_n852 ) );
  NAND2_X1 us02_U350 (.A1( us02_n698 ) , .A2( us02_n728 ) , .ZN( us02_n781 ) );
  AOI21_X1 us02_U351 (.ZN( us02_n638 ) , .B2( us02_n748 ) , .A( us02_n787 ) , .B1( us02_n811 ) );
  AOI21_X1 us02_U352 (.ZN( us02_n639 ) , .B2( us02_n746 ) , .A( us02_n791 ) , .B1( us02_n802 ) );
  AOI21_X1 us02_U353 (.ZN( us02_n640 ) , .B1( us02_n679 ) , .A( us02_n790 ) , .B2( us02_n816 ) );
  NOR2_X1 us02_U354 (.ZN( us02_n517 ) , .A1( us02_n707 ) , .A2( us02_n787 ) );
  OAI21_X1 us02_U355 (.A( us02_n697 ) , .ZN( us02_n701 ) , .B2( us02_n749 ) , .B1( us02_n803 ) );
  OAI21_X1 us02_U356 (.ZN( us02_n697 ) , .B2( us02_n832 ) , .B1( us02_n837 ) , .A( us02_n859 ) );
  OAI21_X1 us02_U357 (.A( us02_n730 ) , .B1( us02_n731 ) , .ZN( us02_n735 ) , .B2( us02_n804 ) );
  OAI21_X1 us02_U358 (.ZN( us02_n730 ) , .A( us02_n832 ) , .B2( us02_n851 ) , .B1( us02_n872 ) );
  NAND2_X1 us02_U359 (.A2( us02_n748 ) , .A1( us02_n785 ) , .ZN( us02_n808 ) );
  NOR3_X1 us02_U36 (.A3( us02_n740 ) , .A2( us02_n741 ) , .A1( us02_n742 ) , .ZN( us02_n759 ) );
  INV_X1 us02_U360 (.A( us02_n816 ) , .ZN( us02_n843 ) );
  INV_X1 us02_U361 (.A( us02_n723 ) , .ZN( us02_n855 ) );
  AND2_X1 us02_U362 (.ZN( us02_n731 ) , .A1( us02_n778 ) , .A2( us02_n784 ) );
  NAND2_X1 us02_U363 (.A1( us02_n446 ) , .A2( us02_n448 ) , .ZN( us02_n804 ) );
  NAND2_X1 us02_U364 (.A1( us02_n454 ) , .A2( us02_n470 ) , .ZN( us02_n802 ) );
  NAND2_X1 us02_U365 (.A1( us02_n450 ) , .A2( us02_n453 ) , .ZN( us02_n813 ) );
  NAND2_X1 us02_U366 (.A1( us02_n450 ) , .A2( us02_n470 ) , .ZN( us02_n815 ) );
  NAND2_X1 us02_U367 (.A1( us02_n453 ) , .A2( us02_n460 ) , .ZN( us02_n812 ) );
  NAND2_X1 us02_U368 (.A1( us02_n452 ) , .A2( us02_n460 ) , .ZN( us02_n743 ) );
  NAND2_X1 us02_U369 (.A1( us02_n451 ) , .A2( us02_n464 ) , .ZN( us02_n668 ) );
  NOR4_X1 us02_U37 (.A4( us02_n733 ) , .A3( us02_n734 ) , .A2( us02_n735 ) , .A1( us02_n736 ) , .ZN( us02_n737 ) );
  NAND2_X1 us02_U370 (.A2( us02_n447 ) , .A1( us02_n459 ) , .ZN( us02_n727 ) );
  NAND2_X1 us02_U371 (.A1( us02_n454 ) , .A2( us02_n461 ) , .ZN( us02_n749 ) );
  NAND2_X1 us02_U372 (.A2( us02_n452 ) , .A1( us02_n454 ) , .ZN( us02_n805 ) );
  NAND2_X1 us02_U373 (.A2( us02_n453 ) , .A1( us02_n471 ) , .ZN( us02_n778 ) );
  NAND2_X1 us02_U374 (.A1( us02_n452 ) , .A2( us02_n471 ) , .ZN( us02_n784 ) );
  NAND2_X1 us02_U375 (.A2( us02_n463 ) , .A1( us02_n464 ) , .ZN( us02_n811 ) );
  NAND2_X1 us02_U376 (.A1( us02_n440 ) , .A2( us02_n459 ) , .ZN( us02_n698 ) );
  NAND2_X1 us02_U377 (.A2( us02_n448 ) , .A1( us02_n451 ) , .ZN( us02_n762 ) );
  NAND2_X1 us02_U378 (.A2( us02_n447 ) , .A1( us02_n451 ) , .ZN( us02_n728 ) );
  NAND2_X1 us02_U379 (.A2( us02_n460 ) , .A1( us02_n461 ) , .ZN( us02_n746 ) );
  AOI211_X1 us02_U38 (.B( us02_n724 ) , .A( us02_n725 ) , .ZN( us02_n738 ) , .C1( us02_n842 ) , .C2( us02_n854 ) );
  NAND2_X2 us02_U380 (.A2( us02_n460 ) , .A1( us02_n470 ) , .ZN( us02_n696 ) );
  NAND2_X1 us02_U381 (.A1( us02_n461 ) , .A2( us02_n471 ) , .ZN( us02_n787 ) );
  NOR2_X1 us02_U382 (.ZN( us02_n464 ) , .A2( us02_n846 ) , .A1( us02_n847 ) );
  NOR2_X1 us02_U383 (.ZN( us02_n452 ) , .A1( us02_n825 ) , .A2( us02_n826 ) );
  NOR2_X1 us02_U384 (.ZN( us02_n450 ) , .A1( us02_n827 ) , .A2( us02_n828 ) );
  NOR2_X1 us02_U385 (.ZN( us02_n446 ) , .A2( us02_n848 ) , .A1( us02_n857 ) );
  NAND2_X1 us02_U386 (.A2( us02_n453 ) , .A1( us02_n454 ) , .ZN( us02_n729 ) );
  NAND2_X1 us02_U387 (.A1( us02_n450 ) , .A2( us02_n461 ) , .ZN( us02_n789 ) );
  NAND2_X2 us02_U388 (.A2( us02_n447 ) , .A1( us02_n463 ) , .ZN( us02_n814 ) );
  NAND2_X2 us02_U389 (.A2( us02_n440 ) , .A1( us02_n451 ) , .ZN( us02_n790 ) );
  NOR3_X1 us02_U39 (.A3( us02_n721 ) , .A1( us02_n722 ) , .ZN( us02_n739 ) , .A2( us02_n740 ) );
  NAND2_X2 us02_U390 (.A1( us02_n448 ) , .A2( us02_n463 ) , .ZN( us02_n723 ) );
  NAND2_X1 us02_U391 (.A2( us02_n440 ) , .A1( us02_n446 ) , .ZN( us02_n783 ) );
  NAND2_X2 us02_U392 (.A1( us02_n448 ) , .A2( us02_n459 ) , .ZN( us02_n791 ) );
  NAND2_X2 us02_U393 (.A2( us02_n459 ) , .A1( us02_n464 ) , .ZN( us02_n779 ) );
  NAND2_X1 us02_U394 (.A1( us02_n446 ) , .A2( us02_n447 ) , .ZN( us02_n785 ) );
  NOR2_X1 us02_U395 (.A2( sa02_6 ) , .A1( sa02_7 ) , .ZN( us02_n463 ) );
  NOR2_X1 us02_U396 (.A2( sa02_5 ) , .ZN( us02_n447 ) , .A1( us02_n846 ) );
  NOR2_X1 us02_U397 (.A2( sa02_7 ) , .ZN( us02_n459 ) , .A1( us02_n848 ) );
  NOR2_X1 us02_U398 (.A2( sa02_4 ) , .ZN( us02_n448 ) , .A1( us02_n847 ) );
  NOR2_X1 us02_U399 (.A2( sa02_4 ) , .A1( sa02_5 ) , .ZN( us02_n440 ) );
  NAND2_X1 us02_U4 (.A2( us02_n470 ) , .A1( us02_n471 ) , .ZN( us02_n816 ) );
  AOI221_X1 us02_U40 (.A( us02_n780 ) , .ZN( us02_n797 ) , .C2( us02_n836 ) , .B2( us02_n837 ) , .B1( us02_n864 ) , .C1( us02_n865 ) );
  NOR2_X1 us02_U400 (.A2( sa02_1 ) , .ZN( us02_n470 ) , .A1( us02_n825 ) );
  NOR2_X1 us02_U401 (.A2( sa02_2 ) , .A1( sa02_3 ) , .ZN( us02_n471 ) );
  NOR2_X1 us02_U402 (.A2( sa02_6 ) , .ZN( us02_n451 ) , .A1( us02_n857 ) );
  NOR2_X1 us02_U403 (.A2( sa02_2 ) , .ZN( us02_n460 ) , .A1( us02_n828 ) );
  NOR2_X1 us02_U404 (.A2( sa02_0 ) , .ZN( us02_n453 ) , .A1( us02_n826 ) );
  NOR2_X1 us02_U405 (.A2( sa02_0 ) , .A1( sa02_1 ) , .ZN( us02_n461 ) );
  NOR2_X1 us02_U406 (.A2( sa02_3 ) , .ZN( us02_n454 ) , .A1( us02_n827 ) );
  INV_X1 us02_U407 (.A( sa02_6 ) , .ZN( us02_n848 ) );
  INV_X1 us02_U408 (.A( sa02_1 ) , .ZN( us02_n826 ) );
  INV_X1 us02_U409 (.A( sa02_3 ) , .ZN( us02_n828 ) );
  NOR4_X1 us02_U41 (.A4( us02_n792 ) , .A3( us02_n793 ) , .A2( us02_n794 ) , .A1( us02_n795 ) , .ZN( us02_n796 ) );
  INV_X1 us02_U410 (.A( sa02_2 ) , .ZN( us02_n827 ) );
  INV_X1 us02_U411 (.A( sa02_0 ) , .ZN( us02_n825 ) );
  INV_X1 us02_U412 (.A( sa02_5 ) , .ZN( us02_n847 ) );
  INV_X1 us02_U413 (.A( sa02_7 ) , .ZN( us02_n857 ) );
  OAI221_X1 us02_U414 (.A( us02_n782 ) , .C2( us02_n783 ) , .B2( us02_n784 ) , .B1( us02_n785 ) , .ZN( us02_n795 ) , .C1( us02_n812 ) );
  OAI22_X1 us02_U415 (.ZN( us02_n587 ) , .A2( us02_n746 ) , .B2( us02_n761 ) , .A1( us02_n762 ) , .B1( us02_n783 ) );
  AOI21_X1 us02_U416 (.ZN( us02_n591 ) , .B1( us02_n727 ) , .B2( us02_n783 ) , .A( us02_n789 ) );
  OAI221_X1 us02_U417 (.A( us02_n695 ) , .ZN( us02_n702 ) , .C2( us02_n783 ) , .C1( us02_n784 ) , .B1( us02_n785 ) , .B2( us02_n805 ) );
  NAND2_X1 us02_U418 (.A1( us02_n728 ) , .A2( us02_n783 ) , .ZN( us02_n810 ) );
  AOI21_X1 us02_U419 (.ZN( us02_n622 ) , .B1( us02_n698 ) , .A( us02_n778 ) , .B2( us02_n783 ) );
  NOR4_X1 us02_U42 (.A4( us02_n775 ) , .A3( us02_n776 ) , .A1( us02_n777 ) , .ZN( us02_n798 ) , .A2( us02_n800 ) );
  OAI22_X1 us02_U420 (.ZN( us02_n680 ) , .A1( us02_n698 ) , .A2( us02_n729 ) , .B2( us02_n783 ) , .B1( us02_n816 ) );
  AOI21_X1 us02_U421 (.ZN( us02_n647 ) , .A( us02_n761 ) , .B2( us02_n783 ) , .B1( us02_n791 ) );
  OAI21_X1 us02_U422 (.A( us02_n612 ) , .ZN( us02_n615 ) , .B1( us02_n624 ) , .B2( us02_n783 ) );
  NOR2_X1 us02_U423 (.ZN( us02_n650 ) , .A1( us02_n783 ) , .A2( us02_n787 ) );
  NOR2_X1 us02_U424 (.ZN( us02_n552 ) , .A2( us02_n743 ) , .A1( us02_n783 ) );
  NOR2_X1 us02_U425 (.ZN( us02_n609 ) , .A1( us02_n783 ) , .A2( us02_n815 ) );
  OAI222_X1 us02_U426 (.A2( us02_n668 ) , .ZN( us02_n673 ) , .B1( us02_n746 ) , .B2( us02_n783 ) , .C2( us02_n787 ) , .C1( us02_n814 ) , .A1( us02_n816 ) );
  NOR2_X1 us02_U427 (.ZN( us02_n599 ) , .A2( us02_n696 ) , .A1( us02_n783 ) );
  INV_X1 us02_U428 (.A( us02_n783 ) , .ZN( us02_n860 ) );
  AOI221_X1 us02_U429 (.A( us02_n575 ) , .ZN( us02_n586 ) , .B2( us02_n830 ) , .C2( us02_n842 ) , .B1( us02_n853 ) , .C1( us02_n860 ) );
  NOR2_X1 us02_U43 (.ZN( us02_n803 ) , .A1( us02_n853 ) , .A2( us02_n860 ) );
  AOI21_X1 us02_U430 (.ZN( us02_n575 ) , .B2( us02_n723 ) , .B1( us02_n747 ) , .A( us02_n784 ) );
  INV_X1 us02_U431 (.A( sa02_4 ) , .ZN( us02_n846 ) );
  NAND2_X1 us02_U432 (.ZN( sa02_sr_2 ) , .A2( us02_n438 ) , .A1( us02_n644 ) );
  NOR3_X1 us02_U433 (.A2( us02_n606 ) , .A1( us02_n607 ) , .ZN( us02_n645 ) , .A3( us02_n721 ) );
  AOI222_X1 us02_U434 (.B2( us02_n637 ) , .ZN( us02_n643 ) , .B1( us02_n840 ) , .A1( us02_n841 ) , .C2( us02_n845 ) , .C1( us02_n862 ) , .A2( us02_n864 ) );
  NOR4_X1 us02_U435 (.A4( us02_n638 ) , .A3( us02_n639 ) , .A2( us02_n640 ) , .A1( us02_n641 ) , .ZN( us02_n642 ) );
  AOI211_X1 us02_U436 (.A( us02_n636 ) , .ZN( us02_n644 ) , .B( us02_n742 ) , .C2( us02_n838 ) , .C1( us02_n853 ) );
  NAND3_X1 us02_U437 (.ZN( sa02_sr_6 ) , .A3( us02_n796 ) , .A2( us02_n797 ) , .A1( us02_n798 ) );
  NAND3_X1 us02_U438 (.ZN( sa02_sr_5 ) , .A3( us02_n757 ) , .A2( us02_n758 ) , .A1( us02_n759 ) );
  NAND3_X1 us02_U439 (.ZN( sa02_sr_4 ) , .A3( us02_n737 ) , .A2( us02_n738 ) , .A1( us02_n739 ) );
  NAND4_X1 us02_U44 (.ZN( sa02_sr_3 ) , .A4( us02_n703 ) , .A3( us02_n704 ) , .A2( us02_n705 ) , .A1( us02_n706 ) );
  NAND3_X1 us02_U440 (.A3( us02_n674 ) , .A2( us02_n675 ) , .A1( us02_n676 ) , .ZN( us02_n806 ) );
  NAND3_X1 us02_U441 (.ZN( us02_n637 ) , .A3( us02_n707 ) , .A2( us02_n723 ) , .A1( us02_n791 ) );
  NAND3_X1 us02_U442 (.A3( us02_n617 ) , .A2( us02_n618 ) , .A1( us02_n619 ) , .ZN( us02_n724 ) );
  NAND3_X1 us02_U443 (.A3( us02_n584 ) , .A2( us02_n585 ) , .A1( us02_n586 ) , .ZN( us02_n620 ) );
  NAND3_X1 us02_U444 (.ZN( us02_n564 ) , .A3( us02_n679 ) , .A2( us02_n749 ) , .A1( us02_n784 ) );
  NAND3_X1 us02_U445 (.A3( us02_n522 ) , .A2( us02_n523 ) , .A1( us02_n524 ) , .ZN( us02_n741 ) );
  NAND3_X1 us02_U446 (.A3( us02_n511 ) , .A1( us02_n512 ) , .ZN( us02_n607 ) , .A2( us02_n870 ) );
  NAND3_X1 us02_U447 (.A3( us02_n466 ) , .A2( us02_n467 ) , .A1( us02_n468 ) , .ZN( us02_n776 ) );
  NAND4_X1 us02_U448 (.A4( us02_n632 ) , .A3( us02_n633 ) , .A2( us02_n634 ) , .A1( us02_n635 ) , .ZN( us02_n742 ) );
  NOR4_X1 us02_U45 (.A4( us02_n699 ) , .A3( us02_n700 ) , .A2( us02_n701 ) , .A1( us02_n702 ) , .ZN( us02_n703 ) );
  AOI211_X1 us02_U46 (.B( us02_n693 ) , .A( us02_n694 ) , .ZN( us02_n704 ) , .C2( us02_n830 ) , .C1( us02_n850 ) );
  NOR2_X1 us02_U47 (.ZN( us02_n706 ) , .A2( us02_n775 ) , .A1( us02_n799 ) );
  NAND4_X1 us02_U48 (.ZN( sa02_sr_7 ) , .A4( us02_n821 ) , .A3( us02_n822 ) , .A2( us02_n823 ) , .A1( us02_n824 ) );
  NOR4_X1 us02_U49 (.A4( us02_n817 ) , .A3( us02_n818 ) , .A2( us02_n819 ) , .A1( us02_n820 ) , .ZN( us02_n821 ) );
  NOR3_X1 us02_U5 (.ZN( us02_n597 ) , .A1( us02_n607 ) , .A3( us02_n722 ) , .A2( us02_n741 ) );
  AOI222_X1 us02_U50 (.C2( us02_n808 ) , .B2( us02_n809 ) , .A2( us02_n810 ) , .ZN( us02_n822 ) , .C1( us02_n831 ) , .A1( us02_n838 ) , .B1( us02_n852 ) );
  AOI211_X1 us02_U51 (.B( us02_n806 ) , .A( us02_n807 ) , .ZN( us02_n823 ) , .C1( us02_n841 ) , .C2( us02_n849 ) );
  NOR2_X1 us02_U52 (.ZN( us02_n747 ) , .A1( us02_n860 ) , .A2( us02_n861 ) );
  NAND4_X1 us02_U53 (.ZN( sa02_sr_0 ) , .A4( us02_n500 ) , .A3( us02_n501 ) , .A2( us02_n502 ) , .A1( us02_n503 ) );
  AOI221_X1 us02_U54 (.A( us02_n496 ) , .ZN( us02_n501 ) , .B2( us02_n842 ) , .C1( us02_n845 ) , .C2( us02_n859 ) , .B1( us02_n861 ) );
  NOR4_X1 us02_U55 (.A4( us02_n497 ) , .A3( us02_n498 ) , .A2( us02_n499 ) , .ZN( us02_n500 ) , .A1( us02_n526 ) );
  AOI211_X1 us02_U56 (.A( us02_n495 ) , .ZN( us02_n502 ) , .B( us02_n801 ) , .C2( us02_n838 ) , .C1( us02_n850 ) );
  NAND4_X1 us02_U57 (.ZN( sa02_sr_1 ) , .A4( us02_n594 ) , .A3( us02_n595 ) , .A2( us02_n596 ) , .A1( us02_n597 ) );
  NOR4_X1 us02_U58 (.A4( us02_n590 ) , .A3( us02_n591 ) , .A2( us02_n592 ) , .A1( us02_n593 ) , .ZN( us02_n594 ) );
  AOI211_X1 us02_U59 (.B( us02_n588 ) , .A( us02_n589 ) , .ZN( us02_n595 ) , .C2( us02_n810 ) , .C1( us02_n832 ) );
  NOR3_X1 us02_U6 (.A3( us02_n799 ) , .A2( us02_n800 ) , .A1( us02_n801 ) , .ZN( us02_n824 ) );
  AOI211_X1 us02_U60 (.A( us02_n587 ) , .ZN( us02_n596 ) , .B( us02_n620 ) , .C1( us02_n844 ) , .C2( us02_n854 ) );
  NOR2_X1 us02_U61 (.ZN( us02_n624 ) , .A2( us02_n835 ) , .A1( us02_n838 ) );
  AND3_X1 us02_U62 (.ZN( us02_n438 ) , .A2( us02_n642 ) , .A3( us02_n643 ) , .A1( us02_n645 ) );
  NOR4_X1 us02_U63 (.A4( us02_n576 ) , .A3( us02_n577 ) , .A2( us02_n578 ) , .ZN( us02_n585 ) , .A1( us02_n682 ) );
  NOR4_X1 us02_U64 (.A1( us02_n583 ) , .ZN( us02_n584 ) , .A3( us02_n651 ) , .A2( us02_n661 ) , .A4( us02_n766 ) );
  AOI211_X1 us02_U65 (.B( us02_n622 ) , .A( us02_n623 ) , .ZN( us02_n634 ) , .C2( us02_n835 ) , .C1( us02_n862 ) );
  NOR4_X1 us02_U66 (.A4( us02_n628 ) , .A3( us02_n629 ) , .A2( us02_n630 ) , .A1( us02_n631 ) , .ZN( us02_n632 ) );
  NOR4_X1 us02_U67 (.A4( us02_n625 ) , .A3( us02_n626 ) , .A2( us02_n627 ) , .ZN( us02_n633 ) , .A1( us02_n663 ) );
  NAND4_X1 us02_U68 (.A4( us02_n656 ) , .A3( us02_n657 ) , .A2( us02_n658 ) , .A1( us02_n659 ) , .ZN( us02_n799 ) );
  NOR3_X1 us02_U69 (.A3( us02_n647 ) , .A2( us02_n648 ) , .A1( us02_n649 ) , .ZN( us02_n658 ) );
  NOR3_X1 us02_U7 (.ZN( us02_n503 ) , .A2( us02_n678 ) , .A3( us02_n776 ) , .A1( us02_n875 ) );
  NOR3_X1 us02_U70 (.A3( us02_n650 ) , .A2( us02_n651 ) , .A1( us02_n652 ) , .ZN( us02_n657 ) );
  NOR3_X1 us02_U71 (.A3( us02_n653 ) , .A2( us02_n654 ) , .A1( us02_n655 ) , .ZN( us02_n656 ) );
  NAND4_X1 us02_U72 (.A4( us02_n771 ) , .A3( us02_n772 ) , .A2( us02_n773 ) , .A1( us02_n774 ) , .ZN( us02_n800 ) );
  NOR3_X1 us02_U73 (.A3( us02_n764 ) , .A2( us02_n765 ) , .A1( us02_n766 ) , .ZN( us02_n772 ) );
  NOR4_X1 us02_U74 (.A4( us02_n767 ) , .A3( us02_n768 ) , .A2( us02_n769 ) , .A1( us02_n770 ) , .ZN( us02_n771 ) );
  AOI222_X1 us02_U75 (.ZN( us02_n774 ) , .A1( us02_n829 ) , .C1( us02_n833 ) , .B2( us02_n840 ) , .A2( us02_n849 ) , .B1( us02_n860 ) , .C2( us02_n872 ) );
  NOR4_X1 us02_U76 (.A4( us02_n664 ) , .A3( us02_n665 ) , .A2( us02_n666 ) , .A1( us02_n667 ) , .ZN( us02_n675 ) );
  NOR4_X1 us02_U77 (.A4( us02_n660 ) , .A3( us02_n661 ) , .A2( us02_n662 ) , .A1( us02_n663 ) , .ZN( us02_n676 ) );
  NOR4_X1 us02_U78 (.A3( us02_n672 ) , .A1( us02_n673 ) , .ZN( us02_n674 ) , .A4( us02_n714 ) , .A2( us02_n858 ) );
  NOR2_X1 us02_U79 (.ZN( us02_n760 ) , .A1( us02_n832 ) , .A2( us02_n833 ) );
  INV_X1 us02_U8 (.A( us02_n705 ) , .ZN( us02_n875 ) );
  NAND4_X1 us02_U80 (.A4( us02_n455 ) , .A3( us02_n456 ) , .A2( us02_n457 ) , .A1( us02_n458 ) , .ZN( us02_n678 ) );
  NOR3_X1 us02_U81 (.ZN( us02_n456 ) , .A3( us02_n529 ) , .A1( us02_n554 ) , .A2( us02_n569 ) );
  AOI221_X1 us02_U82 (.A( us02_n449 ) , .ZN( us02_n458 ) , .C2( us02_n752 ) , .B1( us02_n831 ) , .C1( us02_n841 ) , .B2( us02_n860 ) );
  NOR4_X1 us02_U83 (.ZN( us02_n457 ) , .A2( us02_n508 ) , .A1( us02_n598 ) , .A4( us02_n627 ) , .A3( us02_n710 ) );
  NAND4_X1 us02_U84 (.A4( us02_n602 ) , .A3( us02_n603 ) , .A2( us02_n604 ) , .A1( us02_n605 ) , .ZN( us02_n721 ) );
  NOR3_X1 us02_U85 (.A1( us02_n598 ) , .ZN( us02_n603 ) , .A3( us02_n662 ) , .A2( us02_n769 ) );
  NOR4_X1 us02_U86 (.A3( us02_n599 ) , .A2( us02_n600 ) , .A1( us02_n601 ) , .ZN( us02_n602 ) , .A4( us02_n654 ) );
  AOI222_X1 us02_U87 (.ZN( us02_n605 ) , .A1( us02_n829 ) , .C2( us02_n836 ) , .B1( us02_n841 ) , .A2( us02_n855 ) , .B2( us02_n860 ) , .C1( us02_n867 ) );
  NAND4_X1 us02_U88 (.A4( us02_n534 ) , .A3( us02_n535 ) , .A2( us02_n536 ) , .A1( us02_n537 ) , .ZN( us02_n621 ) );
  NOR4_X1 us02_U89 (.A4( us02_n525 ) , .A2( us02_n526 ) , .A1( us02_n527 ) , .ZN( us02_n537 ) , .A3( us02_n700 ) );
  NOR3_X1 us02_U9 (.A3( us02_n620 ) , .A2( us02_n621 ) , .ZN( us02_n635 ) , .A1( us02_n724 ) );
  NOR4_X1 us02_U90 (.A1( us02_n530 ) , .ZN( us02_n535 ) , .A2( us02_n653 ) , .A4( us02_n667 ) , .A3( us02_n764 ) );
  NOR4_X1 us02_U91 (.A4( us02_n528 ) , .A3( us02_n529 ) , .ZN( us02_n536 ) , .A2( us02_n683 ) , .A1( us02_n793 ) );
  NAND4_X1 us02_U92 (.A4( us02_n547 ) , .A3( us02_n548 ) , .A2( us02_n549 ) , .A1( us02_n550 ) , .ZN( us02_n744 ) );
  NOR3_X1 us02_U93 (.ZN( us02_n548 ) , .A2( us02_n650 ) , .A1( us02_n666 ) , .A3( us02_n770 ) );
  AOI211_X1 us02_U94 (.B( us02_n538 ) , .A( us02_n539 ) , .ZN( us02_n550 ) , .C2( us02_n838 ) , .C1( us02_n850 ) );
  NOR4_X1 us02_U95 (.A4( us02_n543 ) , .A3( us02_n544 ) , .A2( us02_n545 ) , .A1( us02_n546 ) , .ZN( us02_n547 ) );
  NAND4_X1 us02_U96 (.A4( us02_n478 ) , .A3( us02_n479 ) , .A2( us02_n480 ) , .A1( us02_n481 ) , .ZN( us02_n693 ) );
  NOR3_X1 us02_U97 (.ZN( us02_n479 ) , .A2( us02_n507 ) , .A3( us02_n600 ) , .A1( us02_n609 ) );
  AOI211_X1 us02_U98 (.B( us02_n476 ) , .A( us02_n477 ) , .ZN( us02_n481 ) , .C2( us02_n832 ) , .C1( us02_n860 ) );
  NOR4_X1 us02_U99 (.ZN( us02_n480 ) , .A3( us02_n531 ) , .A4( us02_n544 ) , .A2( us02_n566 ) , .A1( us02_n716 ) );
  NOR3_X1 us21_U10 (.A3( us21_n619 ) , .A2( us21_n620 ) , .ZN( us21_n634 ) , .A1( us21_n723 ) );
  NOR4_X1 us21_U100 (.A4( us21_n524 ) , .A2( us21_n525 ) , .A1( us21_n526 ) , .ZN( us21_n536 ) , .A3( us21_n699 ) );
  NOR4_X1 us21_U101 (.A1( us21_n529 ) , .ZN( us21_n534 ) , .A2( us21_n652 ) , .A4( us21_n666 ) , .A3( us21_n763 ) );
  NOR4_X1 us21_U102 (.A4( us21_n527 ) , .A3( us21_n528 ) , .ZN( us21_n535 ) , .A2( us21_n682 ) , .A1( us21_n792 ) );
  NAND4_X1 us21_U103 (.A4( us21_n546 ) , .A3( us21_n547 ) , .A2( us21_n548 ) , .A1( us21_n549 ) , .ZN( us21_n743 ) );
  NOR3_X1 us21_U104 (.ZN( us21_n547 ) , .A2( us21_n649 ) , .A1( us21_n665 ) , .A3( us21_n769 ) );
  AOI211_X1 us21_U105 (.B( us21_n537 ) , .A( us21_n538 ) , .ZN( us21_n549 ) , .C2( us21_n837 ) , .C1( us21_n849 ) );
  NOR4_X1 us21_U106 (.A4( us21_n539 ) , .A3( us21_n540 ) , .A2( us21_n541 ) , .ZN( us21_n548 ) , .A1( us21_n686 ) );
  NAND4_X1 us21_U107 (.A4( us21_n477 ) , .A3( us21_n478 ) , .A2( us21_n479 ) , .A1( us21_n480 ) , .ZN( us21_n692 ) );
  NOR3_X1 us21_U108 (.ZN( us21_n478 ) , .A2( us21_n506 ) , .A3( us21_n599 ) , .A1( us21_n608 ) );
  AOI211_X1 us21_U109 (.B( us21_n475 ) , .A( us21_n476 ) , .ZN( us21_n480 ) , .C2( us21_n831 ) , .C1( us21_n859 ) );
  NOR2_X1 us21_U11 (.ZN( us21_n493 ) , .A1( us21_n676 ) , .A2( us21_n692 ) );
  NOR4_X1 us21_U110 (.ZN( us21_n479 ) , .A3( us21_n530 ) , .A4( us21_n543 ) , .A2( us21_n565 ) , .A1( us21_n715 ) );
  NOR4_X1 us21_U111 (.A4( us21_n607 ) , .A3( us21_n608 ) , .A2( us21_n609 ) , .A1( us21_n610 ) , .ZN( us21_n617 ) );
  NOR4_X1 us21_U112 (.ZN( us21_n618 ) , .A1( us21_n654 ) , .A3( us21_n664 ) , .A4( us21_n680 ) , .A2( us21_n764 ) );
  NOR4_X1 us21_U113 (.A4( us21_n612 ) , .A3( us21_n613 ) , .A2( us21_n614 ) , .A1( us21_n615 ) , .ZN( us21_n616 ) );
  NOR2_X1 us21_U114 (.ZN( us21_n684 ) , .A1( us21_n829 ) , .A2( us21_n830 ) );
  NAND4_X1 us21_U115 (.A4( us21_n471 ) , .A3( us21_n472 ) , .A2( us21_n473 ) , .A1( us21_n474 ) , .ZN( us21_n676 ) );
  NOR4_X1 us21_U116 (.A4( us21_n468 ) , .ZN( us21_n474 ) , .A3( us21_n554 ) , .A1( us21_n733 ) , .A2( us21_n753 ) );
  NOR4_X1 us21_U117 (.ZN( us21_n473 ) , .A1( us21_n529 ) , .A3( us21_n566 ) , .A4( us21_n598 ) , .A2( us21_n640 ) );
  NOR4_X1 us21_U118 (.ZN( us21_n472 ) , .A1( us21_n504 ) , .A3( us21_n542 ) , .A2( us21_n581 ) , .A4( us21_n714 ) );
  NAND4_X1 us21_U119 (.A4( us21_n689 ) , .A3( us21_n690 ) , .A1( us21_n691 ) , .ZN( us21_n774 ) , .A2( us21_n870 ) );
  NOR2_X1 us21_U12 (.A1( us21_n676 ) , .ZN( us21_n691 ) , .A2( us21_n805 ) );
  INV_X1 us21_U120 (.A( us21_n677 ) , .ZN( us21_n870 ) );
  AOI221_X1 us21_U121 (.A( us21_n679 ) , .ZN( us21_n690 ) , .B2( us21_n838 ) , .C1( us21_n840 ) , .C2( us21_n860 ) , .B1( us21_n863 ) );
  NOR4_X1 us21_U122 (.A4( us21_n685 ) , .A3( us21_n686 ) , .A2( us21_n687 ) , .A1( us21_n688 ) , .ZN( us21_n689 ) );
  NOR2_X1 us21_U123 (.ZN( us21_n731 ) , .A2( us21_n830 ) , .A1( us21_n843 ) );
  NAND4_X1 us21_U124 (.A4( us21_n717 ) , .A3( us21_n718 ) , .A2( us21_n719 ) , .ZN( us21_n739 ) , .A1( us21_n855 ) );
  INV_X1 us21_U125 (.A( us21_n707 ) , .ZN( us21_n855 ) );
  NOR4_X1 us21_U126 (.A4( us21_n713 ) , .A3( us21_n714 ) , .A2( us21_n715 ) , .A1( us21_n716 ) , .ZN( us21_n717 ) );
  AOI221_X1 us21_U127 (.A( us21_n708 ) , .ZN( us21_n719 ) , .C2( us21_n842 ) , .B2( us21_n843 ) , .C1( us21_n859 ) , .B1( us21_n860 ) );
  NAND4_X1 us21_U128 (.A4( us21_n571 ) , .A3( us21_n572 ) , .A1( us21_n573 ) , .ZN( us21_n721 ) , .A2( us21_n872 ) );
  NOR4_X1 us21_U129 (.A4( us21_n567 ) , .A3( us21_n568 ) , .A2( us21_n569 ) , .A1( us21_n570 ) , .ZN( us21_n571 ) );
  INV_X1 us21_U13 (.A( us21_n605 ) , .ZN( us21_n872 ) );
  AOI221_X1 us21_U130 (.A( us21_n562 ) , .C2( us21_n563 ) , .ZN( us21_n572 ) , .B2( us21_n843 ) , .B1( us21_n850 ) , .C1( us21_n851 ) );
  NOR2_X1 us21_U131 (.ZN( us21_n573 ) , .A1( us21_n620 ) , .A2( us21_n743 ) );
  NAND4_X1 us21_U132 (.A4( us21_n491 ) , .A3( us21_n492 ) , .A1( us21_n493 ) , .ZN( us21_n800 ) , .A2( us21_n865 ) );
  AOI221_X1 us21_U133 (.A( us21_n487 ) , .ZN( us21_n492 ) , .B2( us21_n834 ) , .C2( us21_n839 ) , .C1( us21_n849 ) , .B1( us21_n858 ) );
  INV_X1 us21_U134 (.A( us21_n776 ) , .ZN( us21_n865 ) );
  NOR4_X1 us21_U135 (.A2( us21_n489 ) , .A1( us21_n490 ) , .ZN( us21_n491 ) , .A3( us21_n578 ) , .A4( us21_n610 ) );
  INV_X1 us21_U136 (.A( us21_n760 ) , .ZN( us21_n828 ) );
  NOR2_X1 us21_U137 (.ZN( us21_n645 ) , .A1( us21_n852 ) , .A2( us21_n866 ) );
  INV_X1 us21_U138 (.A( us21_n461 ) , .ZN( us21_n862 ) );
  OAI21_X1 us21_U139 (.ZN( us21_n461 ) , .B1( us21_n807 ) , .A( us21_n832 ) , .B2( us21_n849 ) );
  INV_X1 us21_U14 (.A( us21_n678 ) , .ZN( us21_n838 ) );
  OR4_X1 us21_U140 (.ZN( us21_n490 ) , .A4( us21_n532 ) , .A2( us21_n545 ) , .A1( us21_n557 ) , .A3( us21_n630 ) );
  OR4_X1 us21_U141 (.A4( us21_n564 ) , .A3( us21_n565 ) , .A2( us21_n566 ) , .ZN( us21_n570 ) , .A1( us21_n663 ) );
  OR4_X1 us21_U142 (.A4( us21_n680 ) , .A3( us21_n681 ) , .A2( us21_n682 ) , .A1( us21_n683 ) , .ZN( us21_n688 ) );
  OR4_X1 us21_U143 (.ZN( us21_n464 ) , .A4( us21_n516 ) , .A3( us21_n527 ) , .A2( us21_n576 ) , .A1( us21_n710 ) );
  OR4_X1 us21_U144 (.A4( us21_n516 ) , .A2( us21_n517 ) , .A1( us21_n518 ) , .ZN( us21_n520 ) , .A3( us21_n819 ) );
  OR4_X1 us21_U145 (.A4( us21_n578 ) , .A3( us21_n579 ) , .A2( us21_n580 ) , .A1( us21_n581 ) , .ZN( us21_n582 ) );
  NAND2_X1 us21_U146 (.ZN( us21_n611 ) , .A2( us21_n835 ) , .A1( us21_n871 ) );
  OR3_X1 us21_U147 (.A3( us21_n504 ) , .A2( us21_n505 ) , .A1( us21_n506 ) , .ZN( us21_n509 ) );
  AOI221_X1 us21_U148 (.A( us21_n711 ) , .B2( us21_n712 ) , .ZN( us21_n718 ) , .C1( us21_n830 ) , .B1( us21_n837 ) , .C2( us21_n861 ) );
  OR2_X1 us21_U149 (.A2( us21_n709 ) , .A1( us21_n710 ) , .ZN( us21_n711 ) );
  NOR4_X1 us21_U15 (.A4( us21_n443 ) , .A3( us21_n444 ) , .A2( us21_n514 ) , .A1( us21_n539 ) , .ZN( us21_n704 ) );
  INV_X1 us21_U150 (.A( us21_n752 ) , .ZN( us21_n867 ) );
  OAI21_X1 us21_U151 (.B1( us21_n751 ) , .ZN( us21_n752 ) , .A( us21_n843 ) , .B2( us21_n866 ) );
  INV_X1 us21_U152 (.A( us21_n670 ) , .ZN( us21_n857 ) );
  AOI21_X1 us21_U153 (.A( us21_n668 ) , .B1( us21_n669 ) , .ZN( us21_n670 ) , .B2( us21_n854 ) );
  AOI222_X1 us21_U154 (.ZN( us21_n658 ) , .A2( us21_n837 ) , .B1( us21_n839 ) , .C2( us21_n843 ) , .A1( us21_n858 ) , .C1( us21_n861 ) , .B2( us21_n868 ) );
  INV_X1 us21_U155 (.A( us21_n645 ) , .ZN( us21_n868 ) );
  OAI22_X1 us21_U156 (.ZN( us21_n481 ) , .A1( us21_n706 ) , .B2( us21_n783 ) , .A2( us21_n804 ) , .B1( us21_n810 ) );
  OAI22_X1 us21_U157 (.ZN( us21_n635 ) , .A1( us21_n697 ) , .B2( us21_n726 ) , .A2( us21_n760 ) , .B1( us21_n814 ) );
  OAI222_X1 us21_U158 (.B2( us21_n706 ) , .ZN( us21_n707 ) , .C2( us21_n722 ) , .B1( us21_n745 ) , .A1( us21_n804 ) , .C1( us21_n812 ) , .A2( us21_n813 ) );
  NAND2_X1 us21_U159 (.A1( us21_n445 ) , .A2( us21_n463 ) , .ZN( us21_n747 ) );
  OR3_X1 us21_U16 (.ZN( us21_n444 ) , .A1( us21_n526 ) , .A3( us21_n575 ) , .A2( us21_n873 ) );
  AOI22_X1 us21_U160 (.ZN( us21_n694 ) , .A1( us21_n828 ) , .B2( us21_n841 ) , .A2( us21_n863 ) , .B1( us21_n866 ) );
  INV_X1 us21_U161 (.A( us21_n728 ) , .ZN( us21_n837 ) );
  NAND2_X1 us21_U162 (.A1( us21_n449 ) , .A2( us21_n451 ) , .ZN( us21_n760 ) );
  INV_X1 us21_U163 (.A( us21_n788 ) , .ZN( us21_n830 ) );
  OAI221_X1 us21_U164 (.A( us21_n725 ) , .C2( us21_n726 ) , .B2( us21_n727 ) , .B1( us21_n728 ) , .ZN( us21_n735 ) , .C1( us21_n815 ) );
  AOI22_X1 us21_U165 (.ZN( us21_n725 ) , .B1( us21_n830 ) , .A2( us21_n836 ) , .A1( us21_n861 ) , .B2( us21_n864 ) );
  AND2_X1 us21_U166 (.ZN( us21_n746 ) , .A1( us21_n782 ) , .A2( us21_n784 ) );
  OAI22_X1 us21_U167 (.ZN( us21_n487 ) , .A1( us21_n722 ) , .B2( us21_n726 ) , .B1( us21_n728 ) , .A2( us21_n777 ) );
  OAI22_X1 us21_U168 (.ZN( us21_n622 ) , .B1( us21_n667 ) , .B2( us21_n745 ) , .A1( us21_n813 ) , .A2( us21_n814 ) );
  OAI22_X1 us21_U169 (.B2( us21_n777 ) , .B1( us21_n778 ) , .ZN( us21_n779 ) , .A2( us21_n812 ) , .A1( us21_n813 ) );
  OR4_X1 us21_U17 (.A4( us21_n440 ) , .A2( us21_n441 ) , .A1( us21_n442 ) , .ZN( us21_n443 ) , .A3( us21_n551 ) );
  OAI22_X1 us21_U170 (.A1( us21_n722 ) , .ZN( us21_n724 ) , .B2( us21_n748 ) , .B1( us21_n810 ) , .A2( us21_n814 ) );
  OAI22_X1 us21_U171 (.B2( us21_n742 ) , .ZN( us21_n744 ) , .A2( us21_n760 ) , .B1( us21_n778 ) , .A1( us21_n790 ) );
  OAI22_X1 us21_U172 (.B2( us21_n801 ) , .B1( us21_n802 ) , .A2( us21_n803 ) , .A1( us21_n804 ) , .ZN( us21_n806 ) );
  OAI22_X1 us21_U173 (.ZN( us21_n494 ) , .A2( us21_n742 ) , .A1( us21_n778 ) , .B1( us21_n789 ) , .B2( us21_n804 ) );
  INV_X1 us21_U174 (.A( us21_n742 ) , .ZN( us21_n835 ) );
  INV_X1 us21_U175 (.A( us21_n786 ) , .ZN( us21_n843 ) );
  INV_X1 us21_U176 (.A( us21_n814 ) , .ZN( us21_n829 ) );
  OAI22_X1 us21_U177 (.B1( us21_n488 ) , .ZN( us21_n489 ) , .A1( us21_n684 ) , .A2( us21_n761 ) , .B2( us21_n815 ) );
  NOR3_X1 us21_U178 (.ZN( us21_n488 ) , .A1( us21_n780 ) , .A2( us21_n848 ) , .A3( us21_n861 ) );
  OAI22_X1 us21_U179 (.ZN( us21_n588 ) , .B1( us21_n728 ) , .B2( us21_n747 ) , .A2( us21_n784 ) , .A1( us21_n801 ) );
  INV_X1 us21_U18 (.A( us21_n611 ) , .ZN( us21_n873 ) );
  OAI22_X1 us21_U180 (.ZN( us21_n693 ) , .A2( us21_n728 ) , .A1( us21_n778 ) , .B1( us21_n789 ) , .B2( us21_n815 ) );
  OAI22_X1 us21_U181 (.ZN( us21_n708 ) , .A2( us21_n726 ) , .B2( us21_n727 ) , .A1( us21_n742 ) , .B1( us21_n811 ) );
  INV_X1 us21_U182 (.A( us21_n812 ) , .ZN( us21_n831 ) );
  INV_X1 us21_U183 (.A( us21_n667 ) , .ZN( us21_n863 ) );
  NOR2_X1 us21_U184 (.ZN( us21_n716 ) , .A2( us21_n722 ) , .A1( us21_n742 ) );
  NOR2_X1 us21_U185 (.ZN( us21_n664 ) , .A1( us21_n726 ) , .A2( us21_n801 ) );
  NOR2_X1 us21_U186 (.ZN( us21_n568 ) , .A1( us21_n726 ) , .A2( us21_n804 ) );
  NOR2_X1 us21_U187 (.ZN( us21_n544 ) , .A2( us21_n778 ) , .A1( us21_n812 ) );
  INV_X1 us21_U188 (.A( us21_n748 ) , .ZN( us21_n840 ) );
  NOR2_X1 us21_U189 (.ZN( us21_n530 ) , .A2( us21_n747 ) , .A1( us21_n748 ) );
  INV_X1 us21_U19 (.A( us21_n747 ) , .ZN( us21_n861 ) );
  NOR2_X1 us21_U190 (.ZN( us21_n575 ) , .A2( us21_n697 ) , .A1( us21_n812 ) );
  NOR2_X1 us21_U191 (.ZN( us21_n652 ) , .A1( us21_n726 ) , .A2( us21_n811 ) );
  NOR2_X1 us21_U192 (.ZN( us21_n613 ) , .A1( us21_n783 ) , .A2( us21_n813 ) );
  NOR2_X1 us21_U193 (.ZN( us21_n627 ) , .A2( us21_n726 ) , .A1( us21_n783 ) );
  NOR2_X1 us21_U194 (.ZN( us21_n599 ) , .A2( us21_n778 ) , .A1( us21_n801 ) );
  NOR2_X1 us21_U195 (.ZN( us21_n610 ) , .A1( us21_n777 ) , .A2( us21_n784 ) );
  NOR2_X1 us21_U196 (.ZN( us21_n526 ) , .A2( us21_n722 ) , .A1( us21_n801 ) );
  NOR2_X1 us21_U197 (.ZN( us21_n626 ) , .A2( us21_n667 ) , .A1( us21_n783 ) );
  INV_X1 us21_U198 (.A( us21_n790 ) , .ZN( us21_n849 ) );
  NOR2_X1 us21_U199 (.A2( us21_n742 ) , .ZN( us21_n767 ) , .A1( us21_n810 ) );
  AOI222_X1 us21_U20 (.ZN( us21_n561 ) , .B1( us21_n828 ) , .C1( us21_n839 ) , .A2( us21_n841 ) , .A1( us21_n852 ) , .B2( us21_n861 ) , .C2( us21_n871 ) );
  NOR2_X1 us21_U200 (.ZN( us21_n529 ) , .A2( us21_n778 ) , .A1( us21_n814 ) );
  NOR2_X1 us21_U201 (.A2( us21_n706 ) , .A1( us21_n748 ) , .ZN( us21_n769 ) );
  NOR2_X1 us21_U202 (.ZN( us21_n597 ) , .A2( us21_n789 ) , .A1( us21_n814 ) );
  NOR2_X1 us21_U203 (.ZN( us21_n609 ) , .A2( us21_n778 ) , .A1( us21_n804 ) );
  NOR2_X1 us21_U204 (.ZN( us21_n650 ) , .A1( us21_n667 ) , .A2( us21_n812 ) );
  INV_X1 us21_U205 (.A( us21_n745 ) , .ZN( us21_n832 ) );
  NOR2_X1 us21_U206 (.A1( us21_n667 ) , .ZN( us21_n671 ) , .A2( us21_n742 ) );
  NOR2_X1 us21_U207 (.ZN( us21_n600 ) , .A1( us21_n667 ) , .A2( us21_n801 ) );
  NOR2_X1 us21_U208 (.A1( us21_n667 ) , .ZN( us21_n686 ) , .A2( us21_n814 ) );
  NOR2_X1 us21_U209 (.ZN( us21_n665 ) , .A1( us21_n748 ) , .A2( us21_n813 ) );
  NOR4_X1 us21_U21 (.ZN( us21_n471 ) , .A2( us21_n519 ) , .A4( us21_n592 ) , .A1( us21_n607 ) , .A3( us21_n627 ) );
  NOR2_X1 us21_U210 (.ZN( us21_n553 ) , .A1( us21_n748 ) , .A2( us21_n789 ) );
  NOR2_X1 us21_U211 (.ZN( us21_n506 ) , .A2( us21_n778 ) , .A1( us21_n783 ) );
  NOR2_X1 us21_U212 (.ZN( us21_n541 ) , .A2( us21_n706 ) , .A1( us21_n783 ) );
  NOR2_X1 us21_U213 (.ZN( us21_n662 ) , .A1( us21_n783 ) , .A2( us21_n789 ) );
  NOR2_X1 us21_U214 (.A1( us21_n667 ) , .ZN( us21_n764 ) , .A2( us21_n811 ) );
  NOR2_X1 us21_U215 (.A1( us21_n697 ) , .ZN( us21_n766 ) , .A2( us21_n811 ) );
  OAI22_X1 us21_U216 (.B1( us21_n438 ) , .ZN( us21_n442 ) , .A2( us21_n726 ) , .A1( us21_n742 ) , .B2( us21_n747 ) );
  NOR3_X1 us21_U217 (.ZN( us21_n438 ) , .A2( us21_n834 ) , .A3( us21_n835 ) , .A1( us21_n844 ) );
  NOR2_X1 us21_U218 (.ZN( us21_n525 ) , .A1( us21_n667 ) , .A2( us21_n777 ) );
  NOR2_X1 us21_U219 (.ZN( us21_n505 ) , .A1( us21_n810 ) , .A2( us21_n815 ) );
  NOR4_X1 us21_U22 (.A4( us21_n542 ) , .A3( us21_n543 ) , .A2( us21_n544 ) , .A1( us21_n545 ) , .ZN( us21_n546 ) );
  NOR2_X1 us21_U220 (.ZN( us21_n659 ) , .A1( us21_n727 ) , .A2( us21_n788 ) );
  INV_X1 us21_U221 (.A( us21_n801 ) , .ZN( us21_n841 ) );
  NOR2_X1 us21_U222 (.ZN( us21_n555 ) , .A1( us21_n790 ) , .A2( us21_n812 ) );
  NOR2_X1 us21_U223 (.ZN( us21_n543 ) , .A1( us21_n747 ) , .A2( us21_n812 ) );
  NOR2_X1 us21_U224 (.ZN( us21_n507 ) , .A1( us21_n727 ) , .A2( us21_n777 ) );
  NOR2_X1 us21_U225 (.ZN( us21_n528 ) , .A2( us21_n742 ) , .A1( us21_n790 ) );
  NOR2_X1 us21_U226 (.A1( us21_n747 ) , .ZN( us21_n765 ) , .A2( us21_n801 ) );
  NOR2_X1 us21_U227 (.A2( us21_n742 ) , .ZN( us21_n753 ) , .A1( us21_n803 ) );
  OAI22_X1 us21_U228 (.B2( us21_n748 ) , .B1( us21_n749 ) , .A1( us21_n750 ) , .ZN( us21_n754 ) , .A2( us21_n804 ) );
  NOR2_X1 us21_U229 (.ZN( us21_n749 ) , .A2( us21_n850 ) , .A1( us21_n858 ) );
  NOR4_X1 us21_U23 (.ZN( us21_n477 ) , .A1( us21_n518 ) , .A4( us21_n555 ) , .A3( us21_n580 ) , .A2( us21_n628 ) );
  NOR3_X1 us21_U230 (.ZN( us21_n750 ) , .A2( us21_n851 ) , .A1( us21_n861 ) , .A3( us21_n863 ) );
  NOR2_X1 us21_U231 (.ZN( us21_n542 ) , .A2( us21_n783 ) , .A1( us21_n790 ) );
  INV_X1 us21_U232 (.A( us21_n804 ) , .ZN( us21_n839 ) );
  NOR2_X1 us21_U233 (.ZN( us21_n629 ) , .A1( us21_n722 ) , .A2( us21_n811 ) );
  NOR2_X1 us21_U234 (.ZN( us21_n733 ) , .A2( us21_n801 ) , .A1( us21_n803 ) );
  NOR2_X1 us21_U235 (.ZN( us21_n514 ) , .A1( us21_n706 ) , .A2( us21_n742 ) );
  NOR2_X1 us21_U236 (.ZN( us21_n661 ) , .A1( us21_n727 ) , .A2( us21_n783 ) );
  NOR2_X1 us21_U237 (.ZN( us21_n715 ) , .A2( us21_n742 ) , .A1( us21_n784 ) );
  NOR2_X1 us21_U238 (.ZN( us21_n612 ) , .A1( us21_n760 ) , .A2( us21_n810 ) );
  INV_X1 us21_U239 (.A( us21_n726 ) , .ZN( us21_n850 ) );
  NOR4_X1 us21_U24 (.ZN( us21_n454 ) , .A2( us21_n515 ) , .A1( us21_n541 ) , .A3( us21_n577 ) , .A4( us21_n613 ) );
  NOR2_X1 us21_U240 (.ZN( us21_n552 ) , .A1( us21_n784 ) , .A2( us21_n811 ) );
  NOR2_X1 us21_U241 (.ZN( us21_n515 ) , .A1( us21_n706 ) , .A2( us21_n801 ) );
  NOR2_X1 us21_U242 (.ZN( us21_n504 ) , .A2( us21_n726 ) , .A1( us21_n760 ) );
  NOR2_X1 us21_U243 (.ZN( us21_n556 ) , .A1( us21_n706 ) , .A2( us21_n814 ) );
  NOR2_X1 us21_U244 (.ZN( us21_n519 ) , .A1( us21_n788 ) , .A2( us21_n810 ) );
  INV_X1 us21_U245 (.A( us21_n803 ) , .ZN( us21_n858 ) );
  NOR2_X1 us21_U246 (.ZN( us21_n713 ) , .A1( us21_n803 ) , .A2( us21_n815 ) );
  NOR2_X1 us21_U247 (.ZN( us21_n653 ) , .A1( us21_n788 ) , .A2( us21_n813 ) );
  NOR2_X1 us21_U248 (.ZN( us21_n666 ) , .A2( us21_n706 ) , .A1( us21_n788 ) );
  NOR2_X1 us21_U249 (.ZN( us21_n628 ) , .A1( us21_n745 ) , .A2( us21_n813 ) );
  NOR4_X1 us21_U25 (.A4( us21_n530 ) , .A3( us21_n531 ) , .A2( us21_n532 ) , .ZN( us21_n533 ) , .A1( us21_n818 ) );
  NOR2_X1 us21_U250 (.ZN( us21_n554 ) , .A1( us21_n760 ) , .A2( us21_n803 ) );
  NOR2_X1 us21_U251 (.ZN( us21_n540 ) , .A1( us21_n760 ) , .A2( us21_n789 ) );
  NOR2_X1 us21_U252 (.ZN( us21_n699 ) , .A2( us21_n784 ) , .A1( us21_n815 ) );
  NOR2_X1 us21_U253 (.A1( us21_n728 ) , .ZN( us21_n763 ) , .A2( us21_n784 ) );
  NOR2_X1 us21_U254 (.ZN( us21_n607 ) , .A2( us21_n722 ) , .A1( us21_n815 ) );
  NOR2_X1 us21_U255 (.ZN( us21_n577 ) , .A2( us21_n706 ) , .A1( us21_n728 ) );
  NOR2_X1 us21_U256 (.ZN( us21_n531 ) , .A2( us21_n722 ) , .A1( us21_n728 ) );
  AOI21_X1 us21_U257 (.A( us21_n810 ) , .B2( us21_n811 ) , .B1( us21_n812 ) , .ZN( us21_n817 ) );
  AOI21_X1 us21_U258 (.ZN( us21_n513 ) , .A( us21_n727 ) , .B1( us21_n748 ) , .B2( us21_n801 ) );
  NOR2_X1 us21_U259 (.ZN( us21_n654 ) , .A1( us21_n745 ) , .A2( us21_n778 ) );
  NOR2_X1 us21_U26 (.ZN( us21_n678 ) , .A2( us21_n832 ) , .A1( us21_n837 ) );
  AOI21_X1 us21_U260 (.A( us21_n813 ) , .B2( us21_n814 ) , .B1( us21_n815 ) , .ZN( us21_n816 ) );
  NOR2_X1 us21_U261 (.ZN( us21_n580 ) , .A1( us21_n742 ) , .A2( us21_n813 ) );
  AOI21_X1 us21_U262 (.ZN( us21_n591 ) , .B1( us21_n748 ) , .A( us21_n790 ) , .B2( us21_n811 ) );
  AOI21_X1 us21_U263 (.B1( us21_n623 ) , .ZN( us21_n625 ) , .A( us21_n761 ) , .B2( us21_n812 ) );
  NOR2_X1 us21_U264 (.A2( us21_n706 ) , .A1( us21_n760 ) , .ZN( us21_n792 ) );
  NOR2_X1 us21_U265 (.ZN( us21_n640 ) , .A2( us21_n786 ) , .A1( us21_n789 ) );
  AOI21_X1 us21_U266 (.ZN( us21_n497 ) , .B1( us21_n678 ) , .A( us21_n810 ) , .B2( us21_n814 ) );
  NOR2_X1 us21_U267 (.ZN( us21_n668 ) , .A1( us21_n788 ) , .A2( us21_n803 ) );
  NOR2_X1 us21_U268 (.ZN( us21_n557 ) , .A2( us21_n789 ) , .A1( us21_n801 ) );
  AOI21_X1 us21_U269 (.ZN( us21_n624 ) , .B2( us21_n667 ) , .A( us21_n788 ) , .B1( us21_n789 ) );
  NOR4_X1 us21_U27 (.A4( us21_n575 ) , .A3( us21_n576 ) , .A2( us21_n577 ) , .ZN( us21_n584 ) , .A1( us21_n681 ) );
  NOR2_X1 us21_U270 (.ZN( us21_n681 ) , .A2( us21_n697 ) , .A1( us21_n801 ) );
  NOR2_X1 us21_U271 (.ZN( us21_n651 ) , .A1( us21_n760 ) , .A2( us21_n784 ) );
  NOR2_X1 us21_U272 (.ZN( us21_n518 ) , .A2( us21_n706 ) , .A1( us21_n812 ) );
  INV_X1 us21_U273 (.A( us21_n811 ) , .ZN( us21_n834 ) );
  NOR2_X1 us21_U274 (.ZN( us21_n517 ) , .A2( us21_n697 ) , .A1( us21_n814 ) );
  AOI21_X1 us21_U275 (.ZN( us21_n475 ) , .A( us21_n667 ) , .B1( us21_n748 ) , .B2( us21_n804 ) );
  AOI21_X1 us21_U276 (.ZN( us21_n508 ) , .B2( us21_n667 ) , .A( us21_n728 ) , .B1( us21_n813 ) );
  AOI21_X1 us21_U277 (.ZN( us21_n537 ) , .B2( us21_n810 ) , .A( us21_n812 ) , .B1( us21_n813 ) );
  INV_X1 us21_U278 (.A( us21_n761 ) , .ZN( us21_n864 ) );
  AOI21_X1 us21_U279 (.ZN( us21_n538 ) , .A( us21_n761 ) , .B2( us21_n777 ) , .B1( us21_n815 ) );
  NOR4_X1 us21_U28 (.A1( us21_n582 ) , .ZN( us21_n583 ) , .A3( us21_n650 ) , .A2( us21_n660 ) , .A4( us21_n765 ) );
  NOR2_X1 us21_U280 (.ZN( us21_n579 ) , .A1( us21_n667 ) , .A2( us21_n786 ) );
  AOI21_X1 us21_U281 (.ZN( us21_n587 ) , .B2( us21_n697 ) , .B1( us21_n813 ) , .A( us21_n815 ) );
  AOI21_X1 us21_U282 (.ZN( us21_n589 ) , .B2( us21_n761 ) , .A( us21_n783 ) , .B1( us21_n810 ) );
  AOI21_X1 us21_U283 (.B1( us21_n697 ) , .ZN( us21_n698 ) , .A( us21_n730 ) , .B2( us21_n761 ) );
  AOI21_X1 us21_U284 (.ZN( us21_n638 ) , .B2( us21_n745 ) , .A( us21_n790 ) , .B1( us21_n801 ) );
  AOI21_X1 us21_U285 (.ZN( us21_n496 ) , .A( us21_n722 ) , .B2( us21_n760 ) , .B1( us21_n812 ) );
  INV_X1 us21_U286 (.A( us21_n789 ) , .ZN( us21_n871 ) );
  NOR2_X1 us21_U287 (.ZN( us21_n545 ) , .A1( us21_n697 ) , .A2( us21_n742 ) );
  INV_X1 us21_U288 (.A( us21_n727 ) , .ZN( us21_n866 ) );
  AOI21_X1 us21_U289 (.ZN( us21_n647 ) , .B1( us21_n727 ) , .B2( us21_n761 ) , .A( us21_n811 ) );
  AOI221_X1 us21_U29 (.A( us21_n779 ) , .ZN( us21_n796 ) , .C2( us21_n835 ) , .B2( us21_n836 ) , .B1( us21_n863 ) , .C1( us21_n864 ) );
  AOI21_X1 us21_U290 (.ZN( us21_n567 ) , .B1( us21_n748 ) , .B2( us21_n760 ) , .A( us21_n778 ) );
  INV_X1 us21_U291 (.A( us21_n810 ) , .ZN( us21_n852 ) );
  NOR2_X1 us21_U292 (.ZN( us21_n683 ) , .A1( us21_n727 ) , .A2( us21_n814 ) );
  AOI21_X1 us21_U293 (.B1( us21_n684 ) , .ZN( us21_n685 ) , .A( us21_n726 ) , .B2( us21_n759 ) );
  NOR2_X1 us21_U294 (.ZN( us21_n566 ) , .A1( us21_n727 ) , .A2( us21_n760 ) );
  NOR2_X1 us21_U295 (.ZN( us21_n663 ) , .A1( us21_n778 ) , .A2( us21_n811 ) );
  AOI21_X1 us21_U296 (.ZN( us21_n448 ) , .B2( us21_n790 ) , .A( us21_n801 ) , .B1( us21_n813 ) );
  AOI21_X1 us21_U297 (.ZN( us21_n512 ) , .A( us21_n777 ) , .B2( us21_n790 ) , .B1( us21_n810 ) );
  AOI21_X1 us21_U298 (.ZN( us21_n637 ) , .B2( us21_n747 ) , .A( us21_n786 ) , .B1( us21_n810 ) );
  INV_X1 us21_U299 (.A( us21_n697 ) , .ZN( us21_n851 ) );
  NAND2_X2 us21_U3 (.A2( us21_n458 ) , .A1( us21_n463 ) , .ZN( us21_n778 ) );
  NOR4_X1 us21_U30 (.A4( us21_n791 ) , .A3( us21_n792 ) , .A2( us21_n793 ) , .A1( us21_n794 ) , .ZN( us21_n795 ) );
  AOI21_X1 us21_U300 (.ZN( us21_n562 ) , .B1( us21_n722 ) , .A( us21_n777 ) , .B2( us21_n789 ) );
  NOR2_X1 us21_U301 (.ZN( us21_n576 ) , .A1( us21_n706 ) , .A2( us21_n811 ) );
  NOR2_X1 us21_U302 (.ZN( us21_n527 ) , .A1( us21_n706 ) , .A2( us21_n777 ) );
  AOI21_X1 us21_U303 (.ZN( us21_n687 ) , .B2( us21_n747 ) , .B1( us21_n761 ) , .A( us21_n804 ) );
  NOR2_X1 us21_U304 (.ZN( us21_n682 ) , .A1( us21_n789 ) , .A2( us21_n811 ) );
  AOI21_X1 us21_U305 (.ZN( us21_n648 ) , .A( us21_n777 ) , .B1( us21_n790 ) , .B2( us21_n803 ) );
  NOR2_X1 us21_U306 (.A2( us21_n811 ) , .A1( us21_n813 ) , .ZN( us21_n819 ) );
  AOI21_X1 us21_U307 (.A( us21_n788 ) , .B2( us21_n789 ) , .B1( us21_n790 ) , .ZN( us21_n791 ) );
  AOI21_X1 us21_U308 (.A( us21_n731 ) , .ZN( us21_n732 ) , .B2( us21_n778 ) , .B1( us21_n790 ) );
  NOR2_X1 us21_U309 (.ZN( us21_n581 ) , .A1( us21_n790 ) , .A2( us21_n815 ) );
  NOR4_X1 us21_U31 (.A4( us21_n774 ) , .A3( us21_n775 ) , .A1( us21_n776 ) , .ZN( us21_n797 ) , .A2( us21_n799 ) );
  NOR2_X1 us21_U310 (.ZN( us21_n532 ) , .A1( us21_n722 ) , .A2( us21_n786 ) );
  AOI21_X1 us21_U311 (.ZN( us21_n639 ) , .B1( us21_n678 ) , .A( us21_n789 ) , .B2( us21_n815 ) );
  NOR2_X1 us21_U312 (.ZN( us21_n709 ) , .A1( us21_n760 ) , .A2( us21_n761 ) );
  NOR2_X1 us21_U313 (.ZN( us21_n565 ) , .A1( us21_n745 ) , .A2( us21_n803 ) );
  NOR2_X1 us21_U314 (.ZN( us21_n680 ) , .A2( us21_n706 ) , .A1( us21_n815 ) );
  INV_X1 us21_U315 (.A( us21_n813 ) , .ZN( us21_n853 ) );
  AOI21_X1 us21_U316 (.ZN( us21_n440 ) , .A( us21_n697 ) , .B1( us21_n731 ) , .B2( us21_n748 ) );
  INV_X1 us21_U317 (.A( us21_n778 ) , .ZN( us21_n848 ) );
  AOI22_X1 us21_U318 (.A2( us21_n780 ) , .ZN( us21_n781 ) , .B2( us21_n829 ) , .A1( us21_n832 ) , .B1( us21_n861 ) );
  NAND2_X1 us21_U319 (.ZN( us21_n712 ) , .A1( us21_n726 ) , .A2( us21_n778 ) );
  NOR4_X1 us21_U32 (.A3( us21_n753 ) , .A2( us21_n754 ) , .A1( us21_n755 ) , .ZN( us21_n756 ) , .A4( us21_n867 ) );
  NAND2_X1 us21_U320 (.ZN( us21_n751 ) , .A1( us21_n761 ) , .A2( us21_n803 ) );
  AOI21_X1 us21_U321 (.ZN( us21_n441 ) , .B1( us21_n787 ) , .B2( us21_n789 ) , .A( us21_n812 ) );
  INV_X1 us21_U322 (.A( us21_n783 ) , .ZN( us21_n844 ) );
  AOI21_X1 us21_U323 (.ZN( us21_n495 ) , .A( us21_n777 ) , .B2( us21_n789 ) , .B1( us21_n802 ) );
  NAND2_X1 us21_U324 (.A2( us21_n760 ) , .A1( us21_n804 ) , .ZN( us21_n808 ) );
  NOR2_X1 us21_U325 (.ZN( us21_n468 ) , .A2( us21_n777 ) , .A1( us21_n813 ) );
  NOR2_X1 us21_U326 (.ZN( us21_n710 ) , .A2( us21_n722 ) , .A1( us21_n788 ) );
  NOR2_X1 us21_U327 (.ZN( us21_n482 ) , .A1( us21_n786 ) , .A2( us21_n803 ) );
  NOR2_X1 us21_U328 (.ZN( us21_n524 ) , .A1( us21_n722 ) , .A2( us21_n748 ) );
  OAI21_X1 us21_U329 (.A( us21_n729 ) , .B1( us21_n730 ) , .ZN( us21_n734 ) , .B2( us21_n803 ) );
  AOI211_X1 us21_U33 (.B( us21_n743 ) , .A( us21_n744 ) , .ZN( us21_n757 ) , .C1( us21_n830 ) , .C2( us21_n851 ) );
  OAI21_X1 us21_U330 (.ZN( us21_n729 ) , .A( us21_n831 ) , .B2( us21_n850 ) , .B1( us21_n871 ) );
  OAI21_X1 us21_U331 (.A( us21_n785 ) , .B2( us21_n786 ) , .B1( us21_n787 ) , .ZN( us21_n793 ) );
  OAI21_X1 us21_U332 (.ZN( us21_n785 ) , .A( us21_n837 ) , .B1( us21_n861 ) , .B2( us21_n871 ) );
  NAND2_X1 us21_U333 (.A1( us21_n697 ) , .A2( us21_n727 ) , .ZN( us21_n780 ) );
  NOR2_X1 us21_U334 (.ZN( us21_n516 ) , .A1( us21_n706 ) , .A2( us21_n786 ) );
  NAND2_X1 us21_U335 (.ZN( us21_n669 ) , .A1( us21_n804 ) , .A2( us21_n814 ) );
  OAI21_X1 us21_U336 (.A( us21_n696 ) , .ZN( us21_n700 ) , .B2( us21_n748 ) , .B1( us21_n802 ) );
  OAI21_X1 us21_U337 (.ZN( us21_n696 ) , .B2( us21_n831 ) , .B1( us21_n836 ) , .A( us21_n858 ) );
  NAND2_X1 us21_U338 (.A2( us21_n747 ) , .A1( us21_n784 ) , .ZN( us21_n807 ) );
  INV_X1 us21_U339 (.A( us21_n722 ) , .ZN( us21_n854 ) );
  NOR3_X1 us21_U34 (.A3( us21_n739 ) , .A2( us21_n740 ) , .A1( us21_n741 ) , .ZN( us21_n758 ) );
  INV_X1 us21_U340 (.A( us21_n815 ) , .ZN( us21_n842 ) );
  AND2_X1 us21_U341 (.ZN( us21_n730 ) , .A1( us21_n777 ) , .A2( us21_n783 ) );
  OAI222_X1 us21_U342 (.ZN( us21_n615 ) , .B1( us21_n695 ) , .C1( us21_n722 ) , .C2( us21_n745 ) , .B2( us21_n784 ) , .A2( us21_n790 ) , .A1( us21_n814 ) );
  AOI221_X1 us21_U343 (.A( us21_n762 ) , .ZN( us21_n772 ) , .C2( us21_n808 ) , .B2( us21_n833 ) , .C1( us21_n853 ) , .B1( us21_n864 ) );
  AOI21_X1 us21_U344 (.B2( us21_n761 ) , .ZN( us21_n762 ) , .A( us21_n786 ) , .B1( us21_n790 ) );
  INV_X1 us21_U345 (.A( us21_n759 ) , .ZN( us21_n833 ) );
  NAND2_X2 us21_U346 (.A2( us21_n439 ) , .A1( us21_n445 ) , .ZN( us21_n782 ) );
  NAND2_X1 us21_U347 (.A1( us21_n453 ) , .A2( us21_n469 ) , .ZN( us21_n801 ) );
  NAND2_X1 us21_U348 (.A1( us21_n452 ) , .A2( us21_n459 ) , .ZN( us21_n811 ) );
  NAND2_X1 us21_U349 (.A1( us21_n451 ) , .A2( us21_n459 ) , .ZN( us21_n742 ) );
  NOR4_X1 us21_U35 (.A4( us21_n732 ) , .A3( us21_n733 ) , .A2( us21_n734 ) , .A1( us21_n735 ) , .ZN( us21_n736 ) );
  NAND2_X1 us21_U350 (.A1( us21_n449 ) , .A2( us21_n452 ) , .ZN( us21_n812 ) );
  NAND2_X1 us21_U351 (.A1( us21_n453 ) , .A2( us21_n460 ) , .ZN( us21_n748 ) );
  NAND2_X1 us21_U352 (.A1( us21_n449 ) , .A2( us21_n469 ) , .ZN( us21_n814 ) );
  NAND2_X1 us21_U353 (.A1( us21_n450 ) , .A2( us21_n463 ) , .ZN( us21_n667 ) );
  NAND2_X1 us21_U354 (.A2( us21_n446 ) , .A1( us21_n458 ) , .ZN( us21_n726 ) );
  NAND2_X1 us21_U355 (.A1( us21_n451 ) , .A2( us21_n470 ) , .ZN( us21_n783 ) );
  NAND2_X1 us21_U356 (.A2( us21_n452 ) , .A1( us21_n470 ) , .ZN( us21_n777 ) );
  NAND2_X1 us21_U357 (.A2( us21_n451 ) , .A1( us21_n453 ) , .ZN( us21_n804 ) );
  NAND2_X1 us21_U358 (.A2( us21_n462 ) , .A1( us21_n463 ) , .ZN( us21_n810 ) );
  NAND2_X1 us21_U359 (.A1( us21_n439 ) , .A2( us21_n458 ) , .ZN( us21_n697 ) );
  AOI211_X1 us21_U36 (.B( us21_n723 ) , .A( us21_n724 ) , .ZN( us21_n737 ) , .C1( us21_n841 ) , .C2( us21_n853 ) );
  NAND2_X1 us21_U360 (.A2( us21_n447 ) , .A1( us21_n450 ) , .ZN( us21_n761 ) );
  NAND2_X1 us21_U361 (.A2( us21_n446 ) , .A1( us21_n450 ) , .ZN( us21_n727 ) );
  NOR2_X1 us21_U362 (.ZN( us21_n445 ) , .A2( us21_n847 ) , .A1( us21_n856 ) );
  NAND2_X1 us21_U363 (.A1( us21_n460 ) , .A2( us21_n470 ) , .ZN( us21_n786 ) );
  NOR2_X1 us21_U364 (.ZN( us21_n463 ) , .A2( us21_n845 ) , .A1( us21_n846 ) );
  NOR2_X1 us21_U365 (.ZN( us21_n451 ) , .A1( us21_n824 ) , .A2( us21_n825 ) );
  NAND2_X1 us21_U366 (.A2( us21_n459 ) , .A1( us21_n460 ) , .ZN( us21_n745 ) );
  NOR2_X1 us21_U367 (.ZN( us21_n449 ) , .A1( us21_n826 ) , .A2( us21_n827 ) );
  NAND2_X1 us21_U368 (.A2( us21_n459 ) , .A1( us21_n469 ) , .ZN( us21_n695 ) );
  NAND2_X1 us21_U369 (.A2( us21_n452 ) , .A1( us21_n453 ) , .ZN( us21_n728 ) );
  NOR3_X1 us21_U37 (.A3( us21_n720 ) , .A1( us21_n721 ) , .ZN( us21_n738 ) , .A2( us21_n739 ) );
  NAND2_X1 us21_U370 (.A1( us21_n449 ) , .A2( us21_n460 ) , .ZN( us21_n788 ) );
  NAND2_X2 us21_U371 (.A2( us21_n446 ) , .A1( us21_n462 ) , .ZN( us21_n813 ) );
  NAND2_X2 us21_U372 (.A2( us21_n439 ) , .A1( us21_n450 ) , .ZN( us21_n789 ) );
  NAND2_X2 us21_U373 (.A1( us21_n447 ) , .A2( us21_n458 ) , .ZN( us21_n790 ) );
  NAND2_X2 us21_U374 (.A1( us21_n439 ) , .A2( us21_n462 ) , .ZN( us21_n706 ) );
  NAND2_X2 us21_U375 (.A2( us21_n469 ) , .A1( us21_n470 ) , .ZN( us21_n815 ) );
  NAND2_X2 us21_U376 (.A1( us21_n445 ) , .A2( us21_n446 ) , .ZN( us21_n784 ) );
  NOR2_X1 us21_U377 (.A2( sa21_6 ) , .A1( sa21_7 ) , .ZN( us21_n462 ) );
  NOR2_X1 us21_U378 (.A2( sa21_4 ) , .ZN( us21_n447 ) , .A1( us21_n846 ) );
  NOR2_X1 us21_U379 (.A2( sa21_5 ) , .ZN( us21_n446 ) , .A1( us21_n845 ) );
  NAND4_X1 us21_U38 (.ZN( sa23_sr_3 ) , .A4( us21_n702 ) , .A3( us21_n703 ) , .A2( us21_n704 ) , .A1( us21_n705 ) );
  NOR2_X1 us21_U380 (.A2( sa21_7 ) , .ZN( us21_n458 ) , .A1( us21_n847 ) );
  NOR2_X1 us21_U381 (.A2( sa21_4 ) , .A1( sa21_5 ) , .ZN( us21_n439 ) );
  NOR2_X1 us21_U382 (.A2( sa21_1 ) , .ZN( us21_n469 ) , .A1( us21_n824 ) );
  NOR2_X1 us21_U383 (.A2( sa21_2 ) , .A1( sa21_3 ) , .ZN( us21_n470 ) );
  NOR2_X1 us21_U384 (.A2( sa21_6 ) , .ZN( us21_n450 ) , .A1( us21_n856 ) );
  NOR2_X1 us21_U385 (.A2( sa21_2 ) , .ZN( us21_n459 ) , .A1( us21_n827 ) );
  NOR2_X1 us21_U386 (.A2( sa21_0 ) , .ZN( us21_n452 ) , .A1( us21_n825 ) );
  NOR2_X1 us21_U387 (.A2( sa21_0 ) , .A1( sa21_1 ) , .ZN( us21_n460 ) );
  NOR2_X1 us21_U388 (.A2( sa21_3 ) , .ZN( us21_n453 ) , .A1( us21_n826 ) );
  INV_X1 us21_U389 (.A( sa21_6 ) , .ZN( us21_n847 ) );
  NOR4_X1 us21_U39 (.A4( us21_n698 ) , .A3( us21_n699 ) , .A2( us21_n700 ) , .A1( us21_n701 ) , .ZN( us21_n702 ) );
  INV_X1 us21_U390 (.A( sa21_3 ) , .ZN( us21_n827 ) );
  INV_X1 us21_U391 (.A( sa21_1 ) , .ZN( us21_n825 ) );
  INV_X1 us21_U392 (.A( sa21_0 ) , .ZN( us21_n824 ) );
  INV_X1 us21_U393 (.A( sa21_2 ) , .ZN( us21_n826 ) );
  INV_X1 us21_U394 (.A( sa21_5 ) , .ZN( us21_n846 ) );
  INV_X1 us21_U395 (.A( sa21_7 ) , .ZN( us21_n856 ) );
  INV_X1 us21_U396 (.A( us21_n784 ) , .ZN( us21_n860 ) );
  AOI21_X1 us21_U397 (.ZN( us21_n498 ) , .A( us21_n695 ) , .B1( us21_n706 ) , .B2( us21_n784 ) );
  INV_X1 us21_U398 (.A( us21_n695 ) , .ZN( us21_n836 ) );
  NOR2_X1 us21_U399 (.A1( us21_n695 ) , .ZN( us21_n768 ) , .A2( us21_n813 ) );
  NAND2_X1 us21_U4 (.A1( us21_n447 ) , .A2( us21_n462 ) , .ZN( us21_n722 ) );
  AOI211_X1 us21_U40 (.B( us21_n692 ) , .A( us21_n693 ) , .ZN( us21_n703 ) , .C2( us21_n829 ) , .C1( us21_n849 ) );
  AOI21_X1 us21_U400 (.ZN( us21_n569 ) , .B2( us21_n695 ) , .B1( us21_n804 ) , .A( us21_n810 ) );
  NOR2_X1 us21_U401 (.ZN( us21_n630 ) , .A2( us21_n695 ) , .A1( us21_n722 ) );
  AOI21_X1 us21_U402 (.ZN( us21_n476 ) , .B2( us21_n695 ) , .A( us21_n747 ) , .B1( us21_n777 ) );
  NOR2_X1 us21_U403 (.ZN( us21_n660 ) , .A2( us21_n695 ) , .A1( us21_n727 ) );
  NOR2_X1 us21_U404 (.A2( us21_n695 ) , .A1( us21_n778 ) , .ZN( us21_n818 ) );
  NOR2_X1 us21_U405 (.A2( us21_n695 ) , .ZN( us21_n714 ) , .A1( us21_n790 ) );
  NOR2_X1 us21_U406 (.ZN( us21_n564 ) , .A2( us21_n695 ) , .A1( us21_n761 ) );
  NOR2_X1 us21_U407 (.ZN( us21_n592 ) , .A2( us21_n695 ) , .A1( us21_n726 ) );
  AOI21_X1 us21_U408 (.ZN( us21_n550 ) , .B1( us21_n667 ) , .A( us21_n695 ) , .B2( us21_n803 ) );
  NOR2_X1 us21_U409 (.ZN( us21_n539 ) , .A2( us21_n695 ) , .A1( us21_n697 ) );
  NOR2_X1 us21_U41 (.ZN( us21_n705 ) , .A2( us21_n774 ) , .A1( us21_n798 ) );
  NOR2_X1 us21_U410 (.ZN( us21_n578 ) , .A2( us21_n695 ) , .A1( us21_n789 ) );
  OAI222_X1 us21_U411 (.B2( us21_n745 ) , .B1( us21_n746 ) , .A2( us21_n747 ) , .ZN( us21_n755 ) , .C2( us21_n803 ) , .C1( us21_n812 ) , .A1( us21_n815 ) );
  OAI222_X1 us21_U412 (.ZN( us21_n503 ) , .C2( us21_n623 ) , .B2( us21_n645 ) , .B1( us21_n745 ) , .A2( us21_n746 ) , .C1( us21_n803 ) , .A1( us21_n804 ) );
  AOI222_X1 us21_U413 (.ZN( us21_n511 ) , .C1( us21_n830 ) , .B2( us21_n835 ) , .A2( us21_n841 ) , .C2( us21_n860 ) , .B1( us21_n861 ) , .A1( us21_n864 ) );
  AOI222_X1 us21_U414 (.ZN( us21_n603 ) , .B2( us21_n669 ) , .B1( us21_n751 ) , .C2( us21_n829 ) , .A1( us21_n831 ) , .A2( us21_n860 ) , .C1( us21_n861 ) );
  AOI221_X1 us21_U415 (.A( us21_n481 ) , .ZN( us21_n486 ) , .B1( us21_n829 ) , .C2( us21_n842 ) , .C1( us21_n850 ) , .B2( us21_n860 ) );
  NOR2_X1 us21_U416 (.ZN( us21_n787 ) , .A2( us21_n860 ) , .A1( us21_n866 ) );
  OAI221_X1 us21_U417 (.A( us21_n781 ) , .C2( us21_n782 ) , .B2( us21_n783 ) , .B1( us21_n784 ) , .ZN( us21_n794 ) , .C1( us21_n811 ) );
  NAND2_X1 us21_U418 (.A1( us21_n727 ) , .A2( us21_n782 ) , .ZN( us21_n809 ) );
  OAI22_X1 us21_U419 (.ZN( us21_n586 ) , .A2( us21_n745 ) , .B2( us21_n760 ) , .A1( us21_n761 ) , .B1( us21_n782 ) );
  NOR2_X1 us21_U42 (.ZN( us21_n802 ) , .A1( us21_n852 ) , .A2( us21_n859 ) );
  OAI221_X1 us21_U420 (.A( us21_n694 ) , .ZN( us21_n701 ) , .C2( us21_n782 ) , .C1( us21_n783 ) , .B1( us21_n784 ) , .B2( us21_n804 ) );
  AOI21_X1 us21_U421 (.ZN( us21_n590 ) , .B1( us21_n726 ) , .B2( us21_n782 ) , .A( us21_n788 ) );
  AOI21_X1 us21_U422 (.ZN( us21_n646 ) , .A( us21_n760 ) , .B2( us21_n782 ) , .B1( us21_n790 ) );
  AOI21_X1 us21_U423 (.ZN( us21_n621 ) , .B1( us21_n697 ) , .A( us21_n777 ) , .B2( us21_n782 ) );
  OAI22_X1 us21_U424 (.ZN( us21_n679 ) , .A1( us21_n697 ) , .A2( us21_n728 ) , .B2( us21_n782 ) , .B1( us21_n815 ) );
  OAI21_X1 us21_U425 (.A( us21_n611 ) , .ZN( us21_n614 ) , .B1( us21_n623 ) , .B2( us21_n782 ) );
  NOR2_X1 us21_U426 (.ZN( us21_n608 ) , .A1( us21_n782 ) , .A2( us21_n814 ) );
  OAI222_X1 us21_U427 (.A2( us21_n667 ) , .ZN( us21_n672 ) , .B1( us21_n745 ) , .B2( us21_n782 ) , .C2( us21_n786 ) , .C1( us21_n813 ) , .A1( us21_n815 ) );
  NOR2_X1 us21_U428 (.ZN( us21_n649 ) , .A1( us21_n782 ) , .A2( us21_n786 ) );
  NOR2_X1 us21_U429 (.ZN( us21_n598 ) , .A2( us21_n695 ) , .A1( us21_n782 ) );
  NAND4_X1 us21_U43 (.ZN( sa23_sr_2 ) , .A4( us21_n641 ) , .A3( us21_n642 ) , .A2( us21_n643 ) , .A1( us21_n644 ) );
  NOR2_X1 us21_U430 (.ZN( us21_n551 ) , .A2( us21_n742 ) , .A1( us21_n782 ) );
  INV_X1 us21_U431 (.A( us21_n782 ) , .ZN( us21_n859 ) );
  AOI221_X1 us21_U432 (.A( us21_n574 ) , .ZN( us21_n585 ) , .B2( us21_n829 ) , .C2( us21_n841 ) , .B1( us21_n852 ) , .C1( us21_n859 ) );
  AOI21_X1 us21_U433 (.ZN( us21_n574 ) , .B2( us21_n722 ) , .B1( us21_n746 ) , .A( us21_n783 ) );
  INV_X1 us21_U434 (.A( sa21_4 ) , .ZN( us21_n845 ) );
  AOI211_X1 us21_U435 (.A( us21_n635 ) , .ZN( us21_n643 ) , .B( us21_n741 ) , .C2( us21_n837 ) , .C1( us21_n852 ) );
  NAND4_X1 us21_U436 (.A4( us21_n631 ) , .A3( us21_n632 ) , .A2( us21_n633 ) , .A1( us21_n634 ) , .ZN( us21_n741 ) );
  NAND3_X1 us21_U437 (.ZN( sa23_sr_6 ) , .A3( us21_n795 ) , .A2( us21_n796 ) , .A1( us21_n797 ) );
  NAND3_X1 us21_U438 (.ZN( sa23_sr_5 ) , .A3( us21_n756 ) , .A2( us21_n757 ) , .A1( us21_n758 ) );
  NAND3_X1 us21_U439 (.ZN( sa23_sr_4 ) , .A3( us21_n736 ) , .A2( us21_n737 ) , .A1( us21_n738 ) );
  AOI222_X1 us21_U44 (.B2( us21_n636 ) , .ZN( us21_n642 ) , .B1( us21_n839 ) , .A1( us21_n840 ) , .C2( us21_n844 ) , .C1( us21_n861 ) , .A2( us21_n863 ) );
  NAND3_X1 us21_U440 (.A3( us21_n673 ) , .A2( us21_n674 ) , .A1( us21_n675 ) , .ZN( us21_n805 ) );
  NAND3_X1 us21_U441 (.ZN( us21_n636 ) , .A3( us21_n706 ) , .A2( us21_n722 ) , .A1( us21_n790 ) );
  NAND3_X1 us21_U442 (.A3( us21_n616 ) , .A2( us21_n617 ) , .A1( us21_n618 ) , .ZN( us21_n723 ) );
  NAND3_X1 us21_U443 (.A3( us21_n583 ) , .A2( us21_n584 ) , .A1( us21_n585 ) , .ZN( us21_n619 ) );
  NAND3_X1 us21_U444 (.ZN( us21_n563 ) , .A3( us21_n678 ) , .A2( us21_n748 ) , .A1( us21_n783 ) );
  NAND3_X1 us21_U445 (.A3( us21_n521 ) , .A2( us21_n522 ) , .A1( us21_n523 ) , .ZN( us21_n740 ) );
  NAND3_X1 us21_U446 (.A3( us21_n510 ) , .A1( us21_n511 ) , .ZN( us21_n606 ) , .A2( us21_n869 ) );
  NAND3_X1 us21_U447 (.A3( us21_n465 ) , .A2( us21_n466 ) , .A1( us21_n467 ) , .ZN( us21_n775 ) );
  NOR4_X1 us21_U45 (.A4( us21_n637 ) , .A3( us21_n638 ) , .A2( us21_n639 ) , .A1( us21_n640 ) , .ZN( us21_n641 ) );
  NOR3_X1 us21_U46 (.A2( us21_n605 ) , .A1( us21_n606 ) , .ZN( us21_n644 ) , .A3( us21_n720 ) );
  NAND4_X1 us21_U47 (.ZN( sa23_sr_0 ) , .A4( us21_n499 ) , .A3( us21_n500 ) , .A2( us21_n501 ) , .A1( us21_n502 ) );
  NOR4_X1 us21_U48 (.A4( us21_n496 ) , .A3( us21_n497 ) , .A2( us21_n498 ) , .ZN( us21_n499 ) , .A1( us21_n525 ) );
  AOI221_X1 us21_U49 (.A( us21_n495 ) , .ZN( us21_n500 ) , .B2( us21_n841 ) , .C1( us21_n844 ) , .C2( us21_n858 ) , .B1( us21_n860 ) );
  NAND2_X1 us21_U5 (.A1( us21_n445 ) , .A2( us21_n447 ) , .ZN( us21_n803 ) );
  AOI211_X1 us21_U50 (.A( us21_n494 ) , .ZN( us21_n501 ) , .B( us21_n800 ) , .C2( us21_n837 ) , .C1( us21_n849 ) );
  NAND4_X1 us21_U51 (.ZN( sa23_sr_1 ) , .A4( us21_n593 ) , .A3( us21_n594 ) , .A2( us21_n595 ) , .A1( us21_n596 ) );
  AOI211_X1 us21_U52 (.B( us21_n587 ) , .A( us21_n588 ) , .ZN( us21_n594 ) , .C2( us21_n809 ) , .C1( us21_n831 ) );
  NOR4_X1 us21_U53 (.A4( us21_n589 ) , .A3( us21_n590 ) , .A2( us21_n591 ) , .A1( us21_n592 ) , .ZN( us21_n593 ) );
  AOI211_X1 us21_U54 (.A( us21_n586 ) , .ZN( us21_n595 ) , .B( us21_n619 ) , .C1( us21_n843 ) , .C2( us21_n853 ) );
  NAND4_X1 us21_U55 (.A4( us21_n601 ) , .A3( us21_n602 ) , .A2( us21_n603 ) , .A1( us21_n604 ) , .ZN( us21_n720 ) );
  NOR3_X1 us21_U56 (.A1( us21_n597 ) , .ZN( us21_n602 ) , .A3( us21_n661 ) , .A2( us21_n768 ) );
  NOR4_X1 us21_U57 (.A3( us21_n598 ) , .A2( us21_n599 ) , .A1( us21_n600 ) , .ZN( us21_n601 ) , .A4( us21_n653 ) );
  AOI222_X1 us21_U58 (.ZN( us21_n604 ) , .A1( us21_n828 ) , .C2( us21_n835 ) , .B1( us21_n840 ) , .A2( us21_n854 ) , .B2( us21_n859 ) , .C1( us21_n866 ) );
  AOI222_X1 us21_U59 (.ZN( us21_n467 ) , .B1( us21_n830 ) , .A1( us21_n837 ) , .C1( us21_n840 ) , .C2( us21_n849 ) , .A2( us21_n853 ) , .B2( us21_n863 ) );
  NOR3_X1 us21_U6 (.ZN( us21_n596 ) , .A1( us21_n606 ) , .A3( us21_n721 ) , .A2( us21_n740 ) );
  NOR4_X1 us21_U60 (.A1( us21_n464 ) , .ZN( us21_n465 ) , .A4( us21_n540 ) , .A2( us21_n552 ) , .A3( us21_n612 ) );
  AOI221_X1 us21_U61 (.ZN( us21_n466 ) , .C2( us21_n712 ) , .B2( us21_n829 ) , .C1( us21_n843 ) , .B1( us21_n858 ) , .A( us21_n862 ) );
  NAND4_X1 us21_U62 (.A4( us21_n483 ) , .A3( us21_n484 ) , .A2( us21_n485 ) , .A1( us21_n486 ) , .ZN( us21_n776 ) );
  NOR4_X1 us21_U63 (.ZN( us21_n484 ) , .A1( us21_n505 ) , .A2( us21_n517 ) , .A4( us21_n544 ) , .A3( us21_n609 ) );
  NOR4_X1 us21_U64 (.A4( us21_n482 ) , .ZN( us21_n485 ) , .A1( us21_n564 ) , .A2( us21_n579 ) , .A3( us21_n600 ) );
  NOR4_X1 us21_U65 (.ZN( us21_n483 ) , .A2( us21_n531 ) , .A1( us21_n556 ) , .A3( us21_n629 ) , .A4( us21_n716 ) );
  AOI211_X1 us21_U66 (.B( us21_n621 ) , .A( us21_n622 ) , .ZN( us21_n633 ) , .C2( us21_n834 ) , .C1( us21_n861 ) );
  NOR4_X1 us21_U67 (.A4( us21_n627 ) , .A3( us21_n628 ) , .A2( us21_n629 ) , .A1( us21_n630 ) , .ZN( us21_n631 ) );
  NOR4_X1 us21_U68 (.A4( us21_n624 ) , .A3( us21_n625 ) , .A2( us21_n626 ) , .ZN( us21_n632 ) , .A1( us21_n662 ) );
  NOR4_X1 us21_U69 (.A4( us21_n512 ) , .A3( us21_n513 ) , .A2( us21_n514 ) , .A1( us21_n515 ) , .ZN( us21_n522 ) );
  NOR3_X1 us21_U7 (.A3( us21_n798 ) , .A2( us21_n799 ) , .A1( us21_n800 ) , .ZN( us21_n823 ) );
  AOI222_X1 us21_U70 (.ZN( us21_n523 ) , .A1( us21_n832 ) , .B2( us21_n835 ) , .C1( us21_n842 ) , .C2( us21_n848 ) , .A2( us21_n850 ) , .B1( us21_n864 ) );
  NOR4_X1 us21_U71 (.A3( us21_n519 ) , .A1( us21_n520 ) , .ZN( us21_n521 ) , .A2( us21_n671 ) , .A4( us21_n767 ) );
  NAND4_X1 us21_U72 (.A4( us21_n655 ) , .A3( us21_n656 ) , .A2( us21_n657 ) , .A1( us21_n658 ) , .ZN( us21_n798 ) );
  NOR3_X1 us21_U73 (.A3( us21_n646 ) , .A2( us21_n647 ) , .A1( us21_n648 ) , .ZN( us21_n657 ) );
  NOR3_X1 us21_U74 (.A3( us21_n649 ) , .A2( us21_n650 ) , .A1( us21_n651 ) , .ZN( us21_n656 ) );
  NOR3_X1 us21_U75 (.A3( us21_n652 ) , .A2( us21_n653 ) , .A1( us21_n654 ) , .ZN( us21_n655 ) );
  NAND4_X1 us21_U76 (.A4( us21_n558 ) , .A3( us21_n559 ) , .A2( us21_n560 ) , .A1( us21_n561 ) , .ZN( us21_n605 ) );
  NOR4_X1 us21_U77 (.A4( us21_n550 ) , .A3( us21_n551 ) , .A2( us21_n552 ) , .A1( us21_n553 ) , .ZN( us21_n560 ) );
  NOR4_X1 us21_U78 (.A4( us21_n554 ) , .A3( us21_n555 ) , .A2( us21_n556 ) , .A1( us21_n557 ) , .ZN( us21_n558 ) );
  NOR4_X1 us21_U79 (.ZN( us21_n559 ) , .A1( us21_n651 ) , .A3( us21_n659 ) , .A4( us21_n683 ) , .A2( us21_n766 ) );
  NOR3_X1 us21_U8 (.ZN( us21_n502 ) , .A2( us21_n677 ) , .A3( us21_n775 ) , .A1( us21_n874 ) );
  NAND4_X1 us21_U80 (.A4( us21_n770 ) , .A3( us21_n771 ) , .A2( us21_n772 ) , .A1( us21_n773 ) , .ZN( us21_n799 ) );
  NOR3_X1 us21_U81 (.A3( us21_n763 ) , .A2( us21_n764 ) , .A1( us21_n765 ) , .ZN( us21_n771 ) );
  NOR4_X1 us21_U82 (.A4( us21_n766 ) , .A3( us21_n767 ) , .A2( us21_n768 ) , .A1( us21_n769 ) , .ZN( us21_n770 ) );
  AOI222_X1 us21_U83 (.ZN( us21_n773 ) , .A1( us21_n828 ) , .C1( us21_n832 ) , .B2( us21_n839 ) , .A2( us21_n848 ) , .B1( us21_n859 ) , .C2( us21_n871 ) );
  NOR4_X1 us21_U84 (.A4( us21_n507 ) , .A2( us21_n508 ) , .A1( us21_n509 ) , .ZN( us21_n510 ) , .A3( us21_n668 ) );
  INV_X1 us21_U85 (.A( us21_n503 ) , .ZN( us21_n869 ) );
  NOR4_X1 us21_U86 (.A4( us21_n659 ) , .A3( us21_n660 ) , .A2( us21_n661 ) , .A1( us21_n662 ) , .ZN( us21_n675 ) );
  NOR4_X1 us21_U87 (.A4( us21_n663 ) , .A3( us21_n664 ) , .A2( us21_n665 ) , .A1( us21_n666 ) , .ZN( us21_n674 ) );
  NOR4_X1 us21_U88 (.A3( us21_n671 ) , .A1( us21_n672 ) , .ZN( us21_n673 ) , .A4( us21_n713 ) , .A2( us21_n857 ) );
  NOR2_X1 us21_U89 (.ZN( us21_n623 ) , .A2( us21_n834 ) , .A1( us21_n837 ) );
  INV_X1 us21_U9 (.A( us21_n704 ) , .ZN( us21_n874 ) );
  NOR2_X1 us21_U90 (.ZN( us21_n759 ) , .A1( us21_n831 ) , .A2( us21_n832 ) );
  NAND4_X1 us21_U91 (.A4( us21_n454 ) , .A3( us21_n455 ) , .A2( us21_n456 ) , .A1( us21_n457 ) , .ZN( us21_n677 ) );
  NOR3_X1 us21_U92 (.ZN( us21_n455 ) , .A3( us21_n528 ) , .A1( us21_n553 ) , .A2( us21_n568 ) );
  AOI221_X1 us21_U93 (.A( us21_n448 ) , .ZN( us21_n457 ) , .C2( us21_n751 ) , .B1( us21_n830 ) , .C1( us21_n840 ) , .B2( us21_n859 ) );
  NOR4_X1 us21_U94 (.ZN( us21_n456 ) , .A2( us21_n507 ) , .A1( us21_n597 ) , .A4( us21_n626 ) , .A3( us21_n709 ) );
  NAND4_X1 us21_U95 (.ZN( sa23_sr_7 ) , .A4( us21_n820 ) , .A3( us21_n821 ) , .A2( us21_n822 ) , .A1( us21_n823 ) );
  NOR4_X1 us21_U96 (.A4( us21_n816 ) , .A3( us21_n817 ) , .A2( us21_n818 ) , .A1( us21_n819 ) , .ZN( us21_n820 ) );
  AOI222_X1 us21_U97 (.C2( us21_n807 ) , .B2( us21_n808 ) , .A2( us21_n809 ) , .ZN( us21_n821 ) , .C1( us21_n830 ) , .A1( us21_n837 ) , .B1( us21_n851 ) );
  AOI211_X1 us21_U98 (.B( us21_n805 ) , .A( us21_n806 ) , .ZN( us21_n822 ) , .C1( us21_n840 ) , .C2( us21_n848 ) );
  NAND4_X1 us21_U99 (.A4( us21_n533 ) , .A3( us21_n534 ) , .A2( us21_n535 ) , .A1( us21_n536 ) , .ZN( us21_n620 ) );
  INV_X1 us23_U10 (.A( us23_n679 ) , .ZN( us23_n839 ) );
  NOR4_X1 us23_U100 (.A4( us23_n483 ) , .ZN( us23_n486 ) , .A1( us23_n565 ) , .A2( us23_n580 ) , .A3( us23_n601 ) );
  NOR4_X1 us23_U101 (.ZN( us23_n485 ) , .A1( us23_n506 ) , .A2( us23_n518 ) , .A4( us23_n545 ) , .A3( us23_n610 ) );
  NOR4_X1 us23_U102 (.ZN( us23_n484 ) , .A2( us23_n532 ) , .A1( us23_n557 ) , .A3( us23_n630 ) , .A4( us23_n717 ) );
  NAND4_X1 us23_U103 (.A4( us23_n690 ) , .A3( us23_n691 ) , .A1( us23_n692 ) , .ZN( us23_n775 ) , .A2( us23_n871 ) );
  AOI221_X1 us23_U104 (.A( us23_n680 ) , .ZN( us23_n691 ) , .B2( us23_n839 ) , .C1( us23_n841 ) , .C2( us23_n861 ) , .B1( us23_n864 ) );
  INV_X1 us23_U105 (.A( us23_n678 ) , .ZN( us23_n871 ) );
  NOR4_X1 us23_U106 (.A4( us23_n686 ) , .A3( us23_n687 ) , .A2( us23_n688 ) , .A1( us23_n689 ) , .ZN( us23_n690 ) );
  NAND4_X1 us23_U107 (.A4( us23_n559 ) , .A3( us23_n560 ) , .A2( us23_n561 ) , .A1( us23_n562 ) , .ZN( us23_n606 ) );
  NOR4_X1 us23_U108 (.ZN( us23_n560 ) , .A1( us23_n652 ) , .A3( us23_n660 ) , .A4( us23_n684 ) , .A2( us23_n767 ) );
  NOR4_X1 us23_U109 (.A4( us23_n551 ) , .A3( us23_n552 ) , .A2( us23_n553 ) , .A1( us23_n554 ) , .ZN( us23_n561 ) );
  NOR4_X1 us23_U11 (.A4( us23_n444 ) , .A3( us23_n445 ) , .A2( us23_n515 ) , .A1( us23_n540 ) , .ZN( us23_n705 ) );
  NOR4_X1 us23_U110 (.A4( us23_n555 ) , .A3( us23_n556 ) , .A2( us23_n557 ) , .A1( us23_n558 ) , .ZN( us23_n559 ) );
  NAND4_X1 us23_U111 (.A4( us23_n718 ) , .A3( us23_n719 ) , .A2( us23_n720 ) , .ZN( us23_n740 ) , .A1( us23_n856 ) );
  INV_X1 us23_U112 (.A( us23_n708 ) , .ZN( us23_n856 ) );
  AOI221_X1 us23_U113 (.A( us23_n709 ) , .ZN( us23_n720 ) , .C2( us23_n843 ) , .B2( us23_n844 ) , .C1( us23_n860 ) , .B1( us23_n861 ) );
  NOR4_X1 us23_U114 (.A4( us23_n714 ) , .A3( us23_n715 ) , .A2( us23_n716 ) , .A1( us23_n717 ) , .ZN( us23_n718 ) );
  NAND4_X1 us23_U115 (.A4( us23_n472 ) , .A3( us23_n473 ) , .A2( us23_n474 ) , .A1( us23_n475 ) , .ZN( us23_n677 ) );
  NOR4_X1 us23_U116 (.A4( us23_n469 ) , .ZN( us23_n475 ) , .A3( us23_n555 ) , .A1( us23_n734 ) , .A2( us23_n754 ) );
  NOR4_X1 us23_U117 (.ZN( us23_n474 ) , .A1( us23_n530 ) , .A3( us23_n567 ) , .A4( us23_n599 ) , .A2( us23_n641 ) );
  NOR4_X1 us23_U118 (.ZN( us23_n473 ) , .A1( us23_n505 ) , .A3( us23_n543 ) , .A2( us23_n582 ) , .A4( us23_n715 ) );
  NOR2_X1 us23_U119 (.ZN( us23_n732 ) , .A2( us23_n831 ) , .A1( us23_n844 ) );
  OR3_X1 us23_U12 (.ZN( us23_n445 ) , .A1( us23_n527 ) , .A3( us23_n576 ) , .A2( us23_n874 ) );
  NOR2_X1 us23_U120 (.ZN( us23_n788 ) , .A2( us23_n861 ) , .A1( us23_n867 ) );
  NAND4_X1 us23_U121 (.A4( us23_n572 ) , .A3( us23_n573 ) , .A1( us23_n574 ) , .ZN( us23_n722 ) , .A2( us23_n873 ) );
  NOR4_X1 us23_U122 (.A4( us23_n568 ) , .A3( us23_n569 ) , .A2( us23_n570 ) , .A1( us23_n571 ) , .ZN( us23_n572 ) );
  AOI221_X1 us23_U123 (.A( us23_n563 ) , .C2( us23_n564 ) , .ZN( us23_n573 ) , .B2( us23_n844 ) , .B1( us23_n851 ) , .C1( us23_n852 ) );
  INV_X1 us23_U124 (.A( us23_n606 ) , .ZN( us23_n873 ) );
  NAND4_X1 us23_U125 (.A4( us23_n492 ) , .A3( us23_n493 ) , .A1( us23_n494 ) , .ZN( us23_n801 ) , .A2( us23_n866 ) );
  AOI221_X1 us23_U126 (.A( us23_n488 ) , .ZN( us23_n493 ) , .B2( us23_n835 ) , .C2( us23_n840 ) , .C1( us23_n850 ) , .B1( us23_n859 ) );
  INV_X1 us23_U127 (.A( us23_n777 ) , .ZN( us23_n866 ) );
  NOR2_X1 us23_U128 (.ZN( us23_n494 ) , .A1( us23_n677 ) , .A2( us23_n693 ) );
  NOR2_X1 us23_U129 (.ZN( us23_n747 ) , .A1( us23_n860 ) , .A2( us23_n861 ) );
  OR4_X1 us23_U13 (.A4( us23_n441 ) , .A2( us23_n442 ) , .A1( us23_n443 ) , .ZN( us23_n444 ) , .A3( us23_n552 ) );
  AOI222_X1 us23_U130 (.ZN( us23_n512 ) , .C1( us23_n831 ) , .B2( us23_n836 ) , .A2( us23_n842 ) , .C2( us23_n861 ) , .B1( us23_n862 ) , .A1( us23_n865 ) );
  NOR4_X1 us23_U131 (.A4( us23_n508 ) , .A2( us23_n509 ) , .A1( us23_n510 ) , .ZN( us23_n511 ) , .A3( us23_n669 ) );
  INV_X1 us23_U132 (.A( us23_n504 ) , .ZN( us23_n870 ) );
  INV_X1 us23_U133 (.A( us23_n761 ) , .ZN( us23_n829 ) );
  NOR2_X1 us23_U134 (.ZN( us23_n646 ) , .A1( us23_n853 ) , .A2( us23_n867 ) );
  OR4_X1 us23_U135 (.A4( us23_n579 ) , .A3( us23_n580 ) , .A2( us23_n581 ) , .A1( us23_n582 ) , .ZN( us23_n583 ) );
  OR4_X1 us23_U136 (.A4( us23_n681 ) , .A3( us23_n682 ) , .A2( us23_n683 ) , .A1( us23_n684 ) , .ZN( us23_n689 ) );
  OR4_X1 us23_U137 (.A4( us23_n565 ) , .A3( us23_n566 ) , .A2( us23_n567 ) , .ZN( us23_n571 ) , .A1( us23_n664 ) );
  OR4_X1 us23_U138 (.A4( us23_n517 ) , .A2( us23_n518 ) , .A1( us23_n519 ) , .ZN( us23_n521 ) , .A3( us23_n820 ) );
  OR4_X1 us23_U139 (.ZN( us23_n465 ) , .A4( us23_n517 ) , .A3( us23_n528 ) , .A2( us23_n577 ) , .A1( us23_n711 ) );
  INV_X1 us23_U14 (.A( us23_n612 ) , .ZN( us23_n874 ) );
  NAND2_X1 us23_U140 (.ZN( us23_n612 ) , .A2( us23_n836 ) , .A1( us23_n872 ) );
  OR3_X1 us23_U141 (.A3( us23_n505 ) , .A2( us23_n506 ) , .A1( us23_n507 ) , .ZN( us23_n510 ) );
  AOI221_X1 us23_U142 (.A( us23_n712 ) , .B2( us23_n713 ) , .ZN( us23_n719 ) , .C1( us23_n831 ) , .B1( us23_n838 ) , .C2( us23_n862 ) );
  OR2_X1 us23_U143 (.A2( us23_n710 ) , .A1( us23_n711 ) , .ZN( us23_n712 ) );
  INV_X1 us23_U144 (.A( us23_n462 ) , .ZN( us23_n863 ) );
  OAI21_X1 us23_U145 (.ZN( us23_n462 ) , .B1( us23_n808 ) , .A( us23_n833 ) , .B2( us23_n850 ) );
  INV_X1 us23_U146 (.A( us23_n753 ) , .ZN( us23_n868 ) );
  OAI21_X1 us23_U147 (.B1( us23_n752 ) , .ZN( us23_n753 ) , .A( us23_n844 ) , .B2( us23_n867 ) );
  INV_X1 us23_U148 (.A( us23_n671 ) , .ZN( us23_n858 ) );
  AOI21_X1 us23_U149 (.A( us23_n669 ) , .B1( us23_n670 ) , .ZN( us23_n671 ) , .B2( us23_n855 ) );
  INV_X1 us23_U15 (.A( us23_n748 ) , .ZN( us23_n862 ) );
  AOI222_X1 us23_U150 (.ZN( us23_n659 ) , .A2( us23_n838 ) , .B1( us23_n840 ) , .C2( us23_n844 ) , .A1( us23_n859 ) , .C1( us23_n862 ) , .B2( us23_n869 ) );
  INV_X1 us23_U151 (.A( us23_n646 ) , .ZN( us23_n869 ) );
  OAI222_X1 us23_U152 (.B2( us23_n707 ) , .ZN( us23_n708 ) , .C2( us23_n723 ) , .B1( us23_n746 ) , .A1( us23_n805 ) , .C1( us23_n813 ) , .A2( us23_n814 ) );
  OAI222_X1 us23_U153 (.A2( us23_n668 ) , .ZN( us23_n673 ) , .B1( us23_n746 ) , .B2( us23_n783 ) , .C2( us23_n787 ) , .C1( us23_n814 ) , .A1( us23_n816 ) );
  NAND2_X1 us23_U154 (.A1( us23_n446 ) , .A2( us23_n464 ) , .ZN( us23_n748 ) );
  NOR4_X1 us23_U155 (.A2( us23_n490 ) , .A1( us23_n491 ) , .ZN( us23_n492 ) , .A3( us23_n579 ) , .A4( us23_n611 ) );
  OR4_X1 us23_U156 (.ZN( us23_n491 ) , .A4( us23_n533 ) , .A2( us23_n546 ) , .A1( us23_n558 ) , .A3( us23_n631 ) );
  OAI22_X1 us23_U157 (.B1( us23_n489 ) , .ZN( us23_n490 ) , .A1( us23_n685 ) , .A2( us23_n762 ) , .B2( us23_n816 ) );
  NOR3_X1 us23_U158 (.ZN( us23_n489 ) , .A1( us23_n781 ) , .A2( us23_n849 ) , .A3( us23_n862 ) );
  AOI22_X1 us23_U159 (.ZN( us23_n695 ) , .A1( us23_n829 ) , .B2( us23_n842 ) , .A2( us23_n864 ) , .B1( us23_n867 ) );
  AOI222_X1 us23_U16 (.ZN( us23_n604 ) , .B2( us23_n670 ) , .B1( us23_n752 ) , .C2( us23_n830 ) , .A1( us23_n832 ) , .A2( us23_n861 ) , .C1( us23_n862 ) );
  AOI21_X1 us23_U160 (.ZN( us23_n638 ) , .B2( us23_n748 ) , .A( us23_n787 ) , .B1( us23_n811 ) );
  AOI21_X1 us23_U161 (.ZN( us23_n639 ) , .B2( us23_n746 ) , .A( us23_n791 ) , .B1( us23_n802 ) );
  AOI21_X1 us23_U162 (.ZN( us23_n640 ) , .B1( us23_n679 ) , .A( us23_n790 ) , .B2( us23_n816 ) );
  INV_X1 us23_U163 (.A( us23_n729 ) , .ZN( us23_n838 ) );
  AOI221_X1 us23_U164 (.A( us23_n763 ) , .ZN( us23_n773 ) , .C2( us23_n809 ) , .B2( us23_n834 ) , .C1( us23_n854 ) , .B1( us23_n865 ) );
  AOI21_X1 us23_U165 (.B2( us23_n762 ) , .ZN( us23_n763 ) , .A( us23_n787 ) , .B1( us23_n791 ) );
  INV_X1 us23_U166 (.A( us23_n760 ) , .ZN( us23_n834 ) );
  AOI221_X1 us23_U167 (.A( us23_n449 ) , .ZN( us23_n458 ) , .C2( us23_n752 ) , .B1( us23_n831 ) , .C1( us23_n841 ) , .B2( us23_n860 ) );
  AOI21_X1 us23_U168 (.ZN( us23_n449 ) , .B2( us23_n791 ) , .A( us23_n802 ) , .B1( us23_n814 ) );
  AOI221_X1 us23_U169 (.A( us23_n482 ) , .ZN( us23_n487 ) , .B1( us23_n830 ) , .C2( us23_n843 ) , .C1( us23_n851 ) , .B2( us23_n861 ) );
  AOI222_X1 us23_U17 (.ZN( us23_n562 ) , .B1( us23_n829 ) , .C1( us23_n840 ) , .A2( us23_n842 ) , .A1( us23_n853 ) , .B2( us23_n862 ) , .C2( us23_n872 ) );
  OAI22_X1 us23_U170 (.ZN( us23_n482 ) , .A1( us23_n707 ) , .B2( us23_n784 ) , .A2( us23_n805 ) , .B1( us23_n811 ) );
  INV_X1 us23_U171 (.A( us23_n789 ) , .ZN( us23_n831 ) );
  NAND2_X1 us23_U172 (.A1( us23_n450 ) , .A2( us23_n452 ) , .ZN( us23_n761 ) );
  INV_X1 us23_U173 (.A( us23_n783 ) , .ZN( us23_n860 ) );
  INV_X1 us23_U174 (.A( us23_n785 ) , .ZN( us23_n861 ) );
  INV_X1 us23_U175 (.A( us23_n815 ) , .ZN( us23_n830 ) );
  OAI22_X1 us23_U176 (.ZN( us23_n709 ) , .A2( us23_n727 ) , .B2( us23_n728 ) , .A1( us23_n743 ) , .B1( us23_n812 ) );
  OAI22_X1 us23_U177 (.ZN( us23_n623 ) , .B1( us23_n668 ) , .B2( us23_n746 ) , .A1( us23_n814 ) , .A2( us23_n815 ) );
  OAI22_X1 us23_U178 (.ZN( us23_n587 ) , .A2( us23_n746 ) , .B2( us23_n761 ) , .A1( us23_n762 ) , .B1( us23_n783 ) );
  INV_X1 us23_U179 (.A( us23_n743 ) , .ZN( us23_n836 ) );
  NOR4_X1 us23_U18 (.ZN( us23_n472 ) , .A2( us23_n520 ) , .A4( us23_n593 ) , .A1( us23_n608 ) , .A3( us23_n628 ) );
  INV_X1 us23_U180 (.A( us23_n787 ) , .ZN( us23_n844 ) );
  OAI22_X1 us23_U181 (.A1( us23_n723 ) , .ZN( us23_n725 ) , .B2( us23_n749 ) , .B1( us23_n811 ) , .A2( us23_n815 ) );
  OAI22_X1 us23_U182 (.B2( us23_n778 ) , .B1( us23_n779 ) , .ZN( us23_n780 ) , .A2( us23_n813 ) , .A1( us23_n814 ) );
  OAI22_X1 us23_U183 (.ZN( us23_n680 ) , .A1( us23_n698 ) , .A2( us23_n729 ) , .B2( us23_n783 ) , .B1( us23_n816 ) );
  OAI22_X1 us23_U184 (.B2( us23_n749 ) , .B1( us23_n750 ) , .A1( us23_n751 ) , .ZN( us23_n755 ) , .A2( us23_n805 ) );
  NOR2_X1 us23_U185 (.ZN( us23_n750 ) , .A2( us23_n851 ) , .A1( us23_n859 ) );
  NOR3_X1 us23_U186 (.ZN( us23_n751 ) , .A2( us23_n852 ) , .A1( us23_n862 ) , .A3( us23_n864 ) );
  OAI22_X1 us23_U187 (.B2( us23_n743 ) , .ZN( us23_n745 ) , .A2( us23_n761 ) , .B1( us23_n779 ) , .A1( us23_n791 ) );
  INV_X1 us23_U188 (.A( us23_n802 ) , .ZN( us23_n842 ) );
  INV_X1 us23_U189 (.A( us23_n813 ) , .ZN( us23_n832 ) );
  NOR4_X1 us23_U19 (.A4( us23_n531 ) , .A3( us23_n532 ) , .A2( us23_n533 ) , .ZN( us23_n534 ) , .A1( us23_n819 ) );
  INV_X1 us23_U190 (.A( us23_n804 ) , .ZN( us23_n859 ) );
  OAI22_X1 us23_U191 (.B2( us23_n802 ) , .B1( us23_n803 ) , .A2( us23_n804 ) , .A1( us23_n805 ) , .ZN( us23_n807 ) );
  OAI22_X1 us23_U192 (.ZN( us23_n495 ) , .A2( us23_n743 ) , .A1( us23_n779 ) , .B1( us23_n790 ) , .B2( us23_n805 ) );
  OAI22_X1 us23_U193 (.ZN( us23_n488 ) , .A1( us23_n723 ) , .B2( us23_n727 ) , .B1( us23_n729 ) , .A2( us23_n778 ) );
  INV_X1 us23_U194 (.A( us23_n668 ) , .ZN( us23_n864 ) );
  OAI22_X1 us23_U195 (.ZN( us23_n694 ) , .A2( us23_n729 ) , .A1( us23_n779 ) , .B1( us23_n790 ) , .B2( us23_n816 ) );
  OAI22_X1 us23_U196 (.ZN( us23_n636 ) , .A1( us23_n698 ) , .B2( us23_n727 ) , .A2( us23_n761 ) , .B1( us23_n815 ) );
  NOR2_X1 us23_U197 (.A1( us23_n696 ) , .ZN( us23_n769 ) , .A2( us23_n814 ) );
  NOR2_X1 us23_U198 (.ZN( us23_n714 ) , .A1( us23_n804 ) , .A2( us23_n816 ) );
  NOR2_X1 us23_U199 (.ZN( us23_n717 ) , .A2( us23_n723 ) , .A1( us23_n743 ) );
  NOR4_X1 us23_U20 (.ZN( us23_n478 ) , .A1( us23_n519 ) , .A4( us23_n556 ) , .A3( us23_n581 ) , .A2( us23_n629 ) );
  NOR2_X1 us23_U200 (.ZN( us23_n545 ) , .A2( us23_n779 ) , .A1( us23_n813 ) );
  INV_X1 us23_U201 (.A( us23_n749 ) , .ZN( us23_n841 ) );
  NOR2_X1 us23_U202 (.ZN( us23_n651 ) , .A1( us23_n668 ) , .A2( us23_n813 ) );
  NOR2_X1 us23_U203 (.ZN( us23_n531 ) , .A2( us23_n748 ) , .A1( us23_n749 ) );
  NOR2_X1 us23_U204 (.ZN( us23_n576 ) , .A2( us23_n698 ) , .A1( us23_n813 ) );
  NOR2_X1 us23_U205 (.ZN( us23_n599 ) , .A2( us23_n696 ) , .A1( us23_n783 ) );
  NOR2_X1 us23_U206 (.A1( us23_n668 ) , .ZN( us23_n672 ) , .A2( us23_n743 ) );
  NOR2_X1 us23_U207 (.ZN( us23_n601 ) , .A1( us23_n668 ) , .A2( us23_n802 ) );
  NOR2_X1 us23_U208 (.A1( us23_n668 ) , .ZN( us23_n687 ) , .A2( us23_n815 ) );
  NOR2_X1 us23_U209 (.ZN( us23_n628 ) , .A2( us23_n727 ) , .A1( us23_n784 ) );
  NOR4_X1 us23_U21 (.A4( us23_n540 ) , .A3( us23_n541 ) , .A2( us23_n542 ) , .ZN( us23_n549 ) , .A1( us23_n687 ) );
  NOR2_X1 us23_U210 (.ZN( us23_n614 ) , .A1( us23_n784 ) , .A2( us23_n814 ) );
  NOR2_X1 us23_U211 (.A2( us23_n743 ) , .ZN( us23_n754 ) , .A1( us23_n804 ) );
  NOR2_X1 us23_U212 (.A1( us23_n668 ) , .ZN( us23_n765 ) , .A2( us23_n812 ) );
  NOR2_X1 us23_U213 (.ZN( us23_n734 ) , .A2( us23_n802 ) , .A1( us23_n804 ) );
  NOR2_X1 us23_U214 (.A1( us23_n698 ) , .ZN( us23_n767 ) , .A2( us23_n812 ) );
  NOR2_X1 us23_U215 (.A2( us23_n743 ) , .ZN( us23_n768 ) , .A1( us23_n811 ) );
  NOR2_X1 us23_U216 (.ZN( us23_n530 ) , .A2( us23_n779 ) , .A1( us23_n815 ) );
  NOR2_X1 us23_U217 (.ZN( us23_n526 ) , .A1( us23_n668 ) , .A2( us23_n778 ) );
  NOR2_X1 us23_U218 (.ZN( us23_n540 ) , .A2( us23_n696 ) , .A1( us23_n698 ) );
  NOR2_X1 us23_U219 (.ZN( us23_n598 ) , .A2( us23_n790 ) , .A1( us23_n815 ) );
  NOR2_X1 us23_U22 (.ZN( us23_n679 ) , .A2( us23_n833 ) , .A1( us23_n838 ) );
  NOR2_X1 us23_U220 (.ZN( us23_n627 ) , .A2( us23_n668 ) , .A1( us23_n784 ) );
  NOR2_X1 us23_U221 (.ZN( us23_n600 ) , .A2( us23_n779 ) , .A1( us23_n802 ) );
  INV_X1 us23_U222 (.A( us23_n746 ) , .ZN( us23_n833 ) );
  NOR2_X1 us23_U223 (.ZN( us23_n610 ) , .A2( us23_n779 ) , .A1( us23_n805 ) );
  NOR2_X1 us23_U224 (.ZN( us23_n527 ) , .A2( us23_n723 ) , .A1( us23_n802 ) );
  NOR2_X1 us23_U225 (.ZN( us23_n609 ) , .A1( us23_n783 ) , .A2( us23_n815 ) );
  INV_X1 us23_U226 (.A( us23_n791 ) , .ZN( us23_n850 ) );
  NOR2_X1 us23_U227 (.ZN( us23_n650 ) , .A1( us23_n783 ) , .A2( us23_n787 ) );
  NOR2_X1 us23_U228 (.A2( us23_n707 ) , .A1( us23_n749 ) , .ZN( us23_n770 ) );
  NOR2_X1 us23_U229 (.ZN( us23_n666 ) , .A1( us23_n749 ) , .A2( us23_n814 ) );
  AOI222_X1 us23_U23 (.ZN( us23_n468 ) , .B1( us23_n831 ) , .A1( us23_n838 ) , .C1( us23_n841 ) , .C2( us23_n850 ) , .A2( us23_n854 ) , .B2( us23_n864 ) );
  NOR2_X1 us23_U230 (.ZN( us23_n554 ) , .A1( us23_n749 ) , .A2( us23_n790 ) );
  NOR2_X1 us23_U231 (.ZN( us23_n507 ) , .A2( us23_n779 ) , .A1( us23_n784 ) );
  NOR2_X1 us23_U232 (.ZN( us23_n542 ) , .A2( us23_n707 ) , .A1( us23_n784 ) );
  NOR2_X1 us23_U233 (.ZN( us23_n663 ) , .A1( us23_n784 ) , .A2( us23_n790 ) );
  OAI22_X1 us23_U234 (.B1( us23_n439 ) , .ZN( us23_n443 ) , .A2( us23_n727 ) , .A1( us23_n743 ) , .B2( us23_n748 ) );
  NOR3_X1 us23_U235 (.ZN( us23_n439 ) , .A2( us23_n835 ) , .A3( us23_n836 ) , .A1( us23_n845 ) );
  NOR2_X1 us23_U236 (.A2( us23_n696 ) , .ZN( us23_n715 ) , .A1( us23_n791 ) );
  NOR2_X1 us23_U237 (.ZN( us23_n506 ) , .A1( us23_n811 ) , .A2( us23_n816 ) );
  NOR2_X1 us23_U238 (.ZN( us23_n593 ) , .A2( us23_n696 ) , .A1( us23_n727 ) );
  NOR2_X1 us23_U239 (.ZN( us23_n661 ) , .A2( us23_n696 ) , .A1( us23_n728 ) );
  NOR4_X1 us23_U24 (.A1( us23_n465 ) , .ZN( us23_n466 ) , .A4( us23_n541 ) , .A2( us23_n553 ) , .A3( us23_n613 ) );
  NOR2_X1 us23_U240 (.ZN( us23_n556 ) , .A1( us23_n791 ) , .A2( us23_n813 ) );
  NOR2_X1 us23_U241 (.ZN( us23_n544 ) , .A1( us23_n748 ) , .A2( us23_n813 ) );
  NOR2_X1 us23_U242 (.ZN( us23_n555 ) , .A1( us23_n761 ) , .A2( us23_n804 ) );
  NOR2_X1 us23_U243 (.ZN( us23_n529 ) , .A2( us23_n743 ) , .A1( us23_n791 ) );
  NOR2_X1 us23_U244 (.A2( us23_n696 ) , .A1( us23_n779 ) , .ZN( us23_n819 ) );
  NOR2_X1 us23_U245 (.ZN( us23_n508 ) , .A1( us23_n728 ) , .A2( us23_n778 ) );
  NOR2_X1 us23_U246 (.ZN( us23_n665 ) , .A1( us23_n727 ) , .A2( us23_n802 ) );
  NOR2_X1 us23_U247 (.ZN( us23_n543 ) , .A2( us23_n784 ) , .A1( us23_n791 ) );
  NOR2_X1 us23_U248 (.A1( us23_n748 ) , .ZN( us23_n766 ) , .A2( us23_n802 ) );
  NOR2_X1 us23_U249 (.ZN( us23_n613 ) , .A1( us23_n761 ) , .A2( us23_n811 ) );
  AOI221_X1 us23_U25 (.ZN( us23_n467 ) , .C2( us23_n713 ) , .B2( us23_n830 ) , .C1( us23_n844 ) , .B1( us23_n859 ) , .A( us23_n863 ) );
  NOR2_X1 us23_U250 (.ZN( us23_n515 ) , .A1( us23_n707 ) , .A2( us23_n743 ) );
  NOR2_X1 us23_U251 (.ZN( us23_n630 ) , .A1( us23_n723 ) , .A2( us23_n812 ) );
  NOR2_X1 us23_U252 (.ZN( us23_n569 ) , .A1( us23_n727 ) , .A2( us23_n805 ) );
  NOR2_X1 us23_U253 (.ZN( us23_n557 ) , .A1( us23_n707 ) , .A2( us23_n815 ) );
  INV_X1 us23_U254 (.A( us23_n762 ) , .ZN( us23_n865 ) );
  NOR2_X1 us23_U255 (.ZN( us23_n653 ) , .A1( us23_n727 ) , .A2( us23_n812 ) );
  NOR2_X1 us23_U256 (.ZN( us23_n516 ) , .A1( us23_n707 ) , .A2( us23_n802 ) );
  NOR2_X1 us23_U257 (.ZN( us23_n520 ) , .A1( us23_n789 ) , .A2( us23_n811 ) );
  NOR2_X1 us23_U258 (.ZN( us23_n662 ) , .A1( us23_n728 ) , .A2( us23_n784 ) );
  NOR2_X1 us23_U259 (.ZN( us23_n654 ) , .A1( us23_n789 ) , .A2( us23_n814 ) );
  NOR4_X1 us23_U26 (.A4( us23_n664 ) , .A3( us23_n665 ) , .A2( us23_n666 ) , .A1( us23_n667 ) , .ZN( us23_n675 ) );
  NOR2_X1 us23_U260 (.ZN( us23_n629 ) , .A1( us23_n746 ) , .A2( us23_n814 ) );
  NOR2_X1 us23_U261 (.ZN( us23_n667 ) , .A2( us23_n707 ) , .A1( us23_n789 ) );
  NOR2_X1 us23_U262 (.ZN( us23_n669 ) , .A1( us23_n789 ) , .A2( us23_n804 ) );
  AOI21_X1 us23_U263 (.ZN( us23_n570 ) , .B2( us23_n696 ) , .B1( us23_n805 ) , .A( us23_n811 ) );
  NOR2_X1 us23_U264 (.ZN( us23_n541 ) , .A1( us23_n761 ) , .A2( us23_n790 ) );
  NOR2_X1 us23_U265 (.ZN( us23_n655 ) , .A1( us23_n746 ) , .A2( us23_n779 ) );
  INV_X1 us23_U266 (.A( us23_n805 ) , .ZN( us23_n840 ) );
  NOR2_X1 us23_U267 (.ZN( us23_n608 ) , .A2( us23_n723 ) , .A1( us23_n816 ) );
  AOI21_X1 us23_U268 (.A( us23_n814 ) , .B2( us23_n815 ) , .B1( us23_n816 ) , .ZN( us23_n817 ) );
  AOI21_X1 us23_U269 (.ZN( us23_n625 ) , .B2( us23_n668 ) , .A( us23_n789 ) , .B1( us23_n790 ) );
  NOR4_X1 us23_U27 (.A4( us23_n660 ) , .A3( us23_n661 ) , .A2( us23_n662 ) , .A1( us23_n663 ) , .ZN( us23_n676 ) );
  NOR2_X1 us23_U270 (.ZN( us23_n660 ) , .A1( us23_n728 ) , .A2( us23_n789 ) );
  INV_X1 us23_U271 (.A( us23_n811 ) , .ZN( us23_n853 ) );
  NOR2_X1 us23_U272 (.ZN( us23_n578 ) , .A2( us23_n707 ) , .A1( us23_n729 ) );
  NOR2_X1 us23_U273 (.ZN( us23_n532 ) , .A2( us23_n723 ) , .A1( us23_n729 ) );
  AOI21_X1 us23_U274 (.ZN( us23_n498 ) , .B1( us23_n679 ) , .A( us23_n811 ) , .B2( us23_n815 ) );
  AOI21_X1 us23_U275 (.ZN( us23_n551 ) , .B1( us23_n668 ) , .A( us23_n696 ) , .B2( us23_n804 ) );
  NOR2_X1 us23_U276 (.ZN( us23_n581 ) , .A1( us23_n743 ) , .A2( us23_n814 ) );
  NOR2_X1 us23_U277 (.A2( us23_n707 ) , .A1( us23_n761 ) , .ZN( us23_n793 ) );
  AOI21_X1 us23_U278 (.B1( us23_n624 ) , .ZN( us23_n626 ) , .A( us23_n762 ) , .B2( us23_n813 ) );
  AOI21_X1 us23_U279 (.ZN( us23_n514 ) , .A( us23_n728 ) , .B1( us23_n749 ) , .B2( us23_n802 ) );
  NOR4_X1 us23_U28 (.A3( us23_n672 ) , .A1( us23_n673 ) , .ZN( us23_n674 ) , .A4( us23_n714 ) , .A2( us23_n858 ) );
  AOI21_X1 us23_U280 (.A( us23_n811 ) , .B2( us23_n812 ) , .B1( us23_n813 ) , .ZN( us23_n818 ) );
  AOI21_X1 us23_U281 (.ZN( us23_n477 ) , .B2( us23_n696 ) , .A( us23_n748 ) , .B1( us23_n778 ) );
  AOI21_X1 us23_U282 (.ZN( us23_n509 ) , .B2( us23_n668 ) , .A( us23_n729 ) , .B1( us23_n814 ) );
  NOR2_X1 us23_U283 (.ZN( us23_n505 ) , .A2( us23_n727 ) , .A1( us23_n761 ) );
  AOI21_X1 us23_U284 (.ZN( us23_n591 ) , .B1( us23_n727 ) , .B2( us23_n783 ) , .A( us23_n789 ) );
  NOR2_X1 us23_U285 (.ZN( us23_n518 ) , .A2( us23_n698 ) , .A1( us23_n815 ) );
  AOI21_X1 us23_U286 (.ZN( us23_n592 ) , .B1( us23_n749 ) , .A( us23_n791 ) , .B2( us23_n812 ) );
  AOI21_X1 us23_U287 (.ZN( us23_n649 ) , .A( us23_n778 ) , .B1( us23_n791 ) , .B2( us23_n804 ) );
  NOR2_X1 us23_U288 (.ZN( us23_n580 ) , .A1( us23_n668 ) , .A2( us23_n787 ) );
  NOR2_X1 us23_U289 (.ZN( us23_n519 ) , .A2( us23_n707 ) , .A1( us23_n813 ) );
  NOR4_X1 us23_U29 (.A4( us23_n513 ) , .A3( us23_n514 ) , .A2( us23_n515 ) , .A1( us23_n516 ) , .ZN( us23_n523 ) );
  AOI21_X1 us23_U290 (.ZN( us23_n476 ) , .A( us23_n668 ) , .B1( us23_n749 ) , .B2( us23_n805 ) );
  NOR2_X1 us23_U291 (.ZN( us23_n558 ) , .A2( us23_n790 ) , .A1( us23_n802 ) );
  AOI21_X1 us23_U292 (.ZN( us23_n647 ) , .A( us23_n761 ) , .B2( us23_n783 ) , .B1( us23_n791 ) );
  AOI21_X1 us23_U293 (.ZN( us23_n622 ) , .B1( us23_n698 ) , .A( us23_n778 ) , .B2( us23_n783 ) );
  AOI21_X1 us23_U294 (.ZN( us23_n588 ) , .B2( us23_n698 ) , .B1( us23_n814 ) , .A( us23_n816 ) );
  NOR2_X1 us23_U295 (.ZN( us23_n552 ) , .A2( us23_n743 ) , .A1( us23_n783 ) );
  NOR2_X1 us23_U296 (.ZN( us23_n682 ) , .A2( us23_n698 ) , .A1( us23_n802 ) );
  AOI21_X1 us23_U297 (.B1( us23_n698 ) , .ZN( us23_n699 ) , .A( us23_n731 ) , .B2( us23_n762 ) );
  AOI21_X1 us23_U298 (.ZN( us23_n590 ) , .B2( us23_n762 ) , .A( us23_n784 ) , .B1( us23_n811 ) );
  AOI21_X1 us23_U299 (.ZN( us23_n538 ) , .B2( us23_n811 ) , .A( us23_n813 ) , .B1( us23_n814 ) );
  NOR3_X1 us23_U3 (.ZN( us23_n597 ) , .A1( us23_n607 ) , .A3( us23_n722 ) , .A2( us23_n741 ) );
  AOI222_X1 us23_U30 (.ZN( us23_n524 ) , .A1( us23_n833 ) , .B2( us23_n836 ) , .C1( us23_n843 ) , .C2( us23_n849 ) , .A2( us23_n851 ) , .B1( us23_n865 ) );
  AOI21_X1 us23_U300 (.ZN( us23_n539 ) , .A( us23_n762 ) , .B2( us23_n778 ) , .B1( us23_n816 ) );
  NOR2_X1 us23_U301 (.ZN( us23_n546 ) , .A1( us23_n698 ) , .A2( us23_n743 ) );
  INV_X1 us23_U302 (.A( us23_n812 ) , .ZN( us23_n835 ) );
  INV_X1 us23_U303 (.A( us23_n727 ) , .ZN( us23_n851 ) );
  AOI21_X1 us23_U304 (.ZN( us23_n648 ) , .B1( us23_n728 ) , .B2( us23_n762 ) , .A( us23_n812 ) );
  INV_X1 us23_U305 (.A( us23_n790 ) , .ZN( us23_n872 ) );
  OAI221_X1 us23_U306 (.A( us23_n726 ) , .C2( us23_n727 ) , .B2( us23_n728 ) , .B1( us23_n729 ) , .ZN( us23_n736 ) , .C1( us23_n816 ) );
  AOI22_X1 us23_U307 (.ZN( us23_n726 ) , .B1( us23_n831 ) , .A2( us23_n837 ) , .A1( us23_n862 ) , .B2( us23_n865 ) );
  AOI21_X1 us23_U308 (.ZN( us23_n497 ) , .A( us23_n723 ) , .B2( us23_n761 ) , .B1( us23_n813 ) );
  NOR2_X1 us23_U309 (.ZN( us23_n565 ) , .A2( us23_n696 ) , .A1( us23_n762 ) );
  NOR4_X1 us23_U31 (.A3( us23_n520 ) , .A1( us23_n521 ) , .ZN( us23_n522 ) , .A2( us23_n672 ) , .A4( us23_n768 ) );
  INV_X1 us23_U310 (.A( us23_n698 ) , .ZN( us23_n852 ) );
  AOI21_X1 us23_U311 (.ZN( us23_n568 ) , .B1( us23_n749 ) , .B2( us23_n761 ) , .A( us23_n779 ) );
  AOI21_X1 us23_U312 (.ZN( us23_n513 ) , .A( us23_n778 ) , .B2( us23_n791 ) , .B1( us23_n811 ) );
  NOR2_X1 us23_U313 (.ZN( us23_n579 ) , .A2( us23_n696 ) , .A1( us23_n790 ) );
  NOR2_X1 us23_U314 (.ZN( us23_n684 ) , .A1( us23_n728 ) , .A2( us23_n815 ) );
  AOI21_X1 us23_U315 (.ZN( us23_n563 ) , .B1( us23_n723 ) , .A( us23_n778 ) , .B2( us23_n790 ) );
  AOI21_X1 us23_U316 (.ZN( us23_n496 ) , .A( us23_n778 ) , .B2( us23_n790 ) , .B1( us23_n803 ) );
  INV_X1 us23_U317 (.A( us23_n728 ) , .ZN( us23_n867 ) );
  NOR2_X1 us23_U318 (.ZN( us23_n664 ) , .A1( us23_n779 ) , .A2( us23_n812 ) );
  NOR2_X1 us23_U319 (.ZN( us23_n631 ) , .A2( us23_n696 ) , .A1( us23_n723 ) );
  AOI221_X1 us23_U32 (.A( us23_n780 ) , .ZN( us23_n797 ) , .C2( us23_n836 ) , .B2( us23_n837 ) , .B1( us23_n864 ) , .C1( us23_n865 ) );
  NOR2_X1 us23_U320 (.ZN( us23_n528 ) , .A1( us23_n707 ) , .A2( us23_n778 ) );
  NOR2_X1 us23_U321 (.ZN( us23_n577 ) , .A1( us23_n707 ) , .A2( us23_n812 ) );
  AOI21_X1 us23_U322 (.A( us23_n789 ) , .B2( us23_n790 ) , .B1( us23_n791 ) , .ZN( us23_n792 ) );
  AOI21_X1 us23_U323 (.ZN( us23_n688 ) , .B2( us23_n748 ) , .B1( us23_n762 ) , .A( us23_n805 ) );
  NOR2_X1 us23_U324 (.ZN( us23_n683 ) , .A1( us23_n790 ) , .A2( us23_n812 ) );
  NOR2_X1 us23_U325 (.ZN( us23_n566 ) , .A1( us23_n746 ) , .A2( us23_n804 ) );
  NAND2_X1 us23_U326 (.ZN( us23_n752 ) , .A1( us23_n762 ) , .A2( us23_n804 ) );
  AOI21_X1 us23_U327 (.A( us23_n732 ) , .ZN( us23_n733 ) , .B2( us23_n779 ) , .B1( us23_n791 ) );
  NOR2_X1 us23_U328 (.A2( us23_n812 ) , .A1( us23_n814 ) , .ZN( us23_n820 ) );
  NOR2_X1 us23_U329 (.ZN( us23_n710 ) , .A1( us23_n761 ) , .A2( us23_n762 ) );
  NOR4_X1 us23_U33 (.A4( us23_n792 ) , .A3( us23_n793 ) , .A2( us23_n794 ) , .A1( us23_n795 ) , .ZN( us23_n796 ) );
  NOR2_X1 us23_U330 (.ZN( us23_n641 ) , .A2( us23_n787 ) , .A1( us23_n790 ) );
  NOR2_X1 us23_U331 (.ZN( us23_n582 ) , .A1( us23_n791 ) , .A2( us23_n816 ) );
  NOR2_X1 us23_U332 (.ZN( us23_n681 ) , .A2( us23_n707 ) , .A1( us23_n816 ) );
  NOR2_X1 us23_U333 (.ZN( us23_n533 ) , .A1( us23_n723 ) , .A2( us23_n787 ) );
  AOI21_X1 us23_U334 (.B1( us23_n685 ) , .ZN( us23_n686 ) , .A( us23_n727 ) , .B2( us23_n760 ) );
  INV_X1 us23_U335 (.A( us23_n696 ) , .ZN( us23_n837 ) );
  INV_X1 us23_U336 (.A( us23_n814 ) , .ZN( us23_n854 ) );
  NOR2_X1 us23_U337 (.ZN( us23_n567 ) , .A1( us23_n728 ) , .A2( us23_n761 ) );
  AOI21_X1 us23_U338 (.ZN( us23_n441 ) , .A( us23_n698 ) , .B1( us23_n732 ) , .B2( us23_n749 ) );
  OAI21_X1 us23_U339 (.A( us23_n730 ) , .B1( us23_n731 ) , .ZN( us23_n735 ) , .B2( us23_n804 ) );
  NOR4_X1 us23_U34 (.A4( us23_n775 ) , .A3( us23_n776 ) , .A1( us23_n777 ) , .ZN( us23_n798 ) , .A2( us23_n800 ) );
  OAI21_X1 us23_U340 (.ZN( us23_n730 ) , .A( us23_n832 ) , .B2( us23_n851 ) , .B1( us23_n872 ) );
  OAI21_X1 us23_U341 (.A( us23_n697 ) , .ZN( us23_n701 ) , .B2( us23_n749 ) , .B1( us23_n803 ) );
  OAI21_X1 us23_U342 (.ZN( us23_n697 ) , .B2( us23_n832 ) , .B1( us23_n837 ) , .A( us23_n859 ) );
  OAI21_X1 us23_U343 (.A( us23_n612 ) , .ZN( us23_n615 ) , .B1( us23_n624 ) , .B2( us23_n783 ) );
  INV_X1 us23_U344 (.A( us23_n779 ) , .ZN( us23_n849 ) );
  AOI22_X1 us23_U345 (.A2( us23_n781 ) , .ZN( us23_n782 ) , .B2( us23_n830 ) , .A1( us23_n833 ) , .B1( us23_n862 ) );
  NAND2_X1 us23_U346 (.ZN( us23_n670 ) , .A1( us23_n805 ) , .A2( us23_n815 ) );
  OAI21_X1 us23_U347 (.A( us23_n786 ) , .B2( us23_n787 ) , .B1( us23_n788 ) , .ZN( us23_n794 ) );
  OAI21_X1 us23_U348 (.ZN( us23_n786 ) , .A( us23_n838 ) , .B1( us23_n862 ) , .B2( us23_n872 ) );
  NAND2_X1 us23_U349 (.A1( us23_n728 ) , .A2( us23_n783 ) , .ZN( us23_n810 ) );
  NOR4_X1 us23_U35 (.A4( us23_n733 ) , .A3( us23_n734 ) , .A2( us23_n735 ) , .A1( us23_n736 ) , .ZN( us23_n737 ) );
  NOR2_X1 us23_U350 (.ZN( us23_n483 ) , .A1( us23_n787 ) , .A2( us23_n804 ) );
  AOI21_X1 us23_U351 (.ZN( us23_n442 ) , .B1( us23_n788 ) , .B2( us23_n790 ) , .A( us23_n813 ) );
  NAND2_X1 us23_U352 (.A2( us23_n761 ) , .A1( us23_n805 ) , .ZN( us23_n809 ) );
  NOR2_X1 us23_U353 (.ZN( us23_n469 ) , .A2( us23_n778 ) , .A1( us23_n814 ) );
  NAND2_X1 us23_U354 (.A1( us23_n698 ) , .A2( us23_n728 ) , .ZN( us23_n781 ) );
  NOR2_X1 us23_U355 (.ZN( us23_n711 ) , .A2( us23_n723 ) , .A1( us23_n789 ) );
  INV_X1 us23_U356 (.A( us23_n784 ) , .ZN( us23_n845 ) );
  NOR2_X1 us23_U357 (.ZN( us23_n525 ) , .A1( us23_n723 ) , .A2( us23_n749 ) );
  NOR2_X1 us23_U358 (.ZN( us23_n517 ) , .A1( us23_n707 ) , .A2( us23_n787 ) );
  INV_X1 us23_U359 (.A( us23_n816 ) , .ZN( us23_n843 ) );
  AOI211_X1 us23_U36 (.B( us23_n724 ) , .A( us23_n725 ) , .ZN( us23_n738 ) , .C1( us23_n842 ) , .C2( us23_n854 ) );
  NAND2_X1 us23_U360 (.ZN( us23_n713 ) , .A1( us23_n727 ) , .A2( us23_n779 ) );
  INV_X1 us23_U361 (.A( us23_n723 ) , .ZN( us23_n855 ) );
  AND2_X1 us23_U362 (.ZN( us23_n731 ) , .A1( us23_n778 ) , .A2( us23_n784 ) );
  NAND2_X1 us23_U363 (.A2( us23_n460 ) , .A1( us23_n470 ) , .ZN( us23_n696 ) );
  NAND2_X1 us23_U364 (.A1( us23_n451 ) , .A2( us23_n464 ) , .ZN( us23_n668 ) );
  NAND2_X1 us23_U365 (.A1( us23_n450 ) , .A2( us23_n470 ) , .ZN( us23_n815 ) );
  NAND2_X1 us23_U366 (.A1( us23_n452 ) , .A2( us23_n460 ) , .ZN( us23_n743 ) );
  NAND2_X1 us23_U367 (.A1( us23_n454 ) , .A2( us23_n470 ) , .ZN( us23_n802 ) );
  NAND2_X1 us23_U368 (.A1( us23_n450 ) , .A2( us23_n453 ) , .ZN( us23_n813 ) );
  NAND2_X1 us23_U369 (.A1( us23_n454 ) , .A2( us23_n461 ) , .ZN( us23_n749 ) );
  NOR3_X1 us23_U37 (.A3( us23_n721 ) , .A1( us23_n722 ) , .ZN( us23_n739 ) , .A2( us23_n740 ) );
  NAND2_X1 us23_U370 (.A1( us23_n446 ) , .A2( us23_n448 ) , .ZN( us23_n804 ) );
  NAND2_X1 us23_U371 (.A1( us23_n453 ) , .A2( us23_n460 ) , .ZN( us23_n812 ) );
  NAND2_X1 us23_U372 (.A2( us23_n440 ) , .A1( us23_n446 ) , .ZN( us23_n783 ) );
  NAND2_X1 us23_U373 (.A2( us23_n453 ) , .A1( us23_n471 ) , .ZN( us23_n778 ) );
  NAND2_X1 us23_U374 (.A2( us23_n452 ) , .A1( us23_n454 ) , .ZN( us23_n805 ) );
  NAND2_X1 us23_U375 (.A1( us23_n452 ) , .A2( us23_n471 ) , .ZN( us23_n784 ) );
  NAND2_X1 us23_U376 (.A1( us23_n440 ) , .A2( us23_n459 ) , .ZN( us23_n698 ) );
  NAND2_X1 us23_U377 (.A2( us23_n463 ) , .A1( us23_n464 ) , .ZN( us23_n811 ) );
  NAND2_X1 us23_U378 (.A2( us23_n448 ) , .A1( us23_n451 ) , .ZN( us23_n762 ) );
  NAND2_X1 us23_U379 (.A1( us23_n461 ) , .A2( us23_n471 ) , .ZN( us23_n787 ) );
  NOR4_X1 us23_U38 (.A3( us23_n754 ) , .A2( us23_n755 ) , .A1( us23_n756 ) , .ZN( us23_n757 ) , .A4( us23_n868 ) );
  NAND2_X1 us23_U380 (.A2( us23_n460 ) , .A1( us23_n461 ) , .ZN( us23_n746 ) );
  NOR2_X1 us23_U381 (.ZN( us23_n464 ) , .A2( us23_n846 ) , .A1( us23_n847 ) );
  NOR2_X1 us23_U382 (.ZN( us23_n452 ) , .A1( us23_n825 ) , .A2( us23_n826 ) );
  NAND2_X1 us23_U383 (.A1( us23_n450 ) , .A2( us23_n461 ) , .ZN( us23_n789 ) );
  NOR2_X1 us23_U384 (.ZN( us23_n450 ) , .A1( us23_n827 ) , .A2( us23_n828 ) );
  NAND2_X2 us23_U385 (.A2( us23_n447 ) , .A1( us23_n463 ) , .ZN( us23_n814 ) );
  NAND2_X1 us23_U386 (.A2( us23_n453 ) , .A1( us23_n454 ) , .ZN( us23_n729 ) );
  NAND2_X2 us23_U387 (.A2( us23_n440 ) , .A1( us23_n451 ) , .ZN( us23_n790 ) );
  NAND2_X2 us23_U388 (.A1( us23_n448 ) , .A2( us23_n459 ) , .ZN( us23_n791 ) );
  NAND2_X2 us23_U389 (.A1( us23_n448 ) , .A2( us23_n463 ) , .ZN( us23_n723 ) );
  AOI211_X1 us23_U39 (.B( us23_n744 ) , .A( us23_n745 ) , .ZN( us23_n758 ) , .C1( us23_n831 ) , .C2( us23_n852 ) );
  NAND2_X2 us23_U390 (.A1( us23_n440 ) , .A2( us23_n463 ) , .ZN( us23_n707 ) );
  NAND2_X2 us23_U391 (.A2( us23_n470 ) , .A1( us23_n471 ) , .ZN( us23_n816 ) );
  NAND2_X2 us23_U392 (.A2( us23_n459 ) , .A1( us23_n464 ) , .ZN( us23_n779 ) );
  NOR2_X1 us23_U393 (.ZN( us23_n446 ) , .A2( us23_n848 ) , .A1( us23_n857 ) );
  NAND2_X1 us23_U394 (.A1( us23_n446 ) , .A2( us23_n447 ) , .ZN( us23_n785 ) );
  NAND2_X1 us23_U395 (.A2( us23_n447 ) , .A1( us23_n459 ) , .ZN( us23_n727 ) );
  NAND2_X1 us23_U396 (.A2( us23_n447 ) , .A1( us23_n451 ) , .ZN( us23_n728 ) );
  NOR2_X1 us23_U397 (.A2( sa23_5 ) , .ZN( us23_n447 ) , .A1( us23_n846 ) );
  NOR2_X1 us23_U398 (.A2( sa23_7 ) , .ZN( us23_n459 ) , .A1( us23_n848 ) );
  NOR2_X1 us23_U399 (.A2( sa23_6 ) , .A1( sa23_7 ) , .ZN( us23_n463 ) );
  NOR3_X1 us23_U4 (.A3( us23_n799 ) , .A2( us23_n800 ) , .A1( us23_n801 ) , .ZN( us23_n824 ) );
  NOR3_X1 us23_U40 (.A3( us23_n740 ) , .A2( us23_n741 ) , .A1( us23_n742 ) , .ZN( us23_n759 ) );
  NOR2_X1 us23_U400 (.A2( sa23_4 ) , .ZN( us23_n448 ) , .A1( us23_n847 ) );
  NOR2_X1 us23_U401 (.A2( sa23_4 ) , .A1( sa23_5 ) , .ZN( us23_n440 ) );
  NOR2_X1 us23_U402 (.A2( sa23_6 ) , .ZN( us23_n451 ) , .A1( us23_n857 ) );
  NOR2_X1 us23_U403 (.A2( sa23_1 ) , .ZN( us23_n470 ) , .A1( us23_n825 ) );
  NOR2_X1 us23_U404 (.A2( sa23_2 ) , .A1( sa23_3 ) , .ZN( us23_n471 ) );
  NOR2_X1 us23_U405 (.A2( sa23_2 ) , .ZN( us23_n460 ) , .A1( us23_n828 ) );
  NOR2_X1 us23_U406 (.A2( sa23_0 ) , .ZN( us23_n453 ) , .A1( us23_n826 ) );
  NOR2_X1 us23_U407 (.A2( sa23_0 ) , .A1( sa23_1 ) , .ZN( us23_n461 ) );
  NOR2_X1 us23_U408 (.A2( sa23_3 ) , .ZN( us23_n454 ) , .A1( us23_n827 ) );
  INV_X1 us23_U409 (.A( sa23_6 ) , .ZN( us23_n848 ) );
  NAND4_X1 us23_U41 (.ZN( sa21_sr_3 ) , .A4( us23_n703 ) , .A3( us23_n704 ) , .A2( us23_n705 ) , .A1( us23_n706 ) );
  INV_X1 us23_U410 (.A( sa23_4 ) , .ZN( us23_n846 ) );
  INV_X1 us23_U411 (.A( sa23_1 ) , .ZN( us23_n826 ) );
  INV_X1 us23_U412 (.A( sa23_3 ) , .ZN( us23_n828 ) );
  INV_X1 us23_U413 (.A( sa23_2 ) , .ZN( us23_n827 ) );
  INV_X1 us23_U414 (.A( sa23_0 ) , .ZN( us23_n825 ) );
  INV_X1 us23_U415 (.A( sa23_7 ) , .ZN( us23_n857 ) );
  INV_X1 us23_U416 (.A( sa23_5 ) , .ZN( us23_n847 ) );
  OAI221_X1 us23_U417 (.A( us23_n782 ) , .C2( us23_n783 ) , .B2( us23_n784 ) , .B1( us23_n785 ) , .ZN( us23_n795 ) , .C1( us23_n812 ) );
  OAI222_X1 us23_U418 (.B2( us23_n746 ) , .B1( us23_n747 ) , .A2( us23_n748 ) , .ZN( us23_n756 ) , .C2( us23_n804 ) , .C1( us23_n813 ) , .A1( us23_n816 ) );
  AOI21_X1 us23_U419 (.ZN( us23_n499 ) , .A( us23_n696 ) , .B1( us23_n707 ) , .B2( us23_n785 ) );
  NOR4_X1 us23_U42 (.A4( us23_n699 ) , .A3( us23_n700 ) , .A2( us23_n701 ) , .A1( us23_n702 ) , .ZN( us23_n703 ) );
  OAI221_X1 us23_U420 (.A( us23_n695 ) , .ZN( us23_n702 ) , .C2( us23_n783 ) , .C1( us23_n784 ) , .B1( us23_n785 ) , .B2( us23_n805 ) );
  OAI22_X1 us23_U421 (.ZN( us23_n589 ) , .B1( us23_n729 ) , .B2( us23_n748 ) , .A2( us23_n785 ) , .A1( us23_n802 ) );
  OAI222_X1 us23_U422 (.ZN( us23_n504 ) , .C2( us23_n624 ) , .B2( us23_n646 ) , .B1( us23_n746 ) , .A2( us23_n747 ) , .C1( us23_n804 ) , .A1( us23_n805 ) );
  NOR2_X1 us23_U423 (.ZN( us23_n611 ) , .A1( us23_n778 ) , .A2( us23_n785 ) );
  OAI222_X1 us23_U424 (.ZN( us23_n616 ) , .B1( us23_n696 ) , .C1( us23_n723 ) , .C2( us23_n746 ) , .B2( us23_n785 ) , .A2( us23_n791 ) , .A1( us23_n815 ) );
  NAND2_X1 us23_U425 (.A2( us23_n748 ) , .A1( us23_n785 ) , .ZN( us23_n808 ) );
  AOI21_X1 us23_U426 (.ZN( us23_n575 ) , .B2( us23_n723 ) , .B1( us23_n747 ) , .A( us23_n784 ) );
  NOR2_X1 us23_U427 (.ZN( us23_n716 ) , .A2( us23_n743 ) , .A1( us23_n785 ) );
  NOR2_X1 us23_U428 (.ZN( us23_n652 ) , .A1( us23_n761 ) , .A2( us23_n785 ) );
  NOR2_X1 us23_U429 (.ZN( us23_n553 ) , .A1( us23_n785 ) , .A2( us23_n812 ) );
  AOI211_X1 us23_U43 (.B( us23_n693 ) , .A( us23_n694 ) , .ZN( us23_n704 ) , .C2( us23_n830 ) , .C1( us23_n850 ) );
  NOR2_X1 us23_U430 (.ZN( us23_n700 ) , .A2( us23_n785 ) , .A1( us23_n816 ) );
  NOR2_X1 us23_U431 (.A1( us23_n729 ) , .ZN( us23_n764 ) , .A2( us23_n785 ) );
  NAND2_X1 us23_U432 (.ZN( sa21_sr_2 ) , .A1( us23_n438 ) , .A2( us23_n644 ) );
  NOR3_X1 us23_U433 (.A2( us23_n606 ) , .A1( us23_n607 ) , .ZN( us23_n645 ) , .A3( us23_n721 ) );
  AOI222_X1 us23_U434 (.B2( us23_n637 ) , .ZN( us23_n643 ) , .B1( us23_n840 ) , .A1( us23_n841 ) , .C2( us23_n845 ) , .C1( us23_n862 ) , .A2( us23_n864 ) );
  NOR4_X1 us23_U435 (.A4( us23_n638 ) , .A3( us23_n639 ) , .A2( us23_n640 ) , .A1( us23_n641 ) , .ZN( us23_n642 ) );
  AOI211_X1 us23_U436 (.A( us23_n636 ) , .ZN( us23_n644 ) , .B( us23_n742 ) , .C2( us23_n838 ) , .C1( us23_n853 ) );
  NAND3_X1 us23_U437 (.ZN( sa21_sr_6 ) , .A3( us23_n796 ) , .A2( us23_n797 ) , .A1( us23_n798 ) );
  NAND3_X1 us23_U438 (.ZN( sa21_sr_5 ) , .A3( us23_n757 ) , .A2( us23_n758 ) , .A1( us23_n759 ) );
  NAND3_X1 us23_U439 (.ZN( sa21_sr_4 ) , .A3( us23_n737 ) , .A2( us23_n738 ) , .A1( us23_n739 ) );
  NOR2_X1 us23_U44 (.ZN( us23_n706 ) , .A2( us23_n775 ) , .A1( us23_n799 ) );
  NAND3_X1 us23_U440 (.A3( us23_n674 ) , .A2( us23_n675 ) , .A1( us23_n676 ) , .ZN( us23_n806 ) );
  NAND3_X1 us23_U441 (.ZN( us23_n637 ) , .A3( us23_n707 ) , .A2( us23_n723 ) , .A1( us23_n791 ) );
  NAND3_X1 us23_U442 (.A3( us23_n617 ) , .A2( us23_n618 ) , .A1( us23_n619 ) , .ZN( us23_n724 ) );
  NAND3_X1 us23_U443 (.A3( us23_n584 ) , .A2( us23_n585 ) , .A1( us23_n586 ) , .ZN( us23_n620 ) );
  NAND3_X1 us23_U444 (.ZN( us23_n564 ) , .A3( us23_n679 ) , .A2( us23_n749 ) , .A1( us23_n784 ) );
  NAND3_X1 us23_U445 (.A3( us23_n522 ) , .A2( us23_n523 ) , .A1( us23_n524 ) , .ZN( us23_n741 ) );
  NAND3_X1 us23_U446 (.A3( us23_n511 ) , .A1( us23_n512 ) , .ZN( us23_n607 ) , .A2( us23_n870 ) );
  NAND3_X1 us23_U447 (.A3( us23_n466 ) , .A2( us23_n467 ) , .A1( us23_n468 ) , .ZN( us23_n776 ) );
  NAND4_X1 us23_U448 (.A4( us23_n632 ) , .A3( us23_n633 ) , .A2( us23_n634 ) , .A1( us23_n635 ) , .ZN( us23_n742 ) );
  NOR2_X1 us23_U45 (.ZN( us23_n803 ) , .A1( us23_n853 ) , .A2( us23_n860 ) );
  NAND4_X1 us23_U46 (.ZN( sa21_sr_7 ) , .A4( us23_n821 ) , .A3( us23_n822 ) , .A2( us23_n823 ) , .A1( us23_n824 ) );
  AOI222_X1 us23_U47 (.C2( us23_n808 ) , .B2( us23_n809 ) , .A2( us23_n810 ) , .ZN( us23_n822 ) , .C1( us23_n831 ) , .A1( us23_n838 ) , .B1( us23_n852 ) );
  NOR4_X1 us23_U48 (.A4( us23_n817 ) , .A3( us23_n818 ) , .A2( us23_n819 ) , .A1( us23_n820 ) , .ZN( us23_n821 ) );
  AOI211_X1 us23_U49 (.B( us23_n806 ) , .A( us23_n807 ) , .ZN( us23_n823 ) , .C1( us23_n841 ) , .C2( us23_n849 ) );
  NOR3_X1 us23_U5 (.ZN( us23_n503 ) , .A2( us23_n678 ) , .A3( us23_n776 ) , .A1( us23_n875 ) );
  NAND4_X1 us23_U50 (.ZN( sa21_sr_0 ) , .A4( us23_n500 ) , .A3( us23_n501 ) , .A2( us23_n502 ) , .A1( us23_n503 ) );
  NOR4_X1 us23_U51 (.A4( us23_n497 ) , .A3( us23_n498 ) , .A2( us23_n499 ) , .ZN( us23_n500 ) , .A1( us23_n526 ) );
  AOI221_X1 us23_U52 (.A( us23_n496 ) , .ZN( us23_n501 ) , .B2( us23_n842 ) , .C1( us23_n845 ) , .C2( us23_n859 ) , .B1( us23_n861 ) );
  AOI211_X1 us23_U53 (.A( us23_n495 ) , .ZN( us23_n502 ) , .B( us23_n801 ) , .C2( us23_n838 ) , .C1( us23_n850 ) );
  AND3_X1 us23_U54 (.ZN( us23_n438 ) , .A2( us23_n642 ) , .A3( us23_n643 ) , .A1( us23_n645 ) );
  NAND4_X1 us23_U55 (.ZN( sa21_sr_1 ) , .A4( us23_n594 ) , .A3( us23_n595 ) , .A2( us23_n596 ) , .A1( us23_n597 ) );
  NOR4_X1 us23_U56 (.A4( us23_n590 ) , .A3( us23_n591 ) , .A2( us23_n592 ) , .A1( us23_n593 ) , .ZN( us23_n594 ) );
  AOI211_X1 us23_U57 (.B( us23_n588 ) , .A( us23_n589 ) , .ZN( us23_n595 ) , .C2( us23_n810 ) , .C1( us23_n832 ) );
  AOI211_X1 us23_U58 (.A( us23_n587 ) , .ZN( us23_n596 ) , .B( us23_n620 ) , .C1( us23_n844 ) , .C2( us23_n854 ) );
  NOR2_X1 us23_U59 (.ZN( us23_n624 ) , .A2( us23_n835 ) , .A1( us23_n838 ) );
  INV_X1 us23_U6 (.A( us23_n705 ) , .ZN( us23_n875 ) );
  NOR4_X1 us23_U60 (.A4( us23_n628 ) , .A3( us23_n629 ) , .A2( us23_n630 ) , .A1( us23_n631 ) , .ZN( us23_n632 ) );
  AOI211_X1 us23_U61 (.B( us23_n622 ) , .A( us23_n623 ) , .ZN( us23_n634 ) , .C2( us23_n835 ) , .C1( us23_n862 ) );
  NOR4_X1 us23_U62 (.A4( us23_n625 ) , .A3( us23_n626 ) , .A2( us23_n627 ) , .ZN( us23_n633 ) , .A1( us23_n663 ) );
  NAND4_X1 us23_U63 (.A4( us23_n656 ) , .A3( us23_n657 ) , .A2( us23_n658 ) , .A1( us23_n659 ) , .ZN( us23_n799 ) );
  NOR3_X1 us23_U64 (.A3( us23_n650 ) , .A2( us23_n651 ) , .A1( us23_n652 ) , .ZN( us23_n657 ) );
  NOR3_X1 us23_U65 (.A3( us23_n647 ) , .A2( us23_n648 ) , .A1( us23_n649 ) , .ZN( us23_n658 ) );
  NOR3_X1 us23_U66 (.A3( us23_n653 ) , .A2( us23_n654 ) , .A1( us23_n655 ) , .ZN( us23_n656 ) );
  NAND4_X1 us23_U67 (.A4( us23_n771 ) , .A3( us23_n772 ) , .A2( us23_n773 ) , .A1( us23_n774 ) , .ZN( us23_n800 ) );
  NOR3_X1 us23_U68 (.A3( us23_n764 ) , .A2( us23_n765 ) , .A1( us23_n766 ) , .ZN( us23_n772 ) );
  NOR4_X1 us23_U69 (.A4( us23_n767 ) , .A3( us23_n768 ) , .A2( us23_n769 ) , .A1( us23_n770 ) , .ZN( us23_n771 ) );
  NOR3_X1 us23_U7 (.A3( us23_n620 ) , .A2( us23_n621 ) , .ZN( us23_n635 ) , .A1( us23_n724 ) );
  AOI222_X1 us23_U70 (.ZN( us23_n774 ) , .A1( us23_n829 ) , .C1( us23_n833 ) , .B2( us23_n840 ) , .A2( us23_n849 ) , .B1( us23_n860 ) , .C2( us23_n872 ) );
  NOR4_X1 us23_U71 (.A4( us23_n576 ) , .A3( us23_n577 ) , .A2( us23_n578 ) , .ZN( us23_n585 ) , .A1( us23_n682 ) );
  NOR4_X1 us23_U72 (.A1( us23_n583 ) , .ZN( us23_n584 ) , .A3( us23_n651 ) , .A2( us23_n661 ) , .A4( us23_n766 ) );
  AOI221_X1 us23_U73 (.A( us23_n575 ) , .ZN( us23_n586 ) , .B2( us23_n830 ) , .C2( us23_n842 ) , .B1( us23_n853 ) , .C1( us23_n860 ) );
  NOR2_X1 us23_U74 (.ZN( us23_n760 ) , .A1( us23_n832 ) , .A2( us23_n833 ) );
  NAND4_X1 us23_U75 (.A4( us23_n455 ) , .A3( us23_n456 ) , .A2( us23_n457 ) , .A1( us23_n458 ) , .ZN( us23_n678 ) );
  NOR3_X1 us23_U76 (.ZN( us23_n456 ) , .A3( us23_n529 ) , .A1( us23_n554 ) , .A2( us23_n569 ) );
  NOR4_X1 us23_U77 (.ZN( us23_n457 ) , .A2( us23_n508 ) , .A1( us23_n598 ) , .A4( us23_n627 ) , .A3( us23_n710 ) );
  NOR4_X1 us23_U78 (.ZN( us23_n455 ) , .A2( us23_n516 ) , .A1( us23_n542 ) , .A3( us23_n578 ) , .A4( us23_n614 ) );
  NAND4_X1 us23_U79 (.A4( us23_n602 ) , .A3( us23_n603 ) , .A2( us23_n604 ) , .A1( us23_n605 ) , .ZN( us23_n721 ) );
  NOR2_X1 us23_U8 (.ZN( us23_n574 ) , .A1( us23_n621 ) , .A2( us23_n744 ) );
  NOR3_X1 us23_U80 (.A1( us23_n598 ) , .ZN( us23_n603 ) , .A3( us23_n662 ) , .A2( us23_n769 ) );
  NOR4_X1 us23_U81 (.A3( us23_n599 ) , .A2( us23_n600 ) , .A1( us23_n601 ) , .ZN( us23_n602 ) , .A4( us23_n654 ) );
  AOI222_X1 us23_U82 (.ZN( us23_n605 ) , .A1( us23_n829 ) , .C2( us23_n836 ) , .B1( us23_n841 ) , .A2( us23_n855 ) , .B2( us23_n860 ) , .C1( us23_n867 ) );
  NAND4_X1 us23_U83 (.A4( us23_n534 ) , .A3( us23_n535 ) , .A2( us23_n536 ) , .A1( us23_n537 ) , .ZN( us23_n621 ) );
  NOR4_X1 us23_U84 (.A4( us23_n525 ) , .A2( us23_n526 ) , .A1( us23_n527 ) , .ZN( us23_n537 ) , .A3( us23_n700 ) );
  NOR4_X1 us23_U85 (.A1( us23_n530 ) , .ZN( us23_n535 ) , .A2( us23_n653 ) , .A4( us23_n667 ) , .A3( us23_n764 ) );
  NOR4_X1 us23_U86 (.A4( us23_n528 ) , .A3( us23_n529 ) , .ZN( us23_n536 ) , .A2( us23_n683 ) , .A1( us23_n793 ) );
  NOR2_X1 us23_U87 (.ZN( us23_n685 ) , .A1( us23_n830 ) , .A2( us23_n831 ) );
  NAND4_X1 us23_U88 (.A4( us23_n547 ) , .A3( us23_n548 ) , .A2( us23_n549 ) , .A1( us23_n550 ) , .ZN( us23_n744 ) );
  NOR3_X1 us23_U89 (.ZN( us23_n548 ) , .A2( us23_n650 ) , .A1( us23_n666 ) , .A3( us23_n770 ) );
  NOR2_X1 us23_U9 (.A1( us23_n677 ) , .ZN( us23_n692 ) , .A2( us23_n806 ) );
  AOI211_X1 us23_U90 (.B( us23_n538 ) , .A( us23_n539 ) , .ZN( us23_n550 ) , .C2( us23_n838 ) , .C1( us23_n850 ) );
  NOR4_X1 us23_U91 (.A4( us23_n543 ) , .A3( us23_n544 ) , .A2( us23_n545 ) , .A1( us23_n546 ) , .ZN( us23_n547 ) );
  NAND4_X1 us23_U92 (.A4( us23_n478 ) , .A3( us23_n479 ) , .A2( us23_n480 ) , .A1( us23_n481 ) , .ZN( us23_n693 ) );
  NOR3_X1 us23_U93 (.ZN( us23_n479 ) , .A2( us23_n507 ) , .A3( us23_n600 ) , .A1( us23_n609 ) );
  AOI211_X1 us23_U94 (.B( us23_n476 ) , .A( us23_n477 ) , .ZN( us23_n481 ) , .C2( us23_n832 ) , .C1( us23_n860 ) );
  NOR4_X1 us23_U95 (.ZN( us23_n480 ) , .A3( us23_n531 ) , .A4( us23_n544 ) , .A2( us23_n566 ) , .A1( us23_n716 ) );
  NOR4_X1 us23_U96 (.ZN( us23_n619 ) , .A1( us23_n655 ) , .A3( us23_n665 ) , .A4( us23_n681 ) , .A2( us23_n765 ) );
  NOR4_X1 us23_U97 (.A4( us23_n608 ) , .A3( us23_n609 ) , .A2( us23_n610 ) , .A1( us23_n611 ) , .ZN( us23_n618 ) );
  NOR4_X1 us23_U98 (.A4( us23_n613 ) , .A3( us23_n614 ) , .A2( us23_n615 ) , .A1( us23_n616 ) , .ZN( us23_n617 ) );
  NAND4_X1 us23_U99 (.A4( us23_n484 ) , .A3( us23_n485 ) , .A2( us23_n486 ) , .A1( us23_n487 ) , .ZN( us23_n777 ) );
  NOR2_X1 us30_U10 (.ZN( us30_n575 ) , .A1( us30_n622 ) , .A2( us30_n745 ) );
  NOR2_X1 us30_U100 (.ZN( us30_n647 ) , .A1( us30_n854 ) , .A2( us30_n868 ) );
  NAND4_X1 us30_U101 (.A4( us30_n479 ) , .A3( us30_n480 ) , .A2( us30_n481 ) , .A1( us30_n482 ) , .ZN( us30_n694 ) );
  NOR3_X1 us30_U102 (.ZN( us30_n480 ) , .A2( us30_n508 ) , .A3( us30_n601 ) , .A1( us30_n610 ) );
  AOI211_X1 us30_U103 (.B( us30_n477 ) , .A( us30_n478 ) , .ZN( us30_n482 ) , .C2( us30_n833 ) , .C1( us30_n861 ) );
  NOR4_X1 us30_U104 (.ZN( us30_n481 ) , .A3( us30_n532 ) , .A4( us30_n545 ) , .A2( us30_n567 ) , .A1( us30_n717 ) );
  NAND4_X1 us30_U105 (.A4( us30_n548 ) , .A3( us30_n549 ) , .A2( us30_n550 ) , .A1( us30_n551 ) , .ZN( us30_n745 ) );
  NOR3_X1 us30_U106 (.ZN( us30_n549 ) , .A2( us30_n651 ) , .A1( us30_n667 ) , .A3( us30_n771 ) );
  AOI211_X1 us30_U107 (.B( us30_n539 ) , .A( us30_n540 ) , .ZN( us30_n551 ) , .C2( us30_n839 ) , .C1( us30_n851 ) );
  NOR4_X1 us30_U108 (.A4( us30_n544 ) , .A3( us30_n545 ) , .A2( us30_n546 ) , .A1( us30_n547 ) , .ZN( us30_n548 ) );
  NOR4_X1 us30_U109 (.ZN( us30_n620 ) , .A1( us30_n656 ) , .A3( us30_n666 ) , .A4( us30_n682 ) , .A2( us30_n766 ) );
  NOR2_X1 us30_U11 (.ZN( us30_n495 ) , .A1( us30_n678 ) , .A2( us30_n694 ) );
  NOR4_X1 us30_U110 (.A4( us30_n609 ) , .A3( us30_n610 ) , .A2( us30_n611 ) , .A1( us30_n612 ) , .ZN( us30_n619 ) );
  NOR4_X1 us30_U111 (.A4( us30_n614 ) , .A3( us30_n615 ) , .A2( us30_n616 ) , .A1( us30_n617 ) , .ZN( us30_n618 ) );
  NOR2_X1 us30_U112 (.ZN( us30_n686 ) , .A1( us30_n831 ) , .A2( us30_n832 ) );
  NAND4_X1 us30_U113 (.A4( us30_n485 ) , .A3( us30_n486 ) , .A2( us30_n487 ) , .A1( us30_n488 ) , .ZN( us30_n778 ) );
  NOR4_X1 us30_U114 (.A4( us30_n484 ) , .ZN( us30_n487 ) , .A1( us30_n566 ) , .A2( us30_n581 ) , .A3( us30_n602 ) );
  NOR4_X1 us30_U115 (.ZN( us30_n486 ) , .A1( us30_n507 ) , .A2( us30_n519 ) , .A4( us30_n546 ) , .A3( us30_n611 ) );
  NOR4_X1 us30_U116 (.ZN( us30_n485 ) , .A2( us30_n533 ) , .A1( us30_n558 ) , .A3( us30_n631 ) , .A4( us30_n718 ) );
  NAND4_X1 us30_U117 (.A4( us30_n691 ) , .A3( us30_n692 ) , .A1( us30_n693 ) , .ZN( us30_n776 ) , .A2( us30_n872 ) );
  AOI221_X1 us30_U118 (.A( us30_n681 ) , .ZN( us30_n692 ) , .B2( us30_n840 ) , .C1( us30_n842 ) , .C2( us30_n862 ) , .B1( us30_n865 ) );
  INV_X1 us30_U119 (.A( us30_n679 ) , .ZN( us30_n872 ) );
  NOR2_X1 us30_U12 (.A1( us30_n678 ) , .ZN( us30_n693 ) , .A2( us30_n807 ) );
  NOR4_X1 us30_U120 (.A4( us30_n687 ) , .A3( us30_n688 ) , .A2( us30_n689 ) , .A1( us30_n690 ) , .ZN( us30_n691 ) );
  NAND4_X1 us30_U121 (.A4( us30_n719 ) , .A3( us30_n720 ) , .A2( us30_n721 ) , .ZN( us30_n741 ) , .A1( us30_n857 ) );
  INV_X1 us30_U122 (.A( us30_n709 ) , .ZN( us30_n857 ) );
  AOI221_X1 us30_U123 (.A( us30_n710 ) , .ZN( us30_n721 ) , .C2( us30_n844 ) , .B2( us30_n845 ) , .C1( us30_n861 ) , .B1( us30_n862 ) );
  NOR4_X1 us30_U124 (.A4( us30_n715 ) , .A3( us30_n716 ) , .A2( us30_n717 ) , .A1( us30_n718 ) , .ZN( us30_n719 ) );
  NAND4_X1 us30_U125 (.A4( us30_n473 ) , .A3( us30_n474 ) , .A2( us30_n475 ) , .A1( us30_n476 ) , .ZN( us30_n678 ) );
  NOR4_X1 us30_U126 (.ZN( us30_n475 ) , .A1( us30_n531 ) , .A3( us30_n568 ) , .A4( us30_n600 ) , .A2( us30_n642 ) );
  NOR4_X1 us30_U127 (.A4( us30_n470 ) , .ZN( us30_n476 ) , .A3( us30_n556 ) , .A1( us30_n735 ) , .A2( us30_n755 ) );
  NOR4_X1 us30_U128 (.ZN( us30_n474 ) , .A1( us30_n506 ) , .A3( us30_n544 ) , .A2( us30_n583 ) , .A4( us30_n716 ) );
  NOR2_X1 us30_U129 (.ZN( us30_n733 ) , .A2( us30_n832 ) , .A1( us30_n845 ) );
  NOR3_X1 us30_U13 (.ZN( us30_n504 ) , .A2( us30_n679 ) , .A3( us30_n777 ) , .A1( us30_n876 ) );
  NOR2_X1 us30_U130 (.ZN( us30_n789 ) , .A2( us30_n862 ) , .A1( us30_n868 ) );
  NAND4_X1 us30_U131 (.A4( us30_n573 ) , .A3( us30_n574 ) , .A1( us30_n575 ) , .ZN( us30_n723 ) , .A2( us30_n874 ) );
  AOI221_X1 us30_U132 (.A( us30_n564 ) , .C2( us30_n565 ) , .ZN( us30_n574 ) , .B2( us30_n845 ) , .B1( us30_n852 ) , .C1( us30_n853 ) );
  NOR4_X1 us30_U133 (.A4( us30_n569 ) , .A3( us30_n570 ) , .A2( us30_n571 ) , .A1( us30_n572 ) , .ZN( us30_n573 ) );
  INV_X1 us30_U134 (.A( us30_n607 ) , .ZN( us30_n874 ) );
  NAND4_X1 us30_U135 (.A4( us30_n633 ) , .A3( us30_n634 ) , .A2( us30_n635 ) , .A1( us30_n636 ) , .ZN( us30_n743 ) );
  AOI211_X1 us30_U136 (.B( us30_n623 ) , .A( us30_n624 ) , .ZN( us30_n635 ) , .C2( us30_n836 ) , .C1( us30_n863 ) );
  NOR4_X1 us30_U137 (.A4( us30_n629 ) , .A3( us30_n630 ) , .A2( us30_n631 ) , .A1( us30_n632 ) , .ZN( us30_n633 ) );
  NOR4_X1 us30_U138 (.A4( us30_n626 ) , .A3( us30_n627 ) , .A2( us30_n628 ) , .ZN( us30_n634 ) , .A1( us30_n664 ) );
  NAND4_X1 us30_U139 (.A4( us30_n493 ) , .A3( us30_n494 ) , .A1( us30_n495 ) , .ZN( us30_n802 ) , .A2( us30_n867 ) );
  INV_X1 us30_U14 (.A( us30_n706 ) , .ZN( us30_n876 ) );
  AOI221_X1 us30_U140 (.A( us30_n489 ) , .ZN( us30_n494 ) , .B2( us30_n836 ) , .C2( us30_n841 ) , .C1( us30_n851 ) , .B1( us30_n860 ) );
  INV_X1 us30_U141 (.A( us30_n778 ) , .ZN( us30_n867 ) );
  NOR4_X1 us30_U142 (.A2( us30_n491 ) , .A1( us30_n492 ) , .ZN( us30_n493 ) , .A3( us30_n580 ) , .A4( us30_n612 ) );
  NOR4_X1 us30_U143 (.A4( us30_n734 ) , .A3( us30_n735 ) , .A2( us30_n736 ) , .A1( us30_n737 ) , .ZN( us30_n738 ) );
  AOI211_X1 us30_U144 (.B( us30_n725 ) , .A( us30_n726 ) , .ZN( us30_n739 ) , .C1( us30_n843 ) , .C2( us30_n855 ) );
  NOR3_X1 us30_U145 (.A3( us30_n722 ) , .A1( us30_n723 ) , .ZN( us30_n740 ) , .A2( us30_n741 ) );
  INV_X1 us30_U146 (.A( us30_n762 ) , .ZN( us30_n830 ) );
  OR4_X1 us30_U147 (.A4( us30_n566 ) , .A3( us30_n567 ) , .A2( us30_n568 ) , .ZN( us30_n572 ) , .A1( us30_n665 ) );
  OR4_X1 us30_U148 (.A4( us30_n682 ) , .A3( us30_n683 ) , .A2( us30_n684 ) , .A1( us30_n685 ) , .ZN( us30_n690 ) );
  OR4_X1 us30_U149 (.ZN( us30_n466 ) , .A4( us30_n518 ) , .A3( us30_n529 ) , .A2( us30_n578 ) , .A1( us30_n712 ) );
  INV_X1 us30_U15 (.A( us30_n680 ) , .ZN( us30_n840 ) );
  OR4_X1 us30_U150 (.A4( us30_n518 ) , .A2( us30_n519 ) , .A1( us30_n520 ) , .ZN( us30_n522 ) , .A3( us30_n821 ) );
  OR4_X1 us30_U151 (.ZN( us30_n492 ) , .A4( us30_n534 ) , .A2( us30_n547 ) , .A1( us30_n559 ) , .A3( us30_n632 ) );
  OR4_X1 us30_U152 (.A4( us30_n580 ) , .A3( us30_n581 ) , .A2( us30_n582 ) , .A1( us30_n583 ) , .ZN( us30_n584 ) );
  INV_X1 us30_U153 (.A( us30_n697 ) , .ZN( us30_n838 ) );
  NAND2_X1 us30_U154 (.ZN( us30_n613 ) , .A2( us30_n837 ) , .A1( us30_n873 ) );
  OR3_X1 us30_U155 (.A3( us30_n506 ) , .A2( us30_n507 ) , .A1( us30_n508 ) , .ZN( us30_n511 ) );
  INV_X1 us30_U156 (.A( us30_n754 ) , .ZN( us30_n869 ) );
  OAI21_X1 us30_U157 (.B1( us30_n753 ) , .ZN( us30_n754 ) , .A( us30_n845 ) , .B2( us30_n868 ) );
  INV_X1 us30_U158 (.A( us30_n463 ) , .ZN( us30_n864 ) );
  OAI21_X1 us30_U159 (.ZN( us30_n463 ) , .B1( us30_n809 ) , .A( us30_n834 ) , .B2( us30_n851 ) );
  NOR4_X1 us30_U16 (.A4( us30_n445 ) , .A3( us30_n446 ) , .A2( us30_n516 ) , .A1( us30_n541 ) , .ZN( us30_n706 ) );
  INV_X1 us30_U160 (.A( us30_n672 ) , .ZN( us30_n859 ) );
  AOI21_X1 us30_U161 (.A( us30_n670 ) , .B1( us30_n671 ) , .ZN( us30_n672 ) , .B2( us30_n856 ) );
  OAI222_X1 us30_U162 (.B2( us30_n747 ) , .B1( us30_n748 ) , .A2( us30_n749 ) , .ZN( us30_n757 ) , .C2( us30_n805 ) , .C1( us30_n814 ) , .A1( us30_n817 ) );
  OAI222_X1 us30_U163 (.ZN( us30_n505 ) , .C2( us30_n625 ) , .B2( us30_n647 ) , .B1( us30_n747 ) , .A2( us30_n748 ) , .C1( us30_n805 ) , .A1( us30_n806 ) );
  OAI222_X1 us30_U164 (.B2( us30_n708 ) , .ZN( us30_n709 ) , .C2( us30_n724 ) , .B1( us30_n747 ) , .A1( us30_n806 ) , .C1( us30_n814 ) , .A2( us30_n815 ) );
  NAND2_X1 us30_U165 (.A1( us30_n447 ) , .A2( us30_n465 ) , .ZN( us30_n749 ) );
  AOI22_X1 us30_U166 (.ZN( us30_n696 ) , .A1( us30_n830 ) , .B2( us30_n843 ) , .A2( us30_n865 ) , .B1( us30_n868 ) );
  AOI22_X1 us30_U167 (.A2( us30_n782 ) , .ZN( us30_n783 ) , .B2( us30_n831 ) , .A1( us30_n834 ) , .B1( us30_n863 ) );
  INV_X1 us30_U168 (.A( us30_n730 ) , .ZN( us30_n839 ) );
  AOI221_X1 us30_U169 (.A( us30_n764 ) , .ZN( us30_n774 ) , .C2( us30_n810 ) , .B2( us30_n835 ) , .C1( us30_n855 ) , .B1( us30_n866 ) );
  OR3_X1 us30_U17 (.ZN( us30_n446 ) , .A1( us30_n528 ) , .A3( us30_n577 ) , .A2( us30_n875 ) );
  AOI21_X1 us30_U170 (.B2( us30_n763 ) , .ZN( us30_n764 ) , .A( us30_n788 ) , .B1( us30_n792 ) );
  INV_X1 us30_U171 (.A( us30_n761 ) , .ZN( us30_n835 ) );
  AOI221_X1 us30_U172 (.A( us30_n483 ) , .ZN( us30_n488 ) , .B1( us30_n831 ) , .C2( us30_n844 ) , .C1( us30_n852 ) , .B2( us30_n862 ) );
  OAI22_X1 us30_U173 (.ZN( us30_n483 ) , .A1( us30_n708 ) , .B2( us30_n785 ) , .A2( us30_n806 ) , .B1( us30_n812 ) );
  INV_X1 us30_U174 (.A( us30_n790 ) , .ZN( us30_n832 ) );
  NAND2_X1 us30_U175 (.A1( us30_n451 ) , .A2( us30_n453 ) , .ZN( us30_n762 ) );
  OAI221_X1 us30_U176 (.A( us30_n727 ) , .C2( us30_n728 ) , .B2( us30_n729 ) , .B1( us30_n730 ) , .ZN( us30_n737 ) , .C1( us30_n817 ) );
  AOI22_X1 us30_U177 (.ZN( us30_n727 ) , .B1( us30_n832 ) , .A2( us30_n838 ) , .A1( us30_n863 ) , .B2( us30_n866 ) );
  INV_X1 us30_U178 (.A( us30_n786 ) , .ZN( us30_n862 ) );
  OAI22_X1 us30_U179 (.ZN( us30_n710 ) , .A2( us30_n728 ) , .B2( us30_n729 ) , .A1( us30_n744 ) , .B1( us30_n813 ) );
  OR4_X1 us30_U18 (.A4( us30_n442 ) , .A2( us30_n443 ) , .A1( us30_n444 ) , .ZN( us30_n445 ) , .A3( us30_n553 ) );
  INV_X1 us30_U180 (.A( us30_n816 ) , .ZN( us30_n831 ) );
  OAI22_X1 us30_U181 (.ZN( us30_n489 ) , .A1( us30_n724 ) , .B2( us30_n728 ) , .B1( us30_n730 ) , .A2( us30_n779 ) );
  OAI22_X1 us30_U182 (.ZN( us30_n624 ) , .B1( us30_n669 ) , .B2( us30_n747 ) , .A1( us30_n815 ) , .A2( us30_n816 ) );
  INV_X1 us30_U183 (.A( us30_n744 ) , .ZN( us30_n837 ) );
  INV_X1 us30_U184 (.A( us30_n788 ) , .ZN( us30_n845 ) );
  OAI22_X1 us30_U185 (.B2( us30_n779 ) , .B1( us30_n780 ) , .ZN( us30_n781 ) , .A2( us30_n814 ) , .A1( us30_n815 ) );
  OAI22_X1 us30_U186 (.A1( us30_n724 ) , .ZN( us30_n726 ) , .B2( us30_n750 ) , .B1( us30_n812 ) , .A2( us30_n816 ) );
  INV_X1 us30_U187 (.A( us30_n805 ) , .ZN( us30_n860 ) );
  INV_X1 us30_U188 (.A( us30_n814 ) , .ZN( us30_n833 ) );
  INV_X1 us30_U189 (.A( us30_n669 ) , .ZN( us30_n865 ) );
  INV_X1 us30_U19 (.A( us30_n613 ) , .ZN( us30_n875 ) );
  OAI22_X1 us30_U190 (.B2( us30_n744 ) , .ZN( us30_n746 ) , .A2( us30_n762 ) , .B1( us30_n780 ) , .A1( us30_n792 ) );
  OAI22_X1 us30_U191 (.ZN( us30_n496 ) , .A2( us30_n744 ) , .A1( us30_n780 ) , .B1( us30_n791 ) , .B2( us30_n806 ) );
  OAI22_X1 us30_U192 (.B2( us30_n803 ) , .B1( us30_n804 ) , .A2( us30_n805 ) , .A1( us30_n806 ) , .ZN( us30_n808 ) );
  AOI211_X1 us30_U193 (.A( us30_n637 ) , .ZN( us30_n645 ) , .B( us30_n743 ) , .C2( us30_n839 ) , .C1( us30_n854 ) );
  OAI22_X1 us30_U194 (.ZN( us30_n637 ) , .A1( us30_n699 ) , .B2( us30_n728 ) , .A2( us30_n762 ) , .B1( us30_n816 ) );
  OAI22_X1 us30_U195 (.B1( us30_n490 ) , .ZN( us30_n491 ) , .A1( us30_n686 ) , .A2( us30_n763 ) , .B2( us30_n817 ) );
  NOR3_X1 us30_U196 (.ZN( us30_n490 ) , .A1( us30_n782 ) , .A2( us30_n850 ) , .A3( us30_n863 ) );
  INV_X1 us30_U197 (.A( us30_n750 ) , .ZN( us30_n842 ) );
  OAI22_X1 us30_U198 (.ZN( us30_n695 ) , .A2( us30_n730 ) , .A1( us30_n780 ) , .B1( us30_n791 ) , .B2( us30_n817 ) );
  NOR2_X1 us30_U199 (.ZN( us30_n715 ) , .A1( us30_n805 ) , .A2( us30_n817 ) );
  INV_X1 us30_U20 (.A( us30_n749 ) , .ZN( us30_n863 ) );
  NOR2_X1 us30_U200 (.ZN( us30_n666 ) , .A1( us30_n728 ) , .A2( us30_n803 ) );
  NOR2_X1 us30_U201 (.ZN( us30_n594 ) , .A2( us30_n697 ) , .A1( us30_n728 ) );
  NOR2_X1 us30_U202 (.ZN( us30_n570 ) , .A1( us30_n728 ) , .A2( us30_n806 ) );
  NOR2_X1 us30_U203 (.A2( us30_n744 ) , .ZN( us30_n755 ) , .A1( us30_n805 ) );
  NOR2_X1 us30_U204 (.ZN( us30_n735 ) , .A2( us30_n803 ) , .A1( us30_n805 ) );
  NOR2_X1 us30_U205 (.ZN( us30_n546 ) , .A2( us30_n780 ) , .A1( us30_n814 ) );
  NOR2_X1 us30_U206 (.ZN( us30_n577 ) , .A2( us30_n699 ) , .A1( us30_n814 ) );
  NOR2_X1 us30_U207 (.ZN( us30_n654 ) , .A1( us30_n728 ) , .A2( us30_n813 ) );
  NOR2_X1 us30_U208 (.ZN( us30_n718 ) , .A2( us30_n724 ) , .A1( us30_n744 ) );
  NOR2_X1 us30_U209 (.ZN( us30_n532 ) , .A2( us30_n749 ) , .A1( us30_n750 ) );
  AOI222_X1 us30_U21 (.ZN( us30_n605 ) , .B2( us30_n671 ) , .B1( us30_n753 ) , .C2( us30_n831 ) , .A1( us30_n833 ) , .A2( us30_n862 ) , .C1( us30_n863 ) );
  NOR2_X1 us30_U210 (.ZN( us30_n615 ) , .A1( us30_n785 ) , .A2( us30_n815 ) );
  NOR2_X1 us30_U211 (.ZN( us30_n629 ) , .A2( us30_n728 ) , .A1( us30_n785 ) );
  NOR2_X1 us30_U212 (.ZN( us30_n611 ) , .A2( us30_n780 ) , .A1( us30_n806 ) );
  NOR2_X1 us30_U213 (.ZN( us30_n628 ) , .A2( us30_n669 ) , .A1( us30_n785 ) );
  INV_X1 us30_U214 (.A( us30_n747 ) , .ZN( us30_n834 ) );
  INV_X1 us30_U215 (.A( us30_n728 ) , .ZN( us30_n852 ) );
  NOR2_X1 us30_U216 (.ZN( us30_n652 ) , .A1( us30_n669 ) , .A2( us30_n814 ) );
  NOR2_X1 us30_U217 (.A1( us30_n669 ) , .ZN( us30_n673 ) , .A2( us30_n744 ) );
  NOR2_X1 us30_U218 (.ZN( us30_n602 ) , .A1( us30_n669 ) , .A2( us30_n803 ) );
  NOR2_X1 us30_U219 (.A1( us30_n669 ) , .ZN( us30_n688 ) , .A2( us30_n816 ) );
  AOI222_X1 us30_U22 (.ZN( us30_n563 ) , .B1( us30_n830 ) , .C1( us30_n841 ) , .A2( us30_n843 ) , .A1( us30_n854 ) , .B2( us30_n863 ) , .C2( us30_n873 ) );
  NOR2_X1 us30_U220 (.A2( us30_n744 ) , .ZN( us30_n769 ) , .A1( us30_n812 ) );
  NOR2_X1 us30_U221 (.ZN( us30_n531 ) , .A2( us30_n780 ) , .A1( us30_n816 ) );
  INV_X1 us30_U222 (.A( us30_n792 ) , .ZN( us30_n851 ) );
  NOR2_X1 us30_U223 (.A2( us30_n708 ) , .A1( us30_n750 ) , .ZN( us30_n771 ) );
  NOR2_X1 us30_U224 (.ZN( us30_n599 ) , .A2( us30_n791 ) , .A1( us30_n816 ) );
  NOR2_X1 us30_U225 (.A1( us30_n669 ) , .ZN( us30_n766 ) , .A2( us30_n813 ) );
  NOR2_X1 us30_U226 (.ZN( us30_n601 ) , .A2( us30_n780 ) , .A1( us30_n803 ) );
  NOR2_X1 us30_U227 (.A1( us30_n699 ) , .ZN( us30_n768 ) , .A2( us30_n813 ) );
  NOR2_X1 us30_U228 (.ZN( us30_n541 ) , .A2( us30_n697 ) , .A1( us30_n699 ) );
  NOR2_X1 us30_U229 (.ZN( us30_n527 ) , .A1( us30_n669 ) , .A2( us30_n779 ) );
  AOI222_X1 us30_U23 (.ZN( us30_n660 ) , .A2( us30_n839 ) , .B1( us30_n841 ) , .C2( us30_n845 ) , .A1( us30_n860 ) , .C1( us30_n863 ) , .B2( us30_n870 ) );
  NOR2_X1 us30_U230 (.ZN( us30_n667 ) , .A1( us30_n750 ) , .A2( us30_n815 ) );
  NOR2_X1 us30_U231 (.ZN( us30_n555 ) , .A1( us30_n750 ) , .A2( us30_n791 ) );
  NOR2_X1 us30_U232 (.ZN( us30_n508 ) , .A2( us30_n780 ) , .A1( us30_n785 ) );
  NOR2_X1 us30_U233 (.ZN( us30_n543 ) , .A2( us30_n708 ) , .A1( us30_n785 ) );
  NOR2_X1 us30_U234 (.ZN( us30_n528 ) , .A2( us30_n724 ) , .A1( us30_n803 ) );
  NOR2_X1 us30_U235 (.ZN( us30_n664 ) , .A1( us30_n785 ) , .A2( us30_n791 ) );
  NOR2_X1 us30_U236 (.ZN( us30_n556 ) , .A1( us30_n762 ) , .A2( us30_n805 ) );
  INV_X1 us30_U237 (.A( us30_n806 ) , .ZN( us30_n841 ) );
  NOR2_X1 us30_U238 (.ZN( us30_n661 ) , .A1( us30_n729 ) , .A2( us30_n790 ) );
  OAI22_X1 us30_U239 (.B1( us30_n440 ) , .ZN( us30_n444 ) , .A2( us30_n728 ) , .A1( us30_n744 ) , .B2( us30_n749 ) );
  INV_X1 us30_U24 (.A( us30_n647 ) , .ZN( us30_n870 ) );
  NOR3_X1 us30_U240 (.ZN( us30_n440 ) , .A2( us30_n836 ) , .A3( us30_n837 ) , .A1( us30_n846 ) );
  NOR2_X1 us30_U241 (.ZN( us30_n507 ) , .A1( us30_n812 ) , .A2( us30_n817 ) );
  NOR2_X1 us30_U242 (.ZN( us30_n557 ) , .A1( us30_n792 ) , .A2( us30_n814 ) );
  NOR2_X1 us30_U243 (.ZN( us30_n545 ) , .A1( us30_n749 ) , .A2( us30_n814 ) );
  NOR2_X1 us30_U244 (.ZN( us30_n509 ) , .A1( us30_n729 ) , .A2( us30_n779 ) );
  NOR2_X1 us30_U245 (.ZN( us30_n662 ) , .A2( us30_n697 ) , .A1( us30_n729 ) );
  OAI22_X1 us30_U246 (.B2( us30_n750 ) , .B1( us30_n751 ) , .A1( us30_n752 ) , .ZN( us30_n756 ) , .A2( us30_n806 ) );
  NOR2_X1 us30_U247 (.ZN( us30_n751 ) , .A2( us30_n852 ) , .A1( us30_n860 ) );
  NOR3_X1 us30_U248 (.ZN( us30_n752 ) , .A2( us30_n853 ) , .A1( us30_n863 ) , .A3( us30_n865 ) );
  NOR2_X1 us30_U249 (.ZN( us30_n544 ) , .A2( us30_n785 ) , .A1( us30_n792 ) );
  NOR4_X1 us30_U25 (.ZN( us30_n473 ) , .A2( us30_n521 ) , .A4( us30_n594 ) , .A1( us30_n609 ) , .A3( us30_n629 ) );
  NOR2_X1 us30_U250 (.ZN( us30_n663 ) , .A1( us30_n729 ) , .A2( us30_n785 ) );
  NOR2_X1 us30_U251 (.ZN( us30_n530 ) , .A2( us30_n744 ) , .A1( us30_n792 ) );
  NOR2_X1 us30_U252 (.ZN( us30_n506 ) , .A2( us30_n728 ) , .A1( us30_n762 ) );
  NOR2_X1 us30_U253 (.ZN( us30_n631 ) , .A1( us30_n724 ) , .A2( us30_n813 ) );
  NOR2_X1 us30_U254 (.ZN( us30_n614 ) , .A1( us30_n762 ) , .A2( us30_n812 ) );
  NOR2_X1 us30_U255 (.A1( us30_n749 ) , .ZN( us30_n767 ) , .A2( us30_n803 ) );
  NOR2_X1 us30_U256 (.ZN( us30_n516 ) , .A1( us30_n708 ) , .A2( us30_n744 ) );
  NOR2_X1 us30_U257 (.ZN( us30_n670 ) , .A1( us30_n790 ) , .A2( us30_n805 ) );
  NOR2_X1 us30_U258 (.ZN( us30_n558 ) , .A1( us30_n708 ) , .A2( us30_n816 ) );
  NOR2_X1 us30_U259 (.A2( us30_n697 ) , .ZN( us30_n716 ) , .A1( us30_n792 ) );
  NOR4_X1 us30_U26 (.ZN( us30_n479 ) , .A1( us30_n520 ) , .A4( us30_n557 ) , .A3( us30_n582 ) , .A2( us30_n630 ) );
  NOR2_X1 us30_U260 (.ZN( us30_n517 ) , .A1( us30_n708 ) , .A2( us30_n803 ) );
  NOR2_X1 us30_U261 (.ZN( us30_n521 ) , .A1( us30_n790 ) , .A2( us30_n812 ) );
  NOR2_X1 us30_U262 (.ZN( us30_n630 ) , .A1( us30_n747 ) , .A2( us30_n815 ) );
  NOR2_X1 us30_U263 (.ZN( us30_n655 ) , .A1( us30_n790 ) , .A2( us30_n815 ) );
  INV_X1 us30_U264 (.A( us30_n763 ) , .ZN( us30_n866 ) );
  AOI21_X1 us30_U265 (.ZN( us30_n552 ) , .B1( us30_n669 ) , .A( us30_n697 ) , .B2( us30_n805 ) );
  NOR2_X1 us30_U266 (.ZN( us30_n668 ) , .A2( us30_n708 ) , .A1( us30_n790 ) );
  NOR2_X1 us30_U267 (.ZN( us30_n542 ) , .A1( us30_n762 ) , .A2( us30_n791 ) );
  NOR2_X1 us30_U268 (.ZN( us30_n656 ) , .A1( us30_n747 ) , .A2( us30_n780 ) );
  NOR2_X1 us30_U269 (.ZN( us30_n609 ) , .A2( us30_n724 ) , .A1( us30_n817 ) );
  NOR4_X1 us30_U27 (.A4( us30_n532 ) , .A3( us30_n533 ) , .A2( us30_n534 ) , .ZN( us30_n535 ) , .A1( us30_n820 ) );
  INV_X1 us30_U270 (.A( us30_n729 ) , .ZN( us30_n868 ) );
  AOI21_X1 us30_U271 (.B1( us30_n625 ) , .ZN( us30_n627 ) , .A( us30_n763 ) , .B2( us30_n814 ) );
  AOI21_X1 us30_U272 (.ZN( us30_n650 ) , .A( us30_n779 ) , .B1( us30_n792 ) , .B2( us30_n805 ) );
  AOI21_X1 us30_U273 (.A( us30_n815 ) , .B2( us30_n816 ) , .B1( us30_n817 ) , .ZN( us30_n818 ) );
  NOR2_X1 us30_U274 (.ZN( us30_n579 ) , .A2( us30_n708 ) , .A1( us30_n730 ) );
  NOR2_X1 us30_U275 (.ZN( us30_n533 ) , .A2( us30_n724 ) , .A1( us30_n730 ) );
  NOR2_X1 us30_U276 (.ZN( us30_n642 ) , .A2( us30_n788 ) , .A1( us30_n791 ) );
  AOI21_X1 us30_U277 (.A( us30_n812 ) , .B2( us30_n813 ) , .B1( us30_n814 ) , .ZN( us30_n819 ) );
  NOR2_X1 us30_U278 (.A2( us30_n708 ) , .A1( us30_n762 ) , .ZN( us30_n794 ) );
  NOR2_X1 us30_U279 (.A2( us30_n697 ) , .A1( us30_n780 ) , .ZN( us30_n820 ) );
  NOR4_X1 us30_U28 (.ZN( us30_n456 ) , .A2( us30_n517 ) , .A1( us30_n543 ) , .A3( us30_n579 ) , .A4( us30_n615 ) );
  AOI21_X1 us30_U280 (.ZN( us30_n626 ) , .B2( us30_n669 ) , .A( us30_n790 ) , .B1( us30_n791 ) );
  AOI21_X1 us30_U281 (.ZN( us30_n499 ) , .B1( us30_n680 ) , .A( us30_n812 ) , .B2( us30_n816 ) );
  NOR2_X1 us30_U282 (.ZN( us30_n520 ) , .A2( us30_n708 ) , .A1( us30_n814 ) );
  AOI21_X1 us30_U283 (.ZN( us30_n477 ) , .A( us30_n669 ) , .B1( us30_n750 ) , .B2( us30_n806 ) );
  NOR2_X1 us30_U284 (.ZN( us30_n582 ) , .A1( us30_n744 ) , .A2( us30_n815 ) );
  AOI21_X1 us30_U285 (.ZN( us30_n593 ) , .B1( us30_n750 ) , .A( us30_n792 ) , .B2( us30_n813 ) );
  AOI21_X1 us30_U286 (.ZN( us30_n515 ) , .A( us30_n729 ) , .B1( us30_n750 ) , .B2( us30_n803 ) );
  NOR2_X1 us30_U287 (.A1( us30_n697 ) , .ZN( us30_n770 ) , .A2( us30_n815 ) );
  AOI21_X1 us30_U288 (.ZN( us30_n510 ) , .B2( us30_n669 ) , .A( us30_n730 ) , .B1( us30_n815 ) );
  NOR2_X1 us30_U289 (.ZN( us30_n519 ) , .A2( us30_n699 ) , .A1( us30_n816 ) );
  NOR4_X1 us30_U29 (.A4( us30_n541 ) , .A3( us30_n542 ) , .A2( us30_n543 ) , .ZN( us30_n550 ) , .A1( us30_n688 ) );
  NOR2_X1 us30_U290 (.ZN( us30_n559 ) , .A2( us30_n791 ) , .A1( us30_n803 ) );
  NOR2_X1 us30_U291 (.ZN( us30_n581 ) , .A1( us30_n669 ) , .A2( us30_n788 ) );
  INV_X1 us30_U292 (.A( us30_n813 ) , .ZN( us30_n836 ) );
  NOR2_X1 us30_U293 (.ZN( us30_n683 ) , .A2( us30_n699 ) , .A1( us30_n803 ) );
  AOI21_X1 us30_U294 (.ZN( us30_n589 ) , .B2( us30_n699 ) , .B1( us30_n815 ) , .A( us30_n817 ) );
  AOI21_X1 us30_U295 (.ZN( us30_n539 ) , .B2( us30_n812 ) , .A( us30_n814 ) , .B1( us30_n815 ) );
  AOI21_X1 us30_U296 (.ZN( us30_n540 ) , .A( us30_n763 ) , .B2( us30_n779 ) , .B1( us30_n817 ) );
  AOI21_X1 us30_U297 (.B1( us30_n699 ) , .ZN( us30_n700 ) , .A( us30_n732 ) , .B2( us30_n763 ) );
  AOI21_X1 us30_U298 (.ZN( us30_n591 ) , .B2( us30_n763 ) , .A( us30_n785 ) , .B1( us30_n812 ) );
  AOI21_X1 us30_U299 (.ZN( us30_n498 ) , .A( us30_n724 ) , .B2( us30_n762 ) , .B1( us30_n814 ) );
  NAND2_X1 us30_U3 (.A2( us30_n448 ) , .A1( us30_n464 ) , .ZN( us30_n815 ) );
  AOI221_X1 us30_U30 (.A( us30_n713 ) , .B2( us30_n714 ) , .ZN( us30_n720 ) , .C1( us30_n832 ) , .B1( us30_n839 ) , .C2( us30_n863 ) );
  NOR2_X1 us30_U300 (.ZN( us30_n547 ) , .A1( us30_n699 ) , .A2( us30_n744 ) );
  INV_X1 us30_U301 (.A( us30_n791 ) , .ZN( us30_n873 ) );
  AOI21_X1 us30_U302 (.ZN( us30_n649 ) , .B1( us30_n729 ) , .B2( us30_n763 ) , .A( us30_n813 ) );
  NOR2_X1 us30_U303 (.ZN( us30_n685 ) , .A1( us30_n729 ) , .A2( us30_n816 ) );
  AOI21_X1 us30_U304 (.B1( us30_n686 ) , .ZN( us30_n687 ) , .A( us30_n728 ) , .B2( us30_n761 ) );
  AOI21_X1 us30_U305 (.ZN( us30_n569 ) , .B1( us30_n750 ) , .B2( us30_n762 ) , .A( us30_n780 ) );
  AOI21_X1 us30_U306 (.ZN( us30_n571 ) , .B2( us30_n697 ) , .B1( us30_n806 ) , .A( us30_n812 ) );
  NOR2_X1 us30_U307 (.ZN( us30_n568 ) , .A1( us30_n729 ) , .A2( us30_n762 ) );
  NOR2_X1 us30_U308 (.ZN( us30_n566 ) , .A2( us30_n697 ) , .A1( us30_n763 ) );
  AOI21_X1 us30_U309 (.ZN( us30_n640 ) , .B2( us30_n747 ) , .A( us30_n792 ) , .B1( us30_n803 ) );
  OR2_X1 us30_U31 (.A2( us30_n711 ) , .A1( us30_n712 ) , .ZN( us30_n713 ) );
  INV_X1 us30_U310 (.A( us30_n699 ) , .ZN( us30_n853 ) );
  AOI21_X1 us30_U311 (.ZN( us30_n514 ) , .A( us30_n779 ) , .B2( us30_n792 ) , .B1( us30_n812 ) );
  AOI21_X1 us30_U312 (.ZN( us30_n639 ) , .B2( us30_n749 ) , .A( us30_n788 ) , .B1( us30_n812 ) );
  NAND2_X1 us30_U313 (.ZN( us30_n753 ) , .A1( us30_n763 ) , .A2( us30_n805 ) );
  NOR2_X1 us30_U314 (.ZN( us30_n665 ) , .A1( us30_n780 ) , .A2( us30_n813 ) );
  AOI21_X1 us30_U315 (.ZN( us30_n564 ) , .B1( us30_n724 ) , .A( us30_n779 ) , .B2( us30_n791 ) );
  AOI21_X1 us30_U316 (.ZN( us30_n497 ) , .A( us30_n779 ) , .B2( us30_n791 ) , .B1( us30_n804 ) );
  AOI21_X1 us30_U317 (.ZN( us30_n689 ) , .B2( us30_n749 ) , .B1( us30_n763 ) , .A( us30_n806 ) );
  AOI21_X1 us30_U318 (.ZN( us30_n450 ) , .B2( us30_n792 ) , .A( us30_n803 ) , .B1( us30_n815 ) );
  NOR2_X1 us30_U319 (.ZN( us30_n567 ) , .A1( us30_n747 ) , .A2( us30_n805 ) );
  NOR2_X1 us30_U32 (.ZN( us30_n680 ) , .A2( us30_n834 ) , .A1( us30_n839 ) );
  NOR2_X1 us30_U320 (.ZN( us30_n529 ) , .A1( us30_n708 ) , .A2( us30_n779 ) );
  NOR2_X1 us30_U321 (.ZN( us30_n578 ) , .A1( us30_n708 ) , .A2( us30_n813 ) );
  AOI21_X1 us30_U322 (.ZN( us30_n478 ) , .B2( us30_n697 ) , .A( us30_n749 ) , .B1( us30_n779 ) );
  AOI21_X1 us30_U323 (.A( us30_n790 ) , .B2( us30_n791 ) , .B1( us30_n792 ) , .ZN( us30_n793 ) );
  NOR2_X1 us30_U324 (.ZN( us30_n684 ) , .A1( us30_n791 ) , .A2( us30_n813 ) );
  AOI21_X1 us30_U325 (.A( us30_n733 ) , .ZN( us30_n734 ) , .B2( us30_n780 ) , .B1( us30_n792 ) );
  NOR2_X1 us30_U326 (.A2( us30_n813 ) , .A1( us30_n815 ) , .ZN( us30_n821 ) );
  AOI21_X1 us30_U327 (.ZN( us30_n641 ) , .B1( us30_n680 ) , .A( us30_n791 ) , .B2( us30_n817 ) );
  NOR2_X1 us30_U328 (.ZN( us30_n711 ) , .A1( us30_n762 ) , .A2( us30_n763 ) );
  NOR2_X1 us30_U329 (.ZN( us30_n583 ) , .A1( us30_n792 ) , .A2( us30_n817 ) );
  AOI222_X1 us30_U33 (.ZN( us30_n469 ) , .B1( us30_n832 ) , .A1( us30_n839 ) , .C1( us30_n842 ) , .C2( us30_n851 ) , .A2( us30_n855 ) , .B2( us30_n865 ) );
  NOR2_X1 us30_U330 (.ZN( us30_n534 ) , .A1( us30_n724 ) , .A2( us30_n788 ) );
  NOR2_X1 us30_U331 (.ZN( us30_n632 ) , .A2( us30_n697 ) , .A1( us30_n724 ) );
  NOR2_X1 us30_U332 (.ZN( us30_n682 ) , .A2( us30_n708 ) , .A1( us30_n817 ) );
  NOR2_X1 us30_U333 (.ZN( us30_n580 ) , .A2( us30_n697 ) , .A1( us30_n791 ) );
  INV_X1 us30_U334 (.A( us30_n815 ) , .ZN( us30_n855 ) );
  AOI21_X1 us30_U335 (.ZN( us30_n442 ) , .A( us30_n699 ) , .B1( us30_n733 ) , .B2( us30_n750 ) );
  INV_X1 us30_U336 (.A( us30_n780 ) , .ZN( us30_n850 ) );
  INV_X1 us30_U337 (.A( us30_n785 ) , .ZN( us30_n846 ) );
  NAND2_X1 us30_U338 (.ZN( us30_n714 ) , .A1( us30_n728 ) , .A2( us30_n780 ) );
  NAND2_X1 us30_U339 (.A2( us30_n762 ) , .A1( us30_n806 ) , .ZN( us30_n810 ) );
  NOR4_X1 us30_U34 (.A1( us30_n466 ) , .ZN( us30_n467 ) , .A4( us30_n542 ) , .A2( us30_n554 ) , .A3( us30_n614 ) );
  AOI21_X1 us30_U340 (.ZN( us30_n443 ) , .B1( us30_n789 ) , .B2( us30_n791 ) , .A( us30_n814 ) );
  NAND2_X1 us30_U341 (.ZN( us30_n671 ) , .A1( us30_n806 ) , .A2( us30_n816 ) );
  NOR2_X1 us30_U342 (.ZN( us30_n484 ) , .A1( us30_n788 ) , .A2( us30_n805 ) );
  NOR2_X1 us30_U343 (.ZN( us30_n470 ) , .A2( us30_n779 ) , .A1( us30_n815 ) );
  NOR2_X1 us30_U344 (.ZN( us30_n712 ) , .A2( us30_n724 ) , .A1( us30_n790 ) );
  OAI21_X1 us30_U345 (.A( us30_n787 ) , .B2( us30_n788 ) , .B1( us30_n789 ) , .ZN( us30_n795 ) );
  OAI21_X1 us30_U346 (.ZN( us30_n787 ) , .A( us30_n839 ) , .B1( us30_n863 ) , .B2( us30_n873 ) );
  NOR2_X1 us30_U347 (.ZN( us30_n526 ) , .A1( us30_n724 ) , .A2( us30_n750 ) );
  NAND2_X1 us30_U348 (.A1( us30_n699 ) , .A2( us30_n729 ) , .ZN( us30_n782 ) );
  NOR2_X1 us30_U349 (.ZN( us30_n518 ) , .A1( us30_n708 ) , .A2( us30_n788 ) );
  AOI221_X1 us30_U35 (.ZN( us30_n468 ) , .C2( us30_n714 ) , .B2( us30_n831 ) , .C1( us30_n845 ) , .B1( us30_n860 ) , .A( us30_n864 ) );
  OAI21_X1 us30_U350 (.A( us30_n698 ) , .ZN( us30_n702 ) , .B2( us30_n750 ) , .B1( us30_n804 ) );
  OAI21_X1 us30_U351 (.ZN( us30_n698 ) , .B2( us30_n833 ) , .B1( us30_n838 ) , .A( us30_n860 ) );
  OAI21_X1 us30_U352 (.A( us30_n731 ) , .B1( us30_n732 ) , .ZN( us30_n736 ) , .B2( us30_n805 ) );
  OAI21_X1 us30_U353 (.ZN( us30_n731 ) , .A( us30_n833 ) , .B2( us30_n852 ) , .B1( us30_n873 ) );
  INV_X1 us30_U354 (.A( us30_n817 ) , .ZN( us30_n844 ) );
  INV_X1 us30_U355 (.A( us30_n724 ) , .ZN( us30_n856 ) );
  AND2_X1 us30_U356 (.ZN( us30_n732 ) , .A1( us30_n779 ) , .A2( us30_n785 ) );
  NAND2_X1 us30_U357 (.A1( us30_n447 ) , .A2( us30_n449 ) , .ZN( us30_n805 ) );
  NAND2_X1 us30_U358 (.A1( us30_n451 ) , .A2( us30_n454 ) , .ZN( us30_n814 ) );
  NAND2_X1 us30_U359 (.A1( us30_n452 ) , .A2( us30_n465 ) , .ZN( us30_n669 ) );
  NOR4_X1 us30_U36 (.A4( us30_n514 ) , .A3( us30_n515 ) , .A2( us30_n516 ) , .A1( us30_n517 ) , .ZN( us30_n524 ) );
  NAND2_X1 us30_U360 (.A2( us30_n448 ) , .A1( us30_n460 ) , .ZN( us30_n728 ) );
  NAND2_X1 us30_U361 (.A1( us30_n455 ) , .A2( us30_n462 ) , .ZN( us30_n750 ) );
  NAND2_X1 us30_U362 (.A2( us30_n453 ) , .A1( us30_n455 ) , .ZN( us30_n806 ) );
  NAND2_X1 us30_U363 (.A1( us30_n451 ) , .A2( us30_n471 ) , .ZN( us30_n816 ) );
  NAND2_X1 us30_U364 (.A1( us30_n454 ) , .A2( us30_n461 ) , .ZN( us30_n813 ) );
  NAND2_X1 us30_U365 (.A1( us30_n455 ) , .A2( us30_n471 ) , .ZN( us30_n803 ) );
  NAND2_X1 us30_U366 (.A1( us30_n453 ) , .A2( us30_n461 ) , .ZN( us30_n744 ) );
  NAND2_X1 us30_U367 (.A1( us30_n453 ) , .A2( us30_n472 ) , .ZN( us30_n785 ) );
  NAND2_X1 us30_U368 (.A2( us30_n454 ) , .A1( us30_n472 ) , .ZN( us30_n779 ) );
  NAND2_X1 us30_U369 (.A2( us30_n464 ) , .A1( us30_n465 ) , .ZN( us30_n812 ) );
  AOI222_X1 us30_U37 (.ZN( us30_n525 ) , .A1( us30_n834 ) , .B2( us30_n837 ) , .C1( us30_n844 ) , .C2( us30_n850 ) , .A2( us30_n852 ) , .B1( us30_n866 ) );
  NAND2_X1 us30_U370 (.A1( us30_n441 ) , .A2( us30_n460 ) , .ZN( us30_n699 ) );
  NAND2_X1 us30_U371 (.A2( us30_n449 ) , .A1( us30_n452 ) , .ZN( us30_n763 ) );
  NAND2_X1 us30_U372 (.A2( us30_n448 ) , .A1( us30_n452 ) , .ZN( us30_n729 ) );
  NAND2_X1 us30_U373 (.A2( us30_n461 ) , .A1( us30_n462 ) , .ZN( us30_n747 ) );
  NAND2_X1 us30_U374 (.A1( us30_n462 ) , .A2( us30_n472 ) , .ZN( us30_n788 ) );
  NOR2_X1 us30_U375 (.ZN( us30_n465 ) , .A2( us30_n847 ) , .A1( us30_n848 ) );
  NOR2_X1 us30_U376 (.ZN( us30_n453 ) , .A1( us30_n826 ) , .A2( us30_n827 ) );
  NOR2_X1 us30_U377 (.ZN( us30_n451 ) , .A1( us30_n828 ) , .A2( us30_n829 ) );
  NAND2_X1 us30_U378 (.A1( us30_n451 ) , .A2( us30_n462 ) , .ZN( us30_n790 ) );
  NAND2_X1 us30_U379 (.A2( us30_n441 ) , .A1( us30_n447 ) , .ZN( us30_n784 ) );
  NOR4_X1 us30_U38 (.A3( us30_n521 ) , .A1( us30_n522 ) , .ZN( us30_n523 ) , .A2( us30_n673 ) , .A4( us30_n769 ) );
  NAND2_X1 us30_U380 (.A2( us30_n454 ) , .A1( us30_n455 ) , .ZN( us30_n730 ) );
  NAND2_X2 us30_U381 (.A1( us30_n449 ) , .A2( us30_n464 ) , .ZN( us30_n724 ) );
  NAND2_X2 us30_U382 (.A1( us30_n449 ) , .A2( us30_n460 ) , .ZN( us30_n792 ) );
  NAND2_X2 us30_U383 (.A2( us30_n460 ) , .A1( us30_n465 ) , .ZN( us30_n780 ) );
  NOR2_X1 us30_U384 (.ZN( us30_n447 ) , .A2( us30_n849 ) , .A1( us30_n858 ) );
  NAND2_X1 us30_U385 (.A1( us30_n447 ) , .A2( us30_n448 ) , .ZN( us30_n786 ) );
  NOR2_X1 us30_U386 (.A2( sa30_6 ) , .A1( sa30_7 ) , .ZN( us30_n464 ) );
  NOR2_X1 us30_U387 (.A2( sa30_7 ) , .ZN( us30_n460 ) , .A1( us30_n849 ) );
  NOR2_X1 us30_U388 (.A2( sa30_4 ) , .ZN( us30_n449 ) , .A1( us30_n848 ) );
  NOR2_X1 us30_U389 (.A2( sa30_4 ) , .A1( sa30_5 ) , .ZN( us30_n441 ) );
  AOI221_X1 us30_U39 (.A( us30_n781 ) , .ZN( us30_n798 ) , .C2( us30_n837 ) , .B2( us30_n838 ) , .B1( us30_n865 ) , .C1( us30_n866 ) );
  NOR2_X1 us30_U390 (.A2( sa30_5 ) , .ZN( us30_n448 ) , .A1( us30_n847 ) );
  NOR2_X1 us30_U391 (.A2( sa30_2 ) , .A1( sa30_3 ) , .ZN( us30_n472 ) );
  NOR2_X1 us30_U392 (.A2( sa30_6 ) , .ZN( us30_n452 ) , .A1( us30_n858 ) );
  NOR2_X1 us30_U393 (.A2( sa30_1 ) , .ZN( us30_n471 ) , .A1( us30_n826 ) );
  NOR2_X1 us30_U394 (.A2( sa30_0 ) , .ZN( us30_n454 ) , .A1( us30_n827 ) );
  NOR2_X1 us30_U395 (.A2( sa30_0 ) , .A1( sa30_1 ) , .ZN( us30_n462 ) );
  NOR2_X1 us30_U396 (.A2( sa30_3 ) , .ZN( us30_n455 ) , .A1( us30_n828 ) );
  NOR2_X1 us30_U397 (.A2( sa30_2 ) , .ZN( us30_n461 ) , .A1( us30_n829 ) );
  INV_X1 us30_U398 (.A( sa30_6 ) , .ZN( us30_n849 ) );
  INV_X1 us30_U399 (.A( sa30_4 ) , .ZN( us30_n847 ) );
  NAND2_X1 us30_U4 (.A1( us30_n441 ) , .A2( us30_n464 ) , .ZN( us30_n708 ) );
  NOR4_X1 us30_U40 (.A4( us30_n793 ) , .A3( us30_n794 ) , .A2( us30_n795 ) , .A1( us30_n796 ) , .ZN( us30_n797 ) );
  INV_X1 us30_U400 (.A( sa30_3 ) , .ZN( us30_n829 ) );
  INV_X1 us30_U401 (.A( sa30_1 ) , .ZN( us30_n827 ) );
  INV_X1 us30_U402 (.A( sa30_0 ) , .ZN( us30_n826 ) );
  INV_X1 us30_U403 (.A( sa30_2 ) , .ZN( us30_n828 ) );
  INV_X1 us30_U404 (.A( sa30_7 ) , .ZN( us30_n858 ) );
  INV_X1 us30_U405 (.A( sa30_5 ) , .ZN( us30_n848 ) );
  NAND2_X1 us30_U406 (.A2( us30_n461 ) , .A1( us30_n471 ) , .ZN( us30_n697 ) );
  OAI221_X1 us30_U407 (.A( us30_n783 ) , .C2( us30_n784 ) , .B2( us30_n785 ) , .B1( us30_n786 ) , .ZN( us30_n796 ) , .C1( us30_n813 ) );
  NAND2_X1 us30_U408 (.A1( us30_n729 ) , .A2( us30_n784 ) , .ZN( us30_n811 ) );
  OAI22_X1 us30_U409 (.ZN( us30_n588 ) , .A2( us30_n747 ) , .B2( us30_n762 ) , .A1( us30_n763 ) , .B1( us30_n784 ) );
  NOR4_X1 us30_U41 (.A4( us30_n776 ) , .A3( us30_n777 ) , .A1( us30_n778 ) , .ZN( us30_n799 ) , .A2( us30_n801 ) );
  AOI21_X1 us30_U410 (.ZN( us30_n592 ) , .B1( us30_n728 ) , .B2( us30_n784 ) , .A( us30_n790 ) );
  AOI21_X1 us30_U411 (.ZN( us30_n623 ) , .B1( us30_n699 ) , .A( us30_n779 ) , .B2( us30_n784 ) );
  AOI21_X1 us30_U412 (.ZN( us30_n648 ) , .A( us30_n762 ) , .B2( us30_n784 ) , .B1( us30_n792 ) );
  OAI22_X1 us30_U413 (.ZN( us30_n681 ) , .A1( us30_n699 ) , .A2( us30_n730 ) , .B2( us30_n784 ) , .B1( us30_n817 ) );
  OAI21_X1 us30_U414 (.A( us30_n613 ) , .ZN( us30_n616 ) , .B1( us30_n625 ) , .B2( us30_n784 ) );
  NOR2_X1 us30_U415 (.ZN( us30_n610 ) , .A1( us30_n784 ) , .A2( us30_n816 ) );
  OAI222_X1 us30_U416 (.A2( us30_n669 ) , .ZN( us30_n674 ) , .B1( us30_n747 ) , .B2( us30_n784 ) , .C2( us30_n788 ) , .C1( us30_n815 ) , .A1( us30_n817 ) );
  NOR2_X1 us30_U417 (.ZN( us30_n651 ) , .A1( us30_n784 ) , .A2( us30_n788 ) );
  NOR2_X1 us30_U418 (.ZN( us30_n600 ) , .A2( us30_n697 ) , .A1( us30_n784 ) );
  NOR2_X1 us30_U419 (.ZN( us30_n553 ) , .A2( us30_n744 ) , .A1( us30_n784 ) );
  NOR4_X1 us30_U42 (.A3( us30_n755 ) , .A2( us30_n756 ) , .A1( us30_n757 ) , .ZN( us30_n758 ) , .A4( us30_n869 ) );
  INV_X1 us30_U420 (.A( us30_n784 ) , .ZN( us30_n861 ) );
  AOI21_X1 us30_U421 (.ZN( us30_n500 ) , .A( us30_n697 ) , .B1( us30_n708 ) , .B2( us30_n786 ) );
  OAI221_X1 us30_U422 (.A( us30_n696 ) , .ZN( us30_n703 ) , .C2( us30_n784 ) , .C1( us30_n785 ) , .B1( us30_n786 ) , .B2( us30_n806 ) );
  OAI22_X1 us30_U423 (.ZN( us30_n590 ) , .B1( us30_n730 ) , .B2( us30_n749 ) , .A2( us30_n786 ) , .A1( us30_n803 ) );
  NOR2_X1 us30_U424 (.ZN( us30_n612 ) , .A1( us30_n779 ) , .A2( us30_n786 ) );
  NAND2_X1 us30_U425 (.A2( us30_n749 ) , .A1( us30_n786 ) , .ZN( us30_n809 ) );
  OAI222_X1 us30_U426 (.ZN( us30_n617 ) , .B1( us30_n697 ) , .C1( us30_n724 ) , .C2( us30_n747 ) , .B2( us30_n786 ) , .A2( us30_n792 ) , .A1( us30_n816 ) );
  NOR2_X1 us30_U427 (.ZN( us30_n717 ) , .A2( us30_n744 ) , .A1( us30_n786 ) );
  NOR2_X1 us30_U428 (.ZN( us30_n653 ) , .A1( us30_n762 ) , .A2( us30_n786 ) );
  NOR2_X1 us30_U429 (.ZN( us30_n554 ) , .A1( us30_n786 ) , .A2( us30_n813 ) );
  AOI211_X1 us30_U43 (.B( us30_n745 ) , .A( us30_n746 ) , .ZN( us30_n759 ) , .C1( us30_n832 ) , .C2( us30_n853 ) );
  NOR2_X1 us30_U430 (.ZN( us30_n701 ) , .A2( us30_n786 ) , .A1( us30_n817 ) );
  NOR2_X1 us30_U431 (.A1( us30_n730 ) , .ZN( us30_n765 ) , .A2( us30_n786 ) );
  AND2_X1 us30_U432 (.ZN( us30_n438 ) , .A2( us30_n831 ) , .A1( us30_n854 ) );
  AND2_X1 us30_U433 (.ZN( us30_n439 ) , .A2( us30_n843 ) , .A1( us30_n861 ) );
  NOR3_X1 us30_U434 (.A1( us30_n438 ) , .A2( us30_n439 ) , .A3( us30_n576 ) , .ZN( us30_n587 ) );
  NAND4_X1 us30_U435 (.ZN( sa31_sr_2 ) , .A4( us30_n643 ) , .A3( us30_n644 ) , .A2( us30_n645 ) , .A1( us30_n646 ) );
  INV_X1 us30_U436 (.A( us30_n812 ) , .ZN( us30_n854 ) );
  NAND3_X1 us30_U437 (.ZN( sa31_sr_6 ) , .A3( us30_n797 ) , .A2( us30_n798 ) , .A1( us30_n799 ) );
  NAND3_X1 us30_U438 (.ZN( sa31_sr_5 ) , .A3( us30_n758 ) , .A2( us30_n759 ) , .A1( us30_n760 ) );
  NAND3_X1 us30_U439 (.ZN( sa31_sr_4 ) , .A3( us30_n738 ) , .A2( us30_n739 ) , .A1( us30_n740 ) );
  NOR3_X1 us30_U44 (.A3( us30_n741 ) , .A2( us30_n742 ) , .A1( us30_n743 ) , .ZN( us30_n760 ) );
  NAND3_X1 us30_U440 (.A3( us30_n675 ) , .A2( us30_n676 ) , .A1( us30_n677 ) , .ZN( us30_n807 ) );
  NAND3_X1 us30_U441 (.ZN( us30_n638 ) , .A3( us30_n708 ) , .A2( us30_n724 ) , .A1( us30_n792 ) );
  NAND3_X1 us30_U442 (.A3( us30_n618 ) , .A2( us30_n619 ) , .A1( us30_n620 ) , .ZN( us30_n725 ) );
  NAND3_X1 us30_U443 (.A3( us30_n585 ) , .A2( us30_n586 ) , .A1( us30_n587 ) , .ZN( us30_n621 ) );
  NAND3_X1 us30_U444 (.ZN( us30_n565 ) , .A3( us30_n680 ) , .A2( us30_n750 ) , .A1( us30_n785 ) );
  NAND3_X1 us30_U445 (.A3( us30_n523 ) , .A2( us30_n524 ) , .A1( us30_n525 ) , .ZN( us30_n742 ) );
  NAND3_X1 us30_U446 (.A3( us30_n512 ) , .A1( us30_n513 ) , .ZN( us30_n608 ) , .A2( us30_n871 ) );
  NAND3_X1 us30_U447 (.A3( us30_n467 ) , .A2( us30_n468 ) , .A1( us30_n469 ) , .ZN( us30_n777 ) );
  INV_X1 us30_U448 (.A( us30_n803 ) , .ZN( us30_n843 ) );
  AOI21_X1 us30_U449 (.ZN( us30_n576 ) , .B2( us30_n724 ) , .B1( us30_n748 ) , .A( us30_n785 ) );
  NAND4_X1 us30_U45 (.ZN( sa31_sr_3 ) , .A4( us30_n704 ) , .A3( us30_n705 ) , .A2( us30_n706 ) , .A1( us30_n707 ) );
  NOR4_X1 us30_U46 (.A4( us30_n700 ) , .A3( us30_n701 ) , .A2( us30_n702 ) , .A1( us30_n703 ) , .ZN( us30_n704 ) );
  AOI211_X1 us30_U47 (.B( us30_n694 ) , .A( us30_n695 ) , .ZN( us30_n705 ) , .C2( us30_n831 ) , .C1( us30_n851 ) );
  NOR2_X1 us30_U48 (.ZN( us30_n707 ) , .A2( us30_n776 ) , .A1( us30_n800 ) );
  AOI222_X1 us30_U49 (.B2( us30_n638 ) , .ZN( us30_n644 ) , .B1( us30_n841 ) , .A1( us30_n842 ) , .C2( us30_n846 ) , .C1( us30_n863 ) , .A2( us30_n865 ) );
  NAND2_X1 us30_U5 (.A2( us30_n441 ) , .A1( us30_n452 ) , .ZN( us30_n791 ) );
  NOR4_X1 us30_U50 (.A4( us30_n639 ) , .A3( us30_n640 ) , .A2( us30_n641 ) , .A1( us30_n642 ) , .ZN( us30_n643 ) );
  NOR3_X1 us30_U51 (.A2( us30_n607 ) , .A1( us30_n608 ) , .ZN( us30_n646 ) , .A3( us30_n722 ) );
  NOR2_X1 us30_U52 (.ZN( us30_n804 ) , .A1( us30_n854 ) , .A2( us30_n861 ) );
  NAND4_X1 us30_U53 (.ZN( sa31_sr_7 ) , .A4( us30_n822 ) , .A3( us30_n823 ) , .A2( us30_n824 ) , .A1( us30_n825 ) );
  NOR4_X1 us30_U54 (.A4( us30_n818 ) , .A3( us30_n819 ) , .A2( us30_n820 ) , .A1( us30_n821 ) , .ZN( us30_n822 ) );
  AOI222_X1 us30_U55 (.C2( us30_n809 ) , .B2( us30_n810 ) , .A2( us30_n811 ) , .ZN( us30_n823 ) , .C1( us30_n832 ) , .A1( us30_n839 ) , .B1( us30_n853 ) );
  AOI211_X1 us30_U56 (.B( us30_n807 ) , .A( us30_n808 ) , .ZN( us30_n824 ) , .C1( us30_n842 ) , .C2( us30_n850 ) );
  NAND4_X1 us30_U57 (.ZN( sa31_sr_0 ) , .A4( us30_n501 ) , .A3( us30_n502 ) , .A2( us30_n503 ) , .A1( us30_n504 ) );
  AOI221_X1 us30_U58 (.A( us30_n497 ) , .ZN( us30_n502 ) , .B2( us30_n843 ) , .C1( us30_n846 ) , .C2( us30_n860 ) , .B1( us30_n862 ) );
  NOR4_X1 us30_U59 (.A4( us30_n498 ) , .A3( us30_n499 ) , .A2( us30_n500 ) , .ZN( us30_n501 ) , .A1( us30_n527 ) );
  NAND2_X1 us30_U6 (.A2( us30_n471 ) , .A1( us30_n472 ) , .ZN( us30_n817 ) );
  AOI211_X1 us30_U60 (.A( us30_n496 ) , .ZN( us30_n503 ) , .B( us30_n802 ) , .C2( us30_n839 ) , .C1( us30_n851 ) );
  NAND4_X1 us30_U61 (.ZN( sa31_sr_1 ) , .A4( us30_n595 ) , .A3( us30_n596 ) , .A2( us30_n597 ) , .A1( us30_n598 ) );
  NOR4_X1 us30_U62 (.A4( us30_n591 ) , .A3( us30_n592 ) , .A2( us30_n593 ) , .A1( us30_n594 ) , .ZN( us30_n595 ) );
  AOI211_X1 us30_U63 (.B( us30_n589 ) , .A( us30_n590 ) , .ZN( us30_n596 ) , .C2( us30_n811 ) , .C1( us30_n833 ) );
  AOI211_X1 us30_U64 (.A( us30_n588 ) , .ZN( us30_n597 ) , .B( us30_n621 ) , .C1( us30_n845 ) , .C2( us30_n855 ) );
  NOR2_X1 us30_U65 (.ZN( us30_n748 ) , .A1( us30_n861 ) , .A2( us30_n862 ) );
  NOR2_X1 us30_U66 (.ZN( us30_n625 ) , .A2( us30_n836 ) , .A1( us30_n839 ) );
  NAND4_X1 us30_U67 (.A4( us30_n603 ) , .A3( us30_n604 ) , .A2( us30_n605 ) , .A1( us30_n606 ) , .ZN( us30_n722 ) );
  NOR3_X1 us30_U68 (.A1( us30_n599 ) , .ZN( us30_n604 ) , .A3( us30_n663 ) , .A2( us30_n770 ) );
  NOR4_X1 us30_U69 (.A3( us30_n600 ) , .A2( us30_n601 ) , .A1( us30_n602 ) , .ZN( us30_n603 ) , .A4( us30_n655 ) );
  NOR3_X1 us30_U7 (.ZN( us30_n598 ) , .A1( us30_n608 ) , .A3( us30_n723 ) , .A2( us30_n742 ) );
  AOI222_X1 us30_U70 (.ZN( us30_n606 ) , .A1( us30_n830 ) , .C2( us30_n837 ) , .B1( us30_n842 ) , .A2( us30_n856 ) , .B2( us30_n861 ) , .C1( us30_n868 ) );
  NAND4_X1 us30_U71 (.A4( us30_n657 ) , .A3( us30_n658 ) , .A2( us30_n659 ) , .A1( us30_n660 ) , .ZN( us30_n800 ) );
  NOR3_X1 us30_U72 (.A3( us30_n648 ) , .A2( us30_n649 ) , .A1( us30_n650 ) , .ZN( us30_n659 ) );
  NOR3_X1 us30_U73 (.A3( us30_n651 ) , .A2( us30_n652 ) , .A1( us30_n653 ) , .ZN( us30_n658 ) );
  NOR3_X1 us30_U74 (.A3( us30_n654 ) , .A2( us30_n655 ) , .A1( us30_n656 ) , .ZN( us30_n657 ) );
  NAND4_X1 us30_U75 (.A4( us30_n560 ) , .A3( us30_n561 ) , .A2( us30_n562 ) , .A1( us30_n563 ) , .ZN( us30_n607 ) );
  NOR4_X1 us30_U76 (.ZN( us30_n561 ) , .A1( us30_n653 ) , .A3( us30_n661 ) , .A4( us30_n685 ) , .A2( us30_n768 ) );
  NOR4_X1 us30_U77 (.A4( us30_n552 ) , .A3( us30_n553 ) , .A2( us30_n554 ) , .A1( us30_n555 ) , .ZN( us30_n562 ) );
  NOR4_X1 us30_U78 (.A4( us30_n556 ) , .A3( us30_n557 ) , .A2( us30_n558 ) , .A1( us30_n559 ) , .ZN( us30_n560 ) );
  NAND4_X1 us30_U79 (.A4( us30_n772 ) , .A3( us30_n773 ) , .A2( us30_n774 ) , .A1( us30_n775 ) , .ZN( us30_n801 ) );
  NOR3_X1 us30_U8 (.A3( us30_n800 ) , .A2( us30_n801 ) , .A1( us30_n802 ) , .ZN( us30_n825 ) );
  NOR3_X1 us30_U80 (.A3( us30_n765 ) , .A2( us30_n766 ) , .A1( us30_n767 ) , .ZN( us30_n773 ) );
  NOR4_X1 us30_U81 (.A4( us30_n768 ) , .A3( us30_n769 ) , .A2( us30_n770 ) , .A1( us30_n771 ) , .ZN( us30_n772 ) );
  AOI222_X1 us30_U82 (.ZN( us30_n775 ) , .A1( us30_n830 ) , .C1( us30_n834 ) , .B2( us30_n841 ) , .A2( us30_n850 ) , .B1( us30_n861 ) , .C2( us30_n873 ) );
  NOR4_X1 us30_U83 (.A4( us30_n665 ) , .A3( us30_n666 ) , .A2( us30_n667 ) , .A1( us30_n668 ) , .ZN( us30_n676 ) );
  NOR4_X1 us30_U84 (.A4( us30_n661 ) , .A3( us30_n662 ) , .A2( us30_n663 ) , .A1( us30_n664 ) , .ZN( us30_n677 ) );
  NOR4_X1 us30_U85 (.A3( us30_n673 ) , .A1( us30_n674 ) , .ZN( us30_n675 ) , .A4( us30_n715 ) , .A2( us30_n859 ) );
  NOR2_X1 us30_U86 (.ZN( us30_n761 ) , .A1( us30_n833 ) , .A2( us30_n834 ) );
  NOR4_X1 us30_U87 (.A4( us30_n577 ) , .A3( us30_n578 ) , .A2( us30_n579 ) , .ZN( us30_n586 ) , .A1( us30_n683 ) );
  NOR4_X1 us30_U88 (.A1( us30_n584 ) , .ZN( us30_n585 ) , .A3( us30_n652 ) , .A2( us30_n662 ) , .A4( us30_n767 ) );
  AOI222_X1 us30_U89 (.ZN( us30_n513 ) , .C1( us30_n832 ) , .B2( us30_n837 ) , .A2( us30_n843 ) , .C2( us30_n862 ) , .B1( us30_n863 ) , .A1( us30_n866 ) );
  NOR3_X1 us30_U9 (.A3( us30_n621 ) , .A2( us30_n622 ) , .ZN( us30_n636 ) , .A1( us30_n725 ) );
  NOR4_X1 us30_U90 (.A4( us30_n509 ) , .A2( us30_n510 ) , .A1( us30_n511 ) , .ZN( us30_n512 ) , .A3( us30_n670 ) );
  INV_X1 us30_U91 (.A( us30_n505 ) , .ZN( us30_n871 ) );
  NAND4_X1 us30_U92 (.A4( us30_n456 ) , .A3( us30_n457 ) , .A2( us30_n458 ) , .A1( us30_n459 ) , .ZN( us30_n679 ) );
  NOR3_X1 us30_U93 (.ZN( us30_n457 ) , .A3( us30_n530 ) , .A1( us30_n555 ) , .A2( us30_n570 ) );
  AOI221_X1 us30_U94 (.A( us30_n450 ) , .ZN( us30_n459 ) , .C2( us30_n753 ) , .B1( us30_n832 ) , .C1( us30_n842 ) , .B2( us30_n861 ) );
  NOR4_X1 us30_U95 (.ZN( us30_n458 ) , .A2( us30_n509 ) , .A1( us30_n599 ) , .A4( us30_n628 ) , .A3( us30_n711 ) );
  NAND4_X1 us30_U96 (.A4( us30_n535 ) , .A3( us30_n536 ) , .A2( us30_n537 ) , .A1( us30_n538 ) , .ZN( us30_n622 ) );
  NOR4_X1 us30_U97 (.A4( us30_n526 ) , .A2( us30_n527 ) , .A1( us30_n528 ) , .ZN( us30_n538 ) , .A3( us30_n701 ) );
  NOR4_X1 us30_U98 (.A1( us30_n531 ) , .ZN( us30_n536 ) , .A2( us30_n654 ) , .A4( us30_n668 ) , .A3( us30_n765 ) );
  NOR4_X1 us30_U99 (.A4( us30_n529 ) , .A3( us30_n530 ) , .ZN( us30_n537 ) , .A2( us30_n684 ) , .A1( us30_n794 ) );
  NOR2_X1 us32_U10 (.A1( us32_n678 ) , .ZN( us32_n693 ) , .A2( us32_n807 ) );
  AOI211_X1 us32_U100 (.B( us32_n477 ) , .A( us32_n478 ) , .ZN( us32_n482 ) , .C2( us32_n833 ) , .C1( us32_n861 ) );
  NOR4_X1 us32_U101 (.ZN( us32_n481 ) , .A3( us32_n532 ) , .A4( us32_n545 ) , .A2( us32_n567 ) , .A1( us32_n717 ) );
  NAND4_X1 us32_U102 (.A4( us32_n548 ) , .A3( us32_n549 ) , .A2( us32_n550 ) , .A1( us32_n551 ) , .ZN( us32_n745 ) );
  NOR3_X1 us32_U103 (.ZN( us32_n549 ) , .A2( us32_n651 ) , .A1( us32_n667 ) , .A3( us32_n771 ) );
  AOI211_X1 us32_U104 (.B( us32_n539 ) , .A( us32_n540 ) , .ZN( us32_n551 ) , .C2( us32_n839 ) , .C1( us32_n851 ) );
  NOR4_X1 us32_U105 (.A4( us32_n541 ) , .A3( us32_n542 ) , .A2( us32_n543 ) , .ZN( us32_n550 ) , .A1( us32_n688 ) );
  NOR4_X1 us32_U106 (.ZN( us32_n620 ) , .A1( us32_n656 ) , .A3( us32_n666 ) , .A4( us32_n682 ) , .A2( us32_n766 ) );
  NOR4_X1 us32_U107 (.A4( us32_n609 ) , .A3( us32_n610 ) , .A2( us32_n611 ) , .A1( us32_n612 ) , .ZN( us32_n619 ) );
  NOR4_X1 us32_U108 (.A4( us32_n614 ) , .A3( us32_n615 ) , .A2( us32_n616 ) , .A1( us32_n617 ) , .ZN( us32_n618 ) );
  NOR2_X1 us32_U109 (.ZN( us32_n686 ) , .A1( us32_n831 ) , .A2( us32_n832 ) );
  NOR3_X1 us32_U11 (.ZN( us32_n504 ) , .A2( us32_n679 ) , .A3( us32_n777 ) , .A1( us32_n876 ) );
  NAND4_X1 us32_U110 (.A4( us32_n485 ) , .A3( us32_n486 ) , .A2( us32_n487 ) , .A1( us32_n488 ) , .ZN( us32_n778 ) );
  NOR4_X1 us32_U111 (.A4( us32_n484 ) , .ZN( us32_n487 ) , .A1( us32_n566 ) , .A2( us32_n581 ) , .A3( us32_n602 ) );
  NOR4_X1 us32_U112 (.ZN( us32_n486 ) , .A1( us32_n507 ) , .A2( us32_n519 ) , .A4( us32_n546 ) , .A3( us32_n611 ) );
  NOR4_X1 us32_U113 (.ZN( us32_n485 ) , .A2( us32_n533 ) , .A1( us32_n558 ) , .A3( us32_n631 ) , .A4( us32_n718 ) );
  NAND4_X1 us32_U114 (.A4( us32_n691 ) , .A3( us32_n692 ) , .A1( us32_n693 ) , .ZN( us32_n776 ) , .A2( us32_n872 ) );
  AOI221_X1 us32_U115 (.A( us32_n681 ) , .ZN( us32_n692 ) , .B2( us32_n840 ) , .C1( us32_n842 ) , .C2( us32_n862 ) , .B1( us32_n865 ) );
  INV_X1 us32_U116 (.A( us32_n679 ) , .ZN( us32_n872 ) );
  NOR4_X1 us32_U117 (.A4( us32_n687 ) , .A3( us32_n688 ) , .A2( us32_n689 ) , .A1( us32_n690 ) , .ZN( us32_n691 ) );
  NAND4_X1 us32_U118 (.A4( us32_n473 ) , .A3( us32_n474 ) , .A2( us32_n475 ) , .A1( us32_n476 ) , .ZN( us32_n678 ) );
  NOR4_X1 us32_U119 (.ZN( us32_n475 ) , .A1( us32_n531 ) , .A3( us32_n568 ) , .A4( us32_n600 ) , .A2( us32_n642 ) );
  INV_X1 us32_U12 (.A( us32_n706 ) , .ZN( us32_n876 ) );
  NOR4_X1 us32_U120 (.A4( us32_n470 ) , .ZN( us32_n476 ) , .A3( us32_n556 ) , .A1( us32_n735 ) , .A2( us32_n755 ) );
  NOR4_X1 us32_U121 (.ZN( us32_n473 ) , .A2( us32_n521 ) , .A4( us32_n594 ) , .A1( us32_n609 ) , .A3( us32_n629 ) );
  NAND4_X1 us32_U122 (.A4( us32_n719 ) , .A3( us32_n720 ) , .A2( us32_n721 ) , .ZN( us32_n741 ) , .A1( us32_n857 ) );
  INV_X1 us32_U123 (.A( us32_n709 ) , .ZN( us32_n857 ) );
  AOI221_X1 us32_U124 (.A( us32_n710 ) , .ZN( us32_n721 ) , .C2( us32_n844 ) , .B2( us32_n845 ) , .C1( us32_n861 ) , .B1( us32_n862 ) );
  NOR4_X1 us32_U125 (.A4( us32_n715 ) , .A3( us32_n716 ) , .A2( us32_n717 ) , .A1( us32_n718 ) , .ZN( us32_n719 ) );
  NOR2_X1 us32_U126 (.ZN( us32_n733 ) , .A2( us32_n832 ) , .A1( us32_n845 ) );
  NOR2_X1 us32_U127 (.ZN( us32_n789 ) , .A2( us32_n862 ) , .A1( us32_n868 ) );
  NAND4_X1 us32_U128 (.A4( us32_n573 ) , .A3( us32_n574 ) , .A1( us32_n575 ) , .ZN( us32_n723 ) , .A2( us32_n874 ) );
  AOI221_X1 us32_U129 (.A( us32_n564 ) , .C2( us32_n565 ) , .ZN( us32_n574 ) , .B2( us32_n845 ) , .B1( us32_n852 ) , .C1( us32_n853 ) );
  INV_X1 us32_U13 (.A( us32_n607 ) , .ZN( us32_n874 ) );
  NOR4_X1 us32_U130 (.A4( us32_n569 ) , .A3( us32_n570 ) , .A2( us32_n571 ) , .A1( us32_n572 ) , .ZN( us32_n573 ) );
  NOR2_X1 us32_U131 (.ZN( us32_n575 ) , .A1( us32_n622 ) , .A2( us32_n745 ) );
  NOR2_X1 us32_U132 (.ZN( us32_n748 ) , .A1( us32_n861 ) , .A2( us32_n862 ) );
  NAND4_X1 us32_U133 (.A4( us32_n633 ) , .A3( us32_n634 ) , .A2( us32_n635 ) , .A1( us32_n636 ) , .ZN( us32_n743 ) );
  AOI211_X1 us32_U134 (.B( us32_n623 ) , .A( us32_n624 ) , .ZN( us32_n635 ) , .C2( us32_n836 ) , .C1( us32_n863 ) );
  NOR4_X1 us32_U135 (.A4( us32_n629 ) , .A3( us32_n630 ) , .A2( us32_n631 ) , .A1( us32_n632 ) , .ZN( us32_n633 ) );
  NOR4_X1 us32_U136 (.A4( us32_n626 ) , .A3( us32_n627 ) , .A2( us32_n628 ) , .ZN( us32_n634 ) , .A1( us32_n664 ) );
  NAND4_X1 us32_U137 (.A4( us32_n493 ) , .A3( us32_n494 ) , .A1( us32_n495 ) , .ZN( us32_n802 ) , .A2( us32_n867 ) );
  AOI221_X1 us32_U138 (.A( us32_n489 ) , .ZN( us32_n494 ) , .B2( us32_n836 ) , .C2( us32_n841 ) , .C1( us32_n851 ) , .B1( us32_n860 ) );
  INV_X1 us32_U139 (.A( us32_n778 ) , .ZN( us32_n867 ) );
  INV_X1 us32_U14 (.A( us32_n680 ) , .ZN( us32_n840 ) );
  NOR4_X1 us32_U140 (.A2( us32_n491 ) , .A1( us32_n492 ) , .ZN( us32_n493 ) , .A3( us32_n580 ) , .A4( us32_n612 ) );
  NOR4_X1 us32_U141 (.A4( us32_n734 ) , .A3( us32_n735 ) , .A2( us32_n736 ) , .A1( us32_n737 ) , .ZN( us32_n738 ) );
  AOI211_X1 us32_U142 (.B( us32_n725 ) , .A( us32_n726 ) , .ZN( us32_n739 ) , .C1( us32_n843 ) , .C2( us32_n855 ) );
  NOR3_X1 us32_U143 (.A3( us32_n722 ) , .A1( us32_n723 ) , .ZN( us32_n740 ) , .A2( us32_n741 ) );
  NOR2_X1 us32_U144 (.ZN( us32_n647 ) , .A1( us32_n854 ) , .A2( us32_n868 ) );
  INV_X1 us32_U145 (.A( us32_n762 ) , .ZN( us32_n830 ) );
  INV_X1 us32_U146 (.A( us32_n754 ) , .ZN( us32_n869 ) );
  OAI21_X1 us32_U147 (.B1( us32_n753 ) , .ZN( us32_n754 ) , .A( us32_n845 ) , .B2( us32_n868 ) );
  INV_X1 us32_U148 (.A( us32_n697 ) , .ZN( us32_n838 ) );
  OR4_X1 us32_U149 (.ZN( us32_n492 ) , .A4( us32_n534 ) , .A2( us32_n547 ) , .A1( us32_n559 ) , .A3( us32_n632 ) );
  NOR4_X1 us32_U15 (.A4( us32_n445 ) , .A3( us32_n446 ) , .A2( us32_n516 ) , .A1( us32_n541 ) , .ZN( us32_n706 ) );
  OR4_X1 us32_U150 (.A4( us32_n566 ) , .A3( us32_n567 ) , .A2( us32_n568 ) , .ZN( us32_n572 ) , .A1( us32_n665 ) );
  OR4_X1 us32_U151 (.A4( us32_n682 ) , .A3( us32_n683 ) , .A2( us32_n684 ) , .A1( us32_n685 ) , .ZN( us32_n690 ) );
  OR4_X1 us32_U152 (.ZN( us32_n466 ) , .A4( us32_n518 ) , .A3( us32_n529 ) , .A2( us32_n578 ) , .A1( us32_n712 ) );
  OR4_X1 us32_U153 (.A4( us32_n518 ) , .A2( us32_n519 ) , .A1( us32_n520 ) , .ZN( us32_n522 ) , .A3( us32_n821 ) );
  OR4_X1 us32_U154 (.A4( us32_n580 ) , .A3( us32_n581 ) , .A2( us32_n582 ) , .A1( us32_n583 ) , .ZN( us32_n584 ) );
  NAND2_X1 us32_U155 (.ZN( us32_n613 ) , .A2( us32_n837 ) , .A1( us32_n873 ) );
  OR3_X1 us32_U156 (.A3( us32_n506 ) , .A2( us32_n507 ) , .A1( us32_n508 ) , .ZN( us32_n511 ) );
  INV_X1 us32_U157 (.A( us32_n672 ) , .ZN( us32_n859 ) );
  AOI21_X1 us32_U158 (.A( us32_n670 ) , .B1( us32_n671 ) , .ZN( us32_n672 ) , .B2( us32_n856 ) );
  INV_X1 us32_U159 (.A( us32_n463 ) , .ZN( us32_n864 ) );
  OR3_X1 us32_U16 (.ZN( us32_n446 ) , .A1( us32_n528 ) , .A3( us32_n577 ) , .A2( us32_n875 ) );
  OAI21_X1 us32_U160 (.ZN( us32_n463 ) , .B1( us32_n809 ) , .A( us32_n834 ) , .B2( us32_n851 ) );
  OAI222_X1 us32_U161 (.B2( us32_n708 ) , .ZN( us32_n709 ) , .C2( us32_n724 ) , .B1( us32_n747 ) , .A1( us32_n806 ) , .C1( us32_n814 ) , .A2( us32_n815 ) );
  NAND2_X1 us32_U162 (.A1( us32_n447 ) , .A2( us32_n465 ) , .ZN( us32_n749 ) );
  AOI22_X1 us32_U163 (.A2( us32_n782 ) , .ZN( us32_n783 ) , .B2( us32_n831 ) , .A1( us32_n834 ) , .B1( us32_n863 ) );
  AOI22_X1 us32_U164 (.ZN( us32_n696 ) , .A1( us32_n830 ) , .B2( us32_n843 ) , .A2( us32_n865 ) , .B1( us32_n868 ) );
  INV_X1 us32_U165 (.A( us32_n730 ) , .ZN( us32_n839 ) );
  AOI221_X1 us32_U166 (.A( us32_n483 ) , .ZN( us32_n488 ) , .B1( us32_n831 ) , .C2( us32_n844 ) , .C1( us32_n852 ) , .B2( us32_n862 ) );
  OAI22_X1 us32_U167 (.ZN( us32_n483 ) , .A1( us32_n708 ) , .B2( us32_n785 ) , .A2( us32_n806 ) , .B1( us32_n812 ) );
  INV_X1 us32_U168 (.A( us32_n790 ) , .ZN( us32_n832 ) );
  OAI221_X1 us32_U169 (.A( us32_n727 ) , .C2( us32_n728 ) , .B2( us32_n729 ) , .B1( us32_n730 ) , .ZN( us32_n737 ) , .C1( us32_n817 ) );
  OR4_X1 us32_U17 (.A4( us32_n442 ) , .A2( us32_n443 ) , .A1( us32_n444 ) , .ZN( us32_n445 ) , .A3( us32_n553 ) );
  AOI22_X1 us32_U170 (.ZN( us32_n727 ) , .B1( us32_n832 ) , .A2( us32_n838 ) , .A1( us32_n863 ) , .B2( us32_n866 ) );
  NAND2_X1 us32_U171 (.A1( us32_n451 ) , .A2( us32_n453 ) , .ZN( us32_n762 ) );
  INV_X1 us32_U172 (.A( us32_n786 ) , .ZN( us32_n862 ) );
  OAI22_X1 us32_U173 (.ZN( us32_n710 ) , .A2( us32_n728 ) , .B2( us32_n729 ) , .A1( us32_n744 ) , .B1( us32_n813 ) );
  INV_X1 us32_U174 (.A( us32_n816 ) , .ZN( us32_n831 ) );
  OAI22_X1 us32_U175 (.ZN( us32_n489 ) , .A1( us32_n724 ) , .B2( us32_n728 ) , .B1( us32_n730 ) , .A2( us32_n779 ) );
  OAI22_X1 us32_U176 (.ZN( us32_n624 ) , .B1( us32_n669 ) , .B2( us32_n747 ) , .A1( us32_n815 ) , .A2( us32_n816 ) );
  INV_X1 us32_U177 (.A( us32_n788 ) , .ZN( us32_n845 ) );
  OAI22_X1 us32_U178 (.A1( us32_n724 ) , .ZN( us32_n726 ) , .B2( us32_n750 ) , .B1( us32_n812 ) , .A2( us32_n816 ) );
  INV_X1 us32_U179 (.A( us32_n744 ) , .ZN( us32_n837 ) );
  INV_X1 us32_U18 (.A( us32_n613 ) , .ZN( us32_n875 ) );
  OAI22_X1 us32_U180 (.B2( us32_n779 ) , .B1( us32_n780 ) , .ZN( us32_n781 ) , .A2( us32_n814 ) , .A1( us32_n815 ) );
  INV_X1 us32_U181 (.A( us32_n814 ) , .ZN( us32_n833 ) );
  INV_X1 us32_U182 (.A( us32_n669 ) , .ZN( us32_n865 ) );
  OAI22_X1 us32_U183 (.B2( us32_n744 ) , .ZN( us32_n746 ) , .A2( us32_n762 ) , .B1( us32_n780 ) , .A1( us32_n792 ) );
  OAI22_X1 us32_U184 (.ZN( us32_n496 ) , .A2( us32_n744 ) , .A1( us32_n780 ) , .B1( us32_n791 ) , .B2( us32_n806 ) );
  AOI211_X1 us32_U185 (.A( us32_n637 ) , .ZN( us32_n645 ) , .B( us32_n743 ) , .C2( us32_n839 ) , .C1( us32_n854 ) );
  OAI22_X1 us32_U186 (.ZN( us32_n637 ) , .A1( us32_n699 ) , .B2( us32_n728 ) , .A2( us32_n762 ) , .B1( us32_n816 ) );
  INV_X1 us32_U187 (.A( us32_n750 ) , .ZN( us32_n842 ) );
  OAI22_X1 us32_U188 (.B1( us32_n490 ) , .ZN( us32_n491 ) , .A1( us32_n686 ) , .A2( us32_n763 ) , .B2( us32_n817 ) );
  NOR3_X1 us32_U189 (.ZN( us32_n490 ) , .A1( us32_n782 ) , .A2( us32_n850 ) , .A3( us32_n863 ) );
  INV_X1 us32_U19 (.A( us32_n749 ) , .ZN( us32_n863 ) );
  OAI22_X1 us32_U190 (.ZN( us32_n695 ) , .A2( us32_n730 ) , .A1( us32_n780 ) , .B1( us32_n791 ) , .B2( us32_n817 ) );
  NOR2_X1 us32_U191 (.ZN( us32_n666 ) , .A1( us32_n728 ) , .A2( us32_n803 ) );
  NOR2_X1 us32_U192 (.ZN( us32_n594 ) , .A2( us32_n697 ) , .A1( us32_n728 ) );
  NOR2_X1 us32_U193 (.ZN( us32_n570 ) , .A1( us32_n728 ) , .A2( us32_n806 ) );
  NOR2_X1 us32_U194 (.ZN( us32_n654 ) , .A1( us32_n728 ) , .A2( us32_n813 ) );
  NOR2_X1 us32_U195 (.ZN( us32_n546 ) , .A2( us32_n780 ) , .A1( us32_n814 ) );
  NOR2_X1 us32_U196 (.ZN( us32_n532 ) , .A2( us32_n749 ) , .A1( us32_n750 ) );
  NOR2_X1 us32_U197 (.ZN( us32_n577 ) , .A2( us32_n699 ) , .A1( us32_n814 ) );
  NOR2_X1 us32_U198 (.ZN( us32_n615 ) , .A1( us32_n785 ) , .A2( us32_n815 ) );
  NOR2_X1 us32_U199 (.ZN( us32_n629 ) , .A2( us32_n728 ) , .A1( us32_n785 ) );
  AOI222_X1 us32_U20 (.ZN( us32_n605 ) , .B2( us32_n671 ) , .B1( us32_n753 ) , .C2( us32_n831 ) , .A1( us32_n833 ) , .A2( us32_n862 ) , .C1( us32_n863 ) );
  NOR2_X1 us32_U200 (.ZN( us32_n718 ) , .A2( us32_n724 ) , .A1( us32_n744 ) );
  NOR2_X1 us32_U201 (.ZN( us32_n628 ) , .A2( us32_n669 ) , .A1( us32_n785 ) );
  INV_X1 us32_U202 (.A( us32_n728 ) , .ZN( us32_n852 ) );
  NOR2_X1 us32_U203 (.A2( us32_n744 ) , .ZN( us32_n769 ) , .A1( us32_n812 ) );
  NOR2_X1 us32_U204 (.ZN( us32_n531 ) , .A2( us32_n780 ) , .A1( us32_n816 ) );
  NOR2_X1 us32_U205 (.A2( us32_n708 ) , .A1( us32_n750 ) , .ZN( us32_n771 ) );
  NOR2_X1 us32_U206 (.ZN( us32_n599 ) , .A2( us32_n791 ) , .A1( us32_n816 ) );
  NOR2_X1 us32_U207 (.ZN( us32_n611 ) , .A2( us32_n780 ) , .A1( us32_n806 ) );
  NOR2_X1 us32_U208 (.ZN( us32_n652 ) , .A1( us32_n669 ) , .A2( us32_n814 ) );
  INV_X1 us32_U209 (.A( us32_n792 ) , .ZN( us32_n851 ) );
  AOI222_X1 us32_U21 (.ZN( us32_n563 ) , .B1( us32_n830 ) , .C1( us32_n841 ) , .A2( us32_n843 ) , .A1( us32_n854 ) , .B2( us32_n863 ) , .C2( us32_n873 ) );
  NOR2_X1 us32_U210 (.A1( us32_n699 ) , .ZN( us32_n768 ) , .A2( us32_n813 ) );
  NOR2_X1 us32_U211 (.A1( us32_n669 ) , .ZN( us32_n673 ) , .A2( us32_n744 ) );
  NOR2_X1 us32_U212 (.ZN( us32_n541 ) , .A2( us32_n697 ) , .A1( us32_n699 ) );
  NOR2_X1 us32_U213 (.ZN( us32_n602 ) , .A1( us32_n669 ) , .A2( us32_n803 ) );
  NOR2_X1 us32_U214 (.A1( us32_n669 ) , .ZN( us32_n688 ) , .A2( us32_n816 ) );
  NOR2_X1 us32_U215 (.ZN( us32_n667 ) , .A1( us32_n750 ) , .A2( us32_n815 ) );
  NOR2_X1 us32_U216 (.ZN( us32_n555 ) , .A1( us32_n750 ) , .A2( us32_n791 ) );
  NOR2_X1 us32_U217 (.ZN( us32_n508 ) , .A2( us32_n780 ) , .A1( us32_n785 ) );
  NOR2_X1 us32_U218 (.ZN( us32_n543 ) , .A2( us32_n708 ) , .A1( us32_n785 ) );
  INV_X1 us32_U219 (.A( us32_n747 ) , .ZN( us32_n834 ) );
  AOI222_X1 us32_U22 (.ZN( us32_n660 ) , .A2( us32_n839 ) , .B1( us32_n841 ) , .C2( us32_n845 ) , .A1( us32_n860 ) , .C1( us32_n863 ) , .B2( us32_n870 ) );
  NOR2_X1 us32_U220 (.ZN( us32_n664 ) , .A1( us32_n785 ) , .A2( us32_n791 ) );
  NOR2_X1 us32_U221 (.A1( us32_n669 ) , .ZN( us32_n766 ) , .A2( us32_n813 ) );
  NOR2_X1 us32_U222 (.ZN( us32_n527 ) , .A1( us32_n669 ) , .A2( us32_n779 ) );
  NOR2_X1 us32_U223 (.ZN( us32_n661 ) , .A1( us32_n729 ) , .A2( us32_n790 ) );
  NOR2_X1 us32_U224 (.ZN( us32_n601 ) , .A2( us32_n780 ) , .A1( us32_n803 ) );
  NOR2_X1 us32_U225 (.ZN( us32_n507 ) , .A1( us32_n812 ) , .A2( us32_n817 ) );
  NOR2_X1 us32_U226 (.ZN( us32_n528 ) , .A2( us32_n724 ) , .A1( us32_n803 ) );
  NOR2_X1 us32_U227 (.ZN( us32_n509 ) , .A1( us32_n729 ) , .A2( us32_n779 ) );
  NOR2_X1 us32_U228 (.ZN( us32_n557 ) , .A1( us32_n792 ) , .A2( us32_n814 ) );
  NOR2_X1 us32_U229 (.ZN( us32_n545 ) , .A1( us32_n749 ) , .A2( us32_n814 ) );
  INV_X1 us32_U23 (.A( us32_n647 ) , .ZN( us32_n870 ) );
  OAI22_X1 us32_U230 (.B1( us32_n440 ) , .ZN( us32_n444 ) , .A2( us32_n728 ) , .A1( us32_n744 ) , .B2( us32_n749 ) );
  NOR3_X1 us32_U231 (.ZN( us32_n440 ) , .A2( us32_n836 ) , .A3( us32_n837 ) , .A1( us32_n846 ) );
  NOR2_X1 us32_U232 (.ZN( us32_n662 ) , .A2( us32_n697 ) , .A1( us32_n729 ) );
  OAI22_X1 us32_U233 (.B2( us32_n750 ) , .B1( us32_n751 ) , .A1( us32_n752 ) , .ZN( us32_n756 ) , .A2( us32_n806 ) );
  NOR2_X1 us32_U234 (.ZN( us32_n751 ) , .A2( us32_n852 ) , .A1( us32_n860 ) );
  NOR3_X1 us32_U235 (.ZN( us32_n752 ) , .A2( us32_n853 ) , .A1( us32_n863 ) , .A3( us32_n865 ) );
  NOR2_X1 us32_U236 (.ZN( us32_n544 ) , .A2( us32_n785 ) , .A1( us32_n792 ) );
  NOR2_X1 us32_U237 (.ZN( us32_n663 ) , .A1( us32_n729 ) , .A2( us32_n785 ) );
  INV_X1 us32_U238 (.A( us32_n806 ) , .ZN( us32_n841 ) );
  NOR2_X1 us32_U239 (.ZN( us32_n506 ) , .A2( us32_n728 ) , .A1( us32_n762 ) );
  NOR4_X1 us32_U24 (.A4( us32_n544 ) , .A3( us32_n545 ) , .A2( us32_n546 ) , .A1( us32_n547 ) , .ZN( us32_n548 ) );
  NOR2_X1 us32_U240 (.ZN( us32_n631 ) , .A1( us32_n724 ) , .A2( us32_n813 ) );
  NOR2_X1 us32_U241 (.ZN( us32_n614 ) , .A1( us32_n762 ) , .A2( us32_n812 ) );
  NOR2_X1 us32_U242 (.ZN( us32_n530 ) , .A2( us32_n744 ) , .A1( us32_n792 ) );
  NOR2_X1 us32_U243 (.ZN( us32_n558 ) , .A1( us32_n708 ) , .A2( us32_n816 ) );
  NOR2_X1 us32_U244 (.ZN( us32_n516 ) , .A1( us32_n708 ) , .A2( us32_n744 ) );
  NOR2_X1 us32_U245 (.A2( us32_n697 ) , .ZN( us32_n716 ) , .A1( us32_n792 ) );
  NOR2_X1 us32_U246 (.A1( us32_n749 ) , .ZN( us32_n767 ) , .A2( us32_n803 ) );
  NOR2_X1 us32_U247 (.ZN( us32_n521 ) , .A1( us32_n790 ) , .A2( us32_n812 ) );
  NOR2_X1 us32_U248 (.ZN( us32_n655 ) , .A1( us32_n790 ) , .A2( us32_n815 ) );
  NOR2_X1 us32_U249 (.ZN( us32_n668 ) , .A2( us32_n708 ) , .A1( us32_n790 ) );
  NOR4_X1 us32_U25 (.ZN( us32_n479 ) , .A1( us32_n520 ) , .A4( us32_n557 ) , .A3( us32_n582 ) , .A2( us32_n630 ) );
  NOR2_X1 us32_U250 (.ZN( us32_n517 ) , .A1( us32_n708 ) , .A2( us32_n803 ) );
  INV_X1 us32_U251 (.A( us32_n763 ) , .ZN( us32_n866 ) );
  NOR2_X1 us32_U252 (.ZN( us32_n542 ) , .A1( us32_n762 ) , .A2( us32_n791 ) );
  NOR2_X1 us32_U253 (.ZN( us32_n630 ) , .A1( us32_n747 ) , .A2( us32_n815 ) );
  INV_X1 us32_U254 (.A( us32_n729 ) , .ZN( us32_n868 ) );
  NOR2_X1 us32_U255 (.ZN( us32_n609 ) , .A2( us32_n724 ) , .A1( us32_n817 ) );
  AOI21_X1 us32_U256 (.A( us32_n815 ) , .B2( us32_n816 ) , .B1( us32_n817 ) , .ZN( us32_n818 ) );
  NOR2_X1 us32_U257 (.ZN( us32_n579 ) , .A2( us32_n708 ) , .A1( us32_n730 ) );
  NOR2_X1 us32_U258 (.ZN( us32_n533 ) , .A2( us32_n724 ) , .A1( us32_n730 ) );
  NOR2_X1 us32_U259 (.ZN( us32_n642 ) , .A2( us32_n788 ) , .A1( us32_n791 ) );
  NOR4_X1 us32_U26 (.ZN( us32_n456 ) , .A2( us32_n517 ) , .A1( us32_n543 ) , .A3( us32_n579 ) , .A4( us32_n615 ) );
  AOI21_X1 us32_U260 (.B1( us32_n625 ) , .ZN( us32_n627 ) , .A( us32_n763 ) , .B2( us32_n814 ) );
  NOR2_X1 us32_U261 (.ZN( us32_n656 ) , .A1( us32_n747 ) , .A2( us32_n780 ) );
  AOI21_X1 us32_U262 (.A( us32_n812 ) , .B2( us32_n813 ) , .B1( us32_n814 ) , .ZN( us32_n819 ) );
  NOR2_X1 us32_U263 (.A2( us32_n697 ) , .A1( us32_n780 ) , .ZN( us32_n820 ) );
  AOI21_X1 us32_U264 (.ZN( us32_n499 ) , .B1( us32_n680 ) , .A( us32_n812 ) , .B2( us32_n816 ) );
  NOR2_X1 us32_U265 (.A2( us32_n708 ) , .A1( us32_n762 ) , .ZN( us32_n794 ) );
  AOI21_X1 us32_U266 (.ZN( us32_n593 ) , .B1( us32_n750 ) , .A( us32_n792 ) , .B2( us32_n813 ) );
  AOI21_X1 us32_U267 (.ZN( us32_n626 ) , .B2( us32_n669 ) , .A( us32_n790 ) , .B1( us32_n791 ) );
  NOR2_X1 us32_U268 (.ZN( us32_n520 ) , .A2( us32_n708 ) , .A1( us32_n814 ) );
  NOR2_X1 us32_U269 (.A1( us32_n697 ) , .ZN( us32_n770 ) , .A2( us32_n815 ) );
  NOR4_X1 us32_U27 (.A4( us32_n532 ) , .A3( us32_n533 ) , .A2( us32_n534 ) , .ZN( us32_n535 ) , .A1( us32_n820 ) );
  NOR2_X1 us32_U270 (.ZN( us32_n582 ) , .A1( us32_n744 ) , .A2( us32_n815 ) );
  NOR2_X1 us32_U271 (.ZN( us32_n519 ) , .A2( us32_n699 ) , .A1( us32_n816 ) );
  AOI21_X1 us32_U272 (.ZN( us32_n477 ) , .A( us32_n669 ) , .B1( us32_n750 ) , .B2( us32_n806 ) );
  AOI21_X1 us32_U273 (.ZN( us32_n510 ) , .B2( us32_n669 ) , .A( us32_n730 ) , .B1( us32_n815 ) );
  INV_X1 us32_U274 (.A( us32_n813 ) , .ZN( us32_n836 ) );
  AOI21_X1 us32_U275 (.ZN( us32_n589 ) , .B2( us32_n699 ) , .B1( us32_n815 ) , .A( us32_n817 ) );
  AOI21_X1 us32_U276 (.ZN( us32_n515 ) , .A( us32_n729 ) , .B1( us32_n750 ) , .B2( us32_n803 ) );
  AOI21_X1 us32_U277 (.ZN( us32_n539 ) , .B2( us32_n812 ) , .A( us32_n814 ) , .B1( us32_n815 ) );
  NOR2_X1 us32_U278 (.ZN( us32_n581 ) , .A1( us32_n669 ) , .A2( us32_n788 ) );
  NOR2_X1 us32_U279 (.ZN( us32_n547 ) , .A1( us32_n699 ) , .A2( us32_n744 ) );
  NOR4_X1 us32_U28 (.ZN( us32_n474 ) , .A1( us32_n506 ) , .A3( us32_n544 ) , .A2( us32_n583 ) , .A4( us32_n716 ) );
  AOI21_X1 us32_U280 (.ZN( us32_n540 ) , .A( us32_n763 ) , .B2( us32_n779 ) , .B1( us32_n817 ) );
  AOI21_X1 us32_U281 (.B1( us32_n699 ) , .ZN( us32_n700 ) , .A( us32_n732 ) , .B2( us32_n763 ) );
  AOI21_X1 us32_U282 (.ZN( us32_n591 ) , .B2( us32_n763 ) , .A( us32_n785 ) , .B1( us32_n812 ) );
  INV_X1 us32_U283 (.A( us32_n791 ) , .ZN( us32_n873 ) );
  NOR2_X1 us32_U284 (.ZN( us32_n559 ) , .A2( us32_n791 ) , .A1( us32_n803 ) );
  AOI21_X1 us32_U285 (.ZN( us32_n498 ) , .A( us32_n724 ) , .B2( us32_n762 ) , .B1( us32_n814 ) );
  NOR2_X1 us32_U286 (.ZN( us32_n683 ) , .A2( us32_n699 ) , .A1( us32_n803 ) );
  NOR2_X1 us32_U287 (.ZN( us32_n685 ) , .A1( us32_n729 ) , .A2( us32_n816 ) );
  AOI21_X1 us32_U288 (.B1( us32_n686 ) , .ZN( us32_n687 ) , .A( us32_n728 ) , .B2( us32_n761 ) );
  AOI21_X1 us32_U289 (.ZN( us32_n569 ) , .B1( us32_n750 ) , .B2( us32_n762 ) , .A( us32_n780 ) );
  AOI221_X1 us32_U29 (.A( us32_n713 ) , .B2( us32_n714 ) , .ZN( us32_n720 ) , .C1( us32_n832 ) , .B1( us32_n839 ) , .C2( us32_n863 ) );
  AOI21_X1 us32_U290 (.ZN( us32_n649 ) , .B1( us32_n729 ) , .B2( us32_n763 ) , .A( us32_n813 ) );
  NOR2_X1 us32_U291 (.ZN( us32_n568 ) , .A1( us32_n729 ) , .A2( us32_n762 ) );
  INV_X1 us32_U292 (.A( us32_n699 ) , .ZN( us32_n853 ) );
  NOR2_X1 us32_U293 (.ZN( us32_n566 ) , .A2( us32_n697 ) , .A1( us32_n763 ) );
  AOI21_X1 us32_U294 (.ZN( us32_n514 ) , .A( us32_n779 ) , .B2( us32_n792 ) , .B1( us32_n812 ) );
  AOI21_X1 us32_U295 (.ZN( us32_n639 ) , .B2( us32_n749 ) , .A( us32_n788 ) , .B1( us32_n812 ) );
  NOR2_X1 us32_U296 (.ZN( us32_n665 ) , .A1( us32_n780 ) , .A2( us32_n813 ) );
  AOI21_X1 us32_U297 (.ZN( us32_n571 ) , .B2( us32_n697 ) , .B1( us32_n806 ) , .A( us32_n812 ) );
  AOI21_X1 us32_U298 (.ZN( us32_n564 ) , .B1( us32_n724 ) , .A( us32_n779 ) , .B2( us32_n791 ) );
  AOI21_X1 us32_U299 (.ZN( us32_n497 ) , .A( us32_n779 ) , .B2( us32_n791 ) , .B1( us32_n804 ) );
  NAND2_X1 us32_U3 (.A1( us32_n449 ) , .A2( us32_n464 ) , .ZN( us32_n724 ) );
  OR2_X1 us32_U30 (.A2( us32_n711 ) , .A1( us32_n712 ) , .ZN( us32_n713 ) );
  AOI21_X1 us32_U300 (.ZN( us32_n640 ) , .B2( us32_n747 ) , .A( us32_n792 ) , .B1( us32_n803 ) );
  NOR2_X1 us32_U301 (.ZN( us32_n578 ) , .A1( us32_n708 ) , .A2( us32_n813 ) );
  NOR2_X1 us32_U302 (.ZN( us32_n529 ) , .A1( us32_n708 ) , .A2( us32_n779 ) );
  AOI21_X1 us32_U303 (.ZN( us32_n689 ) , .B2( us32_n749 ) , .B1( us32_n763 ) , .A( us32_n806 ) );
  AOI21_X1 us32_U304 (.A( us32_n790 ) , .B2( us32_n791 ) , .B1( us32_n792 ) , .ZN( us32_n793 ) );
  AOI21_X1 us32_U305 (.ZN( us32_n478 ) , .B2( us32_n697 ) , .A( us32_n749 ) , .B1( us32_n779 ) );
  NOR2_X1 us32_U306 (.ZN( us32_n684 ) , .A1( us32_n791 ) , .A2( us32_n813 ) );
  AOI21_X1 us32_U307 (.ZN( us32_n450 ) , .B2( us32_n792 ) , .A( us32_n803 ) , .B1( us32_n815 ) );
  AOI21_X1 us32_U308 (.A( us32_n733 ) , .ZN( us32_n734 ) , .B2( us32_n780 ) , .B1( us32_n792 ) );
  NOR2_X1 us32_U309 (.A2( us32_n813 ) , .A1( us32_n815 ) , .ZN( us32_n821 ) );
  NOR2_X1 us32_U31 (.ZN( us32_n680 ) , .A2( us32_n834 ) , .A1( us32_n839 ) );
  AOI21_X1 us32_U310 (.ZN( us32_n641 ) , .B1( us32_n680 ) , .A( us32_n791 ) , .B2( us32_n817 ) );
  NOR2_X1 us32_U311 (.ZN( us32_n583 ) , .A1( us32_n792 ) , .A2( us32_n817 ) );
  NOR2_X1 us32_U312 (.ZN( us32_n711 ) , .A1( us32_n762 ) , .A2( us32_n763 ) );
  NOR2_X1 us32_U313 (.ZN( us32_n534 ) , .A1( us32_n724 ) , .A2( us32_n788 ) );
  NOR2_X1 us32_U314 (.ZN( us32_n632 ) , .A2( us32_n697 ) , .A1( us32_n724 ) );
  NOR2_X1 us32_U315 (.ZN( us32_n580 ) , .A2( us32_n697 ) , .A1( us32_n791 ) );
  NOR2_X1 us32_U316 (.ZN( us32_n682 ) , .A2( us32_n708 ) , .A1( us32_n817 ) );
  INV_X1 us32_U317 (.A( us32_n815 ) , .ZN( us32_n855 ) );
  AOI21_X1 us32_U318 (.ZN( us32_n442 ) , .A( us32_n699 ) , .B1( us32_n733 ) , .B2( us32_n750 ) );
  INV_X1 us32_U319 (.A( us32_n780 ) , .ZN( us32_n850 ) );
  NOR4_X1 us32_U32 (.A4( us32_n514 ) , .A3( us32_n515 ) , .A2( us32_n516 ) , .A1( us32_n517 ) , .ZN( us32_n524 ) );
  INV_X1 us32_U320 (.A( us32_n785 ) , .ZN( us32_n846 ) );
  NAND2_X1 us32_U321 (.ZN( us32_n714 ) , .A1( us32_n728 ) , .A2( us32_n780 ) );
  NAND2_X1 us32_U322 (.ZN( us32_n671 ) , .A1( us32_n806 ) , .A2( us32_n816 ) );
  AOI21_X1 us32_U323 (.ZN( us32_n443 ) , .B1( us32_n789 ) , .B2( us32_n791 ) , .A( us32_n814 ) );
  NOR2_X1 us32_U324 (.ZN( us32_n470 ) , .A2( us32_n779 ) , .A1( us32_n815 ) );
  NAND2_X1 us32_U325 (.A2( us32_n762 ) , .A1( us32_n806 ) , .ZN( us32_n810 ) );
  NOR2_X1 us32_U326 (.ZN( us32_n526 ) , .A1( us32_n724 ) , .A2( us32_n750 ) );
  OAI21_X1 us32_U327 (.A( us32_n787 ) , .B2( us32_n788 ) , .B1( us32_n789 ) , .ZN( us32_n795 ) );
  OAI21_X1 us32_U328 (.ZN( us32_n787 ) , .A( us32_n839 ) , .B1( us32_n863 ) , .B2( us32_n873 ) );
  NAND2_X1 us32_U329 (.A1( us32_n699 ) , .A2( us32_n729 ) , .ZN( us32_n782 ) );
  AOI222_X1 us32_U33 (.ZN( us32_n525 ) , .A1( us32_n834 ) , .B2( us32_n837 ) , .C1( us32_n844 ) , .C2( us32_n850 ) , .A2( us32_n852 ) , .B1( us32_n866 ) );
  NOR2_X1 us32_U330 (.ZN( us32_n712 ) , .A2( us32_n724 ) , .A1( us32_n790 ) );
  NOR2_X1 us32_U331 (.ZN( us32_n518 ) , .A1( us32_n708 ) , .A2( us32_n788 ) );
  OAI21_X1 us32_U332 (.A( us32_n698 ) , .ZN( us32_n702 ) , .B2( us32_n750 ) , .B1( us32_n804 ) );
  OAI21_X1 us32_U333 (.ZN( us32_n698 ) , .B2( us32_n833 ) , .B1( us32_n838 ) , .A( us32_n860 ) );
  INV_X1 us32_U334 (.A( us32_n817 ) , .ZN( us32_n844 ) );
  INV_X1 us32_U335 (.A( us32_n724 ) , .ZN( us32_n856 ) );
  OAI21_X1 us32_U336 (.ZN( us32_n731 ) , .A( us32_n833 ) , .B2( us32_n852 ) , .B1( us32_n873 ) );
  AND2_X1 us32_U337 (.ZN( us32_n732 ) , .A1( us32_n779 ) , .A2( us32_n785 ) );
  AOI221_X1 us32_U338 (.A( us32_n764 ) , .ZN( us32_n774 ) , .C2( us32_n810 ) , .B2( us32_n835 ) , .C1( us32_n855 ) , .B1( us32_n866 ) );
  AOI21_X1 us32_U339 (.B2( us32_n763 ) , .ZN( us32_n764 ) , .A( us32_n788 ) , .B1( us32_n792 ) );
  NOR4_X1 us32_U34 (.A3( us32_n521 ) , .A1( us32_n522 ) , .ZN( us32_n523 ) , .A2( us32_n673 ) , .A4( us32_n769 ) );
  INV_X1 us32_U340 (.A( us32_n761 ) , .ZN( us32_n835 ) );
  NAND2_X1 us32_U341 (.A2( us32_n448 ) , .A1( us32_n460 ) , .ZN( us32_n728 ) );
  NAND2_X1 us32_U342 (.A1( us32_n451 ) , .A2( us32_n454 ) , .ZN( us32_n814 ) );
  NAND2_X1 us32_U343 (.A1( us32_n455 ) , .A2( us32_n462 ) , .ZN( us32_n750 ) );
  NAND2_X1 us32_U344 (.A1( us32_n451 ) , .A2( us32_n471 ) , .ZN( us32_n816 ) );
  NAND2_X1 us32_U345 (.A1( us32_n454 ) , .A2( us32_n461 ) , .ZN( us32_n813 ) );
  NAND2_X1 us32_U346 (.A1( us32_n452 ) , .A2( us32_n465 ) , .ZN( us32_n669 ) );
  NAND2_X1 us32_U347 (.A1( us32_n453 ) , .A2( us32_n472 ) , .ZN( us32_n785 ) );
  NAND2_X1 us32_U348 (.A1( us32_n453 ) , .A2( us32_n461 ) , .ZN( us32_n744 ) );
  NAND2_X1 us32_U349 (.A2( us32_n453 ) , .A1( us32_n455 ) , .ZN( us32_n806 ) );
  AOI221_X1 us32_U35 (.A( us32_n781 ) , .ZN( us32_n798 ) , .C2( us32_n837 ) , .B2( us32_n838 ) , .B1( us32_n865 ) , .C1( us32_n866 ) );
  NAND2_X1 us32_U350 (.A1( us32_n455 ) , .A2( us32_n471 ) , .ZN( us32_n803 ) );
  NAND2_X1 us32_U351 (.A2( us32_n454 ) , .A1( us32_n472 ) , .ZN( us32_n779 ) );
  NAND2_X1 us32_U352 (.A2( us32_n464 ) , .A1( us32_n465 ) , .ZN( us32_n812 ) );
  NAND2_X1 us32_U353 (.A1( us32_n441 ) , .A2( us32_n460 ) , .ZN( us32_n699 ) );
  NAND2_X1 us32_U354 (.A2( us32_n448 ) , .A1( us32_n452 ) , .ZN( us32_n729 ) );
  NAND2_X1 us32_U355 (.A2( us32_n449 ) , .A1( us32_n452 ) , .ZN( us32_n763 ) );
  NOR2_X1 us32_U356 (.ZN( us32_n465 ) , .A2( us32_n847 ) , .A1( us32_n848 ) );
  NOR2_X1 us32_U357 (.ZN( us32_n453 ) , .A1( us32_n826 ) , .A2( us32_n827 ) );
  NAND2_X1 us32_U358 (.A1( us32_n462 ) , .A2( us32_n472 ) , .ZN( us32_n788 ) );
  NOR2_X1 us32_U359 (.ZN( us32_n451 ) , .A1( us32_n828 ) , .A2( us32_n829 ) );
  NOR4_X1 us32_U36 (.A4( us32_n793 ) , .A3( us32_n794 ) , .A2( us32_n795 ) , .A1( us32_n796 ) , .ZN( us32_n797 ) );
  NAND2_X1 us32_U360 (.A2( us32_n461 ) , .A1( us32_n462 ) , .ZN( us32_n747 ) );
  NAND2_X1 us32_U361 (.A1( us32_n451 ) , .A2( us32_n462 ) , .ZN( us32_n790 ) );
  NAND2_X2 us32_U362 (.A2( us32_n448 ) , .A1( us32_n464 ) , .ZN( us32_n815 ) );
  NAND2_X1 us32_U363 (.A2( us32_n441 ) , .A1( us32_n447 ) , .ZN( us32_n784 ) );
  NAND2_X1 us32_U364 (.A1( us32_n447 ) , .A2( us32_n449 ) , .ZN( us32_n805 ) );
  NAND2_X1 us32_U365 (.A2( us32_n454 ) , .A1( us32_n455 ) , .ZN( us32_n730 ) );
  NAND2_X2 us32_U366 (.A1( us32_n449 ) , .A2( us32_n460 ) , .ZN( us32_n792 ) );
  NAND2_X2 us32_U367 (.A2( us32_n460 ) , .A1( us32_n465 ) , .ZN( us32_n780 ) );
  NOR2_X1 us32_U368 (.ZN( us32_n447 ) , .A2( us32_n849 ) , .A1( us32_n858 ) );
  NAND2_X1 us32_U369 (.A1( us32_n447 ) , .A2( us32_n448 ) , .ZN( us32_n786 ) );
  NOR4_X1 us32_U37 (.A4( us32_n776 ) , .A3( us32_n777 ) , .A1( us32_n778 ) , .ZN( us32_n799 ) , .A2( us32_n801 ) );
  NAND2_X1 us32_U370 (.A2( us32_n471 ) , .A1( us32_n472 ) , .ZN( us32_n817 ) );
  NOR2_X1 us32_U371 (.A2( sa32_6 ) , .A1( sa32_7 ) , .ZN( us32_n464 ) );
  NOR2_X1 us32_U372 (.A2( sa32_7 ) , .ZN( us32_n460 ) , .A1( us32_n849 ) );
  NOR2_X1 us32_U373 (.A2( sa32_4 ) , .ZN( us32_n449 ) , .A1( us32_n848 ) );
  NOR2_X1 us32_U374 (.A2( sa32_4 ) , .A1( sa32_5 ) , .ZN( us32_n441 ) );
  NOR2_X1 us32_U375 (.A2( sa32_5 ) , .ZN( us32_n448 ) , .A1( us32_n847 ) );
  NOR2_X1 us32_U376 (.A2( sa32_2 ) , .A1( sa32_3 ) , .ZN( us32_n472 ) );
  NOR2_X1 us32_U377 (.A2( sa32_6 ) , .ZN( us32_n452 ) , .A1( us32_n858 ) );
  NOR2_X1 us32_U378 (.A2( sa32_1 ) , .ZN( us32_n471 ) , .A1( us32_n826 ) );
  NOR2_X1 us32_U379 (.A2( sa32_0 ) , .ZN( us32_n454 ) , .A1( us32_n827 ) );
  NOR4_X1 us32_U38 (.A3( us32_n755 ) , .A2( us32_n756 ) , .A1( us32_n757 ) , .ZN( us32_n758 ) , .A4( us32_n869 ) );
  NOR2_X1 us32_U380 (.A2( sa32_0 ) , .A1( sa32_1 ) , .ZN( us32_n462 ) );
  NOR2_X1 us32_U381 (.A2( sa32_3 ) , .ZN( us32_n455 ) , .A1( us32_n828 ) );
  NOR2_X1 us32_U382 (.A2( sa32_2 ) , .ZN( us32_n461 ) , .A1( us32_n829 ) );
  INV_X1 us32_U383 (.A( sa32_4 ) , .ZN( us32_n847 ) );
  INV_X1 us32_U384 (.A( sa32_6 ) , .ZN( us32_n849 ) );
  INV_X1 us32_U385 (.A( sa32_3 ) , .ZN( us32_n829 ) );
  INV_X1 us32_U386 (.A( sa32_1 ) , .ZN( us32_n827 ) );
  INV_X1 us32_U387 (.A( sa32_0 ) , .ZN( us32_n826 ) );
  INV_X1 us32_U388 (.A( sa32_2 ) , .ZN( us32_n828 ) );
  INV_X1 us32_U389 (.A( sa32_5 ) , .ZN( us32_n848 ) );
  AOI211_X1 us32_U39 (.B( us32_n745 ) , .A( us32_n746 ) , .ZN( us32_n759 ) , .C1( us32_n832 ) , .C2( us32_n853 ) );
  INV_X1 us32_U390 (.A( sa32_7 ) , .ZN( us32_n858 ) );
  NAND2_X1 us32_U391 (.A2( us32_n461 ) , .A1( us32_n471 ) , .ZN( us32_n697 ) );
  OAI222_X1 us32_U392 (.B2( us32_n747 ) , .B1( us32_n748 ) , .A2( us32_n749 ) , .ZN( us32_n757 ) , .C2( us32_n805 ) , .C1( us32_n814 ) , .A1( us32_n817 ) );
  OAI22_X1 us32_U393 (.B2( us32_n803 ) , .B1( us32_n804 ) , .A2( us32_n805 ) , .A1( us32_n806 ) , .ZN( us32_n808 ) );
  OAI21_X1 us32_U394 (.A( us32_n731 ) , .B1( us32_n732 ) , .ZN( us32_n736 ) , .B2( us32_n805 ) );
  OAI222_X1 us32_U395 (.ZN( us32_n505 ) , .C2( us32_n625 ) , .B2( us32_n647 ) , .B1( us32_n747 ) , .A2( us32_n748 ) , .C1( us32_n805 ) , .A1( us32_n806 ) );
  AOI21_X1 us32_U396 (.ZN( us32_n650 ) , .A( us32_n779 ) , .B1( us32_n792 ) , .B2( us32_n805 ) );
  INV_X1 us32_U397 (.A( us32_n805 ) , .ZN( us32_n860 ) );
  NOR2_X1 us32_U398 (.ZN( us32_n735 ) , .A2( us32_n803 ) , .A1( us32_n805 ) );
  NOR2_X1 us32_U399 (.ZN( us32_n484 ) , .A1( us32_n788 ) , .A2( us32_n805 ) );
  NAND2_X1 us32_U4 (.A1( us32_n441 ) , .A2( us32_n464 ) , .ZN( us32_n708 ) );
  NOR3_X1 us32_U40 (.A3( us32_n741 ) , .A2( us32_n742 ) , .A1( us32_n743 ) , .ZN( us32_n760 ) );
  NOR2_X1 us32_U400 (.A2( us32_n744 ) , .ZN( us32_n755 ) , .A1( us32_n805 ) );
  NAND2_X1 us32_U401 (.ZN( us32_n753 ) , .A1( us32_n763 ) , .A2( us32_n805 ) );
  NOR2_X1 us32_U402 (.ZN( us32_n715 ) , .A1( us32_n805 ) , .A2( us32_n817 ) );
  NOR2_X1 us32_U403 (.ZN( us32_n567 ) , .A1( us32_n747 ) , .A2( us32_n805 ) );
  AOI21_X1 us32_U404 (.ZN( us32_n552 ) , .B1( us32_n669 ) , .A( us32_n697 ) , .B2( us32_n805 ) );
  NOR2_X1 us32_U405 (.ZN( us32_n556 ) , .A1( us32_n762 ) , .A2( us32_n805 ) );
  NOR2_X1 us32_U406 (.ZN( us32_n670 ) , .A1( us32_n790 ) , .A2( us32_n805 ) );
  OAI221_X1 us32_U407 (.A( us32_n783 ) , .C2( us32_n784 ) , .B2( us32_n785 ) , .B1( us32_n786 ) , .ZN( us32_n796 ) , .C1( us32_n813 ) );
  NAND2_X1 us32_U408 (.A1( us32_n729 ) , .A2( us32_n784 ) , .ZN( us32_n811 ) );
  OAI22_X1 us32_U409 (.ZN( us32_n588 ) , .A2( us32_n747 ) , .B2( us32_n762 ) , .A1( us32_n763 ) , .B1( us32_n784 ) );
  NAND4_X1 us32_U41 (.ZN( sa33_sr_3 ) , .A4( us32_n704 ) , .A3( us32_n705 ) , .A2( us32_n706 ) , .A1( us32_n707 ) );
  AOI21_X1 us32_U410 (.ZN( us32_n592 ) , .B1( us32_n728 ) , .B2( us32_n784 ) , .A( us32_n790 ) );
  AOI21_X1 us32_U411 (.ZN( us32_n623 ) , .B1( us32_n699 ) , .A( us32_n779 ) , .B2( us32_n784 ) );
  AOI21_X1 us32_U412 (.ZN( us32_n648 ) , .A( us32_n762 ) , .B2( us32_n784 ) , .B1( us32_n792 ) );
  OAI22_X1 us32_U413 (.ZN( us32_n681 ) , .A1( us32_n699 ) , .A2( us32_n730 ) , .B2( us32_n784 ) , .B1( us32_n817 ) );
  OAI21_X1 us32_U414 (.A( us32_n613 ) , .ZN( us32_n616 ) , .B1( us32_n625 ) , .B2( us32_n784 ) );
  NOR2_X1 us32_U415 (.ZN( us32_n610 ) , .A1( us32_n784 ) , .A2( us32_n816 ) );
  OAI222_X1 us32_U416 (.A2( us32_n669 ) , .ZN( us32_n674 ) , .B1( us32_n747 ) , .B2( us32_n784 ) , .C2( us32_n788 ) , .C1( us32_n815 ) , .A1( us32_n817 ) );
  NOR2_X1 us32_U417 (.ZN( us32_n651 ) , .A1( us32_n784 ) , .A2( us32_n788 ) );
  NOR2_X1 us32_U418 (.ZN( us32_n600 ) , .A2( us32_n697 ) , .A1( us32_n784 ) );
  NOR2_X1 us32_U419 (.ZN( us32_n553 ) , .A2( us32_n744 ) , .A1( us32_n784 ) );
  NOR4_X1 us32_U42 (.A4( us32_n700 ) , .A3( us32_n701 ) , .A2( us32_n702 ) , .A1( us32_n703 ) , .ZN( us32_n704 ) );
  INV_X1 us32_U420 (.A( us32_n784 ) , .ZN( us32_n861 ) );
  AOI21_X1 us32_U421 (.ZN( us32_n500 ) , .A( us32_n697 ) , .B1( us32_n708 ) , .B2( us32_n786 ) );
  OAI221_X1 us32_U422 (.A( us32_n696 ) , .ZN( us32_n703 ) , .C2( us32_n784 ) , .C1( us32_n785 ) , .B1( us32_n786 ) , .B2( us32_n806 ) );
  OAI22_X1 us32_U423 (.ZN( us32_n590 ) , .B1( us32_n730 ) , .B2( us32_n749 ) , .A2( us32_n786 ) , .A1( us32_n803 ) );
  NOR2_X1 us32_U424 (.ZN( us32_n612 ) , .A1( us32_n779 ) , .A2( us32_n786 ) );
  NAND2_X1 us32_U425 (.A2( us32_n749 ) , .A1( us32_n786 ) , .ZN( us32_n809 ) );
  OAI222_X1 us32_U426 (.ZN( us32_n617 ) , .B1( us32_n697 ) , .C1( us32_n724 ) , .C2( us32_n747 ) , .B2( us32_n786 ) , .A2( us32_n792 ) , .A1( us32_n816 ) );
  NOR2_X1 us32_U427 (.ZN( us32_n717 ) , .A2( us32_n744 ) , .A1( us32_n786 ) );
  NOR2_X1 us32_U428 (.ZN( us32_n653 ) , .A1( us32_n762 ) , .A2( us32_n786 ) );
  NOR2_X1 us32_U429 (.ZN( us32_n554 ) , .A1( us32_n786 ) , .A2( us32_n813 ) );
  AOI211_X1 us32_U43 (.B( us32_n694 ) , .A( us32_n695 ) , .ZN( us32_n705 ) , .C2( us32_n831 ) , .C1( us32_n851 ) );
  NOR2_X1 us32_U430 (.ZN( us32_n701 ) , .A2( us32_n786 ) , .A1( us32_n817 ) );
  NOR2_X1 us32_U431 (.A1( us32_n730 ) , .ZN( us32_n765 ) , .A2( us32_n786 ) );
  AND2_X1 us32_U432 (.ZN( us32_n438 ) , .A2( us32_n831 ) , .A1( us32_n854 ) );
  AND2_X1 us32_U433 (.ZN( us32_n439 ) , .A2( us32_n843 ) , .A1( us32_n861 ) );
  NOR3_X1 us32_U434 (.A1( us32_n438 ) , .A2( us32_n439 ) , .A3( us32_n576 ) , .ZN( us32_n587 ) );
  NAND4_X1 us32_U435 (.ZN( sa33_sr_2 ) , .A4( us32_n643 ) , .A3( us32_n644 ) , .A2( us32_n645 ) , .A1( us32_n646 ) );
  INV_X1 us32_U436 (.A( us32_n812 ) , .ZN( us32_n854 ) );
  NAND3_X1 us32_U437 (.ZN( sa33_sr_6 ) , .A3( us32_n797 ) , .A2( us32_n798 ) , .A1( us32_n799 ) );
  NAND3_X1 us32_U438 (.ZN( sa33_sr_5 ) , .A3( us32_n758 ) , .A2( us32_n759 ) , .A1( us32_n760 ) );
  NAND3_X1 us32_U439 (.ZN( sa33_sr_4 ) , .A3( us32_n738 ) , .A2( us32_n739 ) , .A1( us32_n740 ) );
  NOR2_X1 us32_U44 (.ZN( us32_n707 ) , .A2( us32_n776 ) , .A1( us32_n800 ) );
  NAND3_X1 us32_U440 (.A3( us32_n675 ) , .A2( us32_n676 ) , .A1( us32_n677 ) , .ZN( us32_n807 ) );
  NAND3_X1 us32_U441 (.ZN( us32_n638 ) , .A3( us32_n708 ) , .A2( us32_n724 ) , .A1( us32_n792 ) );
  NAND3_X1 us32_U442 (.A3( us32_n618 ) , .A2( us32_n619 ) , .A1( us32_n620 ) , .ZN( us32_n725 ) );
  NAND3_X1 us32_U443 (.A3( us32_n585 ) , .A2( us32_n586 ) , .A1( us32_n587 ) , .ZN( us32_n621 ) );
  NAND3_X1 us32_U444 (.ZN( us32_n565 ) , .A3( us32_n680 ) , .A2( us32_n750 ) , .A1( us32_n785 ) );
  NAND3_X1 us32_U445 (.A3( us32_n523 ) , .A2( us32_n524 ) , .A1( us32_n525 ) , .ZN( us32_n742 ) );
  NAND3_X1 us32_U446 (.A3( us32_n512 ) , .A1( us32_n513 ) , .ZN( us32_n608 ) , .A2( us32_n871 ) );
  NAND3_X1 us32_U447 (.A3( us32_n467 ) , .A2( us32_n468 ) , .A1( us32_n469 ) , .ZN( us32_n777 ) );
  INV_X1 us32_U448 (.A( us32_n803 ) , .ZN( us32_n843 ) );
  AOI21_X1 us32_U449 (.ZN( us32_n576 ) , .B2( us32_n724 ) , .B1( us32_n748 ) , .A( us32_n785 ) );
  AOI222_X1 us32_U45 (.B2( us32_n638 ) , .ZN( us32_n644 ) , .B1( us32_n841 ) , .A1( us32_n842 ) , .C2( us32_n846 ) , .C1( us32_n863 ) , .A2( us32_n865 ) );
  NOR4_X1 us32_U46 (.A4( us32_n639 ) , .A3( us32_n640 ) , .A2( us32_n641 ) , .A1( us32_n642 ) , .ZN( us32_n643 ) );
  NOR3_X1 us32_U47 (.A2( us32_n607 ) , .A1( us32_n608 ) , .ZN( us32_n646 ) , .A3( us32_n722 ) );
  NAND4_X1 us32_U48 (.ZN( sa33_sr_7 ) , .A4( us32_n822 ) , .A3( us32_n823 ) , .A2( us32_n824 ) , .A1( us32_n825 ) );
  NOR4_X1 us32_U49 (.A4( us32_n818 ) , .A3( us32_n819 ) , .A2( us32_n820 ) , .A1( us32_n821 ) , .ZN( us32_n822 ) );
  NAND2_X1 us32_U5 (.A2( us32_n441 ) , .A1( us32_n452 ) , .ZN( us32_n791 ) );
  AOI222_X1 us32_U50 (.C2( us32_n809 ) , .B2( us32_n810 ) , .A2( us32_n811 ) , .ZN( us32_n823 ) , .C1( us32_n832 ) , .A1( us32_n839 ) , .B1( us32_n853 ) );
  AOI211_X1 us32_U51 (.B( us32_n807 ) , .A( us32_n808 ) , .ZN( us32_n824 ) , .C1( us32_n842 ) , .C2( us32_n850 ) );
  NAND4_X1 us32_U52 (.ZN( sa33_sr_0 ) , .A4( us32_n501 ) , .A3( us32_n502 ) , .A2( us32_n503 ) , .A1( us32_n504 ) );
  AOI221_X1 us32_U53 (.A( us32_n497 ) , .ZN( us32_n502 ) , .B2( us32_n843 ) , .C1( us32_n846 ) , .C2( us32_n860 ) , .B1( us32_n862 ) );
  NOR4_X1 us32_U54 (.A4( us32_n498 ) , .A3( us32_n499 ) , .A2( us32_n500 ) , .ZN( us32_n501 ) , .A1( us32_n527 ) );
  AOI211_X1 us32_U55 (.A( us32_n496 ) , .ZN( us32_n503 ) , .B( us32_n802 ) , .C2( us32_n839 ) , .C1( us32_n851 ) );
  NAND4_X1 us32_U56 (.ZN( sa33_sr_1 ) , .A4( us32_n595 ) , .A3( us32_n596 ) , .A2( us32_n597 ) , .A1( us32_n598 ) );
  NOR4_X1 us32_U57 (.A4( us32_n591 ) , .A3( us32_n592 ) , .A2( us32_n593 ) , .A1( us32_n594 ) , .ZN( us32_n595 ) );
  AOI211_X1 us32_U58 (.B( us32_n589 ) , .A( us32_n590 ) , .ZN( us32_n596 ) , .C2( us32_n811 ) , .C1( us32_n833 ) );
  AOI211_X1 us32_U59 (.A( us32_n588 ) , .ZN( us32_n597 ) , .B( us32_n621 ) , .C1( us32_n845 ) , .C2( us32_n855 ) );
  NOR3_X1 us32_U6 (.ZN( us32_n598 ) , .A1( us32_n608 ) , .A3( us32_n723 ) , .A2( us32_n742 ) );
  NOR2_X1 us32_U60 (.ZN( us32_n804 ) , .A1( us32_n854 ) , .A2( us32_n861 ) );
  AOI222_X1 us32_U61 (.ZN( us32_n469 ) , .B1( us32_n832 ) , .A1( us32_n839 ) , .C1( us32_n842 ) , .C2( us32_n851 ) , .A2( us32_n855 ) , .B2( us32_n865 ) );
  NOR4_X1 us32_U62 (.A1( us32_n466 ) , .ZN( us32_n467 ) , .A4( us32_n542 ) , .A2( us32_n554 ) , .A3( us32_n614 ) );
  AOI221_X1 us32_U63 (.ZN( us32_n468 ) , .C2( us32_n714 ) , .B2( us32_n831 ) , .C1( us32_n845 ) , .B1( us32_n860 ) , .A( us32_n864 ) );
  NAND4_X1 us32_U64 (.A4( us32_n603 ) , .A3( us32_n604 ) , .A2( us32_n605 ) , .A1( us32_n606 ) , .ZN( us32_n722 ) );
  NOR3_X1 us32_U65 (.A1( us32_n599 ) , .ZN( us32_n604 ) , .A3( us32_n663 ) , .A2( us32_n770 ) );
  NOR4_X1 us32_U66 (.A3( us32_n600 ) , .A2( us32_n601 ) , .A1( us32_n602 ) , .ZN( us32_n603 ) , .A4( us32_n655 ) );
  AOI222_X1 us32_U67 (.ZN( us32_n606 ) , .A1( us32_n830 ) , .C2( us32_n837 ) , .B1( us32_n842 ) , .A2( us32_n856 ) , .B2( us32_n861 ) , .C1( us32_n868 ) );
  NAND4_X1 us32_U68 (.A4( us32_n657 ) , .A3( us32_n658 ) , .A2( us32_n659 ) , .A1( us32_n660 ) , .ZN( us32_n800 ) );
  NOR3_X1 us32_U69 (.A3( us32_n648 ) , .A2( us32_n649 ) , .A1( us32_n650 ) , .ZN( us32_n659 ) );
  NOR3_X1 us32_U7 (.A3( us32_n800 ) , .A2( us32_n801 ) , .A1( us32_n802 ) , .ZN( us32_n825 ) );
  NOR3_X1 us32_U70 (.A3( us32_n651 ) , .A2( us32_n652 ) , .A1( us32_n653 ) , .ZN( us32_n658 ) );
  NOR3_X1 us32_U71 (.A3( us32_n654 ) , .A2( us32_n655 ) , .A1( us32_n656 ) , .ZN( us32_n657 ) );
  NAND4_X1 us32_U72 (.A4( us32_n560 ) , .A3( us32_n561 ) , .A2( us32_n562 ) , .A1( us32_n563 ) , .ZN( us32_n607 ) );
  NOR4_X1 us32_U73 (.A4( us32_n556 ) , .A3( us32_n557 ) , .A2( us32_n558 ) , .A1( us32_n559 ) , .ZN( us32_n560 ) );
  NOR4_X1 us32_U74 (.ZN( us32_n561 ) , .A1( us32_n653 ) , .A3( us32_n661 ) , .A4( us32_n685 ) , .A2( us32_n768 ) );
  NOR4_X1 us32_U75 (.A4( us32_n552 ) , .A3( us32_n553 ) , .A2( us32_n554 ) , .A1( us32_n555 ) , .ZN( us32_n562 ) );
  NAND4_X1 us32_U76 (.A4( us32_n772 ) , .A3( us32_n773 ) , .A2( us32_n774 ) , .A1( us32_n775 ) , .ZN( us32_n801 ) );
  NOR3_X1 us32_U77 (.A3( us32_n765 ) , .A2( us32_n766 ) , .A1( us32_n767 ) , .ZN( us32_n773 ) );
  NOR4_X1 us32_U78 (.A4( us32_n768 ) , .A3( us32_n769 ) , .A2( us32_n770 ) , .A1( us32_n771 ) , .ZN( us32_n772 ) );
  AOI222_X1 us32_U79 (.ZN( us32_n775 ) , .A1( us32_n830 ) , .C1( us32_n834 ) , .B2( us32_n841 ) , .A2( us32_n850 ) , .B1( us32_n861 ) , .C2( us32_n873 ) );
  NOR3_X1 us32_U8 (.A3( us32_n621 ) , .A2( us32_n622 ) , .ZN( us32_n636 ) , .A1( us32_n725 ) );
  NOR4_X1 us32_U80 (.A4( us32_n665 ) , .A3( us32_n666 ) , .A2( us32_n667 ) , .A1( us32_n668 ) , .ZN( us32_n676 ) );
  NOR4_X1 us32_U81 (.A4( us32_n661 ) , .A3( us32_n662 ) , .A2( us32_n663 ) , .A1( us32_n664 ) , .ZN( us32_n677 ) );
  NOR4_X1 us32_U82 (.A3( us32_n673 ) , .A1( us32_n674 ) , .ZN( us32_n675 ) , .A4( us32_n715 ) , .A2( us32_n859 ) );
  NOR2_X1 us32_U83 (.ZN( us32_n625 ) , .A2( us32_n836 ) , .A1( us32_n839 ) );
  NOR2_X1 us32_U84 (.ZN( us32_n761 ) , .A1( us32_n833 ) , .A2( us32_n834 ) );
  NOR4_X1 us32_U85 (.A4( us32_n577 ) , .A3( us32_n578 ) , .A2( us32_n579 ) , .ZN( us32_n586 ) , .A1( us32_n683 ) );
  NOR4_X1 us32_U86 (.A1( us32_n584 ) , .ZN( us32_n585 ) , .A3( us32_n652 ) , .A2( us32_n662 ) , .A4( us32_n767 ) );
  AOI222_X1 us32_U87 (.ZN( us32_n513 ) , .C1( us32_n832 ) , .B2( us32_n837 ) , .A2( us32_n843 ) , .C2( us32_n862 ) , .B1( us32_n863 ) , .A1( us32_n866 ) );
  NOR4_X1 us32_U88 (.A4( us32_n509 ) , .A2( us32_n510 ) , .A1( us32_n511 ) , .ZN( us32_n512 ) , .A3( us32_n670 ) );
  INV_X1 us32_U89 (.A( us32_n505 ) , .ZN( us32_n871 ) );
  NOR2_X1 us32_U9 (.ZN( us32_n495 ) , .A1( us32_n678 ) , .A2( us32_n694 ) );
  NAND4_X1 us32_U90 (.A4( us32_n456 ) , .A3( us32_n457 ) , .A2( us32_n458 ) , .A1( us32_n459 ) , .ZN( us32_n679 ) );
  NOR3_X1 us32_U91 (.ZN( us32_n457 ) , .A3( us32_n530 ) , .A1( us32_n555 ) , .A2( us32_n570 ) );
  AOI221_X1 us32_U92 (.A( us32_n450 ) , .ZN( us32_n459 ) , .C2( us32_n753 ) , .B1( us32_n832 ) , .C1( us32_n842 ) , .B2( us32_n861 ) );
  NOR4_X1 us32_U93 (.ZN( us32_n458 ) , .A2( us32_n509 ) , .A1( us32_n599 ) , .A4( us32_n628 ) , .A3( us32_n711 ) );
  NAND4_X1 us32_U94 (.A4( us32_n535 ) , .A3( us32_n536 ) , .A2( us32_n537 ) , .A1( us32_n538 ) , .ZN( us32_n622 ) );
  NOR4_X1 us32_U95 (.A4( us32_n526 ) , .A2( us32_n527 ) , .A1( us32_n528 ) , .ZN( us32_n538 ) , .A3( us32_n701 ) );
  NOR4_X1 us32_U96 (.A1( us32_n531 ) , .ZN( us32_n536 ) , .A2( us32_n654 ) , .A4( us32_n668 ) , .A3( us32_n765 ) );
  NOR4_X1 us32_U97 (.A4( us32_n529 ) , .A3( us32_n530 ) , .ZN( us32_n537 ) , .A2( us32_n684 ) , .A1( us32_n794 ) );
  NAND4_X1 us32_U98 (.A4( us32_n479 ) , .A3( us32_n480 ) , .A2( us32_n481 ) , .A1( us32_n482 ) , .ZN( us32_n694 ) );
  NOR3_X1 us32_U99 (.ZN( us32_n480 ) , .A2( us32_n508 ) , .A3( us32_n601 ) , .A1( us32_n610 ) );
endmodule

