module aes_aes_die_12 ( sa01_0, sa01_1, sa01_6, sa01_7, sa11_0, sa11_1, sa11_2, sa11_3, sa11_4, 
       sa11_5, sa11_6, sa11_7, us01_n439, us01_n445, us01_n446, us01_n447, us01_n449, us01_n450, 
       us01_n453, us01_n459, us01_n463, us01_n470, us01_n784, us01_n815, sa01_sr_0, sa01_sr_1, sa01_sr_2, sa01_sr_3, sa01_sr_4, sa01_sr_5, sa01_sr_6, sa01_sr_7, sa10_sr_0, 
        sa10_sr_1, sa10_sr_2, sa10_sr_3, sa10_sr_4, sa10_sr_5, sa10_sr_6, sa10_sr_7, us01_n469, us01_n847 );
  input sa01_0, sa01_1, sa01_6, sa01_7, sa11_0, sa11_1, sa11_2, sa11_3, sa11_4, 
        sa11_5, sa11_6, sa11_7, us01_n439, us01_n445, us01_n446, us01_n447, us01_n449, us01_n450, 
        us01_n453, us01_n459, us01_n463, us01_n470, us01_n784, us01_n815;
  output sa01_sr_0, sa01_sr_1, sa01_sr_2, sa01_sr_3, sa01_sr_4, sa01_sr_5, sa01_sr_6, sa01_sr_7, sa10_sr_0, 
        sa10_sr_1, sa10_sr_2, sa10_sr_3, sa10_sr_4, sa10_sr_5, sa10_sr_6, sa10_sr_7, us01_n469, us01_n847;
  wire us01_n438, us01_n440, us01_n441, us01_n442, us01_n443, us01_n444, us01_n448, us01_n451, us01_n452, 
       us01_n454, us01_n455, us01_n456, us01_n457, us01_n458, us01_n460, us01_n461, us01_n462, us01_n464, 
       us01_n465, us01_n466, us01_n467, us01_n468, us01_n471, us01_n472, us01_n473, us01_n474, us01_n475, 
       us01_n476, us01_n477, us01_n478, us01_n479, us01_n480, us01_n481, us01_n482, us01_n483, us01_n484, 
       us01_n485, us01_n486, us01_n487, us01_n488, us01_n489, us01_n490, us01_n491, us01_n492, us01_n493, 
       us01_n494, us01_n495, us01_n496, us01_n497, us01_n498, us01_n499, us01_n500, us01_n501, us01_n502, 
       us01_n503, us01_n504, us01_n505, us01_n506, us01_n507, us01_n508, us01_n509, us01_n510, us01_n511, 
       us01_n512, us01_n513, us01_n514, us01_n515, us01_n516, us01_n517, us01_n518, us01_n519, us01_n520, 
       us01_n521, us01_n522, us01_n523, us01_n524, us01_n525, us01_n526, us01_n527, us01_n528, us01_n529, 
       us01_n530, us01_n531, us01_n532, us01_n533, us01_n534, us01_n535, us01_n536, us01_n537, us01_n538, 
       us01_n539, us01_n540, us01_n541, us01_n542, us01_n543, us01_n544, us01_n545, us01_n546, us01_n547, 
       us01_n548, us01_n549, us01_n550, us01_n551, us01_n552, us01_n553, us01_n554, us01_n555, us01_n556, 
       us01_n557, us01_n558, us01_n559, us01_n560, us01_n561, us01_n562, us01_n563, us01_n564, us01_n565, 
       us01_n566, us01_n567, us01_n568, us01_n569, us01_n570, us01_n571, us01_n572, us01_n573, us01_n574, 
       us01_n575, us01_n576, us01_n577, us01_n578, us01_n579, us01_n580, us01_n581, us01_n582, us01_n583, 
       us01_n584, us01_n585, us01_n586, us01_n587, us01_n588, us01_n589, us01_n590, us01_n591, us01_n592, 
       us01_n593, us01_n594, us01_n595, us01_n596, us01_n597, us01_n598, us01_n599, us01_n600, us01_n601, 
       us01_n602, us01_n603, us01_n604, us01_n605, us01_n606, us01_n607, us01_n608, us01_n609, us01_n610, 
       us01_n611, us01_n612, us01_n613, us01_n614, us01_n615, us01_n616, us01_n617, us01_n618, us01_n619, 
       us01_n620, us01_n621, us01_n622, us01_n623, us01_n624, us01_n625, us01_n626, us01_n627, us01_n628, 
       us01_n629, us01_n630, us01_n631, us01_n632, us01_n633, us01_n634, us01_n635, us01_n636, us01_n637, 
       us01_n638, us01_n639, us01_n640, us01_n641, us01_n642, us01_n643, us01_n644, us01_n645, us01_n646, 
       us01_n647, us01_n648, us01_n649, us01_n650, us01_n651, us01_n652, us01_n653, us01_n654, us01_n655, 
       us01_n656, us01_n657, us01_n658, us01_n659, us01_n660, us01_n661, us01_n662, us01_n663, us01_n664, 
       us01_n665, us01_n666, us01_n667, us01_n668, us01_n669, us01_n670, us01_n671, us01_n672, us01_n673, 
       us01_n674, us01_n675, us01_n676, us01_n677, us01_n678, us01_n679, us01_n680, us01_n681, us01_n682, 
       us01_n683, us01_n684, us01_n685, us01_n686, us01_n687, us01_n688, us01_n689, us01_n690, us01_n691, 
       us01_n692, us01_n693, us01_n694, us01_n695, us01_n696, us01_n697, us01_n698, us01_n699, us01_n700, 
       us01_n701, us01_n702, us01_n703, us01_n704, us01_n705, us01_n706, us01_n707, us01_n708, us01_n709, 
       us01_n710, us01_n711, us01_n712, us01_n713, us01_n714, us01_n715, us01_n716, us01_n717, us01_n718, 
       us01_n719, us01_n720, us01_n721, us01_n722, us01_n723, us01_n724, us01_n725, us01_n726, us01_n727, 
       us01_n728, us01_n729, us01_n730, us01_n731, us01_n732, us01_n733, us01_n734, us01_n735, us01_n736, 
       us01_n737, us01_n738, us01_n739, us01_n740, us01_n741, us01_n742, us01_n743, us01_n744, us01_n745, 
       us01_n746, us01_n747, us01_n748, us01_n749, us01_n750, us01_n751, us01_n752, us01_n753, us01_n754, 
       us01_n755, us01_n756, us01_n757, us01_n758, us01_n759, us01_n760, us01_n761, us01_n762, us01_n763, 
       us01_n764, us01_n765, us01_n766, us01_n767, us01_n768, us01_n769, us01_n770, us01_n771, us01_n772, 
       us01_n773, us01_n774, us01_n775, us01_n776, us01_n777, us01_n778, us01_n779, us01_n780, us01_n781, 
       us01_n782, us01_n783, us01_n785, us01_n786, us01_n787, us01_n788, us01_n789, us01_n790, us01_n791, 
       us01_n792, us01_n793, us01_n794, us01_n795, us01_n796, us01_n797, us01_n798, us01_n799, us01_n800, 
       us01_n801, us01_n802, us01_n803, us01_n804, us01_n805, us01_n806, us01_n807, us01_n808, us01_n809, 
       us01_n810, us01_n811, us01_n812, us01_n813, us01_n814, us01_n816, us01_n817, us01_n818, us01_n819, 
       us01_n820, us01_n821, us01_n822, us01_n823, us01_n824, us01_n825, us01_n828, us01_n829, us01_n830, 
       us01_n831, us01_n832, us01_n833, us01_n834, us01_n835, us01_n836, us01_n837, us01_n838, us01_n839, 
       us01_n840, us01_n841, us01_n842, us01_n843, us01_n844, us01_n848, us01_n849, us01_n850, us01_n851, 
       us01_n852, us01_n853, us01_n854, us01_n855, us01_n857, us01_n858, us01_n859, us01_n860, us01_n861, 
       us01_n862, us01_n863, us01_n864, us01_n865, us01_n866, us01_n867, us01_n868, us01_n869, us01_n870, 
       us01_n871, us01_n872, us01_n873, us01_n874, us11_n438, us11_n439, us11_n440, us11_n441, us11_n442, 
       us11_n443, us11_n444, us11_n445, us11_n446, us11_n447, us11_n448, us11_n449, us11_n450, us11_n451, 
       us11_n452, us11_n453, us11_n454, us11_n455, us11_n456, us11_n457, us11_n458, us11_n459, us11_n460, 
       us11_n461, us11_n462, us11_n463, us11_n464, us11_n465, us11_n466, us11_n467, us11_n468, us11_n469, 
       us11_n470, us11_n471, us11_n472, us11_n473, us11_n474, us11_n475, us11_n476, us11_n477, us11_n478, 
       us11_n479, us11_n480, us11_n481, us11_n482, us11_n483, us11_n484, us11_n485, us11_n486, us11_n487, 
       us11_n488, us11_n489, us11_n490, us11_n491, us11_n492, us11_n493, us11_n494, us11_n495, us11_n496, 
       us11_n497, us11_n498, us11_n499, us11_n500, us11_n501, us11_n502, us11_n503, us11_n504, us11_n505, 
       us11_n506, us11_n507, us11_n508, us11_n509, us11_n510, us11_n511, us11_n512, us11_n513, us11_n514, 
       us11_n515, us11_n516, us11_n517, us11_n518, us11_n519, us11_n520, us11_n521, us11_n522, us11_n523, 
       us11_n524, us11_n525, us11_n526, us11_n527, us11_n528, us11_n529, us11_n530, us11_n531, us11_n532, 
       us11_n533, us11_n534, us11_n535, us11_n536, us11_n537, us11_n538, us11_n539, us11_n540, us11_n541, 
       us11_n542, us11_n543, us11_n544, us11_n545, us11_n546, us11_n547, us11_n548, us11_n549, us11_n550, 
       us11_n551, us11_n552, us11_n553, us11_n554, us11_n555, us11_n556, us11_n557, us11_n558, us11_n559, 
       us11_n560, us11_n561, us11_n562, us11_n563, us11_n564, us11_n565, us11_n566, us11_n567, us11_n568, 
       us11_n569, us11_n570, us11_n571, us11_n572, us11_n573, us11_n574, us11_n575, us11_n576, us11_n577, 
       us11_n578, us11_n579, us11_n580, us11_n581, us11_n582, us11_n583, us11_n584, us11_n585, us11_n586, 
       us11_n587, us11_n588, us11_n589, us11_n590, us11_n591, us11_n592, us11_n593, us11_n594, us11_n595, 
       us11_n596, us11_n597, us11_n598, us11_n599, us11_n600, us11_n601, us11_n602, us11_n603, us11_n604, 
       us11_n605, us11_n606, us11_n607, us11_n608, us11_n609, us11_n610, us11_n611, us11_n612, us11_n613, 
       us11_n614, us11_n615, us11_n616, us11_n617, us11_n618, us11_n619, us11_n620, us11_n621, us11_n622, 
       us11_n623, us11_n624, us11_n625, us11_n626, us11_n627, us11_n628, us11_n629, us11_n630, us11_n631, 
       us11_n632, us11_n633, us11_n634, us11_n635, us11_n636, us11_n637, us11_n638, us11_n639, us11_n640, 
       us11_n641, us11_n642, us11_n643, us11_n644, us11_n645, us11_n646, us11_n647, us11_n648, us11_n649, 
       us11_n650, us11_n651, us11_n652, us11_n653, us11_n654, us11_n655, us11_n656, us11_n657, us11_n658, 
       us11_n659, us11_n660, us11_n661, us11_n662, us11_n663, us11_n664, us11_n665, us11_n666, us11_n667, 
       us11_n668, us11_n669, us11_n670, us11_n671, us11_n672, us11_n673, us11_n674, us11_n675, us11_n676, 
       us11_n677, us11_n678, us11_n679, us11_n680, us11_n681, us11_n682, us11_n683, us11_n684, us11_n685, 
       us11_n686, us11_n687, us11_n688, us11_n689, us11_n690, us11_n691, us11_n692, us11_n693, us11_n694, 
       us11_n695, us11_n696, us11_n697, us11_n698, us11_n699, us11_n700, us11_n701, us11_n702, us11_n703, 
       us11_n704, us11_n705, us11_n706, us11_n707, us11_n708, us11_n709, us11_n710, us11_n711, us11_n712, 
       us11_n713, us11_n714, us11_n715, us11_n716, us11_n717, us11_n718, us11_n719, us11_n720, us11_n721, 
       us11_n722, us11_n723, us11_n724, us11_n725, us11_n726, us11_n727, us11_n728, us11_n729, us11_n730, 
       us11_n731, us11_n732, us11_n733, us11_n734, us11_n735, us11_n736, us11_n737, us11_n738, us11_n739, 
       us11_n740, us11_n741, us11_n742, us11_n743, us11_n744, us11_n745, us11_n746, us11_n747, us11_n748, 
       us11_n749, us11_n750, us11_n751, us11_n752, us11_n753, us11_n754, us11_n755, us11_n756, us11_n757, 
       us11_n758, us11_n759, us11_n760, us11_n761, us11_n762, us11_n763, us11_n764, us11_n765, us11_n766, 
       us11_n767, us11_n768, us11_n769, us11_n770, us11_n771, us11_n772, us11_n773, us11_n774, us11_n775, 
       us11_n776, us11_n777, us11_n778, us11_n779, us11_n780, us11_n781, us11_n782, us11_n783, us11_n784, 
       us11_n785, us11_n786, us11_n787, us11_n788, us11_n789, us11_n790, us11_n791, us11_n792, us11_n793, 
       us11_n794, us11_n795, us11_n796, us11_n797, us11_n798, us11_n799, us11_n800, us11_n801, us11_n802, 
       us11_n803, us11_n804, us11_n805, us11_n806, us11_n807, us11_n808, us11_n809, us11_n810, us11_n811, 
       us11_n812, us11_n813, us11_n814, us11_n815, us11_n816, us11_n817, us11_n818, us11_n819, us11_n820, 
       us11_n821, us11_n822, us11_n823, us11_n824, us11_n825, us11_n826, us11_n827, us11_n828, us11_n829, 
       us11_n830, us11_n831, us11_n832, us11_n833, us11_n834, us11_n835, us11_n836, us11_n837, us11_n838, 
       us11_n839, us11_n840, us11_n841, us11_n842, us11_n843, us11_n844, us11_n845, us11_n846, us11_n847, 
       us11_n848, us11_n849, us11_n850, us11_n851, us11_n852, us11_n853, us11_n854, us11_n855, us11_n856, 
       us11_n857, us11_n858, us11_n859, us11_n860, us11_n861, us11_n862, us11_n863, us11_n864, us11_n865, 
       us11_n866, us11_n867, us11_n868, us11_n869, us11_n870, us11_n871, us11_n872, us11_n873, us11_n874, 
       us11_n875,  us11_n876;
  NOR2_X1 us01_U10 (.ZN( us01_n573 ) , .A1( us01_n620 ) , .A2( us01_n743 ) );
  AOI211_X1 us01_U100 (.B( us01_n537 ) , .A( us01_n538 ) , .ZN( us01_n549 ) , .C2( us01_n837 ) , .C1( us01_n849 ) );
  NOR4_X1 us01_U101 (.A4( us01_n542 ) , .A3( us01_n543 ) , .A2( us01_n544 ) , .A1( us01_n545 ) , .ZN( us01_n546 ) );
  NOR4_X1 us01_U102 (.A4( us01_n607 ) , .A3( us01_n608 ) , .A2( us01_n609 ) , .A1( us01_n610 ) , .ZN( us01_n617 ) );
  NOR4_X1 us01_U103 (.ZN( us01_n618 ) , .A1( us01_n654 ) , .A3( us01_n664 ) , .A4( us01_n680 ) , .A2( us01_n764 ) );
  NOR4_X1 us01_U104 (.A4( us01_n612 ) , .A3( us01_n613 ) , .A2( us01_n614 ) , .A1( us01_n615 ) , .ZN( us01_n616 ) );
  NOR2_X1 us01_U105 (.ZN( us01_n684 ) , .A1( us01_n829 ) , .A2( us01_n830 ) );
  NAND4_X1 us01_U106 (.A4( us01_n471 ) , .A3( us01_n472 ) , .A2( us01_n473 ) , .A1( us01_n474 ) , .ZN( us01_n676 ) );
  NOR4_X1 us01_U107 (.A4( us01_n468 ) , .ZN( us01_n474 ) , .A3( us01_n554 ) , .A1( us01_n733 ) , .A2( us01_n753 ) );
  NOR4_X1 us01_U108 (.ZN( us01_n473 ) , .A1( us01_n529 ) , .A3( us01_n566 ) , .A4( us01_n598 ) , .A2( us01_n640 ) );
  NOR4_X1 us01_U109 (.ZN( us01_n472 ) , .A1( us01_n504 ) , .A3( us01_n542 ) , .A2( us01_n581 ) , .A4( us01_n714 ) );
  NOR2_X1 us01_U11 (.ZN( us01_n493 ) , .A1( us01_n676 ) , .A2( us01_n692 ) );
  NAND4_X1 us01_U110 (.A4( us01_n689 ) , .A3( us01_n690 ) , .A1( us01_n691 ) , .ZN( us01_n774 ) , .A2( us01_n870 ) );
  INV_X1 us01_U111 (.A( us01_n677 ) , .ZN( us01_n870 ) );
  AOI221_X1 us01_U112 (.A( us01_n679 ) , .ZN( us01_n690 ) , .B2( us01_n838 ) , .C1( us01_n840 ) , .C2( us01_n860 ) , .B1( us01_n863 ) );
  NOR4_X1 us01_U113 (.A4( us01_n685 ) , .A3( us01_n686 ) , .A2( us01_n687 ) , .A1( us01_n688 ) , .ZN( us01_n689 ) );
  NOR2_X1 us01_U114 (.ZN( us01_n731 ) , .A2( us01_n830 ) , .A1( us01_n843 ) );
  NAND4_X1 us01_U115 (.A4( us01_n717 ) , .A3( us01_n718 ) , .A2( us01_n719 ) , .ZN( us01_n739 ) , .A1( us01_n855 ) );
  AOI221_X1 us01_U116 (.A( us01_n708 ) , .ZN( us01_n719 ) , .C2( us01_n842 ) , .B2( us01_n843 ) , .C1( us01_n859 ) , .B1( us01_n860 ) );
  INV_X1 us01_U117 (.A( us01_n707 ) , .ZN( us01_n855 ) );
  NOR4_X1 us01_U118 (.A4( us01_n713 ) , .A3( us01_n714 ) , .A2( us01_n715 ) , .A1( us01_n716 ) , .ZN( us01_n717 ) );
  NOR2_X1 us01_U119 (.ZN( us01_n645 ) , .A1( us01_n852 ) , .A2( us01_n866 ) );
  NOR2_X1 us01_U12 (.A1( us01_n676 ) , .ZN( us01_n691 ) , .A2( us01_n805 ) );
  NAND4_X1 us01_U120 (.A4( us01_n571 ) , .A3( us01_n572 ) , .A1( us01_n573 ) , .ZN( us01_n721 ) , .A2( us01_n872 ) );
  AOI221_X1 us01_U121 (.A( us01_n562 ) , .C2( us01_n563 ) , .ZN( us01_n572 ) , .B2( us01_n843 ) , .B1( us01_n850 ) , .C1( us01_n851 ) );
  NOR4_X1 us01_U122 (.A4( us01_n567 ) , .A3( us01_n568 ) , .A2( us01_n569 ) , .A1( us01_n570 ) , .ZN( us01_n571 ) );
  INV_X1 us01_U123 (.A( us01_n605 ) , .ZN( us01_n872 ) );
  NAND4_X1 us01_U124 (.A4( us01_n491 ) , .A3( us01_n492 ) , .A1( us01_n493 ) , .ZN( us01_n800 ) , .A2( us01_n865 ) );
  AOI221_X1 us01_U125 (.A( us01_n487 ) , .ZN( us01_n492 ) , .B2( us01_n834 ) , .C2( us01_n839 ) , .C1( us01_n849 ) , .B1( us01_n858 ) );
  INV_X1 us01_U126 (.A( us01_n776 ) , .ZN( us01_n865 ) );
  NOR4_X1 us01_U127 (.A2( us01_n489 ) , .A1( us01_n490 ) , .ZN( us01_n491 ) , .A3( us01_n578 ) , .A4( us01_n610 ) );
  NOR4_X1 us01_U128 (.A3( us01_n753 ) , .A2( us01_n754 ) , .A1( us01_n755 ) , .ZN( us01_n756 ) , .A4( us01_n867 ) );
  AOI211_X1 us01_U129 (.B( us01_n743 ) , .A( us01_n744 ) , .ZN( us01_n757 ) , .C1( us01_n830 ) , .C2( us01_n851 ) );
  NOR3_X1 us01_U13 (.ZN( us01_n502 ) , .A2( us01_n677 ) , .A3( us01_n775 ) , .A1( us01_n874 ) );
  NOR3_X1 us01_U130 (.A3( us01_n739 ) , .A2( us01_n740 ) , .A1( us01_n741 ) , .ZN( us01_n758 ) );
  NOR4_X1 us01_U131 (.A4( us01_n732 ) , .A3( us01_n733 ) , .A2( us01_n734 ) , .A1( us01_n735 ) , .ZN( us01_n736 ) );
  AOI211_X1 us01_U132 (.B( us01_n723 ) , .A( us01_n724 ) , .ZN( us01_n737 ) , .C1( us01_n841 ) , .C2( us01_n853 ) );
  NOR3_X1 us01_U133 (.A3( us01_n720 ) , .A1( us01_n721 ) , .ZN( us01_n738 ) , .A2( us01_n739 ) );
  INV_X1 us01_U134 (.A( us01_n760 ) , .ZN( us01_n828 ) );
  NAND4_X1 us01_U135 (.ZN( sa01_sr_3 ) , .A4( us01_n702 ) , .A3( us01_n703 ) , .A2( us01_n704 ) , .A1( us01_n705 ) );
  NOR4_X1 us01_U136 (.A4( us01_n698 ) , .A3( us01_n699 ) , .A2( us01_n700 ) , .A1( us01_n701 ) , .ZN( us01_n702 ) );
  AOI211_X1 us01_U137 (.B( us01_n692 ) , .A( us01_n693 ) , .ZN( us01_n703 ) , .C2( us01_n829 ) , .C1( us01_n849 ) );
  NOR2_X1 us01_U138 (.ZN( us01_n705 ) , .A2( us01_n774 ) , .A1( us01_n798 ) );
  OR4_X1 us01_U139 (.A4( us01_n680 ) , .A3( us01_n681 ) , .A2( us01_n682 ) , .A1( us01_n683 ) , .ZN( us01_n688 ) );
  INV_X1 us01_U14 (.A( us01_n704 ) , .ZN( us01_n874 ) );
  OR4_X1 us01_U140 (.ZN( us01_n464 ) , .A4( us01_n516 ) , .A3( us01_n527 ) , .A2( us01_n576 ) , .A1( us01_n710 ) );
  OR4_X1 us01_U141 (.A4( us01_n564 ) , .A3( us01_n565 ) , .A2( us01_n566 ) , .ZN( us01_n570 ) , .A1( us01_n663 ) );
  OR4_X1 us01_U142 (.A4( us01_n516 ) , .A2( us01_n517 ) , .A1( us01_n518 ) , .ZN( us01_n520 ) , .A3( us01_n819 ) );
  OR4_X1 us01_U143 (.ZN( us01_n490 ) , .A4( us01_n532 ) , .A2( us01_n545 ) , .A1( us01_n557 ) , .A3( us01_n630 ) );
  OR4_X1 us01_U144 (.A4( us01_n578 ) , .A3( us01_n579 ) , .A2( us01_n580 ) , .A1( us01_n581 ) , .ZN( us01_n582 ) );
  INV_X1 us01_U145 (.A( us01_n695 ) , .ZN( us01_n836 ) );
  NAND2_X1 us01_U146 (.ZN( us01_n611 ) , .A2( us01_n835 ) , .A1( us01_n871 ) );
  OR3_X1 us01_U147 (.A3( us01_n504 ) , .A2( us01_n505 ) , .A1( us01_n506 ) , .ZN( us01_n509 ) );
  AOI221_X1 us01_U148 (.A( us01_n711 ) , .B2( us01_n712 ) , .ZN( us01_n718 ) , .C1( us01_n830 ) , .B1( us01_n837 ) , .C2( us01_n861 ) );
  OR2_X1 us01_U149 (.A2( us01_n709 ) , .A1( us01_n710 ) , .ZN( us01_n711 ) );
  INV_X1 us01_U15 (.A( us01_n678 ) , .ZN( us01_n838 ) );
  INV_X1 us01_U150 (.A( us01_n461 ) , .ZN( us01_n862 ) );
  OAI21_X1 us01_U151 (.ZN( us01_n461 ) , .B1( us01_n807 ) , .A( us01_n832 ) , .B2( us01_n849 ) );
  INV_X1 us01_U152 (.A( us01_n752 ) , .ZN( us01_n867 ) );
  OAI21_X1 us01_U153 (.B1( us01_n751 ) , .ZN( us01_n752 ) , .A( us01_n843 ) , .B2( us01_n866 ) );
  INV_X1 us01_U154 (.A( us01_n670 ) , .ZN( us01_n857 ) );
  AOI21_X1 us01_U155 (.A( us01_n668 ) , .B1( us01_n669 ) , .ZN( us01_n670 ) , .B2( us01_n854 ) );
  AOI222_X1 us01_U156 (.ZN( us01_n658 ) , .A2( us01_n837 ) , .B1( us01_n839 ) , .C2( us01_n843 ) , .A1( us01_n858 ) , .C1( us01_n861 ) , .B2( us01_n868 ) );
  INV_X1 us01_U157 (.A( us01_n645 ) , .ZN( us01_n868 ) );
  OAI22_X1 us01_U158 (.ZN( us01_n481 ) , .A1( us01_n706 ) , .B2( us01_n783 ) , .A2( us01_n804 ) , .B1( us01_n810 ) );
  OAI22_X1 us01_U159 (.ZN( us01_n635 ) , .A1( us01_n697 ) , .B2( us01_n726 ) , .A2( us01_n760 ) , .B1( us01_n814 ) );
  NOR4_X1 us01_U16 (.A4( us01_n443 ) , .A3( us01_n444 ) , .A2( us01_n514 ) , .A1( us01_n539 ) , .ZN( us01_n704 ) );
  OAI222_X1 us01_U160 (.ZN( us01_n503 ) , .C2( us01_n623 ) , .B2( us01_n645 ) , .B1( us01_n745 ) , .A2( us01_n746 ) , .C1( us01_n803 ) , .A1( us01_n804 ) );
  OAI222_X1 us01_U161 (.B2( us01_n745 ) , .B1( us01_n746 ) , .A2( us01_n747 ) , .ZN( us01_n755 ) , .C2( us01_n803 ) , .C1( us01_n812 ) , .A1( us01_n815 ) );
  OAI222_X1 us01_U162 (.B2( us01_n706 ) , .ZN( us01_n707 ) , .C2( us01_n722 ) , .B1( us01_n745 ) , .A1( us01_n804 ) , .C1( us01_n812 ) , .A2( us01_n813 ) );
  AOI22_X1 us01_U163 (.ZN( us01_n694 ) , .A1( us01_n828 ) , .B2( us01_n841 ) , .A2( us01_n863 ) , .B1( us01_n866 ) );
  AOI22_X1 us01_U164 (.A2( us01_n780 ) , .ZN( us01_n781 ) , .B2( us01_n829 ) , .A1( us01_n832 ) , .B1( us01_n861 ) );
  INV_X1 us01_U165 (.A( us01_n728 ) , .ZN( us01_n837 ) );
  AOI221_X1 us01_U166 (.A( us01_n762 ) , .ZN( us01_n772 ) , .C2( us01_n808 ) , .B2( us01_n833 ) , .C1( us01_n853 ) , .B1( us01_n864 ) );
  AOI21_X1 us01_U167 (.B2( us01_n761 ) , .ZN( us01_n762 ) , .A( us01_n786 ) , .B1( us01_n790 ) );
  INV_X1 us01_U168 (.A( us01_n759 ) , .ZN( us01_n833 ) );
  INV_X1 us01_U169 (.A( us01_n788 ) , .ZN( us01_n830 ) );
  OR3_X1 us01_U17 (.ZN( us01_n444 ) , .A1( us01_n526 ) , .A3( us01_n575 ) , .A2( us01_n873 ) );
  OAI221_X1 us01_U170 (.A( us01_n725 ) , .C2( us01_n726 ) , .B2( us01_n727 ) , .B1( us01_n728 ) , .ZN( us01_n735 ) , .C1( us01_n815 ) );
  AOI22_X1 us01_U171 (.ZN( us01_n725 ) , .B1( us01_n830 ) , .A2( us01_n836 ) , .A1( us01_n861 ) , .B2( us01_n864 ) );
  NAND2_X1 us01_U172 (.A1( us01_n449 ) , .A2( us01_n451 ) , .ZN( us01_n760 ) );
  OAI22_X1 us01_U173 (.ZN( us01_n622 ) , .B1( us01_n667 ) , .B2( us01_n745 ) , .A1( us01_n813 ) , .A2( us01_n814 ) );
  OAI22_X1 us01_U174 (.A1( us01_n722 ) , .ZN( us01_n724 ) , .B2( us01_n748 ) , .B1( us01_n810 ) , .A2( us01_n814 ) );
  OAI22_X1 us01_U175 (.ZN( us01_n487 ) , .A1( us01_n722 ) , .B2( us01_n726 ) , .B1( us01_n728 ) , .A2( us01_n777 ) );
  OAI22_X1 us01_U176 (.B2( us01_n777 ) , .B1( us01_n778 ) , .ZN( us01_n779 ) , .A2( us01_n812 ) , .A1( us01_n813 ) );
  OAI22_X1 us01_U177 (.B2( us01_n748 ) , .B1( us01_n749 ) , .A1( us01_n750 ) , .ZN( us01_n754 ) , .A2( us01_n804 ) );
  NOR3_X1 us01_U178 (.ZN( us01_n750 ) , .A2( us01_n851 ) , .A1( us01_n861 ) , .A3( us01_n863 ) );
  NOR2_X1 us01_U179 (.ZN( us01_n749 ) , .A2( us01_n850 ) , .A1( us01_n858 ) );
  OR4_X1 us01_U18 (.A4( us01_n440 ) , .A2( us01_n441 ) , .A1( us01_n442 ) , .ZN( us01_n443 ) , .A3( us01_n551 ) );
  INV_X1 us01_U180 (.A( us01_n803 ) , .ZN( us01_n858 ) );
  OAI22_X1 us01_U181 (.B2( us01_n742 ) , .ZN( us01_n744 ) , .A2( us01_n760 ) , .B1( us01_n778 ) , .A1( us01_n790 ) );
  OAI22_X1 us01_U182 (.ZN( us01_n494 ) , .A2( us01_n742 ) , .A1( us01_n778 ) , .B1( us01_n789 ) , .B2( us01_n804 ) );
  OAI22_X1 us01_U183 (.B2( us01_n801 ) , .B1( us01_n802 ) , .A2( us01_n803 ) , .A1( us01_n804 ) , .ZN( us01_n806 ) );
  OAI22_X1 us01_U184 (.ZN( us01_n693 ) , .A2( us01_n728 ) , .A1( us01_n778 ) , .B1( us01_n789 ) , .B2( us01_n815 ) );
  NOR2_X1 us01_U185 (.ZN( us01_n713 ) , .A1( us01_n803 ) , .A2( us01_n815 ) );
  NOR2_X1 us01_U186 (.A1( us01_n697 ) , .ZN( us01_n766 ) , .A2( us01_n811 ) );
  INV_X1 us01_U187 (.A( us01_n786 ) , .ZN( us01_n843 ) );
  NOR2_X1 us01_U188 (.ZN( us01_n539 ) , .A2( us01_n695 ) , .A1( us01_n697 ) );
  INV_X1 us01_U189 (.A( us01_n742 ) , .ZN( us01_n835 ) );
  INV_X1 us01_U19 (.A( us01_n611 ) , .ZN( us01_n873 ) );
  INV_X1 us01_U190 (.A( us01_n814 ) , .ZN( us01_n829 ) );
  INV_X1 us01_U191 (.A( us01_n812 ) , .ZN( us01_n831 ) );
  OAI22_X1 us01_U192 (.B1( us01_n488 ) , .ZN( us01_n489 ) , .A1( us01_n684 ) , .A2( us01_n761 ) , .B2( us01_n815 ) );
  NOR3_X1 us01_U193 (.ZN( us01_n488 ) , .A1( us01_n780 ) , .A2( us01_n848 ) , .A3( us01_n861 ) );
  NOR2_X1 us01_U194 (.A2( us01_n742 ) , .ZN( us01_n753 ) , .A1( us01_n803 ) );
  NOR2_X1 us01_U195 (.ZN( us01_n733 ) , .A2( us01_n801 ) , .A1( us01_n803 ) );
  INV_X1 us01_U196 (.A( us01_n790 ) , .ZN( us01_n849 ) );
  NOR2_X1 us01_U197 (.A2( us01_n742 ) , .ZN( us01_n767 ) , .A1( us01_n810 ) );
  NOR2_X1 us01_U198 (.ZN( us01_n664 ) , .A1( us01_n726 ) , .A2( us01_n801 ) );
  OAI22_X1 us01_U199 (.ZN( us01_n708 ) , .A2( us01_n726 ) , .B2( us01_n727 ) , .A1( us01_n742 ) , .B1( us01_n811 ) );
  AOI222_X1 us01_U20 (.ZN( us01_n561 ) , .B1( us01_n828 ) , .C1( us01_n839 ) , .A2( us01_n841 ) , .A1( us01_n852 ) , .B2( us01_n861 ) , .C2( us01_n871 ) );
  NOR2_X1 us01_U200 (.ZN( us01_n650 ) , .A1( us01_n667 ) , .A2( us01_n812 ) );
  NOR2_X1 us01_U201 (.ZN( us01_n592 ) , .A2( us01_n695 ) , .A1( us01_n726 ) );
  NOR2_X1 us01_U202 (.A1( us01_n667 ) , .ZN( us01_n671 ) , .A2( us01_n742 ) );
  NOR2_X1 us01_U203 (.ZN( us01_n600 ) , .A1( us01_n667 ) , .A2( us01_n801 ) );
  NOR2_X1 us01_U204 (.A1( us01_n667 ) , .ZN( us01_n686 ) , .A2( us01_n814 ) );
  NOR2_X1 us01_U205 (.ZN( us01_n568 ) , .A1( us01_n726 ) , .A2( us01_n804 ) );
  NOR2_X1 us01_U206 (.A1( us01_n667 ) , .ZN( us01_n764 ) , .A2( us01_n811 ) );
  NOR2_X1 us01_U207 (.ZN( us01_n525 ) , .A1( us01_n667 ) , .A2( us01_n777 ) );
  NOR2_X1 us01_U208 (.ZN( us01_n652 ) , .A1( us01_n726 ) , .A2( us01_n811 ) );
  NOR2_X1 us01_U209 (.ZN( us01_n505 ) , .A1( us01_n810 ) , .A2( us01_n815 ) );
  NOR4_X1 us01_U21 (.ZN( us01_n471 ) , .A2( us01_n519 ) , .A4( us01_n592 ) , .A1( us01_n607 ) , .A3( us01_n627 ) );
  NOR2_X1 us01_U210 (.ZN( us01_n659 ) , .A1( us01_n727 ) , .A2( us01_n788 ) );
  NOR2_X1 us01_U211 (.ZN( us01_n544 ) , .A2( us01_n778 ) , .A1( us01_n812 ) );
  NOR2_X1 us01_U212 (.ZN( us01_n575 ) , .A2( us01_n697 ) , .A1( us01_n812 ) );
  NOR2_X1 us01_U213 (.ZN( us01_n507 ) , .A1( us01_n727 ) , .A2( us01_n777 ) );
  NOR2_X1 us01_U214 (.ZN( us01_n716 ) , .A2( us01_n722 ) , .A1( us01_n742 ) );
  INV_X1 us01_U215 (.A( us01_n748 ) , .ZN( us01_n840 ) );
  NOR2_X1 us01_U216 (.ZN( us01_n530 ) , .A2( us01_n747 ) , .A1( us01_n748 ) );
  NOR2_X1 us01_U217 (.ZN( us01_n660 ) , .A2( us01_n695 ) , .A1( us01_n727 ) );
  NOR2_X1 us01_U218 (.ZN( us01_n613 ) , .A1( us01_n783 ) , .A2( us01_n813 ) );
  NOR2_X1 us01_U219 (.ZN( us01_n627 ) , .A2( us01_n726 ) , .A1( us01_n783 ) );
  NOR4_X1 us01_U22 (.ZN( us01_n477 ) , .A1( us01_n518 ) , .A4( us01_n555 ) , .A3( us01_n580 ) , .A2( us01_n628 ) );
  NOR2_X1 us01_U220 (.ZN( us01_n609 ) , .A2( us01_n778 ) , .A1( us01_n804 ) );
  NOR2_X1 us01_U221 (.ZN( us01_n661 ) , .A1( us01_n727 ) , .A2( us01_n783 ) );
  NOR2_X1 us01_U222 (.ZN( us01_n626 ) , .A2( us01_n667 ) , .A1( us01_n783 ) );
  NOR2_X1 us01_U223 (.ZN( us01_n599 ) , .A2( us01_n778 ) , .A1( us01_n801 ) );
  INV_X1 us01_U224 (.A( us01_n745 ) , .ZN( us01_n832 ) );
  NOR2_X1 us01_U225 (.ZN( us01_n554 ) , .A1( us01_n760 ) , .A2( us01_n803 ) );
  NOR2_X1 us01_U226 (.ZN( us01_n529 ) , .A2( us01_n778 ) , .A1( us01_n814 ) );
  NOR2_X1 us01_U227 (.ZN( us01_n526 ) , .A2( us01_n722 ) , .A1( us01_n801 ) );
  NOR2_X1 us01_U228 (.A2( us01_n706 ) , .A1( us01_n748 ) , .ZN( us01_n769 ) );
  NOR2_X1 us01_U229 (.ZN( us01_n597 ) , .A2( us01_n789 ) , .A1( us01_n814 ) );
  NOR4_X1 us01_U23 (.ZN( us01_n454 ) , .A2( us01_n515 ) , .A1( us01_n541 ) , .A3( us01_n577 ) , .A4( us01_n613 ) );
  NOR2_X1 us01_U230 (.ZN( us01_n555 ) , .A1( us01_n790 ) , .A2( us01_n812 ) );
  NOR2_X1 us01_U231 (.ZN( us01_n542 ) , .A2( us01_n783 ) , .A1( us01_n790 ) );
  NOR2_X1 us01_U232 (.A2( us01_n695 ) , .ZN( us01_n714 ) , .A1( us01_n790 ) );
  NOR2_X1 us01_U233 (.ZN( us01_n665 ) , .A1( us01_n748 ) , .A2( us01_n813 ) );
  NOR2_X1 us01_U234 (.ZN( us01_n543 ) , .A1( us01_n747 ) , .A2( us01_n812 ) );
  NOR2_X1 us01_U235 (.ZN( us01_n553 ) , .A1( us01_n748 ) , .A2( us01_n789 ) );
  NOR2_X1 us01_U236 (.ZN( us01_n506 ) , .A2( us01_n778 ) , .A1( us01_n783 ) );
  NOR2_X1 us01_U237 (.ZN( us01_n541 ) , .A2( us01_n706 ) , .A1( us01_n783 ) );
  NOR2_X1 us01_U238 (.ZN( us01_n514 ) , .A1( us01_n706 ) , .A2( us01_n742 ) );
  NOR2_X1 us01_U239 (.ZN( us01_n662 ) , .A1( us01_n783 ) , .A2( us01_n789 ) );
  NOR4_X1 us01_U24 (.A4( us01_n530 ) , .A3( us01_n531 ) , .A2( us01_n532 ) , .ZN( us01_n533 ) , .A1( us01_n818 ) );
  NOR2_X1 us01_U240 (.ZN( us01_n556 ) , .A1( us01_n706 ) , .A2( us01_n814 ) );
  NOR2_X1 us01_U241 (.ZN( us01_n515 ) , .A1( us01_n706 ) , .A2( us01_n801 ) );
  NOR2_X1 us01_U242 (.ZN( us01_n612 ) , .A1( us01_n760 ) , .A2( us01_n810 ) );
  NOR2_X1 us01_U243 (.ZN( us01_n629 ) , .A1( us01_n722 ) , .A2( us01_n811 ) );
  NOR2_X1 us01_U244 (.A1( us01_n747 ) , .ZN( us01_n765 ) , .A2( us01_n801 ) );
  NOR2_X1 us01_U245 (.ZN( us01_n528 ) , .A2( us01_n742 ) , .A1( us01_n790 ) );
  INV_X1 us01_U246 (.A( us01_n804 ) , .ZN( us01_n839 ) );
  OAI22_X1 us01_U247 (.B1( us01_n438 ) , .ZN( us01_n442 ) , .A2( us01_n726 ) , .A1( us01_n742 ) , .B2( us01_n747 ) );
  NOR3_X1 us01_U248 (.ZN( us01_n438 ) , .A2( us01_n834 ) , .A3( us01_n835 ) , .A1( us01_n844 ) );
  INV_X1 us01_U249 (.A( us01_n726 ) , .ZN( us01_n850 ) );
  NOR4_X1 us01_U25 (.A4( us01_n539 ) , .A3( us01_n540 ) , .A2( us01_n541 ) , .ZN( us01_n548 ) , .A1( us01_n686 ) );
  NOR2_X1 us01_U250 (.ZN( us01_n519 ) , .A1( us01_n788 ) , .A2( us01_n810 ) );
  NOR2_X1 us01_U251 (.ZN( us01_n668 ) , .A1( us01_n788 ) , .A2( us01_n803 ) );
  AOI21_X1 us01_U252 (.ZN( us01_n550 ) , .B1( us01_n667 ) , .A( us01_n695 ) , .B2( us01_n803 ) );
  AOI21_X1 us01_U253 (.ZN( us01_n587 ) , .B2( us01_n697 ) , .B1( us01_n813 ) , .A( us01_n815 ) );
  NOR2_X1 us01_U254 (.ZN( us01_n504 ) , .A2( us01_n726 ) , .A1( us01_n760 ) );
  NOR2_X1 us01_U255 (.ZN( us01_n653 ) , .A1( us01_n788 ) , .A2( us01_n813 ) );
  INV_X1 us01_U256 (.A( us01_n801 ) , .ZN( us01_n841 ) );
  NOR2_X1 us01_U257 (.ZN( us01_n628 ) , .A1( us01_n745 ) , .A2( us01_n813 ) );
  NOR2_X1 us01_U258 (.ZN( us01_n545 ) , .A1( us01_n697 ) , .A2( us01_n742 ) );
  INV_X1 us01_U259 (.A( us01_n697 ) , .ZN( us01_n851 ) );
  NOR2_X1 us01_U26 (.ZN( us01_n678 ) , .A2( us01_n832 ) , .A1( us01_n837 ) );
  NOR2_X1 us01_U260 (.ZN( us01_n640 ) , .A2( us01_n786 ) , .A1( us01_n789 ) );
  AOI21_X1 us01_U261 (.ZN( us01_n648 ) , .A( us01_n777 ) , .B1( us01_n790 ) , .B2( us01_n803 ) );
  NOR2_X1 us01_U262 (.ZN( us01_n666 ) , .A2( us01_n706 ) , .A1( us01_n788 ) );
  NOR2_X1 us01_U263 (.A2( us01_n695 ) , .A1( us01_n778 ) , .ZN( us01_n818 ) );
  NOR2_X1 us01_U264 (.A1( us01_n695 ) , .ZN( us01_n768 ) , .A2( us01_n813 ) );
  AOI21_X1 us01_U265 (.ZN( us01_n624 ) , .B2( us01_n667 ) , .A( us01_n788 ) , .B1( us01_n789 ) );
  NOR2_X1 us01_U266 (.ZN( us01_n577 ) , .A2( us01_n706 ) , .A1( us01_n728 ) );
  INV_X1 us01_U267 (.A( us01_n761 ) , .ZN( us01_n864 ) );
  NOR2_X1 us01_U268 (.A2( us01_n706 ) , .A1( us01_n760 ) , .ZN( us01_n792 ) );
  NOR2_X1 us01_U269 (.ZN( us01_n607 ) , .A2( us01_n722 ) , .A1( us01_n815 ) );
  AOI222_X1 us01_U27 (.ZN( us01_n467 ) , .B1( us01_n830 ) , .A1( us01_n837 ) , .C1( us01_n840 ) , .C2( us01_n849 ) , .A2( us01_n853 ) , .B2( us01_n863 ) );
  NOR2_X1 us01_U270 (.ZN( us01_n531 ) , .A2( us01_n722 ) , .A1( us01_n728 ) );
  AOI21_X1 us01_U271 (.ZN( us01_n508 ) , .B2( us01_n667 ) , .A( us01_n728 ) , .B1( us01_n813 ) );
  AOI21_X1 us01_U272 (.ZN( us01_n537 ) , .B2( us01_n810 ) , .A( us01_n812 ) , .B1( us01_n813 ) );
  INV_X1 us01_U273 (.A( us01_n727 ) , .ZN( us01_n866 ) );
  NOR2_X1 us01_U274 (.ZN( us01_n540 ) , .A1( us01_n760 ) , .A2( us01_n789 ) );
  INV_X1 us01_U275 (.A( us01_n810 ) , .ZN( us01_n852 ) );
  AOI21_X1 us01_U276 (.B1( us01_n697 ) , .ZN( us01_n698 ) , .A( us01_n730 ) , .B2( us01_n761 ) );
  NOR2_X1 us01_U277 (.ZN( us01_n579 ) , .A1( us01_n667 ) , .A2( us01_n786 ) );
  AOI21_X1 us01_U278 (.ZN( us01_n589 ) , .B2( us01_n761 ) , .A( us01_n783 ) , .B1( us01_n810 ) );
  NOR2_X1 us01_U279 (.ZN( us01_n654 ) , .A1( us01_n745 ) , .A2( us01_n778 ) );
  NOR4_X1 us01_U28 (.A1( us01_n464 ) , .ZN( us01_n465 ) , .A4( us01_n540 ) , .A2( us01_n552 ) , .A3( us01_n612 ) );
  INV_X1 us01_U280 (.A( us01_n789 ) , .ZN( us01_n871 ) );
  AOI21_X1 us01_U281 (.B1( us01_n623 ) , .ZN( us01_n625 ) , .A( us01_n761 ) , .B2( us01_n812 ) );
  NOR2_X1 us01_U282 (.ZN( us01_n683 ) , .A1( us01_n727 ) , .A2( us01_n814 ) );
  AOI21_X1 us01_U283 (.A( us01_n813 ) , .B2( us01_n814 ) , .B1( us01_n815 ) , .ZN( us01_n816 ) );
  AOI21_X1 us01_U284 (.ZN( us01_n647 ) , .B1( us01_n727 ) , .B2( us01_n761 ) , .A( us01_n811 ) );
  AOI21_X1 us01_U285 (.A( us01_n810 ) , .B2( us01_n811 ) , .B1( us01_n812 ) , .ZN( us01_n817 ) );
  AOI21_X1 us01_U286 (.ZN( us01_n513 ) , .A( us01_n727 ) , .B1( us01_n748 ) , .B2( us01_n801 ) );
  AOI21_X1 us01_U287 (.ZN( us01_n497 ) , .B1( us01_n678 ) , .A( us01_n810 ) , .B2( us01_n814 ) );
  NOR2_X1 us01_U288 (.ZN( us01_n518 ) , .A2( us01_n706 ) , .A1( us01_n812 ) );
  AOI21_X1 us01_U289 (.ZN( us01_n475 ) , .A( us01_n667 ) , .B1( us01_n748 ) , .B2( us01_n804 ) );
  AOI221_X1 us01_U29 (.ZN( us01_n466 ) , .C2( us01_n712 ) , .B2( us01_n829 ) , .C1( us01_n843 ) , .B1( us01_n858 ) , .A( us01_n862 ) );
  NOR2_X1 us01_U290 (.ZN( us01_n566 ) , .A1( us01_n727 ) , .A2( us01_n760 ) );
  NOR2_X1 us01_U291 (.ZN( us01_n580 ) , .A1( us01_n742 ) , .A2( us01_n813 ) );
  AOI21_X1 us01_U292 (.ZN( us01_n591 ) , .B1( us01_n748 ) , .A( us01_n790 ) , .B2( us01_n811 ) );
  NOR2_X1 us01_U293 (.ZN( us01_n564 ) , .A2( us01_n695 ) , .A1( us01_n761 ) );
  AOI21_X1 us01_U294 (.ZN( us01_n512 ) , .A( us01_n777 ) , .B2( us01_n790 ) , .B1( us01_n810 ) );
  NAND2_X2 us01_U295 (.A2( us01_n462 ) , .A1( us01_n463 ) , .ZN( us01_n810 ) );
  AOI21_X1 us01_U296 (.ZN( us01_n637 ) , .B2( us01_n747 ) , .A( us01_n786 ) , .B1( us01_n810 ) );
  NOR2_X1 us01_U297 (.ZN( us01_n557 ) , .A2( us01_n789 ) , .A1( us01_n801 ) );
  NOR2_X1 us01_U298 (.A2( us01_n811 ) , .A1( us01_n813 ) , .ZN( us01_n819 ) );
  NOR2_X1 us01_U299 (.ZN( us01_n527 ) , .A1( us01_n706 ) , .A2( us01_n777 ) );
  NAND2_X2 us01_U3 (.A1( us01_n447 ) , .A2( us01_n462 ) , .ZN( us01_n722 ) );
  NOR4_X1 us01_U30 (.A4( us01_n512 ) , .A3( us01_n513 ) , .A2( us01_n514 ) , .A1( us01_n515 ) , .ZN( us01_n522 ) );
  NOR2_X1 us01_U300 (.ZN( us01_n517 ) , .A2( us01_n697 ) , .A1( us01_n814 ) );
  NOR2_X1 us01_U301 (.ZN( us01_n681 ) , .A2( us01_n697 ) , .A1( us01_n801 ) );
  NOR2_X1 us01_U302 (.ZN( us01_n576 ) , .A1( us01_n706 ) , .A2( us01_n811 ) );
  INV_X1 us01_U303 (.A( us01_n813 ) , .ZN( us01_n853 ) );
  INV_X1 us01_U304 (.A( us01_n811 ) , .ZN( us01_n834 ) );
  AOI21_X1 us01_U305 (.ZN( us01_n448 ) , .B2( us01_n790 ) , .A( us01_n801 ) , .B1( us01_n813 ) );
  AOI21_X1 us01_U306 (.ZN( us01_n538 ) , .A( us01_n761 ) , .B2( us01_n777 ) , .B1( us01_n815 ) );
  AOI21_X1 us01_U307 (.ZN( us01_n496 ) , .A( us01_n722 ) , .B2( us01_n760 ) , .B1( us01_n812 ) );
  AOI21_X1 us01_U308 (.ZN( us01_n687 ) , .B2( us01_n747 ) , .B1( us01_n761 ) , .A( us01_n804 ) );
  AOI21_X1 us01_U309 (.B1( us01_n684 ) , .ZN( us01_n685 ) , .A( us01_n726 ) , .B2( us01_n759 ) );
  AOI222_X1 us01_U31 (.ZN( us01_n523 ) , .A1( us01_n832 ) , .B2( us01_n835 ) , .C1( us01_n842 ) , .C2( us01_n848 ) , .A2( us01_n850 ) , .B1( us01_n864 ) );
  NOR2_X1 us01_U310 (.ZN( us01_n581 ) , .A1( us01_n790 ) , .A2( us01_n815 ) );
  NOR2_X1 us01_U311 (.ZN( us01_n532 ) , .A1( us01_n722 ) , .A2( us01_n786 ) );
  NOR2_X1 us01_U312 (.ZN( us01_n630 ) , .A2( us01_n695 ) , .A1( us01_n722 ) );
  AOI21_X1 us01_U313 (.A( us01_n788 ) , .B2( us01_n789 ) , .B1( us01_n790 ) , .ZN( us01_n791 ) );
  AOI21_X1 us01_U314 (.A( us01_n731 ) , .ZN( us01_n732 ) , .B2( us01_n778 ) , .B1( us01_n790 ) );
  NOR2_X1 us01_U315 (.ZN( us01_n565 ) , .A1( us01_n745 ) , .A2( us01_n803 ) );
  AOI21_X1 us01_U316 (.ZN( us01_n567 ) , .B1( us01_n748 ) , .B2( us01_n760 ) , .A( us01_n778 ) );
  AOI21_X1 us01_U317 (.ZN( us01_n638 ) , .B2( us01_n745 ) , .A( us01_n790 ) , .B1( us01_n801 ) );
  AOI21_X1 us01_U318 (.ZN( us01_n562 ) , .B1( us01_n722 ) , .A( us01_n777 ) , .B2( us01_n789 ) );
  AOI21_X1 us01_U319 (.ZN( us01_n569 ) , .B2( us01_n695 ) , .B1( us01_n804 ) , .A( us01_n810 ) );
  NOR4_X1 us01_U32 (.A3( us01_n519 ) , .A1( us01_n520 ) , .ZN( us01_n521 ) , .A2( us01_n671 ) , .A4( us01_n767 ) );
  NOR2_X1 us01_U320 (.ZN( us01_n663 ) , .A1( us01_n778 ) , .A2( us01_n811 ) );
  NOR2_X1 us01_U321 (.ZN( us01_n578 ) , .A2( us01_n695 ) , .A1( us01_n789 ) );
  NOR2_X1 us01_U322 (.ZN( us01_n682 ) , .A1( us01_n789 ) , .A2( us01_n811 ) );
  NAND2_X2 us01_U323 (.A1( us01_n450 ) , .A2( us01_n463 ) , .ZN( us01_n667 ) );
  NAND2_X1 us01_U324 (.ZN( us01_n751 ) , .A1( us01_n761 ) , .A2( us01_n803 ) );
  NOR2_X1 us01_U325 (.ZN( us01_n709 ) , .A1( us01_n760 ) , .A2( us01_n761 ) );
  AOI21_X1 us01_U326 (.ZN( us01_n476 ) , .B2( us01_n695 ) , .A( us01_n747 ) , .B1( us01_n777 ) );
  NOR2_X1 us01_U327 (.ZN( us01_n680 ) , .A2( us01_n706 ) , .A1( us01_n815 ) );
  INV_X1 us01_U328 (.A( us01_n778 ) , .ZN( us01_n848 ) );
  OAI21_X1 us01_U329 (.A( us01_n729 ) , .B1( us01_n730 ) , .ZN( us01_n734 ) , .B2( us01_n803 ) );
  AOI221_X1 us01_U33 (.A( us01_n779 ) , .ZN( us01_n796 ) , .C2( us01_n835 ) , .B2( us01_n836 ) , .B1( us01_n863 ) , .C1( us01_n864 ) );
  OAI21_X1 us01_U330 (.ZN( us01_n729 ) , .A( us01_n831 ) , .B2( us01_n850 ) , .B1( us01_n871 ) );
  AOI21_X1 us01_U331 (.ZN( us01_n639 ) , .B1( us01_n678 ) , .A( us01_n789 ) , .B2( us01_n815 ) );
  AOI21_X1 us01_U332 (.ZN( us01_n440 ) , .A( us01_n697 ) , .B1( us01_n731 ) , .B2( us01_n748 ) );
  NAND2_X1 us01_U333 (.A1( us01_n697 ) , .A2( us01_n727 ) , .ZN( us01_n780 ) );
  NOR2_X1 us01_U334 (.ZN( us01_n468 ) , .A2( us01_n777 ) , .A1( us01_n813 ) );
  NOR2_X1 us01_U335 (.ZN( us01_n516 ) , .A1( us01_n706 ) , .A2( us01_n786 ) );
  NAND2_X2 us01_U336 (.A2( us01_n447 ) , .A1( us01_n450 ) , .ZN( us01_n761 ) );
  OAI21_X1 us01_U337 (.A( us01_n696 ) , .ZN( us01_n700 ) , .B2( us01_n748 ) , .B1( us01_n802 ) );
  OAI21_X1 us01_U338 (.ZN( us01_n696 ) , .B2( us01_n831 ) , .B1( us01_n836 ) , .A( us01_n858 ) );
  NOR2_X1 us01_U339 (.ZN( us01_n524 ) , .A1( us01_n722 ) , .A2( us01_n748 ) );
  NOR4_X1 us01_U34 (.A4( us01_n791 ) , .A3( us01_n792 ) , .A2( us01_n793 ) , .A1( us01_n794 ) , .ZN( us01_n795 ) );
  AOI21_X1 us01_U340 (.ZN( us01_n441 ) , .B1( us01_n787 ) , .B2( us01_n789 ) , .A( us01_n812 ) );
  AOI21_X1 us01_U341 (.ZN( us01_n495 ) , .A( us01_n777 ) , .B2( us01_n789 ) , .B1( us01_n802 ) );
  NAND2_X1 us01_U342 (.ZN( us01_n712 ) , .A1( us01_n726 ) , .A2( us01_n778 ) );
  NOR2_X1 us01_U343 (.ZN( us01_n482 ) , .A1( us01_n786 ) , .A2( us01_n803 ) );
  NAND2_X1 us01_U344 (.A2( us01_n760 ) , .A1( us01_n804 ) , .ZN( us01_n808 ) );
  OAI21_X1 us01_U345 (.A( us01_n785 ) , .B2( us01_n786 ) , .B1( us01_n787 ) , .ZN( us01_n793 ) );
  OAI21_X1 us01_U346 (.ZN( us01_n785 ) , .A( us01_n837 ) , .B1( us01_n861 ) , .B2( us01_n871 ) );
  INV_X1 us01_U347 (.A( us01_n783 ) , .ZN( us01_n844 ) );
  NOR2_X1 us01_U348 (.ZN( us01_n710 ) , .A2( us01_n722 ) , .A1( us01_n788 ) );
  NAND2_X1 us01_U349 (.ZN( us01_n669 ) , .A1( us01_n804 ) , .A2( us01_n814 ) );
  NOR4_X1 us01_U35 (.A4( us01_n774 ) , .A3( us01_n775 ) , .A1( us01_n776 ) , .ZN( us01_n797 ) , .A2( us01_n799 ) );
  NAND2_X2 us01_U350 (.A2( us01_n446 ) , .A1( us01_n450 ) , .ZN( us01_n727 ) );
  INV_X1 us01_U351 (.A( us01_n722 ) , .ZN( us01_n854 ) );
  NAND2_X2 us01_U352 (.A1( us01_n445 ) , .A2( us01_n463 ) , .ZN( us01_n747 ) );
  INV_X1 us01_U353 (.A( us01_n815 ) , .ZN( us01_n842 ) );
  AND2_X1 us01_U354 (.ZN( us01_n730 ) , .A1( us01_n777 ) , .A2( us01_n783 ) );
  NAND2_X1 us01_U355 (.A1( us01_n445 ) , .A2( us01_n447 ) , .ZN( us01_n803 ) );
  NAND2_X1 us01_U356 (.A1( us01_n449 ) , .A2( us01_n452 ) , .ZN( us01_n812 ) );
  NAND2_X1 us01_U357 (.A1( us01_n453 ) , .A2( us01_n469 ) , .ZN( us01_n801 ) );
  NAND2_X1 us01_U358 (.A1( us01_n453 ) , .A2( us01_n460 ) , .ZN( us01_n748 ) );
  NAND2_X2 us01_U359 (.A2( us01_n446 ) , .A1( us01_n458 ) , .ZN( us01_n726 ) );
  NOR2_X1 us01_U36 (.ZN( us01_n802 ) , .A1( us01_n852 ) , .A2( us01_n859 ) );
  NAND2_X1 us01_U360 (.A2( us01_n451 ) , .A1( us01_n453 ) , .ZN( us01_n804 ) );
  NAND2_X1 us01_U361 (.A1( us01_n449 ) , .A2( us01_n469 ) , .ZN( us01_n814 ) );
  NAND2_X1 us01_U362 (.A1( us01_n452 ) , .A2( us01_n459 ) , .ZN( us01_n811 ) );
  NAND2_X1 us01_U363 (.A1( us01_n451 ) , .A2( us01_n459 ) , .ZN( us01_n742 ) );
  NAND2_X1 us01_U364 (.A1( us01_n451 ) , .A2( us01_n470 ) , .ZN( us01_n783 ) );
  NAND2_X1 us01_U365 (.A2( us01_n452 ) , .A1( us01_n470 ) , .ZN( us01_n777 ) );
  NAND2_X1 us01_U366 (.A2( us01_n459 ) , .A1( us01_n460 ) , .ZN( us01_n745 ) );
  NAND2_X2 us01_U367 (.A2( us01_n446 ) , .A1( us01_n462 ) , .ZN( us01_n813 ) );
  NAND2_X1 us01_U368 (.A1( us01_n460 ) , .A2( us01_n470 ) , .ZN( us01_n786 ) );
  NOR2_X1 us01_U369 (.ZN( us01_n451 ) , .A1( us01_n824 ) , .A2( us01_n825 ) );
  NAND4_X1 us01_U37 (.ZN( sa01_sr_2 ) , .A4( us01_n641 ) , .A3( us01_n642 ) , .A2( us01_n643 ) , .A1( us01_n644 ) );
  NAND2_X1 us01_U371 (.A1( us01_n449 ) , .A2( us01_n460 ) , .ZN( us01_n788 ) );
  NAND2_X2 us01_U372 (.A1( us01_n447 ) , .A2( us01_n458 ) , .ZN( us01_n790 ) );
  NAND2_X2 us01_U373 (.A2( us01_n439 ) , .A1( us01_n450 ) , .ZN( us01_n789 ) );
  NAND2_X1 us01_U374 (.A2( us01_n452 ) , .A1( us01_n453 ) , .ZN( us01_n728 ) );
  NAND2_X2 us01_U377 (.A2( us01_n439 ) , .A1( us01_n445 ) , .ZN( us01_n782 ) );
  NOR2_X1 us01_U378 (.A2( sa01_7 ) , .ZN( us01_n458 ) , .A1( us01_n847 ) );
  AOI222_X1 us01_U38 (.B2( us01_n636 ) , .ZN( us01_n642 ) , .B1( us01_n839 ) , .A1( us01_n840 ) , .C2( us01_n844 ) , .C1( us01_n861 ) , .A2( us01_n863 ) );
  NOR2_X1 us01_U380 (.A2( sa01_1 ) , .ZN( us01_n469 ) , .A1( us01_n824 ) );
  NOR2_X1 us01_U381 (.A2( sa01_0 ) , .ZN( us01_n452 ) , .A1( us01_n825 ) );
  NOR2_X1 us01_U382 (.A2( sa01_0 ) , .A1( sa01_1 ) , .ZN( us01_n460 ) );
  NAND2_X2 us01_U383 (.A1( us01_n439 ) , .A2( us01_n458 ) , .ZN( us01_n697 ) );
  INV_X1 us01_U387 (.A( sa01_1 ) , .ZN( us01_n825 ) );
  INV_X1 us01_U388 (.A( sa01_0 ) , .ZN( us01_n824 ) );
  NOR4_X1 us01_U39 (.A4( us01_n637 ) , .A3( us01_n638 ) , .A2( us01_n639 ) , .A1( us01_n640 ) , .ZN( us01_n641 ) );
  NAND2_X1 us01_U391 (.A1( us01_n727 ) , .A2( us01_n782 ) , .ZN( us01_n809 ) );
  OAI22_X1 us01_U392 (.ZN( us01_n586 ) , .A2( us01_n745 ) , .B2( us01_n760 ) , .A1( us01_n761 ) , .B1( us01_n782 ) );
  AOI21_X1 us01_U393 (.ZN( us01_n590 ) , .B1( us01_n726 ) , .B2( us01_n782 ) , .A( us01_n788 ) );
  AOI21_X1 us01_U394 (.ZN( us01_n646 ) , .A( us01_n760 ) , .B2( us01_n782 ) , .B1( us01_n790 ) );
  AOI21_X1 us01_U395 (.ZN( us01_n621 ) , .B1( us01_n697 ) , .A( us01_n777 ) , .B2( us01_n782 ) );
  OAI22_X1 us01_U396 (.ZN( us01_n679 ) , .A1( us01_n697 ) , .A2( us01_n728 ) , .B2( us01_n782 ) , .B1( us01_n815 ) );
  OAI21_X1 us01_U397 (.A( us01_n611 ) , .ZN( us01_n614 ) , .B1( us01_n623 ) , .B2( us01_n782 ) );
  NOR2_X1 us01_U398 (.ZN( us01_n608 ) , .A1( us01_n782 ) , .A2( us01_n814 ) );
  INV_X2 us01_U399 (.A( us01_n747 ) , .ZN( us01_n861 ) );
  NAND2_X2 us01_U4 (.A1( us01_n439 ) , .A2( us01_n462 ) , .ZN( us01_n706 ) );
  NOR3_X1 us01_U40 (.A2( us01_n605 ) , .A1( us01_n606 ) , .ZN( us01_n644 ) , .A3( us01_n720 ) );
  OAI222_X1 us01_U400 (.A2( us01_n667 ) , .ZN( us01_n672 ) , .B1( us01_n745 ) , .B2( us01_n782 ) , .C2( us01_n786 ) , .C1( us01_n813 ) , .A1( us01_n815 ) );
  NOR2_X1 us01_U401 (.ZN( us01_n649 ) , .A1( us01_n782 ) , .A2( us01_n786 ) );
  NOR2_X1 us01_U402 (.ZN( us01_n598 ) , .A2( us01_n695 ) , .A1( us01_n782 ) );
  NOR2_X1 us01_U403 (.ZN( us01_n551 ) , .A2( us01_n742 ) , .A1( us01_n782 ) );
  INV_X1 us01_U404 (.A( us01_n782 ) , .ZN( us01_n859 ) );
  NAND2_X1 us01_U405 (.A2( us01_n459 ) , .A1( us01_n469 ) , .ZN( us01_n695 ) );
  OAI221_X1 us01_U407 (.A( us01_n781 ) , .C2( us01_n782 ) , .B2( us01_n783 ) , .B1( us01_n784 ) , .ZN( us01_n794 ) , .C1( us01_n811 ) );
  AOI21_X1 us01_U408 (.ZN( us01_n498 ) , .A( us01_n695 ) , .B1( us01_n706 ) , .B2( us01_n784 ) );
  OAI221_X1 us01_U409 (.A( us01_n694 ) , .ZN( us01_n701 ) , .C2( us01_n782 ) , .C1( us01_n783 ) , .B1( us01_n784 ) , .B2( us01_n804 ) );
  NAND4_X1 us01_U41 (.ZN( sa01_sr_7 ) , .A4( us01_n820 ) , .A3( us01_n821 ) , .A2( us01_n822 ) , .A1( us01_n823 ) );
  OAI22_X1 us01_U410 (.ZN( us01_n588 ) , .B1( us01_n728 ) , .B2( us01_n747 ) , .A2( us01_n784 ) , .A1( us01_n801 ) );
  AOI222_X1 us01_U411 (.ZN( us01_n511 ) , .C1( us01_n830 ) , .B2( us01_n835 ) , .A2( us01_n841 ) , .C2( us01_n860 ) , .B1( us01_n861 ) , .A1( us01_n864 ) );
  AOI222_X1 us01_U412 (.ZN( us01_n603 ) , .B2( us01_n669 ) , .B1( us01_n751 ) , .C2( us01_n829 ) , .A1( us01_n831 ) , .A2( us01_n860 ) , .C1( us01_n861 ) );
  AOI221_X1 us01_U413 (.A( us01_n481 ) , .ZN( us01_n486 ) , .B1( us01_n829 ) , .C2( us01_n842 ) , .C1( us01_n850 ) , .B2( us01_n860 ) );
  NAND2_X1 us01_U414 (.A2( us01_n747 ) , .A1( us01_n784 ) , .ZN( us01_n807 ) );
  NOR2_X1 us01_U415 (.ZN( us01_n610 ) , .A1( us01_n777 ) , .A2( us01_n784 ) );
  NOR2_X1 us01_U416 (.ZN( us01_n715 ) , .A2( us01_n742 ) , .A1( us01_n784 ) );
  OAI222_X1 us01_U417 (.ZN( us01_n615 ) , .B1( us01_n695 ) , .C1( us01_n722 ) , .C2( us01_n745 ) , .B2( us01_n784 ) , .A2( us01_n790 ) , .A1( us01_n814 ) );
  NOR2_X1 us01_U418 (.ZN( us01_n651 ) , .A1( us01_n760 ) , .A2( us01_n784 ) );
  NOR2_X1 us01_U419 (.ZN( us01_n552 ) , .A1( us01_n784 ) , .A2( us01_n811 ) );
  AOI222_X1 us01_U42 (.C2( us01_n807 ) , .B2( us01_n808 ) , .A2( us01_n809 ) , .ZN( us01_n821 ) , .C1( us01_n830 ) , .A1( us01_n837 ) , .B1( us01_n851 ) );
  NOR2_X1 us01_U420 (.ZN( us01_n787 ) , .A2( us01_n860 ) , .A1( us01_n866 ) );
  NOR2_X1 us01_U421 (.ZN( us01_n699 ) , .A2( us01_n784 ) , .A1( us01_n815 ) );
  NOR2_X1 us01_U422 (.A1( us01_n728 ) , .ZN( us01_n763 ) , .A2( us01_n784 ) );
  INV_X1 us01_U423 (.A( us01_n784 ) , .ZN( us01_n860 ) );
  INV_X1 us01_U428 (.A( sa01_6 ) , .ZN( us01_n847 ) );
  NOR4_X1 us01_U43 (.A4( us01_n816 ) , .A3( us01_n817 ) , .A2( us01_n818 ) , .A1( us01_n819 ) , .ZN( us01_n820 ) );
  NOR2_X1 us01_U431 (.A2( sa01_6 ) , .A1( sa01_7 ) , .ZN( us01_n462 ) );
  AOI221_X1 us01_U432 (.A( us01_n574 ) , .ZN( us01_n585 ) , .B2( us01_n829 ) , .C2( us01_n841 ) , .B1( us01_n852 ) , .C1( us01_n859 ) );
  AOI21_X1 us01_U433 (.ZN( us01_n574 ) , .B2( us01_n722 ) , .B1( us01_n746 ) , .A( us01_n783 ) );
  AOI211_X1 us01_U435 (.A( us01_n635 ) , .ZN( us01_n643 ) , .B( us01_n741 ) , .C2( us01_n837 ) , .C1( us01_n852 ) );
  NAND4_X1 us01_U436 (.A4( us01_n631 ) , .A3( us01_n632 ) , .A2( us01_n633 ) , .A1( us01_n634 ) , .ZN( us01_n741 ) );
  NAND3_X1 us01_U437 (.ZN( sa01_sr_6 ) , .A3( us01_n795 ) , .A2( us01_n796 ) , .A1( us01_n797 ) );
  NAND3_X1 us01_U438 (.ZN( sa01_sr_5 ) , .A3( us01_n756 ) , .A2( us01_n757 ) , .A1( us01_n758 ) );
  NAND3_X1 us01_U439 (.ZN( sa01_sr_4 ) , .A3( us01_n736 ) , .A2( us01_n737 ) , .A1( us01_n738 ) );
  AOI211_X1 us01_U44 (.B( us01_n805 ) , .A( us01_n806 ) , .ZN( us01_n822 ) , .C1( us01_n840 ) , .C2( us01_n848 ) );
  NAND3_X1 us01_U440 (.A3( us01_n673 ) , .A2( us01_n674 ) , .A1( us01_n675 ) , .ZN( us01_n805 ) );
  NAND3_X1 us01_U441 (.ZN( us01_n636 ) , .A3( us01_n706 ) , .A2( us01_n722 ) , .A1( us01_n790 ) );
  NAND3_X1 us01_U442 (.A3( us01_n616 ) , .A2( us01_n617 ) , .A1( us01_n618 ) , .ZN( us01_n723 ) );
  NAND3_X1 us01_U443 (.A3( us01_n583 ) , .A2( us01_n584 ) , .A1( us01_n585 ) , .ZN( us01_n619 ) );
  NAND3_X1 us01_U444 (.ZN( us01_n563 ) , .A3( us01_n678 ) , .A2( us01_n748 ) , .A1( us01_n783 ) );
  NAND3_X1 us01_U445 (.A3( us01_n521 ) , .A2( us01_n522 ) , .A1( us01_n523 ) , .ZN( us01_n740 ) );
  NAND3_X1 us01_U446 (.A3( us01_n510 ) , .A1( us01_n511 ) , .ZN( us01_n606 ) , .A2( us01_n869 ) );
  NAND3_X1 us01_U447 (.A3( us01_n465 ) , .A2( us01_n466 ) , .A1( us01_n467 ) , .ZN( us01_n775 ) );
  NAND4_X1 us01_U45 (.ZN( sa01_sr_0 ) , .A4( us01_n499 ) , .A3( us01_n500 ) , .A2( us01_n501 ) , .A1( us01_n502 ) );
  NOR4_X1 us01_U46 (.A4( us01_n496 ) , .A3( us01_n497 ) , .A2( us01_n498 ) , .ZN( us01_n499 ) , .A1( us01_n525 ) );
  AOI221_X1 us01_U47 (.A( us01_n495 ) , .ZN( us01_n500 ) , .B2( us01_n841 ) , .C1( us01_n844 ) , .C2( us01_n858 ) , .B1( us01_n860 ) );
  AOI211_X1 us01_U48 (.A( us01_n494 ) , .ZN( us01_n501 ) , .B( us01_n800 ) , .C2( us01_n837 ) , .C1( us01_n849 ) );
  NOR2_X1 us01_U49 (.ZN( us01_n746 ) , .A1( us01_n859 ) , .A2( us01_n860 ) );
  NAND2_X2 us01_U5 (.A2( us01_n458 ) , .A1( us01_n463 ) , .ZN( us01_n778 ) );
  NAND4_X1 us01_U50 (.ZN( sa01_sr_1 ) , .A4( us01_n593 ) , .A3( us01_n594 ) , .A2( us01_n595 ) , .A1( us01_n596 ) );
  AOI211_X1 us01_U51 (.B( us01_n587 ) , .A( us01_n588 ) , .ZN( us01_n594 ) , .C2( us01_n809 ) , .C1( us01_n831 ) );
  NOR4_X1 us01_U52 (.A4( us01_n589 ) , .A3( us01_n590 ) , .A2( us01_n591 ) , .A1( us01_n592 ) , .ZN( us01_n593 ) );
  AOI211_X1 us01_U53 (.A( us01_n586 ) , .ZN( us01_n595 ) , .B( us01_n619 ) , .C1( us01_n843 ) , .C2( us01_n853 ) );
  NOR2_X1 us01_U54 (.ZN( us01_n623 ) , .A2( us01_n834 ) , .A1( us01_n837 ) );
  NAND4_X1 us01_U55 (.A4( us01_n601 ) , .A3( us01_n602 ) , .A2( us01_n603 ) , .A1( us01_n604 ) , .ZN( us01_n720 ) );
  NOR3_X1 us01_U56 (.A1( us01_n597 ) , .ZN( us01_n602 ) , .A3( us01_n661 ) , .A2( us01_n768 ) );
  NOR4_X1 us01_U57 (.A3( us01_n598 ) , .A2( us01_n599 ) , .A1( us01_n600 ) , .ZN( us01_n601 ) , .A4( us01_n653 ) );
  AOI222_X1 us01_U58 (.ZN( us01_n604 ) , .A1( us01_n828 ) , .C2( us01_n835 ) , .B1( us01_n840 ) , .A2( us01_n854 ) , .B2( us01_n859 ) , .C1( us01_n866 ) );
  NOR4_X1 us01_U59 (.A4( us01_n575 ) , .A3( us01_n576 ) , .A2( us01_n577 ) , .ZN( us01_n584 ) , .A1( us01_n681 ) );
  INV_X1 us01_U6 (.A( us01_n667 ) , .ZN( us01_n863 ) );
  NOR4_X1 us01_U60 (.A1( us01_n582 ) , .ZN( us01_n583 ) , .A3( us01_n650 ) , .A2( us01_n660 ) , .A4( us01_n765 ) );
  NAND4_X1 us01_U61 (.A4( us01_n483 ) , .A3( us01_n484 ) , .A2( us01_n485 ) , .A1( us01_n486 ) , .ZN( us01_n776 ) );
  NOR4_X1 us01_U62 (.A4( us01_n482 ) , .ZN( us01_n485 ) , .A1( us01_n564 ) , .A2( us01_n579 ) , .A3( us01_n600 ) );
  NOR4_X1 us01_U63 (.ZN( us01_n483 ) , .A2( us01_n531 ) , .A1( us01_n556 ) , .A3( us01_n629 ) , .A4( us01_n716 ) );
  NOR4_X1 us01_U64 (.ZN( us01_n484 ) , .A1( us01_n505 ) , .A2( us01_n517 ) , .A4( us01_n544 ) , .A3( us01_n609 ) );
  NOR4_X1 us01_U65 (.A4( us01_n627 ) , .A3( us01_n628 ) , .A2( us01_n629 ) , .A1( us01_n630 ) , .ZN( us01_n631 ) );
  AOI211_X1 us01_U66 (.B( us01_n621 ) , .A( us01_n622 ) , .ZN( us01_n633 ) , .C2( us01_n834 ) , .C1( us01_n861 ) );
  NOR4_X1 us01_U67 (.A4( us01_n624 ) , .A3( us01_n625 ) , .A2( us01_n626 ) , .ZN( us01_n632 ) , .A1( us01_n662 ) );
  NAND4_X1 us01_U68 (.A4( us01_n655 ) , .A3( us01_n656 ) , .A2( us01_n657 ) , .A1( us01_n658 ) , .ZN( us01_n798 ) );
  NOR3_X1 us01_U69 (.A3( us01_n649 ) , .A2( us01_n650 ) , .A1( us01_n651 ) , .ZN( us01_n656 ) );
  NOR3_X1 us01_U7 (.ZN( us01_n596 ) , .A1( us01_n606 ) , .A3( us01_n721 ) , .A2( us01_n740 ) );
  NOR3_X1 us01_U70 (.A3( us01_n652 ) , .A2( us01_n653 ) , .A1( us01_n654 ) , .ZN( us01_n655 ) );
  NOR3_X1 us01_U71 (.A3( us01_n646 ) , .A2( us01_n647 ) , .A1( us01_n648 ) , .ZN( us01_n657 ) );
  NAND4_X1 us01_U72 (.A4( us01_n558 ) , .A3( us01_n559 ) , .A2( us01_n560 ) , .A1( us01_n561 ) , .ZN( us01_n605 ) );
  NOR4_X1 us01_U73 (.ZN( us01_n559 ) , .A1( us01_n651 ) , .A3( us01_n659 ) , .A4( us01_n683 ) , .A2( us01_n766 ) );
  NOR4_X1 us01_U74 (.A4( us01_n550 ) , .A3( us01_n551 ) , .A2( us01_n552 ) , .A1( us01_n553 ) , .ZN( us01_n560 ) );
  NOR4_X1 us01_U75 (.A4( us01_n554 ) , .A3( us01_n555 ) , .A2( us01_n556 ) , .A1( us01_n557 ) , .ZN( us01_n558 ) );
  NAND4_X1 us01_U76 (.A4( us01_n770 ) , .A3( us01_n771 ) , .A2( us01_n772 ) , .A1( us01_n773 ) , .ZN( us01_n799 ) );
  NOR3_X1 us01_U77 (.A3( us01_n763 ) , .A2( us01_n764 ) , .A1( us01_n765 ) , .ZN( us01_n771 ) );
  NOR4_X1 us01_U78 (.A4( us01_n766 ) , .A3( us01_n767 ) , .A2( us01_n768 ) , .A1( us01_n769 ) , .ZN( us01_n770 ) );
  AOI222_X1 us01_U79 (.ZN( us01_n773 ) , .A1( us01_n828 ) , .C1( us01_n832 ) , .B2( us01_n839 ) , .A2( us01_n848 ) , .B1( us01_n859 ) , .C2( us01_n871 ) );
  NOR3_X1 us01_U8 (.A3( us01_n798 ) , .A2( us01_n799 ) , .A1( us01_n800 ) , .ZN( us01_n823 ) );
  NOR4_X1 us01_U80 (.A4( us01_n507 ) , .A2( us01_n508 ) , .A1( us01_n509 ) , .ZN( us01_n510 ) , .A3( us01_n668 ) );
  INV_X1 us01_U81 (.A( us01_n503 ) , .ZN( us01_n869 ) );
  NOR4_X1 us01_U82 (.A4( us01_n663 ) , .A3( us01_n664 ) , .A2( us01_n665 ) , .A1( us01_n666 ) , .ZN( us01_n674 ) );
  NOR4_X1 us01_U83 (.A4( us01_n659 ) , .A3( us01_n660 ) , .A2( us01_n661 ) , .A1( us01_n662 ) , .ZN( us01_n675 ) );
  NOR4_X1 us01_U84 (.A3( us01_n671 ) , .A1( us01_n672 ) , .ZN( us01_n673 ) , .A4( us01_n713 ) , .A2( us01_n857 ) );
  NOR2_X1 us01_U85 (.ZN( us01_n759 ) , .A1( us01_n831 ) , .A2( us01_n832 ) );
  NAND4_X1 us01_U86 (.A4( us01_n454 ) , .A3( us01_n455 ) , .A2( us01_n456 ) , .A1( us01_n457 ) , .ZN( us01_n677 ) );
  NOR3_X1 us01_U87 (.ZN( us01_n455 ) , .A3( us01_n528 ) , .A1( us01_n553 ) , .A2( us01_n568 ) );
  AOI221_X1 us01_U88 (.A( us01_n448 ) , .ZN( us01_n457 ) , .C2( us01_n751 ) , .B1( us01_n830 ) , .C1( us01_n840 ) , .B2( us01_n859 ) );
  NOR4_X1 us01_U89 (.ZN( us01_n456 ) , .A2( us01_n507 ) , .A1( us01_n597 ) , .A4( us01_n626 ) , .A3( us01_n709 ) );
  NOR3_X1 us01_U9 (.A3( us01_n619 ) , .A2( us01_n620 ) , .ZN( us01_n634 ) , .A1( us01_n723 ) );
  NAND4_X1 us01_U90 (.A4( us01_n533 ) , .A3( us01_n534 ) , .A2( us01_n535 ) , .A1( us01_n536 ) , .ZN( us01_n620 ) );
  NOR4_X1 us01_U91 (.A4( us01_n524 ) , .A2( us01_n525 ) , .A1( us01_n526 ) , .ZN( us01_n536 ) , .A3( us01_n699 ) );
  NOR4_X1 us01_U92 (.A1( us01_n529 ) , .ZN( us01_n534 ) , .A2( us01_n652 ) , .A4( us01_n666 ) , .A3( us01_n763 ) );
  NOR4_X1 us01_U93 (.A4( us01_n527 ) , .A3( us01_n528 ) , .ZN( us01_n535 ) , .A2( us01_n682 ) , .A1( us01_n792 ) );
  NAND4_X1 us01_U94 (.A4( us01_n477 ) , .A3( us01_n478 ) , .A2( us01_n479 ) , .A1( us01_n480 ) , .ZN( us01_n692 ) );
  NOR3_X1 us01_U95 (.ZN( us01_n478 ) , .A2( us01_n506 ) , .A3( us01_n599 ) , .A1( us01_n608 ) );
  AOI211_X1 us01_U96 (.B( us01_n475 ) , .A( us01_n476 ) , .ZN( us01_n480 ) , .C2( us01_n831 ) , .C1( us01_n859 ) );
  NOR4_X1 us01_U97 (.ZN( us01_n479 ) , .A3( us01_n530 ) , .A4( us01_n543 ) , .A2( us01_n565 ) , .A1( us01_n715 ) );
  NAND4_X1 us01_U98 (.A4( us01_n546 ) , .A3( us01_n547 ) , .A2( us01_n548 ) , .A1( us01_n549 ) , .ZN( us01_n743 ) );
  NOR3_X1 us01_U99 (.ZN( us01_n547 ) , .A2( us01_n649 ) , .A1( us01_n665 ) , .A3( us01_n769 ) );
  NOR3_X1 us11_U10 (.ZN( us11_n504 ) , .A2( us11_n679 ) , .A3( us11_n777 ) , .A1( us11_n876 ) );
  NOR4_X1 us11_U100 (.A4( us11_n529 ) , .A3( us11_n530 ) , .ZN( us11_n537 ) , .A2( us11_n684 ) , .A1( us11_n794 ) );
  NAND4_X1 us11_U101 (.A4( us11_n479 ) , .A3( us11_n480 ) , .A2( us11_n481 ) , .A1( us11_n482 ) , .ZN( us11_n694 ) );
  NOR3_X1 us11_U102 (.ZN( us11_n480 ) , .A2( us11_n508 ) , .A3( us11_n601 ) , .A1( us11_n610 ) );
  AOI211_X1 us11_U103 (.B( us11_n477 ) , .A( us11_n478 ) , .ZN( us11_n482 ) , .C2( us11_n833 ) , .C1( us11_n861 ) );
  NOR4_X1 us11_U104 (.ZN( us11_n481 ) , .A3( us11_n532 ) , .A4( us11_n545 ) , .A2( us11_n567 ) , .A1( us11_n717 ) );
  NAND4_X1 us11_U105 (.A4( us11_n548 ) , .A3( us11_n549 ) , .A2( us11_n550 ) , .A1( us11_n551 ) , .ZN( us11_n745 ) );
  NOR3_X1 us11_U106 (.ZN( us11_n549 ) , .A2( us11_n651 ) , .A1( us11_n667 ) , .A3( us11_n771 ) );
  AOI211_X1 us11_U107 (.B( us11_n539 ) , .A( us11_n540 ) , .ZN( us11_n551 ) , .C2( us11_n839 ) , .C1( us11_n851 ) );
  NOR4_X1 us11_U108 (.A4( us11_n544 ) , .A3( us11_n545 ) , .A2( us11_n546 ) , .A1( us11_n547 ) , .ZN( us11_n548 ) );
  NOR4_X1 us11_U109 (.ZN( us11_n620 ) , .A1( us11_n656 ) , .A3( us11_n666 ) , .A4( us11_n682 ) , .A2( us11_n766 ) );
  INV_X1 us11_U11 (.A( us11_n706 ) , .ZN( us11_n876 ) );
  NOR4_X1 us11_U110 (.A4( us11_n609 ) , .A3( us11_n610 ) , .A2( us11_n611 ) , .A1( us11_n612 ) , .ZN( us11_n619 ) );
  NOR4_X1 us11_U111 (.A4( us11_n614 ) , .A3( us11_n615 ) , .A2( us11_n616 ) , .A1( us11_n617 ) , .ZN( us11_n618 ) );
  NOR2_X1 us11_U112 (.ZN( us11_n686 ) , .A1( us11_n831 ) , .A2( us11_n832 ) );
  NAND4_X1 us11_U113 (.A4( us11_n473 ) , .A3( us11_n474 ) , .A2( us11_n475 ) , .A1( us11_n476 ) , .ZN( us11_n678 ) );
  NOR4_X1 us11_U114 (.A4( us11_n470 ) , .ZN( us11_n476 ) , .A3( us11_n556 ) , .A1( us11_n735 ) , .A2( us11_n755 ) );
  NOR4_X1 us11_U115 (.ZN( us11_n475 ) , .A1( us11_n531 ) , .A3( us11_n568 ) , .A4( us11_n600 ) , .A2( us11_n642 ) );
  NOR4_X1 us11_U116 (.ZN( us11_n474 ) , .A1( us11_n506 ) , .A3( us11_n544 ) , .A2( us11_n583 ) , .A4( us11_n716 ) );
  NAND4_X1 us11_U117 (.A4( us11_n691 ) , .A3( us11_n692 ) , .A1( us11_n693 ) , .ZN( us11_n776 ) , .A2( us11_n872 ) );
  INV_X1 us11_U118 (.A( us11_n679 ) , .ZN( us11_n872 ) );
  NOR4_X1 us11_U119 (.A4( us11_n687 ) , .A3( us11_n688 ) , .A2( us11_n689 ) , .A1( us11_n690 ) , .ZN( us11_n691 ) );
  NOR3_X1 us11_U12 (.A3( us11_n621 ) , .A2( us11_n622 ) , .ZN( us11_n636 ) , .A1( us11_n725 ) );
  AOI221_X1 us11_U120 (.A( us11_n681 ) , .ZN( us11_n692 ) , .B2( us11_n840 ) , .C1( us11_n842 ) , .C2( us11_n862 ) , .B1( us11_n865 ) );
  NOR2_X1 us11_U121 (.ZN( us11_n733 ) , .A2( us11_n832 ) , .A1( us11_n845 ) );
  NAND4_X1 us11_U122 (.A4( us11_n719 ) , .A3( us11_n720 ) , .A2( us11_n721 ) , .ZN( us11_n741 ) , .A1( us11_n857 ) );
  AOI221_X1 us11_U123 (.A( us11_n710 ) , .ZN( us11_n721 ) , .C2( us11_n844 ) , .B2( us11_n845 ) , .C1( us11_n861 ) , .B1( us11_n862 ) );
  INV_X1 us11_U124 (.A( us11_n709 ) , .ZN( us11_n857 ) );
  NOR4_X1 us11_U125 (.A4( us11_n715 ) , .A3( us11_n716 ) , .A2( us11_n717 ) , .A1( us11_n718 ) , .ZN( us11_n719 ) );
  NAND4_X1 us11_U126 (.A4( us11_n573 ) , .A3( us11_n574 ) , .A1( us11_n575 ) , .ZN( us11_n723 ) , .A2( us11_n874 ) );
  NOR4_X1 us11_U127 (.A4( us11_n569 ) , .A3( us11_n570 ) , .A2( us11_n571 ) , .A1( us11_n572 ) , .ZN( us11_n573 ) );
  INV_X1 us11_U128 (.A( us11_n607 ) , .ZN( us11_n874 ) );
  NOR2_X1 us11_U129 (.ZN( us11_n575 ) , .A1( us11_n622 ) , .A2( us11_n745 ) );
  NOR2_X1 us11_U13 (.ZN( us11_n495 ) , .A1( us11_n678 ) , .A2( us11_n694 ) );
  NAND4_X1 us11_U130 (.A4( us11_n493 ) , .A3( us11_n494 ) , .A1( us11_n495 ) , .ZN( us11_n802 ) , .A2( us11_n867 ) );
  AOI221_X1 us11_U131 (.A( us11_n489 ) , .ZN( us11_n494 ) , .B2( us11_n836 ) , .C2( us11_n841 ) , .C1( us11_n851 ) , .B1( us11_n860 ) );
  INV_X1 us11_U132 (.A( us11_n778 ) , .ZN( us11_n867 ) );
  NOR4_X1 us11_U133 (.A2( us11_n491 ) , .A1( us11_n492 ) , .ZN( us11_n493 ) , .A3( us11_n580 ) , .A4( us11_n612 ) );
  NOR2_X1 us11_U134 (.ZN( us11_n647 ) , .A1( us11_n854 ) , .A2( us11_n868 ) );
  INV_X1 us11_U135 (.A( us11_n762 ) , .ZN( us11_n830 ) );
  NAND4_X1 us11_U136 (.A4( us11_n633 ) , .A3( us11_n634 ) , .A2( us11_n635 ) , .A1( us11_n636 ) , .ZN( us11_n743 ) );
  AOI211_X1 us11_U137 (.B( us11_n623 ) , .A( us11_n624 ) , .ZN( us11_n635 ) , .C2( us11_n836 ) , .C1( us11_n863 ) );
  NOR4_X1 us11_U138 (.A4( us11_n629 ) , .A3( us11_n630 ) , .A2( us11_n631 ) , .A1( us11_n632 ) , .ZN( us11_n633 ) );
  NOR4_X1 us11_U139 (.A4( us11_n626 ) , .A3( us11_n627 ) , .A2( us11_n628 ) , .ZN( us11_n634 ) , .A1( us11_n664 ) );
  NOR2_X1 us11_U14 (.A1( us11_n678 ) , .ZN( us11_n693 ) , .A2( us11_n807 ) );
  OR4_X1 us11_U140 (.A4( us11_n566 ) , .A3( us11_n567 ) , .A2( us11_n568 ) , .ZN( us11_n572 ) , .A1( us11_n665 ) );
  OR4_X1 us11_U141 (.A4( us11_n518 ) , .A2( us11_n519 ) , .A1( us11_n520 ) , .ZN( us11_n522 ) , .A3( us11_n821 ) );
  OR4_X1 us11_U142 (.ZN( us11_n492 ) , .A4( us11_n534 ) , .A2( us11_n547 ) , .A1( us11_n559 ) , .A3( us11_n632 ) );
  OR4_X1 us11_U143 (.A4( us11_n682 ) , .A3( us11_n683 ) , .A2( us11_n684 ) , .A1( us11_n685 ) , .ZN( us11_n690 ) );
  OR4_X1 us11_U144 (.ZN( us11_n466 ) , .A4( us11_n518 ) , .A3( us11_n529 ) , .A2( us11_n578 ) , .A1( us11_n712 ) );
  INV_X1 us11_U145 (.A( us11_n697 ) , .ZN( us11_n838 ) );
  OR4_X1 us11_U146 (.A4( us11_n580 ) , .A3( us11_n581 ) , .A2( us11_n582 ) , .A1( us11_n583 ) , .ZN( us11_n584 ) );
  NAND2_X1 us11_U147 (.ZN( us11_n613 ) , .A2( us11_n837 ) , .A1( us11_n873 ) );
  OR3_X1 us11_U148 (.A3( us11_n506 ) , .A2( us11_n507 ) , .A1( us11_n508 ) , .ZN( us11_n511 ) );
  INV_X1 us11_U149 (.A( us11_n463 ) , .ZN( us11_n864 ) );
  INV_X1 us11_U15 (.A( us11_n680 ) , .ZN( us11_n840 ) );
  OAI21_X1 us11_U150 (.ZN( us11_n463 ) , .B1( us11_n809 ) , .A( us11_n834 ) , .B2( us11_n851 ) );
  INV_X1 us11_U151 (.A( us11_n754 ) , .ZN( us11_n869 ) );
  OAI21_X1 us11_U152 (.B1( us11_n753 ) , .ZN( us11_n754 ) , .A( us11_n845 ) , .B2( us11_n868 ) );
  INV_X1 us11_U153 (.A( us11_n672 ) , .ZN( us11_n859 ) );
  AOI21_X1 us11_U154 (.A( us11_n670 ) , .B1( us11_n671 ) , .ZN( us11_n672 ) , .B2( us11_n856 ) );
  AOI222_X1 us11_U155 (.ZN( us11_n660 ) , .A2( us11_n839 ) , .B1( us11_n841 ) , .C2( us11_n845 ) , .A1( us11_n860 ) , .C1( us11_n863 ) , .B2( us11_n870 ) );
  INV_X1 us11_U156 (.A( us11_n647 ) , .ZN( us11_n870 ) );
  NAND2_X1 us11_U157 (.A1( us11_n447 ) , .A2( us11_n465 ) , .ZN( us11_n749 ) );
  OAI222_X1 us11_U158 (.ZN( us11_n617 ) , .B1( us11_n697 ) , .C1( us11_n724 ) , .C2( us11_n747 ) , .B2( us11_n786 ) , .A2( us11_n792 ) , .A1( us11_n816 ) );
  OAI222_X1 us11_U159 (.B2( us11_n708 ) , .ZN( us11_n709 ) , .C2( us11_n724 ) , .B1( us11_n747 ) , .A1( us11_n806 ) , .C1( us11_n814 ) , .A2( us11_n815 ) );
  NOR4_X1 us11_U16 (.A4( us11_n445 ) , .A3( us11_n446 ) , .A2( us11_n516 ) , .A1( us11_n541 ) , .ZN( us11_n706 ) );
  AOI22_X1 us11_U160 (.ZN( us11_n696 ) , .A1( us11_n830 ) , .B2( us11_n843 ) , .A2( us11_n865 ) , .B1( us11_n868 ) );
  AOI22_X1 us11_U161 (.A2( us11_n782 ) , .ZN( us11_n783 ) , .B2( us11_n831 ) , .A1( us11_n834 ) , .B1( us11_n863 ) );
  INV_X1 us11_U162 (.A( us11_n730 ) , .ZN( us11_n839 ) );
  AOI221_X1 us11_U163 (.A( us11_n564 ) , .C2( us11_n565 ) , .ZN( us11_n574 ) , .B2( us11_n845 ) , .B1( us11_n852 ) , .C1( us11_n853 ) );
  AOI21_X1 us11_U164 (.ZN( us11_n564 ) , .B1( us11_n724 ) , .A( us11_n779 ) , .B2( us11_n791 ) );
  NAND2_X1 us11_U165 (.A1( us11_n451 ) , .A2( us11_n453 ) , .ZN( us11_n762 ) );
  INV_X1 us11_U166 (.A( us11_n790 ) , .ZN( us11_n832 ) );
  OAI22_X1 us11_U167 (.ZN( us11_n637 ) , .A1( us11_n699 ) , .B2( us11_n728 ) , .A2( us11_n762 ) , .B1( us11_n816 ) );
  OAI221_X1 us11_U168 (.A( us11_n727 ) , .C2( us11_n728 ) , .B2( us11_n729 ) , .B1( us11_n730 ) , .ZN( us11_n737 ) , .C1( us11_n817 ) );
  AOI22_X1 us11_U169 (.ZN( us11_n727 ) , .B1( us11_n832 ) , .A2( us11_n838 ) , .A1( us11_n863 ) , .B2( us11_n866 ) );
  OR3_X1 us11_U17 (.ZN( us11_n446 ) , .A1( us11_n528 ) , .A3( us11_n577 ) , .A2( us11_n875 ) );
  INV_X1 us11_U170 (.A( us11_n747 ) , .ZN( us11_n834 ) );
  OAI22_X1 us11_U171 (.ZN( us11_n624 ) , .B1( us11_n669 ) , .B2( us11_n747 ) , .A1( us11_n815 ) , .A2( us11_n816 ) );
  OAI22_X1 us11_U172 (.ZN( us11_n489 ) , .A1( us11_n724 ) , .B2( us11_n728 ) , .B1( us11_n730 ) , .A2( us11_n779 ) );
  OAI22_X1 us11_U173 (.B2( us11_n779 ) , .B1( us11_n780 ) , .ZN( us11_n781 ) , .A2( us11_n814 ) , .A1( us11_n815 ) );
  OAI22_X1 us11_U174 (.A1( us11_n724 ) , .ZN( us11_n726 ) , .B2( us11_n750 ) , .B1( us11_n812 ) , .A2( us11_n816 ) );
  NOR2_X1 us11_U175 (.ZN( us11_n630 ) , .A1( us11_n747 ) , .A2( us11_n815 ) );
  OAI22_X1 us11_U176 (.B2( us11_n750 ) , .B1( us11_n751 ) , .A1( us11_n752 ) , .ZN( us11_n756 ) , .A2( us11_n806 ) );
  NOR3_X1 us11_U177 (.ZN( us11_n752 ) , .A2( us11_n853 ) , .A1( us11_n863 ) , .A3( us11_n865 ) );
  NOR2_X1 us11_U178 (.ZN( us11_n751 ) , .A2( us11_n852 ) , .A1( us11_n860 ) );
  OAI22_X1 us11_U179 (.B2( us11_n803 ) , .B1( us11_n804 ) , .A2( us11_n805 ) , .A1( us11_n806 ) , .ZN( us11_n808 ) );
  OR4_X1 us11_U18 (.A4( us11_n442 ) , .A2( us11_n443 ) , .A1( us11_n444 ) , .ZN( us11_n445 ) , .A3( us11_n553 ) );
  NOR2_X1 us11_U180 (.ZN( us11_n656 ) , .A1( us11_n747 ) , .A2( us11_n780 ) );
  OAI22_X1 us11_U181 (.B2( us11_n744 ) , .ZN( us11_n746 ) , .A2( us11_n762 ) , .B1( us11_n780 ) , .A1( us11_n792 ) );
  OAI22_X1 us11_U182 (.ZN( us11_n496 ) , .A2( us11_n744 ) , .A1( us11_n780 ) , .B1( us11_n791 ) , .B2( us11_n806 ) );
  OAI22_X1 us11_U183 (.ZN( us11_n695 ) , .A2( us11_n730 ) , .A1( us11_n780 ) , .B1( us11_n791 ) , .B2( us11_n817 ) );
  INV_X1 us11_U184 (.A( us11_n744 ) , .ZN( us11_n837 ) );
  INV_X1 us11_U185 (.A( us11_n805 ) , .ZN( us11_n860 ) );
  INV_X1 us11_U186 (.A( us11_n816 ) , .ZN( us11_n831 ) );
  INV_X1 us11_U187 (.A( us11_n788 ) , .ZN( us11_n845 ) );
  OAI22_X1 us11_U188 (.ZN( us11_n590 ) , .B1( us11_n730 ) , .B2( us11_n749 ) , .A2( us11_n786 ) , .A1( us11_n803 ) );
  OAI22_X1 us11_U189 (.B1( us11_n490 ) , .ZN( us11_n491 ) , .A1( us11_n686 ) , .A2( us11_n763 ) , .B2( us11_n817 ) );
  INV_X1 us11_U19 (.A( us11_n613 ) , .ZN( us11_n875 ) );
  NOR3_X1 us11_U190 (.ZN( us11_n490 ) , .A1( us11_n782 ) , .A2( us11_n850 ) , .A3( us11_n863 ) );
  OAI22_X1 us11_U191 (.ZN( us11_n710 ) , .A2( us11_n728 ) , .B2( us11_n729 ) , .A1( us11_n744 ) , .B1( us11_n813 ) );
  INV_X1 us11_U192 (.A( us11_n792 ) , .ZN( us11_n851 ) );
  NOR2_X1 us11_U193 (.ZN( us11_n715 ) , .A1( us11_n805 ) , .A2( us11_n817 ) );
  NOR2_X1 us11_U194 (.A1( us11_n699 ) , .ZN( us11_n768 ) , .A2( us11_n813 ) );
  NOR2_X1 us11_U195 (.ZN( us11_n541 ) , .A2( us11_n697 ) , .A1( us11_n699 ) );
  INV_X1 us11_U196 (.A( us11_n814 ) , .ZN( us11_n833 ) );
  NOR2_X1 us11_U197 (.A1( us11_n669 ) , .ZN( us11_n673 ) , .A2( us11_n744 ) );
  NOR2_X1 us11_U198 (.ZN( us11_n602 ) , .A1( us11_n669 ) , .A2( us11_n803 ) );
  NOR2_X1 us11_U199 (.A1( us11_n669 ) , .ZN( us11_n688 ) , .A2( us11_n816 ) );
  INV_X1 us11_U20 (.A( us11_n749 ) , .ZN( us11_n863 ) );
  NOR2_X1 us11_U200 (.A2( us11_n744 ) , .ZN( us11_n755 ) , .A1( us11_n805 ) );
  NOR2_X1 us11_U201 (.ZN( us11_n735 ) , .A2( us11_n803 ) , .A1( us11_n805 ) );
  NOR2_X1 us11_U202 (.A1( us11_n669 ) , .ZN( us11_n766 ) , .A2( us11_n813 ) );
  NOR2_X1 us11_U203 (.ZN( us11_n527 ) , .A1( us11_n669 ) , .A2( us11_n779 ) );
  NOR2_X1 us11_U204 (.ZN( us11_n666 ) , .A1( us11_n728 ) , .A2( us11_n803 ) );
  NOR2_X1 us11_U205 (.ZN( us11_n594 ) , .A2( us11_n697 ) , .A1( us11_n728 ) );
  NOR2_X1 us11_U206 (.ZN( us11_n718 ) , .A2( us11_n724 ) , .A1( us11_n744 ) );
  NOR2_X1 us11_U207 (.ZN( us11_n570 ) , .A1( us11_n728 ) , .A2( us11_n806 ) );
  NOR2_X1 us11_U208 (.ZN( us11_n661 ) , .A1( us11_n729 ) , .A2( us11_n790 ) );
  OAI22_X1 us11_U209 (.ZN( us11_n483 ) , .A1( us11_n708 ) , .B2( us11_n785 ) , .A2( us11_n806 ) , .B1( us11_n812 ) );
  AOI222_X1 us11_U21 (.ZN( us11_n563 ) , .B1( us11_n830 ) , .C1( us11_n841 ) , .A2( us11_n843 ) , .A1( us11_n854 ) , .B2( us11_n863 ) , .C2( us11_n873 ) );
  NOR2_X1 us11_U210 (.ZN( us11_n601 ) , .A2( us11_n780 ) , .A1( us11_n803 ) );
  NOR2_X1 us11_U211 (.ZN( us11_n531 ) , .A2( us11_n780 ) , .A1( us11_n816 ) );
  NOR2_X1 us11_U212 (.ZN( us11_n654 ) , .A1( us11_n728 ) , .A2( us11_n813 ) );
  NOR2_X1 us11_U213 (.ZN( us11_n509 ) , .A1( us11_n729 ) , .A2( us11_n779 ) );
  NOR2_X1 us11_U214 (.ZN( us11_n599 ) , .A2( us11_n791 ) , .A1( us11_n816 ) );
  NOR2_X1 us11_U215 (.ZN( us11_n612 ) , .A1( us11_n779 ) , .A2( us11_n786 ) );
  NOR2_X1 us11_U216 (.ZN( us11_n546 ) , .A2( us11_n780 ) , .A1( us11_n814 ) );
  INV_X1 us11_U217 (.A( us11_n750 ) , .ZN( us11_n842 ) );
  NOR2_X1 us11_U218 (.ZN( us11_n532 ) , .A2( us11_n749 ) , .A1( us11_n750 ) );
  NOR2_X1 us11_U219 (.ZN( us11_n528 ) , .A2( us11_n724 ) , .A1( us11_n803 ) );
  NOR4_X1 us11_U22 (.ZN( us11_n479 ) , .A1( us11_n520 ) , .A4( us11_n557 ) , .A3( us11_n582 ) , .A2( us11_n630 ) );
  NOR2_X1 us11_U220 (.ZN( us11_n577 ) , .A2( us11_n699 ) , .A1( us11_n814 ) );
  AOI21_X1 us11_U221 (.ZN( us11_n640 ) , .B2( us11_n747 ) , .A( us11_n792 ) , .B1( us11_n803 ) );
  NOR2_X1 us11_U222 (.ZN( us11_n615 ) , .A1( us11_n785 ) , .A2( us11_n815 ) );
  NOR2_X1 us11_U223 (.ZN( us11_n629 ) , .A2( us11_n728 ) , .A1( us11_n785 ) );
  NOR2_X1 us11_U224 (.ZN( us11_n663 ) , .A1( us11_n729 ) , .A2( us11_n785 ) );
  NOR2_X1 us11_U225 (.ZN( us11_n628 ) , .A2( us11_n669 ) , .A1( us11_n785 ) );
  NOR2_X1 us11_U226 (.ZN( us11_n611 ) , .A2( us11_n780 ) , .A1( us11_n806 ) );
  NOR2_X1 us11_U227 (.A2( us11_n744 ) , .ZN( us11_n769 ) , .A1( us11_n812 ) );
  NOR2_X1 us11_U228 (.ZN( us11_n567 ) , .A1( us11_n747 ) , .A2( us11_n805 ) );
  NOR2_X1 us11_U229 (.A2( us11_n708 ) , .A1( us11_n750 ) , .ZN( us11_n771 ) );
  NOR4_X1 us11_U23 (.ZN( us11_n473 ) , .A2( us11_n521 ) , .A4( us11_n594 ) , .A1( us11_n609 ) , .A3( us11_n629 ) );
  NOR2_X1 us11_U230 (.ZN( us11_n557 ) , .A1( us11_n792 ) , .A2( us11_n814 ) );
  NOR2_X1 us11_U231 (.A2( us11_n697 ) , .ZN( us11_n716 ) , .A1( us11_n792 ) );
  NOR2_X1 us11_U232 (.ZN( us11_n544 ) , .A2( us11_n785 ) , .A1( us11_n792 ) );
  NOR2_X1 us11_U233 (.ZN( us11_n667 ) , .A1( us11_n750 ) , .A2( us11_n815 ) );
  NOR2_X1 us11_U234 (.ZN( us11_n555 ) , .A1( us11_n750 ) , .A2( us11_n791 ) );
  NOR2_X1 us11_U235 (.ZN( us11_n508 ) , .A2( us11_n780 ) , .A1( us11_n785 ) );
  NOR2_X1 us11_U236 (.ZN( us11_n543 ) , .A2( us11_n708 ) , .A1( us11_n785 ) );
  NOR2_X1 us11_U237 (.ZN( us11_n664 ) , .A1( us11_n785 ) , .A2( us11_n791 ) );
  OAI22_X1 us11_U238 (.B1( us11_n440 ) , .ZN( us11_n444 ) , .A2( us11_n728 ) , .A1( us11_n744 ) , .B2( us11_n749 ) );
  NOR3_X1 us11_U239 (.ZN( us11_n440 ) , .A2( us11_n836 ) , .A3( us11_n837 ) , .A1( us11_n846 ) );
  NOR4_X1 us11_U24 (.ZN( us11_n485 ) , .A2( us11_n533 ) , .A1( us11_n558 ) , .A3( us11_n631 ) , .A4( us11_n718 ) );
  NOR2_X1 us11_U240 (.ZN( us11_n631 ) , .A1( us11_n724 ) , .A2( us11_n813 ) );
  NOR2_X1 us11_U241 (.ZN( us11_n556 ) , .A1( us11_n762 ) , .A2( us11_n805 ) );
  NOR2_X1 us11_U242 (.ZN( us11_n530 ) , .A2( us11_n744 ) , .A1( us11_n792 ) );
  NOR2_X1 us11_U243 (.ZN( us11_n507 ) , .A1( us11_n812 ) , .A2( us11_n817 ) );
  NOR2_X1 us11_U244 (.ZN( us11_n516 ) , .A1( us11_n708 ) , .A2( us11_n744 ) );
  NOR2_X1 us11_U245 (.ZN( us11_n558 ) , .A1( us11_n708 ) , .A2( us11_n816 ) );
  NOR2_X1 us11_U246 (.ZN( us11_n517 ) , .A1( us11_n708 ) , .A2( us11_n803 ) );
  INV_X1 us11_U247 (.A( us11_n806 ) , .ZN( us11_n841 ) );
  NOR2_X1 us11_U248 (.ZN( us11_n545 ) , .A1( us11_n749 ) , .A2( us11_n814 ) );
  INV_X1 us11_U249 (.A( us11_n728 ) , .ZN( us11_n852 ) );
  NOR4_X1 us11_U25 (.A4( us11_n532 ) , .A3( us11_n533 ) , .A2( us11_n534 ) , .ZN( us11_n535 ) , .A1( us11_n820 ) );
  NOR2_X1 us11_U250 (.ZN( us11_n554 ) , .A1( us11_n786 ) , .A2( us11_n813 ) );
  NOR2_X1 us11_U251 (.ZN( us11_n670 ) , .A1( us11_n790 ) , .A2( us11_n805 ) );
  NOR2_X1 us11_U252 (.ZN( us11_n717 ) , .A2( us11_n744 ) , .A1( us11_n786 ) );
  NOR2_X1 us11_U253 (.ZN( us11_n506 ) , .A2( us11_n728 ) , .A1( us11_n762 ) );
  NOR2_X1 us11_U254 (.ZN( us11_n642 ) , .A2( us11_n788 ) , .A1( us11_n791 ) );
  NOR2_X1 us11_U255 (.ZN( us11_n614 ) , .A1( us11_n762 ) , .A2( us11_n812 ) );
  AOI21_X1 us11_U256 (.ZN( us11_n626 ) , .B2( us11_n669 ) , .A( us11_n790 ) , .B1( us11_n791 ) );
  AOI21_X1 us11_U257 (.ZN( us11_n552 ) , .B1( us11_n669 ) , .A( us11_n697 ) , .B2( us11_n805 ) );
  AOI21_X1 us11_U258 (.ZN( us11_n589 ) , .B2( us11_n699 ) , .B1( us11_n815 ) , .A( us11_n817 ) );
  INV_X1 us11_U259 (.A( us11_n763 ) , .ZN( us11_n866 ) );
  NOR4_X1 us11_U26 (.ZN( us11_n456 ) , .A2( us11_n517 ) , .A1( us11_n543 ) , .A3( us11_n579 ) , .A4( us11_n615 ) );
  NOR2_X1 us11_U260 (.ZN( us11_n609 ) , .A2( us11_n724 ) , .A1( us11_n817 ) );
  NOR2_X1 us11_U261 (.ZN( us11_n668 ) , .A2( us11_n708 ) , .A1( us11_n790 ) );
  NOR2_X1 us11_U262 (.ZN( us11_n533 ) , .A2( us11_n724 ) , .A1( us11_n730 ) );
  NOR2_X1 us11_U263 (.ZN( us11_n521 ) , .A1( us11_n790 ) , .A2( us11_n812 ) );
  AOI21_X1 us11_U264 (.A( us11_n815 ) , .B2( us11_n816 ) , .B1( us11_n817 ) , .ZN( us11_n818 ) );
  NOR2_X1 us11_U265 (.ZN( us11_n547 ) , .A1( us11_n699 ) , .A2( us11_n744 ) );
  AOI21_X1 us11_U266 (.ZN( us11_n510 ) , .B2( us11_n669 ) , .A( us11_n730 ) , .B1( us11_n815 ) );
  NOR2_X1 us11_U267 (.ZN( us11_n655 ) , .A1( us11_n790 ) , .A2( us11_n815 ) );
  NOR2_X1 us11_U268 (.ZN( us11_n579 ) , .A2( us11_n708 ) , .A1( us11_n730 ) );
  INV_X1 us11_U269 (.A( us11_n729 ) , .ZN( us11_n868 ) );
  NOR4_X1 us11_U27 (.A4( us11_n577 ) , .A3( us11_n578 ) , .A2( us11_n579 ) , .ZN( us11_n586 ) , .A1( us11_n683 ) );
  NOR2_X1 us11_U270 (.ZN( us11_n542 ) , .A1( us11_n762 ) , .A2( us11_n791 ) );
  NOR2_X1 us11_U271 (.ZN( us11_n701 ) , .A2( us11_n786 ) , .A1( us11_n817 ) );
  NOR2_X1 us11_U272 (.A2( us11_n708 ) , .A1( us11_n762 ) , .ZN( us11_n794 ) );
  AOI21_X1 us11_U273 (.ZN( us11_n499 ) , .B1( us11_n680 ) , .A( us11_n812 ) , .B2( us11_n816 ) );
  AOI21_X1 us11_U274 (.ZN( us11_n650 ) , .A( us11_n779 ) , .B1( us11_n792 ) , .B2( us11_n805 ) );
  INV_X1 us11_U275 (.A( us11_n699 ) , .ZN( us11_n853 ) );
  NOR2_X1 us11_U276 (.ZN( us11_n652 ) , .A1( us11_n669 ) , .A2( us11_n814 ) );
  NOR2_X1 us11_U277 (.ZN( us11_n581 ) , .A1( us11_n669 ) , .A2( us11_n788 ) );
  AOI21_X1 us11_U278 (.ZN( us11_n515 ) , .A( us11_n729 ) , .B1( us11_n750 ) , .B2( us11_n803 ) );
  AOI21_X1 us11_U279 (.B1( us11_n699 ) , .ZN( us11_n700 ) , .A( us11_n732 ) , .B2( us11_n763 ) );
  AOI222_X1 us11_U28 (.B2( us11_n638 ) , .ZN( us11_n644 ) , .B1( us11_n841 ) , .A1( us11_n842 ) , .C2( us11_n846 ) , .C1( us11_n863 ) , .A2( us11_n865 ) );
  AOI21_X1 us11_U280 (.ZN( us11_n591 ) , .B2( us11_n763 ) , .A( us11_n785 ) , .B1( us11_n812 ) );
  AOI21_X1 us11_U281 (.A( us11_n812 ) , .B2( us11_n813 ) , .B1( us11_n814 ) , .ZN( us11_n819 ) );
  NOR2_X1 us11_U282 (.A1( us11_n730 ) , .ZN( us11_n765 ) , .A2( us11_n786 ) );
  INV_X1 us11_U283 (.A( us11_n791 ) , .ZN( us11_n873 ) );
  AOI21_X1 us11_U284 (.ZN( us11_n593 ) , .B1( us11_n750 ) , .A( us11_n792 ) , .B2( us11_n813 ) );
  NOR2_X1 us11_U285 (.ZN( us11_n582 ) , .A1( us11_n744 ) , .A2( us11_n815 ) );
  NOR2_X1 us11_U286 (.ZN( us11_n519 ) , .A2( us11_n699 ) , .A1( us11_n816 ) );
  NOR2_X1 us11_U287 (.ZN( us11_n685 ) , .A1( us11_n729 ) , .A2( us11_n816 ) );
  NOR2_X1 us11_U288 (.ZN( us11_n559 ) , .A2( us11_n791 ) , .A1( us11_n803 ) );
  AOI21_X1 us11_U289 (.ZN( us11_n649 ) , .B1( us11_n729 ) , .B2( us11_n763 ) , .A( us11_n813 ) );
  NOR4_X1 us11_U29 (.A4( us11_n639 ) , .A3( us11_n640 ) , .A2( us11_n641 ) , .A1( us11_n642 ) , .ZN( us11_n643 ) );
  AOI21_X1 us11_U290 (.B1( us11_n625 ) , .ZN( us11_n627 ) , .A( us11_n763 ) , .B2( us11_n814 ) );
  NOR2_X1 us11_U291 (.ZN( us11_n683 ) , .A2( us11_n699 ) , .A1( us11_n803 ) );
  NOR2_X1 us11_U292 (.A2( us11_n697 ) , .A1( us11_n780 ) , .ZN( us11_n820 ) );
  NOR2_X1 us11_U293 (.ZN( us11_n653 ) , .A1( us11_n762 ) , .A2( us11_n786 ) );
  NOR2_X1 us11_U294 (.ZN( us11_n568 ) , .A1( us11_n729 ) , .A2( us11_n762 ) );
  NOR2_X1 us11_U295 (.ZN( us11_n662 ) , .A2( us11_n697 ) , .A1( us11_n729 ) );
  INV_X1 us11_U296 (.A( us11_n813 ) , .ZN( us11_n836 ) );
  NOR2_X1 us11_U297 (.ZN( us11_n566 ) , .A2( us11_n697 ) , .A1( us11_n763 ) );
  NOR2_X1 us11_U298 (.ZN( us11_n520 ) , .A2( us11_n708 ) , .A1( us11_n814 ) );
  AOI21_X1 us11_U299 (.ZN( us11_n477 ) , .A( us11_n669 ) , .B1( us11_n750 ) , .B2( us11_n806 ) );
  NAND2_X2 us11_U3 (.A2( us11_n460 ) , .A1( us11_n465 ) , .ZN( us11_n780 ) );
  NOR3_X1 us11_U30 (.A2( us11_n607 ) , .A1( us11_n608 ) , .ZN( us11_n646 ) , .A3( us11_n722 ) );
  NOR2_X1 us11_U300 (.A1( us11_n697 ) , .ZN( us11_n770 ) , .A2( us11_n815 ) );
  AOI21_X1 us11_U301 (.ZN( us11_n514 ) , .A( us11_n779 ) , .B2( us11_n792 ) , .B1( us11_n812 ) );
  INV_X1 us11_U302 (.A( us11_n786 ) , .ZN( us11_n862 ) );
  AOI21_X1 us11_U303 (.ZN( us11_n540 ) , .A( us11_n763 ) , .B2( us11_n779 ) , .B1( us11_n817 ) );
  AOI21_X1 us11_U304 (.ZN( us11_n450 ) , .B2( us11_n792 ) , .A( us11_n803 ) , .B1( us11_n815 ) );
  AOI21_X1 us11_U305 (.ZN( us11_n539 ) , .B2( us11_n812 ) , .A( us11_n814 ) , .B1( us11_n815 ) );
  NOR2_X1 us11_U306 (.ZN( us11_n529 ) , .A1( us11_n708 ) , .A2( us11_n779 ) );
  NOR2_X1 us11_U307 (.ZN( us11_n578 ) , .A1( us11_n708 ) , .A2( us11_n813 ) );
  NOR2_X1 us11_U308 (.ZN( us11_n583 ) , .A1( us11_n792 ) , .A2( us11_n817 ) );
  NOR2_X1 us11_U309 (.ZN( us11_n534 ) , .A1( us11_n724 ) , .A2( us11_n788 ) );
  NOR4_X1 us11_U31 (.A4( us11_n541 ) , .A3( us11_n542 ) , .A2( us11_n543 ) , .ZN( us11_n550 ) , .A1( us11_n688 ) );
  NOR2_X1 us11_U310 (.ZN( us11_n632 ) , .A2( us11_n697 ) , .A1( us11_n724 ) );
  AOI21_X1 us11_U311 (.ZN( us11_n498 ) , .A( us11_n724 ) , .B2( us11_n762 ) , .B1( us11_n814 ) );
  AOI21_X1 us11_U312 (.A( us11_n790 ) , .B2( us11_n791 ) , .B1( us11_n792 ) , .ZN( us11_n793 ) );
  AOI21_X1 us11_U313 (.ZN( us11_n689 ) , .B2( us11_n749 ) , .B1( us11_n763 ) , .A( us11_n806 ) );
  AOI21_X1 us11_U314 (.B1( us11_n686 ) , .ZN( us11_n687 ) , .A( us11_n728 ) , .B2( us11_n761 ) );
  AOI21_X1 us11_U315 (.ZN( us11_n569 ) , .B1( us11_n750 ) , .B2( us11_n762 ) , .A( us11_n780 ) );
  AOI21_X1 us11_U316 (.ZN( us11_n500 ) , .A( us11_n697 ) , .B1( us11_n708 ) , .B2( us11_n786 ) );
  NOR2_X1 us11_U317 (.ZN( us11_n665 ) , .A1( us11_n780 ) , .A2( us11_n813 ) );
  NOR2_X1 us11_U318 (.ZN( us11_n580 ) , .A2( us11_n697 ) , .A1( us11_n791 ) );
  AOI21_X1 us11_U319 (.ZN( us11_n571 ) , .B2( us11_n697 ) , .B1( us11_n806 ) , .A( us11_n812 ) );
  AOI221_X1 us11_U32 (.A( us11_n713 ) , .B2( us11_n714 ) , .ZN( us11_n720 ) , .C1( us11_n832 ) , .B1( us11_n839 ) , .C2( us11_n863 ) );
  NOR2_X1 us11_U320 (.ZN( us11_n684 ) , .A1( us11_n791 ) , .A2( us11_n813 ) );
  AOI21_X1 us11_U321 (.ZN( us11_n639 ) , .B2( us11_n749 ) , .A( us11_n788 ) , .B1( us11_n812 ) );
  AOI21_X1 us11_U322 (.A( us11_n733 ) , .ZN( us11_n734 ) , .B2( us11_n780 ) , .B1( us11_n792 ) );
  NAND2_X2 us11_U323 (.A1( us11_n452 ) , .A2( us11_n465 ) , .ZN( us11_n669 ) );
  NOR2_X1 us11_U324 (.ZN( us11_n711 ) , .A1( us11_n762 ) , .A2( us11_n763 ) );
  AOI21_X1 us11_U325 (.ZN( us11_n478 ) , .B2( us11_n697 ) , .A( us11_n749 ) , .B1( us11_n779 ) );
  NOR2_X1 us11_U326 (.A2( us11_n813 ) , .A1( us11_n815 ) , .ZN( us11_n821 ) );
  NOR2_X1 us11_U327 (.A1( us11_n749 ) , .ZN( us11_n767 ) , .A2( us11_n803 ) );
  NOR2_X1 us11_U328 (.ZN( us11_n682 ) , .A2( us11_n708 ) , .A1( us11_n817 ) );
  NAND2_X2 us11_U329 (.A1( us11_n451 ) , .A2( us11_n471 ) , .ZN( us11_n816 ) );
  OR2_X1 us11_U33 (.A2( us11_n711 ) , .A1( us11_n712 ) , .ZN( us11_n713 ) );
  AOI21_X1 us11_U330 (.ZN( us11_n641 ) , .B1( us11_n680 ) , .A( us11_n791 ) , .B2( us11_n817 ) );
  NAND2_X1 us11_U331 (.ZN( us11_n753 ) , .A1( us11_n763 ) , .A2( us11_n805 ) );
  OAI21_X1 us11_U332 (.A( us11_n731 ) , .B1( us11_n732 ) , .ZN( us11_n736 ) , .B2( us11_n805 ) );
  OAI21_X1 us11_U333 (.ZN( us11_n731 ) , .A( us11_n833 ) , .B2( us11_n852 ) , .B1( us11_n873 ) );
  INV_X1 us11_U334 (.A( us11_n815 ) , .ZN( us11_n855 ) );
  NAND2_X2 us11_U335 (.A1( us11_n447 ) , .A2( us11_n449 ) , .ZN( us11_n805 ) );
  NAND2_X2 us11_U336 (.A2( us11_n449 ) , .A1( us11_n452 ) , .ZN( us11_n763 ) );
  AOI21_X1 us11_U337 (.ZN( us11_n442 ) , .A( us11_n699 ) , .B1( us11_n733 ) , .B2( us11_n750 ) );
  OAI21_X1 us11_U338 (.A( us11_n698 ) , .ZN( us11_n702 ) , .B2( us11_n750 ) , .B1( us11_n804 ) );
  OAI21_X1 us11_U339 (.ZN( us11_n698 ) , .B2( us11_n833 ) , .B1( us11_n838 ) , .A( us11_n860 ) );
  NOR2_X1 us11_U34 (.ZN( us11_n680 ) , .A2( us11_n834 ) , .A1( us11_n839 ) );
  NAND2_X1 us11_U340 (.A1( us11_n699 ) , .A2( us11_n729 ) , .ZN( us11_n782 ) );
  NOR2_X1 us11_U341 (.ZN( us11_n526 ) , .A1( us11_n724 ) , .A2( us11_n750 ) );
  INV_X1 us11_U342 (.A( us11_n780 ) , .ZN( us11_n850 ) );
  NOR2_X1 us11_U343 (.ZN( us11_n518 ) , .A1( us11_n708 ) , .A2( us11_n788 ) );
  AOI21_X1 us11_U344 (.ZN( us11_n443 ) , .B1( us11_n789 ) , .B2( us11_n791 ) , .A( us11_n814 ) );
  AOI21_X1 us11_U345 (.ZN( us11_n497 ) , .A( us11_n779 ) , .B2( us11_n791 ) , .B1( us11_n804 ) );
  NAND2_X2 us11_U346 (.A2( us11_n441 ) , .A1( us11_n447 ) , .ZN( us11_n784 ) );
  NAND2_X1 us11_U347 (.ZN( us11_n714 ) , .A1( us11_n728 ) , .A2( us11_n780 ) );
  NOR2_X1 us11_U348 (.ZN( us11_n484 ) , .A1( us11_n788 ) , .A2( us11_n805 ) );
  OAI21_X1 us11_U349 (.A( us11_n787 ) , .B2( us11_n788 ) , .B1( us11_n789 ) , .ZN( us11_n795 ) );
  AOI222_X1 us11_U35 (.ZN( us11_n469 ) , .B1( us11_n832 ) , .A1( us11_n839 ) , .C1( us11_n842 ) , .C2( us11_n851 ) , .A2( us11_n855 ) , .B2( us11_n865 ) );
  NAND2_X2 us11_U350 (.A2( us11_n448 ) , .A1( us11_n452 ) , .ZN( us11_n729 ) );
  OAI21_X1 us11_U351 (.ZN( us11_n787 ) , .A( us11_n839 ) , .B1( us11_n863 ) , .B2( us11_n873 ) );
  NAND2_X1 us11_U352 (.A2( us11_n762 ) , .A1( us11_n806 ) , .ZN( us11_n810 ) );
  INV_X1 us11_U353 (.A( us11_n785 ) , .ZN( us11_n846 ) );
  NOR2_X1 us11_U354 (.ZN( us11_n470 ) , .A2( us11_n779 ) , .A1( us11_n815 ) );
  NOR2_X1 us11_U355 (.ZN( us11_n712 ) , .A2( us11_n724 ) , .A1( us11_n790 ) );
  NAND2_X1 us11_U356 (.ZN( us11_n671 ) , .A1( us11_n806 ) , .A2( us11_n816 ) );
  NAND2_X1 us11_U357 (.A2( us11_n749 ) , .A1( us11_n786 ) , .ZN( us11_n809 ) );
  INV_X1 us11_U358 (.A( us11_n724 ) , .ZN( us11_n856 ) );
  INV_X1 us11_U359 (.A( us11_n817 ) , .ZN( us11_n844 ) );
  NOR4_X1 us11_U36 (.A1( us11_n466 ) , .ZN( us11_n467 ) , .A4( us11_n542 ) , .A2( us11_n554 ) , .A3( us11_n614 ) );
  AND2_X1 us11_U360 (.ZN( us11_n732 ) , .A1( us11_n779 ) , .A2( us11_n785 ) );
  AOI221_X1 us11_U361 (.A( us11_n764 ) , .ZN( us11_n774 ) , .C2( us11_n810 ) , .B2( us11_n835 ) , .C1( us11_n855 ) , .B1( us11_n866 ) );
  AOI21_X1 us11_U362 (.B2( us11_n763 ) , .ZN( us11_n764 ) , .A( us11_n788 ) , .B1( us11_n792 ) );
  INV_X1 us11_U363 (.A( us11_n761 ) , .ZN( us11_n835 ) );
  NAND2_X1 us11_U364 (.A2( us11_n448 ) , .A1( us11_n460 ) , .ZN( us11_n728 ) );
  NAND2_X1 us11_U365 (.A1( us11_n451 ) , .A2( us11_n454 ) , .ZN( us11_n814 ) );
  NAND2_X1 us11_U366 (.A1( us11_n455 ) , .A2( us11_n462 ) , .ZN( us11_n750 ) );
  NAND2_X1 us11_U367 (.A2( us11_n454 ) , .A1( us11_n472 ) , .ZN( us11_n779 ) );
  NAND2_X1 us11_U368 (.A2( us11_n453 ) , .A1( us11_n455 ) , .ZN( us11_n806 ) );
  NAND2_X1 us11_U369 (.A1( us11_n453 ) , .A2( us11_n472 ) , .ZN( us11_n785 ) );
  AOI221_X1 us11_U37 (.ZN( us11_n468 ) , .C2( us11_n714 ) , .B2( us11_n831 ) , .C1( us11_n845 ) , .B1( us11_n860 ) , .A( us11_n864 ) );
  NAND2_X1 us11_U370 (.A2( us11_n464 ) , .A1( us11_n465 ) , .ZN( us11_n812 ) );
  NAND2_X1 us11_U371 (.A1( us11_n447 ) , .A2( us11_n448 ) , .ZN( us11_n786 ) );
  NAND2_X2 us11_U372 (.A1( us11_n455 ) , .A2( us11_n471 ) , .ZN( us11_n803 ) );
  NAND2_X1 us11_U373 (.A1( us11_n462 ) , .A2( us11_n472 ) , .ZN( us11_n788 ) );
  NOR2_X1 us11_U374 (.ZN( us11_n465 ) , .A2( us11_n847 ) , .A1( us11_n848 ) );
  NAND2_X2 us11_U375 (.A1( us11_n453 ) , .A2( us11_n461 ) , .ZN( us11_n744 ) );
  NOR2_X1 us11_U376 (.ZN( us11_n453 ) , .A1( us11_n826 ) , .A2( us11_n827 ) );
  NOR2_X1 us11_U377 (.ZN( us11_n451 ) , .A1( us11_n828 ) , .A2( us11_n829 ) );
  NAND2_X1 us11_U378 (.A2( us11_n454 ) , .A1( us11_n455 ) , .ZN( us11_n730 ) );
  NAND2_X1 us11_U379 (.A1( us11_n451 ) , .A2( us11_n462 ) , .ZN( us11_n790 ) );
  NOR4_X1 us11_U38 (.A4( us11_n514 ) , .A3( us11_n515 ) , .A2( us11_n516 ) , .A1( us11_n517 ) , .ZN( us11_n524 ) );
  NAND2_X2 us11_U380 (.A1( us11_n449 ) , .A2( us11_n460 ) , .ZN( us11_n792 ) );
  NAND2_X2 us11_U381 (.A2( us11_n448 ) , .A1( us11_n464 ) , .ZN( us11_n815 ) );
  NAND2_X2 us11_U382 (.A2( us11_n471 ) , .A1( us11_n472 ) , .ZN( us11_n817 ) );
  NAND2_X2 us11_U383 (.A1( us11_n441 ) , .A2( us11_n460 ) , .ZN( us11_n699 ) );
  NOR2_X1 us11_U384 (.ZN( us11_n447 ) , .A2( us11_n849 ) , .A1( us11_n858 ) );
  NOR2_X1 us11_U385 (.A2( sa11_6 ) , .A1( sa11_7 ) , .ZN( us11_n464 ) );
  NOR2_X1 us11_U386 (.A2( sa11_7 ) , .ZN( us11_n460 ) , .A1( us11_n849 ) );
  NOR2_X1 us11_U387 (.A2( sa11_5 ) , .ZN( us11_n448 ) , .A1( us11_n847 ) );
  NOR2_X1 us11_U388 (.A2( sa11_2 ) , .A1( sa11_3 ) , .ZN( us11_n472 ) );
  NOR2_X1 us11_U389 (.A2( sa11_0 ) , .ZN( us11_n454 ) , .A1( us11_n827 ) );
  AOI222_X1 us11_U39 (.ZN( us11_n525 ) , .A1( us11_n834 ) , .B2( us11_n837 ) , .C1( us11_n844 ) , .C2( us11_n850 ) , .A2( us11_n852 ) , .B1( us11_n866 ) );
  NOR2_X1 us11_U390 (.A2( sa11_3 ) , .ZN( us11_n455 ) , .A1( us11_n828 ) );
  NOR2_X1 us11_U391 (.A2( sa11_0 ) , .A1( sa11_1 ) , .ZN( us11_n462 ) );
  INV_X1 us11_U392 (.A( sa11_6 ) , .ZN( us11_n849 ) );
  INV_X1 us11_U393 (.A( sa11_1 ) , .ZN( us11_n827 ) );
  INV_X1 us11_U394 (.A( sa11_2 ) , .ZN( us11_n828 ) );
  INV_X1 us11_U395 (.A( sa11_5 ) , .ZN( us11_n848 ) );
  NAND2_X1 us11_U396 (.A2( us11_n461 ) , .A1( us11_n471 ) , .ZN( us11_n697 ) );
  NOR2_X1 us11_U397 (.A2( sa11_6 ) , .ZN( us11_n452 ) , .A1( us11_n858 ) );
  INV_X1 us11_U398 (.A( sa11_7 ) , .ZN( us11_n858 ) );
  NAND2_X1 us11_U399 (.A2( us11_n461 ) , .A1( us11_n462 ) , .ZN( us11_n747 ) );
  NAND2_X2 us11_U4 (.A1( us11_n441 ) , .A2( us11_n464 ) , .ZN( us11_n708 ) );
  NOR4_X1 us11_U40 (.A3( us11_n521 ) , .A1( us11_n522 ) , .ZN( us11_n523 ) , .A2( us11_n673 ) , .A4( us11_n769 ) );
  NAND2_X2 us11_U400 (.A1( us11_n454 ) , .A2( us11_n461 ) , .ZN( us11_n813 ) );
  NOR2_X1 us11_U401 (.A2( sa11_1 ) , .ZN( us11_n471 ) , .A1( us11_n826 ) );
  INV_X1 us11_U402 (.A( sa11_0 ) , .ZN( us11_n826 ) );
  OAI221_X1 us11_U403 (.A( us11_n783 ) , .C2( us11_n784 ) , .B2( us11_n785 ) , .B1( us11_n786 ) , .ZN( us11_n796 ) , .C1( us11_n813 ) );
  NAND2_X1 us11_U404 (.A1( us11_n729 ) , .A2( us11_n784 ) , .ZN( us11_n811 ) );
  OAI22_X1 us11_U405 (.ZN( us11_n588 ) , .A2( us11_n747 ) , .B2( us11_n762 ) , .A1( us11_n763 ) , .B1( us11_n784 ) );
  OAI221_X1 us11_U406 (.A( us11_n696 ) , .ZN( us11_n703 ) , .C2( us11_n784 ) , .C1( us11_n785 ) , .B1( us11_n786 ) , .B2( us11_n806 ) );
  AOI21_X1 us11_U407 (.ZN( us11_n592 ) , .B1( us11_n728 ) , .B2( us11_n784 ) , .A( us11_n790 ) );
  AOI21_X1 us11_U408 (.ZN( us11_n648 ) , .A( us11_n762 ) , .B2( us11_n784 ) , .B1( us11_n792 ) );
  AOI21_X1 us11_U409 (.ZN( us11_n623 ) , .B1( us11_n699 ) , .A( us11_n779 ) , .B2( us11_n784 ) );
  AOI221_X1 us11_U41 (.A( us11_n781 ) , .ZN( us11_n798 ) , .C2( us11_n837 ) , .B2( us11_n838 ) , .B1( us11_n865 ) , .C1( us11_n866 ) );
  OAI22_X1 us11_U410 (.ZN( us11_n681 ) , .A1( us11_n699 ) , .A2( us11_n730 ) , .B2( us11_n784 ) , .B1( us11_n817 ) );
  OAI21_X1 us11_U411 (.A( us11_n613 ) , .ZN( us11_n616 ) , .B1( us11_n625 ) , .B2( us11_n784 ) );
  NOR2_X1 us11_U412 (.ZN( us11_n610 ) , .A1( us11_n784 ) , .A2( us11_n816 ) );
  NOR2_X1 us11_U413 (.ZN( us11_n651 ) , .A1( us11_n784 ) , .A2( us11_n788 ) );
  OAI222_X1 us11_U414 (.A2( us11_n669 ) , .ZN( us11_n674 ) , .B1( us11_n747 ) , .B2( us11_n784 ) , .C2( us11_n788 ) , .C1( us11_n815 ) , .A1( us11_n817 ) );
  NOR2_X1 us11_U415 (.ZN( us11_n600 ) , .A2( us11_n697 ) , .A1( us11_n784 ) );
  NOR2_X1 us11_U416 (.ZN( us11_n553 ) , .A2( us11_n744 ) , .A1( us11_n784 ) );
  INV_X1 us11_U417 (.A( us11_n784 ) , .ZN( us11_n861 ) );
  NAND4_X1 us11_U418 (.ZN( sa10_sr_2 ) , .A4( us11_n643 ) , .A3( us11_n644 ) , .A2( us11_n645 ) , .A1( us11_n646 ) );
  AOI211_X1 us11_U419 (.A( us11_n637 ) , .ZN( us11_n645 ) , .B( us11_n743 ) , .C2( us11_n839 ) , .C1( us11_n854 ) );
  NOR4_X1 us11_U42 (.A4( us11_n793 ) , .A3( us11_n794 ) , .A2( us11_n795 ) , .A1( us11_n796 ) , .ZN( us11_n797 ) );
  NOR4_X1 us11_U420 (.A1( us11_n584 ) , .ZN( us11_n585 ) , .A3( us11_n652 ) , .A2( us11_n662 ) , .A4( us11_n767 ) );
  NOR2_X1 us11_U421 (.A2( sa11_2 ) , .ZN( us11_n461 ) , .A1( us11_n829 ) );
  INV_X1 us11_U422 (.A( sa11_3 ) , .ZN( us11_n829 ) );
  OAI222_X1 us11_U423 (.B2( us11_n747 ) , .B1( us11_n748 ) , .A2( us11_n749 ) , .ZN( us11_n757 ) , .C2( us11_n805 ) , .C1( us11_n814 ) , .A1( us11_n817 ) );
  OAI222_X1 us11_U424 (.ZN( us11_n505 ) , .C2( us11_n625 ) , .B2( us11_n647 ) , .B1( us11_n747 ) , .A2( us11_n748 ) , .C1( us11_n805 ) , .A1( us11_n806 ) );
  AOI222_X1 us11_U425 (.ZN( us11_n605 ) , .B2( us11_n671 ) , .B1( us11_n753 ) , .C2( us11_n831 ) , .A1( us11_n833 ) , .A2( us11_n862 ) , .C1( us11_n863 ) );
  AOI222_X1 us11_U426 (.ZN( us11_n513 ) , .C1( us11_n832 ) , .B2( us11_n837 ) , .A2( us11_n843 ) , .C2( us11_n862 ) , .B1( us11_n863 ) , .A1( us11_n866 ) );
  AOI221_X1 us11_U427 (.A( us11_n483 ) , .ZN( us11_n488 ) , .B1( us11_n831 ) , .C2( us11_n844 ) , .C1( us11_n852 ) , .B2( us11_n862 ) );
  NOR2_X1 us11_U428 (.ZN( us11_n789 ) , .A2( us11_n862 ) , .A1( us11_n868 ) );
  NOR2_X1 us11_U429 (.ZN( us11_n748 ) , .A1( us11_n861 ) , .A2( us11_n862 ) );
  NOR4_X1 us11_U43 (.A4( us11_n776 ) , .A3( us11_n777 ) , .A1( us11_n778 ) , .ZN( us11_n799 ) , .A2( us11_n801 ) );
  NOR2_X1 us11_U430 (.A2( sa11_4 ) , .ZN( us11_n449 ) , .A1( us11_n848 ) );
  NOR2_X1 us11_U431 (.A2( sa11_4 ) , .A1( sa11_5 ) , .ZN( us11_n441 ) );
  INV_X1 us11_U432 (.A( sa11_4 ) , .ZN( us11_n847 ) );
  AND2_X1 us11_U433 (.ZN( us11_n438 ) , .A2( us11_n831 ) , .A1( us11_n854 ) );
  AND2_X1 us11_U434 (.ZN( us11_n439 ) , .A2( us11_n843 ) , .A1( us11_n861 ) );
  NOR3_X1 us11_U435 (.A1( us11_n438 ) , .A2( us11_n439 ) , .A3( us11_n576 ) , .ZN( us11_n587 ) );
  INV_X1 us11_U436 (.A( us11_n812 ) , .ZN( us11_n854 ) );
  NAND3_X1 us11_U437 (.ZN( sa10_sr_6 ) , .A3( us11_n797 ) , .A2( us11_n798 ) , .A1( us11_n799 ) );
  NAND3_X1 us11_U438 (.ZN( sa10_sr_5 ) , .A3( us11_n758 ) , .A2( us11_n759 ) , .A1( us11_n760 ) );
  NAND3_X1 us11_U439 (.ZN( sa10_sr_4 ) , .A3( us11_n738 ) , .A2( us11_n739 ) , .A1( us11_n740 ) );
  NOR4_X1 us11_U44 (.A4( us11_n734 ) , .A3( us11_n735 ) , .A2( us11_n736 ) , .A1( us11_n737 ) , .ZN( us11_n738 ) );
  NAND3_X1 us11_U440 (.A3( us11_n675 ) , .A2( us11_n676 ) , .A1( us11_n677 ) , .ZN( us11_n807 ) );
  NAND3_X1 us11_U441 (.ZN( us11_n638 ) , .A3( us11_n708 ) , .A2( us11_n724 ) , .A1( us11_n792 ) );
  NAND3_X1 us11_U442 (.A3( us11_n618 ) , .A2( us11_n619 ) , .A1( us11_n620 ) , .ZN( us11_n725 ) );
  NAND3_X1 us11_U443 (.A3( us11_n585 ) , .A2( us11_n586 ) , .A1( us11_n587 ) , .ZN( us11_n621 ) );
  NAND3_X1 us11_U444 (.ZN( us11_n565 ) , .A3( us11_n680 ) , .A2( us11_n750 ) , .A1( us11_n785 ) );
  NAND3_X1 us11_U445 (.A3( us11_n523 ) , .A2( us11_n524 ) , .A1( us11_n525 ) , .ZN( us11_n742 ) );
  NAND3_X1 us11_U446 (.A3( us11_n512 ) , .A1( us11_n513 ) , .ZN( us11_n608 ) , .A2( us11_n871 ) );
  NAND3_X1 us11_U447 (.A3( us11_n467 ) , .A2( us11_n468 ) , .A1( us11_n469 ) , .ZN( us11_n777 ) );
  INV_X1 us11_U448 (.A( us11_n803 ) , .ZN( us11_n843 ) );
  AOI21_X1 us11_U449 (.ZN( us11_n576 ) , .B2( us11_n724 ) , .B1( us11_n748 ) , .A( us11_n785 ) );
  AOI211_X1 us11_U45 (.B( us11_n725 ) , .A( us11_n726 ) , .ZN( us11_n739 ) , .C1( us11_n843 ) , .C2( us11_n855 ) );
  NOR3_X1 us11_U46 (.A3( us11_n722 ) , .A1( us11_n723 ) , .ZN( us11_n740 ) , .A2( us11_n741 ) );
  NOR4_X1 us11_U47 (.A3( us11_n755 ) , .A2( us11_n756 ) , .A1( us11_n757 ) , .ZN( us11_n758 ) , .A4( us11_n869 ) );
  AOI211_X1 us11_U48 (.B( us11_n745 ) , .A( us11_n746 ) , .ZN( us11_n759 ) , .C1( us11_n832 ) , .C2( us11_n853 ) );
  NOR3_X1 us11_U49 (.A3( us11_n741 ) , .A2( us11_n742 ) , .A1( us11_n743 ) , .ZN( us11_n760 ) );
  NAND2_X2 us11_U5 (.A2( us11_n441 ) , .A1( us11_n452 ) , .ZN( us11_n791 ) );
  NAND4_X1 us11_U50 (.ZN( sa10_sr_3 ) , .A4( us11_n704 ) , .A3( us11_n705 ) , .A2( us11_n706 ) , .A1( us11_n707 ) );
  NOR4_X1 us11_U51 (.A4( us11_n700 ) , .A3( us11_n701 ) , .A2( us11_n702 ) , .A1( us11_n703 ) , .ZN( us11_n704 ) );
  AOI211_X1 us11_U52 (.B( us11_n694 ) , .A( us11_n695 ) , .ZN( us11_n705 ) , .C2( us11_n831 ) , .C1( us11_n851 ) );
  NOR2_X1 us11_U53 (.ZN( us11_n707 ) , .A2( us11_n776 ) , .A1( us11_n800 ) );
  NOR2_X1 us11_U54 (.ZN( us11_n804 ) , .A1( us11_n854 ) , .A2( us11_n861 ) );
  NAND4_X1 us11_U55 (.ZN( sa10_sr_1 ) , .A4( us11_n595 ) , .A3( us11_n596 ) , .A2( us11_n597 ) , .A1( us11_n598 ) );
  AOI211_X1 us11_U56 (.B( us11_n589 ) , .A( us11_n590 ) , .ZN( us11_n596 ) , .C2( us11_n811 ) , .C1( us11_n833 ) );
  NOR4_X1 us11_U57 (.A4( us11_n591 ) , .A3( us11_n592 ) , .A2( us11_n593 ) , .A1( us11_n594 ) , .ZN( us11_n595 ) );
  AOI211_X1 us11_U58 (.A( us11_n588 ) , .ZN( us11_n597 ) , .B( us11_n621 ) , .C1( us11_n845 ) , .C2( us11_n855 ) );
  NAND4_X1 us11_U59 (.ZN( sa10_sr_0 ) , .A4( us11_n501 ) , .A3( us11_n502 ) , .A2( us11_n503 ) , .A1( us11_n504 ) );
  INV_X1 us11_U6 (.A( us11_n669 ) , .ZN( us11_n865 ) );
  AOI221_X1 us11_U60 (.A( us11_n497 ) , .ZN( us11_n502 ) , .B2( us11_n843 ) , .C1( us11_n846 ) , .C2( us11_n860 ) , .B1( us11_n862 ) );
  NOR4_X1 us11_U61 (.A4( us11_n498 ) , .A3( us11_n499 ) , .A2( us11_n500 ) , .ZN( us11_n501 ) , .A1( us11_n527 ) );
  AOI211_X1 us11_U62 (.A( us11_n496 ) , .ZN( us11_n503 ) , .B( us11_n802 ) , .C2( us11_n839 ) , .C1( us11_n851 ) );
  NAND4_X1 us11_U63 (.ZN( sa10_sr_7 ) , .A4( us11_n822 ) , .A3( us11_n823 ) , .A2( us11_n824 ) , .A1( us11_n825 ) );
  AOI222_X1 us11_U64 (.C2( us11_n809 ) , .B2( us11_n810 ) , .A2( us11_n811 ) , .ZN( us11_n823 ) , .C1( us11_n832 ) , .A1( us11_n839 ) , .B1( us11_n853 ) );
  NOR4_X1 us11_U65 (.A4( us11_n818 ) , .A3( us11_n819 ) , .A2( us11_n820 ) , .A1( us11_n821 ) , .ZN( us11_n822 ) );
  AOI211_X1 us11_U66 (.B( us11_n807 ) , .A( us11_n808 ) , .ZN( us11_n824 ) , .C1( us11_n842 ) , .C2( us11_n850 ) );
  NAND4_X1 us11_U67 (.A4( us11_n603 ) , .A3( us11_n604 ) , .A2( us11_n605 ) , .A1( us11_n606 ) , .ZN( us11_n722 ) );
  NOR3_X1 us11_U68 (.A1( us11_n599 ) , .ZN( us11_n604 ) , .A3( us11_n663 ) , .A2( us11_n770 ) );
  NOR4_X1 us11_U69 (.A3( us11_n600 ) , .A2( us11_n601 ) , .A1( us11_n602 ) , .ZN( us11_n603 ) , .A4( us11_n655 ) );
  NAND2_X1 us11_U7 (.A1( us11_n449 ) , .A2( us11_n464 ) , .ZN( us11_n724 ) );
  AOI222_X1 us11_U70 (.ZN( us11_n606 ) , .A1( us11_n830 ) , .C2( us11_n837 ) , .B1( us11_n842 ) , .A2( us11_n856 ) , .B2( us11_n861 ) , .C1( us11_n868 ) );
  NAND4_X1 us11_U71 (.A4( us11_n485 ) , .A3( us11_n486 ) , .A2( us11_n487 ) , .A1( us11_n488 ) , .ZN( us11_n778 ) );
  NOR4_X1 us11_U72 (.A4( us11_n484 ) , .ZN( us11_n487 ) , .A1( us11_n566 ) , .A2( us11_n581 ) , .A3( us11_n602 ) );
  NOR4_X1 us11_U73 (.ZN( us11_n486 ) , .A1( us11_n507 ) , .A2( us11_n519 ) , .A4( us11_n546 ) , .A3( us11_n611 ) );
  NAND4_X1 us11_U74 (.A4( us11_n657 ) , .A3( us11_n658 ) , .A2( us11_n659 ) , .A1( us11_n660 ) , .ZN( us11_n800 ) );
  NOR3_X1 us11_U75 (.A3( us11_n654 ) , .A2( us11_n655 ) , .A1( us11_n656 ) , .ZN( us11_n657 ) );
  NOR3_X1 us11_U76 (.A3( us11_n651 ) , .A2( us11_n652 ) , .A1( us11_n653 ) , .ZN( us11_n658 ) );
  NOR3_X1 us11_U77 (.A3( us11_n648 ) , .A2( us11_n649 ) , .A1( us11_n650 ) , .ZN( us11_n659 ) );
  NAND4_X1 us11_U78 (.A4( us11_n560 ) , .A3( us11_n561 ) , .A2( us11_n562 ) , .A1( us11_n563 ) , .ZN( us11_n607 ) );
  NOR4_X1 us11_U79 (.ZN( us11_n561 ) , .A1( us11_n653 ) , .A3( us11_n661 ) , .A4( us11_n685 ) , .A2( us11_n768 ) );
  NOR3_X1 us11_U8 (.ZN( us11_n598 ) , .A1( us11_n608 ) , .A3( us11_n723 ) , .A2( us11_n742 ) );
  NOR4_X1 us11_U80 (.A4( us11_n552 ) , .A3( us11_n553 ) , .A2( us11_n554 ) , .A1( us11_n555 ) , .ZN( us11_n562 ) );
  NOR4_X1 us11_U81 (.A4( us11_n556 ) , .A3( us11_n557 ) , .A2( us11_n558 ) , .A1( us11_n559 ) , .ZN( us11_n560 ) );
  NAND4_X1 us11_U82 (.A4( us11_n772 ) , .A3( us11_n773 ) , .A2( us11_n774 ) , .A1( us11_n775 ) , .ZN( us11_n801 ) );
  NOR3_X1 us11_U83 (.A3( us11_n765 ) , .A2( us11_n766 ) , .A1( us11_n767 ) , .ZN( us11_n773 ) );
  NOR4_X1 us11_U84 (.A4( us11_n768 ) , .A3( us11_n769 ) , .A2( us11_n770 ) , .A1( us11_n771 ) , .ZN( us11_n772 ) );
  AOI222_X1 us11_U85 (.ZN( us11_n775 ) , .A1( us11_n830 ) , .C1( us11_n834 ) , .B2( us11_n841 ) , .A2( us11_n850 ) , .B1( us11_n861 ) , .C2( us11_n873 ) );
  NOR4_X1 us11_U86 (.A4( us11_n509 ) , .A2( us11_n510 ) , .A1( us11_n511 ) , .ZN( us11_n512 ) , .A3( us11_n670 ) );
  INV_X1 us11_U87 (.A( us11_n505 ) , .ZN( us11_n871 ) );
  NOR4_X1 us11_U88 (.A4( us11_n665 ) , .A3( us11_n666 ) , .A2( us11_n667 ) , .A1( us11_n668 ) , .ZN( us11_n676 ) );
  NOR4_X1 us11_U89 (.A4( us11_n661 ) , .A3( us11_n662 ) , .A2( us11_n663 ) , .A1( us11_n664 ) , .ZN( us11_n677 ) );
  NOR3_X1 us11_U9 (.A3( us11_n800 ) , .A2( us11_n801 ) , .A1( us11_n802 ) , .ZN( us11_n825 ) );
  NOR4_X1 us11_U90 (.A3( us11_n673 ) , .A1( us11_n674 ) , .ZN( us11_n675 ) , .A4( us11_n715 ) , .A2( us11_n859 ) );
  NOR2_X1 us11_U91 (.ZN( us11_n625 ) , .A2( us11_n836 ) , .A1( us11_n839 ) );
  NOR2_X1 us11_U92 (.ZN( us11_n761 ) , .A1( us11_n833 ) , .A2( us11_n834 ) );
  NAND4_X1 us11_U93 (.A4( us11_n456 ) , .A3( us11_n457 ) , .A2( us11_n458 ) , .A1( us11_n459 ) , .ZN( us11_n679 ) );
  AOI221_X1 us11_U94 (.A( us11_n450 ) , .ZN( us11_n459 ) , .C2( us11_n753 ) , .B1( us11_n832 ) , .C1( us11_n842 ) , .B2( us11_n861 ) );
  NOR3_X1 us11_U95 (.ZN( us11_n457 ) , .A3( us11_n530 ) , .A1( us11_n555 ) , .A2( us11_n570 ) );
  NOR4_X1 us11_U96 (.ZN( us11_n458 ) , .A2( us11_n509 ) , .A1( us11_n599 ) , .A4( us11_n628 ) , .A3( us11_n711 ) );
  NAND4_X1 us11_U97 (.A4( us11_n535 ) , .A3( us11_n536 ) , .A2( us11_n537 ) , .A1( us11_n538 ) , .ZN( us11_n622 ) );
  NOR4_X1 us11_U98 (.A1( us11_n531 ) , .ZN( us11_n536 ) , .A2( us11_n654 ) , .A4( us11_n668 ) , .A3( us11_n765 ) );
  NOR4_X1 us11_U99 (.A4( us11_n526 ) , .A2( us11_n527 ) , .A1( us11_n528 ) , .ZN( us11_n538 ) , .A3( us11_n701 ) );
endmodule

