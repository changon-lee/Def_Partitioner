module aes_aes ( clk, key, ld, rst, text_in, done, text_out );
  input clk;
  input [127:0] key;
  input ld;
  input rst;
  input [127:0] text_in;
  output done;
  output [127:0] text_out;

  wire N100, N102, N105, N114, N116, N132, N133, N134, 
       N147, N148, N149, N150, N169, N227, N228, N229, N230, 
       N231, N233, N242, N244, N245, N246, N247, N258, N261, 
       N277, N278, N280, N35, N36, N37, N38, N40, N41, 
       N430, N434, N435, N436, N437, N438, N439, N440, N441, 
       N463, N52, N53, N54, N57, N66, N67, N68, N73, 
       N82, N83, N84, N85, N86, N87, N88, N89, N98, 
       N99, n101, n103, n105, n1109, n1114, n1145, n115, n117, 
       n1183, n119, n121, n1212, n1213, n1214, n1215, n1216, n1217, 
       n1219, n1220, n1221, n13, n143, n15, n195, n197, n199, 
       n201, n203, n207, n209, n21, n213, n215, n217, n219, 
       n225, n23, n231, n247, n249, n25, n253, n3, n31, 
       n33, n342, n348, n35, n354, n362, n37, n394, n396, 
       n414, n419, n433, n462, n469, n47, n481, n482, n49, 
       n5, n500, n506, n51, n515, n524, n53, n534, n547, 
       n55, n562, n57, n59, n590, n61, n63, n636, n65, 
       n657, n665, n67, n69, n7, n73, n786, n79, n791, 
       n81, n817, n823, n830, n85, n861, n870, n9, n900, 
       n905, n911, n917, n923, n927, n937, n957, sa00_0, sa00_1, 
       sa00_2, sa00_3, sa00_4, sa00_5, sa00_6, sa00_7, sa00_sr_0, sa00_sr_1, sa00_sr_2, 
       sa00_sr_3, sa00_sr_4, sa00_sr_5, sa00_sr_6, sa00_sr_7, sa01_0, sa01_1, sa01_2, sa01_3, 
       sa01_4, sa01_5, sa01_6, sa01_7, sa01_sr_0, sa01_sr_1, sa01_sr_2, sa01_sr_3, sa01_sr_4, 
       sa01_sr_5, sa01_sr_6, sa01_sr_7, sa02_0, sa02_1, sa02_2, sa02_3, sa02_4, sa02_5, 
       sa02_6, sa02_7, sa02_sr_0, sa02_sr_1, sa02_sr_2, sa02_sr_3, sa02_sr_4, sa02_sr_5, sa02_sr_6, 
       sa02_sr_7, sa03_0, sa03_1, sa03_2, sa03_3, sa03_4, sa03_5, sa03_6, sa03_7, 
       sa03_sr_0, sa03_sr_1, sa03_sr_2, sa03_sr_3, sa03_sr_4, sa03_sr_5, sa03_sr_6, sa03_sr_7, sa10_0, 
       sa10_1, sa10_2, sa10_3, sa10_4, sa10_5, sa10_6, sa10_7, sa10_sr_0, sa10_sr_1, 
       sa10_sr_2, sa10_sr_3, sa10_sr_4, sa10_sr_5, sa10_sr_6, sa10_sr_7, sa11_0, sa11_1, sa11_2, 
       sa11_3, sa11_4, sa11_5, sa11_6, sa11_7, sa11_sr_0, sa11_sr_1, sa11_sr_2, sa11_sr_3, 
       sa11_sr_4, sa11_sr_5, sa11_sr_6, sa11_sr_7, sa12_0, sa12_1, sa12_2, sa12_3, sa12_4, 
       sa12_5, sa12_6, sa12_7, sa12_sr_0, sa12_sr_1, sa12_sr_2, sa12_sr_3, sa12_sr_4, sa12_sr_5, 
       sa12_sr_6, sa12_sr_7, sa13_0, sa13_1, sa13_2, sa13_3, sa13_4, sa13_5, sa13_6, 
       sa13_7, sa20_0, sa20_1, sa20_2, sa20_3, sa20_4, sa20_5, sa20_6, sa20_7, 
       sa20_sr_0, sa20_sr_1, sa20_sr_2, sa20_sr_3, sa20_sr_4, sa20_sr_5, sa20_sr_6, sa20_sr_7, sa21_0, 
       sa21_1, sa21_2, sa21_3, sa21_4, sa21_5, sa21_6, sa21_7, sa21_sr_0, sa21_sr_1, 
       sa21_sr_2, sa21_sr_3, sa21_sr_4, sa21_sr_5, sa21_sr_6, sa21_sr_7, sa22_0, sa22_1, sa22_2, 
       sa22_3, sa22_4, sa22_5, sa22_6, sa22_7, sa22_sr_0, sa22_sr_1, sa22_sr_2, sa22_sr_3, 
       sa22_sr_4, sa22_sr_5, sa22_sr_6, sa22_sr_7, sa23_0, sa23_1, sa23_2, sa23_3, sa23_4, 
       sa23_5, sa23_6, sa23_7, sa23_sr_0, sa23_sr_1, sa23_sr_2, sa23_sr_3, sa23_sr_4, sa23_sr_5, 
       sa23_sr_6, sa23_sr_7, sa30_0, sa30_1, sa30_2, sa30_3, sa30_4, sa30_5, sa30_6, 
       sa30_7, sa30_sr_0, sa30_sr_1, sa30_sr_2, sa30_sr_3, sa30_sr_4, sa30_sr_5, sa30_sr_6, sa30_sr_7, 
       sa31_0, sa31_1, sa31_2, sa31_3, sa31_4, sa31_5, sa31_6, sa31_7, sa31_sr_0, 
       sa31_sr_1, sa31_sr_2, sa31_sr_3, sa31_sr_4, sa31_sr_5, sa31_sr_6, sa31_sr_7, sa32_0, sa32_1, 
       sa32_2, sa32_3, sa32_4, sa32_5, sa32_6, sa32_7, sa32_sr_0, sa32_sr_1, sa32_sr_2, 
       sa32_sr_3, sa32_sr_4, sa32_sr_5, sa32_sr_6, sa32_sr_7, sa33_0, sa33_1, sa33_2, sa33_3, 
       sa33_4, sa33_5, sa33_6, sa33_7, sa33_sr_0, sa33_sr_1, sa33_sr_2, sa33_sr_3, sa33_sr_4, 
       sa33_sr_5, sa33_sr_6, sa33_sr_7, u0_n268, u0_n270, u0_n272, u0_n274, u0_n49, u0_n53, 
       u0_n55, u0_n57, u0_n59, u0_n61, u0_n63, u0_subword_10, u0_subword_11, u0_subword_12, u0_subword_13, 
       u0_subword_14, u0_subword_15, u0_subword_16, u0_subword_17, u0_subword_18, u0_subword_19, u0_subword_20, u0_subword_21, u0_subword_22, 
       u0_subword_23, u0_subword_24, u0_subword_25, u0_subword_26, u0_subword_27, u0_subword_28, u0_subword_29, u0_subword_30, u0_subword_31, 
       u0_subword_6, u0_subword_8, u0_subword_9, w0_0, w0_1, w0_10, w0_11, w0_12, w0_13, 
       w0_15, w0_16, w0_18, w0_19, w0_2, w0_20, w0_25, w0_26, w0_27, 
       w0_28, w0_3, w0_30, w0_4, w0_5, w0_7, w0_8, w1_4, w1_7, 
       w2_0, w2_1, w2_10, w2_11, w2_13, w2_16, w2_18, w2_19, w2_2, 
       w2_20, w2_25, w2_26, w2_27, w2_28, w2_4, w2_7, w2_8, w2_9, 
       w3_0, w3_1, w3_10, w3_11, w3_12, w3_13, w3_15, w3_16, w3_17, 
       w3_18, w3_19, w3_2, w3_20, w3_21, w3_22, w3_23, w3_24, w3_25, 
       w3_26, w3_27, w3_28, w3_29, w3_3, w3_30, w3_31, w3_4, w3_5, 
       w3_6, w3_7, w3_8, w3_9 ;

  aes_aes_die_0 u0 ( clk, key, ld, rst, text_in, done, text_out, N100, N102, N105, N114, N116, N132, N133, N134, 
      N147, N148, N149, N150, N169, N227, N228, N229, N230, 
      N231, N233, N242, N244, N245, N246, N247, N258, N261, 
      N277, N278, N280, N35, N36, N37, N38, N40, N41, 
      N430, N434, N435, N436, N437, N438, N439, N440, N441, 
      N463, N52, N53, N54, N57, N66, N67, N68, N73, 
      N82, N83, N84, N85, N86, N87, N88, N89, N98, 
      N99, n1145, n1183, n1212, n1213, n1214, n1215, n1216, n1217, 
      n1219, n1220, n1221, n342, n348, n354, n362, n394, n396, 
      n414, n419, n433, n462, n469, n481, n482, n500, n506, 
      n515, n524, n534, n547, n562, n590, n636, n657, n665, 
      n786, n791, n817, n823, n830, n861, n870, n900, n905, 
      n911, n917, n923, n927, n937, n957, sa00_sr_0, sa00_sr_1, sa00_sr_2, 
      sa00_sr_3, sa00_sr_4, sa00_sr_5, sa00_sr_6, sa00_sr_7, sa01_sr_0, sa01_sr_1, sa01_sr_2, sa01_sr_3, 
      sa01_sr_4, sa01_sr_5, sa01_sr_6, sa01_sr_7, sa02_sr_0, sa02_sr_1, sa02_sr_2, sa02_sr_3, sa02_sr_4, 
      sa02_sr_5, sa02_sr_6, sa02_sr_7, sa03_sr_0, sa03_sr_1, sa03_sr_2, sa03_sr_3, sa03_sr_4, sa03_sr_5, 
      sa03_sr_6, sa03_sr_7, sa10_sr_0, sa10_sr_1, sa10_sr_2, sa10_sr_3, sa10_sr_4, sa10_sr_5, sa10_sr_6, 
      sa10_sr_7, sa11_sr_0, sa11_sr_1, sa11_sr_2, sa11_sr_3, sa11_sr_4, sa11_sr_5, sa11_sr_6, sa11_sr_7, 
      sa12_sr_0, sa12_sr_1, sa12_sr_2, sa12_sr_4, sa12_sr_5, sa12_sr_6, sa12_sr_7, sa20_sr_0, sa20_sr_1, 
      sa20_sr_2, sa20_sr_3, sa20_sr_4, sa20_sr_5, sa20_sr_6, sa20_sr_7, sa21_sr_0, sa21_sr_1, sa21_sr_2, 
      sa21_sr_3, sa21_sr_4, sa21_sr_5, sa21_sr_6, sa21_sr_7, sa22_sr_0, sa22_sr_1, sa22_sr_3, sa22_sr_4, 
      sa22_sr_5, sa22_sr_6, sa22_sr_7, sa23_sr_0, sa23_sr_1, sa23_sr_2, sa23_sr_3, sa23_sr_4, sa23_sr_5, 
      sa23_sr_6, sa23_sr_7, sa30_sr_0, sa30_sr_1, sa30_sr_2, sa30_sr_3, sa30_sr_4, sa30_sr_5, sa30_sr_6, 
      sa30_sr_7, sa31_sr_0, sa31_sr_1, sa31_sr_2, sa31_sr_3, sa31_sr_4, sa31_sr_5, sa31_sr_6, sa31_sr_7, 
      sa32_sr_0, sa32_sr_1, sa32_sr_2, sa32_sr_3, sa32_sr_4, sa32_sr_5, sa32_sr_6, sa32_sr_7, sa33_sr_0, 
      sa33_sr_1, sa33_sr_2, sa33_sr_3, sa33_sr_4, sa33_sr_5, sa33_sr_6, sa33_sr_7, u0_n49, u0_n53, 
      u0_n55, u0_n57, u0_n59, u0_n61, u0_n63, u0_subword_10, u0_subword_11, u0_subword_12, u0_subword_13, 
      u0_subword_14, u0_subword_15, u0_subword_16, u0_subword_17, u0_subword_18, u0_subword_19, u0_subword_20, u0_subword_21, u0_subword_22, 
      u0_subword_23, u0_subword_24, u0_subword_25, u0_subword_26, u0_subword_27, u0_subword_28, u0_subword_29, u0_subword_30, u0_subword_31, 
      u0_subword_6, u0_subword_8, u0_subword_9, n101, n103, n105, n1109, n1114, n115, 
      n117, n119, n121, n13, n143, n15, n195, n197, n199, 
      n201, n203, n207, n209, n21, n213, n215, n217, n219, 
      n225, n23, n231, n247, n249, n25, n253, n3, n31, 
      n33, n35, n37, n47, n49, n5, n51, n53, n55, 
      n57, n59, n61, n63, n65, n67, n69, n7, n73, 
      n79, n81, n85, n9, sa00_0, sa00_1, sa00_2, sa00_3, sa00_4, 
      sa00_5, sa00_6, sa00_7, sa01_0, sa01_1, sa01_2, sa01_3, sa01_4, sa01_5, 
      sa01_6, sa01_7, sa02_0, sa02_1, sa02_2, sa02_3, sa02_4, sa02_5, sa02_6, 
      sa02_7, sa03_0, sa03_1, sa03_2, sa03_3, sa03_4, sa03_5, sa03_6, sa03_7, 
      sa10_0, sa10_1, sa10_2, sa10_3, sa10_4, sa10_5, sa10_6, sa10_7, sa11_0, 
      sa11_1, sa11_2, sa11_3, sa11_4, sa11_5, sa11_6, sa11_7, sa12_0, sa12_1, 
      sa12_2, sa12_3, sa12_4, sa12_5, sa12_6, sa12_7, sa13_0, sa13_1, sa13_2, 
      sa13_3, sa13_4, sa13_5, sa13_6, sa13_7, sa20_0, sa20_1, sa20_2, sa20_3, 
      sa20_4, sa20_5, sa20_6, sa20_7, sa21_0, sa21_1, sa21_2, sa21_3, sa21_4, 
      sa21_5, sa21_6, sa21_7, sa22_0, sa22_1, sa22_2, sa22_3, sa22_4, sa22_5, 
      sa22_6, sa22_7, sa23_0, sa23_1, sa23_2, sa23_3, sa23_4, sa23_5, sa23_6, 
      sa23_7, sa30_0, sa30_1, sa30_2, sa30_3, sa30_4, sa30_5, sa30_6, sa30_7, 
      sa31_0, sa31_1, sa31_2, sa31_3, sa31_4, sa31_5, sa31_6, sa31_7, sa32_0, 
      sa32_1, sa32_2, sa32_3, sa32_4, sa32_5, sa32_6, sa32_7, sa33_0, sa33_1, 
      sa33_2, sa33_3, sa33_4, sa33_5, sa33_6, sa33_7, u0_n268, u0_n270, u0_n272, 
      u0_n274, w0_0, w0_1, w0_10, w0_11, w0_12, w0_13, w0_15, w0_16, 
      w0_18, w0_19, w0_2, w0_20, w0_25, w0_26, w0_27, w0_28, w0_3, 
      w0_30, w0_4, w0_5, w0_7, w0_8, w1_4, w1_7, w2_0, w2_1, 
      w2_10, w2_11, w2_13, w2_16, w2_18, w2_19, w2_2, w2_20, w2_25, 
      w2_26, w2_27, w2_28, w2_4, w2_7, w2_8, w2_9, w3_0, w3_1, 
      w3_10, w3_11, w3_12, w3_13, w3_15, w3_16, w3_17, w3_18, w3_19, 
      w3_2, w3_20, w3_21, w3_22, w3_23, w3_24, w3_25, w3_26, w3_27, 
      w3_28, w3_29, w3_3, w3_30, w3_31, w3_4, w3_5, w3_6, w3_7, 
      w3_8, w3_9 );
  aes_aes_die_1 u1 ( sa01_sr_3, sa01_sr_4, sa01_sr_7, sa03_0, sa03_1, sa03_2, sa03_3, sa03_4, sa03_5, 
      sa03_6, sa03_7, sa12_0, sa12_1, sa12_2, sa12_3, sa12_4, sa12_5, sa12_6, 
      sa12_7, sa21_0, sa21_1, sa21_2, sa21_3, sa21_4, sa21_5, sa21_6, sa21_7, 
      sa21_sr_4, sa31_sr_3, sa31_sr_7, w1_4, n657, n665, n786, n791, sa03_sr_0, 
      sa03_sr_1, sa03_sr_2, sa03_sr_3, sa03_sr_4, sa03_sr_5, sa03_sr_6, sa03_sr_7, sa11_sr_0, sa11_sr_1, 
      sa11_sr_2, sa11_sr_3, sa11_sr_4, sa11_sr_5, sa11_sr_6, sa11_sr_7, sa23_sr_0, sa23_sr_1, sa23_sr_2, 
      sa23_sr_3, sa23_sr_4, sa23_sr_5, sa23_sr_6, sa23_sr_7 );
  aes_aes_die_2 u2 ( sa02_0, sa02_1, sa02_2, sa02_3, sa02_4, sa02_5, sa02_6, sa02_7, sa30_0, 
      sa30_1, sa30_2, sa30_3, sa30_4, sa30_5, sa30_6, sa30_7, sa33_0, sa33_1, 
      sa33_2, sa33_3, sa33_4, sa33_5, sa33_6, sa33_7, sa02_sr_0, sa02_sr_1, sa02_sr_2, 
      sa02_sr_3, sa02_sr_4, sa02_sr_5, sa02_sr_6, sa02_sr_7, sa30_sr_0, sa30_sr_1, sa30_sr_2, sa30_sr_3, 
      sa30_sr_4, sa30_sr_5, sa30_sr_6, sa30_sr_7, sa31_sr_0, sa31_sr_1, sa31_sr_2, sa31_sr_3, sa31_sr_4, 
      sa31_sr_5, sa31_sr_6, sa31_sr_7 );
  aes_aes_die_3 u3 ( sa01_0, sa01_1, sa01_2, sa01_3, sa01_4, sa01_5, sa01_6, sa01_7, sa20_0, 
      sa20_1, sa20_2, sa20_3, sa20_4, sa20_5, sa20_6, sa20_7, sa32_0, sa32_1, 
      sa32_2, sa32_3, sa32_4, sa32_5, sa32_6, sa32_7, sa01_sr_0, sa01_sr_1, sa01_sr_2, 
      sa01_sr_3, sa01_sr_4, sa01_sr_5, sa01_sr_6, sa01_sr_7, sa22_sr_0, sa22_sr_1, sa22_sr_2, sa22_sr_3, 
      sa22_sr_4, sa22_sr_5, sa22_sr_6, sa22_sr_7, sa33_sr_0, sa33_sr_1, sa33_sr_2, sa33_sr_3, sa33_sr_4, 
      sa33_sr_5, sa33_sr_6, sa33_sr_7 );
  aes_aes_die_4 u4 ( sa00_0, sa00_1, sa00_2, sa00_3, sa00_4, sa00_5, sa00_6, sa00_7, sa23_0, 
      sa23_1, sa23_2, sa23_3, sa23_4, sa23_5, sa23_6, sa23_7, w3_0, w3_1, 
      w3_2, w3_3, w3_4, w3_5, w3_6, w3_7, sa00_sr_0, sa00_sr_1, sa00_sr_2, 
      sa00_sr_3, sa00_sr_4, sa00_sr_5, sa00_sr_6, sa00_sr_7, sa21_sr_0, sa21_sr_1, sa21_sr_2, sa21_sr_3, 
      sa21_sr_4, sa21_sr_5, sa21_sr_6, sa21_sr_7, u0_subword_10, u0_subword_11, u0_subword_12, u0_subword_13, u0_subword_14, 
      u0_subword_15, u0_subword_8, u0_subword_9 );
  aes_aes_die_5 u5 ( n101, n103, n105, n1109, n1114, n115, n117, n119, n121, 
      n13, n143, n15, n195, n197, n199, n201, n203, n207, 
      n209, n21, n213, n215, n217, n219, n225, n23, n231, 
      n247, n249, n25, n253, n3, n31, n33, n35, n37, 
      n47, n49, n5, n51, n53, n55, n57, n59, n61, 
      n63, n65, n665, n67, n69, n7, n73, n79, n81, 
      n85, n9, sa00_sr_0, sa00_sr_1, sa00_sr_2, sa00_sr_3, sa00_sr_4, sa00_sr_5, sa00_sr_6, 
      sa00_sr_7, sa01_sr_6, sa02_sr_0, sa02_sr_1, sa02_sr_2, sa02_sr_3, sa02_sr_4, sa02_sr_5, sa02_sr_6, 
      sa02_sr_7, sa03_sr_0, sa03_sr_1, sa03_sr_2, sa03_sr_3, sa03_sr_4, sa03_sr_5, sa03_sr_6, sa03_sr_7, 
      sa10_0, sa10_1, sa10_2, sa10_3, sa10_4, sa10_5, sa10_6, sa10_7, sa10_sr_0, 
      sa10_sr_1, sa10_sr_2, sa10_sr_3, sa10_sr_4, sa10_sr_5, sa10_sr_6, sa10_sr_7, sa12_sr_0, sa12_sr_1, 
      sa12_sr_2, sa12_sr_3, sa12_sr_4, sa12_sr_5, sa12_sr_7, sa20_sr_0, sa20_sr_1, sa20_sr_2, sa20_sr_3, 
      sa20_sr_4, sa20_sr_5, sa20_sr_6, sa20_sr_7, sa21_sr_7, sa22_sr_0, sa22_sr_1, sa22_sr_2, sa22_sr_3, 
      sa22_sr_4, sa22_sr_6, sa22_sr_7, sa23_sr_0, sa23_sr_1, sa23_sr_2, sa23_sr_3, sa23_sr_4, sa23_sr_5, 
      sa23_sr_6, sa23_sr_7, sa30_sr_0, sa30_sr_1, sa30_sr_2, sa30_sr_3, sa30_sr_4, sa30_sr_5, sa30_sr_6, 
      sa30_sr_7, sa31_sr_6, sa32_sr_0, sa32_sr_1, sa32_sr_2, sa32_sr_3, sa32_sr_4, sa32_sr_5, sa32_sr_6, 
      sa32_sr_7, sa33_sr_0, sa33_sr_1, sa33_sr_2, sa33_sr_3, sa33_sr_4, sa33_sr_5, sa33_sr_6, sa33_sr_7, 
      w0_0, w0_1, w0_10, w0_11, w0_12, w0_13, w0_15, w0_16, w0_18, 
      w0_19, w0_2, w0_20, w0_25, w0_26, w0_27, w0_28, w0_3, w0_30, 
      w0_4, w0_5, w0_7, w0_8, w1_7, w2_0, w2_1, w2_10, w2_11, 
      w2_13, w2_16, w2_18, w2_19, w2_2, w2_20, w2_25, w2_26, w2_27, 
      w2_28, w2_4, w2_7, w2_8, w2_9, w3_0, w3_1, w3_10, w3_11, 
      w3_12, w3_13, w3_15, w3_16, w3_17, w3_18, w3_19, w3_2, w3_20, 
      w3_21, w3_22, w3_23, w3_24, w3_25, w3_26, w3_27, w3_28, w3_29, 
      w3_3, w3_30, w3_31, w3_4, w3_5, w3_6, w3_7, w3_8, w3_9, 
      N100, N102, N105, N114, N116, N132, N133, N134, N147, 
      N148, N149, N150, N169, N227, N228, N229, N230, N231, 
      N233, N242, N244, N245, N246, N247, N258, N261, N277, 
      N278, N280, N35, N36, N37, N38, N40, N41, N430, 
      N434, N435, N436, N437, N438, N439, N440, N441, N463, 
      N52, N53, N54, N57, N66, N67, N68, N73, N82, 
      N83, N84, N85, N86, N87, N88, N89, N98, N99, 
      n1145, n1183, n1212, n1213, n1214, n1215, n1216, n1217, n1219, 
      n1220, n1221, n342, n348, n354, n362, n394, n396, n414, 
      n419, n433, n462, n469, n481, n482, n500, n506, n515, 
      n524, n534, n547, n562, n590, n636, n817, n823, n830, 
      n861, n870, n900, n905, n911, n917, n923, n927, n937, 
      n957, u0_n49, u0_n53, u0_n55, u0_n57, u0_n59, u0_n61, u0_n63, u0_subword_6 );
  aes_aes_die_6 u6 ( sa11_0, sa11_1, sa11_2, sa11_3, sa11_4, sa11_5, sa11_6, sa11_7, sa22_0, 
      sa22_1, sa22_2, sa22_3, sa22_4, sa22_5, sa22_6, sa22_7, u0_n268, u0_n270, 
      u0_n272, u0_n274, w3_10, w3_11, w3_8, w3_9, sa10_sr_0, sa10_sr_1, sa10_sr_2, 
      sa10_sr_3, sa10_sr_4, sa10_sr_5, sa10_sr_6, sa10_sr_7, sa20_sr_0, sa20_sr_1, sa20_sr_2, sa20_sr_3, 
      sa20_sr_4, sa20_sr_5, sa20_sr_6, sa20_sr_7, u0_subword_16, u0_subword_17, u0_subword_18, u0_subword_19, u0_subword_20, 
      u0_subword_21, u0_subword_22, u0_subword_23 );
  aes_aes_die_7 u7 ( sa13_0, sa13_1, sa13_2, sa13_3, sa13_4, sa13_5, sa13_6, sa13_7, sa31_0, 
      sa31_1, sa31_2, sa31_3, sa31_4, sa31_5, sa31_6, sa31_7, w3_16, w3_17, 
      w3_18, w3_19, w3_20, w3_21, w3_22, w3_23, sa12_sr_0, sa12_sr_1, sa12_sr_2, 
      sa12_sr_3, sa12_sr_4, sa12_sr_5, sa12_sr_6, sa12_sr_7, sa32_sr_0, sa32_sr_1, sa32_sr_2, sa32_sr_3, 
      sa32_sr_4, sa32_sr_5, sa32_sr_6, sa32_sr_7, u0_subword_24, u0_subword_25, u0_subword_26, u0_subword_27, u0_subword_28, 
      u0_subword_29, u0_subword_30, u0_subword_31 );
endmodule
