module aes_aes_die_5 ( n101, n103, n105, n107, n1109, n111, n1114, n113, n115, 
       n117, n119, n121, n1212, n1213, n1214, n1215, n1216, n1217, 
       n1218, n1219, n1220, n1221, n123, n125, n127, n193, n197, 
       n199, n201, n203, n207, n209, n211, n213, n215, n217, 
       n219, n223, n227, n229, n231, n233, n235, n237, n245, 
       n247, n251, n253, n482, n488, n65, n69, n71, n73, 
       n77, n79, n81, n83, n85, n87, n89, n91, n93, 
       n95, n97, n99, sa00_sr_0, sa00_sr_1, sa00_sr_2, sa00_sr_3, sa00_sr_4, sa00_sr_5, 
       sa00_sr_6, sa00_sr_7, sa02_sr_0, sa02_sr_1, sa02_sr_2, sa02_sr_3, sa02_sr_4, sa02_sr_5, sa02_sr_6, 
       sa02_sr_7, sa10_sr_0, sa10_sr_1, sa10_sr_2, sa10_sr_3, sa10_sr_4, sa10_sr_5, sa10_sr_6, sa10_sr_7, 
       sa12_sr_0, sa12_sr_1, sa12_sr_2, sa12_sr_3, sa12_sr_4, sa12_sr_5, sa12_sr_6, sa12_sr_7, sa20_sr_0, 
       sa20_sr_1, sa20_sr_2, sa20_sr_3, sa20_sr_4, sa20_sr_5, sa20_sr_6, sa20_sr_7, sa22_sr_0, sa22_sr_1, 
       sa22_sr_2, sa22_sr_3, sa22_sr_4, sa22_sr_5, sa22_sr_6, sa22_sr_7, sa30_sr_0, sa30_sr_1, sa30_sr_2, 
       sa30_sr_3, sa30_sr_4, sa30_sr_5, sa30_sr_6, sa30_sr_7, sa32_sr_0, sa32_sr_1, sa32_sr_2, sa32_sr_3, 
       sa32_sr_4, sa32_sr_5, sa32_sr_6, sa32_sr_7, u0_n162, u0_n164, u0_n166, u0_n168, u0_n170, 
       u0_n174, w0_0, w0_1, w0_10, w0_11, w0_12, w0_13, w0_15, w0_17, 
       w0_18, w0_19, w0_2, w0_20, w0_21, w0_22, w0_26, w0_27, w0_28, 
       w0_29, w0_3, w0_30, w0_4, w0_5, w0_6, w0_7, w0_8, w0_9, 
       w1_3, w1_6, w1_7, w2_0, w2_10, w2_11, w2_12, w2_13, w2_14, 
       w2_15, w2_16, w2_17, w2_18, w2_19, w2_2, w2_20, w2_21, w2_23, 
       w2_24, w2_25, w2_26, w2_27, w2_28, w2_29, w2_3, w2_30, w2_31, 
       w2_4, w2_5, w2_6, w2_7, w2_8, w2_9, w3_24, w3_25, w3_26, 
       w3_27, w3_28, w3_29, w3_30, w3_31, N100, N101, N102, N104, N105, N114, N115, N116, N117, 
        N118, N119, N120, N121, N130, N131, N132, N133, N134, 
        N135, N137, N146, N147, N148, N149, N150, N151, N152, 
        N153, N226, N228, N229, N230, N231, N233, N242, N243, 
        N244, N245, N246, N247, N249, N259, N260, N261, N262, 
        N263, N264, N276, N277, N279, N280, N379, N380, N381, 
        N382, N383, N394, N395, N396, N397, N398, N399, N400, 
        N401, N411, N412, N413, N414, N415, N416, N426, N429, 
        N430, N431, N432, N433, N442, N444, N445, N446, N447, 
        N448, N449, N458, N459, N461, N462, N463, N464, N465, 
        N474, N477, N478, N479, N480, N481, N490, N491, N492, 
        N493, N494, N495, N98, n1133, n469, n485, n508, n515, 
        n560, n630, n870, n956, u0_n139, u0_n142, u0_n151, u0_n210, u0_n212, 
        u0_n218, u0_n49, u0_n51, u0_n53, u0_n55, u0_n57, u0_n59, u0_n61, u0_n63, 
        u0_n65, u0_n67, u0_n68, u0_n70, u0_n71, u0_n73, u0_n74, u0_n76, u0_n77, 
        u0_n79, u0_n83, u0_n85 );
  input n101, n103, n105, n107, n1109, n111, n1114, n113, n115, 
        n117, n119, n121, n1212, n1213, n1214, n1215, n1216, n1217, 
        n1218, n1219, n1220, n1221, n123, n125, n127, n193, n197, 
        n199, n201, n203, n207, n209, n211, n213, n215, n217, 
        n219, n223, n227, n229, n231, n233, n235, n237, n245, 
        n247, n251, n253, n482, n488, n65, n69, n71, n73, 
        n77, n79, n81, n83, n85, n87, n89, n91, n93, 
        n95, n97, n99, sa00_sr_0, sa00_sr_1, sa00_sr_2, sa00_sr_3, sa00_sr_4, sa00_sr_5, 
        sa00_sr_6, sa00_sr_7, sa02_sr_0, sa02_sr_1, sa02_sr_2, sa02_sr_3, sa02_sr_4, sa02_sr_5, sa02_sr_6, 
        sa02_sr_7, sa10_sr_0, sa10_sr_1, sa10_sr_2, sa10_sr_3, sa10_sr_4, sa10_sr_5, sa10_sr_6, sa10_sr_7, 
        sa12_sr_0, sa12_sr_1, sa12_sr_2, sa12_sr_3, sa12_sr_4, sa12_sr_5, sa12_sr_6, sa12_sr_7, sa20_sr_0, 
        sa20_sr_1, sa20_sr_2, sa20_sr_3, sa20_sr_4, sa20_sr_5, sa20_sr_6, sa20_sr_7, sa22_sr_0, sa22_sr_1, 
        sa22_sr_2, sa22_sr_3, sa22_sr_4, sa22_sr_5, sa22_sr_6, sa22_sr_7, sa30_sr_0, sa30_sr_1, sa30_sr_2, 
        sa30_sr_3, sa30_sr_4, sa30_sr_5, sa30_sr_6, sa30_sr_7, sa32_sr_0, sa32_sr_1, sa32_sr_2, sa32_sr_3, 
        sa32_sr_4, sa32_sr_5, sa32_sr_6, sa32_sr_7, u0_n162, u0_n164, u0_n166, u0_n168, u0_n170, 
        u0_n174, w0_0, w0_1, w0_10, w0_11, w0_12, w0_13, w0_15, w0_17, 
        w0_18, w0_19, w0_2, w0_20, w0_21, w0_22, w0_26, w0_27, w0_28, 
        w0_29, w0_3, w0_30, w0_4, w0_5, w0_6, w0_7, w0_8, w0_9, 
        w1_3, w1_6, w1_7, w2_0, w2_10, w2_11, w2_12, w2_13, w2_14, 
        w2_15, w2_16, w2_17, w2_18, w2_19, w2_2, w2_20, w2_21, w2_23, 
        w2_24, w2_25, w2_26, w2_27, w2_28, w2_29, w2_3, w2_30, w2_31, 
        w2_4, w2_5, w2_6, w2_7, w2_8, w2_9, w3_24, w3_25, w3_26, 
        w3_27, w3_28, w3_29, w3_30, w3_31;
  output N100, N101, N102, N104, N105, N114, N115, N116, N117, 
        N118, N119, N120, N121, N130, N131, N132, N133, N134, 
        N135, N137, N146, N147, N148, N149, N150, N151, N152, 
        N153, N226, N228, N229, N230, N231, N233, N242, N243, 
        N244, N245, N246, N247, N249, N259, N260, N261, N262, 
        N263, N264, N276, N277, N279, N280, N379, N380, N381, 
        N382, N383, N394, N395, N396, N397, N398, N399, N400, 
        N401, N411, N412, N413, N414, N415, N416, N426, N429, 
        N430, N431, N432, N433, N442, N444, N445, N446, N447, 
        N448, N449, N458, N459, N461, N462, N463, N464, N465, 
        N474, N477, N478, N479, N480, N481, N490, N491, N492, 
        N493, N494, N495, N98, n1133, n469, n485, n508, n515, 
        n560, n630, n870, n956, u0_n139, u0_n142, u0_n151, u0_n210, u0_n212, 
        u0_n218, u0_n49, u0_n51, u0_n53, u0_n55, u0_n57, u0_n59, u0_n61, u0_n63, 
        u0_n65, u0_n67, u0_n68, u0_n70, u0_n71, u0_n73, u0_n74, u0_n76, u0_n77, 
        u0_n79, u0_n83, u0_n85;
  wire n1117, n1118, n1126, n1127, n1128, n1130, n1132, n1135, n1136, 
       n1138, n1139, n1144, n1145, n1148, n1149, n1150, n1151, n1153, 
       n1154, n1155, n1156, n1158, n1160, n1164, n1168, n1172, n1173, 
       n1178, n1179, n1181, n1183, n1186, n1188, n1194, n1196, n1204, 
       n1206, n1208, n1209, n1210, n1211, n277, n278, n279, n280, 
       n281, n283, n284, n472, n473, n475, n476, n477, n478, 
       n479, n481, n483, n486, n487, n489, n490, n491, n492, 
       n493, n495, n496, n497, n498, n499, n500, n502, n503, 
       n504, n509, n510, n516, n522, n523, n524, n526, n528, 
       n529, n530, n531, n532, n533, n534, n535, n536, n537, 
       n538, n539, n540, n541, n542, n543, n544, n546, n547, 
       n548, n550, n551, n552, n554, n555, n556, n561, n562, 
       n564, n569, n570, n571, n572, n573, n574, n575, n576, 
       n577, n578, n579, n581, n582, n583, n584, n586, n587, 
       n588, n590, n591, n592, n593, n595, n596, n597, n598, 
       n599, n600, n606, n607, n608, n609, n610, n611, n612, 
       n613, n614, n615, n616, n617, n618, n619, n620, n622, 
       n623, n624, n625, n626, n628, n632, n633, n634, n635, 
       n636, n638, n813, n814, n816, n817, n818, n819, n820, 
       n821, n823, n824, n825, n826, n827, n828, n829, n830, 
       n831, n832, n833, n834, n835, n836, n837, n838, n839, 
       n840, n841, n843, n844, n845, n846, n847, n848, n850, 
       n851, n852, n853, n854, n856, n857, n858, n859, n861, 
       n862, n863, n864, n865, n866, n867, n874, n875, n876, 
       n877, n878, n879, n880, n881, n882, n883, n884, n885, 
       n886, n887, n888, n889, n890, n892, n893, n894, n896, 
       n898, n899, n900, n901, n902, n903, n904, n905, n907, 
       n908, n909, n911, n912, n913, n915, n916, n917, n918, 
       n919, n920, n921, n922, n923, n924, n925, n926, n927, 
       n929, n930, n931, n932, n933, n935, n936, n937, n939, 
       n940, n941, n942, n944, n945, n946, n947, n948, n949, 
       n950, n951, n952, n954, n957, n958, n959, n960, n961, 
       n962, n964, n965, n966, n967, n969, n970, n971, n972, 
       n973, n974, n975, n976, u0_subword_0, u0_subword_1, u0_subword_2, u0_subword_3, u0_subword_4, 
       u0_subword_5, u0_subword_6, u0_subword_7, u0_u3_n41, u0_u3_n438, u0_u3_n439, u0_u3_n440, u0_u3_n441, u0_u3_n442, 
       u0_u3_n443, u0_u3_n444, u0_u3_n445, u0_u3_n446, u0_u3_n447, u0_u3_n448, u0_u3_n449, u0_u3_n450, u0_u3_n451, 
       u0_u3_n452, u0_u3_n453, u0_u3_n454, u0_u3_n455, u0_u3_n456, u0_u3_n457, u0_u3_n458, u0_u3_n459, u0_u3_n460, 
       u0_u3_n461, u0_u3_n462, u0_u3_n463, u0_u3_n464, u0_u3_n465, u0_u3_n466, u0_u3_n467, u0_u3_n468, u0_u3_n469, 
       u0_u3_n470, u0_u3_n471, u0_u3_n472, u0_u3_n473, u0_u3_n474, u0_u3_n475, u0_u3_n476, u0_u3_n477, u0_u3_n478, 
       u0_u3_n479, u0_u3_n480, u0_u3_n481, u0_u3_n482, u0_u3_n483, u0_u3_n484, u0_u3_n485, u0_u3_n486, u0_u3_n487, 
       u0_u3_n488, u0_u3_n489, u0_u3_n490, u0_u3_n491, u0_u3_n492, u0_u3_n493, u0_u3_n494, u0_u3_n495, u0_u3_n496, 
       u0_u3_n497, u0_u3_n498, u0_u3_n499, u0_u3_n500, u0_u3_n501, u0_u3_n502, u0_u3_n503, u0_u3_n504, u0_u3_n505, 
       u0_u3_n506, u0_u3_n507, u0_u3_n508, u0_u3_n509, u0_u3_n510, u0_u3_n511, u0_u3_n512, u0_u3_n513, u0_u3_n514, 
       u0_u3_n515, u0_u3_n516, u0_u3_n517, u0_u3_n518, u0_u3_n519, u0_u3_n520, u0_u3_n521, u0_u3_n522, u0_u3_n523, 
       u0_u3_n524, u0_u3_n525, u0_u3_n526, u0_u3_n527, u0_u3_n528, u0_u3_n529, u0_u3_n530, u0_u3_n531, u0_u3_n532, 
       u0_u3_n533, u0_u3_n534, u0_u3_n535, u0_u3_n536, u0_u3_n537, u0_u3_n538, u0_u3_n539, u0_u3_n540, u0_u3_n541, 
       u0_u3_n542, u0_u3_n543, u0_u3_n544, u0_u3_n545, u0_u3_n546, u0_u3_n547, u0_u3_n548, u0_u3_n549, u0_u3_n550, 
       u0_u3_n551, u0_u3_n552, u0_u3_n553, u0_u3_n554, u0_u3_n555, u0_u3_n556, u0_u3_n557, u0_u3_n558, u0_u3_n559, 
       u0_u3_n560, u0_u3_n561, u0_u3_n562, u0_u3_n563, u0_u3_n564, u0_u3_n565, u0_u3_n566, u0_u3_n567, u0_u3_n568, 
       u0_u3_n569, u0_u3_n570, u0_u3_n571, u0_u3_n572, u0_u3_n573, u0_u3_n574, u0_u3_n575, u0_u3_n576, u0_u3_n577, 
       u0_u3_n578, u0_u3_n579, u0_u3_n580, u0_u3_n581, u0_u3_n582, u0_u3_n583, u0_u3_n584, u0_u3_n585, u0_u3_n586, 
       u0_u3_n587, u0_u3_n588, u0_u3_n589, u0_u3_n590, u0_u3_n591, u0_u3_n592, u0_u3_n593, u0_u3_n594, u0_u3_n595, 
       u0_u3_n596, u0_u3_n597, u0_u3_n598, u0_u3_n599, u0_u3_n600, u0_u3_n601, u0_u3_n602, u0_u3_n603, u0_u3_n604, 
       u0_u3_n605, u0_u3_n606, u0_u3_n607, u0_u3_n608, u0_u3_n609, u0_u3_n610, u0_u3_n611, u0_u3_n612, u0_u3_n613, 
       u0_u3_n614, u0_u3_n615, u0_u3_n616, u0_u3_n617, u0_u3_n618, u0_u3_n619, u0_u3_n620, u0_u3_n621, u0_u3_n622, 
       u0_u3_n623, u0_u3_n624, u0_u3_n625, u0_u3_n626, u0_u3_n627, u0_u3_n628, u0_u3_n629, u0_u3_n630, u0_u3_n631, 
       u0_u3_n632, u0_u3_n633, u0_u3_n634, u0_u3_n635, u0_u3_n636, u0_u3_n637, u0_u3_n638, u0_u3_n639, u0_u3_n640, 
       u0_u3_n641, u0_u3_n642, u0_u3_n643, u0_u3_n644, u0_u3_n645, u0_u3_n646, u0_u3_n647, u0_u3_n648, u0_u3_n649, 
       u0_u3_n650, u0_u3_n651, u0_u3_n652, u0_u3_n653, u0_u3_n654, u0_u3_n655, u0_u3_n656, u0_u3_n657, u0_u3_n658, 
       u0_u3_n659, u0_u3_n660, u0_u3_n661, u0_u3_n662, u0_u3_n663, u0_u3_n664, u0_u3_n665, u0_u3_n666, u0_u3_n667, 
       u0_u3_n668, u0_u3_n669, u0_u3_n670, u0_u3_n671, u0_u3_n672, u0_u3_n673, u0_u3_n674, u0_u3_n675, u0_u3_n676, 
       u0_u3_n677, u0_u3_n678, u0_u3_n679, u0_u3_n680, u0_u3_n681, u0_u3_n682, u0_u3_n683, u0_u3_n684, u0_u3_n685, 
       u0_u3_n686, u0_u3_n687, u0_u3_n688, u0_u3_n689, u0_u3_n690, u0_u3_n691, u0_u3_n692, u0_u3_n693, u0_u3_n694, 
       u0_u3_n695, u0_u3_n696, u0_u3_n697, u0_u3_n698, u0_u3_n699, u0_u3_n700, u0_u3_n701, u0_u3_n702, u0_u3_n703, 
       u0_u3_n704, u0_u3_n705, u0_u3_n706, u0_u3_n707, u0_u3_n708, u0_u3_n709, u0_u3_n710, u0_u3_n711, u0_u3_n712, 
       u0_u3_n713, u0_u3_n714, u0_u3_n715, u0_u3_n716, u0_u3_n717, u0_u3_n718, u0_u3_n719, u0_u3_n720, u0_u3_n721, 
       u0_u3_n722, u0_u3_n723, u0_u3_n724, u0_u3_n725, u0_u3_n726, u0_u3_n727, u0_u3_n728, u0_u3_n729, u0_u3_n730, 
       u0_u3_n731, u0_u3_n732, u0_u3_n733, u0_u3_n734, u0_u3_n735, u0_u3_n736, u0_u3_n737, u0_u3_n738, u0_u3_n739, 
       u0_u3_n740, u0_u3_n741, u0_u3_n742, u0_u3_n743, u0_u3_n744, u0_u3_n745, u0_u3_n746, u0_u3_n747, u0_u3_n748, 
       u0_u3_n749, u0_u3_n750, u0_u3_n751, u0_u3_n752, u0_u3_n753, u0_u3_n754, u0_u3_n755, u0_u3_n756, u0_u3_n757, 
       u0_u3_n758, u0_u3_n759, u0_u3_n760, u0_u3_n761, u0_u3_n762, u0_u3_n763, u0_u3_n764, u0_u3_n765, u0_u3_n766, 
       u0_u3_n767, u0_u3_n768, u0_u3_n769, u0_u3_n770, u0_u3_n771, u0_u3_n772, u0_u3_n773, u0_u3_n774, u0_u3_n775, 
       u0_u3_n776, u0_u3_n777, u0_u3_n778, u0_u3_n779, u0_u3_n780, u0_u3_n781, u0_u3_n782, u0_u3_n783, u0_u3_n784, 
       u0_u3_n785, u0_u3_n786, u0_u3_n787, u0_u3_n788, u0_u3_n789, u0_u3_n790, u0_u3_n791, u0_u3_n792, u0_u3_n793, 
       u0_u3_n794, u0_u3_n795, u0_u3_n796, u0_u3_n797, u0_u3_n798, u0_u3_n799, u0_u3_n800, u0_u3_n801, u0_u3_n802, 
       u0_u3_n803, u0_u3_n804, u0_u3_n805, u0_u3_n806, u0_u3_n807, u0_u3_n808, u0_u3_n809, u0_u3_n810, u0_u3_n811, 
       u0_u3_n812, u0_u3_n813, u0_u3_n814, u0_u3_n815, u0_u3_n816, u0_u3_n817, u0_u3_n818, u0_u3_n819, u0_u3_n820, 
       u0_u3_n821, u0_u3_n822, u0_u3_n823, u0_u3_n824, u0_u3_n825, u0_u3_n826, u0_u3_n827, u0_u3_n828, u0_u3_n829, 
       u0_u3_n830, u0_u3_n831, u0_u3_n832, u0_u3_n833, u0_u3_n834, u0_u3_n835, u0_u3_n836, u0_u3_n837, u0_u3_n838, 
       u0_u3_n839, u0_u3_n840, u0_u3_n841, u0_u3_n842, u0_u3_n843, u0_u3_n844, u0_u3_n845, u0_u3_n846, u0_u3_n847, 
       u0_u3_n848, u0_u3_n849, u0_u3_n850, u0_u3_n851, u0_u3_n852, u0_u3_n853, u0_u3_n854, u0_u3_n855, u0_u3_n856, 
       u0_u3_n857, u0_u3_n858, u0_u3_n859, u0_u3_n860, u0_u3_n861, u0_u3_n862, u0_u3_n863, u0_u3_n864, u0_u3_n865, 
       u0_u3_n866, u0_u3_n867, u0_u3_n868, u0_u3_n869, u0_u3_n870, u0_u3_n871, u0_u3_n872, u0_u3_n873, u0_u3_n874, 
       u0_u3_n875, u0_u3_n876, u0_u3_n877,  u0_u3_n878;
  OAI22_X1 U1140 (.ZN( N153 ) , .A1( n1215 ) , .B2( n1218 ) , .A2( n813 ) , .B1( n814 ) );
  XOR2_X1 U1142 (.Z( n816 ) , .A( n817 ) , .B( n818 ) );
  INV_X1 U1144 (.ZN( n819 ) , .A( sa12_sr_7 ) );
  XOR2_X1 U1145 (.A( n127 ) , .Z( n813 ) , .B( w2_31 ) );
  OAI22_X1 U1147 (.ZN( N152 ) , .A1( n1215 ) , .B2( n1217 ) , .A2( n820 ) , .B1( n821 ) );
  XOR2_X1 U1149 (.Z( n823 ) , .A( n824 ) , .B( n825 ) );
  XOR2_X1 U1151 (.A( n125 ) , .Z( n820 ) , .B( w2_30 ) );
  OAI22_X1 U1153 (.ZN( N151 ) , .A1( n1215 ) , .B2( n1218 ) , .A2( n826 ) , .B1( n827 ) );
  XOR2_X1 U1154 (.Z( n827 ) , .A( n828 ) , .B( n829 ) );
  XOR2_X1 U1155 (.Z( n829 ) , .A( n830 ) , .B( n831 ) );
  XNOR2_X1 U1156 (.ZN( n828 ) , .B( sa12_sr_5 ) , .A( w2_29 ) );
  XOR2_X1 U1157 (.A( n123 ) , .Z( n826 ) , .B( w2_29 ) );
  OAI22_X1 U1159 (.ZN( N150 ) , .A1( n1215 ) , .B2( n1221 ) , .A2( n832 ) , .B1( n833 ) );
  XOR2_X1 U1160 (.Z( n833 ) , .A( n834 ) , .B( n835 ) );
  XOR2_X1 U1161 (.Z( n835 ) , .A( n836 ) , .B( n837 ) );
  XOR2_X1 U1162 (.Z( n834 ) , .A( n838 ) , .B( n839 ) );
  XNOR2_X1 U1163 (.ZN( n838 ) , .B( sa12_sr_4 ) , .A( w2_28 ) );
  XOR2_X1 U1164 (.A( n121 ) , .Z( n832 ) , .B( w2_28 ) );
  OAI22_X1 U1166 (.ZN( N149 ) , .A1( n1215 ) , .B2( n1221 ) , .A2( n840 ) , .B1( n841 ) );
  XOR2_X1 U1168 (.Z( n843 ) , .B( n844 ) , .A( n845 ) );
  XNOR2_X1 U1170 (.ZN( n846 ) , .B( sa12_sr_3 ) , .A( w2_27 ) );
  XOR2_X1 U1171 (.A( n119 ) , .Z( n840 ) , .B( w2_27 ) );
  OAI22_X1 U1173 (.ZN( N148 ) , .A1( n1215 ) , .B2( n1219 ) , .A2( n847 ) , .B1( n848 ) );
  XOR2_X1 U1175 (.A( n277 ) , .Z( n850 ) , .B( n851 ) );
  XOR2_X1 U1177 (.A( n117 ) , .Z( n847 ) , .B( w2_26 ) );
  OAI22_X1 U1179 (.ZN( N147 ) , .A1( n1215 ) , .B2( n1221 ) , .A2( n852 ) , .B1( n853 ) );
  XOR2_X1 U1182 (.B( n284 ) , .Z( n854 ) , .A( n857 ) );
  XNOR2_X1 U1183 (.ZN( n857 ) , .B( sa12_sr_1 ) , .A( w2_25 ) );
  XOR2_X1 U1184 (.A( n115 ) , .Z( n852 ) , .B( w2_25 ) );
  OAI22_X1 U1186 (.ZN( N146 ) , .A1( n1215 ) , .B2( n1217 ) , .A2( n858 ) , .B1( n859 ) );
  XOR2_X1 U1188 (.A( n836 ) , .Z( n861 ) , .B( n862 ) );
  XOR2_X1 U1190 (.A( n113 ) , .Z( n858 ) , .B( w2_24 ) );
  OAI22_X1 U1192 (.ZN( N137 ) , .A1( n1215 ) , .B2( n1218 ) , .A2( n863 ) , .B1( n864 ) );
  XOR2_X1 U1193 (.Z( n864 ) , .A( n865 ) , .B( n866 ) );
  XOR2_X1 U1194 (.B( n817 ) , .Z( n866 ) , .A( sa02_sr_7 ) );
  XNOR2_X1 U1195 (.ZN( n865 ) , .B( n867 ) , .A( sa12_sr_6 ) );
  XOR2_X1 U1196 (.Z( n867 ) , .B( sa22_sr_6 ) , .A( w2_23 ) );
  XOR2_X1 U1197 (.A( n111 ) , .Z( n863 ) , .B( w2_23 ) );
  OAI22_X1 U1207 (.ZN( N135 ) , .A1( n1213 ) , .B2( n1219 ) , .A2( n874 ) , .B1( n875 ) );
  XOR2_X1 U1208 (.Z( n875 ) , .A( n876 ) , .B( n877 ) );
  XOR2_X1 U1209 (.Z( n877 ) , .B( n878 ) , .A( sa12_sr_4 ) );
  XOR2_X1 U1210 (.Z( n878 ) , .B( sa22_sr_4 ) , .A( w2_21 ) );
  XNOR2_X1 U1211 (.B( n831 ) , .ZN( n876 ) , .A( sa02_sr_5 ) );
  XOR2_X1 U1212 (.A( n107 ) , .Z( n874 ) , .B( w2_21 ) );
  OAI22_X1 U1214 (.ZN( N134 ) , .A1( n1212 ) , .B2( n1219 ) , .A2( n879 ) , .B1( n880 ) );
  XOR2_X1 U1215 (.Z( n880 ) , .A( n881 ) , .B( n882 ) );
  XOR2_X1 U1216 (.Z( n882 ) , .B( n883 ) , .A( sa12_sr_3 ) );
  XOR2_X1 U1217 (.Z( n883 ) , .B( sa22_sr_3 ) , .A( w2_20 ) );
  XOR2_X1 U1218 (.Z( n881 ) , .A( n884 ) , .B( n885 ) );
  XNOR2_X1 U1219 (.B( n839 ) , .ZN( n884 ) , .A( sa02_sr_4 ) );
  XOR2_X1 U1220 (.A( n105 ) , .Z( n879 ) , .B( w2_20 ) );
  OAI22_X1 U1222 (.ZN( N133 ) , .A1( n1213 ) , .B2( n1219 ) , .A2( n886 ) , .B1( n887 ) );
  XOR2_X1 U1223 (.Z( n887 ) , .A( n888 ) , .B( n889 ) );
  XOR2_X1 U1224 (.Z( n889 ) , .B( n890 ) , .A( sa12_sr_2 ) );
  XOR2_X1 U1225 (.Z( n890 ) , .B( sa22_sr_2 ) , .A( w2_19 ) );
  XOR2_X1 U1228 (.A( n103 ) , .Z( n886 ) , .B( w2_19 ) );
  OAI22_X1 U1230 (.ZN( N132 ) , .A1( n1212 ) , .B2( n1219 ) , .A2( n892 ) , .B1( n893 ) );
  XOR2_X1 U1233 (.Z( n896 ) , .B( sa22_sr_1 ) , .A( w2_18 ) );
  XOR2_X1 U1236 (.A( n101 ) , .Z( n892 ) , .B( w2_18 ) );
  OAI22_X1 U1238 (.ZN( N131 ) , .A1( n1212 ) , .B2( n1219 ) , .A2( n898 ) , .B1( n899 ) );
  XOR2_X1 U1239 (.Z( n899 ) , .A( n900 ) , .B( n901 ) );
  XOR2_X1 U1240 (.Z( n901 ) , .B( n902 ) , .A( sa12_sr_0 ) );
  XOR2_X1 U1241 (.Z( n902 ) , .B( sa22_sr_0 ) , .A( w2_17 ) );
  XOR2_X1 U1242 (.B( n885 ) , .Z( n900 ) , .A( n903 ) );
  XNOR2_X1 U1243 (.B( n856 ) , .ZN( n903 ) , .A( sa02_sr_1 ) );
  XOR2_X1 U1244 (.Z( n898 ) , .A( n99 ) , .B( w2_17 ) );
  OAI22_X1 U1246 (.ZN( N130 ) , .A1( n1213 ) , .B2( n1219 ) , .A2( n904 ) , .B1( n905 ) );
  XOR2_X1 U1248 (.A( n862 ) , .B( n885 ) , .Z( n907 ) );
  XOR2_X1 U1249 (.Z( n885 ) , .A( sa12_sr_7 ) , .B( sa22_sr_7 ) );
  XOR2_X1 U1251 (.Z( n904 ) , .A( n97 ) , .B( w2_16 ) );
  OAI22_X1 U1253 (.ZN( N121 ) , .A1( n1109 ) , .B2( n1219 ) , .A2( n908 ) , .B1( n909 ) );
  XOR2_X1 U1255 (.A( n824 ) , .B( n836 ) , .Z( n911 ) );
  XOR2_X1 U1256 (.Z( n824 ) , .A( sa22_sr_6 ) , .B( sa32_sr_6 ) );
  XOR2_X1 U1258 (.Z( n908 ) , .A( n95 ) , .B( w2_15 ) );
  OAI22_X1 U1260 (.ZN( N120 ) , .A1( n1109 ) , .B2( n1220 ) , .A2( n912 ) , .B1( n913 ) );
  XOR2_X1 U1262 (.A( n818 ) , .B( n831 ) , .Z( n915 ) );
  XOR2_X1 U1263 (.Z( n831 ) , .A( sa22_sr_5 ) , .B( sa32_sr_5 ) );
  XOR2_X1 U1265 (.Z( n912 ) , .A( n93 ) , .B( w2_14 ) );
  OAI22_X1 U1267 (.ZN( N119 ) , .A1( n1109 ) , .B2( n1218 ) , .A2( n916 ) , .B1( n917 ) );
  XOR2_X1 U1268 (.Z( n917 ) , .A( n918 ) , .B( n919 ) );
  XOR2_X1 U1269 (.A( n825 ) , .B( n839 ) , .Z( n919 ) );
  XOR2_X1 U1270 (.Z( n839 ) , .A( sa22_sr_4 ) , .B( sa32_sr_4 ) );
  XNOR2_X1 U1271 (.ZN( n918 ) , .B( sa32_sr_5 ) , .A( w2_13 ) );
  XOR2_X1 U1272 (.A( n91 ) , .Z( n916 ) , .B( w2_13 ) );
  OAI22_X1 U1274 (.ZN( N118 ) , .A1( n1109 ) , .B2( n1220 ) , .A2( n920 ) , .B1( n921 ) );
  XOR2_X1 U1275 (.Z( n921 ) , .A( n922 ) , .B( n923 ) );
  XOR2_X1 U1276 (.A( n830 ) , .B( n844 ) , .Z( n923 ) );
  XOR2_X1 U1277 (.Z( n844 ) , .A( sa22_sr_3 ) , .B( sa32_sr_3 ) );
  INV_X1 U1278 (.ZN( n830 ) , .A( n924 ) );
  XOR2_X1 U1279 (.B( n817 ) , .Z( n922 ) , .A( n925 ) );
  XNOR2_X1 U1280 (.ZN( n925 ) , .B( sa32_sr_4 ) , .A( w2_12 ) );
  XOR2_X1 U1281 (.A( n89 ) , .Z( n920 ) , .B( w2_12 ) );
  OAI22_X1 U1283 (.ZN( N117 ) , .A1( n1212 ) , .B2( n1220 ) , .A2( n926 ) , .B1( n927 ) );
  XOR2_X1 U1285 (.A( n837 ) , .B( n851 ) , .Z( n929 ) );
  INV_X1 U1287 (.ZN( n837 ) , .A( n930 ) );
  XNOR2_X1 U1289 (.ZN( n931 ) , .B( sa32_sr_3 ) , .A( w2_11 ) );
  XOR2_X1 U1290 (.A( n87 ) , .Z( n926 ) , .B( w2_11 ) );
  OAI22_X1 U1292 (.ZN( N116 ) , .A1( n1213 ) , .B2( n1217 ) , .A2( n932 ) , .B1( n933 ) );
  XOR2_X1 U1294 (.A( n845 ) , .B( n856 ) , .Z( n935 ) );
  XOR2_X1 U1295 (.Z( n856 ) , .A( sa22_sr_1 ) , .B( sa32_sr_1 ) );
  XOR2_X1 U1297 (.A( n85 ) , .Z( n932 ) , .B( w2_10 ) );
  OAI22_X1 U1299 (.ZN( N115 ) , .B2( n1114 ) , .A1( n1216 ) , .A2( n936 ) , .B1( n937 ) );
  XOR2_X1 U1301 (.A( n817 ) , .B( n862 ) , .Z( n939 ) );
  XOR2_X1 U1302 (.Z( n862 ) , .A( sa22_sr_0 ) , .B( sa32_sr_0 ) );
  XOR2_X1 U1304 (.Z( n277 ) , .A( sa02_sr_1 ) , .B( sa12_sr_1 ) );
  XNOR2_X1 U1305 (.ZN( n940 ) , .B( sa32_sr_1 ) , .A( w2_9 ) );
  XOR2_X1 U1306 (.A( n83 ) , .Z( n936 ) , .B( w2_9 ) );
  OAI22_X1 U1308 (.ZN( N114 ) , .B2( n1114 ) , .A1( n1216 ) , .A2( n941 ) , .B1( n942 ) );
  XOR2_X1 U1310 (.A( n284 ) , .B( n817 ) , .Z( n944 ) );
  XOR2_X1 U1311 (.Z( n817 ) , .A( sa22_sr_7 ) , .B( sa32_sr_7 ) );
  XOR2_X1 U1312 (.Z( n284 ) , .A( sa02_sr_0 ) , .B( sa12_sr_0 ) );
  XOR2_X1 U1314 (.A( n81 ) , .Z( n941 ) , .B( w2_8 ) );
  OAI22_X1 U1316 (.ZN( N105 ) , .B2( n1114 ) , .A1( n1216 ) , .A2( n945 ) , .B1( n946 ) );
  XOR2_X1 U1317 (.Z( n946 ) , .A( n947 ) , .B( n948 ) );
  XOR2_X1 U1318 (.B( n836 ) , .Z( n948 ) , .A( sa02_sr_6 ) );
  XOR2_X1 U1319 (.Z( n836 ) , .A( sa02_sr_7 ) , .B( sa12_sr_7 ) );
  XNOR2_X1 U1320 (.ZN( n947 ) , .B( n949 ) , .A( sa22_sr_7 ) );
  XOR2_X1 U1321 (.Z( n949 ) , .B( sa32_sr_6 ) , .A( w2_7 ) );
  XOR2_X1 U1322 (.A( n79 ) , .Z( n945 ) , .B( w2_7 ) );
  OAI22_X1 U1324 (.ZN( N104 ) , .B2( n1114 ) , .A1( n1216 ) , .A2( n950 ) , .B1( n951 ) );
  XOR2_X1 U1327 (.Z( n954 ) , .B( sa32_sr_5 ) , .A( w2_6 ) );
  XNOR2_X1 U1328 (.B( n818 ) , .ZN( n952 ) , .A( sa02_sr_5 ) );
  XOR2_X1 U1329 (.Z( n818 ) , .A( sa02_sr_6 ) , .B( sa12_sr_6 ) );
  XOR2_X1 U1330 (.A( n77 ) , .Z( n950 ) , .B( w2_6 ) );
  XOR2_X1 U1333 (.Z( n956 ) , .A( n957 ) , .B( n958 ) );
  XOR2_X1 U1334 (.Z( n958 ) , .B( n959 ) , .A( sa22_sr_5 ) );
  XOR2_X1 U1335 (.Z( n959 ) , .B( sa32_sr_4 ) , .A( w2_5 ) );
  XNOR2_X1 U1336 (.B( n825 ) , .ZN( n957 ) , .A( sa02_sr_4 ) );
  XOR2_X1 U1337 (.Z( n825 ) , .A( sa02_sr_5 ) , .B( sa12_sr_5 ) );
  OAI22_X1 U1340 (.ZN( N102 ) , .B2( n1114 ) , .A1( n1216 ) , .A2( n960 ) , .B1( n961 ) );
  XOR2_X1 U1343 (.Z( n964 ) , .B( sa32_sr_3 ) , .A( w2_4 ) );
  XOR2_X1 U1344 (.A( n924 ) , .Z( n962 ) , .B( n965 ) );
  XOR2_X1 U1345 (.B( n279 ) , .Z( n965 ) , .A( sa02_sr_3 ) );
  XNOR2_X1 U1346 (.ZN( n924 ) , .A( sa02_sr_4 ) , .B( sa12_sr_4 ) );
  XOR2_X1 U1347 (.A( n73 ) , .Z( n960 ) , .B( w2_4 ) );
  OAI22_X1 U1349 (.ZN( N101 ) , .B2( n1114 ) , .A1( n1216 ) , .A2( n966 ) , .B1( n967 ) );
  XOR2_X1 U1351 (.Z( n969 ) , .B( n970 ) , .A( sa22_sr_3 ) );
  XOR2_X1 U1352 (.Z( n970 ) , .B( sa32_sr_2 ) , .A( w2_3 ) );
  XOR2_X1 U1354 (.B( n279 ) , .Z( n971 ) , .A( sa02_sr_2 ) );
  XOR2_X1 U1355 (.Z( n279 ) , .A( sa02_sr_7 ) , .B( sa32_sr_7 ) );
  XNOR2_X1 U1356 (.ZN( n930 ) , .A( sa02_sr_3 ) , .B( sa12_sr_3 ) );
  XOR2_X1 U1357 (.A( n71 ) , .Z( n966 ) , .B( w2_3 ) );
  OAI22_X1 U1359 (.ZN( N100 ) , .B2( n1114 ) , .A1( n1216 ) , .A2( n972 ) , .B1( n973 ) );
  XOR2_X1 U1361 (.Z( n973 ) , .A( n974 ) , .B( n975 ) );
  XOR2_X1 U1362 (.Z( n975 ) , .B( n976 ) , .A( sa22_sr_2 ) );
  XOR2_X1 U1363 (.Z( n976 ) , .B( sa32_sr_1 ) , .A( w2_2 ) );
  XNOR2_X1 U1364 (.B( n845 ) , .ZN( n974 ) , .A( sa02_sr_1 ) );
  XOR2_X1 U1365 (.Z( n845 ) , .B( sa02_sr_2 ) , .A( sa12_sr_2 ) );
  XOR2_X1 U1366 (.A( n69 ) , .Z( n972 ) , .B( w2_2 ) );
  XOR2_X1 U1374 (.Z( N495 ) , .B( sa32_sr_2 ) , .A( w2_2 ) );
  XNOR2_X1 U1375 (.A( n1117 ) , .B( n885 ) , .ZN( n888 ) );
  XOR2_X1 U1376 (.Z( n1117 ) , .B( n844 ) , .A( sa02_sr_3 ) );
  XNOR2_X1 U1377 (.A( n1118 ) , .B( n539 ) , .ZN( n542 ) );
  XOR2_X1 U1378 (.Z( n1118 ) , .B( n496 ) , .A( sa00_sr_3 ) );
  XNOR2_X1 U1379 (.B( n476 ) , .ZN( n524 ) , .A( sa00_sr_6 ) );
  XNOR2_X1 U1380 (.B( n824 ) , .ZN( n870 ) , .A( sa02_sr_6 ) );
  XNOR2_X1 U1383 (.B( n851 ) , .ZN( n894 ) , .A( sa02_sr_2 ) );
  XNOR2_X1 U1403 (.A( n1126 ) , .ZN( n493 ) , .B( n495 ) );
  XNOR2_X1 U1404 (.ZN( n1126 ) , .B( n488 ) , .A( n498 ) );
  XNOR2_X1 U1405 (.A( n1127 ) , .ZN( n841 ) , .B( n843 ) );
  XNOR2_X1 U1406 (.ZN( n1127 ) , .B( n836 ) , .A( n846 ) );
  XNOR2_X1 U1407 (.A( n1128 ) , .ZN( n933 ) , .B( n935 ) );
  XOR2_X1 U1408 (.Z( n1128 ) , .B( sa32_sr_2 ) , .A( w2_10 ) );
  XNOR2_X1 U1411 (.A( n1130 ) , .ZN( n848 ) , .B( n850 ) );
  XOR2_X1 U1412 (.Z( n1130 ) , .B( sa12_sr_2 ) , .A( w2_26 ) );
  XNOR2_X1 U1415 (.A( n1132 ) , .ZN( n479 ) , .B( n481 ) );
  XOR2_X1 U1416 (.Z( n1132 ) , .B( sa10_sr_5 ) , .A( w0_29 ) );
  XOR2_X1 U1418 (.Z( n1133 ) , .A( n277 ) , .B( n278 ) );
  XNOR2_X1 U1421 (.A( n1135 ) , .ZN( n579 ) , .B( n581 ) );
  XNOR2_X1 U1422 (.ZN( n1135 ) , .B( n469 ) , .A( n582 ) );
  XNOR2_X1 U1423 (.A( n1136 ) , .ZN( n814 ) , .B( n816 ) );
  XNOR2_X1 U1424 (.ZN( n1136 ) , .B( n819 ) , .A( w2_31 ) );
  XNOR2_X1 U1427 (.A( n1138 ) , .ZN( n927 ) , .B( n929 ) );
  XNOR2_X1 U1428 (.ZN( n1138 ) , .B( n817 ) , .A( n931 ) );
  XNOR2_X1 U1429 (.B( n1139 ) , .ZN( n893 ) , .A( n894 ) );
  XNOR2_X1 U1430 (.ZN( n1139 ) , .B( n896 ) , .A( sa12_sr_1 ) );
  XNOR2_X1 U1439 (.A( n1144 ) , .ZN( n500 ) , .B( n502 ) );
  XOR2_X1 U1440 (.Z( n1144 ) , .B( sa10_sr_2 ) , .A( w0_26 ) );
  XNOR2_X1 U1441 (.A( n1145 ) , .ZN( n967 ) , .B( n969 ) );
  XNOR2_X1 U1442 (.ZN( n1145 ) , .A( n930 ) , .B( n971 ) );
  XNOR2_X1 U1447 (.A( n1148 ) , .ZN( n281 ) , .B( n283 ) );
  XOR2_X1 U1448 (.Z( n1148 ) , .B( sa22_sr_0 ) , .A( w2_0 ) );
  XNOR2_X1 U1449 (.B( n1149 ) , .ZN( n619 ) , .A( n620 ) );
  XNOR2_X1 U1450 (.ZN( n1149 ) , .B( n622 ) , .A( sa20_sr_3 ) );
  XNOR2_X1 U1451 (.A( n1150 ) , .ZN( n937 ) , .B( n939 ) );
  XNOR2_X1 U1452 (.ZN( n1150 ) , .B( n277 ) , .A( n940 ) );
  XNOR2_X1 U1453 (.A( n1151 ) , .ZN( n859 ) , .B( n861 ) );
  XOR2_X1 U1454 (.Z( n1151 ) , .B( sa12_sr_0 ) , .A( w2_24 ) );
  XNOR2_X1 U1457 (.A( n1153 ) , .ZN( n562 ) , .B( n564 ) );
  XOR2_X1 U1458 (.Z( n1153 ) , .B( sa30_sr_7 ) , .A( w0_15 ) );
  XNOR2_X1 U1459 (.A( n1154 ) , .ZN( n909 ) , .B( n911 ) );
  XOR2_X1 U1460 (.Z( n1154 ) , .B( sa32_sr_7 ) , .A( w2_15 ) );
  XNOR2_X1 U1461 (.A( n1155 ) , .ZN( n473 ) , .B( n475 ) );
  XOR2_X1 U1462 (.Z( n1155 ) , .B( sa10_sr_6 ) , .A( w0_30 ) );
  XNOR2_X1 U1463 (.A( n1156 ) , .ZN( n821 ) , .B( n823 ) );
  XOR2_X1 U1464 (.Z( n1156 ) , .B( sa12_sr_6 ) , .A( w2_30 ) );
  XNOR2_X1 U1467 (.A( n1158 ) , .ZN( n588 ) , .B( n590 ) );
  XNOR2_X1 U1468 (.ZN( n1158 ) , .B( n469 ) , .A( n591 ) );
  XNOR2_X1 U1471 (.B( n1160 ) , .ZN( n523 ) , .A( n524 ) );
  XNOR2_X1 U1472 (.ZN( n1160 ) , .B( n526 ) , .A( sa10_sr_5 ) );
  XNOR2_X1 U1479 (.A( n1164 ) , .ZN( n913 ) , .B( n915 ) );
  XOR2_X1 U1480 (.Z( n1164 ) , .B( sa32_sr_6 ) , .A( w2_14 ) );
  XNOR2_X1 U1487 (.A( n1168 ) , .ZN( n942 ) , .B( n944 ) );
  XOR2_X1 U1488 (.Z( n1168 ) , .B( sa32_sr_0 ) , .A( w2_8 ) );
  XNOR2_X1 U1495 (.B( n1172 ) , .ZN( n853 ) , .A( n854 ) );
  XNOR2_X1 U1496 (.ZN( n1172 ) , .A( n836 ) , .B( n856 ) );
  XNOR2_X1 U1497 (.A( n1173 ) , .ZN( n905 ) , .B( n907 ) );
  XOR2_X1 U1498 (.Z( n1173 ) , .B( sa02_sr_0 ) , .A( w2_16 ) );
  XNOR2_X1 U1507 (.B( n1178 ) , .ZN( n625 ) , .A( n626 ) );
  XNOR2_X1 U1508 (.ZN( n1178 ) , .B( n628 ) , .A( sa20_sr_2 ) );
  XNOR2_X1 U1509 (.B( n1179 ) , .ZN( n547 ) , .A( n548 ) );
  XNOR2_X1 U1510 (.ZN( n1179 ) , .B( n550 ) , .A( sa10_sr_1 ) );
  XNOR2_X1 U1513 (.B( n1181 ) , .ZN( n961 ) , .A( n962 ) );
  XNOR2_X1 U1514 (.ZN( n1181 ) , .B( n964 ) , .A( sa22_sr_4 ) );
  XNOR2_X1 U1517 (.A( n1183 ) , .ZN( n552 ) , .B( n554 ) );
  XNOR2_X1 U1518 (.ZN( n1183 ) , .B( n539 ) , .A( n556 ) );
  XNOR2_X1 U1523 (.B( n1186 ) , .ZN( n951 ) , .A( n952 ) );
  XNOR2_X1 U1524 (.ZN( n1186 ) , .B( n954 ) , .A( sa22_sr_6 ) );
  XNOR2_X1 U1527 (.A( n1188 ) , .ZN( n630 ) , .B( n632 ) );
  XNOR2_X1 U1528 (.ZN( n1188 ) , .B( n617 ) , .A( n634 ) );
  XNOR2_X1 U1539 (.A( n1194 ) , .ZN( n593 ) , .B( n595 ) );
  XOR2_X1 U1540 (.Z( n1194 ) , .B( sa30_sr_0 ) , .A( w0_8 ) );
  XNOR2_X1 U1543 (.A( n1196 ) , .ZN( n584 ) , .B( n586 ) );
  XOR2_X1 U1544 (.Z( n1196 ) , .B( sa30_sr_2 ) , .A( w0_10 ) );
  XNOR2_X1 U1559 (.A( n1204 ) , .ZN( n636 ) , .B( n638 ) );
  XOR2_X1 U1560 (.Z( n1204 ) , .B( sa20_sr_0 ) , .A( w0_0 ) );
  XNOR2_X1 U1563 (.ZN( N415 ) , .B( n1206 ) , .A( w0_18 ) );
  XNOR2_X1 U1564 (.ZN( N463 ) , .B( n1208 ) , .A( w2_10 ) );
  INV_X1 U1567 (.ZN( n1206 ) , .A( sa10_sr_2 ) );
  NAND2_X1 U1569 (.A2( n1209 ) , .ZN( n1210 ) , .A1( sa22_sr_2 ) );
  NAND2_X1 U1570 (.A1( n1208 ) , .ZN( n1211 ) , .A2( sa32_sr_2 ) );
  NAND2_X1 U1571 (.A1( n1210 ) , .A2( n1211 ) , .ZN( n851 ) );
  INV_X1 U1572 (.ZN( n1208 ) , .A( sa22_sr_2 ) );
  INV_X1 U1573 (.ZN( n1209 ) , .A( sa32_sr_2 ) );
  XOR2_X1 U281 (.Z( n278 ) , .B( n279 ) , .A( sa02_sr_0 ) );
  OAI22_X1 U284 (.ZN( N98 ) , .A1( n1215 ) , .B2( n1220 ) , .A2( n280 ) , .B1( n281 ) );
  XOR2_X1 U286 (.A( n279 ) , .Z( n283 ) , .B( n284 ) );
  XOR2_X1 U288 (.Z( n280 ) , .A( n65 ) , .B( w2_0 ) );
  XOR2_X1 U471 (.Z( N494 ) , .B( sa32_sr_3 ) , .A( w2_3 ) );
  XOR2_X1 U472 (.Z( N493 ) , .B( sa32_sr_4 ) , .A( w2_4 ) );
  XOR2_X1 U473 (.Z( N492 ) , .B( sa32_sr_5 ) , .A( w2_5 ) );
  XOR2_X1 U474 (.Z( N491 ) , .B( sa32_sr_6 ) , .A( w2_6 ) );
  XOR2_X1 U475 (.Z( N490 ) , .B( sa32_sr_7 ) , .A( w2_7 ) );
  XOR2_X1 U484 (.Z( N481 ) , .B( sa30_sr_0 ) , .A( w0_0 ) );
  XOR2_X1 U485 (.Z( N480 ) , .B( sa30_sr_1 ) , .A( w0_1 ) );
  XOR2_X1 U486 (.Z( N479 ) , .B( sa30_sr_2 ) , .A( w0_2 ) );
  XOR2_X1 U487 (.Z( N478 ) , .B( sa30_sr_3 ) , .A( w0_3 ) );
  XOR2_X1 U488 (.Z( N477 ) , .B( sa30_sr_4 ) , .A( w0_4 ) );
  XOR2_X1 U491 (.Z( N474 ) , .B( sa30_sr_7 ) , .A( w0_7 ) );
  XOR2_X1 U500 (.Z( N465 ) , .B( sa22_sr_0 ) , .A( w2_8 ) );
  XOR2_X1 U501 (.Z( N464 ) , .B( sa22_sr_1 ) , .A( w2_9 ) );
  XOR2_X1 U503 (.Z( N462 ) , .B( sa22_sr_3 ) , .A( w2_11 ) );
  XOR2_X1 U504 (.Z( N461 ) , .B( sa22_sr_4 ) , .A( w2_12 ) );
  XOR2_X1 U506 (.Z( N459 ) , .B( sa22_sr_6 ) , .A( w2_14 ) );
  XOR2_X1 U507 (.Z( N458 ) , .B( sa22_sr_7 ) , .A( w2_15 ) );
  XOR2_X1 U516 (.Z( N449 ) , .B( sa20_sr_0 ) , .A( w0_8 ) );
  XOR2_X1 U517 (.Z( N448 ) , .B( sa20_sr_1 ) , .A( w0_9 ) );
  XOR2_X1 U518 (.Z( N447 ) , .B( sa20_sr_2 ) , .A( w0_10 ) );
  XOR2_X1 U519 (.Z( N446 ) , .B( sa20_sr_3 ) , .A( w0_11 ) );
  XOR2_X1 U520 (.Z( N445 ) , .B( sa20_sr_4 ) , .A( w0_12 ) );
  XOR2_X1 U521 (.Z( N444 ) , .B( sa20_sr_5 ) , .A( w0_13 ) );
  XOR2_X1 U523 (.Z( N442 ) , .B( sa20_sr_7 ) , .A( w0_15 ) );
  XOR2_X1 U532 (.Z( N433 ) , .B( sa12_sr_0 ) , .A( w2_16 ) );
  XOR2_X1 U533 (.Z( N432 ) , .B( sa12_sr_1 ) , .A( w2_17 ) );
  XOR2_X1 U534 (.Z( N431 ) , .B( sa12_sr_2 ) , .A( w2_18 ) );
  XOR2_X1 U535 (.Z( N430 ) , .B( sa12_sr_3 ) , .A( w2_19 ) );
  XOR2_X1 U536 (.Z( N429 ) , .B( sa12_sr_4 ) , .A( w2_20 ) );
  XOR2_X1 U539 (.Z( N426 ) , .B( sa12_sr_7 ) , .A( w2_23 ) );
  XOR2_X1 U549 (.Z( N416 ) , .B( sa10_sr_1 ) , .A( w0_17 ) );
  XOR2_X1 U551 (.Z( N414 ) , .B( sa10_sr_3 ) , .A( w0_19 ) );
  XOR2_X1 U552 (.Z( N413 ) , .B( sa10_sr_4 ) , .A( w0_20 ) );
  XOR2_X1 U553 (.Z( N412 ) , .B( sa10_sr_5 ) , .A( w0_21 ) );
  XOR2_X1 U554 (.Z( N411 ) , .B( sa10_sr_6 ) , .A( w0_22 ) );
  XOR2_X1 U573 (.Z( N401 ) , .B( sa02_sr_0 ) , .A( w2_24 ) );
  XOR2_X1 U574 (.Z( N400 ) , .B( sa02_sr_1 ) , .A( w2_25 ) );
  XOR2_X1 U584 (.Z( N399 ) , .B( sa02_sr_2 ) , .A( w2_26 ) );
  XOR2_X1 U585 (.Z( N398 ) , .B( sa02_sr_3 ) , .A( w2_27 ) );
  XOR2_X1 U586 (.Z( N397 ) , .B( sa02_sr_4 ) , .A( w2_28 ) );
  XOR2_X1 U587 (.Z( N396 ) , .B( sa02_sr_5 ) , .A( w2_29 ) );
  XOR2_X1 U588 (.Z( N395 ) , .B( sa02_sr_6 ) , .A( w2_30 ) );
  XOR2_X1 U589 (.Z( N394 ) , .B( sa02_sr_7 ) , .A( w2_31 ) );
  XOR2_X1 U609 (.Z( N383 ) , .B( sa00_sr_2 ) , .A( w0_26 ) );
  XOR2_X1 U610 (.Z( N382 ) , .B( sa00_sr_3 ) , .A( w0_27 ) );
  XOR2_X1 U611 (.Z( N381 ) , .B( sa00_sr_4 ) , .A( w0_28 ) );
  XOR2_X1 U612 (.Z( N380 ) , .B( sa00_sr_5 ) , .A( w0_29 ) );
  XOR2_X1 U623 (.Z( N379 ) , .B( sa00_sr_6 ) , .A( w0_30 ) );
  OAI22_X1 U669 (.ZN( N280 ) , .B2( n1114 ) , .A1( n1214 ) , .A2( n472 ) , .B1( n473 ) );
  XOR2_X1 U671 (.Z( n475 ) , .A( n476 ) , .B( n477 ) );
  XOR2_X1 U673 (.A( n253 ) , .Z( n472 ) , .B( w0_30 ) );
  OAI22_X1 U675 (.ZN( N279 ) , .A1( n1212 ) , .B2( n1218 ) , .A2( n478 ) , .B1( n479 ) );
  XOR2_X1 U677 (.Z( n481 ) , .A( n482 ) , .B( n483 ) );
  XOR2_X1 U679 (.A( n251 ) , .Z( n478 ) , .B( w0_29 ) );
  XOR2_X1 U682 (.Z( n485 ) , .A( n486 ) , .B( n487 ) );
  XOR2_X1 U683 (.Z( n487 ) , .A( n488 ) , .B( n489 ) );
  XOR2_X1 U684 (.Z( n486 ) , .A( n490 ) , .B( n491 ) );
  XNOR2_X1 U685 (.ZN( n490 ) , .B( sa10_sr_4 ) , .A( w0_28 ) );
  OAI22_X1 U688 (.ZN( N277 ) , .A1( n1212 ) , .B2( n1219 ) , .A2( n492 ) , .B1( n493 ) );
  XOR2_X1 U690 (.Z( n495 ) , .A( n496 ) , .B( n497 ) );
  XNOR2_X1 U692 (.ZN( n498 ) , .B( sa10_sr_3 ) , .A( w0_27 ) );
  XOR2_X1 U693 (.A( n247 ) , .Z( n492 ) , .B( w0_27 ) );
  OAI22_X1 U695 (.ZN( N276 ) , .A1( n1212 ) , .B2( n1220 ) , .A2( n499 ) , .B1( n500 ) );
  XOR2_X1 U697 (.Z( n502 ) , .A( n503 ) , .B( n504 ) );
  XOR2_X1 U699 (.A( n245 ) , .Z( n499 ) , .B( w0_26 ) );
  XOR2_X1 U703 (.Z( n508 ) , .A( n509 ) , .B( n510 ) );
  XOR2_X1 U710 (.A( n488 ) , .Z( n515 ) , .B( n516 ) );
  OAI22_X1 U721 (.ZN( N264 ) , .A1( n1213 ) , .B2( n1220 ) , .A2( n522 ) , .B1( n523 ) );
  XOR2_X1 U724 (.Z( n526 ) , .B( sa20_sr_5 ) , .A( w0_22 ) );
  XOR2_X1 U727 (.A( n237 ) , .Z( n522 ) , .B( w0_22 ) );
  OAI22_X1 U729 (.ZN( N263 ) , .A1( n1213 ) , .B2( n1221 ) , .A2( n528 ) , .B1( n529 ) );
  XOR2_X1 U730 (.Z( n529 ) , .A( n530 ) , .B( n531 ) );
  XOR2_X1 U731 (.Z( n531 ) , .B( n532 ) , .A( sa10_sr_4 ) );
  XOR2_X1 U732 (.Z( n532 ) , .B( sa20_sr_4 ) , .A( w0_21 ) );
  XNOR2_X1 U733 (.B( n482 ) , .ZN( n530 ) , .A( sa00_sr_5 ) );
  XOR2_X1 U734 (.A( n235 ) , .Z( n528 ) , .B( w0_21 ) );
  OAI22_X1 U736 (.ZN( N262 ) , .A1( n1213 ) , .B2( n1218 ) , .A2( n533 ) , .B1( n534 ) );
  XOR2_X1 U737 (.Z( n534 ) , .A( n535 ) , .B( n536 ) );
  XOR2_X1 U738 (.Z( n536 ) , .B( n537 ) , .A( sa10_sr_3 ) );
  XOR2_X1 U739 (.Z( n537 ) , .B( sa20_sr_3 ) , .A( w0_20 ) );
  XOR2_X1 U740 (.Z( n535 ) , .A( n538 ) , .B( n539 ) );
  XNOR2_X1 U741 (.B( n491 ) , .ZN( n538 ) , .A( sa00_sr_4 ) );
  XOR2_X1 U742 (.A( n233 ) , .Z( n533 ) , .B( w0_20 ) );
  OAI22_X1 U744 (.ZN( N261 ) , .A1( n1213 ) , .B2( n1220 ) , .A2( n540 ) , .B1( n541 ) );
  XOR2_X1 U745 (.Z( n541 ) , .A( n542 ) , .B( n543 ) );
  XOR2_X1 U746 (.Z( n543 ) , .B( n544 ) , .A( sa10_sr_2 ) );
  XOR2_X1 U747 (.Z( n544 ) , .B( sa20_sr_2 ) , .A( w0_19 ) );
  XOR2_X1 U750 (.A( n231 ) , .Z( n540 ) , .B( w0_19 ) );
  OAI22_X1 U752 (.ZN( N260 ) , .A1( n1213 ) , .B2( n1218 ) , .A2( n546 ) , .B1( n547 ) );
  XOR2_X1 U755 (.Z( n550 ) , .B( sa20_sr_1 ) , .A( w0_18 ) );
  XNOR2_X1 U756 (.B( n503 ) , .ZN( n548 ) , .A( sa00_sr_2 ) );
  XOR2_X1 U757 (.A( n229 ) , .Z( n546 ) , .B( w0_18 ) );
  OAI22_X1 U759 (.ZN( N259 ) , .A1( n1109 ) , .B2( n1218 ) , .A2( n551 ) , .B1( n552 ) );
  XOR2_X1 U761 (.Z( n554 ) , .B( n555 ) , .A( sa10_sr_0 ) );
  XOR2_X1 U762 (.Z( n555 ) , .B( sa20_sr_0 ) , .A( w0_17 ) );
  XNOR2_X1 U764 (.B( n509 ) , .ZN( n556 ) , .A( sa00_sr_1 ) );
  XOR2_X1 U765 (.A( n227 ) , .Z( n551 ) , .B( w0_17 ) );
  XOR2_X1 U769 (.A( n516 ) , .B( n539 ) , .Z( n560 ) );
  XOR2_X1 U770 (.Z( n539 ) , .A( sa10_sr_7 ) , .B( sa20_sr_7 ) );
  OAI22_X1 U774 (.ZN( N249 ) , .A1( n1109 ) , .B2( n1217 ) , .A2( n561 ) , .B1( n562 ) );
  XOR2_X1 U776 (.A( n476 ) , .B( n488 ) , .Z( n564 ) );
  XOR2_X1 U777 (.Z( n476 ) , .A( sa20_sr_6 ) , .B( sa30_sr_6 ) );
  XOR2_X1 U779 (.A( n223 ) , .Z( n561 ) , .B( w0_15 ) );
  OAI22_X1 U788 (.ZN( N247 ) , .A1( n1212 ) , .B2( n1221 ) , .A2( n569 ) , .B1( n570 ) );
  XOR2_X1 U789 (.Z( n570 ) , .A( n571 ) , .B( n572 ) );
  XOR2_X1 U790 (.A( n477 ) , .B( n491 ) , .Z( n572 ) );
  XOR2_X1 U791 (.Z( n491 ) , .A( sa20_sr_4 ) , .B( sa30_sr_4 ) );
  XNOR2_X1 U792 (.ZN( n571 ) , .B( sa30_sr_5 ) , .A( w0_13 ) );
  XOR2_X1 U793 (.A( n219 ) , .Z( n569 ) , .B( w0_13 ) );
  OAI22_X1 U795 (.ZN( N246 ) , .A1( n1213 ) , .B2( n1217 ) , .A2( n573 ) , .B1( n574 ) );
  XOR2_X1 U796 (.Z( n574 ) , .A( n575 ) , .B( n576 ) );
  XOR2_X1 U797 (.A( n483 ) , .B( n496 ) , .Z( n576 ) );
  XOR2_X1 U798 (.Z( n496 ) , .A( sa20_sr_3 ) , .B( sa30_sr_3 ) );
  XOR2_X1 U799 (.B( n469 ) , .Z( n575 ) , .A( n577 ) );
  XNOR2_X1 U800 (.ZN( n577 ) , .B( sa30_sr_4 ) , .A( w0_12 ) );
  XOR2_X1 U801 (.A( n217 ) , .Z( n573 ) , .B( w0_12 ) );
  OAI22_X1 U803 (.ZN( N245 ) , .B2( n1114 ) , .A1( n1216 ) , .A2( n578 ) , .B1( n579 ) );
  XOR2_X1 U805 (.A( n489 ) , .B( n503 ) , .Z( n581 ) );
  XOR2_X1 U806 (.Z( n503 ) , .A( sa20_sr_2 ) , .B( sa30_sr_2 ) );
  XNOR2_X1 U808 (.ZN( n582 ) , .B( sa30_sr_3 ) , .A( w0_11 ) );
  XOR2_X1 U809 (.A( n215 ) , .Z( n578 ) , .B( w0_11 ) );
  OAI22_X1 U811 (.ZN( N244 ) , .A1( n1212 ) , .B2( n1220 ) , .A2( n583 ) , .B1( n584 ) );
  XOR2_X1 U813 (.A( n497 ) , .B( n509 ) , .Z( n586 ) );
  XOR2_X1 U814 (.Z( n509 ) , .A( sa20_sr_1 ) , .B( sa30_sr_1 ) );
  XOR2_X1 U816 (.A( n213 ) , .Z( n583 ) , .B( w0_10 ) );
  OAI22_X1 U818 (.ZN( N243 ) , .A1( n1212 ) , .B2( n1220 ) , .A2( n587 ) , .B1( n588 ) );
  XOR2_X1 U820 (.A( n504 ) , .B( n516 ) , .Z( n590 ) );
  XOR2_X1 U821 (.Z( n516 ) , .A( sa20_sr_0 ) , .B( sa30_sr_0 ) );
  XNOR2_X1 U823 (.ZN( n591 ) , .B( sa30_sr_1 ) , .A( w0_9 ) );
  XOR2_X1 U824 (.A( n211 ) , .Z( n587 ) , .B( w0_9 ) );
  OAI22_X1 U826 (.ZN( N242 ) , .A1( n1215 ) , .B2( n1220 ) , .A2( n592 ) , .B1( n593 ) );
  XOR2_X1 U828 (.A( n469 ) , .B( n510 ) , .Z( n595 ) );
  XOR2_X1 U829 (.Z( n469 ) , .A( sa20_sr_7 ) , .B( sa30_sr_7 ) );
  XOR2_X1 U831 (.A( n209 ) , .Z( n592 ) , .B( w0_8 ) );
  OAI22_X1 U833 (.ZN( N233 ) , .A1( n1213 ) , .B2( n1221 ) , .A2( n596 ) , .B1( n597 ) );
  XOR2_X1 U834 (.Z( n597 ) , .A( n598 ) , .B( n599 ) );
  XOR2_X1 U835 (.B( n488 ) , .Z( n599 ) , .A( sa00_sr_6 ) );
  XNOR2_X1 U837 (.ZN( n598 ) , .B( n600 ) , .A( sa20_sr_7 ) );
  XOR2_X1 U838 (.Z( n600 ) , .B( sa30_sr_6 ) , .A( w0_7 ) );
  XOR2_X1 U839 (.A( n207 ) , .Z( n596 ) , .B( w0_7 ) );
  OAI22_X1 U849 (.ZN( N231 ) , .A1( n1109 ) , .B2( n1217 ) , .A2( n606 ) , .B1( n607 ) );
  XOR2_X1 U850 (.Z( n607 ) , .A( n608 ) , .B( n609 ) );
  XOR2_X1 U851 (.Z( n609 ) , .B( n610 ) , .A( sa20_sr_5 ) );
  XOR2_X1 U852 (.Z( n610 ) , .B( sa30_sr_4 ) , .A( w0_5 ) );
  XNOR2_X1 U853 (.B( n477 ) , .ZN( n608 ) , .A( sa00_sr_4 ) );
  XOR2_X1 U854 (.Z( n477 ) , .A( sa00_sr_5 ) , .B( sa10_sr_5 ) );
  XOR2_X1 U855 (.A( n203 ) , .Z( n606 ) , .B( w0_5 ) );
  OAI22_X1 U857 (.ZN( N230 ) , .A1( n1109 ) , .B2( n1217 ) , .A2( n611 ) , .B1( n612 ) );
  XOR2_X1 U858 (.Z( n612 ) , .A( n613 ) , .B( n614 ) );
  XOR2_X1 U859 (.Z( n614 ) , .B( n615 ) , .A( sa20_sr_4 ) );
  XOR2_X1 U860 (.Z( n615 ) , .B( sa30_sr_3 ) , .A( w0_4 ) );
  XOR2_X1 U861 (.Z( n613 ) , .A( n616 ) , .B( n617 ) );
  XNOR2_X1 U862 (.B( n483 ) , .ZN( n616 ) , .A( sa00_sr_3 ) );
  XOR2_X1 U863 (.Z( n483 ) , .A( sa00_sr_4 ) , .B( sa10_sr_4 ) );
  XOR2_X1 U864 (.A( n201 ) , .Z( n611 ) , .B( w0_4 ) );
  OAI22_X1 U868 (.ZN( N229 ) , .A1( n1109 ) , .B2( n1217 ) , .A2( n618 ) , .B1( n619 ) );
  XOR2_X1 U871 (.Z( n622 ) , .B( sa30_sr_2 ) , .A( w0_3 ) );
  XOR2_X1 U872 (.B( n617 ) , .Z( n620 ) , .A( n623 ) );
  XNOR2_X1 U873 (.B( n489 ) , .ZN( n623 ) , .A( sa00_sr_2 ) );
  XOR2_X1 U874 (.Z( n489 ) , .A( sa00_sr_3 ) , .B( sa10_sr_3 ) );
  XOR2_X1 U875 (.A( n199 ) , .Z( n618 ) , .B( w0_3 ) );
  OAI22_X1 U877 (.ZN( N228 ) , .A1( n1109 ) , .B2( n1217 ) , .A2( n624 ) , .B1( n625 ) );
  XOR2_X1 U880 (.Z( n628 ) , .B( sa30_sr_1 ) , .A( w0_2 ) );
  XNOR2_X1 U881 (.B( n497 ) , .ZN( n626 ) , .A( sa00_sr_1 ) );
  XOR2_X1 U882 (.Z( n497 ) , .A( sa00_sr_2 ) , .B( sa10_sr_2 ) );
  XOR2_X1 U883 (.A( n197 ) , .Z( n624 ) , .B( w0_2 ) );
  XOR2_X1 U887 (.Z( n632 ) , .B( n633 ) , .A( sa20_sr_1 ) );
  XOR2_X1 U888 (.Z( n633 ) , .B( sa30_sr_0 ) , .A( w0_1 ) );
  XNOR2_X1 U890 (.B( n504 ) , .ZN( n634 ) , .A( sa00_sr_0 ) );
  XOR2_X1 U891 (.Z( n504 ) , .A( sa00_sr_1 ) , .B( sa10_sr_1 ) );
  OAI22_X1 U894 (.ZN( N226 ) , .A1( n1109 ) , .B2( n1217 ) , .A2( n635 ) , .B1( n636 ) );
  XOR2_X1 U896 (.A( n510 ) , .B( n617 ) , .Z( n638 ) );
  XOR2_X1 U897 (.Z( n617 ) , .A( sa00_sr_7 ) , .B( sa30_sr_7 ) );
  XOR2_X1 U898 (.Z( n510 ) , .A( sa00_sr_0 ) , .B( sa10_sr_0 ) );
  XOR2_X1 U900 (.A( n193 ) , .Z( n635 ) , .B( w0_0 ) );
  XNOR2_X1 u0_U10 (.ZN( u0_n57 ) , .B( u0_subword_3 ) , .A( w0_3 ) );
  XNOR2_X1 u0_U17 (.ZN( u0_n53 ) , .B( u0_subword_5 ) , .A( w0_5 ) );
  XNOR2_X1 u0_U183 (.ZN( u0_n61 ) , .B( u0_subword_1 ) , .A( w0_1 ) );
  XNOR2_X1 u0_U185 (.ZN( u0_n55 ) , .B( u0_subword_4 ) , .A( w0_4 ) );
  XNOR2_X1 u0_U21 (.ZN( u0_n49 ) , .B( u0_subword_7 ) , .A( w0_7 ) );
  XNOR2_X1 u0_U212 (.ZN( u0_n59 ) , .A( u0_subword_2 ) , .B( w0_2 ) );
  XNOR2_X1 u0_U248 (.ZN( u0_n63 ) , .B( u0_subword_0 ) , .A( w0_0 ) );
  XNOR2_X1 u0_U259 (.ZN( u0_n51 ) , .B( u0_subword_6 ) , .A( w0_6 ) );
  XOR2_X1 u0_U291 (.Z( u0_n65 ) , .A( u0_n67 ) , .B( w3_31 ) );
  XOR2_X1 u0_U292 (.Z( u0_n68 ) , .A( u0_n70 ) , .B( w3_30 ) );
  XOR2_X1 u0_U293 (.Z( u0_n71 ) , .A( u0_n73 ) , .B( w3_29 ) );
  XOR2_X1 u0_U294 (.Z( u0_n74 ) , .A( u0_n76 ) , .B( w3_28 ) );
  XOR2_X1 u0_U295 (.Z( u0_n77 ) , .A( u0_n79 ) , .B( w3_27 ) );
  XOR2_X1 u0_U297 (.Z( u0_n83 ) , .A( u0_n85 ) , .B( w3_25 ) );
  XOR2_X1 u0_U323 (.A( u0_n162 ) , .Z( u0_n67 ) , .B( w2_31 ) );
  XOR2_X1 u0_U324 (.A( u0_n164 ) , .Z( u0_n70 ) , .B( w2_30 ) );
  XOR2_X1 u0_U325 (.A( u0_n166 ) , .Z( u0_n73 ) , .B( w2_29 ) );
  XOR2_X1 u0_U326 (.A( u0_n168 ) , .Z( u0_n76 ) , .B( w2_28 ) );
  XOR2_X1 u0_U327 (.A( u0_n170 ) , .Z( u0_n79 ) , .B( w2_27 ) );
  XOR2_X1 u0_U329 (.A( u0_n174 ) , .Z( u0_n85 ) , .B( w2_25 ) );
  XOR2_X1 u0_U347 (.Z( u0_n139 ) , .A( u0_n210 ) , .B( w2_7 ) );
  XOR2_X1 u0_U348 (.Z( u0_n142 ) , .A( u0_n212 ) , .B( w2_6 ) );
  XOR2_X1 u0_U351 (.Z( u0_n151 ) , .A( u0_n218 ) , .B( w2_3 ) );
  XOR2_X1 u0_U403 (.Z( u0_n210 ) , .A( u0_n49 ) , .B( w1_7 ) );
  XOR2_X1 u0_U405 (.Z( u0_n212 ) , .A( u0_n51 ) , .B( w1_6 ) );
  XOR2_X1 u0_U411 (.Z( u0_n218 ) , .A( u0_n57 ) , .B( w1_3 ) );
  NOR2_X1 u0_u3_U10 (.ZN( u0_u3_n578 ) , .A1( u0_u3_n625 ) , .A2( u0_u3_n748 ) );
  NOR2_X1 u0_u3_U100 (.ZN( u0_u3_n669 ) , .A1( u0_u3_n731 ) , .A2( u0_u3_n806 ) );
  NOR2_X1 u0_u3_U101 (.ZN( u0_u3_n535 ) , .A2( u0_u3_n752 ) , .A1( u0_u3_n753 ) );
  NOR2_X1 u0_u3_U102 (.A2( u0_u3_n711 ) , .A1( u0_u3_n765 ) , .ZN( u0_u3_n797 ) );
  OAI22_X1 u0_u3_U103 (.B1( u0_u3_n493 ) , .ZN( u0_u3_n494 ) , .A1( u0_u3_n689 ) , .A2( u0_u3_n766 ) , .B2( u0_u3_n820 ) );
  NOR3_X1 u0_u3_U104 (.ZN( u0_u3_n493 ) , .A1( u0_u3_n785 ) , .A2( u0_u3_n852 ) , .A3( u0_u3_n865 ) );
  NOR2_X1 u0_u3_U105 (.ZN( u0_u3_n509 ) , .A2( u0_u3_n731 ) , .A1( u0_u3_n765 ) );
  NOR2_X1 u0_u3_U106 (.ZN( u0_u3_n520 ) , .A1( u0_u3_n711 ) , .A2( u0_u3_n806 ) );
  OAI21_X1 u0_u3_U107 (.ZN( u0_u3_n734 ) , .A( u0_u3_n836 ) , .B2( u0_u3_n854 ) , .B1( u0_u3_n875 ) );
  NOR2_X1 u0_u3_U108 (.ZN( u0_u3_n604 ) , .A2( u0_u3_n783 ) , .A1( u0_u3_n806 ) );
  NOR2_X1 u0_u3_U109 (.A2( u0_u3_n711 ) , .A1( u0_u3_n753 ) , .ZN( u0_u3_n774 ) );
  NOR2_X1 u0_u3_U11 (.A1( u0_u3_n681 ) , .ZN( u0_u3_n696 ) , .A2( u0_u3_n810 ) );
  NOR2_X1 u0_u3_U110 (.A2( u0_u3_n438 ) , .ZN( u0_u3_n670 ) , .A1( u0_u3_n753 ) );
  BUF_X2 u0_u3_U111 (.Z( u0_u3_n439 ) , .A( u0_u3_n794 ) );
  OAI21_X1 u0_u3_U112 (.ZN( u0_u3_n790 ) , .A( u0_u3_n841 ) , .B1( u0_u3_n865 ) , .B2( u0_u3_n875 ) );
  BUF_X2 u0_u3_U113 (.Z( u0_u3_n41 ) , .A( u0_u3_n700 ) );
  NOR2_X1 u0_u3_U114 (.ZN( u0_u3_n632 ) , .A2( u0_u3_n731 ) , .A1( u0_u3_n788 ) );
  NOR2_X1 u0_u3_U115 (.ZN( u0_u3_n512 ) , .A1( u0_u3_n732 ) , .A2( u0_u3_n782 ) );
  NOR2_X1 u0_u3_U116 (.ZN( u0_u3_n510 ) , .A1( u0_u3_n815 ) , .A2( u0_u3_n820 ) );
  NOR2_X1 u0_u3_U117 (.ZN( u0_u3_n666 ) , .A1( u0_u3_n732 ) , .A2( u0_u3_n788 ) );
  NOR2_X1 u0_u3_U118 (.ZN( u0_u3_n546 ) , .A2( u0_u3_n711 ) , .A1( u0_u3_n788 ) );
  NOR2_X1 u0_u3_U119 (.ZN( u0_u3_n511 ) , .A2( u0_u3_n783 ) , .A1( u0_u3_n788 ) );
  INV_X1 u0_u3_U12 (.A( u0_u3_n683 ) , .ZN( u0_u3_n842 ) );
  NOR2_X1 u0_u3_U120 (.ZN( u0_u3_n547 ) , .A2( u0_u3_n788 ) , .A1( u0_u3_n795 ) );
  NOR2_X1 u0_u3_U121 (.ZN( u0_u3_n685 ) , .A2( u0_u3_n711 ) , .A1( u0_u3_n820 ) );
  AOI21_X1 u0_u3_U122 (.ZN( u0_u3_n572 ) , .B1( u0_u3_n753 ) , .B2( u0_u3_n765 ) , .A( u0_u3_n783 ) );
  NOR2_X1 u0_u3_U123 (.ZN( u0_u3_n714 ) , .A1( u0_u3_n765 ) , .A2( u0_u3_n766 ) );
  NOR2_X1 u0_u3_U124 (.ZN( u0_u3_n532 ) , .A1( u0_u3_n711 ) , .A2( u0_u3_n782 ) );
  AOI21_X1 u0_u3_U125 (.ZN( u0_u3_n518 ) , .A( u0_u3_n732 ) , .B1( u0_u3_n753 ) , .B2( u0_u3_n806 ) );
  NOR2_X1 u0_u3_U126 (.ZN( u0_u3_n617 ) , .A1( u0_u3_n765 ) , .A2( u0_u3_n815 ) );
  INV_X1 u0_u3_U127 (.A( u0_u3_n753 ) , .ZN( u0_u3_n844 ) );
  AOI21_X1 u0_u3_U128 (.ZN( u0_u3_n594 ) , .B2( u0_u3_n766 ) , .A( u0_u3_n788 ) , .B1( u0_u3_n815 ) );
  AOI21_X1 u0_u3_U129 (.ZN( u0_u3_n517 ) , .A( u0_u3_n782 ) , .B2( u0_u3_n795 ) , .B1( u0_u3_n815 ) );
  INV_X1 u0_u3_U13 (.A( u0_u3_n650 ) , .ZN( u0_u3_n872 ) );
  AOI21_X1 u0_u3_U130 (.B1( u0_u3_n689 ) , .ZN( u0_u3_n690 ) , .A( u0_u3_n731 ) , .B2( u0_u3_n764 ) );
  INV_X1 u0_u3_U131 (.A( u0_u3_n731 ) , .ZN( u0_u3_n854 ) );
  NOR2_X1 u0_u3_U132 (.ZN( u0_u3_n571 ) , .A1( u0_u3_n732 ) , .A2( u0_u3_n765 ) );
  INV_X1 u0_u3_U133 (.A( u0_u3_n795 ) , .ZN( u0_u3_n853 ) );
  NOR2_X1 u0_u3_U134 (.A1( u0_u3_n752 ) , .ZN( u0_u3_n770 ) , .A2( u0_u3_n806 ) );
  NOR2_X1 u0_u3_U135 (.A2( u0_u3_n438 ) , .ZN( u0_u3_n618 ) , .A1( u0_u3_n788 ) );
  AOI211_X1 u0_u3_U136 (.C2( u0_u3_n440 ) , .B( u0_u3_n626 ) , .A( u0_u3_n627 ) , .ZN( u0_u3_n638 ) , .C1( u0_u3_n865 ) );
  NOR4_X1 u0_u3_U137 (.A4( u0_u3_n632 ) , .A3( u0_u3_n633 ) , .A2( u0_u3_n634 ) , .A1( u0_u3_n635 ) , .ZN( u0_u3_n636 ) );
  NOR4_X1 u0_u3_U138 (.A4( u0_u3_n629 ) , .A3( u0_u3_n630 ) , .A2( u0_u3_n631 ) , .ZN( u0_u3_n637 ) , .A1( u0_u3_n667 ) );
  INV_X1 u0_u3_U139 (.A( u0_u3_n783 ) , .ZN( u0_u3_n852 ) );
  NOR4_X1 u0_u3_U14 (.A4( u0_u3_n547 ) , .A3( u0_u3_n548 ) , .A2( u0_u3_n549 ) , .A1( u0_u3_n550 ) , .ZN( u0_u3_n551 ) );
  OAI21_X1 u0_u3_U140 (.A( u0_u3_n701 ) , .ZN( u0_u3_n705 ) , .B2( u0_u3_n753 ) , .B1( u0_u3_n807 ) );
  OAI21_X1 u0_u3_U141 (.ZN( u0_u3_n701 ) , .B2( u0_u3_n836 ) , .B1( u0_u3_n840 ) , .A( u0_u3_n862 ) );
  INV_X1 u0_u3_U142 (.A( u0_u3_n732 ) , .ZN( u0_u3_n870 ) );
  NOR2_X1 u0_u3_U143 (.A2( u0_u3_n440 ) , .ZN( u0_u3_n628 ) , .A1( u0_u3_n841 ) );
  INV_X1 u0_u3_U144 (.A( u0_u3_n766 ) , .ZN( u0_u3_n868 ) );
  NOR2_X1 u0_u3_U145 (.ZN( u0_u3_n473 ) , .A2( u0_u3_n782 ) , .A1( u0_u3_n818 ) );
  INV_X1 u0_u3_U146 (.A( u0_u3_n440 ) , .ZN( u0_u3_n816 ) );
  INV_X1 u0_u3_U147 (.A( u0_u3_n820 ) , .ZN( u0_u3_n846 ) );
  NAND2_X1 u0_u3_U148 (.ZN( u0_u3_n717 ) , .A1( u0_u3_n731 ) , .A2( u0_u3_n783 ) );
  INV_X1 u0_u3_U149 (.A( u0_u3_n788 ) , .ZN( u0_u3_n848 ) );
  NOR4_X1 u0_u3_U15 (.A4( u0_u3_n448 ) , .A3( u0_u3_n449 ) , .A2( u0_u3_n519 ) , .A1( u0_u3_n544 ) , .ZN( u0_u3_n709 ) );
  AOI221_X1 u0_u3_U150 (.A( u0_u3_n767 ) , .ZN( u0_u3_n777 ) , .C2( u0_u3_n813 ) , .B2( u0_u3_n838 ) , .C1( u0_u3_n857 ) , .B1( u0_u3_n868 ) );
  INV_X1 u0_u3_U151 (.A( u0_u3_n764 ) , .ZN( u0_u3_n838 ) );
  AND2_X1 u0_u3_U152 (.ZN( u0_u3_n735 ) , .A1( u0_u3_n782 ) , .A2( u0_u3_n788 ) );
  AOI221_X1 u0_u3_U153 (.A( u0_u3_n453 ) , .ZN( u0_u3_n462 ) , .C2( u0_u3_n756 ) , .B1( u0_u3_n835 ) , .C1( u0_u3_n844 ) , .B2( u0_u3_n863 ) );
  AOI21_X1 u0_u3_U154 (.ZN( u0_u3_n453 ) , .B2( u0_u3_n795 ) , .A( u0_u3_n806 ) , .B1( u0_u3_n818 ) );
  AOI211_X1 u0_u3_U155 (.A( u0_u3_n591 ) , .ZN( u0_u3_n600 ) , .B( u0_u3_n624 ) , .C1( u0_u3_n847 ) , .C2( u0_u3_n857 ) );
  OAI221_X1 u0_u3_U156 (.A( u0_u3_n730 ) , .C2( u0_u3_n731 ) , .B2( u0_u3_n732 ) , .B1( u0_u3_n733 ) , .ZN( u0_u3_n740 ) , .C1( u0_u3_n820 ) );
  NAND2_X1 u0_u3_U157 (.A1( u0_u3_n444 ) , .A2( u0_u3_n467 ) , .ZN( u0_u3_n711 ) );
  NAND2_X1 u0_u3_U158 (.A2( u0_u3_n474 ) , .A1( u0_u3_n475 ) , .ZN( u0_u3_n820 ) );
  NAND2_X1 u0_u3_U159 (.A2( u0_u3_n463 ) , .A1( u0_u3_n468 ) , .ZN( u0_u3_n783 ) );
  OR3_X1 u0_u3_U16 (.ZN( u0_u3_n449 ) , .A1( u0_u3_n531 ) , .A3( u0_u3_n580 ) , .A2( u0_u3_n877 ) );
  NAND2_X1 u0_u3_U160 (.A1( u0_u3_n458 ) , .A2( u0_u3_n474 ) , .ZN( u0_u3_n806 ) );
  NAND2_X1 u0_u3_U161 (.A2( u0_u3_n451 ) , .A1( u0_u3_n463 ) , .ZN( u0_u3_n731 ) );
  NAND2_X1 u0_u3_U162 (.A1( u0_u3_n452 ) , .A2( u0_u3_n467 ) , .ZN( u0_u3_n727 ) );
  NAND2_X1 u0_u3_U163 (.A2( u0_u3_n457 ) , .A1( u0_u3_n475 ) , .ZN( u0_u3_n782 ) );
  NOR2_X1 u0_u3_U164 (.ZN( u0_u3_n456 ) , .A1( u0_u3_n829 ) , .A2( u0_u3_n830 ) );
  NAND2_X1 u0_u3_U165 (.A2( u0_u3_n467 ) , .A1( u0_u3_n468 ) , .ZN( u0_u3_n815 ) );
  NAND2_X1 u0_u3_U166 (.A2( u0_u3_n451 ) , .A1( u0_u3_n455 ) , .ZN( u0_u3_n732 ) );
  NAND2_X1 u0_u3_U167 (.A2( u0_u3_n452 ) , .A1( u0_u3_n455 ) , .ZN( u0_u3_n766 ) );
  NAND2_X1 u0_u3_U168 (.A1( u0_u3_n454 ) , .A2( u0_u3_n474 ) , .ZN( u0_u3_n819 ) );
  NAND2_X1 u0_u3_U169 (.A1( u0_u3_n456 ) , .A2( u0_u3_n464 ) , .ZN( u0_u3_n747 ) );
  OR4_X1 u0_u3_U17 (.A4( u0_u3_n445 ) , .A2( u0_u3_n446 ) , .A1( u0_u3_n447 ) , .ZN( u0_u3_n448 ) , .A3( u0_u3_n556 ) );
  NAND2_X1 u0_u3_U170 (.A2( u0_u3_n444 ) , .A1( u0_u3_n450 ) , .ZN( u0_u3_n787 ) );
  NAND2_X1 u0_u3_U171 (.A1( u0_u3_n454 ) , .A2( u0_u3_n457 ) , .ZN( u0_u3_n817 ) );
  NAND2_X1 u0_u3_U172 (.A1( u0_u3_n450 ) , .A2( u0_u3_n452 ) , .ZN( u0_u3_n808 ) );
  NAND2_X1 u0_u3_U173 (.A2( u0_u3_n456 ) , .A1( u0_u3_n458 ) , .ZN( u0_u3_n809 ) );
  NAND2_X1 u0_u3_U174 (.A1( u0_u3_n450 ) , .A2( u0_u3_n451 ) , .ZN( u0_u3_n789 ) );
  NAND2_X1 u0_u3_U175 (.A2( u0_u3_n464 ) , .A1( u0_u3_n465 ) , .ZN( u0_u3_n750 ) );
  NAND2_X1 u0_u3_U176 (.A1( u0_u3_n465 ) , .A2( u0_u3_n475 ) , .ZN( u0_u3_n791 ) );
  NAND2_X1 u0_u3_U177 (.A2( u0_u3_n457 ) , .A1( u0_u3_n458 ) , .ZN( u0_u3_n733 ) );
  NAND2_X1 u0_u3_U178 (.A1( u0_u3_n454 ) , .A2( u0_u3_n465 ) , .ZN( u0_u3_n793 ) );
  AND2_X1 u0_u3_U179 (.ZN( u0_u3_n440 ) , .A1( u0_u3_n457 ) , .A2( u0_u3_n464 ) );
  INV_X1 u0_u3_U18 (.A( u0_u3_n616 ) , .ZN( u0_u3_n877 ) );
  NOR2_X1 u0_u3_U180 (.ZN( u0_u3_n452 ) , .A1( u0_u3_n850 ) , .A2( w3_28 ) );
  NAND4_X1 u0_u3_U181 (.ZN( u0_subword_1 ) , .A4( u0_u3_n598 ) , .A3( u0_u3_n599 ) , .A2( u0_u3_n600 ) , .A1( u0_u3_n601 ) );
  AOI211_X1 u0_u3_U182 (.B( u0_u3_n592 ) , .A( u0_u3_n593 ) , .ZN( u0_u3_n599 ) , .C2( u0_u3_n814 ) , .C1( u0_u3_n836 ) );
  NOR4_X1 u0_u3_U183 (.A4( u0_u3_n594 ) , .A3( u0_u3_n595 ) , .A2( u0_u3_n596 ) , .A1( u0_u3_n597 ) , .ZN( u0_u3_n598 ) );
  NOR4_X1 u0_u3_U184 (.A4( u0_u3_n737 ) , .A3( u0_u3_n738 ) , .A2( u0_u3_n739 ) , .A1( u0_u3_n740 ) , .ZN( u0_u3_n741 ) );
  AOI211_X1 u0_u3_U185 (.B( u0_u3_n728 ) , .A( u0_u3_n729 ) , .ZN( u0_u3_n742 ) , .C1( u0_u3_n845 ) , .C2( u0_u3_n857 ) );
  AOI222_X1 u0_u3_U186 (.B2( u0_u3_n641 ) , .ZN( u0_u3_n647 ) , .B1( u0_u3_n843 ) , .A1( u0_u3_n844 ) , .C2( u0_u3_n848 ) , .C1( u0_u3_n865 ) , .A2( u0_u3_n867 ) );
  NOR4_X1 u0_u3_U187 (.A4( u0_u3_n642 ) , .A3( u0_u3_n643 ) , .A2( u0_u3_n644 ) , .A1( u0_u3_n645 ) , .ZN( u0_u3_n646 ) );
  AOI221_X1 u0_u3_U188 (.A( u0_u3_n784 ) , .ZN( u0_u3_n801 ) , .C2( u0_u3_n839 ) , .B2( u0_u3_n840 ) , .B1( u0_u3_n867 ) , .C1( u0_u3_n868 ) );
  NOR4_X1 u0_u3_U189 (.A4( u0_u3_n796 ) , .A3( u0_u3_n797 ) , .A2( u0_u3_n798 ) , .A1( u0_u3_n799 ) , .ZN( u0_u3_n800 ) );
  NOR4_X1 u0_u3_U19 (.ZN( u0_u3_n478 ) , .A1( u0_u3_n534 ) , .A3( u0_u3_n571 ) , .A4( u0_u3_n603 ) , .A2( u0_u3_n645 ) );
  NAND4_X1 u0_u3_U190 (.ZN( u0_subword_0 ) , .A4( u0_u3_n504 ) , .A3( u0_u3_n505 ) , .A2( u0_u3_n506 ) , .A1( u0_u3_n507 ) );
  NOR4_X1 u0_u3_U191 (.A4( u0_u3_n501 ) , .A3( u0_u3_n502 ) , .A2( u0_u3_n503 ) , .ZN( u0_u3_n504 ) , .A1( u0_u3_n530 ) );
  AOI221_X1 u0_u3_U192 (.A( u0_u3_n500 ) , .ZN( u0_u3_n505 ) , .B2( u0_u3_n845 ) , .C1( u0_u3_n848 ) , .C2( u0_u3_n862 ) , .B1( u0_u3_n864 ) );
  NOR4_X1 u0_u3_U193 (.A4( u0_u3_n703 ) , .A3( u0_u3_n704 ) , .A2( u0_u3_n705 ) , .A1( u0_u3_n706 ) , .ZN( u0_u3_n707 ) );
  NOR4_X1 u0_u3_U194 (.A3( u0_u3_n758 ) , .A2( u0_u3_n759 ) , .A1( u0_u3_n760 ) , .ZN( u0_u3_n761 ) , .A4( u0_u3_n871 ) );
  AOI211_X1 u0_u3_U195 (.B( u0_u3_n748 ) , .A( u0_u3_n749 ) , .ZN( u0_u3_n762 ) , .C1( u0_u3_n835 ) , .C2( u0_u3_n855 ) );
  NAND4_X1 u0_u3_U196 (.ZN( u0_subword_7 ) , .A4( u0_u3_n825 ) , .A3( u0_u3_n826 ) , .A2( u0_u3_n827 ) , .A1( u0_u3_n828 ) );
  NOR4_X1 u0_u3_U197 (.A4( u0_u3_n821 ) , .A3( u0_u3_n822 ) , .A2( u0_u3_n823 ) , .A1( u0_u3_n824 ) , .ZN( u0_u3_n825 ) );
  NAND2_X1 u0_u3_U198 (.A2( u0_u3_n464 ) , .A1( u0_u3_n474 ) , .ZN( u0_u3_n700 ) );
  NAND2_X1 u0_u3_U199 (.A2( u0_u3_n451 ) , .A1( u0_u3_n467 ) , .ZN( u0_u3_n818 ) );
  INV_X1 u0_u3_U20 (.A( u0_u3_n752 ) , .ZN( u0_u3_n865 ) );
  OAI21_X1 u0_u3_U200 (.B1( u0_u3_n756 ) , .ZN( u0_u3_n757 ) , .A( u0_u3_n847 ) , .B2( u0_u3_n870 ) );
  AOI221_X1 u0_u3_U201 (.A( u0_u3_n567 ) , .C2( u0_u3_n568 ) , .ZN( u0_u3_n577 ) , .B2( u0_u3_n847 ) , .B1( u0_u3_n854 ) , .C1( u0_u3_n855 ) );
  AOI222_X1 u0_u3_U202 (.ZN( u0_u3_n663 ) , .A2( u0_u3_n841 ) , .B1( u0_u3_n843 ) , .C2( u0_u3_n847 ) , .A1( u0_u3_n862 ) , .C1( u0_u3_n865 ) , .B2( u0_u3_n872 ) );
  AOI221_X1 u0_u3_U203 (.A( u0_u3_n713 ) , .ZN( u0_u3_n724 ) , .C2( u0_u3_n846 ) , .B2( u0_u3_n847 ) , .C1( u0_u3_n863 ) , .B1( u0_u3_n864 ) );
  NAND4_X1 u0_u3_U204 (.A4( u0_u3_n538 ) , .A3( u0_u3_n539 ) , .A2( u0_u3_n540 ) , .A1( u0_u3_n541 ) , .ZN( u0_u3_n625 ) );
  NOR4_X1 u0_u3_U205 (.A1( u0_u3_n534 ) , .ZN( u0_u3_n539 ) , .A2( u0_u3_n657 ) , .A4( u0_u3_n671 ) , .A3( u0_u3_n768 ) );
  NAND4_X1 u0_u3_U206 (.A4( u0_u3_n496 ) , .A3( u0_u3_n497 ) , .A1( u0_u3_n498 ) , .ZN( u0_u3_n805 ) , .A2( u0_u3_n869 ) );
  NOR4_X1 u0_u3_U207 (.A2( u0_u3_n494 ) , .A1( u0_u3_n495 ) , .ZN( u0_u3_n496 ) , .A3( u0_u3_n583 ) , .A4( u0_u3_n615 ) );
  NAND2_X1 u0_u3_U208 (.A1( u0_u3_n444 ) , .A2( u0_u3_n463 ) , .ZN( u0_u3_n702 ) );
  NAND2_X1 u0_u3_U209 (.A1( u0_u3_n455 ) , .A2( u0_u3_n468 ) , .ZN( u0_u3_n672 ) );
  AOI222_X1 u0_u3_U21 (.ZN( u0_u3_n566 ) , .B1( u0_u3_n833 ) , .C1( u0_u3_n843 ) , .A2( u0_u3_n845 ) , .A1( u0_u3_n856 ) , .B2( u0_u3_n865 ) , .C2( u0_u3_n875 ) );
  NAND4_X1 u0_u3_U210 (.A4( u0_u3_n563 ) , .A3( u0_u3_n564 ) , .A2( u0_u3_n565 ) , .A1( u0_u3_n566 ) , .ZN( u0_u3_n610 ) );
  NOR4_X1 u0_u3_U211 (.ZN( u0_u3_n564 ) , .A1( u0_u3_n656 ) , .A3( u0_u3_n664 ) , .A4( u0_u3_n688 ) , .A2( u0_u3_n771 ) );
  NOR2_X1 u0_u3_U212 (.ZN( u0_u3_n454 ) , .A1( u0_u3_n831 ) , .A2( u0_u3_n832 ) );
  INV_X1 u0_u3_U213 (.ZN( u0_u3_n831 ) , .A( w3_26 ) );
  NOR2_X1 u0_u3_U214 (.ZN( u0_u3_n710 ) , .A2( u0_u3_n779 ) , .A1( u0_u3_n803 ) );
  OAI21_X1 u0_u3_U215 (.A( u0_u3_n734 ) , .B1( u0_u3_n735 ) , .ZN( u0_u3_n739 ) , .B2( u0_u3_n808 ) );
  AOI21_X1 u0_u3_U216 (.ZN( u0_u3_n653 ) , .A( u0_u3_n782 ) , .B1( u0_u3_n795 ) , .B2( u0_u3_n808 ) );
  INV_X1 u0_u3_U217 (.A( u0_u3_n808 ) , .ZN( u0_u3_n862 ) );
  NOR2_X1 u0_u3_U218 (.ZN( u0_u3_n738 ) , .A2( u0_u3_n806 ) , .A1( u0_u3_n808 ) );
  NAND2_X1 u0_u3_U219 (.ZN( u0_u3_n756 ) , .A1( u0_u3_n766 ) , .A2( u0_u3_n808 ) );
  NOR4_X1 u0_u3_U22 (.ZN( u0_u3_n482 ) , .A1( u0_u3_n523 ) , .A4( u0_u3_n560 ) , .A3( u0_u3_n585 ) , .A2( u0_u3_n633 ) );
  NOR2_X1 u0_u3_U220 (.ZN( u0_u3_n559 ) , .A1( u0_u3_n765 ) , .A2( u0_u3_n808 ) );
  OAI221_X1 u0_u3_U221 (.A( u0_u3_n699 ) , .ZN( u0_u3_n706 ) , .C2( u0_u3_n787 ) , .C1( u0_u3_n788 ) , .B1( u0_u3_n789 ) , .B2( u0_u3_n809 ) );
  OAI222_X1 u0_u3_U222 (.B1( u0_u3_n41 ) , .ZN( u0_u3_n620 ) , .C1( u0_u3_n727 ) , .C2( u0_u3_n750 ) , .B2( u0_u3_n789 ) , .A2( u0_u3_n795 ) , .A1( u0_u3_n819 ) );
  NAND2_X1 u0_u3_U223 (.A2( u0_u3_n444 ) , .A1( u0_u3_n455 ) , .ZN( u0_u3_n794 ) );
  OAI222_X1 u0_u3_U224 (.B2( u0_u3_n711 ) , .ZN( u0_u3_n712 ) , .C2( u0_u3_n727 ) , .B1( u0_u3_n750 ) , .A1( u0_u3_n809 ) , .C1( u0_u3_n817 ) , .A2( u0_u3_n818 ) );
  INV_X1 u0_u3_U225 (.A( u0_u3_n675 ) , .ZN( u0_u3_n861 ) );
  NOR2_X1 u0_u3_U226 (.ZN( u0_u3_n531 ) , .A2( u0_u3_n727 ) , .A1( u0_u3_n806 ) );
  NOR2_X1 u0_u3_U227 (.ZN( u0_u3_n529 ) , .A1( u0_u3_n727 ) , .A2( u0_u3_n753 ) );
  INV_X1 u0_u3_U228 (.A( u0_u3_n727 ) , .ZN( u0_u3_n858 ) );
  NOR2_X1 u0_u3_U229 (.ZN( u0_u3_n450 ) , .A2( u0_u3_n851 ) , .A1( u0_u3_n860 ) );
  NOR4_X1 u0_u3_U23 (.A4( u0_u3_n559 ) , .A3( u0_u3_n560 ) , .A2( u0_u3_n561 ) , .A1( u0_u3_n562 ) , .ZN( u0_u3_n563 ) );
  AOI222_X1 u0_u3_U230 (.ZN( u0_u3_n528 ) , .A1( u0_u3_n837 ) , .B2( u0_u3_n839 ) , .C1( u0_u3_n846 ) , .C2( u0_u3_n852 ) , .A2( u0_u3_n854 ) , .B1( u0_u3_n868 ) );
  NOR3_X1 u0_u3_U231 (.A2( u0_u3_n440 ) , .ZN( u0_u3_n443 ) , .A3( u0_u3_n839 ) , .A1( u0_u3_n848 ) );
  NAND2_X1 u0_u3_U232 (.ZN( u0_u3_n616 ) , .A2( u0_u3_n839 ) , .A1( u0_u3_n875 ) );
  NOR2_X1 u0_u3_U233 (.ZN( u0_u3_n498 ) , .A1( u0_u3_n681 ) , .A2( u0_u3_n697 ) );
  AOI211_X1 u0_u3_U234 (.B( u0_u3_n697 ) , .A( u0_u3_n698 ) , .ZN( u0_u3_n708 ) , .C2( u0_u3_n834 ) , .C1( u0_u3_n853 ) );
  NOR2_X1 u0_u3_U235 (.ZN( u0_u3_n586 ) , .A1( u0_u3_n795 ) , .A2( u0_u3_n820 ) );
  AOI21_X1 u0_u3_U236 (.ZN( u0_u3_n543 ) , .A( u0_u3_n766 ) , .B2( u0_u3_n782 ) , .B1( u0_u3_n820 ) );
  NOR2_X1 u0_u3_U237 (.ZN( u0_u3_n612 ) , .A2( u0_u3_n727 ) , .A1( u0_u3_n820 ) );
  NOR2_X1 u0_u3_U238 (.ZN( u0_u3_n718 ) , .A1( u0_u3_n808 ) , .A2( u0_u3_n820 ) );
  OAI21_X1 u0_u3_U239 (.A( u0_u3_n790 ) , .B2( u0_u3_n791 ) , .B1( u0_u3_n792 ) , .ZN( u0_u3_n798 ) );
  NOR4_X1 u0_u3_U24 (.A4( u0_u3_n555 ) , .A3( u0_u3_n556 ) , .A2( u0_u3_n557 ) , .A1( u0_u3_n558 ) , .ZN( u0_u3_n565 ) );
  AOI21_X1 u0_u3_U240 (.ZN( u0_u3_n642 ) , .B2( u0_u3_n752 ) , .A( u0_u3_n791 ) , .B1( u0_u3_n815 ) );
  AOI21_X1 u0_u3_U241 (.A( u0_u3_n736 ) , .ZN( u0_u3_n737 ) , .B2( u0_u3_n783 ) , .B1( u0_u3_n795 ) );
  AOI21_X1 u0_u3_U242 (.B2( u0_u3_n766 ) , .ZN( u0_u3_n767 ) , .A( u0_u3_n791 ) , .B1( u0_u3_n795 ) );
  NOR2_X1 u0_u3_U243 (.ZN( u0_u3_n521 ) , .A1( u0_u3_n711 ) , .A2( u0_u3_n791 ) );
  NOR2_X1 u0_u3_U244 (.ZN( u0_u3_n487 ) , .A1( u0_u3_n791 ) , .A2( u0_u3_n808 ) );
  NOR2_X1 u0_u3_U245 (.ZN( u0_u3_n537 ) , .A1( u0_u3_n727 ) , .A2( u0_u3_n791 ) );
  INV_X1 u0_u3_U246 (.A( u0_u3_n791 ) , .ZN( u0_u3_n847 ) );
  OAI22_X1 u0_u3_U247 (.B2( u0_u3_n782 ) , .B1( u0_u3_n783 ) , .ZN( u0_u3_n784 ) , .A2( u0_u3_n817 ) , .A1( u0_u3_n818 ) );
  AOI21_X1 u0_u3_U248 (.ZN( u0_u3_n501 ) , .A( u0_u3_n727 ) , .B2( u0_u3_n765 ) , .B1( u0_u3_n817 ) );
  NAND4_X1 u0_u3_U249 (.A4( u0_u3_n482 ) , .A3( u0_u3_n483 ) , .A2( u0_u3_n484 ) , .A1( u0_u3_n485 ) , .ZN( u0_u3_n697 ) );
  NOR4_X1 u0_u3_U25 (.A4( u0_u3_n771 ) , .A3( u0_u3_n772 ) , .A2( u0_u3_n773 ) , .A1( u0_u3_n774 ) , .ZN( u0_u3_n775 ) );
  AOI21_X1 u0_u3_U250 (.ZN( u0_u3_n542 ) , .B2( u0_u3_n815 ) , .A( u0_u3_n817 ) , .B1( u0_u3_n818 ) );
  NOR2_X1 u0_u3_U251 (.ZN( u0_u3_n523 ) , .A2( u0_u3_n711 ) , .A1( u0_u3_n817 ) );
  NOR2_X1 u0_u3_U252 (.ZN( u0_u3_n549 ) , .A2( u0_u3_n783 ) , .A1( u0_u3_n817 ) );
  INV_X1 u0_u3_U253 (.A( u0_u3_n817 ) , .ZN( u0_u3_n836 ) );
  NOR2_X1 u0_u3_U254 (.ZN( u0_u3_n548 ) , .A1( u0_u3_n752 ) , .A2( u0_u3_n817 ) );
  NOR2_X1 u0_u3_U255 (.ZN( u0_u3_n560 ) , .A1( u0_u3_n795 ) , .A2( u0_u3_n817 ) );
  AOI21_X1 u0_u3_U256 (.A( u0_u3_n673 ) , .B1( u0_u3_n674 ) , .ZN( u0_u3_n675 ) , .B2( u0_u3_n858 ) );
  AOI22_X1 u0_u3_U257 (.A2( u0_u3_n785 ) , .ZN( u0_u3_n786 ) , .B2( u0_u3_n834 ) , .A1( u0_u3_n837 ) , .B1( u0_u3_n865 ) );
  AOI21_X1 u0_u3_U258 (.ZN( u0_u3_n643 ) , .B2( u0_u3_n750 ) , .A( u0_u3_n795 ) , .B1( u0_u3_n806 ) );
  NAND4_X1 u0_u3_U259 (.A4( u0_u3_n775 ) , .A3( u0_u3_n776 ) , .A2( u0_u3_n777 ) , .A1( u0_u3_n778 ) , .ZN( u0_u3_n804 ) );
  NOR3_X1 u0_u3_U26 (.A3( u0_u3_n768 ) , .A2( u0_u3_n769 ) , .A1( u0_u3_n770 ) , .ZN( u0_u3_n776 ) );
  OAI21_X1 u0_u3_U260 (.ZN( u0_u3_n466 ) , .B1( u0_u3_n812 ) , .A( u0_u3_n837 ) , .B2( u0_u3_n853 ) );
  NOR2_X1 u0_u3_U261 (.ZN( u0_u3_n659 ) , .A1( u0_u3_n750 ) , .A2( u0_u3_n783 ) );
  NOR2_X1 u0_u3_U262 (.ZN( u0_u3_n683 ) , .A2( u0_u3_n837 ) , .A1( u0_u3_n841 ) );
  NOR2_X1 u0_u3_U263 (.ZN( u0_u3_n764 ) , .A1( u0_u3_n836 ) , .A2( u0_u3_n837 ) );
  NOR2_X1 u0_u3_U264 (.ZN( u0_u3_n570 ) , .A1( u0_u3_n750 ) , .A2( u0_u3_n808 ) );
  NOR2_X1 u0_u3_U265 (.A2( u0_u3_n438 ) , .ZN( u0_u3_n633 ) , .A1( u0_u3_n750 ) );
  INV_X1 u0_u3_U266 (.A( u0_u3_n750 ) , .ZN( u0_u3_n837 ) );
  NOR4_X1 u0_u3_U267 (.ZN( u0_u3_n488 ) , .A2( u0_u3_n536 ) , .A1( u0_u3_n561 ) , .A3( u0_u3_n634 ) , .A4( u0_u3_n721 ) );
  NAND4_X1 u0_u3_U268 (.A4( u0_u3_n488 ) , .A3( u0_u3_n489 ) , .A2( u0_u3_n490 ) , .A1( u0_u3_n491 ) , .ZN( u0_u3_n781 ) );
  AOI21_X1 u0_u3_U269 (.B1( u0_u3_n438 ) , .ZN( u0_u3_n592 ) , .B2( u0_u3_n702 ) , .A( u0_u3_n820 ) );
  NAND4_X1 u0_u3_U27 (.A4( u0_u3_n606 ) , .A3( u0_u3_n607 ) , .A2( u0_u3_n608 ) , .A1( u0_u3_n609 ) , .ZN( u0_u3_n725 ) );
  AOI21_X1 u0_u3_U270 (.B1( u0_u3_n702 ) , .ZN( u0_u3_n703 ) , .A( u0_u3_n735 ) , .B2( u0_u3_n766 ) );
  INV_X1 u0_u3_U271 (.A( u0_u3_n702 ) , .ZN( u0_u3_n855 ) );
  AOI21_X1 u0_u3_U272 (.ZN( u0_u3_n445 ) , .A( u0_u3_n702 ) , .B1( u0_u3_n736 ) , .B2( u0_u3_n753 ) );
  NOR2_X1 u0_u3_U273 (.ZN( u0_u3_n686 ) , .A2( u0_u3_n702 ) , .A1( u0_u3_n806 ) );
  NOR2_X1 u0_u3_U274 (.ZN( u0_u3_n580 ) , .A2( u0_u3_n702 ) , .A1( u0_u3_n817 ) );
  NAND2_X1 u0_u3_U275 (.A1( u0_u3_n702 ) , .A2( u0_u3_n732 ) , .ZN( u0_u3_n785 ) );
  NOR3_X1 u0_u3_U276 (.A3( u0_u3_n744 ) , .A2( u0_u3_n745 ) , .A1( u0_u3_n746 ) , .ZN( u0_u3_n763 ) );
  OAI22_X1 u0_u3_U277 (.ZN( u0_u3_n492 ) , .A1( u0_u3_n727 ) , .B2( u0_u3_n731 ) , .B1( u0_u3_n733 ) , .A2( u0_u3_n782 ) );
  NOR2_X1 u0_u3_U278 (.ZN( u0_u3_n582 ) , .A2( u0_u3_n711 ) , .A1( u0_u3_n733 ) );
  NOR2_X1 u0_u3_U279 (.ZN( u0_u3_n536 ) , .A2( u0_u3_n727 ) , .A1( u0_u3_n733 ) );
  NOR3_X1 u0_u3_U28 (.A1( u0_u3_n602 ) , .ZN( u0_u3_n607 ) , .A3( u0_u3_n666 ) , .A2( u0_u3_n773 ) );
  AOI222_X1 u0_u3_U280 (.ZN( u0_u3_n608 ) , .B2( u0_u3_n674 ) , .B1( u0_u3_n756 ) , .C2( u0_u3_n834 ) , .A1( u0_u3_n836 ) , .A2( u0_u3_n864 ) , .C1( u0_u3_n865 ) );
  AOI221_X1 u0_u3_U281 (.A( u0_u3_n486 ) , .ZN( u0_u3_n491 ) , .B1( u0_u3_n834 ) , .C2( u0_u3_n846 ) , .C1( u0_u3_n854 ) , .B2( u0_u3_n864 ) );
  NOR2_X1 u0_u3_U282 (.ZN( u0_u3_n792 ) , .A2( u0_u3_n864 ) , .A1( u0_u3_n870 ) );
  NOR2_X1 u0_u3_U283 (.ZN( u0_u3_n464 ) , .A1( u0_u3_n832 ) , .A2( w3_26 ) );
  NOR2_X1 u0_u3_U284 (.ZN( u0_u3_n474 ) , .A1( u0_u3_n829 ) , .A2( w3_25 ) );
  AOI21_X1 u0_u3_U285 (.A( u0_u3_n439 ) , .ZN( u0_u3_n644 ) , .B1( u0_u3_n683 ) , .B2( u0_u3_n820 ) );
  AOI21_X1 u0_u3_U286 (.B2( u0_u3_n439 ) , .ZN( u0_u3_n500 ) , .A( u0_u3_n782 ) , .B1( u0_u3_n807 ) );
  OAI22_X1 u0_u3_U287 (.B1( u0_u3_n439 ) , .ZN( u0_u3_n698 ) , .A2( u0_u3_n733 ) , .A1( u0_u3_n783 ) , .B2( u0_u3_n820 ) );
  AOI21_X1 u0_u3_U288 (.B2( u0_u3_n439 ) , .ZN( u0_u3_n567 ) , .B1( u0_u3_n727 ) , .A( u0_u3_n782 ) );
  AOI21_X1 u0_u3_U289 (.B2( u0_u3_n439 ) , .ZN( u0_u3_n446 ) , .B1( u0_u3_n792 ) , .A( u0_u3_n817 ) );
  NOR4_X1 u0_u3_U29 (.A3( u0_u3_n603 ) , .A2( u0_u3_n604 ) , .A1( u0_u3_n605 ) , .ZN( u0_u3_n606 ) , .A4( u0_u3_n658 ) );
  NOR2_X1 u0_u3_U290 (.A2( u0_u3_n439 ) , .ZN( u0_u3_n667 ) , .A1( u0_u3_n788 ) );
  NOR2_X1 u0_u3_U291 (.A2( u0_u3_n439 ) , .ZN( u0_u3_n558 ) , .A1( u0_u3_n753 ) );
  NOR2_X1 u0_u3_U292 (.A2( u0_u3_n439 ) , .ZN( u0_u3_n562 ) , .A1( u0_u3_n806 ) );
  NOR2_X1 u0_u3_U293 (.A1( u0_u3_n439 ) , .ZN( u0_u3_n645 ) , .A2( u0_u3_n791 ) );
  NOR2_X1 u0_u3_U294 (.A2( u0_u3_n439 ) , .ZN( u0_u3_n545 ) , .A1( u0_u3_n765 ) );
  INV_X1 u0_u3_U295 (.A( u0_u3_n794 ) , .ZN( u0_u3_n875 ) );
  NOR2_X1 u0_u3_U296 (.ZN( u0_u3_n463 ) , .A1( u0_u3_n851 ) , .A2( w3_31 ) );
  AOI21_X1 u0_u3_U297 (.B2( u0_u3_n439 ) , .A( u0_u3_n793 ) , .B1( u0_u3_n795 ) , .ZN( u0_u3_n796 ) );
  AOI222_X1 u0_u3_U298 (.C2( u0_u3_n812 ) , .B2( u0_u3_n813 ) , .A2( u0_u3_n814 ) , .ZN( u0_u3_n826 ) , .C1( u0_u3_n835 ) , .A1( u0_u3_n841 ) , .B1( u0_u3_n855 ) );
  AOI22_X1 u0_u3_U299 (.ZN( u0_u3_n730 ) , .B1( u0_u3_n835 ) , .A2( u0_u3_n840 ) , .A1( u0_u3_n865 ) , .B2( u0_u3_n868 ) );
  BUF_X1 u0_u3_U3 (.Z( u0_u3_n438 ) , .A( u0_u3_n818 ) );
  NOR4_X1 u0_u3_U30 (.A4( u0_u3_n487 ) , .ZN( u0_u3_n490 ) , .A1( u0_u3_n569 ) , .A2( u0_u3_n584 ) , .A3( u0_u3_n605 ) );
  AOI222_X1 u0_u3_U300 (.ZN( u0_u3_n516 ) , .C1( u0_u3_n835 ) , .B2( u0_u3_n839 ) , .A2( u0_u3_n845 ) , .C2( u0_u3_n864 ) , .B1( u0_u3_n865 ) , .A1( u0_u3_n868 ) );
  AOI222_X1 u0_u3_U301 (.ZN( u0_u3_n472 ) , .B1( u0_u3_n835 ) , .A1( u0_u3_n841 ) , .C1( u0_u3_n844 ) , .C2( u0_u3_n853 ) , .A2( u0_u3_n857 ) , .B2( u0_u3_n867 ) );
  NOR2_X1 u0_u3_U302 (.A2( u0_u3_n438 ) , .ZN( u0_u3_n658 ) , .A1( u0_u3_n793 ) );
  NOR2_X1 u0_u3_U303 (.ZN( u0_u3_n715 ) , .A2( u0_u3_n727 ) , .A1( u0_u3_n793 ) );
  NOR2_X1 u0_u3_U304 (.ZN( u0_u3_n689 ) , .A1( u0_u3_n834 ) , .A2( u0_u3_n835 ) );
  NOR2_X1 u0_u3_U305 (.ZN( u0_u3_n524 ) , .A1( u0_u3_n793 ) , .A2( u0_u3_n815 ) );
  NOR2_X1 u0_u3_U306 (.ZN( u0_u3_n664 ) , .A1( u0_u3_n732 ) , .A2( u0_u3_n793 ) );
  NOR2_X1 u0_u3_U307 (.ZN( u0_u3_n736 ) , .A2( u0_u3_n835 ) , .A1( u0_u3_n847 ) );
  NOR2_X1 u0_u3_U308 (.ZN( u0_u3_n671 ) , .A2( u0_u3_n711 ) , .A1( u0_u3_n793 ) );
  NOR2_X1 u0_u3_U309 (.ZN( u0_u3_n673 ) , .A1( u0_u3_n793 ) , .A2( u0_u3_n808 ) );
  NOR4_X1 u0_u3_U31 (.ZN( u0_u3_n489 ) , .A1( u0_u3_n510 ) , .A2( u0_u3_n522 ) , .A4( u0_u3_n549 ) , .A3( u0_u3_n614 ) );
  INV_X1 u0_u3_U310 (.A( u0_u3_n793 ) , .ZN( u0_u3_n835 ) );
  AOI21_X1 u0_u3_U311 (.B1( u0_u3_n438 ) , .ZN( u0_u3_n513 ) , .B2( u0_u3_n672 ) , .A( u0_u3_n733 ) );
  AOI21_X1 u0_u3_U312 (.B1( u0_u3_n439 ) , .ZN( u0_u3_n629 ) , .B2( u0_u3_n672 ) , .A( u0_u3_n793 ) );
  INV_X1 u0_u3_U313 (.A( u0_u3_n672 ) , .ZN( u0_u3_n867 ) );
  NOR2_X1 u0_u3_U314 (.ZN( u0_u3_n655 ) , .A1( u0_u3_n672 ) , .A2( u0_u3_n817 ) );
  NOR2_X1 u0_u3_U315 (.ZN( u0_u3_n631 ) , .A2( u0_u3_n672 ) , .A1( u0_u3_n788 ) );
  NOR2_X1 u0_u3_U316 (.ZN( u0_u3_n605 ) , .A1( u0_u3_n672 ) , .A2( u0_u3_n806 ) );
  NOR2_X1 u0_u3_U317 (.ZN( u0_u3_n530 ) , .A1( u0_u3_n672 ) , .A2( u0_u3_n782 ) );
  NOR2_X1 u0_u3_U318 (.ZN( u0_u3_n584 ) , .A1( u0_u3_n672 ) , .A2( u0_u3_n791 ) );
  NOR2_X1 u0_u3_U319 (.ZN( u0_u3_n444 ) , .A2( w3_28 ) , .A1( w3_29 ) );
  NOR4_X1 u0_u3_U32 (.A4( u0_u3_n529 ) , .A2( u0_u3_n530 ) , .A1( u0_u3_n531 ) , .ZN( u0_u3_n541 ) , .A3( u0_u3_n704 ) );
  NOR2_X1 u0_u3_U320 (.ZN( u0_u3_n468 ) , .A2( u0_u3_n849 ) , .A1( u0_u3_n850 ) );
  OAI222_X1 u0_u3_U321 (.B2( u0_u3_n750 ) , .B1( u0_u3_n751 ) , .A2( u0_u3_n752 ) , .ZN( u0_u3_n760 ) , .C2( u0_u3_n808 ) , .C1( u0_u3_n817 ) , .A1( u0_u3_n820 ) );
  INV_X1 u0_u3_U322 (.A( u0_u3_n789 ) , .ZN( u0_u3_n864 ) );
  NOR4_X1 u0_u3_U323 (.A4( u0_u3_n617 ) , .A3( u0_u3_n618 ) , .A1( u0_u3_n619 ) , .A2( u0_u3_n620 ) , .ZN( u0_u3_n621 ) );
  INV_X1 u0_u3_U324 (.ZN( u0_u3_n830 ) , .A( w3_25 ) );
  OAI22_X1 u0_u3_U325 (.B2( u0_u3_n753 ) , .B1( u0_u3_n754 ) , .A1( u0_u3_n755 ) , .ZN( u0_u3_n759 ) , .A2( u0_u3_n809 ) );
  OAI22_X1 u0_u3_U326 (.B2( u0_u3_n806 ) , .B1( u0_u3_n807 ) , .A2( u0_u3_n808 ) , .A1( u0_u3_n809 ) , .ZN( u0_u3_n811 ) );
  AOI21_X1 u0_u3_U327 (.ZN( u0_u3_n692 ) , .B2( u0_u3_n752 ) , .B1( u0_u3_n766 ) , .A( u0_u3_n809 ) );
  NAND2_X1 u0_u3_U328 (.A2( u0_u3_n765 ) , .A1( u0_u3_n809 ) , .ZN( u0_u3_n813 ) );
  NOR2_X1 u0_u3_U329 (.ZN( u0_u3_n573 ) , .A1( u0_u3_n731 ) , .A2( u0_u3_n809 ) );
  NOR4_X1 u0_u3_U33 (.A4( u0_u3_n535 ) , .A3( u0_u3_n536 ) , .A2( u0_u3_n537 ) , .ZN( u0_u3_n538 ) , .A1( u0_u3_n823 ) );
  NOR2_X1 u0_u3_U330 (.ZN( u0_u3_n614 ) , .A2( u0_u3_n783 ) , .A1( u0_u3_n809 ) );
  OAI22_X1 u0_u3_U331 (.ZN( u0_u3_n486 ) , .A1( u0_u3_n711 ) , .B2( u0_u3_n788 ) , .A2( u0_u3_n809 ) , .B1( u0_u3_n815 ) );
  AOI21_X1 u0_u3_U332 (.ZN( u0_u3_n480 ) , .A( u0_u3_n672 ) , .B1( u0_u3_n753 ) , .B2( u0_u3_n809 ) );
  INV_X1 u0_u3_U333 (.A( u0_u3_n809 ) , .ZN( u0_u3_n843 ) );
  OAI221_X1 u0_u3_U334 (.A( u0_u3_n786 ) , .C2( u0_u3_n787 ) , .B2( u0_u3_n788 ) , .B1( u0_u3_n789 ) , .ZN( u0_u3_n799 ) , .C1( u0_u3_n816 ) );
  NAND2_X1 u0_u3_U335 (.A1( u0_u3_n732 ) , .A2( u0_u3_n787 ) , .ZN( u0_u3_n814 ) );
  OAI22_X1 u0_u3_U336 (.ZN( u0_u3_n591 ) , .A2( u0_u3_n750 ) , .B2( u0_u3_n765 ) , .A1( u0_u3_n766 ) , .B1( u0_u3_n787 ) );
  AOI21_X1 u0_u3_U337 (.ZN( u0_u3_n595 ) , .B1( u0_u3_n731 ) , .B2( u0_u3_n787 ) , .A( u0_u3_n793 ) );
  NOR2_X1 u0_u3_U338 (.ZN( u0_u3_n807 ) , .A1( u0_u3_n856 ) , .A2( u0_u3_n863 ) );
  AOI21_X1 u0_u3_U339 (.ZN( u0_u3_n626 ) , .B1( u0_u3_n702 ) , .A( u0_u3_n782 ) , .B2( u0_u3_n787 ) );
  NOR4_X1 u0_u3_U34 (.A4( u0_u3_n532 ) , .A3( u0_u3_n533 ) , .ZN( u0_u3_n540 ) , .A2( u0_u3_n687 ) , .A1( u0_u3_n797 ) );
  NAND2_X2 u0_u3_U340 (.A1( u0_u3_n458 ) , .A2( u0_u3_n465 ) , .ZN( u0_u3_n753 ) );
  AOI222_X1 u0_u3_U341 (.ZN( u0_u3_n778 ) , .A1( u0_u3_n833 ) , .C1( u0_u3_n837 ) , .B2( u0_u3_n843 ) , .A2( u0_u3_n852 ) , .B1( u0_u3_n863 ) , .C2( u0_u3_n875 ) );
  AOI222_X1 u0_u3_U342 (.ZN( u0_u3_n609 ) , .A1( u0_u3_n833 ) , .C2( u0_u3_n839 ) , .B1( u0_u3_n844 ) , .A2( u0_u3_n858 ) , .B2( u0_u3_n863 ) , .C1( u0_u3_n870 ) );
  AOI21_X1 u0_u3_U343 (.ZN( u0_u3_n651 ) , .A( u0_u3_n765 ) , .B2( u0_u3_n787 ) , .B1( u0_u3_n795 ) );
  OAI22_X1 u0_u3_U344 (.ZN( u0_u3_n684 ) , .A1( u0_u3_n702 ) , .A2( u0_u3_n733 ) , .B2( u0_u3_n787 ) , .B1( u0_u3_n820 ) );
  NOR2_X1 u0_u3_U345 (.ZN( u0_u3_n654 ) , .A1( u0_u3_n787 ) , .A2( u0_u3_n791 ) );
  NOR2_X1 u0_u3_U346 (.ZN( u0_u3_n751 ) , .A1( u0_u3_n863 ) , .A2( u0_u3_n864 ) );
  NOR2_X1 u0_u3_U347 (.ZN( u0_u3_n455 ) , .A1( u0_u3_n860 ) , .A2( w3_30 ) );
  NOR2_X1 u0_u3_U348 (.ZN( u0_u3_n467 ) , .A2( w3_30 ) , .A1( w3_31 ) );
  AND2_X1 u0_u3_U349 (.ZN( u0_u3_n441 ) , .A2( u0_u3_n834 ) , .A1( u0_u3_n856 ) );
  NOR3_X1 u0_u3_U35 (.A3( u0_u3_n803 ) , .A2( u0_u3_n804 ) , .A1( u0_u3_n805 ) , .ZN( u0_u3_n828 ) );
  AND2_X1 u0_u3_U350 (.ZN( u0_u3_n442 ) , .A2( u0_u3_n845 ) , .A1( u0_u3_n863 ) );
  NOR3_X1 u0_u3_U351 (.A3( u0_u3_n441 ) , .A2( u0_u3_n442 ) , .A1( u0_u3_n579 ) , .ZN( u0_u3_n590 ) );
  INV_X1 u0_u3_U352 (.A( u0_u3_n815 ) , .ZN( u0_u3_n856 ) );
  INV_X1 u0_u3_U353 (.A( u0_u3_n787 ) , .ZN( u0_u3_n863 ) );
  INV_X1 u0_u3_U354 (.A( u0_u3_n806 ) , .ZN( u0_u3_n845 ) );
  INV_X1 u0_u3_U355 (.A( u0_u3_n41 ) , .ZN( u0_u3_n840 ) );
  NOR2_X1 u0_u3_U356 (.A1( u0_u3_n41 ) , .ZN( u0_u3_n773 ) , .A2( u0_u3_n818 ) );
  AOI21_X1 u0_u3_U357 (.B2( u0_u3_n41 ) , .ZN( u0_u3_n574 ) , .B1( u0_u3_n809 ) , .A( u0_u3_n815 ) );
  NOR2_X1 u0_u3_U358 (.A2( u0_u3_n41 ) , .ZN( u0_u3_n665 ) , .A1( u0_u3_n732 ) );
  NOR2_X1 u0_u3_U359 (.A2( u0_u3_n41 ) , .ZN( u0_u3_n635 ) , .A1( u0_u3_n727 ) );
  NAND4_X1 u0_u3_U36 (.A4( u0_u3_n660 ) , .A3( u0_u3_n661 ) , .A2( u0_u3_n662 ) , .A1( u0_u3_n663 ) , .ZN( u0_u3_n803 ) );
  NOR2_X1 u0_u3_U360 (.A2( u0_u3_n41 ) , .A1( u0_u3_n783 ) , .ZN( u0_u3_n823 ) );
  AOI21_X1 u0_u3_U361 (.B2( u0_u3_n41 ) , .ZN( u0_u3_n481 ) , .A( u0_u3_n752 ) , .B1( u0_u3_n782 ) );
  NOR2_X1 u0_u3_U362 (.A2( u0_u3_n41 ) , .ZN( u0_u3_n569 ) , .A1( u0_u3_n766 ) );
  NOR2_X1 u0_u3_U363 (.A2( u0_u3_n41 ) , .ZN( u0_u3_n719 ) , .A1( u0_u3_n795 ) );
  NOR2_X1 u0_u3_U364 (.A2( u0_u3_n41 ) , .ZN( u0_u3_n597 ) , .A1( u0_u3_n731 ) );
  AOI21_X1 u0_u3_U365 (.A( u0_u3_n41 ) , .ZN( u0_u3_n555 ) , .B1( u0_u3_n672 ) , .B2( u0_u3_n808 ) );
  NOR2_X1 u0_u3_U366 (.A2( u0_u3_n41 ) , .ZN( u0_u3_n544 ) , .A1( u0_u3_n702 ) );
  NOR2_X1 u0_u3_U367 (.ZN( u0_u3_n583 ) , .A2( u0_u3_n700 ) , .A1( u0_u3_n794 ) );
  NOR4_X1 u0_u3_U368 (.A4( u0_u3_n779 ) , .A3( u0_u3_n780 ) , .A1( u0_u3_n781 ) , .ZN( u0_u3_n802 ) , .A2( u0_u3_n804 ) );
  NAND4_X1 u0_u3_U369 (.A4( u0_u3_n694 ) , .A3( u0_u3_n695 ) , .A1( u0_u3_n696 ) , .ZN( u0_u3_n779 ) , .A2( u0_u3_n874 ) );
  NOR3_X1 u0_u3_U37 (.A3( u0_u3_n654 ) , .A2( u0_u3_n655 ) , .A1( u0_u3_n656 ) , .ZN( u0_u3_n661 ) );
  AOI21_X1 u0_u3_U370 (.ZN( u0_u3_n596 ) , .B1( u0_u3_n753 ) , .A( u0_u3_n795 ) , .B2( u0_u3_n816 ) );
  AOI21_X1 u0_u3_U371 (.A( u0_u3_n815 ) , .B2( u0_u3_n816 ) , .B1( u0_u3_n817 ) , .ZN( u0_u3_n822 ) );
  OAI222_X1 u0_u3_U372 (.ZN( u0_u3_n508 ) , .C2( u0_u3_n628 ) , .B2( u0_u3_n650 ) , .B1( u0_u3_n750 ) , .A2( u0_u3_n751 ) , .C1( u0_u3_n808 ) , .A1( u0_u3_n809 ) );
  AOI21_X1 u0_u3_U373 (.B1( u0_u3_n628 ) , .ZN( u0_u3_n630 ) , .A( u0_u3_n766 ) , .B2( u0_u3_n817 ) );
  AOI21_X1 u0_u3_U374 (.ZN( u0_u3_n652 ) , .B1( u0_u3_n732 ) , .B2( u0_u3_n766 ) , .A( u0_u3_n816 ) );
  OAI21_X1 u0_u3_U375 (.A( u0_u3_n616 ) , .ZN( u0_u3_n619 ) , .B1( u0_u3_n628 ) , .B2( u0_u3_n787 ) );
  NOR2_X1 u0_u3_U376 (.A1( u0_u3_n672 ) , .ZN( u0_u3_n769 ) , .A2( u0_u3_n816 ) );
  NOR2_X1 u0_u3_U377 (.A2( u0_u3_n816 ) , .A1( u0_u3_n818 ) , .ZN( u0_u3_n824 ) );
  NOR2_X1 u0_u3_U378 (.ZN( u0_u3_n581 ) , .A1( u0_u3_n711 ) , .A2( u0_u3_n816 ) );
  NOR2_X1 u0_u3_U379 (.A1( u0_u3_n439 ) , .ZN( u0_u3_n687 ) , .A2( u0_u3_n816 ) );
  NOR3_X1 u0_u3_U38 (.A3( u0_u3_n651 ) , .A2( u0_u3_n652 ) , .A1( u0_u3_n653 ) , .ZN( u0_u3_n662 ) );
  NOR2_X1 u0_u3_U380 (.ZN( u0_u3_n657 ) , .A1( u0_u3_n731 ) , .A2( u0_u3_n816 ) );
  NOR2_X1 u0_u3_U381 (.A1( u0_u3_n702 ) , .ZN( u0_u3_n771 ) , .A2( u0_u3_n816 ) );
  NOR2_X1 u0_u3_U382 (.ZN( u0_u3_n668 ) , .A1( u0_u3_n783 ) , .A2( u0_u3_n816 ) );
  NOR2_X1 u0_u3_U383 (.ZN( u0_u3_n634 ) , .A1( u0_u3_n727 ) , .A2( u0_u3_n816 ) );
  NOR2_X1 u0_u3_U384 (.ZN( u0_u3_n475 ) , .A2( w3_26 ) , .A1( w3_27 ) );
  NOR2_X1 u0_u3_U385 (.ZN( u0_u3_n458 ) , .A1( u0_u3_n831 ) , .A2( w3_27 ) );
  INV_X1 u0_u3_U386 (.ZN( u0_u3_n832 ) , .A( w3_27 ) );
  NOR3_X1 u0_u3_U387 (.A3( u0_u3_n624 ) , .A2( u0_u3_n625 ) , .ZN( u0_u3_n639 ) , .A1( u0_u3_n728 ) );
  NOR4_X1 u0_u3_U388 (.A1( u0_u3_n587 ) , .ZN( u0_u3_n588 ) , .A3( u0_u3_n655 ) , .A2( u0_u3_n665 ) , .A4( u0_u3_n770 ) );
  OAI22_X1 u0_u3_U389 (.ZN( u0_u3_n640 ) , .A1( u0_u3_n702 ) , .B2( u0_u3_n731 ) , .A2( u0_u3_n765 ) , .B1( u0_u3_n819 ) );
  NOR3_X1 u0_u3_U39 (.A3( u0_u3_n657 ) , .A2( u0_u3_n658 ) , .A1( u0_u3_n659 ) , .ZN( u0_u3_n660 ) );
  AOI21_X1 u0_u3_U390 (.ZN( u0_u3_n502 ) , .B1( u0_u3_n683 ) , .A( u0_u3_n815 ) , .B2( u0_u3_n819 ) );
  OAI22_X1 u0_u3_U391 (.A1( u0_u3_n727 ) , .ZN( u0_u3_n729 ) , .B2( u0_u3_n753 ) , .B1( u0_u3_n815 ) , .A2( u0_u3_n819 ) );
  AOI21_X1 u0_u3_U392 (.A( u0_u3_n438 ) , .B2( u0_u3_n819 ) , .B1( u0_u3_n820 ) , .ZN( u0_u3_n821 ) );
  OAI22_X1 u0_u3_U393 (.A1( u0_u3_n438 ) , .ZN( u0_u3_n627 ) , .B1( u0_u3_n672 ) , .B2( u0_u3_n750 ) , .A2( u0_u3_n819 ) );
  NOR2_X1 u0_u3_U394 (.ZN( u0_u3_n522 ) , .A2( u0_u3_n702 ) , .A1( u0_u3_n819 ) );
  NOR2_X1 u0_u3_U395 (.A1( u0_u3_n672 ) , .ZN( u0_u3_n691 ) , .A2( u0_u3_n819 ) );
  NOR2_X1 u0_u3_U396 (.A2( u0_u3_n439 ) , .ZN( u0_u3_n602 ) , .A1( u0_u3_n819 ) );
  NOR2_X1 u0_u3_U397 (.ZN( u0_u3_n534 ) , .A2( u0_u3_n783 ) , .A1( u0_u3_n819 ) );
  NOR2_X1 u0_u3_U398 (.ZN( u0_u3_n561 ) , .A1( u0_u3_n711 ) , .A2( u0_u3_n819 ) );
  NOR2_X1 u0_u3_U399 (.ZN( u0_u3_n688 ) , .A1( u0_u3_n732 ) , .A2( u0_u3_n819 ) );
  NAND2_X1 u0_u3_U4 (.A1( u0_u3_n452 ) , .A2( u0_u3_n463 ) , .ZN( u0_u3_n795 ) );
  NOR4_X1 u0_u3_U40 (.A4( u0_u3_n664 ) , .A3( u0_u3_n665 ) , .A2( u0_u3_n666 ) , .A1( u0_u3_n667 ) , .ZN( u0_u3_n680 ) );
  INV_X1 u0_u3_U400 (.A( u0_u3_n819 ) , .ZN( u0_u3_n834 ) );
  NAND2_X1 u0_u3_U401 (.ZN( u0_u3_n674 ) , .A1( u0_u3_n809 ) , .A2( u0_u3_n819 ) );
  NOR2_X1 u0_u3_U402 (.ZN( u0_u3_n465 ) , .A2( w3_24 ) , .A1( w3_25 ) );
  NOR2_X1 u0_u3_U403 (.ZN( u0_u3_n457 ) , .A1( u0_u3_n830 ) , .A2( w3_24 ) );
  INV_X1 u0_u3_U404 (.ZN( u0_u3_n829 ) , .A( w3_24 ) );
  INV_X1 u0_u3_U405 (.ZN( u0_u3_n850 ) , .A( w3_29 ) );
  NOR2_X1 u0_u3_U406 (.ZN( u0_u3_n451 ) , .A1( u0_u3_n849 ) , .A2( w3_29 ) );
  NAND4_X1 u0_u3_U407 (.ZN( u0_subword_3 ) , .A4( u0_u3_n707 ) , .A3( u0_u3_n708 ) , .A2( u0_u3_n709 ) , .A1( u0_u3_n710 ) );
  INV_X1 u0_u3_U408 (.A( u0_u3_n709 ) , .ZN( u0_u3_n878 ) );
  OAI22_X1 u0_u3_U409 (.B2( u0_u3_n747 ) , .ZN( u0_u3_n749 ) , .A2( u0_u3_n765 ) , .B1( u0_u3_n783 ) , .A1( u0_u3_n795 ) );
  NOR4_X1 u0_u3_U41 (.A4( u0_u3_n668 ) , .A3( u0_u3_n669 ) , .A2( u0_u3_n670 ) , .A1( u0_u3_n671 ) , .ZN( u0_u3_n679 ) );
  OAI22_X1 u0_u3_U410 (.B1( u0_u3_n439 ) , .ZN( u0_u3_n499 ) , .A2( u0_u3_n747 ) , .A1( u0_u3_n783 ) , .B2( u0_u3_n809 ) );
  NOR2_X1 u0_u3_U411 (.ZN( u0_u3_n519 ) , .A1( u0_u3_n711 ) , .A2( u0_u3_n747 ) );
  OAI22_X1 u0_u3_U412 (.ZN( u0_u3_n713 ) , .A2( u0_u3_n731 ) , .B2( u0_u3_n732 ) , .A1( u0_u3_n747 ) , .B1( u0_u3_n816 ) );
  NOR2_X1 u0_u3_U413 (.A2( u0_u3_n747 ) , .ZN( u0_u3_n772 ) , .A1( u0_u3_n815 ) );
  OAI22_X1 u0_u3_U414 (.B1( u0_u3_n443 ) , .ZN( u0_u3_n447 ) , .A2( u0_u3_n731 ) , .A1( u0_u3_n747 ) , .B2( u0_u3_n752 ) );
  NOR2_X1 u0_u3_U415 (.ZN( u0_u3_n550 ) , .A1( u0_u3_n702 ) , .A2( u0_u3_n747 ) );
  NOR2_X1 u0_u3_U416 (.ZN( u0_u3_n556 ) , .A2( u0_u3_n747 ) , .A1( u0_u3_n787 ) );
  NOR2_X1 u0_u3_U417 (.A2( u0_u3_n747 ) , .ZN( u0_u3_n758 ) , .A1( u0_u3_n808 ) );
  NOR2_X1 u0_u3_U418 (.A1( u0_u3_n672 ) , .ZN( u0_u3_n676 ) , .A2( u0_u3_n747 ) );
  NOR2_X1 u0_u3_U419 (.ZN( u0_u3_n533 ) , .A2( u0_u3_n747 ) , .A1( u0_u3_n795 ) );
  NOR4_X1 u0_u3_U42 (.A3( u0_u3_n676 ) , .A1( u0_u3_n677 ) , .ZN( u0_u3_n678 ) , .A4( u0_u3_n718 ) , .A2( u0_u3_n861 ) );
  NOR2_X1 u0_u3_U420 (.ZN( u0_u3_n721 ) , .A2( u0_u3_n727 ) , .A1( u0_u3_n747 ) );
  NOR2_X1 u0_u3_U421 (.ZN( u0_u3_n585 ) , .A1( u0_u3_n747 ) , .A2( u0_u3_n818 ) );
  INV_X1 u0_u3_U422 (.A( u0_u3_n747 ) , .ZN( u0_u3_n839 ) );
  AOI21_X1 u0_u3_U423 (.ZN( u0_u3_n579 ) , .B2( u0_u3_n727 ) , .B1( u0_u3_n751 ) , .A( u0_u3_n788 ) );
  NAND4_X1 u0_u3_U424 (.A4( u0_u3_n636 ) , .A3( u0_u3_n637 ) , .A2( u0_u3_n638 ) , .A1( u0_u3_n639 ) , .ZN( u0_u3_n746 ) );
  INV_X1 u0_u3_U425 (.ZN( u0_u3_n851 ) , .A( w3_30 ) );
  INV_X1 u0_u3_U426 (.ZN( u0_u3_n860 ) , .A( w3_31 ) );
  NAND4_X1 u0_u3_U427 (.ZN( u0_subword_2 ) , .A4( u0_u3_n646 ) , .A3( u0_u3_n647 ) , .A2( u0_u3_n648 ) , .A1( u0_u3_n649 ) );
  AOI211_X1 u0_u3_U428 (.A( u0_u3_n640 ) , .ZN( u0_u3_n648 ) , .B( u0_u3_n746 ) , .C2( u0_u3_n841 ) , .C1( u0_u3_n856 ) );
  NOR2_X1 u0_u3_U429 (.A2( u0_u3_n41 ) , .ZN( u0_u3_n603 ) , .A1( u0_u3_n787 ) );
  NOR4_X1 u0_u3_U43 (.A1( u0_u3_n469 ) , .ZN( u0_u3_n470 ) , .A4( u0_u3_n545 ) , .A2( u0_u3_n557 ) , .A3( u0_u3_n617 ) );
  OAI222_X1 u0_u3_U430 (.A2( u0_u3_n672 ) , .ZN( u0_u3_n677 ) , .B1( u0_u3_n750 ) , .B2( u0_u3_n787 ) , .C2( u0_u3_n791 ) , .C1( u0_u3_n818 ) , .A1( u0_u3_n820 ) );
  NOR2_X1 u0_u3_U431 (.ZN( u0_u3_n613 ) , .A1( u0_u3_n787 ) , .A2( u0_u3_n819 ) );
  AOI21_X1 u0_u3_U432 (.A( u0_u3_n41 ) , .ZN( u0_u3_n503 ) , .B1( u0_u3_n711 ) , .B2( u0_u3_n789 ) );
  OAI22_X1 u0_u3_U433 (.ZN( u0_u3_n593 ) , .B1( u0_u3_n733 ) , .B2( u0_u3_n752 ) , .A2( u0_u3_n789 ) , .A1( u0_u3_n806 ) );
  NOR2_X1 u0_u3_U434 (.ZN( u0_u3_n656 ) , .A1( u0_u3_n765 ) , .A2( u0_u3_n789 ) );
  NAND2_X1 u0_u3_U435 (.A2( u0_u3_n752 ) , .A1( u0_u3_n789 ) , .ZN( u0_u3_n812 ) );
  NOR2_X1 u0_u3_U436 (.ZN( u0_u3_n557 ) , .A1( u0_u3_n789 ) , .A2( u0_u3_n816 ) );
  NAND3_X1 u0_u3_U437 (.ZN( u0_subword_6 ) , .A3( u0_u3_n800 ) , .A2( u0_u3_n801 ) , .A1( u0_u3_n802 ) );
  NAND3_X1 u0_u3_U438 (.ZN( u0_subword_5 ) , .A3( u0_u3_n761 ) , .A2( u0_u3_n762 ) , .A1( u0_u3_n763 ) );
  NAND3_X1 u0_u3_U439 (.ZN( u0_subword_4 ) , .A3( u0_u3_n741 ) , .A2( u0_u3_n742 ) , .A1( u0_u3_n743 ) );
  AOI221_X1 u0_u3_U44 (.ZN( u0_u3_n471 ) , .C2( u0_u3_n717 ) , .B2( u0_u3_n834 ) , .C1( u0_u3_n847 ) , .B1( u0_u3_n862 ) , .A( u0_u3_n866 ) );
  NAND3_X1 u0_u3_U440 (.A3( u0_u3_n678 ) , .A2( u0_u3_n679 ) , .A1( u0_u3_n680 ) , .ZN( u0_u3_n810 ) );
  NAND3_X1 u0_u3_U441 (.ZN( u0_u3_n641 ) , .A3( u0_u3_n711 ) , .A2( u0_u3_n727 ) , .A1( u0_u3_n795 ) );
  NAND3_X1 u0_u3_U442 (.A3( u0_u3_n621 ) , .A2( u0_u3_n622 ) , .A1( u0_u3_n623 ) , .ZN( u0_u3_n728 ) );
  NAND3_X1 u0_u3_U443 (.A3( u0_u3_n588 ) , .A2( u0_u3_n589 ) , .A1( u0_u3_n590 ) , .ZN( u0_u3_n624 ) );
  NAND3_X1 u0_u3_U444 (.ZN( u0_u3_n568 ) , .A3( u0_u3_n683 ) , .A2( u0_u3_n753 ) , .A1( u0_u3_n788 ) );
  NAND3_X1 u0_u3_U445 (.A3( u0_u3_n526 ) , .A2( u0_u3_n527 ) , .A1( u0_u3_n528 ) , .ZN( u0_u3_n745 ) );
  NAND3_X1 u0_u3_U446 (.A3( u0_u3_n515 ) , .A1( u0_u3_n516 ) , .ZN( u0_u3_n611 ) , .A2( u0_u3_n873 ) );
  NAND3_X1 u0_u3_U447 (.A3( u0_u3_n470 ) , .A2( u0_u3_n471 ) , .A1( u0_u3_n472 ) , .ZN( u0_u3_n780 ) );
  NOR2_X1 u0_u3_U448 (.ZN( u0_u3_n615 ) , .A1( u0_u3_n782 ) , .A2( u0_u3_n789 ) );
  NOR2_X1 u0_u3_U449 (.ZN( u0_u3_n720 ) , .A2( u0_u3_n747 ) , .A1( u0_u3_n789 ) );
  NOR4_X1 u0_u3_U45 (.A4( u0_u3_n517 ) , .A3( u0_u3_n518 ) , .A2( u0_u3_n519 ) , .A1( u0_u3_n520 ) , .ZN( u0_u3_n527 ) );
  NOR2_X1 u0_u3_U450 (.ZN( u0_u3_n704 ) , .A2( u0_u3_n789 ) , .A1( u0_u3_n820 ) );
  NOR2_X1 u0_u3_U451 (.A1( u0_u3_n733 ) , .ZN( u0_u3_n768 ) , .A2( u0_u3_n789 ) );
  INV_X1 u0_u3_U452 (.ZN( u0_u3_n849 ) , .A( w3_28 ) );
  NOR4_X1 u0_u3_U46 (.A3( u0_u3_n524 ) , .A1( u0_u3_n525 ) , .ZN( u0_u3_n526 ) , .A2( u0_u3_n676 ) , .A4( u0_u3_n772 ) );
  NAND4_X1 u0_u3_U47 (.A4( u0_u3_n576 ) , .A3( u0_u3_n577 ) , .A1( u0_u3_n578 ) , .ZN( u0_u3_n726 ) , .A2( u0_u3_n876 ) );
  NOR4_X1 u0_u3_U48 (.A4( u0_u3_n572 ) , .A3( u0_u3_n573 ) , .A2( u0_u3_n574 ) , .A1( u0_u3_n575 ) , .ZN( u0_u3_n576 ) );
  INV_X1 u0_u3_U49 (.A( u0_u3_n610 ) , .ZN( u0_u3_n876 ) );
  NAND2_X1 u0_u3_U5 (.A1( u0_u3_n456 ) , .A2( u0_u3_n475 ) , .ZN( u0_u3_n788 ) );
  NAND4_X1 u0_u3_U50 (.A4( u0_u3_n459 ) , .A3( u0_u3_n460 ) , .A2( u0_u3_n461 ) , .A1( u0_u3_n462 ) , .ZN( u0_u3_n682 ) );
  NOR3_X1 u0_u3_U51 (.ZN( u0_u3_n460 ) , .A3( u0_u3_n533 ) , .A1( u0_u3_n558 ) , .A2( u0_u3_n573 ) );
  NOR4_X1 u0_u3_U52 (.ZN( u0_u3_n459 ) , .A2( u0_u3_n520 ) , .A1( u0_u3_n546 ) , .A3( u0_u3_n582 ) , .A4( u0_u3_n618 ) );
  NOR4_X1 u0_u3_U53 (.ZN( u0_u3_n461 ) , .A2( u0_u3_n512 ) , .A1( u0_u3_n602 ) , .A4( u0_u3_n631 ) , .A3( u0_u3_n714 ) );
  NAND4_X1 u0_u3_U54 (.A4( u0_u3_n722 ) , .A3( u0_u3_n723 ) , .A2( u0_u3_n724 ) , .ZN( u0_u3_n744 ) , .A1( u0_u3_n859 ) );
  INV_X1 u0_u3_U55 (.A( u0_u3_n712 ) , .ZN( u0_u3_n859 ) );
  NOR4_X1 u0_u3_U56 (.A4( u0_u3_n718 ) , .A3( u0_u3_n719 ) , .A2( u0_u3_n720 ) , .A1( u0_u3_n721 ) , .ZN( u0_u3_n722 ) );
  NOR3_X1 u0_u3_U57 (.ZN( u0_u3_n483 ) , .A2( u0_u3_n511 ) , .A3( u0_u3_n604 ) , .A1( u0_u3_n613 ) );
  NOR4_X1 u0_u3_U58 (.ZN( u0_u3_n484 ) , .A3( u0_u3_n535 ) , .A4( u0_u3_n548 ) , .A2( u0_u3_n570 ) , .A1( u0_u3_n720 ) );
  AOI211_X1 u0_u3_U59 (.B( u0_u3_n480 ) , .A( u0_u3_n481 ) , .ZN( u0_u3_n485 ) , .C2( u0_u3_n836 ) , .C1( u0_u3_n863 ) );
  NOR3_X1 u0_u3_U6 (.ZN( u0_u3_n601 ) , .A1( u0_u3_n611 ) , .A3( u0_u3_n726 ) , .A2( u0_u3_n745 ) );
  INV_X1 u0_u3_U60 (.A( u0_u3_n682 ) , .ZN( u0_u3_n874 ) );
  NOR4_X1 u0_u3_U61 (.A4( u0_u3_n690 ) , .A3( u0_u3_n691 ) , .A2( u0_u3_n692 ) , .A1( u0_u3_n693 ) , .ZN( u0_u3_n694 ) );
  AOI221_X1 u0_u3_U62 (.A( u0_u3_n684 ) , .ZN( u0_u3_n695 ) , .B2( u0_u3_n842 ) , .C1( u0_u3_n844 ) , .C2( u0_u3_n864 ) , .B1( u0_u3_n867 ) );
  NAND4_X1 u0_u3_U63 (.A4( u0_u3_n476 ) , .A3( u0_u3_n477 ) , .A2( u0_u3_n478 ) , .A1( u0_u3_n479 ) , .ZN( u0_u3_n681 ) );
  NOR4_X1 u0_u3_U64 (.A4( u0_u3_n473 ) , .ZN( u0_u3_n479 ) , .A3( u0_u3_n559 ) , .A1( u0_u3_n738 ) , .A2( u0_u3_n758 ) );
  NOR4_X1 u0_u3_U65 (.ZN( u0_u3_n477 ) , .A1( u0_u3_n509 ) , .A3( u0_u3_n547 ) , .A2( u0_u3_n586 ) , .A4( u0_u3_n719 ) );
  NOR4_X1 u0_u3_U66 (.ZN( u0_u3_n476 ) , .A2( u0_u3_n524 ) , .A4( u0_u3_n597 ) , .A1( u0_u3_n612 ) , .A3( u0_u3_n632 ) );
  NAND4_X1 u0_u3_U67 (.A4( u0_u3_n551 ) , .A3( u0_u3_n552 ) , .A2( u0_u3_n553 ) , .A1( u0_u3_n554 ) , .ZN( u0_u3_n748 ) );
  AOI211_X1 u0_u3_U68 (.B( u0_u3_n542 ) , .A( u0_u3_n543 ) , .ZN( u0_u3_n554 ) , .C2( u0_u3_n841 ) , .C1( u0_u3_n853 ) );
  NOR3_X1 u0_u3_U69 (.ZN( u0_u3_n552 ) , .A2( u0_u3_n654 ) , .A1( u0_u3_n670 ) , .A3( u0_u3_n774 ) );
  NOR3_X1 u0_u3_U7 (.ZN( u0_u3_n507 ) , .A2( u0_u3_n682 ) , .A3( u0_u3_n780 ) , .A1( u0_u3_n878 ) );
  NOR4_X1 u0_u3_U70 (.A4( u0_u3_n544 ) , .A3( u0_u3_n545 ) , .A2( u0_u3_n546 ) , .ZN( u0_u3_n553 ) , .A1( u0_u3_n691 ) );
  NOR4_X1 u0_u3_U71 (.A4( u0_u3_n612 ) , .A3( u0_u3_n613 ) , .A2( u0_u3_n614 ) , .A1( u0_u3_n615 ) , .ZN( u0_u3_n622 ) );
  NOR4_X1 u0_u3_U72 (.ZN( u0_u3_n623 ) , .A1( u0_u3_n659 ) , .A3( u0_u3_n669 ) , .A4( u0_u3_n685 ) , .A2( u0_u3_n769 ) );
  INV_X1 u0_u3_U73 (.A( u0_u3_n765 ) , .ZN( u0_u3_n833 ) );
  NOR2_X1 u0_u3_U74 (.ZN( u0_u3_n650 ) , .A1( u0_u3_n856 ) , .A2( u0_u3_n870 ) );
  NOR4_X1 u0_u3_U75 (.A4( u0_u3_n580 ) , .A3( u0_u3_n581 ) , .A2( u0_u3_n582 ) , .ZN( u0_u3_n589 ) , .A1( u0_u3_n686 ) );
  INV_X1 u0_u3_U76 (.A( u0_u3_n818 ) , .ZN( u0_u3_n857 ) );
  OR4_X1 u0_u3_U77 (.A4( u0_u3_n685 ) , .A3( u0_u3_n686 ) , .A2( u0_u3_n687 ) , .A1( u0_u3_n688 ) , .ZN( u0_u3_n693 ) );
  OR4_X1 u0_u3_U78 (.ZN( u0_u3_n469 ) , .A4( u0_u3_n521 ) , .A3( u0_u3_n532 ) , .A2( u0_u3_n581 ) , .A1( u0_u3_n715 ) );
  OR4_X1 u0_u3_U79 (.A4( u0_u3_n569 ) , .A3( u0_u3_n570 ) , .A2( u0_u3_n571 ) , .ZN( u0_u3_n575 ) , .A1( u0_u3_n668 ) );
  NOR3_X1 u0_u3_U8 (.A2( u0_u3_n610 ) , .A1( u0_u3_n611 ) , .ZN( u0_u3_n649 ) , .A3( u0_u3_n725 ) );
  OR4_X1 u0_u3_U80 (.A4( u0_u3_n521 ) , .A2( u0_u3_n522 ) , .A1( u0_u3_n523 ) , .ZN( u0_u3_n525 ) , .A3( u0_u3_n824 ) );
  OR4_X1 u0_u3_U81 (.A4( u0_u3_n583 ) , .A3( u0_u3_n584 ) , .A2( u0_u3_n585 ) , .A1( u0_u3_n586 ) , .ZN( u0_u3_n587 ) );
  OR4_X1 u0_u3_U82 (.ZN( u0_u3_n495 ) , .A4( u0_u3_n537 ) , .A2( u0_u3_n550 ) , .A1( u0_u3_n562 ) , .A3( u0_u3_n635 ) );
  NOR4_X1 u0_u3_U83 (.A4( u0_u3_n512 ) , .A2( u0_u3_n513 ) , .A1( u0_u3_n514 ) , .ZN( u0_u3_n515 ) , .A3( u0_u3_n673 ) );
  INV_X1 u0_u3_U84 (.A( u0_u3_n508 ) , .ZN( u0_u3_n873 ) );
  OR3_X1 u0_u3_U85 (.A3( u0_u3_n509 ) , .A2( u0_u3_n510 ) , .A1( u0_u3_n511 ) , .ZN( u0_u3_n514 ) );
  INV_X1 u0_u3_U86 (.A( u0_u3_n757 ) , .ZN( u0_u3_n871 ) );
  AOI221_X1 u0_u3_U87 (.A( u0_u3_n716 ) , .B2( u0_u3_n717 ) , .ZN( u0_u3_n723 ) , .C1( u0_u3_n835 ) , .B1( u0_u3_n841 ) , .C2( u0_u3_n865 ) );
  OR2_X1 u0_u3_U88 (.A2( u0_u3_n714 ) , .A1( u0_u3_n715 ) , .ZN( u0_u3_n716 ) );
  INV_X1 u0_u3_U89 (.A( u0_u3_n466 ) , .ZN( u0_u3_n866 ) );
  NOR3_X1 u0_u3_U9 (.A3( u0_u3_n725 ) , .A1( u0_u3_n726 ) , .ZN( u0_u3_n743 ) , .A2( u0_u3_n744 ) );
  NAND2_X1 u0_u3_U90 (.A1( u0_u3_n454 ) , .A2( u0_u3_n456 ) , .ZN( u0_u3_n765 ) );
  AOI22_X1 u0_u3_U91 (.ZN( u0_u3_n699 ) , .A1( u0_u3_n833 ) , .B2( u0_u3_n845 ) , .A2( u0_u3_n867 ) , .B1( u0_u3_n870 ) );
  NOR3_X1 u0_u3_U92 (.ZN( u0_u3_n755 ) , .A2( u0_u3_n855 ) , .A1( u0_u3_n865 ) , .A3( u0_u3_n867 ) );
  NOR2_X1 u0_u3_U93 (.ZN( u0_u3_n754 ) , .A2( u0_u3_n854 ) , .A1( u0_u3_n862 ) );
  AOI211_X1 u0_u3_U94 (.A( u0_u3_n499 ) , .ZN( u0_u3_n506 ) , .B( u0_u3_n805 ) , .C2( u0_u3_n841 ) , .C1( u0_u3_n853 ) );
  AOI211_X1 u0_u3_U95 (.B( u0_u3_n810 ) , .A( u0_u3_n811 ) , .ZN( u0_u3_n827 ) , .C1( u0_u3_n844 ) , .C2( u0_u3_n852 ) );
  NAND2_X1 u0_u3_U96 (.A1( u0_u3_n450 ) , .A2( u0_u3_n468 ) , .ZN( u0_u3_n752 ) );
  INV_X1 u0_u3_U97 (.A( u0_u3_n733 ) , .ZN( u0_u3_n841 ) );
  AOI221_X1 u0_u3_U98 (.B2( u0_u3_n440 ) , .A( u0_u3_n492 ) , .ZN( u0_u3_n497 ) , .C2( u0_u3_n843 ) , .C1( u0_u3_n853 ) , .B1( u0_u3_n862 ) );
  INV_X1 u0_u3_U99 (.A( u0_u3_n781 ) , .ZN( u0_u3_n869 ) );
endmodule

