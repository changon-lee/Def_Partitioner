module aes_aes_die_4 ( sa03_0, sa03_1, sa03_2, sa03_3, sa03_4, sa03_5, sa03_6, sa03_7, sa20_0, 
       sa20_1, sa20_2, sa20_3, sa20_4, sa20_5, sa20_6, sa20_7, sa23_0, sa23_1, 
       sa23_2, sa23_3, sa23_4, sa23_5, sa23_6, sa23_7, sa30_0, sa30_1, sa30_2, 
       sa30_3, sa30_4, sa30_5, sa30_6, sa30_7, w3_0, w3_1, w3_2, w3_3, 
       w3_4, w3_5, w3_6, w3_7, sa03_sr_0, sa03_sr_1, sa03_sr_2, sa03_sr_3, sa03_sr_4, sa03_sr_5, sa03_sr_6, sa03_sr_7, sa21_sr_0, 
        sa21_sr_1, sa21_sr_2, sa21_sr_3, sa21_sr_4, sa21_sr_5, sa21_sr_6, sa21_sr_7, sa22_sr_0, sa22_sr_1, 
        sa22_sr_2, sa22_sr_3, sa22_sr_4, sa22_sr_5, sa22_sr_6, sa22_sr_7, sa31_sr_0, sa31_sr_1, sa31_sr_2, 
        sa31_sr_3, sa31_sr_4, sa31_sr_5, sa31_sr_6, sa31_sr_7, u0_subword_10, u0_subword_11, u0_subword_12, u0_subword_13, 
        u0_subword_14, u0_subword_15, u0_subword_8, u0_subword_9 );
  input sa03_0, sa03_1, sa03_2, sa03_3, sa03_4, sa03_5, sa03_6, sa03_7, sa20_0, 
        sa20_1, sa20_2, sa20_3, sa20_4, sa20_5, sa20_6, sa20_7, sa23_0, sa23_1, 
        sa23_2, sa23_3, sa23_4, sa23_5, sa23_6, sa23_7, sa30_0, sa30_1, sa30_2, 
        sa30_3, sa30_4, sa30_5, sa30_6, sa30_7, w3_0, w3_1, w3_2, w3_3, 
        w3_4, w3_5, w3_6, w3_7;
  output sa03_sr_0, sa03_sr_1, sa03_sr_2, sa03_sr_3, sa03_sr_4, sa03_sr_5, sa03_sr_6, sa03_sr_7, sa21_sr_0, 
        sa21_sr_1, sa21_sr_2, sa21_sr_3, sa21_sr_4, sa21_sr_5, sa21_sr_6, sa21_sr_7, sa22_sr_0, sa22_sr_1, 
        sa22_sr_2, sa22_sr_3, sa22_sr_4, sa22_sr_5, sa22_sr_6, sa22_sr_7, sa31_sr_0, sa31_sr_1, sa31_sr_2, 
        sa31_sr_3, sa31_sr_4, sa31_sr_5, sa31_sr_6, sa31_sr_7, u0_subword_10, u0_subword_11, u0_subword_12, u0_subword_13, 
        u0_subword_14, u0_subword_15, u0_subword_8, u0_subword_9;
  wire u0_u2_n438, u0_u2_n439, u0_u2_n440, u0_u2_n441, u0_u2_n442, u0_u2_n443, u0_u2_n444, u0_u2_n445, u0_u2_n446, 
       u0_u2_n447, u0_u2_n448, u0_u2_n449, u0_u2_n450, u0_u2_n451, u0_u2_n452, u0_u2_n453, u0_u2_n454, u0_u2_n455, 
       u0_u2_n456, u0_u2_n457, u0_u2_n458, u0_u2_n459, u0_u2_n460, u0_u2_n461, u0_u2_n462, u0_u2_n463, u0_u2_n464, 
       u0_u2_n465, u0_u2_n466, u0_u2_n467, u0_u2_n468, u0_u2_n469, u0_u2_n470, u0_u2_n471, u0_u2_n472, u0_u2_n473, 
       u0_u2_n474, u0_u2_n475, u0_u2_n476, u0_u2_n477, u0_u2_n478, u0_u2_n479, u0_u2_n480, u0_u2_n481, u0_u2_n482, 
       u0_u2_n483, u0_u2_n484, u0_u2_n485, u0_u2_n486, u0_u2_n487, u0_u2_n488, u0_u2_n489, u0_u2_n490, u0_u2_n491, 
       u0_u2_n492, u0_u2_n493, u0_u2_n494, u0_u2_n495, u0_u2_n496, u0_u2_n497, u0_u2_n498, u0_u2_n499, u0_u2_n500, 
       u0_u2_n501, u0_u2_n502, u0_u2_n503, u0_u2_n504, u0_u2_n505, u0_u2_n506, u0_u2_n507, u0_u2_n508, u0_u2_n509, 
       u0_u2_n510, u0_u2_n511, u0_u2_n512, u0_u2_n513, u0_u2_n514, u0_u2_n515, u0_u2_n516, u0_u2_n517, u0_u2_n518, 
       u0_u2_n519, u0_u2_n520, u0_u2_n521, u0_u2_n522, u0_u2_n523, u0_u2_n524, u0_u2_n525, u0_u2_n526, u0_u2_n527, 
       u0_u2_n528, u0_u2_n529, u0_u2_n530, u0_u2_n531, u0_u2_n532, u0_u2_n533, u0_u2_n534, u0_u2_n535, u0_u2_n536, 
       u0_u2_n537, u0_u2_n538, u0_u2_n539, u0_u2_n540, u0_u2_n541, u0_u2_n542, u0_u2_n543, u0_u2_n544, u0_u2_n545, 
       u0_u2_n546, u0_u2_n547, u0_u2_n548, u0_u2_n549, u0_u2_n550, u0_u2_n551, u0_u2_n552, u0_u2_n553, u0_u2_n554, 
       u0_u2_n555, u0_u2_n556, u0_u2_n557, u0_u2_n558, u0_u2_n559, u0_u2_n560, u0_u2_n561, u0_u2_n562, u0_u2_n563, 
       u0_u2_n564, u0_u2_n565, u0_u2_n566, u0_u2_n567, u0_u2_n568, u0_u2_n569, u0_u2_n570, u0_u2_n571, u0_u2_n572, 
       u0_u2_n573, u0_u2_n574, u0_u2_n575, u0_u2_n576, u0_u2_n577, u0_u2_n578, u0_u2_n579, u0_u2_n580, u0_u2_n581, 
       u0_u2_n582, u0_u2_n583, u0_u2_n584, u0_u2_n585, u0_u2_n586, u0_u2_n587, u0_u2_n588, u0_u2_n589, u0_u2_n590, 
       u0_u2_n591, u0_u2_n592, u0_u2_n593, u0_u2_n594, u0_u2_n595, u0_u2_n596, u0_u2_n597, u0_u2_n598, u0_u2_n599, 
       u0_u2_n600, u0_u2_n601, u0_u2_n602, u0_u2_n603, u0_u2_n604, u0_u2_n605, u0_u2_n606, u0_u2_n607, u0_u2_n608, 
       u0_u2_n609, u0_u2_n610, u0_u2_n611, u0_u2_n612, u0_u2_n613, u0_u2_n614, u0_u2_n615, u0_u2_n616, u0_u2_n617, 
       u0_u2_n618, u0_u2_n619, u0_u2_n620, u0_u2_n621, u0_u2_n622, u0_u2_n623, u0_u2_n624, u0_u2_n625, u0_u2_n626, 
       u0_u2_n627, u0_u2_n628, u0_u2_n629, u0_u2_n630, u0_u2_n631, u0_u2_n632, u0_u2_n633, u0_u2_n634, u0_u2_n635, 
       u0_u2_n636, u0_u2_n637, u0_u2_n638, u0_u2_n639, u0_u2_n640, u0_u2_n641, u0_u2_n642, u0_u2_n643, u0_u2_n644, 
       u0_u2_n645, u0_u2_n646, u0_u2_n647, u0_u2_n648, u0_u2_n649, u0_u2_n650, u0_u2_n651, u0_u2_n652, u0_u2_n653, 
       u0_u2_n654, u0_u2_n655, u0_u2_n656, u0_u2_n657, u0_u2_n658, u0_u2_n659, u0_u2_n660, u0_u2_n661, u0_u2_n662, 
       u0_u2_n663, u0_u2_n664, u0_u2_n665, u0_u2_n666, u0_u2_n667, u0_u2_n668, u0_u2_n669, u0_u2_n670, u0_u2_n671, 
       u0_u2_n672, u0_u2_n673, u0_u2_n674, u0_u2_n675, u0_u2_n676, u0_u2_n677, u0_u2_n678, u0_u2_n679, u0_u2_n680, 
       u0_u2_n681, u0_u2_n682, u0_u2_n683, u0_u2_n684, u0_u2_n685, u0_u2_n686, u0_u2_n687, u0_u2_n688, u0_u2_n689, 
       u0_u2_n690, u0_u2_n691, u0_u2_n692, u0_u2_n693, u0_u2_n694, u0_u2_n695, u0_u2_n696, u0_u2_n697, u0_u2_n698, 
       u0_u2_n699, u0_u2_n700, u0_u2_n701, u0_u2_n702, u0_u2_n703, u0_u2_n704, u0_u2_n705, u0_u2_n706, u0_u2_n707, 
       u0_u2_n708, u0_u2_n709, u0_u2_n710, u0_u2_n711, u0_u2_n712, u0_u2_n713, u0_u2_n714, u0_u2_n715, u0_u2_n716, 
       u0_u2_n717, u0_u2_n718, u0_u2_n719, u0_u2_n720, u0_u2_n721, u0_u2_n722, u0_u2_n723, u0_u2_n724, u0_u2_n725, 
       u0_u2_n726, u0_u2_n727, u0_u2_n728, u0_u2_n729, u0_u2_n730, u0_u2_n731, u0_u2_n732, u0_u2_n733, u0_u2_n734, 
       u0_u2_n735, u0_u2_n736, u0_u2_n737, u0_u2_n738, u0_u2_n739, u0_u2_n740, u0_u2_n741, u0_u2_n742, u0_u2_n743, 
       u0_u2_n744, u0_u2_n745, u0_u2_n746, u0_u2_n747, u0_u2_n748, u0_u2_n749, u0_u2_n750, u0_u2_n751, u0_u2_n752, 
       u0_u2_n753, u0_u2_n754, u0_u2_n755, u0_u2_n756, u0_u2_n757, u0_u2_n758, u0_u2_n759, u0_u2_n760, u0_u2_n761, 
       u0_u2_n762, u0_u2_n763, u0_u2_n764, u0_u2_n765, u0_u2_n766, u0_u2_n767, u0_u2_n768, u0_u2_n769, u0_u2_n770, 
       u0_u2_n771, u0_u2_n772, u0_u2_n773, u0_u2_n774, u0_u2_n775, u0_u2_n776, u0_u2_n777, u0_u2_n778, u0_u2_n779, 
       u0_u2_n780, u0_u2_n781, u0_u2_n782, u0_u2_n783, u0_u2_n784, u0_u2_n785, u0_u2_n786, u0_u2_n787, u0_u2_n788, 
       u0_u2_n789, u0_u2_n790, u0_u2_n791, u0_u2_n792, u0_u2_n793, u0_u2_n794, u0_u2_n795, u0_u2_n796, u0_u2_n797, 
       u0_u2_n798, u0_u2_n799, u0_u2_n800, u0_u2_n801, u0_u2_n802, u0_u2_n803, u0_u2_n804, u0_u2_n805, u0_u2_n806, 
       u0_u2_n807, u0_u2_n808, u0_u2_n809, u0_u2_n810, u0_u2_n811, u0_u2_n812, u0_u2_n813, u0_u2_n814, u0_u2_n815, 
       u0_u2_n816, u0_u2_n817, u0_u2_n818, u0_u2_n819, u0_u2_n820, u0_u2_n821, u0_u2_n822, u0_u2_n823, u0_u2_n824, 
       u0_u2_n825, u0_u2_n826, u0_u2_n827, u0_u2_n828, u0_u2_n829, u0_u2_n830, u0_u2_n831, u0_u2_n832, u0_u2_n833, 
       u0_u2_n834, u0_u2_n835, u0_u2_n836, u0_u2_n837, u0_u2_n838, u0_u2_n839, u0_u2_n840, u0_u2_n841, u0_u2_n842, 
       u0_u2_n843, u0_u2_n844, u0_u2_n845, u0_u2_n846, u0_u2_n847, u0_u2_n848, u0_u2_n849, u0_u2_n850, u0_u2_n851, 
       u0_u2_n852, u0_u2_n853, u0_u2_n854, u0_u2_n855, u0_u2_n856, u0_u2_n857, u0_u2_n858, u0_u2_n859, u0_u2_n860, 
       u0_u2_n861, u0_u2_n862, u0_u2_n863, u0_u2_n864, u0_u2_n865, u0_u2_n866, u0_u2_n867, u0_u2_n868, u0_u2_n869, 
       u0_u2_n870, u0_u2_n871, u0_u2_n872, u0_u2_n873, u0_u2_n874, u0_u2_n875, u0_u2_n876, u0_u2_n877, u0_u2_n878, 
       u0_u2_n879, u0_u2_n880, u0_u2_n881, u0_u2_n882, u0_u2_n883, us03_n438, us03_n439, us03_n440, us03_n441, 
       us03_n442, us03_n443, us03_n444, us03_n445, us03_n446, us03_n447, us03_n448, us03_n449, us03_n450, 
       us03_n451, us03_n452, us03_n453, us03_n454, us03_n455, us03_n456, us03_n457, us03_n458, us03_n459, 
       us03_n460, us03_n461, us03_n462, us03_n463, us03_n464, us03_n465, us03_n466, us03_n467, us03_n468, 
       us03_n469, us03_n470, us03_n471, us03_n472, us03_n473, us03_n474, us03_n475, us03_n476, us03_n477, 
       us03_n478, us03_n479, us03_n480, us03_n481, us03_n482, us03_n483, us03_n484, us03_n485, us03_n486, 
       us03_n487, us03_n488, us03_n489, us03_n490, us03_n491, us03_n492, us03_n493, us03_n494, us03_n495, 
       us03_n496, us03_n497, us03_n498, us03_n499, us03_n500, us03_n501, us03_n502, us03_n503, us03_n504, 
       us03_n505, us03_n506, us03_n507, us03_n508, us03_n509, us03_n510, us03_n511, us03_n512, us03_n513, 
       us03_n514, us03_n515, us03_n516, us03_n517, us03_n518, us03_n519, us03_n520, us03_n521, us03_n522, 
       us03_n523, us03_n524, us03_n525, us03_n526, us03_n527, us03_n528, us03_n529, us03_n530, us03_n531, 
       us03_n532, us03_n533, us03_n534, us03_n535, us03_n536, us03_n537, us03_n538, us03_n539, us03_n540, 
       us03_n541, us03_n542, us03_n543, us03_n544, us03_n545, us03_n546, us03_n547, us03_n548, us03_n549, 
       us03_n550, us03_n551, us03_n552, us03_n553, us03_n554, us03_n555, us03_n556, us03_n557, us03_n558, 
       us03_n559, us03_n560, us03_n561, us03_n562, us03_n563, us03_n564, us03_n565, us03_n566, us03_n567, 
       us03_n568, us03_n569, us03_n570, us03_n571, us03_n572, us03_n573, us03_n574, us03_n575, us03_n576, 
       us03_n577, us03_n578, us03_n579, us03_n580, us03_n581, us03_n582, us03_n583, us03_n584, us03_n585, 
       us03_n586, us03_n587, us03_n588, us03_n589, us03_n590, us03_n591, us03_n592, us03_n593, us03_n594, 
       us03_n595, us03_n596, us03_n597, us03_n598, us03_n599, us03_n600, us03_n601, us03_n602, us03_n603, 
       us03_n604, us03_n605, us03_n606, us03_n607, us03_n608, us03_n609, us03_n610, us03_n611, us03_n612, 
       us03_n613, us03_n614, us03_n615, us03_n616, us03_n617, us03_n618, us03_n619, us03_n620, us03_n621, 
       us03_n622, us03_n623, us03_n624, us03_n625, us03_n626, us03_n627, us03_n628, us03_n629, us03_n630, 
       us03_n631, us03_n632, us03_n633, us03_n634, us03_n635, us03_n636, us03_n637, us03_n638, us03_n639, 
       us03_n640, us03_n641, us03_n642, us03_n643, us03_n644, us03_n645, us03_n646, us03_n647, us03_n648, 
       us03_n649, us03_n650, us03_n651, us03_n652, us03_n653, us03_n654, us03_n655, us03_n656, us03_n657, 
       us03_n658, us03_n659, us03_n660, us03_n661, us03_n662, us03_n663, us03_n664, us03_n665, us03_n666, 
       us03_n667, us03_n668, us03_n669, us03_n670, us03_n671, us03_n672, us03_n673, us03_n674, us03_n675, 
       us03_n676, us03_n677, us03_n678, us03_n679, us03_n680, us03_n681, us03_n682, us03_n683, us03_n684, 
       us03_n685, us03_n686, us03_n687, us03_n688, us03_n689, us03_n690, us03_n691, us03_n692, us03_n693, 
       us03_n694, us03_n695, us03_n696, us03_n697, us03_n698, us03_n699, us03_n700, us03_n701, us03_n702, 
       us03_n703, us03_n704, us03_n705, us03_n706, us03_n707, us03_n708, us03_n709, us03_n710, us03_n711, 
       us03_n712, us03_n713, us03_n714, us03_n715, us03_n716, us03_n717, us03_n718, us03_n719, us03_n720, 
       us03_n721, us03_n722, us03_n723, us03_n724, us03_n725, us03_n726, us03_n727, us03_n728, us03_n729, 
       us03_n730, us03_n731, us03_n732, us03_n733, us03_n734, us03_n735, us03_n736, us03_n737, us03_n738, 
       us03_n739, us03_n740, us03_n741, us03_n742, us03_n743, us03_n744, us03_n745, us03_n746, us03_n747, 
       us03_n748, us03_n749, us03_n750, us03_n751, us03_n752, us03_n753, us03_n754, us03_n755, us03_n756, 
       us03_n757, us03_n758, us03_n759, us03_n760, us03_n761, us03_n762, us03_n763, us03_n764, us03_n765, 
       us03_n766, us03_n767, us03_n768, us03_n769, us03_n770, us03_n771, us03_n772, us03_n773, us03_n774, 
       us03_n775, us03_n776, us03_n777, us03_n778, us03_n779, us03_n780, us03_n781, us03_n782, us03_n783, 
       us03_n784, us03_n785, us03_n786, us03_n787, us03_n788, us03_n789, us03_n790, us03_n791, us03_n792, 
       us03_n793, us03_n794, us03_n795, us03_n796, us03_n797, us03_n798, us03_n799, us03_n800, us03_n801, 
       us03_n802, us03_n803, us03_n804, us03_n805, us03_n806, us03_n807, us03_n808, us03_n809, us03_n810, 
       us03_n811, us03_n812, us03_n813, us03_n814, us03_n815, us03_n816, us03_n817, us03_n818, us03_n819, 
       us03_n820, us03_n821, us03_n822, us03_n823, us03_n824, us03_n825, us03_n826, us03_n827, us03_n828, 
       us03_n829, us03_n830, us03_n831, us03_n832, us03_n833, us03_n834, us03_n835, us03_n836, us03_n837, 
       us03_n838, us03_n839, us03_n840, us03_n841, us03_n842, us03_n843, us03_n844, us03_n845, us03_n846, 
       us03_n847, us03_n848, us03_n849, us03_n850, us03_n851, us03_n852, us03_n853, us03_n854, us03_n855, 
       us03_n856, us03_n857, us03_n858, us03_n859, us03_n860, us03_n861, us03_n862, us03_n863, us03_n864, 
       us03_n865, us03_n866, us03_n867, us03_n868, us03_n869, us03_n870, us03_n871, us03_n872, us03_n873, 
       us03_n874, us20_n438, us20_n439, us20_n440, us20_n441, us20_n442, us20_n443, us20_n444, us20_n445, 
       us20_n446, us20_n447, us20_n448, us20_n449, us20_n450, us20_n451, us20_n452, us20_n453, us20_n454, 
       us20_n455, us20_n456, us20_n457, us20_n458, us20_n459, us20_n460, us20_n461, us20_n462, us20_n463, 
       us20_n464, us20_n465, us20_n466, us20_n467, us20_n468, us20_n469, us20_n470, us20_n471, us20_n472, 
       us20_n473, us20_n474, us20_n475, us20_n476, us20_n477, us20_n478, us20_n479, us20_n480, us20_n481, 
       us20_n482, us20_n483, us20_n484, us20_n485, us20_n486, us20_n487, us20_n488, us20_n489, us20_n490, 
       us20_n491, us20_n492, us20_n493, us20_n494, us20_n495, us20_n496, us20_n497, us20_n498, us20_n499, 
       us20_n500, us20_n501, us20_n502, us20_n503, us20_n504, us20_n505, us20_n506, us20_n507, us20_n508, 
       us20_n509, us20_n510, us20_n511, us20_n512, us20_n513, us20_n514, us20_n515, us20_n516, us20_n517, 
       us20_n518, us20_n519, us20_n520, us20_n521, us20_n522, us20_n523, us20_n524, us20_n525, us20_n526, 
       us20_n527, us20_n528, us20_n529, us20_n530, us20_n531, us20_n532, us20_n533, us20_n534, us20_n535, 
       us20_n536, us20_n537, us20_n538, us20_n539, us20_n540, us20_n541, us20_n542, us20_n543, us20_n544, 
       us20_n545, us20_n546, us20_n547, us20_n548, us20_n549, us20_n550, us20_n551, us20_n552, us20_n553, 
       us20_n554, us20_n555, us20_n556, us20_n557, us20_n558, us20_n559, us20_n560, us20_n561, us20_n562, 
       us20_n563, us20_n564, us20_n565, us20_n566, us20_n567, us20_n568, us20_n569, us20_n570, us20_n571, 
       us20_n572, us20_n573, us20_n574, us20_n575, us20_n576, us20_n577, us20_n578, us20_n579, us20_n580, 
       us20_n581, us20_n582, us20_n583, us20_n584, us20_n585, us20_n586, us20_n587, us20_n588, us20_n589, 
       us20_n590, us20_n591, us20_n592, us20_n593, us20_n594, us20_n595, us20_n596, us20_n597, us20_n598, 
       us20_n599, us20_n600, us20_n601, us20_n602, us20_n603, us20_n604, us20_n605, us20_n606, us20_n607, 
       us20_n608, us20_n609, us20_n610, us20_n611, us20_n612, us20_n613, us20_n614, us20_n615, us20_n616, 
       us20_n617, us20_n618, us20_n619, us20_n620, us20_n621, us20_n622, us20_n623, us20_n624, us20_n625, 
       us20_n626, us20_n627, us20_n628, us20_n629, us20_n630, us20_n631, us20_n632, us20_n633, us20_n634, 
       us20_n635, us20_n636, us20_n637, us20_n638, us20_n639, us20_n640, us20_n641, us20_n642, us20_n643, 
       us20_n644, us20_n645, us20_n646, us20_n647, us20_n648, us20_n649, us20_n650, us20_n651, us20_n652, 
       us20_n653, us20_n654, us20_n655, us20_n656, us20_n657, us20_n658, us20_n659, us20_n660, us20_n661, 
       us20_n662, us20_n663, us20_n664, us20_n665, us20_n666, us20_n667, us20_n668, us20_n669, us20_n670, 
       us20_n671, us20_n672, us20_n673, us20_n674, us20_n675, us20_n676, us20_n677, us20_n678, us20_n679, 
       us20_n680, us20_n681, us20_n682, us20_n683, us20_n684, us20_n685, us20_n686, us20_n687, us20_n688, 
       us20_n689, us20_n690, us20_n691, us20_n692, us20_n693, us20_n694, us20_n695, us20_n696, us20_n697, 
       us20_n698, us20_n699, us20_n700, us20_n701, us20_n702, us20_n703, us20_n704, us20_n705, us20_n706, 
       us20_n707, us20_n708, us20_n709, us20_n710, us20_n711, us20_n712, us20_n713, us20_n714, us20_n715, 
       us20_n716, us20_n717, us20_n718, us20_n719, us20_n720, us20_n721, us20_n722, us20_n723, us20_n724, 
       us20_n725, us20_n726, us20_n727, us20_n728, us20_n729, us20_n730, us20_n731, us20_n732, us20_n733, 
       us20_n734, us20_n735, us20_n736, us20_n737, us20_n738, us20_n739, us20_n740, us20_n741, us20_n742, 
       us20_n743, us20_n744, us20_n745, us20_n746, us20_n747, us20_n748, us20_n749, us20_n750, us20_n751, 
       us20_n752, us20_n753, us20_n754, us20_n755, us20_n756, us20_n757, us20_n758, us20_n759, us20_n760, 
       us20_n761, us20_n762, us20_n763, us20_n764, us20_n765, us20_n766, us20_n767, us20_n768, us20_n769, 
       us20_n770, us20_n771, us20_n772, us20_n773, us20_n774, us20_n775, us20_n776, us20_n777, us20_n778, 
       us20_n779, us20_n780, us20_n781, us20_n782, us20_n783, us20_n784, us20_n785, us20_n786, us20_n787, 
       us20_n788, us20_n789, us20_n790, us20_n791, us20_n792, us20_n793, us20_n794, us20_n795, us20_n796, 
       us20_n797, us20_n798, us20_n799, us20_n800, us20_n801, us20_n802, us20_n803, us20_n804, us20_n805, 
       us20_n806, us20_n807, us20_n808, us20_n809, us20_n810, us20_n811, us20_n812, us20_n813, us20_n814, 
       us20_n815, us20_n816, us20_n817, us20_n818, us20_n819, us20_n820, us20_n821, us20_n822, us20_n823, 
       us20_n824, us20_n825, us20_n826, us20_n827, us20_n828, us20_n829, us20_n830, us20_n831, us20_n832, 
       us20_n833, us20_n834, us20_n835, us20_n836, us20_n837, us20_n838, us20_n839, us20_n840, us20_n841, 
       us20_n842, us20_n843, us20_n844, us20_n845, us20_n846, us20_n847, us20_n848, us20_n849, us20_n850, 
       us20_n851, us20_n852, us20_n853, us20_n854, us20_n855, us20_n856, us20_n857, us20_n858, us20_n859, 
       us20_n860, us20_n861, us20_n862, us20_n863, us20_n864, us20_n865, us20_n866, us20_n867, us20_n868, 
       us20_n869, us20_n870, us20_n871, us20_n872, us20_n873, us20_n874, us20_n875, us20_n876, us23_n438, 
       us23_n439, us23_n440, us23_n441, us23_n442, us23_n443, us23_n444, us23_n445, us23_n446, us23_n447, 
       us23_n448, us23_n449, us23_n450, us23_n451, us23_n452, us23_n453, us23_n454, us23_n455, us23_n456, 
       us23_n457, us23_n458, us23_n459, us23_n460, us23_n461, us23_n462, us23_n463, us23_n464, us23_n465, 
       us23_n466, us23_n467, us23_n468, us23_n469, us23_n470, us23_n471, us23_n472, us23_n473, us23_n474, 
       us23_n475, us23_n476, us23_n477, us23_n478, us23_n479, us23_n480, us23_n481, us23_n482, us23_n483, 
       us23_n484, us23_n485, us23_n486, us23_n487, us23_n488, us23_n489, us23_n490, us23_n491, us23_n492, 
       us23_n493, us23_n494, us23_n495, us23_n496, us23_n497, us23_n498, us23_n499, us23_n500, us23_n501, 
       us23_n502, us23_n503, us23_n504, us23_n505, us23_n506, us23_n507, us23_n508, us23_n509, us23_n510, 
       us23_n511, us23_n512, us23_n513, us23_n514, us23_n515, us23_n516, us23_n517, us23_n518, us23_n519, 
       us23_n520, us23_n521, us23_n522, us23_n523, us23_n524, us23_n525, us23_n526, us23_n527, us23_n528, 
       us23_n529, us23_n530, us23_n531, us23_n532, us23_n533, us23_n534, us23_n535, us23_n536, us23_n537, 
       us23_n538, us23_n539, us23_n540, us23_n541, us23_n542, us23_n543, us23_n544, us23_n545, us23_n546, 
       us23_n547, us23_n548, us23_n549, us23_n550, us23_n551, us23_n552, us23_n553, us23_n554, us23_n555, 
       us23_n556, us23_n557, us23_n558, us23_n559, us23_n560, us23_n561, us23_n562, us23_n563, us23_n564, 
       us23_n565, us23_n566, us23_n567, us23_n568, us23_n569, us23_n570, us23_n571, us23_n572, us23_n573, 
       us23_n574, us23_n575, us23_n576, us23_n577, us23_n578, us23_n579, us23_n580, us23_n581, us23_n582, 
       us23_n583, us23_n584, us23_n585, us23_n586, us23_n587, us23_n588, us23_n589, us23_n590, us23_n591, 
       us23_n592, us23_n593, us23_n594, us23_n595, us23_n596, us23_n597, us23_n598, us23_n599, us23_n600, 
       us23_n601, us23_n602, us23_n603, us23_n604, us23_n605, us23_n606, us23_n607, us23_n608, us23_n609, 
       us23_n610, us23_n611, us23_n612, us23_n613, us23_n614, us23_n615, us23_n616, us23_n617, us23_n618, 
       us23_n619, us23_n620, us23_n621, us23_n622, us23_n623, us23_n624, us23_n625, us23_n626, us23_n627, 
       us23_n628, us23_n629, us23_n630, us23_n631, us23_n632, us23_n633, us23_n634, us23_n635, us23_n636, 
       us23_n637, us23_n638, us23_n639, us23_n640, us23_n641, us23_n642, us23_n643, us23_n644, us23_n645, 
       us23_n646, us23_n647, us23_n648, us23_n649, us23_n650, us23_n651, us23_n652, us23_n653, us23_n654, 
       us23_n655, us23_n656, us23_n657, us23_n658, us23_n659, us23_n660, us23_n661, us23_n662, us23_n663, 
       us23_n664, us23_n665, us23_n666, us23_n667, us23_n668, us23_n669, us23_n670, us23_n671, us23_n672, 
       us23_n673, us23_n674, us23_n675, us23_n676, us23_n677, us23_n678, us23_n679, us23_n680, us23_n681, 
       us23_n682, us23_n683, us23_n684, us23_n685, us23_n686, us23_n687, us23_n688, us23_n689, us23_n690, 
       us23_n691, us23_n692, us23_n693, us23_n694, us23_n695, us23_n696, us23_n697, us23_n698, us23_n699, 
       us23_n700, us23_n701, us23_n702, us23_n703, us23_n704, us23_n705, us23_n706, us23_n707, us23_n708, 
       us23_n709, us23_n710, us23_n711, us23_n712, us23_n713, us23_n714, us23_n715, us23_n716, us23_n717, 
       us23_n718, us23_n719, us23_n720, us23_n721, us23_n722, us23_n723, us23_n724, us23_n725, us23_n726, 
       us23_n727, us23_n728, us23_n729, us23_n730, us23_n731, us23_n732, us23_n733, us23_n734, us23_n735, 
       us23_n736, us23_n737, us23_n738, us23_n739, us23_n740, us23_n741, us23_n742, us23_n743, us23_n744, 
       us23_n745, us23_n746, us23_n747, us23_n748, us23_n749, us23_n750, us23_n751, us23_n752, us23_n753, 
       us23_n754, us23_n755, us23_n756, us23_n757, us23_n758, us23_n759, us23_n760, us23_n761, us23_n762, 
       us23_n763, us23_n764, us23_n765, us23_n766, us23_n767, us23_n768, us23_n769, us23_n770, us23_n771, 
       us23_n772, us23_n773, us23_n774, us23_n775, us23_n776, us23_n777, us23_n778, us23_n779, us23_n780, 
       us23_n781, us23_n782, us23_n783, us23_n784, us23_n785, us23_n786, us23_n787, us23_n788, us23_n789, 
       us23_n790, us23_n791, us23_n792, us23_n793, us23_n794, us23_n795, us23_n796, us23_n797, us23_n798, 
       us23_n799, us23_n800, us23_n801, us23_n802, us23_n803, us23_n804, us23_n805, us23_n806, us23_n807, 
       us23_n808, us23_n809, us23_n810, us23_n811, us23_n812, us23_n813, us23_n814, us23_n815, us23_n816, 
       us23_n817, us23_n818, us23_n819, us23_n820, us23_n821, us23_n822, us23_n823, us23_n824, us23_n825, 
       us23_n826, us23_n827, us23_n828, us23_n829, us23_n830, us23_n831, us23_n832, us23_n833, us23_n834, 
       us23_n835, us23_n836, us23_n837, us23_n838, us23_n839, us23_n840, us23_n841, us23_n842, us23_n843, 
       us23_n844, us23_n845, us23_n846, us23_n847, us23_n848, us23_n849, us23_n850, us23_n851, us23_n852, 
       us23_n853, us23_n854, us23_n855, us23_n856, us23_n857, us23_n858, us23_n859, us23_n860, us23_n861, 
       us23_n862, us23_n863, us23_n864, us23_n865, us23_n866, us23_n867, us23_n868, us23_n869, us23_n870, 
       us23_n871, us23_n872, us23_n873, us23_n874, us23_n875, us30_n438, us30_n439, us30_n440, us30_n441, 
       us30_n442, us30_n443, us30_n444, us30_n445, us30_n446, us30_n447, us30_n448, us30_n449, us30_n450, 
       us30_n451, us30_n452, us30_n453, us30_n454, us30_n455, us30_n456, us30_n457, us30_n458, us30_n459, 
       us30_n460, us30_n461, us30_n462, us30_n463, us30_n464, us30_n465, us30_n466, us30_n467, us30_n468, 
       us30_n469, us30_n470, us30_n471, us30_n472, us30_n473, us30_n474, us30_n475, us30_n476, us30_n477, 
       us30_n478, us30_n479, us30_n480, us30_n481, us30_n482, us30_n483, us30_n484, us30_n485, us30_n486, 
       us30_n487, us30_n488, us30_n489, us30_n490, us30_n491, us30_n492, us30_n493, us30_n494, us30_n495, 
       us30_n496, us30_n497, us30_n498, us30_n499, us30_n500, us30_n501, us30_n502, us30_n503, us30_n504, 
       us30_n505, us30_n506, us30_n507, us30_n508, us30_n509, us30_n510, us30_n511, us30_n512, us30_n513, 
       us30_n514, us30_n515, us30_n516, us30_n517, us30_n518, us30_n519, us30_n520, us30_n521, us30_n522, 
       us30_n523, us30_n524, us30_n525, us30_n526, us30_n527, us30_n528, us30_n529, us30_n530, us30_n531, 
       us30_n532, us30_n533, us30_n534, us30_n535, us30_n536, us30_n537, us30_n538, us30_n539, us30_n540, 
       us30_n541, us30_n542, us30_n543, us30_n544, us30_n545, us30_n546, us30_n547, us30_n548, us30_n549, 
       us30_n550, us30_n551, us30_n552, us30_n553, us30_n554, us30_n555, us30_n556, us30_n557, us30_n558, 
       us30_n559, us30_n560, us30_n561, us30_n562, us30_n563, us30_n564, us30_n565, us30_n566, us30_n567, 
       us30_n568, us30_n569, us30_n570, us30_n571, us30_n572, us30_n573, us30_n574, us30_n575, us30_n576, 
       us30_n577, us30_n578, us30_n579, us30_n580, us30_n581, us30_n582, us30_n583, us30_n584, us30_n585, 
       us30_n586, us30_n587, us30_n588, us30_n589, us30_n590, us30_n591, us30_n592, us30_n593, us30_n594, 
       us30_n595, us30_n596, us30_n597, us30_n598, us30_n599, us30_n600, us30_n601, us30_n602, us30_n603, 
       us30_n604, us30_n605, us30_n606, us30_n607, us30_n608, us30_n609, us30_n610, us30_n611, us30_n612, 
       us30_n613, us30_n614, us30_n615, us30_n616, us30_n617, us30_n618, us30_n619, us30_n620, us30_n621, 
       us30_n622, us30_n623, us30_n624, us30_n625, us30_n626, us30_n627, us30_n628, us30_n629, us30_n630, 
       us30_n631, us30_n632, us30_n633, us30_n634, us30_n635, us30_n636, us30_n637, us30_n638, us30_n639, 
       us30_n640, us30_n641, us30_n642, us30_n643, us30_n644, us30_n645, us30_n646, us30_n647, us30_n648, 
       us30_n649, us30_n650, us30_n651, us30_n652, us30_n653, us30_n654, us30_n655, us30_n656, us30_n657, 
       us30_n658, us30_n659, us30_n660, us30_n661, us30_n662, us30_n663, us30_n664, us30_n665, us30_n666, 
       us30_n667, us30_n668, us30_n669, us30_n670, us30_n671, us30_n672, us30_n673, us30_n674, us30_n675, 
       us30_n676, us30_n677, us30_n678, us30_n679, us30_n680, us30_n681, us30_n682, us30_n683, us30_n684, 
       us30_n685, us30_n686, us30_n687, us30_n688, us30_n689, us30_n690, us30_n691, us30_n692, us30_n693, 
       us30_n694, us30_n695, us30_n696, us30_n697, us30_n698, us30_n699, us30_n700, us30_n701, us30_n702, 
       us30_n703, us30_n704, us30_n705, us30_n706, us30_n707, us30_n708, us30_n709, us30_n710, us30_n711, 
       us30_n712, us30_n713, us30_n714, us30_n715, us30_n716, us30_n717, us30_n718, us30_n719, us30_n720, 
       us30_n721, us30_n722, us30_n723, us30_n724, us30_n725, us30_n726, us30_n727, us30_n728, us30_n729, 
       us30_n730, us30_n731, us30_n732, us30_n733, us30_n734, us30_n735, us30_n736, us30_n737, us30_n738, 
       us30_n739, us30_n740, us30_n741, us30_n742, us30_n743, us30_n744, us30_n745, us30_n746, us30_n747, 
       us30_n748, us30_n749, us30_n750, us30_n751, us30_n752, us30_n753, us30_n754, us30_n755, us30_n756, 
       us30_n757, us30_n758, us30_n759, us30_n760, us30_n761, us30_n762, us30_n763, us30_n764, us30_n765, 
       us30_n766, us30_n767, us30_n768, us30_n769, us30_n770, us30_n771, us30_n772, us30_n773, us30_n774, 
       us30_n775, us30_n776, us30_n777, us30_n778, us30_n779, us30_n780, us30_n781, us30_n782, us30_n783, 
       us30_n784, us30_n785, us30_n786, us30_n787, us30_n788, us30_n789, us30_n790, us30_n791, us30_n792, 
       us30_n793, us30_n794, us30_n795, us30_n796, us30_n797, us30_n798, us30_n799, us30_n800, us30_n801, 
       us30_n802, us30_n803, us30_n804, us30_n805, us30_n806, us30_n807, us30_n808, us30_n809, us30_n810, 
       us30_n811, us30_n812, us30_n813, us30_n814, us30_n815, us30_n816, us30_n817, us30_n818, us30_n819, 
       us30_n820, us30_n821, us30_n822, us30_n823, us30_n824, us30_n825, us30_n826, us30_n827, us30_n828, 
       us30_n829, us30_n830, us30_n831, us30_n832, us30_n833, us30_n834, us30_n835, us30_n836, us30_n837, 
       us30_n838, us30_n839, us30_n840, us30_n841, us30_n842, us30_n843, us30_n844, us30_n845, us30_n846, 
       us30_n847, us30_n848, us30_n849, us30_n850, us30_n851, us30_n852, us30_n853, us30_n854, us30_n855, 
       us30_n856, us30_n857, us30_n858, us30_n859, us30_n860, us30_n861, us30_n862, us30_n863, us30_n864, 
       us30_n865, us30_n866, us30_n867, us30_n868, us30_n869, us30_n870, us30_n871, us30_n872, us30_n873, 
       us30_n874, us30_n875,  us30_n876;
  NOR2_X1 u0_u2_U10 (.ZN( u0_u2_n714 ) , .A2( u0_u2_n783 ) , .A1( u0_u2_n807 ) );
  OR4_X1 u0_u2_U100 (.ZN( u0_u2_n473 ) , .A4( u0_u2_n525 ) , .A3( u0_u2_n536 ) , .A2( u0_u2_n585 ) , .A1( u0_u2_n719 ) );
  NOR4_X1 u0_u2_U101 (.A4( u0_u2_n584 ) , .A3( u0_u2_n585 ) , .A2( u0_u2_n586 ) , .ZN( u0_u2_n593 ) , .A1( u0_u2_n690 ) );
  NOR4_X1 u0_u2_U102 (.A1( u0_u2_n591 ) , .ZN( u0_u2_n592 ) , .A3( u0_u2_n659 ) , .A2( u0_u2_n669 ) , .A4( u0_u2_n774 ) );
  OR4_X1 u0_u2_U103 (.ZN( u0_u2_n499 ) , .A4( u0_u2_n541 ) , .A2( u0_u2_n554 ) , .A1( u0_u2_n566 ) , .A3( u0_u2_n639 ) );
  OR3_X1 u0_u2_U104 (.A3( u0_u2_n513 ) , .A2( u0_u2_n514 ) , .A1( u0_u2_n515 ) , .ZN( u0_u2_n518 ) );
  AOI21_X1 u0_u2_U105 (.A( u0_u2_n677 ) , .B1( u0_u2_n678 ) , .ZN( u0_u2_n679 ) , .B2( u0_u2_n863 ) );
  INV_X1 u0_u2_U106 (.A( u0_u2_n761 ) , .ZN( u0_u2_n876 ) );
  OAI21_X1 u0_u2_U107 (.B1( u0_u2_n760 ) , .ZN( u0_u2_n761 ) , .A( u0_u2_n852 ) , .B2( u0_u2_n875 ) );
  AOI221_X1 u0_u2_U108 (.A( u0_u2_n720 ) , .B2( u0_u2_n721 ) , .ZN( u0_u2_n727 ) , .C1( u0_u2_n839 ) , .B1( u0_u2_n846 ) , .C2( u0_u2_n870 ) );
  OR2_X1 u0_u2_U109 (.A2( u0_u2_n718 ) , .A1( u0_u2_n719 ) , .ZN( u0_u2_n720 ) );
  INV_X1 u0_u2_U11 (.A( u0_u2_n785 ) , .ZN( u0_u2_n874 ) );
  INV_X1 u0_u2_U110 (.A( u0_u2_n470 ) , .ZN( u0_u2_n871 ) );
  OAI21_X1 u0_u2_U111 (.ZN( u0_u2_n470 ) , .B1( u0_u2_n816 ) , .A( u0_u2_n841 ) , .B2( u0_u2_n858 ) );
  NAND2_X1 u0_u2_U112 (.ZN( u0_u2_n439 ) , .A2( u0_u2_n850 ) , .A1( u0_u2_n868 ) );
  NAND2_X1 u0_u2_U113 (.ZN( u0_u2_n440 ) , .A2( u0_u2_n838 ) , .A1( u0_u2_n861 ) );
  AOI221_X1 u0_u2_U114 (.A( u0_u2_n771 ) , .ZN( u0_u2_n781 ) , .C2( u0_u2_n817 ) , .B2( u0_u2_n842 ) , .C1( u0_u2_n862 ) , .B1( u0_u2_n873 ) );
  INV_X1 u0_u2_U115 (.A( u0_u2_n768 ) , .ZN( u0_u2_n842 ) );
  NAND2_X1 u0_u2_U116 (.A1( u0_u2_n454 ) , .A2( u0_u2_n472 ) , .ZN( u0_u2_n756 ) );
  AOI211_X1 u0_u2_U117 (.B( u0_u2_n814 ) , .A( u0_u2_n815 ) , .ZN( u0_u2_n831 ) , .C1( u0_u2_n849 ) , .C2( u0_u2_n857 ) );
  AOI211_X1 u0_u2_U118 (.A( u0_u2_n595 ) , .ZN( u0_u2_n604 ) , .B( u0_u2_n628 ) , .C1( u0_u2_n852 ) , .C2( u0_u2_n862 ) );
  INV_X1 u0_u2_U119 (.A( u0_u2_n737 ) , .ZN( u0_u2_n846 ) );
  INV_X1 u0_u2_U12 (.A( u0_u2_n686 ) , .ZN( u0_u2_n879 ) );
  NAND2_X1 u0_u2_U120 (.A1( u0_u2_n458 ) , .A2( u0_u2_n460 ) , .ZN( u0_u2_n769 ) );
  NOR3_X1 u0_u2_U121 (.ZN( u0_u2_n497 ) , .A1( u0_u2_n789 ) , .A2( u0_u2_n857 ) , .A3( u0_u2_n870 ) );
  OAI22_X1 u0_u2_U122 (.B2( u0_u2_n757 ) , .B1( u0_u2_n758 ) , .A1( u0_u2_n759 ) , .ZN( u0_u2_n763 ) , .A2( u0_u2_n813 ) );
  NOR2_X1 u0_u2_U123 (.ZN( u0_u2_n758 ) , .A2( u0_u2_n859 ) , .A1( u0_u2_n867 ) );
  NOR3_X1 u0_u2_U124 (.ZN( u0_u2_n759 ) , .A2( u0_u2_n860 ) , .A1( u0_u2_n870 ) , .A3( u0_u2_n872 ) );
  NOR2_X1 u0_u2_U125 (.ZN( u0_u2_n539 ) , .A2( u0_u2_n756 ) , .A1( u0_u2_n757 ) );
  NOR2_X1 u0_u2_U126 (.ZN( u0_u2_n577 ) , .A1( u0_u2_n735 ) , .A2( u0_u2_n813 ) );
  OAI21_X1 u0_u2_U127 (.ZN( u0_u2_n794 ) , .A( u0_u2_n846 ) , .B1( u0_u2_n870 ) , .B2( u0_u2_n880 ) );
  NOR2_X1 u0_u2_U128 (.A2( u0_u2_n715 ) , .A1( u0_u2_n757 ) , .ZN( u0_u2_n778 ) );
  NOR2_X1 u0_u2_U129 (.ZN( u0_u2_n516 ) , .A1( u0_u2_n736 ) , .A2( u0_u2_n786 ) );
  INV_X1 u0_u2_U13 (.A( u0_u2_n687 ) , .ZN( u0_u2_n847 ) );
  NOR2_X1 u0_u2_U130 (.ZN( u0_u2_n553 ) , .A2( u0_u2_n787 ) , .A1( u0_u2_n821 ) );
  NOR2_X1 u0_u2_U131 (.ZN( u0_u2_n618 ) , .A2( u0_u2_n787 ) , .A1( u0_u2_n813 ) );
  NOR2_X1 u0_u2_U132 (.ZN( u0_u2_n514 ) , .A1( u0_u2_n819 ) , .A2( u0_u2_n824 ) );
  NOR2_X1 u0_u2_U133 (.A2( u0_u2_n715 ) , .A1( u0_u2_n769 ) , .ZN( u0_u2_n801 ) );
  NOR2_X1 u0_u2_U134 (.ZN( u0_u2_n663 ) , .A1( u0_u2_n754 ) , .A2( u0_u2_n787 ) );
  NOR2_X1 u0_u2_U135 (.ZN( u0_u2_n513 ) , .A2( u0_u2_n735 ) , .A1( u0_u2_n769 ) );
  INV_X1 u0_u2_U136 (.A( u0_u2_n754 ) , .ZN( u0_u2_n841 ) );
  NOR2_X1 u0_u2_U137 (.ZN( u0_u2_n689 ) , .A2( u0_u2_n715 ) , .A1( u0_u2_n824 ) );
  INV_X1 u0_u2_U138 (.A( u0_u2_n735 ) , .ZN( u0_u2_n859 ) );
  AOI21_X1 u0_u2_U139 (.B1( u0_u2_n706 ) , .ZN( u0_u2_n707 ) , .A( u0_u2_n739 ) , .B2( u0_u2_n770 ) );
  AOI222_X1 u0_u2_U14 (.ZN( u0_u2_n570 ) , .B1( u0_u2_n837 ) , .C1( u0_u2_n848 ) , .A2( u0_u2_n850 ) , .A1( u0_u2_n861 ) , .B2( u0_u2_n870 ) , .C2( u0_u2_n880 ) );
  INV_X1 u0_u2_U140 (.A( u0_u2_n757 ) , .ZN( u0_u2_n849 ) );
  AOI21_X1 u0_u2_U141 (.ZN( u0_u2_n547 ) , .A( u0_u2_n770 ) , .B2( u0_u2_n786 ) , .B1( u0_u2_n824 ) );
  AOI21_X1 u0_u2_U142 (.ZN( u0_u2_n576 ) , .B1( u0_u2_n757 ) , .B2( u0_u2_n769 ) , .A( u0_u2_n787 ) );
  AOI21_X1 u0_u2_U143 (.B1( u0_u2_n693 ) , .ZN( u0_u2_n694 ) , .A( u0_u2_n735 ) , .B2( u0_u2_n768 ) );
  NOR2_X1 u0_u2_U144 (.ZN( u0_u2_n575 ) , .A1( u0_u2_n736 ) , .A2( u0_u2_n769 ) );
  NOR2_X1 u0_u2_U145 (.ZN( u0_u2_n536 ) , .A1( u0_u2_n715 ) , .A2( u0_u2_n786 ) );
  AOI21_X1 u0_u2_U146 (.ZN( u0_u2_n696 ) , .B2( u0_u2_n756 ) , .B1( u0_u2_n770 ) , .A( u0_u2_n813 ) );
  NOR2_X1 u0_u2_U147 (.ZN( u0_u2_n718 ) , .A1( u0_u2_n769 ) , .A2( u0_u2_n770 ) );
  INV_X1 u0_u2_U148 (.A( u0_u2_n787 ) , .ZN( u0_u2_n857 ) );
  NOR2_X1 u0_u2_U149 (.ZN( u0_u2_n621 ) , .A1( u0_u2_n769 ) , .A2( u0_u2_n819 ) );
  AOI222_X1 u0_u2_U15 (.ZN( u0_u2_n667 ) , .A2( u0_u2_n846 ) , .B1( u0_u2_n848 ) , .C2( u0_u2_n852 ) , .A1( u0_u2_n867 ) , .C1( u0_u2_n870 ) , .B2( u0_u2_n877 ) );
  AOI21_X1 u0_u2_U150 (.B1( u0_u2_n444 ) , .ZN( u0_u2_n634 ) , .A( u0_u2_n770 ) , .B2( u0_u2_n821 ) );
  INV_X1 u0_u2_U151 (.A( u0_u2_n736 ) , .ZN( u0_u2_n875 ) );
  NOR2_X1 u0_u2_U152 (.ZN( u0_u2_n527 ) , .A2( u0_u2_n715 ) , .A1( u0_u2_n821 ) );
  NOR2_X1 u0_u2_U153 (.ZN( u0_u2_n584 ) , .A2( u0_u2_n706 ) , .A1( u0_u2_n821 ) );
  INV_X1 u0_u2_U154 (.A( u0_u2_n706 ) , .ZN( u0_u2_n860 ) );
  OAI21_X1 u0_u2_U155 (.A( u0_u2_n705 ) , .ZN( u0_u2_n709 ) , .B2( u0_u2_n757 ) , .B1( u0_u2_n811 ) );
  OAI21_X1 u0_u2_U156 (.ZN( u0_u2_n705 ) , .B2( u0_u2_n840 ) , .B1( u0_u2_n845 ) , .A( u0_u2_n867 ) );
  INV_X1 u0_u2_U157 (.A( u0_u2_n770 ) , .ZN( u0_u2_n873 ) );
  NAND2_X1 u0_u2_U158 (.A1( u0_u2_n706 ) , .A2( u0_u2_n736 ) , .ZN( u0_u2_n789 ) );
  BUF_X1 u0_u2_U159 (.Z( u0_u2_n443 ) , .A( u0_u2_n822 ) );
  INV_X1 u0_u2_U16 (.A( u0_u2_n654 ) , .ZN( u0_u2_n877 ) );
  INV_X1 u0_u2_U160 (.A( u0_u2_n824 ) , .ZN( u0_u2_n851 ) );
  NAND2_X1 u0_u2_U161 (.ZN( u0_u2_n721 ) , .A1( u0_u2_n735 ) , .A2( u0_u2_n787 ) );
  BUF_X1 u0_u2_U162 (.Z( u0_u2_n442 ) , .A( u0_u2_n676 ) );
  BUF_X1 u0_u2_U163 (.Z( u0_u2_n441 ) , .A( u0_u2_n704 ) );
  OR4_X1 u0_u2_U164 (.A3( u0_u2_n587 ) , .A4( u0_u2_n588 ) , .A2( u0_u2_n589 ) , .A1( u0_u2_n590 ) , .ZN( u0_u2_n591 ) );
  OAI222_X1 u0_u2_U165 (.A2( u0_u2_n443 ) , .B2( u0_u2_n715 ) , .ZN( u0_u2_n716 ) , .C2( u0_u2_n731 ) , .B1( u0_u2_n754 ) , .A1( u0_u2_n813 ) , .C1( u0_u2_n821 ) );
  AOI221_X1 u0_u2_U166 (.A( u0_u2_n457 ) , .ZN( u0_u2_n466 ) , .C2( u0_u2_n760 ) , .B1( u0_u2_n839 ) , .C1( u0_u2_n849 ) , .B2( u0_u2_n868 ) );
  OAI221_X1 u0_u2_U167 (.A( u0_u2_n790 ) , .C2( u0_u2_n791 ) , .B2( u0_u2_n792 ) , .B1( u0_u2_n793 ) , .ZN( u0_u2_n803 ) , .C1( u0_u2_n820 ) );
  OAI221_X1 u0_u2_U168 (.A( u0_u2_n703 ) , .ZN( u0_u2_n710 ) , .C2( u0_u2_n791 ) , .C1( u0_u2_n792 ) , .B1( u0_u2_n793 ) , .B2( u0_u2_n813 ) );
  AOI22_X1 u0_u2_U169 (.ZN( u0_u2_n703 ) , .A1( u0_u2_n837 ) , .B2( u0_u2_n850 ) , .A2( u0_u2_n872 ) , .B1( u0_u2_n875 ) );
  NOR4_X1 u0_u2_U17 (.A4( u0_u2_n551 ) , .A3( u0_u2_n552 ) , .A2( u0_u2_n553 ) , .A1( u0_u2_n554 ) , .ZN( u0_u2_n555 ) );
  OAI221_X1 u0_u2_U170 (.A( u0_u2_n734 ) , .C2( u0_u2_n735 ) , .B2( u0_u2_n736 ) , .B1( u0_u2_n737 ) , .ZN( u0_u2_n744 ) , .C1( u0_u2_n824 ) );
  NAND2_X1 u0_u2_U171 (.A2( u0_u2_n467 ) , .A1( u0_u2_n472 ) , .ZN( u0_u2_n787 ) );
  NAND2_X1 u0_u2_U172 (.A2( u0_u2_n478 ) , .A1( u0_u2_n479 ) , .ZN( u0_u2_n824 ) );
  NAND2_X1 u0_u2_U173 (.A1( u0_u2_n456 ) , .A2( u0_u2_n467 ) , .ZN( u0_u2_n799 ) );
  NAND2_X1 u0_u2_U174 (.A2( u0_u2_n455 ) , .A1( u0_u2_n467 ) , .ZN( u0_u2_n735 ) );
  NAND2_X1 u0_u2_U175 (.A2( u0_u2_n456 ) , .A1( u0_u2_n459 ) , .ZN( u0_u2_n770 ) );
  NAND2_X1 u0_u2_U176 (.A2( u0_u2_n461 ) , .A1( u0_u2_n479 ) , .ZN( u0_u2_n786 ) );
  NAND2_X1 u0_u2_U177 (.A1( u0_u2_n448 ) , .A2( u0_u2_n467 ) , .ZN( u0_u2_n706 ) );
  NAND2_X1 u0_u2_U178 (.A1( u0_u2_n460 ) , .A2( u0_u2_n479 ) , .ZN( u0_u2_n792 ) );
  NAND2_X1 u0_u2_U179 (.A2( u0_u2_n455 ) , .A1( u0_u2_n459 ) , .ZN( u0_u2_n736 ) );
  NOR4_X1 u0_u2_U18 (.A4( u0_u2_n539 ) , .A3( u0_u2_n540 ) , .A2( u0_u2_n541 ) , .ZN( u0_u2_n542 ) , .A1( u0_u2_n827 ) );
  NAND2_X1 u0_u2_U180 (.A2( u0_u2_n471 ) , .A1( u0_u2_n472 ) , .ZN( u0_u2_n819 ) );
  NAND2_X1 u0_u2_U181 (.A1( u0_u2_n462 ) , .A2( u0_u2_n478 ) , .ZN( u0_u2_n810 ) );
  NAND2_X1 u0_u2_U182 (.A1( u0_u2_n458 ) , .A2( u0_u2_n478 ) , .ZN( u0_u2_n823 ) );
  NAND2_X1 u0_u2_U183 (.A2( u0_u2_n448 ) , .A1( u0_u2_n454 ) , .ZN( u0_u2_n791 ) );
  NAND2_X1 u0_u2_U184 (.A1( u0_u2_n461 ) , .A2( u0_u2_n468 ) , .ZN( u0_u2_n820 ) );
  NOR2_X1 u0_u2_U185 (.ZN( u0_u2_n460 ) , .A1( u0_u2_n833 ) , .A2( u0_u2_n834 ) );
  NAND2_X1 u0_u2_U186 (.A2( u0_u2_n468 ) , .A1( u0_u2_n469 ) , .ZN( u0_u2_n754 ) );
  NAND2_X1 u0_u2_U187 (.A1( u0_u2_n454 ) , .A2( u0_u2_n455 ) , .ZN( u0_u2_n793 ) );
  NAND2_X1 u0_u2_U188 (.A1( u0_u2_n448 ) , .A2( u0_u2_n471 ) , .ZN( u0_u2_n715 ) );
  NAND2_X1 u0_u2_U189 (.A1( u0_u2_n469 ) , .A2( u0_u2_n479 ) , .ZN( u0_u2_n795 ) );
  NOR4_X1 u0_u2_U19 (.A4( u0_u2_n452 ) , .A3( u0_u2_n453 ) , .A2( u0_u2_n523 ) , .A1( u0_u2_n548 ) , .ZN( u0_u2_n713 ) );
  NAND2_X1 u0_u2_U190 (.A2( u0_u2_n448 ) , .A1( u0_u2_n459 ) , .ZN( u0_u2_n798 ) );
  NAND2_X1 u0_u2_U191 (.A1( u0_u2_n458 ) , .A2( u0_u2_n469 ) , .ZN( u0_u2_n797 ) );
  NAND2_X1 u0_u2_U192 (.A2( u0_u2_n461 ) , .A1( u0_u2_n462 ) , .ZN( u0_u2_n737 ) );
  AOI222_X1 u0_u2_U193 (.B2( u0_u2_n645 ) , .ZN( u0_u2_n651 ) , .B1( u0_u2_n848 ) , .A1( u0_u2_n849 ) , .C2( u0_u2_n853 ) , .C1( u0_u2_n870 ) , .A2( u0_u2_n872 ) );
  NOR4_X1 u0_u2_U194 (.A4( u0_u2_n646 ) , .A3( u0_u2_n647 ) , .A2( u0_u2_n648 ) , .A1( u0_u2_n649 ) , .ZN( u0_u2_n650 ) );
  NAND4_X1 u0_u2_U195 (.ZN( u0_subword_8 ) , .A4( u0_u2_n508 ) , .A3( u0_u2_n509 ) , .A2( u0_u2_n510 ) , .A1( u0_u2_n511 ) );
  NOR4_X1 u0_u2_U196 (.A4( u0_u2_n505 ) , .A3( u0_u2_n506 ) , .A2( u0_u2_n507 ) , .ZN( u0_u2_n508 ) , .A1( u0_u2_n534 ) );
  AOI221_X1 u0_u2_U197 (.A( u0_u2_n504 ) , .ZN( u0_u2_n509 ) , .B2( u0_u2_n850 ) , .C1( u0_u2_n853 ) , .C2( u0_u2_n867 ) , .B1( u0_u2_n869 ) );
  AOI221_X1 u0_u2_U198 (.A( u0_u2_n788 ) , .ZN( u0_u2_n805 ) , .C2( u0_u2_n844 ) , .B2( u0_u2_n845 ) , .B1( u0_u2_n872 ) , .C1( u0_u2_n873 ) );
  NOR4_X1 u0_u2_U199 (.A4( u0_u2_n800 ) , .A3( u0_u2_n801 ) , .A2( u0_u2_n802 ) , .A1( u0_u2_n803 ) , .ZN( u0_u2_n804 ) );
  OR4_X1 u0_u2_U20 (.A4( u0_u2_n449 ) , .A2( u0_u2_n450 ) , .A1( u0_u2_n451 ) , .ZN( u0_u2_n452 ) , .A3( u0_u2_n560 ) );
  NOR4_X1 u0_u2_U200 (.A4( u0_u2_n707 ) , .A3( u0_u2_n708 ) , .A2( u0_u2_n709 ) , .A1( u0_u2_n710 ) , .ZN( u0_u2_n711 ) );
  AOI211_X1 u0_u2_U201 (.B( u0_u2_n701 ) , .A( u0_u2_n702 ) , .ZN( u0_u2_n712 ) , .C2( u0_u2_n838 ) , .C1( u0_u2_n858 ) );
  NAND4_X1 u0_u2_U202 (.ZN( u0_subword_15 ) , .A4( u0_u2_n829 ) , .A3( u0_u2_n830 ) , .A2( u0_u2_n831 ) , .A1( u0_u2_n832 ) );
  NOR4_X1 u0_u2_U203 (.A4( u0_u2_n825 ) , .A3( u0_u2_n826 ) , .A2( u0_u2_n827 ) , .A1( u0_u2_n828 ) , .ZN( u0_u2_n829 ) );
  NAND4_X1 u0_u2_U204 (.ZN( u0_subword_9 ) , .A4( u0_u2_n602 ) , .A3( u0_u2_n603 ) , .A2( u0_u2_n604 ) , .A1( u0_u2_n605 ) );
  NOR4_X1 u0_u2_U205 (.A4( u0_u2_n598 ) , .A3( u0_u2_n599 ) , .A2( u0_u2_n600 ) , .A1( u0_u2_n601 ) , .ZN( u0_u2_n602 ) );
  AOI211_X1 u0_u2_U206 (.B( u0_u2_n596 ) , .A( u0_u2_n597 ) , .ZN( u0_u2_n603 ) , .C2( u0_u2_n818 ) , .C1( u0_u2_n840 ) );
  NOR4_X1 u0_u2_U207 (.A3( u0_u2_n762 ) , .A2( u0_u2_n763 ) , .A1( u0_u2_n764 ) , .ZN( u0_u2_n765 ) , .A4( u0_u2_n876 ) );
  AOI211_X1 u0_u2_U208 (.B( u0_u2_n752 ) , .A( u0_u2_n753 ) , .ZN( u0_u2_n766 ) , .C1( u0_u2_n839 ) , .C2( u0_u2_n860 ) );
  NOR4_X1 u0_u2_U209 (.A4( u0_u2_n741 ) , .A3( u0_u2_n742 ) , .A2( u0_u2_n743 ) , .A1( u0_u2_n744 ) , .ZN( u0_u2_n745 ) );
  INV_X1 u0_u2_U21 (.A( u0_u2_n620 ) , .ZN( u0_u2_n882 ) );
  AOI211_X1 u0_u2_U210 (.B( u0_u2_n732 ) , .A( u0_u2_n733 ) , .ZN( u0_u2_n746 ) , .C1( u0_u2_n850 ) , .C2( u0_u2_n862 ) );
  AOI221_X1 u0_u2_U211 (.ZN( u0_u2_n475 ) , .C2( u0_u2_n721 ) , .B2( u0_u2_n838 ) , .C1( u0_u2_n852 ) , .B1( u0_u2_n867 ) , .A( u0_u2_n871 ) );
  AOI22_X1 u0_u2_U212 (.A2( u0_u2_n789 ) , .ZN( u0_u2_n790 ) , .B2( u0_u2_n838 ) , .A1( u0_u2_n841 ) , .B1( u0_u2_n870 ) );
  NAND2_X1 u0_u2_U213 (.A1( u0_u2_n460 ) , .A2( u0_u2_n468 ) , .ZN( u0_u2_n751 ) );
  NAND2_X1 u0_u2_U214 (.A1( u0_u2_n454 ) , .A2( u0_u2_n456 ) , .ZN( u0_u2_n812 ) );
  NAND2_X1 u0_u2_U215 (.A2( u0_u2_n460 ) , .A1( u0_u2_n462 ) , .ZN( u0_u2_n813 ) );
  NAND2_X1 u0_u2_U216 (.A1( u0_u2_n456 ) , .A2( u0_u2_n471 ) , .ZN( u0_u2_n731 ) );
  AOI21_X1 u0_u2_U217 (.ZN( u0_u2_n522 ) , .A( u0_u2_n736 ) , .B1( u0_u2_n757 ) , .B2( u0_u2_n810 ) );
  NOR2_X1 u0_u2_U218 (.ZN( u0_u2_n690 ) , .A2( u0_u2_n706 ) , .A1( u0_u2_n810 ) );
  NOR2_X1 u0_u2_U219 (.A1( u0_u2_n756 ) , .ZN( u0_u2_n774 ) , .A2( u0_u2_n810 ) );
  NOR4_X1 u0_u2_U22 (.ZN( u0_u2_n493 ) , .A1( u0_u2_n514 ) , .A2( u0_u2_n526 ) , .A4( u0_u2_n553 ) , .A3( u0_u2_n618 ) );
  NOR2_X1 u0_u2_U220 (.ZN( u0_u2_n524 ) , .A1( u0_u2_n715 ) , .A2( u0_u2_n810 ) );
  NOR2_X1 u0_u2_U221 (.ZN( u0_u2_n673 ) , .A1( u0_u2_n735 ) , .A2( u0_u2_n810 ) );
  NOR2_X1 u0_u2_U222 (.ZN( u0_u2_n608 ) , .A2( u0_u2_n787 ) , .A1( u0_u2_n810 ) );
  NAND2_X1 u0_u2_U223 (.A2( u0_u2_n468 ) , .A1( u0_u2_n478 ) , .ZN( u0_u2_n704 ) );
  NAND2_X1 u0_u2_U224 (.A1( u0_u2_n459 ) , .A2( u0_u2_n472 ) , .ZN( u0_u2_n676 ) );
  NAND2_X1 u0_u2_U225 (.A2( u0_u2_n455 ) , .A1( u0_u2_n471 ) , .ZN( u0_u2_n822 ) );
  NOR2_X1 u0_u2_U226 (.ZN( u0_u2_n458 ) , .A1( u0_u2_n835 ) , .A2( u0_u2_n836 ) );
  OR3_X1 u0_u2_U227 (.ZN( u0_u2_n453 ) , .A1( u0_u2_n535 ) , .A3( u0_u2_n584 ) , .A2( u0_u2_n882 ) );
  NAND2_X1 u0_u2_U228 (.A1( u0_u2_n458 ) , .A2( u0_u2_n461 ) , .ZN( u0_u2_n821 ) );
  AOI211_X1 u0_u2_U229 (.A( u0_u2_n503 ) , .ZN( u0_u2_n510 ) , .B( u0_u2_n809 ) , .C2( u0_u2_n846 ) , .C1( u0_u2_n858 ) );
  NOR4_X1 u0_u2_U23 (.ZN( u0_u2_n482 ) , .A1( u0_u2_n538 ) , .A3( u0_u2_n575 ) , .A4( u0_u2_n607 ) , .A2( u0_u2_n649 ) );
  NAND4_X1 u0_u2_U230 (.A4( u0_u2_n500 ) , .A3( u0_u2_n501 ) , .A1( u0_u2_n502 ) , .ZN( u0_u2_n809 ) , .A2( u0_u2_n874 ) );
  NOR4_X1 u0_u2_U231 (.A3( u0_u2_n445 ) , .A2( u0_u2_n498 ) , .A1( u0_u2_n499 ) , .ZN( u0_u2_n500 ) , .A4( u0_u2_n619 ) );
  OAI22_X1 u0_u2_U232 (.B1( u0_u2_n497 ) , .ZN( u0_u2_n498 ) , .A1( u0_u2_n693 ) , .A2( u0_u2_n770 ) , .B2( u0_u2_n824 ) );
  NOR2_X1 u0_u2_U233 (.ZN( u0_u2_n444 ) , .A2( u0_u2_n843 ) , .A1( u0_u2_n846 ) );
  NOR2_X1 u0_u2_U234 (.ZN( u0_u2_n632 ) , .A2( u0_u2_n843 ) , .A1( u0_u2_n846 ) );
  NOR2_X1 u0_u2_U235 (.ZN( u0_u2_n445 ) , .A2( u0_u2_n704 ) , .A1( u0_u2_n798 ) );
  OAI222_X1 u0_u2_U236 (.A2( u0_u2_n442 ) , .C1( u0_u2_n443 ) , .ZN( u0_u2_n681 ) , .B1( u0_u2_n754 ) , .B2( u0_u2_n791 ) , .C2( u0_u2_n795 ) , .A1( u0_u2_n824 ) );
  NOR4_X1 u0_u2_U237 (.A4( u0_u2_n491 ) , .ZN( u0_u2_n494 ) , .A1( u0_u2_n573 ) , .A2( u0_u2_n588 ) , .A3( u0_u2_n609 ) );
  AOI222_X1 u0_u2_U238 (.ZN( u0_u2_n613 ) , .A1( u0_u2_n837 ) , .C2( u0_u2_n844 ) , .B1( u0_u2_n849 ) , .A2( u0_u2_n863 ) , .B2( u0_u2_n868 ) , .C1( u0_u2_n875 ) );
  AOI222_X1 u0_u2_U239 (.ZN( u0_u2_n532 ) , .A1( u0_u2_n841 ) , .B2( u0_u2_n844 ) , .C1( u0_u2_n851 ) , .C2( u0_u2_n857 ) , .A2( u0_u2_n859 ) , .B1( u0_u2_n873 ) );
  INV_X1 u0_u2_U24 (.A( u0_u2_n756 ) , .ZN( u0_u2_n870 ) );
  NAND2_X1 u0_u2_U240 (.ZN( u0_u2_n620 ) , .A2( u0_u2_n844 ) , .A1( u0_u2_n880 ) );
  NAND4_X1 u0_u2_U241 (.A4( u0_u2_n486 ) , .A3( u0_u2_n487 ) , .A2( u0_u2_n488 ) , .A1( u0_u2_n489 ) , .ZN( u0_u2_n701 ) );
  NOR2_X1 u0_u2_U242 (.ZN( u0_u2_n586 ) , .A2( u0_u2_n715 ) , .A1( u0_u2_n737 ) );
  OAI21_X1 u0_u2_U243 (.A( u0_u2_n794 ) , .B2( u0_u2_n795 ) , .B1( u0_u2_n796 ) , .ZN( u0_u2_n802 ) );
  AOI21_X1 u0_u2_U244 (.ZN( u0_u2_n646 ) , .B2( u0_u2_n756 ) , .A( u0_u2_n795 ) , .B1( u0_u2_n819 ) );
  AOI21_X1 u0_u2_U245 (.ZN( u0_u2_n449 ) , .A( u0_u2_n706 ) , .B1( u0_u2_n740 ) , .B2( u0_u2_n757 ) );
  NOR2_X1 u0_u2_U246 (.ZN( u0_u2_n525 ) , .A1( u0_u2_n715 ) , .A2( u0_u2_n795 ) );
  INV_X1 u0_u2_U247 (.A( u0_u2_n795 ) , .ZN( u0_u2_n852 ) );
  NOR2_X1 u0_u2_U248 (.ZN( u0_u2_n456 ) , .A1( u0_u2_n855 ) , .A2( w3_4 ) );
  NOR2_X1 u0_u2_U249 (.ZN( u0_u2_n472 ) , .A2( u0_u2_n854 ) , .A1( u0_u2_n855 ) );
  NOR4_X1 u0_u2_U25 (.ZN( u0_u2_n486 ) , .A1( u0_u2_n527 ) , .A4( u0_u2_n564 ) , .A3( u0_u2_n589 ) , .A2( u0_u2_n637 ) );
  OAI222_X1 u0_u2_U250 (.B1( u0_u2_n441 ) , .ZN( u0_u2_n624 ) , .C1( u0_u2_n731 ) , .C2( u0_u2_n754 ) , .B2( u0_u2_n793 ) , .A2( u0_u2_n799 ) , .A1( u0_u2_n823 ) );
  NOR2_X1 u0_u2_U251 (.ZN( u0_u2_n467 ) , .A1( u0_u2_n856 ) , .A2( w3_7 ) );
  AOI21_X1 u0_u2_U252 (.ZN( u0_u2_n647 ) , .B2( u0_u2_n754 ) , .A( u0_u2_n799 ) , .B1( u0_u2_n810 ) );
  AOI21_X1 u0_u2_U253 (.A( u0_u2_n740 ) , .ZN( u0_u2_n741 ) , .B2( u0_u2_n787 ) , .B1( u0_u2_n799 ) );
  AOI21_X1 u0_u2_U254 (.ZN( u0_u2_n521 ) , .A( u0_u2_n786 ) , .B2( u0_u2_n799 ) , .B1( u0_u2_n819 ) );
  AOI21_X1 u0_u2_U255 (.B2( u0_u2_n770 ) , .ZN( u0_u2_n771 ) , .A( u0_u2_n795 ) , .B1( u0_u2_n799 ) );
  INV_X1 u0_u2_U256 (.A( u0_u2_n799 ) , .ZN( u0_u2_n858 ) );
  NOR2_X1 u0_u2_U257 (.ZN( u0_u2_n564 ) , .A1( u0_u2_n799 ) , .A2( u0_u2_n821 ) );
  NOR2_X1 u0_u2_U258 (.ZN( u0_u2_n590 ) , .A1( u0_u2_n799 ) , .A2( u0_u2_n824 ) );
  AOI221_X1 u0_u2_U259 (.A( u0_u2_n496 ) , .ZN( u0_u2_n501 ) , .B2( u0_u2_n843 ) , .C2( u0_u2_n848 ) , .C1( u0_u2_n858 ) , .B1( u0_u2_n867 ) );
  NOR3_X1 u0_u2_U26 (.ZN( u0_u2_n487 ) , .A2( u0_u2_n515 ) , .A3( u0_u2_n608 ) , .A1( u0_u2_n617 ) );
  NOR3_X1 u0_u2_U260 (.ZN( u0_u2_n447 ) , .A2( u0_u2_n843 ) , .A3( u0_u2_n844 ) , .A1( u0_u2_n853 ) );
  NOR4_X1 u0_u2_U261 (.A3( u0_u2_n680 ) , .A1( u0_u2_n681 ) , .ZN( u0_u2_n682 ) , .A4( u0_u2_n722 ) , .A2( u0_u2_n866 ) );
  INV_X1 u0_u2_U262 (.A( u0_u2_n679 ) , .ZN( u0_u2_n866 ) );
  NOR2_X1 u0_u2_U263 (.ZN( u0_u2_n478 ) , .A1( u0_u2_n833 ) , .A2( w3_1 ) );
  INV_X1 u0_u2_U264 (.ZN( u0_u2_n834 ) , .A( w3_1 ) );
  CLKBUF_X1 u0_u2_U265 (.Z( u0_u2_n446 ) , .A( u0_u2_n798 ) );
  NOR2_X1 u0_u2_U266 (.A2( u0_u2_n438 ) , .A1( u0_u2_n583 ) , .ZN( u0_u2_n594 ) );
  OAI22_X1 u0_u2_U267 (.B2( u0_u2_n786 ) , .B1( u0_u2_n787 ) , .ZN( u0_u2_n788 ) , .A2( u0_u2_n821 ) , .A1( u0_u2_n822 ) );
  AOI21_X1 u0_u2_U268 (.B1( u0_u2_n443 ) , .ZN( u0_u2_n596 ) , .B2( u0_u2_n706 ) , .A( u0_u2_n824 ) );
  INV_X1 u0_u2_U269 (.A( u0_u2_n822 ) , .ZN( u0_u2_n862 ) );
  AOI211_X1 u0_u2_U27 (.B( u0_u2_n484 ) , .A( u0_u2_n485 ) , .ZN( u0_u2_n489 ) , .C2( u0_u2_n840 ) , .C1( u0_u2_n868 ) );
  NOR2_X1 u0_u2_U270 (.ZN( u0_u2_n674 ) , .A1( u0_u2_n757 ) , .A2( u0_u2_n822 ) );
  NOR2_X1 u0_u2_U271 (.A1( u0_u2_n443 ) , .ZN( u0_u2_n477 ) , .A2( u0_u2_n786 ) );
  AOI21_X1 u0_u2_U272 (.B1( u0_u2_n443 ) , .ZN( u0_u2_n546 ) , .B2( u0_u2_n819 ) , .A( u0_u2_n821 ) );
  AOI21_X1 u0_u2_U273 (.B1( u0_u2_n443 ) , .ZN( u0_u2_n457 ) , .B2( u0_u2_n799 ) , .A( u0_u2_n810 ) );
  NOR2_X1 u0_u2_U274 (.A2( u0_u2_n443 ) , .ZN( u0_u2_n637 ) , .A1( u0_u2_n754 ) );
  INV_X1 u0_u2_U275 (.ZN( u0_u2_n865 ) , .A( w3_7 ) );
  AOI222_X1 u0_u2_U276 (.C2( u0_u2_n816 ) , .B2( u0_u2_n817 ) , .A2( u0_u2_n818 ) , .ZN( u0_u2_n830 ) , .C1( u0_u2_n839 ) , .A1( u0_u2_n846 ) , .B1( u0_u2_n860 ) );
  AOI22_X1 u0_u2_U277 (.ZN( u0_u2_n734 ) , .B1( u0_u2_n839 ) , .A2( u0_u2_n845 ) , .A1( u0_u2_n870 ) , .B2( u0_u2_n873 ) );
  AOI222_X1 u0_u2_U278 (.ZN( u0_u2_n476 ) , .B1( u0_u2_n839 ) , .A1( u0_u2_n846 ) , .C1( u0_u2_n849 ) , .C2( u0_u2_n858 ) , .A2( u0_u2_n862 ) , .B2( u0_u2_n872 ) );
  NOR2_X1 u0_u2_U279 (.A2( u0_u2_n443 ) , .ZN( u0_u2_n662 ) , .A1( u0_u2_n797 ) );
  NOR4_X1 u0_u2_U28 (.ZN( u0_u2_n488 ) , .A3( u0_u2_n539 ) , .A4( u0_u2_n552 ) , .A2( u0_u2_n574 ) , .A1( u0_u2_n724 ) );
  NOR2_X1 u0_u2_U280 (.ZN( u0_u2_n693 ) , .A1( u0_u2_n838 ) , .A2( u0_u2_n839 ) );
  NOR2_X1 u0_u2_U281 (.ZN( u0_u2_n528 ) , .A1( u0_u2_n797 ) , .A2( u0_u2_n819 ) );
  NOR2_X1 u0_u2_U282 (.ZN( u0_u2_n740 ) , .A2( u0_u2_n839 ) , .A1( u0_u2_n852 ) );
  NOR2_X1 u0_u2_U283 (.ZN( u0_u2_n668 ) , .A1( u0_u2_n736 ) , .A2( u0_u2_n797 ) );
  NOR2_X1 u0_u2_U284 (.ZN( u0_u2_n675 ) , .A2( u0_u2_n715 ) , .A1( u0_u2_n797 ) );
  INV_X1 u0_u2_U285 (.A( u0_u2_n797 ) , .ZN( u0_u2_n839 ) );
  NOR2_X1 u0_u2_U286 (.ZN( u0_u2_n468 ) , .A1( u0_u2_n836 ) , .A2( w3_2 ) );
  INV_X1 u0_u2_U287 (.ZN( u0_u2_n835 ) , .A( w3_2 ) );
  AOI21_X1 u0_u2_U288 (.ZN( u0_u2_n600 ) , .B1( u0_u2_n757 ) , .A( u0_u2_n799 ) , .B2( u0_u2_n820 ) );
  AOI21_X1 u0_u2_U289 (.A( u0_u2_n819 ) , .B2( u0_u2_n820 ) , .B1( u0_u2_n821 ) , .ZN( u0_u2_n826 ) );
  NOR2_X1 u0_u2_U29 (.ZN( u0_u2_n687 ) , .A2( u0_u2_n841 ) , .A1( u0_u2_n846 ) );
  AOI21_X1 u0_u2_U290 (.ZN( u0_u2_n656 ) , .B1( u0_u2_n736 ) , .B2( u0_u2_n770 ) , .A( u0_u2_n820 ) );
  NOR2_X1 u0_u2_U291 (.A2( u0_u2_n820 ) , .A1( u0_u2_n822 ) , .ZN( u0_u2_n828 ) );
  NOR2_X1 u0_u2_U292 (.ZN( u0_u2_n585 ) , .A1( u0_u2_n715 ) , .A2( u0_u2_n820 ) );
  NOR2_X1 u0_u2_U293 (.ZN( u0_u2_n672 ) , .A1( u0_u2_n787 ) , .A2( u0_u2_n820 ) );
  NOR2_X1 u0_u2_U294 (.A1( u0_u2_n706 ) , .ZN( u0_u2_n775 ) , .A2( u0_u2_n820 ) );
  NOR2_X1 u0_u2_U295 (.ZN( u0_u2_n661 ) , .A1( u0_u2_n735 ) , .A2( u0_u2_n820 ) );
  INV_X1 u0_u2_U296 (.A( u0_u2_n820 ) , .ZN( u0_u2_n843 ) );
  AOI21_X1 u0_u2_U297 (.ZN( u0_u2_n598 ) , .B2( u0_u2_n770 ) , .A( u0_u2_n792 ) , .B1( u0_u2_n819 ) );
  AND2_X1 u0_u2_U298 (.ZN( u0_u2_n739 ) , .A1( u0_u2_n786 ) , .A2( u0_u2_n792 ) );
  NOR2_X1 u0_u2_U299 (.ZN( u0_u2_n670 ) , .A1( u0_u2_n736 ) , .A2( u0_u2_n792 ) );
  NAND2_X1 u0_u2_U3 (.ZN( u0_u2_n438 ) , .A1( u0_u2_n439 ) , .A2( u0_u2_n440 ) );
  NAND4_X1 u0_u2_U30 (.A4( u0_u2_n610 ) , .A3( u0_u2_n611 ) , .A2( u0_u2_n612 ) , .A1( u0_u2_n613 ) , .ZN( u0_u2_n729 ) );
  NOR2_X1 u0_u2_U300 (.ZN( u0_u2_n515 ) , .A2( u0_u2_n787 ) , .A1( u0_u2_n792 ) );
  NOR2_X1 u0_u2_U301 (.A2( u0_u2_n443 ) , .ZN( u0_u2_n622 ) , .A1( u0_u2_n792 ) );
  INV_X1 u0_u2_U302 (.A( u0_u2_n792 ) , .ZN( u0_u2_n853 ) );
  OAI22_X1 u0_u2_U303 (.ZN( u0_u2_n490 ) , .A1( u0_u2_n715 ) , .B2( u0_u2_n792 ) , .A2( u0_u2_n813 ) , .B1( u0_u2_n819 ) );
  NOR2_X1 u0_u2_U304 (.ZN( u0_u2_n636 ) , .A2( u0_u2_n735 ) , .A1( u0_u2_n792 ) );
  NOR2_X1 u0_u2_U305 (.ZN( u0_u2_n550 ) , .A2( u0_u2_n715 ) , .A1( u0_u2_n792 ) );
  NOR2_X1 u0_u2_U306 (.ZN( u0_u2_n551 ) , .A2( u0_u2_n792 ) , .A1( u0_u2_n799 ) );
  NAND4_X1 u0_u2_U307 (.A4( u0_u2_n698 ) , .A3( u0_u2_n699 ) , .A1( u0_u2_n700 ) , .ZN( u0_u2_n783 ) , .A2( u0_u2_n879 ) );
  NOR4_X1 u0_u2_U308 (.A4( u0_u2_n783 ) , .A3( u0_u2_n784 ) , .A1( u0_u2_n785 ) , .ZN( u0_u2_n806 ) , .A2( u0_u2_n808 ) );
  AOI211_X1 u0_u2_U309 (.A( u0_u2_n644 ) , .ZN( u0_u2_n652 ) , .B( u0_u2_n750 ) , .C2( u0_u2_n846 ) , .C1( u0_u2_n861 ) );
  NOR3_X1 u0_u2_U31 (.A1( u0_u2_n606 ) , .ZN( u0_u2_n611 ) , .A3( u0_u2_n670 ) , .A2( u0_u2_n777 ) );
  NOR3_X1 u0_u2_U310 (.A3( u0_u2_n748 ) , .A2( u0_u2_n749 ) , .A1( u0_u2_n750 ) , .ZN( u0_u2_n767 ) );
  NAND4_X1 u0_u2_U311 (.A4( u0_u2_n640 ) , .A3( u0_u2_n641 ) , .A2( u0_u2_n642 ) , .A1( u0_u2_n643 ) , .ZN( u0_u2_n750 ) );
  NOR3_X1 u0_u2_U312 (.A3( u0_u2_n628 ) , .A2( u0_u2_n629 ) , .ZN( u0_u2_n643 ) , .A1( u0_u2_n732 ) );
  NOR4_X1 u0_u2_U313 (.A4( u0_u2_n621 ) , .A3( u0_u2_n622 ) , .A2( u0_u2_n623 ) , .A1( u0_u2_n624 ) , .ZN( u0_u2_n625 ) );
  NOR2_X1 u0_u2_U314 (.ZN( u0_u2_n459 ) , .A1( u0_u2_n865 ) , .A2( w3_6 ) );
  NOR2_X1 u0_u2_U315 (.ZN( u0_u2_n454 ) , .A2( u0_u2_n856 ) , .A1( u0_u2_n865 ) );
  NOR2_X1 u0_u2_U316 (.ZN( u0_u2_n471 ) , .A2( w3_6 ) , .A1( w3_7 ) );
  INV_X1 u0_u2_U317 (.ZN( u0_u2_n856 ) , .A( w3_6 ) );
  AOI21_X1 u0_u2_U318 (.ZN( u0_u2_n505 ) , .A( u0_u2_n731 ) , .B2( u0_u2_n769 ) , .B1( u0_u2_n821 ) );
  OAI22_X1 u0_u2_U319 (.ZN( u0_u2_n496 ) , .A1( u0_u2_n731 ) , .B2( u0_u2_n735 ) , .B1( u0_u2_n737 ) , .A2( u0_u2_n786 ) );
  NOR4_X1 u0_u2_U32 (.A3( u0_u2_n607 ) , .A2( u0_u2_n608 ) , .A1( u0_u2_n609 ) , .ZN( u0_u2_n610 ) , .A4( u0_u2_n662 ) );
  NOR2_X1 u0_u2_U320 (.ZN( u0_u2_n719 ) , .A2( u0_u2_n731 ) , .A1( u0_u2_n797 ) );
  NOR2_X1 u0_u2_U321 (.ZN( u0_u2_n535 ) , .A2( u0_u2_n731 ) , .A1( u0_u2_n810 ) );
  NOR2_X1 u0_u2_U322 (.ZN( u0_u2_n616 ) , .A2( u0_u2_n731 ) , .A1( u0_u2_n824 ) );
  NOR2_X1 u0_u2_U323 (.ZN( u0_u2_n533 ) , .A1( u0_u2_n731 ) , .A2( u0_u2_n757 ) );
  NOR2_X1 u0_u2_U324 (.ZN( u0_u2_n541 ) , .A1( u0_u2_n731 ) , .A2( u0_u2_n795 ) );
  NOR2_X1 u0_u2_U325 (.ZN( u0_u2_n638 ) , .A1( u0_u2_n731 ) , .A2( u0_u2_n820 ) );
  NOR2_X1 u0_u2_U326 (.ZN( u0_u2_n540 ) , .A2( u0_u2_n731 ) , .A1( u0_u2_n737 ) );
  INV_X1 u0_u2_U327 (.A( u0_u2_n731 ) , .ZN( u0_u2_n863 ) );
  NOR2_X1 u0_u2_U328 (.ZN( u0_u2_n455 ) , .A1( u0_u2_n854 ) , .A2( w3_5 ) );
  NOR2_X1 u0_u2_U329 (.ZN( u0_u2_n448 ) , .A2( w3_4 ) , .A1( w3_5 ) );
  NOR4_X1 u0_u2_U33 (.A4( u0_u2_n694 ) , .A3( u0_u2_n695 ) , .A2( u0_u2_n696 ) , .A1( u0_u2_n697 ) , .ZN( u0_u2_n698 ) );
  INV_X1 u0_u2_U330 (.ZN( u0_u2_n855 ) , .A( w3_5 ) );
  AOI21_X1 u0_u2_U331 (.A( u0_u2_n446 ) , .ZN( u0_u2_n648 ) , .B1( u0_u2_n687 ) , .B2( u0_u2_n824 ) );
  AOI21_X1 u0_u2_U332 (.B2( u0_u2_n446 ) , .A( u0_u2_n797 ) , .B1( u0_u2_n799 ) , .ZN( u0_u2_n800 ) );
  OAI22_X1 u0_u2_U333 (.B1( u0_u2_n446 ) , .ZN( u0_u2_n702 ) , .A2( u0_u2_n737 ) , .A1( u0_u2_n787 ) , .B2( u0_u2_n824 ) );
  AOI21_X1 u0_u2_U334 (.B2( u0_u2_n446 ) , .ZN( u0_u2_n504 ) , .A( u0_u2_n786 ) , .B1( u0_u2_n811 ) );
  AOI21_X1 u0_u2_U335 (.B2( u0_u2_n446 ) , .ZN( u0_u2_n571 ) , .B1( u0_u2_n731 ) , .A( u0_u2_n786 ) );
  AOI21_X1 u0_u2_U336 (.ZN( u0_u2_n450 ) , .B1( u0_u2_n796 ) , .B2( u0_u2_n798 ) , .A( u0_u2_n821 ) );
  NOR2_X1 u0_u2_U337 (.ZN( u0_u2_n671 ) , .A1( u0_u2_n792 ) , .A2( u0_u2_n798 ) );
  NOR2_X1 u0_u2_U338 (.ZN( u0_u2_n562 ) , .A1( u0_u2_n757 ) , .A2( u0_u2_n798 ) );
  NOR2_X1 u0_u2_U339 (.ZN( u0_u2_n566 ) , .A2( u0_u2_n798 ) , .A1( u0_u2_n810 ) );
  AOI221_X1 u0_u2_U34 (.A( u0_u2_n688 ) , .ZN( u0_u2_n699 ) , .B2( u0_u2_n847 ) , .C1( u0_u2_n849 ) , .C2( u0_u2_n869 ) , .B1( u0_u2_n872 ) );
  NAND2_X2 u0_u2_U340 (.A1( u0_u2_n462 ) , .A2( u0_u2_n469 ) , .ZN( u0_u2_n757 ) );
  NOR2_X1 u0_u2_U341 (.ZN( u0_u2_n649 ) , .A2( u0_u2_n795 ) , .A1( u0_u2_n798 ) );
  NOR2_X1 u0_u2_U342 (.ZN( u0_u2_n691 ) , .A1( u0_u2_n798 ) , .A2( u0_u2_n820 ) );
  NOR2_X1 u0_u2_U343 (.ZN( u0_u2_n549 ) , .A1( u0_u2_n769 ) , .A2( u0_u2_n798 ) );
  INV_X1 u0_u2_U344 (.A( u0_u2_n798 ) , .ZN( u0_u2_n880 ) );
  AOI21_X1 u0_u2_U345 (.B2( u0_u2_n442 ) , .ZN( u0_u2_n517 ) , .A( u0_u2_n737 ) , .B1( u0_u2_n822 ) );
  AOI21_X1 u0_u2_U346 (.B1( u0_u2_n446 ) , .ZN( u0_u2_n633 ) , .B2( u0_u2_n676 ) , .A( u0_u2_n797 ) );
  INV_X1 u0_u2_U347 (.A( u0_u2_n676 ) , .ZN( u0_u2_n872 ) );
  NOR2_X1 u0_u2_U348 (.A1( u0_u2_n442 ) , .ZN( u0_u2_n773 ) , .A2( u0_u2_n820 ) );
  NOR2_X1 u0_u2_U349 (.A1( u0_u2_n442 ) , .ZN( u0_u2_n659 ) , .A2( u0_u2_n821 ) );
  NOR2_X1 u0_u2_U35 (.A1( u0_u2_n685 ) , .ZN( u0_u2_n700 ) , .A2( u0_u2_n814 ) );
  AOI21_X1 u0_u2_U350 (.A( u0_u2_n442 ) , .ZN( u0_u2_n484 ) , .B1( u0_u2_n757 ) , .B2( u0_u2_n813 ) );
  NOR2_X1 u0_u2_U351 (.A1( u0_u2_n442 ) , .ZN( u0_u2_n534 ) , .A2( u0_u2_n786 ) );
  NOR2_X1 u0_u2_U352 (.A1( u0_u2_n442 ) , .ZN( u0_u2_n609 ) , .A2( u0_u2_n810 ) );
  NOR2_X1 u0_u2_U353 (.A2( u0_u2_n442 ) , .ZN( u0_u2_n635 ) , .A1( u0_u2_n792 ) );
  NOR2_X1 u0_u2_U354 (.ZN( u0_u2_n588 ) , .A1( u0_u2_n676 ) , .A2( u0_u2_n795 ) );
  OAI22_X1 u0_u2_U355 (.ZN( u0_u2_n644 ) , .A1( u0_u2_n706 ) , .B2( u0_u2_n735 ) , .A2( u0_u2_n769 ) , .B1( u0_u2_n823 ) );
  AOI21_X1 u0_u2_U356 (.ZN( u0_u2_n506 ) , .B1( u0_u2_n687 ) , .A( u0_u2_n819 ) , .B2( u0_u2_n823 ) );
  OAI22_X1 u0_u2_U357 (.A1( u0_u2_n731 ) , .ZN( u0_u2_n733 ) , .B2( u0_u2_n757 ) , .B1( u0_u2_n819 ) , .A2( u0_u2_n823 ) );
  AOI21_X1 u0_u2_U358 (.A( u0_u2_n443 ) , .B2( u0_u2_n823 ) , .B1( u0_u2_n824 ) , .ZN( u0_u2_n825 ) );
  OAI22_X1 u0_u2_U359 (.B1( u0_u2_n442 ) , .A1( u0_u2_n443 ) , .ZN( u0_u2_n631 ) , .B2( u0_u2_n754 ) , .A2( u0_u2_n823 ) );
  NOR2_X1 u0_u2_U36 (.ZN( u0_u2_n552 ) , .A1( u0_u2_n756 ) , .A2( u0_u2_n821 ) );
  NOR2_X1 u0_u2_U360 (.ZN( u0_u2_n606 ) , .A2( u0_u2_n798 ) , .A1( u0_u2_n823 ) );
  NOR2_X1 u0_u2_U361 (.ZN( u0_u2_n538 ) , .A2( u0_u2_n787 ) , .A1( u0_u2_n823 ) );
  NOR2_X1 u0_u2_U362 (.ZN( u0_u2_n526 ) , .A2( u0_u2_n706 ) , .A1( u0_u2_n823 ) );
  NOR2_X1 u0_u2_U363 (.A1( u0_u2_n442 ) , .ZN( u0_u2_n695 ) , .A2( u0_u2_n823 ) );
  NOR2_X1 u0_u2_U364 (.ZN( u0_u2_n565 ) , .A1( u0_u2_n715 ) , .A2( u0_u2_n823 ) );
  NOR2_X1 u0_u2_U365 (.ZN( u0_u2_n692 ) , .A1( u0_u2_n736 ) , .A2( u0_u2_n823 ) );
  NAND2_X1 u0_u2_U366 (.ZN( u0_u2_n678 ) , .A1( u0_u2_n813 ) , .A2( u0_u2_n823 ) );
  NOR2_X1 u0_u2_U367 (.ZN( u0_u2_n469 ) , .A2( w3_0 ) , .A1( w3_1 ) );
  NOR2_X1 u0_u2_U368 (.ZN( u0_u2_n461 ) , .A1( u0_u2_n834 ) , .A2( w3_0 ) );
  INV_X1 u0_u2_U369 (.ZN( u0_u2_n833 ) , .A( w3_0 ) );
  NOR2_X1 u0_u2_U37 (.ZN( u0_u2_n502 ) , .A1( u0_u2_n685 ) , .A2( u0_u2_n701 ) );
  INV_X1 u0_u2_U370 (.A( u0_u2_n819 ) , .ZN( u0_u2_n861 ) );
  INV_X1 u0_u2_U371 (.A( u0_u2_n823 ) , .ZN( u0_u2_n838 ) );
  INV_X1 u0_u2_U372 (.A( u0_u2_n810 ) , .ZN( u0_u2_n850 ) );
  INV_X1 u0_u2_U373 (.ZN( u0_u2_n854 ) , .A( w3_4 ) );
  INV_X1 u0_u2_U374 (.A( u0_u2_n441 ) , .ZN( u0_u2_n845 ) );
  NOR2_X1 u0_u2_U375 (.A1( u0_u2_n704 ) , .ZN( u0_u2_n777 ) , .A2( u0_u2_n822 ) );
  AOI21_X1 u0_u2_U376 (.B2( u0_u2_n441 ) , .ZN( u0_u2_n578 ) , .B1( u0_u2_n813 ) , .A( u0_u2_n819 ) );
  NOR2_X1 u0_u2_U377 (.ZN( u0_u2_n639 ) , .A2( u0_u2_n704 ) , .A1( u0_u2_n731 ) );
  NOR2_X1 u0_u2_U378 (.A2( u0_u2_n441 ) , .A1( u0_u2_n787 ) , .ZN( u0_u2_n827 ) );
  AOI21_X1 u0_u2_U379 (.B2( u0_u2_n441 ) , .ZN( u0_u2_n485 ) , .A( u0_u2_n756 ) , .B1( u0_u2_n786 ) );
  INV_X1 u0_u2_U38 (.A( u0_u2_n821 ) , .ZN( u0_u2_n840 ) );
  NOR2_X1 u0_u2_U380 (.A2( u0_u2_n441 ) , .ZN( u0_u2_n573 ) , .A1( u0_u2_n770 ) );
  NOR2_X1 u0_u2_U381 (.ZN( u0_u2_n669 ) , .A2( u0_u2_n704 ) , .A1( u0_u2_n736 ) );
  NOR2_X1 u0_u2_U382 (.A2( u0_u2_n441 ) , .ZN( u0_u2_n723 ) , .A1( u0_u2_n799 ) );
  NOR2_X1 u0_u2_U383 (.A2( u0_u2_n441 ) , .ZN( u0_u2_n601 ) , .A1( u0_u2_n735 ) );
  NOR2_X1 u0_u2_U384 (.A2( u0_u2_n441 ) , .ZN( u0_u2_n548 ) , .A1( u0_u2_n706 ) );
  NOR2_X1 u0_u2_U385 (.ZN( u0_u2_n587 ) , .A2( u0_u2_n704 ) , .A1( u0_u2_n798 ) );
  NOR2_X1 u0_u2_U386 (.ZN( u0_u2_n479 ) , .A2( w3_2 ) , .A1( w3_3 ) );
  NOR2_X1 u0_u2_U387 (.ZN( u0_u2_n462 ) , .A1( u0_u2_n835 ) , .A2( w3_3 ) );
  INV_X1 u0_u2_U388 (.ZN( u0_u2_n836 ) , .A( w3_3 ) );
  AOI21_X1 u0_u2_U389 (.ZN( u0_u2_n583 ) , .B2( u0_u2_n731 ) , .B1( u0_u2_n755 ) , .A( u0_u2_n792 ) );
  NAND4_X1 u0_u2_U39 (.A4( u0_u2_n664 ) , .A3( u0_u2_n665 ) , .A2( u0_u2_n666 ) , .A1( u0_u2_n667 ) , .ZN( u0_u2_n807 ) );
  OAI222_X1 u0_u2_U390 (.B2( u0_u2_n754 ) , .B1( u0_u2_n755 ) , .A2( u0_u2_n756 ) , .ZN( u0_u2_n764 ) , .C2( u0_u2_n812 ) , .C1( u0_u2_n821 ) , .A1( u0_u2_n824 ) );
  OAI21_X1 u0_u2_U391 (.A( u0_u2_n738 ) , .B1( u0_u2_n739 ) , .ZN( u0_u2_n743 ) , .B2( u0_u2_n812 ) );
  OAI22_X1 u0_u2_U392 (.B2( u0_u2_n810 ) , .B1( u0_u2_n811 ) , .A2( u0_u2_n812 ) , .A1( u0_u2_n813 ) , .ZN( u0_u2_n815 ) );
  OAI222_X1 u0_u2_U393 (.C2( u0_u2_n444 ) , .ZN( u0_u2_n512 ) , .B2( u0_u2_n654 ) , .B1( u0_u2_n754 ) , .A2( u0_u2_n755 ) , .C1( u0_u2_n812 ) , .A1( u0_u2_n813 ) );
  AOI21_X1 u0_u2_U394 (.ZN( u0_u2_n657 ) , .A( u0_u2_n786 ) , .B1( u0_u2_n799 ) , .B2( u0_u2_n812 ) );
  INV_X1 u0_u2_U395 (.A( u0_u2_n812 ) , .ZN( u0_u2_n867 ) );
  NOR2_X1 u0_u2_U396 (.ZN( u0_u2_n742 ) , .A2( u0_u2_n810 ) , .A1( u0_u2_n812 ) );
  NOR2_X1 u0_u2_U397 (.ZN( u0_u2_n491 ) , .A1( u0_u2_n795 ) , .A2( u0_u2_n812 ) );
  NOR2_X1 u0_u2_U398 (.ZN( u0_u2_n574 ) , .A1( u0_u2_n754 ) , .A2( u0_u2_n812 ) );
  AOI21_X1 u0_u2_U399 (.A( u0_u2_n441 ) , .B1( u0_u2_n442 ) , .ZN( u0_u2_n559 ) , .B2( u0_u2_n812 ) );
  NOR3_X1 u0_u2_U4 (.A3( u0_u2_n807 ) , .A2( u0_u2_n808 ) , .A1( u0_u2_n809 ) , .ZN( u0_u2_n832 ) );
  NOR3_X1 u0_u2_U40 (.A3( u0_u2_n661 ) , .A2( u0_u2_n662 ) , .A1( u0_u2_n663 ) , .ZN( u0_u2_n664 ) );
  NAND2_X1 u0_u2_U400 (.ZN( u0_u2_n760 ) , .A1( u0_u2_n770 ) , .A2( u0_u2_n812 ) );
  NOR2_X1 u0_u2_U401 (.ZN( u0_u2_n722 ) , .A1( u0_u2_n812 ) , .A2( u0_u2_n824 ) );
  NOR2_X1 u0_u2_U402 (.ZN( u0_u2_n563 ) , .A1( u0_u2_n769 ) , .A2( u0_u2_n812 ) );
  NOR2_X1 u0_u2_U403 (.ZN( u0_u2_n677 ) , .A1( u0_u2_n797 ) , .A2( u0_u2_n812 ) );
  NAND4_X1 u0_u2_U404 (.ZN( u0_subword_11 ) , .A4( u0_u2_n711 ) , .A3( u0_u2_n712 ) , .A2( u0_u2_n713 ) , .A1( u0_u2_n714 ) );
  INV_X1 u0_u2_U405 (.A( u0_u2_n713 ) , .ZN( u0_u2_n883 ) );
  OAI22_X1 u0_u2_U406 (.B2( u0_u2_n751 ) , .ZN( u0_u2_n753 ) , .A2( u0_u2_n769 ) , .B1( u0_u2_n787 ) , .A1( u0_u2_n799 ) );
  OAI22_X1 u0_u2_U407 (.B1( u0_u2_n446 ) , .ZN( u0_u2_n503 ) , .A2( u0_u2_n751 ) , .A1( u0_u2_n787 ) , .B2( u0_u2_n813 ) );
  NOR2_X1 u0_u2_U408 (.ZN( u0_u2_n523 ) , .A1( u0_u2_n715 ) , .A2( u0_u2_n751 ) );
  OAI22_X1 u0_u2_U409 (.ZN( u0_u2_n717 ) , .A2( u0_u2_n735 ) , .B2( u0_u2_n736 ) , .A1( u0_u2_n751 ) , .B1( u0_u2_n820 ) );
  NOR3_X1 u0_u2_U41 (.A3( u0_u2_n655 ) , .A2( u0_u2_n656 ) , .A1( u0_u2_n657 ) , .ZN( u0_u2_n666 ) );
  NOR2_X1 u0_u2_U410 (.A2( u0_u2_n751 ) , .ZN( u0_u2_n776 ) , .A1( u0_u2_n819 ) );
  OAI22_X1 u0_u2_U411 (.B1( u0_u2_n447 ) , .ZN( u0_u2_n451 ) , .A2( u0_u2_n735 ) , .A1( u0_u2_n751 ) , .B2( u0_u2_n756 ) );
  NOR2_X1 u0_u2_U412 (.ZN( u0_u2_n554 ) , .A1( u0_u2_n706 ) , .A2( u0_u2_n751 ) );
  NOR2_X1 u0_u2_U413 (.ZN( u0_u2_n537 ) , .A2( u0_u2_n751 ) , .A1( u0_u2_n799 ) );
  NOR2_X1 u0_u2_U414 (.A2( u0_u2_n751 ) , .ZN( u0_u2_n762 ) , .A1( u0_u2_n812 ) );
  NOR2_X1 u0_u2_U415 (.A1( u0_u2_n442 ) , .ZN( u0_u2_n680 ) , .A2( u0_u2_n751 ) );
  NOR2_X1 u0_u2_U416 (.ZN( u0_u2_n725 ) , .A2( u0_u2_n731 ) , .A1( u0_u2_n751 ) );
  NOR2_X1 u0_u2_U417 (.ZN( u0_u2_n589 ) , .A1( u0_u2_n751 ) , .A2( u0_u2_n822 ) );
  INV_X1 u0_u2_U418 (.A( u0_u2_n751 ) , .ZN( u0_u2_n844 ) );
  NAND4_X1 u0_u2_U419 (.ZN( u0_subword_10 ) , .A4( u0_u2_n650 ) , .A3( u0_u2_n651 ) , .A2( u0_u2_n652 ) , .A1( u0_u2_n653 ) );
  NOR3_X1 u0_u2_U42 (.A3( u0_u2_n658 ) , .A2( u0_u2_n659 ) , .A1( u0_u2_n660 ) , .ZN( u0_u2_n665 ) );
  OAI22_X1 u0_u2_U420 (.ZN( u0_u2_n595 ) , .A2( u0_u2_n754 ) , .B2( u0_u2_n769 ) , .A1( u0_u2_n770 ) , .B1( u0_u2_n791 ) );
  NAND2_X1 u0_u2_U421 (.A1( u0_u2_n736 ) , .A2( u0_u2_n791 ) , .ZN( u0_u2_n818 ) );
  AOI21_X1 u0_u2_U422 (.ZN( u0_u2_n599 ) , .B1( u0_u2_n735 ) , .B2( u0_u2_n791 ) , .A( u0_u2_n797 ) );
  AOI21_X1 u0_u2_U423 (.ZN( u0_u2_n655 ) , .A( u0_u2_n769 ) , .B2( u0_u2_n791 ) , .B1( u0_u2_n799 ) );
  AOI21_X1 u0_u2_U424 (.ZN( u0_u2_n630 ) , .B1( u0_u2_n706 ) , .A( u0_u2_n786 ) , .B2( u0_u2_n791 ) );
  OAI22_X1 u0_u2_U425 (.ZN( u0_u2_n688 ) , .A1( u0_u2_n706 ) , .A2( u0_u2_n737 ) , .B2( u0_u2_n791 ) , .B1( u0_u2_n824 ) );
  OAI21_X1 u0_u2_U426 (.A( u0_u2_n620 ) , .ZN( u0_u2_n623 ) , .B1( u0_u2_n632 ) , .B2( u0_u2_n791 ) );
  NOR2_X1 u0_u2_U427 (.ZN( u0_u2_n658 ) , .A1( u0_u2_n791 ) , .A2( u0_u2_n795 ) );
  NOR2_X1 u0_u2_U428 (.ZN( u0_u2_n617 ) , .A1( u0_u2_n791 ) , .A2( u0_u2_n823 ) );
  NOR2_X1 u0_u2_U429 (.ZN( u0_u2_n560 ) , .A2( u0_u2_n751 ) , .A1( u0_u2_n791 ) );
  NAND4_X1 u0_u2_U43 (.A4( u0_u2_n567 ) , .A3( u0_u2_n568 ) , .A2( u0_u2_n569 ) , .A1( u0_u2_n570 ) , .ZN( u0_u2_n614 ) );
  NOR2_X1 u0_u2_U430 (.A2( u0_u2_n441 ) , .ZN( u0_u2_n607 ) , .A1( u0_u2_n791 ) );
  INV_X1 u0_u2_U431 (.A( u0_u2_n791 ) , .ZN( u0_u2_n868 ) );
  AOI21_X1 u0_u2_U432 (.ZN( u0_u2_n507 ) , .A( u0_u2_n704 ) , .B1( u0_u2_n715 ) , .B2( u0_u2_n793 ) );
  OAI22_X1 u0_u2_U433 (.ZN( u0_u2_n597 ) , .B1( u0_u2_n737 ) , .B2( u0_u2_n756 ) , .A2( u0_u2_n793 ) , .A1( u0_u2_n810 ) );
  AOI222_X1 u0_u2_U434 (.ZN( u0_u2_n520 ) , .C1( u0_u2_n839 ) , .B2( u0_u2_n844 ) , .A2( u0_u2_n850 ) , .C2( u0_u2_n869 ) , .B1( u0_u2_n870 ) , .A1( u0_u2_n873 ) );
  AOI222_X1 u0_u2_U435 (.ZN( u0_u2_n612 ) , .B2( u0_u2_n678 ) , .B1( u0_u2_n760 ) , .C2( u0_u2_n838 ) , .A1( u0_u2_n840 ) , .A2( u0_u2_n869 ) , .C1( u0_u2_n870 ) );
  AOI221_X1 u0_u2_U436 (.A( u0_u2_n490 ) , .ZN( u0_u2_n495 ) , .B1( u0_u2_n838 ) , .C2( u0_u2_n851 ) , .C1( u0_u2_n859 ) , .B2( u0_u2_n869 ) );
  NAND3_X1 u0_u2_U437 (.ZN( u0_subword_14 ) , .A3( u0_u2_n804 ) , .A2( u0_u2_n805 ) , .A1( u0_u2_n806 ) );
  NAND3_X1 u0_u2_U438 (.ZN( u0_subword_13 ) , .A3( u0_u2_n765 ) , .A2( u0_u2_n766 ) , .A1( u0_u2_n767 ) );
  NAND3_X1 u0_u2_U439 (.ZN( u0_subword_12 ) , .A3( u0_u2_n745 ) , .A2( u0_u2_n746 ) , .A1( u0_u2_n747 ) );
  NOR4_X1 u0_u2_U44 (.ZN( u0_u2_n568 ) , .A1( u0_u2_n660 ) , .A3( u0_u2_n668 ) , .A4( u0_u2_n692 ) , .A2( u0_u2_n775 ) );
  NAND3_X1 u0_u2_U440 (.A3( u0_u2_n682 ) , .A2( u0_u2_n683 ) , .A1( u0_u2_n684 ) , .ZN( u0_u2_n814 ) );
  NAND3_X1 u0_u2_U441 (.ZN( u0_u2_n645 ) , .A3( u0_u2_n715 ) , .A2( u0_u2_n731 ) , .A1( u0_u2_n799 ) );
  NAND3_X1 u0_u2_U442 (.A3( u0_u2_n625 ) , .A2( u0_u2_n626 ) , .A1( u0_u2_n627 ) , .ZN( u0_u2_n732 ) );
  NAND3_X1 u0_u2_U443 (.A3( u0_u2_n592 ) , .A2( u0_u2_n593 ) , .A1( u0_u2_n594 ) , .ZN( u0_u2_n628 ) );
  NAND3_X1 u0_u2_U444 (.ZN( u0_u2_n572 ) , .A3( u0_u2_n687 ) , .A2( u0_u2_n757 ) , .A1( u0_u2_n792 ) );
  NAND3_X1 u0_u2_U445 (.A3( u0_u2_n530 ) , .A2( u0_u2_n531 ) , .A1( u0_u2_n532 ) , .ZN( u0_u2_n749 ) );
  NAND3_X1 u0_u2_U446 (.A3( u0_u2_n519 ) , .A1( u0_u2_n520 ) , .ZN( u0_u2_n615 ) , .A2( u0_u2_n878 ) );
  NAND3_X1 u0_u2_U447 (.A3( u0_u2_n474 ) , .A2( u0_u2_n475 ) , .A1( u0_u2_n476 ) , .ZN( u0_u2_n784 ) );
  NOR2_X1 u0_u2_U448 (.ZN( u0_u2_n660 ) , .A1( u0_u2_n769 ) , .A2( u0_u2_n793 ) );
  NAND2_X1 u0_u2_U449 (.A2( u0_u2_n756 ) , .A1( u0_u2_n793 ) , .ZN( u0_u2_n816 ) );
  NOR4_X1 u0_u2_U45 (.A4( u0_u2_n559 ) , .A3( u0_u2_n560 ) , .A2( u0_u2_n561 ) , .A1( u0_u2_n562 ) , .ZN( u0_u2_n569 ) );
  NOR2_X1 u0_u2_U450 (.ZN( u0_u2_n561 ) , .A1( u0_u2_n793 ) , .A2( u0_u2_n820 ) );
  NOR2_X1 u0_u2_U451 (.ZN( u0_u2_n619 ) , .A1( u0_u2_n786 ) , .A2( u0_u2_n793 ) );
  NOR2_X1 u0_u2_U452 (.ZN( u0_u2_n724 ) , .A2( u0_u2_n751 ) , .A1( u0_u2_n793 ) );
  NOR2_X1 u0_u2_U453 (.ZN( u0_u2_n796 ) , .A2( u0_u2_n869 ) , .A1( u0_u2_n875 ) );
  NOR2_X1 u0_u2_U454 (.ZN( u0_u2_n708 ) , .A2( u0_u2_n793 ) , .A1( u0_u2_n824 ) );
  NOR2_X1 u0_u2_U455 (.A1( u0_u2_n737 ) , .ZN( u0_u2_n772 ) , .A2( u0_u2_n793 ) );
  INV_X1 u0_u2_U456 (.A( u0_u2_n793 ) , .ZN( u0_u2_n869 ) );
  NOR4_X1 u0_u2_U46 (.A4( u0_u2_n563 ) , .A3( u0_u2_n564 ) , .A2( u0_u2_n565 ) , .A1( u0_u2_n566 ) , .ZN( u0_u2_n567 ) );
  NOR4_X1 u0_u2_U47 (.A4( u0_u2_n516 ) , .A2( u0_u2_n517 ) , .A1( u0_u2_n518 ) , .ZN( u0_u2_n519 ) , .A3( u0_u2_n677 ) );
  INV_X1 u0_u2_U48 (.A( u0_u2_n512 ) , .ZN( u0_u2_n878 ) );
  NOR4_X1 u0_u2_U49 (.A4( u0_u2_n668 ) , .A3( u0_u2_n669 ) , .A2( u0_u2_n670 ) , .A1( u0_u2_n671 ) , .ZN( u0_u2_n684 ) );
  NOR3_X1 u0_u2_U5 (.ZN( u0_u2_n605 ) , .A1( u0_u2_n615 ) , .A3( u0_u2_n730 ) , .A2( u0_u2_n749 ) );
  NOR4_X1 u0_u2_U50 (.A4( u0_u2_n672 ) , .A3( u0_u2_n673 ) , .A2( u0_u2_n674 ) , .A1( u0_u2_n675 ) , .ZN( u0_u2_n683 ) );
  NOR2_X1 u0_u2_U51 (.ZN( u0_u2_n811 ) , .A1( u0_u2_n861 ) , .A2( u0_u2_n868 ) );
  NOR4_X1 u0_u2_U52 (.A1( u0_u2_n473 ) , .ZN( u0_u2_n474 ) , .A4( u0_u2_n549 ) , .A2( u0_u2_n561 ) , .A3( u0_u2_n621 ) );
  NAND4_X1 u0_u2_U53 (.A4( u0_u2_n492 ) , .A3( u0_u2_n493 ) , .A2( u0_u2_n494 ) , .A1( u0_u2_n495 ) , .ZN( u0_u2_n785 ) );
  NOR4_X1 u0_u2_U54 (.ZN( u0_u2_n492 ) , .A2( u0_u2_n540 ) , .A1( u0_u2_n565 ) , .A3( u0_u2_n638 ) , .A4( u0_u2_n725 ) );
  NOR4_X1 u0_u2_U55 (.A4( u0_u2_n521 ) , .A3( u0_u2_n522 ) , .A2( u0_u2_n523 ) , .A1( u0_u2_n524 ) , .ZN( u0_u2_n531 ) );
  NOR4_X1 u0_u2_U56 (.A3( u0_u2_n528 ) , .A1( u0_u2_n529 ) , .ZN( u0_u2_n530 ) , .A2( u0_u2_n680 ) , .A4( u0_u2_n776 ) );
  NOR2_X1 u0_u2_U57 (.ZN( u0_u2_n768 ) , .A1( u0_u2_n840 ) , .A2( u0_u2_n841 ) );
  NAND4_X1 u0_u2_U58 (.A4( u0_u2_n779 ) , .A3( u0_u2_n780 ) , .A2( u0_u2_n781 ) , .A1( u0_u2_n782 ) , .ZN( u0_u2_n808 ) );
  NOR3_X1 u0_u2_U59 (.A3( u0_u2_n772 ) , .A2( u0_u2_n773 ) , .A1( u0_u2_n774 ) , .ZN( u0_u2_n780 ) );
  NOR3_X1 u0_u2_U6 (.ZN( u0_u2_n511 ) , .A2( u0_u2_n686 ) , .A3( u0_u2_n784 ) , .A1( u0_u2_n883 ) );
  NOR4_X1 u0_u2_U60 (.A4( u0_u2_n775 ) , .A3( u0_u2_n776 ) , .A2( u0_u2_n777 ) , .A1( u0_u2_n778 ) , .ZN( u0_u2_n779 ) );
  AOI222_X1 u0_u2_U61 (.ZN( u0_u2_n782 ) , .A1( u0_u2_n837 ) , .C1( u0_u2_n841 ) , .B2( u0_u2_n848 ) , .A2( u0_u2_n857 ) , .B1( u0_u2_n868 ) , .C2( u0_u2_n880 ) );
  NAND4_X1 u0_u2_U62 (.A4( u0_u2_n480 ) , .A3( u0_u2_n481 ) , .A2( u0_u2_n482 ) , .A1( u0_u2_n483 ) , .ZN( u0_u2_n685 ) );
  NOR4_X1 u0_u2_U63 (.A4( u0_u2_n477 ) , .ZN( u0_u2_n483 ) , .A3( u0_u2_n563 ) , .A1( u0_u2_n742 ) , .A2( u0_u2_n762 ) );
  NOR4_X1 u0_u2_U64 (.ZN( u0_u2_n480 ) , .A2( u0_u2_n528 ) , .A4( u0_u2_n601 ) , .A1( u0_u2_n616 ) , .A3( u0_u2_n636 ) );
  NOR4_X1 u0_u2_U65 (.ZN( u0_u2_n481 ) , .A1( u0_u2_n513 ) , .A3( u0_u2_n551 ) , .A2( u0_u2_n590 ) , .A4( u0_u2_n723 ) );
  NAND4_X1 u0_u2_U66 (.A4( u0_u2_n463 ) , .A3( u0_u2_n464 ) , .A2( u0_u2_n465 ) , .A1( u0_u2_n466 ) , .ZN( u0_u2_n686 ) );
  NOR3_X1 u0_u2_U67 (.ZN( u0_u2_n464 ) , .A3( u0_u2_n537 ) , .A1( u0_u2_n562 ) , .A2( u0_u2_n577 ) );
  NOR4_X1 u0_u2_U68 (.ZN( u0_u2_n463 ) , .A2( u0_u2_n524 ) , .A1( u0_u2_n550 ) , .A3( u0_u2_n586 ) , .A4( u0_u2_n622 ) );
  NOR4_X1 u0_u2_U69 (.ZN( u0_u2_n465 ) , .A2( u0_u2_n516 ) , .A1( u0_u2_n606 ) , .A4( u0_u2_n635 ) , .A3( u0_u2_n718 ) );
  NOR3_X1 u0_u2_U7 (.A2( u0_u2_n614 ) , .A1( u0_u2_n615 ) , .ZN( u0_u2_n653 ) , .A3( u0_u2_n729 ) );
  NAND4_X1 u0_u2_U70 (.A4( u0_u2_n580 ) , .A3( u0_u2_n581 ) , .A1( u0_u2_n582 ) , .ZN( u0_u2_n730 ) , .A2( u0_u2_n881 ) );
  NOR4_X1 u0_u2_U71 (.A4( u0_u2_n576 ) , .A3( u0_u2_n577 ) , .A2( u0_u2_n578 ) , .A1( u0_u2_n579 ) , .ZN( u0_u2_n580 ) );
  AOI221_X1 u0_u2_U72 (.A( u0_u2_n571 ) , .C2( u0_u2_n572 ) , .ZN( u0_u2_n581 ) , .B2( u0_u2_n852 ) , .B1( u0_u2_n859 ) , .C1( u0_u2_n860 ) );
  INV_X1 u0_u2_U73 (.A( u0_u2_n614 ) , .ZN( u0_u2_n881 ) );
  NOR4_X1 u0_u2_U74 (.A4( u0_u2_n636 ) , .A3( u0_u2_n637 ) , .A2( u0_u2_n638 ) , .A1( u0_u2_n639 ) , .ZN( u0_u2_n640 ) );
  AOI211_X1 u0_u2_U75 (.B( u0_u2_n630 ) , .A( u0_u2_n631 ) , .ZN( u0_u2_n642 ) , .C2( u0_u2_n843 ) , .C1( u0_u2_n870 ) );
  NOR4_X1 u0_u2_U76 (.A4( u0_u2_n633 ) , .A3( u0_u2_n634 ) , .A2( u0_u2_n635 ) , .ZN( u0_u2_n641 ) , .A1( u0_u2_n671 ) );
  NAND4_X1 u0_u2_U77 (.A4( u0_u2_n542 ) , .A3( u0_u2_n543 ) , .A2( u0_u2_n544 ) , .A1( u0_u2_n545 ) , .ZN( u0_u2_n629 ) );
  NOR4_X1 u0_u2_U78 (.A4( u0_u2_n533 ) , .A2( u0_u2_n534 ) , .A1( u0_u2_n535 ) , .ZN( u0_u2_n545 ) , .A3( u0_u2_n708 ) );
  NOR4_X1 u0_u2_U79 (.A1( u0_u2_n538 ) , .ZN( u0_u2_n543 ) , .A2( u0_u2_n661 ) , .A4( u0_u2_n675 ) , .A3( u0_u2_n772 ) );
  NOR3_X1 u0_u2_U8 (.A3( u0_u2_n729 ) , .A1( u0_u2_n730 ) , .ZN( u0_u2_n747 ) , .A2( u0_u2_n748 ) );
  NOR4_X1 u0_u2_U80 (.A4( u0_u2_n536 ) , .A3( u0_u2_n537 ) , .ZN( u0_u2_n544 ) , .A2( u0_u2_n691 ) , .A1( u0_u2_n801 ) );
  NOR2_X1 u0_u2_U81 (.ZN( u0_u2_n755 ) , .A1( u0_u2_n868 ) , .A2( u0_u2_n869 ) );
  NAND4_X1 u0_u2_U82 (.A4( u0_u2_n555 ) , .A3( u0_u2_n556 ) , .A2( u0_u2_n557 ) , .A1( u0_u2_n558 ) , .ZN( u0_u2_n752 ) );
  NOR3_X1 u0_u2_U83 (.ZN( u0_u2_n556 ) , .A2( u0_u2_n658 ) , .A1( u0_u2_n674 ) , .A3( u0_u2_n778 ) );
  AOI211_X1 u0_u2_U84 (.B( u0_u2_n546 ) , .A( u0_u2_n547 ) , .ZN( u0_u2_n558 ) , .C2( u0_u2_n846 ) , .C1( u0_u2_n858 ) );
  NOR4_X1 u0_u2_U85 (.A4( u0_u2_n548 ) , .A3( u0_u2_n549 ) , .A2( u0_u2_n550 ) , .ZN( u0_u2_n557 ) , .A1( u0_u2_n695 ) );
  NOR4_X1 u0_u2_U86 (.A4( u0_u2_n616 ) , .A3( u0_u2_n617 ) , .A2( u0_u2_n618 ) , .A1( u0_u2_n619 ) , .ZN( u0_u2_n626 ) );
  NOR4_X1 u0_u2_U87 (.ZN( u0_u2_n627 ) , .A1( u0_u2_n663 ) , .A3( u0_u2_n673 ) , .A4( u0_u2_n689 ) , .A2( u0_u2_n773 ) );
  NOR2_X1 u0_u2_U88 (.ZN( u0_u2_n654 ) , .A1( u0_u2_n861 ) , .A2( u0_u2_n875 ) );
  INV_X1 u0_u2_U89 (.A( u0_u2_n813 ) , .ZN( u0_u2_n848 ) );
  NOR2_X1 u0_u2_U9 (.ZN( u0_u2_n582 ) , .A1( u0_u2_n629 ) , .A2( u0_u2_n752 ) );
  NAND4_X1 u0_u2_U90 (.A4( u0_u2_n726 ) , .A3( u0_u2_n727 ) , .A2( u0_u2_n728 ) , .ZN( u0_u2_n748 ) , .A1( u0_u2_n864 ) );
  NOR4_X1 u0_u2_U91 (.A4( u0_u2_n722 ) , .A3( u0_u2_n723 ) , .A2( u0_u2_n724 ) , .A1( u0_u2_n725 ) , .ZN( u0_u2_n726 ) );
  AOI221_X1 u0_u2_U92 (.A( u0_u2_n717 ) , .ZN( u0_u2_n728 ) , .C2( u0_u2_n851 ) , .B2( u0_u2_n852 ) , .C1( u0_u2_n868 ) , .B1( u0_u2_n869 ) );
  INV_X1 u0_u2_U93 (.A( u0_u2_n716 ) , .ZN( u0_u2_n864 ) );
  INV_X1 u0_u2_U94 (.A( u0_u2_n769 ) , .ZN( u0_u2_n837 ) );
  NAND2_X1 u0_u2_U95 (.A2( u0_u2_n769 ) , .A1( u0_u2_n813 ) , .ZN( u0_u2_n817 ) );
  OAI21_X1 u0_u2_U96 (.ZN( u0_u2_n738 ) , .A( u0_u2_n840 ) , .B2( u0_u2_n859 ) , .B1( u0_u2_n880 ) );
  OR4_X1 u0_u2_U97 (.A4( u0_u2_n525 ) , .A2( u0_u2_n526 ) , .A1( u0_u2_n527 ) , .ZN( u0_u2_n529 ) , .A3( u0_u2_n828 ) );
  OR4_X1 u0_u2_U98 (.A4( u0_u2_n573 ) , .A3( u0_u2_n574 ) , .A2( u0_u2_n575 ) , .ZN( u0_u2_n579 ) , .A1( u0_u2_n672 ) );
  OR4_X1 u0_u2_U99 (.A4( u0_u2_n689 ) , .A3( u0_u2_n690 ) , .A2( u0_u2_n691 ) , .A1( u0_u2_n692 ) , .ZN( u0_u2_n697 ) );
  INV_X1 us03_U10 (.A( us03_n678 ) , .ZN( us03_n838 ) );
  NOR4_X1 us03_U100 (.A4( us03_n607 ) , .A3( us03_n608 ) , .A2( us03_n609 ) , .A1( us03_n610 ) , .ZN( us03_n617 ) );
  NOR4_X1 us03_U101 (.A4( us03_n612 ) , .A3( us03_n613 ) , .A2( us03_n614 ) , .A1( us03_n615 ) , .ZN( us03_n616 ) );
  NOR2_X1 us03_U102 (.ZN( us03_n684 ) , .A1( us03_n829 ) , .A2( us03_n830 ) );
  NAND4_X1 us03_U103 (.A4( us03_n471 ) , .A3( us03_n472 ) , .A2( us03_n473 ) , .A1( us03_n474 ) , .ZN( us03_n676 ) );
  NOR4_X1 us03_U104 (.A4( us03_n468 ) , .ZN( us03_n474 ) , .A3( us03_n554 ) , .A1( us03_n733 ) , .A2( us03_n753 ) );
  NOR4_X1 us03_U105 (.ZN( us03_n473 ) , .A1( us03_n529 ) , .A3( us03_n566 ) , .A4( us03_n598 ) , .A2( us03_n640 ) );
  NOR4_X1 us03_U106 (.ZN( us03_n472 ) , .A1( us03_n504 ) , .A3( us03_n542 ) , .A2( us03_n581 ) , .A4( us03_n714 ) );
  NAND4_X1 us03_U107 (.ZN( sa03_sr_1 ) , .A4( us03_n593 ) , .A3( us03_n594 ) , .A2( us03_n595 ) , .A1( us03_n596 ) );
  AOI211_X1 us03_U108 (.B( us03_n587 ) , .A( us03_n588 ) , .ZN( us03_n594 ) , .C2( us03_n809 ) , .C1( us03_n831 ) );
  NOR4_X1 us03_U109 (.A4( us03_n589 ) , .A3( us03_n590 ) , .A2( us03_n591 ) , .A1( us03_n592 ) , .ZN( us03_n593 ) );
  NOR4_X1 us03_U11 (.A4( us03_n443 ) , .A3( us03_n444 ) , .A2( us03_n514 ) , .A1( us03_n539 ) , .ZN( us03_n704 ) );
  AOI211_X1 us03_U110 (.A( us03_n586 ) , .ZN( us03_n595 ) , .B( us03_n619 ) , .C1( us03_n843 ) , .C2( us03_n853 ) );
  NAND4_X1 us03_U111 (.ZN( sa03_sr_0 ) , .A4( us03_n499 ) , .A3( us03_n500 ) , .A2( us03_n501 ) , .A1( us03_n502 ) );
  NOR4_X1 us03_U112 (.A4( us03_n496 ) , .A3( us03_n497 ) , .A2( us03_n498 ) , .ZN( us03_n499 ) , .A1( us03_n525 ) );
  AOI221_X1 us03_U113 (.A( us03_n495 ) , .ZN( us03_n500 ) , .B2( us03_n841 ) , .C1( us03_n844 ) , .C2( us03_n858 ) , .B1( us03_n860 ) );
  AOI211_X1 us03_U114 (.A( us03_n494 ) , .ZN( us03_n501 ) , .B( us03_n800 ) , .C2( us03_n837 ) , .C1( us03_n849 ) );
  NAND4_X1 us03_U115 (.A4( us03_n689 ) , .A3( us03_n690 ) , .A1( us03_n691 ) , .ZN( us03_n774 ) , .A2( us03_n870 ) );
  INV_X1 us03_U116 (.A( us03_n677 ) , .ZN( us03_n870 ) );
  AOI221_X1 us03_U117 (.A( us03_n679 ) , .ZN( us03_n690 ) , .B2( us03_n838 ) , .C1( us03_n840 ) , .C2( us03_n860 ) , .B1( us03_n863 ) );
  NOR4_X1 us03_U118 (.A4( us03_n685 ) , .A3( us03_n686 ) , .A2( us03_n687 ) , .A1( us03_n688 ) , .ZN( us03_n689 ) );
  NOR2_X1 us03_U119 (.ZN( us03_n731 ) , .A2( us03_n830 ) , .A1( us03_n843 ) );
  OR3_X1 us03_U12 (.ZN( us03_n444 ) , .A1( us03_n526 ) , .A3( us03_n575 ) , .A2( us03_n873 ) );
  NAND4_X1 us03_U120 (.A4( us03_n717 ) , .A3( us03_n718 ) , .A2( us03_n719 ) , .ZN( us03_n739 ) , .A1( us03_n855 ) );
  INV_X1 us03_U121 (.A( us03_n707 ) , .ZN( us03_n855 ) );
  NOR4_X1 us03_U122 (.A4( us03_n713 ) , .A3( us03_n714 ) , .A2( us03_n715 ) , .A1( us03_n716 ) , .ZN( us03_n717 ) );
  AOI221_X1 us03_U123 (.A( us03_n708 ) , .ZN( us03_n719 ) , .C2( us03_n842 ) , .B2( us03_n843 ) , .C1( us03_n859 ) , .B1( us03_n860 ) );
  NOR2_X1 us03_U124 (.ZN( us03_n645 ) , .A1( us03_n852 ) , .A2( us03_n866 ) );
  NAND4_X1 us03_U125 (.A4( us03_n571 ) , .A3( us03_n572 ) , .A1( us03_n573 ) , .ZN( us03_n721 ) , .A2( us03_n872 ) );
  NOR4_X1 us03_U126 (.A4( us03_n567 ) , .A3( us03_n568 ) , .A2( us03_n569 ) , .A1( us03_n570 ) , .ZN( us03_n571 ) );
  AOI221_X1 us03_U127 (.A( us03_n562 ) , .C2( us03_n563 ) , .ZN( us03_n572 ) , .B2( us03_n843 ) , .B1( us03_n850 ) , .C1( us03_n851 ) );
  INV_X1 us03_U128 (.A( us03_n605 ) , .ZN( us03_n872 ) );
  NAND4_X1 us03_U129 (.A4( us03_n491 ) , .A3( us03_n492 ) , .A1( us03_n493 ) , .ZN( us03_n800 ) , .A2( us03_n865 ) );
  OR4_X1 us03_U13 (.A4( us03_n440 ) , .A2( us03_n441 ) , .A1( us03_n442 ) , .ZN( us03_n443 ) , .A3( us03_n551 ) );
  AOI221_X1 us03_U130 (.A( us03_n487 ) , .ZN( us03_n492 ) , .B2( us03_n834 ) , .C2( us03_n839 ) , .C1( us03_n849 ) , .B1( us03_n858 ) );
  INV_X1 us03_U131 (.A( us03_n776 ) , .ZN( us03_n865 ) );
  NOR2_X1 us03_U132 (.ZN( us03_n493 ) , .A1( us03_n676 ) , .A2( us03_n692 ) );
  INV_X1 us03_U133 (.A( us03_n760 ) , .ZN( us03_n828 ) );
  INV_X1 us03_U134 (.A( us03_n461 ) , .ZN( us03_n862 ) );
  OAI21_X1 us03_U135 (.ZN( us03_n461 ) , .B1( us03_n807 ) , .A( us03_n832 ) , .B2( us03_n849 ) );
  OR4_X1 us03_U136 (.A4( us03_n578 ) , .A3( us03_n579 ) , .A2( us03_n580 ) , .A1( us03_n581 ) , .ZN( us03_n582 ) );
  OR4_X1 us03_U137 (.A4( us03_n564 ) , .A3( us03_n565 ) , .A2( us03_n566 ) , .ZN( us03_n570 ) , .A1( us03_n663 ) );
  OR4_X1 us03_U138 (.A4( us03_n516 ) , .A2( us03_n517 ) , .A1( us03_n518 ) , .ZN( us03_n520 ) , .A3( us03_n819 ) );
  OR4_X1 us03_U139 (.A4( us03_n680 ) , .A3( us03_n681 ) , .A2( us03_n682 ) , .A1( us03_n683 ) , .ZN( us03_n688 ) );
  INV_X1 us03_U14 (.A( us03_n611 ) , .ZN( us03_n873 ) );
  OR4_X1 us03_U140 (.ZN( us03_n464 ) , .A4( us03_n516 ) , .A3( us03_n527 ) , .A2( us03_n576 ) , .A1( us03_n710 ) );
  NAND2_X1 us03_U141 (.ZN( us03_n611 ) , .A2( us03_n835 ) , .A1( us03_n871 ) );
  OR3_X1 us03_U142 (.A3( us03_n504 ) , .A2( us03_n505 ) , .A1( us03_n506 ) , .ZN( us03_n509 ) );
  AOI221_X1 us03_U143 (.A( us03_n711 ) , .B2( us03_n712 ) , .ZN( us03_n718 ) , .C1( us03_n830 ) , .B1( us03_n837 ) , .C2( us03_n861 ) );
  OR2_X1 us03_U144 (.A2( us03_n709 ) , .A1( us03_n710 ) , .ZN( us03_n711 ) );
  INV_X1 us03_U145 (.A( us03_n752 ) , .ZN( us03_n867 ) );
  OAI21_X1 us03_U146 (.B1( us03_n751 ) , .ZN( us03_n752 ) , .A( us03_n843 ) , .B2( us03_n866 ) );
  INV_X1 us03_U147 (.A( us03_n670 ) , .ZN( us03_n857 ) );
  AOI21_X1 us03_U148 (.A( us03_n668 ) , .B1( us03_n669 ) , .ZN( us03_n670 ) , .B2( us03_n854 ) );
  AOI222_X1 us03_U149 (.ZN( us03_n658 ) , .A2( us03_n837 ) , .B1( us03_n839 ) , .C2( us03_n843 ) , .A1( us03_n858 ) , .C1( us03_n861 ) , .B2( us03_n868 ) );
  INV_X1 us03_U15 (.A( us03_n747 ) , .ZN( us03_n861 ) );
  INV_X1 us03_U150 (.A( us03_n645 ) , .ZN( us03_n868 ) );
  OAI22_X1 us03_U151 (.ZN( us03_n481 ) , .A1( us03_n706 ) , .B2( us03_n783 ) , .A2( us03_n804 ) , .B1( us03_n810 ) );
  NAND2_X1 us03_U152 (.A1( us03_n445 ) , .A2( us03_n463 ) , .ZN( us03_n747 ) );
  OAI222_X1 us03_U153 (.B2( us03_n745 ) , .B1( us03_n746 ) , .A2( us03_n747 ) , .ZN( us03_n755 ) , .C2( us03_n803 ) , .C1( us03_n812 ) , .A1( us03_n815 ) );
  OAI222_X1 us03_U154 (.B2( us03_n706 ) , .ZN( us03_n707 ) , .C2( us03_n722 ) , .B1( us03_n745 ) , .A1( us03_n804 ) , .C1( us03_n812 ) , .A2( us03_n813 ) );
  OAI222_X1 us03_U155 (.ZN( us03_n615 ) , .B1( us03_n695 ) , .C1( us03_n722 ) , .C2( us03_n745 ) , .B2( us03_n784 ) , .A2( us03_n790 ) , .A1( us03_n814 ) );
  OAI222_X1 us03_U156 (.ZN( us03_n503 ) , .C2( us03_n623 ) , .B2( us03_n645 ) , .B1( us03_n745 ) , .A2( us03_n746 ) , .C1( us03_n803 ) , .A1( us03_n804 ) );
  AOI22_X1 us03_U157 (.ZN( us03_n694 ) , .A1( us03_n828 ) , .B2( us03_n841 ) , .A2( us03_n863 ) , .B1( us03_n866 ) );
  INV_X1 us03_U158 (.A( us03_n728 ) , .ZN( us03_n837 ) );
  AOI221_X1 us03_U159 (.A( us03_n762 ) , .ZN( us03_n772 ) , .C2( us03_n808 ) , .B2( us03_n833 ) , .C1( us03_n853 ) , .B1( us03_n864 ) );
  AOI222_X1 us03_U16 (.ZN( us03_n561 ) , .B1( us03_n828 ) , .C1( us03_n839 ) , .A2( us03_n841 ) , .A1( us03_n852 ) , .B2( us03_n861 ) , .C2( us03_n871 ) );
  AOI21_X1 us03_U160 (.B2( us03_n761 ) , .ZN( us03_n762 ) , .A( us03_n786 ) , .B1( us03_n790 ) );
  INV_X1 us03_U161 (.A( us03_n759 ) , .ZN( us03_n833 ) );
  NAND2_X1 us03_U162 (.A1( us03_n449 ) , .A2( us03_n451 ) , .ZN( us03_n760 ) );
  INV_X1 us03_U163 (.A( us03_n788 ) , .ZN( us03_n830 ) );
  OAI22_X1 us03_U164 (.ZN( us03_n635 ) , .A1( us03_n697 ) , .B2( us03_n726 ) , .A2( us03_n760 ) , .B1( us03_n814 ) );
  OAI221_X1 us03_U165 (.A( us03_n725 ) , .C2( us03_n726 ) , .B2( us03_n727 ) , .B1( us03_n728 ) , .ZN( us03_n735 ) , .C1( us03_n815 ) );
  AOI22_X1 us03_U166 (.ZN( us03_n725 ) , .B1( us03_n830 ) , .A2( us03_n836 ) , .A1( us03_n861 ) , .B2( us03_n864 ) );
  OAI22_X1 us03_U167 (.ZN( us03_n487 ) , .A1( us03_n722 ) , .B2( us03_n726 ) , .B1( us03_n728 ) , .A2( us03_n777 ) );
  OAI22_X1 us03_U168 (.ZN( us03_n622 ) , .B1( us03_n667 ) , .B2( us03_n745 ) , .A1( us03_n813 ) , .A2( us03_n814 ) );
  OAI22_X1 us03_U169 (.A1( us03_n722 ) , .ZN( us03_n724 ) , .B2( us03_n748 ) , .B1( us03_n810 ) , .A2( us03_n814 ) );
  NOR4_X1 us03_U17 (.ZN( us03_n471 ) , .A2( us03_n519 ) , .A4( us03_n592 ) , .A1( us03_n607 ) , .A3( us03_n627 ) );
  OAI22_X1 us03_U170 (.B2( us03_n777 ) , .B1( us03_n778 ) , .ZN( us03_n779 ) , .A2( us03_n812 ) , .A1( us03_n813 ) );
  OAI22_X1 us03_U171 (.B2( us03_n742 ) , .ZN( us03_n744 ) , .A2( us03_n760 ) , .B1( us03_n778 ) , .A1( us03_n790 ) );
  OAI22_X1 us03_U172 (.B2( us03_n801 ) , .B1( us03_n802 ) , .A2( us03_n803 ) , .A1( us03_n804 ) , .ZN( us03_n806 ) );
  OAI22_X1 us03_U173 (.ZN( us03_n494 ) , .A2( us03_n742 ) , .A1( us03_n778 ) , .B1( us03_n789 ) , .B2( us03_n804 ) );
  INV_X1 us03_U174 (.A( us03_n742 ) , .ZN( us03_n835 ) );
  INV_X1 us03_U175 (.A( us03_n814 ) , .ZN( us03_n829 ) );
  INV_X1 us03_U176 (.A( us03_n786 ) , .ZN( us03_n843 ) );
  INV_X1 us03_U177 (.A( us03_n812 ) , .ZN( us03_n831 ) );
  OAI22_X1 us03_U178 (.ZN( us03_n588 ) , .B1( us03_n728 ) , .B2( us03_n747 ) , .A2( us03_n784 ) , .A1( us03_n801 ) );
  OAI22_X1 us03_U179 (.ZN( us03_n693 ) , .A2( us03_n728 ) , .A1( us03_n778 ) , .B1( us03_n789 ) , .B2( us03_n815 ) );
  NOR4_X1 us03_U18 (.ZN( us03_n477 ) , .A1( us03_n518 ) , .A4( us03_n555 ) , .A3( us03_n580 ) , .A2( us03_n628 ) );
  OAI22_X1 us03_U180 (.ZN( us03_n708 ) , .A2( us03_n726 ) , .B2( us03_n727 ) , .A1( us03_n742 ) , .B1( us03_n811 ) );
  INV_X1 us03_U181 (.A( us03_n667 ) , .ZN( us03_n863 ) );
  NOR2_X1 us03_U182 (.A1( us03_n695 ) , .ZN( us03_n768 ) , .A2( us03_n813 ) );
  NOR2_X1 us03_U183 (.ZN( us03_n664 ) , .A1( us03_n726 ) , .A2( us03_n801 ) );
  NOR2_X1 us03_U184 (.ZN( us03_n592 ) , .A2( us03_n695 ) , .A1( us03_n726 ) );
  NOR2_X1 us03_U185 (.ZN( us03_n568 ) , .A1( us03_n726 ) , .A2( us03_n804 ) );
  NOR2_X1 us03_U186 (.ZN( us03_n716 ) , .A2( us03_n722 ) , .A1( us03_n742 ) );
  NOR2_X1 us03_U187 (.ZN( us03_n544 ) , .A2( us03_n778 ) , .A1( us03_n812 ) );
  NOR2_X1 us03_U188 (.ZN( us03_n575 ) , .A2( us03_n697 ) , .A1( us03_n812 ) );
  NOR2_X1 us03_U189 (.ZN( us03_n652 ) , .A1( us03_n726 ) , .A2( us03_n811 ) );
  NOR4_X1 us03_U19 (.A4( us03_n530 ) , .A3( us03_n531 ) , .A2( us03_n532 ) , .ZN( us03_n533 ) , .A1( us03_n818 ) );
  NOR2_X1 us03_U190 (.ZN( us03_n610 ) , .A1( us03_n777 ) , .A2( us03_n784 ) );
  INV_X1 us03_U191 (.A( us03_n748 ) , .ZN( us03_n840 ) );
  NOR2_X1 us03_U192 (.ZN( us03_n530 ) , .A2( us03_n747 ) , .A1( us03_n748 ) );
  NOR2_X1 us03_U193 (.ZN( us03_n627 ) , .A2( us03_n726 ) , .A1( us03_n783 ) );
  NOR2_X1 us03_U194 (.ZN( us03_n613 ) , .A1( us03_n783 ) , .A2( us03_n813 ) );
  NOR2_X1 us03_U195 (.ZN( us03_n599 ) , .A2( us03_n778 ) , .A1( us03_n801 ) );
  NOR2_X1 us03_U196 (.ZN( us03_n609 ) , .A2( us03_n778 ) , .A1( us03_n804 ) );
  INV_X1 us03_U197 (.A( us03_n745 ) , .ZN( us03_n832 ) );
  NOR2_X1 us03_U198 (.A2( us03_n742 ) , .ZN( us03_n767 ) , .A1( us03_n810 ) );
  NOR2_X1 us03_U199 (.ZN( us03_n526 ) , .A2( us03_n722 ) , .A1( us03_n801 ) );
  NOR4_X1 us03_U20 (.ZN( us03_n454 ) , .A2( us03_n515 ) , .A1( us03_n541 ) , .A3( us03_n577 ) , .A4( us03_n613 ) );
  NOR2_X1 us03_U200 (.ZN( us03_n529 ) , .A2( us03_n778 ) , .A1( us03_n814 ) );
  NOR2_X1 us03_U201 (.ZN( us03_n626 ) , .A2( us03_n667 ) , .A1( us03_n783 ) );
  NOR2_X1 us03_U202 (.ZN( us03_n597 ) , .A2( us03_n789 ) , .A1( us03_n814 ) );
  INV_X1 us03_U203 (.A( us03_n790 ) , .ZN( us03_n849 ) );
  NOR2_X1 us03_U204 (.ZN( us03_n650 ) , .A1( us03_n667 ) , .A2( us03_n812 ) );
  NOR2_X1 us03_U205 (.A1( us03_n667 ) , .ZN( us03_n671 ) , .A2( us03_n742 ) );
  NOR2_X1 us03_U206 (.ZN( us03_n600 ) , .A1( us03_n667 ) , .A2( us03_n801 ) );
  NOR2_X1 us03_U207 (.A1( us03_n667 ) , .ZN( us03_n686 ) , .A2( us03_n814 ) );
  NOR2_X1 us03_U208 (.A2( us03_n706 ) , .A1( us03_n748 ) , .ZN( us03_n769 ) );
  NOR2_X1 us03_U209 (.A1( us03_n667 ) , .ZN( us03_n764 ) , .A2( us03_n811 ) );
  NOR4_X1 us03_U21 (.A4( us03_n539 ) , .A3( us03_n540 ) , .A2( us03_n541 ) , .ZN( us03_n548 ) , .A1( us03_n686 ) );
  NOR2_X1 us03_U210 (.A1( us03_n697 ) , .ZN( us03_n766 ) , .A2( us03_n811 ) );
  NOR2_X1 us03_U211 (.ZN( us03_n539 ) , .A2( us03_n695 ) , .A1( us03_n697 ) );
  NOR2_X1 us03_U212 (.ZN( us03_n525 ) , .A1( us03_n667 ) , .A2( us03_n777 ) );
  NOR2_X1 us03_U213 (.ZN( us03_n665 ) , .A1( us03_n748 ) , .A2( us03_n813 ) );
  NOR2_X1 us03_U214 (.ZN( us03_n553 ) , .A1( us03_n748 ) , .A2( us03_n789 ) );
  NOR2_X1 us03_U215 (.ZN( us03_n506 ) , .A2( us03_n778 ) , .A1( us03_n783 ) );
  NOR2_X1 us03_U216 (.ZN( us03_n541 ) , .A2( us03_n706 ) , .A1( us03_n783 ) );
  NOR2_X1 us03_U217 (.ZN( us03_n662 ) , .A1( us03_n783 ) , .A2( us03_n789 ) );
  NOR2_X1 us03_U218 (.A2( us03_n695 ) , .ZN( us03_n714 ) , .A1( us03_n790 ) );
  OAI22_X1 us03_U219 (.B1( us03_n438 ) , .ZN( us03_n442 ) , .A2( us03_n726 ) , .A1( us03_n742 ) , .B2( us03_n747 ) );
  NOR2_X1 us03_U22 (.ZN( us03_n678 ) , .A2( us03_n832 ) , .A1( us03_n837 ) );
  NOR3_X1 us03_U220 (.ZN( us03_n438 ) , .A2( us03_n834 ) , .A3( us03_n835 ) , .A1( us03_n844 ) );
  NOR2_X1 us03_U221 (.ZN( us03_n505 ) , .A1( us03_n810 ) , .A2( us03_n815 ) );
  INV_X1 us03_U222 (.A( us03_n804 ) , .ZN( us03_n839 ) );
  NOR2_X1 us03_U223 (.ZN( us03_n659 ) , .A1( us03_n727 ) , .A2( us03_n788 ) );
  NOR2_X1 us03_U224 (.ZN( us03_n660 ) , .A2( us03_n695 ) , .A1( us03_n727 ) );
  NOR2_X1 us03_U225 (.ZN( us03_n555 ) , .A1( us03_n790 ) , .A2( us03_n812 ) );
  NOR2_X1 us03_U226 (.ZN( us03_n543 ) , .A1( us03_n747 ) , .A2( us03_n812 ) );
  NOR2_X1 us03_U227 (.ZN( us03_n507 ) , .A1( us03_n727 ) , .A2( us03_n777 ) );
  INV_X1 us03_U228 (.A( us03_n801 ) , .ZN( us03_n841 ) );
  NOR2_X1 us03_U229 (.A2( us03_n695 ) , .A1( us03_n778 ) , .ZN( us03_n818 ) );
  NOR4_X1 us03_U23 (.A4( us03_n512 ) , .A3( us03_n513 ) , .A2( us03_n514 ) , .A1( us03_n515 ) , .ZN( us03_n522 ) );
  NOR2_X1 us03_U230 (.ZN( us03_n528 ) , .A2( us03_n742 ) , .A1( us03_n790 ) );
  OAI22_X1 us03_U231 (.B2( us03_n748 ) , .B1( us03_n749 ) , .A1( us03_n750 ) , .ZN( us03_n754 ) , .A2( us03_n804 ) );
  NOR2_X1 us03_U232 (.ZN( us03_n749 ) , .A2( us03_n850 ) , .A1( us03_n858 ) );
  NOR3_X1 us03_U233 (.ZN( us03_n750 ) , .A2( us03_n851 ) , .A1( us03_n861 ) , .A3( us03_n863 ) );
  NOR2_X1 us03_U234 (.A1( us03_n747 ) , .ZN( us03_n765 ) , .A2( us03_n801 ) );
  NOR2_X1 us03_U235 (.A2( us03_n742 ) , .ZN( us03_n753 ) , .A1( us03_n803 ) );
  NOR2_X1 us03_U236 (.ZN( us03_n542 ) , .A2( us03_n783 ) , .A1( us03_n790 ) );
  NOR2_X1 us03_U237 (.ZN( us03_n661 ) , .A1( us03_n727 ) , .A2( us03_n783 ) );
  INV_X1 us03_U238 (.A( us03_n726 ) , .ZN( us03_n850 ) );
  NOR2_X1 us03_U239 (.ZN( us03_n629 ) , .A1( us03_n722 ) , .A2( us03_n811 ) );
  AOI222_X1 us03_U24 (.ZN( us03_n523 ) , .A1( us03_n832 ) , .B2( us03_n835 ) , .C1( us03_n842 ) , .C2( us03_n848 ) , .A2( us03_n850 ) , .B1( us03_n864 ) );
  NOR2_X1 us03_U240 (.ZN( us03_n733 ) , .A2( us03_n801 ) , .A1( us03_n803 ) );
  NOR2_X1 us03_U241 (.ZN( us03_n612 ) , .A1( us03_n760 ) , .A2( us03_n810 ) );
  NOR4_X1 us03_U242 (.A2( us03_n489 ) , .A1( us03_n490 ) , .ZN( us03_n491 ) , .A3( us03_n578 ) , .A4( us03_n610 ) );
  OR4_X1 us03_U243 (.ZN( us03_n490 ) , .A4( us03_n532 ) , .A2( us03_n545 ) , .A1( us03_n557 ) , .A3( us03_n630 ) );
  OAI22_X1 us03_U244 (.B1( us03_n488 ) , .ZN( us03_n489 ) , .A1( us03_n684 ) , .A2( us03_n761 ) , .B2( us03_n815 ) );
  NOR3_X1 us03_U245 (.ZN( us03_n488 ) , .A1( us03_n780 ) , .A2( us03_n848 ) , .A3( us03_n861 ) );
  NOR2_X1 us03_U246 (.ZN( us03_n504 ) , .A2( us03_n726 ) , .A1( us03_n760 ) );
  NOR2_X1 us03_U247 (.ZN( us03_n514 ) , .A1( us03_n706 ) , .A2( us03_n742 ) );
  NOR2_X1 us03_U248 (.ZN( us03_n715 ) , .A2( us03_n742 ) , .A1( us03_n784 ) );
  NOR2_X1 us03_U249 (.ZN( us03_n552 ) , .A1( us03_n784 ) , .A2( us03_n811 ) );
  NOR4_X1 us03_U25 (.A3( us03_n519 ) , .A1( us03_n520 ) , .ZN( us03_n521 ) , .A2( us03_n671 ) , .A4( us03_n767 ) );
  NOR2_X1 us03_U250 (.ZN( us03_n515 ) , .A1( us03_n706 ) , .A2( us03_n801 ) );
  NOR2_X1 us03_U251 (.ZN( us03_n556 ) , .A1( us03_n706 ) , .A2( us03_n814 ) );
  NOR2_X1 us03_U252 (.ZN( us03_n519 ) , .A1( us03_n788 ) , .A2( us03_n810 ) );
  INV_X1 us03_U253 (.A( us03_n803 ) , .ZN( us03_n858 ) );
  NOR2_X1 us03_U254 (.ZN( us03_n628 ) , .A1( us03_n745 ) , .A2( us03_n813 ) );
  NOR2_X1 us03_U255 (.ZN( us03_n713 ) , .A1( us03_n803 ) , .A2( us03_n815 ) );
  AOI21_X1 us03_U256 (.ZN( us03_n569 ) , .B2( us03_n695 ) , .B1( us03_n804 ) , .A( us03_n810 ) );
  NOR2_X1 us03_U257 (.ZN( us03_n653 ) , .A1( us03_n788 ) , .A2( us03_n813 ) );
  NOR2_X1 us03_U258 (.ZN( us03_n666 ) , .A2( us03_n706 ) , .A1( us03_n788 ) );
  NOR2_X1 us03_U259 (.ZN( us03_n654 ) , .A1( us03_n745 ) , .A2( us03_n778 ) );
  AOI222_X1 us03_U26 (.B2( us03_n636 ) , .ZN( us03_n642 ) , .B1( us03_n839 ) , .A1( us03_n840 ) , .C2( us03_n844 ) , .C1( us03_n861 ) , .A2( us03_n863 ) );
  NOR2_X1 us03_U260 (.ZN( us03_n554 ) , .A1( us03_n760 ) , .A2( us03_n803 ) );
  NOR2_X1 us03_U261 (.ZN( us03_n540 ) , .A1( us03_n760 ) , .A2( us03_n789 ) );
  NOR2_X1 us03_U262 (.ZN( us03_n699 ) , .A2( us03_n784 ) , .A1( us03_n815 ) );
  NOR2_X1 us03_U263 (.ZN( us03_n607 ) , .A2( us03_n722 ) , .A1( us03_n815 ) );
  NOR2_X1 us03_U264 (.A1( us03_n728 ) , .ZN( us03_n763 ) , .A2( us03_n784 ) );
  AOI21_X1 us03_U265 (.A( us03_n813 ) , .B2( us03_n814 ) , .B1( us03_n815 ) , .ZN( us03_n816 ) );
  NOR2_X1 us03_U266 (.ZN( us03_n577 ) , .A2( us03_n706 ) , .A1( us03_n728 ) );
  NOR2_X1 us03_U267 (.ZN( us03_n531 ) , .A2( us03_n722 ) , .A1( us03_n728 ) );
  AOI21_X1 us03_U268 (.B1( us03_n623 ) , .ZN( us03_n625 ) , .A( us03_n761 ) , .B2( us03_n812 ) );
  AOI21_X1 us03_U269 (.A( us03_n810 ) , .B2( us03_n811 ) , .B1( us03_n812 ) , .ZN( us03_n817 ) );
  NOR4_X1 us03_U27 (.A4( us03_n637 ) , .A3( us03_n638 ) , .A2( us03_n639 ) , .A1( us03_n640 ) , .ZN( us03_n641 ) );
  AOI21_X1 us03_U270 (.ZN( us03_n513 ) , .A( us03_n727 ) , .B1( us03_n748 ) , .B2( us03_n801 ) );
  AOI21_X1 us03_U271 (.ZN( us03_n497 ) , .B1( us03_n678 ) , .A( us03_n810 ) , .B2( us03_n814 ) );
  AOI21_X1 us03_U272 (.ZN( us03_n476 ) , .B2( us03_n695 ) , .A( us03_n747 ) , .B1( us03_n777 ) );
  NOR2_X1 us03_U273 (.ZN( us03_n580 ) , .A1( us03_n742 ) , .A2( us03_n813 ) );
  NOR2_X1 us03_U274 (.ZN( us03_n640 ) , .A2( us03_n786 ) , .A1( us03_n789 ) );
  AOI21_X1 us03_U275 (.ZN( us03_n591 ) , .B1( us03_n748 ) , .A( us03_n790 ) , .B2( us03_n811 ) );
  NOR2_X1 us03_U276 (.A2( us03_n706 ) , .A1( us03_n760 ) , .ZN( us03_n792 ) );
  AOI21_X1 us03_U277 (.ZN( us03_n624 ) , .B2( us03_n667 ) , .A( us03_n788 ) , .B1( us03_n789 ) );
  NOR2_X1 us03_U278 (.ZN( us03_n668 ) , .A1( us03_n788 ) , .A2( us03_n803 ) );
  NOR2_X1 us03_U279 (.ZN( us03_n518 ) , .A2( us03_n706 ) , .A1( us03_n812 ) );
  NOR3_X1 us03_U28 (.A2( us03_n605 ) , .A1( us03_n606 ) , .ZN( us03_n644 ) , .A3( us03_n720 ) );
  AOI21_X1 us03_U280 (.ZN( us03_n475 ) , .A( us03_n667 ) , .B1( us03_n748 ) , .B2( us03_n804 ) );
  NOR2_X1 us03_U281 (.ZN( us03_n557 ) , .A2( us03_n789 ) , .A1( us03_n801 ) );
  NOR2_X1 us03_U282 (.ZN( us03_n517 ) , .A2( us03_n697 ) , .A1( us03_n814 ) );
  NOR2_X1 us03_U283 (.ZN( us03_n681 ) , .A2( us03_n697 ) , .A1( us03_n801 ) );
  NOR2_X1 us03_U284 (.ZN( us03_n651 ) , .A1( us03_n760 ) , .A2( us03_n784 ) );
  INV_X1 us03_U285 (.A( us03_n811 ) , .ZN( us03_n834 ) );
  AOI21_X1 us03_U286 (.ZN( us03_n508 ) , .B2( us03_n667 ) , .A( us03_n728 ) , .B1( us03_n813 ) );
  AOI21_X1 us03_U287 (.ZN( us03_n537 ) , .B2( us03_n810 ) , .A( us03_n812 ) , .B1( us03_n813 ) );
  INV_X1 us03_U288 (.A( us03_n761 ) , .ZN( us03_n864 ) );
  AOI21_X1 us03_U289 (.ZN( us03_n538 ) , .A( us03_n761 ) , .B2( us03_n777 ) , .B1( us03_n815 ) );
  AOI221_X1 us03_U29 (.A( us03_n779 ) , .ZN( us03_n796 ) , .C2( us03_n835 ) , .B2( us03_n836 ) , .B1( us03_n863 ) , .C1( us03_n864 ) );
  NOR2_X1 us03_U290 (.ZN( us03_n579 ) , .A1( us03_n667 ) , .A2( us03_n786 ) );
  AOI21_X1 us03_U291 (.ZN( us03_n587 ) , .B2( us03_n697 ) , .B1( us03_n813 ) , .A( us03_n815 ) );
  AOI21_X1 us03_U292 (.B1( us03_n697 ) , .ZN( us03_n698 ) , .A( us03_n730 ) , .B2( us03_n761 ) );
  AOI21_X1 us03_U293 (.ZN( us03_n589 ) , .B2( us03_n761 ) , .A( us03_n783 ) , .B1( us03_n810 ) );
  AOI21_X1 us03_U294 (.ZN( us03_n496 ) , .A( us03_n722 ) , .B2( us03_n760 ) , .B1( us03_n812 ) );
  AOI21_X1 us03_U295 (.ZN( us03_n550 ) , .B1( us03_n667 ) , .A( us03_n695 ) , .B2( us03_n803 ) );
  NOR2_X1 us03_U296 (.ZN( us03_n545 ) , .A1( us03_n697 ) , .A2( us03_n742 ) );
  INV_X1 us03_U297 (.A( us03_n727 ) , .ZN( us03_n866 ) );
  INV_X1 us03_U298 (.A( us03_n789 ) , .ZN( us03_n871 ) );
  INV_X1 us03_U299 (.A( us03_n810 ) , .ZN( us03_n852 ) );
  NOR3_X1 us03_U3 (.ZN( us03_n596 ) , .A1( us03_n606 ) , .A3( us03_n721 ) , .A2( us03_n740 ) );
  NOR4_X1 us03_U30 (.A4( us03_n791 ) , .A3( us03_n792 ) , .A2( us03_n793 ) , .A1( us03_n794 ) , .ZN( us03_n795 ) );
  AOI21_X1 us03_U300 (.ZN( us03_n638 ) , .B2( us03_n745 ) , .A( us03_n790 ) , .B1( us03_n801 ) );
  AOI21_X1 us03_U301 (.ZN( us03_n647 ) , .B1( us03_n727 ) , .B2( us03_n761 ) , .A( us03_n811 ) );
  INV_X1 us03_U302 (.A( us03_n784 ) , .ZN( us03_n860 ) );
  NOR2_X1 us03_U303 (.ZN( us03_n683 ) , .A1( us03_n727 ) , .A2( us03_n814 ) );
  AOI21_X1 us03_U304 (.B1( us03_n684 ) , .ZN( us03_n685 ) , .A( us03_n726 ) , .B2( us03_n759 ) );
  AOI21_X1 us03_U305 (.ZN( us03_n567 ) , .B1( us03_n748 ) , .B2( us03_n760 ) , .A( us03_n778 ) );
  AOI21_X1 us03_U306 (.ZN( us03_n498 ) , .A( us03_n695 ) , .B1( us03_n706 ) , .B2( us03_n784 ) );
  NOR2_X1 us03_U307 (.ZN( us03_n566 ) , .A1( us03_n727 ) , .A2( us03_n760 ) );
  AOI21_X1 us03_U308 (.ZN( us03_n637 ) , .B2( us03_n747 ) , .A( us03_n786 ) , .B1( us03_n810 ) );
  NOR2_X1 us03_U309 (.ZN( us03_n564 ) , .A2( us03_n695 ) , .A1( us03_n761 ) );
  NOR4_X1 us03_U31 (.A4( us03_n774 ) , .A3( us03_n775 ) , .A1( us03_n776 ) , .ZN( us03_n797 ) , .A2( us03_n799 ) );
  NOR2_X1 us03_U310 (.ZN( us03_n578 ) , .A2( us03_n695 ) , .A1( us03_n789 ) );
  AOI21_X1 us03_U311 (.ZN( us03_n512 ) , .A( us03_n777 ) , .B2( us03_n790 ) , .B1( us03_n810 ) );
  INV_X1 us03_U312 (.A( us03_n697 ) , .ZN( us03_n851 ) );
  NOR2_X1 us03_U313 (.ZN( us03_n663 ) , .A1( us03_n778 ) , .A2( us03_n811 ) );
  AOI21_X1 us03_U314 (.ZN( us03_n448 ) , .B2( us03_n790 ) , .A( us03_n801 ) , .B1( us03_n813 ) );
  NOR2_X1 us03_U315 (.ZN( us03_n630 ) , .A2( us03_n695 ) , .A1( us03_n722 ) );
  AOI21_X1 us03_U316 (.ZN( us03_n562 ) , .B1( us03_n722 ) , .A( us03_n777 ) , .B2( us03_n789 ) );
  AOI21_X1 us03_U317 (.ZN( us03_n687 ) , .B2( us03_n747 ) , .B1( us03_n761 ) , .A( us03_n804 ) );
  NOR2_X1 us03_U318 (.ZN( us03_n527 ) , .A1( us03_n706 ) , .A2( us03_n777 ) );
  NOR2_X1 us03_U319 (.ZN( us03_n576 ) , .A1( us03_n706 ) , .A2( us03_n811 ) );
  NOR2_X1 us03_U32 (.ZN( us03_n802 ) , .A1( us03_n852 ) , .A2( us03_n859 ) );
  AOI21_X1 us03_U320 (.ZN( us03_n648 ) , .A( us03_n777 ) , .B1( us03_n790 ) , .B2( us03_n803 ) );
  NOR2_X1 us03_U321 (.ZN( us03_n682 ) , .A1( us03_n789 ) , .A2( us03_n811 ) );
  NOR2_X1 us03_U322 (.A2( us03_n811 ) , .A1( us03_n813 ) , .ZN( us03_n819 ) );
  AOI21_X1 us03_U323 (.A( us03_n788 ) , .B2( us03_n789 ) , .B1( us03_n790 ) , .ZN( us03_n791 ) );
  AOI21_X1 us03_U324 (.A( us03_n731 ) , .ZN( us03_n732 ) , .B2( us03_n778 ) , .B1( us03_n790 ) );
  NOR2_X1 us03_U325 (.ZN( us03_n565 ) , .A1( us03_n745 ) , .A2( us03_n803 ) );
  NOR2_X1 us03_U326 (.ZN( us03_n581 ) , .A1( us03_n790 ) , .A2( us03_n815 ) );
  NOR2_X1 us03_U327 (.ZN( us03_n532 ) , .A1( us03_n722 ) , .A2( us03_n786 ) );
  AOI21_X1 us03_U328 (.ZN( us03_n639 ) , .B1( us03_n678 ) , .A( us03_n789 ) , .B2( us03_n815 ) );
  NOR2_X1 us03_U329 (.ZN( us03_n709 ) , .A1( us03_n760 ) , .A2( us03_n761 ) );
  NAND4_X1 us03_U33 (.ZN( sa03_sr_7 ) , .A4( us03_n820 ) , .A3( us03_n821 ) , .A2( us03_n822 ) , .A1( us03_n823 ) );
  NOR2_X1 us03_U330 (.ZN( us03_n680 ) , .A2( us03_n706 ) , .A1( us03_n815 ) );
  INV_X1 us03_U331 (.A( us03_n695 ) , .ZN( us03_n836 ) );
  INV_X1 us03_U332 (.A( us03_n813 ) , .ZN( us03_n853 ) );
  AOI21_X1 us03_U333 (.ZN( us03_n440 ) , .A( us03_n697 ) , .B1( us03_n731 ) , .B2( us03_n748 ) );
  OAI21_X1 us03_U334 (.A( us03_n696 ) , .ZN( us03_n700 ) , .B2( us03_n748 ) , .B1( us03_n802 ) );
  OAI21_X1 us03_U335 (.ZN( us03_n696 ) , .B2( us03_n831 ) , .B1( us03_n836 ) , .A( us03_n858 ) );
  INV_X1 us03_U336 (.A( us03_n778 ) , .ZN( us03_n848 ) );
  AOI22_X1 us03_U337 (.A2( us03_n780 ) , .ZN( us03_n781 ) , .B2( us03_n829 ) , .A1( us03_n832 ) , .B1( us03_n861 ) );
  NAND2_X1 us03_U338 (.ZN( us03_n712 ) , .A1( us03_n726 ) , .A2( us03_n778 ) );
  NAND2_X1 us03_U339 (.ZN( us03_n751 ) , .A1( us03_n761 ) , .A2( us03_n803 ) );
  NOR4_X1 us03_U34 (.A4( us03_n816 ) , .A3( us03_n817 ) , .A2( us03_n818 ) , .A1( us03_n819 ) , .ZN( us03_n820 ) );
  NAND2_X1 us03_U340 (.A2( us03_n760 ) , .A1( us03_n804 ) , .ZN( us03_n808 ) );
  AOI21_X1 us03_U341 (.ZN( us03_n441 ) , .B1( us03_n787 ) , .B2( us03_n789 ) , .A( us03_n812 ) );
  NAND2_X2 us03_U342 (.A1( us03_n449 ) , .A2( us03_n460 ) , .ZN( us03_n788 ) );
  OAI21_X1 us03_U343 (.A( us03_n785 ) , .B2( us03_n786 ) , .B1( us03_n787 ) , .ZN( us03_n793 ) );
  OAI21_X1 us03_U344 (.ZN( us03_n785 ) , .A( us03_n837 ) , .B1( us03_n861 ) , .B2( us03_n871 ) );
  AOI21_X1 us03_U345 (.ZN( us03_n495 ) , .A( us03_n777 ) , .B2( us03_n789 ) , .B1( us03_n802 ) );
  NAND2_X2 us03_U346 (.A2( us03_n439 ) , .A1( us03_n445 ) , .ZN( us03_n782 ) );
  INV_X1 us03_U347 (.A( us03_n783 ) , .ZN( us03_n844 ) );
  NOR2_X1 us03_U348 (.ZN( us03_n468 ) , .A2( us03_n777 ) , .A1( us03_n813 ) );
  OAI21_X1 us03_U349 (.A( us03_n729 ) , .B1( us03_n730 ) , .ZN( us03_n734 ) , .B2( us03_n803 ) );
  AOI222_X1 us03_U35 (.C2( us03_n807 ) , .B2( us03_n808 ) , .A2( us03_n809 ) , .ZN( us03_n821 ) , .C1( us03_n830 ) , .A1( us03_n837 ) , .B1( us03_n851 ) );
  OAI21_X1 us03_U350 (.ZN( us03_n729 ) , .A( us03_n831 ) , .B2( us03_n850 ) , .B1( us03_n871 ) );
  NOR2_X1 us03_U351 (.ZN( us03_n524 ) , .A1( us03_n722 ) , .A2( us03_n748 ) );
  NOR2_X1 us03_U352 (.ZN( us03_n710 ) , .A2( us03_n722 ) , .A1( us03_n788 ) );
  NOR2_X1 us03_U353 (.ZN( us03_n482 ) , .A1( us03_n786 ) , .A2( us03_n803 ) );
  NAND2_X1 us03_U354 (.A1( us03_n697 ) , .A2( us03_n727 ) , .ZN( us03_n780 ) );
  NOR2_X1 us03_U355 (.ZN( us03_n516 ) , .A1( us03_n706 ) , .A2( us03_n786 ) );
  NAND2_X1 us03_U356 (.ZN( us03_n669 ) , .A1( us03_n804 ) , .A2( us03_n814 ) );
  NAND2_X1 us03_U357 (.A2( us03_n747 ) , .A1( us03_n784 ) , .ZN( us03_n807 ) );
  INV_X1 us03_U358 (.A( us03_n722 ) , .ZN( us03_n854 ) );
  INV_X1 us03_U359 (.A( us03_n815 ) , .ZN( us03_n842 ) );
  AOI211_X1 us03_U36 (.B( us03_n805 ) , .A( us03_n806 ) , .ZN( us03_n822 ) , .C1( us03_n840 ) , .C2( us03_n848 ) );
  AND2_X1 us03_U360 (.ZN( us03_n730 ) , .A1( us03_n777 ) , .A2( us03_n783 ) );
  NAND2_X1 us03_U361 (.A1( us03_n453 ) , .A2( us03_n469 ) , .ZN( us03_n801 ) );
  NAND2_X1 us03_U362 (.A1( us03_n449 ) , .A2( us03_n452 ) , .ZN( us03_n812 ) );
  NAND2_X1 us03_U363 (.A1( us03_n449 ) , .A2( us03_n469 ) , .ZN( us03_n814 ) );
  NAND2_X1 us03_U364 (.A1( us03_n452 ) , .A2( us03_n459 ) , .ZN( us03_n811 ) );
  NAND2_X1 us03_U365 (.A1( us03_n451 ) , .A2( us03_n459 ) , .ZN( us03_n742 ) );
  NAND2_X1 us03_U366 (.A1( us03_n450 ) , .A2( us03_n463 ) , .ZN( us03_n667 ) );
  NAND2_X1 us03_U367 (.A2( us03_n446 ) , .A1( us03_n458 ) , .ZN( us03_n726 ) );
  NAND2_X1 us03_U368 (.A1( us03_n453 ) , .A2( us03_n460 ) , .ZN( us03_n748 ) );
  NAND2_X1 us03_U369 (.A2( us03_n451 ) , .A1( us03_n453 ) , .ZN( us03_n804 ) );
  NOR2_X1 us03_U37 (.ZN( us03_n746 ) , .A1( us03_n859 ) , .A2( us03_n860 ) );
  NAND2_X1 us03_U370 (.A2( us03_n452 ) , .A1( us03_n470 ) , .ZN( us03_n777 ) );
  NAND2_X1 us03_U371 (.A1( us03_n451 ) , .A2( us03_n470 ) , .ZN( us03_n783 ) );
  NAND2_X1 us03_U372 (.A2( us03_n462 ) , .A1( us03_n463 ) , .ZN( us03_n810 ) );
  NAND2_X1 us03_U373 (.A1( us03_n439 ) , .A2( us03_n458 ) , .ZN( us03_n697 ) );
  NAND2_X1 us03_U374 (.A2( us03_n447 ) , .A1( us03_n450 ) , .ZN( us03_n761 ) );
  NAND2_X1 us03_U375 (.A2( us03_n446 ) , .A1( us03_n450 ) , .ZN( us03_n727 ) );
  NOR2_X1 us03_U376 (.ZN( us03_n445 ) , .A2( us03_n847 ) , .A1( us03_n856 ) );
  NAND2_X1 us03_U377 (.A2( us03_n459 ) , .A1( us03_n460 ) , .ZN( us03_n745 ) );
  NAND2_X1 us03_U378 (.A1( us03_n460 ) , .A2( us03_n470 ) , .ZN( us03_n786 ) );
  NOR2_X1 us03_U379 (.ZN( us03_n463 ) , .A2( us03_n845 ) , .A1( us03_n846 ) );
  NOR2_X1 us03_U38 (.ZN( us03_n623 ) , .A2( us03_n834 ) , .A1( us03_n837 ) );
  NAND2_X2 us03_U380 (.A2( us03_n459 ) , .A1( us03_n469 ) , .ZN( us03_n695 ) );
  NOR2_X1 us03_U381 (.ZN( us03_n451 ) , .A1( us03_n824 ) , .A2( us03_n825 ) );
  NOR2_X1 us03_U382 (.ZN( us03_n449 ) , .A1( us03_n826 ) , .A2( us03_n827 ) );
  NAND2_X1 us03_U383 (.A2( us03_n452 ) , .A1( us03_n453 ) , .ZN( us03_n728 ) );
  NAND2_X2 us03_U384 (.A2( us03_n446 ) , .A1( us03_n462 ) , .ZN( us03_n813 ) );
  NAND2_X2 us03_U385 (.A2( us03_n439 ) , .A1( us03_n450 ) , .ZN( us03_n789 ) );
  NAND2_X2 us03_U386 (.A1( us03_n447 ) , .A2( us03_n462 ) , .ZN( us03_n722 ) );
  NAND2_X2 us03_U387 (.A1( us03_n447 ) , .A2( us03_n458 ) , .ZN( us03_n790 ) );
  NAND2_X2 us03_U388 (.A1( us03_n439 ) , .A2( us03_n462 ) , .ZN( us03_n706 ) );
  NAND2_X2 us03_U389 (.A2( us03_n469 ) , .A1( us03_n470 ) , .ZN( us03_n815 ) );
  NAND4_X1 us03_U39 (.A4( us03_n601 ) , .A3( us03_n602 ) , .A2( us03_n603 ) , .A1( us03_n604 ) , .ZN( us03_n720 ) );
  NAND2_X2 us03_U390 (.A2( us03_n458 ) , .A1( us03_n463 ) , .ZN( us03_n778 ) );
  NAND2_X1 us03_U391 (.A1( us03_n445 ) , .A2( us03_n447 ) , .ZN( us03_n803 ) );
  NAND2_X2 us03_U392 (.A1( us03_n445 ) , .A2( us03_n446 ) , .ZN( us03_n784 ) );
  NOR2_X1 us03_U393 (.A2( sa03_6 ) , .A1( sa03_7 ) , .ZN( us03_n462 ) );
  NOR2_X1 us03_U394 (.A2( sa03_4 ) , .ZN( us03_n447 ) , .A1( us03_n846 ) );
  NOR2_X1 us03_U395 (.A2( sa03_5 ) , .ZN( us03_n446 ) , .A1( us03_n845 ) );
  NOR2_X1 us03_U396 (.A2( sa03_7 ) , .ZN( us03_n458 ) , .A1( us03_n847 ) );
  NOR2_X1 us03_U397 (.A2( sa03_4 ) , .A1( sa03_5 ) , .ZN( us03_n439 ) );
  NOR2_X1 us03_U398 (.A2( sa03_1 ) , .ZN( us03_n469 ) , .A1( us03_n824 ) );
  NOR2_X1 us03_U399 (.A2( sa03_2 ) , .A1( sa03_3 ) , .ZN( us03_n470 ) );
  NOR3_X1 us03_U4 (.A3( us03_n798 ) , .A2( us03_n799 ) , .A1( us03_n800 ) , .ZN( us03_n823 ) );
  NOR3_X1 us03_U40 (.A1( us03_n597 ) , .ZN( us03_n602 ) , .A3( us03_n661 ) , .A2( us03_n768 ) );
  NOR2_X1 us03_U400 (.A2( sa03_6 ) , .ZN( us03_n450 ) , .A1( us03_n856 ) );
  NOR2_X1 us03_U401 (.A2( sa03_2 ) , .ZN( us03_n459 ) , .A1( us03_n827 ) );
  NOR2_X1 us03_U402 (.A2( sa03_0 ) , .ZN( us03_n452 ) , .A1( us03_n825 ) );
  NOR2_X1 us03_U403 (.A2( sa03_0 ) , .A1( sa03_1 ) , .ZN( us03_n460 ) );
  NOR2_X1 us03_U404 (.A2( sa03_3 ) , .ZN( us03_n453 ) , .A1( us03_n826 ) );
  INV_X1 us03_U405 (.A( sa03_6 ) , .ZN( us03_n847 ) );
  INV_X1 us03_U406 (.A( sa03_3 ) , .ZN( us03_n827 ) );
  INV_X1 us03_U407 (.A( sa03_1 ) , .ZN( us03_n825 ) );
  INV_X1 us03_U408 (.A( sa03_0 ) , .ZN( us03_n824 ) );
  INV_X1 us03_U409 (.A( sa03_2 ) , .ZN( us03_n826 ) );
  NOR4_X1 us03_U41 (.A3( us03_n598 ) , .A2( us03_n599 ) , .A1( us03_n600 ) , .ZN( us03_n601 ) , .A4( us03_n653 ) );
  INV_X1 us03_U410 (.A( sa03_7 ) , .ZN( us03_n856 ) );
  INV_X1 us03_U411 (.A( sa03_5 ) , .ZN( us03_n846 ) );
  AOI222_X1 us03_U412 (.ZN( us03_n603 ) , .B2( us03_n669 ) , .B1( us03_n751 ) , .C2( us03_n829 ) , .A1( us03_n831 ) , .A2( us03_n860 ) , .C1( us03_n861 ) );
  AOI222_X1 us03_U413 (.ZN( us03_n511 ) , .C1( us03_n830 ) , .B2( us03_n835 ) , .A2( us03_n841 ) , .C2( us03_n860 ) , .B1( us03_n861 ) , .A1( us03_n864 ) );
  AOI221_X1 us03_U414 (.A( us03_n481 ) , .ZN( us03_n486 ) , .B1( us03_n829 ) , .C2( us03_n842 ) , .C1( us03_n850 ) , .B2( us03_n860 ) );
  NOR2_X1 us03_U415 (.ZN( us03_n787 ) , .A2( us03_n860 ) , .A1( us03_n866 ) );
  NAND4_X1 us03_U416 (.ZN( sa03_sr_2 ) , .A4( us03_n641 ) , .A3( us03_n642 ) , .A2( us03_n643 ) , .A1( us03_n644 ) );
  OAI221_X1 us03_U417 (.A( us03_n781 ) , .C2( us03_n782 ) , .B2( us03_n783 ) , .B1( us03_n784 ) , .ZN( us03_n794 ) , .C1( us03_n811 ) );
  NAND2_X1 us03_U418 (.A1( us03_n727 ) , .A2( us03_n782 ) , .ZN( us03_n809 ) );
  OAI22_X1 us03_U419 (.ZN( us03_n586 ) , .A2( us03_n745 ) , .B2( us03_n760 ) , .A1( us03_n761 ) , .B1( us03_n782 ) );
  AOI222_X1 us03_U42 (.ZN( us03_n604 ) , .A1( us03_n828 ) , .C2( us03_n835 ) , .B1( us03_n840 ) , .A2( us03_n854 ) , .B2( us03_n859 ) , .C1( us03_n866 ) );
  OAI221_X1 us03_U420 (.A( us03_n694 ) , .ZN( us03_n701 ) , .C2( us03_n782 ) , .C1( us03_n783 ) , .B1( us03_n784 ) , .B2( us03_n804 ) );
  AOI21_X1 us03_U421 (.ZN( us03_n590 ) , .B1( us03_n726 ) , .B2( us03_n782 ) , .A( us03_n788 ) );
  AOI21_X1 us03_U422 (.ZN( us03_n621 ) , .B1( us03_n697 ) , .A( us03_n777 ) , .B2( us03_n782 ) );
  AOI21_X1 us03_U423 (.ZN( us03_n646 ) , .A( us03_n760 ) , .B2( us03_n782 ) , .B1( us03_n790 ) );
  OAI22_X1 us03_U424 (.ZN( us03_n679 ) , .A1( us03_n697 ) , .A2( us03_n728 ) , .B2( us03_n782 ) , .B1( us03_n815 ) );
  OAI21_X1 us03_U425 (.A( us03_n611 ) , .ZN( us03_n614 ) , .B1( us03_n623 ) , .B2( us03_n782 ) );
  NOR2_X1 us03_U426 (.ZN( us03_n608 ) , .A1( us03_n782 ) , .A2( us03_n814 ) );
  OAI222_X1 us03_U427 (.A2( us03_n667 ) , .ZN( us03_n672 ) , .B1( us03_n745 ) , .B2( us03_n782 ) , .C2( us03_n786 ) , .C1( us03_n813 ) , .A1( us03_n815 ) );
  NOR2_X1 us03_U428 (.ZN( us03_n649 ) , .A1( us03_n782 ) , .A2( us03_n786 ) );
  NOR2_X1 us03_U429 (.ZN( us03_n598 ) , .A2( us03_n695 ) , .A1( us03_n782 ) );
  NAND4_X1 us03_U43 (.ZN( sa03_sr_3 ) , .A4( us03_n702 ) , .A3( us03_n703 ) , .A2( us03_n704 ) , .A1( us03_n705 ) );
  NOR2_X1 us03_U430 (.ZN( us03_n551 ) , .A2( us03_n742 ) , .A1( us03_n782 ) );
  INV_X1 us03_U431 (.A( us03_n782 ) , .ZN( us03_n859 ) );
  AOI221_X1 us03_U432 (.A( us03_n574 ) , .ZN( us03_n585 ) , .B2( us03_n829 ) , .C2( us03_n841 ) , .B1( us03_n852 ) , .C1( us03_n859 ) );
  AOI21_X1 us03_U433 (.ZN( us03_n574 ) , .B2( us03_n722 ) , .B1( us03_n746 ) , .A( us03_n783 ) );
  AOI211_X1 us03_U434 (.A( us03_n635 ) , .ZN( us03_n643 ) , .B( us03_n741 ) , .C2( us03_n837 ) , .C1( us03_n852 ) );
  NAND4_X1 us03_U435 (.A4( us03_n631 ) , .A3( us03_n632 ) , .A2( us03_n633 ) , .A1( us03_n634 ) , .ZN( us03_n741 ) );
  INV_X1 us03_U436 (.A( sa03_4 ) , .ZN( us03_n845 ) );
  NAND3_X1 us03_U437 (.ZN( sa03_sr_6 ) , .A3( us03_n795 ) , .A2( us03_n796 ) , .A1( us03_n797 ) );
  NAND3_X1 us03_U438 (.ZN( sa03_sr_5 ) , .A3( us03_n756 ) , .A2( us03_n757 ) , .A1( us03_n758 ) );
  NAND3_X1 us03_U439 (.ZN( sa03_sr_4 ) , .A3( us03_n736 ) , .A2( us03_n737 ) , .A1( us03_n738 ) );
  NOR4_X1 us03_U44 (.A4( us03_n698 ) , .A3( us03_n699 ) , .A2( us03_n700 ) , .A1( us03_n701 ) , .ZN( us03_n702 ) );
  NAND3_X1 us03_U440 (.A3( us03_n673 ) , .A2( us03_n674 ) , .A1( us03_n675 ) , .ZN( us03_n805 ) );
  NAND3_X1 us03_U441 (.ZN( us03_n636 ) , .A3( us03_n706 ) , .A2( us03_n722 ) , .A1( us03_n790 ) );
  NAND3_X1 us03_U442 (.A3( us03_n616 ) , .A2( us03_n617 ) , .A1( us03_n618 ) , .ZN( us03_n723 ) );
  NAND3_X1 us03_U443 (.A3( us03_n583 ) , .A2( us03_n584 ) , .A1( us03_n585 ) , .ZN( us03_n619 ) );
  NAND3_X1 us03_U444 (.ZN( us03_n563 ) , .A3( us03_n678 ) , .A2( us03_n748 ) , .A1( us03_n783 ) );
  NAND3_X1 us03_U445 (.A3( us03_n521 ) , .A2( us03_n522 ) , .A1( us03_n523 ) , .ZN( us03_n740 ) );
  NAND3_X1 us03_U446 (.A3( us03_n510 ) , .A1( us03_n511 ) , .ZN( us03_n606 ) , .A2( us03_n869 ) );
  NAND3_X1 us03_U447 (.A3( us03_n465 ) , .A2( us03_n466 ) , .A1( us03_n467 ) , .ZN( us03_n775 ) );
  AOI211_X1 us03_U45 (.B( us03_n692 ) , .A( us03_n693 ) , .ZN( us03_n703 ) , .C2( us03_n829 ) , .C1( us03_n849 ) );
  NOR2_X1 us03_U46 (.ZN( us03_n705 ) , .A2( us03_n774 ) , .A1( us03_n798 ) );
  AOI222_X1 us03_U47 (.ZN( us03_n467 ) , .B1( us03_n830 ) , .A1( us03_n837 ) , .C1( us03_n840 ) , .C2( us03_n849 ) , .A2( us03_n853 ) , .B2( us03_n863 ) );
  NOR4_X1 us03_U48 (.A1( us03_n464 ) , .ZN( us03_n465 ) , .A4( us03_n540 ) , .A2( us03_n552 ) , .A3( us03_n612 ) );
  AOI221_X1 us03_U49 (.ZN( us03_n466 ) , .C2( us03_n712 ) , .B2( us03_n829 ) , .C1( us03_n843 ) , .B1( us03_n858 ) , .A( us03_n862 ) );
  NOR3_X1 us03_U5 (.ZN( us03_n502 ) , .A2( us03_n677 ) , .A3( us03_n775 ) , .A1( us03_n874 ) );
  NOR4_X1 us03_U50 (.A4( us03_n575 ) , .A3( us03_n576 ) , .A2( us03_n577 ) , .ZN( us03_n584 ) , .A1( us03_n681 ) );
  NOR4_X1 us03_U51 (.A1( us03_n582 ) , .ZN( us03_n583 ) , .A3( us03_n650 ) , .A2( us03_n660 ) , .A4( us03_n765 ) );
  NAND4_X1 us03_U52 (.A4( us03_n483 ) , .A3( us03_n484 ) , .A2( us03_n485 ) , .A1( us03_n486 ) , .ZN( us03_n776 ) );
  NOR4_X1 us03_U53 (.A4( us03_n482 ) , .ZN( us03_n485 ) , .A1( us03_n564 ) , .A2( us03_n579 ) , .A3( us03_n600 ) );
  NOR4_X1 us03_U54 (.ZN( us03_n484 ) , .A1( us03_n505 ) , .A2( us03_n517 ) , .A4( us03_n544 ) , .A3( us03_n609 ) );
  NOR4_X1 us03_U55 (.ZN( us03_n483 ) , .A2( us03_n531 ) , .A1( us03_n556 ) , .A3( us03_n629 ) , .A4( us03_n716 ) );
  AOI211_X1 us03_U56 (.B( us03_n621 ) , .A( us03_n622 ) , .ZN( us03_n633 ) , .C2( us03_n834 ) , .C1( us03_n861 ) );
  NOR4_X1 us03_U57 (.A4( us03_n627 ) , .A3( us03_n628 ) , .A2( us03_n629 ) , .A1( us03_n630 ) , .ZN( us03_n631 ) );
  NOR4_X1 us03_U58 (.A4( us03_n624 ) , .A3( us03_n625 ) , .A2( us03_n626 ) , .ZN( us03_n632 ) , .A1( us03_n662 ) );
  NAND4_X1 us03_U59 (.A4( us03_n655 ) , .A3( us03_n656 ) , .A2( us03_n657 ) , .A1( us03_n658 ) , .ZN( us03_n798 ) );
  INV_X1 us03_U6 (.A( us03_n704 ) , .ZN( us03_n874 ) );
  NOR3_X1 us03_U60 (.A3( us03_n646 ) , .A2( us03_n647 ) , .A1( us03_n648 ) , .ZN( us03_n657 ) );
  NOR3_X1 us03_U61 (.A3( us03_n649 ) , .A2( us03_n650 ) , .A1( us03_n651 ) , .ZN( us03_n656 ) );
  NOR3_X1 us03_U62 (.A3( us03_n652 ) , .A2( us03_n653 ) , .A1( us03_n654 ) , .ZN( us03_n655 ) );
  NAND4_X1 us03_U63 (.A4( us03_n558 ) , .A3( us03_n559 ) , .A2( us03_n560 ) , .A1( us03_n561 ) , .ZN( us03_n605 ) );
  NOR4_X1 us03_U64 (.A4( us03_n554 ) , .A3( us03_n555 ) , .A2( us03_n556 ) , .A1( us03_n557 ) , .ZN( us03_n558 ) );
  NOR4_X1 us03_U65 (.ZN( us03_n559 ) , .A1( us03_n651 ) , .A3( us03_n659 ) , .A4( us03_n683 ) , .A2( us03_n766 ) );
  NOR4_X1 us03_U66 (.A4( us03_n550 ) , .A3( us03_n551 ) , .A2( us03_n552 ) , .A1( us03_n553 ) , .ZN( us03_n560 ) );
  NAND4_X1 us03_U67 (.A4( us03_n770 ) , .A3( us03_n771 ) , .A2( us03_n772 ) , .A1( us03_n773 ) , .ZN( us03_n799 ) );
  NOR3_X1 us03_U68 (.A3( us03_n763 ) , .A2( us03_n764 ) , .A1( us03_n765 ) , .ZN( us03_n771 ) );
  NOR4_X1 us03_U69 (.A4( us03_n766 ) , .A3( us03_n767 ) , .A2( us03_n768 ) , .A1( us03_n769 ) , .ZN( us03_n770 ) );
  NOR3_X1 us03_U7 (.A3( us03_n619 ) , .A2( us03_n620 ) , .ZN( us03_n634 ) , .A1( us03_n723 ) );
  AOI222_X1 us03_U70 (.ZN( us03_n773 ) , .A1( us03_n828 ) , .C1( us03_n832 ) , .B2( us03_n839 ) , .A2( us03_n848 ) , .B1( us03_n859 ) , .C2( us03_n871 ) );
  NOR4_X1 us03_U71 (.A4( us03_n507 ) , .A2( us03_n508 ) , .A1( us03_n509 ) , .ZN( us03_n510 ) , .A3( us03_n668 ) );
  INV_X1 us03_U72 (.A( us03_n503 ) , .ZN( us03_n869 ) );
  NOR4_X1 us03_U73 (.A4( us03_n663 ) , .A3( us03_n664 ) , .A2( us03_n665 ) , .A1( us03_n666 ) , .ZN( us03_n674 ) );
  NOR4_X1 us03_U74 (.A4( us03_n659 ) , .A3( us03_n660 ) , .A2( us03_n661 ) , .A1( us03_n662 ) , .ZN( us03_n675 ) );
  NOR4_X1 us03_U75 (.A3( us03_n671 ) , .A1( us03_n672 ) , .ZN( us03_n673 ) , .A4( us03_n713 ) , .A2( us03_n857 ) );
  NOR2_X1 us03_U76 (.ZN( us03_n759 ) , .A1( us03_n831 ) , .A2( us03_n832 ) );
  NOR4_X1 us03_U77 (.A4( us03_n732 ) , .A3( us03_n733 ) , .A2( us03_n734 ) , .A1( us03_n735 ) , .ZN( us03_n736 ) );
  AOI211_X1 us03_U78 (.B( us03_n723 ) , .A( us03_n724 ) , .ZN( us03_n737 ) , .C1( us03_n841 ) , .C2( us03_n853 ) );
  NOR3_X1 us03_U79 (.A3( us03_n720 ) , .A1( us03_n721 ) , .ZN( us03_n738 ) , .A2( us03_n739 ) );
  NOR2_X1 us03_U8 (.ZN( us03_n573 ) , .A1( us03_n620 ) , .A2( us03_n743 ) );
  NOR4_X1 us03_U80 (.A3( us03_n753 ) , .A2( us03_n754 ) , .A1( us03_n755 ) , .ZN( us03_n756 ) , .A4( us03_n867 ) );
  AOI211_X1 us03_U81 (.B( us03_n743 ) , .A( us03_n744 ) , .ZN( us03_n757 ) , .C1( us03_n830 ) , .C2( us03_n851 ) );
  NOR3_X1 us03_U82 (.A3( us03_n739 ) , .A2( us03_n740 ) , .A1( us03_n741 ) , .ZN( us03_n758 ) );
  NAND4_X1 us03_U83 (.A4( us03_n454 ) , .A3( us03_n455 ) , .A2( us03_n456 ) , .A1( us03_n457 ) , .ZN( us03_n677 ) );
  NOR3_X1 us03_U84 (.ZN( us03_n455 ) , .A3( us03_n528 ) , .A1( us03_n553 ) , .A2( us03_n568 ) );
  AOI221_X1 us03_U85 (.A( us03_n448 ) , .ZN( us03_n457 ) , .C2( us03_n751 ) , .B1( us03_n830 ) , .C1( us03_n840 ) , .B2( us03_n859 ) );
  NOR4_X1 us03_U86 (.ZN( us03_n456 ) , .A2( us03_n507 ) , .A1( us03_n597 ) , .A4( us03_n626 ) , .A3( us03_n709 ) );
  NAND4_X1 us03_U87 (.A4( us03_n533 ) , .A3( us03_n534 ) , .A2( us03_n535 ) , .A1( us03_n536 ) , .ZN( us03_n620 ) );
  NOR4_X1 us03_U88 (.A4( us03_n524 ) , .A2( us03_n525 ) , .A1( us03_n526 ) , .ZN( us03_n536 ) , .A3( us03_n699 ) );
  NOR4_X1 us03_U89 (.A1( us03_n529 ) , .ZN( us03_n534 ) , .A2( us03_n652 ) , .A4( us03_n666 ) , .A3( us03_n763 ) );
  NOR2_X1 us03_U9 (.A1( us03_n676 ) , .ZN( us03_n691 ) , .A2( us03_n805 ) );
  NOR4_X1 us03_U90 (.A4( us03_n527 ) , .A3( us03_n528 ) , .ZN( us03_n535 ) , .A2( us03_n682 ) , .A1( us03_n792 ) );
  NAND4_X1 us03_U91 (.A4( us03_n477 ) , .A3( us03_n478 ) , .A2( us03_n479 ) , .A1( us03_n480 ) , .ZN( us03_n692 ) );
  NOR3_X1 us03_U92 (.ZN( us03_n478 ) , .A2( us03_n506 ) , .A3( us03_n599 ) , .A1( us03_n608 ) );
  AOI211_X1 us03_U93 (.B( us03_n475 ) , .A( us03_n476 ) , .ZN( us03_n480 ) , .C2( us03_n831 ) , .C1( us03_n859 ) );
  NOR4_X1 us03_U94 (.ZN( us03_n479 ) , .A3( us03_n530 ) , .A4( us03_n543 ) , .A2( us03_n565 ) , .A1( us03_n715 ) );
  NAND4_X1 us03_U95 (.A4( us03_n546 ) , .A3( us03_n547 ) , .A2( us03_n548 ) , .A1( us03_n549 ) , .ZN( us03_n743 ) );
  NOR3_X1 us03_U96 (.ZN( us03_n547 ) , .A2( us03_n649 ) , .A1( us03_n665 ) , .A3( us03_n769 ) );
  AOI211_X1 us03_U97 (.B( us03_n537 ) , .A( us03_n538 ) , .ZN( us03_n549 ) , .C2( us03_n837 ) , .C1( us03_n849 ) );
  NOR4_X1 us03_U98 (.A4( us03_n542 ) , .A3( us03_n543 ) , .A2( us03_n544 ) , .A1( us03_n545 ) , .ZN( us03_n546 ) );
  NOR4_X1 us03_U99 (.ZN( us03_n618 ) , .A1( us03_n654 ) , .A3( us03_n664 ) , .A4( us03_n680 ) , .A2( us03_n764 ) );
  INV_X1 us20_U10 (.A( us20_n706 ) , .ZN( us20_n876 ) );
  NOR4_X1 us20_U100 (.A1( us20_n531 ) , .ZN( us20_n536 ) , .A2( us20_n654 ) , .A4( us20_n668 ) , .A3( us20_n765 ) );
  NOR4_X1 us20_U101 (.A4( us20_n529 ) , .A3( us20_n530 ) , .ZN( us20_n537 ) , .A2( us20_n684 ) , .A1( us20_n794 ) );
  NAND4_X1 us20_U102 (.A4( us20_n548 ) , .A3( us20_n549 ) , .A2( us20_n550 ) , .A1( us20_n551 ) , .ZN( us20_n745 ) );
  NOR3_X1 us20_U103 (.ZN( us20_n549 ) , .A2( us20_n651 ) , .A1( us20_n667 ) , .A3( us20_n771 ) );
  AOI211_X1 us20_U104 (.B( us20_n539 ) , .A( us20_n540 ) , .ZN( us20_n551 ) , .C2( us20_n839 ) , .C1( us20_n851 ) );
  NOR4_X1 us20_U105 (.A4( us20_n541 ) , .A3( us20_n542 ) , .A2( us20_n543 ) , .ZN( us20_n550 ) , .A1( us20_n688 ) );
  NAND4_X1 us20_U106 (.A4( us20_n479 ) , .A3( us20_n480 ) , .A2( us20_n481 ) , .A1( us20_n482 ) , .ZN( us20_n694 ) );
  NOR3_X1 us20_U107 (.ZN( us20_n480 ) , .A2( us20_n508 ) , .A3( us20_n601 ) , .A1( us20_n610 ) );
  AOI211_X1 us20_U108 (.B( us20_n477 ) , .A( us20_n478 ) , .ZN( us20_n482 ) , .C2( us20_n833 ) , .C1( us20_n861 ) );
  NOR4_X1 us20_U109 (.ZN( us20_n481 ) , .A3( us20_n532 ) , .A4( us20_n545 ) , .A2( us20_n567 ) , .A1( us20_n717 ) );
  INV_X1 us20_U11 (.A( us20_n607 ) , .ZN( us20_n874 ) );
  NOR2_X1 us20_U110 (.ZN( us20_n647 ) , .A1( us20_n854 ) , .A2( us20_n868 ) );
  NAND4_X1 us20_U111 (.A4( us20_n473 ) , .A3( us20_n474 ) , .A2( us20_n475 ) , .A1( us20_n476 ) , .ZN( us20_n678 ) );
  NOR4_X1 us20_U112 (.ZN( us20_n475 ) , .A1( us20_n531 ) , .A3( us20_n568 ) , .A4( us20_n600 ) , .A2( us20_n642 ) );
  NOR4_X1 us20_U113 (.A4( us20_n470 ) , .ZN( us20_n476 ) , .A3( us20_n556 ) , .A1( us20_n735 ) , .A2( us20_n755 ) );
  NOR4_X1 us20_U114 (.ZN( us20_n474 ) , .A1( us20_n506 ) , .A3( us20_n544 ) , .A2( us20_n583 ) , .A4( us20_n716 ) );
  NAND4_X1 us20_U115 (.A4( us20_n691 ) , .A3( us20_n692 ) , .A1( us20_n693 ) , .ZN( us20_n776 ) , .A2( us20_n872 ) );
  INV_X1 us20_U116 (.A( us20_n679 ) , .ZN( us20_n872 ) );
  AOI221_X1 us20_U117 (.A( us20_n681 ) , .ZN( us20_n692 ) , .B2( us20_n840 ) , .C1( us20_n842 ) , .C2( us20_n862 ) , .B1( us20_n865 ) );
  NOR4_X1 us20_U118 (.A4( us20_n687 ) , .A3( us20_n688 ) , .A2( us20_n689 ) , .A1( us20_n690 ) , .ZN( us20_n691 ) );
  NOR2_X1 us20_U119 (.ZN( us20_n733 ) , .A2( us20_n832 ) , .A1( us20_n845 ) );
  INV_X1 us20_U12 (.A( us20_n680 ) , .ZN( us20_n840 ) );
  NAND4_X1 us20_U120 (.A4( us20_n719 ) , .A3( us20_n720 ) , .A2( us20_n721 ) , .ZN( us20_n741 ) , .A1( us20_n857 ) );
  INV_X1 us20_U121 (.A( us20_n709 ) , .ZN( us20_n857 ) );
  NOR4_X1 us20_U122 (.A4( us20_n715 ) , .A3( us20_n716 ) , .A2( us20_n717 ) , .A1( us20_n718 ) , .ZN( us20_n719 ) );
  AOI221_X1 us20_U123 (.A( us20_n710 ) , .ZN( us20_n721 ) , .C2( us20_n844 ) , .B2( us20_n845 ) , .C1( us20_n861 ) , .B1( us20_n862 ) );
  NAND4_X1 us20_U124 (.A4( us20_n573 ) , .A3( us20_n574 ) , .A1( us20_n575 ) , .ZN( us20_n723 ) , .A2( us20_n874 ) );
  NOR4_X1 us20_U125 (.A4( us20_n569 ) , .A3( us20_n570 ) , .A2( us20_n571 ) , .A1( us20_n572 ) , .ZN( us20_n573 ) );
  AOI221_X1 us20_U126 (.A( us20_n564 ) , .C2( us20_n565 ) , .ZN( us20_n574 ) , .B2( us20_n845 ) , .B1( us20_n852 ) , .C1( us20_n853 ) );
  NOR2_X1 us20_U127 (.ZN( us20_n575 ) , .A1( us20_n622 ) , .A2( us20_n745 ) );
  NAND4_X1 us20_U128 (.A4( us20_n633 ) , .A3( us20_n634 ) , .A2( us20_n635 ) , .A1( us20_n636 ) , .ZN( us20_n743 ) );
  AOI211_X1 us20_U129 (.B( us20_n623 ) , .A( us20_n624 ) , .ZN( us20_n635 ) , .C2( us20_n836 ) , .C1( us20_n863 ) );
  NOR4_X1 us20_U13 (.A4( us20_n445 ) , .A3( us20_n446 ) , .A2( us20_n516 ) , .A1( us20_n541 ) , .ZN( us20_n706 ) );
  NOR4_X1 us20_U130 (.A4( us20_n629 ) , .A3( us20_n630 ) , .A2( us20_n631 ) , .A1( us20_n632 ) , .ZN( us20_n633 ) );
  NOR4_X1 us20_U131 (.A4( us20_n626 ) , .A3( us20_n627 ) , .A2( us20_n628 ) , .ZN( us20_n634 ) , .A1( us20_n664 ) );
  NAND4_X1 us20_U132 (.A4( us20_n493 ) , .A3( us20_n494 ) , .A1( us20_n495 ) , .ZN( us20_n802 ) , .A2( us20_n867 ) );
  AOI221_X1 us20_U133 (.A( us20_n489 ) , .ZN( us20_n494 ) , .B2( us20_n836 ) , .C2( us20_n841 ) , .C1( us20_n851 ) , .B1( us20_n860 ) );
  INV_X1 us20_U134 (.A( us20_n778 ) , .ZN( us20_n867 ) );
  NOR4_X1 us20_U135 (.A2( us20_n491 ) , .A1( us20_n492 ) , .ZN( us20_n493 ) , .A3( us20_n580 ) , .A4( us20_n612 ) );
  INV_X1 us20_U136 (.A( us20_n762 ) , .ZN( us20_n830 ) );
  OR4_X1 us20_U137 (.A4( us20_n580 ) , .A3( us20_n581 ) , .A2( us20_n582 ) , .A1( us20_n583 ) , .ZN( us20_n584 ) );
  OR4_X1 us20_U138 (.A4( us20_n566 ) , .A3( us20_n567 ) , .A2( us20_n568 ) , .ZN( us20_n572 ) , .A1( us20_n665 ) );
  OR4_X1 us20_U139 (.A4( us20_n682 ) , .A3( us20_n683 ) , .A2( us20_n684 ) , .A1( us20_n685 ) , .ZN( us20_n690 ) );
  OR3_X1 us20_U14 (.ZN( us20_n446 ) , .A1( us20_n528 ) , .A3( us20_n577 ) , .A2( us20_n875 ) );
  OR4_X1 us20_U140 (.ZN( us20_n466 ) , .A4( us20_n518 ) , .A3( us20_n529 ) , .A2( us20_n578 ) , .A1( us20_n712 ) );
  OR4_X1 us20_U141 (.A4( us20_n518 ) , .A2( us20_n519 ) , .A1( us20_n520 ) , .ZN( us20_n522 ) , .A3( us20_n821 ) );
  OR4_X1 us20_U142 (.ZN( us20_n492 ) , .A4( us20_n534 ) , .A2( us20_n547 ) , .A1( us20_n559 ) , .A3( us20_n632 ) );
  NAND2_X1 us20_U143 (.ZN( us20_n613 ) , .A2( us20_n837 ) , .A1( us20_n873 ) );
  OR3_X1 us20_U144 (.A3( us20_n506 ) , .A2( us20_n507 ) , .A1( us20_n508 ) , .ZN( us20_n511 ) );
  AOI221_X1 us20_U145 (.A( us20_n713 ) , .B2( us20_n714 ) , .ZN( us20_n720 ) , .C1( us20_n832 ) , .B1( us20_n839 ) , .C2( us20_n863 ) );
  OR2_X1 us20_U146 (.A2( us20_n711 ) , .A1( us20_n712 ) , .ZN( us20_n713 ) );
  INV_X1 us20_U147 (.A( us20_n463 ) , .ZN( us20_n864 ) );
  OAI21_X1 us20_U148 (.ZN( us20_n463 ) , .B1( us20_n809 ) , .A( us20_n834 ) , .B2( us20_n851 ) );
  INV_X1 us20_U149 (.A( us20_n754 ) , .ZN( us20_n869 ) );
  OR4_X1 us20_U15 (.A4( us20_n442 ) , .A2( us20_n443 ) , .A1( us20_n444 ) , .ZN( us20_n445 ) , .A3( us20_n553 ) );
  OAI21_X1 us20_U150 (.B1( us20_n753 ) , .ZN( us20_n754 ) , .A( us20_n845 ) , .B2( us20_n868 ) );
  AOI222_X1 us20_U151 (.ZN( us20_n660 ) , .A2( us20_n839 ) , .B1( us20_n841 ) , .C2( us20_n845 ) , .A1( us20_n860 ) , .C1( us20_n863 ) , .B2( us20_n870 ) );
  INV_X1 us20_U152 (.A( us20_n647 ) , .ZN( us20_n870 ) );
  INV_X1 us20_U153 (.A( us20_n672 ) , .ZN( us20_n859 ) );
  AOI21_X1 us20_U154 (.A( us20_n670 ) , .B1( us20_n671 ) , .ZN( us20_n672 ) , .B2( us20_n856 ) );
  OAI22_X1 us20_U155 (.ZN( us20_n483 ) , .A1( us20_n708 ) , .B2( us20_n785 ) , .A2( us20_n806 ) , .B1( us20_n812 ) );
  OAI222_X1 us20_U156 (.B2( us20_n747 ) , .B1( us20_n748 ) , .A2( us20_n749 ) , .ZN( us20_n757 ) , .C2( us20_n805 ) , .C1( us20_n814 ) , .A1( us20_n817 ) );
  OAI222_X1 us20_U157 (.B2( us20_n708 ) , .ZN( us20_n709 ) , .C2( us20_n724 ) , .B1( us20_n747 ) , .A1( us20_n806 ) , .C1( us20_n814 ) , .A2( us20_n815 ) );
  OAI222_X1 us20_U158 (.ZN( us20_n505 ) , .C2( us20_n625 ) , .B2( us20_n647 ) , .B1( us20_n747 ) , .A2( us20_n748 ) , .C1( us20_n805 ) , .A1( us20_n806 ) );
  NAND2_X1 us20_U159 (.A1( us20_n447 ) , .A2( us20_n465 ) , .ZN( us20_n749 ) );
  INV_X1 us20_U16 (.A( us20_n613 ) , .ZN( us20_n875 ) );
  AOI22_X1 us20_U160 (.ZN( us20_n696 ) , .A1( us20_n830 ) , .B2( us20_n843 ) , .A2( us20_n865 ) , .B1( us20_n868 ) );
  AOI22_X1 us20_U161 (.A2( us20_n782 ) , .ZN( us20_n783 ) , .B2( us20_n831 ) , .A1( us20_n834 ) , .B1( us20_n863 ) );
  INV_X1 us20_U162 (.A( us20_n730 ) , .ZN( us20_n839 ) );
  INV_X1 us20_U163 (.A( us20_n790 ) , .ZN( us20_n832 ) );
  NAND2_X1 us20_U164 (.A1( us20_n451 ) , .A2( us20_n453 ) , .ZN( us20_n762 ) );
  AOI211_X1 us20_U165 (.A( us20_n637 ) , .ZN( us20_n645 ) , .B( us20_n743 ) , .C2( us20_n839 ) , .C1( us20_n854 ) );
  OAI22_X1 us20_U166 (.ZN( us20_n637 ) , .A1( us20_n699 ) , .B2( us20_n728 ) , .A2( us20_n762 ) , .B1( us20_n816 ) );
  OAI221_X1 us20_U167 (.A( us20_n727 ) , .C2( us20_n728 ) , .B2( us20_n729 ) , .B1( us20_n730 ) , .ZN( us20_n737 ) , .C1( us20_n817 ) );
  AOI22_X1 us20_U168 (.ZN( us20_n727 ) , .B1( us20_n832 ) , .A2( us20_n838 ) , .A1( us20_n863 ) , .B2( us20_n866 ) );
  OAI22_X1 us20_U169 (.ZN( us20_n489 ) , .A1( us20_n724 ) , .B2( us20_n728 ) , .B1( us20_n730 ) , .A2( us20_n779 ) );
  INV_X1 us20_U17 (.A( us20_n749 ) , .ZN( us20_n863 ) );
  OAI22_X1 us20_U170 (.ZN( us20_n624 ) , .B1( us20_n669 ) , .B2( us20_n747 ) , .A1( us20_n815 ) , .A2( us20_n816 ) );
  OAI22_X1 us20_U171 (.B2( us20_n779 ) , .B1( us20_n780 ) , .ZN( us20_n781 ) , .A2( us20_n814 ) , .A1( us20_n815 ) );
  OAI22_X1 us20_U172 (.A1( us20_n724 ) , .ZN( us20_n726 ) , .B2( us20_n750 ) , .B1( us20_n812 ) , .A2( us20_n816 ) );
  OAI22_X1 us20_U173 (.B2( us20_n744 ) , .ZN( us20_n746 ) , .A2( us20_n762 ) , .B1( us20_n780 ) , .A1( us20_n792 ) );
  OAI22_X1 us20_U174 (.ZN( us20_n496 ) , .A2( us20_n744 ) , .A1( us20_n780 ) , .B1( us20_n791 ) , .B2( us20_n806 ) );
  OAI22_X1 us20_U175 (.B2( us20_n803 ) , .B1( us20_n804 ) , .A2( us20_n805 ) , .A1( us20_n806 ) , .ZN( us20_n808 ) );
  INV_X1 us20_U176 (.A( us20_n788 ) , .ZN( us20_n845 ) );
  INV_X1 us20_U177 (.A( us20_n744 ) , .ZN( us20_n837 ) );
  INV_X1 us20_U178 (.A( us20_n814 ) , .ZN( us20_n833 ) );
  OAI22_X1 us20_U179 (.B1( us20_n490 ) , .ZN( us20_n491 ) , .A1( us20_n686 ) , .A2( us20_n763 ) , .B2( us20_n817 ) );
  AOI222_X1 us20_U18 (.ZN( us20_n563 ) , .B1( us20_n830 ) , .C1( us20_n841 ) , .A2( us20_n843 ) , .A1( us20_n854 ) , .B2( us20_n863 ) , .C2( us20_n873 ) );
  NOR3_X1 us20_U180 (.ZN( us20_n490 ) , .A1( us20_n782 ) , .A2( us20_n850 ) , .A3( us20_n863 ) );
  OAI22_X1 us20_U181 (.ZN( us20_n695 ) , .A2( us20_n730 ) , .A1( us20_n780 ) , .B1( us20_n791 ) , .B2( us20_n817 ) );
  INV_X1 us20_U182 (.A( us20_n805 ) , .ZN( us20_n860 ) );
  INV_X1 us20_U183 (.A( us20_n669 ) , .ZN( us20_n865 ) );
  NOR2_X1 us20_U184 (.ZN( us20_n715 ) , .A1( us20_n805 ) , .A2( us20_n817 ) );
  NOR2_X1 us20_U185 (.ZN( us20_n666 ) , .A1( us20_n728 ) , .A2( us20_n803 ) );
  NOR2_X1 us20_U186 (.ZN( us20_n546 ) , .A2( us20_n780 ) , .A1( us20_n814 ) );
  NOR2_X1 us20_U187 (.ZN( us20_n577 ) , .A2( us20_n699 ) , .A1( us20_n814 ) );
  NOR2_X1 us20_U188 (.ZN( us20_n570 ) , .A1( us20_n728 ) , .A2( us20_n806 ) );
  NOR2_X1 us20_U189 (.A2( us20_n744 ) , .ZN( us20_n755 ) , .A1( us20_n805 ) );
  NOR4_X1 us20_U19 (.ZN( us20_n473 ) , .A2( us20_n521 ) , .A4( us20_n594 ) , .A1( us20_n609 ) , .A3( us20_n629 ) );
  NOR2_X1 us20_U190 (.ZN( us20_n718 ) , .A2( us20_n724 ) , .A1( us20_n744 ) );
  NOR2_X1 us20_U191 (.ZN( us20_n735 ) , .A2( us20_n803 ) , .A1( us20_n805 ) );
  INV_X1 us20_U192 (.A( us20_n750 ) , .ZN( us20_n842 ) );
  NOR2_X1 us20_U193 (.ZN( us20_n532 ) , .A2( us20_n749 ) , .A1( us20_n750 ) );
  NOR2_X1 us20_U194 (.ZN( us20_n654 ) , .A1( us20_n728 ) , .A2( us20_n813 ) );
  NOR2_X1 us20_U195 (.ZN( us20_n615 ) , .A1( us20_n785 ) , .A2( us20_n815 ) );
  NOR2_X1 us20_U196 (.ZN( us20_n629 ) , .A2( us20_n728 ) , .A1( us20_n785 ) );
  NOR2_X1 us20_U197 (.ZN( us20_n628 ) , .A2( us20_n669 ) , .A1( us20_n785 ) );
  NOR2_X1 us20_U198 (.ZN( us20_n611 ) , .A2( us20_n780 ) , .A1( us20_n806 ) );
  INV_X1 us20_U199 (.A( us20_n747 ) , .ZN( us20_n834 ) );
  NOR4_X1 us20_U20 (.A4( us20_n544 ) , .A3( us20_n545 ) , .A2( us20_n546 ) , .A1( us20_n547 ) , .ZN( us20_n548 ) );
  NOR2_X1 us20_U200 (.ZN( us20_n601 ) , .A2( us20_n780 ) , .A1( us20_n803 ) );
  NOR2_X1 us20_U201 (.A2( us20_n708 ) , .A1( us20_n750 ) , .ZN( us20_n771 ) );
  NOR2_X1 us20_U202 (.ZN( us20_n652 ) , .A1( us20_n669 ) , .A2( us20_n814 ) );
  INV_X1 us20_U203 (.A( us20_n792 ) , .ZN( us20_n851 ) );
  NOR2_X1 us20_U204 (.A1( us20_n669 ) , .ZN( us20_n673 ) , .A2( us20_n744 ) );
  NOR2_X1 us20_U205 (.ZN( us20_n602 ) , .A1( us20_n669 ) , .A2( us20_n803 ) );
  NOR2_X1 us20_U206 (.A1( us20_n669 ) , .ZN( us20_n688 ) , .A2( us20_n816 ) );
  NOR2_X1 us20_U207 (.ZN( us20_n667 ) , .A1( us20_n750 ) , .A2( us20_n815 ) );
  NOR2_X1 us20_U208 (.A2( us20_n744 ) , .ZN( us20_n769 ) , .A1( us20_n812 ) );
  NOR2_X1 us20_U209 (.ZN( us20_n555 ) , .A1( us20_n750 ) , .A2( us20_n791 ) );
  NOR4_X1 us20_U21 (.ZN( us20_n479 ) , .A1( us20_n520 ) , .A4( us20_n557 ) , .A3( us20_n582 ) , .A2( us20_n630 ) );
  NOR2_X1 us20_U210 (.ZN( us20_n528 ) , .A2( us20_n724 ) , .A1( us20_n803 ) );
  NOR2_X1 us20_U211 (.ZN( us20_n508 ) , .A2( us20_n780 ) , .A1( us20_n785 ) );
  NOR2_X1 us20_U212 (.ZN( us20_n543 ) , .A2( us20_n708 ) , .A1( us20_n785 ) );
  NOR2_X1 us20_U213 (.ZN( us20_n531 ) , .A2( us20_n780 ) , .A1( us20_n816 ) );
  NOR2_X1 us20_U214 (.ZN( us20_n664 ) , .A1( us20_n785 ) , .A2( us20_n791 ) );
  NOR2_X1 us20_U215 (.ZN( us20_n599 ) , .A2( us20_n791 ) , .A1( us20_n816 ) );
  NOR2_X1 us20_U216 (.A1( us20_n669 ) , .ZN( us20_n766 ) , .A2( us20_n813 ) );
  NOR2_X1 us20_U217 (.A1( us20_n699 ) , .ZN( us20_n768 ) , .A2( us20_n813 ) );
  NOR2_X1 us20_U218 (.ZN( us20_n527 ) , .A1( us20_n669 ) , .A2( us20_n779 ) );
  OAI22_X1 us20_U219 (.B1( us20_n440 ) , .ZN( us20_n444 ) , .A2( us20_n728 ) , .A1( us20_n744 ) , .B2( us20_n749 ) );
  NOR4_X1 us20_U22 (.A4( us20_n532 ) , .A3( us20_n533 ) , .A2( us20_n534 ) , .ZN( us20_n535 ) , .A1( us20_n820 ) );
  NOR3_X1 us20_U220 (.ZN( us20_n440 ) , .A2( us20_n836 ) , .A3( us20_n837 ) , .A1( us20_n846 ) );
  OAI22_X1 us20_U221 (.ZN( us20_n710 ) , .A2( us20_n728 ) , .B2( us20_n729 ) , .A1( us20_n744 ) , .B1( us20_n813 ) );
  NOR2_X1 us20_U222 (.ZN( us20_n557 ) , .A1( us20_n792 ) , .A2( us20_n814 ) );
  NOR2_X1 us20_U223 (.ZN( us20_n545 ) , .A1( us20_n749 ) , .A2( us20_n814 ) );
  NOR2_X1 us20_U224 (.ZN( us20_n556 ) , .A1( us20_n762 ) , .A2( us20_n805 ) );
  NOR2_X1 us20_U225 (.ZN( us20_n661 ) , .A1( us20_n729 ) , .A2( us20_n790 ) );
  NOR2_X1 us20_U226 (.ZN( us20_n507 ) , .A1( us20_n812 ) , .A2( us20_n817 ) );
  INV_X1 us20_U227 (.A( us20_n806 ) , .ZN( us20_n841 ) );
  NOR2_X1 us20_U228 (.ZN( us20_n509 ) , .A1( us20_n729 ) , .A2( us20_n779 ) );
  NOR2_X1 us20_U229 (.ZN( us20_n544 ) , .A2( us20_n785 ) , .A1( us20_n792 ) );
  NOR4_X1 us20_U23 (.ZN( us20_n456 ) , .A2( us20_n517 ) , .A1( us20_n543 ) , .A3( us20_n579 ) , .A4( us20_n615 ) );
  OAI22_X1 us20_U230 (.B2( us20_n750 ) , .B1( us20_n751 ) , .A1( us20_n752 ) , .ZN( us20_n756 ) , .A2( us20_n806 ) );
  NOR2_X1 us20_U231 (.ZN( us20_n751 ) , .A2( us20_n852 ) , .A1( us20_n860 ) );
  NOR3_X1 us20_U232 (.ZN( us20_n752 ) , .A2( us20_n853 ) , .A1( us20_n863 ) , .A3( us20_n865 ) );
  NOR2_X1 us20_U233 (.ZN( us20_n530 ) , .A2( us20_n744 ) , .A1( us20_n792 ) );
  NOR2_X1 us20_U234 (.ZN( us20_n663 ) , .A1( us20_n729 ) , .A2( us20_n785 ) );
  INV_X1 us20_U235 (.A( us20_n728 ) , .ZN( us20_n852 ) );
  NOR2_X1 us20_U236 (.A1( us20_n749 ) , .ZN( us20_n767 ) , .A2( us20_n803 ) );
  NOR2_X1 us20_U237 (.ZN( us20_n506 ) , .A2( us20_n728 ) , .A1( us20_n762 ) );
  NOR2_X1 us20_U238 (.ZN( us20_n516 ) , .A1( us20_n708 ) , .A2( us20_n744 ) );
  NOR2_X1 us20_U239 (.ZN( us20_n614 ) , .A1( us20_n762 ) , .A2( us20_n812 ) );
  NOR2_X1 us20_U24 (.ZN( us20_n680 ) , .A2( us20_n834 ) , .A1( us20_n839 ) );
  NOR2_X1 us20_U240 (.ZN( us20_n670 ) , .A1( us20_n790 ) , .A2( us20_n805 ) );
  NOR2_X1 us20_U241 (.ZN( us20_n517 ) , .A1( us20_n708 ) , .A2( us20_n803 ) );
  NOR2_X1 us20_U242 (.ZN( us20_n558 ) , .A1( us20_n708 ) , .A2( us20_n816 ) );
  NOR2_X1 us20_U243 (.ZN( us20_n630 ) , .A1( us20_n747 ) , .A2( us20_n815 ) );
  NOR2_X1 us20_U244 (.ZN( us20_n655 ) , .A1( us20_n790 ) , .A2( us20_n815 ) );
  NOR2_X1 us20_U245 (.ZN( us20_n521 ) , .A1( us20_n790 ) , .A2( us20_n812 ) );
  NOR2_X1 us20_U246 (.ZN( us20_n668 ) , .A2( us20_n708 ) , .A1( us20_n790 ) );
  NOR2_X1 us20_U247 (.ZN( us20_n631 ) , .A1( us20_n724 ) , .A2( us20_n813 ) );
  NOR2_X1 us20_U248 (.ZN( us20_n656 ) , .A1( us20_n747 ) , .A2( us20_n780 ) );
  NOR2_X1 us20_U249 (.ZN( us20_n542 ) , .A1( us20_n762 ) , .A2( us20_n791 ) );
  NOR4_X1 us20_U25 (.ZN( us20_n620 ) , .A1( us20_n656 ) , .A3( us20_n666 ) , .A4( us20_n682 ) , .A2( us20_n766 ) );
  NOR2_X1 us20_U250 (.ZN( us20_n609 ) , .A2( us20_n724 ) , .A1( us20_n817 ) );
  AOI21_X1 us20_U251 (.B1( us20_n625 ) , .ZN( us20_n627 ) , .A( us20_n763 ) , .B2( us20_n814 ) );
  NOR2_X1 us20_U252 (.ZN( us20_n579 ) , .A2( us20_n708 ) , .A1( us20_n730 ) );
  NOR2_X1 us20_U253 (.ZN( us20_n533 ) , .A2( us20_n724 ) , .A1( us20_n730 ) );
  NOR2_X1 us20_U254 (.ZN( us20_n642 ) , .A2( us20_n788 ) , .A1( us20_n791 ) );
  NOR2_X1 us20_U255 (.A2( us20_n708 ) , .A1( us20_n762 ) , .ZN( us20_n794 ) );
  AOI21_X1 us20_U256 (.ZN( us20_n650 ) , .A( us20_n779 ) , .B1( us20_n792 ) , .B2( us20_n805 ) );
  AOI21_X1 us20_U257 (.A( us20_n815 ) , .B2( us20_n816 ) , .B1( us20_n817 ) , .ZN( us20_n818 ) );
  NOR2_X1 us20_U258 (.ZN( us20_n520 ) , .A2( us20_n708 ) , .A1( us20_n814 ) );
  NOR2_X1 us20_U259 (.ZN( us20_n582 ) , .A1( us20_n744 ) , .A2( us20_n815 ) );
  NOR4_X1 us20_U26 (.A4( us20_n609 ) , .A3( us20_n610 ) , .A2( us20_n611 ) , .A1( us20_n612 ) , .ZN( us20_n619 ) );
  AOI21_X1 us20_U260 (.ZN( us20_n515 ) , .A( us20_n729 ) , .B1( us20_n750 ) , .B2( us20_n803 ) );
  AOI21_X1 us20_U261 (.ZN( us20_n626 ) , .B2( us20_n669 ) , .A( us20_n790 ) , .B1( us20_n791 ) );
  AOI21_X1 us20_U262 (.ZN( us20_n499 ) , .B1( us20_n680 ) , .A( us20_n812 ) , .B2( us20_n816 ) );
  AOI21_X1 us20_U263 (.ZN( us20_n477 ) , .A( us20_n669 ) , .B1( us20_n750 ) , .B2( us20_n806 ) );
  NOR2_X1 us20_U264 (.ZN( us20_n559 ) , .A2( us20_n791 ) , .A1( us20_n803 ) );
  AOI21_X1 us20_U265 (.ZN( us20_n510 ) , .B2( us20_n669 ) , .A( us20_n730 ) , .B1( us20_n815 ) );
  NOR2_X1 us20_U266 (.ZN( us20_n519 ) , .A2( us20_n699 ) , .A1( us20_n816 ) );
  NOR2_X1 us20_U267 (.ZN( us20_n683 ) , .A2( us20_n699 ) , .A1( us20_n803 ) );
  NOR2_X1 us20_U268 (.ZN( us20_n581 ) , .A1( us20_n669 ) , .A2( us20_n788 ) );
  AOI21_X1 us20_U269 (.ZN( us20_n589 ) , .B2( us20_n699 ) , .B1( us20_n815 ) , .A( us20_n817 ) );
  NOR4_X1 us20_U27 (.A4( us20_n614 ) , .A3( us20_n615 ) , .A2( us20_n616 ) , .A1( us20_n617 ) , .ZN( us20_n618 ) );
  INV_X1 us20_U270 (.A( us20_n763 ) , .ZN( us20_n866 ) );
  AOI21_X1 us20_U271 (.ZN( us20_n498 ) , .A( us20_n724 ) , .B2( us20_n762 ) , .B1( us20_n814 ) );
  AOI21_X1 us20_U272 (.ZN( us20_n539 ) , .B2( us20_n812 ) , .A( us20_n814 ) , .B1( us20_n815 ) );
  AOI21_X1 us20_U273 (.ZN( us20_n540 ) , .A( us20_n763 ) , .B2( us20_n779 ) , .B1( us20_n817 ) );
  AOI21_X1 us20_U274 (.B1( us20_n699 ) , .ZN( us20_n700 ) , .A( us20_n732 ) , .B2( us20_n763 ) );
  AOI21_X1 us20_U275 (.ZN( us20_n591 ) , .B2( us20_n763 ) , .A( us20_n785 ) , .B1( us20_n812 ) );
  AOI21_X1 us20_U276 (.A( us20_n812 ) , .B2( us20_n813 ) , .B1( us20_n814 ) , .ZN( us20_n819 ) );
  INV_X1 us20_U277 (.A( us20_n791 ) , .ZN( us20_n873 ) );
  NOR2_X1 us20_U278 (.ZN( us20_n547 ) , .A1( us20_n699 ) , .A2( us20_n744 ) );
  INV_X1 us20_U279 (.A( us20_n729 ) , .ZN( us20_n868 ) );
  NOR4_X1 us20_U28 (.A4( us20_n514 ) , .A3( us20_n515 ) , .A2( us20_n516 ) , .A1( us20_n517 ) , .ZN( us20_n524 ) );
  AOI21_X1 us20_U280 (.ZN( us20_n569 ) , .B1( us20_n750 ) , .B2( us20_n762 ) , .A( us20_n780 ) );
  AOI21_X1 us20_U281 (.ZN( us20_n649 ) , .B1( us20_n729 ) , .B2( us20_n763 ) , .A( us20_n813 ) );
  NOR2_X1 us20_U282 (.ZN( us20_n685 ) , .A1( us20_n729 ) , .A2( us20_n816 ) );
  AOI21_X1 us20_U283 (.B1( us20_n686 ) , .ZN( us20_n687 ) , .A( us20_n728 ) , .B2( us20_n761 ) );
  AOI21_X1 us20_U284 (.ZN( us20_n640 ) , .B2( us20_n747 ) , .A( us20_n792 ) , .B1( us20_n803 ) );
  NOR2_X1 us20_U285 (.ZN( us20_n568 ) , .A1( us20_n729 ) , .A2( us20_n762 ) );
  AOI21_X1 us20_U286 (.ZN( us20_n593 ) , .B1( us20_n750 ) , .A( us20_n792 ) , .B2( us20_n813 ) );
  AOI21_X1 us20_U287 (.ZN( us20_n514 ) , .A( us20_n779 ) , .B2( us20_n792 ) , .B1( us20_n812 ) );
  INV_X1 us20_U288 (.A( us20_n699 ) , .ZN( us20_n853 ) );
  AOI21_X1 us20_U289 (.ZN( us20_n450 ) , .B2( us20_n792 ) , .A( us20_n803 ) , .B1( us20_n815 ) );
  AOI222_X1 us20_U29 (.ZN( us20_n525 ) , .A1( us20_n834 ) , .B2( us20_n837 ) , .C1( us20_n844 ) , .C2( us20_n850 ) , .A2( us20_n852 ) , .B1( us20_n866 ) );
  AOI21_X1 us20_U290 (.ZN( us20_n639 ) , .B2( us20_n749 ) , .A( us20_n788 ) , .B1( us20_n812 ) );
  AOI21_X1 us20_U291 (.ZN( us20_n564 ) , .B1( us20_n724 ) , .A( us20_n779 ) , .B2( us20_n791 ) );
  AOI21_X1 us20_U292 (.ZN( us20_n689 ) , .B2( us20_n749 ) , .B1( us20_n763 ) , .A( us20_n806 ) );
  NOR2_X1 us20_U293 (.ZN( us20_n529 ) , .A1( us20_n708 ) , .A2( us20_n779 ) );
  NOR2_X1 us20_U294 (.ZN( us20_n567 ) , .A1( us20_n747 ) , .A2( us20_n805 ) );
  AOI21_X1 us20_U295 (.A( us20_n790 ) , .B2( us20_n791 ) , .B1( us20_n792 ) , .ZN( us20_n793 ) );
  AOI21_X1 us20_U296 (.A( us20_n733 ) , .ZN( us20_n734 ) , .B2( us20_n780 ) , .B1( us20_n792 ) );
  NOR2_X1 us20_U297 (.A2( us20_n813 ) , .A1( us20_n815 ) , .ZN( us20_n821 ) );
  AOI21_X1 us20_U298 (.ZN( us20_n641 ) , .B1( us20_n680 ) , .A( us20_n791 ) , .B2( us20_n817 ) );
  NOR2_X1 us20_U299 (.ZN( us20_n578 ) , .A1( us20_n708 ) , .A2( us20_n813 ) );
  NAND4_X1 us20_U3 (.ZN( sa22_sr_2 ) , .A4( us20_n643 ) , .A3( us20_n644 ) , .A2( us20_n645 ) , .A1( us20_n646 ) );
  NOR4_X1 us20_U30 (.A3( us20_n521 ) , .A1( us20_n522 ) , .ZN( us20_n523 ) , .A2( us20_n673 ) , .A4( us20_n769 ) );
  NOR2_X1 us20_U300 (.ZN( us20_n665 ) , .A1( us20_n780 ) , .A2( us20_n813 ) );
  NOR2_X1 us20_U301 (.ZN( us20_n711 ) , .A1( us20_n762 ) , .A2( us20_n763 ) );
  NOR2_X1 us20_U302 (.ZN( us20_n583 ) , .A1( us20_n792 ) , .A2( us20_n817 ) );
  NOR2_X1 us20_U303 (.ZN( us20_n682 ) , .A2( us20_n708 ) , .A1( us20_n817 ) );
  NOR2_X1 us20_U304 (.ZN( us20_n534 ) , .A1( us20_n724 ) , .A2( us20_n788 ) );
  NOR2_X1 us20_U305 (.ZN( us20_n684 ) , .A1( us20_n791 ) , .A2( us20_n813 ) );
  NAND2_X1 us20_U306 (.ZN( us20_n753 ) , .A1( us20_n763 ) , .A2( us20_n805 ) );
  INV_X1 us20_U307 (.A( us20_n815 ) , .ZN( us20_n855 ) );
  AOI21_X1 us20_U308 (.ZN( us20_n442 ) , .A( us20_n699 ) , .B1( us20_n733 ) , .B2( us20_n750 ) );
  OAI21_X1 us20_U309 (.A( us20_n731 ) , .B1( us20_n732 ) , .ZN( us20_n736 ) , .B2( us20_n805 ) );
  AOI221_X1 us20_U31 (.A( us20_n781 ) , .ZN( us20_n798 ) , .C2( us20_n837 ) , .B2( us20_n838 ) , .B1( us20_n865 ) , .C1( us20_n866 ) );
  OAI21_X1 us20_U310 (.ZN( us20_n731 ) , .A( us20_n833 ) , .B2( us20_n852 ) , .B1( us20_n873 ) );
  INV_X1 us20_U311 (.A( us20_n780 ) , .ZN( us20_n850 ) );
  AOI21_X1 us20_U312 (.ZN( us20_n443 ) , .B1( us20_n789 ) , .B2( us20_n791 ) , .A( us20_n814 ) );
  NAND2_X1 us20_U313 (.ZN( us20_n714 ) , .A1( us20_n728 ) , .A2( us20_n780 ) );
  NAND2_X1 us20_U314 (.A2( us20_n762 ) , .A1( us20_n806 ) , .ZN( us20_n810 ) );
  INV_X1 us20_U315 (.A( us20_n785 ) , .ZN( us20_n846 ) );
  NOR2_X1 us20_U316 (.ZN( us20_n484 ) , .A1( us20_n788 ) , .A2( us20_n805 ) );
  AOI21_X1 us20_U317 (.ZN( us20_n497 ) , .A( us20_n779 ) , .B2( us20_n791 ) , .B1( us20_n804 ) );
  NOR2_X1 us20_U318 (.ZN( us20_n470 ) , .A2( us20_n779 ) , .A1( us20_n815 ) );
  NOR2_X1 us20_U319 (.ZN( us20_n712 ) , .A2( us20_n724 ) , .A1( us20_n790 ) );
  NOR4_X1 us20_U32 (.A4( us20_n793 ) , .A3( us20_n794 ) , .A2( us20_n795 ) , .A1( us20_n796 ) , .ZN( us20_n797 ) );
  NOR2_X1 us20_U320 (.ZN( us20_n526 ) , .A1( us20_n724 ) , .A2( us20_n750 ) );
  OAI21_X1 us20_U321 (.A( us20_n787 ) , .B2( us20_n788 ) , .B1( us20_n789 ) , .ZN( us20_n795 ) );
  OAI21_X1 us20_U322 (.ZN( us20_n787 ) , .A( us20_n839 ) , .B1( us20_n863 ) , .B2( us20_n873 ) );
  NAND2_X1 us20_U323 (.A1( us20_n699 ) , .A2( us20_n729 ) , .ZN( us20_n782 ) );
  NOR2_X1 us20_U324 (.ZN( us20_n518 ) , .A1( us20_n708 ) , .A2( us20_n788 ) );
  INV_X1 us20_U325 (.A( us20_n813 ) , .ZN( us20_n836 ) );
  NAND2_X1 us20_U326 (.ZN( us20_n671 ) , .A1( us20_n806 ) , .A2( us20_n816 ) );
  OAI21_X1 us20_U327 (.A( us20_n698 ) , .ZN( us20_n702 ) , .B2( us20_n750 ) , .B1( us20_n804 ) );
  OAI21_X1 us20_U328 (.ZN( us20_n698 ) , .B2( us20_n833 ) , .B1( us20_n838 ) , .A( us20_n860 ) );
  INV_X1 us20_U329 (.A( us20_n724 ) , .ZN( us20_n856 ) );
  NOR4_X1 us20_U33 (.A4( us20_n776 ) , .A3( us20_n777 ) , .A1( us20_n778 ) , .ZN( us20_n799 ) , .A2( us20_n801 ) );
  INV_X1 us20_U330 (.A( us20_n817 ) , .ZN( us20_n844 ) );
  AND2_X1 us20_U331 (.ZN( us20_n732 ) , .A1( us20_n779 ) , .A2( us20_n785 ) );
  OAI222_X1 us20_U332 (.ZN( us20_n617 ) , .B1( us20_n697 ) , .C1( us20_n724 ) , .C2( us20_n747 ) , .B2( us20_n786 ) , .A2( us20_n792 ) , .A1( us20_n816 ) );
  AOI221_X1 us20_U333 (.A( us20_n764 ) , .ZN( us20_n774 ) , .C2( us20_n810 ) , .B2( us20_n835 ) , .C1( us20_n855 ) , .B1( us20_n866 ) );
  AOI21_X1 us20_U334 (.B2( us20_n763 ) , .ZN( us20_n764 ) , .A( us20_n788 ) , .B1( us20_n792 ) );
  INV_X1 us20_U335 (.A( us20_n761 ) , .ZN( us20_n835 ) );
  NAND2_X1 us20_U336 (.A1( us20_n451 ) , .A2( us20_n454 ) , .ZN( us20_n814 ) );
  NAND2_X1 us20_U337 (.A1( us20_n447 ) , .A2( us20_n449 ) , .ZN( us20_n805 ) );
  NAND2_X1 us20_U338 (.A1( us20_n455 ) , .A2( us20_n462 ) , .ZN( us20_n750 ) );
  NAND2_X1 us20_U339 (.A1( us20_n455 ) , .A2( us20_n471 ) , .ZN( us20_n803 ) );
  NOR4_X1 us20_U34 (.A4( us20_n734 ) , .A3( us20_n735 ) , .A2( us20_n736 ) , .A1( us20_n737 ) , .ZN( us20_n738 ) );
  NAND2_X1 us20_U340 (.A1( us20_n453 ) , .A2( us20_n461 ) , .ZN( us20_n744 ) );
  NAND2_X1 us20_U341 (.A1( us20_n452 ) , .A2( us20_n465 ) , .ZN( us20_n669 ) );
  NAND2_X1 us20_U342 (.A2( us20_n448 ) , .A1( us20_n460 ) , .ZN( us20_n728 ) );
  NAND2_X1 us20_U343 (.A2( us20_n453 ) , .A1( us20_n455 ) , .ZN( us20_n806 ) );
  NAND2_X1 us20_U344 (.A1( us20_n451 ) , .A2( us20_n471 ) , .ZN( us20_n816 ) );
  NAND2_X1 us20_U345 (.A1( us20_n453 ) , .A2( us20_n472 ) , .ZN( us20_n785 ) );
  NAND2_X1 us20_U346 (.A2( us20_n454 ) , .A1( us20_n472 ) , .ZN( us20_n779 ) );
  NAND2_X1 us20_U347 (.A2( us20_n464 ) , .A1( us20_n465 ) , .ZN( us20_n812 ) );
  NAND2_X1 us20_U348 (.A1( us20_n441 ) , .A2( us20_n460 ) , .ZN( us20_n699 ) );
  NAND2_X1 us20_U349 (.A2( us20_n449 ) , .A1( us20_n452 ) , .ZN( us20_n763 ) );
  AOI211_X1 us20_U35 (.B( us20_n725 ) , .A( us20_n726 ) , .ZN( us20_n739 ) , .C1( us20_n843 ) , .C2( us20_n855 ) );
  NAND2_X1 us20_U350 (.A2( us20_n448 ) , .A1( us20_n452 ) , .ZN( us20_n729 ) );
  NAND2_X1 us20_U351 (.A2( us20_n461 ) , .A1( us20_n462 ) , .ZN( us20_n747 ) );
  NAND2_X1 us20_U352 (.A1( us20_n462 ) , .A2( us20_n472 ) , .ZN( us20_n788 ) );
  NOR2_X1 us20_U353 (.ZN( us20_n465 ) , .A2( us20_n847 ) , .A1( us20_n848 ) );
  NOR2_X1 us20_U354 (.ZN( us20_n453 ) , .A1( us20_n826 ) , .A2( us20_n827 ) );
  NOR2_X1 us20_U355 (.ZN( us20_n451 ) , .A1( us20_n828 ) , .A2( us20_n829 ) );
  NAND2_X1 us20_U356 (.A2( us20_n461 ) , .A1( us20_n471 ) , .ZN( us20_n697 ) );
  NAND2_X1 us20_U357 (.A1( us20_n451 ) , .A2( us20_n462 ) , .ZN( us20_n790 ) );
  NAND2_X1 us20_U358 (.A2( us20_n441 ) , .A1( us20_n447 ) , .ZN( us20_n784 ) );
  NAND2_X2 us20_U359 (.A2( us20_n448 ) , .A1( us20_n464 ) , .ZN( us20_n815 ) );
  NOR3_X1 us20_U36 (.A3( us20_n722 ) , .A1( us20_n723 ) , .ZN( us20_n740 ) , .A2( us20_n741 ) );
  NAND2_X1 us20_U360 (.A2( us20_n454 ) , .A1( us20_n455 ) , .ZN( us20_n730 ) );
  NAND2_X2 us20_U361 (.A2( us20_n441 ) , .A1( us20_n452 ) , .ZN( us20_n791 ) );
  NAND2_X2 us20_U362 (.A1( us20_n449 ) , .A2( us20_n464 ) , .ZN( us20_n724 ) );
  NAND2_X2 us20_U363 (.A1( us20_n449 ) , .A2( us20_n460 ) , .ZN( us20_n792 ) );
  NAND2_X2 us20_U364 (.A1( us20_n441 ) , .A2( us20_n464 ) , .ZN( us20_n708 ) );
  NAND2_X2 us20_U365 (.A2( us20_n471 ) , .A1( us20_n472 ) , .ZN( us20_n817 ) );
  NAND2_X2 us20_U366 (.A2( us20_n460 ) , .A1( us20_n465 ) , .ZN( us20_n780 ) );
  NOR2_X1 us20_U367 (.ZN( us20_n447 ) , .A2( us20_n849 ) , .A1( us20_n858 ) );
  NAND2_X1 us20_U368 (.A1( us20_n447 ) , .A2( us20_n448 ) , .ZN( us20_n786 ) );
  NOR2_X1 us20_U369 (.A2( sa20_6 ) , .A1( sa20_7 ) , .ZN( us20_n464 ) );
  NOR4_X1 us20_U37 (.A3( us20_n755 ) , .A2( us20_n756 ) , .A1( us20_n757 ) , .ZN( us20_n758 ) , .A4( us20_n869 ) );
  NOR2_X1 us20_U370 (.A2( sa20_7 ) , .ZN( us20_n460 ) , .A1( us20_n849 ) );
  NOR2_X1 us20_U371 (.A2( sa20_4 ) , .ZN( us20_n449 ) , .A1( us20_n848 ) );
  NOR2_X1 us20_U372 (.A2( sa20_4 ) , .A1( sa20_5 ) , .ZN( us20_n441 ) );
  NOR2_X1 us20_U373 (.A2( sa20_5 ) , .ZN( us20_n448 ) , .A1( us20_n847 ) );
  NOR2_X1 us20_U374 (.A2( sa20_1 ) , .ZN( us20_n471 ) , .A1( us20_n826 ) );
  NOR2_X1 us20_U375 (.A2( sa20_2 ) , .A1( sa20_3 ) , .ZN( us20_n472 ) );
  NOR2_X1 us20_U376 (.A2( sa20_6 ) , .ZN( us20_n452 ) , .A1( us20_n858 ) );
  NOR2_X1 us20_U377 (.A2( sa20_0 ) , .A1( sa20_1 ) , .ZN( us20_n462 ) );
  NOR2_X1 us20_U378 (.A2( sa20_3 ) , .ZN( us20_n455 ) , .A1( us20_n828 ) );
  NOR2_X1 us20_U379 (.A2( sa20_2 ) , .ZN( us20_n461 ) , .A1( us20_n829 ) );
  AOI211_X1 us20_U38 (.B( us20_n745 ) , .A( us20_n746 ) , .ZN( us20_n759 ) , .C1( us20_n832 ) , .C2( us20_n853 ) );
  NOR2_X1 us20_U380 (.A2( sa20_0 ) , .ZN( us20_n454 ) , .A1( us20_n827 ) );
  INV_X1 us20_U381 (.A( sa20_4 ) , .ZN( us20_n847 ) );
  INV_X1 us20_U382 (.A( sa20_6 ) , .ZN( us20_n849 ) );
  INV_X1 us20_U383 (.A( sa20_3 ) , .ZN( us20_n829 ) );
  INV_X1 us20_U384 (.A( sa20_1 ) , .ZN( us20_n827 ) );
  INV_X1 us20_U385 (.A( sa20_2 ) , .ZN( us20_n828 ) );
  INV_X1 us20_U386 (.A( sa20_0 ) , .ZN( us20_n826 ) );
  INV_X1 us20_U387 (.A( sa20_5 ) , .ZN( us20_n848 ) );
  INV_X1 us20_U388 (.A( sa20_7 ) , .ZN( us20_n858 ) );
  NAND2_X1 us20_U389 (.A1( us20_n729 ) , .A2( us20_n784 ) , .ZN( us20_n811 ) );
  NOR3_X1 us20_U39 (.A3( us20_n741 ) , .A2( us20_n742 ) , .A1( us20_n743 ) , .ZN( us20_n760 ) );
  OAI22_X1 us20_U390 (.ZN( us20_n588 ) , .A2( us20_n747 ) , .B2( us20_n762 ) , .A1( us20_n763 ) , .B1( us20_n784 ) );
  AOI21_X1 us20_U391 (.ZN( us20_n592 ) , .B1( us20_n728 ) , .B2( us20_n784 ) , .A( us20_n790 ) );
  AOI21_X1 us20_U392 (.ZN( us20_n648 ) , .A( us20_n762 ) , .B2( us20_n784 ) , .B1( us20_n792 ) );
  AOI21_X1 us20_U393 (.ZN( us20_n623 ) , .B1( us20_n699 ) , .A( us20_n779 ) , .B2( us20_n784 ) );
  OAI22_X1 us20_U394 (.ZN( us20_n681 ) , .A1( us20_n699 ) , .A2( us20_n730 ) , .B2( us20_n784 ) , .B1( us20_n817 ) );
  OAI21_X1 us20_U395 (.A( us20_n613 ) , .ZN( us20_n616 ) , .B1( us20_n625 ) , .B2( us20_n784 ) );
  NOR2_X1 us20_U396 (.ZN( us20_n610 ) , .A1( us20_n784 ) , .A2( us20_n816 ) );
  OAI222_X1 us20_U397 (.A2( us20_n669 ) , .ZN( us20_n674 ) , .B1( us20_n747 ) , .B2( us20_n784 ) , .C2( us20_n788 ) , .C1( us20_n815 ) , .A1( us20_n817 ) );
  NOR2_X1 us20_U398 (.ZN( us20_n651 ) , .A1( us20_n784 ) , .A2( us20_n788 ) );
  NOR2_X1 us20_U399 (.ZN( us20_n553 ) , .A2( us20_n744 ) , .A1( us20_n784 ) );
  NOR3_X1 us20_U4 (.ZN( us20_n598 ) , .A1( us20_n608 ) , .A3( us20_n723 ) , .A2( us20_n742 ) );
  NOR2_X1 us20_U40 (.ZN( us20_n804 ) , .A1( us20_n854 ) , .A2( us20_n861 ) );
  INV_X1 us20_U400 (.A( us20_n784 ) , .ZN( us20_n861 ) );
  INV_X1 us20_U401 (.A( us20_n697 ) , .ZN( us20_n838 ) );
  NOR2_X1 us20_U402 (.A1( us20_n697 ) , .ZN( us20_n770 ) , .A2( us20_n815 ) );
  AOI21_X1 us20_U403 (.ZN( us20_n571 ) , .B2( us20_n697 ) , .B1( us20_n806 ) , .A( us20_n812 ) );
  NOR2_X1 us20_U404 (.ZN( us20_n632 ) , .A2( us20_n697 ) , .A1( us20_n724 ) );
  AOI21_X1 us20_U405 (.ZN( us20_n478 ) , .B2( us20_n697 ) , .A( us20_n749 ) , .B1( us20_n779 ) );
  NOR2_X1 us20_U406 (.ZN( us20_n662 ) , .A2( us20_n697 ) , .A1( us20_n729 ) );
  NOR2_X1 us20_U407 (.A2( us20_n697 ) , .A1( us20_n780 ) , .ZN( us20_n820 ) );
  NOR2_X1 us20_U408 (.ZN( us20_n600 ) , .A2( us20_n697 ) , .A1( us20_n784 ) );
  NOR2_X1 us20_U409 (.A2( us20_n697 ) , .ZN( us20_n716 ) , .A1( us20_n792 ) );
  NAND4_X1 us20_U41 (.ZN( sa22_sr_3 ) , .A4( us20_n704 ) , .A3( us20_n705 ) , .A2( us20_n706 ) , .A1( us20_n707 ) );
  NOR2_X1 us20_U410 (.ZN( us20_n566 ) , .A2( us20_n697 ) , .A1( us20_n763 ) );
  NOR2_X1 us20_U411 (.ZN( us20_n594 ) , .A2( us20_n697 ) , .A1( us20_n728 ) );
  AOI21_X1 us20_U412 (.ZN( us20_n552 ) , .B1( us20_n669 ) , .A( us20_n697 ) , .B2( us20_n805 ) );
  NOR2_X1 us20_U413 (.ZN( us20_n541 ) , .A2( us20_n697 ) , .A1( us20_n699 ) );
  NOR2_X1 us20_U414 (.ZN( us20_n580 ) , .A2( us20_n697 ) , .A1( us20_n791 ) );
  NAND2_X1 us20_U415 (.A1( us20_n454 ) , .A2( us20_n461 ) , .ZN( us20_n813 ) );
  AND2_X1 us20_U416 (.ZN( us20_n438 ) , .A2( us20_n831 ) , .A1( us20_n854 ) );
  AND2_X1 us20_U417 (.ZN( us20_n439 ) , .A2( us20_n843 ) , .A1( us20_n861 ) );
  NOR3_X1 us20_U418 (.A1( us20_n438 ) , .A2( us20_n439 ) , .A3( us20_n576 ) , .ZN( us20_n587 ) );
  INV_X1 us20_U419 (.A( us20_n812 ) , .ZN( us20_n854 ) );
  NOR4_X1 us20_U42 (.A4( us20_n700 ) , .A3( us20_n701 ) , .A2( us20_n702 ) , .A1( us20_n703 ) , .ZN( us20_n704 ) );
  INV_X1 us20_U420 (.A( us20_n816 ) , .ZN( us20_n831 ) );
  INV_X1 us20_U421 (.A( us20_n803 ) , .ZN( us20_n843 ) );
  AOI21_X1 us20_U422 (.ZN( us20_n576 ) , .B2( us20_n724 ) , .B1( us20_n748 ) , .A( us20_n785 ) );
  OAI221_X1 us20_U423 (.A( us20_n783 ) , .C2( us20_n784 ) , .B2( us20_n785 ) , .B1( us20_n786 ) , .ZN( us20_n796 ) , .C1( us20_n813 ) );
  AOI21_X1 us20_U424 (.ZN( us20_n500 ) , .A( us20_n697 ) , .B1( us20_n708 ) , .B2( us20_n786 ) );
  OAI221_X1 us20_U425 (.A( us20_n696 ) , .ZN( us20_n703 ) , .C2( us20_n784 ) , .C1( us20_n785 ) , .B1( us20_n786 ) , .B2( us20_n806 ) );
  OAI22_X1 us20_U426 (.ZN( us20_n590 ) , .B1( us20_n730 ) , .B2( us20_n749 ) , .A2( us20_n786 ) , .A1( us20_n803 ) );
  AOI222_X1 us20_U427 (.ZN( us20_n605 ) , .B2( us20_n671 ) , .B1( us20_n753 ) , .C2( us20_n831 ) , .A1( us20_n833 ) , .A2( us20_n862 ) , .C1( us20_n863 ) );
  AOI222_X1 us20_U428 (.ZN( us20_n513 ) , .C1( us20_n832 ) , .B2( us20_n837 ) , .A2( us20_n843 ) , .C2( us20_n862 ) , .B1( us20_n863 ) , .A1( us20_n866 ) );
  AOI221_X1 us20_U429 (.A( us20_n483 ) , .ZN( us20_n488 ) , .B1( us20_n831 ) , .C2( us20_n844 ) , .C1( us20_n852 ) , .B2( us20_n862 ) );
  AOI211_X1 us20_U43 (.B( us20_n694 ) , .A( us20_n695 ) , .ZN( us20_n705 ) , .C2( us20_n831 ) , .C1( us20_n851 ) );
  NAND2_X1 us20_U430 (.A2( us20_n749 ) , .A1( us20_n786 ) , .ZN( us20_n809 ) );
  NOR2_X1 us20_U431 (.ZN( us20_n612 ) , .A1( us20_n779 ) , .A2( us20_n786 ) );
  NOR2_X1 us20_U432 (.ZN( us20_n717 ) , .A2( us20_n744 ) , .A1( us20_n786 ) );
  NOR2_X1 us20_U433 (.ZN( us20_n653 ) , .A1( us20_n762 ) , .A2( us20_n786 ) );
  NOR2_X1 us20_U434 (.ZN( us20_n554 ) , .A1( us20_n786 ) , .A2( us20_n813 ) );
  NOR2_X1 us20_U435 (.ZN( us20_n789 ) , .A2( us20_n862 ) , .A1( us20_n868 ) );
  NOR2_X1 us20_U436 (.ZN( us20_n701 ) , .A2( us20_n786 ) , .A1( us20_n817 ) );
  NAND3_X1 us20_U437 (.ZN( sa22_sr_6 ) , .A3( us20_n797 ) , .A2( us20_n798 ) , .A1( us20_n799 ) );
  NAND3_X1 us20_U438 (.ZN( sa22_sr_5 ) , .A3( us20_n758 ) , .A2( us20_n759 ) , .A1( us20_n760 ) );
  NAND3_X1 us20_U439 (.ZN( sa22_sr_4 ) , .A3( us20_n738 ) , .A2( us20_n739 ) , .A1( us20_n740 ) );
  NOR2_X1 us20_U44 (.ZN( us20_n707 ) , .A2( us20_n776 ) , .A1( us20_n800 ) );
  NAND3_X1 us20_U440 (.A3( us20_n675 ) , .A2( us20_n676 ) , .A1( us20_n677 ) , .ZN( us20_n807 ) );
  NAND3_X1 us20_U441 (.ZN( us20_n638 ) , .A3( us20_n708 ) , .A2( us20_n724 ) , .A1( us20_n792 ) );
  NAND3_X1 us20_U442 (.A3( us20_n618 ) , .A2( us20_n619 ) , .A1( us20_n620 ) , .ZN( us20_n725 ) );
  NAND3_X1 us20_U443 (.A3( us20_n585 ) , .A2( us20_n586 ) , .A1( us20_n587 ) , .ZN( us20_n621 ) );
  NAND3_X1 us20_U444 (.ZN( us20_n565 ) , .A3( us20_n680 ) , .A2( us20_n750 ) , .A1( us20_n785 ) );
  NAND3_X1 us20_U445 (.A3( us20_n523 ) , .A2( us20_n524 ) , .A1( us20_n525 ) , .ZN( us20_n742 ) );
  NAND3_X1 us20_U446 (.A3( us20_n512 ) , .A1( us20_n513 ) , .ZN( us20_n608 ) , .A2( us20_n871 ) );
  NAND3_X1 us20_U447 (.A3( us20_n467 ) , .A2( us20_n468 ) , .A1( us20_n469 ) , .ZN( us20_n777 ) );
  NOR2_X1 us20_U448 (.A1( us20_n730 ) , .ZN( us20_n765 ) , .A2( us20_n786 ) );
  INV_X1 us20_U449 (.A( us20_n786 ) , .ZN( us20_n862 ) );
  NAND4_X1 us20_U45 (.ZN( sa22_sr_7 ) , .A4( us20_n822 ) , .A3( us20_n823 ) , .A2( us20_n824 ) , .A1( us20_n825 ) );
  NOR4_X1 us20_U46 (.A4( us20_n818 ) , .A3( us20_n819 ) , .A2( us20_n820 ) , .A1( us20_n821 ) , .ZN( us20_n822 ) );
  AOI222_X1 us20_U47 (.C2( us20_n809 ) , .B2( us20_n810 ) , .A2( us20_n811 ) , .ZN( us20_n823 ) , .C1( us20_n832 ) , .A1( us20_n839 ) , .B1( us20_n853 ) );
  AOI211_X1 us20_U48 (.B( us20_n807 ) , .A( us20_n808 ) , .ZN( us20_n824 ) , .C1( us20_n842 ) , .C2( us20_n850 ) );
  NAND4_X1 us20_U49 (.ZN( sa22_sr_0 ) , .A4( us20_n501 ) , .A3( us20_n502 ) , .A2( us20_n503 ) , .A1( us20_n504 ) );
  NOR3_X1 us20_U5 (.A3( us20_n800 ) , .A2( us20_n801 ) , .A1( us20_n802 ) , .ZN( us20_n825 ) );
  NOR4_X1 us20_U50 (.A4( us20_n498 ) , .A3( us20_n499 ) , .A2( us20_n500 ) , .ZN( us20_n501 ) , .A1( us20_n527 ) );
  AOI221_X1 us20_U51 (.A( us20_n497 ) , .ZN( us20_n502 ) , .B2( us20_n843 ) , .C1( us20_n846 ) , .C2( us20_n860 ) , .B1( us20_n862 ) );
  AOI211_X1 us20_U52 (.A( us20_n496 ) , .ZN( us20_n503 ) , .B( us20_n802 ) , .C2( us20_n839 ) , .C1( us20_n851 ) );
  NAND4_X1 us20_U53 (.ZN( sa22_sr_1 ) , .A4( us20_n595 ) , .A3( us20_n596 ) , .A2( us20_n597 ) , .A1( us20_n598 ) );
  NOR4_X1 us20_U54 (.A4( us20_n591 ) , .A3( us20_n592 ) , .A2( us20_n593 ) , .A1( us20_n594 ) , .ZN( us20_n595 ) );
  AOI211_X1 us20_U55 (.B( us20_n589 ) , .A( us20_n590 ) , .ZN( us20_n596 ) , .C2( us20_n811 ) , .C1( us20_n833 ) );
  AOI211_X1 us20_U56 (.A( us20_n588 ) , .ZN( us20_n597 ) , .B( us20_n621 ) , .C1( us20_n845 ) , .C2( us20_n855 ) );
  NOR2_X1 us20_U57 (.ZN( us20_n748 ) , .A1( us20_n861 ) , .A2( us20_n862 ) );
  NOR2_X1 us20_U58 (.ZN( us20_n625 ) , .A2( us20_n836 ) , .A1( us20_n839 ) );
  AOI222_X1 us20_U59 (.B2( us20_n638 ) , .ZN( us20_n644 ) , .B1( us20_n841 ) , .A1( us20_n842 ) , .C2( us20_n846 ) , .C1( us20_n863 ) , .A2( us20_n865 ) );
  NOR3_X1 us20_U6 (.A3( us20_n621 ) , .A2( us20_n622 ) , .ZN( us20_n636 ) , .A1( us20_n725 ) );
  NOR4_X1 us20_U60 (.A4( us20_n639 ) , .A3( us20_n640 ) , .A2( us20_n641 ) , .A1( us20_n642 ) , .ZN( us20_n643 ) );
  NOR3_X1 us20_U61 (.A2( us20_n607 ) , .A1( us20_n608 ) , .ZN( us20_n646 ) , .A3( us20_n722 ) );
  NAND4_X1 us20_U62 (.A4( us20_n603 ) , .A3( us20_n604 ) , .A2( us20_n605 ) , .A1( us20_n606 ) , .ZN( us20_n722 ) );
  NOR3_X1 us20_U63 (.A1( us20_n599 ) , .ZN( us20_n604 ) , .A3( us20_n663 ) , .A2( us20_n770 ) );
  NOR4_X1 us20_U64 (.A3( us20_n600 ) , .A2( us20_n601 ) , .A1( us20_n602 ) , .ZN( us20_n603 ) , .A4( us20_n655 ) );
  AOI222_X1 us20_U65 (.ZN( us20_n606 ) , .A1( us20_n830 ) , .C2( us20_n837 ) , .B1( us20_n842 ) , .A2( us20_n856 ) , .B2( us20_n861 ) , .C1( us20_n868 ) );
  AOI222_X1 us20_U66 (.ZN( us20_n469 ) , .B1( us20_n832 ) , .A1( us20_n839 ) , .C1( us20_n842 ) , .C2( us20_n851 ) , .A2( us20_n855 ) , .B2( us20_n865 ) );
  NOR4_X1 us20_U67 (.A1( us20_n466 ) , .ZN( us20_n467 ) , .A4( us20_n542 ) , .A2( us20_n554 ) , .A3( us20_n614 ) );
  AOI221_X1 us20_U68 (.ZN( us20_n468 ) , .C2( us20_n714 ) , .B2( us20_n831 ) , .C1( us20_n845 ) , .B1( us20_n860 ) , .A( us20_n864 ) );
  NAND4_X1 us20_U69 (.A4( us20_n485 ) , .A3( us20_n486 ) , .A2( us20_n487 ) , .A1( us20_n488 ) , .ZN( us20_n778 ) );
  NOR2_X1 us20_U7 (.ZN( us20_n495 ) , .A1( us20_n678 ) , .A2( us20_n694 ) );
  NOR4_X1 us20_U70 (.A4( us20_n484 ) , .ZN( us20_n487 ) , .A1( us20_n566 ) , .A2( us20_n581 ) , .A3( us20_n602 ) );
  NOR4_X1 us20_U71 (.ZN( us20_n486 ) , .A1( us20_n507 ) , .A2( us20_n519 ) , .A4( us20_n546 ) , .A3( us20_n611 ) );
  NOR4_X1 us20_U72 (.ZN( us20_n485 ) , .A2( us20_n533 ) , .A1( us20_n558 ) , .A3( us20_n631 ) , .A4( us20_n718 ) );
  NAND4_X1 us20_U73 (.A4( us20_n657 ) , .A3( us20_n658 ) , .A2( us20_n659 ) , .A1( us20_n660 ) , .ZN( us20_n800 ) );
  NOR3_X1 us20_U74 (.A3( us20_n648 ) , .A2( us20_n649 ) , .A1( us20_n650 ) , .ZN( us20_n659 ) );
  NOR3_X1 us20_U75 (.A3( us20_n651 ) , .A2( us20_n652 ) , .A1( us20_n653 ) , .ZN( us20_n658 ) );
  NOR3_X1 us20_U76 (.A3( us20_n654 ) , .A2( us20_n655 ) , .A1( us20_n656 ) , .ZN( us20_n657 ) );
  NAND4_X1 us20_U77 (.A4( us20_n560 ) , .A3( us20_n561 ) , .A2( us20_n562 ) , .A1( us20_n563 ) , .ZN( us20_n607 ) );
  NOR4_X1 us20_U78 (.A4( us20_n552 ) , .A3( us20_n553 ) , .A2( us20_n554 ) , .A1( us20_n555 ) , .ZN( us20_n562 ) );
  NOR4_X1 us20_U79 (.ZN( us20_n561 ) , .A1( us20_n653 ) , .A3( us20_n661 ) , .A4( us20_n685 ) , .A2( us20_n768 ) );
  NOR2_X1 us20_U8 (.A1( us20_n678 ) , .ZN( us20_n693 ) , .A2( us20_n807 ) );
  NOR4_X1 us20_U80 (.A4( us20_n556 ) , .A3( us20_n557 ) , .A2( us20_n558 ) , .A1( us20_n559 ) , .ZN( us20_n560 ) );
  NAND4_X1 us20_U81 (.A4( us20_n772 ) , .A3( us20_n773 ) , .A2( us20_n774 ) , .A1( us20_n775 ) , .ZN( us20_n801 ) );
  NOR3_X1 us20_U82 (.A3( us20_n765 ) , .A2( us20_n766 ) , .A1( us20_n767 ) , .ZN( us20_n773 ) );
  NOR4_X1 us20_U83 (.A4( us20_n768 ) , .A3( us20_n769 ) , .A2( us20_n770 ) , .A1( us20_n771 ) , .ZN( us20_n772 ) );
  AOI222_X1 us20_U84 (.ZN( us20_n775 ) , .A1( us20_n830 ) , .C1( us20_n834 ) , .B2( us20_n841 ) , .A2( us20_n850 ) , .B1( us20_n861 ) , .C2( us20_n873 ) );
  NOR4_X1 us20_U85 (.A4( us20_n509 ) , .A2( us20_n510 ) , .A1( us20_n511 ) , .ZN( us20_n512 ) , .A3( us20_n670 ) );
  INV_X1 us20_U86 (.A( us20_n505 ) , .ZN( us20_n871 ) );
  NOR4_X1 us20_U87 (.A4( us20_n661 ) , .A3( us20_n662 ) , .A2( us20_n663 ) , .A1( us20_n664 ) , .ZN( us20_n677 ) );
  NOR4_X1 us20_U88 (.A4( us20_n665 ) , .A3( us20_n666 ) , .A2( us20_n667 ) , .A1( us20_n668 ) , .ZN( us20_n676 ) );
  NOR4_X1 us20_U89 (.A3( us20_n673 ) , .A1( us20_n674 ) , .ZN( us20_n675 ) , .A4( us20_n715 ) , .A2( us20_n859 ) );
  NOR3_X1 us20_U9 (.ZN( us20_n504 ) , .A2( us20_n679 ) , .A3( us20_n777 ) , .A1( us20_n876 ) );
  NOR2_X1 us20_U90 (.ZN( us20_n761 ) , .A1( us20_n833 ) , .A2( us20_n834 ) );
  NOR2_X1 us20_U91 (.ZN( us20_n686 ) , .A1( us20_n831 ) , .A2( us20_n832 ) );
  NOR4_X1 us20_U92 (.A4( us20_n577 ) , .A3( us20_n578 ) , .A2( us20_n579 ) , .ZN( us20_n586 ) , .A1( us20_n683 ) );
  NOR4_X1 us20_U93 (.A1( us20_n584 ) , .ZN( us20_n585 ) , .A3( us20_n652 ) , .A2( us20_n662 ) , .A4( us20_n767 ) );
  NAND4_X1 us20_U94 (.A4( us20_n456 ) , .A3( us20_n457 ) , .A2( us20_n458 ) , .A1( us20_n459 ) , .ZN( us20_n679 ) );
  NOR3_X1 us20_U95 (.ZN( us20_n457 ) , .A3( us20_n530 ) , .A1( us20_n555 ) , .A2( us20_n570 ) );
  AOI221_X1 us20_U96 (.A( us20_n450 ) , .ZN( us20_n459 ) , .C2( us20_n753 ) , .B1( us20_n832 ) , .C1( us20_n842 ) , .B2( us20_n861 ) );
  NOR4_X1 us20_U97 (.ZN( us20_n458 ) , .A2( us20_n509 ) , .A1( us20_n599 ) , .A4( us20_n628 ) , .A3( us20_n711 ) );
  NAND4_X1 us20_U98 (.A4( us20_n535 ) , .A3( us20_n536 ) , .A2( us20_n537 ) , .A1( us20_n538 ) , .ZN( us20_n622 ) );
  NOR4_X1 us20_U99 (.A4( us20_n526 ) , .A2( us20_n527 ) , .A1( us20_n528 ) , .ZN( us20_n538 ) , .A3( us20_n701 ) );
  INV_X1 us23_U10 (.A( us23_n679 ) , .ZN( us23_n839 ) );
  NOR4_X1 us23_U100 (.A4( us23_n483 ) , .ZN( us23_n486 ) , .A1( us23_n565 ) , .A2( us23_n580 ) , .A3( us23_n601 ) );
  NOR4_X1 us23_U101 (.ZN( us23_n485 ) , .A1( us23_n506 ) , .A2( us23_n518 ) , .A4( us23_n545 ) , .A3( us23_n610 ) );
  NOR4_X1 us23_U102 (.ZN( us23_n484 ) , .A2( us23_n532 ) , .A1( us23_n557 ) , .A3( us23_n630 ) , .A4( us23_n717 ) );
  NAND4_X1 us23_U103 (.A4( us23_n690 ) , .A3( us23_n691 ) , .A1( us23_n692 ) , .ZN( us23_n775 ) , .A2( us23_n871 ) );
  AOI221_X1 us23_U104 (.A( us23_n680 ) , .ZN( us23_n691 ) , .B2( us23_n839 ) , .C1( us23_n841 ) , .C2( us23_n861 ) , .B1( us23_n864 ) );
  INV_X1 us23_U105 (.A( us23_n678 ) , .ZN( us23_n871 ) );
  NOR4_X1 us23_U106 (.A4( us23_n686 ) , .A3( us23_n687 ) , .A2( us23_n688 ) , .A1( us23_n689 ) , .ZN( us23_n690 ) );
  NAND4_X1 us23_U107 (.A4( us23_n559 ) , .A3( us23_n560 ) , .A2( us23_n561 ) , .A1( us23_n562 ) , .ZN( us23_n606 ) );
  NOR4_X1 us23_U108 (.ZN( us23_n560 ) , .A1( us23_n652 ) , .A3( us23_n660 ) , .A4( us23_n684 ) , .A2( us23_n767 ) );
  NOR4_X1 us23_U109 (.A4( us23_n551 ) , .A3( us23_n552 ) , .A2( us23_n553 ) , .A1( us23_n554 ) , .ZN( us23_n561 ) );
  NOR4_X1 us23_U11 (.A4( us23_n444 ) , .A3( us23_n445 ) , .A2( us23_n515 ) , .A1( us23_n540 ) , .ZN( us23_n705 ) );
  NOR4_X1 us23_U110 (.A4( us23_n555 ) , .A3( us23_n556 ) , .A2( us23_n557 ) , .A1( us23_n558 ) , .ZN( us23_n559 ) );
  NAND4_X1 us23_U111 (.A4( us23_n718 ) , .A3( us23_n719 ) , .A2( us23_n720 ) , .ZN( us23_n740 ) , .A1( us23_n856 ) );
  INV_X1 us23_U112 (.A( us23_n708 ) , .ZN( us23_n856 ) );
  AOI221_X1 us23_U113 (.A( us23_n709 ) , .ZN( us23_n720 ) , .C2( us23_n843 ) , .B2( us23_n844 ) , .C1( us23_n860 ) , .B1( us23_n861 ) );
  NOR4_X1 us23_U114 (.A4( us23_n714 ) , .A3( us23_n715 ) , .A2( us23_n716 ) , .A1( us23_n717 ) , .ZN( us23_n718 ) );
  NAND4_X1 us23_U115 (.A4( us23_n472 ) , .A3( us23_n473 ) , .A2( us23_n474 ) , .A1( us23_n475 ) , .ZN( us23_n677 ) );
  NOR4_X1 us23_U116 (.A4( us23_n469 ) , .ZN( us23_n475 ) , .A3( us23_n555 ) , .A1( us23_n734 ) , .A2( us23_n754 ) );
  NOR4_X1 us23_U117 (.ZN( us23_n474 ) , .A1( us23_n530 ) , .A3( us23_n567 ) , .A4( us23_n599 ) , .A2( us23_n641 ) );
  NOR4_X1 us23_U118 (.ZN( us23_n473 ) , .A1( us23_n505 ) , .A3( us23_n543 ) , .A2( us23_n582 ) , .A4( us23_n715 ) );
  NOR2_X1 us23_U119 (.ZN( us23_n732 ) , .A2( us23_n831 ) , .A1( us23_n844 ) );
  OR3_X1 us23_U12 (.ZN( us23_n445 ) , .A1( us23_n527 ) , .A3( us23_n576 ) , .A2( us23_n874 ) );
  NOR2_X1 us23_U120 (.ZN( us23_n788 ) , .A2( us23_n861 ) , .A1( us23_n867 ) );
  NAND4_X1 us23_U121 (.A4( us23_n572 ) , .A3( us23_n573 ) , .A1( us23_n574 ) , .ZN( us23_n722 ) , .A2( us23_n873 ) );
  NOR4_X1 us23_U122 (.A4( us23_n568 ) , .A3( us23_n569 ) , .A2( us23_n570 ) , .A1( us23_n571 ) , .ZN( us23_n572 ) );
  AOI221_X1 us23_U123 (.A( us23_n563 ) , .C2( us23_n564 ) , .ZN( us23_n573 ) , .B2( us23_n844 ) , .B1( us23_n851 ) , .C1( us23_n852 ) );
  INV_X1 us23_U124 (.A( us23_n606 ) , .ZN( us23_n873 ) );
  NAND4_X1 us23_U125 (.A4( us23_n492 ) , .A3( us23_n493 ) , .A1( us23_n494 ) , .ZN( us23_n801 ) , .A2( us23_n866 ) );
  AOI221_X1 us23_U126 (.A( us23_n488 ) , .ZN( us23_n493 ) , .B2( us23_n835 ) , .C2( us23_n840 ) , .C1( us23_n850 ) , .B1( us23_n859 ) );
  INV_X1 us23_U127 (.A( us23_n777 ) , .ZN( us23_n866 ) );
  NOR2_X1 us23_U128 (.ZN( us23_n494 ) , .A1( us23_n677 ) , .A2( us23_n693 ) );
  NOR2_X1 us23_U129 (.ZN( us23_n747 ) , .A1( us23_n860 ) , .A2( us23_n861 ) );
  OR4_X1 us23_U13 (.A4( us23_n441 ) , .A2( us23_n442 ) , .A1( us23_n443 ) , .ZN( us23_n444 ) , .A3( us23_n552 ) );
  AOI222_X1 us23_U130 (.ZN( us23_n512 ) , .C1( us23_n831 ) , .B2( us23_n836 ) , .A2( us23_n842 ) , .C2( us23_n861 ) , .B1( us23_n862 ) , .A1( us23_n865 ) );
  NOR4_X1 us23_U131 (.A4( us23_n508 ) , .A2( us23_n509 ) , .A1( us23_n510 ) , .ZN( us23_n511 ) , .A3( us23_n669 ) );
  INV_X1 us23_U132 (.A( us23_n504 ) , .ZN( us23_n870 ) );
  INV_X1 us23_U133 (.A( us23_n761 ) , .ZN( us23_n829 ) );
  NOR2_X1 us23_U134 (.ZN( us23_n646 ) , .A1( us23_n853 ) , .A2( us23_n867 ) );
  OR4_X1 us23_U135 (.A4( us23_n579 ) , .A3( us23_n580 ) , .A2( us23_n581 ) , .A1( us23_n582 ) , .ZN( us23_n583 ) );
  OR4_X1 us23_U136 (.A4( us23_n681 ) , .A3( us23_n682 ) , .A2( us23_n683 ) , .A1( us23_n684 ) , .ZN( us23_n689 ) );
  OR4_X1 us23_U137 (.A4( us23_n565 ) , .A3( us23_n566 ) , .A2( us23_n567 ) , .ZN( us23_n571 ) , .A1( us23_n664 ) );
  OR4_X1 us23_U138 (.A4( us23_n517 ) , .A2( us23_n518 ) , .A1( us23_n519 ) , .ZN( us23_n521 ) , .A3( us23_n820 ) );
  OR4_X1 us23_U139 (.ZN( us23_n465 ) , .A4( us23_n517 ) , .A3( us23_n528 ) , .A2( us23_n577 ) , .A1( us23_n711 ) );
  INV_X1 us23_U14 (.A( us23_n612 ) , .ZN( us23_n874 ) );
  NAND2_X1 us23_U140 (.ZN( us23_n612 ) , .A2( us23_n836 ) , .A1( us23_n872 ) );
  OR3_X1 us23_U141 (.A3( us23_n505 ) , .A2( us23_n506 ) , .A1( us23_n507 ) , .ZN( us23_n510 ) );
  AOI221_X1 us23_U142 (.A( us23_n712 ) , .B2( us23_n713 ) , .ZN( us23_n719 ) , .C1( us23_n831 ) , .B1( us23_n838 ) , .C2( us23_n862 ) );
  OR2_X1 us23_U143 (.A2( us23_n710 ) , .A1( us23_n711 ) , .ZN( us23_n712 ) );
  INV_X1 us23_U144 (.A( us23_n462 ) , .ZN( us23_n863 ) );
  OAI21_X1 us23_U145 (.ZN( us23_n462 ) , .B1( us23_n808 ) , .A( us23_n833 ) , .B2( us23_n850 ) );
  INV_X1 us23_U146 (.A( us23_n753 ) , .ZN( us23_n868 ) );
  OAI21_X1 us23_U147 (.B1( us23_n752 ) , .ZN( us23_n753 ) , .A( us23_n844 ) , .B2( us23_n867 ) );
  INV_X1 us23_U148 (.A( us23_n671 ) , .ZN( us23_n858 ) );
  AOI21_X1 us23_U149 (.A( us23_n669 ) , .B1( us23_n670 ) , .ZN( us23_n671 ) , .B2( us23_n855 ) );
  INV_X1 us23_U15 (.A( us23_n748 ) , .ZN( us23_n862 ) );
  AOI222_X1 us23_U150 (.ZN( us23_n659 ) , .A2( us23_n838 ) , .B1( us23_n840 ) , .C2( us23_n844 ) , .A1( us23_n859 ) , .C1( us23_n862 ) , .B2( us23_n869 ) );
  INV_X1 us23_U151 (.A( us23_n646 ) , .ZN( us23_n869 ) );
  OAI222_X1 us23_U152 (.B2( us23_n707 ) , .ZN( us23_n708 ) , .C2( us23_n723 ) , .B1( us23_n746 ) , .A1( us23_n805 ) , .C1( us23_n813 ) , .A2( us23_n814 ) );
  OAI222_X1 us23_U153 (.A2( us23_n668 ) , .ZN( us23_n673 ) , .B1( us23_n746 ) , .B2( us23_n783 ) , .C2( us23_n787 ) , .C1( us23_n814 ) , .A1( us23_n816 ) );
  NAND2_X1 us23_U154 (.A1( us23_n446 ) , .A2( us23_n464 ) , .ZN( us23_n748 ) );
  NOR4_X1 us23_U155 (.A2( us23_n490 ) , .A1( us23_n491 ) , .ZN( us23_n492 ) , .A3( us23_n579 ) , .A4( us23_n611 ) );
  OR4_X1 us23_U156 (.ZN( us23_n491 ) , .A4( us23_n533 ) , .A2( us23_n546 ) , .A1( us23_n558 ) , .A3( us23_n631 ) );
  OAI22_X1 us23_U157 (.B1( us23_n489 ) , .ZN( us23_n490 ) , .A1( us23_n685 ) , .A2( us23_n762 ) , .B2( us23_n816 ) );
  NOR3_X1 us23_U158 (.ZN( us23_n489 ) , .A1( us23_n781 ) , .A2( us23_n849 ) , .A3( us23_n862 ) );
  AOI22_X1 us23_U159 (.ZN( us23_n695 ) , .A1( us23_n829 ) , .B2( us23_n842 ) , .A2( us23_n864 ) , .B1( us23_n867 ) );
  AOI222_X1 us23_U16 (.ZN( us23_n604 ) , .B2( us23_n670 ) , .B1( us23_n752 ) , .C2( us23_n830 ) , .A1( us23_n832 ) , .A2( us23_n861 ) , .C1( us23_n862 ) );
  AOI21_X1 us23_U160 (.ZN( us23_n638 ) , .B2( us23_n748 ) , .A( us23_n787 ) , .B1( us23_n811 ) );
  AOI21_X1 us23_U161 (.ZN( us23_n639 ) , .B2( us23_n746 ) , .A( us23_n791 ) , .B1( us23_n802 ) );
  AOI21_X1 us23_U162 (.ZN( us23_n640 ) , .B1( us23_n679 ) , .A( us23_n790 ) , .B2( us23_n816 ) );
  INV_X1 us23_U163 (.A( us23_n729 ) , .ZN( us23_n838 ) );
  AOI221_X1 us23_U164 (.A( us23_n763 ) , .ZN( us23_n773 ) , .C2( us23_n809 ) , .B2( us23_n834 ) , .C1( us23_n854 ) , .B1( us23_n865 ) );
  AOI21_X1 us23_U165 (.B2( us23_n762 ) , .ZN( us23_n763 ) , .A( us23_n787 ) , .B1( us23_n791 ) );
  INV_X1 us23_U166 (.A( us23_n760 ) , .ZN( us23_n834 ) );
  AOI221_X1 us23_U167 (.A( us23_n449 ) , .ZN( us23_n458 ) , .C2( us23_n752 ) , .B1( us23_n831 ) , .C1( us23_n841 ) , .B2( us23_n860 ) );
  AOI21_X1 us23_U168 (.ZN( us23_n449 ) , .B2( us23_n791 ) , .A( us23_n802 ) , .B1( us23_n814 ) );
  AOI221_X1 us23_U169 (.A( us23_n482 ) , .ZN( us23_n487 ) , .B1( us23_n830 ) , .C2( us23_n843 ) , .C1( us23_n851 ) , .B2( us23_n861 ) );
  AOI222_X1 us23_U17 (.ZN( us23_n562 ) , .B1( us23_n829 ) , .C1( us23_n840 ) , .A2( us23_n842 ) , .A1( us23_n853 ) , .B2( us23_n862 ) , .C2( us23_n872 ) );
  OAI22_X1 us23_U170 (.ZN( us23_n482 ) , .A1( us23_n707 ) , .B2( us23_n784 ) , .A2( us23_n805 ) , .B1( us23_n811 ) );
  INV_X1 us23_U171 (.A( us23_n789 ) , .ZN( us23_n831 ) );
  NAND2_X1 us23_U172 (.A1( us23_n450 ) , .A2( us23_n452 ) , .ZN( us23_n761 ) );
  INV_X1 us23_U173 (.A( us23_n783 ) , .ZN( us23_n860 ) );
  INV_X1 us23_U174 (.A( us23_n785 ) , .ZN( us23_n861 ) );
  INV_X1 us23_U175 (.A( us23_n815 ) , .ZN( us23_n830 ) );
  OAI22_X1 us23_U176 (.ZN( us23_n709 ) , .A2( us23_n727 ) , .B2( us23_n728 ) , .A1( us23_n743 ) , .B1( us23_n812 ) );
  OAI22_X1 us23_U177 (.ZN( us23_n623 ) , .B1( us23_n668 ) , .B2( us23_n746 ) , .A1( us23_n814 ) , .A2( us23_n815 ) );
  OAI22_X1 us23_U178 (.ZN( us23_n587 ) , .A2( us23_n746 ) , .B2( us23_n761 ) , .A1( us23_n762 ) , .B1( us23_n783 ) );
  INV_X1 us23_U179 (.A( us23_n743 ) , .ZN( us23_n836 ) );
  NOR4_X1 us23_U18 (.ZN( us23_n472 ) , .A2( us23_n520 ) , .A4( us23_n593 ) , .A1( us23_n608 ) , .A3( us23_n628 ) );
  INV_X1 us23_U180 (.A( us23_n787 ) , .ZN( us23_n844 ) );
  OAI22_X1 us23_U181 (.A1( us23_n723 ) , .ZN( us23_n725 ) , .B2( us23_n749 ) , .B1( us23_n811 ) , .A2( us23_n815 ) );
  OAI22_X1 us23_U182 (.B2( us23_n778 ) , .B1( us23_n779 ) , .ZN( us23_n780 ) , .A2( us23_n813 ) , .A1( us23_n814 ) );
  OAI22_X1 us23_U183 (.ZN( us23_n680 ) , .A1( us23_n698 ) , .A2( us23_n729 ) , .B2( us23_n783 ) , .B1( us23_n816 ) );
  OAI22_X1 us23_U184 (.B2( us23_n749 ) , .B1( us23_n750 ) , .A1( us23_n751 ) , .ZN( us23_n755 ) , .A2( us23_n805 ) );
  NOR2_X1 us23_U185 (.ZN( us23_n750 ) , .A2( us23_n851 ) , .A1( us23_n859 ) );
  NOR3_X1 us23_U186 (.ZN( us23_n751 ) , .A2( us23_n852 ) , .A1( us23_n862 ) , .A3( us23_n864 ) );
  OAI22_X1 us23_U187 (.B2( us23_n743 ) , .ZN( us23_n745 ) , .A2( us23_n761 ) , .B1( us23_n779 ) , .A1( us23_n791 ) );
  INV_X1 us23_U188 (.A( us23_n802 ) , .ZN( us23_n842 ) );
  INV_X1 us23_U189 (.A( us23_n813 ) , .ZN( us23_n832 ) );
  NOR4_X1 us23_U19 (.A4( us23_n531 ) , .A3( us23_n532 ) , .A2( us23_n533 ) , .ZN( us23_n534 ) , .A1( us23_n819 ) );
  INV_X1 us23_U190 (.A( us23_n804 ) , .ZN( us23_n859 ) );
  OAI22_X1 us23_U191 (.B2( us23_n802 ) , .B1( us23_n803 ) , .A2( us23_n804 ) , .A1( us23_n805 ) , .ZN( us23_n807 ) );
  OAI22_X1 us23_U192 (.ZN( us23_n495 ) , .A2( us23_n743 ) , .A1( us23_n779 ) , .B1( us23_n790 ) , .B2( us23_n805 ) );
  OAI22_X1 us23_U193 (.ZN( us23_n488 ) , .A1( us23_n723 ) , .B2( us23_n727 ) , .B1( us23_n729 ) , .A2( us23_n778 ) );
  INV_X1 us23_U194 (.A( us23_n668 ) , .ZN( us23_n864 ) );
  OAI22_X1 us23_U195 (.ZN( us23_n694 ) , .A2( us23_n729 ) , .A1( us23_n779 ) , .B1( us23_n790 ) , .B2( us23_n816 ) );
  OAI22_X1 us23_U196 (.ZN( us23_n636 ) , .A1( us23_n698 ) , .B2( us23_n727 ) , .A2( us23_n761 ) , .B1( us23_n815 ) );
  NOR2_X1 us23_U197 (.A1( us23_n696 ) , .ZN( us23_n769 ) , .A2( us23_n814 ) );
  NOR2_X1 us23_U198 (.ZN( us23_n714 ) , .A1( us23_n804 ) , .A2( us23_n816 ) );
  NOR2_X1 us23_U199 (.ZN( us23_n717 ) , .A2( us23_n723 ) , .A1( us23_n743 ) );
  NOR4_X1 us23_U20 (.ZN( us23_n478 ) , .A1( us23_n519 ) , .A4( us23_n556 ) , .A3( us23_n581 ) , .A2( us23_n629 ) );
  NOR2_X1 us23_U200 (.ZN( us23_n545 ) , .A2( us23_n779 ) , .A1( us23_n813 ) );
  INV_X1 us23_U201 (.A( us23_n749 ) , .ZN( us23_n841 ) );
  NOR2_X1 us23_U202 (.ZN( us23_n651 ) , .A1( us23_n668 ) , .A2( us23_n813 ) );
  NOR2_X1 us23_U203 (.ZN( us23_n531 ) , .A2( us23_n748 ) , .A1( us23_n749 ) );
  NOR2_X1 us23_U204 (.ZN( us23_n576 ) , .A2( us23_n698 ) , .A1( us23_n813 ) );
  NOR2_X1 us23_U205 (.ZN( us23_n599 ) , .A2( us23_n696 ) , .A1( us23_n783 ) );
  NOR2_X1 us23_U206 (.A1( us23_n668 ) , .ZN( us23_n672 ) , .A2( us23_n743 ) );
  NOR2_X1 us23_U207 (.ZN( us23_n601 ) , .A1( us23_n668 ) , .A2( us23_n802 ) );
  NOR2_X1 us23_U208 (.A1( us23_n668 ) , .ZN( us23_n687 ) , .A2( us23_n815 ) );
  NOR2_X1 us23_U209 (.ZN( us23_n628 ) , .A2( us23_n727 ) , .A1( us23_n784 ) );
  NOR4_X1 us23_U21 (.A4( us23_n540 ) , .A3( us23_n541 ) , .A2( us23_n542 ) , .ZN( us23_n549 ) , .A1( us23_n687 ) );
  NOR2_X1 us23_U210 (.ZN( us23_n614 ) , .A1( us23_n784 ) , .A2( us23_n814 ) );
  NOR2_X1 us23_U211 (.A2( us23_n743 ) , .ZN( us23_n754 ) , .A1( us23_n804 ) );
  NOR2_X1 us23_U212 (.A1( us23_n668 ) , .ZN( us23_n765 ) , .A2( us23_n812 ) );
  NOR2_X1 us23_U213 (.ZN( us23_n734 ) , .A2( us23_n802 ) , .A1( us23_n804 ) );
  NOR2_X1 us23_U214 (.A1( us23_n698 ) , .ZN( us23_n767 ) , .A2( us23_n812 ) );
  NOR2_X1 us23_U215 (.A2( us23_n743 ) , .ZN( us23_n768 ) , .A1( us23_n811 ) );
  NOR2_X1 us23_U216 (.ZN( us23_n530 ) , .A2( us23_n779 ) , .A1( us23_n815 ) );
  NOR2_X1 us23_U217 (.ZN( us23_n526 ) , .A1( us23_n668 ) , .A2( us23_n778 ) );
  NOR2_X1 us23_U218 (.ZN( us23_n540 ) , .A2( us23_n696 ) , .A1( us23_n698 ) );
  NOR2_X1 us23_U219 (.ZN( us23_n598 ) , .A2( us23_n790 ) , .A1( us23_n815 ) );
  NOR2_X1 us23_U22 (.ZN( us23_n679 ) , .A2( us23_n833 ) , .A1( us23_n838 ) );
  NOR2_X1 us23_U220 (.ZN( us23_n627 ) , .A2( us23_n668 ) , .A1( us23_n784 ) );
  NOR2_X1 us23_U221 (.ZN( us23_n600 ) , .A2( us23_n779 ) , .A1( us23_n802 ) );
  INV_X1 us23_U222 (.A( us23_n746 ) , .ZN( us23_n833 ) );
  NOR2_X1 us23_U223 (.ZN( us23_n610 ) , .A2( us23_n779 ) , .A1( us23_n805 ) );
  NOR2_X1 us23_U224 (.ZN( us23_n527 ) , .A2( us23_n723 ) , .A1( us23_n802 ) );
  NOR2_X1 us23_U225 (.ZN( us23_n609 ) , .A1( us23_n783 ) , .A2( us23_n815 ) );
  INV_X1 us23_U226 (.A( us23_n791 ) , .ZN( us23_n850 ) );
  NOR2_X1 us23_U227 (.ZN( us23_n650 ) , .A1( us23_n783 ) , .A2( us23_n787 ) );
  NOR2_X1 us23_U228 (.A2( us23_n707 ) , .A1( us23_n749 ) , .ZN( us23_n770 ) );
  NOR2_X1 us23_U229 (.ZN( us23_n666 ) , .A1( us23_n749 ) , .A2( us23_n814 ) );
  AOI222_X1 us23_U23 (.ZN( us23_n468 ) , .B1( us23_n831 ) , .A1( us23_n838 ) , .C1( us23_n841 ) , .C2( us23_n850 ) , .A2( us23_n854 ) , .B2( us23_n864 ) );
  NOR2_X1 us23_U230 (.ZN( us23_n554 ) , .A1( us23_n749 ) , .A2( us23_n790 ) );
  NOR2_X1 us23_U231 (.ZN( us23_n507 ) , .A2( us23_n779 ) , .A1( us23_n784 ) );
  NOR2_X1 us23_U232 (.ZN( us23_n542 ) , .A2( us23_n707 ) , .A1( us23_n784 ) );
  NOR2_X1 us23_U233 (.ZN( us23_n663 ) , .A1( us23_n784 ) , .A2( us23_n790 ) );
  OAI22_X1 us23_U234 (.B1( us23_n439 ) , .ZN( us23_n443 ) , .A2( us23_n727 ) , .A1( us23_n743 ) , .B2( us23_n748 ) );
  NOR3_X1 us23_U235 (.ZN( us23_n439 ) , .A2( us23_n835 ) , .A3( us23_n836 ) , .A1( us23_n845 ) );
  NOR2_X1 us23_U236 (.A2( us23_n696 ) , .ZN( us23_n715 ) , .A1( us23_n791 ) );
  NOR2_X1 us23_U237 (.ZN( us23_n506 ) , .A1( us23_n811 ) , .A2( us23_n816 ) );
  NOR2_X1 us23_U238 (.ZN( us23_n593 ) , .A2( us23_n696 ) , .A1( us23_n727 ) );
  NOR2_X1 us23_U239 (.ZN( us23_n661 ) , .A2( us23_n696 ) , .A1( us23_n728 ) );
  NOR4_X1 us23_U24 (.A1( us23_n465 ) , .ZN( us23_n466 ) , .A4( us23_n541 ) , .A2( us23_n553 ) , .A3( us23_n613 ) );
  NOR2_X1 us23_U240 (.ZN( us23_n556 ) , .A1( us23_n791 ) , .A2( us23_n813 ) );
  NOR2_X1 us23_U241 (.ZN( us23_n544 ) , .A1( us23_n748 ) , .A2( us23_n813 ) );
  NOR2_X1 us23_U242 (.ZN( us23_n555 ) , .A1( us23_n761 ) , .A2( us23_n804 ) );
  NOR2_X1 us23_U243 (.ZN( us23_n529 ) , .A2( us23_n743 ) , .A1( us23_n791 ) );
  NOR2_X1 us23_U244 (.A2( us23_n696 ) , .A1( us23_n779 ) , .ZN( us23_n819 ) );
  NOR2_X1 us23_U245 (.ZN( us23_n508 ) , .A1( us23_n728 ) , .A2( us23_n778 ) );
  NOR2_X1 us23_U246 (.ZN( us23_n665 ) , .A1( us23_n727 ) , .A2( us23_n802 ) );
  NOR2_X1 us23_U247 (.ZN( us23_n543 ) , .A2( us23_n784 ) , .A1( us23_n791 ) );
  NOR2_X1 us23_U248 (.A1( us23_n748 ) , .ZN( us23_n766 ) , .A2( us23_n802 ) );
  NOR2_X1 us23_U249 (.ZN( us23_n613 ) , .A1( us23_n761 ) , .A2( us23_n811 ) );
  AOI221_X1 us23_U25 (.ZN( us23_n467 ) , .C2( us23_n713 ) , .B2( us23_n830 ) , .C1( us23_n844 ) , .B1( us23_n859 ) , .A( us23_n863 ) );
  NOR2_X1 us23_U250 (.ZN( us23_n515 ) , .A1( us23_n707 ) , .A2( us23_n743 ) );
  NOR2_X1 us23_U251 (.ZN( us23_n630 ) , .A1( us23_n723 ) , .A2( us23_n812 ) );
  NOR2_X1 us23_U252 (.ZN( us23_n569 ) , .A1( us23_n727 ) , .A2( us23_n805 ) );
  NOR2_X1 us23_U253 (.ZN( us23_n557 ) , .A1( us23_n707 ) , .A2( us23_n815 ) );
  INV_X1 us23_U254 (.A( us23_n762 ) , .ZN( us23_n865 ) );
  NOR2_X1 us23_U255 (.ZN( us23_n653 ) , .A1( us23_n727 ) , .A2( us23_n812 ) );
  NOR2_X1 us23_U256 (.ZN( us23_n516 ) , .A1( us23_n707 ) , .A2( us23_n802 ) );
  NOR2_X1 us23_U257 (.ZN( us23_n520 ) , .A1( us23_n789 ) , .A2( us23_n811 ) );
  NOR2_X1 us23_U258 (.ZN( us23_n662 ) , .A1( us23_n728 ) , .A2( us23_n784 ) );
  NOR2_X1 us23_U259 (.ZN( us23_n654 ) , .A1( us23_n789 ) , .A2( us23_n814 ) );
  NOR4_X1 us23_U26 (.A4( us23_n664 ) , .A3( us23_n665 ) , .A2( us23_n666 ) , .A1( us23_n667 ) , .ZN( us23_n675 ) );
  NOR2_X1 us23_U260 (.ZN( us23_n629 ) , .A1( us23_n746 ) , .A2( us23_n814 ) );
  NOR2_X1 us23_U261 (.ZN( us23_n667 ) , .A2( us23_n707 ) , .A1( us23_n789 ) );
  NOR2_X1 us23_U262 (.ZN( us23_n669 ) , .A1( us23_n789 ) , .A2( us23_n804 ) );
  AOI21_X1 us23_U263 (.ZN( us23_n570 ) , .B2( us23_n696 ) , .B1( us23_n805 ) , .A( us23_n811 ) );
  NOR2_X1 us23_U264 (.ZN( us23_n541 ) , .A1( us23_n761 ) , .A2( us23_n790 ) );
  NOR2_X1 us23_U265 (.ZN( us23_n655 ) , .A1( us23_n746 ) , .A2( us23_n779 ) );
  INV_X1 us23_U266 (.A( us23_n805 ) , .ZN( us23_n840 ) );
  NOR2_X1 us23_U267 (.ZN( us23_n608 ) , .A2( us23_n723 ) , .A1( us23_n816 ) );
  AOI21_X1 us23_U268 (.A( us23_n814 ) , .B2( us23_n815 ) , .B1( us23_n816 ) , .ZN( us23_n817 ) );
  AOI21_X1 us23_U269 (.ZN( us23_n625 ) , .B2( us23_n668 ) , .A( us23_n789 ) , .B1( us23_n790 ) );
  NOR4_X1 us23_U27 (.A4( us23_n660 ) , .A3( us23_n661 ) , .A2( us23_n662 ) , .A1( us23_n663 ) , .ZN( us23_n676 ) );
  NOR2_X1 us23_U270 (.ZN( us23_n660 ) , .A1( us23_n728 ) , .A2( us23_n789 ) );
  INV_X1 us23_U271 (.A( us23_n811 ) , .ZN( us23_n853 ) );
  NOR2_X1 us23_U272 (.ZN( us23_n578 ) , .A2( us23_n707 ) , .A1( us23_n729 ) );
  NOR2_X1 us23_U273 (.ZN( us23_n532 ) , .A2( us23_n723 ) , .A1( us23_n729 ) );
  AOI21_X1 us23_U274 (.ZN( us23_n498 ) , .B1( us23_n679 ) , .A( us23_n811 ) , .B2( us23_n815 ) );
  AOI21_X1 us23_U275 (.ZN( us23_n551 ) , .B1( us23_n668 ) , .A( us23_n696 ) , .B2( us23_n804 ) );
  NOR2_X1 us23_U276 (.ZN( us23_n581 ) , .A1( us23_n743 ) , .A2( us23_n814 ) );
  NOR2_X1 us23_U277 (.A2( us23_n707 ) , .A1( us23_n761 ) , .ZN( us23_n793 ) );
  AOI21_X1 us23_U278 (.B1( us23_n624 ) , .ZN( us23_n626 ) , .A( us23_n762 ) , .B2( us23_n813 ) );
  AOI21_X1 us23_U279 (.ZN( us23_n514 ) , .A( us23_n728 ) , .B1( us23_n749 ) , .B2( us23_n802 ) );
  NOR4_X1 us23_U28 (.A3( us23_n672 ) , .A1( us23_n673 ) , .ZN( us23_n674 ) , .A4( us23_n714 ) , .A2( us23_n858 ) );
  AOI21_X1 us23_U280 (.A( us23_n811 ) , .B2( us23_n812 ) , .B1( us23_n813 ) , .ZN( us23_n818 ) );
  AOI21_X1 us23_U281 (.ZN( us23_n477 ) , .B2( us23_n696 ) , .A( us23_n748 ) , .B1( us23_n778 ) );
  AOI21_X1 us23_U282 (.ZN( us23_n509 ) , .B2( us23_n668 ) , .A( us23_n729 ) , .B1( us23_n814 ) );
  NOR2_X1 us23_U283 (.ZN( us23_n505 ) , .A2( us23_n727 ) , .A1( us23_n761 ) );
  AOI21_X1 us23_U284 (.ZN( us23_n591 ) , .B1( us23_n727 ) , .B2( us23_n783 ) , .A( us23_n789 ) );
  NOR2_X1 us23_U285 (.ZN( us23_n518 ) , .A2( us23_n698 ) , .A1( us23_n815 ) );
  AOI21_X1 us23_U286 (.ZN( us23_n592 ) , .B1( us23_n749 ) , .A( us23_n791 ) , .B2( us23_n812 ) );
  AOI21_X1 us23_U287 (.ZN( us23_n649 ) , .A( us23_n778 ) , .B1( us23_n791 ) , .B2( us23_n804 ) );
  NOR2_X1 us23_U288 (.ZN( us23_n580 ) , .A1( us23_n668 ) , .A2( us23_n787 ) );
  NOR2_X1 us23_U289 (.ZN( us23_n519 ) , .A2( us23_n707 ) , .A1( us23_n813 ) );
  NOR4_X1 us23_U29 (.A4( us23_n513 ) , .A3( us23_n514 ) , .A2( us23_n515 ) , .A1( us23_n516 ) , .ZN( us23_n523 ) );
  AOI21_X1 us23_U290 (.ZN( us23_n476 ) , .A( us23_n668 ) , .B1( us23_n749 ) , .B2( us23_n805 ) );
  NOR2_X1 us23_U291 (.ZN( us23_n558 ) , .A2( us23_n790 ) , .A1( us23_n802 ) );
  AOI21_X1 us23_U292 (.ZN( us23_n647 ) , .A( us23_n761 ) , .B2( us23_n783 ) , .B1( us23_n791 ) );
  AOI21_X1 us23_U293 (.ZN( us23_n622 ) , .B1( us23_n698 ) , .A( us23_n778 ) , .B2( us23_n783 ) );
  AOI21_X1 us23_U294 (.ZN( us23_n588 ) , .B2( us23_n698 ) , .B1( us23_n814 ) , .A( us23_n816 ) );
  NOR2_X1 us23_U295 (.ZN( us23_n552 ) , .A2( us23_n743 ) , .A1( us23_n783 ) );
  NOR2_X1 us23_U296 (.ZN( us23_n682 ) , .A2( us23_n698 ) , .A1( us23_n802 ) );
  AOI21_X1 us23_U297 (.B1( us23_n698 ) , .ZN( us23_n699 ) , .A( us23_n731 ) , .B2( us23_n762 ) );
  AOI21_X1 us23_U298 (.ZN( us23_n590 ) , .B2( us23_n762 ) , .A( us23_n784 ) , .B1( us23_n811 ) );
  AOI21_X1 us23_U299 (.ZN( us23_n538 ) , .B2( us23_n811 ) , .A( us23_n813 ) , .B1( us23_n814 ) );
  NOR3_X1 us23_U3 (.ZN( us23_n597 ) , .A1( us23_n607 ) , .A3( us23_n722 ) , .A2( us23_n741 ) );
  AOI222_X1 us23_U30 (.ZN( us23_n524 ) , .A1( us23_n833 ) , .B2( us23_n836 ) , .C1( us23_n843 ) , .C2( us23_n849 ) , .A2( us23_n851 ) , .B1( us23_n865 ) );
  AOI21_X1 us23_U300 (.ZN( us23_n539 ) , .A( us23_n762 ) , .B2( us23_n778 ) , .B1( us23_n816 ) );
  NOR2_X1 us23_U301 (.ZN( us23_n546 ) , .A1( us23_n698 ) , .A2( us23_n743 ) );
  INV_X1 us23_U302 (.A( us23_n812 ) , .ZN( us23_n835 ) );
  INV_X1 us23_U303 (.A( us23_n727 ) , .ZN( us23_n851 ) );
  AOI21_X1 us23_U304 (.ZN( us23_n648 ) , .B1( us23_n728 ) , .B2( us23_n762 ) , .A( us23_n812 ) );
  INV_X1 us23_U305 (.A( us23_n790 ) , .ZN( us23_n872 ) );
  OAI221_X1 us23_U306 (.A( us23_n726 ) , .C2( us23_n727 ) , .B2( us23_n728 ) , .B1( us23_n729 ) , .ZN( us23_n736 ) , .C1( us23_n816 ) );
  AOI22_X1 us23_U307 (.ZN( us23_n726 ) , .B1( us23_n831 ) , .A2( us23_n837 ) , .A1( us23_n862 ) , .B2( us23_n865 ) );
  AOI21_X1 us23_U308 (.ZN( us23_n497 ) , .A( us23_n723 ) , .B2( us23_n761 ) , .B1( us23_n813 ) );
  NOR2_X1 us23_U309 (.ZN( us23_n565 ) , .A2( us23_n696 ) , .A1( us23_n762 ) );
  NOR4_X1 us23_U31 (.A3( us23_n520 ) , .A1( us23_n521 ) , .ZN( us23_n522 ) , .A2( us23_n672 ) , .A4( us23_n768 ) );
  INV_X1 us23_U310 (.A( us23_n698 ) , .ZN( us23_n852 ) );
  AOI21_X1 us23_U311 (.ZN( us23_n568 ) , .B1( us23_n749 ) , .B2( us23_n761 ) , .A( us23_n779 ) );
  AOI21_X1 us23_U312 (.ZN( us23_n513 ) , .A( us23_n778 ) , .B2( us23_n791 ) , .B1( us23_n811 ) );
  NOR2_X1 us23_U313 (.ZN( us23_n579 ) , .A2( us23_n696 ) , .A1( us23_n790 ) );
  NOR2_X1 us23_U314 (.ZN( us23_n684 ) , .A1( us23_n728 ) , .A2( us23_n815 ) );
  AOI21_X1 us23_U315 (.ZN( us23_n563 ) , .B1( us23_n723 ) , .A( us23_n778 ) , .B2( us23_n790 ) );
  AOI21_X1 us23_U316 (.ZN( us23_n496 ) , .A( us23_n778 ) , .B2( us23_n790 ) , .B1( us23_n803 ) );
  INV_X1 us23_U317 (.A( us23_n728 ) , .ZN( us23_n867 ) );
  NOR2_X1 us23_U318 (.ZN( us23_n664 ) , .A1( us23_n779 ) , .A2( us23_n812 ) );
  NOR2_X1 us23_U319 (.ZN( us23_n631 ) , .A2( us23_n696 ) , .A1( us23_n723 ) );
  AOI221_X1 us23_U32 (.A( us23_n780 ) , .ZN( us23_n797 ) , .C2( us23_n836 ) , .B2( us23_n837 ) , .B1( us23_n864 ) , .C1( us23_n865 ) );
  NOR2_X1 us23_U320 (.ZN( us23_n528 ) , .A1( us23_n707 ) , .A2( us23_n778 ) );
  NOR2_X1 us23_U321 (.ZN( us23_n577 ) , .A1( us23_n707 ) , .A2( us23_n812 ) );
  AOI21_X1 us23_U322 (.A( us23_n789 ) , .B2( us23_n790 ) , .B1( us23_n791 ) , .ZN( us23_n792 ) );
  AOI21_X1 us23_U323 (.ZN( us23_n688 ) , .B2( us23_n748 ) , .B1( us23_n762 ) , .A( us23_n805 ) );
  NOR2_X1 us23_U324 (.ZN( us23_n683 ) , .A1( us23_n790 ) , .A2( us23_n812 ) );
  NOR2_X1 us23_U325 (.ZN( us23_n566 ) , .A1( us23_n746 ) , .A2( us23_n804 ) );
  NAND2_X1 us23_U326 (.ZN( us23_n752 ) , .A1( us23_n762 ) , .A2( us23_n804 ) );
  AOI21_X1 us23_U327 (.A( us23_n732 ) , .ZN( us23_n733 ) , .B2( us23_n779 ) , .B1( us23_n791 ) );
  NOR2_X1 us23_U328 (.A2( us23_n812 ) , .A1( us23_n814 ) , .ZN( us23_n820 ) );
  NOR2_X1 us23_U329 (.ZN( us23_n710 ) , .A1( us23_n761 ) , .A2( us23_n762 ) );
  NOR4_X1 us23_U33 (.A4( us23_n792 ) , .A3( us23_n793 ) , .A2( us23_n794 ) , .A1( us23_n795 ) , .ZN( us23_n796 ) );
  NOR2_X1 us23_U330 (.ZN( us23_n641 ) , .A2( us23_n787 ) , .A1( us23_n790 ) );
  NOR2_X1 us23_U331 (.ZN( us23_n582 ) , .A1( us23_n791 ) , .A2( us23_n816 ) );
  NOR2_X1 us23_U332 (.ZN( us23_n681 ) , .A2( us23_n707 ) , .A1( us23_n816 ) );
  NOR2_X1 us23_U333 (.ZN( us23_n533 ) , .A1( us23_n723 ) , .A2( us23_n787 ) );
  AOI21_X1 us23_U334 (.B1( us23_n685 ) , .ZN( us23_n686 ) , .A( us23_n727 ) , .B2( us23_n760 ) );
  INV_X1 us23_U335 (.A( us23_n696 ) , .ZN( us23_n837 ) );
  INV_X1 us23_U336 (.A( us23_n814 ) , .ZN( us23_n854 ) );
  NOR2_X1 us23_U337 (.ZN( us23_n567 ) , .A1( us23_n728 ) , .A2( us23_n761 ) );
  AOI21_X1 us23_U338 (.ZN( us23_n441 ) , .A( us23_n698 ) , .B1( us23_n732 ) , .B2( us23_n749 ) );
  OAI21_X1 us23_U339 (.A( us23_n730 ) , .B1( us23_n731 ) , .ZN( us23_n735 ) , .B2( us23_n804 ) );
  NOR4_X1 us23_U34 (.A4( us23_n775 ) , .A3( us23_n776 ) , .A1( us23_n777 ) , .ZN( us23_n798 ) , .A2( us23_n800 ) );
  OAI21_X1 us23_U340 (.ZN( us23_n730 ) , .A( us23_n832 ) , .B2( us23_n851 ) , .B1( us23_n872 ) );
  OAI21_X1 us23_U341 (.A( us23_n697 ) , .ZN( us23_n701 ) , .B2( us23_n749 ) , .B1( us23_n803 ) );
  OAI21_X1 us23_U342 (.ZN( us23_n697 ) , .B2( us23_n832 ) , .B1( us23_n837 ) , .A( us23_n859 ) );
  OAI21_X1 us23_U343 (.A( us23_n612 ) , .ZN( us23_n615 ) , .B1( us23_n624 ) , .B2( us23_n783 ) );
  INV_X1 us23_U344 (.A( us23_n779 ) , .ZN( us23_n849 ) );
  AOI22_X1 us23_U345 (.A2( us23_n781 ) , .ZN( us23_n782 ) , .B2( us23_n830 ) , .A1( us23_n833 ) , .B1( us23_n862 ) );
  NAND2_X1 us23_U346 (.ZN( us23_n670 ) , .A1( us23_n805 ) , .A2( us23_n815 ) );
  OAI21_X1 us23_U347 (.A( us23_n786 ) , .B2( us23_n787 ) , .B1( us23_n788 ) , .ZN( us23_n794 ) );
  OAI21_X1 us23_U348 (.ZN( us23_n786 ) , .A( us23_n838 ) , .B1( us23_n862 ) , .B2( us23_n872 ) );
  NAND2_X1 us23_U349 (.A1( us23_n728 ) , .A2( us23_n783 ) , .ZN( us23_n810 ) );
  NOR4_X1 us23_U35 (.A4( us23_n733 ) , .A3( us23_n734 ) , .A2( us23_n735 ) , .A1( us23_n736 ) , .ZN( us23_n737 ) );
  NOR2_X1 us23_U350 (.ZN( us23_n483 ) , .A1( us23_n787 ) , .A2( us23_n804 ) );
  AOI21_X1 us23_U351 (.ZN( us23_n442 ) , .B1( us23_n788 ) , .B2( us23_n790 ) , .A( us23_n813 ) );
  NAND2_X1 us23_U352 (.A2( us23_n761 ) , .A1( us23_n805 ) , .ZN( us23_n809 ) );
  NOR2_X1 us23_U353 (.ZN( us23_n469 ) , .A2( us23_n778 ) , .A1( us23_n814 ) );
  NAND2_X1 us23_U354 (.A1( us23_n698 ) , .A2( us23_n728 ) , .ZN( us23_n781 ) );
  NOR2_X1 us23_U355 (.ZN( us23_n711 ) , .A2( us23_n723 ) , .A1( us23_n789 ) );
  INV_X1 us23_U356 (.A( us23_n784 ) , .ZN( us23_n845 ) );
  NOR2_X1 us23_U357 (.ZN( us23_n525 ) , .A1( us23_n723 ) , .A2( us23_n749 ) );
  NOR2_X1 us23_U358 (.ZN( us23_n517 ) , .A1( us23_n707 ) , .A2( us23_n787 ) );
  INV_X1 us23_U359 (.A( us23_n816 ) , .ZN( us23_n843 ) );
  AOI211_X1 us23_U36 (.B( us23_n724 ) , .A( us23_n725 ) , .ZN( us23_n738 ) , .C1( us23_n842 ) , .C2( us23_n854 ) );
  NAND2_X1 us23_U360 (.ZN( us23_n713 ) , .A1( us23_n727 ) , .A2( us23_n779 ) );
  INV_X1 us23_U361 (.A( us23_n723 ) , .ZN( us23_n855 ) );
  AND2_X1 us23_U362 (.ZN( us23_n731 ) , .A1( us23_n778 ) , .A2( us23_n784 ) );
  NAND2_X1 us23_U363 (.A2( us23_n460 ) , .A1( us23_n470 ) , .ZN( us23_n696 ) );
  NAND2_X1 us23_U364 (.A1( us23_n451 ) , .A2( us23_n464 ) , .ZN( us23_n668 ) );
  NAND2_X1 us23_U365 (.A1( us23_n450 ) , .A2( us23_n470 ) , .ZN( us23_n815 ) );
  NAND2_X1 us23_U366 (.A1( us23_n452 ) , .A2( us23_n460 ) , .ZN( us23_n743 ) );
  NAND2_X1 us23_U367 (.A1( us23_n454 ) , .A2( us23_n470 ) , .ZN( us23_n802 ) );
  NAND2_X1 us23_U368 (.A1( us23_n450 ) , .A2( us23_n453 ) , .ZN( us23_n813 ) );
  NAND2_X1 us23_U369 (.A1( us23_n454 ) , .A2( us23_n461 ) , .ZN( us23_n749 ) );
  NOR3_X1 us23_U37 (.A3( us23_n721 ) , .A1( us23_n722 ) , .ZN( us23_n739 ) , .A2( us23_n740 ) );
  NAND2_X1 us23_U370 (.A1( us23_n446 ) , .A2( us23_n448 ) , .ZN( us23_n804 ) );
  NAND2_X1 us23_U371 (.A1( us23_n453 ) , .A2( us23_n460 ) , .ZN( us23_n812 ) );
  NAND2_X1 us23_U372 (.A2( us23_n440 ) , .A1( us23_n446 ) , .ZN( us23_n783 ) );
  NAND2_X1 us23_U373 (.A2( us23_n453 ) , .A1( us23_n471 ) , .ZN( us23_n778 ) );
  NAND2_X1 us23_U374 (.A2( us23_n452 ) , .A1( us23_n454 ) , .ZN( us23_n805 ) );
  NAND2_X1 us23_U375 (.A1( us23_n452 ) , .A2( us23_n471 ) , .ZN( us23_n784 ) );
  NAND2_X1 us23_U376 (.A1( us23_n440 ) , .A2( us23_n459 ) , .ZN( us23_n698 ) );
  NAND2_X1 us23_U377 (.A2( us23_n463 ) , .A1( us23_n464 ) , .ZN( us23_n811 ) );
  NAND2_X1 us23_U378 (.A2( us23_n448 ) , .A1( us23_n451 ) , .ZN( us23_n762 ) );
  NAND2_X1 us23_U379 (.A1( us23_n461 ) , .A2( us23_n471 ) , .ZN( us23_n787 ) );
  NOR4_X1 us23_U38 (.A3( us23_n754 ) , .A2( us23_n755 ) , .A1( us23_n756 ) , .ZN( us23_n757 ) , .A4( us23_n868 ) );
  NAND2_X1 us23_U380 (.A2( us23_n460 ) , .A1( us23_n461 ) , .ZN( us23_n746 ) );
  NOR2_X1 us23_U381 (.ZN( us23_n464 ) , .A2( us23_n846 ) , .A1( us23_n847 ) );
  NOR2_X1 us23_U382 (.ZN( us23_n452 ) , .A1( us23_n825 ) , .A2( us23_n826 ) );
  NAND2_X1 us23_U383 (.A1( us23_n450 ) , .A2( us23_n461 ) , .ZN( us23_n789 ) );
  NOR2_X1 us23_U384 (.ZN( us23_n450 ) , .A1( us23_n827 ) , .A2( us23_n828 ) );
  NAND2_X2 us23_U385 (.A2( us23_n447 ) , .A1( us23_n463 ) , .ZN( us23_n814 ) );
  NAND2_X1 us23_U386 (.A2( us23_n453 ) , .A1( us23_n454 ) , .ZN( us23_n729 ) );
  NAND2_X2 us23_U387 (.A2( us23_n440 ) , .A1( us23_n451 ) , .ZN( us23_n790 ) );
  NAND2_X2 us23_U388 (.A1( us23_n448 ) , .A2( us23_n459 ) , .ZN( us23_n791 ) );
  NAND2_X2 us23_U389 (.A1( us23_n448 ) , .A2( us23_n463 ) , .ZN( us23_n723 ) );
  AOI211_X1 us23_U39 (.B( us23_n744 ) , .A( us23_n745 ) , .ZN( us23_n758 ) , .C1( us23_n831 ) , .C2( us23_n852 ) );
  NAND2_X2 us23_U390 (.A1( us23_n440 ) , .A2( us23_n463 ) , .ZN( us23_n707 ) );
  NAND2_X2 us23_U391 (.A2( us23_n470 ) , .A1( us23_n471 ) , .ZN( us23_n816 ) );
  NAND2_X2 us23_U392 (.A2( us23_n459 ) , .A1( us23_n464 ) , .ZN( us23_n779 ) );
  NOR2_X1 us23_U393 (.ZN( us23_n446 ) , .A2( us23_n848 ) , .A1( us23_n857 ) );
  NAND2_X1 us23_U394 (.A1( us23_n446 ) , .A2( us23_n447 ) , .ZN( us23_n785 ) );
  NAND2_X1 us23_U395 (.A2( us23_n447 ) , .A1( us23_n459 ) , .ZN( us23_n727 ) );
  NAND2_X1 us23_U396 (.A2( us23_n447 ) , .A1( us23_n451 ) , .ZN( us23_n728 ) );
  NOR2_X1 us23_U397 (.A2( sa23_5 ) , .ZN( us23_n447 ) , .A1( us23_n846 ) );
  NOR2_X1 us23_U398 (.A2( sa23_7 ) , .ZN( us23_n459 ) , .A1( us23_n848 ) );
  NOR2_X1 us23_U399 (.A2( sa23_6 ) , .A1( sa23_7 ) , .ZN( us23_n463 ) );
  NOR3_X1 us23_U4 (.A3( us23_n799 ) , .A2( us23_n800 ) , .A1( us23_n801 ) , .ZN( us23_n824 ) );
  NOR3_X1 us23_U40 (.A3( us23_n740 ) , .A2( us23_n741 ) , .A1( us23_n742 ) , .ZN( us23_n759 ) );
  NOR2_X1 us23_U400 (.A2( sa23_4 ) , .ZN( us23_n448 ) , .A1( us23_n847 ) );
  NOR2_X1 us23_U401 (.A2( sa23_4 ) , .A1( sa23_5 ) , .ZN( us23_n440 ) );
  NOR2_X1 us23_U402 (.A2( sa23_6 ) , .ZN( us23_n451 ) , .A1( us23_n857 ) );
  NOR2_X1 us23_U403 (.A2( sa23_1 ) , .ZN( us23_n470 ) , .A1( us23_n825 ) );
  NOR2_X1 us23_U404 (.A2( sa23_2 ) , .A1( sa23_3 ) , .ZN( us23_n471 ) );
  NOR2_X1 us23_U405 (.A2( sa23_2 ) , .ZN( us23_n460 ) , .A1( us23_n828 ) );
  NOR2_X1 us23_U406 (.A2( sa23_0 ) , .ZN( us23_n453 ) , .A1( us23_n826 ) );
  NOR2_X1 us23_U407 (.A2( sa23_0 ) , .A1( sa23_1 ) , .ZN( us23_n461 ) );
  NOR2_X1 us23_U408 (.A2( sa23_3 ) , .ZN( us23_n454 ) , .A1( us23_n827 ) );
  INV_X1 us23_U409 (.A( sa23_6 ) , .ZN( us23_n848 ) );
  NAND4_X1 us23_U41 (.ZN( sa21_sr_3 ) , .A4( us23_n703 ) , .A3( us23_n704 ) , .A2( us23_n705 ) , .A1( us23_n706 ) );
  INV_X1 us23_U410 (.A( sa23_4 ) , .ZN( us23_n846 ) );
  INV_X1 us23_U411 (.A( sa23_1 ) , .ZN( us23_n826 ) );
  INV_X1 us23_U412 (.A( sa23_3 ) , .ZN( us23_n828 ) );
  INV_X1 us23_U413 (.A( sa23_2 ) , .ZN( us23_n827 ) );
  INV_X1 us23_U414 (.A( sa23_0 ) , .ZN( us23_n825 ) );
  INV_X1 us23_U415 (.A( sa23_7 ) , .ZN( us23_n857 ) );
  INV_X1 us23_U416 (.A( sa23_5 ) , .ZN( us23_n847 ) );
  OAI221_X1 us23_U417 (.A( us23_n782 ) , .C2( us23_n783 ) , .B2( us23_n784 ) , .B1( us23_n785 ) , .ZN( us23_n795 ) , .C1( us23_n812 ) );
  OAI222_X1 us23_U418 (.B2( us23_n746 ) , .B1( us23_n747 ) , .A2( us23_n748 ) , .ZN( us23_n756 ) , .C2( us23_n804 ) , .C1( us23_n813 ) , .A1( us23_n816 ) );
  AOI21_X1 us23_U419 (.ZN( us23_n499 ) , .A( us23_n696 ) , .B1( us23_n707 ) , .B2( us23_n785 ) );
  NOR4_X1 us23_U42 (.A4( us23_n699 ) , .A3( us23_n700 ) , .A2( us23_n701 ) , .A1( us23_n702 ) , .ZN( us23_n703 ) );
  OAI221_X1 us23_U420 (.A( us23_n695 ) , .ZN( us23_n702 ) , .C2( us23_n783 ) , .C1( us23_n784 ) , .B1( us23_n785 ) , .B2( us23_n805 ) );
  OAI22_X1 us23_U421 (.ZN( us23_n589 ) , .B1( us23_n729 ) , .B2( us23_n748 ) , .A2( us23_n785 ) , .A1( us23_n802 ) );
  OAI222_X1 us23_U422 (.ZN( us23_n504 ) , .C2( us23_n624 ) , .B2( us23_n646 ) , .B1( us23_n746 ) , .A2( us23_n747 ) , .C1( us23_n804 ) , .A1( us23_n805 ) );
  NOR2_X1 us23_U423 (.ZN( us23_n611 ) , .A1( us23_n778 ) , .A2( us23_n785 ) );
  OAI222_X1 us23_U424 (.ZN( us23_n616 ) , .B1( us23_n696 ) , .C1( us23_n723 ) , .C2( us23_n746 ) , .B2( us23_n785 ) , .A2( us23_n791 ) , .A1( us23_n815 ) );
  NAND2_X1 us23_U425 (.A2( us23_n748 ) , .A1( us23_n785 ) , .ZN( us23_n808 ) );
  AOI21_X1 us23_U426 (.ZN( us23_n575 ) , .B2( us23_n723 ) , .B1( us23_n747 ) , .A( us23_n784 ) );
  NOR2_X1 us23_U427 (.ZN( us23_n716 ) , .A2( us23_n743 ) , .A1( us23_n785 ) );
  NOR2_X1 us23_U428 (.ZN( us23_n652 ) , .A1( us23_n761 ) , .A2( us23_n785 ) );
  NOR2_X1 us23_U429 (.ZN( us23_n553 ) , .A1( us23_n785 ) , .A2( us23_n812 ) );
  AOI211_X1 us23_U43 (.B( us23_n693 ) , .A( us23_n694 ) , .ZN( us23_n704 ) , .C2( us23_n830 ) , .C1( us23_n850 ) );
  NOR2_X1 us23_U430 (.ZN( us23_n700 ) , .A2( us23_n785 ) , .A1( us23_n816 ) );
  NOR2_X1 us23_U431 (.A1( us23_n729 ) , .ZN( us23_n764 ) , .A2( us23_n785 ) );
  NAND2_X1 us23_U432 (.ZN( sa21_sr_2 ) , .A1( us23_n438 ) , .A2( us23_n644 ) );
  NOR3_X1 us23_U433 (.A2( us23_n606 ) , .A1( us23_n607 ) , .ZN( us23_n645 ) , .A3( us23_n721 ) );
  AOI222_X1 us23_U434 (.B2( us23_n637 ) , .ZN( us23_n643 ) , .B1( us23_n840 ) , .A1( us23_n841 ) , .C2( us23_n845 ) , .C1( us23_n862 ) , .A2( us23_n864 ) );
  NOR4_X1 us23_U435 (.A4( us23_n638 ) , .A3( us23_n639 ) , .A2( us23_n640 ) , .A1( us23_n641 ) , .ZN( us23_n642 ) );
  AOI211_X1 us23_U436 (.A( us23_n636 ) , .ZN( us23_n644 ) , .B( us23_n742 ) , .C2( us23_n838 ) , .C1( us23_n853 ) );
  NAND3_X1 us23_U437 (.ZN( sa21_sr_6 ) , .A3( us23_n796 ) , .A2( us23_n797 ) , .A1( us23_n798 ) );
  NAND3_X1 us23_U438 (.ZN( sa21_sr_5 ) , .A3( us23_n757 ) , .A2( us23_n758 ) , .A1( us23_n759 ) );
  NAND3_X1 us23_U439 (.ZN( sa21_sr_4 ) , .A3( us23_n737 ) , .A2( us23_n738 ) , .A1( us23_n739 ) );
  NOR2_X1 us23_U44 (.ZN( us23_n706 ) , .A2( us23_n775 ) , .A1( us23_n799 ) );
  NAND3_X1 us23_U440 (.A3( us23_n674 ) , .A2( us23_n675 ) , .A1( us23_n676 ) , .ZN( us23_n806 ) );
  NAND3_X1 us23_U441 (.ZN( us23_n637 ) , .A3( us23_n707 ) , .A2( us23_n723 ) , .A1( us23_n791 ) );
  NAND3_X1 us23_U442 (.A3( us23_n617 ) , .A2( us23_n618 ) , .A1( us23_n619 ) , .ZN( us23_n724 ) );
  NAND3_X1 us23_U443 (.A3( us23_n584 ) , .A2( us23_n585 ) , .A1( us23_n586 ) , .ZN( us23_n620 ) );
  NAND3_X1 us23_U444 (.ZN( us23_n564 ) , .A3( us23_n679 ) , .A2( us23_n749 ) , .A1( us23_n784 ) );
  NAND3_X1 us23_U445 (.A3( us23_n522 ) , .A2( us23_n523 ) , .A1( us23_n524 ) , .ZN( us23_n741 ) );
  NAND3_X1 us23_U446 (.A3( us23_n511 ) , .A1( us23_n512 ) , .ZN( us23_n607 ) , .A2( us23_n870 ) );
  NAND3_X1 us23_U447 (.A3( us23_n466 ) , .A2( us23_n467 ) , .A1( us23_n468 ) , .ZN( us23_n776 ) );
  NAND4_X1 us23_U448 (.A4( us23_n632 ) , .A3( us23_n633 ) , .A2( us23_n634 ) , .A1( us23_n635 ) , .ZN( us23_n742 ) );
  NOR2_X1 us23_U45 (.ZN( us23_n803 ) , .A1( us23_n853 ) , .A2( us23_n860 ) );
  NAND4_X1 us23_U46 (.ZN( sa21_sr_7 ) , .A4( us23_n821 ) , .A3( us23_n822 ) , .A2( us23_n823 ) , .A1( us23_n824 ) );
  AOI222_X1 us23_U47 (.C2( us23_n808 ) , .B2( us23_n809 ) , .A2( us23_n810 ) , .ZN( us23_n822 ) , .C1( us23_n831 ) , .A1( us23_n838 ) , .B1( us23_n852 ) );
  NOR4_X1 us23_U48 (.A4( us23_n817 ) , .A3( us23_n818 ) , .A2( us23_n819 ) , .A1( us23_n820 ) , .ZN( us23_n821 ) );
  AOI211_X1 us23_U49 (.B( us23_n806 ) , .A( us23_n807 ) , .ZN( us23_n823 ) , .C1( us23_n841 ) , .C2( us23_n849 ) );
  NOR3_X1 us23_U5 (.ZN( us23_n503 ) , .A2( us23_n678 ) , .A3( us23_n776 ) , .A1( us23_n875 ) );
  NAND4_X1 us23_U50 (.ZN( sa21_sr_0 ) , .A4( us23_n500 ) , .A3( us23_n501 ) , .A2( us23_n502 ) , .A1( us23_n503 ) );
  NOR4_X1 us23_U51 (.A4( us23_n497 ) , .A3( us23_n498 ) , .A2( us23_n499 ) , .ZN( us23_n500 ) , .A1( us23_n526 ) );
  AOI221_X1 us23_U52 (.A( us23_n496 ) , .ZN( us23_n501 ) , .B2( us23_n842 ) , .C1( us23_n845 ) , .C2( us23_n859 ) , .B1( us23_n861 ) );
  AOI211_X1 us23_U53 (.A( us23_n495 ) , .ZN( us23_n502 ) , .B( us23_n801 ) , .C2( us23_n838 ) , .C1( us23_n850 ) );
  AND3_X1 us23_U54 (.ZN( us23_n438 ) , .A2( us23_n642 ) , .A3( us23_n643 ) , .A1( us23_n645 ) );
  NAND4_X1 us23_U55 (.ZN( sa21_sr_1 ) , .A4( us23_n594 ) , .A3( us23_n595 ) , .A2( us23_n596 ) , .A1( us23_n597 ) );
  NOR4_X1 us23_U56 (.A4( us23_n590 ) , .A3( us23_n591 ) , .A2( us23_n592 ) , .A1( us23_n593 ) , .ZN( us23_n594 ) );
  AOI211_X1 us23_U57 (.B( us23_n588 ) , .A( us23_n589 ) , .ZN( us23_n595 ) , .C2( us23_n810 ) , .C1( us23_n832 ) );
  AOI211_X1 us23_U58 (.A( us23_n587 ) , .ZN( us23_n596 ) , .B( us23_n620 ) , .C1( us23_n844 ) , .C2( us23_n854 ) );
  NOR2_X1 us23_U59 (.ZN( us23_n624 ) , .A2( us23_n835 ) , .A1( us23_n838 ) );
  INV_X1 us23_U6 (.A( us23_n705 ) , .ZN( us23_n875 ) );
  NOR4_X1 us23_U60 (.A4( us23_n628 ) , .A3( us23_n629 ) , .A2( us23_n630 ) , .A1( us23_n631 ) , .ZN( us23_n632 ) );
  AOI211_X1 us23_U61 (.B( us23_n622 ) , .A( us23_n623 ) , .ZN( us23_n634 ) , .C2( us23_n835 ) , .C1( us23_n862 ) );
  NOR4_X1 us23_U62 (.A4( us23_n625 ) , .A3( us23_n626 ) , .A2( us23_n627 ) , .ZN( us23_n633 ) , .A1( us23_n663 ) );
  NAND4_X1 us23_U63 (.A4( us23_n656 ) , .A3( us23_n657 ) , .A2( us23_n658 ) , .A1( us23_n659 ) , .ZN( us23_n799 ) );
  NOR3_X1 us23_U64 (.A3( us23_n650 ) , .A2( us23_n651 ) , .A1( us23_n652 ) , .ZN( us23_n657 ) );
  NOR3_X1 us23_U65 (.A3( us23_n647 ) , .A2( us23_n648 ) , .A1( us23_n649 ) , .ZN( us23_n658 ) );
  NOR3_X1 us23_U66 (.A3( us23_n653 ) , .A2( us23_n654 ) , .A1( us23_n655 ) , .ZN( us23_n656 ) );
  NAND4_X1 us23_U67 (.A4( us23_n771 ) , .A3( us23_n772 ) , .A2( us23_n773 ) , .A1( us23_n774 ) , .ZN( us23_n800 ) );
  NOR3_X1 us23_U68 (.A3( us23_n764 ) , .A2( us23_n765 ) , .A1( us23_n766 ) , .ZN( us23_n772 ) );
  NOR4_X1 us23_U69 (.A4( us23_n767 ) , .A3( us23_n768 ) , .A2( us23_n769 ) , .A1( us23_n770 ) , .ZN( us23_n771 ) );
  NOR3_X1 us23_U7 (.A3( us23_n620 ) , .A2( us23_n621 ) , .ZN( us23_n635 ) , .A1( us23_n724 ) );
  AOI222_X1 us23_U70 (.ZN( us23_n774 ) , .A1( us23_n829 ) , .C1( us23_n833 ) , .B2( us23_n840 ) , .A2( us23_n849 ) , .B1( us23_n860 ) , .C2( us23_n872 ) );
  NOR4_X1 us23_U71 (.A4( us23_n576 ) , .A3( us23_n577 ) , .A2( us23_n578 ) , .ZN( us23_n585 ) , .A1( us23_n682 ) );
  NOR4_X1 us23_U72 (.A1( us23_n583 ) , .ZN( us23_n584 ) , .A3( us23_n651 ) , .A2( us23_n661 ) , .A4( us23_n766 ) );
  AOI221_X1 us23_U73 (.A( us23_n575 ) , .ZN( us23_n586 ) , .B2( us23_n830 ) , .C2( us23_n842 ) , .B1( us23_n853 ) , .C1( us23_n860 ) );
  NOR2_X1 us23_U74 (.ZN( us23_n760 ) , .A1( us23_n832 ) , .A2( us23_n833 ) );
  NAND4_X1 us23_U75 (.A4( us23_n455 ) , .A3( us23_n456 ) , .A2( us23_n457 ) , .A1( us23_n458 ) , .ZN( us23_n678 ) );
  NOR3_X1 us23_U76 (.ZN( us23_n456 ) , .A3( us23_n529 ) , .A1( us23_n554 ) , .A2( us23_n569 ) );
  NOR4_X1 us23_U77 (.ZN( us23_n457 ) , .A2( us23_n508 ) , .A1( us23_n598 ) , .A4( us23_n627 ) , .A3( us23_n710 ) );
  NOR4_X1 us23_U78 (.ZN( us23_n455 ) , .A2( us23_n516 ) , .A1( us23_n542 ) , .A3( us23_n578 ) , .A4( us23_n614 ) );
  NAND4_X1 us23_U79 (.A4( us23_n602 ) , .A3( us23_n603 ) , .A2( us23_n604 ) , .A1( us23_n605 ) , .ZN( us23_n721 ) );
  NOR2_X1 us23_U8 (.ZN( us23_n574 ) , .A1( us23_n621 ) , .A2( us23_n744 ) );
  NOR3_X1 us23_U80 (.A1( us23_n598 ) , .ZN( us23_n603 ) , .A3( us23_n662 ) , .A2( us23_n769 ) );
  NOR4_X1 us23_U81 (.A3( us23_n599 ) , .A2( us23_n600 ) , .A1( us23_n601 ) , .ZN( us23_n602 ) , .A4( us23_n654 ) );
  AOI222_X1 us23_U82 (.ZN( us23_n605 ) , .A1( us23_n829 ) , .C2( us23_n836 ) , .B1( us23_n841 ) , .A2( us23_n855 ) , .B2( us23_n860 ) , .C1( us23_n867 ) );
  NAND4_X1 us23_U83 (.A4( us23_n534 ) , .A3( us23_n535 ) , .A2( us23_n536 ) , .A1( us23_n537 ) , .ZN( us23_n621 ) );
  NOR4_X1 us23_U84 (.A4( us23_n525 ) , .A2( us23_n526 ) , .A1( us23_n527 ) , .ZN( us23_n537 ) , .A3( us23_n700 ) );
  NOR4_X1 us23_U85 (.A1( us23_n530 ) , .ZN( us23_n535 ) , .A2( us23_n653 ) , .A4( us23_n667 ) , .A3( us23_n764 ) );
  NOR4_X1 us23_U86 (.A4( us23_n528 ) , .A3( us23_n529 ) , .ZN( us23_n536 ) , .A2( us23_n683 ) , .A1( us23_n793 ) );
  NOR2_X1 us23_U87 (.ZN( us23_n685 ) , .A1( us23_n830 ) , .A2( us23_n831 ) );
  NAND4_X1 us23_U88 (.A4( us23_n547 ) , .A3( us23_n548 ) , .A2( us23_n549 ) , .A1( us23_n550 ) , .ZN( us23_n744 ) );
  NOR3_X1 us23_U89 (.ZN( us23_n548 ) , .A2( us23_n650 ) , .A1( us23_n666 ) , .A3( us23_n770 ) );
  NOR2_X1 us23_U9 (.A1( us23_n677 ) , .ZN( us23_n692 ) , .A2( us23_n806 ) );
  AOI211_X1 us23_U90 (.B( us23_n538 ) , .A( us23_n539 ) , .ZN( us23_n550 ) , .C2( us23_n838 ) , .C1( us23_n850 ) );
  NOR4_X1 us23_U91 (.A4( us23_n543 ) , .A3( us23_n544 ) , .A2( us23_n545 ) , .A1( us23_n546 ) , .ZN( us23_n547 ) );
  NAND4_X1 us23_U92 (.A4( us23_n478 ) , .A3( us23_n479 ) , .A2( us23_n480 ) , .A1( us23_n481 ) , .ZN( us23_n693 ) );
  NOR3_X1 us23_U93 (.ZN( us23_n479 ) , .A2( us23_n507 ) , .A3( us23_n600 ) , .A1( us23_n609 ) );
  AOI211_X1 us23_U94 (.B( us23_n476 ) , .A( us23_n477 ) , .ZN( us23_n481 ) , .C2( us23_n832 ) , .C1( us23_n860 ) );
  NOR4_X1 us23_U95 (.ZN( us23_n480 ) , .A3( us23_n531 ) , .A4( us23_n544 ) , .A2( us23_n566 ) , .A1( us23_n716 ) );
  NOR4_X1 us23_U96 (.ZN( us23_n619 ) , .A1( us23_n655 ) , .A3( us23_n665 ) , .A4( us23_n681 ) , .A2( us23_n765 ) );
  NOR4_X1 us23_U97 (.A4( us23_n608 ) , .A3( us23_n609 ) , .A2( us23_n610 ) , .A1( us23_n611 ) , .ZN( us23_n618 ) );
  NOR4_X1 us23_U98 (.A4( us23_n613 ) , .A3( us23_n614 ) , .A2( us23_n615 ) , .A1( us23_n616 ) , .ZN( us23_n617 ) );
  NAND4_X1 us23_U99 (.A4( us23_n484 ) , .A3( us23_n485 ) , .A2( us23_n486 ) , .A1( us23_n487 ) , .ZN( us23_n777 ) );
  NOR2_X1 us30_U10 (.ZN( us30_n575 ) , .A1( us30_n622 ) , .A2( us30_n745 ) );
  NOR2_X1 us30_U100 (.ZN( us30_n647 ) , .A1( us30_n854 ) , .A2( us30_n868 ) );
  NAND4_X1 us30_U101 (.A4( us30_n479 ) , .A3( us30_n480 ) , .A2( us30_n481 ) , .A1( us30_n482 ) , .ZN( us30_n694 ) );
  NOR3_X1 us30_U102 (.ZN( us30_n480 ) , .A2( us30_n508 ) , .A3( us30_n601 ) , .A1( us30_n610 ) );
  AOI211_X1 us30_U103 (.B( us30_n477 ) , .A( us30_n478 ) , .ZN( us30_n482 ) , .C2( us30_n833 ) , .C1( us30_n861 ) );
  NOR4_X1 us30_U104 (.ZN( us30_n481 ) , .A3( us30_n532 ) , .A4( us30_n545 ) , .A2( us30_n567 ) , .A1( us30_n717 ) );
  NAND4_X1 us30_U105 (.A4( us30_n548 ) , .A3( us30_n549 ) , .A2( us30_n550 ) , .A1( us30_n551 ) , .ZN( us30_n745 ) );
  NOR3_X1 us30_U106 (.ZN( us30_n549 ) , .A2( us30_n651 ) , .A1( us30_n667 ) , .A3( us30_n771 ) );
  AOI211_X1 us30_U107 (.B( us30_n539 ) , .A( us30_n540 ) , .ZN( us30_n551 ) , .C2( us30_n839 ) , .C1( us30_n851 ) );
  NOR4_X1 us30_U108 (.A4( us30_n544 ) , .A3( us30_n545 ) , .A2( us30_n546 ) , .A1( us30_n547 ) , .ZN( us30_n548 ) );
  NOR4_X1 us30_U109 (.ZN( us30_n620 ) , .A1( us30_n656 ) , .A3( us30_n666 ) , .A4( us30_n682 ) , .A2( us30_n766 ) );
  NOR2_X1 us30_U11 (.ZN( us30_n495 ) , .A1( us30_n678 ) , .A2( us30_n694 ) );
  NOR4_X1 us30_U110 (.A4( us30_n609 ) , .A3( us30_n610 ) , .A2( us30_n611 ) , .A1( us30_n612 ) , .ZN( us30_n619 ) );
  NOR4_X1 us30_U111 (.A4( us30_n614 ) , .A3( us30_n615 ) , .A2( us30_n616 ) , .A1( us30_n617 ) , .ZN( us30_n618 ) );
  NOR2_X1 us30_U112 (.ZN( us30_n686 ) , .A1( us30_n831 ) , .A2( us30_n832 ) );
  NAND4_X1 us30_U113 (.A4( us30_n485 ) , .A3( us30_n486 ) , .A2( us30_n487 ) , .A1( us30_n488 ) , .ZN( us30_n778 ) );
  NOR4_X1 us30_U114 (.A4( us30_n484 ) , .ZN( us30_n487 ) , .A1( us30_n566 ) , .A2( us30_n581 ) , .A3( us30_n602 ) );
  NOR4_X1 us30_U115 (.ZN( us30_n486 ) , .A1( us30_n507 ) , .A2( us30_n519 ) , .A4( us30_n546 ) , .A3( us30_n611 ) );
  NOR4_X1 us30_U116 (.ZN( us30_n485 ) , .A2( us30_n533 ) , .A1( us30_n558 ) , .A3( us30_n631 ) , .A4( us30_n718 ) );
  NAND4_X1 us30_U117 (.A4( us30_n691 ) , .A3( us30_n692 ) , .A1( us30_n693 ) , .ZN( us30_n776 ) , .A2( us30_n872 ) );
  AOI221_X1 us30_U118 (.A( us30_n681 ) , .ZN( us30_n692 ) , .B2( us30_n840 ) , .C1( us30_n842 ) , .C2( us30_n862 ) , .B1( us30_n865 ) );
  INV_X1 us30_U119 (.A( us30_n679 ) , .ZN( us30_n872 ) );
  NOR2_X1 us30_U12 (.A1( us30_n678 ) , .ZN( us30_n693 ) , .A2( us30_n807 ) );
  NOR4_X1 us30_U120 (.A4( us30_n687 ) , .A3( us30_n688 ) , .A2( us30_n689 ) , .A1( us30_n690 ) , .ZN( us30_n691 ) );
  NAND4_X1 us30_U121 (.A4( us30_n719 ) , .A3( us30_n720 ) , .A2( us30_n721 ) , .ZN( us30_n741 ) , .A1( us30_n857 ) );
  INV_X1 us30_U122 (.A( us30_n709 ) , .ZN( us30_n857 ) );
  AOI221_X1 us30_U123 (.A( us30_n710 ) , .ZN( us30_n721 ) , .C2( us30_n844 ) , .B2( us30_n845 ) , .C1( us30_n861 ) , .B1( us30_n862 ) );
  NOR4_X1 us30_U124 (.A4( us30_n715 ) , .A3( us30_n716 ) , .A2( us30_n717 ) , .A1( us30_n718 ) , .ZN( us30_n719 ) );
  NAND4_X1 us30_U125 (.A4( us30_n473 ) , .A3( us30_n474 ) , .A2( us30_n475 ) , .A1( us30_n476 ) , .ZN( us30_n678 ) );
  NOR4_X1 us30_U126 (.ZN( us30_n475 ) , .A1( us30_n531 ) , .A3( us30_n568 ) , .A4( us30_n600 ) , .A2( us30_n642 ) );
  NOR4_X1 us30_U127 (.A4( us30_n470 ) , .ZN( us30_n476 ) , .A3( us30_n556 ) , .A1( us30_n735 ) , .A2( us30_n755 ) );
  NOR4_X1 us30_U128 (.ZN( us30_n474 ) , .A1( us30_n506 ) , .A3( us30_n544 ) , .A2( us30_n583 ) , .A4( us30_n716 ) );
  NOR2_X1 us30_U129 (.ZN( us30_n733 ) , .A2( us30_n832 ) , .A1( us30_n845 ) );
  NOR3_X1 us30_U13 (.ZN( us30_n504 ) , .A2( us30_n679 ) , .A3( us30_n777 ) , .A1( us30_n876 ) );
  NOR2_X1 us30_U130 (.ZN( us30_n789 ) , .A2( us30_n862 ) , .A1( us30_n868 ) );
  NAND4_X1 us30_U131 (.A4( us30_n573 ) , .A3( us30_n574 ) , .A1( us30_n575 ) , .ZN( us30_n723 ) , .A2( us30_n874 ) );
  AOI221_X1 us30_U132 (.A( us30_n564 ) , .C2( us30_n565 ) , .ZN( us30_n574 ) , .B2( us30_n845 ) , .B1( us30_n852 ) , .C1( us30_n853 ) );
  NOR4_X1 us30_U133 (.A4( us30_n569 ) , .A3( us30_n570 ) , .A2( us30_n571 ) , .A1( us30_n572 ) , .ZN( us30_n573 ) );
  INV_X1 us30_U134 (.A( us30_n607 ) , .ZN( us30_n874 ) );
  NAND4_X1 us30_U135 (.A4( us30_n633 ) , .A3( us30_n634 ) , .A2( us30_n635 ) , .A1( us30_n636 ) , .ZN( us30_n743 ) );
  AOI211_X1 us30_U136 (.B( us30_n623 ) , .A( us30_n624 ) , .ZN( us30_n635 ) , .C2( us30_n836 ) , .C1( us30_n863 ) );
  NOR4_X1 us30_U137 (.A4( us30_n629 ) , .A3( us30_n630 ) , .A2( us30_n631 ) , .A1( us30_n632 ) , .ZN( us30_n633 ) );
  NOR4_X1 us30_U138 (.A4( us30_n626 ) , .A3( us30_n627 ) , .A2( us30_n628 ) , .ZN( us30_n634 ) , .A1( us30_n664 ) );
  NAND4_X1 us30_U139 (.A4( us30_n493 ) , .A3( us30_n494 ) , .A1( us30_n495 ) , .ZN( us30_n802 ) , .A2( us30_n867 ) );
  INV_X1 us30_U14 (.A( us30_n706 ) , .ZN( us30_n876 ) );
  AOI221_X1 us30_U140 (.A( us30_n489 ) , .ZN( us30_n494 ) , .B2( us30_n836 ) , .C2( us30_n841 ) , .C1( us30_n851 ) , .B1( us30_n860 ) );
  INV_X1 us30_U141 (.A( us30_n778 ) , .ZN( us30_n867 ) );
  NOR4_X1 us30_U142 (.A2( us30_n491 ) , .A1( us30_n492 ) , .ZN( us30_n493 ) , .A3( us30_n580 ) , .A4( us30_n612 ) );
  NOR4_X1 us30_U143 (.A4( us30_n734 ) , .A3( us30_n735 ) , .A2( us30_n736 ) , .A1( us30_n737 ) , .ZN( us30_n738 ) );
  AOI211_X1 us30_U144 (.B( us30_n725 ) , .A( us30_n726 ) , .ZN( us30_n739 ) , .C1( us30_n843 ) , .C2( us30_n855 ) );
  NOR3_X1 us30_U145 (.A3( us30_n722 ) , .A1( us30_n723 ) , .ZN( us30_n740 ) , .A2( us30_n741 ) );
  INV_X1 us30_U146 (.A( us30_n762 ) , .ZN( us30_n830 ) );
  OR4_X1 us30_U147 (.A4( us30_n566 ) , .A3( us30_n567 ) , .A2( us30_n568 ) , .ZN( us30_n572 ) , .A1( us30_n665 ) );
  OR4_X1 us30_U148 (.A4( us30_n682 ) , .A3( us30_n683 ) , .A2( us30_n684 ) , .A1( us30_n685 ) , .ZN( us30_n690 ) );
  OR4_X1 us30_U149 (.ZN( us30_n466 ) , .A4( us30_n518 ) , .A3( us30_n529 ) , .A2( us30_n578 ) , .A1( us30_n712 ) );
  INV_X1 us30_U15 (.A( us30_n680 ) , .ZN( us30_n840 ) );
  OR4_X1 us30_U150 (.A4( us30_n518 ) , .A2( us30_n519 ) , .A1( us30_n520 ) , .ZN( us30_n522 ) , .A3( us30_n821 ) );
  OR4_X1 us30_U151 (.ZN( us30_n492 ) , .A4( us30_n534 ) , .A2( us30_n547 ) , .A1( us30_n559 ) , .A3( us30_n632 ) );
  OR4_X1 us30_U152 (.A4( us30_n580 ) , .A3( us30_n581 ) , .A2( us30_n582 ) , .A1( us30_n583 ) , .ZN( us30_n584 ) );
  INV_X1 us30_U153 (.A( us30_n697 ) , .ZN( us30_n838 ) );
  NAND2_X1 us30_U154 (.ZN( us30_n613 ) , .A2( us30_n837 ) , .A1( us30_n873 ) );
  OR3_X1 us30_U155 (.A3( us30_n506 ) , .A2( us30_n507 ) , .A1( us30_n508 ) , .ZN( us30_n511 ) );
  INV_X1 us30_U156 (.A( us30_n754 ) , .ZN( us30_n869 ) );
  OAI21_X1 us30_U157 (.B1( us30_n753 ) , .ZN( us30_n754 ) , .A( us30_n845 ) , .B2( us30_n868 ) );
  INV_X1 us30_U158 (.A( us30_n463 ) , .ZN( us30_n864 ) );
  OAI21_X1 us30_U159 (.ZN( us30_n463 ) , .B1( us30_n809 ) , .A( us30_n834 ) , .B2( us30_n851 ) );
  NOR4_X1 us30_U16 (.A4( us30_n445 ) , .A3( us30_n446 ) , .A2( us30_n516 ) , .A1( us30_n541 ) , .ZN( us30_n706 ) );
  INV_X1 us30_U160 (.A( us30_n672 ) , .ZN( us30_n859 ) );
  AOI21_X1 us30_U161 (.A( us30_n670 ) , .B1( us30_n671 ) , .ZN( us30_n672 ) , .B2( us30_n856 ) );
  OAI222_X1 us30_U162 (.B2( us30_n747 ) , .B1( us30_n748 ) , .A2( us30_n749 ) , .ZN( us30_n757 ) , .C2( us30_n805 ) , .C1( us30_n814 ) , .A1( us30_n817 ) );
  OAI222_X1 us30_U163 (.ZN( us30_n505 ) , .C2( us30_n625 ) , .B2( us30_n647 ) , .B1( us30_n747 ) , .A2( us30_n748 ) , .C1( us30_n805 ) , .A1( us30_n806 ) );
  OAI222_X1 us30_U164 (.B2( us30_n708 ) , .ZN( us30_n709 ) , .C2( us30_n724 ) , .B1( us30_n747 ) , .A1( us30_n806 ) , .C1( us30_n814 ) , .A2( us30_n815 ) );
  NAND2_X1 us30_U165 (.A1( us30_n447 ) , .A2( us30_n465 ) , .ZN( us30_n749 ) );
  AOI22_X1 us30_U166 (.ZN( us30_n696 ) , .A1( us30_n830 ) , .B2( us30_n843 ) , .A2( us30_n865 ) , .B1( us30_n868 ) );
  AOI22_X1 us30_U167 (.A2( us30_n782 ) , .ZN( us30_n783 ) , .B2( us30_n831 ) , .A1( us30_n834 ) , .B1( us30_n863 ) );
  INV_X1 us30_U168 (.A( us30_n730 ) , .ZN( us30_n839 ) );
  AOI221_X1 us30_U169 (.A( us30_n764 ) , .ZN( us30_n774 ) , .C2( us30_n810 ) , .B2( us30_n835 ) , .C1( us30_n855 ) , .B1( us30_n866 ) );
  OR3_X1 us30_U17 (.ZN( us30_n446 ) , .A1( us30_n528 ) , .A3( us30_n577 ) , .A2( us30_n875 ) );
  AOI21_X1 us30_U170 (.B2( us30_n763 ) , .ZN( us30_n764 ) , .A( us30_n788 ) , .B1( us30_n792 ) );
  INV_X1 us30_U171 (.A( us30_n761 ) , .ZN( us30_n835 ) );
  AOI221_X1 us30_U172 (.A( us30_n483 ) , .ZN( us30_n488 ) , .B1( us30_n831 ) , .C2( us30_n844 ) , .C1( us30_n852 ) , .B2( us30_n862 ) );
  OAI22_X1 us30_U173 (.ZN( us30_n483 ) , .A1( us30_n708 ) , .B2( us30_n785 ) , .A2( us30_n806 ) , .B1( us30_n812 ) );
  INV_X1 us30_U174 (.A( us30_n790 ) , .ZN( us30_n832 ) );
  NAND2_X1 us30_U175 (.A1( us30_n451 ) , .A2( us30_n453 ) , .ZN( us30_n762 ) );
  OAI221_X1 us30_U176 (.A( us30_n727 ) , .C2( us30_n728 ) , .B2( us30_n729 ) , .B1( us30_n730 ) , .ZN( us30_n737 ) , .C1( us30_n817 ) );
  AOI22_X1 us30_U177 (.ZN( us30_n727 ) , .B1( us30_n832 ) , .A2( us30_n838 ) , .A1( us30_n863 ) , .B2( us30_n866 ) );
  INV_X1 us30_U178 (.A( us30_n786 ) , .ZN( us30_n862 ) );
  OAI22_X1 us30_U179 (.ZN( us30_n710 ) , .A2( us30_n728 ) , .B2( us30_n729 ) , .A1( us30_n744 ) , .B1( us30_n813 ) );
  OR4_X1 us30_U18 (.A4( us30_n442 ) , .A2( us30_n443 ) , .A1( us30_n444 ) , .ZN( us30_n445 ) , .A3( us30_n553 ) );
  INV_X1 us30_U180 (.A( us30_n816 ) , .ZN( us30_n831 ) );
  OAI22_X1 us30_U181 (.ZN( us30_n489 ) , .A1( us30_n724 ) , .B2( us30_n728 ) , .B1( us30_n730 ) , .A2( us30_n779 ) );
  OAI22_X1 us30_U182 (.ZN( us30_n624 ) , .B1( us30_n669 ) , .B2( us30_n747 ) , .A1( us30_n815 ) , .A2( us30_n816 ) );
  INV_X1 us30_U183 (.A( us30_n744 ) , .ZN( us30_n837 ) );
  INV_X1 us30_U184 (.A( us30_n788 ) , .ZN( us30_n845 ) );
  OAI22_X1 us30_U185 (.B2( us30_n779 ) , .B1( us30_n780 ) , .ZN( us30_n781 ) , .A2( us30_n814 ) , .A1( us30_n815 ) );
  OAI22_X1 us30_U186 (.A1( us30_n724 ) , .ZN( us30_n726 ) , .B2( us30_n750 ) , .B1( us30_n812 ) , .A2( us30_n816 ) );
  INV_X1 us30_U187 (.A( us30_n805 ) , .ZN( us30_n860 ) );
  INV_X1 us30_U188 (.A( us30_n814 ) , .ZN( us30_n833 ) );
  INV_X1 us30_U189 (.A( us30_n669 ) , .ZN( us30_n865 ) );
  INV_X1 us30_U19 (.A( us30_n613 ) , .ZN( us30_n875 ) );
  OAI22_X1 us30_U190 (.B2( us30_n744 ) , .ZN( us30_n746 ) , .A2( us30_n762 ) , .B1( us30_n780 ) , .A1( us30_n792 ) );
  OAI22_X1 us30_U191 (.ZN( us30_n496 ) , .A2( us30_n744 ) , .A1( us30_n780 ) , .B1( us30_n791 ) , .B2( us30_n806 ) );
  OAI22_X1 us30_U192 (.B2( us30_n803 ) , .B1( us30_n804 ) , .A2( us30_n805 ) , .A1( us30_n806 ) , .ZN( us30_n808 ) );
  AOI211_X1 us30_U193 (.A( us30_n637 ) , .ZN( us30_n645 ) , .B( us30_n743 ) , .C2( us30_n839 ) , .C1( us30_n854 ) );
  OAI22_X1 us30_U194 (.ZN( us30_n637 ) , .A1( us30_n699 ) , .B2( us30_n728 ) , .A2( us30_n762 ) , .B1( us30_n816 ) );
  OAI22_X1 us30_U195 (.B1( us30_n490 ) , .ZN( us30_n491 ) , .A1( us30_n686 ) , .A2( us30_n763 ) , .B2( us30_n817 ) );
  NOR3_X1 us30_U196 (.ZN( us30_n490 ) , .A1( us30_n782 ) , .A2( us30_n850 ) , .A3( us30_n863 ) );
  INV_X1 us30_U197 (.A( us30_n750 ) , .ZN( us30_n842 ) );
  OAI22_X1 us30_U198 (.ZN( us30_n695 ) , .A2( us30_n730 ) , .A1( us30_n780 ) , .B1( us30_n791 ) , .B2( us30_n817 ) );
  NOR2_X1 us30_U199 (.ZN( us30_n715 ) , .A1( us30_n805 ) , .A2( us30_n817 ) );
  INV_X1 us30_U20 (.A( us30_n749 ) , .ZN( us30_n863 ) );
  NOR2_X1 us30_U200 (.ZN( us30_n666 ) , .A1( us30_n728 ) , .A2( us30_n803 ) );
  NOR2_X1 us30_U201 (.ZN( us30_n594 ) , .A2( us30_n697 ) , .A1( us30_n728 ) );
  NOR2_X1 us30_U202 (.ZN( us30_n570 ) , .A1( us30_n728 ) , .A2( us30_n806 ) );
  NOR2_X1 us30_U203 (.A2( us30_n744 ) , .ZN( us30_n755 ) , .A1( us30_n805 ) );
  NOR2_X1 us30_U204 (.ZN( us30_n735 ) , .A2( us30_n803 ) , .A1( us30_n805 ) );
  NOR2_X1 us30_U205 (.ZN( us30_n546 ) , .A2( us30_n780 ) , .A1( us30_n814 ) );
  NOR2_X1 us30_U206 (.ZN( us30_n577 ) , .A2( us30_n699 ) , .A1( us30_n814 ) );
  NOR2_X1 us30_U207 (.ZN( us30_n654 ) , .A1( us30_n728 ) , .A2( us30_n813 ) );
  NOR2_X1 us30_U208 (.ZN( us30_n718 ) , .A2( us30_n724 ) , .A1( us30_n744 ) );
  NOR2_X1 us30_U209 (.ZN( us30_n532 ) , .A2( us30_n749 ) , .A1( us30_n750 ) );
  AOI222_X1 us30_U21 (.ZN( us30_n605 ) , .B2( us30_n671 ) , .B1( us30_n753 ) , .C2( us30_n831 ) , .A1( us30_n833 ) , .A2( us30_n862 ) , .C1( us30_n863 ) );
  NOR2_X1 us30_U210 (.ZN( us30_n615 ) , .A1( us30_n785 ) , .A2( us30_n815 ) );
  NOR2_X1 us30_U211 (.ZN( us30_n629 ) , .A2( us30_n728 ) , .A1( us30_n785 ) );
  NOR2_X1 us30_U212 (.ZN( us30_n611 ) , .A2( us30_n780 ) , .A1( us30_n806 ) );
  NOR2_X1 us30_U213 (.ZN( us30_n628 ) , .A2( us30_n669 ) , .A1( us30_n785 ) );
  INV_X1 us30_U214 (.A( us30_n747 ) , .ZN( us30_n834 ) );
  INV_X1 us30_U215 (.A( us30_n728 ) , .ZN( us30_n852 ) );
  NOR2_X1 us30_U216 (.ZN( us30_n652 ) , .A1( us30_n669 ) , .A2( us30_n814 ) );
  NOR2_X1 us30_U217 (.A1( us30_n669 ) , .ZN( us30_n673 ) , .A2( us30_n744 ) );
  NOR2_X1 us30_U218 (.ZN( us30_n602 ) , .A1( us30_n669 ) , .A2( us30_n803 ) );
  NOR2_X1 us30_U219 (.A1( us30_n669 ) , .ZN( us30_n688 ) , .A2( us30_n816 ) );
  AOI222_X1 us30_U22 (.ZN( us30_n563 ) , .B1( us30_n830 ) , .C1( us30_n841 ) , .A2( us30_n843 ) , .A1( us30_n854 ) , .B2( us30_n863 ) , .C2( us30_n873 ) );
  NOR2_X1 us30_U220 (.A2( us30_n744 ) , .ZN( us30_n769 ) , .A1( us30_n812 ) );
  NOR2_X1 us30_U221 (.ZN( us30_n531 ) , .A2( us30_n780 ) , .A1( us30_n816 ) );
  INV_X1 us30_U222 (.A( us30_n792 ) , .ZN( us30_n851 ) );
  NOR2_X1 us30_U223 (.A2( us30_n708 ) , .A1( us30_n750 ) , .ZN( us30_n771 ) );
  NOR2_X1 us30_U224 (.ZN( us30_n599 ) , .A2( us30_n791 ) , .A1( us30_n816 ) );
  NOR2_X1 us30_U225 (.A1( us30_n669 ) , .ZN( us30_n766 ) , .A2( us30_n813 ) );
  NOR2_X1 us30_U226 (.ZN( us30_n601 ) , .A2( us30_n780 ) , .A1( us30_n803 ) );
  NOR2_X1 us30_U227 (.A1( us30_n699 ) , .ZN( us30_n768 ) , .A2( us30_n813 ) );
  NOR2_X1 us30_U228 (.ZN( us30_n541 ) , .A2( us30_n697 ) , .A1( us30_n699 ) );
  NOR2_X1 us30_U229 (.ZN( us30_n527 ) , .A1( us30_n669 ) , .A2( us30_n779 ) );
  AOI222_X1 us30_U23 (.ZN( us30_n660 ) , .A2( us30_n839 ) , .B1( us30_n841 ) , .C2( us30_n845 ) , .A1( us30_n860 ) , .C1( us30_n863 ) , .B2( us30_n870 ) );
  NOR2_X1 us30_U230 (.ZN( us30_n667 ) , .A1( us30_n750 ) , .A2( us30_n815 ) );
  NOR2_X1 us30_U231 (.ZN( us30_n555 ) , .A1( us30_n750 ) , .A2( us30_n791 ) );
  NOR2_X1 us30_U232 (.ZN( us30_n508 ) , .A2( us30_n780 ) , .A1( us30_n785 ) );
  NOR2_X1 us30_U233 (.ZN( us30_n543 ) , .A2( us30_n708 ) , .A1( us30_n785 ) );
  NOR2_X1 us30_U234 (.ZN( us30_n528 ) , .A2( us30_n724 ) , .A1( us30_n803 ) );
  NOR2_X1 us30_U235 (.ZN( us30_n664 ) , .A1( us30_n785 ) , .A2( us30_n791 ) );
  NOR2_X1 us30_U236 (.ZN( us30_n556 ) , .A1( us30_n762 ) , .A2( us30_n805 ) );
  INV_X1 us30_U237 (.A( us30_n806 ) , .ZN( us30_n841 ) );
  NOR2_X1 us30_U238 (.ZN( us30_n661 ) , .A1( us30_n729 ) , .A2( us30_n790 ) );
  OAI22_X1 us30_U239 (.B1( us30_n440 ) , .ZN( us30_n444 ) , .A2( us30_n728 ) , .A1( us30_n744 ) , .B2( us30_n749 ) );
  INV_X1 us30_U24 (.A( us30_n647 ) , .ZN( us30_n870 ) );
  NOR3_X1 us30_U240 (.ZN( us30_n440 ) , .A2( us30_n836 ) , .A3( us30_n837 ) , .A1( us30_n846 ) );
  NOR2_X1 us30_U241 (.ZN( us30_n507 ) , .A1( us30_n812 ) , .A2( us30_n817 ) );
  NOR2_X1 us30_U242 (.ZN( us30_n557 ) , .A1( us30_n792 ) , .A2( us30_n814 ) );
  NOR2_X1 us30_U243 (.ZN( us30_n545 ) , .A1( us30_n749 ) , .A2( us30_n814 ) );
  NOR2_X1 us30_U244 (.ZN( us30_n509 ) , .A1( us30_n729 ) , .A2( us30_n779 ) );
  NOR2_X1 us30_U245 (.ZN( us30_n662 ) , .A2( us30_n697 ) , .A1( us30_n729 ) );
  OAI22_X1 us30_U246 (.B2( us30_n750 ) , .B1( us30_n751 ) , .A1( us30_n752 ) , .ZN( us30_n756 ) , .A2( us30_n806 ) );
  NOR2_X1 us30_U247 (.ZN( us30_n751 ) , .A2( us30_n852 ) , .A1( us30_n860 ) );
  NOR3_X1 us30_U248 (.ZN( us30_n752 ) , .A2( us30_n853 ) , .A1( us30_n863 ) , .A3( us30_n865 ) );
  NOR2_X1 us30_U249 (.ZN( us30_n544 ) , .A2( us30_n785 ) , .A1( us30_n792 ) );
  NOR4_X1 us30_U25 (.ZN( us30_n473 ) , .A2( us30_n521 ) , .A4( us30_n594 ) , .A1( us30_n609 ) , .A3( us30_n629 ) );
  NOR2_X1 us30_U250 (.ZN( us30_n663 ) , .A1( us30_n729 ) , .A2( us30_n785 ) );
  NOR2_X1 us30_U251 (.ZN( us30_n530 ) , .A2( us30_n744 ) , .A1( us30_n792 ) );
  NOR2_X1 us30_U252 (.ZN( us30_n506 ) , .A2( us30_n728 ) , .A1( us30_n762 ) );
  NOR2_X1 us30_U253 (.ZN( us30_n631 ) , .A1( us30_n724 ) , .A2( us30_n813 ) );
  NOR2_X1 us30_U254 (.ZN( us30_n614 ) , .A1( us30_n762 ) , .A2( us30_n812 ) );
  NOR2_X1 us30_U255 (.A1( us30_n749 ) , .ZN( us30_n767 ) , .A2( us30_n803 ) );
  NOR2_X1 us30_U256 (.ZN( us30_n516 ) , .A1( us30_n708 ) , .A2( us30_n744 ) );
  NOR2_X1 us30_U257 (.ZN( us30_n670 ) , .A1( us30_n790 ) , .A2( us30_n805 ) );
  NOR2_X1 us30_U258 (.ZN( us30_n558 ) , .A1( us30_n708 ) , .A2( us30_n816 ) );
  NOR2_X1 us30_U259 (.A2( us30_n697 ) , .ZN( us30_n716 ) , .A1( us30_n792 ) );
  NOR4_X1 us30_U26 (.ZN( us30_n479 ) , .A1( us30_n520 ) , .A4( us30_n557 ) , .A3( us30_n582 ) , .A2( us30_n630 ) );
  NOR2_X1 us30_U260 (.ZN( us30_n517 ) , .A1( us30_n708 ) , .A2( us30_n803 ) );
  NOR2_X1 us30_U261 (.ZN( us30_n521 ) , .A1( us30_n790 ) , .A2( us30_n812 ) );
  NOR2_X1 us30_U262 (.ZN( us30_n630 ) , .A1( us30_n747 ) , .A2( us30_n815 ) );
  NOR2_X1 us30_U263 (.ZN( us30_n655 ) , .A1( us30_n790 ) , .A2( us30_n815 ) );
  INV_X1 us30_U264 (.A( us30_n763 ) , .ZN( us30_n866 ) );
  AOI21_X1 us30_U265 (.ZN( us30_n552 ) , .B1( us30_n669 ) , .A( us30_n697 ) , .B2( us30_n805 ) );
  NOR2_X1 us30_U266 (.ZN( us30_n668 ) , .A2( us30_n708 ) , .A1( us30_n790 ) );
  NOR2_X1 us30_U267 (.ZN( us30_n542 ) , .A1( us30_n762 ) , .A2( us30_n791 ) );
  NOR2_X1 us30_U268 (.ZN( us30_n656 ) , .A1( us30_n747 ) , .A2( us30_n780 ) );
  NOR2_X1 us30_U269 (.ZN( us30_n609 ) , .A2( us30_n724 ) , .A1( us30_n817 ) );
  NOR4_X1 us30_U27 (.A4( us30_n532 ) , .A3( us30_n533 ) , .A2( us30_n534 ) , .ZN( us30_n535 ) , .A1( us30_n820 ) );
  INV_X1 us30_U270 (.A( us30_n729 ) , .ZN( us30_n868 ) );
  AOI21_X1 us30_U271 (.B1( us30_n625 ) , .ZN( us30_n627 ) , .A( us30_n763 ) , .B2( us30_n814 ) );
  AOI21_X1 us30_U272 (.ZN( us30_n650 ) , .A( us30_n779 ) , .B1( us30_n792 ) , .B2( us30_n805 ) );
  AOI21_X1 us30_U273 (.A( us30_n815 ) , .B2( us30_n816 ) , .B1( us30_n817 ) , .ZN( us30_n818 ) );
  NOR2_X1 us30_U274 (.ZN( us30_n579 ) , .A2( us30_n708 ) , .A1( us30_n730 ) );
  NOR2_X1 us30_U275 (.ZN( us30_n533 ) , .A2( us30_n724 ) , .A1( us30_n730 ) );
  NOR2_X1 us30_U276 (.ZN( us30_n642 ) , .A2( us30_n788 ) , .A1( us30_n791 ) );
  AOI21_X1 us30_U277 (.A( us30_n812 ) , .B2( us30_n813 ) , .B1( us30_n814 ) , .ZN( us30_n819 ) );
  NOR2_X1 us30_U278 (.A2( us30_n708 ) , .A1( us30_n762 ) , .ZN( us30_n794 ) );
  NOR2_X1 us30_U279 (.A2( us30_n697 ) , .A1( us30_n780 ) , .ZN( us30_n820 ) );
  NOR4_X1 us30_U28 (.ZN( us30_n456 ) , .A2( us30_n517 ) , .A1( us30_n543 ) , .A3( us30_n579 ) , .A4( us30_n615 ) );
  AOI21_X1 us30_U280 (.ZN( us30_n626 ) , .B2( us30_n669 ) , .A( us30_n790 ) , .B1( us30_n791 ) );
  AOI21_X1 us30_U281 (.ZN( us30_n499 ) , .B1( us30_n680 ) , .A( us30_n812 ) , .B2( us30_n816 ) );
  NOR2_X1 us30_U282 (.ZN( us30_n520 ) , .A2( us30_n708 ) , .A1( us30_n814 ) );
  AOI21_X1 us30_U283 (.ZN( us30_n477 ) , .A( us30_n669 ) , .B1( us30_n750 ) , .B2( us30_n806 ) );
  NOR2_X1 us30_U284 (.ZN( us30_n582 ) , .A1( us30_n744 ) , .A2( us30_n815 ) );
  AOI21_X1 us30_U285 (.ZN( us30_n593 ) , .B1( us30_n750 ) , .A( us30_n792 ) , .B2( us30_n813 ) );
  AOI21_X1 us30_U286 (.ZN( us30_n515 ) , .A( us30_n729 ) , .B1( us30_n750 ) , .B2( us30_n803 ) );
  NOR2_X1 us30_U287 (.A1( us30_n697 ) , .ZN( us30_n770 ) , .A2( us30_n815 ) );
  AOI21_X1 us30_U288 (.ZN( us30_n510 ) , .B2( us30_n669 ) , .A( us30_n730 ) , .B1( us30_n815 ) );
  NOR2_X1 us30_U289 (.ZN( us30_n519 ) , .A2( us30_n699 ) , .A1( us30_n816 ) );
  NOR4_X1 us30_U29 (.A4( us30_n541 ) , .A3( us30_n542 ) , .A2( us30_n543 ) , .ZN( us30_n550 ) , .A1( us30_n688 ) );
  NOR2_X1 us30_U290 (.ZN( us30_n559 ) , .A2( us30_n791 ) , .A1( us30_n803 ) );
  NOR2_X1 us30_U291 (.ZN( us30_n581 ) , .A1( us30_n669 ) , .A2( us30_n788 ) );
  INV_X1 us30_U292 (.A( us30_n813 ) , .ZN( us30_n836 ) );
  NOR2_X1 us30_U293 (.ZN( us30_n683 ) , .A2( us30_n699 ) , .A1( us30_n803 ) );
  AOI21_X1 us30_U294 (.ZN( us30_n589 ) , .B2( us30_n699 ) , .B1( us30_n815 ) , .A( us30_n817 ) );
  AOI21_X1 us30_U295 (.ZN( us30_n539 ) , .B2( us30_n812 ) , .A( us30_n814 ) , .B1( us30_n815 ) );
  AOI21_X1 us30_U296 (.ZN( us30_n540 ) , .A( us30_n763 ) , .B2( us30_n779 ) , .B1( us30_n817 ) );
  AOI21_X1 us30_U297 (.B1( us30_n699 ) , .ZN( us30_n700 ) , .A( us30_n732 ) , .B2( us30_n763 ) );
  AOI21_X1 us30_U298 (.ZN( us30_n591 ) , .B2( us30_n763 ) , .A( us30_n785 ) , .B1( us30_n812 ) );
  AOI21_X1 us30_U299 (.ZN( us30_n498 ) , .A( us30_n724 ) , .B2( us30_n762 ) , .B1( us30_n814 ) );
  NAND2_X1 us30_U3 (.A2( us30_n448 ) , .A1( us30_n464 ) , .ZN( us30_n815 ) );
  AOI221_X1 us30_U30 (.A( us30_n713 ) , .B2( us30_n714 ) , .ZN( us30_n720 ) , .C1( us30_n832 ) , .B1( us30_n839 ) , .C2( us30_n863 ) );
  NOR2_X1 us30_U300 (.ZN( us30_n547 ) , .A1( us30_n699 ) , .A2( us30_n744 ) );
  INV_X1 us30_U301 (.A( us30_n791 ) , .ZN( us30_n873 ) );
  AOI21_X1 us30_U302 (.ZN( us30_n649 ) , .B1( us30_n729 ) , .B2( us30_n763 ) , .A( us30_n813 ) );
  NOR2_X1 us30_U303 (.ZN( us30_n685 ) , .A1( us30_n729 ) , .A2( us30_n816 ) );
  AOI21_X1 us30_U304 (.B1( us30_n686 ) , .ZN( us30_n687 ) , .A( us30_n728 ) , .B2( us30_n761 ) );
  AOI21_X1 us30_U305 (.ZN( us30_n569 ) , .B1( us30_n750 ) , .B2( us30_n762 ) , .A( us30_n780 ) );
  AOI21_X1 us30_U306 (.ZN( us30_n571 ) , .B2( us30_n697 ) , .B1( us30_n806 ) , .A( us30_n812 ) );
  NOR2_X1 us30_U307 (.ZN( us30_n568 ) , .A1( us30_n729 ) , .A2( us30_n762 ) );
  NOR2_X1 us30_U308 (.ZN( us30_n566 ) , .A2( us30_n697 ) , .A1( us30_n763 ) );
  AOI21_X1 us30_U309 (.ZN( us30_n640 ) , .B2( us30_n747 ) , .A( us30_n792 ) , .B1( us30_n803 ) );
  OR2_X1 us30_U31 (.A2( us30_n711 ) , .A1( us30_n712 ) , .ZN( us30_n713 ) );
  INV_X1 us30_U310 (.A( us30_n699 ) , .ZN( us30_n853 ) );
  AOI21_X1 us30_U311 (.ZN( us30_n514 ) , .A( us30_n779 ) , .B2( us30_n792 ) , .B1( us30_n812 ) );
  AOI21_X1 us30_U312 (.ZN( us30_n639 ) , .B2( us30_n749 ) , .A( us30_n788 ) , .B1( us30_n812 ) );
  NAND2_X1 us30_U313 (.ZN( us30_n753 ) , .A1( us30_n763 ) , .A2( us30_n805 ) );
  NOR2_X1 us30_U314 (.ZN( us30_n665 ) , .A1( us30_n780 ) , .A2( us30_n813 ) );
  AOI21_X1 us30_U315 (.ZN( us30_n564 ) , .B1( us30_n724 ) , .A( us30_n779 ) , .B2( us30_n791 ) );
  AOI21_X1 us30_U316 (.ZN( us30_n497 ) , .A( us30_n779 ) , .B2( us30_n791 ) , .B1( us30_n804 ) );
  AOI21_X1 us30_U317 (.ZN( us30_n689 ) , .B2( us30_n749 ) , .B1( us30_n763 ) , .A( us30_n806 ) );
  AOI21_X1 us30_U318 (.ZN( us30_n450 ) , .B2( us30_n792 ) , .A( us30_n803 ) , .B1( us30_n815 ) );
  NOR2_X1 us30_U319 (.ZN( us30_n567 ) , .A1( us30_n747 ) , .A2( us30_n805 ) );
  NOR2_X1 us30_U32 (.ZN( us30_n680 ) , .A2( us30_n834 ) , .A1( us30_n839 ) );
  NOR2_X1 us30_U320 (.ZN( us30_n529 ) , .A1( us30_n708 ) , .A2( us30_n779 ) );
  NOR2_X1 us30_U321 (.ZN( us30_n578 ) , .A1( us30_n708 ) , .A2( us30_n813 ) );
  AOI21_X1 us30_U322 (.ZN( us30_n478 ) , .B2( us30_n697 ) , .A( us30_n749 ) , .B1( us30_n779 ) );
  AOI21_X1 us30_U323 (.A( us30_n790 ) , .B2( us30_n791 ) , .B1( us30_n792 ) , .ZN( us30_n793 ) );
  NOR2_X1 us30_U324 (.ZN( us30_n684 ) , .A1( us30_n791 ) , .A2( us30_n813 ) );
  AOI21_X1 us30_U325 (.A( us30_n733 ) , .ZN( us30_n734 ) , .B2( us30_n780 ) , .B1( us30_n792 ) );
  NOR2_X1 us30_U326 (.A2( us30_n813 ) , .A1( us30_n815 ) , .ZN( us30_n821 ) );
  AOI21_X1 us30_U327 (.ZN( us30_n641 ) , .B1( us30_n680 ) , .A( us30_n791 ) , .B2( us30_n817 ) );
  NOR2_X1 us30_U328 (.ZN( us30_n711 ) , .A1( us30_n762 ) , .A2( us30_n763 ) );
  NOR2_X1 us30_U329 (.ZN( us30_n583 ) , .A1( us30_n792 ) , .A2( us30_n817 ) );
  AOI222_X1 us30_U33 (.ZN( us30_n469 ) , .B1( us30_n832 ) , .A1( us30_n839 ) , .C1( us30_n842 ) , .C2( us30_n851 ) , .A2( us30_n855 ) , .B2( us30_n865 ) );
  NOR2_X1 us30_U330 (.ZN( us30_n534 ) , .A1( us30_n724 ) , .A2( us30_n788 ) );
  NOR2_X1 us30_U331 (.ZN( us30_n632 ) , .A2( us30_n697 ) , .A1( us30_n724 ) );
  NOR2_X1 us30_U332 (.ZN( us30_n682 ) , .A2( us30_n708 ) , .A1( us30_n817 ) );
  NOR2_X1 us30_U333 (.ZN( us30_n580 ) , .A2( us30_n697 ) , .A1( us30_n791 ) );
  INV_X1 us30_U334 (.A( us30_n815 ) , .ZN( us30_n855 ) );
  AOI21_X1 us30_U335 (.ZN( us30_n442 ) , .A( us30_n699 ) , .B1( us30_n733 ) , .B2( us30_n750 ) );
  INV_X1 us30_U336 (.A( us30_n780 ) , .ZN( us30_n850 ) );
  INV_X1 us30_U337 (.A( us30_n785 ) , .ZN( us30_n846 ) );
  NAND2_X1 us30_U338 (.ZN( us30_n714 ) , .A1( us30_n728 ) , .A2( us30_n780 ) );
  NAND2_X1 us30_U339 (.A2( us30_n762 ) , .A1( us30_n806 ) , .ZN( us30_n810 ) );
  NOR4_X1 us30_U34 (.A1( us30_n466 ) , .ZN( us30_n467 ) , .A4( us30_n542 ) , .A2( us30_n554 ) , .A3( us30_n614 ) );
  AOI21_X1 us30_U340 (.ZN( us30_n443 ) , .B1( us30_n789 ) , .B2( us30_n791 ) , .A( us30_n814 ) );
  NAND2_X1 us30_U341 (.ZN( us30_n671 ) , .A1( us30_n806 ) , .A2( us30_n816 ) );
  NOR2_X1 us30_U342 (.ZN( us30_n484 ) , .A1( us30_n788 ) , .A2( us30_n805 ) );
  NOR2_X1 us30_U343 (.ZN( us30_n470 ) , .A2( us30_n779 ) , .A1( us30_n815 ) );
  NOR2_X1 us30_U344 (.ZN( us30_n712 ) , .A2( us30_n724 ) , .A1( us30_n790 ) );
  OAI21_X1 us30_U345 (.A( us30_n787 ) , .B2( us30_n788 ) , .B1( us30_n789 ) , .ZN( us30_n795 ) );
  OAI21_X1 us30_U346 (.ZN( us30_n787 ) , .A( us30_n839 ) , .B1( us30_n863 ) , .B2( us30_n873 ) );
  NOR2_X1 us30_U347 (.ZN( us30_n526 ) , .A1( us30_n724 ) , .A2( us30_n750 ) );
  NAND2_X1 us30_U348 (.A1( us30_n699 ) , .A2( us30_n729 ) , .ZN( us30_n782 ) );
  NOR2_X1 us30_U349 (.ZN( us30_n518 ) , .A1( us30_n708 ) , .A2( us30_n788 ) );
  AOI221_X1 us30_U35 (.ZN( us30_n468 ) , .C2( us30_n714 ) , .B2( us30_n831 ) , .C1( us30_n845 ) , .B1( us30_n860 ) , .A( us30_n864 ) );
  OAI21_X1 us30_U350 (.A( us30_n698 ) , .ZN( us30_n702 ) , .B2( us30_n750 ) , .B1( us30_n804 ) );
  OAI21_X1 us30_U351 (.ZN( us30_n698 ) , .B2( us30_n833 ) , .B1( us30_n838 ) , .A( us30_n860 ) );
  OAI21_X1 us30_U352 (.A( us30_n731 ) , .B1( us30_n732 ) , .ZN( us30_n736 ) , .B2( us30_n805 ) );
  OAI21_X1 us30_U353 (.ZN( us30_n731 ) , .A( us30_n833 ) , .B2( us30_n852 ) , .B1( us30_n873 ) );
  INV_X1 us30_U354 (.A( us30_n817 ) , .ZN( us30_n844 ) );
  INV_X1 us30_U355 (.A( us30_n724 ) , .ZN( us30_n856 ) );
  AND2_X1 us30_U356 (.ZN( us30_n732 ) , .A1( us30_n779 ) , .A2( us30_n785 ) );
  NAND2_X1 us30_U357 (.A1( us30_n447 ) , .A2( us30_n449 ) , .ZN( us30_n805 ) );
  NAND2_X1 us30_U358 (.A1( us30_n451 ) , .A2( us30_n454 ) , .ZN( us30_n814 ) );
  NAND2_X1 us30_U359 (.A1( us30_n452 ) , .A2( us30_n465 ) , .ZN( us30_n669 ) );
  NOR4_X1 us30_U36 (.A4( us30_n514 ) , .A3( us30_n515 ) , .A2( us30_n516 ) , .A1( us30_n517 ) , .ZN( us30_n524 ) );
  NAND2_X1 us30_U360 (.A2( us30_n448 ) , .A1( us30_n460 ) , .ZN( us30_n728 ) );
  NAND2_X1 us30_U361 (.A1( us30_n455 ) , .A2( us30_n462 ) , .ZN( us30_n750 ) );
  NAND2_X1 us30_U362 (.A2( us30_n453 ) , .A1( us30_n455 ) , .ZN( us30_n806 ) );
  NAND2_X1 us30_U363 (.A1( us30_n451 ) , .A2( us30_n471 ) , .ZN( us30_n816 ) );
  NAND2_X1 us30_U364 (.A1( us30_n454 ) , .A2( us30_n461 ) , .ZN( us30_n813 ) );
  NAND2_X1 us30_U365 (.A1( us30_n455 ) , .A2( us30_n471 ) , .ZN( us30_n803 ) );
  NAND2_X1 us30_U366 (.A1( us30_n453 ) , .A2( us30_n461 ) , .ZN( us30_n744 ) );
  NAND2_X1 us30_U367 (.A1( us30_n453 ) , .A2( us30_n472 ) , .ZN( us30_n785 ) );
  NAND2_X1 us30_U368 (.A2( us30_n454 ) , .A1( us30_n472 ) , .ZN( us30_n779 ) );
  NAND2_X1 us30_U369 (.A2( us30_n464 ) , .A1( us30_n465 ) , .ZN( us30_n812 ) );
  AOI222_X1 us30_U37 (.ZN( us30_n525 ) , .A1( us30_n834 ) , .B2( us30_n837 ) , .C1( us30_n844 ) , .C2( us30_n850 ) , .A2( us30_n852 ) , .B1( us30_n866 ) );
  NAND2_X1 us30_U370 (.A1( us30_n441 ) , .A2( us30_n460 ) , .ZN( us30_n699 ) );
  NAND2_X1 us30_U371 (.A2( us30_n449 ) , .A1( us30_n452 ) , .ZN( us30_n763 ) );
  NAND2_X1 us30_U372 (.A2( us30_n448 ) , .A1( us30_n452 ) , .ZN( us30_n729 ) );
  NAND2_X1 us30_U373 (.A2( us30_n461 ) , .A1( us30_n462 ) , .ZN( us30_n747 ) );
  NAND2_X1 us30_U374 (.A1( us30_n462 ) , .A2( us30_n472 ) , .ZN( us30_n788 ) );
  NOR2_X1 us30_U375 (.ZN( us30_n465 ) , .A2( us30_n847 ) , .A1( us30_n848 ) );
  NOR2_X1 us30_U376 (.ZN( us30_n453 ) , .A1( us30_n826 ) , .A2( us30_n827 ) );
  NOR2_X1 us30_U377 (.ZN( us30_n451 ) , .A1( us30_n828 ) , .A2( us30_n829 ) );
  NAND2_X1 us30_U378 (.A1( us30_n451 ) , .A2( us30_n462 ) , .ZN( us30_n790 ) );
  NAND2_X1 us30_U379 (.A2( us30_n441 ) , .A1( us30_n447 ) , .ZN( us30_n784 ) );
  NOR4_X1 us30_U38 (.A3( us30_n521 ) , .A1( us30_n522 ) , .ZN( us30_n523 ) , .A2( us30_n673 ) , .A4( us30_n769 ) );
  NAND2_X1 us30_U380 (.A2( us30_n454 ) , .A1( us30_n455 ) , .ZN( us30_n730 ) );
  NAND2_X2 us30_U381 (.A1( us30_n449 ) , .A2( us30_n464 ) , .ZN( us30_n724 ) );
  NAND2_X2 us30_U382 (.A1( us30_n449 ) , .A2( us30_n460 ) , .ZN( us30_n792 ) );
  NAND2_X2 us30_U383 (.A2( us30_n460 ) , .A1( us30_n465 ) , .ZN( us30_n780 ) );
  NOR2_X1 us30_U384 (.ZN( us30_n447 ) , .A2( us30_n849 ) , .A1( us30_n858 ) );
  NAND2_X1 us30_U385 (.A1( us30_n447 ) , .A2( us30_n448 ) , .ZN( us30_n786 ) );
  NOR2_X1 us30_U386 (.A2( sa30_6 ) , .A1( sa30_7 ) , .ZN( us30_n464 ) );
  NOR2_X1 us30_U387 (.A2( sa30_7 ) , .ZN( us30_n460 ) , .A1( us30_n849 ) );
  NOR2_X1 us30_U388 (.A2( sa30_4 ) , .ZN( us30_n449 ) , .A1( us30_n848 ) );
  NOR2_X1 us30_U389 (.A2( sa30_4 ) , .A1( sa30_5 ) , .ZN( us30_n441 ) );
  AOI221_X1 us30_U39 (.A( us30_n781 ) , .ZN( us30_n798 ) , .C2( us30_n837 ) , .B2( us30_n838 ) , .B1( us30_n865 ) , .C1( us30_n866 ) );
  NOR2_X1 us30_U390 (.A2( sa30_5 ) , .ZN( us30_n448 ) , .A1( us30_n847 ) );
  NOR2_X1 us30_U391 (.A2( sa30_2 ) , .A1( sa30_3 ) , .ZN( us30_n472 ) );
  NOR2_X1 us30_U392 (.A2( sa30_6 ) , .ZN( us30_n452 ) , .A1( us30_n858 ) );
  NOR2_X1 us30_U393 (.A2( sa30_1 ) , .ZN( us30_n471 ) , .A1( us30_n826 ) );
  NOR2_X1 us30_U394 (.A2( sa30_0 ) , .ZN( us30_n454 ) , .A1( us30_n827 ) );
  NOR2_X1 us30_U395 (.A2( sa30_0 ) , .A1( sa30_1 ) , .ZN( us30_n462 ) );
  NOR2_X1 us30_U396 (.A2( sa30_3 ) , .ZN( us30_n455 ) , .A1( us30_n828 ) );
  NOR2_X1 us30_U397 (.A2( sa30_2 ) , .ZN( us30_n461 ) , .A1( us30_n829 ) );
  INV_X1 us30_U398 (.A( sa30_6 ) , .ZN( us30_n849 ) );
  INV_X1 us30_U399 (.A( sa30_4 ) , .ZN( us30_n847 ) );
  NAND2_X1 us30_U4 (.A1( us30_n441 ) , .A2( us30_n464 ) , .ZN( us30_n708 ) );
  NOR4_X1 us30_U40 (.A4( us30_n793 ) , .A3( us30_n794 ) , .A2( us30_n795 ) , .A1( us30_n796 ) , .ZN( us30_n797 ) );
  INV_X1 us30_U400 (.A( sa30_3 ) , .ZN( us30_n829 ) );
  INV_X1 us30_U401 (.A( sa30_1 ) , .ZN( us30_n827 ) );
  INV_X1 us30_U402 (.A( sa30_0 ) , .ZN( us30_n826 ) );
  INV_X1 us30_U403 (.A( sa30_2 ) , .ZN( us30_n828 ) );
  INV_X1 us30_U404 (.A( sa30_7 ) , .ZN( us30_n858 ) );
  INV_X1 us30_U405 (.A( sa30_5 ) , .ZN( us30_n848 ) );
  NAND2_X1 us30_U406 (.A2( us30_n461 ) , .A1( us30_n471 ) , .ZN( us30_n697 ) );
  OAI221_X1 us30_U407 (.A( us30_n783 ) , .C2( us30_n784 ) , .B2( us30_n785 ) , .B1( us30_n786 ) , .ZN( us30_n796 ) , .C1( us30_n813 ) );
  NAND2_X1 us30_U408 (.A1( us30_n729 ) , .A2( us30_n784 ) , .ZN( us30_n811 ) );
  OAI22_X1 us30_U409 (.ZN( us30_n588 ) , .A2( us30_n747 ) , .B2( us30_n762 ) , .A1( us30_n763 ) , .B1( us30_n784 ) );
  NOR4_X1 us30_U41 (.A4( us30_n776 ) , .A3( us30_n777 ) , .A1( us30_n778 ) , .ZN( us30_n799 ) , .A2( us30_n801 ) );
  AOI21_X1 us30_U410 (.ZN( us30_n592 ) , .B1( us30_n728 ) , .B2( us30_n784 ) , .A( us30_n790 ) );
  AOI21_X1 us30_U411 (.ZN( us30_n623 ) , .B1( us30_n699 ) , .A( us30_n779 ) , .B2( us30_n784 ) );
  AOI21_X1 us30_U412 (.ZN( us30_n648 ) , .A( us30_n762 ) , .B2( us30_n784 ) , .B1( us30_n792 ) );
  OAI22_X1 us30_U413 (.ZN( us30_n681 ) , .A1( us30_n699 ) , .A2( us30_n730 ) , .B2( us30_n784 ) , .B1( us30_n817 ) );
  OAI21_X1 us30_U414 (.A( us30_n613 ) , .ZN( us30_n616 ) , .B1( us30_n625 ) , .B2( us30_n784 ) );
  NOR2_X1 us30_U415 (.ZN( us30_n610 ) , .A1( us30_n784 ) , .A2( us30_n816 ) );
  OAI222_X1 us30_U416 (.A2( us30_n669 ) , .ZN( us30_n674 ) , .B1( us30_n747 ) , .B2( us30_n784 ) , .C2( us30_n788 ) , .C1( us30_n815 ) , .A1( us30_n817 ) );
  NOR2_X1 us30_U417 (.ZN( us30_n651 ) , .A1( us30_n784 ) , .A2( us30_n788 ) );
  NOR2_X1 us30_U418 (.ZN( us30_n600 ) , .A2( us30_n697 ) , .A1( us30_n784 ) );
  NOR2_X1 us30_U419 (.ZN( us30_n553 ) , .A2( us30_n744 ) , .A1( us30_n784 ) );
  NOR4_X1 us30_U42 (.A3( us30_n755 ) , .A2( us30_n756 ) , .A1( us30_n757 ) , .ZN( us30_n758 ) , .A4( us30_n869 ) );
  INV_X1 us30_U420 (.A( us30_n784 ) , .ZN( us30_n861 ) );
  AOI21_X1 us30_U421 (.ZN( us30_n500 ) , .A( us30_n697 ) , .B1( us30_n708 ) , .B2( us30_n786 ) );
  OAI221_X1 us30_U422 (.A( us30_n696 ) , .ZN( us30_n703 ) , .C2( us30_n784 ) , .C1( us30_n785 ) , .B1( us30_n786 ) , .B2( us30_n806 ) );
  OAI22_X1 us30_U423 (.ZN( us30_n590 ) , .B1( us30_n730 ) , .B2( us30_n749 ) , .A2( us30_n786 ) , .A1( us30_n803 ) );
  NOR2_X1 us30_U424 (.ZN( us30_n612 ) , .A1( us30_n779 ) , .A2( us30_n786 ) );
  NAND2_X1 us30_U425 (.A2( us30_n749 ) , .A1( us30_n786 ) , .ZN( us30_n809 ) );
  OAI222_X1 us30_U426 (.ZN( us30_n617 ) , .B1( us30_n697 ) , .C1( us30_n724 ) , .C2( us30_n747 ) , .B2( us30_n786 ) , .A2( us30_n792 ) , .A1( us30_n816 ) );
  NOR2_X1 us30_U427 (.ZN( us30_n717 ) , .A2( us30_n744 ) , .A1( us30_n786 ) );
  NOR2_X1 us30_U428 (.ZN( us30_n653 ) , .A1( us30_n762 ) , .A2( us30_n786 ) );
  NOR2_X1 us30_U429 (.ZN( us30_n554 ) , .A1( us30_n786 ) , .A2( us30_n813 ) );
  AOI211_X1 us30_U43 (.B( us30_n745 ) , .A( us30_n746 ) , .ZN( us30_n759 ) , .C1( us30_n832 ) , .C2( us30_n853 ) );
  NOR2_X1 us30_U430 (.ZN( us30_n701 ) , .A2( us30_n786 ) , .A1( us30_n817 ) );
  NOR2_X1 us30_U431 (.A1( us30_n730 ) , .ZN( us30_n765 ) , .A2( us30_n786 ) );
  AND2_X1 us30_U432 (.ZN( us30_n438 ) , .A2( us30_n831 ) , .A1( us30_n854 ) );
  AND2_X1 us30_U433 (.ZN( us30_n439 ) , .A2( us30_n843 ) , .A1( us30_n861 ) );
  NOR3_X1 us30_U434 (.A1( us30_n438 ) , .A2( us30_n439 ) , .A3( us30_n576 ) , .ZN( us30_n587 ) );
  NAND4_X1 us30_U435 (.ZN( sa31_sr_2 ) , .A4( us30_n643 ) , .A3( us30_n644 ) , .A2( us30_n645 ) , .A1( us30_n646 ) );
  INV_X1 us30_U436 (.A( us30_n812 ) , .ZN( us30_n854 ) );
  NAND3_X1 us30_U437 (.ZN( sa31_sr_6 ) , .A3( us30_n797 ) , .A2( us30_n798 ) , .A1( us30_n799 ) );
  NAND3_X1 us30_U438 (.ZN( sa31_sr_5 ) , .A3( us30_n758 ) , .A2( us30_n759 ) , .A1( us30_n760 ) );
  NAND3_X1 us30_U439 (.ZN( sa31_sr_4 ) , .A3( us30_n738 ) , .A2( us30_n739 ) , .A1( us30_n740 ) );
  NOR3_X1 us30_U44 (.A3( us30_n741 ) , .A2( us30_n742 ) , .A1( us30_n743 ) , .ZN( us30_n760 ) );
  NAND3_X1 us30_U440 (.A3( us30_n675 ) , .A2( us30_n676 ) , .A1( us30_n677 ) , .ZN( us30_n807 ) );
  NAND3_X1 us30_U441 (.ZN( us30_n638 ) , .A3( us30_n708 ) , .A2( us30_n724 ) , .A1( us30_n792 ) );
  NAND3_X1 us30_U442 (.A3( us30_n618 ) , .A2( us30_n619 ) , .A1( us30_n620 ) , .ZN( us30_n725 ) );
  NAND3_X1 us30_U443 (.A3( us30_n585 ) , .A2( us30_n586 ) , .A1( us30_n587 ) , .ZN( us30_n621 ) );
  NAND3_X1 us30_U444 (.ZN( us30_n565 ) , .A3( us30_n680 ) , .A2( us30_n750 ) , .A1( us30_n785 ) );
  NAND3_X1 us30_U445 (.A3( us30_n523 ) , .A2( us30_n524 ) , .A1( us30_n525 ) , .ZN( us30_n742 ) );
  NAND3_X1 us30_U446 (.A3( us30_n512 ) , .A1( us30_n513 ) , .ZN( us30_n608 ) , .A2( us30_n871 ) );
  NAND3_X1 us30_U447 (.A3( us30_n467 ) , .A2( us30_n468 ) , .A1( us30_n469 ) , .ZN( us30_n777 ) );
  INV_X1 us30_U448 (.A( us30_n803 ) , .ZN( us30_n843 ) );
  AOI21_X1 us30_U449 (.ZN( us30_n576 ) , .B2( us30_n724 ) , .B1( us30_n748 ) , .A( us30_n785 ) );
  NAND4_X1 us30_U45 (.ZN( sa31_sr_3 ) , .A4( us30_n704 ) , .A3( us30_n705 ) , .A2( us30_n706 ) , .A1( us30_n707 ) );
  NOR4_X1 us30_U46 (.A4( us30_n700 ) , .A3( us30_n701 ) , .A2( us30_n702 ) , .A1( us30_n703 ) , .ZN( us30_n704 ) );
  AOI211_X1 us30_U47 (.B( us30_n694 ) , .A( us30_n695 ) , .ZN( us30_n705 ) , .C2( us30_n831 ) , .C1( us30_n851 ) );
  NOR2_X1 us30_U48 (.ZN( us30_n707 ) , .A2( us30_n776 ) , .A1( us30_n800 ) );
  AOI222_X1 us30_U49 (.B2( us30_n638 ) , .ZN( us30_n644 ) , .B1( us30_n841 ) , .A1( us30_n842 ) , .C2( us30_n846 ) , .C1( us30_n863 ) , .A2( us30_n865 ) );
  NAND2_X1 us30_U5 (.A2( us30_n441 ) , .A1( us30_n452 ) , .ZN( us30_n791 ) );
  NOR4_X1 us30_U50 (.A4( us30_n639 ) , .A3( us30_n640 ) , .A2( us30_n641 ) , .A1( us30_n642 ) , .ZN( us30_n643 ) );
  NOR3_X1 us30_U51 (.A2( us30_n607 ) , .A1( us30_n608 ) , .ZN( us30_n646 ) , .A3( us30_n722 ) );
  NOR2_X1 us30_U52 (.ZN( us30_n804 ) , .A1( us30_n854 ) , .A2( us30_n861 ) );
  NAND4_X1 us30_U53 (.ZN( sa31_sr_7 ) , .A4( us30_n822 ) , .A3( us30_n823 ) , .A2( us30_n824 ) , .A1( us30_n825 ) );
  NOR4_X1 us30_U54 (.A4( us30_n818 ) , .A3( us30_n819 ) , .A2( us30_n820 ) , .A1( us30_n821 ) , .ZN( us30_n822 ) );
  AOI222_X1 us30_U55 (.C2( us30_n809 ) , .B2( us30_n810 ) , .A2( us30_n811 ) , .ZN( us30_n823 ) , .C1( us30_n832 ) , .A1( us30_n839 ) , .B1( us30_n853 ) );
  AOI211_X1 us30_U56 (.B( us30_n807 ) , .A( us30_n808 ) , .ZN( us30_n824 ) , .C1( us30_n842 ) , .C2( us30_n850 ) );
  NAND4_X1 us30_U57 (.ZN( sa31_sr_0 ) , .A4( us30_n501 ) , .A3( us30_n502 ) , .A2( us30_n503 ) , .A1( us30_n504 ) );
  AOI221_X1 us30_U58 (.A( us30_n497 ) , .ZN( us30_n502 ) , .B2( us30_n843 ) , .C1( us30_n846 ) , .C2( us30_n860 ) , .B1( us30_n862 ) );
  NOR4_X1 us30_U59 (.A4( us30_n498 ) , .A3( us30_n499 ) , .A2( us30_n500 ) , .ZN( us30_n501 ) , .A1( us30_n527 ) );
  NAND2_X1 us30_U6 (.A2( us30_n471 ) , .A1( us30_n472 ) , .ZN( us30_n817 ) );
  AOI211_X1 us30_U60 (.A( us30_n496 ) , .ZN( us30_n503 ) , .B( us30_n802 ) , .C2( us30_n839 ) , .C1( us30_n851 ) );
  NAND4_X1 us30_U61 (.ZN( sa31_sr_1 ) , .A4( us30_n595 ) , .A3( us30_n596 ) , .A2( us30_n597 ) , .A1( us30_n598 ) );
  NOR4_X1 us30_U62 (.A4( us30_n591 ) , .A3( us30_n592 ) , .A2( us30_n593 ) , .A1( us30_n594 ) , .ZN( us30_n595 ) );
  AOI211_X1 us30_U63 (.B( us30_n589 ) , .A( us30_n590 ) , .ZN( us30_n596 ) , .C2( us30_n811 ) , .C1( us30_n833 ) );
  AOI211_X1 us30_U64 (.A( us30_n588 ) , .ZN( us30_n597 ) , .B( us30_n621 ) , .C1( us30_n845 ) , .C2( us30_n855 ) );
  NOR2_X1 us30_U65 (.ZN( us30_n748 ) , .A1( us30_n861 ) , .A2( us30_n862 ) );
  NOR2_X1 us30_U66 (.ZN( us30_n625 ) , .A2( us30_n836 ) , .A1( us30_n839 ) );
  NAND4_X1 us30_U67 (.A4( us30_n603 ) , .A3( us30_n604 ) , .A2( us30_n605 ) , .A1( us30_n606 ) , .ZN( us30_n722 ) );
  NOR3_X1 us30_U68 (.A1( us30_n599 ) , .ZN( us30_n604 ) , .A3( us30_n663 ) , .A2( us30_n770 ) );
  NOR4_X1 us30_U69 (.A3( us30_n600 ) , .A2( us30_n601 ) , .A1( us30_n602 ) , .ZN( us30_n603 ) , .A4( us30_n655 ) );
  NOR3_X1 us30_U7 (.ZN( us30_n598 ) , .A1( us30_n608 ) , .A3( us30_n723 ) , .A2( us30_n742 ) );
  AOI222_X1 us30_U70 (.ZN( us30_n606 ) , .A1( us30_n830 ) , .C2( us30_n837 ) , .B1( us30_n842 ) , .A2( us30_n856 ) , .B2( us30_n861 ) , .C1( us30_n868 ) );
  NAND4_X1 us30_U71 (.A4( us30_n657 ) , .A3( us30_n658 ) , .A2( us30_n659 ) , .A1( us30_n660 ) , .ZN( us30_n800 ) );
  NOR3_X1 us30_U72 (.A3( us30_n648 ) , .A2( us30_n649 ) , .A1( us30_n650 ) , .ZN( us30_n659 ) );
  NOR3_X1 us30_U73 (.A3( us30_n651 ) , .A2( us30_n652 ) , .A1( us30_n653 ) , .ZN( us30_n658 ) );
  NOR3_X1 us30_U74 (.A3( us30_n654 ) , .A2( us30_n655 ) , .A1( us30_n656 ) , .ZN( us30_n657 ) );
  NAND4_X1 us30_U75 (.A4( us30_n560 ) , .A3( us30_n561 ) , .A2( us30_n562 ) , .A1( us30_n563 ) , .ZN( us30_n607 ) );
  NOR4_X1 us30_U76 (.ZN( us30_n561 ) , .A1( us30_n653 ) , .A3( us30_n661 ) , .A4( us30_n685 ) , .A2( us30_n768 ) );
  NOR4_X1 us30_U77 (.A4( us30_n552 ) , .A3( us30_n553 ) , .A2( us30_n554 ) , .A1( us30_n555 ) , .ZN( us30_n562 ) );
  NOR4_X1 us30_U78 (.A4( us30_n556 ) , .A3( us30_n557 ) , .A2( us30_n558 ) , .A1( us30_n559 ) , .ZN( us30_n560 ) );
  NAND4_X1 us30_U79 (.A4( us30_n772 ) , .A3( us30_n773 ) , .A2( us30_n774 ) , .A1( us30_n775 ) , .ZN( us30_n801 ) );
  NOR3_X1 us30_U8 (.A3( us30_n800 ) , .A2( us30_n801 ) , .A1( us30_n802 ) , .ZN( us30_n825 ) );
  NOR3_X1 us30_U80 (.A3( us30_n765 ) , .A2( us30_n766 ) , .A1( us30_n767 ) , .ZN( us30_n773 ) );
  NOR4_X1 us30_U81 (.A4( us30_n768 ) , .A3( us30_n769 ) , .A2( us30_n770 ) , .A1( us30_n771 ) , .ZN( us30_n772 ) );
  AOI222_X1 us30_U82 (.ZN( us30_n775 ) , .A1( us30_n830 ) , .C1( us30_n834 ) , .B2( us30_n841 ) , .A2( us30_n850 ) , .B1( us30_n861 ) , .C2( us30_n873 ) );
  NOR4_X1 us30_U83 (.A4( us30_n665 ) , .A3( us30_n666 ) , .A2( us30_n667 ) , .A1( us30_n668 ) , .ZN( us30_n676 ) );
  NOR4_X1 us30_U84 (.A4( us30_n661 ) , .A3( us30_n662 ) , .A2( us30_n663 ) , .A1( us30_n664 ) , .ZN( us30_n677 ) );
  NOR4_X1 us30_U85 (.A3( us30_n673 ) , .A1( us30_n674 ) , .ZN( us30_n675 ) , .A4( us30_n715 ) , .A2( us30_n859 ) );
  NOR2_X1 us30_U86 (.ZN( us30_n761 ) , .A1( us30_n833 ) , .A2( us30_n834 ) );
  NOR4_X1 us30_U87 (.A4( us30_n577 ) , .A3( us30_n578 ) , .A2( us30_n579 ) , .ZN( us30_n586 ) , .A1( us30_n683 ) );
  NOR4_X1 us30_U88 (.A1( us30_n584 ) , .ZN( us30_n585 ) , .A3( us30_n652 ) , .A2( us30_n662 ) , .A4( us30_n767 ) );
  AOI222_X1 us30_U89 (.ZN( us30_n513 ) , .C1( us30_n832 ) , .B2( us30_n837 ) , .A2( us30_n843 ) , .C2( us30_n862 ) , .B1( us30_n863 ) , .A1( us30_n866 ) );
  NOR3_X1 us30_U9 (.A3( us30_n621 ) , .A2( us30_n622 ) , .ZN( us30_n636 ) , .A1( us30_n725 ) );
  NOR4_X1 us30_U90 (.A4( us30_n509 ) , .A2( us30_n510 ) , .A1( us30_n511 ) , .ZN( us30_n512 ) , .A3( us30_n670 ) );
  INV_X1 us30_U91 (.A( us30_n505 ) , .ZN( us30_n871 ) );
  NAND4_X1 us30_U92 (.A4( us30_n456 ) , .A3( us30_n457 ) , .A2( us30_n458 ) , .A1( us30_n459 ) , .ZN( us30_n679 ) );
  NOR3_X1 us30_U93 (.ZN( us30_n457 ) , .A3( us30_n530 ) , .A1( us30_n555 ) , .A2( us30_n570 ) );
  AOI221_X1 us30_U94 (.A( us30_n450 ) , .ZN( us30_n459 ) , .C2( us30_n753 ) , .B1( us30_n832 ) , .C1( us30_n842 ) , .B2( us30_n861 ) );
  NOR4_X1 us30_U95 (.ZN( us30_n458 ) , .A2( us30_n509 ) , .A1( us30_n599 ) , .A4( us30_n628 ) , .A3( us30_n711 ) );
  NAND4_X1 us30_U96 (.A4( us30_n535 ) , .A3( us30_n536 ) , .A2( us30_n537 ) , .A1( us30_n538 ) , .ZN( us30_n622 ) );
  NOR4_X1 us30_U97 (.A4( us30_n526 ) , .A2( us30_n527 ) , .A1( us30_n528 ) , .ZN( us30_n538 ) , .A3( us30_n701 ) );
  NOR4_X1 us30_U98 (.A1( us30_n531 ) , .ZN( us30_n536 ) , .A2( us30_n654 ) , .A4( us30_n668 ) , .A3( us30_n765 ) );
  NOR4_X1 us30_U99 (.A4( us30_n529 ) , .A3( us30_n530 ) , .ZN( us30_n537 ) , .A2( us30_n684 ) , .A1( us30_n794 ) );
endmodule

