module aes_aes_die_21 ( w0_10, w0_12, w0_13, w0_14, w0_15, w3_0, w3_1, w3_2, w3_3, 
       w3_4, w3_5, w3_6, w3_7, u0_n33, u0_n35, u0_n37, u0_n39, u0_n43, u0_subword_11, u0_subword_8, u0_subword_9 );
  input w0_10, w0_12, w0_13, w0_14, w0_15, w3_0, w3_1, w3_2, w3_3, 
        w3_4, w3_5, w3_6, w3_7;
  output u0_n33, u0_n35, u0_n37, u0_n39, u0_n43, u0_subword_11, u0_subword_8, u0_subword_9;
  wire u0_subword_10, u0_subword_12, u0_subword_13, u0_subword_14, u0_subword_15, u0_u2_n438, u0_u2_n439, u0_u2_n440, u0_u2_n441, 
       u0_u2_n442, u0_u2_n443, u0_u2_n444, u0_u2_n445, u0_u2_n446, u0_u2_n447, u0_u2_n448, u0_u2_n449, u0_u2_n450, 
       u0_u2_n451, u0_u2_n452, u0_u2_n453, u0_u2_n454, u0_u2_n455, u0_u2_n456, u0_u2_n457, u0_u2_n458, u0_u2_n459, 
       u0_u2_n460, u0_u2_n461, u0_u2_n462, u0_u2_n463, u0_u2_n464, u0_u2_n465, u0_u2_n466, u0_u2_n467, u0_u2_n468, 
       u0_u2_n469, u0_u2_n470, u0_u2_n471, u0_u2_n472, u0_u2_n473, u0_u2_n474, u0_u2_n475, u0_u2_n476, u0_u2_n477, 
       u0_u2_n478, u0_u2_n479, u0_u2_n480, u0_u2_n481, u0_u2_n482, u0_u2_n483, u0_u2_n484, u0_u2_n485, u0_u2_n486, 
       u0_u2_n487, u0_u2_n488, u0_u2_n489, u0_u2_n490, u0_u2_n491, u0_u2_n492, u0_u2_n493, u0_u2_n494, u0_u2_n495, 
       u0_u2_n496, u0_u2_n497, u0_u2_n498, u0_u2_n499, u0_u2_n500, u0_u2_n501, u0_u2_n502, u0_u2_n503, u0_u2_n504, 
       u0_u2_n505, u0_u2_n506, u0_u2_n507, u0_u2_n508, u0_u2_n509, u0_u2_n510, u0_u2_n511, u0_u2_n512, u0_u2_n513, 
       u0_u2_n514, u0_u2_n515, u0_u2_n516, u0_u2_n517, u0_u2_n518, u0_u2_n519, u0_u2_n520, u0_u2_n521, u0_u2_n522, 
       u0_u2_n523, u0_u2_n524, u0_u2_n525, u0_u2_n526, u0_u2_n527, u0_u2_n528, u0_u2_n529, u0_u2_n530, u0_u2_n531, 
       u0_u2_n532, u0_u2_n533, u0_u2_n534, u0_u2_n535, u0_u2_n536, u0_u2_n537, u0_u2_n538, u0_u2_n539, u0_u2_n540, 
       u0_u2_n541, u0_u2_n542, u0_u2_n543, u0_u2_n544, u0_u2_n545, u0_u2_n546, u0_u2_n547, u0_u2_n548, u0_u2_n549, 
       u0_u2_n550, u0_u2_n551, u0_u2_n552, u0_u2_n553, u0_u2_n554, u0_u2_n555, u0_u2_n556, u0_u2_n557, u0_u2_n558, 
       u0_u2_n559, u0_u2_n560, u0_u2_n561, u0_u2_n562, u0_u2_n563, u0_u2_n564, u0_u2_n565, u0_u2_n566, u0_u2_n567, 
       u0_u2_n568, u0_u2_n569, u0_u2_n570, u0_u2_n571, u0_u2_n572, u0_u2_n573, u0_u2_n574, u0_u2_n575, u0_u2_n576, 
       u0_u2_n577, u0_u2_n578, u0_u2_n579, u0_u2_n580, u0_u2_n581, u0_u2_n582, u0_u2_n583, u0_u2_n584, u0_u2_n585, 
       u0_u2_n586, u0_u2_n587, u0_u2_n588, u0_u2_n589, u0_u2_n590, u0_u2_n591, u0_u2_n592, u0_u2_n593, u0_u2_n594, 
       u0_u2_n595, u0_u2_n596, u0_u2_n597, u0_u2_n598, u0_u2_n599, u0_u2_n600, u0_u2_n601, u0_u2_n602, u0_u2_n603, 
       u0_u2_n604, u0_u2_n605, u0_u2_n606, u0_u2_n607, u0_u2_n608, u0_u2_n609, u0_u2_n610, u0_u2_n611, u0_u2_n612, 
       u0_u2_n613, u0_u2_n614, u0_u2_n615, u0_u2_n616, u0_u2_n617, u0_u2_n618, u0_u2_n619, u0_u2_n620, u0_u2_n621, 
       u0_u2_n622, u0_u2_n623, u0_u2_n624, u0_u2_n625, u0_u2_n626, u0_u2_n627, u0_u2_n628, u0_u2_n629, u0_u2_n630, 
       u0_u2_n631, u0_u2_n632, u0_u2_n633, u0_u2_n634, u0_u2_n635, u0_u2_n636, u0_u2_n637, u0_u2_n638, u0_u2_n639, 
       u0_u2_n640, u0_u2_n641, u0_u2_n642, u0_u2_n643, u0_u2_n644, u0_u2_n645, u0_u2_n646, u0_u2_n647, u0_u2_n648, 
       u0_u2_n649, u0_u2_n650, u0_u2_n651, u0_u2_n652, u0_u2_n653, u0_u2_n654, u0_u2_n655, u0_u2_n656, u0_u2_n657, 
       u0_u2_n658, u0_u2_n659, u0_u2_n660, u0_u2_n661, u0_u2_n662, u0_u2_n663, u0_u2_n664, u0_u2_n665, u0_u2_n666, 
       u0_u2_n667, u0_u2_n668, u0_u2_n669, u0_u2_n670, u0_u2_n671, u0_u2_n672, u0_u2_n673, u0_u2_n674, u0_u2_n675, 
       u0_u2_n676, u0_u2_n677, u0_u2_n678, u0_u2_n679, u0_u2_n680, u0_u2_n681, u0_u2_n682, u0_u2_n683, u0_u2_n684, 
       u0_u2_n685, u0_u2_n686, u0_u2_n687, u0_u2_n688, u0_u2_n689, u0_u2_n690, u0_u2_n691, u0_u2_n692, u0_u2_n693, 
       u0_u2_n694, u0_u2_n695, u0_u2_n696, u0_u2_n697, u0_u2_n698, u0_u2_n699, u0_u2_n700, u0_u2_n701, u0_u2_n702, 
       u0_u2_n703, u0_u2_n704, u0_u2_n705, u0_u2_n706, u0_u2_n707, u0_u2_n708, u0_u2_n709, u0_u2_n710, u0_u2_n711, 
       u0_u2_n712, u0_u2_n713, u0_u2_n714, u0_u2_n715, u0_u2_n716, u0_u2_n717, u0_u2_n718, u0_u2_n719, u0_u2_n720, 
       u0_u2_n721, u0_u2_n722, u0_u2_n723, u0_u2_n724, u0_u2_n725, u0_u2_n726, u0_u2_n727, u0_u2_n728, u0_u2_n729, 
       u0_u2_n730, u0_u2_n731, u0_u2_n732, u0_u2_n733, u0_u2_n734, u0_u2_n735, u0_u2_n736, u0_u2_n737, u0_u2_n738, 
       u0_u2_n739, u0_u2_n740, u0_u2_n741, u0_u2_n742, u0_u2_n743, u0_u2_n744, u0_u2_n745, u0_u2_n746, u0_u2_n747, 
       u0_u2_n748, u0_u2_n749, u0_u2_n750, u0_u2_n751, u0_u2_n752, u0_u2_n753, u0_u2_n754, u0_u2_n755, u0_u2_n756, 
       u0_u2_n757, u0_u2_n758, u0_u2_n759, u0_u2_n760, u0_u2_n761, u0_u2_n762, u0_u2_n763, u0_u2_n764, u0_u2_n765, 
       u0_u2_n766, u0_u2_n767, u0_u2_n768, u0_u2_n769, u0_u2_n770, u0_u2_n771, u0_u2_n772, u0_u2_n773, u0_u2_n774, 
       u0_u2_n775, u0_u2_n776, u0_u2_n777, u0_u2_n778, u0_u2_n779, u0_u2_n780, u0_u2_n781, u0_u2_n782, u0_u2_n783, 
       u0_u2_n784, u0_u2_n785, u0_u2_n786, u0_u2_n787, u0_u2_n788, u0_u2_n789, u0_u2_n790, u0_u2_n791, u0_u2_n792, 
       u0_u2_n793, u0_u2_n794, u0_u2_n795, u0_u2_n796, u0_u2_n797, u0_u2_n798, u0_u2_n799, u0_u2_n800, u0_u2_n801, 
       u0_u2_n802, u0_u2_n803, u0_u2_n804, u0_u2_n805, u0_u2_n806, u0_u2_n807, u0_u2_n808, u0_u2_n809, u0_u2_n810, 
       u0_u2_n811, u0_u2_n812, u0_u2_n813, u0_u2_n814, u0_u2_n815, u0_u2_n816, u0_u2_n817, u0_u2_n818, u0_u2_n819, 
       u0_u2_n820, u0_u2_n821, u0_u2_n822, u0_u2_n823, u0_u2_n824, u0_u2_n825, u0_u2_n826, u0_u2_n827, u0_u2_n828, 
       u0_u2_n829, u0_u2_n830, u0_u2_n831, u0_u2_n832, u0_u2_n833, u0_u2_n834, u0_u2_n835, u0_u2_n836, u0_u2_n837, 
       u0_u2_n838, u0_u2_n839, u0_u2_n840, u0_u2_n841, u0_u2_n842, u0_u2_n843, u0_u2_n844, u0_u2_n845, u0_u2_n846, 
       u0_u2_n847, u0_u2_n848, u0_u2_n849, u0_u2_n850, u0_u2_n851, u0_u2_n852, u0_u2_n853, u0_u2_n854, u0_u2_n855, 
       u0_u2_n856, u0_u2_n857, u0_u2_n858, u0_u2_n859, u0_u2_n860, u0_u2_n861, u0_u2_n862, u0_u2_n863, u0_u2_n864, 
       u0_u2_n865, u0_u2_n866, u0_u2_n867, u0_u2_n868, u0_u2_n869, u0_u2_n870, u0_u2_n871, u0_u2_n872, u0_u2_n873, 
       u0_u2_n874, u0_u2_n875, u0_u2_n876, u0_u2_n877, u0_u2_n878, u0_u2_n879, u0_u2_n880, u0_u2_n881, u0_u2_n882, 
        u0_u2_n883;
  XNOR2_X1 u0_U12 (.ZN( u0_n33 ) , .B( u0_subword_15 ) , .A( w0_15 ) );
  XNOR2_X1 u0_U16 (.ZN( u0_n37 ) , .B( u0_subword_13 ) , .A( w0_13 ) );
  XNOR2_X1 u0_U211 (.ZN( u0_n43 ) , .B( u0_subword_10 ) , .A( w0_10 ) );
  XNOR2_X1 u0_U23 (.ZN( u0_n39 ) , .B( u0_subword_12 ) , .A( w0_12 ) );
  XNOR2_X1 u0_U240 (.ZN( u0_n35 ) , .B( u0_subword_14 ) , .A( w0_14 ) );
  NOR2_X1 u0_u2_U10 (.ZN( u0_u2_n714 ) , .A2( u0_u2_n783 ) , .A1( u0_u2_n807 ) );
  OR4_X1 u0_u2_U100 (.ZN( u0_u2_n473 ) , .A4( u0_u2_n525 ) , .A3( u0_u2_n536 ) , .A2( u0_u2_n585 ) , .A1( u0_u2_n719 ) );
  NOR4_X1 u0_u2_U101 (.A4( u0_u2_n584 ) , .A3( u0_u2_n585 ) , .A2( u0_u2_n586 ) , .ZN( u0_u2_n593 ) , .A1( u0_u2_n690 ) );
  NOR4_X1 u0_u2_U102 (.A1( u0_u2_n591 ) , .ZN( u0_u2_n592 ) , .A3( u0_u2_n659 ) , .A2( u0_u2_n669 ) , .A4( u0_u2_n774 ) );
  OR4_X1 u0_u2_U103 (.ZN( u0_u2_n499 ) , .A4( u0_u2_n541 ) , .A2( u0_u2_n554 ) , .A1( u0_u2_n566 ) , .A3( u0_u2_n639 ) );
  OR3_X1 u0_u2_U104 (.A3( u0_u2_n513 ) , .A2( u0_u2_n514 ) , .A1( u0_u2_n515 ) , .ZN( u0_u2_n518 ) );
  AOI21_X1 u0_u2_U105 (.A( u0_u2_n677 ) , .B1( u0_u2_n678 ) , .ZN( u0_u2_n679 ) , .B2( u0_u2_n863 ) );
  INV_X1 u0_u2_U106 (.A( u0_u2_n761 ) , .ZN( u0_u2_n876 ) );
  OAI21_X1 u0_u2_U107 (.B1( u0_u2_n760 ) , .ZN( u0_u2_n761 ) , .A( u0_u2_n852 ) , .B2( u0_u2_n875 ) );
  AOI221_X1 u0_u2_U108 (.A( u0_u2_n720 ) , .B2( u0_u2_n721 ) , .ZN( u0_u2_n727 ) , .C1( u0_u2_n839 ) , .B1( u0_u2_n846 ) , .C2( u0_u2_n870 ) );
  OR2_X1 u0_u2_U109 (.A2( u0_u2_n718 ) , .A1( u0_u2_n719 ) , .ZN( u0_u2_n720 ) );
  INV_X1 u0_u2_U11 (.A( u0_u2_n785 ) , .ZN( u0_u2_n874 ) );
  INV_X1 u0_u2_U110 (.A( u0_u2_n470 ) , .ZN( u0_u2_n871 ) );
  OAI21_X1 u0_u2_U111 (.ZN( u0_u2_n470 ) , .B1( u0_u2_n816 ) , .A( u0_u2_n841 ) , .B2( u0_u2_n858 ) );
  NAND2_X1 u0_u2_U112 (.ZN( u0_u2_n439 ) , .A2( u0_u2_n850 ) , .A1( u0_u2_n868 ) );
  NAND2_X1 u0_u2_U113 (.ZN( u0_u2_n440 ) , .A2( u0_u2_n838 ) , .A1( u0_u2_n861 ) );
  AOI221_X1 u0_u2_U114 (.A( u0_u2_n771 ) , .ZN( u0_u2_n781 ) , .C2( u0_u2_n817 ) , .B2( u0_u2_n842 ) , .C1( u0_u2_n862 ) , .B1( u0_u2_n873 ) );
  INV_X1 u0_u2_U115 (.A( u0_u2_n768 ) , .ZN( u0_u2_n842 ) );
  NAND2_X1 u0_u2_U116 (.A1( u0_u2_n454 ) , .A2( u0_u2_n472 ) , .ZN( u0_u2_n756 ) );
  AOI211_X1 u0_u2_U117 (.B( u0_u2_n814 ) , .A( u0_u2_n815 ) , .ZN( u0_u2_n831 ) , .C1( u0_u2_n849 ) , .C2( u0_u2_n857 ) );
  AOI211_X1 u0_u2_U118 (.A( u0_u2_n595 ) , .ZN( u0_u2_n604 ) , .B( u0_u2_n628 ) , .C1( u0_u2_n852 ) , .C2( u0_u2_n862 ) );
  INV_X1 u0_u2_U119 (.A( u0_u2_n737 ) , .ZN( u0_u2_n846 ) );
  INV_X1 u0_u2_U12 (.A( u0_u2_n686 ) , .ZN( u0_u2_n879 ) );
  NAND2_X1 u0_u2_U120 (.A1( u0_u2_n458 ) , .A2( u0_u2_n460 ) , .ZN( u0_u2_n769 ) );
  NOR3_X1 u0_u2_U121 (.ZN( u0_u2_n497 ) , .A1( u0_u2_n789 ) , .A2( u0_u2_n857 ) , .A3( u0_u2_n870 ) );
  OAI22_X1 u0_u2_U122 (.B2( u0_u2_n757 ) , .B1( u0_u2_n758 ) , .A1( u0_u2_n759 ) , .ZN( u0_u2_n763 ) , .A2( u0_u2_n813 ) );
  NOR2_X1 u0_u2_U123 (.ZN( u0_u2_n758 ) , .A2( u0_u2_n859 ) , .A1( u0_u2_n867 ) );
  NOR3_X1 u0_u2_U124 (.ZN( u0_u2_n759 ) , .A2( u0_u2_n860 ) , .A1( u0_u2_n870 ) , .A3( u0_u2_n872 ) );
  NOR2_X1 u0_u2_U125 (.ZN( u0_u2_n539 ) , .A2( u0_u2_n756 ) , .A1( u0_u2_n757 ) );
  NOR2_X1 u0_u2_U126 (.ZN( u0_u2_n577 ) , .A1( u0_u2_n735 ) , .A2( u0_u2_n813 ) );
  OAI21_X1 u0_u2_U127 (.ZN( u0_u2_n794 ) , .A( u0_u2_n846 ) , .B1( u0_u2_n870 ) , .B2( u0_u2_n880 ) );
  NOR2_X1 u0_u2_U128 (.A2( u0_u2_n715 ) , .A1( u0_u2_n757 ) , .ZN( u0_u2_n778 ) );
  NOR2_X1 u0_u2_U129 (.ZN( u0_u2_n516 ) , .A1( u0_u2_n736 ) , .A2( u0_u2_n786 ) );
  INV_X1 u0_u2_U13 (.A( u0_u2_n687 ) , .ZN( u0_u2_n847 ) );
  NOR2_X1 u0_u2_U130 (.ZN( u0_u2_n553 ) , .A2( u0_u2_n787 ) , .A1( u0_u2_n821 ) );
  NOR2_X1 u0_u2_U131 (.ZN( u0_u2_n618 ) , .A2( u0_u2_n787 ) , .A1( u0_u2_n813 ) );
  NOR2_X1 u0_u2_U132 (.ZN( u0_u2_n514 ) , .A1( u0_u2_n819 ) , .A2( u0_u2_n824 ) );
  NOR2_X1 u0_u2_U133 (.A2( u0_u2_n715 ) , .A1( u0_u2_n769 ) , .ZN( u0_u2_n801 ) );
  NOR2_X1 u0_u2_U134 (.ZN( u0_u2_n663 ) , .A1( u0_u2_n754 ) , .A2( u0_u2_n787 ) );
  NOR2_X1 u0_u2_U135 (.ZN( u0_u2_n513 ) , .A2( u0_u2_n735 ) , .A1( u0_u2_n769 ) );
  INV_X1 u0_u2_U136 (.A( u0_u2_n754 ) , .ZN( u0_u2_n841 ) );
  NOR2_X1 u0_u2_U137 (.ZN( u0_u2_n689 ) , .A2( u0_u2_n715 ) , .A1( u0_u2_n824 ) );
  INV_X1 u0_u2_U138 (.A( u0_u2_n735 ) , .ZN( u0_u2_n859 ) );
  AOI21_X1 u0_u2_U139 (.B1( u0_u2_n706 ) , .ZN( u0_u2_n707 ) , .A( u0_u2_n739 ) , .B2( u0_u2_n770 ) );
  AOI222_X1 u0_u2_U14 (.ZN( u0_u2_n570 ) , .B1( u0_u2_n837 ) , .C1( u0_u2_n848 ) , .A2( u0_u2_n850 ) , .A1( u0_u2_n861 ) , .B2( u0_u2_n870 ) , .C2( u0_u2_n880 ) );
  INV_X1 u0_u2_U140 (.A( u0_u2_n757 ) , .ZN( u0_u2_n849 ) );
  AOI21_X1 u0_u2_U141 (.ZN( u0_u2_n547 ) , .A( u0_u2_n770 ) , .B2( u0_u2_n786 ) , .B1( u0_u2_n824 ) );
  AOI21_X1 u0_u2_U142 (.ZN( u0_u2_n576 ) , .B1( u0_u2_n757 ) , .B2( u0_u2_n769 ) , .A( u0_u2_n787 ) );
  AOI21_X1 u0_u2_U143 (.B1( u0_u2_n693 ) , .ZN( u0_u2_n694 ) , .A( u0_u2_n735 ) , .B2( u0_u2_n768 ) );
  NOR2_X1 u0_u2_U144 (.ZN( u0_u2_n575 ) , .A1( u0_u2_n736 ) , .A2( u0_u2_n769 ) );
  NOR2_X1 u0_u2_U145 (.ZN( u0_u2_n536 ) , .A1( u0_u2_n715 ) , .A2( u0_u2_n786 ) );
  AOI21_X1 u0_u2_U146 (.ZN( u0_u2_n696 ) , .B2( u0_u2_n756 ) , .B1( u0_u2_n770 ) , .A( u0_u2_n813 ) );
  NOR2_X1 u0_u2_U147 (.ZN( u0_u2_n718 ) , .A1( u0_u2_n769 ) , .A2( u0_u2_n770 ) );
  INV_X1 u0_u2_U148 (.A( u0_u2_n787 ) , .ZN( u0_u2_n857 ) );
  NOR2_X1 u0_u2_U149 (.ZN( u0_u2_n621 ) , .A1( u0_u2_n769 ) , .A2( u0_u2_n819 ) );
  AOI222_X1 u0_u2_U15 (.ZN( u0_u2_n667 ) , .A2( u0_u2_n846 ) , .B1( u0_u2_n848 ) , .C2( u0_u2_n852 ) , .A1( u0_u2_n867 ) , .C1( u0_u2_n870 ) , .B2( u0_u2_n877 ) );
  AOI21_X1 u0_u2_U150 (.B1( u0_u2_n444 ) , .ZN( u0_u2_n634 ) , .A( u0_u2_n770 ) , .B2( u0_u2_n821 ) );
  INV_X1 u0_u2_U151 (.A( u0_u2_n736 ) , .ZN( u0_u2_n875 ) );
  NOR2_X1 u0_u2_U152 (.ZN( u0_u2_n527 ) , .A2( u0_u2_n715 ) , .A1( u0_u2_n821 ) );
  NOR2_X1 u0_u2_U153 (.ZN( u0_u2_n584 ) , .A2( u0_u2_n706 ) , .A1( u0_u2_n821 ) );
  INV_X1 u0_u2_U154 (.A( u0_u2_n706 ) , .ZN( u0_u2_n860 ) );
  OAI21_X1 u0_u2_U155 (.A( u0_u2_n705 ) , .ZN( u0_u2_n709 ) , .B2( u0_u2_n757 ) , .B1( u0_u2_n811 ) );
  OAI21_X1 u0_u2_U156 (.ZN( u0_u2_n705 ) , .B2( u0_u2_n840 ) , .B1( u0_u2_n845 ) , .A( u0_u2_n867 ) );
  INV_X1 u0_u2_U157 (.A( u0_u2_n770 ) , .ZN( u0_u2_n873 ) );
  NAND2_X1 u0_u2_U158 (.A1( u0_u2_n706 ) , .A2( u0_u2_n736 ) , .ZN( u0_u2_n789 ) );
  BUF_X1 u0_u2_U159 (.Z( u0_u2_n443 ) , .A( u0_u2_n822 ) );
  INV_X1 u0_u2_U16 (.A( u0_u2_n654 ) , .ZN( u0_u2_n877 ) );
  INV_X1 u0_u2_U160 (.A( u0_u2_n824 ) , .ZN( u0_u2_n851 ) );
  NAND2_X1 u0_u2_U161 (.ZN( u0_u2_n721 ) , .A1( u0_u2_n735 ) , .A2( u0_u2_n787 ) );
  BUF_X1 u0_u2_U162 (.Z( u0_u2_n442 ) , .A( u0_u2_n676 ) );
  BUF_X1 u0_u2_U163 (.Z( u0_u2_n441 ) , .A( u0_u2_n704 ) );
  OR4_X1 u0_u2_U164 (.A3( u0_u2_n587 ) , .A4( u0_u2_n588 ) , .A2( u0_u2_n589 ) , .A1( u0_u2_n590 ) , .ZN( u0_u2_n591 ) );
  OAI222_X1 u0_u2_U165 (.A2( u0_u2_n443 ) , .B2( u0_u2_n715 ) , .ZN( u0_u2_n716 ) , .C2( u0_u2_n731 ) , .B1( u0_u2_n754 ) , .A1( u0_u2_n813 ) , .C1( u0_u2_n821 ) );
  AOI221_X1 u0_u2_U166 (.A( u0_u2_n457 ) , .ZN( u0_u2_n466 ) , .C2( u0_u2_n760 ) , .B1( u0_u2_n839 ) , .C1( u0_u2_n849 ) , .B2( u0_u2_n868 ) );
  OAI221_X1 u0_u2_U167 (.A( u0_u2_n790 ) , .C2( u0_u2_n791 ) , .B2( u0_u2_n792 ) , .B1( u0_u2_n793 ) , .ZN( u0_u2_n803 ) , .C1( u0_u2_n820 ) );
  OAI221_X1 u0_u2_U168 (.A( u0_u2_n703 ) , .ZN( u0_u2_n710 ) , .C2( u0_u2_n791 ) , .C1( u0_u2_n792 ) , .B1( u0_u2_n793 ) , .B2( u0_u2_n813 ) );
  AOI22_X1 u0_u2_U169 (.ZN( u0_u2_n703 ) , .A1( u0_u2_n837 ) , .B2( u0_u2_n850 ) , .A2( u0_u2_n872 ) , .B1( u0_u2_n875 ) );
  NOR4_X1 u0_u2_U17 (.A4( u0_u2_n551 ) , .A3( u0_u2_n552 ) , .A2( u0_u2_n553 ) , .A1( u0_u2_n554 ) , .ZN( u0_u2_n555 ) );
  OAI221_X1 u0_u2_U170 (.A( u0_u2_n734 ) , .C2( u0_u2_n735 ) , .B2( u0_u2_n736 ) , .B1( u0_u2_n737 ) , .ZN( u0_u2_n744 ) , .C1( u0_u2_n824 ) );
  NAND2_X1 u0_u2_U171 (.A2( u0_u2_n467 ) , .A1( u0_u2_n472 ) , .ZN( u0_u2_n787 ) );
  NAND2_X1 u0_u2_U172 (.A2( u0_u2_n478 ) , .A1( u0_u2_n479 ) , .ZN( u0_u2_n824 ) );
  NAND2_X1 u0_u2_U173 (.A1( u0_u2_n456 ) , .A2( u0_u2_n467 ) , .ZN( u0_u2_n799 ) );
  NAND2_X1 u0_u2_U174 (.A2( u0_u2_n455 ) , .A1( u0_u2_n467 ) , .ZN( u0_u2_n735 ) );
  NAND2_X1 u0_u2_U175 (.A2( u0_u2_n456 ) , .A1( u0_u2_n459 ) , .ZN( u0_u2_n770 ) );
  NAND2_X1 u0_u2_U176 (.A2( u0_u2_n461 ) , .A1( u0_u2_n479 ) , .ZN( u0_u2_n786 ) );
  NAND2_X1 u0_u2_U177 (.A1( u0_u2_n448 ) , .A2( u0_u2_n467 ) , .ZN( u0_u2_n706 ) );
  NAND2_X1 u0_u2_U178 (.A1( u0_u2_n460 ) , .A2( u0_u2_n479 ) , .ZN( u0_u2_n792 ) );
  NAND2_X1 u0_u2_U179 (.A2( u0_u2_n455 ) , .A1( u0_u2_n459 ) , .ZN( u0_u2_n736 ) );
  NOR4_X1 u0_u2_U18 (.A4( u0_u2_n539 ) , .A3( u0_u2_n540 ) , .A2( u0_u2_n541 ) , .ZN( u0_u2_n542 ) , .A1( u0_u2_n827 ) );
  NAND2_X1 u0_u2_U180 (.A2( u0_u2_n471 ) , .A1( u0_u2_n472 ) , .ZN( u0_u2_n819 ) );
  NAND2_X1 u0_u2_U181 (.A1( u0_u2_n462 ) , .A2( u0_u2_n478 ) , .ZN( u0_u2_n810 ) );
  NAND2_X1 u0_u2_U182 (.A1( u0_u2_n458 ) , .A2( u0_u2_n478 ) , .ZN( u0_u2_n823 ) );
  NAND2_X1 u0_u2_U183 (.A2( u0_u2_n448 ) , .A1( u0_u2_n454 ) , .ZN( u0_u2_n791 ) );
  NAND2_X1 u0_u2_U184 (.A1( u0_u2_n461 ) , .A2( u0_u2_n468 ) , .ZN( u0_u2_n820 ) );
  NOR2_X1 u0_u2_U185 (.ZN( u0_u2_n460 ) , .A1( u0_u2_n833 ) , .A2( u0_u2_n834 ) );
  NAND2_X1 u0_u2_U186 (.A2( u0_u2_n468 ) , .A1( u0_u2_n469 ) , .ZN( u0_u2_n754 ) );
  NAND2_X1 u0_u2_U187 (.A1( u0_u2_n454 ) , .A2( u0_u2_n455 ) , .ZN( u0_u2_n793 ) );
  NAND2_X1 u0_u2_U188 (.A1( u0_u2_n448 ) , .A2( u0_u2_n471 ) , .ZN( u0_u2_n715 ) );
  NAND2_X1 u0_u2_U189 (.A1( u0_u2_n469 ) , .A2( u0_u2_n479 ) , .ZN( u0_u2_n795 ) );
  NOR4_X1 u0_u2_U19 (.A4( u0_u2_n452 ) , .A3( u0_u2_n453 ) , .A2( u0_u2_n523 ) , .A1( u0_u2_n548 ) , .ZN( u0_u2_n713 ) );
  NAND2_X1 u0_u2_U190 (.A2( u0_u2_n448 ) , .A1( u0_u2_n459 ) , .ZN( u0_u2_n798 ) );
  NAND2_X1 u0_u2_U191 (.A1( u0_u2_n458 ) , .A2( u0_u2_n469 ) , .ZN( u0_u2_n797 ) );
  NAND2_X1 u0_u2_U192 (.A2( u0_u2_n461 ) , .A1( u0_u2_n462 ) , .ZN( u0_u2_n737 ) );
  AOI222_X1 u0_u2_U193 (.B2( u0_u2_n645 ) , .ZN( u0_u2_n651 ) , .B1( u0_u2_n848 ) , .A1( u0_u2_n849 ) , .C2( u0_u2_n853 ) , .C1( u0_u2_n870 ) , .A2( u0_u2_n872 ) );
  NOR4_X1 u0_u2_U194 (.A4( u0_u2_n646 ) , .A3( u0_u2_n647 ) , .A2( u0_u2_n648 ) , .A1( u0_u2_n649 ) , .ZN( u0_u2_n650 ) );
  NAND4_X1 u0_u2_U195 (.ZN( u0_subword_8 ) , .A4( u0_u2_n508 ) , .A3( u0_u2_n509 ) , .A2( u0_u2_n510 ) , .A1( u0_u2_n511 ) );
  NOR4_X1 u0_u2_U196 (.A4( u0_u2_n505 ) , .A3( u0_u2_n506 ) , .A2( u0_u2_n507 ) , .ZN( u0_u2_n508 ) , .A1( u0_u2_n534 ) );
  AOI221_X1 u0_u2_U197 (.A( u0_u2_n504 ) , .ZN( u0_u2_n509 ) , .B2( u0_u2_n850 ) , .C1( u0_u2_n853 ) , .C2( u0_u2_n867 ) , .B1( u0_u2_n869 ) );
  AOI221_X1 u0_u2_U198 (.A( u0_u2_n788 ) , .ZN( u0_u2_n805 ) , .C2( u0_u2_n844 ) , .B2( u0_u2_n845 ) , .B1( u0_u2_n872 ) , .C1( u0_u2_n873 ) );
  NOR4_X1 u0_u2_U199 (.A4( u0_u2_n800 ) , .A3( u0_u2_n801 ) , .A2( u0_u2_n802 ) , .A1( u0_u2_n803 ) , .ZN( u0_u2_n804 ) );
  OR4_X1 u0_u2_U20 (.A4( u0_u2_n449 ) , .A2( u0_u2_n450 ) , .A1( u0_u2_n451 ) , .ZN( u0_u2_n452 ) , .A3( u0_u2_n560 ) );
  NOR4_X1 u0_u2_U200 (.A4( u0_u2_n707 ) , .A3( u0_u2_n708 ) , .A2( u0_u2_n709 ) , .A1( u0_u2_n710 ) , .ZN( u0_u2_n711 ) );
  AOI211_X1 u0_u2_U201 (.B( u0_u2_n701 ) , .A( u0_u2_n702 ) , .ZN( u0_u2_n712 ) , .C2( u0_u2_n838 ) , .C1( u0_u2_n858 ) );
  NAND4_X1 u0_u2_U202 (.ZN( u0_subword_15 ) , .A4( u0_u2_n829 ) , .A3( u0_u2_n830 ) , .A2( u0_u2_n831 ) , .A1( u0_u2_n832 ) );
  NOR4_X1 u0_u2_U203 (.A4( u0_u2_n825 ) , .A3( u0_u2_n826 ) , .A2( u0_u2_n827 ) , .A1( u0_u2_n828 ) , .ZN( u0_u2_n829 ) );
  NAND4_X1 u0_u2_U204 (.ZN( u0_subword_9 ) , .A4( u0_u2_n602 ) , .A3( u0_u2_n603 ) , .A2( u0_u2_n604 ) , .A1( u0_u2_n605 ) );
  NOR4_X1 u0_u2_U205 (.A4( u0_u2_n598 ) , .A3( u0_u2_n599 ) , .A2( u0_u2_n600 ) , .A1( u0_u2_n601 ) , .ZN( u0_u2_n602 ) );
  AOI211_X1 u0_u2_U206 (.B( u0_u2_n596 ) , .A( u0_u2_n597 ) , .ZN( u0_u2_n603 ) , .C2( u0_u2_n818 ) , .C1( u0_u2_n840 ) );
  NOR4_X1 u0_u2_U207 (.A3( u0_u2_n762 ) , .A2( u0_u2_n763 ) , .A1( u0_u2_n764 ) , .ZN( u0_u2_n765 ) , .A4( u0_u2_n876 ) );
  AOI211_X1 u0_u2_U208 (.B( u0_u2_n752 ) , .A( u0_u2_n753 ) , .ZN( u0_u2_n766 ) , .C1( u0_u2_n839 ) , .C2( u0_u2_n860 ) );
  NOR4_X1 u0_u2_U209 (.A4( u0_u2_n741 ) , .A3( u0_u2_n742 ) , .A2( u0_u2_n743 ) , .A1( u0_u2_n744 ) , .ZN( u0_u2_n745 ) );
  INV_X1 u0_u2_U21 (.A( u0_u2_n620 ) , .ZN( u0_u2_n882 ) );
  AOI211_X1 u0_u2_U210 (.B( u0_u2_n732 ) , .A( u0_u2_n733 ) , .ZN( u0_u2_n746 ) , .C1( u0_u2_n850 ) , .C2( u0_u2_n862 ) );
  AOI221_X1 u0_u2_U211 (.ZN( u0_u2_n475 ) , .C2( u0_u2_n721 ) , .B2( u0_u2_n838 ) , .C1( u0_u2_n852 ) , .B1( u0_u2_n867 ) , .A( u0_u2_n871 ) );
  AOI22_X1 u0_u2_U212 (.A2( u0_u2_n789 ) , .ZN( u0_u2_n790 ) , .B2( u0_u2_n838 ) , .A1( u0_u2_n841 ) , .B1( u0_u2_n870 ) );
  NAND2_X1 u0_u2_U213 (.A1( u0_u2_n460 ) , .A2( u0_u2_n468 ) , .ZN( u0_u2_n751 ) );
  NAND2_X1 u0_u2_U214 (.A1( u0_u2_n454 ) , .A2( u0_u2_n456 ) , .ZN( u0_u2_n812 ) );
  NAND2_X1 u0_u2_U215 (.A2( u0_u2_n460 ) , .A1( u0_u2_n462 ) , .ZN( u0_u2_n813 ) );
  NAND2_X1 u0_u2_U216 (.A1( u0_u2_n456 ) , .A2( u0_u2_n471 ) , .ZN( u0_u2_n731 ) );
  AOI21_X1 u0_u2_U217 (.ZN( u0_u2_n522 ) , .A( u0_u2_n736 ) , .B1( u0_u2_n757 ) , .B2( u0_u2_n810 ) );
  NOR2_X1 u0_u2_U218 (.ZN( u0_u2_n690 ) , .A2( u0_u2_n706 ) , .A1( u0_u2_n810 ) );
  NOR2_X1 u0_u2_U219 (.A1( u0_u2_n756 ) , .ZN( u0_u2_n774 ) , .A2( u0_u2_n810 ) );
  NOR4_X1 u0_u2_U22 (.ZN( u0_u2_n493 ) , .A1( u0_u2_n514 ) , .A2( u0_u2_n526 ) , .A4( u0_u2_n553 ) , .A3( u0_u2_n618 ) );
  NOR2_X1 u0_u2_U220 (.ZN( u0_u2_n524 ) , .A1( u0_u2_n715 ) , .A2( u0_u2_n810 ) );
  NOR2_X1 u0_u2_U221 (.ZN( u0_u2_n673 ) , .A1( u0_u2_n735 ) , .A2( u0_u2_n810 ) );
  NOR2_X1 u0_u2_U222 (.ZN( u0_u2_n608 ) , .A2( u0_u2_n787 ) , .A1( u0_u2_n810 ) );
  NAND2_X1 u0_u2_U223 (.A2( u0_u2_n468 ) , .A1( u0_u2_n478 ) , .ZN( u0_u2_n704 ) );
  NAND2_X1 u0_u2_U224 (.A1( u0_u2_n459 ) , .A2( u0_u2_n472 ) , .ZN( u0_u2_n676 ) );
  NAND2_X1 u0_u2_U225 (.A2( u0_u2_n455 ) , .A1( u0_u2_n471 ) , .ZN( u0_u2_n822 ) );
  NOR2_X1 u0_u2_U226 (.ZN( u0_u2_n458 ) , .A1( u0_u2_n835 ) , .A2( u0_u2_n836 ) );
  OR3_X1 u0_u2_U227 (.ZN( u0_u2_n453 ) , .A1( u0_u2_n535 ) , .A3( u0_u2_n584 ) , .A2( u0_u2_n882 ) );
  NAND2_X1 u0_u2_U228 (.A1( u0_u2_n458 ) , .A2( u0_u2_n461 ) , .ZN( u0_u2_n821 ) );
  AOI211_X1 u0_u2_U229 (.A( u0_u2_n503 ) , .ZN( u0_u2_n510 ) , .B( u0_u2_n809 ) , .C2( u0_u2_n846 ) , .C1( u0_u2_n858 ) );
  NOR4_X1 u0_u2_U23 (.ZN( u0_u2_n482 ) , .A1( u0_u2_n538 ) , .A3( u0_u2_n575 ) , .A4( u0_u2_n607 ) , .A2( u0_u2_n649 ) );
  NAND4_X1 u0_u2_U230 (.A4( u0_u2_n500 ) , .A3( u0_u2_n501 ) , .A1( u0_u2_n502 ) , .ZN( u0_u2_n809 ) , .A2( u0_u2_n874 ) );
  NOR4_X1 u0_u2_U231 (.A3( u0_u2_n445 ) , .A2( u0_u2_n498 ) , .A1( u0_u2_n499 ) , .ZN( u0_u2_n500 ) , .A4( u0_u2_n619 ) );
  OAI22_X1 u0_u2_U232 (.B1( u0_u2_n497 ) , .ZN( u0_u2_n498 ) , .A1( u0_u2_n693 ) , .A2( u0_u2_n770 ) , .B2( u0_u2_n824 ) );
  NOR2_X1 u0_u2_U233 (.ZN( u0_u2_n444 ) , .A2( u0_u2_n843 ) , .A1( u0_u2_n846 ) );
  NOR2_X1 u0_u2_U234 (.ZN( u0_u2_n632 ) , .A2( u0_u2_n843 ) , .A1( u0_u2_n846 ) );
  NOR2_X1 u0_u2_U235 (.ZN( u0_u2_n445 ) , .A2( u0_u2_n704 ) , .A1( u0_u2_n798 ) );
  OAI222_X1 u0_u2_U236 (.A2( u0_u2_n442 ) , .C1( u0_u2_n443 ) , .ZN( u0_u2_n681 ) , .B1( u0_u2_n754 ) , .B2( u0_u2_n791 ) , .C2( u0_u2_n795 ) , .A1( u0_u2_n824 ) );
  NOR4_X1 u0_u2_U237 (.A4( u0_u2_n491 ) , .ZN( u0_u2_n494 ) , .A1( u0_u2_n573 ) , .A2( u0_u2_n588 ) , .A3( u0_u2_n609 ) );
  AOI222_X1 u0_u2_U238 (.ZN( u0_u2_n613 ) , .A1( u0_u2_n837 ) , .C2( u0_u2_n844 ) , .B1( u0_u2_n849 ) , .A2( u0_u2_n863 ) , .B2( u0_u2_n868 ) , .C1( u0_u2_n875 ) );
  AOI222_X1 u0_u2_U239 (.ZN( u0_u2_n532 ) , .A1( u0_u2_n841 ) , .B2( u0_u2_n844 ) , .C1( u0_u2_n851 ) , .C2( u0_u2_n857 ) , .A2( u0_u2_n859 ) , .B1( u0_u2_n873 ) );
  INV_X1 u0_u2_U24 (.A( u0_u2_n756 ) , .ZN( u0_u2_n870 ) );
  NAND2_X1 u0_u2_U240 (.ZN( u0_u2_n620 ) , .A2( u0_u2_n844 ) , .A1( u0_u2_n880 ) );
  NAND4_X1 u0_u2_U241 (.A4( u0_u2_n486 ) , .A3( u0_u2_n487 ) , .A2( u0_u2_n488 ) , .A1( u0_u2_n489 ) , .ZN( u0_u2_n701 ) );
  NOR2_X1 u0_u2_U242 (.ZN( u0_u2_n586 ) , .A2( u0_u2_n715 ) , .A1( u0_u2_n737 ) );
  OAI21_X1 u0_u2_U243 (.A( u0_u2_n794 ) , .B2( u0_u2_n795 ) , .B1( u0_u2_n796 ) , .ZN( u0_u2_n802 ) );
  AOI21_X1 u0_u2_U244 (.ZN( u0_u2_n646 ) , .B2( u0_u2_n756 ) , .A( u0_u2_n795 ) , .B1( u0_u2_n819 ) );
  AOI21_X1 u0_u2_U245 (.ZN( u0_u2_n449 ) , .A( u0_u2_n706 ) , .B1( u0_u2_n740 ) , .B2( u0_u2_n757 ) );
  NOR2_X1 u0_u2_U246 (.ZN( u0_u2_n525 ) , .A1( u0_u2_n715 ) , .A2( u0_u2_n795 ) );
  INV_X1 u0_u2_U247 (.A( u0_u2_n795 ) , .ZN( u0_u2_n852 ) );
  NOR2_X1 u0_u2_U248 (.ZN( u0_u2_n456 ) , .A1( u0_u2_n855 ) , .A2( w3_4 ) );
  NOR2_X1 u0_u2_U249 (.ZN( u0_u2_n472 ) , .A2( u0_u2_n854 ) , .A1( u0_u2_n855 ) );
  NOR4_X1 u0_u2_U25 (.ZN( u0_u2_n486 ) , .A1( u0_u2_n527 ) , .A4( u0_u2_n564 ) , .A3( u0_u2_n589 ) , .A2( u0_u2_n637 ) );
  OAI222_X1 u0_u2_U250 (.B1( u0_u2_n441 ) , .ZN( u0_u2_n624 ) , .C1( u0_u2_n731 ) , .C2( u0_u2_n754 ) , .B2( u0_u2_n793 ) , .A2( u0_u2_n799 ) , .A1( u0_u2_n823 ) );
  NOR2_X1 u0_u2_U251 (.ZN( u0_u2_n467 ) , .A1( u0_u2_n856 ) , .A2( w3_7 ) );
  AOI21_X1 u0_u2_U252 (.ZN( u0_u2_n647 ) , .B2( u0_u2_n754 ) , .A( u0_u2_n799 ) , .B1( u0_u2_n810 ) );
  AOI21_X1 u0_u2_U253 (.A( u0_u2_n740 ) , .ZN( u0_u2_n741 ) , .B2( u0_u2_n787 ) , .B1( u0_u2_n799 ) );
  AOI21_X1 u0_u2_U254 (.ZN( u0_u2_n521 ) , .A( u0_u2_n786 ) , .B2( u0_u2_n799 ) , .B1( u0_u2_n819 ) );
  AOI21_X1 u0_u2_U255 (.B2( u0_u2_n770 ) , .ZN( u0_u2_n771 ) , .A( u0_u2_n795 ) , .B1( u0_u2_n799 ) );
  INV_X1 u0_u2_U256 (.A( u0_u2_n799 ) , .ZN( u0_u2_n858 ) );
  NOR2_X1 u0_u2_U257 (.ZN( u0_u2_n564 ) , .A1( u0_u2_n799 ) , .A2( u0_u2_n821 ) );
  NOR2_X1 u0_u2_U258 (.ZN( u0_u2_n590 ) , .A1( u0_u2_n799 ) , .A2( u0_u2_n824 ) );
  AOI221_X1 u0_u2_U259 (.A( u0_u2_n496 ) , .ZN( u0_u2_n501 ) , .B2( u0_u2_n843 ) , .C2( u0_u2_n848 ) , .C1( u0_u2_n858 ) , .B1( u0_u2_n867 ) );
  NOR3_X1 u0_u2_U26 (.ZN( u0_u2_n487 ) , .A2( u0_u2_n515 ) , .A3( u0_u2_n608 ) , .A1( u0_u2_n617 ) );
  NOR3_X1 u0_u2_U260 (.ZN( u0_u2_n447 ) , .A2( u0_u2_n843 ) , .A3( u0_u2_n844 ) , .A1( u0_u2_n853 ) );
  NOR4_X1 u0_u2_U261 (.A3( u0_u2_n680 ) , .A1( u0_u2_n681 ) , .ZN( u0_u2_n682 ) , .A4( u0_u2_n722 ) , .A2( u0_u2_n866 ) );
  INV_X1 u0_u2_U262 (.A( u0_u2_n679 ) , .ZN( u0_u2_n866 ) );
  NOR2_X1 u0_u2_U263 (.ZN( u0_u2_n478 ) , .A1( u0_u2_n833 ) , .A2( w3_1 ) );
  INV_X1 u0_u2_U264 (.ZN( u0_u2_n834 ) , .A( w3_1 ) );
  CLKBUF_X1 u0_u2_U265 (.Z( u0_u2_n446 ) , .A( u0_u2_n798 ) );
  NOR2_X1 u0_u2_U266 (.A2( u0_u2_n438 ) , .A1( u0_u2_n583 ) , .ZN( u0_u2_n594 ) );
  OAI22_X1 u0_u2_U267 (.B2( u0_u2_n786 ) , .B1( u0_u2_n787 ) , .ZN( u0_u2_n788 ) , .A2( u0_u2_n821 ) , .A1( u0_u2_n822 ) );
  AOI21_X1 u0_u2_U268 (.B1( u0_u2_n443 ) , .ZN( u0_u2_n596 ) , .B2( u0_u2_n706 ) , .A( u0_u2_n824 ) );
  INV_X1 u0_u2_U269 (.A( u0_u2_n822 ) , .ZN( u0_u2_n862 ) );
  AOI211_X1 u0_u2_U27 (.B( u0_u2_n484 ) , .A( u0_u2_n485 ) , .ZN( u0_u2_n489 ) , .C2( u0_u2_n840 ) , .C1( u0_u2_n868 ) );
  NOR2_X1 u0_u2_U270 (.ZN( u0_u2_n674 ) , .A1( u0_u2_n757 ) , .A2( u0_u2_n822 ) );
  NOR2_X1 u0_u2_U271 (.A1( u0_u2_n443 ) , .ZN( u0_u2_n477 ) , .A2( u0_u2_n786 ) );
  AOI21_X1 u0_u2_U272 (.B1( u0_u2_n443 ) , .ZN( u0_u2_n546 ) , .B2( u0_u2_n819 ) , .A( u0_u2_n821 ) );
  AOI21_X1 u0_u2_U273 (.B1( u0_u2_n443 ) , .ZN( u0_u2_n457 ) , .B2( u0_u2_n799 ) , .A( u0_u2_n810 ) );
  NOR2_X1 u0_u2_U274 (.A2( u0_u2_n443 ) , .ZN( u0_u2_n637 ) , .A1( u0_u2_n754 ) );
  INV_X1 u0_u2_U275 (.ZN( u0_u2_n865 ) , .A( w3_7 ) );
  AOI222_X1 u0_u2_U276 (.C2( u0_u2_n816 ) , .B2( u0_u2_n817 ) , .A2( u0_u2_n818 ) , .ZN( u0_u2_n830 ) , .C1( u0_u2_n839 ) , .A1( u0_u2_n846 ) , .B1( u0_u2_n860 ) );
  AOI22_X1 u0_u2_U277 (.ZN( u0_u2_n734 ) , .B1( u0_u2_n839 ) , .A2( u0_u2_n845 ) , .A1( u0_u2_n870 ) , .B2( u0_u2_n873 ) );
  AOI222_X1 u0_u2_U278 (.ZN( u0_u2_n476 ) , .B1( u0_u2_n839 ) , .A1( u0_u2_n846 ) , .C1( u0_u2_n849 ) , .C2( u0_u2_n858 ) , .A2( u0_u2_n862 ) , .B2( u0_u2_n872 ) );
  NOR2_X1 u0_u2_U279 (.A2( u0_u2_n443 ) , .ZN( u0_u2_n662 ) , .A1( u0_u2_n797 ) );
  NOR4_X1 u0_u2_U28 (.ZN( u0_u2_n488 ) , .A3( u0_u2_n539 ) , .A4( u0_u2_n552 ) , .A2( u0_u2_n574 ) , .A1( u0_u2_n724 ) );
  NOR2_X1 u0_u2_U280 (.ZN( u0_u2_n693 ) , .A1( u0_u2_n838 ) , .A2( u0_u2_n839 ) );
  NOR2_X1 u0_u2_U281 (.ZN( u0_u2_n528 ) , .A1( u0_u2_n797 ) , .A2( u0_u2_n819 ) );
  NOR2_X1 u0_u2_U282 (.ZN( u0_u2_n740 ) , .A2( u0_u2_n839 ) , .A1( u0_u2_n852 ) );
  NOR2_X1 u0_u2_U283 (.ZN( u0_u2_n668 ) , .A1( u0_u2_n736 ) , .A2( u0_u2_n797 ) );
  NOR2_X1 u0_u2_U284 (.ZN( u0_u2_n675 ) , .A2( u0_u2_n715 ) , .A1( u0_u2_n797 ) );
  INV_X1 u0_u2_U285 (.A( u0_u2_n797 ) , .ZN( u0_u2_n839 ) );
  NOR2_X1 u0_u2_U286 (.ZN( u0_u2_n468 ) , .A1( u0_u2_n836 ) , .A2( w3_2 ) );
  INV_X1 u0_u2_U287 (.ZN( u0_u2_n835 ) , .A( w3_2 ) );
  AOI21_X1 u0_u2_U288 (.ZN( u0_u2_n600 ) , .B1( u0_u2_n757 ) , .A( u0_u2_n799 ) , .B2( u0_u2_n820 ) );
  AOI21_X1 u0_u2_U289 (.A( u0_u2_n819 ) , .B2( u0_u2_n820 ) , .B1( u0_u2_n821 ) , .ZN( u0_u2_n826 ) );
  NOR2_X1 u0_u2_U29 (.ZN( u0_u2_n687 ) , .A2( u0_u2_n841 ) , .A1( u0_u2_n846 ) );
  AOI21_X1 u0_u2_U290 (.ZN( u0_u2_n656 ) , .B1( u0_u2_n736 ) , .B2( u0_u2_n770 ) , .A( u0_u2_n820 ) );
  NOR2_X1 u0_u2_U291 (.A2( u0_u2_n820 ) , .A1( u0_u2_n822 ) , .ZN( u0_u2_n828 ) );
  NOR2_X1 u0_u2_U292 (.ZN( u0_u2_n585 ) , .A1( u0_u2_n715 ) , .A2( u0_u2_n820 ) );
  NOR2_X1 u0_u2_U293 (.ZN( u0_u2_n672 ) , .A1( u0_u2_n787 ) , .A2( u0_u2_n820 ) );
  NOR2_X1 u0_u2_U294 (.A1( u0_u2_n706 ) , .ZN( u0_u2_n775 ) , .A2( u0_u2_n820 ) );
  NOR2_X1 u0_u2_U295 (.ZN( u0_u2_n661 ) , .A1( u0_u2_n735 ) , .A2( u0_u2_n820 ) );
  INV_X1 u0_u2_U296 (.A( u0_u2_n820 ) , .ZN( u0_u2_n843 ) );
  AOI21_X1 u0_u2_U297 (.ZN( u0_u2_n598 ) , .B2( u0_u2_n770 ) , .A( u0_u2_n792 ) , .B1( u0_u2_n819 ) );
  AND2_X1 u0_u2_U298 (.ZN( u0_u2_n739 ) , .A1( u0_u2_n786 ) , .A2( u0_u2_n792 ) );
  NOR2_X1 u0_u2_U299 (.ZN( u0_u2_n670 ) , .A1( u0_u2_n736 ) , .A2( u0_u2_n792 ) );
  NAND2_X1 u0_u2_U3 (.ZN( u0_u2_n438 ) , .A1( u0_u2_n439 ) , .A2( u0_u2_n440 ) );
  NAND4_X1 u0_u2_U30 (.A4( u0_u2_n610 ) , .A3( u0_u2_n611 ) , .A2( u0_u2_n612 ) , .A1( u0_u2_n613 ) , .ZN( u0_u2_n729 ) );
  NOR2_X1 u0_u2_U300 (.ZN( u0_u2_n515 ) , .A2( u0_u2_n787 ) , .A1( u0_u2_n792 ) );
  NOR2_X1 u0_u2_U301 (.A2( u0_u2_n443 ) , .ZN( u0_u2_n622 ) , .A1( u0_u2_n792 ) );
  INV_X1 u0_u2_U302 (.A( u0_u2_n792 ) , .ZN( u0_u2_n853 ) );
  OAI22_X1 u0_u2_U303 (.ZN( u0_u2_n490 ) , .A1( u0_u2_n715 ) , .B2( u0_u2_n792 ) , .A2( u0_u2_n813 ) , .B1( u0_u2_n819 ) );
  NOR2_X1 u0_u2_U304 (.ZN( u0_u2_n636 ) , .A2( u0_u2_n735 ) , .A1( u0_u2_n792 ) );
  NOR2_X1 u0_u2_U305 (.ZN( u0_u2_n550 ) , .A2( u0_u2_n715 ) , .A1( u0_u2_n792 ) );
  NOR2_X1 u0_u2_U306 (.ZN( u0_u2_n551 ) , .A2( u0_u2_n792 ) , .A1( u0_u2_n799 ) );
  NAND4_X1 u0_u2_U307 (.A4( u0_u2_n698 ) , .A3( u0_u2_n699 ) , .A1( u0_u2_n700 ) , .ZN( u0_u2_n783 ) , .A2( u0_u2_n879 ) );
  NOR4_X1 u0_u2_U308 (.A4( u0_u2_n783 ) , .A3( u0_u2_n784 ) , .A1( u0_u2_n785 ) , .ZN( u0_u2_n806 ) , .A2( u0_u2_n808 ) );
  AOI211_X1 u0_u2_U309 (.A( u0_u2_n644 ) , .ZN( u0_u2_n652 ) , .B( u0_u2_n750 ) , .C2( u0_u2_n846 ) , .C1( u0_u2_n861 ) );
  NOR3_X1 u0_u2_U31 (.A1( u0_u2_n606 ) , .ZN( u0_u2_n611 ) , .A3( u0_u2_n670 ) , .A2( u0_u2_n777 ) );
  NOR3_X1 u0_u2_U310 (.A3( u0_u2_n748 ) , .A2( u0_u2_n749 ) , .A1( u0_u2_n750 ) , .ZN( u0_u2_n767 ) );
  NAND4_X1 u0_u2_U311 (.A4( u0_u2_n640 ) , .A3( u0_u2_n641 ) , .A2( u0_u2_n642 ) , .A1( u0_u2_n643 ) , .ZN( u0_u2_n750 ) );
  NOR3_X1 u0_u2_U312 (.A3( u0_u2_n628 ) , .A2( u0_u2_n629 ) , .ZN( u0_u2_n643 ) , .A1( u0_u2_n732 ) );
  NOR4_X1 u0_u2_U313 (.A4( u0_u2_n621 ) , .A3( u0_u2_n622 ) , .A2( u0_u2_n623 ) , .A1( u0_u2_n624 ) , .ZN( u0_u2_n625 ) );
  NOR2_X1 u0_u2_U314 (.ZN( u0_u2_n459 ) , .A1( u0_u2_n865 ) , .A2( w3_6 ) );
  NOR2_X1 u0_u2_U315 (.ZN( u0_u2_n454 ) , .A2( u0_u2_n856 ) , .A1( u0_u2_n865 ) );
  NOR2_X1 u0_u2_U316 (.ZN( u0_u2_n471 ) , .A2( w3_6 ) , .A1( w3_7 ) );
  INV_X1 u0_u2_U317 (.ZN( u0_u2_n856 ) , .A( w3_6 ) );
  AOI21_X1 u0_u2_U318 (.ZN( u0_u2_n505 ) , .A( u0_u2_n731 ) , .B2( u0_u2_n769 ) , .B1( u0_u2_n821 ) );
  OAI22_X1 u0_u2_U319 (.ZN( u0_u2_n496 ) , .A1( u0_u2_n731 ) , .B2( u0_u2_n735 ) , .B1( u0_u2_n737 ) , .A2( u0_u2_n786 ) );
  NOR4_X1 u0_u2_U32 (.A3( u0_u2_n607 ) , .A2( u0_u2_n608 ) , .A1( u0_u2_n609 ) , .ZN( u0_u2_n610 ) , .A4( u0_u2_n662 ) );
  NOR2_X1 u0_u2_U320 (.ZN( u0_u2_n719 ) , .A2( u0_u2_n731 ) , .A1( u0_u2_n797 ) );
  NOR2_X1 u0_u2_U321 (.ZN( u0_u2_n535 ) , .A2( u0_u2_n731 ) , .A1( u0_u2_n810 ) );
  NOR2_X1 u0_u2_U322 (.ZN( u0_u2_n616 ) , .A2( u0_u2_n731 ) , .A1( u0_u2_n824 ) );
  NOR2_X1 u0_u2_U323 (.ZN( u0_u2_n533 ) , .A1( u0_u2_n731 ) , .A2( u0_u2_n757 ) );
  NOR2_X1 u0_u2_U324 (.ZN( u0_u2_n541 ) , .A1( u0_u2_n731 ) , .A2( u0_u2_n795 ) );
  NOR2_X1 u0_u2_U325 (.ZN( u0_u2_n638 ) , .A1( u0_u2_n731 ) , .A2( u0_u2_n820 ) );
  NOR2_X1 u0_u2_U326 (.ZN( u0_u2_n540 ) , .A2( u0_u2_n731 ) , .A1( u0_u2_n737 ) );
  INV_X1 u0_u2_U327 (.A( u0_u2_n731 ) , .ZN( u0_u2_n863 ) );
  NOR2_X1 u0_u2_U328 (.ZN( u0_u2_n455 ) , .A1( u0_u2_n854 ) , .A2( w3_5 ) );
  NOR2_X1 u0_u2_U329 (.ZN( u0_u2_n448 ) , .A2( w3_4 ) , .A1( w3_5 ) );
  NOR4_X1 u0_u2_U33 (.A4( u0_u2_n694 ) , .A3( u0_u2_n695 ) , .A2( u0_u2_n696 ) , .A1( u0_u2_n697 ) , .ZN( u0_u2_n698 ) );
  INV_X1 u0_u2_U330 (.ZN( u0_u2_n855 ) , .A( w3_5 ) );
  AOI21_X1 u0_u2_U331 (.A( u0_u2_n446 ) , .ZN( u0_u2_n648 ) , .B1( u0_u2_n687 ) , .B2( u0_u2_n824 ) );
  AOI21_X1 u0_u2_U332 (.B2( u0_u2_n446 ) , .A( u0_u2_n797 ) , .B1( u0_u2_n799 ) , .ZN( u0_u2_n800 ) );
  OAI22_X1 u0_u2_U333 (.B1( u0_u2_n446 ) , .ZN( u0_u2_n702 ) , .A2( u0_u2_n737 ) , .A1( u0_u2_n787 ) , .B2( u0_u2_n824 ) );
  AOI21_X1 u0_u2_U334 (.B2( u0_u2_n446 ) , .ZN( u0_u2_n504 ) , .A( u0_u2_n786 ) , .B1( u0_u2_n811 ) );
  AOI21_X1 u0_u2_U335 (.B2( u0_u2_n446 ) , .ZN( u0_u2_n571 ) , .B1( u0_u2_n731 ) , .A( u0_u2_n786 ) );
  AOI21_X1 u0_u2_U336 (.ZN( u0_u2_n450 ) , .B1( u0_u2_n796 ) , .B2( u0_u2_n798 ) , .A( u0_u2_n821 ) );
  NOR2_X1 u0_u2_U337 (.ZN( u0_u2_n671 ) , .A1( u0_u2_n792 ) , .A2( u0_u2_n798 ) );
  NOR2_X1 u0_u2_U338 (.ZN( u0_u2_n562 ) , .A1( u0_u2_n757 ) , .A2( u0_u2_n798 ) );
  NOR2_X1 u0_u2_U339 (.ZN( u0_u2_n566 ) , .A2( u0_u2_n798 ) , .A1( u0_u2_n810 ) );
  AOI221_X1 u0_u2_U34 (.A( u0_u2_n688 ) , .ZN( u0_u2_n699 ) , .B2( u0_u2_n847 ) , .C1( u0_u2_n849 ) , .C2( u0_u2_n869 ) , .B1( u0_u2_n872 ) );
  NAND2_X2 u0_u2_U340 (.A1( u0_u2_n462 ) , .A2( u0_u2_n469 ) , .ZN( u0_u2_n757 ) );
  NOR2_X1 u0_u2_U341 (.ZN( u0_u2_n649 ) , .A2( u0_u2_n795 ) , .A1( u0_u2_n798 ) );
  NOR2_X1 u0_u2_U342 (.ZN( u0_u2_n691 ) , .A1( u0_u2_n798 ) , .A2( u0_u2_n820 ) );
  NOR2_X1 u0_u2_U343 (.ZN( u0_u2_n549 ) , .A1( u0_u2_n769 ) , .A2( u0_u2_n798 ) );
  INV_X1 u0_u2_U344 (.A( u0_u2_n798 ) , .ZN( u0_u2_n880 ) );
  AOI21_X1 u0_u2_U345 (.B2( u0_u2_n442 ) , .ZN( u0_u2_n517 ) , .A( u0_u2_n737 ) , .B1( u0_u2_n822 ) );
  AOI21_X1 u0_u2_U346 (.B1( u0_u2_n446 ) , .ZN( u0_u2_n633 ) , .B2( u0_u2_n676 ) , .A( u0_u2_n797 ) );
  INV_X1 u0_u2_U347 (.A( u0_u2_n676 ) , .ZN( u0_u2_n872 ) );
  NOR2_X1 u0_u2_U348 (.A1( u0_u2_n442 ) , .ZN( u0_u2_n773 ) , .A2( u0_u2_n820 ) );
  NOR2_X1 u0_u2_U349 (.A1( u0_u2_n442 ) , .ZN( u0_u2_n659 ) , .A2( u0_u2_n821 ) );
  NOR2_X1 u0_u2_U35 (.A1( u0_u2_n685 ) , .ZN( u0_u2_n700 ) , .A2( u0_u2_n814 ) );
  AOI21_X1 u0_u2_U350 (.A( u0_u2_n442 ) , .ZN( u0_u2_n484 ) , .B1( u0_u2_n757 ) , .B2( u0_u2_n813 ) );
  NOR2_X1 u0_u2_U351 (.A1( u0_u2_n442 ) , .ZN( u0_u2_n534 ) , .A2( u0_u2_n786 ) );
  NOR2_X1 u0_u2_U352 (.A1( u0_u2_n442 ) , .ZN( u0_u2_n609 ) , .A2( u0_u2_n810 ) );
  NOR2_X1 u0_u2_U353 (.A2( u0_u2_n442 ) , .ZN( u0_u2_n635 ) , .A1( u0_u2_n792 ) );
  NOR2_X1 u0_u2_U354 (.ZN( u0_u2_n588 ) , .A1( u0_u2_n676 ) , .A2( u0_u2_n795 ) );
  OAI22_X1 u0_u2_U355 (.ZN( u0_u2_n644 ) , .A1( u0_u2_n706 ) , .B2( u0_u2_n735 ) , .A2( u0_u2_n769 ) , .B1( u0_u2_n823 ) );
  AOI21_X1 u0_u2_U356 (.ZN( u0_u2_n506 ) , .B1( u0_u2_n687 ) , .A( u0_u2_n819 ) , .B2( u0_u2_n823 ) );
  OAI22_X1 u0_u2_U357 (.A1( u0_u2_n731 ) , .ZN( u0_u2_n733 ) , .B2( u0_u2_n757 ) , .B1( u0_u2_n819 ) , .A2( u0_u2_n823 ) );
  AOI21_X1 u0_u2_U358 (.A( u0_u2_n443 ) , .B2( u0_u2_n823 ) , .B1( u0_u2_n824 ) , .ZN( u0_u2_n825 ) );
  OAI22_X1 u0_u2_U359 (.B1( u0_u2_n442 ) , .A1( u0_u2_n443 ) , .ZN( u0_u2_n631 ) , .B2( u0_u2_n754 ) , .A2( u0_u2_n823 ) );
  NOR2_X1 u0_u2_U36 (.ZN( u0_u2_n552 ) , .A1( u0_u2_n756 ) , .A2( u0_u2_n821 ) );
  NOR2_X1 u0_u2_U360 (.ZN( u0_u2_n606 ) , .A2( u0_u2_n798 ) , .A1( u0_u2_n823 ) );
  NOR2_X1 u0_u2_U361 (.ZN( u0_u2_n538 ) , .A2( u0_u2_n787 ) , .A1( u0_u2_n823 ) );
  NOR2_X1 u0_u2_U362 (.ZN( u0_u2_n526 ) , .A2( u0_u2_n706 ) , .A1( u0_u2_n823 ) );
  NOR2_X1 u0_u2_U363 (.A1( u0_u2_n442 ) , .ZN( u0_u2_n695 ) , .A2( u0_u2_n823 ) );
  NOR2_X1 u0_u2_U364 (.ZN( u0_u2_n565 ) , .A1( u0_u2_n715 ) , .A2( u0_u2_n823 ) );
  NOR2_X1 u0_u2_U365 (.ZN( u0_u2_n692 ) , .A1( u0_u2_n736 ) , .A2( u0_u2_n823 ) );
  NAND2_X1 u0_u2_U366 (.ZN( u0_u2_n678 ) , .A1( u0_u2_n813 ) , .A2( u0_u2_n823 ) );
  NOR2_X1 u0_u2_U367 (.ZN( u0_u2_n469 ) , .A2( w3_0 ) , .A1( w3_1 ) );
  NOR2_X1 u0_u2_U368 (.ZN( u0_u2_n461 ) , .A1( u0_u2_n834 ) , .A2( w3_0 ) );
  INV_X1 u0_u2_U369 (.ZN( u0_u2_n833 ) , .A( w3_0 ) );
  NOR2_X1 u0_u2_U37 (.ZN( u0_u2_n502 ) , .A1( u0_u2_n685 ) , .A2( u0_u2_n701 ) );
  INV_X1 u0_u2_U370 (.A( u0_u2_n819 ) , .ZN( u0_u2_n861 ) );
  INV_X1 u0_u2_U371 (.A( u0_u2_n823 ) , .ZN( u0_u2_n838 ) );
  INV_X1 u0_u2_U372 (.A( u0_u2_n810 ) , .ZN( u0_u2_n850 ) );
  INV_X1 u0_u2_U373 (.ZN( u0_u2_n854 ) , .A( w3_4 ) );
  INV_X1 u0_u2_U374 (.A( u0_u2_n441 ) , .ZN( u0_u2_n845 ) );
  NOR2_X1 u0_u2_U375 (.A1( u0_u2_n704 ) , .ZN( u0_u2_n777 ) , .A2( u0_u2_n822 ) );
  AOI21_X1 u0_u2_U376 (.B2( u0_u2_n441 ) , .ZN( u0_u2_n578 ) , .B1( u0_u2_n813 ) , .A( u0_u2_n819 ) );
  NOR2_X1 u0_u2_U377 (.ZN( u0_u2_n639 ) , .A2( u0_u2_n704 ) , .A1( u0_u2_n731 ) );
  NOR2_X1 u0_u2_U378 (.A2( u0_u2_n441 ) , .A1( u0_u2_n787 ) , .ZN( u0_u2_n827 ) );
  AOI21_X1 u0_u2_U379 (.B2( u0_u2_n441 ) , .ZN( u0_u2_n485 ) , .A( u0_u2_n756 ) , .B1( u0_u2_n786 ) );
  INV_X1 u0_u2_U38 (.A( u0_u2_n821 ) , .ZN( u0_u2_n840 ) );
  NOR2_X1 u0_u2_U380 (.A2( u0_u2_n441 ) , .ZN( u0_u2_n573 ) , .A1( u0_u2_n770 ) );
  NOR2_X1 u0_u2_U381 (.ZN( u0_u2_n669 ) , .A2( u0_u2_n704 ) , .A1( u0_u2_n736 ) );
  NOR2_X1 u0_u2_U382 (.A2( u0_u2_n441 ) , .ZN( u0_u2_n723 ) , .A1( u0_u2_n799 ) );
  NOR2_X1 u0_u2_U383 (.A2( u0_u2_n441 ) , .ZN( u0_u2_n601 ) , .A1( u0_u2_n735 ) );
  NOR2_X1 u0_u2_U384 (.A2( u0_u2_n441 ) , .ZN( u0_u2_n548 ) , .A1( u0_u2_n706 ) );
  NOR2_X1 u0_u2_U385 (.ZN( u0_u2_n587 ) , .A2( u0_u2_n704 ) , .A1( u0_u2_n798 ) );
  NOR2_X1 u0_u2_U386 (.ZN( u0_u2_n479 ) , .A2( w3_2 ) , .A1( w3_3 ) );
  NOR2_X1 u0_u2_U387 (.ZN( u0_u2_n462 ) , .A1( u0_u2_n835 ) , .A2( w3_3 ) );
  INV_X1 u0_u2_U388 (.ZN( u0_u2_n836 ) , .A( w3_3 ) );
  AOI21_X1 u0_u2_U389 (.ZN( u0_u2_n583 ) , .B2( u0_u2_n731 ) , .B1( u0_u2_n755 ) , .A( u0_u2_n792 ) );
  NAND4_X1 u0_u2_U39 (.A4( u0_u2_n664 ) , .A3( u0_u2_n665 ) , .A2( u0_u2_n666 ) , .A1( u0_u2_n667 ) , .ZN( u0_u2_n807 ) );
  OAI222_X1 u0_u2_U390 (.B2( u0_u2_n754 ) , .B1( u0_u2_n755 ) , .A2( u0_u2_n756 ) , .ZN( u0_u2_n764 ) , .C2( u0_u2_n812 ) , .C1( u0_u2_n821 ) , .A1( u0_u2_n824 ) );
  OAI21_X1 u0_u2_U391 (.A( u0_u2_n738 ) , .B1( u0_u2_n739 ) , .ZN( u0_u2_n743 ) , .B2( u0_u2_n812 ) );
  OAI22_X1 u0_u2_U392 (.B2( u0_u2_n810 ) , .B1( u0_u2_n811 ) , .A2( u0_u2_n812 ) , .A1( u0_u2_n813 ) , .ZN( u0_u2_n815 ) );
  OAI222_X1 u0_u2_U393 (.C2( u0_u2_n444 ) , .ZN( u0_u2_n512 ) , .B2( u0_u2_n654 ) , .B1( u0_u2_n754 ) , .A2( u0_u2_n755 ) , .C1( u0_u2_n812 ) , .A1( u0_u2_n813 ) );
  AOI21_X1 u0_u2_U394 (.ZN( u0_u2_n657 ) , .A( u0_u2_n786 ) , .B1( u0_u2_n799 ) , .B2( u0_u2_n812 ) );
  INV_X1 u0_u2_U395 (.A( u0_u2_n812 ) , .ZN( u0_u2_n867 ) );
  NOR2_X1 u0_u2_U396 (.ZN( u0_u2_n742 ) , .A2( u0_u2_n810 ) , .A1( u0_u2_n812 ) );
  NOR2_X1 u0_u2_U397 (.ZN( u0_u2_n491 ) , .A1( u0_u2_n795 ) , .A2( u0_u2_n812 ) );
  NOR2_X1 u0_u2_U398 (.ZN( u0_u2_n574 ) , .A1( u0_u2_n754 ) , .A2( u0_u2_n812 ) );
  AOI21_X1 u0_u2_U399 (.A( u0_u2_n441 ) , .B1( u0_u2_n442 ) , .ZN( u0_u2_n559 ) , .B2( u0_u2_n812 ) );
  NOR3_X1 u0_u2_U4 (.A3( u0_u2_n807 ) , .A2( u0_u2_n808 ) , .A1( u0_u2_n809 ) , .ZN( u0_u2_n832 ) );
  NOR3_X1 u0_u2_U40 (.A3( u0_u2_n661 ) , .A2( u0_u2_n662 ) , .A1( u0_u2_n663 ) , .ZN( u0_u2_n664 ) );
  NAND2_X1 u0_u2_U400 (.ZN( u0_u2_n760 ) , .A1( u0_u2_n770 ) , .A2( u0_u2_n812 ) );
  NOR2_X1 u0_u2_U401 (.ZN( u0_u2_n722 ) , .A1( u0_u2_n812 ) , .A2( u0_u2_n824 ) );
  NOR2_X1 u0_u2_U402 (.ZN( u0_u2_n563 ) , .A1( u0_u2_n769 ) , .A2( u0_u2_n812 ) );
  NOR2_X1 u0_u2_U403 (.ZN( u0_u2_n677 ) , .A1( u0_u2_n797 ) , .A2( u0_u2_n812 ) );
  NAND4_X1 u0_u2_U404 (.ZN( u0_subword_11 ) , .A4( u0_u2_n711 ) , .A3( u0_u2_n712 ) , .A2( u0_u2_n713 ) , .A1( u0_u2_n714 ) );
  INV_X1 u0_u2_U405 (.A( u0_u2_n713 ) , .ZN( u0_u2_n883 ) );
  OAI22_X1 u0_u2_U406 (.B2( u0_u2_n751 ) , .ZN( u0_u2_n753 ) , .A2( u0_u2_n769 ) , .B1( u0_u2_n787 ) , .A1( u0_u2_n799 ) );
  OAI22_X1 u0_u2_U407 (.B1( u0_u2_n446 ) , .ZN( u0_u2_n503 ) , .A2( u0_u2_n751 ) , .A1( u0_u2_n787 ) , .B2( u0_u2_n813 ) );
  NOR2_X1 u0_u2_U408 (.ZN( u0_u2_n523 ) , .A1( u0_u2_n715 ) , .A2( u0_u2_n751 ) );
  OAI22_X1 u0_u2_U409 (.ZN( u0_u2_n717 ) , .A2( u0_u2_n735 ) , .B2( u0_u2_n736 ) , .A1( u0_u2_n751 ) , .B1( u0_u2_n820 ) );
  NOR3_X1 u0_u2_U41 (.A3( u0_u2_n655 ) , .A2( u0_u2_n656 ) , .A1( u0_u2_n657 ) , .ZN( u0_u2_n666 ) );
  NOR2_X1 u0_u2_U410 (.A2( u0_u2_n751 ) , .ZN( u0_u2_n776 ) , .A1( u0_u2_n819 ) );
  OAI22_X1 u0_u2_U411 (.B1( u0_u2_n447 ) , .ZN( u0_u2_n451 ) , .A2( u0_u2_n735 ) , .A1( u0_u2_n751 ) , .B2( u0_u2_n756 ) );
  NOR2_X1 u0_u2_U412 (.ZN( u0_u2_n554 ) , .A1( u0_u2_n706 ) , .A2( u0_u2_n751 ) );
  NOR2_X1 u0_u2_U413 (.ZN( u0_u2_n537 ) , .A2( u0_u2_n751 ) , .A1( u0_u2_n799 ) );
  NOR2_X1 u0_u2_U414 (.A2( u0_u2_n751 ) , .ZN( u0_u2_n762 ) , .A1( u0_u2_n812 ) );
  NOR2_X1 u0_u2_U415 (.A1( u0_u2_n442 ) , .ZN( u0_u2_n680 ) , .A2( u0_u2_n751 ) );
  NOR2_X1 u0_u2_U416 (.ZN( u0_u2_n725 ) , .A2( u0_u2_n731 ) , .A1( u0_u2_n751 ) );
  NOR2_X1 u0_u2_U417 (.ZN( u0_u2_n589 ) , .A1( u0_u2_n751 ) , .A2( u0_u2_n822 ) );
  INV_X1 u0_u2_U418 (.A( u0_u2_n751 ) , .ZN( u0_u2_n844 ) );
  NAND4_X1 u0_u2_U419 (.ZN( u0_subword_10 ) , .A4( u0_u2_n650 ) , .A3( u0_u2_n651 ) , .A2( u0_u2_n652 ) , .A1( u0_u2_n653 ) );
  NOR3_X1 u0_u2_U42 (.A3( u0_u2_n658 ) , .A2( u0_u2_n659 ) , .A1( u0_u2_n660 ) , .ZN( u0_u2_n665 ) );
  OAI22_X1 u0_u2_U420 (.ZN( u0_u2_n595 ) , .A2( u0_u2_n754 ) , .B2( u0_u2_n769 ) , .A1( u0_u2_n770 ) , .B1( u0_u2_n791 ) );
  NAND2_X1 u0_u2_U421 (.A1( u0_u2_n736 ) , .A2( u0_u2_n791 ) , .ZN( u0_u2_n818 ) );
  AOI21_X1 u0_u2_U422 (.ZN( u0_u2_n599 ) , .B1( u0_u2_n735 ) , .B2( u0_u2_n791 ) , .A( u0_u2_n797 ) );
  AOI21_X1 u0_u2_U423 (.ZN( u0_u2_n655 ) , .A( u0_u2_n769 ) , .B2( u0_u2_n791 ) , .B1( u0_u2_n799 ) );
  AOI21_X1 u0_u2_U424 (.ZN( u0_u2_n630 ) , .B1( u0_u2_n706 ) , .A( u0_u2_n786 ) , .B2( u0_u2_n791 ) );
  OAI22_X1 u0_u2_U425 (.ZN( u0_u2_n688 ) , .A1( u0_u2_n706 ) , .A2( u0_u2_n737 ) , .B2( u0_u2_n791 ) , .B1( u0_u2_n824 ) );
  OAI21_X1 u0_u2_U426 (.A( u0_u2_n620 ) , .ZN( u0_u2_n623 ) , .B1( u0_u2_n632 ) , .B2( u0_u2_n791 ) );
  NOR2_X1 u0_u2_U427 (.ZN( u0_u2_n658 ) , .A1( u0_u2_n791 ) , .A2( u0_u2_n795 ) );
  NOR2_X1 u0_u2_U428 (.ZN( u0_u2_n617 ) , .A1( u0_u2_n791 ) , .A2( u0_u2_n823 ) );
  NOR2_X1 u0_u2_U429 (.ZN( u0_u2_n560 ) , .A2( u0_u2_n751 ) , .A1( u0_u2_n791 ) );
  NAND4_X1 u0_u2_U43 (.A4( u0_u2_n567 ) , .A3( u0_u2_n568 ) , .A2( u0_u2_n569 ) , .A1( u0_u2_n570 ) , .ZN( u0_u2_n614 ) );
  NOR2_X1 u0_u2_U430 (.A2( u0_u2_n441 ) , .ZN( u0_u2_n607 ) , .A1( u0_u2_n791 ) );
  INV_X1 u0_u2_U431 (.A( u0_u2_n791 ) , .ZN( u0_u2_n868 ) );
  AOI21_X1 u0_u2_U432 (.ZN( u0_u2_n507 ) , .A( u0_u2_n704 ) , .B1( u0_u2_n715 ) , .B2( u0_u2_n793 ) );
  OAI22_X1 u0_u2_U433 (.ZN( u0_u2_n597 ) , .B1( u0_u2_n737 ) , .B2( u0_u2_n756 ) , .A2( u0_u2_n793 ) , .A1( u0_u2_n810 ) );
  AOI222_X1 u0_u2_U434 (.ZN( u0_u2_n520 ) , .C1( u0_u2_n839 ) , .B2( u0_u2_n844 ) , .A2( u0_u2_n850 ) , .C2( u0_u2_n869 ) , .B1( u0_u2_n870 ) , .A1( u0_u2_n873 ) );
  AOI222_X1 u0_u2_U435 (.ZN( u0_u2_n612 ) , .B2( u0_u2_n678 ) , .B1( u0_u2_n760 ) , .C2( u0_u2_n838 ) , .A1( u0_u2_n840 ) , .A2( u0_u2_n869 ) , .C1( u0_u2_n870 ) );
  AOI221_X1 u0_u2_U436 (.A( u0_u2_n490 ) , .ZN( u0_u2_n495 ) , .B1( u0_u2_n838 ) , .C2( u0_u2_n851 ) , .C1( u0_u2_n859 ) , .B2( u0_u2_n869 ) );
  NAND3_X1 u0_u2_U437 (.ZN( u0_subword_14 ) , .A3( u0_u2_n804 ) , .A2( u0_u2_n805 ) , .A1( u0_u2_n806 ) );
  NAND3_X1 u0_u2_U438 (.ZN( u0_subword_13 ) , .A3( u0_u2_n765 ) , .A2( u0_u2_n766 ) , .A1( u0_u2_n767 ) );
  NAND3_X1 u0_u2_U439 (.ZN( u0_subword_12 ) , .A3( u0_u2_n745 ) , .A2( u0_u2_n746 ) , .A1( u0_u2_n747 ) );
  NOR4_X1 u0_u2_U44 (.ZN( u0_u2_n568 ) , .A1( u0_u2_n660 ) , .A3( u0_u2_n668 ) , .A4( u0_u2_n692 ) , .A2( u0_u2_n775 ) );
  NAND3_X1 u0_u2_U440 (.A3( u0_u2_n682 ) , .A2( u0_u2_n683 ) , .A1( u0_u2_n684 ) , .ZN( u0_u2_n814 ) );
  NAND3_X1 u0_u2_U441 (.ZN( u0_u2_n645 ) , .A3( u0_u2_n715 ) , .A2( u0_u2_n731 ) , .A1( u0_u2_n799 ) );
  NAND3_X1 u0_u2_U442 (.A3( u0_u2_n625 ) , .A2( u0_u2_n626 ) , .A1( u0_u2_n627 ) , .ZN( u0_u2_n732 ) );
  NAND3_X1 u0_u2_U443 (.A3( u0_u2_n592 ) , .A2( u0_u2_n593 ) , .A1( u0_u2_n594 ) , .ZN( u0_u2_n628 ) );
  NAND3_X1 u0_u2_U444 (.ZN( u0_u2_n572 ) , .A3( u0_u2_n687 ) , .A2( u0_u2_n757 ) , .A1( u0_u2_n792 ) );
  NAND3_X1 u0_u2_U445 (.A3( u0_u2_n530 ) , .A2( u0_u2_n531 ) , .A1( u0_u2_n532 ) , .ZN( u0_u2_n749 ) );
  NAND3_X1 u0_u2_U446 (.A3( u0_u2_n519 ) , .A1( u0_u2_n520 ) , .ZN( u0_u2_n615 ) , .A2( u0_u2_n878 ) );
  NAND3_X1 u0_u2_U447 (.A3( u0_u2_n474 ) , .A2( u0_u2_n475 ) , .A1( u0_u2_n476 ) , .ZN( u0_u2_n784 ) );
  NOR2_X1 u0_u2_U448 (.ZN( u0_u2_n660 ) , .A1( u0_u2_n769 ) , .A2( u0_u2_n793 ) );
  NAND2_X1 u0_u2_U449 (.A2( u0_u2_n756 ) , .A1( u0_u2_n793 ) , .ZN( u0_u2_n816 ) );
  NOR4_X1 u0_u2_U45 (.A4( u0_u2_n559 ) , .A3( u0_u2_n560 ) , .A2( u0_u2_n561 ) , .A1( u0_u2_n562 ) , .ZN( u0_u2_n569 ) );
  NOR2_X1 u0_u2_U450 (.ZN( u0_u2_n561 ) , .A1( u0_u2_n793 ) , .A2( u0_u2_n820 ) );
  NOR2_X1 u0_u2_U451 (.ZN( u0_u2_n619 ) , .A1( u0_u2_n786 ) , .A2( u0_u2_n793 ) );
  NOR2_X1 u0_u2_U452 (.ZN( u0_u2_n724 ) , .A2( u0_u2_n751 ) , .A1( u0_u2_n793 ) );
  NOR2_X1 u0_u2_U453 (.ZN( u0_u2_n796 ) , .A2( u0_u2_n869 ) , .A1( u0_u2_n875 ) );
  NOR2_X1 u0_u2_U454 (.ZN( u0_u2_n708 ) , .A2( u0_u2_n793 ) , .A1( u0_u2_n824 ) );
  NOR2_X1 u0_u2_U455 (.A1( u0_u2_n737 ) , .ZN( u0_u2_n772 ) , .A2( u0_u2_n793 ) );
  INV_X1 u0_u2_U456 (.A( u0_u2_n793 ) , .ZN( u0_u2_n869 ) );
  NOR4_X1 u0_u2_U46 (.A4( u0_u2_n563 ) , .A3( u0_u2_n564 ) , .A2( u0_u2_n565 ) , .A1( u0_u2_n566 ) , .ZN( u0_u2_n567 ) );
  NOR4_X1 u0_u2_U47 (.A4( u0_u2_n516 ) , .A2( u0_u2_n517 ) , .A1( u0_u2_n518 ) , .ZN( u0_u2_n519 ) , .A3( u0_u2_n677 ) );
  INV_X1 u0_u2_U48 (.A( u0_u2_n512 ) , .ZN( u0_u2_n878 ) );
  NOR4_X1 u0_u2_U49 (.A4( u0_u2_n668 ) , .A3( u0_u2_n669 ) , .A2( u0_u2_n670 ) , .A1( u0_u2_n671 ) , .ZN( u0_u2_n684 ) );
  NOR3_X1 u0_u2_U5 (.ZN( u0_u2_n605 ) , .A1( u0_u2_n615 ) , .A3( u0_u2_n730 ) , .A2( u0_u2_n749 ) );
  NOR4_X1 u0_u2_U50 (.A4( u0_u2_n672 ) , .A3( u0_u2_n673 ) , .A2( u0_u2_n674 ) , .A1( u0_u2_n675 ) , .ZN( u0_u2_n683 ) );
  NOR2_X1 u0_u2_U51 (.ZN( u0_u2_n811 ) , .A1( u0_u2_n861 ) , .A2( u0_u2_n868 ) );
  NOR4_X1 u0_u2_U52 (.A1( u0_u2_n473 ) , .ZN( u0_u2_n474 ) , .A4( u0_u2_n549 ) , .A2( u0_u2_n561 ) , .A3( u0_u2_n621 ) );
  NAND4_X1 u0_u2_U53 (.A4( u0_u2_n492 ) , .A3( u0_u2_n493 ) , .A2( u0_u2_n494 ) , .A1( u0_u2_n495 ) , .ZN( u0_u2_n785 ) );
  NOR4_X1 u0_u2_U54 (.ZN( u0_u2_n492 ) , .A2( u0_u2_n540 ) , .A1( u0_u2_n565 ) , .A3( u0_u2_n638 ) , .A4( u0_u2_n725 ) );
  NOR4_X1 u0_u2_U55 (.A4( u0_u2_n521 ) , .A3( u0_u2_n522 ) , .A2( u0_u2_n523 ) , .A1( u0_u2_n524 ) , .ZN( u0_u2_n531 ) );
  NOR4_X1 u0_u2_U56 (.A3( u0_u2_n528 ) , .A1( u0_u2_n529 ) , .ZN( u0_u2_n530 ) , .A2( u0_u2_n680 ) , .A4( u0_u2_n776 ) );
  NOR2_X1 u0_u2_U57 (.ZN( u0_u2_n768 ) , .A1( u0_u2_n840 ) , .A2( u0_u2_n841 ) );
  NAND4_X1 u0_u2_U58 (.A4( u0_u2_n779 ) , .A3( u0_u2_n780 ) , .A2( u0_u2_n781 ) , .A1( u0_u2_n782 ) , .ZN( u0_u2_n808 ) );
  NOR3_X1 u0_u2_U59 (.A3( u0_u2_n772 ) , .A2( u0_u2_n773 ) , .A1( u0_u2_n774 ) , .ZN( u0_u2_n780 ) );
  NOR3_X1 u0_u2_U6 (.ZN( u0_u2_n511 ) , .A2( u0_u2_n686 ) , .A3( u0_u2_n784 ) , .A1( u0_u2_n883 ) );
  NOR4_X1 u0_u2_U60 (.A4( u0_u2_n775 ) , .A3( u0_u2_n776 ) , .A2( u0_u2_n777 ) , .A1( u0_u2_n778 ) , .ZN( u0_u2_n779 ) );
  AOI222_X1 u0_u2_U61 (.ZN( u0_u2_n782 ) , .A1( u0_u2_n837 ) , .C1( u0_u2_n841 ) , .B2( u0_u2_n848 ) , .A2( u0_u2_n857 ) , .B1( u0_u2_n868 ) , .C2( u0_u2_n880 ) );
  NAND4_X1 u0_u2_U62 (.A4( u0_u2_n480 ) , .A3( u0_u2_n481 ) , .A2( u0_u2_n482 ) , .A1( u0_u2_n483 ) , .ZN( u0_u2_n685 ) );
  NOR4_X1 u0_u2_U63 (.A4( u0_u2_n477 ) , .ZN( u0_u2_n483 ) , .A3( u0_u2_n563 ) , .A1( u0_u2_n742 ) , .A2( u0_u2_n762 ) );
  NOR4_X1 u0_u2_U64 (.ZN( u0_u2_n480 ) , .A2( u0_u2_n528 ) , .A4( u0_u2_n601 ) , .A1( u0_u2_n616 ) , .A3( u0_u2_n636 ) );
  NOR4_X1 u0_u2_U65 (.ZN( u0_u2_n481 ) , .A1( u0_u2_n513 ) , .A3( u0_u2_n551 ) , .A2( u0_u2_n590 ) , .A4( u0_u2_n723 ) );
  NAND4_X1 u0_u2_U66 (.A4( u0_u2_n463 ) , .A3( u0_u2_n464 ) , .A2( u0_u2_n465 ) , .A1( u0_u2_n466 ) , .ZN( u0_u2_n686 ) );
  NOR3_X1 u0_u2_U67 (.ZN( u0_u2_n464 ) , .A3( u0_u2_n537 ) , .A1( u0_u2_n562 ) , .A2( u0_u2_n577 ) );
  NOR4_X1 u0_u2_U68 (.ZN( u0_u2_n463 ) , .A2( u0_u2_n524 ) , .A1( u0_u2_n550 ) , .A3( u0_u2_n586 ) , .A4( u0_u2_n622 ) );
  NOR4_X1 u0_u2_U69 (.ZN( u0_u2_n465 ) , .A2( u0_u2_n516 ) , .A1( u0_u2_n606 ) , .A4( u0_u2_n635 ) , .A3( u0_u2_n718 ) );
  NOR3_X1 u0_u2_U7 (.A2( u0_u2_n614 ) , .A1( u0_u2_n615 ) , .ZN( u0_u2_n653 ) , .A3( u0_u2_n729 ) );
  NAND4_X1 u0_u2_U70 (.A4( u0_u2_n580 ) , .A3( u0_u2_n581 ) , .A1( u0_u2_n582 ) , .ZN( u0_u2_n730 ) , .A2( u0_u2_n881 ) );
  NOR4_X1 u0_u2_U71 (.A4( u0_u2_n576 ) , .A3( u0_u2_n577 ) , .A2( u0_u2_n578 ) , .A1( u0_u2_n579 ) , .ZN( u0_u2_n580 ) );
  AOI221_X1 u0_u2_U72 (.A( u0_u2_n571 ) , .C2( u0_u2_n572 ) , .ZN( u0_u2_n581 ) , .B2( u0_u2_n852 ) , .B1( u0_u2_n859 ) , .C1( u0_u2_n860 ) );
  INV_X1 u0_u2_U73 (.A( u0_u2_n614 ) , .ZN( u0_u2_n881 ) );
  NOR4_X1 u0_u2_U74 (.A4( u0_u2_n636 ) , .A3( u0_u2_n637 ) , .A2( u0_u2_n638 ) , .A1( u0_u2_n639 ) , .ZN( u0_u2_n640 ) );
  AOI211_X1 u0_u2_U75 (.B( u0_u2_n630 ) , .A( u0_u2_n631 ) , .ZN( u0_u2_n642 ) , .C2( u0_u2_n843 ) , .C1( u0_u2_n870 ) );
  NOR4_X1 u0_u2_U76 (.A4( u0_u2_n633 ) , .A3( u0_u2_n634 ) , .A2( u0_u2_n635 ) , .ZN( u0_u2_n641 ) , .A1( u0_u2_n671 ) );
  NAND4_X1 u0_u2_U77 (.A4( u0_u2_n542 ) , .A3( u0_u2_n543 ) , .A2( u0_u2_n544 ) , .A1( u0_u2_n545 ) , .ZN( u0_u2_n629 ) );
  NOR4_X1 u0_u2_U78 (.A4( u0_u2_n533 ) , .A2( u0_u2_n534 ) , .A1( u0_u2_n535 ) , .ZN( u0_u2_n545 ) , .A3( u0_u2_n708 ) );
  NOR4_X1 u0_u2_U79 (.A1( u0_u2_n538 ) , .ZN( u0_u2_n543 ) , .A2( u0_u2_n661 ) , .A4( u0_u2_n675 ) , .A3( u0_u2_n772 ) );
  NOR3_X1 u0_u2_U8 (.A3( u0_u2_n729 ) , .A1( u0_u2_n730 ) , .ZN( u0_u2_n747 ) , .A2( u0_u2_n748 ) );
  NOR4_X1 u0_u2_U80 (.A4( u0_u2_n536 ) , .A3( u0_u2_n537 ) , .ZN( u0_u2_n544 ) , .A2( u0_u2_n691 ) , .A1( u0_u2_n801 ) );
  NOR2_X1 u0_u2_U81 (.ZN( u0_u2_n755 ) , .A1( u0_u2_n868 ) , .A2( u0_u2_n869 ) );
  NAND4_X1 u0_u2_U82 (.A4( u0_u2_n555 ) , .A3( u0_u2_n556 ) , .A2( u0_u2_n557 ) , .A1( u0_u2_n558 ) , .ZN( u0_u2_n752 ) );
  NOR3_X1 u0_u2_U83 (.ZN( u0_u2_n556 ) , .A2( u0_u2_n658 ) , .A1( u0_u2_n674 ) , .A3( u0_u2_n778 ) );
  AOI211_X1 u0_u2_U84 (.B( u0_u2_n546 ) , .A( u0_u2_n547 ) , .ZN( u0_u2_n558 ) , .C2( u0_u2_n846 ) , .C1( u0_u2_n858 ) );
  NOR4_X1 u0_u2_U85 (.A4( u0_u2_n548 ) , .A3( u0_u2_n549 ) , .A2( u0_u2_n550 ) , .ZN( u0_u2_n557 ) , .A1( u0_u2_n695 ) );
  NOR4_X1 u0_u2_U86 (.A4( u0_u2_n616 ) , .A3( u0_u2_n617 ) , .A2( u0_u2_n618 ) , .A1( u0_u2_n619 ) , .ZN( u0_u2_n626 ) );
  NOR4_X1 u0_u2_U87 (.ZN( u0_u2_n627 ) , .A1( u0_u2_n663 ) , .A3( u0_u2_n673 ) , .A4( u0_u2_n689 ) , .A2( u0_u2_n773 ) );
  NOR2_X1 u0_u2_U88 (.ZN( u0_u2_n654 ) , .A1( u0_u2_n861 ) , .A2( u0_u2_n875 ) );
  INV_X1 u0_u2_U89 (.A( u0_u2_n813 ) , .ZN( u0_u2_n848 ) );
  NOR2_X1 u0_u2_U9 (.ZN( u0_u2_n582 ) , .A1( u0_u2_n629 ) , .A2( u0_u2_n752 ) );
  NAND4_X1 u0_u2_U90 (.A4( u0_u2_n726 ) , .A3( u0_u2_n727 ) , .A2( u0_u2_n728 ) , .ZN( u0_u2_n748 ) , .A1( u0_u2_n864 ) );
  NOR4_X1 u0_u2_U91 (.A4( u0_u2_n722 ) , .A3( u0_u2_n723 ) , .A2( u0_u2_n724 ) , .A1( u0_u2_n725 ) , .ZN( u0_u2_n726 ) );
  AOI221_X1 u0_u2_U92 (.A( u0_u2_n717 ) , .ZN( u0_u2_n728 ) , .C2( u0_u2_n851 ) , .B2( u0_u2_n852 ) , .C1( u0_u2_n868 ) , .B1( u0_u2_n869 ) );
  INV_X1 u0_u2_U93 (.A( u0_u2_n716 ) , .ZN( u0_u2_n864 ) );
  INV_X1 u0_u2_U94 (.A( u0_u2_n769 ) , .ZN( u0_u2_n837 ) );
  NAND2_X1 u0_u2_U95 (.A2( u0_u2_n769 ) , .A1( u0_u2_n813 ) , .ZN( u0_u2_n817 ) );
  OAI21_X1 u0_u2_U96 (.ZN( u0_u2_n738 ) , .A( u0_u2_n840 ) , .B2( u0_u2_n859 ) , .B1( u0_u2_n880 ) );
  OR4_X1 u0_u2_U97 (.A4( u0_u2_n525 ) , .A2( u0_u2_n526 ) , .A1( u0_u2_n527 ) , .ZN( u0_u2_n529 ) , .A3( u0_u2_n828 ) );
  OR4_X1 u0_u2_U98 (.A4( u0_u2_n573 ) , .A3( u0_u2_n574 ) , .A2( u0_u2_n575 ) , .ZN( u0_u2_n579 ) , .A1( u0_u2_n672 ) );
  OR4_X1 u0_u2_U99 (.A4( u0_u2_n689 ) , .A3( u0_u2_n690 ) , .A2( u0_u2_n691 ) , .A1( u0_u2_n692 ) , .ZN( u0_u2_n697 ) );
endmodule

