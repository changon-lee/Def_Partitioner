module des_des_die_1 ( u0_K10_10, u0_K10_13, u0_K10_14, u0_K10_18, u0_K10_41, u0_K8_19, u0_L0_1, u0_L0_10, u0_L0_16, 
       u0_L0_20, u0_L0_24, u0_L0_26, u0_L0_30, u0_L0_6, u0_L6_1, u0_L6_10, u0_L6_16, u0_L6_20, 
       u0_L6_24, u0_L6_26, u0_L6_30, u0_L6_6, u0_L8_12, u0_L8_13, u0_L8_16, u0_L8_17, u0_L8_18, 
       u0_L8_2, u0_L8_22, u0_L8_23, u0_L8_24, u0_L8_28, u0_L8_30, u0_L8_31, u0_L8_32, u0_L8_6, 
       u0_L8_7, u0_L8_9, u0_R0_10, u0_R0_11, u0_R0_12, u0_R0_13, u0_R0_14, u0_R0_15, u0_R0_16, 
       u0_R0_17, u0_R0_8, u0_R0_9, u0_R6_10, u0_R6_11, u0_R6_12, u0_R6_13, u0_R6_14, u0_R6_15, 
       u0_R6_16, u0_R6_17, u0_R6_8, u0_R6_9, u0_R8_1, u0_R8_10, u0_R8_11, u0_R8_12, u0_R8_13, 
       u0_R8_2, u0_R8_24, u0_R8_25, u0_R8_26, u0_R8_27, u0_R8_28, u0_R8_29, u0_R8_3, u0_R8_32, 
       u0_R8_4, u0_R8_5, u0_R8_6, u0_R8_7, u0_R8_8, u0_R8_9, u0_uk_K_r0_11, u0_uk_K_r0_19, u0_uk_K_r0_32, 
       u0_uk_K_r0_47, u0_uk_K_r11_8, u0_uk_K_r6_26, u0_uk_K_r6_34, u0_uk_K_r6_46, u0_uk_K_r8_17, u0_uk_K_r8_2, u0_uk_K_r8_22, u0_uk_K_r8_27, 
       u0_uk_K_r8_28, u0_uk_K_r8_32, u0_uk_K_r8_41, u0_uk_K_r8_44, u0_uk_K_r8_52, u0_uk_K_r8_8, u0_uk_n10, u0_uk_n100, u0_uk_n1009, 
       u0_uk_n102, u0_uk_n1021, u0_uk_n1024, u0_uk_n109, u0_uk_n11, u0_uk_n110, u0_uk_n117, u0_uk_n141, u0_uk_n142, 
       u0_uk_n146, u0_uk_n161, u0_uk_n162, u0_uk_n164, u0_uk_n182, u0_uk_n188, u0_uk_n202, u0_uk_n213, u0_uk_n214, 
       u0_uk_n217, u0_uk_n220, u0_uk_n223, u0_uk_n227, u0_uk_n228, u0_uk_n229, u0_uk_n230, u0_uk_n231, u0_uk_n234, 
       u0_uk_n235, u0_uk_n238, u0_uk_n239, u0_uk_n240, u0_uk_n243, u0_uk_n245, u0_uk_n246, u0_uk_n250, u0_uk_n251, 
       u0_uk_n252, u0_uk_n253, u0_uk_n254, u0_uk_n255, u0_uk_n257, u0_uk_n258, u0_uk_n262, u0_uk_n263, u0_uk_n266, 
       u0_uk_n267, u0_uk_n269, u0_uk_n318, u0_uk_n323, u0_uk_n329, u0_uk_n330, u0_uk_n331, u0_uk_n336, u0_uk_n337, 
       u0_uk_n340, u0_uk_n344, u0_uk_n345, u0_uk_n351, u0_uk_n352, u0_uk_n357, u0_uk_n358, u0_uk_n588, u0_uk_n589, 
       u0_uk_n596, u0_uk_n597, u0_uk_n598, u0_uk_n609, u0_uk_n610, u0_uk_n611, u0_uk_n614, u0_uk_n615, u0_uk_n619, 
       u0_uk_n620, u0_uk_n624, u0_uk_n625, u0_uk_n627, u0_uk_n63, u0_uk_n759, u0_uk_n83, u0_uk_n92, u0_uk_n93, 
       u0_uk_n94, u0_uk_n99, u1_L10_13, u1_L10_18, u1_L10_2, u1_L10_28, u1_L11_11, u1_L11_14, u1_L11_19, 
       u1_L11_25, u1_L11_29, u1_L11_3, u1_L11_4, u1_L11_8, u1_L12_12, u1_L12_15, u1_L12_21, u1_L12_22, 
       u1_L12_27, u1_L12_32, u1_L12_5, u1_L12_7, u1_L5_14, u1_L5_25, u1_L5_3, u1_L5_8, u1_L6_12, 
       u1_L6_22, u1_L6_32, u1_L6_7, u1_L7_11, u1_L7_12, u1_L7_19, u1_L7_22, u1_L7_29, u1_L7_32, 
       u1_L7_4, u1_L7_7, u1_L9_1, u1_L9_10, u1_L9_14, u1_L9_15, u1_L9_20, u1_L9_21, u1_L9_25, 
       u1_L9_26, u1_L9_27, u1_L9_3, u1_L9_5, u1_L9_8, u1_R10_4, u1_R10_5, u1_R10_6, u1_R10_7, 
       u1_R10_8, u1_R10_9, u1_R11_16, u1_R11_17, u1_R11_18, u1_R11_19, u1_R11_20, u1_R11_21, u1_R11_22, 
       u1_R11_23, u1_R11_24, u1_R11_25, u1_R12_1, u1_R12_24, u1_R12_25, u1_R12_26, u1_R12_27, u1_R12_28, 
       u1_R12_29, u1_R12_30, u1_R12_31, u1_R12_32, u1_R5_16, u1_R5_17, u1_R5_18, u1_R5_19, u1_R5_20, 
       u1_R5_21, u1_R6_24, u1_R6_25, u1_R6_26, u1_R6_27, u1_R6_28, u1_R6_29, u1_R7_20, u1_R7_21, 
       u1_R7_22, u1_R7_23, u1_R7_24, u1_R7_25, u1_R7_26, u1_R7_27, u1_R7_28, u1_R7_29, u1_R9_1, 
       u1_R9_12, u1_R9_13, u1_R9_14, u1_R9_15, u1_R9_16, u1_R9_17, u1_R9_18, u1_R9_19, u1_R9_20, 
       u1_R9_21, u1_R9_28, u1_R9_29, u1_R9_30, u1_R9_31, u1_R9_32, u1_uk_K_r10_11, u1_uk_K_r10_19, u1_uk_K_r11_21, 
       u1_uk_K_r11_28, u1_uk_K_r11_7, u1_uk_K_r12_15, u1_uk_K_r12_16, u1_uk_K_r12_21, u1_uk_K_r12_22, u1_uk_K_r5_23, u1_uk_K_r5_31, u1_uk_K_r5_43, 
       u1_uk_K_r5_7, u1_uk_K_r6_14, u1_uk_K_r6_22, u1_uk_K_r6_30, u1_uk_K_r6_31, u1_uk_K_r6_7, u1_uk_K_r7_1, u1_uk_K_r7_15, u1_uk_K_r7_16, 
       u1_uk_K_r7_22, u1_uk_K_r7_23, u1_uk_K_r7_30, u1_uk_K_r7_31, u1_uk_K_r7_7, u1_uk_K_r7_8, u1_uk_K_r9_0, u1_uk_K_r9_1, u1_uk_K_r9_10, 
       u1_uk_K_r9_13, u1_uk_K_r9_15, u1_uk_K_r9_19, u1_uk_K_r9_23, u1_uk_K_r9_27, u1_uk_K_r9_35, u1_uk_K_r9_4, u1_uk_K_r9_45, u1_uk_K_r9_48, 
       u1_uk_K_r9_5, u1_uk_K_r9_9, u1_uk_n10, u1_uk_n100, u1_uk_n11, u1_uk_n117, u1_uk_n118, u1_uk_n128, u1_uk_n141, 
       u1_uk_n145, u1_uk_n147, u1_uk_n148, u1_uk_n1489, u1_uk_n1490, u1_uk_n1500, u1_uk_n1501, u1_uk_n1510, u1_uk_n1520, 
       u1_uk_n1521, u1_uk_n1540, u1_uk_n1547, u1_uk_n155, u1_uk_n1555, u1_uk_n1556, u1_uk_n1560, u1_uk_n1561, u1_uk_n1566, 
       u1_uk_n1572, u1_uk_n1581, u1_uk_n1588, u1_uk_n1599, u1_uk_n1600, u1_uk_n1601, u1_uk_n1605, u1_uk_n1606, u1_uk_n1608, 
       u1_uk_n1612, u1_uk_n1613, u1_uk_n162, u1_uk_n163, u1_uk_n164, u1_uk_n1662, u1_uk_n1664, u1_uk_n1667, u1_uk_n1672, 
       u1_uk_n1677, u1_uk_n1682, u1_uk_n1683, u1_uk_n1684, u1_uk_n1687, u1_uk_n1689, u1_uk_n1690, u1_uk_n1695, u1_uk_n1696, 
       u1_uk_n1698, u1_uk_n17, u1_uk_n1703, u1_uk_n1704, u1_uk_n1713, u1_uk_n1718, u1_uk_n1719, u1_uk_n1731, u1_uk_n1739, 
       u1_uk_n1745, u1_uk_n1750, u1_uk_n1752, u1_uk_n1753, u1_uk_n1754, u1_uk_n1758, u1_uk_n1764, u1_uk_n1765, u1_uk_n1768, 
       u1_uk_n1772, u1_uk_n1775, u1_uk_n1776, u1_uk_n1777, u1_uk_n1782, u1_uk_n1783, u1_uk_n1784, u1_uk_n1790, u1_uk_n1793, 
       u1_uk_n1798, u1_uk_n1806, u1_uk_n1807, u1_uk_n1811, u1_uk_n1815, u1_uk_n1820, u1_uk_n1821, u1_uk_n1823, u1_uk_n1829, 
       u1_uk_n1830, u1_uk_n1832, u1_uk_n1836, u1_uk_n187, u1_uk_n191, u1_uk_n202, u1_uk_n203, u1_uk_n207, u1_uk_n208, 
       u1_uk_n213, u1_uk_n214, u1_uk_n222, u1_uk_n223, u1_uk_n238, u1_uk_n250, u1_uk_n27, u1_uk_n277, u1_uk_n279, 
       u1_uk_n286, u1_uk_n291, u1_uk_n292, u1_uk_n294, u1_uk_n297, u1_uk_n298, u1_uk_n31, u1_uk_n60, u1_uk_n63, 
       u1_uk_n83, u1_uk_n92, u1_uk_n93, u1_uk_n94, u1_uk_n99, u2_L8_1, u2_L8_10, u2_L8_20, u2_L8_26, 
       u2_R8_12, u2_R8_13, u2_R8_14, u2_R8_15, u2_R8_16, u2_R8_17, u2_uk_K_r8_13, u2_uk_K_r8_19, u2_uk_K_r8_40, 
       u2_uk_n10, u2_uk_n102, u2_uk_n117, u2_uk_n118, u2_uk_n129, u2_uk_n1590, u2_uk_n1599, u2_uk_n1603, u2_uk_n1613, 
       u2_uk_n1629, u2_uk_n1630, u2_uk_n182, u2_uk_n187, u2_uk_n257, u2_uk_n27, u0_N224, u0_N229, u0_N233, u0_N239, u0_N243, u0_N247, u0_N249, u0_N253, u0_N289, 
        u0_N293, u0_N294, u0_N296, u0_N299, u0_N300, u0_N303, u0_N304, u0_N305, u0_N309, 
        u0_N310, u0_N311, u0_N315, u0_N317, u0_N318, u0_N319, u0_N32, u0_N37, u0_N41, 
        u0_N47, u0_N51, u0_N55, u0_N57, u0_N61, u0_uk_n942, u1_N194, u1_N199, u1_N205, 
        u1_N216, u1_N230, u1_N235, u1_N245, u1_N255, u1_N259, u1_N262, u1_N266, u1_N267, 
        u1_N274, u1_N277, u1_N284, u1_N287, u1_N320, u1_N322, u1_N324, u1_N327, u1_N329, 
        u1_N333, u1_N334, u1_N339, u1_N340, u1_N344, u1_N345, u1_N346, u1_N353, u1_N364, 
        u1_N369, u1_N379, u1_N386, u1_N387, u1_N391, u1_N394, u1_N397, u1_N402, u1_N408, 
        u1_N412, u1_N420, u1_N422, u1_N427, u1_N430, u1_N436, u1_N437, u1_N442, u1_N447, 
        u1_uk_n102, u1_uk_n109, u1_uk_n129, u1_uk_n146, u1_uk_n161, u1_uk_n182, u1_uk_n188, u1_uk_n230, u1_uk_n231, 
        u1_uk_n251, u1_uk_n252, u1_uk_n257, u2_N288, u2_N297, u2_N307, u2_N313 );
  input u0_K10_10, u0_K10_13, u0_K10_14, u0_K10_18, u0_K10_41, u0_K8_19, u0_L0_1, u0_L0_10, u0_L0_16, 
        u0_L0_20, u0_L0_24, u0_L0_26, u0_L0_30, u0_L0_6, u0_L6_1, u0_L6_10, u0_L6_16, u0_L6_20, 
        u0_L6_24, u0_L6_26, u0_L6_30, u0_L6_6, u0_L8_12, u0_L8_13, u0_L8_16, u0_L8_17, u0_L8_18, 
        u0_L8_2, u0_L8_22, u0_L8_23, u0_L8_24, u0_L8_28, u0_L8_30, u0_L8_31, u0_L8_32, u0_L8_6, 
        u0_L8_7, u0_L8_9, u0_R0_10, u0_R0_11, u0_R0_12, u0_R0_13, u0_R0_14, u0_R0_15, u0_R0_16, 
        u0_R0_17, u0_R0_8, u0_R0_9, u0_R6_10, u0_R6_11, u0_R6_12, u0_R6_13, u0_R6_14, u0_R6_15, 
        u0_R6_16, u0_R6_17, u0_R6_8, u0_R6_9, u0_R8_1, u0_R8_10, u0_R8_11, u0_R8_12, u0_R8_13, 
        u0_R8_2, u0_R8_24, u0_R8_25, u0_R8_26, u0_R8_27, u0_R8_28, u0_R8_29, u0_R8_3, u0_R8_32, 
        u0_R8_4, u0_R8_5, u0_R8_6, u0_R8_7, u0_R8_8, u0_R8_9, u0_uk_K_r0_11, u0_uk_K_r0_19, u0_uk_K_r0_32, 
        u0_uk_K_r0_47, u0_uk_K_r11_8, u0_uk_K_r6_26, u0_uk_K_r6_34, u0_uk_K_r6_46, u0_uk_K_r8_17, u0_uk_K_r8_2, u0_uk_K_r8_22, u0_uk_K_r8_27, 
        u0_uk_K_r8_28, u0_uk_K_r8_32, u0_uk_K_r8_41, u0_uk_K_r8_44, u0_uk_K_r8_52, u0_uk_K_r8_8, u0_uk_n10, u0_uk_n100, u0_uk_n1009, 
        u0_uk_n102, u0_uk_n1021, u0_uk_n1024, u0_uk_n109, u0_uk_n11, u0_uk_n110, u0_uk_n117, u0_uk_n141, u0_uk_n142, 
        u0_uk_n146, u0_uk_n161, u0_uk_n162, u0_uk_n164, u0_uk_n182, u0_uk_n188, u0_uk_n202, u0_uk_n213, u0_uk_n214, 
        u0_uk_n217, u0_uk_n220, u0_uk_n223, u0_uk_n227, u0_uk_n228, u0_uk_n229, u0_uk_n230, u0_uk_n231, u0_uk_n234, 
        u0_uk_n235, u0_uk_n238, u0_uk_n239, u0_uk_n240, u0_uk_n243, u0_uk_n245, u0_uk_n246, u0_uk_n250, u0_uk_n251, 
        u0_uk_n252, u0_uk_n253, u0_uk_n254, u0_uk_n255, u0_uk_n257, u0_uk_n258, u0_uk_n262, u0_uk_n263, u0_uk_n266, 
        u0_uk_n267, u0_uk_n269, u0_uk_n318, u0_uk_n323, u0_uk_n329, u0_uk_n330, u0_uk_n331, u0_uk_n336, u0_uk_n337, 
        u0_uk_n340, u0_uk_n344, u0_uk_n345, u0_uk_n351, u0_uk_n352, u0_uk_n357, u0_uk_n358, u0_uk_n588, u0_uk_n589, 
        u0_uk_n596, u0_uk_n597, u0_uk_n598, u0_uk_n609, u0_uk_n610, u0_uk_n611, u0_uk_n614, u0_uk_n615, u0_uk_n619, 
        u0_uk_n620, u0_uk_n624, u0_uk_n625, u0_uk_n627, u0_uk_n63, u0_uk_n759, u0_uk_n83, u0_uk_n92, u0_uk_n93, 
        u0_uk_n94, u0_uk_n99, u1_L10_13, u1_L10_18, u1_L10_2, u1_L10_28, u1_L11_11, u1_L11_14, u1_L11_19, 
        u1_L11_25, u1_L11_29, u1_L11_3, u1_L11_4, u1_L11_8, u1_L12_12, u1_L12_15, u1_L12_21, u1_L12_22, 
        u1_L12_27, u1_L12_32, u1_L12_5, u1_L12_7, u1_L5_14, u1_L5_25, u1_L5_3, u1_L5_8, u1_L6_12, 
        u1_L6_22, u1_L6_32, u1_L6_7, u1_L7_11, u1_L7_12, u1_L7_19, u1_L7_22, u1_L7_29, u1_L7_32, 
        u1_L7_4, u1_L7_7, u1_L9_1, u1_L9_10, u1_L9_14, u1_L9_15, u1_L9_20, u1_L9_21, u1_L9_25, 
        u1_L9_26, u1_L9_27, u1_L9_3, u1_L9_5, u1_L9_8, u1_R10_4, u1_R10_5, u1_R10_6, u1_R10_7, 
        u1_R10_8, u1_R10_9, u1_R11_16, u1_R11_17, u1_R11_18, u1_R11_19, u1_R11_20, u1_R11_21, u1_R11_22, 
        u1_R11_23, u1_R11_24, u1_R11_25, u1_R12_1, u1_R12_24, u1_R12_25, u1_R12_26, u1_R12_27, u1_R12_28, 
        u1_R12_29, u1_R12_30, u1_R12_31, u1_R12_32, u1_R5_16, u1_R5_17, u1_R5_18, u1_R5_19, u1_R5_20, 
        u1_R5_21, u1_R6_24, u1_R6_25, u1_R6_26, u1_R6_27, u1_R6_28, u1_R6_29, u1_R7_20, u1_R7_21, 
        u1_R7_22, u1_R7_23, u1_R7_24, u1_R7_25, u1_R7_26, u1_R7_27, u1_R7_28, u1_R7_29, u1_R9_1, 
        u1_R9_12, u1_R9_13, u1_R9_14, u1_R9_15, u1_R9_16, u1_R9_17, u1_R9_18, u1_R9_19, u1_R9_20, 
        u1_R9_21, u1_R9_28, u1_R9_29, u1_R9_30, u1_R9_31, u1_R9_32, u1_uk_K_r10_11, u1_uk_K_r10_19, u1_uk_K_r11_21, 
        u1_uk_K_r11_28, u1_uk_K_r11_7, u1_uk_K_r12_15, u1_uk_K_r12_16, u1_uk_K_r12_21, u1_uk_K_r12_22, u1_uk_K_r5_23, u1_uk_K_r5_31, u1_uk_K_r5_43, 
        u1_uk_K_r5_7, u1_uk_K_r6_14, u1_uk_K_r6_22, u1_uk_K_r6_30, u1_uk_K_r6_31, u1_uk_K_r6_7, u1_uk_K_r7_1, u1_uk_K_r7_15, u1_uk_K_r7_16, 
        u1_uk_K_r7_22, u1_uk_K_r7_23, u1_uk_K_r7_30, u1_uk_K_r7_31, u1_uk_K_r7_7, u1_uk_K_r7_8, u1_uk_K_r9_0, u1_uk_K_r9_1, u1_uk_K_r9_10, 
        u1_uk_K_r9_13, u1_uk_K_r9_15, u1_uk_K_r9_19, u1_uk_K_r9_23, u1_uk_K_r9_27, u1_uk_K_r9_35, u1_uk_K_r9_4, u1_uk_K_r9_45, u1_uk_K_r9_48, 
        u1_uk_K_r9_5, u1_uk_K_r9_9, u1_uk_n10, u1_uk_n100, u1_uk_n11, u1_uk_n117, u1_uk_n118, u1_uk_n128, u1_uk_n141, 
        u1_uk_n145, u1_uk_n147, u1_uk_n148, u1_uk_n1489, u1_uk_n1490, u1_uk_n1500, u1_uk_n1501, u1_uk_n1510, u1_uk_n1520, 
        u1_uk_n1521, u1_uk_n1540, u1_uk_n1547, u1_uk_n155, u1_uk_n1555, u1_uk_n1556, u1_uk_n1560, u1_uk_n1561, u1_uk_n1566, 
        u1_uk_n1572, u1_uk_n1581, u1_uk_n1588, u1_uk_n1599, u1_uk_n1600, u1_uk_n1601, u1_uk_n1605, u1_uk_n1606, u1_uk_n1608, 
        u1_uk_n1612, u1_uk_n1613, u1_uk_n162, u1_uk_n163, u1_uk_n164, u1_uk_n1662, u1_uk_n1664, u1_uk_n1667, u1_uk_n1672, 
        u1_uk_n1677, u1_uk_n1682, u1_uk_n1683, u1_uk_n1684, u1_uk_n1687, u1_uk_n1689, u1_uk_n1690, u1_uk_n1695, u1_uk_n1696, 
        u1_uk_n1698, u1_uk_n17, u1_uk_n1703, u1_uk_n1704, u1_uk_n1713, u1_uk_n1718, u1_uk_n1719, u1_uk_n1731, u1_uk_n1739, 
        u1_uk_n1745, u1_uk_n1750, u1_uk_n1752, u1_uk_n1753, u1_uk_n1754, u1_uk_n1758, u1_uk_n1764, u1_uk_n1765, u1_uk_n1768, 
        u1_uk_n1772, u1_uk_n1775, u1_uk_n1776, u1_uk_n1777, u1_uk_n1782, u1_uk_n1783, u1_uk_n1784, u1_uk_n1790, u1_uk_n1793, 
        u1_uk_n1798, u1_uk_n1806, u1_uk_n1807, u1_uk_n1811, u1_uk_n1815, u1_uk_n1820, u1_uk_n1821, u1_uk_n1823, u1_uk_n1829, 
        u1_uk_n1830, u1_uk_n1832, u1_uk_n1836, u1_uk_n187, u1_uk_n191, u1_uk_n202, u1_uk_n203, u1_uk_n207, u1_uk_n208, 
        u1_uk_n213, u1_uk_n214, u1_uk_n222, u1_uk_n223, u1_uk_n238, u1_uk_n250, u1_uk_n27, u1_uk_n277, u1_uk_n279, 
        u1_uk_n286, u1_uk_n291, u1_uk_n292, u1_uk_n294, u1_uk_n297, u1_uk_n298, u1_uk_n31, u1_uk_n60, u1_uk_n63, 
        u1_uk_n83, u1_uk_n92, u1_uk_n93, u1_uk_n94, u1_uk_n99, u2_L8_1, u2_L8_10, u2_L8_20, u2_L8_26, 
        u2_R8_12, u2_R8_13, u2_R8_14, u2_R8_15, u2_R8_16, u2_R8_17, u2_uk_K_r8_13, u2_uk_K_r8_19, u2_uk_K_r8_40, 
        u2_uk_n10, u2_uk_n102, u2_uk_n117, u2_uk_n118, u2_uk_n129, u2_uk_n1590, u2_uk_n1599, u2_uk_n1603, u2_uk_n1613, 
        u2_uk_n1629, u2_uk_n1630, u2_uk_n182, u2_uk_n187, u2_uk_n257, u2_uk_n27;
  output u0_N224, u0_N229, u0_N233, u0_N239, u0_N243, u0_N247, u0_N249, u0_N253, u0_N289, 
        u0_N293, u0_N294, u0_N296, u0_N299, u0_N300, u0_N303, u0_N304, u0_N305, u0_N309, 
        u0_N310, u0_N311, u0_N315, u0_N317, u0_N318, u0_N319, u0_N32, u0_N37, u0_N41, 
        u0_N47, u0_N51, u0_N55, u0_N57, u0_N61, u0_uk_n942, u1_N194, u1_N199, u1_N205, 
        u1_N216, u1_N230, u1_N235, u1_N245, u1_N255, u1_N259, u1_N262, u1_N266, u1_N267, 
        u1_N274, u1_N277, u1_N284, u1_N287, u1_N320, u1_N322, u1_N324, u1_N327, u1_N329, 
        u1_N333, u1_N334, u1_N339, u1_N340, u1_N344, u1_N345, u1_N346, u1_N353, u1_N364, 
        u1_N369, u1_N379, u1_N386, u1_N387, u1_N391, u1_N394, u1_N397, u1_N402, u1_N408, 
        u1_N412, u1_N420, u1_N422, u1_N427, u1_N430, u1_N436, u1_N437, u1_N442, u1_N447, 
        u1_uk_n102, u1_uk_n109, u1_uk_n129, u1_uk_n146, u1_uk_n161, u1_uk_n182, u1_uk_n188, u1_uk_n230, u1_uk_n231, 
        u1_uk_n251, u1_uk_n252, u1_uk_n257, u2_N288, u2_N297, u2_N307, u2_N313;
  wire u0_K10_1, u0_K10_11, u0_K10_12, u0_K10_15, u0_K10_16, u0_K10_17, u0_K10_2, u0_K10_3, u0_K10_37, 
       u0_K10_38, u0_K10_39, u0_K10_4, u0_K10_40, u0_K10_42, u0_K10_5, u0_K10_6, u0_K10_7, u0_K10_8, 
       u0_K10_9, u0_K2_13, u0_K2_14, u0_K2_15, u0_K2_16, u0_K2_17, u0_K2_18, u0_K2_19, u0_K2_20, 
       u0_K2_21, u0_K2_22, u0_K2_23, u0_K2_24, u0_K8_13, u0_K8_14, u0_K8_15, u0_K8_16, u0_K8_17, 
       u0_K8_18, u0_K8_20, u0_K8_21, u0_K8_22, u0_K8_23, u0_K8_24, u0_out1_1, u0_out1_10, u0_out1_16, 
       u0_out1_20, u0_out1_24, u0_out1_26, u0_out1_30, u0_out1_6, u0_out7_1, u0_out7_10, u0_out7_16, u0_out7_20, 
       u0_out7_24, u0_out7_26, u0_out7_30, u0_out7_6, u0_out9_12, u0_out9_13, u0_out9_16, u0_out9_17, u0_out9_18, 
       u0_out9_2, u0_out9_22, u0_out9_23, u0_out9_24, u0_out9_28, u0_out9_30, u0_out9_31, u0_out9_32, u0_out9_6, 
       u0_out9_7, u0_out9_9, u0_u1_X_13, u0_u1_X_14, u0_u1_X_15, u0_u1_X_16, u0_u1_X_17, u0_u1_X_18, u0_u1_X_19, 
       u0_u1_X_20, u0_u1_X_21, u0_u1_X_22, u0_u1_X_23, u0_u1_X_24, u0_u1_u2_n100, u0_u1_u2_n101, u0_u1_u2_n102, u0_u1_u2_n103, 
       u0_u1_u2_n104, u0_u1_u2_n105, u0_u1_u2_n106, u0_u1_u2_n107, u0_u1_u2_n108, u0_u1_u2_n109, u0_u1_u2_n110, u0_u1_u2_n111, u0_u1_u2_n112, 
       u0_u1_u2_n113, u0_u1_u2_n114, u0_u1_u2_n115, u0_u1_u2_n116, u0_u1_u2_n117, u0_u1_u2_n118, u0_u1_u2_n119, u0_u1_u2_n120, u0_u1_u2_n121, 
       u0_u1_u2_n122, u0_u1_u2_n123, u0_u1_u2_n124, u0_u1_u2_n125, u0_u1_u2_n126, u0_u1_u2_n127, u0_u1_u2_n128, u0_u1_u2_n129, u0_u1_u2_n130, 
       u0_u1_u2_n131, u0_u1_u2_n132, u0_u1_u2_n133, u0_u1_u2_n134, u0_u1_u2_n135, u0_u1_u2_n136, u0_u1_u2_n137, u0_u1_u2_n138, u0_u1_u2_n139, 
       u0_u1_u2_n140, u0_u1_u2_n141, u0_u1_u2_n142, u0_u1_u2_n143, u0_u1_u2_n144, u0_u1_u2_n145, u0_u1_u2_n146, u0_u1_u2_n147, u0_u1_u2_n148, 
       u0_u1_u2_n149, u0_u1_u2_n150, u0_u1_u2_n151, u0_u1_u2_n152, u0_u1_u2_n153, u0_u1_u2_n154, u0_u1_u2_n155, u0_u1_u2_n156, u0_u1_u2_n157, 
       u0_u1_u2_n158, u0_u1_u2_n159, u0_u1_u2_n160, u0_u1_u2_n161, u0_u1_u2_n162, u0_u1_u2_n163, u0_u1_u2_n164, u0_u1_u2_n165, u0_u1_u2_n166, 
       u0_u1_u2_n167, u0_u1_u2_n168, u0_u1_u2_n169, u0_u1_u2_n170, u0_u1_u2_n171, u0_u1_u2_n172, u0_u1_u2_n173, u0_u1_u2_n174, u0_u1_u2_n175, 
       u0_u1_u2_n176, u0_u1_u2_n177, u0_u1_u2_n178, u0_u1_u2_n179, u0_u1_u2_n180, u0_u1_u2_n181, u0_u1_u2_n182, u0_u1_u2_n183, u0_u1_u2_n184, 
       u0_u1_u2_n185, u0_u1_u2_n186, u0_u1_u2_n187, u0_u1_u2_n188, u0_u1_u2_n95, u0_u1_u2_n96, u0_u1_u2_n97, u0_u1_u2_n98, u0_u1_u2_n99, 
       u0_u1_u3_n100, u0_u1_u3_n101, u0_u1_u3_n102, u0_u1_u3_n103, u0_u1_u3_n104, u0_u1_u3_n105, u0_u1_u3_n106, u0_u1_u3_n107, u0_u1_u3_n108, 
       u0_u1_u3_n109, u0_u1_u3_n110, u0_u1_u3_n111, u0_u1_u3_n112, u0_u1_u3_n113, u0_u1_u3_n114, u0_u1_u3_n115, u0_u1_u3_n116, u0_u1_u3_n117, 
       u0_u1_u3_n118, u0_u1_u3_n119, u0_u1_u3_n120, u0_u1_u3_n121, u0_u1_u3_n122, u0_u1_u3_n123, u0_u1_u3_n124, u0_u1_u3_n125, u0_u1_u3_n126, 
       u0_u1_u3_n127, u0_u1_u3_n128, u0_u1_u3_n129, u0_u1_u3_n130, u0_u1_u3_n131, u0_u1_u3_n132, u0_u1_u3_n133, u0_u1_u3_n134, u0_u1_u3_n135, 
       u0_u1_u3_n136, u0_u1_u3_n137, u0_u1_u3_n138, u0_u1_u3_n139, u0_u1_u3_n140, u0_u1_u3_n141, u0_u1_u3_n142, u0_u1_u3_n143, u0_u1_u3_n144, 
       u0_u1_u3_n145, u0_u1_u3_n146, u0_u1_u3_n147, u0_u1_u3_n148, u0_u1_u3_n149, u0_u1_u3_n150, u0_u1_u3_n151, u0_u1_u3_n152, u0_u1_u3_n153, 
       u0_u1_u3_n154, u0_u1_u3_n155, u0_u1_u3_n156, u0_u1_u3_n157, u0_u1_u3_n158, u0_u1_u3_n159, u0_u1_u3_n160, u0_u1_u3_n161, u0_u1_u3_n162, 
       u0_u1_u3_n163, u0_u1_u3_n164, u0_u1_u3_n165, u0_u1_u3_n166, u0_u1_u3_n167, u0_u1_u3_n168, u0_u1_u3_n169, u0_u1_u3_n170, u0_u1_u3_n171, 
       u0_u1_u3_n172, u0_u1_u3_n173, u0_u1_u3_n174, u0_u1_u3_n175, u0_u1_u3_n176, u0_u1_u3_n177, u0_u1_u3_n178, u0_u1_u3_n179, u0_u1_u3_n180, 
       u0_u1_u3_n181, u0_u1_u3_n182, u0_u1_u3_n183, u0_u1_u3_n184, u0_u1_u3_n185, u0_u1_u3_n186, u0_u1_u3_n94, u0_u1_u3_n95, u0_u1_u3_n96, 
       u0_u1_u3_n97, u0_u1_u3_n98, u0_u1_u3_n99, u0_u7_X_13, u0_u7_X_14, u0_u7_X_15, u0_u7_X_16, u0_u7_X_17, u0_u7_X_18, 
       u0_u7_X_19, u0_u7_X_20, u0_u7_X_21, u0_u7_X_22, u0_u7_X_23, u0_u7_X_24, u0_u7_u2_n100, u0_u7_u2_n101, u0_u7_u2_n102, 
       u0_u7_u2_n103, u0_u7_u2_n104, u0_u7_u2_n105, u0_u7_u2_n106, u0_u7_u2_n107, u0_u7_u2_n108, u0_u7_u2_n109, u0_u7_u2_n110, u0_u7_u2_n111, 
       u0_u7_u2_n112, u0_u7_u2_n113, u0_u7_u2_n114, u0_u7_u2_n115, u0_u7_u2_n116, u0_u7_u2_n117, u0_u7_u2_n118, u0_u7_u2_n119, u0_u7_u2_n120, 
       u0_u7_u2_n121, u0_u7_u2_n122, u0_u7_u2_n123, u0_u7_u2_n124, u0_u7_u2_n125, u0_u7_u2_n126, u0_u7_u2_n127, u0_u7_u2_n128, u0_u7_u2_n129, 
       u0_u7_u2_n130, u0_u7_u2_n131, u0_u7_u2_n132, u0_u7_u2_n133, u0_u7_u2_n134, u0_u7_u2_n135, u0_u7_u2_n136, u0_u7_u2_n137, u0_u7_u2_n138, 
       u0_u7_u2_n139, u0_u7_u2_n140, u0_u7_u2_n141, u0_u7_u2_n142, u0_u7_u2_n143, u0_u7_u2_n144, u0_u7_u2_n145, u0_u7_u2_n146, u0_u7_u2_n147, 
       u0_u7_u2_n148, u0_u7_u2_n149, u0_u7_u2_n150, u0_u7_u2_n151, u0_u7_u2_n152, u0_u7_u2_n153, u0_u7_u2_n154, u0_u7_u2_n155, u0_u7_u2_n156, 
       u0_u7_u2_n157, u0_u7_u2_n158, u0_u7_u2_n159, u0_u7_u2_n160, u0_u7_u2_n161, u0_u7_u2_n162, u0_u7_u2_n163, u0_u7_u2_n164, u0_u7_u2_n165, 
       u0_u7_u2_n166, u0_u7_u2_n167, u0_u7_u2_n168, u0_u7_u2_n169, u0_u7_u2_n170, u0_u7_u2_n171, u0_u7_u2_n172, u0_u7_u2_n173, u0_u7_u2_n174, 
       u0_u7_u2_n175, u0_u7_u2_n176, u0_u7_u2_n177, u0_u7_u2_n178, u0_u7_u2_n179, u0_u7_u2_n180, u0_u7_u2_n181, u0_u7_u2_n182, u0_u7_u2_n183, 
       u0_u7_u2_n184, u0_u7_u2_n185, u0_u7_u2_n186, u0_u7_u2_n187, u0_u7_u2_n188, u0_u7_u2_n95, u0_u7_u2_n96, u0_u7_u2_n97, u0_u7_u2_n98, 
       u0_u7_u2_n99, u0_u7_u3_n100, u0_u7_u3_n101, u0_u7_u3_n102, u0_u7_u3_n103, u0_u7_u3_n104, u0_u7_u3_n105, u0_u7_u3_n106, u0_u7_u3_n107, 
       u0_u7_u3_n108, u0_u7_u3_n109, u0_u7_u3_n110, u0_u7_u3_n111, u0_u7_u3_n112, u0_u7_u3_n113, u0_u7_u3_n114, u0_u7_u3_n115, u0_u7_u3_n116, 
       u0_u7_u3_n117, u0_u7_u3_n118, u0_u7_u3_n119, u0_u7_u3_n120, u0_u7_u3_n121, u0_u7_u3_n122, u0_u7_u3_n123, u0_u7_u3_n124, u0_u7_u3_n125, 
       u0_u7_u3_n126, u0_u7_u3_n127, u0_u7_u3_n128, u0_u7_u3_n129, u0_u7_u3_n130, u0_u7_u3_n131, u0_u7_u3_n132, u0_u7_u3_n133, u0_u7_u3_n134, 
       u0_u7_u3_n135, u0_u7_u3_n136, u0_u7_u3_n137, u0_u7_u3_n138, u0_u7_u3_n139, u0_u7_u3_n140, u0_u7_u3_n141, u0_u7_u3_n142, u0_u7_u3_n143, 
       u0_u7_u3_n144, u0_u7_u3_n145, u0_u7_u3_n146, u0_u7_u3_n147, u0_u7_u3_n148, u0_u7_u3_n149, u0_u7_u3_n150, u0_u7_u3_n151, u0_u7_u3_n152, 
       u0_u7_u3_n153, u0_u7_u3_n154, u0_u7_u3_n155, u0_u7_u3_n156, u0_u7_u3_n157, u0_u7_u3_n158, u0_u7_u3_n159, u0_u7_u3_n160, u0_u7_u3_n161, 
       u0_u7_u3_n162, u0_u7_u3_n163, u0_u7_u3_n164, u0_u7_u3_n165, u0_u7_u3_n166, u0_u7_u3_n167, u0_u7_u3_n168, u0_u7_u3_n169, u0_u7_u3_n170, 
       u0_u7_u3_n171, u0_u7_u3_n172, u0_u7_u3_n173, u0_u7_u3_n174, u0_u7_u3_n175, u0_u7_u3_n176, u0_u7_u3_n177, u0_u7_u3_n178, u0_u7_u3_n179, 
       u0_u7_u3_n180, u0_u7_u3_n181, u0_u7_u3_n182, u0_u7_u3_n183, u0_u7_u3_n184, u0_u7_u3_n185, u0_u7_u3_n186, u0_u7_u3_n94, u0_u7_u3_n95, 
       u0_u7_u3_n96, u0_u7_u3_n97, u0_u7_u3_n98, u0_u7_u3_n99, u0_u9_X_1, u0_u9_X_10, u0_u9_X_11, u0_u9_X_12, u0_u9_X_13, 
       u0_u9_X_14, u0_u9_X_15, u0_u9_X_16, u0_u9_X_17, u0_u9_X_18, u0_u9_X_2, u0_u9_X_3, u0_u9_X_37, u0_u9_X_38, 
       u0_u9_X_39, u0_u9_X_4, u0_u9_X_40, u0_u9_X_41, u0_u9_X_42, u0_u9_X_5, u0_u9_X_6, u0_u9_X_7, u0_u9_X_8, 
       u0_u9_X_9, u0_u9_u0_n100, u0_u9_u0_n101, u0_u9_u0_n102, u0_u9_u0_n103, u0_u9_u0_n104, u0_u9_u0_n105, u0_u9_u0_n106, u0_u9_u0_n107, 
       u0_u9_u0_n108, u0_u9_u0_n109, u0_u9_u0_n110, u0_u9_u0_n111, u0_u9_u0_n112, u0_u9_u0_n113, u0_u9_u0_n114, u0_u9_u0_n115, u0_u9_u0_n116, 
       u0_u9_u0_n117, u0_u9_u0_n118, u0_u9_u0_n119, u0_u9_u0_n120, u0_u9_u0_n121, u0_u9_u0_n122, u0_u9_u0_n123, u0_u9_u0_n124, u0_u9_u0_n125, 
       u0_u9_u0_n126, u0_u9_u0_n127, u0_u9_u0_n128, u0_u9_u0_n129, u0_u9_u0_n130, u0_u9_u0_n131, u0_u9_u0_n132, u0_u9_u0_n133, u0_u9_u0_n134, 
       u0_u9_u0_n135, u0_u9_u0_n136, u0_u9_u0_n137, u0_u9_u0_n138, u0_u9_u0_n139, u0_u9_u0_n140, u0_u9_u0_n141, u0_u9_u0_n142, u0_u9_u0_n143, 
       u0_u9_u0_n144, u0_u9_u0_n145, u0_u9_u0_n146, u0_u9_u0_n147, u0_u9_u0_n148, u0_u9_u0_n149, u0_u9_u0_n150, u0_u9_u0_n151, u0_u9_u0_n152, 
       u0_u9_u0_n153, u0_u9_u0_n154, u0_u9_u0_n155, u0_u9_u0_n156, u0_u9_u0_n157, u0_u9_u0_n158, u0_u9_u0_n159, u0_u9_u0_n160, u0_u9_u0_n161, 
       u0_u9_u0_n162, u0_u9_u0_n163, u0_u9_u0_n164, u0_u9_u0_n165, u0_u9_u0_n166, u0_u9_u0_n167, u0_u9_u0_n168, u0_u9_u0_n169, u0_u9_u0_n170, 
       u0_u9_u0_n171, u0_u9_u0_n172, u0_u9_u0_n173, u0_u9_u0_n174, u0_u9_u0_n88, u0_u9_u0_n89, u0_u9_u0_n90, u0_u9_u0_n91, u0_u9_u0_n92, 
       u0_u9_u0_n93, u0_u9_u0_n94, u0_u9_u0_n95, u0_u9_u0_n96, u0_u9_u0_n97, u0_u9_u0_n98, u0_u9_u0_n99, u0_u9_u1_n100, u0_u9_u1_n101, 
       u0_u9_u1_n102, u0_u9_u1_n103, u0_u9_u1_n104, u0_u9_u1_n105, u0_u9_u1_n106, u0_u9_u1_n107, u0_u9_u1_n108, u0_u9_u1_n109, u0_u9_u1_n110, 
       u0_u9_u1_n111, u0_u9_u1_n112, u0_u9_u1_n113, u0_u9_u1_n114, u0_u9_u1_n115, u0_u9_u1_n116, u0_u9_u1_n117, u0_u9_u1_n118, u0_u9_u1_n119, 
       u0_u9_u1_n120, u0_u9_u1_n121, u0_u9_u1_n122, u0_u9_u1_n123, u0_u9_u1_n124, u0_u9_u1_n125, u0_u9_u1_n126, u0_u9_u1_n127, u0_u9_u1_n128, 
       u0_u9_u1_n129, u0_u9_u1_n130, u0_u9_u1_n131, u0_u9_u1_n132, u0_u9_u1_n133, u0_u9_u1_n134, u0_u9_u1_n135, u0_u9_u1_n136, u0_u9_u1_n137, 
       u0_u9_u1_n138, u0_u9_u1_n139, u0_u9_u1_n140, u0_u9_u1_n141, u0_u9_u1_n142, u0_u9_u1_n143, u0_u9_u1_n144, u0_u9_u1_n145, u0_u9_u1_n146, 
       u0_u9_u1_n147, u0_u9_u1_n148, u0_u9_u1_n149, u0_u9_u1_n150, u0_u9_u1_n151, u0_u9_u1_n152, u0_u9_u1_n153, u0_u9_u1_n154, u0_u9_u1_n155, 
       u0_u9_u1_n156, u0_u9_u1_n157, u0_u9_u1_n158, u0_u9_u1_n159, u0_u9_u1_n160, u0_u9_u1_n161, u0_u9_u1_n162, u0_u9_u1_n163, u0_u9_u1_n164, 
       u0_u9_u1_n165, u0_u9_u1_n166, u0_u9_u1_n167, u0_u9_u1_n168, u0_u9_u1_n169, u0_u9_u1_n170, u0_u9_u1_n171, u0_u9_u1_n172, u0_u9_u1_n173, 
       u0_u9_u1_n174, u0_u9_u1_n175, u0_u9_u1_n176, u0_u9_u1_n177, u0_u9_u1_n178, u0_u9_u1_n179, u0_u9_u1_n180, u0_u9_u1_n181, u0_u9_u1_n182, 
       u0_u9_u1_n183, u0_u9_u1_n184, u0_u9_u1_n185, u0_u9_u1_n186, u0_u9_u1_n187, u0_u9_u1_n188, u0_u9_u1_n95, u0_u9_u1_n96, u0_u9_u1_n97, 
       u0_u9_u1_n98, u0_u9_u1_n99, u0_u9_u2_n100, u0_u9_u2_n101, u0_u9_u2_n102, u0_u9_u2_n103, u0_u9_u2_n104, u0_u9_u2_n105, u0_u9_u2_n106, 
       u0_u9_u2_n107, u0_u9_u2_n108, u0_u9_u2_n109, u0_u9_u2_n110, u0_u9_u2_n111, u0_u9_u2_n112, u0_u9_u2_n113, u0_u9_u2_n114, u0_u9_u2_n115, 
       u0_u9_u2_n116, u0_u9_u2_n117, u0_u9_u2_n118, u0_u9_u2_n119, u0_u9_u2_n120, u0_u9_u2_n121, u0_u9_u2_n122, u0_u9_u2_n123, u0_u9_u2_n124, 
       u0_u9_u2_n125, u0_u9_u2_n126, u0_u9_u2_n127, u0_u9_u2_n128, u0_u9_u2_n129, u0_u9_u2_n130, u0_u9_u2_n131, u0_u9_u2_n132, u0_u9_u2_n133, 
       u0_u9_u2_n134, u0_u9_u2_n135, u0_u9_u2_n136, u0_u9_u2_n137, u0_u9_u2_n138, u0_u9_u2_n139, u0_u9_u2_n140, u0_u9_u2_n141, u0_u9_u2_n142, 
       u0_u9_u2_n143, u0_u9_u2_n144, u0_u9_u2_n145, u0_u9_u2_n146, u0_u9_u2_n147, u0_u9_u2_n148, u0_u9_u2_n149, u0_u9_u2_n150, u0_u9_u2_n151, 
       u0_u9_u2_n152, u0_u9_u2_n153, u0_u9_u2_n154, u0_u9_u2_n155, u0_u9_u2_n156, u0_u9_u2_n157, u0_u9_u2_n158, u0_u9_u2_n159, u0_u9_u2_n160, 
       u0_u9_u2_n161, u0_u9_u2_n162, u0_u9_u2_n163, u0_u9_u2_n164, u0_u9_u2_n165, u0_u9_u2_n166, u0_u9_u2_n167, u0_u9_u2_n168, u0_u9_u2_n169, 
       u0_u9_u2_n170, u0_u9_u2_n171, u0_u9_u2_n172, u0_u9_u2_n173, u0_u9_u2_n174, u0_u9_u2_n175, u0_u9_u2_n176, u0_u9_u2_n177, u0_u9_u2_n178, 
       u0_u9_u2_n179, u0_u9_u2_n180, u0_u9_u2_n181, u0_u9_u2_n182, u0_u9_u2_n183, u0_u9_u2_n184, u0_u9_u2_n185, u0_u9_u2_n186, u0_u9_u2_n187, 
       u0_u9_u2_n188, u0_u9_u2_n95, u0_u9_u2_n96, u0_u9_u2_n97, u0_u9_u2_n98, u0_u9_u2_n99, u0_u9_u6_n100, u0_u9_u6_n101, u0_u9_u6_n102, 
       u0_u9_u6_n103, u0_u9_u6_n104, u0_u9_u6_n105, u0_u9_u6_n106, u0_u9_u6_n107, u0_u9_u6_n108, u0_u9_u6_n109, u0_u9_u6_n110, u0_u9_u6_n111, 
       u0_u9_u6_n112, u0_u9_u6_n113, u0_u9_u6_n114, u0_u9_u6_n115, u0_u9_u6_n116, u0_u9_u6_n117, u0_u9_u6_n118, u0_u9_u6_n119, u0_u9_u6_n120, 
       u0_u9_u6_n121, u0_u9_u6_n122, u0_u9_u6_n123, u0_u9_u6_n124, u0_u9_u6_n125, u0_u9_u6_n126, u0_u9_u6_n127, u0_u9_u6_n128, u0_u9_u6_n129, 
       u0_u9_u6_n130, u0_u9_u6_n131, u0_u9_u6_n132, u0_u9_u6_n133, u0_u9_u6_n134, u0_u9_u6_n135, u0_u9_u6_n136, u0_u9_u6_n137, u0_u9_u6_n138, 
       u0_u9_u6_n139, u0_u9_u6_n140, u0_u9_u6_n141, u0_u9_u6_n142, u0_u9_u6_n143, u0_u9_u6_n144, u0_u9_u6_n145, u0_u9_u6_n146, u0_u9_u6_n147, 
       u0_u9_u6_n148, u0_u9_u6_n149, u0_u9_u6_n150, u0_u9_u6_n151, u0_u9_u6_n152, u0_u9_u6_n153, u0_u9_u6_n154, u0_u9_u6_n155, u0_u9_u6_n156, 
       u0_u9_u6_n157, u0_u9_u6_n158, u0_u9_u6_n159, u0_u9_u6_n160, u0_u9_u6_n161, u0_u9_u6_n162, u0_u9_u6_n163, u0_u9_u6_n164, u0_u9_u6_n165, 
       u0_u9_u6_n166, u0_u9_u6_n167, u0_u9_u6_n168, u0_u9_u6_n169, u0_u9_u6_n170, u0_u9_u6_n171, u0_u9_u6_n172, u0_u9_u6_n173, u0_u9_u6_n174, 
       u0_u9_u6_n88, u0_u9_u6_n89, u0_u9_u6_n90, u0_u9_u6_n91, u0_u9_u6_n92, u0_u9_u6_n93, u0_u9_u6_n94, u0_u9_u6_n95, u0_u9_u6_n96, 
       u0_u9_u6_n97, u0_u9_u6_n98, u0_u9_u6_n99, u0_uk_n1005, u0_uk_n1006, u0_uk_n1007, u0_uk_n1008, u0_uk_n1015, u0_uk_n1022, 
       u0_uk_n757, u0_uk_n758, u0_uk_n760, u0_uk_n864, u0_uk_n865, u0_uk_n866, u1_K11_19, u1_K11_20, u1_K11_21, 
       u1_K11_22, u1_K11_23, u1_K11_24, u1_K11_25, u1_K11_26, u1_K11_27, u1_K11_28, u1_K11_29, u1_K11_30, 
       u1_K11_43, u1_K11_44, u1_K11_45, u1_K11_46, u1_K11_47, u1_K11_48, u1_K12_10, u1_K12_11, u1_K12_12, 
       u1_K12_7, u1_K12_8, u1_K12_9, u1_K13_25, u1_K13_26, u1_K13_27, u1_K13_28, u1_K13_29, u1_K13_30, 
       u1_K13_31, u1_K13_32, u1_K13_33, u1_K13_34, u1_K13_35, u1_K13_36, u1_K14_37, u1_K14_38, u1_K14_39, 
       u1_K14_40, u1_K14_41, u1_K14_42, u1_K14_43, u1_K14_44, u1_K14_45, u1_K14_46, u1_K14_47, u1_K14_48, 
       u1_K7_25, u1_K7_26, u1_K7_27, u1_K7_28, u1_K7_29, u1_K7_30, u1_K8_37, u1_K8_38, u1_K8_39, 
       u1_K8_40, u1_K8_41, u1_K8_42, u1_K9_31, u1_K9_32, u1_K9_33, u1_K9_34, u1_K9_35, u1_K9_36, 
       u1_K9_37, u1_K9_38, u1_K9_39, u1_K9_40, u1_K9_41, u1_K9_42, u1_out10_1, u1_out10_10, u1_out10_14, 
       u1_out10_15, u1_out10_20, u1_out10_21, u1_out10_25, u1_out10_26, u1_out10_27, u1_out10_3, u1_out10_5, u1_out10_8, 
       u1_out11_13, u1_out11_18, u1_out11_2, u1_out11_28, u1_out12_11, u1_out12_14, u1_out12_19, u1_out12_25, u1_out12_29, 
       u1_out12_3, u1_out12_4, u1_out12_8, u1_out13_12, u1_out13_15, u1_out13_21, u1_out13_22, u1_out13_27, u1_out13_32, 
       u1_out13_5, u1_out13_7, u1_out6_14, u1_out6_25, u1_out6_3, u1_out6_8, u1_out7_12, u1_out7_22, u1_out7_32, 
       u1_out7_7, u1_out8_11, u1_out8_12, u1_out8_19, u1_out8_22, u1_out8_29, u1_out8_32, u1_out8_4, u1_out8_7, 
       u1_u10_X_19, u1_u10_X_20, u1_u10_X_21, u1_u10_X_22, u1_u10_X_23, u1_u10_X_24, u1_u10_X_25, u1_u10_X_26, u1_u10_X_27, 
       u1_u10_X_28, u1_u10_X_29, u1_u10_X_30, u1_u10_X_43, u1_u10_X_44, u1_u10_X_45, u1_u10_X_46, u1_u10_X_47, u1_u10_X_48, 
       u1_u10_u3_n100, u1_u10_u3_n101, u1_u10_u3_n102, u1_u10_u3_n103, u1_u10_u3_n104, u1_u10_u3_n105, u1_u10_u3_n106, u1_u10_u3_n107, u1_u10_u3_n108, 
       u1_u10_u3_n109, u1_u10_u3_n110, u1_u10_u3_n111, u1_u10_u3_n112, u1_u10_u3_n113, u1_u10_u3_n114, u1_u10_u3_n115, u1_u10_u3_n116, u1_u10_u3_n117, 
       u1_u10_u3_n118, u1_u10_u3_n119, u1_u10_u3_n120, u1_u10_u3_n121, u1_u10_u3_n122, u1_u10_u3_n123, u1_u10_u3_n124, u1_u10_u3_n125, u1_u10_u3_n126, 
       u1_u10_u3_n127, u1_u10_u3_n128, u1_u10_u3_n129, u1_u10_u3_n130, u1_u10_u3_n131, u1_u10_u3_n132, u1_u10_u3_n133, u1_u10_u3_n134, u1_u10_u3_n135, 
       u1_u10_u3_n136, u1_u10_u3_n137, u1_u10_u3_n138, u1_u10_u3_n139, u1_u10_u3_n140, u1_u10_u3_n141, u1_u10_u3_n142, u1_u10_u3_n143, u1_u10_u3_n144, 
       u1_u10_u3_n145, u1_u10_u3_n146, u1_u10_u3_n147, u1_u10_u3_n148, u1_u10_u3_n149, u1_u10_u3_n150, u1_u10_u3_n151, u1_u10_u3_n152, u1_u10_u3_n153, 
       u1_u10_u3_n154, u1_u10_u3_n155, u1_u10_u3_n156, u1_u10_u3_n157, u1_u10_u3_n158, u1_u10_u3_n159, u1_u10_u3_n160, u1_u10_u3_n161, u1_u10_u3_n162, 
       u1_u10_u3_n163, u1_u10_u3_n164, u1_u10_u3_n165, u1_u10_u3_n166, u1_u10_u3_n167, u1_u10_u3_n168, u1_u10_u3_n169, u1_u10_u3_n170, u1_u10_u3_n171, 
       u1_u10_u3_n172, u1_u10_u3_n173, u1_u10_u3_n174, u1_u10_u3_n175, u1_u10_u3_n176, u1_u10_u3_n177, u1_u10_u3_n178, u1_u10_u3_n179, u1_u10_u3_n180, 
       u1_u10_u3_n181, u1_u10_u3_n182, u1_u10_u3_n183, u1_u10_u3_n184, u1_u10_u3_n185, u1_u10_u3_n186, u1_u10_u3_n94, u1_u10_u3_n95, u1_u10_u3_n96, 
       u1_u10_u3_n97, u1_u10_u3_n98, u1_u10_u3_n99, u1_u10_u4_n100, u1_u10_u4_n101, u1_u10_u4_n102, u1_u10_u4_n103, u1_u10_u4_n104, u1_u10_u4_n105, 
       u1_u10_u4_n106, u1_u10_u4_n107, u1_u10_u4_n108, u1_u10_u4_n109, u1_u10_u4_n110, u1_u10_u4_n111, u1_u10_u4_n112, u1_u10_u4_n113, u1_u10_u4_n114, 
       u1_u10_u4_n115, u1_u10_u4_n116, u1_u10_u4_n117, u1_u10_u4_n118, u1_u10_u4_n119, u1_u10_u4_n120, u1_u10_u4_n121, u1_u10_u4_n122, u1_u10_u4_n123, 
       u1_u10_u4_n124, u1_u10_u4_n125, u1_u10_u4_n126, u1_u10_u4_n127, u1_u10_u4_n128, u1_u10_u4_n129, u1_u10_u4_n130, u1_u10_u4_n131, u1_u10_u4_n132, 
       u1_u10_u4_n133, u1_u10_u4_n134, u1_u10_u4_n135, u1_u10_u4_n136, u1_u10_u4_n137, u1_u10_u4_n138, u1_u10_u4_n139, u1_u10_u4_n140, u1_u10_u4_n141, 
       u1_u10_u4_n142, u1_u10_u4_n143, u1_u10_u4_n144, u1_u10_u4_n145, u1_u10_u4_n146, u1_u10_u4_n147, u1_u10_u4_n148, u1_u10_u4_n149, u1_u10_u4_n150, 
       u1_u10_u4_n151, u1_u10_u4_n152, u1_u10_u4_n153, u1_u10_u4_n154, u1_u10_u4_n155, u1_u10_u4_n156, u1_u10_u4_n157, u1_u10_u4_n158, u1_u10_u4_n159, 
       u1_u10_u4_n160, u1_u10_u4_n161, u1_u10_u4_n162, u1_u10_u4_n163, u1_u10_u4_n164, u1_u10_u4_n165, u1_u10_u4_n166, u1_u10_u4_n167, u1_u10_u4_n168, 
       u1_u10_u4_n169, u1_u10_u4_n170, u1_u10_u4_n171, u1_u10_u4_n172, u1_u10_u4_n173, u1_u10_u4_n174, u1_u10_u4_n175, u1_u10_u4_n176, u1_u10_u4_n177, 
       u1_u10_u4_n178, u1_u10_u4_n179, u1_u10_u4_n180, u1_u10_u4_n181, u1_u10_u4_n182, u1_u10_u4_n183, u1_u10_u4_n184, u1_u10_u4_n185, u1_u10_u4_n186, 
       u1_u10_u4_n94, u1_u10_u4_n95, u1_u10_u4_n96, u1_u10_u4_n97, u1_u10_u4_n98, u1_u10_u4_n99, u1_u10_u7_n100, u1_u10_u7_n101, u1_u10_u7_n102, 
       u1_u10_u7_n103, u1_u10_u7_n104, u1_u10_u7_n105, u1_u10_u7_n106, u1_u10_u7_n107, u1_u10_u7_n108, u1_u10_u7_n109, u1_u10_u7_n110, u1_u10_u7_n111, 
       u1_u10_u7_n112, u1_u10_u7_n113, u1_u10_u7_n114, u1_u10_u7_n115, u1_u10_u7_n116, u1_u10_u7_n117, u1_u10_u7_n118, u1_u10_u7_n119, u1_u10_u7_n120, 
       u1_u10_u7_n121, u1_u10_u7_n122, u1_u10_u7_n123, u1_u10_u7_n124, u1_u10_u7_n125, u1_u10_u7_n126, u1_u10_u7_n127, u1_u10_u7_n128, u1_u10_u7_n129, 
       u1_u10_u7_n130, u1_u10_u7_n131, u1_u10_u7_n132, u1_u10_u7_n133, u1_u10_u7_n134, u1_u10_u7_n135, u1_u10_u7_n136, u1_u10_u7_n137, u1_u10_u7_n138, 
       u1_u10_u7_n139, u1_u10_u7_n140, u1_u10_u7_n141, u1_u10_u7_n142, u1_u10_u7_n143, u1_u10_u7_n144, u1_u10_u7_n145, u1_u10_u7_n146, u1_u10_u7_n147, 
       u1_u10_u7_n148, u1_u10_u7_n149, u1_u10_u7_n150, u1_u10_u7_n151, u1_u10_u7_n152, u1_u10_u7_n153, u1_u10_u7_n154, u1_u10_u7_n155, u1_u10_u7_n156, 
       u1_u10_u7_n157, u1_u10_u7_n158, u1_u10_u7_n159, u1_u10_u7_n160, u1_u10_u7_n161, u1_u10_u7_n162, u1_u10_u7_n163, u1_u10_u7_n164, u1_u10_u7_n165, 
       u1_u10_u7_n166, u1_u10_u7_n167, u1_u10_u7_n168, u1_u10_u7_n169, u1_u10_u7_n170, u1_u10_u7_n171, u1_u10_u7_n172, u1_u10_u7_n173, u1_u10_u7_n174, 
       u1_u10_u7_n175, u1_u10_u7_n176, u1_u10_u7_n177, u1_u10_u7_n178, u1_u10_u7_n179, u1_u10_u7_n180, u1_u10_u7_n91, u1_u10_u7_n92, u1_u10_u7_n93, 
       u1_u10_u7_n94, u1_u10_u7_n95, u1_u10_u7_n96, u1_u10_u7_n97, u1_u10_u7_n98, u1_u10_u7_n99, u1_u11_X_10, u1_u11_X_11, u1_u11_X_12, 
       u1_u11_X_7, u1_u11_X_8, u1_u11_X_9, u1_u11_u1_n100, u1_u11_u1_n101, u1_u11_u1_n102, u1_u11_u1_n103, u1_u11_u1_n104, u1_u11_u1_n105, 
       u1_u11_u1_n106, u1_u11_u1_n107, u1_u11_u1_n108, u1_u11_u1_n109, u1_u11_u1_n110, u1_u11_u1_n111, u1_u11_u1_n112, u1_u11_u1_n113, u1_u11_u1_n114, 
       u1_u11_u1_n115, u1_u11_u1_n116, u1_u11_u1_n117, u1_u11_u1_n118, u1_u11_u1_n119, u1_u11_u1_n120, u1_u11_u1_n121, u1_u11_u1_n122, u1_u11_u1_n123, 
       u1_u11_u1_n124, u1_u11_u1_n125, u1_u11_u1_n126, u1_u11_u1_n127, u1_u11_u1_n128, u1_u11_u1_n129, u1_u11_u1_n130, u1_u11_u1_n131, u1_u11_u1_n132, 
       u1_u11_u1_n133, u1_u11_u1_n134, u1_u11_u1_n135, u1_u11_u1_n136, u1_u11_u1_n137, u1_u11_u1_n138, u1_u11_u1_n139, u1_u11_u1_n140, u1_u11_u1_n141, 
       u1_u11_u1_n142, u1_u11_u1_n143, u1_u11_u1_n144, u1_u11_u1_n145, u1_u11_u1_n146, u1_u11_u1_n147, u1_u11_u1_n148, u1_u11_u1_n149, u1_u11_u1_n150, 
       u1_u11_u1_n151, u1_u11_u1_n152, u1_u11_u1_n153, u1_u11_u1_n154, u1_u11_u1_n155, u1_u11_u1_n156, u1_u11_u1_n157, u1_u11_u1_n158, u1_u11_u1_n159, 
       u1_u11_u1_n160, u1_u11_u1_n161, u1_u11_u1_n162, u1_u11_u1_n163, u1_u11_u1_n164, u1_u11_u1_n165, u1_u11_u1_n166, u1_u11_u1_n167, u1_u11_u1_n168, 
       u1_u11_u1_n169, u1_u11_u1_n170, u1_u11_u1_n171, u1_u11_u1_n172, u1_u11_u1_n173, u1_u11_u1_n174, u1_u11_u1_n175, u1_u11_u1_n176, u1_u11_u1_n177, 
       u1_u11_u1_n178, u1_u11_u1_n179, u1_u11_u1_n180, u1_u11_u1_n181, u1_u11_u1_n182, u1_u11_u1_n183, u1_u11_u1_n184, u1_u11_u1_n185, u1_u11_u1_n186, 
       u1_u11_u1_n187, u1_u11_u1_n188, u1_u11_u1_n95, u1_u11_u1_n96, u1_u11_u1_n97, u1_u11_u1_n98, u1_u11_u1_n99, u1_u12_X_25, u1_u12_X_26, 
       u1_u12_X_27, u1_u12_X_28, u1_u12_X_29, u1_u12_X_30, u1_u12_X_31, u1_u12_X_32, u1_u12_X_33, u1_u12_X_34, u1_u12_X_35, 
       u1_u12_X_36, u1_u12_u4_n100, u1_u12_u4_n101, u1_u12_u4_n102, u1_u12_u4_n103, u1_u12_u4_n104, u1_u12_u4_n105, u1_u12_u4_n106, u1_u12_u4_n107, 
       u1_u12_u4_n108, u1_u12_u4_n109, u1_u12_u4_n110, u1_u12_u4_n111, u1_u12_u4_n112, u1_u12_u4_n113, u1_u12_u4_n114, u1_u12_u4_n115, u1_u12_u4_n116, 
       u1_u12_u4_n117, u1_u12_u4_n118, u1_u12_u4_n119, u1_u12_u4_n120, u1_u12_u4_n121, u1_u12_u4_n122, u1_u12_u4_n123, u1_u12_u4_n124, u1_u12_u4_n125, 
       u1_u12_u4_n126, u1_u12_u4_n127, u1_u12_u4_n128, u1_u12_u4_n129, u1_u12_u4_n130, u1_u12_u4_n131, u1_u12_u4_n132, u1_u12_u4_n133, u1_u12_u4_n134, 
       u1_u12_u4_n135, u1_u12_u4_n136, u1_u12_u4_n137, u1_u12_u4_n138, u1_u12_u4_n139, u1_u12_u4_n140, u1_u12_u4_n141, u1_u12_u4_n142, u1_u12_u4_n143, 
       u1_u12_u4_n144, u1_u12_u4_n145, u1_u12_u4_n146, u1_u12_u4_n147, u1_u12_u4_n148, u1_u12_u4_n149, u1_u12_u4_n150, u1_u12_u4_n151, u1_u12_u4_n152, 
       u1_u12_u4_n153, u1_u12_u4_n154, u1_u12_u4_n155, u1_u12_u4_n156, u1_u12_u4_n157, u1_u12_u4_n158, u1_u12_u4_n159, u1_u12_u4_n160, u1_u12_u4_n161, 
       u1_u12_u4_n162, u1_u12_u4_n163, u1_u12_u4_n164, u1_u12_u4_n165, u1_u12_u4_n166, u1_u12_u4_n167, u1_u12_u4_n168, u1_u12_u4_n169, u1_u12_u4_n170, 
       u1_u12_u4_n171, u1_u12_u4_n172, u1_u12_u4_n173, u1_u12_u4_n174, u1_u12_u4_n175, u1_u12_u4_n176, u1_u12_u4_n177, u1_u12_u4_n178, u1_u12_u4_n179, 
       u1_u12_u4_n180, u1_u12_u4_n181, u1_u12_u4_n182, u1_u12_u4_n183, u1_u12_u4_n184, u1_u12_u4_n185, u1_u12_u4_n186, u1_u12_u4_n94, u1_u12_u4_n95, 
       u1_u12_u4_n96, u1_u12_u4_n97, u1_u12_u4_n98, u1_u12_u4_n99, u1_u12_u5_n100, u1_u12_u5_n101, u1_u12_u5_n102, u1_u12_u5_n103, u1_u12_u5_n104, 
       u1_u12_u5_n105, u1_u12_u5_n106, u1_u12_u5_n107, u1_u12_u5_n108, u1_u12_u5_n109, u1_u12_u5_n110, u1_u12_u5_n111, u1_u12_u5_n112, u1_u12_u5_n113, 
       u1_u12_u5_n114, u1_u12_u5_n115, u1_u12_u5_n116, u1_u12_u5_n117, u1_u12_u5_n118, u1_u12_u5_n119, u1_u12_u5_n120, u1_u12_u5_n121, u1_u12_u5_n122, 
       u1_u12_u5_n123, u1_u12_u5_n124, u1_u12_u5_n125, u1_u12_u5_n126, u1_u12_u5_n127, u1_u12_u5_n128, u1_u12_u5_n129, u1_u12_u5_n130, u1_u12_u5_n131, 
       u1_u12_u5_n132, u1_u12_u5_n133, u1_u12_u5_n134, u1_u12_u5_n135, u1_u12_u5_n136, u1_u12_u5_n137, u1_u12_u5_n138, u1_u12_u5_n139, u1_u12_u5_n140, 
       u1_u12_u5_n141, u1_u12_u5_n142, u1_u12_u5_n143, u1_u12_u5_n144, u1_u12_u5_n145, u1_u12_u5_n146, u1_u12_u5_n147, u1_u12_u5_n148, u1_u12_u5_n149, 
       u1_u12_u5_n150, u1_u12_u5_n151, u1_u12_u5_n152, u1_u12_u5_n153, u1_u12_u5_n154, u1_u12_u5_n155, u1_u12_u5_n156, u1_u12_u5_n157, u1_u12_u5_n158, 
       u1_u12_u5_n159, u1_u12_u5_n160, u1_u12_u5_n161, u1_u12_u5_n162, u1_u12_u5_n163, u1_u12_u5_n164, u1_u12_u5_n165, u1_u12_u5_n166, u1_u12_u5_n167, 
       u1_u12_u5_n168, u1_u12_u5_n169, u1_u12_u5_n170, u1_u12_u5_n171, u1_u12_u5_n172, u1_u12_u5_n173, u1_u12_u5_n174, u1_u12_u5_n175, u1_u12_u5_n176, 
       u1_u12_u5_n177, u1_u12_u5_n178, u1_u12_u5_n179, u1_u12_u5_n180, u1_u12_u5_n181, u1_u12_u5_n182, u1_u12_u5_n183, u1_u12_u5_n184, u1_u12_u5_n185, 
       u1_u12_u5_n186, u1_u12_u5_n187, u1_u12_u5_n188, u1_u12_u5_n189, u1_u12_u5_n190, u1_u12_u5_n191, u1_u12_u5_n192, u1_u12_u5_n193, u1_u12_u5_n194, 
       u1_u12_u5_n195, u1_u12_u5_n196, u1_u12_u5_n99, u1_u13_X_37, u1_u13_X_38, u1_u13_X_39, u1_u13_X_40, u1_u13_X_41, u1_u13_X_42, 
       u1_u13_X_43, u1_u13_X_44, u1_u13_X_45, u1_u13_X_46, u1_u13_X_47, u1_u13_X_48, u1_u13_u6_n100, u1_u13_u6_n101, u1_u13_u6_n102, 
       u1_u13_u6_n103, u1_u13_u6_n104, u1_u13_u6_n105, u1_u13_u6_n106, u1_u13_u6_n107, u1_u13_u6_n108, u1_u13_u6_n109, u1_u13_u6_n110, u1_u13_u6_n111, 
       u1_u13_u6_n112, u1_u13_u6_n113, u1_u13_u6_n114, u1_u13_u6_n115, u1_u13_u6_n116, u1_u13_u6_n117, u1_u13_u6_n118, u1_u13_u6_n119, u1_u13_u6_n120, 
       u1_u13_u6_n121, u1_u13_u6_n122, u1_u13_u6_n123, u1_u13_u6_n124, u1_u13_u6_n125, u1_u13_u6_n126, u1_u13_u6_n127, u1_u13_u6_n128, u1_u13_u6_n129, 
       u1_u13_u6_n130, u1_u13_u6_n131, u1_u13_u6_n132, u1_u13_u6_n133, u1_u13_u6_n134, u1_u13_u6_n135, u1_u13_u6_n136, u1_u13_u6_n137, u1_u13_u6_n138, 
       u1_u13_u6_n139, u1_u13_u6_n140, u1_u13_u6_n141, u1_u13_u6_n142, u1_u13_u6_n143, u1_u13_u6_n144, u1_u13_u6_n145, u1_u13_u6_n146, u1_u13_u6_n147, 
       u1_u13_u6_n148, u1_u13_u6_n149, u1_u13_u6_n150, u1_u13_u6_n151, u1_u13_u6_n152, u1_u13_u6_n153, u1_u13_u6_n154, u1_u13_u6_n155, u1_u13_u6_n156, 
       u1_u13_u6_n157, u1_u13_u6_n158, u1_u13_u6_n159, u1_u13_u6_n160, u1_u13_u6_n161, u1_u13_u6_n162, u1_u13_u6_n163, u1_u13_u6_n164, u1_u13_u6_n165, 
       u1_u13_u6_n166, u1_u13_u6_n167, u1_u13_u6_n168, u1_u13_u6_n169, u1_u13_u6_n170, u1_u13_u6_n171, u1_u13_u6_n172, u1_u13_u6_n173, u1_u13_u6_n174, 
       u1_u13_u6_n88, u1_u13_u6_n89, u1_u13_u6_n90, u1_u13_u6_n91, u1_u13_u6_n92, u1_u13_u6_n93, u1_u13_u6_n94, u1_u13_u6_n95, u1_u13_u6_n96, 
       u1_u13_u6_n97, u1_u13_u6_n98, u1_u13_u6_n99, u1_u13_u7_n100, u1_u13_u7_n101, u1_u13_u7_n102, u1_u13_u7_n103, u1_u13_u7_n104, u1_u13_u7_n105, 
       u1_u13_u7_n106, u1_u13_u7_n107, u1_u13_u7_n108, u1_u13_u7_n109, u1_u13_u7_n110, u1_u13_u7_n111, u1_u13_u7_n112, u1_u13_u7_n113, u1_u13_u7_n114, 
       u1_u13_u7_n115, u1_u13_u7_n116, u1_u13_u7_n117, u1_u13_u7_n118, u1_u13_u7_n119, u1_u13_u7_n120, u1_u13_u7_n121, u1_u13_u7_n122, u1_u13_u7_n123, 
       u1_u13_u7_n124, u1_u13_u7_n125, u1_u13_u7_n126, u1_u13_u7_n127, u1_u13_u7_n128, u1_u13_u7_n129, u1_u13_u7_n130, u1_u13_u7_n131, u1_u13_u7_n132, 
       u1_u13_u7_n133, u1_u13_u7_n134, u1_u13_u7_n135, u1_u13_u7_n136, u1_u13_u7_n137, u1_u13_u7_n138, u1_u13_u7_n139, u1_u13_u7_n140, u1_u13_u7_n141, 
       u1_u13_u7_n142, u1_u13_u7_n143, u1_u13_u7_n144, u1_u13_u7_n145, u1_u13_u7_n146, u1_u13_u7_n147, u1_u13_u7_n148, u1_u13_u7_n149, u1_u13_u7_n150, 
       u1_u13_u7_n151, u1_u13_u7_n152, u1_u13_u7_n153, u1_u13_u7_n154, u1_u13_u7_n155, u1_u13_u7_n156, u1_u13_u7_n157, u1_u13_u7_n158, u1_u13_u7_n159, 
       u1_u13_u7_n160, u1_u13_u7_n161, u1_u13_u7_n162, u1_u13_u7_n163, u1_u13_u7_n164, u1_u13_u7_n165, u1_u13_u7_n166, u1_u13_u7_n167, u1_u13_u7_n168, 
       u1_u13_u7_n169, u1_u13_u7_n170, u1_u13_u7_n171, u1_u13_u7_n172, u1_u13_u7_n173, u1_u13_u7_n174, u1_u13_u7_n175, u1_u13_u7_n176, u1_u13_u7_n177, 
       u1_u13_u7_n178, u1_u13_u7_n179, u1_u13_u7_n180, u1_u13_u7_n91, u1_u13_u7_n92, u1_u13_u7_n93, u1_u13_u7_n94, u1_u13_u7_n95, u1_u13_u7_n96, 
       u1_u13_u7_n97, u1_u13_u7_n98, u1_u13_u7_n99, u1_u6_X_25, u1_u6_X_26, u1_u6_X_27, u1_u6_X_28, u1_u6_X_29, u1_u6_X_30, 
       u1_u6_u4_n100, u1_u6_u4_n101, u1_u6_u4_n102, u1_u6_u4_n103, u1_u6_u4_n104, u1_u6_u4_n105, u1_u6_u4_n106, u1_u6_u4_n107, u1_u6_u4_n108, 
       u1_u6_u4_n109, u1_u6_u4_n110, u1_u6_u4_n111, u1_u6_u4_n112, u1_u6_u4_n113, u1_u6_u4_n114, u1_u6_u4_n115, u1_u6_u4_n116, u1_u6_u4_n117, 
       u1_u6_u4_n118, u1_u6_u4_n119, u1_u6_u4_n120, u1_u6_u4_n121, u1_u6_u4_n122, u1_u6_u4_n123, u1_u6_u4_n124, u1_u6_u4_n125, u1_u6_u4_n126, 
       u1_u6_u4_n127, u1_u6_u4_n128, u1_u6_u4_n129, u1_u6_u4_n130, u1_u6_u4_n131, u1_u6_u4_n132, u1_u6_u4_n133, u1_u6_u4_n134, u1_u6_u4_n135, 
       u1_u6_u4_n136, u1_u6_u4_n137, u1_u6_u4_n138, u1_u6_u4_n139, u1_u6_u4_n140, u1_u6_u4_n141, u1_u6_u4_n142, u1_u6_u4_n143, u1_u6_u4_n144, 
       u1_u6_u4_n145, u1_u6_u4_n146, u1_u6_u4_n147, u1_u6_u4_n148, u1_u6_u4_n149, u1_u6_u4_n150, u1_u6_u4_n151, u1_u6_u4_n152, u1_u6_u4_n153, 
       u1_u6_u4_n154, u1_u6_u4_n155, u1_u6_u4_n156, u1_u6_u4_n157, u1_u6_u4_n158, u1_u6_u4_n159, u1_u6_u4_n160, u1_u6_u4_n161, u1_u6_u4_n162, 
       u1_u6_u4_n163, u1_u6_u4_n164, u1_u6_u4_n165, u1_u6_u4_n166, u1_u6_u4_n167, u1_u6_u4_n168, u1_u6_u4_n169, u1_u6_u4_n170, u1_u6_u4_n171, 
       u1_u6_u4_n172, u1_u6_u4_n173, u1_u6_u4_n174, u1_u6_u4_n175, u1_u6_u4_n176, u1_u6_u4_n177, u1_u6_u4_n178, u1_u6_u4_n179, u1_u6_u4_n180, 
       u1_u6_u4_n181, u1_u6_u4_n182, u1_u6_u4_n183, u1_u6_u4_n184, u1_u6_u4_n185, u1_u6_u4_n186, u1_u6_u4_n94, u1_u6_u4_n95, u1_u6_u4_n96, 
       u1_u6_u4_n97, u1_u6_u4_n98, u1_u6_u4_n99, u1_u7_X_37, u1_u7_X_38, u1_u7_X_39, u1_u7_X_40, u1_u7_X_41, u1_u7_X_42, 
       u1_u7_u6_n100, u1_u7_u6_n101, u1_u7_u6_n102, u1_u7_u6_n103, u1_u7_u6_n104, u1_u7_u6_n105, u1_u7_u6_n106, u1_u7_u6_n107, u1_u7_u6_n108, 
       u1_u7_u6_n109, u1_u7_u6_n110, u1_u7_u6_n111, u1_u7_u6_n112, u1_u7_u6_n113, u1_u7_u6_n114, u1_u7_u6_n115, u1_u7_u6_n116, u1_u7_u6_n117, 
       u1_u7_u6_n118, u1_u7_u6_n119, u1_u7_u6_n120, u1_u7_u6_n121, u1_u7_u6_n122, u1_u7_u6_n123, u1_u7_u6_n124, u1_u7_u6_n125, u1_u7_u6_n126, 
       u1_u7_u6_n127, u1_u7_u6_n128, u1_u7_u6_n129, u1_u7_u6_n130, u1_u7_u6_n131, u1_u7_u6_n132, u1_u7_u6_n133, u1_u7_u6_n134, u1_u7_u6_n135, 
       u1_u7_u6_n136, u1_u7_u6_n137, u1_u7_u6_n138, u1_u7_u6_n139, u1_u7_u6_n140, u1_u7_u6_n141, u1_u7_u6_n142, u1_u7_u6_n143, u1_u7_u6_n144, 
       u1_u7_u6_n145, u1_u7_u6_n146, u1_u7_u6_n147, u1_u7_u6_n148, u1_u7_u6_n149, u1_u7_u6_n150, u1_u7_u6_n151, u1_u7_u6_n152, u1_u7_u6_n153, 
       u1_u7_u6_n154, u1_u7_u6_n155, u1_u7_u6_n156, u1_u7_u6_n157, u1_u7_u6_n158, u1_u7_u6_n159, u1_u7_u6_n160, u1_u7_u6_n161, u1_u7_u6_n162, 
       u1_u7_u6_n163, u1_u7_u6_n164, u1_u7_u6_n165, u1_u7_u6_n166, u1_u7_u6_n167, u1_u7_u6_n168, u1_u7_u6_n169, u1_u7_u6_n170, u1_u7_u6_n171, 
       u1_u7_u6_n172, u1_u7_u6_n173, u1_u7_u6_n174, u1_u7_u6_n88, u1_u7_u6_n89, u1_u7_u6_n90, u1_u7_u6_n91, u1_u7_u6_n92, u1_u7_u6_n93, 
       u1_u7_u6_n94, u1_u7_u6_n95, u1_u7_u6_n96, u1_u7_u6_n97, u1_u7_u6_n98, u1_u7_u6_n99, u1_u8_X_31, u1_u8_X_32, u1_u8_X_33, 
       u1_u8_X_34, u1_u8_X_35, u1_u8_X_36, u1_u8_X_37, u1_u8_X_38, u1_u8_X_39, u1_u8_X_40, u1_u8_X_41, u1_u8_X_42, 
       u1_u8_u5_n100, u1_u8_u5_n101, u1_u8_u5_n102, u1_u8_u5_n103, u1_u8_u5_n104, u1_u8_u5_n105, u1_u8_u5_n106, u1_u8_u5_n107, u1_u8_u5_n108, 
       u1_u8_u5_n109, u1_u8_u5_n110, u1_u8_u5_n111, u1_u8_u5_n112, u1_u8_u5_n113, u1_u8_u5_n114, u1_u8_u5_n115, u1_u8_u5_n116, u1_u8_u5_n117, 
       u1_u8_u5_n118, u1_u8_u5_n119, u1_u8_u5_n120, u1_u8_u5_n121, u1_u8_u5_n122, u1_u8_u5_n123, u1_u8_u5_n124, u1_u8_u5_n125, u1_u8_u5_n126, 
       u1_u8_u5_n127, u1_u8_u5_n128, u1_u8_u5_n129, u1_u8_u5_n130, u1_u8_u5_n131, u1_u8_u5_n132, u1_u8_u5_n133, u1_u8_u5_n134, u1_u8_u5_n135, 
       u1_u8_u5_n136, u1_u8_u5_n137, u1_u8_u5_n138, u1_u8_u5_n139, u1_u8_u5_n140, u1_u8_u5_n141, u1_u8_u5_n142, u1_u8_u5_n143, u1_u8_u5_n144, 
       u1_u8_u5_n145, u1_u8_u5_n146, u1_u8_u5_n147, u1_u8_u5_n148, u1_u8_u5_n149, u1_u8_u5_n150, u1_u8_u5_n151, u1_u8_u5_n152, u1_u8_u5_n153, 
       u1_u8_u5_n154, u1_u8_u5_n155, u1_u8_u5_n156, u1_u8_u5_n157, u1_u8_u5_n158, u1_u8_u5_n159, u1_u8_u5_n160, u1_u8_u5_n161, u1_u8_u5_n162, 
       u1_u8_u5_n163, u1_u8_u5_n164, u1_u8_u5_n165, u1_u8_u5_n166, u1_u8_u5_n167, u1_u8_u5_n168, u1_u8_u5_n169, u1_u8_u5_n170, u1_u8_u5_n171, 
       u1_u8_u5_n172, u1_u8_u5_n173, u1_u8_u5_n174, u1_u8_u5_n175, u1_u8_u5_n176, u1_u8_u5_n177, u1_u8_u5_n178, u1_u8_u5_n179, u1_u8_u5_n180, 
       u1_u8_u5_n181, u1_u8_u5_n182, u1_u8_u5_n183, u1_u8_u5_n184, u1_u8_u5_n185, u1_u8_u5_n186, u1_u8_u5_n187, u1_u8_u5_n188, u1_u8_u5_n189, 
       u1_u8_u5_n190, u1_u8_u5_n191, u1_u8_u5_n192, u1_u8_u5_n193, u1_u8_u5_n194, u1_u8_u5_n195, u1_u8_u5_n196, u1_u8_u5_n99, u1_u8_u6_n100, 
       u1_u8_u6_n101, u1_u8_u6_n102, u1_u8_u6_n103, u1_u8_u6_n104, u1_u8_u6_n105, u1_u8_u6_n106, u1_u8_u6_n107, u1_u8_u6_n108, u1_u8_u6_n109, 
       u1_u8_u6_n110, u1_u8_u6_n111, u1_u8_u6_n112, u1_u8_u6_n113, u1_u8_u6_n114, u1_u8_u6_n115, u1_u8_u6_n116, u1_u8_u6_n117, u1_u8_u6_n118, 
       u1_u8_u6_n119, u1_u8_u6_n120, u1_u8_u6_n121, u1_u8_u6_n122, u1_u8_u6_n123, u1_u8_u6_n124, u1_u8_u6_n125, u1_u8_u6_n126, u1_u8_u6_n127, 
       u1_u8_u6_n128, u1_u8_u6_n129, u1_u8_u6_n130, u1_u8_u6_n131, u1_u8_u6_n132, u1_u8_u6_n133, u1_u8_u6_n134, u1_u8_u6_n135, u1_u8_u6_n136, 
       u1_u8_u6_n137, u1_u8_u6_n138, u1_u8_u6_n139, u1_u8_u6_n140, u1_u8_u6_n141, u1_u8_u6_n142, u1_u8_u6_n143, u1_u8_u6_n144, u1_u8_u6_n145, 
       u1_u8_u6_n146, u1_u8_u6_n147, u1_u8_u6_n148, u1_u8_u6_n149, u1_u8_u6_n150, u1_u8_u6_n151, u1_u8_u6_n152, u1_u8_u6_n153, u1_u8_u6_n154, 
       u1_u8_u6_n155, u1_u8_u6_n156, u1_u8_u6_n157, u1_u8_u6_n158, u1_u8_u6_n159, u1_u8_u6_n160, u1_u8_u6_n161, u1_u8_u6_n162, u1_u8_u6_n163, 
       u1_u8_u6_n164, u1_u8_u6_n165, u1_u8_u6_n166, u1_u8_u6_n167, u1_u8_u6_n168, u1_u8_u6_n169, u1_u8_u6_n170, u1_u8_u6_n171, u1_u8_u6_n172, 
       u1_u8_u6_n173, u1_u8_u6_n174, u1_u8_u6_n88, u1_u8_u6_n89, u1_u8_u6_n90, u1_u8_u6_n91, u1_u8_u6_n92, u1_u8_u6_n93, u1_u8_u6_n94, 
       u1_u8_u6_n95, u1_u8_u6_n96, u1_u8_u6_n97, u1_u8_u6_n98, u1_u8_u6_n99, u1_uk_n1114, u1_uk_n1115, u1_uk_n1138, u1_uk_n1139, 
       u1_uk_n1141, u1_uk_n1142, u1_uk_n1162, u1_uk_n1163, u1_uk_n1164, u1_uk_n1165, u1_uk_n1166, u1_uk_n1167, u1_uk_n386, 
       u1_uk_n391, u1_uk_n395, u1_uk_n407, u1_uk_n408, u1_uk_n409, u1_uk_n415, u1_uk_n421, u1_uk_n468, u1_uk_n472, 
       u1_uk_n503, u1_uk_n665, u1_uk_n694, u1_uk_n695, u1_uk_n717, u1_uk_n958, u1_uk_n959, u1_uk_n960, u1_uk_n961, 
       u2_K10_19, u2_K10_20, u2_K10_21, u2_K10_22, u2_K10_23, u2_K10_24, u2_out9_1, u2_out9_10, u2_out9_20, 
       u2_out9_26, u2_u9_X_19, u2_u9_X_20, u2_u9_X_21, u2_u9_X_22, u2_u9_X_23, u2_u9_X_24, u2_u9_u3_n100, u2_u9_u3_n101, 
       u2_u9_u3_n102, u2_u9_u3_n103, u2_u9_u3_n104, u2_u9_u3_n105, u2_u9_u3_n106, u2_u9_u3_n107, u2_u9_u3_n108, u2_u9_u3_n109, u2_u9_u3_n110, 
       u2_u9_u3_n111, u2_u9_u3_n112, u2_u9_u3_n113, u2_u9_u3_n114, u2_u9_u3_n115, u2_u9_u3_n116, u2_u9_u3_n117, u2_u9_u3_n118, u2_u9_u3_n119, 
       u2_u9_u3_n120, u2_u9_u3_n121, u2_u9_u3_n122, u2_u9_u3_n123, u2_u9_u3_n124, u2_u9_u3_n125, u2_u9_u3_n126, u2_u9_u3_n127, u2_u9_u3_n128, 
       u2_u9_u3_n129, u2_u9_u3_n130, u2_u9_u3_n131, u2_u9_u3_n132, u2_u9_u3_n133, u2_u9_u3_n134, u2_u9_u3_n135, u2_u9_u3_n136, u2_u9_u3_n137, 
       u2_u9_u3_n138, u2_u9_u3_n139, u2_u9_u3_n140, u2_u9_u3_n141, u2_u9_u3_n142, u2_u9_u3_n143, u2_u9_u3_n144, u2_u9_u3_n145, u2_u9_u3_n146, 
       u2_u9_u3_n147, u2_u9_u3_n148, u2_u9_u3_n149, u2_u9_u3_n150, u2_u9_u3_n151, u2_u9_u3_n152, u2_u9_u3_n153, u2_u9_u3_n154, u2_u9_u3_n155, 
       u2_u9_u3_n156, u2_u9_u3_n157, u2_u9_u3_n158, u2_u9_u3_n159, u2_u9_u3_n160, u2_u9_u3_n161, u2_u9_u3_n162, u2_u9_u3_n163, u2_u9_u3_n164, 
       u2_u9_u3_n165, u2_u9_u3_n166, u2_u9_u3_n167, u2_u9_u3_n168, u2_u9_u3_n169, u2_u9_u3_n170, u2_u9_u3_n171, u2_u9_u3_n172, u2_u9_u3_n173, 
       u2_u9_u3_n174, u2_u9_u3_n175, u2_u9_u3_n176, u2_u9_u3_n177, u2_u9_u3_n178, u2_u9_u3_n179, u2_u9_u3_n180, u2_u9_u3_n181, u2_u9_u3_n182, 
       u2_u9_u3_n183, u2_u9_u3_n184, u2_u9_u3_n185, u2_u9_u3_n186, u2_u9_u3_n94, u2_u9_u3_n95, u2_u9_u3_n96, u2_u9_u3_n97, u2_u9_u3_n98, 
       u2_u9_u3_n99, u2_uk_n252, u2_uk_n271,  u2_uk_n277;
  XOR2_X1 u0_U136 (.B( u0_L0_10 ) , .Z( u0_N41 ) , .A( u0_out1_10 ) );
  XOR2_X1 u0_U181 (.B( u0_L0_6 ) , .Z( u0_N37 ) , .A( u0_out1_6 ) );
  XOR2_X1 u0_U236 (.B( u0_L0_1 ) , .Z( u0_N32 ) , .A( u0_out1_1 ) );
  XOR2_X1 u0_U237 (.B( u0_L8_32 ) , .Z( u0_N319 ) , .A( u0_out9_32 ) );
  XOR2_X1 u0_U238 (.B( u0_L8_31 ) , .Z( u0_N318 ) , .A( u0_out9_31 ) );
  XOR2_X1 u0_U239 (.B( u0_L8_30 ) , .Z( u0_N317 ) , .A( u0_out9_30 ) );
  XOR2_X1 u0_U241 (.B( u0_L8_28 ) , .Z( u0_N315 ) , .A( u0_out9_28 ) );
  XOR2_X1 u0_U245 (.B( u0_L8_24 ) , .Z( u0_N311 ) , .A( u0_out9_24 ) );
  XOR2_X1 u0_U246 (.B( u0_L8_23 ) , .Z( u0_N310 ) , .A( u0_out9_23 ) );
  XOR2_X1 u0_U248 (.B( u0_L8_22 ) , .Z( u0_N309 ) , .A( u0_out9_22 ) );
  XOR2_X1 u0_U252 (.B( u0_L8_18 ) , .Z( u0_N305 ) , .A( u0_out9_18 ) );
  XOR2_X1 u0_U253 (.B( u0_L8_17 ) , .Z( u0_N304 ) , .A( u0_out9_17 ) );
  XOR2_X1 u0_U254 (.B( u0_L8_16 ) , .Z( u0_N303 ) , .A( u0_out9_16 ) );
  XOR2_X1 u0_U257 (.B( u0_L8_13 ) , .Z( u0_N300 ) , .A( u0_out9_13 ) );
  XOR2_X1 u0_U260 (.B( u0_L8_12 ) , .Z( u0_N299 ) , .A( u0_out9_12 ) );
  XOR2_X1 u0_U263 (.B( u0_L8_9 ) , .Z( u0_N296 ) , .A( u0_out9_9 ) );
  XOR2_X1 u0_U265 (.B( u0_L8_7 ) , .Z( u0_N294 ) , .A( u0_out9_7 ) );
  XOR2_X1 u0_U266 (.B( u0_L8_6 ) , .Z( u0_N293 ) , .A( u0_out9_6 ) );
  XOR2_X1 u0_U271 (.B( u0_L8_2 ) , .Z( u0_N289 ) , .A( u0_out9_2 ) );
  XOR2_X1 u0_U310 (.B( u0_L6_30 ) , .Z( u0_N253 ) , .A( u0_out7_30 ) );
  XOR2_X1 u0_U315 (.B( u0_L6_26 ) , .Z( u0_N249 ) , .A( u0_out7_26 ) );
  XOR2_X1 u0_U317 (.B( u0_L6_24 ) , .Z( u0_N247 ) , .A( u0_out7_24 ) );
  XOR2_X1 u0_U321 (.B( u0_L6_20 ) , .Z( u0_N243 ) , .A( u0_out7_20 ) );
  XOR2_X1 u0_U326 (.B( u0_L6_16 ) , .Z( u0_N239 ) , .A( u0_out7_16 ) );
  XOR2_X1 u0_U332 (.B( u0_L6_10 ) , .Z( u0_N233 ) , .A( u0_out7_10 ) );
  XOR2_X1 u0_U337 (.B( u0_L6_6 ) , .Z( u0_N229 ) , .A( u0_out7_6 ) );
  XOR2_X1 u0_U342 (.B( u0_L6_1 ) , .Z( u0_N224 ) , .A( u0_out7_1 ) );
  XOR2_X1 u0_U44 (.B( u0_L0_30 ) , .Z( u0_N61 ) , .A( u0_out1_30 ) );
  XOR2_X1 u0_U49 (.B( u0_L0_26 ) , .Z( u0_N57 ) , .A( u0_out1_26 ) );
  XOR2_X1 u0_U51 (.B( u0_L0_24 ) , .Z( u0_N55 ) , .A( u0_out1_24 ) );
  XOR2_X1 u0_U55 (.B( u0_L0_20 ) , .Z( u0_N51 ) , .A( u0_out1_20 ) );
  XOR2_X1 u0_U70 (.B( u0_L0_16 ) , .Z( u0_N47 ) , .A( u0_out1_16 ) );
  XOR2_X1 u0_u1_U33 (.B( u0_K2_24 ) , .A( u0_R0_17 ) , .Z( u0_u1_X_24 ) );
  XOR2_X1 u0_u1_U34 (.B( u0_K2_23 ) , .A( u0_R0_16 ) , .Z( u0_u1_X_23 ) );
  XOR2_X1 u0_u1_U35 (.B( u0_K2_22 ) , .A( u0_R0_15 ) , .Z( u0_u1_X_22 ) );
  XOR2_X1 u0_u1_U36 (.B( u0_K2_21 ) , .A( u0_R0_14 ) , .Z( u0_u1_X_21 ) );
  XOR2_X1 u0_u1_U37 (.B( u0_K2_20 ) , .A( u0_R0_13 ) , .Z( u0_u1_X_20 ) );
  XOR2_X1 u0_u1_U39 (.B( u0_K2_19 ) , .A( u0_R0_12 ) , .Z( u0_u1_X_19 ) );
  XOR2_X1 u0_u1_U40 (.B( u0_K2_18 ) , .A( u0_R0_13 ) , .Z( u0_u1_X_18 ) );
  XOR2_X1 u0_u1_U41 (.B( u0_K2_17 ) , .A( u0_R0_12 ) , .Z( u0_u1_X_17 ) );
  XOR2_X1 u0_u1_U42 (.B( u0_K2_16 ) , .A( u0_R0_11 ) , .Z( u0_u1_X_16 ) );
  XOR2_X1 u0_u1_U43 (.B( u0_K2_15 ) , .A( u0_R0_10 ) , .Z( u0_u1_X_15 ) );
  XOR2_X1 u0_u1_U44 (.B( u0_K2_14 ) , .A( u0_R0_9 ) , .Z( u0_u1_X_14 ) );
  XOR2_X1 u0_u1_U45 (.B( u0_K2_13 ) , .A( u0_R0_8 ) , .Z( u0_u1_X_13 ) );
  OAI22_X1 u0_u1_u2_U10 (.ZN( u0_u1_u2_n109 ) , .A2( u0_u1_u2_n113 ) , .B2( u0_u1_u2_n133 ) , .B1( u0_u1_u2_n167 ) , .A1( u0_u1_u2_n168 ) );
  NAND3_X1 u0_u1_u2_U100 (.A2( u0_u1_u2_n100 ) , .A1( u0_u1_u2_n104 ) , .A3( u0_u1_u2_n138 ) , .ZN( u0_u1_u2_n98 ) );
  OAI22_X1 u0_u1_u2_U11 (.B1( u0_u1_u2_n151 ) , .A2( u0_u1_u2_n152 ) , .A1( u0_u1_u2_n153 ) , .ZN( u0_u1_u2_n160 ) , .B2( u0_u1_u2_n168 ) );
  NOR3_X1 u0_u1_u2_U12 (.A1( u0_u1_u2_n150 ) , .ZN( u0_u1_u2_n151 ) , .A3( u0_u1_u2_n175 ) , .A2( u0_u1_u2_n188 ) );
  AOI21_X1 u0_u1_u2_U13 (.ZN( u0_u1_u2_n144 ) , .B2( u0_u1_u2_n155 ) , .A( u0_u1_u2_n172 ) , .B1( u0_u1_u2_n185 ) );
  AOI21_X1 u0_u1_u2_U14 (.B2( u0_u1_u2_n143 ) , .ZN( u0_u1_u2_n145 ) , .B1( u0_u1_u2_n152 ) , .A( u0_u1_u2_n171 ) );
  AOI21_X1 u0_u1_u2_U15 (.B2( u0_u1_u2_n120 ) , .B1( u0_u1_u2_n121 ) , .ZN( u0_u1_u2_n126 ) , .A( u0_u1_u2_n167 ) );
  INV_X1 u0_u1_u2_U16 (.A( u0_u1_u2_n156 ) , .ZN( u0_u1_u2_n171 ) );
  INV_X1 u0_u1_u2_U17 (.A( u0_u1_u2_n120 ) , .ZN( u0_u1_u2_n188 ) );
  NAND2_X1 u0_u1_u2_U18 (.A2( u0_u1_u2_n122 ) , .ZN( u0_u1_u2_n150 ) , .A1( u0_u1_u2_n152 ) );
  INV_X1 u0_u1_u2_U19 (.A( u0_u1_u2_n153 ) , .ZN( u0_u1_u2_n170 ) );
  INV_X1 u0_u1_u2_U20 (.A( u0_u1_u2_n137 ) , .ZN( u0_u1_u2_n173 ) );
  NAND2_X1 u0_u1_u2_U21 (.A1( u0_u1_u2_n132 ) , .A2( u0_u1_u2_n139 ) , .ZN( u0_u1_u2_n157 ) );
  INV_X1 u0_u1_u2_U22 (.A( u0_u1_u2_n113 ) , .ZN( u0_u1_u2_n178 ) );
  INV_X1 u0_u1_u2_U23 (.A( u0_u1_u2_n139 ) , .ZN( u0_u1_u2_n175 ) );
  INV_X1 u0_u1_u2_U24 (.A( u0_u1_u2_n155 ) , .ZN( u0_u1_u2_n181 ) );
  INV_X1 u0_u1_u2_U25 (.A( u0_u1_u2_n119 ) , .ZN( u0_u1_u2_n177 ) );
  INV_X1 u0_u1_u2_U26 (.A( u0_u1_u2_n116 ) , .ZN( u0_u1_u2_n180 ) );
  INV_X1 u0_u1_u2_U27 (.A( u0_u1_u2_n131 ) , .ZN( u0_u1_u2_n179 ) );
  INV_X1 u0_u1_u2_U28 (.A( u0_u1_u2_n154 ) , .ZN( u0_u1_u2_n176 ) );
  NAND2_X1 u0_u1_u2_U29 (.A2( u0_u1_u2_n116 ) , .A1( u0_u1_u2_n117 ) , .ZN( u0_u1_u2_n118 ) );
  NOR2_X1 u0_u1_u2_U3 (.ZN( u0_u1_u2_n121 ) , .A2( u0_u1_u2_n177 ) , .A1( u0_u1_u2_n180 ) );
  INV_X1 u0_u1_u2_U30 (.A( u0_u1_u2_n132 ) , .ZN( u0_u1_u2_n182 ) );
  INV_X1 u0_u1_u2_U31 (.A( u0_u1_u2_n158 ) , .ZN( u0_u1_u2_n183 ) );
  OAI21_X1 u0_u1_u2_U32 (.A( u0_u1_u2_n156 ) , .B1( u0_u1_u2_n157 ) , .ZN( u0_u1_u2_n158 ) , .B2( u0_u1_u2_n179 ) );
  NOR2_X1 u0_u1_u2_U33 (.ZN( u0_u1_u2_n156 ) , .A1( u0_u1_u2_n166 ) , .A2( u0_u1_u2_n169 ) );
  NOR2_X1 u0_u1_u2_U34 (.A2( u0_u1_u2_n114 ) , .ZN( u0_u1_u2_n137 ) , .A1( u0_u1_u2_n140 ) );
  NOR2_X1 u0_u1_u2_U35 (.A2( u0_u1_u2_n138 ) , .ZN( u0_u1_u2_n153 ) , .A1( u0_u1_u2_n156 ) );
  AOI211_X1 u0_u1_u2_U36 (.ZN( u0_u1_u2_n130 ) , .C1( u0_u1_u2_n138 ) , .C2( u0_u1_u2_n179 ) , .B( u0_u1_u2_n96 ) , .A( u0_u1_u2_n97 ) );
  OAI22_X1 u0_u1_u2_U37 (.B1( u0_u1_u2_n133 ) , .A2( u0_u1_u2_n137 ) , .A1( u0_u1_u2_n152 ) , .B2( u0_u1_u2_n168 ) , .ZN( u0_u1_u2_n97 ) );
  OAI221_X1 u0_u1_u2_U38 (.B1( u0_u1_u2_n113 ) , .C1( u0_u1_u2_n132 ) , .A( u0_u1_u2_n149 ) , .B2( u0_u1_u2_n171 ) , .C2( u0_u1_u2_n172 ) , .ZN( u0_u1_u2_n96 ) );
  OAI221_X1 u0_u1_u2_U39 (.A( u0_u1_u2_n115 ) , .C2( u0_u1_u2_n123 ) , .B2( u0_u1_u2_n143 ) , .B1( u0_u1_u2_n153 ) , .ZN( u0_u1_u2_n163 ) , .C1( u0_u1_u2_n168 ) );
  INV_X1 u0_u1_u2_U4 (.A( u0_u1_u2_n134 ) , .ZN( u0_u1_u2_n185 ) );
  OAI21_X1 u0_u1_u2_U40 (.A( u0_u1_u2_n114 ) , .ZN( u0_u1_u2_n115 ) , .B1( u0_u1_u2_n176 ) , .B2( u0_u1_u2_n178 ) );
  OAI221_X1 u0_u1_u2_U41 (.A( u0_u1_u2_n135 ) , .B2( u0_u1_u2_n136 ) , .B1( u0_u1_u2_n137 ) , .ZN( u0_u1_u2_n162 ) , .C2( u0_u1_u2_n167 ) , .C1( u0_u1_u2_n185 ) );
  AND3_X1 u0_u1_u2_U42 (.A3( u0_u1_u2_n131 ) , .A2( u0_u1_u2_n132 ) , .A1( u0_u1_u2_n133 ) , .ZN( u0_u1_u2_n136 ) );
  AOI22_X1 u0_u1_u2_U43 (.ZN( u0_u1_u2_n135 ) , .B1( u0_u1_u2_n140 ) , .A1( u0_u1_u2_n156 ) , .B2( u0_u1_u2_n180 ) , .A2( u0_u1_u2_n188 ) );
  AOI21_X1 u0_u1_u2_U44 (.ZN( u0_u1_u2_n149 ) , .B1( u0_u1_u2_n173 ) , .B2( u0_u1_u2_n188 ) , .A( u0_u1_u2_n95 ) );
  AND3_X1 u0_u1_u2_U45 (.A2( u0_u1_u2_n100 ) , .A1( u0_u1_u2_n104 ) , .A3( u0_u1_u2_n156 ) , .ZN( u0_u1_u2_n95 ) );
  OAI21_X1 u0_u1_u2_U46 (.A( u0_u1_u2_n101 ) , .B2( u0_u1_u2_n121 ) , .B1( u0_u1_u2_n153 ) , .ZN( u0_u1_u2_n164 ) );
  NAND2_X1 u0_u1_u2_U47 (.A2( u0_u1_u2_n100 ) , .A1( u0_u1_u2_n107 ) , .ZN( u0_u1_u2_n155 ) );
  NAND2_X1 u0_u1_u2_U48 (.A2( u0_u1_u2_n105 ) , .A1( u0_u1_u2_n108 ) , .ZN( u0_u1_u2_n143 ) );
  NAND2_X1 u0_u1_u2_U49 (.A1( u0_u1_u2_n104 ) , .A2( u0_u1_u2_n106 ) , .ZN( u0_u1_u2_n152 ) );
  INV_X1 u0_u1_u2_U5 (.A( u0_u1_u2_n150 ) , .ZN( u0_u1_u2_n184 ) );
  NAND2_X1 u0_u1_u2_U50 (.A1( u0_u1_u2_n100 ) , .A2( u0_u1_u2_n105 ) , .ZN( u0_u1_u2_n132 ) );
  INV_X1 u0_u1_u2_U51 (.A( u0_u1_u2_n140 ) , .ZN( u0_u1_u2_n168 ) );
  INV_X1 u0_u1_u2_U52 (.A( u0_u1_u2_n138 ) , .ZN( u0_u1_u2_n167 ) );
  OAI21_X1 u0_u1_u2_U53 (.A( u0_u1_u2_n141 ) , .B2( u0_u1_u2_n142 ) , .ZN( u0_u1_u2_n146 ) , .B1( u0_u1_u2_n153 ) );
  OAI21_X1 u0_u1_u2_U54 (.A( u0_u1_u2_n140 ) , .ZN( u0_u1_u2_n141 ) , .B1( u0_u1_u2_n176 ) , .B2( u0_u1_u2_n177 ) );
  NOR3_X1 u0_u1_u2_U55 (.ZN( u0_u1_u2_n142 ) , .A3( u0_u1_u2_n175 ) , .A2( u0_u1_u2_n178 ) , .A1( u0_u1_u2_n181 ) );
  NAND2_X1 u0_u1_u2_U56 (.A1( u0_u1_u2_n102 ) , .A2( u0_u1_u2_n106 ) , .ZN( u0_u1_u2_n113 ) );
  NAND2_X1 u0_u1_u2_U57 (.A1( u0_u1_u2_n106 ) , .A2( u0_u1_u2_n107 ) , .ZN( u0_u1_u2_n131 ) );
  NAND2_X1 u0_u1_u2_U58 (.A1( u0_u1_u2_n103 ) , .A2( u0_u1_u2_n107 ) , .ZN( u0_u1_u2_n139 ) );
  NAND2_X1 u0_u1_u2_U59 (.A1( u0_u1_u2_n103 ) , .A2( u0_u1_u2_n105 ) , .ZN( u0_u1_u2_n133 ) );
  NOR4_X1 u0_u1_u2_U6 (.A4( u0_u1_u2_n124 ) , .A3( u0_u1_u2_n125 ) , .A2( u0_u1_u2_n126 ) , .A1( u0_u1_u2_n127 ) , .ZN( u0_u1_u2_n128 ) );
  NAND2_X1 u0_u1_u2_U60 (.A1( u0_u1_u2_n102 ) , .A2( u0_u1_u2_n103 ) , .ZN( u0_u1_u2_n154 ) );
  NAND2_X1 u0_u1_u2_U61 (.A2( u0_u1_u2_n103 ) , .A1( u0_u1_u2_n104 ) , .ZN( u0_u1_u2_n119 ) );
  NAND2_X1 u0_u1_u2_U62 (.A2( u0_u1_u2_n107 ) , .A1( u0_u1_u2_n108 ) , .ZN( u0_u1_u2_n123 ) );
  NAND2_X1 u0_u1_u2_U63 (.A1( u0_u1_u2_n104 ) , .A2( u0_u1_u2_n108 ) , .ZN( u0_u1_u2_n122 ) );
  INV_X1 u0_u1_u2_U64 (.A( u0_u1_u2_n114 ) , .ZN( u0_u1_u2_n172 ) );
  NAND2_X1 u0_u1_u2_U65 (.A2( u0_u1_u2_n100 ) , .A1( u0_u1_u2_n102 ) , .ZN( u0_u1_u2_n116 ) );
  NAND2_X1 u0_u1_u2_U66 (.A1( u0_u1_u2_n102 ) , .A2( u0_u1_u2_n108 ) , .ZN( u0_u1_u2_n120 ) );
  NAND2_X1 u0_u1_u2_U67 (.A2( u0_u1_u2_n105 ) , .A1( u0_u1_u2_n106 ) , .ZN( u0_u1_u2_n117 ) );
  INV_X1 u0_u1_u2_U68 (.ZN( u0_u1_u2_n187 ) , .A( u0_u1_u2_n99 ) );
  OAI21_X1 u0_u1_u2_U69 (.B1( u0_u1_u2_n137 ) , .B2( u0_u1_u2_n143 ) , .A( u0_u1_u2_n98 ) , .ZN( u0_u1_u2_n99 ) );
  AOI21_X1 u0_u1_u2_U7 (.B2( u0_u1_u2_n119 ) , .ZN( u0_u1_u2_n127 ) , .A( u0_u1_u2_n137 ) , .B1( u0_u1_u2_n155 ) );
  NOR2_X1 u0_u1_u2_U70 (.A2( u0_u1_X_16 ) , .ZN( u0_u1_u2_n140 ) , .A1( u0_u1_u2_n166 ) );
  NOR2_X1 u0_u1_u2_U71 (.A2( u0_u1_X_13 ) , .A1( u0_u1_X_14 ) , .ZN( u0_u1_u2_n100 ) );
  NOR2_X1 u0_u1_u2_U72 (.A2( u0_u1_X_16 ) , .A1( u0_u1_X_17 ) , .ZN( u0_u1_u2_n138 ) );
  NOR2_X1 u0_u1_u2_U73 (.A2( u0_u1_X_15 ) , .A1( u0_u1_X_18 ) , .ZN( u0_u1_u2_n104 ) );
  NOR2_X1 u0_u1_u2_U74 (.A2( u0_u1_X_14 ) , .ZN( u0_u1_u2_n103 ) , .A1( u0_u1_u2_n174 ) );
  NOR2_X1 u0_u1_u2_U75 (.A2( u0_u1_X_15 ) , .ZN( u0_u1_u2_n102 ) , .A1( u0_u1_u2_n165 ) );
  NOR2_X1 u0_u1_u2_U76 (.A2( u0_u1_X_17 ) , .ZN( u0_u1_u2_n114 ) , .A1( u0_u1_u2_n169 ) );
  AND2_X1 u0_u1_u2_U77 (.A1( u0_u1_X_15 ) , .ZN( u0_u1_u2_n105 ) , .A2( u0_u1_u2_n165 ) );
  AND2_X1 u0_u1_u2_U78 (.A2( u0_u1_X_15 ) , .A1( u0_u1_X_18 ) , .ZN( u0_u1_u2_n107 ) );
  AND2_X1 u0_u1_u2_U79 (.A1( u0_u1_X_14 ) , .ZN( u0_u1_u2_n106 ) , .A2( u0_u1_u2_n174 ) );
  AOI21_X1 u0_u1_u2_U8 (.ZN( u0_u1_u2_n124 ) , .B1( u0_u1_u2_n131 ) , .B2( u0_u1_u2_n143 ) , .A( u0_u1_u2_n172 ) );
  AND2_X1 u0_u1_u2_U80 (.A1( u0_u1_X_13 ) , .A2( u0_u1_X_14 ) , .ZN( u0_u1_u2_n108 ) );
  INV_X1 u0_u1_u2_U81 (.A( u0_u1_X_16 ) , .ZN( u0_u1_u2_n169 ) );
  INV_X1 u0_u1_u2_U82 (.A( u0_u1_X_17 ) , .ZN( u0_u1_u2_n166 ) );
  INV_X1 u0_u1_u2_U83 (.A( u0_u1_X_13 ) , .ZN( u0_u1_u2_n174 ) );
  INV_X1 u0_u1_u2_U84 (.A( u0_u1_X_18 ) , .ZN( u0_u1_u2_n165 ) );
  NAND4_X1 u0_u1_u2_U85 (.ZN( u0_out1_30 ) , .A4( u0_u1_u2_n147 ) , .A3( u0_u1_u2_n148 ) , .A2( u0_u1_u2_n149 ) , .A1( u0_u1_u2_n187 ) );
  NOR3_X1 u0_u1_u2_U86 (.A3( u0_u1_u2_n144 ) , .A2( u0_u1_u2_n145 ) , .A1( u0_u1_u2_n146 ) , .ZN( u0_u1_u2_n147 ) );
  AOI21_X1 u0_u1_u2_U87 (.B2( u0_u1_u2_n138 ) , .ZN( u0_u1_u2_n148 ) , .A( u0_u1_u2_n162 ) , .B1( u0_u1_u2_n182 ) );
  NAND4_X1 u0_u1_u2_U88 (.ZN( u0_out1_24 ) , .A4( u0_u1_u2_n111 ) , .A3( u0_u1_u2_n112 ) , .A1( u0_u1_u2_n130 ) , .A2( u0_u1_u2_n187 ) );
  AOI221_X1 u0_u1_u2_U89 (.A( u0_u1_u2_n109 ) , .B1( u0_u1_u2_n110 ) , .ZN( u0_u1_u2_n111 ) , .C1( u0_u1_u2_n134 ) , .C2( u0_u1_u2_n170 ) , .B2( u0_u1_u2_n173 ) );
  AOI21_X1 u0_u1_u2_U9 (.B2( u0_u1_u2_n123 ) , .ZN( u0_u1_u2_n125 ) , .A( u0_u1_u2_n171 ) , .B1( u0_u1_u2_n184 ) );
  AOI21_X1 u0_u1_u2_U90 (.ZN( u0_u1_u2_n112 ) , .B2( u0_u1_u2_n156 ) , .A( u0_u1_u2_n164 ) , .B1( u0_u1_u2_n181 ) );
  NAND4_X1 u0_u1_u2_U91 (.ZN( u0_out1_16 ) , .A4( u0_u1_u2_n128 ) , .A3( u0_u1_u2_n129 ) , .A1( u0_u1_u2_n130 ) , .A2( u0_u1_u2_n186 ) );
  AOI22_X1 u0_u1_u2_U92 (.A2( u0_u1_u2_n118 ) , .ZN( u0_u1_u2_n129 ) , .A1( u0_u1_u2_n140 ) , .B1( u0_u1_u2_n157 ) , .B2( u0_u1_u2_n170 ) );
  INV_X1 u0_u1_u2_U93 (.A( u0_u1_u2_n163 ) , .ZN( u0_u1_u2_n186 ) );
  OR4_X1 u0_u1_u2_U94 (.ZN( u0_out1_6 ) , .A4( u0_u1_u2_n161 ) , .A3( u0_u1_u2_n162 ) , .A2( u0_u1_u2_n163 ) , .A1( u0_u1_u2_n164 ) );
  OR3_X1 u0_u1_u2_U95 (.A2( u0_u1_u2_n159 ) , .A1( u0_u1_u2_n160 ) , .ZN( u0_u1_u2_n161 ) , .A3( u0_u1_u2_n183 ) );
  AOI21_X1 u0_u1_u2_U96 (.B2( u0_u1_u2_n154 ) , .B1( u0_u1_u2_n155 ) , .ZN( u0_u1_u2_n159 ) , .A( u0_u1_u2_n167 ) );
  NAND3_X1 u0_u1_u2_U97 (.A2( u0_u1_u2_n117 ) , .A1( u0_u1_u2_n122 ) , .A3( u0_u1_u2_n123 ) , .ZN( u0_u1_u2_n134 ) );
  NAND3_X1 u0_u1_u2_U98 (.ZN( u0_u1_u2_n110 ) , .A2( u0_u1_u2_n131 ) , .A3( u0_u1_u2_n139 ) , .A1( u0_u1_u2_n154 ) );
  NAND3_X1 u0_u1_u2_U99 (.A2( u0_u1_u2_n100 ) , .ZN( u0_u1_u2_n101 ) , .A1( u0_u1_u2_n104 ) , .A3( u0_u1_u2_n114 ) );
  OAI22_X1 u0_u1_u3_U10 (.B1( u0_u1_u3_n113 ) , .A2( u0_u1_u3_n135 ) , .A1( u0_u1_u3_n150 ) , .B2( u0_u1_u3_n164 ) , .ZN( u0_u1_u3_n98 ) );
  OAI211_X1 u0_u1_u3_U11 (.B( u0_u1_u3_n106 ) , .ZN( u0_u1_u3_n119 ) , .C2( u0_u1_u3_n128 ) , .C1( u0_u1_u3_n167 ) , .A( u0_u1_u3_n181 ) );
  AOI221_X1 u0_u1_u3_U12 (.C1( u0_u1_u3_n105 ) , .ZN( u0_u1_u3_n106 ) , .A( u0_u1_u3_n131 ) , .B2( u0_u1_u3_n132 ) , .C2( u0_u1_u3_n133 ) , .B1( u0_u1_u3_n169 ) );
  INV_X1 u0_u1_u3_U13 (.ZN( u0_u1_u3_n181 ) , .A( u0_u1_u3_n98 ) );
  NAND2_X1 u0_u1_u3_U14 (.ZN( u0_u1_u3_n105 ) , .A2( u0_u1_u3_n130 ) , .A1( u0_u1_u3_n155 ) );
  AOI22_X1 u0_u1_u3_U15 (.B1( u0_u1_u3_n115 ) , .A2( u0_u1_u3_n116 ) , .ZN( u0_u1_u3_n123 ) , .B2( u0_u1_u3_n133 ) , .A1( u0_u1_u3_n169 ) );
  NAND2_X1 u0_u1_u3_U16 (.ZN( u0_u1_u3_n116 ) , .A2( u0_u1_u3_n151 ) , .A1( u0_u1_u3_n182 ) );
  NOR2_X1 u0_u1_u3_U17 (.ZN( u0_u1_u3_n126 ) , .A2( u0_u1_u3_n150 ) , .A1( u0_u1_u3_n164 ) );
  AOI21_X1 u0_u1_u3_U18 (.ZN( u0_u1_u3_n112 ) , .B2( u0_u1_u3_n146 ) , .B1( u0_u1_u3_n155 ) , .A( u0_u1_u3_n167 ) );
  NAND2_X1 u0_u1_u3_U19 (.A1( u0_u1_u3_n135 ) , .ZN( u0_u1_u3_n142 ) , .A2( u0_u1_u3_n164 ) );
  NAND2_X1 u0_u1_u3_U20 (.ZN( u0_u1_u3_n132 ) , .A2( u0_u1_u3_n152 ) , .A1( u0_u1_u3_n156 ) );
  AND2_X1 u0_u1_u3_U21 (.A2( u0_u1_u3_n113 ) , .A1( u0_u1_u3_n114 ) , .ZN( u0_u1_u3_n151 ) );
  INV_X1 u0_u1_u3_U22 (.A( u0_u1_u3_n133 ) , .ZN( u0_u1_u3_n165 ) );
  INV_X1 u0_u1_u3_U23 (.A( u0_u1_u3_n135 ) , .ZN( u0_u1_u3_n170 ) );
  NAND2_X1 u0_u1_u3_U24 (.A1( u0_u1_u3_n107 ) , .A2( u0_u1_u3_n108 ) , .ZN( u0_u1_u3_n140 ) );
  NAND2_X1 u0_u1_u3_U25 (.ZN( u0_u1_u3_n117 ) , .A1( u0_u1_u3_n124 ) , .A2( u0_u1_u3_n148 ) );
  NAND2_X1 u0_u1_u3_U26 (.ZN( u0_u1_u3_n143 ) , .A1( u0_u1_u3_n165 ) , .A2( u0_u1_u3_n167 ) );
  INV_X1 u0_u1_u3_U27 (.A( u0_u1_u3_n130 ) , .ZN( u0_u1_u3_n177 ) );
  INV_X1 u0_u1_u3_U28 (.A( u0_u1_u3_n128 ) , .ZN( u0_u1_u3_n176 ) );
  INV_X1 u0_u1_u3_U29 (.A( u0_u1_u3_n155 ) , .ZN( u0_u1_u3_n174 ) );
  INV_X1 u0_u1_u3_U3 (.A( u0_u1_u3_n129 ) , .ZN( u0_u1_u3_n183 ) );
  INV_X1 u0_u1_u3_U30 (.A( u0_u1_u3_n139 ) , .ZN( u0_u1_u3_n185 ) );
  NOR2_X1 u0_u1_u3_U31 (.ZN( u0_u1_u3_n135 ) , .A2( u0_u1_u3_n141 ) , .A1( u0_u1_u3_n169 ) );
  OAI222_X1 u0_u1_u3_U32 (.C2( u0_u1_u3_n107 ) , .A2( u0_u1_u3_n108 ) , .B1( u0_u1_u3_n135 ) , .ZN( u0_u1_u3_n138 ) , .B2( u0_u1_u3_n146 ) , .C1( u0_u1_u3_n154 ) , .A1( u0_u1_u3_n164 ) );
  NOR4_X1 u0_u1_u3_U33 (.A4( u0_u1_u3_n157 ) , .A3( u0_u1_u3_n158 ) , .A2( u0_u1_u3_n159 ) , .A1( u0_u1_u3_n160 ) , .ZN( u0_u1_u3_n161 ) );
  AOI21_X1 u0_u1_u3_U34 (.B2( u0_u1_u3_n152 ) , .B1( u0_u1_u3_n153 ) , .ZN( u0_u1_u3_n158 ) , .A( u0_u1_u3_n164 ) );
  AOI21_X1 u0_u1_u3_U35 (.A( u0_u1_u3_n154 ) , .B2( u0_u1_u3_n155 ) , .B1( u0_u1_u3_n156 ) , .ZN( u0_u1_u3_n157 ) );
  AOI21_X1 u0_u1_u3_U36 (.A( u0_u1_u3_n149 ) , .B2( u0_u1_u3_n150 ) , .B1( u0_u1_u3_n151 ) , .ZN( u0_u1_u3_n159 ) );
  AOI211_X1 u0_u1_u3_U37 (.ZN( u0_u1_u3_n109 ) , .A( u0_u1_u3_n119 ) , .C2( u0_u1_u3_n129 ) , .B( u0_u1_u3_n138 ) , .C1( u0_u1_u3_n141 ) );
  AOI211_X1 u0_u1_u3_U38 (.B( u0_u1_u3_n119 ) , .A( u0_u1_u3_n120 ) , .C2( u0_u1_u3_n121 ) , .ZN( u0_u1_u3_n122 ) , .C1( u0_u1_u3_n179 ) );
  INV_X1 u0_u1_u3_U39 (.A( u0_u1_u3_n156 ) , .ZN( u0_u1_u3_n179 ) );
  INV_X1 u0_u1_u3_U4 (.A( u0_u1_u3_n140 ) , .ZN( u0_u1_u3_n182 ) );
  OAI22_X1 u0_u1_u3_U40 (.B1( u0_u1_u3_n118 ) , .ZN( u0_u1_u3_n120 ) , .A1( u0_u1_u3_n135 ) , .B2( u0_u1_u3_n154 ) , .A2( u0_u1_u3_n178 ) );
  AND3_X1 u0_u1_u3_U41 (.ZN( u0_u1_u3_n118 ) , .A2( u0_u1_u3_n124 ) , .A1( u0_u1_u3_n144 ) , .A3( u0_u1_u3_n152 ) );
  INV_X1 u0_u1_u3_U42 (.A( u0_u1_u3_n121 ) , .ZN( u0_u1_u3_n164 ) );
  NAND2_X1 u0_u1_u3_U43 (.ZN( u0_u1_u3_n133 ) , .A1( u0_u1_u3_n154 ) , .A2( u0_u1_u3_n164 ) );
  OAI211_X1 u0_u1_u3_U44 (.B( u0_u1_u3_n127 ) , .ZN( u0_u1_u3_n139 ) , .C1( u0_u1_u3_n150 ) , .C2( u0_u1_u3_n154 ) , .A( u0_u1_u3_n184 ) );
  INV_X1 u0_u1_u3_U45 (.A( u0_u1_u3_n125 ) , .ZN( u0_u1_u3_n184 ) );
  AOI221_X1 u0_u1_u3_U46 (.A( u0_u1_u3_n126 ) , .ZN( u0_u1_u3_n127 ) , .C2( u0_u1_u3_n132 ) , .C1( u0_u1_u3_n169 ) , .B2( u0_u1_u3_n170 ) , .B1( u0_u1_u3_n174 ) );
  OAI22_X1 u0_u1_u3_U47 (.A1( u0_u1_u3_n124 ) , .ZN( u0_u1_u3_n125 ) , .B2( u0_u1_u3_n145 ) , .A2( u0_u1_u3_n165 ) , .B1( u0_u1_u3_n167 ) );
  NOR2_X1 u0_u1_u3_U48 (.A1( u0_u1_u3_n113 ) , .ZN( u0_u1_u3_n131 ) , .A2( u0_u1_u3_n154 ) );
  NAND2_X1 u0_u1_u3_U49 (.A1( u0_u1_u3_n103 ) , .ZN( u0_u1_u3_n150 ) , .A2( u0_u1_u3_n99 ) );
  INV_X1 u0_u1_u3_U5 (.A( u0_u1_u3_n117 ) , .ZN( u0_u1_u3_n178 ) );
  NAND2_X1 u0_u1_u3_U50 (.A2( u0_u1_u3_n102 ) , .ZN( u0_u1_u3_n155 ) , .A1( u0_u1_u3_n97 ) );
  INV_X1 u0_u1_u3_U51 (.A( u0_u1_u3_n141 ) , .ZN( u0_u1_u3_n167 ) );
  AOI21_X1 u0_u1_u3_U52 (.B2( u0_u1_u3_n114 ) , .B1( u0_u1_u3_n146 ) , .A( u0_u1_u3_n154 ) , .ZN( u0_u1_u3_n94 ) );
  AOI21_X1 u0_u1_u3_U53 (.ZN( u0_u1_u3_n110 ) , .B2( u0_u1_u3_n142 ) , .B1( u0_u1_u3_n186 ) , .A( u0_u1_u3_n95 ) );
  INV_X1 u0_u1_u3_U54 (.A( u0_u1_u3_n145 ) , .ZN( u0_u1_u3_n186 ) );
  AOI21_X1 u0_u1_u3_U55 (.B1( u0_u1_u3_n124 ) , .A( u0_u1_u3_n149 ) , .B2( u0_u1_u3_n155 ) , .ZN( u0_u1_u3_n95 ) );
  INV_X1 u0_u1_u3_U56 (.A( u0_u1_u3_n149 ) , .ZN( u0_u1_u3_n169 ) );
  NAND2_X1 u0_u1_u3_U57 (.ZN( u0_u1_u3_n124 ) , .A1( u0_u1_u3_n96 ) , .A2( u0_u1_u3_n97 ) );
  NAND2_X1 u0_u1_u3_U58 (.A2( u0_u1_u3_n100 ) , .ZN( u0_u1_u3_n146 ) , .A1( u0_u1_u3_n96 ) );
  NAND2_X1 u0_u1_u3_U59 (.A1( u0_u1_u3_n101 ) , .ZN( u0_u1_u3_n145 ) , .A2( u0_u1_u3_n99 ) );
  AOI221_X1 u0_u1_u3_U6 (.A( u0_u1_u3_n131 ) , .C2( u0_u1_u3_n132 ) , .C1( u0_u1_u3_n133 ) , .ZN( u0_u1_u3_n134 ) , .B1( u0_u1_u3_n143 ) , .B2( u0_u1_u3_n177 ) );
  NAND2_X1 u0_u1_u3_U60 (.A1( u0_u1_u3_n100 ) , .ZN( u0_u1_u3_n156 ) , .A2( u0_u1_u3_n99 ) );
  NAND2_X1 u0_u1_u3_U61 (.A2( u0_u1_u3_n101 ) , .A1( u0_u1_u3_n104 ) , .ZN( u0_u1_u3_n148 ) );
  NAND2_X1 u0_u1_u3_U62 (.A1( u0_u1_u3_n100 ) , .A2( u0_u1_u3_n102 ) , .ZN( u0_u1_u3_n128 ) );
  NAND2_X1 u0_u1_u3_U63 (.A2( u0_u1_u3_n101 ) , .A1( u0_u1_u3_n102 ) , .ZN( u0_u1_u3_n152 ) );
  NAND2_X1 u0_u1_u3_U64 (.A2( u0_u1_u3_n101 ) , .ZN( u0_u1_u3_n114 ) , .A1( u0_u1_u3_n96 ) );
  NAND2_X1 u0_u1_u3_U65 (.ZN( u0_u1_u3_n107 ) , .A1( u0_u1_u3_n97 ) , .A2( u0_u1_u3_n99 ) );
  NAND2_X1 u0_u1_u3_U66 (.A2( u0_u1_u3_n100 ) , .A1( u0_u1_u3_n104 ) , .ZN( u0_u1_u3_n113 ) );
  NAND2_X1 u0_u1_u3_U67 (.A1( u0_u1_u3_n104 ) , .ZN( u0_u1_u3_n153 ) , .A2( u0_u1_u3_n97 ) );
  NAND2_X1 u0_u1_u3_U68 (.A2( u0_u1_u3_n103 ) , .A1( u0_u1_u3_n104 ) , .ZN( u0_u1_u3_n130 ) );
  NAND2_X1 u0_u1_u3_U69 (.A2( u0_u1_u3_n103 ) , .ZN( u0_u1_u3_n144 ) , .A1( u0_u1_u3_n96 ) );
  OAI22_X1 u0_u1_u3_U7 (.B2( u0_u1_u3_n147 ) , .A2( u0_u1_u3_n148 ) , .ZN( u0_u1_u3_n160 ) , .B1( u0_u1_u3_n165 ) , .A1( u0_u1_u3_n168 ) );
  NAND2_X1 u0_u1_u3_U70 (.A1( u0_u1_u3_n102 ) , .A2( u0_u1_u3_n103 ) , .ZN( u0_u1_u3_n108 ) );
  NOR2_X1 u0_u1_u3_U71 (.A2( u0_u1_X_19 ) , .A1( u0_u1_X_20 ) , .ZN( u0_u1_u3_n99 ) );
  NOR2_X1 u0_u1_u3_U72 (.A2( u0_u1_X_21 ) , .A1( u0_u1_X_24 ) , .ZN( u0_u1_u3_n103 ) );
  NOR2_X1 u0_u1_u3_U73 (.A2( u0_u1_X_24 ) , .A1( u0_u1_u3_n171 ) , .ZN( u0_u1_u3_n97 ) );
  NOR2_X1 u0_u1_u3_U74 (.A2( u0_u1_X_23 ) , .ZN( u0_u1_u3_n141 ) , .A1( u0_u1_u3_n166 ) );
  NOR2_X1 u0_u1_u3_U75 (.A2( u0_u1_X_19 ) , .A1( u0_u1_u3_n172 ) , .ZN( u0_u1_u3_n96 ) );
  NAND2_X1 u0_u1_u3_U76 (.A1( u0_u1_X_22 ) , .A2( u0_u1_X_23 ) , .ZN( u0_u1_u3_n154 ) );
  NAND2_X1 u0_u1_u3_U77 (.A1( u0_u1_X_23 ) , .ZN( u0_u1_u3_n149 ) , .A2( u0_u1_u3_n166 ) );
  NOR2_X1 u0_u1_u3_U78 (.A2( u0_u1_X_22 ) , .A1( u0_u1_X_23 ) , .ZN( u0_u1_u3_n121 ) );
  AND2_X1 u0_u1_u3_U79 (.A1( u0_u1_X_24 ) , .ZN( u0_u1_u3_n101 ) , .A2( u0_u1_u3_n171 ) );
  AND3_X1 u0_u1_u3_U8 (.A3( u0_u1_u3_n144 ) , .A2( u0_u1_u3_n145 ) , .A1( u0_u1_u3_n146 ) , .ZN( u0_u1_u3_n147 ) );
  AND2_X1 u0_u1_u3_U80 (.A1( u0_u1_X_19 ) , .ZN( u0_u1_u3_n102 ) , .A2( u0_u1_u3_n172 ) );
  AND2_X1 u0_u1_u3_U81 (.A1( u0_u1_X_21 ) , .A2( u0_u1_X_24 ) , .ZN( u0_u1_u3_n100 ) );
  AND2_X1 u0_u1_u3_U82 (.A2( u0_u1_X_19 ) , .A1( u0_u1_X_20 ) , .ZN( u0_u1_u3_n104 ) );
  INV_X1 u0_u1_u3_U83 (.A( u0_u1_X_22 ) , .ZN( u0_u1_u3_n166 ) );
  INV_X1 u0_u1_u3_U84 (.A( u0_u1_X_21 ) , .ZN( u0_u1_u3_n171 ) );
  INV_X1 u0_u1_u3_U85 (.A( u0_u1_X_20 ) , .ZN( u0_u1_u3_n172 ) );
  OR4_X1 u0_u1_u3_U86 (.ZN( u0_out1_10 ) , .A4( u0_u1_u3_n136 ) , .A3( u0_u1_u3_n137 ) , .A1( u0_u1_u3_n138 ) , .A2( u0_u1_u3_n139 ) );
  OAI222_X1 u0_u1_u3_U87 (.C1( u0_u1_u3_n128 ) , .ZN( u0_u1_u3_n137 ) , .B1( u0_u1_u3_n148 ) , .A2( u0_u1_u3_n150 ) , .B2( u0_u1_u3_n154 ) , .C2( u0_u1_u3_n164 ) , .A1( u0_u1_u3_n167 ) );
  OAI221_X1 u0_u1_u3_U88 (.A( u0_u1_u3_n134 ) , .B2( u0_u1_u3_n135 ) , .ZN( u0_u1_u3_n136 ) , .C1( u0_u1_u3_n149 ) , .B1( u0_u1_u3_n151 ) , .C2( u0_u1_u3_n183 ) );
  NAND4_X1 u0_u1_u3_U89 (.ZN( u0_out1_26 ) , .A4( u0_u1_u3_n109 ) , .A3( u0_u1_u3_n110 ) , .A2( u0_u1_u3_n111 ) , .A1( u0_u1_u3_n173 ) );
  INV_X1 u0_u1_u3_U9 (.A( u0_u1_u3_n143 ) , .ZN( u0_u1_u3_n168 ) );
  INV_X1 u0_u1_u3_U90 (.ZN( u0_u1_u3_n173 ) , .A( u0_u1_u3_n94 ) );
  OAI21_X1 u0_u1_u3_U91 (.ZN( u0_u1_u3_n111 ) , .B2( u0_u1_u3_n117 ) , .A( u0_u1_u3_n133 ) , .B1( u0_u1_u3_n176 ) );
  NAND4_X1 u0_u1_u3_U92 (.ZN( u0_out1_20 ) , .A4( u0_u1_u3_n122 ) , .A3( u0_u1_u3_n123 ) , .A1( u0_u1_u3_n175 ) , .A2( u0_u1_u3_n180 ) );
  INV_X1 u0_u1_u3_U93 (.A( u0_u1_u3_n112 ) , .ZN( u0_u1_u3_n175 ) );
  INV_X1 u0_u1_u3_U94 (.A( u0_u1_u3_n126 ) , .ZN( u0_u1_u3_n180 ) );
  NAND4_X1 u0_u1_u3_U95 (.ZN( u0_out1_1 ) , .A4( u0_u1_u3_n161 ) , .A3( u0_u1_u3_n162 ) , .A2( u0_u1_u3_n163 ) , .A1( u0_u1_u3_n185 ) );
  NAND2_X1 u0_u1_u3_U96 (.ZN( u0_u1_u3_n163 ) , .A2( u0_u1_u3_n170 ) , .A1( u0_u1_u3_n176 ) );
  AOI22_X1 u0_u1_u3_U97 (.B2( u0_u1_u3_n140 ) , .B1( u0_u1_u3_n141 ) , .A2( u0_u1_u3_n142 ) , .ZN( u0_u1_u3_n162 ) , .A1( u0_u1_u3_n177 ) );
  NAND3_X1 u0_u1_u3_U98 (.A1( u0_u1_u3_n114 ) , .ZN( u0_u1_u3_n115 ) , .A2( u0_u1_u3_n145 ) , .A3( u0_u1_u3_n153 ) );
  NAND3_X1 u0_u1_u3_U99 (.ZN( u0_u1_u3_n129 ) , .A2( u0_u1_u3_n144 ) , .A1( u0_u1_u3_n153 ) , .A3( u0_u1_u3_n182 ) );
  XOR2_X1 u0_u7_U33 (.B( u0_K8_24 ) , .A( u0_R6_17 ) , .Z( u0_u7_X_24 ) );
  XOR2_X1 u0_u7_U34 (.B( u0_K8_23 ) , .A( u0_R6_16 ) , .Z( u0_u7_X_23 ) );
  XOR2_X1 u0_u7_U35 (.B( u0_K8_22 ) , .A( u0_R6_15 ) , .Z( u0_u7_X_22 ) );
  XOR2_X1 u0_u7_U36 (.B( u0_K8_21 ) , .A( u0_R6_14 ) , .Z( u0_u7_X_21 ) );
  XOR2_X1 u0_u7_U37 (.B( u0_K8_20 ) , .A( u0_R6_13 ) , .Z( u0_u7_X_20 ) );
  XOR2_X1 u0_u7_U39 (.B( u0_K8_19 ) , .A( u0_R6_12 ) , .Z( u0_u7_X_19 ) );
  XOR2_X1 u0_u7_U40 (.B( u0_K8_18 ) , .A( u0_R6_13 ) , .Z( u0_u7_X_18 ) );
  XOR2_X1 u0_u7_U41 (.B( u0_K8_17 ) , .A( u0_R6_12 ) , .Z( u0_u7_X_17 ) );
  XOR2_X1 u0_u7_U42 (.B( u0_K8_16 ) , .A( u0_R6_11 ) , .Z( u0_u7_X_16 ) );
  XOR2_X1 u0_u7_U43 (.B( u0_K8_15 ) , .A( u0_R6_10 ) , .Z( u0_u7_X_15 ) );
  XOR2_X1 u0_u7_U44 (.B( u0_K8_14 ) , .A( u0_R6_9 ) , .Z( u0_u7_X_14 ) );
  XOR2_X1 u0_u7_U45 (.B( u0_K8_13 ) , .A( u0_R6_8 ) , .Z( u0_u7_X_13 ) );
  OAI22_X1 u0_u7_u2_U10 (.ZN( u0_u7_u2_n109 ) , .A2( u0_u7_u2_n113 ) , .B2( u0_u7_u2_n133 ) , .B1( u0_u7_u2_n167 ) , .A1( u0_u7_u2_n168 ) );
  NAND3_X1 u0_u7_u2_U100 (.A2( u0_u7_u2_n100 ) , .A1( u0_u7_u2_n104 ) , .A3( u0_u7_u2_n138 ) , .ZN( u0_u7_u2_n98 ) );
  OAI22_X1 u0_u7_u2_U11 (.B1( u0_u7_u2_n151 ) , .A2( u0_u7_u2_n152 ) , .A1( u0_u7_u2_n153 ) , .ZN( u0_u7_u2_n160 ) , .B2( u0_u7_u2_n168 ) );
  NOR3_X1 u0_u7_u2_U12 (.A1( u0_u7_u2_n150 ) , .ZN( u0_u7_u2_n151 ) , .A3( u0_u7_u2_n175 ) , .A2( u0_u7_u2_n188 ) );
  AOI21_X1 u0_u7_u2_U13 (.ZN( u0_u7_u2_n144 ) , .B2( u0_u7_u2_n155 ) , .A( u0_u7_u2_n172 ) , .B1( u0_u7_u2_n185 ) );
  AOI21_X1 u0_u7_u2_U14 (.B2( u0_u7_u2_n143 ) , .ZN( u0_u7_u2_n145 ) , .B1( u0_u7_u2_n152 ) , .A( u0_u7_u2_n171 ) );
  AOI21_X1 u0_u7_u2_U15 (.B2( u0_u7_u2_n120 ) , .B1( u0_u7_u2_n121 ) , .ZN( u0_u7_u2_n126 ) , .A( u0_u7_u2_n167 ) );
  INV_X1 u0_u7_u2_U16 (.A( u0_u7_u2_n156 ) , .ZN( u0_u7_u2_n171 ) );
  INV_X1 u0_u7_u2_U17 (.A( u0_u7_u2_n120 ) , .ZN( u0_u7_u2_n188 ) );
  NAND2_X1 u0_u7_u2_U18 (.A2( u0_u7_u2_n122 ) , .ZN( u0_u7_u2_n150 ) , .A1( u0_u7_u2_n152 ) );
  INV_X1 u0_u7_u2_U19 (.A( u0_u7_u2_n153 ) , .ZN( u0_u7_u2_n170 ) );
  INV_X1 u0_u7_u2_U20 (.A( u0_u7_u2_n137 ) , .ZN( u0_u7_u2_n173 ) );
  NAND2_X1 u0_u7_u2_U21 (.A1( u0_u7_u2_n132 ) , .A2( u0_u7_u2_n139 ) , .ZN( u0_u7_u2_n157 ) );
  INV_X1 u0_u7_u2_U22 (.A( u0_u7_u2_n113 ) , .ZN( u0_u7_u2_n178 ) );
  INV_X1 u0_u7_u2_U23 (.A( u0_u7_u2_n139 ) , .ZN( u0_u7_u2_n175 ) );
  INV_X1 u0_u7_u2_U24 (.A( u0_u7_u2_n155 ) , .ZN( u0_u7_u2_n181 ) );
  INV_X1 u0_u7_u2_U25 (.A( u0_u7_u2_n119 ) , .ZN( u0_u7_u2_n177 ) );
  INV_X1 u0_u7_u2_U26 (.A( u0_u7_u2_n116 ) , .ZN( u0_u7_u2_n180 ) );
  INV_X1 u0_u7_u2_U27 (.A( u0_u7_u2_n131 ) , .ZN( u0_u7_u2_n179 ) );
  INV_X1 u0_u7_u2_U28 (.A( u0_u7_u2_n154 ) , .ZN( u0_u7_u2_n176 ) );
  NAND2_X1 u0_u7_u2_U29 (.A2( u0_u7_u2_n116 ) , .A1( u0_u7_u2_n117 ) , .ZN( u0_u7_u2_n118 ) );
  NOR2_X1 u0_u7_u2_U3 (.ZN( u0_u7_u2_n121 ) , .A2( u0_u7_u2_n177 ) , .A1( u0_u7_u2_n180 ) );
  INV_X1 u0_u7_u2_U30 (.A( u0_u7_u2_n132 ) , .ZN( u0_u7_u2_n182 ) );
  INV_X1 u0_u7_u2_U31 (.A( u0_u7_u2_n158 ) , .ZN( u0_u7_u2_n183 ) );
  OAI21_X1 u0_u7_u2_U32 (.A( u0_u7_u2_n156 ) , .B1( u0_u7_u2_n157 ) , .ZN( u0_u7_u2_n158 ) , .B2( u0_u7_u2_n179 ) );
  NOR2_X1 u0_u7_u2_U33 (.ZN( u0_u7_u2_n156 ) , .A1( u0_u7_u2_n166 ) , .A2( u0_u7_u2_n169 ) );
  NOR2_X1 u0_u7_u2_U34 (.A2( u0_u7_u2_n114 ) , .ZN( u0_u7_u2_n137 ) , .A1( u0_u7_u2_n140 ) );
  NOR2_X1 u0_u7_u2_U35 (.A2( u0_u7_u2_n138 ) , .ZN( u0_u7_u2_n153 ) , .A1( u0_u7_u2_n156 ) );
  AOI211_X1 u0_u7_u2_U36 (.ZN( u0_u7_u2_n130 ) , .C1( u0_u7_u2_n138 ) , .C2( u0_u7_u2_n179 ) , .B( u0_u7_u2_n96 ) , .A( u0_u7_u2_n97 ) );
  OAI22_X1 u0_u7_u2_U37 (.B1( u0_u7_u2_n133 ) , .A2( u0_u7_u2_n137 ) , .A1( u0_u7_u2_n152 ) , .B2( u0_u7_u2_n168 ) , .ZN( u0_u7_u2_n97 ) );
  OAI221_X1 u0_u7_u2_U38 (.B1( u0_u7_u2_n113 ) , .C1( u0_u7_u2_n132 ) , .A( u0_u7_u2_n149 ) , .B2( u0_u7_u2_n171 ) , .C2( u0_u7_u2_n172 ) , .ZN( u0_u7_u2_n96 ) );
  OAI221_X1 u0_u7_u2_U39 (.A( u0_u7_u2_n115 ) , .C2( u0_u7_u2_n123 ) , .B2( u0_u7_u2_n143 ) , .B1( u0_u7_u2_n153 ) , .ZN( u0_u7_u2_n163 ) , .C1( u0_u7_u2_n168 ) );
  INV_X1 u0_u7_u2_U4 (.A( u0_u7_u2_n134 ) , .ZN( u0_u7_u2_n185 ) );
  OAI21_X1 u0_u7_u2_U40 (.A( u0_u7_u2_n114 ) , .ZN( u0_u7_u2_n115 ) , .B1( u0_u7_u2_n176 ) , .B2( u0_u7_u2_n178 ) );
  OAI221_X1 u0_u7_u2_U41 (.A( u0_u7_u2_n135 ) , .B2( u0_u7_u2_n136 ) , .B1( u0_u7_u2_n137 ) , .ZN( u0_u7_u2_n162 ) , .C2( u0_u7_u2_n167 ) , .C1( u0_u7_u2_n185 ) );
  AND3_X1 u0_u7_u2_U42 (.A3( u0_u7_u2_n131 ) , .A2( u0_u7_u2_n132 ) , .A1( u0_u7_u2_n133 ) , .ZN( u0_u7_u2_n136 ) );
  AOI22_X1 u0_u7_u2_U43 (.ZN( u0_u7_u2_n135 ) , .B1( u0_u7_u2_n140 ) , .A1( u0_u7_u2_n156 ) , .B2( u0_u7_u2_n180 ) , .A2( u0_u7_u2_n188 ) );
  AOI21_X1 u0_u7_u2_U44 (.ZN( u0_u7_u2_n149 ) , .B1( u0_u7_u2_n173 ) , .B2( u0_u7_u2_n188 ) , .A( u0_u7_u2_n95 ) );
  AND3_X1 u0_u7_u2_U45 (.A2( u0_u7_u2_n100 ) , .A1( u0_u7_u2_n104 ) , .A3( u0_u7_u2_n156 ) , .ZN( u0_u7_u2_n95 ) );
  OAI21_X1 u0_u7_u2_U46 (.A( u0_u7_u2_n101 ) , .B2( u0_u7_u2_n121 ) , .B1( u0_u7_u2_n153 ) , .ZN( u0_u7_u2_n164 ) );
  NAND2_X1 u0_u7_u2_U47 (.A2( u0_u7_u2_n100 ) , .A1( u0_u7_u2_n107 ) , .ZN( u0_u7_u2_n155 ) );
  NAND2_X1 u0_u7_u2_U48 (.A2( u0_u7_u2_n105 ) , .A1( u0_u7_u2_n108 ) , .ZN( u0_u7_u2_n143 ) );
  NAND2_X1 u0_u7_u2_U49 (.A1( u0_u7_u2_n104 ) , .A2( u0_u7_u2_n106 ) , .ZN( u0_u7_u2_n152 ) );
  INV_X1 u0_u7_u2_U5 (.A( u0_u7_u2_n150 ) , .ZN( u0_u7_u2_n184 ) );
  NAND2_X1 u0_u7_u2_U50 (.A1( u0_u7_u2_n100 ) , .A2( u0_u7_u2_n105 ) , .ZN( u0_u7_u2_n132 ) );
  INV_X1 u0_u7_u2_U51 (.A( u0_u7_u2_n140 ) , .ZN( u0_u7_u2_n168 ) );
  INV_X1 u0_u7_u2_U52 (.A( u0_u7_u2_n138 ) , .ZN( u0_u7_u2_n167 ) );
  OAI21_X1 u0_u7_u2_U53 (.A( u0_u7_u2_n141 ) , .B2( u0_u7_u2_n142 ) , .ZN( u0_u7_u2_n146 ) , .B1( u0_u7_u2_n153 ) );
  OAI21_X1 u0_u7_u2_U54 (.A( u0_u7_u2_n140 ) , .ZN( u0_u7_u2_n141 ) , .B1( u0_u7_u2_n176 ) , .B2( u0_u7_u2_n177 ) );
  NOR3_X1 u0_u7_u2_U55 (.ZN( u0_u7_u2_n142 ) , .A3( u0_u7_u2_n175 ) , .A2( u0_u7_u2_n178 ) , .A1( u0_u7_u2_n181 ) );
  INV_X1 u0_u7_u2_U56 (.ZN( u0_u7_u2_n187 ) , .A( u0_u7_u2_n99 ) );
  OAI21_X1 u0_u7_u2_U57 (.B1( u0_u7_u2_n137 ) , .B2( u0_u7_u2_n143 ) , .A( u0_u7_u2_n98 ) , .ZN( u0_u7_u2_n99 ) );
  NAND2_X1 u0_u7_u2_U58 (.A1( u0_u7_u2_n102 ) , .A2( u0_u7_u2_n106 ) , .ZN( u0_u7_u2_n113 ) );
  NAND2_X1 u0_u7_u2_U59 (.A1( u0_u7_u2_n106 ) , .A2( u0_u7_u2_n107 ) , .ZN( u0_u7_u2_n131 ) );
  NOR4_X1 u0_u7_u2_U6 (.A4( u0_u7_u2_n124 ) , .A3( u0_u7_u2_n125 ) , .A2( u0_u7_u2_n126 ) , .A1( u0_u7_u2_n127 ) , .ZN( u0_u7_u2_n128 ) );
  NAND2_X1 u0_u7_u2_U60 (.A1( u0_u7_u2_n103 ) , .A2( u0_u7_u2_n107 ) , .ZN( u0_u7_u2_n139 ) );
  NAND2_X1 u0_u7_u2_U61 (.A1( u0_u7_u2_n103 ) , .A2( u0_u7_u2_n105 ) , .ZN( u0_u7_u2_n133 ) );
  NAND2_X1 u0_u7_u2_U62 (.A1( u0_u7_u2_n102 ) , .A2( u0_u7_u2_n103 ) , .ZN( u0_u7_u2_n154 ) );
  NAND2_X1 u0_u7_u2_U63 (.A2( u0_u7_u2_n103 ) , .A1( u0_u7_u2_n104 ) , .ZN( u0_u7_u2_n119 ) );
  NAND2_X1 u0_u7_u2_U64 (.A2( u0_u7_u2_n107 ) , .A1( u0_u7_u2_n108 ) , .ZN( u0_u7_u2_n123 ) );
  NAND2_X1 u0_u7_u2_U65 (.A1( u0_u7_u2_n104 ) , .A2( u0_u7_u2_n108 ) , .ZN( u0_u7_u2_n122 ) );
  INV_X1 u0_u7_u2_U66 (.A( u0_u7_u2_n114 ) , .ZN( u0_u7_u2_n172 ) );
  NAND2_X1 u0_u7_u2_U67 (.A2( u0_u7_u2_n100 ) , .A1( u0_u7_u2_n102 ) , .ZN( u0_u7_u2_n116 ) );
  NAND2_X1 u0_u7_u2_U68 (.A1( u0_u7_u2_n102 ) , .A2( u0_u7_u2_n108 ) , .ZN( u0_u7_u2_n120 ) );
  NAND2_X1 u0_u7_u2_U69 (.A2( u0_u7_u2_n105 ) , .A1( u0_u7_u2_n106 ) , .ZN( u0_u7_u2_n117 ) );
  AOI21_X1 u0_u7_u2_U7 (.B2( u0_u7_u2_n119 ) , .ZN( u0_u7_u2_n127 ) , .A( u0_u7_u2_n137 ) , .B1( u0_u7_u2_n155 ) );
  NOR2_X1 u0_u7_u2_U70 (.A2( u0_u7_X_16 ) , .ZN( u0_u7_u2_n140 ) , .A1( u0_u7_u2_n166 ) );
  NOR2_X1 u0_u7_u2_U71 (.A2( u0_u7_X_13 ) , .A1( u0_u7_X_14 ) , .ZN( u0_u7_u2_n100 ) );
  NOR2_X1 u0_u7_u2_U72 (.A2( u0_u7_X_16 ) , .A1( u0_u7_X_17 ) , .ZN( u0_u7_u2_n138 ) );
  NOR2_X1 u0_u7_u2_U73 (.A2( u0_u7_X_15 ) , .A1( u0_u7_X_18 ) , .ZN( u0_u7_u2_n104 ) );
  NOR2_X1 u0_u7_u2_U74 (.A2( u0_u7_X_14 ) , .ZN( u0_u7_u2_n103 ) , .A1( u0_u7_u2_n174 ) );
  NOR2_X1 u0_u7_u2_U75 (.A2( u0_u7_X_15 ) , .ZN( u0_u7_u2_n102 ) , .A1( u0_u7_u2_n165 ) );
  NOR2_X1 u0_u7_u2_U76 (.A2( u0_u7_X_17 ) , .ZN( u0_u7_u2_n114 ) , .A1( u0_u7_u2_n169 ) );
  AND2_X1 u0_u7_u2_U77 (.A1( u0_u7_X_15 ) , .ZN( u0_u7_u2_n105 ) , .A2( u0_u7_u2_n165 ) );
  AND2_X1 u0_u7_u2_U78 (.A2( u0_u7_X_15 ) , .A1( u0_u7_X_18 ) , .ZN( u0_u7_u2_n107 ) );
  AND2_X1 u0_u7_u2_U79 (.A1( u0_u7_X_14 ) , .ZN( u0_u7_u2_n106 ) , .A2( u0_u7_u2_n174 ) );
  AOI21_X1 u0_u7_u2_U8 (.ZN( u0_u7_u2_n124 ) , .B1( u0_u7_u2_n131 ) , .B2( u0_u7_u2_n143 ) , .A( u0_u7_u2_n172 ) );
  AND2_X1 u0_u7_u2_U80 (.A1( u0_u7_X_13 ) , .A2( u0_u7_X_14 ) , .ZN( u0_u7_u2_n108 ) );
  INV_X1 u0_u7_u2_U81 (.A( u0_u7_X_16 ) , .ZN( u0_u7_u2_n169 ) );
  INV_X1 u0_u7_u2_U82 (.A( u0_u7_X_17 ) , .ZN( u0_u7_u2_n166 ) );
  INV_X1 u0_u7_u2_U83 (.A( u0_u7_X_13 ) , .ZN( u0_u7_u2_n174 ) );
  INV_X1 u0_u7_u2_U84 (.A( u0_u7_X_18 ) , .ZN( u0_u7_u2_n165 ) );
  NAND4_X1 u0_u7_u2_U85 (.ZN( u0_out7_30 ) , .A4( u0_u7_u2_n147 ) , .A3( u0_u7_u2_n148 ) , .A2( u0_u7_u2_n149 ) , .A1( u0_u7_u2_n187 ) );
  NOR3_X1 u0_u7_u2_U86 (.A3( u0_u7_u2_n144 ) , .A2( u0_u7_u2_n145 ) , .A1( u0_u7_u2_n146 ) , .ZN( u0_u7_u2_n147 ) );
  AOI21_X1 u0_u7_u2_U87 (.B2( u0_u7_u2_n138 ) , .ZN( u0_u7_u2_n148 ) , .A( u0_u7_u2_n162 ) , .B1( u0_u7_u2_n182 ) );
  NAND4_X1 u0_u7_u2_U88 (.ZN( u0_out7_24 ) , .A4( u0_u7_u2_n111 ) , .A3( u0_u7_u2_n112 ) , .A1( u0_u7_u2_n130 ) , .A2( u0_u7_u2_n187 ) );
  AOI221_X1 u0_u7_u2_U89 (.A( u0_u7_u2_n109 ) , .B1( u0_u7_u2_n110 ) , .ZN( u0_u7_u2_n111 ) , .C1( u0_u7_u2_n134 ) , .C2( u0_u7_u2_n170 ) , .B2( u0_u7_u2_n173 ) );
  AOI21_X1 u0_u7_u2_U9 (.B2( u0_u7_u2_n123 ) , .ZN( u0_u7_u2_n125 ) , .A( u0_u7_u2_n171 ) , .B1( u0_u7_u2_n184 ) );
  AOI21_X1 u0_u7_u2_U90 (.ZN( u0_u7_u2_n112 ) , .B2( u0_u7_u2_n156 ) , .A( u0_u7_u2_n164 ) , .B1( u0_u7_u2_n181 ) );
  NAND4_X1 u0_u7_u2_U91 (.ZN( u0_out7_16 ) , .A4( u0_u7_u2_n128 ) , .A3( u0_u7_u2_n129 ) , .A1( u0_u7_u2_n130 ) , .A2( u0_u7_u2_n186 ) );
  AOI22_X1 u0_u7_u2_U92 (.A2( u0_u7_u2_n118 ) , .ZN( u0_u7_u2_n129 ) , .A1( u0_u7_u2_n140 ) , .B1( u0_u7_u2_n157 ) , .B2( u0_u7_u2_n170 ) );
  INV_X1 u0_u7_u2_U93 (.A( u0_u7_u2_n163 ) , .ZN( u0_u7_u2_n186 ) );
  OR4_X1 u0_u7_u2_U94 (.ZN( u0_out7_6 ) , .A4( u0_u7_u2_n161 ) , .A3( u0_u7_u2_n162 ) , .A2( u0_u7_u2_n163 ) , .A1( u0_u7_u2_n164 ) );
  OR3_X1 u0_u7_u2_U95 (.A2( u0_u7_u2_n159 ) , .A1( u0_u7_u2_n160 ) , .ZN( u0_u7_u2_n161 ) , .A3( u0_u7_u2_n183 ) );
  AOI21_X1 u0_u7_u2_U96 (.B2( u0_u7_u2_n154 ) , .B1( u0_u7_u2_n155 ) , .ZN( u0_u7_u2_n159 ) , .A( u0_u7_u2_n167 ) );
  NAND3_X1 u0_u7_u2_U97 (.A2( u0_u7_u2_n117 ) , .A1( u0_u7_u2_n122 ) , .A3( u0_u7_u2_n123 ) , .ZN( u0_u7_u2_n134 ) );
  NAND3_X1 u0_u7_u2_U98 (.ZN( u0_u7_u2_n110 ) , .A2( u0_u7_u2_n131 ) , .A3( u0_u7_u2_n139 ) , .A1( u0_u7_u2_n154 ) );
  NAND3_X1 u0_u7_u2_U99 (.A2( u0_u7_u2_n100 ) , .ZN( u0_u7_u2_n101 ) , .A1( u0_u7_u2_n104 ) , .A3( u0_u7_u2_n114 ) );
  OAI22_X1 u0_u7_u3_U10 (.B1( u0_u7_u3_n113 ) , .A2( u0_u7_u3_n135 ) , .A1( u0_u7_u3_n150 ) , .B2( u0_u7_u3_n164 ) , .ZN( u0_u7_u3_n98 ) );
  OAI211_X1 u0_u7_u3_U11 (.B( u0_u7_u3_n106 ) , .ZN( u0_u7_u3_n119 ) , .C2( u0_u7_u3_n128 ) , .C1( u0_u7_u3_n167 ) , .A( u0_u7_u3_n181 ) );
  AOI221_X1 u0_u7_u3_U12 (.C1( u0_u7_u3_n105 ) , .ZN( u0_u7_u3_n106 ) , .A( u0_u7_u3_n131 ) , .B2( u0_u7_u3_n132 ) , .C2( u0_u7_u3_n133 ) , .B1( u0_u7_u3_n169 ) );
  INV_X1 u0_u7_u3_U13 (.ZN( u0_u7_u3_n181 ) , .A( u0_u7_u3_n98 ) );
  NAND2_X1 u0_u7_u3_U14 (.ZN( u0_u7_u3_n105 ) , .A2( u0_u7_u3_n130 ) , .A1( u0_u7_u3_n155 ) );
  AOI22_X1 u0_u7_u3_U15 (.B1( u0_u7_u3_n115 ) , .A2( u0_u7_u3_n116 ) , .ZN( u0_u7_u3_n123 ) , .B2( u0_u7_u3_n133 ) , .A1( u0_u7_u3_n169 ) );
  NAND2_X1 u0_u7_u3_U16 (.ZN( u0_u7_u3_n116 ) , .A2( u0_u7_u3_n151 ) , .A1( u0_u7_u3_n182 ) );
  NOR2_X1 u0_u7_u3_U17 (.ZN( u0_u7_u3_n126 ) , .A2( u0_u7_u3_n150 ) , .A1( u0_u7_u3_n164 ) );
  AOI21_X1 u0_u7_u3_U18 (.ZN( u0_u7_u3_n112 ) , .B2( u0_u7_u3_n146 ) , .B1( u0_u7_u3_n155 ) , .A( u0_u7_u3_n167 ) );
  NAND2_X1 u0_u7_u3_U19 (.A1( u0_u7_u3_n135 ) , .ZN( u0_u7_u3_n142 ) , .A2( u0_u7_u3_n164 ) );
  NAND2_X1 u0_u7_u3_U20 (.ZN( u0_u7_u3_n132 ) , .A2( u0_u7_u3_n152 ) , .A1( u0_u7_u3_n156 ) );
  AND2_X1 u0_u7_u3_U21 (.A2( u0_u7_u3_n113 ) , .A1( u0_u7_u3_n114 ) , .ZN( u0_u7_u3_n151 ) );
  INV_X1 u0_u7_u3_U22 (.A( u0_u7_u3_n133 ) , .ZN( u0_u7_u3_n165 ) );
  INV_X1 u0_u7_u3_U23 (.A( u0_u7_u3_n135 ) , .ZN( u0_u7_u3_n170 ) );
  NAND2_X1 u0_u7_u3_U24 (.A1( u0_u7_u3_n107 ) , .A2( u0_u7_u3_n108 ) , .ZN( u0_u7_u3_n140 ) );
  NAND2_X1 u0_u7_u3_U25 (.ZN( u0_u7_u3_n117 ) , .A1( u0_u7_u3_n124 ) , .A2( u0_u7_u3_n148 ) );
  NAND2_X1 u0_u7_u3_U26 (.ZN( u0_u7_u3_n143 ) , .A1( u0_u7_u3_n165 ) , .A2( u0_u7_u3_n167 ) );
  INV_X1 u0_u7_u3_U27 (.A( u0_u7_u3_n130 ) , .ZN( u0_u7_u3_n177 ) );
  INV_X1 u0_u7_u3_U28 (.A( u0_u7_u3_n128 ) , .ZN( u0_u7_u3_n176 ) );
  INV_X1 u0_u7_u3_U29 (.A( u0_u7_u3_n155 ) , .ZN( u0_u7_u3_n174 ) );
  INV_X1 u0_u7_u3_U3 (.A( u0_u7_u3_n129 ) , .ZN( u0_u7_u3_n183 ) );
  INV_X1 u0_u7_u3_U30 (.A( u0_u7_u3_n139 ) , .ZN( u0_u7_u3_n185 ) );
  NOR2_X1 u0_u7_u3_U31 (.ZN( u0_u7_u3_n135 ) , .A2( u0_u7_u3_n141 ) , .A1( u0_u7_u3_n169 ) );
  OAI222_X1 u0_u7_u3_U32 (.C2( u0_u7_u3_n107 ) , .A2( u0_u7_u3_n108 ) , .B1( u0_u7_u3_n135 ) , .ZN( u0_u7_u3_n138 ) , .B2( u0_u7_u3_n146 ) , .C1( u0_u7_u3_n154 ) , .A1( u0_u7_u3_n164 ) );
  NOR4_X1 u0_u7_u3_U33 (.A4( u0_u7_u3_n157 ) , .A3( u0_u7_u3_n158 ) , .A2( u0_u7_u3_n159 ) , .A1( u0_u7_u3_n160 ) , .ZN( u0_u7_u3_n161 ) );
  AOI21_X1 u0_u7_u3_U34 (.B2( u0_u7_u3_n152 ) , .B1( u0_u7_u3_n153 ) , .ZN( u0_u7_u3_n158 ) , .A( u0_u7_u3_n164 ) );
  AOI21_X1 u0_u7_u3_U35 (.A( u0_u7_u3_n154 ) , .B2( u0_u7_u3_n155 ) , .B1( u0_u7_u3_n156 ) , .ZN( u0_u7_u3_n157 ) );
  AOI21_X1 u0_u7_u3_U36 (.A( u0_u7_u3_n149 ) , .B2( u0_u7_u3_n150 ) , .B1( u0_u7_u3_n151 ) , .ZN( u0_u7_u3_n159 ) );
  AOI211_X1 u0_u7_u3_U37 (.ZN( u0_u7_u3_n109 ) , .A( u0_u7_u3_n119 ) , .C2( u0_u7_u3_n129 ) , .B( u0_u7_u3_n138 ) , .C1( u0_u7_u3_n141 ) );
  AOI211_X1 u0_u7_u3_U38 (.B( u0_u7_u3_n119 ) , .A( u0_u7_u3_n120 ) , .C2( u0_u7_u3_n121 ) , .ZN( u0_u7_u3_n122 ) , .C1( u0_u7_u3_n179 ) );
  INV_X1 u0_u7_u3_U39 (.A( u0_u7_u3_n156 ) , .ZN( u0_u7_u3_n179 ) );
  INV_X1 u0_u7_u3_U4 (.A( u0_u7_u3_n140 ) , .ZN( u0_u7_u3_n182 ) );
  OAI22_X1 u0_u7_u3_U40 (.B1( u0_u7_u3_n118 ) , .ZN( u0_u7_u3_n120 ) , .A1( u0_u7_u3_n135 ) , .B2( u0_u7_u3_n154 ) , .A2( u0_u7_u3_n178 ) );
  AND3_X1 u0_u7_u3_U41 (.ZN( u0_u7_u3_n118 ) , .A2( u0_u7_u3_n124 ) , .A1( u0_u7_u3_n144 ) , .A3( u0_u7_u3_n152 ) );
  INV_X1 u0_u7_u3_U42 (.A( u0_u7_u3_n121 ) , .ZN( u0_u7_u3_n164 ) );
  NAND2_X1 u0_u7_u3_U43 (.ZN( u0_u7_u3_n133 ) , .A1( u0_u7_u3_n154 ) , .A2( u0_u7_u3_n164 ) );
  OAI211_X1 u0_u7_u3_U44 (.B( u0_u7_u3_n127 ) , .ZN( u0_u7_u3_n139 ) , .C1( u0_u7_u3_n150 ) , .C2( u0_u7_u3_n154 ) , .A( u0_u7_u3_n184 ) );
  INV_X1 u0_u7_u3_U45 (.A( u0_u7_u3_n125 ) , .ZN( u0_u7_u3_n184 ) );
  AOI221_X1 u0_u7_u3_U46 (.A( u0_u7_u3_n126 ) , .ZN( u0_u7_u3_n127 ) , .C2( u0_u7_u3_n132 ) , .C1( u0_u7_u3_n169 ) , .B2( u0_u7_u3_n170 ) , .B1( u0_u7_u3_n174 ) );
  OAI22_X1 u0_u7_u3_U47 (.A1( u0_u7_u3_n124 ) , .ZN( u0_u7_u3_n125 ) , .B2( u0_u7_u3_n145 ) , .A2( u0_u7_u3_n165 ) , .B1( u0_u7_u3_n167 ) );
  NOR2_X1 u0_u7_u3_U48 (.A1( u0_u7_u3_n113 ) , .ZN( u0_u7_u3_n131 ) , .A2( u0_u7_u3_n154 ) );
  NAND2_X1 u0_u7_u3_U49 (.A1( u0_u7_u3_n103 ) , .ZN( u0_u7_u3_n150 ) , .A2( u0_u7_u3_n99 ) );
  INV_X1 u0_u7_u3_U5 (.A( u0_u7_u3_n117 ) , .ZN( u0_u7_u3_n178 ) );
  NAND2_X1 u0_u7_u3_U50 (.A2( u0_u7_u3_n102 ) , .ZN( u0_u7_u3_n155 ) , .A1( u0_u7_u3_n97 ) );
  INV_X1 u0_u7_u3_U51 (.A( u0_u7_u3_n141 ) , .ZN( u0_u7_u3_n167 ) );
  AOI21_X1 u0_u7_u3_U52 (.B2( u0_u7_u3_n114 ) , .B1( u0_u7_u3_n146 ) , .A( u0_u7_u3_n154 ) , .ZN( u0_u7_u3_n94 ) );
  AOI21_X1 u0_u7_u3_U53 (.ZN( u0_u7_u3_n110 ) , .B2( u0_u7_u3_n142 ) , .B1( u0_u7_u3_n186 ) , .A( u0_u7_u3_n95 ) );
  INV_X1 u0_u7_u3_U54 (.A( u0_u7_u3_n145 ) , .ZN( u0_u7_u3_n186 ) );
  AOI21_X1 u0_u7_u3_U55 (.B1( u0_u7_u3_n124 ) , .A( u0_u7_u3_n149 ) , .B2( u0_u7_u3_n155 ) , .ZN( u0_u7_u3_n95 ) );
  INV_X1 u0_u7_u3_U56 (.A( u0_u7_u3_n149 ) , .ZN( u0_u7_u3_n169 ) );
  NAND2_X1 u0_u7_u3_U57 (.ZN( u0_u7_u3_n124 ) , .A1( u0_u7_u3_n96 ) , .A2( u0_u7_u3_n97 ) );
  NAND2_X1 u0_u7_u3_U58 (.A2( u0_u7_u3_n100 ) , .ZN( u0_u7_u3_n146 ) , .A1( u0_u7_u3_n96 ) );
  NAND2_X1 u0_u7_u3_U59 (.A1( u0_u7_u3_n101 ) , .ZN( u0_u7_u3_n145 ) , .A2( u0_u7_u3_n99 ) );
  AOI221_X1 u0_u7_u3_U6 (.A( u0_u7_u3_n131 ) , .C2( u0_u7_u3_n132 ) , .C1( u0_u7_u3_n133 ) , .ZN( u0_u7_u3_n134 ) , .B1( u0_u7_u3_n143 ) , .B2( u0_u7_u3_n177 ) );
  NAND2_X1 u0_u7_u3_U60 (.A1( u0_u7_u3_n100 ) , .ZN( u0_u7_u3_n156 ) , .A2( u0_u7_u3_n99 ) );
  NAND2_X1 u0_u7_u3_U61 (.A2( u0_u7_u3_n101 ) , .A1( u0_u7_u3_n104 ) , .ZN( u0_u7_u3_n148 ) );
  NAND2_X1 u0_u7_u3_U62 (.A1( u0_u7_u3_n100 ) , .A2( u0_u7_u3_n102 ) , .ZN( u0_u7_u3_n128 ) );
  NAND2_X1 u0_u7_u3_U63 (.A2( u0_u7_u3_n101 ) , .A1( u0_u7_u3_n102 ) , .ZN( u0_u7_u3_n152 ) );
  NAND2_X1 u0_u7_u3_U64 (.A2( u0_u7_u3_n101 ) , .ZN( u0_u7_u3_n114 ) , .A1( u0_u7_u3_n96 ) );
  NAND2_X1 u0_u7_u3_U65 (.ZN( u0_u7_u3_n107 ) , .A1( u0_u7_u3_n97 ) , .A2( u0_u7_u3_n99 ) );
  NAND2_X1 u0_u7_u3_U66 (.A2( u0_u7_u3_n100 ) , .A1( u0_u7_u3_n104 ) , .ZN( u0_u7_u3_n113 ) );
  NAND2_X1 u0_u7_u3_U67 (.A1( u0_u7_u3_n104 ) , .ZN( u0_u7_u3_n153 ) , .A2( u0_u7_u3_n97 ) );
  NAND2_X1 u0_u7_u3_U68 (.A2( u0_u7_u3_n103 ) , .A1( u0_u7_u3_n104 ) , .ZN( u0_u7_u3_n130 ) );
  NAND2_X1 u0_u7_u3_U69 (.A2( u0_u7_u3_n103 ) , .ZN( u0_u7_u3_n144 ) , .A1( u0_u7_u3_n96 ) );
  OAI22_X1 u0_u7_u3_U7 (.B2( u0_u7_u3_n147 ) , .A2( u0_u7_u3_n148 ) , .ZN( u0_u7_u3_n160 ) , .B1( u0_u7_u3_n165 ) , .A1( u0_u7_u3_n168 ) );
  NAND2_X1 u0_u7_u3_U70 (.A1( u0_u7_u3_n102 ) , .A2( u0_u7_u3_n103 ) , .ZN( u0_u7_u3_n108 ) );
  NOR2_X1 u0_u7_u3_U71 (.A2( u0_u7_X_19 ) , .A1( u0_u7_X_20 ) , .ZN( u0_u7_u3_n99 ) );
  NOR2_X1 u0_u7_u3_U72 (.A2( u0_u7_X_21 ) , .A1( u0_u7_X_24 ) , .ZN( u0_u7_u3_n103 ) );
  NOR2_X1 u0_u7_u3_U73 (.A2( u0_u7_X_24 ) , .A1( u0_u7_u3_n171 ) , .ZN( u0_u7_u3_n97 ) );
  NOR2_X1 u0_u7_u3_U74 (.A2( u0_u7_X_23 ) , .ZN( u0_u7_u3_n141 ) , .A1( u0_u7_u3_n166 ) );
  NOR2_X1 u0_u7_u3_U75 (.A2( u0_u7_X_19 ) , .A1( u0_u7_u3_n172 ) , .ZN( u0_u7_u3_n96 ) );
  NAND2_X1 u0_u7_u3_U76 (.A1( u0_u7_X_22 ) , .A2( u0_u7_X_23 ) , .ZN( u0_u7_u3_n154 ) );
  NAND2_X1 u0_u7_u3_U77 (.A1( u0_u7_X_23 ) , .ZN( u0_u7_u3_n149 ) , .A2( u0_u7_u3_n166 ) );
  NOR2_X1 u0_u7_u3_U78 (.A2( u0_u7_X_22 ) , .A1( u0_u7_X_23 ) , .ZN( u0_u7_u3_n121 ) );
  AND2_X1 u0_u7_u3_U79 (.A1( u0_u7_X_24 ) , .ZN( u0_u7_u3_n101 ) , .A2( u0_u7_u3_n171 ) );
  AND3_X1 u0_u7_u3_U8 (.A3( u0_u7_u3_n144 ) , .A2( u0_u7_u3_n145 ) , .A1( u0_u7_u3_n146 ) , .ZN( u0_u7_u3_n147 ) );
  AND2_X1 u0_u7_u3_U80 (.A1( u0_u7_X_19 ) , .ZN( u0_u7_u3_n102 ) , .A2( u0_u7_u3_n172 ) );
  AND2_X1 u0_u7_u3_U81 (.A1( u0_u7_X_21 ) , .A2( u0_u7_X_24 ) , .ZN( u0_u7_u3_n100 ) );
  AND2_X1 u0_u7_u3_U82 (.A2( u0_u7_X_19 ) , .A1( u0_u7_X_20 ) , .ZN( u0_u7_u3_n104 ) );
  INV_X1 u0_u7_u3_U83 (.A( u0_u7_X_22 ) , .ZN( u0_u7_u3_n166 ) );
  INV_X1 u0_u7_u3_U84 (.A( u0_u7_X_21 ) , .ZN( u0_u7_u3_n171 ) );
  INV_X1 u0_u7_u3_U85 (.A( u0_u7_X_20 ) , .ZN( u0_u7_u3_n172 ) );
  OR4_X1 u0_u7_u3_U86 (.ZN( u0_out7_10 ) , .A4( u0_u7_u3_n136 ) , .A3( u0_u7_u3_n137 ) , .A1( u0_u7_u3_n138 ) , .A2( u0_u7_u3_n139 ) );
  OAI222_X1 u0_u7_u3_U87 (.C1( u0_u7_u3_n128 ) , .ZN( u0_u7_u3_n137 ) , .B1( u0_u7_u3_n148 ) , .A2( u0_u7_u3_n150 ) , .B2( u0_u7_u3_n154 ) , .C2( u0_u7_u3_n164 ) , .A1( u0_u7_u3_n167 ) );
  OAI221_X1 u0_u7_u3_U88 (.A( u0_u7_u3_n134 ) , .B2( u0_u7_u3_n135 ) , .ZN( u0_u7_u3_n136 ) , .C1( u0_u7_u3_n149 ) , .B1( u0_u7_u3_n151 ) , .C2( u0_u7_u3_n183 ) );
  NAND4_X1 u0_u7_u3_U89 (.ZN( u0_out7_26 ) , .A4( u0_u7_u3_n109 ) , .A3( u0_u7_u3_n110 ) , .A2( u0_u7_u3_n111 ) , .A1( u0_u7_u3_n173 ) );
  INV_X1 u0_u7_u3_U9 (.A( u0_u7_u3_n143 ) , .ZN( u0_u7_u3_n168 ) );
  INV_X1 u0_u7_u3_U90 (.ZN( u0_u7_u3_n173 ) , .A( u0_u7_u3_n94 ) );
  OAI21_X1 u0_u7_u3_U91 (.ZN( u0_u7_u3_n111 ) , .B2( u0_u7_u3_n117 ) , .A( u0_u7_u3_n133 ) , .B1( u0_u7_u3_n176 ) );
  NAND4_X1 u0_u7_u3_U92 (.ZN( u0_out7_20 ) , .A4( u0_u7_u3_n122 ) , .A3( u0_u7_u3_n123 ) , .A1( u0_u7_u3_n175 ) , .A2( u0_u7_u3_n180 ) );
  INV_X1 u0_u7_u3_U93 (.A( u0_u7_u3_n126 ) , .ZN( u0_u7_u3_n180 ) );
  INV_X1 u0_u7_u3_U94 (.A( u0_u7_u3_n112 ) , .ZN( u0_u7_u3_n175 ) );
  NAND4_X1 u0_u7_u3_U95 (.ZN( u0_out7_1 ) , .A4( u0_u7_u3_n161 ) , .A3( u0_u7_u3_n162 ) , .A2( u0_u7_u3_n163 ) , .A1( u0_u7_u3_n185 ) );
  NAND2_X1 u0_u7_u3_U96 (.ZN( u0_u7_u3_n163 ) , .A2( u0_u7_u3_n170 ) , .A1( u0_u7_u3_n176 ) );
  AOI22_X1 u0_u7_u3_U97 (.B2( u0_u7_u3_n140 ) , .B1( u0_u7_u3_n141 ) , .A2( u0_u7_u3_n142 ) , .ZN( u0_u7_u3_n162 ) , .A1( u0_u7_u3_n177 ) );
  NAND3_X1 u0_u7_u3_U98 (.A1( u0_u7_u3_n114 ) , .ZN( u0_u7_u3_n115 ) , .A2( u0_u7_u3_n145 ) , .A3( u0_u7_u3_n153 ) );
  NAND3_X1 u0_u7_u3_U99 (.ZN( u0_u7_u3_n129 ) , .A2( u0_u7_u3_n144 ) , .A1( u0_u7_u3_n153 ) , .A3( u0_u7_u3_n182 ) );
  XOR2_X1 u0_u9_U1 (.B( u0_K10_9 ) , .A( u0_R8_6 ) , .Z( u0_u9_X_9 ) );
  XOR2_X1 u0_u9_U13 (.B( u0_K10_42 ) , .A( u0_R8_29 ) , .Z( u0_u9_X_42 ) );
  XOR2_X1 u0_u9_U14 (.B( u0_K10_41 ) , .A( u0_R8_28 ) , .Z( u0_u9_X_41 ) );
  XOR2_X1 u0_u9_U15 (.B( u0_K10_40 ) , .A( u0_R8_27 ) , .Z( u0_u9_X_40 ) );
  XOR2_X1 u0_u9_U16 (.B( u0_K10_3 ) , .A( u0_R8_2 ) , .Z( u0_u9_X_3 ) );
  XOR2_X1 u0_u9_U17 (.B( u0_K10_39 ) , .A( u0_R8_26 ) , .Z( u0_u9_X_39 ) );
  XOR2_X1 u0_u9_U18 (.B( u0_K10_38 ) , .A( u0_R8_25 ) , .Z( u0_u9_X_38 ) );
  XOR2_X1 u0_u9_U19 (.B( u0_K10_37 ) , .A( u0_R8_24 ) , .Z( u0_u9_X_37 ) );
  XOR2_X1 u0_u9_U2 (.B( u0_K10_8 ) , .A( u0_R8_5 ) , .Z( u0_u9_X_8 ) );
  XOR2_X1 u0_u9_U27 (.B( u0_K10_2 ) , .A( u0_R8_1 ) , .Z( u0_u9_X_2 ) );
  XOR2_X1 u0_u9_U3 (.B( u0_K10_7 ) , .A( u0_R8_4 ) , .Z( u0_u9_X_7 ) );
  XOR2_X1 u0_u9_U38 (.B( u0_K10_1 ) , .A( u0_R8_32 ) , .Z( u0_u9_X_1 ) );
  XOR2_X1 u0_u9_U4 (.B( u0_K10_6 ) , .A( u0_R8_5 ) , .Z( u0_u9_X_6 ) );
  XOR2_X1 u0_u9_U40 (.B( u0_K10_18 ) , .A( u0_R8_13 ) , .Z( u0_u9_X_18 ) );
  XOR2_X1 u0_u9_U41 (.B( u0_K10_17 ) , .A( u0_R8_12 ) , .Z( u0_u9_X_17 ) );
  XOR2_X1 u0_u9_U42 (.B( u0_K10_16 ) , .A( u0_R8_11 ) , .Z( u0_u9_X_16 ) );
  XOR2_X1 u0_u9_U43 (.B( u0_K10_15 ) , .A( u0_R8_10 ) , .Z( u0_u9_X_15 ) );
  XOR2_X1 u0_u9_U44 (.B( u0_K10_14 ) , .A( u0_R8_9 ) , .Z( u0_u9_X_14 ) );
  XOR2_X1 u0_u9_U45 (.B( u0_K10_13 ) , .A( u0_R8_8 ) , .Z( u0_u9_X_13 ) );
  XOR2_X1 u0_u9_U46 (.B( u0_K10_12 ) , .A( u0_R8_9 ) , .Z( u0_u9_X_12 ) );
  XOR2_X1 u0_u9_U47 (.B( u0_K10_11 ) , .A( u0_R8_8 ) , .Z( u0_u9_X_11 ) );
  XOR2_X1 u0_u9_U48 (.B( u0_K10_10 ) , .A( u0_R8_7 ) , .Z( u0_u9_X_10 ) );
  XOR2_X1 u0_u9_U5 (.B( u0_K10_5 ) , .A( u0_R8_4 ) , .Z( u0_u9_X_5 ) );
  XOR2_X1 u0_u9_U6 (.B( u0_K10_4 ) , .A( u0_R8_3 ) , .Z( u0_u9_X_4 ) );
  AND3_X1 u0_u9_u0_U10 (.A2( u0_u9_u0_n112 ) , .ZN( u0_u9_u0_n127 ) , .A3( u0_u9_u0_n130 ) , .A1( u0_u9_u0_n148 ) );
  NAND2_X1 u0_u9_u0_U11 (.ZN( u0_u9_u0_n113 ) , .A1( u0_u9_u0_n139 ) , .A2( u0_u9_u0_n149 ) );
  AND2_X1 u0_u9_u0_U12 (.ZN( u0_u9_u0_n107 ) , .A1( u0_u9_u0_n130 ) , .A2( u0_u9_u0_n140 ) );
  AND2_X1 u0_u9_u0_U13 (.A2( u0_u9_u0_n129 ) , .A1( u0_u9_u0_n130 ) , .ZN( u0_u9_u0_n151 ) );
  AND2_X1 u0_u9_u0_U14 (.A1( u0_u9_u0_n108 ) , .A2( u0_u9_u0_n125 ) , .ZN( u0_u9_u0_n145 ) );
  INV_X1 u0_u9_u0_U15 (.A( u0_u9_u0_n143 ) , .ZN( u0_u9_u0_n173 ) );
  NOR2_X1 u0_u9_u0_U16 (.A2( u0_u9_u0_n136 ) , .ZN( u0_u9_u0_n147 ) , .A1( u0_u9_u0_n160 ) );
  AOI21_X1 u0_u9_u0_U17 (.B1( u0_u9_u0_n103 ) , .ZN( u0_u9_u0_n132 ) , .A( u0_u9_u0_n165 ) , .B2( u0_u9_u0_n93 ) );
  INV_X1 u0_u9_u0_U18 (.A( u0_u9_u0_n142 ) , .ZN( u0_u9_u0_n165 ) );
  OAI221_X1 u0_u9_u0_U19 (.C1( u0_u9_u0_n121 ) , .ZN( u0_u9_u0_n122 ) , .B2( u0_u9_u0_n127 ) , .A( u0_u9_u0_n143 ) , .B1( u0_u9_u0_n144 ) , .C2( u0_u9_u0_n147 ) );
  OAI22_X1 u0_u9_u0_U20 (.B1( u0_u9_u0_n131 ) , .A1( u0_u9_u0_n144 ) , .B2( u0_u9_u0_n147 ) , .A2( u0_u9_u0_n90 ) , .ZN( u0_u9_u0_n91 ) );
  AND3_X1 u0_u9_u0_U21 (.A3( u0_u9_u0_n121 ) , .A2( u0_u9_u0_n125 ) , .A1( u0_u9_u0_n148 ) , .ZN( u0_u9_u0_n90 ) );
  OAI22_X1 u0_u9_u0_U22 (.B1( u0_u9_u0_n125 ) , .ZN( u0_u9_u0_n126 ) , .A1( u0_u9_u0_n138 ) , .A2( u0_u9_u0_n146 ) , .B2( u0_u9_u0_n147 ) );
  NOR2_X1 u0_u9_u0_U23 (.A1( u0_u9_u0_n163 ) , .A2( u0_u9_u0_n164 ) , .ZN( u0_u9_u0_n95 ) );
  INV_X1 u0_u9_u0_U24 (.A( u0_u9_u0_n136 ) , .ZN( u0_u9_u0_n161 ) );
  NOR2_X1 u0_u9_u0_U25 (.A1( u0_u9_u0_n120 ) , .ZN( u0_u9_u0_n143 ) , .A2( u0_u9_u0_n167 ) );
  OAI221_X1 u0_u9_u0_U26 (.C1( u0_u9_u0_n112 ) , .ZN( u0_u9_u0_n120 ) , .B1( u0_u9_u0_n138 ) , .B2( u0_u9_u0_n141 ) , .C2( u0_u9_u0_n147 ) , .A( u0_u9_u0_n172 ) );
  AOI211_X1 u0_u9_u0_U27 (.B( u0_u9_u0_n115 ) , .A( u0_u9_u0_n116 ) , .C2( u0_u9_u0_n117 ) , .C1( u0_u9_u0_n118 ) , .ZN( u0_u9_u0_n119 ) );
  NAND2_X1 u0_u9_u0_U28 (.A1( u0_u9_u0_n101 ) , .A2( u0_u9_u0_n102 ) , .ZN( u0_u9_u0_n150 ) );
  AOI22_X1 u0_u9_u0_U29 (.B2( u0_u9_u0_n109 ) , .A2( u0_u9_u0_n110 ) , .ZN( u0_u9_u0_n111 ) , .B1( u0_u9_u0_n118 ) , .A1( u0_u9_u0_n160 ) );
  INV_X1 u0_u9_u0_U3 (.A( u0_u9_u0_n113 ) , .ZN( u0_u9_u0_n166 ) );
  INV_X1 u0_u9_u0_U30 (.A( u0_u9_u0_n118 ) , .ZN( u0_u9_u0_n158 ) );
  NAND2_X1 u0_u9_u0_U31 (.A2( u0_u9_u0_n100 ) , .A1( u0_u9_u0_n101 ) , .ZN( u0_u9_u0_n139 ) );
  NAND2_X1 u0_u9_u0_U32 (.A2( u0_u9_u0_n100 ) , .ZN( u0_u9_u0_n131 ) , .A1( u0_u9_u0_n92 ) );
  NAND2_X1 u0_u9_u0_U33 (.ZN( u0_u9_u0_n108 ) , .A1( u0_u9_u0_n92 ) , .A2( u0_u9_u0_n94 ) );
  AOI21_X1 u0_u9_u0_U34 (.ZN( u0_u9_u0_n104 ) , .B1( u0_u9_u0_n107 ) , .B2( u0_u9_u0_n141 ) , .A( u0_u9_u0_n144 ) );
  AOI21_X1 u0_u9_u0_U35 (.B1( u0_u9_u0_n127 ) , .B2( u0_u9_u0_n129 ) , .A( u0_u9_u0_n138 ) , .ZN( u0_u9_u0_n96 ) );
  NAND2_X1 u0_u9_u0_U36 (.A2( u0_u9_u0_n102 ) , .ZN( u0_u9_u0_n114 ) , .A1( u0_u9_u0_n92 ) );
  AOI21_X1 u0_u9_u0_U37 (.ZN( u0_u9_u0_n116 ) , .B2( u0_u9_u0_n142 ) , .A( u0_u9_u0_n144 ) , .B1( u0_u9_u0_n166 ) );
  NAND2_X1 u0_u9_u0_U38 (.A1( u0_u9_u0_n101 ) , .ZN( u0_u9_u0_n130 ) , .A2( u0_u9_u0_n94 ) );
  NAND2_X1 u0_u9_u0_U39 (.A1( u0_u9_u0_n100 ) , .A2( u0_u9_u0_n103 ) , .ZN( u0_u9_u0_n125 ) );
  AOI21_X1 u0_u9_u0_U4 (.B1( u0_u9_u0_n114 ) , .ZN( u0_u9_u0_n115 ) , .B2( u0_u9_u0_n129 ) , .A( u0_u9_u0_n161 ) );
  NAND2_X1 u0_u9_u0_U40 (.A2( u0_u9_u0_n103 ) , .ZN( u0_u9_u0_n140 ) , .A1( u0_u9_u0_n94 ) );
  INV_X1 u0_u9_u0_U41 (.A( u0_u9_u0_n138 ) , .ZN( u0_u9_u0_n160 ) );
  NAND2_X1 u0_u9_u0_U42 (.A2( u0_u9_u0_n102 ) , .A1( u0_u9_u0_n103 ) , .ZN( u0_u9_u0_n149 ) );
  NAND2_X1 u0_u9_u0_U43 (.A2( u0_u9_u0_n101 ) , .ZN( u0_u9_u0_n121 ) , .A1( u0_u9_u0_n93 ) );
  NAND2_X1 u0_u9_u0_U44 (.ZN( u0_u9_u0_n112 ) , .A2( u0_u9_u0_n92 ) , .A1( u0_u9_u0_n93 ) );
  INV_X1 u0_u9_u0_U45 (.ZN( u0_u9_u0_n172 ) , .A( u0_u9_u0_n88 ) );
  OAI222_X1 u0_u9_u0_U46 (.C1( u0_u9_u0_n108 ) , .A1( u0_u9_u0_n125 ) , .B2( u0_u9_u0_n128 ) , .B1( u0_u9_u0_n144 ) , .A2( u0_u9_u0_n158 ) , .C2( u0_u9_u0_n161 ) , .ZN( u0_u9_u0_n88 ) );
  OR3_X1 u0_u9_u0_U47 (.A3( u0_u9_u0_n152 ) , .A2( u0_u9_u0_n153 ) , .A1( u0_u9_u0_n154 ) , .ZN( u0_u9_u0_n155 ) );
  AOI21_X1 u0_u9_u0_U48 (.A( u0_u9_u0_n144 ) , .B2( u0_u9_u0_n145 ) , .B1( u0_u9_u0_n146 ) , .ZN( u0_u9_u0_n154 ) );
  AOI21_X1 u0_u9_u0_U49 (.B2( u0_u9_u0_n150 ) , .B1( u0_u9_u0_n151 ) , .ZN( u0_u9_u0_n152 ) , .A( u0_u9_u0_n158 ) );
  AOI21_X1 u0_u9_u0_U5 (.B2( u0_u9_u0_n131 ) , .ZN( u0_u9_u0_n134 ) , .B1( u0_u9_u0_n151 ) , .A( u0_u9_u0_n158 ) );
  AOI21_X1 u0_u9_u0_U50 (.A( u0_u9_u0_n147 ) , .B2( u0_u9_u0_n148 ) , .B1( u0_u9_u0_n149 ) , .ZN( u0_u9_u0_n153 ) );
  INV_X1 u0_u9_u0_U51 (.ZN( u0_u9_u0_n171 ) , .A( u0_u9_u0_n99 ) );
  OAI211_X1 u0_u9_u0_U52 (.C2( u0_u9_u0_n140 ) , .C1( u0_u9_u0_n161 ) , .A( u0_u9_u0_n169 ) , .B( u0_u9_u0_n98 ) , .ZN( u0_u9_u0_n99 ) );
  INV_X1 u0_u9_u0_U53 (.ZN( u0_u9_u0_n169 ) , .A( u0_u9_u0_n91 ) );
  AOI211_X1 u0_u9_u0_U54 (.C1( u0_u9_u0_n118 ) , .A( u0_u9_u0_n123 ) , .B( u0_u9_u0_n96 ) , .C2( u0_u9_u0_n97 ) , .ZN( u0_u9_u0_n98 ) );
  NOR2_X1 u0_u9_u0_U55 (.A2( u0_u9_X_2 ) , .ZN( u0_u9_u0_n103 ) , .A1( u0_u9_u0_n164 ) );
  NOR2_X1 u0_u9_u0_U56 (.A2( u0_u9_X_4 ) , .A1( u0_u9_X_5 ) , .ZN( u0_u9_u0_n118 ) );
  NOR2_X1 u0_u9_u0_U57 (.A2( u0_u9_X_3 ) , .A1( u0_u9_X_6 ) , .ZN( u0_u9_u0_n94 ) );
  NOR2_X1 u0_u9_u0_U58 (.A2( u0_u9_X_6 ) , .ZN( u0_u9_u0_n100 ) , .A1( u0_u9_u0_n162 ) );
  NAND2_X1 u0_u9_u0_U59 (.A2( u0_u9_X_4 ) , .A1( u0_u9_X_5 ) , .ZN( u0_u9_u0_n144 ) );
  NOR2_X1 u0_u9_u0_U6 (.A1( u0_u9_u0_n108 ) , .ZN( u0_u9_u0_n123 ) , .A2( u0_u9_u0_n158 ) );
  NOR2_X1 u0_u9_u0_U60 (.A2( u0_u9_X_5 ) , .ZN( u0_u9_u0_n136 ) , .A1( u0_u9_u0_n159 ) );
  NAND2_X1 u0_u9_u0_U61 (.A1( u0_u9_X_5 ) , .ZN( u0_u9_u0_n138 ) , .A2( u0_u9_u0_n159 ) );
  AND2_X1 u0_u9_u0_U62 (.A2( u0_u9_X_3 ) , .A1( u0_u9_X_6 ) , .ZN( u0_u9_u0_n102 ) );
  AND2_X1 u0_u9_u0_U63 (.A1( u0_u9_X_6 ) , .A2( u0_u9_u0_n162 ) , .ZN( u0_u9_u0_n93 ) );
  INV_X1 u0_u9_u0_U64 (.A( u0_u9_X_4 ) , .ZN( u0_u9_u0_n159 ) );
  INV_X1 u0_u9_u0_U65 (.A( u0_u9_X_3 ) , .ZN( u0_u9_u0_n162 ) );
  INV_X1 u0_u9_u0_U66 (.A( u0_u9_X_2 ) , .ZN( u0_u9_u0_n163 ) );
  INV_X1 u0_u9_u0_U67 (.A( u0_u9_u0_n126 ) , .ZN( u0_u9_u0_n168 ) );
  AOI211_X1 u0_u9_u0_U68 (.B( u0_u9_u0_n133 ) , .A( u0_u9_u0_n134 ) , .C2( u0_u9_u0_n135 ) , .C1( u0_u9_u0_n136 ) , .ZN( u0_u9_u0_n137 ) );
  INV_X1 u0_u9_u0_U69 (.ZN( u0_u9_u0_n174 ) , .A( u0_u9_u0_n89 ) );
  OAI21_X1 u0_u9_u0_U7 (.B1( u0_u9_u0_n150 ) , .B2( u0_u9_u0_n158 ) , .A( u0_u9_u0_n172 ) , .ZN( u0_u9_u0_n89 ) );
  AOI211_X1 u0_u9_u0_U70 (.B( u0_u9_u0_n104 ) , .A( u0_u9_u0_n105 ) , .ZN( u0_u9_u0_n106 ) , .C2( u0_u9_u0_n113 ) , .C1( u0_u9_u0_n160 ) );
  OR4_X1 u0_u9_u0_U71 (.ZN( u0_out9_17 ) , .A4( u0_u9_u0_n122 ) , .A2( u0_u9_u0_n123 ) , .A1( u0_u9_u0_n124 ) , .A3( u0_u9_u0_n170 ) );
  AOI21_X1 u0_u9_u0_U72 (.B2( u0_u9_u0_n107 ) , .ZN( u0_u9_u0_n124 ) , .B1( u0_u9_u0_n128 ) , .A( u0_u9_u0_n161 ) );
  INV_X1 u0_u9_u0_U73 (.A( u0_u9_u0_n111 ) , .ZN( u0_u9_u0_n170 ) );
  OR4_X1 u0_u9_u0_U74 (.ZN( u0_out9_31 ) , .A4( u0_u9_u0_n155 ) , .A2( u0_u9_u0_n156 ) , .A1( u0_u9_u0_n157 ) , .A3( u0_u9_u0_n173 ) );
  AOI21_X1 u0_u9_u0_U75 (.A( u0_u9_u0_n138 ) , .B2( u0_u9_u0_n139 ) , .B1( u0_u9_u0_n140 ) , .ZN( u0_u9_u0_n157 ) );
  AOI21_X1 u0_u9_u0_U76 (.B2( u0_u9_u0_n141 ) , .B1( u0_u9_u0_n142 ) , .ZN( u0_u9_u0_n156 ) , .A( u0_u9_u0_n161 ) );
  AOI21_X1 u0_u9_u0_U77 (.B1( u0_u9_u0_n132 ) , .ZN( u0_u9_u0_n133 ) , .A( u0_u9_u0_n144 ) , .B2( u0_u9_u0_n166 ) );
  OAI22_X1 u0_u9_u0_U78 (.ZN( u0_u9_u0_n105 ) , .A2( u0_u9_u0_n132 ) , .B1( u0_u9_u0_n146 ) , .A1( u0_u9_u0_n147 ) , .B2( u0_u9_u0_n161 ) );
  NAND2_X1 u0_u9_u0_U79 (.ZN( u0_u9_u0_n110 ) , .A2( u0_u9_u0_n132 ) , .A1( u0_u9_u0_n145 ) );
  AND2_X1 u0_u9_u0_U8 (.A1( u0_u9_u0_n114 ) , .A2( u0_u9_u0_n121 ) , .ZN( u0_u9_u0_n146 ) );
  INV_X1 u0_u9_u0_U80 (.A( u0_u9_u0_n119 ) , .ZN( u0_u9_u0_n167 ) );
  NAND2_X1 u0_u9_u0_U81 (.ZN( u0_u9_u0_n148 ) , .A1( u0_u9_u0_n93 ) , .A2( u0_u9_u0_n95 ) );
  NAND2_X1 u0_u9_u0_U82 (.A1( u0_u9_u0_n100 ) , .ZN( u0_u9_u0_n129 ) , .A2( u0_u9_u0_n95 ) );
  NAND2_X1 u0_u9_u0_U83 (.A1( u0_u9_u0_n102 ) , .ZN( u0_u9_u0_n128 ) , .A2( u0_u9_u0_n95 ) );
  NOR2_X1 u0_u9_u0_U84 (.A2( u0_u9_X_1 ) , .A1( u0_u9_X_2 ) , .ZN( u0_u9_u0_n92 ) );
  NAND2_X1 u0_u9_u0_U85 (.ZN( u0_u9_u0_n142 ) , .A1( u0_u9_u0_n94 ) , .A2( u0_u9_u0_n95 ) );
  NOR2_X1 u0_u9_u0_U86 (.A2( u0_u9_X_1 ) , .ZN( u0_u9_u0_n101 ) , .A1( u0_u9_u0_n163 ) );
  INV_X1 u0_u9_u0_U87 (.A( u0_u9_X_1 ) , .ZN( u0_u9_u0_n164 ) );
  NAND3_X1 u0_u9_u0_U88 (.ZN( u0_out9_23 ) , .A3( u0_u9_u0_n137 ) , .A1( u0_u9_u0_n168 ) , .A2( u0_u9_u0_n171 ) );
  NAND3_X1 u0_u9_u0_U89 (.A3( u0_u9_u0_n127 ) , .A2( u0_u9_u0_n128 ) , .ZN( u0_u9_u0_n135 ) , .A1( u0_u9_u0_n150 ) );
  AND2_X1 u0_u9_u0_U9 (.A1( u0_u9_u0_n131 ) , .ZN( u0_u9_u0_n141 ) , .A2( u0_u9_u0_n150 ) );
  NAND3_X1 u0_u9_u0_U90 (.ZN( u0_u9_u0_n117 ) , .A3( u0_u9_u0_n132 ) , .A2( u0_u9_u0_n139 ) , .A1( u0_u9_u0_n148 ) );
  NAND3_X1 u0_u9_u0_U91 (.ZN( u0_u9_u0_n109 ) , .A2( u0_u9_u0_n114 ) , .A3( u0_u9_u0_n140 ) , .A1( u0_u9_u0_n149 ) );
  NAND3_X1 u0_u9_u0_U92 (.ZN( u0_out9_9 ) , .A3( u0_u9_u0_n106 ) , .A2( u0_u9_u0_n171 ) , .A1( u0_u9_u0_n174 ) );
  NAND3_X1 u0_u9_u0_U93 (.A2( u0_u9_u0_n128 ) , .A1( u0_u9_u0_n132 ) , .A3( u0_u9_u0_n146 ) , .ZN( u0_u9_u0_n97 ) );
  NOR2_X1 u0_u9_u1_U10 (.A1( u0_u9_u1_n112 ) , .A2( u0_u9_u1_n116 ) , .ZN( u0_u9_u1_n118 ) );
  NAND3_X1 u0_u9_u1_U100 (.ZN( u0_u9_u1_n113 ) , .A1( u0_u9_u1_n120 ) , .A3( u0_u9_u1_n133 ) , .A2( u0_u9_u1_n155 ) );
  OAI21_X1 u0_u9_u1_U11 (.ZN( u0_u9_u1_n101 ) , .B1( u0_u9_u1_n141 ) , .A( u0_u9_u1_n146 ) , .B2( u0_u9_u1_n183 ) );
  AOI21_X1 u0_u9_u1_U12 (.B2( u0_u9_u1_n155 ) , .B1( u0_u9_u1_n156 ) , .ZN( u0_u9_u1_n157 ) , .A( u0_u9_u1_n174 ) );
  NAND2_X1 u0_u9_u1_U13 (.ZN( u0_u9_u1_n140 ) , .A2( u0_u9_u1_n150 ) , .A1( u0_u9_u1_n155 ) );
  NAND2_X1 u0_u9_u1_U14 (.A1( u0_u9_u1_n131 ) , .ZN( u0_u9_u1_n147 ) , .A2( u0_u9_u1_n153 ) );
  INV_X1 u0_u9_u1_U15 (.A( u0_u9_u1_n139 ) , .ZN( u0_u9_u1_n174 ) );
  OR4_X1 u0_u9_u1_U16 (.A4( u0_u9_u1_n106 ) , .A3( u0_u9_u1_n107 ) , .ZN( u0_u9_u1_n108 ) , .A1( u0_u9_u1_n117 ) , .A2( u0_u9_u1_n184 ) );
  AOI21_X1 u0_u9_u1_U17 (.ZN( u0_u9_u1_n106 ) , .A( u0_u9_u1_n112 ) , .B1( u0_u9_u1_n154 ) , .B2( u0_u9_u1_n156 ) );
  AOI21_X1 u0_u9_u1_U18 (.ZN( u0_u9_u1_n107 ) , .B1( u0_u9_u1_n134 ) , .B2( u0_u9_u1_n149 ) , .A( u0_u9_u1_n174 ) );
  INV_X1 u0_u9_u1_U19 (.A( u0_u9_u1_n101 ) , .ZN( u0_u9_u1_n184 ) );
  INV_X1 u0_u9_u1_U20 (.A( u0_u9_u1_n112 ) , .ZN( u0_u9_u1_n171 ) );
  NAND2_X1 u0_u9_u1_U21 (.ZN( u0_u9_u1_n141 ) , .A1( u0_u9_u1_n153 ) , .A2( u0_u9_u1_n156 ) );
  AND2_X1 u0_u9_u1_U22 (.A1( u0_u9_u1_n123 ) , .ZN( u0_u9_u1_n134 ) , .A2( u0_u9_u1_n161 ) );
  NAND2_X1 u0_u9_u1_U23 (.A2( u0_u9_u1_n115 ) , .A1( u0_u9_u1_n116 ) , .ZN( u0_u9_u1_n148 ) );
  NAND2_X1 u0_u9_u1_U24 (.A2( u0_u9_u1_n133 ) , .A1( u0_u9_u1_n135 ) , .ZN( u0_u9_u1_n159 ) );
  NAND2_X1 u0_u9_u1_U25 (.A2( u0_u9_u1_n115 ) , .A1( u0_u9_u1_n120 ) , .ZN( u0_u9_u1_n132 ) );
  INV_X1 u0_u9_u1_U26 (.A( u0_u9_u1_n154 ) , .ZN( u0_u9_u1_n178 ) );
  INV_X1 u0_u9_u1_U27 (.A( u0_u9_u1_n151 ) , .ZN( u0_u9_u1_n183 ) );
  AND2_X1 u0_u9_u1_U28 (.A1( u0_u9_u1_n129 ) , .A2( u0_u9_u1_n133 ) , .ZN( u0_u9_u1_n149 ) );
  INV_X1 u0_u9_u1_U29 (.A( u0_u9_u1_n131 ) , .ZN( u0_u9_u1_n180 ) );
  INV_X1 u0_u9_u1_U3 (.A( u0_u9_u1_n159 ) , .ZN( u0_u9_u1_n182 ) );
  OAI221_X1 u0_u9_u1_U30 (.A( u0_u9_u1_n119 ) , .C2( u0_u9_u1_n129 ) , .ZN( u0_u9_u1_n138 ) , .B2( u0_u9_u1_n152 ) , .C1( u0_u9_u1_n174 ) , .B1( u0_u9_u1_n187 ) );
  INV_X1 u0_u9_u1_U31 (.A( u0_u9_u1_n148 ) , .ZN( u0_u9_u1_n187 ) );
  AOI211_X1 u0_u9_u1_U32 (.B( u0_u9_u1_n117 ) , .A( u0_u9_u1_n118 ) , .ZN( u0_u9_u1_n119 ) , .C2( u0_u9_u1_n146 ) , .C1( u0_u9_u1_n159 ) );
  NOR2_X1 u0_u9_u1_U33 (.A1( u0_u9_u1_n168 ) , .A2( u0_u9_u1_n176 ) , .ZN( u0_u9_u1_n98 ) );
  AOI211_X1 u0_u9_u1_U34 (.B( u0_u9_u1_n162 ) , .A( u0_u9_u1_n163 ) , .C2( u0_u9_u1_n164 ) , .ZN( u0_u9_u1_n165 ) , .C1( u0_u9_u1_n171 ) );
  AOI21_X1 u0_u9_u1_U35 (.A( u0_u9_u1_n160 ) , .B2( u0_u9_u1_n161 ) , .ZN( u0_u9_u1_n162 ) , .B1( u0_u9_u1_n182 ) );
  OR2_X1 u0_u9_u1_U36 (.A2( u0_u9_u1_n157 ) , .A1( u0_u9_u1_n158 ) , .ZN( u0_u9_u1_n163 ) );
  NAND2_X1 u0_u9_u1_U37 (.A1( u0_u9_u1_n128 ) , .ZN( u0_u9_u1_n146 ) , .A2( u0_u9_u1_n160 ) );
  NAND2_X1 u0_u9_u1_U38 (.A2( u0_u9_u1_n112 ) , .ZN( u0_u9_u1_n139 ) , .A1( u0_u9_u1_n152 ) );
  NAND2_X1 u0_u9_u1_U39 (.A1( u0_u9_u1_n105 ) , .ZN( u0_u9_u1_n156 ) , .A2( u0_u9_u1_n99 ) );
  AOI221_X1 u0_u9_u1_U4 (.A( u0_u9_u1_n138 ) , .C2( u0_u9_u1_n139 ) , .C1( u0_u9_u1_n140 ) , .B2( u0_u9_u1_n141 ) , .ZN( u0_u9_u1_n142 ) , .B1( u0_u9_u1_n175 ) );
  AOI221_X1 u0_u9_u1_U40 (.B1( u0_u9_u1_n140 ) , .ZN( u0_u9_u1_n167 ) , .B2( u0_u9_u1_n172 ) , .C2( u0_u9_u1_n175 ) , .C1( u0_u9_u1_n178 ) , .A( u0_u9_u1_n188 ) );
  INV_X1 u0_u9_u1_U41 (.ZN( u0_u9_u1_n188 ) , .A( u0_u9_u1_n97 ) );
  AOI211_X1 u0_u9_u1_U42 (.A( u0_u9_u1_n118 ) , .C1( u0_u9_u1_n132 ) , .C2( u0_u9_u1_n139 ) , .B( u0_u9_u1_n96 ) , .ZN( u0_u9_u1_n97 ) );
  AOI21_X1 u0_u9_u1_U43 (.B2( u0_u9_u1_n121 ) , .B1( u0_u9_u1_n135 ) , .A( u0_u9_u1_n152 ) , .ZN( u0_u9_u1_n96 ) );
  NOR2_X1 u0_u9_u1_U44 (.ZN( u0_u9_u1_n117 ) , .A1( u0_u9_u1_n121 ) , .A2( u0_u9_u1_n160 ) );
  OAI21_X1 u0_u9_u1_U45 (.B2( u0_u9_u1_n123 ) , .ZN( u0_u9_u1_n145 ) , .B1( u0_u9_u1_n160 ) , .A( u0_u9_u1_n185 ) );
  INV_X1 u0_u9_u1_U46 (.A( u0_u9_u1_n122 ) , .ZN( u0_u9_u1_n185 ) );
  AOI21_X1 u0_u9_u1_U47 (.B2( u0_u9_u1_n120 ) , .B1( u0_u9_u1_n121 ) , .ZN( u0_u9_u1_n122 ) , .A( u0_u9_u1_n128 ) );
  AOI21_X1 u0_u9_u1_U48 (.A( u0_u9_u1_n128 ) , .B2( u0_u9_u1_n129 ) , .ZN( u0_u9_u1_n130 ) , .B1( u0_u9_u1_n150 ) );
  NAND2_X1 u0_u9_u1_U49 (.ZN( u0_u9_u1_n112 ) , .A1( u0_u9_u1_n169 ) , .A2( u0_u9_u1_n170 ) );
  AOI211_X1 u0_u9_u1_U5 (.ZN( u0_u9_u1_n124 ) , .A( u0_u9_u1_n138 ) , .C2( u0_u9_u1_n139 ) , .B( u0_u9_u1_n145 ) , .C1( u0_u9_u1_n147 ) );
  NAND2_X1 u0_u9_u1_U50 (.ZN( u0_u9_u1_n129 ) , .A2( u0_u9_u1_n95 ) , .A1( u0_u9_u1_n98 ) );
  NAND2_X1 u0_u9_u1_U51 (.A1( u0_u9_u1_n102 ) , .ZN( u0_u9_u1_n154 ) , .A2( u0_u9_u1_n99 ) );
  NAND2_X1 u0_u9_u1_U52 (.A2( u0_u9_u1_n100 ) , .ZN( u0_u9_u1_n135 ) , .A1( u0_u9_u1_n99 ) );
  AOI21_X1 u0_u9_u1_U53 (.A( u0_u9_u1_n152 ) , .B2( u0_u9_u1_n153 ) , .B1( u0_u9_u1_n154 ) , .ZN( u0_u9_u1_n158 ) );
  INV_X1 u0_u9_u1_U54 (.A( u0_u9_u1_n160 ) , .ZN( u0_u9_u1_n175 ) );
  NAND2_X1 u0_u9_u1_U55 (.A1( u0_u9_u1_n100 ) , .ZN( u0_u9_u1_n116 ) , .A2( u0_u9_u1_n95 ) );
  NAND2_X1 u0_u9_u1_U56 (.A1( u0_u9_u1_n102 ) , .ZN( u0_u9_u1_n131 ) , .A2( u0_u9_u1_n95 ) );
  NAND2_X1 u0_u9_u1_U57 (.A2( u0_u9_u1_n104 ) , .ZN( u0_u9_u1_n121 ) , .A1( u0_u9_u1_n98 ) );
  NAND2_X1 u0_u9_u1_U58 (.A1( u0_u9_u1_n103 ) , .ZN( u0_u9_u1_n153 ) , .A2( u0_u9_u1_n98 ) );
  NAND2_X1 u0_u9_u1_U59 (.A2( u0_u9_u1_n104 ) , .A1( u0_u9_u1_n105 ) , .ZN( u0_u9_u1_n133 ) );
  AOI22_X1 u0_u9_u1_U6 (.B2( u0_u9_u1_n136 ) , .A2( u0_u9_u1_n137 ) , .ZN( u0_u9_u1_n143 ) , .A1( u0_u9_u1_n171 ) , .B1( u0_u9_u1_n173 ) );
  NAND2_X1 u0_u9_u1_U60 (.ZN( u0_u9_u1_n150 ) , .A2( u0_u9_u1_n98 ) , .A1( u0_u9_u1_n99 ) );
  NAND2_X1 u0_u9_u1_U61 (.A1( u0_u9_u1_n105 ) , .ZN( u0_u9_u1_n155 ) , .A2( u0_u9_u1_n95 ) );
  OAI21_X1 u0_u9_u1_U62 (.ZN( u0_u9_u1_n109 ) , .B1( u0_u9_u1_n129 ) , .B2( u0_u9_u1_n160 ) , .A( u0_u9_u1_n167 ) );
  NAND2_X1 u0_u9_u1_U63 (.A2( u0_u9_u1_n100 ) , .A1( u0_u9_u1_n103 ) , .ZN( u0_u9_u1_n120 ) );
  NAND2_X1 u0_u9_u1_U64 (.A1( u0_u9_u1_n102 ) , .A2( u0_u9_u1_n104 ) , .ZN( u0_u9_u1_n115 ) );
  NAND2_X1 u0_u9_u1_U65 (.A2( u0_u9_u1_n100 ) , .A1( u0_u9_u1_n104 ) , .ZN( u0_u9_u1_n151 ) );
  NAND2_X1 u0_u9_u1_U66 (.A2( u0_u9_u1_n103 ) , .A1( u0_u9_u1_n105 ) , .ZN( u0_u9_u1_n161 ) );
  INV_X1 u0_u9_u1_U67 (.A( u0_u9_u1_n152 ) , .ZN( u0_u9_u1_n173 ) );
  INV_X1 u0_u9_u1_U68 (.A( u0_u9_u1_n128 ) , .ZN( u0_u9_u1_n172 ) );
  NAND2_X1 u0_u9_u1_U69 (.A2( u0_u9_u1_n102 ) , .A1( u0_u9_u1_n103 ) , .ZN( u0_u9_u1_n123 ) );
  INV_X1 u0_u9_u1_U7 (.A( u0_u9_u1_n147 ) , .ZN( u0_u9_u1_n181 ) );
  NOR2_X1 u0_u9_u1_U70 (.A2( u0_u9_X_7 ) , .A1( u0_u9_X_8 ) , .ZN( u0_u9_u1_n95 ) );
  NOR2_X1 u0_u9_u1_U71 (.A1( u0_u9_X_12 ) , .A2( u0_u9_X_9 ) , .ZN( u0_u9_u1_n100 ) );
  NOR2_X1 u0_u9_u1_U72 (.A2( u0_u9_X_8 ) , .A1( u0_u9_u1_n177 ) , .ZN( u0_u9_u1_n99 ) );
  NOR2_X1 u0_u9_u1_U73 (.A2( u0_u9_X_12 ) , .ZN( u0_u9_u1_n102 ) , .A1( u0_u9_u1_n176 ) );
  NOR2_X1 u0_u9_u1_U74 (.A2( u0_u9_X_9 ) , .ZN( u0_u9_u1_n105 ) , .A1( u0_u9_u1_n168 ) );
  NAND2_X1 u0_u9_u1_U75 (.A1( u0_u9_X_10 ) , .ZN( u0_u9_u1_n160 ) , .A2( u0_u9_u1_n169 ) );
  NAND2_X1 u0_u9_u1_U76 (.A2( u0_u9_X_10 ) , .A1( u0_u9_X_11 ) , .ZN( u0_u9_u1_n152 ) );
  NAND2_X1 u0_u9_u1_U77 (.A1( u0_u9_X_11 ) , .ZN( u0_u9_u1_n128 ) , .A2( u0_u9_u1_n170 ) );
  AND2_X1 u0_u9_u1_U78 (.A2( u0_u9_X_7 ) , .A1( u0_u9_X_8 ) , .ZN( u0_u9_u1_n104 ) );
  AND2_X1 u0_u9_u1_U79 (.A1( u0_u9_X_8 ) , .ZN( u0_u9_u1_n103 ) , .A2( u0_u9_u1_n177 ) );
  AOI22_X1 u0_u9_u1_U8 (.B2( u0_u9_u1_n113 ) , .A2( u0_u9_u1_n114 ) , .ZN( u0_u9_u1_n125 ) , .A1( u0_u9_u1_n171 ) , .B1( u0_u9_u1_n173 ) );
  INV_X1 u0_u9_u1_U80 (.A( u0_u9_X_10 ) , .ZN( u0_u9_u1_n170 ) );
  INV_X1 u0_u9_u1_U81 (.A( u0_u9_X_9 ) , .ZN( u0_u9_u1_n176 ) );
  INV_X1 u0_u9_u1_U82 (.A( u0_u9_X_11 ) , .ZN( u0_u9_u1_n169 ) );
  INV_X1 u0_u9_u1_U83 (.A( u0_u9_X_12 ) , .ZN( u0_u9_u1_n168 ) );
  INV_X1 u0_u9_u1_U84 (.A( u0_u9_X_7 ) , .ZN( u0_u9_u1_n177 ) );
  NAND4_X1 u0_u9_u1_U85 (.ZN( u0_out9_28 ) , .A4( u0_u9_u1_n124 ) , .A3( u0_u9_u1_n125 ) , .A2( u0_u9_u1_n126 ) , .A1( u0_u9_u1_n127 ) );
  OAI21_X1 u0_u9_u1_U86 (.ZN( u0_u9_u1_n127 ) , .B2( u0_u9_u1_n139 ) , .B1( u0_u9_u1_n175 ) , .A( u0_u9_u1_n183 ) );
  OAI21_X1 u0_u9_u1_U87 (.ZN( u0_u9_u1_n126 ) , .B2( u0_u9_u1_n140 ) , .A( u0_u9_u1_n146 ) , .B1( u0_u9_u1_n178 ) );
  NAND4_X1 u0_u9_u1_U88 (.ZN( u0_out9_18 ) , .A4( u0_u9_u1_n165 ) , .A3( u0_u9_u1_n166 ) , .A1( u0_u9_u1_n167 ) , .A2( u0_u9_u1_n186 ) );
  AOI22_X1 u0_u9_u1_U89 (.B2( u0_u9_u1_n146 ) , .B1( u0_u9_u1_n147 ) , .A2( u0_u9_u1_n148 ) , .ZN( u0_u9_u1_n166 ) , .A1( u0_u9_u1_n172 ) );
  NAND2_X1 u0_u9_u1_U9 (.ZN( u0_u9_u1_n114 ) , .A1( u0_u9_u1_n134 ) , .A2( u0_u9_u1_n156 ) );
  INV_X1 u0_u9_u1_U90 (.A( u0_u9_u1_n145 ) , .ZN( u0_u9_u1_n186 ) );
  NAND4_X1 u0_u9_u1_U91 (.ZN( u0_out9_2 ) , .A4( u0_u9_u1_n142 ) , .A3( u0_u9_u1_n143 ) , .A2( u0_u9_u1_n144 ) , .A1( u0_u9_u1_n179 ) );
  OAI21_X1 u0_u9_u1_U92 (.B2( u0_u9_u1_n132 ) , .ZN( u0_u9_u1_n144 ) , .A( u0_u9_u1_n146 ) , .B1( u0_u9_u1_n180 ) );
  INV_X1 u0_u9_u1_U93 (.A( u0_u9_u1_n130 ) , .ZN( u0_u9_u1_n179 ) );
  OR4_X1 u0_u9_u1_U94 (.ZN( u0_out9_13 ) , .A4( u0_u9_u1_n108 ) , .A3( u0_u9_u1_n109 ) , .A2( u0_u9_u1_n110 ) , .A1( u0_u9_u1_n111 ) );
  AOI21_X1 u0_u9_u1_U95 (.ZN( u0_u9_u1_n110 ) , .A( u0_u9_u1_n116 ) , .B1( u0_u9_u1_n152 ) , .B2( u0_u9_u1_n160 ) );
  AOI21_X1 u0_u9_u1_U96 (.ZN( u0_u9_u1_n111 ) , .A( u0_u9_u1_n128 ) , .B2( u0_u9_u1_n131 ) , .B1( u0_u9_u1_n135 ) );
  NAND3_X1 u0_u9_u1_U97 (.A3( u0_u9_u1_n149 ) , .A2( u0_u9_u1_n150 ) , .A1( u0_u9_u1_n151 ) , .ZN( u0_u9_u1_n164 ) );
  NAND3_X1 u0_u9_u1_U98 (.A3( u0_u9_u1_n134 ) , .A2( u0_u9_u1_n135 ) , .ZN( u0_u9_u1_n136 ) , .A1( u0_u9_u1_n151 ) );
  NAND3_X1 u0_u9_u1_U99 (.A1( u0_u9_u1_n133 ) , .ZN( u0_u9_u1_n137 ) , .A2( u0_u9_u1_n154 ) , .A3( u0_u9_u1_n181 ) );
  OAI22_X1 u0_u9_u2_U10 (.B1( u0_u9_u2_n151 ) , .A2( u0_u9_u2_n152 ) , .A1( u0_u9_u2_n153 ) , .ZN( u0_u9_u2_n160 ) , .B2( u0_u9_u2_n168 ) );
  NAND3_X1 u0_u9_u2_U100 (.A2( u0_u9_u2_n100 ) , .A1( u0_u9_u2_n104 ) , .A3( u0_u9_u2_n138 ) , .ZN( u0_u9_u2_n98 ) );
  NOR3_X1 u0_u9_u2_U11 (.A1( u0_u9_u2_n150 ) , .ZN( u0_u9_u2_n151 ) , .A3( u0_u9_u2_n175 ) , .A2( u0_u9_u2_n188 ) );
  AOI21_X1 u0_u9_u2_U12 (.B2( u0_u9_u2_n123 ) , .ZN( u0_u9_u2_n125 ) , .A( u0_u9_u2_n171 ) , .B1( u0_u9_u2_n184 ) );
  INV_X1 u0_u9_u2_U13 (.A( u0_u9_u2_n150 ) , .ZN( u0_u9_u2_n184 ) );
  AOI21_X1 u0_u9_u2_U14 (.ZN( u0_u9_u2_n144 ) , .B2( u0_u9_u2_n155 ) , .A( u0_u9_u2_n172 ) , .B1( u0_u9_u2_n185 ) );
  AOI21_X1 u0_u9_u2_U15 (.B2( u0_u9_u2_n143 ) , .ZN( u0_u9_u2_n145 ) , .B1( u0_u9_u2_n152 ) , .A( u0_u9_u2_n171 ) );
  INV_X1 u0_u9_u2_U16 (.A( u0_u9_u2_n156 ) , .ZN( u0_u9_u2_n171 ) );
  INV_X1 u0_u9_u2_U17 (.A( u0_u9_u2_n120 ) , .ZN( u0_u9_u2_n188 ) );
  NAND2_X1 u0_u9_u2_U18 (.A2( u0_u9_u2_n122 ) , .ZN( u0_u9_u2_n150 ) , .A1( u0_u9_u2_n152 ) );
  INV_X1 u0_u9_u2_U19 (.A( u0_u9_u2_n153 ) , .ZN( u0_u9_u2_n170 ) );
  INV_X1 u0_u9_u2_U20 (.A( u0_u9_u2_n137 ) , .ZN( u0_u9_u2_n173 ) );
  NAND2_X1 u0_u9_u2_U21 (.A1( u0_u9_u2_n132 ) , .A2( u0_u9_u2_n139 ) , .ZN( u0_u9_u2_n157 ) );
  INV_X1 u0_u9_u2_U22 (.A( u0_u9_u2_n113 ) , .ZN( u0_u9_u2_n178 ) );
  INV_X1 u0_u9_u2_U23 (.A( u0_u9_u2_n139 ) , .ZN( u0_u9_u2_n175 ) );
  INV_X1 u0_u9_u2_U24 (.A( u0_u9_u2_n155 ) , .ZN( u0_u9_u2_n181 ) );
  INV_X1 u0_u9_u2_U25 (.A( u0_u9_u2_n119 ) , .ZN( u0_u9_u2_n177 ) );
  INV_X1 u0_u9_u2_U26 (.A( u0_u9_u2_n116 ) , .ZN( u0_u9_u2_n180 ) );
  INV_X1 u0_u9_u2_U27 (.A( u0_u9_u2_n131 ) , .ZN( u0_u9_u2_n179 ) );
  INV_X1 u0_u9_u2_U28 (.A( u0_u9_u2_n154 ) , .ZN( u0_u9_u2_n176 ) );
  NAND2_X1 u0_u9_u2_U29 (.A2( u0_u9_u2_n116 ) , .A1( u0_u9_u2_n117 ) , .ZN( u0_u9_u2_n118 ) );
  NOR2_X1 u0_u9_u2_U3 (.ZN( u0_u9_u2_n121 ) , .A2( u0_u9_u2_n177 ) , .A1( u0_u9_u2_n180 ) );
  INV_X1 u0_u9_u2_U30 (.A( u0_u9_u2_n132 ) , .ZN( u0_u9_u2_n182 ) );
  INV_X1 u0_u9_u2_U31 (.A( u0_u9_u2_n158 ) , .ZN( u0_u9_u2_n183 ) );
  OAI21_X1 u0_u9_u2_U32 (.A( u0_u9_u2_n156 ) , .B1( u0_u9_u2_n157 ) , .ZN( u0_u9_u2_n158 ) , .B2( u0_u9_u2_n179 ) );
  NOR2_X1 u0_u9_u2_U33 (.ZN( u0_u9_u2_n156 ) , .A1( u0_u9_u2_n166 ) , .A2( u0_u9_u2_n169 ) );
  NOR2_X1 u0_u9_u2_U34 (.A2( u0_u9_u2_n114 ) , .ZN( u0_u9_u2_n137 ) , .A1( u0_u9_u2_n140 ) );
  NOR2_X1 u0_u9_u2_U35 (.A2( u0_u9_u2_n138 ) , .ZN( u0_u9_u2_n153 ) , .A1( u0_u9_u2_n156 ) );
  AOI211_X1 u0_u9_u2_U36 (.ZN( u0_u9_u2_n130 ) , .C1( u0_u9_u2_n138 ) , .C2( u0_u9_u2_n179 ) , .B( u0_u9_u2_n96 ) , .A( u0_u9_u2_n97 ) );
  OAI22_X1 u0_u9_u2_U37 (.B1( u0_u9_u2_n133 ) , .A2( u0_u9_u2_n137 ) , .A1( u0_u9_u2_n152 ) , .B2( u0_u9_u2_n168 ) , .ZN( u0_u9_u2_n97 ) );
  OAI221_X1 u0_u9_u2_U38 (.B1( u0_u9_u2_n113 ) , .C1( u0_u9_u2_n132 ) , .A( u0_u9_u2_n149 ) , .B2( u0_u9_u2_n171 ) , .C2( u0_u9_u2_n172 ) , .ZN( u0_u9_u2_n96 ) );
  OAI221_X1 u0_u9_u2_U39 (.A( u0_u9_u2_n115 ) , .C2( u0_u9_u2_n123 ) , .B2( u0_u9_u2_n143 ) , .B1( u0_u9_u2_n153 ) , .ZN( u0_u9_u2_n163 ) , .C1( u0_u9_u2_n168 ) );
  INV_X1 u0_u9_u2_U4 (.A( u0_u9_u2_n134 ) , .ZN( u0_u9_u2_n185 ) );
  OAI21_X1 u0_u9_u2_U40 (.A( u0_u9_u2_n114 ) , .ZN( u0_u9_u2_n115 ) , .B1( u0_u9_u2_n176 ) , .B2( u0_u9_u2_n178 ) );
  OAI221_X1 u0_u9_u2_U41 (.A( u0_u9_u2_n135 ) , .B2( u0_u9_u2_n136 ) , .B1( u0_u9_u2_n137 ) , .ZN( u0_u9_u2_n162 ) , .C2( u0_u9_u2_n167 ) , .C1( u0_u9_u2_n185 ) );
  AND3_X1 u0_u9_u2_U42 (.A3( u0_u9_u2_n131 ) , .A2( u0_u9_u2_n132 ) , .A1( u0_u9_u2_n133 ) , .ZN( u0_u9_u2_n136 ) );
  AOI22_X1 u0_u9_u2_U43 (.ZN( u0_u9_u2_n135 ) , .B1( u0_u9_u2_n140 ) , .A1( u0_u9_u2_n156 ) , .B2( u0_u9_u2_n180 ) , .A2( u0_u9_u2_n188 ) );
  AOI21_X1 u0_u9_u2_U44 (.ZN( u0_u9_u2_n149 ) , .B1( u0_u9_u2_n173 ) , .B2( u0_u9_u2_n188 ) , .A( u0_u9_u2_n95 ) );
  AND3_X1 u0_u9_u2_U45 (.A2( u0_u9_u2_n100 ) , .A1( u0_u9_u2_n104 ) , .A3( u0_u9_u2_n156 ) , .ZN( u0_u9_u2_n95 ) );
  OAI21_X1 u0_u9_u2_U46 (.A( u0_u9_u2_n141 ) , .B2( u0_u9_u2_n142 ) , .ZN( u0_u9_u2_n146 ) , .B1( u0_u9_u2_n153 ) );
  OAI21_X1 u0_u9_u2_U47 (.A( u0_u9_u2_n140 ) , .ZN( u0_u9_u2_n141 ) , .B1( u0_u9_u2_n176 ) , .B2( u0_u9_u2_n177 ) );
  NOR3_X1 u0_u9_u2_U48 (.ZN( u0_u9_u2_n142 ) , .A3( u0_u9_u2_n175 ) , .A2( u0_u9_u2_n178 ) , .A1( u0_u9_u2_n181 ) );
  OAI21_X1 u0_u9_u2_U49 (.A( u0_u9_u2_n101 ) , .B2( u0_u9_u2_n121 ) , .B1( u0_u9_u2_n153 ) , .ZN( u0_u9_u2_n164 ) );
  NOR4_X1 u0_u9_u2_U5 (.A4( u0_u9_u2_n124 ) , .A3( u0_u9_u2_n125 ) , .A2( u0_u9_u2_n126 ) , .A1( u0_u9_u2_n127 ) , .ZN( u0_u9_u2_n128 ) );
  NAND2_X1 u0_u9_u2_U50 (.A2( u0_u9_u2_n100 ) , .A1( u0_u9_u2_n107 ) , .ZN( u0_u9_u2_n155 ) );
  NAND2_X1 u0_u9_u2_U51 (.A2( u0_u9_u2_n105 ) , .A1( u0_u9_u2_n108 ) , .ZN( u0_u9_u2_n143 ) );
  NAND2_X1 u0_u9_u2_U52 (.A1( u0_u9_u2_n104 ) , .A2( u0_u9_u2_n106 ) , .ZN( u0_u9_u2_n152 ) );
  NAND2_X1 u0_u9_u2_U53 (.A1( u0_u9_u2_n100 ) , .A2( u0_u9_u2_n105 ) , .ZN( u0_u9_u2_n132 ) );
  INV_X1 u0_u9_u2_U54 (.A( u0_u9_u2_n140 ) , .ZN( u0_u9_u2_n168 ) );
  INV_X1 u0_u9_u2_U55 (.A( u0_u9_u2_n138 ) , .ZN( u0_u9_u2_n167 ) );
  NAND2_X1 u0_u9_u2_U56 (.A1( u0_u9_u2_n102 ) , .A2( u0_u9_u2_n106 ) , .ZN( u0_u9_u2_n113 ) );
  NAND2_X1 u0_u9_u2_U57 (.A1( u0_u9_u2_n106 ) , .A2( u0_u9_u2_n107 ) , .ZN( u0_u9_u2_n131 ) );
  NAND2_X1 u0_u9_u2_U58 (.A1( u0_u9_u2_n103 ) , .A2( u0_u9_u2_n107 ) , .ZN( u0_u9_u2_n139 ) );
  NAND2_X1 u0_u9_u2_U59 (.A1( u0_u9_u2_n103 ) , .A2( u0_u9_u2_n105 ) , .ZN( u0_u9_u2_n133 ) );
  AOI21_X1 u0_u9_u2_U6 (.B2( u0_u9_u2_n119 ) , .ZN( u0_u9_u2_n127 ) , .A( u0_u9_u2_n137 ) , .B1( u0_u9_u2_n155 ) );
  NAND2_X1 u0_u9_u2_U60 (.A1( u0_u9_u2_n102 ) , .A2( u0_u9_u2_n103 ) , .ZN( u0_u9_u2_n154 ) );
  NAND2_X1 u0_u9_u2_U61 (.A2( u0_u9_u2_n103 ) , .A1( u0_u9_u2_n104 ) , .ZN( u0_u9_u2_n119 ) );
  NAND2_X1 u0_u9_u2_U62 (.A2( u0_u9_u2_n107 ) , .A1( u0_u9_u2_n108 ) , .ZN( u0_u9_u2_n123 ) );
  NAND2_X1 u0_u9_u2_U63 (.A1( u0_u9_u2_n104 ) , .A2( u0_u9_u2_n108 ) , .ZN( u0_u9_u2_n122 ) );
  INV_X1 u0_u9_u2_U64 (.A( u0_u9_u2_n114 ) , .ZN( u0_u9_u2_n172 ) );
  NAND2_X1 u0_u9_u2_U65 (.A2( u0_u9_u2_n100 ) , .A1( u0_u9_u2_n102 ) , .ZN( u0_u9_u2_n116 ) );
  NAND2_X1 u0_u9_u2_U66 (.A1( u0_u9_u2_n102 ) , .A2( u0_u9_u2_n108 ) , .ZN( u0_u9_u2_n120 ) );
  NAND2_X1 u0_u9_u2_U67 (.A2( u0_u9_u2_n105 ) , .A1( u0_u9_u2_n106 ) , .ZN( u0_u9_u2_n117 ) );
  INV_X1 u0_u9_u2_U68 (.ZN( u0_u9_u2_n187 ) , .A( u0_u9_u2_n99 ) );
  OAI21_X1 u0_u9_u2_U69 (.B1( u0_u9_u2_n137 ) , .B2( u0_u9_u2_n143 ) , .A( u0_u9_u2_n98 ) , .ZN( u0_u9_u2_n99 ) );
  AOI21_X1 u0_u9_u2_U7 (.ZN( u0_u9_u2_n124 ) , .B1( u0_u9_u2_n131 ) , .B2( u0_u9_u2_n143 ) , .A( u0_u9_u2_n172 ) );
  NOR2_X1 u0_u9_u2_U70 (.A2( u0_u9_X_16 ) , .ZN( u0_u9_u2_n140 ) , .A1( u0_u9_u2_n166 ) );
  NOR2_X1 u0_u9_u2_U71 (.A2( u0_u9_X_13 ) , .A1( u0_u9_X_14 ) , .ZN( u0_u9_u2_n100 ) );
  NOR2_X1 u0_u9_u2_U72 (.A2( u0_u9_X_16 ) , .A1( u0_u9_X_17 ) , .ZN( u0_u9_u2_n138 ) );
  NOR2_X1 u0_u9_u2_U73 (.A2( u0_u9_X_15 ) , .A1( u0_u9_X_18 ) , .ZN( u0_u9_u2_n104 ) );
  NOR2_X1 u0_u9_u2_U74 (.A2( u0_u9_X_14 ) , .ZN( u0_u9_u2_n103 ) , .A1( u0_u9_u2_n174 ) );
  NOR2_X1 u0_u9_u2_U75 (.A2( u0_u9_X_15 ) , .ZN( u0_u9_u2_n102 ) , .A1( u0_u9_u2_n165 ) );
  NOR2_X1 u0_u9_u2_U76 (.A2( u0_u9_X_17 ) , .ZN( u0_u9_u2_n114 ) , .A1( u0_u9_u2_n169 ) );
  AND2_X1 u0_u9_u2_U77 (.A1( u0_u9_X_15 ) , .ZN( u0_u9_u2_n105 ) , .A2( u0_u9_u2_n165 ) );
  AND2_X1 u0_u9_u2_U78 (.A2( u0_u9_X_15 ) , .A1( u0_u9_X_18 ) , .ZN( u0_u9_u2_n107 ) );
  AND2_X1 u0_u9_u2_U79 (.A1( u0_u9_X_14 ) , .ZN( u0_u9_u2_n106 ) , .A2( u0_u9_u2_n174 ) );
  AOI21_X1 u0_u9_u2_U8 (.B2( u0_u9_u2_n120 ) , .B1( u0_u9_u2_n121 ) , .ZN( u0_u9_u2_n126 ) , .A( u0_u9_u2_n167 ) );
  AND2_X1 u0_u9_u2_U80 (.A1( u0_u9_X_13 ) , .A2( u0_u9_X_14 ) , .ZN( u0_u9_u2_n108 ) );
  INV_X1 u0_u9_u2_U81 (.A( u0_u9_X_16 ) , .ZN( u0_u9_u2_n169 ) );
  INV_X1 u0_u9_u2_U82 (.A( u0_u9_X_17 ) , .ZN( u0_u9_u2_n166 ) );
  INV_X1 u0_u9_u2_U83 (.A( u0_u9_X_13 ) , .ZN( u0_u9_u2_n174 ) );
  INV_X1 u0_u9_u2_U84 (.A( u0_u9_X_18 ) , .ZN( u0_u9_u2_n165 ) );
  NAND4_X1 u0_u9_u2_U85 (.ZN( u0_out9_30 ) , .A4( u0_u9_u2_n147 ) , .A3( u0_u9_u2_n148 ) , .A2( u0_u9_u2_n149 ) , .A1( u0_u9_u2_n187 ) );
  AOI21_X1 u0_u9_u2_U86 (.B2( u0_u9_u2_n138 ) , .ZN( u0_u9_u2_n148 ) , .A( u0_u9_u2_n162 ) , .B1( u0_u9_u2_n182 ) );
  NOR3_X1 u0_u9_u2_U87 (.A3( u0_u9_u2_n144 ) , .A2( u0_u9_u2_n145 ) , .A1( u0_u9_u2_n146 ) , .ZN( u0_u9_u2_n147 ) );
  NAND4_X1 u0_u9_u2_U88 (.ZN( u0_out9_24 ) , .A4( u0_u9_u2_n111 ) , .A3( u0_u9_u2_n112 ) , .A1( u0_u9_u2_n130 ) , .A2( u0_u9_u2_n187 ) );
  AOI221_X1 u0_u9_u2_U89 (.A( u0_u9_u2_n109 ) , .B1( u0_u9_u2_n110 ) , .ZN( u0_u9_u2_n111 ) , .C1( u0_u9_u2_n134 ) , .C2( u0_u9_u2_n170 ) , .B2( u0_u9_u2_n173 ) );
  OAI22_X1 u0_u9_u2_U9 (.ZN( u0_u9_u2_n109 ) , .A2( u0_u9_u2_n113 ) , .B2( u0_u9_u2_n133 ) , .B1( u0_u9_u2_n167 ) , .A1( u0_u9_u2_n168 ) );
  AOI21_X1 u0_u9_u2_U90 (.ZN( u0_u9_u2_n112 ) , .B2( u0_u9_u2_n156 ) , .A( u0_u9_u2_n164 ) , .B1( u0_u9_u2_n181 ) );
  NAND4_X1 u0_u9_u2_U91 (.ZN( u0_out9_16 ) , .A4( u0_u9_u2_n128 ) , .A3( u0_u9_u2_n129 ) , .A1( u0_u9_u2_n130 ) , .A2( u0_u9_u2_n186 ) );
  AOI22_X1 u0_u9_u2_U92 (.A2( u0_u9_u2_n118 ) , .ZN( u0_u9_u2_n129 ) , .A1( u0_u9_u2_n140 ) , .B1( u0_u9_u2_n157 ) , .B2( u0_u9_u2_n170 ) );
  INV_X1 u0_u9_u2_U93 (.A( u0_u9_u2_n163 ) , .ZN( u0_u9_u2_n186 ) );
  OR4_X1 u0_u9_u2_U94 (.ZN( u0_out9_6 ) , .A4( u0_u9_u2_n161 ) , .A3( u0_u9_u2_n162 ) , .A2( u0_u9_u2_n163 ) , .A1( u0_u9_u2_n164 ) );
  OR3_X1 u0_u9_u2_U95 (.A2( u0_u9_u2_n159 ) , .A1( u0_u9_u2_n160 ) , .ZN( u0_u9_u2_n161 ) , .A3( u0_u9_u2_n183 ) );
  AOI21_X1 u0_u9_u2_U96 (.B2( u0_u9_u2_n154 ) , .B1( u0_u9_u2_n155 ) , .ZN( u0_u9_u2_n159 ) , .A( u0_u9_u2_n167 ) );
  NAND3_X1 u0_u9_u2_U97 (.A2( u0_u9_u2_n117 ) , .A1( u0_u9_u2_n122 ) , .A3( u0_u9_u2_n123 ) , .ZN( u0_u9_u2_n134 ) );
  NAND3_X1 u0_u9_u2_U98 (.ZN( u0_u9_u2_n110 ) , .A2( u0_u9_u2_n131 ) , .A3( u0_u9_u2_n139 ) , .A1( u0_u9_u2_n154 ) );
  NAND3_X1 u0_u9_u2_U99 (.A2( u0_u9_u2_n100 ) , .ZN( u0_u9_u2_n101 ) , .A1( u0_u9_u2_n104 ) , .A3( u0_u9_u2_n114 ) );
  AOI22_X1 u0_u9_u6_U10 (.A2( u0_u9_u6_n151 ) , .B2( u0_u9_u6_n161 ) , .A1( u0_u9_u6_n167 ) , .B1( u0_u9_u6_n170 ) , .ZN( u0_u9_u6_n89 ) );
  AOI21_X1 u0_u9_u6_U11 (.B1( u0_u9_u6_n107 ) , .B2( u0_u9_u6_n132 ) , .A( u0_u9_u6_n158 ) , .ZN( u0_u9_u6_n88 ) );
  AOI21_X1 u0_u9_u6_U12 (.B2( u0_u9_u6_n147 ) , .B1( u0_u9_u6_n148 ) , .ZN( u0_u9_u6_n149 ) , .A( u0_u9_u6_n158 ) );
  AOI21_X1 u0_u9_u6_U13 (.ZN( u0_u9_u6_n106 ) , .A( u0_u9_u6_n142 ) , .B2( u0_u9_u6_n159 ) , .B1( u0_u9_u6_n164 ) );
  INV_X1 u0_u9_u6_U14 (.A( u0_u9_u6_n155 ) , .ZN( u0_u9_u6_n161 ) );
  INV_X1 u0_u9_u6_U15 (.A( u0_u9_u6_n128 ) , .ZN( u0_u9_u6_n164 ) );
  NAND2_X1 u0_u9_u6_U16 (.ZN( u0_u9_u6_n110 ) , .A1( u0_u9_u6_n122 ) , .A2( u0_u9_u6_n129 ) );
  NAND2_X1 u0_u9_u6_U17 (.ZN( u0_u9_u6_n124 ) , .A2( u0_u9_u6_n146 ) , .A1( u0_u9_u6_n148 ) );
  INV_X1 u0_u9_u6_U18 (.A( u0_u9_u6_n132 ) , .ZN( u0_u9_u6_n171 ) );
  AND2_X1 u0_u9_u6_U19 (.A1( u0_u9_u6_n100 ) , .ZN( u0_u9_u6_n130 ) , .A2( u0_u9_u6_n147 ) );
  INV_X1 u0_u9_u6_U20 (.A( u0_u9_u6_n127 ) , .ZN( u0_u9_u6_n173 ) );
  INV_X1 u0_u9_u6_U21 (.A( u0_u9_u6_n121 ) , .ZN( u0_u9_u6_n167 ) );
  INV_X1 u0_u9_u6_U22 (.A( u0_u9_u6_n100 ) , .ZN( u0_u9_u6_n169 ) );
  INV_X1 u0_u9_u6_U23 (.A( u0_u9_u6_n123 ) , .ZN( u0_u9_u6_n170 ) );
  INV_X1 u0_u9_u6_U24 (.A( u0_u9_u6_n113 ) , .ZN( u0_u9_u6_n168 ) );
  AND2_X1 u0_u9_u6_U25 (.A1( u0_u9_u6_n107 ) , .A2( u0_u9_u6_n119 ) , .ZN( u0_u9_u6_n133 ) );
  AND2_X1 u0_u9_u6_U26 (.A2( u0_u9_u6_n121 ) , .A1( u0_u9_u6_n122 ) , .ZN( u0_u9_u6_n131 ) );
  AND3_X1 u0_u9_u6_U27 (.ZN( u0_u9_u6_n120 ) , .A2( u0_u9_u6_n127 ) , .A1( u0_u9_u6_n132 ) , .A3( u0_u9_u6_n145 ) );
  INV_X1 u0_u9_u6_U28 (.A( u0_u9_u6_n146 ) , .ZN( u0_u9_u6_n163 ) );
  AOI222_X1 u0_u9_u6_U29 (.ZN( u0_u9_u6_n114 ) , .A1( u0_u9_u6_n118 ) , .A2( u0_u9_u6_n126 ) , .B2( u0_u9_u6_n151 ) , .C2( u0_u9_u6_n159 ) , .C1( u0_u9_u6_n168 ) , .B1( u0_u9_u6_n169 ) );
  INV_X1 u0_u9_u6_U3 (.A( u0_u9_u6_n110 ) , .ZN( u0_u9_u6_n166 ) );
  NOR2_X1 u0_u9_u6_U30 (.A1( u0_u9_u6_n162 ) , .A2( u0_u9_u6_n165 ) , .ZN( u0_u9_u6_n98 ) );
  NAND2_X1 u0_u9_u6_U31 (.A1( u0_u9_u6_n144 ) , .ZN( u0_u9_u6_n151 ) , .A2( u0_u9_u6_n158 ) );
  NAND2_X1 u0_u9_u6_U32 (.ZN( u0_u9_u6_n132 ) , .A1( u0_u9_u6_n91 ) , .A2( u0_u9_u6_n97 ) );
  AOI22_X1 u0_u9_u6_U33 (.B2( u0_u9_u6_n110 ) , .B1( u0_u9_u6_n111 ) , .A1( u0_u9_u6_n112 ) , .ZN( u0_u9_u6_n115 ) , .A2( u0_u9_u6_n161 ) );
  NAND4_X1 u0_u9_u6_U34 (.A3( u0_u9_u6_n109 ) , .ZN( u0_u9_u6_n112 ) , .A4( u0_u9_u6_n132 ) , .A2( u0_u9_u6_n147 ) , .A1( u0_u9_u6_n166 ) );
  NOR2_X1 u0_u9_u6_U35 (.ZN( u0_u9_u6_n109 ) , .A1( u0_u9_u6_n170 ) , .A2( u0_u9_u6_n173 ) );
  NOR2_X1 u0_u9_u6_U36 (.A2( u0_u9_u6_n126 ) , .ZN( u0_u9_u6_n155 ) , .A1( u0_u9_u6_n160 ) );
  NAND2_X1 u0_u9_u6_U37 (.ZN( u0_u9_u6_n146 ) , .A2( u0_u9_u6_n94 ) , .A1( u0_u9_u6_n99 ) );
  AOI21_X1 u0_u9_u6_U38 (.A( u0_u9_u6_n144 ) , .B2( u0_u9_u6_n145 ) , .B1( u0_u9_u6_n146 ) , .ZN( u0_u9_u6_n150 ) );
  AOI211_X1 u0_u9_u6_U39 (.B( u0_u9_u6_n134 ) , .A( u0_u9_u6_n135 ) , .C1( u0_u9_u6_n136 ) , .ZN( u0_u9_u6_n137 ) , .C2( u0_u9_u6_n151 ) );
  INV_X1 u0_u9_u6_U4 (.A( u0_u9_u6_n142 ) , .ZN( u0_u9_u6_n174 ) );
  NAND4_X1 u0_u9_u6_U40 (.A4( u0_u9_u6_n127 ) , .A3( u0_u9_u6_n128 ) , .A2( u0_u9_u6_n129 ) , .A1( u0_u9_u6_n130 ) , .ZN( u0_u9_u6_n136 ) );
  AOI21_X1 u0_u9_u6_U41 (.B2( u0_u9_u6_n132 ) , .B1( u0_u9_u6_n133 ) , .ZN( u0_u9_u6_n134 ) , .A( u0_u9_u6_n158 ) );
  AOI21_X1 u0_u9_u6_U42 (.B1( u0_u9_u6_n131 ) , .ZN( u0_u9_u6_n135 ) , .A( u0_u9_u6_n144 ) , .B2( u0_u9_u6_n146 ) );
  INV_X1 u0_u9_u6_U43 (.A( u0_u9_u6_n111 ) , .ZN( u0_u9_u6_n158 ) );
  NAND2_X1 u0_u9_u6_U44 (.ZN( u0_u9_u6_n127 ) , .A1( u0_u9_u6_n91 ) , .A2( u0_u9_u6_n92 ) );
  NAND2_X1 u0_u9_u6_U45 (.ZN( u0_u9_u6_n129 ) , .A2( u0_u9_u6_n95 ) , .A1( u0_u9_u6_n96 ) );
  INV_X1 u0_u9_u6_U46 (.A( u0_u9_u6_n144 ) , .ZN( u0_u9_u6_n159 ) );
  NAND2_X1 u0_u9_u6_U47 (.ZN( u0_u9_u6_n145 ) , .A2( u0_u9_u6_n97 ) , .A1( u0_u9_u6_n98 ) );
  NAND2_X1 u0_u9_u6_U48 (.ZN( u0_u9_u6_n148 ) , .A2( u0_u9_u6_n92 ) , .A1( u0_u9_u6_n94 ) );
  NAND2_X1 u0_u9_u6_U49 (.ZN( u0_u9_u6_n108 ) , .A2( u0_u9_u6_n139 ) , .A1( u0_u9_u6_n144 ) );
  NAND2_X1 u0_u9_u6_U5 (.A2( u0_u9_u6_n143 ) , .ZN( u0_u9_u6_n152 ) , .A1( u0_u9_u6_n166 ) );
  NAND2_X1 u0_u9_u6_U50 (.ZN( u0_u9_u6_n121 ) , .A2( u0_u9_u6_n95 ) , .A1( u0_u9_u6_n97 ) );
  NAND2_X1 u0_u9_u6_U51 (.ZN( u0_u9_u6_n107 ) , .A2( u0_u9_u6_n92 ) , .A1( u0_u9_u6_n95 ) );
  AND2_X1 u0_u9_u6_U52 (.ZN( u0_u9_u6_n118 ) , .A2( u0_u9_u6_n91 ) , .A1( u0_u9_u6_n99 ) );
  NAND2_X1 u0_u9_u6_U53 (.ZN( u0_u9_u6_n147 ) , .A2( u0_u9_u6_n98 ) , .A1( u0_u9_u6_n99 ) );
  NAND2_X1 u0_u9_u6_U54 (.ZN( u0_u9_u6_n128 ) , .A1( u0_u9_u6_n94 ) , .A2( u0_u9_u6_n96 ) );
  NAND2_X1 u0_u9_u6_U55 (.ZN( u0_u9_u6_n119 ) , .A2( u0_u9_u6_n95 ) , .A1( u0_u9_u6_n99 ) );
  NAND2_X1 u0_u9_u6_U56 (.ZN( u0_u9_u6_n123 ) , .A2( u0_u9_u6_n91 ) , .A1( u0_u9_u6_n96 ) );
  NAND2_X1 u0_u9_u6_U57 (.ZN( u0_u9_u6_n100 ) , .A2( u0_u9_u6_n92 ) , .A1( u0_u9_u6_n98 ) );
  NAND2_X1 u0_u9_u6_U58 (.ZN( u0_u9_u6_n122 ) , .A1( u0_u9_u6_n94 ) , .A2( u0_u9_u6_n97 ) );
  INV_X1 u0_u9_u6_U59 (.A( u0_u9_u6_n139 ) , .ZN( u0_u9_u6_n160 ) );
  AOI22_X1 u0_u9_u6_U6 (.B2( u0_u9_u6_n101 ) , .A1( u0_u9_u6_n102 ) , .ZN( u0_u9_u6_n103 ) , .B1( u0_u9_u6_n160 ) , .A2( u0_u9_u6_n161 ) );
  NAND2_X1 u0_u9_u6_U60 (.ZN( u0_u9_u6_n113 ) , .A1( u0_u9_u6_n96 ) , .A2( u0_u9_u6_n98 ) );
  NOR2_X1 u0_u9_u6_U61 (.A2( u0_u9_X_40 ) , .A1( u0_u9_X_41 ) , .ZN( u0_u9_u6_n126 ) );
  NOR2_X1 u0_u9_u6_U62 (.A2( u0_u9_X_39 ) , .A1( u0_u9_X_42 ) , .ZN( u0_u9_u6_n92 ) );
  NOR2_X1 u0_u9_u6_U63 (.A2( u0_u9_X_39 ) , .A1( u0_u9_u6_n156 ) , .ZN( u0_u9_u6_n97 ) );
  NOR2_X1 u0_u9_u6_U64 (.A2( u0_u9_X_38 ) , .A1( u0_u9_u6_n165 ) , .ZN( u0_u9_u6_n95 ) );
  NOR2_X1 u0_u9_u6_U65 (.A2( u0_u9_X_41 ) , .ZN( u0_u9_u6_n111 ) , .A1( u0_u9_u6_n157 ) );
  NOR2_X1 u0_u9_u6_U66 (.A2( u0_u9_X_37 ) , .A1( u0_u9_u6_n162 ) , .ZN( u0_u9_u6_n94 ) );
  NOR2_X1 u0_u9_u6_U67 (.A2( u0_u9_X_37 ) , .A1( u0_u9_X_38 ) , .ZN( u0_u9_u6_n91 ) );
  NAND2_X1 u0_u9_u6_U68 (.A1( u0_u9_X_41 ) , .ZN( u0_u9_u6_n144 ) , .A2( u0_u9_u6_n157 ) );
  NAND2_X1 u0_u9_u6_U69 (.A2( u0_u9_X_40 ) , .A1( u0_u9_X_41 ) , .ZN( u0_u9_u6_n139 ) );
  NOR2_X1 u0_u9_u6_U7 (.A1( u0_u9_u6_n118 ) , .ZN( u0_u9_u6_n143 ) , .A2( u0_u9_u6_n168 ) );
  AND2_X1 u0_u9_u6_U70 (.A1( u0_u9_X_39 ) , .A2( u0_u9_u6_n156 ) , .ZN( u0_u9_u6_n96 ) );
  AND2_X1 u0_u9_u6_U71 (.A1( u0_u9_X_39 ) , .A2( u0_u9_X_42 ) , .ZN( u0_u9_u6_n99 ) );
  INV_X1 u0_u9_u6_U72 (.A( u0_u9_X_40 ) , .ZN( u0_u9_u6_n157 ) );
  INV_X1 u0_u9_u6_U73 (.A( u0_u9_X_37 ) , .ZN( u0_u9_u6_n165 ) );
  INV_X1 u0_u9_u6_U74 (.A( u0_u9_X_38 ) , .ZN( u0_u9_u6_n162 ) );
  INV_X1 u0_u9_u6_U75 (.A( u0_u9_X_42 ) , .ZN( u0_u9_u6_n156 ) );
  NAND4_X1 u0_u9_u6_U76 (.ZN( u0_out9_32 ) , .A4( u0_u9_u6_n103 ) , .A3( u0_u9_u6_n104 ) , .A2( u0_u9_u6_n105 ) , .A1( u0_u9_u6_n106 ) );
  AOI22_X1 u0_u9_u6_U77 (.ZN( u0_u9_u6_n105 ) , .A2( u0_u9_u6_n108 ) , .A1( u0_u9_u6_n118 ) , .B2( u0_u9_u6_n126 ) , .B1( u0_u9_u6_n171 ) );
  AOI22_X1 u0_u9_u6_U78 (.ZN( u0_u9_u6_n104 ) , .A1( u0_u9_u6_n111 ) , .B1( u0_u9_u6_n124 ) , .B2( u0_u9_u6_n151 ) , .A2( u0_u9_u6_n93 ) );
  NAND4_X1 u0_u9_u6_U79 (.ZN( u0_out9_12 ) , .A4( u0_u9_u6_n114 ) , .A3( u0_u9_u6_n115 ) , .A2( u0_u9_u6_n116 ) , .A1( u0_u9_u6_n117 ) );
  OAI21_X1 u0_u9_u6_U8 (.A( u0_u9_u6_n159 ) , .B1( u0_u9_u6_n169 ) , .B2( u0_u9_u6_n173 ) , .ZN( u0_u9_u6_n90 ) );
  OAI22_X1 u0_u9_u6_U80 (.B2( u0_u9_u6_n111 ) , .ZN( u0_u9_u6_n116 ) , .B1( u0_u9_u6_n126 ) , .A2( u0_u9_u6_n164 ) , .A1( u0_u9_u6_n167 ) );
  OAI21_X1 u0_u9_u6_U81 (.A( u0_u9_u6_n108 ) , .ZN( u0_u9_u6_n117 ) , .B2( u0_u9_u6_n141 ) , .B1( u0_u9_u6_n163 ) );
  OAI211_X1 u0_u9_u6_U82 (.ZN( u0_out9_7 ) , .B( u0_u9_u6_n153 ) , .C2( u0_u9_u6_n154 ) , .C1( u0_u9_u6_n155 ) , .A( u0_u9_u6_n174 ) );
  NOR3_X1 u0_u9_u6_U83 (.A1( u0_u9_u6_n141 ) , .ZN( u0_u9_u6_n154 ) , .A3( u0_u9_u6_n164 ) , .A2( u0_u9_u6_n171 ) );
  AOI211_X1 u0_u9_u6_U84 (.B( u0_u9_u6_n149 ) , .A( u0_u9_u6_n150 ) , .C2( u0_u9_u6_n151 ) , .C1( u0_u9_u6_n152 ) , .ZN( u0_u9_u6_n153 ) );
  OAI211_X1 u0_u9_u6_U85 (.ZN( u0_out9_22 ) , .B( u0_u9_u6_n137 ) , .A( u0_u9_u6_n138 ) , .C2( u0_u9_u6_n139 ) , .C1( u0_u9_u6_n140 ) );
  AOI22_X1 u0_u9_u6_U86 (.B1( u0_u9_u6_n124 ) , .A2( u0_u9_u6_n125 ) , .A1( u0_u9_u6_n126 ) , .ZN( u0_u9_u6_n138 ) , .B2( u0_u9_u6_n161 ) );
  AND4_X1 u0_u9_u6_U87 (.A3( u0_u9_u6_n119 ) , .A1( u0_u9_u6_n120 ) , .A4( u0_u9_u6_n129 ) , .ZN( u0_u9_u6_n140 ) , .A2( u0_u9_u6_n143 ) );
  NAND3_X1 u0_u9_u6_U88 (.A2( u0_u9_u6_n123 ) , .ZN( u0_u9_u6_n125 ) , .A1( u0_u9_u6_n130 ) , .A3( u0_u9_u6_n131 ) );
  NAND3_X1 u0_u9_u6_U89 (.A3( u0_u9_u6_n133 ) , .ZN( u0_u9_u6_n141 ) , .A1( u0_u9_u6_n145 ) , .A2( u0_u9_u6_n148 ) );
  INV_X1 u0_u9_u6_U9 (.ZN( u0_u9_u6_n172 ) , .A( u0_u9_u6_n88 ) );
  NAND3_X1 u0_u9_u6_U90 (.ZN( u0_u9_u6_n101 ) , .A3( u0_u9_u6_n107 ) , .A2( u0_u9_u6_n121 ) , .A1( u0_u9_u6_n127 ) );
  NAND3_X1 u0_u9_u6_U91 (.ZN( u0_u9_u6_n102 ) , .A3( u0_u9_u6_n130 ) , .A2( u0_u9_u6_n145 ) , .A1( u0_u9_u6_n166 ) );
  NAND3_X1 u0_u9_u6_U92 (.A3( u0_u9_u6_n113 ) , .A1( u0_u9_u6_n119 ) , .A2( u0_u9_u6_n123 ) , .ZN( u0_u9_u6_n93 ) );
  NAND3_X1 u0_u9_u6_U93 (.ZN( u0_u9_u6_n142 ) , .A2( u0_u9_u6_n172 ) , .A3( u0_u9_u6_n89 ) , .A1( u0_u9_u6_n90 ) );
  OAI21_X1 u0_uk_U1087 (.ZN( u0_K8_14 ) , .B1( u0_uk_n250 ) , .B2( u0_uk_n329 ) , .A( u0_uk_n760 ) );
  NAND2_X1 u0_uk_U1088 (.A1( u0_uk_K_r6_34 ) , .A2( u0_uk_n202 ) , .ZN( u0_uk_n760 ) );
  INV_X1 u0_uk_U1141 (.ZN( u0_K10_12 ) , .A( u0_uk_n1024 ) );
  INV_X1 u0_uk_U1145 (.ZN( u0_K8_15 ) , .A( u0_uk_n759 ) );
  OAI21_X1 u0_uk_U142 (.ZN( u0_K2_15 ) , .B1( u0_uk_n11 ) , .B2( u0_uk_n597 ) , .A( u0_uk_n865 ) );
  NAND2_X1 u0_uk_U143 (.A1( u0_uk_K_r0_19 ) , .A2( u0_uk_n102 ) , .ZN( u0_uk_n865 ) );
  OAI22_X1 u0_uk_U146 (.ZN( u0_K10_15 ) , .B1( u0_uk_n214 ) , .B2( u0_uk_n229 ) , .A2( u0_uk_n266 ) , .A1( u0_uk_n94 ) );
  INV_X1 u0_uk_U159 (.ZN( u0_K2_19 ) , .A( u0_uk_n864 ) );
  AOI22_X1 u0_uk_U160 (.B2( u0_uk_K_r0_11 ) , .A2( u0_uk_K_r0_47 ) , .A1( u0_uk_n141 ) , .B1( u0_uk_n217 ) , .ZN( u0_uk_n864 ) );
  INV_X1 u0_uk_U187 (.ZN( u0_K2_14 ) , .A( u0_uk_n866 ) );
  AOI22_X1 u0_uk_U188 (.B2( u0_uk_K_r0_11 ) , .A2( u0_uk_K_r0_32 ) , .B1( u0_uk_n142 ) , .A1( u0_uk_n161 ) , .ZN( u0_uk_n866 ) );
  INV_X1 u0_uk_U223 (.ZN( u0_K10_39 ) , .A( u0_uk_n1007 ) );
  AOI22_X1 u0_uk_U224 (.B2( u0_uk_K_r8_44 ) , .A2( u0_uk_K_r8_52 ) , .ZN( u0_uk_n1007 ) , .B1( u0_uk_n141 ) , .A1( u0_uk_n217 ) );
  NAND2_X1 u0_uk_U257 (.A1( u0_uk_K_r11_8 ) , .A2( u0_uk_n141 ) , .ZN( u0_uk_n942 ) );
  OAI22_X1 u0_uk_U278 (.ZN( u0_K10_6 ) , .B1( u0_uk_n102 ) , .A1( u0_uk_n162 ) , .B2( u0_uk_n239 ) , .A2( u0_uk_n267 ) );
  OAI22_X1 u0_uk_U339 (.ZN( u0_K10_4 ) , .A1( u0_uk_n213 ) , .A2( u0_uk_n227 ) , .B2( u0_uk_n246 ) , .B1( u0_uk_n92 ) );
  INV_X1 u0_uk_U355 (.ZN( u0_K10_40 ) , .A( u0_uk_n1006 ) );
  AOI22_X1 u0_uk_U356 (.A2( u0_uk_K_r8_2 ) , .B2( u0_uk_K_r8_22 ) , .ZN( u0_uk_n1006 ) , .B1( u0_uk_n141 ) , .A1( u0_uk_n217 ) );
  OAI21_X1 u0_uk_U393 (.ZN( u0_K10_16 ) , .A( u0_uk_n1022 ) , .B2( u0_uk_n228 ) , .B1( u0_uk_n250 ) );
  NAND2_X1 u0_uk_U394 (.A1( u0_uk_K_r8_32 ) , .ZN( u0_uk_n1022 ) , .A2( u0_uk_n251 ) );
  OAI22_X1 u0_uk_U396 (.ZN( u0_K8_16 ) , .A1( u0_uk_n213 ) , .A2( u0_uk_n344 ) , .B2( u0_uk_n352 ) , .B1( u0_uk_n63 ) );
  INV_X1 u0_uk_U412 (.ZN( u0_K10_37 ) , .A( u0_uk_n1009 ) );
  INV_X1 u0_uk_U416 (.ZN( u0_K10_9 ) , .A( u0_uk_n1005 ) );
  AOI22_X1 u0_uk_U417 (.B2( u0_uk_K_r8_17 ) , .A2( u0_uk_K_r8_27 ) , .ZN( u0_uk_n1005 ) , .B1( u0_uk_n142 ) , .A1( u0_uk_n220 ) );
  OAI22_X1 u0_uk_U431 (.ZN( u0_K2_16 ) , .B1( u0_uk_n240 ) , .A2( u0_uk_n596 ) , .B2( u0_uk_n614 ) , .A1( u0_uk_n94 ) );
  OAI22_X1 u0_uk_U503 (.ZN( u0_K10_17 ) , .B1( u0_uk_n164 ) , .A2( u0_uk_n234 ) , .B2( u0_uk_n262 ) , .A1( u0_uk_n99 ) );
  OAI21_X1 u0_uk_U510 (.ZN( u0_K8_17 ) , .B1( u0_uk_n252 ) , .B2( u0_uk_n336 ) , .A( u0_uk_n758 ) );
  NAND2_X1 u0_uk_U511 (.A1( u0_uk_K_r6_26 ) , .A2( u0_uk_n220 ) , .ZN( u0_uk_n758 ) );
  INV_X1 u0_uk_U564 (.ZN( u0_K10_38 ) , .A( u0_uk_n1008 ) );
  AOI22_X1 u0_uk_U565 (.B2( u0_uk_K_r8_28 ) , .A2( u0_uk_K_r8_8 ) , .ZN( u0_uk_n1008 ) , .B1( u0_uk_n141 ) , .A1( u0_uk_n251 ) );
  OAI22_X1 u0_uk_U598 (.ZN( u0_K8_22 ) , .A1( u0_uk_n257 ) , .A2( u0_uk_n323 ) , .B2( u0_uk_n329 ) , .B1( u0_uk_n92 ) );
  OAI22_X1 u0_uk_U630 (.ZN( u0_K10_11 ) , .A1( u0_uk_n161 ) , .A2( u0_uk_n245 ) , .B2( u0_uk_n262 ) , .B1( u0_uk_n83 ) );
  OAI22_X1 u0_uk_U678 (.ZN( u0_K10_7 ) , .A1( u0_uk_n223 ) , .A2( u0_uk_n234 ) , .B2( u0_uk_n254 ) , .B1( u0_uk_n94 ) );
  OAI21_X1 u0_uk_U714 (.ZN( u0_K10_2 ) , .A( u0_uk_n1015 ) , .B1( u0_uk_n250 ) , .B2( u0_uk_n266 ) );
  NAND2_X1 u0_uk_U715 (.A1( u0_uk_K_r8_41 ) , .ZN( u0_uk_n1015 ) , .A2( u0_uk_n220 ) );
  OAI22_X1 u0_uk_U730 (.ZN( u0_K10_42 ) , .A1( u0_uk_n102 ) , .B1( u0_uk_n238 ) , .A2( u0_uk_n243 ) , .B2( u0_uk_n269 ) );
  OAI22_X1 u0_uk_U753 (.ZN( u0_K8_13 ) , .A1( u0_uk_n109 ) , .B1( u0_uk_n257 ) , .B2( u0_uk_n351 ) , .A2( u0_uk_n357 ) );
  OAI22_X1 u0_uk_U755 (.ZN( u0_K2_13 ) , .B1( u0_uk_n164 ) , .B2( u0_uk_n598 ) , .A2( u0_uk_n627 ) , .A1( u0_uk_n83 ) );
  OAI22_X1 u0_uk_U767 (.ZN( u0_K2_21 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n230 ) , .B2( u0_uk_n620 ) , .A2( u0_uk_n624 ) );
  OAI22_X1 u0_uk_U79 (.ZN( u0_K8_23 ) , .A1( u0_uk_n223 ) , .A2( u0_uk_n340 ) , .B2( u0_uk_n345 ) , .B1( u0_uk_n93 ) );
  OAI21_X1 u0_uk_U812 (.ZN( u0_K8_18 ) , .B2( u0_uk_n331 ) , .A( u0_uk_n757 ) , .B1( u0_uk_n93 ) );
  NAND2_X1 u0_uk_U813 (.A1( u0_uk_K_r6_46 ) , .A2( u0_uk_n10 ) , .ZN( u0_uk_n757 ) );
  OAI22_X1 u0_uk_U814 (.ZN( u0_K2_18 ) , .A1( u0_uk_n230 ) , .A2( u0_uk_n588 ) , .B2( u0_uk_n619 ) , .B1( u0_uk_n63 ) );
  OAI22_X1 u0_uk_U824 (.ZN( u0_K8_20 ) , .B1( u0_uk_n110 ) , .A1( u0_uk_n213 ) , .A2( u0_uk_n331 ) , .B2( u0_uk_n337 ) );
  OAI22_X1 u0_uk_U83 (.ZN( u0_K2_23 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n231 ) , .A2( u0_uk_n589 ) , .B2( u0_uk_n610 ) );
  OAI21_X1 u0_uk_U864 (.ZN( u0_K10_1 ) , .A( u0_uk_n1021 ) , .B2( u0_uk_n258 ) , .B1( u0_uk_n63 ) );
  OAI22_X1 u0_uk_U869 (.ZN( u0_K10_5 ) , .A1( u0_uk_n223 ) , .A2( u0_uk_n246 ) , .B2( u0_uk_n263 ) , .B1( u0_uk_n94 ) );
  OAI22_X1 u0_uk_U894 (.ZN( u0_K10_3 ) , .A2( u0_uk_n235 ) , .A1( u0_uk_n238 ) , .B2( u0_uk_n255 ) , .B1( u0_uk_n93 ) );
  OAI22_X1 u0_uk_U907 (.ZN( u0_K2_24 ) , .A1( u0_uk_n188 ) , .B2( u0_uk_n609 ) , .A2( u0_uk_n624 ) , .B1( u0_uk_n83 ) );
  OAI22_X1 u0_uk_U909 (.ZN( u0_K8_21 ) , .B1( u0_uk_n102 ) , .A1( u0_uk_n257 ) , .A2( u0_uk_n330 ) , .B2( u0_uk_n336 ) );
  OAI22_X1 u0_uk_U917 (.ZN( u0_K2_17 ) , .B1( u0_uk_n100 ) , .A1( u0_uk_n164 ) , .B2( u0_uk_n611 ) , .A2( u0_uk_n627 ) );
  OAI22_X1 u0_uk_U941 (.ZN( u0_K2_20 ) , .A1( u0_uk_n146 ) , .B1( u0_uk_n238 ) , .B2( u0_uk_n596 ) , .A2( u0_uk_n625 ) );
  OAI22_X1 u0_uk_U944 (.ZN( u0_K8_24 ) , .A1( u0_uk_n102 ) , .B1( u0_uk_n213 ) , .A2( u0_uk_n318 ) , .B2( u0_uk_n358 ) );
  OAI22_X1 u0_uk_U956 (.ZN( u0_K10_8 ) , .A1( u0_uk_n109 ) , .B1( u0_uk_n182 ) , .B2( u0_uk_n253 ) , .A2( u0_uk_n267 ) );
  OAI22_X1 u0_uk_U973 (.ZN( u0_K2_22 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n220 ) , .A2( u0_uk_n598 ) , .B2( u0_uk_n615 ) );
  XOR2_X1 u1_U100 (.B( u1_L12_27 ) , .Z( u1_N442 ) , .A( u1_out13_27 ) );
  XOR2_X1 u1_U106 (.B( u1_L12_22 ) , .Z( u1_N437 ) , .A( u1_out13_22 ) );
  XOR2_X1 u1_U107 (.B( u1_L12_21 ) , .Z( u1_N436 ) , .A( u1_out13_21 ) );
  XOR2_X1 u1_U113 (.B( u1_L12_15 ) , .Z( u1_N430 ) , .A( u1_out13_15 ) );
  XOR2_X1 u1_U117 (.B( u1_L12_12 ) , .Z( u1_N427 ) , .A( u1_out13_12 ) );
  XOR2_X1 u1_U122 (.B( u1_L12_7 ) , .Z( u1_N422 ) , .A( u1_out13_7 ) );
  XOR2_X1 u1_U124 (.B( u1_L12_5 ) , .Z( u1_N420 ) , .A( u1_out13_5 ) );
  XOR2_X1 u1_U133 (.B( u1_L11_29 ) , .Z( u1_N412 ) , .A( u1_out12_29 ) );
  XOR2_X1 u1_U138 (.B( u1_L11_25 ) , .Z( u1_N408 ) , .A( u1_out12_25 ) );
  XOR2_X1 u1_U144 (.B( u1_L11_19 ) , .Z( u1_N402 ) , .A( u1_out12_19 ) );
  XOR2_X1 u1_U151 (.B( u1_L11_14 ) , .Z( u1_N397 ) , .A( u1_out12_14 ) );
  XOR2_X1 u1_U154 (.B( u1_L11_11 ) , .Z( u1_N394 ) , .A( u1_out12_11 ) );
  XOR2_X1 u1_U157 (.B( u1_L11_8 ) , .Z( u1_N391 ) , .A( u1_out12_8 ) );
  XOR2_X1 u1_U162 (.B( u1_L11_4 ) , .Z( u1_N387 ) , .A( u1_out12_4 ) );
  XOR2_X1 u1_U163 (.B( u1_L11_3 ) , .Z( u1_N386 ) , .A( u1_out12_3 ) );
  XOR2_X1 u1_U171 (.B( u1_L10_28 ) , .Z( u1_N379 ) , .A( u1_out11_28 ) );
  XOR2_X1 u1_U182 (.B( u1_L10_18 ) , .Z( u1_N369 ) , .A( u1_out11_18 ) );
  XOR2_X1 u1_U187 (.B( u1_L10_13 ) , .Z( u1_N364 ) , .A( u1_out11_13 ) );
  XOR2_X1 u1_U199 (.B( u1_L10_2 ) , .Z( u1_N353 ) , .A( u1_out11_2 ) );
  XOR2_X1 u1_U207 (.B( u1_L9_27 ) , .Z( u1_N346 ) , .A( u1_out10_27 ) );
  XOR2_X1 u1_U208 (.B( u1_L9_26 ) , .Z( u1_N345 ) , .A( u1_out10_26 ) );
  XOR2_X1 u1_U209 (.B( u1_L9_25 ) , .Z( u1_N344 ) , .A( u1_out10_25 ) );
  XOR2_X1 u1_U213 (.B( u1_L9_21 ) , .Z( u1_N340 ) , .A( u1_out10_21 ) );
  XOR2_X1 u1_U215 (.B( u1_L9_20 ) , .Z( u1_N339 ) , .A( u1_out10_20 ) );
  XOR2_X1 u1_U220 (.B( u1_L9_15 ) , .Z( u1_N334 ) , .A( u1_out10_15 ) );
  XOR2_X1 u1_U221 (.B( u1_L9_14 ) , .Z( u1_N333 ) , .A( u1_out10_14 ) );
  XOR2_X1 u1_U226 (.B( u1_L9_10 ) , .Z( u1_N329 ) , .A( u1_out10_10 ) );
  XOR2_X1 u1_U228 (.B( u1_L9_8 ) , .Z( u1_N327 ) , .A( u1_out10_8 ) );
  XOR2_X1 u1_U231 (.B( u1_L9_5 ) , .Z( u1_N324 ) , .A( u1_out10_5 ) );
  XOR2_X1 u1_U233 (.B( u1_L9_3 ) , .Z( u1_N322 ) , .A( u1_out10_3 ) );
  XOR2_X1 u1_U235 (.B( u1_L9_1 ) , .Z( u1_N320 ) , .A( u1_out10_1 ) );
  XOR2_X1 u1_U273 (.B( u1_L7_32 ) , .Z( u1_N287 ) , .A( u1_out8_32 ) );
  XOR2_X1 u1_U276 (.B( u1_L7_29 ) , .Z( u1_N284 ) , .A( u1_out8_29 ) );
  XOR2_X1 u1_U284 (.B( u1_L7_22 ) , .Z( u1_N277 ) , .A( u1_out8_22 ) );
  XOR2_X1 u1_U287 (.B( u1_L7_19 ) , .Z( u1_N274 ) , .A( u1_out8_19 ) );
  XOR2_X1 u1_U295 (.B( u1_L7_12 ) , .Z( u1_N267 ) , .A( u1_out8_12 ) );
  XOR2_X1 u1_U296 (.B( u1_L7_11 ) , .Z( u1_N266 ) , .A( u1_out8_11 ) );
  XOR2_X1 u1_U300 (.B( u1_L7_7 ) , .Z( u1_N262 ) , .A( u1_out8_7 ) );
  XOR2_X1 u1_U304 (.B( u1_L7_4 ) , .Z( u1_N259 ) , .A( u1_out8_4 ) );
  XOR2_X1 u1_U308 (.B( u1_L6_32 ) , .Z( u1_N255 ) , .A( u1_out7_32 ) );
  XOR2_X1 u1_U319 (.B( u1_L6_22 ) , .Z( u1_N245 ) , .A( u1_out7_22 ) );
  XOR2_X1 u1_U330 (.B( u1_L6_12 ) , .Z( u1_N235 ) , .A( u1_out7_12 ) );
  XOR2_X1 u1_U335 (.B( u1_L6_7 ) , .Z( u1_N230 ) , .A( u1_out7_7 ) );
  XOR2_X1 u1_U351 (.B( u1_L5_25 ) , .Z( u1_N216 ) , .A( u1_out6_25 ) );
  XOR2_X1 u1_U363 (.B( u1_L5_14 ) , .Z( u1_N205 ) , .A( u1_out6_14 ) );
  XOR2_X1 u1_U371 (.B( u1_L5_8 ) , .Z( u1_N199 ) , .A( u1_out6_8 ) );
  XOR2_X1 u1_U376 (.B( u1_L5_3 ) , .Z( u1_N194 ) , .A( u1_out6_3 ) );
  XOR2_X1 u1_U95 (.B( u1_L12_32 ) , .Z( u1_N447 ) , .A( u1_out13_32 ) );
  XOR2_X1 u1_u10_U10 (.B( u1_K11_45 ) , .A( u1_R9_30 ) , .Z( u1_u10_X_45 ) );
  XOR2_X1 u1_u10_U11 (.B( u1_K11_44 ) , .A( u1_R9_29 ) , .Z( u1_u10_X_44 ) );
  XOR2_X1 u1_u10_U12 (.B( u1_K11_43 ) , .A( u1_R9_28 ) , .Z( u1_u10_X_43 ) );
  XOR2_X1 u1_u10_U26 (.B( u1_K11_30 ) , .A( u1_R9_21 ) , .Z( u1_u10_X_30 ) );
  XOR2_X1 u1_u10_U28 (.B( u1_K11_29 ) , .A( u1_R9_20 ) , .Z( u1_u10_X_29 ) );
  XOR2_X1 u1_u10_U29 (.B( u1_K11_28 ) , .A( u1_R9_19 ) , .Z( u1_u10_X_28 ) );
  XOR2_X1 u1_u10_U30 (.B( u1_K11_27 ) , .A( u1_R9_18 ) , .Z( u1_u10_X_27 ) );
  XOR2_X1 u1_u10_U31 (.B( u1_K11_26 ) , .A( u1_R9_17 ) , .Z( u1_u10_X_26 ) );
  XOR2_X1 u1_u10_U32 (.B( u1_K11_25 ) , .A( u1_R9_16 ) , .Z( u1_u10_X_25 ) );
  XOR2_X1 u1_u10_U33 (.B( u1_K11_24 ) , .A( u1_R9_17 ) , .Z( u1_u10_X_24 ) );
  XOR2_X1 u1_u10_U34 (.B( u1_K11_23 ) , .A( u1_R9_16 ) , .Z( u1_u10_X_23 ) );
  XOR2_X1 u1_u10_U35 (.B( u1_K11_22 ) , .A( u1_R9_15 ) , .Z( u1_u10_X_22 ) );
  XOR2_X1 u1_u10_U36 (.B( u1_K11_21 ) , .A( u1_R9_14 ) , .Z( u1_u10_X_21 ) );
  XOR2_X1 u1_u10_U37 (.B( u1_K11_20 ) , .A( u1_R9_13 ) , .Z( u1_u10_X_20 ) );
  XOR2_X1 u1_u10_U39 (.B( u1_K11_19 ) , .A( u1_R9_12 ) , .Z( u1_u10_X_19 ) );
  XOR2_X1 u1_u10_U7 (.B( u1_K11_48 ) , .A( u1_R9_1 ) , .Z( u1_u10_X_48 ) );
  XOR2_X1 u1_u10_U8 (.B( u1_K11_47 ) , .A( u1_R9_32 ) , .Z( u1_u10_X_47 ) );
  XOR2_X1 u1_u10_U9 (.B( u1_K11_46 ) , .A( u1_R9_31 ) , .Z( u1_u10_X_46 ) );
  OAI22_X1 u1_u10_u3_U10 (.B1( u1_u10_u3_n113 ) , .A2( u1_u10_u3_n135 ) , .A1( u1_u10_u3_n150 ) , .B2( u1_u10_u3_n164 ) , .ZN( u1_u10_u3_n98 ) );
  OAI211_X1 u1_u10_u3_U11 (.B( u1_u10_u3_n106 ) , .ZN( u1_u10_u3_n119 ) , .C2( u1_u10_u3_n128 ) , .C1( u1_u10_u3_n167 ) , .A( u1_u10_u3_n181 ) );
  AOI221_X1 u1_u10_u3_U12 (.C1( u1_u10_u3_n105 ) , .ZN( u1_u10_u3_n106 ) , .A( u1_u10_u3_n131 ) , .B2( u1_u10_u3_n132 ) , .C2( u1_u10_u3_n133 ) , .B1( u1_u10_u3_n169 ) );
  INV_X1 u1_u10_u3_U13 (.ZN( u1_u10_u3_n181 ) , .A( u1_u10_u3_n98 ) );
  NAND2_X1 u1_u10_u3_U14 (.ZN( u1_u10_u3_n105 ) , .A2( u1_u10_u3_n130 ) , .A1( u1_u10_u3_n155 ) );
  AOI22_X1 u1_u10_u3_U15 (.B1( u1_u10_u3_n115 ) , .A2( u1_u10_u3_n116 ) , .ZN( u1_u10_u3_n123 ) , .B2( u1_u10_u3_n133 ) , .A1( u1_u10_u3_n169 ) );
  NAND2_X1 u1_u10_u3_U16 (.ZN( u1_u10_u3_n116 ) , .A2( u1_u10_u3_n151 ) , .A1( u1_u10_u3_n182 ) );
  NOR2_X1 u1_u10_u3_U17 (.ZN( u1_u10_u3_n126 ) , .A2( u1_u10_u3_n150 ) , .A1( u1_u10_u3_n164 ) );
  AOI21_X1 u1_u10_u3_U18 (.ZN( u1_u10_u3_n112 ) , .B2( u1_u10_u3_n146 ) , .B1( u1_u10_u3_n155 ) , .A( u1_u10_u3_n167 ) );
  NAND2_X1 u1_u10_u3_U19 (.A1( u1_u10_u3_n135 ) , .ZN( u1_u10_u3_n142 ) , .A2( u1_u10_u3_n164 ) );
  NAND2_X1 u1_u10_u3_U20 (.ZN( u1_u10_u3_n132 ) , .A2( u1_u10_u3_n152 ) , .A1( u1_u10_u3_n156 ) );
  AND2_X1 u1_u10_u3_U21 (.A2( u1_u10_u3_n113 ) , .A1( u1_u10_u3_n114 ) , .ZN( u1_u10_u3_n151 ) );
  INV_X1 u1_u10_u3_U22 (.A( u1_u10_u3_n133 ) , .ZN( u1_u10_u3_n165 ) );
  INV_X1 u1_u10_u3_U23 (.A( u1_u10_u3_n135 ) , .ZN( u1_u10_u3_n170 ) );
  NAND2_X1 u1_u10_u3_U24 (.A1( u1_u10_u3_n107 ) , .A2( u1_u10_u3_n108 ) , .ZN( u1_u10_u3_n140 ) );
  NAND2_X1 u1_u10_u3_U25 (.ZN( u1_u10_u3_n117 ) , .A1( u1_u10_u3_n124 ) , .A2( u1_u10_u3_n148 ) );
  NAND2_X1 u1_u10_u3_U26 (.ZN( u1_u10_u3_n143 ) , .A1( u1_u10_u3_n165 ) , .A2( u1_u10_u3_n167 ) );
  INV_X1 u1_u10_u3_U27 (.A( u1_u10_u3_n130 ) , .ZN( u1_u10_u3_n177 ) );
  INV_X1 u1_u10_u3_U28 (.A( u1_u10_u3_n128 ) , .ZN( u1_u10_u3_n176 ) );
  INV_X1 u1_u10_u3_U29 (.A( u1_u10_u3_n155 ) , .ZN( u1_u10_u3_n174 ) );
  INV_X1 u1_u10_u3_U3 (.A( u1_u10_u3_n129 ) , .ZN( u1_u10_u3_n183 ) );
  INV_X1 u1_u10_u3_U30 (.A( u1_u10_u3_n139 ) , .ZN( u1_u10_u3_n185 ) );
  NOR2_X1 u1_u10_u3_U31 (.ZN( u1_u10_u3_n135 ) , .A2( u1_u10_u3_n141 ) , .A1( u1_u10_u3_n169 ) );
  OAI222_X1 u1_u10_u3_U32 (.C2( u1_u10_u3_n107 ) , .A2( u1_u10_u3_n108 ) , .B1( u1_u10_u3_n135 ) , .ZN( u1_u10_u3_n138 ) , .B2( u1_u10_u3_n146 ) , .C1( u1_u10_u3_n154 ) , .A1( u1_u10_u3_n164 ) );
  NOR4_X1 u1_u10_u3_U33 (.A4( u1_u10_u3_n157 ) , .A3( u1_u10_u3_n158 ) , .A2( u1_u10_u3_n159 ) , .A1( u1_u10_u3_n160 ) , .ZN( u1_u10_u3_n161 ) );
  AOI21_X1 u1_u10_u3_U34 (.B2( u1_u10_u3_n152 ) , .B1( u1_u10_u3_n153 ) , .ZN( u1_u10_u3_n158 ) , .A( u1_u10_u3_n164 ) );
  AOI21_X1 u1_u10_u3_U35 (.A( u1_u10_u3_n154 ) , .B2( u1_u10_u3_n155 ) , .B1( u1_u10_u3_n156 ) , .ZN( u1_u10_u3_n157 ) );
  AOI21_X1 u1_u10_u3_U36 (.A( u1_u10_u3_n149 ) , .B2( u1_u10_u3_n150 ) , .B1( u1_u10_u3_n151 ) , .ZN( u1_u10_u3_n159 ) );
  AOI211_X1 u1_u10_u3_U37 (.ZN( u1_u10_u3_n109 ) , .A( u1_u10_u3_n119 ) , .C2( u1_u10_u3_n129 ) , .B( u1_u10_u3_n138 ) , .C1( u1_u10_u3_n141 ) );
  AOI211_X1 u1_u10_u3_U38 (.B( u1_u10_u3_n119 ) , .A( u1_u10_u3_n120 ) , .C2( u1_u10_u3_n121 ) , .ZN( u1_u10_u3_n122 ) , .C1( u1_u10_u3_n179 ) );
  INV_X1 u1_u10_u3_U39 (.A( u1_u10_u3_n156 ) , .ZN( u1_u10_u3_n179 ) );
  INV_X1 u1_u10_u3_U4 (.A( u1_u10_u3_n140 ) , .ZN( u1_u10_u3_n182 ) );
  OAI22_X1 u1_u10_u3_U40 (.B1( u1_u10_u3_n118 ) , .ZN( u1_u10_u3_n120 ) , .A1( u1_u10_u3_n135 ) , .B2( u1_u10_u3_n154 ) , .A2( u1_u10_u3_n178 ) );
  AND3_X1 u1_u10_u3_U41 (.ZN( u1_u10_u3_n118 ) , .A2( u1_u10_u3_n124 ) , .A1( u1_u10_u3_n144 ) , .A3( u1_u10_u3_n152 ) );
  INV_X1 u1_u10_u3_U42 (.A( u1_u10_u3_n121 ) , .ZN( u1_u10_u3_n164 ) );
  NAND2_X1 u1_u10_u3_U43 (.ZN( u1_u10_u3_n133 ) , .A1( u1_u10_u3_n154 ) , .A2( u1_u10_u3_n164 ) );
  OAI211_X1 u1_u10_u3_U44 (.B( u1_u10_u3_n127 ) , .ZN( u1_u10_u3_n139 ) , .C1( u1_u10_u3_n150 ) , .C2( u1_u10_u3_n154 ) , .A( u1_u10_u3_n184 ) );
  INV_X1 u1_u10_u3_U45 (.A( u1_u10_u3_n125 ) , .ZN( u1_u10_u3_n184 ) );
  AOI221_X1 u1_u10_u3_U46 (.A( u1_u10_u3_n126 ) , .ZN( u1_u10_u3_n127 ) , .C2( u1_u10_u3_n132 ) , .C1( u1_u10_u3_n169 ) , .B2( u1_u10_u3_n170 ) , .B1( u1_u10_u3_n174 ) );
  OAI22_X1 u1_u10_u3_U47 (.A1( u1_u10_u3_n124 ) , .ZN( u1_u10_u3_n125 ) , .B2( u1_u10_u3_n145 ) , .A2( u1_u10_u3_n165 ) , .B1( u1_u10_u3_n167 ) );
  NOR2_X1 u1_u10_u3_U48 (.A1( u1_u10_u3_n113 ) , .ZN( u1_u10_u3_n131 ) , .A2( u1_u10_u3_n154 ) );
  NAND2_X1 u1_u10_u3_U49 (.A1( u1_u10_u3_n103 ) , .ZN( u1_u10_u3_n150 ) , .A2( u1_u10_u3_n99 ) );
  INV_X1 u1_u10_u3_U5 (.A( u1_u10_u3_n117 ) , .ZN( u1_u10_u3_n178 ) );
  NAND2_X1 u1_u10_u3_U50 (.A2( u1_u10_u3_n102 ) , .ZN( u1_u10_u3_n155 ) , .A1( u1_u10_u3_n97 ) );
  INV_X1 u1_u10_u3_U51 (.A( u1_u10_u3_n141 ) , .ZN( u1_u10_u3_n167 ) );
  AOI21_X1 u1_u10_u3_U52 (.B2( u1_u10_u3_n114 ) , .B1( u1_u10_u3_n146 ) , .A( u1_u10_u3_n154 ) , .ZN( u1_u10_u3_n94 ) );
  AOI21_X1 u1_u10_u3_U53 (.ZN( u1_u10_u3_n110 ) , .B2( u1_u10_u3_n142 ) , .B1( u1_u10_u3_n186 ) , .A( u1_u10_u3_n95 ) );
  INV_X1 u1_u10_u3_U54 (.A( u1_u10_u3_n145 ) , .ZN( u1_u10_u3_n186 ) );
  AOI21_X1 u1_u10_u3_U55 (.B1( u1_u10_u3_n124 ) , .A( u1_u10_u3_n149 ) , .B2( u1_u10_u3_n155 ) , .ZN( u1_u10_u3_n95 ) );
  INV_X1 u1_u10_u3_U56 (.A( u1_u10_u3_n149 ) , .ZN( u1_u10_u3_n169 ) );
  NAND2_X1 u1_u10_u3_U57 (.ZN( u1_u10_u3_n124 ) , .A1( u1_u10_u3_n96 ) , .A2( u1_u10_u3_n97 ) );
  NAND2_X1 u1_u10_u3_U58 (.A2( u1_u10_u3_n100 ) , .ZN( u1_u10_u3_n146 ) , .A1( u1_u10_u3_n96 ) );
  NAND2_X1 u1_u10_u3_U59 (.A1( u1_u10_u3_n101 ) , .ZN( u1_u10_u3_n145 ) , .A2( u1_u10_u3_n99 ) );
  AOI221_X1 u1_u10_u3_U6 (.A( u1_u10_u3_n131 ) , .C2( u1_u10_u3_n132 ) , .C1( u1_u10_u3_n133 ) , .ZN( u1_u10_u3_n134 ) , .B1( u1_u10_u3_n143 ) , .B2( u1_u10_u3_n177 ) );
  NAND2_X1 u1_u10_u3_U60 (.A1( u1_u10_u3_n100 ) , .ZN( u1_u10_u3_n156 ) , .A2( u1_u10_u3_n99 ) );
  NAND2_X1 u1_u10_u3_U61 (.A2( u1_u10_u3_n101 ) , .A1( u1_u10_u3_n104 ) , .ZN( u1_u10_u3_n148 ) );
  NAND2_X1 u1_u10_u3_U62 (.A1( u1_u10_u3_n100 ) , .A2( u1_u10_u3_n102 ) , .ZN( u1_u10_u3_n128 ) );
  NAND2_X1 u1_u10_u3_U63 (.A2( u1_u10_u3_n101 ) , .A1( u1_u10_u3_n102 ) , .ZN( u1_u10_u3_n152 ) );
  NAND2_X1 u1_u10_u3_U64 (.A2( u1_u10_u3_n101 ) , .ZN( u1_u10_u3_n114 ) , .A1( u1_u10_u3_n96 ) );
  NAND2_X1 u1_u10_u3_U65 (.ZN( u1_u10_u3_n107 ) , .A1( u1_u10_u3_n97 ) , .A2( u1_u10_u3_n99 ) );
  NAND2_X1 u1_u10_u3_U66 (.A2( u1_u10_u3_n100 ) , .A1( u1_u10_u3_n104 ) , .ZN( u1_u10_u3_n113 ) );
  NAND2_X1 u1_u10_u3_U67 (.A1( u1_u10_u3_n104 ) , .ZN( u1_u10_u3_n153 ) , .A2( u1_u10_u3_n97 ) );
  NAND2_X1 u1_u10_u3_U68 (.A2( u1_u10_u3_n103 ) , .A1( u1_u10_u3_n104 ) , .ZN( u1_u10_u3_n130 ) );
  NAND2_X1 u1_u10_u3_U69 (.A2( u1_u10_u3_n103 ) , .ZN( u1_u10_u3_n144 ) , .A1( u1_u10_u3_n96 ) );
  OAI22_X1 u1_u10_u3_U7 (.B2( u1_u10_u3_n147 ) , .A2( u1_u10_u3_n148 ) , .ZN( u1_u10_u3_n160 ) , .B1( u1_u10_u3_n165 ) , .A1( u1_u10_u3_n168 ) );
  NAND2_X1 u1_u10_u3_U70 (.A1( u1_u10_u3_n102 ) , .A2( u1_u10_u3_n103 ) , .ZN( u1_u10_u3_n108 ) );
  NOR2_X1 u1_u10_u3_U71 (.A2( u1_u10_X_19 ) , .A1( u1_u10_X_20 ) , .ZN( u1_u10_u3_n99 ) );
  NOR2_X1 u1_u10_u3_U72 (.A2( u1_u10_X_21 ) , .A1( u1_u10_X_24 ) , .ZN( u1_u10_u3_n103 ) );
  NOR2_X1 u1_u10_u3_U73 (.A2( u1_u10_X_24 ) , .A1( u1_u10_u3_n171 ) , .ZN( u1_u10_u3_n97 ) );
  NOR2_X1 u1_u10_u3_U74 (.A2( u1_u10_X_23 ) , .ZN( u1_u10_u3_n141 ) , .A1( u1_u10_u3_n166 ) );
  NOR2_X1 u1_u10_u3_U75 (.A2( u1_u10_X_19 ) , .A1( u1_u10_u3_n172 ) , .ZN( u1_u10_u3_n96 ) );
  NAND2_X1 u1_u10_u3_U76 (.A1( u1_u10_X_22 ) , .A2( u1_u10_X_23 ) , .ZN( u1_u10_u3_n154 ) );
  NAND2_X1 u1_u10_u3_U77 (.A1( u1_u10_X_23 ) , .ZN( u1_u10_u3_n149 ) , .A2( u1_u10_u3_n166 ) );
  NOR2_X1 u1_u10_u3_U78 (.A2( u1_u10_X_22 ) , .A1( u1_u10_X_23 ) , .ZN( u1_u10_u3_n121 ) );
  AND2_X1 u1_u10_u3_U79 (.A1( u1_u10_X_24 ) , .ZN( u1_u10_u3_n101 ) , .A2( u1_u10_u3_n171 ) );
  AND3_X1 u1_u10_u3_U8 (.A3( u1_u10_u3_n144 ) , .A2( u1_u10_u3_n145 ) , .A1( u1_u10_u3_n146 ) , .ZN( u1_u10_u3_n147 ) );
  AND2_X1 u1_u10_u3_U80 (.A1( u1_u10_X_19 ) , .ZN( u1_u10_u3_n102 ) , .A2( u1_u10_u3_n172 ) );
  AND2_X1 u1_u10_u3_U81 (.A1( u1_u10_X_21 ) , .A2( u1_u10_X_24 ) , .ZN( u1_u10_u3_n100 ) );
  AND2_X1 u1_u10_u3_U82 (.A2( u1_u10_X_19 ) , .A1( u1_u10_X_20 ) , .ZN( u1_u10_u3_n104 ) );
  INV_X1 u1_u10_u3_U83 (.A( u1_u10_X_22 ) , .ZN( u1_u10_u3_n166 ) );
  INV_X1 u1_u10_u3_U84 (.A( u1_u10_X_21 ) , .ZN( u1_u10_u3_n171 ) );
  INV_X1 u1_u10_u3_U85 (.A( u1_u10_X_20 ) , .ZN( u1_u10_u3_n172 ) );
  OR4_X1 u1_u10_u3_U86 (.ZN( u1_out10_10 ) , .A4( u1_u10_u3_n136 ) , .A3( u1_u10_u3_n137 ) , .A1( u1_u10_u3_n138 ) , .A2( u1_u10_u3_n139 ) );
  OAI222_X1 u1_u10_u3_U87 (.C1( u1_u10_u3_n128 ) , .ZN( u1_u10_u3_n137 ) , .B1( u1_u10_u3_n148 ) , .A2( u1_u10_u3_n150 ) , .B2( u1_u10_u3_n154 ) , .C2( u1_u10_u3_n164 ) , .A1( u1_u10_u3_n167 ) );
  OAI221_X1 u1_u10_u3_U88 (.A( u1_u10_u3_n134 ) , .B2( u1_u10_u3_n135 ) , .ZN( u1_u10_u3_n136 ) , .C1( u1_u10_u3_n149 ) , .B1( u1_u10_u3_n151 ) , .C2( u1_u10_u3_n183 ) );
  NAND4_X1 u1_u10_u3_U89 (.ZN( u1_out10_26 ) , .A4( u1_u10_u3_n109 ) , .A3( u1_u10_u3_n110 ) , .A2( u1_u10_u3_n111 ) , .A1( u1_u10_u3_n173 ) );
  INV_X1 u1_u10_u3_U9 (.A( u1_u10_u3_n143 ) , .ZN( u1_u10_u3_n168 ) );
  INV_X1 u1_u10_u3_U90 (.ZN( u1_u10_u3_n173 ) , .A( u1_u10_u3_n94 ) );
  OAI21_X1 u1_u10_u3_U91 (.ZN( u1_u10_u3_n111 ) , .B2( u1_u10_u3_n117 ) , .A( u1_u10_u3_n133 ) , .B1( u1_u10_u3_n176 ) );
  NAND4_X1 u1_u10_u3_U92 (.ZN( u1_out10_20 ) , .A4( u1_u10_u3_n122 ) , .A3( u1_u10_u3_n123 ) , .A1( u1_u10_u3_n175 ) , .A2( u1_u10_u3_n180 ) );
  INV_X1 u1_u10_u3_U93 (.A( u1_u10_u3_n126 ) , .ZN( u1_u10_u3_n180 ) );
  INV_X1 u1_u10_u3_U94 (.A( u1_u10_u3_n112 ) , .ZN( u1_u10_u3_n175 ) );
  NAND4_X1 u1_u10_u3_U95 (.ZN( u1_out10_1 ) , .A4( u1_u10_u3_n161 ) , .A3( u1_u10_u3_n162 ) , .A2( u1_u10_u3_n163 ) , .A1( u1_u10_u3_n185 ) );
  NAND2_X1 u1_u10_u3_U96 (.ZN( u1_u10_u3_n163 ) , .A2( u1_u10_u3_n170 ) , .A1( u1_u10_u3_n176 ) );
  AOI22_X1 u1_u10_u3_U97 (.B2( u1_u10_u3_n140 ) , .B1( u1_u10_u3_n141 ) , .A2( u1_u10_u3_n142 ) , .ZN( u1_u10_u3_n162 ) , .A1( u1_u10_u3_n177 ) );
  NAND3_X1 u1_u10_u3_U98 (.A1( u1_u10_u3_n114 ) , .ZN( u1_u10_u3_n115 ) , .A2( u1_u10_u3_n145 ) , .A3( u1_u10_u3_n153 ) );
  NAND3_X1 u1_u10_u3_U99 (.ZN( u1_u10_u3_n129 ) , .A2( u1_u10_u3_n144 ) , .A1( u1_u10_u3_n153 ) , .A3( u1_u10_u3_n182 ) );
  OAI22_X1 u1_u10_u4_U10 (.B2( u1_u10_u4_n135 ) , .ZN( u1_u10_u4_n137 ) , .B1( u1_u10_u4_n153 ) , .A1( u1_u10_u4_n155 ) , .A2( u1_u10_u4_n171 ) );
  AND3_X1 u1_u10_u4_U11 (.A2( u1_u10_u4_n134 ) , .ZN( u1_u10_u4_n135 ) , .A3( u1_u10_u4_n145 ) , .A1( u1_u10_u4_n157 ) );
  NAND2_X1 u1_u10_u4_U12 (.ZN( u1_u10_u4_n132 ) , .A2( u1_u10_u4_n170 ) , .A1( u1_u10_u4_n173 ) );
  AOI21_X1 u1_u10_u4_U13 (.B2( u1_u10_u4_n160 ) , .B1( u1_u10_u4_n161 ) , .ZN( u1_u10_u4_n162 ) , .A( u1_u10_u4_n170 ) );
  AOI21_X1 u1_u10_u4_U14 (.ZN( u1_u10_u4_n107 ) , .B2( u1_u10_u4_n143 ) , .A( u1_u10_u4_n174 ) , .B1( u1_u10_u4_n184 ) );
  AOI21_X1 u1_u10_u4_U15 (.B2( u1_u10_u4_n158 ) , .B1( u1_u10_u4_n159 ) , .ZN( u1_u10_u4_n163 ) , .A( u1_u10_u4_n174 ) );
  AOI21_X1 u1_u10_u4_U16 (.A( u1_u10_u4_n153 ) , .B2( u1_u10_u4_n154 ) , .B1( u1_u10_u4_n155 ) , .ZN( u1_u10_u4_n165 ) );
  AOI21_X1 u1_u10_u4_U17 (.A( u1_u10_u4_n156 ) , .B2( u1_u10_u4_n157 ) , .ZN( u1_u10_u4_n164 ) , .B1( u1_u10_u4_n184 ) );
  INV_X1 u1_u10_u4_U18 (.A( u1_u10_u4_n138 ) , .ZN( u1_u10_u4_n170 ) );
  AND2_X1 u1_u10_u4_U19 (.A2( u1_u10_u4_n120 ) , .ZN( u1_u10_u4_n155 ) , .A1( u1_u10_u4_n160 ) );
  INV_X1 u1_u10_u4_U20 (.A( u1_u10_u4_n156 ) , .ZN( u1_u10_u4_n175 ) );
  NAND2_X1 u1_u10_u4_U21 (.A2( u1_u10_u4_n118 ) , .ZN( u1_u10_u4_n131 ) , .A1( u1_u10_u4_n147 ) );
  NAND2_X1 u1_u10_u4_U22 (.A1( u1_u10_u4_n119 ) , .A2( u1_u10_u4_n120 ) , .ZN( u1_u10_u4_n130 ) );
  NAND2_X1 u1_u10_u4_U23 (.ZN( u1_u10_u4_n117 ) , .A2( u1_u10_u4_n118 ) , .A1( u1_u10_u4_n148 ) );
  NAND2_X1 u1_u10_u4_U24 (.ZN( u1_u10_u4_n129 ) , .A1( u1_u10_u4_n134 ) , .A2( u1_u10_u4_n148 ) );
  AND3_X1 u1_u10_u4_U25 (.A1( u1_u10_u4_n119 ) , .A2( u1_u10_u4_n143 ) , .A3( u1_u10_u4_n154 ) , .ZN( u1_u10_u4_n161 ) );
  AND2_X1 u1_u10_u4_U26 (.A1( u1_u10_u4_n145 ) , .A2( u1_u10_u4_n147 ) , .ZN( u1_u10_u4_n159 ) );
  OR3_X1 u1_u10_u4_U27 (.A3( u1_u10_u4_n114 ) , .A2( u1_u10_u4_n115 ) , .A1( u1_u10_u4_n116 ) , .ZN( u1_u10_u4_n136 ) );
  AOI21_X1 u1_u10_u4_U28 (.A( u1_u10_u4_n113 ) , .ZN( u1_u10_u4_n116 ) , .B2( u1_u10_u4_n173 ) , .B1( u1_u10_u4_n174 ) );
  AOI21_X1 u1_u10_u4_U29 (.ZN( u1_u10_u4_n115 ) , .B2( u1_u10_u4_n145 ) , .B1( u1_u10_u4_n146 ) , .A( u1_u10_u4_n156 ) );
  NOR2_X1 u1_u10_u4_U3 (.ZN( u1_u10_u4_n121 ) , .A1( u1_u10_u4_n181 ) , .A2( u1_u10_u4_n182 ) );
  OAI22_X1 u1_u10_u4_U30 (.ZN( u1_u10_u4_n114 ) , .A2( u1_u10_u4_n121 ) , .B1( u1_u10_u4_n160 ) , .B2( u1_u10_u4_n170 ) , .A1( u1_u10_u4_n171 ) );
  INV_X1 u1_u10_u4_U31 (.A( u1_u10_u4_n158 ) , .ZN( u1_u10_u4_n182 ) );
  INV_X1 u1_u10_u4_U32 (.ZN( u1_u10_u4_n181 ) , .A( u1_u10_u4_n96 ) );
  INV_X1 u1_u10_u4_U33 (.A( u1_u10_u4_n144 ) , .ZN( u1_u10_u4_n179 ) );
  INV_X1 u1_u10_u4_U34 (.A( u1_u10_u4_n157 ) , .ZN( u1_u10_u4_n178 ) );
  NAND2_X1 u1_u10_u4_U35 (.A2( u1_u10_u4_n154 ) , .A1( u1_u10_u4_n96 ) , .ZN( u1_u10_u4_n97 ) );
  INV_X1 u1_u10_u4_U36 (.ZN( u1_u10_u4_n186 ) , .A( u1_u10_u4_n95 ) );
  OAI221_X1 u1_u10_u4_U37 (.C1( u1_u10_u4_n134 ) , .B1( u1_u10_u4_n158 ) , .B2( u1_u10_u4_n171 ) , .C2( u1_u10_u4_n173 ) , .A( u1_u10_u4_n94 ) , .ZN( u1_u10_u4_n95 ) );
  AOI222_X1 u1_u10_u4_U38 (.B2( u1_u10_u4_n132 ) , .A1( u1_u10_u4_n138 ) , .C2( u1_u10_u4_n175 ) , .A2( u1_u10_u4_n179 ) , .C1( u1_u10_u4_n181 ) , .B1( u1_u10_u4_n185 ) , .ZN( u1_u10_u4_n94 ) );
  INV_X1 u1_u10_u4_U39 (.A( u1_u10_u4_n113 ) , .ZN( u1_u10_u4_n185 ) );
  INV_X1 u1_u10_u4_U4 (.A( u1_u10_u4_n117 ) , .ZN( u1_u10_u4_n184 ) );
  INV_X1 u1_u10_u4_U40 (.A( u1_u10_u4_n143 ) , .ZN( u1_u10_u4_n183 ) );
  NOR2_X1 u1_u10_u4_U41 (.ZN( u1_u10_u4_n138 ) , .A1( u1_u10_u4_n168 ) , .A2( u1_u10_u4_n169 ) );
  NOR2_X1 u1_u10_u4_U42 (.A1( u1_u10_u4_n150 ) , .A2( u1_u10_u4_n152 ) , .ZN( u1_u10_u4_n153 ) );
  NOR2_X1 u1_u10_u4_U43 (.A2( u1_u10_u4_n128 ) , .A1( u1_u10_u4_n138 ) , .ZN( u1_u10_u4_n156 ) );
  AOI22_X1 u1_u10_u4_U44 (.B2( u1_u10_u4_n122 ) , .A1( u1_u10_u4_n123 ) , .ZN( u1_u10_u4_n124 ) , .B1( u1_u10_u4_n128 ) , .A2( u1_u10_u4_n172 ) );
  INV_X1 u1_u10_u4_U45 (.A( u1_u10_u4_n153 ) , .ZN( u1_u10_u4_n172 ) );
  NAND2_X1 u1_u10_u4_U46 (.A2( u1_u10_u4_n120 ) , .ZN( u1_u10_u4_n123 ) , .A1( u1_u10_u4_n161 ) );
  AOI22_X1 u1_u10_u4_U47 (.B2( u1_u10_u4_n132 ) , .A2( u1_u10_u4_n133 ) , .ZN( u1_u10_u4_n140 ) , .A1( u1_u10_u4_n150 ) , .B1( u1_u10_u4_n179 ) );
  NAND2_X1 u1_u10_u4_U48 (.ZN( u1_u10_u4_n133 ) , .A2( u1_u10_u4_n146 ) , .A1( u1_u10_u4_n154 ) );
  NAND2_X1 u1_u10_u4_U49 (.A1( u1_u10_u4_n103 ) , .ZN( u1_u10_u4_n154 ) , .A2( u1_u10_u4_n98 ) );
  NOR4_X1 u1_u10_u4_U5 (.A4( u1_u10_u4_n106 ) , .A3( u1_u10_u4_n107 ) , .A2( u1_u10_u4_n108 ) , .A1( u1_u10_u4_n109 ) , .ZN( u1_u10_u4_n110 ) );
  NAND2_X1 u1_u10_u4_U50 (.A1( u1_u10_u4_n101 ) , .ZN( u1_u10_u4_n158 ) , .A2( u1_u10_u4_n99 ) );
  AOI21_X1 u1_u10_u4_U51 (.ZN( u1_u10_u4_n127 ) , .A( u1_u10_u4_n136 ) , .B2( u1_u10_u4_n150 ) , .B1( u1_u10_u4_n180 ) );
  INV_X1 u1_u10_u4_U52 (.A( u1_u10_u4_n160 ) , .ZN( u1_u10_u4_n180 ) );
  NAND2_X1 u1_u10_u4_U53 (.A2( u1_u10_u4_n104 ) , .A1( u1_u10_u4_n105 ) , .ZN( u1_u10_u4_n146 ) );
  NAND2_X1 u1_u10_u4_U54 (.A2( u1_u10_u4_n101 ) , .A1( u1_u10_u4_n102 ) , .ZN( u1_u10_u4_n160 ) );
  NAND2_X1 u1_u10_u4_U55 (.ZN( u1_u10_u4_n134 ) , .A1( u1_u10_u4_n98 ) , .A2( u1_u10_u4_n99 ) );
  NAND2_X1 u1_u10_u4_U56 (.A1( u1_u10_u4_n103 ) , .A2( u1_u10_u4_n104 ) , .ZN( u1_u10_u4_n143 ) );
  NAND2_X1 u1_u10_u4_U57 (.A2( u1_u10_u4_n105 ) , .ZN( u1_u10_u4_n145 ) , .A1( u1_u10_u4_n98 ) );
  NAND2_X1 u1_u10_u4_U58 (.A1( u1_u10_u4_n100 ) , .A2( u1_u10_u4_n105 ) , .ZN( u1_u10_u4_n120 ) );
  NAND2_X1 u1_u10_u4_U59 (.A1( u1_u10_u4_n102 ) , .A2( u1_u10_u4_n104 ) , .ZN( u1_u10_u4_n148 ) );
  AOI21_X1 u1_u10_u4_U6 (.ZN( u1_u10_u4_n106 ) , .B2( u1_u10_u4_n146 ) , .B1( u1_u10_u4_n158 ) , .A( u1_u10_u4_n170 ) );
  NAND2_X1 u1_u10_u4_U60 (.A2( u1_u10_u4_n100 ) , .A1( u1_u10_u4_n103 ) , .ZN( u1_u10_u4_n157 ) );
  INV_X1 u1_u10_u4_U61 (.A( u1_u10_u4_n150 ) , .ZN( u1_u10_u4_n173 ) );
  INV_X1 u1_u10_u4_U62 (.A( u1_u10_u4_n152 ) , .ZN( u1_u10_u4_n171 ) );
  NAND2_X1 u1_u10_u4_U63 (.A1( u1_u10_u4_n100 ) , .ZN( u1_u10_u4_n118 ) , .A2( u1_u10_u4_n99 ) );
  NAND2_X1 u1_u10_u4_U64 (.A2( u1_u10_u4_n100 ) , .A1( u1_u10_u4_n102 ) , .ZN( u1_u10_u4_n144 ) );
  NAND2_X1 u1_u10_u4_U65 (.A2( u1_u10_u4_n101 ) , .A1( u1_u10_u4_n105 ) , .ZN( u1_u10_u4_n96 ) );
  INV_X1 u1_u10_u4_U66 (.A( u1_u10_u4_n128 ) , .ZN( u1_u10_u4_n174 ) );
  NAND2_X1 u1_u10_u4_U67 (.A2( u1_u10_u4_n102 ) , .ZN( u1_u10_u4_n119 ) , .A1( u1_u10_u4_n98 ) );
  NAND2_X1 u1_u10_u4_U68 (.A2( u1_u10_u4_n101 ) , .A1( u1_u10_u4_n103 ) , .ZN( u1_u10_u4_n147 ) );
  NAND2_X1 u1_u10_u4_U69 (.A2( u1_u10_u4_n104 ) , .ZN( u1_u10_u4_n113 ) , .A1( u1_u10_u4_n99 ) );
  AOI21_X1 u1_u10_u4_U7 (.ZN( u1_u10_u4_n108 ) , .B2( u1_u10_u4_n134 ) , .B1( u1_u10_u4_n155 ) , .A( u1_u10_u4_n156 ) );
  NOR2_X1 u1_u10_u4_U70 (.A2( u1_u10_X_28 ) , .ZN( u1_u10_u4_n150 ) , .A1( u1_u10_u4_n168 ) );
  NOR2_X1 u1_u10_u4_U71 (.A2( u1_u10_X_29 ) , .ZN( u1_u10_u4_n152 ) , .A1( u1_u10_u4_n169 ) );
  NOR2_X1 u1_u10_u4_U72 (.A2( u1_u10_X_30 ) , .ZN( u1_u10_u4_n105 ) , .A1( u1_u10_u4_n176 ) );
  NOR2_X1 u1_u10_u4_U73 (.A2( u1_u10_X_26 ) , .ZN( u1_u10_u4_n100 ) , .A1( u1_u10_u4_n177 ) );
  NOR2_X1 u1_u10_u4_U74 (.A2( u1_u10_X_28 ) , .A1( u1_u10_X_29 ) , .ZN( u1_u10_u4_n128 ) );
  NOR2_X1 u1_u10_u4_U75 (.A2( u1_u10_X_27 ) , .A1( u1_u10_X_30 ) , .ZN( u1_u10_u4_n102 ) );
  NOR2_X1 u1_u10_u4_U76 (.A2( u1_u10_X_25 ) , .A1( u1_u10_X_26 ) , .ZN( u1_u10_u4_n98 ) );
  AND2_X1 u1_u10_u4_U77 (.A2( u1_u10_X_25 ) , .A1( u1_u10_X_26 ) , .ZN( u1_u10_u4_n104 ) );
  AND2_X1 u1_u10_u4_U78 (.A1( u1_u10_X_30 ) , .A2( u1_u10_u4_n176 ) , .ZN( u1_u10_u4_n99 ) );
  AND2_X1 u1_u10_u4_U79 (.A1( u1_u10_X_26 ) , .ZN( u1_u10_u4_n101 ) , .A2( u1_u10_u4_n177 ) );
  AOI21_X1 u1_u10_u4_U8 (.ZN( u1_u10_u4_n109 ) , .A( u1_u10_u4_n153 ) , .B1( u1_u10_u4_n159 ) , .B2( u1_u10_u4_n184 ) );
  AND2_X1 u1_u10_u4_U80 (.A1( u1_u10_X_27 ) , .A2( u1_u10_X_30 ) , .ZN( u1_u10_u4_n103 ) );
  INV_X1 u1_u10_u4_U81 (.A( u1_u10_X_28 ) , .ZN( u1_u10_u4_n169 ) );
  INV_X1 u1_u10_u4_U82 (.A( u1_u10_X_29 ) , .ZN( u1_u10_u4_n168 ) );
  INV_X1 u1_u10_u4_U83 (.A( u1_u10_X_25 ) , .ZN( u1_u10_u4_n177 ) );
  INV_X1 u1_u10_u4_U84 (.A( u1_u10_X_27 ) , .ZN( u1_u10_u4_n176 ) );
  NAND4_X1 u1_u10_u4_U85 (.ZN( u1_out10_25 ) , .A4( u1_u10_u4_n139 ) , .A3( u1_u10_u4_n140 ) , .A2( u1_u10_u4_n141 ) , .A1( u1_u10_u4_n142 ) );
  OAI21_X1 u1_u10_u4_U86 (.A( u1_u10_u4_n128 ) , .B2( u1_u10_u4_n129 ) , .B1( u1_u10_u4_n130 ) , .ZN( u1_u10_u4_n142 ) );
  OAI21_X1 u1_u10_u4_U87 (.B2( u1_u10_u4_n131 ) , .ZN( u1_u10_u4_n141 ) , .A( u1_u10_u4_n175 ) , .B1( u1_u10_u4_n183 ) );
  NAND4_X1 u1_u10_u4_U88 (.ZN( u1_out10_14 ) , .A4( u1_u10_u4_n124 ) , .A3( u1_u10_u4_n125 ) , .A2( u1_u10_u4_n126 ) , .A1( u1_u10_u4_n127 ) );
  AOI22_X1 u1_u10_u4_U89 (.B2( u1_u10_u4_n117 ) , .ZN( u1_u10_u4_n126 ) , .A1( u1_u10_u4_n129 ) , .B1( u1_u10_u4_n152 ) , .A2( u1_u10_u4_n175 ) );
  AOI211_X1 u1_u10_u4_U9 (.B( u1_u10_u4_n136 ) , .A( u1_u10_u4_n137 ) , .C2( u1_u10_u4_n138 ) , .ZN( u1_u10_u4_n139 ) , .C1( u1_u10_u4_n182 ) );
  AOI22_X1 u1_u10_u4_U90 (.ZN( u1_u10_u4_n125 ) , .B2( u1_u10_u4_n131 ) , .A2( u1_u10_u4_n132 ) , .B1( u1_u10_u4_n138 ) , .A1( u1_u10_u4_n178 ) );
  NAND4_X1 u1_u10_u4_U91 (.ZN( u1_out10_8 ) , .A4( u1_u10_u4_n110 ) , .A3( u1_u10_u4_n111 ) , .A2( u1_u10_u4_n112 ) , .A1( u1_u10_u4_n186 ) );
  NAND2_X1 u1_u10_u4_U92 (.ZN( u1_u10_u4_n112 ) , .A2( u1_u10_u4_n130 ) , .A1( u1_u10_u4_n150 ) );
  AOI22_X1 u1_u10_u4_U93 (.ZN( u1_u10_u4_n111 ) , .B2( u1_u10_u4_n132 ) , .A1( u1_u10_u4_n152 ) , .B1( u1_u10_u4_n178 ) , .A2( u1_u10_u4_n97 ) );
  AOI22_X1 u1_u10_u4_U94 (.B2( u1_u10_u4_n149 ) , .B1( u1_u10_u4_n150 ) , .A2( u1_u10_u4_n151 ) , .A1( u1_u10_u4_n152 ) , .ZN( u1_u10_u4_n167 ) );
  NOR4_X1 u1_u10_u4_U95 (.A4( u1_u10_u4_n162 ) , .A3( u1_u10_u4_n163 ) , .A2( u1_u10_u4_n164 ) , .A1( u1_u10_u4_n165 ) , .ZN( u1_u10_u4_n166 ) );
  NAND3_X1 u1_u10_u4_U96 (.ZN( u1_out10_3 ) , .A3( u1_u10_u4_n166 ) , .A1( u1_u10_u4_n167 ) , .A2( u1_u10_u4_n186 ) );
  NAND3_X1 u1_u10_u4_U97 (.A3( u1_u10_u4_n146 ) , .A2( u1_u10_u4_n147 ) , .A1( u1_u10_u4_n148 ) , .ZN( u1_u10_u4_n149 ) );
  NAND3_X1 u1_u10_u4_U98 (.A3( u1_u10_u4_n143 ) , .A2( u1_u10_u4_n144 ) , .A1( u1_u10_u4_n145 ) , .ZN( u1_u10_u4_n151 ) );
  NAND3_X1 u1_u10_u4_U99 (.A3( u1_u10_u4_n121 ) , .ZN( u1_u10_u4_n122 ) , .A2( u1_u10_u4_n144 ) , .A1( u1_u10_u4_n154 ) );
  AND3_X1 u1_u10_u7_U10 (.A3( u1_u10_u7_n110 ) , .A2( u1_u10_u7_n127 ) , .A1( u1_u10_u7_n132 ) , .ZN( u1_u10_u7_n92 ) );
  OAI21_X1 u1_u10_u7_U11 (.A( u1_u10_u7_n161 ) , .B1( u1_u10_u7_n168 ) , .B2( u1_u10_u7_n173 ) , .ZN( u1_u10_u7_n91 ) );
  AOI211_X1 u1_u10_u7_U12 (.A( u1_u10_u7_n117 ) , .ZN( u1_u10_u7_n118 ) , .C2( u1_u10_u7_n126 ) , .C1( u1_u10_u7_n177 ) , .B( u1_u10_u7_n180 ) );
  OAI22_X1 u1_u10_u7_U13 (.B1( u1_u10_u7_n115 ) , .ZN( u1_u10_u7_n117 ) , .A2( u1_u10_u7_n133 ) , .A1( u1_u10_u7_n137 ) , .B2( u1_u10_u7_n162 ) );
  INV_X1 u1_u10_u7_U14 (.A( u1_u10_u7_n116 ) , .ZN( u1_u10_u7_n180 ) );
  NOR3_X1 u1_u10_u7_U15 (.ZN( u1_u10_u7_n115 ) , .A3( u1_u10_u7_n145 ) , .A2( u1_u10_u7_n168 ) , .A1( u1_u10_u7_n169 ) );
  OAI211_X1 u1_u10_u7_U16 (.B( u1_u10_u7_n122 ) , .A( u1_u10_u7_n123 ) , .C2( u1_u10_u7_n124 ) , .ZN( u1_u10_u7_n154 ) , .C1( u1_u10_u7_n162 ) );
  AOI222_X1 u1_u10_u7_U17 (.ZN( u1_u10_u7_n122 ) , .C2( u1_u10_u7_n126 ) , .C1( u1_u10_u7_n145 ) , .B1( u1_u10_u7_n161 ) , .A2( u1_u10_u7_n165 ) , .B2( u1_u10_u7_n170 ) , .A1( u1_u10_u7_n176 ) );
  INV_X1 u1_u10_u7_U18 (.A( u1_u10_u7_n133 ) , .ZN( u1_u10_u7_n176 ) );
  NOR3_X1 u1_u10_u7_U19 (.A2( u1_u10_u7_n134 ) , .A1( u1_u10_u7_n135 ) , .ZN( u1_u10_u7_n136 ) , .A3( u1_u10_u7_n171 ) );
  NOR2_X1 u1_u10_u7_U20 (.A1( u1_u10_u7_n130 ) , .A2( u1_u10_u7_n134 ) , .ZN( u1_u10_u7_n153 ) );
  INV_X1 u1_u10_u7_U21 (.A( u1_u10_u7_n101 ) , .ZN( u1_u10_u7_n165 ) );
  NOR2_X1 u1_u10_u7_U22 (.ZN( u1_u10_u7_n111 ) , .A2( u1_u10_u7_n134 ) , .A1( u1_u10_u7_n169 ) );
  AOI21_X1 u1_u10_u7_U23 (.ZN( u1_u10_u7_n104 ) , .B2( u1_u10_u7_n112 ) , .B1( u1_u10_u7_n127 ) , .A( u1_u10_u7_n164 ) );
  AOI21_X1 u1_u10_u7_U24 (.ZN( u1_u10_u7_n106 ) , .B1( u1_u10_u7_n133 ) , .B2( u1_u10_u7_n146 ) , .A( u1_u10_u7_n162 ) );
  AOI21_X1 u1_u10_u7_U25 (.A( u1_u10_u7_n101 ) , .ZN( u1_u10_u7_n107 ) , .B2( u1_u10_u7_n128 ) , .B1( u1_u10_u7_n175 ) );
  INV_X1 u1_u10_u7_U26 (.A( u1_u10_u7_n138 ) , .ZN( u1_u10_u7_n171 ) );
  INV_X1 u1_u10_u7_U27 (.A( u1_u10_u7_n131 ) , .ZN( u1_u10_u7_n177 ) );
  INV_X1 u1_u10_u7_U28 (.A( u1_u10_u7_n110 ) , .ZN( u1_u10_u7_n174 ) );
  NAND2_X1 u1_u10_u7_U29 (.A1( u1_u10_u7_n129 ) , .A2( u1_u10_u7_n132 ) , .ZN( u1_u10_u7_n149 ) );
  OAI21_X1 u1_u10_u7_U3 (.ZN( u1_u10_u7_n159 ) , .A( u1_u10_u7_n165 ) , .B2( u1_u10_u7_n171 ) , .B1( u1_u10_u7_n174 ) );
  NAND2_X1 u1_u10_u7_U30 (.A1( u1_u10_u7_n113 ) , .A2( u1_u10_u7_n124 ) , .ZN( u1_u10_u7_n130 ) );
  INV_X1 u1_u10_u7_U31 (.A( u1_u10_u7_n112 ) , .ZN( u1_u10_u7_n173 ) );
  INV_X1 u1_u10_u7_U32 (.A( u1_u10_u7_n128 ) , .ZN( u1_u10_u7_n168 ) );
  INV_X1 u1_u10_u7_U33 (.A( u1_u10_u7_n148 ) , .ZN( u1_u10_u7_n169 ) );
  INV_X1 u1_u10_u7_U34 (.A( u1_u10_u7_n127 ) , .ZN( u1_u10_u7_n179 ) );
  NOR2_X1 u1_u10_u7_U35 (.ZN( u1_u10_u7_n101 ) , .A2( u1_u10_u7_n150 ) , .A1( u1_u10_u7_n156 ) );
  AOI211_X1 u1_u10_u7_U36 (.B( u1_u10_u7_n154 ) , .A( u1_u10_u7_n155 ) , .C1( u1_u10_u7_n156 ) , .ZN( u1_u10_u7_n157 ) , .C2( u1_u10_u7_n172 ) );
  INV_X1 u1_u10_u7_U37 (.A( u1_u10_u7_n153 ) , .ZN( u1_u10_u7_n172 ) );
  AOI211_X1 u1_u10_u7_U38 (.B( u1_u10_u7_n139 ) , .A( u1_u10_u7_n140 ) , .C2( u1_u10_u7_n141 ) , .ZN( u1_u10_u7_n142 ) , .C1( u1_u10_u7_n156 ) );
  NAND4_X1 u1_u10_u7_U39 (.A3( u1_u10_u7_n127 ) , .A2( u1_u10_u7_n128 ) , .A1( u1_u10_u7_n129 ) , .ZN( u1_u10_u7_n141 ) , .A4( u1_u10_u7_n147 ) );
  INV_X1 u1_u10_u7_U4 (.A( u1_u10_u7_n111 ) , .ZN( u1_u10_u7_n170 ) );
  AOI21_X1 u1_u10_u7_U40 (.A( u1_u10_u7_n137 ) , .B1( u1_u10_u7_n138 ) , .ZN( u1_u10_u7_n139 ) , .B2( u1_u10_u7_n146 ) );
  OAI22_X1 u1_u10_u7_U41 (.B1( u1_u10_u7_n136 ) , .ZN( u1_u10_u7_n140 ) , .A1( u1_u10_u7_n153 ) , .B2( u1_u10_u7_n162 ) , .A2( u1_u10_u7_n164 ) );
  AOI21_X1 u1_u10_u7_U42 (.ZN( u1_u10_u7_n123 ) , .B1( u1_u10_u7_n165 ) , .B2( u1_u10_u7_n177 ) , .A( u1_u10_u7_n97 ) );
  AOI21_X1 u1_u10_u7_U43 (.B2( u1_u10_u7_n113 ) , .B1( u1_u10_u7_n124 ) , .A( u1_u10_u7_n125 ) , .ZN( u1_u10_u7_n97 ) );
  INV_X1 u1_u10_u7_U44 (.A( u1_u10_u7_n125 ) , .ZN( u1_u10_u7_n161 ) );
  INV_X1 u1_u10_u7_U45 (.A( u1_u10_u7_n152 ) , .ZN( u1_u10_u7_n162 ) );
  AOI22_X1 u1_u10_u7_U46 (.A2( u1_u10_u7_n114 ) , .ZN( u1_u10_u7_n119 ) , .B1( u1_u10_u7_n130 ) , .A1( u1_u10_u7_n156 ) , .B2( u1_u10_u7_n165 ) );
  NAND2_X1 u1_u10_u7_U47 (.A2( u1_u10_u7_n112 ) , .ZN( u1_u10_u7_n114 ) , .A1( u1_u10_u7_n175 ) );
  AND2_X1 u1_u10_u7_U48 (.ZN( u1_u10_u7_n145 ) , .A2( u1_u10_u7_n98 ) , .A1( u1_u10_u7_n99 ) );
  NOR2_X1 u1_u10_u7_U49 (.ZN( u1_u10_u7_n137 ) , .A1( u1_u10_u7_n150 ) , .A2( u1_u10_u7_n161 ) );
  INV_X1 u1_u10_u7_U5 (.A( u1_u10_u7_n149 ) , .ZN( u1_u10_u7_n175 ) );
  AOI21_X1 u1_u10_u7_U50 (.ZN( u1_u10_u7_n105 ) , .B2( u1_u10_u7_n110 ) , .A( u1_u10_u7_n125 ) , .B1( u1_u10_u7_n147 ) );
  NAND2_X1 u1_u10_u7_U51 (.ZN( u1_u10_u7_n146 ) , .A1( u1_u10_u7_n95 ) , .A2( u1_u10_u7_n98 ) );
  NAND2_X1 u1_u10_u7_U52 (.A2( u1_u10_u7_n103 ) , .ZN( u1_u10_u7_n147 ) , .A1( u1_u10_u7_n93 ) );
  NAND2_X1 u1_u10_u7_U53 (.A1( u1_u10_u7_n103 ) , .ZN( u1_u10_u7_n127 ) , .A2( u1_u10_u7_n99 ) );
  OR2_X1 u1_u10_u7_U54 (.ZN( u1_u10_u7_n126 ) , .A2( u1_u10_u7_n152 ) , .A1( u1_u10_u7_n156 ) );
  NAND2_X1 u1_u10_u7_U55 (.A2( u1_u10_u7_n102 ) , .A1( u1_u10_u7_n103 ) , .ZN( u1_u10_u7_n133 ) );
  NAND2_X1 u1_u10_u7_U56 (.ZN( u1_u10_u7_n112 ) , .A2( u1_u10_u7_n96 ) , .A1( u1_u10_u7_n99 ) );
  NAND2_X1 u1_u10_u7_U57 (.A2( u1_u10_u7_n102 ) , .ZN( u1_u10_u7_n128 ) , .A1( u1_u10_u7_n98 ) );
  NAND2_X1 u1_u10_u7_U58 (.A1( u1_u10_u7_n100 ) , .ZN( u1_u10_u7_n113 ) , .A2( u1_u10_u7_n93 ) );
  NAND2_X1 u1_u10_u7_U59 (.A2( u1_u10_u7_n102 ) , .ZN( u1_u10_u7_n124 ) , .A1( u1_u10_u7_n96 ) );
  INV_X1 u1_u10_u7_U6 (.A( u1_u10_u7_n154 ) , .ZN( u1_u10_u7_n178 ) );
  NAND2_X1 u1_u10_u7_U60 (.ZN( u1_u10_u7_n110 ) , .A1( u1_u10_u7_n95 ) , .A2( u1_u10_u7_n96 ) );
  INV_X1 u1_u10_u7_U61 (.A( u1_u10_u7_n150 ) , .ZN( u1_u10_u7_n164 ) );
  AND2_X1 u1_u10_u7_U62 (.ZN( u1_u10_u7_n134 ) , .A1( u1_u10_u7_n93 ) , .A2( u1_u10_u7_n98 ) );
  NAND2_X1 u1_u10_u7_U63 (.A1( u1_u10_u7_n100 ) , .A2( u1_u10_u7_n102 ) , .ZN( u1_u10_u7_n129 ) );
  NAND2_X1 u1_u10_u7_U64 (.A2( u1_u10_u7_n103 ) , .ZN( u1_u10_u7_n131 ) , .A1( u1_u10_u7_n95 ) );
  NAND2_X1 u1_u10_u7_U65 (.A1( u1_u10_u7_n100 ) , .ZN( u1_u10_u7_n138 ) , .A2( u1_u10_u7_n99 ) );
  NAND2_X1 u1_u10_u7_U66 (.ZN( u1_u10_u7_n132 ) , .A1( u1_u10_u7_n93 ) , .A2( u1_u10_u7_n96 ) );
  NAND2_X1 u1_u10_u7_U67 (.A1( u1_u10_u7_n100 ) , .ZN( u1_u10_u7_n148 ) , .A2( u1_u10_u7_n95 ) );
  NOR2_X1 u1_u10_u7_U68 (.A2( u1_u10_X_47 ) , .ZN( u1_u10_u7_n150 ) , .A1( u1_u10_u7_n163 ) );
  NOR2_X1 u1_u10_u7_U69 (.A2( u1_u10_X_43 ) , .A1( u1_u10_X_44 ) , .ZN( u1_u10_u7_n103 ) );
  AOI211_X1 u1_u10_u7_U7 (.ZN( u1_u10_u7_n116 ) , .A( u1_u10_u7_n155 ) , .C1( u1_u10_u7_n161 ) , .C2( u1_u10_u7_n171 ) , .B( u1_u10_u7_n94 ) );
  NOR2_X1 u1_u10_u7_U70 (.A2( u1_u10_X_48 ) , .A1( u1_u10_u7_n166 ) , .ZN( u1_u10_u7_n95 ) );
  NOR2_X1 u1_u10_u7_U71 (.A2( u1_u10_X_45 ) , .A1( u1_u10_X_48 ) , .ZN( u1_u10_u7_n99 ) );
  NOR2_X1 u1_u10_u7_U72 (.A2( u1_u10_X_44 ) , .A1( u1_u10_u7_n167 ) , .ZN( u1_u10_u7_n98 ) );
  NOR2_X1 u1_u10_u7_U73 (.A2( u1_u10_X_46 ) , .A1( u1_u10_X_47 ) , .ZN( u1_u10_u7_n152 ) );
  AND2_X1 u1_u10_u7_U74 (.A1( u1_u10_X_47 ) , .ZN( u1_u10_u7_n156 ) , .A2( u1_u10_u7_n163 ) );
  NAND2_X1 u1_u10_u7_U75 (.A2( u1_u10_X_46 ) , .A1( u1_u10_X_47 ) , .ZN( u1_u10_u7_n125 ) );
  AND2_X1 u1_u10_u7_U76 (.A2( u1_u10_X_45 ) , .A1( u1_u10_X_48 ) , .ZN( u1_u10_u7_n102 ) );
  AND2_X1 u1_u10_u7_U77 (.A2( u1_u10_X_43 ) , .A1( u1_u10_X_44 ) , .ZN( u1_u10_u7_n96 ) );
  AND2_X1 u1_u10_u7_U78 (.A1( u1_u10_X_44 ) , .ZN( u1_u10_u7_n100 ) , .A2( u1_u10_u7_n167 ) );
  AND2_X1 u1_u10_u7_U79 (.A1( u1_u10_X_48 ) , .A2( u1_u10_u7_n166 ) , .ZN( u1_u10_u7_n93 ) );
  OAI222_X1 u1_u10_u7_U8 (.C2( u1_u10_u7_n101 ) , .B2( u1_u10_u7_n111 ) , .A1( u1_u10_u7_n113 ) , .C1( u1_u10_u7_n146 ) , .A2( u1_u10_u7_n162 ) , .B1( u1_u10_u7_n164 ) , .ZN( u1_u10_u7_n94 ) );
  INV_X1 u1_u10_u7_U80 (.A( u1_u10_X_46 ) , .ZN( u1_u10_u7_n163 ) );
  INV_X1 u1_u10_u7_U81 (.A( u1_u10_X_43 ) , .ZN( u1_u10_u7_n167 ) );
  INV_X1 u1_u10_u7_U82 (.A( u1_u10_X_45 ) , .ZN( u1_u10_u7_n166 ) );
  NAND4_X1 u1_u10_u7_U83 (.ZN( u1_out10_27 ) , .A4( u1_u10_u7_n118 ) , .A3( u1_u10_u7_n119 ) , .A2( u1_u10_u7_n120 ) , .A1( u1_u10_u7_n121 ) );
  OAI21_X1 u1_u10_u7_U84 (.ZN( u1_u10_u7_n121 ) , .B2( u1_u10_u7_n145 ) , .A( u1_u10_u7_n150 ) , .B1( u1_u10_u7_n174 ) );
  OAI21_X1 u1_u10_u7_U85 (.ZN( u1_u10_u7_n120 ) , .A( u1_u10_u7_n161 ) , .B2( u1_u10_u7_n170 ) , .B1( u1_u10_u7_n179 ) );
  NAND4_X1 u1_u10_u7_U86 (.ZN( u1_out10_21 ) , .A4( u1_u10_u7_n157 ) , .A3( u1_u10_u7_n158 ) , .A2( u1_u10_u7_n159 ) , .A1( u1_u10_u7_n160 ) );
  OAI21_X1 u1_u10_u7_U87 (.B1( u1_u10_u7_n145 ) , .ZN( u1_u10_u7_n160 ) , .A( u1_u10_u7_n161 ) , .B2( u1_u10_u7_n177 ) );
  AOI22_X1 u1_u10_u7_U88 (.B2( u1_u10_u7_n149 ) , .B1( u1_u10_u7_n150 ) , .A2( u1_u10_u7_n151 ) , .A1( u1_u10_u7_n152 ) , .ZN( u1_u10_u7_n158 ) );
  NAND4_X1 u1_u10_u7_U89 (.ZN( u1_out10_15 ) , .A4( u1_u10_u7_n142 ) , .A3( u1_u10_u7_n143 ) , .A2( u1_u10_u7_n144 ) , .A1( u1_u10_u7_n178 ) );
  OAI221_X1 u1_u10_u7_U9 (.C1( u1_u10_u7_n101 ) , .C2( u1_u10_u7_n147 ) , .ZN( u1_u10_u7_n155 ) , .B2( u1_u10_u7_n162 ) , .A( u1_u10_u7_n91 ) , .B1( u1_u10_u7_n92 ) );
  OR2_X1 u1_u10_u7_U90 (.A2( u1_u10_u7_n125 ) , .A1( u1_u10_u7_n129 ) , .ZN( u1_u10_u7_n144 ) );
  AOI22_X1 u1_u10_u7_U91 (.A2( u1_u10_u7_n126 ) , .ZN( u1_u10_u7_n143 ) , .B2( u1_u10_u7_n165 ) , .B1( u1_u10_u7_n173 ) , .A1( u1_u10_u7_n174 ) );
  NAND4_X1 u1_u10_u7_U92 (.ZN( u1_out10_5 ) , .A4( u1_u10_u7_n108 ) , .A3( u1_u10_u7_n109 ) , .A1( u1_u10_u7_n116 ) , .A2( u1_u10_u7_n123 ) );
  AOI22_X1 u1_u10_u7_U93 (.ZN( u1_u10_u7_n109 ) , .A2( u1_u10_u7_n126 ) , .B2( u1_u10_u7_n145 ) , .B1( u1_u10_u7_n156 ) , .A1( u1_u10_u7_n171 ) );
  NOR4_X1 u1_u10_u7_U94 (.A4( u1_u10_u7_n104 ) , .A3( u1_u10_u7_n105 ) , .A2( u1_u10_u7_n106 ) , .A1( u1_u10_u7_n107 ) , .ZN( u1_u10_u7_n108 ) );
  NAND3_X1 u1_u10_u7_U95 (.A3( u1_u10_u7_n146 ) , .A2( u1_u10_u7_n147 ) , .A1( u1_u10_u7_n148 ) , .ZN( u1_u10_u7_n151 ) );
  NAND3_X1 u1_u10_u7_U96 (.A3( u1_u10_u7_n131 ) , .A2( u1_u10_u7_n132 ) , .A1( u1_u10_u7_n133 ) , .ZN( u1_u10_u7_n135 ) );
  XOR2_X1 u1_u11_U1 (.B( u1_K12_9 ) , .A( u1_R10_6 ) , .Z( u1_u11_X_9 ) );
  XOR2_X1 u1_u11_U2 (.B( u1_K12_8 ) , .A( u1_R10_5 ) , .Z( u1_u11_X_8 ) );
  XOR2_X1 u1_u11_U3 (.B( u1_K12_7 ) , .A( u1_R10_4 ) , .Z( u1_u11_X_7 ) );
  XOR2_X1 u1_u11_U46 (.B( u1_K12_12 ) , .A( u1_R10_9 ) , .Z( u1_u11_X_12 ) );
  XOR2_X1 u1_u11_U47 (.B( u1_K12_11 ) , .A( u1_R10_8 ) , .Z( u1_u11_X_11 ) );
  XOR2_X1 u1_u11_U48 (.B( u1_K12_10 ) , .A( u1_R10_7 ) , .Z( u1_u11_X_10 ) );
  NOR2_X1 u1_u11_u1_U10 (.A1( u1_u11_u1_n112 ) , .A2( u1_u11_u1_n116 ) , .ZN( u1_u11_u1_n118 ) );
  NAND3_X1 u1_u11_u1_U100 (.ZN( u1_u11_u1_n113 ) , .A1( u1_u11_u1_n120 ) , .A3( u1_u11_u1_n133 ) , .A2( u1_u11_u1_n155 ) );
  OAI21_X1 u1_u11_u1_U11 (.ZN( u1_u11_u1_n101 ) , .B1( u1_u11_u1_n141 ) , .A( u1_u11_u1_n146 ) , .B2( u1_u11_u1_n183 ) );
  AOI21_X1 u1_u11_u1_U12 (.B2( u1_u11_u1_n155 ) , .B1( u1_u11_u1_n156 ) , .ZN( u1_u11_u1_n157 ) , .A( u1_u11_u1_n174 ) );
  NAND2_X1 u1_u11_u1_U13 (.ZN( u1_u11_u1_n140 ) , .A2( u1_u11_u1_n150 ) , .A1( u1_u11_u1_n155 ) );
  NAND2_X1 u1_u11_u1_U14 (.A1( u1_u11_u1_n131 ) , .ZN( u1_u11_u1_n147 ) , .A2( u1_u11_u1_n153 ) );
  INV_X1 u1_u11_u1_U15 (.A( u1_u11_u1_n139 ) , .ZN( u1_u11_u1_n174 ) );
  OR4_X1 u1_u11_u1_U16 (.A4( u1_u11_u1_n106 ) , .A3( u1_u11_u1_n107 ) , .ZN( u1_u11_u1_n108 ) , .A1( u1_u11_u1_n117 ) , .A2( u1_u11_u1_n184 ) );
  AOI21_X1 u1_u11_u1_U17 (.ZN( u1_u11_u1_n106 ) , .A( u1_u11_u1_n112 ) , .B1( u1_u11_u1_n154 ) , .B2( u1_u11_u1_n156 ) );
  AOI21_X1 u1_u11_u1_U18 (.ZN( u1_u11_u1_n107 ) , .B1( u1_u11_u1_n134 ) , .B2( u1_u11_u1_n149 ) , .A( u1_u11_u1_n174 ) );
  INV_X1 u1_u11_u1_U19 (.A( u1_u11_u1_n101 ) , .ZN( u1_u11_u1_n184 ) );
  INV_X1 u1_u11_u1_U20 (.A( u1_u11_u1_n112 ) , .ZN( u1_u11_u1_n171 ) );
  NAND2_X1 u1_u11_u1_U21 (.ZN( u1_u11_u1_n141 ) , .A1( u1_u11_u1_n153 ) , .A2( u1_u11_u1_n156 ) );
  AND2_X1 u1_u11_u1_U22 (.A1( u1_u11_u1_n123 ) , .ZN( u1_u11_u1_n134 ) , .A2( u1_u11_u1_n161 ) );
  NAND2_X1 u1_u11_u1_U23 (.A2( u1_u11_u1_n115 ) , .A1( u1_u11_u1_n116 ) , .ZN( u1_u11_u1_n148 ) );
  NAND2_X1 u1_u11_u1_U24 (.A2( u1_u11_u1_n133 ) , .A1( u1_u11_u1_n135 ) , .ZN( u1_u11_u1_n159 ) );
  NAND2_X1 u1_u11_u1_U25 (.A2( u1_u11_u1_n115 ) , .A1( u1_u11_u1_n120 ) , .ZN( u1_u11_u1_n132 ) );
  INV_X1 u1_u11_u1_U26 (.A( u1_u11_u1_n154 ) , .ZN( u1_u11_u1_n178 ) );
  INV_X1 u1_u11_u1_U27 (.A( u1_u11_u1_n151 ) , .ZN( u1_u11_u1_n183 ) );
  AND2_X1 u1_u11_u1_U28 (.A1( u1_u11_u1_n129 ) , .A2( u1_u11_u1_n133 ) , .ZN( u1_u11_u1_n149 ) );
  INV_X1 u1_u11_u1_U29 (.A( u1_u11_u1_n131 ) , .ZN( u1_u11_u1_n180 ) );
  INV_X1 u1_u11_u1_U3 (.A( u1_u11_u1_n159 ) , .ZN( u1_u11_u1_n182 ) );
  OAI221_X1 u1_u11_u1_U30 (.A( u1_u11_u1_n119 ) , .C2( u1_u11_u1_n129 ) , .ZN( u1_u11_u1_n138 ) , .B2( u1_u11_u1_n152 ) , .C1( u1_u11_u1_n174 ) , .B1( u1_u11_u1_n187 ) );
  INV_X1 u1_u11_u1_U31 (.A( u1_u11_u1_n148 ) , .ZN( u1_u11_u1_n187 ) );
  AOI211_X1 u1_u11_u1_U32 (.B( u1_u11_u1_n117 ) , .A( u1_u11_u1_n118 ) , .ZN( u1_u11_u1_n119 ) , .C2( u1_u11_u1_n146 ) , .C1( u1_u11_u1_n159 ) );
  NOR2_X1 u1_u11_u1_U33 (.A1( u1_u11_u1_n168 ) , .A2( u1_u11_u1_n176 ) , .ZN( u1_u11_u1_n98 ) );
  AOI211_X1 u1_u11_u1_U34 (.B( u1_u11_u1_n162 ) , .A( u1_u11_u1_n163 ) , .C2( u1_u11_u1_n164 ) , .ZN( u1_u11_u1_n165 ) , .C1( u1_u11_u1_n171 ) );
  AOI21_X1 u1_u11_u1_U35 (.A( u1_u11_u1_n160 ) , .B2( u1_u11_u1_n161 ) , .ZN( u1_u11_u1_n162 ) , .B1( u1_u11_u1_n182 ) );
  OR2_X1 u1_u11_u1_U36 (.A2( u1_u11_u1_n157 ) , .A1( u1_u11_u1_n158 ) , .ZN( u1_u11_u1_n163 ) );
  NAND2_X1 u1_u11_u1_U37 (.A1( u1_u11_u1_n128 ) , .ZN( u1_u11_u1_n146 ) , .A2( u1_u11_u1_n160 ) );
  NAND2_X1 u1_u11_u1_U38 (.A2( u1_u11_u1_n112 ) , .ZN( u1_u11_u1_n139 ) , .A1( u1_u11_u1_n152 ) );
  NAND2_X1 u1_u11_u1_U39 (.A1( u1_u11_u1_n105 ) , .ZN( u1_u11_u1_n156 ) , .A2( u1_u11_u1_n99 ) );
  AOI221_X1 u1_u11_u1_U4 (.A( u1_u11_u1_n138 ) , .C2( u1_u11_u1_n139 ) , .C1( u1_u11_u1_n140 ) , .B2( u1_u11_u1_n141 ) , .ZN( u1_u11_u1_n142 ) , .B1( u1_u11_u1_n175 ) );
  AOI221_X1 u1_u11_u1_U40 (.B1( u1_u11_u1_n140 ) , .ZN( u1_u11_u1_n167 ) , .B2( u1_u11_u1_n172 ) , .C2( u1_u11_u1_n175 ) , .C1( u1_u11_u1_n178 ) , .A( u1_u11_u1_n188 ) );
  INV_X1 u1_u11_u1_U41 (.ZN( u1_u11_u1_n188 ) , .A( u1_u11_u1_n97 ) );
  AOI211_X1 u1_u11_u1_U42 (.A( u1_u11_u1_n118 ) , .C1( u1_u11_u1_n132 ) , .C2( u1_u11_u1_n139 ) , .B( u1_u11_u1_n96 ) , .ZN( u1_u11_u1_n97 ) );
  AOI21_X1 u1_u11_u1_U43 (.B2( u1_u11_u1_n121 ) , .B1( u1_u11_u1_n135 ) , .A( u1_u11_u1_n152 ) , .ZN( u1_u11_u1_n96 ) );
  NOR2_X1 u1_u11_u1_U44 (.ZN( u1_u11_u1_n117 ) , .A1( u1_u11_u1_n121 ) , .A2( u1_u11_u1_n160 ) );
  OAI21_X1 u1_u11_u1_U45 (.B2( u1_u11_u1_n123 ) , .ZN( u1_u11_u1_n145 ) , .B1( u1_u11_u1_n160 ) , .A( u1_u11_u1_n185 ) );
  INV_X1 u1_u11_u1_U46 (.A( u1_u11_u1_n122 ) , .ZN( u1_u11_u1_n185 ) );
  AOI21_X1 u1_u11_u1_U47 (.B2( u1_u11_u1_n120 ) , .B1( u1_u11_u1_n121 ) , .ZN( u1_u11_u1_n122 ) , .A( u1_u11_u1_n128 ) );
  AOI21_X1 u1_u11_u1_U48 (.A( u1_u11_u1_n128 ) , .B2( u1_u11_u1_n129 ) , .ZN( u1_u11_u1_n130 ) , .B1( u1_u11_u1_n150 ) );
  NAND2_X1 u1_u11_u1_U49 (.ZN( u1_u11_u1_n112 ) , .A1( u1_u11_u1_n169 ) , .A2( u1_u11_u1_n170 ) );
  AOI211_X1 u1_u11_u1_U5 (.ZN( u1_u11_u1_n124 ) , .A( u1_u11_u1_n138 ) , .C2( u1_u11_u1_n139 ) , .B( u1_u11_u1_n145 ) , .C1( u1_u11_u1_n147 ) );
  NAND2_X1 u1_u11_u1_U50 (.ZN( u1_u11_u1_n129 ) , .A2( u1_u11_u1_n95 ) , .A1( u1_u11_u1_n98 ) );
  NAND2_X1 u1_u11_u1_U51 (.A1( u1_u11_u1_n102 ) , .ZN( u1_u11_u1_n154 ) , .A2( u1_u11_u1_n99 ) );
  NAND2_X1 u1_u11_u1_U52 (.A2( u1_u11_u1_n100 ) , .ZN( u1_u11_u1_n135 ) , .A1( u1_u11_u1_n99 ) );
  AOI21_X1 u1_u11_u1_U53 (.A( u1_u11_u1_n152 ) , .B2( u1_u11_u1_n153 ) , .B1( u1_u11_u1_n154 ) , .ZN( u1_u11_u1_n158 ) );
  INV_X1 u1_u11_u1_U54 (.A( u1_u11_u1_n160 ) , .ZN( u1_u11_u1_n175 ) );
  NAND2_X1 u1_u11_u1_U55 (.A1( u1_u11_u1_n100 ) , .ZN( u1_u11_u1_n116 ) , .A2( u1_u11_u1_n95 ) );
  NAND2_X1 u1_u11_u1_U56 (.A1( u1_u11_u1_n102 ) , .ZN( u1_u11_u1_n131 ) , .A2( u1_u11_u1_n95 ) );
  NAND2_X1 u1_u11_u1_U57 (.A2( u1_u11_u1_n104 ) , .ZN( u1_u11_u1_n121 ) , .A1( u1_u11_u1_n98 ) );
  NAND2_X1 u1_u11_u1_U58 (.A1( u1_u11_u1_n103 ) , .ZN( u1_u11_u1_n153 ) , .A2( u1_u11_u1_n98 ) );
  NAND2_X1 u1_u11_u1_U59 (.A2( u1_u11_u1_n104 ) , .A1( u1_u11_u1_n105 ) , .ZN( u1_u11_u1_n133 ) );
  AOI22_X1 u1_u11_u1_U6 (.B2( u1_u11_u1_n113 ) , .A2( u1_u11_u1_n114 ) , .ZN( u1_u11_u1_n125 ) , .A1( u1_u11_u1_n171 ) , .B1( u1_u11_u1_n173 ) );
  NAND2_X1 u1_u11_u1_U60 (.ZN( u1_u11_u1_n150 ) , .A2( u1_u11_u1_n98 ) , .A1( u1_u11_u1_n99 ) );
  NAND2_X1 u1_u11_u1_U61 (.A1( u1_u11_u1_n105 ) , .ZN( u1_u11_u1_n155 ) , .A2( u1_u11_u1_n95 ) );
  OAI21_X1 u1_u11_u1_U62 (.ZN( u1_u11_u1_n109 ) , .B1( u1_u11_u1_n129 ) , .B2( u1_u11_u1_n160 ) , .A( u1_u11_u1_n167 ) );
  NAND2_X1 u1_u11_u1_U63 (.A2( u1_u11_u1_n100 ) , .A1( u1_u11_u1_n103 ) , .ZN( u1_u11_u1_n120 ) );
  NAND2_X1 u1_u11_u1_U64 (.A1( u1_u11_u1_n102 ) , .A2( u1_u11_u1_n104 ) , .ZN( u1_u11_u1_n115 ) );
  NAND2_X1 u1_u11_u1_U65 (.A2( u1_u11_u1_n100 ) , .A1( u1_u11_u1_n104 ) , .ZN( u1_u11_u1_n151 ) );
  NAND2_X1 u1_u11_u1_U66 (.A2( u1_u11_u1_n103 ) , .A1( u1_u11_u1_n105 ) , .ZN( u1_u11_u1_n161 ) );
  INV_X1 u1_u11_u1_U67 (.A( u1_u11_u1_n152 ) , .ZN( u1_u11_u1_n173 ) );
  INV_X1 u1_u11_u1_U68 (.A( u1_u11_u1_n128 ) , .ZN( u1_u11_u1_n172 ) );
  NAND2_X1 u1_u11_u1_U69 (.A2( u1_u11_u1_n102 ) , .A1( u1_u11_u1_n103 ) , .ZN( u1_u11_u1_n123 ) );
  NAND2_X1 u1_u11_u1_U7 (.ZN( u1_u11_u1_n114 ) , .A1( u1_u11_u1_n134 ) , .A2( u1_u11_u1_n156 ) );
  NOR2_X1 u1_u11_u1_U70 (.A2( u1_u11_X_7 ) , .A1( u1_u11_X_8 ) , .ZN( u1_u11_u1_n95 ) );
  NOR2_X1 u1_u11_u1_U71 (.A1( u1_u11_X_12 ) , .A2( u1_u11_X_9 ) , .ZN( u1_u11_u1_n100 ) );
  NOR2_X1 u1_u11_u1_U72 (.A2( u1_u11_X_8 ) , .A1( u1_u11_u1_n177 ) , .ZN( u1_u11_u1_n99 ) );
  NOR2_X1 u1_u11_u1_U73 (.A2( u1_u11_X_12 ) , .ZN( u1_u11_u1_n102 ) , .A1( u1_u11_u1_n176 ) );
  NOR2_X1 u1_u11_u1_U74 (.A2( u1_u11_X_9 ) , .ZN( u1_u11_u1_n105 ) , .A1( u1_u11_u1_n168 ) );
  NAND2_X1 u1_u11_u1_U75 (.A1( u1_u11_X_10 ) , .ZN( u1_u11_u1_n160 ) , .A2( u1_u11_u1_n169 ) );
  NAND2_X1 u1_u11_u1_U76 (.A2( u1_u11_X_10 ) , .A1( u1_u11_X_11 ) , .ZN( u1_u11_u1_n152 ) );
  NAND2_X1 u1_u11_u1_U77 (.A1( u1_u11_X_11 ) , .ZN( u1_u11_u1_n128 ) , .A2( u1_u11_u1_n170 ) );
  AND2_X1 u1_u11_u1_U78 (.A2( u1_u11_X_7 ) , .A1( u1_u11_X_8 ) , .ZN( u1_u11_u1_n104 ) );
  AND2_X1 u1_u11_u1_U79 (.A1( u1_u11_X_8 ) , .ZN( u1_u11_u1_n103 ) , .A2( u1_u11_u1_n177 ) );
  AOI22_X1 u1_u11_u1_U8 (.B2( u1_u11_u1_n136 ) , .A2( u1_u11_u1_n137 ) , .ZN( u1_u11_u1_n143 ) , .A1( u1_u11_u1_n171 ) , .B1( u1_u11_u1_n173 ) );
  INV_X1 u1_u11_u1_U80 (.A( u1_u11_X_10 ) , .ZN( u1_u11_u1_n170 ) );
  INV_X1 u1_u11_u1_U81 (.A( u1_u11_X_9 ) , .ZN( u1_u11_u1_n176 ) );
  INV_X1 u1_u11_u1_U82 (.A( u1_u11_X_11 ) , .ZN( u1_u11_u1_n169 ) );
  INV_X1 u1_u11_u1_U83 (.A( u1_u11_X_12 ) , .ZN( u1_u11_u1_n168 ) );
  INV_X1 u1_u11_u1_U84 (.A( u1_u11_X_7 ) , .ZN( u1_u11_u1_n177 ) );
  NAND4_X1 u1_u11_u1_U85 (.ZN( u1_out11_18 ) , .A4( u1_u11_u1_n165 ) , .A3( u1_u11_u1_n166 ) , .A1( u1_u11_u1_n167 ) , .A2( u1_u11_u1_n186 ) );
  AOI22_X1 u1_u11_u1_U86 (.B2( u1_u11_u1_n146 ) , .B1( u1_u11_u1_n147 ) , .A2( u1_u11_u1_n148 ) , .ZN( u1_u11_u1_n166 ) , .A1( u1_u11_u1_n172 ) );
  INV_X1 u1_u11_u1_U87 (.A( u1_u11_u1_n145 ) , .ZN( u1_u11_u1_n186 ) );
  NAND4_X1 u1_u11_u1_U88 (.ZN( u1_out11_2 ) , .A4( u1_u11_u1_n142 ) , .A3( u1_u11_u1_n143 ) , .A2( u1_u11_u1_n144 ) , .A1( u1_u11_u1_n179 ) );
  OAI21_X1 u1_u11_u1_U89 (.B2( u1_u11_u1_n132 ) , .ZN( u1_u11_u1_n144 ) , .A( u1_u11_u1_n146 ) , .B1( u1_u11_u1_n180 ) );
  INV_X1 u1_u11_u1_U9 (.A( u1_u11_u1_n147 ) , .ZN( u1_u11_u1_n181 ) );
  INV_X1 u1_u11_u1_U90 (.A( u1_u11_u1_n130 ) , .ZN( u1_u11_u1_n179 ) );
  NAND4_X1 u1_u11_u1_U91 (.ZN( u1_out11_28 ) , .A4( u1_u11_u1_n124 ) , .A3( u1_u11_u1_n125 ) , .A2( u1_u11_u1_n126 ) , .A1( u1_u11_u1_n127 ) );
  OAI21_X1 u1_u11_u1_U92 (.ZN( u1_u11_u1_n127 ) , .B2( u1_u11_u1_n139 ) , .B1( u1_u11_u1_n175 ) , .A( u1_u11_u1_n183 ) );
  OAI21_X1 u1_u11_u1_U93 (.ZN( u1_u11_u1_n126 ) , .B2( u1_u11_u1_n140 ) , .A( u1_u11_u1_n146 ) , .B1( u1_u11_u1_n178 ) );
  OR4_X1 u1_u11_u1_U94 (.ZN( u1_out11_13 ) , .A4( u1_u11_u1_n108 ) , .A3( u1_u11_u1_n109 ) , .A2( u1_u11_u1_n110 ) , .A1( u1_u11_u1_n111 ) );
  AOI21_X1 u1_u11_u1_U95 (.ZN( u1_u11_u1_n111 ) , .A( u1_u11_u1_n128 ) , .B2( u1_u11_u1_n131 ) , .B1( u1_u11_u1_n135 ) );
  AOI21_X1 u1_u11_u1_U96 (.ZN( u1_u11_u1_n110 ) , .A( u1_u11_u1_n116 ) , .B1( u1_u11_u1_n152 ) , .B2( u1_u11_u1_n160 ) );
  NAND3_X1 u1_u11_u1_U97 (.A3( u1_u11_u1_n149 ) , .A2( u1_u11_u1_n150 ) , .A1( u1_u11_u1_n151 ) , .ZN( u1_u11_u1_n164 ) );
  NAND3_X1 u1_u11_u1_U98 (.A3( u1_u11_u1_n134 ) , .A2( u1_u11_u1_n135 ) , .ZN( u1_u11_u1_n136 ) , .A1( u1_u11_u1_n151 ) );
  NAND3_X1 u1_u11_u1_U99 (.A1( u1_u11_u1_n133 ) , .ZN( u1_u11_u1_n137 ) , .A2( u1_u11_u1_n154 ) , .A3( u1_u11_u1_n181 ) );
  XOR2_X1 u1_u12_U20 (.B( u1_K13_36 ) , .A( u1_R11_25 ) , .Z( u1_u12_X_36 ) );
  XOR2_X1 u1_u12_U21 (.B( u1_K13_35 ) , .A( u1_R11_24 ) , .Z( u1_u12_X_35 ) );
  XOR2_X1 u1_u12_U22 (.B( u1_K13_34 ) , .A( u1_R11_23 ) , .Z( u1_u12_X_34 ) );
  XOR2_X1 u1_u12_U23 (.B( u1_K13_33 ) , .A( u1_R11_22 ) , .Z( u1_u12_X_33 ) );
  XOR2_X1 u1_u12_U24 (.B( u1_K13_32 ) , .A( u1_R11_21 ) , .Z( u1_u12_X_32 ) );
  XOR2_X1 u1_u12_U25 (.B( u1_K13_31 ) , .A( u1_R11_20 ) , .Z( u1_u12_X_31 ) );
  XOR2_X1 u1_u12_U26 (.B( u1_K13_30 ) , .A( u1_R11_21 ) , .Z( u1_u12_X_30 ) );
  XOR2_X1 u1_u12_U28 (.B( u1_K13_29 ) , .A( u1_R11_20 ) , .Z( u1_u12_X_29 ) );
  XOR2_X1 u1_u12_U29 (.B( u1_K13_28 ) , .A( u1_R11_19 ) , .Z( u1_u12_X_28 ) );
  XOR2_X1 u1_u12_U30 (.B( u1_K13_27 ) , .A( u1_R11_18 ) , .Z( u1_u12_X_27 ) );
  XOR2_X1 u1_u12_U31 (.B( u1_K13_26 ) , .A( u1_R11_17 ) , .Z( u1_u12_X_26 ) );
  XOR2_X1 u1_u12_U32 (.B( u1_K13_25 ) , .A( u1_R11_16 ) , .Z( u1_u12_X_25 ) );
  OAI22_X1 u1_u12_u4_U10 (.B2( u1_u12_u4_n135 ) , .ZN( u1_u12_u4_n137 ) , .B1( u1_u12_u4_n153 ) , .A1( u1_u12_u4_n155 ) , .A2( u1_u12_u4_n171 ) );
  AND3_X1 u1_u12_u4_U11 (.A2( u1_u12_u4_n134 ) , .ZN( u1_u12_u4_n135 ) , .A3( u1_u12_u4_n145 ) , .A1( u1_u12_u4_n157 ) );
  NAND2_X1 u1_u12_u4_U12 (.ZN( u1_u12_u4_n132 ) , .A2( u1_u12_u4_n170 ) , .A1( u1_u12_u4_n173 ) );
  AOI21_X1 u1_u12_u4_U13 (.B2( u1_u12_u4_n160 ) , .B1( u1_u12_u4_n161 ) , .ZN( u1_u12_u4_n162 ) , .A( u1_u12_u4_n170 ) );
  AOI21_X1 u1_u12_u4_U14 (.ZN( u1_u12_u4_n107 ) , .B2( u1_u12_u4_n143 ) , .A( u1_u12_u4_n174 ) , .B1( u1_u12_u4_n184 ) );
  AOI21_X1 u1_u12_u4_U15 (.B2( u1_u12_u4_n158 ) , .B1( u1_u12_u4_n159 ) , .ZN( u1_u12_u4_n163 ) , .A( u1_u12_u4_n174 ) );
  AOI21_X1 u1_u12_u4_U16 (.A( u1_u12_u4_n153 ) , .B2( u1_u12_u4_n154 ) , .B1( u1_u12_u4_n155 ) , .ZN( u1_u12_u4_n165 ) );
  AOI21_X1 u1_u12_u4_U17 (.A( u1_u12_u4_n156 ) , .B2( u1_u12_u4_n157 ) , .ZN( u1_u12_u4_n164 ) , .B1( u1_u12_u4_n184 ) );
  INV_X1 u1_u12_u4_U18 (.A( u1_u12_u4_n138 ) , .ZN( u1_u12_u4_n170 ) );
  AND2_X1 u1_u12_u4_U19 (.A2( u1_u12_u4_n120 ) , .ZN( u1_u12_u4_n155 ) , .A1( u1_u12_u4_n160 ) );
  INV_X1 u1_u12_u4_U20 (.A( u1_u12_u4_n156 ) , .ZN( u1_u12_u4_n175 ) );
  NAND2_X1 u1_u12_u4_U21 (.A2( u1_u12_u4_n118 ) , .ZN( u1_u12_u4_n131 ) , .A1( u1_u12_u4_n147 ) );
  NAND2_X1 u1_u12_u4_U22 (.A1( u1_u12_u4_n119 ) , .A2( u1_u12_u4_n120 ) , .ZN( u1_u12_u4_n130 ) );
  NAND2_X1 u1_u12_u4_U23 (.ZN( u1_u12_u4_n117 ) , .A2( u1_u12_u4_n118 ) , .A1( u1_u12_u4_n148 ) );
  NAND2_X1 u1_u12_u4_U24 (.ZN( u1_u12_u4_n129 ) , .A1( u1_u12_u4_n134 ) , .A2( u1_u12_u4_n148 ) );
  AND3_X1 u1_u12_u4_U25 (.A1( u1_u12_u4_n119 ) , .A2( u1_u12_u4_n143 ) , .A3( u1_u12_u4_n154 ) , .ZN( u1_u12_u4_n161 ) );
  AND2_X1 u1_u12_u4_U26 (.A1( u1_u12_u4_n145 ) , .A2( u1_u12_u4_n147 ) , .ZN( u1_u12_u4_n159 ) );
  OR3_X1 u1_u12_u4_U27 (.A3( u1_u12_u4_n114 ) , .A2( u1_u12_u4_n115 ) , .A1( u1_u12_u4_n116 ) , .ZN( u1_u12_u4_n136 ) );
  AOI21_X1 u1_u12_u4_U28 (.A( u1_u12_u4_n113 ) , .ZN( u1_u12_u4_n116 ) , .B2( u1_u12_u4_n173 ) , .B1( u1_u12_u4_n174 ) );
  AOI21_X1 u1_u12_u4_U29 (.ZN( u1_u12_u4_n115 ) , .B2( u1_u12_u4_n145 ) , .B1( u1_u12_u4_n146 ) , .A( u1_u12_u4_n156 ) );
  NOR2_X1 u1_u12_u4_U3 (.ZN( u1_u12_u4_n121 ) , .A1( u1_u12_u4_n181 ) , .A2( u1_u12_u4_n182 ) );
  OAI22_X1 u1_u12_u4_U30 (.ZN( u1_u12_u4_n114 ) , .A2( u1_u12_u4_n121 ) , .B1( u1_u12_u4_n160 ) , .B2( u1_u12_u4_n170 ) , .A1( u1_u12_u4_n171 ) );
  INV_X1 u1_u12_u4_U31 (.A( u1_u12_u4_n158 ) , .ZN( u1_u12_u4_n182 ) );
  INV_X1 u1_u12_u4_U32 (.ZN( u1_u12_u4_n181 ) , .A( u1_u12_u4_n96 ) );
  INV_X1 u1_u12_u4_U33 (.A( u1_u12_u4_n144 ) , .ZN( u1_u12_u4_n179 ) );
  INV_X1 u1_u12_u4_U34 (.A( u1_u12_u4_n157 ) , .ZN( u1_u12_u4_n178 ) );
  NAND2_X1 u1_u12_u4_U35 (.A2( u1_u12_u4_n154 ) , .A1( u1_u12_u4_n96 ) , .ZN( u1_u12_u4_n97 ) );
  INV_X1 u1_u12_u4_U36 (.ZN( u1_u12_u4_n186 ) , .A( u1_u12_u4_n95 ) );
  OAI221_X1 u1_u12_u4_U37 (.C1( u1_u12_u4_n134 ) , .B1( u1_u12_u4_n158 ) , .B2( u1_u12_u4_n171 ) , .C2( u1_u12_u4_n173 ) , .A( u1_u12_u4_n94 ) , .ZN( u1_u12_u4_n95 ) );
  AOI222_X1 u1_u12_u4_U38 (.B2( u1_u12_u4_n132 ) , .A1( u1_u12_u4_n138 ) , .C2( u1_u12_u4_n175 ) , .A2( u1_u12_u4_n179 ) , .C1( u1_u12_u4_n181 ) , .B1( u1_u12_u4_n185 ) , .ZN( u1_u12_u4_n94 ) );
  INV_X1 u1_u12_u4_U39 (.A( u1_u12_u4_n113 ) , .ZN( u1_u12_u4_n185 ) );
  INV_X1 u1_u12_u4_U4 (.A( u1_u12_u4_n117 ) , .ZN( u1_u12_u4_n184 ) );
  INV_X1 u1_u12_u4_U40 (.A( u1_u12_u4_n143 ) , .ZN( u1_u12_u4_n183 ) );
  NOR2_X1 u1_u12_u4_U41 (.ZN( u1_u12_u4_n138 ) , .A1( u1_u12_u4_n168 ) , .A2( u1_u12_u4_n169 ) );
  NOR2_X1 u1_u12_u4_U42 (.A1( u1_u12_u4_n150 ) , .A2( u1_u12_u4_n152 ) , .ZN( u1_u12_u4_n153 ) );
  NOR2_X1 u1_u12_u4_U43 (.A2( u1_u12_u4_n128 ) , .A1( u1_u12_u4_n138 ) , .ZN( u1_u12_u4_n156 ) );
  AOI22_X1 u1_u12_u4_U44 (.B2( u1_u12_u4_n122 ) , .A1( u1_u12_u4_n123 ) , .ZN( u1_u12_u4_n124 ) , .B1( u1_u12_u4_n128 ) , .A2( u1_u12_u4_n172 ) );
  INV_X1 u1_u12_u4_U45 (.A( u1_u12_u4_n153 ) , .ZN( u1_u12_u4_n172 ) );
  NAND2_X1 u1_u12_u4_U46 (.A2( u1_u12_u4_n120 ) , .ZN( u1_u12_u4_n123 ) , .A1( u1_u12_u4_n161 ) );
  AOI22_X1 u1_u12_u4_U47 (.B2( u1_u12_u4_n132 ) , .A2( u1_u12_u4_n133 ) , .ZN( u1_u12_u4_n140 ) , .A1( u1_u12_u4_n150 ) , .B1( u1_u12_u4_n179 ) );
  NAND2_X1 u1_u12_u4_U48 (.ZN( u1_u12_u4_n133 ) , .A2( u1_u12_u4_n146 ) , .A1( u1_u12_u4_n154 ) );
  NAND2_X1 u1_u12_u4_U49 (.A1( u1_u12_u4_n103 ) , .ZN( u1_u12_u4_n154 ) , .A2( u1_u12_u4_n98 ) );
  NOR4_X1 u1_u12_u4_U5 (.A4( u1_u12_u4_n106 ) , .A3( u1_u12_u4_n107 ) , .A2( u1_u12_u4_n108 ) , .A1( u1_u12_u4_n109 ) , .ZN( u1_u12_u4_n110 ) );
  NAND2_X1 u1_u12_u4_U50 (.A1( u1_u12_u4_n101 ) , .ZN( u1_u12_u4_n158 ) , .A2( u1_u12_u4_n99 ) );
  AOI21_X1 u1_u12_u4_U51 (.ZN( u1_u12_u4_n127 ) , .A( u1_u12_u4_n136 ) , .B2( u1_u12_u4_n150 ) , .B1( u1_u12_u4_n180 ) );
  INV_X1 u1_u12_u4_U52 (.A( u1_u12_u4_n160 ) , .ZN( u1_u12_u4_n180 ) );
  NAND2_X1 u1_u12_u4_U53 (.A2( u1_u12_u4_n104 ) , .A1( u1_u12_u4_n105 ) , .ZN( u1_u12_u4_n146 ) );
  NAND2_X1 u1_u12_u4_U54 (.A2( u1_u12_u4_n101 ) , .A1( u1_u12_u4_n102 ) , .ZN( u1_u12_u4_n160 ) );
  NAND2_X1 u1_u12_u4_U55 (.ZN( u1_u12_u4_n134 ) , .A1( u1_u12_u4_n98 ) , .A2( u1_u12_u4_n99 ) );
  NAND2_X1 u1_u12_u4_U56 (.A1( u1_u12_u4_n103 ) , .A2( u1_u12_u4_n104 ) , .ZN( u1_u12_u4_n143 ) );
  NAND2_X1 u1_u12_u4_U57 (.A2( u1_u12_u4_n105 ) , .ZN( u1_u12_u4_n145 ) , .A1( u1_u12_u4_n98 ) );
  NAND2_X1 u1_u12_u4_U58 (.A1( u1_u12_u4_n100 ) , .A2( u1_u12_u4_n105 ) , .ZN( u1_u12_u4_n120 ) );
  NAND2_X1 u1_u12_u4_U59 (.A1( u1_u12_u4_n102 ) , .A2( u1_u12_u4_n104 ) , .ZN( u1_u12_u4_n148 ) );
  AOI21_X1 u1_u12_u4_U6 (.ZN( u1_u12_u4_n106 ) , .B2( u1_u12_u4_n146 ) , .B1( u1_u12_u4_n158 ) , .A( u1_u12_u4_n170 ) );
  NAND2_X1 u1_u12_u4_U60 (.A2( u1_u12_u4_n100 ) , .A1( u1_u12_u4_n103 ) , .ZN( u1_u12_u4_n157 ) );
  INV_X1 u1_u12_u4_U61 (.A( u1_u12_u4_n150 ) , .ZN( u1_u12_u4_n173 ) );
  INV_X1 u1_u12_u4_U62 (.A( u1_u12_u4_n152 ) , .ZN( u1_u12_u4_n171 ) );
  NAND2_X1 u1_u12_u4_U63 (.A1( u1_u12_u4_n100 ) , .ZN( u1_u12_u4_n118 ) , .A2( u1_u12_u4_n99 ) );
  NAND2_X1 u1_u12_u4_U64 (.A2( u1_u12_u4_n100 ) , .A1( u1_u12_u4_n102 ) , .ZN( u1_u12_u4_n144 ) );
  NAND2_X1 u1_u12_u4_U65 (.A2( u1_u12_u4_n101 ) , .A1( u1_u12_u4_n105 ) , .ZN( u1_u12_u4_n96 ) );
  INV_X1 u1_u12_u4_U66 (.A( u1_u12_u4_n128 ) , .ZN( u1_u12_u4_n174 ) );
  NAND2_X1 u1_u12_u4_U67 (.A2( u1_u12_u4_n102 ) , .ZN( u1_u12_u4_n119 ) , .A1( u1_u12_u4_n98 ) );
  NAND2_X1 u1_u12_u4_U68 (.A2( u1_u12_u4_n101 ) , .A1( u1_u12_u4_n103 ) , .ZN( u1_u12_u4_n147 ) );
  NAND2_X1 u1_u12_u4_U69 (.A2( u1_u12_u4_n104 ) , .ZN( u1_u12_u4_n113 ) , .A1( u1_u12_u4_n99 ) );
  AOI21_X1 u1_u12_u4_U7 (.ZN( u1_u12_u4_n108 ) , .B2( u1_u12_u4_n134 ) , .B1( u1_u12_u4_n155 ) , .A( u1_u12_u4_n156 ) );
  NOR2_X1 u1_u12_u4_U70 (.A2( u1_u12_X_28 ) , .ZN( u1_u12_u4_n150 ) , .A1( u1_u12_u4_n168 ) );
  NOR2_X1 u1_u12_u4_U71 (.A2( u1_u12_X_29 ) , .ZN( u1_u12_u4_n152 ) , .A1( u1_u12_u4_n169 ) );
  NOR2_X1 u1_u12_u4_U72 (.A2( u1_u12_X_30 ) , .ZN( u1_u12_u4_n105 ) , .A1( u1_u12_u4_n176 ) );
  NOR2_X1 u1_u12_u4_U73 (.A2( u1_u12_X_26 ) , .ZN( u1_u12_u4_n100 ) , .A1( u1_u12_u4_n177 ) );
  NOR2_X1 u1_u12_u4_U74 (.A2( u1_u12_X_28 ) , .A1( u1_u12_X_29 ) , .ZN( u1_u12_u4_n128 ) );
  NOR2_X1 u1_u12_u4_U75 (.A2( u1_u12_X_27 ) , .A1( u1_u12_X_30 ) , .ZN( u1_u12_u4_n102 ) );
  NOR2_X1 u1_u12_u4_U76 (.A2( u1_u12_X_25 ) , .A1( u1_u12_X_26 ) , .ZN( u1_u12_u4_n98 ) );
  AND2_X1 u1_u12_u4_U77 (.A2( u1_u12_X_25 ) , .A1( u1_u12_X_26 ) , .ZN( u1_u12_u4_n104 ) );
  AND2_X1 u1_u12_u4_U78 (.A1( u1_u12_X_30 ) , .A2( u1_u12_u4_n176 ) , .ZN( u1_u12_u4_n99 ) );
  AND2_X1 u1_u12_u4_U79 (.A1( u1_u12_X_26 ) , .ZN( u1_u12_u4_n101 ) , .A2( u1_u12_u4_n177 ) );
  AOI21_X1 u1_u12_u4_U8 (.ZN( u1_u12_u4_n109 ) , .A( u1_u12_u4_n153 ) , .B1( u1_u12_u4_n159 ) , .B2( u1_u12_u4_n184 ) );
  AND2_X1 u1_u12_u4_U80 (.A1( u1_u12_X_27 ) , .A2( u1_u12_X_30 ) , .ZN( u1_u12_u4_n103 ) );
  INV_X1 u1_u12_u4_U81 (.A( u1_u12_X_28 ) , .ZN( u1_u12_u4_n169 ) );
  INV_X1 u1_u12_u4_U82 (.A( u1_u12_X_29 ) , .ZN( u1_u12_u4_n168 ) );
  INV_X1 u1_u12_u4_U83 (.A( u1_u12_X_25 ) , .ZN( u1_u12_u4_n177 ) );
  INV_X1 u1_u12_u4_U84 (.A( u1_u12_X_27 ) , .ZN( u1_u12_u4_n176 ) );
  NAND4_X1 u1_u12_u4_U85 (.ZN( u1_out12_25 ) , .A4( u1_u12_u4_n139 ) , .A3( u1_u12_u4_n140 ) , .A2( u1_u12_u4_n141 ) , .A1( u1_u12_u4_n142 ) );
  OAI21_X1 u1_u12_u4_U86 (.A( u1_u12_u4_n128 ) , .B2( u1_u12_u4_n129 ) , .B1( u1_u12_u4_n130 ) , .ZN( u1_u12_u4_n142 ) );
  OAI21_X1 u1_u12_u4_U87 (.B2( u1_u12_u4_n131 ) , .ZN( u1_u12_u4_n141 ) , .A( u1_u12_u4_n175 ) , .B1( u1_u12_u4_n183 ) );
  NAND4_X1 u1_u12_u4_U88 (.ZN( u1_out12_14 ) , .A4( u1_u12_u4_n124 ) , .A3( u1_u12_u4_n125 ) , .A2( u1_u12_u4_n126 ) , .A1( u1_u12_u4_n127 ) );
  AOI22_X1 u1_u12_u4_U89 (.B2( u1_u12_u4_n117 ) , .ZN( u1_u12_u4_n126 ) , .A1( u1_u12_u4_n129 ) , .B1( u1_u12_u4_n152 ) , .A2( u1_u12_u4_n175 ) );
  AOI211_X1 u1_u12_u4_U9 (.B( u1_u12_u4_n136 ) , .A( u1_u12_u4_n137 ) , .C2( u1_u12_u4_n138 ) , .ZN( u1_u12_u4_n139 ) , .C1( u1_u12_u4_n182 ) );
  AOI22_X1 u1_u12_u4_U90 (.ZN( u1_u12_u4_n125 ) , .B2( u1_u12_u4_n131 ) , .A2( u1_u12_u4_n132 ) , .B1( u1_u12_u4_n138 ) , .A1( u1_u12_u4_n178 ) );
  NAND4_X1 u1_u12_u4_U91 (.ZN( u1_out12_8 ) , .A4( u1_u12_u4_n110 ) , .A3( u1_u12_u4_n111 ) , .A2( u1_u12_u4_n112 ) , .A1( u1_u12_u4_n186 ) );
  NAND2_X1 u1_u12_u4_U92 (.ZN( u1_u12_u4_n112 ) , .A2( u1_u12_u4_n130 ) , .A1( u1_u12_u4_n150 ) );
  AOI22_X1 u1_u12_u4_U93 (.ZN( u1_u12_u4_n111 ) , .B2( u1_u12_u4_n132 ) , .A1( u1_u12_u4_n152 ) , .B1( u1_u12_u4_n178 ) , .A2( u1_u12_u4_n97 ) );
  AOI22_X1 u1_u12_u4_U94 (.B2( u1_u12_u4_n149 ) , .B1( u1_u12_u4_n150 ) , .A2( u1_u12_u4_n151 ) , .A1( u1_u12_u4_n152 ) , .ZN( u1_u12_u4_n167 ) );
  NOR4_X1 u1_u12_u4_U95 (.A4( u1_u12_u4_n162 ) , .A3( u1_u12_u4_n163 ) , .A2( u1_u12_u4_n164 ) , .A1( u1_u12_u4_n165 ) , .ZN( u1_u12_u4_n166 ) );
  NAND3_X1 u1_u12_u4_U96 (.ZN( u1_out12_3 ) , .A3( u1_u12_u4_n166 ) , .A1( u1_u12_u4_n167 ) , .A2( u1_u12_u4_n186 ) );
  NAND3_X1 u1_u12_u4_U97 (.A3( u1_u12_u4_n146 ) , .A2( u1_u12_u4_n147 ) , .A1( u1_u12_u4_n148 ) , .ZN( u1_u12_u4_n149 ) );
  NAND3_X1 u1_u12_u4_U98 (.A3( u1_u12_u4_n143 ) , .A2( u1_u12_u4_n144 ) , .A1( u1_u12_u4_n145 ) , .ZN( u1_u12_u4_n151 ) );
  NAND3_X1 u1_u12_u4_U99 (.A3( u1_u12_u4_n121 ) , .ZN( u1_u12_u4_n122 ) , .A2( u1_u12_u4_n144 ) , .A1( u1_u12_u4_n154 ) );
  INV_X1 u1_u12_u5_U10 (.A( u1_u12_u5_n121 ) , .ZN( u1_u12_u5_n177 ) );
  NOR3_X1 u1_u12_u5_U100 (.A3( u1_u12_u5_n141 ) , .A1( u1_u12_u5_n142 ) , .ZN( u1_u12_u5_n143 ) , .A2( u1_u12_u5_n191 ) );
  NAND4_X1 u1_u12_u5_U101 (.ZN( u1_out12_4 ) , .A4( u1_u12_u5_n112 ) , .A2( u1_u12_u5_n113 ) , .A1( u1_u12_u5_n114 ) , .A3( u1_u12_u5_n195 ) );
  AOI211_X1 u1_u12_u5_U102 (.A( u1_u12_u5_n110 ) , .C1( u1_u12_u5_n111 ) , .ZN( u1_u12_u5_n112 ) , .B( u1_u12_u5_n118 ) , .C2( u1_u12_u5_n177 ) );
  AOI222_X1 u1_u12_u5_U103 (.ZN( u1_u12_u5_n113 ) , .A1( u1_u12_u5_n131 ) , .C1( u1_u12_u5_n148 ) , .B2( u1_u12_u5_n174 ) , .C2( u1_u12_u5_n178 ) , .A2( u1_u12_u5_n179 ) , .B1( u1_u12_u5_n99 ) );
  NAND3_X1 u1_u12_u5_U104 (.A2( u1_u12_u5_n154 ) , .A3( u1_u12_u5_n158 ) , .A1( u1_u12_u5_n161 ) , .ZN( u1_u12_u5_n99 ) );
  NOR2_X1 u1_u12_u5_U11 (.ZN( u1_u12_u5_n160 ) , .A2( u1_u12_u5_n173 ) , .A1( u1_u12_u5_n177 ) );
  INV_X1 u1_u12_u5_U12 (.A( u1_u12_u5_n150 ) , .ZN( u1_u12_u5_n174 ) );
  AOI21_X1 u1_u12_u5_U13 (.A( u1_u12_u5_n160 ) , .B2( u1_u12_u5_n161 ) , .ZN( u1_u12_u5_n162 ) , .B1( u1_u12_u5_n192 ) );
  INV_X1 u1_u12_u5_U14 (.A( u1_u12_u5_n159 ) , .ZN( u1_u12_u5_n192 ) );
  AOI21_X1 u1_u12_u5_U15 (.A( u1_u12_u5_n156 ) , .B2( u1_u12_u5_n157 ) , .B1( u1_u12_u5_n158 ) , .ZN( u1_u12_u5_n163 ) );
  AOI21_X1 u1_u12_u5_U16 (.B2( u1_u12_u5_n139 ) , .B1( u1_u12_u5_n140 ) , .ZN( u1_u12_u5_n141 ) , .A( u1_u12_u5_n150 ) );
  OAI21_X1 u1_u12_u5_U17 (.A( u1_u12_u5_n133 ) , .B2( u1_u12_u5_n134 ) , .B1( u1_u12_u5_n135 ) , .ZN( u1_u12_u5_n142 ) );
  OAI21_X1 u1_u12_u5_U18 (.ZN( u1_u12_u5_n133 ) , .B2( u1_u12_u5_n147 ) , .A( u1_u12_u5_n173 ) , .B1( u1_u12_u5_n188 ) );
  NAND2_X1 u1_u12_u5_U19 (.A2( u1_u12_u5_n119 ) , .A1( u1_u12_u5_n123 ) , .ZN( u1_u12_u5_n137 ) );
  INV_X1 u1_u12_u5_U20 (.A( u1_u12_u5_n155 ) , .ZN( u1_u12_u5_n194 ) );
  NAND2_X1 u1_u12_u5_U21 (.A1( u1_u12_u5_n121 ) , .ZN( u1_u12_u5_n132 ) , .A2( u1_u12_u5_n172 ) );
  NAND2_X1 u1_u12_u5_U22 (.A2( u1_u12_u5_n122 ) , .ZN( u1_u12_u5_n136 ) , .A1( u1_u12_u5_n154 ) );
  NAND2_X1 u1_u12_u5_U23 (.A2( u1_u12_u5_n119 ) , .A1( u1_u12_u5_n120 ) , .ZN( u1_u12_u5_n159 ) );
  INV_X1 u1_u12_u5_U24 (.A( u1_u12_u5_n156 ) , .ZN( u1_u12_u5_n175 ) );
  INV_X1 u1_u12_u5_U25 (.A( u1_u12_u5_n158 ) , .ZN( u1_u12_u5_n188 ) );
  INV_X1 u1_u12_u5_U26 (.A( u1_u12_u5_n152 ) , .ZN( u1_u12_u5_n179 ) );
  INV_X1 u1_u12_u5_U27 (.A( u1_u12_u5_n140 ) , .ZN( u1_u12_u5_n182 ) );
  INV_X1 u1_u12_u5_U28 (.A( u1_u12_u5_n151 ) , .ZN( u1_u12_u5_n183 ) );
  INV_X1 u1_u12_u5_U29 (.A( u1_u12_u5_n123 ) , .ZN( u1_u12_u5_n185 ) );
  NOR2_X1 u1_u12_u5_U3 (.ZN( u1_u12_u5_n134 ) , .A1( u1_u12_u5_n183 ) , .A2( u1_u12_u5_n190 ) );
  INV_X1 u1_u12_u5_U30 (.A( u1_u12_u5_n161 ) , .ZN( u1_u12_u5_n184 ) );
  INV_X1 u1_u12_u5_U31 (.A( u1_u12_u5_n139 ) , .ZN( u1_u12_u5_n189 ) );
  INV_X1 u1_u12_u5_U32 (.A( u1_u12_u5_n157 ) , .ZN( u1_u12_u5_n190 ) );
  INV_X1 u1_u12_u5_U33 (.A( u1_u12_u5_n120 ) , .ZN( u1_u12_u5_n193 ) );
  NAND2_X1 u1_u12_u5_U34 (.ZN( u1_u12_u5_n111 ) , .A1( u1_u12_u5_n140 ) , .A2( u1_u12_u5_n155 ) );
  NOR2_X1 u1_u12_u5_U35 (.ZN( u1_u12_u5_n100 ) , .A1( u1_u12_u5_n170 ) , .A2( u1_u12_u5_n180 ) );
  INV_X1 u1_u12_u5_U36 (.A( u1_u12_u5_n117 ) , .ZN( u1_u12_u5_n196 ) );
  OAI221_X1 u1_u12_u5_U37 (.A( u1_u12_u5_n116 ) , .ZN( u1_u12_u5_n117 ) , .B2( u1_u12_u5_n119 ) , .C1( u1_u12_u5_n153 ) , .C2( u1_u12_u5_n158 ) , .B1( u1_u12_u5_n172 ) );
  AOI222_X1 u1_u12_u5_U38 (.ZN( u1_u12_u5_n116 ) , .B2( u1_u12_u5_n145 ) , .C1( u1_u12_u5_n148 ) , .A2( u1_u12_u5_n174 ) , .C2( u1_u12_u5_n177 ) , .B1( u1_u12_u5_n187 ) , .A1( u1_u12_u5_n193 ) );
  INV_X1 u1_u12_u5_U39 (.A( u1_u12_u5_n115 ) , .ZN( u1_u12_u5_n187 ) );
  INV_X1 u1_u12_u5_U4 (.A( u1_u12_u5_n138 ) , .ZN( u1_u12_u5_n191 ) );
  AOI22_X1 u1_u12_u5_U40 (.B2( u1_u12_u5_n131 ) , .A2( u1_u12_u5_n146 ) , .ZN( u1_u12_u5_n169 ) , .B1( u1_u12_u5_n174 ) , .A1( u1_u12_u5_n185 ) );
  NOR2_X1 u1_u12_u5_U41 (.A1( u1_u12_u5_n146 ) , .ZN( u1_u12_u5_n150 ) , .A2( u1_u12_u5_n173 ) );
  AOI21_X1 u1_u12_u5_U42 (.A( u1_u12_u5_n118 ) , .B2( u1_u12_u5_n145 ) , .ZN( u1_u12_u5_n168 ) , .B1( u1_u12_u5_n186 ) );
  INV_X1 u1_u12_u5_U43 (.A( u1_u12_u5_n122 ) , .ZN( u1_u12_u5_n186 ) );
  NOR2_X1 u1_u12_u5_U44 (.A1( u1_u12_u5_n146 ) , .ZN( u1_u12_u5_n152 ) , .A2( u1_u12_u5_n176 ) );
  NOR2_X1 u1_u12_u5_U45 (.A1( u1_u12_u5_n115 ) , .ZN( u1_u12_u5_n118 ) , .A2( u1_u12_u5_n153 ) );
  NOR2_X1 u1_u12_u5_U46 (.A2( u1_u12_u5_n145 ) , .ZN( u1_u12_u5_n156 ) , .A1( u1_u12_u5_n174 ) );
  NOR2_X1 u1_u12_u5_U47 (.ZN( u1_u12_u5_n121 ) , .A2( u1_u12_u5_n145 ) , .A1( u1_u12_u5_n176 ) );
  AOI22_X1 u1_u12_u5_U48 (.ZN( u1_u12_u5_n114 ) , .A2( u1_u12_u5_n137 ) , .A1( u1_u12_u5_n145 ) , .B2( u1_u12_u5_n175 ) , .B1( u1_u12_u5_n193 ) );
  OAI211_X1 u1_u12_u5_U49 (.B( u1_u12_u5_n124 ) , .A( u1_u12_u5_n125 ) , .C2( u1_u12_u5_n126 ) , .C1( u1_u12_u5_n127 ) , .ZN( u1_u12_u5_n128 ) );
  OAI21_X1 u1_u12_u5_U5 (.B2( u1_u12_u5_n136 ) , .B1( u1_u12_u5_n137 ) , .ZN( u1_u12_u5_n138 ) , .A( u1_u12_u5_n177 ) );
  NOR3_X1 u1_u12_u5_U50 (.ZN( u1_u12_u5_n127 ) , .A1( u1_u12_u5_n136 ) , .A3( u1_u12_u5_n148 ) , .A2( u1_u12_u5_n182 ) );
  OAI21_X1 u1_u12_u5_U51 (.ZN( u1_u12_u5_n124 ) , .A( u1_u12_u5_n177 ) , .B2( u1_u12_u5_n183 ) , .B1( u1_u12_u5_n189 ) );
  OAI21_X1 u1_u12_u5_U52 (.ZN( u1_u12_u5_n125 ) , .A( u1_u12_u5_n174 ) , .B2( u1_u12_u5_n185 ) , .B1( u1_u12_u5_n190 ) );
  AOI21_X1 u1_u12_u5_U53 (.A( u1_u12_u5_n153 ) , .B2( u1_u12_u5_n154 ) , .B1( u1_u12_u5_n155 ) , .ZN( u1_u12_u5_n164 ) );
  AOI21_X1 u1_u12_u5_U54 (.ZN( u1_u12_u5_n110 ) , .B1( u1_u12_u5_n122 ) , .B2( u1_u12_u5_n139 ) , .A( u1_u12_u5_n153 ) );
  INV_X1 u1_u12_u5_U55 (.A( u1_u12_u5_n153 ) , .ZN( u1_u12_u5_n176 ) );
  INV_X1 u1_u12_u5_U56 (.A( u1_u12_u5_n126 ) , .ZN( u1_u12_u5_n173 ) );
  AND2_X1 u1_u12_u5_U57 (.A2( u1_u12_u5_n104 ) , .A1( u1_u12_u5_n107 ) , .ZN( u1_u12_u5_n147 ) );
  AND2_X1 u1_u12_u5_U58 (.A2( u1_u12_u5_n104 ) , .A1( u1_u12_u5_n108 ) , .ZN( u1_u12_u5_n148 ) );
  NAND2_X1 u1_u12_u5_U59 (.A1( u1_u12_u5_n105 ) , .A2( u1_u12_u5_n106 ) , .ZN( u1_u12_u5_n158 ) );
  INV_X1 u1_u12_u5_U6 (.A( u1_u12_u5_n135 ) , .ZN( u1_u12_u5_n178 ) );
  NAND2_X1 u1_u12_u5_U60 (.A2( u1_u12_u5_n108 ) , .A1( u1_u12_u5_n109 ) , .ZN( u1_u12_u5_n139 ) );
  NAND2_X1 u1_u12_u5_U61 (.A1( u1_u12_u5_n106 ) , .A2( u1_u12_u5_n108 ) , .ZN( u1_u12_u5_n119 ) );
  NAND2_X1 u1_u12_u5_U62 (.A2( u1_u12_u5_n103 ) , .A1( u1_u12_u5_n105 ) , .ZN( u1_u12_u5_n140 ) );
  NAND2_X1 u1_u12_u5_U63 (.A2( u1_u12_u5_n104 ) , .A1( u1_u12_u5_n105 ) , .ZN( u1_u12_u5_n155 ) );
  NAND2_X1 u1_u12_u5_U64 (.A2( u1_u12_u5_n106 ) , .A1( u1_u12_u5_n107 ) , .ZN( u1_u12_u5_n122 ) );
  NAND2_X1 u1_u12_u5_U65 (.A2( u1_u12_u5_n100 ) , .A1( u1_u12_u5_n106 ) , .ZN( u1_u12_u5_n115 ) );
  NAND2_X1 u1_u12_u5_U66 (.A2( u1_u12_u5_n100 ) , .A1( u1_u12_u5_n103 ) , .ZN( u1_u12_u5_n161 ) );
  NAND2_X1 u1_u12_u5_U67 (.A1( u1_u12_u5_n105 ) , .A2( u1_u12_u5_n109 ) , .ZN( u1_u12_u5_n154 ) );
  INV_X1 u1_u12_u5_U68 (.A( u1_u12_u5_n146 ) , .ZN( u1_u12_u5_n172 ) );
  NAND2_X1 u1_u12_u5_U69 (.A1( u1_u12_u5_n103 ) , .A2( u1_u12_u5_n108 ) , .ZN( u1_u12_u5_n123 ) );
  OAI22_X1 u1_u12_u5_U7 (.B2( u1_u12_u5_n149 ) , .B1( u1_u12_u5_n150 ) , .A2( u1_u12_u5_n151 ) , .A1( u1_u12_u5_n152 ) , .ZN( u1_u12_u5_n165 ) );
  NAND2_X1 u1_u12_u5_U70 (.A2( u1_u12_u5_n103 ) , .A1( u1_u12_u5_n107 ) , .ZN( u1_u12_u5_n151 ) );
  NAND2_X1 u1_u12_u5_U71 (.A2( u1_u12_u5_n107 ) , .A1( u1_u12_u5_n109 ) , .ZN( u1_u12_u5_n120 ) );
  NAND2_X1 u1_u12_u5_U72 (.A2( u1_u12_u5_n100 ) , .A1( u1_u12_u5_n109 ) , .ZN( u1_u12_u5_n157 ) );
  AND2_X1 u1_u12_u5_U73 (.A2( u1_u12_u5_n100 ) , .A1( u1_u12_u5_n104 ) , .ZN( u1_u12_u5_n131 ) );
  INV_X1 u1_u12_u5_U74 (.A( u1_u12_u5_n102 ) , .ZN( u1_u12_u5_n195 ) );
  OAI221_X1 u1_u12_u5_U75 (.A( u1_u12_u5_n101 ) , .ZN( u1_u12_u5_n102 ) , .C2( u1_u12_u5_n115 ) , .C1( u1_u12_u5_n126 ) , .B1( u1_u12_u5_n134 ) , .B2( u1_u12_u5_n160 ) );
  OAI21_X1 u1_u12_u5_U76 (.ZN( u1_u12_u5_n101 ) , .B1( u1_u12_u5_n137 ) , .A( u1_u12_u5_n146 ) , .B2( u1_u12_u5_n147 ) );
  NOR2_X1 u1_u12_u5_U77 (.A2( u1_u12_X_34 ) , .A1( u1_u12_X_35 ) , .ZN( u1_u12_u5_n145 ) );
  NOR2_X1 u1_u12_u5_U78 (.A2( u1_u12_X_34 ) , .ZN( u1_u12_u5_n146 ) , .A1( u1_u12_u5_n171 ) );
  NOR2_X1 u1_u12_u5_U79 (.A2( u1_u12_X_31 ) , .A1( u1_u12_X_32 ) , .ZN( u1_u12_u5_n103 ) );
  NOR3_X1 u1_u12_u5_U8 (.A2( u1_u12_u5_n147 ) , .A1( u1_u12_u5_n148 ) , .ZN( u1_u12_u5_n149 ) , .A3( u1_u12_u5_n194 ) );
  NOR2_X1 u1_u12_u5_U80 (.A2( u1_u12_X_36 ) , .ZN( u1_u12_u5_n105 ) , .A1( u1_u12_u5_n180 ) );
  NOR2_X1 u1_u12_u5_U81 (.A2( u1_u12_X_33 ) , .ZN( u1_u12_u5_n108 ) , .A1( u1_u12_u5_n170 ) );
  NOR2_X1 u1_u12_u5_U82 (.A2( u1_u12_X_33 ) , .A1( u1_u12_X_36 ) , .ZN( u1_u12_u5_n107 ) );
  NOR2_X1 u1_u12_u5_U83 (.A2( u1_u12_X_31 ) , .ZN( u1_u12_u5_n104 ) , .A1( u1_u12_u5_n181 ) );
  NAND2_X1 u1_u12_u5_U84 (.A2( u1_u12_X_34 ) , .A1( u1_u12_X_35 ) , .ZN( u1_u12_u5_n153 ) );
  NAND2_X1 u1_u12_u5_U85 (.A1( u1_u12_X_34 ) , .ZN( u1_u12_u5_n126 ) , .A2( u1_u12_u5_n171 ) );
  AND2_X1 u1_u12_u5_U86 (.A1( u1_u12_X_31 ) , .A2( u1_u12_X_32 ) , .ZN( u1_u12_u5_n106 ) );
  AND2_X1 u1_u12_u5_U87 (.A1( u1_u12_X_31 ) , .ZN( u1_u12_u5_n109 ) , .A2( u1_u12_u5_n181 ) );
  INV_X1 u1_u12_u5_U88 (.A( u1_u12_X_33 ) , .ZN( u1_u12_u5_n180 ) );
  INV_X1 u1_u12_u5_U89 (.A( u1_u12_X_35 ) , .ZN( u1_u12_u5_n171 ) );
  NOR2_X1 u1_u12_u5_U9 (.ZN( u1_u12_u5_n135 ) , .A1( u1_u12_u5_n173 ) , .A2( u1_u12_u5_n176 ) );
  INV_X1 u1_u12_u5_U90 (.A( u1_u12_X_36 ) , .ZN( u1_u12_u5_n170 ) );
  INV_X1 u1_u12_u5_U91 (.A( u1_u12_X_32 ) , .ZN( u1_u12_u5_n181 ) );
  NAND4_X1 u1_u12_u5_U92 (.ZN( u1_out12_29 ) , .A4( u1_u12_u5_n129 ) , .A3( u1_u12_u5_n130 ) , .A2( u1_u12_u5_n168 ) , .A1( u1_u12_u5_n196 ) );
  AOI221_X1 u1_u12_u5_U93 (.A( u1_u12_u5_n128 ) , .ZN( u1_u12_u5_n129 ) , .C2( u1_u12_u5_n132 ) , .B2( u1_u12_u5_n159 ) , .B1( u1_u12_u5_n176 ) , .C1( u1_u12_u5_n184 ) );
  AOI222_X1 u1_u12_u5_U94 (.ZN( u1_u12_u5_n130 ) , .A2( u1_u12_u5_n146 ) , .B1( u1_u12_u5_n147 ) , .C2( u1_u12_u5_n175 ) , .B2( u1_u12_u5_n179 ) , .A1( u1_u12_u5_n188 ) , .C1( u1_u12_u5_n194 ) );
  NAND4_X1 u1_u12_u5_U95 (.ZN( u1_out12_19 ) , .A4( u1_u12_u5_n166 ) , .A3( u1_u12_u5_n167 ) , .A2( u1_u12_u5_n168 ) , .A1( u1_u12_u5_n169 ) );
  AOI22_X1 u1_u12_u5_U96 (.B2( u1_u12_u5_n145 ) , .A2( u1_u12_u5_n146 ) , .ZN( u1_u12_u5_n167 ) , .B1( u1_u12_u5_n182 ) , .A1( u1_u12_u5_n189 ) );
  NOR4_X1 u1_u12_u5_U97 (.A4( u1_u12_u5_n162 ) , .A3( u1_u12_u5_n163 ) , .A2( u1_u12_u5_n164 ) , .A1( u1_u12_u5_n165 ) , .ZN( u1_u12_u5_n166 ) );
  NAND4_X1 u1_u12_u5_U98 (.ZN( u1_out12_11 ) , .A4( u1_u12_u5_n143 ) , .A3( u1_u12_u5_n144 ) , .A2( u1_u12_u5_n169 ) , .A1( u1_u12_u5_n196 ) );
  AOI22_X1 u1_u12_u5_U99 (.A2( u1_u12_u5_n132 ) , .ZN( u1_u12_u5_n144 ) , .B2( u1_u12_u5_n145 ) , .B1( u1_u12_u5_n184 ) , .A1( u1_u12_u5_n194 ) );
  XOR2_X1 u1_u13_U10 (.B( u1_K14_45 ) , .A( u1_R12_30 ) , .Z( u1_u13_X_45 ) );
  XOR2_X1 u1_u13_U11 (.B( u1_K14_44 ) , .A( u1_R12_29 ) , .Z( u1_u13_X_44 ) );
  XOR2_X1 u1_u13_U12 (.B( u1_K14_43 ) , .A( u1_R12_28 ) , .Z( u1_u13_X_43 ) );
  XOR2_X1 u1_u13_U13 (.B( u1_K14_42 ) , .A( u1_R12_29 ) , .Z( u1_u13_X_42 ) );
  XOR2_X1 u1_u13_U14 (.B( u1_K14_41 ) , .A( u1_R12_28 ) , .Z( u1_u13_X_41 ) );
  XOR2_X1 u1_u13_U15 (.B( u1_K14_40 ) , .A( u1_R12_27 ) , .Z( u1_u13_X_40 ) );
  XOR2_X1 u1_u13_U17 (.B( u1_K14_39 ) , .A( u1_R12_26 ) , .Z( u1_u13_X_39 ) );
  XOR2_X1 u1_u13_U18 (.B( u1_K14_38 ) , .A( u1_R12_25 ) , .Z( u1_u13_X_38 ) );
  XOR2_X1 u1_u13_U19 (.B( u1_K14_37 ) , .A( u1_R12_24 ) , .Z( u1_u13_X_37 ) );
  XOR2_X1 u1_u13_U7 (.B( u1_K14_48 ) , .A( u1_R12_1 ) , .Z( u1_u13_X_48 ) );
  XOR2_X1 u1_u13_U8 (.B( u1_K14_47 ) , .A( u1_R12_32 ) , .Z( u1_u13_X_47 ) );
  XOR2_X1 u1_u13_U9 (.B( u1_K14_46 ) , .A( u1_R12_31 ) , .Z( u1_u13_X_46 ) );
  AOI22_X1 u1_u13_u6_U10 (.A2( u1_u13_u6_n151 ) , .B2( u1_u13_u6_n161 ) , .A1( u1_u13_u6_n167 ) , .B1( u1_u13_u6_n170 ) , .ZN( u1_u13_u6_n89 ) );
  AOI21_X1 u1_u13_u6_U11 (.B1( u1_u13_u6_n107 ) , .B2( u1_u13_u6_n132 ) , .A( u1_u13_u6_n158 ) , .ZN( u1_u13_u6_n88 ) );
  AOI21_X1 u1_u13_u6_U12 (.B2( u1_u13_u6_n147 ) , .B1( u1_u13_u6_n148 ) , .ZN( u1_u13_u6_n149 ) , .A( u1_u13_u6_n158 ) );
  AOI21_X1 u1_u13_u6_U13 (.ZN( u1_u13_u6_n106 ) , .A( u1_u13_u6_n142 ) , .B2( u1_u13_u6_n159 ) , .B1( u1_u13_u6_n164 ) );
  INV_X1 u1_u13_u6_U14 (.A( u1_u13_u6_n155 ) , .ZN( u1_u13_u6_n161 ) );
  INV_X1 u1_u13_u6_U15 (.A( u1_u13_u6_n128 ) , .ZN( u1_u13_u6_n164 ) );
  NAND2_X1 u1_u13_u6_U16 (.ZN( u1_u13_u6_n110 ) , .A1( u1_u13_u6_n122 ) , .A2( u1_u13_u6_n129 ) );
  NAND2_X1 u1_u13_u6_U17 (.ZN( u1_u13_u6_n124 ) , .A2( u1_u13_u6_n146 ) , .A1( u1_u13_u6_n148 ) );
  INV_X1 u1_u13_u6_U18 (.A( u1_u13_u6_n132 ) , .ZN( u1_u13_u6_n171 ) );
  AND2_X1 u1_u13_u6_U19 (.A1( u1_u13_u6_n100 ) , .ZN( u1_u13_u6_n130 ) , .A2( u1_u13_u6_n147 ) );
  INV_X1 u1_u13_u6_U20 (.A( u1_u13_u6_n127 ) , .ZN( u1_u13_u6_n173 ) );
  INV_X1 u1_u13_u6_U21 (.A( u1_u13_u6_n121 ) , .ZN( u1_u13_u6_n167 ) );
  INV_X1 u1_u13_u6_U22 (.A( u1_u13_u6_n100 ) , .ZN( u1_u13_u6_n169 ) );
  INV_X1 u1_u13_u6_U23 (.A( u1_u13_u6_n123 ) , .ZN( u1_u13_u6_n170 ) );
  INV_X1 u1_u13_u6_U24 (.A( u1_u13_u6_n113 ) , .ZN( u1_u13_u6_n168 ) );
  AND2_X1 u1_u13_u6_U25 (.A1( u1_u13_u6_n107 ) , .A2( u1_u13_u6_n119 ) , .ZN( u1_u13_u6_n133 ) );
  AND2_X1 u1_u13_u6_U26 (.A2( u1_u13_u6_n121 ) , .A1( u1_u13_u6_n122 ) , .ZN( u1_u13_u6_n131 ) );
  AND3_X1 u1_u13_u6_U27 (.ZN( u1_u13_u6_n120 ) , .A2( u1_u13_u6_n127 ) , .A1( u1_u13_u6_n132 ) , .A3( u1_u13_u6_n145 ) );
  INV_X1 u1_u13_u6_U28 (.A( u1_u13_u6_n146 ) , .ZN( u1_u13_u6_n163 ) );
  AOI222_X1 u1_u13_u6_U29 (.ZN( u1_u13_u6_n114 ) , .A1( u1_u13_u6_n118 ) , .A2( u1_u13_u6_n126 ) , .B2( u1_u13_u6_n151 ) , .C2( u1_u13_u6_n159 ) , .C1( u1_u13_u6_n168 ) , .B1( u1_u13_u6_n169 ) );
  INV_X1 u1_u13_u6_U3 (.A( u1_u13_u6_n110 ) , .ZN( u1_u13_u6_n166 ) );
  NOR2_X1 u1_u13_u6_U30 (.A1( u1_u13_u6_n162 ) , .A2( u1_u13_u6_n165 ) , .ZN( u1_u13_u6_n98 ) );
  AOI211_X1 u1_u13_u6_U31 (.B( u1_u13_u6_n134 ) , .A( u1_u13_u6_n135 ) , .C1( u1_u13_u6_n136 ) , .ZN( u1_u13_u6_n137 ) , .C2( u1_u13_u6_n151 ) );
  AOI21_X1 u1_u13_u6_U32 (.B2( u1_u13_u6_n132 ) , .B1( u1_u13_u6_n133 ) , .ZN( u1_u13_u6_n134 ) , .A( u1_u13_u6_n158 ) );
  AOI21_X1 u1_u13_u6_U33 (.B1( u1_u13_u6_n131 ) , .ZN( u1_u13_u6_n135 ) , .A( u1_u13_u6_n144 ) , .B2( u1_u13_u6_n146 ) );
  NAND4_X1 u1_u13_u6_U34 (.A4( u1_u13_u6_n127 ) , .A3( u1_u13_u6_n128 ) , .A2( u1_u13_u6_n129 ) , .A1( u1_u13_u6_n130 ) , .ZN( u1_u13_u6_n136 ) );
  NAND2_X1 u1_u13_u6_U35 (.A1( u1_u13_u6_n144 ) , .ZN( u1_u13_u6_n151 ) , .A2( u1_u13_u6_n158 ) );
  NAND2_X1 u1_u13_u6_U36 (.ZN( u1_u13_u6_n132 ) , .A1( u1_u13_u6_n91 ) , .A2( u1_u13_u6_n97 ) );
  AOI22_X1 u1_u13_u6_U37 (.B2( u1_u13_u6_n110 ) , .B1( u1_u13_u6_n111 ) , .A1( u1_u13_u6_n112 ) , .ZN( u1_u13_u6_n115 ) , .A2( u1_u13_u6_n161 ) );
  NAND4_X1 u1_u13_u6_U38 (.A3( u1_u13_u6_n109 ) , .ZN( u1_u13_u6_n112 ) , .A4( u1_u13_u6_n132 ) , .A2( u1_u13_u6_n147 ) , .A1( u1_u13_u6_n166 ) );
  NOR2_X1 u1_u13_u6_U39 (.ZN( u1_u13_u6_n109 ) , .A1( u1_u13_u6_n170 ) , .A2( u1_u13_u6_n173 ) );
  INV_X1 u1_u13_u6_U4 (.A( u1_u13_u6_n142 ) , .ZN( u1_u13_u6_n174 ) );
  NOR2_X1 u1_u13_u6_U40 (.A2( u1_u13_u6_n126 ) , .ZN( u1_u13_u6_n155 ) , .A1( u1_u13_u6_n160 ) );
  NAND2_X1 u1_u13_u6_U41 (.ZN( u1_u13_u6_n146 ) , .A2( u1_u13_u6_n94 ) , .A1( u1_u13_u6_n99 ) );
  AOI21_X1 u1_u13_u6_U42 (.A( u1_u13_u6_n144 ) , .B2( u1_u13_u6_n145 ) , .B1( u1_u13_u6_n146 ) , .ZN( u1_u13_u6_n150 ) );
  INV_X1 u1_u13_u6_U43 (.A( u1_u13_u6_n111 ) , .ZN( u1_u13_u6_n158 ) );
  NAND2_X1 u1_u13_u6_U44 (.ZN( u1_u13_u6_n127 ) , .A1( u1_u13_u6_n91 ) , .A2( u1_u13_u6_n92 ) );
  NAND2_X1 u1_u13_u6_U45 (.ZN( u1_u13_u6_n129 ) , .A2( u1_u13_u6_n95 ) , .A1( u1_u13_u6_n96 ) );
  INV_X1 u1_u13_u6_U46 (.A( u1_u13_u6_n144 ) , .ZN( u1_u13_u6_n159 ) );
  NAND2_X1 u1_u13_u6_U47 (.ZN( u1_u13_u6_n145 ) , .A2( u1_u13_u6_n97 ) , .A1( u1_u13_u6_n98 ) );
  NAND2_X1 u1_u13_u6_U48 (.ZN( u1_u13_u6_n148 ) , .A2( u1_u13_u6_n92 ) , .A1( u1_u13_u6_n94 ) );
  NAND2_X1 u1_u13_u6_U49 (.ZN( u1_u13_u6_n108 ) , .A2( u1_u13_u6_n139 ) , .A1( u1_u13_u6_n144 ) );
  NAND2_X1 u1_u13_u6_U5 (.A2( u1_u13_u6_n143 ) , .ZN( u1_u13_u6_n152 ) , .A1( u1_u13_u6_n166 ) );
  NAND2_X1 u1_u13_u6_U50 (.ZN( u1_u13_u6_n121 ) , .A2( u1_u13_u6_n95 ) , .A1( u1_u13_u6_n97 ) );
  NAND2_X1 u1_u13_u6_U51 (.ZN( u1_u13_u6_n107 ) , .A2( u1_u13_u6_n92 ) , .A1( u1_u13_u6_n95 ) );
  AND2_X1 u1_u13_u6_U52 (.ZN( u1_u13_u6_n118 ) , .A2( u1_u13_u6_n91 ) , .A1( u1_u13_u6_n99 ) );
  NAND2_X1 u1_u13_u6_U53 (.ZN( u1_u13_u6_n147 ) , .A2( u1_u13_u6_n98 ) , .A1( u1_u13_u6_n99 ) );
  NAND2_X1 u1_u13_u6_U54 (.ZN( u1_u13_u6_n128 ) , .A1( u1_u13_u6_n94 ) , .A2( u1_u13_u6_n96 ) );
  NAND2_X1 u1_u13_u6_U55 (.ZN( u1_u13_u6_n119 ) , .A2( u1_u13_u6_n95 ) , .A1( u1_u13_u6_n99 ) );
  NAND2_X1 u1_u13_u6_U56 (.ZN( u1_u13_u6_n123 ) , .A2( u1_u13_u6_n91 ) , .A1( u1_u13_u6_n96 ) );
  NAND2_X1 u1_u13_u6_U57 (.ZN( u1_u13_u6_n100 ) , .A2( u1_u13_u6_n92 ) , .A1( u1_u13_u6_n98 ) );
  NAND2_X1 u1_u13_u6_U58 (.ZN( u1_u13_u6_n122 ) , .A1( u1_u13_u6_n94 ) , .A2( u1_u13_u6_n97 ) );
  INV_X1 u1_u13_u6_U59 (.A( u1_u13_u6_n139 ) , .ZN( u1_u13_u6_n160 ) );
  AOI22_X1 u1_u13_u6_U6 (.B2( u1_u13_u6_n101 ) , .A1( u1_u13_u6_n102 ) , .ZN( u1_u13_u6_n103 ) , .B1( u1_u13_u6_n160 ) , .A2( u1_u13_u6_n161 ) );
  NAND2_X1 u1_u13_u6_U60 (.ZN( u1_u13_u6_n113 ) , .A1( u1_u13_u6_n96 ) , .A2( u1_u13_u6_n98 ) );
  NOR2_X1 u1_u13_u6_U61 (.A2( u1_u13_X_40 ) , .A1( u1_u13_X_41 ) , .ZN( u1_u13_u6_n126 ) );
  NOR2_X1 u1_u13_u6_U62 (.A2( u1_u13_X_39 ) , .A1( u1_u13_X_42 ) , .ZN( u1_u13_u6_n92 ) );
  NOR2_X1 u1_u13_u6_U63 (.A2( u1_u13_X_39 ) , .A1( u1_u13_u6_n156 ) , .ZN( u1_u13_u6_n97 ) );
  NOR2_X1 u1_u13_u6_U64 (.A2( u1_u13_X_38 ) , .A1( u1_u13_u6_n165 ) , .ZN( u1_u13_u6_n95 ) );
  NOR2_X1 u1_u13_u6_U65 (.A2( u1_u13_X_41 ) , .ZN( u1_u13_u6_n111 ) , .A1( u1_u13_u6_n157 ) );
  NOR2_X1 u1_u13_u6_U66 (.A2( u1_u13_X_37 ) , .A1( u1_u13_u6_n162 ) , .ZN( u1_u13_u6_n94 ) );
  NOR2_X1 u1_u13_u6_U67 (.A2( u1_u13_X_37 ) , .A1( u1_u13_X_38 ) , .ZN( u1_u13_u6_n91 ) );
  NAND2_X1 u1_u13_u6_U68 (.A1( u1_u13_X_41 ) , .ZN( u1_u13_u6_n144 ) , .A2( u1_u13_u6_n157 ) );
  NAND2_X1 u1_u13_u6_U69 (.A2( u1_u13_X_40 ) , .A1( u1_u13_X_41 ) , .ZN( u1_u13_u6_n139 ) );
  NOR2_X1 u1_u13_u6_U7 (.A1( u1_u13_u6_n118 ) , .ZN( u1_u13_u6_n143 ) , .A2( u1_u13_u6_n168 ) );
  AND2_X1 u1_u13_u6_U70 (.A1( u1_u13_X_39 ) , .A2( u1_u13_u6_n156 ) , .ZN( u1_u13_u6_n96 ) );
  AND2_X1 u1_u13_u6_U71 (.A1( u1_u13_X_39 ) , .A2( u1_u13_X_42 ) , .ZN( u1_u13_u6_n99 ) );
  INV_X1 u1_u13_u6_U72 (.A( u1_u13_X_40 ) , .ZN( u1_u13_u6_n157 ) );
  INV_X1 u1_u13_u6_U73 (.A( u1_u13_X_37 ) , .ZN( u1_u13_u6_n165 ) );
  INV_X1 u1_u13_u6_U74 (.A( u1_u13_X_38 ) , .ZN( u1_u13_u6_n162 ) );
  INV_X1 u1_u13_u6_U75 (.A( u1_u13_X_42 ) , .ZN( u1_u13_u6_n156 ) );
  NAND4_X1 u1_u13_u6_U76 (.ZN( u1_out13_32 ) , .A4( u1_u13_u6_n103 ) , .A3( u1_u13_u6_n104 ) , .A2( u1_u13_u6_n105 ) , .A1( u1_u13_u6_n106 ) );
  AOI22_X1 u1_u13_u6_U77 (.ZN( u1_u13_u6_n105 ) , .A2( u1_u13_u6_n108 ) , .A1( u1_u13_u6_n118 ) , .B2( u1_u13_u6_n126 ) , .B1( u1_u13_u6_n171 ) );
  AOI22_X1 u1_u13_u6_U78 (.ZN( u1_u13_u6_n104 ) , .A1( u1_u13_u6_n111 ) , .B1( u1_u13_u6_n124 ) , .B2( u1_u13_u6_n151 ) , .A2( u1_u13_u6_n93 ) );
  NAND4_X1 u1_u13_u6_U79 (.ZN( u1_out13_12 ) , .A4( u1_u13_u6_n114 ) , .A3( u1_u13_u6_n115 ) , .A2( u1_u13_u6_n116 ) , .A1( u1_u13_u6_n117 ) );
  OAI21_X1 u1_u13_u6_U8 (.A( u1_u13_u6_n159 ) , .B1( u1_u13_u6_n169 ) , .B2( u1_u13_u6_n173 ) , .ZN( u1_u13_u6_n90 ) );
  OAI22_X1 u1_u13_u6_U80 (.B2( u1_u13_u6_n111 ) , .ZN( u1_u13_u6_n116 ) , .B1( u1_u13_u6_n126 ) , .A2( u1_u13_u6_n164 ) , .A1( u1_u13_u6_n167 ) );
  OAI21_X1 u1_u13_u6_U81 (.A( u1_u13_u6_n108 ) , .ZN( u1_u13_u6_n117 ) , .B2( u1_u13_u6_n141 ) , .B1( u1_u13_u6_n163 ) );
  OAI211_X1 u1_u13_u6_U82 (.ZN( u1_out13_7 ) , .B( u1_u13_u6_n153 ) , .C2( u1_u13_u6_n154 ) , .C1( u1_u13_u6_n155 ) , .A( u1_u13_u6_n174 ) );
  NOR3_X1 u1_u13_u6_U83 (.A1( u1_u13_u6_n141 ) , .ZN( u1_u13_u6_n154 ) , .A3( u1_u13_u6_n164 ) , .A2( u1_u13_u6_n171 ) );
  AOI211_X1 u1_u13_u6_U84 (.B( u1_u13_u6_n149 ) , .A( u1_u13_u6_n150 ) , .C2( u1_u13_u6_n151 ) , .C1( u1_u13_u6_n152 ) , .ZN( u1_u13_u6_n153 ) );
  OAI211_X1 u1_u13_u6_U85 (.ZN( u1_out13_22 ) , .B( u1_u13_u6_n137 ) , .A( u1_u13_u6_n138 ) , .C2( u1_u13_u6_n139 ) , .C1( u1_u13_u6_n140 ) );
  AOI22_X1 u1_u13_u6_U86 (.B1( u1_u13_u6_n124 ) , .A2( u1_u13_u6_n125 ) , .A1( u1_u13_u6_n126 ) , .ZN( u1_u13_u6_n138 ) , .B2( u1_u13_u6_n161 ) );
  AND4_X1 u1_u13_u6_U87 (.A3( u1_u13_u6_n119 ) , .A1( u1_u13_u6_n120 ) , .A4( u1_u13_u6_n129 ) , .ZN( u1_u13_u6_n140 ) , .A2( u1_u13_u6_n143 ) );
  NAND3_X1 u1_u13_u6_U88 (.A2( u1_u13_u6_n123 ) , .ZN( u1_u13_u6_n125 ) , .A1( u1_u13_u6_n130 ) , .A3( u1_u13_u6_n131 ) );
  NAND3_X1 u1_u13_u6_U89 (.A3( u1_u13_u6_n133 ) , .ZN( u1_u13_u6_n141 ) , .A1( u1_u13_u6_n145 ) , .A2( u1_u13_u6_n148 ) );
  INV_X1 u1_u13_u6_U9 (.ZN( u1_u13_u6_n172 ) , .A( u1_u13_u6_n88 ) );
  NAND3_X1 u1_u13_u6_U90 (.ZN( u1_u13_u6_n101 ) , .A3( u1_u13_u6_n107 ) , .A2( u1_u13_u6_n121 ) , .A1( u1_u13_u6_n127 ) );
  NAND3_X1 u1_u13_u6_U91 (.ZN( u1_u13_u6_n102 ) , .A3( u1_u13_u6_n130 ) , .A2( u1_u13_u6_n145 ) , .A1( u1_u13_u6_n166 ) );
  NAND3_X1 u1_u13_u6_U92 (.A3( u1_u13_u6_n113 ) , .A1( u1_u13_u6_n119 ) , .A2( u1_u13_u6_n123 ) , .ZN( u1_u13_u6_n93 ) );
  NAND3_X1 u1_u13_u6_U93 (.ZN( u1_u13_u6_n142 ) , .A2( u1_u13_u6_n172 ) , .A3( u1_u13_u6_n89 ) , .A1( u1_u13_u6_n90 ) );
  AND3_X1 u1_u13_u7_U10 (.A3( u1_u13_u7_n110 ) , .A2( u1_u13_u7_n127 ) , .A1( u1_u13_u7_n132 ) , .ZN( u1_u13_u7_n92 ) );
  OAI21_X1 u1_u13_u7_U11 (.A( u1_u13_u7_n161 ) , .B1( u1_u13_u7_n168 ) , .B2( u1_u13_u7_n173 ) , .ZN( u1_u13_u7_n91 ) );
  AOI211_X1 u1_u13_u7_U12 (.A( u1_u13_u7_n117 ) , .ZN( u1_u13_u7_n118 ) , .C2( u1_u13_u7_n126 ) , .C1( u1_u13_u7_n177 ) , .B( u1_u13_u7_n180 ) );
  OAI22_X1 u1_u13_u7_U13 (.B1( u1_u13_u7_n115 ) , .ZN( u1_u13_u7_n117 ) , .A2( u1_u13_u7_n133 ) , .A1( u1_u13_u7_n137 ) , .B2( u1_u13_u7_n162 ) );
  INV_X1 u1_u13_u7_U14 (.A( u1_u13_u7_n116 ) , .ZN( u1_u13_u7_n180 ) );
  NOR3_X1 u1_u13_u7_U15 (.ZN( u1_u13_u7_n115 ) , .A3( u1_u13_u7_n145 ) , .A2( u1_u13_u7_n168 ) , .A1( u1_u13_u7_n169 ) );
  OAI211_X1 u1_u13_u7_U16 (.B( u1_u13_u7_n122 ) , .A( u1_u13_u7_n123 ) , .C2( u1_u13_u7_n124 ) , .ZN( u1_u13_u7_n154 ) , .C1( u1_u13_u7_n162 ) );
  AOI222_X1 u1_u13_u7_U17 (.ZN( u1_u13_u7_n122 ) , .C2( u1_u13_u7_n126 ) , .C1( u1_u13_u7_n145 ) , .B1( u1_u13_u7_n161 ) , .A2( u1_u13_u7_n165 ) , .B2( u1_u13_u7_n170 ) , .A1( u1_u13_u7_n176 ) );
  INV_X1 u1_u13_u7_U18 (.A( u1_u13_u7_n133 ) , .ZN( u1_u13_u7_n176 ) );
  NOR3_X1 u1_u13_u7_U19 (.A2( u1_u13_u7_n134 ) , .A1( u1_u13_u7_n135 ) , .ZN( u1_u13_u7_n136 ) , .A3( u1_u13_u7_n171 ) );
  NOR2_X1 u1_u13_u7_U20 (.A1( u1_u13_u7_n130 ) , .A2( u1_u13_u7_n134 ) , .ZN( u1_u13_u7_n153 ) );
  INV_X1 u1_u13_u7_U21 (.A( u1_u13_u7_n101 ) , .ZN( u1_u13_u7_n165 ) );
  NOR2_X1 u1_u13_u7_U22 (.ZN( u1_u13_u7_n111 ) , .A2( u1_u13_u7_n134 ) , .A1( u1_u13_u7_n169 ) );
  AOI21_X1 u1_u13_u7_U23 (.ZN( u1_u13_u7_n104 ) , .B2( u1_u13_u7_n112 ) , .B1( u1_u13_u7_n127 ) , .A( u1_u13_u7_n164 ) );
  AOI21_X1 u1_u13_u7_U24 (.ZN( u1_u13_u7_n106 ) , .B1( u1_u13_u7_n133 ) , .B2( u1_u13_u7_n146 ) , .A( u1_u13_u7_n162 ) );
  AOI21_X1 u1_u13_u7_U25 (.A( u1_u13_u7_n101 ) , .ZN( u1_u13_u7_n107 ) , .B2( u1_u13_u7_n128 ) , .B1( u1_u13_u7_n175 ) );
  INV_X1 u1_u13_u7_U26 (.A( u1_u13_u7_n138 ) , .ZN( u1_u13_u7_n171 ) );
  INV_X1 u1_u13_u7_U27 (.A( u1_u13_u7_n131 ) , .ZN( u1_u13_u7_n177 ) );
  INV_X1 u1_u13_u7_U28 (.A( u1_u13_u7_n110 ) , .ZN( u1_u13_u7_n174 ) );
  NAND2_X1 u1_u13_u7_U29 (.A1( u1_u13_u7_n129 ) , .A2( u1_u13_u7_n132 ) , .ZN( u1_u13_u7_n149 ) );
  OAI21_X1 u1_u13_u7_U3 (.ZN( u1_u13_u7_n159 ) , .A( u1_u13_u7_n165 ) , .B2( u1_u13_u7_n171 ) , .B1( u1_u13_u7_n174 ) );
  NAND2_X1 u1_u13_u7_U30 (.A1( u1_u13_u7_n113 ) , .A2( u1_u13_u7_n124 ) , .ZN( u1_u13_u7_n130 ) );
  INV_X1 u1_u13_u7_U31 (.A( u1_u13_u7_n112 ) , .ZN( u1_u13_u7_n173 ) );
  INV_X1 u1_u13_u7_U32 (.A( u1_u13_u7_n128 ) , .ZN( u1_u13_u7_n168 ) );
  INV_X1 u1_u13_u7_U33 (.A( u1_u13_u7_n148 ) , .ZN( u1_u13_u7_n169 ) );
  INV_X1 u1_u13_u7_U34 (.A( u1_u13_u7_n127 ) , .ZN( u1_u13_u7_n179 ) );
  NOR2_X1 u1_u13_u7_U35 (.ZN( u1_u13_u7_n101 ) , .A2( u1_u13_u7_n150 ) , .A1( u1_u13_u7_n156 ) );
  AOI211_X1 u1_u13_u7_U36 (.B( u1_u13_u7_n154 ) , .A( u1_u13_u7_n155 ) , .C1( u1_u13_u7_n156 ) , .ZN( u1_u13_u7_n157 ) , .C2( u1_u13_u7_n172 ) );
  INV_X1 u1_u13_u7_U37 (.A( u1_u13_u7_n153 ) , .ZN( u1_u13_u7_n172 ) );
  AOI211_X1 u1_u13_u7_U38 (.B( u1_u13_u7_n139 ) , .A( u1_u13_u7_n140 ) , .C2( u1_u13_u7_n141 ) , .ZN( u1_u13_u7_n142 ) , .C1( u1_u13_u7_n156 ) );
  NAND4_X1 u1_u13_u7_U39 (.A3( u1_u13_u7_n127 ) , .A2( u1_u13_u7_n128 ) , .A1( u1_u13_u7_n129 ) , .ZN( u1_u13_u7_n141 ) , .A4( u1_u13_u7_n147 ) );
  INV_X1 u1_u13_u7_U4 (.A( u1_u13_u7_n111 ) , .ZN( u1_u13_u7_n170 ) );
  AOI21_X1 u1_u13_u7_U40 (.A( u1_u13_u7_n137 ) , .B1( u1_u13_u7_n138 ) , .ZN( u1_u13_u7_n139 ) , .B2( u1_u13_u7_n146 ) );
  OAI22_X1 u1_u13_u7_U41 (.B1( u1_u13_u7_n136 ) , .ZN( u1_u13_u7_n140 ) , .A1( u1_u13_u7_n153 ) , .B2( u1_u13_u7_n162 ) , .A2( u1_u13_u7_n164 ) );
  AOI21_X1 u1_u13_u7_U42 (.ZN( u1_u13_u7_n123 ) , .B1( u1_u13_u7_n165 ) , .B2( u1_u13_u7_n177 ) , .A( u1_u13_u7_n97 ) );
  AOI21_X1 u1_u13_u7_U43 (.B2( u1_u13_u7_n113 ) , .B1( u1_u13_u7_n124 ) , .A( u1_u13_u7_n125 ) , .ZN( u1_u13_u7_n97 ) );
  INV_X1 u1_u13_u7_U44 (.A( u1_u13_u7_n125 ) , .ZN( u1_u13_u7_n161 ) );
  INV_X1 u1_u13_u7_U45 (.A( u1_u13_u7_n152 ) , .ZN( u1_u13_u7_n162 ) );
  AOI22_X1 u1_u13_u7_U46 (.A2( u1_u13_u7_n114 ) , .ZN( u1_u13_u7_n119 ) , .B1( u1_u13_u7_n130 ) , .A1( u1_u13_u7_n156 ) , .B2( u1_u13_u7_n165 ) );
  NAND2_X1 u1_u13_u7_U47 (.A2( u1_u13_u7_n112 ) , .ZN( u1_u13_u7_n114 ) , .A1( u1_u13_u7_n175 ) );
  AND2_X1 u1_u13_u7_U48 (.ZN( u1_u13_u7_n145 ) , .A2( u1_u13_u7_n98 ) , .A1( u1_u13_u7_n99 ) );
  NOR2_X1 u1_u13_u7_U49 (.ZN( u1_u13_u7_n137 ) , .A1( u1_u13_u7_n150 ) , .A2( u1_u13_u7_n161 ) );
  INV_X1 u1_u13_u7_U5 (.A( u1_u13_u7_n149 ) , .ZN( u1_u13_u7_n175 ) );
  AOI21_X1 u1_u13_u7_U50 (.ZN( u1_u13_u7_n105 ) , .B2( u1_u13_u7_n110 ) , .A( u1_u13_u7_n125 ) , .B1( u1_u13_u7_n147 ) );
  NAND2_X1 u1_u13_u7_U51 (.ZN( u1_u13_u7_n146 ) , .A1( u1_u13_u7_n95 ) , .A2( u1_u13_u7_n98 ) );
  NAND2_X1 u1_u13_u7_U52 (.A2( u1_u13_u7_n103 ) , .ZN( u1_u13_u7_n147 ) , .A1( u1_u13_u7_n93 ) );
  NAND2_X1 u1_u13_u7_U53 (.A1( u1_u13_u7_n103 ) , .ZN( u1_u13_u7_n127 ) , .A2( u1_u13_u7_n99 ) );
  OR2_X1 u1_u13_u7_U54 (.ZN( u1_u13_u7_n126 ) , .A2( u1_u13_u7_n152 ) , .A1( u1_u13_u7_n156 ) );
  NAND2_X1 u1_u13_u7_U55 (.A2( u1_u13_u7_n102 ) , .A1( u1_u13_u7_n103 ) , .ZN( u1_u13_u7_n133 ) );
  NAND2_X1 u1_u13_u7_U56 (.ZN( u1_u13_u7_n112 ) , .A2( u1_u13_u7_n96 ) , .A1( u1_u13_u7_n99 ) );
  NAND2_X1 u1_u13_u7_U57 (.A2( u1_u13_u7_n102 ) , .ZN( u1_u13_u7_n128 ) , .A1( u1_u13_u7_n98 ) );
  NAND2_X1 u1_u13_u7_U58 (.A1( u1_u13_u7_n100 ) , .ZN( u1_u13_u7_n113 ) , .A2( u1_u13_u7_n93 ) );
  NAND2_X1 u1_u13_u7_U59 (.A2( u1_u13_u7_n102 ) , .ZN( u1_u13_u7_n124 ) , .A1( u1_u13_u7_n96 ) );
  INV_X1 u1_u13_u7_U6 (.A( u1_u13_u7_n154 ) , .ZN( u1_u13_u7_n178 ) );
  NAND2_X1 u1_u13_u7_U60 (.ZN( u1_u13_u7_n110 ) , .A1( u1_u13_u7_n95 ) , .A2( u1_u13_u7_n96 ) );
  INV_X1 u1_u13_u7_U61 (.A( u1_u13_u7_n150 ) , .ZN( u1_u13_u7_n164 ) );
  AND2_X1 u1_u13_u7_U62 (.ZN( u1_u13_u7_n134 ) , .A1( u1_u13_u7_n93 ) , .A2( u1_u13_u7_n98 ) );
  NAND2_X1 u1_u13_u7_U63 (.A1( u1_u13_u7_n100 ) , .A2( u1_u13_u7_n102 ) , .ZN( u1_u13_u7_n129 ) );
  NAND2_X1 u1_u13_u7_U64 (.A2( u1_u13_u7_n103 ) , .ZN( u1_u13_u7_n131 ) , .A1( u1_u13_u7_n95 ) );
  NAND2_X1 u1_u13_u7_U65 (.A1( u1_u13_u7_n100 ) , .ZN( u1_u13_u7_n138 ) , .A2( u1_u13_u7_n99 ) );
  NAND2_X1 u1_u13_u7_U66 (.ZN( u1_u13_u7_n132 ) , .A1( u1_u13_u7_n93 ) , .A2( u1_u13_u7_n96 ) );
  NAND2_X1 u1_u13_u7_U67 (.A1( u1_u13_u7_n100 ) , .ZN( u1_u13_u7_n148 ) , .A2( u1_u13_u7_n95 ) );
  NOR2_X1 u1_u13_u7_U68 (.A2( u1_u13_X_47 ) , .ZN( u1_u13_u7_n150 ) , .A1( u1_u13_u7_n163 ) );
  NOR2_X1 u1_u13_u7_U69 (.A2( u1_u13_X_43 ) , .A1( u1_u13_X_44 ) , .ZN( u1_u13_u7_n103 ) );
  AOI211_X1 u1_u13_u7_U7 (.ZN( u1_u13_u7_n116 ) , .A( u1_u13_u7_n155 ) , .C1( u1_u13_u7_n161 ) , .C2( u1_u13_u7_n171 ) , .B( u1_u13_u7_n94 ) );
  NOR2_X1 u1_u13_u7_U70 (.A2( u1_u13_X_48 ) , .A1( u1_u13_u7_n166 ) , .ZN( u1_u13_u7_n95 ) );
  NOR2_X1 u1_u13_u7_U71 (.A2( u1_u13_X_45 ) , .A1( u1_u13_X_48 ) , .ZN( u1_u13_u7_n99 ) );
  NOR2_X1 u1_u13_u7_U72 (.A2( u1_u13_X_44 ) , .A1( u1_u13_u7_n167 ) , .ZN( u1_u13_u7_n98 ) );
  NOR2_X1 u1_u13_u7_U73 (.A2( u1_u13_X_46 ) , .A1( u1_u13_X_47 ) , .ZN( u1_u13_u7_n152 ) );
  AND2_X1 u1_u13_u7_U74 (.A1( u1_u13_X_47 ) , .ZN( u1_u13_u7_n156 ) , .A2( u1_u13_u7_n163 ) );
  NAND2_X1 u1_u13_u7_U75 (.A2( u1_u13_X_46 ) , .A1( u1_u13_X_47 ) , .ZN( u1_u13_u7_n125 ) );
  AND2_X1 u1_u13_u7_U76 (.A2( u1_u13_X_45 ) , .A1( u1_u13_X_48 ) , .ZN( u1_u13_u7_n102 ) );
  AND2_X1 u1_u13_u7_U77 (.A2( u1_u13_X_43 ) , .A1( u1_u13_X_44 ) , .ZN( u1_u13_u7_n96 ) );
  AND2_X1 u1_u13_u7_U78 (.A1( u1_u13_X_44 ) , .ZN( u1_u13_u7_n100 ) , .A2( u1_u13_u7_n167 ) );
  AND2_X1 u1_u13_u7_U79 (.A1( u1_u13_X_48 ) , .A2( u1_u13_u7_n166 ) , .ZN( u1_u13_u7_n93 ) );
  OAI222_X1 u1_u13_u7_U8 (.C2( u1_u13_u7_n101 ) , .B2( u1_u13_u7_n111 ) , .A1( u1_u13_u7_n113 ) , .C1( u1_u13_u7_n146 ) , .A2( u1_u13_u7_n162 ) , .B1( u1_u13_u7_n164 ) , .ZN( u1_u13_u7_n94 ) );
  INV_X1 u1_u13_u7_U80 (.A( u1_u13_X_46 ) , .ZN( u1_u13_u7_n163 ) );
  INV_X1 u1_u13_u7_U81 (.A( u1_u13_X_43 ) , .ZN( u1_u13_u7_n167 ) );
  INV_X1 u1_u13_u7_U82 (.A( u1_u13_X_45 ) , .ZN( u1_u13_u7_n166 ) );
  NAND4_X1 u1_u13_u7_U83 (.ZN( u1_out13_5 ) , .A4( u1_u13_u7_n108 ) , .A3( u1_u13_u7_n109 ) , .A1( u1_u13_u7_n116 ) , .A2( u1_u13_u7_n123 ) );
  AOI22_X1 u1_u13_u7_U84 (.ZN( u1_u13_u7_n109 ) , .A2( u1_u13_u7_n126 ) , .B2( u1_u13_u7_n145 ) , .B1( u1_u13_u7_n156 ) , .A1( u1_u13_u7_n171 ) );
  NOR4_X1 u1_u13_u7_U85 (.A4( u1_u13_u7_n104 ) , .A3( u1_u13_u7_n105 ) , .A2( u1_u13_u7_n106 ) , .A1( u1_u13_u7_n107 ) , .ZN( u1_u13_u7_n108 ) );
  NAND4_X1 u1_u13_u7_U86 (.ZN( u1_out13_27 ) , .A4( u1_u13_u7_n118 ) , .A3( u1_u13_u7_n119 ) , .A2( u1_u13_u7_n120 ) , .A1( u1_u13_u7_n121 ) );
  OAI21_X1 u1_u13_u7_U87 (.ZN( u1_u13_u7_n121 ) , .B2( u1_u13_u7_n145 ) , .A( u1_u13_u7_n150 ) , .B1( u1_u13_u7_n174 ) );
  OAI21_X1 u1_u13_u7_U88 (.ZN( u1_u13_u7_n120 ) , .A( u1_u13_u7_n161 ) , .B2( u1_u13_u7_n170 ) , .B1( u1_u13_u7_n179 ) );
  NAND4_X1 u1_u13_u7_U89 (.ZN( u1_out13_21 ) , .A4( u1_u13_u7_n157 ) , .A3( u1_u13_u7_n158 ) , .A2( u1_u13_u7_n159 ) , .A1( u1_u13_u7_n160 ) );
  OAI221_X1 u1_u13_u7_U9 (.C1( u1_u13_u7_n101 ) , .C2( u1_u13_u7_n147 ) , .ZN( u1_u13_u7_n155 ) , .B2( u1_u13_u7_n162 ) , .A( u1_u13_u7_n91 ) , .B1( u1_u13_u7_n92 ) );
  OAI21_X1 u1_u13_u7_U90 (.B1( u1_u13_u7_n145 ) , .ZN( u1_u13_u7_n160 ) , .A( u1_u13_u7_n161 ) , .B2( u1_u13_u7_n177 ) );
  AOI22_X1 u1_u13_u7_U91 (.B2( u1_u13_u7_n149 ) , .B1( u1_u13_u7_n150 ) , .A2( u1_u13_u7_n151 ) , .A1( u1_u13_u7_n152 ) , .ZN( u1_u13_u7_n158 ) );
  NAND4_X1 u1_u13_u7_U92 (.ZN( u1_out13_15 ) , .A4( u1_u13_u7_n142 ) , .A3( u1_u13_u7_n143 ) , .A2( u1_u13_u7_n144 ) , .A1( u1_u13_u7_n178 ) );
  OR2_X1 u1_u13_u7_U93 (.A2( u1_u13_u7_n125 ) , .A1( u1_u13_u7_n129 ) , .ZN( u1_u13_u7_n144 ) );
  AOI22_X1 u1_u13_u7_U94 (.A2( u1_u13_u7_n126 ) , .ZN( u1_u13_u7_n143 ) , .B2( u1_u13_u7_n165 ) , .B1( u1_u13_u7_n173 ) , .A1( u1_u13_u7_n174 ) );
  NAND3_X1 u1_u13_u7_U95 (.A3( u1_u13_u7_n146 ) , .A2( u1_u13_u7_n147 ) , .A1( u1_u13_u7_n148 ) , .ZN( u1_u13_u7_n151 ) );
  NAND3_X1 u1_u13_u7_U96 (.A3( u1_u13_u7_n131 ) , .A2( u1_u13_u7_n132 ) , .A1( u1_u13_u7_n133 ) , .ZN( u1_u13_u7_n135 ) );
  XOR2_X1 u1_u6_U26 (.B( u1_K7_30 ) , .A( u1_R5_21 ) , .Z( u1_u6_X_30 ) );
  XOR2_X1 u1_u6_U28 (.B( u1_K7_29 ) , .A( u1_R5_20 ) , .Z( u1_u6_X_29 ) );
  XOR2_X1 u1_u6_U29 (.B( u1_K7_28 ) , .A( u1_R5_19 ) , .Z( u1_u6_X_28 ) );
  XOR2_X1 u1_u6_U30 (.B( u1_K7_27 ) , .A( u1_R5_18 ) , .Z( u1_u6_X_27 ) );
  XOR2_X1 u1_u6_U31 (.B( u1_K7_26 ) , .A( u1_R5_17 ) , .Z( u1_u6_X_26 ) );
  XOR2_X1 u1_u6_U32 (.B( u1_K7_25 ) , .A( u1_R5_16 ) , .Z( u1_u6_X_25 ) );
  OAI22_X1 u1_u6_u4_U10 (.B2( u1_u6_u4_n135 ) , .ZN( u1_u6_u4_n137 ) , .B1( u1_u6_u4_n153 ) , .A1( u1_u6_u4_n155 ) , .A2( u1_u6_u4_n171 ) );
  AND3_X1 u1_u6_u4_U11 (.A2( u1_u6_u4_n134 ) , .ZN( u1_u6_u4_n135 ) , .A3( u1_u6_u4_n145 ) , .A1( u1_u6_u4_n157 ) );
  NAND2_X1 u1_u6_u4_U12 (.ZN( u1_u6_u4_n132 ) , .A2( u1_u6_u4_n170 ) , .A1( u1_u6_u4_n173 ) );
  AOI21_X1 u1_u6_u4_U13 (.B2( u1_u6_u4_n160 ) , .B1( u1_u6_u4_n161 ) , .ZN( u1_u6_u4_n162 ) , .A( u1_u6_u4_n170 ) );
  AOI21_X1 u1_u6_u4_U14 (.ZN( u1_u6_u4_n107 ) , .B2( u1_u6_u4_n143 ) , .A( u1_u6_u4_n174 ) , .B1( u1_u6_u4_n184 ) );
  AOI21_X1 u1_u6_u4_U15 (.B2( u1_u6_u4_n158 ) , .B1( u1_u6_u4_n159 ) , .ZN( u1_u6_u4_n163 ) , .A( u1_u6_u4_n174 ) );
  AOI21_X1 u1_u6_u4_U16 (.A( u1_u6_u4_n153 ) , .B2( u1_u6_u4_n154 ) , .B1( u1_u6_u4_n155 ) , .ZN( u1_u6_u4_n165 ) );
  AOI21_X1 u1_u6_u4_U17 (.A( u1_u6_u4_n156 ) , .B2( u1_u6_u4_n157 ) , .ZN( u1_u6_u4_n164 ) , .B1( u1_u6_u4_n184 ) );
  INV_X1 u1_u6_u4_U18 (.A( u1_u6_u4_n138 ) , .ZN( u1_u6_u4_n170 ) );
  AND2_X1 u1_u6_u4_U19 (.A2( u1_u6_u4_n120 ) , .ZN( u1_u6_u4_n155 ) , .A1( u1_u6_u4_n160 ) );
  INV_X1 u1_u6_u4_U20 (.A( u1_u6_u4_n156 ) , .ZN( u1_u6_u4_n175 ) );
  NAND2_X1 u1_u6_u4_U21 (.A2( u1_u6_u4_n118 ) , .ZN( u1_u6_u4_n131 ) , .A1( u1_u6_u4_n147 ) );
  NAND2_X1 u1_u6_u4_U22 (.A1( u1_u6_u4_n119 ) , .A2( u1_u6_u4_n120 ) , .ZN( u1_u6_u4_n130 ) );
  NAND2_X1 u1_u6_u4_U23 (.ZN( u1_u6_u4_n117 ) , .A2( u1_u6_u4_n118 ) , .A1( u1_u6_u4_n148 ) );
  NAND2_X1 u1_u6_u4_U24 (.ZN( u1_u6_u4_n129 ) , .A1( u1_u6_u4_n134 ) , .A2( u1_u6_u4_n148 ) );
  AND3_X1 u1_u6_u4_U25 (.A1( u1_u6_u4_n119 ) , .A2( u1_u6_u4_n143 ) , .A3( u1_u6_u4_n154 ) , .ZN( u1_u6_u4_n161 ) );
  AND2_X1 u1_u6_u4_U26 (.A1( u1_u6_u4_n145 ) , .A2( u1_u6_u4_n147 ) , .ZN( u1_u6_u4_n159 ) );
  OR3_X1 u1_u6_u4_U27 (.A3( u1_u6_u4_n114 ) , .A2( u1_u6_u4_n115 ) , .A1( u1_u6_u4_n116 ) , .ZN( u1_u6_u4_n136 ) );
  AOI21_X1 u1_u6_u4_U28 (.A( u1_u6_u4_n113 ) , .ZN( u1_u6_u4_n116 ) , .B2( u1_u6_u4_n173 ) , .B1( u1_u6_u4_n174 ) );
  AOI21_X1 u1_u6_u4_U29 (.ZN( u1_u6_u4_n115 ) , .B2( u1_u6_u4_n145 ) , .B1( u1_u6_u4_n146 ) , .A( u1_u6_u4_n156 ) );
  NOR2_X1 u1_u6_u4_U3 (.ZN( u1_u6_u4_n121 ) , .A1( u1_u6_u4_n181 ) , .A2( u1_u6_u4_n182 ) );
  OAI22_X1 u1_u6_u4_U30 (.ZN( u1_u6_u4_n114 ) , .A2( u1_u6_u4_n121 ) , .B1( u1_u6_u4_n160 ) , .B2( u1_u6_u4_n170 ) , .A1( u1_u6_u4_n171 ) );
  INV_X1 u1_u6_u4_U31 (.A( u1_u6_u4_n158 ) , .ZN( u1_u6_u4_n182 ) );
  INV_X1 u1_u6_u4_U32 (.ZN( u1_u6_u4_n181 ) , .A( u1_u6_u4_n96 ) );
  INV_X1 u1_u6_u4_U33 (.A( u1_u6_u4_n144 ) , .ZN( u1_u6_u4_n179 ) );
  INV_X1 u1_u6_u4_U34 (.A( u1_u6_u4_n157 ) , .ZN( u1_u6_u4_n178 ) );
  NAND2_X1 u1_u6_u4_U35 (.A2( u1_u6_u4_n154 ) , .A1( u1_u6_u4_n96 ) , .ZN( u1_u6_u4_n97 ) );
  INV_X1 u1_u6_u4_U36 (.ZN( u1_u6_u4_n186 ) , .A( u1_u6_u4_n95 ) );
  OAI221_X1 u1_u6_u4_U37 (.C1( u1_u6_u4_n134 ) , .B1( u1_u6_u4_n158 ) , .B2( u1_u6_u4_n171 ) , .C2( u1_u6_u4_n173 ) , .A( u1_u6_u4_n94 ) , .ZN( u1_u6_u4_n95 ) );
  AOI222_X1 u1_u6_u4_U38 (.B2( u1_u6_u4_n132 ) , .A1( u1_u6_u4_n138 ) , .C2( u1_u6_u4_n175 ) , .A2( u1_u6_u4_n179 ) , .C1( u1_u6_u4_n181 ) , .B1( u1_u6_u4_n185 ) , .ZN( u1_u6_u4_n94 ) );
  INV_X1 u1_u6_u4_U39 (.A( u1_u6_u4_n113 ) , .ZN( u1_u6_u4_n185 ) );
  INV_X1 u1_u6_u4_U4 (.A( u1_u6_u4_n117 ) , .ZN( u1_u6_u4_n184 ) );
  INV_X1 u1_u6_u4_U40 (.A( u1_u6_u4_n143 ) , .ZN( u1_u6_u4_n183 ) );
  NOR2_X1 u1_u6_u4_U41 (.ZN( u1_u6_u4_n138 ) , .A1( u1_u6_u4_n168 ) , .A2( u1_u6_u4_n169 ) );
  NOR2_X1 u1_u6_u4_U42 (.A1( u1_u6_u4_n150 ) , .A2( u1_u6_u4_n152 ) , .ZN( u1_u6_u4_n153 ) );
  NOR2_X1 u1_u6_u4_U43 (.A2( u1_u6_u4_n128 ) , .A1( u1_u6_u4_n138 ) , .ZN( u1_u6_u4_n156 ) );
  AOI22_X1 u1_u6_u4_U44 (.B2( u1_u6_u4_n122 ) , .A1( u1_u6_u4_n123 ) , .ZN( u1_u6_u4_n124 ) , .B1( u1_u6_u4_n128 ) , .A2( u1_u6_u4_n172 ) );
  INV_X1 u1_u6_u4_U45 (.A( u1_u6_u4_n153 ) , .ZN( u1_u6_u4_n172 ) );
  NAND2_X1 u1_u6_u4_U46 (.A2( u1_u6_u4_n120 ) , .ZN( u1_u6_u4_n123 ) , .A1( u1_u6_u4_n161 ) );
  AOI22_X1 u1_u6_u4_U47 (.B2( u1_u6_u4_n132 ) , .A2( u1_u6_u4_n133 ) , .ZN( u1_u6_u4_n140 ) , .A1( u1_u6_u4_n150 ) , .B1( u1_u6_u4_n179 ) );
  NAND2_X1 u1_u6_u4_U48 (.ZN( u1_u6_u4_n133 ) , .A2( u1_u6_u4_n146 ) , .A1( u1_u6_u4_n154 ) );
  NAND2_X1 u1_u6_u4_U49 (.A1( u1_u6_u4_n103 ) , .ZN( u1_u6_u4_n154 ) , .A2( u1_u6_u4_n98 ) );
  NOR4_X1 u1_u6_u4_U5 (.A4( u1_u6_u4_n106 ) , .A3( u1_u6_u4_n107 ) , .A2( u1_u6_u4_n108 ) , .A1( u1_u6_u4_n109 ) , .ZN( u1_u6_u4_n110 ) );
  NAND2_X1 u1_u6_u4_U50 (.A1( u1_u6_u4_n101 ) , .ZN( u1_u6_u4_n158 ) , .A2( u1_u6_u4_n99 ) );
  AOI21_X1 u1_u6_u4_U51 (.ZN( u1_u6_u4_n127 ) , .A( u1_u6_u4_n136 ) , .B2( u1_u6_u4_n150 ) , .B1( u1_u6_u4_n180 ) );
  INV_X1 u1_u6_u4_U52 (.A( u1_u6_u4_n160 ) , .ZN( u1_u6_u4_n180 ) );
  NAND2_X1 u1_u6_u4_U53 (.A2( u1_u6_u4_n104 ) , .A1( u1_u6_u4_n105 ) , .ZN( u1_u6_u4_n146 ) );
  NAND2_X1 u1_u6_u4_U54 (.A2( u1_u6_u4_n101 ) , .A1( u1_u6_u4_n102 ) , .ZN( u1_u6_u4_n160 ) );
  NAND2_X1 u1_u6_u4_U55 (.ZN( u1_u6_u4_n134 ) , .A1( u1_u6_u4_n98 ) , .A2( u1_u6_u4_n99 ) );
  NAND2_X1 u1_u6_u4_U56 (.A1( u1_u6_u4_n103 ) , .A2( u1_u6_u4_n104 ) , .ZN( u1_u6_u4_n143 ) );
  NAND2_X1 u1_u6_u4_U57 (.A2( u1_u6_u4_n105 ) , .ZN( u1_u6_u4_n145 ) , .A1( u1_u6_u4_n98 ) );
  NAND2_X1 u1_u6_u4_U58 (.A1( u1_u6_u4_n100 ) , .A2( u1_u6_u4_n105 ) , .ZN( u1_u6_u4_n120 ) );
  NAND2_X1 u1_u6_u4_U59 (.A1( u1_u6_u4_n102 ) , .A2( u1_u6_u4_n104 ) , .ZN( u1_u6_u4_n148 ) );
  AOI21_X1 u1_u6_u4_U6 (.ZN( u1_u6_u4_n106 ) , .B2( u1_u6_u4_n146 ) , .B1( u1_u6_u4_n158 ) , .A( u1_u6_u4_n170 ) );
  NAND2_X1 u1_u6_u4_U60 (.A2( u1_u6_u4_n100 ) , .A1( u1_u6_u4_n103 ) , .ZN( u1_u6_u4_n157 ) );
  INV_X1 u1_u6_u4_U61 (.A( u1_u6_u4_n150 ) , .ZN( u1_u6_u4_n173 ) );
  INV_X1 u1_u6_u4_U62 (.A( u1_u6_u4_n152 ) , .ZN( u1_u6_u4_n171 ) );
  NAND2_X1 u1_u6_u4_U63 (.A1( u1_u6_u4_n100 ) , .ZN( u1_u6_u4_n118 ) , .A2( u1_u6_u4_n99 ) );
  NAND2_X1 u1_u6_u4_U64 (.A2( u1_u6_u4_n100 ) , .A1( u1_u6_u4_n102 ) , .ZN( u1_u6_u4_n144 ) );
  NAND2_X1 u1_u6_u4_U65 (.A2( u1_u6_u4_n101 ) , .A1( u1_u6_u4_n105 ) , .ZN( u1_u6_u4_n96 ) );
  INV_X1 u1_u6_u4_U66 (.A( u1_u6_u4_n128 ) , .ZN( u1_u6_u4_n174 ) );
  NAND2_X1 u1_u6_u4_U67 (.A2( u1_u6_u4_n102 ) , .ZN( u1_u6_u4_n119 ) , .A1( u1_u6_u4_n98 ) );
  NAND2_X1 u1_u6_u4_U68 (.A2( u1_u6_u4_n101 ) , .A1( u1_u6_u4_n103 ) , .ZN( u1_u6_u4_n147 ) );
  NAND2_X1 u1_u6_u4_U69 (.A2( u1_u6_u4_n104 ) , .ZN( u1_u6_u4_n113 ) , .A1( u1_u6_u4_n99 ) );
  AOI21_X1 u1_u6_u4_U7 (.ZN( u1_u6_u4_n108 ) , .B2( u1_u6_u4_n134 ) , .B1( u1_u6_u4_n155 ) , .A( u1_u6_u4_n156 ) );
  NOR2_X1 u1_u6_u4_U70 (.A2( u1_u6_X_28 ) , .ZN( u1_u6_u4_n150 ) , .A1( u1_u6_u4_n168 ) );
  NOR2_X1 u1_u6_u4_U71 (.A2( u1_u6_X_29 ) , .ZN( u1_u6_u4_n152 ) , .A1( u1_u6_u4_n169 ) );
  NOR2_X1 u1_u6_u4_U72 (.A2( u1_u6_X_30 ) , .ZN( u1_u6_u4_n105 ) , .A1( u1_u6_u4_n176 ) );
  NOR2_X1 u1_u6_u4_U73 (.A2( u1_u6_X_26 ) , .ZN( u1_u6_u4_n100 ) , .A1( u1_u6_u4_n177 ) );
  NOR2_X1 u1_u6_u4_U74 (.A2( u1_u6_X_28 ) , .A1( u1_u6_X_29 ) , .ZN( u1_u6_u4_n128 ) );
  NOR2_X1 u1_u6_u4_U75 (.A2( u1_u6_X_27 ) , .A1( u1_u6_X_30 ) , .ZN( u1_u6_u4_n102 ) );
  NOR2_X1 u1_u6_u4_U76 (.A2( u1_u6_X_25 ) , .A1( u1_u6_X_26 ) , .ZN( u1_u6_u4_n98 ) );
  AND2_X1 u1_u6_u4_U77 (.A2( u1_u6_X_25 ) , .A1( u1_u6_X_26 ) , .ZN( u1_u6_u4_n104 ) );
  AND2_X1 u1_u6_u4_U78 (.A1( u1_u6_X_30 ) , .A2( u1_u6_u4_n176 ) , .ZN( u1_u6_u4_n99 ) );
  AND2_X1 u1_u6_u4_U79 (.A1( u1_u6_X_26 ) , .ZN( u1_u6_u4_n101 ) , .A2( u1_u6_u4_n177 ) );
  AOI21_X1 u1_u6_u4_U8 (.ZN( u1_u6_u4_n109 ) , .A( u1_u6_u4_n153 ) , .B1( u1_u6_u4_n159 ) , .B2( u1_u6_u4_n184 ) );
  AND2_X1 u1_u6_u4_U80 (.A1( u1_u6_X_27 ) , .A2( u1_u6_X_30 ) , .ZN( u1_u6_u4_n103 ) );
  INV_X1 u1_u6_u4_U81 (.A( u1_u6_X_28 ) , .ZN( u1_u6_u4_n169 ) );
  INV_X1 u1_u6_u4_U82 (.A( u1_u6_X_29 ) , .ZN( u1_u6_u4_n168 ) );
  INV_X1 u1_u6_u4_U83 (.A( u1_u6_X_25 ) , .ZN( u1_u6_u4_n177 ) );
  INV_X1 u1_u6_u4_U84 (.A( u1_u6_X_27 ) , .ZN( u1_u6_u4_n176 ) );
  NAND4_X1 u1_u6_u4_U85 (.ZN( u1_out6_8 ) , .A4( u1_u6_u4_n110 ) , .A3( u1_u6_u4_n111 ) , .A2( u1_u6_u4_n112 ) , .A1( u1_u6_u4_n186 ) );
  NAND2_X1 u1_u6_u4_U86 (.ZN( u1_u6_u4_n112 ) , .A2( u1_u6_u4_n130 ) , .A1( u1_u6_u4_n150 ) );
  AOI22_X1 u1_u6_u4_U87 (.ZN( u1_u6_u4_n111 ) , .B2( u1_u6_u4_n132 ) , .A1( u1_u6_u4_n152 ) , .B1( u1_u6_u4_n178 ) , .A2( u1_u6_u4_n97 ) );
  NAND4_X1 u1_u6_u4_U88 (.ZN( u1_out6_25 ) , .A4( u1_u6_u4_n139 ) , .A3( u1_u6_u4_n140 ) , .A2( u1_u6_u4_n141 ) , .A1( u1_u6_u4_n142 ) );
  OAI21_X1 u1_u6_u4_U89 (.B2( u1_u6_u4_n131 ) , .ZN( u1_u6_u4_n141 ) , .A( u1_u6_u4_n175 ) , .B1( u1_u6_u4_n183 ) );
  AOI211_X1 u1_u6_u4_U9 (.B( u1_u6_u4_n136 ) , .A( u1_u6_u4_n137 ) , .C2( u1_u6_u4_n138 ) , .ZN( u1_u6_u4_n139 ) , .C1( u1_u6_u4_n182 ) );
  OAI21_X1 u1_u6_u4_U90 (.A( u1_u6_u4_n128 ) , .B2( u1_u6_u4_n129 ) , .B1( u1_u6_u4_n130 ) , .ZN( u1_u6_u4_n142 ) );
  NAND4_X1 u1_u6_u4_U91 (.ZN( u1_out6_14 ) , .A4( u1_u6_u4_n124 ) , .A3( u1_u6_u4_n125 ) , .A2( u1_u6_u4_n126 ) , .A1( u1_u6_u4_n127 ) );
  AOI22_X1 u1_u6_u4_U92 (.B2( u1_u6_u4_n117 ) , .ZN( u1_u6_u4_n126 ) , .A1( u1_u6_u4_n129 ) , .B1( u1_u6_u4_n152 ) , .A2( u1_u6_u4_n175 ) );
  AOI22_X1 u1_u6_u4_U93 (.ZN( u1_u6_u4_n125 ) , .B2( u1_u6_u4_n131 ) , .A2( u1_u6_u4_n132 ) , .B1( u1_u6_u4_n138 ) , .A1( u1_u6_u4_n178 ) );
  AOI22_X1 u1_u6_u4_U94 (.B2( u1_u6_u4_n149 ) , .B1( u1_u6_u4_n150 ) , .A2( u1_u6_u4_n151 ) , .A1( u1_u6_u4_n152 ) , .ZN( u1_u6_u4_n167 ) );
  NOR4_X1 u1_u6_u4_U95 (.A4( u1_u6_u4_n162 ) , .A3( u1_u6_u4_n163 ) , .A2( u1_u6_u4_n164 ) , .A1( u1_u6_u4_n165 ) , .ZN( u1_u6_u4_n166 ) );
  NAND3_X1 u1_u6_u4_U96 (.ZN( u1_out6_3 ) , .A3( u1_u6_u4_n166 ) , .A1( u1_u6_u4_n167 ) , .A2( u1_u6_u4_n186 ) );
  NAND3_X1 u1_u6_u4_U97 (.A3( u1_u6_u4_n146 ) , .A2( u1_u6_u4_n147 ) , .A1( u1_u6_u4_n148 ) , .ZN( u1_u6_u4_n149 ) );
  NAND3_X1 u1_u6_u4_U98 (.A3( u1_u6_u4_n143 ) , .A2( u1_u6_u4_n144 ) , .A1( u1_u6_u4_n145 ) , .ZN( u1_u6_u4_n151 ) );
  NAND3_X1 u1_u6_u4_U99 (.A3( u1_u6_u4_n121 ) , .ZN( u1_u6_u4_n122 ) , .A2( u1_u6_u4_n144 ) , .A1( u1_u6_u4_n154 ) );
  XOR2_X1 u1_u7_U13 (.B( u1_K8_42 ) , .A( u1_R6_29 ) , .Z( u1_u7_X_42 ) );
  XOR2_X1 u1_u7_U14 (.B( u1_K8_41 ) , .A( u1_R6_28 ) , .Z( u1_u7_X_41 ) );
  XOR2_X1 u1_u7_U15 (.B( u1_K8_40 ) , .A( u1_R6_27 ) , .Z( u1_u7_X_40 ) );
  XOR2_X1 u1_u7_U17 (.B( u1_K8_39 ) , .A( u1_R6_26 ) , .Z( u1_u7_X_39 ) );
  XOR2_X1 u1_u7_U18 (.B( u1_K8_38 ) , .A( u1_R6_25 ) , .Z( u1_u7_X_38 ) );
  XOR2_X1 u1_u7_U19 (.B( u1_K8_37 ) , .A( u1_R6_24 ) , .Z( u1_u7_X_37 ) );
  INV_X1 u1_u7_u6_U10 (.ZN( u1_u7_u6_n172 ) , .A( u1_u7_u6_n88 ) );
  OAI21_X1 u1_u7_u6_U11 (.A( u1_u7_u6_n159 ) , .B1( u1_u7_u6_n169 ) , .B2( u1_u7_u6_n173 ) , .ZN( u1_u7_u6_n90 ) );
  AOI22_X1 u1_u7_u6_U12 (.A2( u1_u7_u6_n151 ) , .B2( u1_u7_u6_n161 ) , .A1( u1_u7_u6_n167 ) , .B1( u1_u7_u6_n170 ) , .ZN( u1_u7_u6_n89 ) );
  AOI21_X1 u1_u7_u6_U13 (.ZN( u1_u7_u6_n106 ) , .A( u1_u7_u6_n142 ) , .B2( u1_u7_u6_n159 ) , .B1( u1_u7_u6_n164 ) );
  INV_X1 u1_u7_u6_U14 (.A( u1_u7_u6_n155 ) , .ZN( u1_u7_u6_n161 ) );
  INV_X1 u1_u7_u6_U15 (.A( u1_u7_u6_n128 ) , .ZN( u1_u7_u6_n164 ) );
  NAND2_X1 u1_u7_u6_U16 (.ZN( u1_u7_u6_n110 ) , .A1( u1_u7_u6_n122 ) , .A2( u1_u7_u6_n129 ) );
  NAND2_X1 u1_u7_u6_U17 (.ZN( u1_u7_u6_n124 ) , .A2( u1_u7_u6_n146 ) , .A1( u1_u7_u6_n148 ) );
  INV_X1 u1_u7_u6_U18 (.A( u1_u7_u6_n132 ) , .ZN( u1_u7_u6_n171 ) );
  AND2_X1 u1_u7_u6_U19 (.A1( u1_u7_u6_n100 ) , .ZN( u1_u7_u6_n130 ) , .A2( u1_u7_u6_n147 ) );
  INV_X1 u1_u7_u6_U20 (.A( u1_u7_u6_n127 ) , .ZN( u1_u7_u6_n173 ) );
  INV_X1 u1_u7_u6_U21 (.A( u1_u7_u6_n121 ) , .ZN( u1_u7_u6_n167 ) );
  INV_X1 u1_u7_u6_U22 (.A( u1_u7_u6_n100 ) , .ZN( u1_u7_u6_n169 ) );
  INV_X1 u1_u7_u6_U23 (.A( u1_u7_u6_n123 ) , .ZN( u1_u7_u6_n170 ) );
  INV_X1 u1_u7_u6_U24 (.A( u1_u7_u6_n113 ) , .ZN( u1_u7_u6_n168 ) );
  AND2_X1 u1_u7_u6_U25 (.A1( u1_u7_u6_n107 ) , .A2( u1_u7_u6_n119 ) , .ZN( u1_u7_u6_n133 ) );
  AND2_X1 u1_u7_u6_U26 (.A2( u1_u7_u6_n121 ) , .A1( u1_u7_u6_n122 ) , .ZN( u1_u7_u6_n131 ) );
  AND3_X1 u1_u7_u6_U27 (.ZN( u1_u7_u6_n120 ) , .A2( u1_u7_u6_n127 ) , .A1( u1_u7_u6_n132 ) , .A3( u1_u7_u6_n145 ) );
  INV_X1 u1_u7_u6_U28 (.A( u1_u7_u6_n146 ) , .ZN( u1_u7_u6_n163 ) );
  AOI222_X1 u1_u7_u6_U29 (.ZN( u1_u7_u6_n114 ) , .A1( u1_u7_u6_n118 ) , .A2( u1_u7_u6_n126 ) , .B2( u1_u7_u6_n151 ) , .C2( u1_u7_u6_n159 ) , .C1( u1_u7_u6_n168 ) , .B1( u1_u7_u6_n169 ) );
  INV_X1 u1_u7_u6_U3 (.A( u1_u7_u6_n110 ) , .ZN( u1_u7_u6_n166 ) );
  NOR2_X1 u1_u7_u6_U30 (.A1( u1_u7_u6_n162 ) , .A2( u1_u7_u6_n165 ) , .ZN( u1_u7_u6_n98 ) );
  NAND2_X1 u1_u7_u6_U31 (.A1( u1_u7_u6_n144 ) , .ZN( u1_u7_u6_n151 ) , .A2( u1_u7_u6_n158 ) );
  NAND2_X1 u1_u7_u6_U32 (.ZN( u1_u7_u6_n132 ) , .A1( u1_u7_u6_n91 ) , .A2( u1_u7_u6_n97 ) );
  AOI22_X1 u1_u7_u6_U33 (.B2( u1_u7_u6_n110 ) , .B1( u1_u7_u6_n111 ) , .A1( u1_u7_u6_n112 ) , .ZN( u1_u7_u6_n115 ) , .A2( u1_u7_u6_n161 ) );
  NAND4_X1 u1_u7_u6_U34 (.A3( u1_u7_u6_n109 ) , .ZN( u1_u7_u6_n112 ) , .A4( u1_u7_u6_n132 ) , .A2( u1_u7_u6_n147 ) , .A1( u1_u7_u6_n166 ) );
  NOR2_X1 u1_u7_u6_U35 (.ZN( u1_u7_u6_n109 ) , .A1( u1_u7_u6_n170 ) , .A2( u1_u7_u6_n173 ) );
  NOR2_X1 u1_u7_u6_U36 (.A2( u1_u7_u6_n126 ) , .ZN( u1_u7_u6_n155 ) , .A1( u1_u7_u6_n160 ) );
  NAND2_X1 u1_u7_u6_U37 (.ZN( u1_u7_u6_n146 ) , .A2( u1_u7_u6_n94 ) , .A1( u1_u7_u6_n99 ) );
  AOI21_X1 u1_u7_u6_U38 (.A( u1_u7_u6_n144 ) , .B2( u1_u7_u6_n145 ) , .B1( u1_u7_u6_n146 ) , .ZN( u1_u7_u6_n150 ) );
  AOI211_X1 u1_u7_u6_U39 (.B( u1_u7_u6_n134 ) , .A( u1_u7_u6_n135 ) , .C1( u1_u7_u6_n136 ) , .ZN( u1_u7_u6_n137 ) , .C2( u1_u7_u6_n151 ) );
  INV_X1 u1_u7_u6_U4 (.A( u1_u7_u6_n142 ) , .ZN( u1_u7_u6_n174 ) );
  NAND4_X1 u1_u7_u6_U40 (.A4( u1_u7_u6_n127 ) , .A3( u1_u7_u6_n128 ) , .A2( u1_u7_u6_n129 ) , .A1( u1_u7_u6_n130 ) , .ZN( u1_u7_u6_n136 ) );
  AOI21_X1 u1_u7_u6_U41 (.B2( u1_u7_u6_n132 ) , .B1( u1_u7_u6_n133 ) , .ZN( u1_u7_u6_n134 ) , .A( u1_u7_u6_n158 ) );
  AOI21_X1 u1_u7_u6_U42 (.B1( u1_u7_u6_n131 ) , .ZN( u1_u7_u6_n135 ) , .A( u1_u7_u6_n144 ) , .B2( u1_u7_u6_n146 ) );
  INV_X1 u1_u7_u6_U43 (.A( u1_u7_u6_n111 ) , .ZN( u1_u7_u6_n158 ) );
  NAND2_X1 u1_u7_u6_U44 (.ZN( u1_u7_u6_n127 ) , .A1( u1_u7_u6_n91 ) , .A2( u1_u7_u6_n92 ) );
  NAND2_X1 u1_u7_u6_U45 (.ZN( u1_u7_u6_n129 ) , .A2( u1_u7_u6_n95 ) , .A1( u1_u7_u6_n96 ) );
  INV_X1 u1_u7_u6_U46 (.A( u1_u7_u6_n144 ) , .ZN( u1_u7_u6_n159 ) );
  NAND2_X1 u1_u7_u6_U47 (.ZN( u1_u7_u6_n145 ) , .A2( u1_u7_u6_n97 ) , .A1( u1_u7_u6_n98 ) );
  NAND2_X1 u1_u7_u6_U48 (.ZN( u1_u7_u6_n148 ) , .A2( u1_u7_u6_n92 ) , .A1( u1_u7_u6_n94 ) );
  NAND2_X1 u1_u7_u6_U49 (.ZN( u1_u7_u6_n108 ) , .A2( u1_u7_u6_n139 ) , .A1( u1_u7_u6_n144 ) );
  NAND2_X1 u1_u7_u6_U5 (.A2( u1_u7_u6_n143 ) , .ZN( u1_u7_u6_n152 ) , .A1( u1_u7_u6_n166 ) );
  NAND2_X1 u1_u7_u6_U50 (.ZN( u1_u7_u6_n121 ) , .A2( u1_u7_u6_n95 ) , .A1( u1_u7_u6_n97 ) );
  NAND2_X1 u1_u7_u6_U51 (.ZN( u1_u7_u6_n107 ) , .A2( u1_u7_u6_n92 ) , .A1( u1_u7_u6_n95 ) );
  AND2_X1 u1_u7_u6_U52 (.ZN( u1_u7_u6_n118 ) , .A2( u1_u7_u6_n91 ) , .A1( u1_u7_u6_n99 ) );
  NAND2_X1 u1_u7_u6_U53 (.ZN( u1_u7_u6_n147 ) , .A2( u1_u7_u6_n98 ) , .A1( u1_u7_u6_n99 ) );
  NAND2_X1 u1_u7_u6_U54 (.ZN( u1_u7_u6_n128 ) , .A1( u1_u7_u6_n94 ) , .A2( u1_u7_u6_n96 ) );
  NAND2_X1 u1_u7_u6_U55 (.ZN( u1_u7_u6_n119 ) , .A2( u1_u7_u6_n95 ) , .A1( u1_u7_u6_n99 ) );
  NAND2_X1 u1_u7_u6_U56 (.ZN( u1_u7_u6_n123 ) , .A2( u1_u7_u6_n91 ) , .A1( u1_u7_u6_n96 ) );
  NAND2_X1 u1_u7_u6_U57 (.ZN( u1_u7_u6_n100 ) , .A2( u1_u7_u6_n92 ) , .A1( u1_u7_u6_n98 ) );
  NAND2_X1 u1_u7_u6_U58 (.ZN( u1_u7_u6_n122 ) , .A1( u1_u7_u6_n94 ) , .A2( u1_u7_u6_n97 ) );
  INV_X1 u1_u7_u6_U59 (.A( u1_u7_u6_n139 ) , .ZN( u1_u7_u6_n160 ) );
  AOI22_X1 u1_u7_u6_U6 (.B2( u1_u7_u6_n101 ) , .A1( u1_u7_u6_n102 ) , .ZN( u1_u7_u6_n103 ) , .B1( u1_u7_u6_n160 ) , .A2( u1_u7_u6_n161 ) );
  NAND2_X1 u1_u7_u6_U60 (.ZN( u1_u7_u6_n113 ) , .A1( u1_u7_u6_n96 ) , .A2( u1_u7_u6_n98 ) );
  NOR2_X1 u1_u7_u6_U61 (.A2( u1_u7_X_40 ) , .A1( u1_u7_X_41 ) , .ZN( u1_u7_u6_n126 ) );
  NOR2_X1 u1_u7_u6_U62 (.A2( u1_u7_X_39 ) , .A1( u1_u7_X_42 ) , .ZN( u1_u7_u6_n92 ) );
  NOR2_X1 u1_u7_u6_U63 (.A2( u1_u7_X_39 ) , .A1( u1_u7_u6_n156 ) , .ZN( u1_u7_u6_n97 ) );
  NOR2_X1 u1_u7_u6_U64 (.A2( u1_u7_X_38 ) , .A1( u1_u7_u6_n165 ) , .ZN( u1_u7_u6_n95 ) );
  NOR2_X1 u1_u7_u6_U65 (.A2( u1_u7_X_41 ) , .ZN( u1_u7_u6_n111 ) , .A1( u1_u7_u6_n157 ) );
  NOR2_X1 u1_u7_u6_U66 (.A2( u1_u7_X_37 ) , .A1( u1_u7_u6_n162 ) , .ZN( u1_u7_u6_n94 ) );
  NOR2_X1 u1_u7_u6_U67 (.A2( u1_u7_X_37 ) , .A1( u1_u7_X_38 ) , .ZN( u1_u7_u6_n91 ) );
  NAND2_X1 u1_u7_u6_U68 (.A1( u1_u7_X_41 ) , .ZN( u1_u7_u6_n144 ) , .A2( u1_u7_u6_n157 ) );
  NAND2_X1 u1_u7_u6_U69 (.A2( u1_u7_X_40 ) , .A1( u1_u7_X_41 ) , .ZN( u1_u7_u6_n139 ) );
  NOR2_X1 u1_u7_u6_U7 (.A1( u1_u7_u6_n118 ) , .ZN( u1_u7_u6_n143 ) , .A2( u1_u7_u6_n168 ) );
  AND2_X1 u1_u7_u6_U70 (.A1( u1_u7_X_39 ) , .A2( u1_u7_u6_n156 ) , .ZN( u1_u7_u6_n96 ) );
  AND2_X1 u1_u7_u6_U71 (.A1( u1_u7_X_39 ) , .A2( u1_u7_X_42 ) , .ZN( u1_u7_u6_n99 ) );
  INV_X1 u1_u7_u6_U72 (.A( u1_u7_X_40 ) , .ZN( u1_u7_u6_n157 ) );
  INV_X1 u1_u7_u6_U73 (.A( u1_u7_X_37 ) , .ZN( u1_u7_u6_n165 ) );
  INV_X1 u1_u7_u6_U74 (.A( u1_u7_X_38 ) , .ZN( u1_u7_u6_n162 ) );
  INV_X1 u1_u7_u6_U75 (.A( u1_u7_X_42 ) , .ZN( u1_u7_u6_n156 ) );
  NAND4_X1 u1_u7_u6_U76 (.ZN( u1_out7_12 ) , .A4( u1_u7_u6_n114 ) , .A3( u1_u7_u6_n115 ) , .A2( u1_u7_u6_n116 ) , .A1( u1_u7_u6_n117 ) );
  OAI22_X1 u1_u7_u6_U77 (.B2( u1_u7_u6_n111 ) , .ZN( u1_u7_u6_n116 ) , .B1( u1_u7_u6_n126 ) , .A2( u1_u7_u6_n164 ) , .A1( u1_u7_u6_n167 ) );
  OAI21_X1 u1_u7_u6_U78 (.A( u1_u7_u6_n108 ) , .ZN( u1_u7_u6_n117 ) , .B2( u1_u7_u6_n141 ) , .B1( u1_u7_u6_n163 ) );
  NAND4_X1 u1_u7_u6_U79 (.ZN( u1_out7_32 ) , .A4( u1_u7_u6_n103 ) , .A3( u1_u7_u6_n104 ) , .A2( u1_u7_u6_n105 ) , .A1( u1_u7_u6_n106 ) );
  AOI21_X1 u1_u7_u6_U8 (.B1( u1_u7_u6_n107 ) , .B2( u1_u7_u6_n132 ) , .A( u1_u7_u6_n158 ) , .ZN( u1_u7_u6_n88 ) );
  AOI22_X1 u1_u7_u6_U80 (.ZN( u1_u7_u6_n105 ) , .A2( u1_u7_u6_n108 ) , .A1( u1_u7_u6_n118 ) , .B2( u1_u7_u6_n126 ) , .B1( u1_u7_u6_n171 ) );
  AOI22_X1 u1_u7_u6_U81 (.ZN( u1_u7_u6_n104 ) , .A1( u1_u7_u6_n111 ) , .B1( u1_u7_u6_n124 ) , .B2( u1_u7_u6_n151 ) , .A2( u1_u7_u6_n93 ) );
  OAI211_X1 u1_u7_u6_U82 (.ZN( u1_out7_7 ) , .B( u1_u7_u6_n153 ) , .C2( u1_u7_u6_n154 ) , .C1( u1_u7_u6_n155 ) , .A( u1_u7_u6_n174 ) );
  NOR3_X1 u1_u7_u6_U83 (.A1( u1_u7_u6_n141 ) , .ZN( u1_u7_u6_n154 ) , .A3( u1_u7_u6_n164 ) , .A2( u1_u7_u6_n171 ) );
  AOI211_X1 u1_u7_u6_U84 (.B( u1_u7_u6_n149 ) , .A( u1_u7_u6_n150 ) , .C2( u1_u7_u6_n151 ) , .C1( u1_u7_u6_n152 ) , .ZN( u1_u7_u6_n153 ) );
  OAI211_X1 u1_u7_u6_U85 (.ZN( u1_out7_22 ) , .B( u1_u7_u6_n137 ) , .A( u1_u7_u6_n138 ) , .C2( u1_u7_u6_n139 ) , .C1( u1_u7_u6_n140 ) );
  AOI22_X1 u1_u7_u6_U86 (.B1( u1_u7_u6_n124 ) , .A2( u1_u7_u6_n125 ) , .A1( u1_u7_u6_n126 ) , .ZN( u1_u7_u6_n138 ) , .B2( u1_u7_u6_n161 ) );
  AND4_X1 u1_u7_u6_U87 (.A3( u1_u7_u6_n119 ) , .A1( u1_u7_u6_n120 ) , .A4( u1_u7_u6_n129 ) , .ZN( u1_u7_u6_n140 ) , .A2( u1_u7_u6_n143 ) );
  NAND3_X1 u1_u7_u6_U88 (.A2( u1_u7_u6_n123 ) , .ZN( u1_u7_u6_n125 ) , .A1( u1_u7_u6_n130 ) , .A3( u1_u7_u6_n131 ) );
  NAND3_X1 u1_u7_u6_U89 (.A3( u1_u7_u6_n133 ) , .ZN( u1_u7_u6_n141 ) , .A1( u1_u7_u6_n145 ) , .A2( u1_u7_u6_n148 ) );
  AOI21_X1 u1_u7_u6_U9 (.B2( u1_u7_u6_n147 ) , .B1( u1_u7_u6_n148 ) , .ZN( u1_u7_u6_n149 ) , .A( u1_u7_u6_n158 ) );
  NAND3_X1 u1_u7_u6_U90 (.ZN( u1_u7_u6_n101 ) , .A3( u1_u7_u6_n107 ) , .A2( u1_u7_u6_n121 ) , .A1( u1_u7_u6_n127 ) );
  NAND3_X1 u1_u7_u6_U91 (.ZN( u1_u7_u6_n102 ) , .A3( u1_u7_u6_n130 ) , .A2( u1_u7_u6_n145 ) , .A1( u1_u7_u6_n166 ) );
  NAND3_X1 u1_u7_u6_U92 (.A3( u1_u7_u6_n113 ) , .A1( u1_u7_u6_n119 ) , .A2( u1_u7_u6_n123 ) , .ZN( u1_u7_u6_n93 ) );
  NAND3_X1 u1_u7_u6_U93 (.ZN( u1_u7_u6_n142 ) , .A2( u1_u7_u6_n172 ) , .A3( u1_u7_u6_n89 ) , .A1( u1_u7_u6_n90 ) );
  XOR2_X1 u1_u8_U13 (.B( u1_K9_42 ) , .A( u1_R7_29 ) , .Z( u1_u8_X_42 ) );
  XOR2_X1 u1_u8_U14 (.B( u1_K9_41 ) , .A( u1_R7_28 ) , .Z( u1_u8_X_41 ) );
  XOR2_X1 u1_u8_U15 (.B( u1_K9_40 ) , .A( u1_R7_27 ) , .Z( u1_u8_X_40 ) );
  XOR2_X1 u1_u8_U17 (.B( u1_K9_39 ) , .A( u1_R7_26 ) , .Z( u1_u8_X_39 ) );
  XOR2_X1 u1_u8_U18 (.B( u1_K9_38 ) , .A( u1_R7_25 ) , .Z( u1_u8_X_38 ) );
  XOR2_X1 u1_u8_U19 (.B( u1_K9_37 ) , .A( u1_R7_24 ) , .Z( u1_u8_X_37 ) );
  XOR2_X1 u1_u8_U20 (.B( u1_K9_36 ) , .A( u1_R7_25 ) , .Z( u1_u8_X_36 ) );
  XOR2_X1 u1_u8_U21 (.B( u1_K9_35 ) , .A( u1_R7_24 ) , .Z( u1_u8_X_35 ) );
  XOR2_X1 u1_u8_U22 (.B( u1_K9_34 ) , .A( u1_R7_23 ) , .Z( u1_u8_X_34 ) );
  XOR2_X1 u1_u8_U23 (.B( u1_K9_33 ) , .A( u1_R7_22 ) , .Z( u1_u8_X_33 ) );
  XOR2_X1 u1_u8_U24 (.B( u1_K9_32 ) , .A( u1_R7_21 ) , .Z( u1_u8_X_32 ) );
  XOR2_X1 u1_u8_U25 (.B( u1_K9_31 ) , .A( u1_R7_20 ) , .Z( u1_u8_X_31 ) );
  NOR2_X1 u1_u8_u5_U10 (.ZN( u1_u8_u5_n135 ) , .A1( u1_u8_u5_n173 ) , .A2( u1_u8_u5_n176 ) );
  NOR3_X1 u1_u8_u5_U100 (.A3( u1_u8_u5_n141 ) , .A1( u1_u8_u5_n142 ) , .ZN( u1_u8_u5_n143 ) , .A2( u1_u8_u5_n191 ) );
  NAND4_X1 u1_u8_u5_U101 (.ZN( u1_out8_4 ) , .A4( u1_u8_u5_n112 ) , .A2( u1_u8_u5_n113 ) , .A1( u1_u8_u5_n114 ) , .A3( u1_u8_u5_n195 ) );
  AOI211_X1 u1_u8_u5_U102 (.A( u1_u8_u5_n110 ) , .C1( u1_u8_u5_n111 ) , .ZN( u1_u8_u5_n112 ) , .B( u1_u8_u5_n118 ) , .C2( u1_u8_u5_n177 ) );
  INV_X1 u1_u8_u5_U103 (.A( u1_u8_u5_n102 ) , .ZN( u1_u8_u5_n195 ) );
  NAND3_X1 u1_u8_u5_U104 (.A2( u1_u8_u5_n154 ) , .A3( u1_u8_u5_n158 ) , .A1( u1_u8_u5_n161 ) , .ZN( u1_u8_u5_n99 ) );
  INV_X1 u1_u8_u5_U11 (.A( u1_u8_u5_n121 ) , .ZN( u1_u8_u5_n177 ) );
  NOR2_X1 u1_u8_u5_U12 (.ZN( u1_u8_u5_n160 ) , .A2( u1_u8_u5_n173 ) , .A1( u1_u8_u5_n177 ) );
  INV_X1 u1_u8_u5_U13 (.A( u1_u8_u5_n150 ) , .ZN( u1_u8_u5_n174 ) );
  AOI21_X1 u1_u8_u5_U14 (.A( u1_u8_u5_n160 ) , .B2( u1_u8_u5_n161 ) , .ZN( u1_u8_u5_n162 ) , .B1( u1_u8_u5_n192 ) );
  INV_X1 u1_u8_u5_U15 (.A( u1_u8_u5_n159 ) , .ZN( u1_u8_u5_n192 ) );
  AOI21_X1 u1_u8_u5_U16 (.A( u1_u8_u5_n156 ) , .B2( u1_u8_u5_n157 ) , .B1( u1_u8_u5_n158 ) , .ZN( u1_u8_u5_n163 ) );
  AOI21_X1 u1_u8_u5_U17 (.B2( u1_u8_u5_n139 ) , .B1( u1_u8_u5_n140 ) , .ZN( u1_u8_u5_n141 ) , .A( u1_u8_u5_n150 ) );
  OAI21_X1 u1_u8_u5_U18 (.A( u1_u8_u5_n133 ) , .B2( u1_u8_u5_n134 ) , .B1( u1_u8_u5_n135 ) , .ZN( u1_u8_u5_n142 ) );
  OAI21_X1 u1_u8_u5_U19 (.ZN( u1_u8_u5_n133 ) , .B2( u1_u8_u5_n147 ) , .A( u1_u8_u5_n173 ) , .B1( u1_u8_u5_n188 ) );
  NAND2_X1 u1_u8_u5_U20 (.A2( u1_u8_u5_n119 ) , .A1( u1_u8_u5_n123 ) , .ZN( u1_u8_u5_n137 ) );
  INV_X1 u1_u8_u5_U21 (.A( u1_u8_u5_n155 ) , .ZN( u1_u8_u5_n194 ) );
  NAND2_X1 u1_u8_u5_U22 (.A1( u1_u8_u5_n121 ) , .ZN( u1_u8_u5_n132 ) , .A2( u1_u8_u5_n172 ) );
  NAND2_X1 u1_u8_u5_U23 (.A2( u1_u8_u5_n122 ) , .ZN( u1_u8_u5_n136 ) , .A1( u1_u8_u5_n154 ) );
  NAND2_X1 u1_u8_u5_U24 (.A2( u1_u8_u5_n119 ) , .A1( u1_u8_u5_n120 ) , .ZN( u1_u8_u5_n159 ) );
  INV_X1 u1_u8_u5_U25 (.A( u1_u8_u5_n156 ) , .ZN( u1_u8_u5_n175 ) );
  INV_X1 u1_u8_u5_U26 (.A( u1_u8_u5_n158 ) , .ZN( u1_u8_u5_n188 ) );
  INV_X1 u1_u8_u5_U27 (.A( u1_u8_u5_n152 ) , .ZN( u1_u8_u5_n179 ) );
  INV_X1 u1_u8_u5_U28 (.A( u1_u8_u5_n140 ) , .ZN( u1_u8_u5_n182 ) );
  INV_X1 u1_u8_u5_U29 (.A( u1_u8_u5_n151 ) , .ZN( u1_u8_u5_n183 ) );
  NOR2_X1 u1_u8_u5_U3 (.ZN( u1_u8_u5_n134 ) , .A1( u1_u8_u5_n183 ) , .A2( u1_u8_u5_n190 ) );
  INV_X1 u1_u8_u5_U30 (.A( u1_u8_u5_n123 ) , .ZN( u1_u8_u5_n185 ) );
  INV_X1 u1_u8_u5_U31 (.A( u1_u8_u5_n161 ) , .ZN( u1_u8_u5_n184 ) );
  INV_X1 u1_u8_u5_U32 (.A( u1_u8_u5_n139 ) , .ZN( u1_u8_u5_n189 ) );
  INV_X1 u1_u8_u5_U33 (.A( u1_u8_u5_n157 ) , .ZN( u1_u8_u5_n190 ) );
  INV_X1 u1_u8_u5_U34 (.A( u1_u8_u5_n120 ) , .ZN( u1_u8_u5_n193 ) );
  NAND2_X1 u1_u8_u5_U35 (.ZN( u1_u8_u5_n111 ) , .A1( u1_u8_u5_n140 ) , .A2( u1_u8_u5_n155 ) );
  INV_X1 u1_u8_u5_U36 (.A( u1_u8_u5_n117 ) , .ZN( u1_u8_u5_n196 ) );
  OAI221_X1 u1_u8_u5_U37 (.A( u1_u8_u5_n116 ) , .ZN( u1_u8_u5_n117 ) , .B2( u1_u8_u5_n119 ) , .C1( u1_u8_u5_n153 ) , .C2( u1_u8_u5_n158 ) , .B1( u1_u8_u5_n172 ) );
  AOI222_X1 u1_u8_u5_U38 (.ZN( u1_u8_u5_n116 ) , .B2( u1_u8_u5_n145 ) , .C1( u1_u8_u5_n148 ) , .A2( u1_u8_u5_n174 ) , .C2( u1_u8_u5_n177 ) , .B1( u1_u8_u5_n187 ) , .A1( u1_u8_u5_n193 ) );
  INV_X1 u1_u8_u5_U39 (.A( u1_u8_u5_n115 ) , .ZN( u1_u8_u5_n187 ) );
  INV_X1 u1_u8_u5_U4 (.A( u1_u8_u5_n138 ) , .ZN( u1_u8_u5_n191 ) );
  NOR2_X1 u1_u8_u5_U40 (.ZN( u1_u8_u5_n100 ) , .A1( u1_u8_u5_n170 ) , .A2( u1_u8_u5_n180 ) );
  OAI221_X1 u1_u8_u5_U41 (.A( u1_u8_u5_n101 ) , .ZN( u1_u8_u5_n102 ) , .C2( u1_u8_u5_n115 ) , .C1( u1_u8_u5_n126 ) , .B1( u1_u8_u5_n134 ) , .B2( u1_u8_u5_n160 ) );
  OAI21_X1 u1_u8_u5_U42 (.ZN( u1_u8_u5_n101 ) , .B1( u1_u8_u5_n137 ) , .A( u1_u8_u5_n146 ) , .B2( u1_u8_u5_n147 ) );
  AOI22_X1 u1_u8_u5_U43 (.B2( u1_u8_u5_n131 ) , .A2( u1_u8_u5_n146 ) , .ZN( u1_u8_u5_n169 ) , .B1( u1_u8_u5_n174 ) , .A1( u1_u8_u5_n185 ) );
  NOR2_X1 u1_u8_u5_U44 (.A1( u1_u8_u5_n146 ) , .ZN( u1_u8_u5_n150 ) , .A2( u1_u8_u5_n173 ) );
  AOI21_X1 u1_u8_u5_U45 (.A( u1_u8_u5_n118 ) , .B2( u1_u8_u5_n145 ) , .ZN( u1_u8_u5_n168 ) , .B1( u1_u8_u5_n186 ) );
  INV_X1 u1_u8_u5_U46 (.A( u1_u8_u5_n122 ) , .ZN( u1_u8_u5_n186 ) );
  NOR2_X1 u1_u8_u5_U47 (.A1( u1_u8_u5_n146 ) , .ZN( u1_u8_u5_n152 ) , .A2( u1_u8_u5_n176 ) );
  NOR2_X1 u1_u8_u5_U48 (.A1( u1_u8_u5_n115 ) , .ZN( u1_u8_u5_n118 ) , .A2( u1_u8_u5_n153 ) );
  NOR2_X1 u1_u8_u5_U49 (.A2( u1_u8_u5_n145 ) , .ZN( u1_u8_u5_n156 ) , .A1( u1_u8_u5_n174 ) );
  OAI21_X1 u1_u8_u5_U5 (.B2( u1_u8_u5_n136 ) , .B1( u1_u8_u5_n137 ) , .ZN( u1_u8_u5_n138 ) , .A( u1_u8_u5_n177 ) );
  NOR2_X1 u1_u8_u5_U50 (.ZN( u1_u8_u5_n121 ) , .A2( u1_u8_u5_n145 ) , .A1( u1_u8_u5_n176 ) );
  AOI22_X1 u1_u8_u5_U51 (.ZN( u1_u8_u5_n114 ) , .A2( u1_u8_u5_n137 ) , .A1( u1_u8_u5_n145 ) , .B2( u1_u8_u5_n175 ) , .B1( u1_u8_u5_n193 ) );
  OAI211_X1 u1_u8_u5_U52 (.B( u1_u8_u5_n124 ) , .A( u1_u8_u5_n125 ) , .C2( u1_u8_u5_n126 ) , .C1( u1_u8_u5_n127 ) , .ZN( u1_u8_u5_n128 ) );
  NOR3_X1 u1_u8_u5_U53 (.ZN( u1_u8_u5_n127 ) , .A1( u1_u8_u5_n136 ) , .A3( u1_u8_u5_n148 ) , .A2( u1_u8_u5_n182 ) );
  OAI21_X1 u1_u8_u5_U54 (.ZN( u1_u8_u5_n124 ) , .A( u1_u8_u5_n177 ) , .B2( u1_u8_u5_n183 ) , .B1( u1_u8_u5_n189 ) );
  OAI21_X1 u1_u8_u5_U55 (.ZN( u1_u8_u5_n125 ) , .A( u1_u8_u5_n174 ) , .B2( u1_u8_u5_n185 ) , .B1( u1_u8_u5_n190 ) );
  AOI21_X1 u1_u8_u5_U56 (.A( u1_u8_u5_n153 ) , .B2( u1_u8_u5_n154 ) , .B1( u1_u8_u5_n155 ) , .ZN( u1_u8_u5_n164 ) );
  AOI21_X1 u1_u8_u5_U57 (.ZN( u1_u8_u5_n110 ) , .B1( u1_u8_u5_n122 ) , .B2( u1_u8_u5_n139 ) , .A( u1_u8_u5_n153 ) );
  INV_X1 u1_u8_u5_U58 (.A( u1_u8_u5_n153 ) , .ZN( u1_u8_u5_n176 ) );
  INV_X1 u1_u8_u5_U59 (.A( u1_u8_u5_n126 ) , .ZN( u1_u8_u5_n173 ) );
  AOI222_X1 u1_u8_u5_U6 (.ZN( u1_u8_u5_n113 ) , .A1( u1_u8_u5_n131 ) , .C1( u1_u8_u5_n148 ) , .B2( u1_u8_u5_n174 ) , .C2( u1_u8_u5_n178 ) , .A2( u1_u8_u5_n179 ) , .B1( u1_u8_u5_n99 ) );
  AND2_X1 u1_u8_u5_U60 (.A2( u1_u8_u5_n104 ) , .A1( u1_u8_u5_n107 ) , .ZN( u1_u8_u5_n147 ) );
  AND2_X1 u1_u8_u5_U61 (.A2( u1_u8_u5_n104 ) , .A1( u1_u8_u5_n108 ) , .ZN( u1_u8_u5_n148 ) );
  NAND2_X1 u1_u8_u5_U62 (.A1( u1_u8_u5_n105 ) , .A2( u1_u8_u5_n106 ) , .ZN( u1_u8_u5_n158 ) );
  NAND2_X1 u1_u8_u5_U63 (.A2( u1_u8_u5_n108 ) , .A1( u1_u8_u5_n109 ) , .ZN( u1_u8_u5_n139 ) );
  NAND2_X1 u1_u8_u5_U64 (.A1( u1_u8_u5_n106 ) , .A2( u1_u8_u5_n108 ) , .ZN( u1_u8_u5_n119 ) );
  NAND2_X1 u1_u8_u5_U65 (.A2( u1_u8_u5_n103 ) , .A1( u1_u8_u5_n105 ) , .ZN( u1_u8_u5_n140 ) );
  NAND2_X1 u1_u8_u5_U66 (.A2( u1_u8_u5_n104 ) , .A1( u1_u8_u5_n105 ) , .ZN( u1_u8_u5_n155 ) );
  NAND2_X1 u1_u8_u5_U67 (.A2( u1_u8_u5_n106 ) , .A1( u1_u8_u5_n107 ) , .ZN( u1_u8_u5_n122 ) );
  NAND2_X1 u1_u8_u5_U68 (.A2( u1_u8_u5_n100 ) , .A1( u1_u8_u5_n106 ) , .ZN( u1_u8_u5_n115 ) );
  NAND2_X1 u1_u8_u5_U69 (.A2( u1_u8_u5_n100 ) , .A1( u1_u8_u5_n103 ) , .ZN( u1_u8_u5_n161 ) );
  INV_X1 u1_u8_u5_U7 (.A( u1_u8_u5_n135 ) , .ZN( u1_u8_u5_n178 ) );
  NAND2_X1 u1_u8_u5_U70 (.A1( u1_u8_u5_n105 ) , .A2( u1_u8_u5_n109 ) , .ZN( u1_u8_u5_n154 ) );
  INV_X1 u1_u8_u5_U71 (.A( u1_u8_u5_n146 ) , .ZN( u1_u8_u5_n172 ) );
  NAND2_X1 u1_u8_u5_U72 (.A1( u1_u8_u5_n103 ) , .A2( u1_u8_u5_n108 ) , .ZN( u1_u8_u5_n123 ) );
  NAND2_X1 u1_u8_u5_U73 (.A2( u1_u8_u5_n103 ) , .A1( u1_u8_u5_n107 ) , .ZN( u1_u8_u5_n151 ) );
  NAND2_X1 u1_u8_u5_U74 (.A2( u1_u8_u5_n107 ) , .A1( u1_u8_u5_n109 ) , .ZN( u1_u8_u5_n120 ) );
  NAND2_X1 u1_u8_u5_U75 (.A2( u1_u8_u5_n100 ) , .A1( u1_u8_u5_n109 ) , .ZN( u1_u8_u5_n157 ) );
  AND2_X1 u1_u8_u5_U76 (.A2( u1_u8_u5_n100 ) , .A1( u1_u8_u5_n104 ) , .ZN( u1_u8_u5_n131 ) );
  NOR2_X1 u1_u8_u5_U77 (.A2( u1_u8_X_34 ) , .A1( u1_u8_X_35 ) , .ZN( u1_u8_u5_n145 ) );
  NOR2_X1 u1_u8_u5_U78 (.A2( u1_u8_X_34 ) , .ZN( u1_u8_u5_n146 ) , .A1( u1_u8_u5_n171 ) );
  NOR2_X1 u1_u8_u5_U79 (.A2( u1_u8_X_31 ) , .A1( u1_u8_X_32 ) , .ZN( u1_u8_u5_n103 ) );
  OAI22_X1 u1_u8_u5_U8 (.B2( u1_u8_u5_n149 ) , .B1( u1_u8_u5_n150 ) , .A2( u1_u8_u5_n151 ) , .A1( u1_u8_u5_n152 ) , .ZN( u1_u8_u5_n165 ) );
  NOR2_X1 u1_u8_u5_U80 (.A2( u1_u8_X_36 ) , .ZN( u1_u8_u5_n105 ) , .A1( u1_u8_u5_n180 ) );
  NOR2_X1 u1_u8_u5_U81 (.A2( u1_u8_X_33 ) , .ZN( u1_u8_u5_n108 ) , .A1( u1_u8_u5_n170 ) );
  NOR2_X1 u1_u8_u5_U82 (.A2( u1_u8_X_33 ) , .A1( u1_u8_X_36 ) , .ZN( u1_u8_u5_n107 ) );
  NOR2_X1 u1_u8_u5_U83 (.A2( u1_u8_X_31 ) , .ZN( u1_u8_u5_n104 ) , .A1( u1_u8_u5_n181 ) );
  NAND2_X1 u1_u8_u5_U84 (.A2( u1_u8_X_34 ) , .A1( u1_u8_X_35 ) , .ZN( u1_u8_u5_n153 ) );
  NAND2_X1 u1_u8_u5_U85 (.A1( u1_u8_X_34 ) , .ZN( u1_u8_u5_n126 ) , .A2( u1_u8_u5_n171 ) );
  AND2_X1 u1_u8_u5_U86 (.A1( u1_u8_X_31 ) , .A2( u1_u8_X_32 ) , .ZN( u1_u8_u5_n106 ) );
  AND2_X1 u1_u8_u5_U87 (.A1( u1_u8_X_31 ) , .ZN( u1_u8_u5_n109 ) , .A2( u1_u8_u5_n181 ) );
  INV_X1 u1_u8_u5_U88 (.A( u1_u8_X_33 ) , .ZN( u1_u8_u5_n180 ) );
  INV_X1 u1_u8_u5_U89 (.A( u1_u8_X_35 ) , .ZN( u1_u8_u5_n171 ) );
  NOR3_X1 u1_u8_u5_U9 (.A2( u1_u8_u5_n147 ) , .A1( u1_u8_u5_n148 ) , .ZN( u1_u8_u5_n149 ) , .A3( u1_u8_u5_n194 ) );
  INV_X1 u1_u8_u5_U90 (.A( u1_u8_X_36 ) , .ZN( u1_u8_u5_n170 ) );
  INV_X1 u1_u8_u5_U91 (.A( u1_u8_X_32 ) , .ZN( u1_u8_u5_n181 ) );
  NAND4_X1 u1_u8_u5_U92 (.ZN( u1_out8_29 ) , .A4( u1_u8_u5_n129 ) , .A3( u1_u8_u5_n130 ) , .A2( u1_u8_u5_n168 ) , .A1( u1_u8_u5_n196 ) );
  AOI221_X1 u1_u8_u5_U93 (.A( u1_u8_u5_n128 ) , .ZN( u1_u8_u5_n129 ) , .C2( u1_u8_u5_n132 ) , .B2( u1_u8_u5_n159 ) , .B1( u1_u8_u5_n176 ) , .C1( u1_u8_u5_n184 ) );
  AOI222_X1 u1_u8_u5_U94 (.ZN( u1_u8_u5_n130 ) , .A2( u1_u8_u5_n146 ) , .B1( u1_u8_u5_n147 ) , .C2( u1_u8_u5_n175 ) , .B2( u1_u8_u5_n179 ) , .A1( u1_u8_u5_n188 ) , .C1( u1_u8_u5_n194 ) );
  NAND4_X1 u1_u8_u5_U95 (.ZN( u1_out8_19 ) , .A4( u1_u8_u5_n166 ) , .A3( u1_u8_u5_n167 ) , .A2( u1_u8_u5_n168 ) , .A1( u1_u8_u5_n169 ) );
  AOI22_X1 u1_u8_u5_U96 (.B2( u1_u8_u5_n145 ) , .A2( u1_u8_u5_n146 ) , .ZN( u1_u8_u5_n167 ) , .B1( u1_u8_u5_n182 ) , .A1( u1_u8_u5_n189 ) );
  NOR4_X1 u1_u8_u5_U97 (.A4( u1_u8_u5_n162 ) , .A3( u1_u8_u5_n163 ) , .A2( u1_u8_u5_n164 ) , .A1( u1_u8_u5_n165 ) , .ZN( u1_u8_u5_n166 ) );
  NAND4_X1 u1_u8_u5_U98 (.ZN( u1_out8_11 ) , .A4( u1_u8_u5_n143 ) , .A3( u1_u8_u5_n144 ) , .A2( u1_u8_u5_n169 ) , .A1( u1_u8_u5_n196 ) );
  AOI22_X1 u1_u8_u5_U99 (.A2( u1_u8_u5_n132 ) , .ZN( u1_u8_u5_n144 ) , .B2( u1_u8_u5_n145 ) , .B1( u1_u8_u5_n184 ) , .A1( u1_u8_u5_n194 ) );
  AOI22_X1 u1_u8_u6_U10 (.A2( u1_u8_u6_n151 ) , .B2( u1_u8_u6_n161 ) , .A1( u1_u8_u6_n167 ) , .B1( u1_u8_u6_n170 ) , .ZN( u1_u8_u6_n89 ) );
  AOI21_X1 u1_u8_u6_U11 (.B1( u1_u8_u6_n107 ) , .B2( u1_u8_u6_n132 ) , .A( u1_u8_u6_n158 ) , .ZN( u1_u8_u6_n88 ) );
  AOI21_X1 u1_u8_u6_U12 (.B2( u1_u8_u6_n147 ) , .B1( u1_u8_u6_n148 ) , .ZN( u1_u8_u6_n149 ) , .A( u1_u8_u6_n158 ) );
  AOI21_X1 u1_u8_u6_U13 (.ZN( u1_u8_u6_n106 ) , .A( u1_u8_u6_n142 ) , .B2( u1_u8_u6_n159 ) , .B1( u1_u8_u6_n164 ) );
  INV_X1 u1_u8_u6_U14 (.A( u1_u8_u6_n155 ) , .ZN( u1_u8_u6_n161 ) );
  INV_X1 u1_u8_u6_U15 (.A( u1_u8_u6_n128 ) , .ZN( u1_u8_u6_n164 ) );
  NAND2_X1 u1_u8_u6_U16 (.ZN( u1_u8_u6_n110 ) , .A1( u1_u8_u6_n122 ) , .A2( u1_u8_u6_n129 ) );
  NAND2_X1 u1_u8_u6_U17 (.ZN( u1_u8_u6_n124 ) , .A2( u1_u8_u6_n146 ) , .A1( u1_u8_u6_n148 ) );
  INV_X1 u1_u8_u6_U18 (.A( u1_u8_u6_n132 ) , .ZN( u1_u8_u6_n171 ) );
  AND2_X1 u1_u8_u6_U19 (.A1( u1_u8_u6_n100 ) , .ZN( u1_u8_u6_n130 ) , .A2( u1_u8_u6_n147 ) );
  INV_X1 u1_u8_u6_U20 (.A( u1_u8_u6_n127 ) , .ZN( u1_u8_u6_n173 ) );
  INV_X1 u1_u8_u6_U21 (.A( u1_u8_u6_n121 ) , .ZN( u1_u8_u6_n167 ) );
  INV_X1 u1_u8_u6_U22 (.A( u1_u8_u6_n100 ) , .ZN( u1_u8_u6_n169 ) );
  INV_X1 u1_u8_u6_U23 (.A( u1_u8_u6_n123 ) , .ZN( u1_u8_u6_n170 ) );
  INV_X1 u1_u8_u6_U24 (.A( u1_u8_u6_n113 ) , .ZN( u1_u8_u6_n168 ) );
  AND2_X1 u1_u8_u6_U25 (.A1( u1_u8_u6_n107 ) , .A2( u1_u8_u6_n119 ) , .ZN( u1_u8_u6_n133 ) );
  AND2_X1 u1_u8_u6_U26 (.A2( u1_u8_u6_n121 ) , .A1( u1_u8_u6_n122 ) , .ZN( u1_u8_u6_n131 ) );
  AND3_X1 u1_u8_u6_U27 (.ZN( u1_u8_u6_n120 ) , .A2( u1_u8_u6_n127 ) , .A1( u1_u8_u6_n132 ) , .A3( u1_u8_u6_n145 ) );
  INV_X1 u1_u8_u6_U28 (.A( u1_u8_u6_n146 ) , .ZN( u1_u8_u6_n163 ) );
  AOI222_X1 u1_u8_u6_U29 (.ZN( u1_u8_u6_n114 ) , .A1( u1_u8_u6_n118 ) , .A2( u1_u8_u6_n126 ) , .B2( u1_u8_u6_n151 ) , .C2( u1_u8_u6_n159 ) , .C1( u1_u8_u6_n168 ) , .B1( u1_u8_u6_n169 ) );
  INV_X1 u1_u8_u6_U3 (.A( u1_u8_u6_n110 ) , .ZN( u1_u8_u6_n166 ) );
  NOR2_X1 u1_u8_u6_U30 (.A1( u1_u8_u6_n162 ) , .A2( u1_u8_u6_n165 ) , .ZN( u1_u8_u6_n98 ) );
  AOI211_X1 u1_u8_u6_U31 (.B( u1_u8_u6_n134 ) , .A( u1_u8_u6_n135 ) , .C1( u1_u8_u6_n136 ) , .ZN( u1_u8_u6_n137 ) , .C2( u1_u8_u6_n151 ) );
  AOI21_X1 u1_u8_u6_U32 (.B2( u1_u8_u6_n132 ) , .B1( u1_u8_u6_n133 ) , .ZN( u1_u8_u6_n134 ) , .A( u1_u8_u6_n158 ) );
  NAND4_X1 u1_u8_u6_U33 (.A4( u1_u8_u6_n127 ) , .A3( u1_u8_u6_n128 ) , .A2( u1_u8_u6_n129 ) , .A1( u1_u8_u6_n130 ) , .ZN( u1_u8_u6_n136 ) );
  AOI21_X1 u1_u8_u6_U34 (.B1( u1_u8_u6_n131 ) , .ZN( u1_u8_u6_n135 ) , .A( u1_u8_u6_n144 ) , .B2( u1_u8_u6_n146 ) );
  NAND2_X1 u1_u8_u6_U35 (.A1( u1_u8_u6_n144 ) , .ZN( u1_u8_u6_n151 ) , .A2( u1_u8_u6_n158 ) );
  NAND2_X1 u1_u8_u6_U36 (.ZN( u1_u8_u6_n132 ) , .A1( u1_u8_u6_n91 ) , .A2( u1_u8_u6_n97 ) );
  AOI22_X1 u1_u8_u6_U37 (.B2( u1_u8_u6_n110 ) , .B1( u1_u8_u6_n111 ) , .A1( u1_u8_u6_n112 ) , .ZN( u1_u8_u6_n115 ) , .A2( u1_u8_u6_n161 ) );
  NAND4_X1 u1_u8_u6_U38 (.A3( u1_u8_u6_n109 ) , .ZN( u1_u8_u6_n112 ) , .A4( u1_u8_u6_n132 ) , .A2( u1_u8_u6_n147 ) , .A1( u1_u8_u6_n166 ) );
  NOR2_X1 u1_u8_u6_U39 (.ZN( u1_u8_u6_n109 ) , .A1( u1_u8_u6_n170 ) , .A2( u1_u8_u6_n173 ) );
  INV_X1 u1_u8_u6_U4 (.A( u1_u8_u6_n142 ) , .ZN( u1_u8_u6_n174 ) );
  NOR2_X1 u1_u8_u6_U40 (.A2( u1_u8_u6_n126 ) , .ZN( u1_u8_u6_n155 ) , .A1( u1_u8_u6_n160 ) );
  NAND2_X1 u1_u8_u6_U41 (.ZN( u1_u8_u6_n146 ) , .A2( u1_u8_u6_n94 ) , .A1( u1_u8_u6_n99 ) );
  AOI21_X1 u1_u8_u6_U42 (.A( u1_u8_u6_n144 ) , .B2( u1_u8_u6_n145 ) , .B1( u1_u8_u6_n146 ) , .ZN( u1_u8_u6_n150 ) );
  INV_X1 u1_u8_u6_U43 (.A( u1_u8_u6_n111 ) , .ZN( u1_u8_u6_n158 ) );
  NAND2_X1 u1_u8_u6_U44 (.ZN( u1_u8_u6_n127 ) , .A1( u1_u8_u6_n91 ) , .A2( u1_u8_u6_n92 ) );
  NAND2_X1 u1_u8_u6_U45 (.ZN( u1_u8_u6_n129 ) , .A2( u1_u8_u6_n95 ) , .A1( u1_u8_u6_n96 ) );
  INV_X1 u1_u8_u6_U46 (.A( u1_u8_u6_n144 ) , .ZN( u1_u8_u6_n159 ) );
  NAND2_X1 u1_u8_u6_U47 (.ZN( u1_u8_u6_n145 ) , .A2( u1_u8_u6_n97 ) , .A1( u1_u8_u6_n98 ) );
  NAND2_X1 u1_u8_u6_U48 (.ZN( u1_u8_u6_n148 ) , .A2( u1_u8_u6_n92 ) , .A1( u1_u8_u6_n94 ) );
  NAND2_X1 u1_u8_u6_U49 (.ZN( u1_u8_u6_n108 ) , .A2( u1_u8_u6_n139 ) , .A1( u1_u8_u6_n144 ) );
  NAND2_X1 u1_u8_u6_U5 (.A2( u1_u8_u6_n143 ) , .ZN( u1_u8_u6_n152 ) , .A1( u1_u8_u6_n166 ) );
  NAND2_X1 u1_u8_u6_U50 (.ZN( u1_u8_u6_n121 ) , .A2( u1_u8_u6_n95 ) , .A1( u1_u8_u6_n97 ) );
  NAND2_X1 u1_u8_u6_U51 (.ZN( u1_u8_u6_n107 ) , .A2( u1_u8_u6_n92 ) , .A1( u1_u8_u6_n95 ) );
  AND2_X1 u1_u8_u6_U52 (.ZN( u1_u8_u6_n118 ) , .A2( u1_u8_u6_n91 ) , .A1( u1_u8_u6_n99 ) );
  NAND2_X1 u1_u8_u6_U53 (.ZN( u1_u8_u6_n147 ) , .A2( u1_u8_u6_n98 ) , .A1( u1_u8_u6_n99 ) );
  NAND2_X1 u1_u8_u6_U54 (.ZN( u1_u8_u6_n128 ) , .A1( u1_u8_u6_n94 ) , .A2( u1_u8_u6_n96 ) );
  NAND2_X1 u1_u8_u6_U55 (.ZN( u1_u8_u6_n119 ) , .A2( u1_u8_u6_n95 ) , .A1( u1_u8_u6_n99 ) );
  NAND2_X1 u1_u8_u6_U56 (.ZN( u1_u8_u6_n123 ) , .A2( u1_u8_u6_n91 ) , .A1( u1_u8_u6_n96 ) );
  NAND2_X1 u1_u8_u6_U57 (.ZN( u1_u8_u6_n100 ) , .A2( u1_u8_u6_n92 ) , .A1( u1_u8_u6_n98 ) );
  NAND2_X1 u1_u8_u6_U58 (.ZN( u1_u8_u6_n122 ) , .A1( u1_u8_u6_n94 ) , .A2( u1_u8_u6_n97 ) );
  INV_X1 u1_u8_u6_U59 (.A( u1_u8_u6_n139 ) , .ZN( u1_u8_u6_n160 ) );
  AOI22_X1 u1_u8_u6_U6 (.B2( u1_u8_u6_n101 ) , .A1( u1_u8_u6_n102 ) , .ZN( u1_u8_u6_n103 ) , .B1( u1_u8_u6_n160 ) , .A2( u1_u8_u6_n161 ) );
  NAND2_X1 u1_u8_u6_U60 (.ZN( u1_u8_u6_n113 ) , .A1( u1_u8_u6_n96 ) , .A2( u1_u8_u6_n98 ) );
  NOR2_X1 u1_u8_u6_U61 (.A2( u1_u8_X_40 ) , .A1( u1_u8_X_41 ) , .ZN( u1_u8_u6_n126 ) );
  NOR2_X1 u1_u8_u6_U62 (.A2( u1_u8_X_39 ) , .A1( u1_u8_X_42 ) , .ZN( u1_u8_u6_n92 ) );
  NOR2_X1 u1_u8_u6_U63 (.A2( u1_u8_X_39 ) , .A1( u1_u8_u6_n156 ) , .ZN( u1_u8_u6_n97 ) );
  NOR2_X1 u1_u8_u6_U64 (.A2( u1_u8_X_38 ) , .A1( u1_u8_u6_n165 ) , .ZN( u1_u8_u6_n95 ) );
  NOR2_X1 u1_u8_u6_U65 (.A2( u1_u8_X_41 ) , .ZN( u1_u8_u6_n111 ) , .A1( u1_u8_u6_n157 ) );
  NOR2_X1 u1_u8_u6_U66 (.A2( u1_u8_X_37 ) , .A1( u1_u8_u6_n162 ) , .ZN( u1_u8_u6_n94 ) );
  NOR2_X1 u1_u8_u6_U67 (.A2( u1_u8_X_37 ) , .A1( u1_u8_X_38 ) , .ZN( u1_u8_u6_n91 ) );
  NAND2_X1 u1_u8_u6_U68 (.A1( u1_u8_X_41 ) , .ZN( u1_u8_u6_n144 ) , .A2( u1_u8_u6_n157 ) );
  NAND2_X1 u1_u8_u6_U69 (.A2( u1_u8_X_40 ) , .A1( u1_u8_X_41 ) , .ZN( u1_u8_u6_n139 ) );
  NOR2_X1 u1_u8_u6_U7 (.A1( u1_u8_u6_n118 ) , .ZN( u1_u8_u6_n143 ) , .A2( u1_u8_u6_n168 ) );
  AND2_X1 u1_u8_u6_U70 (.A1( u1_u8_X_39 ) , .A2( u1_u8_u6_n156 ) , .ZN( u1_u8_u6_n96 ) );
  AND2_X1 u1_u8_u6_U71 (.A1( u1_u8_X_39 ) , .A2( u1_u8_X_42 ) , .ZN( u1_u8_u6_n99 ) );
  INV_X1 u1_u8_u6_U72 (.A( u1_u8_X_40 ) , .ZN( u1_u8_u6_n157 ) );
  INV_X1 u1_u8_u6_U73 (.A( u1_u8_X_37 ) , .ZN( u1_u8_u6_n165 ) );
  INV_X1 u1_u8_u6_U74 (.A( u1_u8_X_38 ) , .ZN( u1_u8_u6_n162 ) );
  INV_X1 u1_u8_u6_U75 (.A( u1_u8_X_42 ) , .ZN( u1_u8_u6_n156 ) );
  NAND4_X1 u1_u8_u6_U76 (.ZN( u1_out8_12 ) , .A4( u1_u8_u6_n114 ) , .A3( u1_u8_u6_n115 ) , .A2( u1_u8_u6_n116 ) , .A1( u1_u8_u6_n117 ) );
  OAI22_X1 u1_u8_u6_U77 (.B2( u1_u8_u6_n111 ) , .ZN( u1_u8_u6_n116 ) , .B1( u1_u8_u6_n126 ) , .A2( u1_u8_u6_n164 ) , .A1( u1_u8_u6_n167 ) );
  OAI21_X1 u1_u8_u6_U78 (.A( u1_u8_u6_n108 ) , .ZN( u1_u8_u6_n117 ) , .B2( u1_u8_u6_n141 ) , .B1( u1_u8_u6_n163 ) );
  NAND4_X1 u1_u8_u6_U79 (.ZN( u1_out8_32 ) , .A4( u1_u8_u6_n103 ) , .A3( u1_u8_u6_n104 ) , .A2( u1_u8_u6_n105 ) , .A1( u1_u8_u6_n106 ) );
  OAI21_X1 u1_u8_u6_U8 (.A( u1_u8_u6_n159 ) , .B1( u1_u8_u6_n169 ) , .B2( u1_u8_u6_n173 ) , .ZN( u1_u8_u6_n90 ) );
  AOI22_X1 u1_u8_u6_U80 (.ZN( u1_u8_u6_n105 ) , .A2( u1_u8_u6_n108 ) , .A1( u1_u8_u6_n118 ) , .B2( u1_u8_u6_n126 ) , .B1( u1_u8_u6_n171 ) );
  AOI22_X1 u1_u8_u6_U81 (.ZN( u1_u8_u6_n104 ) , .A1( u1_u8_u6_n111 ) , .B1( u1_u8_u6_n124 ) , .B2( u1_u8_u6_n151 ) , .A2( u1_u8_u6_n93 ) );
  OAI211_X1 u1_u8_u6_U82 (.ZN( u1_out8_7 ) , .B( u1_u8_u6_n153 ) , .C2( u1_u8_u6_n154 ) , .C1( u1_u8_u6_n155 ) , .A( u1_u8_u6_n174 ) );
  NOR3_X1 u1_u8_u6_U83 (.A1( u1_u8_u6_n141 ) , .ZN( u1_u8_u6_n154 ) , .A3( u1_u8_u6_n164 ) , .A2( u1_u8_u6_n171 ) );
  AOI211_X1 u1_u8_u6_U84 (.B( u1_u8_u6_n149 ) , .A( u1_u8_u6_n150 ) , .C2( u1_u8_u6_n151 ) , .C1( u1_u8_u6_n152 ) , .ZN( u1_u8_u6_n153 ) );
  OAI211_X1 u1_u8_u6_U85 (.ZN( u1_out8_22 ) , .B( u1_u8_u6_n137 ) , .A( u1_u8_u6_n138 ) , .C2( u1_u8_u6_n139 ) , .C1( u1_u8_u6_n140 ) );
  AOI22_X1 u1_u8_u6_U86 (.B1( u1_u8_u6_n124 ) , .A2( u1_u8_u6_n125 ) , .A1( u1_u8_u6_n126 ) , .ZN( u1_u8_u6_n138 ) , .B2( u1_u8_u6_n161 ) );
  AND4_X1 u1_u8_u6_U87 (.A3( u1_u8_u6_n119 ) , .A1( u1_u8_u6_n120 ) , .A4( u1_u8_u6_n129 ) , .ZN( u1_u8_u6_n140 ) , .A2( u1_u8_u6_n143 ) );
  NAND3_X1 u1_u8_u6_U88 (.A2( u1_u8_u6_n123 ) , .ZN( u1_u8_u6_n125 ) , .A1( u1_u8_u6_n130 ) , .A3( u1_u8_u6_n131 ) );
  NAND3_X1 u1_u8_u6_U89 (.A3( u1_u8_u6_n133 ) , .ZN( u1_u8_u6_n141 ) , .A1( u1_u8_u6_n145 ) , .A2( u1_u8_u6_n148 ) );
  INV_X1 u1_u8_u6_U9 (.ZN( u1_u8_u6_n172 ) , .A( u1_u8_u6_n88 ) );
  NAND3_X1 u1_u8_u6_U90 (.ZN( u1_u8_u6_n101 ) , .A3( u1_u8_u6_n107 ) , .A2( u1_u8_u6_n121 ) , .A1( u1_u8_u6_n127 ) );
  NAND3_X1 u1_u8_u6_U91 (.ZN( u1_u8_u6_n102 ) , .A3( u1_u8_u6_n130 ) , .A2( u1_u8_u6_n145 ) , .A1( u1_u8_u6_n166 ) );
  NAND3_X1 u1_u8_u6_U92 (.A3( u1_u8_u6_n113 ) , .A1( u1_u8_u6_n119 ) , .A2( u1_u8_u6_n123 ) , .ZN( u1_u8_u6_n93 ) );
  NAND3_X1 u1_u8_u6_U93 (.ZN( u1_u8_u6_n142 ) , .A2( u1_u8_u6_n172 ) , .A3( u1_u8_u6_n89 ) , .A1( u1_u8_u6_n90 ) );
  OAI21_X1 u1_uk_U1004 (.ZN( u1_K14_46 ) , .B2( u1_uk_n1820 ) , .B1( u1_uk_n63 ) , .A( u1_uk_n961 ) );
  NAND2_X1 u1_uk_U1005 (.A1( u1_uk_K_r12_22 ) , .A2( u1_uk_n17 ) , .ZN( u1_uk_n961 ) );
  OAI21_X1 u1_uk_U1028 (.ZN( u1_K9_39 ) , .A( u1_uk_n1165 ) , .B2( u1_uk_n1601 ) , .B1( u1_uk_n60 ) );
  NAND2_X1 u1_uk_U1029 (.A1( u1_uk_K_r7_31 ) , .ZN( u1_uk_n1165 ) , .A2( u1_uk_n31 ) );
  OAI21_X1 u1_uk_U1030 (.ZN( u1_K14_44 ) , .B2( u1_uk_n1807 ) , .B1( u1_uk_n251 ) , .A( u1_uk_n959 ) );
  NAND2_X1 u1_uk_U1031 (.A1( u1_uk_K_r12_15 ) , .A2( u1_uk_n279 ) , .ZN( u1_uk_n959 ) );
  OAI21_X1 u1_uk_U1044 (.ZN( u1_K8_41 ) , .A( u1_uk_n1141 ) , .B2( u1_uk_n1547 ) , .B1( u1_uk_n155 ) );
  NAND2_X1 u1_uk_U1045 (.A1( u1_uk_K_r6_30 ) , .ZN( u1_uk_n1141 ) , .A2( u1_uk_n93 ) );
  OAI21_X1 u1_uk_U1058 (.ZN( u1_K14_40 ) , .B1( u1_uk_n109 ) , .B2( u1_uk_n1823 ) , .A( u1_uk_n958 ) );
  NAND2_X1 u1_uk_U1059 (.A1( u1_uk_K_r12_21 ) , .A2( u1_uk_n11 ) , .ZN( u1_uk_n958 ) );
  OAI21_X1 u1_uk_U1070 (.ZN( u1_K8_42 ) , .A( u1_uk_n1142 ) , .B2( u1_uk_n1540 ) , .B1( u1_uk_n155 ) );
  NAND2_X1 u1_uk_U1071 (.A1( u1_uk_K_r6_22 ) , .ZN( u1_uk_n1142 ) , .A2( u1_uk_n117 ) );
  OAI21_X1 u1_uk_U1103 (.ZN( u1_K13_28 ) , .B2( u1_uk_n1783 ) , .B1( u1_uk_n230 ) , .A( u1_uk_n695 ) );
  NAND2_X1 u1_uk_U1104 (.A1( u1_uk_K_r11_21 ) , .A2( u1_uk_n277 ) , .ZN( u1_uk_n695 ) );
  OAI21_X1 u1_uk_U1113 (.ZN( u1_K8_39 ) , .A( u1_uk_n1139 ) , .B2( u1_uk_n1556 ) , .B1( u1_uk_n203 ) );
  NAND2_X1 u1_uk_U1114 (.A1( u1_uk_K_r6_31 ) , .ZN( u1_uk_n1139 ) , .A2( u1_uk_n286 ) );
  INV_X1 u1_uk_U1139 (.ZN( u1_K11_30 ) , .A( u1_uk_n421 ) );
  AOI22_X1 u1_uk_U1140 (.B2( u1_uk_K_r9_1 ) , .A2( u1_uk_K_r9_9 ) , .B1( u1_uk_n182 ) , .A1( u1_uk_n231 ) , .ZN( u1_uk_n421 ) );
  INV_X1 u1_uk_U1161 (.ZN( u1_K7_25 ) , .A( u1_uk_n1114 ) );
  AOI22_X1 u1_uk_U1162 (.B2( u1_uk_K_r5_31 ) , .A2( u1_uk_K_r5_7 ) , .A1( u1_uk_n10 ) , .ZN( u1_uk_n1114 ) , .B1( u1_uk_n208 ) );
  OAI22_X1 u1_uk_U120 (.ZN( u1_K14_41 ) , .B1( u1_uk_n102 ) , .A2( u1_uk_n1806 ) , .B2( u1_uk_n1811 ) , .A1( u1_uk_n257 ) );
  INV_X1 u1_uk_U126 (.ZN( u1_K11_47 ) , .A( u1_uk_n472 ) );
  AOI22_X1 u1_uk_U127 (.B2( u1_uk_K_r9_15 ) , .A2( u1_uk_K_r9_23 ) , .B1( u1_uk_n164 ) , .A1( u1_uk_n223 ) , .ZN( u1_uk_n472 ) );
  INV_X1 u1_uk_U16 (.ZN( u1_uk_n109 ) , .A( u1_uk_n231 ) );
  INV_X1 u1_uk_U161 (.ZN( u1_K11_19 ) , .A( u1_uk_n386 ) );
  AOI22_X1 u1_uk_U162 (.B2( u1_uk_K_r9_10 ) , .A2( u1_uk_K_r9_48 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n222 ) , .ZN( u1_uk_n386 ) );
  OAI21_X1 u1_uk_U199 (.ZN( u1_K13_30 ) , .B2( u1_uk_n1776 ) , .A( u1_uk_n717 ) , .B1( u1_uk_n83 ) );
  NAND2_X1 u1_uk_U200 (.A1( u1_uk_K_r11_28 ) , .A2( u1_uk_n27 ) , .ZN( u1_uk_n717 ) );
  OAI22_X1 u1_uk_U233 (.ZN( u1_K13_31 ) , .B1( u1_uk_n100 ) , .B2( u1_uk_n1772 ) , .A2( u1_uk_n1790 ) , .A1( u1_uk_n207 ) );
  INV_X1 u1_uk_U24 (.ZN( u1_uk_n129 ) , .A( u1_uk_n223 ) );
  OAI22_X1 u1_uk_U245 (.ZN( u1_K9_31 ) , .B1( u1_uk_n148 ) , .B2( u1_uk_n1572 ) , .A2( u1_uk_n1613 ) , .A1( u1_uk_n202 ) );
  OAI22_X1 u1_uk_U247 (.ZN( u1_K14_39 ) , .A1( u1_uk_n148 ) , .B2( u1_uk_n1832 ) , .A2( u1_uk_n1836 ) , .B1( u1_uk_n231 ) );
  INV_X1 u1_uk_U25 (.ZN( u1_uk_n146 ) , .A( u1_uk_n251 ) );
  OAI22_X1 u1_uk_U266 (.ZN( u1_K14_48 ) , .B1( u1_uk_n148 ) , .B2( u1_uk_n1798 ) , .A2( u1_uk_n1836 ) , .A1( u1_uk_n297 ) );
  OAI22_X1 u1_uk_U273 (.ZN( u1_K11_44 ) , .B1( u1_uk_n102 ) , .B2( u1_uk_n1683 ) , .A2( u1_uk_n1703 ) , .A1( u1_uk_n257 ) );
  OAI22_X1 u1_uk_U301 (.ZN( u1_K12_8 ) , .B2( u1_uk_n1731 ) , .A2( u1_uk_n1752 ) , .A1( u1_uk_n230 ) , .B1( u1_uk_n99 ) );
  OAI22_X1 u1_uk_U311 (.ZN( u1_K7_26 ) , .A1( u1_uk_n141 ) , .B2( u1_uk_n1500 ) , .A2( u1_uk_n1520 ) , .B1( u1_uk_n230 ) );
  OAI21_X1 u1_uk_U323 (.ZN( u1_K11_26 ) , .B1( u1_uk_n161 ) , .B2( u1_uk_n1695 ) , .A( u1_uk_n409 ) );
  NAND2_X1 u1_uk_U324 (.A1( u1_uk_K_r9_35 ) , .A2( u1_uk_n11 ) , .ZN( u1_uk_n409 ) );
  OAI21_X1 u1_uk_U325 (.ZN( u1_K13_26 ) , .B1( u1_uk_n148 ) , .B2( u1_uk_n1765 ) , .A( u1_uk_n694 ) );
  NAND2_X1 u1_uk_U326 (.A1( u1_uk_K_r11_7 ) , .A2( u1_uk_n31 ) , .ZN( u1_uk_n694 ) );
  INV_X1 u1_uk_U33 (.ZN( u1_uk_n161 ) , .A( u1_uk_n230 ) );
  BUF_X1 u1_uk_U36 (.Z( u1_uk_n230 ) , .A( u1_uk_n277 ) );
  INV_X1 u1_uk_U365 (.ZN( u1_K11_46 ) , .A( u1_uk_n468 ) );
  AOI22_X1 u1_uk_U366 (.B2( u1_uk_K_r9_45 ) , .A2( u1_uk_K_r9_9 ) , .A1( u1_uk_n164 ) , .B1( u1_uk_n292 ) , .ZN( u1_uk_n468 ) );
  OAI22_X1 u1_uk_U374 (.ZN( u1_K8_40 ) , .B2( u1_uk_n1555 ) , .A2( u1_uk_n1561 ) , .A1( u1_uk_n250 ) , .B1( u1_uk_n63 ) );
  OAI22_X1 u1_uk_U385 (.ZN( u1_K11_28 ) , .A1( u1_uk_n129 ) , .B2( u1_uk_n1672 ) , .A2( u1_uk_n1704 ) , .B1( u1_uk_n298 ) );
  OAI22_X1 u1_uk_U394 (.ZN( u1_K7_28 ) , .B2( u1_uk_n1501 ) , .A2( u1_uk_n1510 ) , .A1( u1_uk_n251 ) , .B1( u1_uk_n92 ) );
  OAI22_X1 u1_uk_U421 (.ZN( u1_K12_9 ) , .A1( u1_uk_n10 ) , .B2( u1_uk_n1745 ) , .A2( u1_uk_n1752 ) , .B1( u1_uk_n207 ) );
  OAI22_X1 u1_uk_U438 (.ZN( u1_K14_37 ) , .A1( u1_uk_n163 ) , .B2( u1_uk_n1815 ) , .A2( u1_uk_n1821 ) , .B1( u1_uk_n230 ) );
  INV_X1 u1_uk_U443 (.ZN( u1_K8_37 ) , .A( u1_uk_n1138 ) );
  AOI22_X1 u1_uk_U444 (.B2( u1_uk_K_r6_14 ) , .A2( u1_uk_K_r6_7 ) , .ZN( u1_uk_n1138 ) , .B1( u1_uk_n163 ) , .A1( u1_uk_n203 ) );
  OAI22_X1 u1_uk_U457 (.ZN( u1_K13_33 ) , .A1( u1_uk_n129 ) , .B2( u1_uk_n1753 ) , .A2( u1_uk_n1758 ) , .B1( u1_uk_n188 ) );
  INV_X1 u1_uk_U461 (.ZN( u1_K9_33 ) , .A( u1_uk_n1162 ) );
  AOI22_X1 u1_uk_U462 (.B2( u1_uk_K_r7_1 ) , .A2( u1_uk_K_r7_8 ) , .ZN( u1_uk_n1162 ) , .B1( u1_uk_n162 ) , .A1( u1_uk_n286 ) );
  OAI21_X1 u1_uk_U475 (.ZN( u1_K9_37 ) , .A( u1_uk_n1164 ) , .B2( u1_uk_n1581 ) , .B1( u1_uk_n92 ) );
  NAND2_X1 u1_uk_U476 (.A1( u1_uk_K_r7_7 ) , .A2( u1_uk_n102 ) , .ZN( u1_uk_n1164 ) );
  OAI22_X1 u1_uk_U485 (.ZN( u1_K13_29 ) , .A1( u1_uk_n145 ) , .B2( u1_uk_n1772 ) , .A2( u1_uk_n1775 ) , .B1( u1_uk_n188 ) );
  OAI21_X1 u1_uk_U486 (.ZN( u1_K11_29 ) , .B1( u1_uk_n161 ) , .B2( u1_uk_n1664 ) , .A( u1_uk_n415 ) );
  NAND2_X1 u1_uk_U487 (.A1( u1_uk_K_r9_0 ) , .A2( u1_uk_n11 ) , .ZN( u1_uk_n415 ) );
  BUF_X1 u1_uk_U49 (.Z( u1_uk_n231 ) , .A( u1_uk_n277 ) );
  OAI22_X1 u1_uk_U504 (.ZN( u1_K7_29 ) , .B2( u1_uk_n1489 ) , .A2( u1_uk_n1520 ) , .A1( u1_uk_n208 ) , .B1( u1_uk_n92 ) );
  BUF_X1 u1_uk_U53 (.Z( u1_uk_n188 ) , .A( u1_uk_n292 ) );
  OAI21_X1 u1_uk_U531 (.ZN( u1_K12_12 ) , .B2( u1_uk_n1719 ) , .A( u1_uk_n503 ) , .B1( u1_uk_n63 ) );
  NAND2_X1 u1_uk_U532 (.A1( u1_uk_K_r10_11 ) , .A2( u1_uk_n27 ) , .ZN( u1_uk_n503 ) );
  BUF_X1 u1_uk_U55 (.Z( u1_uk_n251 ) , .A( u1_uk_n257 ) );
  OAI22_X1 u1_uk_U550 (.ZN( u1_K9_36 ) , .A1( u1_uk_n117 ) , .B2( u1_uk_n1599 ) , .A2( u1_uk_n1605 ) , .B1( u1_uk_n291 ) );
  OAI22_X1 u1_uk_U558 (.ZN( u1_K13_36 ) , .A1( u1_uk_n146 ) , .B2( u1_uk_n1777 ) , .A2( u1_uk_n1783 ) , .B1( u1_uk_n251 ) );
  BUF_X1 u1_uk_U56 (.A( u1_uk_n251 ) , .Z( u1_uk_n252 ) );
  OAI22_X1 u1_uk_U565 (.ZN( u1_K9_38 ) , .B2( u1_uk_n1605 ) , .A2( u1_uk_n1612 ) , .B1( u1_uk_n214 ) , .A1( u1_uk_n92 ) );
  INV_X1 u1_uk_U6 (.ZN( u1_uk_n182 ) , .A( u1_uk_n223 ) );
  INV_X1 u1_uk_U601 (.ZN( u1_K11_22 ) , .A( u1_uk_n407 ) );
  AOI22_X1 u1_uk_U602 (.B2( u1_uk_K_r9_13 ) , .A2( u1_uk_K_r9_19 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n230 ) , .ZN( u1_uk_n407 ) );
  OAI22_X1 u1_uk_U618 (.ZN( u1_K13_35 ) , .A1( u1_uk_n146 ) , .B2( u1_uk_n1764 ) , .A2( u1_uk_n1793 ) , .B1( u1_uk_n223 ) );
  INV_X1 u1_uk_U624 (.ZN( u1_K9_35 ) , .A( u1_uk_n1163 ) );
  AOI22_X1 u1_uk_U625 (.B2( u1_uk_K_r7_16 ) , .A2( u1_uk_K_r7_23 ) , .ZN( u1_uk_n1163 ) , .B1( u1_uk_n129 ) , .A1( u1_uk_n292 ) );
  BUF_X1 u1_uk_U63 (.Z( u1_uk_n257 ) , .A( u1_uk_n292 ) );
  OAI22_X1 u1_uk_U655 (.ZN( u1_K14_43 ) , .A1( u1_uk_n146 ) , .B2( u1_uk_n1829 ) , .A2( u1_uk_n1832 ) , .B1( u1_uk_n231 ) );
  OAI21_X1 u1_uk_U669 (.ZN( u1_K14_45 ) , .B2( u1_uk_n1830 ) , .B1( u1_uk_n251 ) , .A( u1_uk_n960 ) );
  NAND2_X1 u1_uk_U670 (.A1( u1_uk_K_r12_16 ) , .A2( u1_uk_n292 ) , .ZN( u1_uk_n960 ) );
  OAI22_X1 u1_uk_U675 (.ZN( u1_K11_43 ) , .B1( u1_uk_n146 ) , .B2( u1_uk_n1662 ) , .A2( u1_uk_n1704 ) , .A1( u1_uk_n298 ) );
  OAI21_X1 u1_uk_U684 (.ZN( u1_K12_7 ) , .B1( u1_uk_n161 ) , .B2( u1_uk_n1750 ) , .A( u1_uk_n665 ) );
  NAND2_X1 u1_uk_U685 (.A1( u1_uk_K_r10_19 ) , .A2( u1_uk_n11 ) , .ZN( u1_uk_n665 ) );
  OAI22_X1 u1_uk_U690 (.ZN( u1_K11_25 ) , .B1( u1_uk_n109 ) , .B2( u1_uk_n1677 ) , .A2( u1_uk_n1696 ) , .A1( u1_uk_n213 ) );
  OAI22_X1 u1_uk_U691 (.ZN( u1_K13_25 ) , .A1( u1_uk_n147 ) , .B2( u1_uk_n1765 ) , .A2( u1_uk_n1790 ) , .B1( u1_uk_n191 ) );
  INV_X1 u1_uk_U7 (.ZN( u1_uk_n102 ) , .A( u1_uk_n230 ) );
  OAI22_X1 u1_uk_U726 (.ZN( u1_K13_32 ) , .B1( u1_uk_n100 ) , .A2( u1_uk_n1758 ) , .B2( u1_uk_n1782 ) , .A1( u1_uk_n291 ) );
  OAI22_X1 u1_uk_U731 (.ZN( u1_K9_32 ) , .A1( u1_uk_n117 ) , .B2( u1_uk_n1601 ) , .A2( u1_uk_n1608 ) , .B1( u1_uk_n257 ) );
  OAI22_X1 u1_uk_U733 (.ZN( u1_K14_42 ) , .A1( u1_uk_n145 ) , .B2( u1_uk_n1798 ) , .A2( u1_uk_n1829 ) , .B1( u1_uk_n231 ) );
  INV_X1 u1_uk_U742 (.ZN( u1_K9_42 ) , .A( u1_uk_n1167 ) );
  AOI22_X1 u1_uk_U743 (.B2( u1_uk_K_r7_15 ) , .A2( u1_uk_K_r7_22 ) , .ZN( u1_uk_n1167 ) , .B1( u1_uk_n162 ) , .A1( u1_uk_n291 ) );
  OAI22_X1 u1_uk_U763 (.ZN( u1_K11_27 ) , .A1( u1_uk_n129 ) , .B2( u1_uk_n1684 ) , .A2( u1_uk_n1690 ) , .B1( u1_uk_n279 ) );
  OAI22_X1 u1_uk_U764 (.ZN( u1_K13_27 ) , .A1( u1_uk_n117 ) , .B2( u1_uk_n1754 ) , .A2( u1_uk_n1777 ) , .B1( u1_uk_n191 ) );
  OAI21_X1 u1_uk_U766 (.ZN( u1_K11_21 ) , .B1( u1_uk_n161 ) , .B2( u1_uk_n1667 ) , .A( u1_uk_n395 ) );
  NAND2_X1 u1_uk_U767 (.A1( u1_uk_K_r9_5 ) , .A2( u1_uk_n11 ) , .ZN( u1_uk_n395 ) );
  INV_X1 u1_uk_U796 (.ZN( u1_K7_27 ) , .A( u1_uk_n1115 ) );
  AOI22_X1 u1_uk_U797 (.B2( u1_uk_K_r5_23 ) , .A2( u1_uk_K_r5_43 ) , .ZN( u1_uk_n1115 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n203 ) );
  INV_X1 u1_uk_U835 (.ZN( u1_K11_20 ) , .A( u1_uk_n391 ) );
  AOI22_X1 u1_uk_U836 (.B2( u1_uk_K_r9_10 ) , .A2( u1_uk_K_r9_4 ) , .A1( u1_uk_n100 ) , .B1( u1_uk_n292 ) , .ZN( u1_uk_n391 ) );
  OAI22_X1 u1_uk_U875 (.ZN( u1_K13_34 ) , .B1( u1_uk_n100 ) , .B2( u1_uk_n1768 ) , .A2( u1_uk_n1784 ) , .A1( u1_uk_n294 ) );
  OAI21_X1 u1_uk_U88 (.ZN( u1_K11_23 ) , .B2( u1_uk_n1698 ) , .B1( u1_uk_n292 ) , .A( u1_uk_n408 ) );
  OAI22_X1 u1_uk_U880 (.ZN( u1_K12_10 ) , .B1( u1_uk_n118 ) , .B2( u1_uk_n1718 ) , .A2( u1_uk_n1739 ) , .A1( u1_uk_n207 ) );
  OAI22_X1 u1_uk_U881 (.ZN( u1_K12_11 ) , .B1( u1_uk_n102 ) , .A2( u1_uk_n1713 ) , .B2( u1_uk_n1739 ) , .A1( u1_uk_n279 ) );
  NAND2_X1 u1_uk_U89 (.A1( u1_uk_K_r9_27 ) , .A2( u1_uk_n298 ) , .ZN( u1_uk_n408 ) );
  OAI22_X1 u1_uk_U910 (.ZN( u1_K7_30 ) , .B2( u1_uk_n1490 ) , .A2( u1_uk_n1521 ) , .A1( u1_uk_n213 ) , .B1( u1_uk_n92 ) );
  OAI22_X1 u1_uk_U920 (.ZN( u1_K8_38 ) , .B1( u1_uk_n145 ) , .B2( u1_uk_n1560 ) , .A2( u1_uk_n1566 ) , .A1( u1_uk_n202 ) );
  OAI22_X1 u1_uk_U933 (.ZN( u1_K11_48 ) , .A1( u1_uk_n128 ) , .B2( u1_uk_n1689 ) , .A2( u1_uk_n1696 ) , .B1( u1_uk_n223 ) );
  OAI22_X1 u1_uk_U941 (.ZN( u1_K11_24 ) , .A1( u1_uk_n129 ) , .B2( u1_uk_n1682 ) , .A2( u1_uk_n1687 ) , .B1( u1_uk_n231 ) );
  OAI22_X1 u1_uk_U946 (.ZN( u1_K14_47 ) , .A1( u1_uk_n146 ) , .B2( u1_uk_n1820 ) , .A2( u1_uk_n1830 ) , .B1( u1_uk_n238 ) );
  OAI22_X1 u1_uk_U949 (.ZN( u1_K9_34 ) , .A1( u1_uk_n117 ) , .B2( u1_uk_n1581 ) , .A2( u1_uk_n1588 ) , .B1( u1_uk_n286 ) );
  OAI22_X1 u1_uk_U966 (.ZN( u1_K14_38 ) , .A2( u1_uk_n1807 ) , .B2( u1_uk_n1823 ) , .B1( u1_uk_n230 ) , .A1( u1_uk_n94 ) );
  INV_X1 u1_uk_U97 (.ZN( u1_K9_41 ) , .A( u1_uk_n1166 ) );
  OAI22_X1 u1_uk_U971 (.ZN( u1_K9_40 ) , .B2( u1_uk_n1600 ) , .A2( u1_uk_n1606 ) , .A1( u1_uk_n17 ) , .B1( u1_uk_n231 ) );
  OAI22_X1 u1_uk_U975 (.ZN( u1_K11_45 ) , .A1( u1_uk_n161 ) , .B2( u1_uk_n1677 ) , .A2( u1_uk_n1684 ) , .B1( u1_uk_n231 ) );
  AOI22_X1 u1_uk_U98 (.B2( u1_uk_K_r7_23 ) , .A2( u1_uk_K_r7_30 ) , .ZN( u1_uk_n1166 ) , .B1( u1_uk_n162 ) , .A1( u1_uk_n252 ) );
  XOR2_X1 u2_U243 (.B( u2_L8_26 ) , .Z( u2_N313 ) , .A( u2_out9_26 ) );
  XOR2_X1 u2_U250 (.B( u2_L8_20 ) , .Z( u2_N307 ) , .A( u2_out9_20 ) );
  XOR2_X1 u2_U262 (.B( u2_L8_10 ) , .Z( u2_N297 ) , .A( u2_out9_10 ) );
  XOR2_X1 u2_U272 (.B( u2_L8_1 ) , .Z( u2_N288 ) , .A( u2_out9_1 ) );
  XOR2_X1 u2_u9_U33 (.B( u2_K10_24 ) , .A( u2_R8_17 ) , .Z( u2_u9_X_24 ) );
  XOR2_X1 u2_u9_U34 (.B( u2_K10_23 ) , .A( u2_R8_16 ) , .Z( u2_u9_X_23 ) );
  XOR2_X1 u2_u9_U35 (.B( u2_K10_22 ) , .A( u2_R8_15 ) , .Z( u2_u9_X_22 ) );
  XOR2_X1 u2_u9_U36 (.B( u2_K10_21 ) , .A( u2_R8_14 ) , .Z( u2_u9_X_21 ) );
  XOR2_X1 u2_u9_U37 (.B( u2_K10_20 ) , .A( u2_R8_13 ) , .Z( u2_u9_X_20 ) );
  XOR2_X1 u2_u9_U39 (.B( u2_K10_19 ) , .A( u2_R8_12 ) , .Z( u2_u9_X_19 ) );
  OAI22_X1 u2_u9_u3_U10 (.B1( u2_u9_u3_n113 ) , .A2( u2_u9_u3_n135 ) , .A1( u2_u9_u3_n150 ) , .B2( u2_u9_u3_n164 ) , .ZN( u2_u9_u3_n98 ) );
  OAI211_X1 u2_u9_u3_U11 (.B( u2_u9_u3_n106 ) , .ZN( u2_u9_u3_n119 ) , .C2( u2_u9_u3_n128 ) , .C1( u2_u9_u3_n167 ) , .A( u2_u9_u3_n181 ) );
  AOI221_X1 u2_u9_u3_U12 (.C1( u2_u9_u3_n105 ) , .ZN( u2_u9_u3_n106 ) , .A( u2_u9_u3_n131 ) , .B2( u2_u9_u3_n132 ) , .C2( u2_u9_u3_n133 ) , .B1( u2_u9_u3_n169 ) );
  INV_X1 u2_u9_u3_U13 (.ZN( u2_u9_u3_n181 ) , .A( u2_u9_u3_n98 ) );
  NAND2_X1 u2_u9_u3_U14 (.ZN( u2_u9_u3_n105 ) , .A2( u2_u9_u3_n130 ) , .A1( u2_u9_u3_n155 ) );
  AOI22_X1 u2_u9_u3_U15 (.B1( u2_u9_u3_n115 ) , .A2( u2_u9_u3_n116 ) , .ZN( u2_u9_u3_n123 ) , .B2( u2_u9_u3_n133 ) , .A1( u2_u9_u3_n169 ) );
  NAND2_X1 u2_u9_u3_U16 (.ZN( u2_u9_u3_n116 ) , .A2( u2_u9_u3_n151 ) , .A1( u2_u9_u3_n182 ) );
  NOR2_X1 u2_u9_u3_U17 (.ZN( u2_u9_u3_n126 ) , .A2( u2_u9_u3_n150 ) , .A1( u2_u9_u3_n164 ) );
  AOI21_X1 u2_u9_u3_U18 (.ZN( u2_u9_u3_n112 ) , .B2( u2_u9_u3_n146 ) , .B1( u2_u9_u3_n155 ) , .A( u2_u9_u3_n167 ) );
  NAND2_X1 u2_u9_u3_U19 (.A1( u2_u9_u3_n135 ) , .ZN( u2_u9_u3_n142 ) , .A2( u2_u9_u3_n164 ) );
  NAND2_X1 u2_u9_u3_U20 (.ZN( u2_u9_u3_n132 ) , .A2( u2_u9_u3_n152 ) , .A1( u2_u9_u3_n156 ) );
  AND2_X1 u2_u9_u3_U21 (.A2( u2_u9_u3_n113 ) , .A1( u2_u9_u3_n114 ) , .ZN( u2_u9_u3_n151 ) );
  INV_X1 u2_u9_u3_U22 (.A( u2_u9_u3_n133 ) , .ZN( u2_u9_u3_n165 ) );
  INV_X1 u2_u9_u3_U23 (.A( u2_u9_u3_n135 ) , .ZN( u2_u9_u3_n170 ) );
  NAND2_X1 u2_u9_u3_U24 (.A1( u2_u9_u3_n107 ) , .A2( u2_u9_u3_n108 ) , .ZN( u2_u9_u3_n140 ) );
  NAND2_X1 u2_u9_u3_U25 (.ZN( u2_u9_u3_n117 ) , .A1( u2_u9_u3_n124 ) , .A2( u2_u9_u3_n148 ) );
  NAND2_X1 u2_u9_u3_U26 (.ZN( u2_u9_u3_n143 ) , .A1( u2_u9_u3_n165 ) , .A2( u2_u9_u3_n167 ) );
  INV_X1 u2_u9_u3_U27 (.A( u2_u9_u3_n130 ) , .ZN( u2_u9_u3_n177 ) );
  INV_X1 u2_u9_u3_U28 (.A( u2_u9_u3_n128 ) , .ZN( u2_u9_u3_n176 ) );
  INV_X1 u2_u9_u3_U29 (.A( u2_u9_u3_n155 ) , .ZN( u2_u9_u3_n174 ) );
  INV_X1 u2_u9_u3_U3 (.A( u2_u9_u3_n129 ) , .ZN( u2_u9_u3_n183 ) );
  INV_X1 u2_u9_u3_U30 (.A( u2_u9_u3_n139 ) , .ZN( u2_u9_u3_n185 ) );
  NOR2_X1 u2_u9_u3_U31 (.ZN( u2_u9_u3_n135 ) , .A2( u2_u9_u3_n141 ) , .A1( u2_u9_u3_n169 ) );
  OAI222_X1 u2_u9_u3_U32 (.C2( u2_u9_u3_n107 ) , .A2( u2_u9_u3_n108 ) , .B1( u2_u9_u3_n135 ) , .ZN( u2_u9_u3_n138 ) , .B2( u2_u9_u3_n146 ) , .C1( u2_u9_u3_n154 ) , .A1( u2_u9_u3_n164 ) );
  NOR4_X1 u2_u9_u3_U33 (.A4( u2_u9_u3_n157 ) , .A3( u2_u9_u3_n158 ) , .A2( u2_u9_u3_n159 ) , .A1( u2_u9_u3_n160 ) , .ZN( u2_u9_u3_n161 ) );
  AOI21_X1 u2_u9_u3_U34 (.B2( u2_u9_u3_n152 ) , .B1( u2_u9_u3_n153 ) , .ZN( u2_u9_u3_n158 ) , .A( u2_u9_u3_n164 ) );
  AOI21_X1 u2_u9_u3_U35 (.A( u2_u9_u3_n154 ) , .B2( u2_u9_u3_n155 ) , .B1( u2_u9_u3_n156 ) , .ZN( u2_u9_u3_n157 ) );
  AOI21_X1 u2_u9_u3_U36 (.A( u2_u9_u3_n149 ) , .B2( u2_u9_u3_n150 ) , .B1( u2_u9_u3_n151 ) , .ZN( u2_u9_u3_n159 ) );
  AOI211_X1 u2_u9_u3_U37 (.ZN( u2_u9_u3_n109 ) , .A( u2_u9_u3_n119 ) , .C2( u2_u9_u3_n129 ) , .B( u2_u9_u3_n138 ) , .C1( u2_u9_u3_n141 ) );
  AOI211_X1 u2_u9_u3_U38 (.B( u2_u9_u3_n119 ) , .A( u2_u9_u3_n120 ) , .C2( u2_u9_u3_n121 ) , .ZN( u2_u9_u3_n122 ) , .C1( u2_u9_u3_n179 ) );
  INV_X1 u2_u9_u3_U39 (.A( u2_u9_u3_n156 ) , .ZN( u2_u9_u3_n179 ) );
  INV_X1 u2_u9_u3_U4 (.A( u2_u9_u3_n140 ) , .ZN( u2_u9_u3_n182 ) );
  OAI22_X1 u2_u9_u3_U40 (.B1( u2_u9_u3_n118 ) , .ZN( u2_u9_u3_n120 ) , .A1( u2_u9_u3_n135 ) , .B2( u2_u9_u3_n154 ) , .A2( u2_u9_u3_n178 ) );
  AND3_X1 u2_u9_u3_U41 (.ZN( u2_u9_u3_n118 ) , .A2( u2_u9_u3_n124 ) , .A1( u2_u9_u3_n144 ) , .A3( u2_u9_u3_n152 ) );
  INV_X1 u2_u9_u3_U42 (.A( u2_u9_u3_n121 ) , .ZN( u2_u9_u3_n164 ) );
  NAND2_X1 u2_u9_u3_U43 (.ZN( u2_u9_u3_n133 ) , .A1( u2_u9_u3_n154 ) , .A2( u2_u9_u3_n164 ) );
  OAI211_X1 u2_u9_u3_U44 (.B( u2_u9_u3_n127 ) , .ZN( u2_u9_u3_n139 ) , .C1( u2_u9_u3_n150 ) , .C2( u2_u9_u3_n154 ) , .A( u2_u9_u3_n184 ) );
  INV_X1 u2_u9_u3_U45 (.A( u2_u9_u3_n125 ) , .ZN( u2_u9_u3_n184 ) );
  AOI221_X1 u2_u9_u3_U46 (.A( u2_u9_u3_n126 ) , .ZN( u2_u9_u3_n127 ) , .C2( u2_u9_u3_n132 ) , .C1( u2_u9_u3_n169 ) , .B2( u2_u9_u3_n170 ) , .B1( u2_u9_u3_n174 ) );
  OAI22_X1 u2_u9_u3_U47 (.A1( u2_u9_u3_n124 ) , .ZN( u2_u9_u3_n125 ) , .B2( u2_u9_u3_n145 ) , .A2( u2_u9_u3_n165 ) , .B1( u2_u9_u3_n167 ) );
  NOR2_X1 u2_u9_u3_U48 (.A1( u2_u9_u3_n113 ) , .ZN( u2_u9_u3_n131 ) , .A2( u2_u9_u3_n154 ) );
  NAND2_X1 u2_u9_u3_U49 (.A1( u2_u9_u3_n103 ) , .ZN( u2_u9_u3_n150 ) , .A2( u2_u9_u3_n99 ) );
  INV_X1 u2_u9_u3_U5 (.A( u2_u9_u3_n117 ) , .ZN( u2_u9_u3_n178 ) );
  NAND2_X1 u2_u9_u3_U50 (.A2( u2_u9_u3_n102 ) , .ZN( u2_u9_u3_n155 ) , .A1( u2_u9_u3_n97 ) );
  INV_X1 u2_u9_u3_U51 (.A( u2_u9_u3_n141 ) , .ZN( u2_u9_u3_n167 ) );
  AOI21_X1 u2_u9_u3_U52 (.B2( u2_u9_u3_n114 ) , .B1( u2_u9_u3_n146 ) , .A( u2_u9_u3_n154 ) , .ZN( u2_u9_u3_n94 ) );
  AOI21_X1 u2_u9_u3_U53 (.ZN( u2_u9_u3_n110 ) , .B2( u2_u9_u3_n142 ) , .B1( u2_u9_u3_n186 ) , .A( u2_u9_u3_n95 ) );
  INV_X1 u2_u9_u3_U54 (.A( u2_u9_u3_n145 ) , .ZN( u2_u9_u3_n186 ) );
  AOI21_X1 u2_u9_u3_U55 (.B1( u2_u9_u3_n124 ) , .A( u2_u9_u3_n149 ) , .B2( u2_u9_u3_n155 ) , .ZN( u2_u9_u3_n95 ) );
  INV_X1 u2_u9_u3_U56 (.A( u2_u9_u3_n149 ) , .ZN( u2_u9_u3_n169 ) );
  NAND2_X1 u2_u9_u3_U57 (.ZN( u2_u9_u3_n124 ) , .A1( u2_u9_u3_n96 ) , .A2( u2_u9_u3_n97 ) );
  NAND2_X1 u2_u9_u3_U58 (.A2( u2_u9_u3_n100 ) , .ZN( u2_u9_u3_n146 ) , .A1( u2_u9_u3_n96 ) );
  NAND2_X1 u2_u9_u3_U59 (.A1( u2_u9_u3_n101 ) , .ZN( u2_u9_u3_n145 ) , .A2( u2_u9_u3_n99 ) );
  AOI221_X1 u2_u9_u3_U6 (.A( u2_u9_u3_n131 ) , .C2( u2_u9_u3_n132 ) , .C1( u2_u9_u3_n133 ) , .ZN( u2_u9_u3_n134 ) , .B1( u2_u9_u3_n143 ) , .B2( u2_u9_u3_n177 ) );
  NAND2_X1 u2_u9_u3_U60 (.A1( u2_u9_u3_n100 ) , .ZN( u2_u9_u3_n156 ) , .A2( u2_u9_u3_n99 ) );
  NAND2_X1 u2_u9_u3_U61 (.A2( u2_u9_u3_n101 ) , .A1( u2_u9_u3_n104 ) , .ZN( u2_u9_u3_n148 ) );
  NAND2_X1 u2_u9_u3_U62 (.A1( u2_u9_u3_n100 ) , .A2( u2_u9_u3_n102 ) , .ZN( u2_u9_u3_n128 ) );
  NAND2_X1 u2_u9_u3_U63 (.A2( u2_u9_u3_n101 ) , .A1( u2_u9_u3_n102 ) , .ZN( u2_u9_u3_n152 ) );
  NAND2_X1 u2_u9_u3_U64 (.A2( u2_u9_u3_n101 ) , .ZN( u2_u9_u3_n114 ) , .A1( u2_u9_u3_n96 ) );
  NAND2_X1 u2_u9_u3_U65 (.ZN( u2_u9_u3_n107 ) , .A1( u2_u9_u3_n97 ) , .A2( u2_u9_u3_n99 ) );
  NAND2_X1 u2_u9_u3_U66 (.A2( u2_u9_u3_n100 ) , .A1( u2_u9_u3_n104 ) , .ZN( u2_u9_u3_n113 ) );
  NAND2_X1 u2_u9_u3_U67 (.A1( u2_u9_u3_n104 ) , .ZN( u2_u9_u3_n153 ) , .A2( u2_u9_u3_n97 ) );
  NAND2_X1 u2_u9_u3_U68 (.A2( u2_u9_u3_n103 ) , .A1( u2_u9_u3_n104 ) , .ZN( u2_u9_u3_n130 ) );
  NAND2_X1 u2_u9_u3_U69 (.A2( u2_u9_u3_n103 ) , .ZN( u2_u9_u3_n144 ) , .A1( u2_u9_u3_n96 ) );
  OAI22_X1 u2_u9_u3_U7 (.B2( u2_u9_u3_n147 ) , .A2( u2_u9_u3_n148 ) , .ZN( u2_u9_u3_n160 ) , .B1( u2_u9_u3_n165 ) , .A1( u2_u9_u3_n168 ) );
  NAND2_X1 u2_u9_u3_U70 (.A1( u2_u9_u3_n102 ) , .A2( u2_u9_u3_n103 ) , .ZN( u2_u9_u3_n108 ) );
  NOR2_X1 u2_u9_u3_U71 (.A2( u2_u9_X_19 ) , .A1( u2_u9_X_20 ) , .ZN( u2_u9_u3_n99 ) );
  NOR2_X1 u2_u9_u3_U72 (.A2( u2_u9_X_21 ) , .A1( u2_u9_X_24 ) , .ZN( u2_u9_u3_n103 ) );
  NOR2_X1 u2_u9_u3_U73 (.A2( u2_u9_X_24 ) , .A1( u2_u9_u3_n171 ) , .ZN( u2_u9_u3_n97 ) );
  NOR2_X1 u2_u9_u3_U74 (.A2( u2_u9_X_23 ) , .ZN( u2_u9_u3_n141 ) , .A1( u2_u9_u3_n166 ) );
  NOR2_X1 u2_u9_u3_U75 (.A2( u2_u9_X_19 ) , .A1( u2_u9_u3_n172 ) , .ZN( u2_u9_u3_n96 ) );
  NAND2_X1 u2_u9_u3_U76 (.A1( u2_u9_X_22 ) , .A2( u2_u9_X_23 ) , .ZN( u2_u9_u3_n154 ) );
  NAND2_X1 u2_u9_u3_U77 (.A1( u2_u9_X_23 ) , .ZN( u2_u9_u3_n149 ) , .A2( u2_u9_u3_n166 ) );
  NOR2_X1 u2_u9_u3_U78 (.A2( u2_u9_X_22 ) , .A1( u2_u9_X_23 ) , .ZN( u2_u9_u3_n121 ) );
  AND2_X1 u2_u9_u3_U79 (.A1( u2_u9_X_24 ) , .ZN( u2_u9_u3_n101 ) , .A2( u2_u9_u3_n171 ) );
  AND3_X1 u2_u9_u3_U8 (.A3( u2_u9_u3_n144 ) , .A2( u2_u9_u3_n145 ) , .A1( u2_u9_u3_n146 ) , .ZN( u2_u9_u3_n147 ) );
  AND2_X1 u2_u9_u3_U80 (.A1( u2_u9_X_19 ) , .ZN( u2_u9_u3_n102 ) , .A2( u2_u9_u3_n172 ) );
  AND2_X1 u2_u9_u3_U81 (.A1( u2_u9_X_21 ) , .A2( u2_u9_X_24 ) , .ZN( u2_u9_u3_n100 ) );
  AND2_X1 u2_u9_u3_U82 (.A2( u2_u9_X_19 ) , .A1( u2_u9_X_20 ) , .ZN( u2_u9_u3_n104 ) );
  INV_X1 u2_u9_u3_U83 (.A( u2_u9_X_22 ) , .ZN( u2_u9_u3_n166 ) );
  INV_X1 u2_u9_u3_U84 (.A( u2_u9_X_21 ) , .ZN( u2_u9_u3_n171 ) );
  INV_X1 u2_u9_u3_U85 (.A( u2_u9_X_20 ) , .ZN( u2_u9_u3_n172 ) );
  OR4_X1 u2_u9_u3_U86 (.ZN( u2_out9_10 ) , .A4( u2_u9_u3_n136 ) , .A3( u2_u9_u3_n137 ) , .A1( u2_u9_u3_n138 ) , .A2( u2_u9_u3_n139 ) );
  OAI222_X1 u2_u9_u3_U87 (.C1( u2_u9_u3_n128 ) , .ZN( u2_u9_u3_n137 ) , .B1( u2_u9_u3_n148 ) , .A2( u2_u9_u3_n150 ) , .B2( u2_u9_u3_n154 ) , .C2( u2_u9_u3_n164 ) , .A1( u2_u9_u3_n167 ) );
  OAI221_X1 u2_u9_u3_U88 (.A( u2_u9_u3_n134 ) , .B2( u2_u9_u3_n135 ) , .ZN( u2_u9_u3_n136 ) , .C1( u2_u9_u3_n149 ) , .B1( u2_u9_u3_n151 ) , .C2( u2_u9_u3_n183 ) );
  NAND4_X1 u2_u9_u3_U89 (.ZN( u2_out9_26 ) , .A4( u2_u9_u3_n109 ) , .A3( u2_u9_u3_n110 ) , .A2( u2_u9_u3_n111 ) , .A1( u2_u9_u3_n173 ) );
  INV_X1 u2_u9_u3_U9 (.A( u2_u9_u3_n143 ) , .ZN( u2_u9_u3_n168 ) );
  INV_X1 u2_u9_u3_U90 (.ZN( u2_u9_u3_n173 ) , .A( u2_u9_u3_n94 ) );
  OAI21_X1 u2_u9_u3_U91 (.ZN( u2_u9_u3_n111 ) , .B2( u2_u9_u3_n117 ) , .A( u2_u9_u3_n133 ) , .B1( u2_u9_u3_n176 ) );
  NAND4_X1 u2_u9_u3_U92 (.ZN( u2_out9_20 ) , .A4( u2_u9_u3_n122 ) , .A3( u2_u9_u3_n123 ) , .A1( u2_u9_u3_n175 ) , .A2( u2_u9_u3_n180 ) );
  INV_X1 u2_u9_u3_U93 (.A( u2_u9_u3_n126 ) , .ZN( u2_u9_u3_n180 ) );
  INV_X1 u2_u9_u3_U94 (.A( u2_u9_u3_n112 ) , .ZN( u2_u9_u3_n175 ) );
  NAND4_X1 u2_u9_u3_U95 (.ZN( u2_out9_1 ) , .A4( u2_u9_u3_n161 ) , .A3( u2_u9_u3_n162 ) , .A2( u2_u9_u3_n163 ) , .A1( u2_u9_u3_n185 ) );
  NAND2_X1 u2_u9_u3_U96 (.ZN( u2_u9_u3_n163 ) , .A2( u2_u9_u3_n170 ) , .A1( u2_u9_u3_n176 ) );
  AOI22_X1 u2_u9_u3_U97 (.B2( u2_u9_u3_n140 ) , .B1( u2_u9_u3_n141 ) , .A2( u2_u9_u3_n142 ) , .ZN( u2_u9_u3_n162 ) , .A1( u2_u9_u3_n177 ) );
  NAND3_X1 u2_u9_u3_U98 (.A1( u2_u9_u3_n114 ) , .ZN( u2_u9_u3_n115 ) , .A2( u2_u9_u3_n145 ) , .A3( u2_u9_u3_n153 ) );
  NAND3_X1 u2_u9_u3_U99 (.ZN( u2_u9_u3_n129 ) , .A2( u2_u9_u3_n144 ) , .A1( u2_u9_u3_n153 ) , .A3( u2_u9_u3_n182 ) );
  OAI21_X1 u2_uk_U1005 (.ZN( u2_K10_21 ) , .B1( u2_uk_n102 ) , .B2( u2_uk_n1630 ) , .A( u2_uk_n252 ) );
  NAND2_X1 u2_uk_U1006 (.A1( u2_uk_K_r8_19 ) , .A2( u2_uk_n10 ) , .ZN( u2_uk_n252 ) );
  OAI22_X1 u2_uk_U160 (.ZN( u2_K10_19 ) , .A1( u2_uk_n117 ) , .B2( u2_uk_n1603 ) , .A2( u2_uk_n1613 ) , .B1( u2_uk_n187 ) );
  OAI21_X1 u2_uk_U179 (.ZN( u2_K10_24 ) , .B1( u2_uk_n102 ) , .B2( u2_uk_n1599 ) , .A( u2_uk_n277 ) );
  NAND2_X1 u2_uk_U180 (.A1( u2_uk_K_r8_40 ) , .A2( u2_uk_n27 ) , .ZN( u2_uk_n277 ) );
  INV_X1 u2_uk_U593 (.ZN( u2_K10_22 ) , .A( u2_uk_n257 ) );
  OAI21_X1 u2_uk_U73 (.ZN( u2_K10_23 ) , .B2( u2_uk_n1590 ) , .B1( u2_uk_n187 ) , .A( u2_uk_n271 ) );
  NAND2_X1 u2_uk_U74 (.A1( u2_uk_K_r8_13 ) , .A2( u2_uk_n129 ) , .ZN( u2_uk_n271 ) );
  OAI22_X1 u2_uk_U940 (.ZN( u2_K10_20 ) , .A1( u2_uk_n118 ) , .B2( u2_uk_n1599 ) , .A2( u2_uk_n1629 ) , .B1( u2_uk_n182 ) );
endmodule

