module aes_aes_die_23 ( sa02_0, sa02_1, sa02_2, sa02_3, sa02_4, sa02_5, sa02_6, sa02_7, sa02_sr_0, sa02_sr_1, sa02_sr_2, sa02_sr_3, sa02_sr_4, sa02_sr_5, sa02_sr_6, sa02_sr_7 );
  input sa02_0, sa02_1, sa02_2, sa02_3, sa02_4, sa02_5, sa02_6, sa02_7;
  output sa02_sr_0, sa02_sr_1, sa02_sr_2, sa02_sr_3, sa02_sr_4, sa02_sr_5, sa02_sr_6, sa02_sr_7;
  wire us02_n438, us02_n439, us02_n440, us02_n441, us02_n442, us02_n443, us02_n444, us02_n445, us02_n446, 
       us02_n447, us02_n448, us02_n449, us02_n450, us02_n451, us02_n452, us02_n453, us02_n454, us02_n455, 
       us02_n456, us02_n457, us02_n458, us02_n459, us02_n460, us02_n461, us02_n462, us02_n463, us02_n464, 
       us02_n465, us02_n466, us02_n467, us02_n468, us02_n469, us02_n470, us02_n471, us02_n472, us02_n473, 
       us02_n474, us02_n475, us02_n476, us02_n477, us02_n478, us02_n479, us02_n480, us02_n481, us02_n482, 
       us02_n483, us02_n484, us02_n485, us02_n486, us02_n487, us02_n488, us02_n489, us02_n490, us02_n491, 
       us02_n492, us02_n493, us02_n494, us02_n495, us02_n496, us02_n497, us02_n498, us02_n499, us02_n500, 
       us02_n501, us02_n502, us02_n503, us02_n504, us02_n505, us02_n506, us02_n507, us02_n508, us02_n509, 
       us02_n510, us02_n511, us02_n512, us02_n513, us02_n514, us02_n515, us02_n516, us02_n517, us02_n518, 
       us02_n519, us02_n520, us02_n521, us02_n522, us02_n523, us02_n524, us02_n525, us02_n526, us02_n527, 
       us02_n528, us02_n529, us02_n530, us02_n531, us02_n532, us02_n533, us02_n534, us02_n535, us02_n536, 
       us02_n537, us02_n538, us02_n539, us02_n540, us02_n541, us02_n542, us02_n543, us02_n544, us02_n545, 
       us02_n546, us02_n547, us02_n548, us02_n549, us02_n550, us02_n551, us02_n552, us02_n553, us02_n554, 
       us02_n555, us02_n556, us02_n557, us02_n558, us02_n559, us02_n560, us02_n561, us02_n562, us02_n563, 
       us02_n564, us02_n565, us02_n566, us02_n567, us02_n568, us02_n569, us02_n570, us02_n571, us02_n572, 
       us02_n573, us02_n574, us02_n575, us02_n576, us02_n577, us02_n578, us02_n579, us02_n580, us02_n581, 
       us02_n582, us02_n583, us02_n584, us02_n585, us02_n586, us02_n587, us02_n588, us02_n589, us02_n590, 
       us02_n591, us02_n592, us02_n593, us02_n594, us02_n595, us02_n596, us02_n597, us02_n598, us02_n599, 
       us02_n600, us02_n601, us02_n602, us02_n603, us02_n604, us02_n605, us02_n606, us02_n607, us02_n608, 
       us02_n609, us02_n610, us02_n611, us02_n612, us02_n613, us02_n614, us02_n615, us02_n616, us02_n617, 
       us02_n618, us02_n619, us02_n620, us02_n621, us02_n622, us02_n623, us02_n624, us02_n625, us02_n626, 
       us02_n627, us02_n628, us02_n629, us02_n630, us02_n631, us02_n632, us02_n633, us02_n634, us02_n635, 
       us02_n636, us02_n637, us02_n638, us02_n639, us02_n640, us02_n641, us02_n642, us02_n643, us02_n644, 
       us02_n645, us02_n646, us02_n647, us02_n648, us02_n649, us02_n650, us02_n651, us02_n652, us02_n653, 
       us02_n654, us02_n655, us02_n656, us02_n657, us02_n658, us02_n659, us02_n660, us02_n661, us02_n662, 
       us02_n663, us02_n664, us02_n665, us02_n666, us02_n667, us02_n668, us02_n669, us02_n670, us02_n671, 
       us02_n672, us02_n673, us02_n674, us02_n675, us02_n676, us02_n677, us02_n678, us02_n679, us02_n680, 
       us02_n681, us02_n682, us02_n683, us02_n684, us02_n685, us02_n686, us02_n687, us02_n688, us02_n689, 
       us02_n690, us02_n691, us02_n692, us02_n693, us02_n694, us02_n695, us02_n696, us02_n697, us02_n698, 
       us02_n699, us02_n700, us02_n701, us02_n702, us02_n703, us02_n704, us02_n705, us02_n706, us02_n707, 
       us02_n708, us02_n709, us02_n710, us02_n711, us02_n712, us02_n713, us02_n714, us02_n715, us02_n716, 
       us02_n717, us02_n718, us02_n719, us02_n720, us02_n721, us02_n722, us02_n723, us02_n724, us02_n725, 
       us02_n726, us02_n727, us02_n728, us02_n729, us02_n730, us02_n731, us02_n732, us02_n733, us02_n734, 
       us02_n735, us02_n736, us02_n737, us02_n738, us02_n739, us02_n740, us02_n741, us02_n742, us02_n743, 
       us02_n744, us02_n745, us02_n746, us02_n747, us02_n748, us02_n749, us02_n750, us02_n751, us02_n752, 
       us02_n753, us02_n754, us02_n755, us02_n756, us02_n757, us02_n758, us02_n759, us02_n760, us02_n761, 
       us02_n762, us02_n763, us02_n764, us02_n765, us02_n766, us02_n767, us02_n768, us02_n769, us02_n770, 
       us02_n771, us02_n772, us02_n773, us02_n774, us02_n775, us02_n776, us02_n777, us02_n778, us02_n779, 
       us02_n780, us02_n781, us02_n782, us02_n783, us02_n784, us02_n785, us02_n786, us02_n787, us02_n788, 
       us02_n789, us02_n790, us02_n791, us02_n792, us02_n793, us02_n794, us02_n795, us02_n796, us02_n797, 
       us02_n798, us02_n799, us02_n800, us02_n801, us02_n802, us02_n803, us02_n804, us02_n805, us02_n806, 
       us02_n807, us02_n808, us02_n809, us02_n810, us02_n811, us02_n812, us02_n813, us02_n814, us02_n815, 
       us02_n816, us02_n817, us02_n818, us02_n819, us02_n820, us02_n821, us02_n822, us02_n823, us02_n824, 
       us02_n825, us02_n826, us02_n827, us02_n828, us02_n829, us02_n830, us02_n831, us02_n832, us02_n833, 
       us02_n834, us02_n835, us02_n836, us02_n837, us02_n838, us02_n839, us02_n840, us02_n841, us02_n842, 
       us02_n843, us02_n844, us02_n845, us02_n846, us02_n847, us02_n848, us02_n849, us02_n850, us02_n851, 
       us02_n852, us02_n853, us02_n854, us02_n855, us02_n856, us02_n857, us02_n858, us02_n859, us02_n860, 
       us02_n861, us02_n862, us02_n863, us02_n864, us02_n865, us02_n866, us02_n867, us02_n868, us02_n869, 
       us02_n870, us02_n871, us02_n872, us02_n873, us02_n874,  us02_n875;
  NOR2_X1 us02_U10 (.ZN( us02_n574 ) , .A1( us02_n621 ) , .A2( us02_n744 ) );
  NOR2_X1 us02_U100 (.ZN( us02_n685 ) , .A1( us02_n830 ) , .A2( us02_n831 ) );
  NOR4_X1 us02_U101 (.ZN( us02_n619 ) , .A1( us02_n655 ) , .A3( us02_n665 ) , .A4( us02_n681 ) , .A2( us02_n765 ) );
  NOR4_X1 us02_U102 (.A4( us02_n608 ) , .A3( us02_n609 ) , .A2( us02_n610 ) , .A1( us02_n611 ) , .ZN( us02_n618 ) );
  NOR4_X1 us02_U103 (.A4( us02_n613 ) , .A3( us02_n614 ) , .A2( us02_n615 ) , .A1( us02_n616 ) , .ZN( us02_n617 ) );
  NAND4_X1 us02_U104 (.A4( us02_n484 ) , .A3( us02_n485 ) , .A2( us02_n486 ) , .A1( us02_n487 ) , .ZN( us02_n777 ) );
  NOR4_X1 us02_U105 (.A4( us02_n483 ) , .ZN( us02_n486 ) , .A1( us02_n565 ) , .A2( us02_n580 ) , .A3( us02_n601 ) );
  NOR4_X1 us02_U106 (.ZN( us02_n485 ) , .A1( us02_n506 ) , .A2( us02_n518 ) , .A4( us02_n545 ) , .A3( us02_n610 ) );
  NOR4_X1 us02_U107 (.ZN( us02_n484 ) , .A2( us02_n532 ) , .A1( us02_n557 ) , .A3( us02_n630 ) , .A4( us02_n717 ) );
  NAND4_X1 us02_U108 (.A4( us02_n690 ) , .A3( us02_n691 ) , .A1( us02_n692 ) , .ZN( us02_n775 ) , .A2( us02_n871 ) );
  AOI221_X1 us02_U109 (.A( us02_n680 ) , .ZN( us02_n691 ) , .B2( us02_n839 ) , .C1( us02_n841 ) , .C2( us02_n861 ) , .B1( us02_n864 ) );
  NOR2_X1 us02_U11 (.A1( us02_n677 ) , .ZN( us02_n692 ) , .A2( us02_n806 ) );
  INV_X1 us02_U110 (.A( us02_n678 ) , .ZN( us02_n871 ) );
  NOR4_X1 us02_U111 (.A4( us02_n686 ) , .A3( us02_n687 ) , .A2( us02_n688 ) , .A1( us02_n689 ) , .ZN( us02_n690 ) );
  NAND4_X1 us02_U112 (.A4( us02_n559 ) , .A3( us02_n560 ) , .A2( us02_n561 ) , .A1( us02_n562 ) , .ZN( us02_n606 ) );
  NOR4_X1 us02_U113 (.ZN( us02_n560 ) , .A1( us02_n652 ) , .A3( us02_n660 ) , .A4( us02_n684 ) , .A2( us02_n767 ) );
  NOR4_X1 us02_U114 (.A4( us02_n551 ) , .A3( us02_n552 ) , .A2( us02_n553 ) , .A1( us02_n554 ) , .ZN( us02_n561 ) );
  NOR4_X1 us02_U115 (.A4( us02_n555 ) , .A3( us02_n556 ) , .A2( us02_n557 ) , .A1( us02_n558 ) , .ZN( us02_n559 ) );
  NAND4_X1 us02_U116 (.A4( us02_n718 ) , .A3( us02_n719 ) , .A2( us02_n720 ) , .ZN( us02_n740 ) , .A1( us02_n856 ) );
  INV_X1 us02_U117 (.A( us02_n708 ) , .ZN( us02_n856 ) );
  AOI221_X1 us02_U118 (.A( us02_n709 ) , .ZN( us02_n720 ) , .C2( us02_n843 ) , .B2( us02_n844 ) , .C1( us02_n860 ) , .B1( us02_n861 ) );
  NOR4_X1 us02_U119 (.A4( us02_n714 ) , .A3( us02_n715 ) , .A2( us02_n716 ) , .A1( us02_n717 ) , .ZN( us02_n718 ) );
  INV_X1 us02_U12 (.A( us02_n679 ) , .ZN( us02_n839 ) );
  NAND4_X1 us02_U120 (.A4( us02_n472 ) , .A3( us02_n473 ) , .A2( us02_n474 ) , .A1( us02_n475 ) , .ZN( us02_n677 ) );
  NOR4_X1 us02_U121 (.A4( us02_n469 ) , .ZN( us02_n475 ) , .A3( us02_n555 ) , .A1( us02_n734 ) , .A2( us02_n754 ) );
  NOR4_X1 us02_U122 (.ZN( us02_n474 ) , .A1( us02_n530 ) , .A3( us02_n567 ) , .A4( us02_n599 ) , .A2( us02_n641 ) );
  NOR4_X1 us02_U123 (.ZN( us02_n473 ) , .A1( us02_n505 ) , .A3( us02_n543 ) , .A2( us02_n582 ) , .A4( us02_n715 ) );
  NOR2_X1 us02_U124 (.ZN( us02_n732 ) , .A2( us02_n831 ) , .A1( us02_n844 ) );
  NOR2_X1 us02_U125 (.ZN( us02_n788 ) , .A2( us02_n861 ) , .A1( us02_n867 ) );
  NOR2_X1 us02_U126 (.ZN( us02_n646 ) , .A1( us02_n853 ) , .A2( us02_n867 ) );
  NAND4_X1 us02_U127 (.A4( us02_n572 ) , .A3( us02_n573 ) , .A1( us02_n574 ) , .ZN( us02_n722 ) , .A2( us02_n873 ) );
  NOR4_X1 us02_U128 (.A4( us02_n568 ) , .A3( us02_n569 ) , .A2( us02_n570 ) , .A1( us02_n571 ) , .ZN( us02_n572 ) );
  AOI221_X1 us02_U129 (.A( us02_n563 ) , .C2( us02_n564 ) , .ZN( us02_n573 ) , .B2( us02_n844 ) , .B1( us02_n851 ) , .C1( us02_n852 ) );
  NOR4_X1 us02_U13 (.A4( us02_n444 ) , .A3( us02_n445 ) , .A2( us02_n515 ) , .A1( us02_n540 ) , .ZN( us02_n705 ) );
  INV_X1 us02_U130 (.A( us02_n606 ) , .ZN( us02_n873 ) );
  NAND4_X1 us02_U131 (.A4( us02_n492 ) , .A3( us02_n493 ) , .A1( us02_n494 ) , .ZN( us02_n801 ) , .A2( us02_n866 ) );
  AOI221_X1 us02_U132 (.A( us02_n488 ) , .ZN( us02_n493 ) , .B2( us02_n835 ) , .C2( us02_n840 ) , .C1( us02_n850 ) , .B1( us02_n859 ) );
  INV_X1 us02_U133 (.A( us02_n777 ) , .ZN( us02_n866 ) );
  NOR2_X1 us02_U134 (.ZN( us02_n494 ) , .A1( us02_n677 ) , .A2( us02_n693 ) );
  AOI222_X1 us02_U135 (.ZN( us02_n512 ) , .C1( us02_n831 ) , .B2( us02_n836 ) , .A2( us02_n842 ) , .C2( us02_n861 ) , .B1( us02_n862 ) , .A1( us02_n865 ) );
  NOR4_X1 us02_U136 (.A4( us02_n508 ) , .A2( us02_n509 ) , .A1( us02_n510 ) , .ZN( us02_n511 ) , .A3( us02_n669 ) );
  INV_X1 us02_U137 (.A( us02_n504 ) , .ZN( us02_n870 ) );
  INV_X1 us02_U138 (.A( us02_n761 ) , .ZN( us02_n829 ) );
  INV_X1 us02_U139 (.A( us02_n462 ) , .ZN( us02_n863 ) );
  OR3_X1 us02_U14 (.ZN( us02_n445 ) , .A1( us02_n527 ) , .A3( us02_n576 ) , .A2( us02_n874 ) );
  OAI21_X1 us02_U140 (.ZN( us02_n462 ) , .B1( us02_n808 ) , .A( us02_n833 ) , .B2( us02_n850 ) );
  OR4_X1 us02_U141 (.A4( us02_n565 ) , .A3( us02_n566 ) , .A2( us02_n567 ) , .ZN( us02_n571 ) , .A1( us02_n664 ) );
  OR4_X1 us02_U142 (.A4( us02_n517 ) , .A2( us02_n518 ) , .A1( us02_n519 ) , .ZN( us02_n521 ) , .A3( us02_n820 ) );
  OR4_X1 us02_U143 (.ZN( us02_n465 ) , .A4( us02_n517 ) , .A3( us02_n528 ) , .A2( us02_n577 ) , .A1( us02_n711 ) );
  OR4_X1 us02_U144 (.A4( us02_n681 ) , .A3( us02_n682 ) , .A2( us02_n683 ) , .A1( us02_n684 ) , .ZN( us02_n689 ) );
  OR4_X1 us02_U145 (.A4( us02_n579 ) , .A3( us02_n580 ) , .A2( us02_n581 ) , .A1( us02_n582 ) , .ZN( us02_n583 ) );
  NAND2_X1 us02_U146 (.ZN( us02_n612 ) , .A2( us02_n836 ) , .A1( us02_n872 ) );
  OR3_X1 us02_U147 (.A3( us02_n505 ) , .A2( us02_n506 ) , .A1( us02_n507 ) , .ZN( us02_n510 ) );
  AOI221_X1 us02_U148 (.A( us02_n712 ) , .B2( us02_n713 ) , .ZN( us02_n719 ) , .C1( us02_n831 ) , .B1( us02_n838 ) , .C2( us02_n862 ) );
  OR2_X1 us02_U149 (.A2( us02_n710 ) , .A1( us02_n711 ) , .ZN( us02_n712 ) );
  OR4_X1 us02_U15 (.A4( us02_n441 ) , .A2( us02_n442 ) , .A1( us02_n443 ) , .ZN( us02_n444 ) , .A3( us02_n552 ) );
  INV_X1 us02_U150 (.A( us02_n753 ) , .ZN( us02_n868 ) );
  OAI21_X1 us02_U151 (.B1( us02_n752 ) , .ZN( us02_n753 ) , .A( us02_n844 ) , .B2( us02_n867 ) );
  INV_X1 us02_U152 (.A( us02_n671 ) , .ZN( us02_n858 ) );
  AOI21_X1 us02_U153 (.A( us02_n669 ) , .B1( us02_n670 ) , .ZN( us02_n671 ) , .B2( us02_n855 ) );
  NAND2_X1 us02_U154 (.A1( us02_n446 ) , .A2( us02_n464 ) , .ZN( us02_n748 ) );
  OAI222_X1 us02_U155 (.B2( us02_n746 ) , .B1( us02_n747 ) , .A2( us02_n748 ) , .ZN( us02_n756 ) , .C2( us02_n804 ) , .C1( us02_n813 ) , .A1( us02_n816 ) );
  OAI222_X1 us02_U156 (.ZN( us02_n504 ) , .C2( us02_n624 ) , .B2( us02_n646 ) , .B1( us02_n746 ) , .A2( us02_n747 ) , .C1( us02_n804 ) , .A1( us02_n805 ) );
  OAI222_X1 us02_U157 (.B2( us02_n707 ) , .ZN( us02_n708 ) , .C2( us02_n723 ) , .B1( us02_n746 ) , .A1( us02_n805 ) , .C1( us02_n813 ) , .A2( us02_n814 ) );
  OAI222_X1 us02_U158 (.ZN( us02_n616 ) , .B1( us02_n696 ) , .C1( us02_n723 ) , .C2( us02_n746 ) , .B2( us02_n785 ) , .A2( us02_n791 ) , .A1( us02_n815 ) );
  NOR4_X1 us02_U159 (.A2( us02_n490 ) , .A1( us02_n491 ) , .ZN( us02_n492 ) , .A3( us02_n579 ) , .A4( us02_n611 ) );
  INV_X1 us02_U16 (.A( us02_n612 ) , .ZN( us02_n874 ) );
  OR4_X1 us02_U160 (.ZN( us02_n491 ) , .A4( us02_n533 ) , .A2( us02_n546 ) , .A1( us02_n558 ) , .A3( us02_n631 ) );
  OAI22_X1 us02_U161 (.B1( us02_n489 ) , .ZN( us02_n490 ) , .A1( us02_n685 ) , .A2( us02_n762 ) , .B2( us02_n816 ) );
  NOR3_X1 us02_U162 (.ZN( us02_n489 ) , .A1( us02_n781 ) , .A2( us02_n849 ) , .A3( us02_n862 ) );
  AOI22_X1 us02_U163 (.ZN( us02_n695 ) , .A1( us02_n829 ) , .B2( us02_n842 ) , .A2( us02_n864 ) , .B1( us02_n867 ) );
  INV_X1 us02_U164 (.A( us02_n729 ) , .ZN( us02_n838 ) );
  AOI221_X1 us02_U165 (.A( us02_n763 ) , .ZN( us02_n773 ) , .C2( us02_n809 ) , .B2( us02_n834 ) , .C1( us02_n854 ) , .B1( us02_n865 ) );
  AOI21_X1 us02_U166 (.B2( us02_n762 ) , .ZN( us02_n763 ) , .A( us02_n787 ) , .B1( us02_n791 ) );
  INV_X1 us02_U167 (.A( us02_n760 ) , .ZN( us02_n834 ) );
  AOI221_X1 us02_U168 (.A( us02_n482 ) , .ZN( us02_n487 ) , .B1( us02_n830 ) , .C2( us02_n843 ) , .C1( us02_n851 ) , .B2( us02_n861 ) );
  OAI22_X1 us02_U169 (.ZN( us02_n482 ) , .A1( us02_n707 ) , .B2( us02_n784 ) , .A2( us02_n805 ) , .B1( us02_n811 ) );
  INV_X1 us02_U17 (.A( us02_n748 ) , .ZN( us02_n862 ) );
  INV_X1 us02_U170 (.A( us02_n789 ) , .ZN( us02_n831 ) );
  NAND2_X1 us02_U171 (.A1( us02_n450 ) , .A2( us02_n452 ) , .ZN( us02_n761 ) );
  OAI221_X1 us02_U172 (.A( us02_n726 ) , .C2( us02_n727 ) , .B2( us02_n728 ) , .B1( us02_n729 ) , .ZN( us02_n736 ) , .C1( us02_n816 ) );
  AOI22_X1 us02_U173 (.ZN( us02_n726 ) , .B1( us02_n831 ) , .A2( us02_n837 ) , .A1( us02_n862 ) , .B2( us02_n865 ) );
  INV_X1 us02_U174 (.A( us02_n785 ) , .ZN( us02_n861 ) );
  OAI22_X1 us02_U175 (.ZN( us02_n709 ) , .A2( us02_n727 ) , .B2( us02_n728 ) , .A1( us02_n743 ) , .B1( us02_n812 ) );
  INV_X1 us02_U176 (.A( us02_n815 ) , .ZN( us02_n830 ) );
  OAI22_X1 us02_U177 (.ZN( us02_n488 ) , .A1( us02_n723 ) , .B2( us02_n727 ) , .B1( us02_n729 ) , .A2( us02_n778 ) );
  OAI22_X1 us02_U178 (.ZN( us02_n623 ) , .B1( us02_n668 ) , .B2( us02_n746 ) , .A1( us02_n814 ) , .A2( us02_n815 ) );
  INV_X1 us02_U179 (.A( us02_n743 ) , .ZN( us02_n836 ) );
  AOI222_X1 us02_U18 (.ZN( us02_n604 ) , .B2( us02_n670 ) , .B1( us02_n752 ) , .C2( us02_n830 ) , .A1( us02_n832 ) , .A2( us02_n861 ) , .C1( us02_n862 ) );
  OAI22_X1 us02_U180 (.A1( us02_n723 ) , .ZN( us02_n725 ) , .B2( us02_n749 ) , .B1( us02_n811 ) , .A2( us02_n815 ) );
  OAI22_X1 us02_U181 (.B2( us02_n778 ) , .B1( us02_n779 ) , .ZN( us02_n780 ) , .A2( us02_n813 ) , .A1( us02_n814 ) );
  INV_X1 us02_U182 (.A( us02_n787 ) , .ZN( us02_n844 ) );
  INV_X1 us02_U183 (.A( us02_n804 ) , .ZN( us02_n859 ) );
  INV_X1 us02_U184 (.A( us02_n813 ) , .ZN( us02_n832 ) );
  OAI22_X1 us02_U185 (.B2( us02_n743 ) , .ZN( us02_n745 ) , .A2( us02_n761 ) , .B1( us02_n779 ) , .A1( us02_n791 ) );
  OAI22_X1 us02_U186 (.B2( us02_n802 ) , .B1( us02_n803 ) , .A2( us02_n804 ) , .A1( us02_n805 ) , .ZN( us02_n807 ) );
  OAI22_X1 us02_U187 (.ZN( us02_n495 ) , .A2( us02_n743 ) , .A1( us02_n779 ) , .B1( us02_n790 ) , .B2( us02_n805 ) );
  OAI22_X1 us02_U188 (.ZN( us02_n589 ) , .B1( us02_n729 ) , .B2( us02_n748 ) , .A2( us02_n785 ) , .A1( us02_n802 ) );
  OAI22_X1 us02_U189 (.ZN( us02_n694 ) , .A2( us02_n729 ) , .A1( us02_n779 ) , .B1( us02_n790 ) , .B2( us02_n816 ) );
  AOI222_X1 us02_U19 (.ZN( us02_n562 ) , .B1( us02_n829 ) , .C1( us02_n840 ) , .A2( us02_n842 ) , .A1( us02_n853 ) , .B2( us02_n862 ) , .C2( us02_n872 ) );
  INV_X1 us02_U190 (.A( us02_n802 ) , .ZN( us02_n842 ) );
  INV_X1 us02_U191 (.A( us02_n668 ) , .ZN( us02_n864 ) );
  OAI22_X1 us02_U192 (.ZN( us02_n636 ) , .A1( us02_n698 ) , .B2( us02_n727 ) , .A2( us02_n761 ) , .B1( us02_n815 ) );
  NOR2_X1 us02_U193 (.ZN( us02_n714 ) , .A1( us02_n804 ) , .A2( us02_n816 ) );
  NOR2_X1 us02_U194 (.A1( us02_n696 ) , .ZN( us02_n769 ) , .A2( us02_n814 ) );
  NOR2_X1 us02_U195 (.ZN( us02_n665 ) , .A1( us02_n727 ) , .A2( us02_n802 ) );
  NOR2_X1 us02_U196 (.ZN( us02_n593 ) , .A2( us02_n696 ) , .A1( us02_n727 ) );
  NOR2_X1 us02_U197 (.ZN( us02_n569 ) , .A1( us02_n727 ) , .A2( us02_n805 ) );
  NOR2_X1 us02_U198 (.A2( us02_n743 ) , .ZN( us02_n754 ) , .A1( us02_n804 ) );
  NOR2_X1 us02_U199 (.ZN( us02_n717 ) , .A2( us02_n723 ) , .A1( us02_n743 ) );
  AOI222_X1 us02_U20 (.ZN( us02_n659 ) , .A2( us02_n838 ) , .B1( us02_n840 ) , .C2( us02_n844 ) , .A1( us02_n859 ) , .C1( us02_n862 ) , .B2( us02_n869 ) );
  NOR2_X1 us02_U200 (.ZN( us02_n734 ) , .A2( us02_n802 ) , .A1( us02_n804 ) );
  NOR2_X1 us02_U201 (.ZN( us02_n545 ) , .A2( us02_n779 ) , .A1( us02_n813 ) );
  NOR2_X1 us02_U202 (.ZN( us02_n576 ) , .A2( us02_n698 ) , .A1( us02_n813 ) );
  NOR2_X1 us02_U203 (.ZN( us02_n653 ) , .A1( us02_n727 ) , .A2( us02_n812 ) );
  NOR2_X1 us02_U204 (.ZN( us02_n611 ) , .A1( us02_n778 ) , .A2( us02_n785 ) );
  INV_X1 us02_U205 (.A( us02_n749 ) , .ZN( us02_n841 ) );
  NOR2_X1 us02_U206 (.ZN( us02_n531 ) , .A2( us02_n748 ) , .A1( us02_n749 ) );
  NOR2_X1 us02_U207 (.ZN( us02_n628 ) , .A2( us02_n727 ) , .A1( us02_n784 ) );
  NOR2_X1 us02_U208 (.ZN( us02_n614 ) , .A1( us02_n784 ) , .A2( us02_n814 ) );
  NOR2_X1 us02_U209 (.ZN( us02_n600 ) , .A2( us02_n779 ) , .A1( us02_n802 ) );
  INV_X1 us02_U21 (.A( us02_n646 ) , .ZN( us02_n869 ) );
  NOR2_X1 us02_U210 (.ZN( us02_n610 ) , .A2( us02_n779 ) , .A1( us02_n805 ) );
  INV_X1 us02_U211 (.A( us02_n746 ) , .ZN( us02_n833 ) );
  NOR2_X1 us02_U212 (.A2( us02_n743 ) , .ZN( us02_n768 ) , .A1( us02_n811 ) );
  NOR2_X1 us02_U213 (.ZN( us02_n527 ) , .A2( us02_n723 ) , .A1( us02_n802 ) );
  NOR2_X1 us02_U214 (.ZN( us02_n530 ) , .A2( us02_n779 ) , .A1( us02_n815 ) );
  NOR2_X1 us02_U215 (.ZN( us02_n627 ) , .A2( us02_n668 ) , .A1( us02_n784 ) );
  NOR2_X1 us02_U216 (.ZN( us02_n598 ) , .A2( us02_n790 ) , .A1( us02_n815 ) );
  INV_X1 us02_U217 (.A( us02_n727 ) , .ZN( us02_n851 ) );
  NOR2_X1 us02_U218 (.ZN( us02_n651 ) , .A1( us02_n668 ) , .A2( us02_n813 ) );
  NOR2_X1 us02_U219 (.A1( us02_n668 ) , .ZN( us02_n672 ) , .A2( us02_n743 ) );
  NOR4_X1 us02_U22 (.ZN( us02_n472 ) , .A2( us02_n520 ) , .A4( us02_n593 ) , .A1( us02_n608 ) , .A3( us02_n628 ) );
  NOR2_X1 us02_U220 (.ZN( us02_n601 ) , .A1( us02_n668 ) , .A2( us02_n802 ) );
  NOR2_X1 us02_U221 (.A1( us02_n668 ) , .ZN( us02_n687 ) , .A2( us02_n815 ) );
  INV_X1 us02_U222 (.A( us02_n791 ) , .ZN( us02_n850 ) );
  NOR2_X1 us02_U223 (.A2( us02_n707 ) , .A1( us02_n749 ) , .ZN( us02_n770 ) );
  NOR2_X1 us02_U224 (.A1( us02_n668 ) , .ZN( us02_n765 ) , .A2( us02_n812 ) );
  NOR2_X1 us02_U225 (.A1( us02_n698 ) , .ZN( us02_n767 ) , .A2( us02_n812 ) );
  NOR2_X1 us02_U226 (.ZN( us02_n540 ) , .A2( us02_n696 ) , .A1( us02_n698 ) );
  NOR2_X1 us02_U227 (.ZN( us02_n526 ) , .A1( us02_n668 ) , .A2( us02_n778 ) );
  NOR2_X1 us02_U228 (.ZN( us02_n666 ) , .A1( us02_n749 ) , .A2( us02_n814 ) );
  NOR2_X1 us02_U229 (.ZN( us02_n554 ) , .A1( us02_n749 ) , .A2( us02_n790 ) );
  NOR4_X1 us02_U23 (.ZN( us02_n478 ) , .A1( us02_n519 ) , .A4( us02_n556 ) , .A3( us02_n581 ) , .A2( us02_n629 ) );
  NOR2_X1 us02_U230 (.ZN( us02_n507 ) , .A2( us02_n779 ) , .A1( us02_n784 ) );
  NOR2_X1 us02_U231 (.ZN( us02_n542 ) , .A2( us02_n707 ) , .A1( us02_n784 ) );
  NOR2_X1 us02_U232 (.ZN( us02_n663 ) , .A1( us02_n784 ) , .A2( us02_n790 ) );
  NOR2_X1 us02_U233 (.A2( us02_n696 ) , .ZN( us02_n715 ) , .A1( us02_n791 ) );
  NOR2_X1 us02_U234 (.ZN( us02_n506 ) , .A1( us02_n811 ) , .A2( us02_n816 ) );
  NOR2_X1 us02_U235 (.ZN( us02_n555 ) , .A1( us02_n761 ) , .A2( us02_n804 ) );
  NOR2_X1 us02_U236 (.ZN( us02_n660 ) , .A1( us02_n728 ) , .A2( us02_n789 ) );
  NOR2_X1 us02_U237 (.ZN( us02_n661 ) , .A2( us02_n696 ) , .A1( us02_n728 ) );
  NOR2_X1 us02_U238 (.ZN( us02_n556 ) , .A1( us02_n791 ) , .A2( us02_n813 ) );
  NOR2_X1 us02_U239 (.ZN( us02_n544 ) , .A1( us02_n748 ) , .A2( us02_n813 ) );
  NOR4_X1 us02_U24 (.A4( us02_n531 ) , .A3( us02_n532 ) , .A2( us02_n533 ) , .ZN( us02_n534 ) , .A1( us02_n819 ) );
  NOR2_X1 us02_U240 (.ZN( us02_n508 ) , .A1( us02_n728 ) , .A2( us02_n778 ) );
  NOR2_X1 us02_U241 (.A2( us02_n696 ) , .A1( us02_n779 ) , .ZN( us02_n819 ) );
  OAI22_X1 us02_U242 (.B2( us02_n749 ) , .B1( us02_n750 ) , .A1( us02_n751 ) , .ZN( us02_n755 ) , .A2( us02_n805 ) );
  NOR2_X1 us02_U243 (.ZN( us02_n750 ) , .A2( us02_n851 ) , .A1( us02_n859 ) );
  NOR3_X1 us02_U244 (.ZN( us02_n751 ) , .A2( us02_n852 ) , .A1( us02_n862 ) , .A3( us02_n864 ) );
  NOR2_X1 us02_U245 (.ZN( us02_n529 ) , .A2( us02_n743 ) , .A1( us02_n791 ) );
  NOR2_X1 us02_U246 (.A1( us02_n748 ) , .ZN( us02_n766 ) , .A2( us02_n802 ) );
  NOR2_X1 us02_U247 (.ZN( us02_n543 ) , .A2( us02_n784 ) , .A1( us02_n791 ) );
  NOR2_X1 us02_U248 (.ZN( us02_n662 ) , .A1( us02_n728 ) , .A2( us02_n784 ) );
  NOR2_X1 us02_U249 (.ZN( us02_n630 ) , .A1( us02_n723 ) , .A2( us02_n812 ) );
  NOR4_X1 us02_U25 (.ZN( us02_n455 ) , .A2( us02_n516 ) , .A1( us02_n542 ) , .A3( us02_n578 ) , .A4( us02_n614 ) );
  NOR2_X1 us02_U250 (.ZN( us02_n613 ) , .A1( us02_n761 ) , .A2( us02_n811 ) );
  OAI22_X1 us02_U251 (.B1( us02_n439 ) , .ZN( us02_n443 ) , .A2( us02_n727 ) , .A1( us02_n743 ) , .B2( us02_n748 ) );
  NOR3_X1 us02_U252 (.ZN( us02_n439 ) , .A2( us02_n835 ) , .A3( us02_n836 ) , .A1( us02_n845 ) );
  NOR2_X1 us02_U253 (.ZN( us02_n505 ) , .A2( us02_n727 ) , .A1( us02_n761 ) );
  NOR2_X1 us02_U254 (.ZN( us02_n515 ) , .A1( us02_n707 ) , .A2( us02_n743 ) );
  NOR2_X1 us02_U255 (.ZN( us02_n716 ) , .A2( us02_n743 ) , .A1( us02_n785 ) );
  NOR2_X1 us02_U256 (.ZN( us02_n553 ) , .A1( us02_n785 ) , .A2( us02_n812 ) );
  NOR2_X1 us02_U257 (.ZN( us02_n516 ) , .A1( us02_n707 ) , .A2( us02_n802 ) );
  NOR2_X1 us02_U258 (.ZN( us02_n557 ) , .A1( us02_n707 ) , .A2( us02_n815 ) );
  NOR2_X1 us02_U259 (.ZN( us02_n669 ) , .A1( us02_n789 ) , .A2( us02_n804 ) );
  NOR4_X1 us02_U26 (.A4( us02_n540 ) , .A3( us02_n541 ) , .A2( us02_n542 ) , .ZN( us02_n549 ) , .A1( us02_n687 ) );
  NOR2_X1 us02_U260 (.ZN( us02_n520 ) , .A1( us02_n789 ) , .A2( us02_n811 ) );
  NOR2_X1 us02_U261 (.ZN( us02_n629 ) , .A1( us02_n746 ) , .A2( us02_n814 ) );
  INV_X1 us02_U262 (.A( us02_n805 ) , .ZN( us02_n840 ) );
  AOI21_X1 us02_U263 (.ZN( us02_n570 ) , .B2( us02_n696 ) , .B1( us02_n805 ) , .A( us02_n811 ) );
  NOR2_X1 us02_U264 (.ZN( us02_n654 ) , .A1( us02_n789 ) , .A2( us02_n814 ) );
  INV_X1 us02_U265 (.A( us02_n762 ) , .ZN( us02_n865 ) );
  AOI21_X1 us02_U266 (.ZN( us02_n551 ) , .B1( us02_n668 ) , .A( us02_n696 ) , .B2( us02_n804 ) );
  NOR2_X1 us02_U267 (.ZN( us02_n667 ) , .A2( us02_n707 ) , .A1( us02_n789 ) );
  NOR2_X1 us02_U268 (.ZN( us02_n655 ) , .A1( us02_n746 ) , .A2( us02_n779 ) );
  NOR2_X1 us02_U269 (.ZN( us02_n541 ) , .A1( us02_n761 ) , .A2( us02_n790 ) );
  NOR2_X1 us02_U27 (.ZN( us02_n679 ) , .A2( us02_n833 ) , .A1( us02_n838 ) );
  NOR2_X1 us02_U270 (.ZN( us02_n700 ) , .A2( us02_n785 ) , .A1( us02_n816 ) );
  NOR2_X1 us02_U271 (.ZN( us02_n608 ) , .A2( us02_n723 ) , .A1( us02_n816 ) );
  NOR2_X1 us02_U272 (.A1( us02_n729 ) , .ZN( us02_n764 ) , .A2( us02_n785 ) );
  AOI21_X1 us02_U273 (.A( us02_n814 ) , .B2( us02_n815 ) , .B1( us02_n816 ) , .ZN( us02_n817 ) );
  INV_X1 us02_U274 (.A( us02_n728 ) , .ZN( us02_n867 ) );
  NOR2_X1 us02_U275 (.ZN( us02_n578 ) , .A2( us02_n707 ) , .A1( us02_n729 ) );
  NOR2_X1 us02_U276 (.ZN( us02_n532 ) , .A2( us02_n723 ) , .A1( us02_n729 ) );
  AOI21_X1 us02_U277 (.B1( us02_n624 ) , .ZN( us02_n626 ) , .A( us02_n762 ) , .B2( us02_n813 ) );
  AOI21_X1 us02_U278 (.A( us02_n811 ) , .B2( us02_n812 ) , .B1( us02_n813 ) , .ZN( us02_n818 ) );
  AOI21_X1 us02_U279 (.ZN( us02_n514 ) , .A( us02_n728 ) , .B1( us02_n749 ) , .B2( us02_n802 ) );
  AOI222_X1 us02_U28 (.ZN( us02_n468 ) , .B1( us02_n831 ) , .A1( us02_n838 ) , .C1( us02_n841 ) , .C2( us02_n850 ) , .A2( us02_n854 ) , .B2( us02_n864 ) );
  AOI21_X1 us02_U280 (.ZN( us02_n498 ) , .B1( us02_n679 ) , .A( us02_n811 ) , .B2( us02_n815 ) );
  AOI21_X1 us02_U281 (.ZN( us02_n649 ) , .A( us02_n778 ) , .B1( us02_n791 ) , .B2( us02_n804 ) );
  AOI21_X1 us02_U282 (.ZN( us02_n477 ) , .B2( us02_n696 ) , .A( us02_n748 ) , .B1( us02_n778 ) );
  NOR2_X1 us02_U283 (.ZN( us02_n581 ) , .A1( us02_n743 ) , .A2( us02_n814 ) );
  AOI21_X1 us02_U284 (.ZN( us02_n592 ) , .B1( us02_n749 ) , .A( us02_n791 ) , .B2( us02_n812 ) );
  NOR2_X1 us02_U285 (.A2( us02_n707 ) , .A1( us02_n761 ) , .ZN( us02_n793 ) );
  AOI21_X1 us02_U286 (.ZN( us02_n625 ) , .B2( us02_n668 ) , .A( us02_n789 ) , .B1( us02_n790 ) );
  NOR2_X1 us02_U287 (.ZN( us02_n519 ) , .A2( us02_n707 ) , .A1( us02_n813 ) );
  AOI21_X1 us02_U288 (.ZN( us02_n476 ) , .A( us02_n668 ) , .B1( us02_n749 ) , .B2( us02_n805 ) );
  NOR2_X1 us02_U289 (.ZN( us02_n558 ) , .A2( us02_n790 ) , .A1( us02_n802 ) );
  NOR4_X1 us02_U29 (.A1( us02_n465 ) , .ZN( us02_n466 ) , .A4( us02_n541 ) , .A2( us02_n553 ) , .A3( us02_n613 ) );
  NOR2_X1 us02_U290 (.ZN( us02_n518 ) , .A2( us02_n698 ) , .A1( us02_n815 ) );
  NOR2_X1 us02_U291 (.ZN( us02_n682 ) , .A2( us02_n698 ) , .A1( us02_n802 ) );
  NOR2_X1 us02_U292 (.ZN( us02_n652 ) , .A1( us02_n761 ) , .A2( us02_n785 ) );
  INV_X1 us02_U293 (.A( us02_n812 ) , .ZN( us02_n835 ) );
  AOI21_X1 us02_U294 (.ZN( us02_n509 ) , .B2( us02_n668 ) , .A( us02_n729 ) , .B1( us02_n814 ) );
  AOI21_X1 us02_U295 (.ZN( us02_n538 ) , .B2( us02_n811 ) , .A( us02_n813 ) , .B1( us02_n814 ) );
  AOI21_X1 us02_U296 (.ZN( us02_n539 ) , .A( us02_n762 ) , .B2( us02_n778 ) , .B1( us02_n816 ) );
  NOR2_X1 us02_U297 (.ZN( us02_n580 ) , .A1( us02_n668 ) , .A2( us02_n787 ) );
  AOI21_X1 us02_U298 (.ZN( us02_n588 ) , .B2( us02_n698 ) , .B1( us02_n814 ) , .A( us02_n816 ) );
  AOI21_X1 us02_U299 (.B1( us02_n698 ) , .ZN( us02_n699 ) , .A( us02_n731 ) , .B2( us02_n762 ) );
  NAND2_X1 us02_U3 (.A1( us02_n440 ) , .A2( us02_n463 ) , .ZN( us02_n707 ) );
  AOI221_X1 us02_U30 (.ZN( us02_n467 ) , .C2( us02_n713 ) , .B2( us02_n830 ) , .C1( us02_n844 ) , .B1( us02_n859 ) , .A( us02_n863 ) );
  AOI21_X1 us02_U300 (.ZN( us02_n590 ) , .B2( us02_n762 ) , .A( us02_n784 ) , .B1( us02_n811 ) );
  AOI21_X1 us02_U301 (.ZN( us02_n497 ) , .A( us02_n723 ) , .B2( us02_n761 ) , .B1( us02_n813 ) );
  NOR2_X1 us02_U302 (.ZN( us02_n546 ) , .A1( us02_n698 ) , .A2( us02_n743 ) );
  INV_X1 us02_U303 (.A( us02_n790 ) , .ZN( us02_n872 ) );
  INV_X1 us02_U304 (.A( us02_n811 ) , .ZN( us02_n853 ) );
  AOI21_X1 us02_U305 (.ZN( us02_n648 ) , .B1( us02_n728 ) , .B2( us02_n762 ) , .A( us02_n812 ) );
  NOR2_X1 us02_U306 (.ZN( us02_n684 ) , .A1( us02_n728 ) , .A2( us02_n815 ) );
  AOI21_X1 us02_U307 (.B1( us02_n685 ) , .ZN( us02_n686 ) , .A( us02_n727 ) , .B2( us02_n760 ) );
  AOI21_X1 us02_U308 (.ZN( us02_n568 ) , .B1( us02_n749 ) , .B2( us02_n761 ) , .A( us02_n779 ) );
  AOI21_X1 us02_U309 (.ZN( us02_n499 ) , .A( us02_n696 ) , .B1( us02_n707 ) , .B2( us02_n785 ) );
  NOR4_X1 us02_U31 (.A4( us02_n513 ) , .A3( us02_n514 ) , .A2( us02_n515 ) , .A1( us02_n516 ) , .ZN( us02_n523 ) );
  NOR2_X1 us02_U310 (.ZN( us02_n567 ) , .A1( us02_n728 ) , .A2( us02_n761 ) );
  NOR2_X1 us02_U311 (.ZN( us02_n579 ) , .A2( us02_n696 ) , .A1( us02_n790 ) );
  NOR2_X1 us02_U312 (.ZN( us02_n565 ) , .A2( us02_n696 ) , .A1( us02_n762 ) );
  AOI21_X1 us02_U313 (.ZN( us02_n513 ) , .A( us02_n778 ) , .B2( us02_n791 ) , .B1( us02_n811 ) );
  INV_X1 us02_U314 (.A( us02_n698 ) , .ZN( us02_n852 ) );
  NOR2_X1 us02_U315 (.ZN( us02_n664 ) , .A1( us02_n779 ) , .A2( us02_n812 ) );
  AOI21_X1 us02_U316 (.ZN( us02_n449 ) , .B2( us02_n791 ) , .A( us02_n802 ) , .B1( us02_n814 ) );
  NOR2_X1 us02_U317 (.ZN( us02_n631 ) , .A2( us02_n696 ) , .A1( us02_n723 ) );
  AOI21_X1 us02_U318 (.ZN( us02_n563 ) , .B1( us02_n723 ) , .A( us02_n778 ) , .B2( us02_n790 ) );
  AOI21_X1 us02_U319 (.ZN( us02_n496 ) , .A( us02_n778 ) , .B2( us02_n790 ) , .B1( us02_n803 ) );
  AOI222_X1 us02_U32 (.ZN( us02_n524 ) , .A1( us02_n833 ) , .B2( us02_n836 ) , .C1( us02_n843 ) , .C2( us02_n849 ) , .A2( us02_n851 ) , .B1( us02_n865 ) );
  NAND2_X1 us02_U320 (.ZN( us02_n752 ) , .A1( us02_n762 ) , .A2( us02_n804 ) );
  NOR2_X1 us02_U321 (.ZN( us02_n528 ) , .A1( us02_n707 ) , .A2( us02_n778 ) );
  NOR2_X1 us02_U322 (.ZN( us02_n577 ) , .A1( us02_n707 ) , .A2( us02_n812 ) );
  AOI21_X1 us02_U323 (.ZN( us02_n688 ) , .B2( us02_n748 ) , .B1( us02_n762 ) , .A( us02_n805 ) );
  NOR2_X1 us02_U324 (.ZN( us02_n566 ) , .A1( us02_n746 ) , .A2( us02_n804 ) );
  NOR2_X1 us02_U325 (.ZN( us02_n683 ) , .A1( us02_n790 ) , .A2( us02_n812 ) );
  NOR2_X1 us02_U326 (.A2( us02_n812 ) , .A1( us02_n814 ) , .ZN( us02_n820 ) );
  AOI21_X1 us02_U327 (.A( us02_n789 ) , .B2( us02_n790 ) , .B1( us02_n791 ) , .ZN( us02_n792 ) );
  AOI21_X1 us02_U328 (.A( us02_n732 ) , .ZN( us02_n733 ) , .B2( us02_n779 ) , .B1( us02_n791 ) );
  NOR2_X1 us02_U329 (.ZN( us02_n710 ) , .A1( us02_n761 ) , .A2( us02_n762 ) );
  NOR4_X1 us02_U33 (.A3( us02_n520 ) , .A1( us02_n521 ) , .ZN( us02_n522 ) , .A2( us02_n672 ) , .A4( us02_n768 ) );
  NOR2_X1 us02_U330 (.ZN( us02_n582 ) , .A1( us02_n791 ) , .A2( us02_n816 ) );
  NOR2_X1 us02_U331 (.ZN( us02_n533 ) , .A1( us02_n723 ) , .A2( us02_n787 ) );
  NOR2_X1 us02_U332 (.ZN( us02_n681 ) , .A2( us02_n707 ) , .A1( us02_n816 ) );
  INV_X1 us02_U333 (.A( us02_n696 ) , .ZN( us02_n837 ) );
  NOR2_X1 us02_U334 (.ZN( us02_n641 ) , .A2( us02_n787 ) , .A1( us02_n790 ) );
  INV_X1 us02_U335 (.A( us02_n814 ) , .ZN( us02_n854 ) );
  AOI21_X1 us02_U336 (.ZN( us02_n441 ) , .A( us02_n698 ) , .B1( us02_n732 ) , .B2( us02_n749 ) );
  INV_X1 us02_U337 (.A( us02_n779 ) , .ZN( us02_n849 ) );
  AOI22_X1 us02_U338 (.A2( us02_n781 ) , .ZN( us02_n782 ) , .B2( us02_n830 ) , .A1( us02_n833 ) , .B1( us02_n862 ) );
  NAND2_X1 us02_U339 (.ZN( us02_n670 ) , .A1( us02_n805 ) , .A2( us02_n815 ) );
  NOR4_X1 us02_U34 (.A3( us02_n754 ) , .A2( us02_n755 ) , .A1( us02_n756 ) , .ZN( us02_n757 ) , .A4( us02_n868 ) );
  NAND2_X1 us02_U340 (.ZN( us02_n713 ) , .A1( us02_n727 ) , .A2( us02_n779 ) );
  NAND2_X1 us02_U341 (.A2( us02_n761 ) , .A1( us02_n805 ) , .ZN( us02_n809 ) );
  AOI21_X1 us02_U342 (.ZN( us02_n442 ) , .B1( us02_n788 ) , .B2( us02_n790 ) , .A( us02_n813 ) );
  NOR2_X1 us02_U343 (.ZN( us02_n483 ) , .A1( us02_n787 ) , .A2( us02_n804 ) );
  NOR2_X1 us02_U344 (.ZN( us02_n469 ) , .A2( us02_n778 ) , .A1( us02_n814 ) );
  INV_X1 us02_U345 (.A( us02_n784 ) , .ZN( us02_n845 ) );
  OAI21_X1 us02_U346 (.A( us02_n786 ) , .B2( us02_n787 ) , .B1( us02_n788 ) , .ZN( us02_n794 ) );
  OAI21_X1 us02_U347 (.ZN( us02_n786 ) , .A( us02_n838 ) , .B1( us02_n862 ) , .B2( us02_n872 ) );
  NOR2_X1 us02_U348 (.ZN( us02_n711 ) , .A2( us02_n723 ) , .A1( us02_n789 ) );
  NOR2_X1 us02_U349 (.ZN( us02_n525 ) , .A1( us02_n723 ) , .A2( us02_n749 ) );
  AOI211_X1 us02_U35 (.B( us02_n744 ) , .A( us02_n745 ) , .ZN( us02_n758 ) , .C1( us02_n831 ) , .C2( us02_n852 ) );
  NAND2_X1 us02_U350 (.A1( us02_n698 ) , .A2( us02_n728 ) , .ZN( us02_n781 ) );
  AOI21_X1 us02_U351 (.ZN( us02_n638 ) , .B2( us02_n748 ) , .A( us02_n787 ) , .B1( us02_n811 ) );
  AOI21_X1 us02_U352 (.ZN( us02_n639 ) , .B2( us02_n746 ) , .A( us02_n791 ) , .B1( us02_n802 ) );
  AOI21_X1 us02_U353 (.ZN( us02_n640 ) , .B1( us02_n679 ) , .A( us02_n790 ) , .B2( us02_n816 ) );
  NOR2_X1 us02_U354 (.ZN( us02_n517 ) , .A1( us02_n707 ) , .A2( us02_n787 ) );
  OAI21_X1 us02_U355 (.A( us02_n697 ) , .ZN( us02_n701 ) , .B2( us02_n749 ) , .B1( us02_n803 ) );
  OAI21_X1 us02_U356 (.ZN( us02_n697 ) , .B2( us02_n832 ) , .B1( us02_n837 ) , .A( us02_n859 ) );
  OAI21_X1 us02_U357 (.A( us02_n730 ) , .B1( us02_n731 ) , .ZN( us02_n735 ) , .B2( us02_n804 ) );
  OAI21_X1 us02_U358 (.ZN( us02_n730 ) , .A( us02_n832 ) , .B2( us02_n851 ) , .B1( us02_n872 ) );
  NAND2_X1 us02_U359 (.A2( us02_n748 ) , .A1( us02_n785 ) , .ZN( us02_n808 ) );
  NOR3_X1 us02_U36 (.A3( us02_n740 ) , .A2( us02_n741 ) , .A1( us02_n742 ) , .ZN( us02_n759 ) );
  INV_X1 us02_U360 (.A( us02_n816 ) , .ZN( us02_n843 ) );
  INV_X1 us02_U361 (.A( us02_n723 ) , .ZN( us02_n855 ) );
  AND2_X1 us02_U362 (.ZN( us02_n731 ) , .A1( us02_n778 ) , .A2( us02_n784 ) );
  NAND2_X1 us02_U363 (.A1( us02_n446 ) , .A2( us02_n448 ) , .ZN( us02_n804 ) );
  NAND2_X1 us02_U364 (.A1( us02_n454 ) , .A2( us02_n470 ) , .ZN( us02_n802 ) );
  NAND2_X1 us02_U365 (.A1( us02_n450 ) , .A2( us02_n453 ) , .ZN( us02_n813 ) );
  NAND2_X1 us02_U366 (.A1( us02_n450 ) , .A2( us02_n470 ) , .ZN( us02_n815 ) );
  NAND2_X1 us02_U367 (.A1( us02_n453 ) , .A2( us02_n460 ) , .ZN( us02_n812 ) );
  NAND2_X1 us02_U368 (.A1( us02_n452 ) , .A2( us02_n460 ) , .ZN( us02_n743 ) );
  NAND2_X1 us02_U369 (.A1( us02_n451 ) , .A2( us02_n464 ) , .ZN( us02_n668 ) );
  NOR4_X1 us02_U37 (.A4( us02_n733 ) , .A3( us02_n734 ) , .A2( us02_n735 ) , .A1( us02_n736 ) , .ZN( us02_n737 ) );
  NAND2_X1 us02_U370 (.A2( us02_n447 ) , .A1( us02_n459 ) , .ZN( us02_n727 ) );
  NAND2_X1 us02_U371 (.A1( us02_n454 ) , .A2( us02_n461 ) , .ZN( us02_n749 ) );
  NAND2_X1 us02_U372 (.A2( us02_n452 ) , .A1( us02_n454 ) , .ZN( us02_n805 ) );
  NAND2_X1 us02_U373 (.A2( us02_n453 ) , .A1( us02_n471 ) , .ZN( us02_n778 ) );
  NAND2_X1 us02_U374 (.A1( us02_n452 ) , .A2( us02_n471 ) , .ZN( us02_n784 ) );
  NAND2_X1 us02_U375 (.A2( us02_n463 ) , .A1( us02_n464 ) , .ZN( us02_n811 ) );
  NAND2_X1 us02_U376 (.A1( us02_n440 ) , .A2( us02_n459 ) , .ZN( us02_n698 ) );
  NAND2_X1 us02_U377 (.A2( us02_n448 ) , .A1( us02_n451 ) , .ZN( us02_n762 ) );
  NAND2_X1 us02_U378 (.A2( us02_n447 ) , .A1( us02_n451 ) , .ZN( us02_n728 ) );
  NAND2_X1 us02_U379 (.A2( us02_n460 ) , .A1( us02_n461 ) , .ZN( us02_n746 ) );
  AOI211_X1 us02_U38 (.B( us02_n724 ) , .A( us02_n725 ) , .ZN( us02_n738 ) , .C1( us02_n842 ) , .C2( us02_n854 ) );
  NAND2_X2 us02_U380 (.A2( us02_n460 ) , .A1( us02_n470 ) , .ZN( us02_n696 ) );
  NAND2_X1 us02_U381 (.A1( us02_n461 ) , .A2( us02_n471 ) , .ZN( us02_n787 ) );
  NOR2_X1 us02_U382 (.ZN( us02_n464 ) , .A2( us02_n846 ) , .A1( us02_n847 ) );
  NOR2_X1 us02_U383 (.ZN( us02_n452 ) , .A1( us02_n825 ) , .A2( us02_n826 ) );
  NOR2_X1 us02_U384 (.ZN( us02_n450 ) , .A1( us02_n827 ) , .A2( us02_n828 ) );
  NOR2_X1 us02_U385 (.ZN( us02_n446 ) , .A2( us02_n848 ) , .A1( us02_n857 ) );
  NAND2_X1 us02_U386 (.A2( us02_n453 ) , .A1( us02_n454 ) , .ZN( us02_n729 ) );
  NAND2_X1 us02_U387 (.A1( us02_n450 ) , .A2( us02_n461 ) , .ZN( us02_n789 ) );
  NAND2_X2 us02_U388 (.A2( us02_n447 ) , .A1( us02_n463 ) , .ZN( us02_n814 ) );
  NAND2_X2 us02_U389 (.A2( us02_n440 ) , .A1( us02_n451 ) , .ZN( us02_n790 ) );
  NOR3_X1 us02_U39 (.A3( us02_n721 ) , .A1( us02_n722 ) , .ZN( us02_n739 ) , .A2( us02_n740 ) );
  NAND2_X2 us02_U390 (.A1( us02_n448 ) , .A2( us02_n463 ) , .ZN( us02_n723 ) );
  NAND2_X1 us02_U391 (.A2( us02_n440 ) , .A1( us02_n446 ) , .ZN( us02_n783 ) );
  NAND2_X2 us02_U392 (.A1( us02_n448 ) , .A2( us02_n459 ) , .ZN( us02_n791 ) );
  NAND2_X2 us02_U393 (.A2( us02_n459 ) , .A1( us02_n464 ) , .ZN( us02_n779 ) );
  NAND2_X1 us02_U394 (.A1( us02_n446 ) , .A2( us02_n447 ) , .ZN( us02_n785 ) );
  NOR2_X1 us02_U395 (.A2( sa02_6 ) , .A1( sa02_7 ) , .ZN( us02_n463 ) );
  NOR2_X1 us02_U396 (.A2( sa02_5 ) , .ZN( us02_n447 ) , .A1( us02_n846 ) );
  NOR2_X1 us02_U397 (.A2( sa02_7 ) , .ZN( us02_n459 ) , .A1( us02_n848 ) );
  NOR2_X1 us02_U398 (.A2( sa02_4 ) , .ZN( us02_n448 ) , .A1( us02_n847 ) );
  NOR2_X1 us02_U399 (.A2( sa02_4 ) , .A1( sa02_5 ) , .ZN( us02_n440 ) );
  NAND2_X1 us02_U4 (.A2( us02_n470 ) , .A1( us02_n471 ) , .ZN( us02_n816 ) );
  AOI221_X1 us02_U40 (.A( us02_n780 ) , .ZN( us02_n797 ) , .C2( us02_n836 ) , .B2( us02_n837 ) , .B1( us02_n864 ) , .C1( us02_n865 ) );
  NOR2_X1 us02_U400 (.A2( sa02_1 ) , .ZN( us02_n470 ) , .A1( us02_n825 ) );
  NOR2_X1 us02_U401 (.A2( sa02_2 ) , .A1( sa02_3 ) , .ZN( us02_n471 ) );
  NOR2_X1 us02_U402 (.A2( sa02_6 ) , .ZN( us02_n451 ) , .A1( us02_n857 ) );
  NOR2_X1 us02_U403 (.A2( sa02_2 ) , .ZN( us02_n460 ) , .A1( us02_n828 ) );
  NOR2_X1 us02_U404 (.A2( sa02_0 ) , .ZN( us02_n453 ) , .A1( us02_n826 ) );
  NOR2_X1 us02_U405 (.A2( sa02_0 ) , .A1( sa02_1 ) , .ZN( us02_n461 ) );
  NOR2_X1 us02_U406 (.A2( sa02_3 ) , .ZN( us02_n454 ) , .A1( us02_n827 ) );
  INV_X1 us02_U407 (.A( sa02_6 ) , .ZN( us02_n848 ) );
  INV_X1 us02_U408 (.A( sa02_1 ) , .ZN( us02_n826 ) );
  INV_X1 us02_U409 (.A( sa02_3 ) , .ZN( us02_n828 ) );
  NOR4_X1 us02_U41 (.A4( us02_n792 ) , .A3( us02_n793 ) , .A2( us02_n794 ) , .A1( us02_n795 ) , .ZN( us02_n796 ) );
  INV_X1 us02_U410 (.A( sa02_2 ) , .ZN( us02_n827 ) );
  INV_X1 us02_U411 (.A( sa02_0 ) , .ZN( us02_n825 ) );
  INV_X1 us02_U412 (.A( sa02_5 ) , .ZN( us02_n847 ) );
  INV_X1 us02_U413 (.A( sa02_7 ) , .ZN( us02_n857 ) );
  OAI221_X1 us02_U414 (.A( us02_n782 ) , .C2( us02_n783 ) , .B2( us02_n784 ) , .B1( us02_n785 ) , .ZN( us02_n795 ) , .C1( us02_n812 ) );
  OAI22_X1 us02_U415 (.ZN( us02_n587 ) , .A2( us02_n746 ) , .B2( us02_n761 ) , .A1( us02_n762 ) , .B1( us02_n783 ) );
  AOI21_X1 us02_U416 (.ZN( us02_n591 ) , .B1( us02_n727 ) , .B2( us02_n783 ) , .A( us02_n789 ) );
  OAI221_X1 us02_U417 (.A( us02_n695 ) , .ZN( us02_n702 ) , .C2( us02_n783 ) , .C1( us02_n784 ) , .B1( us02_n785 ) , .B2( us02_n805 ) );
  NAND2_X1 us02_U418 (.A1( us02_n728 ) , .A2( us02_n783 ) , .ZN( us02_n810 ) );
  AOI21_X1 us02_U419 (.ZN( us02_n622 ) , .B1( us02_n698 ) , .A( us02_n778 ) , .B2( us02_n783 ) );
  NOR4_X1 us02_U42 (.A4( us02_n775 ) , .A3( us02_n776 ) , .A1( us02_n777 ) , .ZN( us02_n798 ) , .A2( us02_n800 ) );
  OAI22_X1 us02_U420 (.ZN( us02_n680 ) , .A1( us02_n698 ) , .A2( us02_n729 ) , .B2( us02_n783 ) , .B1( us02_n816 ) );
  AOI21_X1 us02_U421 (.ZN( us02_n647 ) , .A( us02_n761 ) , .B2( us02_n783 ) , .B1( us02_n791 ) );
  OAI21_X1 us02_U422 (.A( us02_n612 ) , .ZN( us02_n615 ) , .B1( us02_n624 ) , .B2( us02_n783 ) );
  NOR2_X1 us02_U423 (.ZN( us02_n650 ) , .A1( us02_n783 ) , .A2( us02_n787 ) );
  NOR2_X1 us02_U424 (.ZN( us02_n552 ) , .A2( us02_n743 ) , .A1( us02_n783 ) );
  NOR2_X1 us02_U425 (.ZN( us02_n609 ) , .A1( us02_n783 ) , .A2( us02_n815 ) );
  OAI222_X1 us02_U426 (.A2( us02_n668 ) , .ZN( us02_n673 ) , .B1( us02_n746 ) , .B2( us02_n783 ) , .C2( us02_n787 ) , .C1( us02_n814 ) , .A1( us02_n816 ) );
  NOR2_X1 us02_U427 (.ZN( us02_n599 ) , .A2( us02_n696 ) , .A1( us02_n783 ) );
  INV_X1 us02_U428 (.A( us02_n783 ) , .ZN( us02_n860 ) );
  AOI221_X1 us02_U429 (.A( us02_n575 ) , .ZN( us02_n586 ) , .B2( us02_n830 ) , .C2( us02_n842 ) , .B1( us02_n853 ) , .C1( us02_n860 ) );
  NOR2_X1 us02_U43 (.ZN( us02_n803 ) , .A1( us02_n853 ) , .A2( us02_n860 ) );
  AOI21_X1 us02_U430 (.ZN( us02_n575 ) , .B2( us02_n723 ) , .B1( us02_n747 ) , .A( us02_n784 ) );
  INV_X1 us02_U431 (.A( sa02_4 ) , .ZN( us02_n846 ) );
  NAND2_X1 us02_U432 (.ZN( sa02_sr_2 ) , .A2( us02_n438 ) , .A1( us02_n644 ) );
  NOR3_X1 us02_U433 (.A2( us02_n606 ) , .A1( us02_n607 ) , .ZN( us02_n645 ) , .A3( us02_n721 ) );
  AOI222_X1 us02_U434 (.B2( us02_n637 ) , .ZN( us02_n643 ) , .B1( us02_n840 ) , .A1( us02_n841 ) , .C2( us02_n845 ) , .C1( us02_n862 ) , .A2( us02_n864 ) );
  NOR4_X1 us02_U435 (.A4( us02_n638 ) , .A3( us02_n639 ) , .A2( us02_n640 ) , .A1( us02_n641 ) , .ZN( us02_n642 ) );
  AOI211_X1 us02_U436 (.A( us02_n636 ) , .ZN( us02_n644 ) , .B( us02_n742 ) , .C2( us02_n838 ) , .C1( us02_n853 ) );
  NAND3_X1 us02_U437 (.ZN( sa02_sr_6 ) , .A3( us02_n796 ) , .A2( us02_n797 ) , .A1( us02_n798 ) );
  NAND3_X1 us02_U438 (.ZN( sa02_sr_5 ) , .A3( us02_n757 ) , .A2( us02_n758 ) , .A1( us02_n759 ) );
  NAND3_X1 us02_U439 (.ZN( sa02_sr_4 ) , .A3( us02_n737 ) , .A2( us02_n738 ) , .A1( us02_n739 ) );
  NAND4_X1 us02_U44 (.ZN( sa02_sr_3 ) , .A4( us02_n703 ) , .A3( us02_n704 ) , .A2( us02_n705 ) , .A1( us02_n706 ) );
  NAND3_X1 us02_U440 (.A3( us02_n674 ) , .A2( us02_n675 ) , .A1( us02_n676 ) , .ZN( us02_n806 ) );
  NAND3_X1 us02_U441 (.ZN( us02_n637 ) , .A3( us02_n707 ) , .A2( us02_n723 ) , .A1( us02_n791 ) );
  NAND3_X1 us02_U442 (.A3( us02_n617 ) , .A2( us02_n618 ) , .A1( us02_n619 ) , .ZN( us02_n724 ) );
  NAND3_X1 us02_U443 (.A3( us02_n584 ) , .A2( us02_n585 ) , .A1( us02_n586 ) , .ZN( us02_n620 ) );
  NAND3_X1 us02_U444 (.ZN( us02_n564 ) , .A3( us02_n679 ) , .A2( us02_n749 ) , .A1( us02_n784 ) );
  NAND3_X1 us02_U445 (.A3( us02_n522 ) , .A2( us02_n523 ) , .A1( us02_n524 ) , .ZN( us02_n741 ) );
  NAND3_X1 us02_U446 (.A3( us02_n511 ) , .A1( us02_n512 ) , .ZN( us02_n607 ) , .A2( us02_n870 ) );
  NAND3_X1 us02_U447 (.A3( us02_n466 ) , .A2( us02_n467 ) , .A1( us02_n468 ) , .ZN( us02_n776 ) );
  NAND4_X1 us02_U448 (.A4( us02_n632 ) , .A3( us02_n633 ) , .A2( us02_n634 ) , .A1( us02_n635 ) , .ZN( us02_n742 ) );
  NOR4_X1 us02_U45 (.A4( us02_n699 ) , .A3( us02_n700 ) , .A2( us02_n701 ) , .A1( us02_n702 ) , .ZN( us02_n703 ) );
  AOI211_X1 us02_U46 (.B( us02_n693 ) , .A( us02_n694 ) , .ZN( us02_n704 ) , .C2( us02_n830 ) , .C1( us02_n850 ) );
  NOR2_X1 us02_U47 (.ZN( us02_n706 ) , .A2( us02_n775 ) , .A1( us02_n799 ) );
  NAND4_X1 us02_U48 (.ZN( sa02_sr_7 ) , .A4( us02_n821 ) , .A3( us02_n822 ) , .A2( us02_n823 ) , .A1( us02_n824 ) );
  NOR4_X1 us02_U49 (.A4( us02_n817 ) , .A3( us02_n818 ) , .A2( us02_n819 ) , .A1( us02_n820 ) , .ZN( us02_n821 ) );
  NOR3_X1 us02_U5 (.ZN( us02_n597 ) , .A1( us02_n607 ) , .A3( us02_n722 ) , .A2( us02_n741 ) );
  AOI222_X1 us02_U50 (.C2( us02_n808 ) , .B2( us02_n809 ) , .A2( us02_n810 ) , .ZN( us02_n822 ) , .C1( us02_n831 ) , .A1( us02_n838 ) , .B1( us02_n852 ) );
  AOI211_X1 us02_U51 (.B( us02_n806 ) , .A( us02_n807 ) , .ZN( us02_n823 ) , .C1( us02_n841 ) , .C2( us02_n849 ) );
  NOR2_X1 us02_U52 (.ZN( us02_n747 ) , .A1( us02_n860 ) , .A2( us02_n861 ) );
  NAND4_X1 us02_U53 (.ZN( sa02_sr_0 ) , .A4( us02_n500 ) , .A3( us02_n501 ) , .A2( us02_n502 ) , .A1( us02_n503 ) );
  AOI221_X1 us02_U54 (.A( us02_n496 ) , .ZN( us02_n501 ) , .B2( us02_n842 ) , .C1( us02_n845 ) , .C2( us02_n859 ) , .B1( us02_n861 ) );
  NOR4_X1 us02_U55 (.A4( us02_n497 ) , .A3( us02_n498 ) , .A2( us02_n499 ) , .ZN( us02_n500 ) , .A1( us02_n526 ) );
  AOI211_X1 us02_U56 (.A( us02_n495 ) , .ZN( us02_n502 ) , .B( us02_n801 ) , .C2( us02_n838 ) , .C1( us02_n850 ) );
  NAND4_X1 us02_U57 (.ZN( sa02_sr_1 ) , .A4( us02_n594 ) , .A3( us02_n595 ) , .A2( us02_n596 ) , .A1( us02_n597 ) );
  NOR4_X1 us02_U58 (.A4( us02_n590 ) , .A3( us02_n591 ) , .A2( us02_n592 ) , .A1( us02_n593 ) , .ZN( us02_n594 ) );
  AOI211_X1 us02_U59 (.B( us02_n588 ) , .A( us02_n589 ) , .ZN( us02_n595 ) , .C2( us02_n810 ) , .C1( us02_n832 ) );
  NOR3_X1 us02_U6 (.A3( us02_n799 ) , .A2( us02_n800 ) , .A1( us02_n801 ) , .ZN( us02_n824 ) );
  AOI211_X1 us02_U60 (.A( us02_n587 ) , .ZN( us02_n596 ) , .B( us02_n620 ) , .C1( us02_n844 ) , .C2( us02_n854 ) );
  NOR2_X1 us02_U61 (.ZN( us02_n624 ) , .A2( us02_n835 ) , .A1( us02_n838 ) );
  AND3_X1 us02_U62 (.ZN( us02_n438 ) , .A2( us02_n642 ) , .A3( us02_n643 ) , .A1( us02_n645 ) );
  NOR4_X1 us02_U63 (.A4( us02_n576 ) , .A3( us02_n577 ) , .A2( us02_n578 ) , .ZN( us02_n585 ) , .A1( us02_n682 ) );
  NOR4_X1 us02_U64 (.A1( us02_n583 ) , .ZN( us02_n584 ) , .A3( us02_n651 ) , .A2( us02_n661 ) , .A4( us02_n766 ) );
  AOI211_X1 us02_U65 (.B( us02_n622 ) , .A( us02_n623 ) , .ZN( us02_n634 ) , .C2( us02_n835 ) , .C1( us02_n862 ) );
  NOR4_X1 us02_U66 (.A4( us02_n628 ) , .A3( us02_n629 ) , .A2( us02_n630 ) , .A1( us02_n631 ) , .ZN( us02_n632 ) );
  NOR4_X1 us02_U67 (.A4( us02_n625 ) , .A3( us02_n626 ) , .A2( us02_n627 ) , .ZN( us02_n633 ) , .A1( us02_n663 ) );
  NAND4_X1 us02_U68 (.A4( us02_n656 ) , .A3( us02_n657 ) , .A2( us02_n658 ) , .A1( us02_n659 ) , .ZN( us02_n799 ) );
  NOR3_X1 us02_U69 (.A3( us02_n647 ) , .A2( us02_n648 ) , .A1( us02_n649 ) , .ZN( us02_n658 ) );
  NOR3_X1 us02_U7 (.ZN( us02_n503 ) , .A2( us02_n678 ) , .A3( us02_n776 ) , .A1( us02_n875 ) );
  NOR3_X1 us02_U70 (.A3( us02_n650 ) , .A2( us02_n651 ) , .A1( us02_n652 ) , .ZN( us02_n657 ) );
  NOR3_X1 us02_U71 (.A3( us02_n653 ) , .A2( us02_n654 ) , .A1( us02_n655 ) , .ZN( us02_n656 ) );
  NAND4_X1 us02_U72 (.A4( us02_n771 ) , .A3( us02_n772 ) , .A2( us02_n773 ) , .A1( us02_n774 ) , .ZN( us02_n800 ) );
  NOR3_X1 us02_U73 (.A3( us02_n764 ) , .A2( us02_n765 ) , .A1( us02_n766 ) , .ZN( us02_n772 ) );
  NOR4_X1 us02_U74 (.A4( us02_n767 ) , .A3( us02_n768 ) , .A2( us02_n769 ) , .A1( us02_n770 ) , .ZN( us02_n771 ) );
  AOI222_X1 us02_U75 (.ZN( us02_n774 ) , .A1( us02_n829 ) , .C1( us02_n833 ) , .B2( us02_n840 ) , .A2( us02_n849 ) , .B1( us02_n860 ) , .C2( us02_n872 ) );
  NOR4_X1 us02_U76 (.A4( us02_n664 ) , .A3( us02_n665 ) , .A2( us02_n666 ) , .A1( us02_n667 ) , .ZN( us02_n675 ) );
  NOR4_X1 us02_U77 (.A4( us02_n660 ) , .A3( us02_n661 ) , .A2( us02_n662 ) , .A1( us02_n663 ) , .ZN( us02_n676 ) );
  NOR4_X1 us02_U78 (.A3( us02_n672 ) , .A1( us02_n673 ) , .ZN( us02_n674 ) , .A4( us02_n714 ) , .A2( us02_n858 ) );
  NOR2_X1 us02_U79 (.ZN( us02_n760 ) , .A1( us02_n832 ) , .A2( us02_n833 ) );
  INV_X1 us02_U8 (.A( us02_n705 ) , .ZN( us02_n875 ) );
  NAND4_X1 us02_U80 (.A4( us02_n455 ) , .A3( us02_n456 ) , .A2( us02_n457 ) , .A1( us02_n458 ) , .ZN( us02_n678 ) );
  NOR3_X1 us02_U81 (.ZN( us02_n456 ) , .A3( us02_n529 ) , .A1( us02_n554 ) , .A2( us02_n569 ) );
  AOI221_X1 us02_U82 (.A( us02_n449 ) , .ZN( us02_n458 ) , .C2( us02_n752 ) , .B1( us02_n831 ) , .C1( us02_n841 ) , .B2( us02_n860 ) );
  NOR4_X1 us02_U83 (.ZN( us02_n457 ) , .A2( us02_n508 ) , .A1( us02_n598 ) , .A4( us02_n627 ) , .A3( us02_n710 ) );
  NAND4_X1 us02_U84 (.A4( us02_n602 ) , .A3( us02_n603 ) , .A2( us02_n604 ) , .A1( us02_n605 ) , .ZN( us02_n721 ) );
  NOR3_X1 us02_U85 (.A1( us02_n598 ) , .ZN( us02_n603 ) , .A3( us02_n662 ) , .A2( us02_n769 ) );
  NOR4_X1 us02_U86 (.A3( us02_n599 ) , .A2( us02_n600 ) , .A1( us02_n601 ) , .ZN( us02_n602 ) , .A4( us02_n654 ) );
  AOI222_X1 us02_U87 (.ZN( us02_n605 ) , .A1( us02_n829 ) , .C2( us02_n836 ) , .B1( us02_n841 ) , .A2( us02_n855 ) , .B2( us02_n860 ) , .C1( us02_n867 ) );
  NAND4_X1 us02_U88 (.A4( us02_n534 ) , .A3( us02_n535 ) , .A2( us02_n536 ) , .A1( us02_n537 ) , .ZN( us02_n621 ) );
  NOR4_X1 us02_U89 (.A4( us02_n525 ) , .A2( us02_n526 ) , .A1( us02_n527 ) , .ZN( us02_n537 ) , .A3( us02_n700 ) );
  NOR3_X1 us02_U9 (.A3( us02_n620 ) , .A2( us02_n621 ) , .ZN( us02_n635 ) , .A1( us02_n724 ) );
  NOR4_X1 us02_U90 (.A1( us02_n530 ) , .ZN( us02_n535 ) , .A2( us02_n653 ) , .A4( us02_n667 ) , .A3( us02_n764 ) );
  NOR4_X1 us02_U91 (.A4( us02_n528 ) , .A3( us02_n529 ) , .ZN( us02_n536 ) , .A2( us02_n683 ) , .A1( us02_n793 ) );
  NAND4_X1 us02_U92 (.A4( us02_n547 ) , .A3( us02_n548 ) , .A2( us02_n549 ) , .A1( us02_n550 ) , .ZN( us02_n744 ) );
  NOR3_X1 us02_U93 (.ZN( us02_n548 ) , .A2( us02_n650 ) , .A1( us02_n666 ) , .A3( us02_n770 ) );
  AOI211_X1 us02_U94 (.B( us02_n538 ) , .A( us02_n539 ) , .ZN( us02_n550 ) , .C2( us02_n838 ) , .C1( us02_n850 ) );
  NOR4_X1 us02_U95 (.A4( us02_n543 ) , .A3( us02_n544 ) , .A2( us02_n545 ) , .A1( us02_n546 ) , .ZN( us02_n547 ) );
  NAND4_X1 us02_U96 (.A4( us02_n478 ) , .A3( us02_n479 ) , .A2( us02_n480 ) , .A1( us02_n481 ) , .ZN( us02_n693 ) );
  NOR3_X1 us02_U97 (.ZN( us02_n479 ) , .A2( us02_n507 ) , .A3( us02_n600 ) , .A1( us02_n609 ) );
  AOI211_X1 us02_U98 (.B( us02_n476 ) , .A( us02_n477 ) , .ZN( us02_n481 ) , .C2( us02_n832 ) , .C1( us02_n860 ) );
  NOR4_X1 us02_U99 (.ZN( us02_n480 ) , .A3( us02_n531 ) , .A4( us02_n544 ) , .A2( us02_n566 ) , .A1( us02_n716 ) );
endmodule

