module des_des_die_6 ( u0_K14_10, u0_K14_12, u0_K14_13, u0_K14_14, u0_K14_15, u0_K14_18, u0_K14_21, u0_K14_24, u0_K14_27, 
       u0_K14_4, u0_K14_9, u0_K1_13, u0_K1_14, u0_K1_15, u0_K1_16, u0_K1_17, u0_K1_23, u0_K5_13, 
       u0_K5_14, u0_K5_15, u0_K5_16, u0_K5_18, u0_K5_19, u0_K5_23, u0_K5_24, u0_K5_9, u0_L12_1, 
       u0_L12_10, u0_L12_11, u0_L12_13, u0_L12_14, u0_L12_16, u0_L12_17, u0_L12_18, u0_L12_19, u0_L12_2, 
       u0_L12_20, u0_L12_23, u0_L12_24, u0_L12_25, u0_L12_26, u0_L12_28, u0_L12_29, u0_L12_3, u0_L12_30, 
       u0_L12_31, u0_L12_4, u0_L12_6, u0_L12_8, u0_L12_9, u0_L3_1, u0_L3_10, u0_L3_13, u0_L3_16, 
       u0_L3_18, u0_L3_2, u0_L3_20, u0_L3_24, u0_L3_26, u0_L3_28, u0_L3_30, u0_L3_6, u0_R12_1, 
       u0_R12_10, u0_R12_11, u0_R12_12, u0_R12_13, u0_R12_14, u0_R12_15, u0_R12_16, u0_R12_17, u0_R12_18, 
       u0_R12_19, u0_R12_2, u0_R12_20, u0_R12_21, u0_R12_22, u0_R12_23, u0_R12_24, u0_R12_25, u0_R12_3, 
       u0_R12_32, u0_R12_4, u0_R12_5, u0_R12_6, u0_R12_7, u0_R12_8, u0_R12_9, u0_R3_10, u0_R3_11, 
       u0_R3_12, u0_R3_13, u0_R3_14, u0_R3_15, u0_R3_16, u0_R3_17, u0_R3_4, u0_R3_5, u0_R3_6, 
       u0_R3_7, u0_R3_8, u0_R3_9, u0_desIn_r_10, u0_desIn_r_12, u0_desIn_r_13, u0_desIn_r_14, u0_desIn_r_15, u0_desIn_r_2, 
       u0_desIn_r_21, u0_desIn_r_23, u0_desIn_r_24, u0_desIn_r_26, u0_desIn_r_29, u0_desIn_r_3, u0_desIn_r_31, u0_desIn_r_36, u0_desIn_r_37, 
       u0_desIn_r_39, u0_desIn_r_4, u0_desIn_r_40, u0_desIn_r_45, u0_desIn_r_46, u0_desIn_r_47, u0_desIn_r_48, u0_desIn_r_5, u0_desIn_r_50, 
       u0_desIn_r_53, u0_desIn_r_55, u0_desIn_r_57, u0_desIn_r_58, u0_desIn_r_6, u0_desIn_r_60, u0_desIn_r_61, u0_desIn_r_63, u0_desIn_r_7, 
       u0_desIn_r_8, u0_key_r_11, u0_key_r_12, u0_key_r_13, u0_key_r_17, u0_key_r_19, u0_key_r_20, u0_key_r_24, u0_key_r_25, 
       u0_key_r_26, u0_key_r_27, u0_key_r_3, u0_key_r_32, u0_key_r_34, u0_key_r_39, u0_key_r_4, u0_key_r_40, u0_key_r_41, 
       u0_key_r_47, u0_key_r_48, u0_key_r_49, u0_key_r_5, u0_key_r_53, u0_key_r_54, u0_key_r_55, u0_key_r_6, u0_uk_K_r12_1, 
       u0_uk_K_r12_10, u0_uk_K_r12_25, u0_uk_K_r12_30, u0_uk_K_r12_33, u0_uk_K_r12_36, u0_uk_K_r12_44, u0_uk_K_r12_47, u0_uk_K_r12_7, u0_uk_K_r3_11, 
       u0_uk_K_r3_19, u0_uk_K_r3_24, u0_uk_K_r3_47, u0_uk_n10, u0_uk_n100, u0_uk_n109, u0_uk_n11, u0_uk_n110, u0_uk_n117, 
       u0_uk_n118, u0_uk_n128, u0_uk_n129, u0_uk_n141, u0_uk_n142, u0_uk_n145, u0_uk_n146, u0_uk_n147, u0_uk_n163, 
       u0_uk_n164, u0_uk_n17, u0_uk_n182, u0_uk_n187, u0_uk_n188, u0_uk_n202, u0_uk_n203, u0_uk_n207, u0_uk_n208, 
       u0_uk_n213, u0_uk_n217, u0_uk_n220, u0_uk_n222, u0_uk_n230, u0_uk_n231, u0_uk_n240, u0_uk_n242, u0_uk_n250, 
       u0_uk_n251, u0_uk_n257, u0_uk_n451, u0_uk_n453, u0_uk_n459, u0_uk_n46, u0_uk_n464, u0_uk_n465, u0_uk_n473, 
       u0_uk_n479, u0_uk_n48, u0_uk_n483, u0_uk_n484, u0_uk_n485, u0_uk_n489, u0_uk_n49, u0_uk_n50, u0_uk_n51, 
       u0_uk_n53, u0_uk_n54, u0_uk_n55, u0_uk_n57, u0_uk_n61, u0_uk_n62, u0_uk_n63, u0_uk_n64, u0_uk_n66, 
       u0_uk_n67, u0_uk_n69, u0_uk_n72, u0_uk_n73, u0_uk_n75, u0_uk_n77, u0_uk_n78, u0_uk_n79, u0_uk_n80, 
       u0_uk_n815, u0_uk_n82, u0_uk_n83, u0_uk_n84, u0_uk_n85, u0_uk_n86, u0_uk_n87, u0_uk_n88, u0_uk_n89, 
       u0_uk_n92, u0_uk_n93, u0_uk_n94, u0_uk_n99, u2_FP_33, u2_FP_34, u2_FP_35, u2_FP_36, u2_FP_37, 
       u2_FP_48, u2_FP_49, u2_FP_50, u2_FP_51, u2_FP_52, u2_FP_53, u2_FP_54, u2_FP_55, u2_FP_56, 
       u2_FP_57, u2_FP_58, u2_FP_59, u2_FP_60, u2_FP_61, u2_FP_62, u2_FP_63, u2_FP_64, u2_K10_10, 
       u2_K10_11, u2_K10_15, u2_K10_17, u2_K10_4, u2_K10_43, u2_K10_44, u2_K10_46, u2_K10_6, u2_K12_2, 
       u2_K12_8, u2_K14_25, u2_K14_28, u2_K15_1, u2_K15_2, u2_K15_28, u2_K15_29, u2_K15_31, u2_K15_34, 
       u2_K15_35, u2_K15_39, u2_K15_5, u2_K16_26, u2_K16_31, u2_K16_42, u2_K16_44, u2_K16_47, u2_K16_5, 
       u2_K16_6, u2_K1_15, u2_K1_16, u2_K1_19, u2_K1_24, u2_K1_5, u2_K1_9, u2_K2_40, u2_K3_13, 
       u2_K3_15, u2_K3_16, u2_K3_20, u2_K3_23, u2_K3_32, u2_K3_35, u2_K3_42, u2_K3_43, u2_K3_47, 
       u2_K3_48, u2_K3_7, u2_K4_14, u2_K4_21, u2_K4_22, u2_K4_27, u2_K4_33, u2_K4_34, u2_K4_35, 
       u2_K5_10, u2_K5_11, u2_K5_13, u2_K5_14, u2_K5_16, u2_K5_17, u2_K5_18, u2_K5_19, u2_K5_21, 
       u2_K5_23, u2_K5_24, u2_K5_8, u2_K5_9, u2_K6_20, u2_K6_22, u2_K6_24, u2_K6_25, u2_K6_27, 
       u2_K7_26, u2_K7_3, u2_K7_37, u2_K7_38, u2_K7_4, u2_K7_43, u2_K7_45, u2_K7_48, u2_K7_5, 
       u2_K7_7, u2_K8_41, u2_K8_45, u2_L0_12, u2_L0_14, u2_L0_22, u2_L0_25, u2_L0_3, u2_L0_32, 
       u2_L0_7, u2_L0_8, u2_L10_13, u2_L10_16, u2_L10_17, u2_L10_18, u2_L10_2, u2_L10_23, u2_L10_24, 
       u2_L10_28, u2_L10_30, u2_L10_31, u2_L10_6, u2_L10_9, u2_L12_11, u2_L12_14, u2_L12_19, u2_L12_25, 
       u2_L12_29, u2_L12_3, u2_L12_4, u2_L12_8, u2_L13_11, u2_L13_12, u2_L13_13, u2_L13_14, u2_L13_17, 
       u2_L13_18, u2_L13_19, u2_L13_2, u2_L13_22, u2_L13_23, u2_L13_25, u2_L13_28, u2_L13_29, u2_L13_3, 
       u2_L13_31, u2_L13_32, u2_L13_4, u2_L13_7, u2_L13_8, u2_L13_9, u2_L14_11, u2_L14_12, u2_L14_14, 
       u2_L14_15, u2_L14_17, u2_L14_19, u2_L14_21, u2_L14_22, u2_L14_23, u2_L14_25, u2_L14_27, u2_L14_29, 
       u2_L14_3, u2_L14_31, u2_L14_32, u2_L14_4, u2_L14_5, u2_L14_7, u2_L14_8, u2_L14_9, u2_L1_1, 
       u2_L1_10, u2_L1_11, u2_L1_12, u2_L1_13, u2_L1_15, u2_L1_16, u2_L1_17, u2_L1_18, u2_L1_19, 
       u2_L1_2, u2_L1_20, u2_L1_21, u2_L1_22, u2_L1_23, u2_L1_24, u2_L1_26, u2_L1_27, u2_L1_28, 
       u2_L1_29, u2_L1_30, u2_L1_31, u2_L1_32, u2_L1_4, u2_L1_5, u2_L1_6, u2_L1_7, u2_L1_9, 
       u2_L2_1, u2_L2_10, u2_L2_11, u2_L2_14, u2_L2_16, u2_L2_19, u2_L2_20, u2_L2_24, u2_L2_25, 
       u2_L2_26, u2_L2_29, u2_L2_3, u2_L2_30, u2_L2_4, u2_L2_6, u2_L2_8, u2_L3_1, u2_L3_10, 
       u2_L3_13, u2_L3_16, u2_L3_18, u2_L3_2, u2_L3_20, u2_L3_24, u2_L3_26, u2_L3_28, u2_L3_30, 
       u2_L3_6, u2_L4_1, u2_L4_10, u2_L4_14, u2_L4_20, u2_L4_25, u2_L4_26, u2_L4_3, u2_L4_8, 
       u2_L5_1, u2_L5_10, u2_L5_12, u2_L5_13, u2_L5_14, u2_L5_15, u2_L5_16, u2_L5_17, u2_L5_18, 
       u2_L5_2, u2_L5_20, u2_L5_21, u2_L5_22, u2_L5_23, u2_L5_24, u2_L5_25, u2_L5_26, u2_L5_27, 
       u2_L5_28, u2_L5_3, u2_L5_30, u2_L5_31, u2_L5_32, u2_L5_5, u2_L5_6, u2_L5_7, u2_L5_8, 
       u2_L5_9, u2_L6_12, u2_L6_15, u2_L6_21, u2_L6_22, u2_L6_27, u2_L6_32, u2_L6_5, u2_L6_7, 
       u2_L8_13, u2_L8_15, u2_L8_16, u2_L8_17, u2_L8_18, u2_L8_2, u2_L8_21, u2_L8_23, u2_L8_24, 
       u2_L8_27, u2_L8_28, u2_L8_30, u2_L8_31, u2_L8_5, u2_L8_6, u2_L8_9, u2_R0_16, u2_R0_17, 
       u2_R0_18, u2_R0_19, u2_R0_20, u2_R0_21, u2_R0_24, u2_R0_25, u2_R0_26, u2_R0_27, u2_R0_28, 
       u2_R0_29, u2_R10_1, u2_R10_10, u2_R10_11, u2_R10_12, u2_R10_13, u2_R10_2, u2_R10_3, u2_R10_32, 
       u2_R10_4, u2_R10_5, u2_R10_6, u2_R10_7, u2_R10_8, u2_R10_9, u2_R12_16, u2_R12_17, u2_R12_18, 
       u2_R12_19, u2_R12_20, u2_R12_21, u2_R12_22, u2_R12_23, u2_R12_24, u2_R12_25, u2_R13_1, u2_R13_16, 
       u2_R13_17, u2_R13_18, u2_R13_19, u2_R13_2, u2_R13_20, u2_R13_21, u2_R13_22, u2_R13_23, u2_R13_24, 
       u2_R13_25, u2_R13_26, u2_R13_27, u2_R13_28, u2_R13_29, u2_R13_3, u2_R13_32, u2_R13_4, u2_R13_5, 
       u2_R13_6, u2_R13_7, u2_R13_8, u2_R13_9, u2_R1_1, u2_R1_10, u2_R1_11, u2_R1_12, u2_R1_13, 
       u2_R1_14, u2_R1_15, u2_R1_16, u2_R1_17, u2_R1_2, u2_R1_20, u2_R1_21, u2_R1_22, u2_R1_23, 
       u2_R1_24, u2_R1_25, u2_R1_26, u2_R1_27, u2_R1_28, u2_R1_29, u2_R1_3, u2_R1_30, u2_R1_31, 
       u2_R1_32, u2_R1_4, u2_R1_5, u2_R1_6, u2_R1_7, u2_R1_8, u2_R1_9, u2_R2_10, u2_R2_11, 
       u2_R2_12, u2_R2_13, u2_R2_14, u2_R2_15, u2_R2_16, u2_R2_17, u2_R2_18, u2_R2_19, u2_R2_20, 
       u2_R2_21, u2_R2_22, u2_R2_23, u2_R2_24, u2_R2_25, u2_R2_8, u2_R2_9, u2_R3_10, u2_R3_11, 
       u2_R3_12, u2_R3_13, u2_R3_14, u2_R3_15, u2_R3_16, u2_R3_17, u2_R3_4, u2_R3_5, u2_R3_6, 
       u2_R3_7, u2_R3_8, u2_R3_9, u2_R4_12, u2_R4_13, u2_R4_14, u2_R4_15, u2_R4_16, u2_R4_17, 
       u2_R4_18, u2_R4_19, u2_R4_20, u2_R4_21, u2_R5_1, u2_R5_10, u2_R5_11, u2_R5_12, u2_R5_13, 
       u2_R5_14, u2_R5_15, u2_R5_16, u2_R5_17, u2_R5_18, u2_R5_19, u2_R5_2, u2_R5_20, u2_R5_21, 
       u2_R5_24, u2_R5_25, u2_R5_26, u2_R5_27, u2_R5_28, u2_R5_29, u2_R5_3, u2_R5_30, u2_R5_31, 
       u2_R5_32, u2_R5_4, u2_R5_5, u2_R5_6, u2_R5_7, u2_R5_8, u2_R5_9, u2_R6_1, u2_R6_24, 
       u2_R6_25, u2_R6_26, u2_R6_27, u2_R6_28, u2_R6_29, u2_R6_30, u2_R6_31, u2_R6_32, u2_R8_1, 
       u2_R8_10, u2_R8_11, u2_R8_12, u2_R8_13, u2_R8_2, u2_R8_28, u2_R8_29, u2_R8_3, u2_R8_30, 
       u2_R8_31, u2_R8_32, u2_R8_4, u2_R8_5, u2_R8_6, u2_R8_7, u2_R8_8, u2_R8_9, u2_desIn_r_10, 
       u2_desIn_r_12, u2_desIn_r_13, u2_desIn_r_14, u2_desIn_r_15, u2_desIn_r_2, u2_desIn_r_21, u2_desIn_r_23, u2_desIn_r_24, u2_desIn_r_26, 
       u2_desIn_r_29, u2_desIn_r_3, u2_desIn_r_31, u2_desIn_r_36, u2_desIn_r_37, u2_desIn_r_39, u2_desIn_r_4, u2_desIn_r_40, u2_desIn_r_45, 
       u2_desIn_r_46, u2_desIn_r_47, u2_desIn_r_48, u2_desIn_r_5, u2_desIn_r_50, u2_desIn_r_53, u2_desIn_r_55, u2_desIn_r_57, u2_desIn_r_58, 
       u2_desIn_r_6, u2_desIn_r_60, u2_desIn_r_61, u2_desIn_r_63, u2_desIn_r_7, u2_desIn_r_8, u2_key_r_10, u2_key_r_11, u2_key_r_12, 
       u2_key_r_17, u2_key_r_19, u2_key_r_20, u2_key_r_24, u2_key_r_25, u2_key_r_26, u2_key_r_27, u2_key_r_3, u2_key_r_32, 
       u2_key_r_33, u2_key_r_34, u2_key_r_4, u2_key_r_40, u2_key_r_41, u2_key_r_46, u2_key_r_47, u2_key_r_48, u2_key_r_49, 
       u2_key_r_50, u2_key_r_53, u2_key_r_55, u2_key_r_6, u2_uk_K_r0_15, u2_uk_K_r0_49, u2_uk_K_r10_10, u2_uk_K_r10_25, u2_uk_K_r10_27, 
       u2_uk_K_r10_34, u2_uk_K_r10_4, u2_uk_K_r11_7, u2_uk_K_r12_1, u2_uk_K_r12_30, u2_uk_K_r12_36, u2_uk_K_r12_42, u2_uk_K_r12_7, u2_uk_K_r13_0, 
       u2_uk_K_r13_13, u2_uk_K_r13_17, u2_uk_K_r13_22, u2_uk_K_r13_25, u2_uk_K_r13_38, u2_uk_K_r13_55, u2_uk_K_r14_15, u2_uk_K_r14_16, u2_uk_K_r14_2, 
       u2_uk_K_r14_3, u2_uk_K_r14_45, u2_uk_K_r14_50, u2_uk_K_r14_9, u2_uk_K_r1_15, u2_uk_K_r1_16, u2_uk_K_r1_17, u2_uk_K_r1_18, u2_uk_K_r1_21, 
       u2_uk_K_r1_22, u2_uk_K_r1_41, u2_uk_K_r1_47, u2_uk_K_r1_7, u2_uk_K_r2_18, u2_uk_K_r2_21, u2_uk_K_r2_27, u2_uk_K_r2_28, u2_uk_K_r2_31, 
       u2_uk_K_r2_36, u2_uk_K_r2_49, u2_uk_K_r2_55, u2_uk_K_r3_11, u2_uk_K_r3_19, u2_uk_K_r4_0, u2_uk_K_r4_11, u2_uk_K_r4_35, u2_uk_K_r4_5, 
       u2_uk_K_r5_10, u2_uk_K_r5_16, u2_uk_K_r5_17, u2_uk_K_r5_18, u2_uk_K_r5_19, u2_uk_K_r5_23, u2_uk_K_r5_26, u2_uk_K_r5_31, u2_uk_K_r5_37, 
       u2_uk_K_r5_39, u2_uk_K_r5_4, u2_uk_K_r5_40, u2_uk_K_r5_41, u2_uk_K_r5_43, u2_uk_K_r5_48, u2_uk_K_r5_7, u2_uk_K_r6_0, u2_uk_K_r6_14, 
       u2_uk_K_r6_31, u2_uk_K_r6_37, u2_uk_K_r6_46, u2_uk_K_r6_7, u2_uk_K_r8_17, u2_uk_K_r8_21, u2_uk_K_r8_27, u2_uk_K_r8_32, u2_uk_K_r8_41, 
       u2_uk_K_r8_48, u2_uk_K_r9_0, u2_uk_n1001, u2_uk_n1007, u2_uk_n1011, u2_uk_n1018, u2_uk_n102, u2_uk_n1022, u2_uk_n1024, 
       u2_uk_n1027, u2_uk_n1028, u2_uk_n1042, u2_uk_n1043, u2_uk_n1044, u2_uk_n1061, u2_uk_n1063, u2_uk_n1077, u2_uk_n1079, 
       u2_uk_n1081, u2_uk_n1082, u2_uk_n109, u2_uk_n1093, u2_uk_n1094, u2_uk_n1096, u2_uk_n110, u2_uk_n1112, u2_uk_n1113, 
       u2_uk_n1188, u2_uk_n1189, u2_uk_n1190, u2_uk_n1195, u2_uk_n1198, u2_uk_n1200, u2_uk_n1201, u2_uk_n1203, u2_uk_n1206, 
       u2_uk_n1208, u2_uk_n1209, u2_uk_n1210, u2_uk_n1215, u2_uk_n1216, u2_uk_n1217, u2_uk_n1218, u2_uk_n1220, u2_uk_n1221, 
       u2_uk_n1223, u2_uk_n1225, u2_uk_n1226, u2_uk_n1227, u2_uk_n1230, u2_uk_n1236, u2_uk_n1237, u2_uk_n1246, u2_uk_n1251, 
       u2_uk_n1252, u2_uk_n1259, u2_uk_n1264, u2_uk_n1265, u2_uk_n1266, u2_uk_n1274, u2_uk_n1279, u2_uk_n128, u2_uk_n1280, 
       u2_uk_n1281, u2_uk_n1282, u2_uk_n1283, u2_uk_n1284, u2_uk_n1285, u2_uk_n1286, u2_uk_n1287, u2_uk_n1288, u2_uk_n1290, 
       u2_uk_n1291, u2_uk_n1292, u2_uk_n1293, u2_uk_n1294, u2_uk_n1295, u2_uk_n1296, u2_uk_n1297, u2_uk_n1298, u2_uk_n1299, 
       u2_uk_n1300, u2_uk_n1301, u2_uk_n1302, u2_uk_n1303, u2_uk_n1305, u2_uk_n1306, u2_uk_n1308, u2_uk_n1309, u2_uk_n1310, 
       u2_uk_n1311, u2_uk_n1312, u2_uk_n1314, u2_uk_n1316, u2_uk_n1317, u2_uk_n1318, u2_uk_n1322, u2_uk_n1324, u2_uk_n1326, 
       u2_uk_n1328, u2_uk_n1329, u2_uk_n1333, u2_uk_n1335, u2_uk_n1339, u2_uk_n1345, u2_uk_n1346, u2_uk_n1347, u2_uk_n1348, 
       u2_uk_n1350, u2_uk_n1351, u2_uk_n1356, u2_uk_n1363, u2_uk_n1375, u2_uk_n1379, u2_uk_n1405, u2_uk_n1408, u2_uk_n1412, 
       u2_uk_n1413, u2_uk_n1414, u2_uk_n1420, u2_uk_n1439, u2_uk_n1442, u2_uk_n1447, u2_uk_n145, u2_uk_n1452, u2_uk_n1453, 
       u2_uk_n1454, u2_uk_n1456, u2_uk_n1457, u2_uk_n1458, u2_uk_n1459, u2_uk_n1460, u2_uk_n1461, u2_uk_n1462, u2_uk_n1464, 
       u2_uk_n1465, u2_uk_n1466, u2_uk_n1468, u2_uk_n147, u2_uk_n1470, u2_uk_n1471, u2_uk_n1475, u2_uk_n148, u2_uk_n1480, 
       u2_uk_n1486, u2_uk_n1487, u2_uk_n1488, u2_uk_n1490, u2_uk_n1491, u2_uk_n1493, u2_uk_n1494, u2_uk_n1496, u2_uk_n1497, 
       u2_uk_n1504, u2_uk_n1510, u2_uk_n1511, u2_uk_n1525, u2_uk_n1526, u2_uk_n1530, u2_uk_n1531, u2_uk_n1532, u2_uk_n1536, 
       u2_uk_n1537, u2_uk_n1538, u2_uk_n155, u2_uk_n1590, u2_uk_n1591, u2_uk_n1592, u2_uk_n1594, u2_uk_n1595, u2_uk_n1598, 
       u2_uk_n1600, u2_uk_n1603, u2_uk_n1604, u2_uk_n1605, u2_uk_n1609, u2_uk_n1610, u2_uk_n1612, u2_uk_n1614, u2_uk_n162, 
       u2_uk_n1623, u2_uk_n1624, u2_uk_n1626, u2_uk_n163, u2_uk_n1630, u2_uk_n1631, u2_uk_n1681, u2_uk_n1682, u2_uk_n1683, 
       u2_uk_n1688, u2_uk_n1689, u2_uk_n1693, u2_uk_n17, u2_uk_n1702, u2_uk_n1708, u2_uk_n1709, u2_uk_n1715, u2_uk_n1720, 
       u2_uk_n1721, u2_uk_n1722, u2_uk_n1769, u2_uk_n1770, u2_uk_n1781, u2_uk_n1785, u2_uk_n1792, u2_uk_n1797, u2_uk_n1803, 
       u2_uk_n1807, u2_uk_n1808, u2_uk_n1809, u2_uk_n1815, u2_uk_n1817, u2_uk_n1819, u2_uk_n1820, u2_uk_n1822, u2_uk_n1823, 
       u2_uk_n1825, u2_uk_n1826, u2_uk_n1833, u2_uk_n1834, u2_uk_n1835, u2_uk_n1838, u2_uk_n1839, u2_uk_n1840, u2_uk_n1843, 
       u2_uk_n1846, u2_uk_n1849, u2_uk_n1850, u2_uk_n1852, u2_uk_n1853, u2_uk_n1855, u2_uk_n188, u2_uk_n191, u2_uk_n203, 
       u2_uk_n207, u2_uk_n209, u2_uk_n214, u2_uk_n217, u2_uk_n223, u2_uk_n230, u2_uk_n231, u2_uk_n238, u2_uk_n240, 
       u2_uk_n251, u2_uk_n27, u2_uk_n408, u2_uk_n415, u2_uk_n421, u2_uk_n500, u2_uk_n520, u2_uk_n60, u2_uk_n63, 
       u2_uk_n689, u2_uk_n939, u2_uk_n941, u2_uk_n942, u2_uk_n943, u2_uk_n947, u2_uk_n954, u2_uk_n955, u2_uk_n956, 
       u2_uk_n961, u2_uk_n967, u2_uk_n970, u2_uk_n972, u2_uk_n99, u2_uk_n996, u2_uk_n997, u0_N0, u0_N1, u0_N12, u0_N128, u0_N129, u0_N133, u0_N137, u0_N140, u0_N143, 
        u0_N145, u0_N147, u0_N15, u0_N151, u0_N153, u0_N155, u0_N157, u0_N16, u0_N17, 
        u0_N19, u0_N22, u0_N23, u0_N25, u0_N27, u0_N29, u0_N30, u0_N416, u0_N417, 
        u0_N418, u0_N419, u0_N421, u0_N423, u0_N424, u0_N425, u0_N426, u0_N428, u0_N429, 
        u0_N431, u0_N432, u0_N433, u0_N434, u0_N435, u0_N438, u0_N439, u0_N440, u0_N441, 
        u0_N443, u0_N444, u0_N445, u0_N446, u0_N5, u0_N8, u0_N9, u0_uk_n674, u0_uk_n684, 
        u0_uk_n690, u0_uk_n696, u0_uk_n697, u0_uk_n698, u0_uk_n705, u0_uk_n871, u2_FP_11, u2_FP_12, u2_FP_14, 
        u2_FP_15, u2_FP_17, u2_FP_19, u2_FP_21, u2_FP_22, u2_FP_23, u2_FP_25, u2_FP_27, u2_FP_29, 
        u2_FP_3, u2_FP_31, u2_FP_32, u2_FP_4, u2_FP_5, u2_FP_7, u2_FP_8, u2_FP_9, u2_N0, 
        u2_N1, u2_N101, u2_N103, u2_N105, u2_N106, u2_N109, u2_N111, u2_N114, u2_N115, 
        u2_N119, u2_N12, u2_N120, u2_N121, u2_N124, u2_N125, u2_N128, u2_N129, u2_N133, 
        u2_N137, u2_N140, u2_N143, u2_N145, u2_N147, u2_N15, u2_N151, u2_N153, u2_N155, 
        u2_N157, u2_N16, u2_N160, u2_N162, u2_N167, u2_N169, u2_N17, u2_N173, u2_N179, 
        u2_N184, u2_N185, u2_N19, u2_N192, u2_N193, u2_N194, u2_N196, u2_N197, u2_N198, 
        u2_N199, u2_N200, u2_N201, u2_N203, u2_N204, u2_N205, u2_N206, u2_N207, u2_N208, 
        u2_N209, u2_N211, u2_N212, u2_N213, u2_N214, u2_N215, u2_N216, u2_N217, u2_N218, 
        u2_N219, u2_N22, u2_N221, u2_N222, u2_N223, u2_N228, u2_N23, u2_N230, u2_N235, 
        u2_N238, u2_N244, u2_N245, u2_N25, u2_N250, u2_N255, u2_N27, u2_N289, u2_N29, 
        u2_N292, u2_N293, u2_N296, u2_N30, u2_N300, u2_N302, u2_N303, u2_N304, u2_N305, 
        u2_N308, u2_N310, u2_N311, u2_N314, u2_N315, u2_N317, u2_N318, u2_N34, u2_N353, 
        u2_N357, u2_N360, u2_N364, u2_N367, u2_N368, u2_N369, u2_N374, u2_N375, u2_N379, 
        u2_N38, u2_N381, u2_N382, u2_N39, u2_N418, u2_N419, u2_N423, u2_N426, u2_N429, 
        u2_N43, u2_N434, u2_N440, u2_N444, u2_N449, u2_N45, u2_N450, u2_N451, u2_N454, 
        u2_N455, u2_N456, u2_N458, u2_N459, u2_N460, u2_N461, u2_N464, u2_N465, u2_N466, 
        u2_N469, u2_N470, u2_N472, u2_N475, u2_N476, u2_N478, u2_N479, u2_N5, u2_N53, 
        u2_N56, u2_N63, u2_N64, u2_N65, u2_N67, u2_N68, u2_N69, u2_N70, u2_N72, 
        u2_N73, u2_N74, u2_N75, u2_N76, u2_N78, u2_N79, u2_N8, u2_N80, u2_N81, 
        u2_N82, u2_N83, u2_N84, u2_N85, u2_N86, u2_N87, u2_N89, u2_N9, u2_N90, 
        u2_N91, u2_N92, u2_N93, u2_N94, u2_N95, u2_N96, u2_N98, u2_N99, u2_uk_n10, 
        u2_uk_n100, u2_uk_n1012, u2_uk_n1087, u2_uk_n1090, u2_uk_n11, u2_uk_n1102, u2_uk_n1145, u2_uk_n1146, u2_uk_n1155, 
        u2_uk_n1161, u2_uk_n1162, u2_uk_n1167, u2_uk_n1168, u2_uk_n117, u2_uk_n1179, u2_uk_n118, u2_uk_n129, u2_uk_n141, 
        u2_uk_n142, u2_uk_n146, u2_uk_n161, u2_uk_n164, u2_uk_n182, u2_uk_n187, u2_uk_n202, u2_uk_n208, u2_uk_n213, 
        u2_uk_n220, u2_uk_n222, u2_uk_n298, u2_uk_n31, u2_uk_n366, u2_uk_n656, u2_uk_n83, u2_uk_n92, u2_uk_n93, 
        u2_uk_n94, u2_uk_n983, u2_uk_n988 );
  input u0_K14_10, u0_K14_12, u0_K14_13, u0_K14_14, u0_K14_15, u0_K14_18, u0_K14_21, u0_K14_24, u0_K14_27, 
        u0_K14_4, u0_K14_9, u0_K1_13, u0_K1_14, u0_K1_15, u0_K1_16, u0_K1_17, u0_K1_23, u0_K5_13, 
        u0_K5_14, u0_K5_15, u0_K5_16, u0_K5_18, u0_K5_19, u0_K5_23, u0_K5_24, u0_K5_9, u0_L12_1, 
        u0_L12_10, u0_L12_11, u0_L12_13, u0_L12_14, u0_L12_16, u0_L12_17, u0_L12_18, u0_L12_19, u0_L12_2, 
        u0_L12_20, u0_L12_23, u0_L12_24, u0_L12_25, u0_L12_26, u0_L12_28, u0_L12_29, u0_L12_3, u0_L12_30, 
        u0_L12_31, u0_L12_4, u0_L12_6, u0_L12_8, u0_L12_9, u0_L3_1, u0_L3_10, u0_L3_13, u0_L3_16, 
        u0_L3_18, u0_L3_2, u0_L3_20, u0_L3_24, u0_L3_26, u0_L3_28, u0_L3_30, u0_L3_6, u0_R12_1, 
        u0_R12_10, u0_R12_11, u0_R12_12, u0_R12_13, u0_R12_14, u0_R12_15, u0_R12_16, u0_R12_17, u0_R12_18, 
        u0_R12_19, u0_R12_2, u0_R12_20, u0_R12_21, u0_R12_22, u0_R12_23, u0_R12_24, u0_R12_25, u0_R12_3, 
        u0_R12_32, u0_R12_4, u0_R12_5, u0_R12_6, u0_R12_7, u0_R12_8, u0_R12_9, u0_R3_10, u0_R3_11, 
        u0_R3_12, u0_R3_13, u0_R3_14, u0_R3_15, u0_R3_16, u0_R3_17, u0_R3_4, u0_R3_5, u0_R3_6, 
        u0_R3_7, u0_R3_8, u0_R3_9, u0_desIn_r_10, u0_desIn_r_12, u0_desIn_r_13, u0_desIn_r_14, u0_desIn_r_15, u0_desIn_r_2, 
        u0_desIn_r_21, u0_desIn_r_23, u0_desIn_r_24, u0_desIn_r_26, u0_desIn_r_29, u0_desIn_r_3, u0_desIn_r_31, u0_desIn_r_36, u0_desIn_r_37, 
        u0_desIn_r_39, u0_desIn_r_4, u0_desIn_r_40, u0_desIn_r_45, u0_desIn_r_46, u0_desIn_r_47, u0_desIn_r_48, u0_desIn_r_5, u0_desIn_r_50, 
        u0_desIn_r_53, u0_desIn_r_55, u0_desIn_r_57, u0_desIn_r_58, u0_desIn_r_6, u0_desIn_r_60, u0_desIn_r_61, u0_desIn_r_63, u0_desIn_r_7, 
        u0_desIn_r_8, u0_key_r_11, u0_key_r_12, u0_key_r_13, u0_key_r_17, u0_key_r_19, u0_key_r_20, u0_key_r_24, u0_key_r_25, 
        u0_key_r_26, u0_key_r_27, u0_key_r_3, u0_key_r_32, u0_key_r_34, u0_key_r_39, u0_key_r_4, u0_key_r_40, u0_key_r_41, 
        u0_key_r_47, u0_key_r_48, u0_key_r_49, u0_key_r_5, u0_key_r_53, u0_key_r_54, u0_key_r_55, u0_key_r_6, u0_uk_K_r12_1, 
        u0_uk_K_r12_10, u0_uk_K_r12_25, u0_uk_K_r12_30, u0_uk_K_r12_33, u0_uk_K_r12_36, u0_uk_K_r12_44, u0_uk_K_r12_47, u0_uk_K_r12_7, u0_uk_K_r3_11, 
        u0_uk_K_r3_19, u0_uk_K_r3_24, u0_uk_K_r3_47, u0_uk_n10, u0_uk_n100, u0_uk_n109, u0_uk_n11, u0_uk_n110, u0_uk_n117, 
        u0_uk_n118, u0_uk_n128, u0_uk_n129, u0_uk_n141, u0_uk_n142, u0_uk_n145, u0_uk_n146, u0_uk_n147, u0_uk_n163, 
        u0_uk_n164, u0_uk_n17, u0_uk_n182, u0_uk_n187, u0_uk_n188, u0_uk_n202, u0_uk_n203, u0_uk_n207, u0_uk_n208, 
        u0_uk_n213, u0_uk_n217, u0_uk_n220, u0_uk_n222, u0_uk_n230, u0_uk_n231, u0_uk_n240, u0_uk_n242, u0_uk_n250, 
        u0_uk_n251, u0_uk_n257, u0_uk_n451, u0_uk_n453, u0_uk_n459, u0_uk_n46, u0_uk_n464, u0_uk_n465, u0_uk_n473, 
        u0_uk_n479, u0_uk_n48, u0_uk_n483, u0_uk_n484, u0_uk_n485, u0_uk_n489, u0_uk_n49, u0_uk_n50, u0_uk_n51, 
        u0_uk_n53, u0_uk_n54, u0_uk_n55, u0_uk_n57, u0_uk_n61, u0_uk_n62, u0_uk_n63, u0_uk_n64, u0_uk_n66, 
        u0_uk_n67, u0_uk_n69, u0_uk_n72, u0_uk_n73, u0_uk_n75, u0_uk_n77, u0_uk_n78, u0_uk_n79, u0_uk_n80, 
        u0_uk_n815, u0_uk_n82, u0_uk_n83, u0_uk_n84, u0_uk_n85, u0_uk_n86, u0_uk_n87, u0_uk_n88, u0_uk_n89, 
        u0_uk_n92, u0_uk_n93, u0_uk_n94, u0_uk_n99, u2_FP_33, u2_FP_34, u2_FP_35, u2_FP_36, u2_FP_37, 
        u2_FP_48, u2_FP_49, u2_FP_50, u2_FP_51, u2_FP_52, u2_FP_53, u2_FP_54, u2_FP_55, u2_FP_56, 
        u2_FP_57, u2_FP_58, u2_FP_59, u2_FP_60, u2_FP_61, u2_FP_62, u2_FP_63, u2_FP_64, u2_K10_10, 
        u2_K10_11, u2_K10_15, u2_K10_17, u2_K10_4, u2_K10_43, u2_K10_44, u2_K10_46, u2_K10_6, u2_K12_2, 
        u2_K12_8, u2_K14_25, u2_K14_28, u2_K15_1, u2_K15_2, u2_K15_28, u2_K15_29, u2_K15_31, u2_K15_34, 
        u2_K15_35, u2_K15_39, u2_K15_5, u2_K16_26, u2_K16_31, u2_K16_42, u2_K16_44, u2_K16_47, u2_K16_5, 
        u2_K16_6, u2_K1_15, u2_K1_16, u2_K1_19, u2_K1_24, u2_K1_5, u2_K1_9, u2_K2_40, u2_K3_13, 
        u2_K3_15, u2_K3_16, u2_K3_20, u2_K3_23, u2_K3_32, u2_K3_35, u2_K3_42, u2_K3_43, u2_K3_47, 
        u2_K3_48, u2_K3_7, u2_K4_14, u2_K4_21, u2_K4_22, u2_K4_27, u2_K4_33, u2_K4_34, u2_K4_35, 
        u2_K5_10, u2_K5_11, u2_K5_13, u2_K5_14, u2_K5_16, u2_K5_17, u2_K5_18, u2_K5_19, u2_K5_21, 
        u2_K5_23, u2_K5_24, u2_K5_8, u2_K5_9, u2_K6_20, u2_K6_22, u2_K6_24, u2_K6_25, u2_K6_27, 
        u2_K7_26, u2_K7_3, u2_K7_37, u2_K7_38, u2_K7_4, u2_K7_43, u2_K7_45, u2_K7_48, u2_K7_5, 
        u2_K7_7, u2_K8_41, u2_K8_45, u2_L0_12, u2_L0_14, u2_L0_22, u2_L0_25, u2_L0_3, u2_L0_32, 
        u2_L0_7, u2_L0_8, u2_L10_13, u2_L10_16, u2_L10_17, u2_L10_18, u2_L10_2, u2_L10_23, u2_L10_24, 
        u2_L10_28, u2_L10_30, u2_L10_31, u2_L10_6, u2_L10_9, u2_L12_11, u2_L12_14, u2_L12_19, u2_L12_25, 
        u2_L12_29, u2_L12_3, u2_L12_4, u2_L12_8, u2_L13_11, u2_L13_12, u2_L13_13, u2_L13_14, u2_L13_17, 
        u2_L13_18, u2_L13_19, u2_L13_2, u2_L13_22, u2_L13_23, u2_L13_25, u2_L13_28, u2_L13_29, u2_L13_3, 
        u2_L13_31, u2_L13_32, u2_L13_4, u2_L13_7, u2_L13_8, u2_L13_9, u2_L14_11, u2_L14_12, u2_L14_14, 
        u2_L14_15, u2_L14_17, u2_L14_19, u2_L14_21, u2_L14_22, u2_L14_23, u2_L14_25, u2_L14_27, u2_L14_29, 
        u2_L14_3, u2_L14_31, u2_L14_32, u2_L14_4, u2_L14_5, u2_L14_7, u2_L14_8, u2_L14_9, u2_L1_1, 
        u2_L1_10, u2_L1_11, u2_L1_12, u2_L1_13, u2_L1_15, u2_L1_16, u2_L1_17, u2_L1_18, u2_L1_19, 
        u2_L1_2, u2_L1_20, u2_L1_21, u2_L1_22, u2_L1_23, u2_L1_24, u2_L1_26, u2_L1_27, u2_L1_28, 
        u2_L1_29, u2_L1_30, u2_L1_31, u2_L1_32, u2_L1_4, u2_L1_5, u2_L1_6, u2_L1_7, u2_L1_9, 
        u2_L2_1, u2_L2_10, u2_L2_11, u2_L2_14, u2_L2_16, u2_L2_19, u2_L2_20, u2_L2_24, u2_L2_25, 
        u2_L2_26, u2_L2_29, u2_L2_3, u2_L2_30, u2_L2_4, u2_L2_6, u2_L2_8, u2_L3_1, u2_L3_10, 
        u2_L3_13, u2_L3_16, u2_L3_18, u2_L3_2, u2_L3_20, u2_L3_24, u2_L3_26, u2_L3_28, u2_L3_30, 
        u2_L3_6, u2_L4_1, u2_L4_10, u2_L4_14, u2_L4_20, u2_L4_25, u2_L4_26, u2_L4_3, u2_L4_8, 
        u2_L5_1, u2_L5_10, u2_L5_12, u2_L5_13, u2_L5_14, u2_L5_15, u2_L5_16, u2_L5_17, u2_L5_18, 
        u2_L5_2, u2_L5_20, u2_L5_21, u2_L5_22, u2_L5_23, u2_L5_24, u2_L5_25, u2_L5_26, u2_L5_27, 
        u2_L5_28, u2_L5_3, u2_L5_30, u2_L5_31, u2_L5_32, u2_L5_5, u2_L5_6, u2_L5_7, u2_L5_8, 
        u2_L5_9, u2_L6_12, u2_L6_15, u2_L6_21, u2_L6_22, u2_L6_27, u2_L6_32, u2_L6_5, u2_L6_7, 
        u2_L8_13, u2_L8_15, u2_L8_16, u2_L8_17, u2_L8_18, u2_L8_2, u2_L8_21, u2_L8_23, u2_L8_24, 
        u2_L8_27, u2_L8_28, u2_L8_30, u2_L8_31, u2_L8_5, u2_L8_6, u2_L8_9, u2_R0_16, u2_R0_17, 
        u2_R0_18, u2_R0_19, u2_R0_20, u2_R0_21, u2_R0_24, u2_R0_25, u2_R0_26, u2_R0_27, u2_R0_28, 
        u2_R0_29, u2_R10_1, u2_R10_10, u2_R10_11, u2_R10_12, u2_R10_13, u2_R10_2, u2_R10_3, u2_R10_32, 
        u2_R10_4, u2_R10_5, u2_R10_6, u2_R10_7, u2_R10_8, u2_R10_9, u2_R12_16, u2_R12_17, u2_R12_18, 
        u2_R12_19, u2_R12_20, u2_R12_21, u2_R12_22, u2_R12_23, u2_R12_24, u2_R12_25, u2_R13_1, u2_R13_16, 
        u2_R13_17, u2_R13_18, u2_R13_19, u2_R13_2, u2_R13_20, u2_R13_21, u2_R13_22, u2_R13_23, u2_R13_24, 
        u2_R13_25, u2_R13_26, u2_R13_27, u2_R13_28, u2_R13_29, u2_R13_3, u2_R13_32, u2_R13_4, u2_R13_5, 
        u2_R13_6, u2_R13_7, u2_R13_8, u2_R13_9, u2_R1_1, u2_R1_10, u2_R1_11, u2_R1_12, u2_R1_13, 
        u2_R1_14, u2_R1_15, u2_R1_16, u2_R1_17, u2_R1_2, u2_R1_20, u2_R1_21, u2_R1_22, u2_R1_23, 
        u2_R1_24, u2_R1_25, u2_R1_26, u2_R1_27, u2_R1_28, u2_R1_29, u2_R1_3, u2_R1_30, u2_R1_31, 
        u2_R1_32, u2_R1_4, u2_R1_5, u2_R1_6, u2_R1_7, u2_R1_8, u2_R1_9, u2_R2_10, u2_R2_11, 
        u2_R2_12, u2_R2_13, u2_R2_14, u2_R2_15, u2_R2_16, u2_R2_17, u2_R2_18, u2_R2_19, u2_R2_20, 
        u2_R2_21, u2_R2_22, u2_R2_23, u2_R2_24, u2_R2_25, u2_R2_8, u2_R2_9, u2_R3_10, u2_R3_11, 
        u2_R3_12, u2_R3_13, u2_R3_14, u2_R3_15, u2_R3_16, u2_R3_17, u2_R3_4, u2_R3_5, u2_R3_6, 
        u2_R3_7, u2_R3_8, u2_R3_9, u2_R4_12, u2_R4_13, u2_R4_14, u2_R4_15, u2_R4_16, u2_R4_17, 
        u2_R4_18, u2_R4_19, u2_R4_20, u2_R4_21, u2_R5_1, u2_R5_10, u2_R5_11, u2_R5_12, u2_R5_13, 
        u2_R5_14, u2_R5_15, u2_R5_16, u2_R5_17, u2_R5_18, u2_R5_19, u2_R5_2, u2_R5_20, u2_R5_21, 
        u2_R5_24, u2_R5_25, u2_R5_26, u2_R5_27, u2_R5_28, u2_R5_29, u2_R5_3, u2_R5_30, u2_R5_31, 
        u2_R5_32, u2_R5_4, u2_R5_5, u2_R5_6, u2_R5_7, u2_R5_8, u2_R5_9, u2_R6_1, u2_R6_24, 
        u2_R6_25, u2_R6_26, u2_R6_27, u2_R6_28, u2_R6_29, u2_R6_30, u2_R6_31, u2_R6_32, u2_R8_1, 
        u2_R8_10, u2_R8_11, u2_R8_12, u2_R8_13, u2_R8_2, u2_R8_28, u2_R8_29, u2_R8_3, u2_R8_30, 
        u2_R8_31, u2_R8_32, u2_R8_4, u2_R8_5, u2_R8_6, u2_R8_7, u2_R8_8, u2_R8_9, u2_desIn_r_10, 
        u2_desIn_r_12, u2_desIn_r_13, u2_desIn_r_14, u2_desIn_r_15, u2_desIn_r_2, u2_desIn_r_21, u2_desIn_r_23, u2_desIn_r_24, u2_desIn_r_26, 
        u2_desIn_r_29, u2_desIn_r_3, u2_desIn_r_31, u2_desIn_r_36, u2_desIn_r_37, u2_desIn_r_39, u2_desIn_r_4, u2_desIn_r_40, u2_desIn_r_45, 
        u2_desIn_r_46, u2_desIn_r_47, u2_desIn_r_48, u2_desIn_r_5, u2_desIn_r_50, u2_desIn_r_53, u2_desIn_r_55, u2_desIn_r_57, u2_desIn_r_58, 
        u2_desIn_r_6, u2_desIn_r_60, u2_desIn_r_61, u2_desIn_r_63, u2_desIn_r_7, u2_desIn_r_8, u2_key_r_10, u2_key_r_11, u2_key_r_12, 
        u2_key_r_17, u2_key_r_19, u2_key_r_20, u2_key_r_24, u2_key_r_25, u2_key_r_26, u2_key_r_27, u2_key_r_3, u2_key_r_32, 
        u2_key_r_33, u2_key_r_34, u2_key_r_4, u2_key_r_40, u2_key_r_41, u2_key_r_46, u2_key_r_47, u2_key_r_48, u2_key_r_49, 
        u2_key_r_50, u2_key_r_53, u2_key_r_55, u2_key_r_6, u2_uk_K_r0_15, u2_uk_K_r0_49, u2_uk_K_r10_10, u2_uk_K_r10_25, u2_uk_K_r10_27, 
        u2_uk_K_r10_34, u2_uk_K_r10_4, u2_uk_K_r11_7, u2_uk_K_r12_1, u2_uk_K_r12_30, u2_uk_K_r12_36, u2_uk_K_r12_42, u2_uk_K_r12_7, u2_uk_K_r13_0, 
        u2_uk_K_r13_13, u2_uk_K_r13_17, u2_uk_K_r13_22, u2_uk_K_r13_25, u2_uk_K_r13_38, u2_uk_K_r13_55, u2_uk_K_r14_15, u2_uk_K_r14_16, u2_uk_K_r14_2, 
        u2_uk_K_r14_3, u2_uk_K_r14_45, u2_uk_K_r14_50, u2_uk_K_r14_9, u2_uk_K_r1_15, u2_uk_K_r1_16, u2_uk_K_r1_17, u2_uk_K_r1_18, u2_uk_K_r1_21, 
        u2_uk_K_r1_22, u2_uk_K_r1_41, u2_uk_K_r1_47, u2_uk_K_r1_7, u2_uk_K_r2_18, u2_uk_K_r2_21, u2_uk_K_r2_27, u2_uk_K_r2_28, u2_uk_K_r2_31, 
        u2_uk_K_r2_36, u2_uk_K_r2_49, u2_uk_K_r2_55, u2_uk_K_r3_11, u2_uk_K_r3_19, u2_uk_K_r4_0, u2_uk_K_r4_11, u2_uk_K_r4_35, u2_uk_K_r4_5, 
        u2_uk_K_r5_10, u2_uk_K_r5_16, u2_uk_K_r5_17, u2_uk_K_r5_18, u2_uk_K_r5_19, u2_uk_K_r5_23, u2_uk_K_r5_26, u2_uk_K_r5_31, u2_uk_K_r5_37, 
        u2_uk_K_r5_39, u2_uk_K_r5_4, u2_uk_K_r5_40, u2_uk_K_r5_41, u2_uk_K_r5_43, u2_uk_K_r5_48, u2_uk_K_r5_7, u2_uk_K_r6_0, u2_uk_K_r6_14, 
        u2_uk_K_r6_31, u2_uk_K_r6_37, u2_uk_K_r6_46, u2_uk_K_r6_7, u2_uk_K_r8_17, u2_uk_K_r8_21, u2_uk_K_r8_27, u2_uk_K_r8_32, u2_uk_K_r8_41, 
        u2_uk_K_r8_48, u2_uk_K_r9_0, u2_uk_n1001, u2_uk_n1007, u2_uk_n1011, u2_uk_n1018, u2_uk_n102, u2_uk_n1022, u2_uk_n1024, 
        u2_uk_n1027, u2_uk_n1028, u2_uk_n1042, u2_uk_n1043, u2_uk_n1044, u2_uk_n1061, u2_uk_n1063, u2_uk_n1077, u2_uk_n1079, 
        u2_uk_n1081, u2_uk_n1082, u2_uk_n109, u2_uk_n1093, u2_uk_n1094, u2_uk_n1096, u2_uk_n110, u2_uk_n1112, u2_uk_n1113, 
        u2_uk_n1188, u2_uk_n1189, u2_uk_n1190, u2_uk_n1195, u2_uk_n1198, u2_uk_n1200, u2_uk_n1201, u2_uk_n1203, u2_uk_n1206, 
        u2_uk_n1208, u2_uk_n1209, u2_uk_n1210, u2_uk_n1215, u2_uk_n1216, u2_uk_n1217, u2_uk_n1218, u2_uk_n1220, u2_uk_n1221, 
        u2_uk_n1223, u2_uk_n1225, u2_uk_n1226, u2_uk_n1227, u2_uk_n1230, u2_uk_n1236, u2_uk_n1237, u2_uk_n1246, u2_uk_n1251, 
        u2_uk_n1252, u2_uk_n1259, u2_uk_n1264, u2_uk_n1265, u2_uk_n1266, u2_uk_n1274, u2_uk_n1279, u2_uk_n128, u2_uk_n1280, 
        u2_uk_n1281, u2_uk_n1282, u2_uk_n1283, u2_uk_n1284, u2_uk_n1285, u2_uk_n1286, u2_uk_n1287, u2_uk_n1288, u2_uk_n1290, 
        u2_uk_n1291, u2_uk_n1292, u2_uk_n1293, u2_uk_n1294, u2_uk_n1295, u2_uk_n1296, u2_uk_n1297, u2_uk_n1298, u2_uk_n1299, 
        u2_uk_n1300, u2_uk_n1301, u2_uk_n1302, u2_uk_n1303, u2_uk_n1305, u2_uk_n1306, u2_uk_n1308, u2_uk_n1309, u2_uk_n1310, 
        u2_uk_n1311, u2_uk_n1312, u2_uk_n1314, u2_uk_n1316, u2_uk_n1317, u2_uk_n1318, u2_uk_n1322, u2_uk_n1324, u2_uk_n1326, 
        u2_uk_n1328, u2_uk_n1329, u2_uk_n1333, u2_uk_n1335, u2_uk_n1339, u2_uk_n1345, u2_uk_n1346, u2_uk_n1347, u2_uk_n1348, 
        u2_uk_n1350, u2_uk_n1351, u2_uk_n1356, u2_uk_n1363, u2_uk_n1375, u2_uk_n1379, u2_uk_n1405, u2_uk_n1408, u2_uk_n1412, 
        u2_uk_n1413, u2_uk_n1414, u2_uk_n1420, u2_uk_n1439, u2_uk_n1442, u2_uk_n1447, u2_uk_n145, u2_uk_n1452, u2_uk_n1453, 
        u2_uk_n1454, u2_uk_n1456, u2_uk_n1457, u2_uk_n1458, u2_uk_n1459, u2_uk_n1460, u2_uk_n1461, u2_uk_n1462, u2_uk_n1464, 
        u2_uk_n1465, u2_uk_n1466, u2_uk_n1468, u2_uk_n147, u2_uk_n1470, u2_uk_n1471, u2_uk_n1475, u2_uk_n148, u2_uk_n1480, 
        u2_uk_n1486, u2_uk_n1487, u2_uk_n1488, u2_uk_n1490, u2_uk_n1491, u2_uk_n1493, u2_uk_n1494, u2_uk_n1496, u2_uk_n1497, 
        u2_uk_n1504, u2_uk_n1510, u2_uk_n1511, u2_uk_n1525, u2_uk_n1526, u2_uk_n1530, u2_uk_n1531, u2_uk_n1532, u2_uk_n1536, 
        u2_uk_n1537, u2_uk_n1538, u2_uk_n155, u2_uk_n1590, u2_uk_n1591, u2_uk_n1592, u2_uk_n1594, u2_uk_n1595, u2_uk_n1598, 
        u2_uk_n1600, u2_uk_n1603, u2_uk_n1604, u2_uk_n1605, u2_uk_n1609, u2_uk_n1610, u2_uk_n1612, u2_uk_n1614, u2_uk_n162, 
        u2_uk_n1623, u2_uk_n1624, u2_uk_n1626, u2_uk_n163, u2_uk_n1630, u2_uk_n1631, u2_uk_n1681, u2_uk_n1682, u2_uk_n1683, 
        u2_uk_n1688, u2_uk_n1689, u2_uk_n1693, u2_uk_n17, u2_uk_n1702, u2_uk_n1708, u2_uk_n1709, u2_uk_n1715, u2_uk_n1720, 
        u2_uk_n1721, u2_uk_n1722, u2_uk_n1769, u2_uk_n1770, u2_uk_n1781, u2_uk_n1785, u2_uk_n1792, u2_uk_n1797, u2_uk_n1803, 
        u2_uk_n1807, u2_uk_n1808, u2_uk_n1809, u2_uk_n1815, u2_uk_n1817, u2_uk_n1819, u2_uk_n1820, u2_uk_n1822, u2_uk_n1823, 
        u2_uk_n1825, u2_uk_n1826, u2_uk_n1833, u2_uk_n1834, u2_uk_n1835, u2_uk_n1838, u2_uk_n1839, u2_uk_n1840, u2_uk_n1843, 
        u2_uk_n1846, u2_uk_n1849, u2_uk_n1850, u2_uk_n1852, u2_uk_n1853, u2_uk_n1855, u2_uk_n188, u2_uk_n191, u2_uk_n203, 
        u2_uk_n207, u2_uk_n209, u2_uk_n214, u2_uk_n217, u2_uk_n223, u2_uk_n230, u2_uk_n231, u2_uk_n238, u2_uk_n240, 
        u2_uk_n251, u2_uk_n27, u2_uk_n408, u2_uk_n415, u2_uk_n421, u2_uk_n500, u2_uk_n520, u2_uk_n60, u2_uk_n63, 
        u2_uk_n689, u2_uk_n939, u2_uk_n941, u2_uk_n942, u2_uk_n943, u2_uk_n947, u2_uk_n954, u2_uk_n955, u2_uk_n956, 
        u2_uk_n961, u2_uk_n967, u2_uk_n970, u2_uk_n972, u2_uk_n99, u2_uk_n996, u2_uk_n997;
  output u0_N0, u0_N1, u0_N12, u0_N128, u0_N129, u0_N133, u0_N137, u0_N140, u0_N143, 
        u0_N145, u0_N147, u0_N15, u0_N151, u0_N153, u0_N155, u0_N157, u0_N16, u0_N17, 
        u0_N19, u0_N22, u0_N23, u0_N25, u0_N27, u0_N29, u0_N30, u0_N416, u0_N417, 
        u0_N418, u0_N419, u0_N421, u0_N423, u0_N424, u0_N425, u0_N426, u0_N428, u0_N429, 
        u0_N431, u0_N432, u0_N433, u0_N434, u0_N435, u0_N438, u0_N439, u0_N440, u0_N441, 
        u0_N443, u0_N444, u0_N445, u0_N446, u0_N5, u0_N8, u0_N9, u0_uk_n674, u0_uk_n684, 
        u0_uk_n690, u0_uk_n696, u0_uk_n697, u0_uk_n698, u0_uk_n705, u0_uk_n871, u2_FP_11, u2_FP_12, u2_FP_14, 
        u2_FP_15, u2_FP_17, u2_FP_19, u2_FP_21, u2_FP_22, u2_FP_23, u2_FP_25, u2_FP_27, u2_FP_29, 
        u2_FP_3, u2_FP_31, u2_FP_32, u2_FP_4, u2_FP_5, u2_FP_7, u2_FP_8, u2_FP_9, u2_N0, 
        u2_N1, u2_N101, u2_N103, u2_N105, u2_N106, u2_N109, u2_N111, u2_N114, u2_N115, 
        u2_N119, u2_N12, u2_N120, u2_N121, u2_N124, u2_N125, u2_N128, u2_N129, u2_N133, 
        u2_N137, u2_N140, u2_N143, u2_N145, u2_N147, u2_N15, u2_N151, u2_N153, u2_N155, 
        u2_N157, u2_N16, u2_N160, u2_N162, u2_N167, u2_N169, u2_N17, u2_N173, u2_N179, 
        u2_N184, u2_N185, u2_N19, u2_N192, u2_N193, u2_N194, u2_N196, u2_N197, u2_N198, 
        u2_N199, u2_N200, u2_N201, u2_N203, u2_N204, u2_N205, u2_N206, u2_N207, u2_N208, 
        u2_N209, u2_N211, u2_N212, u2_N213, u2_N214, u2_N215, u2_N216, u2_N217, u2_N218, 
        u2_N219, u2_N22, u2_N221, u2_N222, u2_N223, u2_N228, u2_N23, u2_N230, u2_N235, 
        u2_N238, u2_N244, u2_N245, u2_N25, u2_N250, u2_N255, u2_N27, u2_N289, u2_N29, 
        u2_N292, u2_N293, u2_N296, u2_N30, u2_N300, u2_N302, u2_N303, u2_N304, u2_N305, 
        u2_N308, u2_N310, u2_N311, u2_N314, u2_N315, u2_N317, u2_N318, u2_N34, u2_N353, 
        u2_N357, u2_N360, u2_N364, u2_N367, u2_N368, u2_N369, u2_N374, u2_N375, u2_N379, 
        u2_N38, u2_N381, u2_N382, u2_N39, u2_N418, u2_N419, u2_N423, u2_N426, u2_N429, 
        u2_N43, u2_N434, u2_N440, u2_N444, u2_N449, u2_N45, u2_N450, u2_N451, u2_N454, 
        u2_N455, u2_N456, u2_N458, u2_N459, u2_N460, u2_N461, u2_N464, u2_N465, u2_N466, 
        u2_N469, u2_N470, u2_N472, u2_N475, u2_N476, u2_N478, u2_N479, u2_N5, u2_N53, 
        u2_N56, u2_N63, u2_N64, u2_N65, u2_N67, u2_N68, u2_N69, u2_N70, u2_N72, 
        u2_N73, u2_N74, u2_N75, u2_N76, u2_N78, u2_N79, u2_N8, u2_N80, u2_N81, 
        u2_N82, u2_N83, u2_N84, u2_N85, u2_N86, u2_N87, u2_N89, u2_N9, u2_N90, 
        u2_N91, u2_N92, u2_N93, u2_N94, u2_N95, u2_N96, u2_N98, u2_N99, u2_uk_n10, 
        u2_uk_n100, u2_uk_n1012, u2_uk_n1087, u2_uk_n1090, u2_uk_n11, u2_uk_n1102, u2_uk_n1145, u2_uk_n1146, u2_uk_n1155, 
        u2_uk_n1161, u2_uk_n1162, u2_uk_n1167, u2_uk_n1168, u2_uk_n117, u2_uk_n1179, u2_uk_n118, u2_uk_n129, u2_uk_n141, 
        u2_uk_n142, u2_uk_n146, u2_uk_n161, u2_uk_n164, u2_uk_n182, u2_uk_n187, u2_uk_n202, u2_uk_n208, u2_uk_n213, 
        u2_uk_n220, u2_uk_n222, u2_uk_n298, u2_uk_n31, u2_uk_n366, u2_uk_n656, u2_uk_n83, u2_uk_n92, u2_uk_n93, 
        u2_uk_n94, u2_uk_n983, u2_uk_n988;
  wire u0_K14_1, u0_K14_11, u0_K14_16, u0_K14_17, u0_K14_19, u0_K14_2, u0_K14_20, u0_K14_22, u0_K14_23, 
       u0_K14_25, u0_K14_26, u0_K14_28, u0_K14_29, u0_K14_3, u0_K14_30, u0_K14_31, u0_K14_32, u0_K14_33, 
       u0_K14_34, u0_K14_35, u0_K14_36, u0_K14_5, u0_K14_6, u0_K14_7, u0_K14_8, u0_K1_1, u0_K1_10, 
       u0_K1_11, u0_K1_12, u0_K1_18, u0_K1_19, u0_K1_2, u0_K1_20, u0_K1_21, u0_K1_22, u0_K1_24, 
       u0_K1_3, u0_K1_4, u0_K1_5, u0_K1_6, u0_K1_7, u0_K1_8, u0_K1_9, u0_K5_10, u0_K5_11, 
       u0_K5_12, u0_K5_17, u0_K5_20, u0_K5_21, u0_K5_22, u0_K5_7, u0_K5_8, u0_out0_1, u0_out0_10, 
       u0_out0_13, u0_out0_16, u0_out0_17, u0_out0_18, u0_out0_2, u0_out0_20, u0_out0_23, u0_out0_24, u0_out0_26, 
       u0_out0_28, u0_out0_30, u0_out0_31, u0_out0_6, u0_out0_9, u0_out13_1, u0_out13_10, u0_out13_11, u0_out13_13, 
       u0_out13_14, u0_out13_16, u0_out13_17, u0_out13_18, u0_out13_19, u0_out13_2, u0_out13_20, u0_out13_23, u0_out13_24, 
       u0_out13_25, u0_out13_26, u0_out13_28, u0_out13_29, u0_out13_3, u0_out13_30, u0_out13_31, u0_out13_4, u0_out13_6, 
       u0_out13_8, u0_out13_9, u0_out4_1, u0_out4_10, u0_out4_13, u0_out4_16, u0_out4_18, u0_out4_2, u0_out4_20, 
       u0_out4_24, u0_out4_26, u0_out4_28, u0_out4_30, u0_out4_6, u0_u0_X_1, u0_u0_X_10, u0_u0_X_11, u0_u0_X_12, 
       u0_u0_X_13, u0_u0_X_14, u0_u0_X_15, u0_u0_X_16, u0_u0_X_17, u0_u0_X_18, u0_u0_X_19, u0_u0_X_2, u0_u0_X_20, 
       u0_u0_X_21, u0_u0_X_22, u0_u0_X_23, u0_u0_X_24, u0_u0_X_3, u0_u0_X_4, u0_u0_X_5, u0_u0_X_6, u0_u0_X_7, 
       u0_u0_X_8, u0_u0_X_9, u0_u0_u0_n1, u0_u0_u0_n10, u0_u0_u0_n11, u0_u0_u0_n12, u0_u0_u0_n13, u0_u0_u0_n14, u0_u0_u0_n15, 
       u0_u0_u0_n16, u0_u0_u0_n17, u0_u0_u0_n18, u0_u0_u0_n19, u0_u0_u0_n2, u0_u0_u0_n20, u0_u0_u0_n21, u0_u0_u0_n22, u0_u0_u0_n23, 
       u0_u0_u0_n24, u0_u0_u0_n25, u0_u0_u0_n26, u0_u0_u0_n27, u0_u0_u0_n28, u0_u0_u0_n29, u0_u0_u0_n3, u0_u0_u0_n30, u0_u0_u0_n31, 
       u0_u0_u0_n32, u0_u0_u0_n33, u0_u0_u0_n34, u0_u0_u0_n35, u0_u0_u0_n36, u0_u0_u0_n37, u0_u0_u0_n38, u0_u0_u0_n39, u0_u0_u0_n4, 
       u0_u0_u0_n40, u0_u0_u0_n41, u0_u0_u0_n42, u0_u0_u0_n43, u0_u0_u0_n44, u0_u0_u0_n45, u0_u0_u0_n46, u0_u0_u0_n47, u0_u0_u0_n48, 
       u0_u0_u0_n49, u0_u0_u0_n5, u0_u0_u0_n50, u0_u0_u0_n51, u0_u0_u0_n52, u0_u0_u0_n53, u0_u0_u0_n54, u0_u0_u0_n55, u0_u0_u0_n56, 
       u0_u0_u0_n57, u0_u0_u0_n58, u0_u0_u0_n59, u0_u0_u0_n6, u0_u0_u0_n60, u0_u0_u0_n61, u0_u0_u0_n62, u0_u0_u0_n63, u0_u0_u0_n64, 
       u0_u0_u0_n65, u0_u0_u0_n66, u0_u0_u0_n67, u0_u0_u0_n68, u0_u0_u0_n69, u0_u0_u0_n7, u0_u0_u0_n70, u0_u0_u0_n71, u0_u0_u0_n72, 
       u0_u0_u0_n73, u0_u0_u0_n74, u0_u0_u0_n75, u0_u0_u0_n76, u0_u0_u0_n77, u0_u0_u0_n78, u0_u0_u0_n79, u0_u0_u0_n8, u0_u0_u0_n80, 
       u0_u0_u0_n81, u0_u0_u0_n82, u0_u0_u0_n83, u0_u0_u0_n84, u0_u0_u0_n85, u0_u0_u0_n86, u0_u0_u0_n87, u0_u0_u0_n9, u0_u0_u1_n1, 
       u0_u0_u1_n10, u0_u0_u1_n11, u0_u0_u1_n12, u0_u0_u1_n13, u0_u0_u1_n14, u0_u0_u1_n15, u0_u0_u1_n16, u0_u0_u1_n17, u0_u0_u1_n18, 
       u0_u0_u1_n19, u0_u0_u1_n2, u0_u0_u1_n20, u0_u0_u1_n21, u0_u0_u1_n22, u0_u0_u1_n23, u0_u0_u1_n24, u0_u0_u1_n25, u0_u0_u1_n26, 
       u0_u0_u1_n27, u0_u0_u1_n28, u0_u0_u1_n29, u0_u0_u1_n3, u0_u0_u1_n30, u0_u0_u1_n31, u0_u0_u1_n32, u0_u0_u1_n33, u0_u0_u1_n34, 
       u0_u0_u1_n35, u0_u0_u1_n36, u0_u0_u1_n37, u0_u0_u1_n38, u0_u0_u1_n39, u0_u0_u1_n4, u0_u0_u1_n40, u0_u0_u1_n41, u0_u0_u1_n42, 
       u0_u0_u1_n43, u0_u0_u1_n44, u0_u0_u1_n45, u0_u0_u1_n46, u0_u0_u1_n47, u0_u0_u1_n48, u0_u0_u1_n49, u0_u0_u1_n5, u0_u0_u1_n50, 
       u0_u0_u1_n51, u0_u0_u1_n52, u0_u0_u1_n53, u0_u0_u1_n54, u0_u0_u1_n55, u0_u0_u1_n56, u0_u0_u1_n57, u0_u0_u1_n58, u0_u0_u1_n59, 
       u0_u0_u1_n6, u0_u0_u1_n60, u0_u0_u1_n61, u0_u0_u1_n62, u0_u0_u1_n63, u0_u0_u1_n64, u0_u0_u1_n65, u0_u0_u1_n66, u0_u0_u1_n67, 
       u0_u0_u1_n68, u0_u0_u1_n69, u0_u0_u1_n7, u0_u0_u1_n70, u0_u0_u1_n71, u0_u0_u1_n72, u0_u0_u1_n73, u0_u0_u1_n74, u0_u0_u1_n75, 
       u0_u0_u1_n76, u0_u0_u1_n77, u0_u0_u1_n78, u0_u0_u1_n79, u0_u0_u1_n8, u0_u0_u1_n80, u0_u0_u1_n81, u0_u0_u1_n82, u0_u0_u1_n83, 
       u0_u0_u1_n84, u0_u0_u1_n85, u0_u0_u1_n86, u0_u0_u1_n87, u0_u0_u1_n88, u0_u0_u1_n89, u0_u0_u1_n9, u0_u0_u1_n90, u0_u0_u1_n91, 
       u0_u0_u1_n92, u0_u0_u1_n93, u0_u0_u1_n94, u0_u0_u2_n1, u0_u0_u2_n10, u0_u0_u2_n11, u0_u0_u2_n12, u0_u0_u2_n13, u0_u0_u2_n14, 
       u0_u0_u2_n15, u0_u0_u2_n16, u0_u0_u2_n17, u0_u0_u2_n18, u0_u0_u2_n19, u0_u0_u2_n2, u0_u0_u2_n20, u0_u0_u2_n21, u0_u0_u2_n22, 
       u0_u0_u2_n23, u0_u0_u2_n24, u0_u0_u2_n25, u0_u0_u2_n26, u0_u0_u2_n27, u0_u0_u2_n28, u0_u0_u2_n29, u0_u0_u2_n3, u0_u0_u2_n30, 
       u0_u0_u2_n31, u0_u0_u2_n32, u0_u0_u2_n33, u0_u0_u2_n34, u0_u0_u2_n35, u0_u0_u2_n36, u0_u0_u2_n37, u0_u0_u2_n38, u0_u0_u2_n39, 
       u0_u0_u2_n4, u0_u0_u2_n40, u0_u0_u2_n41, u0_u0_u2_n42, u0_u0_u2_n43, u0_u0_u2_n44, u0_u0_u2_n45, u0_u0_u2_n46, u0_u0_u2_n47, 
       u0_u0_u2_n48, u0_u0_u2_n49, u0_u0_u2_n5, u0_u0_u2_n50, u0_u0_u2_n51, u0_u0_u2_n52, u0_u0_u2_n53, u0_u0_u2_n54, u0_u0_u2_n55, 
       u0_u0_u2_n56, u0_u0_u2_n57, u0_u0_u2_n58, u0_u0_u2_n59, u0_u0_u2_n6, u0_u0_u2_n60, u0_u0_u2_n61, u0_u0_u2_n62, u0_u0_u2_n63, 
       u0_u0_u2_n64, u0_u0_u2_n65, u0_u0_u2_n66, u0_u0_u2_n67, u0_u0_u2_n68, u0_u0_u2_n69, u0_u0_u2_n7, u0_u0_u2_n70, u0_u0_u2_n71, 
       u0_u0_u2_n72, u0_u0_u2_n73, u0_u0_u2_n74, u0_u0_u2_n75, u0_u0_u2_n76, u0_u0_u2_n77, u0_u0_u2_n78, u0_u0_u2_n79, u0_u0_u2_n8, 
       u0_u0_u2_n80, u0_u0_u2_n81, u0_u0_u2_n82, u0_u0_u2_n83, u0_u0_u2_n84, u0_u0_u2_n85, u0_u0_u2_n86, u0_u0_u2_n87, u0_u0_u2_n88, 
       u0_u0_u2_n89, u0_u0_u2_n9, u0_u0_u2_n90, u0_u0_u2_n91, u0_u0_u2_n92, u0_u0_u2_n93, u0_u0_u2_n94, u0_u0_u3_n1, u0_u0_u3_n10, 
       u0_u0_u3_n11, u0_u0_u3_n12, u0_u0_u3_n13, u0_u0_u3_n14, u0_u0_u3_n15, u0_u0_u3_n16, u0_u0_u3_n17, u0_u0_u3_n18, u0_u0_u3_n19, 
       u0_u0_u3_n2, u0_u0_u3_n20, u0_u0_u3_n21, u0_u0_u3_n22, u0_u0_u3_n23, u0_u0_u3_n24, u0_u0_u3_n25, u0_u0_u3_n26, u0_u0_u3_n27, 
       u0_u0_u3_n28, u0_u0_u3_n29, u0_u0_u3_n3, u0_u0_u3_n30, u0_u0_u3_n31, u0_u0_u3_n32, u0_u0_u3_n33, u0_u0_u3_n34, u0_u0_u3_n35, 
       u0_u0_u3_n36, u0_u0_u3_n37, u0_u0_u3_n38, u0_u0_u3_n39, u0_u0_u3_n4, u0_u0_u3_n40, u0_u0_u3_n41, u0_u0_u3_n42, u0_u0_u3_n43, 
       u0_u0_u3_n44, u0_u0_u3_n45, u0_u0_u3_n46, u0_u0_u3_n47, u0_u0_u3_n48, u0_u0_u3_n49, u0_u0_u3_n5, u0_u0_u3_n50, u0_u0_u3_n51, 
       u0_u0_u3_n52, u0_u0_u3_n53, u0_u0_u3_n54, u0_u0_u3_n55, u0_u0_u3_n56, u0_u0_u3_n57, u0_u0_u3_n58, u0_u0_u3_n59, u0_u0_u3_n6, 
       u0_u0_u3_n60, u0_u0_u3_n61, u0_u0_u3_n62, u0_u0_u3_n63, u0_u0_u3_n64, u0_u0_u3_n65, u0_u0_u3_n66, u0_u0_u3_n67, u0_u0_u3_n68, 
       u0_u0_u3_n69, u0_u0_u3_n7, u0_u0_u3_n70, u0_u0_u3_n71, u0_u0_u3_n72, u0_u0_u3_n73, u0_u0_u3_n74, u0_u0_u3_n75, u0_u0_u3_n76, 
       u0_u0_u3_n77, u0_u0_u3_n78, u0_u0_u3_n79, u0_u0_u3_n8, u0_u0_u3_n80, u0_u0_u3_n81, u0_u0_u3_n82, u0_u0_u3_n83, u0_u0_u3_n84, 
       u0_u0_u3_n85, u0_u0_u3_n86, u0_u0_u3_n87, u0_u0_u3_n88, u0_u0_u3_n89, u0_u0_u3_n9, u0_u0_u3_n90, u0_u0_u3_n91, u0_u0_u3_n92, 
       u0_u0_u3_n93, u0_u13_X_1, u0_u13_X_10, u0_u13_X_11, u0_u13_X_12, u0_u13_X_13, u0_u13_X_14, u0_u13_X_15, u0_u13_X_16, 
       u0_u13_X_17, u0_u13_X_18, u0_u13_X_19, u0_u13_X_2, u0_u13_X_20, u0_u13_X_21, u0_u13_X_22, u0_u13_X_23, u0_u13_X_24, 
       u0_u13_X_25, u0_u13_X_26, u0_u13_X_27, u0_u13_X_28, u0_u13_X_29, u0_u13_X_3, u0_u13_X_30, u0_u13_X_31, u0_u13_X_32, 
       u0_u13_X_33, u0_u13_X_34, u0_u13_X_35, u0_u13_X_36, u0_u13_X_4, u0_u13_X_5, u0_u13_X_6, u0_u13_X_7, u0_u13_X_8, 
       u0_u13_X_9, u0_u13_u0_n100, u0_u13_u0_n101, u0_u13_u0_n102, u0_u13_u0_n103, u0_u13_u0_n104, u0_u13_u0_n105, u0_u13_u0_n106, u0_u13_u0_n107, 
       u0_u13_u0_n108, u0_u13_u0_n109, u0_u13_u0_n110, u0_u13_u0_n111, u0_u13_u0_n112, u0_u13_u0_n113, u0_u13_u0_n114, u0_u13_u0_n115, u0_u13_u0_n116, 
       u0_u13_u0_n117, u0_u13_u0_n118, u0_u13_u0_n119, u0_u13_u0_n120, u0_u13_u0_n121, u0_u13_u0_n122, u0_u13_u0_n123, u0_u13_u0_n124, u0_u13_u0_n125, 
       u0_u13_u0_n126, u0_u13_u0_n127, u0_u13_u0_n128, u0_u13_u0_n129, u0_u13_u0_n130, u0_u13_u0_n131, u0_u13_u0_n132, u0_u13_u0_n133, u0_u13_u0_n134, 
       u0_u13_u0_n135, u0_u13_u0_n136, u0_u13_u0_n137, u0_u13_u0_n138, u0_u13_u0_n139, u0_u13_u0_n140, u0_u13_u0_n141, u0_u13_u0_n142, u0_u13_u0_n143, 
       u0_u13_u0_n144, u0_u13_u0_n145, u0_u13_u0_n146, u0_u13_u0_n147, u0_u13_u0_n148, u0_u13_u0_n149, u0_u13_u0_n150, u0_u13_u0_n151, u0_u13_u0_n152, 
       u0_u13_u0_n153, u0_u13_u0_n154, u0_u13_u0_n155, u0_u13_u0_n156, u0_u13_u0_n157, u0_u13_u0_n158, u0_u13_u0_n159, u0_u13_u0_n160, u0_u13_u0_n161, 
       u0_u13_u0_n162, u0_u13_u0_n163, u0_u13_u0_n164, u0_u13_u0_n165, u0_u13_u0_n166, u0_u13_u0_n167, u0_u13_u0_n168, u0_u13_u0_n169, u0_u13_u0_n170, 
       u0_u13_u0_n171, u0_u13_u0_n172, u0_u13_u0_n173, u0_u13_u0_n174, u0_u13_u0_n88, u0_u13_u0_n89, u0_u13_u0_n90, u0_u13_u0_n91, u0_u13_u0_n92, 
       u0_u13_u0_n93, u0_u13_u0_n94, u0_u13_u0_n95, u0_u13_u0_n96, u0_u13_u0_n97, u0_u13_u0_n98, u0_u13_u0_n99, u0_u13_u1_n100, u0_u13_u1_n101, 
       u0_u13_u1_n102, u0_u13_u1_n103, u0_u13_u1_n104, u0_u13_u1_n105, u0_u13_u1_n106, u0_u13_u1_n107, u0_u13_u1_n108, u0_u13_u1_n109, u0_u13_u1_n110, 
       u0_u13_u1_n111, u0_u13_u1_n112, u0_u13_u1_n113, u0_u13_u1_n114, u0_u13_u1_n115, u0_u13_u1_n116, u0_u13_u1_n117, u0_u13_u1_n118, u0_u13_u1_n119, 
       u0_u13_u1_n120, u0_u13_u1_n121, u0_u13_u1_n122, u0_u13_u1_n123, u0_u13_u1_n124, u0_u13_u1_n125, u0_u13_u1_n126, u0_u13_u1_n127, u0_u13_u1_n128, 
       u0_u13_u1_n129, u0_u13_u1_n130, u0_u13_u1_n131, u0_u13_u1_n132, u0_u13_u1_n133, u0_u13_u1_n134, u0_u13_u1_n135, u0_u13_u1_n136, u0_u13_u1_n137, 
       u0_u13_u1_n138, u0_u13_u1_n139, u0_u13_u1_n140, u0_u13_u1_n141, u0_u13_u1_n142, u0_u13_u1_n143, u0_u13_u1_n144, u0_u13_u1_n145, u0_u13_u1_n146, 
       u0_u13_u1_n147, u0_u13_u1_n148, u0_u13_u1_n149, u0_u13_u1_n150, u0_u13_u1_n151, u0_u13_u1_n152, u0_u13_u1_n153, u0_u13_u1_n154, u0_u13_u1_n155, 
       u0_u13_u1_n156, u0_u13_u1_n157, u0_u13_u1_n158, u0_u13_u1_n159, u0_u13_u1_n160, u0_u13_u1_n161, u0_u13_u1_n162, u0_u13_u1_n163, u0_u13_u1_n164, 
       u0_u13_u1_n165, u0_u13_u1_n166, u0_u13_u1_n167, u0_u13_u1_n168, u0_u13_u1_n169, u0_u13_u1_n170, u0_u13_u1_n171, u0_u13_u1_n172, u0_u13_u1_n173, 
       u0_u13_u1_n174, u0_u13_u1_n175, u0_u13_u1_n176, u0_u13_u1_n177, u0_u13_u1_n178, u0_u13_u1_n179, u0_u13_u1_n180, u0_u13_u1_n181, u0_u13_u1_n182, 
       u0_u13_u1_n183, u0_u13_u1_n184, u0_u13_u1_n185, u0_u13_u1_n186, u0_u13_u1_n187, u0_u13_u1_n188, u0_u13_u1_n95, u0_u13_u1_n96, u0_u13_u1_n97, 
       u0_u13_u1_n98, u0_u13_u1_n99, u0_u13_u2_n100, u0_u13_u2_n101, u0_u13_u2_n102, u0_u13_u2_n103, u0_u13_u2_n104, u0_u13_u2_n105, u0_u13_u2_n106, 
       u0_u13_u2_n107, u0_u13_u2_n108, u0_u13_u2_n109, u0_u13_u2_n110, u0_u13_u2_n111, u0_u13_u2_n112, u0_u13_u2_n113, u0_u13_u2_n114, u0_u13_u2_n115, 
       u0_u13_u2_n116, u0_u13_u2_n117, u0_u13_u2_n118, u0_u13_u2_n119, u0_u13_u2_n120, u0_u13_u2_n121, u0_u13_u2_n122, u0_u13_u2_n123, u0_u13_u2_n124, 
       u0_u13_u2_n125, u0_u13_u2_n126, u0_u13_u2_n127, u0_u13_u2_n128, u0_u13_u2_n129, u0_u13_u2_n130, u0_u13_u2_n131, u0_u13_u2_n132, u0_u13_u2_n133, 
       u0_u13_u2_n134, u0_u13_u2_n135, u0_u13_u2_n136, u0_u13_u2_n137, u0_u13_u2_n138, u0_u13_u2_n139, u0_u13_u2_n140, u0_u13_u2_n141, u0_u13_u2_n142, 
       u0_u13_u2_n143, u0_u13_u2_n144, u0_u13_u2_n145, u0_u13_u2_n146, u0_u13_u2_n147, u0_u13_u2_n148, u0_u13_u2_n149, u0_u13_u2_n150, u0_u13_u2_n151, 
       u0_u13_u2_n152, u0_u13_u2_n153, u0_u13_u2_n154, u0_u13_u2_n155, u0_u13_u2_n156, u0_u13_u2_n157, u0_u13_u2_n158, u0_u13_u2_n159, u0_u13_u2_n160, 
       u0_u13_u2_n161, u0_u13_u2_n162, u0_u13_u2_n163, u0_u13_u2_n164, u0_u13_u2_n165, u0_u13_u2_n166, u0_u13_u2_n167, u0_u13_u2_n168, u0_u13_u2_n169, 
       u0_u13_u2_n170, u0_u13_u2_n171, u0_u13_u2_n172, u0_u13_u2_n173, u0_u13_u2_n174, u0_u13_u2_n175, u0_u13_u2_n176, u0_u13_u2_n177, u0_u13_u2_n178, 
       u0_u13_u2_n179, u0_u13_u2_n180, u0_u13_u2_n181, u0_u13_u2_n182, u0_u13_u2_n183, u0_u13_u2_n184, u0_u13_u2_n185, u0_u13_u2_n186, u0_u13_u2_n187, 
       u0_u13_u2_n188, u0_u13_u2_n95, u0_u13_u2_n96, u0_u13_u2_n97, u0_u13_u2_n98, u0_u13_u2_n99, u0_u13_u3_n100, u0_u13_u3_n101, u0_u13_u3_n102, 
       u0_u13_u3_n103, u0_u13_u3_n104, u0_u13_u3_n105, u0_u13_u3_n106, u0_u13_u3_n107, u0_u13_u3_n108, u0_u13_u3_n109, u0_u13_u3_n110, u0_u13_u3_n111, 
       u0_u13_u3_n112, u0_u13_u3_n113, u0_u13_u3_n114, u0_u13_u3_n115, u0_u13_u3_n116, u0_u13_u3_n117, u0_u13_u3_n118, u0_u13_u3_n119, u0_u13_u3_n120, 
       u0_u13_u3_n121, u0_u13_u3_n122, u0_u13_u3_n123, u0_u13_u3_n124, u0_u13_u3_n125, u0_u13_u3_n126, u0_u13_u3_n127, u0_u13_u3_n128, u0_u13_u3_n129, 
       u0_u13_u3_n130, u0_u13_u3_n131, u0_u13_u3_n132, u0_u13_u3_n133, u0_u13_u3_n134, u0_u13_u3_n135, u0_u13_u3_n136, u0_u13_u3_n137, u0_u13_u3_n138, 
       u0_u13_u3_n139, u0_u13_u3_n140, u0_u13_u3_n141, u0_u13_u3_n142, u0_u13_u3_n143, u0_u13_u3_n144, u0_u13_u3_n145, u0_u13_u3_n146, u0_u13_u3_n147, 
       u0_u13_u3_n148, u0_u13_u3_n149, u0_u13_u3_n150, u0_u13_u3_n151, u0_u13_u3_n152, u0_u13_u3_n153, u0_u13_u3_n154, u0_u13_u3_n155, u0_u13_u3_n156, 
       u0_u13_u3_n157, u0_u13_u3_n158, u0_u13_u3_n159, u0_u13_u3_n160, u0_u13_u3_n161, u0_u13_u3_n162, u0_u13_u3_n163, u0_u13_u3_n164, u0_u13_u3_n165, 
       u0_u13_u3_n166, u0_u13_u3_n167, u0_u13_u3_n168, u0_u13_u3_n169, u0_u13_u3_n170, u0_u13_u3_n171, u0_u13_u3_n172, u0_u13_u3_n173, u0_u13_u3_n174, 
       u0_u13_u3_n175, u0_u13_u3_n176, u0_u13_u3_n177, u0_u13_u3_n178, u0_u13_u3_n179, u0_u13_u3_n180, u0_u13_u3_n181, u0_u13_u3_n182, u0_u13_u3_n183, 
       u0_u13_u3_n184, u0_u13_u3_n185, u0_u13_u3_n186, u0_u13_u3_n94, u0_u13_u3_n95, u0_u13_u3_n96, u0_u13_u3_n97, u0_u13_u3_n98, u0_u13_u3_n99, 
       u0_u13_u4_n100, u0_u13_u4_n101, u0_u13_u4_n102, u0_u13_u4_n103, u0_u13_u4_n104, u0_u13_u4_n105, u0_u13_u4_n106, u0_u13_u4_n107, u0_u13_u4_n108, 
       u0_u13_u4_n109, u0_u13_u4_n110, u0_u13_u4_n111, u0_u13_u4_n112, u0_u13_u4_n113, u0_u13_u4_n114, u0_u13_u4_n115, u0_u13_u4_n116, u0_u13_u4_n117, 
       u0_u13_u4_n118, u0_u13_u4_n119, u0_u13_u4_n120, u0_u13_u4_n121, u0_u13_u4_n122, u0_u13_u4_n123, u0_u13_u4_n124, u0_u13_u4_n125, u0_u13_u4_n126, 
       u0_u13_u4_n127, u0_u13_u4_n128, u0_u13_u4_n129, u0_u13_u4_n130, u0_u13_u4_n131, u0_u13_u4_n132, u0_u13_u4_n133, u0_u13_u4_n134, u0_u13_u4_n135, 
       u0_u13_u4_n136, u0_u13_u4_n137, u0_u13_u4_n138, u0_u13_u4_n139, u0_u13_u4_n140, u0_u13_u4_n141, u0_u13_u4_n142, u0_u13_u4_n143, u0_u13_u4_n144, 
       u0_u13_u4_n145, u0_u13_u4_n146, u0_u13_u4_n147, u0_u13_u4_n148, u0_u13_u4_n149, u0_u13_u4_n150, u0_u13_u4_n151, u0_u13_u4_n152, u0_u13_u4_n153, 
       u0_u13_u4_n154, u0_u13_u4_n155, u0_u13_u4_n156, u0_u13_u4_n157, u0_u13_u4_n158, u0_u13_u4_n159, u0_u13_u4_n160, u0_u13_u4_n161, u0_u13_u4_n162, 
       u0_u13_u4_n163, u0_u13_u4_n164, u0_u13_u4_n165, u0_u13_u4_n166, u0_u13_u4_n167, u0_u13_u4_n168, u0_u13_u4_n169, u0_u13_u4_n170, u0_u13_u4_n171, 
       u0_u13_u4_n172, u0_u13_u4_n173, u0_u13_u4_n174, u0_u13_u4_n175, u0_u13_u4_n176, u0_u13_u4_n177, u0_u13_u4_n178, u0_u13_u4_n179, u0_u13_u4_n180, 
       u0_u13_u4_n181, u0_u13_u4_n182, u0_u13_u4_n183, u0_u13_u4_n184, u0_u13_u4_n185, u0_u13_u4_n186, u0_u13_u4_n94, u0_u13_u4_n95, u0_u13_u4_n96, 
       u0_u13_u4_n97, u0_u13_u4_n98, u0_u13_u4_n99, u0_u13_u5_n100, u0_u13_u5_n101, u0_u13_u5_n102, u0_u13_u5_n103, u0_u13_u5_n104, u0_u13_u5_n105, 
       u0_u13_u5_n106, u0_u13_u5_n107, u0_u13_u5_n108, u0_u13_u5_n109, u0_u13_u5_n110, u0_u13_u5_n111, u0_u13_u5_n112, u0_u13_u5_n113, u0_u13_u5_n114, 
       u0_u13_u5_n115, u0_u13_u5_n116, u0_u13_u5_n117, u0_u13_u5_n118, u0_u13_u5_n119, u0_u13_u5_n120, u0_u13_u5_n121, u0_u13_u5_n122, u0_u13_u5_n123, 
       u0_u13_u5_n124, u0_u13_u5_n125, u0_u13_u5_n126, u0_u13_u5_n127, u0_u13_u5_n128, u0_u13_u5_n129, u0_u13_u5_n130, u0_u13_u5_n131, u0_u13_u5_n132, 
       u0_u13_u5_n133, u0_u13_u5_n134, u0_u13_u5_n135, u0_u13_u5_n136, u0_u13_u5_n137, u0_u13_u5_n138, u0_u13_u5_n139, u0_u13_u5_n140, u0_u13_u5_n141, 
       u0_u13_u5_n142, u0_u13_u5_n143, u0_u13_u5_n144, u0_u13_u5_n145, u0_u13_u5_n146, u0_u13_u5_n147, u0_u13_u5_n148, u0_u13_u5_n149, u0_u13_u5_n150, 
       u0_u13_u5_n151, u0_u13_u5_n152, u0_u13_u5_n153, u0_u13_u5_n154, u0_u13_u5_n155, u0_u13_u5_n156, u0_u13_u5_n157, u0_u13_u5_n158, u0_u13_u5_n159, 
       u0_u13_u5_n160, u0_u13_u5_n161, u0_u13_u5_n162, u0_u13_u5_n163, u0_u13_u5_n164, u0_u13_u5_n165, u0_u13_u5_n166, u0_u13_u5_n167, u0_u13_u5_n168, 
       u0_u13_u5_n169, u0_u13_u5_n170, u0_u13_u5_n171, u0_u13_u5_n172, u0_u13_u5_n173, u0_u13_u5_n174, u0_u13_u5_n175, u0_u13_u5_n176, u0_u13_u5_n177, 
       u0_u13_u5_n178, u0_u13_u5_n179, u0_u13_u5_n180, u0_u13_u5_n181, u0_u13_u5_n182, u0_u13_u5_n183, u0_u13_u5_n184, u0_u13_u5_n185, u0_u13_u5_n186, 
       u0_u13_u5_n187, u0_u13_u5_n188, u0_u13_u5_n189, u0_u13_u5_n190, u0_u13_u5_n191, u0_u13_u5_n192, u0_u13_u5_n193, u0_u13_u5_n194, u0_u13_u5_n195, 
       u0_u13_u5_n196, u0_u13_u5_n99, u0_u4_X_10, u0_u4_X_11, u0_u4_X_12, u0_u4_X_13, u0_u4_X_14, u0_u4_X_15, u0_u4_X_16, 
       u0_u4_X_17, u0_u4_X_18, u0_u4_X_19, u0_u4_X_20, u0_u4_X_21, u0_u4_X_22, u0_u4_X_23, u0_u4_X_24, u0_u4_X_7, 
       u0_u4_X_8, u0_u4_X_9, u0_u4_u1_n100, u0_u4_u1_n101, u0_u4_u1_n102, u0_u4_u1_n103, u0_u4_u1_n104, u0_u4_u1_n105, u0_u4_u1_n106, 
       u0_u4_u1_n107, u0_u4_u1_n108, u0_u4_u1_n109, u0_u4_u1_n110, u0_u4_u1_n111, u0_u4_u1_n112, u0_u4_u1_n113, u0_u4_u1_n114, u0_u4_u1_n115, 
       u0_u4_u1_n116, u0_u4_u1_n117, u0_u4_u1_n118, u0_u4_u1_n119, u0_u4_u1_n120, u0_u4_u1_n121, u0_u4_u1_n122, u0_u4_u1_n123, u0_u4_u1_n124, 
       u0_u4_u1_n125, u0_u4_u1_n126, u0_u4_u1_n127, u0_u4_u1_n128, u0_u4_u1_n129, u0_u4_u1_n130, u0_u4_u1_n131, u0_u4_u1_n132, u0_u4_u1_n133, 
       u0_u4_u1_n134, u0_u4_u1_n135, u0_u4_u1_n136, u0_u4_u1_n137, u0_u4_u1_n138, u0_u4_u1_n139, u0_u4_u1_n140, u0_u4_u1_n141, u0_u4_u1_n142, 
       u0_u4_u1_n143, u0_u4_u1_n144, u0_u4_u1_n145, u0_u4_u1_n146, u0_u4_u1_n147, u0_u4_u1_n148, u0_u4_u1_n149, u0_u4_u1_n150, u0_u4_u1_n151, 
       u0_u4_u1_n152, u0_u4_u1_n153, u0_u4_u1_n154, u0_u4_u1_n155, u0_u4_u1_n156, u0_u4_u1_n157, u0_u4_u1_n158, u0_u4_u1_n159, u0_u4_u1_n160, 
       u0_u4_u1_n161, u0_u4_u1_n162, u0_u4_u1_n163, u0_u4_u1_n164, u0_u4_u1_n165, u0_u4_u1_n166, u0_u4_u1_n167, u0_u4_u1_n168, u0_u4_u1_n169, 
       u0_u4_u1_n170, u0_u4_u1_n171, u0_u4_u1_n172, u0_u4_u1_n173, u0_u4_u1_n174, u0_u4_u1_n175, u0_u4_u1_n176, u0_u4_u1_n177, u0_u4_u1_n178, 
       u0_u4_u1_n179, u0_u4_u1_n180, u0_u4_u1_n181, u0_u4_u1_n182, u0_u4_u1_n183, u0_u4_u1_n184, u0_u4_u1_n185, u0_u4_u1_n186, u0_u4_u1_n187, 
       u0_u4_u1_n188, u0_u4_u1_n95, u0_u4_u1_n96, u0_u4_u1_n97, u0_u4_u1_n98, u0_u4_u1_n99, u0_u4_u2_n100, u0_u4_u2_n101, u0_u4_u2_n102, 
       u0_u4_u2_n103, u0_u4_u2_n104, u0_u4_u2_n105, u0_u4_u2_n106, u0_u4_u2_n107, u0_u4_u2_n108, u0_u4_u2_n109, u0_u4_u2_n110, u0_u4_u2_n111, 
       u0_u4_u2_n112, u0_u4_u2_n113, u0_u4_u2_n114, u0_u4_u2_n115, u0_u4_u2_n116, u0_u4_u2_n117, u0_u4_u2_n118, u0_u4_u2_n119, u0_u4_u2_n120, 
       u0_u4_u2_n121, u0_u4_u2_n122, u0_u4_u2_n123, u0_u4_u2_n124, u0_u4_u2_n125, u0_u4_u2_n126, u0_u4_u2_n127, u0_u4_u2_n128, u0_u4_u2_n129, 
       u0_u4_u2_n130, u0_u4_u2_n131, u0_u4_u2_n132, u0_u4_u2_n133, u0_u4_u2_n134, u0_u4_u2_n135, u0_u4_u2_n136, u0_u4_u2_n137, u0_u4_u2_n138, 
       u0_u4_u2_n139, u0_u4_u2_n140, u0_u4_u2_n141, u0_u4_u2_n142, u0_u4_u2_n143, u0_u4_u2_n144, u0_u4_u2_n145, u0_u4_u2_n146, u0_u4_u2_n147, 
       u0_u4_u2_n148, u0_u4_u2_n149, u0_u4_u2_n150, u0_u4_u2_n151, u0_u4_u2_n152, u0_u4_u2_n153, u0_u4_u2_n154, u0_u4_u2_n155, u0_u4_u2_n156, 
       u0_u4_u2_n157, u0_u4_u2_n158, u0_u4_u2_n159, u0_u4_u2_n160, u0_u4_u2_n161, u0_u4_u2_n162, u0_u4_u2_n163, u0_u4_u2_n164, u0_u4_u2_n165, 
       u0_u4_u2_n166, u0_u4_u2_n167, u0_u4_u2_n168, u0_u4_u2_n169, u0_u4_u2_n170, u0_u4_u2_n171, u0_u4_u2_n172, u0_u4_u2_n173, u0_u4_u2_n174, 
       u0_u4_u2_n175, u0_u4_u2_n176, u0_u4_u2_n177, u0_u4_u2_n178, u0_u4_u2_n179, u0_u4_u2_n180, u0_u4_u2_n181, u0_u4_u2_n182, u0_u4_u2_n183, 
       u0_u4_u2_n184, u0_u4_u2_n185, u0_u4_u2_n186, u0_u4_u2_n187, u0_u4_u2_n188, u0_u4_u2_n95, u0_u4_u2_n96, u0_u4_u2_n97, u0_u4_u2_n98, 
       u0_u4_u2_n99, u0_u4_u3_n100, u0_u4_u3_n101, u0_u4_u3_n102, u0_u4_u3_n103, u0_u4_u3_n104, u0_u4_u3_n105, u0_u4_u3_n106, u0_u4_u3_n107, 
       u0_u4_u3_n108, u0_u4_u3_n109, u0_u4_u3_n110, u0_u4_u3_n111, u0_u4_u3_n112, u0_u4_u3_n113, u0_u4_u3_n114, u0_u4_u3_n115, u0_u4_u3_n116, 
       u0_u4_u3_n117, u0_u4_u3_n118, u0_u4_u3_n119, u0_u4_u3_n120, u0_u4_u3_n121, u0_u4_u3_n122, u0_u4_u3_n123, u0_u4_u3_n124, u0_u4_u3_n125, 
       u0_u4_u3_n126, u0_u4_u3_n127, u0_u4_u3_n128, u0_u4_u3_n129, u0_u4_u3_n130, u0_u4_u3_n131, u0_u4_u3_n132, u0_u4_u3_n133, u0_u4_u3_n134, 
       u0_u4_u3_n135, u0_u4_u3_n136, u0_u4_u3_n137, u0_u4_u3_n138, u0_u4_u3_n139, u0_u4_u3_n140, u0_u4_u3_n141, u0_u4_u3_n142, u0_u4_u3_n143, 
       u0_u4_u3_n144, u0_u4_u3_n145, u0_u4_u3_n146, u0_u4_u3_n147, u0_u4_u3_n148, u0_u4_u3_n149, u0_u4_u3_n150, u0_u4_u3_n151, u0_u4_u3_n152, 
       u0_u4_u3_n153, u0_u4_u3_n154, u0_u4_u3_n155, u0_u4_u3_n156, u0_u4_u3_n157, u0_u4_u3_n158, u0_u4_u3_n159, u0_u4_u3_n160, u0_u4_u3_n161, 
       u0_u4_u3_n162, u0_u4_u3_n163, u0_u4_u3_n164, u0_u4_u3_n165, u0_u4_u3_n166, u0_u4_u3_n167, u0_u4_u3_n168, u0_u4_u3_n169, u0_u4_u3_n170, 
       u0_u4_u3_n171, u0_u4_u3_n172, u0_u4_u3_n173, u0_u4_u3_n174, u0_u4_u3_n175, u0_u4_u3_n176, u0_u4_u3_n177, u0_u4_u3_n178, u0_u4_u3_n179, 
       u0_u4_u3_n180, u0_u4_u3_n181, u0_u4_u3_n182, u0_u4_u3_n183, u0_u4_u3_n184, u0_u4_u3_n185, u0_u4_u3_n186, u0_u4_u3_n94, u0_u4_u3_n95, 
       u0_u4_u3_n96, u0_u4_u3_n97, u0_u4_u3_n98, u0_u4_u3_n99, u0_uk_n673, u0_uk_n679, u0_uk_n683, u0_uk_n699, u0_uk_n703, 
       u0_uk_n704, u0_uk_n708, u0_uk_n712, u0_uk_n713, u0_uk_n802, u0_uk_n816, u0_uk_n818, u0_uk_n869, u0_uk_n881, 
       u0_uk_n885, u0_uk_n886, u0_uk_n887, u0_uk_n891, u0_uk_n892, u0_uk_n893, u0_uk_n927, u0_uk_n932, u0_uk_n933, 
       u0_uk_n934, u0_uk_n935, u0_uk_n938, u2_K10_1, u2_K10_12, u2_K10_13, u2_K10_14, u2_K10_16, u2_K10_18, 
       u2_K10_2, u2_K10_3, u2_K10_45, u2_K10_47, u2_K10_48, u2_K10_5, u2_K10_7, u2_K10_8, u2_K10_9, 
       u2_K12_1, u2_K12_10, u2_K12_11, u2_K12_12, u2_K12_13, u2_K12_14, u2_K12_15, u2_K12_16, u2_K12_17, 
       u2_K12_18, u2_K12_3, u2_K12_4, u2_K12_5, u2_K12_6, u2_K12_7, u2_K12_9, u2_K14_26, u2_K14_27, 
       u2_K14_29, u2_K14_30, u2_K14_31, u2_K14_32, u2_K14_33, u2_K14_34, u2_K14_35, u2_K14_36, u2_K15_10, 
       u2_K15_11, u2_K15_12, u2_K15_25, u2_K15_26, u2_K15_27, u2_K15_3, u2_K15_30, u2_K15_32, u2_K15_33, 
       u2_K15_36, u2_K15_37, u2_K15_38, u2_K15_4, u2_K15_40, u2_K15_41, u2_K15_42, u2_K15_6, u2_K15_7, 
       u2_K15_8, u2_K15_9, u2_K16_1, u2_K16_2, u2_K16_25, u2_K16_27, u2_K16_28, u2_K16_29, u2_K16_3, 
       u2_K16_30, u2_K16_32, u2_K16_33, u2_K16_34, u2_K16_35, u2_K16_36, u2_K16_37, u2_K16_38, u2_K16_39, 
       u2_K16_4, u2_K16_40, u2_K16_41, u2_K16_43, u2_K16_45, u2_K16_46, u2_K16_48, u2_K1_1, u2_K1_10, 
       u2_K1_11, u2_K1_12, u2_K1_13, u2_K1_14, u2_K1_17, u2_K1_18, u2_K1_2, u2_K1_20, u2_K1_21, 
       u2_K1_22, u2_K1_23, u2_K1_3, u2_K1_4, u2_K1_6, u2_K1_7, u2_K1_8, u2_K2_25, u2_K2_26, 
       u2_K2_27, u2_K2_28, u2_K2_29, u2_K2_30, u2_K2_37, u2_K2_38, u2_K2_39, u2_K2_41, u2_K2_42, 
       u2_K3_1, u2_K3_10, u2_K3_11, u2_K3_12, u2_K3_14, u2_K3_17, u2_K3_18, u2_K3_19, u2_K3_2, 
       u2_K3_21, u2_K3_22, u2_K3_24, u2_K3_3, u2_K3_31, u2_K3_33, u2_K3_34, u2_K3_36, u2_K3_37, 
       u2_K3_38, u2_K3_39, u2_K3_4, u2_K3_40, u2_K3_41, u2_K3_44, u2_K3_45, u2_K3_46, u2_K3_5, 
       u2_K3_6, u2_K3_8, u2_K3_9, u2_K4_13, u2_K4_15, u2_K4_16, u2_K4_17, u2_K4_18, u2_K4_19, 
       u2_K4_20, u2_K4_23, u2_K4_24, u2_K4_25, u2_K4_26, u2_K4_28, u2_K4_29, u2_K4_30, u2_K4_31, 
       u2_K4_32, u2_K4_36, u2_K5_12, u2_K5_15, u2_K5_20, u2_K5_22, u2_K5_7, u2_K6_19, u2_K6_21, 
       u2_K6_23, u2_K6_26, u2_K6_28, u2_K6_29, u2_K6_30, u2_K7_1, u2_K7_10, u2_K7_11, u2_K7_12, 
       u2_K7_13, u2_K7_14, u2_K7_15, u2_K7_16, u2_K7_17, u2_K7_18, u2_K7_19, u2_K7_2, u2_K7_20, 
       u2_K7_21, u2_K7_22, u2_K7_23, u2_K7_24, u2_K7_25, u2_K7_27, u2_K7_28, u2_K7_29, u2_K7_30, 
       u2_K7_39, u2_K7_40, u2_K7_41, u2_K7_42, u2_K7_44, u2_K7_46, u2_K7_47, u2_K7_6, u2_K7_8, 
       u2_K7_9, u2_K8_37, u2_K8_38, u2_K8_39, u2_K8_40, u2_K8_42, u2_K8_43, u2_K8_44, u2_K8_46, 
       u2_K8_47, u2_K8_48, u2_out0_1, u2_out0_10, u2_out0_13, u2_out0_16, u2_out0_17, u2_out0_18, u2_out0_2, 
       u2_out0_20, u2_out0_23, u2_out0_24, u2_out0_26, u2_out0_28, u2_out0_30, u2_out0_31, u2_out0_6, u2_out0_9, 
       u2_out11_13, u2_out11_16, u2_out11_17, u2_out11_18, u2_out11_2, u2_out11_23, u2_out11_24, u2_out11_28, u2_out11_30, 
       u2_out11_31, u2_out11_6, u2_out11_9, u2_out13_11, u2_out13_14, u2_out13_19, u2_out13_25, u2_out13_29, u2_out13_3, 
       u2_out13_4, u2_out13_8, u2_out14_11, u2_out14_12, u2_out14_13, u2_out14_14, u2_out14_17, u2_out14_18, u2_out14_19, 
       u2_out14_2, u2_out14_22, u2_out14_23, u2_out14_25, u2_out14_28, u2_out14_29, u2_out14_3, u2_out14_31, u2_out14_32, 
       u2_out14_4, u2_out14_7, u2_out14_8, u2_out14_9, u2_out15_11, u2_out15_12, u2_out15_14, u2_out15_15, u2_out15_17, 
       u2_out15_19, u2_out15_21, u2_out15_22, u2_out15_23, u2_out15_25, u2_out15_27, u2_out15_29, u2_out15_3, u2_out15_31, 
       u2_out15_32, u2_out15_4, u2_out15_5, u2_out15_7, u2_out15_8, u2_out15_9, u2_out1_12, u2_out1_14, u2_out1_22, 
       u2_out1_25, u2_out1_3, u2_out1_32, u2_out1_7, u2_out1_8, u2_out2_1, u2_out2_10, u2_out2_11, u2_out2_12, 
       u2_out2_13, u2_out2_15, u2_out2_16, u2_out2_17, u2_out2_18, u2_out2_19, u2_out2_2, u2_out2_20, u2_out2_21, 
       u2_out2_22, u2_out2_23, u2_out2_24, u2_out2_26, u2_out2_27, u2_out2_28, u2_out2_29, u2_out2_30, u2_out2_31, 
       u2_out2_32, u2_out2_4, u2_out2_5, u2_out2_6, u2_out2_7, u2_out2_9, u2_out3_1, u2_out3_10, u2_out3_11, 
       u2_out3_14, u2_out3_16, u2_out3_19, u2_out3_20, u2_out3_24, u2_out3_25, u2_out3_26, u2_out3_29, u2_out3_3, 
       u2_out3_30, u2_out3_4, u2_out3_6, u2_out3_8, u2_out4_1, u2_out4_10, u2_out4_13, u2_out4_16, u2_out4_18, 
       u2_out4_2, u2_out4_20, u2_out4_24, u2_out4_26, u2_out4_28, u2_out4_30, u2_out4_6, u2_out5_1, u2_out5_10, 
       u2_out5_14, u2_out5_20, u2_out5_25, u2_out5_26, u2_out5_3, u2_out5_8, u2_out6_1, u2_out6_10, u2_out6_12, 
       u2_out6_13, u2_out6_14, u2_out6_15, u2_out6_16, u2_out6_17, u2_out6_18, u2_out6_2, u2_out6_20, u2_out6_21, 
       u2_out6_22, u2_out6_23, u2_out6_24, u2_out6_25, u2_out6_26, u2_out6_27, u2_out6_28, u2_out6_3, u2_out6_30, 
       u2_out6_31, u2_out6_32, u2_out6_5, u2_out6_6, u2_out6_7, u2_out6_8, u2_out6_9, u2_out7_12, u2_out7_15, 
       u2_out7_21, u2_out7_22, u2_out7_27, u2_out7_32, u2_out7_5, u2_out7_7, u2_out9_13, u2_out9_15, u2_out9_16, 
       u2_out9_17, u2_out9_18, u2_out9_2, u2_out9_21, u2_out9_23, u2_out9_24, u2_out9_27, u2_out9_28, u2_out9_30, 
       u2_out9_31, u2_out9_5, u2_out9_6, u2_out9_9, u2_u0_X_1, u2_u0_X_10, u2_u0_X_11, u2_u0_X_12, u2_u0_X_13, 
       u2_u0_X_14, u2_u0_X_15, u2_u0_X_16, u2_u0_X_17, u2_u0_X_18, u2_u0_X_19, u2_u0_X_2, u2_u0_X_20, u2_u0_X_21, 
       u2_u0_X_22, u2_u0_X_23, u2_u0_X_24, u2_u0_X_3, u2_u0_X_4, u2_u0_X_5, u2_u0_X_6, u2_u0_X_7, u2_u0_X_8, 
       u2_u0_X_9, u2_u0_u0_n100, u2_u0_u0_n101, u2_u0_u0_n102, u2_u0_u0_n103, u2_u0_u0_n104, u2_u0_u0_n105, u2_u0_u0_n106, u2_u0_u0_n107, 
       u2_u0_u0_n108, u2_u0_u0_n109, u2_u0_u0_n110, u2_u0_u0_n111, u2_u0_u0_n112, u2_u0_u0_n113, u2_u0_u0_n114, u2_u0_u0_n115, u2_u0_u0_n116, 
       u2_u0_u0_n117, u2_u0_u0_n118, u2_u0_u0_n119, u2_u0_u0_n120, u2_u0_u0_n121, u2_u0_u0_n122, u2_u0_u0_n123, u2_u0_u0_n124, u2_u0_u0_n125, 
       u2_u0_u0_n126, u2_u0_u0_n127, u2_u0_u0_n128, u2_u0_u0_n129, u2_u0_u0_n130, u2_u0_u0_n131, u2_u0_u0_n132, u2_u0_u0_n133, u2_u0_u0_n134, 
       u2_u0_u0_n135, u2_u0_u0_n136, u2_u0_u0_n137, u2_u0_u0_n138, u2_u0_u0_n139, u2_u0_u0_n140, u2_u0_u0_n141, u2_u0_u0_n142, u2_u0_u0_n143, 
       u2_u0_u0_n144, u2_u0_u0_n145, u2_u0_u0_n146, u2_u0_u0_n147, u2_u0_u0_n148, u2_u0_u0_n149, u2_u0_u0_n150, u2_u0_u0_n151, u2_u0_u0_n152, 
       u2_u0_u0_n153, u2_u0_u0_n154, u2_u0_u0_n155, u2_u0_u0_n156, u2_u0_u0_n157, u2_u0_u0_n158, u2_u0_u0_n159, u2_u0_u0_n160, u2_u0_u0_n161, 
       u2_u0_u0_n162, u2_u0_u0_n163, u2_u0_u0_n164, u2_u0_u0_n165, u2_u0_u0_n166, u2_u0_u0_n167, u2_u0_u0_n168, u2_u0_u0_n169, u2_u0_u0_n170, 
       u2_u0_u0_n171, u2_u0_u0_n172, u2_u0_u0_n173, u2_u0_u0_n174, u2_u0_u0_n88, u2_u0_u0_n89, u2_u0_u0_n90, u2_u0_u0_n91, u2_u0_u0_n92, 
       u2_u0_u0_n93, u2_u0_u0_n94, u2_u0_u0_n95, u2_u0_u0_n96, u2_u0_u0_n97, u2_u0_u0_n98, u2_u0_u0_n99, u2_u0_u1_n100, u2_u0_u1_n101, 
       u2_u0_u1_n102, u2_u0_u1_n103, u2_u0_u1_n104, u2_u0_u1_n105, u2_u0_u1_n106, u2_u0_u1_n107, u2_u0_u1_n108, u2_u0_u1_n109, u2_u0_u1_n110, 
       u2_u0_u1_n111, u2_u0_u1_n112, u2_u0_u1_n113, u2_u0_u1_n114, u2_u0_u1_n115, u2_u0_u1_n116, u2_u0_u1_n117, u2_u0_u1_n118, u2_u0_u1_n119, 
       u2_u0_u1_n120, u2_u0_u1_n121, u2_u0_u1_n122, u2_u0_u1_n123, u2_u0_u1_n124, u2_u0_u1_n125, u2_u0_u1_n126, u2_u0_u1_n127, u2_u0_u1_n128, 
       u2_u0_u1_n129, u2_u0_u1_n130, u2_u0_u1_n131, u2_u0_u1_n132, u2_u0_u1_n133, u2_u0_u1_n134, u2_u0_u1_n135, u2_u0_u1_n136, u2_u0_u1_n137, 
       u2_u0_u1_n138, u2_u0_u1_n139, u2_u0_u1_n140, u2_u0_u1_n141, u2_u0_u1_n142, u2_u0_u1_n143, u2_u0_u1_n144, u2_u0_u1_n145, u2_u0_u1_n146, 
       u2_u0_u1_n147, u2_u0_u1_n148, u2_u0_u1_n149, u2_u0_u1_n150, u2_u0_u1_n151, u2_u0_u1_n152, u2_u0_u1_n153, u2_u0_u1_n154, u2_u0_u1_n155, 
       u2_u0_u1_n156, u2_u0_u1_n157, u2_u0_u1_n158, u2_u0_u1_n159, u2_u0_u1_n160, u2_u0_u1_n161, u2_u0_u1_n162, u2_u0_u1_n163, u2_u0_u1_n164, 
       u2_u0_u1_n165, u2_u0_u1_n166, u2_u0_u1_n167, u2_u0_u1_n168, u2_u0_u1_n169, u2_u0_u1_n170, u2_u0_u1_n171, u2_u0_u1_n172, u2_u0_u1_n173, 
       u2_u0_u1_n174, u2_u0_u1_n175, u2_u0_u1_n176, u2_u0_u1_n177, u2_u0_u1_n178, u2_u0_u1_n179, u2_u0_u1_n180, u2_u0_u1_n181, u2_u0_u1_n182, 
       u2_u0_u1_n183, u2_u0_u1_n184, u2_u0_u1_n185, u2_u0_u1_n186, u2_u0_u1_n187, u2_u0_u1_n188, u2_u0_u1_n95, u2_u0_u1_n96, u2_u0_u1_n97, 
       u2_u0_u1_n98, u2_u0_u1_n99, u2_u0_u2_n100, u2_u0_u2_n101, u2_u0_u2_n102, u2_u0_u2_n103, u2_u0_u2_n104, u2_u0_u2_n105, u2_u0_u2_n106, 
       u2_u0_u2_n107, u2_u0_u2_n108, u2_u0_u2_n109, u2_u0_u2_n110, u2_u0_u2_n111, u2_u0_u2_n112, u2_u0_u2_n113, u2_u0_u2_n114, u2_u0_u2_n115, 
       u2_u0_u2_n116, u2_u0_u2_n117, u2_u0_u2_n118, u2_u0_u2_n119, u2_u0_u2_n120, u2_u0_u2_n121, u2_u0_u2_n122, u2_u0_u2_n123, u2_u0_u2_n124, 
       u2_u0_u2_n125, u2_u0_u2_n126, u2_u0_u2_n127, u2_u0_u2_n128, u2_u0_u2_n129, u2_u0_u2_n130, u2_u0_u2_n131, u2_u0_u2_n132, u2_u0_u2_n133, 
       u2_u0_u2_n134, u2_u0_u2_n135, u2_u0_u2_n136, u2_u0_u2_n137, u2_u0_u2_n138, u2_u0_u2_n139, u2_u0_u2_n140, u2_u0_u2_n141, u2_u0_u2_n142, 
       u2_u0_u2_n143, u2_u0_u2_n144, u2_u0_u2_n145, u2_u0_u2_n146, u2_u0_u2_n147, u2_u0_u2_n148, u2_u0_u2_n149, u2_u0_u2_n150, u2_u0_u2_n151, 
       u2_u0_u2_n152, u2_u0_u2_n153, u2_u0_u2_n154, u2_u0_u2_n155, u2_u0_u2_n156, u2_u0_u2_n157, u2_u0_u2_n158, u2_u0_u2_n159, u2_u0_u2_n160, 
       u2_u0_u2_n161, u2_u0_u2_n162, u2_u0_u2_n163, u2_u0_u2_n164, u2_u0_u2_n165, u2_u0_u2_n166, u2_u0_u2_n167, u2_u0_u2_n168, u2_u0_u2_n169, 
       u2_u0_u2_n170, u2_u0_u2_n171, u2_u0_u2_n172, u2_u0_u2_n173, u2_u0_u2_n174, u2_u0_u2_n175, u2_u0_u2_n176, u2_u0_u2_n177, u2_u0_u2_n178, 
       u2_u0_u2_n179, u2_u0_u2_n180, u2_u0_u2_n181, u2_u0_u2_n182, u2_u0_u2_n183, u2_u0_u2_n184, u2_u0_u2_n185, u2_u0_u2_n186, u2_u0_u2_n187, 
       u2_u0_u2_n188, u2_u0_u2_n95, u2_u0_u2_n96, u2_u0_u2_n97, u2_u0_u2_n98, u2_u0_u2_n99, u2_u0_u3_n100, u2_u0_u3_n101, u2_u0_u3_n102, 
       u2_u0_u3_n103, u2_u0_u3_n104, u2_u0_u3_n105, u2_u0_u3_n106, u2_u0_u3_n107, u2_u0_u3_n108, u2_u0_u3_n109, u2_u0_u3_n110, u2_u0_u3_n111, 
       u2_u0_u3_n112, u2_u0_u3_n113, u2_u0_u3_n114, u2_u0_u3_n115, u2_u0_u3_n116, u2_u0_u3_n117, u2_u0_u3_n118, u2_u0_u3_n119, u2_u0_u3_n120, 
       u2_u0_u3_n121, u2_u0_u3_n122, u2_u0_u3_n123, u2_u0_u3_n124, u2_u0_u3_n125, u2_u0_u3_n126, u2_u0_u3_n127, u2_u0_u3_n128, u2_u0_u3_n129, 
       u2_u0_u3_n130, u2_u0_u3_n131, u2_u0_u3_n132, u2_u0_u3_n133, u2_u0_u3_n134, u2_u0_u3_n135, u2_u0_u3_n136, u2_u0_u3_n137, u2_u0_u3_n138, 
       u2_u0_u3_n139, u2_u0_u3_n140, u2_u0_u3_n141, u2_u0_u3_n142, u2_u0_u3_n143, u2_u0_u3_n144, u2_u0_u3_n145, u2_u0_u3_n146, u2_u0_u3_n147, 
       u2_u0_u3_n148, u2_u0_u3_n149, u2_u0_u3_n150, u2_u0_u3_n151, u2_u0_u3_n152, u2_u0_u3_n153, u2_u0_u3_n154, u2_u0_u3_n155, u2_u0_u3_n156, 
       u2_u0_u3_n157, u2_u0_u3_n158, u2_u0_u3_n159, u2_u0_u3_n160, u2_u0_u3_n161, u2_u0_u3_n162, u2_u0_u3_n163, u2_u0_u3_n164, u2_u0_u3_n165, 
       u2_u0_u3_n166, u2_u0_u3_n167, u2_u0_u3_n168, u2_u0_u3_n169, u2_u0_u3_n170, u2_u0_u3_n171, u2_u0_u3_n172, u2_u0_u3_n173, u2_u0_u3_n174, 
       u2_u0_u3_n175, u2_u0_u3_n176, u2_u0_u3_n177, u2_u0_u3_n178, u2_u0_u3_n179, u2_u0_u3_n180, u2_u0_u3_n181, u2_u0_u3_n182, u2_u0_u3_n183, 
       u2_u0_u3_n184, u2_u0_u3_n185, u2_u0_u3_n186, u2_u0_u3_n94, u2_u0_u3_n95, u2_u0_u3_n96, u2_u0_u3_n97, u2_u0_u3_n98, u2_u0_u3_n99, 
       u2_u11_X_1, u2_u11_X_10, u2_u11_X_11, u2_u11_X_12, u2_u11_X_13, u2_u11_X_14, u2_u11_X_15, u2_u11_X_16, u2_u11_X_17, 
       u2_u11_X_18, u2_u11_X_2, u2_u11_X_3, u2_u11_X_4, u2_u11_X_5, u2_u11_X_6, u2_u11_X_7, u2_u11_X_8, u2_u11_X_9, 
       u2_u11_u0_n100, u2_u11_u0_n101, u2_u11_u0_n102, u2_u11_u0_n103, u2_u11_u0_n104, u2_u11_u0_n105, u2_u11_u0_n106, u2_u11_u0_n107, u2_u11_u0_n108, 
       u2_u11_u0_n109, u2_u11_u0_n110, u2_u11_u0_n111, u2_u11_u0_n112, u2_u11_u0_n113, u2_u11_u0_n114, u2_u11_u0_n115, u2_u11_u0_n116, u2_u11_u0_n117, 
       u2_u11_u0_n118, u2_u11_u0_n119, u2_u11_u0_n120, u2_u11_u0_n121, u2_u11_u0_n122, u2_u11_u0_n123, u2_u11_u0_n124, u2_u11_u0_n125, u2_u11_u0_n126, 
       u2_u11_u0_n127, u2_u11_u0_n128, u2_u11_u0_n129, u2_u11_u0_n130, u2_u11_u0_n131, u2_u11_u0_n132, u2_u11_u0_n133, u2_u11_u0_n134, u2_u11_u0_n135, 
       u2_u11_u0_n136, u2_u11_u0_n137, u2_u11_u0_n138, u2_u11_u0_n139, u2_u11_u0_n140, u2_u11_u0_n141, u2_u11_u0_n142, u2_u11_u0_n143, u2_u11_u0_n144, 
       u2_u11_u0_n145, u2_u11_u0_n146, u2_u11_u0_n147, u2_u11_u0_n148, u2_u11_u0_n149, u2_u11_u0_n150, u2_u11_u0_n151, u2_u11_u0_n152, u2_u11_u0_n153, 
       u2_u11_u0_n154, u2_u11_u0_n155, u2_u11_u0_n156, u2_u11_u0_n157, u2_u11_u0_n158, u2_u11_u0_n159, u2_u11_u0_n160, u2_u11_u0_n161, u2_u11_u0_n162, 
       u2_u11_u0_n163, u2_u11_u0_n164, u2_u11_u0_n165, u2_u11_u0_n166, u2_u11_u0_n167, u2_u11_u0_n168, u2_u11_u0_n169, u2_u11_u0_n170, u2_u11_u0_n171, 
       u2_u11_u0_n172, u2_u11_u0_n173, u2_u11_u0_n174, u2_u11_u0_n88, u2_u11_u0_n89, u2_u11_u0_n90, u2_u11_u0_n91, u2_u11_u0_n92, u2_u11_u0_n93, 
       u2_u11_u0_n94, u2_u11_u0_n95, u2_u11_u0_n96, u2_u11_u0_n97, u2_u11_u0_n98, u2_u11_u0_n99, u2_u11_u1_n100, u2_u11_u1_n101, u2_u11_u1_n102, 
       u2_u11_u1_n103, u2_u11_u1_n104, u2_u11_u1_n105, u2_u11_u1_n106, u2_u11_u1_n107, u2_u11_u1_n108, u2_u11_u1_n109, u2_u11_u1_n110, u2_u11_u1_n111, 
       u2_u11_u1_n112, u2_u11_u1_n113, u2_u11_u1_n114, u2_u11_u1_n115, u2_u11_u1_n116, u2_u11_u1_n117, u2_u11_u1_n118, u2_u11_u1_n119, u2_u11_u1_n120, 
       u2_u11_u1_n121, u2_u11_u1_n122, u2_u11_u1_n123, u2_u11_u1_n124, u2_u11_u1_n125, u2_u11_u1_n126, u2_u11_u1_n127, u2_u11_u1_n128, u2_u11_u1_n129, 
       u2_u11_u1_n130, u2_u11_u1_n131, u2_u11_u1_n132, u2_u11_u1_n133, u2_u11_u1_n134, u2_u11_u1_n135, u2_u11_u1_n136, u2_u11_u1_n137, u2_u11_u1_n138, 
       u2_u11_u1_n139, u2_u11_u1_n140, u2_u11_u1_n141, u2_u11_u1_n142, u2_u11_u1_n143, u2_u11_u1_n144, u2_u11_u1_n145, u2_u11_u1_n146, u2_u11_u1_n147, 
       u2_u11_u1_n148, u2_u11_u1_n149, u2_u11_u1_n150, u2_u11_u1_n151, u2_u11_u1_n152, u2_u11_u1_n153, u2_u11_u1_n154, u2_u11_u1_n155, u2_u11_u1_n156, 
       u2_u11_u1_n157, u2_u11_u1_n158, u2_u11_u1_n159, u2_u11_u1_n160, u2_u11_u1_n161, u2_u11_u1_n162, u2_u11_u1_n163, u2_u11_u1_n164, u2_u11_u1_n165, 
       u2_u11_u1_n166, u2_u11_u1_n167, u2_u11_u1_n168, u2_u11_u1_n169, u2_u11_u1_n170, u2_u11_u1_n171, u2_u11_u1_n172, u2_u11_u1_n173, u2_u11_u1_n174, 
       u2_u11_u1_n175, u2_u11_u1_n176, u2_u11_u1_n177, u2_u11_u1_n178, u2_u11_u1_n179, u2_u11_u1_n180, u2_u11_u1_n181, u2_u11_u1_n182, u2_u11_u1_n183, 
       u2_u11_u1_n184, u2_u11_u1_n185, u2_u11_u1_n186, u2_u11_u1_n187, u2_u11_u1_n188, u2_u11_u1_n95, u2_u11_u1_n96, u2_u11_u1_n97, u2_u11_u1_n98, 
       u2_u11_u1_n99, u2_u11_u2_n100, u2_u11_u2_n101, u2_u11_u2_n102, u2_u11_u2_n103, u2_u11_u2_n104, u2_u11_u2_n105, u2_u11_u2_n106, u2_u11_u2_n107, 
       u2_u11_u2_n108, u2_u11_u2_n109, u2_u11_u2_n110, u2_u11_u2_n111, u2_u11_u2_n112, u2_u11_u2_n113, u2_u11_u2_n114, u2_u11_u2_n115, u2_u11_u2_n116, 
       u2_u11_u2_n117, u2_u11_u2_n118, u2_u11_u2_n119, u2_u11_u2_n120, u2_u11_u2_n121, u2_u11_u2_n122, u2_u11_u2_n123, u2_u11_u2_n124, u2_u11_u2_n125, 
       u2_u11_u2_n126, u2_u11_u2_n127, u2_u11_u2_n128, u2_u11_u2_n129, u2_u11_u2_n130, u2_u11_u2_n131, u2_u11_u2_n132, u2_u11_u2_n133, u2_u11_u2_n134, 
       u2_u11_u2_n135, u2_u11_u2_n136, u2_u11_u2_n137, u2_u11_u2_n138, u2_u11_u2_n139, u2_u11_u2_n140, u2_u11_u2_n141, u2_u11_u2_n142, u2_u11_u2_n143, 
       u2_u11_u2_n144, u2_u11_u2_n145, u2_u11_u2_n146, u2_u11_u2_n147, u2_u11_u2_n148, u2_u11_u2_n149, u2_u11_u2_n150, u2_u11_u2_n151, u2_u11_u2_n152, 
       u2_u11_u2_n153, u2_u11_u2_n154, u2_u11_u2_n155, u2_u11_u2_n156, u2_u11_u2_n157, u2_u11_u2_n158, u2_u11_u2_n159, u2_u11_u2_n160, u2_u11_u2_n161, 
       u2_u11_u2_n162, u2_u11_u2_n163, u2_u11_u2_n164, u2_u11_u2_n165, u2_u11_u2_n166, u2_u11_u2_n167, u2_u11_u2_n168, u2_u11_u2_n169, u2_u11_u2_n170, 
       u2_u11_u2_n171, u2_u11_u2_n172, u2_u11_u2_n173, u2_u11_u2_n174, u2_u11_u2_n175, u2_u11_u2_n176, u2_u11_u2_n177, u2_u11_u2_n178, u2_u11_u2_n179, 
       u2_u11_u2_n180, u2_u11_u2_n181, u2_u11_u2_n182, u2_u11_u2_n183, u2_u11_u2_n184, u2_u11_u2_n185, u2_u11_u2_n186, u2_u11_u2_n187, u2_u11_u2_n188, 
       u2_u11_u2_n95, u2_u11_u2_n96, u2_u11_u2_n97, u2_u11_u2_n98, u2_u11_u2_n99, u2_u13_X_25, u2_u13_X_26, u2_u13_X_27, u2_u13_X_28, 
       u2_u13_X_29, u2_u13_X_30, u2_u13_X_31, u2_u13_X_32, u2_u13_X_33, u2_u13_X_34, u2_u13_X_35, u2_u13_X_36, u2_u13_u4_n100, 
       u2_u13_u4_n101, u2_u13_u4_n102, u2_u13_u4_n103, u2_u13_u4_n104, u2_u13_u4_n105, u2_u13_u4_n106, u2_u13_u4_n107, u2_u13_u4_n108, u2_u13_u4_n109, 
       u2_u13_u4_n110, u2_u13_u4_n111, u2_u13_u4_n112, u2_u13_u4_n113, u2_u13_u4_n114, u2_u13_u4_n115, u2_u13_u4_n116, u2_u13_u4_n117, u2_u13_u4_n118, 
       u2_u13_u4_n119, u2_u13_u4_n120, u2_u13_u4_n121, u2_u13_u4_n122, u2_u13_u4_n123, u2_u13_u4_n124, u2_u13_u4_n125, u2_u13_u4_n126, u2_u13_u4_n127, 
       u2_u13_u4_n128, u2_u13_u4_n129, u2_u13_u4_n130, u2_u13_u4_n131, u2_u13_u4_n132, u2_u13_u4_n133, u2_u13_u4_n134, u2_u13_u4_n135, u2_u13_u4_n136, 
       u2_u13_u4_n137, u2_u13_u4_n138, u2_u13_u4_n139, u2_u13_u4_n140, u2_u13_u4_n141, u2_u13_u4_n142, u2_u13_u4_n143, u2_u13_u4_n144, u2_u13_u4_n145, 
       u2_u13_u4_n146, u2_u13_u4_n147, u2_u13_u4_n148, u2_u13_u4_n149, u2_u13_u4_n150, u2_u13_u4_n151, u2_u13_u4_n152, u2_u13_u4_n153, u2_u13_u4_n154, 
       u2_u13_u4_n155, u2_u13_u4_n156, u2_u13_u4_n157, u2_u13_u4_n158, u2_u13_u4_n159, u2_u13_u4_n160, u2_u13_u4_n161, u2_u13_u4_n162, u2_u13_u4_n163, 
       u2_u13_u4_n164, u2_u13_u4_n165, u2_u13_u4_n166, u2_u13_u4_n167, u2_u13_u4_n168, u2_u13_u4_n169, u2_u13_u4_n170, u2_u13_u4_n171, u2_u13_u4_n172, 
       u2_u13_u4_n173, u2_u13_u4_n174, u2_u13_u4_n175, u2_u13_u4_n176, u2_u13_u4_n177, u2_u13_u4_n178, u2_u13_u4_n179, u2_u13_u4_n180, u2_u13_u4_n181, 
       u2_u13_u4_n182, u2_u13_u4_n183, u2_u13_u4_n184, u2_u13_u4_n185, u2_u13_u4_n186, u2_u13_u4_n94, u2_u13_u4_n95, u2_u13_u4_n96, u2_u13_u4_n97, 
       u2_u13_u4_n98, u2_u13_u4_n99, u2_u13_u5_n100, u2_u13_u5_n101, u2_u13_u5_n102, u2_u13_u5_n103, u2_u13_u5_n104, u2_u13_u5_n105, u2_u13_u5_n106, 
       u2_u13_u5_n107, u2_u13_u5_n108, u2_u13_u5_n109, u2_u13_u5_n110, u2_u13_u5_n111, u2_u13_u5_n112, u2_u13_u5_n113, u2_u13_u5_n114, u2_u13_u5_n115, 
       u2_u13_u5_n116, u2_u13_u5_n117, u2_u13_u5_n118, u2_u13_u5_n119, u2_u13_u5_n120, u2_u13_u5_n121, u2_u13_u5_n122, u2_u13_u5_n123, u2_u13_u5_n124, 
       u2_u13_u5_n125, u2_u13_u5_n126, u2_u13_u5_n127, u2_u13_u5_n128, u2_u13_u5_n129, u2_u13_u5_n130, u2_u13_u5_n131, u2_u13_u5_n132, u2_u13_u5_n133, 
       u2_u13_u5_n134, u2_u13_u5_n135, u2_u13_u5_n136, u2_u13_u5_n137, u2_u13_u5_n138, u2_u13_u5_n139, u2_u13_u5_n140, u2_u13_u5_n141, u2_u13_u5_n142, 
       u2_u13_u5_n143, u2_u13_u5_n144, u2_u13_u5_n145, u2_u13_u5_n146, u2_u13_u5_n147, u2_u13_u5_n148, u2_u13_u5_n149, u2_u13_u5_n150, u2_u13_u5_n151, 
       u2_u13_u5_n152, u2_u13_u5_n153, u2_u13_u5_n154, u2_u13_u5_n155, u2_u13_u5_n156, u2_u13_u5_n157, u2_u13_u5_n158, u2_u13_u5_n159, u2_u13_u5_n160, 
       u2_u13_u5_n161, u2_u13_u5_n162, u2_u13_u5_n163, u2_u13_u5_n164, u2_u13_u5_n165, u2_u13_u5_n166, u2_u13_u5_n167, u2_u13_u5_n168, u2_u13_u5_n169, 
       u2_u13_u5_n170, u2_u13_u5_n171, u2_u13_u5_n172, u2_u13_u5_n173, u2_u13_u5_n174, u2_u13_u5_n175, u2_u13_u5_n176, u2_u13_u5_n177, u2_u13_u5_n178, 
       u2_u13_u5_n179, u2_u13_u5_n180, u2_u13_u5_n181, u2_u13_u5_n182, u2_u13_u5_n183, u2_u13_u5_n184, u2_u13_u5_n185, u2_u13_u5_n186, u2_u13_u5_n187, 
       u2_u13_u5_n188, u2_u13_u5_n189, u2_u13_u5_n190, u2_u13_u5_n191, u2_u13_u5_n192, u2_u13_u5_n193, u2_u13_u5_n194, u2_u13_u5_n195, u2_u13_u5_n196, 
       u2_u13_u5_n99, u2_u14_X_1, u2_u14_X_10, u2_u14_X_11, u2_u14_X_12, u2_u14_X_2, u2_u14_X_25, u2_u14_X_26, u2_u14_X_27, 
       u2_u14_X_28, u2_u14_X_29, u2_u14_X_3, u2_u14_X_30, u2_u14_X_31, u2_u14_X_32, u2_u14_X_33, u2_u14_X_34, u2_u14_X_35, 
       u2_u14_X_36, u2_u14_X_37, u2_u14_X_38, u2_u14_X_39, u2_u14_X_4, u2_u14_X_40, u2_u14_X_41, u2_u14_X_42, u2_u14_X_5, 
       u2_u14_X_6, u2_u14_X_7, u2_u14_X_8, u2_u14_X_9, u2_u14_u0_n100, u2_u14_u0_n101, u2_u14_u0_n102, u2_u14_u0_n103, u2_u14_u0_n104, 
       u2_u14_u0_n105, u2_u14_u0_n106, u2_u14_u0_n107, u2_u14_u0_n108, u2_u14_u0_n109, u2_u14_u0_n110, u2_u14_u0_n111, u2_u14_u0_n112, u2_u14_u0_n113, 
       u2_u14_u0_n114, u2_u14_u0_n115, u2_u14_u0_n116, u2_u14_u0_n117, u2_u14_u0_n118, u2_u14_u0_n119, u2_u14_u0_n120, u2_u14_u0_n121, u2_u14_u0_n122, 
       u2_u14_u0_n123, u2_u14_u0_n124, u2_u14_u0_n125, u2_u14_u0_n126, u2_u14_u0_n127, u2_u14_u0_n128, u2_u14_u0_n129, u2_u14_u0_n130, u2_u14_u0_n131, 
       u2_u14_u0_n132, u2_u14_u0_n133, u2_u14_u0_n134, u2_u14_u0_n135, u2_u14_u0_n136, u2_u14_u0_n137, u2_u14_u0_n138, u2_u14_u0_n139, u2_u14_u0_n140, 
       u2_u14_u0_n141, u2_u14_u0_n142, u2_u14_u0_n143, u2_u14_u0_n144, u2_u14_u0_n145, u2_u14_u0_n146, u2_u14_u0_n147, u2_u14_u0_n148, u2_u14_u0_n149, 
       u2_u14_u0_n150, u2_u14_u0_n151, u2_u14_u0_n152, u2_u14_u0_n153, u2_u14_u0_n154, u2_u14_u0_n155, u2_u14_u0_n156, u2_u14_u0_n157, u2_u14_u0_n158, 
       u2_u14_u0_n159, u2_u14_u0_n160, u2_u14_u0_n161, u2_u14_u0_n162, u2_u14_u0_n163, u2_u14_u0_n164, u2_u14_u0_n165, u2_u14_u0_n166, u2_u14_u0_n167, 
       u2_u14_u0_n168, u2_u14_u0_n169, u2_u14_u0_n170, u2_u14_u0_n171, u2_u14_u0_n172, u2_u14_u0_n173, u2_u14_u0_n174, u2_u14_u0_n88, u2_u14_u0_n89, 
       u2_u14_u0_n90, u2_u14_u0_n91, u2_u14_u0_n92, u2_u14_u0_n93, u2_u14_u0_n94, u2_u14_u0_n95, u2_u14_u0_n96, u2_u14_u0_n97, u2_u14_u0_n98, 
       u2_u14_u0_n99, u2_u14_u1_n100, u2_u14_u1_n101, u2_u14_u1_n102, u2_u14_u1_n103, u2_u14_u1_n104, u2_u14_u1_n105, u2_u14_u1_n106, u2_u14_u1_n107, 
       u2_u14_u1_n108, u2_u14_u1_n109, u2_u14_u1_n110, u2_u14_u1_n111, u2_u14_u1_n112, u2_u14_u1_n113, u2_u14_u1_n114, u2_u14_u1_n115, u2_u14_u1_n116, 
       u2_u14_u1_n117, u2_u14_u1_n118, u2_u14_u1_n119, u2_u14_u1_n120, u2_u14_u1_n121, u2_u14_u1_n122, u2_u14_u1_n123, u2_u14_u1_n124, u2_u14_u1_n125, 
       u2_u14_u1_n126, u2_u14_u1_n127, u2_u14_u1_n128, u2_u14_u1_n129, u2_u14_u1_n130, u2_u14_u1_n131, u2_u14_u1_n132, u2_u14_u1_n133, u2_u14_u1_n134, 
       u2_u14_u1_n135, u2_u14_u1_n136, u2_u14_u1_n137, u2_u14_u1_n138, u2_u14_u1_n139, u2_u14_u1_n140, u2_u14_u1_n141, u2_u14_u1_n142, u2_u14_u1_n143, 
       u2_u14_u1_n144, u2_u14_u1_n145, u2_u14_u1_n146, u2_u14_u1_n147, u2_u14_u1_n148, u2_u14_u1_n149, u2_u14_u1_n150, u2_u14_u1_n151, u2_u14_u1_n152, 
       u2_u14_u1_n153, u2_u14_u1_n154, u2_u14_u1_n155, u2_u14_u1_n156, u2_u14_u1_n157, u2_u14_u1_n158, u2_u14_u1_n159, u2_u14_u1_n160, u2_u14_u1_n161, 
       u2_u14_u1_n162, u2_u14_u1_n163, u2_u14_u1_n164, u2_u14_u1_n165, u2_u14_u1_n166, u2_u14_u1_n167, u2_u14_u1_n168, u2_u14_u1_n169, u2_u14_u1_n170, 
       u2_u14_u1_n171, u2_u14_u1_n172, u2_u14_u1_n173, u2_u14_u1_n174, u2_u14_u1_n175, u2_u14_u1_n176, u2_u14_u1_n177, u2_u14_u1_n178, u2_u14_u1_n179, 
       u2_u14_u1_n180, u2_u14_u1_n181, u2_u14_u1_n182, u2_u14_u1_n183, u2_u14_u1_n184, u2_u14_u1_n185, u2_u14_u1_n186, u2_u14_u1_n187, u2_u14_u1_n188, 
       u2_u14_u1_n95, u2_u14_u1_n96, u2_u14_u1_n97, u2_u14_u1_n98, u2_u14_u1_n99, u2_u14_u4_n100, u2_u14_u4_n101, u2_u14_u4_n102, u2_u14_u4_n103, 
       u2_u14_u4_n104, u2_u14_u4_n105, u2_u14_u4_n106, u2_u14_u4_n107, u2_u14_u4_n108, u2_u14_u4_n109, u2_u14_u4_n110, u2_u14_u4_n111, u2_u14_u4_n112, 
       u2_u14_u4_n113, u2_u14_u4_n114, u2_u14_u4_n115, u2_u14_u4_n116, u2_u14_u4_n117, u2_u14_u4_n118, u2_u14_u4_n119, u2_u14_u4_n120, u2_u14_u4_n121, 
       u2_u14_u4_n122, u2_u14_u4_n123, u2_u14_u4_n124, u2_u14_u4_n125, u2_u14_u4_n126, u2_u14_u4_n127, u2_u14_u4_n128, u2_u14_u4_n129, u2_u14_u4_n130, 
       u2_u14_u4_n131, u2_u14_u4_n132, u2_u14_u4_n133, u2_u14_u4_n134, u2_u14_u4_n135, u2_u14_u4_n136, u2_u14_u4_n137, u2_u14_u4_n138, u2_u14_u4_n139, 
       u2_u14_u4_n140, u2_u14_u4_n141, u2_u14_u4_n142, u2_u14_u4_n143, u2_u14_u4_n144, u2_u14_u4_n145, u2_u14_u4_n146, u2_u14_u4_n147, u2_u14_u4_n148, 
       u2_u14_u4_n149, u2_u14_u4_n150, u2_u14_u4_n151, u2_u14_u4_n152, u2_u14_u4_n153, u2_u14_u4_n154, u2_u14_u4_n155, u2_u14_u4_n156, u2_u14_u4_n157, 
       u2_u14_u4_n158, u2_u14_u4_n159, u2_u14_u4_n160, u2_u14_u4_n161, u2_u14_u4_n162, u2_u14_u4_n163, u2_u14_u4_n164, u2_u14_u4_n165, u2_u14_u4_n166, 
       u2_u14_u4_n167, u2_u14_u4_n168, u2_u14_u4_n169, u2_u14_u4_n170, u2_u14_u4_n171, u2_u14_u4_n172, u2_u14_u4_n173, u2_u14_u4_n174, u2_u14_u4_n175, 
       u2_u14_u4_n176, u2_u14_u4_n177, u2_u14_u4_n178, u2_u14_u4_n179, u2_u14_u4_n180, u2_u14_u4_n181, u2_u14_u4_n182, u2_u14_u4_n183, u2_u14_u4_n184, 
       u2_u14_u4_n185, u2_u14_u4_n186, u2_u14_u4_n94, u2_u14_u4_n95, u2_u14_u4_n96, u2_u14_u4_n97, u2_u14_u4_n98, u2_u14_u4_n99, u2_u14_u5_n100, 
       u2_u14_u5_n101, u2_u14_u5_n102, u2_u14_u5_n103, u2_u14_u5_n104, u2_u14_u5_n105, u2_u14_u5_n106, u2_u14_u5_n107, u2_u14_u5_n108, u2_u14_u5_n109, 
       u2_u14_u5_n110, u2_u14_u5_n111, u2_u14_u5_n112, u2_u14_u5_n113, u2_u14_u5_n114, u2_u14_u5_n115, u2_u14_u5_n116, u2_u14_u5_n117, u2_u14_u5_n118, 
       u2_u14_u5_n119, u2_u14_u5_n120, u2_u14_u5_n121, u2_u14_u5_n122, u2_u14_u5_n123, u2_u14_u5_n124, u2_u14_u5_n125, u2_u14_u5_n126, u2_u14_u5_n127, 
       u2_u14_u5_n128, u2_u14_u5_n129, u2_u14_u5_n130, u2_u14_u5_n131, u2_u14_u5_n132, u2_u14_u5_n133, u2_u14_u5_n134, u2_u14_u5_n135, u2_u14_u5_n136, 
       u2_u14_u5_n137, u2_u14_u5_n138, u2_u14_u5_n139, u2_u14_u5_n140, u2_u14_u5_n141, u2_u14_u5_n142, u2_u14_u5_n143, u2_u14_u5_n144, u2_u14_u5_n145, 
       u2_u14_u5_n146, u2_u14_u5_n147, u2_u14_u5_n148, u2_u14_u5_n149, u2_u14_u5_n150, u2_u14_u5_n151, u2_u14_u5_n152, u2_u14_u5_n153, u2_u14_u5_n154, 
       u2_u14_u5_n155, u2_u14_u5_n156, u2_u14_u5_n157, u2_u14_u5_n158, u2_u14_u5_n159, u2_u14_u5_n160, u2_u14_u5_n161, u2_u14_u5_n162, u2_u14_u5_n163, 
       u2_u14_u5_n164, u2_u14_u5_n165, u2_u14_u5_n166, u2_u14_u5_n167, u2_u14_u5_n168, u2_u14_u5_n169, u2_u14_u5_n170, u2_u14_u5_n171, u2_u14_u5_n172, 
       u2_u14_u5_n173, u2_u14_u5_n174, u2_u14_u5_n175, u2_u14_u5_n176, u2_u14_u5_n177, u2_u14_u5_n178, u2_u14_u5_n179, u2_u14_u5_n180, u2_u14_u5_n181, 
       u2_u14_u5_n182, u2_u14_u5_n183, u2_u14_u5_n184, u2_u14_u5_n185, u2_u14_u5_n186, u2_u14_u5_n187, u2_u14_u5_n188, u2_u14_u5_n189, u2_u14_u5_n190, 
       u2_u14_u5_n191, u2_u14_u5_n192, u2_u14_u5_n193, u2_u14_u5_n194, u2_u14_u5_n195, u2_u14_u5_n196, u2_u14_u5_n99, u2_u14_u6_n100, u2_u14_u6_n101, 
       u2_u14_u6_n102, u2_u14_u6_n103, u2_u14_u6_n104, u2_u14_u6_n105, u2_u14_u6_n106, u2_u14_u6_n107, u2_u14_u6_n108, u2_u14_u6_n109, u2_u14_u6_n110, 
       u2_u14_u6_n111, u2_u14_u6_n112, u2_u14_u6_n113, u2_u14_u6_n114, u2_u14_u6_n115, u2_u14_u6_n116, u2_u14_u6_n117, u2_u14_u6_n118, u2_u14_u6_n119, 
       u2_u14_u6_n120, u2_u14_u6_n121, u2_u14_u6_n122, u2_u14_u6_n123, u2_u14_u6_n124, u2_u14_u6_n125, u2_u14_u6_n126, u2_u14_u6_n127, u2_u14_u6_n128, 
       u2_u14_u6_n129, u2_u14_u6_n130, u2_u14_u6_n131, u2_u14_u6_n132, u2_u14_u6_n133, u2_u14_u6_n134, u2_u14_u6_n135, u2_u14_u6_n136, u2_u14_u6_n137, 
       u2_u14_u6_n138, u2_u14_u6_n139, u2_u14_u6_n140, u2_u14_u6_n141, u2_u14_u6_n142, u2_u14_u6_n143, u2_u14_u6_n144, u2_u14_u6_n145, u2_u14_u6_n146, 
       u2_u14_u6_n147, u2_u14_u6_n148, u2_u14_u6_n149, u2_u14_u6_n150, u2_u14_u6_n151, u2_u14_u6_n152, u2_u14_u6_n153, u2_u14_u6_n154, u2_u14_u6_n155, 
       u2_u14_u6_n156, u2_u14_u6_n157, u2_u14_u6_n158, u2_u14_u6_n159, u2_u14_u6_n160, u2_u14_u6_n161, u2_u14_u6_n162, u2_u14_u6_n163, u2_u14_u6_n164, 
       u2_u14_u6_n165, u2_u14_u6_n166, u2_u14_u6_n167, u2_u14_u6_n168, u2_u14_u6_n169, u2_u14_u6_n170, u2_u14_u6_n171, u2_u14_u6_n172, u2_u14_u6_n173, 
       u2_u14_u6_n174, u2_u14_u6_n88, u2_u14_u6_n89, u2_u14_u6_n90, u2_u14_u6_n91, u2_u14_u6_n92, u2_u14_u6_n93, u2_u14_u6_n94, u2_u14_u6_n95, 
       u2_u14_u6_n96, u2_u14_u6_n97, u2_u14_u6_n98, u2_u14_u6_n99, u2_u15_X_1, u2_u15_X_2, u2_u15_X_25, u2_u15_X_26, u2_u15_X_27, 
       u2_u15_X_28, u2_u15_X_29, u2_u15_X_3, u2_u15_X_30, u2_u15_X_31, u2_u15_X_32, u2_u15_X_33, u2_u15_X_34, u2_u15_X_35, 
       u2_u15_X_36, u2_u15_X_37, u2_u15_X_38, u2_u15_X_39, u2_u15_X_4, u2_u15_X_40, u2_u15_X_41, u2_u15_X_42, u2_u15_X_43, 
       u2_u15_X_44, u2_u15_X_45, u2_u15_X_46, u2_u15_X_47, u2_u15_X_48, u2_u15_X_5, u2_u15_X_6, u2_u15_u0_n100, u2_u15_u0_n101, 
       u2_u15_u0_n102, u2_u15_u0_n103, u2_u15_u0_n104, u2_u15_u0_n105, u2_u15_u0_n106, u2_u15_u0_n107, u2_u15_u0_n108, u2_u15_u0_n109, u2_u15_u0_n110, 
       u2_u15_u0_n111, u2_u15_u0_n112, u2_u15_u0_n113, u2_u15_u0_n114, u2_u15_u0_n115, u2_u15_u0_n116, u2_u15_u0_n117, u2_u15_u0_n118, u2_u15_u0_n119, 
       u2_u15_u0_n120, u2_u15_u0_n121, u2_u15_u0_n122, u2_u15_u0_n123, u2_u15_u0_n124, u2_u15_u0_n125, u2_u15_u0_n126, u2_u15_u0_n127, u2_u15_u0_n128, 
       u2_u15_u0_n129, u2_u15_u0_n130, u2_u15_u0_n131, u2_u15_u0_n132, u2_u15_u0_n133, u2_u15_u0_n134, u2_u15_u0_n135, u2_u15_u0_n136, u2_u15_u0_n137, 
       u2_u15_u0_n138, u2_u15_u0_n139, u2_u15_u0_n140, u2_u15_u0_n141, u2_u15_u0_n142, u2_u15_u0_n143, u2_u15_u0_n144, u2_u15_u0_n145, u2_u15_u0_n146, 
       u2_u15_u0_n147, u2_u15_u0_n148, u2_u15_u0_n149, u2_u15_u0_n150, u2_u15_u0_n151, u2_u15_u0_n152, u2_u15_u0_n153, u2_u15_u0_n154, u2_u15_u0_n155, 
       u2_u15_u0_n156, u2_u15_u0_n157, u2_u15_u0_n158, u2_u15_u0_n159, u2_u15_u0_n160, u2_u15_u0_n161, u2_u15_u0_n162, u2_u15_u0_n163, u2_u15_u0_n164, 
       u2_u15_u0_n165, u2_u15_u0_n166, u2_u15_u0_n167, u2_u15_u0_n168, u2_u15_u0_n169, u2_u15_u0_n170, u2_u15_u0_n171, u2_u15_u0_n172, u2_u15_u0_n173, 
       u2_u15_u0_n174, u2_u15_u0_n88, u2_u15_u0_n89, u2_u15_u0_n90, u2_u15_u0_n91, u2_u15_u0_n92, u2_u15_u0_n93, u2_u15_u0_n94, u2_u15_u0_n95, 
       u2_u15_u0_n96, u2_u15_u0_n97, u2_u15_u0_n98, u2_u15_u0_n99, u2_u15_u4_n100, u2_u15_u4_n101, u2_u15_u4_n102, u2_u15_u4_n103, u2_u15_u4_n104, 
       u2_u15_u4_n105, u2_u15_u4_n106, u2_u15_u4_n107, u2_u15_u4_n108, u2_u15_u4_n109, u2_u15_u4_n110, u2_u15_u4_n111, u2_u15_u4_n112, u2_u15_u4_n113, 
       u2_u15_u4_n114, u2_u15_u4_n115, u2_u15_u4_n116, u2_u15_u4_n117, u2_u15_u4_n118, u2_u15_u4_n119, u2_u15_u4_n120, u2_u15_u4_n121, u2_u15_u4_n122, 
       u2_u15_u4_n123, u2_u15_u4_n124, u2_u15_u4_n125, u2_u15_u4_n126, u2_u15_u4_n127, u2_u15_u4_n128, u2_u15_u4_n129, u2_u15_u4_n130, u2_u15_u4_n131, 
       u2_u15_u4_n132, u2_u15_u4_n133, u2_u15_u4_n134, u2_u15_u4_n135, u2_u15_u4_n136, u2_u15_u4_n137, u2_u15_u4_n138, u2_u15_u4_n139, u2_u15_u4_n140, 
       u2_u15_u4_n141, u2_u15_u4_n142, u2_u15_u4_n143, u2_u15_u4_n144, u2_u15_u4_n145, u2_u15_u4_n146, u2_u15_u4_n147, u2_u15_u4_n148, u2_u15_u4_n149, 
       u2_u15_u4_n150, u2_u15_u4_n151, u2_u15_u4_n152, u2_u15_u4_n153, u2_u15_u4_n154, u2_u15_u4_n155, u2_u15_u4_n156, u2_u15_u4_n157, u2_u15_u4_n158, 
       u2_u15_u4_n159, u2_u15_u4_n160, u2_u15_u4_n161, u2_u15_u4_n162, u2_u15_u4_n163, u2_u15_u4_n164, u2_u15_u4_n165, u2_u15_u4_n166, u2_u15_u4_n167, 
       u2_u15_u4_n168, u2_u15_u4_n169, u2_u15_u4_n170, u2_u15_u4_n171, u2_u15_u4_n172, u2_u15_u4_n173, u2_u15_u4_n174, u2_u15_u4_n175, u2_u15_u4_n176, 
       u2_u15_u4_n177, u2_u15_u4_n178, u2_u15_u4_n179, u2_u15_u4_n180, u2_u15_u4_n181, u2_u15_u4_n182, u2_u15_u4_n183, u2_u15_u4_n184, u2_u15_u4_n185, 
       u2_u15_u4_n186, u2_u15_u4_n94, u2_u15_u4_n95, u2_u15_u4_n96, u2_u15_u4_n97, u2_u15_u4_n98, u2_u15_u4_n99, u2_u15_u5_n100, u2_u15_u5_n101, 
       u2_u15_u5_n102, u2_u15_u5_n103, u2_u15_u5_n104, u2_u15_u5_n105, u2_u15_u5_n106, u2_u15_u5_n107, u2_u15_u5_n108, u2_u15_u5_n109, u2_u15_u5_n110, 
       u2_u15_u5_n111, u2_u15_u5_n112, u2_u15_u5_n113, u2_u15_u5_n114, u2_u15_u5_n115, u2_u15_u5_n116, u2_u15_u5_n117, u2_u15_u5_n118, u2_u15_u5_n119, 
       u2_u15_u5_n120, u2_u15_u5_n121, u2_u15_u5_n122, u2_u15_u5_n123, u2_u15_u5_n124, u2_u15_u5_n125, u2_u15_u5_n126, u2_u15_u5_n127, u2_u15_u5_n128, 
       u2_u15_u5_n129, u2_u15_u5_n130, u2_u15_u5_n131, u2_u15_u5_n132, u2_u15_u5_n133, u2_u15_u5_n134, u2_u15_u5_n135, u2_u15_u5_n136, u2_u15_u5_n137, 
       u2_u15_u5_n138, u2_u15_u5_n139, u2_u15_u5_n140, u2_u15_u5_n141, u2_u15_u5_n142, u2_u15_u5_n143, u2_u15_u5_n144, u2_u15_u5_n145, u2_u15_u5_n146, 
       u2_u15_u5_n147, u2_u15_u5_n148, u2_u15_u5_n149, u2_u15_u5_n150, u2_u15_u5_n151, u2_u15_u5_n152, u2_u15_u5_n153, u2_u15_u5_n154, u2_u15_u5_n155, 
       u2_u15_u5_n156, u2_u15_u5_n157, u2_u15_u5_n158, u2_u15_u5_n159, u2_u15_u5_n160, u2_u15_u5_n161, u2_u15_u5_n162, u2_u15_u5_n163, u2_u15_u5_n164, 
       u2_u15_u5_n165, u2_u15_u5_n166, u2_u15_u5_n167, u2_u15_u5_n168, u2_u15_u5_n169, u2_u15_u5_n170, u2_u15_u5_n171, u2_u15_u5_n172, u2_u15_u5_n173, 
       u2_u15_u5_n174, u2_u15_u5_n175, u2_u15_u5_n176, u2_u15_u5_n177, u2_u15_u5_n178, u2_u15_u5_n179, u2_u15_u5_n180, u2_u15_u5_n181, u2_u15_u5_n182, 
       u2_u15_u5_n183, u2_u15_u5_n184, u2_u15_u5_n185, u2_u15_u5_n186, u2_u15_u5_n187, u2_u15_u5_n188, u2_u15_u5_n189, u2_u15_u5_n190, u2_u15_u5_n191, 
       u2_u15_u5_n192, u2_u15_u5_n193, u2_u15_u5_n194, u2_u15_u5_n195, u2_u15_u5_n196, u2_u15_u5_n99, u2_u15_u6_n100, u2_u15_u6_n101, u2_u15_u6_n102, 
       u2_u15_u6_n103, u2_u15_u6_n104, u2_u15_u6_n105, u2_u15_u6_n106, u2_u15_u6_n107, u2_u15_u6_n108, u2_u15_u6_n109, u2_u15_u6_n110, u2_u15_u6_n111, 
       u2_u15_u6_n112, u2_u15_u6_n113, u2_u15_u6_n114, u2_u15_u6_n115, u2_u15_u6_n116, u2_u15_u6_n117, u2_u15_u6_n118, u2_u15_u6_n119, u2_u15_u6_n120, 
       u2_u15_u6_n121, u2_u15_u6_n122, u2_u15_u6_n123, u2_u15_u6_n124, u2_u15_u6_n125, u2_u15_u6_n126, u2_u15_u6_n127, u2_u15_u6_n128, u2_u15_u6_n129, 
       u2_u15_u6_n130, u2_u15_u6_n131, u2_u15_u6_n132, u2_u15_u6_n133, u2_u15_u6_n134, u2_u15_u6_n135, u2_u15_u6_n136, u2_u15_u6_n137, u2_u15_u6_n138, 
       u2_u15_u6_n139, u2_u15_u6_n140, u2_u15_u6_n141, u2_u15_u6_n142, u2_u15_u6_n143, u2_u15_u6_n144, u2_u15_u6_n145, u2_u15_u6_n146, u2_u15_u6_n147, 
       u2_u15_u6_n148, u2_u15_u6_n149, u2_u15_u6_n150, u2_u15_u6_n151, u2_u15_u6_n152, u2_u15_u6_n153, u2_u15_u6_n154, u2_u15_u6_n155, u2_u15_u6_n156, 
       u2_u15_u6_n157, u2_u15_u6_n158, u2_u15_u6_n159, u2_u15_u6_n160, u2_u15_u6_n161, u2_u15_u6_n162, u2_u15_u6_n163, u2_u15_u6_n164, u2_u15_u6_n165, 
       u2_u15_u6_n166, u2_u15_u6_n167, u2_u15_u6_n168, u2_u15_u6_n169, u2_u15_u6_n170, u2_u15_u6_n171, u2_u15_u6_n172, u2_u15_u6_n173, u2_u15_u6_n174, 
       u2_u15_u6_n88, u2_u15_u6_n89, u2_u15_u6_n90, u2_u15_u6_n91, u2_u15_u6_n92, u2_u15_u6_n93, u2_u15_u6_n94, u2_u15_u6_n95, u2_u15_u6_n96, 
       u2_u15_u6_n97, u2_u15_u6_n98, u2_u15_u6_n99, u2_u15_u7_n100, u2_u15_u7_n101, u2_u15_u7_n102, u2_u15_u7_n103, u2_u15_u7_n104, u2_u15_u7_n105, 
       u2_u15_u7_n106, u2_u15_u7_n107, u2_u15_u7_n108, u2_u15_u7_n109, u2_u15_u7_n110, u2_u15_u7_n111, u2_u15_u7_n112, u2_u15_u7_n113, u2_u15_u7_n114, 
       u2_u15_u7_n115, u2_u15_u7_n116, u2_u15_u7_n117, u2_u15_u7_n118, u2_u15_u7_n119, u2_u15_u7_n120, u2_u15_u7_n121, u2_u15_u7_n122, u2_u15_u7_n123, 
       u2_u15_u7_n124, u2_u15_u7_n125, u2_u15_u7_n126, u2_u15_u7_n127, u2_u15_u7_n128, u2_u15_u7_n129, u2_u15_u7_n130, u2_u15_u7_n131, u2_u15_u7_n132, 
       u2_u15_u7_n133, u2_u15_u7_n134, u2_u15_u7_n135, u2_u15_u7_n136, u2_u15_u7_n137, u2_u15_u7_n138, u2_u15_u7_n139, u2_u15_u7_n140, u2_u15_u7_n141, 
       u2_u15_u7_n142, u2_u15_u7_n143, u2_u15_u7_n144, u2_u15_u7_n145, u2_u15_u7_n146, u2_u15_u7_n147, u2_u15_u7_n148, u2_u15_u7_n149, u2_u15_u7_n150, 
       u2_u15_u7_n151, u2_u15_u7_n152, u2_u15_u7_n153, u2_u15_u7_n154, u2_u15_u7_n155, u2_u15_u7_n156, u2_u15_u7_n157, u2_u15_u7_n158, u2_u15_u7_n159, 
       u2_u15_u7_n160, u2_u15_u7_n161, u2_u15_u7_n162, u2_u15_u7_n163, u2_u15_u7_n164, u2_u15_u7_n165, u2_u15_u7_n166, u2_u15_u7_n167, u2_u15_u7_n168, 
       u2_u15_u7_n169, u2_u15_u7_n170, u2_u15_u7_n171, u2_u15_u7_n172, u2_u15_u7_n173, u2_u15_u7_n174, u2_u15_u7_n175, u2_u15_u7_n176, u2_u15_u7_n177, 
       u2_u15_u7_n178, u2_u15_u7_n179, u2_u15_u7_n180, u2_u15_u7_n91, u2_u15_u7_n92, u2_u15_u7_n93, u2_u15_u7_n94, u2_u15_u7_n95, u2_u15_u7_n96, 
       u2_u15_u7_n97, u2_u15_u7_n98, u2_u15_u7_n99, u2_u1_X_25, u2_u1_X_26, u2_u1_X_27, u2_u1_X_28, u2_u1_X_29, u2_u1_X_30, 
       u2_u1_X_37, u2_u1_X_38, u2_u1_X_39, u2_u1_X_40, u2_u1_X_41, u2_u1_X_42, u2_u1_u4_n100, u2_u1_u4_n101, u2_u1_u4_n102, 
       u2_u1_u4_n103, u2_u1_u4_n104, u2_u1_u4_n105, u2_u1_u4_n106, u2_u1_u4_n107, u2_u1_u4_n108, u2_u1_u4_n109, u2_u1_u4_n110, u2_u1_u4_n111, 
       u2_u1_u4_n112, u2_u1_u4_n113, u2_u1_u4_n114, u2_u1_u4_n115, u2_u1_u4_n116, u2_u1_u4_n117, u2_u1_u4_n118, u2_u1_u4_n119, u2_u1_u4_n120, 
       u2_u1_u4_n121, u2_u1_u4_n122, u2_u1_u4_n123, u2_u1_u4_n124, u2_u1_u4_n125, u2_u1_u4_n126, u2_u1_u4_n127, u2_u1_u4_n128, u2_u1_u4_n129, 
       u2_u1_u4_n130, u2_u1_u4_n131, u2_u1_u4_n132, u2_u1_u4_n133, u2_u1_u4_n134, u2_u1_u4_n135, u2_u1_u4_n136, u2_u1_u4_n137, u2_u1_u4_n138, 
       u2_u1_u4_n139, u2_u1_u4_n140, u2_u1_u4_n141, u2_u1_u4_n142, u2_u1_u4_n143, u2_u1_u4_n144, u2_u1_u4_n145, u2_u1_u4_n146, u2_u1_u4_n147, 
       u2_u1_u4_n148, u2_u1_u4_n149, u2_u1_u4_n150, u2_u1_u4_n151, u2_u1_u4_n152, u2_u1_u4_n153, u2_u1_u4_n154, u2_u1_u4_n155, u2_u1_u4_n156, 
       u2_u1_u4_n157, u2_u1_u4_n158, u2_u1_u4_n159, u2_u1_u4_n160, u2_u1_u4_n161, u2_u1_u4_n162, u2_u1_u4_n163, u2_u1_u4_n164, u2_u1_u4_n165, 
       u2_u1_u4_n166, u2_u1_u4_n167, u2_u1_u4_n168, u2_u1_u4_n169, u2_u1_u4_n170, u2_u1_u4_n171, u2_u1_u4_n172, u2_u1_u4_n173, u2_u1_u4_n174, 
       u2_u1_u4_n175, u2_u1_u4_n176, u2_u1_u4_n177, u2_u1_u4_n178, u2_u1_u4_n179, u2_u1_u4_n180, u2_u1_u4_n181, u2_u1_u4_n182, u2_u1_u4_n183, 
       u2_u1_u4_n184, u2_u1_u4_n185, u2_u1_u4_n186, u2_u1_u4_n94, u2_u1_u4_n95, u2_u1_u4_n96, u2_u1_u4_n97, u2_u1_u4_n98, u2_u1_u4_n99, 
       u2_u1_u6_n100, u2_u1_u6_n101, u2_u1_u6_n102, u2_u1_u6_n103, u2_u1_u6_n104, u2_u1_u6_n105, u2_u1_u6_n106, u2_u1_u6_n107, u2_u1_u6_n108, 
       u2_u1_u6_n109, u2_u1_u6_n110, u2_u1_u6_n111, u2_u1_u6_n112, u2_u1_u6_n113, u2_u1_u6_n114, u2_u1_u6_n115, u2_u1_u6_n116, u2_u1_u6_n117, 
       u2_u1_u6_n118, u2_u1_u6_n119, u2_u1_u6_n120, u2_u1_u6_n121, u2_u1_u6_n122, u2_u1_u6_n123, u2_u1_u6_n124, u2_u1_u6_n125, u2_u1_u6_n126, 
       u2_u1_u6_n127, u2_u1_u6_n128, u2_u1_u6_n129, u2_u1_u6_n130, u2_u1_u6_n131, u2_u1_u6_n132, u2_u1_u6_n133, u2_u1_u6_n134, u2_u1_u6_n135, 
       u2_u1_u6_n136, u2_u1_u6_n137, u2_u1_u6_n138, u2_u1_u6_n139, u2_u1_u6_n140, u2_u1_u6_n141, u2_u1_u6_n142, u2_u1_u6_n143, u2_u1_u6_n144, 
       u2_u1_u6_n145, u2_u1_u6_n146, u2_u1_u6_n147, u2_u1_u6_n148, u2_u1_u6_n149, u2_u1_u6_n150, u2_u1_u6_n151, u2_u1_u6_n152, u2_u1_u6_n153, 
       u2_u1_u6_n154, u2_u1_u6_n155, u2_u1_u6_n156, u2_u1_u6_n157, u2_u1_u6_n158, u2_u1_u6_n159, u2_u1_u6_n160, u2_u1_u6_n161, u2_u1_u6_n162, 
       u2_u1_u6_n163, u2_u1_u6_n164, u2_u1_u6_n165, u2_u1_u6_n166, u2_u1_u6_n167, u2_u1_u6_n168, u2_u1_u6_n169, u2_u1_u6_n170, u2_u1_u6_n171, 
       u2_u1_u6_n172, u2_u1_u6_n173, u2_u1_u6_n174, u2_u1_u6_n88, u2_u1_u6_n89, u2_u1_u6_n90, u2_u1_u6_n91, u2_u1_u6_n92, u2_u1_u6_n93, 
       u2_u1_u6_n94, u2_u1_u6_n95, u2_u1_u6_n96, u2_u1_u6_n97, u2_u1_u6_n98, u2_u1_u6_n99, u2_u2_X_1, u2_u2_X_10, u2_u2_X_11, 
       u2_u2_X_12, u2_u2_X_13, u2_u2_X_14, u2_u2_X_15, u2_u2_X_16, u2_u2_X_17, u2_u2_X_18, u2_u2_X_19, u2_u2_X_2, 
       u2_u2_X_20, u2_u2_X_21, u2_u2_X_22, u2_u2_X_23, u2_u2_X_24, u2_u2_X_3, u2_u2_X_31, u2_u2_X_32, u2_u2_X_33, 
       u2_u2_X_34, u2_u2_X_35, u2_u2_X_36, u2_u2_X_37, u2_u2_X_38, u2_u2_X_39, u2_u2_X_4, u2_u2_X_40, u2_u2_X_41, 
       u2_u2_X_42, u2_u2_X_43, u2_u2_X_44, u2_u2_X_45, u2_u2_X_46, u2_u2_X_47, u2_u2_X_48, u2_u2_X_5, u2_u2_X_6, 
       u2_u2_X_7, u2_u2_X_8, u2_u2_X_9, u2_u2_u0_n100, u2_u2_u0_n101, u2_u2_u0_n102, u2_u2_u0_n103, u2_u2_u0_n104, u2_u2_u0_n105, 
       u2_u2_u0_n106, u2_u2_u0_n107, u2_u2_u0_n108, u2_u2_u0_n109, u2_u2_u0_n110, u2_u2_u0_n111, u2_u2_u0_n112, u2_u2_u0_n113, u2_u2_u0_n114, 
       u2_u2_u0_n115, u2_u2_u0_n116, u2_u2_u0_n117, u2_u2_u0_n118, u2_u2_u0_n119, u2_u2_u0_n120, u2_u2_u0_n121, u2_u2_u0_n122, u2_u2_u0_n123, 
       u2_u2_u0_n124, u2_u2_u0_n125, u2_u2_u0_n126, u2_u2_u0_n127, u2_u2_u0_n128, u2_u2_u0_n129, u2_u2_u0_n130, u2_u2_u0_n131, u2_u2_u0_n132, 
       u2_u2_u0_n133, u2_u2_u0_n134, u2_u2_u0_n135, u2_u2_u0_n136, u2_u2_u0_n137, u2_u2_u0_n138, u2_u2_u0_n139, u2_u2_u0_n140, u2_u2_u0_n141, 
       u2_u2_u0_n142, u2_u2_u0_n143, u2_u2_u0_n144, u2_u2_u0_n145, u2_u2_u0_n146, u2_u2_u0_n147, u2_u2_u0_n148, u2_u2_u0_n149, u2_u2_u0_n150, 
       u2_u2_u0_n151, u2_u2_u0_n152, u2_u2_u0_n153, u2_u2_u0_n154, u2_u2_u0_n155, u2_u2_u0_n156, u2_u2_u0_n157, u2_u2_u0_n158, u2_u2_u0_n159, 
       u2_u2_u0_n160, u2_u2_u0_n161, u2_u2_u0_n162, u2_u2_u0_n163, u2_u2_u0_n164, u2_u2_u0_n165, u2_u2_u0_n166, u2_u2_u0_n167, u2_u2_u0_n168, 
       u2_u2_u0_n169, u2_u2_u0_n170, u2_u2_u0_n171, u2_u2_u0_n172, u2_u2_u0_n173, u2_u2_u0_n174, u2_u2_u0_n88, u2_u2_u0_n89, u2_u2_u0_n90, 
       u2_u2_u0_n91, u2_u2_u0_n92, u2_u2_u0_n93, u2_u2_u0_n94, u2_u2_u0_n95, u2_u2_u0_n96, u2_u2_u0_n97, u2_u2_u0_n98, u2_u2_u0_n99, 
       u2_u2_u1_n100, u2_u2_u1_n101, u2_u2_u1_n102, u2_u2_u1_n103, u2_u2_u1_n104, u2_u2_u1_n105, u2_u2_u1_n106, u2_u2_u1_n107, u2_u2_u1_n108, 
       u2_u2_u1_n109, u2_u2_u1_n110, u2_u2_u1_n111, u2_u2_u1_n112, u2_u2_u1_n113, u2_u2_u1_n114, u2_u2_u1_n115, u2_u2_u1_n116, u2_u2_u1_n117, 
       u2_u2_u1_n118, u2_u2_u1_n119, u2_u2_u1_n120, u2_u2_u1_n121, u2_u2_u1_n122, u2_u2_u1_n123, u2_u2_u1_n124, u2_u2_u1_n125, u2_u2_u1_n126, 
       u2_u2_u1_n127, u2_u2_u1_n128, u2_u2_u1_n129, u2_u2_u1_n130, u2_u2_u1_n131, u2_u2_u1_n132, u2_u2_u1_n133, u2_u2_u1_n134, u2_u2_u1_n135, 
       u2_u2_u1_n136, u2_u2_u1_n137, u2_u2_u1_n138, u2_u2_u1_n139, u2_u2_u1_n140, u2_u2_u1_n141, u2_u2_u1_n142, u2_u2_u1_n143, u2_u2_u1_n144, 
       u2_u2_u1_n145, u2_u2_u1_n146, u2_u2_u1_n147, u2_u2_u1_n148, u2_u2_u1_n149, u2_u2_u1_n150, u2_u2_u1_n151, u2_u2_u1_n152, u2_u2_u1_n153, 
       u2_u2_u1_n154, u2_u2_u1_n155, u2_u2_u1_n156, u2_u2_u1_n157, u2_u2_u1_n158, u2_u2_u1_n159, u2_u2_u1_n160, u2_u2_u1_n161, u2_u2_u1_n162, 
       u2_u2_u1_n163, u2_u2_u1_n164, u2_u2_u1_n165, u2_u2_u1_n166, u2_u2_u1_n167, u2_u2_u1_n168, u2_u2_u1_n169, u2_u2_u1_n170, u2_u2_u1_n171, 
       u2_u2_u1_n172, u2_u2_u1_n173, u2_u2_u1_n174, u2_u2_u1_n175, u2_u2_u1_n176, u2_u2_u1_n177, u2_u2_u1_n178, u2_u2_u1_n179, u2_u2_u1_n180, 
       u2_u2_u1_n181, u2_u2_u1_n182, u2_u2_u1_n183, u2_u2_u1_n184, u2_u2_u1_n185, u2_u2_u1_n186, u2_u2_u1_n187, u2_u2_u1_n188, u2_u2_u1_n95, 
       u2_u2_u1_n96, u2_u2_u1_n97, u2_u2_u1_n98, u2_u2_u1_n99, u2_u2_u2_n100, u2_u2_u2_n101, u2_u2_u2_n102, u2_u2_u2_n103, u2_u2_u2_n104, 
       u2_u2_u2_n105, u2_u2_u2_n106, u2_u2_u2_n107, u2_u2_u2_n108, u2_u2_u2_n109, u2_u2_u2_n110, u2_u2_u2_n111, u2_u2_u2_n112, u2_u2_u2_n113, 
       u2_u2_u2_n114, u2_u2_u2_n115, u2_u2_u2_n116, u2_u2_u2_n117, u2_u2_u2_n118, u2_u2_u2_n119, u2_u2_u2_n120, u2_u2_u2_n121, u2_u2_u2_n122, 
       u2_u2_u2_n123, u2_u2_u2_n124, u2_u2_u2_n125, u2_u2_u2_n126, u2_u2_u2_n127, u2_u2_u2_n128, u2_u2_u2_n129, u2_u2_u2_n130, u2_u2_u2_n131, 
       u2_u2_u2_n132, u2_u2_u2_n133, u2_u2_u2_n134, u2_u2_u2_n135, u2_u2_u2_n136, u2_u2_u2_n137, u2_u2_u2_n138, u2_u2_u2_n139, u2_u2_u2_n140, 
       u2_u2_u2_n141, u2_u2_u2_n142, u2_u2_u2_n143, u2_u2_u2_n144, u2_u2_u2_n145, u2_u2_u2_n146, u2_u2_u2_n147, u2_u2_u2_n148, u2_u2_u2_n149, 
       u2_u2_u2_n150, u2_u2_u2_n151, u2_u2_u2_n152, u2_u2_u2_n153, u2_u2_u2_n154, u2_u2_u2_n155, u2_u2_u2_n156, u2_u2_u2_n157, u2_u2_u2_n158, 
       u2_u2_u2_n159, u2_u2_u2_n160, u2_u2_u2_n161, u2_u2_u2_n162, u2_u2_u2_n163, u2_u2_u2_n164, u2_u2_u2_n165, u2_u2_u2_n166, u2_u2_u2_n167, 
       u2_u2_u2_n168, u2_u2_u2_n169, u2_u2_u2_n170, u2_u2_u2_n171, u2_u2_u2_n172, u2_u2_u2_n173, u2_u2_u2_n174, u2_u2_u2_n175, u2_u2_u2_n176, 
       u2_u2_u2_n177, u2_u2_u2_n178, u2_u2_u2_n179, u2_u2_u2_n180, u2_u2_u2_n181, u2_u2_u2_n182, u2_u2_u2_n183, u2_u2_u2_n184, u2_u2_u2_n185, 
       u2_u2_u2_n186, u2_u2_u2_n187, u2_u2_u2_n188, u2_u2_u2_n95, u2_u2_u2_n96, u2_u2_u2_n97, u2_u2_u2_n98, u2_u2_u2_n99, u2_u2_u3_n100, 
       u2_u2_u3_n101, u2_u2_u3_n102, u2_u2_u3_n103, u2_u2_u3_n104, u2_u2_u3_n105, u2_u2_u3_n106, u2_u2_u3_n107, u2_u2_u3_n108, u2_u2_u3_n109, 
       u2_u2_u3_n110, u2_u2_u3_n111, u2_u2_u3_n112, u2_u2_u3_n113, u2_u2_u3_n114, u2_u2_u3_n115, u2_u2_u3_n116, u2_u2_u3_n117, u2_u2_u3_n118, 
       u2_u2_u3_n119, u2_u2_u3_n120, u2_u2_u3_n121, u2_u2_u3_n122, u2_u2_u3_n123, u2_u2_u3_n124, u2_u2_u3_n125, u2_u2_u3_n126, u2_u2_u3_n127, 
       u2_u2_u3_n128, u2_u2_u3_n129, u2_u2_u3_n130, u2_u2_u3_n131, u2_u2_u3_n132, u2_u2_u3_n133, u2_u2_u3_n134, u2_u2_u3_n135, u2_u2_u3_n136, 
       u2_u2_u3_n137, u2_u2_u3_n138, u2_u2_u3_n139, u2_u2_u3_n140, u2_u2_u3_n141, u2_u2_u3_n142, u2_u2_u3_n143, u2_u2_u3_n144, u2_u2_u3_n145, 
       u2_u2_u3_n146, u2_u2_u3_n147, u2_u2_u3_n148, u2_u2_u3_n149, u2_u2_u3_n150, u2_u2_u3_n151, u2_u2_u3_n152, u2_u2_u3_n153, u2_u2_u3_n154, 
       u2_u2_u3_n155, u2_u2_u3_n156, u2_u2_u3_n157, u2_u2_u3_n158, u2_u2_u3_n159, u2_u2_u3_n160, u2_u2_u3_n161, u2_u2_u3_n162, u2_u2_u3_n163, 
       u2_u2_u3_n164, u2_u2_u3_n165, u2_u2_u3_n166, u2_u2_u3_n167, u2_u2_u3_n168, u2_u2_u3_n169, u2_u2_u3_n170, u2_u2_u3_n171, u2_u2_u3_n172, 
       u2_u2_u3_n173, u2_u2_u3_n174, u2_u2_u3_n175, u2_u2_u3_n176, u2_u2_u3_n177, u2_u2_u3_n178, u2_u2_u3_n179, u2_u2_u3_n180, u2_u2_u3_n181, 
       u2_u2_u3_n182, u2_u2_u3_n183, u2_u2_u3_n184, u2_u2_u3_n185, u2_u2_u3_n186, u2_u2_u3_n94, u2_u2_u3_n95, u2_u2_u3_n96, u2_u2_u3_n97, 
       u2_u2_u3_n98, u2_u2_u3_n99, u2_u2_u5_n100, u2_u2_u5_n101, u2_u2_u5_n102, u2_u2_u5_n103, u2_u2_u5_n104, u2_u2_u5_n105, u2_u2_u5_n106, 
       u2_u2_u5_n107, u2_u2_u5_n108, u2_u2_u5_n109, u2_u2_u5_n110, u2_u2_u5_n111, u2_u2_u5_n112, u2_u2_u5_n113, u2_u2_u5_n114, u2_u2_u5_n115, 
       u2_u2_u5_n116, u2_u2_u5_n117, u2_u2_u5_n118, u2_u2_u5_n119, u2_u2_u5_n120, u2_u2_u5_n121, u2_u2_u5_n122, u2_u2_u5_n123, u2_u2_u5_n124, 
       u2_u2_u5_n125, u2_u2_u5_n126, u2_u2_u5_n127, u2_u2_u5_n128, u2_u2_u5_n129, u2_u2_u5_n130, u2_u2_u5_n131, u2_u2_u5_n132, u2_u2_u5_n133, 
       u2_u2_u5_n134, u2_u2_u5_n135, u2_u2_u5_n136, u2_u2_u5_n137, u2_u2_u5_n138, u2_u2_u5_n139, u2_u2_u5_n140, u2_u2_u5_n141, u2_u2_u5_n142, 
       u2_u2_u5_n143, u2_u2_u5_n144, u2_u2_u5_n145, u2_u2_u5_n146, u2_u2_u5_n147, u2_u2_u5_n148, u2_u2_u5_n149, u2_u2_u5_n150, u2_u2_u5_n151, 
       u2_u2_u5_n152, u2_u2_u5_n153, u2_u2_u5_n154, u2_u2_u5_n155, u2_u2_u5_n156, u2_u2_u5_n157, u2_u2_u5_n158, u2_u2_u5_n159, u2_u2_u5_n160, 
       u2_u2_u5_n161, u2_u2_u5_n162, u2_u2_u5_n163, u2_u2_u5_n164, u2_u2_u5_n165, u2_u2_u5_n166, u2_u2_u5_n167, u2_u2_u5_n168, u2_u2_u5_n169, 
       u2_u2_u5_n170, u2_u2_u5_n171, u2_u2_u5_n172, u2_u2_u5_n173, u2_u2_u5_n174, u2_u2_u5_n175, u2_u2_u5_n176, u2_u2_u5_n177, u2_u2_u5_n178, 
       u2_u2_u5_n179, u2_u2_u5_n180, u2_u2_u5_n181, u2_u2_u5_n182, u2_u2_u5_n183, u2_u2_u5_n184, u2_u2_u5_n185, u2_u2_u5_n186, u2_u2_u5_n187, 
       u2_u2_u5_n188, u2_u2_u5_n189, u2_u2_u5_n190, u2_u2_u5_n191, u2_u2_u5_n192, u2_u2_u5_n193, u2_u2_u5_n194, u2_u2_u5_n195, u2_u2_u5_n196, 
       u2_u2_u5_n99, u2_u2_u6_n100, u2_u2_u6_n101, u2_u2_u6_n102, u2_u2_u6_n103, u2_u2_u6_n104, u2_u2_u6_n105, u2_u2_u6_n106, u2_u2_u6_n107, 
       u2_u2_u6_n108, u2_u2_u6_n109, u2_u2_u6_n110, u2_u2_u6_n111, u2_u2_u6_n112, u2_u2_u6_n113, u2_u2_u6_n114, u2_u2_u6_n115, u2_u2_u6_n116, 
       u2_u2_u6_n117, u2_u2_u6_n118, u2_u2_u6_n119, u2_u2_u6_n120, u2_u2_u6_n121, u2_u2_u6_n122, u2_u2_u6_n123, u2_u2_u6_n124, u2_u2_u6_n125, 
       u2_u2_u6_n126, u2_u2_u6_n127, u2_u2_u6_n128, u2_u2_u6_n129, u2_u2_u6_n130, u2_u2_u6_n131, u2_u2_u6_n132, u2_u2_u6_n133, u2_u2_u6_n134, 
       u2_u2_u6_n135, u2_u2_u6_n136, u2_u2_u6_n137, u2_u2_u6_n138, u2_u2_u6_n139, u2_u2_u6_n140, u2_u2_u6_n141, u2_u2_u6_n142, u2_u2_u6_n143, 
       u2_u2_u6_n144, u2_u2_u6_n145, u2_u2_u6_n146, u2_u2_u6_n147, u2_u2_u6_n148, u2_u2_u6_n149, u2_u2_u6_n150, u2_u2_u6_n151, u2_u2_u6_n152, 
       u2_u2_u6_n153, u2_u2_u6_n154, u2_u2_u6_n155, u2_u2_u6_n156, u2_u2_u6_n157, u2_u2_u6_n158, u2_u2_u6_n159, u2_u2_u6_n160, u2_u2_u6_n161, 
       u2_u2_u6_n162, u2_u2_u6_n163, u2_u2_u6_n164, u2_u2_u6_n165, u2_u2_u6_n166, u2_u2_u6_n167, u2_u2_u6_n168, u2_u2_u6_n169, u2_u2_u6_n170, 
       u2_u2_u6_n171, u2_u2_u6_n172, u2_u2_u6_n173, u2_u2_u6_n174, u2_u2_u6_n88, u2_u2_u6_n89, u2_u2_u6_n90, u2_u2_u6_n91, u2_u2_u6_n92, 
       u2_u2_u6_n93, u2_u2_u6_n94, u2_u2_u6_n95, u2_u2_u6_n96, u2_u2_u6_n97, u2_u2_u6_n98, u2_u2_u6_n99, u2_u2_u7_n100, u2_u2_u7_n101, 
       u2_u2_u7_n102, u2_u2_u7_n103, u2_u2_u7_n104, u2_u2_u7_n105, u2_u2_u7_n106, u2_u2_u7_n107, u2_u2_u7_n108, u2_u2_u7_n109, u2_u2_u7_n110, 
       u2_u2_u7_n111, u2_u2_u7_n112, u2_u2_u7_n113, u2_u2_u7_n114, u2_u2_u7_n115, u2_u2_u7_n116, u2_u2_u7_n117, u2_u2_u7_n118, u2_u2_u7_n119, 
       u2_u2_u7_n120, u2_u2_u7_n121, u2_u2_u7_n122, u2_u2_u7_n123, u2_u2_u7_n124, u2_u2_u7_n125, u2_u2_u7_n126, u2_u2_u7_n127, u2_u2_u7_n128, 
       u2_u2_u7_n129, u2_u2_u7_n130, u2_u2_u7_n131, u2_u2_u7_n132, u2_u2_u7_n133, u2_u2_u7_n134, u2_u2_u7_n135, u2_u2_u7_n136, u2_u2_u7_n137, 
       u2_u2_u7_n138, u2_u2_u7_n139, u2_u2_u7_n140, u2_u2_u7_n141, u2_u2_u7_n142, u2_u2_u7_n143, u2_u2_u7_n144, u2_u2_u7_n145, u2_u2_u7_n146, 
       u2_u2_u7_n147, u2_u2_u7_n148, u2_u2_u7_n149, u2_u2_u7_n150, u2_u2_u7_n151, u2_u2_u7_n152, u2_u2_u7_n153, u2_u2_u7_n154, u2_u2_u7_n155, 
       u2_u2_u7_n156, u2_u2_u7_n157, u2_u2_u7_n158, u2_u2_u7_n159, u2_u2_u7_n160, u2_u2_u7_n161, u2_u2_u7_n162, u2_u2_u7_n163, u2_u2_u7_n164, 
       u2_u2_u7_n165, u2_u2_u7_n166, u2_u2_u7_n167, u2_u2_u7_n168, u2_u2_u7_n169, u2_u2_u7_n170, u2_u2_u7_n171, u2_u2_u7_n172, u2_u2_u7_n173, 
       u2_u2_u7_n174, u2_u2_u7_n175, u2_u2_u7_n176, u2_u2_u7_n177, u2_u2_u7_n178, u2_u2_u7_n179, u2_u2_u7_n180, u2_u2_u7_n91, u2_u2_u7_n92, 
       u2_u2_u7_n93, u2_u2_u7_n94, u2_u2_u7_n95, u2_u2_u7_n96, u2_u2_u7_n97, u2_u2_u7_n98, u2_u2_u7_n99, u2_u3_X_13, u2_u3_X_14, 
       u2_u3_X_15, u2_u3_X_16, u2_u3_X_17, u2_u3_X_18, u2_u3_X_19, u2_u3_X_20, u2_u3_X_21, u2_u3_X_22, u2_u3_X_23, 
       u2_u3_X_24, u2_u3_X_25, u2_u3_X_26, u2_u3_X_27, u2_u3_X_28, u2_u3_X_29, u2_u3_X_30, u2_u3_X_31, u2_u3_X_32, 
       u2_u3_X_33, u2_u3_X_34, u2_u3_X_35, u2_u3_X_36, u2_u3_u2_n100, u2_u3_u2_n101, u2_u3_u2_n102, u2_u3_u2_n103, u2_u3_u2_n104, 
       u2_u3_u2_n105, u2_u3_u2_n106, u2_u3_u2_n107, u2_u3_u2_n108, u2_u3_u2_n109, u2_u3_u2_n110, u2_u3_u2_n111, u2_u3_u2_n112, u2_u3_u2_n113, 
       u2_u3_u2_n114, u2_u3_u2_n115, u2_u3_u2_n116, u2_u3_u2_n117, u2_u3_u2_n118, u2_u3_u2_n119, u2_u3_u2_n120, u2_u3_u2_n121, u2_u3_u2_n122, 
       u2_u3_u2_n123, u2_u3_u2_n124, u2_u3_u2_n125, u2_u3_u2_n126, u2_u3_u2_n127, u2_u3_u2_n128, u2_u3_u2_n129, u2_u3_u2_n130, u2_u3_u2_n131, 
       u2_u3_u2_n132, u2_u3_u2_n133, u2_u3_u2_n134, u2_u3_u2_n135, u2_u3_u2_n136, u2_u3_u2_n137, u2_u3_u2_n138, u2_u3_u2_n139, u2_u3_u2_n140, 
       u2_u3_u2_n141, u2_u3_u2_n142, u2_u3_u2_n143, u2_u3_u2_n144, u2_u3_u2_n145, u2_u3_u2_n146, u2_u3_u2_n147, u2_u3_u2_n148, u2_u3_u2_n149, 
       u2_u3_u2_n150, u2_u3_u2_n151, u2_u3_u2_n152, u2_u3_u2_n153, u2_u3_u2_n154, u2_u3_u2_n155, u2_u3_u2_n156, u2_u3_u2_n157, u2_u3_u2_n158, 
       u2_u3_u2_n159, u2_u3_u2_n160, u2_u3_u2_n161, u2_u3_u2_n162, u2_u3_u2_n163, u2_u3_u2_n164, u2_u3_u2_n165, u2_u3_u2_n166, u2_u3_u2_n167, 
       u2_u3_u2_n168, u2_u3_u2_n169, u2_u3_u2_n170, u2_u3_u2_n171, u2_u3_u2_n172, u2_u3_u2_n173, u2_u3_u2_n174, u2_u3_u2_n175, u2_u3_u2_n176, 
       u2_u3_u2_n177, u2_u3_u2_n178, u2_u3_u2_n179, u2_u3_u2_n180, u2_u3_u2_n181, u2_u3_u2_n182, u2_u3_u2_n183, u2_u3_u2_n184, u2_u3_u2_n185, 
       u2_u3_u2_n186, u2_u3_u2_n187, u2_u3_u2_n188, u2_u3_u2_n95, u2_u3_u2_n96, u2_u3_u2_n97, u2_u3_u2_n98, u2_u3_u2_n99, u2_u3_u3_n100, 
       u2_u3_u3_n101, u2_u3_u3_n102, u2_u3_u3_n103, u2_u3_u3_n104, u2_u3_u3_n105, u2_u3_u3_n106, u2_u3_u3_n107, u2_u3_u3_n108, u2_u3_u3_n109, 
       u2_u3_u3_n110, u2_u3_u3_n111, u2_u3_u3_n112, u2_u3_u3_n113, u2_u3_u3_n114, u2_u3_u3_n115, u2_u3_u3_n116, u2_u3_u3_n117, u2_u3_u3_n118, 
       u2_u3_u3_n119, u2_u3_u3_n120, u2_u3_u3_n121, u2_u3_u3_n122, u2_u3_u3_n123, u2_u3_u3_n124, u2_u3_u3_n125, u2_u3_u3_n126, u2_u3_u3_n127, 
       u2_u3_u3_n128, u2_u3_u3_n129, u2_u3_u3_n130, u2_u3_u3_n131, u2_u3_u3_n132, u2_u3_u3_n133, u2_u3_u3_n134, u2_u3_u3_n135, u2_u3_u3_n136, 
       u2_u3_u3_n137, u2_u3_u3_n138, u2_u3_u3_n139, u2_u3_u3_n140, u2_u3_u3_n141, u2_u3_u3_n142, u2_u3_u3_n143, u2_u3_u3_n144, u2_u3_u3_n145, 
       u2_u3_u3_n146, u2_u3_u3_n147, u2_u3_u3_n148, u2_u3_u3_n149, u2_u3_u3_n150, u2_u3_u3_n151, u2_u3_u3_n152, u2_u3_u3_n153, u2_u3_u3_n154, 
       u2_u3_u3_n155, u2_u3_u3_n156, u2_u3_u3_n157, u2_u3_u3_n158, u2_u3_u3_n159, u2_u3_u3_n160, u2_u3_u3_n161, u2_u3_u3_n162, u2_u3_u3_n163, 
       u2_u3_u3_n164, u2_u3_u3_n165, u2_u3_u3_n166, u2_u3_u3_n167, u2_u3_u3_n168, u2_u3_u3_n169, u2_u3_u3_n170, u2_u3_u3_n171, u2_u3_u3_n172, 
       u2_u3_u3_n173, u2_u3_u3_n174, u2_u3_u3_n175, u2_u3_u3_n176, u2_u3_u3_n177, u2_u3_u3_n178, u2_u3_u3_n179, u2_u3_u3_n180, u2_u3_u3_n181, 
       u2_u3_u3_n182, u2_u3_u3_n183, u2_u3_u3_n184, u2_u3_u3_n185, u2_u3_u3_n186, u2_u3_u3_n94, u2_u3_u3_n95, u2_u3_u3_n96, u2_u3_u3_n97, 
       u2_u3_u3_n98, u2_u3_u3_n99, u2_u3_u4_n100, u2_u3_u4_n101, u2_u3_u4_n102, u2_u3_u4_n103, u2_u3_u4_n104, u2_u3_u4_n105, u2_u3_u4_n106, 
       u2_u3_u4_n107, u2_u3_u4_n108, u2_u3_u4_n109, u2_u3_u4_n110, u2_u3_u4_n111, u2_u3_u4_n112, u2_u3_u4_n113, u2_u3_u4_n114, u2_u3_u4_n115, 
       u2_u3_u4_n116, u2_u3_u4_n117, u2_u3_u4_n118, u2_u3_u4_n119, u2_u3_u4_n120, u2_u3_u4_n121, u2_u3_u4_n122, u2_u3_u4_n123, u2_u3_u4_n124, 
       u2_u3_u4_n125, u2_u3_u4_n126, u2_u3_u4_n127, u2_u3_u4_n128, u2_u3_u4_n129, u2_u3_u4_n130, u2_u3_u4_n131, u2_u3_u4_n132, u2_u3_u4_n133, 
       u2_u3_u4_n134, u2_u3_u4_n135, u2_u3_u4_n136, u2_u3_u4_n137, u2_u3_u4_n138, u2_u3_u4_n139, u2_u3_u4_n140, u2_u3_u4_n141, u2_u3_u4_n142, 
       u2_u3_u4_n143, u2_u3_u4_n144, u2_u3_u4_n145, u2_u3_u4_n146, u2_u3_u4_n147, u2_u3_u4_n148, u2_u3_u4_n149, u2_u3_u4_n150, u2_u3_u4_n151, 
       u2_u3_u4_n152, u2_u3_u4_n153, u2_u3_u4_n154, u2_u3_u4_n155, u2_u3_u4_n156, u2_u3_u4_n157, u2_u3_u4_n158, u2_u3_u4_n159, u2_u3_u4_n160, 
       u2_u3_u4_n161, u2_u3_u4_n162, u2_u3_u4_n163, u2_u3_u4_n164, u2_u3_u4_n165, u2_u3_u4_n166, u2_u3_u4_n167, u2_u3_u4_n168, u2_u3_u4_n169, 
       u2_u3_u4_n170, u2_u3_u4_n171, u2_u3_u4_n172, u2_u3_u4_n173, u2_u3_u4_n174, u2_u3_u4_n175, u2_u3_u4_n176, u2_u3_u4_n177, u2_u3_u4_n178, 
       u2_u3_u4_n179, u2_u3_u4_n180, u2_u3_u4_n181, u2_u3_u4_n182, u2_u3_u4_n183, u2_u3_u4_n184, u2_u3_u4_n185, u2_u3_u4_n186, u2_u3_u4_n94, 
       u2_u3_u4_n95, u2_u3_u4_n96, u2_u3_u4_n97, u2_u3_u4_n98, u2_u3_u4_n99, u2_u3_u5_n100, u2_u3_u5_n101, u2_u3_u5_n102, u2_u3_u5_n103, 
       u2_u3_u5_n104, u2_u3_u5_n105, u2_u3_u5_n106, u2_u3_u5_n107, u2_u3_u5_n108, u2_u3_u5_n109, u2_u3_u5_n110, u2_u3_u5_n111, u2_u3_u5_n112, 
       u2_u3_u5_n113, u2_u3_u5_n114, u2_u3_u5_n115, u2_u3_u5_n116, u2_u3_u5_n117, u2_u3_u5_n118, u2_u3_u5_n119, u2_u3_u5_n120, u2_u3_u5_n121, 
       u2_u3_u5_n122, u2_u3_u5_n123, u2_u3_u5_n124, u2_u3_u5_n125, u2_u3_u5_n126, u2_u3_u5_n127, u2_u3_u5_n128, u2_u3_u5_n129, u2_u3_u5_n130, 
       u2_u3_u5_n131, u2_u3_u5_n132, u2_u3_u5_n133, u2_u3_u5_n134, u2_u3_u5_n135, u2_u3_u5_n136, u2_u3_u5_n137, u2_u3_u5_n138, u2_u3_u5_n139, 
       u2_u3_u5_n140, u2_u3_u5_n141, u2_u3_u5_n142, u2_u3_u5_n143, u2_u3_u5_n144, u2_u3_u5_n145, u2_u3_u5_n146, u2_u3_u5_n147, u2_u3_u5_n148, 
       u2_u3_u5_n149, u2_u3_u5_n150, u2_u3_u5_n151, u2_u3_u5_n152, u2_u3_u5_n153, u2_u3_u5_n154, u2_u3_u5_n155, u2_u3_u5_n156, u2_u3_u5_n157, 
       u2_u3_u5_n158, u2_u3_u5_n159, u2_u3_u5_n160, u2_u3_u5_n161, u2_u3_u5_n162, u2_u3_u5_n163, u2_u3_u5_n164, u2_u3_u5_n165, u2_u3_u5_n166, 
       u2_u3_u5_n167, u2_u3_u5_n168, u2_u3_u5_n169, u2_u3_u5_n170, u2_u3_u5_n171, u2_u3_u5_n172, u2_u3_u5_n173, u2_u3_u5_n174, u2_u3_u5_n175, 
       u2_u3_u5_n176, u2_u3_u5_n177, u2_u3_u5_n178, u2_u3_u5_n179, u2_u3_u5_n180, u2_u3_u5_n181, u2_u3_u5_n182, u2_u3_u5_n183, u2_u3_u5_n184, 
       u2_u3_u5_n185, u2_u3_u5_n186, u2_u3_u5_n187, u2_u3_u5_n188, u2_u3_u5_n189, u2_u3_u5_n190, u2_u3_u5_n191, u2_u3_u5_n192, u2_u3_u5_n193, 
       u2_u3_u5_n194, u2_u3_u5_n195, u2_u3_u5_n196, u2_u3_u5_n99, u2_u4_X_10, u2_u4_X_11, u2_u4_X_12, u2_u4_X_13, u2_u4_X_14, 
       u2_u4_X_15, u2_u4_X_16, u2_u4_X_17, u2_u4_X_18, u2_u4_X_19, u2_u4_X_20, u2_u4_X_21, u2_u4_X_22, u2_u4_X_23, 
       u2_u4_X_24, u2_u4_X_7, u2_u4_X_8, u2_u4_X_9, u2_u4_u1_n100, u2_u4_u1_n101, u2_u4_u1_n102, u2_u4_u1_n103, u2_u4_u1_n104, 
       u2_u4_u1_n105, u2_u4_u1_n106, u2_u4_u1_n107, u2_u4_u1_n108, u2_u4_u1_n109, u2_u4_u1_n110, u2_u4_u1_n111, u2_u4_u1_n112, u2_u4_u1_n113, 
       u2_u4_u1_n114, u2_u4_u1_n115, u2_u4_u1_n116, u2_u4_u1_n117, u2_u4_u1_n118, u2_u4_u1_n119, u2_u4_u1_n120, u2_u4_u1_n121, u2_u4_u1_n122, 
       u2_u4_u1_n123, u2_u4_u1_n124, u2_u4_u1_n125, u2_u4_u1_n126, u2_u4_u1_n127, u2_u4_u1_n128, u2_u4_u1_n129, u2_u4_u1_n130, u2_u4_u1_n131, 
       u2_u4_u1_n132, u2_u4_u1_n133, u2_u4_u1_n134, u2_u4_u1_n135, u2_u4_u1_n136, u2_u4_u1_n137, u2_u4_u1_n138, u2_u4_u1_n139, u2_u4_u1_n140, 
       u2_u4_u1_n141, u2_u4_u1_n142, u2_u4_u1_n143, u2_u4_u1_n144, u2_u4_u1_n145, u2_u4_u1_n146, u2_u4_u1_n147, u2_u4_u1_n148, u2_u4_u1_n149, 
       u2_u4_u1_n150, u2_u4_u1_n151, u2_u4_u1_n152, u2_u4_u1_n153, u2_u4_u1_n154, u2_u4_u1_n155, u2_u4_u1_n156, u2_u4_u1_n157, u2_u4_u1_n158, 
       u2_u4_u1_n159, u2_u4_u1_n160, u2_u4_u1_n161, u2_u4_u1_n162, u2_u4_u1_n163, u2_u4_u1_n164, u2_u4_u1_n165, u2_u4_u1_n166, u2_u4_u1_n167, 
       u2_u4_u1_n168, u2_u4_u1_n169, u2_u4_u1_n170, u2_u4_u1_n171, u2_u4_u1_n172, u2_u4_u1_n173, u2_u4_u1_n174, u2_u4_u1_n175, u2_u4_u1_n176, 
       u2_u4_u1_n177, u2_u4_u1_n178, u2_u4_u1_n179, u2_u4_u1_n180, u2_u4_u1_n181, u2_u4_u1_n182, u2_u4_u1_n183, u2_u4_u1_n184, u2_u4_u1_n185, 
       u2_u4_u1_n186, u2_u4_u1_n187, u2_u4_u1_n188, u2_u4_u1_n95, u2_u4_u1_n96, u2_u4_u1_n97, u2_u4_u1_n98, u2_u4_u1_n99, u2_u4_u2_n100, 
       u2_u4_u2_n101, u2_u4_u2_n102, u2_u4_u2_n103, u2_u4_u2_n104, u2_u4_u2_n105, u2_u4_u2_n106, u2_u4_u2_n107, u2_u4_u2_n108, u2_u4_u2_n109, 
       u2_u4_u2_n110, u2_u4_u2_n111, u2_u4_u2_n112, u2_u4_u2_n113, u2_u4_u2_n114, u2_u4_u2_n115, u2_u4_u2_n116, u2_u4_u2_n117, u2_u4_u2_n118, 
       u2_u4_u2_n119, u2_u4_u2_n120, u2_u4_u2_n121, u2_u4_u2_n122, u2_u4_u2_n123, u2_u4_u2_n124, u2_u4_u2_n125, u2_u4_u2_n126, u2_u4_u2_n127, 
       u2_u4_u2_n128, u2_u4_u2_n129, u2_u4_u2_n130, u2_u4_u2_n131, u2_u4_u2_n132, u2_u4_u2_n133, u2_u4_u2_n134, u2_u4_u2_n135, u2_u4_u2_n136, 
       u2_u4_u2_n137, u2_u4_u2_n138, u2_u4_u2_n139, u2_u4_u2_n140, u2_u4_u2_n141, u2_u4_u2_n142, u2_u4_u2_n143, u2_u4_u2_n144, u2_u4_u2_n145, 
       u2_u4_u2_n146, u2_u4_u2_n147, u2_u4_u2_n148, u2_u4_u2_n149, u2_u4_u2_n150, u2_u4_u2_n151, u2_u4_u2_n152, u2_u4_u2_n153, u2_u4_u2_n154, 
       u2_u4_u2_n155, u2_u4_u2_n156, u2_u4_u2_n157, u2_u4_u2_n158, u2_u4_u2_n159, u2_u4_u2_n160, u2_u4_u2_n161, u2_u4_u2_n162, u2_u4_u2_n163, 
       u2_u4_u2_n164, u2_u4_u2_n165, u2_u4_u2_n166, u2_u4_u2_n167, u2_u4_u2_n168, u2_u4_u2_n169, u2_u4_u2_n170, u2_u4_u2_n171, u2_u4_u2_n172, 
       u2_u4_u2_n173, u2_u4_u2_n174, u2_u4_u2_n175, u2_u4_u2_n176, u2_u4_u2_n177, u2_u4_u2_n178, u2_u4_u2_n179, u2_u4_u2_n180, u2_u4_u2_n181, 
       u2_u4_u2_n182, u2_u4_u2_n183, u2_u4_u2_n184, u2_u4_u2_n185, u2_u4_u2_n186, u2_u4_u2_n187, u2_u4_u2_n188, u2_u4_u2_n95, u2_u4_u2_n96, 
       u2_u4_u2_n97, u2_u4_u2_n98, u2_u4_u2_n99, u2_u4_u3_n100, u2_u4_u3_n101, u2_u4_u3_n102, u2_u4_u3_n103, u2_u4_u3_n104, u2_u4_u3_n105, 
       u2_u4_u3_n106, u2_u4_u3_n107, u2_u4_u3_n108, u2_u4_u3_n109, u2_u4_u3_n110, u2_u4_u3_n111, u2_u4_u3_n112, u2_u4_u3_n113, u2_u4_u3_n114, 
       u2_u4_u3_n115, u2_u4_u3_n116, u2_u4_u3_n117, u2_u4_u3_n118, u2_u4_u3_n119, u2_u4_u3_n120, u2_u4_u3_n121, u2_u4_u3_n122, u2_u4_u3_n123, 
       u2_u4_u3_n124, u2_u4_u3_n125, u2_u4_u3_n126, u2_u4_u3_n127, u2_u4_u3_n128, u2_u4_u3_n129, u2_u4_u3_n130, u2_u4_u3_n131, u2_u4_u3_n132, 
       u2_u4_u3_n133, u2_u4_u3_n134, u2_u4_u3_n135, u2_u4_u3_n136, u2_u4_u3_n137, u2_u4_u3_n138, u2_u4_u3_n139, u2_u4_u3_n140, u2_u4_u3_n141, 
       u2_u4_u3_n142, u2_u4_u3_n143, u2_u4_u3_n144, u2_u4_u3_n145, u2_u4_u3_n146, u2_u4_u3_n147, u2_u4_u3_n148, u2_u4_u3_n149, u2_u4_u3_n150, 
       u2_u4_u3_n151, u2_u4_u3_n152, u2_u4_u3_n153, u2_u4_u3_n154, u2_u4_u3_n155, u2_u4_u3_n156, u2_u4_u3_n157, u2_u4_u3_n158, u2_u4_u3_n159, 
       u2_u4_u3_n160, u2_u4_u3_n161, u2_u4_u3_n162, u2_u4_u3_n163, u2_u4_u3_n164, u2_u4_u3_n165, u2_u4_u3_n166, u2_u4_u3_n167, u2_u4_u3_n168, 
       u2_u4_u3_n169, u2_u4_u3_n170, u2_u4_u3_n171, u2_u4_u3_n172, u2_u4_u3_n173, u2_u4_u3_n174, u2_u4_u3_n175, u2_u4_u3_n176, u2_u4_u3_n177, 
       u2_u4_u3_n178, u2_u4_u3_n179, u2_u4_u3_n180, u2_u4_u3_n181, u2_u4_u3_n182, u2_u4_u3_n183, u2_u4_u3_n184, u2_u4_u3_n185, u2_u4_u3_n186, 
       u2_u4_u3_n94, u2_u4_u3_n95, u2_u4_u3_n96, u2_u4_u3_n97, u2_u4_u3_n98, u2_u4_u3_n99, u2_u5_X_19, u2_u5_X_20, u2_u5_X_21, 
       u2_u5_X_22, u2_u5_X_23, u2_u5_X_24, u2_u5_X_25, u2_u5_X_26, u2_u5_X_27, u2_u5_X_28, u2_u5_X_29, u2_u5_X_30, 
       u2_u5_u3_n100, u2_u5_u3_n101, u2_u5_u3_n102, u2_u5_u3_n103, u2_u5_u3_n104, u2_u5_u3_n105, u2_u5_u3_n106, u2_u5_u3_n107, u2_u5_u3_n108, 
       u2_u5_u3_n109, u2_u5_u3_n110, u2_u5_u3_n111, u2_u5_u3_n112, u2_u5_u3_n113, u2_u5_u3_n114, u2_u5_u3_n115, u2_u5_u3_n116, u2_u5_u3_n117, 
       u2_u5_u3_n118, u2_u5_u3_n119, u2_u5_u3_n120, u2_u5_u3_n121, u2_u5_u3_n122, u2_u5_u3_n123, u2_u5_u3_n124, u2_u5_u3_n125, u2_u5_u3_n126, 
       u2_u5_u3_n127, u2_u5_u3_n128, u2_u5_u3_n129, u2_u5_u3_n130, u2_u5_u3_n131, u2_u5_u3_n132, u2_u5_u3_n133, u2_u5_u3_n134, u2_u5_u3_n135, 
       u2_u5_u3_n136, u2_u5_u3_n137, u2_u5_u3_n138, u2_u5_u3_n139, u2_u5_u3_n140, u2_u5_u3_n141, u2_u5_u3_n142, u2_u5_u3_n143, u2_u5_u3_n144, 
       u2_u5_u3_n145, u2_u5_u3_n146, u2_u5_u3_n147, u2_u5_u3_n148, u2_u5_u3_n149, u2_u5_u3_n150, u2_u5_u3_n151, u2_u5_u3_n152, u2_u5_u3_n153, 
       u2_u5_u3_n154, u2_u5_u3_n155, u2_u5_u3_n156, u2_u5_u3_n157, u2_u5_u3_n158, u2_u5_u3_n159, u2_u5_u3_n160, u2_u5_u3_n161, u2_u5_u3_n162, 
       u2_u5_u3_n163, u2_u5_u3_n164, u2_u5_u3_n165, u2_u5_u3_n166, u2_u5_u3_n167, u2_u5_u3_n168, u2_u5_u3_n169, u2_u5_u3_n170, u2_u5_u3_n171, 
       u2_u5_u3_n172, u2_u5_u3_n173, u2_u5_u3_n174, u2_u5_u3_n175, u2_u5_u3_n176, u2_u5_u3_n177, u2_u5_u3_n178, u2_u5_u3_n179, u2_u5_u3_n180, 
       u2_u5_u3_n181, u2_u5_u3_n182, u2_u5_u3_n183, u2_u5_u3_n184, u2_u5_u3_n185, u2_u5_u3_n186, u2_u5_u3_n94, u2_u5_u3_n95, u2_u5_u3_n96, 
       u2_u5_u3_n97, u2_u5_u3_n98, u2_u5_u3_n99, u2_u5_u4_n100, u2_u5_u4_n101, u2_u5_u4_n102, u2_u5_u4_n103, u2_u5_u4_n104, u2_u5_u4_n105, 
       u2_u5_u4_n106, u2_u5_u4_n107, u2_u5_u4_n108, u2_u5_u4_n109, u2_u5_u4_n110, u2_u5_u4_n111, u2_u5_u4_n112, u2_u5_u4_n113, u2_u5_u4_n114, 
       u2_u5_u4_n115, u2_u5_u4_n116, u2_u5_u4_n117, u2_u5_u4_n118, u2_u5_u4_n119, u2_u5_u4_n120, u2_u5_u4_n121, u2_u5_u4_n122, u2_u5_u4_n123, 
       u2_u5_u4_n124, u2_u5_u4_n125, u2_u5_u4_n126, u2_u5_u4_n127, u2_u5_u4_n128, u2_u5_u4_n129, u2_u5_u4_n130, u2_u5_u4_n131, u2_u5_u4_n132, 
       u2_u5_u4_n133, u2_u5_u4_n134, u2_u5_u4_n135, u2_u5_u4_n136, u2_u5_u4_n137, u2_u5_u4_n138, u2_u5_u4_n139, u2_u5_u4_n140, u2_u5_u4_n141, 
       u2_u5_u4_n142, u2_u5_u4_n143, u2_u5_u4_n144, u2_u5_u4_n145, u2_u5_u4_n146, u2_u5_u4_n147, u2_u5_u4_n148, u2_u5_u4_n149, u2_u5_u4_n150, 
       u2_u5_u4_n151, u2_u5_u4_n152, u2_u5_u4_n153, u2_u5_u4_n154, u2_u5_u4_n155, u2_u5_u4_n156, u2_u5_u4_n157, u2_u5_u4_n158, u2_u5_u4_n159, 
       u2_u5_u4_n160, u2_u5_u4_n161, u2_u5_u4_n162, u2_u5_u4_n163, u2_u5_u4_n164, u2_u5_u4_n165, u2_u5_u4_n166, u2_u5_u4_n167, u2_u5_u4_n168, 
       u2_u5_u4_n169, u2_u5_u4_n170, u2_u5_u4_n171, u2_u5_u4_n172, u2_u5_u4_n173, u2_u5_u4_n174, u2_u5_u4_n175, u2_u5_u4_n176, u2_u5_u4_n177, 
       u2_u5_u4_n178, u2_u5_u4_n179, u2_u5_u4_n180, u2_u5_u4_n181, u2_u5_u4_n182, u2_u5_u4_n183, u2_u5_u4_n184, u2_u5_u4_n185, u2_u5_u4_n186, 
       u2_u5_u4_n94, u2_u5_u4_n95, u2_u5_u4_n96, u2_u5_u4_n97, u2_u5_u4_n98, u2_u5_u4_n99, u2_u6_X_1, u2_u6_X_10, u2_u6_X_11, 
       u2_u6_X_12, u2_u6_X_13, u2_u6_X_14, u2_u6_X_15, u2_u6_X_16, u2_u6_X_17, u2_u6_X_18, u2_u6_X_19, u2_u6_X_2, 
       u2_u6_X_20, u2_u6_X_21, u2_u6_X_22, u2_u6_X_23, u2_u6_X_24, u2_u6_X_25, u2_u6_X_26, u2_u6_X_27, u2_u6_X_28, 
       u2_u6_X_29, u2_u6_X_3, u2_u6_X_30, u2_u6_X_37, u2_u6_X_38, u2_u6_X_39, u2_u6_X_4, u2_u6_X_40, u2_u6_X_41, 
       u2_u6_X_42, u2_u6_X_43, u2_u6_X_44, u2_u6_X_45, u2_u6_X_46, u2_u6_X_47, u2_u6_X_48, u2_u6_X_5, u2_u6_X_6, 
       u2_u6_X_7, u2_u6_X_8, u2_u6_X_9, u2_u6_u0_n100, u2_u6_u0_n101, u2_u6_u0_n102, u2_u6_u0_n103, u2_u6_u0_n104, u2_u6_u0_n105, 
       u2_u6_u0_n106, u2_u6_u0_n107, u2_u6_u0_n108, u2_u6_u0_n109, u2_u6_u0_n110, u2_u6_u0_n111, u2_u6_u0_n112, u2_u6_u0_n113, u2_u6_u0_n114, 
       u2_u6_u0_n115, u2_u6_u0_n116, u2_u6_u0_n117, u2_u6_u0_n118, u2_u6_u0_n119, u2_u6_u0_n120, u2_u6_u0_n121, u2_u6_u0_n122, u2_u6_u0_n123, 
       u2_u6_u0_n124, u2_u6_u0_n125, u2_u6_u0_n126, u2_u6_u0_n127, u2_u6_u0_n128, u2_u6_u0_n129, u2_u6_u0_n130, u2_u6_u0_n131, u2_u6_u0_n132, 
       u2_u6_u0_n133, u2_u6_u0_n134, u2_u6_u0_n135, u2_u6_u0_n136, u2_u6_u0_n137, u2_u6_u0_n138, u2_u6_u0_n139, u2_u6_u0_n140, u2_u6_u0_n141, 
       u2_u6_u0_n142, u2_u6_u0_n143, u2_u6_u0_n144, u2_u6_u0_n145, u2_u6_u0_n146, u2_u6_u0_n147, u2_u6_u0_n148, u2_u6_u0_n149, u2_u6_u0_n150, 
       u2_u6_u0_n151, u2_u6_u0_n152, u2_u6_u0_n153, u2_u6_u0_n154, u2_u6_u0_n155, u2_u6_u0_n156, u2_u6_u0_n157, u2_u6_u0_n158, u2_u6_u0_n159, 
       u2_u6_u0_n160, u2_u6_u0_n161, u2_u6_u0_n162, u2_u6_u0_n163, u2_u6_u0_n164, u2_u6_u0_n165, u2_u6_u0_n166, u2_u6_u0_n167, u2_u6_u0_n168, 
       u2_u6_u0_n169, u2_u6_u0_n170, u2_u6_u0_n171, u2_u6_u0_n172, u2_u6_u0_n173, u2_u6_u0_n174, u2_u6_u0_n88, u2_u6_u0_n89, u2_u6_u0_n90, 
       u2_u6_u0_n91, u2_u6_u0_n92, u2_u6_u0_n93, u2_u6_u0_n94, u2_u6_u0_n95, u2_u6_u0_n96, u2_u6_u0_n97, u2_u6_u0_n98, u2_u6_u0_n99, 
       u2_u6_u1_n100, u2_u6_u1_n101, u2_u6_u1_n102, u2_u6_u1_n103, u2_u6_u1_n104, u2_u6_u1_n105, u2_u6_u1_n106, u2_u6_u1_n107, u2_u6_u1_n108, 
       u2_u6_u1_n109, u2_u6_u1_n110, u2_u6_u1_n111, u2_u6_u1_n112, u2_u6_u1_n113, u2_u6_u1_n114, u2_u6_u1_n115, u2_u6_u1_n116, u2_u6_u1_n117, 
       u2_u6_u1_n118, u2_u6_u1_n119, u2_u6_u1_n120, u2_u6_u1_n121, u2_u6_u1_n122, u2_u6_u1_n123, u2_u6_u1_n124, u2_u6_u1_n125, u2_u6_u1_n126, 
       u2_u6_u1_n127, u2_u6_u1_n128, u2_u6_u1_n129, u2_u6_u1_n130, u2_u6_u1_n131, u2_u6_u1_n132, u2_u6_u1_n133, u2_u6_u1_n134, u2_u6_u1_n135, 
       u2_u6_u1_n136, u2_u6_u1_n137, u2_u6_u1_n138, u2_u6_u1_n139, u2_u6_u1_n140, u2_u6_u1_n141, u2_u6_u1_n142, u2_u6_u1_n143, u2_u6_u1_n144, 
       u2_u6_u1_n145, u2_u6_u1_n146, u2_u6_u1_n147, u2_u6_u1_n148, u2_u6_u1_n149, u2_u6_u1_n150, u2_u6_u1_n151, u2_u6_u1_n152, u2_u6_u1_n153, 
       u2_u6_u1_n154, u2_u6_u1_n155, u2_u6_u1_n156, u2_u6_u1_n157, u2_u6_u1_n158, u2_u6_u1_n159, u2_u6_u1_n160, u2_u6_u1_n161, u2_u6_u1_n162, 
       u2_u6_u1_n163, u2_u6_u1_n164, u2_u6_u1_n165, u2_u6_u1_n166, u2_u6_u1_n167, u2_u6_u1_n168, u2_u6_u1_n169, u2_u6_u1_n170, u2_u6_u1_n171, 
       u2_u6_u1_n172, u2_u6_u1_n173, u2_u6_u1_n174, u2_u6_u1_n175, u2_u6_u1_n176, u2_u6_u1_n177, u2_u6_u1_n178, u2_u6_u1_n179, u2_u6_u1_n180, 
       u2_u6_u1_n181, u2_u6_u1_n182, u2_u6_u1_n183, u2_u6_u1_n184, u2_u6_u1_n185, u2_u6_u1_n186, u2_u6_u1_n187, u2_u6_u1_n188, u2_u6_u1_n95, 
       u2_u6_u1_n96, u2_u6_u1_n97, u2_u6_u1_n98, u2_u6_u1_n99, u2_u6_u2_n100, u2_u6_u2_n101, u2_u6_u2_n102, u2_u6_u2_n103, u2_u6_u2_n104, 
       u2_u6_u2_n105, u2_u6_u2_n106, u2_u6_u2_n107, u2_u6_u2_n108, u2_u6_u2_n109, u2_u6_u2_n110, u2_u6_u2_n111, u2_u6_u2_n112, u2_u6_u2_n113, 
       u2_u6_u2_n114, u2_u6_u2_n115, u2_u6_u2_n116, u2_u6_u2_n117, u2_u6_u2_n118, u2_u6_u2_n119, u2_u6_u2_n120, u2_u6_u2_n121, u2_u6_u2_n122, 
       u2_u6_u2_n123, u2_u6_u2_n124, u2_u6_u2_n125, u2_u6_u2_n126, u2_u6_u2_n127, u2_u6_u2_n128, u2_u6_u2_n129, u2_u6_u2_n130, u2_u6_u2_n131, 
       u2_u6_u2_n132, u2_u6_u2_n133, u2_u6_u2_n134, u2_u6_u2_n135, u2_u6_u2_n136, u2_u6_u2_n137, u2_u6_u2_n138, u2_u6_u2_n139, u2_u6_u2_n140, 
       u2_u6_u2_n141, u2_u6_u2_n142, u2_u6_u2_n143, u2_u6_u2_n144, u2_u6_u2_n145, u2_u6_u2_n146, u2_u6_u2_n147, u2_u6_u2_n148, u2_u6_u2_n149, 
       u2_u6_u2_n150, u2_u6_u2_n151, u2_u6_u2_n152, u2_u6_u2_n153, u2_u6_u2_n154, u2_u6_u2_n155, u2_u6_u2_n156, u2_u6_u2_n157, u2_u6_u2_n158, 
       u2_u6_u2_n159, u2_u6_u2_n160, u2_u6_u2_n161, u2_u6_u2_n162, u2_u6_u2_n163, u2_u6_u2_n164, u2_u6_u2_n165, u2_u6_u2_n166, u2_u6_u2_n167, 
       u2_u6_u2_n168, u2_u6_u2_n169, u2_u6_u2_n170, u2_u6_u2_n171, u2_u6_u2_n172, u2_u6_u2_n173, u2_u6_u2_n174, u2_u6_u2_n175, u2_u6_u2_n176, 
       u2_u6_u2_n177, u2_u6_u2_n178, u2_u6_u2_n179, u2_u6_u2_n180, u2_u6_u2_n181, u2_u6_u2_n182, u2_u6_u2_n183, u2_u6_u2_n184, u2_u6_u2_n185, 
       u2_u6_u2_n186, u2_u6_u2_n187, u2_u6_u2_n188, u2_u6_u2_n95, u2_u6_u2_n96, u2_u6_u2_n97, u2_u6_u2_n98, u2_u6_u2_n99, u2_u6_u3_n100, 
       u2_u6_u3_n101, u2_u6_u3_n102, u2_u6_u3_n103, u2_u6_u3_n104, u2_u6_u3_n105, u2_u6_u3_n106, u2_u6_u3_n107, u2_u6_u3_n108, u2_u6_u3_n109, 
       u2_u6_u3_n110, u2_u6_u3_n111, u2_u6_u3_n112, u2_u6_u3_n113, u2_u6_u3_n114, u2_u6_u3_n115, u2_u6_u3_n116, u2_u6_u3_n117, u2_u6_u3_n118, 
       u2_u6_u3_n119, u2_u6_u3_n120, u2_u6_u3_n121, u2_u6_u3_n122, u2_u6_u3_n123, u2_u6_u3_n124, u2_u6_u3_n125, u2_u6_u3_n126, u2_u6_u3_n127, 
       u2_u6_u3_n128, u2_u6_u3_n129, u2_u6_u3_n130, u2_u6_u3_n131, u2_u6_u3_n132, u2_u6_u3_n133, u2_u6_u3_n134, u2_u6_u3_n135, u2_u6_u3_n136, 
       u2_u6_u3_n137, u2_u6_u3_n138, u2_u6_u3_n139, u2_u6_u3_n140, u2_u6_u3_n141, u2_u6_u3_n142, u2_u6_u3_n143, u2_u6_u3_n144, u2_u6_u3_n145, 
       u2_u6_u3_n146, u2_u6_u3_n147, u2_u6_u3_n148, u2_u6_u3_n149, u2_u6_u3_n150, u2_u6_u3_n151, u2_u6_u3_n152, u2_u6_u3_n153, u2_u6_u3_n154, 
       u2_u6_u3_n155, u2_u6_u3_n156, u2_u6_u3_n157, u2_u6_u3_n158, u2_u6_u3_n159, u2_u6_u3_n160, u2_u6_u3_n161, u2_u6_u3_n162, u2_u6_u3_n163, 
       u2_u6_u3_n164, u2_u6_u3_n165, u2_u6_u3_n166, u2_u6_u3_n167, u2_u6_u3_n168, u2_u6_u3_n169, u2_u6_u3_n170, u2_u6_u3_n171, u2_u6_u3_n172, 
       u2_u6_u3_n173, u2_u6_u3_n174, u2_u6_u3_n175, u2_u6_u3_n176, u2_u6_u3_n177, u2_u6_u3_n178, u2_u6_u3_n179, u2_u6_u3_n180, u2_u6_u3_n181, 
       u2_u6_u3_n182, u2_u6_u3_n183, u2_u6_u3_n184, u2_u6_u3_n185, u2_u6_u3_n186, u2_u6_u3_n94, u2_u6_u3_n95, u2_u6_u3_n96, u2_u6_u3_n97, 
       u2_u6_u3_n98, u2_u6_u3_n99, u2_u6_u4_n100, u2_u6_u4_n101, u2_u6_u4_n102, u2_u6_u4_n103, u2_u6_u4_n104, u2_u6_u4_n105, u2_u6_u4_n106, 
       u2_u6_u4_n107, u2_u6_u4_n108, u2_u6_u4_n109, u2_u6_u4_n110, u2_u6_u4_n111, u2_u6_u4_n112, u2_u6_u4_n113, u2_u6_u4_n114, u2_u6_u4_n115, 
       u2_u6_u4_n116, u2_u6_u4_n117, u2_u6_u4_n118, u2_u6_u4_n119, u2_u6_u4_n120, u2_u6_u4_n121, u2_u6_u4_n122, u2_u6_u4_n123, u2_u6_u4_n124, 
       u2_u6_u4_n125, u2_u6_u4_n126, u2_u6_u4_n127, u2_u6_u4_n128, u2_u6_u4_n129, u2_u6_u4_n130, u2_u6_u4_n131, u2_u6_u4_n132, u2_u6_u4_n133, 
       u2_u6_u4_n134, u2_u6_u4_n135, u2_u6_u4_n136, u2_u6_u4_n137, u2_u6_u4_n138, u2_u6_u4_n139, u2_u6_u4_n140, u2_u6_u4_n141, u2_u6_u4_n142, 
       u2_u6_u4_n143, u2_u6_u4_n144, u2_u6_u4_n145, u2_u6_u4_n146, u2_u6_u4_n147, u2_u6_u4_n148, u2_u6_u4_n149, u2_u6_u4_n150, u2_u6_u4_n151, 
       u2_u6_u4_n152, u2_u6_u4_n153, u2_u6_u4_n154, u2_u6_u4_n155, u2_u6_u4_n156, u2_u6_u4_n157, u2_u6_u4_n158, u2_u6_u4_n159, u2_u6_u4_n160, 
       u2_u6_u4_n161, u2_u6_u4_n162, u2_u6_u4_n163, u2_u6_u4_n164, u2_u6_u4_n165, u2_u6_u4_n166, u2_u6_u4_n167, u2_u6_u4_n168, u2_u6_u4_n169, 
       u2_u6_u4_n170, u2_u6_u4_n171, u2_u6_u4_n172, u2_u6_u4_n173, u2_u6_u4_n174, u2_u6_u4_n175, u2_u6_u4_n176, u2_u6_u4_n177, u2_u6_u4_n178, 
       u2_u6_u4_n179, u2_u6_u4_n180, u2_u6_u4_n181, u2_u6_u4_n182, u2_u6_u4_n183, u2_u6_u4_n184, u2_u6_u4_n185, u2_u6_u4_n186, u2_u6_u4_n94, 
       u2_u6_u4_n95, u2_u6_u4_n96, u2_u6_u4_n97, u2_u6_u4_n98, u2_u6_u4_n99, u2_u6_u6_n100, u2_u6_u6_n101, u2_u6_u6_n102, u2_u6_u6_n103, 
       u2_u6_u6_n104, u2_u6_u6_n105, u2_u6_u6_n106, u2_u6_u6_n107, u2_u6_u6_n108, u2_u6_u6_n109, u2_u6_u6_n110, u2_u6_u6_n111, u2_u6_u6_n112, 
       u2_u6_u6_n113, u2_u6_u6_n114, u2_u6_u6_n115, u2_u6_u6_n116, u2_u6_u6_n117, u2_u6_u6_n118, u2_u6_u6_n119, u2_u6_u6_n120, u2_u6_u6_n121, 
       u2_u6_u6_n122, u2_u6_u6_n123, u2_u6_u6_n124, u2_u6_u6_n125, u2_u6_u6_n126, u2_u6_u6_n127, u2_u6_u6_n128, u2_u6_u6_n129, u2_u6_u6_n130, 
       u2_u6_u6_n131, u2_u6_u6_n132, u2_u6_u6_n133, u2_u6_u6_n134, u2_u6_u6_n135, u2_u6_u6_n136, u2_u6_u6_n137, u2_u6_u6_n138, u2_u6_u6_n139, 
       u2_u6_u6_n140, u2_u6_u6_n141, u2_u6_u6_n142, u2_u6_u6_n143, u2_u6_u6_n144, u2_u6_u6_n145, u2_u6_u6_n146, u2_u6_u6_n147, u2_u6_u6_n148, 
       u2_u6_u6_n149, u2_u6_u6_n150, u2_u6_u6_n151, u2_u6_u6_n152, u2_u6_u6_n153, u2_u6_u6_n154, u2_u6_u6_n155, u2_u6_u6_n156, u2_u6_u6_n157, 
       u2_u6_u6_n158, u2_u6_u6_n159, u2_u6_u6_n160, u2_u6_u6_n161, u2_u6_u6_n162, u2_u6_u6_n163, u2_u6_u6_n164, u2_u6_u6_n165, u2_u6_u6_n166, 
       u2_u6_u6_n167, u2_u6_u6_n168, u2_u6_u6_n169, u2_u6_u6_n170, u2_u6_u6_n171, u2_u6_u6_n172, u2_u6_u6_n173, u2_u6_u6_n174, u2_u6_u6_n88, 
       u2_u6_u6_n89, u2_u6_u6_n90, u2_u6_u6_n91, u2_u6_u6_n92, u2_u6_u6_n93, u2_u6_u6_n94, u2_u6_u6_n95, u2_u6_u6_n96, u2_u6_u6_n97, 
       u2_u6_u6_n98, u2_u6_u6_n99, u2_u6_u7_n100, u2_u6_u7_n101, u2_u6_u7_n102, u2_u6_u7_n103, u2_u6_u7_n104, u2_u6_u7_n105, u2_u6_u7_n106, 
       u2_u6_u7_n107, u2_u6_u7_n108, u2_u6_u7_n109, u2_u6_u7_n110, u2_u6_u7_n111, u2_u6_u7_n112, u2_u6_u7_n113, u2_u6_u7_n114, u2_u6_u7_n115, 
       u2_u6_u7_n116, u2_u6_u7_n117, u2_u6_u7_n118, u2_u6_u7_n119, u2_u6_u7_n120, u2_u6_u7_n121, u2_u6_u7_n122, u2_u6_u7_n123, u2_u6_u7_n124, 
       u2_u6_u7_n125, u2_u6_u7_n126, u2_u6_u7_n127, u2_u6_u7_n128, u2_u6_u7_n129, u2_u6_u7_n130, u2_u6_u7_n131, u2_u6_u7_n132, u2_u6_u7_n133, 
       u2_u6_u7_n134, u2_u6_u7_n135, u2_u6_u7_n136, u2_u6_u7_n137, u2_u6_u7_n138, u2_u6_u7_n139, u2_u6_u7_n140, u2_u6_u7_n141, u2_u6_u7_n142, 
       u2_u6_u7_n143, u2_u6_u7_n144, u2_u6_u7_n145, u2_u6_u7_n146, u2_u6_u7_n147, u2_u6_u7_n148, u2_u6_u7_n149, u2_u6_u7_n150, u2_u6_u7_n151, 
       u2_u6_u7_n152, u2_u6_u7_n153, u2_u6_u7_n154, u2_u6_u7_n155, u2_u6_u7_n156, u2_u6_u7_n157, u2_u6_u7_n158, u2_u6_u7_n159, u2_u6_u7_n160, 
       u2_u6_u7_n161, u2_u6_u7_n162, u2_u6_u7_n163, u2_u6_u7_n164, u2_u6_u7_n165, u2_u6_u7_n166, u2_u6_u7_n167, u2_u6_u7_n168, u2_u6_u7_n169, 
       u2_u6_u7_n170, u2_u6_u7_n171, u2_u6_u7_n172, u2_u6_u7_n173, u2_u6_u7_n174, u2_u6_u7_n175, u2_u6_u7_n176, u2_u6_u7_n177, u2_u6_u7_n178, 
       u2_u6_u7_n179, u2_u6_u7_n180, u2_u6_u7_n91, u2_u6_u7_n92, u2_u6_u7_n93, u2_u6_u7_n94, u2_u6_u7_n95, u2_u6_u7_n96, u2_u6_u7_n97, 
       u2_u6_u7_n98, u2_u6_u7_n99, u2_u7_X_37, u2_u7_X_38, u2_u7_X_39, u2_u7_X_40, u2_u7_X_41, u2_u7_X_42, u2_u7_X_43, 
       u2_u7_X_44, u2_u7_X_45, u2_u7_X_46, u2_u7_X_47, u2_u7_X_48, u2_u7_u6_n100, u2_u7_u6_n101, u2_u7_u6_n102, u2_u7_u6_n103, 
       u2_u7_u6_n104, u2_u7_u6_n105, u2_u7_u6_n106, u2_u7_u6_n107, u2_u7_u6_n108, u2_u7_u6_n109, u2_u7_u6_n110, u2_u7_u6_n111, u2_u7_u6_n112, 
       u2_u7_u6_n113, u2_u7_u6_n114, u2_u7_u6_n115, u2_u7_u6_n116, u2_u7_u6_n117, u2_u7_u6_n118, u2_u7_u6_n119, u2_u7_u6_n120, u2_u7_u6_n121, 
       u2_u7_u6_n122, u2_u7_u6_n123, u2_u7_u6_n124, u2_u7_u6_n125, u2_u7_u6_n126, u2_u7_u6_n127, u2_u7_u6_n128, u2_u7_u6_n129, u2_u7_u6_n130, 
       u2_u7_u6_n131, u2_u7_u6_n132, u2_u7_u6_n133, u2_u7_u6_n134, u2_u7_u6_n135, u2_u7_u6_n136, u2_u7_u6_n137, u2_u7_u6_n138, u2_u7_u6_n139, 
       u2_u7_u6_n140, u2_u7_u6_n141, u2_u7_u6_n142, u2_u7_u6_n143, u2_u7_u6_n144, u2_u7_u6_n145, u2_u7_u6_n146, u2_u7_u6_n147, u2_u7_u6_n148, 
       u2_u7_u6_n149, u2_u7_u6_n150, u2_u7_u6_n151, u2_u7_u6_n152, u2_u7_u6_n153, u2_u7_u6_n154, u2_u7_u6_n155, u2_u7_u6_n156, u2_u7_u6_n157, 
       u2_u7_u6_n158, u2_u7_u6_n159, u2_u7_u6_n160, u2_u7_u6_n161, u2_u7_u6_n162, u2_u7_u6_n163, u2_u7_u6_n164, u2_u7_u6_n165, u2_u7_u6_n166, 
       u2_u7_u6_n167, u2_u7_u6_n168, u2_u7_u6_n169, u2_u7_u6_n170, u2_u7_u6_n171, u2_u7_u6_n172, u2_u7_u6_n173, u2_u7_u6_n174, u2_u7_u6_n88, 
       u2_u7_u6_n89, u2_u7_u6_n90, u2_u7_u6_n91, u2_u7_u6_n92, u2_u7_u6_n93, u2_u7_u6_n94, u2_u7_u6_n95, u2_u7_u6_n96, u2_u7_u6_n97, 
       u2_u7_u6_n98, u2_u7_u6_n99, u2_u7_u7_n100, u2_u7_u7_n101, u2_u7_u7_n102, u2_u7_u7_n103, u2_u7_u7_n104, u2_u7_u7_n105, u2_u7_u7_n106, 
       u2_u7_u7_n107, u2_u7_u7_n108, u2_u7_u7_n109, u2_u7_u7_n110, u2_u7_u7_n111, u2_u7_u7_n112, u2_u7_u7_n113, u2_u7_u7_n114, u2_u7_u7_n115, 
       u2_u7_u7_n116, u2_u7_u7_n117, u2_u7_u7_n118, u2_u7_u7_n119, u2_u7_u7_n120, u2_u7_u7_n121, u2_u7_u7_n122, u2_u7_u7_n123, u2_u7_u7_n124, 
       u2_u7_u7_n125, u2_u7_u7_n126, u2_u7_u7_n127, u2_u7_u7_n128, u2_u7_u7_n129, u2_u7_u7_n130, u2_u7_u7_n131, u2_u7_u7_n132, u2_u7_u7_n133, 
       u2_u7_u7_n134, u2_u7_u7_n135, u2_u7_u7_n136, u2_u7_u7_n137, u2_u7_u7_n138, u2_u7_u7_n139, u2_u7_u7_n140, u2_u7_u7_n141, u2_u7_u7_n142, 
       u2_u7_u7_n143, u2_u7_u7_n144, u2_u7_u7_n145, u2_u7_u7_n146, u2_u7_u7_n147, u2_u7_u7_n148, u2_u7_u7_n149, u2_u7_u7_n150, u2_u7_u7_n151, 
       u2_u7_u7_n152, u2_u7_u7_n153, u2_u7_u7_n154, u2_u7_u7_n155, u2_u7_u7_n156, u2_u7_u7_n157, u2_u7_u7_n158, u2_u7_u7_n159, u2_u7_u7_n160, 
       u2_u7_u7_n161, u2_u7_u7_n162, u2_u7_u7_n163, u2_u7_u7_n164, u2_u7_u7_n165, u2_u7_u7_n166, u2_u7_u7_n167, u2_u7_u7_n168, u2_u7_u7_n169, 
       u2_u7_u7_n170, u2_u7_u7_n171, u2_u7_u7_n172, u2_u7_u7_n173, u2_u7_u7_n174, u2_u7_u7_n175, u2_u7_u7_n176, u2_u7_u7_n177, u2_u7_u7_n178, 
       u2_u7_u7_n179, u2_u7_u7_n180, u2_u7_u7_n91, u2_u7_u7_n92, u2_u7_u7_n93, u2_u7_u7_n94, u2_u7_u7_n95, u2_u7_u7_n96, u2_u7_u7_n97, 
       u2_u7_u7_n98, u2_u7_u7_n99, u2_u9_X_1, u2_u9_X_10, u2_u9_X_11, u2_u9_X_12, u2_u9_X_13, u2_u9_X_14, u2_u9_X_15, 
       u2_u9_X_16, u2_u9_X_17, u2_u9_X_18, u2_u9_X_2, u2_u9_X_3, u2_u9_X_4, u2_u9_X_43, u2_u9_X_44, u2_u9_X_45, 
       u2_u9_X_46, u2_u9_X_47, u2_u9_X_48, u2_u9_X_5, u2_u9_X_6, u2_u9_X_7, u2_u9_X_8, u2_u9_X_9, u2_u9_u0_n100, 
       u2_u9_u0_n101, u2_u9_u0_n102, u2_u9_u0_n103, u2_u9_u0_n104, u2_u9_u0_n105, u2_u9_u0_n106, u2_u9_u0_n107, u2_u9_u0_n108, u2_u9_u0_n109, 
       u2_u9_u0_n110, u2_u9_u0_n111, u2_u9_u0_n112, u2_u9_u0_n113, u2_u9_u0_n114, u2_u9_u0_n115, u2_u9_u0_n116, u2_u9_u0_n117, u2_u9_u0_n118, 
       u2_u9_u0_n119, u2_u9_u0_n120, u2_u9_u0_n121, u2_u9_u0_n122, u2_u9_u0_n123, u2_u9_u0_n124, u2_u9_u0_n125, u2_u9_u0_n126, u2_u9_u0_n127, 
       u2_u9_u0_n128, u2_u9_u0_n129, u2_u9_u0_n130, u2_u9_u0_n131, u2_u9_u0_n132, u2_u9_u0_n133, u2_u9_u0_n134, u2_u9_u0_n135, u2_u9_u0_n136, 
       u2_u9_u0_n137, u2_u9_u0_n138, u2_u9_u0_n139, u2_u9_u0_n140, u2_u9_u0_n141, u2_u9_u0_n142, u2_u9_u0_n143, u2_u9_u0_n144, u2_u9_u0_n145, 
       u2_u9_u0_n146, u2_u9_u0_n147, u2_u9_u0_n148, u2_u9_u0_n149, u2_u9_u0_n150, u2_u9_u0_n151, u2_u9_u0_n152, u2_u9_u0_n153, u2_u9_u0_n154, 
       u2_u9_u0_n155, u2_u9_u0_n156, u2_u9_u0_n157, u2_u9_u0_n158, u2_u9_u0_n159, u2_u9_u0_n160, u2_u9_u0_n161, u2_u9_u0_n162, u2_u9_u0_n163, 
       u2_u9_u0_n164, u2_u9_u0_n165, u2_u9_u0_n166, u2_u9_u0_n167, u2_u9_u0_n168, u2_u9_u0_n169, u2_u9_u0_n170, u2_u9_u0_n171, u2_u9_u0_n172, 
       u2_u9_u0_n173, u2_u9_u0_n174, u2_u9_u0_n88, u2_u9_u0_n89, u2_u9_u0_n90, u2_u9_u0_n91, u2_u9_u0_n92, u2_u9_u0_n93, u2_u9_u0_n94, 
       u2_u9_u0_n95, u2_u9_u0_n96, u2_u9_u0_n97, u2_u9_u0_n98, u2_u9_u0_n99, u2_u9_u1_n100, u2_u9_u1_n101, u2_u9_u1_n102, u2_u9_u1_n103, 
       u2_u9_u1_n104, u2_u9_u1_n105, u2_u9_u1_n106, u2_u9_u1_n107, u2_u9_u1_n108, u2_u9_u1_n109, u2_u9_u1_n110, u2_u9_u1_n111, u2_u9_u1_n112, 
       u2_u9_u1_n113, u2_u9_u1_n114, u2_u9_u1_n115, u2_u9_u1_n116, u2_u9_u1_n117, u2_u9_u1_n118, u2_u9_u1_n119, u2_u9_u1_n120, u2_u9_u1_n121, 
       u2_u9_u1_n122, u2_u9_u1_n123, u2_u9_u1_n124, u2_u9_u1_n125, u2_u9_u1_n126, u2_u9_u1_n127, u2_u9_u1_n128, u2_u9_u1_n129, u2_u9_u1_n130, 
       u2_u9_u1_n131, u2_u9_u1_n132, u2_u9_u1_n133, u2_u9_u1_n134, u2_u9_u1_n135, u2_u9_u1_n136, u2_u9_u1_n137, u2_u9_u1_n138, u2_u9_u1_n139, 
       u2_u9_u1_n140, u2_u9_u1_n141, u2_u9_u1_n142, u2_u9_u1_n143, u2_u9_u1_n144, u2_u9_u1_n145, u2_u9_u1_n146, u2_u9_u1_n147, u2_u9_u1_n148, 
       u2_u9_u1_n149, u2_u9_u1_n150, u2_u9_u1_n151, u2_u9_u1_n152, u2_u9_u1_n153, u2_u9_u1_n154, u2_u9_u1_n155, u2_u9_u1_n156, u2_u9_u1_n157, 
       u2_u9_u1_n158, u2_u9_u1_n159, u2_u9_u1_n160, u2_u9_u1_n161, u2_u9_u1_n162, u2_u9_u1_n163, u2_u9_u1_n164, u2_u9_u1_n165, u2_u9_u1_n166, 
       u2_u9_u1_n167, u2_u9_u1_n168, u2_u9_u1_n169, u2_u9_u1_n170, u2_u9_u1_n171, u2_u9_u1_n172, u2_u9_u1_n173, u2_u9_u1_n174, u2_u9_u1_n175, 
       u2_u9_u1_n176, u2_u9_u1_n177, u2_u9_u1_n178, u2_u9_u1_n179, u2_u9_u1_n180, u2_u9_u1_n181, u2_u9_u1_n182, u2_u9_u1_n183, u2_u9_u1_n184, 
       u2_u9_u1_n185, u2_u9_u1_n186, u2_u9_u1_n187, u2_u9_u1_n188, u2_u9_u1_n95, u2_u9_u1_n96, u2_u9_u1_n97, u2_u9_u1_n98, u2_u9_u1_n99, 
       u2_u9_u2_n100, u2_u9_u2_n101, u2_u9_u2_n102, u2_u9_u2_n103, u2_u9_u2_n104, u2_u9_u2_n105, u2_u9_u2_n106, u2_u9_u2_n107, u2_u9_u2_n108, 
       u2_u9_u2_n109, u2_u9_u2_n110, u2_u9_u2_n111, u2_u9_u2_n112, u2_u9_u2_n113, u2_u9_u2_n114, u2_u9_u2_n115, u2_u9_u2_n116, u2_u9_u2_n117, 
       u2_u9_u2_n118, u2_u9_u2_n119, u2_u9_u2_n120, u2_u9_u2_n121, u2_u9_u2_n122, u2_u9_u2_n123, u2_u9_u2_n124, u2_u9_u2_n125, u2_u9_u2_n126, 
       u2_u9_u2_n127, u2_u9_u2_n128, u2_u9_u2_n129, u2_u9_u2_n130, u2_u9_u2_n131, u2_u9_u2_n132, u2_u9_u2_n133, u2_u9_u2_n134, u2_u9_u2_n135, 
       u2_u9_u2_n136, u2_u9_u2_n137, u2_u9_u2_n138, u2_u9_u2_n139, u2_u9_u2_n140, u2_u9_u2_n141, u2_u9_u2_n142, u2_u9_u2_n143, u2_u9_u2_n144, 
       u2_u9_u2_n145, u2_u9_u2_n146, u2_u9_u2_n147, u2_u9_u2_n148, u2_u9_u2_n149, u2_u9_u2_n150, u2_u9_u2_n151, u2_u9_u2_n152, u2_u9_u2_n153, 
       u2_u9_u2_n154, u2_u9_u2_n155, u2_u9_u2_n156, u2_u9_u2_n157, u2_u9_u2_n158, u2_u9_u2_n159, u2_u9_u2_n160, u2_u9_u2_n161, u2_u9_u2_n162, 
       u2_u9_u2_n163, u2_u9_u2_n164, u2_u9_u2_n165, u2_u9_u2_n166, u2_u9_u2_n167, u2_u9_u2_n168, u2_u9_u2_n169, u2_u9_u2_n170, u2_u9_u2_n171, 
       u2_u9_u2_n172, u2_u9_u2_n173, u2_u9_u2_n174, u2_u9_u2_n175, u2_u9_u2_n176, u2_u9_u2_n177, u2_u9_u2_n178, u2_u9_u2_n179, u2_u9_u2_n180, 
       u2_u9_u2_n181, u2_u9_u2_n182, u2_u9_u2_n183, u2_u9_u2_n184, u2_u9_u2_n185, u2_u9_u2_n186, u2_u9_u2_n187, u2_u9_u2_n188, u2_u9_u2_n95, 
       u2_u9_u2_n96, u2_u9_u2_n97, u2_u9_u2_n98, u2_u9_u2_n99, u2_u9_u7_n100, u2_u9_u7_n101, u2_u9_u7_n102, u2_u9_u7_n103, u2_u9_u7_n104, 
       u2_u9_u7_n105, u2_u9_u7_n106, u2_u9_u7_n107, u2_u9_u7_n108, u2_u9_u7_n109, u2_u9_u7_n110, u2_u9_u7_n111, u2_u9_u7_n112, u2_u9_u7_n113, 
       u2_u9_u7_n114, u2_u9_u7_n115, u2_u9_u7_n116, u2_u9_u7_n117, u2_u9_u7_n118, u2_u9_u7_n119, u2_u9_u7_n120, u2_u9_u7_n121, u2_u9_u7_n122, 
       u2_u9_u7_n123, u2_u9_u7_n124, u2_u9_u7_n125, u2_u9_u7_n126, u2_u9_u7_n127, u2_u9_u7_n128, u2_u9_u7_n129, u2_u9_u7_n130, u2_u9_u7_n131, 
       u2_u9_u7_n132, u2_u9_u7_n133, u2_u9_u7_n134, u2_u9_u7_n135, u2_u9_u7_n136, u2_u9_u7_n137, u2_u9_u7_n138, u2_u9_u7_n139, u2_u9_u7_n140, 
       u2_u9_u7_n141, u2_u9_u7_n142, u2_u9_u7_n143, u2_u9_u7_n144, u2_u9_u7_n145, u2_u9_u7_n146, u2_u9_u7_n147, u2_u9_u7_n148, u2_u9_u7_n149, 
       u2_u9_u7_n150, u2_u9_u7_n151, u2_u9_u7_n152, u2_u9_u7_n153, u2_u9_u7_n154, u2_u9_u7_n155, u2_u9_u7_n156, u2_u9_u7_n157, u2_u9_u7_n158, 
       u2_u9_u7_n159, u2_u9_u7_n160, u2_u9_u7_n161, u2_u9_u7_n162, u2_u9_u7_n163, u2_u9_u7_n164, u2_u9_u7_n165, u2_u9_u7_n166, u2_u9_u7_n167, 
       u2_u9_u7_n168, u2_u9_u7_n169, u2_u9_u7_n170, u2_u9_u7_n171, u2_u9_u7_n172, u2_u9_u7_n173, u2_u9_u7_n174, u2_u9_u7_n175, u2_u9_u7_n176, 
       u2_u9_u7_n177, u2_u9_u7_n178, u2_u9_u7_n179, u2_u9_u7_n180, u2_u9_u7_n91, u2_u9_u7_n92, u2_u9_u7_n93, u2_u9_u7_n94, u2_u9_u7_n95, 
       u2_u9_u7_n96, u2_u9_u7_n97, u2_u9_u7_n98, u2_u9_u7_n99, u2_uk_n1008, u2_uk_n1013, u2_uk_n1014, u2_uk_n1015, u2_uk_n1016, 
       u2_uk_n1017, u2_uk_n1019, u2_uk_n1021, u2_uk_n1026, u2_uk_n1029, u2_uk_n1030, u2_uk_n1032, u2_uk_n1033, u2_uk_n1041, 
       u2_uk_n1057, u2_uk_n1062, u2_uk_n1064, u2_uk_n1065, u2_uk_n1075, u2_uk_n1076, u2_uk_n1078, u2_uk_n1080, u2_uk_n1083, 
       u2_uk_n1084, u2_uk_n1085, u2_uk_n1086, u2_uk_n1095, u2_uk_n1108, u2_uk_n1109, u2_uk_n1114, u2_uk_n1115, u2_uk_n1153, 
       u2_uk_n1154, u2_uk_n1159, u2_uk_n1160, u2_uk_n1174, u2_uk_n1175, u2_uk_n1184, u2_uk_n242, u2_uk_n250, u2_uk_n286, 
       u2_uk_n308, u2_uk_n409, u2_uk_n515, u2_uk_n518, u2_uk_n688, u2_uk_n692, u2_uk_n694, u2_uk_n934, u2_uk_n935, 
       u2_uk_n938, u2_uk_n940, u2_uk_n946, u2_uk_n957, u2_uk_n958, u2_uk_n959, u2_uk_n960, u2_uk_n963, u2_uk_n965, 
       u2_uk_n966, u2_uk_n968, u2_uk_n969, u2_uk_n971, u2_uk_n973, u2_uk_n974, u2_uk_n978, u2_uk_n990,  u2_uk_n998;
  XOR2_X1 u0_U101 (.B( u0_L12_26 ) , .Z( u0_N441 ) , .A( u0_out13_26 ) );
  XOR2_X1 u0_U102 (.B( u0_L12_25 ) , .Z( u0_N440 ) , .A( u0_out13_25 ) );
  XOR2_X1 u0_U104 (.B( u0_L12_24 ) , .Z( u0_N439 ) , .A( u0_out13_24 ) );
  XOR2_X1 u0_U105 (.B( u0_L12_23 ) , .Z( u0_N438 ) , .A( u0_out13_23 ) );
  XOR2_X1 u0_U108 (.B( u0_L12_20 ) , .Z( u0_N435 ) , .A( u0_out13_20 ) );
  XOR2_X1 u0_U109 (.B( u0_L12_19 ) , .Z( u0_N434 ) , .A( u0_out13_19 ) );
  XOR2_X1 u0_U110 (.B( u0_L12_18 ) , .Z( u0_N433 ) , .A( u0_out13_18 ) );
  XOR2_X1 u0_U111 (.B( u0_L12_17 ) , .Z( u0_N432 ) , .A( u0_out13_17 ) );
  XOR2_X1 u0_U112 (.B( u0_L12_16 ) , .Z( u0_N431 ) , .A( u0_out13_16 ) );
  XOR2_X1 u0_U115 (.B( u0_L12_14 ) , .Z( u0_N429 ) , .A( u0_out13_14 ) );
  XOR2_X1 u0_U116 (.B( u0_L12_13 ) , .Z( u0_N428 ) , .A( u0_out13_13 ) );
  XOR2_X1 u0_U118 (.B( u0_L12_11 ) , .Z( u0_N426 ) , .A( u0_out13_11 ) );
  XOR2_X1 u0_U119 (.B( u0_L12_10 ) , .Z( u0_N425 ) , .A( u0_out13_10 ) );
  XOR2_X1 u0_U120 (.B( u0_L12_9 ) , .Z( u0_N424 ) , .A( u0_out13_9 ) );
  XOR2_X1 u0_U121 (.B( u0_L12_8 ) , .Z( u0_N423 ) , .A( u0_out13_8 ) );
  XOR2_X1 u0_U123 (.B( u0_L12_6 ) , .Z( u0_N421 ) , .A( u0_out13_6 ) );
  XOR2_X1 u0_U126 (.B( u0_L12_4 ) , .Z( u0_N419 ) , .A( u0_out13_4 ) );
  XOR2_X1 u0_U127 (.B( u0_L12_3 ) , .Z( u0_N418 ) , .A( u0_out13_3 ) );
  XOR2_X1 u0_U128 (.B( u0_L12_2 ) , .Z( u0_N417 ) , .A( u0_out13_2 ) );
  XOR2_X1 u0_U129 (.B( u0_L12_1 ) , .Z( u0_N416 ) , .A( u0_out13_1 ) );
  XOR2_X1 u0_U13 (.Z( u0_N9 ) , .B( u0_desIn_r_12 ) , .A( u0_out0_10 ) );
  XOR2_X1 u0_U24 (.Z( u0_N8 ) , .B( u0_desIn_r_4 ) , .A( u0_out0_9 ) );
  XOR2_X1 u0_U258 (.Z( u0_N30 ) , .B( u0_desIn_r_48 ) , .A( u0_out0_31 ) );
  XOR2_X1 u0_U270 (.Z( u0_N29 ) , .B( u0_desIn_r_40 ) , .A( u0_out0_30 ) );
  XOR2_X1 u0_U292 (.Z( u0_N27 ) , .B( u0_desIn_r_24 ) , .A( u0_out0_28 ) );
  XOR2_X1 u0_U314 (.Z( u0_N25 ) , .B( u0_desIn_r_8 ) , .A( u0_out0_26 ) );
  XOR2_X1 u0_U336 (.Z( u0_N23 ) , .B( u0_desIn_r_58 ) , .A( u0_out0_24 ) );
  XOR2_X1 u0_U347 (.Z( u0_N22 ) , .B( u0_desIn_r_50 ) , .A( u0_out0_23 ) );
  XOR2_X1 u0_U381 (.Z( u0_N19 ) , .B( u0_desIn_r_26 ) , .A( u0_out0_20 ) );
  XOR2_X1 u0_U403 (.Z( u0_N17 ) , .B( u0_desIn_r_10 ) , .A( u0_out0_18 ) );
  XOR2_X1 u0_U414 (.Z( u0_N16 ) , .B( u0_desIn_r_2 ) , .A( u0_out0_17 ) );
  XOR2_X1 u0_U417 (.B( u0_L3_30 ) , .Z( u0_N157 ) , .A( u0_out4_30 ) );
  XOR2_X1 u0_U419 (.B( u0_L3_28 ) , .Z( u0_N155 ) , .A( u0_out4_28 ) );
  XOR2_X1 u0_U421 (.B( u0_L3_26 ) , .Z( u0_N153 ) , .A( u0_out4_26 ) );
  XOR2_X1 u0_U423 (.B( u0_L3_24 ) , .Z( u0_N151 ) , .A( u0_out4_24 ) );
  XOR2_X1 u0_U425 (.Z( u0_N15 ) , .B( u0_desIn_r_60 ) , .A( u0_out0_16 ) );
  XOR2_X1 u0_U428 (.B( u0_L3_20 ) , .Z( u0_N147 ) , .A( u0_out4_20 ) );
  XOR2_X1 u0_U430 (.B( u0_L3_18 ) , .Z( u0_N145 ) , .A( u0_out4_18 ) );
  XOR2_X1 u0_U432 (.B( u0_L3_16 ) , .Z( u0_N143 ) , .A( u0_out4_16 ) );
  XOR2_X1 u0_U435 (.B( u0_L3_13 ) , .Z( u0_N140 ) , .A( u0_out4_13 ) );
  XOR2_X1 u0_U439 (.B( u0_L3_10 ) , .Z( u0_N137 ) , .A( u0_out4_10 ) );
  XOR2_X1 u0_U443 (.B( u0_L3_6 ) , .Z( u0_N133 ) , .A( u0_out4_6 ) );
  XOR2_X1 u0_U448 (.B( u0_L3_2 ) , .Z( u0_N129 ) , .A( u0_out4_2 ) );
  XOR2_X1 u0_U449 (.B( u0_L3_1 ) , .Z( u0_N128 ) , .A( u0_out4_1 ) );
  XOR2_X1 u0_U458 (.Z( u0_N12 ) , .B( u0_desIn_r_36 ) , .A( u0_out0_13 ) );
  XOR2_X1 u0_U481 (.Z( u0_N1 ) , .B( u0_desIn_r_14 ) , .A( u0_out0_2 ) );
  XOR2_X1 u0_U482 (.Z( u0_N0 ) , .B( u0_desIn_r_6 ) , .A( u0_out0_1 ) );
  XOR2_X1 u0_U57 (.Z( u0_N5 ) , .B( u0_desIn_r_46 ) , .A( u0_out0_6 ) );
  XOR2_X1 u0_U96 (.B( u0_L12_31 ) , .Z( u0_N446 ) , .A( u0_out13_31 ) );
  XOR2_X1 u0_U97 (.B( u0_L12_30 ) , .Z( u0_N445 ) , .A( u0_out13_30 ) );
  XOR2_X1 u0_U98 (.B( u0_L12_29 ) , .Z( u0_N444 ) , .A( u0_out13_29 ) );
  XOR2_X1 u0_U99 (.B( u0_L12_28 ) , .Z( u0_N443 ) , .A( u0_out13_28 ) );
  XOR2_X1 u0_u0_U1 (.B( u0_K1_9 ) , .A( u0_desIn_r_47 ) , .Z( u0_u0_X_9 ) );
  XOR2_X1 u0_u0_U16 (.B( u0_K1_3 ) , .A( u0_desIn_r_15 ) , .Z( u0_u0_X_3 ) );
  XOR2_X1 u0_u0_U2 (.B( u0_K1_8 ) , .A( u0_desIn_r_39 ) , .Z( u0_u0_X_8 ) );
  XOR2_X1 u0_u0_U27 (.B( u0_K1_2 ) , .A( u0_desIn_r_7 ) , .Z( u0_u0_X_2 ) );
  XOR2_X1 u0_u0_U3 (.B( u0_K1_7 ) , .A( u0_desIn_r_31 ) , .Z( u0_u0_X_7 ) );
  XOR2_X1 u0_u0_U33 (.B( u0_K1_24 ) , .A( u0_desIn_r_3 ) , .Z( u0_u0_X_24 ) );
  XOR2_X1 u0_u0_U34 (.B( u0_K1_23 ) , .A( u0_desIn_r_61 ) , .Z( u0_u0_X_23 ) );
  XOR2_X1 u0_u0_U35 (.B( u0_K1_22 ) , .A( u0_desIn_r_53 ) , .Z( u0_u0_X_22 ) );
  XOR2_X1 u0_u0_U36 (.B( u0_K1_21 ) , .A( u0_desIn_r_45 ) , .Z( u0_u0_X_21 ) );
  XOR2_X1 u0_u0_U37 (.B( u0_K1_20 ) , .A( u0_desIn_r_37 ) , .Z( u0_u0_X_20 ) );
  XOR2_X1 u0_u0_U38 (.B( u0_K1_1 ) , .A( u0_desIn_r_57 ) , .Z( u0_u0_X_1 ) );
  XOR2_X1 u0_u0_U39 (.B( u0_K1_19 ) , .A( u0_desIn_r_29 ) , .Z( u0_u0_X_19 ) );
  XOR2_X1 u0_u0_U4 (.B( u0_K1_6 ) , .A( u0_desIn_r_39 ) , .Z( u0_u0_X_6 ) );
  XOR2_X1 u0_u0_U40 (.B( u0_K1_18 ) , .A( u0_desIn_r_37 ) , .Z( u0_u0_X_18 ) );
  XOR2_X1 u0_u0_U41 (.B( u0_K1_17 ) , .A( u0_desIn_r_29 ) , .Z( u0_u0_X_17 ) );
  XOR2_X1 u0_u0_U42 (.B( u0_K1_16 ) , .A( u0_desIn_r_21 ) , .Z( u0_u0_X_16 ) );
  XOR2_X1 u0_u0_U43 (.B( u0_K1_15 ) , .A( u0_desIn_r_13 ) , .Z( u0_u0_X_15 ) );
  XOR2_X1 u0_u0_U44 (.B( u0_K1_14 ) , .A( u0_desIn_r_5 ) , .Z( u0_u0_X_14 ) );
  XOR2_X1 u0_u0_U45 (.B( u0_K1_13 ) , .A( u0_desIn_r_63 ) , .Z( u0_u0_X_13 ) );
  XOR2_X1 u0_u0_U46 (.B( u0_K1_12 ) , .A( u0_desIn_r_5 ) , .Z( u0_u0_X_12 ) );
  XOR2_X1 u0_u0_U47 (.B( u0_K1_11 ) , .A( u0_desIn_r_63 ) , .Z( u0_u0_X_11 ) );
  XOR2_X1 u0_u0_U48 (.B( u0_K1_10 ) , .A( u0_desIn_r_55 ) , .Z( u0_u0_X_10 ) );
  XOR2_X1 u0_u0_U5 (.B( u0_K1_5 ) , .A( u0_desIn_r_31 ) , .Z( u0_u0_X_5 ) );
  XOR2_X1 u0_u0_U6 (.B( u0_K1_4 ) , .A( u0_desIn_r_23 ) , .Z( u0_u0_X_4 ) );
  AND3_X1 u0_u0_u0_U10 (.A1( u0_u0_u0_n27 ) , .A3( u0_u0_u0_n45 ) , .ZN( u0_u0_u0_n48 ) , .A2( u0_u0_u0_n63 ) );
  NAND2_X1 u0_u0_u0_U11 (.A2( u0_u0_u0_n26 ) , .A1( u0_u0_u0_n36 ) , .ZN( u0_u0_u0_n62 ) );
  AND2_X1 u0_u0_u0_U12 (.A2( u0_u0_u0_n35 ) , .A1( u0_u0_u0_n45 ) , .ZN( u0_u0_u0_n68 ) );
  AND2_X1 u0_u0_u0_U13 (.ZN( u0_u0_u0_n24 ) , .A1( u0_u0_u0_n45 ) , .A2( u0_u0_u0_n46 ) );
  AND2_X1 u0_u0_u0_U14 (.ZN( u0_u0_u0_n30 ) , .A2( u0_u0_u0_n50 ) , .A1( u0_u0_u0_n67 ) );
  INV_X1 u0_u0_u0_U15 (.ZN( u0_u0_u0_n2 ) , .A( u0_u0_u0_n32 ) );
  NOR2_X1 u0_u0_u0_U16 (.A1( u0_u0_u0_n15 ) , .ZN( u0_u0_u0_n28 ) , .A2( u0_u0_u0_n39 ) );
  AOI21_X1 u0_u0_u0_U17 (.A( u0_u0_u0_n10 ) , .ZN( u0_u0_u0_n43 ) , .B1( u0_u0_u0_n72 ) , .B2( u0_u0_u0_n82 ) );
  INV_X1 u0_u0_u0_U18 (.ZN( u0_u0_u0_n10 ) , .A( u0_u0_u0_n33 ) );
  OAI22_X1 u0_u0_u0_U19 (.B2( u0_u0_u0_n28 ) , .A2( u0_u0_u0_n29 ) , .A1( u0_u0_u0_n37 ) , .ZN( u0_u0_u0_n49 ) , .B1( u0_u0_u0_n50 ) );
  OAI22_X1 u0_u0_u0_U20 (.B2( u0_u0_u0_n28 ) , .A1( u0_u0_u0_n31 ) , .B1( u0_u0_u0_n44 ) , .ZN( u0_u0_u0_n84 ) , .A2( u0_u0_u0_n85 ) );
  AND3_X1 u0_u0_u0_U21 (.A1( u0_u0_u0_n27 ) , .A2( u0_u0_u0_n50 ) , .A3( u0_u0_u0_n54 ) , .ZN( u0_u0_u0_n85 ) );
  NAND2_X1 u0_u0_u0_U22 (.ZN( u0_u0_u0_n50 ) , .A2( u0_u0_u0_n72 ) , .A1( u0_u0_u0_n75 ) );
  INV_X1 u0_u0_u0_U23 (.ZN( u0_u0_u0_n14 ) , .A( u0_u0_u0_n39 ) );
  AOI22_X1 u0_u0_u0_U24 (.A1( u0_u0_u0_n15 ) , .B1( u0_u0_u0_n57 ) , .ZN( u0_u0_u0_n64 ) , .A2( u0_u0_u0_n65 ) , .B2( u0_u0_u0_n66 ) );
  NAND2_X1 u0_u0_u0_U25 (.ZN( u0_u0_u0_n46 ) , .A1( u0_u0_u0_n75 ) , .A2( u0_u0_u0_n80 ) );
  INV_X1 u0_u0_u0_U26 (.ZN( u0_u0_u0_n17 ) , .A( u0_u0_u0_n57 ) );
  AOI21_X1 u0_u0_u0_U27 (.A( u0_u0_u0_n31 ) , .B2( u0_u0_u0_n34 ) , .B1( u0_u0_u0_n68 ) , .ZN( u0_u0_u0_n71 ) );
  AOI21_X1 u0_u0_u0_U28 (.A( u0_u0_u0_n37 ) , .B2( u0_u0_u0_n46 ) , .B1( u0_u0_u0_n48 ) , .ZN( u0_u0_u0_n79 ) );
  AOI21_X1 u0_u0_u0_U29 (.A( u0_u0_u0_n31 ) , .B2( u0_u0_u0_n33 ) , .ZN( u0_u0_u0_n59 ) , .B1( u0_u0_u0_n9 ) );
  INV_X1 u0_u0_u0_U3 (.A( u0_u0_u0_n62 ) , .ZN( u0_u0_u0_n9 ) );
  NOR2_X1 u0_u0_u0_U30 (.ZN( u0_u0_u0_n32 ) , .A1( u0_u0_u0_n55 ) , .A2( u0_u0_u0_n8 ) );
  OAI221_X1 u0_u0_u0_U31 (.C2( u0_u0_u0_n28 ) , .A( u0_u0_u0_n3 ) , .B2( u0_u0_u0_n34 ) , .B1( u0_u0_u0_n37 ) , .ZN( u0_u0_u0_n55 ) , .C1( u0_u0_u0_n63 ) );
  AOI211_X1 u0_u0_u0_U32 (.ZN( u0_u0_u0_n56 ) , .C1( u0_u0_u0_n57 ) , .C2( u0_u0_u0_n58 ) , .A( u0_u0_u0_n59 ) , .B( u0_u0_u0_n60 ) );
  NAND2_X1 u0_u0_u0_U33 (.ZN( u0_u0_u0_n47 ) , .A1( u0_u0_u0_n73 ) , .A2( u0_u0_u0_n80 ) );
  NAND2_X1 u0_u0_u0_U34 (.ZN( u0_u0_u0_n36 ) , .A1( u0_u0_u0_n74 ) , .A2( u0_u0_u0_n75 ) );
  NAND2_X1 u0_u0_u0_U35 (.ZN( u0_u0_u0_n27 ) , .A2( u0_u0_u0_n80 ) , .A1( u0_u0_u0_n82 ) );
  NAND2_X1 u0_u0_u0_U36 (.ZN( u0_u0_u0_n44 ) , .A2( u0_u0_u0_n75 ) , .A1( u0_u0_u0_n83 ) );
  NAND2_X1 u0_u0_u0_U37 (.ZN( u0_u0_u0_n25 ) , .A2( u0_u0_u0_n73 ) , .A1( u0_u0_u0_n74 ) );
  INV_X1 u0_u0_u0_U38 (.ZN( u0_u0_u0_n15 ) , .A( u0_u0_u0_n37 ) );
  NAND2_X1 u0_u0_u0_U39 (.ZN( u0_u0_u0_n26 ) , .A1( u0_u0_u0_n72 ) , .A2( u0_u0_u0_n73 ) );
  AOI21_X1 u0_u0_u0_U4 (.A( u0_u0_u0_n14 ) , .B2( u0_u0_u0_n46 ) , .ZN( u0_u0_u0_n60 ) , .B1( u0_u0_u0_n61 ) );
  NAND2_X1 u0_u0_u0_U40 (.ZN( u0_u0_u0_n61 ) , .A2( u0_u0_u0_n73 ) , .A1( u0_u0_u0_n83 ) );
  INV_X1 u0_u0_u0_U41 (.ZN( u0_u0_u0_n3 ) , .A( u0_u0_u0_n87 ) );
  OAI222_X1 u0_u0_u0_U42 (.C2( u0_u0_u0_n14 ) , .A2( u0_u0_u0_n17 ) , .B1( u0_u0_u0_n31 ) , .B2( u0_u0_u0_n47 ) , .A1( u0_u0_u0_n50 ) , .C1( u0_u0_u0_n67 ) , .ZN( u0_u0_u0_n87 ) );
  NAND2_X1 u0_u0_u0_U43 (.ZN( u0_u0_u0_n54 ) , .A2( u0_u0_u0_n74 ) , .A1( u0_u0_u0_n82 ) );
  NAND2_X1 u0_u0_u0_U44 (.ZN( u0_u0_u0_n63 ) , .A1( u0_u0_u0_n82 ) , .A2( u0_u0_u0_n83 ) );
  OR3_X1 u0_u0_u0_U45 (.ZN( u0_u0_u0_n20 ) , .A1( u0_u0_u0_n21 ) , .A2( u0_u0_u0_n22 ) , .A3( u0_u0_u0_n23 ) );
  AOI21_X1 u0_u0_u0_U46 (.A( u0_u0_u0_n17 ) , .ZN( u0_u0_u0_n23 ) , .B1( u0_u0_u0_n24 ) , .B2( u0_u0_u0_n25 ) );
  AOI21_X1 u0_u0_u0_U47 (.ZN( u0_u0_u0_n21 ) , .B1( u0_u0_u0_n29 ) , .B2( u0_u0_u0_n30 ) , .A( u0_u0_u0_n31 ) );
  AOI21_X1 u0_u0_u0_U48 (.ZN( u0_u0_u0_n22 ) , .B1( u0_u0_u0_n26 ) , .B2( u0_u0_u0_n27 ) , .A( u0_u0_u0_n28 ) );
  INV_X1 u0_u0_u0_U49 (.ZN( u0_u0_u0_n4 ) , .A( u0_u0_u0_n76 ) );
  AOI21_X1 u0_u0_u0_U5 (.A( u0_u0_u0_n17 ) , .B1( u0_u0_u0_n24 ) , .ZN( u0_u0_u0_n41 ) , .B2( u0_u0_u0_n44 ) );
  OAI211_X1 u0_u0_u0_U50 (.C1( u0_u0_u0_n14 ) , .C2( u0_u0_u0_n35 ) , .A( u0_u0_u0_n6 ) , .ZN( u0_u0_u0_n76 ) , .B( u0_u0_u0_n77 ) );
  INV_X1 u0_u0_u0_U51 (.ZN( u0_u0_u0_n6 ) , .A( u0_u0_u0_n84 ) );
  AOI211_X1 u0_u0_u0_U52 (.A( u0_u0_u0_n52 ) , .C1( u0_u0_u0_n57 ) , .ZN( u0_u0_u0_n77 ) , .C2( u0_u0_u0_n78 ) , .B( u0_u0_u0_n79 ) );
  NOR2_X1 u0_u0_u0_U53 (.A2( u0_u0_X_4 ) , .A1( u0_u0_X_5 ) , .ZN( u0_u0_u0_n57 ) );
  NOR2_X1 u0_u0_u0_U54 (.A2( u0_u0_X_2 ) , .A1( u0_u0_u0_n11 ) , .ZN( u0_u0_u0_n72 ) );
  NOR2_X1 u0_u0_u0_U55 (.A2( u0_u0_X_1 ) , .A1( u0_u0_X_2 ) , .ZN( u0_u0_u0_n83 ) );
  NOR2_X1 u0_u0_u0_U56 (.A2( u0_u0_X_1 ) , .A1( u0_u0_u0_n12 ) , .ZN( u0_u0_u0_n74 ) );
  NAND2_X1 u0_u0_u0_U57 (.A2( u0_u0_X_4 ) , .A1( u0_u0_X_5 ) , .ZN( u0_u0_u0_n31 ) );
  NOR2_X1 u0_u0_u0_U58 (.A2( u0_u0_X_5 ) , .A1( u0_u0_u0_n16 ) , .ZN( u0_u0_u0_n39 ) );
  NAND2_X1 u0_u0_u0_U59 (.A1( u0_u0_X_5 ) , .A2( u0_u0_u0_n16 ) , .ZN( u0_u0_u0_n37 ) );
  NOR2_X1 u0_u0_u0_U6 (.A2( u0_u0_u0_n17 ) , .ZN( u0_u0_u0_n52 ) , .A1( u0_u0_u0_n67 ) );
  AND2_X1 u0_u0_u0_U60 (.A2( u0_u0_X_3 ) , .A1( u0_u0_X_6 ) , .ZN( u0_u0_u0_n73 ) );
  AND2_X1 u0_u0_u0_U61 (.A1( u0_u0_X_6 ) , .A2( u0_u0_u0_n13 ) , .ZN( u0_u0_u0_n82 ) );
  INV_X1 u0_u0_u0_U62 (.A( u0_u0_X_4 ) , .ZN( u0_u0_u0_n16 ) );
  INV_X1 u0_u0_u0_U63 (.A( u0_u0_X_2 ) , .ZN( u0_u0_u0_n12 ) );
  INV_X1 u0_u0_u0_U64 (.A( u0_u0_X_3 ) , .ZN( u0_u0_u0_n13 ) );
  AOI211_X1 u0_u0_u0_U65 (.C1( u0_u0_u0_n15 ) , .C2( u0_u0_u0_n62 ) , .ZN( u0_u0_u0_n69 ) , .A( u0_u0_u0_n70 ) , .B( u0_u0_u0_n71 ) );
  INV_X1 u0_u0_u0_U66 (.ZN( u0_u0_u0_n1 ) , .A( u0_u0_u0_n86 ) );
  OR4_X1 u0_u0_u0_U67 (.ZN( u0_out0_17 ) , .A3( u0_u0_u0_n5 ) , .A1( u0_u0_u0_n51 ) , .A2( u0_u0_u0_n52 ) , .A4( u0_u0_u0_n53 ) );
  AOI21_X1 u0_u0_u0_U68 (.A( u0_u0_u0_n14 ) , .B1( u0_u0_u0_n47 ) , .ZN( u0_u0_u0_n51 ) , .B2( u0_u0_u0_n68 ) );
  INV_X1 u0_u0_u0_U69 (.ZN( u0_u0_u0_n5 ) , .A( u0_u0_u0_n64 ) );
  OAI21_X1 u0_u0_u0_U7 (.B2( u0_u0_u0_n17 ) , .B1( u0_u0_u0_n25 ) , .A( u0_u0_u0_n3 ) , .ZN( u0_u0_u0_n86 ) );
  OR4_X1 u0_u0_u0_U70 (.ZN( u0_out0_31 ) , .A1( u0_u0_u0_n18 ) , .A2( u0_u0_u0_n19 ) , .A3( u0_u0_u0_n2 ) , .A4( u0_u0_u0_n20 ) );
  AOI21_X1 u0_u0_u0_U71 (.ZN( u0_u0_u0_n18 ) , .B1( u0_u0_u0_n35 ) , .B2( u0_u0_u0_n36 ) , .A( u0_u0_u0_n37 ) );
  AOI21_X1 u0_u0_u0_U72 (.A( u0_u0_u0_n14 ) , .ZN( u0_u0_u0_n19 ) , .B1( u0_u0_u0_n33 ) , .B2( u0_u0_u0_n34 ) );
  INV_X1 u0_u0_u0_U73 (.A( u0_u0_u0_n49 ) , .ZN( u0_u0_u0_n7 ) );
  AOI211_X1 u0_u0_u0_U74 (.ZN( u0_u0_u0_n38 ) , .C1( u0_u0_u0_n39 ) , .C2( u0_u0_u0_n40 ) , .A( u0_u0_u0_n41 ) , .B( u0_u0_u0_n42 ) );
  NOR2_X1 u0_u0_u0_U75 (.A2( u0_u0_u0_n11 ) , .A1( u0_u0_u0_n12 ) , .ZN( u0_u0_u0_n80 ) );
  OAI221_X1 u0_u0_u0_U76 (.C2( u0_u0_u0_n28 ) , .B1( u0_u0_u0_n31 ) , .A( u0_u0_u0_n32 ) , .B2( u0_u0_u0_n48 ) , .ZN( u0_u0_u0_n53 ) , .C1( u0_u0_u0_n54 ) );
  INV_X1 u0_u0_u0_U77 (.A( u0_u0_X_1 ) , .ZN( u0_u0_u0_n11 ) );
  AOI21_X1 u0_u0_u0_U78 (.A( u0_u0_u0_n31 ) , .ZN( u0_u0_u0_n42 ) , .B1( u0_u0_u0_n43 ) , .B2( u0_u0_u0_n9 ) );
  OAI22_X1 u0_u0_u0_U79 (.B2( u0_u0_u0_n14 ) , .A1( u0_u0_u0_n28 ) , .B1( u0_u0_u0_n29 ) , .A2( u0_u0_u0_n43 ) , .ZN( u0_u0_u0_n70 ) );
  AND2_X1 u0_u0_u0_U8 (.ZN( u0_u0_u0_n29 ) , .A2( u0_u0_u0_n54 ) , .A1( u0_u0_u0_n61 ) );
  NAND2_X1 u0_u0_u0_U80 (.A1( u0_u0_u0_n30 ) , .A2( u0_u0_u0_n43 ) , .ZN( u0_u0_u0_n65 ) );
  INV_X1 u0_u0_u0_U81 (.A( u0_u0_u0_n56 ) , .ZN( u0_u0_u0_n8 ) );
  NAND2_X1 u0_u0_u0_U82 (.ZN( u0_u0_u0_n35 ) , .A2( u0_u0_u0_n72 ) , .A1( u0_u0_u0_n81 ) );
  NAND2_X1 u0_u0_u0_U83 (.ZN( u0_u0_u0_n45 ) , .A1( u0_u0_u0_n74 ) , .A2( u0_u0_u0_n81 ) );
  NAND2_X1 u0_u0_u0_U84 (.ZN( u0_u0_u0_n67 ) , .A2( u0_u0_u0_n81 ) , .A1( u0_u0_u0_n83 ) );
  NAND2_X1 u0_u0_u0_U85 (.ZN( u0_u0_u0_n33 ) , .A2( u0_u0_u0_n80 ) , .A1( u0_u0_u0_n81 ) );
  NOR2_X1 u0_u0_u0_U86 (.A2( u0_u0_X_6 ) , .A1( u0_u0_u0_n13 ) , .ZN( u0_u0_u0_n75 ) );
  NOR2_X1 u0_u0_u0_U87 (.A2( u0_u0_X_3 ) , .A1( u0_u0_X_6 ) , .ZN( u0_u0_u0_n81 ) );
  NAND3_X1 u0_u0_u0_U88 (.ZN( u0_out0_23 ) , .A3( u0_u0_u0_n38 ) , .A2( u0_u0_u0_n4 ) , .A1( u0_u0_u0_n7 ) );
  NAND3_X1 u0_u0_u0_U89 (.A1( u0_u0_u0_n25 ) , .ZN( u0_u0_u0_n40 ) , .A2( u0_u0_u0_n47 ) , .A3( u0_u0_u0_n48 ) );
  AND2_X1 u0_u0_u0_U9 (.A2( u0_u0_u0_n25 ) , .ZN( u0_u0_u0_n34 ) , .A1( u0_u0_u0_n44 ) );
  NAND3_X1 u0_u0_u0_U90 (.A1( u0_u0_u0_n27 ) , .A2( u0_u0_u0_n36 ) , .A3( u0_u0_u0_n43 ) , .ZN( u0_u0_u0_n58 ) );
  NAND3_X1 u0_u0_u0_U91 (.A1( u0_u0_u0_n26 ) , .A3( u0_u0_u0_n35 ) , .A2( u0_u0_u0_n61 ) , .ZN( u0_u0_u0_n66 ) );
  NAND3_X1 u0_u0_u0_U92 (.ZN( u0_out0_9 ) , .A1( u0_u0_u0_n1 ) , .A2( u0_u0_u0_n4 ) , .A3( u0_u0_u0_n69 ) );
  NAND3_X1 u0_u0_u0_U93 (.A3( u0_u0_u0_n29 ) , .A1( u0_u0_u0_n43 ) , .A2( u0_u0_u0_n47 ) , .ZN( u0_u0_u0_n78 ) );
  AOI21_X1 u0_u0_u1_U10 (.A( u0_u0_u1_n15 ) , .ZN( u0_u0_u1_n32 ) , .B1( u0_u0_u1_n33 ) , .B2( u0_u0_u1_n34 ) );
  NAND3_X1 u0_u0_u1_U100 (.A2( u0_u0_u1_n34 ) , .A3( u0_u0_u1_n56 ) , .A1( u0_u0_u1_n69 ) , .ZN( u0_u0_u1_n76 ) );
  NAND2_X1 u0_u0_u1_U11 (.A1( u0_u0_u1_n34 ) , .A2( u0_u0_u1_n39 ) , .ZN( u0_u0_u1_n49 ) );
  NAND2_X1 u0_u0_u1_U12 (.A2( u0_u0_u1_n36 ) , .ZN( u0_u0_u1_n42 ) , .A1( u0_u0_u1_n58 ) );
  AOI22_X1 u0_u0_u1_U13 (.B1( u0_u0_u1_n16 ) , .A1( u0_u0_u1_n18 ) , .ZN( u0_u0_u1_n46 ) , .A2( u0_u0_u1_n52 ) , .B2( u0_u0_u1_n53 ) );
  INV_X1 u0_u0_u1_U14 (.A( u0_u0_u1_n42 ) , .ZN( u0_u0_u1_n8 ) );
  INV_X1 u0_u0_u1_U15 (.ZN( u0_u0_u1_n15 ) , .A( u0_u0_u1_n50 ) );
  OR4_X1 u0_u0_u1_U16 (.A2( u0_u0_u1_n5 ) , .A1( u0_u0_u1_n72 ) , .ZN( u0_u0_u1_n81 ) , .A3( u0_u0_u1_n82 ) , .A4( u0_u0_u1_n83 ) );
  AOI21_X1 u0_u0_u1_U17 (.B2( u0_u0_u1_n33 ) , .B1( u0_u0_u1_n35 ) , .A( u0_u0_u1_n77 ) , .ZN( u0_u0_u1_n83 ) );
  AOI21_X1 u0_u0_u1_U18 (.A( u0_u0_u1_n15 ) , .B2( u0_u0_u1_n40 ) , .B1( u0_u0_u1_n55 ) , .ZN( u0_u0_u1_n82 ) );
  INV_X1 u0_u0_u1_U19 (.ZN( u0_u0_u1_n5 ) , .A( u0_u0_u1_n88 ) );
  INV_X1 u0_u0_u1_U20 (.ZN( u0_u0_u1_n18 ) , .A( u0_u0_u1_n77 ) );
  NAND2_X1 u0_u0_u1_U21 (.A2( u0_u0_u1_n33 ) , .A1( u0_u0_u1_n36 ) , .ZN( u0_u0_u1_n48 ) );
  AND2_X1 u0_u0_u1_U22 (.A2( u0_u0_u1_n28 ) , .ZN( u0_u0_u1_n55 ) , .A1( u0_u0_u1_n66 ) );
  NAND2_X1 u0_u0_u1_U23 (.ZN( u0_u0_u1_n41 ) , .A1( u0_u0_u1_n73 ) , .A2( u0_u0_u1_n74 ) );
  NAND2_X1 u0_u0_u1_U24 (.ZN( u0_u0_u1_n30 ) , .A1( u0_u0_u1_n54 ) , .A2( u0_u0_u1_n56 ) );
  NAND2_X1 u0_u0_u1_U25 (.ZN( u0_u0_u1_n57 ) , .A1( u0_u0_u1_n69 ) , .A2( u0_u0_u1_n74 ) );
  INV_X1 u0_u0_u1_U26 (.ZN( u0_u0_u1_n11 ) , .A( u0_u0_u1_n35 ) );
  INV_X1 u0_u0_u1_U27 (.A( u0_u0_u1_n38 ) , .ZN( u0_u0_u1_n6 ) );
  AND2_X1 u0_u0_u1_U28 (.ZN( u0_u0_u1_n40 ) , .A2( u0_u0_u1_n56 ) , .A1( u0_u0_u1_n60 ) );
  INV_X1 u0_u0_u1_U29 (.A( u0_u0_u1_n58 ) , .ZN( u0_u0_u1_n9 ) );
  INV_X1 u0_u0_u1_U3 (.A( u0_u0_u1_n30 ) , .ZN( u0_u0_u1_n7 ) );
  AOI221_X1 u0_u0_u1_U30 (.A( u0_u0_u1_n1 ) , .C1( u0_u0_u1_n11 ) , .C2( u0_u0_u1_n14 ) , .B2( u0_u0_u1_n17 ) , .ZN( u0_u0_u1_n22 ) , .B1( u0_u0_u1_n49 ) );
  INV_X1 u0_u0_u1_U31 (.ZN( u0_u0_u1_n1 ) , .A( u0_u0_u1_n92 ) );
  AOI211_X1 u0_u0_u1_U32 (.C2( u0_u0_u1_n50 ) , .C1( u0_u0_u1_n57 ) , .A( u0_u0_u1_n71 ) , .ZN( u0_u0_u1_n92 ) , .B( u0_u0_u1_n93 ) );
  AOI21_X1 u0_u0_u1_U33 (.A( u0_u0_u1_n37 ) , .B1( u0_u0_u1_n54 ) , .B2( u0_u0_u1_n68 ) , .ZN( u0_u0_u1_n93 ) );
  OAI221_X1 u0_u0_u1_U34 (.C1( u0_u0_u1_n15 ) , .B1( u0_u0_u1_n2 ) , .B2( u0_u0_u1_n37 ) , .ZN( u0_u0_u1_n51 ) , .C2( u0_u0_u1_n60 ) , .A( u0_u0_u1_n70 ) );
  INV_X1 u0_u0_u1_U35 (.ZN( u0_u0_u1_n2 ) , .A( u0_u0_u1_n41 ) );
  AOI211_X1 u0_u0_u1_U36 (.C1( u0_u0_u1_n30 ) , .C2( u0_u0_u1_n43 ) , .ZN( u0_u0_u1_n70 ) , .A( u0_u0_u1_n71 ) , .B( u0_u0_u1_n72 ) );
  NOR2_X1 u0_u0_u1_U37 (.A2( u0_u0_u1_n13 ) , .A1( u0_u0_u1_n21 ) , .ZN( u0_u0_u1_n91 ) );
  AOI211_X1 u0_u0_u1_U38 (.C1( u0_u0_u1_n18 ) , .ZN( u0_u0_u1_n24 ) , .C2( u0_u0_u1_n25 ) , .A( u0_u0_u1_n26 ) , .B( u0_u0_u1_n27 ) );
  AOI21_X1 u0_u0_u1_U39 (.ZN( u0_u0_u1_n27 ) , .B2( u0_u0_u1_n28 ) , .A( u0_u0_u1_n29 ) , .B1( u0_u0_u1_n7 ) );
  AOI221_X1 u0_u0_u1_U4 (.B1( u0_u0_u1_n14 ) , .ZN( u0_u0_u1_n47 ) , .B2( u0_u0_u1_n48 ) , .C1( u0_u0_u1_n49 ) , .C2( u0_u0_u1_n50 ) , .A( u0_u0_u1_n51 ) );
  OR2_X1 u0_u0_u1_U40 (.ZN( u0_u0_u1_n26 ) , .A1( u0_u0_u1_n31 ) , .A2( u0_u0_u1_n32 ) );
  NAND2_X1 u0_u0_u1_U41 (.A2( u0_u0_u1_n29 ) , .ZN( u0_u0_u1_n43 ) , .A1( u0_u0_u1_n61 ) );
  NAND2_X1 u0_u0_u1_U42 (.A1( u0_u0_u1_n37 ) , .ZN( u0_u0_u1_n50 ) , .A2( u0_u0_u1_n77 ) );
  NAND2_X1 u0_u0_u1_U43 (.ZN( u0_u0_u1_n33 ) , .A1( u0_u0_u1_n84 ) , .A2( u0_u0_u1_n90 ) );
  NOR2_X1 u0_u0_u1_U44 (.A2( u0_u0_u1_n29 ) , .A1( u0_u0_u1_n68 ) , .ZN( u0_u0_u1_n72 ) );
  AOI21_X1 u0_u0_u1_U45 (.B1( u0_u0_u1_n39 ) , .ZN( u0_u0_u1_n59 ) , .B2( u0_u0_u1_n60 ) , .A( u0_u0_u1_n61 ) );
  NAND2_X1 u0_u0_u1_U46 (.A2( u0_u0_u1_n19 ) , .A1( u0_u0_u1_n20 ) , .ZN( u0_u0_u1_n77 ) );
  NAND2_X1 u0_u0_u1_U47 (.ZN( u0_u0_u1_n60 ) , .A1( u0_u0_u1_n91 ) , .A2( u0_u0_u1_n94 ) );
  NAND2_X1 u0_u0_u1_U48 (.ZN( u0_u0_u1_n35 ) , .A1( u0_u0_u1_n87 ) , .A2( u0_u0_u1_n90 ) );
  NAND2_X1 u0_u0_u1_U49 (.ZN( u0_u0_u1_n54 ) , .A2( u0_u0_u1_n89 ) , .A1( u0_u0_u1_n90 ) );
  AOI211_X1 u0_u0_u1_U5 (.C1( u0_u0_u1_n42 ) , .B( u0_u0_u1_n44 ) , .C2( u0_u0_u1_n50 ) , .A( u0_u0_u1_n51 ) , .ZN( u0_u0_u1_n65 ) );
  AOI21_X1 u0_u0_u1_U50 (.ZN( u0_u0_u1_n31 ) , .B1( u0_u0_u1_n35 ) , .B2( u0_u0_u1_n36 ) , .A( u0_u0_u1_n37 ) );
  INV_X1 u0_u0_u1_U51 (.ZN( u0_u0_u1_n14 ) , .A( u0_u0_u1_n29 ) );
  NAND2_X1 u0_u0_u1_U52 (.ZN( u0_u0_u1_n73 ) , .A1( u0_u0_u1_n89 ) , .A2( u0_u0_u1_n94 ) );
  NAND2_X1 u0_u0_u1_U53 (.ZN( u0_u0_u1_n58 ) , .A1( u0_u0_u1_n87 ) , .A2( u0_u0_u1_n94 ) );
  NAND2_X1 u0_u0_u1_U54 (.ZN( u0_u0_u1_n68 ) , .A2( u0_u0_u1_n85 ) , .A1( u0_u0_u1_n91 ) );
  NAND2_X1 u0_u0_u1_U55 (.ZN( u0_u0_u1_n36 ) , .A1( u0_u0_u1_n86 ) , .A2( u0_u0_u1_n91 ) );
  NAND2_X1 u0_u0_u1_U56 (.ZN( u0_u0_u1_n56 ) , .A1( u0_u0_u1_n84 ) , .A2( u0_u0_u1_n85 ) );
  NAND2_X1 u0_u0_u1_U57 (.ZN( u0_u0_u1_n39 ) , .A1( u0_u0_u1_n90 ) , .A2( u0_u0_u1_n91 ) );
  NAND2_X1 u0_u0_u1_U58 (.ZN( u0_u0_u1_n34 ) , .A1( u0_u0_u1_n84 ) , .A2( u0_u0_u1_n94 ) );
  OAI21_X1 u0_u0_u1_U59 (.A( u0_u0_u1_n22 ) , .B2( u0_u0_u1_n29 ) , .B1( u0_u0_u1_n60 ) , .ZN( u0_u0_u1_n80 ) );
  AOI22_X1 u0_u0_u1_U6 (.B1( u0_u0_u1_n16 ) , .A1( u0_u0_u1_n18 ) , .ZN( u0_u0_u1_n64 ) , .A2( u0_u0_u1_n75 ) , .B2( u0_u0_u1_n76 ) );
  NAND2_X1 u0_u0_u1_U60 (.ZN( u0_u0_u1_n69 ) , .A1( u0_u0_u1_n86 ) , .A2( u0_u0_u1_n89 ) );
  NAND2_X1 u0_u0_u1_U61 (.ZN( u0_u0_u1_n74 ) , .A2( u0_u0_u1_n85 ) , .A1( u0_u0_u1_n87 ) );
  NAND2_X1 u0_u0_u1_U62 (.ZN( u0_u0_u1_n38 ) , .A1( u0_u0_u1_n85 ) , .A2( u0_u0_u1_n89 ) );
  NAND2_X1 u0_u0_u1_U63 (.ZN( u0_u0_u1_n28 ) , .A1( u0_u0_u1_n84 ) , .A2( u0_u0_u1_n86 ) );
  INV_X1 u0_u0_u1_U64 (.ZN( u0_u0_u1_n16 ) , .A( u0_u0_u1_n37 ) );
  INV_X1 u0_u0_u1_U65 (.ZN( u0_u0_u1_n17 ) , .A( u0_u0_u1_n61 ) );
  NAND2_X1 u0_u0_u1_U66 (.ZN( u0_u0_u1_n66 ) , .A1( u0_u0_u1_n86 ) , .A2( u0_u0_u1_n87 ) );
  OAI21_X1 u0_u0_u1_U67 (.B1( u0_u0_u1_n29 ) , .A( u0_u0_u1_n4 ) , .ZN( u0_u0_u1_n44 ) , .B2( u0_u0_u1_n66 ) );
  INV_X1 u0_u0_u1_U68 (.ZN( u0_u0_u1_n4 ) , .A( u0_u0_u1_n67 ) );
  AOI21_X1 u0_u0_u1_U69 (.A( u0_u0_u1_n61 ) , .ZN( u0_u0_u1_n67 ) , .B1( u0_u0_u1_n68 ) , .B2( u0_u0_u1_n69 ) );
  NAND2_X1 u0_u0_u1_U7 (.A2( u0_u0_u1_n33 ) , .A1( u0_u0_u1_n55 ) , .ZN( u0_u0_u1_n75 ) );
  NOR2_X1 u0_u0_u1_U70 (.A2( u0_u0_X_7 ) , .A1( u0_u0_X_8 ) , .ZN( u0_u0_u1_n94 ) );
  NOR2_X1 u0_u0_u1_U71 (.A1( u0_u0_X_12 ) , .A2( u0_u0_X_9 ) , .ZN( u0_u0_u1_n89 ) );
  NOR2_X1 u0_u0_u1_U72 (.A2( u0_u0_X_8 ) , .A1( u0_u0_u1_n12 ) , .ZN( u0_u0_u1_n90 ) );
  NOR2_X1 u0_u0_u1_U73 (.A2( u0_u0_X_12 ) , .A1( u0_u0_u1_n13 ) , .ZN( u0_u0_u1_n87 ) );
  NOR2_X1 u0_u0_u1_U74 (.A2( u0_u0_X_9 ) , .A1( u0_u0_u1_n21 ) , .ZN( u0_u0_u1_n84 ) );
  NAND2_X1 u0_u0_u1_U75 (.A1( u0_u0_X_10 ) , .A2( u0_u0_u1_n20 ) , .ZN( u0_u0_u1_n29 ) );
  NAND2_X1 u0_u0_u1_U76 (.A2( u0_u0_X_10 ) , .A1( u0_u0_X_11 ) , .ZN( u0_u0_u1_n37 ) );
  NAND2_X1 u0_u0_u1_U77 (.A1( u0_u0_X_11 ) , .A2( u0_u0_u1_n19 ) , .ZN( u0_u0_u1_n61 ) );
  AND2_X1 u0_u0_u1_U78 (.A2( u0_u0_X_7 ) , .A1( u0_u0_X_8 ) , .ZN( u0_u0_u1_n85 ) );
  AND2_X1 u0_u0_u1_U79 (.A1( u0_u0_X_8 ) , .A2( u0_u0_u1_n12 ) , .ZN( u0_u0_u1_n86 ) );
  NOR2_X1 u0_u0_u1_U8 (.ZN( u0_u0_u1_n71 ) , .A2( u0_u0_u1_n73 ) , .A1( u0_u0_u1_n77 ) );
  INV_X1 u0_u0_u1_U80 (.A( u0_u0_X_10 ) , .ZN( u0_u0_u1_n19 ) );
  INV_X1 u0_u0_u1_U81 (.A( u0_u0_X_9 ) , .ZN( u0_u0_u1_n13 ) );
  INV_X1 u0_u0_u1_U82 (.A( u0_u0_X_11 ) , .ZN( u0_u0_u1_n20 ) );
  INV_X1 u0_u0_u1_U83 (.A( u0_u0_X_12 ) , .ZN( u0_u0_u1_n21 ) );
  INV_X1 u0_u0_u1_U84 (.A( u0_u0_X_7 ) , .ZN( u0_u0_u1_n12 ) );
  NAND4_X1 u0_u0_u1_U85 (.ZN( u0_out0_18 ) , .A1( u0_u0_u1_n22 ) , .A3( u0_u0_u1_n23 ) , .A4( u0_u0_u1_n24 ) , .A2( u0_u0_u1_n3 ) );
  AOI22_X1 u0_u0_u1_U86 (.A1( u0_u0_u1_n17 ) , .ZN( u0_u0_u1_n23 ) , .A2( u0_u0_u1_n41 ) , .B1( u0_u0_u1_n42 ) , .B2( u0_u0_u1_n43 ) );
  INV_X1 u0_u0_u1_U87 (.ZN( u0_u0_u1_n3 ) , .A( u0_u0_u1_n44 ) );
  NAND4_X1 u0_u0_u1_U88 (.ZN( u0_out0_2 ) , .A1( u0_u0_u1_n10 ) , .A2( u0_u0_u1_n45 ) , .A3( u0_u0_u1_n46 ) , .A4( u0_u0_u1_n47 ) );
  OAI21_X1 u0_u0_u1_U89 (.A( u0_u0_u1_n43 ) , .ZN( u0_u0_u1_n45 ) , .B2( u0_u0_u1_n57 ) , .B1( u0_u0_u1_n9 ) );
  OAI21_X1 u0_u0_u1_U9 (.A( u0_u0_u1_n43 ) , .B1( u0_u0_u1_n48 ) , .B2( u0_u0_u1_n6 ) , .ZN( u0_u0_u1_n88 ) );
  INV_X1 u0_u0_u1_U90 (.ZN( u0_u0_u1_n10 ) , .A( u0_u0_u1_n59 ) );
  NAND4_X1 u0_u0_u1_U91 (.ZN( u0_out0_28 ) , .A1( u0_u0_u1_n62 ) , .A2( u0_u0_u1_n63 ) , .A3( u0_u0_u1_n64 ) , .A4( u0_u0_u1_n65 ) );
  OAI21_X1 u0_u0_u1_U92 (.B1( u0_u0_u1_n14 ) , .B2( u0_u0_u1_n50 ) , .A( u0_u0_u1_n6 ) , .ZN( u0_u0_u1_n62 ) );
  OAI21_X1 u0_u0_u1_U93 (.B1( u0_u0_u1_n11 ) , .A( u0_u0_u1_n43 ) , .B2( u0_u0_u1_n49 ) , .ZN( u0_u0_u1_n63 ) );
  OR4_X1 u0_u0_u1_U94 (.ZN( u0_out0_13 ) , .A1( u0_u0_u1_n78 ) , .A2( u0_u0_u1_n79 ) , .A3( u0_u0_u1_n80 ) , .A4( u0_u0_u1_n81 ) );
  AOI21_X1 u0_u0_u1_U95 (.B1( u0_u0_u1_n54 ) , .B2( u0_u0_u1_n58 ) , .A( u0_u0_u1_n61 ) , .ZN( u0_u0_u1_n78 ) );
  AOI21_X1 u0_u0_u1_U96 (.B2( u0_u0_u1_n29 ) , .B1( u0_u0_u1_n37 ) , .A( u0_u0_u1_n73 ) , .ZN( u0_u0_u1_n79 ) );
  NAND3_X1 u0_u0_u1_U97 (.ZN( u0_u0_u1_n25 ) , .A1( u0_u0_u1_n38 ) , .A2( u0_u0_u1_n39 ) , .A3( u0_u0_u1_n40 ) );
  NAND3_X1 u0_u0_u1_U98 (.A1( u0_u0_u1_n38 ) , .ZN( u0_u0_u1_n53 ) , .A2( u0_u0_u1_n54 ) , .A3( u0_u0_u1_n55 ) );
  NAND3_X1 u0_u0_u1_U99 (.A2( u0_u0_u1_n35 ) , .ZN( u0_u0_u1_n52 ) , .A1( u0_u0_u1_n56 ) , .A3( u0_u0_u1_n8 ) );
  OAI22_X1 u0_u0_u2_U10 (.B2( u0_u0_u2_n21 ) , .ZN( u0_u0_u2_n29 ) , .A1( u0_u0_u2_n36 ) , .A2( u0_u0_u2_n37 ) , .B1( u0_u0_u2_n38 ) );
  NAND3_X1 u0_u0_u2_U100 (.A3( u0_u0_u2_n51 ) , .A1( u0_u0_u2_n85 ) , .A2( u0_u0_u2_n89 ) , .ZN( u0_u0_u2_n91 ) );
  NOR3_X1 u0_u0_u2_U11 (.A2( u0_u0_u2_n1 ) , .A3( u0_u0_u2_n14 ) , .ZN( u0_u0_u2_n38 ) , .A1( u0_u0_u2_n39 ) );
  AOI21_X1 u0_u0_u2_U12 (.A( u0_u0_u2_n18 ) , .B1( u0_u0_u2_n5 ) , .ZN( u0_u0_u2_n64 ) , .B2( u0_u0_u2_n66 ) );
  INV_X1 u0_u0_u2_U13 (.A( u0_u0_u2_n39 ) , .ZN( u0_u0_u2_n5 ) );
  AOI21_X1 u0_u0_u2_U14 (.A( u0_u0_u2_n17 ) , .B2( u0_u0_u2_n34 ) , .B1( u0_u0_u2_n4 ) , .ZN( u0_u0_u2_n45 ) );
  AOI21_X1 u0_u0_u2_U15 (.A( u0_u0_u2_n18 ) , .B1( u0_u0_u2_n37 ) , .ZN( u0_u0_u2_n44 ) , .B2( u0_u0_u2_n46 ) );
  INV_X1 u0_u0_u2_U16 (.ZN( u0_u0_u2_n18 ) , .A( u0_u0_u2_n33 ) );
  INV_X1 u0_u0_u2_U17 (.ZN( u0_u0_u2_n1 ) , .A( u0_u0_u2_n69 ) );
  NAND2_X1 u0_u0_u2_U18 (.A1( u0_u0_u2_n37 ) , .ZN( u0_u0_u2_n39 ) , .A2( u0_u0_u2_n67 ) );
  INV_X1 u0_u0_u2_U19 (.ZN( u0_u0_u2_n19 ) , .A( u0_u0_u2_n36 ) );
  INV_X1 u0_u0_u2_U20 (.ZN( u0_u0_u2_n16 ) , .A( u0_u0_u2_n52 ) );
  NAND2_X1 u0_u0_u2_U21 (.ZN( u0_u0_u2_n32 ) , .A2( u0_u0_u2_n50 ) , .A1( u0_u0_u2_n57 ) );
  INV_X1 u0_u0_u2_U22 (.ZN( u0_u0_u2_n11 ) , .A( u0_u0_u2_n76 ) );
  INV_X1 u0_u0_u2_U23 (.ZN( u0_u0_u2_n14 ) , .A( u0_u0_u2_n50 ) );
  INV_X1 u0_u0_u2_U24 (.A( u0_u0_u2_n34 ) , .ZN( u0_u0_u2_n8 ) );
  INV_X1 u0_u0_u2_U25 (.ZN( u0_u0_u2_n12 ) , .A( u0_u0_u2_n70 ) );
  INV_X1 u0_u0_u2_U26 (.A( u0_u0_u2_n73 ) , .ZN( u0_u0_u2_n9 ) );
  INV_X1 u0_u0_u2_U27 (.ZN( u0_u0_u2_n10 ) , .A( u0_u0_u2_n58 ) );
  INV_X1 u0_u0_u2_U28 (.ZN( u0_u0_u2_n13 ) , .A( u0_u0_u2_n35 ) );
  NAND2_X1 u0_u0_u2_U29 (.ZN( u0_u0_u2_n71 ) , .A1( u0_u0_u2_n72 ) , .A2( u0_u0_u2_n73 ) );
  NOR2_X1 u0_u0_u2_U3 (.A2( u0_u0_u2_n12 ) , .ZN( u0_u0_u2_n68 ) , .A1( u0_u0_u2_n9 ) );
  INV_X1 u0_u0_u2_U30 (.A( u0_u0_u2_n57 ) , .ZN( u0_u0_u2_n7 ) );
  INV_X1 u0_u0_u2_U31 (.A( u0_u0_u2_n31 ) , .ZN( u0_u0_u2_n6 ) );
  OAI21_X1 u0_u0_u2_U32 (.B2( u0_u0_u2_n10 ) , .ZN( u0_u0_u2_n31 ) , .B1( u0_u0_u2_n32 ) , .A( u0_u0_u2_n33 ) );
  NOR2_X1 u0_u0_u2_U33 (.A2( u0_u0_u2_n20 ) , .A1( u0_u0_u2_n23 ) , .ZN( u0_u0_u2_n33 ) );
  NOR2_X1 u0_u0_u2_U34 (.A1( u0_u0_u2_n49 ) , .ZN( u0_u0_u2_n52 ) , .A2( u0_u0_u2_n75 ) );
  NOR2_X1 u0_u0_u2_U35 (.A1( u0_u0_u2_n33 ) , .ZN( u0_u0_u2_n36 ) , .A2( u0_u0_u2_n51 ) );
  AOI211_X1 u0_u0_u2_U36 (.C2( u0_u0_u2_n10 ) , .C1( u0_u0_u2_n51 ) , .ZN( u0_u0_u2_n59 ) , .A( u0_u0_u2_n92 ) , .B( u0_u0_u2_n93 ) );
  OAI22_X1 u0_u0_u2_U37 (.B2( u0_u0_u2_n21 ) , .A1( u0_u0_u2_n37 ) , .A2( u0_u0_u2_n52 ) , .B1( u0_u0_u2_n56 ) , .ZN( u0_u0_u2_n92 ) );
  OAI221_X1 u0_u0_u2_U38 (.C2( u0_u0_u2_n17 ) , .B2( u0_u0_u2_n18 ) , .A( u0_u0_u2_n40 ) , .C1( u0_u0_u2_n57 ) , .B1( u0_u0_u2_n76 ) , .ZN( u0_u0_u2_n93 ) );
  OAI221_X1 u0_u0_u2_U39 (.C1( u0_u0_u2_n21 ) , .ZN( u0_u0_u2_n26 ) , .B1( u0_u0_u2_n36 ) , .B2( u0_u0_u2_n46 ) , .C2( u0_u0_u2_n66 ) , .A( u0_u0_u2_n74 ) );
  INV_X1 u0_u0_u2_U4 (.ZN( u0_u0_u2_n4 ) , .A( u0_u0_u2_n55 ) );
  OAI21_X1 u0_u0_u2_U40 (.B2( u0_u0_u2_n11 ) , .B1( u0_u0_u2_n13 ) , .ZN( u0_u0_u2_n74 ) , .A( u0_u0_u2_n75 ) );
  OAI221_X1 u0_u0_u2_U41 (.C2( u0_u0_u2_n22 ) , .ZN( u0_u0_u2_n27 ) , .C1( u0_u0_u2_n4 ) , .B1( u0_u0_u2_n52 ) , .B2( u0_u0_u2_n53 ) , .A( u0_u0_u2_n54 ) );
  AND3_X1 u0_u0_u2_U42 (.ZN( u0_u0_u2_n53 ) , .A1( u0_u0_u2_n56 ) , .A2( u0_u0_u2_n57 ) , .A3( u0_u0_u2_n58 ) );
  AOI22_X1 u0_u0_u2_U43 (.A2( u0_u0_u2_n1 ) , .A1( u0_u0_u2_n33 ) , .B1( u0_u0_u2_n49 ) , .ZN( u0_u0_u2_n54 ) , .B2( u0_u0_u2_n9 ) );
  AOI21_X1 u0_u0_u2_U44 (.B2( u0_u0_u2_n1 ) , .B1( u0_u0_u2_n16 ) , .ZN( u0_u0_u2_n40 ) , .A( u0_u0_u2_n94 ) );
  AND3_X1 u0_u0_u2_U45 (.A3( u0_u0_u2_n33 ) , .A1( u0_u0_u2_n85 ) , .A2( u0_u0_u2_n89 ) , .ZN( u0_u0_u2_n94 ) );
  OAI21_X1 u0_u0_u2_U46 (.B1( u0_u0_u2_n36 ) , .ZN( u0_u0_u2_n43 ) , .B2( u0_u0_u2_n47 ) , .A( u0_u0_u2_n48 ) );
  OAI21_X1 u0_u0_u2_U47 (.B2( u0_u0_u2_n12 ) , .B1( u0_u0_u2_n13 ) , .ZN( u0_u0_u2_n48 ) , .A( u0_u0_u2_n49 ) );
  NOR3_X1 u0_u0_u2_U48 (.A2( u0_u0_u2_n11 ) , .A3( u0_u0_u2_n14 ) , .ZN( u0_u0_u2_n47 ) , .A1( u0_u0_u2_n8 ) );
  OAI21_X1 u0_u0_u2_U49 (.ZN( u0_u0_u2_n25 ) , .B1( u0_u0_u2_n36 ) , .B2( u0_u0_u2_n68 ) , .A( u0_u0_u2_n88 ) );
  NOR4_X1 u0_u0_u2_U5 (.ZN( u0_u0_u2_n61 ) , .A1( u0_u0_u2_n62 ) , .A2( u0_u0_u2_n63 ) , .A3( u0_u0_u2_n64 ) , .A4( u0_u0_u2_n65 ) );
  NAND2_X1 u0_u0_u2_U50 (.ZN( u0_u0_u2_n34 ) , .A1( u0_u0_u2_n82 ) , .A2( u0_u0_u2_n89 ) );
  NAND2_X1 u0_u0_u2_U51 (.ZN( u0_u0_u2_n46 ) , .A1( u0_u0_u2_n81 ) , .A2( u0_u0_u2_n84 ) );
  NAND2_X1 u0_u0_u2_U52 (.ZN( u0_u0_u2_n37 ) , .A2( u0_u0_u2_n83 ) , .A1( u0_u0_u2_n85 ) );
  NAND2_X1 u0_u0_u2_U53 (.ZN( u0_u0_u2_n57 ) , .A2( u0_u0_u2_n84 ) , .A1( u0_u0_u2_n89 ) );
  INV_X1 u0_u0_u2_U54 (.ZN( u0_u0_u2_n21 ) , .A( u0_u0_u2_n49 ) );
  INV_X1 u0_u0_u2_U55 (.ZN( u0_u0_u2_n22 ) , .A( u0_u0_u2_n51 ) );
  NAND2_X1 u0_u0_u2_U56 (.ZN( u0_u0_u2_n76 ) , .A2( u0_u0_u2_n83 ) , .A1( u0_u0_u2_n87 ) );
  NAND2_X1 u0_u0_u2_U57 (.ZN( u0_u0_u2_n58 ) , .A2( u0_u0_u2_n82 ) , .A1( u0_u0_u2_n83 ) );
  NAND2_X1 u0_u0_u2_U58 (.ZN( u0_u0_u2_n50 ) , .A2( u0_u0_u2_n82 ) , .A1( u0_u0_u2_n86 ) );
  NAND2_X1 u0_u0_u2_U59 (.ZN( u0_u0_u2_n56 ) , .A2( u0_u0_u2_n84 ) , .A1( u0_u0_u2_n86 ) );
  AOI21_X1 u0_u0_u2_U6 (.B1( u0_u0_u2_n34 ) , .A( u0_u0_u2_n52 ) , .ZN( u0_u0_u2_n62 ) , .B2( u0_u0_u2_n70 ) );
  NAND2_X1 u0_u0_u2_U60 (.ZN( u0_u0_u2_n35 ) , .A2( u0_u0_u2_n86 ) , .A1( u0_u0_u2_n87 ) );
  NAND2_X1 u0_u0_u2_U61 (.ZN( u0_u0_u2_n70 ) , .A1( u0_u0_u2_n85 ) , .A2( u0_u0_u2_n86 ) );
  NAND2_X1 u0_u0_u2_U62 (.ZN( u0_u0_u2_n66 ) , .A1( u0_u0_u2_n81 ) , .A2( u0_u0_u2_n82 ) );
  NAND2_X1 u0_u0_u2_U63 (.ZN( u0_u0_u2_n67 ) , .A2( u0_u0_u2_n81 ) , .A1( u0_u0_u2_n85 ) );
  INV_X1 u0_u0_u2_U64 (.ZN( u0_u0_u2_n17 ) , .A( u0_u0_u2_n75 ) );
  NAND2_X1 u0_u0_u2_U65 (.ZN( u0_u0_u2_n73 ) , .A1( u0_u0_u2_n87 ) , .A2( u0_u0_u2_n89 ) );
  NAND2_X1 u0_u0_u2_U66 (.ZN( u0_u0_u2_n69 ) , .A2( u0_u0_u2_n81 ) , .A1( u0_u0_u2_n87 ) );
  NAND2_X1 u0_u0_u2_U67 (.ZN( u0_u0_u2_n72 ) , .A1( u0_u0_u2_n83 ) , .A2( u0_u0_u2_n84 ) );
  INV_X1 u0_u0_u2_U68 (.ZN( u0_u0_u2_n2 ) , .A( u0_u0_u2_n90 ) );
  OAI21_X1 u0_u0_u2_U69 (.B2( u0_u0_u2_n46 ) , .B1( u0_u0_u2_n52 ) , .ZN( u0_u0_u2_n90 ) , .A( u0_u0_u2_n91 ) );
  AOI21_X1 u0_u0_u2_U7 (.A( u0_u0_u2_n17 ) , .B2( u0_u0_u2_n46 ) , .B1( u0_u0_u2_n58 ) , .ZN( u0_u0_u2_n65 ) );
  NOR2_X1 u0_u0_u2_U70 (.A2( u0_u0_X_16 ) , .A1( u0_u0_u2_n23 ) , .ZN( u0_u0_u2_n49 ) );
  NOR2_X1 u0_u0_u2_U71 (.A2( u0_u0_X_13 ) , .A1( u0_u0_X_14 ) , .ZN( u0_u0_u2_n89 ) );
  NOR2_X1 u0_u0_u2_U72 (.A2( u0_u0_X_16 ) , .A1( u0_u0_X_17 ) , .ZN( u0_u0_u2_n51 ) );
  NOR2_X1 u0_u0_u2_U73 (.A2( u0_u0_X_15 ) , .A1( u0_u0_X_18 ) , .ZN( u0_u0_u2_n85 ) );
  NOR2_X1 u0_u0_u2_U74 (.A2( u0_u0_X_14 ) , .A1( u0_u0_u2_n15 ) , .ZN( u0_u0_u2_n86 ) );
  NOR2_X1 u0_u0_u2_U75 (.A2( u0_u0_X_15 ) , .A1( u0_u0_u2_n24 ) , .ZN( u0_u0_u2_n87 ) );
  NOR2_X1 u0_u0_u2_U76 (.A2( u0_u0_X_17 ) , .A1( u0_u0_u2_n20 ) , .ZN( u0_u0_u2_n75 ) );
  AND2_X1 u0_u0_u2_U77 (.A1( u0_u0_X_15 ) , .A2( u0_u0_u2_n24 ) , .ZN( u0_u0_u2_n84 ) );
  AND2_X1 u0_u0_u2_U78 (.A2( u0_u0_X_15 ) , .A1( u0_u0_X_18 ) , .ZN( u0_u0_u2_n82 ) );
  AND2_X1 u0_u0_u2_U79 (.A1( u0_u0_X_14 ) , .A2( u0_u0_u2_n15 ) , .ZN( u0_u0_u2_n83 ) );
  AOI21_X1 u0_u0_u2_U8 (.A( u0_u0_u2_n22 ) , .ZN( u0_u0_u2_n63 ) , .B1( u0_u0_u2_n68 ) , .B2( u0_u0_u2_n69 ) );
  AND2_X1 u0_u0_u2_U80 (.A1( u0_u0_X_13 ) , .A2( u0_u0_X_14 ) , .ZN( u0_u0_u2_n81 ) );
  INV_X1 u0_u0_u2_U81 (.A( u0_u0_X_16 ) , .ZN( u0_u0_u2_n20 ) );
  INV_X1 u0_u0_u2_U82 (.A( u0_u0_X_17 ) , .ZN( u0_u0_u2_n23 ) );
  INV_X1 u0_u0_u2_U83 (.A( u0_u0_X_13 ) , .ZN( u0_u0_u2_n15 ) );
  INV_X1 u0_u0_u2_U84 (.A( u0_u0_X_18 ) , .ZN( u0_u0_u2_n24 ) );
  NAND4_X1 u0_u0_u2_U85 (.ZN( u0_out0_30 ) , .A1( u0_u0_u2_n2 ) , .A2( u0_u0_u2_n40 ) , .A3( u0_u0_u2_n41 ) , .A4( u0_u0_u2_n42 ) );
  NOR3_X1 u0_u0_u2_U86 (.ZN( u0_u0_u2_n42 ) , .A1( u0_u0_u2_n43 ) , .A2( u0_u0_u2_n44 ) , .A3( u0_u0_u2_n45 ) );
  AOI21_X1 u0_u0_u2_U87 (.A( u0_u0_u2_n27 ) , .ZN( u0_u0_u2_n41 ) , .B2( u0_u0_u2_n51 ) , .B1( u0_u0_u2_n7 ) );
  NAND4_X1 u0_u0_u2_U88 (.ZN( u0_out0_24 ) , .A2( u0_u0_u2_n2 ) , .A1( u0_u0_u2_n59 ) , .A3( u0_u0_u2_n77 ) , .A4( u0_u0_u2_n78 ) );
  AOI221_X1 u0_u0_u2_U89 (.B2( u0_u0_u2_n16 ) , .C2( u0_u0_u2_n19 ) , .C1( u0_u0_u2_n55 ) , .ZN( u0_u0_u2_n78 ) , .B1( u0_u0_u2_n79 ) , .A( u0_u0_u2_n80 ) );
  OAI22_X1 u0_u0_u2_U9 (.A1( u0_u0_u2_n21 ) , .B1( u0_u0_u2_n22 ) , .B2( u0_u0_u2_n56 ) , .A2( u0_u0_u2_n76 ) , .ZN( u0_u0_u2_n80 ) );
  AOI21_X1 u0_u0_u2_U90 (.A( u0_u0_u2_n25 ) , .B2( u0_u0_u2_n33 ) , .ZN( u0_u0_u2_n77 ) , .B1( u0_u0_u2_n8 ) );
  NAND4_X1 u0_u0_u2_U91 (.ZN( u0_out0_16 ) , .A2( u0_u0_u2_n3 ) , .A1( u0_u0_u2_n59 ) , .A3( u0_u0_u2_n60 ) , .A4( u0_u0_u2_n61 ) );
  AOI22_X1 u0_u0_u2_U92 (.B2( u0_u0_u2_n19 ) , .B1( u0_u0_u2_n32 ) , .A1( u0_u0_u2_n49 ) , .ZN( u0_u0_u2_n60 ) , .A2( u0_u0_u2_n71 ) );
  INV_X1 u0_u0_u2_U93 (.A( u0_u0_u2_n26 ) , .ZN( u0_u0_u2_n3 ) );
  OR4_X1 u0_u0_u2_U94 (.ZN( u0_out0_6 ) , .A1( u0_u0_u2_n25 ) , .A2( u0_u0_u2_n26 ) , .A3( u0_u0_u2_n27 ) , .A4( u0_u0_u2_n28 ) );
  OR3_X1 u0_u0_u2_U95 (.ZN( u0_u0_u2_n28 ) , .A1( u0_u0_u2_n29 ) , .A2( u0_u0_u2_n30 ) , .A3( u0_u0_u2_n6 ) );
  AOI21_X1 u0_u0_u2_U96 (.A( u0_u0_u2_n22 ) , .ZN( u0_u0_u2_n30 ) , .B1( u0_u0_u2_n34 ) , .B2( u0_u0_u2_n35 ) );
  NAND3_X1 u0_u0_u2_U97 (.ZN( u0_u0_u2_n55 ) , .A3( u0_u0_u2_n66 ) , .A1( u0_u0_u2_n67 ) , .A2( u0_u0_u2_n72 ) );
  NAND3_X1 u0_u0_u2_U98 (.A1( u0_u0_u2_n35 ) , .A3( u0_u0_u2_n50 ) , .A2( u0_u0_u2_n58 ) , .ZN( u0_u0_u2_n79 ) );
  NAND3_X1 u0_u0_u2_U99 (.A3( u0_u0_u2_n75 ) , .A1( u0_u0_u2_n85 ) , .ZN( u0_u0_u2_n88 ) , .A2( u0_u0_u2_n89 ) );
  OAI22_X1 u0_u0_u3_U10 (.B2( u0_u0_u3_n23 ) , .A1( u0_u0_u3_n37 ) , .A2( u0_u0_u3_n52 ) , .B1( u0_u0_u3_n74 ) , .ZN( u0_u0_u3_n89 ) );
  OAI211_X1 u0_u0_u3_U11 (.C1( u0_u0_u3_n20 ) , .C2( u0_u0_u3_n59 ) , .A( u0_u0_u3_n6 ) , .ZN( u0_u0_u3_n68 ) , .B( u0_u0_u3_n81 ) );
  AOI221_X1 u0_u0_u3_U12 (.B1( u0_u0_u3_n18 ) , .C2( u0_u0_u3_n54 ) , .B2( u0_u0_u3_n55 ) , .A( u0_u0_u3_n56 ) , .ZN( u0_u0_u3_n81 ) , .C1( u0_u0_u3_n82 ) );
  INV_X1 u0_u0_u3_U13 (.ZN( u0_u0_u3_n6 ) , .A( u0_u0_u3_n89 ) );
  NAND2_X1 u0_u0_u3_U14 (.A1( u0_u0_u3_n32 ) , .A2( u0_u0_u3_n57 ) , .ZN( u0_u0_u3_n82 ) );
  AOI22_X1 u0_u0_u3_U15 (.A1( u0_u0_u3_n18 ) , .B2( u0_u0_u3_n54 ) , .ZN( u0_u0_u3_n64 ) , .A2( u0_u0_u3_n71 ) , .B1( u0_u0_u3_n72 ) );
  NAND2_X1 u0_u0_u3_U16 (.A2( u0_u0_u3_n36 ) , .A1( u0_u0_u3_n5 ) , .ZN( u0_u0_u3_n71 ) );
  NOR2_X1 u0_u0_u3_U17 (.A1( u0_u0_u3_n23 ) , .A2( u0_u0_u3_n37 ) , .ZN( u0_u0_u3_n61 ) );
  AOI21_X1 u0_u0_u3_U18 (.A( u0_u0_u3_n20 ) , .B1( u0_u0_u3_n32 ) , .B2( u0_u0_u3_n41 ) , .ZN( u0_u0_u3_n75 ) );
  NAND2_X1 u0_u0_u3_U19 (.A2( u0_u0_u3_n23 ) , .ZN( u0_u0_u3_n45 ) , .A1( u0_u0_u3_n52 ) );
  NAND2_X1 u0_u0_u3_U20 (.A1( u0_u0_u3_n31 ) , .A2( u0_u0_u3_n35 ) , .ZN( u0_u0_u3_n55 ) );
  INV_X1 u0_u0_u3_U21 (.ZN( u0_u0_u3_n22 ) , .A( u0_u0_u3_n54 ) );
  AND2_X1 u0_u0_u3_U22 (.ZN( u0_u0_u3_n36 ) , .A1( u0_u0_u3_n73 ) , .A2( u0_u0_u3_n74 ) );
  INV_X1 u0_u0_u3_U23 (.ZN( u0_u0_u3_n17 ) , .A( u0_u0_u3_n52 ) );
  NAND2_X1 u0_u0_u3_U24 (.ZN( u0_u0_u3_n47 ) , .A2( u0_u0_u3_n79 ) , .A1( u0_u0_u3_n80 ) );
  NAND2_X1 u0_u0_u3_U25 (.A2( u0_u0_u3_n39 ) , .A1( u0_u0_u3_n63 ) , .ZN( u0_u0_u3_n70 ) );
  NAND2_X1 u0_u0_u3_U26 (.A2( u0_u0_u3_n20 ) , .A1( u0_u0_u3_n22 ) , .ZN( u0_u0_u3_n44 ) );
  INV_X1 u0_u0_u3_U27 (.ZN( u0_u0_u3_n10 ) , .A( u0_u0_u3_n57 ) );
  INV_X1 u0_u0_u3_U28 (.ZN( u0_u0_u3_n11 ) , .A( u0_u0_u3_n59 ) );
  INV_X1 u0_u0_u3_U29 (.ZN( u0_u0_u3_n13 ) , .A( u0_u0_u3_n32 ) );
  INV_X1 u0_u0_u3_U3 (.A( u0_u0_u3_n47 ) , .ZN( u0_u0_u3_n5 ) );
  INV_X1 u0_u0_u3_U30 (.ZN( u0_u0_u3_n2 ) , .A( u0_u0_u3_n48 ) );
  NOR2_X1 u0_u0_u3_U31 (.A1( u0_u0_u3_n18 ) , .A2( u0_u0_u3_n46 ) , .ZN( u0_u0_u3_n52 ) );
  OAI222_X1 u0_u0_u3_U32 (.A1( u0_u0_u3_n23 ) , .C1( u0_u0_u3_n33 ) , .B2( u0_u0_u3_n41 ) , .ZN( u0_u0_u3_n49 ) , .B1( u0_u0_u3_n52 ) , .A2( u0_u0_u3_n79 ) , .C2( u0_u0_u3_n80 ) );
  NOR4_X1 u0_u0_u3_U33 (.ZN( u0_u0_u3_n26 ) , .A1( u0_u0_u3_n27 ) , .A2( u0_u0_u3_n28 ) , .A3( u0_u0_u3_n29 ) , .A4( u0_u0_u3_n30 ) );
  AOI21_X1 u0_u0_u3_U34 (.A( u0_u0_u3_n23 ) , .ZN( u0_u0_u3_n29 ) , .B1( u0_u0_u3_n34 ) , .B2( u0_u0_u3_n35 ) );
  AOI21_X1 u0_u0_u3_U35 (.ZN( u0_u0_u3_n30 ) , .B1( u0_u0_u3_n31 ) , .B2( u0_u0_u3_n32 ) , .A( u0_u0_u3_n33 ) );
  AOI21_X1 u0_u0_u3_U36 (.ZN( u0_u0_u3_n28 ) , .B1( u0_u0_u3_n36 ) , .B2( u0_u0_u3_n37 ) , .A( u0_u0_u3_n38 ) );
  OAI211_X1 u0_u0_u3_U37 (.A( u0_u0_u3_n3 ) , .C2( u0_u0_u3_n33 ) , .C1( u0_u0_u3_n37 ) , .ZN( u0_u0_u3_n48 ) , .B( u0_u0_u3_n60 ) );
  INV_X1 u0_u0_u3_U38 (.ZN( u0_u0_u3_n3 ) , .A( u0_u0_u3_n62 ) );
  AOI221_X1 u0_u0_u3_U39 (.B1( u0_u0_u3_n13 ) , .B2( u0_u0_u3_n17 ) , .C1( u0_u0_u3_n18 ) , .C2( u0_u0_u3_n55 ) , .ZN( u0_u0_u3_n60 ) , .A( u0_u0_u3_n61 ) );
  INV_X1 u0_u0_u3_U4 (.ZN( u0_u0_u3_n4 ) , .A( u0_u0_u3_n58 ) );
  OAI22_X1 u0_u0_u3_U40 (.B1( u0_u0_u3_n20 ) , .A2( u0_u0_u3_n22 ) , .B2( u0_u0_u3_n42 ) , .ZN( u0_u0_u3_n62 ) , .A1( u0_u0_u3_n63 ) );
  AOI211_X1 u0_u0_u3_U41 (.C1( u0_u0_u3_n46 ) , .B( u0_u0_u3_n49 ) , .C2( u0_u0_u3_n58 ) , .A( u0_u0_u3_n68 ) , .ZN( u0_u0_u3_n78 ) );
  AOI211_X1 u0_u0_u3_U42 (.ZN( u0_u0_u3_n65 ) , .C2( u0_u0_u3_n66 ) , .A( u0_u0_u3_n67 ) , .B( u0_u0_u3_n68 ) , .C1( u0_u0_u3_n8 ) );
  INV_X1 u0_u0_u3_U43 (.A( u0_u0_u3_n31 ) , .ZN( u0_u0_u3_n8 ) );
  OAI22_X1 u0_u0_u3_U44 (.B2( u0_u0_u3_n33 ) , .A1( u0_u0_u3_n52 ) , .ZN( u0_u0_u3_n67 ) , .B1( u0_u0_u3_n69 ) , .A2( u0_u0_u3_n9 ) );
  AND3_X1 u0_u0_u3_U45 (.A3( u0_u0_u3_n35 ) , .A1( u0_u0_u3_n43 ) , .A2( u0_u0_u3_n63 ) , .ZN( u0_u0_u3_n69 ) );
  INV_X1 u0_u0_u3_U46 (.ZN( u0_u0_u3_n23 ) , .A( u0_u0_u3_n66 ) );
  NAND2_X1 u0_u0_u3_U47 (.A2( u0_u0_u3_n23 ) , .A1( u0_u0_u3_n33 ) , .ZN( u0_u0_u3_n54 ) );
  NOR2_X1 u0_u0_u3_U48 (.A2( u0_u0_u3_n33 ) , .ZN( u0_u0_u3_n56 ) , .A1( u0_u0_u3_n74 ) );
  NAND2_X1 u0_u0_u3_U49 (.ZN( u0_u0_u3_n37 ) , .A1( u0_u0_u3_n84 ) , .A2( u0_u0_u3_n88 ) );
  INV_X1 u0_u0_u3_U5 (.A( u0_u0_u3_n70 ) , .ZN( u0_u0_u3_n9 ) );
  NAND2_X1 u0_u0_u3_U50 (.ZN( u0_u0_u3_n32 ) , .A2( u0_u0_u3_n85 ) , .A1( u0_u0_u3_n90 ) );
  INV_X1 u0_u0_u3_U51 (.ZN( u0_u0_u3_n20 ) , .A( u0_u0_u3_n46 ) );
  AOI21_X1 u0_u0_u3_U52 (.A( u0_u0_u3_n33 ) , .B1( u0_u0_u3_n41 ) , .B2( u0_u0_u3_n73 ) , .ZN( u0_u0_u3_n93 ) );
  AOI21_X1 u0_u0_u3_U53 (.B1( u0_u0_u3_n1 ) , .B2( u0_u0_u3_n45 ) , .ZN( u0_u0_u3_n77 ) , .A( u0_u0_u3_n92 ) );
  INV_X1 u0_u0_u3_U54 (.ZN( u0_u0_u3_n1 ) , .A( u0_u0_u3_n42 ) );
  AOI21_X1 u0_u0_u3_U55 (.B2( u0_u0_u3_n32 ) , .A( u0_u0_u3_n38 ) , .B1( u0_u0_u3_n63 ) , .ZN( u0_u0_u3_n92 ) );
  INV_X1 u0_u0_u3_U56 (.ZN( u0_u0_u3_n18 ) , .A( u0_u0_u3_n38 ) );
  NAND2_X1 u0_u0_u3_U57 (.ZN( u0_u0_u3_n63 ) , .A2( u0_u0_u3_n90 ) , .A1( u0_u0_u3_n91 ) );
  NAND2_X1 u0_u0_u3_U58 (.ZN( u0_u0_u3_n41 ) , .A2( u0_u0_u3_n87 ) , .A1( u0_u0_u3_n91 ) );
  NAND2_X1 u0_u0_u3_U59 (.ZN( u0_u0_u3_n42 ) , .A1( u0_u0_u3_n86 ) , .A2( u0_u0_u3_n88 ) );
  AOI221_X1 u0_u0_u3_U6 (.B2( u0_u0_u3_n10 ) , .B1( u0_u0_u3_n44 ) , .ZN( u0_u0_u3_n53 ) , .C1( u0_u0_u3_n54 ) , .C2( u0_u0_u3_n55 ) , .A( u0_u0_u3_n56 ) );
  NAND2_X1 u0_u0_u3_U60 (.ZN( u0_u0_u3_n31 ) , .A1( u0_u0_u3_n87 ) , .A2( u0_u0_u3_n88 ) );
  NAND2_X1 u0_u0_u3_U61 (.ZN( u0_u0_u3_n39 ) , .A1( u0_u0_u3_n83 ) , .A2( u0_u0_u3_n86 ) );
  NAND2_X1 u0_u0_u3_U62 (.ZN( u0_u0_u3_n59 ) , .A2( u0_u0_u3_n85 ) , .A1( u0_u0_u3_n87 ) );
  NAND2_X1 u0_u0_u3_U63 (.ZN( u0_u0_u3_n35 ) , .A1( u0_u0_u3_n85 ) , .A2( u0_u0_u3_n86 ) );
  NAND2_X1 u0_u0_u3_U64 (.ZN( u0_u0_u3_n73 ) , .A2( u0_u0_u3_n86 ) , .A1( u0_u0_u3_n91 ) );
  NAND2_X1 u0_u0_u3_U65 (.ZN( u0_u0_u3_n80 ) , .A2( u0_u0_u3_n88 ) , .A1( u0_u0_u3_n90 ) );
  NAND2_X1 u0_u0_u3_U66 (.ZN( u0_u0_u3_n74 ) , .A1( u0_u0_u3_n83 ) , .A2( u0_u0_u3_n87 ) );
  NAND2_X1 u0_u0_u3_U67 (.ZN( u0_u0_u3_n34 ) , .A1( u0_u0_u3_n83 ) , .A2( u0_u0_u3_n90 ) );
  NAND2_X1 u0_u0_u3_U68 (.ZN( u0_u0_u3_n57 ) , .A1( u0_u0_u3_n83 ) , .A2( u0_u0_u3_n84 ) );
  NAND2_X1 u0_u0_u3_U69 (.ZN( u0_u0_u3_n43 ) , .A2( u0_u0_u3_n84 ) , .A1( u0_u0_u3_n91 ) );
  OAI22_X1 u0_u0_u3_U7 (.A1( u0_u0_u3_n19 ) , .B1( u0_u0_u3_n22 ) , .ZN( u0_u0_u3_n27 ) , .A2( u0_u0_u3_n39 ) , .B2( u0_u0_u3_n40 ) );
  NAND2_X1 u0_u0_u3_U70 (.ZN( u0_u0_u3_n79 ) , .A2( u0_u0_u3_n84 ) , .A1( u0_u0_u3_n85 ) );
  NOR2_X1 u0_u0_u3_U71 (.A2( u0_u0_X_19 ) , .A1( u0_u0_X_20 ) , .ZN( u0_u0_u3_n88 ) );
  NOR2_X1 u0_u0_u3_U72 (.A2( u0_u0_X_21 ) , .A1( u0_u0_X_24 ) , .ZN( u0_u0_u3_n84 ) );
  NOR2_X1 u0_u0_u3_U73 (.A2( u0_u0_X_24 ) , .A1( u0_u0_u3_n16 ) , .ZN( u0_u0_u3_n90 ) );
  NOR2_X1 u0_u0_u3_U74 (.A2( u0_u0_X_23 ) , .A1( u0_u0_u3_n21 ) , .ZN( u0_u0_u3_n46 ) );
  NOR2_X1 u0_u0_u3_U75 (.A2( u0_u0_X_19 ) , .A1( u0_u0_u3_n15 ) , .ZN( u0_u0_u3_n91 ) );
  NAND2_X1 u0_u0_u3_U76 (.A1( u0_u0_X_22 ) , .A2( u0_u0_X_23 ) , .ZN( u0_u0_u3_n33 ) );
  NAND2_X1 u0_u0_u3_U77 (.A1( u0_u0_X_23 ) , .A2( u0_u0_u3_n21 ) , .ZN( u0_u0_u3_n38 ) );
  NOR2_X1 u0_u0_u3_U78 (.A2( u0_u0_X_22 ) , .A1( u0_u0_X_23 ) , .ZN( u0_u0_u3_n66 ) );
  AND2_X1 u0_u0_u3_U79 (.A1( u0_u0_X_24 ) , .A2( u0_u0_u3_n16 ) , .ZN( u0_u0_u3_n86 ) );
  AND3_X1 u0_u0_u3_U8 (.ZN( u0_u0_u3_n40 ) , .A1( u0_u0_u3_n41 ) , .A2( u0_u0_u3_n42 ) , .A3( u0_u0_u3_n43 ) );
  AND2_X1 u0_u0_u3_U80 (.A1( u0_u0_X_19 ) , .A2( u0_u0_u3_n15 ) , .ZN( u0_u0_u3_n85 ) );
  AND2_X1 u0_u0_u3_U81 (.A1( u0_u0_X_21 ) , .A2( u0_u0_X_24 ) , .ZN( u0_u0_u3_n87 ) );
  AND2_X1 u0_u0_u3_U82 (.A2( u0_u0_X_19 ) , .A1( u0_u0_X_20 ) , .ZN( u0_u0_u3_n83 ) );
  INV_X1 u0_u0_u3_U83 (.A( u0_u0_X_22 ) , .ZN( u0_u0_u3_n21 ) );
  INV_X1 u0_u0_u3_U84 (.A( u0_u0_X_21 ) , .ZN( u0_u0_u3_n16 ) );
  INV_X1 u0_u0_u3_U85 (.A( u0_u0_X_20 ) , .ZN( u0_u0_u3_n15 ) );
  NAND4_X1 u0_u0_u3_U86 (.ZN( u0_out0_26 ) , .A1( u0_u0_u3_n14 ) , .A2( u0_u0_u3_n76 ) , .A3( u0_u0_u3_n77 ) , .A4( u0_u0_u3_n78 ) );
  INV_X1 u0_u0_u3_U87 (.ZN( u0_u0_u3_n14 ) , .A( u0_u0_u3_n93 ) );
  OAI21_X1 u0_u0_u3_U88 (.B1( u0_u0_u3_n11 ) , .A( u0_u0_u3_n54 ) , .B2( u0_u0_u3_n70 ) , .ZN( u0_u0_u3_n76 ) );
  NAND4_X1 u0_u0_u3_U89 (.ZN( u0_out0_1 ) , .A1( u0_u0_u3_n2 ) , .A2( u0_u0_u3_n24 ) , .A3( u0_u0_u3_n25 ) , .A4( u0_u0_u3_n26 ) );
  INV_X1 u0_u0_u3_U9 (.ZN( u0_u0_u3_n19 ) , .A( u0_u0_u3_n44 ) );
  NAND2_X1 u0_u0_u3_U90 (.A1( u0_u0_u3_n11 ) , .A2( u0_u0_u3_n17 ) , .ZN( u0_u0_u3_n24 ) );
  AOI22_X1 u0_u0_u3_U91 (.A1( u0_u0_u3_n10 ) , .ZN( u0_u0_u3_n25 ) , .A2( u0_u0_u3_n45 ) , .B1( u0_u0_u3_n46 ) , .B2( u0_u0_u3_n47 ) );
  NAND4_X1 u0_u0_u3_U92 (.ZN( u0_out0_20 ) , .A1( u0_u0_u3_n12 ) , .A3( u0_u0_u3_n64 ) , .A4( u0_u0_u3_n65 ) , .A2( u0_u0_u3_n7 ) );
  INV_X1 u0_u0_u3_U93 (.A( u0_u0_u3_n61 ) , .ZN( u0_u0_u3_n7 ) );
  INV_X1 u0_u0_u3_U94 (.ZN( u0_u0_u3_n12 ) , .A( u0_u0_u3_n75 ) );
  OR4_X1 u0_u0_u3_U95 (.ZN( u0_out0_10 ) , .A2( u0_u0_u3_n48 ) , .A1( u0_u0_u3_n49 ) , .A3( u0_u0_u3_n50 ) , .A4( u0_u0_u3_n51 ) );
  OAI222_X1 u0_u0_u3_U96 (.A1( u0_u0_u3_n20 ) , .C2( u0_u0_u3_n23 ) , .B2( u0_u0_u3_n33 ) , .A2( u0_u0_u3_n37 ) , .B1( u0_u0_u3_n39 ) , .ZN( u0_u0_u3_n50 ) , .C1( u0_u0_u3_n59 ) );
  OAI221_X1 u0_u0_u3_U97 (.B1( u0_u0_u3_n36 ) , .C1( u0_u0_u3_n38 ) , .C2( u0_u0_u3_n4 ) , .ZN( u0_u0_u3_n51 ) , .B2( u0_u0_u3_n52 ) , .A( u0_u0_u3_n53 ) );
  NAND3_X1 u0_u0_u3_U98 (.A3( u0_u0_u3_n34 ) , .A2( u0_u0_u3_n42 ) , .ZN( u0_u0_u3_n72 ) , .A1( u0_u0_u3_n73 ) );
  NAND3_X1 u0_u0_u3_U99 (.A1( u0_u0_u3_n34 ) , .A2( u0_u0_u3_n43 ) , .A3( u0_u0_u3_n5 ) , .ZN( u0_u0_u3_n58 ) );
  XOR2_X1 u0_u13_U1 (.B( u0_K14_9 ) , .A( u0_R12_6 ) , .Z( u0_u13_X_9 ) );
  XOR2_X1 u0_u13_U16 (.B( u0_K14_3 ) , .A( u0_R12_2 ) , .Z( u0_u13_X_3 ) );
  XOR2_X1 u0_u13_U2 (.B( u0_K14_8 ) , .A( u0_R12_5 ) , .Z( u0_u13_X_8 ) );
  XOR2_X1 u0_u13_U20 (.B( u0_K14_36 ) , .A( u0_R12_25 ) , .Z( u0_u13_X_36 ) );
  XOR2_X1 u0_u13_U21 (.B( u0_K14_35 ) , .A( u0_R12_24 ) , .Z( u0_u13_X_35 ) );
  XOR2_X1 u0_u13_U22 (.B( u0_K14_34 ) , .A( u0_R12_23 ) , .Z( u0_u13_X_34 ) );
  XOR2_X1 u0_u13_U23 (.B( u0_K14_33 ) , .A( u0_R12_22 ) , .Z( u0_u13_X_33 ) );
  XOR2_X1 u0_u13_U24 (.B( u0_K14_32 ) , .A( u0_R12_21 ) , .Z( u0_u13_X_32 ) );
  XOR2_X1 u0_u13_U25 (.B( u0_K14_31 ) , .A( u0_R12_20 ) , .Z( u0_u13_X_31 ) );
  XOR2_X1 u0_u13_U26 (.B( u0_K14_30 ) , .A( u0_R12_21 ) , .Z( u0_u13_X_30 ) );
  XOR2_X1 u0_u13_U27 (.B( u0_K14_2 ) , .A( u0_R12_1 ) , .Z( u0_u13_X_2 ) );
  XOR2_X1 u0_u13_U28 (.B( u0_K14_29 ) , .A( u0_R12_20 ) , .Z( u0_u13_X_29 ) );
  XOR2_X1 u0_u13_U29 (.B( u0_K14_28 ) , .A( u0_R12_19 ) , .Z( u0_u13_X_28 ) );
  XOR2_X1 u0_u13_U3 (.B( u0_K14_7 ) , .A( u0_R12_4 ) , .Z( u0_u13_X_7 ) );
  XOR2_X1 u0_u13_U30 (.B( u0_K14_27 ) , .A( u0_R12_18 ) , .Z( u0_u13_X_27 ) );
  XOR2_X1 u0_u13_U31 (.B( u0_K14_26 ) , .A( u0_R12_17 ) , .Z( u0_u13_X_26 ) );
  XOR2_X1 u0_u13_U32 (.B( u0_K14_25 ) , .A( u0_R12_16 ) , .Z( u0_u13_X_25 ) );
  XOR2_X1 u0_u13_U33 (.B( u0_K14_24 ) , .A( u0_R12_17 ) , .Z( u0_u13_X_24 ) );
  XOR2_X1 u0_u13_U34 (.B( u0_K14_23 ) , .A( u0_R12_16 ) , .Z( u0_u13_X_23 ) );
  XOR2_X1 u0_u13_U35 (.B( u0_K14_22 ) , .A( u0_R12_15 ) , .Z( u0_u13_X_22 ) );
  XOR2_X1 u0_u13_U36 (.B( u0_K14_21 ) , .A( u0_R12_14 ) , .Z( u0_u13_X_21 ) );
  XOR2_X1 u0_u13_U37 (.B( u0_K14_20 ) , .A( u0_R12_13 ) , .Z( u0_u13_X_20 ) );
  XOR2_X1 u0_u13_U38 (.B( u0_K14_1 ) , .A( u0_R12_32 ) , .Z( u0_u13_X_1 ) );
  XOR2_X1 u0_u13_U39 (.B( u0_K14_19 ) , .A( u0_R12_12 ) , .Z( u0_u13_X_19 ) );
  XOR2_X1 u0_u13_U4 (.B( u0_K14_6 ) , .A( u0_R12_5 ) , .Z( u0_u13_X_6 ) );
  XOR2_X1 u0_u13_U40 (.B( u0_K14_18 ) , .A( u0_R12_13 ) , .Z( u0_u13_X_18 ) );
  XOR2_X1 u0_u13_U41 (.B( u0_K14_17 ) , .A( u0_R12_12 ) , .Z( u0_u13_X_17 ) );
  XOR2_X1 u0_u13_U42 (.B( u0_K14_16 ) , .A( u0_R12_11 ) , .Z( u0_u13_X_16 ) );
  XOR2_X1 u0_u13_U43 (.B( u0_K14_15 ) , .A( u0_R12_10 ) , .Z( u0_u13_X_15 ) );
  XOR2_X1 u0_u13_U44 (.B( u0_K14_14 ) , .A( u0_R12_9 ) , .Z( u0_u13_X_14 ) );
  XOR2_X1 u0_u13_U45 (.B( u0_K14_13 ) , .A( u0_R12_8 ) , .Z( u0_u13_X_13 ) );
  XOR2_X1 u0_u13_U46 (.B( u0_K14_12 ) , .A( u0_R12_9 ) , .Z( u0_u13_X_12 ) );
  XOR2_X1 u0_u13_U47 (.B( u0_K14_11 ) , .A( u0_R12_8 ) , .Z( u0_u13_X_11 ) );
  XOR2_X1 u0_u13_U48 (.B( u0_K14_10 ) , .A( u0_R12_7 ) , .Z( u0_u13_X_10 ) );
  XOR2_X1 u0_u13_U5 (.B( u0_K14_5 ) , .A( u0_R12_4 ) , .Z( u0_u13_X_5 ) );
  XOR2_X1 u0_u13_U6 (.B( u0_K14_4 ) , .A( u0_R12_3 ) , .Z( u0_u13_X_4 ) );
  AND3_X1 u0_u13_u0_U10 (.A2( u0_u13_u0_n112 ) , .ZN( u0_u13_u0_n127 ) , .A3( u0_u13_u0_n130 ) , .A1( u0_u13_u0_n148 ) );
  NAND2_X1 u0_u13_u0_U11 (.ZN( u0_u13_u0_n113 ) , .A1( u0_u13_u0_n139 ) , .A2( u0_u13_u0_n149 ) );
  AND2_X1 u0_u13_u0_U12 (.ZN( u0_u13_u0_n107 ) , .A1( u0_u13_u0_n130 ) , .A2( u0_u13_u0_n140 ) );
  AND2_X1 u0_u13_u0_U13 (.A2( u0_u13_u0_n129 ) , .A1( u0_u13_u0_n130 ) , .ZN( u0_u13_u0_n151 ) );
  AND2_X1 u0_u13_u0_U14 (.A1( u0_u13_u0_n108 ) , .A2( u0_u13_u0_n125 ) , .ZN( u0_u13_u0_n145 ) );
  INV_X1 u0_u13_u0_U15 (.A( u0_u13_u0_n143 ) , .ZN( u0_u13_u0_n173 ) );
  NOR2_X1 u0_u13_u0_U16 (.A2( u0_u13_u0_n136 ) , .ZN( u0_u13_u0_n147 ) , .A1( u0_u13_u0_n160 ) );
  INV_X1 u0_u13_u0_U17 (.ZN( u0_u13_u0_n172 ) , .A( u0_u13_u0_n88 ) );
  OAI222_X1 u0_u13_u0_U18 (.C1( u0_u13_u0_n108 ) , .A1( u0_u13_u0_n125 ) , .B2( u0_u13_u0_n128 ) , .B1( u0_u13_u0_n144 ) , .A2( u0_u13_u0_n158 ) , .C2( u0_u13_u0_n161 ) , .ZN( u0_u13_u0_n88 ) );
  NOR2_X1 u0_u13_u0_U19 (.A1( u0_u13_u0_n163 ) , .A2( u0_u13_u0_n164 ) , .ZN( u0_u13_u0_n95 ) );
  AOI21_X1 u0_u13_u0_U20 (.B1( u0_u13_u0_n103 ) , .ZN( u0_u13_u0_n132 ) , .A( u0_u13_u0_n165 ) , .B2( u0_u13_u0_n93 ) );
  INV_X1 u0_u13_u0_U21 (.A( u0_u13_u0_n142 ) , .ZN( u0_u13_u0_n165 ) );
  OAI221_X1 u0_u13_u0_U22 (.C1( u0_u13_u0_n121 ) , .ZN( u0_u13_u0_n122 ) , .B2( u0_u13_u0_n127 ) , .A( u0_u13_u0_n143 ) , .B1( u0_u13_u0_n144 ) , .C2( u0_u13_u0_n147 ) );
  OAI22_X1 u0_u13_u0_U23 (.B1( u0_u13_u0_n125 ) , .ZN( u0_u13_u0_n126 ) , .A1( u0_u13_u0_n138 ) , .A2( u0_u13_u0_n146 ) , .B2( u0_u13_u0_n147 ) );
  OAI22_X1 u0_u13_u0_U24 (.B1( u0_u13_u0_n131 ) , .A1( u0_u13_u0_n144 ) , .B2( u0_u13_u0_n147 ) , .A2( u0_u13_u0_n90 ) , .ZN( u0_u13_u0_n91 ) );
  AND3_X1 u0_u13_u0_U25 (.A3( u0_u13_u0_n121 ) , .A2( u0_u13_u0_n125 ) , .A1( u0_u13_u0_n148 ) , .ZN( u0_u13_u0_n90 ) );
  INV_X1 u0_u13_u0_U26 (.A( u0_u13_u0_n136 ) , .ZN( u0_u13_u0_n161 ) );
  NOR2_X1 u0_u13_u0_U27 (.A1( u0_u13_u0_n120 ) , .ZN( u0_u13_u0_n143 ) , .A2( u0_u13_u0_n167 ) );
  OAI221_X1 u0_u13_u0_U28 (.C1( u0_u13_u0_n112 ) , .ZN( u0_u13_u0_n120 ) , .B1( u0_u13_u0_n138 ) , .B2( u0_u13_u0_n141 ) , .C2( u0_u13_u0_n147 ) , .A( u0_u13_u0_n172 ) );
  AOI211_X1 u0_u13_u0_U29 (.B( u0_u13_u0_n115 ) , .A( u0_u13_u0_n116 ) , .C2( u0_u13_u0_n117 ) , .C1( u0_u13_u0_n118 ) , .ZN( u0_u13_u0_n119 ) );
  INV_X1 u0_u13_u0_U3 (.A( u0_u13_u0_n113 ) , .ZN( u0_u13_u0_n166 ) );
  AOI22_X1 u0_u13_u0_U30 (.B2( u0_u13_u0_n109 ) , .A2( u0_u13_u0_n110 ) , .ZN( u0_u13_u0_n111 ) , .B1( u0_u13_u0_n118 ) , .A1( u0_u13_u0_n160 ) );
  INV_X1 u0_u13_u0_U31 (.A( u0_u13_u0_n118 ) , .ZN( u0_u13_u0_n158 ) );
  AOI21_X1 u0_u13_u0_U32 (.ZN( u0_u13_u0_n104 ) , .B1( u0_u13_u0_n107 ) , .B2( u0_u13_u0_n141 ) , .A( u0_u13_u0_n144 ) );
  AOI21_X1 u0_u13_u0_U33 (.B1( u0_u13_u0_n127 ) , .B2( u0_u13_u0_n129 ) , .A( u0_u13_u0_n138 ) , .ZN( u0_u13_u0_n96 ) );
  AOI21_X1 u0_u13_u0_U34 (.ZN( u0_u13_u0_n116 ) , .B2( u0_u13_u0_n142 ) , .A( u0_u13_u0_n144 ) , .B1( u0_u13_u0_n166 ) );
  NAND2_X1 u0_u13_u0_U35 (.A1( u0_u13_u0_n100 ) , .A2( u0_u13_u0_n103 ) , .ZN( u0_u13_u0_n125 ) );
  NAND2_X1 u0_u13_u0_U36 (.A1( u0_u13_u0_n101 ) , .A2( u0_u13_u0_n102 ) , .ZN( u0_u13_u0_n150 ) );
  INV_X1 u0_u13_u0_U37 (.A( u0_u13_u0_n138 ) , .ZN( u0_u13_u0_n160 ) );
  NAND2_X1 u0_u13_u0_U38 (.A1( u0_u13_u0_n102 ) , .ZN( u0_u13_u0_n128 ) , .A2( u0_u13_u0_n95 ) );
  NAND2_X1 u0_u13_u0_U39 (.A1( u0_u13_u0_n100 ) , .ZN( u0_u13_u0_n129 ) , .A2( u0_u13_u0_n95 ) );
  AOI21_X1 u0_u13_u0_U4 (.B1( u0_u13_u0_n114 ) , .ZN( u0_u13_u0_n115 ) , .B2( u0_u13_u0_n129 ) , .A( u0_u13_u0_n161 ) );
  NAND2_X1 u0_u13_u0_U40 (.A2( u0_u13_u0_n100 ) , .ZN( u0_u13_u0_n131 ) , .A1( u0_u13_u0_n92 ) );
  NAND2_X1 u0_u13_u0_U41 (.A2( u0_u13_u0_n100 ) , .A1( u0_u13_u0_n101 ) , .ZN( u0_u13_u0_n139 ) );
  NAND2_X1 u0_u13_u0_U42 (.ZN( u0_u13_u0_n148 ) , .A1( u0_u13_u0_n93 ) , .A2( u0_u13_u0_n95 ) );
  NAND2_X1 u0_u13_u0_U43 (.A2( u0_u13_u0_n102 ) , .A1( u0_u13_u0_n103 ) , .ZN( u0_u13_u0_n149 ) );
  NAND2_X1 u0_u13_u0_U44 (.A2( u0_u13_u0_n102 ) , .ZN( u0_u13_u0_n114 ) , .A1( u0_u13_u0_n92 ) );
  NAND2_X1 u0_u13_u0_U45 (.A2( u0_u13_u0_n101 ) , .ZN( u0_u13_u0_n121 ) , .A1( u0_u13_u0_n93 ) );
  NAND2_X1 u0_u13_u0_U46 (.ZN( u0_u13_u0_n112 ) , .A2( u0_u13_u0_n92 ) , .A1( u0_u13_u0_n93 ) );
  OR3_X1 u0_u13_u0_U47 (.A3( u0_u13_u0_n152 ) , .A2( u0_u13_u0_n153 ) , .A1( u0_u13_u0_n154 ) , .ZN( u0_u13_u0_n155 ) );
  AOI21_X1 u0_u13_u0_U48 (.B2( u0_u13_u0_n150 ) , .B1( u0_u13_u0_n151 ) , .ZN( u0_u13_u0_n152 ) , .A( u0_u13_u0_n158 ) );
  AOI21_X1 u0_u13_u0_U49 (.A( u0_u13_u0_n144 ) , .B2( u0_u13_u0_n145 ) , .B1( u0_u13_u0_n146 ) , .ZN( u0_u13_u0_n154 ) );
  AOI21_X1 u0_u13_u0_U5 (.B2( u0_u13_u0_n131 ) , .ZN( u0_u13_u0_n134 ) , .B1( u0_u13_u0_n151 ) , .A( u0_u13_u0_n158 ) );
  AOI21_X1 u0_u13_u0_U50 (.A( u0_u13_u0_n147 ) , .B2( u0_u13_u0_n148 ) , .B1( u0_u13_u0_n149 ) , .ZN( u0_u13_u0_n153 ) );
  INV_X1 u0_u13_u0_U51 (.ZN( u0_u13_u0_n171 ) , .A( u0_u13_u0_n99 ) );
  OAI211_X1 u0_u13_u0_U52 (.C2( u0_u13_u0_n140 ) , .C1( u0_u13_u0_n161 ) , .A( u0_u13_u0_n169 ) , .B( u0_u13_u0_n98 ) , .ZN( u0_u13_u0_n99 ) );
  AOI211_X1 u0_u13_u0_U53 (.C1( u0_u13_u0_n118 ) , .A( u0_u13_u0_n123 ) , .B( u0_u13_u0_n96 ) , .C2( u0_u13_u0_n97 ) , .ZN( u0_u13_u0_n98 ) );
  INV_X1 u0_u13_u0_U54 (.ZN( u0_u13_u0_n169 ) , .A( u0_u13_u0_n91 ) );
  NOR2_X1 u0_u13_u0_U55 (.A2( u0_u13_X_6 ) , .ZN( u0_u13_u0_n100 ) , .A1( u0_u13_u0_n162 ) );
  NOR2_X1 u0_u13_u0_U56 (.A2( u0_u13_X_4 ) , .A1( u0_u13_X_5 ) , .ZN( u0_u13_u0_n118 ) );
  NOR2_X1 u0_u13_u0_U57 (.A2( u0_u13_X_2 ) , .ZN( u0_u13_u0_n103 ) , .A1( u0_u13_u0_n164 ) );
  NOR2_X1 u0_u13_u0_U58 (.A2( u0_u13_X_1 ) , .A1( u0_u13_X_2 ) , .ZN( u0_u13_u0_n92 ) );
  NOR2_X1 u0_u13_u0_U59 (.A2( u0_u13_X_1 ) , .ZN( u0_u13_u0_n101 ) , .A1( u0_u13_u0_n163 ) );
  NOR2_X1 u0_u13_u0_U6 (.A1( u0_u13_u0_n108 ) , .ZN( u0_u13_u0_n123 ) , .A2( u0_u13_u0_n158 ) );
  NAND2_X1 u0_u13_u0_U60 (.A2( u0_u13_X_4 ) , .A1( u0_u13_X_5 ) , .ZN( u0_u13_u0_n144 ) );
  NOR2_X1 u0_u13_u0_U61 (.A2( u0_u13_X_5 ) , .ZN( u0_u13_u0_n136 ) , .A1( u0_u13_u0_n159 ) );
  NAND2_X1 u0_u13_u0_U62 (.A1( u0_u13_X_5 ) , .ZN( u0_u13_u0_n138 ) , .A2( u0_u13_u0_n159 ) );
  AND2_X1 u0_u13_u0_U63 (.A2( u0_u13_X_3 ) , .A1( u0_u13_X_6 ) , .ZN( u0_u13_u0_n102 ) );
  AND2_X1 u0_u13_u0_U64 (.A1( u0_u13_X_6 ) , .A2( u0_u13_u0_n162 ) , .ZN( u0_u13_u0_n93 ) );
  INV_X1 u0_u13_u0_U65 (.A( u0_u13_X_4 ) , .ZN( u0_u13_u0_n159 ) );
  INV_X1 u0_u13_u0_U66 (.A( u0_u13_X_1 ) , .ZN( u0_u13_u0_n164 ) );
  INV_X1 u0_u13_u0_U67 (.A( u0_u13_X_2 ) , .ZN( u0_u13_u0_n163 ) );
  INV_X1 u0_u13_u0_U68 (.A( u0_u13_u0_n126 ) , .ZN( u0_u13_u0_n168 ) );
  AOI211_X1 u0_u13_u0_U69 (.B( u0_u13_u0_n133 ) , .A( u0_u13_u0_n134 ) , .C2( u0_u13_u0_n135 ) , .C1( u0_u13_u0_n136 ) , .ZN( u0_u13_u0_n137 ) );
  OAI21_X1 u0_u13_u0_U7 (.B1( u0_u13_u0_n150 ) , .B2( u0_u13_u0_n158 ) , .A( u0_u13_u0_n172 ) , .ZN( u0_u13_u0_n89 ) );
  INV_X1 u0_u13_u0_U70 (.ZN( u0_u13_u0_n174 ) , .A( u0_u13_u0_n89 ) );
  AOI211_X1 u0_u13_u0_U71 (.B( u0_u13_u0_n104 ) , .A( u0_u13_u0_n105 ) , .ZN( u0_u13_u0_n106 ) , .C2( u0_u13_u0_n113 ) , .C1( u0_u13_u0_n160 ) );
  OR4_X1 u0_u13_u0_U72 (.ZN( u0_out13_17 ) , .A4( u0_u13_u0_n122 ) , .A2( u0_u13_u0_n123 ) , .A1( u0_u13_u0_n124 ) , .A3( u0_u13_u0_n170 ) );
  AOI21_X1 u0_u13_u0_U73 (.B2( u0_u13_u0_n107 ) , .ZN( u0_u13_u0_n124 ) , .B1( u0_u13_u0_n128 ) , .A( u0_u13_u0_n161 ) );
  INV_X1 u0_u13_u0_U74 (.A( u0_u13_u0_n111 ) , .ZN( u0_u13_u0_n170 ) );
  OR4_X1 u0_u13_u0_U75 (.ZN( u0_out13_31 ) , .A4( u0_u13_u0_n155 ) , .A2( u0_u13_u0_n156 ) , .A1( u0_u13_u0_n157 ) , .A3( u0_u13_u0_n173 ) );
  AOI21_X1 u0_u13_u0_U76 (.A( u0_u13_u0_n138 ) , .B2( u0_u13_u0_n139 ) , .B1( u0_u13_u0_n140 ) , .ZN( u0_u13_u0_n157 ) );
  AOI21_X1 u0_u13_u0_U77 (.B2( u0_u13_u0_n141 ) , .B1( u0_u13_u0_n142 ) , .ZN( u0_u13_u0_n156 ) , .A( u0_u13_u0_n161 ) );
  AOI21_X1 u0_u13_u0_U78 (.B1( u0_u13_u0_n132 ) , .ZN( u0_u13_u0_n133 ) , .A( u0_u13_u0_n144 ) , .B2( u0_u13_u0_n166 ) );
  OAI22_X1 u0_u13_u0_U79 (.ZN( u0_u13_u0_n105 ) , .A2( u0_u13_u0_n132 ) , .B1( u0_u13_u0_n146 ) , .A1( u0_u13_u0_n147 ) , .B2( u0_u13_u0_n161 ) );
  AND2_X1 u0_u13_u0_U8 (.A1( u0_u13_u0_n114 ) , .A2( u0_u13_u0_n121 ) , .ZN( u0_u13_u0_n146 ) );
  NAND2_X1 u0_u13_u0_U80 (.ZN( u0_u13_u0_n110 ) , .A2( u0_u13_u0_n132 ) , .A1( u0_u13_u0_n145 ) );
  INV_X1 u0_u13_u0_U81 (.A( u0_u13_u0_n119 ) , .ZN( u0_u13_u0_n167 ) );
  NAND2_X1 u0_u13_u0_U82 (.A2( u0_u13_u0_n103 ) , .ZN( u0_u13_u0_n140 ) , .A1( u0_u13_u0_n94 ) );
  NAND2_X1 u0_u13_u0_U83 (.A1( u0_u13_u0_n101 ) , .ZN( u0_u13_u0_n130 ) , .A2( u0_u13_u0_n94 ) );
  NAND2_X1 u0_u13_u0_U84 (.ZN( u0_u13_u0_n108 ) , .A1( u0_u13_u0_n92 ) , .A2( u0_u13_u0_n94 ) );
  NAND2_X1 u0_u13_u0_U85 (.ZN( u0_u13_u0_n142 ) , .A1( u0_u13_u0_n94 ) , .A2( u0_u13_u0_n95 ) );
  INV_X1 u0_u13_u0_U86 (.A( u0_u13_X_3 ) , .ZN( u0_u13_u0_n162 ) );
  NOR2_X1 u0_u13_u0_U87 (.A2( u0_u13_X_3 ) , .A1( u0_u13_X_6 ) , .ZN( u0_u13_u0_n94 ) );
  NAND3_X1 u0_u13_u0_U88 (.ZN( u0_out13_23 ) , .A3( u0_u13_u0_n137 ) , .A1( u0_u13_u0_n168 ) , .A2( u0_u13_u0_n171 ) );
  NAND3_X1 u0_u13_u0_U89 (.A3( u0_u13_u0_n127 ) , .A2( u0_u13_u0_n128 ) , .ZN( u0_u13_u0_n135 ) , .A1( u0_u13_u0_n150 ) );
  AND2_X1 u0_u13_u0_U9 (.A1( u0_u13_u0_n131 ) , .ZN( u0_u13_u0_n141 ) , .A2( u0_u13_u0_n150 ) );
  NAND3_X1 u0_u13_u0_U90 (.ZN( u0_u13_u0_n117 ) , .A3( u0_u13_u0_n132 ) , .A2( u0_u13_u0_n139 ) , .A1( u0_u13_u0_n148 ) );
  NAND3_X1 u0_u13_u0_U91 (.ZN( u0_u13_u0_n109 ) , .A2( u0_u13_u0_n114 ) , .A3( u0_u13_u0_n140 ) , .A1( u0_u13_u0_n149 ) );
  NAND3_X1 u0_u13_u0_U92 (.ZN( u0_out13_9 ) , .A3( u0_u13_u0_n106 ) , .A2( u0_u13_u0_n171 ) , .A1( u0_u13_u0_n174 ) );
  NAND3_X1 u0_u13_u0_U93 (.A2( u0_u13_u0_n128 ) , .A1( u0_u13_u0_n132 ) , .A3( u0_u13_u0_n146 ) , .ZN( u0_u13_u0_n97 ) );
  AOI21_X1 u0_u13_u1_U10 (.B2( u0_u13_u1_n155 ) , .B1( u0_u13_u1_n156 ) , .ZN( u0_u13_u1_n157 ) , .A( u0_u13_u1_n174 ) );
  NAND3_X1 u0_u13_u1_U100 (.ZN( u0_u13_u1_n113 ) , .A1( u0_u13_u1_n120 ) , .A3( u0_u13_u1_n133 ) , .A2( u0_u13_u1_n155 ) );
  NAND2_X1 u0_u13_u1_U11 (.ZN( u0_u13_u1_n140 ) , .A2( u0_u13_u1_n150 ) , .A1( u0_u13_u1_n155 ) );
  NAND2_X1 u0_u13_u1_U12 (.A1( u0_u13_u1_n131 ) , .ZN( u0_u13_u1_n147 ) , .A2( u0_u13_u1_n153 ) );
  INV_X1 u0_u13_u1_U13 (.A( u0_u13_u1_n139 ) , .ZN( u0_u13_u1_n174 ) );
  OR4_X1 u0_u13_u1_U14 (.A4( u0_u13_u1_n106 ) , .A3( u0_u13_u1_n107 ) , .ZN( u0_u13_u1_n108 ) , .A1( u0_u13_u1_n117 ) , .A2( u0_u13_u1_n184 ) );
  AOI21_X1 u0_u13_u1_U15 (.ZN( u0_u13_u1_n106 ) , .A( u0_u13_u1_n112 ) , .B1( u0_u13_u1_n154 ) , .B2( u0_u13_u1_n156 ) );
  AOI21_X1 u0_u13_u1_U16 (.ZN( u0_u13_u1_n107 ) , .B1( u0_u13_u1_n134 ) , .B2( u0_u13_u1_n149 ) , .A( u0_u13_u1_n174 ) );
  INV_X1 u0_u13_u1_U17 (.A( u0_u13_u1_n101 ) , .ZN( u0_u13_u1_n184 ) );
  INV_X1 u0_u13_u1_U18 (.A( u0_u13_u1_n112 ) , .ZN( u0_u13_u1_n171 ) );
  NAND2_X1 u0_u13_u1_U19 (.ZN( u0_u13_u1_n141 ) , .A1( u0_u13_u1_n153 ) , .A2( u0_u13_u1_n156 ) );
  AND2_X1 u0_u13_u1_U20 (.A1( u0_u13_u1_n123 ) , .ZN( u0_u13_u1_n134 ) , .A2( u0_u13_u1_n161 ) );
  NAND2_X1 u0_u13_u1_U21 (.A2( u0_u13_u1_n115 ) , .A1( u0_u13_u1_n116 ) , .ZN( u0_u13_u1_n148 ) );
  NAND2_X1 u0_u13_u1_U22 (.A2( u0_u13_u1_n133 ) , .A1( u0_u13_u1_n135 ) , .ZN( u0_u13_u1_n159 ) );
  NAND2_X1 u0_u13_u1_U23 (.A2( u0_u13_u1_n115 ) , .A1( u0_u13_u1_n120 ) , .ZN( u0_u13_u1_n132 ) );
  INV_X1 u0_u13_u1_U24 (.A( u0_u13_u1_n154 ) , .ZN( u0_u13_u1_n178 ) );
  AOI22_X1 u0_u13_u1_U25 (.B2( u0_u13_u1_n113 ) , .A2( u0_u13_u1_n114 ) , .ZN( u0_u13_u1_n125 ) , .A1( u0_u13_u1_n171 ) , .B1( u0_u13_u1_n173 ) );
  NAND2_X1 u0_u13_u1_U26 (.ZN( u0_u13_u1_n114 ) , .A1( u0_u13_u1_n134 ) , .A2( u0_u13_u1_n156 ) );
  INV_X1 u0_u13_u1_U27 (.A( u0_u13_u1_n151 ) , .ZN( u0_u13_u1_n183 ) );
  AND2_X1 u0_u13_u1_U28 (.A1( u0_u13_u1_n129 ) , .A2( u0_u13_u1_n133 ) , .ZN( u0_u13_u1_n149 ) );
  INV_X1 u0_u13_u1_U29 (.A( u0_u13_u1_n131 ) , .ZN( u0_u13_u1_n180 ) );
  INV_X1 u0_u13_u1_U3 (.A( u0_u13_u1_n159 ) , .ZN( u0_u13_u1_n182 ) );
  OAI221_X1 u0_u13_u1_U30 (.A( u0_u13_u1_n119 ) , .C2( u0_u13_u1_n129 ) , .ZN( u0_u13_u1_n138 ) , .B2( u0_u13_u1_n152 ) , .C1( u0_u13_u1_n174 ) , .B1( u0_u13_u1_n187 ) );
  INV_X1 u0_u13_u1_U31 (.A( u0_u13_u1_n148 ) , .ZN( u0_u13_u1_n187 ) );
  AOI211_X1 u0_u13_u1_U32 (.B( u0_u13_u1_n117 ) , .A( u0_u13_u1_n118 ) , .ZN( u0_u13_u1_n119 ) , .C2( u0_u13_u1_n146 ) , .C1( u0_u13_u1_n159 ) );
  NOR2_X1 u0_u13_u1_U33 (.A1( u0_u13_u1_n168 ) , .A2( u0_u13_u1_n176 ) , .ZN( u0_u13_u1_n98 ) );
  AOI211_X1 u0_u13_u1_U34 (.B( u0_u13_u1_n162 ) , .A( u0_u13_u1_n163 ) , .C2( u0_u13_u1_n164 ) , .ZN( u0_u13_u1_n165 ) , .C1( u0_u13_u1_n171 ) );
  AOI21_X1 u0_u13_u1_U35 (.A( u0_u13_u1_n160 ) , .B2( u0_u13_u1_n161 ) , .ZN( u0_u13_u1_n162 ) , .B1( u0_u13_u1_n182 ) );
  OR2_X1 u0_u13_u1_U36 (.A2( u0_u13_u1_n157 ) , .A1( u0_u13_u1_n158 ) , .ZN( u0_u13_u1_n163 ) );
  OAI21_X1 u0_u13_u1_U37 (.B2( u0_u13_u1_n123 ) , .ZN( u0_u13_u1_n145 ) , .B1( u0_u13_u1_n160 ) , .A( u0_u13_u1_n185 ) );
  INV_X1 u0_u13_u1_U38 (.A( u0_u13_u1_n122 ) , .ZN( u0_u13_u1_n185 ) );
  AOI21_X1 u0_u13_u1_U39 (.B2( u0_u13_u1_n120 ) , .B1( u0_u13_u1_n121 ) , .ZN( u0_u13_u1_n122 ) , .A( u0_u13_u1_n128 ) );
  AOI221_X1 u0_u13_u1_U4 (.A( u0_u13_u1_n138 ) , .C2( u0_u13_u1_n139 ) , .C1( u0_u13_u1_n140 ) , .B2( u0_u13_u1_n141 ) , .ZN( u0_u13_u1_n142 ) , .B1( u0_u13_u1_n175 ) );
  NAND2_X1 u0_u13_u1_U40 (.A1( u0_u13_u1_n128 ) , .ZN( u0_u13_u1_n146 ) , .A2( u0_u13_u1_n160 ) );
  NAND2_X1 u0_u13_u1_U41 (.A2( u0_u13_u1_n112 ) , .ZN( u0_u13_u1_n139 ) , .A1( u0_u13_u1_n152 ) );
  NAND2_X1 u0_u13_u1_U42 (.A1( u0_u13_u1_n105 ) , .ZN( u0_u13_u1_n156 ) , .A2( u0_u13_u1_n99 ) );
  AOI221_X1 u0_u13_u1_U43 (.B1( u0_u13_u1_n140 ) , .ZN( u0_u13_u1_n167 ) , .B2( u0_u13_u1_n172 ) , .C2( u0_u13_u1_n175 ) , .C1( u0_u13_u1_n178 ) , .A( u0_u13_u1_n188 ) );
  INV_X1 u0_u13_u1_U44 (.ZN( u0_u13_u1_n188 ) , .A( u0_u13_u1_n97 ) );
  AOI211_X1 u0_u13_u1_U45 (.A( u0_u13_u1_n118 ) , .C1( u0_u13_u1_n132 ) , .C2( u0_u13_u1_n139 ) , .B( u0_u13_u1_n96 ) , .ZN( u0_u13_u1_n97 ) );
  AOI21_X1 u0_u13_u1_U46 (.B2( u0_u13_u1_n121 ) , .B1( u0_u13_u1_n135 ) , .A( u0_u13_u1_n152 ) , .ZN( u0_u13_u1_n96 ) );
  NOR2_X1 u0_u13_u1_U47 (.ZN( u0_u13_u1_n117 ) , .A1( u0_u13_u1_n121 ) , .A2( u0_u13_u1_n160 ) );
  AOI21_X1 u0_u13_u1_U48 (.A( u0_u13_u1_n128 ) , .B2( u0_u13_u1_n129 ) , .ZN( u0_u13_u1_n130 ) , .B1( u0_u13_u1_n150 ) );
  NAND2_X1 u0_u13_u1_U49 (.ZN( u0_u13_u1_n112 ) , .A1( u0_u13_u1_n169 ) , .A2( u0_u13_u1_n170 ) );
  AOI211_X1 u0_u13_u1_U5 (.ZN( u0_u13_u1_n124 ) , .A( u0_u13_u1_n138 ) , .C2( u0_u13_u1_n139 ) , .B( u0_u13_u1_n145 ) , .C1( u0_u13_u1_n147 ) );
  NAND2_X1 u0_u13_u1_U50 (.ZN( u0_u13_u1_n129 ) , .A2( u0_u13_u1_n95 ) , .A1( u0_u13_u1_n98 ) );
  NAND2_X1 u0_u13_u1_U51 (.A1( u0_u13_u1_n102 ) , .ZN( u0_u13_u1_n154 ) , .A2( u0_u13_u1_n99 ) );
  NAND2_X1 u0_u13_u1_U52 (.A2( u0_u13_u1_n100 ) , .ZN( u0_u13_u1_n135 ) , .A1( u0_u13_u1_n99 ) );
  AOI21_X1 u0_u13_u1_U53 (.A( u0_u13_u1_n152 ) , .B2( u0_u13_u1_n153 ) , .B1( u0_u13_u1_n154 ) , .ZN( u0_u13_u1_n158 ) );
  INV_X1 u0_u13_u1_U54 (.A( u0_u13_u1_n160 ) , .ZN( u0_u13_u1_n175 ) );
  NAND2_X1 u0_u13_u1_U55 (.A1( u0_u13_u1_n100 ) , .ZN( u0_u13_u1_n116 ) , .A2( u0_u13_u1_n95 ) );
  NAND2_X1 u0_u13_u1_U56 (.A1( u0_u13_u1_n102 ) , .ZN( u0_u13_u1_n131 ) , .A2( u0_u13_u1_n95 ) );
  NAND2_X1 u0_u13_u1_U57 (.A2( u0_u13_u1_n104 ) , .ZN( u0_u13_u1_n121 ) , .A1( u0_u13_u1_n98 ) );
  NAND2_X1 u0_u13_u1_U58 (.A1( u0_u13_u1_n103 ) , .ZN( u0_u13_u1_n153 ) , .A2( u0_u13_u1_n98 ) );
  NAND2_X1 u0_u13_u1_U59 (.A2( u0_u13_u1_n104 ) , .A1( u0_u13_u1_n105 ) , .ZN( u0_u13_u1_n133 ) );
  AOI22_X1 u0_u13_u1_U6 (.B2( u0_u13_u1_n136 ) , .A2( u0_u13_u1_n137 ) , .ZN( u0_u13_u1_n143 ) , .A1( u0_u13_u1_n171 ) , .B1( u0_u13_u1_n173 ) );
  NAND2_X1 u0_u13_u1_U60 (.ZN( u0_u13_u1_n150 ) , .A2( u0_u13_u1_n98 ) , .A1( u0_u13_u1_n99 ) );
  NAND2_X1 u0_u13_u1_U61 (.A1( u0_u13_u1_n105 ) , .ZN( u0_u13_u1_n155 ) , .A2( u0_u13_u1_n95 ) );
  OAI21_X1 u0_u13_u1_U62 (.ZN( u0_u13_u1_n109 ) , .B1( u0_u13_u1_n129 ) , .B2( u0_u13_u1_n160 ) , .A( u0_u13_u1_n167 ) );
  NAND2_X1 u0_u13_u1_U63 (.A2( u0_u13_u1_n100 ) , .A1( u0_u13_u1_n103 ) , .ZN( u0_u13_u1_n120 ) );
  NAND2_X1 u0_u13_u1_U64 (.A1( u0_u13_u1_n102 ) , .A2( u0_u13_u1_n104 ) , .ZN( u0_u13_u1_n115 ) );
  NAND2_X1 u0_u13_u1_U65 (.A2( u0_u13_u1_n100 ) , .A1( u0_u13_u1_n104 ) , .ZN( u0_u13_u1_n151 ) );
  NAND2_X1 u0_u13_u1_U66 (.A2( u0_u13_u1_n103 ) , .A1( u0_u13_u1_n105 ) , .ZN( u0_u13_u1_n161 ) );
  INV_X1 u0_u13_u1_U67 (.A( u0_u13_u1_n152 ) , .ZN( u0_u13_u1_n173 ) );
  INV_X1 u0_u13_u1_U68 (.A( u0_u13_u1_n128 ) , .ZN( u0_u13_u1_n172 ) );
  NAND2_X1 u0_u13_u1_U69 (.A2( u0_u13_u1_n102 ) , .A1( u0_u13_u1_n103 ) , .ZN( u0_u13_u1_n123 ) );
  INV_X1 u0_u13_u1_U7 (.A( u0_u13_u1_n147 ) , .ZN( u0_u13_u1_n181 ) );
  NOR2_X1 u0_u13_u1_U70 (.A2( u0_u13_X_7 ) , .A1( u0_u13_X_8 ) , .ZN( u0_u13_u1_n95 ) );
  NOR2_X1 u0_u13_u1_U71 (.A1( u0_u13_X_12 ) , .A2( u0_u13_X_9 ) , .ZN( u0_u13_u1_n100 ) );
  NOR2_X1 u0_u13_u1_U72 (.A2( u0_u13_X_8 ) , .A1( u0_u13_u1_n177 ) , .ZN( u0_u13_u1_n99 ) );
  NOR2_X1 u0_u13_u1_U73 (.A2( u0_u13_X_12 ) , .ZN( u0_u13_u1_n102 ) , .A1( u0_u13_u1_n176 ) );
  NOR2_X1 u0_u13_u1_U74 (.A2( u0_u13_X_9 ) , .ZN( u0_u13_u1_n105 ) , .A1( u0_u13_u1_n168 ) );
  NAND2_X1 u0_u13_u1_U75 (.A1( u0_u13_X_10 ) , .ZN( u0_u13_u1_n160 ) , .A2( u0_u13_u1_n169 ) );
  NAND2_X1 u0_u13_u1_U76 (.A2( u0_u13_X_10 ) , .A1( u0_u13_X_11 ) , .ZN( u0_u13_u1_n152 ) );
  NAND2_X1 u0_u13_u1_U77 (.A1( u0_u13_X_11 ) , .ZN( u0_u13_u1_n128 ) , .A2( u0_u13_u1_n170 ) );
  AND2_X1 u0_u13_u1_U78 (.A2( u0_u13_X_7 ) , .A1( u0_u13_X_8 ) , .ZN( u0_u13_u1_n104 ) );
  AND2_X1 u0_u13_u1_U79 (.A1( u0_u13_X_8 ) , .ZN( u0_u13_u1_n103 ) , .A2( u0_u13_u1_n177 ) );
  NOR2_X1 u0_u13_u1_U8 (.A1( u0_u13_u1_n112 ) , .A2( u0_u13_u1_n116 ) , .ZN( u0_u13_u1_n118 ) );
  INV_X1 u0_u13_u1_U80 (.A( u0_u13_X_10 ) , .ZN( u0_u13_u1_n170 ) );
  INV_X1 u0_u13_u1_U81 (.A( u0_u13_X_9 ) , .ZN( u0_u13_u1_n176 ) );
  INV_X1 u0_u13_u1_U82 (.A( u0_u13_X_11 ) , .ZN( u0_u13_u1_n169 ) );
  INV_X1 u0_u13_u1_U83 (.A( u0_u13_X_12 ) , .ZN( u0_u13_u1_n168 ) );
  INV_X1 u0_u13_u1_U84 (.A( u0_u13_X_7 ) , .ZN( u0_u13_u1_n177 ) );
  NAND4_X1 u0_u13_u1_U85 (.ZN( u0_out13_28 ) , .A4( u0_u13_u1_n124 ) , .A3( u0_u13_u1_n125 ) , .A2( u0_u13_u1_n126 ) , .A1( u0_u13_u1_n127 ) );
  OAI21_X1 u0_u13_u1_U86 (.ZN( u0_u13_u1_n127 ) , .B2( u0_u13_u1_n139 ) , .B1( u0_u13_u1_n175 ) , .A( u0_u13_u1_n183 ) );
  OAI21_X1 u0_u13_u1_U87 (.ZN( u0_u13_u1_n126 ) , .B2( u0_u13_u1_n140 ) , .A( u0_u13_u1_n146 ) , .B1( u0_u13_u1_n178 ) );
  NAND4_X1 u0_u13_u1_U88 (.ZN( u0_out13_18 ) , .A4( u0_u13_u1_n165 ) , .A3( u0_u13_u1_n166 ) , .A1( u0_u13_u1_n167 ) , .A2( u0_u13_u1_n186 ) );
  AOI22_X1 u0_u13_u1_U89 (.B2( u0_u13_u1_n146 ) , .B1( u0_u13_u1_n147 ) , .A2( u0_u13_u1_n148 ) , .ZN( u0_u13_u1_n166 ) , .A1( u0_u13_u1_n172 ) );
  OAI21_X1 u0_u13_u1_U9 (.ZN( u0_u13_u1_n101 ) , .B1( u0_u13_u1_n141 ) , .A( u0_u13_u1_n146 ) , .B2( u0_u13_u1_n183 ) );
  INV_X1 u0_u13_u1_U90 (.A( u0_u13_u1_n145 ) , .ZN( u0_u13_u1_n186 ) );
  NAND4_X1 u0_u13_u1_U91 (.ZN( u0_out13_2 ) , .A4( u0_u13_u1_n142 ) , .A3( u0_u13_u1_n143 ) , .A2( u0_u13_u1_n144 ) , .A1( u0_u13_u1_n179 ) );
  OAI21_X1 u0_u13_u1_U92 (.B2( u0_u13_u1_n132 ) , .ZN( u0_u13_u1_n144 ) , .A( u0_u13_u1_n146 ) , .B1( u0_u13_u1_n180 ) );
  INV_X1 u0_u13_u1_U93 (.A( u0_u13_u1_n130 ) , .ZN( u0_u13_u1_n179 ) );
  OR4_X1 u0_u13_u1_U94 (.ZN( u0_out13_13 ) , .A4( u0_u13_u1_n108 ) , .A3( u0_u13_u1_n109 ) , .A2( u0_u13_u1_n110 ) , .A1( u0_u13_u1_n111 ) );
  AOI21_X1 u0_u13_u1_U95 (.ZN( u0_u13_u1_n111 ) , .A( u0_u13_u1_n128 ) , .B2( u0_u13_u1_n131 ) , .B1( u0_u13_u1_n135 ) );
  AOI21_X1 u0_u13_u1_U96 (.ZN( u0_u13_u1_n110 ) , .A( u0_u13_u1_n116 ) , .B1( u0_u13_u1_n152 ) , .B2( u0_u13_u1_n160 ) );
  NAND3_X1 u0_u13_u1_U97 (.A3( u0_u13_u1_n149 ) , .A2( u0_u13_u1_n150 ) , .A1( u0_u13_u1_n151 ) , .ZN( u0_u13_u1_n164 ) );
  NAND3_X1 u0_u13_u1_U98 (.A3( u0_u13_u1_n134 ) , .A2( u0_u13_u1_n135 ) , .ZN( u0_u13_u1_n136 ) , .A1( u0_u13_u1_n151 ) );
  NAND3_X1 u0_u13_u1_U99 (.A1( u0_u13_u1_n133 ) , .ZN( u0_u13_u1_n137 ) , .A2( u0_u13_u1_n154 ) , .A3( u0_u13_u1_n181 ) );
  OAI22_X1 u0_u13_u2_U10 (.B1( u0_u13_u2_n151 ) , .A2( u0_u13_u2_n152 ) , .A1( u0_u13_u2_n153 ) , .ZN( u0_u13_u2_n160 ) , .B2( u0_u13_u2_n168 ) );
  NAND3_X1 u0_u13_u2_U100 (.A2( u0_u13_u2_n100 ) , .A1( u0_u13_u2_n104 ) , .A3( u0_u13_u2_n138 ) , .ZN( u0_u13_u2_n98 ) );
  NOR3_X1 u0_u13_u2_U11 (.A1( u0_u13_u2_n150 ) , .ZN( u0_u13_u2_n151 ) , .A3( u0_u13_u2_n175 ) , .A2( u0_u13_u2_n188 ) );
  AOI21_X1 u0_u13_u2_U12 (.B2( u0_u13_u2_n123 ) , .ZN( u0_u13_u2_n125 ) , .A( u0_u13_u2_n171 ) , .B1( u0_u13_u2_n184 ) );
  INV_X1 u0_u13_u2_U13 (.A( u0_u13_u2_n150 ) , .ZN( u0_u13_u2_n184 ) );
  AOI21_X1 u0_u13_u2_U14 (.ZN( u0_u13_u2_n144 ) , .B2( u0_u13_u2_n155 ) , .A( u0_u13_u2_n172 ) , .B1( u0_u13_u2_n185 ) );
  AOI21_X1 u0_u13_u2_U15 (.B2( u0_u13_u2_n143 ) , .ZN( u0_u13_u2_n145 ) , .B1( u0_u13_u2_n152 ) , .A( u0_u13_u2_n171 ) );
  INV_X1 u0_u13_u2_U16 (.A( u0_u13_u2_n156 ) , .ZN( u0_u13_u2_n171 ) );
  INV_X1 u0_u13_u2_U17 (.A( u0_u13_u2_n120 ) , .ZN( u0_u13_u2_n188 ) );
  NAND2_X1 u0_u13_u2_U18 (.A2( u0_u13_u2_n122 ) , .ZN( u0_u13_u2_n150 ) , .A1( u0_u13_u2_n152 ) );
  INV_X1 u0_u13_u2_U19 (.A( u0_u13_u2_n153 ) , .ZN( u0_u13_u2_n170 ) );
  INV_X1 u0_u13_u2_U20 (.A( u0_u13_u2_n137 ) , .ZN( u0_u13_u2_n173 ) );
  NAND2_X1 u0_u13_u2_U21 (.A1( u0_u13_u2_n132 ) , .A2( u0_u13_u2_n139 ) , .ZN( u0_u13_u2_n157 ) );
  INV_X1 u0_u13_u2_U22 (.A( u0_u13_u2_n113 ) , .ZN( u0_u13_u2_n178 ) );
  INV_X1 u0_u13_u2_U23 (.A( u0_u13_u2_n139 ) , .ZN( u0_u13_u2_n175 ) );
  INV_X1 u0_u13_u2_U24 (.A( u0_u13_u2_n155 ) , .ZN( u0_u13_u2_n181 ) );
  INV_X1 u0_u13_u2_U25 (.A( u0_u13_u2_n119 ) , .ZN( u0_u13_u2_n177 ) );
  INV_X1 u0_u13_u2_U26 (.A( u0_u13_u2_n116 ) , .ZN( u0_u13_u2_n180 ) );
  INV_X1 u0_u13_u2_U27 (.A( u0_u13_u2_n131 ) , .ZN( u0_u13_u2_n179 ) );
  INV_X1 u0_u13_u2_U28 (.A( u0_u13_u2_n154 ) , .ZN( u0_u13_u2_n176 ) );
  NAND2_X1 u0_u13_u2_U29 (.A2( u0_u13_u2_n116 ) , .A1( u0_u13_u2_n117 ) , .ZN( u0_u13_u2_n118 ) );
  NOR2_X1 u0_u13_u2_U3 (.ZN( u0_u13_u2_n121 ) , .A2( u0_u13_u2_n177 ) , .A1( u0_u13_u2_n180 ) );
  INV_X1 u0_u13_u2_U30 (.A( u0_u13_u2_n132 ) , .ZN( u0_u13_u2_n182 ) );
  INV_X1 u0_u13_u2_U31 (.A( u0_u13_u2_n158 ) , .ZN( u0_u13_u2_n183 ) );
  OAI21_X1 u0_u13_u2_U32 (.A( u0_u13_u2_n156 ) , .B1( u0_u13_u2_n157 ) , .ZN( u0_u13_u2_n158 ) , .B2( u0_u13_u2_n179 ) );
  NOR2_X1 u0_u13_u2_U33 (.ZN( u0_u13_u2_n156 ) , .A1( u0_u13_u2_n166 ) , .A2( u0_u13_u2_n169 ) );
  NOR2_X1 u0_u13_u2_U34 (.A2( u0_u13_u2_n114 ) , .ZN( u0_u13_u2_n137 ) , .A1( u0_u13_u2_n140 ) );
  NOR2_X1 u0_u13_u2_U35 (.A2( u0_u13_u2_n138 ) , .ZN( u0_u13_u2_n153 ) , .A1( u0_u13_u2_n156 ) );
  AOI211_X1 u0_u13_u2_U36 (.ZN( u0_u13_u2_n130 ) , .C1( u0_u13_u2_n138 ) , .C2( u0_u13_u2_n179 ) , .B( u0_u13_u2_n96 ) , .A( u0_u13_u2_n97 ) );
  OAI22_X1 u0_u13_u2_U37 (.B1( u0_u13_u2_n133 ) , .A2( u0_u13_u2_n137 ) , .A1( u0_u13_u2_n152 ) , .B2( u0_u13_u2_n168 ) , .ZN( u0_u13_u2_n97 ) );
  OAI221_X1 u0_u13_u2_U38 (.B1( u0_u13_u2_n113 ) , .C1( u0_u13_u2_n132 ) , .A( u0_u13_u2_n149 ) , .B2( u0_u13_u2_n171 ) , .C2( u0_u13_u2_n172 ) , .ZN( u0_u13_u2_n96 ) );
  OAI221_X1 u0_u13_u2_U39 (.A( u0_u13_u2_n115 ) , .C2( u0_u13_u2_n123 ) , .B2( u0_u13_u2_n143 ) , .B1( u0_u13_u2_n153 ) , .ZN( u0_u13_u2_n163 ) , .C1( u0_u13_u2_n168 ) );
  INV_X1 u0_u13_u2_U4 (.A( u0_u13_u2_n134 ) , .ZN( u0_u13_u2_n185 ) );
  OAI21_X1 u0_u13_u2_U40 (.A( u0_u13_u2_n114 ) , .ZN( u0_u13_u2_n115 ) , .B1( u0_u13_u2_n176 ) , .B2( u0_u13_u2_n178 ) );
  OAI221_X1 u0_u13_u2_U41 (.A( u0_u13_u2_n135 ) , .B2( u0_u13_u2_n136 ) , .B1( u0_u13_u2_n137 ) , .ZN( u0_u13_u2_n162 ) , .C2( u0_u13_u2_n167 ) , .C1( u0_u13_u2_n185 ) );
  AND3_X1 u0_u13_u2_U42 (.A3( u0_u13_u2_n131 ) , .A2( u0_u13_u2_n132 ) , .A1( u0_u13_u2_n133 ) , .ZN( u0_u13_u2_n136 ) );
  AOI22_X1 u0_u13_u2_U43 (.ZN( u0_u13_u2_n135 ) , .B1( u0_u13_u2_n140 ) , .A1( u0_u13_u2_n156 ) , .B2( u0_u13_u2_n180 ) , .A2( u0_u13_u2_n188 ) );
  AOI21_X1 u0_u13_u2_U44 (.ZN( u0_u13_u2_n149 ) , .B1( u0_u13_u2_n173 ) , .B2( u0_u13_u2_n188 ) , .A( u0_u13_u2_n95 ) );
  AND3_X1 u0_u13_u2_U45 (.A2( u0_u13_u2_n100 ) , .A1( u0_u13_u2_n104 ) , .A3( u0_u13_u2_n156 ) , .ZN( u0_u13_u2_n95 ) );
  OAI21_X1 u0_u13_u2_U46 (.A( u0_u13_u2_n141 ) , .B2( u0_u13_u2_n142 ) , .ZN( u0_u13_u2_n146 ) , .B1( u0_u13_u2_n153 ) );
  OAI21_X1 u0_u13_u2_U47 (.A( u0_u13_u2_n140 ) , .ZN( u0_u13_u2_n141 ) , .B1( u0_u13_u2_n176 ) , .B2( u0_u13_u2_n177 ) );
  NOR3_X1 u0_u13_u2_U48 (.ZN( u0_u13_u2_n142 ) , .A3( u0_u13_u2_n175 ) , .A2( u0_u13_u2_n178 ) , .A1( u0_u13_u2_n181 ) );
  OAI21_X1 u0_u13_u2_U49 (.A( u0_u13_u2_n101 ) , .B2( u0_u13_u2_n121 ) , .B1( u0_u13_u2_n153 ) , .ZN( u0_u13_u2_n164 ) );
  NOR4_X1 u0_u13_u2_U5 (.A4( u0_u13_u2_n124 ) , .A3( u0_u13_u2_n125 ) , .A2( u0_u13_u2_n126 ) , .A1( u0_u13_u2_n127 ) , .ZN( u0_u13_u2_n128 ) );
  NAND2_X1 u0_u13_u2_U50 (.A2( u0_u13_u2_n100 ) , .A1( u0_u13_u2_n107 ) , .ZN( u0_u13_u2_n155 ) );
  NAND2_X1 u0_u13_u2_U51 (.A2( u0_u13_u2_n105 ) , .A1( u0_u13_u2_n108 ) , .ZN( u0_u13_u2_n143 ) );
  NAND2_X1 u0_u13_u2_U52 (.A1( u0_u13_u2_n104 ) , .A2( u0_u13_u2_n106 ) , .ZN( u0_u13_u2_n152 ) );
  NAND2_X1 u0_u13_u2_U53 (.A1( u0_u13_u2_n100 ) , .A2( u0_u13_u2_n105 ) , .ZN( u0_u13_u2_n132 ) );
  INV_X1 u0_u13_u2_U54 (.A( u0_u13_u2_n140 ) , .ZN( u0_u13_u2_n168 ) );
  INV_X1 u0_u13_u2_U55 (.A( u0_u13_u2_n138 ) , .ZN( u0_u13_u2_n167 ) );
  NAND2_X1 u0_u13_u2_U56 (.A1( u0_u13_u2_n102 ) , .A2( u0_u13_u2_n106 ) , .ZN( u0_u13_u2_n113 ) );
  NAND2_X1 u0_u13_u2_U57 (.A1( u0_u13_u2_n106 ) , .A2( u0_u13_u2_n107 ) , .ZN( u0_u13_u2_n131 ) );
  NAND2_X1 u0_u13_u2_U58 (.A1( u0_u13_u2_n103 ) , .A2( u0_u13_u2_n107 ) , .ZN( u0_u13_u2_n139 ) );
  NAND2_X1 u0_u13_u2_U59 (.A1( u0_u13_u2_n103 ) , .A2( u0_u13_u2_n105 ) , .ZN( u0_u13_u2_n133 ) );
  AOI21_X1 u0_u13_u2_U6 (.B2( u0_u13_u2_n119 ) , .ZN( u0_u13_u2_n127 ) , .A( u0_u13_u2_n137 ) , .B1( u0_u13_u2_n155 ) );
  NAND2_X1 u0_u13_u2_U60 (.A1( u0_u13_u2_n102 ) , .A2( u0_u13_u2_n103 ) , .ZN( u0_u13_u2_n154 ) );
  NAND2_X1 u0_u13_u2_U61 (.A2( u0_u13_u2_n103 ) , .A1( u0_u13_u2_n104 ) , .ZN( u0_u13_u2_n119 ) );
  NAND2_X1 u0_u13_u2_U62 (.A2( u0_u13_u2_n107 ) , .A1( u0_u13_u2_n108 ) , .ZN( u0_u13_u2_n123 ) );
  NAND2_X1 u0_u13_u2_U63 (.A1( u0_u13_u2_n104 ) , .A2( u0_u13_u2_n108 ) , .ZN( u0_u13_u2_n122 ) );
  INV_X1 u0_u13_u2_U64 (.A( u0_u13_u2_n114 ) , .ZN( u0_u13_u2_n172 ) );
  NAND2_X1 u0_u13_u2_U65 (.A2( u0_u13_u2_n100 ) , .A1( u0_u13_u2_n102 ) , .ZN( u0_u13_u2_n116 ) );
  NAND2_X1 u0_u13_u2_U66 (.A1( u0_u13_u2_n102 ) , .A2( u0_u13_u2_n108 ) , .ZN( u0_u13_u2_n120 ) );
  NAND2_X1 u0_u13_u2_U67 (.A2( u0_u13_u2_n105 ) , .A1( u0_u13_u2_n106 ) , .ZN( u0_u13_u2_n117 ) );
  INV_X1 u0_u13_u2_U68 (.ZN( u0_u13_u2_n187 ) , .A( u0_u13_u2_n99 ) );
  OAI21_X1 u0_u13_u2_U69 (.B1( u0_u13_u2_n137 ) , .B2( u0_u13_u2_n143 ) , .A( u0_u13_u2_n98 ) , .ZN( u0_u13_u2_n99 ) );
  AOI21_X1 u0_u13_u2_U7 (.ZN( u0_u13_u2_n124 ) , .B1( u0_u13_u2_n131 ) , .B2( u0_u13_u2_n143 ) , .A( u0_u13_u2_n172 ) );
  NOR2_X1 u0_u13_u2_U70 (.A2( u0_u13_X_16 ) , .ZN( u0_u13_u2_n140 ) , .A1( u0_u13_u2_n166 ) );
  NOR2_X1 u0_u13_u2_U71 (.A2( u0_u13_X_13 ) , .A1( u0_u13_X_14 ) , .ZN( u0_u13_u2_n100 ) );
  NOR2_X1 u0_u13_u2_U72 (.A2( u0_u13_X_16 ) , .A1( u0_u13_X_17 ) , .ZN( u0_u13_u2_n138 ) );
  NOR2_X1 u0_u13_u2_U73 (.A2( u0_u13_X_15 ) , .A1( u0_u13_X_18 ) , .ZN( u0_u13_u2_n104 ) );
  NOR2_X1 u0_u13_u2_U74 (.A2( u0_u13_X_14 ) , .ZN( u0_u13_u2_n103 ) , .A1( u0_u13_u2_n174 ) );
  NOR2_X1 u0_u13_u2_U75 (.A2( u0_u13_X_15 ) , .ZN( u0_u13_u2_n102 ) , .A1( u0_u13_u2_n165 ) );
  NOR2_X1 u0_u13_u2_U76 (.A2( u0_u13_X_17 ) , .ZN( u0_u13_u2_n114 ) , .A1( u0_u13_u2_n169 ) );
  AND2_X1 u0_u13_u2_U77 (.A1( u0_u13_X_15 ) , .ZN( u0_u13_u2_n105 ) , .A2( u0_u13_u2_n165 ) );
  AND2_X1 u0_u13_u2_U78 (.A2( u0_u13_X_15 ) , .A1( u0_u13_X_18 ) , .ZN( u0_u13_u2_n107 ) );
  AND2_X1 u0_u13_u2_U79 (.A1( u0_u13_X_14 ) , .ZN( u0_u13_u2_n106 ) , .A2( u0_u13_u2_n174 ) );
  AOI21_X1 u0_u13_u2_U8 (.B2( u0_u13_u2_n120 ) , .B1( u0_u13_u2_n121 ) , .ZN( u0_u13_u2_n126 ) , .A( u0_u13_u2_n167 ) );
  AND2_X1 u0_u13_u2_U80 (.A1( u0_u13_X_13 ) , .A2( u0_u13_X_14 ) , .ZN( u0_u13_u2_n108 ) );
  INV_X1 u0_u13_u2_U81 (.A( u0_u13_X_16 ) , .ZN( u0_u13_u2_n169 ) );
  INV_X1 u0_u13_u2_U82 (.A( u0_u13_X_17 ) , .ZN( u0_u13_u2_n166 ) );
  INV_X1 u0_u13_u2_U83 (.A( u0_u13_X_13 ) , .ZN( u0_u13_u2_n174 ) );
  INV_X1 u0_u13_u2_U84 (.A( u0_u13_X_18 ) , .ZN( u0_u13_u2_n165 ) );
  NAND4_X1 u0_u13_u2_U85 (.ZN( u0_out13_30 ) , .A4( u0_u13_u2_n147 ) , .A3( u0_u13_u2_n148 ) , .A2( u0_u13_u2_n149 ) , .A1( u0_u13_u2_n187 ) );
  NOR3_X1 u0_u13_u2_U86 (.A3( u0_u13_u2_n144 ) , .A2( u0_u13_u2_n145 ) , .A1( u0_u13_u2_n146 ) , .ZN( u0_u13_u2_n147 ) );
  AOI21_X1 u0_u13_u2_U87 (.B2( u0_u13_u2_n138 ) , .ZN( u0_u13_u2_n148 ) , .A( u0_u13_u2_n162 ) , .B1( u0_u13_u2_n182 ) );
  NAND4_X1 u0_u13_u2_U88 (.ZN( u0_out13_24 ) , .A4( u0_u13_u2_n111 ) , .A3( u0_u13_u2_n112 ) , .A1( u0_u13_u2_n130 ) , .A2( u0_u13_u2_n187 ) );
  AOI221_X1 u0_u13_u2_U89 (.A( u0_u13_u2_n109 ) , .B1( u0_u13_u2_n110 ) , .ZN( u0_u13_u2_n111 ) , .C1( u0_u13_u2_n134 ) , .C2( u0_u13_u2_n170 ) , .B2( u0_u13_u2_n173 ) );
  OAI22_X1 u0_u13_u2_U9 (.ZN( u0_u13_u2_n109 ) , .A2( u0_u13_u2_n113 ) , .B2( u0_u13_u2_n133 ) , .B1( u0_u13_u2_n167 ) , .A1( u0_u13_u2_n168 ) );
  AOI21_X1 u0_u13_u2_U90 (.ZN( u0_u13_u2_n112 ) , .B2( u0_u13_u2_n156 ) , .A( u0_u13_u2_n164 ) , .B1( u0_u13_u2_n181 ) );
  NAND4_X1 u0_u13_u2_U91 (.ZN( u0_out13_16 ) , .A4( u0_u13_u2_n128 ) , .A3( u0_u13_u2_n129 ) , .A1( u0_u13_u2_n130 ) , .A2( u0_u13_u2_n186 ) );
  AOI22_X1 u0_u13_u2_U92 (.A2( u0_u13_u2_n118 ) , .ZN( u0_u13_u2_n129 ) , .A1( u0_u13_u2_n140 ) , .B1( u0_u13_u2_n157 ) , .B2( u0_u13_u2_n170 ) );
  INV_X1 u0_u13_u2_U93 (.A( u0_u13_u2_n163 ) , .ZN( u0_u13_u2_n186 ) );
  OR4_X1 u0_u13_u2_U94 (.ZN( u0_out13_6 ) , .A4( u0_u13_u2_n161 ) , .A3( u0_u13_u2_n162 ) , .A2( u0_u13_u2_n163 ) , .A1( u0_u13_u2_n164 ) );
  OR3_X1 u0_u13_u2_U95 (.A2( u0_u13_u2_n159 ) , .A1( u0_u13_u2_n160 ) , .ZN( u0_u13_u2_n161 ) , .A3( u0_u13_u2_n183 ) );
  AOI21_X1 u0_u13_u2_U96 (.B2( u0_u13_u2_n154 ) , .B1( u0_u13_u2_n155 ) , .ZN( u0_u13_u2_n159 ) , .A( u0_u13_u2_n167 ) );
  NAND3_X1 u0_u13_u2_U97 (.A2( u0_u13_u2_n117 ) , .A1( u0_u13_u2_n122 ) , .A3( u0_u13_u2_n123 ) , .ZN( u0_u13_u2_n134 ) );
  NAND3_X1 u0_u13_u2_U98 (.ZN( u0_u13_u2_n110 ) , .A2( u0_u13_u2_n131 ) , .A3( u0_u13_u2_n139 ) , .A1( u0_u13_u2_n154 ) );
  NAND3_X1 u0_u13_u2_U99 (.A2( u0_u13_u2_n100 ) , .ZN( u0_u13_u2_n101 ) , .A1( u0_u13_u2_n104 ) , .A3( u0_u13_u2_n114 ) );
  OAI22_X1 u0_u13_u3_U10 (.B1( u0_u13_u3_n113 ) , .A2( u0_u13_u3_n135 ) , .A1( u0_u13_u3_n150 ) , .B2( u0_u13_u3_n164 ) , .ZN( u0_u13_u3_n98 ) );
  OAI211_X1 u0_u13_u3_U11 (.B( u0_u13_u3_n106 ) , .ZN( u0_u13_u3_n119 ) , .C2( u0_u13_u3_n128 ) , .C1( u0_u13_u3_n167 ) , .A( u0_u13_u3_n181 ) );
  AOI221_X1 u0_u13_u3_U12 (.C1( u0_u13_u3_n105 ) , .ZN( u0_u13_u3_n106 ) , .A( u0_u13_u3_n131 ) , .B2( u0_u13_u3_n132 ) , .C2( u0_u13_u3_n133 ) , .B1( u0_u13_u3_n169 ) );
  INV_X1 u0_u13_u3_U13 (.ZN( u0_u13_u3_n181 ) , .A( u0_u13_u3_n98 ) );
  NAND2_X1 u0_u13_u3_U14 (.ZN( u0_u13_u3_n105 ) , .A2( u0_u13_u3_n130 ) , .A1( u0_u13_u3_n155 ) );
  AOI22_X1 u0_u13_u3_U15 (.B1( u0_u13_u3_n115 ) , .A2( u0_u13_u3_n116 ) , .ZN( u0_u13_u3_n123 ) , .B2( u0_u13_u3_n133 ) , .A1( u0_u13_u3_n169 ) );
  NAND2_X1 u0_u13_u3_U16 (.ZN( u0_u13_u3_n116 ) , .A2( u0_u13_u3_n151 ) , .A1( u0_u13_u3_n182 ) );
  NOR2_X1 u0_u13_u3_U17 (.ZN( u0_u13_u3_n126 ) , .A2( u0_u13_u3_n150 ) , .A1( u0_u13_u3_n164 ) );
  AOI21_X1 u0_u13_u3_U18 (.ZN( u0_u13_u3_n112 ) , .B2( u0_u13_u3_n146 ) , .B1( u0_u13_u3_n155 ) , .A( u0_u13_u3_n167 ) );
  NAND2_X1 u0_u13_u3_U19 (.A1( u0_u13_u3_n135 ) , .ZN( u0_u13_u3_n142 ) , .A2( u0_u13_u3_n164 ) );
  NAND2_X1 u0_u13_u3_U20 (.ZN( u0_u13_u3_n132 ) , .A2( u0_u13_u3_n152 ) , .A1( u0_u13_u3_n156 ) );
  AND2_X1 u0_u13_u3_U21 (.A2( u0_u13_u3_n113 ) , .A1( u0_u13_u3_n114 ) , .ZN( u0_u13_u3_n151 ) );
  INV_X1 u0_u13_u3_U22 (.A( u0_u13_u3_n133 ) , .ZN( u0_u13_u3_n165 ) );
  INV_X1 u0_u13_u3_U23 (.A( u0_u13_u3_n135 ) , .ZN( u0_u13_u3_n170 ) );
  NAND2_X1 u0_u13_u3_U24 (.A1( u0_u13_u3_n107 ) , .A2( u0_u13_u3_n108 ) , .ZN( u0_u13_u3_n140 ) );
  NAND2_X1 u0_u13_u3_U25 (.ZN( u0_u13_u3_n117 ) , .A1( u0_u13_u3_n124 ) , .A2( u0_u13_u3_n148 ) );
  NAND2_X1 u0_u13_u3_U26 (.ZN( u0_u13_u3_n143 ) , .A1( u0_u13_u3_n165 ) , .A2( u0_u13_u3_n167 ) );
  INV_X1 u0_u13_u3_U27 (.A( u0_u13_u3_n130 ) , .ZN( u0_u13_u3_n177 ) );
  INV_X1 u0_u13_u3_U28 (.A( u0_u13_u3_n128 ) , .ZN( u0_u13_u3_n176 ) );
  INV_X1 u0_u13_u3_U29 (.A( u0_u13_u3_n155 ) , .ZN( u0_u13_u3_n174 ) );
  INV_X1 u0_u13_u3_U3 (.A( u0_u13_u3_n129 ) , .ZN( u0_u13_u3_n183 ) );
  INV_X1 u0_u13_u3_U30 (.A( u0_u13_u3_n139 ) , .ZN( u0_u13_u3_n185 ) );
  NOR2_X1 u0_u13_u3_U31 (.ZN( u0_u13_u3_n135 ) , .A2( u0_u13_u3_n141 ) , .A1( u0_u13_u3_n169 ) );
  OAI222_X1 u0_u13_u3_U32 (.C2( u0_u13_u3_n107 ) , .A2( u0_u13_u3_n108 ) , .B1( u0_u13_u3_n135 ) , .ZN( u0_u13_u3_n138 ) , .B2( u0_u13_u3_n146 ) , .C1( u0_u13_u3_n154 ) , .A1( u0_u13_u3_n164 ) );
  NOR4_X1 u0_u13_u3_U33 (.A4( u0_u13_u3_n157 ) , .A3( u0_u13_u3_n158 ) , .A2( u0_u13_u3_n159 ) , .A1( u0_u13_u3_n160 ) , .ZN( u0_u13_u3_n161 ) );
  AOI21_X1 u0_u13_u3_U34 (.B2( u0_u13_u3_n152 ) , .B1( u0_u13_u3_n153 ) , .ZN( u0_u13_u3_n158 ) , .A( u0_u13_u3_n164 ) );
  AOI21_X1 u0_u13_u3_U35 (.A( u0_u13_u3_n154 ) , .B2( u0_u13_u3_n155 ) , .B1( u0_u13_u3_n156 ) , .ZN( u0_u13_u3_n157 ) );
  AOI21_X1 u0_u13_u3_U36 (.A( u0_u13_u3_n149 ) , .B2( u0_u13_u3_n150 ) , .B1( u0_u13_u3_n151 ) , .ZN( u0_u13_u3_n159 ) );
  AOI211_X1 u0_u13_u3_U37 (.ZN( u0_u13_u3_n109 ) , .A( u0_u13_u3_n119 ) , .C2( u0_u13_u3_n129 ) , .B( u0_u13_u3_n138 ) , .C1( u0_u13_u3_n141 ) );
  AOI211_X1 u0_u13_u3_U38 (.B( u0_u13_u3_n119 ) , .A( u0_u13_u3_n120 ) , .C2( u0_u13_u3_n121 ) , .ZN( u0_u13_u3_n122 ) , .C1( u0_u13_u3_n179 ) );
  INV_X1 u0_u13_u3_U39 (.A( u0_u13_u3_n156 ) , .ZN( u0_u13_u3_n179 ) );
  INV_X1 u0_u13_u3_U4 (.A( u0_u13_u3_n140 ) , .ZN( u0_u13_u3_n182 ) );
  OAI22_X1 u0_u13_u3_U40 (.B1( u0_u13_u3_n118 ) , .ZN( u0_u13_u3_n120 ) , .A1( u0_u13_u3_n135 ) , .B2( u0_u13_u3_n154 ) , .A2( u0_u13_u3_n178 ) );
  AND3_X1 u0_u13_u3_U41 (.ZN( u0_u13_u3_n118 ) , .A2( u0_u13_u3_n124 ) , .A1( u0_u13_u3_n144 ) , .A3( u0_u13_u3_n152 ) );
  INV_X1 u0_u13_u3_U42 (.A( u0_u13_u3_n121 ) , .ZN( u0_u13_u3_n164 ) );
  NAND2_X1 u0_u13_u3_U43 (.ZN( u0_u13_u3_n133 ) , .A1( u0_u13_u3_n154 ) , .A2( u0_u13_u3_n164 ) );
  OAI211_X1 u0_u13_u3_U44 (.B( u0_u13_u3_n127 ) , .ZN( u0_u13_u3_n139 ) , .C1( u0_u13_u3_n150 ) , .C2( u0_u13_u3_n154 ) , .A( u0_u13_u3_n184 ) );
  INV_X1 u0_u13_u3_U45 (.A( u0_u13_u3_n125 ) , .ZN( u0_u13_u3_n184 ) );
  AOI221_X1 u0_u13_u3_U46 (.A( u0_u13_u3_n126 ) , .ZN( u0_u13_u3_n127 ) , .C2( u0_u13_u3_n132 ) , .C1( u0_u13_u3_n169 ) , .B2( u0_u13_u3_n170 ) , .B1( u0_u13_u3_n174 ) );
  OAI22_X1 u0_u13_u3_U47 (.A1( u0_u13_u3_n124 ) , .ZN( u0_u13_u3_n125 ) , .B2( u0_u13_u3_n145 ) , .A2( u0_u13_u3_n165 ) , .B1( u0_u13_u3_n167 ) );
  NOR2_X1 u0_u13_u3_U48 (.A1( u0_u13_u3_n113 ) , .ZN( u0_u13_u3_n131 ) , .A2( u0_u13_u3_n154 ) );
  NAND2_X1 u0_u13_u3_U49 (.A1( u0_u13_u3_n103 ) , .ZN( u0_u13_u3_n150 ) , .A2( u0_u13_u3_n99 ) );
  INV_X1 u0_u13_u3_U5 (.A( u0_u13_u3_n117 ) , .ZN( u0_u13_u3_n178 ) );
  NAND2_X1 u0_u13_u3_U50 (.A2( u0_u13_u3_n102 ) , .ZN( u0_u13_u3_n155 ) , .A1( u0_u13_u3_n97 ) );
  INV_X1 u0_u13_u3_U51 (.A( u0_u13_u3_n141 ) , .ZN( u0_u13_u3_n167 ) );
  AOI21_X1 u0_u13_u3_U52 (.B2( u0_u13_u3_n114 ) , .B1( u0_u13_u3_n146 ) , .A( u0_u13_u3_n154 ) , .ZN( u0_u13_u3_n94 ) );
  AOI21_X1 u0_u13_u3_U53 (.ZN( u0_u13_u3_n110 ) , .B2( u0_u13_u3_n142 ) , .B1( u0_u13_u3_n186 ) , .A( u0_u13_u3_n95 ) );
  INV_X1 u0_u13_u3_U54 (.A( u0_u13_u3_n145 ) , .ZN( u0_u13_u3_n186 ) );
  AOI21_X1 u0_u13_u3_U55 (.B1( u0_u13_u3_n124 ) , .A( u0_u13_u3_n149 ) , .B2( u0_u13_u3_n155 ) , .ZN( u0_u13_u3_n95 ) );
  INV_X1 u0_u13_u3_U56 (.A( u0_u13_u3_n149 ) , .ZN( u0_u13_u3_n169 ) );
  NAND2_X1 u0_u13_u3_U57 (.ZN( u0_u13_u3_n124 ) , .A1( u0_u13_u3_n96 ) , .A2( u0_u13_u3_n97 ) );
  NAND2_X1 u0_u13_u3_U58 (.A2( u0_u13_u3_n100 ) , .ZN( u0_u13_u3_n146 ) , .A1( u0_u13_u3_n96 ) );
  NAND2_X1 u0_u13_u3_U59 (.A1( u0_u13_u3_n101 ) , .ZN( u0_u13_u3_n145 ) , .A2( u0_u13_u3_n99 ) );
  AOI221_X1 u0_u13_u3_U6 (.A( u0_u13_u3_n131 ) , .C2( u0_u13_u3_n132 ) , .C1( u0_u13_u3_n133 ) , .ZN( u0_u13_u3_n134 ) , .B1( u0_u13_u3_n143 ) , .B2( u0_u13_u3_n177 ) );
  NAND2_X1 u0_u13_u3_U60 (.A1( u0_u13_u3_n100 ) , .ZN( u0_u13_u3_n156 ) , .A2( u0_u13_u3_n99 ) );
  NAND2_X1 u0_u13_u3_U61 (.A2( u0_u13_u3_n101 ) , .A1( u0_u13_u3_n104 ) , .ZN( u0_u13_u3_n148 ) );
  NAND2_X1 u0_u13_u3_U62 (.A1( u0_u13_u3_n100 ) , .A2( u0_u13_u3_n102 ) , .ZN( u0_u13_u3_n128 ) );
  NAND2_X1 u0_u13_u3_U63 (.A2( u0_u13_u3_n101 ) , .A1( u0_u13_u3_n102 ) , .ZN( u0_u13_u3_n152 ) );
  NAND2_X1 u0_u13_u3_U64 (.A2( u0_u13_u3_n101 ) , .ZN( u0_u13_u3_n114 ) , .A1( u0_u13_u3_n96 ) );
  NAND2_X1 u0_u13_u3_U65 (.ZN( u0_u13_u3_n107 ) , .A1( u0_u13_u3_n97 ) , .A2( u0_u13_u3_n99 ) );
  NAND2_X1 u0_u13_u3_U66 (.A2( u0_u13_u3_n100 ) , .A1( u0_u13_u3_n104 ) , .ZN( u0_u13_u3_n113 ) );
  NAND2_X1 u0_u13_u3_U67 (.A1( u0_u13_u3_n104 ) , .ZN( u0_u13_u3_n153 ) , .A2( u0_u13_u3_n97 ) );
  NAND2_X1 u0_u13_u3_U68 (.A2( u0_u13_u3_n103 ) , .A1( u0_u13_u3_n104 ) , .ZN( u0_u13_u3_n130 ) );
  NAND2_X1 u0_u13_u3_U69 (.A2( u0_u13_u3_n103 ) , .ZN( u0_u13_u3_n144 ) , .A1( u0_u13_u3_n96 ) );
  OAI22_X1 u0_u13_u3_U7 (.B2( u0_u13_u3_n147 ) , .A2( u0_u13_u3_n148 ) , .ZN( u0_u13_u3_n160 ) , .B1( u0_u13_u3_n165 ) , .A1( u0_u13_u3_n168 ) );
  NAND2_X1 u0_u13_u3_U70 (.A1( u0_u13_u3_n102 ) , .A2( u0_u13_u3_n103 ) , .ZN( u0_u13_u3_n108 ) );
  NOR2_X1 u0_u13_u3_U71 (.A2( u0_u13_X_19 ) , .A1( u0_u13_X_20 ) , .ZN( u0_u13_u3_n99 ) );
  NOR2_X1 u0_u13_u3_U72 (.A2( u0_u13_X_21 ) , .A1( u0_u13_X_24 ) , .ZN( u0_u13_u3_n103 ) );
  NOR2_X1 u0_u13_u3_U73 (.A2( u0_u13_X_24 ) , .A1( u0_u13_u3_n171 ) , .ZN( u0_u13_u3_n97 ) );
  NOR2_X1 u0_u13_u3_U74 (.A2( u0_u13_X_23 ) , .ZN( u0_u13_u3_n141 ) , .A1( u0_u13_u3_n166 ) );
  NOR2_X1 u0_u13_u3_U75 (.A2( u0_u13_X_19 ) , .A1( u0_u13_u3_n172 ) , .ZN( u0_u13_u3_n96 ) );
  NAND2_X1 u0_u13_u3_U76 (.A1( u0_u13_X_22 ) , .A2( u0_u13_X_23 ) , .ZN( u0_u13_u3_n154 ) );
  NAND2_X1 u0_u13_u3_U77 (.A1( u0_u13_X_23 ) , .ZN( u0_u13_u3_n149 ) , .A2( u0_u13_u3_n166 ) );
  NOR2_X1 u0_u13_u3_U78 (.A2( u0_u13_X_22 ) , .A1( u0_u13_X_23 ) , .ZN( u0_u13_u3_n121 ) );
  AND2_X1 u0_u13_u3_U79 (.A1( u0_u13_X_24 ) , .ZN( u0_u13_u3_n101 ) , .A2( u0_u13_u3_n171 ) );
  AND3_X1 u0_u13_u3_U8 (.A3( u0_u13_u3_n144 ) , .A2( u0_u13_u3_n145 ) , .A1( u0_u13_u3_n146 ) , .ZN( u0_u13_u3_n147 ) );
  AND2_X1 u0_u13_u3_U80 (.A1( u0_u13_X_19 ) , .ZN( u0_u13_u3_n102 ) , .A2( u0_u13_u3_n172 ) );
  AND2_X1 u0_u13_u3_U81 (.A1( u0_u13_X_21 ) , .A2( u0_u13_X_24 ) , .ZN( u0_u13_u3_n100 ) );
  AND2_X1 u0_u13_u3_U82 (.A2( u0_u13_X_19 ) , .A1( u0_u13_X_20 ) , .ZN( u0_u13_u3_n104 ) );
  INV_X1 u0_u13_u3_U83 (.A( u0_u13_X_22 ) , .ZN( u0_u13_u3_n166 ) );
  INV_X1 u0_u13_u3_U84 (.A( u0_u13_X_21 ) , .ZN( u0_u13_u3_n171 ) );
  INV_X1 u0_u13_u3_U85 (.A( u0_u13_X_20 ) , .ZN( u0_u13_u3_n172 ) );
  NAND4_X1 u0_u13_u3_U86 (.ZN( u0_out13_26 ) , .A4( u0_u13_u3_n109 ) , .A3( u0_u13_u3_n110 ) , .A2( u0_u13_u3_n111 ) , .A1( u0_u13_u3_n173 ) );
  INV_X1 u0_u13_u3_U87 (.ZN( u0_u13_u3_n173 ) , .A( u0_u13_u3_n94 ) );
  OAI21_X1 u0_u13_u3_U88 (.ZN( u0_u13_u3_n111 ) , .B2( u0_u13_u3_n117 ) , .A( u0_u13_u3_n133 ) , .B1( u0_u13_u3_n176 ) );
  NAND4_X1 u0_u13_u3_U89 (.ZN( u0_out13_20 ) , .A4( u0_u13_u3_n122 ) , .A3( u0_u13_u3_n123 ) , .A1( u0_u13_u3_n175 ) , .A2( u0_u13_u3_n180 ) );
  INV_X1 u0_u13_u3_U9 (.A( u0_u13_u3_n143 ) , .ZN( u0_u13_u3_n168 ) );
  INV_X1 u0_u13_u3_U90 (.A( u0_u13_u3_n112 ) , .ZN( u0_u13_u3_n175 ) );
  INV_X1 u0_u13_u3_U91 (.A( u0_u13_u3_n126 ) , .ZN( u0_u13_u3_n180 ) );
  NAND4_X1 u0_u13_u3_U92 (.ZN( u0_out13_1 ) , .A4( u0_u13_u3_n161 ) , .A3( u0_u13_u3_n162 ) , .A2( u0_u13_u3_n163 ) , .A1( u0_u13_u3_n185 ) );
  NAND2_X1 u0_u13_u3_U93 (.ZN( u0_u13_u3_n163 ) , .A2( u0_u13_u3_n170 ) , .A1( u0_u13_u3_n176 ) );
  AOI22_X1 u0_u13_u3_U94 (.B2( u0_u13_u3_n140 ) , .B1( u0_u13_u3_n141 ) , .A2( u0_u13_u3_n142 ) , .ZN( u0_u13_u3_n162 ) , .A1( u0_u13_u3_n177 ) );
  OR4_X1 u0_u13_u3_U95 (.ZN( u0_out13_10 ) , .A4( u0_u13_u3_n136 ) , .A3( u0_u13_u3_n137 ) , .A1( u0_u13_u3_n138 ) , .A2( u0_u13_u3_n139 ) );
  OAI222_X1 u0_u13_u3_U96 (.C1( u0_u13_u3_n128 ) , .ZN( u0_u13_u3_n137 ) , .B1( u0_u13_u3_n148 ) , .A2( u0_u13_u3_n150 ) , .B2( u0_u13_u3_n154 ) , .C2( u0_u13_u3_n164 ) , .A1( u0_u13_u3_n167 ) );
  OAI221_X1 u0_u13_u3_U97 (.A( u0_u13_u3_n134 ) , .B2( u0_u13_u3_n135 ) , .ZN( u0_u13_u3_n136 ) , .C1( u0_u13_u3_n149 ) , .B1( u0_u13_u3_n151 ) , .C2( u0_u13_u3_n183 ) );
  NAND3_X1 u0_u13_u3_U98 (.A1( u0_u13_u3_n114 ) , .ZN( u0_u13_u3_n115 ) , .A2( u0_u13_u3_n145 ) , .A3( u0_u13_u3_n153 ) );
  NAND3_X1 u0_u13_u3_U99 (.ZN( u0_u13_u3_n129 ) , .A2( u0_u13_u3_n144 ) , .A1( u0_u13_u3_n153 ) , .A3( u0_u13_u3_n182 ) );
  AOI21_X1 u0_u13_u4_U10 (.ZN( u0_u13_u4_n106 ) , .B2( u0_u13_u4_n146 ) , .B1( u0_u13_u4_n158 ) , .A( u0_u13_u4_n170 ) );
  AOI21_X1 u0_u13_u4_U11 (.ZN( u0_u13_u4_n108 ) , .B2( u0_u13_u4_n134 ) , .B1( u0_u13_u4_n155 ) , .A( u0_u13_u4_n156 ) );
  AOI21_X1 u0_u13_u4_U12 (.ZN( u0_u13_u4_n109 ) , .A( u0_u13_u4_n153 ) , .B1( u0_u13_u4_n159 ) , .B2( u0_u13_u4_n184 ) );
  AOI211_X1 u0_u13_u4_U13 (.B( u0_u13_u4_n136 ) , .A( u0_u13_u4_n137 ) , .C2( u0_u13_u4_n138 ) , .ZN( u0_u13_u4_n139 ) , .C1( u0_u13_u4_n182 ) );
  OAI22_X1 u0_u13_u4_U14 (.B2( u0_u13_u4_n135 ) , .ZN( u0_u13_u4_n137 ) , .B1( u0_u13_u4_n153 ) , .A1( u0_u13_u4_n155 ) , .A2( u0_u13_u4_n171 ) );
  AND3_X1 u0_u13_u4_U15 (.A2( u0_u13_u4_n134 ) , .ZN( u0_u13_u4_n135 ) , .A3( u0_u13_u4_n145 ) , .A1( u0_u13_u4_n157 ) );
  NAND2_X1 u0_u13_u4_U16 (.ZN( u0_u13_u4_n132 ) , .A2( u0_u13_u4_n170 ) , .A1( u0_u13_u4_n173 ) );
  AOI21_X1 u0_u13_u4_U17 (.B2( u0_u13_u4_n160 ) , .B1( u0_u13_u4_n161 ) , .ZN( u0_u13_u4_n162 ) , .A( u0_u13_u4_n170 ) );
  AOI21_X1 u0_u13_u4_U18 (.ZN( u0_u13_u4_n107 ) , .B2( u0_u13_u4_n143 ) , .A( u0_u13_u4_n174 ) , .B1( u0_u13_u4_n184 ) );
  AOI21_X1 u0_u13_u4_U19 (.B2( u0_u13_u4_n158 ) , .B1( u0_u13_u4_n159 ) , .ZN( u0_u13_u4_n163 ) , .A( u0_u13_u4_n174 ) );
  AOI21_X1 u0_u13_u4_U20 (.A( u0_u13_u4_n153 ) , .B2( u0_u13_u4_n154 ) , .B1( u0_u13_u4_n155 ) , .ZN( u0_u13_u4_n165 ) );
  AOI21_X1 u0_u13_u4_U21 (.A( u0_u13_u4_n156 ) , .B2( u0_u13_u4_n157 ) , .ZN( u0_u13_u4_n164 ) , .B1( u0_u13_u4_n184 ) );
  INV_X1 u0_u13_u4_U22 (.A( u0_u13_u4_n138 ) , .ZN( u0_u13_u4_n170 ) );
  AND2_X1 u0_u13_u4_U23 (.A2( u0_u13_u4_n120 ) , .ZN( u0_u13_u4_n155 ) , .A1( u0_u13_u4_n160 ) );
  INV_X1 u0_u13_u4_U24 (.A( u0_u13_u4_n156 ) , .ZN( u0_u13_u4_n175 ) );
  NAND2_X1 u0_u13_u4_U25 (.A2( u0_u13_u4_n118 ) , .ZN( u0_u13_u4_n131 ) , .A1( u0_u13_u4_n147 ) );
  NAND2_X1 u0_u13_u4_U26 (.A1( u0_u13_u4_n119 ) , .A2( u0_u13_u4_n120 ) , .ZN( u0_u13_u4_n130 ) );
  NAND2_X1 u0_u13_u4_U27 (.ZN( u0_u13_u4_n117 ) , .A2( u0_u13_u4_n118 ) , .A1( u0_u13_u4_n148 ) );
  NAND2_X1 u0_u13_u4_U28 (.ZN( u0_u13_u4_n129 ) , .A1( u0_u13_u4_n134 ) , .A2( u0_u13_u4_n148 ) );
  AND3_X1 u0_u13_u4_U29 (.A1( u0_u13_u4_n119 ) , .A2( u0_u13_u4_n143 ) , .A3( u0_u13_u4_n154 ) , .ZN( u0_u13_u4_n161 ) );
  NOR2_X1 u0_u13_u4_U3 (.ZN( u0_u13_u4_n121 ) , .A1( u0_u13_u4_n181 ) , .A2( u0_u13_u4_n182 ) );
  AND2_X1 u0_u13_u4_U30 (.A1( u0_u13_u4_n145 ) , .A2( u0_u13_u4_n147 ) , .ZN( u0_u13_u4_n159 ) );
  OR3_X1 u0_u13_u4_U31 (.A3( u0_u13_u4_n114 ) , .A2( u0_u13_u4_n115 ) , .A1( u0_u13_u4_n116 ) , .ZN( u0_u13_u4_n136 ) );
  AOI21_X1 u0_u13_u4_U32 (.A( u0_u13_u4_n113 ) , .ZN( u0_u13_u4_n116 ) , .B2( u0_u13_u4_n173 ) , .B1( u0_u13_u4_n174 ) );
  AOI21_X1 u0_u13_u4_U33 (.ZN( u0_u13_u4_n115 ) , .B2( u0_u13_u4_n145 ) , .B1( u0_u13_u4_n146 ) , .A( u0_u13_u4_n156 ) );
  OAI22_X1 u0_u13_u4_U34 (.ZN( u0_u13_u4_n114 ) , .A2( u0_u13_u4_n121 ) , .B1( u0_u13_u4_n160 ) , .B2( u0_u13_u4_n170 ) , .A1( u0_u13_u4_n171 ) );
  INV_X1 u0_u13_u4_U35 (.A( u0_u13_u4_n158 ) , .ZN( u0_u13_u4_n182 ) );
  INV_X1 u0_u13_u4_U36 (.ZN( u0_u13_u4_n181 ) , .A( u0_u13_u4_n96 ) );
  INV_X1 u0_u13_u4_U37 (.A( u0_u13_u4_n144 ) , .ZN( u0_u13_u4_n179 ) );
  INV_X1 u0_u13_u4_U38 (.A( u0_u13_u4_n157 ) , .ZN( u0_u13_u4_n178 ) );
  NAND2_X1 u0_u13_u4_U39 (.A2( u0_u13_u4_n154 ) , .A1( u0_u13_u4_n96 ) , .ZN( u0_u13_u4_n97 ) );
  INV_X1 u0_u13_u4_U4 (.A( u0_u13_u4_n117 ) , .ZN( u0_u13_u4_n184 ) );
  INV_X1 u0_u13_u4_U40 (.A( u0_u13_u4_n143 ) , .ZN( u0_u13_u4_n183 ) );
  NOR2_X1 u0_u13_u4_U41 (.ZN( u0_u13_u4_n138 ) , .A1( u0_u13_u4_n168 ) , .A2( u0_u13_u4_n169 ) );
  NOR2_X1 u0_u13_u4_U42 (.A1( u0_u13_u4_n150 ) , .A2( u0_u13_u4_n152 ) , .ZN( u0_u13_u4_n153 ) );
  NOR2_X1 u0_u13_u4_U43 (.A2( u0_u13_u4_n128 ) , .A1( u0_u13_u4_n138 ) , .ZN( u0_u13_u4_n156 ) );
  AOI22_X1 u0_u13_u4_U44 (.B2( u0_u13_u4_n122 ) , .A1( u0_u13_u4_n123 ) , .ZN( u0_u13_u4_n124 ) , .B1( u0_u13_u4_n128 ) , .A2( u0_u13_u4_n172 ) );
  NAND2_X1 u0_u13_u4_U45 (.A2( u0_u13_u4_n120 ) , .ZN( u0_u13_u4_n123 ) , .A1( u0_u13_u4_n161 ) );
  INV_X1 u0_u13_u4_U46 (.A( u0_u13_u4_n153 ) , .ZN( u0_u13_u4_n172 ) );
  AOI22_X1 u0_u13_u4_U47 (.B2( u0_u13_u4_n132 ) , .A2( u0_u13_u4_n133 ) , .ZN( u0_u13_u4_n140 ) , .A1( u0_u13_u4_n150 ) , .B1( u0_u13_u4_n179 ) );
  NAND2_X1 u0_u13_u4_U48 (.ZN( u0_u13_u4_n133 ) , .A2( u0_u13_u4_n146 ) , .A1( u0_u13_u4_n154 ) );
  NAND2_X1 u0_u13_u4_U49 (.A1( u0_u13_u4_n103 ) , .ZN( u0_u13_u4_n154 ) , .A2( u0_u13_u4_n98 ) );
  INV_X1 u0_u13_u4_U5 (.ZN( u0_u13_u4_n186 ) , .A( u0_u13_u4_n95 ) );
  NAND2_X1 u0_u13_u4_U50 (.A1( u0_u13_u4_n101 ) , .ZN( u0_u13_u4_n158 ) , .A2( u0_u13_u4_n99 ) );
  AOI21_X1 u0_u13_u4_U51 (.ZN( u0_u13_u4_n127 ) , .A( u0_u13_u4_n136 ) , .B2( u0_u13_u4_n150 ) , .B1( u0_u13_u4_n180 ) );
  INV_X1 u0_u13_u4_U52 (.A( u0_u13_u4_n160 ) , .ZN( u0_u13_u4_n180 ) );
  NAND2_X1 u0_u13_u4_U53 (.A2( u0_u13_u4_n104 ) , .A1( u0_u13_u4_n105 ) , .ZN( u0_u13_u4_n146 ) );
  NAND2_X1 u0_u13_u4_U54 (.A2( u0_u13_u4_n101 ) , .A1( u0_u13_u4_n102 ) , .ZN( u0_u13_u4_n160 ) );
  NAND2_X1 u0_u13_u4_U55 (.ZN( u0_u13_u4_n134 ) , .A1( u0_u13_u4_n98 ) , .A2( u0_u13_u4_n99 ) );
  NAND2_X1 u0_u13_u4_U56 (.A1( u0_u13_u4_n103 ) , .A2( u0_u13_u4_n104 ) , .ZN( u0_u13_u4_n143 ) );
  NAND2_X1 u0_u13_u4_U57 (.A2( u0_u13_u4_n105 ) , .ZN( u0_u13_u4_n145 ) , .A1( u0_u13_u4_n98 ) );
  NAND2_X1 u0_u13_u4_U58 (.A1( u0_u13_u4_n100 ) , .A2( u0_u13_u4_n105 ) , .ZN( u0_u13_u4_n120 ) );
  NAND2_X1 u0_u13_u4_U59 (.A1( u0_u13_u4_n102 ) , .A2( u0_u13_u4_n104 ) , .ZN( u0_u13_u4_n148 ) );
  OAI221_X1 u0_u13_u4_U6 (.C1( u0_u13_u4_n134 ) , .B1( u0_u13_u4_n158 ) , .B2( u0_u13_u4_n171 ) , .C2( u0_u13_u4_n173 ) , .A( u0_u13_u4_n94 ) , .ZN( u0_u13_u4_n95 ) );
  NAND2_X1 u0_u13_u4_U60 (.A2( u0_u13_u4_n100 ) , .A1( u0_u13_u4_n103 ) , .ZN( u0_u13_u4_n157 ) );
  INV_X1 u0_u13_u4_U61 (.A( u0_u13_u4_n150 ) , .ZN( u0_u13_u4_n173 ) );
  INV_X1 u0_u13_u4_U62 (.A( u0_u13_u4_n152 ) , .ZN( u0_u13_u4_n171 ) );
  NAND2_X1 u0_u13_u4_U63 (.A1( u0_u13_u4_n100 ) , .ZN( u0_u13_u4_n118 ) , .A2( u0_u13_u4_n99 ) );
  NAND2_X1 u0_u13_u4_U64 (.A2( u0_u13_u4_n100 ) , .A1( u0_u13_u4_n102 ) , .ZN( u0_u13_u4_n144 ) );
  NAND2_X1 u0_u13_u4_U65 (.A2( u0_u13_u4_n101 ) , .A1( u0_u13_u4_n105 ) , .ZN( u0_u13_u4_n96 ) );
  INV_X1 u0_u13_u4_U66 (.A( u0_u13_u4_n128 ) , .ZN( u0_u13_u4_n174 ) );
  NAND2_X1 u0_u13_u4_U67 (.A2( u0_u13_u4_n102 ) , .ZN( u0_u13_u4_n119 ) , .A1( u0_u13_u4_n98 ) );
  NAND2_X1 u0_u13_u4_U68 (.A2( u0_u13_u4_n101 ) , .A1( u0_u13_u4_n103 ) , .ZN( u0_u13_u4_n147 ) );
  NAND2_X1 u0_u13_u4_U69 (.A2( u0_u13_u4_n104 ) , .ZN( u0_u13_u4_n113 ) , .A1( u0_u13_u4_n99 ) );
  AOI222_X1 u0_u13_u4_U7 (.B2( u0_u13_u4_n132 ) , .A1( u0_u13_u4_n138 ) , .C2( u0_u13_u4_n175 ) , .A2( u0_u13_u4_n179 ) , .C1( u0_u13_u4_n181 ) , .B1( u0_u13_u4_n185 ) , .ZN( u0_u13_u4_n94 ) );
  NOR2_X1 u0_u13_u4_U70 (.A2( u0_u13_X_28 ) , .ZN( u0_u13_u4_n150 ) , .A1( u0_u13_u4_n168 ) );
  NOR2_X1 u0_u13_u4_U71 (.A2( u0_u13_X_29 ) , .ZN( u0_u13_u4_n152 ) , .A1( u0_u13_u4_n169 ) );
  NOR2_X1 u0_u13_u4_U72 (.A2( u0_u13_X_30 ) , .ZN( u0_u13_u4_n105 ) , .A1( u0_u13_u4_n176 ) );
  NOR2_X1 u0_u13_u4_U73 (.A2( u0_u13_X_26 ) , .ZN( u0_u13_u4_n100 ) , .A1( u0_u13_u4_n177 ) );
  NOR2_X1 u0_u13_u4_U74 (.A2( u0_u13_X_28 ) , .A1( u0_u13_X_29 ) , .ZN( u0_u13_u4_n128 ) );
  NOR2_X1 u0_u13_u4_U75 (.A2( u0_u13_X_27 ) , .A1( u0_u13_X_30 ) , .ZN( u0_u13_u4_n102 ) );
  NOR2_X1 u0_u13_u4_U76 (.A2( u0_u13_X_25 ) , .A1( u0_u13_X_26 ) , .ZN( u0_u13_u4_n98 ) );
  AND2_X1 u0_u13_u4_U77 (.A2( u0_u13_X_25 ) , .A1( u0_u13_X_26 ) , .ZN( u0_u13_u4_n104 ) );
  AND2_X1 u0_u13_u4_U78 (.A1( u0_u13_X_30 ) , .A2( u0_u13_u4_n176 ) , .ZN( u0_u13_u4_n99 ) );
  AND2_X1 u0_u13_u4_U79 (.A1( u0_u13_X_26 ) , .ZN( u0_u13_u4_n101 ) , .A2( u0_u13_u4_n177 ) );
  INV_X1 u0_u13_u4_U8 (.A( u0_u13_u4_n113 ) , .ZN( u0_u13_u4_n185 ) );
  AND2_X1 u0_u13_u4_U80 (.A1( u0_u13_X_27 ) , .A2( u0_u13_X_30 ) , .ZN( u0_u13_u4_n103 ) );
  INV_X1 u0_u13_u4_U81 (.A( u0_u13_X_28 ) , .ZN( u0_u13_u4_n169 ) );
  INV_X1 u0_u13_u4_U82 (.A( u0_u13_X_29 ) , .ZN( u0_u13_u4_n168 ) );
  INV_X1 u0_u13_u4_U83 (.A( u0_u13_X_25 ) , .ZN( u0_u13_u4_n177 ) );
  INV_X1 u0_u13_u4_U84 (.A( u0_u13_X_27 ) , .ZN( u0_u13_u4_n176 ) );
  NAND4_X1 u0_u13_u4_U85 (.ZN( u0_out13_25 ) , .A4( u0_u13_u4_n139 ) , .A3( u0_u13_u4_n140 ) , .A2( u0_u13_u4_n141 ) , .A1( u0_u13_u4_n142 ) );
  OAI21_X1 u0_u13_u4_U86 (.A( u0_u13_u4_n128 ) , .B2( u0_u13_u4_n129 ) , .B1( u0_u13_u4_n130 ) , .ZN( u0_u13_u4_n142 ) );
  OAI21_X1 u0_u13_u4_U87 (.B2( u0_u13_u4_n131 ) , .ZN( u0_u13_u4_n141 ) , .A( u0_u13_u4_n175 ) , .B1( u0_u13_u4_n183 ) );
  NAND4_X1 u0_u13_u4_U88 (.ZN( u0_out13_14 ) , .A4( u0_u13_u4_n124 ) , .A3( u0_u13_u4_n125 ) , .A2( u0_u13_u4_n126 ) , .A1( u0_u13_u4_n127 ) );
  AOI22_X1 u0_u13_u4_U89 (.B2( u0_u13_u4_n117 ) , .ZN( u0_u13_u4_n126 ) , .A1( u0_u13_u4_n129 ) , .B1( u0_u13_u4_n152 ) , .A2( u0_u13_u4_n175 ) );
  NOR4_X1 u0_u13_u4_U9 (.A4( u0_u13_u4_n106 ) , .A3( u0_u13_u4_n107 ) , .A2( u0_u13_u4_n108 ) , .A1( u0_u13_u4_n109 ) , .ZN( u0_u13_u4_n110 ) );
  AOI22_X1 u0_u13_u4_U90 (.ZN( u0_u13_u4_n125 ) , .B2( u0_u13_u4_n131 ) , .A2( u0_u13_u4_n132 ) , .B1( u0_u13_u4_n138 ) , .A1( u0_u13_u4_n178 ) );
  NAND4_X1 u0_u13_u4_U91 (.ZN( u0_out13_8 ) , .A4( u0_u13_u4_n110 ) , .A3( u0_u13_u4_n111 ) , .A2( u0_u13_u4_n112 ) , .A1( u0_u13_u4_n186 ) );
  NAND2_X1 u0_u13_u4_U92 (.ZN( u0_u13_u4_n112 ) , .A2( u0_u13_u4_n130 ) , .A1( u0_u13_u4_n150 ) );
  AOI22_X1 u0_u13_u4_U93 (.ZN( u0_u13_u4_n111 ) , .B2( u0_u13_u4_n132 ) , .A1( u0_u13_u4_n152 ) , .B1( u0_u13_u4_n178 ) , .A2( u0_u13_u4_n97 ) );
  AOI22_X1 u0_u13_u4_U94 (.B2( u0_u13_u4_n149 ) , .B1( u0_u13_u4_n150 ) , .A2( u0_u13_u4_n151 ) , .A1( u0_u13_u4_n152 ) , .ZN( u0_u13_u4_n167 ) );
  NOR4_X1 u0_u13_u4_U95 (.A4( u0_u13_u4_n162 ) , .A3( u0_u13_u4_n163 ) , .A2( u0_u13_u4_n164 ) , .A1( u0_u13_u4_n165 ) , .ZN( u0_u13_u4_n166 ) );
  NAND3_X1 u0_u13_u4_U96 (.ZN( u0_out13_3 ) , .A3( u0_u13_u4_n166 ) , .A1( u0_u13_u4_n167 ) , .A2( u0_u13_u4_n186 ) );
  NAND3_X1 u0_u13_u4_U97 (.A3( u0_u13_u4_n146 ) , .A2( u0_u13_u4_n147 ) , .A1( u0_u13_u4_n148 ) , .ZN( u0_u13_u4_n149 ) );
  NAND3_X1 u0_u13_u4_U98 (.A3( u0_u13_u4_n143 ) , .A2( u0_u13_u4_n144 ) , .A1( u0_u13_u4_n145 ) , .ZN( u0_u13_u4_n151 ) );
  NAND3_X1 u0_u13_u4_U99 (.A3( u0_u13_u4_n121 ) , .ZN( u0_u13_u4_n122 ) , .A2( u0_u13_u4_n144 ) , .A1( u0_u13_u4_n154 ) );
  INV_X1 u0_u13_u5_U10 (.A( u0_u13_u5_n121 ) , .ZN( u0_u13_u5_n177 ) );
  NOR3_X1 u0_u13_u5_U100 (.A3( u0_u13_u5_n141 ) , .A1( u0_u13_u5_n142 ) , .ZN( u0_u13_u5_n143 ) , .A2( u0_u13_u5_n191 ) );
  NAND4_X1 u0_u13_u5_U101 (.ZN( u0_out13_4 ) , .A4( u0_u13_u5_n112 ) , .A2( u0_u13_u5_n113 ) , .A1( u0_u13_u5_n114 ) , .A3( u0_u13_u5_n195 ) );
  AOI211_X1 u0_u13_u5_U102 (.A( u0_u13_u5_n110 ) , .C1( u0_u13_u5_n111 ) , .ZN( u0_u13_u5_n112 ) , .B( u0_u13_u5_n118 ) , .C2( u0_u13_u5_n177 ) );
  AOI222_X1 u0_u13_u5_U103 (.ZN( u0_u13_u5_n113 ) , .A1( u0_u13_u5_n131 ) , .C1( u0_u13_u5_n148 ) , .B2( u0_u13_u5_n174 ) , .C2( u0_u13_u5_n178 ) , .A2( u0_u13_u5_n179 ) , .B1( u0_u13_u5_n99 ) );
  NAND3_X1 u0_u13_u5_U104 (.A2( u0_u13_u5_n154 ) , .A3( u0_u13_u5_n158 ) , .A1( u0_u13_u5_n161 ) , .ZN( u0_u13_u5_n99 ) );
  NOR2_X1 u0_u13_u5_U11 (.ZN( u0_u13_u5_n160 ) , .A2( u0_u13_u5_n173 ) , .A1( u0_u13_u5_n177 ) );
  INV_X1 u0_u13_u5_U12 (.A( u0_u13_u5_n150 ) , .ZN( u0_u13_u5_n174 ) );
  AOI21_X1 u0_u13_u5_U13 (.A( u0_u13_u5_n160 ) , .B2( u0_u13_u5_n161 ) , .ZN( u0_u13_u5_n162 ) , .B1( u0_u13_u5_n192 ) );
  INV_X1 u0_u13_u5_U14 (.A( u0_u13_u5_n159 ) , .ZN( u0_u13_u5_n192 ) );
  AOI21_X1 u0_u13_u5_U15 (.A( u0_u13_u5_n156 ) , .B2( u0_u13_u5_n157 ) , .B1( u0_u13_u5_n158 ) , .ZN( u0_u13_u5_n163 ) );
  AOI21_X1 u0_u13_u5_U16 (.B2( u0_u13_u5_n139 ) , .B1( u0_u13_u5_n140 ) , .ZN( u0_u13_u5_n141 ) , .A( u0_u13_u5_n150 ) );
  OAI21_X1 u0_u13_u5_U17 (.A( u0_u13_u5_n133 ) , .B2( u0_u13_u5_n134 ) , .B1( u0_u13_u5_n135 ) , .ZN( u0_u13_u5_n142 ) );
  OAI21_X1 u0_u13_u5_U18 (.ZN( u0_u13_u5_n133 ) , .B2( u0_u13_u5_n147 ) , .A( u0_u13_u5_n173 ) , .B1( u0_u13_u5_n188 ) );
  NAND2_X1 u0_u13_u5_U19 (.A2( u0_u13_u5_n119 ) , .A1( u0_u13_u5_n123 ) , .ZN( u0_u13_u5_n137 ) );
  INV_X1 u0_u13_u5_U20 (.A( u0_u13_u5_n155 ) , .ZN( u0_u13_u5_n194 ) );
  NAND2_X1 u0_u13_u5_U21 (.A1( u0_u13_u5_n121 ) , .ZN( u0_u13_u5_n132 ) , .A2( u0_u13_u5_n172 ) );
  NAND2_X1 u0_u13_u5_U22 (.A2( u0_u13_u5_n122 ) , .ZN( u0_u13_u5_n136 ) , .A1( u0_u13_u5_n154 ) );
  NAND2_X1 u0_u13_u5_U23 (.A2( u0_u13_u5_n119 ) , .A1( u0_u13_u5_n120 ) , .ZN( u0_u13_u5_n159 ) );
  INV_X1 u0_u13_u5_U24 (.A( u0_u13_u5_n156 ) , .ZN( u0_u13_u5_n175 ) );
  INV_X1 u0_u13_u5_U25 (.A( u0_u13_u5_n158 ) , .ZN( u0_u13_u5_n188 ) );
  INV_X1 u0_u13_u5_U26 (.A( u0_u13_u5_n152 ) , .ZN( u0_u13_u5_n179 ) );
  INV_X1 u0_u13_u5_U27 (.A( u0_u13_u5_n140 ) , .ZN( u0_u13_u5_n182 ) );
  INV_X1 u0_u13_u5_U28 (.A( u0_u13_u5_n151 ) , .ZN( u0_u13_u5_n183 ) );
  INV_X1 u0_u13_u5_U29 (.A( u0_u13_u5_n123 ) , .ZN( u0_u13_u5_n185 ) );
  NOR2_X1 u0_u13_u5_U3 (.ZN( u0_u13_u5_n134 ) , .A1( u0_u13_u5_n183 ) , .A2( u0_u13_u5_n190 ) );
  INV_X1 u0_u13_u5_U30 (.A( u0_u13_u5_n161 ) , .ZN( u0_u13_u5_n184 ) );
  INV_X1 u0_u13_u5_U31 (.A( u0_u13_u5_n139 ) , .ZN( u0_u13_u5_n189 ) );
  INV_X1 u0_u13_u5_U32 (.A( u0_u13_u5_n157 ) , .ZN( u0_u13_u5_n190 ) );
  INV_X1 u0_u13_u5_U33 (.A( u0_u13_u5_n120 ) , .ZN( u0_u13_u5_n193 ) );
  NAND2_X1 u0_u13_u5_U34 (.ZN( u0_u13_u5_n111 ) , .A1( u0_u13_u5_n140 ) , .A2( u0_u13_u5_n155 ) );
  INV_X1 u0_u13_u5_U35 (.A( u0_u13_u5_n117 ) , .ZN( u0_u13_u5_n196 ) );
  OAI221_X1 u0_u13_u5_U36 (.A( u0_u13_u5_n116 ) , .ZN( u0_u13_u5_n117 ) , .B2( u0_u13_u5_n119 ) , .C1( u0_u13_u5_n153 ) , .C2( u0_u13_u5_n158 ) , .B1( u0_u13_u5_n172 ) );
  AOI222_X1 u0_u13_u5_U37 (.ZN( u0_u13_u5_n116 ) , .B2( u0_u13_u5_n145 ) , .C1( u0_u13_u5_n148 ) , .A2( u0_u13_u5_n174 ) , .C2( u0_u13_u5_n177 ) , .B1( u0_u13_u5_n187 ) , .A1( u0_u13_u5_n193 ) );
  INV_X1 u0_u13_u5_U38 (.A( u0_u13_u5_n115 ) , .ZN( u0_u13_u5_n187 ) );
  NOR2_X1 u0_u13_u5_U39 (.ZN( u0_u13_u5_n100 ) , .A1( u0_u13_u5_n170 ) , .A2( u0_u13_u5_n180 ) );
  INV_X1 u0_u13_u5_U4 (.A( u0_u13_u5_n138 ) , .ZN( u0_u13_u5_n191 ) );
  AOI22_X1 u0_u13_u5_U40 (.B2( u0_u13_u5_n131 ) , .A2( u0_u13_u5_n146 ) , .ZN( u0_u13_u5_n169 ) , .B1( u0_u13_u5_n174 ) , .A1( u0_u13_u5_n185 ) );
  NOR2_X1 u0_u13_u5_U41 (.A1( u0_u13_u5_n146 ) , .ZN( u0_u13_u5_n150 ) , .A2( u0_u13_u5_n173 ) );
  AOI21_X1 u0_u13_u5_U42 (.A( u0_u13_u5_n118 ) , .B2( u0_u13_u5_n145 ) , .ZN( u0_u13_u5_n168 ) , .B1( u0_u13_u5_n186 ) );
  INV_X1 u0_u13_u5_U43 (.A( u0_u13_u5_n122 ) , .ZN( u0_u13_u5_n186 ) );
  NOR2_X1 u0_u13_u5_U44 (.A1( u0_u13_u5_n146 ) , .ZN( u0_u13_u5_n152 ) , .A2( u0_u13_u5_n176 ) );
  NOR2_X1 u0_u13_u5_U45 (.A1( u0_u13_u5_n115 ) , .ZN( u0_u13_u5_n118 ) , .A2( u0_u13_u5_n153 ) );
  NOR2_X1 u0_u13_u5_U46 (.A2( u0_u13_u5_n145 ) , .ZN( u0_u13_u5_n156 ) , .A1( u0_u13_u5_n174 ) );
  NOR2_X1 u0_u13_u5_U47 (.ZN( u0_u13_u5_n121 ) , .A2( u0_u13_u5_n145 ) , .A1( u0_u13_u5_n176 ) );
  AOI22_X1 u0_u13_u5_U48 (.ZN( u0_u13_u5_n114 ) , .A2( u0_u13_u5_n137 ) , .A1( u0_u13_u5_n145 ) , .B2( u0_u13_u5_n175 ) , .B1( u0_u13_u5_n193 ) );
  OAI211_X1 u0_u13_u5_U49 (.B( u0_u13_u5_n124 ) , .A( u0_u13_u5_n125 ) , .C2( u0_u13_u5_n126 ) , .C1( u0_u13_u5_n127 ) , .ZN( u0_u13_u5_n128 ) );
  OAI21_X1 u0_u13_u5_U5 (.B2( u0_u13_u5_n136 ) , .B1( u0_u13_u5_n137 ) , .ZN( u0_u13_u5_n138 ) , .A( u0_u13_u5_n177 ) );
  NOR3_X1 u0_u13_u5_U50 (.ZN( u0_u13_u5_n127 ) , .A1( u0_u13_u5_n136 ) , .A3( u0_u13_u5_n148 ) , .A2( u0_u13_u5_n182 ) );
  OAI21_X1 u0_u13_u5_U51 (.ZN( u0_u13_u5_n124 ) , .A( u0_u13_u5_n177 ) , .B2( u0_u13_u5_n183 ) , .B1( u0_u13_u5_n189 ) );
  OAI21_X1 u0_u13_u5_U52 (.ZN( u0_u13_u5_n125 ) , .A( u0_u13_u5_n174 ) , .B2( u0_u13_u5_n185 ) , .B1( u0_u13_u5_n190 ) );
  AOI21_X1 u0_u13_u5_U53 (.A( u0_u13_u5_n153 ) , .B2( u0_u13_u5_n154 ) , .B1( u0_u13_u5_n155 ) , .ZN( u0_u13_u5_n164 ) );
  AOI21_X1 u0_u13_u5_U54 (.ZN( u0_u13_u5_n110 ) , .B1( u0_u13_u5_n122 ) , .B2( u0_u13_u5_n139 ) , .A( u0_u13_u5_n153 ) );
  INV_X1 u0_u13_u5_U55 (.A( u0_u13_u5_n153 ) , .ZN( u0_u13_u5_n176 ) );
  INV_X1 u0_u13_u5_U56 (.A( u0_u13_u5_n126 ) , .ZN( u0_u13_u5_n173 ) );
  AND2_X1 u0_u13_u5_U57 (.A2( u0_u13_u5_n104 ) , .A1( u0_u13_u5_n107 ) , .ZN( u0_u13_u5_n147 ) );
  AND2_X1 u0_u13_u5_U58 (.A2( u0_u13_u5_n104 ) , .A1( u0_u13_u5_n108 ) , .ZN( u0_u13_u5_n148 ) );
  NAND2_X1 u0_u13_u5_U59 (.A1( u0_u13_u5_n105 ) , .A2( u0_u13_u5_n106 ) , .ZN( u0_u13_u5_n158 ) );
  INV_X1 u0_u13_u5_U6 (.A( u0_u13_u5_n135 ) , .ZN( u0_u13_u5_n178 ) );
  NAND2_X1 u0_u13_u5_U60 (.A2( u0_u13_u5_n108 ) , .A1( u0_u13_u5_n109 ) , .ZN( u0_u13_u5_n139 ) );
  NAND2_X1 u0_u13_u5_U61 (.A1( u0_u13_u5_n106 ) , .A2( u0_u13_u5_n108 ) , .ZN( u0_u13_u5_n119 ) );
  NAND2_X1 u0_u13_u5_U62 (.A2( u0_u13_u5_n103 ) , .A1( u0_u13_u5_n105 ) , .ZN( u0_u13_u5_n140 ) );
  NAND2_X1 u0_u13_u5_U63 (.A2( u0_u13_u5_n104 ) , .A1( u0_u13_u5_n105 ) , .ZN( u0_u13_u5_n155 ) );
  NAND2_X1 u0_u13_u5_U64 (.A2( u0_u13_u5_n106 ) , .A1( u0_u13_u5_n107 ) , .ZN( u0_u13_u5_n122 ) );
  NAND2_X1 u0_u13_u5_U65 (.A2( u0_u13_u5_n100 ) , .A1( u0_u13_u5_n106 ) , .ZN( u0_u13_u5_n115 ) );
  NAND2_X1 u0_u13_u5_U66 (.A2( u0_u13_u5_n100 ) , .A1( u0_u13_u5_n103 ) , .ZN( u0_u13_u5_n161 ) );
  NAND2_X1 u0_u13_u5_U67 (.A1( u0_u13_u5_n105 ) , .A2( u0_u13_u5_n109 ) , .ZN( u0_u13_u5_n154 ) );
  INV_X1 u0_u13_u5_U68 (.A( u0_u13_u5_n146 ) , .ZN( u0_u13_u5_n172 ) );
  NAND2_X1 u0_u13_u5_U69 (.A1( u0_u13_u5_n103 ) , .A2( u0_u13_u5_n108 ) , .ZN( u0_u13_u5_n123 ) );
  OAI22_X1 u0_u13_u5_U7 (.B2( u0_u13_u5_n149 ) , .B1( u0_u13_u5_n150 ) , .A2( u0_u13_u5_n151 ) , .A1( u0_u13_u5_n152 ) , .ZN( u0_u13_u5_n165 ) );
  NAND2_X1 u0_u13_u5_U70 (.A2( u0_u13_u5_n103 ) , .A1( u0_u13_u5_n107 ) , .ZN( u0_u13_u5_n151 ) );
  NAND2_X1 u0_u13_u5_U71 (.A2( u0_u13_u5_n107 ) , .A1( u0_u13_u5_n109 ) , .ZN( u0_u13_u5_n120 ) );
  NAND2_X1 u0_u13_u5_U72 (.A2( u0_u13_u5_n100 ) , .A1( u0_u13_u5_n109 ) , .ZN( u0_u13_u5_n157 ) );
  AND2_X1 u0_u13_u5_U73 (.A2( u0_u13_u5_n100 ) , .A1( u0_u13_u5_n104 ) , .ZN( u0_u13_u5_n131 ) );
  INV_X1 u0_u13_u5_U74 (.A( u0_u13_u5_n102 ) , .ZN( u0_u13_u5_n195 ) );
  OAI221_X1 u0_u13_u5_U75 (.A( u0_u13_u5_n101 ) , .ZN( u0_u13_u5_n102 ) , .C2( u0_u13_u5_n115 ) , .C1( u0_u13_u5_n126 ) , .B1( u0_u13_u5_n134 ) , .B2( u0_u13_u5_n160 ) );
  OAI21_X1 u0_u13_u5_U76 (.ZN( u0_u13_u5_n101 ) , .B1( u0_u13_u5_n137 ) , .A( u0_u13_u5_n146 ) , .B2( u0_u13_u5_n147 ) );
  NOR2_X1 u0_u13_u5_U77 (.A2( u0_u13_X_34 ) , .A1( u0_u13_X_35 ) , .ZN( u0_u13_u5_n145 ) );
  NOR2_X1 u0_u13_u5_U78 (.A2( u0_u13_X_34 ) , .ZN( u0_u13_u5_n146 ) , .A1( u0_u13_u5_n171 ) );
  NOR2_X1 u0_u13_u5_U79 (.A2( u0_u13_X_31 ) , .A1( u0_u13_X_32 ) , .ZN( u0_u13_u5_n103 ) );
  NOR3_X1 u0_u13_u5_U8 (.A2( u0_u13_u5_n147 ) , .A1( u0_u13_u5_n148 ) , .ZN( u0_u13_u5_n149 ) , .A3( u0_u13_u5_n194 ) );
  NOR2_X1 u0_u13_u5_U80 (.A2( u0_u13_X_36 ) , .ZN( u0_u13_u5_n105 ) , .A1( u0_u13_u5_n180 ) );
  NOR2_X1 u0_u13_u5_U81 (.A2( u0_u13_X_33 ) , .ZN( u0_u13_u5_n108 ) , .A1( u0_u13_u5_n170 ) );
  NOR2_X1 u0_u13_u5_U82 (.A2( u0_u13_X_33 ) , .A1( u0_u13_X_36 ) , .ZN( u0_u13_u5_n107 ) );
  NOR2_X1 u0_u13_u5_U83 (.A2( u0_u13_X_31 ) , .ZN( u0_u13_u5_n104 ) , .A1( u0_u13_u5_n181 ) );
  NAND2_X1 u0_u13_u5_U84 (.A2( u0_u13_X_34 ) , .A1( u0_u13_X_35 ) , .ZN( u0_u13_u5_n153 ) );
  NAND2_X1 u0_u13_u5_U85 (.A1( u0_u13_X_34 ) , .ZN( u0_u13_u5_n126 ) , .A2( u0_u13_u5_n171 ) );
  AND2_X1 u0_u13_u5_U86 (.A1( u0_u13_X_31 ) , .A2( u0_u13_X_32 ) , .ZN( u0_u13_u5_n106 ) );
  AND2_X1 u0_u13_u5_U87 (.A1( u0_u13_X_31 ) , .ZN( u0_u13_u5_n109 ) , .A2( u0_u13_u5_n181 ) );
  INV_X1 u0_u13_u5_U88 (.A( u0_u13_X_33 ) , .ZN( u0_u13_u5_n180 ) );
  INV_X1 u0_u13_u5_U89 (.A( u0_u13_X_35 ) , .ZN( u0_u13_u5_n171 ) );
  NOR2_X1 u0_u13_u5_U9 (.ZN( u0_u13_u5_n135 ) , .A1( u0_u13_u5_n173 ) , .A2( u0_u13_u5_n176 ) );
  INV_X1 u0_u13_u5_U90 (.A( u0_u13_X_36 ) , .ZN( u0_u13_u5_n170 ) );
  INV_X1 u0_u13_u5_U91 (.A( u0_u13_X_32 ) , .ZN( u0_u13_u5_n181 ) );
  NAND4_X1 u0_u13_u5_U92 (.ZN( u0_out13_29 ) , .A4( u0_u13_u5_n129 ) , .A3( u0_u13_u5_n130 ) , .A2( u0_u13_u5_n168 ) , .A1( u0_u13_u5_n196 ) );
  AOI221_X1 u0_u13_u5_U93 (.A( u0_u13_u5_n128 ) , .ZN( u0_u13_u5_n129 ) , .C2( u0_u13_u5_n132 ) , .B2( u0_u13_u5_n159 ) , .B1( u0_u13_u5_n176 ) , .C1( u0_u13_u5_n184 ) );
  AOI222_X1 u0_u13_u5_U94 (.ZN( u0_u13_u5_n130 ) , .A2( u0_u13_u5_n146 ) , .B1( u0_u13_u5_n147 ) , .C2( u0_u13_u5_n175 ) , .B2( u0_u13_u5_n179 ) , .A1( u0_u13_u5_n188 ) , .C1( u0_u13_u5_n194 ) );
  NAND4_X1 u0_u13_u5_U95 (.ZN( u0_out13_19 ) , .A4( u0_u13_u5_n166 ) , .A3( u0_u13_u5_n167 ) , .A2( u0_u13_u5_n168 ) , .A1( u0_u13_u5_n169 ) );
  AOI22_X1 u0_u13_u5_U96 (.B2( u0_u13_u5_n145 ) , .A2( u0_u13_u5_n146 ) , .ZN( u0_u13_u5_n167 ) , .B1( u0_u13_u5_n182 ) , .A1( u0_u13_u5_n189 ) );
  NOR4_X1 u0_u13_u5_U97 (.A4( u0_u13_u5_n162 ) , .A3( u0_u13_u5_n163 ) , .A2( u0_u13_u5_n164 ) , .A1( u0_u13_u5_n165 ) , .ZN( u0_u13_u5_n166 ) );
  NAND4_X1 u0_u13_u5_U98 (.ZN( u0_out13_11 ) , .A4( u0_u13_u5_n143 ) , .A3( u0_u13_u5_n144 ) , .A2( u0_u13_u5_n169 ) , .A1( u0_u13_u5_n196 ) );
  AOI22_X1 u0_u13_u5_U99 (.A2( u0_u13_u5_n132 ) , .ZN( u0_u13_u5_n144 ) , .B2( u0_u13_u5_n145 ) , .B1( u0_u13_u5_n184 ) , .A1( u0_u13_u5_n194 ) );
  XOR2_X1 u0_u4_U1 (.B( u0_K5_9 ) , .A( u0_R3_6 ) , .Z( u0_u4_X_9 ) );
  XOR2_X1 u0_u4_U2 (.B( u0_K5_8 ) , .A( u0_R3_5 ) , .Z( u0_u4_X_8 ) );
  XOR2_X1 u0_u4_U3 (.B( u0_K5_7 ) , .A( u0_R3_4 ) , .Z( u0_u4_X_7 ) );
  XOR2_X1 u0_u4_U33 (.B( u0_K5_24 ) , .A( u0_R3_17 ) , .Z( u0_u4_X_24 ) );
  XOR2_X1 u0_u4_U34 (.B( u0_K5_23 ) , .A( u0_R3_16 ) , .Z( u0_u4_X_23 ) );
  XOR2_X1 u0_u4_U35 (.B( u0_K5_22 ) , .A( u0_R3_15 ) , .Z( u0_u4_X_22 ) );
  XOR2_X1 u0_u4_U36 (.B( u0_K5_21 ) , .A( u0_R3_14 ) , .Z( u0_u4_X_21 ) );
  XOR2_X1 u0_u4_U37 (.B( u0_K5_20 ) , .A( u0_R3_13 ) , .Z( u0_u4_X_20 ) );
  XOR2_X1 u0_u4_U39 (.B( u0_K5_19 ) , .A( u0_R3_12 ) , .Z( u0_u4_X_19 ) );
  XOR2_X1 u0_u4_U40 (.B( u0_K5_18 ) , .A( u0_R3_13 ) , .Z( u0_u4_X_18 ) );
  XOR2_X1 u0_u4_U41 (.B( u0_K5_17 ) , .A( u0_R3_12 ) , .Z( u0_u4_X_17 ) );
  XOR2_X1 u0_u4_U42 (.B( u0_K5_16 ) , .A( u0_R3_11 ) , .Z( u0_u4_X_16 ) );
  XOR2_X1 u0_u4_U43 (.B( u0_K5_15 ) , .A( u0_R3_10 ) , .Z( u0_u4_X_15 ) );
  XOR2_X1 u0_u4_U44 (.B( u0_K5_14 ) , .A( u0_R3_9 ) , .Z( u0_u4_X_14 ) );
  XOR2_X1 u0_u4_U45 (.B( u0_K5_13 ) , .A( u0_R3_8 ) , .Z( u0_u4_X_13 ) );
  XOR2_X1 u0_u4_U46 (.B( u0_K5_12 ) , .A( u0_R3_9 ) , .Z( u0_u4_X_12 ) );
  XOR2_X1 u0_u4_U47 (.B( u0_K5_11 ) , .A( u0_R3_8 ) , .Z( u0_u4_X_11 ) );
  XOR2_X1 u0_u4_U48 (.B( u0_K5_10 ) , .A( u0_R3_7 ) , .Z( u0_u4_X_10 ) );
  NOR2_X1 u0_u4_u1_U10 (.A1( u0_u4_u1_n112 ) , .A2( u0_u4_u1_n116 ) , .ZN( u0_u4_u1_n118 ) );
  NAND3_X1 u0_u4_u1_U100 (.ZN( u0_u4_u1_n113 ) , .A1( u0_u4_u1_n120 ) , .A3( u0_u4_u1_n133 ) , .A2( u0_u4_u1_n155 ) );
  OAI21_X1 u0_u4_u1_U11 (.ZN( u0_u4_u1_n101 ) , .B1( u0_u4_u1_n141 ) , .A( u0_u4_u1_n146 ) , .B2( u0_u4_u1_n183 ) );
  AOI21_X1 u0_u4_u1_U12 (.B2( u0_u4_u1_n155 ) , .B1( u0_u4_u1_n156 ) , .ZN( u0_u4_u1_n157 ) , .A( u0_u4_u1_n174 ) );
  NAND2_X1 u0_u4_u1_U13 (.ZN( u0_u4_u1_n140 ) , .A2( u0_u4_u1_n150 ) , .A1( u0_u4_u1_n155 ) );
  NAND2_X1 u0_u4_u1_U14 (.A1( u0_u4_u1_n131 ) , .ZN( u0_u4_u1_n147 ) , .A2( u0_u4_u1_n153 ) );
  INV_X1 u0_u4_u1_U15 (.A( u0_u4_u1_n139 ) , .ZN( u0_u4_u1_n174 ) );
  OR4_X1 u0_u4_u1_U16 (.A4( u0_u4_u1_n106 ) , .A3( u0_u4_u1_n107 ) , .ZN( u0_u4_u1_n108 ) , .A1( u0_u4_u1_n117 ) , .A2( u0_u4_u1_n184 ) );
  AOI21_X1 u0_u4_u1_U17 (.ZN( u0_u4_u1_n106 ) , .A( u0_u4_u1_n112 ) , .B1( u0_u4_u1_n154 ) , .B2( u0_u4_u1_n156 ) );
  AOI21_X1 u0_u4_u1_U18 (.ZN( u0_u4_u1_n107 ) , .B1( u0_u4_u1_n134 ) , .B2( u0_u4_u1_n149 ) , .A( u0_u4_u1_n174 ) );
  INV_X1 u0_u4_u1_U19 (.A( u0_u4_u1_n101 ) , .ZN( u0_u4_u1_n184 ) );
  INV_X1 u0_u4_u1_U20 (.A( u0_u4_u1_n112 ) , .ZN( u0_u4_u1_n171 ) );
  NAND2_X1 u0_u4_u1_U21 (.ZN( u0_u4_u1_n141 ) , .A1( u0_u4_u1_n153 ) , .A2( u0_u4_u1_n156 ) );
  AND2_X1 u0_u4_u1_U22 (.A1( u0_u4_u1_n123 ) , .ZN( u0_u4_u1_n134 ) , .A2( u0_u4_u1_n161 ) );
  NAND2_X1 u0_u4_u1_U23 (.A2( u0_u4_u1_n115 ) , .A1( u0_u4_u1_n116 ) , .ZN( u0_u4_u1_n148 ) );
  NAND2_X1 u0_u4_u1_U24 (.A2( u0_u4_u1_n133 ) , .A1( u0_u4_u1_n135 ) , .ZN( u0_u4_u1_n159 ) );
  NAND2_X1 u0_u4_u1_U25 (.A2( u0_u4_u1_n115 ) , .A1( u0_u4_u1_n120 ) , .ZN( u0_u4_u1_n132 ) );
  INV_X1 u0_u4_u1_U26 (.A( u0_u4_u1_n154 ) , .ZN( u0_u4_u1_n178 ) );
  INV_X1 u0_u4_u1_U27 (.A( u0_u4_u1_n151 ) , .ZN( u0_u4_u1_n183 ) );
  AND2_X1 u0_u4_u1_U28 (.A1( u0_u4_u1_n129 ) , .A2( u0_u4_u1_n133 ) , .ZN( u0_u4_u1_n149 ) );
  INV_X1 u0_u4_u1_U29 (.A( u0_u4_u1_n131 ) , .ZN( u0_u4_u1_n180 ) );
  INV_X1 u0_u4_u1_U3 (.A( u0_u4_u1_n159 ) , .ZN( u0_u4_u1_n182 ) );
  OAI221_X1 u0_u4_u1_U30 (.A( u0_u4_u1_n119 ) , .C2( u0_u4_u1_n129 ) , .ZN( u0_u4_u1_n138 ) , .B2( u0_u4_u1_n152 ) , .C1( u0_u4_u1_n174 ) , .B1( u0_u4_u1_n187 ) );
  INV_X1 u0_u4_u1_U31 (.A( u0_u4_u1_n148 ) , .ZN( u0_u4_u1_n187 ) );
  AOI211_X1 u0_u4_u1_U32 (.B( u0_u4_u1_n117 ) , .A( u0_u4_u1_n118 ) , .ZN( u0_u4_u1_n119 ) , .C2( u0_u4_u1_n146 ) , .C1( u0_u4_u1_n159 ) );
  NOR2_X1 u0_u4_u1_U33 (.A1( u0_u4_u1_n168 ) , .A2( u0_u4_u1_n176 ) , .ZN( u0_u4_u1_n98 ) );
  AOI211_X1 u0_u4_u1_U34 (.B( u0_u4_u1_n162 ) , .A( u0_u4_u1_n163 ) , .C2( u0_u4_u1_n164 ) , .ZN( u0_u4_u1_n165 ) , .C1( u0_u4_u1_n171 ) );
  AOI21_X1 u0_u4_u1_U35 (.A( u0_u4_u1_n160 ) , .B2( u0_u4_u1_n161 ) , .ZN( u0_u4_u1_n162 ) , .B1( u0_u4_u1_n182 ) );
  OR2_X1 u0_u4_u1_U36 (.A2( u0_u4_u1_n157 ) , .A1( u0_u4_u1_n158 ) , .ZN( u0_u4_u1_n163 ) );
  NAND2_X1 u0_u4_u1_U37 (.A1( u0_u4_u1_n128 ) , .ZN( u0_u4_u1_n146 ) , .A2( u0_u4_u1_n160 ) );
  NAND2_X1 u0_u4_u1_U38 (.A2( u0_u4_u1_n112 ) , .ZN( u0_u4_u1_n139 ) , .A1( u0_u4_u1_n152 ) );
  NAND2_X1 u0_u4_u1_U39 (.A1( u0_u4_u1_n105 ) , .ZN( u0_u4_u1_n156 ) , .A2( u0_u4_u1_n99 ) );
  AOI221_X1 u0_u4_u1_U4 (.A( u0_u4_u1_n138 ) , .C2( u0_u4_u1_n139 ) , .C1( u0_u4_u1_n140 ) , .B2( u0_u4_u1_n141 ) , .ZN( u0_u4_u1_n142 ) , .B1( u0_u4_u1_n175 ) );
  AOI221_X1 u0_u4_u1_U40 (.B1( u0_u4_u1_n140 ) , .ZN( u0_u4_u1_n167 ) , .B2( u0_u4_u1_n172 ) , .C2( u0_u4_u1_n175 ) , .C1( u0_u4_u1_n178 ) , .A( u0_u4_u1_n188 ) );
  INV_X1 u0_u4_u1_U41 (.ZN( u0_u4_u1_n188 ) , .A( u0_u4_u1_n97 ) );
  AOI211_X1 u0_u4_u1_U42 (.A( u0_u4_u1_n118 ) , .C1( u0_u4_u1_n132 ) , .C2( u0_u4_u1_n139 ) , .B( u0_u4_u1_n96 ) , .ZN( u0_u4_u1_n97 ) );
  AOI21_X1 u0_u4_u1_U43 (.B2( u0_u4_u1_n121 ) , .B1( u0_u4_u1_n135 ) , .A( u0_u4_u1_n152 ) , .ZN( u0_u4_u1_n96 ) );
  NOR2_X1 u0_u4_u1_U44 (.ZN( u0_u4_u1_n117 ) , .A1( u0_u4_u1_n121 ) , .A2( u0_u4_u1_n160 ) );
  OAI21_X1 u0_u4_u1_U45 (.B2( u0_u4_u1_n123 ) , .ZN( u0_u4_u1_n145 ) , .B1( u0_u4_u1_n160 ) , .A( u0_u4_u1_n185 ) );
  INV_X1 u0_u4_u1_U46 (.A( u0_u4_u1_n122 ) , .ZN( u0_u4_u1_n185 ) );
  AOI21_X1 u0_u4_u1_U47 (.B2( u0_u4_u1_n120 ) , .B1( u0_u4_u1_n121 ) , .ZN( u0_u4_u1_n122 ) , .A( u0_u4_u1_n128 ) );
  AOI21_X1 u0_u4_u1_U48 (.A( u0_u4_u1_n128 ) , .B2( u0_u4_u1_n129 ) , .ZN( u0_u4_u1_n130 ) , .B1( u0_u4_u1_n150 ) );
  NAND2_X1 u0_u4_u1_U49 (.ZN( u0_u4_u1_n112 ) , .A1( u0_u4_u1_n169 ) , .A2( u0_u4_u1_n170 ) );
  AOI211_X1 u0_u4_u1_U5 (.ZN( u0_u4_u1_n124 ) , .A( u0_u4_u1_n138 ) , .C2( u0_u4_u1_n139 ) , .B( u0_u4_u1_n145 ) , .C1( u0_u4_u1_n147 ) );
  NAND2_X1 u0_u4_u1_U50 (.ZN( u0_u4_u1_n129 ) , .A2( u0_u4_u1_n95 ) , .A1( u0_u4_u1_n98 ) );
  NAND2_X1 u0_u4_u1_U51 (.A1( u0_u4_u1_n102 ) , .ZN( u0_u4_u1_n154 ) , .A2( u0_u4_u1_n99 ) );
  NAND2_X1 u0_u4_u1_U52 (.A2( u0_u4_u1_n100 ) , .ZN( u0_u4_u1_n135 ) , .A1( u0_u4_u1_n99 ) );
  AOI21_X1 u0_u4_u1_U53 (.A( u0_u4_u1_n152 ) , .B2( u0_u4_u1_n153 ) , .B1( u0_u4_u1_n154 ) , .ZN( u0_u4_u1_n158 ) );
  INV_X1 u0_u4_u1_U54 (.A( u0_u4_u1_n160 ) , .ZN( u0_u4_u1_n175 ) );
  NAND2_X1 u0_u4_u1_U55 (.A1( u0_u4_u1_n100 ) , .ZN( u0_u4_u1_n116 ) , .A2( u0_u4_u1_n95 ) );
  NAND2_X1 u0_u4_u1_U56 (.A1( u0_u4_u1_n102 ) , .ZN( u0_u4_u1_n131 ) , .A2( u0_u4_u1_n95 ) );
  NAND2_X1 u0_u4_u1_U57 (.A2( u0_u4_u1_n104 ) , .ZN( u0_u4_u1_n121 ) , .A1( u0_u4_u1_n98 ) );
  NAND2_X1 u0_u4_u1_U58 (.A1( u0_u4_u1_n103 ) , .ZN( u0_u4_u1_n153 ) , .A2( u0_u4_u1_n98 ) );
  NAND2_X1 u0_u4_u1_U59 (.A2( u0_u4_u1_n104 ) , .A1( u0_u4_u1_n105 ) , .ZN( u0_u4_u1_n133 ) );
  AOI22_X1 u0_u4_u1_U6 (.B2( u0_u4_u1_n113 ) , .A2( u0_u4_u1_n114 ) , .ZN( u0_u4_u1_n125 ) , .A1( u0_u4_u1_n171 ) , .B1( u0_u4_u1_n173 ) );
  NAND2_X1 u0_u4_u1_U60 (.ZN( u0_u4_u1_n150 ) , .A2( u0_u4_u1_n98 ) , .A1( u0_u4_u1_n99 ) );
  NAND2_X1 u0_u4_u1_U61 (.A1( u0_u4_u1_n105 ) , .ZN( u0_u4_u1_n155 ) , .A2( u0_u4_u1_n95 ) );
  OAI21_X1 u0_u4_u1_U62 (.ZN( u0_u4_u1_n109 ) , .B1( u0_u4_u1_n129 ) , .B2( u0_u4_u1_n160 ) , .A( u0_u4_u1_n167 ) );
  NAND2_X1 u0_u4_u1_U63 (.A2( u0_u4_u1_n100 ) , .A1( u0_u4_u1_n103 ) , .ZN( u0_u4_u1_n120 ) );
  NAND2_X1 u0_u4_u1_U64 (.A1( u0_u4_u1_n102 ) , .A2( u0_u4_u1_n104 ) , .ZN( u0_u4_u1_n115 ) );
  NAND2_X1 u0_u4_u1_U65 (.A2( u0_u4_u1_n100 ) , .A1( u0_u4_u1_n104 ) , .ZN( u0_u4_u1_n151 ) );
  NAND2_X1 u0_u4_u1_U66 (.A2( u0_u4_u1_n103 ) , .A1( u0_u4_u1_n105 ) , .ZN( u0_u4_u1_n161 ) );
  INV_X1 u0_u4_u1_U67 (.A( u0_u4_u1_n152 ) , .ZN( u0_u4_u1_n173 ) );
  INV_X1 u0_u4_u1_U68 (.A( u0_u4_u1_n128 ) , .ZN( u0_u4_u1_n172 ) );
  NAND2_X1 u0_u4_u1_U69 (.A2( u0_u4_u1_n102 ) , .A1( u0_u4_u1_n103 ) , .ZN( u0_u4_u1_n123 ) );
  NAND2_X1 u0_u4_u1_U7 (.ZN( u0_u4_u1_n114 ) , .A1( u0_u4_u1_n134 ) , .A2( u0_u4_u1_n156 ) );
  NOR2_X1 u0_u4_u1_U70 (.A2( u0_u4_X_7 ) , .A1( u0_u4_X_8 ) , .ZN( u0_u4_u1_n95 ) );
  NOR2_X1 u0_u4_u1_U71 (.A1( u0_u4_X_12 ) , .A2( u0_u4_X_9 ) , .ZN( u0_u4_u1_n100 ) );
  NOR2_X1 u0_u4_u1_U72 (.A2( u0_u4_X_8 ) , .A1( u0_u4_u1_n177 ) , .ZN( u0_u4_u1_n99 ) );
  NOR2_X1 u0_u4_u1_U73 (.A2( u0_u4_X_12 ) , .ZN( u0_u4_u1_n102 ) , .A1( u0_u4_u1_n176 ) );
  NOR2_X1 u0_u4_u1_U74 (.A2( u0_u4_X_9 ) , .ZN( u0_u4_u1_n105 ) , .A1( u0_u4_u1_n168 ) );
  NAND2_X1 u0_u4_u1_U75 (.A1( u0_u4_X_10 ) , .ZN( u0_u4_u1_n160 ) , .A2( u0_u4_u1_n169 ) );
  NAND2_X1 u0_u4_u1_U76 (.A2( u0_u4_X_10 ) , .A1( u0_u4_X_11 ) , .ZN( u0_u4_u1_n152 ) );
  NAND2_X1 u0_u4_u1_U77 (.A1( u0_u4_X_11 ) , .ZN( u0_u4_u1_n128 ) , .A2( u0_u4_u1_n170 ) );
  AND2_X1 u0_u4_u1_U78 (.A2( u0_u4_X_7 ) , .A1( u0_u4_X_8 ) , .ZN( u0_u4_u1_n104 ) );
  AND2_X1 u0_u4_u1_U79 (.A1( u0_u4_X_8 ) , .ZN( u0_u4_u1_n103 ) , .A2( u0_u4_u1_n177 ) );
  AOI22_X1 u0_u4_u1_U8 (.B2( u0_u4_u1_n136 ) , .A2( u0_u4_u1_n137 ) , .ZN( u0_u4_u1_n143 ) , .A1( u0_u4_u1_n171 ) , .B1( u0_u4_u1_n173 ) );
  INV_X1 u0_u4_u1_U80 (.A( u0_u4_X_10 ) , .ZN( u0_u4_u1_n170 ) );
  INV_X1 u0_u4_u1_U81 (.A( u0_u4_X_9 ) , .ZN( u0_u4_u1_n176 ) );
  INV_X1 u0_u4_u1_U82 (.A( u0_u4_X_11 ) , .ZN( u0_u4_u1_n169 ) );
  INV_X1 u0_u4_u1_U83 (.A( u0_u4_X_12 ) , .ZN( u0_u4_u1_n168 ) );
  INV_X1 u0_u4_u1_U84 (.A( u0_u4_X_7 ) , .ZN( u0_u4_u1_n177 ) );
  NAND4_X1 u0_u4_u1_U85 (.ZN( u0_out4_28 ) , .A4( u0_u4_u1_n124 ) , .A3( u0_u4_u1_n125 ) , .A2( u0_u4_u1_n126 ) , .A1( u0_u4_u1_n127 ) );
  OAI21_X1 u0_u4_u1_U86 (.ZN( u0_u4_u1_n127 ) , .B2( u0_u4_u1_n139 ) , .B1( u0_u4_u1_n175 ) , .A( u0_u4_u1_n183 ) );
  OAI21_X1 u0_u4_u1_U87 (.ZN( u0_u4_u1_n126 ) , .B2( u0_u4_u1_n140 ) , .A( u0_u4_u1_n146 ) , .B1( u0_u4_u1_n178 ) );
  NAND4_X1 u0_u4_u1_U88 (.ZN( u0_out4_18 ) , .A4( u0_u4_u1_n165 ) , .A3( u0_u4_u1_n166 ) , .A1( u0_u4_u1_n167 ) , .A2( u0_u4_u1_n186 ) );
  AOI22_X1 u0_u4_u1_U89 (.B2( u0_u4_u1_n146 ) , .B1( u0_u4_u1_n147 ) , .A2( u0_u4_u1_n148 ) , .ZN( u0_u4_u1_n166 ) , .A1( u0_u4_u1_n172 ) );
  INV_X1 u0_u4_u1_U9 (.A( u0_u4_u1_n147 ) , .ZN( u0_u4_u1_n181 ) );
  INV_X1 u0_u4_u1_U90 (.A( u0_u4_u1_n145 ) , .ZN( u0_u4_u1_n186 ) );
  NAND4_X1 u0_u4_u1_U91 (.ZN( u0_out4_2 ) , .A4( u0_u4_u1_n142 ) , .A3( u0_u4_u1_n143 ) , .A2( u0_u4_u1_n144 ) , .A1( u0_u4_u1_n179 ) );
  OAI21_X1 u0_u4_u1_U92 (.B2( u0_u4_u1_n132 ) , .ZN( u0_u4_u1_n144 ) , .A( u0_u4_u1_n146 ) , .B1( u0_u4_u1_n180 ) );
  INV_X1 u0_u4_u1_U93 (.A( u0_u4_u1_n130 ) , .ZN( u0_u4_u1_n179 ) );
  OR4_X1 u0_u4_u1_U94 (.ZN( u0_out4_13 ) , .A4( u0_u4_u1_n108 ) , .A3( u0_u4_u1_n109 ) , .A2( u0_u4_u1_n110 ) , .A1( u0_u4_u1_n111 ) );
  AOI21_X1 u0_u4_u1_U95 (.ZN( u0_u4_u1_n111 ) , .A( u0_u4_u1_n128 ) , .B2( u0_u4_u1_n131 ) , .B1( u0_u4_u1_n135 ) );
  AOI21_X1 u0_u4_u1_U96 (.ZN( u0_u4_u1_n110 ) , .A( u0_u4_u1_n116 ) , .B1( u0_u4_u1_n152 ) , .B2( u0_u4_u1_n160 ) );
  NAND3_X1 u0_u4_u1_U97 (.A3( u0_u4_u1_n149 ) , .A2( u0_u4_u1_n150 ) , .A1( u0_u4_u1_n151 ) , .ZN( u0_u4_u1_n164 ) );
  NAND3_X1 u0_u4_u1_U98 (.A3( u0_u4_u1_n134 ) , .A2( u0_u4_u1_n135 ) , .ZN( u0_u4_u1_n136 ) , .A1( u0_u4_u1_n151 ) );
  NAND3_X1 u0_u4_u1_U99 (.A1( u0_u4_u1_n133 ) , .ZN( u0_u4_u1_n137 ) , .A2( u0_u4_u1_n154 ) , .A3( u0_u4_u1_n181 ) );
  OAI22_X1 u0_u4_u2_U10 (.ZN( u0_u4_u2_n109 ) , .A2( u0_u4_u2_n113 ) , .B2( u0_u4_u2_n133 ) , .B1( u0_u4_u2_n167 ) , .A1( u0_u4_u2_n168 ) );
  NAND3_X1 u0_u4_u2_U100 (.A2( u0_u4_u2_n100 ) , .A1( u0_u4_u2_n104 ) , .A3( u0_u4_u2_n138 ) , .ZN( u0_u4_u2_n98 ) );
  OAI22_X1 u0_u4_u2_U11 (.B1( u0_u4_u2_n151 ) , .A2( u0_u4_u2_n152 ) , .A1( u0_u4_u2_n153 ) , .ZN( u0_u4_u2_n160 ) , .B2( u0_u4_u2_n168 ) );
  NOR3_X1 u0_u4_u2_U12 (.A1( u0_u4_u2_n150 ) , .ZN( u0_u4_u2_n151 ) , .A3( u0_u4_u2_n175 ) , .A2( u0_u4_u2_n188 ) );
  AOI21_X1 u0_u4_u2_U13 (.ZN( u0_u4_u2_n144 ) , .B2( u0_u4_u2_n155 ) , .A( u0_u4_u2_n172 ) , .B1( u0_u4_u2_n185 ) );
  AOI21_X1 u0_u4_u2_U14 (.B2( u0_u4_u2_n143 ) , .ZN( u0_u4_u2_n145 ) , .B1( u0_u4_u2_n152 ) , .A( u0_u4_u2_n171 ) );
  AOI21_X1 u0_u4_u2_U15 (.B2( u0_u4_u2_n120 ) , .B1( u0_u4_u2_n121 ) , .ZN( u0_u4_u2_n126 ) , .A( u0_u4_u2_n167 ) );
  INV_X1 u0_u4_u2_U16 (.A( u0_u4_u2_n156 ) , .ZN( u0_u4_u2_n171 ) );
  INV_X1 u0_u4_u2_U17 (.A( u0_u4_u2_n120 ) , .ZN( u0_u4_u2_n188 ) );
  NAND2_X1 u0_u4_u2_U18 (.A2( u0_u4_u2_n122 ) , .ZN( u0_u4_u2_n150 ) , .A1( u0_u4_u2_n152 ) );
  INV_X1 u0_u4_u2_U19 (.A( u0_u4_u2_n153 ) , .ZN( u0_u4_u2_n170 ) );
  INV_X1 u0_u4_u2_U20 (.A( u0_u4_u2_n137 ) , .ZN( u0_u4_u2_n173 ) );
  NAND2_X1 u0_u4_u2_U21 (.A1( u0_u4_u2_n132 ) , .A2( u0_u4_u2_n139 ) , .ZN( u0_u4_u2_n157 ) );
  INV_X1 u0_u4_u2_U22 (.A( u0_u4_u2_n113 ) , .ZN( u0_u4_u2_n178 ) );
  INV_X1 u0_u4_u2_U23 (.A( u0_u4_u2_n139 ) , .ZN( u0_u4_u2_n175 ) );
  INV_X1 u0_u4_u2_U24 (.A( u0_u4_u2_n155 ) , .ZN( u0_u4_u2_n181 ) );
  INV_X1 u0_u4_u2_U25 (.A( u0_u4_u2_n119 ) , .ZN( u0_u4_u2_n177 ) );
  INV_X1 u0_u4_u2_U26 (.A( u0_u4_u2_n116 ) , .ZN( u0_u4_u2_n180 ) );
  INV_X1 u0_u4_u2_U27 (.A( u0_u4_u2_n131 ) , .ZN( u0_u4_u2_n179 ) );
  INV_X1 u0_u4_u2_U28 (.A( u0_u4_u2_n154 ) , .ZN( u0_u4_u2_n176 ) );
  NAND2_X1 u0_u4_u2_U29 (.A2( u0_u4_u2_n116 ) , .A1( u0_u4_u2_n117 ) , .ZN( u0_u4_u2_n118 ) );
  NOR2_X1 u0_u4_u2_U3 (.ZN( u0_u4_u2_n121 ) , .A2( u0_u4_u2_n177 ) , .A1( u0_u4_u2_n180 ) );
  INV_X1 u0_u4_u2_U30 (.A( u0_u4_u2_n132 ) , .ZN( u0_u4_u2_n182 ) );
  INV_X1 u0_u4_u2_U31 (.A( u0_u4_u2_n158 ) , .ZN( u0_u4_u2_n183 ) );
  OAI21_X1 u0_u4_u2_U32 (.A( u0_u4_u2_n156 ) , .B1( u0_u4_u2_n157 ) , .ZN( u0_u4_u2_n158 ) , .B2( u0_u4_u2_n179 ) );
  NOR2_X1 u0_u4_u2_U33 (.ZN( u0_u4_u2_n156 ) , .A1( u0_u4_u2_n166 ) , .A2( u0_u4_u2_n169 ) );
  NOR2_X1 u0_u4_u2_U34 (.A2( u0_u4_u2_n114 ) , .ZN( u0_u4_u2_n137 ) , .A1( u0_u4_u2_n140 ) );
  NOR2_X1 u0_u4_u2_U35 (.A2( u0_u4_u2_n138 ) , .ZN( u0_u4_u2_n153 ) , .A1( u0_u4_u2_n156 ) );
  AOI211_X1 u0_u4_u2_U36 (.ZN( u0_u4_u2_n130 ) , .C1( u0_u4_u2_n138 ) , .C2( u0_u4_u2_n179 ) , .B( u0_u4_u2_n96 ) , .A( u0_u4_u2_n97 ) );
  OAI22_X1 u0_u4_u2_U37 (.B1( u0_u4_u2_n133 ) , .A2( u0_u4_u2_n137 ) , .A1( u0_u4_u2_n152 ) , .B2( u0_u4_u2_n168 ) , .ZN( u0_u4_u2_n97 ) );
  OAI221_X1 u0_u4_u2_U38 (.B1( u0_u4_u2_n113 ) , .C1( u0_u4_u2_n132 ) , .A( u0_u4_u2_n149 ) , .B2( u0_u4_u2_n171 ) , .C2( u0_u4_u2_n172 ) , .ZN( u0_u4_u2_n96 ) );
  OAI221_X1 u0_u4_u2_U39 (.A( u0_u4_u2_n115 ) , .C2( u0_u4_u2_n123 ) , .B2( u0_u4_u2_n143 ) , .B1( u0_u4_u2_n153 ) , .ZN( u0_u4_u2_n163 ) , .C1( u0_u4_u2_n168 ) );
  INV_X1 u0_u4_u2_U4 (.A( u0_u4_u2_n134 ) , .ZN( u0_u4_u2_n185 ) );
  OAI21_X1 u0_u4_u2_U40 (.A( u0_u4_u2_n114 ) , .ZN( u0_u4_u2_n115 ) , .B1( u0_u4_u2_n176 ) , .B2( u0_u4_u2_n178 ) );
  OAI221_X1 u0_u4_u2_U41 (.A( u0_u4_u2_n135 ) , .B2( u0_u4_u2_n136 ) , .B1( u0_u4_u2_n137 ) , .ZN( u0_u4_u2_n162 ) , .C2( u0_u4_u2_n167 ) , .C1( u0_u4_u2_n185 ) );
  AND3_X1 u0_u4_u2_U42 (.A3( u0_u4_u2_n131 ) , .A2( u0_u4_u2_n132 ) , .A1( u0_u4_u2_n133 ) , .ZN( u0_u4_u2_n136 ) );
  AOI22_X1 u0_u4_u2_U43 (.ZN( u0_u4_u2_n135 ) , .B1( u0_u4_u2_n140 ) , .A1( u0_u4_u2_n156 ) , .B2( u0_u4_u2_n180 ) , .A2( u0_u4_u2_n188 ) );
  AOI21_X1 u0_u4_u2_U44 (.ZN( u0_u4_u2_n149 ) , .B1( u0_u4_u2_n173 ) , .B2( u0_u4_u2_n188 ) , .A( u0_u4_u2_n95 ) );
  AND3_X1 u0_u4_u2_U45 (.A2( u0_u4_u2_n100 ) , .A1( u0_u4_u2_n104 ) , .A3( u0_u4_u2_n156 ) , .ZN( u0_u4_u2_n95 ) );
  OAI21_X1 u0_u4_u2_U46 (.A( u0_u4_u2_n101 ) , .B2( u0_u4_u2_n121 ) , .B1( u0_u4_u2_n153 ) , .ZN( u0_u4_u2_n164 ) );
  NAND2_X1 u0_u4_u2_U47 (.A2( u0_u4_u2_n100 ) , .A1( u0_u4_u2_n107 ) , .ZN( u0_u4_u2_n155 ) );
  NAND2_X1 u0_u4_u2_U48 (.A2( u0_u4_u2_n105 ) , .A1( u0_u4_u2_n108 ) , .ZN( u0_u4_u2_n143 ) );
  NAND2_X1 u0_u4_u2_U49 (.A1( u0_u4_u2_n104 ) , .A2( u0_u4_u2_n106 ) , .ZN( u0_u4_u2_n152 ) );
  INV_X1 u0_u4_u2_U5 (.A( u0_u4_u2_n150 ) , .ZN( u0_u4_u2_n184 ) );
  NAND2_X1 u0_u4_u2_U50 (.A1( u0_u4_u2_n100 ) , .A2( u0_u4_u2_n105 ) , .ZN( u0_u4_u2_n132 ) );
  INV_X1 u0_u4_u2_U51 (.A( u0_u4_u2_n140 ) , .ZN( u0_u4_u2_n168 ) );
  INV_X1 u0_u4_u2_U52 (.A( u0_u4_u2_n138 ) , .ZN( u0_u4_u2_n167 ) );
  OAI21_X1 u0_u4_u2_U53 (.A( u0_u4_u2_n141 ) , .B2( u0_u4_u2_n142 ) , .ZN( u0_u4_u2_n146 ) , .B1( u0_u4_u2_n153 ) );
  OAI21_X1 u0_u4_u2_U54 (.A( u0_u4_u2_n140 ) , .ZN( u0_u4_u2_n141 ) , .B1( u0_u4_u2_n176 ) , .B2( u0_u4_u2_n177 ) );
  NOR3_X1 u0_u4_u2_U55 (.ZN( u0_u4_u2_n142 ) , .A3( u0_u4_u2_n175 ) , .A2( u0_u4_u2_n178 ) , .A1( u0_u4_u2_n181 ) );
  INV_X1 u0_u4_u2_U56 (.ZN( u0_u4_u2_n187 ) , .A( u0_u4_u2_n99 ) );
  OAI21_X1 u0_u4_u2_U57 (.B1( u0_u4_u2_n137 ) , .B2( u0_u4_u2_n143 ) , .A( u0_u4_u2_n98 ) , .ZN( u0_u4_u2_n99 ) );
  NAND2_X1 u0_u4_u2_U58 (.A1( u0_u4_u2_n102 ) , .A2( u0_u4_u2_n106 ) , .ZN( u0_u4_u2_n113 ) );
  NAND2_X1 u0_u4_u2_U59 (.A1( u0_u4_u2_n106 ) , .A2( u0_u4_u2_n107 ) , .ZN( u0_u4_u2_n131 ) );
  NOR4_X1 u0_u4_u2_U6 (.A4( u0_u4_u2_n124 ) , .A3( u0_u4_u2_n125 ) , .A2( u0_u4_u2_n126 ) , .A1( u0_u4_u2_n127 ) , .ZN( u0_u4_u2_n128 ) );
  NAND2_X1 u0_u4_u2_U60 (.A1( u0_u4_u2_n103 ) , .A2( u0_u4_u2_n107 ) , .ZN( u0_u4_u2_n139 ) );
  NAND2_X1 u0_u4_u2_U61 (.A1( u0_u4_u2_n103 ) , .A2( u0_u4_u2_n105 ) , .ZN( u0_u4_u2_n133 ) );
  NAND2_X1 u0_u4_u2_U62 (.A1( u0_u4_u2_n102 ) , .A2( u0_u4_u2_n103 ) , .ZN( u0_u4_u2_n154 ) );
  NAND2_X1 u0_u4_u2_U63 (.A2( u0_u4_u2_n103 ) , .A1( u0_u4_u2_n104 ) , .ZN( u0_u4_u2_n119 ) );
  NAND2_X1 u0_u4_u2_U64 (.A2( u0_u4_u2_n107 ) , .A1( u0_u4_u2_n108 ) , .ZN( u0_u4_u2_n123 ) );
  NAND2_X1 u0_u4_u2_U65 (.A1( u0_u4_u2_n104 ) , .A2( u0_u4_u2_n108 ) , .ZN( u0_u4_u2_n122 ) );
  INV_X1 u0_u4_u2_U66 (.A( u0_u4_u2_n114 ) , .ZN( u0_u4_u2_n172 ) );
  NAND2_X1 u0_u4_u2_U67 (.A2( u0_u4_u2_n100 ) , .A1( u0_u4_u2_n102 ) , .ZN( u0_u4_u2_n116 ) );
  NAND2_X1 u0_u4_u2_U68 (.A1( u0_u4_u2_n102 ) , .A2( u0_u4_u2_n108 ) , .ZN( u0_u4_u2_n120 ) );
  NAND2_X1 u0_u4_u2_U69 (.A2( u0_u4_u2_n105 ) , .A1( u0_u4_u2_n106 ) , .ZN( u0_u4_u2_n117 ) );
  AOI21_X1 u0_u4_u2_U7 (.B2( u0_u4_u2_n119 ) , .ZN( u0_u4_u2_n127 ) , .A( u0_u4_u2_n137 ) , .B1( u0_u4_u2_n155 ) );
  NOR2_X1 u0_u4_u2_U70 (.A2( u0_u4_X_16 ) , .ZN( u0_u4_u2_n140 ) , .A1( u0_u4_u2_n166 ) );
  NOR2_X1 u0_u4_u2_U71 (.A2( u0_u4_X_13 ) , .A1( u0_u4_X_14 ) , .ZN( u0_u4_u2_n100 ) );
  NOR2_X1 u0_u4_u2_U72 (.A2( u0_u4_X_16 ) , .A1( u0_u4_X_17 ) , .ZN( u0_u4_u2_n138 ) );
  NOR2_X1 u0_u4_u2_U73 (.A2( u0_u4_X_15 ) , .A1( u0_u4_X_18 ) , .ZN( u0_u4_u2_n104 ) );
  NOR2_X1 u0_u4_u2_U74 (.A2( u0_u4_X_14 ) , .ZN( u0_u4_u2_n103 ) , .A1( u0_u4_u2_n174 ) );
  NOR2_X1 u0_u4_u2_U75 (.A2( u0_u4_X_15 ) , .ZN( u0_u4_u2_n102 ) , .A1( u0_u4_u2_n165 ) );
  NOR2_X1 u0_u4_u2_U76 (.A2( u0_u4_X_17 ) , .ZN( u0_u4_u2_n114 ) , .A1( u0_u4_u2_n169 ) );
  AND2_X1 u0_u4_u2_U77 (.A1( u0_u4_X_15 ) , .ZN( u0_u4_u2_n105 ) , .A2( u0_u4_u2_n165 ) );
  AND2_X1 u0_u4_u2_U78 (.A2( u0_u4_X_15 ) , .A1( u0_u4_X_18 ) , .ZN( u0_u4_u2_n107 ) );
  AND2_X1 u0_u4_u2_U79 (.A1( u0_u4_X_14 ) , .ZN( u0_u4_u2_n106 ) , .A2( u0_u4_u2_n174 ) );
  AOI21_X1 u0_u4_u2_U8 (.ZN( u0_u4_u2_n124 ) , .B1( u0_u4_u2_n131 ) , .B2( u0_u4_u2_n143 ) , .A( u0_u4_u2_n172 ) );
  AND2_X1 u0_u4_u2_U80 (.A1( u0_u4_X_13 ) , .A2( u0_u4_X_14 ) , .ZN( u0_u4_u2_n108 ) );
  INV_X1 u0_u4_u2_U81 (.A( u0_u4_X_16 ) , .ZN( u0_u4_u2_n169 ) );
  INV_X1 u0_u4_u2_U82 (.A( u0_u4_X_17 ) , .ZN( u0_u4_u2_n166 ) );
  INV_X1 u0_u4_u2_U83 (.A( u0_u4_X_13 ) , .ZN( u0_u4_u2_n174 ) );
  INV_X1 u0_u4_u2_U84 (.A( u0_u4_X_18 ) , .ZN( u0_u4_u2_n165 ) );
  NAND4_X1 u0_u4_u2_U85 (.ZN( u0_out4_30 ) , .A4( u0_u4_u2_n147 ) , .A3( u0_u4_u2_n148 ) , .A2( u0_u4_u2_n149 ) , .A1( u0_u4_u2_n187 ) );
  NOR3_X1 u0_u4_u2_U86 (.A3( u0_u4_u2_n144 ) , .A2( u0_u4_u2_n145 ) , .A1( u0_u4_u2_n146 ) , .ZN( u0_u4_u2_n147 ) );
  AOI21_X1 u0_u4_u2_U87 (.B2( u0_u4_u2_n138 ) , .ZN( u0_u4_u2_n148 ) , .A( u0_u4_u2_n162 ) , .B1( u0_u4_u2_n182 ) );
  NAND4_X1 u0_u4_u2_U88 (.ZN( u0_out4_24 ) , .A4( u0_u4_u2_n111 ) , .A3( u0_u4_u2_n112 ) , .A1( u0_u4_u2_n130 ) , .A2( u0_u4_u2_n187 ) );
  AOI221_X1 u0_u4_u2_U89 (.A( u0_u4_u2_n109 ) , .B1( u0_u4_u2_n110 ) , .ZN( u0_u4_u2_n111 ) , .C1( u0_u4_u2_n134 ) , .C2( u0_u4_u2_n170 ) , .B2( u0_u4_u2_n173 ) );
  AOI21_X1 u0_u4_u2_U9 (.B2( u0_u4_u2_n123 ) , .ZN( u0_u4_u2_n125 ) , .A( u0_u4_u2_n171 ) , .B1( u0_u4_u2_n184 ) );
  AOI21_X1 u0_u4_u2_U90 (.ZN( u0_u4_u2_n112 ) , .B2( u0_u4_u2_n156 ) , .A( u0_u4_u2_n164 ) , .B1( u0_u4_u2_n181 ) );
  NAND4_X1 u0_u4_u2_U91 (.ZN( u0_out4_16 ) , .A4( u0_u4_u2_n128 ) , .A3( u0_u4_u2_n129 ) , .A1( u0_u4_u2_n130 ) , .A2( u0_u4_u2_n186 ) );
  AOI22_X1 u0_u4_u2_U92 (.A2( u0_u4_u2_n118 ) , .ZN( u0_u4_u2_n129 ) , .A1( u0_u4_u2_n140 ) , .B1( u0_u4_u2_n157 ) , .B2( u0_u4_u2_n170 ) );
  INV_X1 u0_u4_u2_U93 (.A( u0_u4_u2_n163 ) , .ZN( u0_u4_u2_n186 ) );
  OR4_X1 u0_u4_u2_U94 (.ZN( u0_out4_6 ) , .A4( u0_u4_u2_n161 ) , .A3( u0_u4_u2_n162 ) , .A2( u0_u4_u2_n163 ) , .A1( u0_u4_u2_n164 ) );
  OR3_X1 u0_u4_u2_U95 (.A2( u0_u4_u2_n159 ) , .A1( u0_u4_u2_n160 ) , .ZN( u0_u4_u2_n161 ) , .A3( u0_u4_u2_n183 ) );
  AOI21_X1 u0_u4_u2_U96 (.B2( u0_u4_u2_n154 ) , .B1( u0_u4_u2_n155 ) , .ZN( u0_u4_u2_n159 ) , .A( u0_u4_u2_n167 ) );
  NAND3_X1 u0_u4_u2_U97 (.A2( u0_u4_u2_n117 ) , .A1( u0_u4_u2_n122 ) , .A3( u0_u4_u2_n123 ) , .ZN( u0_u4_u2_n134 ) );
  NAND3_X1 u0_u4_u2_U98 (.ZN( u0_u4_u2_n110 ) , .A2( u0_u4_u2_n131 ) , .A3( u0_u4_u2_n139 ) , .A1( u0_u4_u2_n154 ) );
  NAND3_X1 u0_u4_u2_U99 (.A2( u0_u4_u2_n100 ) , .ZN( u0_u4_u2_n101 ) , .A1( u0_u4_u2_n104 ) , .A3( u0_u4_u2_n114 ) );
  OAI22_X1 u0_u4_u3_U10 (.B1( u0_u4_u3_n113 ) , .A2( u0_u4_u3_n135 ) , .A1( u0_u4_u3_n150 ) , .B2( u0_u4_u3_n164 ) , .ZN( u0_u4_u3_n98 ) );
  OAI211_X1 u0_u4_u3_U11 (.B( u0_u4_u3_n106 ) , .ZN( u0_u4_u3_n119 ) , .C2( u0_u4_u3_n128 ) , .C1( u0_u4_u3_n167 ) , .A( u0_u4_u3_n181 ) );
  AOI221_X1 u0_u4_u3_U12 (.C1( u0_u4_u3_n105 ) , .ZN( u0_u4_u3_n106 ) , .A( u0_u4_u3_n131 ) , .B2( u0_u4_u3_n132 ) , .C2( u0_u4_u3_n133 ) , .B1( u0_u4_u3_n169 ) );
  INV_X1 u0_u4_u3_U13 (.ZN( u0_u4_u3_n181 ) , .A( u0_u4_u3_n98 ) );
  NAND2_X1 u0_u4_u3_U14 (.ZN( u0_u4_u3_n105 ) , .A2( u0_u4_u3_n130 ) , .A1( u0_u4_u3_n155 ) );
  AOI22_X1 u0_u4_u3_U15 (.B1( u0_u4_u3_n115 ) , .A2( u0_u4_u3_n116 ) , .ZN( u0_u4_u3_n123 ) , .B2( u0_u4_u3_n133 ) , .A1( u0_u4_u3_n169 ) );
  NAND2_X1 u0_u4_u3_U16 (.ZN( u0_u4_u3_n116 ) , .A2( u0_u4_u3_n151 ) , .A1( u0_u4_u3_n182 ) );
  NOR2_X1 u0_u4_u3_U17 (.ZN( u0_u4_u3_n126 ) , .A2( u0_u4_u3_n150 ) , .A1( u0_u4_u3_n164 ) );
  AOI21_X1 u0_u4_u3_U18 (.ZN( u0_u4_u3_n112 ) , .B2( u0_u4_u3_n146 ) , .B1( u0_u4_u3_n155 ) , .A( u0_u4_u3_n167 ) );
  NAND2_X1 u0_u4_u3_U19 (.A1( u0_u4_u3_n135 ) , .ZN( u0_u4_u3_n142 ) , .A2( u0_u4_u3_n164 ) );
  NAND2_X1 u0_u4_u3_U20 (.ZN( u0_u4_u3_n132 ) , .A2( u0_u4_u3_n152 ) , .A1( u0_u4_u3_n156 ) );
  AND2_X1 u0_u4_u3_U21 (.A2( u0_u4_u3_n113 ) , .A1( u0_u4_u3_n114 ) , .ZN( u0_u4_u3_n151 ) );
  INV_X1 u0_u4_u3_U22 (.A( u0_u4_u3_n133 ) , .ZN( u0_u4_u3_n165 ) );
  INV_X1 u0_u4_u3_U23 (.A( u0_u4_u3_n135 ) , .ZN( u0_u4_u3_n170 ) );
  NAND2_X1 u0_u4_u3_U24 (.A1( u0_u4_u3_n107 ) , .A2( u0_u4_u3_n108 ) , .ZN( u0_u4_u3_n140 ) );
  NAND2_X1 u0_u4_u3_U25 (.ZN( u0_u4_u3_n117 ) , .A1( u0_u4_u3_n124 ) , .A2( u0_u4_u3_n148 ) );
  NAND2_X1 u0_u4_u3_U26 (.ZN( u0_u4_u3_n143 ) , .A1( u0_u4_u3_n165 ) , .A2( u0_u4_u3_n167 ) );
  INV_X1 u0_u4_u3_U27 (.A( u0_u4_u3_n130 ) , .ZN( u0_u4_u3_n177 ) );
  INV_X1 u0_u4_u3_U28 (.A( u0_u4_u3_n128 ) , .ZN( u0_u4_u3_n176 ) );
  INV_X1 u0_u4_u3_U29 (.A( u0_u4_u3_n155 ) , .ZN( u0_u4_u3_n174 ) );
  INV_X1 u0_u4_u3_U3 (.A( u0_u4_u3_n129 ) , .ZN( u0_u4_u3_n183 ) );
  INV_X1 u0_u4_u3_U30 (.A( u0_u4_u3_n139 ) , .ZN( u0_u4_u3_n185 ) );
  NOR2_X1 u0_u4_u3_U31 (.ZN( u0_u4_u3_n135 ) , .A2( u0_u4_u3_n141 ) , .A1( u0_u4_u3_n169 ) );
  OAI222_X1 u0_u4_u3_U32 (.C2( u0_u4_u3_n107 ) , .A2( u0_u4_u3_n108 ) , .B1( u0_u4_u3_n135 ) , .ZN( u0_u4_u3_n138 ) , .B2( u0_u4_u3_n146 ) , .C1( u0_u4_u3_n154 ) , .A1( u0_u4_u3_n164 ) );
  NOR4_X1 u0_u4_u3_U33 (.A4( u0_u4_u3_n157 ) , .A3( u0_u4_u3_n158 ) , .A2( u0_u4_u3_n159 ) , .A1( u0_u4_u3_n160 ) , .ZN( u0_u4_u3_n161 ) );
  AOI21_X1 u0_u4_u3_U34 (.B2( u0_u4_u3_n152 ) , .B1( u0_u4_u3_n153 ) , .ZN( u0_u4_u3_n158 ) , .A( u0_u4_u3_n164 ) );
  AOI21_X1 u0_u4_u3_U35 (.A( u0_u4_u3_n149 ) , .B2( u0_u4_u3_n150 ) , .B1( u0_u4_u3_n151 ) , .ZN( u0_u4_u3_n159 ) );
  AOI21_X1 u0_u4_u3_U36 (.A( u0_u4_u3_n154 ) , .B2( u0_u4_u3_n155 ) , .B1( u0_u4_u3_n156 ) , .ZN( u0_u4_u3_n157 ) );
  AOI211_X1 u0_u4_u3_U37 (.ZN( u0_u4_u3_n109 ) , .A( u0_u4_u3_n119 ) , .C2( u0_u4_u3_n129 ) , .B( u0_u4_u3_n138 ) , .C1( u0_u4_u3_n141 ) );
  AOI211_X1 u0_u4_u3_U38 (.B( u0_u4_u3_n119 ) , .A( u0_u4_u3_n120 ) , .C2( u0_u4_u3_n121 ) , .ZN( u0_u4_u3_n122 ) , .C1( u0_u4_u3_n179 ) );
  INV_X1 u0_u4_u3_U39 (.A( u0_u4_u3_n156 ) , .ZN( u0_u4_u3_n179 ) );
  INV_X1 u0_u4_u3_U4 (.A( u0_u4_u3_n140 ) , .ZN( u0_u4_u3_n182 ) );
  OAI22_X1 u0_u4_u3_U40 (.B1( u0_u4_u3_n118 ) , .ZN( u0_u4_u3_n120 ) , .A1( u0_u4_u3_n135 ) , .B2( u0_u4_u3_n154 ) , .A2( u0_u4_u3_n178 ) );
  AND3_X1 u0_u4_u3_U41 (.ZN( u0_u4_u3_n118 ) , .A2( u0_u4_u3_n124 ) , .A1( u0_u4_u3_n144 ) , .A3( u0_u4_u3_n152 ) );
  INV_X1 u0_u4_u3_U42 (.A( u0_u4_u3_n121 ) , .ZN( u0_u4_u3_n164 ) );
  NAND2_X1 u0_u4_u3_U43 (.ZN( u0_u4_u3_n133 ) , .A1( u0_u4_u3_n154 ) , .A2( u0_u4_u3_n164 ) );
  OAI211_X1 u0_u4_u3_U44 (.B( u0_u4_u3_n127 ) , .ZN( u0_u4_u3_n139 ) , .C1( u0_u4_u3_n150 ) , .C2( u0_u4_u3_n154 ) , .A( u0_u4_u3_n184 ) );
  INV_X1 u0_u4_u3_U45 (.A( u0_u4_u3_n125 ) , .ZN( u0_u4_u3_n184 ) );
  AOI221_X1 u0_u4_u3_U46 (.A( u0_u4_u3_n126 ) , .ZN( u0_u4_u3_n127 ) , .C2( u0_u4_u3_n132 ) , .C1( u0_u4_u3_n169 ) , .B2( u0_u4_u3_n170 ) , .B1( u0_u4_u3_n174 ) );
  OAI22_X1 u0_u4_u3_U47 (.A1( u0_u4_u3_n124 ) , .ZN( u0_u4_u3_n125 ) , .B2( u0_u4_u3_n145 ) , .A2( u0_u4_u3_n165 ) , .B1( u0_u4_u3_n167 ) );
  NOR2_X1 u0_u4_u3_U48 (.A1( u0_u4_u3_n113 ) , .ZN( u0_u4_u3_n131 ) , .A2( u0_u4_u3_n154 ) );
  NAND2_X1 u0_u4_u3_U49 (.A1( u0_u4_u3_n103 ) , .ZN( u0_u4_u3_n150 ) , .A2( u0_u4_u3_n99 ) );
  INV_X1 u0_u4_u3_U5 (.A( u0_u4_u3_n117 ) , .ZN( u0_u4_u3_n178 ) );
  NAND2_X1 u0_u4_u3_U50 (.A2( u0_u4_u3_n102 ) , .ZN( u0_u4_u3_n155 ) , .A1( u0_u4_u3_n97 ) );
  INV_X1 u0_u4_u3_U51 (.A( u0_u4_u3_n141 ) , .ZN( u0_u4_u3_n167 ) );
  AOI21_X1 u0_u4_u3_U52 (.B2( u0_u4_u3_n114 ) , .B1( u0_u4_u3_n146 ) , .A( u0_u4_u3_n154 ) , .ZN( u0_u4_u3_n94 ) );
  AOI21_X1 u0_u4_u3_U53 (.ZN( u0_u4_u3_n110 ) , .B2( u0_u4_u3_n142 ) , .B1( u0_u4_u3_n186 ) , .A( u0_u4_u3_n95 ) );
  INV_X1 u0_u4_u3_U54 (.A( u0_u4_u3_n145 ) , .ZN( u0_u4_u3_n186 ) );
  AOI21_X1 u0_u4_u3_U55 (.B1( u0_u4_u3_n124 ) , .A( u0_u4_u3_n149 ) , .B2( u0_u4_u3_n155 ) , .ZN( u0_u4_u3_n95 ) );
  INV_X1 u0_u4_u3_U56 (.A( u0_u4_u3_n149 ) , .ZN( u0_u4_u3_n169 ) );
  NAND2_X1 u0_u4_u3_U57 (.ZN( u0_u4_u3_n124 ) , .A1( u0_u4_u3_n96 ) , .A2( u0_u4_u3_n97 ) );
  NAND2_X1 u0_u4_u3_U58 (.A2( u0_u4_u3_n100 ) , .ZN( u0_u4_u3_n146 ) , .A1( u0_u4_u3_n96 ) );
  NAND2_X1 u0_u4_u3_U59 (.A1( u0_u4_u3_n101 ) , .ZN( u0_u4_u3_n145 ) , .A2( u0_u4_u3_n99 ) );
  AOI221_X1 u0_u4_u3_U6 (.A( u0_u4_u3_n131 ) , .C2( u0_u4_u3_n132 ) , .C1( u0_u4_u3_n133 ) , .ZN( u0_u4_u3_n134 ) , .B1( u0_u4_u3_n143 ) , .B2( u0_u4_u3_n177 ) );
  NAND2_X1 u0_u4_u3_U60 (.A1( u0_u4_u3_n100 ) , .ZN( u0_u4_u3_n156 ) , .A2( u0_u4_u3_n99 ) );
  NAND2_X1 u0_u4_u3_U61 (.A2( u0_u4_u3_n101 ) , .A1( u0_u4_u3_n104 ) , .ZN( u0_u4_u3_n148 ) );
  NAND2_X1 u0_u4_u3_U62 (.A1( u0_u4_u3_n100 ) , .A2( u0_u4_u3_n102 ) , .ZN( u0_u4_u3_n128 ) );
  NAND2_X1 u0_u4_u3_U63 (.A2( u0_u4_u3_n101 ) , .A1( u0_u4_u3_n102 ) , .ZN( u0_u4_u3_n152 ) );
  NAND2_X1 u0_u4_u3_U64 (.A2( u0_u4_u3_n101 ) , .ZN( u0_u4_u3_n114 ) , .A1( u0_u4_u3_n96 ) );
  NAND2_X1 u0_u4_u3_U65 (.ZN( u0_u4_u3_n107 ) , .A1( u0_u4_u3_n97 ) , .A2( u0_u4_u3_n99 ) );
  NAND2_X1 u0_u4_u3_U66 (.A2( u0_u4_u3_n100 ) , .A1( u0_u4_u3_n104 ) , .ZN( u0_u4_u3_n113 ) );
  NAND2_X1 u0_u4_u3_U67 (.A1( u0_u4_u3_n104 ) , .ZN( u0_u4_u3_n153 ) , .A2( u0_u4_u3_n97 ) );
  NAND2_X1 u0_u4_u3_U68 (.A2( u0_u4_u3_n103 ) , .A1( u0_u4_u3_n104 ) , .ZN( u0_u4_u3_n130 ) );
  NAND2_X1 u0_u4_u3_U69 (.A2( u0_u4_u3_n103 ) , .ZN( u0_u4_u3_n144 ) , .A1( u0_u4_u3_n96 ) );
  OAI22_X1 u0_u4_u3_U7 (.B2( u0_u4_u3_n147 ) , .A2( u0_u4_u3_n148 ) , .ZN( u0_u4_u3_n160 ) , .B1( u0_u4_u3_n165 ) , .A1( u0_u4_u3_n168 ) );
  NAND2_X1 u0_u4_u3_U70 (.A1( u0_u4_u3_n102 ) , .A2( u0_u4_u3_n103 ) , .ZN( u0_u4_u3_n108 ) );
  NOR2_X1 u0_u4_u3_U71 (.A2( u0_u4_X_19 ) , .A1( u0_u4_X_20 ) , .ZN( u0_u4_u3_n99 ) );
  NOR2_X1 u0_u4_u3_U72 (.A2( u0_u4_X_21 ) , .A1( u0_u4_X_24 ) , .ZN( u0_u4_u3_n103 ) );
  NOR2_X1 u0_u4_u3_U73 (.A2( u0_u4_X_24 ) , .A1( u0_u4_u3_n171 ) , .ZN( u0_u4_u3_n97 ) );
  NOR2_X1 u0_u4_u3_U74 (.A2( u0_u4_X_23 ) , .ZN( u0_u4_u3_n141 ) , .A1( u0_u4_u3_n166 ) );
  NOR2_X1 u0_u4_u3_U75 (.A2( u0_u4_X_19 ) , .A1( u0_u4_u3_n172 ) , .ZN( u0_u4_u3_n96 ) );
  NAND2_X1 u0_u4_u3_U76 (.A1( u0_u4_X_22 ) , .A2( u0_u4_X_23 ) , .ZN( u0_u4_u3_n154 ) );
  NAND2_X1 u0_u4_u3_U77 (.A1( u0_u4_X_23 ) , .ZN( u0_u4_u3_n149 ) , .A2( u0_u4_u3_n166 ) );
  NOR2_X1 u0_u4_u3_U78 (.A2( u0_u4_X_22 ) , .A1( u0_u4_X_23 ) , .ZN( u0_u4_u3_n121 ) );
  AND2_X1 u0_u4_u3_U79 (.A1( u0_u4_X_24 ) , .ZN( u0_u4_u3_n101 ) , .A2( u0_u4_u3_n171 ) );
  AND3_X1 u0_u4_u3_U8 (.A3( u0_u4_u3_n144 ) , .A2( u0_u4_u3_n145 ) , .A1( u0_u4_u3_n146 ) , .ZN( u0_u4_u3_n147 ) );
  AND2_X1 u0_u4_u3_U80 (.A1( u0_u4_X_19 ) , .ZN( u0_u4_u3_n102 ) , .A2( u0_u4_u3_n172 ) );
  AND2_X1 u0_u4_u3_U81 (.A1( u0_u4_X_21 ) , .A2( u0_u4_X_24 ) , .ZN( u0_u4_u3_n100 ) );
  AND2_X1 u0_u4_u3_U82 (.A2( u0_u4_X_19 ) , .A1( u0_u4_X_20 ) , .ZN( u0_u4_u3_n104 ) );
  INV_X1 u0_u4_u3_U83 (.A( u0_u4_X_22 ) , .ZN( u0_u4_u3_n166 ) );
  INV_X1 u0_u4_u3_U84 (.A( u0_u4_X_21 ) , .ZN( u0_u4_u3_n171 ) );
  INV_X1 u0_u4_u3_U85 (.A( u0_u4_X_20 ) , .ZN( u0_u4_u3_n172 ) );
  OR4_X1 u0_u4_u3_U86 (.ZN( u0_out4_10 ) , .A4( u0_u4_u3_n136 ) , .A3( u0_u4_u3_n137 ) , .A1( u0_u4_u3_n138 ) , .A2( u0_u4_u3_n139 ) );
  OAI222_X1 u0_u4_u3_U87 (.C1( u0_u4_u3_n128 ) , .ZN( u0_u4_u3_n137 ) , .B1( u0_u4_u3_n148 ) , .A2( u0_u4_u3_n150 ) , .B2( u0_u4_u3_n154 ) , .C2( u0_u4_u3_n164 ) , .A1( u0_u4_u3_n167 ) );
  OAI221_X1 u0_u4_u3_U88 (.A( u0_u4_u3_n134 ) , .B2( u0_u4_u3_n135 ) , .ZN( u0_u4_u3_n136 ) , .C1( u0_u4_u3_n149 ) , .B1( u0_u4_u3_n151 ) , .C2( u0_u4_u3_n183 ) );
  NAND4_X1 u0_u4_u3_U89 (.ZN( u0_out4_26 ) , .A4( u0_u4_u3_n109 ) , .A3( u0_u4_u3_n110 ) , .A2( u0_u4_u3_n111 ) , .A1( u0_u4_u3_n173 ) );
  INV_X1 u0_u4_u3_U9 (.A( u0_u4_u3_n143 ) , .ZN( u0_u4_u3_n168 ) );
  INV_X1 u0_u4_u3_U90 (.ZN( u0_u4_u3_n173 ) , .A( u0_u4_u3_n94 ) );
  OAI21_X1 u0_u4_u3_U91 (.ZN( u0_u4_u3_n111 ) , .B2( u0_u4_u3_n117 ) , .A( u0_u4_u3_n133 ) , .B1( u0_u4_u3_n176 ) );
  NAND4_X1 u0_u4_u3_U92 (.ZN( u0_out4_20 ) , .A4( u0_u4_u3_n122 ) , .A3( u0_u4_u3_n123 ) , .A1( u0_u4_u3_n175 ) , .A2( u0_u4_u3_n180 ) );
  INV_X1 u0_u4_u3_U93 (.A( u0_u4_u3_n126 ) , .ZN( u0_u4_u3_n180 ) );
  INV_X1 u0_u4_u3_U94 (.A( u0_u4_u3_n112 ) , .ZN( u0_u4_u3_n175 ) );
  NAND4_X1 u0_u4_u3_U95 (.ZN( u0_out4_1 ) , .A4( u0_u4_u3_n161 ) , .A3( u0_u4_u3_n162 ) , .A2( u0_u4_u3_n163 ) , .A1( u0_u4_u3_n185 ) );
  NAND2_X1 u0_u4_u3_U96 (.ZN( u0_u4_u3_n163 ) , .A2( u0_u4_u3_n170 ) , .A1( u0_u4_u3_n176 ) );
  AOI22_X1 u0_u4_u3_U97 (.B2( u0_u4_u3_n140 ) , .B1( u0_u4_u3_n141 ) , .A2( u0_u4_u3_n142 ) , .ZN( u0_u4_u3_n162 ) , .A1( u0_u4_u3_n177 ) );
  NAND3_X1 u0_u4_u3_U98 (.A1( u0_u4_u3_n114 ) , .ZN( u0_u4_u3_n115 ) , .A2( u0_u4_u3_n145 ) , .A3( u0_u4_u3_n153 ) );
  NAND3_X1 u0_u4_u3_U99 (.ZN( u0_u4_u3_n129 ) , .A2( u0_u4_u3_n144 ) , .A1( u0_u4_u3_n153 ) , .A3( u0_u4_u3_n182 ) );
  INV_X1 u0_uk_U1064 (.A( u0_key_r_6 ) , .ZN( u0_uk_n712 ) );
  INV_X1 u0_uk_U1065 (.A( u0_key_r_54 ) , .ZN( u0_uk_n673 ) );
  INV_X1 u0_uk_U1068 (.A( u0_key_r_26 ) , .ZN( u0_uk_n697 ) );
  OAI22_X1 u0_uk_U107 (.ZN( u0_K1_5 ) , .A1( u0_uk_n188 ) , .B2( u0_uk_n708 ) , .A2( u0_uk_n712 ) , .B1( u0_uk_n99 ) );
  INV_X1 u0_uk_U1070 (.A( u0_key_r_34 ) , .ZN( u0_uk_n690 ) );
  INV_X1 u0_uk_U1071 (.A( u0_key_r_27 ) , .ZN( u0_uk_n696 ) );
  INV_X1 u0_uk_U1072 (.A( u0_key_r_24 ) , .ZN( u0_uk_n699 ) );
  INV_X1 u0_uk_U1073 (.A( u0_key_r_20 ) , .ZN( u0_uk_n703 ) );
  INV_X1 u0_uk_U1078 (.A( u0_key_r_13 ) , .ZN( u0_uk_n708 ) );
  INV_X1 u0_uk_U1081 (.A( u0_key_r_19 ) , .ZN( u0_uk_n704 ) );
  INV_X1 u0_uk_U1082 (.A( u0_key_r_4 ) , .ZN( u0_uk_n713 ) );
  INV_X1 u0_uk_U1083 (.A( u0_key_r_17 ) , .ZN( u0_uk_n705 ) );
  INV_X1 u0_uk_U1084 (.A( u0_key_r_53 ) , .ZN( u0_uk_n674 ) );
  INV_X1 u0_uk_U1099 (.A( u0_key_r_40 ) , .ZN( u0_uk_n684 ) );
  INV_X1 u0_uk_U1100 (.A( u0_key_r_47 ) , .ZN( u0_uk_n679 ) );
  INV_X1 u0_uk_U1103 (.ZN( u0_K1_11 ) , .A( u0_uk_n892 ) );
  AOI22_X1 u0_uk_U1104 (.B2( u0_key_r_32 ) , .A2( u0_key_r_39 ) , .B1( u0_uk_n145 ) , .A1( u0_uk_n240 ) , .ZN( u0_uk_n892 ) );
  INV_X1 u0_uk_U1105 (.ZN( u0_K1_18 ) , .A( u0_uk_n887 ) );
  AOI22_X1 u0_uk_U1106 (.A2( u0_key_r_5 ) , .B2( u0_key_r_55 ) , .B1( u0_uk_n145 ) , .A1( u0_uk_n240 ) , .ZN( u0_uk_n887 ) );
  INV_X1 u0_uk_U1115 (.ZN( u0_K1_20 ) , .A( u0_uk_n886 ) );
  AOI22_X1 u0_uk_U1116 (.B2( u0_key_r_48 ) , .A2( u0_key_r_55 ) , .B1( u0_uk_n145 ) , .A1( u0_uk_n242 ) , .ZN( u0_uk_n886 ) );
  INV_X1 u0_uk_U1121 (.ZN( u0_K5_20 ) , .A( u0_uk_n816 ) );
  AOI22_X1 u0_uk_U1122 (.B2( u0_uk_K_r3_24 ) , .A2( u0_uk_K_r3_47 ) , .B1( u0_uk_n100 ) , .A1( u0_uk_n257 ) , .ZN( u0_uk_n816 ) );
  OAI22_X1 u0_uk_U1157 (.ZN( u0_K1_1 ) , .A1( u0_uk_n142 ) , .B1( u0_uk_n217 ) , .A2( u0_uk_n679 ) , .B2( u0_uk_n684 ) );
  OAI22_X1 u0_uk_U144 (.ZN( u0_K1_19 ) , .B1( u0_uk_n110 ) , .A1( u0_uk_n187 ) , .A2( u0_uk_n673 ) , .B2( u0_uk_n713 ) );
  INV_X1 u0_uk_U149 (.ZN( u0_K14_19 ) , .A( u0_uk_n938 ) );
  AOI22_X1 u0_uk_U150 (.B2( u0_uk_K_r12_25 ) , .A2( u0_uk_K_r12_33 ) , .B1( u0_uk_n146 ) , .A1( u0_uk_n207 ) , .ZN( u0_uk_n938 ) );
  OAI22_X1 u0_uk_U166 (.ZN( u0_K14_30 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n250 ) , .A2( u0_uk_n50 ) , .B2( u0_uk_n77 ) );
  INV_X1 u0_uk_U172 (.A( u0_key_r_25 ) , .ZN( u0_uk_n698 ) );
  OAI22_X1 u0_uk_U189 (.ZN( u0_K1_24 ) , .A1( u0_uk_n118 ) , .B1( u0_uk_n222 ) , .A2( u0_uk_n703 ) , .B2( u0_uk_n708 ) );
  OAI22_X1 u0_uk_U234 (.ZN( u0_K14_31 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n240 ) , .A2( u0_uk_n55 ) , .B2( u0_uk_n61 ) );
  OAI22_X1 u0_uk_U283 (.ZN( u0_K1_8 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n182 ) , .B2( u0_uk_n699 ) , .A2( u0_uk_n712 ) );
  OAI22_X1 u0_uk_U290 (.ZN( u0_K5_8 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n182 ) , .A2( u0_uk_n451 ) , .B2( u0_uk_n473 ) );
  OAI22_X1 u0_uk_U315 (.ZN( u0_K14_26 ) , .A1( u0_uk_n164 ) , .A2( u0_uk_n49 ) , .B2( u0_uk_n66 ) , .B1( u0_uk_n93 ) );
  NAND2_X1 u0_uk_U331 (.A1( u0_key_r_49 ) , .A2( u0_uk_n117 ) , .ZN( u0_uk_n871 ) );
  OAI21_X1 u0_uk_U349 (.ZN( u0_K1_4 ) , .B1( u0_uk_n217 ) , .B2( u0_uk_n674 ) , .A( u0_uk_n869 ) );
  NAND2_X1 u0_uk_U350 (.A1( u0_key_r_3 ) , .A2( u0_uk_n251 ) , .ZN( u0_uk_n869 ) );
  OAI22_X1 u0_uk_U373 (.ZN( u0_K14_28 ) , .A1( u0_uk_n109 ) , .B1( u0_uk_n203 ) , .A2( u0_uk_n61 ) , .B2( u0_uk_n67 ) );
  OAI22_X1 u0_uk_U387 (.ZN( u0_K14_1 ) , .A1( u0_uk_n118 ) , .B1( u0_uk_n240 ) , .A2( u0_uk_n75 ) , .B2( u0_uk_n80 ) );
  OAI22_X1 u0_uk_U391 (.ZN( u0_K1_9 ) , .B1( u0_uk_n231 ) , .A2( u0_uk_n673 ) , .B2( u0_uk_n679 ) , .A1( u0_uk_n94 ) );
  OAI22_X1 u0_uk_U444 (.ZN( u0_K14_33 ) , .A1( u0_uk_n230 ) , .A2( u0_uk_n55 ) , .B2( u0_uk_n73 ) , .B1( u0_uk_n94 ) );
  OAI21_X1 u0_uk_U472 (.ZN( u0_K14_29 ) , .B1( u0_uk_n11 ) , .B2( u0_uk_n51 ) , .A( u0_uk_n935 ) );
  NAND2_X1 u0_uk_U473 (.A1( u0_uk_K_r12_44 ) , .A2( u0_uk_n145 ) , .ZN( u0_uk_n935 ) );
  OAI22_X1 u0_uk_U488 (.ZN( u0_K14_2 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n231 ) , .A2( u0_uk_n57 ) , .B2( u0_uk_n64 ) );
  OAI21_X1 u0_uk_U495 (.ZN( u0_K1_2 ) , .B1( u0_uk_n250 ) , .B2( u0_uk_n713 ) , .A( u0_uk_n881 ) );
  NAND2_X1 u0_uk_U496 (.A1( u0_key_r_11 ) , .A2( u0_uk_n202 ) , .ZN( u0_uk_n881 ) );
  OAI21_X1 u0_uk_U499 (.ZN( u0_K1_12 ) , .B1( u0_uk_n128 ) , .B2( u0_uk_n704 ) , .A( u0_uk_n891 ) );
  NAND2_X1 u0_uk_U500 (.A1( u0_key_r_12 ) , .A2( u0_uk_n10 ) , .ZN( u0_uk_n891 ) );
  OAI21_X1 u0_uk_U524 (.ZN( u0_K5_12 ) , .B1( u0_uk_n202 ) , .B2( u0_uk_n483 ) , .A( u0_uk_n818 ) );
  NAND2_X1 u0_uk_U525 (.A1( u0_uk_K_r3_11 ) , .A2( u0_uk_n208 ) , .ZN( u0_uk_n818 ) );
  OAI22_X1 u0_uk_U538 (.ZN( u0_K14_17 ) , .A1( u0_uk_n118 ) , .B1( u0_uk_n231 ) , .A2( u0_uk_n54 ) , .B2( u0_uk_n78 ) );
  OAI22_X1 u0_uk_U539 (.ZN( u0_K5_17 ) , .B1( u0_uk_n203 ) , .A2( u0_uk_n464 ) , .B2( u0_uk_n484 ) , .A1( u0_uk_n99 ) );
  OAI22_X1 u0_uk_U545 (.ZN( u0_K14_36 ) , .A1( u0_uk_n230 ) , .A2( u0_uk_n50 ) , .B2( u0_uk_n88 ) , .B1( u0_uk_n93 ) );
  OAI22_X1 u0_uk_U570 (.ZN( u0_K5_10 ) , .B1( u0_uk_n208 ) , .A2( u0_uk_n465 ) , .B2( u0_uk_n485 ) , .A1( u0_uk_n99 ) );
  INV_X1 u0_uk_U586 (.ZN( u0_K1_10 ) , .A( u0_uk_n893 ) );
  AOI22_X1 u0_uk_U587 (.B2( u0_key_r_41 ) , .A2( u0_key_r_48 ) , .B1( u0_uk_n142 ) , .A1( u0_uk_n251 ) , .ZN( u0_uk_n893 ) );
  INV_X1 u0_uk_U599 (.ZN( u0_K5_22 ) , .A( u0_uk_n815 ) );
  INV_X1 u0_uk_U601 (.ZN( u0_K1_22 ) , .A( u0_uk_n885 ) );
  AOI22_X1 u0_uk_U602 (.B2( u0_key_r_25 ) , .A2( u0_key_r_32 ) , .B1( u0_uk_n145 ) , .A1( u0_uk_n213 ) , .ZN( u0_uk_n885 ) );
  INV_X1 u0_uk_U612 (.ZN( u0_K14_35 ) , .A( u0_uk_n933 ) );
  AOI22_X1 u0_uk_U613 (.B2( u0_uk_K_r12_1 ) , .A2( u0_uk_K_r12_7 ) , .B1( u0_uk_n141 ) , .A1( u0_uk_n220 ) , .ZN( u0_uk_n933 ) );
  OAI22_X1 u0_uk_U626 (.ZN( u0_K14_11 ) , .A1( u0_uk_n164 ) , .B2( u0_uk_n80 ) , .B1( u0_uk_n83 ) , .A2( u0_uk_n87 ) );
  OAI22_X1 u0_uk_U640 (.ZN( u0_K5_11 ) , .B1( u0_uk_n208 ) , .B2( u0_uk_n465 ) , .A2( u0_uk_n489 ) , .A1( u0_uk_n99 ) );
  INV_X1 u0_uk_U65 (.ZN( u0_K14_34 ) , .A( u0_uk_n934 ) );
  OAI22_X1 u0_uk_U656 (.ZN( u0_K1_7 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n203 ) , .A2( u0_uk_n696 ) , .B2( u0_uk_n703 ) );
  AOI22_X1 u0_uk_U66 (.B2( u0_uk_K_r12_30 ) , .A2( u0_uk_K_r12_36 ) , .B1( u0_uk_n141 ) , .A1( u0_uk_n251 ) , .ZN( u0_uk_n934 ) );
  OAI21_X1 u0_uk_U706 (.ZN( u0_K5_7 ) , .B1( u0_uk_n163 ) , .B2( u0_uk_n453 ) , .A( u0_uk_n802 ) );
  NAND2_X1 u0_uk_U707 (.A1( u0_uk_K_r3_19 ) , .A2( u0_uk_n203 ) , .ZN( u0_uk_n802 ) );
  OAI22_X1 u0_uk_U724 (.ZN( u0_K14_32 ) , .A1( u0_uk_n164 ) , .A2( u0_uk_n51 ) , .B2( u0_uk_n89 ) , .B1( u0_uk_n94 ) );
  OAI22_X1 u0_uk_U756 (.ZN( u0_K1_21 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n147 ) , .A2( u0_uk_n699 ) , .B2( u0_uk_n705 ) );
  OAI22_X1 u0_uk_U765 (.ZN( u0_K5_21 ) , .B1( u0_uk_n163 ) , .A2( u0_uk_n459 ) , .B2( u0_uk_n479 ) , .A1( u0_uk_n99 ) );
  OAI22_X1 u0_uk_U840 (.ZN( u0_K1_6 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n222 ) , .A2( u0_uk_n683 ) , .B2( u0_uk_n690 ) );
  INV_X1 u0_uk_U841 (.A( u0_key_r_41 ) , .ZN( u0_uk_n683 ) );
  OAI21_X1 u0_uk_U856 (.ZN( u0_K14_3 ) , .B1( u0_uk_n17 ) , .B2( u0_uk_n46 ) , .A( u0_uk_n932 ) );
  NAND2_X1 u0_uk_U857 (.A1( u0_uk_K_r12_47 ) , .A2( u0_uk_n63 ) , .ZN( u0_uk_n932 ) );
  OAI22_X1 u0_uk_U868 (.ZN( u0_K14_22 ) , .A1( u0_uk_n188 ) , .A2( u0_uk_n48 ) , .B2( u0_uk_n86 ) , .B1( u0_uk_n94 ) );
  OAI22_X1 u0_uk_U874 (.ZN( u0_K14_23 ) , .A1( u0_uk_n188 ) , .B2( u0_uk_n79 ) , .A2( u0_uk_n86 ) , .B1( u0_uk_n93 ) );
  OAI22_X1 u0_uk_U893 (.ZN( u0_K14_6 ) , .A1( u0_uk_n230 ) , .B2( u0_uk_n78 ) , .A2( u0_uk_n85 ) , .B1( u0_uk_n92 ) );
  OAI22_X1 u0_uk_U899 (.ZN( u0_K14_7 ) , .B1( u0_uk_n146 ) , .A1( u0_uk_n164 ) , .A2( u0_uk_n53 ) , .B2( u0_uk_n72 ) );
  OAI22_X1 u0_uk_U938 (.ZN( u0_K14_8 ) , .A1( u0_uk_n145 ) , .B1( u0_uk_n231 ) , .B2( u0_uk_n69 ) , .A2( u0_uk_n87 ) );
  OAI22_X1 u0_uk_U940 (.ZN( u0_K14_20 ) , .B1( u0_uk_n231 ) , .A2( u0_uk_n69 ) , .B2( u0_uk_n75 ) , .A1( u0_uk_n93 ) );
  OAI21_X1 u0_uk_U96 (.ZN( u0_K14_5 ) , .B1( u0_uk_n203 ) , .B2( u0_uk_n62 ) , .A( u0_uk_n927 ) );
  OAI22_X1 u0_uk_U964 (.ZN( u0_K14_16 ) , .A1( u0_uk_n17 ) , .B1( u0_uk_n231 ) , .B2( u0_uk_n46 ) , .A2( u0_uk_n84 ) );
  NAND2_X1 u0_uk_U97 (.A1( u0_uk_K_r12_10 ) , .A2( u0_uk_n251 ) , .ZN( u0_uk_n927 ) );
  OAI22_X1 u0_uk_U989 (.ZN( u0_K14_25 ) , .A1( u0_uk_n129 ) , .B1( u0_uk_n231 ) , .A2( u0_uk_n82 ) , .B2( u0_uk_n88 ) );
  OAI22_X1 u0_uk_U993 (.ZN( u0_K1_3 ) , .A1( u0_uk_n142 ) , .B1( u0_uk_n188 ) , .A2( u0_uk_n697 ) , .B2( u0_uk_n704 ) );
  XOR2_X1 u2_U10 (.B( u2_L1_29 ) , .Z( u2_N92 ) , .A( u2_out2_29 ) );
  XOR2_X1 u2_U102 (.B( u2_L12_25 ) , .Z( u2_N440 ) , .A( u2_out13_25 ) );
  XOR2_X1 u2_U109 (.B( u2_L12_19 ) , .Z( u2_N434 ) , .A( u2_out13_19 ) );
  XOR2_X1 u2_U11 (.B( u2_L1_28 ) , .Z( u2_N91 ) , .A( u2_out2_28 ) );
  XOR2_X1 u2_U114 (.B( u2_L0_12 ) , .Z( u2_N43 ) , .A( u2_out1_12 ) );
  XOR2_X1 u2_U115 (.B( u2_L12_14 ) , .Z( u2_N429 ) , .A( u2_out13_14 ) );
  XOR2_X1 u2_U118 (.B( u2_L12_11 ) , .Z( u2_N426 ) , .A( u2_out13_11 ) );
  XOR2_X1 u2_U12 (.B( u2_L1_27 ) , .Z( u2_N90 ) , .A( u2_out2_27 ) );
  XOR2_X1 u2_U121 (.B( u2_L12_8 ) , .Z( u2_N423 ) , .A( u2_out13_8 ) );
  XOR2_X1 u2_U126 (.B( u2_L12_4 ) , .Z( u2_N419 ) , .A( u2_out13_4 ) );
  XOR2_X1 u2_U127 (.B( u2_L12_3 ) , .Z( u2_N418 ) , .A( u2_out13_3 ) );
  XOR2_X1 u2_U13 (.Z( u2_N9 ) , .B( u2_desIn_r_12 ) , .A( u2_out0_10 ) );
  XOR2_X1 u2_U14 (.B( u2_L1_26 ) , .Z( u2_N89 ) , .A( u2_out2_26 ) );
  XOR2_X1 u2_U159 (.B( u2_L0_8 ) , .Z( u2_N39 ) , .A( u2_out1_8 ) );
  XOR2_X1 u2_U16 (.B( u2_L1_24 ) , .Z( u2_N87 ) , .A( u2_out2_24 ) );
  XOR2_X1 u2_U167 (.B( u2_L10_31 ) , .Z( u2_N382 ) , .A( u2_out11_31 ) );
  XOR2_X1 u2_U168 (.B( u2_L10_30 ) , .Z( u2_N381 ) , .A( u2_out11_30 ) );
  XOR2_X1 u2_U17 (.B( u2_L1_23 ) , .Z( u2_N86 ) , .A( u2_out2_23 ) );
  XOR2_X1 u2_U170 (.B( u2_L0_7 ) , .Z( u2_N38 ) , .A( u2_out1_7 ) );
  XOR2_X1 u2_U171 (.B( u2_L10_28 ) , .Z( u2_N379 ) , .A( u2_out11_28 ) );
  XOR2_X1 u2_U175 (.B( u2_L10_24 ) , .Z( u2_N375 ) , .A( u2_out11_24 ) );
  XOR2_X1 u2_U176 (.B( u2_L10_23 ) , .Z( u2_N374 ) , .A( u2_out11_23 ) );
  XOR2_X1 u2_U18 (.B( u2_L1_22 ) , .Z( u2_N85 ) , .A( u2_out2_22 ) );
  XOR2_X1 u2_U182 (.B( u2_L10_18 ) , .Z( u2_N369 ) , .A( u2_out11_18 ) );
  XOR2_X1 u2_U183 (.B( u2_L10_17 ) , .Z( u2_N368 ) , .A( u2_out11_17 ) );
  XOR2_X1 u2_U184 (.B( u2_L10_16 ) , .Z( u2_N367 ) , .A( u2_out11_16 ) );
  XOR2_X1 u2_U187 (.B( u2_L10_13 ) , .Z( u2_N364 ) , .A( u2_out11_13 ) );
  XOR2_X1 u2_U19 (.B( u2_L1_21 ) , .Z( u2_N84 ) , .A( u2_out2_21 ) );
  XOR2_X1 u2_U191 (.B( u2_L10_9 ) , .Z( u2_N360 ) , .A( u2_out11_9 ) );
  XOR2_X1 u2_U195 (.B( u2_L10_6 ) , .Z( u2_N357 ) , .A( u2_out11_6 ) );
  XOR2_X1 u2_U199 (.B( u2_L10_2 ) , .Z( u2_N353 ) , .A( u2_out11_2 ) );
  XOR2_X1 u2_U20 (.B( u2_L1_20 ) , .Z( u2_N83 ) , .A( u2_out2_20 ) );
  XOR2_X1 u2_U21 (.B( u2_L1_19 ) , .Z( u2_N82 ) , .A( u2_out2_19 ) );
  XOR2_X1 u2_U214 (.B( u2_L0_3 ) , .Z( u2_N34 ) , .A( u2_out1_3 ) );
  XOR2_X1 u2_U22 (.B( u2_L1_18 ) , .Z( u2_N81 ) , .A( u2_out2_18 ) );
  XOR2_X1 u2_U23 (.B( u2_L1_17 ) , .Z( u2_N80 ) , .A( u2_out2_17 ) );
  XOR2_X1 u2_U238 (.B( u2_L8_31 ) , .Z( u2_N318 ) , .A( u2_out9_31 ) );
  XOR2_X1 u2_U239 (.B( u2_L8_30 ) , .Z( u2_N317 ) , .A( u2_out9_30 ) );
  XOR2_X1 u2_U24 (.Z( u2_N8 ) , .B( u2_desIn_r_4 ) , .A( u2_out0_9 ) );
  XOR2_X1 u2_U241 (.B( u2_L8_28 ) , .Z( u2_N315 ) , .A( u2_out9_28 ) );
  XOR2_X1 u2_U242 (.B( u2_L8_27 ) , .Z( u2_N314 ) , .A( u2_out9_27 ) );
  XOR2_X1 u2_U245 (.B( u2_L8_24 ) , .Z( u2_N311 ) , .A( u2_out9_24 ) );
  XOR2_X1 u2_U246 (.B( u2_L8_23 ) , .Z( u2_N310 ) , .A( u2_out9_23 ) );
  XOR2_X1 u2_U249 (.B( u2_L8_21 ) , .Z( u2_N308 ) , .A( u2_out9_21 ) );
  XOR2_X1 u2_U25 (.B( u2_L1_16 ) , .Z( u2_N79 ) , .A( u2_out2_16 ) );
  XOR2_X1 u2_U252 (.B( u2_L8_18 ) , .Z( u2_N305 ) , .A( u2_out9_18 ) );
  XOR2_X1 u2_U253 (.B( u2_L8_17 ) , .Z( u2_N304 ) , .A( u2_out9_17 ) );
  XOR2_X1 u2_U254 (.B( u2_L8_16 ) , .Z( u2_N303 ) , .A( u2_out9_16 ) );
  XOR2_X1 u2_U255 (.B( u2_L8_15 ) , .Z( u2_N302 ) , .A( u2_out9_15 ) );
  XOR2_X1 u2_U257 (.B( u2_L8_13 ) , .Z( u2_N300 ) , .A( u2_out9_13 ) );
  XOR2_X1 u2_U258 (.Z( u2_N30 ) , .B( u2_desIn_r_48 ) , .A( u2_out0_31 ) );
  XOR2_X1 u2_U26 (.B( u2_L1_15 ) , .Z( u2_N78 ) , .A( u2_out2_15 ) );
  XOR2_X1 u2_U263 (.B( u2_L8_9 ) , .Z( u2_N296 ) , .A( u2_out9_9 ) );
  XOR2_X1 u2_U266 (.B( u2_L8_6 ) , .Z( u2_N293 ) , .A( u2_out9_6 ) );
  XOR2_X1 u2_U267 (.B( u2_L8_5 ) , .Z( u2_N292 ) , .A( u2_out9_5 ) );
  XOR2_X1 u2_U270 (.Z( u2_N29 ) , .B( u2_desIn_r_40 ) , .A( u2_out0_30 ) );
  XOR2_X1 u2_U271 (.B( u2_L8_2 ) , .Z( u2_N289 ) , .A( u2_out9_2 ) );
  XOR2_X1 u2_U28 (.B( u2_L1_13 ) , .Z( u2_N76 ) , .A( u2_out2_13 ) );
  XOR2_X1 u2_U29 (.B( u2_L1_12 ) , .Z( u2_N75 ) , .A( u2_out2_12 ) );
  XOR2_X1 u2_U292 (.Z( u2_N27 ) , .B( u2_desIn_r_24 ) , .A( u2_out0_28 ) );
  XOR2_X1 u2_U3 (.B( u2_L2_4 ) , .Z( u2_N99 ) , .A( u2_out3_4 ) );
  XOR2_X1 u2_U30 (.B( u2_L1_11 ) , .Z( u2_N74 ) , .A( u2_out2_11 ) );
  XOR2_X1 u2_U308 (.B( u2_L6_32 ) , .Z( u2_N255 ) , .A( u2_out7_32 ) );
  XOR2_X1 u2_U31 (.B( u2_L1_10 ) , .Z( u2_N73 ) , .A( u2_out2_10 ) );
  XOR2_X1 u2_U313 (.B( u2_L6_27 ) , .Z( u2_N250 ) , .A( u2_out7_27 ) );
  XOR2_X1 u2_U314 (.Z( u2_N25 ) , .B( u2_desIn_r_8 ) , .A( u2_out0_26 ) );
  XOR2_X1 u2_U319 (.B( u2_L6_22 ) , .Z( u2_N245 ) , .A( u2_out7_22 ) );
  XOR2_X1 u2_U32 (.B( u2_L1_9 ) , .Z( u2_N72 ) , .A( u2_out2_9 ) );
  XOR2_X1 u2_U320 (.B( u2_L6_21 ) , .Z( u2_N244 ) , .A( u2_out7_21 ) );
  XOR2_X1 u2_U327 (.B( u2_L6_15 ) , .Z( u2_N238 ) , .A( u2_out7_15 ) );
  XOR2_X1 u2_U330 (.B( u2_L6_12 ) , .Z( u2_N235 ) , .A( u2_out7_12 ) );
  XOR2_X1 u2_U335 (.B( u2_L6_7 ) , .Z( u2_N230 ) , .A( u2_out7_7 ) );
  XOR2_X1 u2_U336 (.Z( u2_N23 ) , .B( u2_desIn_r_58 ) , .A( u2_out0_24 ) );
  XOR2_X1 u2_U338 (.B( u2_L6_5 ) , .Z( u2_N228 ) , .A( u2_out7_5 ) );
  XOR2_X1 u2_U34 (.B( u2_L1_7 ) , .Z( u2_N70 ) , .A( u2_out2_7 ) );
  XOR2_X1 u2_U343 (.B( u2_L5_32 ) , .Z( u2_N223 ) , .A( u2_out6_32 ) );
  XOR2_X1 u2_U344 (.B( u2_L5_31 ) , .Z( u2_N222 ) , .A( u2_out6_31 ) );
  XOR2_X1 u2_U345 (.B( u2_L5_30 ) , .Z( u2_N221 ) , .A( u2_out6_30 ) );
  XOR2_X1 u2_U347 (.Z( u2_N22 ) , .B( u2_desIn_r_50 ) , .A( u2_out0_23 ) );
  XOR2_X1 u2_U348 (.B( u2_L5_28 ) , .Z( u2_N219 ) , .A( u2_out6_28 ) );
  XOR2_X1 u2_U349 (.B( u2_L5_27 ) , .Z( u2_N218 ) , .A( u2_out6_27 ) );
  XOR2_X1 u2_U350 (.B( u2_L5_26 ) , .Z( u2_N217 ) , .A( u2_out6_26 ) );
  XOR2_X1 u2_U351 (.B( u2_L5_25 ) , .Z( u2_N216 ) , .A( u2_out6_25 ) );
  XOR2_X1 u2_U352 (.B( u2_L5_24 ) , .Z( u2_N215 ) , .A( u2_out6_24 ) );
  XOR2_X1 u2_U353 (.B( u2_L5_23 ) , .Z( u2_N214 ) , .A( u2_out6_23 ) );
  XOR2_X1 u2_U354 (.B( u2_L5_22 ) , .Z( u2_N213 ) , .A( u2_out6_22 ) );
  XOR2_X1 u2_U355 (.B( u2_L5_21 ) , .Z( u2_N212 ) , .A( u2_out6_21 ) );
  XOR2_X1 u2_U356 (.B( u2_L5_20 ) , .Z( u2_N211 ) , .A( u2_out6_20 ) );
  XOR2_X1 u2_U359 (.B( u2_L5_18 ) , .Z( u2_N209 ) , .A( u2_out6_18 ) );
  XOR2_X1 u2_U36 (.B( u2_L1_6 ) , .Z( u2_N69 ) , .A( u2_out2_6 ) );
  XOR2_X1 u2_U360 (.B( u2_L5_17 ) , .Z( u2_N208 ) , .A( u2_out6_17 ) );
  XOR2_X1 u2_U361 (.B( u2_L5_16 ) , .Z( u2_N207 ) , .A( u2_out6_16 ) );
  XOR2_X1 u2_U362 (.B( u2_L5_15 ) , .Z( u2_N206 ) , .A( u2_out6_15 ) );
  XOR2_X1 u2_U363 (.B( u2_L5_14 ) , .Z( u2_N205 ) , .A( u2_out6_14 ) );
  XOR2_X1 u2_U364 (.B( u2_L5_13 ) , .Z( u2_N204 ) , .A( u2_out6_13 ) );
  XOR2_X1 u2_U365 (.B( u2_L5_12 ) , .Z( u2_N203 ) , .A( u2_out6_12 ) );
  XOR2_X1 u2_U367 (.B( u2_L5_10 ) , .Z( u2_N201 ) , .A( u2_out6_10 ) );
  XOR2_X1 u2_U368 (.B( u2_L5_9 ) , .Z( u2_N200 ) , .A( u2_out6_9 ) );
  XOR2_X1 u2_U37 (.B( u2_L1_5 ) , .Z( u2_N68 ) , .A( u2_out2_5 ) );
  XOR2_X1 u2_U371 (.B( u2_L5_8 ) , .Z( u2_N199 ) , .A( u2_out6_8 ) );
  XOR2_X1 u2_U372 (.B( u2_L5_7 ) , .Z( u2_N198 ) , .A( u2_out6_7 ) );
  XOR2_X1 u2_U373 (.B( u2_L5_6 ) , .Z( u2_N197 ) , .A( u2_out6_6 ) );
  XOR2_X1 u2_U374 (.B( u2_L5_5 ) , .Z( u2_N196 ) , .A( u2_out6_5 ) );
  XOR2_X1 u2_U376 (.B( u2_L5_3 ) , .Z( u2_N194 ) , .A( u2_out6_3 ) );
  XOR2_X1 u2_U377 (.B( u2_L5_2 ) , .Z( u2_N193 ) , .A( u2_out6_2 ) );
  XOR2_X1 u2_U378 (.B( u2_L5_1 ) , .Z( u2_N192 ) , .A( u2_out6_1 ) );
  XOR2_X1 u2_U38 (.B( u2_L1_4 ) , .Z( u2_N67 ) , .A( u2_out2_4 ) );
  XOR2_X1 u2_U381 (.Z( u2_N19 ) , .B( u2_desIn_r_26 ) , .A( u2_out0_20 ) );
  XOR2_X1 u2_U386 (.B( u2_L4_26 ) , .Z( u2_N185 ) , .A( u2_out5_26 ) );
  XOR2_X1 u2_U387 (.B( u2_L4_25 ) , .Z( u2_N184 ) , .A( u2_out5_25 ) );
  XOR2_X1 u2_U393 (.B( u2_L4_20 ) , .Z( u2_N179 ) , .A( u2_out5_20 ) );
  XOR2_X1 u2_U399 (.B( u2_L4_14 ) , .Z( u2_N173 ) , .A( u2_out5_14 ) );
  XOR2_X1 u2_U4 (.B( u2_L2_3 ) , .Z( u2_N98 ) , .A( u2_out3_3 ) );
  XOR2_X1 u2_U40 (.B( u2_L1_2 ) , .Z( u2_N65 ) , .A( u2_out2_2 ) );
  XOR2_X1 u2_U403 (.Z( u2_N17 ) , .B( u2_desIn_r_10 ) , .A( u2_out0_18 ) );
  XOR2_X1 u2_U404 (.B( u2_L4_10 ) , .Z( u2_N169 ) , .A( u2_out5_10 ) );
  XOR2_X1 u2_U406 (.B( u2_L4_8 ) , .Z( u2_N167 ) , .A( u2_out5_8 ) );
  XOR2_X1 u2_U41 (.B( u2_L1_1 ) , .Z( u2_N64 ) , .A( u2_out2_1 ) );
  XOR2_X1 u2_U411 (.B( u2_L4_3 ) , .Z( u2_N162 ) , .A( u2_out5_3 ) );
  XOR2_X1 u2_U413 (.B( u2_L4_1 ) , .Z( u2_N160 ) , .A( u2_out5_1 ) );
  XOR2_X1 u2_U414 (.Z( u2_N16 ) , .B( u2_desIn_r_2 ) , .A( u2_out0_17 ) );
  XOR2_X1 u2_U417 (.B( u2_L3_30 ) , .Z( u2_N157 ) , .A( u2_out4_30 ) );
  XOR2_X1 u2_U419 (.B( u2_L3_28 ) , .Z( u2_N155 ) , .A( u2_out4_28 ) );
  XOR2_X1 u2_U42 (.B( u2_L0_32 ) , .Z( u2_N63 ) , .A( u2_out1_32 ) );
  XOR2_X1 u2_U421 (.B( u2_L3_26 ) , .Z( u2_N153 ) , .A( u2_out4_26 ) );
  XOR2_X1 u2_U423 (.B( u2_L3_24 ) , .Z( u2_N151 ) , .A( u2_out4_24 ) );
  XOR2_X1 u2_U425 (.Z( u2_N15 ) , .B( u2_desIn_r_60 ) , .A( u2_out0_16 ) );
  XOR2_X1 u2_U428 (.B( u2_L3_20 ) , .Z( u2_N147 ) , .A( u2_out4_20 ) );
  XOR2_X1 u2_U430 (.B( u2_L3_18 ) , .Z( u2_N145 ) , .A( u2_out4_18 ) );
  XOR2_X1 u2_U432 (.B( u2_L3_16 ) , .Z( u2_N143 ) , .A( u2_out4_16 ) );
  XOR2_X1 u2_U435 (.B( u2_L3_13 ) , .Z( u2_N140 ) , .A( u2_out4_13 ) );
  XOR2_X1 u2_U439 (.B( u2_L3_10 ) , .Z( u2_N137 ) , .A( u2_out4_10 ) );
  XOR2_X1 u2_U443 (.B( u2_L3_6 ) , .Z( u2_N133 ) , .A( u2_out4_6 ) );
  XOR2_X1 u2_U448 (.B( u2_L3_2 ) , .Z( u2_N129 ) , .A( u2_out4_2 ) );
  XOR2_X1 u2_U449 (.B( u2_L3_1 ) , .Z( u2_N128 ) , .A( u2_out4_1 ) );
  XOR2_X1 u2_U452 (.B( u2_L2_30 ) , .Z( u2_N125 ) , .A( u2_out3_30 ) );
  XOR2_X1 u2_U453 (.B( u2_L2_29 ) , .Z( u2_N124 ) , .A( u2_out3_29 ) );
  XOR2_X1 u2_U456 (.B( u2_L2_26 ) , .Z( u2_N121 ) , .A( u2_out3_26 ) );
  XOR2_X1 u2_U457 (.B( u2_L2_25 ) , .Z( u2_N120 ) , .A( u2_out3_25 ) );
  XOR2_X1 u2_U458 (.Z( u2_N12 ) , .B( u2_desIn_r_36 ) , .A( u2_out0_13 ) );
  XOR2_X1 u2_U459 (.B( u2_L2_24 ) , .Z( u2_N119 ) , .A( u2_out3_24 ) );
  XOR2_X1 u2_U463 (.B( u2_L2_20 ) , .Z( u2_N115 ) , .A( u2_out3_20 ) );
  XOR2_X1 u2_U464 (.B( u2_L2_19 ) , .Z( u2_N114 ) , .A( u2_out3_19 ) );
  XOR2_X1 u2_U467 (.B( u2_L2_16 ) , .Z( u2_N111 ) , .A( u2_out3_16 ) );
  XOR2_X1 u2_U470 (.B( u2_L2_14 ) , .Z( u2_N109 ) , .A( u2_out3_14 ) );
  XOR2_X1 u2_U473 (.B( u2_L2_11 ) , .Z( u2_N106 ) , .A( u2_out3_11 ) );
  XOR2_X1 u2_U474 (.B( u2_L2_10 ) , .Z( u2_N105 ) , .A( u2_out3_10 ) );
  XOR2_X1 u2_U476 (.B( u2_L2_8 ) , .Z( u2_N103 ) , .A( u2_out3_8 ) );
  XOR2_X1 u2_U478 (.B( u2_L2_6 ) , .Z( u2_N101 ) , .A( u2_out3_6 ) );
  XOR2_X1 u2_U481 (.Z( u2_N1 ) , .B( u2_desIn_r_14 ) , .A( u2_out0_2 ) );
  XOR2_X1 u2_U482 (.Z( u2_N0 ) , .B( u2_desIn_r_6 ) , .A( u2_out0_1 ) );
  XOR2_X1 u2_U483 (.Z( u2_FP_9 ) , .B( u2_L14_9 ) , .A( u2_out15_9 ) );
  XOR2_X1 u2_U484 (.Z( u2_FP_8 ) , .B( u2_L14_8 ) , .A( u2_out15_8 ) );
  XOR2_X1 u2_U485 (.Z( u2_FP_7 ) , .B( u2_L14_7 ) , .A( u2_out15_7 ) );
  XOR2_X1 u2_U487 (.Z( u2_FP_5 ) , .B( u2_L14_5 ) , .A( u2_out15_5 ) );
  XOR2_X1 u2_U488 (.Z( u2_FP_4 ) , .B( u2_L14_4 ) , .A( u2_out15_4 ) );
  XOR2_X1 u2_U489 (.Z( u2_FP_3 ) , .B( u2_L14_3 ) , .A( u2_out15_3 ) );
  XOR2_X1 u2_U490 (.Z( u2_FP_32 ) , .B( u2_L14_32 ) , .A( u2_out15_32 ) );
  XOR2_X1 u2_U491 (.Z( u2_FP_31 ) , .B( u2_L14_31 ) , .A( u2_out15_31 ) );
  XOR2_X1 u2_U494 (.Z( u2_FP_29 ) , .B( u2_L14_29 ) , .A( u2_out15_29 ) );
  XOR2_X1 u2_U496 (.Z( u2_FP_27 ) , .B( u2_L14_27 ) , .A( u2_out15_27 ) );
  XOR2_X1 u2_U498 (.Z( u2_FP_25 ) , .B( u2_L14_25 ) , .A( u2_out15_25 ) );
  XOR2_X1 u2_U50 (.B( u2_L0_25 ) , .Z( u2_N56 ) , .A( u2_out1_25 ) );
  XOR2_X1 u2_U500 (.Z( u2_FP_23 ) , .B( u2_L14_23 ) , .A( u2_out15_23 ) );
  XOR2_X1 u2_U501 (.Z( u2_FP_22 ) , .B( u2_L14_22 ) , .A( u2_out15_22 ) );
  XOR2_X1 u2_U502 (.Z( u2_FP_21 ) , .B( u2_L14_21 ) , .A( u2_out15_21 ) );
  XOR2_X1 u2_U505 (.Z( u2_FP_19 ) , .B( u2_L14_19 ) , .A( u2_out15_19 ) );
  XOR2_X1 u2_U507 (.Z( u2_FP_17 ) , .B( u2_L14_17 ) , .A( u2_out15_17 ) );
  XOR2_X1 u2_U509 (.Z( u2_FP_15 ) , .B( u2_L14_15 ) , .A( u2_out15_15 ) );
  XOR2_X1 u2_U510 (.Z( u2_FP_14 ) , .B( u2_L14_14 ) , .A( u2_out15_14 ) );
  XOR2_X1 u2_U512 (.Z( u2_FP_12 ) , .B( u2_L14_12 ) , .A( u2_out15_12 ) );
  XOR2_X1 u2_U513 (.Z( u2_FP_11 ) , .B( u2_L14_11 ) , .A( u2_out15_11 ) );
  XOR2_X1 u2_U53 (.B( u2_L0_22 ) , .Z( u2_N53 ) , .A( u2_out1_22 ) );
  XOR2_X1 u2_U57 (.Z( u2_N5 ) , .B( u2_desIn_r_46 ) , .A( u2_out0_6 ) );
  XOR2_X1 u2_U6 (.B( u2_L2_1 ) , .Z( u2_N96 ) , .A( u2_out3_1 ) );
  XOR2_X1 u2_U60 (.B( u2_L13_32 ) , .Z( u2_N479 ) , .A( u2_out14_32 ) );
  XOR2_X1 u2_U61 (.B( u2_L13_31 ) , .Z( u2_N478 ) , .A( u2_out14_31 ) );
  XOR2_X1 u2_U63 (.B( u2_L13_29 ) , .Z( u2_N476 ) , .A( u2_out14_29 ) );
  XOR2_X1 u2_U64 (.B( u2_L13_28 ) , .Z( u2_N475 ) , .A( u2_out14_28 ) );
  XOR2_X1 u2_U67 (.B( u2_L13_25 ) , .Z( u2_N472 ) , .A( u2_out14_25 ) );
  XOR2_X1 u2_U69 (.B( u2_L13_23 ) , .Z( u2_N470 ) , .A( u2_out14_23 ) );
  XOR2_X1 u2_U7 (.B( u2_L1_32 ) , .Z( u2_N95 ) , .A( u2_out2_32 ) );
  XOR2_X1 u2_U71 (.B( u2_L13_22 ) , .Z( u2_N469 ) , .A( u2_out14_22 ) );
  XOR2_X1 u2_U74 (.B( u2_L13_19 ) , .Z( u2_N466 ) , .A( u2_out14_19 ) );
  XOR2_X1 u2_U75 (.B( u2_L13_18 ) , .Z( u2_N465 ) , .A( u2_out14_18 ) );
  XOR2_X1 u2_U76 (.B( u2_L13_17 ) , .Z( u2_N464 ) , .A( u2_out14_17 ) );
  XOR2_X1 u2_U79 (.B( u2_L13_14 ) , .Z( u2_N461 ) , .A( u2_out14_14 ) );
  XOR2_X1 u2_U8 (.B( u2_L1_31 ) , .Z( u2_N94 ) , .A( u2_out2_31 ) );
  XOR2_X1 u2_U80 (.B( u2_L13_13 ) , .Z( u2_N460 ) , .A( u2_out14_13 ) );
  XOR2_X1 u2_U82 (.B( u2_L13_12 ) , .Z( u2_N459 ) , .A( u2_out14_12 ) );
  XOR2_X1 u2_U83 (.B( u2_L13_11 ) , .Z( u2_N458 ) , .A( u2_out14_11 ) );
  XOR2_X1 u2_U85 (.B( u2_L13_9 ) , .Z( u2_N456 ) , .A( u2_out14_9 ) );
  XOR2_X1 u2_U86 (.B( u2_L13_8 ) , .Z( u2_N455 ) , .A( u2_out14_8 ) );
  XOR2_X1 u2_U87 (.B( u2_L13_7 ) , .Z( u2_N454 ) , .A( u2_out14_7 ) );
  XOR2_X1 u2_U9 (.B( u2_L1_30 ) , .Z( u2_N93 ) , .A( u2_out2_30 ) );
  XOR2_X1 u2_U90 (.B( u2_L13_4 ) , .Z( u2_N451 ) , .A( u2_out14_4 ) );
  XOR2_X1 u2_U91 (.B( u2_L13_3 ) , .Z( u2_N450 ) , .A( u2_out14_3 ) );
  XOR2_X1 u2_U92 (.B( u2_L0_14 ) , .Z( u2_N45 ) , .A( u2_out1_14 ) );
  XOR2_X1 u2_U93 (.B( u2_L13_2 ) , .Z( u2_N449 ) , .A( u2_out14_2 ) );
  XOR2_X1 u2_U98 (.B( u2_L12_29 ) , .Z( u2_N444 ) , .A( u2_out13_29 ) );
  XOR2_X1 u2_u0_U1 (.B( u2_K1_9 ) , .A( u2_desIn_r_47 ) , .Z( u2_u0_X_9 ) );
  XOR2_X1 u2_u0_U16 (.B( u2_K1_3 ) , .A( u2_desIn_r_15 ) , .Z( u2_u0_X_3 ) );
  XOR2_X1 u2_u0_U2 (.B( u2_K1_8 ) , .A( u2_desIn_r_39 ) , .Z( u2_u0_X_8 ) );
  XOR2_X1 u2_u0_U27 (.B( u2_K1_2 ) , .A( u2_desIn_r_7 ) , .Z( u2_u0_X_2 ) );
  XOR2_X1 u2_u0_U3 (.B( u2_K1_7 ) , .A( u2_desIn_r_31 ) , .Z( u2_u0_X_7 ) );
  XOR2_X1 u2_u0_U33 (.B( u2_K1_24 ) , .A( u2_desIn_r_3 ) , .Z( u2_u0_X_24 ) );
  XOR2_X1 u2_u0_U34 (.B( u2_K1_23 ) , .A( u2_desIn_r_61 ) , .Z( u2_u0_X_23 ) );
  XOR2_X1 u2_u0_U35 (.B( u2_K1_22 ) , .A( u2_desIn_r_53 ) , .Z( u2_u0_X_22 ) );
  XOR2_X1 u2_u0_U36 (.B( u2_K1_21 ) , .A( u2_desIn_r_45 ) , .Z( u2_u0_X_21 ) );
  XOR2_X1 u2_u0_U37 (.B( u2_K1_20 ) , .A( u2_desIn_r_37 ) , .Z( u2_u0_X_20 ) );
  XOR2_X1 u2_u0_U38 (.B( u2_K1_1 ) , .A( u2_desIn_r_57 ) , .Z( u2_u0_X_1 ) );
  XOR2_X1 u2_u0_U39 (.B( u2_K1_19 ) , .A( u2_desIn_r_29 ) , .Z( u2_u0_X_19 ) );
  XOR2_X1 u2_u0_U4 (.B( u2_K1_6 ) , .A( u2_desIn_r_39 ) , .Z( u2_u0_X_6 ) );
  XOR2_X1 u2_u0_U40 (.B( u2_K1_18 ) , .A( u2_desIn_r_37 ) , .Z( u2_u0_X_18 ) );
  XOR2_X1 u2_u0_U41 (.B( u2_K1_17 ) , .A( u2_desIn_r_29 ) , .Z( u2_u0_X_17 ) );
  XOR2_X1 u2_u0_U42 (.B( u2_K1_16 ) , .A( u2_desIn_r_21 ) , .Z( u2_u0_X_16 ) );
  XOR2_X1 u2_u0_U43 (.B( u2_K1_15 ) , .A( u2_desIn_r_13 ) , .Z( u2_u0_X_15 ) );
  XOR2_X1 u2_u0_U44 (.B( u2_K1_14 ) , .A( u2_desIn_r_5 ) , .Z( u2_u0_X_14 ) );
  XOR2_X1 u2_u0_U45 (.B( u2_K1_13 ) , .A( u2_desIn_r_63 ) , .Z( u2_u0_X_13 ) );
  XOR2_X1 u2_u0_U46 (.B( u2_K1_12 ) , .A( u2_desIn_r_5 ) , .Z( u2_u0_X_12 ) );
  XOR2_X1 u2_u0_U47 (.B( u2_K1_11 ) , .A( u2_desIn_r_63 ) , .Z( u2_u0_X_11 ) );
  XOR2_X1 u2_u0_U48 (.B( u2_K1_10 ) , .A( u2_desIn_r_55 ) , .Z( u2_u0_X_10 ) );
  XOR2_X1 u2_u0_U5 (.B( u2_K1_5 ) , .A( u2_desIn_r_31 ) , .Z( u2_u0_X_5 ) );
  XOR2_X1 u2_u0_U6 (.B( u2_K1_4 ) , .A( u2_desIn_r_23 ) , .Z( u2_u0_X_4 ) );
  AND3_X1 u2_u0_u0_U10 (.A2( u2_u0_u0_n112 ) , .ZN( u2_u0_u0_n127 ) , .A3( u2_u0_u0_n130 ) , .A1( u2_u0_u0_n148 ) );
  NAND2_X1 u2_u0_u0_U11 (.ZN( u2_u0_u0_n113 ) , .A1( u2_u0_u0_n139 ) , .A2( u2_u0_u0_n149 ) );
  AND2_X1 u2_u0_u0_U12 (.ZN( u2_u0_u0_n107 ) , .A1( u2_u0_u0_n130 ) , .A2( u2_u0_u0_n140 ) );
  AND2_X1 u2_u0_u0_U13 (.A2( u2_u0_u0_n129 ) , .A1( u2_u0_u0_n130 ) , .ZN( u2_u0_u0_n151 ) );
  AND2_X1 u2_u0_u0_U14 (.A1( u2_u0_u0_n108 ) , .A2( u2_u0_u0_n125 ) , .ZN( u2_u0_u0_n145 ) );
  INV_X1 u2_u0_u0_U15 (.A( u2_u0_u0_n143 ) , .ZN( u2_u0_u0_n173 ) );
  NOR2_X1 u2_u0_u0_U16 (.A2( u2_u0_u0_n136 ) , .ZN( u2_u0_u0_n147 ) , .A1( u2_u0_u0_n160 ) );
  OAI22_X1 u2_u0_u0_U17 (.B1( u2_u0_u0_n125 ) , .ZN( u2_u0_u0_n126 ) , .A1( u2_u0_u0_n138 ) , .A2( u2_u0_u0_n146 ) , .B2( u2_u0_u0_n147 ) );
  OAI22_X1 u2_u0_u0_U18 (.B1( u2_u0_u0_n131 ) , .A1( u2_u0_u0_n144 ) , .B2( u2_u0_u0_n147 ) , .A2( u2_u0_u0_n90 ) , .ZN( u2_u0_u0_n91 ) );
  AND3_X1 u2_u0_u0_U19 (.A3( u2_u0_u0_n121 ) , .A2( u2_u0_u0_n125 ) , .A1( u2_u0_u0_n148 ) , .ZN( u2_u0_u0_n90 ) );
  NOR2_X1 u2_u0_u0_U20 (.A1( u2_u0_u0_n163 ) , .A2( u2_u0_u0_n164 ) , .ZN( u2_u0_u0_n95 ) );
  AOI22_X1 u2_u0_u0_U21 (.B2( u2_u0_u0_n109 ) , .A2( u2_u0_u0_n110 ) , .ZN( u2_u0_u0_n111 ) , .B1( u2_u0_u0_n118 ) , .A1( u2_u0_u0_n160 ) );
  NAND2_X1 u2_u0_u0_U22 (.A1( u2_u0_u0_n100 ) , .A2( u2_u0_u0_n103 ) , .ZN( u2_u0_u0_n125 ) );
  NAND2_X1 u2_u0_u0_U23 (.A1( u2_u0_u0_n101 ) , .A2( u2_u0_u0_n102 ) , .ZN( u2_u0_u0_n150 ) );
  INV_X1 u2_u0_u0_U24 (.A( u2_u0_u0_n136 ) , .ZN( u2_u0_u0_n161 ) );
  INV_X1 u2_u0_u0_U25 (.A( u2_u0_u0_n118 ) , .ZN( u2_u0_u0_n158 ) );
  AOI21_X1 u2_u0_u0_U26 (.B1( u2_u0_u0_n127 ) , .B2( u2_u0_u0_n129 ) , .A( u2_u0_u0_n138 ) , .ZN( u2_u0_u0_n96 ) );
  AOI21_X1 u2_u0_u0_U27 (.ZN( u2_u0_u0_n104 ) , .B1( u2_u0_u0_n107 ) , .B2( u2_u0_u0_n141 ) , .A( u2_u0_u0_n144 ) );
  NAND2_X1 u2_u0_u0_U28 (.A2( u2_u0_u0_n100 ) , .A1( u2_u0_u0_n101 ) , .ZN( u2_u0_u0_n139 ) );
  NAND2_X1 u2_u0_u0_U29 (.A2( u2_u0_u0_n100 ) , .ZN( u2_u0_u0_n131 ) , .A1( u2_u0_u0_n92 ) );
  INV_X1 u2_u0_u0_U3 (.A( u2_u0_u0_n113 ) , .ZN( u2_u0_u0_n166 ) );
  NAND2_X1 u2_u0_u0_U30 (.A2( u2_u0_u0_n102 ) , .ZN( u2_u0_u0_n114 ) , .A1( u2_u0_u0_n92 ) );
  NOR2_X1 u2_u0_u0_U31 (.A1( u2_u0_u0_n120 ) , .ZN( u2_u0_u0_n143 ) , .A2( u2_u0_u0_n167 ) );
  OAI221_X1 u2_u0_u0_U32 (.C1( u2_u0_u0_n112 ) , .ZN( u2_u0_u0_n120 ) , .B1( u2_u0_u0_n138 ) , .B2( u2_u0_u0_n141 ) , .C2( u2_u0_u0_n147 ) , .A( u2_u0_u0_n172 ) );
  AOI211_X1 u2_u0_u0_U33 (.B( u2_u0_u0_n115 ) , .A( u2_u0_u0_n116 ) , .C2( u2_u0_u0_n117 ) , .C1( u2_u0_u0_n118 ) , .ZN( u2_u0_u0_n119 ) );
  INV_X1 u2_u0_u0_U34 (.A( u2_u0_u0_n138 ) , .ZN( u2_u0_u0_n160 ) );
  NAND2_X1 u2_u0_u0_U35 (.A2( u2_u0_u0_n102 ) , .A1( u2_u0_u0_n103 ) , .ZN( u2_u0_u0_n149 ) );
  NAND2_X1 u2_u0_u0_U36 (.A2( u2_u0_u0_n101 ) , .ZN( u2_u0_u0_n121 ) , .A1( u2_u0_u0_n93 ) );
  NAND2_X1 u2_u0_u0_U37 (.ZN( u2_u0_u0_n112 ) , .A2( u2_u0_u0_n92 ) , .A1( u2_u0_u0_n93 ) );
  INV_X1 u2_u0_u0_U38 (.ZN( u2_u0_u0_n172 ) , .A( u2_u0_u0_n88 ) );
  OAI222_X1 u2_u0_u0_U39 (.C1( u2_u0_u0_n108 ) , .A1( u2_u0_u0_n125 ) , .B2( u2_u0_u0_n128 ) , .B1( u2_u0_u0_n144 ) , .A2( u2_u0_u0_n158 ) , .C2( u2_u0_u0_n161 ) , .ZN( u2_u0_u0_n88 ) );
  AOI21_X1 u2_u0_u0_U4 (.B1( u2_u0_u0_n114 ) , .ZN( u2_u0_u0_n115 ) , .B2( u2_u0_u0_n129 ) , .A( u2_u0_u0_n161 ) );
  AOI21_X1 u2_u0_u0_U40 (.B1( u2_u0_u0_n103 ) , .ZN( u2_u0_u0_n132 ) , .A( u2_u0_u0_n165 ) , .B2( u2_u0_u0_n93 ) );
  OR3_X1 u2_u0_u0_U41 (.A3( u2_u0_u0_n152 ) , .A2( u2_u0_u0_n153 ) , .A1( u2_u0_u0_n154 ) , .ZN( u2_u0_u0_n155 ) );
  AOI21_X1 u2_u0_u0_U42 (.B2( u2_u0_u0_n150 ) , .B1( u2_u0_u0_n151 ) , .ZN( u2_u0_u0_n152 ) , .A( u2_u0_u0_n158 ) );
  AOI21_X1 u2_u0_u0_U43 (.A( u2_u0_u0_n144 ) , .B2( u2_u0_u0_n145 ) , .B1( u2_u0_u0_n146 ) , .ZN( u2_u0_u0_n154 ) );
  AOI21_X1 u2_u0_u0_U44 (.A( u2_u0_u0_n147 ) , .B2( u2_u0_u0_n148 ) , .B1( u2_u0_u0_n149 ) , .ZN( u2_u0_u0_n153 ) );
  INV_X1 u2_u0_u0_U45 (.ZN( u2_u0_u0_n171 ) , .A( u2_u0_u0_n99 ) );
  OAI211_X1 u2_u0_u0_U46 (.C2( u2_u0_u0_n140 ) , .C1( u2_u0_u0_n161 ) , .A( u2_u0_u0_n169 ) , .B( u2_u0_u0_n98 ) , .ZN( u2_u0_u0_n99 ) );
  INV_X1 u2_u0_u0_U47 (.ZN( u2_u0_u0_n169 ) , .A( u2_u0_u0_n91 ) );
  AOI211_X1 u2_u0_u0_U48 (.C1( u2_u0_u0_n118 ) , .A( u2_u0_u0_n123 ) , .B( u2_u0_u0_n96 ) , .C2( u2_u0_u0_n97 ) , .ZN( u2_u0_u0_n98 ) );
  NOR2_X1 u2_u0_u0_U49 (.A2( u2_u0_X_4 ) , .A1( u2_u0_X_5 ) , .ZN( u2_u0_u0_n118 ) );
  NOR2_X1 u2_u0_u0_U5 (.A1( u2_u0_u0_n108 ) , .ZN( u2_u0_u0_n123 ) , .A2( u2_u0_u0_n158 ) );
  NOR2_X1 u2_u0_u0_U50 (.A2( u2_u0_X_2 ) , .ZN( u2_u0_u0_n103 ) , .A1( u2_u0_u0_n164 ) );
  NAND2_X1 u2_u0_u0_U51 (.A2( u2_u0_X_4 ) , .A1( u2_u0_X_5 ) , .ZN( u2_u0_u0_n144 ) );
  NOR2_X1 u2_u0_u0_U52 (.A2( u2_u0_X_5 ) , .ZN( u2_u0_u0_n136 ) , .A1( u2_u0_u0_n159 ) );
  NAND2_X1 u2_u0_u0_U53 (.A1( u2_u0_X_5 ) , .ZN( u2_u0_u0_n138 ) , .A2( u2_u0_u0_n159 ) );
  AND2_X1 u2_u0_u0_U54 (.A2( u2_u0_X_3 ) , .A1( u2_u0_X_6 ) , .ZN( u2_u0_u0_n102 ) );
  INV_X1 u2_u0_u0_U55 (.A( u2_u0_X_4 ) , .ZN( u2_u0_u0_n159 ) );
  INV_X1 u2_u0_u0_U56 (.A( u2_u0_X_2 ) , .ZN( u2_u0_u0_n163 ) );
  INV_X1 u2_u0_u0_U57 (.A( u2_u0_X_3 ) , .ZN( u2_u0_u0_n162 ) );
  INV_X1 u2_u0_u0_U58 (.A( u2_u0_u0_n126 ) , .ZN( u2_u0_u0_n168 ) );
  AOI211_X1 u2_u0_u0_U59 (.B( u2_u0_u0_n133 ) , .A( u2_u0_u0_n134 ) , .C2( u2_u0_u0_n135 ) , .C1( u2_u0_u0_n136 ) , .ZN( u2_u0_u0_n137 ) );
  AOI21_X1 u2_u0_u0_U6 (.B2( u2_u0_u0_n131 ) , .ZN( u2_u0_u0_n134 ) , .B1( u2_u0_u0_n151 ) , .A( u2_u0_u0_n158 ) );
  OR4_X1 u2_u0_u0_U60 (.ZN( u2_out0_17 ) , .A4( u2_u0_u0_n122 ) , .A2( u2_u0_u0_n123 ) , .A1( u2_u0_u0_n124 ) , .A3( u2_u0_u0_n170 ) );
  AOI21_X1 u2_u0_u0_U61 (.B2( u2_u0_u0_n107 ) , .ZN( u2_u0_u0_n124 ) , .B1( u2_u0_u0_n128 ) , .A( u2_u0_u0_n161 ) );
  INV_X1 u2_u0_u0_U62 (.A( u2_u0_u0_n111 ) , .ZN( u2_u0_u0_n170 ) );
  OR4_X1 u2_u0_u0_U63 (.ZN( u2_out0_31 ) , .A4( u2_u0_u0_n155 ) , .A2( u2_u0_u0_n156 ) , .A1( u2_u0_u0_n157 ) , .A3( u2_u0_u0_n173 ) );
  AOI21_X1 u2_u0_u0_U64 (.A( u2_u0_u0_n138 ) , .B2( u2_u0_u0_n139 ) , .B1( u2_u0_u0_n140 ) , .ZN( u2_u0_u0_n157 ) );
  INV_X1 u2_u0_u0_U65 (.ZN( u2_u0_u0_n174 ) , .A( u2_u0_u0_n89 ) );
  AOI211_X1 u2_u0_u0_U66 (.B( u2_u0_u0_n104 ) , .A( u2_u0_u0_n105 ) , .ZN( u2_u0_u0_n106 ) , .C2( u2_u0_u0_n113 ) , .C1( u2_u0_u0_n160 ) );
  AOI21_X1 u2_u0_u0_U67 (.B2( u2_u0_u0_n141 ) , .B1( u2_u0_u0_n142 ) , .ZN( u2_u0_u0_n156 ) , .A( u2_u0_u0_n161 ) );
  AOI21_X1 u2_u0_u0_U68 (.ZN( u2_u0_u0_n116 ) , .B2( u2_u0_u0_n142 ) , .A( u2_u0_u0_n144 ) , .B1( u2_u0_u0_n166 ) );
  NAND2_X1 u2_u0_u0_U69 (.ZN( u2_u0_u0_n148 ) , .A1( u2_u0_u0_n93 ) , .A2( u2_u0_u0_n95 ) );
  OAI21_X1 u2_u0_u0_U7 (.B1( u2_u0_u0_n150 ) , .B2( u2_u0_u0_n158 ) , .A( u2_u0_u0_n172 ) , .ZN( u2_u0_u0_n89 ) );
  NAND2_X1 u2_u0_u0_U70 (.A1( u2_u0_u0_n100 ) , .ZN( u2_u0_u0_n129 ) , .A2( u2_u0_u0_n95 ) );
  NAND2_X1 u2_u0_u0_U71 (.A1( u2_u0_u0_n102 ) , .ZN( u2_u0_u0_n128 ) , .A2( u2_u0_u0_n95 ) );
  INV_X1 u2_u0_u0_U72 (.A( u2_u0_u0_n142 ) , .ZN( u2_u0_u0_n165 ) );
  NOR2_X1 u2_u0_u0_U73 (.A2( u2_u0_X_1 ) , .A1( u2_u0_X_2 ) , .ZN( u2_u0_u0_n92 ) );
  NOR2_X1 u2_u0_u0_U74 (.A2( u2_u0_X_1 ) , .ZN( u2_u0_u0_n101 ) , .A1( u2_u0_u0_n163 ) );
  INV_X1 u2_u0_u0_U75 (.A( u2_u0_X_1 ) , .ZN( u2_u0_u0_n164 ) );
  AND2_X1 u2_u0_u0_U76 (.A1( u2_u0_X_6 ) , .A2( u2_u0_u0_n162 ) , .ZN( u2_u0_u0_n93 ) );
  NOR2_X1 u2_u0_u0_U77 (.A2( u2_u0_X_3 ) , .A1( u2_u0_X_6 ) , .ZN( u2_u0_u0_n94 ) );
  NOR2_X1 u2_u0_u0_U78 (.A2( u2_u0_X_6 ) , .ZN( u2_u0_u0_n100 ) , .A1( u2_u0_u0_n162 ) );
  OAI221_X1 u2_u0_u0_U79 (.C1( u2_u0_u0_n121 ) , .ZN( u2_u0_u0_n122 ) , .B2( u2_u0_u0_n127 ) , .A( u2_u0_u0_n143 ) , .B1( u2_u0_u0_n144 ) , .C2( u2_u0_u0_n147 ) );
  AND2_X1 u2_u0_u0_U8 (.A1( u2_u0_u0_n114 ) , .A2( u2_u0_u0_n121 ) , .ZN( u2_u0_u0_n146 ) );
  AOI21_X1 u2_u0_u0_U80 (.B1( u2_u0_u0_n132 ) , .ZN( u2_u0_u0_n133 ) , .A( u2_u0_u0_n144 ) , .B2( u2_u0_u0_n166 ) );
  OAI22_X1 u2_u0_u0_U81 (.ZN( u2_u0_u0_n105 ) , .A2( u2_u0_u0_n132 ) , .B1( u2_u0_u0_n146 ) , .A1( u2_u0_u0_n147 ) , .B2( u2_u0_u0_n161 ) );
  NAND2_X1 u2_u0_u0_U82 (.ZN( u2_u0_u0_n110 ) , .A2( u2_u0_u0_n132 ) , .A1( u2_u0_u0_n145 ) );
  INV_X1 u2_u0_u0_U83 (.A( u2_u0_u0_n119 ) , .ZN( u2_u0_u0_n167 ) );
  NAND2_X1 u2_u0_u0_U84 (.A2( u2_u0_u0_n103 ) , .ZN( u2_u0_u0_n140 ) , .A1( u2_u0_u0_n94 ) );
  NAND2_X1 u2_u0_u0_U85 (.A1( u2_u0_u0_n101 ) , .ZN( u2_u0_u0_n130 ) , .A2( u2_u0_u0_n94 ) );
  NAND2_X1 u2_u0_u0_U86 (.ZN( u2_u0_u0_n108 ) , .A1( u2_u0_u0_n92 ) , .A2( u2_u0_u0_n94 ) );
  NAND2_X1 u2_u0_u0_U87 (.ZN( u2_u0_u0_n142 ) , .A1( u2_u0_u0_n94 ) , .A2( u2_u0_u0_n95 ) );
  NAND3_X1 u2_u0_u0_U88 (.ZN( u2_out0_23 ) , .A3( u2_u0_u0_n137 ) , .A1( u2_u0_u0_n168 ) , .A2( u2_u0_u0_n171 ) );
  NAND3_X1 u2_u0_u0_U89 (.A3( u2_u0_u0_n127 ) , .A2( u2_u0_u0_n128 ) , .ZN( u2_u0_u0_n135 ) , .A1( u2_u0_u0_n150 ) );
  AND2_X1 u2_u0_u0_U9 (.A1( u2_u0_u0_n131 ) , .ZN( u2_u0_u0_n141 ) , .A2( u2_u0_u0_n150 ) );
  NAND3_X1 u2_u0_u0_U90 (.ZN( u2_u0_u0_n117 ) , .A3( u2_u0_u0_n132 ) , .A2( u2_u0_u0_n139 ) , .A1( u2_u0_u0_n148 ) );
  NAND3_X1 u2_u0_u0_U91 (.ZN( u2_u0_u0_n109 ) , .A2( u2_u0_u0_n114 ) , .A3( u2_u0_u0_n140 ) , .A1( u2_u0_u0_n149 ) );
  NAND3_X1 u2_u0_u0_U92 (.ZN( u2_out0_9 ) , .A3( u2_u0_u0_n106 ) , .A2( u2_u0_u0_n171 ) , .A1( u2_u0_u0_n174 ) );
  NAND3_X1 u2_u0_u0_U93 (.A2( u2_u0_u0_n128 ) , .A1( u2_u0_u0_n132 ) , .A3( u2_u0_u0_n146 ) , .ZN( u2_u0_u0_n97 ) );
  AOI21_X1 u2_u0_u1_U10 (.B2( u2_u0_u1_n155 ) , .B1( u2_u0_u1_n156 ) , .ZN( u2_u0_u1_n157 ) , .A( u2_u0_u1_n174 ) );
  NAND3_X1 u2_u0_u1_U100 (.ZN( u2_u0_u1_n113 ) , .A1( u2_u0_u1_n120 ) , .A3( u2_u0_u1_n133 ) , .A2( u2_u0_u1_n155 ) );
  NAND2_X1 u2_u0_u1_U11 (.ZN( u2_u0_u1_n140 ) , .A2( u2_u0_u1_n150 ) , .A1( u2_u0_u1_n155 ) );
  NAND2_X1 u2_u0_u1_U12 (.A1( u2_u0_u1_n131 ) , .ZN( u2_u0_u1_n147 ) , .A2( u2_u0_u1_n153 ) );
  AOI22_X1 u2_u0_u1_U13 (.B2( u2_u0_u1_n136 ) , .A2( u2_u0_u1_n137 ) , .ZN( u2_u0_u1_n143 ) , .A1( u2_u0_u1_n171 ) , .B1( u2_u0_u1_n173 ) );
  INV_X1 u2_u0_u1_U14 (.A( u2_u0_u1_n147 ) , .ZN( u2_u0_u1_n181 ) );
  INV_X1 u2_u0_u1_U15 (.A( u2_u0_u1_n139 ) , .ZN( u2_u0_u1_n174 ) );
  OR4_X1 u2_u0_u1_U16 (.A4( u2_u0_u1_n106 ) , .A3( u2_u0_u1_n107 ) , .ZN( u2_u0_u1_n108 ) , .A1( u2_u0_u1_n117 ) , .A2( u2_u0_u1_n184 ) );
  AOI21_X1 u2_u0_u1_U17 (.ZN( u2_u0_u1_n106 ) , .A( u2_u0_u1_n112 ) , .B1( u2_u0_u1_n154 ) , .B2( u2_u0_u1_n156 ) );
  AOI21_X1 u2_u0_u1_U18 (.ZN( u2_u0_u1_n107 ) , .B1( u2_u0_u1_n134 ) , .B2( u2_u0_u1_n149 ) , .A( u2_u0_u1_n174 ) );
  INV_X1 u2_u0_u1_U19 (.A( u2_u0_u1_n101 ) , .ZN( u2_u0_u1_n184 ) );
  INV_X1 u2_u0_u1_U20 (.A( u2_u0_u1_n112 ) , .ZN( u2_u0_u1_n171 ) );
  NAND2_X1 u2_u0_u1_U21 (.ZN( u2_u0_u1_n141 ) , .A1( u2_u0_u1_n153 ) , .A2( u2_u0_u1_n156 ) );
  AND2_X1 u2_u0_u1_U22 (.A1( u2_u0_u1_n123 ) , .ZN( u2_u0_u1_n134 ) , .A2( u2_u0_u1_n161 ) );
  NAND2_X1 u2_u0_u1_U23 (.A2( u2_u0_u1_n115 ) , .A1( u2_u0_u1_n116 ) , .ZN( u2_u0_u1_n148 ) );
  NAND2_X1 u2_u0_u1_U24 (.A2( u2_u0_u1_n133 ) , .A1( u2_u0_u1_n135 ) , .ZN( u2_u0_u1_n159 ) );
  NAND2_X1 u2_u0_u1_U25 (.A2( u2_u0_u1_n115 ) , .A1( u2_u0_u1_n120 ) , .ZN( u2_u0_u1_n132 ) );
  INV_X1 u2_u0_u1_U26 (.A( u2_u0_u1_n154 ) , .ZN( u2_u0_u1_n178 ) );
  INV_X1 u2_u0_u1_U27 (.A( u2_u0_u1_n151 ) , .ZN( u2_u0_u1_n183 ) );
  AND2_X1 u2_u0_u1_U28 (.A1( u2_u0_u1_n129 ) , .A2( u2_u0_u1_n133 ) , .ZN( u2_u0_u1_n149 ) );
  INV_X1 u2_u0_u1_U29 (.A( u2_u0_u1_n131 ) , .ZN( u2_u0_u1_n180 ) );
  INV_X1 u2_u0_u1_U3 (.A( u2_u0_u1_n159 ) , .ZN( u2_u0_u1_n182 ) );
  AOI221_X1 u2_u0_u1_U30 (.B1( u2_u0_u1_n140 ) , .ZN( u2_u0_u1_n167 ) , .B2( u2_u0_u1_n172 ) , .C2( u2_u0_u1_n175 ) , .C1( u2_u0_u1_n178 ) , .A( u2_u0_u1_n188 ) );
  INV_X1 u2_u0_u1_U31 (.ZN( u2_u0_u1_n188 ) , .A( u2_u0_u1_n97 ) );
  AOI211_X1 u2_u0_u1_U32 (.A( u2_u0_u1_n118 ) , .C1( u2_u0_u1_n132 ) , .C2( u2_u0_u1_n139 ) , .B( u2_u0_u1_n96 ) , .ZN( u2_u0_u1_n97 ) );
  AOI21_X1 u2_u0_u1_U33 (.B2( u2_u0_u1_n121 ) , .B1( u2_u0_u1_n135 ) , .A( u2_u0_u1_n152 ) , .ZN( u2_u0_u1_n96 ) );
  OAI221_X1 u2_u0_u1_U34 (.A( u2_u0_u1_n119 ) , .C2( u2_u0_u1_n129 ) , .ZN( u2_u0_u1_n138 ) , .B2( u2_u0_u1_n152 ) , .C1( u2_u0_u1_n174 ) , .B1( u2_u0_u1_n187 ) );
  INV_X1 u2_u0_u1_U35 (.A( u2_u0_u1_n148 ) , .ZN( u2_u0_u1_n187 ) );
  AOI211_X1 u2_u0_u1_U36 (.B( u2_u0_u1_n117 ) , .A( u2_u0_u1_n118 ) , .ZN( u2_u0_u1_n119 ) , .C2( u2_u0_u1_n146 ) , .C1( u2_u0_u1_n159 ) );
  NOR2_X1 u2_u0_u1_U37 (.A1( u2_u0_u1_n168 ) , .A2( u2_u0_u1_n176 ) , .ZN( u2_u0_u1_n98 ) );
  AOI211_X1 u2_u0_u1_U38 (.B( u2_u0_u1_n162 ) , .A( u2_u0_u1_n163 ) , .C2( u2_u0_u1_n164 ) , .ZN( u2_u0_u1_n165 ) , .C1( u2_u0_u1_n171 ) );
  AOI21_X1 u2_u0_u1_U39 (.A( u2_u0_u1_n160 ) , .B2( u2_u0_u1_n161 ) , .ZN( u2_u0_u1_n162 ) , .B1( u2_u0_u1_n182 ) );
  AOI221_X1 u2_u0_u1_U4 (.A( u2_u0_u1_n138 ) , .C2( u2_u0_u1_n139 ) , .C1( u2_u0_u1_n140 ) , .B2( u2_u0_u1_n141 ) , .ZN( u2_u0_u1_n142 ) , .B1( u2_u0_u1_n175 ) );
  OR2_X1 u2_u0_u1_U40 (.A2( u2_u0_u1_n157 ) , .A1( u2_u0_u1_n158 ) , .ZN( u2_u0_u1_n163 ) );
  NAND2_X1 u2_u0_u1_U41 (.A1( u2_u0_u1_n128 ) , .ZN( u2_u0_u1_n146 ) , .A2( u2_u0_u1_n160 ) );
  NAND2_X1 u2_u0_u1_U42 (.A2( u2_u0_u1_n112 ) , .ZN( u2_u0_u1_n139 ) , .A1( u2_u0_u1_n152 ) );
  NAND2_X1 u2_u0_u1_U43 (.A1( u2_u0_u1_n105 ) , .ZN( u2_u0_u1_n156 ) , .A2( u2_u0_u1_n99 ) );
  NOR2_X1 u2_u0_u1_U44 (.ZN( u2_u0_u1_n117 ) , .A1( u2_u0_u1_n121 ) , .A2( u2_u0_u1_n160 ) );
  AOI21_X1 u2_u0_u1_U45 (.A( u2_u0_u1_n128 ) , .B2( u2_u0_u1_n129 ) , .ZN( u2_u0_u1_n130 ) , .B1( u2_u0_u1_n150 ) );
  NAND2_X1 u2_u0_u1_U46 (.ZN( u2_u0_u1_n112 ) , .A1( u2_u0_u1_n169 ) , .A2( u2_u0_u1_n170 ) );
  NAND2_X1 u2_u0_u1_U47 (.ZN( u2_u0_u1_n129 ) , .A2( u2_u0_u1_n95 ) , .A1( u2_u0_u1_n98 ) );
  NAND2_X1 u2_u0_u1_U48 (.A1( u2_u0_u1_n102 ) , .ZN( u2_u0_u1_n154 ) , .A2( u2_u0_u1_n99 ) );
  NAND2_X1 u2_u0_u1_U49 (.A2( u2_u0_u1_n100 ) , .ZN( u2_u0_u1_n135 ) , .A1( u2_u0_u1_n99 ) );
  AOI211_X1 u2_u0_u1_U5 (.ZN( u2_u0_u1_n124 ) , .A( u2_u0_u1_n138 ) , .C2( u2_u0_u1_n139 ) , .B( u2_u0_u1_n145 ) , .C1( u2_u0_u1_n147 ) );
  AOI21_X1 u2_u0_u1_U50 (.A( u2_u0_u1_n152 ) , .B2( u2_u0_u1_n153 ) , .B1( u2_u0_u1_n154 ) , .ZN( u2_u0_u1_n158 ) );
  INV_X1 u2_u0_u1_U51 (.A( u2_u0_u1_n160 ) , .ZN( u2_u0_u1_n175 ) );
  NAND2_X1 u2_u0_u1_U52 (.A1( u2_u0_u1_n100 ) , .ZN( u2_u0_u1_n116 ) , .A2( u2_u0_u1_n95 ) );
  NAND2_X1 u2_u0_u1_U53 (.A1( u2_u0_u1_n102 ) , .ZN( u2_u0_u1_n131 ) , .A2( u2_u0_u1_n95 ) );
  NAND2_X1 u2_u0_u1_U54 (.A2( u2_u0_u1_n104 ) , .ZN( u2_u0_u1_n121 ) , .A1( u2_u0_u1_n98 ) );
  NAND2_X1 u2_u0_u1_U55 (.A1( u2_u0_u1_n103 ) , .ZN( u2_u0_u1_n153 ) , .A2( u2_u0_u1_n98 ) );
  NAND2_X1 u2_u0_u1_U56 (.A2( u2_u0_u1_n104 ) , .A1( u2_u0_u1_n105 ) , .ZN( u2_u0_u1_n133 ) );
  NAND2_X1 u2_u0_u1_U57 (.ZN( u2_u0_u1_n150 ) , .A2( u2_u0_u1_n98 ) , .A1( u2_u0_u1_n99 ) );
  NAND2_X1 u2_u0_u1_U58 (.A1( u2_u0_u1_n105 ) , .ZN( u2_u0_u1_n155 ) , .A2( u2_u0_u1_n95 ) );
  OAI21_X1 u2_u0_u1_U59 (.ZN( u2_u0_u1_n109 ) , .B1( u2_u0_u1_n129 ) , .B2( u2_u0_u1_n160 ) , .A( u2_u0_u1_n167 ) );
  AOI22_X1 u2_u0_u1_U6 (.B2( u2_u0_u1_n113 ) , .A2( u2_u0_u1_n114 ) , .ZN( u2_u0_u1_n125 ) , .A1( u2_u0_u1_n171 ) , .B1( u2_u0_u1_n173 ) );
  NAND2_X1 u2_u0_u1_U60 (.A2( u2_u0_u1_n100 ) , .A1( u2_u0_u1_n103 ) , .ZN( u2_u0_u1_n120 ) );
  NAND2_X1 u2_u0_u1_U61 (.A1( u2_u0_u1_n102 ) , .A2( u2_u0_u1_n104 ) , .ZN( u2_u0_u1_n115 ) );
  NAND2_X1 u2_u0_u1_U62 (.A2( u2_u0_u1_n100 ) , .A1( u2_u0_u1_n104 ) , .ZN( u2_u0_u1_n151 ) );
  NAND2_X1 u2_u0_u1_U63 (.A2( u2_u0_u1_n103 ) , .A1( u2_u0_u1_n105 ) , .ZN( u2_u0_u1_n161 ) );
  INV_X1 u2_u0_u1_U64 (.A( u2_u0_u1_n152 ) , .ZN( u2_u0_u1_n173 ) );
  INV_X1 u2_u0_u1_U65 (.A( u2_u0_u1_n128 ) , .ZN( u2_u0_u1_n172 ) );
  NAND2_X1 u2_u0_u1_U66 (.A2( u2_u0_u1_n102 ) , .A1( u2_u0_u1_n103 ) , .ZN( u2_u0_u1_n123 ) );
  OAI21_X1 u2_u0_u1_U67 (.B2( u2_u0_u1_n123 ) , .ZN( u2_u0_u1_n145 ) , .B1( u2_u0_u1_n160 ) , .A( u2_u0_u1_n185 ) );
  INV_X1 u2_u0_u1_U68 (.A( u2_u0_u1_n122 ) , .ZN( u2_u0_u1_n185 ) );
  AOI21_X1 u2_u0_u1_U69 (.B2( u2_u0_u1_n120 ) , .B1( u2_u0_u1_n121 ) , .ZN( u2_u0_u1_n122 ) , .A( u2_u0_u1_n128 ) );
  NAND2_X1 u2_u0_u1_U7 (.ZN( u2_u0_u1_n114 ) , .A1( u2_u0_u1_n134 ) , .A2( u2_u0_u1_n156 ) );
  NOR2_X1 u2_u0_u1_U70 (.A2( u2_u0_X_7 ) , .A1( u2_u0_X_8 ) , .ZN( u2_u0_u1_n95 ) );
  NOR2_X1 u2_u0_u1_U71 (.A1( u2_u0_X_12 ) , .A2( u2_u0_X_9 ) , .ZN( u2_u0_u1_n100 ) );
  NOR2_X1 u2_u0_u1_U72 (.A2( u2_u0_X_8 ) , .A1( u2_u0_u1_n177 ) , .ZN( u2_u0_u1_n99 ) );
  NOR2_X1 u2_u0_u1_U73 (.A2( u2_u0_X_12 ) , .ZN( u2_u0_u1_n102 ) , .A1( u2_u0_u1_n176 ) );
  NOR2_X1 u2_u0_u1_U74 (.A2( u2_u0_X_9 ) , .ZN( u2_u0_u1_n105 ) , .A1( u2_u0_u1_n168 ) );
  NAND2_X1 u2_u0_u1_U75 (.A1( u2_u0_X_10 ) , .ZN( u2_u0_u1_n160 ) , .A2( u2_u0_u1_n169 ) );
  NAND2_X1 u2_u0_u1_U76 (.A2( u2_u0_X_10 ) , .A1( u2_u0_X_11 ) , .ZN( u2_u0_u1_n152 ) );
  NAND2_X1 u2_u0_u1_U77 (.A1( u2_u0_X_11 ) , .ZN( u2_u0_u1_n128 ) , .A2( u2_u0_u1_n170 ) );
  AND2_X1 u2_u0_u1_U78 (.A2( u2_u0_X_7 ) , .A1( u2_u0_X_8 ) , .ZN( u2_u0_u1_n104 ) );
  AND2_X1 u2_u0_u1_U79 (.A1( u2_u0_X_8 ) , .ZN( u2_u0_u1_n103 ) , .A2( u2_u0_u1_n177 ) );
  NOR2_X1 u2_u0_u1_U8 (.A1( u2_u0_u1_n112 ) , .A2( u2_u0_u1_n116 ) , .ZN( u2_u0_u1_n118 ) );
  INV_X1 u2_u0_u1_U80 (.A( u2_u0_X_10 ) , .ZN( u2_u0_u1_n170 ) );
  INV_X1 u2_u0_u1_U81 (.A( u2_u0_X_9 ) , .ZN( u2_u0_u1_n176 ) );
  INV_X1 u2_u0_u1_U82 (.A( u2_u0_X_11 ) , .ZN( u2_u0_u1_n169 ) );
  INV_X1 u2_u0_u1_U83 (.A( u2_u0_X_12 ) , .ZN( u2_u0_u1_n168 ) );
  INV_X1 u2_u0_u1_U84 (.A( u2_u0_X_7 ) , .ZN( u2_u0_u1_n177 ) );
  NAND4_X1 u2_u0_u1_U85 (.ZN( u2_out0_28 ) , .A4( u2_u0_u1_n124 ) , .A3( u2_u0_u1_n125 ) , .A2( u2_u0_u1_n126 ) , .A1( u2_u0_u1_n127 ) );
  OAI21_X1 u2_u0_u1_U86 (.ZN( u2_u0_u1_n127 ) , .B2( u2_u0_u1_n139 ) , .B1( u2_u0_u1_n175 ) , .A( u2_u0_u1_n183 ) );
  OAI21_X1 u2_u0_u1_U87 (.ZN( u2_u0_u1_n126 ) , .B2( u2_u0_u1_n140 ) , .A( u2_u0_u1_n146 ) , .B1( u2_u0_u1_n178 ) );
  NAND4_X1 u2_u0_u1_U88 (.ZN( u2_out0_18 ) , .A4( u2_u0_u1_n165 ) , .A3( u2_u0_u1_n166 ) , .A1( u2_u0_u1_n167 ) , .A2( u2_u0_u1_n186 ) );
  AOI22_X1 u2_u0_u1_U89 (.B2( u2_u0_u1_n146 ) , .B1( u2_u0_u1_n147 ) , .A2( u2_u0_u1_n148 ) , .ZN( u2_u0_u1_n166 ) , .A1( u2_u0_u1_n172 ) );
  OAI21_X1 u2_u0_u1_U9 (.ZN( u2_u0_u1_n101 ) , .B1( u2_u0_u1_n141 ) , .A( u2_u0_u1_n146 ) , .B2( u2_u0_u1_n183 ) );
  INV_X1 u2_u0_u1_U90 (.A( u2_u0_u1_n145 ) , .ZN( u2_u0_u1_n186 ) );
  NAND4_X1 u2_u0_u1_U91 (.ZN( u2_out0_2 ) , .A4( u2_u0_u1_n142 ) , .A3( u2_u0_u1_n143 ) , .A2( u2_u0_u1_n144 ) , .A1( u2_u0_u1_n179 ) );
  OAI21_X1 u2_u0_u1_U92 (.B2( u2_u0_u1_n132 ) , .ZN( u2_u0_u1_n144 ) , .A( u2_u0_u1_n146 ) , .B1( u2_u0_u1_n180 ) );
  INV_X1 u2_u0_u1_U93 (.A( u2_u0_u1_n130 ) , .ZN( u2_u0_u1_n179 ) );
  OR4_X1 u2_u0_u1_U94 (.ZN( u2_out0_13 ) , .A4( u2_u0_u1_n108 ) , .A3( u2_u0_u1_n109 ) , .A2( u2_u0_u1_n110 ) , .A1( u2_u0_u1_n111 ) );
  AOI21_X1 u2_u0_u1_U95 (.ZN( u2_u0_u1_n111 ) , .A( u2_u0_u1_n128 ) , .B2( u2_u0_u1_n131 ) , .B1( u2_u0_u1_n135 ) );
  AOI21_X1 u2_u0_u1_U96 (.ZN( u2_u0_u1_n110 ) , .A( u2_u0_u1_n116 ) , .B1( u2_u0_u1_n152 ) , .B2( u2_u0_u1_n160 ) );
  NAND3_X1 u2_u0_u1_U97 (.A3( u2_u0_u1_n149 ) , .A2( u2_u0_u1_n150 ) , .A1( u2_u0_u1_n151 ) , .ZN( u2_u0_u1_n164 ) );
  NAND3_X1 u2_u0_u1_U98 (.A3( u2_u0_u1_n134 ) , .A2( u2_u0_u1_n135 ) , .ZN( u2_u0_u1_n136 ) , .A1( u2_u0_u1_n151 ) );
  NAND3_X1 u2_u0_u1_U99 (.A1( u2_u0_u1_n133 ) , .ZN( u2_u0_u1_n137 ) , .A2( u2_u0_u1_n154 ) , .A3( u2_u0_u1_n181 ) );
  OAI22_X1 u2_u0_u2_U10 (.B1( u2_u0_u2_n151 ) , .A2( u2_u0_u2_n152 ) , .A1( u2_u0_u2_n153 ) , .ZN( u2_u0_u2_n160 ) , .B2( u2_u0_u2_n168 ) );
  NAND3_X1 u2_u0_u2_U100 (.A2( u2_u0_u2_n100 ) , .A1( u2_u0_u2_n104 ) , .A3( u2_u0_u2_n138 ) , .ZN( u2_u0_u2_n98 ) );
  NOR3_X1 u2_u0_u2_U11 (.A1( u2_u0_u2_n150 ) , .ZN( u2_u0_u2_n151 ) , .A3( u2_u0_u2_n175 ) , .A2( u2_u0_u2_n188 ) );
  AOI21_X1 u2_u0_u2_U12 (.B2( u2_u0_u2_n123 ) , .ZN( u2_u0_u2_n125 ) , .A( u2_u0_u2_n171 ) , .B1( u2_u0_u2_n184 ) );
  INV_X1 u2_u0_u2_U13 (.A( u2_u0_u2_n150 ) , .ZN( u2_u0_u2_n184 ) );
  AOI21_X1 u2_u0_u2_U14 (.ZN( u2_u0_u2_n144 ) , .B2( u2_u0_u2_n155 ) , .A( u2_u0_u2_n172 ) , .B1( u2_u0_u2_n185 ) );
  AOI21_X1 u2_u0_u2_U15 (.B2( u2_u0_u2_n143 ) , .ZN( u2_u0_u2_n145 ) , .B1( u2_u0_u2_n152 ) , .A( u2_u0_u2_n171 ) );
  INV_X1 u2_u0_u2_U16 (.A( u2_u0_u2_n156 ) , .ZN( u2_u0_u2_n171 ) );
  INV_X1 u2_u0_u2_U17 (.A( u2_u0_u2_n120 ) , .ZN( u2_u0_u2_n188 ) );
  NAND2_X1 u2_u0_u2_U18 (.A2( u2_u0_u2_n122 ) , .ZN( u2_u0_u2_n150 ) , .A1( u2_u0_u2_n152 ) );
  INV_X1 u2_u0_u2_U19 (.A( u2_u0_u2_n153 ) , .ZN( u2_u0_u2_n170 ) );
  INV_X1 u2_u0_u2_U20 (.A( u2_u0_u2_n137 ) , .ZN( u2_u0_u2_n173 ) );
  NAND2_X1 u2_u0_u2_U21 (.A1( u2_u0_u2_n132 ) , .A2( u2_u0_u2_n139 ) , .ZN( u2_u0_u2_n157 ) );
  INV_X1 u2_u0_u2_U22 (.A( u2_u0_u2_n113 ) , .ZN( u2_u0_u2_n178 ) );
  INV_X1 u2_u0_u2_U23 (.A( u2_u0_u2_n139 ) , .ZN( u2_u0_u2_n175 ) );
  INV_X1 u2_u0_u2_U24 (.A( u2_u0_u2_n155 ) , .ZN( u2_u0_u2_n181 ) );
  INV_X1 u2_u0_u2_U25 (.A( u2_u0_u2_n119 ) , .ZN( u2_u0_u2_n177 ) );
  INV_X1 u2_u0_u2_U26 (.A( u2_u0_u2_n116 ) , .ZN( u2_u0_u2_n180 ) );
  INV_X1 u2_u0_u2_U27 (.A( u2_u0_u2_n131 ) , .ZN( u2_u0_u2_n179 ) );
  INV_X1 u2_u0_u2_U28 (.A( u2_u0_u2_n154 ) , .ZN( u2_u0_u2_n176 ) );
  NAND2_X1 u2_u0_u2_U29 (.A2( u2_u0_u2_n116 ) , .A1( u2_u0_u2_n117 ) , .ZN( u2_u0_u2_n118 ) );
  NOR2_X1 u2_u0_u2_U3 (.ZN( u2_u0_u2_n121 ) , .A2( u2_u0_u2_n177 ) , .A1( u2_u0_u2_n180 ) );
  INV_X1 u2_u0_u2_U30 (.A( u2_u0_u2_n132 ) , .ZN( u2_u0_u2_n182 ) );
  INV_X1 u2_u0_u2_U31 (.A( u2_u0_u2_n158 ) , .ZN( u2_u0_u2_n183 ) );
  OAI21_X1 u2_u0_u2_U32 (.A( u2_u0_u2_n156 ) , .B1( u2_u0_u2_n157 ) , .ZN( u2_u0_u2_n158 ) , .B2( u2_u0_u2_n179 ) );
  NOR2_X1 u2_u0_u2_U33 (.ZN( u2_u0_u2_n156 ) , .A1( u2_u0_u2_n166 ) , .A2( u2_u0_u2_n169 ) );
  NOR2_X1 u2_u0_u2_U34 (.A2( u2_u0_u2_n114 ) , .ZN( u2_u0_u2_n137 ) , .A1( u2_u0_u2_n140 ) );
  NOR2_X1 u2_u0_u2_U35 (.A2( u2_u0_u2_n138 ) , .ZN( u2_u0_u2_n153 ) , .A1( u2_u0_u2_n156 ) );
  AOI211_X1 u2_u0_u2_U36 (.ZN( u2_u0_u2_n130 ) , .C1( u2_u0_u2_n138 ) , .C2( u2_u0_u2_n179 ) , .B( u2_u0_u2_n96 ) , .A( u2_u0_u2_n97 ) );
  OAI22_X1 u2_u0_u2_U37 (.B1( u2_u0_u2_n133 ) , .A2( u2_u0_u2_n137 ) , .A1( u2_u0_u2_n152 ) , .B2( u2_u0_u2_n168 ) , .ZN( u2_u0_u2_n97 ) );
  OAI221_X1 u2_u0_u2_U38 (.B1( u2_u0_u2_n113 ) , .C1( u2_u0_u2_n132 ) , .A( u2_u0_u2_n149 ) , .B2( u2_u0_u2_n171 ) , .C2( u2_u0_u2_n172 ) , .ZN( u2_u0_u2_n96 ) );
  OAI221_X1 u2_u0_u2_U39 (.A( u2_u0_u2_n115 ) , .C2( u2_u0_u2_n123 ) , .B2( u2_u0_u2_n143 ) , .B1( u2_u0_u2_n153 ) , .ZN( u2_u0_u2_n163 ) , .C1( u2_u0_u2_n168 ) );
  INV_X1 u2_u0_u2_U4 (.A( u2_u0_u2_n134 ) , .ZN( u2_u0_u2_n185 ) );
  OAI21_X1 u2_u0_u2_U40 (.A( u2_u0_u2_n114 ) , .ZN( u2_u0_u2_n115 ) , .B1( u2_u0_u2_n176 ) , .B2( u2_u0_u2_n178 ) );
  OAI221_X1 u2_u0_u2_U41 (.A( u2_u0_u2_n135 ) , .B2( u2_u0_u2_n136 ) , .B1( u2_u0_u2_n137 ) , .ZN( u2_u0_u2_n162 ) , .C2( u2_u0_u2_n167 ) , .C1( u2_u0_u2_n185 ) );
  AND3_X1 u2_u0_u2_U42 (.A3( u2_u0_u2_n131 ) , .A2( u2_u0_u2_n132 ) , .A1( u2_u0_u2_n133 ) , .ZN( u2_u0_u2_n136 ) );
  AOI22_X1 u2_u0_u2_U43 (.ZN( u2_u0_u2_n135 ) , .B1( u2_u0_u2_n140 ) , .A1( u2_u0_u2_n156 ) , .B2( u2_u0_u2_n180 ) , .A2( u2_u0_u2_n188 ) );
  AOI21_X1 u2_u0_u2_U44 (.ZN( u2_u0_u2_n149 ) , .B1( u2_u0_u2_n173 ) , .B2( u2_u0_u2_n188 ) , .A( u2_u0_u2_n95 ) );
  AND3_X1 u2_u0_u2_U45 (.A2( u2_u0_u2_n100 ) , .A1( u2_u0_u2_n104 ) , .A3( u2_u0_u2_n156 ) , .ZN( u2_u0_u2_n95 ) );
  OAI21_X1 u2_u0_u2_U46 (.A( u2_u0_u2_n141 ) , .B2( u2_u0_u2_n142 ) , .ZN( u2_u0_u2_n146 ) , .B1( u2_u0_u2_n153 ) );
  OAI21_X1 u2_u0_u2_U47 (.A( u2_u0_u2_n140 ) , .ZN( u2_u0_u2_n141 ) , .B1( u2_u0_u2_n176 ) , .B2( u2_u0_u2_n177 ) );
  NOR3_X1 u2_u0_u2_U48 (.ZN( u2_u0_u2_n142 ) , .A3( u2_u0_u2_n175 ) , .A2( u2_u0_u2_n178 ) , .A1( u2_u0_u2_n181 ) );
  OAI21_X1 u2_u0_u2_U49 (.A( u2_u0_u2_n101 ) , .B2( u2_u0_u2_n121 ) , .B1( u2_u0_u2_n153 ) , .ZN( u2_u0_u2_n164 ) );
  NOR4_X1 u2_u0_u2_U5 (.A4( u2_u0_u2_n124 ) , .A3( u2_u0_u2_n125 ) , .A2( u2_u0_u2_n126 ) , .A1( u2_u0_u2_n127 ) , .ZN( u2_u0_u2_n128 ) );
  NAND2_X1 u2_u0_u2_U50 (.A2( u2_u0_u2_n100 ) , .A1( u2_u0_u2_n107 ) , .ZN( u2_u0_u2_n155 ) );
  NAND2_X1 u2_u0_u2_U51 (.A2( u2_u0_u2_n105 ) , .A1( u2_u0_u2_n108 ) , .ZN( u2_u0_u2_n143 ) );
  NAND2_X1 u2_u0_u2_U52 (.A1( u2_u0_u2_n104 ) , .A2( u2_u0_u2_n106 ) , .ZN( u2_u0_u2_n152 ) );
  NAND2_X1 u2_u0_u2_U53 (.A1( u2_u0_u2_n100 ) , .A2( u2_u0_u2_n105 ) , .ZN( u2_u0_u2_n132 ) );
  INV_X1 u2_u0_u2_U54 (.A( u2_u0_u2_n140 ) , .ZN( u2_u0_u2_n168 ) );
  INV_X1 u2_u0_u2_U55 (.A( u2_u0_u2_n138 ) , .ZN( u2_u0_u2_n167 ) );
  NAND2_X1 u2_u0_u2_U56 (.A1( u2_u0_u2_n102 ) , .A2( u2_u0_u2_n106 ) , .ZN( u2_u0_u2_n113 ) );
  NAND2_X1 u2_u0_u2_U57 (.A1( u2_u0_u2_n106 ) , .A2( u2_u0_u2_n107 ) , .ZN( u2_u0_u2_n131 ) );
  NAND2_X1 u2_u0_u2_U58 (.A1( u2_u0_u2_n103 ) , .A2( u2_u0_u2_n107 ) , .ZN( u2_u0_u2_n139 ) );
  NAND2_X1 u2_u0_u2_U59 (.A1( u2_u0_u2_n103 ) , .A2( u2_u0_u2_n105 ) , .ZN( u2_u0_u2_n133 ) );
  AOI21_X1 u2_u0_u2_U6 (.B2( u2_u0_u2_n119 ) , .ZN( u2_u0_u2_n127 ) , .A( u2_u0_u2_n137 ) , .B1( u2_u0_u2_n155 ) );
  NAND2_X1 u2_u0_u2_U60 (.A1( u2_u0_u2_n102 ) , .A2( u2_u0_u2_n103 ) , .ZN( u2_u0_u2_n154 ) );
  NAND2_X1 u2_u0_u2_U61 (.A2( u2_u0_u2_n103 ) , .A1( u2_u0_u2_n104 ) , .ZN( u2_u0_u2_n119 ) );
  NAND2_X1 u2_u0_u2_U62 (.A2( u2_u0_u2_n107 ) , .A1( u2_u0_u2_n108 ) , .ZN( u2_u0_u2_n123 ) );
  NAND2_X1 u2_u0_u2_U63 (.A1( u2_u0_u2_n104 ) , .A2( u2_u0_u2_n108 ) , .ZN( u2_u0_u2_n122 ) );
  INV_X1 u2_u0_u2_U64 (.A( u2_u0_u2_n114 ) , .ZN( u2_u0_u2_n172 ) );
  NAND2_X1 u2_u0_u2_U65 (.A2( u2_u0_u2_n100 ) , .A1( u2_u0_u2_n102 ) , .ZN( u2_u0_u2_n116 ) );
  NAND2_X1 u2_u0_u2_U66 (.A1( u2_u0_u2_n102 ) , .A2( u2_u0_u2_n108 ) , .ZN( u2_u0_u2_n120 ) );
  NAND2_X1 u2_u0_u2_U67 (.A2( u2_u0_u2_n105 ) , .A1( u2_u0_u2_n106 ) , .ZN( u2_u0_u2_n117 ) );
  INV_X1 u2_u0_u2_U68 (.ZN( u2_u0_u2_n187 ) , .A( u2_u0_u2_n99 ) );
  OAI21_X1 u2_u0_u2_U69 (.B1( u2_u0_u2_n137 ) , .B2( u2_u0_u2_n143 ) , .A( u2_u0_u2_n98 ) , .ZN( u2_u0_u2_n99 ) );
  AOI21_X1 u2_u0_u2_U7 (.ZN( u2_u0_u2_n124 ) , .B1( u2_u0_u2_n131 ) , .B2( u2_u0_u2_n143 ) , .A( u2_u0_u2_n172 ) );
  NOR2_X1 u2_u0_u2_U70 (.A2( u2_u0_X_16 ) , .ZN( u2_u0_u2_n140 ) , .A1( u2_u0_u2_n166 ) );
  NOR2_X1 u2_u0_u2_U71 (.A2( u2_u0_X_13 ) , .A1( u2_u0_X_14 ) , .ZN( u2_u0_u2_n100 ) );
  NOR2_X1 u2_u0_u2_U72 (.A2( u2_u0_X_16 ) , .A1( u2_u0_X_17 ) , .ZN( u2_u0_u2_n138 ) );
  NOR2_X1 u2_u0_u2_U73 (.A2( u2_u0_X_15 ) , .A1( u2_u0_X_18 ) , .ZN( u2_u0_u2_n104 ) );
  NOR2_X1 u2_u0_u2_U74 (.A2( u2_u0_X_14 ) , .ZN( u2_u0_u2_n103 ) , .A1( u2_u0_u2_n174 ) );
  NOR2_X1 u2_u0_u2_U75 (.A2( u2_u0_X_15 ) , .ZN( u2_u0_u2_n102 ) , .A1( u2_u0_u2_n165 ) );
  NOR2_X1 u2_u0_u2_U76 (.A2( u2_u0_X_17 ) , .ZN( u2_u0_u2_n114 ) , .A1( u2_u0_u2_n169 ) );
  AND2_X1 u2_u0_u2_U77 (.A1( u2_u0_X_15 ) , .ZN( u2_u0_u2_n105 ) , .A2( u2_u0_u2_n165 ) );
  AND2_X1 u2_u0_u2_U78 (.A2( u2_u0_X_15 ) , .A1( u2_u0_X_18 ) , .ZN( u2_u0_u2_n107 ) );
  AND2_X1 u2_u0_u2_U79 (.A1( u2_u0_X_14 ) , .ZN( u2_u0_u2_n106 ) , .A2( u2_u0_u2_n174 ) );
  AOI21_X1 u2_u0_u2_U8 (.B2( u2_u0_u2_n120 ) , .B1( u2_u0_u2_n121 ) , .ZN( u2_u0_u2_n126 ) , .A( u2_u0_u2_n167 ) );
  AND2_X1 u2_u0_u2_U80 (.A1( u2_u0_X_13 ) , .A2( u2_u0_X_14 ) , .ZN( u2_u0_u2_n108 ) );
  INV_X1 u2_u0_u2_U81 (.A( u2_u0_X_16 ) , .ZN( u2_u0_u2_n169 ) );
  INV_X1 u2_u0_u2_U82 (.A( u2_u0_X_17 ) , .ZN( u2_u0_u2_n166 ) );
  INV_X1 u2_u0_u2_U83 (.A( u2_u0_X_13 ) , .ZN( u2_u0_u2_n174 ) );
  INV_X1 u2_u0_u2_U84 (.A( u2_u0_X_18 ) , .ZN( u2_u0_u2_n165 ) );
  NAND4_X1 u2_u0_u2_U85 (.ZN( u2_out0_30 ) , .A4( u2_u0_u2_n147 ) , .A3( u2_u0_u2_n148 ) , .A2( u2_u0_u2_n149 ) , .A1( u2_u0_u2_n187 ) );
  NOR3_X1 u2_u0_u2_U86 (.A3( u2_u0_u2_n144 ) , .A2( u2_u0_u2_n145 ) , .A1( u2_u0_u2_n146 ) , .ZN( u2_u0_u2_n147 ) );
  AOI21_X1 u2_u0_u2_U87 (.B2( u2_u0_u2_n138 ) , .ZN( u2_u0_u2_n148 ) , .A( u2_u0_u2_n162 ) , .B1( u2_u0_u2_n182 ) );
  NAND4_X1 u2_u0_u2_U88 (.ZN( u2_out0_24 ) , .A4( u2_u0_u2_n111 ) , .A3( u2_u0_u2_n112 ) , .A1( u2_u0_u2_n130 ) , .A2( u2_u0_u2_n187 ) );
  AOI221_X1 u2_u0_u2_U89 (.A( u2_u0_u2_n109 ) , .B1( u2_u0_u2_n110 ) , .ZN( u2_u0_u2_n111 ) , .C1( u2_u0_u2_n134 ) , .C2( u2_u0_u2_n170 ) , .B2( u2_u0_u2_n173 ) );
  OAI22_X1 u2_u0_u2_U9 (.ZN( u2_u0_u2_n109 ) , .A2( u2_u0_u2_n113 ) , .B2( u2_u0_u2_n133 ) , .B1( u2_u0_u2_n167 ) , .A1( u2_u0_u2_n168 ) );
  AOI21_X1 u2_u0_u2_U90 (.ZN( u2_u0_u2_n112 ) , .B2( u2_u0_u2_n156 ) , .A( u2_u0_u2_n164 ) , .B1( u2_u0_u2_n181 ) );
  NAND4_X1 u2_u0_u2_U91 (.ZN( u2_out0_16 ) , .A4( u2_u0_u2_n128 ) , .A3( u2_u0_u2_n129 ) , .A1( u2_u0_u2_n130 ) , .A2( u2_u0_u2_n186 ) );
  AOI22_X1 u2_u0_u2_U92 (.A2( u2_u0_u2_n118 ) , .ZN( u2_u0_u2_n129 ) , .A1( u2_u0_u2_n140 ) , .B1( u2_u0_u2_n157 ) , .B2( u2_u0_u2_n170 ) );
  INV_X1 u2_u0_u2_U93 (.A( u2_u0_u2_n163 ) , .ZN( u2_u0_u2_n186 ) );
  OR4_X1 u2_u0_u2_U94 (.ZN( u2_out0_6 ) , .A4( u2_u0_u2_n161 ) , .A3( u2_u0_u2_n162 ) , .A2( u2_u0_u2_n163 ) , .A1( u2_u0_u2_n164 ) );
  OR3_X1 u2_u0_u2_U95 (.A2( u2_u0_u2_n159 ) , .A1( u2_u0_u2_n160 ) , .ZN( u2_u0_u2_n161 ) , .A3( u2_u0_u2_n183 ) );
  AOI21_X1 u2_u0_u2_U96 (.B2( u2_u0_u2_n154 ) , .B1( u2_u0_u2_n155 ) , .ZN( u2_u0_u2_n159 ) , .A( u2_u0_u2_n167 ) );
  NAND3_X1 u2_u0_u2_U97 (.A2( u2_u0_u2_n117 ) , .A1( u2_u0_u2_n122 ) , .A3( u2_u0_u2_n123 ) , .ZN( u2_u0_u2_n134 ) );
  NAND3_X1 u2_u0_u2_U98 (.ZN( u2_u0_u2_n110 ) , .A2( u2_u0_u2_n131 ) , .A3( u2_u0_u2_n139 ) , .A1( u2_u0_u2_n154 ) );
  NAND3_X1 u2_u0_u2_U99 (.A2( u2_u0_u2_n100 ) , .ZN( u2_u0_u2_n101 ) , .A1( u2_u0_u2_n104 ) , .A3( u2_u0_u2_n114 ) );
  OAI211_X1 u2_u0_u3_U10 (.B( u2_u0_u3_n106 ) , .ZN( u2_u0_u3_n119 ) , .C2( u2_u0_u3_n128 ) , .C1( u2_u0_u3_n167 ) , .A( u2_u0_u3_n181 ) );
  AOI221_X1 u2_u0_u3_U11 (.C1( u2_u0_u3_n105 ) , .ZN( u2_u0_u3_n106 ) , .A( u2_u0_u3_n131 ) , .B2( u2_u0_u3_n132 ) , .C2( u2_u0_u3_n133 ) , .B1( u2_u0_u3_n169 ) );
  INV_X1 u2_u0_u3_U12 (.ZN( u2_u0_u3_n181 ) , .A( u2_u0_u3_n98 ) );
  NAND2_X1 u2_u0_u3_U13 (.ZN( u2_u0_u3_n105 ) , .A2( u2_u0_u3_n130 ) , .A1( u2_u0_u3_n155 ) );
  AOI22_X1 u2_u0_u3_U14 (.B1( u2_u0_u3_n115 ) , .A2( u2_u0_u3_n116 ) , .ZN( u2_u0_u3_n123 ) , .B2( u2_u0_u3_n133 ) , .A1( u2_u0_u3_n169 ) );
  NAND2_X1 u2_u0_u3_U15 (.ZN( u2_u0_u3_n116 ) , .A2( u2_u0_u3_n151 ) , .A1( u2_u0_u3_n182 ) );
  NOR2_X1 u2_u0_u3_U16 (.ZN( u2_u0_u3_n126 ) , .A2( u2_u0_u3_n150 ) , .A1( u2_u0_u3_n164 ) );
  AOI21_X1 u2_u0_u3_U17 (.ZN( u2_u0_u3_n112 ) , .B2( u2_u0_u3_n146 ) , .B1( u2_u0_u3_n155 ) , .A( u2_u0_u3_n167 ) );
  NAND2_X1 u2_u0_u3_U18 (.A1( u2_u0_u3_n135 ) , .ZN( u2_u0_u3_n142 ) , .A2( u2_u0_u3_n164 ) );
  NAND2_X1 u2_u0_u3_U19 (.ZN( u2_u0_u3_n132 ) , .A2( u2_u0_u3_n152 ) , .A1( u2_u0_u3_n156 ) );
  INV_X1 u2_u0_u3_U20 (.A( u2_u0_u3_n133 ) , .ZN( u2_u0_u3_n165 ) );
  AND2_X1 u2_u0_u3_U21 (.A2( u2_u0_u3_n113 ) , .A1( u2_u0_u3_n114 ) , .ZN( u2_u0_u3_n151 ) );
  INV_X1 u2_u0_u3_U22 (.A( u2_u0_u3_n135 ) , .ZN( u2_u0_u3_n170 ) );
  NAND2_X1 u2_u0_u3_U23 (.A1( u2_u0_u3_n107 ) , .A2( u2_u0_u3_n108 ) , .ZN( u2_u0_u3_n140 ) );
  NAND2_X1 u2_u0_u3_U24 (.ZN( u2_u0_u3_n117 ) , .A1( u2_u0_u3_n124 ) , .A2( u2_u0_u3_n148 ) );
  INV_X1 u2_u0_u3_U25 (.A( u2_u0_u3_n128 ) , .ZN( u2_u0_u3_n176 ) );
  INV_X1 u2_u0_u3_U26 (.A( u2_u0_u3_n155 ) , .ZN( u2_u0_u3_n174 ) );
  INV_X1 u2_u0_u3_U27 (.A( u2_u0_u3_n130 ) , .ZN( u2_u0_u3_n177 ) );
  INV_X1 u2_u0_u3_U28 (.A( u2_u0_u3_n139 ) , .ZN( u2_u0_u3_n185 ) );
  NOR2_X1 u2_u0_u3_U29 (.ZN( u2_u0_u3_n135 ) , .A2( u2_u0_u3_n141 ) , .A1( u2_u0_u3_n169 ) );
  INV_X1 u2_u0_u3_U3 (.A( u2_u0_u3_n140 ) , .ZN( u2_u0_u3_n182 ) );
  OAI222_X1 u2_u0_u3_U30 (.C2( u2_u0_u3_n107 ) , .A2( u2_u0_u3_n108 ) , .B1( u2_u0_u3_n135 ) , .ZN( u2_u0_u3_n138 ) , .B2( u2_u0_u3_n146 ) , .C1( u2_u0_u3_n154 ) , .A1( u2_u0_u3_n164 ) );
  NOR4_X1 u2_u0_u3_U31 (.A4( u2_u0_u3_n157 ) , .A3( u2_u0_u3_n158 ) , .A2( u2_u0_u3_n159 ) , .A1( u2_u0_u3_n160 ) , .ZN( u2_u0_u3_n161 ) );
  AOI21_X1 u2_u0_u3_U32 (.B2( u2_u0_u3_n152 ) , .B1( u2_u0_u3_n153 ) , .ZN( u2_u0_u3_n158 ) , .A( u2_u0_u3_n164 ) );
  AOI21_X1 u2_u0_u3_U33 (.A( u2_u0_u3_n154 ) , .B2( u2_u0_u3_n155 ) , .B1( u2_u0_u3_n156 ) , .ZN( u2_u0_u3_n157 ) );
  AOI21_X1 u2_u0_u3_U34 (.A( u2_u0_u3_n149 ) , .B2( u2_u0_u3_n150 ) , .B1( u2_u0_u3_n151 ) , .ZN( u2_u0_u3_n159 ) );
  AOI211_X1 u2_u0_u3_U35 (.ZN( u2_u0_u3_n109 ) , .A( u2_u0_u3_n119 ) , .C2( u2_u0_u3_n129 ) , .B( u2_u0_u3_n138 ) , .C1( u2_u0_u3_n141 ) );
  AOI211_X1 u2_u0_u3_U36 (.B( u2_u0_u3_n119 ) , .A( u2_u0_u3_n120 ) , .C2( u2_u0_u3_n121 ) , .ZN( u2_u0_u3_n122 ) , .C1( u2_u0_u3_n179 ) );
  INV_X1 u2_u0_u3_U37 (.A( u2_u0_u3_n156 ) , .ZN( u2_u0_u3_n179 ) );
  OAI22_X1 u2_u0_u3_U38 (.B1( u2_u0_u3_n118 ) , .ZN( u2_u0_u3_n120 ) , .A1( u2_u0_u3_n135 ) , .B2( u2_u0_u3_n154 ) , .A2( u2_u0_u3_n178 ) );
  AND3_X1 u2_u0_u3_U39 (.ZN( u2_u0_u3_n118 ) , .A2( u2_u0_u3_n124 ) , .A1( u2_u0_u3_n144 ) , .A3( u2_u0_u3_n152 ) );
  INV_X1 u2_u0_u3_U4 (.A( u2_u0_u3_n129 ) , .ZN( u2_u0_u3_n183 ) );
  INV_X1 u2_u0_u3_U40 (.A( u2_u0_u3_n121 ) , .ZN( u2_u0_u3_n164 ) );
  OAI211_X1 u2_u0_u3_U41 (.B( u2_u0_u3_n127 ) , .ZN( u2_u0_u3_n139 ) , .C1( u2_u0_u3_n150 ) , .C2( u2_u0_u3_n154 ) , .A( u2_u0_u3_n184 ) );
  INV_X1 u2_u0_u3_U42 (.A( u2_u0_u3_n125 ) , .ZN( u2_u0_u3_n184 ) );
  AOI221_X1 u2_u0_u3_U43 (.A( u2_u0_u3_n126 ) , .ZN( u2_u0_u3_n127 ) , .C2( u2_u0_u3_n132 ) , .C1( u2_u0_u3_n169 ) , .B2( u2_u0_u3_n170 ) , .B1( u2_u0_u3_n174 ) );
  OAI22_X1 u2_u0_u3_U44 (.A1( u2_u0_u3_n124 ) , .ZN( u2_u0_u3_n125 ) , .B2( u2_u0_u3_n145 ) , .A2( u2_u0_u3_n165 ) , .B1( u2_u0_u3_n167 ) );
  NAND2_X1 u2_u0_u3_U45 (.A1( u2_u0_u3_n103 ) , .ZN( u2_u0_u3_n150 ) , .A2( u2_u0_u3_n99 ) );
  NAND2_X1 u2_u0_u3_U46 (.A2( u2_u0_u3_n102 ) , .ZN( u2_u0_u3_n155 ) , .A1( u2_u0_u3_n97 ) );
  NAND2_X1 u2_u0_u3_U47 (.ZN( u2_u0_u3_n133 ) , .A1( u2_u0_u3_n154 ) , .A2( u2_u0_u3_n164 ) );
  NOR2_X1 u2_u0_u3_U48 (.A1( u2_u0_u3_n113 ) , .ZN( u2_u0_u3_n131 ) , .A2( u2_u0_u3_n154 ) );
  AOI21_X1 u2_u0_u3_U49 (.B2( u2_u0_u3_n114 ) , .B1( u2_u0_u3_n146 ) , .A( u2_u0_u3_n154 ) , .ZN( u2_u0_u3_n94 ) );
  INV_X1 u2_u0_u3_U5 (.A( u2_u0_u3_n117 ) , .ZN( u2_u0_u3_n178 ) );
  AOI21_X1 u2_u0_u3_U50 (.ZN( u2_u0_u3_n110 ) , .B2( u2_u0_u3_n142 ) , .B1( u2_u0_u3_n186 ) , .A( u2_u0_u3_n95 ) );
  INV_X1 u2_u0_u3_U51 (.A( u2_u0_u3_n145 ) , .ZN( u2_u0_u3_n186 ) );
  AOI21_X1 u2_u0_u3_U52 (.B1( u2_u0_u3_n124 ) , .A( u2_u0_u3_n149 ) , .B2( u2_u0_u3_n155 ) , .ZN( u2_u0_u3_n95 ) );
  INV_X1 u2_u0_u3_U53 (.A( u2_u0_u3_n141 ) , .ZN( u2_u0_u3_n167 ) );
  NAND2_X1 u2_u0_u3_U54 (.ZN( u2_u0_u3_n124 ) , .A1( u2_u0_u3_n96 ) , .A2( u2_u0_u3_n97 ) );
  NAND2_X1 u2_u0_u3_U55 (.A2( u2_u0_u3_n100 ) , .ZN( u2_u0_u3_n146 ) , .A1( u2_u0_u3_n96 ) );
  INV_X1 u2_u0_u3_U56 (.A( u2_u0_u3_n149 ) , .ZN( u2_u0_u3_n169 ) );
  NAND2_X1 u2_u0_u3_U57 (.A1( u2_u0_u3_n101 ) , .ZN( u2_u0_u3_n145 ) , .A2( u2_u0_u3_n99 ) );
  NAND2_X1 u2_u0_u3_U58 (.A1( u2_u0_u3_n100 ) , .ZN( u2_u0_u3_n156 ) , .A2( u2_u0_u3_n99 ) );
  NAND2_X1 u2_u0_u3_U59 (.A2( u2_u0_u3_n101 ) , .A1( u2_u0_u3_n104 ) , .ZN( u2_u0_u3_n148 ) );
  OAI22_X1 u2_u0_u3_U6 (.B2( u2_u0_u3_n147 ) , .A2( u2_u0_u3_n148 ) , .ZN( u2_u0_u3_n160 ) , .B1( u2_u0_u3_n165 ) , .A1( u2_u0_u3_n168 ) );
  NAND2_X1 u2_u0_u3_U60 (.A1( u2_u0_u3_n100 ) , .A2( u2_u0_u3_n102 ) , .ZN( u2_u0_u3_n128 ) );
  NAND2_X1 u2_u0_u3_U61 (.A2( u2_u0_u3_n101 ) , .A1( u2_u0_u3_n102 ) , .ZN( u2_u0_u3_n152 ) );
  NAND2_X1 u2_u0_u3_U62 (.A2( u2_u0_u3_n101 ) , .ZN( u2_u0_u3_n114 ) , .A1( u2_u0_u3_n96 ) );
  NAND2_X1 u2_u0_u3_U63 (.ZN( u2_u0_u3_n107 ) , .A1( u2_u0_u3_n97 ) , .A2( u2_u0_u3_n99 ) );
  NAND2_X1 u2_u0_u3_U64 (.A2( u2_u0_u3_n100 ) , .A1( u2_u0_u3_n104 ) , .ZN( u2_u0_u3_n113 ) );
  NAND2_X1 u2_u0_u3_U65 (.A1( u2_u0_u3_n104 ) , .ZN( u2_u0_u3_n153 ) , .A2( u2_u0_u3_n97 ) );
  NAND2_X1 u2_u0_u3_U66 (.A2( u2_u0_u3_n103 ) , .A1( u2_u0_u3_n104 ) , .ZN( u2_u0_u3_n130 ) );
  NAND2_X1 u2_u0_u3_U67 (.A2( u2_u0_u3_n103 ) , .ZN( u2_u0_u3_n144 ) , .A1( u2_u0_u3_n96 ) );
  NAND2_X1 u2_u0_u3_U68 (.A1( u2_u0_u3_n102 ) , .A2( u2_u0_u3_n103 ) , .ZN( u2_u0_u3_n108 ) );
  NOR2_X1 u2_u0_u3_U69 (.A2( u2_u0_X_19 ) , .A1( u2_u0_X_20 ) , .ZN( u2_u0_u3_n99 ) );
  AND3_X1 u2_u0_u3_U7 (.A3( u2_u0_u3_n144 ) , .A2( u2_u0_u3_n145 ) , .A1( u2_u0_u3_n146 ) , .ZN( u2_u0_u3_n147 ) );
  NOR2_X1 u2_u0_u3_U70 (.A2( u2_u0_X_21 ) , .A1( u2_u0_X_24 ) , .ZN( u2_u0_u3_n103 ) );
  NOR2_X1 u2_u0_u3_U71 (.A2( u2_u0_X_24 ) , .A1( u2_u0_u3_n171 ) , .ZN( u2_u0_u3_n97 ) );
  NOR2_X1 u2_u0_u3_U72 (.A2( u2_u0_X_23 ) , .ZN( u2_u0_u3_n141 ) , .A1( u2_u0_u3_n166 ) );
  NOR2_X1 u2_u0_u3_U73 (.A2( u2_u0_X_19 ) , .A1( u2_u0_u3_n172 ) , .ZN( u2_u0_u3_n96 ) );
  NAND2_X1 u2_u0_u3_U74 (.A1( u2_u0_X_22 ) , .A2( u2_u0_X_23 ) , .ZN( u2_u0_u3_n154 ) );
  NOR2_X1 u2_u0_u3_U75 (.A2( u2_u0_X_22 ) , .A1( u2_u0_X_23 ) , .ZN( u2_u0_u3_n121 ) );
  AND2_X1 u2_u0_u3_U76 (.A1( u2_u0_X_24 ) , .ZN( u2_u0_u3_n101 ) , .A2( u2_u0_u3_n171 ) );
  NAND2_X1 u2_u0_u3_U77 (.A1( u2_u0_X_23 ) , .ZN( u2_u0_u3_n149 ) , .A2( u2_u0_u3_n166 ) );
  AND2_X1 u2_u0_u3_U78 (.A1( u2_u0_X_19 ) , .ZN( u2_u0_u3_n102 ) , .A2( u2_u0_u3_n172 ) );
  AND2_X1 u2_u0_u3_U79 (.A1( u2_u0_X_21 ) , .A2( u2_u0_X_24 ) , .ZN( u2_u0_u3_n100 ) );
  INV_X1 u2_u0_u3_U8 (.A( u2_u0_u3_n143 ) , .ZN( u2_u0_u3_n168 ) );
  AND2_X1 u2_u0_u3_U80 (.A2( u2_u0_X_19 ) , .A1( u2_u0_X_20 ) , .ZN( u2_u0_u3_n104 ) );
  INV_X1 u2_u0_u3_U81 (.A( u2_u0_X_22 ) , .ZN( u2_u0_u3_n166 ) );
  INV_X1 u2_u0_u3_U82 (.A( u2_u0_X_21 ) , .ZN( u2_u0_u3_n171 ) );
  INV_X1 u2_u0_u3_U83 (.A( u2_u0_X_20 ) , .ZN( u2_u0_u3_n172 ) );
  NAND4_X1 u2_u0_u3_U84 (.ZN( u2_out0_26 ) , .A4( u2_u0_u3_n109 ) , .A3( u2_u0_u3_n110 ) , .A2( u2_u0_u3_n111 ) , .A1( u2_u0_u3_n173 ) );
  INV_X1 u2_u0_u3_U85 (.ZN( u2_u0_u3_n173 ) , .A( u2_u0_u3_n94 ) );
  OAI21_X1 u2_u0_u3_U86 (.ZN( u2_u0_u3_n111 ) , .B2( u2_u0_u3_n117 ) , .A( u2_u0_u3_n133 ) , .B1( u2_u0_u3_n176 ) );
  NAND4_X1 u2_u0_u3_U87 (.ZN( u2_out0_20 ) , .A4( u2_u0_u3_n122 ) , .A3( u2_u0_u3_n123 ) , .A1( u2_u0_u3_n175 ) , .A2( u2_u0_u3_n180 ) );
  INV_X1 u2_u0_u3_U88 (.A( u2_u0_u3_n126 ) , .ZN( u2_u0_u3_n180 ) );
  INV_X1 u2_u0_u3_U89 (.A( u2_u0_u3_n112 ) , .ZN( u2_u0_u3_n175 ) );
  OAI22_X1 u2_u0_u3_U9 (.B1( u2_u0_u3_n113 ) , .A2( u2_u0_u3_n135 ) , .A1( u2_u0_u3_n150 ) , .B2( u2_u0_u3_n164 ) , .ZN( u2_u0_u3_n98 ) );
  NAND4_X1 u2_u0_u3_U90 (.ZN( u2_out0_1 ) , .A4( u2_u0_u3_n161 ) , .A3( u2_u0_u3_n162 ) , .A2( u2_u0_u3_n163 ) , .A1( u2_u0_u3_n185 ) );
  NAND2_X1 u2_u0_u3_U91 (.ZN( u2_u0_u3_n163 ) , .A2( u2_u0_u3_n170 ) , .A1( u2_u0_u3_n176 ) );
  AOI22_X1 u2_u0_u3_U92 (.B2( u2_u0_u3_n140 ) , .B1( u2_u0_u3_n141 ) , .A2( u2_u0_u3_n142 ) , .ZN( u2_u0_u3_n162 ) , .A1( u2_u0_u3_n177 ) );
  OR4_X1 u2_u0_u3_U93 (.ZN( u2_out0_10 ) , .A4( u2_u0_u3_n136 ) , .A3( u2_u0_u3_n137 ) , .A1( u2_u0_u3_n138 ) , .A2( u2_u0_u3_n139 ) );
  OAI222_X1 u2_u0_u3_U94 (.C1( u2_u0_u3_n128 ) , .ZN( u2_u0_u3_n137 ) , .B1( u2_u0_u3_n148 ) , .A2( u2_u0_u3_n150 ) , .B2( u2_u0_u3_n154 ) , .C2( u2_u0_u3_n164 ) , .A1( u2_u0_u3_n167 ) );
  OAI221_X1 u2_u0_u3_U95 (.A( u2_u0_u3_n134 ) , .B2( u2_u0_u3_n135 ) , .ZN( u2_u0_u3_n136 ) , .C1( u2_u0_u3_n149 ) , .B1( u2_u0_u3_n151 ) , .C2( u2_u0_u3_n183 ) );
  AOI221_X1 u2_u0_u3_U96 (.A( u2_u0_u3_n131 ) , .C2( u2_u0_u3_n132 ) , .C1( u2_u0_u3_n133 ) , .ZN( u2_u0_u3_n134 ) , .B1( u2_u0_u3_n143 ) , .B2( u2_u0_u3_n177 ) );
  NAND2_X1 u2_u0_u3_U97 (.ZN( u2_u0_u3_n143 ) , .A1( u2_u0_u3_n165 ) , .A2( u2_u0_u3_n167 ) );
  NAND3_X1 u2_u0_u3_U98 (.A1( u2_u0_u3_n114 ) , .ZN( u2_u0_u3_n115 ) , .A2( u2_u0_u3_n145 ) , .A3( u2_u0_u3_n153 ) );
  NAND3_X1 u2_u0_u3_U99 (.ZN( u2_u0_u3_n129 ) , .A2( u2_u0_u3_n144 ) , .A1( u2_u0_u3_n153 ) , .A3( u2_u0_u3_n182 ) );
  XOR2_X1 u2_u11_U1 (.B( u2_K12_9 ) , .A( u2_R10_6 ) , .Z( u2_u11_X_9 ) );
  XOR2_X1 u2_u11_U16 (.B( u2_K12_3 ) , .A( u2_R10_2 ) , .Z( u2_u11_X_3 ) );
  XOR2_X1 u2_u11_U2 (.B( u2_K12_8 ) , .A( u2_R10_5 ) , .Z( u2_u11_X_8 ) );
  XOR2_X1 u2_u11_U27 (.B( u2_K12_2 ) , .A( u2_R10_1 ) , .Z( u2_u11_X_2 ) );
  XOR2_X1 u2_u11_U3 (.B( u2_K12_7 ) , .A( u2_R10_4 ) , .Z( u2_u11_X_7 ) );
  XOR2_X1 u2_u11_U38 (.B( u2_K12_1 ) , .A( u2_R10_32 ) , .Z( u2_u11_X_1 ) );
  XOR2_X1 u2_u11_U4 (.B( u2_K12_6 ) , .A( u2_R10_5 ) , .Z( u2_u11_X_6 ) );
  XOR2_X1 u2_u11_U40 (.B( u2_K12_18 ) , .A( u2_R10_13 ) , .Z( u2_u11_X_18 ) );
  XOR2_X1 u2_u11_U41 (.B( u2_K12_17 ) , .A( u2_R10_12 ) , .Z( u2_u11_X_17 ) );
  XOR2_X1 u2_u11_U42 (.B( u2_K12_16 ) , .A( u2_R10_11 ) , .Z( u2_u11_X_16 ) );
  XOR2_X1 u2_u11_U43 (.B( u2_K12_15 ) , .A( u2_R10_10 ) , .Z( u2_u11_X_15 ) );
  XOR2_X1 u2_u11_U44 (.B( u2_K12_14 ) , .A( u2_R10_9 ) , .Z( u2_u11_X_14 ) );
  XOR2_X1 u2_u11_U45 (.B( u2_K12_13 ) , .A( u2_R10_8 ) , .Z( u2_u11_X_13 ) );
  XOR2_X1 u2_u11_U46 (.B( u2_K12_12 ) , .A( u2_R10_9 ) , .Z( u2_u11_X_12 ) );
  XOR2_X1 u2_u11_U47 (.B( u2_K12_11 ) , .A( u2_R10_8 ) , .Z( u2_u11_X_11 ) );
  XOR2_X1 u2_u11_U48 (.B( u2_K12_10 ) , .A( u2_R10_7 ) , .Z( u2_u11_X_10 ) );
  XOR2_X1 u2_u11_U5 (.B( u2_K12_5 ) , .A( u2_R10_4 ) , .Z( u2_u11_X_5 ) );
  XOR2_X1 u2_u11_U6 (.B( u2_K12_4 ) , .A( u2_R10_3 ) , .Z( u2_u11_X_4 ) );
  NAND2_X1 u2_u11_u0_U10 (.ZN( u2_u11_u0_n113 ) , .A1( u2_u11_u0_n139 ) , .A2( u2_u11_u0_n149 ) );
  AND3_X1 u2_u11_u0_U11 (.A2( u2_u11_u0_n112 ) , .ZN( u2_u11_u0_n127 ) , .A3( u2_u11_u0_n130 ) , .A1( u2_u11_u0_n148 ) );
  AND2_X1 u2_u11_u0_U12 (.ZN( u2_u11_u0_n107 ) , .A1( u2_u11_u0_n130 ) , .A2( u2_u11_u0_n140 ) );
  AND2_X1 u2_u11_u0_U13 (.A2( u2_u11_u0_n129 ) , .A1( u2_u11_u0_n130 ) , .ZN( u2_u11_u0_n151 ) );
  AND2_X1 u2_u11_u0_U14 (.A1( u2_u11_u0_n108 ) , .A2( u2_u11_u0_n125 ) , .ZN( u2_u11_u0_n145 ) );
  INV_X1 u2_u11_u0_U15 (.A( u2_u11_u0_n143 ) , .ZN( u2_u11_u0_n173 ) );
  NOR2_X1 u2_u11_u0_U16 (.A2( u2_u11_u0_n136 ) , .ZN( u2_u11_u0_n147 ) , .A1( u2_u11_u0_n160 ) );
  OAI22_X1 u2_u11_u0_U17 (.B1( u2_u11_u0_n125 ) , .ZN( u2_u11_u0_n126 ) , .A1( u2_u11_u0_n138 ) , .A2( u2_u11_u0_n146 ) , .B2( u2_u11_u0_n147 ) );
  OAI22_X1 u2_u11_u0_U18 (.B1( u2_u11_u0_n131 ) , .A1( u2_u11_u0_n144 ) , .B2( u2_u11_u0_n147 ) , .A2( u2_u11_u0_n90 ) , .ZN( u2_u11_u0_n91 ) );
  AND3_X1 u2_u11_u0_U19 (.A3( u2_u11_u0_n121 ) , .A2( u2_u11_u0_n125 ) , .A1( u2_u11_u0_n148 ) , .ZN( u2_u11_u0_n90 ) );
  NOR2_X1 u2_u11_u0_U20 (.A1( u2_u11_u0_n163 ) , .A2( u2_u11_u0_n164 ) , .ZN( u2_u11_u0_n95 ) );
  NAND2_X1 u2_u11_u0_U21 (.A1( u2_u11_u0_n101 ) , .A2( u2_u11_u0_n102 ) , .ZN( u2_u11_u0_n150 ) );
  AOI22_X1 u2_u11_u0_U22 (.B2( u2_u11_u0_n109 ) , .A2( u2_u11_u0_n110 ) , .ZN( u2_u11_u0_n111 ) , .B1( u2_u11_u0_n118 ) , .A1( u2_u11_u0_n160 ) );
  NAND2_X1 u2_u11_u0_U23 (.A1( u2_u11_u0_n100 ) , .A2( u2_u11_u0_n103 ) , .ZN( u2_u11_u0_n125 ) );
  INV_X1 u2_u11_u0_U24 (.A( u2_u11_u0_n136 ) , .ZN( u2_u11_u0_n161 ) );
  INV_X1 u2_u11_u0_U25 (.A( u2_u11_u0_n118 ) , .ZN( u2_u11_u0_n158 ) );
  NAND2_X1 u2_u11_u0_U26 (.A2( u2_u11_u0_n100 ) , .A1( u2_u11_u0_n101 ) , .ZN( u2_u11_u0_n139 ) );
  NAND2_X1 u2_u11_u0_U27 (.A2( u2_u11_u0_n100 ) , .ZN( u2_u11_u0_n131 ) , .A1( u2_u11_u0_n92 ) );
  NAND2_X1 u2_u11_u0_U28 (.ZN( u2_u11_u0_n108 ) , .A1( u2_u11_u0_n92 ) , .A2( u2_u11_u0_n94 ) );
  AOI21_X1 u2_u11_u0_U29 (.B1( u2_u11_u0_n127 ) , .B2( u2_u11_u0_n129 ) , .A( u2_u11_u0_n138 ) , .ZN( u2_u11_u0_n96 ) );
  INV_X1 u2_u11_u0_U3 (.A( u2_u11_u0_n113 ) , .ZN( u2_u11_u0_n166 ) );
  AOI21_X1 u2_u11_u0_U30 (.ZN( u2_u11_u0_n104 ) , .B1( u2_u11_u0_n107 ) , .B2( u2_u11_u0_n141 ) , .A( u2_u11_u0_n144 ) );
  NAND2_X1 u2_u11_u0_U31 (.A2( u2_u11_u0_n102 ) , .ZN( u2_u11_u0_n114 ) , .A1( u2_u11_u0_n92 ) );
  NAND2_X1 u2_u11_u0_U32 (.A1( u2_u11_u0_n101 ) , .ZN( u2_u11_u0_n130 ) , .A2( u2_u11_u0_n94 ) );
  NOR2_X1 u2_u11_u0_U33 (.A1( u2_u11_u0_n120 ) , .ZN( u2_u11_u0_n143 ) , .A2( u2_u11_u0_n167 ) );
  OAI221_X1 u2_u11_u0_U34 (.C1( u2_u11_u0_n112 ) , .ZN( u2_u11_u0_n120 ) , .B1( u2_u11_u0_n138 ) , .B2( u2_u11_u0_n141 ) , .C2( u2_u11_u0_n147 ) , .A( u2_u11_u0_n172 ) );
  AOI211_X1 u2_u11_u0_U35 (.B( u2_u11_u0_n115 ) , .A( u2_u11_u0_n116 ) , .C2( u2_u11_u0_n117 ) , .C1( u2_u11_u0_n118 ) , .ZN( u2_u11_u0_n119 ) );
  NAND2_X1 u2_u11_u0_U36 (.A2( u2_u11_u0_n103 ) , .ZN( u2_u11_u0_n140 ) , .A1( u2_u11_u0_n94 ) );
  INV_X1 u2_u11_u0_U37 (.A( u2_u11_u0_n138 ) , .ZN( u2_u11_u0_n160 ) );
  NAND2_X1 u2_u11_u0_U38 (.A2( u2_u11_u0_n102 ) , .A1( u2_u11_u0_n103 ) , .ZN( u2_u11_u0_n149 ) );
  NAND2_X1 u2_u11_u0_U39 (.A2( u2_u11_u0_n101 ) , .ZN( u2_u11_u0_n121 ) , .A1( u2_u11_u0_n93 ) );
  AOI21_X1 u2_u11_u0_U4 (.B1( u2_u11_u0_n114 ) , .ZN( u2_u11_u0_n115 ) , .B2( u2_u11_u0_n129 ) , .A( u2_u11_u0_n161 ) );
  NAND2_X1 u2_u11_u0_U40 (.ZN( u2_u11_u0_n112 ) , .A2( u2_u11_u0_n92 ) , .A1( u2_u11_u0_n93 ) );
  INV_X1 u2_u11_u0_U41 (.ZN( u2_u11_u0_n172 ) , .A( u2_u11_u0_n88 ) );
  OAI222_X1 u2_u11_u0_U42 (.C1( u2_u11_u0_n108 ) , .A1( u2_u11_u0_n125 ) , .B2( u2_u11_u0_n128 ) , .B1( u2_u11_u0_n144 ) , .A2( u2_u11_u0_n158 ) , .C2( u2_u11_u0_n161 ) , .ZN( u2_u11_u0_n88 ) );
  AOI21_X1 u2_u11_u0_U43 (.B1( u2_u11_u0_n103 ) , .ZN( u2_u11_u0_n132 ) , .A( u2_u11_u0_n165 ) , .B2( u2_u11_u0_n93 ) );
  OR3_X1 u2_u11_u0_U44 (.A3( u2_u11_u0_n152 ) , .A2( u2_u11_u0_n153 ) , .A1( u2_u11_u0_n154 ) , .ZN( u2_u11_u0_n155 ) );
  AOI21_X1 u2_u11_u0_U45 (.A( u2_u11_u0_n144 ) , .B2( u2_u11_u0_n145 ) , .B1( u2_u11_u0_n146 ) , .ZN( u2_u11_u0_n154 ) );
  AOI21_X1 u2_u11_u0_U46 (.B2( u2_u11_u0_n150 ) , .B1( u2_u11_u0_n151 ) , .ZN( u2_u11_u0_n152 ) , .A( u2_u11_u0_n158 ) );
  AOI21_X1 u2_u11_u0_U47 (.A( u2_u11_u0_n147 ) , .B2( u2_u11_u0_n148 ) , .B1( u2_u11_u0_n149 ) , .ZN( u2_u11_u0_n153 ) );
  INV_X1 u2_u11_u0_U48 (.ZN( u2_u11_u0_n171 ) , .A( u2_u11_u0_n99 ) );
  OAI211_X1 u2_u11_u0_U49 (.C2( u2_u11_u0_n140 ) , .C1( u2_u11_u0_n161 ) , .A( u2_u11_u0_n169 ) , .B( u2_u11_u0_n98 ) , .ZN( u2_u11_u0_n99 ) );
  AOI21_X1 u2_u11_u0_U5 (.B2( u2_u11_u0_n131 ) , .ZN( u2_u11_u0_n134 ) , .B1( u2_u11_u0_n151 ) , .A( u2_u11_u0_n158 ) );
  AOI211_X1 u2_u11_u0_U50 (.C1( u2_u11_u0_n118 ) , .A( u2_u11_u0_n123 ) , .B( u2_u11_u0_n96 ) , .C2( u2_u11_u0_n97 ) , .ZN( u2_u11_u0_n98 ) );
  INV_X1 u2_u11_u0_U51 (.ZN( u2_u11_u0_n169 ) , .A( u2_u11_u0_n91 ) );
  NOR2_X1 u2_u11_u0_U52 (.A2( u2_u11_X_2 ) , .ZN( u2_u11_u0_n103 ) , .A1( u2_u11_u0_n164 ) );
  NOR2_X1 u2_u11_u0_U53 (.A2( u2_u11_X_4 ) , .A1( u2_u11_X_5 ) , .ZN( u2_u11_u0_n118 ) );
  NOR2_X1 u2_u11_u0_U54 (.A2( u2_u11_X_3 ) , .A1( u2_u11_X_6 ) , .ZN( u2_u11_u0_n94 ) );
  NAND2_X1 u2_u11_u0_U55 (.A2( u2_u11_X_4 ) , .A1( u2_u11_X_5 ) , .ZN( u2_u11_u0_n144 ) );
  NOR2_X1 u2_u11_u0_U56 (.A2( u2_u11_X_5 ) , .ZN( u2_u11_u0_n136 ) , .A1( u2_u11_u0_n159 ) );
  NAND2_X1 u2_u11_u0_U57 (.A1( u2_u11_X_5 ) , .ZN( u2_u11_u0_n138 ) , .A2( u2_u11_u0_n159 ) );
  AND2_X1 u2_u11_u0_U58 (.A2( u2_u11_X_3 ) , .A1( u2_u11_X_6 ) , .ZN( u2_u11_u0_n102 ) );
  AND2_X1 u2_u11_u0_U59 (.A1( u2_u11_X_6 ) , .A2( u2_u11_u0_n162 ) , .ZN( u2_u11_u0_n93 ) );
  NOR2_X1 u2_u11_u0_U6 (.A1( u2_u11_u0_n108 ) , .ZN( u2_u11_u0_n123 ) , .A2( u2_u11_u0_n158 ) );
  INV_X1 u2_u11_u0_U60 (.A( u2_u11_X_4 ) , .ZN( u2_u11_u0_n159 ) );
  INV_X1 u2_u11_u0_U61 (.A( u2_u11_X_2 ) , .ZN( u2_u11_u0_n163 ) );
  INV_X1 u2_u11_u0_U62 (.A( u2_u11_u0_n126 ) , .ZN( u2_u11_u0_n168 ) );
  AOI211_X1 u2_u11_u0_U63 (.B( u2_u11_u0_n133 ) , .A( u2_u11_u0_n134 ) , .C2( u2_u11_u0_n135 ) , .C1( u2_u11_u0_n136 ) , .ZN( u2_u11_u0_n137 ) );
  OR4_X1 u2_u11_u0_U64 (.ZN( u2_out11_17 ) , .A4( u2_u11_u0_n122 ) , .A2( u2_u11_u0_n123 ) , .A1( u2_u11_u0_n124 ) , .A3( u2_u11_u0_n170 ) );
  AOI21_X1 u2_u11_u0_U65 (.B2( u2_u11_u0_n107 ) , .ZN( u2_u11_u0_n124 ) , .B1( u2_u11_u0_n128 ) , .A( u2_u11_u0_n161 ) );
  INV_X1 u2_u11_u0_U66 (.A( u2_u11_u0_n111 ) , .ZN( u2_u11_u0_n170 ) );
  OR4_X1 u2_u11_u0_U67 (.ZN( u2_out11_31 ) , .A4( u2_u11_u0_n155 ) , .A2( u2_u11_u0_n156 ) , .A1( u2_u11_u0_n157 ) , .A3( u2_u11_u0_n173 ) );
  AOI21_X1 u2_u11_u0_U68 (.A( u2_u11_u0_n138 ) , .B2( u2_u11_u0_n139 ) , .B1( u2_u11_u0_n140 ) , .ZN( u2_u11_u0_n157 ) );
  INV_X1 u2_u11_u0_U69 (.ZN( u2_u11_u0_n174 ) , .A( u2_u11_u0_n89 ) );
  OAI21_X1 u2_u11_u0_U7 (.B1( u2_u11_u0_n150 ) , .B2( u2_u11_u0_n158 ) , .A( u2_u11_u0_n172 ) , .ZN( u2_u11_u0_n89 ) );
  AOI211_X1 u2_u11_u0_U70 (.B( u2_u11_u0_n104 ) , .A( u2_u11_u0_n105 ) , .ZN( u2_u11_u0_n106 ) , .C2( u2_u11_u0_n113 ) , .C1( u2_u11_u0_n160 ) );
  INV_X1 u2_u11_u0_U71 (.A( u2_u11_u0_n142 ) , .ZN( u2_u11_u0_n165 ) );
  AOI21_X1 u2_u11_u0_U72 (.ZN( u2_u11_u0_n116 ) , .B2( u2_u11_u0_n142 ) , .A( u2_u11_u0_n144 ) , .B1( u2_u11_u0_n166 ) );
  AOI21_X1 u2_u11_u0_U73 (.B2( u2_u11_u0_n141 ) , .B1( u2_u11_u0_n142 ) , .ZN( u2_u11_u0_n156 ) , .A( u2_u11_u0_n161 ) );
  OAI221_X1 u2_u11_u0_U74 (.C1( u2_u11_u0_n121 ) , .ZN( u2_u11_u0_n122 ) , .B2( u2_u11_u0_n127 ) , .A( u2_u11_u0_n143 ) , .B1( u2_u11_u0_n144 ) , .C2( u2_u11_u0_n147 ) );
  NOR2_X1 u2_u11_u0_U75 (.A2( u2_u11_X_6 ) , .ZN( u2_u11_u0_n100 ) , .A1( u2_u11_u0_n162 ) );
  INV_X1 u2_u11_u0_U76 (.A( u2_u11_X_3 ) , .ZN( u2_u11_u0_n162 ) );
  AOI21_X1 u2_u11_u0_U77 (.B1( u2_u11_u0_n132 ) , .ZN( u2_u11_u0_n133 ) , .A( u2_u11_u0_n144 ) , .B2( u2_u11_u0_n166 ) );
  OAI22_X1 u2_u11_u0_U78 (.ZN( u2_u11_u0_n105 ) , .A2( u2_u11_u0_n132 ) , .B1( u2_u11_u0_n146 ) , .A1( u2_u11_u0_n147 ) , .B2( u2_u11_u0_n161 ) );
  NAND2_X1 u2_u11_u0_U79 (.ZN( u2_u11_u0_n110 ) , .A2( u2_u11_u0_n132 ) , .A1( u2_u11_u0_n145 ) );
  AND2_X1 u2_u11_u0_U8 (.A1( u2_u11_u0_n114 ) , .A2( u2_u11_u0_n121 ) , .ZN( u2_u11_u0_n146 ) );
  INV_X1 u2_u11_u0_U80 (.A( u2_u11_u0_n119 ) , .ZN( u2_u11_u0_n167 ) );
  NAND2_X1 u2_u11_u0_U81 (.ZN( u2_u11_u0_n148 ) , .A1( u2_u11_u0_n93 ) , .A2( u2_u11_u0_n95 ) );
  NAND2_X1 u2_u11_u0_U82 (.A1( u2_u11_u0_n100 ) , .ZN( u2_u11_u0_n129 ) , .A2( u2_u11_u0_n95 ) );
  NAND2_X1 u2_u11_u0_U83 (.A1( u2_u11_u0_n102 ) , .ZN( u2_u11_u0_n128 ) , .A2( u2_u11_u0_n95 ) );
  NOR2_X1 u2_u11_u0_U84 (.A2( u2_u11_X_1 ) , .A1( u2_u11_X_2 ) , .ZN( u2_u11_u0_n92 ) );
  NAND2_X1 u2_u11_u0_U85 (.ZN( u2_u11_u0_n142 ) , .A1( u2_u11_u0_n94 ) , .A2( u2_u11_u0_n95 ) );
  NOR2_X1 u2_u11_u0_U86 (.A2( u2_u11_X_1 ) , .ZN( u2_u11_u0_n101 ) , .A1( u2_u11_u0_n163 ) );
  INV_X1 u2_u11_u0_U87 (.A( u2_u11_X_1 ) , .ZN( u2_u11_u0_n164 ) );
  NAND3_X1 u2_u11_u0_U88 (.ZN( u2_out11_23 ) , .A3( u2_u11_u0_n137 ) , .A1( u2_u11_u0_n168 ) , .A2( u2_u11_u0_n171 ) );
  NAND3_X1 u2_u11_u0_U89 (.A3( u2_u11_u0_n127 ) , .A2( u2_u11_u0_n128 ) , .ZN( u2_u11_u0_n135 ) , .A1( u2_u11_u0_n150 ) );
  AND2_X1 u2_u11_u0_U9 (.A1( u2_u11_u0_n131 ) , .ZN( u2_u11_u0_n141 ) , .A2( u2_u11_u0_n150 ) );
  NAND3_X1 u2_u11_u0_U90 (.ZN( u2_u11_u0_n117 ) , .A3( u2_u11_u0_n132 ) , .A2( u2_u11_u0_n139 ) , .A1( u2_u11_u0_n148 ) );
  NAND3_X1 u2_u11_u0_U91 (.ZN( u2_u11_u0_n109 ) , .A2( u2_u11_u0_n114 ) , .A3( u2_u11_u0_n140 ) , .A1( u2_u11_u0_n149 ) );
  NAND3_X1 u2_u11_u0_U92 (.ZN( u2_out11_9 ) , .A3( u2_u11_u0_n106 ) , .A2( u2_u11_u0_n171 ) , .A1( u2_u11_u0_n174 ) );
  NAND3_X1 u2_u11_u0_U93 (.A2( u2_u11_u0_n128 ) , .A1( u2_u11_u0_n132 ) , .A3( u2_u11_u0_n146 ) , .ZN( u2_u11_u0_n97 ) );
  NOR2_X1 u2_u11_u1_U10 (.A1( u2_u11_u1_n112 ) , .A2( u2_u11_u1_n116 ) , .ZN( u2_u11_u1_n118 ) );
  NAND3_X1 u2_u11_u1_U100 (.ZN( u2_u11_u1_n113 ) , .A1( u2_u11_u1_n120 ) , .A3( u2_u11_u1_n133 ) , .A2( u2_u11_u1_n155 ) );
  OAI21_X1 u2_u11_u1_U11 (.ZN( u2_u11_u1_n101 ) , .B1( u2_u11_u1_n141 ) , .A( u2_u11_u1_n146 ) , .B2( u2_u11_u1_n183 ) );
  AOI21_X1 u2_u11_u1_U12 (.B2( u2_u11_u1_n155 ) , .B1( u2_u11_u1_n156 ) , .ZN( u2_u11_u1_n157 ) , .A( u2_u11_u1_n174 ) );
  NAND2_X1 u2_u11_u1_U13 (.ZN( u2_u11_u1_n140 ) , .A2( u2_u11_u1_n150 ) , .A1( u2_u11_u1_n155 ) );
  NAND2_X1 u2_u11_u1_U14 (.A1( u2_u11_u1_n131 ) , .ZN( u2_u11_u1_n147 ) , .A2( u2_u11_u1_n153 ) );
  INV_X1 u2_u11_u1_U15 (.A( u2_u11_u1_n139 ) , .ZN( u2_u11_u1_n174 ) );
  OR4_X1 u2_u11_u1_U16 (.A4( u2_u11_u1_n106 ) , .A3( u2_u11_u1_n107 ) , .ZN( u2_u11_u1_n108 ) , .A1( u2_u11_u1_n117 ) , .A2( u2_u11_u1_n184 ) );
  AOI21_X1 u2_u11_u1_U17 (.ZN( u2_u11_u1_n106 ) , .A( u2_u11_u1_n112 ) , .B1( u2_u11_u1_n154 ) , .B2( u2_u11_u1_n156 ) );
  AOI21_X1 u2_u11_u1_U18 (.ZN( u2_u11_u1_n107 ) , .B1( u2_u11_u1_n134 ) , .B2( u2_u11_u1_n149 ) , .A( u2_u11_u1_n174 ) );
  INV_X1 u2_u11_u1_U19 (.A( u2_u11_u1_n101 ) , .ZN( u2_u11_u1_n184 ) );
  INV_X1 u2_u11_u1_U20 (.A( u2_u11_u1_n112 ) , .ZN( u2_u11_u1_n171 ) );
  NAND2_X1 u2_u11_u1_U21 (.ZN( u2_u11_u1_n141 ) , .A1( u2_u11_u1_n153 ) , .A2( u2_u11_u1_n156 ) );
  AND2_X1 u2_u11_u1_U22 (.A1( u2_u11_u1_n123 ) , .ZN( u2_u11_u1_n134 ) , .A2( u2_u11_u1_n161 ) );
  NAND2_X1 u2_u11_u1_U23 (.A2( u2_u11_u1_n115 ) , .A1( u2_u11_u1_n116 ) , .ZN( u2_u11_u1_n148 ) );
  NAND2_X1 u2_u11_u1_U24 (.A2( u2_u11_u1_n133 ) , .A1( u2_u11_u1_n135 ) , .ZN( u2_u11_u1_n159 ) );
  NAND2_X1 u2_u11_u1_U25 (.A2( u2_u11_u1_n115 ) , .A1( u2_u11_u1_n120 ) , .ZN( u2_u11_u1_n132 ) );
  INV_X1 u2_u11_u1_U26 (.A( u2_u11_u1_n154 ) , .ZN( u2_u11_u1_n178 ) );
  INV_X1 u2_u11_u1_U27 (.A( u2_u11_u1_n151 ) , .ZN( u2_u11_u1_n183 ) );
  AND2_X1 u2_u11_u1_U28 (.A1( u2_u11_u1_n129 ) , .A2( u2_u11_u1_n133 ) , .ZN( u2_u11_u1_n149 ) );
  INV_X1 u2_u11_u1_U29 (.A( u2_u11_u1_n131 ) , .ZN( u2_u11_u1_n180 ) );
  INV_X1 u2_u11_u1_U3 (.A( u2_u11_u1_n159 ) , .ZN( u2_u11_u1_n182 ) );
  OAI221_X1 u2_u11_u1_U30 (.A( u2_u11_u1_n119 ) , .C2( u2_u11_u1_n129 ) , .ZN( u2_u11_u1_n138 ) , .B2( u2_u11_u1_n152 ) , .C1( u2_u11_u1_n174 ) , .B1( u2_u11_u1_n187 ) );
  INV_X1 u2_u11_u1_U31 (.A( u2_u11_u1_n148 ) , .ZN( u2_u11_u1_n187 ) );
  AOI211_X1 u2_u11_u1_U32 (.B( u2_u11_u1_n117 ) , .A( u2_u11_u1_n118 ) , .ZN( u2_u11_u1_n119 ) , .C2( u2_u11_u1_n146 ) , .C1( u2_u11_u1_n159 ) );
  NOR2_X1 u2_u11_u1_U33 (.A1( u2_u11_u1_n168 ) , .A2( u2_u11_u1_n176 ) , .ZN( u2_u11_u1_n98 ) );
  AOI211_X1 u2_u11_u1_U34 (.B( u2_u11_u1_n162 ) , .A( u2_u11_u1_n163 ) , .C2( u2_u11_u1_n164 ) , .ZN( u2_u11_u1_n165 ) , .C1( u2_u11_u1_n171 ) );
  AOI21_X1 u2_u11_u1_U35 (.A( u2_u11_u1_n160 ) , .B2( u2_u11_u1_n161 ) , .ZN( u2_u11_u1_n162 ) , .B1( u2_u11_u1_n182 ) );
  OR2_X1 u2_u11_u1_U36 (.A2( u2_u11_u1_n157 ) , .A1( u2_u11_u1_n158 ) , .ZN( u2_u11_u1_n163 ) );
  NAND2_X1 u2_u11_u1_U37 (.A1( u2_u11_u1_n128 ) , .ZN( u2_u11_u1_n146 ) , .A2( u2_u11_u1_n160 ) );
  NAND2_X1 u2_u11_u1_U38 (.A2( u2_u11_u1_n112 ) , .ZN( u2_u11_u1_n139 ) , .A1( u2_u11_u1_n152 ) );
  NAND2_X1 u2_u11_u1_U39 (.A1( u2_u11_u1_n105 ) , .ZN( u2_u11_u1_n156 ) , .A2( u2_u11_u1_n99 ) );
  AOI221_X1 u2_u11_u1_U4 (.A( u2_u11_u1_n138 ) , .C2( u2_u11_u1_n139 ) , .C1( u2_u11_u1_n140 ) , .B2( u2_u11_u1_n141 ) , .ZN( u2_u11_u1_n142 ) , .B1( u2_u11_u1_n175 ) );
  AOI221_X1 u2_u11_u1_U40 (.B1( u2_u11_u1_n140 ) , .ZN( u2_u11_u1_n167 ) , .B2( u2_u11_u1_n172 ) , .C2( u2_u11_u1_n175 ) , .C1( u2_u11_u1_n178 ) , .A( u2_u11_u1_n188 ) );
  INV_X1 u2_u11_u1_U41 (.ZN( u2_u11_u1_n188 ) , .A( u2_u11_u1_n97 ) );
  AOI211_X1 u2_u11_u1_U42 (.A( u2_u11_u1_n118 ) , .C1( u2_u11_u1_n132 ) , .C2( u2_u11_u1_n139 ) , .B( u2_u11_u1_n96 ) , .ZN( u2_u11_u1_n97 ) );
  AOI21_X1 u2_u11_u1_U43 (.B2( u2_u11_u1_n121 ) , .B1( u2_u11_u1_n135 ) , .A( u2_u11_u1_n152 ) , .ZN( u2_u11_u1_n96 ) );
  NOR2_X1 u2_u11_u1_U44 (.ZN( u2_u11_u1_n117 ) , .A1( u2_u11_u1_n121 ) , .A2( u2_u11_u1_n160 ) );
  OAI21_X1 u2_u11_u1_U45 (.B2( u2_u11_u1_n123 ) , .ZN( u2_u11_u1_n145 ) , .B1( u2_u11_u1_n160 ) , .A( u2_u11_u1_n185 ) );
  INV_X1 u2_u11_u1_U46 (.A( u2_u11_u1_n122 ) , .ZN( u2_u11_u1_n185 ) );
  AOI21_X1 u2_u11_u1_U47 (.B2( u2_u11_u1_n120 ) , .B1( u2_u11_u1_n121 ) , .ZN( u2_u11_u1_n122 ) , .A( u2_u11_u1_n128 ) );
  AOI21_X1 u2_u11_u1_U48 (.A( u2_u11_u1_n128 ) , .B2( u2_u11_u1_n129 ) , .ZN( u2_u11_u1_n130 ) , .B1( u2_u11_u1_n150 ) );
  NAND2_X1 u2_u11_u1_U49 (.ZN( u2_u11_u1_n112 ) , .A1( u2_u11_u1_n169 ) , .A2( u2_u11_u1_n170 ) );
  AOI211_X1 u2_u11_u1_U5 (.ZN( u2_u11_u1_n124 ) , .A( u2_u11_u1_n138 ) , .C2( u2_u11_u1_n139 ) , .B( u2_u11_u1_n145 ) , .C1( u2_u11_u1_n147 ) );
  NAND2_X1 u2_u11_u1_U50 (.ZN( u2_u11_u1_n129 ) , .A2( u2_u11_u1_n95 ) , .A1( u2_u11_u1_n98 ) );
  NAND2_X1 u2_u11_u1_U51 (.A1( u2_u11_u1_n102 ) , .ZN( u2_u11_u1_n154 ) , .A2( u2_u11_u1_n99 ) );
  NAND2_X1 u2_u11_u1_U52 (.A2( u2_u11_u1_n100 ) , .ZN( u2_u11_u1_n135 ) , .A1( u2_u11_u1_n99 ) );
  AOI21_X1 u2_u11_u1_U53 (.A( u2_u11_u1_n152 ) , .B2( u2_u11_u1_n153 ) , .B1( u2_u11_u1_n154 ) , .ZN( u2_u11_u1_n158 ) );
  INV_X1 u2_u11_u1_U54 (.A( u2_u11_u1_n160 ) , .ZN( u2_u11_u1_n175 ) );
  NAND2_X1 u2_u11_u1_U55 (.A1( u2_u11_u1_n100 ) , .ZN( u2_u11_u1_n116 ) , .A2( u2_u11_u1_n95 ) );
  NAND2_X1 u2_u11_u1_U56 (.A1( u2_u11_u1_n102 ) , .ZN( u2_u11_u1_n131 ) , .A2( u2_u11_u1_n95 ) );
  NAND2_X1 u2_u11_u1_U57 (.A2( u2_u11_u1_n104 ) , .ZN( u2_u11_u1_n121 ) , .A1( u2_u11_u1_n98 ) );
  NAND2_X1 u2_u11_u1_U58 (.A1( u2_u11_u1_n103 ) , .ZN( u2_u11_u1_n153 ) , .A2( u2_u11_u1_n98 ) );
  NAND2_X1 u2_u11_u1_U59 (.A2( u2_u11_u1_n104 ) , .A1( u2_u11_u1_n105 ) , .ZN( u2_u11_u1_n133 ) );
  AOI22_X1 u2_u11_u1_U6 (.B2( u2_u11_u1_n113 ) , .A2( u2_u11_u1_n114 ) , .ZN( u2_u11_u1_n125 ) , .A1( u2_u11_u1_n171 ) , .B1( u2_u11_u1_n173 ) );
  NAND2_X1 u2_u11_u1_U60 (.ZN( u2_u11_u1_n150 ) , .A2( u2_u11_u1_n98 ) , .A1( u2_u11_u1_n99 ) );
  NAND2_X1 u2_u11_u1_U61 (.A1( u2_u11_u1_n105 ) , .ZN( u2_u11_u1_n155 ) , .A2( u2_u11_u1_n95 ) );
  OAI21_X1 u2_u11_u1_U62 (.ZN( u2_u11_u1_n109 ) , .B1( u2_u11_u1_n129 ) , .B2( u2_u11_u1_n160 ) , .A( u2_u11_u1_n167 ) );
  NAND2_X1 u2_u11_u1_U63 (.A2( u2_u11_u1_n100 ) , .A1( u2_u11_u1_n103 ) , .ZN( u2_u11_u1_n120 ) );
  NAND2_X1 u2_u11_u1_U64 (.A1( u2_u11_u1_n102 ) , .A2( u2_u11_u1_n104 ) , .ZN( u2_u11_u1_n115 ) );
  NAND2_X1 u2_u11_u1_U65 (.A2( u2_u11_u1_n100 ) , .A1( u2_u11_u1_n104 ) , .ZN( u2_u11_u1_n151 ) );
  NAND2_X1 u2_u11_u1_U66 (.A2( u2_u11_u1_n103 ) , .A1( u2_u11_u1_n105 ) , .ZN( u2_u11_u1_n161 ) );
  INV_X1 u2_u11_u1_U67 (.A( u2_u11_u1_n152 ) , .ZN( u2_u11_u1_n173 ) );
  INV_X1 u2_u11_u1_U68 (.A( u2_u11_u1_n128 ) , .ZN( u2_u11_u1_n172 ) );
  NAND2_X1 u2_u11_u1_U69 (.A2( u2_u11_u1_n102 ) , .A1( u2_u11_u1_n103 ) , .ZN( u2_u11_u1_n123 ) );
  NAND2_X1 u2_u11_u1_U7 (.ZN( u2_u11_u1_n114 ) , .A1( u2_u11_u1_n134 ) , .A2( u2_u11_u1_n156 ) );
  NOR2_X1 u2_u11_u1_U70 (.A2( u2_u11_X_7 ) , .A1( u2_u11_X_8 ) , .ZN( u2_u11_u1_n95 ) );
  NOR2_X1 u2_u11_u1_U71 (.A1( u2_u11_X_12 ) , .A2( u2_u11_X_9 ) , .ZN( u2_u11_u1_n100 ) );
  NOR2_X1 u2_u11_u1_U72 (.A2( u2_u11_X_8 ) , .A1( u2_u11_u1_n177 ) , .ZN( u2_u11_u1_n99 ) );
  NOR2_X1 u2_u11_u1_U73 (.A2( u2_u11_X_12 ) , .ZN( u2_u11_u1_n102 ) , .A1( u2_u11_u1_n176 ) );
  NOR2_X1 u2_u11_u1_U74 (.A2( u2_u11_X_9 ) , .ZN( u2_u11_u1_n105 ) , .A1( u2_u11_u1_n168 ) );
  NAND2_X1 u2_u11_u1_U75 (.A1( u2_u11_X_10 ) , .ZN( u2_u11_u1_n160 ) , .A2( u2_u11_u1_n169 ) );
  NAND2_X1 u2_u11_u1_U76 (.A2( u2_u11_X_10 ) , .A1( u2_u11_X_11 ) , .ZN( u2_u11_u1_n152 ) );
  NAND2_X1 u2_u11_u1_U77 (.A1( u2_u11_X_11 ) , .ZN( u2_u11_u1_n128 ) , .A2( u2_u11_u1_n170 ) );
  AND2_X1 u2_u11_u1_U78 (.A2( u2_u11_X_7 ) , .A1( u2_u11_X_8 ) , .ZN( u2_u11_u1_n104 ) );
  AND2_X1 u2_u11_u1_U79 (.A1( u2_u11_X_8 ) , .ZN( u2_u11_u1_n103 ) , .A2( u2_u11_u1_n177 ) );
  AOI22_X1 u2_u11_u1_U8 (.B2( u2_u11_u1_n136 ) , .A2( u2_u11_u1_n137 ) , .ZN( u2_u11_u1_n143 ) , .A1( u2_u11_u1_n171 ) , .B1( u2_u11_u1_n173 ) );
  INV_X1 u2_u11_u1_U80 (.A( u2_u11_X_10 ) , .ZN( u2_u11_u1_n170 ) );
  INV_X1 u2_u11_u1_U81 (.A( u2_u11_X_9 ) , .ZN( u2_u11_u1_n176 ) );
  INV_X1 u2_u11_u1_U82 (.A( u2_u11_X_11 ) , .ZN( u2_u11_u1_n169 ) );
  INV_X1 u2_u11_u1_U83 (.A( u2_u11_X_12 ) , .ZN( u2_u11_u1_n168 ) );
  INV_X1 u2_u11_u1_U84 (.A( u2_u11_X_7 ) , .ZN( u2_u11_u1_n177 ) );
  NAND4_X1 u2_u11_u1_U85 (.ZN( u2_out11_28 ) , .A4( u2_u11_u1_n124 ) , .A3( u2_u11_u1_n125 ) , .A2( u2_u11_u1_n126 ) , .A1( u2_u11_u1_n127 ) );
  OAI21_X1 u2_u11_u1_U86 (.ZN( u2_u11_u1_n127 ) , .B2( u2_u11_u1_n139 ) , .B1( u2_u11_u1_n175 ) , .A( u2_u11_u1_n183 ) );
  OAI21_X1 u2_u11_u1_U87 (.ZN( u2_u11_u1_n126 ) , .B2( u2_u11_u1_n140 ) , .A( u2_u11_u1_n146 ) , .B1( u2_u11_u1_n178 ) );
  NAND4_X1 u2_u11_u1_U88 (.ZN( u2_out11_18 ) , .A4( u2_u11_u1_n165 ) , .A3( u2_u11_u1_n166 ) , .A1( u2_u11_u1_n167 ) , .A2( u2_u11_u1_n186 ) );
  AOI22_X1 u2_u11_u1_U89 (.B2( u2_u11_u1_n146 ) , .B1( u2_u11_u1_n147 ) , .A2( u2_u11_u1_n148 ) , .ZN( u2_u11_u1_n166 ) , .A1( u2_u11_u1_n172 ) );
  INV_X1 u2_u11_u1_U9 (.A( u2_u11_u1_n147 ) , .ZN( u2_u11_u1_n181 ) );
  INV_X1 u2_u11_u1_U90 (.A( u2_u11_u1_n145 ) , .ZN( u2_u11_u1_n186 ) );
  NAND4_X1 u2_u11_u1_U91 (.ZN( u2_out11_2 ) , .A4( u2_u11_u1_n142 ) , .A3( u2_u11_u1_n143 ) , .A2( u2_u11_u1_n144 ) , .A1( u2_u11_u1_n179 ) );
  OAI21_X1 u2_u11_u1_U92 (.B2( u2_u11_u1_n132 ) , .ZN( u2_u11_u1_n144 ) , .A( u2_u11_u1_n146 ) , .B1( u2_u11_u1_n180 ) );
  INV_X1 u2_u11_u1_U93 (.A( u2_u11_u1_n130 ) , .ZN( u2_u11_u1_n179 ) );
  OR4_X1 u2_u11_u1_U94 (.ZN( u2_out11_13 ) , .A4( u2_u11_u1_n108 ) , .A3( u2_u11_u1_n109 ) , .A2( u2_u11_u1_n110 ) , .A1( u2_u11_u1_n111 ) );
  AOI21_X1 u2_u11_u1_U95 (.ZN( u2_u11_u1_n111 ) , .A( u2_u11_u1_n128 ) , .B2( u2_u11_u1_n131 ) , .B1( u2_u11_u1_n135 ) );
  AOI21_X1 u2_u11_u1_U96 (.ZN( u2_u11_u1_n110 ) , .A( u2_u11_u1_n116 ) , .B1( u2_u11_u1_n152 ) , .B2( u2_u11_u1_n160 ) );
  NAND3_X1 u2_u11_u1_U97 (.A3( u2_u11_u1_n149 ) , .A2( u2_u11_u1_n150 ) , .A1( u2_u11_u1_n151 ) , .ZN( u2_u11_u1_n164 ) );
  NAND3_X1 u2_u11_u1_U98 (.A3( u2_u11_u1_n134 ) , .A2( u2_u11_u1_n135 ) , .ZN( u2_u11_u1_n136 ) , .A1( u2_u11_u1_n151 ) );
  NAND3_X1 u2_u11_u1_U99 (.A1( u2_u11_u1_n133 ) , .ZN( u2_u11_u1_n137 ) , .A2( u2_u11_u1_n154 ) , .A3( u2_u11_u1_n181 ) );
  OAI22_X1 u2_u11_u2_U10 (.ZN( u2_u11_u2_n109 ) , .A2( u2_u11_u2_n113 ) , .B2( u2_u11_u2_n133 ) , .B1( u2_u11_u2_n167 ) , .A1( u2_u11_u2_n168 ) );
  NAND3_X1 u2_u11_u2_U100 (.A2( u2_u11_u2_n100 ) , .A1( u2_u11_u2_n104 ) , .A3( u2_u11_u2_n138 ) , .ZN( u2_u11_u2_n98 ) );
  OAI22_X1 u2_u11_u2_U11 (.B1( u2_u11_u2_n151 ) , .A2( u2_u11_u2_n152 ) , .A1( u2_u11_u2_n153 ) , .ZN( u2_u11_u2_n160 ) , .B2( u2_u11_u2_n168 ) );
  NOR3_X1 u2_u11_u2_U12 (.A1( u2_u11_u2_n150 ) , .ZN( u2_u11_u2_n151 ) , .A3( u2_u11_u2_n175 ) , .A2( u2_u11_u2_n188 ) );
  AOI21_X1 u2_u11_u2_U13 (.ZN( u2_u11_u2_n144 ) , .B2( u2_u11_u2_n155 ) , .A( u2_u11_u2_n172 ) , .B1( u2_u11_u2_n185 ) );
  AOI21_X1 u2_u11_u2_U14 (.B2( u2_u11_u2_n143 ) , .ZN( u2_u11_u2_n145 ) , .B1( u2_u11_u2_n152 ) , .A( u2_u11_u2_n171 ) );
  AOI21_X1 u2_u11_u2_U15 (.B2( u2_u11_u2_n120 ) , .B1( u2_u11_u2_n121 ) , .ZN( u2_u11_u2_n126 ) , .A( u2_u11_u2_n167 ) );
  INV_X1 u2_u11_u2_U16 (.A( u2_u11_u2_n156 ) , .ZN( u2_u11_u2_n171 ) );
  INV_X1 u2_u11_u2_U17 (.A( u2_u11_u2_n120 ) , .ZN( u2_u11_u2_n188 ) );
  NAND2_X1 u2_u11_u2_U18 (.A2( u2_u11_u2_n122 ) , .ZN( u2_u11_u2_n150 ) , .A1( u2_u11_u2_n152 ) );
  INV_X1 u2_u11_u2_U19 (.A( u2_u11_u2_n153 ) , .ZN( u2_u11_u2_n170 ) );
  INV_X1 u2_u11_u2_U20 (.A( u2_u11_u2_n137 ) , .ZN( u2_u11_u2_n173 ) );
  NAND2_X1 u2_u11_u2_U21 (.A1( u2_u11_u2_n132 ) , .A2( u2_u11_u2_n139 ) , .ZN( u2_u11_u2_n157 ) );
  INV_X1 u2_u11_u2_U22 (.A( u2_u11_u2_n113 ) , .ZN( u2_u11_u2_n178 ) );
  INV_X1 u2_u11_u2_U23 (.A( u2_u11_u2_n139 ) , .ZN( u2_u11_u2_n175 ) );
  INV_X1 u2_u11_u2_U24 (.A( u2_u11_u2_n155 ) , .ZN( u2_u11_u2_n181 ) );
  INV_X1 u2_u11_u2_U25 (.A( u2_u11_u2_n119 ) , .ZN( u2_u11_u2_n177 ) );
  INV_X1 u2_u11_u2_U26 (.A( u2_u11_u2_n116 ) , .ZN( u2_u11_u2_n180 ) );
  INV_X1 u2_u11_u2_U27 (.A( u2_u11_u2_n131 ) , .ZN( u2_u11_u2_n179 ) );
  INV_X1 u2_u11_u2_U28 (.A( u2_u11_u2_n154 ) , .ZN( u2_u11_u2_n176 ) );
  NAND2_X1 u2_u11_u2_U29 (.A2( u2_u11_u2_n116 ) , .A1( u2_u11_u2_n117 ) , .ZN( u2_u11_u2_n118 ) );
  NOR2_X1 u2_u11_u2_U3 (.ZN( u2_u11_u2_n121 ) , .A2( u2_u11_u2_n177 ) , .A1( u2_u11_u2_n180 ) );
  INV_X1 u2_u11_u2_U30 (.A( u2_u11_u2_n132 ) , .ZN( u2_u11_u2_n182 ) );
  INV_X1 u2_u11_u2_U31 (.A( u2_u11_u2_n158 ) , .ZN( u2_u11_u2_n183 ) );
  OAI21_X1 u2_u11_u2_U32 (.A( u2_u11_u2_n156 ) , .B1( u2_u11_u2_n157 ) , .ZN( u2_u11_u2_n158 ) , .B2( u2_u11_u2_n179 ) );
  NOR2_X1 u2_u11_u2_U33 (.ZN( u2_u11_u2_n156 ) , .A1( u2_u11_u2_n166 ) , .A2( u2_u11_u2_n169 ) );
  NOR2_X1 u2_u11_u2_U34 (.A2( u2_u11_u2_n114 ) , .ZN( u2_u11_u2_n137 ) , .A1( u2_u11_u2_n140 ) );
  NOR2_X1 u2_u11_u2_U35 (.A2( u2_u11_u2_n138 ) , .ZN( u2_u11_u2_n153 ) , .A1( u2_u11_u2_n156 ) );
  AOI211_X1 u2_u11_u2_U36 (.ZN( u2_u11_u2_n130 ) , .C1( u2_u11_u2_n138 ) , .C2( u2_u11_u2_n179 ) , .B( u2_u11_u2_n96 ) , .A( u2_u11_u2_n97 ) );
  OAI22_X1 u2_u11_u2_U37 (.B1( u2_u11_u2_n133 ) , .A2( u2_u11_u2_n137 ) , .A1( u2_u11_u2_n152 ) , .B2( u2_u11_u2_n168 ) , .ZN( u2_u11_u2_n97 ) );
  OAI221_X1 u2_u11_u2_U38 (.B1( u2_u11_u2_n113 ) , .C1( u2_u11_u2_n132 ) , .A( u2_u11_u2_n149 ) , .B2( u2_u11_u2_n171 ) , .C2( u2_u11_u2_n172 ) , .ZN( u2_u11_u2_n96 ) );
  OAI221_X1 u2_u11_u2_U39 (.A( u2_u11_u2_n115 ) , .C2( u2_u11_u2_n123 ) , .B2( u2_u11_u2_n143 ) , .B1( u2_u11_u2_n153 ) , .ZN( u2_u11_u2_n163 ) , .C1( u2_u11_u2_n168 ) );
  INV_X1 u2_u11_u2_U4 (.A( u2_u11_u2_n134 ) , .ZN( u2_u11_u2_n185 ) );
  OAI21_X1 u2_u11_u2_U40 (.A( u2_u11_u2_n114 ) , .ZN( u2_u11_u2_n115 ) , .B1( u2_u11_u2_n176 ) , .B2( u2_u11_u2_n178 ) );
  OAI221_X1 u2_u11_u2_U41 (.A( u2_u11_u2_n135 ) , .B2( u2_u11_u2_n136 ) , .B1( u2_u11_u2_n137 ) , .ZN( u2_u11_u2_n162 ) , .C2( u2_u11_u2_n167 ) , .C1( u2_u11_u2_n185 ) );
  AND3_X1 u2_u11_u2_U42 (.A3( u2_u11_u2_n131 ) , .A2( u2_u11_u2_n132 ) , .A1( u2_u11_u2_n133 ) , .ZN( u2_u11_u2_n136 ) );
  AOI22_X1 u2_u11_u2_U43 (.ZN( u2_u11_u2_n135 ) , .B1( u2_u11_u2_n140 ) , .A1( u2_u11_u2_n156 ) , .B2( u2_u11_u2_n180 ) , .A2( u2_u11_u2_n188 ) );
  AOI21_X1 u2_u11_u2_U44 (.ZN( u2_u11_u2_n149 ) , .B1( u2_u11_u2_n173 ) , .B2( u2_u11_u2_n188 ) , .A( u2_u11_u2_n95 ) );
  AND3_X1 u2_u11_u2_U45 (.A2( u2_u11_u2_n100 ) , .A1( u2_u11_u2_n104 ) , .A3( u2_u11_u2_n156 ) , .ZN( u2_u11_u2_n95 ) );
  OAI21_X1 u2_u11_u2_U46 (.A( u2_u11_u2_n101 ) , .B2( u2_u11_u2_n121 ) , .B1( u2_u11_u2_n153 ) , .ZN( u2_u11_u2_n164 ) );
  NAND2_X1 u2_u11_u2_U47 (.A2( u2_u11_u2_n100 ) , .A1( u2_u11_u2_n107 ) , .ZN( u2_u11_u2_n155 ) );
  NAND2_X1 u2_u11_u2_U48 (.A2( u2_u11_u2_n105 ) , .A1( u2_u11_u2_n108 ) , .ZN( u2_u11_u2_n143 ) );
  NAND2_X1 u2_u11_u2_U49 (.A1( u2_u11_u2_n104 ) , .A2( u2_u11_u2_n106 ) , .ZN( u2_u11_u2_n152 ) );
  INV_X1 u2_u11_u2_U5 (.A( u2_u11_u2_n150 ) , .ZN( u2_u11_u2_n184 ) );
  NAND2_X1 u2_u11_u2_U50 (.A1( u2_u11_u2_n100 ) , .A2( u2_u11_u2_n105 ) , .ZN( u2_u11_u2_n132 ) );
  INV_X1 u2_u11_u2_U51 (.A( u2_u11_u2_n140 ) , .ZN( u2_u11_u2_n168 ) );
  INV_X1 u2_u11_u2_U52 (.A( u2_u11_u2_n138 ) , .ZN( u2_u11_u2_n167 ) );
  OAI21_X1 u2_u11_u2_U53 (.A( u2_u11_u2_n141 ) , .B2( u2_u11_u2_n142 ) , .ZN( u2_u11_u2_n146 ) , .B1( u2_u11_u2_n153 ) );
  OAI21_X1 u2_u11_u2_U54 (.A( u2_u11_u2_n140 ) , .ZN( u2_u11_u2_n141 ) , .B1( u2_u11_u2_n176 ) , .B2( u2_u11_u2_n177 ) );
  NOR3_X1 u2_u11_u2_U55 (.ZN( u2_u11_u2_n142 ) , .A3( u2_u11_u2_n175 ) , .A2( u2_u11_u2_n178 ) , .A1( u2_u11_u2_n181 ) );
  NAND2_X1 u2_u11_u2_U56 (.A1( u2_u11_u2_n102 ) , .A2( u2_u11_u2_n106 ) , .ZN( u2_u11_u2_n113 ) );
  NAND2_X1 u2_u11_u2_U57 (.A1( u2_u11_u2_n106 ) , .A2( u2_u11_u2_n107 ) , .ZN( u2_u11_u2_n131 ) );
  NAND2_X1 u2_u11_u2_U58 (.A1( u2_u11_u2_n103 ) , .A2( u2_u11_u2_n107 ) , .ZN( u2_u11_u2_n139 ) );
  NAND2_X1 u2_u11_u2_U59 (.A1( u2_u11_u2_n103 ) , .A2( u2_u11_u2_n105 ) , .ZN( u2_u11_u2_n133 ) );
  NOR4_X1 u2_u11_u2_U6 (.A4( u2_u11_u2_n124 ) , .A3( u2_u11_u2_n125 ) , .A2( u2_u11_u2_n126 ) , .A1( u2_u11_u2_n127 ) , .ZN( u2_u11_u2_n128 ) );
  NAND2_X1 u2_u11_u2_U60 (.A1( u2_u11_u2_n102 ) , .A2( u2_u11_u2_n103 ) , .ZN( u2_u11_u2_n154 ) );
  NAND2_X1 u2_u11_u2_U61 (.A2( u2_u11_u2_n103 ) , .A1( u2_u11_u2_n104 ) , .ZN( u2_u11_u2_n119 ) );
  NAND2_X1 u2_u11_u2_U62 (.A2( u2_u11_u2_n107 ) , .A1( u2_u11_u2_n108 ) , .ZN( u2_u11_u2_n123 ) );
  NAND2_X1 u2_u11_u2_U63 (.A1( u2_u11_u2_n104 ) , .A2( u2_u11_u2_n108 ) , .ZN( u2_u11_u2_n122 ) );
  INV_X1 u2_u11_u2_U64 (.A( u2_u11_u2_n114 ) , .ZN( u2_u11_u2_n172 ) );
  NAND2_X1 u2_u11_u2_U65 (.A2( u2_u11_u2_n100 ) , .A1( u2_u11_u2_n102 ) , .ZN( u2_u11_u2_n116 ) );
  NAND2_X1 u2_u11_u2_U66 (.A1( u2_u11_u2_n102 ) , .A2( u2_u11_u2_n108 ) , .ZN( u2_u11_u2_n120 ) );
  NAND2_X1 u2_u11_u2_U67 (.A2( u2_u11_u2_n105 ) , .A1( u2_u11_u2_n106 ) , .ZN( u2_u11_u2_n117 ) );
  INV_X1 u2_u11_u2_U68 (.ZN( u2_u11_u2_n187 ) , .A( u2_u11_u2_n99 ) );
  OAI21_X1 u2_u11_u2_U69 (.B1( u2_u11_u2_n137 ) , .B2( u2_u11_u2_n143 ) , .A( u2_u11_u2_n98 ) , .ZN( u2_u11_u2_n99 ) );
  AOI21_X1 u2_u11_u2_U7 (.ZN( u2_u11_u2_n124 ) , .B1( u2_u11_u2_n131 ) , .B2( u2_u11_u2_n143 ) , .A( u2_u11_u2_n172 ) );
  NOR2_X1 u2_u11_u2_U70 (.A2( u2_u11_X_16 ) , .ZN( u2_u11_u2_n140 ) , .A1( u2_u11_u2_n166 ) );
  NOR2_X1 u2_u11_u2_U71 (.A2( u2_u11_X_13 ) , .A1( u2_u11_X_14 ) , .ZN( u2_u11_u2_n100 ) );
  NOR2_X1 u2_u11_u2_U72 (.A2( u2_u11_X_16 ) , .A1( u2_u11_X_17 ) , .ZN( u2_u11_u2_n138 ) );
  NOR2_X1 u2_u11_u2_U73 (.A2( u2_u11_X_15 ) , .A1( u2_u11_X_18 ) , .ZN( u2_u11_u2_n104 ) );
  NOR2_X1 u2_u11_u2_U74 (.A2( u2_u11_X_14 ) , .ZN( u2_u11_u2_n103 ) , .A1( u2_u11_u2_n174 ) );
  NOR2_X1 u2_u11_u2_U75 (.A2( u2_u11_X_15 ) , .ZN( u2_u11_u2_n102 ) , .A1( u2_u11_u2_n165 ) );
  NOR2_X1 u2_u11_u2_U76 (.A2( u2_u11_X_17 ) , .ZN( u2_u11_u2_n114 ) , .A1( u2_u11_u2_n169 ) );
  AND2_X1 u2_u11_u2_U77 (.A1( u2_u11_X_15 ) , .ZN( u2_u11_u2_n105 ) , .A2( u2_u11_u2_n165 ) );
  AND2_X1 u2_u11_u2_U78 (.A2( u2_u11_X_15 ) , .A1( u2_u11_X_18 ) , .ZN( u2_u11_u2_n107 ) );
  AND2_X1 u2_u11_u2_U79 (.A1( u2_u11_X_14 ) , .ZN( u2_u11_u2_n106 ) , .A2( u2_u11_u2_n174 ) );
  AOI21_X1 u2_u11_u2_U8 (.B2( u2_u11_u2_n119 ) , .ZN( u2_u11_u2_n127 ) , .A( u2_u11_u2_n137 ) , .B1( u2_u11_u2_n155 ) );
  AND2_X1 u2_u11_u2_U80 (.A1( u2_u11_X_13 ) , .A2( u2_u11_X_14 ) , .ZN( u2_u11_u2_n108 ) );
  INV_X1 u2_u11_u2_U81 (.A( u2_u11_X_16 ) , .ZN( u2_u11_u2_n169 ) );
  INV_X1 u2_u11_u2_U82 (.A( u2_u11_X_17 ) , .ZN( u2_u11_u2_n166 ) );
  INV_X1 u2_u11_u2_U83 (.A( u2_u11_X_13 ) , .ZN( u2_u11_u2_n174 ) );
  INV_X1 u2_u11_u2_U84 (.A( u2_u11_X_18 ) , .ZN( u2_u11_u2_n165 ) );
  NAND4_X1 u2_u11_u2_U85 (.ZN( u2_out11_30 ) , .A4( u2_u11_u2_n147 ) , .A3( u2_u11_u2_n148 ) , .A2( u2_u11_u2_n149 ) , .A1( u2_u11_u2_n187 ) );
  NOR3_X1 u2_u11_u2_U86 (.A3( u2_u11_u2_n144 ) , .A2( u2_u11_u2_n145 ) , .A1( u2_u11_u2_n146 ) , .ZN( u2_u11_u2_n147 ) );
  AOI21_X1 u2_u11_u2_U87 (.B2( u2_u11_u2_n138 ) , .ZN( u2_u11_u2_n148 ) , .A( u2_u11_u2_n162 ) , .B1( u2_u11_u2_n182 ) );
  NAND4_X1 u2_u11_u2_U88 (.ZN( u2_out11_24 ) , .A4( u2_u11_u2_n111 ) , .A3( u2_u11_u2_n112 ) , .A1( u2_u11_u2_n130 ) , .A2( u2_u11_u2_n187 ) );
  AOI221_X1 u2_u11_u2_U89 (.A( u2_u11_u2_n109 ) , .B1( u2_u11_u2_n110 ) , .ZN( u2_u11_u2_n111 ) , .C1( u2_u11_u2_n134 ) , .C2( u2_u11_u2_n170 ) , .B2( u2_u11_u2_n173 ) );
  AOI21_X1 u2_u11_u2_U9 (.B2( u2_u11_u2_n123 ) , .ZN( u2_u11_u2_n125 ) , .A( u2_u11_u2_n171 ) , .B1( u2_u11_u2_n184 ) );
  AOI21_X1 u2_u11_u2_U90 (.ZN( u2_u11_u2_n112 ) , .B2( u2_u11_u2_n156 ) , .A( u2_u11_u2_n164 ) , .B1( u2_u11_u2_n181 ) );
  NAND4_X1 u2_u11_u2_U91 (.ZN( u2_out11_16 ) , .A4( u2_u11_u2_n128 ) , .A3( u2_u11_u2_n129 ) , .A1( u2_u11_u2_n130 ) , .A2( u2_u11_u2_n186 ) );
  AOI22_X1 u2_u11_u2_U92 (.A2( u2_u11_u2_n118 ) , .ZN( u2_u11_u2_n129 ) , .A1( u2_u11_u2_n140 ) , .B1( u2_u11_u2_n157 ) , .B2( u2_u11_u2_n170 ) );
  INV_X1 u2_u11_u2_U93 (.A( u2_u11_u2_n163 ) , .ZN( u2_u11_u2_n186 ) );
  OR4_X1 u2_u11_u2_U94 (.ZN( u2_out11_6 ) , .A4( u2_u11_u2_n161 ) , .A3( u2_u11_u2_n162 ) , .A2( u2_u11_u2_n163 ) , .A1( u2_u11_u2_n164 ) );
  OR3_X1 u2_u11_u2_U95 (.A2( u2_u11_u2_n159 ) , .A1( u2_u11_u2_n160 ) , .ZN( u2_u11_u2_n161 ) , .A3( u2_u11_u2_n183 ) );
  AOI21_X1 u2_u11_u2_U96 (.B2( u2_u11_u2_n154 ) , .B1( u2_u11_u2_n155 ) , .ZN( u2_u11_u2_n159 ) , .A( u2_u11_u2_n167 ) );
  NAND3_X1 u2_u11_u2_U97 (.A2( u2_u11_u2_n117 ) , .A1( u2_u11_u2_n122 ) , .A3( u2_u11_u2_n123 ) , .ZN( u2_u11_u2_n134 ) );
  NAND3_X1 u2_u11_u2_U98 (.ZN( u2_u11_u2_n110 ) , .A2( u2_u11_u2_n131 ) , .A3( u2_u11_u2_n139 ) , .A1( u2_u11_u2_n154 ) );
  NAND3_X1 u2_u11_u2_U99 (.A2( u2_u11_u2_n100 ) , .ZN( u2_u11_u2_n101 ) , .A1( u2_u11_u2_n104 ) , .A3( u2_u11_u2_n114 ) );
  XOR2_X1 u2_u13_U20 (.B( u2_K14_36 ) , .A( u2_R12_25 ) , .Z( u2_u13_X_36 ) );
  XOR2_X1 u2_u13_U21 (.B( u2_K14_35 ) , .A( u2_R12_24 ) , .Z( u2_u13_X_35 ) );
  XOR2_X1 u2_u13_U22 (.B( u2_K14_34 ) , .A( u2_R12_23 ) , .Z( u2_u13_X_34 ) );
  XOR2_X1 u2_u13_U23 (.B( u2_K14_33 ) , .A( u2_R12_22 ) , .Z( u2_u13_X_33 ) );
  XOR2_X1 u2_u13_U24 (.B( u2_K14_32 ) , .A( u2_R12_21 ) , .Z( u2_u13_X_32 ) );
  XOR2_X1 u2_u13_U25 (.B( u2_K14_31 ) , .A( u2_R12_20 ) , .Z( u2_u13_X_31 ) );
  XOR2_X1 u2_u13_U26 (.B( u2_K14_30 ) , .A( u2_R12_21 ) , .Z( u2_u13_X_30 ) );
  XOR2_X1 u2_u13_U28 (.B( u2_K14_29 ) , .A( u2_R12_20 ) , .Z( u2_u13_X_29 ) );
  XOR2_X1 u2_u13_U29 (.B( u2_K14_28 ) , .A( u2_R12_19 ) , .Z( u2_u13_X_28 ) );
  XOR2_X1 u2_u13_U30 (.B( u2_K14_27 ) , .A( u2_R12_18 ) , .Z( u2_u13_X_27 ) );
  XOR2_X1 u2_u13_U31 (.B( u2_K14_26 ) , .A( u2_R12_17 ) , .Z( u2_u13_X_26 ) );
  XOR2_X1 u2_u13_U32 (.B( u2_K14_25 ) , .A( u2_R12_16 ) , .Z( u2_u13_X_25 ) );
  AOI21_X1 u2_u13_u4_U10 (.ZN( u2_u13_u4_n106 ) , .B2( u2_u13_u4_n146 ) , .B1( u2_u13_u4_n158 ) , .A( u2_u13_u4_n170 ) );
  AOI21_X1 u2_u13_u4_U11 (.ZN( u2_u13_u4_n108 ) , .B2( u2_u13_u4_n134 ) , .B1( u2_u13_u4_n155 ) , .A( u2_u13_u4_n156 ) );
  AOI21_X1 u2_u13_u4_U12 (.ZN( u2_u13_u4_n109 ) , .A( u2_u13_u4_n153 ) , .B1( u2_u13_u4_n159 ) , .B2( u2_u13_u4_n184 ) );
  AOI211_X1 u2_u13_u4_U13 (.B( u2_u13_u4_n136 ) , .A( u2_u13_u4_n137 ) , .C2( u2_u13_u4_n138 ) , .ZN( u2_u13_u4_n139 ) , .C1( u2_u13_u4_n182 ) );
  OAI22_X1 u2_u13_u4_U14 (.B2( u2_u13_u4_n135 ) , .ZN( u2_u13_u4_n137 ) , .B1( u2_u13_u4_n153 ) , .A1( u2_u13_u4_n155 ) , .A2( u2_u13_u4_n171 ) );
  AND3_X1 u2_u13_u4_U15 (.A2( u2_u13_u4_n134 ) , .ZN( u2_u13_u4_n135 ) , .A3( u2_u13_u4_n145 ) , .A1( u2_u13_u4_n157 ) );
  NAND2_X1 u2_u13_u4_U16 (.ZN( u2_u13_u4_n132 ) , .A2( u2_u13_u4_n170 ) , .A1( u2_u13_u4_n173 ) );
  AOI21_X1 u2_u13_u4_U17 (.B2( u2_u13_u4_n160 ) , .B1( u2_u13_u4_n161 ) , .ZN( u2_u13_u4_n162 ) , .A( u2_u13_u4_n170 ) );
  AOI21_X1 u2_u13_u4_U18 (.ZN( u2_u13_u4_n107 ) , .B2( u2_u13_u4_n143 ) , .A( u2_u13_u4_n174 ) , .B1( u2_u13_u4_n184 ) );
  AOI21_X1 u2_u13_u4_U19 (.B2( u2_u13_u4_n158 ) , .B1( u2_u13_u4_n159 ) , .ZN( u2_u13_u4_n163 ) , .A( u2_u13_u4_n174 ) );
  AOI21_X1 u2_u13_u4_U20 (.A( u2_u13_u4_n153 ) , .B2( u2_u13_u4_n154 ) , .B1( u2_u13_u4_n155 ) , .ZN( u2_u13_u4_n165 ) );
  AOI21_X1 u2_u13_u4_U21 (.A( u2_u13_u4_n156 ) , .B2( u2_u13_u4_n157 ) , .ZN( u2_u13_u4_n164 ) , .B1( u2_u13_u4_n184 ) );
  INV_X1 u2_u13_u4_U22 (.A( u2_u13_u4_n138 ) , .ZN( u2_u13_u4_n170 ) );
  AND2_X1 u2_u13_u4_U23 (.A2( u2_u13_u4_n120 ) , .ZN( u2_u13_u4_n155 ) , .A1( u2_u13_u4_n160 ) );
  INV_X1 u2_u13_u4_U24 (.A( u2_u13_u4_n156 ) , .ZN( u2_u13_u4_n175 ) );
  NAND2_X1 u2_u13_u4_U25 (.A2( u2_u13_u4_n118 ) , .ZN( u2_u13_u4_n131 ) , .A1( u2_u13_u4_n147 ) );
  NAND2_X1 u2_u13_u4_U26 (.A1( u2_u13_u4_n119 ) , .A2( u2_u13_u4_n120 ) , .ZN( u2_u13_u4_n130 ) );
  NAND2_X1 u2_u13_u4_U27 (.ZN( u2_u13_u4_n117 ) , .A2( u2_u13_u4_n118 ) , .A1( u2_u13_u4_n148 ) );
  NAND2_X1 u2_u13_u4_U28 (.ZN( u2_u13_u4_n129 ) , .A1( u2_u13_u4_n134 ) , .A2( u2_u13_u4_n148 ) );
  AND3_X1 u2_u13_u4_U29 (.A1( u2_u13_u4_n119 ) , .A2( u2_u13_u4_n143 ) , .A3( u2_u13_u4_n154 ) , .ZN( u2_u13_u4_n161 ) );
  NOR2_X1 u2_u13_u4_U3 (.ZN( u2_u13_u4_n121 ) , .A1( u2_u13_u4_n181 ) , .A2( u2_u13_u4_n182 ) );
  AND2_X1 u2_u13_u4_U30 (.A1( u2_u13_u4_n145 ) , .A2( u2_u13_u4_n147 ) , .ZN( u2_u13_u4_n159 ) );
  OR3_X1 u2_u13_u4_U31 (.A3( u2_u13_u4_n114 ) , .A2( u2_u13_u4_n115 ) , .A1( u2_u13_u4_n116 ) , .ZN( u2_u13_u4_n136 ) );
  AOI21_X1 u2_u13_u4_U32 (.A( u2_u13_u4_n113 ) , .ZN( u2_u13_u4_n116 ) , .B2( u2_u13_u4_n173 ) , .B1( u2_u13_u4_n174 ) );
  AOI21_X1 u2_u13_u4_U33 (.ZN( u2_u13_u4_n115 ) , .B2( u2_u13_u4_n145 ) , .B1( u2_u13_u4_n146 ) , .A( u2_u13_u4_n156 ) );
  OAI22_X1 u2_u13_u4_U34 (.ZN( u2_u13_u4_n114 ) , .A2( u2_u13_u4_n121 ) , .B1( u2_u13_u4_n160 ) , .B2( u2_u13_u4_n170 ) , .A1( u2_u13_u4_n171 ) );
  INV_X1 u2_u13_u4_U35 (.A( u2_u13_u4_n158 ) , .ZN( u2_u13_u4_n182 ) );
  INV_X1 u2_u13_u4_U36 (.ZN( u2_u13_u4_n181 ) , .A( u2_u13_u4_n96 ) );
  INV_X1 u2_u13_u4_U37 (.A( u2_u13_u4_n144 ) , .ZN( u2_u13_u4_n179 ) );
  INV_X1 u2_u13_u4_U38 (.A( u2_u13_u4_n157 ) , .ZN( u2_u13_u4_n178 ) );
  NAND2_X1 u2_u13_u4_U39 (.A2( u2_u13_u4_n154 ) , .A1( u2_u13_u4_n96 ) , .ZN( u2_u13_u4_n97 ) );
  INV_X1 u2_u13_u4_U4 (.A( u2_u13_u4_n117 ) , .ZN( u2_u13_u4_n184 ) );
  INV_X1 u2_u13_u4_U40 (.A( u2_u13_u4_n143 ) , .ZN( u2_u13_u4_n183 ) );
  NOR2_X1 u2_u13_u4_U41 (.ZN( u2_u13_u4_n138 ) , .A1( u2_u13_u4_n168 ) , .A2( u2_u13_u4_n169 ) );
  NOR2_X1 u2_u13_u4_U42 (.A1( u2_u13_u4_n150 ) , .A2( u2_u13_u4_n152 ) , .ZN( u2_u13_u4_n153 ) );
  NOR2_X1 u2_u13_u4_U43 (.A2( u2_u13_u4_n128 ) , .A1( u2_u13_u4_n138 ) , .ZN( u2_u13_u4_n156 ) );
  AOI22_X1 u2_u13_u4_U44 (.B2( u2_u13_u4_n122 ) , .A1( u2_u13_u4_n123 ) , .ZN( u2_u13_u4_n124 ) , .B1( u2_u13_u4_n128 ) , .A2( u2_u13_u4_n172 ) );
  NAND2_X1 u2_u13_u4_U45 (.A2( u2_u13_u4_n120 ) , .ZN( u2_u13_u4_n123 ) , .A1( u2_u13_u4_n161 ) );
  INV_X1 u2_u13_u4_U46 (.A( u2_u13_u4_n153 ) , .ZN( u2_u13_u4_n172 ) );
  AOI22_X1 u2_u13_u4_U47 (.B2( u2_u13_u4_n132 ) , .A2( u2_u13_u4_n133 ) , .ZN( u2_u13_u4_n140 ) , .A1( u2_u13_u4_n150 ) , .B1( u2_u13_u4_n179 ) );
  NAND2_X1 u2_u13_u4_U48 (.ZN( u2_u13_u4_n133 ) , .A2( u2_u13_u4_n146 ) , .A1( u2_u13_u4_n154 ) );
  NAND2_X1 u2_u13_u4_U49 (.A1( u2_u13_u4_n103 ) , .ZN( u2_u13_u4_n154 ) , .A2( u2_u13_u4_n98 ) );
  INV_X1 u2_u13_u4_U5 (.ZN( u2_u13_u4_n186 ) , .A( u2_u13_u4_n95 ) );
  NAND2_X1 u2_u13_u4_U50 (.A1( u2_u13_u4_n101 ) , .ZN( u2_u13_u4_n158 ) , .A2( u2_u13_u4_n99 ) );
  AOI21_X1 u2_u13_u4_U51 (.ZN( u2_u13_u4_n127 ) , .A( u2_u13_u4_n136 ) , .B2( u2_u13_u4_n150 ) , .B1( u2_u13_u4_n180 ) );
  INV_X1 u2_u13_u4_U52 (.A( u2_u13_u4_n160 ) , .ZN( u2_u13_u4_n180 ) );
  NAND2_X1 u2_u13_u4_U53 (.A2( u2_u13_u4_n104 ) , .A1( u2_u13_u4_n105 ) , .ZN( u2_u13_u4_n146 ) );
  NAND2_X1 u2_u13_u4_U54 (.A2( u2_u13_u4_n101 ) , .A1( u2_u13_u4_n102 ) , .ZN( u2_u13_u4_n160 ) );
  NAND2_X1 u2_u13_u4_U55 (.ZN( u2_u13_u4_n134 ) , .A1( u2_u13_u4_n98 ) , .A2( u2_u13_u4_n99 ) );
  NAND2_X1 u2_u13_u4_U56 (.A1( u2_u13_u4_n103 ) , .A2( u2_u13_u4_n104 ) , .ZN( u2_u13_u4_n143 ) );
  NAND2_X1 u2_u13_u4_U57 (.A2( u2_u13_u4_n105 ) , .ZN( u2_u13_u4_n145 ) , .A1( u2_u13_u4_n98 ) );
  NAND2_X1 u2_u13_u4_U58 (.A1( u2_u13_u4_n100 ) , .A2( u2_u13_u4_n105 ) , .ZN( u2_u13_u4_n120 ) );
  NAND2_X1 u2_u13_u4_U59 (.A1( u2_u13_u4_n102 ) , .A2( u2_u13_u4_n104 ) , .ZN( u2_u13_u4_n148 ) );
  OAI221_X1 u2_u13_u4_U6 (.C1( u2_u13_u4_n134 ) , .B1( u2_u13_u4_n158 ) , .B2( u2_u13_u4_n171 ) , .C2( u2_u13_u4_n173 ) , .A( u2_u13_u4_n94 ) , .ZN( u2_u13_u4_n95 ) );
  NAND2_X1 u2_u13_u4_U60 (.A2( u2_u13_u4_n100 ) , .A1( u2_u13_u4_n103 ) , .ZN( u2_u13_u4_n157 ) );
  INV_X1 u2_u13_u4_U61 (.A( u2_u13_u4_n150 ) , .ZN( u2_u13_u4_n173 ) );
  INV_X1 u2_u13_u4_U62 (.A( u2_u13_u4_n152 ) , .ZN( u2_u13_u4_n171 ) );
  NAND2_X1 u2_u13_u4_U63 (.A1( u2_u13_u4_n100 ) , .ZN( u2_u13_u4_n118 ) , .A2( u2_u13_u4_n99 ) );
  NAND2_X1 u2_u13_u4_U64 (.A2( u2_u13_u4_n100 ) , .A1( u2_u13_u4_n102 ) , .ZN( u2_u13_u4_n144 ) );
  NAND2_X1 u2_u13_u4_U65 (.A2( u2_u13_u4_n101 ) , .A1( u2_u13_u4_n105 ) , .ZN( u2_u13_u4_n96 ) );
  INV_X1 u2_u13_u4_U66 (.A( u2_u13_u4_n128 ) , .ZN( u2_u13_u4_n174 ) );
  NAND2_X1 u2_u13_u4_U67 (.A2( u2_u13_u4_n102 ) , .ZN( u2_u13_u4_n119 ) , .A1( u2_u13_u4_n98 ) );
  NAND2_X1 u2_u13_u4_U68 (.A2( u2_u13_u4_n101 ) , .A1( u2_u13_u4_n103 ) , .ZN( u2_u13_u4_n147 ) );
  NAND2_X1 u2_u13_u4_U69 (.A2( u2_u13_u4_n104 ) , .ZN( u2_u13_u4_n113 ) , .A1( u2_u13_u4_n99 ) );
  AOI222_X1 u2_u13_u4_U7 (.B2( u2_u13_u4_n132 ) , .A1( u2_u13_u4_n138 ) , .C2( u2_u13_u4_n175 ) , .A2( u2_u13_u4_n179 ) , .C1( u2_u13_u4_n181 ) , .B1( u2_u13_u4_n185 ) , .ZN( u2_u13_u4_n94 ) );
  NOR2_X1 u2_u13_u4_U70 (.A2( u2_u13_X_28 ) , .ZN( u2_u13_u4_n150 ) , .A1( u2_u13_u4_n168 ) );
  NOR2_X1 u2_u13_u4_U71 (.A2( u2_u13_X_29 ) , .ZN( u2_u13_u4_n152 ) , .A1( u2_u13_u4_n169 ) );
  NOR2_X1 u2_u13_u4_U72 (.A2( u2_u13_X_30 ) , .ZN( u2_u13_u4_n105 ) , .A1( u2_u13_u4_n176 ) );
  NOR2_X1 u2_u13_u4_U73 (.A2( u2_u13_X_26 ) , .ZN( u2_u13_u4_n100 ) , .A1( u2_u13_u4_n177 ) );
  NOR2_X1 u2_u13_u4_U74 (.A2( u2_u13_X_28 ) , .A1( u2_u13_X_29 ) , .ZN( u2_u13_u4_n128 ) );
  NOR2_X1 u2_u13_u4_U75 (.A2( u2_u13_X_27 ) , .A1( u2_u13_X_30 ) , .ZN( u2_u13_u4_n102 ) );
  NOR2_X1 u2_u13_u4_U76 (.A2( u2_u13_X_25 ) , .A1( u2_u13_X_26 ) , .ZN( u2_u13_u4_n98 ) );
  AND2_X1 u2_u13_u4_U77 (.A2( u2_u13_X_25 ) , .A1( u2_u13_X_26 ) , .ZN( u2_u13_u4_n104 ) );
  AND2_X1 u2_u13_u4_U78 (.A1( u2_u13_X_30 ) , .A2( u2_u13_u4_n176 ) , .ZN( u2_u13_u4_n99 ) );
  AND2_X1 u2_u13_u4_U79 (.A1( u2_u13_X_26 ) , .ZN( u2_u13_u4_n101 ) , .A2( u2_u13_u4_n177 ) );
  INV_X1 u2_u13_u4_U8 (.A( u2_u13_u4_n113 ) , .ZN( u2_u13_u4_n185 ) );
  AND2_X1 u2_u13_u4_U80 (.A1( u2_u13_X_27 ) , .A2( u2_u13_X_30 ) , .ZN( u2_u13_u4_n103 ) );
  INV_X1 u2_u13_u4_U81 (.A( u2_u13_X_28 ) , .ZN( u2_u13_u4_n169 ) );
  INV_X1 u2_u13_u4_U82 (.A( u2_u13_X_29 ) , .ZN( u2_u13_u4_n168 ) );
  INV_X1 u2_u13_u4_U83 (.A( u2_u13_X_25 ) , .ZN( u2_u13_u4_n177 ) );
  INV_X1 u2_u13_u4_U84 (.A( u2_u13_X_27 ) , .ZN( u2_u13_u4_n176 ) );
  NAND4_X1 u2_u13_u4_U85 (.ZN( u2_out13_25 ) , .A4( u2_u13_u4_n139 ) , .A3( u2_u13_u4_n140 ) , .A2( u2_u13_u4_n141 ) , .A1( u2_u13_u4_n142 ) );
  OAI21_X1 u2_u13_u4_U86 (.A( u2_u13_u4_n128 ) , .B2( u2_u13_u4_n129 ) , .B1( u2_u13_u4_n130 ) , .ZN( u2_u13_u4_n142 ) );
  OAI21_X1 u2_u13_u4_U87 (.B2( u2_u13_u4_n131 ) , .ZN( u2_u13_u4_n141 ) , .A( u2_u13_u4_n175 ) , .B1( u2_u13_u4_n183 ) );
  NAND4_X1 u2_u13_u4_U88 (.ZN( u2_out13_14 ) , .A4( u2_u13_u4_n124 ) , .A3( u2_u13_u4_n125 ) , .A2( u2_u13_u4_n126 ) , .A1( u2_u13_u4_n127 ) );
  AOI22_X1 u2_u13_u4_U89 (.B2( u2_u13_u4_n117 ) , .ZN( u2_u13_u4_n126 ) , .A1( u2_u13_u4_n129 ) , .B1( u2_u13_u4_n152 ) , .A2( u2_u13_u4_n175 ) );
  NOR4_X1 u2_u13_u4_U9 (.A4( u2_u13_u4_n106 ) , .A3( u2_u13_u4_n107 ) , .A2( u2_u13_u4_n108 ) , .A1( u2_u13_u4_n109 ) , .ZN( u2_u13_u4_n110 ) );
  AOI22_X1 u2_u13_u4_U90 (.ZN( u2_u13_u4_n125 ) , .B2( u2_u13_u4_n131 ) , .A2( u2_u13_u4_n132 ) , .B1( u2_u13_u4_n138 ) , .A1( u2_u13_u4_n178 ) );
  NAND4_X1 u2_u13_u4_U91 (.ZN( u2_out13_8 ) , .A4( u2_u13_u4_n110 ) , .A3( u2_u13_u4_n111 ) , .A2( u2_u13_u4_n112 ) , .A1( u2_u13_u4_n186 ) );
  NAND2_X1 u2_u13_u4_U92 (.ZN( u2_u13_u4_n112 ) , .A2( u2_u13_u4_n130 ) , .A1( u2_u13_u4_n150 ) );
  AOI22_X1 u2_u13_u4_U93 (.ZN( u2_u13_u4_n111 ) , .B2( u2_u13_u4_n132 ) , .A1( u2_u13_u4_n152 ) , .B1( u2_u13_u4_n178 ) , .A2( u2_u13_u4_n97 ) );
  AOI22_X1 u2_u13_u4_U94 (.B2( u2_u13_u4_n149 ) , .B1( u2_u13_u4_n150 ) , .A2( u2_u13_u4_n151 ) , .A1( u2_u13_u4_n152 ) , .ZN( u2_u13_u4_n167 ) );
  NOR4_X1 u2_u13_u4_U95 (.A4( u2_u13_u4_n162 ) , .A3( u2_u13_u4_n163 ) , .A2( u2_u13_u4_n164 ) , .A1( u2_u13_u4_n165 ) , .ZN( u2_u13_u4_n166 ) );
  NAND3_X1 u2_u13_u4_U96 (.ZN( u2_out13_3 ) , .A3( u2_u13_u4_n166 ) , .A1( u2_u13_u4_n167 ) , .A2( u2_u13_u4_n186 ) );
  NAND3_X1 u2_u13_u4_U97 (.A3( u2_u13_u4_n146 ) , .A2( u2_u13_u4_n147 ) , .A1( u2_u13_u4_n148 ) , .ZN( u2_u13_u4_n149 ) );
  NAND3_X1 u2_u13_u4_U98 (.A3( u2_u13_u4_n143 ) , .A2( u2_u13_u4_n144 ) , .A1( u2_u13_u4_n145 ) , .ZN( u2_u13_u4_n151 ) );
  NAND3_X1 u2_u13_u4_U99 (.A3( u2_u13_u4_n121 ) , .ZN( u2_u13_u4_n122 ) , .A2( u2_u13_u4_n144 ) , .A1( u2_u13_u4_n154 ) );
  INV_X1 u2_u13_u5_U10 (.A( u2_u13_u5_n121 ) , .ZN( u2_u13_u5_n177 ) );
  NOR3_X1 u2_u13_u5_U100 (.A3( u2_u13_u5_n141 ) , .A1( u2_u13_u5_n142 ) , .ZN( u2_u13_u5_n143 ) , .A2( u2_u13_u5_n191 ) );
  NAND4_X1 u2_u13_u5_U101 (.ZN( u2_out13_4 ) , .A4( u2_u13_u5_n112 ) , .A2( u2_u13_u5_n113 ) , .A1( u2_u13_u5_n114 ) , .A3( u2_u13_u5_n195 ) );
  AOI211_X1 u2_u13_u5_U102 (.A( u2_u13_u5_n110 ) , .C1( u2_u13_u5_n111 ) , .ZN( u2_u13_u5_n112 ) , .B( u2_u13_u5_n118 ) , .C2( u2_u13_u5_n177 ) );
  AOI222_X1 u2_u13_u5_U103 (.ZN( u2_u13_u5_n113 ) , .A1( u2_u13_u5_n131 ) , .C1( u2_u13_u5_n148 ) , .B2( u2_u13_u5_n174 ) , .C2( u2_u13_u5_n178 ) , .A2( u2_u13_u5_n179 ) , .B1( u2_u13_u5_n99 ) );
  NAND3_X1 u2_u13_u5_U104 (.A2( u2_u13_u5_n154 ) , .A3( u2_u13_u5_n158 ) , .A1( u2_u13_u5_n161 ) , .ZN( u2_u13_u5_n99 ) );
  NOR2_X1 u2_u13_u5_U11 (.ZN( u2_u13_u5_n160 ) , .A2( u2_u13_u5_n173 ) , .A1( u2_u13_u5_n177 ) );
  INV_X1 u2_u13_u5_U12 (.A( u2_u13_u5_n150 ) , .ZN( u2_u13_u5_n174 ) );
  AOI21_X1 u2_u13_u5_U13 (.A( u2_u13_u5_n160 ) , .B2( u2_u13_u5_n161 ) , .ZN( u2_u13_u5_n162 ) , .B1( u2_u13_u5_n192 ) );
  INV_X1 u2_u13_u5_U14 (.A( u2_u13_u5_n159 ) , .ZN( u2_u13_u5_n192 ) );
  AOI21_X1 u2_u13_u5_U15 (.A( u2_u13_u5_n156 ) , .B2( u2_u13_u5_n157 ) , .B1( u2_u13_u5_n158 ) , .ZN( u2_u13_u5_n163 ) );
  AOI21_X1 u2_u13_u5_U16 (.B2( u2_u13_u5_n139 ) , .B1( u2_u13_u5_n140 ) , .ZN( u2_u13_u5_n141 ) , .A( u2_u13_u5_n150 ) );
  OAI21_X1 u2_u13_u5_U17 (.A( u2_u13_u5_n133 ) , .B2( u2_u13_u5_n134 ) , .B1( u2_u13_u5_n135 ) , .ZN( u2_u13_u5_n142 ) );
  OAI21_X1 u2_u13_u5_U18 (.ZN( u2_u13_u5_n133 ) , .B2( u2_u13_u5_n147 ) , .A( u2_u13_u5_n173 ) , .B1( u2_u13_u5_n188 ) );
  NAND2_X1 u2_u13_u5_U19 (.A2( u2_u13_u5_n119 ) , .A1( u2_u13_u5_n123 ) , .ZN( u2_u13_u5_n137 ) );
  INV_X1 u2_u13_u5_U20 (.A( u2_u13_u5_n155 ) , .ZN( u2_u13_u5_n194 ) );
  NAND2_X1 u2_u13_u5_U21 (.A1( u2_u13_u5_n121 ) , .ZN( u2_u13_u5_n132 ) , .A2( u2_u13_u5_n172 ) );
  NAND2_X1 u2_u13_u5_U22 (.A2( u2_u13_u5_n122 ) , .ZN( u2_u13_u5_n136 ) , .A1( u2_u13_u5_n154 ) );
  NAND2_X1 u2_u13_u5_U23 (.A2( u2_u13_u5_n119 ) , .A1( u2_u13_u5_n120 ) , .ZN( u2_u13_u5_n159 ) );
  INV_X1 u2_u13_u5_U24 (.A( u2_u13_u5_n156 ) , .ZN( u2_u13_u5_n175 ) );
  INV_X1 u2_u13_u5_U25 (.A( u2_u13_u5_n158 ) , .ZN( u2_u13_u5_n188 ) );
  INV_X1 u2_u13_u5_U26 (.A( u2_u13_u5_n152 ) , .ZN( u2_u13_u5_n179 ) );
  INV_X1 u2_u13_u5_U27 (.A( u2_u13_u5_n140 ) , .ZN( u2_u13_u5_n182 ) );
  INV_X1 u2_u13_u5_U28 (.A( u2_u13_u5_n151 ) , .ZN( u2_u13_u5_n183 ) );
  INV_X1 u2_u13_u5_U29 (.A( u2_u13_u5_n123 ) , .ZN( u2_u13_u5_n185 ) );
  NOR2_X1 u2_u13_u5_U3 (.ZN( u2_u13_u5_n134 ) , .A1( u2_u13_u5_n183 ) , .A2( u2_u13_u5_n190 ) );
  INV_X1 u2_u13_u5_U30 (.A( u2_u13_u5_n161 ) , .ZN( u2_u13_u5_n184 ) );
  INV_X1 u2_u13_u5_U31 (.A( u2_u13_u5_n139 ) , .ZN( u2_u13_u5_n189 ) );
  INV_X1 u2_u13_u5_U32 (.A( u2_u13_u5_n157 ) , .ZN( u2_u13_u5_n190 ) );
  INV_X1 u2_u13_u5_U33 (.A( u2_u13_u5_n120 ) , .ZN( u2_u13_u5_n193 ) );
  NAND2_X1 u2_u13_u5_U34 (.ZN( u2_u13_u5_n111 ) , .A1( u2_u13_u5_n140 ) , .A2( u2_u13_u5_n155 ) );
  NOR2_X1 u2_u13_u5_U35 (.ZN( u2_u13_u5_n100 ) , .A1( u2_u13_u5_n170 ) , .A2( u2_u13_u5_n180 ) );
  INV_X1 u2_u13_u5_U36 (.A( u2_u13_u5_n117 ) , .ZN( u2_u13_u5_n196 ) );
  OAI221_X1 u2_u13_u5_U37 (.A( u2_u13_u5_n116 ) , .ZN( u2_u13_u5_n117 ) , .B2( u2_u13_u5_n119 ) , .C1( u2_u13_u5_n153 ) , .C2( u2_u13_u5_n158 ) , .B1( u2_u13_u5_n172 ) );
  AOI222_X1 u2_u13_u5_U38 (.ZN( u2_u13_u5_n116 ) , .B2( u2_u13_u5_n145 ) , .C1( u2_u13_u5_n148 ) , .A2( u2_u13_u5_n174 ) , .C2( u2_u13_u5_n177 ) , .B1( u2_u13_u5_n187 ) , .A1( u2_u13_u5_n193 ) );
  INV_X1 u2_u13_u5_U39 (.A( u2_u13_u5_n115 ) , .ZN( u2_u13_u5_n187 ) );
  INV_X1 u2_u13_u5_U4 (.A( u2_u13_u5_n138 ) , .ZN( u2_u13_u5_n191 ) );
  AOI22_X1 u2_u13_u5_U40 (.B2( u2_u13_u5_n131 ) , .A2( u2_u13_u5_n146 ) , .ZN( u2_u13_u5_n169 ) , .B1( u2_u13_u5_n174 ) , .A1( u2_u13_u5_n185 ) );
  NOR2_X1 u2_u13_u5_U41 (.A1( u2_u13_u5_n146 ) , .ZN( u2_u13_u5_n150 ) , .A2( u2_u13_u5_n173 ) );
  AOI21_X1 u2_u13_u5_U42 (.A( u2_u13_u5_n118 ) , .B2( u2_u13_u5_n145 ) , .ZN( u2_u13_u5_n168 ) , .B1( u2_u13_u5_n186 ) );
  INV_X1 u2_u13_u5_U43 (.A( u2_u13_u5_n122 ) , .ZN( u2_u13_u5_n186 ) );
  NOR2_X1 u2_u13_u5_U44 (.A1( u2_u13_u5_n146 ) , .ZN( u2_u13_u5_n152 ) , .A2( u2_u13_u5_n176 ) );
  NOR2_X1 u2_u13_u5_U45 (.A1( u2_u13_u5_n115 ) , .ZN( u2_u13_u5_n118 ) , .A2( u2_u13_u5_n153 ) );
  NOR2_X1 u2_u13_u5_U46 (.A2( u2_u13_u5_n145 ) , .ZN( u2_u13_u5_n156 ) , .A1( u2_u13_u5_n174 ) );
  NOR2_X1 u2_u13_u5_U47 (.ZN( u2_u13_u5_n121 ) , .A2( u2_u13_u5_n145 ) , .A1( u2_u13_u5_n176 ) );
  AOI22_X1 u2_u13_u5_U48 (.ZN( u2_u13_u5_n114 ) , .A2( u2_u13_u5_n137 ) , .A1( u2_u13_u5_n145 ) , .B2( u2_u13_u5_n175 ) , .B1( u2_u13_u5_n193 ) );
  OAI211_X1 u2_u13_u5_U49 (.B( u2_u13_u5_n124 ) , .A( u2_u13_u5_n125 ) , .C2( u2_u13_u5_n126 ) , .C1( u2_u13_u5_n127 ) , .ZN( u2_u13_u5_n128 ) );
  OAI21_X1 u2_u13_u5_U5 (.B2( u2_u13_u5_n136 ) , .B1( u2_u13_u5_n137 ) , .ZN( u2_u13_u5_n138 ) , .A( u2_u13_u5_n177 ) );
  NOR3_X1 u2_u13_u5_U50 (.ZN( u2_u13_u5_n127 ) , .A1( u2_u13_u5_n136 ) , .A3( u2_u13_u5_n148 ) , .A2( u2_u13_u5_n182 ) );
  OAI21_X1 u2_u13_u5_U51 (.ZN( u2_u13_u5_n124 ) , .A( u2_u13_u5_n177 ) , .B2( u2_u13_u5_n183 ) , .B1( u2_u13_u5_n189 ) );
  OAI21_X1 u2_u13_u5_U52 (.ZN( u2_u13_u5_n125 ) , .A( u2_u13_u5_n174 ) , .B2( u2_u13_u5_n185 ) , .B1( u2_u13_u5_n190 ) );
  AOI21_X1 u2_u13_u5_U53 (.A( u2_u13_u5_n153 ) , .B2( u2_u13_u5_n154 ) , .B1( u2_u13_u5_n155 ) , .ZN( u2_u13_u5_n164 ) );
  AOI21_X1 u2_u13_u5_U54 (.ZN( u2_u13_u5_n110 ) , .B1( u2_u13_u5_n122 ) , .B2( u2_u13_u5_n139 ) , .A( u2_u13_u5_n153 ) );
  INV_X1 u2_u13_u5_U55 (.A( u2_u13_u5_n153 ) , .ZN( u2_u13_u5_n176 ) );
  INV_X1 u2_u13_u5_U56 (.A( u2_u13_u5_n126 ) , .ZN( u2_u13_u5_n173 ) );
  AND2_X1 u2_u13_u5_U57 (.A2( u2_u13_u5_n104 ) , .A1( u2_u13_u5_n107 ) , .ZN( u2_u13_u5_n147 ) );
  AND2_X1 u2_u13_u5_U58 (.A2( u2_u13_u5_n104 ) , .A1( u2_u13_u5_n108 ) , .ZN( u2_u13_u5_n148 ) );
  NAND2_X1 u2_u13_u5_U59 (.A1( u2_u13_u5_n105 ) , .A2( u2_u13_u5_n106 ) , .ZN( u2_u13_u5_n158 ) );
  INV_X1 u2_u13_u5_U6 (.A( u2_u13_u5_n135 ) , .ZN( u2_u13_u5_n178 ) );
  NAND2_X1 u2_u13_u5_U60 (.A2( u2_u13_u5_n108 ) , .A1( u2_u13_u5_n109 ) , .ZN( u2_u13_u5_n139 ) );
  NAND2_X1 u2_u13_u5_U61 (.A1( u2_u13_u5_n106 ) , .A2( u2_u13_u5_n108 ) , .ZN( u2_u13_u5_n119 ) );
  NAND2_X1 u2_u13_u5_U62 (.A2( u2_u13_u5_n103 ) , .A1( u2_u13_u5_n105 ) , .ZN( u2_u13_u5_n140 ) );
  NAND2_X1 u2_u13_u5_U63 (.A2( u2_u13_u5_n104 ) , .A1( u2_u13_u5_n105 ) , .ZN( u2_u13_u5_n155 ) );
  NAND2_X1 u2_u13_u5_U64 (.A2( u2_u13_u5_n106 ) , .A1( u2_u13_u5_n107 ) , .ZN( u2_u13_u5_n122 ) );
  NAND2_X1 u2_u13_u5_U65 (.A2( u2_u13_u5_n100 ) , .A1( u2_u13_u5_n106 ) , .ZN( u2_u13_u5_n115 ) );
  NAND2_X1 u2_u13_u5_U66 (.A2( u2_u13_u5_n100 ) , .A1( u2_u13_u5_n103 ) , .ZN( u2_u13_u5_n161 ) );
  NAND2_X1 u2_u13_u5_U67 (.A1( u2_u13_u5_n105 ) , .A2( u2_u13_u5_n109 ) , .ZN( u2_u13_u5_n154 ) );
  INV_X1 u2_u13_u5_U68 (.A( u2_u13_u5_n146 ) , .ZN( u2_u13_u5_n172 ) );
  NAND2_X1 u2_u13_u5_U69 (.A1( u2_u13_u5_n103 ) , .A2( u2_u13_u5_n108 ) , .ZN( u2_u13_u5_n123 ) );
  OAI22_X1 u2_u13_u5_U7 (.B2( u2_u13_u5_n149 ) , .B1( u2_u13_u5_n150 ) , .A2( u2_u13_u5_n151 ) , .A1( u2_u13_u5_n152 ) , .ZN( u2_u13_u5_n165 ) );
  NAND2_X1 u2_u13_u5_U70 (.A2( u2_u13_u5_n103 ) , .A1( u2_u13_u5_n107 ) , .ZN( u2_u13_u5_n151 ) );
  NAND2_X1 u2_u13_u5_U71 (.A2( u2_u13_u5_n107 ) , .A1( u2_u13_u5_n109 ) , .ZN( u2_u13_u5_n120 ) );
  NAND2_X1 u2_u13_u5_U72 (.A2( u2_u13_u5_n100 ) , .A1( u2_u13_u5_n109 ) , .ZN( u2_u13_u5_n157 ) );
  AND2_X1 u2_u13_u5_U73 (.A2( u2_u13_u5_n100 ) , .A1( u2_u13_u5_n104 ) , .ZN( u2_u13_u5_n131 ) );
  INV_X1 u2_u13_u5_U74 (.A( u2_u13_u5_n102 ) , .ZN( u2_u13_u5_n195 ) );
  OAI221_X1 u2_u13_u5_U75 (.A( u2_u13_u5_n101 ) , .ZN( u2_u13_u5_n102 ) , .C2( u2_u13_u5_n115 ) , .C1( u2_u13_u5_n126 ) , .B1( u2_u13_u5_n134 ) , .B2( u2_u13_u5_n160 ) );
  OAI21_X1 u2_u13_u5_U76 (.ZN( u2_u13_u5_n101 ) , .B1( u2_u13_u5_n137 ) , .A( u2_u13_u5_n146 ) , .B2( u2_u13_u5_n147 ) );
  NOR2_X1 u2_u13_u5_U77 (.A2( u2_u13_X_34 ) , .A1( u2_u13_X_35 ) , .ZN( u2_u13_u5_n145 ) );
  NOR2_X1 u2_u13_u5_U78 (.A2( u2_u13_X_34 ) , .ZN( u2_u13_u5_n146 ) , .A1( u2_u13_u5_n171 ) );
  NOR2_X1 u2_u13_u5_U79 (.A2( u2_u13_X_31 ) , .A1( u2_u13_X_32 ) , .ZN( u2_u13_u5_n103 ) );
  NOR3_X1 u2_u13_u5_U8 (.A2( u2_u13_u5_n147 ) , .A1( u2_u13_u5_n148 ) , .ZN( u2_u13_u5_n149 ) , .A3( u2_u13_u5_n194 ) );
  NOR2_X1 u2_u13_u5_U80 (.A2( u2_u13_X_36 ) , .ZN( u2_u13_u5_n105 ) , .A1( u2_u13_u5_n180 ) );
  NOR2_X1 u2_u13_u5_U81 (.A2( u2_u13_X_33 ) , .ZN( u2_u13_u5_n108 ) , .A1( u2_u13_u5_n170 ) );
  NOR2_X1 u2_u13_u5_U82 (.A2( u2_u13_X_33 ) , .A1( u2_u13_X_36 ) , .ZN( u2_u13_u5_n107 ) );
  NOR2_X1 u2_u13_u5_U83 (.A2( u2_u13_X_31 ) , .ZN( u2_u13_u5_n104 ) , .A1( u2_u13_u5_n181 ) );
  NAND2_X1 u2_u13_u5_U84 (.A2( u2_u13_X_34 ) , .A1( u2_u13_X_35 ) , .ZN( u2_u13_u5_n153 ) );
  NAND2_X1 u2_u13_u5_U85 (.A1( u2_u13_X_34 ) , .ZN( u2_u13_u5_n126 ) , .A2( u2_u13_u5_n171 ) );
  AND2_X1 u2_u13_u5_U86 (.A1( u2_u13_X_31 ) , .A2( u2_u13_X_32 ) , .ZN( u2_u13_u5_n106 ) );
  AND2_X1 u2_u13_u5_U87 (.A1( u2_u13_X_31 ) , .ZN( u2_u13_u5_n109 ) , .A2( u2_u13_u5_n181 ) );
  INV_X1 u2_u13_u5_U88 (.A( u2_u13_X_33 ) , .ZN( u2_u13_u5_n180 ) );
  INV_X1 u2_u13_u5_U89 (.A( u2_u13_X_35 ) , .ZN( u2_u13_u5_n171 ) );
  NOR2_X1 u2_u13_u5_U9 (.ZN( u2_u13_u5_n135 ) , .A1( u2_u13_u5_n173 ) , .A2( u2_u13_u5_n176 ) );
  INV_X1 u2_u13_u5_U90 (.A( u2_u13_X_36 ) , .ZN( u2_u13_u5_n170 ) );
  INV_X1 u2_u13_u5_U91 (.A( u2_u13_X_32 ) , .ZN( u2_u13_u5_n181 ) );
  NAND4_X1 u2_u13_u5_U92 (.ZN( u2_out13_29 ) , .A4( u2_u13_u5_n129 ) , .A3( u2_u13_u5_n130 ) , .A2( u2_u13_u5_n168 ) , .A1( u2_u13_u5_n196 ) );
  AOI221_X1 u2_u13_u5_U93 (.A( u2_u13_u5_n128 ) , .ZN( u2_u13_u5_n129 ) , .C2( u2_u13_u5_n132 ) , .B2( u2_u13_u5_n159 ) , .B1( u2_u13_u5_n176 ) , .C1( u2_u13_u5_n184 ) );
  AOI222_X1 u2_u13_u5_U94 (.ZN( u2_u13_u5_n130 ) , .A2( u2_u13_u5_n146 ) , .B1( u2_u13_u5_n147 ) , .C2( u2_u13_u5_n175 ) , .B2( u2_u13_u5_n179 ) , .A1( u2_u13_u5_n188 ) , .C1( u2_u13_u5_n194 ) );
  NAND4_X1 u2_u13_u5_U95 (.ZN( u2_out13_19 ) , .A4( u2_u13_u5_n166 ) , .A3( u2_u13_u5_n167 ) , .A2( u2_u13_u5_n168 ) , .A1( u2_u13_u5_n169 ) );
  AOI22_X1 u2_u13_u5_U96 (.B2( u2_u13_u5_n145 ) , .A2( u2_u13_u5_n146 ) , .ZN( u2_u13_u5_n167 ) , .B1( u2_u13_u5_n182 ) , .A1( u2_u13_u5_n189 ) );
  NOR4_X1 u2_u13_u5_U97 (.A4( u2_u13_u5_n162 ) , .A3( u2_u13_u5_n163 ) , .A2( u2_u13_u5_n164 ) , .A1( u2_u13_u5_n165 ) , .ZN( u2_u13_u5_n166 ) );
  NAND4_X1 u2_u13_u5_U98 (.ZN( u2_out13_11 ) , .A4( u2_u13_u5_n143 ) , .A3( u2_u13_u5_n144 ) , .A2( u2_u13_u5_n169 ) , .A1( u2_u13_u5_n196 ) );
  AOI22_X1 u2_u13_u5_U99 (.A2( u2_u13_u5_n132 ) , .ZN( u2_u13_u5_n144 ) , .B2( u2_u13_u5_n145 ) , .B1( u2_u13_u5_n184 ) , .A1( u2_u13_u5_n194 ) );
  XOR2_X1 u2_u14_U1 (.B( u2_K15_9 ) , .A( u2_R13_6 ) , .Z( u2_u14_X_9 ) );
  XOR2_X1 u2_u14_U13 (.B( u2_K15_42 ) , .A( u2_R13_29 ) , .Z( u2_u14_X_42 ) );
  XOR2_X1 u2_u14_U14 (.B( u2_K15_41 ) , .A( u2_R13_28 ) , .Z( u2_u14_X_41 ) );
  XOR2_X1 u2_u14_U15 (.B( u2_K15_40 ) , .A( u2_R13_27 ) , .Z( u2_u14_X_40 ) );
  XOR2_X1 u2_u14_U16 (.B( u2_K15_3 ) , .A( u2_R13_2 ) , .Z( u2_u14_X_3 ) );
  XOR2_X1 u2_u14_U17 (.B( u2_K15_39 ) , .A( u2_R13_26 ) , .Z( u2_u14_X_39 ) );
  XOR2_X1 u2_u14_U18 (.B( u2_K15_38 ) , .A( u2_R13_25 ) , .Z( u2_u14_X_38 ) );
  XOR2_X1 u2_u14_U19 (.B( u2_K15_37 ) , .A( u2_R13_24 ) , .Z( u2_u14_X_37 ) );
  XOR2_X1 u2_u14_U2 (.B( u2_K15_8 ) , .A( u2_R13_5 ) , .Z( u2_u14_X_8 ) );
  XOR2_X1 u2_u14_U20 (.B( u2_K15_36 ) , .A( u2_R13_25 ) , .Z( u2_u14_X_36 ) );
  XOR2_X1 u2_u14_U21 (.B( u2_K15_35 ) , .A( u2_R13_24 ) , .Z( u2_u14_X_35 ) );
  XOR2_X1 u2_u14_U22 (.B( u2_K15_34 ) , .A( u2_R13_23 ) , .Z( u2_u14_X_34 ) );
  XOR2_X1 u2_u14_U23 (.B( u2_K15_33 ) , .A( u2_R13_22 ) , .Z( u2_u14_X_33 ) );
  XOR2_X1 u2_u14_U24 (.B( u2_K15_32 ) , .A( u2_R13_21 ) , .Z( u2_u14_X_32 ) );
  XOR2_X1 u2_u14_U25 (.B( u2_K15_31 ) , .A( u2_R13_20 ) , .Z( u2_u14_X_31 ) );
  XOR2_X1 u2_u14_U26 (.B( u2_K15_30 ) , .A( u2_R13_21 ) , .Z( u2_u14_X_30 ) );
  XOR2_X1 u2_u14_U27 (.B( u2_K15_2 ) , .A( u2_R13_1 ) , .Z( u2_u14_X_2 ) );
  XOR2_X1 u2_u14_U28 (.B( u2_K15_29 ) , .A( u2_R13_20 ) , .Z( u2_u14_X_29 ) );
  XOR2_X1 u2_u14_U29 (.B( u2_K15_28 ) , .A( u2_R13_19 ) , .Z( u2_u14_X_28 ) );
  XOR2_X1 u2_u14_U3 (.B( u2_K15_7 ) , .A( u2_R13_4 ) , .Z( u2_u14_X_7 ) );
  XOR2_X1 u2_u14_U30 (.B( u2_K15_27 ) , .A( u2_R13_18 ) , .Z( u2_u14_X_27 ) );
  XOR2_X1 u2_u14_U31 (.B( u2_K15_26 ) , .A( u2_R13_17 ) , .Z( u2_u14_X_26 ) );
  XOR2_X1 u2_u14_U32 (.B( u2_K15_25 ) , .A( u2_R13_16 ) , .Z( u2_u14_X_25 ) );
  XOR2_X1 u2_u14_U38 (.B( u2_K15_1 ) , .A( u2_R13_32 ) , .Z( u2_u14_X_1 ) );
  XOR2_X1 u2_u14_U4 (.B( u2_K15_6 ) , .A( u2_R13_5 ) , .Z( u2_u14_X_6 ) );
  XOR2_X1 u2_u14_U46 (.B( u2_K15_12 ) , .A( u2_R13_9 ) , .Z( u2_u14_X_12 ) );
  XOR2_X1 u2_u14_U47 (.B( u2_K15_11 ) , .A( u2_R13_8 ) , .Z( u2_u14_X_11 ) );
  XOR2_X1 u2_u14_U48 (.B( u2_K15_10 ) , .A( u2_R13_7 ) , .Z( u2_u14_X_10 ) );
  XOR2_X1 u2_u14_U5 (.B( u2_K15_5 ) , .A( u2_R13_4 ) , .Z( u2_u14_X_5 ) );
  XOR2_X1 u2_u14_U6 (.B( u2_K15_4 ) , .A( u2_R13_3 ) , .Z( u2_u14_X_4 ) );
  AND3_X1 u2_u14_u0_U10 (.A2( u2_u14_u0_n112 ) , .ZN( u2_u14_u0_n127 ) , .A3( u2_u14_u0_n130 ) , .A1( u2_u14_u0_n148 ) );
  NAND2_X1 u2_u14_u0_U11 (.ZN( u2_u14_u0_n113 ) , .A1( u2_u14_u0_n139 ) , .A2( u2_u14_u0_n149 ) );
  AND2_X1 u2_u14_u0_U12 (.ZN( u2_u14_u0_n107 ) , .A1( u2_u14_u0_n130 ) , .A2( u2_u14_u0_n140 ) );
  AND2_X1 u2_u14_u0_U13 (.A2( u2_u14_u0_n129 ) , .A1( u2_u14_u0_n130 ) , .ZN( u2_u14_u0_n151 ) );
  AND2_X1 u2_u14_u0_U14 (.A1( u2_u14_u0_n108 ) , .A2( u2_u14_u0_n125 ) , .ZN( u2_u14_u0_n145 ) );
  INV_X1 u2_u14_u0_U15 (.A( u2_u14_u0_n143 ) , .ZN( u2_u14_u0_n173 ) );
  NOR2_X1 u2_u14_u0_U16 (.A2( u2_u14_u0_n136 ) , .ZN( u2_u14_u0_n147 ) , .A1( u2_u14_u0_n160 ) );
  NOR2_X1 u2_u14_u0_U17 (.A1( u2_u14_u0_n163 ) , .A2( u2_u14_u0_n164 ) , .ZN( u2_u14_u0_n95 ) );
  AOI21_X1 u2_u14_u0_U18 (.B1( u2_u14_u0_n103 ) , .ZN( u2_u14_u0_n132 ) , .A( u2_u14_u0_n165 ) , .B2( u2_u14_u0_n93 ) );
  INV_X1 u2_u14_u0_U19 (.A( u2_u14_u0_n142 ) , .ZN( u2_u14_u0_n165 ) );
  OAI221_X1 u2_u14_u0_U20 (.C1( u2_u14_u0_n121 ) , .ZN( u2_u14_u0_n122 ) , .B2( u2_u14_u0_n127 ) , .A( u2_u14_u0_n143 ) , .B1( u2_u14_u0_n144 ) , .C2( u2_u14_u0_n147 ) );
  OAI22_X1 u2_u14_u0_U21 (.B1( u2_u14_u0_n125 ) , .ZN( u2_u14_u0_n126 ) , .A1( u2_u14_u0_n138 ) , .A2( u2_u14_u0_n146 ) , .B2( u2_u14_u0_n147 ) );
  OAI22_X1 u2_u14_u0_U22 (.B1( u2_u14_u0_n131 ) , .A1( u2_u14_u0_n144 ) , .B2( u2_u14_u0_n147 ) , .A2( u2_u14_u0_n90 ) , .ZN( u2_u14_u0_n91 ) );
  AND3_X1 u2_u14_u0_U23 (.A3( u2_u14_u0_n121 ) , .A2( u2_u14_u0_n125 ) , .A1( u2_u14_u0_n148 ) , .ZN( u2_u14_u0_n90 ) );
  INV_X1 u2_u14_u0_U24 (.A( u2_u14_u0_n136 ) , .ZN( u2_u14_u0_n161 ) );
  NOR2_X1 u2_u14_u0_U25 (.A1( u2_u14_u0_n120 ) , .ZN( u2_u14_u0_n143 ) , .A2( u2_u14_u0_n167 ) );
  OAI221_X1 u2_u14_u0_U26 (.C1( u2_u14_u0_n112 ) , .ZN( u2_u14_u0_n120 ) , .B1( u2_u14_u0_n138 ) , .B2( u2_u14_u0_n141 ) , .C2( u2_u14_u0_n147 ) , .A( u2_u14_u0_n172 ) );
  AOI211_X1 u2_u14_u0_U27 (.B( u2_u14_u0_n115 ) , .A( u2_u14_u0_n116 ) , .C2( u2_u14_u0_n117 ) , .C1( u2_u14_u0_n118 ) , .ZN( u2_u14_u0_n119 ) );
  AOI22_X1 u2_u14_u0_U28 (.B2( u2_u14_u0_n109 ) , .A2( u2_u14_u0_n110 ) , .ZN( u2_u14_u0_n111 ) , .B1( u2_u14_u0_n118 ) , .A1( u2_u14_u0_n160 ) );
  INV_X1 u2_u14_u0_U29 (.A( u2_u14_u0_n118 ) , .ZN( u2_u14_u0_n158 ) );
  INV_X1 u2_u14_u0_U3 (.A( u2_u14_u0_n113 ) , .ZN( u2_u14_u0_n166 ) );
  AOI21_X1 u2_u14_u0_U30 (.ZN( u2_u14_u0_n104 ) , .B1( u2_u14_u0_n107 ) , .B2( u2_u14_u0_n141 ) , .A( u2_u14_u0_n144 ) );
  AOI21_X1 u2_u14_u0_U31 (.B1( u2_u14_u0_n127 ) , .B2( u2_u14_u0_n129 ) , .A( u2_u14_u0_n138 ) , .ZN( u2_u14_u0_n96 ) );
  AOI21_X1 u2_u14_u0_U32 (.ZN( u2_u14_u0_n116 ) , .B2( u2_u14_u0_n142 ) , .A( u2_u14_u0_n144 ) , .B1( u2_u14_u0_n166 ) );
  NAND2_X1 u2_u14_u0_U33 (.A1( u2_u14_u0_n100 ) , .A2( u2_u14_u0_n103 ) , .ZN( u2_u14_u0_n125 ) );
  NAND2_X1 u2_u14_u0_U34 (.A2( u2_u14_u0_n103 ) , .ZN( u2_u14_u0_n140 ) , .A1( u2_u14_u0_n94 ) );
  NAND2_X1 u2_u14_u0_U35 (.A1( u2_u14_u0_n101 ) , .A2( u2_u14_u0_n102 ) , .ZN( u2_u14_u0_n150 ) );
  INV_X1 u2_u14_u0_U36 (.A( u2_u14_u0_n138 ) , .ZN( u2_u14_u0_n160 ) );
  NAND2_X1 u2_u14_u0_U37 (.ZN( u2_u14_u0_n142 ) , .A1( u2_u14_u0_n94 ) , .A2( u2_u14_u0_n95 ) );
  NAND2_X1 u2_u14_u0_U38 (.A1( u2_u14_u0_n102 ) , .ZN( u2_u14_u0_n128 ) , .A2( u2_u14_u0_n95 ) );
  NAND2_X1 u2_u14_u0_U39 (.A2( u2_u14_u0_n102 ) , .A1( u2_u14_u0_n103 ) , .ZN( u2_u14_u0_n149 ) );
  AOI21_X1 u2_u14_u0_U4 (.B1( u2_u14_u0_n114 ) , .ZN( u2_u14_u0_n115 ) , .B2( u2_u14_u0_n129 ) , .A( u2_u14_u0_n161 ) );
  NAND2_X1 u2_u14_u0_U40 (.A1( u2_u14_u0_n100 ) , .ZN( u2_u14_u0_n129 ) , .A2( u2_u14_u0_n95 ) );
  NAND2_X1 u2_u14_u0_U41 (.A2( u2_u14_u0_n100 ) , .A1( u2_u14_u0_n101 ) , .ZN( u2_u14_u0_n139 ) );
  NAND2_X1 u2_u14_u0_U42 (.A2( u2_u14_u0_n100 ) , .ZN( u2_u14_u0_n131 ) , .A1( u2_u14_u0_n92 ) );
  NAND2_X1 u2_u14_u0_U43 (.ZN( u2_u14_u0_n108 ) , .A1( u2_u14_u0_n92 ) , .A2( u2_u14_u0_n94 ) );
  NAND2_X1 u2_u14_u0_U44 (.ZN( u2_u14_u0_n148 ) , .A1( u2_u14_u0_n93 ) , .A2( u2_u14_u0_n95 ) );
  NAND2_X1 u2_u14_u0_U45 (.A2( u2_u14_u0_n102 ) , .ZN( u2_u14_u0_n114 ) , .A1( u2_u14_u0_n92 ) );
  NAND2_X1 u2_u14_u0_U46 (.A1( u2_u14_u0_n101 ) , .ZN( u2_u14_u0_n130 ) , .A2( u2_u14_u0_n94 ) );
  NAND2_X1 u2_u14_u0_U47 (.A2( u2_u14_u0_n101 ) , .ZN( u2_u14_u0_n121 ) , .A1( u2_u14_u0_n93 ) );
  INV_X1 u2_u14_u0_U48 (.ZN( u2_u14_u0_n172 ) , .A( u2_u14_u0_n88 ) );
  OAI222_X1 u2_u14_u0_U49 (.C1( u2_u14_u0_n108 ) , .A1( u2_u14_u0_n125 ) , .B2( u2_u14_u0_n128 ) , .B1( u2_u14_u0_n144 ) , .A2( u2_u14_u0_n158 ) , .C2( u2_u14_u0_n161 ) , .ZN( u2_u14_u0_n88 ) );
  AOI21_X1 u2_u14_u0_U5 (.B2( u2_u14_u0_n131 ) , .ZN( u2_u14_u0_n134 ) , .B1( u2_u14_u0_n151 ) , .A( u2_u14_u0_n158 ) );
  NAND2_X1 u2_u14_u0_U50 (.ZN( u2_u14_u0_n112 ) , .A2( u2_u14_u0_n92 ) , .A1( u2_u14_u0_n93 ) );
  OR3_X1 u2_u14_u0_U51 (.A3( u2_u14_u0_n152 ) , .A2( u2_u14_u0_n153 ) , .A1( u2_u14_u0_n154 ) , .ZN( u2_u14_u0_n155 ) );
  AOI21_X1 u2_u14_u0_U52 (.B2( u2_u14_u0_n150 ) , .B1( u2_u14_u0_n151 ) , .ZN( u2_u14_u0_n152 ) , .A( u2_u14_u0_n158 ) );
  AOI21_X1 u2_u14_u0_U53 (.A( u2_u14_u0_n144 ) , .B2( u2_u14_u0_n145 ) , .B1( u2_u14_u0_n146 ) , .ZN( u2_u14_u0_n154 ) );
  AOI21_X1 u2_u14_u0_U54 (.A( u2_u14_u0_n147 ) , .B2( u2_u14_u0_n148 ) , .B1( u2_u14_u0_n149 ) , .ZN( u2_u14_u0_n153 ) );
  INV_X1 u2_u14_u0_U55 (.ZN( u2_u14_u0_n171 ) , .A( u2_u14_u0_n99 ) );
  OAI211_X1 u2_u14_u0_U56 (.C2( u2_u14_u0_n140 ) , .C1( u2_u14_u0_n161 ) , .A( u2_u14_u0_n169 ) , .B( u2_u14_u0_n98 ) , .ZN( u2_u14_u0_n99 ) );
  INV_X1 u2_u14_u0_U57 (.ZN( u2_u14_u0_n169 ) , .A( u2_u14_u0_n91 ) );
  AOI211_X1 u2_u14_u0_U58 (.C1( u2_u14_u0_n118 ) , .A( u2_u14_u0_n123 ) , .B( u2_u14_u0_n96 ) , .C2( u2_u14_u0_n97 ) , .ZN( u2_u14_u0_n98 ) );
  NOR2_X1 u2_u14_u0_U59 (.A2( u2_u14_X_2 ) , .ZN( u2_u14_u0_n103 ) , .A1( u2_u14_u0_n164 ) );
  NOR2_X1 u2_u14_u0_U6 (.A1( u2_u14_u0_n108 ) , .ZN( u2_u14_u0_n123 ) , .A2( u2_u14_u0_n158 ) );
  NOR2_X1 u2_u14_u0_U60 (.A2( u2_u14_X_3 ) , .A1( u2_u14_X_6 ) , .ZN( u2_u14_u0_n94 ) );
  NOR2_X1 u2_u14_u0_U61 (.A2( u2_u14_X_6 ) , .ZN( u2_u14_u0_n100 ) , .A1( u2_u14_u0_n162 ) );
  NOR2_X1 u2_u14_u0_U62 (.A2( u2_u14_X_4 ) , .A1( u2_u14_X_5 ) , .ZN( u2_u14_u0_n118 ) );
  NOR2_X1 u2_u14_u0_U63 (.A2( u2_u14_X_1 ) , .A1( u2_u14_X_2 ) , .ZN( u2_u14_u0_n92 ) );
  NOR2_X1 u2_u14_u0_U64 (.A2( u2_u14_X_1 ) , .ZN( u2_u14_u0_n101 ) , .A1( u2_u14_u0_n163 ) );
  NAND2_X1 u2_u14_u0_U65 (.A2( u2_u14_X_4 ) , .A1( u2_u14_X_5 ) , .ZN( u2_u14_u0_n144 ) );
  NOR2_X1 u2_u14_u0_U66 (.A2( u2_u14_X_5 ) , .ZN( u2_u14_u0_n136 ) , .A1( u2_u14_u0_n159 ) );
  NAND2_X1 u2_u14_u0_U67 (.A1( u2_u14_X_5 ) , .ZN( u2_u14_u0_n138 ) , .A2( u2_u14_u0_n159 ) );
  AND2_X1 u2_u14_u0_U68 (.A2( u2_u14_X_3 ) , .A1( u2_u14_X_6 ) , .ZN( u2_u14_u0_n102 ) );
  AND2_X1 u2_u14_u0_U69 (.A1( u2_u14_X_6 ) , .A2( u2_u14_u0_n162 ) , .ZN( u2_u14_u0_n93 ) );
  OAI21_X1 u2_u14_u0_U7 (.B1( u2_u14_u0_n150 ) , .B2( u2_u14_u0_n158 ) , .A( u2_u14_u0_n172 ) , .ZN( u2_u14_u0_n89 ) );
  INV_X1 u2_u14_u0_U70 (.A( u2_u14_X_4 ) , .ZN( u2_u14_u0_n159 ) );
  INV_X1 u2_u14_u0_U71 (.A( u2_u14_X_1 ) , .ZN( u2_u14_u0_n164 ) );
  INV_X1 u2_u14_u0_U72 (.A( u2_u14_X_2 ) , .ZN( u2_u14_u0_n163 ) );
  INV_X1 u2_u14_u0_U73 (.A( u2_u14_X_3 ) , .ZN( u2_u14_u0_n162 ) );
  INV_X1 u2_u14_u0_U74 (.A( u2_u14_u0_n126 ) , .ZN( u2_u14_u0_n168 ) );
  AOI211_X1 u2_u14_u0_U75 (.B( u2_u14_u0_n133 ) , .A( u2_u14_u0_n134 ) , .C2( u2_u14_u0_n135 ) , .C1( u2_u14_u0_n136 ) , .ZN( u2_u14_u0_n137 ) );
  INV_X1 u2_u14_u0_U76 (.ZN( u2_u14_u0_n174 ) , .A( u2_u14_u0_n89 ) );
  AOI211_X1 u2_u14_u0_U77 (.B( u2_u14_u0_n104 ) , .A( u2_u14_u0_n105 ) , .ZN( u2_u14_u0_n106 ) , .C2( u2_u14_u0_n113 ) , .C1( u2_u14_u0_n160 ) );
  OR4_X1 u2_u14_u0_U78 (.ZN( u2_out14_17 ) , .A4( u2_u14_u0_n122 ) , .A2( u2_u14_u0_n123 ) , .A1( u2_u14_u0_n124 ) , .A3( u2_u14_u0_n170 ) );
  AOI21_X1 u2_u14_u0_U79 (.B2( u2_u14_u0_n107 ) , .ZN( u2_u14_u0_n124 ) , .B1( u2_u14_u0_n128 ) , .A( u2_u14_u0_n161 ) );
  AND2_X1 u2_u14_u0_U8 (.A1( u2_u14_u0_n114 ) , .A2( u2_u14_u0_n121 ) , .ZN( u2_u14_u0_n146 ) );
  INV_X1 u2_u14_u0_U80 (.A( u2_u14_u0_n111 ) , .ZN( u2_u14_u0_n170 ) );
  OR4_X1 u2_u14_u0_U81 (.ZN( u2_out14_31 ) , .A4( u2_u14_u0_n155 ) , .A2( u2_u14_u0_n156 ) , .A1( u2_u14_u0_n157 ) , .A3( u2_u14_u0_n173 ) );
  AOI21_X1 u2_u14_u0_U82 (.A( u2_u14_u0_n138 ) , .B2( u2_u14_u0_n139 ) , .B1( u2_u14_u0_n140 ) , .ZN( u2_u14_u0_n157 ) );
  AOI21_X1 u2_u14_u0_U83 (.B2( u2_u14_u0_n141 ) , .B1( u2_u14_u0_n142 ) , .ZN( u2_u14_u0_n156 ) , .A( u2_u14_u0_n161 ) );
  AOI21_X1 u2_u14_u0_U84 (.B1( u2_u14_u0_n132 ) , .ZN( u2_u14_u0_n133 ) , .A( u2_u14_u0_n144 ) , .B2( u2_u14_u0_n166 ) );
  OAI22_X1 u2_u14_u0_U85 (.ZN( u2_u14_u0_n105 ) , .A2( u2_u14_u0_n132 ) , .B1( u2_u14_u0_n146 ) , .A1( u2_u14_u0_n147 ) , .B2( u2_u14_u0_n161 ) );
  NAND2_X1 u2_u14_u0_U86 (.ZN( u2_u14_u0_n110 ) , .A2( u2_u14_u0_n132 ) , .A1( u2_u14_u0_n145 ) );
  INV_X1 u2_u14_u0_U87 (.A( u2_u14_u0_n119 ) , .ZN( u2_u14_u0_n167 ) );
  NAND3_X1 u2_u14_u0_U88 (.ZN( u2_out14_23 ) , .A3( u2_u14_u0_n137 ) , .A1( u2_u14_u0_n168 ) , .A2( u2_u14_u0_n171 ) );
  NAND3_X1 u2_u14_u0_U89 (.A3( u2_u14_u0_n127 ) , .A2( u2_u14_u0_n128 ) , .ZN( u2_u14_u0_n135 ) , .A1( u2_u14_u0_n150 ) );
  AND2_X1 u2_u14_u0_U9 (.A1( u2_u14_u0_n131 ) , .ZN( u2_u14_u0_n141 ) , .A2( u2_u14_u0_n150 ) );
  NAND3_X1 u2_u14_u0_U90 (.ZN( u2_u14_u0_n117 ) , .A3( u2_u14_u0_n132 ) , .A2( u2_u14_u0_n139 ) , .A1( u2_u14_u0_n148 ) );
  NAND3_X1 u2_u14_u0_U91 (.ZN( u2_u14_u0_n109 ) , .A2( u2_u14_u0_n114 ) , .A3( u2_u14_u0_n140 ) , .A1( u2_u14_u0_n149 ) );
  NAND3_X1 u2_u14_u0_U92 (.ZN( u2_out14_9 ) , .A3( u2_u14_u0_n106 ) , .A2( u2_u14_u0_n171 ) , .A1( u2_u14_u0_n174 ) );
  NAND3_X1 u2_u14_u0_U93 (.A2( u2_u14_u0_n128 ) , .A1( u2_u14_u0_n132 ) , .A3( u2_u14_u0_n146 ) , .ZN( u2_u14_u0_n97 ) );
  AOI21_X1 u2_u14_u1_U10 (.ZN( u2_u14_u1_n106 ) , .A( u2_u14_u1_n112 ) , .B1( u2_u14_u1_n154 ) , .B2( u2_u14_u1_n156 ) );
  NAND3_X1 u2_u14_u1_U100 (.ZN( u2_u14_u1_n113 ) , .A1( u2_u14_u1_n120 ) , .A3( u2_u14_u1_n133 ) , .A2( u2_u14_u1_n155 ) );
  INV_X1 u2_u14_u1_U11 (.A( u2_u14_u1_n101 ) , .ZN( u2_u14_u1_n184 ) );
  AOI21_X1 u2_u14_u1_U12 (.ZN( u2_u14_u1_n107 ) , .B1( u2_u14_u1_n134 ) , .B2( u2_u14_u1_n149 ) , .A( u2_u14_u1_n174 ) );
  NAND2_X1 u2_u14_u1_U13 (.ZN( u2_u14_u1_n140 ) , .A2( u2_u14_u1_n150 ) , .A1( u2_u14_u1_n155 ) );
  NAND2_X1 u2_u14_u1_U14 (.A1( u2_u14_u1_n131 ) , .ZN( u2_u14_u1_n147 ) , .A2( u2_u14_u1_n153 ) );
  AOI22_X1 u2_u14_u1_U15 (.B2( u2_u14_u1_n136 ) , .A2( u2_u14_u1_n137 ) , .ZN( u2_u14_u1_n143 ) , .A1( u2_u14_u1_n171 ) , .B1( u2_u14_u1_n173 ) );
  INV_X1 u2_u14_u1_U16 (.A( u2_u14_u1_n147 ) , .ZN( u2_u14_u1_n181 ) );
  INV_X1 u2_u14_u1_U17 (.A( u2_u14_u1_n139 ) , .ZN( u2_u14_u1_n174 ) );
  INV_X1 u2_u14_u1_U18 (.A( u2_u14_u1_n112 ) , .ZN( u2_u14_u1_n171 ) );
  NAND2_X1 u2_u14_u1_U19 (.ZN( u2_u14_u1_n141 ) , .A1( u2_u14_u1_n153 ) , .A2( u2_u14_u1_n156 ) );
  AND2_X1 u2_u14_u1_U20 (.A1( u2_u14_u1_n123 ) , .ZN( u2_u14_u1_n134 ) , .A2( u2_u14_u1_n161 ) );
  NAND2_X1 u2_u14_u1_U21 (.A2( u2_u14_u1_n115 ) , .A1( u2_u14_u1_n116 ) , .ZN( u2_u14_u1_n148 ) );
  NAND2_X1 u2_u14_u1_U22 (.A2( u2_u14_u1_n133 ) , .A1( u2_u14_u1_n135 ) , .ZN( u2_u14_u1_n159 ) );
  NAND2_X1 u2_u14_u1_U23 (.A2( u2_u14_u1_n115 ) , .A1( u2_u14_u1_n120 ) , .ZN( u2_u14_u1_n132 ) );
  INV_X1 u2_u14_u1_U24 (.A( u2_u14_u1_n154 ) , .ZN( u2_u14_u1_n178 ) );
  AOI22_X1 u2_u14_u1_U25 (.B2( u2_u14_u1_n113 ) , .A2( u2_u14_u1_n114 ) , .ZN( u2_u14_u1_n125 ) , .A1( u2_u14_u1_n171 ) , .B1( u2_u14_u1_n173 ) );
  NAND2_X1 u2_u14_u1_U26 (.ZN( u2_u14_u1_n114 ) , .A1( u2_u14_u1_n134 ) , .A2( u2_u14_u1_n156 ) );
  INV_X1 u2_u14_u1_U27 (.A( u2_u14_u1_n151 ) , .ZN( u2_u14_u1_n183 ) );
  AND2_X1 u2_u14_u1_U28 (.A1( u2_u14_u1_n129 ) , .A2( u2_u14_u1_n133 ) , .ZN( u2_u14_u1_n149 ) );
  INV_X1 u2_u14_u1_U29 (.A( u2_u14_u1_n131 ) , .ZN( u2_u14_u1_n180 ) );
  INV_X1 u2_u14_u1_U3 (.A( u2_u14_u1_n159 ) , .ZN( u2_u14_u1_n182 ) );
  AOI221_X1 u2_u14_u1_U30 (.B1( u2_u14_u1_n140 ) , .ZN( u2_u14_u1_n167 ) , .B2( u2_u14_u1_n172 ) , .C2( u2_u14_u1_n175 ) , .C1( u2_u14_u1_n178 ) , .A( u2_u14_u1_n188 ) );
  INV_X1 u2_u14_u1_U31 (.ZN( u2_u14_u1_n188 ) , .A( u2_u14_u1_n97 ) );
  AOI211_X1 u2_u14_u1_U32 (.A( u2_u14_u1_n118 ) , .C1( u2_u14_u1_n132 ) , .C2( u2_u14_u1_n139 ) , .B( u2_u14_u1_n96 ) , .ZN( u2_u14_u1_n97 ) );
  AOI21_X1 u2_u14_u1_U33 (.B2( u2_u14_u1_n121 ) , .B1( u2_u14_u1_n135 ) , .A( u2_u14_u1_n152 ) , .ZN( u2_u14_u1_n96 ) );
  OAI221_X1 u2_u14_u1_U34 (.A( u2_u14_u1_n119 ) , .C2( u2_u14_u1_n129 ) , .ZN( u2_u14_u1_n138 ) , .B2( u2_u14_u1_n152 ) , .C1( u2_u14_u1_n174 ) , .B1( u2_u14_u1_n187 ) );
  INV_X1 u2_u14_u1_U35 (.A( u2_u14_u1_n148 ) , .ZN( u2_u14_u1_n187 ) );
  AOI211_X1 u2_u14_u1_U36 (.B( u2_u14_u1_n117 ) , .A( u2_u14_u1_n118 ) , .ZN( u2_u14_u1_n119 ) , .C2( u2_u14_u1_n146 ) , .C1( u2_u14_u1_n159 ) );
  NOR2_X1 u2_u14_u1_U37 (.A1( u2_u14_u1_n168 ) , .A2( u2_u14_u1_n176 ) , .ZN( u2_u14_u1_n98 ) );
  AOI211_X1 u2_u14_u1_U38 (.B( u2_u14_u1_n162 ) , .A( u2_u14_u1_n163 ) , .C2( u2_u14_u1_n164 ) , .ZN( u2_u14_u1_n165 ) , .C1( u2_u14_u1_n171 ) );
  AOI21_X1 u2_u14_u1_U39 (.A( u2_u14_u1_n160 ) , .B2( u2_u14_u1_n161 ) , .ZN( u2_u14_u1_n162 ) , .B1( u2_u14_u1_n182 ) );
  AOI221_X1 u2_u14_u1_U4 (.A( u2_u14_u1_n138 ) , .C2( u2_u14_u1_n139 ) , .C1( u2_u14_u1_n140 ) , .B2( u2_u14_u1_n141 ) , .ZN( u2_u14_u1_n142 ) , .B1( u2_u14_u1_n175 ) );
  OR2_X1 u2_u14_u1_U40 (.A2( u2_u14_u1_n157 ) , .A1( u2_u14_u1_n158 ) , .ZN( u2_u14_u1_n163 ) );
  OAI21_X1 u2_u14_u1_U41 (.B2( u2_u14_u1_n123 ) , .ZN( u2_u14_u1_n145 ) , .B1( u2_u14_u1_n160 ) , .A( u2_u14_u1_n185 ) );
  INV_X1 u2_u14_u1_U42 (.A( u2_u14_u1_n122 ) , .ZN( u2_u14_u1_n185 ) );
  AOI21_X1 u2_u14_u1_U43 (.B2( u2_u14_u1_n120 ) , .B1( u2_u14_u1_n121 ) , .ZN( u2_u14_u1_n122 ) , .A( u2_u14_u1_n128 ) );
  NAND2_X1 u2_u14_u1_U44 (.A1( u2_u14_u1_n128 ) , .ZN( u2_u14_u1_n146 ) , .A2( u2_u14_u1_n160 ) );
  NAND2_X1 u2_u14_u1_U45 (.A2( u2_u14_u1_n112 ) , .ZN( u2_u14_u1_n139 ) , .A1( u2_u14_u1_n152 ) );
  NAND2_X1 u2_u14_u1_U46 (.A1( u2_u14_u1_n105 ) , .ZN( u2_u14_u1_n156 ) , .A2( u2_u14_u1_n99 ) );
  NOR2_X1 u2_u14_u1_U47 (.ZN( u2_u14_u1_n117 ) , .A1( u2_u14_u1_n121 ) , .A2( u2_u14_u1_n160 ) );
  AOI21_X1 u2_u14_u1_U48 (.A( u2_u14_u1_n128 ) , .B2( u2_u14_u1_n129 ) , .ZN( u2_u14_u1_n130 ) , .B1( u2_u14_u1_n150 ) );
  NAND2_X1 u2_u14_u1_U49 (.ZN( u2_u14_u1_n112 ) , .A1( u2_u14_u1_n169 ) , .A2( u2_u14_u1_n170 ) );
  AOI211_X1 u2_u14_u1_U5 (.ZN( u2_u14_u1_n124 ) , .A( u2_u14_u1_n138 ) , .C2( u2_u14_u1_n139 ) , .B( u2_u14_u1_n145 ) , .C1( u2_u14_u1_n147 ) );
  NAND2_X1 u2_u14_u1_U50 (.ZN( u2_u14_u1_n129 ) , .A2( u2_u14_u1_n95 ) , .A1( u2_u14_u1_n98 ) );
  NAND2_X1 u2_u14_u1_U51 (.A1( u2_u14_u1_n102 ) , .ZN( u2_u14_u1_n154 ) , .A2( u2_u14_u1_n99 ) );
  NAND2_X1 u2_u14_u1_U52 (.A2( u2_u14_u1_n100 ) , .ZN( u2_u14_u1_n135 ) , .A1( u2_u14_u1_n99 ) );
  AOI21_X1 u2_u14_u1_U53 (.A( u2_u14_u1_n152 ) , .B2( u2_u14_u1_n153 ) , .B1( u2_u14_u1_n154 ) , .ZN( u2_u14_u1_n158 ) );
  INV_X1 u2_u14_u1_U54 (.A( u2_u14_u1_n160 ) , .ZN( u2_u14_u1_n175 ) );
  NAND2_X1 u2_u14_u1_U55 (.A1( u2_u14_u1_n100 ) , .ZN( u2_u14_u1_n116 ) , .A2( u2_u14_u1_n95 ) );
  NAND2_X1 u2_u14_u1_U56 (.A1( u2_u14_u1_n102 ) , .ZN( u2_u14_u1_n131 ) , .A2( u2_u14_u1_n95 ) );
  NAND2_X1 u2_u14_u1_U57 (.A2( u2_u14_u1_n104 ) , .ZN( u2_u14_u1_n121 ) , .A1( u2_u14_u1_n98 ) );
  NAND2_X1 u2_u14_u1_U58 (.A1( u2_u14_u1_n103 ) , .ZN( u2_u14_u1_n153 ) , .A2( u2_u14_u1_n98 ) );
  NAND2_X1 u2_u14_u1_U59 (.A2( u2_u14_u1_n104 ) , .A1( u2_u14_u1_n105 ) , .ZN( u2_u14_u1_n133 ) );
  NOR2_X1 u2_u14_u1_U6 (.A1( u2_u14_u1_n112 ) , .A2( u2_u14_u1_n116 ) , .ZN( u2_u14_u1_n118 ) );
  NAND2_X1 u2_u14_u1_U60 (.ZN( u2_u14_u1_n150 ) , .A2( u2_u14_u1_n98 ) , .A1( u2_u14_u1_n99 ) );
  NAND2_X1 u2_u14_u1_U61 (.A1( u2_u14_u1_n105 ) , .ZN( u2_u14_u1_n155 ) , .A2( u2_u14_u1_n95 ) );
  OAI21_X1 u2_u14_u1_U62 (.ZN( u2_u14_u1_n109 ) , .B1( u2_u14_u1_n129 ) , .B2( u2_u14_u1_n160 ) , .A( u2_u14_u1_n167 ) );
  NAND2_X1 u2_u14_u1_U63 (.A2( u2_u14_u1_n100 ) , .A1( u2_u14_u1_n103 ) , .ZN( u2_u14_u1_n120 ) );
  NAND2_X1 u2_u14_u1_U64 (.A1( u2_u14_u1_n102 ) , .A2( u2_u14_u1_n104 ) , .ZN( u2_u14_u1_n115 ) );
  NAND2_X1 u2_u14_u1_U65 (.A2( u2_u14_u1_n100 ) , .A1( u2_u14_u1_n104 ) , .ZN( u2_u14_u1_n151 ) );
  NAND2_X1 u2_u14_u1_U66 (.A2( u2_u14_u1_n103 ) , .A1( u2_u14_u1_n105 ) , .ZN( u2_u14_u1_n161 ) );
  INV_X1 u2_u14_u1_U67 (.A( u2_u14_u1_n152 ) , .ZN( u2_u14_u1_n173 ) );
  INV_X1 u2_u14_u1_U68 (.A( u2_u14_u1_n128 ) , .ZN( u2_u14_u1_n172 ) );
  NAND2_X1 u2_u14_u1_U69 (.A2( u2_u14_u1_n102 ) , .A1( u2_u14_u1_n103 ) , .ZN( u2_u14_u1_n123 ) );
  OAI21_X1 u2_u14_u1_U7 (.ZN( u2_u14_u1_n101 ) , .B1( u2_u14_u1_n141 ) , .A( u2_u14_u1_n146 ) , .B2( u2_u14_u1_n183 ) );
  NOR2_X1 u2_u14_u1_U70 (.A2( u2_u14_X_7 ) , .A1( u2_u14_X_8 ) , .ZN( u2_u14_u1_n95 ) );
  NOR2_X1 u2_u14_u1_U71 (.A1( u2_u14_X_12 ) , .A2( u2_u14_X_9 ) , .ZN( u2_u14_u1_n100 ) );
  NOR2_X1 u2_u14_u1_U72 (.A2( u2_u14_X_8 ) , .A1( u2_u14_u1_n177 ) , .ZN( u2_u14_u1_n99 ) );
  NOR2_X1 u2_u14_u1_U73 (.A2( u2_u14_X_12 ) , .ZN( u2_u14_u1_n102 ) , .A1( u2_u14_u1_n176 ) );
  NOR2_X1 u2_u14_u1_U74 (.A2( u2_u14_X_9 ) , .ZN( u2_u14_u1_n105 ) , .A1( u2_u14_u1_n168 ) );
  NAND2_X1 u2_u14_u1_U75 (.A1( u2_u14_X_10 ) , .ZN( u2_u14_u1_n160 ) , .A2( u2_u14_u1_n169 ) );
  NAND2_X1 u2_u14_u1_U76 (.A2( u2_u14_X_10 ) , .A1( u2_u14_X_11 ) , .ZN( u2_u14_u1_n152 ) );
  NAND2_X1 u2_u14_u1_U77 (.A1( u2_u14_X_11 ) , .ZN( u2_u14_u1_n128 ) , .A2( u2_u14_u1_n170 ) );
  AND2_X1 u2_u14_u1_U78 (.A2( u2_u14_X_7 ) , .A1( u2_u14_X_8 ) , .ZN( u2_u14_u1_n104 ) );
  AND2_X1 u2_u14_u1_U79 (.A1( u2_u14_X_8 ) , .ZN( u2_u14_u1_n103 ) , .A2( u2_u14_u1_n177 ) );
  AOI21_X1 u2_u14_u1_U8 (.B2( u2_u14_u1_n155 ) , .B1( u2_u14_u1_n156 ) , .ZN( u2_u14_u1_n157 ) , .A( u2_u14_u1_n174 ) );
  INV_X1 u2_u14_u1_U80 (.A( u2_u14_X_10 ) , .ZN( u2_u14_u1_n170 ) );
  INV_X1 u2_u14_u1_U81 (.A( u2_u14_X_9 ) , .ZN( u2_u14_u1_n176 ) );
  INV_X1 u2_u14_u1_U82 (.A( u2_u14_X_11 ) , .ZN( u2_u14_u1_n169 ) );
  INV_X1 u2_u14_u1_U83 (.A( u2_u14_X_12 ) , .ZN( u2_u14_u1_n168 ) );
  INV_X1 u2_u14_u1_U84 (.A( u2_u14_X_7 ) , .ZN( u2_u14_u1_n177 ) );
  NAND4_X1 u2_u14_u1_U85 (.ZN( u2_out14_28 ) , .A4( u2_u14_u1_n124 ) , .A3( u2_u14_u1_n125 ) , .A2( u2_u14_u1_n126 ) , .A1( u2_u14_u1_n127 ) );
  OAI21_X1 u2_u14_u1_U86 (.ZN( u2_u14_u1_n127 ) , .B2( u2_u14_u1_n139 ) , .B1( u2_u14_u1_n175 ) , .A( u2_u14_u1_n183 ) );
  OAI21_X1 u2_u14_u1_U87 (.ZN( u2_u14_u1_n126 ) , .B2( u2_u14_u1_n140 ) , .A( u2_u14_u1_n146 ) , .B1( u2_u14_u1_n178 ) );
  NAND4_X1 u2_u14_u1_U88 (.ZN( u2_out14_18 ) , .A4( u2_u14_u1_n165 ) , .A3( u2_u14_u1_n166 ) , .A1( u2_u14_u1_n167 ) , .A2( u2_u14_u1_n186 ) );
  AOI22_X1 u2_u14_u1_U89 (.B2( u2_u14_u1_n146 ) , .B1( u2_u14_u1_n147 ) , .A2( u2_u14_u1_n148 ) , .ZN( u2_u14_u1_n166 ) , .A1( u2_u14_u1_n172 ) );
  OR4_X1 u2_u14_u1_U9 (.A4( u2_u14_u1_n106 ) , .A3( u2_u14_u1_n107 ) , .ZN( u2_u14_u1_n108 ) , .A1( u2_u14_u1_n117 ) , .A2( u2_u14_u1_n184 ) );
  INV_X1 u2_u14_u1_U90 (.A( u2_u14_u1_n145 ) , .ZN( u2_u14_u1_n186 ) );
  NAND4_X1 u2_u14_u1_U91 (.ZN( u2_out14_2 ) , .A4( u2_u14_u1_n142 ) , .A3( u2_u14_u1_n143 ) , .A2( u2_u14_u1_n144 ) , .A1( u2_u14_u1_n179 ) );
  OAI21_X1 u2_u14_u1_U92 (.B2( u2_u14_u1_n132 ) , .ZN( u2_u14_u1_n144 ) , .A( u2_u14_u1_n146 ) , .B1( u2_u14_u1_n180 ) );
  INV_X1 u2_u14_u1_U93 (.A( u2_u14_u1_n130 ) , .ZN( u2_u14_u1_n179 ) );
  OR4_X1 u2_u14_u1_U94 (.ZN( u2_out14_13 ) , .A4( u2_u14_u1_n108 ) , .A3( u2_u14_u1_n109 ) , .A2( u2_u14_u1_n110 ) , .A1( u2_u14_u1_n111 ) );
  AOI21_X1 u2_u14_u1_U95 (.ZN( u2_u14_u1_n111 ) , .A( u2_u14_u1_n128 ) , .B2( u2_u14_u1_n131 ) , .B1( u2_u14_u1_n135 ) );
  AOI21_X1 u2_u14_u1_U96 (.ZN( u2_u14_u1_n110 ) , .A( u2_u14_u1_n116 ) , .B1( u2_u14_u1_n152 ) , .B2( u2_u14_u1_n160 ) );
  NAND3_X1 u2_u14_u1_U97 (.A3( u2_u14_u1_n149 ) , .A2( u2_u14_u1_n150 ) , .A1( u2_u14_u1_n151 ) , .ZN( u2_u14_u1_n164 ) );
  NAND3_X1 u2_u14_u1_U98 (.A3( u2_u14_u1_n134 ) , .A2( u2_u14_u1_n135 ) , .ZN( u2_u14_u1_n136 ) , .A1( u2_u14_u1_n151 ) );
  NAND3_X1 u2_u14_u1_U99 (.A1( u2_u14_u1_n133 ) , .ZN( u2_u14_u1_n137 ) , .A2( u2_u14_u1_n154 ) , .A3( u2_u14_u1_n181 ) );
  OAI22_X1 u2_u14_u4_U10 (.B2( u2_u14_u4_n135 ) , .ZN( u2_u14_u4_n137 ) , .B1( u2_u14_u4_n153 ) , .A1( u2_u14_u4_n155 ) , .A2( u2_u14_u4_n171 ) );
  AND3_X1 u2_u14_u4_U11 (.A2( u2_u14_u4_n134 ) , .ZN( u2_u14_u4_n135 ) , .A3( u2_u14_u4_n145 ) , .A1( u2_u14_u4_n157 ) );
  NAND2_X1 u2_u14_u4_U12 (.ZN( u2_u14_u4_n132 ) , .A2( u2_u14_u4_n170 ) , .A1( u2_u14_u4_n173 ) );
  AOI21_X1 u2_u14_u4_U13 (.B2( u2_u14_u4_n160 ) , .B1( u2_u14_u4_n161 ) , .ZN( u2_u14_u4_n162 ) , .A( u2_u14_u4_n170 ) );
  AOI21_X1 u2_u14_u4_U14 (.ZN( u2_u14_u4_n107 ) , .B2( u2_u14_u4_n143 ) , .A( u2_u14_u4_n174 ) , .B1( u2_u14_u4_n184 ) );
  AOI21_X1 u2_u14_u4_U15 (.B2( u2_u14_u4_n158 ) , .B1( u2_u14_u4_n159 ) , .ZN( u2_u14_u4_n163 ) , .A( u2_u14_u4_n174 ) );
  AOI21_X1 u2_u14_u4_U16 (.A( u2_u14_u4_n153 ) , .B2( u2_u14_u4_n154 ) , .B1( u2_u14_u4_n155 ) , .ZN( u2_u14_u4_n165 ) );
  AOI21_X1 u2_u14_u4_U17 (.A( u2_u14_u4_n156 ) , .B2( u2_u14_u4_n157 ) , .ZN( u2_u14_u4_n164 ) , .B1( u2_u14_u4_n184 ) );
  INV_X1 u2_u14_u4_U18 (.A( u2_u14_u4_n138 ) , .ZN( u2_u14_u4_n170 ) );
  AND2_X1 u2_u14_u4_U19 (.A2( u2_u14_u4_n120 ) , .ZN( u2_u14_u4_n155 ) , .A1( u2_u14_u4_n160 ) );
  INV_X1 u2_u14_u4_U20 (.A( u2_u14_u4_n156 ) , .ZN( u2_u14_u4_n175 ) );
  NAND2_X1 u2_u14_u4_U21 (.A2( u2_u14_u4_n118 ) , .ZN( u2_u14_u4_n131 ) , .A1( u2_u14_u4_n147 ) );
  NAND2_X1 u2_u14_u4_U22 (.A1( u2_u14_u4_n119 ) , .A2( u2_u14_u4_n120 ) , .ZN( u2_u14_u4_n130 ) );
  NAND2_X1 u2_u14_u4_U23 (.ZN( u2_u14_u4_n117 ) , .A2( u2_u14_u4_n118 ) , .A1( u2_u14_u4_n148 ) );
  NAND2_X1 u2_u14_u4_U24 (.ZN( u2_u14_u4_n129 ) , .A1( u2_u14_u4_n134 ) , .A2( u2_u14_u4_n148 ) );
  AND3_X1 u2_u14_u4_U25 (.A1( u2_u14_u4_n119 ) , .A2( u2_u14_u4_n143 ) , .A3( u2_u14_u4_n154 ) , .ZN( u2_u14_u4_n161 ) );
  AND2_X1 u2_u14_u4_U26 (.A1( u2_u14_u4_n145 ) , .A2( u2_u14_u4_n147 ) , .ZN( u2_u14_u4_n159 ) );
  OR3_X1 u2_u14_u4_U27 (.A3( u2_u14_u4_n114 ) , .A2( u2_u14_u4_n115 ) , .A1( u2_u14_u4_n116 ) , .ZN( u2_u14_u4_n136 ) );
  AOI21_X1 u2_u14_u4_U28 (.A( u2_u14_u4_n113 ) , .ZN( u2_u14_u4_n116 ) , .B2( u2_u14_u4_n173 ) , .B1( u2_u14_u4_n174 ) );
  AOI21_X1 u2_u14_u4_U29 (.ZN( u2_u14_u4_n115 ) , .B2( u2_u14_u4_n145 ) , .B1( u2_u14_u4_n146 ) , .A( u2_u14_u4_n156 ) );
  NOR2_X1 u2_u14_u4_U3 (.ZN( u2_u14_u4_n121 ) , .A1( u2_u14_u4_n181 ) , .A2( u2_u14_u4_n182 ) );
  OAI22_X1 u2_u14_u4_U30 (.ZN( u2_u14_u4_n114 ) , .A2( u2_u14_u4_n121 ) , .B1( u2_u14_u4_n160 ) , .B2( u2_u14_u4_n170 ) , .A1( u2_u14_u4_n171 ) );
  INV_X1 u2_u14_u4_U31 (.A( u2_u14_u4_n158 ) , .ZN( u2_u14_u4_n182 ) );
  INV_X1 u2_u14_u4_U32 (.ZN( u2_u14_u4_n181 ) , .A( u2_u14_u4_n96 ) );
  INV_X1 u2_u14_u4_U33 (.A( u2_u14_u4_n144 ) , .ZN( u2_u14_u4_n179 ) );
  INV_X1 u2_u14_u4_U34 (.A( u2_u14_u4_n157 ) , .ZN( u2_u14_u4_n178 ) );
  NAND2_X1 u2_u14_u4_U35 (.A2( u2_u14_u4_n154 ) , .A1( u2_u14_u4_n96 ) , .ZN( u2_u14_u4_n97 ) );
  INV_X1 u2_u14_u4_U36 (.ZN( u2_u14_u4_n186 ) , .A( u2_u14_u4_n95 ) );
  OAI221_X1 u2_u14_u4_U37 (.C1( u2_u14_u4_n134 ) , .B1( u2_u14_u4_n158 ) , .B2( u2_u14_u4_n171 ) , .C2( u2_u14_u4_n173 ) , .A( u2_u14_u4_n94 ) , .ZN( u2_u14_u4_n95 ) );
  AOI222_X1 u2_u14_u4_U38 (.B2( u2_u14_u4_n132 ) , .A1( u2_u14_u4_n138 ) , .C2( u2_u14_u4_n175 ) , .A2( u2_u14_u4_n179 ) , .C1( u2_u14_u4_n181 ) , .B1( u2_u14_u4_n185 ) , .ZN( u2_u14_u4_n94 ) );
  INV_X1 u2_u14_u4_U39 (.A( u2_u14_u4_n113 ) , .ZN( u2_u14_u4_n185 ) );
  INV_X1 u2_u14_u4_U4 (.A( u2_u14_u4_n117 ) , .ZN( u2_u14_u4_n184 ) );
  INV_X1 u2_u14_u4_U40 (.A( u2_u14_u4_n143 ) , .ZN( u2_u14_u4_n183 ) );
  NOR2_X1 u2_u14_u4_U41 (.ZN( u2_u14_u4_n138 ) , .A1( u2_u14_u4_n168 ) , .A2( u2_u14_u4_n169 ) );
  NOR2_X1 u2_u14_u4_U42 (.A1( u2_u14_u4_n150 ) , .A2( u2_u14_u4_n152 ) , .ZN( u2_u14_u4_n153 ) );
  NOR2_X1 u2_u14_u4_U43 (.A2( u2_u14_u4_n128 ) , .A1( u2_u14_u4_n138 ) , .ZN( u2_u14_u4_n156 ) );
  AOI22_X1 u2_u14_u4_U44 (.B2( u2_u14_u4_n122 ) , .A1( u2_u14_u4_n123 ) , .ZN( u2_u14_u4_n124 ) , .B1( u2_u14_u4_n128 ) , .A2( u2_u14_u4_n172 ) );
  INV_X1 u2_u14_u4_U45 (.A( u2_u14_u4_n153 ) , .ZN( u2_u14_u4_n172 ) );
  NAND2_X1 u2_u14_u4_U46 (.A2( u2_u14_u4_n120 ) , .ZN( u2_u14_u4_n123 ) , .A1( u2_u14_u4_n161 ) );
  AOI22_X1 u2_u14_u4_U47 (.B2( u2_u14_u4_n132 ) , .A2( u2_u14_u4_n133 ) , .ZN( u2_u14_u4_n140 ) , .A1( u2_u14_u4_n150 ) , .B1( u2_u14_u4_n179 ) );
  NAND2_X1 u2_u14_u4_U48 (.ZN( u2_u14_u4_n133 ) , .A2( u2_u14_u4_n146 ) , .A1( u2_u14_u4_n154 ) );
  NAND2_X1 u2_u14_u4_U49 (.A1( u2_u14_u4_n103 ) , .ZN( u2_u14_u4_n154 ) , .A2( u2_u14_u4_n98 ) );
  NOR4_X1 u2_u14_u4_U5 (.A4( u2_u14_u4_n106 ) , .A3( u2_u14_u4_n107 ) , .A2( u2_u14_u4_n108 ) , .A1( u2_u14_u4_n109 ) , .ZN( u2_u14_u4_n110 ) );
  NAND2_X1 u2_u14_u4_U50 (.A1( u2_u14_u4_n101 ) , .ZN( u2_u14_u4_n158 ) , .A2( u2_u14_u4_n99 ) );
  AOI21_X1 u2_u14_u4_U51 (.ZN( u2_u14_u4_n127 ) , .A( u2_u14_u4_n136 ) , .B2( u2_u14_u4_n150 ) , .B1( u2_u14_u4_n180 ) );
  INV_X1 u2_u14_u4_U52 (.A( u2_u14_u4_n160 ) , .ZN( u2_u14_u4_n180 ) );
  NAND2_X1 u2_u14_u4_U53 (.A2( u2_u14_u4_n104 ) , .A1( u2_u14_u4_n105 ) , .ZN( u2_u14_u4_n146 ) );
  NAND2_X1 u2_u14_u4_U54 (.A2( u2_u14_u4_n101 ) , .A1( u2_u14_u4_n102 ) , .ZN( u2_u14_u4_n160 ) );
  NAND2_X1 u2_u14_u4_U55 (.ZN( u2_u14_u4_n134 ) , .A1( u2_u14_u4_n98 ) , .A2( u2_u14_u4_n99 ) );
  NAND2_X1 u2_u14_u4_U56 (.A1( u2_u14_u4_n103 ) , .A2( u2_u14_u4_n104 ) , .ZN( u2_u14_u4_n143 ) );
  NAND2_X1 u2_u14_u4_U57 (.A2( u2_u14_u4_n105 ) , .ZN( u2_u14_u4_n145 ) , .A1( u2_u14_u4_n98 ) );
  NAND2_X1 u2_u14_u4_U58 (.A1( u2_u14_u4_n100 ) , .A2( u2_u14_u4_n105 ) , .ZN( u2_u14_u4_n120 ) );
  NAND2_X1 u2_u14_u4_U59 (.A1( u2_u14_u4_n102 ) , .A2( u2_u14_u4_n104 ) , .ZN( u2_u14_u4_n148 ) );
  AOI21_X1 u2_u14_u4_U6 (.ZN( u2_u14_u4_n106 ) , .B2( u2_u14_u4_n146 ) , .B1( u2_u14_u4_n158 ) , .A( u2_u14_u4_n170 ) );
  NAND2_X1 u2_u14_u4_U60 (.A2( u2_u14_u4_n100 ) , .A1( u2_u14_u4_n103 ) , .ZN( u2_u14_u4_n157 ) );
  INV_X1 u2_u14_u4_U61 (.A( u2_u14_u4_n150 ) , .ZN( u2_u14_u4_n173 ) );
  INV_X1 u2_u14_u4_U62 (.A( u2_u14_u4_n152 ) , .ZN( u2_u14_u4_n171 ) );
  NAND2_X1 u2_u14_u4_U63 (.A1( u2_u14_u4_n100 ) , .ZN( u2_u14_u4_n118 ) , .A2( u2_u14_u4_n99 ) );
  NAND2_X1 u2_u14_u4_U64 (.A2( u2_u14_u4_n100 ) , .A1( u2_u14_u4_n102 ) , .ZN( u2_u14_u4_n144 ) );
  NAND2_X1 u2_u14_u4_U65 (.A2( u2_u14_u4_n101 ) , .A1( u2_u14_u4_n105 ) , .ZN( u2_u14_u4_n96 ) );
  INV_X1 u2_u14_u4_U66 (.A( u2_u14_u4_n128 ) , .ZN( u2_u14_u4_n174 ) );
  NAND2_X1 u2_u14_u4_U67 (.A2( u2_u14_u4_n102 ) , .ZN( u2_u14_u4_n119 ) , .A1( u2_u14_u4_n98 ) );
  NAND2_X1 u2_u14_u4_U68 (.A2( u2_u14_u4_n101 ) , .A1( u2_u14_u4_n103 ) , .ZN( u2_u14_u4_n147 ) );
  NAND2_X1 u2_u14_u4_U69 (.A2( u2_u14_u4_n104 ) , .ZN( u2_u14_u4_n113 ) , .A1( u2_u14_u4_n99 ) );
  AOI21_X1 u2_u14_u4_U7 (.ZN( u2_u14_u4_n108 ) , .B2( u2_u14_u4_n134 ) , .B1( u2_u14_u4_n155 ) , .A( u2_u14_u4_n156 ) );
  NOR2_X1 u2_u14_u4_U70 (.A2( u2_u14_X_28 ) , .ZN( u2_u14_u4_n150 ) , .A1( u2_u14_u4_n168 ) );
  NOR2_X1 u2_u14_u4_U71 (.A2( u2_u14_X_29 ) , .ZN( u2_u14_u4_n152 ) , .A1( u2_u14_u4_n169 ) );
  NOR2_X1 u2_u14_u4_U72 (.A2( u2_u14_X_30 ) , .ZN( u2_u14_u4_n105 ) , .A1( u2_u14_u4_n176 ) );
  NOR2_X1 u2_u14_u4_U73 (.A2( u2_u14_X_26 ) , .ZN( u2_u14_u4_n100 ) , .A1( u2_u14_u4_n177 ) );
  NOR2_X1 u2_u14_u4_U74 (.A2( u2_u14_X_28 ) , .A1( u2_u14_X_29 ) , .ZN( u2_u14_u4_n128 ) );
  NOR2_X1 u2_u14_u4_U75 (.A2( u2_u14_X_27 ) , .A1( u2_u14_X_30 ) , .ZN( u2_u14_u4_n102 ) );
  NOR2_X1 u2_u14_u4_U76 (.A2( u2_u14_X_25 ) , .A1( u2_u14_X_26 ) , .ZN( u2_u14_u4_n98 ) );
  AND2_X1 u2_u14_u4_U77 (.A2( u2_u14_X_25 ) , .A1( u2_u14_X_26 ) , .ZN( u2_u14_u4_n104 ) );
  AND2_X1 u2_u14_u4_U78 (.A1( u2_u14_X_30 ) , .A2( u2_u14_u4_n176 ) , .ZN( u2_u14_u4_n99 ) );
  AND2_X1 u2_u14_u4_U79 (.A1( u2_u14_X_26 ) , .ZN( u2_u14_u4_n101 ) , .A2( u2_u14_u4_n177 ) );
  AOI21_X1 u2_u14_u4_U8 (.ZN( u2_u14_u4_n109 ) , .A( u2_u14_u4_n153 ) , .B1( u2_u14_u4_n159 ) , .B2( u2_u14_u4_n184 ) );
  AND2_X1 u2_u14_u4_U80 (.A1( u2_u14_X_27 ) , .A2( u2_u14_X_30 ) , .ZN( u2_u14_u4_n103 ) );
  INV_X1 u2_u14_u4_U81 (.A( u2_u14_X_28 ) , .ZN( u2_u14_u4_n169 ) );
  INV_X1 u2_u14_u4_U82 (.A( u2_u14_X_29 ) , .ZN( u2_u14_u4_n168 ) );
  INV_X1 u2_u14_u4_U83 (.A( u2_u14_X_25 ) , .ZN( u2_u14_u4_n177 ) );
  INV_X1 u2_u14_u4_U84 (.A( u2_u14_X_27 ) , .ZN( u2_u14_u4_n176 ) );
  NAND4_X1 u2_u14_u4_U85 (.ZN( u2_out14_25 ) , .A4( u2_u14_u4_n139 ) , .A3( u2_u14_u4_n140 ) , .A2( u2_u14_u4_n141 ) , .A1( u2_u14_u4_n142 ) );
  OAI21_X1 u2_u14_u4_U86 (.A( u2_u14_u4_n128 ) , .B2( u2_u14_u4_n129 ) , .B1( u2_u14_u4_n130 ) , .ZN( u2_u14_u4_n142 ) );
  OAI21_X1 u2_u14_u4_U87 (.B2( u2_u14_u4_n131 ) , .ZN( u2_u14_u4_n141 ) , .A( u2_u14_u4_n175 ) , .B1( u2_u14_u4_n183 ) );
  NAND4_X1 u2_u14_u4_U88 (.ZN( u2_out14_14 ) , .A4( u2_u14_u4_n124 ) , .A3( u2_u14_u4_n125 ) , .A2( u2_u14_u4_n126 ) , .A1( u2_u14_u4_n127 ) );
  AOI22_X1 u2_u14_u4_U89 (.B2( u2_u14_u4_n117 ) , .ZN( u2_u14_u4_n126 ) , .A1( u2_u14_u4_n129 ) , .B1( u2_u14_u4_n152 ) , .A2( u2_u14_u4_n175 ) );
  AOI211_X1 u2_u14_u4_U9 (.B( u2_u14_u4_n136 ) , .A( u2_u14_u4_n137 ) , .C2( u2_u14_u4_n138 ) , .ZN( u2_u14_u4_n139 ) , .C1( u2_u14_u4_n182 ) );
  AOI22_X1 u2_u14_u4_U90 (.ZN( u2_u14_u4_n125 ) , .B2( u2_u14_u4_n131 ) , .A2( u2_u14_u4_n132 ) , .B1( u2_u14_u4_n138 ) , .A1( u2_u14_u4_n178 ) );
  NAND4_X1 u2_u14_u4_U91 (.ZN( u2_out14_8 ) , .A4( u2_u14_u4_n110 ) , .A3( u2_u14_u4_n111 ) , .A2( u2_u14_u4_n112 ) , .A1( u2_u14_u4_n186 ) );
  NAND2_X1 u2_u14_u4_U92 (.ZN( u2_u14_u4_n112 ) , .A2( u2_u14_u4_n130 ) , .A1( u2_u14_u4_n150 ) );
  AOI22_X1 u2_u14_u4_U93 (.ZN( u2_u14_u4_n111 ) , .B2( u2_u14_u4_n132 ) , .A1( u2_u14_u4_n152 ) , .B1( u2_u14_u4_n178 ) , .A2( u2_u14_u4_n97 ) );
  AOI22_X1 u2_u14_u4_U94 (.B2( u2_u14_u4_n149 ) , .B1( u2_u14_u4_n150 ) , .A2( u2_u14_u4_n151 ) , .A1( u2_u14_u4_n152 ) , .ZN( u2_u14_u4_n167 ) );
  NOR4_X1 u2_u14_u4_U95 (.A4( u2_u14_u4_n162 ) , .A3( u2_u14_u4_n163 ) , .A2( u2_u14_u4_n164 ) , .A1( u2_u14_u4_n165 ) , .ZN( u2_u14_u4_n166 ) );
  NAND3_X1 u2_u14_u4_U96 (.ZN( u2_out14_3 ) , .A3( u2_u14_u4_n166 ) , .A1( u2_u14_u4_n167 ) , .A2( u2_u14_u4_n186 ) );
  NAND3_X1 u2_u14_u4_U97 (.A3( u2_u14_u4_n146 ) , .A2( u2_u14_u4_n147 ) , .A1( u2_u14_u4_n148 ) , .ZN( u2_u14_u4_n149 ) );
  NAND3_X1 u2_u14_u4_U98 (.A3( u2_u14_u4_n143 ) , .A2( u2_u14_u4_n144 ) , .A1( u2_u14_u4_n145 ) , .ZN( u2_u14_u4_n151 ) );
  NAND3_X1 u2_u14_u4_U99 (.A3( u2_u14_u4_n121 ) , .ZN( u2_u14_u4_n122 ) , .A2( u2_u14_u4_n144 ) , .A1( u2_u14_u4_n154 ) );
  INV_X1 u2_u14_u5_U10 (.A( u2_u14_u5_n121 ) , .ZN( u2_u14_u5_n177 ) );
  NOR3_X1 u2_u14_u5_U100 (.A3( u2_u14_u5_n141 ) , .A1( u2_u14_u5_n142 ) , .ZN( u2_u14_u5_n143 ) , .A2( u2_u14_u5_n191 ) );
  NAND4_X1 u2_u14_u5_U101 (.ZN( u2_out14_4 ) , .A4( u2_u14_u5_n112 ) , .A2( u2_u14_u5_n113 ) , .A1( u2_u14_u5_n114 ) , .A3( u2_u14_u5_n195 ) );
  AOI211_X1 u2_u14_u5_U102 (.A( u2_u14_u5_n110 ) , .C1( u2_u14_u5_n111 ) , .ZN( u2_u14_u5_n112 ) , .B( u2_u14_u5_n118 ) , .C2( u2_u14_u5_n177 ) );
  AOI222_X1 u2_u14_u5_U103 (.ZN( u2_u14_u5_n113 ) , .A1( u2_u14_u5_n131 ) , .C1( u2_u14_u5_n148 ) , .B2( u2_u14_u5_n174 ) , .C2( u2_u14_u5_n178 ) , .A2( u2_u14_u5_n179 ) , .B1( u2_u14_u5_n99 ) );
  NAND3_X1 u2_u14_u5_U104 (.A2( u2_u14_u5_n154 ) , .A3( u2_u14_u5_n158 ) , .A1( u2_u14_u5_n161 ) , .ZN( u2_u14_u5_n99 ) );
  NOR2_X1 u2_u14_u5_U11 (.ZN( u2_u14_u5_n160 ) , .A2( u2_u14_u5_n173 ) , .A1( u2_u14_u5_n177 ) );
  INV_X1 u2_u14_u5_U12 (.A( u2_u14_u5_n150 ) , .ZN( u2_u14_u5_n174 ) );
  AOI21_X1 u2_u14_u5_U13 (.A( u2_u14_u5_n160 ) , .B2( u2_u14_u5_n161 ) , .ZN( u2_u14_u5_n162 ) , .B1( u2_u14_u5_n192 ) );
  INV_X1 u2_u14_u5_U14 (.A( u2_u14_u5_n159 ) , .ZN( u2_u14_u5_n192 ) );
  AOI21_X1 u2_u14_u5_U15 (.A( u2_u14_u5_n156 ) , .B2( u2_u14_u5_n157 ) , .B1( u2_u14_u5_n158 ) , .ZN( u2_u14_u5_n163 ) );
  AOI21_X1 u2_u14_u5_U16 (.B2( u2_u14_u5_n139 ) , .B1( u2_u14_u5_n140 ) , .ZN( u2_u14_u5_n141 ) , .A( u2_u14_u5_n150 ) );
  OAI21_X1 u2_u14_u5_U17 (.A( u2_u14_u5_n133 ) , .B2( u2_u14_u5_n134 ) , .B1( u2_u14_u5_n135 ) , .ZN( u2_u14_u5_n142 ) );
  OAI21_X1 u2_u14_u5_U18 (.ZN( u2_u14_u5_n133 ) , .B2( u2_u14_u5_n147 ) , .A( u2_u14_u5_n173 ) , .B1( u2_u14_u5_n188 ) );
  NAND2_X1 u2_u14_u5_U19 (.A2( u2_u14_u5_n119 ) , .A1( u2_u14_u5_n123 ) , .ZN( u2_u14_u5_n137 ) );
  INV_X1 u2_u14_u5_U20 (.A( u2_u14_u5_n155 ) , .ZN( u2_u14_u5_n194 ) );
  NAND2_X1 u2_u14_u5_U21 (.A1( u2_u14_u5_n121 ) , .ZN( u2_u14_u5_n132 ) , .A2( u2_u14_u5_n172 ) );
  NAND2_X1 u2_u14_u5_U22 (.A2( u2_u14_u5_n122 ) , .ZN( u2_u14_u5_n136 ) , .A1( u2_u14_u5_n154 ) );
  NAND2_X1 u2_u14_u5_U23 (.A2( u2_u14_u5_n119 ) , .A1( u2_u14_u5_n120 ) , .ZN( u2_u14_u5_n159 ) );
  INV_X1 u2_u14_u5_U24 (.A( u2_u14_u5_n156 ) , .ZN( u2_u14_u5_n175 ) );
  INV_X1 u2_u14_u5_U25 (.A( u2_u14_u5_n158 ) , .ZN( u2_u14_u5_n188 ) );
  INV_X1 u2_u14_u5_U26 (.A( u2_u14_u5_n152 ) , .ZN( u2_u14_u5_n179 ) );
  INV_X1 u2_u14_u5_U27 (.A( u2_u14_u5_n140 ) , .ZN( u2_u14_u5_n182 ) );
  INV_X1 u2_u14_u5_U28 (.A( u2_u14_u5_n151 ) , .ZN( u2_u14_u5_n183 ) );
  INV_X1 u2_u14_u5_U29 (.A( u2_u14_u5_n123 ) , .ZN( u2_u14_u5_n185 ) );
  NOR2_X1 u2_u14_u5_U3 (.ZN( u2_u14_u5_n134 ) , .A1( u2_u14_u5_n183 ) , .A2( u2_u14_u5_n190 ) );
  INV_X1 u2_u14_u5_U30 (.A( u2_u14_u5_n161 ) , .ZN( u2_u14_u5_n184 ) );
  INV_X1 u2_u14_u5_U31 (.A( u2_u14_u5_n139 ) , .ZN( u2_u14_u5_n189 ) );
  INV_X1 u2_u14_u5_U32 (.A( u2_u14_u5_n157 ) , .ZN( u2_u14_u5_n190 ) );
  INV_X1 u2_u14_u5_U33 (.A( u2_u14_u5_n120 ) , .ZN( u2_u14_u5_n193 ) );
  NAND2_X1 u2_u14_u5_U34 (.ZN( u2_u14_u5_n111 ) , .A1( u2_u14_u5_n140 ) , .A2( u2_u14_u5_n155 ) );
  INV_X1 u2_u14_u5_U35 (.A( u2_u14_u5_n117 ) , .ZN( u2_u14_u5_n196 ) );
  OAI221_X1 u2_u14_u5_U36 (.A( u2_u14_u5_n116 ) , .ZN( u2_u14_u5_n117 ) , .B2( u2_u14_u5_n119 ) , .C1( u2_u14_u5_n153 ) , .C2( u2_u14_u5_n158 ) , .B1( u2_u14_u5_n172 ) );
  AOI222_X1 u2_u14_u5_U37 (.ZN( u2_u14_u5_n116 ) , .B2( u2_u14_u5_n145 ) , .C1( u2_u14_u5_n148 ) , .A2( u2_u14_u5_n174 ) , .C2( u2_u14_u5_n177 ) , .B1( u2_u14_u5_n187 ) , .A1( u2_u14_u5_n193 ) );
  INV_X1 u2_u14_u5_U38 (.A( u2_u14_u5_n115 ) , .ZN( u2_u14_u5_n187 ) );
  NOR2_X1 u2_u14_u5_U39 (.ZN( u2_u14_u5_n100 ) , .A1( u2_u14_u5_n170 ) , .A2( u2_u14_u5_n180 ) );
  INV_X1 u2_u14_u5_U4 (.A( u2_u14_u5_n138 ) , .ZN( u2_u14_u5_n191 ) );
  AOI22_X1 u2_u14_u5_U40 (.B2( u2_u14_u5_n131 ) , .A2( u2_u14_u5_n146 ) , .ZN( u2_u14_u5_n169 ) , .B1( u2_u14_u5_n174 ) , .A1( u2_u14_u5_n185 ) );
  NOR2_X1 u2_u14_u5_U41 (.A1( u2_u14_u5_n146 ) , .ZN( u2_u14_u5_n150 ) , .A2( u2_u14_u5_n173 ) );
  AOI21_X1 u2_u14_u5_U42 (.A( u2_u14_u5_n118 ) , .B2( u2_u14_u5_n145 ) , .ZN( u2_u14_u5_n168 ) , .B1( u2_u14_u5_n186 ) );
  INV_X1 u2_u14_u5_U43 (.A( u2_u14_u5_n122 ) , .ZN( u2_u14_u5_n186 ) );
  NOR2_X1 u2_u14_u5_U44 (.A1( u2_u14_u5_n146 ) , .ZN( u2_u14_u5_n152 ) , .A2( u2_u14_u5_n176 ) );
  NOR2_X1 u2_u14_u5_U45 (.A1( u2_u14_u5_n115 ) , .ZN( u2_u14_u5_n118 ) , .A2( u2_u14_u5_n153 ) );
  NOR2_X1 u2_u14_u5_U46 (.A2( u2_u14_u5_n145 ) , .ZN( u2_u14_u5_n156 ) , .A1( u2_u14_u5_n174 ) );
  NOR2_X1 u2_u14_u5_U47 (.ZN( u2_u14_u5_n121 ) , .A2( u2_u14_u5_n145 ) , .A1( u2_u14_u5_n176 ) );
  AOI22_X1 u2_u14_u5_U48 (.ZN( u2_u14_u5_n114 ) , .A2( u2_u14_u5_n137 ) , .A1( u2_u14_u5_n145 ) , .B2( u2_u14_u5_n175 ) , .B1( u2_u14_u5_n193 ) );
  OAI211_X1 u2_u14_u5_U49 (.B( u2_u14_u5_n124 ) , .A( u2_u14_u5_n125 ) , .C2( u2_u14_u5_n126 ) , .C1( u2_u14_u5_n127 ) , .ZN( u2_u14_u5_n128 ) );
  OAI21_X1 u2_u14_u5_U5 (.B2( u2_u14_u5_n136 ) , .B1( u2_u14_u5_n137 ) , .ZN( u2_u14_u5_n138 ) , .A( u2_u14_u5_n177 ) );
  NOR3_X1 u2_u14_u5_U50 (.ZN( u2_u14_u5_n127 ) , .A1( u2_u14_u5_n136 ) , .A3( u2_u14_u5_n148 ) , .A2( u2_u14_u5_n182 ) );
  OAI21_X1 u2_u14_u5_U51 (.ZN( u2_u14_u5_n124 ) , .A( u2_u14_u5_n177 ) , .B2( u2_u14_u5_n183 ) , .B1( u2_u14_u5_n189 ) );
  OAI21_X1 u2_u14_u5_U52 (.ZN( u2_u14_u5_n125 ) , .A( u2_u14_u5_n174 ) , .B2( u2_u14_u5_n185 ) , .B1( u2_u14_u5_n190 ) );
  AOI21_X1 u2_u14_u5_U53 (.A( u2_u14_u5_n153 ) , .B2( u2_u14_u5_n154 ) , .B1( u2_u14_u5_n155 ) , .ZN( u2_u14_u5_n164 ) );
  AOI21_X1 u2_u14_u5_U54 (.ZN( u2_u14_u5_n110 ) , .B1( u2_u14_u5_n122 ) , .B2( u2_u14_u5_n139 ) , .A( u2_u14_u5_n153 ) );
  INV_X1 u2_u14_u5_U55 (.A( u2_u14_u5_n153 ) , .ZN( u2_u14_u5_n176 ) );
  INV_X1 u2_u14_u5_U56 (.A( u2_u14_u5_n126 ) , .ZN( u2_u14_u5_n173 ) );
  AND2_X1 u2_u14_u5_U57 (.A2( u2_u14_u5_n104 ) , .A1( u2_u14_u5_n107 ) , .ZN( u2_u14_u5_n147 ) );
  AND2_X1 u2_u14_u5_U58 (.A2( u2_u14_u5_n104 ) , .A1( u2_u14_u5_n108 ) , .ZN( u2_u14_u5_n148 ) );
  NAND2_X1 u2_u14_u5_U59 (.A1( u2_u14_u5_n105 ) , .A2( u2_u14_u5_n106 ) , .ZN( u2_u14_u5_n158 ) );
  INV_X1 u2_u14_u5_U6 (.A( u2_u14_u5_n135 ) , .ZN( u2_u14_u5_n178 ) );
  NAND2_X1 u2_u14_u5_U60 (.A2( u2_u14_u5_n108 ) , .A1( u2_u14_u5_n109 ) , .ZN( u2_u14_u5_n139 ) );
  NAND2_X1 u2_u14_u5_U61 (.A1( u2_u14_u5_n106 ) , .A2( u2_u14_u5_n108 ) , .ZN( u2_u14_u5_n119 ) );
  NAND2_X1 u2_u14_u5_U62 (.A2( u2_u14_u5_n103 ) , .A1( u2_u14_u5_n105 ) , .ZN( u2_u14_u5_n140 ) );
  NAND2_X1 u2_u14_u5_U63 (.A2( u2_u14_u5_n104 ) , .A1( u2_u14_u5_n105 ) , .ZN( u2_u14_u5_n155 ) );
  NAND2_X1 u2_u14_u5_U64 (.A2( u2_u14_u5_n106 ) , .A1( u2_u14_u5_n107 ) , .ZN( u2_u14_u5_n122 ) );
  NAND2_X1 u2_u14_u5_U65 (.A2( u2_u14_u5_n100 ) , .A1( u2_u14_u5_n106 ) , .ZN( u2_u14_u5_n115 ) );
  NAND2_X1 u2_u14_u5_U66 (.A2( u2_u14_u5_n100 ) , .A1( u2_u14_u5_n103 ) , .ZN( u2_u14_u5_n161 ) );
  NAND2_X1 u2_u14_u5_U67 (.A1( u2_u14_u5_n105 ) , .A2( u2_u14_u5_n109 ) , .ZN( u2_u14_u5_n154 ) );
  INV_X1 u2_u14_u5_U68 (.A( u2_u14_u5_n146 ) , .ZN( u2_u14_u5_n172 ) );
  NAND2_X1 u2_u14_u5_U69 (.A1( u2_u14_u5_n103 ) , .A2( u2_u14_u5_n108 ) , .ZN( u2_u14_u5_n123 ) );
  OAI22_X1 u2_u14_u5_U7 (.B2( u2_u14_u5_n149 ) , .B1( u2_u14_u5_n150 ) , .A2( u2_u14_u5_n151 ) , .A1( u2_u14_u5_n152 ) , .ZN( u2_u14_u5_n165 ) );
  NAND2_X1 u2_u14_u5_U70 (.A2( u2_u14_u5_n103 ) , .A1( u2_u14_u5_n107 ) , .ZN( u2_u14_u5_n151 ) );
  NAND2_X1 u2_u14_u5_U71 (.A2( u2_u14_u5_n107 ) , .A1( u2_u14_u5_n109 ) , .ZN( u2_u14_u5_n120 ) );
  NAND2_X1 u2_u14_u5_U72 (.A2( u2_u14_u5_n100 ) , .A1( u2_u14_u5_n109 ) , .ZN( u2_u14_u5_n157 ) );
  AND2_X1 u2_u14_u5_U73 (.A2( u2_u14_u5_n100 ) , .A1( u2_u14_u5_n104 ) , .ZN( u2_u14_u5_n131 ) );
  INV_X1 u2_u14_u5_U74 (.A( u2_u14_u5_n102 ) , .ZN( u2_u14_u5_n195 ) );
  OAI221_X1 u2_u14_u5_U75 (.A( u2_u14_u5_n101 ) , .ZN( u2_u14_u5_n102 ) , .C2( u2_u14_u5_n115 ) , .C1( u2_u14_u5_n126 ) , .B1( u2_u14_u5_n134 ) , .B2( u2_u14_u5_n160 ) );
  OAI21_X1 u2_u14_u5_U76 (.ZN( u2_u14_u5_n101 ) , .B1( u2_u14_u5_n137 ) , .A( u2_u14_u5_n146 ) , .B2( u2_u14_u5_n147 ) );
  NOR2_X1 u2_u14_u5_U77 (.A2( u2_u14_X_34 ) , .A1( u2_u14_X_35 ) , .ZN( u2_u14_u5_n145 ) );
  NOR2_X1 u2_u14_u5_U78 (.A2( u2_u14_X_34 ) , .ZN( u2_u14_u5_n146 ) , .A1( u2_u14_u5_n171 ) );
  NOR2_X1 u2_u14_u5_U79 (.A2( u2_u14_X_31 ) , .A1( u2_u14_X_32 ) , .ZN( u2_u14_u5_n103 ) );
  NOR3_X1 u2_u14_u5_U8 (.A2( u2_u14_u5_n147 ) , .A1( u2_u14_u5_n148 ) , .ZN( u2_u14_u5_n149 ) , .A3( u2_u14_u5_n194 ) );
  NOR2_X1 u2_u14_u5_U80 (.A2( u2_u14_X_36 ) , .ZN( u2_u14_u5_n105 ) , .A1( u2_u14_u5_n180 ) );
  NOR2_X1 u2_u14_u5_U81 (.A2( u2_u14_X_33 ) , .ZN( u2_u14_u5_n108 ) , .A1( u2_u14_u5_n170 ) );
  NOR2_X1 u2_u14_u5_U82 (.A2( u2_u14_X_33 ) , .A1( u2_u14_X_36 ) , .ZN( u2_u14_u5_n107 ) );
  NOR2_X1 u2_u14_u5_U83 (.A2( u2_u14_X_31 ) , .ZN( u2_u14_u5_n104 ) , .A1( u2_u14_u5_n181 ) );
  NAND2_X1 u2_u14_u5_U84 (.A2( u2_u14_X_34 ) , .A1( u2_u14_X_35 ) , .ZN( u2_u14_u5_n153 ) );
  NAND2_X1 u2_u14_u5_U85 (.A1( u2_u14_X_34 ) , .ZN( u2_u14_u5_n126 ) , .A2( u2_u14_u5_n171 ) );
  AND2_X1 u2_u14_u5_U86 (.A1( u2_u14_X_31 ) , .A2( u2_u14_X_32 ) , .ZN( u2_u14_u5_n106 ) );
  AND2_X1 u2_u14_u5_U87 (.A1( u2_u14_X_31 ) , .ZN( u2_u14_u5_n109 ) , .A2( u2_u14_u5_n181 ) );
  INV_X1 u2_u14_u5_U88 (.A( u2_u14_X_33 ) , .ZN( u2_u14_u5_n180 ) );
  INV_X1 u2_u14_u5_U89 (.A( u2_u14_X_35 ) , .ZN( u2_u14_u5_n171 ) );
  NOR2_X1 u2_u14_u5_U9 (.ZN( u2_u14_u5_n135 ) , .A1( u2_u14_u5_n173 ) , .A2( u2_u14_u5_n176 ) );
  INV_X1 u2_u14_u5_U90 (.A( u2_u14_X_36 ) , .ZN( u2_u14_u5_n170 ) );
  INV_X1 u2_u14_u5_U91 (.A( u2_u14_X_32 ) , .ZN( u2_u14_u5_n181 ) );
  NAND4_X1 u2_u14_u5_U92 (.ZN( u2_out14_29 ) , .A4( u2_u14_u5_n129 ) , .A3( u2_u14_u5_n130 ) , .A2( u2_u14_u5_n168 ) , .A1( u2_u14_u5_n196 ) );
  AOI221_X1 u2_u14_u5_U93 (.A( u2_u14_u5_n128 ) , .ZN( u2_u14_u5_n129 ) , .C2( u2_u14_u5_n132 ) , .B2( u2_u14_u5_n159 ) , .B1( u2_u14_u5_n176 ) , .C1( u2_u14_u5_n184 ) );
  AOI222_X1 u2_u14_u5_U94 (.ZN( u2_u14_u5_n130 ) , .A2( u2_u14_u5_n146 ) , .B1( u2_u14_u5_n147 ) , .C2( u2_u14_u5_n175 ) , .B2( u2_u14_u5_n179 ) , .A1( u2_u14_u5_n188 ) , .C1( u2_u14_u5_n194 ) );
  NAND4_X1 u2_u14_u5_U95 (.ZN( u2_out14_19 ) , .A4( u2_u14_u5_n166 ) , .A3( u2_u14_u5_n167 ) , .A2( u2_u14_u5_n168 ) , .A1( u2_u14_u5_n169 ) );
  AOI22_X1 u2_u14_u5_U96 (.B2( u2_u14_u5_n145 ) , .A2( u2_u14_u5_n146 ) , .ZN( u2_u14_u5_n167 ) , .B1( u2_u14_u5_n182 ) , .A1( u2_u14_u5_n189 ) );
  NOR4_X1 u2_u14_u5_U97 (.A4( u2_u14_u5_n162 ) , .A3( u2_u14_u5_n163 ) , .A2( u2_u14_u5_n164 ) , .A1( u2_u14_u5_n165 ) , .ZN( u2_u14_u5_n166 ) );
  NAND4_X1 u2_u14_u5_U98 (.ZN( u2_out14_11 ) , .A4( u2_u14_u5_n143 ) , .A3( u2_u14_u5_n144 ) , .A2( u2_u14_u5_n169 ) , .A1( u2_u14_u5_n196 ) );
  AOI22_X1 u2_u14_u5_U99 (.A2( u2_u14_u5_n132 ) , .ZN( u2_u14_u5_n144 ) , .B2( u2_u14_u5_n145 ) , .B1( u2_u14_u5_n184 ) , .A1( u2_u14_u5_n194 ) );
  AOI22_X1 u2_u14_u6_U10 (.A2( u2_u14_u6_n151 ) , .B2( u2_u14_u6_n161 ) , .A1( u2_u14_u6_n167 ) , .B1( u2_u14_u6_n170 ) , .ZN( u2_u14_u6_n89 ) );
  AOI21_X1 u2_u14_u6_U11 (.B1( u2_u14_u6_n107 ) , .B2( u2_u14_u6_n132 ) , .A( u2_u14_u6_n158 ) , .ZN( u2_u14_u6_n88 ) );
  AOI21_X1 u2_u14_u6_U12 (.B2( u2_u14_u6_n147 ) , .B1( u2_u14_u6_n148 ) , .ZN( u2_u14_u6_n149 ) , .A( u2_u14_u6_n158 ) );
  AOI21_X1 u2_u14_u6_U13 (.ZN( u2_u14_u6_n106 ) , .A( u2_u14_u6_n142 ) , .B2( u2_u14_u6_n159 ) , .B1( u2_u14_u6_n164 ) );
  INV_X1 u2_u14_u6_U14 (.A( u2_u14_u6_n155 ) , .ZN( u2_u14_u6_n161 ) );
  INV_X1 u2_u14_u6_U15 (.A( u2_u14_u6_n128 ) , .ZN( u2_u14_u6_n164 ) );
  NAND2_X1 u2_u14_u6_U16 (.ZN( u2_u14_u6_n110 ) , .A1( u2_u14_u6_n122 ) , .A2( u2_u14_u6_n129 ) );
  NAND2_X1 u2_u14_u6_U17 (.ZN( u2_u14_u6_n124 ) , .A2( u2_u14_u6_n146 ) , .A1( u2_u14_u6_n148 ) );
  INV_X1 u2_u14_u6_U18 (.A( u2_u14_u6_n132 ) , .ZN( u2_u14_u6_n171 ) );
  AND2_X1 u2_u14_u6_U19 (.A1( u2_u14_u6_n100 ) , .ZN( u2_u14_u6_n130 ) , .A2( u2_u14_u6_n147 ) );
  INV_X1 u2_u14_u6_U20 (.A( u2_u14_u6_n127 ) , .ZN( u2_u14_u6_n173 ) );
  INV_X1 u2_u14_u6_U21 (.A( u2_u14_u6_n121 ) , .ZN( u2_u14_u6_n167 ) );
  INV_X1 u2_u14_u6_U22 (.A( u2_u14_u6_n100 ) , .ZN( u2_u14_u6_n169 ) );
  INV_X1 u2_u14_u6_U23 (.A( u2_u14_u6_n123 ) , .ZN( u2_u14_u6_n170 ) );
  INV_X1 u2_u14_u6_U24 (.A( u2_u14_u6_n113 ) , .ZN( u2_u14_u6_n168 ) );
  AND2_X1 u2_u14_u6_U25 (.A1( u2_u14_u6_n107 ) , .A2( u2_u14_u6_n119 ) , .ZN( u2_u14_u6_n133 ) );
  AND2_X1 u2_u14_u6_U26 (.A2( u2_u14_u6_n121 ) , .A1( u2_u14_u6_n122 ) , .ZN( u2_u14_u6_n131 ) );
  AND3_X1 u2_u14_u6_U27 (.ZN( u2_u14_u6_n120 ) , .A2( u2_u14_u6_n127 ) , .A1( u2_u14_u6_n132 ) , .A3( u2_u14_u6_n145 ) );
  INV_X1 u2_u14_u6_U28 (.A( u2_u14_u6_n146 ) , .ZN( u2_u14_u6_n163 ) );
  AOI222_X1 u2_u14_u6_U29 (.ZN( u2_u14_u6_n114 ) , .A1( u2_u14_u6_n118 ) , .A2( u2_u14_u6_n126 ) , .B2( u2_u14_u6_n151 ) , .C2( u2_u14_u6_n159 ) , .C1( u2_u14_u6_n168 ) , .B1( u2_u14_u6_n169 ) );
  INV_X1 u2_u14_u6_U3 (.A( u2_u14_u6_n110 ) , .ZN( u2_u14_u6_n166 ) );
  NOR2_X1 u2_u14_u6_U30 (.A1( u2_u14_u6_n162 ) , .A2( u2_u14_u6_n165 ) , .ZN( u2_u14_u6_n98 ) );
  NAND2_X1 u2_u14_u6_U31 (.A1( u2_u14_u6_n144 ) , .ZN( u2_u14_u6_n151 ) , .A2( u2_u14_u6_n158 ) );
  NAND2_X1 u2_u14_u6_U32 (.ZN( u2_u14_u6_n132 ) , .A1( u2_u14_u6_n91 ) , .A2( u2_u14_u6_n97 ) );
  AOI22_X1 u2_u14_u6_U33 (.B2( u2_u14_u6_n110 ) , .B1( u2_u14_u6_n111 ) , .A1( u2_u14_u6_n112 ) , .ZN( u2_u14_u6_n115 ) , .A2( u2_u14_u6_n161 ) );
  NAND4_X1 u2_u14_u6_U34 (.A3( u2_u14_u6_n109 ) , .ZN( u2_u14_u6_n112 ) , .A4( u2_u14_u6_n132 ) , .A2( u2_u14_u6_n147 ) , .A1( u2_u14_u6_n166 ) );
  NOR2_X1 u2_u14_u6_U35 (.ZN( u2_u14_u6_n109 ) , .A1( u2_u14_u6_n170 ) , .A2( u2_u14_u6_n173 ) );
  NOR2_X1 u2_u14_u6_U36 (.A2( u2_u14_u6_n126 ) , .ZN( u2_u14_u6_n155 ) , .A1( u2_u14_u6_n160 ) );
  NAND2_X1 u2_u14_u6_U37 (.ZN( u2_u14_u6_n146 ) , .A2( u2_u14_u6_n94 ) , .A1( u2_u14_u6_n99 ) );
  AOI21_X1 u2_u14_u6_U38 (.A( u2_u14_u6_n144 ) , .B2( u2_u14_u6_n145 ) , .B1( u2_u14_u6_n146 ) , .ZN( u2_u14_u6_n150 ) );
  AOI211_X1 u2_u14_u6_U39 (.B( u2_u14_u6_n134 ) , .A( u2_u14_u6_n135 ) , .C1( u2_u14_u6_n136 ) , .ZN( u2_u14_u6_n137 ) , .C2( u2_u14_u6_n151 ) );
  INV_X1 u2_u14_u6_U4 (.A( u2_u14_u6_n142 ) , .ZN( u2_u14_u6_n174 ) );
  AOI21_X1 u2_u14_u6_U40 (.B2( u2_u14_u6_n132 ) , .B1( u2_u14_u6_n133 ) , .ZN( u2_u14_u6_n134 ) , .A( u2_u14_u6_n158 ) );
  NAND4_X1 u2_u14_u6_U41 (.A4( u2_u14_u6_n127 ) , .A3( u2_u14_u6_n128 ) , .A2( u2_u14_u6_n129 ) , .A1( u2_u14_u6_n130 ) , .ZN( u2_u14_u6_n136 ) );
  AOI21_X1 u2_u14_u6_U42 (.B1( u2_u14_u6_n131 ) , .ZN( u2_u14_u6_n135 ) , .A( u2_u14_u6_n144 ) , .B2( u2_u14_u6_n146 ) );
  INV_X1 u2_u14_u6_U43 (.A( u2_u14_u6_n111 ) , .ZN( u2_u14_u6_n158 ) );
  NAND2_X1 u2_u14_u6_U44 (.ZN( u2_u14_u6_n127 ) , .A1( u2_u14_u6_n91 ) , .A2( u2_u14_u6_n92 ) );
  NAND2_X1 u2_u14_u6_U45 (.ZN( u2_u14_u6_n129 ) , .A2( u2_u14_u6_n95 ) , .A1( u2_u14_u6_n96 ) );
  INV_X1 u2_u14_u6_U46 (.A( u2_u14_u6_n144 ) , .ZN( u2_u14_u6_n159 ) );
  NAND2_X1 u2_u14_u6_U47 (.ZN( u2_u14_u6_n145 ) , .A2( u2_u14_u6_n97 ) , .A1( u2_u14_u6_n98 ) );
  NAND2_X1 u2_u14_u6_U48 (.ZN( u2_u14_u6_n148 ) , .A2( u2_u14_u6_n92 ) , .A1( u2_u14_u6_n94 ) );
  NAND2_X1 u2_u14_u6_U49 (.ZN( u2_u14_u6_n108 ) , .A2( u2_u14_u6_n139 ) , .A1( u2_u14_u6_n144 ) );
  NAND2_X1 u2_u14_u6_U5 (.A2( u2_u14_u6_n143 ) , .ZN( u2_u14_u6_n152 ) , .A1( u2_u14_u6_n166 ) );
  NAND2_X1 u2_u14_u6_U50 (.ZN( u2_u14_u6_n121 ) , .A2( u2_u14_u6_n95 ) , .A1( u2_u14_u6_n97 ) );
  NAND2_X1 u2_u14_u6_U51 (.ZN( u2_u14_u6_n107 ) , .A2( u2_u14_u6_n92 ) , .A1( u2_u14_u6_n95 ) );
  AND2_X1 u2_u14_u6_U52 (.ZN( u2_u14_u6_n118 ) , .A2( u2_u14_u6_n91 ) , .A1( u2_u14_u6_n99 ) );
  NAND2_X1 u2_u14_u6_U53 (.ZN( u2_u14_u6_n147 ) , .A2( u2_u14_u6_n98 ) , .A1( u2_u14_u6_n99 ) );
  NAND2_X1 u2_u14_u6_U54 (.ZN( u2_u14_u6_n128 ) , .A1( u2_u14_u6_n94 ) , .A2( u2_u14_u6_n96 ) );
  NAND2_X1 u2_u14_u6_U55 (.ZN( u2_u14_u6_n119 ) , .A2( u2_u14_u6_n95 ) , .A1( u2_u14_u6_n99 ) );
  NAND2_X1 u2_u14_u6_U56 (.ZN( u2_u14_u6_n123 ) , .A2( u2_u14_u6_n91 ) , .A1( u2_u14_u6_n96 ) );
  NAND2_X1 u2_u14_u6_U57 (.ZN( u2_u14_u6_n100 ) , .A2( u2_u14_u6_n92 ) , .A1( u2_u14_u6_n98 ) );
  NAND2_X1 u2_u14_u6_U58 (.ZN( u2_u14_u6_n122 ) , .A1( u2_u14_u6_n94 ) , .A2( u2_u14_u6_n97 ) );
  INV_X1 u2_u14_u6_U59 (.A( u2_u14_u6_n139 ) , .ZN( u2_u14_u6_n160 ) );
  AOI22_X1 u2_u14_u6_U6 (.B2( u2_u14_u6_n101 ) , .A1( u2_u14_u6_n102 ) , .ZN( u2_u14_u6_n103 ) , .B1( u2_u14_u6_n160 ) , .A2( u2_u14_u6_n161 ) );
  NAND2_X1 u2_u14_u6_U60 (.ZN( u2_u14_u6_n113 ) , .A1( u2_u14_u6_n96 ) , .A2( u2_u14_u6_n98 ) );
  NOR2_X1 u2_u14_u6_U61 (.A2( u2_u14_X_40 ) , .A1( u2_u14_X_41 ) , .ZN( u2_u14_u6_n126 ) );
  NOR2_X1 u2_u14_u6_U62 (.A2( u2_u14_X_39 ) , .A1( u2_u14_X_42 ) , .ZN( u2_u14_u6_n92 ) );
  NOR2_X1 u2_u14_u6_U63 (.A2( u2_u14_X_39 ) , .A1( u2_u14_u6_n156 ) , .ZN( u2_u14_u6_n97 ) );
  NOR2_X1 u2_u14_u6_U64 (.A2( u2_u14_X_38 ) , .A1( u2_u14_u6_n165 ) , .ZN( u2_u14_u6_n95 ) );
  NOR2_X1 u2_u14_u6_U65 (.A2( u2_u14_X_41 ) , .ZN( u2_u14_u6_n111 ) , .A1( u2_u14_u6_n157 ) );
  NOR2_X1 u2_u14_u6_U66 (.A2( u2_u14_X_37 ) , .A1( u2_u14_u6_n162 ) , .ZN( u2_u14_u6_n94 ) );
  NOR2_X1 u2_u14_u6_U67 (.A2( u2_u14_X_37 ) , .A1( u2_u14_X_38 ) , .ZN( u2_u14_u6_n91 ) );
  NAND2_X1 u2_u14_u6_U68 (.A1( u2_u14_X_41 ) , .ZN( u2_u14_u6_n144 ) , .A2( u2_u14_u6_n157 ) );
  NAND2_X1 u2_u14_u6_U69 (.A2( u2_u14_X_40 ) , .A1( u2_u14_X_41 ) , .ZN( u2_u14_u6_n139 ) );
  NOR2_X1 u2_u14_u6_U7 (.A1( u2_u14_u6_n118 ) , .ZN( u2_u14_u6_n143 ) , .A2( u2_u14_u6_n168 ) );
  AND2_X1 u2_u14_u6_U70 (.A1( u2_u14_X_39 ) , .A2( u2_u14_u6_n156 ) , .ZN( u2_u14_u6_n96 ) );
  AND2_X1 u2_u14_u6_U71 (.A1( u2_u14_X_39 ) , .A2( u2_u14_X_42 ) , .ZN( u2_u14_u6_n99 ) );
  INV_X1 u2_u14_u6_U72 (.A( u2_u14_X_40 ) , .ZN( u2_u14_u6_n157 ) );
  INV_X1 u2_u14_u6_U73 (.A( u2_u14_X_37 ) , .ZN( u2_u14_u6_n165 ) );
  INV_X1 u2_u14_u6_U74 (.A( u2_u14_X_38 ) , .ZN( u2_u14_u6_n162 ) );
  INV_X1 u2_u14_u6_U75 (.A( u2_u14_X_42 ) , .ZN( u2_u14_u6_n156 ) );
  NAND4_X1 u2_u14_u6_U76 (.ZN( u2_out14_32 ) , .A4( u2_u14_u6_n103 ) , .A3( u2_u14_u6_n104 ) , .A2( u2_u14_u6_n105 ) , .A1( u2_u14_u6_n106 ) );
  AOI22_X1 u2_u14_u6_U77 (.ZN( u2_u14_u6_n105 ) , .A2( u2_u14_u6_n108 ) , .A1( u2_u14_u6_n118 ) , .B2( u2_u14_u6_n126 ) , .B1( u2_u14_u6_n171 ) );
  AOI22_X1 u2_u14_u6_U78 (.ZN( u2_u14_u6_n104 ) , .A1( u2_u14_u6_n111 ) , .B1( u2_u14_u6_n124 ) , .B2( u2_u14_u6_n151 ) , .A2( u2_u14_u6_n93 ) );
  NAND4_X1 u2_u14_u6_U79 (.ZN( u2_out14_12 ) , .A4( u2_u14_u6_n114 ) , .A3( u2_u14_u6_n115 ) , .A2( u2_u14_u6_n116 ) , .A1( u2_u14_u6_n117 ) );
  INV_X1 u2_u14_u6_U8 (.ZN( u2_u14_u6_n172 ) , .A( u2_u14_u6_n88 ) );
  OAI22_X1 u2_u14_u6_U80 (.B2( u2_u14_u6_n111 ) , .ZN( u2_u14_u6_n116 ) , .B1( u2_u14_u6_n126 ) , .A2( u2_u14_u6_n164 ) , .A1( u2_u14_u6_n167 ) );
  OAI21_X1 u2_u14_u6_U81 (.A( u2_u14_u6_n108 ) , .ZN( u2_u14_u6_n117 ) , .B2( u2_u14_u6_n141 ) , .B1( u2_u14_u6_n163 ) );
  OAI211_X1 u2_u14_u6_U82 (.ZN( u2_out14_22 ) , .B( u2_u14_u6_n137 ) , .A( u2_u14_u6_n138 ) , .C2( u2_u14_u6_n139 ) , .C1( u2_u14_u6_n140 ) );
  AOI22_X1 u2_u14_u6_U83 (.B1( u2_u14_u6_n124 ) , .A2( u2_u14_u6_n125 ) , .A1( u2_u14_u6_n126 ) , .ZN( u2_u14_u6_n138 ) , .B2( u2_u14_u6_n161 ) );
  AND4_X1 u2_u14_u6_U84 (.A3( u2_u14_u6_n119 ) , .A1( u2_u14_u6_n120 ) , .A4( u2_u14_u6_n129 ) , .ZN( u2_u14_u6_n140 ) , .A2( u2_u14_u6_n143 ) );
  OAI211_X1 u2_u14_u6_U85 (.ZN( u2_out14_7 ) , .B( u2_u14_u6_n153 ) , .C2( u2_u14_u6_n154 ) , .C1( u2_u14_u6_n155 ) , .A( u2_u14_u6_n174 ) );
  NOR3_X1 u2_u14_u6_U86 (.A1( u2_u14_u6_n141 ) , .ZN( u2_u14_u6_n154 ) , .A3( u2_u14_u6_n164 ) , .A2( u2_u14_u6_n171 ) );
  AOI211_X1 u2_u14_u6_U87 (.B( u2_u14_u6_n149 ) , .A( u2_u14_u6_n150 ) , .C2( u2_u14_u6_n151 ) , .C1( u2_u14_u6_n152 ) , .ZN( u2_u14_u6_n153 ) );
  NAND3_X1 u2_u14_u6_U88 (.A2( u2_u14_u6_n123 ) , .ZN( u2_u14_u6_n125 ) , .A1( u2_u14_u6_n130 ) , .A3( u2_u14_u6_n131 ) );
  NAND3_X1 u2_u14_u6_U89 (.A3( u2_u14_u6_n133 ) , .ZN( u2_u14_u6_n141 ) , .A1( u2_u14_u6_n145 ) , .A2( u2_u14_u6_n148 ) );
  OAI21_X1 u2_u14_u6_U9 (.A( u2_u14_u6_n159 ) , .B1( u2_u14_u6_n169 ) , .B2( u2_u14_u6_n173 ) , .ZN( u2_u14_u6_n90 ) );
  NAND3_X1 u2_u14_u6_U90 (.ZN( u2_u14_u6_n101 ) , .A3( u2_u14_u6_n107 ) , .A2( u2_u14_u6_n121 ) , .A1( u2_u14_u6_n127 ) );
  NAND3_X1 u2_u14_u6_U91 (.ZN( u2_u14_u6_n102 ) , .A3( u2_u14_u6_n130 ) , .A2( u2_u14_u6_n145 ) , .A1( u2_u14_u6_n166 ) );
  NAND3_X1 u2_u14_u6_U92 (.A3( u2_u14_u6_n113 ) , .A1( u2_u14_u6_n119 ) , .A2( u2_u14_u6_n123 ) , .ZN( u2_u14_u6_n93 ) );
  NAND3_X1 u2_u14_u6_U93 (.ZN( u2_u14_u6_n142 ) , .A2( u2_u14_u6_n172 ) , .A3( u2_u14_u6_n89 ) , .A1( u2_u14_u6_n90 ) );
  XOR2_X1 u2_u15_U10 (.A( u2_FP_62 ) , .B( u2_K16_45 ) , .Z( u2_u15_X_45 ) );
  XOR2_X1 u2_u15_U11 (.A( u2_FP_61 ) , .B( u2_K16_44 ) , .Z( u2_u15_X_44 ) );
  XOR2_X1 u2_u15_U12 (.A( u2_FP_60 ) , .B( u2_K16_43 ) , .Z( u2_u15_X_43 ) );
  XOR2_X1 u2_u15_U13 (.A( u2_FP_61 ) , .B( u2_K16_42 ) , .Z( u2_u15_X_42 ) );
  XOR2_X1 u2_u15_U14 (.A( u2_FP_60 ) , .B( u2_K16_41 ) , .Z( u2_u15_X_41 ) );
  XOR2_X1 u2_u15_U15 (.A( u2_FP_59 ) , .B( u2_K16_40 ) , .Z( u2_u15_X_40 ) );
  XOR2_X1 u2_u15_U16 (.A( u2_FP_34 ) , .B( u2_K16_3 ) , .Z( u2_u15_X_3 ) );
  XOR2_X1 u2_u15_U17 (.A( u2_FP_58 ) , .B( u2_K16_39 ) , .Z( u2_u15_X_39 ) );
  XOR2_X1 u2_u15_U18 (.A( u2_FP_57 ) , .B( u2_K16_38 ) , .Z( u2_u15_X_38 ) );
  XOR2_X1 u2_u15_U19 (.A( u2_FP_56 ) , .B( u2_K16_37 ) , .Z( u2_u15_X_37 ) );
  XOR2_X1 u2_u15_U20 (.A( u2_FP_57 ) , .B( u2_K16_36 ) , .Z( u2_u15_X_36 ) );
  XOR2_X1 u2_u15_U21 (.A( u2_FP_56 ) , .B( u2_K16_35 ) , .Z( u2_u15_X_35 ) );
  XOR2_X1 u2_u15_U22 (.A( u2_FP_55 ) , .B( u2_K16_34 ) , .Z( u2_u15_X_34 ) );
  XOR2_X1 u2_u15_U23 (.A( u2_FP_54 ) , .B( u2_K16_33 ) , .Z( u2_u15_X_33 ) );
  XOR2_X1 u2_u15_U24 (.A( u2_FP_53 ) , .B( u2_K16_32 ) , .Z( u2_u15_X_32 ) );
  XOR2_X1 u2_u15_U25 (.A( u2_FP_52 ) , .B( u2_K16_31 ) , .Z( u2_u15_X_31 ) );
  XOR2_X1 u2_u15_U26 (.A( u2_FP_53 ) , .B( u2_K16_30 ) , .Z( u2_u15_X_30 ) );
  XOR2_X1 u2_u15_U27 (.A( u2_FP_33 ) , .B( u2_K16_2 ) , .Z( u2_u15_X_2 ) );
  XOR2_X1 u2_u15_U28 (.A( u2_FP_52 ) , .B( u2_K16_29 ) , .Z( u2_u15_X_29 ) );
  XOR2_X1 u2_u15_U29 (.A( u2_FP_51 ) , .B( u2_K16_28 ) , .Z( u2_u15_X_28 ) );
  XOR2_X1 u2_u15_U30 (.A( u2_FP_50 ) , .B( u2_K16_27 ) , .Z( u2_u15_X_27 ) );
  XOR2_X1 u2_u15_U31 (.A( u2_FP_49 ) , .B( u2_K16_26 ) , .Z( u2_u15_X_26 ) );
  XOR2_X1 u2_u15_U32 (.A( u2_FP_48 ) , .B( u2_K16_25 ) , .Z( u2_u15_X_25 ) );
  XOR2_X1 u2_u15_U38 (.A( u2_FP_64 ) , .B( u2_K16_1 ) , .Z( u2_u15_X_1 ) );
  XOR2_X1 u2_u15_U4 (.A( u2_FP_37 ) , .B( u2_K16_6 ) , .Z( u2_u15_X_6 ) );
  XOR2_X1 u2_u15_U5 (.A( u2_FP_36 ) , .B( u2_K16_5 ) , .Z( u2_u15_X_5 ) );
  XOR2_X1 u2_u15_U6 (.A( u2_FP_35 ) , .B( u2_K16_4 ) , .Z( u2_u15_X_4 ) );
  XOR2_X1 u2_u15_U7 (.A( u2_FP_33 ) , .B( u2_K16_48 ) , .Z( u2_u15_X_48 ) );
  XOR2_X1 u2_u15_U8 (.A( u2_FP_64 ) , .B( u2_K16_47 ) , .Z( u2_u15_X_47 ) );
  XOR2_X1 u2_u15_U9 (.A( u2_FP_63 ) , .B( u2_K16_46 ) , .Z( u2_u15_X_46 ) );
  AND3_X1 u2_u15_u0_U10 (.A2( u2_u15_u0_n112 ) , .ZN( u2_u15_u0_n127 ) , .A3( u2_u15_u0_n130 ) , .A1( u2_u15_u0_n148 ) );
  NAND2_X1 u2_u15_u0_U11 (.ZN( u2_u15_u0_n113 ) , .A1( u2_u15_u0_n139 ) , .A2( u2_u15_u0_n149 ) );
  AND2_X1 u2_u15_u0_U12 (.ZN( u2_u15_u0_n107 ) , .A1( u2_u15_u0_n130 ) , .A2( u2_u15_u0_n140 ) );
  AND2_X1 u2_u15_u0_U13 (.A2( u2_u15_u0_n129 ) , .A1( u2_u15_u0_n130 ) , .ZN( u2_u15_u0_n151 ) );
  AND2_X1 u2_u15_u0_U14 (.A1( u2_u15_u0_n108 ) , .A2( u2_u15_u0_n125 ) , .ZN( u2_u15_u0_n145 ) );
  INV_X1 u2_u15_u0_U15 (.A( u2_u15_u0_n143 ) , .ZN( u2_u15_u0_n173 ) );
  NOR2_X1 u2_u15_u0_U16 (.A2( u2_u15_u0_n136 ) , .ZN( u2_u15_u0_n147 ) , .A1( u2_u15_u0_n160 ) );
  AOI21_X1 u2_u15_u0_U17 (.B1( u2_u15_u0_n103 ) , .ZN( u2_u15_u0_n132 ) , .A( u2_u15_u0_n165 ) , .B2( u2_u15_u0_n93 ) );
  INV_X1 u2_u15_u0_U18 (.A( u2_u15_u0_n142 ) , .ZN( u2_u15_u0_n165 ) );
  OAI221_X1 u2_u15_u0_U19 (.C1( u2_u15_u0_n112 ) , .ZN( u2_u15_u0_n120 ) , .B1( u2_u15_u0_n138 ) , .B2( u2_u15_u0_n141 ) , .C2( u2_u15_u0_n147 ) , .A( u2_u15_u0_n172 ) );
  AOI211_X1 u2_u15_u0_U20 (.B( u2_u15_u0_n115 ) , .A( u2_u15_u0_n116 ) , .C2( u2_u15_u0_n117 ) , .C1( u2_u15_u0_n118 ) , .ZN( u2_u15_u0_n119 ) );
  OAI22_X1 u2_u15_u0_U21 (.B1( u2_u15_u0_n125 ) , .ZN( u2_u15_u0_n126 ) , .A1( u2_u15_u0_n138 ) , .A2( u2_u15_u0_n146 ) , .B2( u2_u15_u0_n147 ) );
  OAI22_X1 u2_u15_u0_U22 (.B1( u2_u15_u0_n131 ) , .A1( u2_u15_u0_n144 ) , .B2( u2_u15_u0_n147 ) , .A2( u2_u15_u0_n90 ) , .ZN( u2_u15_u0_n91 ) );
  AND3_X1 u2_u15_u0_U23 (.A3( u2_u15_u0_n121 ) , .A2( u2_u15_u0_n125 ) , .A1( u2_u15_u0_n148 ) , .ZN( u2_u15_u0_n90 ) );
  INV_X1 u2_u15_u0_U24 (.A( u2_u15_u0_n136 ) , .ZN( u2_u15_u0_n161 ) );
  AOI22_X1 u2_u15_u0_U25 (.B2( u2_u15_u0_n109 ) , .A2( u2_u15_u0_n110 ) , .ZN( u2_u15_u0_n111 ) , .B1( u2_u15_u0_n118 ) , .A1( u2_u15_u0_n160 ) );
  INV_X1 u2_u15_u0_U26 (.A( u2_u15_u0_n118 ) , .ZN( u2_u15_u0_n158 ) );
  AOI21_X1 u2_u15_u0_U27 (.ZN( u2_u15_u0_n104 ) , .B1( u2_u15_u0_n107 ) , .B2( u2_u15_u0_n141 ) , .A( u2_u15_u0_n144 ) );
  AOI21_X1 u2_u15_u0_U28 (.B1( u2_u15_u0_n127 ) , .B2( u2_u15_u0_n129 ) , .A( u2_u15_u0_n138 ) , .ZN( u2_u15_u0_n96 ) );
  AOI21_X1 u2_u15_u0_U29 (.ZN( u2_u15_u0_n116 ) , .B2( u2_u15_u0_n142 ) , .A( u2_u15_u0_n144 ) , .B1( u2_u15_u0_n166 ) );
  INV_X1 u2_u15_u0_U3 (.A( u2_u15_u0_n113 ) , .ZN( u2_u15_u0_n166 ) );
  NAND2_X1 u2_u15_u0_U30 (.A1( u2_u15_u0_n100 ) , .A2( u2_u15_u0_n103 ) , .ZN( u2_u15_u0_n125 ) );
  NAND2_X1 u2_u15_u0_U31 (.A2( u2_u15_u0_n103 ) , .ZN( u2_u15_u0_n140 ) , .A1( u2_u15_u0_n94 ) );
  NAND2_X1 u2_u15_u0_U32 (.A1( u2_u15_u0_n101 ) , .A2( u2_u15_u0_n102 ) , .ZN( u2_u15_u0_n150 ) );
  INV_X1 u2_u15_u0_U33 (.A( u2_u15_u0_n138 ) , .ZN( u2_u15_u0_n160 ) );
  NAND2_X1 u2_u15_u0_U34 (.A2( u2_u15_u0_n102 ) , .A1( u2_u15_u0_n103 ) , .ZN( u2_u15_u0_n149 ) );
  NAND2_X1 u2_u15_u0_U35 (.A2( u2_u15_u0_n100 ) , .A1( u2_u15_u0_n101 ) , .ZN( u2_u15_u0_n139 ) );
  NAND2_X1 u2_u15_u0_U36 (.A2( u2_u15_u0_n100 ) , .ZN( u2_u15_u0_n131 ) , .A1( u2_u15_u0_n92 ) );
  NAND2_X1 u2_u15_u0_U37 (.ZN( u2_u15_u0_n108 ) , .A1( u2_u15_u0_n92 ) , .A2( u2_u15_u0_n94 ) );
  NAND2_X1 u2_u15_u0_U38 (.A2( u2_u15_u0_n102 ) , .ZN( u2_u15_u0_n114 ) , .A1( u2_u15_u0_n92 ) );
  NAND2_X1 u2_u15_u0_U39 (.A1( u2_u15_u0_n101 ) , .ZN( u2_u15_u0_n130 ) , .A2( u2_u15_u0_n94 ) );
  AOI21_X1 u2_u15_u0_U4 (.B1( u2_u15_u0_n114 ) , .ZN( u2_u15_u0_n115 ) , .B2( u2_u15_u0_n129 ) , .A( u2_u15_u0_n161 ) );
  NAND2_X1 u2_u15_u0_U40 (.A2( u2_u15_u0_n101 ) , .ZN( u2_u15_u0_n121 ) , .A1( u2_u15_u0_n93 ) );
  INV_X1 u2_u15_u0_U41 (.ZN( u2_u15_u0_n172 ) , .A( u2_u15_u0_n88 ) );
  OAI222_X1 u2_u15_u0_U42 (.C1( u2_u15_u0_n108 ) , .A1( u2_u15_u0_n125 ) , .B2( u2_u15_u0_n128 ) , .B1( u2_u15_u0_n144 ) , .A2( u2_u15_u0_n158 ) , .C2( u2_u15_u0_n161 ) , .ZN( u2_u15_u0_n88 ) );
  NAND2_X1 u2_u15_u0_U43 (.ZN( u2_u15_u0_n112 ) , .A2( u2_u15_u0_n92 ) , .A1( u2_u15_u0_n93 ) );
  OR3_X1 u2_u15_u0_U44 (.A3( u2_u15_u0_n152 ) , .A2( u2_u15_u0_n153 ) , .A1( u2_u15_u0_n154 ) , .ZN( u2_u15_u0_n155 ) );
  AOI21_X1 u2_u15_u0_U45 (.B2( u2_u15_u0_n150 ) , .B1( u2_u15_u0_n151 ) , .ZN( u2_u15_u0_n152 ) , .A( u2_u15_u0_n158 ) );
  AOI21_X1 u2_u15_u0_U46 (.A( u2_u15_u0_n144 ) , .B2( u2_u15_u0_n145 ) , .B1( u2_u15_u0_n146 ) , .ZN( u2_u15_u0_n154 ) );
  AOI21_X1 u2_u15_u0_U47 (.A( u2_u15_u0_n147 ) , .B2( u2_u15_u0_n148 ) , .B1( u2_u15_u0_n149 ) , .ZN( u2_u15_u0_n153 ) );
  INV_X1 u2_u15_u0_U48 (.ZN( u2_u15_u0_n171 ) , .A( u2_u15_u0_n99 ) );
  OAI211_X1 u2_u15_u0_U49 (.C2( u2_u15_u0_n140 ) , .C1( u2_u15_u0_n161 ) , .A( u2_u15_u0_n169 ) , .B( u2_u15_u0_n98 ) , .ZN( u2_u15_u0_n99 ) );
  AOI21_X1 u2_u15_u0_U5 (.B2( u2_u15_u0_n131 ) , .ZN( u2_u15_u0_n134 ) , .B1( u2_u15_u0_n151 ) , .A( u2_u15_u0_n158 ) );
  AOI211_X1 u2_u15_u0_U50 (.C1( u2_u15_u0_n118 ) , .A( u2_u15_u0_n123 ) , .B( u2_u15_u0_n96 ) , .C2( u2_u15_u0_n97 ) , .ZN( u2_u15_u0_n98 ) );
  INV_X1 u2_u15_u0_U51 (.ZN( u2_u15_u0_n169 ) , .A( u2_u15_u0_n91 ) );
  NOR2_X1 u2_u15_u0_U52 (.A2( u2_u15_X_2 ) , .ZN( u2_u15_u0_n103 ) , .A1( u2_u15_u0_n164 ) );
  NOR2_X1 u2_u15_u0_U53 (.A2( u2_u15_X_4 ) , .A1( u2_u15_X_5 ) , .ZN( u2_u15_u0_n118 ) );
  NOR2_X1 u2_u15_u0_U54 (.A2( u2_u15_X_1 ) , .A1( u2_u15_X_2 ) , .ZN( u2_u15_u0_n92 ) );
  NOR2_X1 u2_u15_u0_U55 (.A2( u2_u15_X_1 ) , .ZN( u2_u15_u0_n101 ) , .A1( u2_u15_u0_n163 ) );
  NOR2_X1 u2_u15_u0_U56 (.A2( u2_u15_X_3 ) , .A1( u2_u15_X_6 ) , .ZN( u2_u15_u0_n94 ) );
  NOR2_X1 u2_u15_u0_U57 (.A2( u2_u15_X_6 ) , .ZN( u2_u15_u0_n100 ) , .A1( u2_u15_u0_n162 ) );
  NAND2_X1 u2_u15_u0_U58 (.A2( u2_u15_X_4 ) , .A1( u2_u15_X_5 ) , .ZN( u2_u15_u0_n144 ) );
  NOR2_X1 u2_u15_u0_U59 (.A2( u2_u15_X_5 ) , .ZN( u2_u15_u0_n136 ) , .A1( u2_u15_u0_n159 ) );
  NOR2_X1 u2_u15_u0_U6 (.A1( u2_u15_u0_n108 ) , .ZN( u2_u15_u0_n123 ) , .A2( u2_u15_u0_n158 ) );
  NAND2_X1 u2_u15_u0_U60 (.A1( u2_u15_X_5 ) , .ZN( u2_u15_u0_n138 ) , .A2( u2_u15_u0_n159 ) );
  AND2_X1 u2_u15_u0_U61 (.A2( u2_u15_X_3 ) , .A1( u2_u15_X_6 ) , .ZN( u2_u15_u0_n102 ) );
  AND2_X1 u2_u15_u0_U62 (.A1( u2_u15_X_6 ) , .A2( u2_u15_u0_n162 ) , .ZN( u2_u15_u0_n93 ) );
  INV_X1 u2_u15_u0_U63 (.A( u2_u15_X_4 ) , .ZN( u2_u15_u0_n159 ) );
  INV_X1 u2_u15_u0_U64 (.A( u2_u15_X_1 ) , .ZN( u2_u15_u0_n164 ) );
  INV_X1 u2_u15_u0_U65 (.A( u2_u15_X_2 ) , .ZN( u2_u15_u0_n163 ) );
  INV_X1 u2_u15_u0_U66 (.A( u2_u15_X_3 ) , .ZN( u2_u15_u0_n162 ) );
  INV_X1 u2_u15_u0_U67 (.A( u2_u15_u0_n126 ) , .ZN( u2_u15_u0_n168 ) );
  AOI211_X1 u2_u15_u0_U68 (.B( u2_u15_u0_n133 ) , .A( u2_u15_u0_n134 ) , .C2( u2_u15_u0_n135 ) , .C1( u2_u15_u0_n136 ) , .ZN( u2_u15_u0_n137 ) );
  OR4_X1 u2_u15_u0_U69 (.ZN( u2_out15_17 ) , .A4( u2_u15_u0_n122 ) , .A2( u2_u15_u0_n123 ) , .A1( u2_u15_u0_n124 ) , .A3( u2_u15_u0_n170 ) );
  OAI21_X1 u2_u15_u0_U7 (.B1( u2_u15_u0_n150 ) , .B2( u2_u15_u0_n158 ) , .A( u2_u15_u0_n172 ) , .ZN( u2_u15_u0_n89 ) );
  AOI21_X1 u2_u15_u0_U70 (.B2( u2_u15_u0_n107 ) , .ZN( u2_u15_u0_n124 ) , .B1( u2_u15_u0_n128 ) , .A( u2_u15_u0_n161 ) );
  INV_X1 u2_u15_u0_U71 (.A( u2_u15_u0_n111 ) , .ZN( u2_u15_u0_n170 ) );
  OR4_X1 u2_u15_u0_U72 (.ZN( u2_out15_31 ) , .A4( u2_u15_u0_n155 ) , .A2( u2_u15_u0_n156 ) , .A1( u2_u15_u0_n157 ) , .A3( u2_u15_u0_n173 ) );
  AOI21_X1 u2_u15_u0_U73 (.A( u2_u15_u0_n138 ) , .B2( u2_u15_u0_n139 ) , .B1( u2_u15_u0_n140 ) , .ZN( u2_u15_u0_n157 ) );
  AOI21_X1 u2_u15_u0_U74 (.B2( u2_u15_u0_n141 ) , .B1( u2_u15_u0_n142 ) , .ZN( u2_u15_u0_n156 ) , .A( u2_u15_u0_n161 ) );
  INV_X1 u2_u15_u0_U75 (.ZN( u2_u15_u0_n174 ) , .A( u2_u15_u0_n89 ) );
  AOI211_X1 u2_u15_u0_U76 (.B( u2_u15_u0_n104 ) , .A( u2_u15_u0_n105 ) , .ZN( u2_u15_u0_n106 ) , .C2( u2_u15_u0_n113 ) , .C1( u2_u15_u0_n160 ) );
  NOR2_X1 u2_u15_u0_U77 (.A1( u2_u15_u0_n163 ) , .A2( u2_u15_u0_n164 ) , .ZN( u2_u15_u0_n95 ) );
  OAI221_X1 u2_u15_u0_U78 (.C1( u2_u15_u0_n121 ) , .ZN( u2_u15_u0_n122 ) , .B2( u2_u15_u0_n127 ) , .A( u2_u15_u0_n143 ) , .B1( u2_u15_u0_n144 ) , .C2( u2_u15_u0_n147 ) );
  NOR2_X1 u2_u15_u0_U79 (.A1( u2_u15_u0_n120 ) , .ZN( u2_u15_u0_n143 ) , .A2( u2_u15_u0_n167 ) );
  AND2_X1 u2_u15_u0_U8 (.A1( u2_u15_u0_n114 ) , .A2( u2_u15_u0_n121 ) , .ZN( u2_u15_u0_n146 ) );
  AOI21_X1 u2_u15_u0_U80 (.B1( u2_u15_u0_n132 ) , .ZN( u2_u15_u0_n133 ) , .A( u2_u15_u0_n144 ) , .B2( u2_u15_u0_n166 ) );
  OAI22_X1 u2_u15_u0_U81 (.ZN( u2_u15_u0_n105 ) , .A2( u2_u15_u0_n132 ) , .B1( u2_u15_u0_n146 ) , .A1( u2_u15_u0_n147 ) , .B2( u2_u15_u0_n161 ) );
  NAND2_X1 u2_u15_u0_U82 (.ZN( u2_u15_u0_n110 ) , .A2( u2_u15_u0_n132 ) , .A1( u2_u15_u0_n145 ) );
  INV_X1 u2_u15_u0_U83 (.A( u2_u15_u0_n119 ) , .ZN( u2_u15_u0_n167 ) );
  NAND2_X1 u2_u15_u0_U84 (.ZN( u2_u15_u0_n148 ) , .A1( u2_u15_u0_n93 ) , .A2( u2_u15_u0_n95 ) );
  NAND2_X1 u2_u15_u0_U85 (.A1( u2_u15_u0_n100 ) , .ZN( u2_u15_u0_n129 ) , .A2( u2_u15_u0_n95 ) );
  NAND2_X1 u2_u15_u0_U86 (.A1( u2_u15_u0_n102 ) , .ZN( u2_u15_u0_n128 ) , .A2( u2_u15_u0_n95 ) );
  NAND2_X1 u2_u15_u0_U87 (.ZN( u2_u15_u0_n142 ) , .A1( u2_u15_u0_n94 ) , .A2( u2_u15_u0_n95 ) );
  NAND3_X1 u2_u15_u0_U88 (.ZN( u2_out15_23 ) , .A3( u2_u15_u0_n137 ) , .A1( u2_u15_u0_n168 ) , .A2( u2_u15_u0_n171 ) );
  NAND3_X1 u2_u15_u0_U89 (.A3( u2_u15_u0_n127 ) , .A2( u2_u15_u0_n128 ) , .ZN( u2_u15_u0_n135 ) , .A1( u2_u15_u0_n150 ) );
  AND2_X1 u2_u15_u0_U9 (.A1( u2_u15_u0_n131 ) , .ZN( u2_u15_u0_n141 ) , .A2( u2_u15_u0_n150 ) );
  NAND3_X1 u2_u15_u0_U90 (.ZN( u2_u15_u0_n117 ) , .A3( u2_u15_u0_n132 ) , .A2( u2_u15_u0_n139 ) , .A1( u2_u15_u0_n148 ) );
  NAND3_X1 u2_u15_u0_U91 (.ZN( u2_u15_u0_n109 ) , .A2( u2_u15_u0_n114 ) , .A3( u2_u15_u0_n140 ) , .A1( u2_u15_u0_n149 ) );
  NAND3_X1 u2_u15_u0_U92 (.ZN( u2_out15_9 ) , .A3( u2_u15_u0_n106 ) , .A2( u2_u15_u0_n171 ) , .A1( u2_u15_u0_n174 ) );
  NAND3_X1 u2_u15_u0_U93 (.A2( u2_u15_u0_n128 ) , .A1( u2_u15_u0_n132 ) , .A3( u2_u15_u0_n146 ) , .ZN( u2_u15_u0_n97 ) );
  OAI22_X1 u2_u15_u4_U10 (.B2( u2_u15_u4_n135 ) , .ZN( u2_u15_u4_n137 ) , .B1( u2_u15_u4_n153 ) , .A1( u2_u15_u4_n155 ) , .A2( u2_u15_u4_n171 ) );
  AND3_X1 u2_u15_u4_U11 (.A2( u2_u15_u4_n134 ) , .ZN( u2_u15_u4_n135 ) , .A3( u2_u15_u4_n145 ) , .A1( u2_u15_u4_n157 ) );
  OR3_X1 u2_u15_u4_U12 (.A3( u2_u15_u4_n114 ) , .A2( u2_u15_u4_n115 ) , .A1( u2_u15_u4_n116 ) , .ZN( u2_u15_u4_n136 ) );
  AOI21_X1 u2_u15_u4_U13 (.A( u2_u15_u4_n113 ) , .ZN( u2_u15_u4_n116 ) , .B2( u2_u15_u4_n173 ) , .B1( u2_u15_u4_n174 ) );
  AOI21_X1 u2_u15_u4_U14 (.ZN( u2_u15_u4_n115 ) , .B2( u2_u15_u4_n145 ) , .B1( u2_u15_u4_n146 ) , .A( u2_u15_u4_n156 ) );
  OAI22_X1 u2_u15_u4_U15 (.ZN( u2_u15_u4_n114 ) , .A2( u2_u15_u4_n121 ) , .B1( u2_u15_u4_n160 ) , .B2( u2_u15_u4_n170 ) , .A1( u2_u15_u4_n171 ) );
  NAND2_X1 u2_u15_u4_U16 (.ZN( u2_u15_u4_n132 ) , .A2( u2_u15_u4_n170 ) , .A1( u2_u15_u4_n173 ) );
  AOI21_X1 u2_u15_u4_U17 (.B2( u2_u15_u4_n160 ) , .B1( u2_u15_u4_n161 ) , .ZN( u2_u15_u4_n162 ) , .A( u2_u15_u4_n170 ) );
  AOI21_X1 u2_u15_u4_U18 (.ZN( u2_u15_u4_n107 ) , .B2( u2_u15_u4_n143 ) , .A( u2_u15_u4_n174 ) , .B1( u2_u15_u4_n184 ) );
  AOI21_X1 u2_u15_u4_U19 (.B2( u2_u15_u4_n158 ) , .B1( u2_u15_u4_n159 ) , .ZN( u2_u15_u4_n163 ) , .A( u2_u15_u4_n174 ) );
  AOI21_X1 u2_u15_u4_U20 (.A( u2_u15_u4_n153 ) , .B2( u2_u15_u4_n154 ) , .B1( u2_u15_u4_n155 ) , .ZN( u2_u15_u4_n165 ) );
  AOI21_X1 u2_u15_u4_U21 (.A( u2_u15_u4_n156 ) , .B2( u2_u15_u4_n157 ) , .ZN( u2_u15_u4_n164 ) , .B1( u2_u15_u4_n184 ) );
  INV_X1 u2_u15_u4_U22 (.A( u2_u15_u4_n138 ) , .ZN( u2_u15_u4_n170 ) );
  AND2_X1 u2_u15_u4_U23 (.A2( u2_u15_u4_n120 ) , .ZN( u2_u15_u4_n155 ) , .A1( u2_u15_u4_n160 ) );
  INV_X1 u2_u15_u4_U24 (.A( u2_u15_u4_n156 ) , .ZN( u2_u15_u4_n175 ) );
  NAND2_X1 u2_u15_u4_U25 (.A2( u2_u15_u4_n118 ) , .ZN( u2_u15_u4_n131 ) , .A1( u2_u15_u4_n147 ) );
  NAND2_X1 u2_u15_u4_U26 (.A1( u2_u15_u4_n119 ) , .A2( u2_u15_u4_n120 ) , .ZN( u2_u15_u4_n130 ) );
  NAND2_X1 u2_u15_u4_U27 (.ZN( u2_u15_u4_n117 ) , .A2( u2_u15_u4_n118 ) , .A1( u2_u15_u4_n148 ) );
  NAND2_X1 u2_u15_u4_U28 (.ZN( u2_u15_u4_n129 ) , .A1( u2_u15_u4_n134 ) , .A2( u2_u15_u4_n148 ) );
  AND3_X1 u2_u15_u4_U29 (.A1( u2_u15_u4_n119 ) , .A2( u2_u15_u4_n143 ) , .A3( u2_u15_u4_n154 ) , .ZN( u2_u15_u4_n161 ) );
  NOR2_X1 u2_u15_u4_U3 (.ZN( u2_u15_u4_n121 ) , .A1( u2_u15_u4_n181 ) , .A2( u2_u15_u4_n182 ) );
  AND2_X1 u2_u15_u4_U30 (.A1( u2_u15_u4_n145 ) , .A2( u2_u15_u4_n147 ) , .ZN( u2_u15_u4_n159 ) );
  INV_X1 u2_u15_u4_U31 (.A( u2_u15_u4_n158 ) , .ZN( u2_u15_u4_n182 ) );
  INV_X1 u2_u15_u4_U32 (.ZN( u2_u15_u4_n181 ) , .A( u2_u15_u4_n96 ) );
  INV_X1 u2_u15_u4_U33 (.A( u2_u15_u4_n144 ) , .ZN( u2_u15_u4_n179 ) );
  INV_X1 u2_u15_u4_U34 (.A( u2_u15_u4_n157 ) , .ZN( u2_u15_u4_n178 ) );
  NAND2_X1 u2_u15_u4_U35 (.A2( u2_u15_u4_n154 ) , .A1( u2_u15_u4_n96 ) , .ZN( u2_u15_u4_n97 ) );
  INV_X1 u2_u15_u4_U36 (.ZN( u2_u15_u4_n186 ) , .A( u2_u15_u4_n95 ) );
  OAI221_X1 u2_u15_u4_U37 (.C1( u2_u15_u4_n134 ) , .B1( u2_u15_u4_n158 ) , .B2( u2_u15_u4_n171 ) , .C2( u2_u15_u4_n173 ) , .A( u2_u15_u4_n94 ) , .ZN( u2_u15_u4_n95 ) );
  AOI222_X1 u2_u15_u4_U38 (.B2( u2_u15_u4_n132 ) , .A1( u2_u15_u4_n138 ) , .C2( u2_u15_u4_n175 ) , .A2( u2_u15_u4_n179 ) , .C1( u2_u15_u4_n181 ) , .B1( u2_u15_u4_n185 ) , .ZN( u2_u15_u4_n94 ) );
  INV_X1 u2_u15_u4_U39 (.A( u2_u15_u4_n113 ) , .ZN( u2_u15_u4_n185 ) );
  INV_X1 u2_u15_u4_U4 (.A( u2_u15_u4_n117 ) , .ZN( u2_u15_u4_n184 ) );
  INV_X1 u2_u15_u4_U40 (.A( u2_u15_u4_n143 ) , .ZN( u2_u15_u4_n183 ) );
  NOR2_X1 u2_u15_u4_U41 (.ZN( u2_u15_u4_n138 ) , .A1( u2_u15_u4_n168 ) , .A2( u2_u15_u4_n169 ) );
  NOR2_X1 u2_u15_u4_U42 (.A1( u2_u15_u4_n150 ) , .A2( u2_u15_u4_n152 ) , .ZN( u2_u15_u4_n153 ) );
  NOR2_X1 u2_u15_u4_U43 (.A2( u2_u15_u4_n128 ) , .A1( u2_u15_u4_n138 ) , .ZN( u2_u15_u4_n156 ) );
  AOI22_X1 u2_u15_u4_U44 (.B2( u2_u15_u4_n122 ) , .A1( u2_u15_u4_n123 ) , .ZN( u2_u15_u4_n124 ) , .B1( u2_u15_u4_n128 ) , .A2( u2_u15_u4_n172 ) );
  NAND2_X1 u2_u15_u4_U45 (.A2( u2_u15_u4_n120 ) , .ZN( u2_u15_u4_n123 ) , .A1( u2_u15_u4_n161 ) );
  INV_X1 u2_u15_u4_U46 (.A( u2_u15_u4_n153 ) , .ZN( u2_u15_u4_n172 ) );
  AOI22_X1 u2_u15_u4_U47 (.B2( u2_u15_u4_n132 ) , .A2( u2_u15_u4_n133 ) , .ZN( u2_u15_u4_n140 ) , .A1( u2_u15_u4_n150 ) , .B1( u2_u15_u4_n179 ) );
  NAND2_X1 u2_u15_u4_U48 (.ZN( u2_u15_u4_n133 ) , .A2( u2_u15_u4_n146 ) , .A1( u2_u15_u4_n154 ) );
  NAND2_X1 u2_u15_u4_U49 (.A1( u2_u15_u4_n103 ) , .ZN( u2_u15_u4_n154 ) , .A2( u2_u15_u4_n98 ) );
  NOR4_X1 u2_u15_u4_U5 (.A4( u2_u15_u4_n106 ) , .A3( u2_u15_u4_n107 ) , .A2( u2_u15_u4_n108 ) , .A1( u2_u15_u4_n109 ) , .ZN( u2_u15_u4_n110 ) );
  NAND2_X1 u2_u15_u4_U50 (.A1( u2_u15_u4_n101 ) , .ZN( u2_u15_u4_n158 ) , .A2( u2_u15_u4_n99 ) );
  AOI21_X1 u2_u15_u4_U51 (.ZN( u2_u15_u4_n127 ) , .A( u2_u15_u4_n136 ) , .B2( u2_u15_u4_n150 ) , .B1( u2_u15_u4_n180 ) );
  INV_X1 u2_u15_u4_U52 (.A( u2_u15_u4_n160 ) , .ZN( u2_u15_u4_n180 ) );
  NAND2_X1 u2_u15_u4_U53 (.A2( u2_u15_u4_n104 ) , .A1( u2_u15_u4_n105 ) , .ZN( u2_u15_u4_n146 ) );
  NAND2_X1 u2_u15_u4_U54 (.A2( u2_u15_u4_n101 ) , .A1( u2_u15_u4_n102 ) , .ZN( u2_u15_u4_n160 ) );
  NAND2_X1 u2_u15_u4_U55 (.ZN( u2_u15_u4_n134 ) , .A1( u2_u15_u4_n98 ) , .A2( u2_u15_u4_n99 ) );
  NAND2_X1 u2_u15_u4_U56 (.A1( u2_u15_u4_n103 ) , .A2( u2_u15_u4_n104 ) , .ZN( u2_u15_u4_n143 ) );
  NAND2_X1 u2_u15_u4_U57 (.A2( u2_u15_u4_n105 ) , .ZN( u2_u15_u4_n145 ) , .A1( u2_u15_u4_n98 ) );
  NAND2_X1 u2_u15_u4_U58 (.A1( u2_u15_u4_n100 ) , .A2( u2_u15_u4_n105 ) , .ZN( u2_u15_u4_n120 ) );
  NAND2_X1 u2_u15_u4_U59 (.A1( u2_u15_u4_n102 ) , .A2( u2_u15_u4_n104 ) , .ZN( u2_u15_u4_n148 ) );
  AOI21_X1 u2_u15_u4_U6 (.ZN( u2_u15_u4_n106 ) , .B2( u2_u15_u4_n146 ) , .B1( u2_u15_u4_n158 ) , .A( u2_u15_u4_n170 ) );
  NAND2_X1 u2_u15_u4_U60 (.A2( u2_u15_u4_n100 ) , .A1( u2_u15_u4_n103 ) , .ZN( u2_u15_u4_n157 ) );
  INV_X1 u2_u15_u4_U61 (.A( u2_u15_u4_n150 ) , .ZN( u2_u15_u4_n173 ) );
  INV_X1 u2_u15_u4_U62 (.A( u2_u15_u4_n152 ) , .ZN( u2_u15_u4_n171 ) );
  NAND2_X1 u2_u15_u4_U63 (.A1( u2_u15_u4_n100 ) , .ZN( u2_u15_u4_n118 ) , .A2( u2_u15_u4_n99 ) );
  NAND2_X1 u2_u15_u4_U64 (.A2( u2_u15_u4_n100 ) , .A1( u2_u15_u4_n102 ) , .ZN( u2_u15_u4_n144 ) );
  NAND2_X1 u2_u15_u4_U65 (.A2( u2_u15_u4_n101 ) , .A1( u2_u15_u4_n105 ) , .ZN( u2_u15_u4_n96 ) );
  INV_X1 u2_u15_u4_U66 (.A( u2_u15_u4_n128 ) , .ZN( u2_u15_u4_n174 ) );
  NAND2_X1 u2_u15_u4_U67 (.A2( u2_u15_u4_n102 ) , .ZN( u2_u15_u4_n119 ) , .A1( u2_u15_u4_n98 ) );
  NAND2_X1 u2_u15_u4_U68 (.A2( u2_u15_u4_n101 ) , .A1( u2_u15_u4_n103 ) , .ZN( u2_u15_u4_n147 ) );
  NAND2_X1 u2_u15_u4_U69 (.A2( u2_u15_u4_n104 ) , .ZN( u2_u15_u4_n113 ) , .A1( u2_u15_u4_n99 ) );
  AOI21_X1 u2_u15_u4_U7 (.ZN( u2_u15_u4_n108 ) , .B2( u2_u15_u4_n134 ) , .B1( u2_u15_u4_n155 ) , .A( u2_u15_u4_n156 ) );
  NOR2_X1 u2_u15_u4_U70 (.A2( u2_u15_X_28 ) , .ZN( u2_u15_u4_n150 ) , .A1( u2_u15_u4_n168 ) );
  NOR2_X1 u2_u15_u4_U71 (.A2( u2_u15_X_29 ) , .ZN( u2_u15_u4_n152 ) , .A1( u2_u15_u4_n169 ) );
  NOR2_X1 u2_u15_u4_U72 (.A2( u2_u15_X_26 ) , .ZN( u2_u15_u4_n100 ) , .A1( u2_u15_u4_n177 ) );
  NOR2_X1 u2_u15_u4_U73 (.A2( u2_u15_X_30 ) , .ZN( u2_u15_u4_n105 ) , .A1( u2_u15_u4_n176 ) );
  NOR2_X1 u2_u15_u4_U74 (.A2( u2_u15_X_28 ) , .A1( u2_u15_X_29 ) , .ZN( u2_u15_u4_n128 ) );
  NOR2_X1 u2_u15_u4_U75 (.A2( u2_u15_X_25 ) , .A1( u2_u15_X_26 ) , .ZN( u2_u15_u4_n98 ) );
  NOR2_X1 u2_u15_u4_U76 (.A2( u2_u15_X_27 ) , .A1( u2_u15_X_30 ) , .ZN( u2_u15_u4_n102 ) );
  AND2_X1 u2_u15_u4_U77 (.A2( u2_u15_X_25 ) , .A1( u2_u15_X_26 ) , .ZN( u2_u15_u4_n104 ) );
  AND2_X1 u2_u15_u4_U78 (.A1( u2_u15_X_30 ) , .A2( u2_u15_u4_n176 ) , .ZN( u2_u15_u4_n99 ) );
  AND2_X1 u2_u15_u4_U79 (.A1( u2_u15_X_26 ) , .ZN( u2_u15_u4_n101 ) , .A2( u2_u15_u4_n177 ) );
  AOI21_X1 u2_u15_u4_U8 (.ZN( u2_u15_u4_n109 ) , .A( u2_u15_u4_n153 ) , .B1( u2_u15_u4_n159 ) , .B2( u2_u15_u4_n184 ) );
  AND2_X1 u2_u15_u4_U80 (.A1( u2_u15_X_27 ) , .A2( u2_u15_X_30 ) , .ZN( u2_u15_u4_n103 ) );
  INV_X1 u2_u15_u4_U81 (.A( u2_u15_X_28 ) , .ZN( u2_u15_u4_n169 ) );
  INV_X1 u2_u15_u4_U82 (.A( u2_u15_X_29 ) , .ZN( u2_u15_u4_n168 ) );
  INV_X1 u2_u15_u4_U83 (.A( u2_u15_X_25 ) , .ZN( u2_u15_u4_n177 ) );
  INV_X1 u2_u15_u4_U84 (.A( u2_u15_X_27 ) , .ZN( u2_u15_u4_n176 ) );
  NAND4_X1 u2_u15_u4_U85 (.ZN( u2_out15_14 ) , .A4( u2_u15_u4_n124 ) , .A3( u2_u15_u4_n125 ) , .A2( u2_u15_u4_n126 ) , .A1( u2_u15_u4_n127 ) );
  AOI22_X1 u2_u15_u4_U86 (.B2( u2_u15_u4_n117 ) , .ZN( u2_u15_u4_n126 ) , .A1( u2_u15_u4_n129 ) , .B1( u2_u15_u4_n152 ) , .A2( u2_u15_u4_n175 ) );
  AOI22_X1 u2_u15_u4_U87 (.ZN( u2_u15_u4_n125 ) , .B2( u2_u15_u4_n131 ) , .A2( u2_u15_u4_n132 ) , .B1( u2_u15_u4_n138 ) , .A1( u2_u15_u4_n178 ) );
  AOI22_X1 u2_u15_u4_U88 (.B2( u2_u15_u4_n149 ) , .B1( u2_u15_u4_n150 ) , .A2( u2_u15_u4_n151 ) , .A1( u2_u15_u4_n152 ) , .ZN( u2_u15_u4_n167 ) );
  NOR4_X1 u2_u15_u4_U89 (.A4( u2_u15_u4_n162 ) , .A3( u2_u15_u4_n163 ) , .A2( u2_u15_u4_n164 ) , .A1( u2_u15_u4_n165 ) , .ZN( u2_u15_u4_n166 ) );
  AOI211_X1 u2_u15_u4_U9 (.B( u2_u15_u4_n136 ) , .A( u2_u15_u4_n137 ) , .C2( u2_u15_u4_n138 ) , .ZN( u2_u15_u4_n139 ) , .C1( u2_u15_u4_n182 ) );
  NAND4_X1 u2_u15_u4_U90 (.ZN( u2_out15_8 ) , .A4( u2_u15_u4_n110 ) , .A3( u2_u15_u4_n111 ) , .A2( u2_u15_u4_n112 ) , .A1( u2_u15_u4_n186 ) );
  NAND2_X1 u2_u15_u4_U91 (.ZN( u2_u15_u4_n112 ) , .A2( u2_u15_u4_n130 ) , .A1( u2_u15_u4_n150 ) );
  AOI22_X1 u2_u15_u4_U92 (.ZN( u2_u15_u4_n111 ) , .B2( u2_u15_u4_n132 ) , .A1( u2_u15_u4_n152 ) , .B1( u2_u15_u4_n178 ) , .A2( u2_u15_u4_n97 ) );
  NAND4_X1 u2_u15_u4_U93 (.ZN( u2_out15_25 ) , .A4( u2_u15_u4_n139 ) , .A3( u2_u15_u4_n140 ) , .A2( u2_u15_u4_n141 ) , .A1( u2_u15_u4_n142 ) );
  OAI21_X1 u2_u15_u4_U94 (.A( u2_u15_u4_n128 ) , .B2( u2_u15_u4_n129 ) , .B1( u2_u15_u4_n130 ) , .ZN( u2_u15_u4_n142 ) );
  OAI21_X1 u2_u15_u4_U95 (.B2( u2_u15_u4_n131 ) , .ZN( u2_u15_u4_n141 ) , .A( u2_u15_u4_n175 ) , .B1( u2_u15_u4_n183 ) );
  NAND3_X1 u2_u15_u4_U96 (.ZN( u2_out15_3 ) , .A3( u2_u15_u4_n166 ) , .A1( u2_u15_u4_n167 ) , .A2( u2_u15_u4_n186 ) );
  NAND3_X1 u2_u15_u4_U97 (.A3( u2_u15_u4_n146 ) , .A2( u2_u15_u4_n147 ) , .A1( u2_u15_u4_n148 ) , .ZN( u2_u15_u4_n149 ) );
  NAND3_X1 u2_u15_u4_U98 (.A3( u2_u15_u4_n143 ) , .A2( u2_u15_u4_n144 ) , .A1( u2_u15_u4_n145 ) , .ZN( u2_u15_u4_n151 ) );
  NAND3_X1 u2_u15_u4_U99 (.A3( u2_u15_u4_n121 ) , .ZN( u2_u15_u4_n122 ) , .A2( u2_u15_u4_n144 ) , .A1( u2_u15_u4_n154 ) );
  INV_X1 u2_u15_u5_U10 (.A( u2_u15_u5_n121 ) , .ZN( u2_u15_u5_n177 ) );
  AOI222_X1 u2_u15_u5_U100 (.ZN( u2_u15_u5_n113 ) , .A1( u2_u15_u5_n131 ) , .C1( u2_u15_u5_n148 ) , .B2( u2_u15_u5_n174 ) , .C2( u2_u15_u5_n178 ) , .A2( u2_u15_u5_n179 ) , .B1( u2_u15_u5_n99 ) );
  NAND4_X1 u2_u15_u5_U101 (.ZN( u2_out15_29 ) , .A4( u2_u15_u5_n129 ) , .A3( u2_u15_u5_n130 ) , .A2( u2_u15_u5_n168 ) , .A1( u2_u15_u5_n196 ) );
  AOI221_X1 u2_u15_u5_U102 (.A( u2_u15_u5_n128 ) , .ZN( u2_u15_u5_n129 ) , .C2( u2_u15_u5_n132 ) , .B2( u2_u15_u5_n159 ) , .B1( u2_u15_u5_n176 ) , .C1( u2_u15_u5_n184 ) );
  AOI222_X1 u2_u15_u5_U103 (.ZN( u2_u15_u5_n130 ) , .A2( u2_u15_u5_n146 ) , .B1( u2_u15_u5_n147 ) , .C2( u2_u15_u5_n175 ) , .B2( u2_u15_u5_n179 ) , .A1( u2_u15_u5_n188 ) , .C1( u2_u15_u5_n194 ) );
  NAND3_X1 u2_u15_u5_U104 (.A2( u2_u15_u5_n154 ) , .A3( u2_u15_u5_n158 ) , .A1( u2_u15_u5_n161 ) , .ZN( u2_u15_u5_n99 ) );
  NOR2_X1 u2_u15_u5_U11 (.ZN( u2_u15_u5_n160 ) , .A2( u2_u15_u5_n173 ) , .A1( u2_u15_u5_n177 ) );
  INV_X1 u2_u15_u5_U12 (.A( u2_u15_u5_n150 ) , .ZN( u2_u15_u5_n174 ) );
  AOI21_X1 u2_u15_u5_U13 (.A( u2_u15_u5_n160 ) , .B2( u2_u15_u5_n161 ) , .ZN( u2_u15_u5_n162 ) , .B1( u2_u15_u5_n192 ) );
  INV_X1 u2_u15_u5_U14 (.A( u2_u15_u5_n159 ) , .ZN( u2_u15_u5_n192 ) );
  AOI21_X1 u2_u15_u5_U15 (.A( u2_u15_u5_n156 ) , .B2( u2_u15_u5_n157 ) , .B1( u2_u15_u5_n158 ) , .ZN( u2_u15_u5_n163 ) );
  AOI21_X1 u2_u15_u5_U16 (.B2( u2_u15_u5_n139 ) , .B1( u2_u15_u5_n140 ) , .ZN( u2_u15_u5_n141 ) , .A( u2_u15_u5_n150 ) );
  OAI21_X1 u2_u15_u5_U17 (.A( u2_u15_u5_n133 ) , .B2( u2_u15_u5_n134 ) , .B1( u2_u15_u5_n135 ) , .ZN( u2_u15_u5_n142 ) );
  OAI21_X1 u2_u15_u5_U18 (.ZN( u2_u15_u5_n133 ) , .B2( u2_u15_u5_n147 ) , .A( u2_u15_u5_n173 ) , .B1( u2_u15_u5_n188 ) );
  NAND2_X1 u2_u15_u5_U19 (.A2( u2_u15_u5_n119 ) , .A1( u2_u15_u5_n123 ) , .ZN( u2_u15_u5_n137 ) );
  INV_X1 u2_u15_u5_U20 (.A( u2_u15_u5_n155 ) , .ZN( u2_u15_u5_n194 ) );
  NAND2_X1 u2_u15_u5_U21 (.A1( u2_u15_u5_n121 ) , .ZN( u2_u15_u5_n132 ) , .A2( u2_u15_u5_n172 ) );
  NAND2_X1 u2_u15_u5_U22 (.A2( u2_u15_u5_n122 ) , .ZN( u2_u15_u5_n136 ) , .A1( u2_u15_u5_n154 ) );
  NAND2_X1 u2_u15_u5_U23 (.A2( u2_u15_u5_n119 ) , .A1( u2_u15_u5_n120 ) , .ZN( u2_u15_u5_n159 ) );
  INV_X1 u2_u15_u5_U24 (.A( u2_u15_u5_n156 ) , .ZN( u2_u15_u5_n175 ) );
  INV_X1 u2_u15_u5_U25 (.A( u2_u15_u5_n158 ) , .ZN( u2_u15_u5_n188 ) );
  INV_X1 u2_u15_u5_U26 (.A( u2_u15_u5_n152 ) , .ZN( u2_u15_u5_n179 ) );
  INV_X1 u2_u15_u5_U27 (.A( u2_u15_u5_n140 ) , .ZN( u2_u15_u5_n182 ) );
  INV_X1 u2_u15_u5_U28 (.A( u2_u15_u5_n151 ) , .ZN( u2_u15_u5_n183 ) );
  INV_X1 u2_u15_u5_U29 (.A( u2_u15_u5_n123 ) , .ZN( u2_u15_u5_n185 ) );
  NOR2_X1 u2_u15_u5_U3 (.ZN( u2_u15_u5_n134 ) , .A1( u2_u15_u5_n183 ) , .A2( u2_u15_u5_n190 ) );
  INV_X1 u2_u15_u5_U30 (.A( u2_u15_u5_n161 ) , .ZN( u2_u15_u5_n184 ) );
  INV_X1 u2_u15_u5_U31 (.A( u2_u15_u5_n139 ) , .ZN( u2_u15_u5_n189 ) );
  INV_X1 u2_u15_u5_U32 (.A( u2_u15_u5_n157 ) , .ZN( u2_u15_u5_n190 ) );
  INV_X1 u2_u15_u5_U33 (.A( u2_u15_u5_n120 ) , .ZN( u2_u15_u5_n193 ) );
  NAND2_X1 u2_u15_u5_U34 (.ZN( u2_u15_u5_n111 ) , .A1( u2_u15_u5_n140 ) , .A2( u2_u15_u5_n155 ) );
  NOR2_X1 u2_u15_u5_U35 (.ZN( u2_u15_u5_n100 ) , .A1( u2_u15_u5_n170 ) , .A2( u2_u15_u5_n180 ) );
  INV_X1 u2_u15_u5_U36 (.A( u2_u15_u5_n117 ) , .ZN( u2_u15_u5_n196 ) );
  OAI221_X1 u2_u15_u5_U37 (.A( u2_u15_u5_n116 ) , .ZN( u2_u15_u5_n117 ) , .B2( u2_u15_u5_n119 ) , .C1( u2_u15_u5_n153 ) , .C2( u2_u15_u5_n158 ) , .B1( u2_u15_u5_n172 ) );
  AOI222_X1 u2_u15_u5_U38 (.ZN( u2_u15_u5_n116 ) , .B2( u2_u15_u5_n145 ) , .C1( u2_u15_u5_n148 ) , .A2( u2_u15_u5_n174 ) , .C2( u2_u15_u5_n177 ) , .B1( u2_u15_u5_n187 ) , .A1( u2_u15_u5_n193 ) );
  INV_X1 u2_u15_u5_U39 (.A( u2_u15_u5_n115 ) , .ZN( u2_u15_u5_n187 ) );
  INV_X1 u2_u15_u5_U4 (.A( u2_u15_u5_n138 ) , .ZN( u2_u15_u5_n191 ) );
  AOI22_X1 u2_u15_u5_U40 (.B2( u2_u15_u5_n131 ) , .A2( u2_u15_u5_n146 ) , .ZN( u2_u15_u5_n169 ) , .B1( u2_u15_u5_n174 ) , .A1( u2_u15_u5_n185 ) );
  NOR2_X1 u2_u15_u5_U41 (.A1( u2_u15_u5_n146 ) , .ZN( u2_u15_u5_n150 ) , .A2( u2_u15_u5_n173 ) );
  AOI21_X1 u2_u15_u5_U42 (.A( u2_u15_u5_n118 ) , .B2( u2_u15_u5_n145 ) , .ZN( u2_u15_u5_n168 ) , .B1( u2_u15_u5_n186 ) );
  INV_X1 u2_u15_u5_U43 (.A( u2_u15_u5_n122 ) , .ZN( u2_u15_u5_n186 ) );
  NOR2_X1 u2_u15_u5_U44 (.A1( u2_u15_u5_n146 ) , .ZN( u2_u15_u5_n152 ) , .A2( u2_u15_u5_n176 ) );
  NOR2_X1 u2_u15_u5_U45 (.A1( u2_u15_u5_n115 ) , .ZN( u2_u15_u5_n118 ) , .A2( u2_u15_u5_n153 ) );
  NOR2_X1 u2_u15_u5_U46 (.A2( u2_u15_u5_n145 ) , .ZN( u2_u15_u5_n156 ) , .A1( u2_u15_u5_n174 ) );
  NOR2_X1 u2_u15_u5_U47 (.ZN( u2_u15_u5_n121 ) , .A2( u2_u15_u5_n145 ) , .A1( u2_u15_u5_n176 ) );
  AOI22_X1 u2_u15_u5_U48 (.ZN( u2_u15_u5_n114 ) , .A2( u2_u15_u5_n137 ) , .A1( u2_u15_u5_n145 ) , .B2( u2_u15_u5_n175 ) , .B1( u2_u15_u5_n193 ) );
  OAI211_X1 u2_u15_u5_U49 (.B( u2_u15_u5_n124 ) , .A( u2_u15_u5_n125 ) , .C2( u2_u15_u5_n126 ) , .C1( u2_u15_u5_n127 ) , .ZN( u2_u15_u5_n128 ) );
  OAI21_X1 u2_u15_u5_U5 (.B2( u2_u15_u5_n136 ) , .B1( u2_u15_u5_n137 ) , .ZN( u2_u15_u5_n138 ) , .A( u2_u15_u5_n177 ) );
  NOR3_X1 u2_u15_u5_U50 (.ZN( u2_u15_u5_n127 ) , .A1( u2_u15_u5_n136 ) , .A3( u2_u15_u5_n148 ) , .A2( u2_u15_u5_n182 ) );
  OAI21_X1 u2_u15_u5_U51 (.ZN( u2_u15_u5_n124 ) , .A( u2_u15_u5_n177 ) , .B2( u2_u15_u5_n183 ) , .B1( u2_u15_u5_n189 ) );
  OAI21_X1 u2_u15_u5_U52 (.ZN( u2_u15_u5_n125 ) , .A( u2_u15_u5_n174 ) , .B2( u2_u15_u5_n185 ) , .B1( u2_u15_u5_n190 ) );
  AOI21_X1 u2_u15_u5_U53 (.A( u2_u15_u5_n153 ) , .B2( u2_u15_u5_n154 ) , .B1( u2_u15_u5_n155 ) , .ZN( u2_u15_u5_n164 ) );
  AOI21_X1 u2_u15_u5_U54 (.ZN( u2_u15_u5_n110 ) , .B1( u2_u15_u5_n122 ) , .B2( u2_u15_u5_n139 ) , .A( u2_u15_u5_n153 ) );
  INV_X1 u2_u15_u5_U55 (.A( u2_u15_u5_n153 ) , .ZN( u2_u15_u5_n176 ) );
  INV_X1 u2_u15_u5_U56 (.A( u2_u15_u5_n126 ) , .ZN( u2_u15_u5_n173 ) );
  AND2_X1 u2_u15_u5_U57 (.A2( u2_u15_u5_n104 ) , .A1( u2_u15_u5_n107 ) , .ZN( u2_u15_u5_n147 ) );
  AND2_X1 u2_u15_u5_U58 (.A2( u2_u15_u5_n104 ) , .A1( u2_u15_u5_n108 ) , .ZN( u2_u15_u5_n148 ) );
  NAND2_X1 u2_u15_u5_U59 (.A1( u2_u15_u5_n105 ) , .A2( u2_u15_u5_n106 ) , .ZN( u2_u15_u5_n158 ) );
  INV_X1 u2_u15_u5_U6 (.A( u2_u15_u5_n135 ) , .ZN( u2_u15_u5_n178 ) );
  NAND2_X1 u2_u15_u5_U60 (.A2( u2_u15_u5_n108 ) , .A1( u2_u15_u5_n109 ) , .ZN( u2_u15_u5_n139 ) );
  NAND2_X1 u2_u15_u5_U61 (.A1( u2_u15_u5_n106 ) , .A2( u2_u15_u5_n108 ) , .ZN( u2_u15_u5_n119 ) );
  NAND2_X1 u2_u15_u5_U62 (.A2( u2_u15_u5_n103 ) , .A1( u2_u15_u5_n105 ) , .ZN( u2_u15_u5_n140 ) );
  NAND2_X1 u2_u15_u5_U63 (.A2( u2_u15_u5_n104 ) , .A1( u2_u15_u5_n105 ) , .ZN( u2_u15_u5_n155 ) );
  NAND2_X1 u2_u15_u5_U64 (.A2( u2_u15_u5_n106 ) , .A1( u2_u15_u5_n107 ) , .ZN( u2_u15_u5_n122 ) );
  NAND2_X1 u2_u15_u5_U65 (.A2( u2_u15_u5_n100 ) , .A1( u2_u15_u5_n106 ) , .ZN( u2_u15_u5_n115 ) );
  NAND2_X1 u2_u15_u5_U66 (.A2( u2_u15_u5_n100 ) , .A1( u2_u15_u5_n103 ) , .ZN( u2_u15_u5_n161 ) );
  NAND2_X1 u2_u15_u5_U67 (.A1( u2_u15_u5_n105 ) , .A2( u2_u15_u5_n109 ) , .ZN( u2_u15_u5_n154 ) );
  INV_X1 u2_u15_u5_U68 (.A( u2_u15_u5_n146 ) , .ZN( u2_u15_u5_n172 ) );
  NAND2_X1 u2_u15_u5_U69 (.A1( u2_u15_u5_n103 ) , .A2( u2_u15_u5_n108 ) , .ZN( u2_u15_u5_n123 ) );
  OAI22_X1 u2_u15_u5_U7 (.B2( u2_u15_u5_n149 ) , .B1( u2_u15_u5_n150 ) , .A2( u2_u15_u5_n151 ) , .A1( u2_u15_u5_n152 ) , .ZN( u2_u15_u5_n165 ) );
  NAND2_X1 u2_u15_u5_U70 (.A2( u2_u15_u5_n103 ) , .A1( u2_u15_u5_n107 ) , .ZN( u2_u15_u5_n151 ) );
  NAND2_X1 u2_u15_u5_U71 (.A2( u2_u15_u5_n107 ) , .A1( u2_u15_u5_n109 ) , .ZN( u2_u15_u5_n120 ) );
  NAND2_X1 u2_u15_u5_U72 (.A2( u2_u15_u5_n100 ) , .A1( u2_u15_u5_n109 ) , .ZN( u2_u15_u5_n157 ) );
  AND2_X1 u2_u15_u5_U73 (.A2( u2_u15_u5_n100 ) , .A1( u2_u15_u5_n104 ) , .ZN( u2_u15_u5_n131 ) );
  INV_X1 u2_u15_u5_U74 (.A( u2_u15_u5_n102 ) , .ZN( u2_u15_u5_n195 ) );
  OAI221_X1 u2_u15_u5_U75 (.A( u2_u15_u5_n101 ) , .ZN( u2_u15_u5_n102 ) , .C2( u2_u15_u5_n115 ) , .C1( u2_u15_u5_n126 ) , .B1( u2_u15_u5_n134 ) , .B2( u2_u15_u5_n160 ) );
  OAI21_X1 u2_u15_u5_U76 (.ZN( u2_u15_u5_n101 ) , .B1( u2_u15_u5_n137 ) , .A( u2_u15_u5_n146 ) , .B2( u2_u15_u5_n147 ) );
  NOR2_X1 u2_u15_u5_U77 (.A2( u2_u15_X_34 ) , .A1( u2_u15_X_35 ) , .ZN( u2_u15_u5_n145 ) );
  NOR2_X1 u2_u15_u5_U78 (.A2( u2_u15_X_34 ) , .ZN( u2_u15_u5_n146 ) , .A1( u2_u15_u5_n171 ) );
  NOR2_X1 u2_u15_u5_U79 (.A2( u2_u15_X_31 ) , .A1( u2_u15_X_32 ) , .ZN( u2_u15_u5_n103 ) );
  NOR3_X1 u2_u15_u5_U8 (.A2( u2_u15_u5_n147 ) , .A1( u2_u15_u5_n148 ) , .ZN( u2_u15_u5_n149 ) , .A3( u2_u15_u5_n194 ) );
  NOR2_X1 u2_u15_u5_U80 (.A2( u2_u15_X_36 ) , .ZN( u2_u15_u5_n105 ) , .A1( u2_u15_u5_n180 ) );
  NOR2_X1 u2_u15_u5_U81 (.A2( u2_u15_X_33 ) , .ZN( u2_u15_u5_n108 ) , .A1( u2_u15_u5_n170 ) );
  NOR2_X1 u2_u15_u5_U82 (.A2( u2_u15_X_33 ) , .A1( u2_u15_X_36 ) , .ZN( u2_u15_u5_n107 ) );
  NOR2_X1 u2_u15_u5_U83 (.A2( u2_u15_X_31 ) , .ZN( u2_u15_u5_n104 ) , .A1( u2_u15_u5_n181 ) );
  NAND2_X1 u2_u15_u5_U84 (.A2( u2_u15_X_34 ) , .A1( u2_u15_X_35 ) , .ZN( u2_u15_u5_n153 ) );
  NAND2_X1 u2_u15_u5_U85 (.A1( u2_u15_X_34 ) , .ZN( u2_u15_u5_n126 ) , .A2( u2_u15_u5_n171 ) );
  AND2_X1 u2_u15_u5_U86 (.A1( u2_u15_X_31 ) , .A2( u2_u15_X_32 ) , .ZN( u2_u15_u5_n106 ) );
  AND2_X1 u2_u15_u5_U87 (.A1( u2_u15_X_31 ) , .ZN( u2_u15_u5_n109 ) , .A2( u2_u15_u5_n181 ) );
  INV_X1 u2_u15_u5_U88 (.A( u2_u15_X_33 ) , .ZN( u2_u15_u5_n180 ) );
  INV_X1 u2_u15_u5_U89 (.A( u2_u15_X_35 ) , .ZN( u2_u15_u5_n171 ) );
  NOR2_X1 u2_u15_u5_U9 (.ZN( u2_u15_u5_n135 ) , .A1( u2_u15_u5_n173 ) , .A2( u2_u15_u5_n176 ) );
  INV_X1 u2_u15_u5_U90 (.A( u2_u15_X_36 ) , .ZN( u2_u15_u5_n170 ) );
  INV_X1 u2_u15_u5_U91 (.A( u2_u15_X_32 ) , .ZN( u2_u15_u5_n181 ) );
  NAND4_X1 u2_u15_u5_U92 (.ZN( u2_out15_19 ) , .A4( u2_u15_u5_n166 ) , .A3( u2_u15_u5_n167 ) , .A2( u2_u15_u5_n168 ) , .A1( u2_u15_u5_n169 ) );
  AOI22_X1 u2_u15_u5_U93 (.B2( u2_u15_u5_n145 ) , .A2( u2_u15_u5_n146 ) , .ZN( u2_u15_u5_n167 ) , .B1( u2_u15_u5_n182 ) , .A1( u2_u15_u5_n189 ) );
  NOR4_X1 u2_u15_u5_U94 (.A4( u2_u15_u5_n162 ) , .A3( u2_u15_u5_n163 ) , .A2( u2_u15_u5_n164 ) , .A1( u2_u15_u5_n165 ) , .ZN( u2_u15_u5_n166 ) );
  NAND4_X1 u2_u15_u5_U95 (.ZN( u2_out15_11 ) , .A4( u2_u15_u5_n143 ) , .A3( u2_u15_u5_n144 ) , .A2( u2_u15_u5_n169 ) , .A1( u2_u15_u5_n196 ) );
  AOI22_X1 u2_u15_u5_U96 (.A2( u2_u15_u5_n132 ) , .ZN( u2_u15_u5_n144 ) , .B2( u2_u15_u5_n145 ) , .B1( u2_u15_u5_n184 ) , .A1( u2_u15_u5_n194 ) );
  NOR3_X1 u2_u15_u5_U97 (.A3( u2_u15_u5_n141 ) , .A1( u2_u15_u5_n142 ) , .ZN( u2_u15_u5_n143 ) , .A2( u2_u15_u5_n191 ) );
  NAND4_X1 u2_u15_u5_U98 (.ZN( u2_out15_4 ) , .A4( u2_u15_u5_n112 ) , .A2( u2_u15_u5_n113 ) , .A1( u2_u15_u5_n114 ) , .A3( u2_u15_u5_n195 ) );
  AOI211_X1 u2_u15_u5_U99 (.A( u2_u15_u5_n110 ) , .C1( u2_u15_u5_n111 ) , .ZN( u2_u15_u5_n112 ) , .B( u2_u15_u5_n118 ) , .C2( u2_u15_u5_n177 ) );
  INV_X1 u2_u15_u6_U10 (.ZN( u2_u15_u6_n172 ) , .A( u2_u15_u6_n88 ) );
  OAI21_X1 u2_u15_u6_U11 (.A( u2_u15_u6_n159 ) , .B1( u2_u15_u6_n169 ) , .B2( u2_u15_u6_n173 ) , .ZN( u2_u15_u6_n90 ) );
  AOI22_X1 u2_u15_u6_U12 (.A2( u2_u15_u6_n151 ) , .B2( u2_u15_u6_n161 ) , .A1( u2_u15_u6_n167 ) , .B1( u2_u15_u6_n170 ) , .ZN( u2_u15_u6_n89 ) );
  AOI21_X1 u2_u15_u6_U13 (.ZN( u2_u15_u6_n106 ) , .A( u2_u15_u6_n142 ) , .B2( u2_u15_u6_n159 ) , .B1( u2_u15_u6_n164 ) );
  INV_X1 u2_u15_u6_U14 (.A( u2_u15_u6_n155 ) , .ZN( u2_u15_u6_n161 ) );
  INV_X1 u2_u15_u6_U15 (.A( u2_u15_u6_n128 ) , .ZN( u2_u15_u6_n164 ) );
  NAND2_X1 u2_u15_u6_U16 (.ZN( u2_u15_u6_n110 ) , .A1( u2_u15_u6_n122 ) , .A2( u2_u15_u6_n129 ) );
  NAND2_X1 u2_u15_u6_U17 (.ZN( u2_u15_u6_n124 ) , .A2( u2_u15_u6_n146 ) , .A1( u2_u15_u6_n148 ) );
  INV_X1 u2_u15_u6_U18 (.A( u2_u15_u6_n132 ) , .ZN( u2_u15_u6_n171 ) );
  AND2_X1 u2_u15_u6_U19 (.A1( u2_u15_u6_n100 ) , .ZN( u2_u15_u6_n130 ) , .A2( u2_u15_u6_n147 ) );
  INV_X1 u2_u15_u6_U20 (.A( u2_u15_u6_n127 ) , .ZN( u2_u15_u6_n173 ) );
  INV_X1 u2_u15_u6_U21 (.A( u2_u15_u6_n121 ) , .ZN( u2_u15_u6_n167 ) );
  INV_X1 u2_u15_u6_U22 (.A( u2_u15_u6_n100 ) , .ZN( u2_u15_u6_n169 ) );
  INV_X1 u2_u15_u6_U23 (.A( u2_u15_u6_n123 ) , .ZN( u2_u15_u6_n170 ) );
  INV_X1 u2_u15_u6_U24 (.A( u2_u15_u6_n113 ) , .ZN( u2_u15_u6_n168 ) );
  AND2_X1 u2_u15_u6_U25 (.A1( u2_u15_u6_n107 ) , .A2( u2_u15_u6_n119 ) , .ZN( u2_u15_u6_n133 ) );
  AND2_X1 u2_u15_u6_U26 (.A2( u2_u15_u6_n121 ) , .A1( u2_u15_u6_n122 ) , .ZN( u2_u15_u6_n131 ) );
  AND3_X1 u2_u15_u6_U27 (.ZN( u2_u15_u6_n120 ) , .A2( u2_u15_u6_n127 ) , .A1( u2_u15_u6_n132 ) , .A3( u2_u15_u6_n145 ) );
  INV_X1 u2_u15_u6_U28 (.A( u2_u15_u6_n146 ) , .ZN( u2_u15_u6_n163 ) );
  AOI222_X1 u2_u15_u6_U29 (.ZN( u2_u15_u6_n114 ) , .A1( u2_u15_u6_n118 ) , .A2( u2_u15_u6_n126 ) , .B2( u2_u15_u6_n151 ) , .C2( u2_u15_u6_n159 ) , .C1( u2_u15_u6_n168 ) , .B1( u2_u15_u6_n169 ) );
  INV_X1 u2_u15_u6_U3 (.A( u2_u15_u6_n110 ) , .ZN( u2_u15_u6_n166 ) );
  NOR2_X1 u2_u15_u6_U30 (.A1( u2_u15_u6_n162 ) , .A2( u2_u15_u6_n165 ) , .ZN( u2_u15_u6_n98 ) );
  NAND2_X1 u2_u15_u6_U31 (.A1( u2_u15_u6_n144 ) , .ZN( u2_u15_u6_n151 ) , .A2( u2_u15_u6_n158 ) );
  NAND2_X1 u2_u15_u6_U32 (.ZN( u2_u15_u6_n132 ) , .A1( u2_u15_u6_n91 ) , .A2( u2_u15_u6_n97 ) );
  AOI22_X1 u2_u15_u6_U33 (.B2( u2_u15_u6_n110 ) , .B1( u2_u15_u6_n111 ) , .A1( u2_u15_u6_n112 ) , .ZN( u2_u15_u6_n115 ) , .A2( u2_u15_u6_n161 ) );
  NAND4_X1 u2_u15_u6_U34 (.A3( u2_u15_u6_n109 ) , .ZN( u2_u15_u6_n112 ) , .A4( u2_u15_u6_n132 ) , .A2( u2_u15_u6_n147 ) , .A1( u2_u15_u6_n166 ) );
  NOR2_X1 u2_u15_u6_U35 (.ZN( u2_u15_u6_n109 ) , .A1( u2_u15_u6_n170 ) , .A2( u2_u15_u6_n173 ) );
  NOR2_X1 u2_u15_u6_U36 (.A2( u2_u15_u6_n126 ) , .ZN( u2_u15_u6_n155 ) , .A1( u2_u15_u6_n160 ) );
  NAND2_X1 u2_u15_u6_U37 (.ZN( u2_u15_u6_n146 ) , .A2( u2_u15_u6_n94 ) , .A1( u2_u15_u6_n99 ) );
  AOI21_X1 u2_u15_u6_U38 (.A( u2_u15_u6_n144 ) , .B2( u2_u15_u6_n145 ) , .B1( u2_u15_u6_n146 ) , .ZN( u2_u15_u6_n150 ) );
  AOI211_X1 u2_u15_u6_U39 (.B( u2_u15_u6_n134 ) , .A( u2_u15_u6_n135 ) , .C1( u2_u15_u6_n136 ) , .ZN( u2_u15_u6_n137 ) , .C2( u2_u15_u6_n151 ) );
  INV_X1 u2_u15_u6_U4 (.A( u2_u15_u6_n142 ) , .ZN( u2_u15_u6_n174 ) );
  NAND4_X1 u2_u15_u6_U40 (.A4( u2_u15_u6_n127 ) , .A3( u2_u15_u6_n128 ) , .A2( u2_u15_u6_n129 ) , .A1( u2_u15_u6_n130 ) , .ZN( u2_u15_u6_n136 ) );
  AOI21_X1 u2_u15_u6_U41 (.B2( u2_u15_u6_n132 ) , .B1( u2_u15_u6_n133 ) , .ZN( u2_u15_u6_n134 ) , .A( u2_u15_u6_n158 ) );
  AOI21_X1 u2_u15_u6_U42 (.B1( u2_u15_u6_n131 ) , .ZN( u2_u15_u6_n135 ) , .A( u2_u15_u6_n144 ) , .B2( u2_u15_u6_n146 ) );
  INV_X1 u2_u15_u6_U43 (.A( u2_u15_u6_n111 ) , .ZN( u2_u15_u6_n158 ) );
  NAND2_X1 u2_u15_u6_U44 (.ZN( u2_u15_u6_n127 ) , .A1( u2_u15_u6_n91 ) , .A2( u2_u15_u6_n92 ) );
  NAND2_X1 u2_u15_u6_U45 (.ZN( u2_u15_u6_n129 ) , .A2( u2_u15_u6_n95 ) , .A1( u2_u15_u6_n96 ) );
  INV_X1 u2_u15_u6_U46 (.A( u2_u15_u6_n144 ) , .ZN( u2_u15_u6_n159 ) );
  NAND2_X1 u2_u15_u6_U47 (.ZN( u2_u15_u6_n145 ) , .A2( u2_u15_u6_n97 ) , .A1( u2_u15_u6_n98 ) );
  NAND2_X1 u2_u15_u6_U48 (.ZN( u2_u15_u6_n148 ) , .A2( u2_u15_u6_n92 ) , .A1( u2_u15_u6_n94 ) );
  NAND2_X1 u2_u15_u6_U49 (.ZN( u2_u15_u6_n108 ) , .A2( u2_u15_u6_n139 ) , .A1( u2_u15_u6_n144 ) );
  NAND2_X1 u2_u15_u6_U5 (.A2( u2_u15_u6_n143 ) , .ZN( u2_u15_u6_n152 ) , .A1( u2_u15_u6_n166 ) );
  NAND2_X1 u2_u15_u6_U50 (.ZN( u2_u15_u6_n121 ) , .A2( u2_u15_u6_n95 ) , .A1( u2_u15_u6_n97 ) );
  NAND2_X1 u2_u15_u6_U51 (.ZN( u2_u15_u6_n107 ) , .A2( u2_u15_u6_n92 ) , .A1( u2_u15_u6_n95 ) );
  AND2_X1 u2_u15_u6_U52 (.ZN( u2_u15_u6_n118 ) , .A2( u2_u15_u6_n91 ) , .A1( u2_u15_u6_n99 ) );
  NAND2_X1 u2_u15_u6_U53 (.ZN( u2_u15_u6_n147 ) , .A2( u2_u15_u6_n98 ) , .A1( u2_u15_u6_n99 ) );
  NAND2_X1 u2_u15_u6_U54 (.ZN( u2_u15_u6_n128 ) , .A1( u2_u15_u6_n94 ) , .A2( u2_u15_u6_n96 ) );
  NAND2_X1 u2_u15_u6_U55 (.ZN( u2_u15_u6_n119 ) , .A2( u2_u15_u6_n95 ) , .A1( u2_u15_u6_n99 ) );
  NAND2_X1 u2_u15_u6_U56 (.ZN( u2_u15_u6_n123 ) , .A2( u2_u15_u6_n91 ) , .A1( u2_u15_u6_n96 ) );
  NAND2_X1 u2_u15_u6_U57 (.ZN( u2_u15_u6_n100 ) , .A2( u2_u15_u6_n92 ) , .A1( u2_u15_u6_n98 ) );
  NAND2_X1 u2_u15_u6_U58 (.ZN( u2_u15_u6_n122 ) , .A1( u2_u15_u6_n94 ) , .A2( u2_u15_u6_n97 ) );
  INV_X1 u2_u15_u6_U59 (.A( u2_u15_u6_n139 ) , .ZN( u2_u15_u6_n160 ) );
  AOI22_X1 u2_u15_u6_U6 (.B2( u2_u15_u6_n101 ) , .A1( u2_u15_u6_n102 ) , .ZN( u2_u15_u6_n103 ) , .B1( u2_u15_u6_n160 ) , .A2( u2_u15_u6_n161 ) );
  NAND2_X1 u2_u15_u6_U60 (.ZN( u2_u15_u6_n113 ) , .A1( u2_u15_u6_n96 ) , .A2( u2_u15_u6_n98 ) );
  NOR2_X1 u2_u15_u6_U61 (.A2( u2_u15_X_40 ) , .A1( u2_u15_X_41 ) , .ZN( u2_u15_u6_n126 ) );
  NOR2_X1 u2_u15_u6_U62 (.A2( u2_u15_X_39 ) , .A1( u2_u15_X_42 ) , .ZN( u2_u15_u6_n92 ) );
  NOR2_X1 u2_u15_u6_U63 (.A2( u2_u15_X_39 ) , .A1( u2_u15_u6_n156 ) , .ZN( u2_u15_u6_n97 ) );
  NOR2_X1 u2_u15_u6_U64 (.A2( u2_u15_X_38 ) , .A1( u2_u15_u6_n165 ) , .ZN( u2_u15_u6_n95 ) );
  NOR2_X1 u2_u15_u6_U65 (.A2( u2_u15_X_41 ) , .ZN( u2_u15_u6_n111 ) , .A1( u2_u15_u6_n157 ) );
  NOR2_X1 u2_u15_u6_U66 (.A2( u2_u15_X_37 ) , .A1( u2_u15_u6_n162 ) , .ZN( u2_u15_u6_n94 ) );
  NOR2_X1 u2_u15_u6_U67 (.A2( u2_u15_X_37 ) , .A1( u2_u15_X_38 ) , .ZN( u2_u15_u6_n91 ) );
  NAND2_X1 u2_u15_u6_U68 (.A1( u2_u15_X_41 ) , .ZN( u2_u15_u6_n144 ) , .A2( u2_u15_u6_n157 ) );
  NAND2_X1 u2_u15_u6_U69 (.A2( u2_u15_X_40 ) , .A1( u2_u15_X_41 ) , .ZN( u2_u15_u6_n139 ) );
  NOR2_X1 u2_u15_u6_U7 (.A1( u2_u15_u6_n118 ) , .ZN( u2_u15_u6_n143 ) , .A2( u2_u15_u6_n168 ) );
  AND2_X1 u2_u15_u6_U70 (.A1( u2_u15_X_39 ) , .A2( u2_u15_u6_n156 ) , .ZN( u2_u15_u6_n96 ) );
  AND2_X1 u2_u15_u6_U71 (.A1( u2_u15_X_39 ) , .A2( u2_u15_X_42 ) , .ZN( u2_u15_u6_n99 ) );
  INV_X1 u2_u15_u6_U72 (.A( u2_u15_X_40 ) , .ZN( u2_u15_u6_n157 ) );
  INV_X1 u2_u15_u6_U73 (.A( u2_u15_X_37 ) , .ZN( u2_u15_u6_n165 ) );
  INV_X1 u2_u15_u6_U74 (.A( u2_u15_X_38 ) , .ZN( u2_u15_u6_n162 ) );
  INV_X1 u2_u15_u6_U75 (.A( u2_u15_X_42 ) , .ZN( u2_u15_u6_n156 ) );
  NAND4_X1 u2_u15_u6_U76 (.ZN( u2_out15_12 ) , .A4( u2_u15_u6_n114 ) , .A3( u2_u15_u6_n115 ) , .A2( u2_u15_u6_n116 ) , .A1( u2_u15_u6_n117 ) );
  OAI22_X1 u2_u15_u6_U77 (.B2( u2_u15_u6_n111 ) , .ZN( u2_u15_u6_n116 ) , .B1( u2_u15_u6_n126 ) , .A2( u2_u15_u6_n164 ) , .A1( u2_u15_u6_n167 ) );
  OAI21_X1 u2_u15_u6_U78 (.A( u2_u15_u6_n108 ) , .ZN( u2_u15_u6_n117 ) , .B2( u2_u15_u6_n141 ) , .B1( u2_u15_u6_n163 ) );
  NAND4_X1 u2_u15_u6_U79 (.ZN( u2_out15_32 ) , .A4( u2_u15_u6_n103 ) , .A3( u2_u15_u6_n104 ) , .A2( u2_u15_u6_n105 ) , .A1( u2_u15_u6_n106 ) );
  AOI21_X1 u2_u15_u6_U8 (.B1( u2_u15_u6_n107 ) , .B2( u2_u15_u6_n132 ) , .A( u2_u15_u6_n158 ) , .ZN( u2_u15_u6_n88 ) );
  AOI22_X1 u2_u15_u6_U80 (.ZN( u2_u15_u6_n105 ) , .A2( u2_u15_u6_n108 ) , .A1( u2_u15_u6_n118 ) , .B2( u2_u15_u6_n126 ) , .B1( u2_u15_u6_n171 ) );
  AOI22_X1 u2_u15_u6_U81 (.ZN( u2_u15_u6_n104 ) , .A1( u2_u15_u6_n111 ) , .B1( u2_u15_u6_n124 ) , .B2( u2_u15_u6_n151 ) , .A2( u2_u15_u6_n93 ) );
  OAI211_X1 u2_u15_u6_U82 (.ZN( u2_out15_22 ) , .B( u2_u15_u6_n137 ) , .A( u2_u15_u6_n138 ) , .C2( u2_u15_u6_n139 ) , .C1( u2_u15_u6_n140 ) );
  AOI22_X1 u2_u15_u6_U83 (.B1( u2_u15_u6_n124 ) , .A2( u2_u15_u6_n125 ) , .A1( u2_u15_u6_n126 ) , .ZN( u2_u15_u6_n138 ) , .B2( u2_u15_u6_n161 ) );
  AND4_X1 u2_u15_u6_U84 (.A3( u2_u15_u6_n119 ) , .A1( u2_u15_u6_n120 ) , .A4( u2_u15_u6_n129 ) , .ZN( u2_u15_u6_n140 ) , .A2( u2_u15_u6_n143 ) );
  OAI211_X1 u2_u15_u6_U85 (.ZN( u2_out15_7 ) , .B( u2_u15_u6_n153 ) , .C2( u2_u15_u6_n154 ) , .C1( u2_u15_u6_n155 ) , .A( u2_u15_u6_n174 ) );
  NOR3_X1 u2_u15_u6_U86 (.A1( u2_u15_u6_n141 ) , .ZN( u2_u15_u6_n154 ) , .A3( u2_u15_u6_n164 ) , .A2( u2_u15_u6_n171 ) );
  AOI211_X1 u2_u15_u6_U87 (.B( u2_u15_u6_n149 ) , .A( u2_u15_u6_n150 ) , .C2( u2_u15_u6_n151 ) , .C1( u2_u15_u6_n152 ) , .ZN( u2_u15_u6_n153 ) );
  NAND3_X1 u2_u15_u6_U88 (.A2( u2_u15_u6_n123 ) , .ZN( u2_u15_u6_n125 ) , .A1( u2_u15_u6_n130 ) , .A3( u2_u15_u6_n131 ) );
  NAND3_X1 u2_u15_u6_U89 (.A3( u2_u15_u6_n133 ) , .ZN( u2_u15_u6_n141 ) , .A1( u2_u15_u6_n145 ) , .A2( u2_u15_u6_n148 ) );
  AOI21_X1 u2_u15_u6_U9 (.B2( u2_u15_u6_n147 ) , .B1( u2_u15_u6_n148 ) , .ZN( u2_u15_u6_n149 ) , .A( u2_u15_u6_n158 ) );
  NAND3_X1 u2_u15_u6_U90 (.ZN( u2_u15_u6_n101 ) , .A3( u2_u15_u6_n107 ) , .A2( u2_u15_u6_n121 ) , .A1( u2_u15_u6_n127 ) );
  NAND3_X1 u2_u15_u6_U91 (.ZN( u2_u15_u6_n102 ) , .A3( u2_u15_u6_n130 ) , .A2( u2_u15_u6_n145 ) , .A1( u2_u15_u6_n166 ) );
  NAND3_X1 u2_u15_u6_U92 (.A3( u2_u15_u6_n113 ) , .A1( u2_u15_u6_n119 ) , .A2( u2_u15_u6_n123 ) , .ZN( u2_u15_u6_n93 ) );
  NAND3_X1 u2_u15_u6_U93 (.ZN( u2_u15_u6_n142 ) , .A2( u2_u15_u6_n172 ) , .A3( u2_u15_u6_n89 ) , .A1( u2_u15_u6_n90 ) );
  OAI21_X1 u2_u15_u7_U10 (.A( u2_u15_u7_n161 ) , .B1( u2_u15_u7_n168 ) , .B2( u2_u15_u7_n173 ) , .ZN( u2_u15_u7_n91 ) );
  AOI211_X1 u2_u15_u7_U11 (.A( u2_u15_u7_n117 ) , .ZN( u2_u15_u7_n118 ) , .C2( u2_u15_u7_n126 ) , .C1( u2_u15_u7_n177 ) , .B( u2_u15_u7_n180 ) );
  OAI22_X1 u2_u15_u7_U12 (.B1( u2_u15_u7_n115 ) , .ZN( u2_u15_u7_n117 ) , .A2( u2_u15_u7_n133 ) , .A1( u2_u15_u7_n137 ) , .B2( u2_u15_u7_n162 ) );
  INV_X1 u2_u15_u7_U13 (.A( u2_u15_u7_n116 ) , .ZN( u2_u15_u7_n180 ) );
  NOR3_X1 u2_u15_u7_U14 (.ZN( u2_u15_u7_n115 ) , .A3( u2_u15_u7_n145 ) , .A2( u2_u15_u7_n168 ) , .A1( u2_u15_u7_n169 ) );
  OAI211_X1 u2_u15_u7_U15 (.B( u2_u15_u7_n122 ) , .A( u2_u15_u7_n123 ) , .C2( u2_u15_u7_n124 ) , .ZN( u2_u15_u7_n154 ) , .C1( u2_u15_u7_n162 ) );
  AOI222_X1 u2_u15_u7_U16 (.ZN( u2_u15_u7_n122 ) , .C2( u2_u15_u7_n126 ) , .C1( u2_u15_u7_n145 ) , .B1( u2_u15_u7_n161 ) , .A2( u2_u15_u7_n165 ) , .B2( u2_u15_u7_n170 ) , .A1( u2_u15_u7_n176 ) );
  INV_X1 u2_u15_u7_U17 (.A( u2_u15_u7_n133 ) , .ZN( u2_u15_u7_n176 ) );
  NOR3_X1 u2_u15_u7_U18 (.A2( u2_u15_u7_n134 ) , .A1( u2_u15_u7_n135 ) , .ZN( u2_u15_u7_n136 ) , .A3( u2_u15_u7_n171 ) );
  NOR2_X1 u2_u15_u7_U19 (.A1( u2_u15_u7_n130 ) , .A2( u2_u15_u7_n134 ) , .ZN( u2_u15_u7_n153 ) );
  INV_X1 u2_u15_u7_U20 (.A( u2_u15_u7_n101 ) , .ZN( u2_u15_u7_n165 ) );
  NOR2_X1 u2_u15_u7_U21 (.ZN( u2_u15_u7_n111 ) , .A2( u2_u15_u7_n134 ) , .A1( u2_u15_u7_n169 ) );
  AOI21_X1 u2_u15_u7_U22 (.ZN( u2_u15_u7_n104 ) , .B2( u2_u15_u7_n112 ) , .B1( u2_u15_u7_n127 ) , .A( u2_u15_u7_n164 ) );
  AOI21_X1 u2_u15_u7_U23 (.ZN( u2_u15_u7_n106 ) , .B1( u2_u15_u7_n133 ) , .B2( u2_u15_u7_n146 ) , .A( u2_u15_u7_n162 ) );
  AOI21_X1 u2_u15_u7_U24 (.A( u2_u15_u7_n101 ) , .ZN( u2_u15_u7_n107 ) , .B2( u2_u15_u7_n128 ) , .B1( u2_u15_u7_n175 ) );
  INV_X1 u2_u15_u7_U25 (.A( u2_u15_u7_n138 ) , .ZN( u2_u15_u7_n171 ) );
  INV_X1 u2_u15_u7_U26 (.A( u2_u15_u7_n131 ) , .ZN( u2_u15_u7_n177 ) );
  INV_X1 u2_u15_u7_U27 (.A( u2_u15_u7_n110 ) , .ZN( u2_u15_u7_n174 ) );
  NAND2_X1 u2_u15_u7_U28 (.A1( u2_u15_u7_n129 ) , .A2( u2_u15_u7_n132 ) , .ZN( u2_u15_u7_n149 ) );
  NAND2_X1 u2_u15_u7_U29 (.A1( u2_u15_u7_n113 ) , .A2( u2_u15_u7_n124 ) , .ZN( u2_u15_u7_n130 ) );
  INV_X1 u2_u15_u7_U3 (.A( u2_u15_u7_n111 ) , .ZN( u2_u15_u7_n170 ) );
  INV_X1 u2_u15_u7_U30 (.A( u2_u15_u7_n112 ) , .ZN( u2_u15_u7_n173 ) );
  INV_X1 u2_u15_u7_U31 (.A( u2_u15_u7_n128 ) , .ZN( u2_u15_u7_n168 ) );
  INV_X1 u2_u15_u7_U32 (.A( u2_u15_u7_n148 ) , .ZN( u2_u15_u7_n169 ) );
  INV_X1 u2_u15_u7_U33 (.A( u2_u15_u7_n127 ) , .ZN( u2_u15_u7_n179 ) );
  NOR2_X1 u2_u15_u7_U34 (.ZN( u2_u15_u7_n101 ) , .A2( u2_u15_u7_n150 ) , .A1( u2_u15_u7_n156 ) );
  AOI211_X1 u2_u15_u7_U35 (.B( u2_u15_u7_n154 ) , .A( u2_u15_u7_n155 ) , .C1( u2_u15_u7_n156 ) , .ZN( u2_u15_u7_n157 ) , .C2( u2_u15_u7_n172 ) );
  INV_X1 u2_u15_u7_U36 (.A( u2_u15_u7_n153 ) , .ZN( u2_u15_u7_n172 ) );
  AOI211_X1 u2_u15_u7_U37 (.B( u2_u15_u7_n139 ) , .A( u2_u15_u7_n140 ) , .C2( u2_u15_u7_n141 ) , .ZN( u2_u15_u7_n142 ) , .C1( u2_u15_u7_n156 ) );
  NAND4_X1 u2_u15_u7_U38 (.A3( u2_u15_u7_n127 ) , .A2( u2_u15_u7_n128 ) , .A1( u2_u15_u7_n129 ) , .ZN( u2_u15_u7_n141 ) , .A4( u2_u15_u7_n147 ) );
  AOI21_X1 u2_u15_u7_U39 (.A( u2_u15_u7_n137 ) , .B1( u2_u15_u7_n138 ) , .ZN( u2_u15_u7_n139 ) , .B2( u2_u15_u7_n146 ) );
  INV_X1 u2_u15_u7_U4 (.A( u2_u15_u7_n149 ) , .ZN( u2_u15_u7_n175 ) );
  OAI22_X1 u2_u15_u7_U40 (.B1( u2_u15_u7_n136 ) , .ZN( u2_u15_u7_n140 ) , .A1( u2_u15_u7_n153 ) , .B2( u2_u15_u7_n162 ) , .A2( u2_u15_u7_n164 ) );
  AOI21_X1 u2_u15_u7_U41 (.ZN( u2_u15_u7_n123 ) , .B1( u2_u15_u7_n165 ) , .B2( u2_u15_u7_n177 ) , .A( u2_u15_u7_n97 ) );
  AOI21_X1 u2_u15_u7_U42 (.B2( u2_u15_u7_n113 ) , .B1( u2_u15_u7_n124 ) , .A( u2_u15_u7_n125 ) , .ZN( u2_u15_u7_n97 ) );
  INV_X1 u2_u15_u7_U43 (.A( u2_u15_u7_n125 ) , .ZN( u2_u15_u7_n161 ) );
  INV_X1 u2_u15_u7_U44 (.A( u2_u15_u7_n152 ) , .ZN( u2_u15_u7_n162 ) );
  AOI22_X1 u2_u15_u7_U45 (.A2( u2_u15_u7_n114 ) , .ZN( u2_u15_u7_n119 ) , .B1( u2_u15_u7_n130 ) , .A1( u2_u15_u7_n156 ) , .B2( u2_u15_u7_n165 ) );
  NAND2_X1 u2_u15_u7_U46 (.A2( u2_u15_u7_n112 ) , .ZN( u2_u15_u7_n114 ) , .A1( u2_u15_u7_n175 ) );
  AOI22_X1 u2_u15_u7_U47 (.B2( u2_u15_u7_n149 ) , .B1( u2_u15_u7_n150 ) , .A2( u2_u15_u7_n151 ) , .A1( u2_u15_u7_n152 ) , .ZN( u2_u15_u7_n158 ) );
  AND2_X1 u2_u15_u7_U48 (.ZN( u2_u15_u7_n145 ) , .A2( u2_u15_u7_n98 ) , .A1( u2_u15_u7_n99 ) );
  NOR2_X1 u2_u15_u7_U49 (.ZN( u2_u15_u7_n137 ) , .A1( u2_u15_u7_n150 ) , .A2( u2_u15_u7_n161 ) );
  INV_X1 u2_u15_u7_U5 (.A( u2_u15_u7_n154 ) , .ZN( u2_u15_u7_n178 ) );
  AOI21_X1 u2_u15_u7_U50 (.ZN( u2_u15_u7_n105 ) , .B2( u2_u15_u7_n110 ) , .A( u2_u15_u7_n125 ) , .B1( u2_u15_u7_n147 ) );
  NAND2_X1 u2_u15_u7_U51 (.ZN( u2_u15_u7_n146 ) , .A1( u2_u15_u7_n95 ) , .A2( u2_u15_u7_n98 ) );
  NAND2_X1 u2_u15_u7_U52 (.A2( u2_u15_u7_n103 ) , .ZN( u2_u15_u7_n147 ) , .A1( u2_u15_u7_n93 ) );
  NAND2_X1 u2_u15_u7_U53 (.A1( u2_u15_u7_n103 ) , .ZN( u2_u15_u7_n127 ) , .A2( u2_u15_u7_n99 ) );
  OR2_X1 u2_u15_u7_U54 (.ZN( u2_u15_u7_n126 ) , .A2( u2_u15_u7_n152 ) , .A1( u2_u15_u7_n156 ) );
  NAND2_X1 u2_u15_u7_U55 (.A2( u2_u15_u7_n102 ) , .A1( u2_u15_u7_n103 ) , .ZN( u2_u15_u7_n133 ) );
  NAND2_X1 u2_u15_u7_U56 (.ZN( u2_u15_u7_n112 ) , .A2( u2_u15_u7_n96 ) , .A1( u2_u15_u7_n99 ) );
  NAND2_X1 u2_u15_u7_U57 (.A2( u2_u15_u7_n102 ) , .ZN( u2_u15_u7_n128 ) , .A1( u2_u15_u7_n98 ) );
  NAND2_X1 u2_u15_u7_U58 (.A1( u2_u15_u7_n100 ) , .ZN( u2_u15_u7_n113 ) , .A2( u2_u15_u7_n93 ) );
  NAND2_X1 u2_u15_u7_U59 (.A2( u2_u15_u7_n102 ) , .ZN( u2_u15_u7_n124 ) , .A1( u2_u15_u7_n96 ) );
  AOI211_X1 u2_u15_u7_U6 (.ZN( u2_u15_u7_n116 ) , .A( u2_u15_u7_n155 ) , .C1( u2_u15_u7_n161 ) , .C2( u2_u15_u7_n171 ) , .B( u2_u15_u7_n94 ) );
  NAND2_X1 u2_u15_u7_U60 (.ZN( u2_u15_u7_n110 ) , .A1( u2_u15_u7_n95 ) , .A2( u2_u15_u7_n96 ) );
  INV_X1 u2_u15_u7_U61 (.A( u2_u15_u7_n150 ) , .ZN( u2_u15_u7_n164 ) );
  AND2_X1 u2_u15_u7_U62 (.ZN( u2_u15_u7_n134 ) , .A1( u2_u15_u7_n93 ) , .A2( u2_u15_u7_n98 ) );
  NAND2_X1 u2_u15_u7_U63 (.A1( u2_u15_u7_n100 ) , .A2( u2_u15_u7_n102 ) , .ZN( u2_u15_u7_n129 ) );
  NAND2_X1 u2_u15_u7_U64 (.A2( u2_u15_u7_n103 ) , .ZN( u2_u15_u7_n131 ) , .A1( u2_u15_u7_n95 ) );
  NAND2_X1 u2_u15_u7_U65 (.A1( u2_u15_u7_n100 ) , .ZN( u2_u15_u7_n138 ) , .A2( u2_u15_u7_n99 ) );
  NAND2_X1 u2_u15_u7_U66 (.ZN( u2_u15_u7_n132 ) , .A1( u2_u15_u7_n93 ) , .A2( u2_u15_u7_n96 ) );
  NAND2_X1 u2_u15_u7_U67 (.A1( u2_u15_u7_n100 ) , .ZN( u2_u15_u7_n148 ) , .A2( u2_u15_u7_n95 ) );
  NOR2_X1 u2_u15_u7_U68 (.A2( u2_u15_X_47 ) , .ZN( u2_u15_u7_n150 ) , .A1( u2_u15_u7_n163 ) );
  NOR2_X1 u2_u15_u7_U69 (.A2( u2_u15_X_43 ) , .A1( u2_u15_X_44 ) , .ZN( u2_u15_u7_n103 ) );
  OAI222_X1 u2_u15_u7_U7 (.C2( u2_u15_u7_n101 ) , .B2( u2_u15_u7_n111 ) , .A1( u2_u15_u7_n113 ) , .C1( u2_u15_u7_n146 ) , .A2( u2_u15_u7_n162 ) , .B1( u2_u15_u7_n164 ) , .ZN( u2_u15_u7_n94 ) );
  NOR2_X1 u2_u15_u7_U70 (.A2( u2_u15_X_48 ) , .A1( u2_u15_u7_n166 ) , .ZN( u2_u15_u7_n95 ) );
  NOR2_X1 u2_u15_u7_U71 (.A2( u2_u15_X_45 ) , .A1( u2_u15_X_48 ) , .ZN( u2_u15_u7_n99 ) );
  NOR2_X1 u2_u15_u7_U72 (.A2( u2_u15_X_44 ) , .A1( u2_u15_u7_n167 ) , .ZN( u2_u15_u7_n98 ) );
  NOR2_X1 u2_u15_u7_U73 (.A2( u2_u15_X_46 ) , .A1( u2_u15_X_47 ) , .ZN( u2_u15_u7_n152 ) );
  AND2_X1 u2_u15_u7_U74 (.A1( u2_u15_X_47 ) , .ZN( u2_u15_u7_n156 ) , .A2( u2_u15_u7_n163 ) );
  NAND2_X1 u2_u15_u7_U75 (.A2( u2_u15_X_46 ) , .A1( u2_u15_X_47 ) , .ZN( u2_u15_u7_n125 ) );
  AND2_X1 u2_u15_u7_U76 (.A2( u2_u15_X_45 ) , .A1( u2_u15_X_48 ) , .ZN( u2_u15_u7_n102 ) );
  AND2_X1 u2_u15_u7_U77 (.A2( u2_u15_X_43 ) , .A1( u2_u15_X_44 ) , .ZN( u2_u15_u7_n96 ) );
  AND2_X1 u2_u15_u7_U78 (.A1( u2_u15_X_44 ) , .ZN( u2_u15_u7_n100 ) , .A2( u2_u15_u7_n167 ) );
  AND2_X1 u2_u15_u7_U79 (.A1( u2_u15_X_48 ) , .A2( u2_u15_u7_n166 ) , .ZN( u2_u15_u7_n93 ) );
  OAI221_X1 u2_u15_u7_U8 (.C1( u2_u15_u7_n101 ) , .C2( u2_u15_u7_n147 ) , .ZN( u2_u15_u7_n155 ) , .B2( u2_u15_u7_n162 ) , .A( u2_u15_u7_n91 ) , .B1( u2_u15_u7_n92 ) );
  INV_X1 u2_u15_u7_U80 (.A( u2_u15_X_46 ) , .ZN( u2_u15_u7_n163 ) );
  INV_X1 u2_u15_u7_U81 (.A( u2_u15_X_45 ) , .ZN( u2_u15_u7_n166 ) );
  INV_X1 u2_u15_u7_U82 (.A( u2_u15_X_43 ) , .ZN( u2_u15_u7_n167 ) );
  NAND4_X1 u2_u15_u7_U83 (.ZN( u2_out15_5 ) , .A4( u2_u15_u7_n108 ) , .A3( u2_u15_u7_n109 ) , .A1( u2_u15_u7_n116 ) , .A2( u2_u15_u7_n123 ) );
  AOI22_X1 u2_u15_u7_U84 (.ZN( u2_u15_u7_n109 ) , .A2( u2_u15_u7_n126 ) , .B2( u2_u15_u7_n145 ) , .B1( u2_u15_u7_n156 ) , .A1( u2_u15_u7_n171 ) );
  NOR4_X1 u2_u15_u7_U85 (.A4( u2_u15_u7_n104 ) , .A3( u2_u15_u7_n105 ) , .A2( u2_u15_u7_n106 ) , .A1( u2_u15_u7_n107 ) , .ZN( u2_u15_u7_n108 ) );
  NAND4_X1 u2_u15_u7_U86 (.ZN( u2_out15_27 ) , .A4( u2_u15_u7_n118 ) , .A3( u2_u15_u7_n119 ) , .A2( u2_u15_u7_n120 ) , .A1( u2_u15_u7_n121 ) );
  OAI21_X1 u2_u15_u7_U87 (.ZN( u2_u15_u7_n121 ) , .B2( u2_u15_u7_n145 ) , .A( u2_u15_u7_n150 ) , .B1( u2_u15_u7_n174 ) );
  OAI21_X1 u2_u15_u7_U88 (.ZN( u2_u15_u7_n120 ) , .A( u2_u15_u7_n161 ) , .B2( u2_u15_u7_n170 ) , .B1( u2_u15_u7_n179 ) );
  NAND4_X1 u2_u15_u7_U89 (.ZN( u2_out15_21 ) , .A4( u2_u15_u7_n157 ) , .A3( u2_u15_u7_n158 ) , .A2( u2_u15_u7_n159 ) , .A1( u2_u15_u7_n160 ) );
  AND3_X1 u2_u15_u7_U9 (.A3( u2_u15_u7_n110 ) , .A2( u2_u15_u7_n127 ) , .A1( u2_u15_u7_n132 ) , .ZN( u2_u15_u7_n92 ) );
  OAI21_X1 u2_u15_u7_U90 (.B1( u2_u15_u7_n145 ) , .ZN( u2_u15_u7_n160 ) , .A( u2_u15_u7_n161 ) , .B2( u2_u15_u7_n177 ) );
  OAI21_X1 u2_u15_u7_U91 (.ZN( u2_u15_u7_n159 ) , .A( u2_u15_u7_n165 ) , .B2( u2_u15_u7_n171 ) , .B1( u2_u15_u7_n174 ) );
  NAND4_X1 u2_u15_u7_U92 (.ZN( u2_out15_15 ) , .A4( u2_u15_u7_n142 ) , .A3( u2_u15_u7_n143 ) , .A2( u2_u15_u7_n144 ) , .A1( u2_u15_u7_n178 ) );
  OR2_X1 u2_u15_u7_U93 (.A2( u2_u15_u7_n125 ) , .A1( u2_u15_u7_n129 ) , .ZN( u2_u15_u7_n144 ) );
  AOI22_X1 u2_u15_u7_U94 (.A2( u2_u15_u7_n126 ) , .ZN( u2_u15_u7_n143 ) , .B2( u2_u15_u7_n165 ) , .B1( u2_u15_u7_n173 ) , .A1( u2_u15_u7_n174 ) );
  NAND3_X1 u2_u15_u7_U95 (.A3( u2_u15_u7_n146 ) , .A2( u2_u15_u7_n147 ) , .A1( u2_u15_u7_n148 ) , .ZN( u2_u15_u7_n151 ) );
  NAND3_X1 u2_u15_u7_U96 (.A3( u2_u15_u7_n131 ) , .A2( u2_u15_u7_n132 ) , .A1( u2_u15_u7_n133 ) , .ZN( u2_u15_u7_n135 ) );
  XOR2_X1 u2_u1_U13 (.B( u2_K2_42 ) , .A( u2_R0_29 ) , .Z( u2_u1_X_42 ) );
  XOR2_X1 u2_u1_U14 (.B( u2_K2_41 ) , .A( u2_R0_28 ) , .Z( u2_u1_X_41 ) );
  XOR2_X1 u2_u1_U15 (.B( u2_K2_40 ) , .A( u2_R0_27 ) , .Z( u2_u1_X_40 ) );
  XOR2_X1 u2_u1_U17 (.B( u2_K2_39 ) , .A( u2_R0_26 ) , .Z( u2_u1_X_39 ) );
  XOR2_X1 u2_u1_U18 (.B( u2_K2_38 ) , .A( u2_R0_25 ) , .Z( u2_u1_X_38 ) );
  XOR2_X1 u2_u1_U19 (.B( u2_K2_37 ) , .A( u2_R0_24 ) , .Z( u2_u1_X_37 ) );
  XOR2_X1 u2_u1_U26 (.B( u2_K2_30 ) , .A( u2_R0_21 ) , .Z( u2_u1_X_30 ) );
  XOR2_X1 u2_u1_U28 (.B( u2_K2_29 ) , .A( u2_R0_20 ) , .Z( u2_u1_X_29 ) );
  XOR2_X1 u2_u1_U29 (.B( u2_K2_28 ) , .A( u2_R0_19 ) , .Z( u2_u1_X_28 ) );
  XOR2_X1 u2_u1_U30 (.B( u2_K2_27 ) , .A( u2_R0_18 ) , .Z( u2_u1_X_27 ) );
  XOR2_X1 u2_u1_U31 (.B( u2_K2_26 ) , .A( u2_R0_17 ) , .Z( u2_u1_X_26 ) );
  XOR2_X1 u2_u1_U32 (.B( u2_K2_25 ) , .A( u2_R0_16 ) , .Z( u2_u1_X_25 ) );
  OAI22_X1 u2_u1_u4_U10 (.B2( u2_u1_u4_n135 ) , .ZN( u2_u1_u4_n137 ) , .B1( u2_u1_u4_n153 ) , .A1( u2_u1_u4_n155 ) , .A2( u2_u1_u4_n171 ) );
  AND3_X1 u2_u1_u4_U11 (.A2( u2_u1_u4_n134 ) , .ZN( u2_u1_u4_n135 ) , .A3( u2_u1_u4_n145 ) , .A1( u2_u1_u4_n157 ) );
  NAND2_X1 u2_u1_u4_U12 (.ZN( u2_u1_u4_n132 ) , .A2( u2_u1_u4_n170 ) , .A1( u2_u1_u4_n173 ) );
  AOI21_X1 u2_u1_u4_U13 (.B2( u2_u1_u4_n160 ) , .B1( u2_u1_u4_n161 ) , .ZN( u2_u1_u4_n162 ) , .A( u2_u1_u4_n170 ) );
  AOI21_X1 u2_u1_u4_U14 (.ZN( u2_u1_u4_n107 ) , .B2( u2_u1_u4_n143 ) , .A( u2_u1_u4_n174 ) , .B1( u2_u1_u4_n184 ) );
  AOI21_X1 u2_u1_u4_U15 (.B2( u2_u1_u4_n158 ) , .B1( u2_u1_u4_n159 ) , .ZN( u2_u1_u4_n163 ) , .A( u2_u1_u4_n174 ) );
  AOI21_X1 u2_u1_u4_U16 (.A( u2_u1_u4_n153 ) , .B2( u2_u1_u4_n154 ) , .B1( u2_u1_u4_n155 ) , .ZN( u2_u1_u4_n165 ) );
  AOI21_X1 u2_u1_u4_U17 (.A( u2_u1_u4_n156 ) , .B2( u2_u1_u4_n157 ) , .ZN( u2_u1_u4_n164 ) , .B1( u2_u1_u4_n184 ) );
  INV_X1 u2_u1_u4_U18 (.A( u2_u1_u4_n138 ) , .ZN( u2_u1_u4_n170 ) );
  AND2_X1 u2_u1_u4_U19 (.A2( u2_u1_u4_n120 ) , .ZN( u2_u1_u4_n155 ) , .A1( u2_u1_u4_n160 ) );
  INV_X1 u2_u1_u4_U20 (.A( u2_u1_u4_n156 ) , .ZN( u2_u1_u4_n175 ) );
  NAND2_X1 u2_u1_u4_U21 (.A2( u2_u1_u4_n118 ) , .ZN( u2_u1_u4_n131 ) , .A1( u2_u1_u4_n147 ) );
  NAND2_X1 u2_u1_u4_U22 (.A1( u2_u1_u4_n119 ) , .A2( u2_u1_u4_n120 ) , .ZN( u2_u1_u4_n130 ) );
  NAND2_X1 u2_u1_u4_U23 (.ZN( u2_u1_u4_n117 ) , .A2( u2_u1_u4_n118 ) , .A1( u2_u1_u4_n148 ) );
  NAND2_X1 u2_u1_u4_U24 (.ZN( u2_u1_u4_n129 ) , .A1( u2_u1_u4_n134 ) , .A2( u2_u1_u4_n148 ) );
  AND3_X1 u2_u1_u4_U25 (.A1( u2_u1_u4_n119 ) , .A2( u2_u1_u4_n143 ) , .A3( u2_u1_u4_n154 ) , .ZN( u2_u1_u4_n161 ) );
  AND2_X1 u2_u1_u4_U26 (.A1( u2_u1_u4_n145 ) , .A2( u2_u1_u4_n147 ) , .ZN( u2_u1_u4_n159 ) );
  OR3_X1 u2_u1_u4_U27 (.A3( u2_u1_u4_n114 ) , .A2( u2_u1_u4_n115 ) , .A1( u2_u1_u4_n116 ) , .ZN( u2_u1_u4_n136 ) );
  AOI21_X1 u2_u1_u4_U28 (.A( u2_u1_u4_n113 ) , .ZN( u2_u1_u4_n116 ) , .B2( u2_u1_u4_n173 ) , .B1( u2_u1_u4_n174 ) );
  AOI21_X1 u2_u1_u4_U29 (.ZN( u2_u1_u4_n115 ) , .B2( u2_u1_u4_n145 ) , .B1( u2_u1_u4_n146 ) , .A( u2_u1_u4_n156 ) );
  NOR2_X1 u2_u1_u4_U3 (.ZN( u2_u1_u4_n121 ) , .A1( u2_u1_u4_n181 ) , .A2( u2_u1_u4_n182 ) );
  OAI22_X1 u2_u1_u4_U30 (.ZN( u2_u1_u4_n114 ) , .A2( u2_u1_u4_n121 ) , .B1( u2_u1_u4_n160 ) , .B2( u2_u1_u4_n170 ) , .A1( u2_u1_u4_n171 ) );
  INV_X1 u2_u1_u4_U31 (.A( u2_u1_u4_n158 ) , .ZN( u2_u1_u4_n182 ) );
  INV_X1 u2_u1_u4_U32 (.ZN( u2_u1_u4_n181 ) , .A( u2_u1_u4_n96 ) );
  INV_X1 u2_u1_u4_U33 (.A( u2_u1_u4_n144 ) , .ZN( u2_u1_u4_n179 ) );
  INV_X1 u2_u1_u4_U34 (.A( u2_u1_u4_n157 ) , .ZN( u2_u1_u4_n178 ) );
  NAND2_X1 u2_u1_u4_U35 (.A2( u2_u1_u4_n154 ) , .A1( u2_u1_u4_n96 ) , .ZN( u2_u1_u4_n97 ) );
  INV_X1 u2_u1_u4_U36 (.ZN( u2_u1_u4_n186 ) , .A( u2_u1_u4_n95 ) );
  OAI221_X1 u2_u1_u4_U37 (.C1( u2_u1_u4_n134 ) , .B1( u2_u1_u4_n158 ) , .B2( u2_u1_u4_n171 ) , .C2( u2_u1_u4_n173 ) , .A( u2_u1_u4_n94 ) , .ZN( u2_u1_u4_n95 ) );
  AOI222_X1 u2_u1_u4_U38 (.B2( u2_u1_u4_n132 ) , .A1( u2_u1_u4_n138 ) , .C2( u2_u1_u4_n175 ) , .A2( u2_u1_u4_n179 ) , .C1( u2_u1_u4_n181 ) , .B1( u2_u1_u4_n185 ) , .ZN( u2_u1_u4_n94 ) );
  INV_X1 u2_u1_u4_U39 (.A( u2_u1_u4_n113 ) , .ZN( u2_u1_u4_n185 ) );
  INV_X1 u2_u1_u4_U4 (.A( u2_u1_u4_n117 ) , .ZN( u2_u1_u4_n184 ) );
  INV_X1 u2_u1_u4_U40 (.A( u2_u1_u4_n143 ) , .ZN( u2_u1_u4_n183 ) );
  NOR2_X1 u2_u1_u4_U41 (.ZN( u2_u1_u4_n138 ) , .A1( u2_u1_u4_n168 ) , .A2( u2_u1_u4_n169 ) );
  NOR2_X1 u2_u1_u4_U42 (.A1( u2_u1_u4_n150 ) , .A2( u2_u1_u4_n152 ) , .ZN( u2_u1_u4_n153 ) );
  NOR2_X1 u2_u1_u4_U43 (.A2( u2_u1_u4_n128 ) , .A1( u2_u1_u4_n138 ) , .ZN( u2_u1_u4_n156 ) );
  AOI22_X1 u2_u1_u4_U44 (.B2( u2_u1_u4_n122 ) , .A1( u2_u1_u4_n123 ) , .ZN( u2_u1_u4_n124 ) , .B1( u2_u1_u4_n128 ) , .A2( u2_u1_u4_n172 ) );
  NAND2_X1 u2_u1_u4_U45 (.A2( u2_u1_u4_n120 ) , .ZN( u2_u1_u4_n123 ) , .A1( u2_u1_u4_n161 ) );
  INV_X1 u2_u1_u4_U46 (.A( u2_u1_u4_n153 ) , .ZN( u2_u1_u4_n172 ) );
  AOI22_X1 u2_u1_u4_U47 (.B2( u2_u1_u4_n132 ) , .A2( u2_u1_u4_n133 ) , .ZN( u2_u1_u4_n140 ) , .A1( u2_u1_u4_n150 ) , .B1( u2_u1_u4_n179 ) );
  NAND2_X1 u2_u1_u4_U48 (.ZN( u2_u1_u4_n133 ) , .A2( u2_u1_u4_n146 ) , .A1( u2_u1_u4_n154 ) );
  NAND2_X1 u2_u1_u4_U49 (.A1( u2_u1_u4_n103 ) , .ZN( u2_u1_u4_n154 ) , .A2( u2_u1_u4_n98 ) );
  NOR4_X1 u2_u1_u4_U5 (.A4( u2_u1_u4_n106 ) , .A3( u2_u1_u4_n107 ) , .A2( u2_u1_u4_n108 ) , .A1( u2_u1_u4_n109 ) , .ZN( u2_u1_u4_n110 ) );
  NAND2_X1 u2_u1_u4_U50 (.A1( u2_u1_u4_n101 ) , .ZN( u2_u1_u4_n158 ) , .A2( u2_u1_u4_n99 ) );
  AOI21_X1 u2_u1_u4_U51 (.ZN( u2_u1_u4_n127 ) , .A( u2_u1_u4_n136 ) , .B2( u2_u1_u4_n150 ) , .B1( u2_u1_u4_n180 ) );
  INV_X1 u2_u1_u4_U52 (.A( u2_u1_u4_n160 ) , .ZN( u2_u1_u4_n180 ) );
  NAND2_X1 u2_u1_u4_U53 (.A2( u2_u1_u4_n104 ) , .A1( u2_u1_u4_n105 ) , .ZN( u2_u1_u4_n146 ) );
  NAND2_X1 u2_u1_u4_U54 (.A2( u2_u1_u4_n101 ) , .A1( u2_u1_u4_n102 ) , .ZN( u2_u1_u4_n160 ) );
  NAND2_X1 u2_u1_u4_U55 (.ZN( u2_u1_u4_n134 ) , .A1( u2_u1_u4_n98 ) , .A2( u2_u1_u4_n99 ) );
  NAND2_X1 u2_u1_u4_U56 (.A1( u2_u1_u4_n103 ) , .A2( u2_u1_u4_n104 ) , .ZN( u2_u1_u4_n143 ) );
  NAND2_X1 u2_u1_u4_U57 (.A2( u2_u1_u4_n105 ) , .ZN( u2_u1_u4_n145 ) , .A1( u2_u1_u4_n98 ) );
  NAND2_X1 u2_u1_u4_U58 (.A1( u2_u1_u4_n100 ) , .A2( u2_u1_u4_n105 ) , .ZN( u2_u1_u4_n120 ) );
  NAND2_X1 u2_u1_u4_U59 (.A1( u2_u1_u4_n102 ) , .A2( u2_u1_u4_n104 ) , .ZN( u2_u1_u4_n148 ) );
  AOI21_X1 u2_u1_u4_U6 (.ZN( u2_u1_u4_n106 ) , .B2( u2_u1_u4_n146 ) , .B1( u2_u1_u4_n158 ) , .A( u2_u1_u4_n170 ) );
  NAND2_X1 u2_u1_u4_U60 (.A2( u2_u1_u4_n100 ) , .A1( u2_u1_u4_n103 ) , .ZN( u2_u1_u4_n157 ) );
  INV_X1 u2_u1_u4_U61 (.A( u2_u1_u4_n150 ) , .ZN( u2_u1_u4_n173 ) );
  INV_X1 u2_u1_u4_U62 (.A( u2_u1_u4_n152 ) , .ZN( u2_u1_u4_n171 ) );
  NAND2_X1 u2_u1_u4_U63 (.A1( u2_u1_u4_n100 ) , .ZN( u2_u1_u4_n118 ) , .A2( u2_u1_u4_n99 ) );
  NAND2_X1 u2_u1_u4_U64 (.A2( u2_u1_u4_n100 ) , .A1( u2_u1_u4_n102 ) , .ZN( u2_u1_u4_n144 ) );
  NAND2_X1 u2_u1_u4_U65 (.A2( u2_u1_u4_n101 ) , .A1( u2_u1_u4_n105 ) , .ZN( u2_u1_u4_n96 ) );
  INV_X1 u2_u1_u4_U66 (.A( u2_u1_u4_n128 ) , .ZN( u2_u1_u4_n174 ) );
  NAND2_X1 u2_u1_u4_U67 (.A2( u2_u1_u4_n102 ) , .ZN( u2_u1_u4_n119 ) , .A1( u2_u1_u4_n98 ) );
  NAND2_X1 u2_u1_u4_U68 (.A2( u2_u1_u4_n101 ) , .A1( u2_u1_u4_n103 ) , .ZN( u2_u1_u4_n147 ) );
  NAND2_X1 u2_u1_u4_U69 (.A2( u2_u1_u4_n104 ) , .ZN( u2_u1_u4_n113 ) , .A1( u2_u1_u4_n99 ) );
  AOI21_X1 u2_u1_u4_U7 (.ZN( u2_u1_u4_n108 ) , .B2( u2_u1_u4_n134 ) , .B1( u2_u1_u4_n155 ) , .A( u2_u1_u4_n156 ) );
  NOR2_X1 u2_u1_u4_U70 (.A2( u2_u1_X_28 ) , .ZN( u2_u1_u4_n150 ) , .A1( u2_u1_u4_n168 ) );
  NOR2_X1 u2_u1_u4_U71 (.A2( u2_u1_X_29 ) , .ZN( u2_u1_u4_n152 ) , .A1( u2_u1_u4_n169 ) );
  NOR2_X1 u2_u1_u4_U72 (.A2( u2_u1_X_30 ) , .ZN( u2_u1_u4_n105 ) , .A1( u2_u1_u4_n176 ) );
  NOR2_X1 u2_u1_u4_U73 (.A2( u2_u1_X_26 ) , .ZN( u2_u1_u4_n100 ) , .A1( u2_u1_u4_n177 ) );
  NOR2_X1 u2_u1_u4_U74 (.A2( u2_u1_X_28 ) , .A1( u2_u1_X_29 ) , .ZN( u2_u1_u4_n128 ) );
  NOR2_X1 u2_u1_u4_U75 (.A2( u2_u1_X_27 ) , .A1( u2_u1_X_30 ) , .ZN( u2_u1_u4_n102 ) );
  NOR2_X1 u2_u1_u4_U76 (.A2( u2_u1_X_25 ) , .A1( u2_u1_X_26 ) , .ZN( u2_u1_u4_n98 ) );
  AND2_X1 u2_u1_u4_U77 (.A2( u2_u1_X_25 ) , .A1( u2_u1_X_26 ) , .ZN( u2_u1_u4_n104 ) );
  AND2_X1 u2_u1_u4_U78 (.A1( u2_u1_X_30 ) , .A2( u2_u1_u4_n176 ) , .ZN( u2_u1_u4_n99 ) );
  AND2_X1 u2_u1_u4_U79 (.A1( u2_u1_X_26 ) , .ZN( u2_u1_u4_n101 ) , .A2( u2_u1_u4_n177 ) );
  AOI21_X1 u2_u1_u4_U8 (.ZN( u2_u1_u4_n109 ) , .A( u2_u1_u4_n153 ) , .B1( u2_u1_u4_n159 ) , .B2( u2_u1_u4_n184 ) );
  AND2_X1 u2_u1_u4_U80 (.A1( u2_u1_X_27 ) , .A2( u2_u1_X_30 ) , .ZN( u2_u1_u4_n103 ) );
  INV_X1 u2_u1_u4_U81 (.A( u2_u1_X_28 ) , .ZN( u2_u1_u4_n169 ) );
  INV_X1 u2_u1_u4_U82 (.A( u2_u1_X_29 ) , .ZN( u2_u1_u4_n168 ) );
  INV_X1 u2_u1_u4_U83 (.A( u2_u1_X_25 ) , .ZN( u2_u1_u4_n177 ) );
  INV_X1 u2_u1_u4_U84 (.A( u2_u1_X_27 ) , .ZN( u2_u1_u4_n176 ) );
  NAND4_X1 u2_u1_u4_U85 (.ZN( u2_out1_25 ) , .A4( u2_u1_u4_n139 ) , .A3( u2_u1_u4_n140 ) , .A2( u2_u1_u4_n141 ) , .A1( u2_u1_u4_n142 ) );
  OAI21_X1 u2_u1_u4_U86 (.A( u2_u1_u4_n128 ) , .B2( u2_u1_u4_n129 ) , .B1( u2_u1_u4_n130 ) , .ZN( u2_u1_u4_n142 ) );
  OAI21_X1 u2_u1_u4_U87 (.B2( u2_u1_u4_n131 ) , .ZN( u2_u1_u4_n141 ) , .A( u2_u1_u4_n175 ) , .B1( u2_u1_u4_n183 ) );
  NAND4_X1 u2_u1_u4_U88 (.ZN( u2_out1_14 ) , .A4( u2_u1_u4_n124 ) , .A3( u2_u1_u4_n125 ) , .A2( u2_u1_u4_n126 ) , .A1( u2_u1_u4_n127 ) );
  AOI22_X1 u2_u1_u4_U89 (.B2( u2_u1_u4_n117 ) , .ZN( u2_u1_u4_n126 ) , .A1( u2_u1_u4_n129 ) , .B1( u2_u1_u4_n152 ) , .A2( u2_u1_u4_n175 ) );
  AOI211_X1 u2_u1_u4_U9 (.B( u2_u1_u4_n136 ) , .A( u2_u1_u4_n137 ) , .C2( u2_u1_u4_n138 ) , .ZN( u2_u1_u4_n139 ) , .C1( u2_u1_u4_n182 ) );
  AOI22_X1 u2_u1_u4_U90 (.ZN( u2_u1_u4_n125 ) , .B2( u2_u1_u4_n131 ) , .A2( u2_u1_u4_n132 ) , .B1( u2_u1_u4_n138 ) , .A1( u2_u1_u4_n178 ) );
  NAND4_X1 u2_u1_u4_U91 (.ZN( u2_out1_8 ) , .A4( u2_u1_u4_n110 ) , .A3( u2_u1_u4_n111 ) , .A2( u2_u1_u4_n112 ) , .A1( u2_u1_u4_n186 ) );
  NAND2_X1 u2_u1_u4_U92 (.ZN( u2_u1_u4_n112 ) , .A2( u2_u1_u4_n130 ) , .A1( u2_u1_u4_n150 ) );
  AOI22_X1 u2_u1_u4_U93 (.ZN( u2_u1_u4_n111 ) , .B2( u2_u1_u4_n132 ) , .A1( u2_u1_u4_n152 ) , .B1( u2_u1_u4_n178 ) , .A2( u2_u1_u4_n97 ) );
  AOI22_X1 u2_u1_u4_U94 (.B2( u2_u1_u4_n149 ) , .B1( u2_u1_u4_n150 ) , .A2( u2_u1_u4_n151 ) , .A1( u2_u1_u4_n152 ) , .ZN( u2_u1_u4_n167 ) );
  NOR4_X1 u2_u1_u4_U95 (.A4( u2_u1_u4_n162 ) , .A3( u2_u1_u4_n163 ) , .A2( u2_u1_u4_n164 ) , .A1( u2_u1_u4_n165 ) , .ZN( u2_u1_u4_n166 ) );
  NAND3_X1 u2_u1_u4_U96 (.ZN( u2_out1_3 ) , .A3( u2_u1_u4_n166 ) , .A1( u2_u1_u4_n167 ) , .A2( u2_u1_u4_n186 ) );
  NAND3_X1 u2_u1_u4_U97 (.A3( u2_u1_u4_n146 ) , .A2( u2_u1_u4_n147 ) , .A1( u2_u1_u4_n148 ) , .ZN( u2_u1_u4_n149 ) );
  NAND3_X1 u2_u1_u4_U98 (.A3( u2_u1_u4_n143 ) , .A2( u2_u1_u4_n144 ) , .A1( u2_u1_u4_n145 ) , .ZN( u2_u1_u4_n151 ) );
  NAND3_X1 u2_u1_u4_U99 (.A3( u2_u1_u4_n121 ) , .ZN( u2_u1_u4_n122 ) , .A2( u2_u1_u4_n144 ) , .A1( u2_u1_u4_n154 ) );
  AOI22_X1 u2_u1_u6_U10 (.A2( u2_u1_u6_n151 ) , .B2( u2_u1_u6_n161 ) , .A1( u2_u1_u6_n167 ) , .B1( u2_u1_u6_n170 ) , .ZN( u2_u1_u6_n89 ) );
  AOI21_X1 u2_u1_u6_U11 (.B1( u2_u1_u6_n107 ) , .B2( u2_u1_u6_n132 ) , .A( u2_u1_u6_n158 ) , .ZN( u2_u1_u6_n88 ) );
  AOI21_X1 u2_u1_u6_U12 (.B2( u2_u1_u6_n147 ) , .B1( u2_u1_u6_n148 ) , .ZN( u2_u1_u6_n149 ) , .A( u2_u1_u6_n158 ) );
  AOI21_X1 u2_u1_u6_U13 (.ZN( u2_u1_u6_n106 ) , .A( u2_u1_u6_n142 ) , .B2( u2_u1_u6_n159 ) , .B1( u2_u1_u6_n164 ) );
  INV_X1 u2_u1_u6_U14 (.A( u2_u1_u6_n155 ) , .ZN( u2_u1_u6_n161 ) );
  INV_X1 u2_u1_u6_U15 (.A( u2_u1_u6_n128 ) , .ZN( u2_u1_u6_n164 ) );
  NAND2_X1 u2_u1_u6_U16 (.ZN( u2_u1_u6_n110 ) , .A1( u2_u1_u6_n122 ) , .A2( u2_u1_u6_n129 ) );
  NAND2_X1 u2_u1_u6_U17 (.ZN( u2_u1_u6_n124 ) , .A2( u2_u1_u6_n146 ) , .A1( u2_u1_u6_n148 ) );
  INV_X1 u2_u1_u6_U18 (.A( u2_u1_u6_n132 ) , .ZN( u2_u1_u6_n171 ) );
  AND2_X1 u2_u1_u6_U19 (.A1( u2_u1_u6_n100 ) , .ZN( u2_u1_u6_n130 ) , .A2( u2_u1_u6_n147 ) );
  INV_X1 u2_u1_u6_U20 (.A( u2_u1_u6_n127 ) , .ZN( u2_u1_u6_n173 ) );
  INV_X1 u2_u1_u6_U21 (.A( u2_u1_u6_n121 ) , .ZN( u2_u1_u6_n167 ) );
  INV_X1 u2_u1_u6_U22 (.A( u2_u1_u6_n100 ) , .ZN( u2_u1_u6_n169 ) );
  INV_X1 u2_u1_u6_U23 (.A( u2_u1_u6_n123 ) , .ZN( u2_u1_u6_n170 ) );
  INV_X1 u2_u1_u6_U24 (.A( u2_u1_u6_n113 ) , .ZN( u2_u1_u6_n168 ) );
  AND2_X1 u2_u1_u6_U25 (.A1( u2_u1_u6_n107 ) , .A2( u2_u1_u6_n119 ) , .ZN( u2_u1_u6_n133 ) );
  AND2_X1 u2_u1_u6_U26 (.A2( u2_u1_u6_n121 ) , .A1( u2_u1_u6_n122 ) , .ZN( u2_u1_u6_n131 ) );
  AND3_X1 u2_u1_u6_U27 (.ZN( u2_u1_u6_n120 ) , .A2( u2_u1_u6_n127 ) , .A1( u2_u1_u6_n132 ) , .A3( u2_u1_u6_n145 ) );
  INV_X1 u2_u1_u6_U28 (.A( u2_u1_u6_n146 ) , .ZN( u2_u1_u6_n163 ) );
  AOI222_X1 u2_u1_u6_U29 (.ZN( u2_u1_u6_n114 ) , .A1( u2_u1_u6_n118 ) , .A2( u2_u1_u6_n126 ) , .B2( u2_u1_u6_n151 ) , .C2( u2_u1_u6_n159 ) , .C1( u2_u1_u6_n168 ) , .B1( u2_u1_u6_n169 ) );
  INV_X1 u2_u1_u6_U3 (.A( u2_u1_u6_n110 ) , .ZN( u2_u1_u6_n166 ) );
  NOR2_X1 u2_u1_u6_U30 (.A1( u2_u1_u6_n162 ) , .A2( u2_u1_u6_n165 ) , .ZN( u2_u1_u6_n98 ) );
  AOI211_X1 u2_u1_u6_U31 (.B( u2_u1_u6_n134 ) , .A( u2_u1_u6_n135 ) , .C1( u2_u1_u6_n136 ) , .ZN( u2_u1_u6_n137 ) , .C2( u2_u1_u6_n151 ) );
  AOI21_X1 u2_u1_u6_U32 (.B1( u2_u1_u6_n131 ) , .ZN( u2_u1_u6_n135 ) , .A( u2_u1_u6_n144 ) , .B2( u2_u1_u6_n146 ) );
  NAND4_X1 u2_u1_u6_U33 (.A4( u2_u1_u6_n127 ) , .A3( u2_u1_u6_n128 ) , .A2( u2_u1_u6_n129 ) , .A1( u2_u1_u6_n130 ) , .ZN( u2_u1_u6_n136 ) );
  AOI21_X1 u2_u1_u6_U34 (.B2( u2_u1_u6_n132 ) , .B1( u2_u1_u6_n133 ) , .ZN( u2_u1_u6_n134 ) , .A( u2_u1_u6_n158 ) );
  NAND2_X1 u2_u1_u6_U35 (.A1( u2_u1_u6_n144 ) , .ZN( u2_u1_u6_n151 ) , .A2( u2_u1_u6_n158 ) );
  NAND2_X1 u2_u1_u6_U36 (.ZN( u2_u1_u6_n132 ) , .A1( u2_u1_u6_n91 ) , .A2( u2_u1_u6_n97 ) );
  AOI22_X1 u2_u1_u6_U37 (.B2( u2_u1_u6_n110 ) , .B1( u2_u1_u6_n111 ) , .A1( u2_u1_u6_n112 ) , .ZN( u2_u1_u6_n115 ) , .A2( u2_u1_u6_n161 ) );
  NAND4_X1 u2_u1_u6_U38 (.A3( u2_u1_u6_n109 ) , .ZN( u2_u1_u6_n112 ) , .A4( u2_u1_u6_n132 ) , .A2( u2_u1_u6_n147 ) , .A1( u2_u1_u6_n166 ) );
  NOR2_X1 u2_u1_u6_U39 (.ZN( u2_u1_u6_n109 ) , .A1( u2_u1_u6_n170 ) , .A2( u2_u1_u6_n173 ) );
  INV_X1 u2_u1_u6_U4 (.A( u2_u1_u6_n142 ) , .ZN( u2_u1_u6_n174 ) );
  NOR2_X1 u2_u1_u6_U40 (.A2( u2_u1_u6_n126 ) , .ZN( u2_u1_u6_n155 ) , .A1( u2_u1_u6_n160 ) );
  NAND2_X1 u2_u1_u6_U41 (.ZN( u2_u1_u6_n146 ) , .A2( u2_u1_u6_n94 ) , .A1( u2_u1_u6_n99 ) );
  AOI21_X1 u2_u1_u6_U42 (.A( u2_u1_u6_n144 ) , .B2( u2_u1_u6_n145 ) , .B1( u2_u1_u6_n146 ) , .ZN( u2_u1_u6_n150 ) );
  INV_X1 u2_u1_u6_U43 (.A( u2_u1_u6_n111 ) , .ZN( u2_u1_u6_n158 ) );
  NAND2_X1 u2_u1_u6_U44 (.ZN( u2_u1_u6_n127 ) , .A1( u2_u1_u6_n91 ) , .A2( u2_u1_u6_n92 ) );
  NAND2_X1 u2_u1_u6_U45 (.ZN( u2_u1_u6_n129 ) , .A2( u2_u1_u6_n95 ) , .A1( u2_u1_u6_n96 ) );
  INV_X1 u2_u1_u6_U46 (.A( u2_u1_u6_n144 ) , .ZN( u2_u1_u6_n159 ) );
  NAND2_X1 u2_u1_u6_U47 (.ZN( u2_u1_u6_n145 ) , .A2( u2_u1_u6_n97 ) , .A1( u2_u1_u6_n98 ) );
  NAND2_X1 u2_u1_u6_U48 (.ZN( u2_u1_u6_n148 ) , .A2( u2_u1_u6_n92 ) , .A1( u2_u1_u6_n94 ) );
  NAND2_X1 u2_u1_u6_U49 (.ZN( u2_u1_u6_n108 ) , .A2( u2_u1_u6_n139 ) , .A1( u2_u1_u6_n144 ) );
  NAND2_X1 u2_u1_u6_U5 (.A2( u2_u1_u6_n143 ) , .ZN( u2_u1_u6_n152 ) , .A1( u2_u1_u6_n166 ) );
  NAND2_X1 u2_u1_u6_U50 (.ZN( u2_u1_u6_n121 ) , .A2( u2_u1_u6_n95 ) , .A1( u2_u1_u6_n97 ) );
  NAND2_X1 u2_u1_u6_U51 (.ZN( u2_u1_u6_n107 ) , .A2( u2_u1_u6_n92 ) , .A1( u2_u1_u6_n95 ) );
  AND2_X1 u2_u1_u6_U52 (.ZN( u2_u1_u6_n118 ) , .A2( u2_u1_u6_n91 ) , .A1( u2_u1_u6_n99 ) );
  NAND2_X1 u2_u1_u6_U53 (.ZN( u2_u1_u6_n147 ) , .A2( u2_u1_u6_n98 ) , .A1( u2_u1_u6_n99 ) );
  NAND2_X1 u2_u1_u6_U54 (.ZN( u2_u1_u6_n128 ) , .A1( u2_u1_u6_n94 ) , .A2( u2_u1_u6_n96 ) );
  NAND2_X1 u2_u1_u6_U55 (.ZN( u2_u1_u6_n119 ) , .A2( u2_u1_u6_n95 ) , .A1( u2_u1_u6_n99 ) );
  NAND2_X1 u2_u1_u6_U56 (.ZN( u2_u1_u6_n123 ) , .A2( u2_u1_u6_n91 ) , .A1( u2_u1_u6_n96 ) );
  NAND2_X1 u2_u1_u6_U57 (.ZN( u2_u1_u6_n100 ) , .A2( u2_u1_u6_n92 ) , .A1( u2_u1_u6_n98 ) );
  NAND2_X1 u2_u1_u6_U58 (.ZN( u2_u1_u6_n122 ) , .A1( u2_u1_u6_n94 ) , .A2( u2_u1_u6_n97 ) );
  INV_X1 u2_u1_u6_U59 (.A( u2_u1_u6_n139 ) , .ZN( u2_u1_u6_n160 ) );
  AOI22_X1 u2_u1_u6_U6 (.B2( u2_u1_u6_n101 ) , .A1( u2_u1_u6_n102 ) , .ZN( u2_u1_u6_n103 ) , .B1( u2_u1_u6_n160 ) , .A2( u2_u1_u6_n161 ) );
  NAND2_X1 u2_u1_u6_U60 (.ZN( u2_u1_u6_n113 ) , .A1( u2_u1_u6_n96 ) , .A2( u2_u1_u6_n98 ) );
  NOR2_X1 u2_u1_u6_U61 (.A2( u2_u1_X_40 ) , .A1( u2_u1_X_41 ) , .ZN( u2_u1_u6_n126 ) );
  NOR2_X1 u2_u1_u6_U62 (.A2( u2_u1_X_39 ) , .A1( u2_u1_X_42 ) , .ZN( u2_u1_u6_n92 ) );
  NOR2_X1 u2_u1_u6_U63 (.A2( u2_u1_X_39 ) , .A1( u2_u1_u6_n156 ) , .ZN( u2_u1_u6_n97 ) );
  NOR2_X1 u2_u1_u6_U64 (.A2( u2_u1_X_38 ) , .A1( u2_u1_u6_n165 ) , .ZN( u2_u1_u6_n95 ) );
  NOR2_X1 u2_u1_u6_U65 (.A2( u2_u1_X_41 ) , .ZN( u2_u1_u6_n111 ) , .A1( u2_u1_u6_n157 ) );
  NOR2_X1 u2_u1_u6_U66 (.A2( u2_u1_X_37 ) , .A1( u2_u1_u6_n162 ) , .ZN( u2_u1_u6_n94 ) );
  NOR2_X1 u2_u1_u6_U67 (.A2( u2_u1_X_37 ) , .A1( u2_u1_X_38 ) , .ZN( u2_u1_u6_n91 ) );
  NAND2_X1 u2_u1_u6_U68 (.A1( u2_u1_X_41 ) , .ZN( u2_u1_u6_n144 ) , .A2( u2_u1_u6_n157 ) );
  NAND2_X1 u2_u1_u6_U69 (.A2( u2_u1_X_40 ) , .A1( u2_u1_X_41 ) , .ZN( u2_u1_u6_n139 ) );
  NOR2_X1 u2_u1_u6_U7 (.A1( u2_u1_u6_n118 ) , .ZN( u2_u1_u6_n143 ) , .A2( u2_u1_u6_n168 ) );
  AND2_X1 u2_u1_u6_U70 (.A1( u2_u1_X_39 ) , .A2( u2_u1_u6_n156 ) , .ZN( u2_u1_u6_n96 ) );
  AND2_X1 u2_u1_u6_U71 (.A1( u2_u1_X_39 ) , .A2( u2_u1_X_42 ) , .ZN( u2_u1_u6_n99 ) );
  INV_X1 u2_u1_u6_U72 (.A( u2_u1_X_40 ) , .ZN( u2_u1_u6_n157 ) );
  INV_X1 u2_u1_u6_U73 (.A( u2_u1_X_37 ) , .ZN( u2_u1_u6_n165 ) );
  INV_X1 u2_u1_u6_U74 (.A( u2_u1_X_38 ) , .ZN( u2_u1_u6_n162 ) );
  INV_X1 u2_u1_u6_U75 (.A( u2_u1_X_42 ) , .ZN( u2_u1_u6_n156 ) );
  NAND4_X1 u2_u1_u6_U76 (.ZN( u2_out1_32 ) , .A4( u2_u1_u6_n103 ) , .A3( u2_u1_u6_n104 ) , .A2( u2_u1_u6_n105 ) , .A1( u2_u1_u6_n106 ) );
  AOI22_X1 u2_u1_u6_U77 (.ZN( u2_u1_u6_n105 ) , .A2( u2_u1_u6_n108 ) , .A1( u2_u1_u6_n118 ) , .B2( u2_u1_u6_n126 ) , .B1( u2_u1_u6_n171 ) );
  AOI22_X1 u2_u1_u6_U78 (.ZN( u2_u1_u6_n104 ) , .A1( u2_u1_u6_n111 ) , .B1( u2_u1_u6_n124 ) , .B2( u2_u1_u6_n151 ) , .A2( u2_u1_u6_n93 ) );
  NAND4_X1 u2_u1_u6_U79 (.ZN( u2_out1_12 ) , .A4( u2_u1_u6_n114 ) , .A3( u2_u1_u6_n115 ) , .A2( u2_u1_u6_n116 ) , .A1( u2_u1_u6_n117 ) );
  OAI21_X1 u2_u1_u6_U8 (.A( u2_u1_u6_n159 ) , .B1( u2_u1_u6_n169 ) , .B2( u2_u1_u6_n173 ) , .ZN( u2_u1_u6_n90 ) );
  OAI22_X1 u2_u1_u6_U80 (.B2( u2_u1_u6_n111 ) , .ZN( u2_u1_u6_n116 ) , .B1( u2_u1_u6_n126 ) , .A2( u2_u1_u6_n164 ) , .A1( u2_u1_u6_n167 ) );
  OAI21_X1 u2_u1_u6_U81 (.A( u2_u1_u6_n108 ) , .ZN( u2_u1_u6_n117 ) , .B2( u2_u1_u6_n141 ) , .B1( u2_u1_u6_n163 ) );
  OAI211_X1 u2_u1_u6_U82 (.ZN( u2_out1_22 ) , .B( u2_u1_u6_n137 ) , .A( u2_u1_u6_n138 ) , .C2( u2_u1_u6_n139 ) , .C1( u2_u1_u6_n140 ) );
  AND4_X1 u2_u1_u6_U83 (.A3( u2_u1_u6_n119 ) , .A1( u2_u1_u6_n120 ) , .A4( u2_u1_u6_n129 ) , .ZN( u2_u1_u6_n140 ) , .A2( u2_u1_u6_n143 ) );
  AOI22_X1 u2_u1_u6_U84 (.B1( u2_u1_u6_n124 ) , .A2( u2_u1_u6_n125 ) , .A1( u2_u1_u6_n126 ) , .ZN( u2_u1_u6_n138 ) , .B2( u2_u1_u6_n161 ) );
  OAI211_X1 u2_u1_u6_U85 (.ZN( u2_out1_7 ) , .B( u2_u1_u6_n153 ) , .C2( u2_u1_u6_n154 ) , .C1( u2_u1_u6_n155 ) , .A( u2_u1_u6_n174 ) );
  NOR3_X1 u2_u1_u6_U86 (.A1( u2_u1_u6_n141 ) , .ZN( u2_u1_u6_n154 ) , .A3( u2_u1_u6_n164 ) , .A2( u2_u1_u6_n171 ) );
  AOI211_X1 u2_u1_u6_U87 (.B( u2_u1_u6_n149 ) , .A( u2_u1_u6_n150 ) , .C2( u2_u1_u6_n151 ) , .C1( u2_u1_u6_n152 ) , .ZN( u2_u1_u6_n153 ) );
  NAND3_X1 u2_u1_u6_U88 (.A2( u2_u1_u6_n123 ) , .ZN( u2_u1_u6_n125 ) , .A1( u2_u1_u6_n130 ) , .A3( u2_u1_u6_n131 ) );
  NAND3_X1 u2_u1_u6_U89 (.A3( u2_u1_u6_n133 ) , .ZN( u2_u1_u6_n141 ) , .A1( u2_u1_u6_n145 ) , .A2( u2_u1_u6_n148 ) );
  INV_X1 u2_u1_u6_U9 (.ZN( u2_u1_u6_n172 ) , .A( u2_u1_u6_n88 ) );
  NAND3_X1 u2_u1_u6_U90 (.ZN( u2_u1_u6_n101 ) , .A3( u2_u1_u6_n107 ) , .A2( u2_u1_u6_n121 ) , .A1( u2_u1_u6_n127 ) );
  NAND3_X1 u2_u1_u6_U91 (.ZN( u2_u1_u6_n102 ) , .A3( u2_u1_u6_n130 ) , .A2( u2_u1_u6_n145 ) , .A1( u2_u1_u6_n166 ) );
  NAND3_X1 u2_u1_u6_U92 (.A3( u2_u1_u6_n113 ) , .A1( u2_u1_u6_n119 ) , .A2( u2_u1_u6_n123 ) , .ZN( u2_u1_u6_n93 ) );
  NAND3_X1 u2_u1_u6_U93 (.ZN( u2_u1_u6_n142 ) , .A2( u2_u1_u6_n172 ) , .A3( u2_u1_u6_n89 ) , .A1( u2_u1_u6_n90 ) );
  XOR2_X1 u2_u2_U1 (.B( u2_K3_9 ) , .A( u2_R1_6 ) , .Z( u2_u2_X_9 ) );
  XOR2_X1 u2_u2_U10 (.B( u2_K3_45 ) , .A( u2_R1_30 ) , .Z( u2_u2_X_45 ) );
  XOR2_X1 u2_u2_U11 (.B( u2_K3_44 ) , .A( u2_R1_29 ) , .Z( u2_u2_X_44 ) );
  XOR2_X1 u2_u2_U12 (.B( u2_K3_43 ) , .A( u2_R1_28 ) , .Z( u2_u2_X_43 ) );
  XOR2_X1 u2_u2_U13 (.B( u2_K3_42 ) , .A( u2_R1_29 ) , .Z( u2_u2_X_42 ) );
  XOR2_X1 u2_u2_U14 (.B( u2_K3_41 ) , .A( u2_R1_28 ) , .Z( u2_u2_X_41 ) );
  XOR2_X1 u2_u2_U15 (.B( u2_K3_40 ) , .A( u2_R1_27 ) , .Z( u2_u2_X_40 ) );
  XOR2_X1 u2_u2_U16 (.B( u2_K3_3 ) , .A( u2_R1_2 ) , .Z( u2_u2_X_3 ) );
  XOR2_X1 u2_u2_U17 (.B( u2_K3_39 ) , .A( u2_R1_26 ) , .Z( u2_u2_X_39 ) );
  XOR2_X1 u2_u2_U18 (.B( u2_K3_38 ) , .A( u2_R1_25 ) , .Z( u2_u2_X_38 ) );
  XOR2_X1 u2_u2_U19 (.B( u2_K3_37 ) , .A( u2_R1_24 ) , .Z( u2_u2_X_37 ) );
  XOR2_X1 u2_u2_U2 (.B( u2_K3_8 ) , .A( u2_R1_5 ) , .Z( u2_u2_X_8 ) );
  XOR2_X1 u2_u2_U20 (.B( u2_K3_36 ) , .A( u2_R1_25 ) , .Z( u2_u2_X_36 ) );
  XOR2_X1 u2_u2_U21 (.B( u2_K3_35 ) , .A( u2_R1_24 ) , .Z( u2_u2_X_35 ) );
  XOR2_X1 u2_u2_U22 (.B( u2_K3_34 ) , .A( u2_R1_23 ) , .Z( u2_u2_X_34 ) );
  XOR2_X1 u2_u2_U23 (.B( u2_K3_33 ) , .A( u2_R1_22 ) , .Z( u2_u2_X_33 ) );
  XOR2_X1 u2_u2_U24 (.B( u2_K3_32 ) , .A( u2_R1_21 ) , .Z( u2_u2_X_32 ) );
  XOR2_X1 u2_u2_U25 (.B( u2_K3_31 ) , .A( u2_R1_20 ) , .Z( u2_u2_X_31 ) );
  XOR2_X1 u2_u2_U27 (.B( u2_K3_2 ) , .A( u2_R1_1 ) , .Z( u2_u2_X_2 ) );
  XOR2_X1 u2_u2_U3 (.B( u2_K3_7 ) , .A( u2_R1_4 ) , .Z( u2_u2_X_7 ) );
  XOR2_X1 u2_u2_U33 (.B( u2_K3_24 ) , .A( u2_R1_17 ) , .Z( u2_u2_X_24 ) );
  XOR2_X1 u2_u2_U34 (.B( u2_K3_23 ) , .A( u2_R1_16 ) , .Z( u2_u2_X_23 ) );
  XOR2_X1 u2_u2_U35 (.B( u2_K3_22 ) , .A( u2_R1_15 ) , .Z( u2_u2_X_22 ) );
  XOR2_X1 u2_u2_U36 (.B( u2_K3_21 ) , .A( u2_R1_14 ) , .Z( u2_u2_X_21 ) );
  XOR2_X1 u2_u2_U37 (.B( u2_K3_20 ) , .A( u2_R1_13 ) , .Z( u2_u2_X_20 ) );
  XOR2_X1 u2_u2_U38 (.B( u2_K3_1 ) , .A( u2_R1_32 ) , .Z( u2_u2_X_1 ) );
  XOR2_X1 u2_u2_U39 (.B( u2_K3_19 ) , .A( u2_R1_12 ) , .Z( u2_u2_X_19 ) );
  XOR2_X1 u2_u2_U4 (.B( u2_K3_6 ) , .A( u2_R1_5 ) , .Z( u2_u2_X_6 ) );
  XOR2_X1 u2_u2_U40 (.B( u2_K3_18 ) , .A( u2_R1_13 ) , .Z( u2_u2_X_18 ) );
  XOR2_X1 u2_u2_U41 (.B( u2_K3_17 ) , .A( u2_R1_12 ) , .Z( u2_u2_X_17 ) );
  XOR2_X1 u2_u2_U42 (.B( u2_K3_16 ) , .A( u2_R1_11 ) , .Z( u2_u2_X_16 ) );
  XOR2_X1 u2_u2_U43 (.B( u2_K3_15 ) , .A( u2_R1_10 ) , .Z( u2_u2_X_15 ) );
  XOR2_X1 u2_u2_U44 (.B( u2_K3_14 ) , .A( u2_R1_9 ) , .Z( u2_u2_X_14 ) );
  XOR2_X1 u2_u2_U45 (.B( u2_K3_13 ) , .A( u2_R1_8 ) , .Z( u2_u2_X_13 ) );
  XOR2_X1 u2_u2_U46 (.B( u2_K3_12 ) , .A( u2_R1_9 ) , .Z( u2_u2_X_12 ) );
  XOR2_X1 u2_u2_U47 (.B( u2_K3_11 ) , .A( u2_R1_8 ) , .Z( u2_u2_X_11 ) );
  XOR2_X1 u2_u2_U48 (.B( u2_K3_10 ) , .A( u2_R1_7 ) , .Z( u2_u2_X_10 ) );
  XOR2_X1 u2_u2_U5 (.B( u2_K3_5 ) , .A( u2_R1_4 ) , .Z( u2_u2_X_5 ) );
  XOR2_X1 u2_u2_U6 (.B( u2_K3_4 ) , .A( u2_R1_3 ) , .Z( u2_u2_X_4 ) );
  XOR2_X1 u2_u2_U7 (.B( u2_K3_48 ) , .A( u2_R1_1 ) , .Z( u2_u2_X_48 ) );
  XOR2_X1 u2_u2_U8 (.B( u2_K3_47 ) , .A( u2_R1_32 ) , .Z( u2_u2_X_47 ) );
  XOR2_X1 u2_u2_U9 (.B( u2_K3_46 ) , .A( u2_R1_31 ) , .Z( u2_u2_X_46 ) );
  AND3_X1 u2_u2_u0_U10 (.A2( u2_u2_u0_n112 ) , .ZN( u2_u2_u0_n127 ) , .A3( u2_u2_u0_n130 ) , .A1( u2_u2_u0_n148 ) );
  NAND2_X1 u2_u2_u0_U11 (.ZN( u2_u2_u0_n113 ) , .A1( u2_u2_u0_n139 ) , .A2( u2_u2_u0_n149 ) );
  AND2_X1 u2_u2_u0_U12 (.ZN( u2_u2_u0_n107 ) , .A1( u2_u2_u0_n130 ) , .A2( u2_u2_u0_n140 ) );
  AND2_X1 u2_u2_u0_U13 (.A2( u2_u2_u0_n129 ) , .A1( u2_u2_u0_n130 ) , .ZN( u2_u2_u0_n151 ) );
  AND2_X1 u2_u2_u0_U14 (.A1( u2_u2_u0_n108 ) , .A2( u2_u2_u0_n125 ) , .ZN( u2_u2_u0_n145 ) );
  INV_X1 u2_u2_u0_U15 (.A( u2_u2_u0_n143 ) , .ZN( u2_u2_u0_n173 ) );
  NOR2_X1 u2_u2_u0_U16 (.A2( u2_u2_u0_n136 ) , .ZN( u2_u2_u0_n147 ) , .A1( u2_u2_u0_n160 ) );
  INV_X1 u2_u2_u0_U17 (.ZN( u2_u2_u0_n172 ) , .A( u2_u2_u0_n88 ) );
  OAI222_X1 u2_u2_u0_U18 (.C1( u2_u2_u0_n108 ) , .A1( u2_u2_u0_n125 ) , .B2( u2_u2_u0_n128 ) , .B1( u2_u2_u0_n144 ) , .A2( u2_u2_u0_n158 ) , .C2( u2_u2_u0_n161 ) , .ZN( u2_u2_u0_n88 ) );
  NOR2_X1 u2_u2_u0_U19 (.A1( u2_u2_u0_n163 ) , .A2( u2_u2_u0_n164 ) , .ZN( u2_u2_u0_n95 ) );
  AOI21_X1 u2_u2_u0_U20 (.B1( u2_u2_u0_n103 ) , .ZN( u2_u2_u0_n132 ) , .A( u2_u2_u0_n165 ) , .B2( u2_u2_u0_n93 ) );
  INV_X1 u2_u2_u0_U21 (.A( u2_u2_u0_n142 ) , .ZN( u2_u2_u0_n165 ) );
  OAI221_X1 u2_u2_u0_U22 (.C1( u2_u2_u0_n121 ) , .ZN( u2_u2_u0_n122 ) , .B2( u2_u2_u0_n127 ) , .A( u2_u2_u0_n143 ) , .B1( u2_u2_u0_n144 ) , .C2( u2_u2_u0_n147 ) );
  OAI22_X1 u2_u2_u0_U23 (.B1( u2_u2_u0_n125 ) , .ZN( u2_u2_u0_n126 ) , .A1( u2_u2_u0_n138 ) , .A2( u2_u2_u0_n146 ) , .B2( u2_u2_u0_n147 ) );
  OAI22_X1 u2_u2_u0_U24 (.B1( u2_u2_u0_n131 ) , .A1( u2_u2_u0_n144 ) , .B2( u2_u2_u0_n147 ) , .A2( u2_u2_u0_n90 ) , .ZN( u2_u2_u0_n91 ) );
  AND3_X1 u2_u2_u0_U25 (.A3( u2_u2_u0_n121 ) , .A2( u2_u2_u0_n125 ) , .A1( u2_u2_u0_n148 ) , .ZN( u2_u2_u0_n90 ) );
  INV_X1 u2_u2_u0_U26 (.A( u2_u2_u0_n136 ) , .ZN( u2_u2_u0_n161 ) );
  NOR2_X1 u2_u2_u0_U27 (.A1( u2_u2_u0_n120 ) , .ZN( u2_u2_u0_n143 ) , .A2( u2_u2_u0_n167 ) );
  OAI221_X1 u2_u2_u0_U28 (.C1( u2_u2_u0_n112 ) , .ZN( u2_u2_u0_n120 ) , .B1( u2_u2_u0_n138 ) , .B2( u2_u2_u0_n141 ) , .C2( u2_u2_u0_n147 ) , .A( u2_u2_u0_n172 ) );
  AOI211_X1 u2_u2_u0_U29 (.B( u2_u2_u0_n115 ) , .A( u2_u2_u0_n116 ) , .C2( u2_u2_u0_n117 ) , .C1( u2_u2_u0_n118 ) , .ZN( u2_u2_u0_n119 ) );
  INV_X1 u2_u2_u0_U3 (.A( u2_u2_u0_n113 ) , .ZN( u2_u2_u0_n166 ) );
  AOI22_X1 u2_u2_u0_U30 (.B2( u2_u2_u0_n109 ) , .A2( u2_u2_u0_n110 ) , .ZN( u2_u2_u0_n111 ) , .B1( u2_u2_u0_n118 ) , .A1( u2_u2_u0_n160 ) );
  INV_X1 u2_u2_u0_U31 (.A( u2_u2_u0_n118 ) , .ZN( u2_u2_u0_n158 ) );
  AOI21_X1 u2_u2_u0_U32 (.ZN( u2_u2_u0_n104 ) , .B1( u2_u2_u0_n107 ) , .B2( u2_u2_u0_n141 ) , .A( u2_u2_u0_n144 ) );
  AOI21_X1 u2_u2_u0_U33 (.B1( u2_u2_u0_n127 ) , .B2( u2_u2_u0_n129 ) , .A( u2_u2_u0_n138 ) , .ZN( u2_u2_u0_n96 ) );
  AOI21_X1 u2_u2_u0_U34 (.ZN( u2_u2_u0_n116 ) , .B2( u2_u2_u0_n142 ) , .A( u2_u2_u0_n144 ) , .B1( u2_u2_u0_n166 ) );
  NAND2_X1 u2_u2_u0_U35 (.A1( u2_u2_u0_n100 ) , .A2( u2_u2_u0_n103 ) , .ZN( u2_u2_u0_n125 ) );
  NAND2_X1 u2_u2_u0_U36 (.A1( u2_u2_u0_n101 ) , .A2( u2_u2_u0_n102 ) , .ZN( u2_u2_u0_n150 ) );
  INV_X1 u2_u2_u0_U37 (.A( u2_u2_u0_n138 ) , .ZN( u2_u2_u0_n160 ) );
  NAND2_X1 u2_u2_u0_U38 (.A1( u2_u2_u0_n102 ) , .ZN( u2_u2_u0_n128 ) , .A2( u2_u2_u0_n95 ) );
  NAND2_X1 u2_u2_u0_U39 (.A1( u2_u2_u0_n100 ) , .ZN( u2_u2_u0_n129 ) , .A2( u2_u2_u0_n95 ) );
  AOI21_X1 u2_u2_u0_U4 (.B1( u2_u2_u0_n114 ) , .ZN( u2_u2_u0_n115 ) , .B2( u2_u2_u0_n129 ) , .A( u2_u2_u0_n161 ) );
  NAND2_X1 u2_u2_u0_U40 (.A2( u2_u2_u0_n100 ) , .ZN( u2_u2_u0_n131 ) , .A1( u2_u2_u0_n92 ) );
  NAND2_X1 u2_u2_u0_U41 (.A2( u2_u2_u0_n100 ) , .A1( u2_u2_u0_n101 ) , .ZN( u2_u2_u0_n139 ) );
  NAND2_X1 u2_u2_u0_U42 (.ZN( u2_u2_u0_n148 ) , .A1( u2_u2_u0_n93 ) , .A2( u2_u2_u0_n95 ) );
  NAND2_X1 u2_u2_u0_U43 (.A2( u2_u2_u0_n102 ) , .A1( u2_u2_u0_n103 ) , .ZN( u2_u2_u0_n149 ) );
  NAND2_X1 u2_u2_u0_U44 (.A2( u2_u2_u0_n102 ) , .ZN( u2_u2_u0_n114 ) , .A1( u2_u2_u0_n92 ) );
  NAND2_X1 u2_u2_u0_U45 (.A2( u2_u2_u0_n101 ) , .ZN( u2_u2_u0_n121 ) , .A1( u2_u2_u0_n93 ) );
  NAND2_X1 u2_u2_u0_U46 (.ZN( u2_u2_u0_n112 ) , .A2( u2_u2_u0_n92 ) , .A1( u2_u2_u0_n93 ) );
  OR3_X1 u2_u2_u0_U47 (.A3( u2_u2_u0_n152 ) , .A2( u2_u2_u0_n153 ) , .A1( u2_u2_u0_n154 ) , .ZN( u2_u2_u0_n155 ) );
  AOI21_X1 u2_u2_u0_U48 (.B2( u2_u2_u0_n150 ) , .B1( u2_u2_u0_n151 ) , .ZN( u2_u2_u0_n152 ) , .A( u2_u2_u0_n158 ) );
  AOI21_X1 u2_u2_u0_U49 (.A( u2_u2_u0_n144 ) , .B2( u2_u2_u0_n145 ) , .B1( u2_u2_u0_n146 ) , .ZN( u2_u2_u0_n154 ) );
  AOI21_X1 u2_u2_u0_U5 (.B2( u2_u2_u0_n131 ) , .ZN( u2_u2_u0_n134 ) , .B1( u2_u2_u0_n151 ) , .A( u2_u2_u0_n158 ) );
  AOI21_X1 u2_u2_u0_U50 (.A( u2_u2_u0_n147 ) , .B2( u2_u2_u0_n148 ) , .B1( u2_u2_u0_n149 ) , .ZN( u2_u2_u0_n153 ) );
  INV_X1 u2_u2_u0_U51 (.ZN( u2_u2_u0_n171 ) , .A( u2_u2_u0_n99 ) );
  OAI211_X1 u2_u2_u0_U52 (.C2( u2_u2_u0_n140 ) , .C1( u2_u2_u0_n161 ) , .A( u2_u2_u0_n169 ) , .B( u2_u2_u0_n98 ) , .ZN( u2_u2_u0_n99 ) );
  INV_X1 u2_u2_u0_U53 (.ZN( u2_u2_u0_n169 ) , .A( u2_u2_u0_n91 ) );
  AOI211_X1 u2_u2_u0_U54 (.C1( u2_u2_u0_n118 ) , .A( u2_u2_u0_n123 ) , .B( u2_u2_u0_n96 ) , .C2( u2_u2_u0_n97 ) , .ZN( u2_u2_u0_n98 ) );
  NOR2_X1 u2_u2_u0_U55 (.A2( u2_u2_X_6 ) , .ZN( u2_u2_u0_n100 ) , .A1( u2_u2_u0_n162 ) );
  NOR2_X1 u2_u2_u0_U56 (.A2( u2_u2_X_4 ) , .A1( u2_u2_X_5 ) , .ZN( u2_u2_u0_n118 ) );
  NOR2_X1 u2_u2_u0_U57 (.A2( u2_u2_X_2 ) , .ZN( u2_u2_u0_n103 ) , .A1( u2_u2_u0_n164 ) );
  NOR2_X1 u2_u2_u0_U58 (.A2( u2_u2_X_1 ) , .A1( u2_u2_X_2 ) , .ZN( u2_u2_u0_n92 ) );
  NOR2_X1 u2_u2_u0_U59 (.A2( u2_u2_X_1 ) , .ZN( u2_u2_u0_n101 ) , .A1( u2_u2_u0_n163 ) );
  NOR2_X1 u2_u2_u0_U6 (.A1( u2_u2_u0_n108 ) , .ZN( u2_u2_u0_n123 ) , .A2( u2_u2_u0_n158 ) );
  NAND2_X1 u2_u2_u0_U60 (.A2( u2_u2_X_4 ) , .A1( u2_u2_X_5 ) , .ZN( u2_u2_u0_n144 ) );
  NOR2_X1 u2_u2_u0_U61 (.A2( u2_u2_X_5 ) , .ZN( u2_u2_u0_n136 ) , .A1( u2_u2_u0_n159 ) );
  NAND2_X1 u2_u2_u0_U62 (.A1( u2_u2_X_5 ) , .ZN( u2_u2_u0_n138 ) , .A2( u2_u2_u0_n159 ) );
  NOR2_X1 u2_u2_u0_U63 (.A2( u2_u2_X_3 ) , .A1( u2_u2_X_6 ) , .ZN( u2_u2_u0_n94 ) );
  AND2_X1 u2_u2_u0_U64 (.A2( u2_u2_X_3 ) , .A1( u2_u2_X_6 ) , .ZN( u2_u2_u0_n102 ) );
  AND2_X1 u2_u2_u0_U65 (.A1( u2_u2_X_6 ) , .A2( u2_u2_u0_n162 ) , .ZN( u2_u2_u0_n93 ) );
  INV_X1 u2_u2_u0_U66 (.A( u2_u2_X_4 ) , .ZN( u2_u2_u0_n159 ) );
  INV_X1 u2_u2_u0_U67 (.A( u2_u2_X_1 ) , .ZN( u2_u2_u0_n164 ) );
  INV_X1 u2_u2_u0_U68 (.A( u2_u2_X_2 ) , .ZN( u2_u2_u0_n163 ) );
  INV_X1 u2_u2_u0_U69 (.A( u2_u2_X_3 ) , .ZN( u2_u2_u0_n162 ) );
  OAI21_X1 u2_u2_u0_U7 (.B1( u2_u2_u0_n150 ) , .B2( u2_u2_u0_n158 ) , .A( u2_u2_u0_n172 ) , .ZN( u2_u2_u0_n89 ) );
  INV_X1 u2_u2_u0_U70 (.A( u2_u2_u0_n126 ) , .ZN( u2_u2_u0_n168 ) );
  AOI211_X1 u2_u2_u0_U71 (.B( u2_u2_u0_n133 ) , .A( u2_u2_u0_n134 ) , .C2( u2_u2_u0_n135 ) , .C1( u2_u2_u0_n136 ) , .ZN( u2_u2_u0_n137 ) );
  INV_X1 u2_u2_u0_U72 (.ZN( u2_u2_u0_n174 ) , .A( u2_u2_u0_n89 ) );
  AOI211_X1 u2_u2_u0_U73 (.B( u2_u2_u0_n104 ) , .A( u2_u2_u0_n105 ) , .ZN( u2_u2_u0_n106 ) , .C2( u2_u2_u0_n113 ) , .C1( u2_u2_u0_n160 ) );
  OR4_X1 u2_u2_u0_U74 (.ZN( u2_out2_17 ) , .A4( u2_u2_u0_n122 ) , .A2( u2_u2_u0_n123 ) , .A1( u2_u2_u0_n124 ) , .A3( u2_u2_u0_n170 ) );
  AOI21_X1 u2_u2_u0_U75 (.B2( u2_u2_u0_n107 ) , .ZN( u2_u2_u0_n124 ) , .B1( u2_u2_u0_n128 ) , .A( u2_u2_u0_n161 ) );
  INV_X1 u2_u2_u0_U76 (.A( u2_u2_u0_n111 ) , .ZN( u2_u2_u0_n170 ) );
  OR4_X1 u2_u2_u0_U77 (.ZN( u2_out2_31 ) , .A4( u2_u2_u0_n155 ) , .A2( u2_u2_u0_n156 ) , .A1( u2_u2_u0_n157 ) , .A3( u2_u2_u0_n173 ) );
  AOI21_X1 u2_u2_u0_U78 (.A( u2_u2_u0_n138 ) , .B2( u2_u2_u0_n139 ) , .B1( u2_u2_u0_n140 ) , .ZN( u2_u2_u0_n157 ) );
  AOI21_X1 u2_u2_u0_U79 (.B2( u2_u2_u0_n141 ) , .B1( u2_u2_u0_n142 ) , .ZN( u2_u2_u0_n156 ) , .A( u2_u2_u0_n161 ) );
  AND2_X1 u2_u2_u0_U8 (.A1( u2_u2_u0_n114 ) , .A2( u2_u2_u0_n121 ) , .ZN( u2_u2_u0_n146 ) );
  AOI21_X1 u2_u2_u0_U80 (.B1( u2_u2_u0_n132 ) , .ZN( u2_u2_u0_n133 ) , .A( u2_u2_u0_n144 ) , .B2( u2_u2_u0_n166 ) );
  OAI22_X1 u2_u2_u0_U81 (.ZN( u2_u2_u0_n105 ) , .A2( u2_u2_u0_n132 ) , .B1( u2_u2_u0_n146 ) , .A1( u2_u2_u0_n147 ) , .B2( u2_u2_u0_n161 ) );
  NAND2_X1 u2_u2_u0_U82 (.ZN( u2_u2_u0_n110 ) , .A2( u2_u2_u0_n132 ) , .A1( u2_u2_u0_n145 ) );
  INV_X1 u2_u2_u0_U83 (.A( u2_u2_u0_n119 ) , .ZN( u2_u2_u0_n167 ) );
  NAND2_X1 u2_u2_u0_U84 (.A2( u2_u2_u0_n103 ) , .ZN( u2_u2_u0_n140 ) , .A1( u2_u2_u0_n94 ) );
  NAND2_X1 u2_u2_u0_U85 (.A1( u2_u2_u0_n101 ) , .ZN( u2_u2_u0_n130 ) , .A2( u2_u2_u0_n94 ) );
  NAND2_X1 u2_u2_u0_U86 (.ZN( u2_u2_u0_n108 ) , .A1( u2_u2_u0_n92 ) , .A2( u2_u2_u0_n94 ) );
  NAND2_X1 u2_u2_u0_U87 (.ZN( u2_u2_u0_n142 ) , .A1( u2_u2_u0_n94 ) , .A2( u2_u2_u0_n95 ) );
  NAND3_X1 u2_u2_u0_U88 (.ZN( u2_out2_23 ) , .A3( u2_u2_u0_n137 ) , .A1( u2_u2_u0_n168 ) , .A2( u2_u2_u0_n171 ) );
  NAND3_X1 u2_u2_u0_U89 (.A3( u2_u2_u0_n127 ) , .A2( u2_u2_u0_n128 ) , .ZN( u2_u2_u0_n135 ) , .A1( u2_u2_u0_n150 ) );
  AND2_X1 u2_u2_u0_U9 (.A1( u2_u2_u0_n131 ) , .ZN( u2_u2_u0_n141 ) , .A2( u2_u2_u0_n150 ) );
  NAND3_X1 u2_u2_u0_U90 (.ZN( u2_u2_u0_n117 ) , .A3( u2_u2_u0_n132 ) , .A2( u2_u2_u0_n139 ) , .A1( u2_u2_u0_n148 ) );
  NAND3_X1 u2_u2_u0_U91 (.ZN( u2_u2_u0_n109 ) , .A2( u2_u2_u0_n114 ) , .A3( u2_u2_u0_n140 ) , .A1( u2_u2_u0_n149 ) );
  NAND3_X1 u2_u2_u0_U92 (.ZN( u2_out2_9 ) , .A3( u2_u2_u0_n106 ) , .A2( u2_u2_u0_n171 ) , .A1( u2_u2_u0_n174 ) );
  NAND3_X1 u2_u2_u0_U93 (.A2( u2_u2_u0_n128 ) , .A1( u2_u2_u0_n132 ) , .A3( u2_u2_u0_n146 ) , .ZN( u2_u2_u0_n97 ) );
  NOR2_X1 u2_u2_u1_U10 (.A1( u2_u2_u1_n112 ) , .A2( u2_u2_u1_n116 ) , .ZN( u2_u2_u1_n118 ) );
  NAND3_X1 u2_u2_u1_U100 (.ZN( u2_u2_u1_n113 ) , .A1( u2_u2_u1_n120 ) , .A3( u2_u2_u1_n133 ) , .A2( u2_u2_u1_n155 ) );
  OAI21_X1 u2_u2_u1_U11 (.ZN( u2_u2_u1_n101 ) , .B1( u2_u2_u1_n141 ) , .A( u2_u2_u1_n146 ) , .B2( u2_u2_u1_n183 ) );
  AOI21_X1 u2_u2_u1_U12 (.B2( u2_u2_u1_n155 ) , .B1( u2_u2_u1_n156 ) , .ZN( u2_u2_u1_n157 ) , .A( u2_u2_u1_n174 ) );
  OR4_X1 u2_u2_u1_U13 (.A4( u2_u2_u1_n106 ) , .A3( u2_u2_u1_n107 ) , .ZN( u2_u2_u1_n108 ) , .A1( u2_u2_u1_n117 ) , .A2( u2_u2_u1_n184 ) );
  AOI21_X1 u2_u2_u1_U14 (.ZN( u2_u2_u1_n106 ) , .A( u2_u2_u1_n112 ) , .B1( u2_u2_u1_n154 ) , .B2( u2_u2_u1_n156 ) );
  INV_X1 u2_u2_u1_U15 (.A( u2_u2_u1_n101 ) , .ZN( u2_u2_u1_n184 ) );
  AOI21_X1 u2_u2_u1_U16 (.ZN( u2_u2_u1_n107 ) , .B1( u2_u2_u1_n134 ) , .B2( u2_u2_u1_n149 ) , .A( u2_u2_u1_n174 ) );
  NAND2_X1 u2_u2_u1_U17 (.ZN( u2_u2_u1_n140 ) , .A2( u2_u2_u1_n150 ) , .A1( u2_u2_u1_n155 ) );
  NAND2_X1 u2_u2_u1_U18 (.A1( u2_u2_u1_n131 ) , .ZN( u2_u2_u1_n147 ) , .A2( u2_u2_u1_n153 ) );
  INV_X1 u2_u2_u1_U19 (.A( u2_u2_u1_n139 ) , .ZN( u2_u2_u1_n174 ) );
  INV_X1 u2_u2_u1_U20 (.A( u2_u2_u1_n112 ) , .ZN( u2_u2_u1_n171 ) );
  NAND2_X1 u2_u2_u1_U21 (.ZN( u2_u2_u1_n141 ) , .A1( u2_u2_u1_n153 ) , .A2( u2_u2_u1_n156 ) );
  AND2_X1 u2_u2_u1_U22 (.A1( u2_u2_u1_n123 ) , .ZN( u2_u2_u1_n134 ) , .A2( u2_u2_u1_n161 ) );
  NAND2_X1 u2_u2_u1_U23 (.A2( u2_u2_u1_n115 ) , .A1( u2_u2_u1_n116 ) , .ZN( u2_u2_u1_n148 ) );
  NAND2_X1 u2_u2_u1_U24 (.A2( u2_u2_u1_n133 ) , .A1( u2_u2_u1_n135 ) , .ZN( u2_u2_u1_n159 ) );
  NAND2_X1 u2_u2_u1_U25 (.A2( u2_u2_u1_n115 ) , .A1( u2_u2_u1_n120 ) , .ZN( u2_u2_u1_n132 ) );
  INV_X1 u2_u2_u1_U26 (.A( u2_u2_u1_n154 ) , .ZN( u2_u2_u1_n178 ) );
  INV_X1 u2_u2_u1_U27 (.A( u2_u2_u1_n151 ) , .ZN( u2_u2_u1_n183 ) );
  AND2_X1 u2_u2_u1_U28 (.A1( u2_u2_u1_n129 ) , .A2( u2_u2_u1_n133 ) , .ZN( u2_u2_u1_n149 ) );
  INV_X1 u2_u2_u1_U29 (.A( u2_u2_u1_n131 ) , .ZN( u2_u2_u1_n180 ) );
  INV_X1 u2_u2_u1_U3 (.A( u2_u2_u1_n159 ) , .ZN( u2_u2_u1_n182 ) );
  OAI221_X1 u2_u2_u1_U30 (.A( u2_u2_u1_n119 ) , .C2( u2_u2_u1_n129 ) , .ZN( u2_u2_u1_n138 ) , .B2( u2_u2_u1_n152 ) , .C1( u2_u2_u1_n174 ) , .B1( u2_u2_u1_n187 ) );
  INV_X1 u2_u2_u1_U31 (.A( u2_u2_u1_n148 ) , .ZN( u2_u2_u1_n187 ) );
  AOI211_X1 u2_u2_u1_U32 (.B( u2_u2_u1_n117 ) , .A( u2_u2_u1_n118 ) , .ZN( u2_u2_u1_n119 ) , .C2( u2_u2_u1_n146 ) , .C1( u2_u2_u1_n159 ) );
  NOR2_X1 u2_u2_u1_U33 (.A1( u2_u2_u1_n168 ) , .A2( u2_u2_u1_n176 ) , .ZN( u2_u2_u1_n98 ) );
  AOI211_X1 u2_u2_u1_U34 (.B( u2_u2_u1_n162 ) , .A( u2_u2_u1_n163 ) , .C2( u2_u2_u1_n164 ) , .ZN( u2_u2_u1_n165 ) , .C1( u2_u2_u1_n171 ) );
  AOI21_X1 u2_u2_u1_U35 (.A( u2_u2_u1_n160 ) , .B2( u2_u2_u1_n161 ) , .ZN( u2_u2_u1_n162 ) , .B1( u2_u2_u1_n182 ) );
  OR2_X1 u2_u2_u1_U36 (.A2( u2_u2_u1_n157 ) , .A1( u2_u2_u1_n158 ) , .ZN( u2_u2_u1_n163 ) );
  OAI21_X1 u2_u2_u1_U37 (.B2( u2_u2_u1_n123 ) , .ZN( u2_u2_u1_n145 ) , .B1( u2_u2_u1_n160 ) , .A( u2_u2_u1_n185 ) );
  INV_X1 u2_u2_u1_U38 (.A( u2_u2_u1_n122 ) , .ZN( u2_u2_u1_n185 ) );
  AOI21_X1 u2_u2_u1_U39 (.B2( u2_u2_u1_n120 ) , .B1( u2_u2_u1_n121 ) , .ZN( u2_u2_u1_n122 ) , .A( u2_u2_u1_n128 ) );
  AOI221_X1 u2_u2_u1_U4 (.A( u2_u2_u1_n138 ) , .C2( u2_u2_u1_n139 ) , .C1( u2_u2_u1_n140 ) , .B2( u2_u2_u1_n141 ) , .ZN( u2_u2_u1_n142 ) , .B1( u2_u2_u1_n175 ) );
  NAND2_X1 u2_u2_u1_U40 (.A1( u2_u2_u1_n128 ) , .ZN( u2_u2_u1_n146 ) , .A2( u2_u2_u1_n160 ) );
  NAND2_X1 u2_u2_u1_U41 (.A2( u2_u2_u1_n112 ) , .ZN( u2_u2_u1_n139 ) , .A1( u2_u2_u1_n152 ) );
  NAND2_X1 u2_u2_u1_U42 (.A1( u2_u2_u1_n105 ) , .ZN( u2_u2_u1_n156 ) , .A2( u2_u2_u1_n99 ) );
  AOI221_X1 u2_u2_u1_U43 (.B1( u2_u2_u1_n140 ) , .ZN( u2_u2_u1_n167 ) , .B2( u2_u2_u1_n172 ) , .C2( u2_u2_u1_n175 ) , .C1( u2_u2_u1_n178 ) , .A( u2_u2_u1_n188 ) );
  INV_X1 u2_u2_u1_U44 (.ZN( u2_u2_u1_n188 ) , .A( u2_u2_u1_n97 ) );
  AOI211_X1 u2_u2_u1_U45 (.A( u2_u2_u1_n118 ) , .C1( u2_u2_u1_n132 ) , .C2( u2_u2_u1_n139 ) , .B( u2_u2_u1_n96 ) , .ZN( u2_u2_u1_n97 ) );
  AOI21_X1 u2_u2_u1_U46 (.B2( u2_u2_u1_n121 ) , .B1( u2_u2_u1_n135 ) , .A( u2_u2_u1_n152 ) , .ZN( u2_u2_u1_n96 ) );
  NOR2_X1 u2_u2_u1_U47 (.ZN( u2_u2_u1_n117 ) , .A1( u2_u2_u1_n121 ) , .A2( u2_u2_u1_n160 ) );
  AOI21_X1 u2_u2_u1_U48 (.A( u2_u2_u1_n128 ) , .B2( u2_u2_u1_n129 ) , .ZN( u2_u2_u1_n130 ) , .B1( u2_u2_u1_n150 ) );
  NAND2_X1 u2_u2_u1_U49 (.ZN( u2_u2_u1_n112 ) , .A1( u2_u2_u1_n169 ) , .A2( u2_u2_u1_n170 ) );
  AOI211_X1 u2_u2_u1_U5 (.ZN( u2_u2_u1_n124 ) , .A( u2_u2_u1_n138 ) , .C2( u2_u2_u1_n139 ) , .B( u2_u2_u1_n145 ) , .C1( u2_u2_u1_n147 ) );
  NAND2_X1 u2_u2_u1_U50 (.ZN( u2_u2_u1_n129 ) , .A2( u2_u2_u1_n95 ) , .A1( u2_u2_u1_n98 ) );
  NAND2_X1 u2_u2_u1_U51 (.A1( u2_u2_u1_n102 ) , .ZN( u2_u2_u1_n154 ) , .A2( u2_u2_u1_n99 ) );
  NAND2_X1 u2_u2_u1_U52 (.A2( u2_u2_u1_n100 ) , .ZN( u2_u2_u1_n135 ) , .A1( u2_u2_u1_n99 ) );
  AOI21_X1 u2_u2_u1_U53 (.A( u2_u2_u1_n152 ) , .B2( u2_u2_u1_n153 ) , .B1( u2_u2_u1_n154 ) , .ZN( u2_u2_u1_n158 ) );
  INV_X1 u2_u2_u1_U54 (.A( u2_u2_u1_n160 ) , .ZN( u2_u2_u1_n175 ) );
  NAND2_X1 u2_u2_u1_U55 (.A1( u2_u2_u1_n100 ) , .ZN( u2_u2_u1_n116 ) , .A2( u2_u2_u1_n95 ) );
  NAND2_X1 u2_u2_u1_U56 (.A1( u2_u2_u1_n102 ) , .ZN( u2_u2_u1_n131 ) , .A2( u2_u2_u1_n95 ) );
  NAND2_X1 u2_u2_u1_U57 (.A2( u2_u2_u1_n104 ) , .ZN( u2_u2_u1_n121 ) , .A1( u2_u2_u1_n98 ) );
  NAND2_X1 u2_u2_u1_U58 (.A1( u2_u2_u1_n103 ) , .ZN( u2_u2_u1_n153 ) , .A2( u2_u2_u1_n98 ) );
  NAND2_X1 u2_u2_u1_U59 (.A2( u2_u2_u1_n104 ) , .A1( u2_u2_u1_n105 ) , .ZN( u2_u2_u1_n133 ) );
  AOI22_X1 u2_u2_u1_U6 (.B2( u2_u2_u1_n113 ) , .A2( u2_u2_u1_n114 ) , .ZN( u2_u2_u1_n125 ) , .A1( u2_u2_u1_n171 ) , .B1( u2_u2_u1_n173 ) );
  NAND2_X1 u2_u2_u1_U60 (.ZN( u2_u2_u1_n150 ) , .A2( u2_u2_u1_n98 ) , .A1( u2_u2_u1_n99 ) );
  NAND2_X1 u2_u2_u1_U61 (.A1( u2_u2_u1_n105 ) , .ZN( u2_u2_u1_n155 ) , .A2( u2_u2_u1_n95 ) );
  OAI21_X1 u2_u2_u1_U62 (.ZN( u2_u2_u1_n109 ) , .B1( u2_u2_u1_n129 ) , .B2( u2_u2_u1_n160 ) , .A( u2_u2_u1_n167 ) );
  NAND2_X1 u2_u2_u1_U63 (.A2( u2_u2_u1_n100 ) , .A1( u2_u2_u1_n103 ) , .ZN( u2_u2_u1_n120 ) );
  NAND2_X1 u2_u2_u1_U64 (.A1( u2_u2_u1_n102 ) , .A2( u2_u2_u1_n104 ) , .ZN( u2_u2_u1_n115 ) );
  NAND2_X1 u2_u2_u1_U65 (.A2( u2_u2_u1_n100 ) , .A1( u2_u2_u1_n104 ) , .ZN( u2_u2_u1_n151 ) );
  NAND2_X1 u2_u2_u1_U66 (.A2( u2_u2_u1_n103 ) , .A1( u2_u2_u1_n105 ) , .ZN( u2_u2_u1_n161 ) );
  INV_X1 u2_u2_u1_U67 (.A( u2_u2_u1_n152 ) , .ZN( u2_u2_u1_n173 ) );
  INV_X1 u2_u2_u1_U68 (.A( u2_u2_u1_n128 ) , .ZN( u2_u2_u1_n172 ) );
  NAND2_X1 u2_u2_u1_U69 (.A2( u2_u2_u1_n102 ) , .A1( u2_u2_u1_n103 ) , .ZN( u2_u2_u1_n123 ) );
  NAND2_X1 u2_u2_u1_U7 (.ZN( u2_u2_u1_n114 ) , .A1( u2_u2_u1_n134 ) , .A2( u2_u2_u1_n156 ) );
  NOR2_X1 u2_u2_u1_U70 (.A2( u2_u2_X_7 ) , .A1( u2_u2_X_8 ) , .ZN( u2_u2_u1_n95 ) );
  NOR2_X1 u2_u2_u1_U71 (.A1( u2_u2_X_12 ) , .A2( u2_u2_X_9 ) , .ZN( u2_u2_u1_n100 ) );
  NOR2_X1 u2_u2_u1_U72 (.A2( u2_u2_X_8 ) , .A1( u2_u2_u1_n177 ) , .ZN( u2_u2_u1_n99 ) );
  NOR2_X1 u2_u2_u1_U73 (.A2( u2_u2_X_12 ) , .ZN( u2_u2_u1_n102 ) , .A1( u2_u2_u1_n176 ) );
  NOR2_X1 u2_u2_u1_U74 (.A2( u2_u2_X_9 ) , .ZN( u2_u2_u1_n105 ) , .A1( u2_u2_u1_n168 ) );
  NAND2_X1 u2_u2_u1_U75 (.A1( u2_u2_X_10 ) , .ZN( u2_u2_u1_n160 ) , .A2( u2_u2_u1_n169 ) );
  NAND2_X1 u2_u2_u1_U76 (.A2( u2_u2_X_10 ) , .A1( u2_u2_X_11 ) , .ZN( u2_u2_u1_n152 ) );
  NAND2_X1 u2_u2_u1_U77 (.A1( u2_u2_X_11 ) , .ZN( u2_u2_u1_n128 ) , .A2( u2_u2_u1_n170 ) );
  AND2_X1 u2_u2_u1_U78 (.A2( u2_u2_X_7 ) , .A1( u2_u2_X_8 ) , .ZN( u2_u2_u1_n104 ) );
  AND2_X1 u2_u2_u1_U79 (.A1( u2_u2_X_8 ) , .ZN( u2_u2_u1_n103 ) , .A2( u2_u2_u1_n177 ) );
  AOI22_X1 u2_u2_u1_U8 (.B2( u2_u2_u1_n136 ) , .A2( u2_u2_u1_n137 ) , .ZN( u2_u2_u1_n143 ) , .A1( u2_u2_u1_n171 ) , .B1( u2_u2_u1_n173 ) );
  INV_X1 u2_u2_u1_U80 (.A( u2_u2_X_10 ) , .ZN( u2_u2_u1_n170 ) );
  INV_X1 u2_u2_u1_U81 (.A( u2_u2_X_9 ) , .ZN( u2_u2_u1_n176 ) );
  INV_X1 u2_u2_u1_U82 (.A( u2_u2_X_11 ) , .ZN( u2_u2_u1_n169 ) );
  INV_X1 u2_u2_u1_U83 (.A( u2_u2_X_12 ) , .ZN( u2_u2_u1_n168 ) );
  INV_X1 u2_u2_u1_U84 (.A( u2_u2_X_7 ) , .ZN( u2_u2_u1_n177 ) );
  NAND4_X1 u2_u2_u1_U85 (.ZN( u2_out2_28 ) , .A4( u2_u2_u1_n124 ) , .A3( u2_u2_u1_n125 ) , .A2( u2_u2_u1_n126 ) , .A1( u2_u2_u1_n127 ) );
  OAI21_X1 u2_u2_u1_U86 (.ZN( u2_u2_u1_n127 ) , .B2( u2_u2_u1_n139 ) , .B1( u2_u2_u1_n175 ) , .A( u2_u2_u1_n183 ) );
  OAI21_X1 u2_u2_u1_U87 (.ZN( u2_u2_u1_n126 ) , .B2( u2_u2_u1_n140 ) , .A( u2_u2_u1_n146 ) , .B1( u2_u2_u1_n178 ) );
  NAND4_X1 u2_u2_u1_U88 (.ZN( u2_out2_18 ) , .A4( u2_u2_u1_n165 ) , .A3( u2_u2_u1_n166 ) , .A1( u2_u2_u1_n167 ) , .A2( u2_u2_u1_n186 ) );
  AOI22_X1 u2_u2_u1_U89 (.B2( u2_u2_u1_n146 ) , .B1( u2_u2_u1_n147 ) , .A2( u2_u2_u1_n148 ) , .ZN( u2_u2_u1_n166 ) , .A1( u2_u2_u1_n172 ) );
  INV_X1 u2_u2_u1_U9 (.A( u2_u2_u1_n147 ) , .ZN( u2_u2_u1_n181 ) );
  INV_X1 u2_u2_u1_U90 (.A( u2_u2_u1_n145 ) , .ZN( u2_u2_u1_n186 ) );
  NAND4_X1 u2_u2_u1_U91 (.ZN( u2_out2_2 ) , .A4( u2_u2_u1_n142 ) , .A3( u2_u2_u1_n143 ) , .A2( u2_u2_u1_n144 ) , .A1( u2_u2_u1_n179 ) );
  OAI21_X1 u2_u2_u1_U92 (.B2( u2_u2_u1_n132 ) , .ZN( u2_u2_u1_n144 ) , .A( u2_u2_u1_n146 ) , .B1( u2_u2_u1_n180 ) );
  INV_X1 u2_u2_u1_U93 (.A( u2_u2_u1_n130 ) , .ZN( u2_u2_u1_n179 ) );
  OR4_X1 u2_u2_u1_U94 (.ZN( u2_out2_13 ) , .A4( u2_u2_u1_n108 ) , .A3( u2_u2_u1_n109 ) , .A2( u2_u2_u1_n110 ) , .A1( u2_u2_u1_n111 ) );
  AOI21_X1 u2_u2_u1_U95 (.ZN( u2_u2_u1_n111 ) , .A( u2_u2_u1_n128 ) , .B2( u2_u2_u1_n131 ) , .B1( u2_u2_u1_n135 ) );
  AOI21_X1 u2_u2_u1_U96 (.ZN( u2_u2_u1_n110 ) , .A( u2_u2_u1_n116 ) , .B1( u2_u2_u1_n152 ) , .B2( u2_u2_u1_n160 ) );
  NAND3_X1 u2_u2_u1_U97 (.A3( u2_u2_u1_n149 ) , .A2( u2_u2_u1_n150 ) , .A1( u2_u2_u1_n151 ) , .ZN( u2_u2_u1_n164 ) );
  NAND3_X1 u2_u2_u1_U98 (.A3( u2_u2_u1_n134 ) , .A2( u2_u2_u1_n135 ) , .ZN( u2_u2_u1_n136 ) , .A1( u2_u2_u1_n151 ) );
  NAND3_X1 u2_u2_u1_U99 (.A1( u2_u2_u1_n133 ) , .ZN( u2_u2_u1_n137 ) , .A2( u2_u2_u1_n154 ) , .A3( u2_u2_u1_n181 ) );
  OAI22_X1 u2_u2_u2_U10 (.B1( u2_u2_u2_n151 ) , .A2( u2_u2_u2_n152 ) , .A1( u2_u2_u2_n153 ) , .ZN( u2_u2_u2_n160 ) , .B2( u2_u2_u2_n168 ) );
  NAND3_X1 u2_u2_u2_U100 (.A2( u2_u2_u2_n100 ) , .A1( u2_u2_u2_n104 ) , .A3( u2_u2_u2_n138 ) , .ZN( u2_u2_u2_n98 ) );
  NOR3_X1 u2_u2_u2_U11 (.A1( u2_u2_u2_n150 ) , .ZN( u2_u2_u2_n151 ) , .A3( u2_u2_u2_n175 ) , .A2( u2_u2_u2_n188 ) );
  AOI21_X1 u2_u2_u2_U12 (.B2( u2_u2_u2_n123 ) , .ZN( u2_u2_u2_n125 ) , .A( u2_u2_u2_n171 ) , .B1( u2_u2_u2_n184 ) );
  INV_X1 u2_u2_u2_U13 (.A( u2_u2_u2_n150 ) , .ZN( u2_u2_u2_n184 ) );
  AOI21_X1 u2_u2_u2_U14 (.ZN( u2_u2_u2_n144 ) , .B2( u2_u2_u2_n155 ) , .A( u2_u2_u2_n172 ) , .B1( u2_u2_u2_n185 ) );
  AOI21_X1 u2_u2_u2_U15 (.B2( u2_u2_u2_n143 ) , .ZN( u2_u2_u2_n145 ) , .B1( u2_u2_u2_n152 ) , .A( u2_u2_u2_n171 ) );
  INV_X1 u2_u2_u2_U16 (.A( u2_u2_u2_n156 ) , .ZN( u2_u2_u2_n171 ) );
  INV_X1 u2_u2_u2_U17 (.A( u2_u2_u2_n120 ) , .ZN( u2_u2_u2_n188 ) );
  NAND2_X1 u2_u2_u2_U18 (.A2( u2_u2_u2_n122 ) , .ZN( u2_u2_u2_n150 ) , .A1( u2_u2_u2_n152 ) );
  INV_X1 u2_u2_u2_U19 (.A( u2_u2_u2_n153 ) , .ZN( u2_u2_u2_n170 ) );
  INV_X1 u2_u2_u2_U20 (.A( u2_u2_u2_n137 ) , .ZN( u2_u2_u2_n173 ) );
  NAND2_X1 u2_u2_u2_U21 (.A1( u2_u2_u2_n132 ) , .A2( u2_u2_u2_n139 ) , .ZN( u2_u2_u2_n157 ) );
  INV_X1 u2_u2_u2_U22 (.A( u2_u2_u2_n113 ) , .ZN( u2_u2_u2_n178 ) );
  INV_X1 u2_u2_u2_U23 (.A( u2_u2_u2_n139 ) , .ZN( u2_u2_u2_n175 ) );
  INV_X1 u2_u2_u2_U24 (.A( u2_u2_u2_n155 ) , .ZN( u2_u2_u2_n181 ) );
  INV_X1 u2_u2_u2_U25 (.A( u2_u2_u2_n119 ) , .ZN( u2_u2_u2_n177 ) );
  INV_X1 u2_u2_u2_U26 (.A( u2_u2_u2_n116 ) , .ZN( u2_u2_u2_n180 ) );
  INV_X1 u2_u2_u2_U27 (.A( u2_u2_u2_n131 ) , .ZN( u2_u2_u2_n179 ) );
  INV_X1 u2_u2_u2_U28 (.A( u2_u2_u2_n154 ) , .ZN( u2_u2_u2_n176 ) );
  NAND2_X1 u2_u2_u2_U29 (.A2( u2_u2_u2_n116 ) , .A1( u2_u2_u2_n117 ) , .ZN( u2_u2_u2_n118 ) );
  NOR2_X1 u2_u2_u2_U3 (.ZN( u2_u2_u2_n121 ) , .A2( u2_u2_u2_n177 ) , .A1( u2_u2_u2_n180 ) );
  INV_X1 u2_u2_u2_U30 (.A( u2_u2_u2_n132 ) , .ZN( u2_u2_u2_n182 ) );
  INV_X1 u2_u2_u2_U31 (.A( u2_u2_u2_n158 ) , .ZN( u2_u2_u2_n183 ) );
  OAI21_X1 u2_u2_u2_U32 (.A( u2_u2_u2_n156 ) , .B1( u2_u2_u2_n157 ) , .ZN( u2_u2_u2_n158 ) , .B2( u2_u2_u2_n179 ) );
  NOR2_X1 u2_u2_u2_U33 (.ZN( u2_u2_u2_n156 ) , .A1( u2_u2_u2_n166 ) , .A2( u2_u2_u2_n169 ) );
  NOR2_X1 u2_u2_u2_U34 (.A2( u2_u2_u2_n114 ) , .ZN( u2_u2_u2_n137 ) , .A1( u2_u2_u2_n140 ) );
  NOR2_X1 u2_u2_u2_U35 (.A2( u2_u2_u2_n138 ) , .ZN( u2_u2_u2_n153 ) , .A1( u2_u2_u2_n156 ) );
  AOI211_X1 u2_u2_u2_U36 (.ZN( u2_u2_u2_n130 ) , .C1( u2_u2_u2_n138 ) , .C2( u2_u2_u2_n179 ) , .B( u2_u2_u2_n96 ) , .A( u2_u2_u2_n97 ) );
  OAI22_X1 u2_u2_u2_U37 (.B1( u2_u2_u2_n133 ) , .A2( u2_u2_u2_n137 ) , .A1( u2_u2_u2_n152 ) , .B2( u2_u2_u2_n168 ) , .ZN( u2_u2_u2_n97 ) );
  OAI221_X1 u2_u2_u2_U38 (.B1( u2_u2_u2_n113 ) , .C1( u2_u2_u2_n132 ) , .A( u2_u2_u2_n149 ) , .B2( u2_u2_u2_n171 ) , .C2( u2_u2_u2_n172 ) , .ZN( u2_u2_u2_n96 ) );
  OAI221_X1 u2_u2_u2_U39 (.A( u2_u2_u2_n115 ) , .C2( u2_u2_u2_n123 ) , .B2( u2_u2_u2_n143 ) , .B1( u2_u2_u2_n153 ) , .ZN( u2_u2_u2_n163 ) , .C1( u2_u2_u2_n168 ) );
  INV_X1 u2_u2_u2_U4 (.A( u2_u2_u2_n134 ) , .ZN( u2_u2_u2_n185 ) );
  OAI21_X1 u2_u2_u2_U40 (.A( u2_u2_u2_n114 ) , .ZN( u2_u2_u2_n115 ) , .B1( u2_u2_u2_n176 ) , .B2( u2_u2_u2_n178 ) );
  OAI221_X1 u2_u2_u2_U41 (.A( u2_u2_u2_n135 ) , .B2( u2_u2_u2_n136 ) , .B1( u2_u2_u2_n137 ) , .ZN( u2_u2_u2_n162 ) , .C2( u2_u2_u2_n167 ) , .C1( u2_u2_u2_n185 ) );
  AND3_X1 u2_u2_u2_U42 (.A3( u2_u2_u2_n131 ) , .A2( u2_u2_u2_n132 ) , .A1( u2_u2_u2_n133 ) , .ZN( u2_u2_u2_n136 ) );
  AOI22_X1 u2_u2_u2_U43 (.ZN( u2_u2_u2_n135 ) , .B1( u2_u2_u2_n140 ) , .A1( u2_u2_u2_n156 ) , .B2( u2_u2_u2_n180 ) , .A2( u2_u2_u2_n188 ) );
  AOI21_X1 u2_u2_u2_U44 (.ZN( u2_u2_u2_n149 ) , .B1( u2_u2_u2_n173 ) , .B2( u2_u2_u2_n188 ) , .A( u2_u2_u2_n95 ) );
  AND3_X1 u2_u2_u2_U45 (.A2( u2_u2_u2_n100 ) , .A1( u2_u2_u2_n104 ) , .A3( u2_u2_u2_n156 ) , .ZN( u2_u2_u2_n95 ) );
  OAI21_X1 u2_u2_u2_U46 (.A( u2_u2_u2_n141 ) , .B2( u2_u2_u2_n142 ) , .ZN( u2_u2_u2_n146 ) , .B1( u2_u2_u2_n153 ) );
  OAI21_X1 u2_u2_u2_U47 (.A( u2_u2_u2_n140 ) , .ZN( u2_u2_u2_n141 ) , .B1( u2_u2_u2_n176 ) , .B2( u2_u2_u2_n177 ) );
  NOR3_X1 u2_u2_u2_U48 (.ZN( u2_u2_u2_n142 ) , .A3( u2_u2_u2_n175 ) , .A2( u2_u2_u2_n178 ) , .A1( u2_u2_u2_n181 ) );
  OAI21_X1 u2_u2_u2_U49 (.A( u2_u2_u2_n101 ) , .B2( u2_u2_u2_n121 ) , .B1( u2_u2_u2_n153 ) , .ZN( u2_u2_u2_n164 ) );
  NOR4_X1 u2_u2_u2_U5 (.A4( u2_u2_u2_n124 ) , .A3( u2_u2_u2_n125 ) , .A2( u2_u2_u2_n126 ) , .A1( u2_u2_u2_n127 ) , .ZN( u2_u2_u2_n128 ) );
  NAND2_X1 u2_u2_u2_U50 (.A2( u2_u2_u2_n100 ) , .A1( u2_u2_u2_n107 ) , .ZN( u2_u2_u2_n155 ) );
  NAND2_X1 u2_u2_u2_U51 (.A2( u2_u2_u2_n105 ) , .A1( u2_u2_u2_n108 ) , .ZN( u2_u2_u2_n143 ) );
  NAND2_X1 u2_u2_u2_U52 (.A1( u2_u2_u2_n104 ) , .A2( u2_u2_u2_n106 ) , .ZN( u2_u2_u2_n152 ) );
  NAND2_X1 u2_u2_u2_U53 (.A1( u2_u2_u2_n100 ) , .A2( u2_u2_u2_n105 ) , .ZN( u2_u2_u2_n132 ) );
  INV_X1 u2_u2_u2_U54 (.A( u2_u2_u2_n140 ) , .ZN( u2_u2_u2_n168 ) );
  INV_X1 u2_u2_u2_U55 (.A( u2_u2_u2_n138 ) , .ZN( u2_u2_u2_n167 ) );
  INV_X1 u2_u2_u2_U56 (.ZN( u2_u2_u2_n187 ) , .A( u2_u2_u2_n99 ) );
  OAI21_X1 u2_u2_u2_U57 (.B1( u2_u2_u2_n137 ) , .B2( u2_u2_u2_n143 ) , .A( u2_u2_u2_n98 ) , .ZN( u2_u2_u2_n99 ) );
  NAND2_X1 u2_u2_u2_U58 (.A1( u2_u2_u2_n102 ) , .A2( u2_u2_u2_n106 ) , .ZN( u2_u2_u2_n113 ) );
  NAND2_X1 u2_u2_u2_U59 (.A1( u2_u2_u2_n106 ) , .A2( u2_u2_u2_n107 ) , .ZN( u2_u2_u2_n131 ) );
  AOI21_X1 u2_u2_u2_U6 (.B2( u2_u2_u2_n119 ) , .ZN( u2_u2_u2_n127 ) , .A( u2_u2_u2_n137 ) , .B1( u2_u2_u2_n155 ) );
  NAND2_X1 u2_u2_u2_U60 (.A1( u2_u2_u2_n103 ) , .A2( u2_u2_u2_n107 ) , .ZN( u2_u2_u2_n139 ) );
  NAND2_X1 u2_u2_u2_U61 (.A1( u2_u2_u2_n103 ) , .A2( u2_u2_u2_n105 ) , .ZN( u2_u2_u2_n133 ) );
  NAND2_X1 u2_u2_u2_U62 (.A1( u2_u2_u2_n102 ) , .A2( u2_u2_u2_n103 ) , .ZN( u2_u2_u2_n154 ) );
  NAND2_X1 u2_u2_u2_U63 (.A2( u2_u2_u2_n103 ) , .A1( u2_u2_u2_n104 ) , .ZN( u2_u2_u2_n119 ) );
  NAND2_X1 u2_u2_u2_U64 (.A2( u2_u2_u2_n107 ) , .A1( u2_u2_u2_n108 ) , .ZN( u2_u2_u2_n123 ) );
  NAND2_X1 u2_u2_u2_U65 (.A1( u2_u2_u2_n104 ) , .A2( u2_u2_u2_n108 ) , .ZN( u2_u2_u2_n122 ) );
  INV_X1 u2_u2_u2_U66 (.A( u2_u2_u2_n114 ) , .ZN( u2_u2_u2_n172 ) );
  NAND2_X1 u2_u2_u2_U67 (.A2( u2_u2_u2_n100 ) , .A1( u2_u2_u2_n102 ) , .ZN( u2_u2_u2_n116 ) );
  NAND2_X1 u2_u2_u2_U68 (.A1( u2_u2_u2_n102 ) , .A2( u2_u2_u2_n108 ) , .ZN( u2_u2_u2_n120 ) );
  NAND2_X1 u2_u2_u2_U69 (.A2( u2_u2_u2_n105 ) , .A1( u2_u2_u2_n106 ) , .ZN( u2_u2_u2_n117 ) );
  AOI21_X1 u2_u2_u2_U7 (.ZN( u2_u2_u2_n124 ) , .B1( u2_u2_u2_n131 ) , .B2( u2_u2_u2_n143 ) , .A( u2_u2_u2_n172 ) );
  NOR2_X1 u2_u2_u2_U70 (.A2( u2_u2_X_16 ) , .ZN( u2_u2_u2_n140 ) , .A1( u2_u2_u2_n166 ) );
  NOR2_X1 u2_u2_u2_U71 (.A2( u2_u2_X_13 ) , .A1( u2_u2_X_14 ) , .ZN( u2_u2_u2_n100 ) );
  NOR2_X1 u2_u2_u2_U72 (.A2( u2_u2_X_16 ) , .A1( u2_u2_X_17 ) , .ZN( u2_u2_u2_n138 ) );
  NOR2_X1 u2_u2_u2_U73 (.A2( u2_u2_X_15 ) , .A1( u2_u2_X_18 ) , .ZN( u2_u2_u2_n104 ) );
  NOR2_X1 u2_u2_u2_U74 (.A2( u2_u2_X_14 ) , .ZN( u2_u2_u2_n103 ) , .A1( u2_u2_u2_n174 ) );
  NOR2_X1 u2_u2_u2_U75 (.A2( u2_u2_X_15 ) , .ZN( u2_u2_u2_n102 ) , .A1( u2_u2_u2_n165 ) );
  NOR2_X1 u2_u2_u2_U76 (.A2( u2_u2_X_17 ) , .ZN( u2_u2_u2_n114 ) , .A1( u2_u2_u2_n169 ) );
  AND2_X1 u2_u2_u2_U77 (.A1( u2_u2_X_15 ) , .ZN( u2_u2_u2_n105 ) , .A2( u2_u2_u2_n165 ) );
  AND2_X1 u2_u2_u2_U78 (.A2( u2_u2_X_15 ) , .A1( u2_u2_X_18 ) , .ZN( u2_u2_u2_n107 ) );
  AND2_X1 u2_u2_u2_U79 (.A1( u2_u2_X_14 ) , .ZN( u2_u2_u2_n106 ) , .A2( u2_u2_u2_n174 ) );
  AOI21_X1 u2_u2_u2_U8 (.B2( u2_u2_u2_n120 ) , .B1( u2_u2_u2_n121 ) , .ZN( u2_u2_u2_n126 ) , .A( u2_u2_u2_n167 ) );
  AND2_X1 u2_u2_u2_U80 (.A1( u2_u2_X_13 ) , .A2( u2_u2_X_14 ) , .ZN( u2_u2_u2_n108 ) );
  INV_X1 u2_u2_u2_U81 (.A( u2_u2_X_16 ) , .ZN( u2_u2_u2_n169 ) );
  INV_X1 u2_u2_u2_U82 (.A( u2_u2_X_17 ) , .ZN( u2_u2_u2_n166 ) );
  INV_X1 u2_u2_u2_U83 (.A( u2_u2_X_13 ) , .ZN( u2_u2_u2_n174 ) );
  INV_X1 u2_u2_u2_U84 (.A( u2_u2_X_18 ) , .ZN( u2_u2_u2_n165 ) );
  NAND4_X1 u2_u2_u2_U85 (.ZN( u2_out2_24 ) , .A4( u2_u2_u2_n111 ) , .A3( u2_u2_u2_n112 ) , .A1( u2_u2_u2_n130 ) , .A2( u2_u2_u2_n187 ) );
  AOI21_X1 u2_u2_u2_U86 (.ZN( u2_u2_u2_n112 ) , .B2( u2_u2_u2_n156 ) , .A( u2_u2_u2_n164 ) , .B1( u2_u2_u2_n181 ) );
  AOI221_X1 u2_u2_u2_U87 (.A( u2_u2_u2_n109 ) , .B1( u2_u2_u2_n110 ) , .ZN( u2_u2_u2_n111 ) , .C1( u2_u2_u2_n134 ) , .C2( u2_u2_u2_n170 ) , .B2( u2_u2_u2_n173 ) );
  NAND4_X1 u2_u2_u2_U88 (.ZN( u2_out2_16 ) , .A4( u2_u2_u2_n128 ) , .A3( u2_u2_u2_n129 ) , .A1( u2_u2_u2_n130 ) , .A2( u2_u2_u2_n186 ) );
  AOI22_X1 u2_u2_u2_U89 (.A2( u2_u2_u2_n118 ) , .ZN( u2_u2_u2_n129 ) , .A1( u2_u2_u2_n140 ) , .B1( u2_u2_u2_n157 ) , .B2( u2_u2_u2_n170 ) );
  OAI22_X1 u2_u2_u2_U9 (.ZN( u2_u2_u2_n109 ) , .A2( u2_u2_u2_n113 ) , .B2( u2_u2_u2_n133 ) , .B1( u2_u2_u2_n167 ) , .A1( u2_u2_u2_n168 ) );
  INV_X1 u2_u2_u2_U90 (.A( u2_u2_u2_n163 ) , .ZN( u2_u2_u2_n186 ) );
  NAND4_X1 u2_u2_u2_U91 (.ZN( u2_out2_30 ) , .A4( u2_u2_u2_n147 ) , .A3( u2_u2_u2_n148 ) , .A2( u2_u2_u2_n149 ) , .A1( u2_u2_u2_n187 ) );
  NOR3_X1 u2_u2_u2_U92 (.A3( u2_u2_u2_n144 ) , .A2( u2_u2_u2_n145 ) , .A1( u2_u2_u2_n146 ) , .ZN( u2_u2_u2_n147 ) );
  AOI21_X1 u2_u2_u2_U93 (.B2( u2_u2_u2_n138 ) , .ZN( u2_u2_u2_n148 ) , .A( u2_u2_u2_n162 ) , .B1( u2_u2_u2_n182 ) );
  OR4_X1 u2_u2_u2_U94 (.ZN( u2_out2_6 ) , .A4( u2_u2_u2_n161 ) , .A3( u2_u2_u2_n162 ) , .A2( u2_u2_u2_n163 ) , .A1( u2_u2_u2_n164 ) );
  OR3_X1 u2_u2_u2_U95 (.A2( u2_u2_u2_n159 ) , .A1( u2_u2_u2_n160 ) , .ZN( u2_u2_u2_n161 ) , .A3( u2_u2_u2_n183 ) );
  AOI21_X1 u2_u2_u2_U96 (.B2( u2_u2_u2_n154 ) , .B1( u2_u2_u2_n155 ) , .ZN( u2_u2_u2_n159 ) , .A( u2_u2_u2_n167 ) );
  NAND3_X1 u2_u2_u2_U97 (.A2( u2_u2_u2_n117 ) , .A1( u2_u2_u2_n122 ) , .A3( u2_u2_u2_n123 ) , .ZN( u2_u2_u2_n134 ) );
  NAND3_X1 u2_u2_u2_U98 (.ZN( u2_u2_u2_n110 ) , .A2( u2_u2_u2_n131 ) , .A3( u2_u2_u2_n139 ) , .A1( u2_u2_u2_n154 ) );
  NAND3_X1 u2_u2_u2_U99 (.A2( u2_u2_u2_n100 ) , .ZN( u2_u2_u2_n101 ) , .A1( u2_u2_u2_n104 ) , .A3( u2_u2_u2_n114 ) );
  OAI22_X1 u2_u2_u3_U10 (.B1( u2_u2_u3_n113 ) , .A2( u2_u2_u3_n135 ) , .A1( u2_u2_u3_n150 ) , .B2( u2_u2_u3_n164 ) , .ZN( u2_u2_u3_n98 ) );
  OAI211_X1 u2_u2_u3_U11 (.B( u2_u2_u3_n106 ) , .ZN( u2_u2_u3_n119 ) , .C2( u2_u2_u3_n128 ) , .C1( u2_u2_u3_n167 ) , .A( u2_u2_u3_n181 ) );
  AOI221_X1 u2_u2_u3_U12 (.C1( u2_u2_u3_n105 ) , .ZN( u2_u2_u3_n106 ) , .A( u2_u2_u3_n131 ) , .B2( u2_u2_u3_n132 ) , .C2( u2_u2_u3_n133 ) , .B1( u2_u2_u3_n169 ) );
  INV_X1 u2_u2_u3_U13 (.ZN( u2_u2_u3_n181 ) , .A( u2_u2_u3_n98 ) );
  NAND2_X1 u2_u2_u3_U14 (.ZN( u2_u2_u3_n105 ) , .A2( u2_u2_u3_n130 ) , .A1( u2_u2_u3_n155 ) );
  AOI22_X1 u2_u2_u3_U15 (.B1( u2_u2_u3_n115 ) , .A2( u2_u2_u3_n116 ) , .ZN( u2_u2_u3_n123 ) , .B2( u2_u2_u3_n133 ) , .A1( u2_u2_u3_n169 ) );
  NAND2_X1 u2_u2_u3_U16 (.ZN( u2_u2_u3_n116 ) , .A2( u2_u2_u3_n151 ) , .A1( u2_u2_u3_n182 ) );
  NOR2_X1 u2_u2_u3_U17 (.ZN( u2_u2_u3_n126 ) , .A2( u2_u2_u3_n150 ) , .A1( u2_u2_u3_n164 ) );
  AOI21_X1 u2_u2_u3_U18 (.ZN( u2_u2_u3_n112 ) , .B2( u2_u2_u3_n146 ) , .B1( u2_u2_u3_n155 ) , .A( u2_u2_u3_n167 ) );
  NAND2_X1 u2_u2_u3_U19 (.A1( u2_u2_u3_n135 ) , .ZN( u2_u2_u3_n142 ) , .A2( u2_u2_u3_n164 ) );
  NAND2_X1 u2_u2_u3_U20 (.ZN( u2_u2_u3_n132 ) , .A2( u2_u2_u3_n152 ) , .A1( u2_u2_u3_n156 ) );
  AND2_X1 u2_u2_u3_U21 (.A2( u2_u2_u3_n113 ) , .A1( u2_u2_u3_n114 ) , .ZN( u2_u2_u3_n151 ) );
  INV_X1 u2_u2_u3_U22 (.A( u2_u2_u3_n133 ) , .ZN( u2_u2_u3_n165 ) );
  INV_X1 u2_u2_u3_U23 (.A( u2_u2_u3_n135 ) , .ZN( u2_u2_u3_n170 ) );
  NAND2_X1 u2_u2_u3_U24 (.A1( u2_u2_u3_n107 ) , .A2( u2_u2_u3_n108 ) , .ZN( u2_u2_u3_n140 ) );
  NAND2_X1 u2_u2_u3_U25 (.ZN( u2_u2_u3_n117 ) , .A1( u2_u2_u3_n124 ) , .A2( u2_u2_u3_n148 ) );
  NAND2_X1 u2_u2_u3_U26 (.ZN( u2_u2_u3_n143 ) , .A1( u2_u2_u3_n165 ) , .A2( u2_u2_u3_n167 ) );
  INV_X1 u2_u2_u3_U27 (.A( u2_u2_u3_n130 ) , .ZN( u2_u2_u3_n177 ) );
  INV_X1 u2_u2_u3_U28 (.A( u2_u2_u3_n128 ) , .ZN( u2_u2_u3_n176 ) );
  INV_X1 u2_u2_u3_U29 (.A( u2_u2_u3_n155 ) , .ZN( u2_u2_u3_n174 ) );
  INV_X1 u2_u2_u3_U3 (.A( u2_u2_u3_n129 ) , .ZN( u2_u2_u3_n183 ) );
  INV_X1 u2_u2_u3_U30 (.A( u2_u2_u3_n139 ) , .ZN( u2_u2_u3_n185 ) );
  NOR2_X1 u2_u2_u3_U31 (.ZN( u2_u2_u3_n135 ) , .A2( u2_u2_u3_n141 ) , .A1( u2_u2_u3_n169 ) );
  OAI222_X1 u2_u2_u3_U32 (.C2( u2_u2_u3_n107 ) , .A2( u2_u2_u3_n108 ) , .B1( u2_u2_u3_n135 ) , .ZN( u2_u2_u3_n138 ) , .B2( u2_u2_u3_n146 ) , .C1( u2_u2_u3_n154 ) , .A1( u2_u2_u3_n164 ) );
  NOR4_X1 u2_u2_u3_U33 (.A4( u2_u2_u3_n157 ) , .A3( u2_u2_u3_n158 ) , .A2( u2_u2_u3_n159 ) , .A1( u2_u2_u3_n160 ) , .ZN( u2_u2_u3_n161 ) );
  AOI21_X1 u2_u2_u3_U34 (.B2( u2_u2_u3_n152 ) , .B1( u2_u2_u3_n153 ) , .ZN( u2_u2_u3_n158 ) , .A( u2_u2_u3_n164 ) );
  AOI21_X1 u2_u2_u3_U35 (.A( u2_u2_u3_n154 ) , .B2( u2_u2_u3_n155 ) , .B1( u2_u2_u3_n156 ) , .ZN( u2_u2_u3_n157 ) );
  AOI21_X1 u2_u2_u3_U36 (.A( u2_u2_u3_n149 ) , .B2( u2_u2_u3_n150 ) , .B1( u2_u2_u3_n151 ) , .ZN( u2_u2_u3_n159 ) );
  AOI211_X1 u2_u2_u3_U37 (.ZN( u2_u2_u3_n109 ) , .A( u2_u2_u3_n119 ) , .C2( u2_u2_u3_n129 ) , .B( u2_u2_u3_n138 ) , .C1( u2_u2_u3_n141 ) );
  AOI211_X1 u2_u2_u3_U38 (.B( u2_u2_u3_n119 ) , .A( u2_u2_u3_n120 ) , .C2( u2_u2_u3_n121 ) , .ZN( u2_u2_u3_n122 ) , .C1( u2_u2_u3_n179 ) );
  INV_X1 u2_u2_u3_U39 (.A( u2_u2_u3_n156 ) , .ZN( u2_u2_u3_n179 ) );
  INV_X1 u2_u2_u3_U4 (.A( u2_u2_u3_n140 ) , .ZN( u2_u2_u3_n182 ) );
  OAI22_X1 u2_u2_u3_U40 (.B1( u2_u2_u3_n118 ) , .ZN( u2_u2_u3_n120 ) , .A1( u2_u2_u3_n135 ) , .B2( u2_u2_u3_n154 ) , .A2( u2_u2_u3_n178 ) );
  AND3_X1 u2_u2_u3_U41 (.ZN( u2_u2_u3_n118 ) , .A2( u2_u2_u3_n124 ) , .A1( u2_u2_u3_n144 ) , .A3( u2_u2_u3_n152 ) );
  INV_X1 u2_u2_u3_U42 (.A( u2_u2_u3_n121 ) , .ZN( u2_u2_u3_n164 ) );
  NAND2_X1 u2_u2_u3_U43 (.ZN( u2_u2_u3_n133 ) , .A1( u2_u2_u3_n154 ) , .A2( u2_u2_u3_n164 ) );
  OAI211_X1 u2_u2_u3_U44 (.B( u2_u2_u3_n127 ) , .ZN( u2_u2_u3_n139 ) , .C1( u2_u2_u3_n150 ) , .C2( u2_u2_u3_n154 ) , .A( u2_u2_u3_n184 ) );
  INV_X1 u2_u2_u3_U45 (.A( u2_u2_u3_n125 ) , .ZN( u2_u2_u3_n184 ) );
  AOI221_X1 u2_u2_u3_U46 (.A( u2_u2_u3_n126 ) , .ZN( u2_u2_u3_n127 ) , .C2( u2_u2_u3_n132 ) , .C1( u2_u2_u3_n169 ) , .B2( u2_u2_u3_n170 ) , .B1( u2_u2_u3_n174 ) );
  OAI22_X1 u2_u2_u3_U47 (.A1( u2_u2_u3_n124 ) , .ZN( u2_u2_u3_n125 ) , .B2( u2_u2_u3_n145 ) , .A2( u2_u2_u3_n165 ) , .B1( u2_u2_u3_n167 ) );
  NOR2_X1 u2_u2_u3_U48 (.A1( u2_u2_u3_n113 ) , .ZN( u2_u2_u3_n131 ) , .A2( u2_u2_u3_n154 ) );
  NAND2_X1 u2_u2_u3_U49 (.A1( u2_u2_u3_n103 ) , .ZN( u2_u2_u3_n150 ) , .A2( u2_u2_u3_n99 ) );
  INV_X1 u2_u2_u3_U5 (.A( u2_u2_u3_n117 ) , .ZN( u2_u2_u3_n178 ) );
  NAND2_X1 u2_u2_u3_U50 (.A2( u2_u2_u3_n102 ) , .ZN( u2_u2_u3_n155 ) , .A1( u2_u2_u3_n97 ) );
  INV_X1 u2_u2_u3_U51 (.A( u2_u2_u3_n141 ) , .ZN( u2_u2_u3_n167 ) );
  AOI21_X1 u2_u2_u3_U52 (.B2( u2_u2_u3_n114 ) , .B1( u2_u2_u3_n146 ) , .A( u2_u2_u3_n154 ) , .ZN( u2_u2_u3_n94 ) );
  AOI21_X1 u2_u2_u3_U53 (.ZN( u2_u2_u3_n110 ) , .B2( u2_u2_u3_n142 ) , .B1( u2_u2_u3_n186 ) , .A( u2_u2_u3_n95 ) );
  INV_X1 u2_u2_u3_U54 (.A( u2_u2_u3_n145 ) , .ZN( u2_u2_u3_n186 ) );
  AOI21_X1 u2_u2_u3_U55 (.B1( u2_u2_u3_n124 ) , .A( u2_u2_u3_n149 ) , .B2( u2_u2_u3_n155 ) , .ZN( u2_u2_u3_n95 ) );
  INV_X1 u2_u2_u3_U56 (.A( u2_u2_u3_n149 ) , .ZN( u2_u2_u3_n169 ) );
  NAND2_X1 u2_u2_u3_U57 (.ZN( u2_u2_u3_n124 ) , .A1( u2_u2_u3_n96 ) , .A2( u2_u2_u3_n97 ) );
  NAND2_X1 u2_u2_u3_U58 (.A2( u2_u2_u3_n100 ) , .ZN( u2_u2_u3_n146 ) , .A1( u2_u2_u3_n96 ) );
  NAND2_X1 u2_u2_u3_U59 (.A1( u2_u2_u3_n101 ) , .ZN( u2_u2_u3_n145 ) , .A2( u2_u2_u3_n99 ) );
  AOI221_X1 u2_u2_u3_U6 (.A( u2_u2_u3_n131 ) , .C2( u2_u2_u3_n132 ) , .C1( u2_u2_u3_n133 ) , .ZN( u2_u2_u3_n134 ) , .B1( u2_u2_u3_n143 ) , .B2( u2_u2_u3_n177 ) );
  NAND2_X1 u2_u2_u3_U60 (.A1( u2_u2_u3_n100 ) , .ZN( u2_u2_u3_n156 ) , .A2( u2_u2_u3_n99 ) );
  NAND2_X1 u2_u2_u3_U61 (.A2( u2_u2_u3_n101 ) , .A1( u2_u2_u3_n104 ) , .ZN( u2_u2_u3_n148 ) );
  NAND2_X1 u2_u2_u3_U62 (.A1( u2_u2_u3_n100 ) , .A2( u2_u2_u3_n102 ) , .ZN( u2_u2_u3_n128 ) );
  NAND2_X1 u2_u2_u3_U63 (.A2( u2_u2_u3_n101 ) , .A1( u2_u2_u3_n102 ) , .ZN( u2_u2_u3_n152 ) );
  NAND2_X1 u2_u2_u3_U64 (.A2( u2_u2_u3_n101 ) , .ZN( u2_u2_u3_n114 ) , .A1( u2_u2_u3_n96 ) );
  NAND2_X1 u2_u2_u3_U65 (.ZN( u2_u2_u3_n107 ) , .A1( u2_u2_u3_n97 ) , .A2( u2_u2_u3_n99 ) );
  NAND2_X1 u2_u2_u3_U66 (.A2( u2_u2_u3_n100 ) , .A1( u2_u2_u3_n104 ) , .ZN( u2_u2_u3_n113 ) );
  NAND2_X1 u2_u2_u3_U67 (.A1( u2_u2_u3_n104 ) , .ZN( u2_u2_u3_n153 ) , .A2( u2_u2_u3_n97 ) );
  NAND2_X1 u2_u2_u3_U68 (.A2( u2_u2_u3_n103 ) , .A1( u2_u2_u3_n104 ) , .ZN( u2_u2_u3_n130 ) );
  NAND2_X1 u2_u2_u3_U69 (.A2( u2_u2_u3_n103 ) , .ZN( u2_u2_u3_n144 ) , .A1( u2_u2_u3_n96 ) );
  OAI22_X1 u2_u2_u3_U7 (.B2( u2_u2_u3_n147 ) , .A2( u2_u2_u3_n148 ) , .ZN( u2_u2_u3_n160 ) , .B1( u2_u2_u3_n165 ) , .A1( u2_u2_u3_n168 ) );
  NAND2_X1 u2_u2_u3_U70 (.A1( u2_u2_u3_n102 ) , .A2( u2_u2_u3_n103 ) , .ZN( u2_u2_u3_n108 ) );
  NOR2_X1 u2_u2_u3_U71 (.A2( u2_u2_X_19 ) , .A1( u2_u2_X_20 ) , .ZN( u2_u2_u3_n99 ) );
  NOR2_X1 u2_u2_u3_U72 (.A2( u2_u2_X_21 ) , .A1( u2_u2_X_24 ) , .ZN( u2_u2_u3_n103 ) );
  NOR2_X1 u2_u2_u3_U73 (.A2( u2_u2_X_24 ) , .A1( u2_u2_u3_n171 ) , .ZN( u2_u2_u3_n97 ) );
  NOR2_X1 u2_u2_u3_U74 (.A2( u2_u2_X_23 ) , .ZN( u2_u2_u3_n141 ) , .A1( u2_u2_u3_n166 ) );
  NOR2_X1 u2_u2_u3_U75 (.A2( u2_u2_X_19 ) , .A1( u2_u2_u3_n172 ) , .ZN( u2_u2_u3_n96 ) );
  NAND2_X1 u2_u2_u3_U76 (.A1( u2_u2_X_22 ) , .A2( u2_u2_X_23 ) , .ZN( u2_u2_u3_n154 ) );
  NAND2_X1 u2_u2_u3_U77 (.A1( u2_u2_X_23 ) , .ZN( u2_u2_u3_n149 ) , .A2( u2_u2_u3_n166 ) );
  NOR2_X1 u2_u2_u3_U78 (.A2( u2_u2_X_22 ) , .A1( u2_u2_X_23 ) , .ZN( u2_u2_u3_n121 ) );
  AND2_X1 u2_u2_u3_U79 (.A1( u2_u2_X_24 ) , .ZN( u2_u2_u3_n101 ) , .A2( u2_u2_u3_n171 ) );
  AND3_X1 u2_u2_u3_U8 (.A3( u2_u2_u3_n144 ) , .A2( u2_u2_u3_n145 ) , .A1( u2_u2_u3_n146 ) , .ZN( u2_u2_u3_n147 ) );
  AND2_X1 u2_u2_u3_U80 (.A1( u2_u2_X_19 ) , .ZN( u2_u2_u3_n102 ) , .A2( u2_u2_u3_n172 ) );
  AND2_X1 u2_u2_u3_U81 (.A1( u2_u2_X_21 ) , .A2( u2_u2_X_24 ) , .ZN( u2_u2_u3_n100 ) );
  AND2_X1 u2_u2_u3_U82 (.A2( u2_u2_X_19 ) , .A1( u2_u2_X_20 ) , .ZN( u2_u2_u3_n104 ) );
  INV_X1 u2_u2_u3_U83 (.A( u2_u2_X_22 ) , .ZN( u2_u2_u3_n166 ) );
  INV_X1 u2_u2_u3_U84 (.A( u2_u2_X_21 ) , .ZN( u2_u2_u3_n171 ) );
  INV_X1 u2_u2_u3_U85 (.A( u2_u2_X_20 ) , .ZN( u2_u2_u3_n172 ) );
  OR4_X1 u2_u2_u3_U86 (.ZN( u2_out2_10 ) , .A4( u2_u2_u3_n136 ) , .A3( u2_u2_u3_n137 ) , .A1( u2_u2_u3_n138 ) , .A2( u2_u2_u3_n139 ) );
  OAI222_X1 u2_u2_u3_U87 (.C1( u2_u2_u3_n128 ) , .ZN( u2_u2_u3_n137 ) , .B1( u2_u2_u3_n148 ) , .A2( u2_u2_u3_n150 ) , .B2( u2_u2_u3_n154 ) , .C2( u2_u2_u3_n164 ) , .A1( u2_u2_u3_n167 ) );
  OAI221_X1 u2_u2_u3_U88 (.A( u2_u2_u3_n134 ) , .B2( u2_u2_u3_n135 ) , .ZN( u2_u2_u3_n136 ) , .C1( u2_u2_u3_n149 ) , .B1( u2_u2_u3_n151 ) , .C2( u2_u2_u3_n183 ) );
  NAND4_X1 u2_u2_u3_U89 (.ZN( u2_out2_26 ) , .A4( u2_u2_u3_n109 ) , .A3( u2_u2_u3_n110 ) , .A2( u2_u2_u3_n111 ) , .A1( u2_u2_u3_n173 ) );
  INV_X1 u2_u2_u3_U9 (.A( u2_u2_u3_n143 ) , .ZN( u2_u2_u3_n168 ) );
  INV_X1 u2_u2_u3_U90 (.ZN( u2_u2_u3_n173 ) , .A( u2_u2_u3_n94 ) );
  OAI21_X1 u2_u2_u3_U91 (.ZN( u2_u2_u3_n111 ) , .B2( u2_u2_u3_n117 ) , .A( u2_u2_u3_n133 ) , .B1( u2_u2_u3_n176 ) );
  NAND4_X1 u2_u2_u3_U92 (.ZN( u2_out2_20 ) , .A4( u2_u2_u3_n122 ) , .A3( u2_u2_u3_n123 ) , .A1( u2_u2_u3_n175 ) , .A2( u2_u2_u3_n180 ) );
  INV_X1 u2_u2_u3_U93 (.A( u2_u2_u3_n112 ) , .ZN( u2_u2_u3_n175 ) );
  INV_X1 u2_u2_u3_U94 (.A( u2_u2_u3_n126 ) , .ZN( u2_u2_u3_n180 ) );
  NAND4_X1 u2_u2_u3_U95 (.ZN( u2_out2_1 ) , .A4( u2_u2_u3_n161 ) , .A3( u2_u2_u3_n162 ) , .A2( u2_u2_u3_n163 ) , .A1( u2_u2_u3_n185 ) );
  NAND2_X1 u2_u2_u3_U96 (.ZN( u2_u2_u3_n163 ) , .A2( u2_u2_u3_n170 ) , .A1( u2_u2_u3_n176 ) );
  AOI22_X1 u2_u2_u3_U97 (.B2( u2_u2_u3_n140 ) , .B1( u2_u2_u3_n141 ) , .A2( u2_u2_u3_n142 ) , .ZN( u2_u2_u3_n162 ) , .A1( u2_u2_u3_n177 ) );
  NAND3_X1 u2_u2_u3_U98 (.A1( u2_u2_u3_n114 ) , .ZN( u2_u2_u3_n115 ) , .A2( u2_u2_u3_n145 ) , .A3( u2_u2_u3_n153 ) );
  NAND3_X1 u2_u2_u3_U99 (.ZN( u2_u2_u3_n129 ) , .A2( u2_u2_u3_n144 ) , .A1( u2_u2_u3_n153 ) , .A3( u2_u2_u3_n182 ) );
  INV_X1 u2_u2_u5_U10 (.A( u2_u2_u5_n121 ) , .ZN( u2_u2_u5_n177 ) );
  NOR3_X1 u2_u2_u5_U100 (.A3( u2_u2_u5_n141 ) , .A1( u2_u2_u5_n142 ) , .ZN( u2_u2_u5_n143 ) , .A2( u2_u2_u5_n191 ) );
  NAND4_X1 u2_u2_u5_U101 (.ZN( u2_out2_4 ) , .A4( u2_u2_u5_n112 ) , .A2( u2_u2_u5_n113 ) , .A1( u2_u2_u5_n114 ) , .A3( u2_u2_u5_n195 ) );
  AOI211_X1 u2_u2_u5_U102 (.A( u2_u2_u5_n110 ) , .C1( u2_u2_u5_n111 ) , .ZN( u2_u2_u5_n112 ) , .B( u2_u2_u5_n118 ) , .C2( u2_u2_u5_n177 ) );
  AOI222_X1 u2_u2_u5_U103 (.ZN( u2_u2_u5_n113 ) , .A1( u2_u2_u5_n131 ) , .C1( u2_u2_u5_n148 ) , .B2( u2_u2_u5_n174 ) , .C2( u2_u2_u5_n178 ) , .A2( u2_u2_u5_n179 ) , .B1( u2_u2_u5_n99 ) );
  NAND3_X1 u2_u2_u5_U104 (.A2( u2_u2_u5_n154 ) , .A3( u2_u2_u5_n158 ) , .A1( u2_u2_u5_n161 ) , .ZN( u2_u2_u5_n99 ) );
  NOR2_X1 u2_u2_u5_U11 (.ZN( u2_u2_u5_n160 ) , .A2( u2_u2_u5_n173 ) , .A1( u2_u2_u5_n177 ) );
  INV_X1 u2_u2_u5_U12 (.A( u2_u2_u5_n150 ) , .ZN( u2_u2_u5_n174 ) );
  AOI21_X1 u2_u2_u5_U13 (.A( u2_u2_u5_n160 ) , .B2( u2_u2_u5_n161 ) , .ZN( u2_u2_u5_n162 ) , .B1( u2_u2_u5_n192 ) );
  INV_X1 u2_u2_u5_U14 (.A( u2_u2_u5_n159 ) , .ZN( u2_u2_u5_n192 ) );
  AOI21_X1 u2_u2_u5_U15 (.A( u2_u2_u5_n156 ) , .B2( u2_u2_u5_n157 ) , .B1( u2_u2_u5_n158 ) , .ZN( u2_u2_u5_n163 ) );
  AOI21_X1 u2_u2_u5_U16 (.B2( u2_u2_u5_n139 ) , .B1( u2_u2_u5_n140 ) , .ZN( u2_u2_u5_n141 ) , .A( u2_u2_u5_n150 ) );
  OAI21_X1 u2_u2_u5_U17 (.A( u2_u2_u5_n133 ) , .B2( u2_u2_u5_n134 ) , .B1( u2_u2_u5_n135 ) , .ZN( u2_u2_u5_n142 ) );
  OAI21_X1 u2_u2_u5_U18 (.ZN( u2_u2_u5_n133 ) , .B2( u2_u2_u5_n147 ) , .A( u2_u2_u5_n173 ) , .B1( u2_u2_u5_n188 ) );
  NAND2_X1 u2_u2_u5_U19 (.A2( u2_u2_u5_n119 ) , .A1( u2_u2_u5_n123 ) , .ZN( u2_u2_u5_n137 ) );
  INV_X1 u2_u2_u5_U20 (.A( u2_u2_u5_n155 ) , .ZN( u2_u2_u5_n194 ) );
  NAND2_X1 u2_u2_u5_U21 (.A1( u2_u2_u5_n121 ) , .ZN( u2_u2_u5_n132 ) , .A2( u2_u2_u5_n172 ) );
  NAND2_X1 u2_u2_u5_U22 (.A2( u2_u2_u5_n122 ) , .ZN( u2_u2_u5_n136 ) , .A1( u2_u2_u5_n154 ) );
  NAND2_X1 u2_u2_u5_U23 (.A2( u2_u2_u5_n119 ) , .A1( u2_u2_u5_n120 ) , .ZN( u2_u2_u5_n159 ) );
  INV_X1 u2_u2_u5_U24 (.A( u2_u2_u5_n156 ) , .ZN( u2_u2_u5_n175 ) );
  INV_X1 u2_u2_u5_U25 (.A( u2_u2_u5_n158 ) , .ZN( u2_u2_u5_n188 ) );
  INV_X1 u2_u2_u5_U26 (.A( u2_u2_u5_n152 ) , .ZN( u2_u2_u5_n179 ) );
  INV_X1 u2_u2_u5_U27 (.A( u2_u2_u5_n140 ) , .ZN( u2_u2_u5_n182 ) );
  INV_X1 u2_u2_u5_U28 (.A( u2_u2_u5_n151 ) , .ZN( u2_u2_u5_n183 ) );
  INV_X1 u2_u2_u5_U29 (.A( u2_u2_u5_n123 ) , .ZN( u2_u2_u5_n185 ) );
  NOR2_X1 u2_u2_u5_U3 (.ZN( u2_u2_u5_n134 ) , .A1( u2_u2_u5_n183 ) , .A2( u2_u2_u5_n190 ) );
  INV_X1 u2_u2_u5_U30 (.A( u2_u2_u5_n161 ) , .ZN( u2_u2_u5_n184 ) );
  INV_X1 u2_u2_u5_U31 (.A( u2_u2_u5_n139 ) , .ZN( u2_u2_u5_n189 ) );
  INV_X1 u2_u2_u5_U32 (.A( u2_u2_u5_n157 ) , .ZN( u2_u2_u5_n190 ) );
  INV_X1 u2_u2_u5_U33 (.A( u2_u2_u5_n120 ) , .ZN( u2_u2_u5_n193 ) );
  NAND2_X1 u2_u2_u5_U34 (.ZN( u2_u2_u5_n111 ) , .A1( u2_u2_u5_n140 ) , .A2( u2_u2_u5_n155 ) );
  INV_X1 u2_u2_u5_U35 (.A( u2_u2_u5_n117 ) , .ZN( u2_u2_u5_n196 ) );
  OAI221_X1 u2_u2_u5_U36 (.A( u2_u2_u5_n116 ) , .ZN( u2_u2_u5_n117 ) , .B2( u2_u2_u5_n119 ) , .C1( u2_u2_u5_n153 ) , .C2( u2_u2_u5_n158 ) , .B1( u2_u2_u5_n172 ) );
  AOI222_X1 u2_u2_u5_U37 (.ZN( u2_u2_u5_n116 ) , .B2( u2_u2_u5_n145 ) , .C1( u2_u2_u5_n148 ) , .A2( u2_u2_u5_n174 ) , .C2( u2_u2_u5_n177 ) , .B1( u2_u2_u5_n187 ) , .A1( u2_u2_u5_n193 ) );
  INV_X1 u2_u2_u5_U38 (.A( u2_u2_u5_n115 ) , .ZN( u2_u2_u5_n187 ) );
  NOR2_X1 u2_u2_u5_U39 (.ZN( u2_u2_u5_n100 ) , .A1( u2_u2_u5_n170 ) , .A2( u2_u2_u5_n180 ) );
  INV_X1 u2_u2_u5_U4 (.A( u2_u2_u5_n138 ) , .ZN( u2_u2_u5_n191 ) );
  AOI22_X1 u2_u2_u5_U40 (.B2( u2_u2_u5_n131 ) , .A2( u2_u2_u5_n146 ) , .ZN( u2_u2_u5_n169 ) , .B1( u2_u2_u5_n174 ) , .A1( u2_u2_u5_n185 ) );
  NOR2_X1 u2_u2_u5_U41 (.A1( u2_u2_u5_n146 ) , .ZN( u2_u2_u5_n150 ) , .A2( u2_u2_u5_n173 ) );
  AOI21_X1 u2_u2_u5_U42 (.A( u2_u2_u5_n118 ) , .B2( u2_u2_u5_n145 ) , .ZN( u2_u2_u5_n168 ) , .B1( u2_u2_u5_n186 ) );
  INV_X1 u2_u2_u5_U43 (.A( u2_u2_u5_n122 ) , .ZN( u2_u2_u5_n186 ) );
  NOR2_X1 u2_u2_u5_U44 (.A1( u2_u2_u5_n146 ) , .ZN( u2_u2_u5_n152 ) , .A2( u2_u2_u5_n176 ) );
  NOR2_X1 u2_u2_u5_U45 (.A1( u2_u2_u5_n115 ) , .ZN( u2_u2_u5_n118 ) , .A2( u2_u2_u5_n153 ) );
  NOR2_X1 u2_u2_u5_U46 (.A2( u2_u2_u5_n145 ) , .ZN( u2_u2_u5_n156 ) , .A1( u2_u2_u5_n174 ) );
  NOR2_X1 u2_u2_u5_U47 (.ZN( u2_u2_u5_n121 ) , .A2( u2_u2_u5_n145 ) , .A1( u2_u2_u5_n176 ) );
  AOI22_X1 u2_u2_u5_U48 (.ZN( u2_u2_u5_n114 ) , .A2( u2_u2_u5_n137 ) , .A1( u2_u2_u5_n145 ) , .B2( u2_u2_u5_n175 ) , .B1( u2_u2_u5_n193 ) );
  AOI21_X1 u2_u2_u5_U49 (.A( u2_u2_u5_n153 ) , .B2( u2_u2_u5_n154 ) , .B1( u2_u2_u5_n155 ) , .ZN( u2_u2_u5_n164 ) );
  OAI21_X1 u2_u2_u5_U5 (.B2( u2_u2_u5_n136 ) , .B1( u2_u2_u5_n137 ) , .ZN( u2_u2_u5_n138 ) , .A( u2_u2_u5_n177 ) );
  AOI21_X1 u2_u2_u5_U50 (.ZN( u2_u2_u5_n110 ) , .B1( u2_u2_u5_n122 ) , .B2( u2_u2_u5_n139 ) , .A( u2_u2_u5_n153 ) );
  INV_X1 u2_u2_u5_U51 (.A( u2_u2_u5_n153 ) , .ZN( u2_u2_u5_n176 ) );
  INV_X1 u2_u2_u5_U52 (.A( u2_u2_u5_n126 ) , .ZN( u2_u2_u5_n173 ) );
  AND2_X1 u2_u2_u5_U53 (.A2( u2_u2_u5_n104 ) , .A1( u2_u2_u5_n107 ) , .ZN( u2_u2_u5_n147 ) );
  AND2_X1 u2_u2_u5_U54 (.A2( u2_u2_u5_n104 ) , .A1( u2_u2_u5_n108 ) , .ZN( u2_u2_u5_n148 ) );
  NAND2_X1 u2_u2_u5_U55 (.A1( u2_u2_u5_n105 ) , .A2( u2_u2_u5_n106 ) , .ZN( u2_u2_u5_n158 ) );
  NAND2_X1 u2_u2_u5_U56 (.A2( u2_u2_u5_n108 ) , .A1( u2_u2_u5_n109 ) , .ZN( u2_u2_u5_n139 ) );
  NAND2_X1 u2_u2_u5_U57 (.A1( u2_u2_u5_n106 ) , .A2( u2_u2_u5_n108 ) , .ZN( u2_u2_u5_n119 ) );
  OAI211_X1 u2_u2_u5_U58 (.B( u2_u2_u5_n124 ) , .A( u2_u2_u5_n125 ) , .C2( u2_u2_u5_n126 ) , .C1( u2_u2_u5_n127 ) , .ZN( u2_u2_u5_n128 ) );
  NOR3_X1 u2_u2_u5_U59 (.ZN( u2_u2_u5_n127 ) , .A1( u2_u2_u5_n136 ) , .A3( u2_u2_u5_n148 ) , .A2( u2_u2_u5_n182 ) );
  INV_X1 u2_u2_u5_U6 (.A( u2_u2_u5_n135 ) , .ZN( u2_u2_u5_n178 ) );
  OAI21_X1 u2_u2_u5_U60 (.ZN( u2_u2_u5_n124 ) , .A( u2_u2_u5_n177 ) , .B2( u2_u2_u5_n183 ) , .B1( u2_u2_u5_n189 ) );
  OAI21_X1 u2_u2_u5_U61 (.ZN( u2_u2_u5_n125 ) , .A( u2_u2_u5_n174 ) , .B2( u2_u2_u5_n185 ) , .B1( u2_u2_u5_n190 ) );
  NAND2_X1 u2_u2_u5_U62 (.A2( u2_u2_u5_n103 ) , .A1( u2_u2_u5_n105 ) , .ZN( u2_u2_u5_n140 ) );
  NAND2_X1 u2_u2_u5_U63 (.A2( u2_u2_u5_n104 ) , .A1( u2_u2_u5_n105 ) , .ZN( u2_u2_u5_n155 ) );
  NAND2_X1 u2_u2_u5_U64 (.A2( u2_u2_u5_n106 ) , .A1( u2_u2_u5_n107 ) , .ZN( u2_u2_u5_n122 ) );
  NAND2_X1 u2_u2_u5_U65 (.A2( u2_u2_u5_n100 ) , .A1( u2_u2_u5_n106 ) , .ZN( u2_u2_u5_n115 ) );
  NAND2_X1 u2_u2_u5_U66 (.A2( u2_u2_u5_n100 ) , .A1( u2_u2_u5_n103 ) , .ZN( u2_u2_u5_n161 ) );
  NAND2_X1 u2_u2_u5_U67 (.A1( u2_u2_u5_n105 ) , .A2( u2_u2_u5_n109 ) , .ZN( u2_u2_u5_n154 ) );
  INV_X1 u2_u2_u5_U68 (.A( u2_u2_u5_n146 ) , .ZN( u2_u2_u5_n172 ) );
  NAND2_X1 u2_u2_u5_U69 (.A1( u2_u2_u5_n103 ) , .A2( u2_u2_u5_n108 ) , .ZN( u2_u2_u5_n123 ) );
  OAI22_X1 u2_u2_u5_U7 (.B2( u2_u2_u5_n149 ) , .B1( u2_u2_u5_n150 ) , .A2( u2_u2_u5_n151 ) , .A1( u2_u2_u5_n152 ) , .ZN( u2_u2_u5_n165 ) );
  NAND2_X1 u2_u2_u5_U70 (.A2( u2_u2_u5_n103 ) , .A1( u2_u2_u5_n107 ) , .ZN( u2_u2_u5_n151 ) );
  NAND2_X1 u2_u2_u5_U71 (.A2( u2_u2_u5_n107 ) , .A1( u2_u2_u5_n109 ) , .ZN( u2_u2_u5_n120 ) );
  NAND2_X1 u2_u2_u5_U72 (.A2( u2_u2_u5_n100 ) , .A1( u2_u2_u5_n109 ) , .ZN( u2_u2_u5_n157 ) );
  AND2_X1 u2_u2_u5_U73 (.A2( u2_u2_u5_n100 ) , .A1( u2_u2_u5_n104 ) , .ZN( u2_u2_u5_n131 ) );
  INV_X1 u2_u2_u5_U74 (.A( u2_u2_u5_n102 ) , .ZN( u2_u2_u5_n195 ) );
  OAI221_X1 u2_u2_u5_U75 (.A( u2_u2_u5_n101 ) , .ZN( u2_u2_u5_n102 ) , .C2( u2_u2_u5_n115 ) , .C1( u2_u2_u5_n126 ) , .B1( u2_u2_u5_n134 ) , .B2( u2_u2_u5_n160 ) );
  OAI21_X1 u2_u2_u5_U76 (.ZN( u2_u2_u5_n101 ) , .B1( u2_u2_u5_n137 ) , .A( u2_u2_u5_n146 ) , .B2( u2_u2_u5_n147 ) );
  NOR2_X1 u2_u2_u5_U77 (.A2( u2_u2_X_34 ) , .A1( u2_u2_X_35 ) , .ZN( u2_u2_u5_n145 ) );
  NOR2_X1 u2_u2_u5_U78 (.A2( u2_u2_X_34 ) , .ZN( u2_u2_u5_n146 ) , .A1( u2_u2_u5_n171 ) );
  NOR2_X1 u2_u2_u5_U79 (.A2( u2_u2_X_31 ) , .A1( u2_u2_X_32 ) , .ZN( u2_u2_u5_n103 ) );
  NOR3_X1 u2_u2_u5_U8 (.A2( u2_u2_u5_n147 ) , .A1( u2_u2_u5_n148 ) , .ZN( u2_u2_u5_n149 ) , .A3( u2_u2_u5_n194 ) );
  NOR2_X1 u2_u2_u5_U80 (.A2( u2_u2_X_36 ) , .ZN( u2_u2_u5_n105 ) , .A1( u2_u2_u5_n180 ) );
  NOR2_X1 u2_u2_u5_U81 (.A2( u2_u2_X_33 ) , .ZN( u2_u2_u5_n108 ) , .A1( u2_u2_u5_n170 ) );
  NOR2_X1 u2_u2_u5_U82 (.A2( u2_u2_X_33 ) , .A1( u2_u2_X_36 ) , .ZN( u2_u2_u5_n107 ) );
  NOR2_X1 u2_u2_u5_U83 (.A2( u2_u2_X_31 ) , .ZN( u2_u2_u5_n104 ) , .A1( u2_u2_u5_n181 ) );
  NAND2_X1 u2_u2_u5_U84 (.A2( u2_u2_X_34 ) , .A1( u2_u2_X_35 ) , .ZN( u2_u2_u5_n153 ) );
  NAND2_X1 u2_u2_u5_U85 (.A1( u2_u2_X_34 ) , .ZN( u2_u2_u5_n126 ) , .A2( u2_u2_u5_n171 ) );
  AND2_X1 u2_u2_u5_U86 (.A1( u2_u2_X_31 ) , .A2( u2_u2_X_32 ) , .ZN( u2_u2_u5_n106 ) );
  AND2_X1 u2_u2_u5_U87 (.A1( u2_u2_X_31 ) , .ZN( u2_u2_u5_n109 ) , .A2( u2_u2_u5_n181 ) );
  INV_X1 u2_u2_u5_U88 (.A( u2_u2_X_33 ) , .ZN( u2_u2_u5_n180 ) );
  INV_X1 u2_u2_u5_U89 (.A( u2_u2_X_35 ) , .ZN( u2_u2_u5_n171 ) );
  NOR2_X1 u2_u2_u5_U9 (.ZN( u2_u2_u5_n135 ) , .A1( u2_u2_u5_n173 ) , .A2( u2_u2_u5_n176 ) );
  INV_X1 u2_u2_u5_U90 (.A( u2_u2_X_36 ) , .ZN( u2_u2_u5_n170 ) );
  INV_X1 u2_u2_u5_U91 (.A( u2_u2_X_32 ) , .ZN( u2_u2_u5_n181 ) );
  NAND4_X1 u2_u2_u5_U92 (.ZN( u2_out2_29 ) , .A4( u2_u2_u5_n129 ) , .A3( u2_u2_u5_n130 ) , .A2( u2_u2_u5_n168 ) , .A1( u2_u2_u5_n196 ) );
  AOI221_X1 u2_u2_u5_U93 (.A( u2_u2_u5_n128 ) , .ZN( u2_u2_u5_n129 ) , .C2( u2_u2_u5_n132 ) , .B2( u2_u2_u5_n159 ) , .B1( u2_u2_u5_n176 ) , .C1( u2_u2_u5_n184 ) );
  AOI222_X1 u2_u2_u5_U94 (.ZN( u2_u2_u5_n130 ) , .A2( u2_u2_u5_n146 ) , .B1( u2_u2_u5_n147 ) , .C2( u2_u2_u5_n175 ) , .B2( u2_u2_u5_n179 ) , .A1( u2_u2_u5_n188 ) , .C1( u2_u2_u5_n194 ) );
  NAND4_X1 u2_u2_u5_U95 (.ZN( u2_out2_19 ) , .A4( u2_u2_u5_n166 ) , .A3( u2_u2_u5_n167 ) , .A2( u2_u2_u5_n168 ) , .A1( u2_u2_u5_n169 ) );
  AOI22_X1 u2_u2_u5_U96 (.B2( u2_u2_u5_n145 ) , .A2( u2_u2_u5_n146 ) , .ZN( u2_u2_u5_n167 ) , .B1( u2_u2_u5_n182 ) , .A1( u2_u2_u5_n189 ) );
  NOR4_X1 u2_u2_u5_U97 (.A4( u2_u2_u5_n162 ) , .A3( u2_u2_u5_n163 ) , .A2( u2_u2_u5_n164 ) , .A1( u2_u2_u5_n165 ) , .ZN( u2_u2_u5_n166 ) );
  NAND4_X1 u2_u2_u5_U98 (.ZN( u2_out2_11 ) , .A4( u2_u2_u5_n143 ) , .A3( u2_u2_u5_n144 ) , .A2( u2_u2_u5_n169 ) , .A1( u2_u2_u5_n196 ) );
  AOI22_X1 u2_u2_u5_U99 (.A2( u2_u2_u5_n132 ) , .ZN( u2_u2_u5_n144 ) , .B2( u2_u2_u5_n145 ) , .B1( u2_u2_u5_n184 ) , .A1( u2_u2_u5_n194 ) );
  OAI21_X1 u2_u2_u6_U10 (.A( u2_u2_u6_n159 ) , .B1( u2_u2_u6_n169 ) , .B2( u2_u2_u6_n173 ) , .ZN( u2_u2_u6_n90 ) );
  INV_X1 u2_u2_u6_U11 (.ZN( u2_u2_u6_n172 ) , .A( u2_u2_u6_n88 ) );
  AOI22_X1 u2_u2_u6_U12 (.A2( u2_u2_u6_n151 ) , .B2( u2_u2_u6_n161 ) , .A1( u2_u2_u6_n167 ) , .B1( u2_u2_u6_n170 ) , .ZN( u2_u2_u6_n89 ) );
  AOI21_X1 u2_u2_u6_U13 (.ZN( u2_u2_u6_n106 ) , .A( u2_u2_u6_n142 ) , .B2( u2_u2_u6_n159 ) , .B1( u2_u2_u6_n164 ) );
  INV_X1 u2_u2_u6_U14 (.A( u2_u2_u6_n155 ) , .ZN( u2_u2_u6_n161 ) );
  INV_X1 u2_u2_u6_U15 (.A( u2_u2_u6_n128 ) , .ZN( u2_u2_u6_n164 ) );
  NAND2_X1 u2_u2_u6_U16 (.ZN( u2_u2_u6_n110 ) , .A1( u2_u2_u6_n122 ) , .A2( u2_u2_u6_n129 ) );
  NAND2_X1 u2_u2_u6_U17 (.ZN( u2_u2_u6_n124 ) , .A2( u2_u2_u6_n146 ) , .A1( u2_u2_u6_n148 ) );
  INV_X1 u2_u2_u6_U18 (.A( u2_u2_u6_n132 ) , .ZN( u2_u2_u6_n171 ) );
  AND2_X1 u2_u2_u6_U19 (.A1( u2_u2_u6_n100 ) , .ZN( u2_u2_u6_n130 ) , .A2( u2_u2_u6_n147 ) );
  INV_X1 u2_u2_u6_U20 (.A( u2_u2_u6_n127 ) , .ZN( u2_u2_u6_n173 ) );
  INV_X1 u2_u2_u6_U21 (.A( u2_u2_u6_n121 ) , .ZN( u2_u2_u6_n167 ) );
  INV_X1 u2_u2_u6_U22 (.A( u2_u2_u6_n100 ) , .ZN( u2_u2_u6_n169 ) );
  INV_X1 u2_u2_u6_U23 (.A( u2_u2_u6_n123 ) , .ZN( u2_u2_u6_n170 ) );
  INV_X1 u2_u2_u6_U24 (.A( u2_u2_u6_n113 ) , .ZN( u2_u2_u6_n168 ) );
  AND2_X1 u2_u2_u6_U25 (.A1( u2_u2_u6_n107 ) , .A2( u2_u2_u6_n119 ) , .ZN( u2_u2_u6_n133 ) );
  AND2_X1 u2_u2_u6_U26 (.A2( u2_u2_u6_n121 ) , .A1( u2_u2_u6_n122 ) , .ZN( u2_u2_u6_n131 ) );
  AND3_X1 u2_u2_u6_U27 (.ZN( u2_u2_u6_n120 ) , .A2( u2_u2_u6_n127 ) , .A1( u2_u2_u6_n132 ) , .A3( u2_u2_u6_n145 ) );
  INV_X1 u2_u2_u6_U28 (.A( u2_u2_u6_n146 ) , .ZN( u2_u2_u6_n163 ) );
  AOI222_X1 u2_u2_u6_U29 (.ZN( u2_u2_u6_n114 ) , .A1( u2_u2_u6_n118 ) , .A2( u2_u2_u6_n126 ) , .B2( u2_u2_u6_n151 ) , .C2( u2_u2_u6_n159 ) , .C1( u2_u2_u6_n168 ) , .B1( u2_u2_u6_n169 ) );
  INV_X1 u2_u2_u6_U3 (.A( u2_u2_u6_n110 ) , .ZN( u2_u2_u6_n166 ) );
  NOR2_X1 u2_u2_u6_U30 (.A1( u2_u2_u6_n162 ) , .A2( u2_u2_u6_n165 ) , .ZN( u2_u2_u6_n98 ) );
  NAND2_X1 u2_u2_u6_U31 (.A1( u2_u2_u6_n144 ) , .ZN( u2_u2_u6_n151 ) , .A2( u2_u2_u6_n158 ) );
  NAND2_X1 u2_u2_u6_U32 (.ZN( u2_u2_u6_n132 ) , .A1( u2_u2_u6_n91 ) , .A2( u2_u2_u6_n97 ) );
  AOI22_X1 u2_u2_u6_U33 (.B2( u2_u2_u6_n110 ) , .B1( u2_u2_u6_n111 ) , .A1( u2_u2_u6_n112 ) , .ZN( u2_u2_u6_n115 ) , .A2( u2_u2_u6_n161 ) );
  NAND4_X1 u2_u2_u6_U34 (.A3( u2_u2_u6_n109 ) , .ZN( u2_u2_u6_n112 ) , .A4( u2_u2_u6_n132 ) , .A2( u2_u2_u6_n147 ) , .A1( u2_u2_u6_n166 ) );
  NOR2_X1 u2_u2_u6_U35 (.ZN( u2_u2_u6_n109 ) , .A1( u2_u2_u6_n170 ) , .A2( u2_u2_u6_n173 ) );
  NOR2_X1 u2_u2_u6_U36 (.A2( u2_u2_u6_n126 ) , .ZN( u2_u2_u6_n155 ) , .A1( u2_u2_u6_n160 ) );
  NAND2_X1 u2_u2_u6_U37 (.ZN( u2_u2_u6_n146 ) , .A2( u2_u2_u6_n94 ) , .A1( u2_u2_u6_n99 ) );
  AOI21_X1 u2_u2_u6_U38 (.A( u2_u2_u6_n144 ) , .B2( u2_u2_u6_n145 ) , .B1( u2_u2_u6_n146 ) , .ZN( u2_u2_u6_n150 ) );
  INV_X1 u2_u2_u6_U39 (.A( u2_u2_u6_n111 ) , .ZN( u2_u2_u6_n158 ) );
  INV_X1 u2_u2_u6_U4 (.A( u2_u2_u6_n142 ) , .ZN( u2_u2_u6_n174 ) );
  NAND2_X1 u2_u2_u6_U40 (.ZN( u2_u2_u6_n127 ) , .A1( u2_u2_u6_n91 ) , .A2( u2_u2_u6_n92 ) );
  NAND2_X1 u2_u2_u6_U41 (.ZN( u2_u2_u6_n129 ) , .A2( u2_u2_u6_n95 ) , .A1( u2_u2_u6_n96 ) );
  INV_X1 u2_u2_u6_U42 (.A( u2_u2_u6_n144 ) , .ZN( u2_u2_u6_n159 ) );
  NAND2_X1 u2_u2_u6_U43 (.ZN( u2_u2_u6_n145 ) , .A2( u2_u2_u6_n97 ) , .A1( u2_u2_u6_n98 ) );
  NAND2_X1 u2_u2_u6_U44 (.ZN( u2_u2_u6_n148 ) , .A2( u2_u2_u6_n92 ) , .A1( u2_u2_u6_n94 ) );
  NAND2_X1 u2_u2_u6_U45 (.ZN( u2_u2_u6_n108 ) , .A2( u2_u2_u6_n139 ) , .A1( u2_u2_u6_n144 ) );
  NAND2_X1 u2_u2_u6_U46 (.ZN( u2_u2_u6_n121 ) , .A2( u2_u2_u6_n95 ) , .A1( u2_u2_u6_n97 ) );
  NAND2_X1 u2_u2_u6_U47 (.ZN( u2_u2_u6_n107 ) , .A2( u2_u2_u6_n92 ) , .A1( u2_u2_u6_n95 ) );
  AND2_X1 u2_u2_u6_U48 (.ZN( u2_u2_u6_n118 ) , .A2( u2_u2_u6_n91 ) , .A1( u2_u2_u6_n99 ) );
  NAND2_X1 u2_u2_u6_U49 (.ZN( u2_u2_u6_n147 ) , .A2( u2_u2_u6_n98 ) , .A1( u2_u2_u6_n99 ) );
  NAND2_X1 u2_u2_u6_U5 (.A2( u2_u2_u6_n143 ) , .ZN( u2_u2_u6_n152 ) , .A1( u2_u2_u6_n166 ) );
  NAND2_X1 u2_u2_u6_U50 (.ZN( u2_u2_u6_n128 ) , .A1( u2_u2_u6_n94 ) , .A2( u2_u2_u6_n96 ) );
  AOI211_X1 u2_u2_u6_U51 (.B( u2_u2_u6_n134 ) , .A( u2_u2_u6_n135 ) , .C1( u2_u2_u6_n136 ) , .ZN( u2_u2_u6_n137 ) , .C2( u2_u2_u6_n151 ) );
  AOI21_X1 u2_u2_u6_U52 (.B2( u2_u2_u6_n132 ) , .B1( u2_u2_u6_n133 ) , .ZN( u2_u2_u6_n134 ) , .A( u2_u2_u6_n158 ) );
  AOI21_X1 u2_u2_u6_U53 (.B1( u2_u2_u6_n131 ) , .ZN( u2_u2_u6_n135 ) , .A( u2_u2_u6_n144 ) , .B2( u2_u2_u6_n146 ) );
  NAND4_X1 u2_u2_u6_U54 (.A4( u2_u2_u6_n127 ) , .A3( u2_u2_u6_n128 ) , .A2( u2_u2_u6_n129 ) , .A1( u2_u2_u6_n130 ) , .ZN( u2_u2_u6_n136 ) );
  NAND2_X1 u2_u2_u6_U55 (.ZN( u2_u2_u6_n119 ) , .A2( u2_u2_u6_n95 ) , .A1( u2_u2_u6_n99 ) );
  NAND2_X1 u2_u2_u6_U56 (.ZN( u2_u2_u6_n123 ) , .A2( u2_u2_u6_n91 ) , .A1( u2_u2_u6_n96 ) );
  NAND2_X1 u2_u2_u6_U57 (.ZN( u2_u2_u6_n100 ) , .A2( u2_u2_u6_n92 ) , .A1( u2_u2_u6_n98 ) );
  NAND2_X1 u2_u2_u6_U58 (.ZN( u2_u2_u6_n122 ) , .A1( u2_u2_u6_n94 ) , .A2( u2_u2_u6_n97 ) );
  INV_X1 u2_u2_u6_U59 (.A( u2_u2_u6_n139 ) , .ZN( u2_u2_u6_n160 ) );
  AOI22_X1 u2_u2_u6_U6 (.B2( u2_u2_u6_n101 ) , .A1( u2_u2_u6_n102 ) , .ZN( u2_u2_u6_n103 ) , .B1( u2_u2_u6_n160 ) , .A2( u2_u2_u6_n161 ) );
  NAND2_X1 u2_u2_u6_U60 (.ZN( u2_u2_u6_n113 ) , .A1( u2_u2_u6_n96 ) , .A2( u2_u2_u6_n98 ) );
  NOR2_X1 u2_u2_u6_U61 (.A2( u2_u2_X_40 ) , .A1( u2_u2_X_41 ) , .ZN( u2_u2_u6_n126 ) );
  NOR2_X1 u2_u2_u6_U62 (.A2( u2_u2_X_39 ) , .A1( u2_u2_X_42 ) , .ZN( u2_u2_u6_n92 ) );
  NOR2_X1 u2_u2_u6_U63 (.A2( u2_u2_X_39 ) , .A1( u2_u2_u6_n156 ) , .ZN( u2_u2_u6_n97 ) );
  NOR2_X1 u2_u2_u6_U64 (.A2( u2_u2_X_38 ) , .A1( u2_u2_u6_n165 ) , .ZN( u2_u2_u6_n95 ) );
  NOR2_X1 u2_u2_u6_U65 (.A2( u2_u2_X_41 ) , .ZN( u2_u2_u6_n111 ) , .A1( u2_u2_u6_n157 ) );
  NOR2_X1 u2_u2_u6_U66 (.A2( u2_u2_X_37 ) , .A1( u2_u2_u6_n162 ) , .ZN( u2_u2_u6_n94 ) );
  NOR2_X1 u2_u2_u6_U67 (.A2( u2_u2_X_37 ) , .A1( u2_u2_X_38 ) , .ZN( u2_u2_u6_n91 ) );
  NAND2_X1 u2_u2_u6_U68 (.A1( u2_u2_X_41 ) , .ZN( u2_u2_u6_n144 ) , .A2( u2_u2_u6_n157 ) );
  NAND2_X1 u2_u2_u6_U69 (.A2( u2_u2_X_40 ) , .A1( u2_u2_X_41 ) , .ZN( u2_u2_u6_n139 ) );
  NOR2_X1 u2_u2_u6_U7 (.A1( u2_u2_u6_n118 ) , .ZN( u2_u2_u6_n143 ) , .A2( u2_u2_u6_n168 ) );
  AND2_X1 u2_u2_u6_U70 (.A1( u2_u2_X_39 ) , .A2( u2_u2_u6_n156 ) , .ZN( u2_u2_u6_n96 ) );
  AND2_X1 u2_u2_u6_U71 (.A1( u2_u2_X_39 ) , .A2( u2_u2_X_42 ) , .ZN( u2_u2_u6_n99 ) );
  INV_X1 u2_u2_u6_U72 (.A( u2_u2_X_40 ) , .ZN( u2_u2_u6_n157 ) );
  INV_X1 u2_u2_u6_U73 (.A( u2_u2_X_37 ) , .ZN( u2_u2_u6_n165 ) );
  INV_X1 u2_u2_u6_U74 (.A( u2_u2_X_38 ) , .ZN( u2_u2_u6_n162 ) );
  INV_X1 u2_u2_u6_U75 (.A( u2_u2_X_42 ) , .ZN( u2_u2_u6_n156 ) );
  NAND4_X1 u2_u2_u6_U76 (.ZN( u2_out2_32 ) , .A4( u2_u2_u6_n103 ) , .A3( u2_u2_u6_n104 ) , .A2( u2_u2_u6_n105 ) , .A1( u2_u2_u6_n106 ) );
  AOI22_X1 u2_u2_u6_U77 (.ZN( u2_u2_u6_n105 ) , .A2( u2_u2_u6_n108 ) , .A1( u2_u2_u6_n118 ) , .B2( u2_u2_u6_n126 ) , .B1( u2_u2_u6_n171 ) );
  AOI22_X1 u2_u2_u6_U78 (.ZN( u2_u2_u6_n104 ) , .A1( u2_u2_u6_n111 ) , .B1( u2_u2_u6_n124 ) , .B2( u2_u2_u6_n151 ) , .A2( u2_u2_u6_n93 ) );
  NAND4_X1 u2_u2_u6_U79 (.ZN( u2_out2_12 ) , .A4( u2_u2_u6_n114 ) , .A3( u2_u2_u6_n115 ) , .A2( u2_u2_u6_n116 ) , .A1( u2_u2_u6_n117 ) );
  AOI21_X1 u2_u2_u6_U8 (.B1( u2_u2_u6_n107 ) , .B2( u2_u2_u6_n132 ) , .A( u2_u2_u6_n158 ) , .ZN( u2_u2_u6_n88 ) );
  OAI22_X1 u2_u2_u6_U80 (.B2( u2_u2_u6_n111 ) , .ZN( u2_u2_u6_n116 ) , .B1( u2_u2_u6_n126 ) , .A2( u2_u2_u6_n164 ) , .A1( u2_u2_u6_n167 ) );
  OAI21_X1 u2_u2_u6_U81 (.A( u2_u2_u6_n108 ) , .ZN( u2_u2_u6_n117 ) , .B2( u2_u2_u6_n141 ) , .B1( u2_u2_u6_n163 ) );
  OAI211_X1 u2_u2_u6_U82 (.ZN( u2_out2_7 ) , .B( u2_u2_u6_n153 ) , .C2( u2_u2_u6_n154 ) , .C1( u2_u2_u6_n155 ) , .A( u2_u2_u6_n174 ) );
  NOR3_X1 u2_u2_u6_U83 (.A1( u2_u2_u6_n141 ) , .ZN( u2_u2_u6_n154 ) , .A3( u2_u2_u6_n164 ) , .A2( u2_u2_u6_n171 ) );
  AOI211_X1 u2_u2_u6_U84 (.B( u2_u2_u6_n149 ) , .A( u2_u2_u6_n150 ) , .C2( u2_u2_u6_n151 ) , .C1( u2_u2_u6_n152 ) , .ZN( u2_u2_u6_n153 ) );
  OAI211_X1 u2_u2_u6_U85 (.ZN( u2_out2_22 ) , .B( u2_u2_u6_n137 ) , .A( u2_u2_u6_n138 ) , .C2( u2_u2_u6_n139 ) , .C1( u2_u2_u6_n140 ) );
  AOI22_X1 u2_u2_u6_U86 (.B1( u2_u2_u6_n124 ) , .A2( u2_u2_u6_n125 ) , .A1( u2_u2_u6_n126 ) , .ZN( u2_u2_u6_n138 ) , .B2( u2_u2_u6_n161 ) );
  AND4_X1 u2_u2_u6_U87 (.A3( u2_u2_u6_n119 ) , .A1( u2_u2_u6_n120 ) , .A4( u2_u2_u6_n129 ) , .ZN( u2_u2_u6_n140 ) , .A2( u2_u2_u6_n143 ) );
  NAND3_X1 u2_u2_u6_U88 (.A2( u2_u2_u6_n123 ) , .ZN( u2_u2_u6_n125 ) , .A1( u2_u2_u6_n130 ) , .A3( u2_u2_u6_n131 ) );
  NAND3_X1 u2_u2_u6_U89 (.A3( u2_u2_u6_n133 ) , .ZN( u2_u2_u6_n141 ) , .A1( u2_u2_u6_n145 ) , .A2( u2_u2_u6_n148 ) );
  AOI21_X1 u2_u2_u6_U9 (.B2( u2_u2_u6_n147 ) , .B1( u2_u2_u6_n148 ) , .ZN( u2_u2_u6_n149 ) , .A( u2_u2_u6_n158 ) );
  NAND3_X1 u2_u2_u6_U90 (.ZN( u2_u2_u6_n101 ) , .A3( u2_u2_u6_n107 ) , .A2( u2_u2_u6_n121 ) , .A1( u2_u2_u6_n127 ) );
  NAND3_X1 u2_u2_u6_U91 (.ZN( u2_u2_u6_n102 ) , .A3( u2_u2_u6_n130 ) , .A2( u2_u2_u6_n145 ) , .A1( u2_u2_u6_n166 ) );
  NAND3_X1 u2_u2_u6_U92 (.A3( u2_u2_u6_n113 ) , .A1( u2_u2_u6_n119 ) , .A2( u2_u2_u6_n123 ) , .ZN( u2_u2_u6_n93 ) );
  NAND3_X1 u2_u2_u6_U93 (.ZN( u2_u2_u6_n142 ) , .A2( u2_u2_u6_n172 ) , .A3( u2_u2_u6_n89 ) , .A1( u2_u2_u6_n90 ) );
  AND3_X1 u2_u2_u7_U10 (.A3( u2_u2_u7_n110 ) , .A2( u2_u2_u7_n127 ) , .A1( u2_u2_u7_n132 ) , .ZN( u2_u2_u7_n92 ) );
  OAI21_X1 u2_u2_u7_U11 (.A( u2_u2_u7_n161 ) , .B1( u2_u2_u7_n168 ) , .B2( u2_u2_u7_n173 ) , .ZN( u2_u2_u7_n91 ) );
  AOI211_X1 u2_u2_u7_U12 (.A( u2_u2_u7_n117 ) , .ZN( u2_u2_u7_n118 ) , .C2( u2_u2_u7_n126 ) , .C1( u2_u2_u7_n177 ) , .B( u2_u2_u7_n180 ) );
  OAI22_X1 u2_u2_u7_U13 (.B1( u2_u2_u7_n115 ) , .ZN( u2_u2_u7_n117 ) , .A2( u2_u2_u7_n133 ) , .A1( u2_u2_u7_n137 ) , .B2( u2_u2_u7_n162 ) );
  INV_X1 u2_u2_u7_U14 (.A( u2_u2_u7_n116 ) , .ZN( u2_u2_u7_n180 ) );
  NOR3_X1 u2_u2_u7_U15 (.ZN( u2_u2_u7_n115 ) , .A3( u2_u2_u7_n145 ) , .A2( u2_u2_u7_n168 ) , .A1( u2_u2_u7_n169 ) );
  OAI211_X1 u2_u2_u7_U16 (.B( u2_u2_u7_n122 ) , .A( u2_u2_u7_n123 ) , .C2( u2_u2_u7_n124 ) , .ZN( u2_u2_u7_n154 ) , .C1( u2_u2_u7_n162 ) );
  AOI222_X1 u2_u2_u7_U17 (.ZN( u2_u2_u7_n122 ) , .C2( u2_u2_u7_n126 ) , .C1( u2_u2_u7_n145 ) , .B1( u2_u2_u7_n161 ) , .A2( u2_u2_u7_n165 ) , .B2( u2_u2_u7_n170 ) , .A1( u2_u2_u7_n176 ) );
  INV_X1 u2_u2_u7_U18 (.A( u2_u2_u7_n133 ) , .ZN( u2_u2_u7_n176 ) );
  NOR3_X1 u2_u2_u7_U19 (.A2( u2_u2_u7_n134 ) , .A1( u2_u2_u7_n135 ) , .ZN( u2_u2_u7_n136 ) , .A3( u2_u2_u7_n171 ) );
  NOR2_X1 u2_u2_u7_U20 (.A1( u2_u2_u7_n130 ) , .A2( u2_u2_u7_n134 ) , .ZN( u2_u2_u7_n153 ) );
  INV_X1 u2_u2_u7_U21 (.A( u2_u2_u7_n101 ) , .ZN( u2_u2_u7_n165 ) );
  NOR2_X1 u2_u2_u7_U22 (.ZN( u2_u2_u7_n111 ) , .A2( u2_u2_u7_n134 ) , .A1( u2_u2_u7_n169 ) );
  AOI21_X1 u2_u2_u7_U23 (.ZN( u2_u2_u7_n104 ) , .B2( u2_u2_u7_n112 ) , .B1( u2_u2_u7_n127 ) , .A( u2_u2_u7_n164 ) );
  AOI21_X1 u2_u2_u7_U24 (.ZN( u2_u2_u7_n106 ) , .B1( u2_u2_u7_n133 ) , .B2( u2_u2_u7_n146 ) , .A( u2_u2_u7_n162 ) );
  AOI21_X1 u2_u2_u7_U25 (.A( u2_u2_u7_n101 ) , .ZN( u2_u2_u7_n107 ) , .B2( u2_u2_u7_n128 ) , .B1( u2_u2_u7_n175 ) );
  INV_X1 u2_u2_u7_U26 (.A( u2_u2_u7_n138 ) , .ZN( u2_u2_u7_n171 ) );
  INV_X1 u2_u2_u7_U27 (.A( u2_u2_u7_n131 ) , .ZN( u2_u2_u7_n177 ) );
  INV_X1 u2_u2_u7_U28 (.A( u2_u2_u7_n110 ) , .ZN( u2_u2_u7_n174 ) );
  NAND2_X1 u2_u2_u7_U29 (.A1( u2_u2_u7_n129 ) , .A2( u2_u2_u7_n132 ) , .ZN( u2_u2_u7_n149 ) );
  OAI21_X1 u2_u2_u7_U3 (.ZN( u2_u2_u7_n159 ) , .A( u2_u2_u7_n165 ) , .B2( u2_u2_u7_n171 ) , .B1( u2_u2_u7_n174 ) );
  NAND2_X1 u2_u2_u7_U30 (.A1( u2_u2_u7_n113 ) , .A2( u2_u2_u7_n124 ) , .ZN( u2_u2_u7_n130 ) );
  INV_X1 u2_u2_u7_U31 (.A( u2_u2_u7_n112 ) , .ZN( u2_u2_u7_n173 ) );
  INV_X1 u2_u2_u7_U32 (.A( u2_u2_u7_n128 ) , .ZN( u2_u2_u7_n168 ) );
  INV_X1 u2_u2_u7_U33 (.A( u2_u2_u7_n148 ) , .ZN( u2_u2_u7_n169 ) );
  INV_X1 u2_u2_u7_U34 (.A( u2_u2_u7_n127 ) , .ZN( u2_u2_u7_n179 ) );
  NOR2_X1 u2_u2_u7_U35 (.ZN( u2_u2_u7_n101 ) , .A2( u2_u2_u7_n150 ) , .A1( u2_u2_u7_n156 ) );
  AOI211_X1 u2_u2_u7_U36 (.B( u2_u2_u7_n154 ) , .A( u2_u2_u7_n155 ) , .C1( u2_u2_u7_n156 ) , .ZN( u2_u2_u7_n157 ) , .C2( u2_u2_u7_n172 ) );
  INV_X1 u2_u2_u7_U37 (.A( u2_u2_u7_n153 ) , .ZN( u2_u2_u7_n172 ) );
  AOI211_X1 u2_u2_u7_U38 (.B( u2_u2_u7_n139 ) , .A( u2_u2_u7_n140 ) , .C2( u2_u2_u7_n141 ) , .ZN( u2_u2_u7_n142 ) , .C1( u2_u2_u7_n156 ) );
  NAND4_X1 u2_u2_u7_U39 (.A3( u2_u2_u7_n127 ) , .A2( u2_u2_u7_n128 ) , .A1( u2_u2_u7_n129 ) , .ZN( u2_u2_u7_n141 ) , .A4( u2_u2_u7_n147 ) );
  INV_X1 u2_u2_u7_U4 (.A( u2_u2_u7_n111 ) , .ZN( u2_u2_u7_n170 ) );
  AOI21_X1 u2_u2_u7_U40 (.A( u2_u2_u7_n137 ) , .B1( u2_u2_u7_n138 ) , .ZN( u2_u2_u7_n139 ) , .B2( u2_u2_u7_n146 ) );
  OAI22_X1 u2_u2_u7_U41 (.B1( u2_u2_u7_n136 ) , .ZN( u2_u2_u7_n140 ) , .A1( u2_u2_u7_n153 ) , .B2( u2_u2_u7_n162 ) , .A2( u2_u2_u7_n164 ) );
  AOI21_X1 u2_u2_u7_U42 (.ZN( u2_u2_u7_n123 ) , .B1( u2_u2_u7_n165 ) , .B2( u2_u2_u7_n177 ) , .A( u2_u2_u7_n97 ) );
  AOI21_X1 u2_u2_u7_U43 (.B2( u2_u2_u7_n113 ) , .B1( u2_u2_u7_n124 ) , .A( u2_u2_u7_n125 ) , .ZN( u2_u2_u7_n97 ) );
  INV_X1 u2_u2_u7_U44 (.A( u2_u2_u7_n125 ) , .ZN( u2_u2_u7_n161 ) );
  INV_X1 u2_u2_u7_U45 (.A( u2_u2_u7_n152 ) , .ZN( u2_u2_u7_n162 ) );
  AOI22_X1 u2_u2_u7_U46 (.A2( u2_u2_u7_n114 ) , .ZN( u2_u2_u7_n119 ) , .B1( u2_u2_u7_n130 ) , .A1( u2_u2_u7_n156 ) , .B2( u2_u2_u7_n165 ) );
  NAND2_X1 u2_u2_u7_U47 (.A2( u2_u2_u7_n112 ) , .ZN( u2_u2_u7_n114 ) , .A1( u2_u2_u7_n175 ) );
  AND2_X1 u2_u2_u7_U48 (.ZN( u2_u2_u7_n145 ) , .A2( u2_u2_u7_n98 ) , .A1( u2_u2_u7_n99 ) );
  NOR2_X1 u2_u2_u7_U49 (.ZN( u2_u2_u7_n137 ) , .A1( u2_u2_u7_n150 ) , .A2( u2_u2_u7_n161 ) );
  INV_X1 u2_u2_u7_U5 (.A( u2_u2_u7_n149 ) , .ZN( u2_u2_u7_n175 ) );
  AOI21_X1 u2_u2_u7_U50 (.ZN( u2_u2_u7_n105 ) , .B2( u2_u2_u7_n110 ) , .A( u2_u2_u7_n125 ) , .B1( u2_u2_u7_n147 ) );
  NAND2_X1 u2_u2_u7_U51 (.ZN( u2_u2_u7_n146 ) , .A1( u2_u2_u7_n95 ) , .A2( u2_u2_u7_n98 ) );
  NAND2_X1 u2_u2_u7_U52 (.A2( u2_u2_u7_n103 ) , .ZN( u2_u2_u7_n147 ) , .A1( u2_u2_u7_n93 ) );
  NAND2_X1 u2_u2_u7_U53 (.A1( u2_u2_u7_n103 ) , .ZN( u2_u2_u7_n127 ) , .A2( u2_u2_u7_n99 ) );
  OR2_X1 u2_u2_u7_U54 (.ZN( u2_u2_u7_n126 ) , .A2( u2_u2_u7_n152 ) , .A1( u2_u2_u7_n156 ) );
  NAND2_X1 u2_u2_u7_U55 (.A2( u2_u2_u7_n102 ) , .A1( u2_u2_u7_n103 ) , .ZN( u2_u2_u7_n133 ) );
  NAND2_X1 u2_u2_u7_U56 (.ZN( u2_u2_u7_n112 ) , .A2( u2_u2_u7_n96 ) , .A1( u2_u2_u7_n99 ) );
  NAND2_X1 u2_u2_u7_U57 (.A2( u2_u2_u7_n102 ) , .ZN( u2_u2_u7_n128 ) , .A1( u2_u2_u7_n98 ) );
  NAND2_X1 u2_u2_u7_U58 (.A1( u2_u2_u7_n100 ) , .ZN( u2_u2_u7_n113 ) , .A2( u2_u2_u7_n93 ) );
  NAND2_X1 u2_u2_u7_U59 (.A2( u2_u2_u7_n102 ) , .ZN( u2_u2_u7_n124 ) , .A1( u2_u2_u7_n96 ) );
  INV_X1 u2_u2_u7_U6 (.A( u2_u2_u7_n154 ) , .ZN( u2_u2_u7_n178 ) );
  NAND2_X1 u2_u2_u7_U60 (.ZN( u2_u2_u7_n110 ) , .A1( u2_u2_u7_n95 ) , .A2( u2_u2_u7_n96 ) );
  INV_X1 u2_u2_u7_U61 (.A( u2_u2_u7_n150 ) , .ZN( u2_u2_u7_n164 ) );
  AND2_X1 u2_u2_u7_U62 (.ZN( u2_u2_u7_n134 ) , .A1( u2_u2_u7_n93 ) , .A2( u2_u2_u7_n98 ) );
  NAND2_X1 u2_u2_u7_U63 (.A1( u2_u2_u7_n100 ) , .A2( u2_u2_u7_n102 ) , .ZN( u2_u2_u7_n129 ) );
  NAND2_X1 u2_u2_u7_U64 (.A2( u2_u2_u7_n103 ) , .ZN( u2_u2_u7_n131 ) , .A1( u2_u2_u7_n95 ) );
  NAND2_X1 u2_u2_u7_U65 (.A1( u2_u2_u7_n100 ) , .ZN( u2_u2_u7_n138 ) , .A2( u2_u2_u7_n99 ) );
  NAND2_X1 u2_u2_u7_U66 (.ZN( u2_u2_u7_n132 ) , .A1( u2_u2_u7_n93 ) , .A2( u2_u2_u7_n96 ) );
  NAND2_X1 u2_u2_u7_U67 (.A1( u2_u2_u7_n100 ) , .ZN( u2_u2_u7_n148 ) , .A2( u2_u2_u7_n95 ) );
  NOR2_X1 u2_u2_u7_U68 (.A2( u2_u2_X_47 ) , .ZN( u2_u2_u7_n150 ) , .A1( u2_u2_u7_n163 ) );
  NOR2_X1 u2_u2_u7_U69 (.A2( u2_u2_X_43 ) , .A1( u2_u2_X_44 ) , .ZN( u2_u2_u7_n103 ) );
  AOI211_X1 u2_u2_u7_U7 (.ZN( u2_u2_u7_n116 ) , .A( u2_u2_u7_n155 ) , .C1( u2_u2_u7_n161 ) , .C2( u2_u2_u7_n171 ) , .B( u2_u2_u7_n94 ) );
  NOR2_X1 u2_u2_u7_U70 (.A2( u2_u2_X_48 ) , .A1( u2_u2_u7_n166 ) , .ZN( u2_u2_u7_n95 ) );
  NOR2_X1 u2_u2_u7_U71 (.A2( u2_u2_X_45 ) , .A1( u2_u2_X_48 ) , .ZN( u2_u2_u7_n99 ) );
  NOR2_X1 u2_u2_u7_U72 (.A2( u2_u2_X_44 ) , .A1( u2_u2_u7_n167 ) , .ZN( u2_u2_u7_n98 ) );
  NOR2_X1 u2_u2_u7_U73 (.A2( u2_u2_X_46 ) , .A1( u2_u2_X_47 ) , .ZN( u2_u2_u7_n152 ) );
  AND2_X1 u2_u2_u7_U74 (.A1( u2_u2_X_47 ) , .ZN( u2_u2_u7_n156 ) , .A2( u2_u2_u7_n163 ) );
  NAND2_X1 u2_u2_u7_U75 (.A2( u2_u2_X_46 ) , .A1( u2_u2_X_47 ) , .ZN( u2_u2_u7_n125 ) );
  AND2_X1 u2_u2_u7_U76 (.A2( u2_u2_X_45 ) , .A1( u2_u2_X_48 ) , .ZN( u2_u2_u7_n102 ) );
  AND2_X1 u2_u2_u7_U77 (.A2( u2_u2_X_43 ) , .A1( u2_u2_X_44 ) , .ZN( u2_u2_u7_n96 ) );
  AND2_X1 u2_u2_u7_U78 (.A1( u2_u2_X_44 ) , .ZN( u2_u2_u7_n100 ) , .A2( u2_u2_u7_n167 ) );
  AND2_X1 u2_u2_u7_U79 (.A1( u2_u2_X_48 ) , .A2( u2_u2_u7_n166 ) , .ZN( u2_u2_u7_n93 ) );
  OAI222_X1 u2_u2_u7_U8 (.C2( u2_u2_u7_n101 ) , .B2( u2_u2_u7_n111 ) , .A1( u2_u2_u7_n113 ) , .C1( u2_u2_u7_n146 ) , .A2( u2_u2_u7_n162 ) , .B1( u2_u2_u7_n164 ) , .ZN( u2_u2_u7_n94 ) );
  INV_X1 u2_u2_u7_U80 (.A( u2_u2_X_46 ) , .ZN( u2_u2_u7_n163 ) );
  INV_X1 u2_u2_u7_U81 (.A( u2_u2_X_43 ) , .ZN( u2_u2_u7_n167 ) );
  INV_X1 u2_u2_u7_U82 (.A( u2_u2_X_45 ) , .ZN( u2_u2_u7_n166 ) );
  NAND4_X1 u2_u2_u7_U83 (.ZN( u2_out2_5 ) , .A4( u2_u2_u7_n108 ) , .A3( u2_u2_u7_n109 ) , .A1( u2_u2_u7_n116 ) , .A2( u2_u2_u7_n123 ) );
  AOI22_X1 u2_u2_u7_U84 (.ZN( u2_u2_u7_n109 ) , .A2( u2_u2_u7_n126 ) , .B2( u2_u2_u7_n145 ) , .B1( u2_u2_u7_n156 ) , .A1( u2_u2_u7_n171 ) );
  NOR4_X1 u2_u2_u7_U85 (.A4( u2_u2_u7_n104 ) , .A3( u2_u2_u7_n105 ) , .A2( u2_u2_u7_n106 ) , .A1( u2_u2_u7_n107 ) , .ZN( u2_u2_u7_n108 ) );
  NAND4_X1 u2_u2_u7_U86 (.ZN( u2_out2_27 ) , .A4( u2_u2_u7_n118 ) , .A3( u2_u2_u7_n119 ) , .A2( u2_u2_u7_n120 ) , .A1( u2_u2_u7_n121 ) );
  OAI21_X1 u2_u2_u7_U87 (.ZN( u2_u2_u7_n121 ) , .B2( u2_u2_u7_n145 ) , .A( u2_u2_u7_n150 ) , .B1( u2_u2_u7_n174 ) );
  OAI21_X1 u2_u2_u7_U88 (.ZN( u2_u2_u7_n120 ) , .A( u2_u2_u7_n161 ) , .B2( u2_u2_u7_n170 ) , .B1( u2_u2_u7_n179 ) );
  NAND4_X1 u2_u2_u7_U89 (.ZN( u2_out2_21 ) , .A4( u2_u2_u7_n157 ) , .A3( u2_u2_u7_n158 ) , .A2( u2_u2_u7_n159 ) , .A1( u2_u2_u7_n160 ) );
  OAI221_X1 u2_u2_u7_U9 (.C1( u2_u2_u7_n101 ) , .C2( u2_u2_u7_n147 ) , .ZN( u2_u2_u7_n155 ) , .B2( u2_u2_u7_n162 ) , .A( u2_u2_u7_n91 ) , .B1( u2_u2_u7_n92 ) );
  OAI21_X1 u2_u2_u7_U90 (.B1( u2_u2_u7_n145 ) , .ZN( u2_u2_u7_n160 ) , .A( u2_u2_u7_n161 ) , .B2( u2_u2_u7_n177 ) );
  AOI22_X1 u2_u2_u7_U91 (.B2( u2_u2_u7_n149 ) , .B1( u2_u2_u7_n150 ) , .A2( u2_u2_u7_n151 ) , .A1( u2_u2_u7_n152 ) , .ZN( u2_u2_u7_n158 ) );
  NAND4_X1 u2_u2_u7_U92 (.ZN( u2_out2_15 ) , .A4( u2_u2_u7_n142 ) , .A3( u2_u2_u7_n143 ) , .A2( u2_u2_u7_n144 ) , .A1( u2_u2_u7_n178 ) );
  OR2_X1 u2_u2_u7_U93 (.A2( u2_u2_u7_n125 ) , .A1( u2_u2_u7_n129 ) , .ZN( u2_u2_u7_n144 ) );
  AOI22_X1 u2_u2_u7_U94 (.A2( u2_u2_u7_n126 ) , .ZN( u2_u2_u7_n143 ) , .B2( u2_u2_u7_n165 ) , .B1( u2_u2_u7_n173 ) , .A1( u2_u2_u7_n174 ) );
  NAND3_X1 u2_u2_u7_U95 (.A3( u2_u2_u7_n146 ) , .A2( u2_u2_u7_n147 ) , .A1( u2_u2_u7_n148 ) , .ZN( u2_u2_u7_n151 ) );
  NAND3_X1 u2_u2_u7_U96 (.A3( u2_u2_u7_n131 ) , .A2( u2_u2_u7_n132 ) , .A1( u2_u2_u7_n133 ) , .ZN( u2_u2_u7_n135 ) );
  XOR2_X1 u2_u3_U20 (.B( u2_K4_36 ) , .A( u2_R2_25 ) , .Z( u2_u3_X_36 ) );
  XOR2_X1 u2_u3_U21 (.B( u2_K4_35 ) , .A( u2_R2_24 ) , .Z( u2_u3_X_35 ) );
  XOR2_X1 u2_u3_U22 (.B( u2_K4_34 ) , .A( u2_R2_23 ) , .Z( u2_u3_X_34 ) );
  XOR2_X1 u2_u3_U23 (.B( u2_K4_33 ) , .A( u2_R2_22 ) , .Z( u2_u3_X_33 ) );
  XOR2_X1 u2_u3_U24 (.B( u2_K4_32 ) , .A( u2_R2_21 ) , .Z( u2_u3_X_32 ) );
  XOR2_X1 u2_u3_U25 (.B( u2_K4_31 ) , .A( u2_R2_20 ) , .Z( u2_u3_X_31 ) );
  XOR2_X1 u2_u3_U26 (.B( u2_K4_30 ) , .A( u2_R2_21 ) , .Z( u2_u3_X_30 ) );
  XOR2_X1 u2_u3_U28 (.B( u2_K4_29 ) , .A( u2_R2_20 ) , .Z( u2_u3_X_29 ) );
  XOR2_X1 u2_u3_U29 (.B( u2_K4_28 ) , .A( u2_R2_19 ) , .Z( u2_u3_X_28 ) );
  XOR2_X1 u2_u3_U30 (.B( u2_K4_27 ) , .A( u2_R2_18 ) , .Z( u2_u3_X_27 ) );
  XOR2_X1 u2_u3_U31 (.B( u2_K4_26 ) , .A( u2_R2_17 ) , .Z( u2_u3_X_26 ) );
  XOR2_X1 u2_u3_U32 (.B( u2_K4_25 ) , .A( u2_R2_16 ) , .Z( u2_u3_X_25 ) );
  XOR2_X1 u2_u3_U33 (.B( u2_K4_24 ) , .A( u2_R2_17 ) , .Z( u2_u3_X_24 ) );
  XOR2_X1 u2_u3_U34 (.B( u2_K4_23 ) , .A( u2_R2_16 ) , .Z( u2_u3_X_23 ) );
  XOR2_X1 u2_u3_U35 (.B( u2_K4_22 ) , .A( u2_R2_15 ) , .Z( u2_u3_X_22 ) );
  XOR2_X1 u2_u3_U36 (.B( u2_K4_21 ) , .A( u2_R2_14 ) , .Z( u2_u3_X_21 ) );
  XOR2_X1 u2_u3_U37 (.B( u2_K4_20 ) , .A( u2_R2_13 ) , .Z( u2_u3_X_20 ) );
  XOR2_X1 u2_u3_U39 (.B( u2_K4_19 ) , .A( u2_R2_12 ) , .Z( u2_u3_X_19 ) );
  XOR2_X1 u2_u3_U40 (.B( u2_K4_18 ) , .A( u2_R2_13 ) , .Z( u2_u3_X_18 ) );
  XOR2_X1 u2_u3_U41 (.B( u2_K4_17 ) , .A( u2_R2_12 ) , .Z( u2_u3_X_17 ) );
  XOR2_X1 u2_u3_U42 (.B( u2_K4_16 ) , .A( u2_R2_11 ) , .Z( u2_u3_X_16 ) );
  XOR2_X1 u2_u3_U43 (.B( u2_K4_15 ) , .A( u2_R2_10 ) , .Z( u2_u3_X_15 ) );
  XOR2_X1 u2_u3_U44 (.B( u2_K4_14 ) , .A( u2_R2_9 ) , .Z( u2_u3_X_14 ) );
  XOR2_X1 u2_u3_U45 (.B( u2_K4_13 ) , .A( u2_R2_8 ) , .Z( u2_u3_X_13 ) );
  OAI22_X1 u2_u3_u2_U10 (.B1( u2_u3_u2_n151 ) , .A2( u2_u3_u2_n152 ) , .A1( u2_u3_u2_n153 ) , .ZN( u2_u3_u2_n160 ) , .B2( u2_u3_u2_n168 ) );
  NAND3_X1 u2_u3_u2_U100 (.A2( u2_u3_u2_n100 ) , .A1( u2_u3_u2_n104 ) , .A3( u2_u3_u2_n138 ) , .ZN( u2_u3_u2_n98 ) );
  NOR3_X1 u2_u3_u2_U11 (.A1( u2_u3_u2_n150 ) , .ZN( u2_u3_u2_n151 ) , .A3( u2_u3_u2_n175 ) , .A2( u2_u3_u2_n188 ) );
  AOI21_X1 u2_u3_u2_U12 (.B2( u2_u3_u2_n123 ) , .ZN( u2_u3_u2_n125 ) , .A( u2_u3_u2_n171 ) , .B1( u2_u3_u2_n184 ) );
  INV_X1 u2_u3_u2_U13 (.A( u2_u3_u2_n150 ) , .ZN( u2_u3_u2_n184 ) );
  AOI21_X1 u2_u3_u2_U14 (.ZN( u2_u3_u2_n144 ) , .B2( u2_u3_u2_n155 ) , .A( u2_u3_u2_n172 ) , .B1( u2_u3_u2_n185 ) );
  AOI21_X1 u2_u3_u2_U15 (.B2( u2_u3_u2_n143 ) , .ZN( u2_u3_u2_n145 ) , .B1( u2_u3_u2_n152 ) , .A( u2_u3_u2_n171 ) );
  INV_X1 u2_u3_u2_U16 (.A( u2_u3_u2_n156 ) , .ZN( u2_u3_u2_n171 ) );
  INV_X1 u2_u3_u2_U17 (.A( u2_u3_u2_n120 ) , .ZN( u2_u3_u2_n188 ) );
  NAND2_X1 u2_u3_u2_U18 (.A2( u2_u3_u2_n122 ) , .ZN( u2_u3_u2_n150 ) , .A1( u2_u3_u2_n152 ) );
  INV_X1 u2_u3_u2_U19 (.A( u2_u3_u2_n153 ) , .ZN( u2_u3_u2_n170 ) );
  INV_X1 u2_u3_u2_U20 (.A( u2_u3_u2_n137 ) , .ZN( u2_u3_u2_n173 ) );
  NAND2_X1 u2_u3_u2_U21 (.A1( u2_u3_u2_n132 ) , .A2( u2_u3_u2_n139 ) , .ZN( u2_u3_u2_n157 ) );
  INV_X1 u2_u3_u2_U22 (.A( u2_u3_u2_n113 ) , .ZN( u2_u3_u2_n178 ) );
  INV_X1 u2_u3_u2_U23 (.A( u2_u3_u2_n139 ) , .ZN( u2_u3_u2_n175 ) );
  INV_X1 u2_u3_u2_U24 (.A( u2_u3_u2_n155 ) , .ZN( u2_u3_u2_n181 ) );
  INV_X1 u2_u3_u2_U25 (.A( u2_u3_u2_n119 ) , .ZN( u2_u3_u2_n177 ) );
  INV_X1 u2_u3_u2_U26 (.A( u2_u3_u2_n116 ) , .ZN( u2_u3_u2_n180 ) );
  INV_X1 u2_u3_u2_U27 (.A( u2_u3_u2_n131 ) , .ZN( u2_u3_u2_n179 ) );
  INV_X1 u2_u3_u2_U28 (.A( u2_u3_u2_n154 ) , .ZN( u2_u3_u2_n176 ) );
  NAND2_X1 u2_u3_u2_U29 (.A2( u2_u3_u2_n116 ) , .A1( u2_u3_u2_n117 ) , .ZN( u2_u3_u2_n118 ) );
  NOR2_X1 u2_u3_u2_U3 (.ZN( u2_u3_u2_n121 ) , .A2( u2_u3_u2_n177 ) , .A1( u2_u3_u2_n180 ) );
  INV_X1 u2_u3_u2_U30 (.A( u2_u3_u2_n132 ) , .ZN( u2_u3_u2_n182 ) );
  INV_X1 u2_u3_u2_U31 (.A( u2_u3_u2_n158 ) , .ZN( u2_u3_u2_n183 ) );
  OAI21_X1 u2_u3_u2_U32 (.A( u2_u3_u2_n156 ) , .B1( u2_u3_u2_n157 ) , .ZN( u2_u3_u2_n158 ) , .B2( u2_u3_u2_n179 ) );
  NOR2_X1 u2_u3_u2_U33 (.ZN( u2_u3_u2_n156 ) , .A1( u2_u3_u2_n166 ) , .A2( u2_u3_u2_n169 ) );
  NOR2_X1 u2_u3_u2_U34 (.A2( u2_u3_u2_n114 ) , .ZN( u2_u3_u2_n137 ) , .A1( u2_u3_u2_n140 ) );
  NOR2_X1 u2_u3_u2_U35 (.A2( u2_u3_u2_n138 ) , .ZN( u2_u3_u2_n153 ) , .A1( u2_u3_u2_n156 ) );
  AOI211_X1 u2_u3_u2_U36 (.ZN( u2_u3_u2_n130 ) , .C1( u2_u3_u2_n138 ) , .C2( u2_u3_u2_n179 ) , .B( u2_u3_u2_n96 ) , .A( u2_u3_u2_n97 ) );
  OAI22_X1 u2_u3_u2_U37 (.B1( u2_u3_u2_n133 ) , .A2( u2_u3_u2_n137 ) , .A1( u2_u3_u2_n152 ) , .B2( u2_u3_u2_n168 ) , .ZN( u2_u3_u2_n97 ) );
  OAI221_X1 u2_u3_u2_U38 (.B1( u2_u3_u2_n113 ) , .C1( u2_u3_u2_n132 ) , .A( u2_u3_u2_n149 ) , .B2( u2_u3_u2_n171 ) , .C2( u2_u3_u2_n172 ) , .ZN( u2_u3_u2_n96 ) );
  OAI221_X1 u2_u3_u2_U39 (.A( u2_u3_u2_n115 ) , .C2( u2_u3_u2_n123 ) , .B2( u2_u3_u2_n143 ) , .B1( u2_u3_u2_n153 ) , .ZN( u2_u3_u2_n163 ) , .C1( u2_u3_u2_n168 ) );
  INV_X1 u2_u3_u2_U4 (.A( u2_u3_u2_n134 ) , .ZN( u2_u3_u2_n185 ) );
  OAI21_X1 u2_u3_u2_U40 (.A( u2_u3_u2_n114 ) , .ZN( u2_u3_u2_n115 ) , .B1( u2_u3_u2_n176 ) , .B2( u2_u3_u2_n178 ) );
  OAI221_X1 u2_u3_u2_U41 (.A( u2_u3_u2_n135 ) , .B2( u2_u3_u2_n136 ) , .B1( u2_u3_u2_n137 ) , .ZN( u2_u3_u2_n162 ) , .C2( u2_u3_u2_n167 ) , .C1( u2_u3_u2_n185 ) );
  AND3_X1 u2_u3_u2_U42 (.A3( u2_u3_u2_n131 ) , .A2( u2_u3_u2_n132 ) , .A1( u2_u3_u2_n133 ) , .ZN( u2_u3_u2_n136 ) );
  AOI22_X1 u2_u3_u2_U43 (.ZN( u2_u3_u2_n135 ) , .B1( u2_u3_u2_n140 ) , .A1( u2_u3_u2_n156 ) , .B2( u2_u3_u2_n180 ) , .A2( u2_u3_u2_n188 ) );
  AOI21_X1 u2_u3_u2_U44 (.ZN( u2_u3_u2_n149 ) , .B1( u2_u3_u2_n173 ) , .B2( u2_u3_u2_n188 ) , .A( u2_u3_u2_n95 ) );
  AND3_X1 u2_u3_u2_U45 (.A2( u2_u3_u2_n100 ) , .A1( u2_u3_u2_n104 ) , .A3( u2_u3_u2_n156 ) , .ZN( u2_u3_u2_n95 ) );
  OAI21_X1 u2_u3_u2_U46 (.A( u2_u3_u2_n141 ) , .B2( u2_u3_u2_n142 ) , .ZN( u2_u3_u2_n146 ) , .B1( u2_u3_u2_n153 ) );
  OAI21_X1 u2_u3_u2_U47 (.A( u2_u3_u2_n140 ) , .ZN( u2_u3_u2_n141 ) , .B1( u2_u3_u2_n176 ) , .B2( u2_u3_u2_n177 ) );
  NOR3_X1 u2_u3_u2_U48 (.ZN( u2_u3_u2_n142 ) , .A3( u2_u3_u2_n175 ) , .A2( u2_u3_u2_n178 ) , .A1( u2_u3_u2_n181 ) );
  OAI21_X1 u2_u3_u2_U49 (.A( u2_u3_u2_n101 ) , .B2( u2_u3_u2_n121 ) , .B1( u2_u3_u2_n153 ) , .ZN( u2_u3_u2_n164 ) );
  NOR4_X1 u2_u3_u2_U5 (.A4( u2_u3_u2_n124 ) , .A3( u2_u3_u2_n125 ) , .A2( u2_u3_u2_n126 ) , .A1( u2_u3_u2_n127 ) , .ZN( u2_u3_u2_n128 ) );
  NAND2_X1 u2_u3_u2_U50 (.A2( u2_u3_u2_n100 ) , .A1( u2_u3_u2_n107 ) , .ZN( u2_u3_u2_n155 ) );
  NAND2_X1 u2_u3_u2_U51 (.A2( u2_u3_u2_n105 ) , .A1( u2_u3_u2_n108 ) , .ZN( u2_u3_u2_n143 ) );
  NAND2_X1 u2_u3_u2_U52 (.A1( u2_u3_u2_n104 ) , .A2( u2_u3_u2_n106 ) , .ZN( u2_u3_u2_n152 ) );
  NAND2_X1 u2_u3_u2_U53 (.A1( u2_u3_u2_n100 ) , .A2( u2_u3_u2_n105 ) , .ZN( u2_u3_u2_n132 ) );
  INV_X1 u2_u3_u2_U54 (.A( u2_u3_u2_n140 ) , .ZN( u2_u3_u2_n168 ) );
  INV_X1 u2_u3_u2_U55 (.A( u2_u3_u2_n138 ) , .ZN( u2_u3_u2_n167 ) );
  INV_X1 u2_u3_u2_U56 (.ZN( u2_u3_u2_n187 ) , .A( u2_u3_u2_n99 ) );
  OAI21_X1 u2_u3_u2_U57 (.B1( u2_u3_u2_n137 ) , .B2( u2_u3_u2_n143 ) , .A( u2_u3_u2_n98 ) , .ZN( u2_u3_u2_n99 ) );
  NAND2_X1 u2_u3_u2_U58 (.A1( u2_u3_u2_n102 ) , .A2( u2_u3_u2_n106 ) , .ZN( u2_u3_u2_n113 ) );
  NAND2_X1 u2_u3_u2_U59 (.A1( u2_u3_u2_n106 ) , .A2( u2_u3_u2_n107 ) , .ZN( u2_u3_u2_n131 ) );
  AOI21_X1 u2_u3_u2_U6 (.B2( u2_u3_u2_n119 ) , .ZN( u2_u3_u2_n127 ) , .A( u2_u3_u2_n137 ) , .B1( u2_u3_u2_n155 ) );
  NAND2_X1 u2_u3_u2_U60 (.A1( u2_u3_u2_n103 ) , .A2( u2_u3_u2_n107 ) , .ZN( u2_u3_u2_n139 ) );
  NAND2_X1 u2_u3_u2_U61 (.A1( u2_u3_u2_n103 ) , .A2( u2_u3_u2_n105 ) , .ZN( u2_u3_u2_n133 ) );
  NAND2_X1 u2_u3_u2_U62 (.A1( u2_u3_u2_n102 ) , .A2( u2_u3_u2_n103 ) , .ZN( u2_u3_u2_n154 ) );
  NAND2_X1 u2_u3_u2_U63 (.A2( u2_u3_u2_n103 ) , .A1( u2_u3_u2_n104 ) , .ZN( u2_u3_u2_n119 ) );
  NAND2_X1 u2_u3_u2_U64 (.A2( u2_u3_u2_n107 ) , .A1( u2_u3_u2_n108 ) , .ZN( u2_u3_u2_n123 ) );
  NAND2_X1 u2_u3_u2_U65 (.A1( u2_u3_u2_n104 ) , .A2( u2_u3_u2_n108 ) , .ZN( u2_u3_u2_n122 ) );
  INV_X1 u2_u3_u2_U66 (.A( u2_u3_u2_n114 ) , .ZN( u2_u3_u2_n172 ) );
  NAND2_X1 u2_u3_u2_U67 (.A2( u2_u3_u2_n100 ) , .A1( u2_u3_u2_n102 ) , .ZN( u2_u3_u2_n116 ) );
  NAND2_X1 u2_u3_u2_U68 (.A1( u2_u3_u2_n102 ) , .A2( u2_u3_u2_n108 ) , .ZN( u2_u3_u2_n120 ) );
  NAND2_X1 u2_u3_u2_U69 (.A2( u2_u3_u2_n105 ) , .A1( u2_u3_u2_n106 ) , .ZN( u2_u3_u2_n117 ) );
  AOI21_X1 u2_u3_u2_U7 (.ZN( u2_u3_u2_n124 ) , .B1( u2_u3_u2_n131 ) , .B2( u2_u3_u2_n143 ) , .A( u2_u3_u2_n172 ) );
  NOR2_X1 u2_u3_u2_U70 (.A2( u2_u3_X_16 ) , .ZN( u2_u3_u2_n140 ) , .A1( u2_u3_u2_n166 ) );
  NOR2_X1 u2_u3_u2_U71 (.A2( u2_u3_X_13 ) , .A1( u2_u3_X_14 ) , .ZN( u2_u3_u2_n100 ) );
  NOR2_X1 u2_u3_u2_U72 (.A2( u2_u3_X_16 ) , .A1( u2_u3_X_17 ) , .ZN( u2_u3_u2_n138 ) );
  NOR2_X1 u2_u3_u2_U73 (.A2( u2_u3_X_15 ) , .A1( u2_u3_X_18 ) , .ZN( u2_u3_u2_n104 ) );
  NOR2_X1 u2_u3_u2_U74 (.A2( u2_u3_X_14 ) , .ZN( u2_u3_u2_n103 ) , .A1( u2_u3_u2_n174 ) );
  NOR2_X1 u2_u3_u2_U75 (.A2( u2_u3_X_15 ) , .ZN( u2_u3_u2_n102 ) , .A1( u2_u3_u2_n165 ) );
  NOR2_X1 u2_u3_u2_U76 (.A2( u2_u3_X_17 ) , .ZN( u2_u3_u2_n114 ) , .A1( u2_u3_u2_n169 ) );
  AND2_X1 u2_u3_u2_U77 (.A1( u2_u3_X_15 ) , .ZN( u2_u3_u2_n105 ) , .A2( u2_u3_u2_n165 ) );
  AND2_X1 u2_u3_u2_U78 (.A2( u2_u3_X_15 ) , .A1( u2_u3_X_18 ) , .ZN( u2_u3_u2_n107 ) );
  AND2_X1 u2_u3_u2_U79 (.A1( u2_u3_X_14 ) , .ZN( u2_u3_u2_n106 ) , .A2( u2_u3_u2_n174 ) );
  AOI21_X1 u2_u3_u2_U8 (.B2( u2_u3_u2_n120 ) , .B1( u2_u3_u2_n121 ) , .ZN( u2_u3_u2_n126 ) , .A( u2_u3_u2_n167 ) );
  AND2_X1 u2_u3_u2_U80 (.A1( u2_u3_X_13 ) , .A2( u2_u3_X_14 ) , .ZN( u2_u3_u2_n108 ) );
  INV_X1 u2_u3_u2_U81 (.A( u2_u3_X_16 ) , .ZN( u2_u3_u2_n169 ) );
  INV_X1 u2_u3_u2_U82 (.A( u2_u3_X_17 ) , .ZN( u2_u3_u2_n166 ) );
  INV_X1 u2_u3_u2_U83 (.A( u2_u3_X_13 ) , .ZN( u2_u3_u2_n174 ) );
  INV_X1 u2_u3_u2_U84 (.A( u2_u3_X_18 ) , .ZN( u2_u3_u2_n165 ) );
  NAND4_X1 u2_u3_u2_U85 (.ZN( u2_out3_24 ) , .A4( u2_u3_u2_n111 ) , .A3( u2_u3_u2_n112 ) , .A1( u2_u3_u2_n130 ) , .A2( u2_u3_u2_n187 ) );
  AOI221_X1 u2_u3_u2_U86 (.A( u2_u3_u2_n109 ) , .B1( u2_u3_u2_n110 ) , .ZN( u2_u3_u2_n111 ) , .C1( u2_u3_u2_n134 ) , .C2( u2_u3_u2_n170 ) , .B2( u2_u3_u2_n173 ) );
  AOI21_X1 u2_u3_u2_U87 (.ZN( u2_u3_u2_n112 ) , .B2( u2_u3_u2_n156 ) , .A( u2_u3_u2_n164 ) , .B1( u2_u3_u2_n181 ) );
  NAND4_X1 u2_u3_u2_U88 (.ZN( u2_out3_16 ) , .A4( u2_u3_u2_n128 ) , .A3( u2_u3_u2_n129 ) , .A1( u2_u3_u2_n130 ) , .A2( u2_u3_u2_n186 ) );
  AOI22_X1 u2_u3_u2_U89 (.A2( u2_u3_u2_n118 ) , .ZN( u2_u3_u2_n129 ) , .A1( u2_u3_u2_n140 ) , .B1( u2_u3_u2_n157 ) , .B2( u2_u3_u2_n170 ) );
  OAI22_X1 u2_u3_u2_U9 (.ZN( u2_u3_u2_n109 ) , .A2( u2_u3_u2_n113 ) , .B2( u2_u3_u2_n133 ) , .B1( u2_u3_u2_n167 ) , .A1( u2_u3_u2_n168 ) );
  INV_X1 u2_u3_u2_U90 (.A( u2_u3_u2_n163 ) , .ZN( u2_u3_u2_n186 ) );
  NAND4_X1 u2_u3_u2_U91 (.ZN( u2_out3_30 ) , .A4( u2_u3_u2_n147 ) , .A3( u2_u3_u2_n148 ) , .A2( u2_u3_u2_n149 ) , .A1( u2_u3_u2_n187 ) );
  AOI21_X1 u2_u3_u2_U92 (.B2( u2_u3_u2_n138 ) , .ZN( u2_u3_u2_n148 ) , .A( u2_u3_u2_n162 ) , .B1( u2_u3_u2_n182 ) );
  NOR3_X1 u2_u3_u2_U93 (.A3( u2_u3_u2_n144 ) , .A2( u2_u3_u2_n145 ) , .A1( u2_u3_u2_n146 ) , .ZN( u2_u3_u2_n147 ) );
  OR4_X1 u2_u3_u2_U94 (.ZN( u2_out3_6 ) , .A4( u2_u3_u2_n161 ) , .A3( u2_u3_u2_n162 ) , .A2( u2_u3_u2_n163 ) , .A1( u2_u3_u2_n164 ) );
  OR3_X1 u2_u3_u2_U95 (.A2( u2_u3_u2_n159 ) , .A1( u2_u3_u2_n160 ) , .ZN( u2_u3_u2_n161 ) , .A3( u2_u3_u2_n183 ) );
  AOI21_X1 u2_u3_u2_U96 (.B2( u2_u3_u2_n154 ) , .B1( u2_u3_u2_n155 ) , .ZN( u2_u3_u2_n159 ) , .A( u2_u3_u2_n167 ) );
  NAND3_X1 u2_u3_u2_U97 (.A2( u2_u3_u2_n117 ) , .A1( u2_u3_u2_n122 ) , .A3( u2_u3_u2_n123 ) , .ZN( u2_u3_u2_n134 ) );
  NAND3_X1 u2_u3_u2_U98 (.ZN( u2_u3_u2_n110 ) , .A2( u2_u3_u2_n131 ) , .A3( u2_u3_u2_n139 ) , .A1( u2_u3_u2_n154 ) );
  NAND3_X1 u2_u3_u2_U99 (.A2( u2_u3_u2_n100 ) , .ZN( u2_u3_u2_n101 ) , .A1( u2_u3_u2_n104 ) , .A3( u2_u3_u2_n114 ) );
  OAI22_X1 u2_u3_u3_U10 (.B1( u2_u3_u3_n113 ) , .A2( u2_u3_u3_n135 ) , .A1( u2_u3_u3_n150 ) , .B2( u2_u3_u3_n164 ) , .ZN( u2_u3_u3_n98 ) );
  OAI211_X1 u2_u3_u3_U11 (.B( u2_u3_u3_n106 ) , .ZN( u2_u3_u3_n119 ) , .C2( u2_u3_u3_n128 ) , .C1( u2_u3_u3_n167 ) , .A( u2_u3_u3_n181 ) );
  AOI221_X1 u2_u3_u3_U12 (.C1( u2_u3_u3_n105 ) , .ZN( u2_u3_u3_n106 ) , .A( u2_u3_u3_n131 ) , .B2( u2_u3_u3_n132 ) , .C2( u2_u3_u3_n133 ) , .B1( u2_u3_u3_n169 ) );
  INV_X1 u2_u3_u3_U13 (.ZN( u2_u3_u3_n181 ) , .A( u2_u3_u3_n98 ) );
  NAND2_X1 u2_u3_u3_U14 (.ZN( u2_u3_u3_n105 ) , .A2( u2_u3_u3_n130 ) , .A1( u2_u3_u3_n155 ) );
  AOI22_X1 u2_u3_u3_U15 (.B1( u2_u3_u3_n115 ) , .A2( u2_u3_u3_n116 ) , .ZN( u2_u3_u3_n123 ) , .B2( u2_u3_u3_n133 ) , .A1( u2_u3_u3_n169 ) );
  NAND2_X1 u2_u3_u3_U16 (.ZN( u2_u3_u3_n116 ) , .A2( u2_u3_u3_n151 ) , .A1( u2_u3_u3_n182 ) );
  NOR2_X1 u2_u3_u3_U17 (.ZN( u2_u3_u3_n126 ) , .A2( u2_u3_u3_n150 ) , .A1( u2_u3_u3_n164 ) );
  AOI21_X1 u2_u3_u3_U18 (.ZN( u2_u3_u3_n112 ) , .B2( u2_u3_u3_n146 ) , .B1( u2_u3_u3_n155 ) , .A( u2_u3_u3_n167 ) );
  NAND2_X1 u2_u3_u3_U19 (.A1( u2_u3_u3_n135 ) , .ZN( u2_u3_u3_n142 ) , .A2( u2_u3_u3_n164 ) );
  NAND2_X1 u2_u3_u3_U20 (.ZN( u2_u3_u3_n132 ) , .A2( u2_u3_u3_n152 ) , .A1( u2_u3_u3_n156 ) );
  INV_X1 u2_u3_u3_U21 (.A( u2_u3_u3_n133 ) , .ZN( u2_u3_u3_n165 ) );
  AND2_X1 u2_u3_u3_U22 (.A2( u2_u3_u3_n113 ) , .A1( u2_u3_u3_n114 ) , .ZN( u2_u3_u3_n151 ) );
  INV_X1 u2_u3_u3_U23 (.A( u2_u3_u3_n135 ) , .ZN( u2_u3_u3_n170 ) );
  NAND2_X1 u2_u3_u3_U24 (.A1( u2_u3_u3_n107 ) , .A2( u2_u3_u3_n108 ) , .ZN( u2_u3_u3_n140 ) );
  NAND2_X1 u2_u3_u3_U25 (.ZN( u2_u3_u3_n117 ) , .A1( u2_u3_u3_n124 ) , .A2( u2_u3_u3_n148 ) );
  NAND2_X1 u2_u3_u3_U26 (.ZN( u2_u3_u3_n143 ) , .A1( u2_u3_u3_n165 ) , .A2( u2_u3_u3_n167 ) );
  INV_X1 u2_u3_u3_U27 (.A( u2_u3_u3_n130 ) , .ZN( u2_u3_u3_n177 ) );
  INV_X1 u2_u3_u3_U28 (.A( u2_u3_u3_n128 ) , .ZN( u2_u3_u3_n176 ) );
  INV_X1 u2_u3_u3_U29 (.A( u2_u3_u3_n155 ) , .ZN( u2_u3_u3_n174 ) );
  INV_X1 u2_u3_u3_U3 (.A( u2_u3_u3_n140 ) , .ZN( u2_u3_u3_n182 ) );
  INV_X1 u2_u3_u3_U30 (.A( u2_u3_u3_n139 ) , .ZN( u2_u3_u3_n185 ) );
  NOR2_X1 u2_u3_u3_U31 (.ZN( u2_u3_u3_n135 ) , .A2( u2_u3_u3_n141 ) , .A1( u2_u3_u3_n169 ) );
  OAI222_X1 u2_u3_u3_U32 (.C2( u2_u3_u3_n107 ) , .A2( u2_u3_u3_n108 ) , .B1( u2_u3_u3_n135 ) , .ZN( u2_u3_u3_n138 ) , .B2( u2_u3_u3_n146 ) , .C1( u2_u3_u3_n154 ) , .A1( u2_u3_u3_n164 ) );
  NOR4_X1 u2_u3_u3_U33 (.A4( u2_u3_u3_n157 ) , .A3( u2_u3_u3_n158 ) , .A2( u2_u3_u3_n159 ) , .A1( u2_u3_u3_n160 ) , .ZN( u2_u3_u3_n161 ) );
  AOI21_X1 u2_u3_u3_U34 (.B2( u2_u3_u3_n152 ) , .B1( u2_u3_u3_n153 ) , .ZN( u2_u3_u3_n158 ) , .A( u2_u3_u3_n164 ) );
  AOI21_X1 u2_u3_u3_U35 (.A( u2_u3_u3_n149 ) , .B2( u2_u3_u3_n150 ) , .B1( u2_u3_u3_n151 ) , .ZN( u2_u3_u3_n159 ) );
  AOI21_X1 u2_u3_u3_U36 (.A( u2_u3_u3_n154 ) , .B2( u2_u3_u3_n155 ) , .B1( u2_u3_u3_n156 ) , .ZN( u2_u3_u3_n157 ) );
  AOI211_X1 u2_u3_u3_U37 (.ZN( u2_u3_u3_n109 ) , .A( u2_u3_u3_n119 ) , .C2( u2_u3_u3_n129 ) , .B( u2_u3_u3_n138 ) , .C1( u2_u3_u3_n141 ) );
  AOI211_X1 u2_u3_u3_U38 (.B( u2_u3_u3_n119 ) , .A( u2_u3_u3_n120 ) , .C2( u2_u3_u3_n121 ) , .ZN( u2_u3_u3_n122 ) , .C1( u2_u3_u3_n179 ) );
  INV_X1 u2_u3_u3_U39 (.A( u2_u3_u3_n156 ) , .ZN( u2_u3_u3_n179 ) );
  INV_X1 u2_u3_u3_U4 (.A( u2_u3_u3_n129 ) , .ZN( u2_u3_u3_n183 ) );
  OAI22_X1 u2_u3_u3_U40 (.B1( u2_u3_u3_n118 ) , .ZN( u2_u3_u3_n120 ) , .A1( u2_u3_u3_n135 ) , .B2( u2_u3_u3_n154 ) , .A2( u2_u3_u3_n178 ) );
  AND3_X1 u2_u3_u3_U41 (.ZN( u2_u3_u3_n118 ) , .A2( u2_u3_u3_n124 ) , .A1( u2_u3_u3_n144 ) , .A3( u2_u3_u3_n152 ) );
  INV_X1 u2_u3_u3_U42 (.A( u2_u3_u3_n121 ) , .ZN( u2_u3_u3_n164 ) );
  NAND2_X1 u2_u3_u3_U43 (.ZN( u2_u3_u3_n133 ) , .A1( u2_u3_u3_n154 ) , .A2( u2_u3_u3_n164 ) );
  NOR2_X1 u2_u3_u3_U44 (.A1( u2_u3_u3_n113 ) , .ZN( u2_u3_u3_n131 ) , .A2( u2_u3_u3_n154 ) );
  NAND2_X1 u2_u3_u3_U45 (.A1( u2_u3_u3_n103 ) , .ZN( u2_u3_u3_n150 ) , .A2( u2_u3_u3_n99 ) );
  NAND2_X1 u2_u3_u3_U46 (.A2( u2_u3_u3_n102 ) , .ZN( u2_u3_u3_n155 ) , .A1( u2_u3_u3_n97 ) );
  OAI211_X1 u2_u3_u3_U47 (.B( u2_u3_u3_n127 ) , .ZN( u2_u3_u3_n139 ) , .C1( u2_u3_u3_n150 ) , .C2( u2_u3_u3_n154 ) , .A( u2_u3_u3_n184 ) );
  INV_X1 u2_u3_u3_U48 (.A( u2_u3_u3_n125 ) , .ZN( u2_u3_u3_n184 ) );
  AOI221_X1 u2_u3_u3_U49 (.A( u2_u3_u3_n126 ) , .ZN( u2_u3_u3_n127 ) , .C2( u2_u3_u3_n132 ) , .C1( u2_u3_u3_n169 ) , .B2( u2_u3_u3_n170 ) , .B1( u2_u3_u3_n174 ) );
  INV_X1 u2_u3_u3_U5 (.A( u2_u3_u3_n117 ) , .ZN( u2_u3_u3_n178 ) );
  OAI22_X1 u2_u3_u3_U50 (.A1( u2_u3_u3_n124 ) , .ZN( u2_u3_u3_n125 ) , .B2( u2_u3_u3_n145 ) , .A2( u2_u3_u3_n165 ) , .B1( u2_u3_u3_n167 ) );
  INV_X1 u2_u3_u3_U51 (.A( u2_u3_u3_n141 ) , .ZN( u2_u3_u3_n167 ) );
  AOI21_X1 u2_u3_u3_U52 (.B2( u2_u3_u3_n114 ) , .B1( u2_u3_u3_n146 ) , .A( u2_u3_u3_n154 ) , .ZN( u2_u3_u3_n94 ) );
  AOI21_X1 u2_u3_u3_U53 (.ZN( u2_u3_u3_n110 ) , .B2( u2_u3_u3_n142 ) , .B1( u2_u3_u3_n186 ) , .A( u2_u3_u3_n95 ) );
  INV_X1 u2_u3_u3_U54 (.A( u2_u3_u3_n145 ) , .ZN( u2_u3_u3_n186 ) );
  AOI21_X1 u2_u3_u3_U55 (.B1( u2_u3_u3_n124 ) , .A( u2_u3_u3_n149 ) , .B2( u2_u3_u3_n155 ) , .ZN( u2_u3_u3_n95 ) );
  INV_X1 u2_u3_u3_U56 (.A( u2_u3_u3_n149 ) , .ZN( u2_u3_u3_n169 ) );
  NAND2_X1 u2_u3_u3_U57 (.ZN( u2_u3_u3_n124 ) , .A1( u2_u3_u3_n96 ) , .A2( u2_u3_u3_n97 ) );
  NAND2_X1 u2_u3_u3_U58 (.A2( u2_u3_u3_n100 ) , .ZN( u2_u3_u3_n146 ) , .A1( u2_u3_u3_n96 ) );
  NAND2_X1 u2_u3_u3_U59 (.A1( u2_u3_u3_n101 ) , .ZN( u2_u3_u3_n145 ) , .A2( u2_u3_u3_n99 ) );
  AOI221_X1 u2_u3_u3_U6 (.A( u2_u3_u3_n131 ) , .C2( u2_u3_u3_n132 ) , .C1( u2_u3_u3_n133 ) , .ZN( u2_u3_u3_n134 ) , .B1( u2_u3_u3_n143 ) , .B2( u2_u3_u3_n177 ) );
  NAND2_X1 u2_u3_u3_U60 (.A1( u2_u3_u3_n100 ) , .ZN( u2_u3_u3_n156 ) , .A2( u2_u3_u3_n99 ) );
  NAND2_X1 u2_u3_u3_U61 (.A2( u2_u3_u3_n101 ) , .A1( u2_u3_u3_n104 ) , .ZN( u2_u3_u3_n148 ) );
  NAND2_X1 u2_u3_u3_U62 (.A1( u2_u3_u3_n100 ) , .A2( u2_u3_u3_n102 ) , .ZN( u2_u3_u3_n128 ) );
  NAND2_X1 u2_u3_u3_U63 (.A2( u2_u3_u3_n101 ) , .A1( u2_u3_u3_n102 ) , .ZN( u2_u3_u3_n152 ) );
  NAND2_X1 u2_u3_u3_U64 (.A2( u2_u3_u3_n101 ) , .ZN( u2_u3_u3_n114 ) , .A1( u2_u3_u3_n96 ) );
  NAND2_X1 u2_u3_u3_U65 (.ZN( u2_u3_u3_n107 ) , .A1( u2_u3_u3_n97 ) , .A2( u2_u3_u3_n99 ) );
  NAND2_X1 u2_u3_u3_U66 (.A2( u2_u3_u3_n100 ) , .A1( u2_u3_u3_n104 ) , .ZN( u2_u3_u3_n113 ) );
  NAND2_X1 u2_u3_u3_U67 (.A1( u2_u3_u3_n104 ) , .ZN( u2_u3_u3_n153 ) , .A2( u2_u3_u3_n97 ) );
  NAND2_X1 u2_u3_u3_U68 (.A2( u2_u3_u3_n103 ) , .A1( u2_u3_u3_n104 ) , .ZN( u2_u3_u3_n130 ) );
  NAND2_X1 u2_u3_u3_U69 (.A2( u2_u3_u3_n103 ) , .ZN( u2_u3_u3_n144 ) , .A1( u2_u3_u3_n96 ) );
  OAI22_X1 u2_u3_u3_U7 (.B2( u2_u3_u3_n147 ) , .A2( u2_u3_u3_n148 ) , .ZN( u2_u3_u3_n160 ) , .B1( u2_u3_u3_n165 ) , .A1( u2_u3_u3_n168 ) );
  NAND2_X1 u2_u3_u3_U70 (.A1( u2_u3_u3_n102 ) , .A2( u2_u3_u3_n103 ) , .ZN( u2_u3_u3_n108 ) );
  NOR2_X1 u2_u3_u3_U71 (.A2( u2_u3_X_19 ) , .A1( u2_u3_X_20 ) , .ZN( u2_u3_u3_n99 ) );
  NOR2_X1 u2_u3_u3_U72 (.A2( u2_u3_X_21 ) , .A1( u2_u3_X_24 ) , .ZN( u2_u3_u3_n103 ) );
  NOR2_X1 u2_u3_u3_U73 (.A2( u2_u3_X_24 ) , .A1( u2_u3_u3_n171 ) , .ZN( u2_u3_u3_n97 ) );
  NOR2_X1 u2_u3_u3_U74 (.A2( u2_u3_X_23 ) , .ZN( u2_u3_u3_n141 ) , .A1( u2_u3_u3_n166 ) );
  NOR2_X1 u2_u3_u3_U75 (.A2( u2_u3_X_19 ) , .A1( u2_u3_u3_n172 ) , .ZN( u2_u3_u3_n96 ) );
  NAND2_X1 u2_u3_u3_U76 (.A1( u2_u3_X_22 ) , .A2( u2_u3_X_23 ) , .ZN( u2_u3_u3_n154 ) );
  NAND2_X1 u2_u3_u3_U77 (.A1( u2_u3_X_23 ) , .ZN( u2_u3_u3_n149 ) , .A2( u2_u3_u3_n166 ) );
  NOR2_X1 u2_u3_u3_U78 (.A2( u2_u3_X_22 ) , .A1( u2_u3_X_23 ) , .ZN( u2_u3_u3_n121 ) );
  AND2_X1 u2_u3_u3_U79 (.A1( u2_u3_X_24 ) , .ZN( u2_u3_u3_n101 ) , .A2( u2_u3_u3_n171 ) );
  AND3_X1 u2_u3_u3_U8 (.A3( u2_u3_u3_n144 ) , .A2( u2_u3_u3_n145 ) , .A1( u2_u3_u3_n146 ) , .ZN( u2_u3_u3_n147 ) );
  AND2_X1 u2_u3_u3_U80 (.A1( u2_u3_X_19 ) , .ZN( u2_u3_u3_n102 ) , .A2( u2_u3_u3_n172 ) );
  AND2_X1 u2_u3_u3_U81 (.A1( u2_u3_X_21 ) , .A2( u2_u3_X_24 ) , .ZN( u2_u3_u3_n100 ) );
  AND2_X1 u2_u3_u3_U82 (.A2( u2_u3_X_19 ) , .A1( u2_u3_X_20 ) , .ZN( u2_u3_u3_n104 ) );
  INV_X1 u2_u3_u3_U83 (.A( u2_u3_X_22 ) , .ZN( u2_u3_u3_n166 ) );
  INV_X1 u2_u3_u3_U84 (.A( u2_u3_X_21 ) , .ZN( u2_u3_u3_n171 ) );
  INV_X1 u2_u3_u3_U85 (.A( u2_u3_X_20 ) , .ZN( u2_u3_u3_n172 ) );
  NAND4_X1 u2_u3_u3_U86 (.ZN( u2_out3_26 ) , .A4( u2_u3_u3_n109 ) , .A3( u2_u3_u3_n110 ) , .A2( u2_u3_u3_n111 ) , .A1( u2_u3_u3_n173 ) );
  INV_X1 u2_u3_u3_U87 (.ZN( u2_u3_u3_n173 ) , .A( u2_u3_u3_n94 ) );
  OAI21_X1 u2_u3_u3_U88 (.ZN( u2_u3_u3_n111 ) , .B2( u2_u3_u3_n117 ) , .A( u2_u3_u3_n133 ) , .B1( u2_u3_u3_n176 ) );
  NAND4_X1 u2_u3_u3_U89 (.ZN( u2_out3_20 ) , .A4( u2_u3_u3_n122 ) , .A3( u2_u3_u3_n123 ) , .A1( u2_u3_u3_n175 ) , .A2( u2_u3_u3_n180 ) );
  INV_X1 u2_u3_u3_U9 (.A( u2_u3_u3_n143 ) , .ZN( u2_u3_u3_n168 ) );
  INV_X1 u2_u3_u3_U90 (.A( u2_u3_u3_n126 ) , .ZN( u2_u3_u3_n180 ) );
  INV_X1 u2_u3_u3_U91 (.A( u2_u3_u3_n112 ) , .ZN( u2_u3_u3_n175 ) );
  NAND4_X1 u2_u3_u3_U92 (.ZN( u2_out3_1 ) , .A4( u2_u3_u3_n161 ) , .A3( u2_u3_u3_n162 ) , .A2( u2_u3_u3_n163 ) , .A1( u2_u3_u3_n185 ) );
  NAND2_X1 u2_u3_u3_U93 (.ZN( u2_u3_u3_n163 ) , .A2( u2_u3_u3_n170 ) , .A1( u2_u3_u3_n176 ) );
  AOI22_X1 u2_u3_u3_U94 (.B2( u2_u3_u3_n140 ) , .B1( u2_u3_u3_n141 ) , .A2( u2_u3_u3_n142 ) , .ZN( u2_u3_u3_n162 ) , .A1( u2_u3_u3_n177 ) );
  OAI222_X1 u2_u3_u3_U95 (.C1( u2_u3_u3_n128 ) , .ZN( u2_u3_u3_n137 ) , .B1( u2_u3_u3_n148 ) , .A2( u2_u3_u3_n150 ) , .B2( u2_u3_u3_n154 ) , .C2( u2_u3_u3_n164 ) , .A1( u2_u3_u3_n167 ) );
  OR4_X1 u2_u3_u3_U96 (.ZN( u2_out3_10 ) , .A4( u2_u3_u3_n136 ) , .A3( u2_u3_u3_n137 ) , .A1( u2_u3_u3_n138 ) , .A2( u2_u3_u3_n139 ) );
  OAI221_X1 u2_u3_u3_U97 (.A( u2_u3_u3_n134 ) , .B2( u2_u3_u3_n135 ) , .ZN( u2_u3_u3_n136 ) , .C1( u2_u3_u3_n149 ) , .B1( u2_u3_u3_n151 ) , .C2( u2_u3_u3_n183 ) );
  NAND3_X1 u2_u3_u3_U98 (.A1( u2_u3_u3_n114 ) , .ZN( u2_u3_u3_n115 ) , .A2( u2_u3_u3_n145 ) , .A3( u2_u3_u3_n153 ) );
  NAND3_X1 u2_u3_u3_U99 (.ZN( u2_u3_u3_n129 ) , .A2( u2_u3_u3_n144 ) , .A1( u2_u3_u3_n153 ) , .A3( u2_u3_u3_n182 ) );
  OAI22_X1 u2_u3_u4_U10 (.B2( u2_u3_u4_n135 ) , .ZN( u2_u3_u4_n137 ) , .B1( u2_u3_u4_n153 ) , .A1( u2_u3_u4_n155 ) , .A2( u2_u3_u4_n171 ) );
  AND3_X1 u2_u3_u4_U11 (.A2( u2_u3_u4_n134 ) , .ZN( u2_u3_u4_n135 ) , .A3( u2_u3_u4_n145 ) , .A1( u2_u3_u4_n157 ) );
  OR3_X1 u2_u3_u4_U12 (.A3( u2_u3_u4_n114 ) , .A2( u2_u3_u4_n115 ) , .A1( u2_u3_u4_n116 ) , .ZN( u2_u3_u4_n136 ) );
  AOI21_X1 u2_u3_u4_U13 (.A( u2_u3_u4_n113 ) , .ZN( u2_u3_u4_n116 ) , .B2( u2_u3_u4_n173 ) , .B1( u2_u3_u4_n174 ) );
  AOI21_X1 u2_u3_u4_U14 (.ZN( u2_u3_u4_n115 ) , .B2( u2_u3_u4_n145 ) , .B1( u2_u3_u4_n146 ) , .A( u2_u3_u4_n156 ) );
  OAI22_X1 u2_u3_u4_U15 (.ZN( u2_u3_u4_n114 ) , .A2( u2_u3_u4_n121 ) , .B1( u2_u3_u4_n160 ) , .B2( u2_u3_u4_n170 ) , .A1( u2_u3_u4_n171 ) );
  NAND2_X1 u2_u3_u4_U16 (.ZN( u2_u3_u4_n132 ) , .A2( u2_u3_u4_n170 ) , .A1( u2_u3_u4_n173 ) );
  AOI21_X1 u2_u3_u4_U17 (.B2( u2_u3_u4_n160 ) , .B1( u2_u3_u4_n161 ) , .ZN( u2_u3_u4_n162 ) , .A( u2_u3_u4_n170 ) );
  AOI21_X1 u2_u3_u4_U18 (.ZN( u2_u3_u4_n107 ) , .B2( u2_u3_u4_n143 ) , .A( u2_u3_u4_n174 ) , .B1( u2_u3_u4_n184 ) );
  AOI21_X1 u2_u3_u4_U19 (.B2( u2_u3_u4_n158 ) , .B1( u2_u3_u4_n159 ) , .ZN( u2_u3_u4_n163 ) , .A( u2_u3_u4_n174 ) );
  AOI21_X1 u2_u3_u4_U20 (.A( u2_u3_u4_n153 ) , .B2( u2_u3_u4_n154 ) , .B1( u2_u3_u4_n155 ) , .ZN( u2_u3_u4_n165 ) );
  AOI21_X1 u2_u3_u4_U21 (.A( u2_u3_u4_n156 ) , .B2( u2_u3_u4_n157 ) , .ZN( u2_u3_u4_n164 ) , .B1( u2_u3_u4_n184 ) );
  INV_X1 u2_u3_u4_U22 (.A( u2_u3_u4_n138 ) , .ZN( u2_u3_u4_n170 ) );
  AND2_X1 u2_u3_u4_U23 (.A2( u2_u3_u4_n120 ) , .ZN( u2_u3_u4_n155 ) , .A1( u2_u3_u4_n160 ) );
  INV_X1 u2_u3_u4_U24 (.A( u2_u3_u4_n156 ) , .ZN( u2_u3_u4_n175 ) );
  NAND2_X1 u2_u3_u4_U25 (.A2( u2_u3_u4_n118 ) , .ZN( u2_u3_u4_n131 ) , .A1( u2_u3_u4_n147 ) );
  NAND2_X1 u2_u3_u4_U26 (.A1( u2_u3_u4_n119 ) , .A2( u2_u3_u4_n120 ) , .ZN( u2_u3_u4_n130 ) );
  NAND2_X1 u2_u3_u4_U27 (.ZN( u2_u3_u4_n117 ) , .A2( u2_u3_u4_n118 ) , .A1( u2_u3_u4_n148 ) );
  NAND2_X1 u2_u3_u4_U28 (.ZN( u2_u3_u4_n129 ) , .A1( u2_u3_u4_n134 ) , .A2( u2_u3_u4_n148 ) );
  AND3_X1 u2_u3_u4_U29 (.A1( u2_u3_u4_n119 ) , .A2( u2_u3_u4_n143 ) , .A3( u2_u3_u4_n154 ) , .ZN( u2_u3_u4_n161 ) );
  NOR2_X1 u2_u3_u4_U3 (.ZN( u2_u3_u4_n121 ) , .A1( u2_u3_u4_n181 ) , .A2( u2_u3_u4_n182 ) );
  AND2_X1 u2_u3_u4_U30 (.A1( u2_u3_u4_n145 ) , .A2( u2_u3_u4_n147 ) , .ZN( u2_u3_u4_n159 ) );
  INV_X1 u2_u3_u4_U31 (.A( u2_u3_u4_n158 ) , .ZN( u2_u3_u4_n182 ) );
  INV_X1 u2_u3_u4_U32 (.ZN( u2_u3_u4_n181 ) , .A( u2_u3_u4_n96 ) );
  INV_X1 u2_u3_u4_U33 (.A( u2_u3_u4_n144 ) , .ZN( u2_u3_u4_n179 ) );
  INV_X1 u2_u3_u4_U34 (.A( u2_u3_u4_n157 ) , .ZN( u2_u3_u4_n178 ) );
  NAND2_X1 u2_u3_u4_U35 (.A2( u2_u3_u4_n154 ) , .A1( u2_u3_u4_n96 ) , .ZN( u2_u3_u4_n97 ) );
  INV_X1 u2_u3_u4_U36 (.ZN( u2_u3_u4_n186 ) , .A( u2_u3_u4_n95 ) );
  OAI221_X1 u2_u3_u4_U37 (.C1( u2_u3_u4_n134 ) , .B1( u2_u3_u4_n158 ) , .B2( u2_u3_u4_n171 ) , .C2( u2_u3_u4_n173 ) , .A( u2_u3_u4_n94 ) , .ZN( u2_u3_u4_n95 ) );
  AOI222_X1 u2_u3_u4_U38 (.B2( u2_u3_u4_n132 ) , .A1( u2_u3_u4_n138 ) , .C2( u2_u3_u4_n175 ) , .A2( u2_u3_u4_n179 ) , .C1( u2_u3_u4_n181 ) , .B1( u2_u3_u4_n185 ) , .ZN( u2_u3_u4_n94 ) );
  INV_X1 u2_u3_u4_U39 (.A( u2_u3_u4_n113 ) , .ZN( u2_u3_u4_n185 ) );
  INV_X1 u2_u3_u4_U4 (.A( u2_u3_u4_n117 ) , .ZN( u2_u3_u4_n184 ) );
  INV_X1 u2_u3_u4_U40 (.A( u2_u3_u4_n143 ) , .ZN( u2_u3_u4_n183 ) );
  NOR2_X1 u2_u3_u4_U41 (.ZN( u2_u3_u4_n138 ) , .A1( u2_u3_u4_n168 ) , .A2( u2_u3_u4_n169 ) );
  NOR2_X1 u2_u3_u4_U42 (.A1( u2_u3_u4_n150 ) , .A2( u2_u3_u4_n152 ) , .ZN( u2_u3_u4_n153 ) );
  NOR2_X1 u2_u3_u4_U43 (.A2( u2_u3_u4_n128 ) , .A1( u2_u3_u4_n138 ) , .ZN( u2_u3_u4_n156 ) );
  AOI22_X1 u2_u3_u4_U44 (.B2( u2_u3_u4_n122 ) , .A1( u2_u3_u4_n123 ) , .ZN( u2_u3_u4_n124 ) , .B1( u2_u3_u4_n128 ) , .A2( u2_u3_u4_n172 ) );
  INV_X1 u2_u3_u4_U45 (.A( u2_u3_u4_n153 ) , .ZN( u2_u3_u4_n172 ) );
  NAND2_X1 u2_u3_u4_U46 (.A2( u2_u3_u4_n120 ) , .ZN( u2_u3_u4_n123 ) , .A1( u2_u3_u4_n161 ) );
  AOI22_X1 u2_u3_u4_U47 (.B2( u2_u3_u4_n132 ) , .A2( u2_u3_u4_n133 ) , .ZN( u2_u3_u4_n140 ) , .A1( u2_u3_u4_n150 ) , .B1( u2_u3_u4_n179 ) );
  NAND2_X1 u2_u3_u4_U48 (.ZN( u2_u3_u4_n133 ) , .A2( u2_u3_u4_n146 ) , .A1( u2_u3_u4_n154 ) );
  NAND2_X1 u2_u3_u4_U49 (.A1( u2_u3_u4_n103 ) , .ZN( u2_u3_u4_n154 ) , .A2( u2_u3_u4_n98 ) );
  NOR4_X1 u2_u3_u4_U5 (.A4( u2_u3_u4_n106 ) , .A3( u2_u3_u4_n107 ) , .A2( u2_u3_u4_n108 ) , .A1( u2_u3_u4_n109 ) , .ZN( u2_u3_u4_n110 ) );
  NAND2_X1 u2_u3_u4_U50 (.A1( u2_u3_u4_n101 ) , .ZN( u2_u3_u4_n158 ) , .A2( u2_u3_u4_n99 ) );
  AOI21_X1 u2_u3_u4_U51 (.ZN( u2_u3_u4_n127 ) , .A( u2_u3_u4_n136 ) , .B2( u2_u3_u4_n150 ) , .B1( u2_u3_u4_n180 ) );
  INV_X1 u2_u3_u4_U52 (.A( u2_u3_u4_n160 ) , .ZN( u2_u3_u4_n180 ) );
  NAND2_X1 u2_u3_u4_U53 (.A2( u2_u3_u4_n104 ) , .A1( u2_u3_u4_n105 ) , .ZN( u2_u3_u4_n146 ) );
  NAND2_X1 u2_u3_u4_U54 (.A2( u2_u3_u4_n101 ) , .A1( u2_u3_u4_n102 ) , .ZN( u2_u3_u4_n160 ) );
  NAND2_X1 u2_u3_u4_U55 (.ZN( u2_u3_u4_n134 ) , .A1( u2_u3_u4_n98 ) , .A2( u2_u3_u4_n99 ) );
  NAND2_X1 u2_u3_u4_U56 (.A1( u2_u3_u4_n103 ) , .A2( u2_u3_u4_n104 ) , .ZN( u2_u3_u4_n143 ) );
  NAND2_X1 u2_u3_u4_U57 (.A2( u2_u3_u4_n105 ) , .ZN( u2_u3_u4_n145 ) , .A1( u2_u3_u4_n98 ) );
  NAND2_X1 u2_u3_u4_U58 (.A1( u2_u3_u4_n100 ) , .A2( u2_u3_u4_n105 ) , .ZN( u2_u3_u4_n120 ) );
  NAND2_X1 u2_u3_u4_U59 (.A1( u2_u3_u4_n102 ) , .A2( u2_u3_u4_n104 ) , .ZN( u2_u3_u4_n148 ) );
  AOI21_X1 u2_u3_u4_U6 (.ZN( u2_u3_u4_n106 ) , .B2( u2_u3_u4_n146 ) , .B1( u2_u3_u4_n158 ) , .A( u2_u3_u4_n170 ) );
  NAND2_X1 u2_u3_u4_U60 (.A2( u2_u3_u4_n100 ) , .A1( u2_u3_u4_n103 ) , .ZN( u2_u3_u4_n157 ) );
  INV_X1 u2_u3_u4_U61 (.A( u2_u3_u4_n150 ) , .ZN( u2_u3_u4_n173 ) );
  INV_X1 u2_u3_u4_U62 (.A( u2_u3_u4_n152 ) , .ZN( u2_u3_u4_n171 ) );
  NAND2_X1 u2_u3_u4_U63 (.A1( u2_u3_u4_n100 ) , .ZN( u2_u3_u4_n118 ) , .A2( u2_u3_u4_n99 ) );
  NAND2_X1 u2_u3_u4_U64 (.A2( u2_u3_u4_n100 ) , .A1( u2_u3_u4_n102 ) , .ZN( u2_u3_u4_n144 ) );
  NAND2_X1 u2_u3_u4_U65 (.A2( u2_u3_u4_n101 ) , .A1( u2_u3_u4_n105 ) , .ZN( u2_u3_u4_n96 ) );
  INV_X1 u2_u3_u4_U66 (.A( u2_u3_u4_n128 ) , .ZN( u2_u3_u4_n174 ) );
  NAND2_X1 u2_u3_u4_U67 (.A2( u2_u3_u4_n102 ) , .ZN( u2_u3_u4_n119 ) , .A1( u2_u3_u4_n98 ) );
  NAND2_X1 u2_u3_u4_U68 (.A2( u2_u3_u4_n101 ) , .A1( u2_u3_u4_n103 ) , .ZN( u2_u3_u4_n147 ) );
  NAND2_X1 u2_u3_u4_U69 (.A2( u2_u3_u4_n104 ) , .ZN( u2_u3_u4_n113 ) , .A1( u2_u3_u4_n99 ) );
  AOI21_X1 u2_u3_u4_U7 (.ZN( u2_u3_u4_n109 ) , .A( u2_u3_u4_n153 ) , .B1( u2_u3_u4_n159 ) , .B2( u2_u3_u4_n184 ) );
  NOR2_X1 u2_u3_u4_U70 (.A2( u2_u3_X_28 ) , .ZN( u2_u3_u4_n150 ) , .A1( u2_u3_u4_n168 ) );
  NOR2_X1 u2_u3_u4_U71 (.A2( u2_u3_X_29 ) , .ZN( u2_u3_u4_n152 ) , .A1( u2_u3_u4_n169 ) );
  NOR2_X1 u2_u3_u4_U72 (.A2( u2_u3_X_30 ) , .ZN( u2_u3_u4_n105 ) , .A1( u2_u3_u4_n176 ) );
  NOR2_X1 u2_u3_u4_U73 (.A2( u2_u3_X_26 ) , .ZN( u2_u3_u4_n100 ) , .A1( u2_u3_u4_n177 ) );
  NOR2_X1 u2_u3_u4_U74 (.A2( u2_u3_X_28 ) , .A1( u2_u3_X_29 ) , .ZN( u2_u3_u4_n128 ) );
  NOR2_X1 u2_u3_u4_U75 (.A2( u2_u3_X_27 ) , .A1( u2_u3_X_30 ) , .ZN( u2_u3_u4_n102 ) );
  NOR2_X1 u2_u3_u4_U76 (.A2( u2_u3_X_25 ) , .A1( u2_u3_X_26 ) , .ZN( u2_u3_u4_n98 ) );
  AND2_X1 u2_u3_u4_U77 (.A2( u2_u3_X_25 ) , .A1( u2_u3_X_26 ) , .ZN( u2_u3_u4_n104 ) );
  AND2_X1 u2_u3_u4_U78 (.A1( u2_u3_X_30 ) , .A2( u2_u3_u4_n176 ) , .ZN( u2_u3_u4_n99 ) );
  AND2_X1 u2_u3_u4_U79 (.A1( u2_u3_X_26 ) , .ZN( u2_u3_u4_n101 ) , .A2( u2_u3_u4_n177 ) );
  AOI21_X1 u2_u3_u4_U8 (.ZN( u2_u3_u4_n108 ) , .B2( u2_u3_u4_n134 ) , .B1( u2_u3_u4_n155 ) , .A( u2_u3_u4_n156 ) );
  AND2_X1 u2_u3_u4_U80 (.A1( u2_u3_X_27 ) , .A2( u2_u3_X_30 ) , .ZN( u2_u3_u4_n103 ) );
  INV_X1 u2_u3_u4_U81 (.A( u2_u3_X_28 ) , .ZN( u2_u3_u4_n169 ) );
  INV_X1 u2_u3_u4_U82 (.A( u2_u3_X_29 ) , .ZN( u2_u3_u4_n168 ) );
  INV_X1 u2_u3_u4_U83 (.A( u2_u3_X_25 ) , .ZN( u2_u3_u4_n177 ) );
  INV_X1 u2_u3_u4_U84 (.A( u2_u3_X_27 ) , .ZN( u2_u3_u4_n176 ) );
  NAND4_X1 u2_u3_u4_U85 (.ZN( u2_out3_25 ) , .A4( u2_u3_u4_n139 ) , .A3( u2_u3_u4_n140 ) , .A2( u2_u3_u4_n141 ) , .A1( u2_u3_u4_n142 ) );
  OAI21_X1 u2_u3_u4_U86 (.A( u2_u3_u4_n128 ) , .B2( u2_u3_u4_n129 ) , .B1( u2_u3_u4_n130 ) , .ZN( u2_u3_u4_n142 ) );
  OAI21_X1 u2_u3_u4_U87 (.B2( u2_u3_u4_n131 ) , .ZN( u2_u3_u4_n141 ) , .A( u2_u3_u4_n175 ) , .B1( u2_u3_u4_n183 ) );
  NAND4_X1 u2_u3_u4_U88 (.ZN( u2_out3_14 ) , .A4( u2_u3_u4_n124 ) , .A3( u2_u3_u4_n125 ) , .A2( u2_u3_u4_n126 ) , .A1( u2_u3_u4_n127 ) );
  AOI22_X1 u2_u3_u4_U89 (.B2( u2_u3_u4_n117 ) , .ZN( u2_u3_u4_n126 ) , .A1( u2_u3_u4_n129 ) , .B1( u2_u3_u4_n152 ) , .A2( u2_u3_u4_n175 ) );
  AOI211_X1 u2_u3_u4_U9 (.B( u2_u3_u4_n136 ) , .A( u2_u3_u4_n137 ) , .C2( u2_u3_u4_n138 ) , .ZN( u2_u3_u4_n139 ) , .C1( u2_u3_u4_n182 ) );
  AOI22_X1 u2_u3_u4_U90 (.ZN( u2_u3_u4_n125 ) , .B2( u2_u3_u4_n131 ) , .A2( u2_u3_u4_n132 ) , .B1( u2_u3_u4_n138 ) , .A1( u2_u3_u4_n178 ) );
  NAND4_X1 u2_u3_u4_U91 (.ZN( u2_out3_8 ) , .A4( u2_u3_u4_n110 ) , .A3( u2_u3_u4_n111 ) , .A2( u2_u3_u4_n112 ) , .A1( u2_u3_u4_n186 ) );
  NAND2_X1 u2_u3_u4_U92 (.ZN( u2_u3_u4_n112 ) , .A2( u2_u3_u4_n130 ) , .A1( u2_u3_u4_n150 ) );
  AOI22_X1 u2_u3_u4_U93 (.ZN( u2_u3_u4_n111 ) , .B2( u2_u3_u4_n132 ) , .A1( u2_u3_u4_n152 ) , .B1( u2_u3_u4_n178 ) , .A2( u2_u3_u4_n97 ) );
  AOI22_X1 u2_u3_u4_U94 (.B2( u2_u3_u4_n149 ) , .B1( u2_u3_u4_n150 ) , .A2( u2_u3_u4_n151 ) , .A1( u2_u3_u4_n152 ) , .ZN( u2_u3_u4_n167 ) );
  NOR4_X1 u2_u3_u4_U95 (.A4( u2_u3_u4_n162 ) , .A3( u2_u3_u4_n163 ) , .A2( u2_u3_u4_n164 ) , .A1( u2_u3_u4_n165 ) , .ZN( u2_u3_u4_n166 ) );
  NAND3_X1 u2_u3_u4_U96 (.ZN( u2_out3_3 ) , .A3( u2_u3_u4_n166 ) , .A1( u2_u3_u4_n167 ) , .A2( u2_u3_u4_n186 ) );
  NAND3_X1 u2_u3_u4_U97 (.A3( u2_u3_u4_n146 ) , .A2( u2_u3_u4_n147 ) , .A1( u2_u3_u4_n148 ) , .ZN( u2_u3_u4_n149 ) );
  NAND3_X1 u2_u3_u4_U98 (.A3( u2_u3_u4_n143 ) , .A2( u2_u3_u4_n144 ) , .A1( u2_u3_u4_n145 ) , .ZN( u2_u3_u4_n151 ) );
  NAND3_X1 u2_u3_u4_U99 (.A3( u2_u3_u4_n121 ) , .ZN( u2_u3_u4_n122 ) , .A2( u2_u3_u4_n144 ) , .A1( u2_u3_u4_n154 ) );
  INV_X1 u2_u3_u5_U10 (.A( u2_u3_u5_n121 ) , .ZN( u2_u3_u5_n177 ) );
  NOR3_X1 u2_u3_u5_U100 (.A3( u2_u3_u5_n141 ) , .A1( u2_u3_u5_n142 ) , .ZN( u2_u3_u5_n143 ) , .A2( u2_u3_u5_n191 ) );
  NAND4_X1 u2_u3_u5_U101 (.ZN( u2_out3_4 ) , .A4( u2_u3_u5_n112 ) , .A2( u2_u3_u5_n113 ) , .A1( u2_u3_u5_n114 ) , .A3( u2_u3_u5_n195 ) );
  AOI211_X1 u2_u3_u5_U102 (.A( u2_u3_u5_n110 ) , .C1( u2_u3_u5_n111 ) , .ZN( u2_u3_u5_n112 ) , .B( u2_u3_u5_n118 ) , .C2( u2_u3_u5_n177 ) );
  AOI222_X1 u2_u3_u5_U103 (.ZN( u2_u3_u5_n113 ) , .A1( u2_u3_u5_n131 ) , .C1( u2_u3_u5_n148 ) , .B2( u2_u3_u5_n174 ) , .C2( u2_u3_u5_n178 ) , .A2( u2_u3_u5_n179 ) , .B1( u2_u3_u5_n99 ) );
  NAND3_X1 u2_u3_u5_U104 (.A2( u2_u3_u5_n154 ) , .A3( u2_u3_u5_n158 ) , .A1( u2_u3_u5_n161 ) , .ZN( u2_u3_u5_n99 ) );
  NOR2_X1 u2_u3_u5_U11 (.ZN( u2_u3_u5_n160 ) , .A2( u2_u3_u5_n173 ) , .A1( u2_u3_u5_n177 ) );
  INV_X1 u2_u3_u5_U12 (.A( u2_u3_u5_n150 ) , .ZN( u2_u3_u5_n174 ) );
  AOI21_X1 u2_u3_u5_U13 (.A( u2_u3_u5_n160 ) , .B2( u2_u3_u5_n161 ) , .ZN( u2_u3_u5_n162 ) , .B1( u2_u3_u5_n192 ) );
  INV_X1 u2_u3_u5_U14 (.A( u2_u3_u5_n159 ) , .ZN( u2_u3_u5_n192 ) );
  AOI21_X1 u2_u3_u5_U15 (.A( u2_u3_u5_n156 ) , .B2( u2_u3_u5_n157 ) , .B1( u2_u3_u5_n158 ) , .ZN( u2_u3_u5_n163 ) );
  AOI21_X1 u2_u3_u5_U16 (.B2( u2_u3_u5_n139 ) , .B1( u2_u3_u5_n140 ) , .ZN( u2_u3_u5_n141 ) , .A( u2_u3_u5_n150 ) );
  OAI21_X1 u2_u3_u5_U17 (.A( u2_u3_u5_n133 ) , .B2( u2_u3_u5_n134 ) , .B1( u2_u3_u5_n135 ) , .ZN( u2_u3_u5_n142 ) );
  OAI21_X1 u2_u3_u5_U18 (.ZN( u2_u3_u5_n133 ) , .B2( u2_u3_u5_n147 ) , .A( u2_u3_u5_n173 ) , .B1( u2_u3_u5_n188 ) );
  NAND2_X1 u2_u3_u5_U19 (.A2( u2_u3_u5_n119 ) , .A1( u2_u3_u5_n123 ) , .ZN( u2_u3_u5_n137 ) );
  INV_X1 u2_u3_u5_U20 (.A( u2_u3_u5_n155 ) , .ZN( u2_u3_u5_n194 ) );
  NAND2_X1 u2_u3_u5_U21 (.A1( u2_u3_u5_n121 ) , .ZN( u2_u3_u5_n132 ) , .A2( u2_u3_u5_n172 ) );
  NAND2_X1 u2_u3_u5_U22 (.A2( u2_u3_u5_n122 ) , .ZN( u2_u3_u5_n136 ) , .A1( u2_u3_u5_n154 ) );
  NAND2_X1 u2_u3_u5_U23 (.A2( u2_u3_u5_n119 ) , .A1( u2_u3_u5_n120 ) , .ZN( u2_u3_u5_n159 ) );
  INV_X1 u2_u3_u5_U24 (.A( u2_u3_u5_n156 ) , .ZN( u2_u3_u5_n175 ) );
  INV_X1 u2_u3_u5_U25 (.A( u2_u3_u5_n158 ) , .ZN( u2_u3_u5_n188 ) );
  INV_X1 u2_u3_u5_U26 (.A( u2_u3_u5_n152 ) , .ZN( u2_u3_u5_n179 ) );
  INV_X1 u2_u3_u5_U27 (.A( u2_u3_u5_n140 ) , .ZN( u2_u3_u5_n182 ) );
  INV_X1 u2_u3_u5_U28 (.A( u2_u3_u5_n151 ) , .ZN( u2_u3_u5_n183 ) );
  INV_X1 u2_u3_u5_U29 (.A( u2_u3_u5_n123 ) , .ZN( u2_u3_u5_n185 ) );
  NOR2_X1 u2_u3_u5_U3 (.ZN( u2_u3_u5_n134 ) , .A1( u2_u3_u5_n183 ) , .A2( u2_u3_u5_n190 ) );
  INV_X1 u2_u3_u5_U30 (.A( u2_u3_u5_n161 ) , .ZN( u2_u3_u5_n184 ) );
  INV_X1 u2_u3_u5_U31 (.A( u2_u3_u5_n139 ) , .ZN( u2_u3_u5_n189 ) );
  INV_X1 u2_u3_u5_U32 (.A( u2_u3_u5_n157 ) , .ZN( u2_u3_u5_n190 ) );
  INV_X1 u2_u3_u5_U33 (.A( u2_u3_u5_n120 ) , .ZN( u2_u3_u5_n193 ) );
  NAND2_X1 u2_u3_u5_U34 (.ZN( u2_u3_u5_n111 ) , .A1( u2_u3_u5_n140 ) , .A2( u2_u3_u5_n155 ) );
  INV_X1 u2_u3_u5_U35 (.A( u2_u3_u5_n117 ) , .ZN( u2_u3_u5_n196 ) );
  OAI221_X1 u2_u3_u5_U36 (.A( u2_u3_u5_n116 ) , .ZN( u2_u3_u5_n117 ) , .B2( u2_u3_u5_n119 ) , .C1( u2_u3_u5_n153 ) , .C2( u2_u3_u5_n158 ) , .B1( u2_u3_u5_n172 ) );
  AOI222_X1 u2_u3_u5_U37 (.ZN( u2_u3_u5_n116 ) , .B2( u2_u3_u5_n145 ) , .C1( u2_u3_u5_n148 ) , .A2( u2_u3_u5_n174 ) , .C2( u2_u3_u5_n177 ) , .B1( u2_u3_u5_n187 ) , .A1( u2_u3_u5_n193 ) );
  INV_X1 u2_u3_u5_U38 (.A( u2_u3_u5_n115 ) , .ZN( u2_u3_u5_n187 ) );
  NOR2_X1 u2_u3_u5_U39 (.ZN( u2_u3_u5_n100 ) , .A1( u2_u3_u5_n170 ) , .A2( u2_u3_u5_n180 ) );
  INV_X1 u2_u3_u5_U4 (.A( u2_u3_u5_n138 ) , .ZN( u2_u3_u5_n191 ) );
  AOI22_X1 u2_u3_u5_U40 (.B2( u2_u3_u5_n131 ) , .A2( u2_u3_u5_n146 ) , .ZN( u2_u3_u5_n169 ) , .B1( u2_u3_u5_n174 ) , .A1( u2_u3_u5_n185 ) );
  NOR2_X1 u2_u3_u5_U41 (.A1( u2_u3_u5_n146 ) , .ZN( u2_u3_u5_n150 ) , .A2( u2_u3_u5_n173 ) );
  AOI21_X1 u2_u3_u5_U42 (.A( u2_u3_u5_n118 ) , .B2( u2_u3_u5_n145 ) , .ZN( u2_u3_u5_n168 ) , .B1( u2_u3_u5_n186 ) );
  INV_X1 u2_u3_u5_U43 (.A( u2_u3_u5_n122 ) , .ZN( u2_u3_u5_n186 ) );
  NOR2_X1 u2_u3_u5_U44 (.A1( u2_u3_u5_n146 ) , .ZN( u2_u3_u5_n152 ) , .A2( u2_u3_u5_n176 ) );
  NOR2_X1 u2_u3_u5_U45 (.A1( u2_u3_u5_n115 ) , .ZN( u2_u3_u5_n118 ) , .A2( u2_u3_u5_n153 ) );
  NOR2_X1 u2_u3_u5_U46 (.A2( u2_u3_u5_n145 ) , .ZN( u2_u3_u5_n156 ) , .A1( u2_u3_u5_n174 ) );
  NOR2_X1 u2_u3_u5_U47 (.ZN( u2_u3_u5_n121 ) , .A2( u2_u3_u5_n145 ) , .A1( u2_u3_u5_n176 ) );
  AOI22_X1 u2_u3_u5_U48 (.ZN( u2_u3_u5_n114 ) , .A2( u2_u3_u5_n137 ) , .A1( u2_u3_u5_n145 ) , .B2( u2_u3_u5_n175 ) , .B1( u2_u3_u5_n193 ) );
  OAI211_X1 u2_u3_u5_U49 (.B( u2_u3_u5_n124 ) , .A( u2_u3_u5_n125 ) , .C2( u2_u3_u5_n126 ) , .C1( u2_u3_u5_n127 ) , .ZN( u2_u3_u5_n128 ) );
  OAI21_X1 u2_u3_u5_U5 (.B2( u2_u3_u5_n136 ) , .B1( u2_u3_u5_n137 ) , .ZN( u2_u3_u5_n138 ) , .A( u2_u3_u5_n177 ) );
  NOR3_X1 u2_u3_u5_U50 (.ZN( u2_u3_u5_n127 ) , .A1( u2_u3_u5_n136 ) , .A3( u2_u3_u5_n148 ) , .A2( u2_u3_u5_n182 ) );
  OAI21_X1 u2_u3_u5_U51 (.ZN( u2_u3_u5_n124 ) , .A( u2_u3_u5_n177 ) , .B2( u2_u3_u5_n183 ) , .B1( u2_u3_u5_n189 ) );
  OAI21_X1 u2_u3_u5_U52 (.ZN( u2_u3_u5_n125 ) , .A( u2_u3_u5_n174 ) , .B2( u2_u3_u5_n185 ) , .B1( u2_u3_u5_n190 ) );
  AOI21_X1 u2_u3_u5_U53 (.A( u2_u3_u5_n153 ) , .B2( u2_u3_u5_n154 ) , .B1( u2_u3_u5_n155 ) , .ZN( u2_u3_u5_n164 ) );
  AOI21_X1 u2_u3_u5_U54 (.ZN( u2_u3_u5_n110 ) , .B1( u2_u3_u5_n122 ) , .B2( u2_u3_u5_n139 ) , .A( u2_u3_u5_n153 ) );
  INV_X1 u2_u3_u5_U55 (.A( u2_u3_u5_n153 ) , .ZN( u2_u3_u5_n176 ) );
  INV_X1 u2_u3_u5_U56 (.A( u2_u3_u5_n126 ) , .ZN( u2_u3_u5_n173 ) );
  AND2_X1 u2_u3_u5_U57 (.A2( u2_u3_u5_n104 ) , .A1( u2_u3_u5_n107 ) , .ZN( u2_u3_u5_n147 ) );
  AND2_X1 u2_u3_u5_U58 (.A2( u2_u3_u5_n104 ) , .A1( u2_u3_u5_n108 ) , .ZN( u2_u3_u5_n148 ) );
  NAND2_X1 u2_u3_u5_U59 (.A1( u2_u3_u5_n105 ) , .A2( u2_u3_u5_n106 ) , .ZN( u2_u3_u5_n158 ) );
  INV_X1 u2_u3_u5_U6 (.A( u2_u3_u5_n135 ) , .ZN( u2_u3_u5_n178 ) );
  NAND2_X1 u2_u3_u5_U60 (.A2( u2_u3_u5_n108 ) , .A1( u2_u3_u5_n109 ) , .ZN( u2_u3_u5_n139 ) );
  NAND2_X1 u2_u3_u5_U61 (.A1( u2_u3_u5_n106 ) , .A2( u2_u3_u5_n108 ) , .ZN( u2_u3_u5_n119 ) );
  NAND2_X1 u2_u3_u5_U62 (.A2( u2_u3_u5_n103 ) , .A1( u2_u3_u5_n105 ) , .ZN( u2_u3_u5_n140 ) );
  NAND2_X1 u2_u3_u5_U63 (.A2( u2_u3_u5_n104 ) , .A1( u2_u3_u5_n105 ) , .ZN( u2_u3_u5_n155 ) );
  NAND2_X1 u2_u3_u5_U64 (.A2( u2_u3_u5_n106 ) , .A1( u2_u3_u5_n107 ) , .ZN( u2_u3_u5_n122 ) );
  NAND2_X1 u2_u3_u5_U65 (.A2( u2_u3_u5_n100 ) , .A1( u2_u3_u5_n106 ) , .ZN( u2_u3_u5_n115 ) );
  NAND2_X1 u2_u3_u5_U66 (.A2( u2_u3_u5_n100 ) , .A1( u2_u3_u5_n103 ) , .ZN( u2_u3_u5_n161 ) );
  NAND2_X1 u2_u3_u5_U67 (.A1( u2_u3_u5_n105 ) , .A2( u2_u3_u5_n109 ) , .ZN( u2_u3_u5_n154 ) );
  INV_X1 u2_u3_u5_U68 (.A( u2_u3_u5_n146 ) , .ZN( u2_u3_u5_n172 ) );
  NAND2_X1 u2_u3_u5_U69 (.A1( u2_u3_u5_n103 ) , .A2( u2_u3_u5_n108 ) , .ZN( u2_u3_u5_n123 ) );
  OAI22_X1 u2_u3_u5_U7 (.B2( u2_u3_u5_n149 ) , .B1( u2_u3_u5_n150 ) , .A2( u2_u3_u5_n151 ) , .A1( u2_u3_u5_n152 ) , .ZN( u2_u3_u5_n165 ) );
  NAND2_X1 u2_u3_u5_U70 (.A2( u2_u3_u5_n103 ) , .A1( u2_u3_u5_n107 ) , .ZN( u2_u3_u5_n151 ) );
  NAND2_X1 u2_u3_u5_U71 (.A2( u2_u3_u5_n107 ) , .A1( u2_u3_u5_n109 ) , .ZN( u2_u3_u5_n120 ) );
  NAND2_X1 u2_u3_u5_U72 (.A2( u2_u3_u5_n100 ) , .A1( u2_u3_u5_n109 ) , .ZN( u2_u3_u5_n157 ) );
  AND2_X1 u2_u3_u5_U73 (.A2( u2_u3_u5_n100 ) , .A1( u2_u3_u5_n104 ) , .ZN( u2_u3_u5_n131 ) );
  INV_X1 u2_u3_u5_U74 (.A( u2_u3_u5_n102 ) , .ZN( u2_u3_u5_n195 ) );
  OAI221_X1 u2_u3_u5_U75 (.A( u2_u3_u5_n101 ) , .ZN( u2_u3_u5_n102 ) , .C2( u2_u3_u5_n115 ) , .C1( u2_u3_u5_n126 ) , .B1( u2_u3_u5_n134 ) , .B2( u2_u3_u5_n160 ) );
  OAI21_X1 u2_u3_u5_U76 (.ZN( u2_u3_u5_n101 ) , .B1( u2_u3_u5_n137 ) , .A( u2_u3_u5_n146 ) , .B2( u2_u3_u5_n147 ) );
  NOR2_X1 u2_u3_u5_U77 (.A2( u2_u3_X_34 ) , .A1( u2_u3_X_35 ) , .ZN( u2_u3_u5_n145 ) );
  NOR2_X1 u2_u3_u5_U78 (.A2( u2_u3_X_34 ) , .ZN( u2_u3_u5_n146 ) , .A1( u2_u3_u5_n171 ) );
  NOR2_X1 u2_u3_u5_U79 (.A2( u2_u3_X_31 ) , .A1( u2_u3_X_32 ) , .ZN( u2_u3_u5_n103 ) );
  NOR3_X1 u2_u3_u5_U8 (.A2( u2_u3_u5_n147 ) , .A1( u2_u3_u5_n148 ) , .ZN( u2_u3_u5_n149 ) , .A3( u2_u3_u5_n194 ) );
  NOR2_X1 u2_u3_u5_U80 (.A2( u2_u3_X_36 ) , .ZN( u2_u3_u5_n105 ) , .A1( u2_u3_u5_n180 ) );
  NOR2_X1 u2_u3_u5_U81 (.A2( u2_u3_X_33 ) , .ZN( u2_u3_u5_n108 ) , .A1( u2_u3_u5_n170 ) );
  NOR2_X1 u2_u3_u5_U82 (.A2( u2_u3_X_33 ) , .A1( u2_u3_X_36 ) , .ZN( u2_u3_u5_n107 ) );
  NOR2_X1 u2_u3_u5_U83 (.A2( u2_u3_X_31 ) , .ZN( u2_u3_u5_n104 ) , .A1( u2_u3_u5_n181 ) );
  NAND2_X1 u2_u3_u5_U84 (.A2( u2_u3_X_34 ) , .A1( u2_u3_X_35 ) , .ZN( u2_u3_u5_n153 ) );
  NAND2_X1 u2_u3_u5_U85 (.A1( u2_u3_X_34 ) , .ZN( u2_u3_u5_n126 ) , .A2( u2_u3_u5_n171 ) );
  AND2_X1 u2_u3_u5_U86 (.A1( u2_u3_X_31 ) , .A2( u2_u3_X_32 ) , .ZN( u2_u3_u5_n106 ) );
  AND2_X1 u2_u3_u5_U87 (.A1( u2_u3_X_31 ) , .ZN( u2_u3_u5_n109 ) , .A2( u2_u3_u5_n181 ) );
  INV_X1 u2_u3_u5_U88 (.A( u2_u3_X_33 ) , .ZN( u2_u3_u5_n180 ) );
  INV_X1 u2_u3_u5_U89 (.A( u2_u3_X_35 ) , .ZN( u2_u3_u5_n171 ) );
  NOR2_X1 u2_u3_u5_U9 (.ZN( u2_u3_u5_n135 ) , .A1( u2_u3_u5_n173 ) , .A2( u2_u3_u5_n176 ) );
  INV_X1 u2_u3_u5_U90 (.A( u2_u3_X_36 ) , .ZN( u2_u3_u5_n170 ) );
  INV_X1 u2_u3_u5_U91 (.A( u2_u3_X_32 ) , .ZN( u2_u3_u5_n181 ) );
  NAND4_X1 u2_u3_u5_U92 (.ZN( u2_out3_29 ) , .A4( u2_u3_u5_n129 ) , .A3( u2_u3_u5_n130 ) , .A2( u2_u3_u5_n168 ) , .A1( u2_u3_u5_n196 ) );
  AOI221_X1 u2_u3_u5_U93 (.A( u2_u3_u5_n128 ) , .ZN( u2_u3_u5_n129 ) , .C2( u2_u3_u5_n132 ) , .B2( u2_u3_u5_n159 ) , .B1( u2_u3_u5_n176 ) , .C1( u2_u3_u5_n184 ) );
  AOI222_X1 u2_u3_u5_U94 (.ZN( u2_u3_u5_n130 ) , .A2( u2_u3_u5_n146 ) , .B1( u2_u3_u5_n147 ) , .C2( u2_u3_u5_n175 ) , .B2( u2_u3_u5_n179 ) , .A1( u2_u3_u5_n188 ) , .C1( u2_u3_u5_n194 ) );
  NAND4_X1 u2_u3_u5_U95 (.ZN( u2_out3_19 ) , .A4( u2_u3_u5_n166 ) , .A3( u2_u3_u5_n167 ) , .A2( u2_u3_u5_n168 ) , .A1( u2_u3_u5_n169 ) );
  AOI22_X1 u2_u3_u5_U96 (.B2( u2_u3_u5_n145 ) , .A2( u2_u3_u5_n146 ) , .ZN( u2_u3_u5_n167 ) , .B1( u2_u3_u5_n182 ) , .A1( u2_u3_u5_n189 ) );
  NOR4_X1 u2_u3_u5_U97 (.A4( u2_u3_u5_n162 ) , .A3( u2_u3_u5_n163 ) , .A2( u2_u3_u5_n164 ) , .A1( u2_u3_u5_n165 ) , .ZN( u2_u3_u5_n166 ) );
  NAND4_X1 u2_u3_u5_U98 (.ZN( u2_out3_11 ) , .A4( u2_u3_u5_n143 ) , .A3( u2_u3_u5_n144 ) , .A2( u2_u3_u5_n169 ) , .A1( u2_u3_u5_n196 ) );
  AOI22_X1 u2_u3_u5_U99 (.A2( u2_u3_u5_n132 ) , .ZN( u2_u3_u5_n144 ) , .B2( u2_u3_u5_n145 ) , .B1( u2_u3_u5_n184 ) , .A1( u2_u3_u5_n194 ) );
  XOR2_X1 u2_u4_U1 (.B( u2_K5_9 ) , .A( u2_R3_6 ) , .Z( u2_u4_X_9 ) );
  XOR2_X1 u2_u4_U2 (.B( u2_K5_8 ) , .A( u2_R3_5 ) , .Z( u2_u4_X_8 ) );
  XOR2_X1 u2_u4_U3 (.B( u2_K5_7 ) , .A( u2_R3_4 ) , .Z( u2_u4_X_7 ) );
  XOR2_X1 u2_u4_U33 (.B( u2_K5_24 ) , .A( u2_R3_17 ) , .Z( u2_u4_X_24 ) );
  XOR2_X1 u2_u4_U34 (.B( u2_K5_23 ) , .A( u2_R3_16 ) , .Z( u2_u4_X_23 ) );
  XOR2_X1 u2_u4_U35 (.B( u2_K5_22 ) , .A( u2_R3_15 ) , .Z( u2_u4_X_22 ) );
  XOR2_X1 u2_u4_U36 (.B( u2_K5_21 ) , .A( u2_R3_14 ) , .Z( u2_u4_X_21 ) );
  XOR2_X1 u2_u4_U37 (.B( u2_K5_20 ) , .A( u2_R3_13 ) , .Z( u2_u4_X_20 ) );
  XOR2_X1 u2_u4_U39 (.B( u2_K5_19 ) , .A( u2_R3_12 ) , .Z( u2_u4_X_19 ) );
  XOR2_X1 u2_u4_U40 (.B( u2_K5_18 ) , .A( u2_R3_13 ) , .Z( u2_u4_X_18 ) );
  XOR2_X1 u2_u4_U41 (.B( u2_K5_17 ) , .A( u2_R3_12 ) , .Z( u2_u4_X_17 ) );
  XOR2_X1 u2_u4_U42 (.B( u2_K5_16 ) , .A( u2_R3_11 ) , .Z( u2_u4_X_16 ) );
  XOR2_X1 u2_u4_U43 (.B( u2_K5_15 ) , .A( u2_R3_10 ) , .Z( u2_u4_X_15 ) );
  XOR2_X1 u2_u4_U44 (.B( u2_K5_14 ) , .A( u2_R3_9 ) , .Z( u2_u4_X_14 ) );
  XOR2_X1 u2_u4_U45 (.B( u2_K5_13 ) , .A( u2_R3_8 ) , .Z( u2_u4_X_13 ) );
  XOR2_X1 u2_u4_U46 (.B( u2_K5_12 ) , .A( u2_R3_9 ) , .Z( u2_u4_X_12 ) );
  XOR2_X1 u2_u4_U47 (.B( u2_K5_11 ) , .A( u2_R3_8 ) , .Z( u2_u4_X_11 ) );
  XOR2_X1 u2_u4_U48 (.B( u2_K5_10 ) , .A( u2_R3_7 ) , .Z( u2_u4_X_10 ) );
  NOR2_X1 u2_u4_u1_U10 (.A1( u2_u4_u1_n112 ) , .A2( u2_u4_u1_n116 ) , .ZN( u2_u4_u1_n118 ) );
  NAND3_X1 u2_u4_u1_U100 (.ZN( u2_u4_u1_n113 ) , .A1( u2_u4_u1_n120 ) , .A3( u2_u4_u1_n133 ) , .A2( u2_u4_u1_n155 ) );
  OAI21_X1 u2_u4_u1_U11 (.ZN( u2_u4_u1_n101 ) , .B1( u2_u4_u1_n141 ) , .A( u2_u4_u1_n146 ) , .B2( u2_u4_u1_n183 ) );
  AOI21_X1 u2_u4_u1_U12 (.B2( u2_u4_u1_n155 ) , .B1( u2_u4_u1_n156 ) , .ZN( u2_u4_u1_n157 ) , .A( u2_u4_u1_n174 ) );
  NAND2_X1 u2_u4_u1_U13 (.ZN( u2_u4_u1_n140 ) , .A2( u2_u4_u1_n150 ) , .A1( u2_u4_u1_n155 ) );
  NAND2_X1 u2_u4_u1_U14 (.A1( u2_u4_u1_n131 ) , .ZN( u2_u4_u1_n147 ) , .A2( u2_u4_u1_n153 ) );
  INV_X1 u2_u4_u1_U15 (.A( u2_u4_u1_n139 ) , .ZN( u2_u4_u1_n174 ) );
  OR4_X1 u2_u4_u1_U16 (.A4( u2_u4_u1_n106 ) , .A3( u2_u4_u1_n107 ) , .ZN( u2_u4_u1_n108 ) , .A1( u2_u4_u1_n117 ) , .A2( u2_u4_u1_n184 ) );
  AOI21_X1 u2_u4_u1_U17 (.ZN( u2_u4_u1_n106 ) , .A( u2_u4_u1_n112 ) , .B1( u2_u4_u1_n154 ) , .B2( u2_u4_u1_n156 ) );
  AOI21_X1 u2_u4_u1_U18 (.ZN( u2_u4_u1_n107 ) , .B1( u2_u4_u1_n134 ) , .B2( u2_u4_u1_n149 ) , .A( u2_u4_u1_n174 ) );
  INV_X1 u2_u4_u1_U19 (.A( u2_u4_u1_n101 ) , .ZN( u2_u4_u1_n184 ) );
  INV_X1 u2_u4_u1_U20 (.A( u2_u4_u1_n112 ) , .ZN( u2_u4_u1_n171 ) );
  NAND2_X1 u2_u4_u1_U21 (.ZN( u2_u4_u1_n141 ) , .A1( u2_u4_u1_n153 ) , .A2( u2_u4_u1_n156 ) );
  AND2_X1 u2_u4_u1_U22 (.A1( u2_u4_u1_n123 ) , .ZN( u2_u4_u1_n134 ) , .A2( u2_u4_u1_n161 ) );
  NAND2_X1 u2_u4_u1_U23 (.A2( u2_u4_u1_n115 ) , .A1( u2_u4_u1_n116 ) , .ZN( u2_u4_u1_n148 ) );
  NAND2_X1 u2_u4_u1_U24 (.A2( u2_u4_u1_n133 ) , .A1( u2_u4_u1_n135 ) , .ZN( u2_u4_u1_n159 ) );
  NAND2_X1 u2_u4_u1_U25 (.A2( u2_u4_u1_n115 ) , .A1( u2_u4_u1_n120 ) , .ZN( u2_u4_u1_n132 ) );
  INV_X1 u2_u4_u1_U26 (.A( u2_u4_u1_n154 ) , .ZN( u2_u4_u1_n178 ) );
  INV_X1 u2_u4_u1_U27 (.A( u2_u4_u1_n151 ) , .ZN( u2_u4_u1_n183 ) );
  AND2_X1 u2_u4_u1_U28 (.A1( u2_u4_u1_n129 ) , .A2( u2_u4_u1_n133 ) , .ZN( u2_u4_u1_n149 ) );
  INV_X1 u2_u4_u1_U29 (.A( u2_u4_u1_n131 ) , .ZN( u2_u4_u1_n180 ) );
  INV_X1 u2_u4_u1_U3 (.A( u2_u4_u1_n159 ) , .ZN( u2_u4_u1_n182 ) );
  OAI221_X1 u2_u4_u1_U30 (.A( u2_u4_u1_n119 ) , .C2( u2_u4_u1_n129 ) , .ZN( u2_u4_u1_n138 ) , .B2( u2_u4_u1_n152 ) , .C1( u2_u4_u1_n174 ) , .B1( u2_u4_u1_n187 ) );
  INV_X1 u2_u4_u1_U31 (.A( u2_u4_u1_n148 ) , .ZN( u2_u4_u1_n187 ) );
  AOI211_X1 u2_u4_u1_U32 (.B( u2_u4_u1_n117 ) , .A( u2_u4_u1_n118 ) , .ZN( u2_u4_u1_n119 ) , .C2( u2_u4_u1_n146 ) , .C1( u2_u4_u1_n159 ) );
  NOR2_X1 u2_u4_u1_U33 (.A1( u2_u4_u1_n168 ) , .A2( u2_u4_u1_n176 ) , .ZN( u2_u4_u1_n98 ) );
  AOI211_X1 u2_u4_u1_U34 (.B( u2_u4_u1_n162 ) , .A( u2_u4_u1_n163 ) , .C2( u2_u4_u1_n164 ) , .ZN( u2_u4_u1_n165 ) , .C1( u2_u4_u1_n171 ) );
  AOI21_X1 u2_u4_u1_U35 (.A( u2_u4_u1_n160 ) , .B2( u2_u4_u1_n161 ) , .ZN( u2_u4_u1_n162 ) , .B1( u2_u4_u1_n182 ) );
  OR2_X1 u2_u4_u1_U36 (.A2( u2_u4_u1_n157 ) , .A1( u2_u4_u1_n158 ) , .ZN( u2_u4_u1_n163 ) );
  NAND2_X1 u2_u4_u1_U37 (.A1( u2_u4_u1_n128 ) , .ZN( u2_u4_u1_n146 ) , .A2( u2_u4_u1_n160 ) );
  NAND2_X1 u2_u4_u1_U38 (.A2( u2_u4_u1_n112 ) , .ZN( u2_u4_u1_n139 ) , .A1( u2_u4_u1_n152 ) );
  NAND2_X1 u2_u4_u1_U39 (.A1( u2_u4_u1_n105 ) , .ZN( u2_u4_u1_n156 ) , .A2( u2_u4_u1_n99 ) );
  AOI221_X1 u2_u4_u1_U4 (.A( u2_u4_u1_n138 ) , .C2( u2_u4_u1_n139 ) , .C1( u2_u4_u1_n140 ) , .B2( u2_u4_u1_n141 ) , .ZN( u2_u4_u1_n142 ) , .B1( u2_u4_u1_n175 ) );
  AOI221_X1 u2_u4_u1_U40 (.B1( u2_u4_u1_n140 ) , .ZN( u2_u4_u1_n167 ) , .B2( u2_u4_u1_n172 ) , .C2( u2_u4_u1_n175 ) , .C1( u2_u4_u1_n178 ) , .A( u2_u4_u1_n188 ) );
  INV_X1 u2_u4_u1_U41 (.ZN( u2_u4_u1_n188 ) , .A( u2_u4_u1_n97 ) );
  AOI211_X1 u2_u4_u1_U42 (.A( u2_u4_u1_n118 ) , .C1( u2_u4_u1_n132 ) , .C2( u2_u4_u1_n139 ) , .B( u2_u4_u1_n96 ) , .ZN( u2_u4_u1_n97 ) );
  AOI21_X1 u2_u4_u1_U43 (.B2( u2_u4_u1_n121 ) , .B1( u2_u4_u1_n135 ) , .A( u2_u4_u1_n152 ) , .ZN( u2_u4_u1_n96 ) );
  NOR2_X1 u2_u4_u1_U44 (.ZN( u2_u4_u1_n117 ) , .A1( u2_u4_u1_n121 ) , .A2( u2_u4_u1_n160 ) );
  OAI21_X1 u2_u4_u1_U45 (.B2( u2_u4_u1_n123 ) , .ZN( u2_u4_u1_n145 ) , .B1( u2_u4_u1_n160 ) , .A( u2_u4_u1_n185 ) );
  INV_X1 u2_u4_u1_U46 (.A( u2_u4_u1_n122 ) , .ZN( u2_u4_u1_n185 ) );
  AOI21_X1 u2_u4_u1_U47 (.B2( u2_u4_u1_n120 ) , .B1( u2_u4_u1_n121 ) , .ZN( u2_u4_u1_n122 ) , .A( u2_u4_u1_n128 ) );
  AOI21_X1 u2_u4_u1_U48 (.A( u2_u4_u1_n128 ) , .B2( u2_u4_u1_n129 ) , .ZN( u2_u4_u1_n130 ) , .B1( u2_u4_u1_n150 ) );
  NAND2_X1 u2_u4_u1_U49 (.ZN( u2_u4_u1_n112 ) , .A1( u2_u4_u1_n169 ) , .A2( u2_u4_u1_n170 ) );
  AOI211_X1 u2_u4_u1_U5 (.ZN( u2_u4_u1_n124 ) , .A( u2_u4_u1_n138 ) , .C2( u2_u4_u1_n139 ) , .B( u2_u4_u1_n145 ) , .C1( u2_u4_u1_n147 ) );
  NAND2_X1 u2_u4_u1_U50 (.ZN( u2_u4_u1_n129 ) , .A2( u2_u4_u1_n95 ) , .A1( u2_u4_u1_n98 ) );
  NAND2_X1 u2_u4_u1_U51 (.A1( u2_u4_u1_n102 ) , .ZN( u2_u4_u1_n154 ) , .A2( u2_u4_u1_n99 ) );
  NAND2_X1 u2_u4_u1_U52 (.A2( u2_u4_u1_n100 ) , .ZN( u2_u4_u1_n135 ) , .A1( u2_u4_u1_n99 ) );
  AOI21_X1 u2_u4_u1_U53 (.A( u2_u4_u1_n152 ) , .B2( u2_u4_u1_n153 ) , .B1( u2_u4_u1_n154 ) , .ZN( u2_u4_u1_n158 ) );
  INV_X1 u2_u4_u1_U54 (.A( u2_u4_u1_n160 ) , .ZN( u2_u4_u1_n175 ) );
  NAND2_X1 u2_u4_u1_U55 (.A1( u2_u4_u1_n100 ) , .ZN( u2_u4_u1_n116 ) , .A2( u2_u4_u1_n95 ) );
  NAND2_X1 u2_u4_u1_U56 (.A1( u2_u4_u1_n102 ) , .ZN( u2_u4_u1_n131 ) , .A2( u2_u4_u1_n95 ) );
  NAND2_X1 u2_u4_u1_U57 (.A2( u2_u4_u1_n104 ) , .ZN( u2_u4_u1_n121 ) , .A1( u2_u4_u1_n98 ) );
  NAND2_X1 u2_u4_u1_U58 (.A1( u2_u4_u1_n103 ) , .ZN( u2_u4_u1_n153 ) , .A2( u2_u4_u1_n98 ) );
  NAND2_X1 u2_u4_u1_U59 (.A2( u2_u4_u1_n104 ) , .A1( u2_u4_u1_n105 ) , .ZN( u2_u4_u1_n133 ) );
  AOI22_X1 u2_u4_u1_U6 (.B2( u2_u4_u1_n113 ) , .A2( u2_u4_u1_n114 ) , .ZN( u2_u4_u1_n125 ) , .A1( u2_u4_u1_n171 ) , .B1( u2_u4_u1_n173 ) );
  NAND2_X1 u2_u4_u1_U60 (.ZN( u2_u4_u1_n150 ) , .A2( u2_u4_u1_n98 ) , .A1( u2_u4_u1_n99 ) );
  NAND2_X1 u2_u4_u1_U61 (.A1( u2_u4_u1_n105 ) , .ZN( u2_u4_u1_n155 ) , .A2( u2_u4_u1_n95 ) );
  OAI21_X1 u2_u4_u1_U62 (.ZN( u2_u4_u1_n109 ) , .B1( u2_u4_u1_n129 ) , .B2( u2_u4_u1_n160 ) , .A( u2_u4_u1_n167 ) );
  NAND2_X1 u2_u4_u1_U63 (.A2( u2_u4_u1_n100 ) , .A1( u2_u4_u1_n103 ) , .ZN( u2_u4_u1_n120 ) );
  NAND2_X1 u2_u4_u1_U64 (.A1( u2_u4_u1_n102 ) , .A2( u2_u4_u1_n104 ) , .ZN( u2_u4_u1_n115 ) );
  NAND2_X1 u2_u4_u1_U65 (.A2( u2_u4_u1_n100 ) , .A1( u2_u4_u1_n104 ) , .ZN( u2_u4_u1_n151 ) );
  NAND2_X1 u2_u4_u1_U66 (.A2( u2_u4_u1_n103 ) , .A1( u2_u4_u1_n105 ) , .ZN( u2_u4_u1_n161 ) );
  INV_X1 u2_u4_u1_U67 (.A( u2_u4_u1_n152 ) , .ZN( u2_u4_u1_n173 ) );
  INV_X1 u2_u4_u1_U68 (.A( u2_u4_u1_n128 ) , .ZN( u2_u4_u1_n172 ) );
  NAND2_X1 u2_u4_u1_U69 (.A2( u2_u4_u1_n102 ) , .A1( u2_u4_u1_n103 ) , .ZN( u2_u4_u1_n123 ) );
  NAND2_X1 u2_u4_u1_U7 (.ZN( u2_u4_u1_n114 ) , .A1( u2_u4_u1_n134 ) , .A2( u2_u4_u1_n156 ) );
  NOR2_X1 u2_u4_u1_U70 (.A2( u2_u4_X_7 ) , .A1( u2_u4_X_8 ) , .ZN( u2_u4_u1_n95 ) );
  NOR2_X1 u2_u4_u1_U71 (.A1( u2_u4_X_12 ) , .A2( u2_u4_X_9 ) , .ZN( u2_u4_u1_n100 ) );
  NOR2_X1 u2_u4_u1_U72 (.A2( u2_u4_X_8 ) , .A1( u2_u4_u1_n177 ) , .ZN( u2_u4_u1_n99 ) );
  NOR2_X1 u2_u4_u1_U73 (.A2( u2_u4_X_12 ) , .ZN( u2_u4_u1_n102 ) , .A1( u2_u4_u1_n176 ) );
  NOR2_X1 u2_u4_u1_U74 (.A2( u2_u4_X_9 ) , .ZN( u2_u4_u1_n105 ) , .A1( u2_u4_u1_n168 ) );
  NAND2_X1 u2_u4_u1_U75 (.A1( u2_u4_X_10 ) , .ZN( u2_u4_u1_n160 ) , .A2( u2_u4_u1_n169 ) );
  NAND2_X1 u2_u4_u1_U76 (.A2( u2_u4_X_10 ) , .A1( u2_u4_X_11 ) , .ZN( u2_u4_u1_n152 ) );
  NAND2_X1 u2_u4_u1_U77 (.A1( u2_u4_X_11 ) , .ZN( u2_u4_u1_n128 ) , .A2( u2_u4_u1_n170 ) );
  AND2_X1 u2_u4_u1_U78 (.A2( u2_u4_X_7 ) , .A1( u2_u4_X_8 ) , .ZN( u2_u4_u1_n104 ) );
  AND2_X1 u2_u4_u1_U79 (.A1( u2_u4_X_8 ) , .ZN( u2_u4_u1_n103 ) , .A2( u2_u4_u1_n177 ) );
  AOI22_X1 u2_u4_u1_U8 (.B2( u2_u4_u1_n136 ) , .A2( u2_u4_u1_n137 ) , .ZN( u2_u4_u1_n143 ) , .A1( u2_u4_u1_n171 ) , .B1( u2_u4_u1_n173 ) );
  INV_X1 u2_u4_u1_U80 (.A( u2_u4_X_10 ) , .ZN( u2_u4_u1_n170 ) );
  INV_X1 u2_u4_u1_U81 (.A( u2_u4_X_9 ) , .ZN( u2_u4_u1_n176 ) );
  INV_X1 u2_u4_u1_U82 (.A( u2_u4_X_11 ) , .ZN( u2_u4_u1_n169 ) );
  INV_X1 u2_u4_u1_U83 (.A( u2_u4_X_12 ) , .ZN( u2_u4_u1_n168 ) );
  INV_X1 u2_u4_u1_U84 (.A( u2_u4_X_7 ) , .ZN( u2_u4_u1_n177 ) );
  NAND4_X1 u2_u4_u1_U85 (.ZN( u2_out4_28 ) , .A4( u2_u4_u1_n124 ) , .A3( u2_u4_u1_n125 ) , .A2( u2_u4_u1_n126 ) , .A1( u2_u4_u1_n127 ) );
  OAI21_X1 u2_u4_u1_U86 (.ZN( u2_u4_u1_n127 ) , .B2( u2_u4_u1_n139 ) , .B1( u2_u4_u1_n175 ) , .A( u2_u4_u1_n183 ) );
  OAI21_X1 u2_u4_u1_U87 (.ZN( u2_u4_u1_n126 ) , .B2( u2_u4_u1_n140 ) , .A( u2_u4_u1_n146 ) , .B1( u2_u4_u1_n178 ) );
  NAND4_X1 u2_u4_u1_U88 (.ZN( u2_out4_18 ) , .A4( u2_u4_u1_n165 ) , .A3( u2_u4_u1_n166 ) , .A1( u2_u4_u1_n167 ) , .A2( u2_u4_u1_n186 ) );
  AOI22_X1 u2_u4_u1_U89 (.B2( u2_u4_u1_n146 ) , .B1( u2_u4_u1_n147 ) , .A2( u2_u4_u1_n148 ) , .ZN( u2_u4_u1_n166 ) , .A1( u2_u4_u1_n172 ) );
  INV_X1 u2_u4_u1_U9 (.A( u2_u4_u1_n147 ) , .ZN( u2_u4_u1_n181 ) );
  INV_X1 u2_u4_u1_U90 (.A( u2_u4_u1_n145 ) , .ZN( u2_u4_u1_n186 ) );
  NAND4_X1 u2_u4_u1_U91 (.ZN( u2_out4_2 ) , .A4( u2_u4_u1_n142 ) , .A3( u2_u4_u1_n143 ) , .A2( u2_u4_u1_n144 ) , .A1( u2_u4_u1_n179 ) );
  OAI21_X1 u2_u4_u1_U92 (.B2( u2_u4_u1_n132 ) , .ZN( u2_u4_u1_n144 ) , .A( u2_u4_u1_n146 ) , .B1( u2_u4_u1_n180 ) );
  INV_X1 u2_u4_u1_U93 (.A( u2_u4_u1_n130 ) , .ZN( u2_u4_u1_n179 ) );
  OR4_X1 u2_u4_u1_U94 (.ZN( u2_out4_13 ) , .A4( u2_u4_u1_n108 ) , .A3( u2_u4_u1_n109 ) , .A2( u2_u4_u1_n110 ) , .A1( u2_u4_u1_n111 ) );
  AOI21_X1 u2_u4_u1_U95 (.ZN( u2_u4_u1_n111 ) , .A( u2_u4_u1_n128 ) , .B2( u2_u4_u1_n131 ) , .B1( u2_u4_u1_n135 ) );
  AOI21_X1 u2_u4_u1_U96 (.ZN( u2_u4_u1_n110 ) , .A( u2_u4_u1_n116 ) , .B1( u2_u4_u1_n152 ) , .B2( u2_u4_u1_n160 ) );
  NAND3_X1 u2_u4_u1_U97 (.A3( u2_u4_u1_n149 ) , .A2( u2_u4_u1_n150 ) , .A1( u2_u4_u1_n151 ) , .ZN( u2_u4_u1_n164 ) );
  NAND3_X1 u2_u4_u1_U98 (.A3( u2_u4_u1_n134 ) , .A2( u2_u4_u1_n135 ) , .ZN( u2_u4_u1_n136 ) , .A1( u2_u4_u1_n151 ) );
  NAND3_X1 u2_u4_u1_U99 (.A1( u2_u4_u1_n133 ) , .ZN( u2_u4_u1_n137 ) , .A2( u2_u4_u1_n154 ) , .A3( u2_u4_u1_n181 ) );
  OAI22_X1 u2_u4_u2_U10 (.ZN( u2_u4_u2_n109 ) , .A2( u2_u4_u2_n113 ) , .B2( u2_u4_u2_n133 ) , .B1( u2_u4_u2_n167 ) , .A1( u2_u4_u2_n168 ) );
  NAND3_X1 u2_u4_u2_U100 (.A2( u2_u4_u2_n100 ) , .A1( u2_u4_u2_n104 ) , .A3( u2_u4_u2_n138 ) , .ZN( u2_u4_u2_n98 ) );
  OAI22_X1 u2_u4_u2_U11 (.B1( u2_u4_u2_n151 ) , .A2( u2_u4_u2_n152 ) , .A1( u2_u4_u2_n153 ) , .ZN( u2_u4_u2_n160 ) , .B2( u2_u4_u2_n168 ) );
  NOR3_X1 u2_u4_u2_U12 (.A1( u2_u4_u2_n150 ) , .ZN( u2_u4_u2_n151 ) , .A3( u2_u4_u2_n175 ) , .A2( u2_u4_u2_n188 ) );
  AOI21_X1 u2_u4_u2_U13 (.ZN( u2_u4_u2_n144 ) , .B2( u2_u4_u2_n155 ) , .A( u2_u4_u2_n172 ) , .B1( u2_u4_u2_n185 ) );
  AOI21_X1 u2_u4_u2_U14 (.B2( u2_u4_u2_n143 ) , .ZN( u2_u4_u2_n145 ) , .B1( u2_u4_u2_n152 ) , .A( u2_u4_u2_n171 ) );
  AOI21_X1 u2_u4_u2_U15 (.B2( u2_u4_u2_n120 ) , .B1( u2_u4_u2_n121 ) , .ZN( u2_u4_u2_n126 ) , .A( u2_u4_u2_n167 ) );
  INV_X1 u2_u4_u2_U16 (.A( u2_u4_u2_n156 ) , .ZN( u2_u4_u2_n171 ) );
  INV_X1 u2_u4_u2_U17 (.A( u2_u4_u2_n120 ) , .ZN( u2_u4_u2_n188 ) );
  NAND2_X1 u2_u4_u2_U18 (.A2( u2_u4_u2_n122 ) , .ZN( u2_u4_u2_n150 ) , .A1( u2_u4_u2_n152 ) );
  INV_X1 u2_u4_u2_U19 (.A( u2_u4_u2_n153 ) , .ZN( u2_u4_u2_n170 ) );
  INV_X1 u2_u4_u2_U20 (.A( u2_u4_u2_n137 ) , .ZN( u2_u4_u2_n173 ) );
  NAND2_X1 u2_u4_u2_U21 (.A1( u2_u4_u2_n132 ) , .A2( u2_u4_u2_n139 ) , .ZN( u2_u4_u2_n157 ) );
  INV_X1 u2_u4_u2_U22 (.A( u2_u4_u2_n113 ) , .ZN( u2_u4_u2_n178 ) );
  INV_X1 u2_u4_u2_U23 (.A( u2_u4_u2_n139 ) , .ZN( u2_u4_u2_n175 ) );
  INV_X1 u2_u4_u2_U24 (.A( u2_u4_u2_n155 ) , .ZN( u2_u4_u2_n181 ) );
  INV_X1 u2_u4_u2_U25 (.A( u2_u4_u2_n119 ) , .ZN( u2_u4_u2_n177 ) );
  INV_X1 u2_u4_u2_U26 (.A( u2_u4_u2_n116 ) , .ZN( u2_u4_u2_n180 ) );
  INV_X1 u2_u4_u2_U27 (.A( u2_u4_u2_n131 ) , .ZN( u2_u4_u2_n179 ) );
  INV_X1 u2_u4_u2_U28 (.A( u2_u4_u2_n154 ) , .ZN( u2_u4_u2_n176 ) );
  NAND2_X1 u2_u4_u2_U29 (.A2( u2_u4_u2_n116 ) , .A1( u2_u4_u2_n117 ) , .ZN( u2_u4_u2_n118 ) );
  NOR2_X1 u2_u4_u2_U3 (.ZN( u2_u4_u2_n121 ) , .A2( u2_u4_u2_n177 ) , .A1( u2_u4_u2_n180 ) );
  INV_X1 u2_u4_u2_U30 (.A( u2_u4_u2_n132 ) , .ZN( u2_u4_u2_n182 ) );
  INV_X1 u2_u4_u2_U31 (.A( u2_u4_u2_n158 ) , .ZN( u2_u4_u2_n183 ) );
  OAI21_X1 u2_u4_u2_U32 (.A( u2_u4_u2_n156 ) , .B1( u2_u4_u2_n157 ) , .ZN( u2_u4_u2_n158 ) , .B2( u2_u4_u2_n179 ) );
  NOR2_X1 u2_u4_u2_U33 (.ZN( u2_u4_u2_n156 ) , .A1( u2_u4_u2_n166 ) , .A2( u2_u4_u2_n169 ) );
  NOR2_X1 u2_u4_u2_U34 (.A2( u2_u4_u2_n114 ) , .ZN( u2_u4_u2_n137 ) , .A1( u2_u4_u2_n140 ) );
  NOR2_X1 u2_u4_u2_U35 (.A2( u2_u4_u2_n138 ) , .ZN( u2_u4_u2_n153 ) , .A1( u2_u4_u2_n156 ) );
  AOI211_X1 u2_u4_u2_U36 (.ZN( u2_u4_u2_n130 ) , .C1( u2_u4_u2_n138 ) , .C2( u2_u4_u2_n179 ) , .B( u2_u4_u2_n96 ) , .A( u2_u4_u2_n97 ) );
  OAI22_X1 u2_u4_u2_U37 (.B1( u2_u4_u2_n133 ) , .A2( u2_u4_u2_n137 ) , .A1( u2_u4_u2_n152 ) , .B2( u2_u4_u2_n168 ) , .ZN( u2_u4_u2_n97 ) );
  OAI221_X1 u2_u4_u2_U38 (.B1( u2_u4_u2_n113 ) , .C1( u2_u4_u2_n132 ) , .A( u2_u4_u2_n149 ) , .B2( u2_u4_u2_n171 ) , .C2( u2_u4_u2_n172 ) , .ZN( u2_u4_u2_n96 ) );
  OAI221_X1 u2_u4_u2_U39 (.A( u2_u4_u2_n115 ) , .C2( u2_u4_u2_n123 ) , .B2( u2_u4_u2_n143 ) , .B1( u2_u4_u2_n153 ) , .ZN( u2_u4_u2_n163 ) , .C1( u2_u4_u2_n168 ) );
  INV_X1 u2_u4_u2_U4 (.A( u2_u4_u2_n134 ) , .ZN( u2_u4_u2_n185 ) );
  OAI21_X1 u2_u4_u2_U40 (.A( u2_u4_u2_n114 ) , .ZN( u2_u4_u2_n115 ) , .B1( u2_u4_u2_n176 ) , .B2( u2_u4_u2_n178 ) );
  OAI221_X1 u2_u4_u2_U41 (.A( u2_u4_u2_n135 ) , .B2( u2_u4_u2_n136 ) , .B1( u2_u4_u2_n137 ) , .ZN( u2_u4_u2_n162 ) , .C2( u2_u4_u2_n167 ) , .C1( u2_u4_u2_n185 ) );
  AND3_X1 u2_u4_u2_U42 (.A3( u2_u4_u2_n131 ) , .A2( u2_u4_u2_n132 ) , .A1( u2_u4_u2_n133 ) , .ZN( u2_u4_u2_n136 ) );
  AOI22_X1 u2_u4_u2_U43 (.ZN( u2_u4_u2_n135 ) , .B1( u2_u4_u2_n140 ) , .A1( u2_u4_u2_n156 ) , .B2( u2_u4_u2_n180 ) , .A2( u2_u4_u2_n188 ) );
  AOI21_X1 u2_u4_u2_U44 (.ZN( u2_u4_u2_n149 ) , .B1( u2_u4_u2_n173 ) , .B2( u2_u4_u2_n188 ) , .A( u2_u4_u2_n95 ) );
  AND3_X1 u2_u4_u2_U45 (.A2( u2_u4_u2_n100 ) , .A1( u2_u4_u2_n104 ) , .A3( u2_u4_u2_n156 ) , .ZN( u2_u4_u2_n95 ) );
  OAI21_X1 u2_u4_u2_U46 (.A( u2_u4_u2_n101 ) , .B2( u2_u4_u2_n121 ) , .B1( u2_u4_u2_n153 ) , .ZN( u2_u4_u2_n164 ) );
  NAND2_X1 u2_u4_u2_U47 (.A2( u2_u4_u2_n100 ) , .A1( u2_u4_u2_n107 ) , .ZN( u2_u4_u2_n155 ) );
  NAND2_X1 u2_u4_u2_U48 (.A2( u2_u4_u2_n105 ) , .A1( u2_u4_u2_n108 ) , .ZN( u2_u4_u2_n143 ) );
  NAND2_X1 u2_u4_u2_U49 (.A1( u2_u4_u2_n104 ) , .A2( u2_u4_u2_n106 ) , .ZN( u2_u4_u2_n152 ) );
  INV_X1 u2_u4_u2_U5 (.A( u2_u4_u2_n150 ) , .ZN( u2_u4_u2_n184 ) );
  NAND2_X1 u2_u4_u2_U50 (.A1( u2_u4_u2_n100 ) , .A2( u2_u4_u2_n105 ) , .ZN( u2_u4_u2_n132 ) );
  INV_X1 u2_u4_u2_U51 (.A( u2_u4_u2_n140 ) , .ZN( u2_u4_u2_n168 ) );
  INV_X1 u2_u4_u2_U52 (.A( u2_u4_u2_n138 ) , .ZN( u2_u4_u2_n167 ) );
  OAI21_X1 u2_u4_u2_U53 (.A( u2_u4_u2_n141 ) , .B2( u2_u4_u2_n142 ) , .ZN( u2_u4_u2_n146 ) , .B1( u2_u4_u2_n153 ) );
  OAI21_X1 u2_u4_u2_U54 (.A( u2_u4_u2_n140 ) , .ZN( u2_u4_u2_n141 ) , .B1( u2_u4_u2_n176 ) , .B2( u2_u4_u2_n177 ) );
  NOR3_X1 u2_u4_u2_U55 (.ZN( u2_u4_u2_n142 ) , .A3( u2_u4_u2_n175 ) , .A2( u2_u4_u2_n178 ) , .A1( u2_u4_u2_n181 ) );
  INV_X1 u2_u4_u2_U56 (.ZN( u2_u4_u2_n187 ) , .A( u2_u4_u2_n99 ) );
  OAI21_X1 u2_u4_u2_U57 (.B1( u2_u4_u2_n137 ) , .B2( u2_u4_u2_n143 ) , .A( u2_u4_u2_n98 ) , .ZN( u2_u4_u2_n99 ) );
  NAND2_X1 u2_u4_u2_U58 (.A1( u2_u4_u2_n102 ) , .A2( u2_u4_u2_n106 ) , .ZN( u2_u4_u2_n113 ) );
  NAND2_X1 u2_u4_u2_U59 (.A1( u2_u4_u2_n106 ) , .A2( u2_u4_u2_n107 ) , .ZN( u2_u4_u2_n131 ) );
  NOR4_X1 u2_u4_u2_U6 (.A4( u2_u4_u2_n124 ) , .A3( u2_u4_u2_n125 ) , .A2( u2_u4_u2_n126 ) , .A1( u2_u4_u2_n127 ) , .ZN( u2_u4_u2_n128 ) );
  NAND2_X1 u2_u4_u2_U60 (.A1( u2_u4_u2_n103 ) , .A2( u2_u4_u2_n107 ) , .ZN( u2_u4_u2_n139 ) );
  NAND2_X1 u2_u4_u2_U61 (.A1( u2_u4_u2_n103 ) , .A2( u2_u4_u2_n105 ) , .ZN( u2_u4_u2_n133 ) );
  NAND2_X1 u2_u4_u2_U62 (.A1( u2_u4_u2_n102 ) , .A2( u2_u4_u2_n103 ) , .ZN( u2_u4_u2_n154 ) );
  NAND2_X1 u2_u4_u2_U63 (.A2( u2_u4_u2_n103 ) , .A1( u2_u4_u2_n104 ) , .ZN( u2_u4_u2_n119 ) );
  NAND2_X1 u2_u4_u2_U64 (.A2( u2_u4_u2_n107 ) , .A1( u2_u4_u2_n108 ) , .ZN( u2_u4_u2_n123 ) );
  NAND2_X1 u2_u4_u2_U65 (.A1( u2_u4_u2_n104 ) , .A2( u2_u4_u2_n108 ) , .ZN( u2_u4_u2_n122 ) );
  INV_X1 u2_u4_u2_U66 (.A( u2_u4_u2_n114 ) , .ZN( u2_u4_u2_n172 ) );
  NAND2_X1 u2_u4_u2_U67 (.A2( u2_u4_u2_n100 ) , .A1( u2_u4_u2_n102 ) , .ZN( u2_u4_u2_n116 ) );
  NAND2_X1 u2_u4_u2_U68 (.A1( u2_u4_u2_n102 ) , .A2( u2_u4_u2_n108 ) , .ZN( u2_u4_u2_n120 ) );
  NAND2_X1 u2_u4_u2_U69 (.A2( u2_u4_u2_n105 ) , .A1( u2_u4_u2_n106 ) , .ZN( u2_u4_u2_n117 ) );
  AOI21_X1 u2_u4_u2_U7 (.B2( u2_u4_u2_n119 ) , .ZN( u2_u4_u2_n127 ) , .A( u2_u4_u2_n137 ) , .B1( u2_u4_u2_n155 ) );
  NOR2_X1 u2_u4_u2_U70 (.A2( u2_u4_X_16 ) , .ZN( u2_u4_u2_n140 ) , .A1( u2_u4_u2_n166 ) );
  NOR2_X1 u2_u4_u2_U71 (.A2( u2_u4_X_13 ) , .A1( u2_u4_X_14 ) , .ZN( u2_u4_u2_n100 ) );
  NOR2_X1 u2_u4_u2_U72 (.A2( u2_u4_X_16 ) , .A1( u2_u4_X_17 ) , .ZN( u2_u4_u2_n138 ) );
  NOR2_X1 u2_u4_u2_U73 (.A2( u2_u4_X_15 ) , .A1( u2_u4_X_18 ) , .ZN( u2_u4_u2_n104 ) );
  NOR2_X1 u2_u4_u2_U74 (.A2( u2_u4_X_14 ) , .ZN( u2_u4_u2_n103 ) , .A1( u2_u4_u2_n174 ) );
  NOR2_X1 u2_u4_u2_U75 (.A2( u2_u4_X_15 ) , .ZN( u2_u4_u2_n102 ) , .A1( u2_u4_u2_n165 ) );
  NOR2_X1 u2_u4_u2_U76 (.A2( u2_u4_X_17 ) , .ZN( u2_u4_u2_n114 ) , .A1( u2_u4_u2_n169 ) );
  AND2_X1 u2_u4_u2_U77 (.A1( u2_u4_X_15 ) , .ZN( u2_u4_u2_n105 ) , .A2( u2_u4_u2_n165 ) );
  AND2_X1 u2_u4_u2_U78 (.A2( u2_u4_X_15 ) , .A1( u2_u4_X_18 ) , .ZN( u2_u4_u2_n107 ) );
  AND2_X1 u2_u4_u2_U79 (.A1( u2_u4_X_14 ) , .ZN( u2_u4_u2_n106 ) , .A2( u2_u4_u2_n174 ) );
  AOI21_X1 u2_u4_u2_U8 (.ZN( u2_u4_u2_n124 ) , .B1( u2_u4_u2_n131 ) , .B2( u2_u4_u2_n143 ) , .A( u2_u4_u2_n172 ) );
  AND2_X1 u2_u4_u2_U80 (.A1( u2_u4_X_13 ) , .A2( u2_u4_X_14 ) , .ZN( u2_u4_u2_n108 ) );
  INV_X1 u2_u4_u2_U81 (.A( u2_u4_X_16 ) , .ZN( u2_u4_u2_n169 ) );
  INV_X1 u2_u4_u2_U82 (.A( u2_u4_X_17 ) , .ZN( u2_u4_u2_n166 ) );
  INV_X1 u2_u4_u2_U83 (.A( u2_u4_X_13 ) , .ZN( u2_u4_u2_n174 ) );
  INV_X1 u2_u4_u2_U84 (.A( u2_u4_X_18 ) , .ZN( u2_u4_u2_n165 ) );
  NAND4_X1 u2_u4_u2_U85 (.ZN( u2_out4_30 ) , .A4( u2_u4_u2_n147 ) , .A3( u2_u4_u2_n148 ) , .A2( u2_u4_u2_n149 ) , .A1( u2_u4_u2_n187 ) );
  NOR3_X1 u2_u4_u2_U86 (.A3( u2_u4_u2_n144 ) , .A2( u2_u4_u2_n145 ) , .A1( u2_u4_u2_n146 ) , .ZN( u2_u4_u2_n147 ) );
  AOI21_X1 u2_u4_u2_U87 (.B2( u2_u4_u2_n138 ) , .ZN( u2_u4_u2_n148 ) , .A( u2_u4_u2_n162 ) , .B1( u2_u4_u2_n182 ) );
  NAND4_X1 u2_u4_u2_U88 (.ZN( u2_out4_24 ) , .A4( u2_u4_u2_n111 ) , .A3( u2_u4_u2_n112 ) , .A1( u2_u4_u2_n130 ) , .A2( u2_u4_u2_n187 ) );
  AOI221_X1 u2_u4_u2_U89 (.A( u2_u4_u2_n109 ) , .B1( u2_u4_u2_n110 ) , .ZN( u2_u4_u2_n111 ) , .C1( u2_u4_u2_n134 ) , .C2( u2_u4_u2_n170 ) , .B2( u2_u4_u2_n173 ) );
  AOI21_X1 u2_u4_u2_U9 (.B2( u2_u4_u2_n123 ) , .ZN( u2_u4_u2_n125 ) , .A( u2_u4_u2_n171 ) , .B1( u2_u4_u2_n184 ) );
  AOI21_X1 u2_u4_u2_U90 (.ZN( u2_u4_u2_n112 ) , .B2( u2_u4_u2_n156 ) , .A( u2_u4_u2_n164 ) , .B1( u2_u4_u2_n181 ) );
  NAND4_X1 u2_u4_u2_U91 (.ZN( u2_out4_16 ) , .A4( u2_u4_u2_n128 ) , .A3( u2_u4_u2_n129 ) , .A1( u2_u4_u2_n130 ) , .A2( u2_u4_u2_n186 ) );
  AOI22_X1 u2_u4_u2_U92 (.A2( u2_u4_u2_n118 ) , .ZN( u2_u4_u2_n129 ) , .A1( u2_u4_u2_n140 ) , .B1( u2_u4_u2_n157 ) , .B2( u2_u4_u2_n170 ) );
  INV_X1 u2_u4_u2_U93 (.A( u2_u4_u2_n163 ) , .ZN( u2_u4_u2_n186 ) );
  OR4_X1 u2_u4_u2_U94 (.ZN( u2_out4_6 ) , .A4( u2_u4_u2_n161 ) , .A3( u2_u4_u2_n162 ) , .A2( u2_u4_u2_n163 ) , .A1( u2_u4_u2_n164 ) );
  OR3_X1 u2_u4_u2_U95 (.A2( u2_u4_u2_n159 ) , .A1( u2_u4_u2_n160 ) , .ZN( u2_u4_u2_n161 ) , .A3( u2_u4_u2_n183 ) );
  AOI21_X1 u2_u4_u2_U96 (.B2( u2_u4_u2_n154 ) , .B1( u2_u4_u2_n155 ) , .ZN( u2_u4_u2_n159 ) , .A( u2_u4_u2_n167 ) );
  NAND3_X1 u2_u4_u2_U97 (.A2( u2_u4_u2_n117 ) , .A1( u2_u4_u2_n122 ) , .A3( u2_u4_u2_n123 ) , .ZN( u2_u4_u2_n134 ) );
  NAND3_X1 u2_u4_u2_U98 (.ZN( u2_u4_u2_n110 ) , .A2( u2_u4_u2_n131 ) , .A3( u2_u4_u2_n139 ) , .A1( u2_u4_u2_n154 ) );
  NAND3_X1 u2_u4_u2_U99 (.A2( u2_u4_u2_n100 ) , .ZN( u2_u4_u2_n101 ) , .A1( u2_u4_u2_n104 ) , .A3( u2_u4_u2_n114 ) );
  OAI22_X1 u2_u4_u3_U10 (.B1( u2_u4_u3_n113 ) , .A2( u2_u4_u3_n135 ) , .A1( u2_u4_u3_n150 ) , .B2( u2_u4_u3_n164 ) , .ZN( u2_u4_u3_n98 ) );
  OAI211_X1 u2_u4_u3_U11 (.B( u2_u4_u3_n106 ) , .ZN( u2_u4_u3_n119 ) , .C2( u2_u4_u3_n128 ) , .C1( u2_u4_u3_n167 ) , .A( u2_u4_u3_n181 ) );
  AOI221_X1 u2_u4_u3_U12 (.C1( u2_u4_u3_n105 ) , .ZN( u2_u4_u3_n106 ) , .A( u2_u4_u3_n131 ) , .B2( u2_u4_u3_n132 ) , .C2( u2_u4_u3_n133 ) , .B1( u2_u4_u3_n169 ) );
  INV_X1 u2_u4_u3_U13 (.ZN( u2_u4_u3_n181 ) , .A( u2_u4_u3_n98 ) );
  NAND2_X1 u2_u4_u3_U14 (.ZN( u2_u4_u3_n105 ) , .A2( u2_u4_u3_n130 ) , .A1( u2_u4_u3_n155 ) );
  AOI22_X1 u2_u4_u3_U15 (.B1( u2_u4_u3_n115 ) , .A2( u2_u4_u3_n116 ) , .ZN( u2_u4_u3_n123 ) , .B2( u2_u4_u3_n133 ) , .A1( u2_u4_u3_n169 ) );
  NAND2_X1 u2_u4_u3_U16 (.ZN( u2_u4_u3_n116 ) , .A2( u2_u4_u3_n151 ) , .A1( u2_u4_u3_n182 ) );
  NOR2_X1 u2_u4_u3_U17 (.ZN( u2_u4_u3_n126 ) , .A2( u2_u4_u3_n150 ) , .A1( u2_u4_u3_n164 ) );
  AOI21_X1 u2_u4_u3_U18 (.ZN( u2_u4_u3_n112 ) , .B2( u2_u4_u3_n146 ) , .B1( u2_u4_u3_n155 ) , .A( u2_u4_u3_n167 ) );
  NAND2_X1 u2_u4_u3_U19 (.A1( u2_u4_u3_n135 ) , .ZN( u2_u4_u3_n142 ) , .A2( u2_u4_u3_n164 ) );
  NAND2_X1 u2_u4_u3_U20 (.ZN( u2_u4_u3_n132 ) , .A2( u2_u4_u3_n152 ) , .A1( u2_u4_u3_n156 ) );
  AND2_X1 u2_u4_u3_U21 (.A2( u2_u4_u3_n113 ) , .A1( u2_u4_u3_n114 ) , .ZN( u2_u4_u3_n151 ) );
  INV_X1 u2_u4_u3_U22 (.A( u2_u4_u3_n133 ) , .ZN( u2_u4_u3_n165 ) );
  INV_X1 u2_u4_u3_U23 (.A( u2_u4_u3_n135 ) , .ZN( u2_u4_u3_n170 ) );
  NAND2_X1 u2_u4_u3_U24 (.A1( u2_u4_u3_n107 ) , .A2( u2_u4_u3_n108 ) , .ZN( u2_u4_u3_n140 ) );
  NAND2_X1 u2_u4_u3_U25 (.ZN( u2_u4_u3_n117 ) , .A1( u2_u4_u3_n124 ) , .A2( u2_u4_u3_n148 ) );
  NAND2_X1 u2_u4_u3_U26 (.ZN( u2_u4_u3_n143 ) , .A1( u2_u4_u3_n165 ) , .A2( u2_u4_u3_n167 ) );
  INV_X1 u2_u4_u3_U27 (.A( u2_u4_u3_n130 ) , .ZN( u2_u4_u3_n177 ) );
  INV_X1 u2_u4_u3_U28 (.A( u2_u4_u3_n128 ) , .ZN( u2_u4_u3_n176 ) );
  INV_X1 u2_u4_u3_U29 (.A( u2_u4_u3_n155 ) , .ZN( u2_u4_u3_n174 ) );
  INV_X1 u2_u4_u3_U3 (.A( u2_u4_u3_n129 ) , .ZN( u2_u4_u3_n183 ) );
  INV_X1 u2_u4_u3_U30 (.A( u2_u4_u3_n139 ) , .ZN( u2_u4_u3_n185 ) );
  NOR2_X1 u2_u4_u3_U31 (.ZN( u2_u4_u3_n135 ) , .A2( u2_u4_u3_n141 ) , .A1( u2_u4_u3_n169 ) );
  OAI222_X1 u2_u4_u3_U32 (.C2( u2_u4_u3_n107 ) , .A2( u2_u4_u3_n108 ) , .B1( u2_u4_u3_n135 ) , .ZN( u2_u4_u3_n138 ) , .B2( u2_u4_u3_n146 ) , .C1( u2_u4_u3_n154 ) , .A1( u2_u4_u3_n164 ) );
  NOR4_X1 u2_u4_u3_U33 (.A4( u2_u4_u3_n157 ) , .A3( u2_u4_u3_n158 ) , .A2( u2_u4_u3_n159 ) , .A1( u2_u4_u3_n160 ) , .ZN( u2_u4_u3_n161 ) );
  AOI21_X1 u2_u4_u3_U34 (.B2( u2_u4_u3_n152 ) , .B1( u2_u4_u3_n153 ) , .ZN( u2_u4_u3_n158 ) , .A( u2_u4_u3_n164 ) );
  AOI21_X1 u2_u4_u3_U35 (.A( u2_u4_u3_n149 ) , .B2( u2_u4_u3_n150 ) , .B1( u2_u4_u3_n151 ) , .ZN( u2_u4_u3_n159 ) );
  AOI21_X1 u2_u4_u3_U36 (.A( u2_u4_u3_n154 ) , .B2( u2_u4_u3_n155 ) , .B1( u2_u4_u3_n156 ) , .ZN( u2_u4_u3_n157 ) );
  AOI211_X1 u2_u4_u3_U37 (.ZN( u2_u4_u3_n109 ) , .A( u2_u4_u3_n119 ) , .C2( u2_u4_u3_n129 ) , .B( u2_u4_u3_n138 ) , .C1( u2_u4_u3_n141 ) );
  AOI211_X1 u2_u4_u3_U38 (.B( u2_u4_u3_n119 ) , .A( u2_u4_u3_n120 ) , .C2( u2_u4_u3_n121 ) , .ZN( u2_u4_u3_n122 ) , .C1( u2_u4_u3_n179 ) );
  INV_X1 u2_u4_u3_U39 (.A( u2_u4_u3_n156 ) , .ZN( u2_u4_u3_n179 ) );
  INV_X1 u2_u4_u3_U4 (.A( u2_u4_u3_n140 ) , .ZN( u2_u4_u3_n182 ) );
  OAI22_X1 u2_u4_u3_U40 (.B1( u2_u4_u3_n118 ) , .ZN( u2_u4_u3_n120 ) , .A1( u2_u4_u3_n135 ) , .B2( u2_u4_u3_n154 ) , .A2( u2_u4_u3_n178 ) );
  AND3_X1 u2_u4_u3_U41 (.ZN( u2_u4_u3_n118 ) , .A2( u2_u4_u3_n124 ) , .A1( u2_u4_u3_n144 ) , .A3( u2_u4_u3_n152 ) );
  INV_X1 u2_u4_u3_U42 (.A( u2_u4_u3_n121 ) , .ZN( u2_u4_u3_n164 ) );
  NAND2_X1 u2_u4_u3_U43 (.ZN( u2_u4_u3_n133 ) , .A1( u2_u4_u3_n154 ) , .A2( u2_u4_u3_n164 ) );
  OAI211_X1 u2_u4_u3_U44 (.B( u2_u4_u3_n127 ) , .ZN( u2_u4_u3_n139 ) , .C1( u2_u4_u3_n150 ) , .C2( u2_u4_u3_n154 ) , .A( u2_u4_u3_n184 ) );
  INV_X1 u2_u4_u3_U45 (.A( u2_u4_u3_n125 ) , .ZN( u2_u4_u3_n184 ) );
  AOI221_X1 u2_u4_u3_U46 (.A( u2_u4_u3_n126 ) , .ZN( u2_u4_u3_n127 ) , .C2( u2_u4_u3_n132 ) , .C1( u2_u4_u3_n169 ) , .B2( u2_u4_u3_n170 ) , .B1( u2_u4_u3_n174 ) );
  OAI22_X1 u2_u4_u3_U47 (.A1( u2_u4_u3_n124 ) , .ZN( u2_u4_u3_n125 ) , .B2( u2_u4_u3_n145 ) , .A2( u2_u4_u3_n165 ) , .B1( u2_u4_u3_n167 ) );
  NOR2_X1 u2_u4_u3_U48 (.A1( u2_u4_u3_n113 ) , .ZN( u2_u4_u3_n131 ) , .A2( u2_u4_u3_n154 ) );
  NAND2_X1 u2_u4_u3_U49 (.A1( u2_u4_u3_n103 ) , .ZN( u2_u4_u3_n150 ) , .A2( u2_u4_u3_n99 ) );
  INV_X1 u2_u4_u3_U5 (.A( u2_u4_u3_n117 ) , .ZN( u2_u4_u3_n178 ) );
  NAND2_X1 u2_u4_u3_U50 (.A2( u2_u4_u3_n102 ) , .ZN( u2_u4_u3_n155 ) , .A1( u2_u4_u3_n97 ) );
  INV_X1 u2_u4_u3_U51 (.A( u2_u4_u3_n141 ) , .ZN( u2_u4_u3_n167 ) );
  AOI21_X1 u2_u4_u3_U52 (.B2( u2_u4_u3_n114 ) , .B1( u2_u4_u3_n146 ) , .A( u2_u4_u3_n154 ) , .ZN( u2_u4_u3_n94 ) );
  AOI21_X1 u2_u4_u3_U53 (.ZN( u2_u4_u3_n110 ) , .B2( u2_u4_u3_n142 ) , .B1( u2_u4_u3_n186 ) , .A( u2_u4_u3_n95 ) );
  INV_X1 u2_u4_u3_U54 (.A( u2_u4_u3_n145 ) , .ZN( u2_u4_u3_n186 ) );
  AOI21_X1 u2_u4_u3_U55 (.B1( u2_u4_u3_n124 ) , .A( u2_u4_u3_n149 ) , .B2( u2_u4_u3_n155 ) , .ZN( u2_u4_u3_n95 ) );
  INV_X1 u2_u4_u3_U56 (.A( u2_u4_u3_n149 ) , .ZN( u2_u4_u3_n169 ) );
  NAND2_X1 u2_u4_u3_U57 (.ZN( u2_u4_u3_n124 ) , .A1( u2_u4_u3_n96 ) , .A2( u2_u4_u3_n97 ) );
  NAND2_X1 u2_u4_u3_U58 (.A2( u2_u4_u3_n100 ) , .ZN( u2_u4_u3_n146 ) , .A1( u2_u4_u3_n96 ) );
  NAND2_X1 u2_u4_u3_U59 (.A1( u2_u4_u3_n101 ) , .ZN( u2_u4_u3_n145 ) , .A2( u2_u4_u3_n99 ) );
  AOI221_X1 u2_u4_u3_U6 (.A( u2_u4_u3_n131 ) , .C2( u2_u4_u3_n132 ) , .C1( u2_u4_u3_n133 ) , .ZN( u2_u4_u3_n134 ) , .B1( u2_u4_u3_n143 ) , .B2( u2_u4_u3_n177 ) );
  NAND2_X1 u2_u4_u3_U60 (.A1( u2_u4_u3_n100 ) , .ZN( u2_u4_u3_n156 ) , .A2( u2_u4_u3_n99 ) );
  NAND2_X1 u2_u4_u3_U61 (.A2( u2_u4_u3_n101 ) , .A1( u2_u4_u3_n104 ) , .ZN( u2_u4_u3_n148 ) );
  NAND2_X1 u2_u4_u3_U62 (.A1( u2_u4_u3_n100 ) , .A2( u2_u4_u3_n102 ) , .ZN( u2_u4_u3_n128 ) );
  NAND2_X1 u2_u4_u3_U63 (.A2( u2_u4_u3_n101 ) , .A1( u2_u4_u3_n102 ) , .ZN( u2_u4_u3_n152 ) );
  NAND2_X1 u2_u4_u3_U64 (.A2( u2_u4_u3_n101 ) , .ZN( u2_u4_u3_n114 ) , .A1( u2_u4_u3_n96 ) );
  NAND2_X1 u2_u4_u3_U65 (.ZN( u2_u4_u3_n107 ) , .A1( u2_u4_u3_n97 ) , .A2( u2_u4_u3_n99 ) );
  NAND2_X1 u2_u4_u3_U66 (.A2( u2_u4_u3_n100 ) , .A1( u2_u4_u3_n104 ) , .ZN( u2_u4_u3_n113 ) );
  NAND2_X1 u2_u4_u3_U67 (.A1( u2_u4_u3_n104 ) , .ZN( u2_u4_u3_n153 ) , .A2( u2_u4_u3_n97 ) );
  NAND2_X1 u2_u4_u3_U68 (.A2( u2_u4_u3_n103 ) , .A1( u2_u4_u3_n104 ) , .ZN( u2_u4_u3_n130 ) );
  NAND2_X1 u2_u4_u3_U69 (.A2( u2_u4_u3_n103 ) , .ZN( u2_u4_u3_n144 ) , .A1( u2_u4_u3_n96 ) );
  OAI22_X1 u2_u4_u3_U7 (.B2( u2_u4_u3_n147 ) , .A2( u2_u4_u3_n148 ) , .ZN( u2_u4_u3_n160 ) , .B1( u2_u4_u3_n165 ) , .A1( u2_u4_u3_n168 ) );
  NAND2_X1 u2_u4_u3_U70 (.A1( u2_u4_u3_n102 ) , .A2( u2_u4_u3_n103 ) , .ZN( u2_u4_u3_n108 ) );
  NOR2_X1 u2_u4_u3_U71 (.A2( u2_u4_X_19 ) , .A1( u2_u4_X_20 ) , .ZN( u2_u4_u3_n99 ) );
  NOR2_X1 u2_u4_u3_U72 (.A2( u2_u4_X_21 ) , .A1( u2_u4_X_24 ) , .ZN( u2_u4_u3_n103 ) );
  NOR2_X1 u2_u4_u3_U73 (.A2( u2_u4_X_24 ) , .A1( u2_u4_u3_n171 ) , .ZN( u2_u4_u3_n97 ) );
  NOR2_X1 u2_u4_u3_U74 (.A2( u2_u4_X_23 ) , .ZN( u2_u4_u3_n141 ) , .A1( u2_u4_u3_n166 ) );
  NOR2_X1 u2_u4_u3_U75 (.A2( u2_u4_X_19 ) , .A1( u2_u4_u3_n172 ) , .ZN( u2_u4_u3_n96 ) );
  NAND2_X1 u2_u4_u3_U76 (.A1( u2_u4_X_22 ) , .A2( u2_u4_X_23 ) , .ZN( u2_u4_u3_n154 ) );
  NAND2_X1 u2_u4_u3_U77 (.A1( u2_u4_X_23 ) , .ZN( u2_u4_u3_n149 ) , .A2( u2_u4_u3_n166 ) );
  NOR2_X1 u2_u4_u3_U78 (.A2( u2_u4_X_22 ) , .A1( u2_u4_X_23 ) , .ZN( u2_u4_u3_n121 ) );
  AND2_X1 u2_u4_u3_U79 (.A1( u2_u4_X_24 ) , .ZN( u2_u4_u3_n101 ) , .A2( u2_u4_u3_n171 ) );
  AND3_X1 u2_u4_u3_U8 (.A3( u2_u4_u3_n144 ) , .A2( u2_u4_u3_n145 ) , .A1( u2_u4_u3_n146 ) , .ZN( u2_u4_u3_n147 ) );
  AND2_X1 u2_u4_u3_U80 (.A1( u2_u4_X_19 ) , .ZN( u2_u4_u3_n102 ) , .A2( u2_u4_u3_n172 ) );
  AND2_X1 u2_u4_u3_U81 (.A1( u2_u4_X_21 ) , .A2( u2_u4_X_24 ) , .ZN( u2_u4_u3_n100 ) );
  AND2_X1 u2_u4_u3_U82 (.A2( u2_u4_X_19 ) , .A1( u2_u4_X_20 ) , .ZN( u2_u4_u3_n104 ) );
  INV_X1 u2_u4_u3_U83 (.A( u2_u4_X_22 ) , .ZN( u2_u4_u3_n166 ) );
  INV_X1 u2_u4_u3_U84 (.A( u2_u4_X_21 ) , .ZN( u2_u4_u3_n171 ) );
  INV_X1 u2_u4_u3_U85 (.A( u2_u4_X_20 ) , .ZN( u2_u4_u3_n172 ) );
  OR4_X1 u2_u4_u3_U86 (.ZN( u2_out4_10 ) , .A4( u2_u4_u3_n136 ) , .A3( u2_u4_u3_n137 ) , .A1( u2_u4_u3_n138 ) , .A2( u2_u4_u3_n139 ) );
  OAI222_X1 u2_u4_u3_U87 (.C1( u2_u4_u3_n128 ) , .ZN( u2_u4_u3_n137 ) , .B1( u2_u4_u3_n148 ) , .A2( u2_u4_u3_n150 ) , .B2( u2_u4_u3_n154 ) , .C2( u2_u4_u3_n164 ) , .A1( u2_u4_u3_n167 ) );
  OAI221_X1 u2_u4_u3_U88 (.A( u2_u4_u3_n134 ) , .B2( u2_u4_u3_n135 ) , .ZN( u2_u4_u3_n136 ) , .C1( u2_u4_u3_n149 ) , .B1( u2_u4_u3_n151 ) , .C2( u2_u4_u3_n183 ) );
  NAND4_X1 u2_u4_u3_U89 (.ZN( u2_out4_26 ) , .A4( u2_u4_u3_n109 ) , .A3( u2_u4_u3_n110 ) , .A2( u2_u4_u3_n111 ) , .A1( u2_u4_u3_n173 ) );
  INV_X1 u2_u4_u3_U9 (.A( u2_u4_u3_n143 ) , .ZN( u2_u4_u3_n168 ) );
  INV_X1 u2_u4_u3_U90 (.ZN( u2_u4_u3_n173 ) , .A( u2_u4_u3_n94 ) );
  OAI21_X1 u2_u4_u3_U91 (.ZN( u2_u4_u3_n111 ) , .B2( u2_u4_u3_n117 ) , .A( u2_u4_u3_n133 ) , .B1( u2_u4_u3_n176 ) );
  NAND4_X1 u2_u4_u3_U92 (.ZN( u2_out4_20 ) , .A4( u2_u4_u3_n122 ) , .A3( u2_u4_u3_n123 ) , .A1( u2_u4_u3_n175 ) , .A2( u2_u4_u3_n180 ) );
  INV_X1 u2_u4_u3_U93 (.A( u2_u4_u3_n126 ) , .ZN( u2_u4_u3_n180 ) );
  INV_X1 u2_u4_u3_U94 (.A( u2_u4_u3_n112 ) , .ZN( u2_u4_u3_n175 ) );
  NAND4_X1 u2_u4_u3_U95 (.ZN( u2_out4_1 ) , .A4( u2_u4_u3_n161 ) , .A3( u2_u4_u3_n162 ) , .A2( u2_u4_u3_n163 ) , .A1( u2_u4_u3_n185 ) );
  NAND2_X1 u2_u4_u3_U96 (.ZN( u2_u4_u3_n163 ) , .A2( u2_u4_u3_n170 ) , .A1( u2_u4_u3_n176 ) );
  AOI22_X1 u2_u4_u3_U97 (.B2( u2_u4_u3_n140 ) , .B1( u2_u4_u3_n141 ) , .A2( u2_u4_u3_n142 ) , .ZN( u2_u4_u3_n162 ) , .A1( u2_u4_u3_n177 ) );
  NAND3_X1 u2_u4_u3_U98 (.A1( u2_u4_u3_n114 ) , .ZN( u2_u4_u3_n115 ) , .A2( u2_u4_u3_n145 ) , .A3( u2_u4_u3_n153 ) );
  NAND3_X1 u2_u4_u3_U99 (.ZN( u2_u4_u3_n129 ) , .A2( u2_u4_u3_n144 ) , .A1( u2_u4_u3_n153 ) , .A3( u2_u4_u3_n182 ) );
  XOR2_X1 u2_u5_U26 (.B( u2_K6_30 ) , .A( u2_R4_21 ) , .Z( u2_u5_X_30 ) );
  XOR2_X1 u2_u5_U28 (.B( u2_K6_29 ) , .A( u2_R4_20 ) , .Z( u2_u5_X_29 ) );
  XOR2_X1 u2_u5_U29 (.B( u2_K6_28 ) , .A( u2_R4_19 ) , .Z( u2_u5_X_28 ) );
  XOR2_X1 u2_u5_U30 (.B( u2_K6_27 ) , .A( u2_R4_18 ) , .Z( u2_u5_X_27 ) );
  XOR2_X1 u2_u5_U31 (.B( u2_K6_26 ) , .A( u2_R4_17 ) , .Z( u2_u5_X_26 ) );
  XOR2_X1 u2_u5_U32 (.B( u2_K6_25 ) , .A( u2_R4_16 ) , .Z( u2_u5_X_25 ) );
  XOR2_X1 u2_u5_U33 (.B( u2_K6_24 ) , .A( u2_R4_17 ) , .Z( u2_u5_X_24 ) );
  XOR2_X1 u2_u5_U34 (.B( u2_K6_23 ) , .A( u2_R4_16 ) , .Z( u2_u5_X_23 ) );
  XOR2_X1 u2_u5_U35 (.B( u2_K6_22 ) , .A( u2_R4_15 ) , .Z( u2_u5_X_22 ) );
  XOR2_X1 u2_u5_U36 (.B( u2_K6_21 ) , .A( u2_R4_14 ) , .Z( u2_u5_X_21 ) );
  XOR2_X1 u2_u5_U37 (.B( u2_K6_20 ) , .A( u2_R4_13 ) , .Z( u2_u5_X_20 ) );
  XOR2_X1 u2_u5_U39 (.B( u2_K6_19 ) , .A( u2_R4_12 ) , .Z( u2_u5_X_19 ) );
  OAI22_X1 u2_u5_u3_U10 (.B1( u2_u5_u3_n113 ) , .A2( u2_u5_u3_n135 ) , .A1( u2_u5_u3_n150 ) , .B2( u2_u5_u3_n164 ) , .ZN( u2_u5_u3_n98 ) );
  OAI211_X1 u2_u5_u3_U11 (.B( u2_u5_u3_n106 ) , .ZN( u2_u5_u3_n119 ) , .C2( u2_u5_u3_n128 ) , .C1( u2_u5_u3_n167 ) , .A( u2_u5_u3_n181 ) );
  AOI221_X1 u2_u5_u3_U12 (.C1( u2_u5_u3_n105 ) , .ZN( u2_u5_u3_n106 ) , .A( u2_u5_u3_n131 ) , .B2( u2_u5_u3_n132 ) , .C2( u2_u5_u3_n133 ) , .B1( u2_u5_u3_n169 ) );
  INV_X1 u2_u5_u3_U13 (.ZN( u2_u5_u3_n181 ) , .A( u2_u5_u3_n98 ) );
  NAND2_X1 u2_u5_u3_U14 (.ZN( u2_u5_u3_n105 ) , .A2( u2_u5_u3_n130 ) , .A1( u2_u5_u3_n155 ) );
  AOI22_X1 u2_u5_u3_U15 (.B1( u2_u5_u3_n115 ) , .A2( u2_u5_u3_n116 ) , .ZN( u2_u5_u3_n123 ) , .B2( u2_u5_u3_n133 ) , .A1( u2_u5_u3_n169 ) );
  NAND2_X1 u2_u5_u3_U16 (.ZN( u2_u5_u3_n116 ) , .A2( u2_u5_u3_n151 ) , .A1( u2_u5_u3_n182 ) );
  NOR2_X1 u2_u5_u3_U17 (.ZN( u2_u5_u3_n126 ) , .A2( u2_u5_u3_n150 ) , .A1( u2_u5_u3_n164 ) );
  AOI21_X1 u2_u5_u3_U18 (.ZN( u2_u5_u3_n112 ) , .B2( u2_u5_u3_n146 ) , .B1( u2_u5_u3_n155 ) , .A( u2_u5_u3_n167 ) );
  NAND2_X1 u2_u5_u3_U19 (.A1( u2_u5_u3_n135 ) , .ZN( u2_u5_u3_n142 ) , .A2( u2_u5_u3_n164 ) );
  NAND2_X1 u2_u5_u3_U20 (.ZN( u2_u5_u3_n132 ) , .A2( u2_u5_u3_n152 ) , .A1( u2_u5_u3_n156 ) );
  AND2_X1 u2_u5_u3_U21 (.A2( u2_u5_u3_n113 ) , .A1( u2_u5_u3_n114 ) , .ZN( u2_u5_u3_n151 ) );
  INV_X1 u2_u5_u3_U22 (.A( u2_u5_u3_n133 ) , .ZN( u2_u5_u3_n165 ) );
  INV_X1 u2_u5_u3_U23 (.A( u2_u5_u3_n135 ) , .ZN( u2_u5_u3_n170 ) );
  NAND2_X1 u2_u5_u3_U24 (.A1( u2_u5_u3_n107 ) , .A2( u2_u5_u3_n108 ) , .ZN( u2_u5_u3_n140 ) );
  NAND2_X1 u2_u5_u3_U25 (.ZN( u2_u5_u3_n117 ) , .A1( u2_u5_u3_n124 ) , .A2( u2_u5_u3_n148 ) );
  NAND2_X1 u2_u5_u3_U26 (.ZN( u2_u5_u3_n143 ) , .A1( u2_u5_u3_n165 ) , .A2( u2_u5_u3_n167 ) );
  INV_X1 u2_u5_u3_U27 (.A( u2_u5_u3_n130 ) , .ZN( u2_u5_u3_n177 ) );
  INV_X1 u2_u5_u3_U28 (.A( u2_u5_u3_n128 ) , .ZN( u2_u5_u3_n176 ) );
  INV_X1 u2_u5_u3_U29 (.A( u2_u5_u3_n155 ) , .ZN( u2_u5_u3_n174 ) );
  INV_X1 u2_u5_u3_U3 (.A( u2_u5_u3_n129 ) , .ZN( u2_u5_u3_n183 ) );
  INV_X1 u2_u5_u3_U30 (.A( u2_u5_u3_n139 ) , .ZN( u2_u5_u3_n185 ) );
  NOR2_X1 u2_u5_u3_U31 (.ZN( u2_u5_u3_n135 ) , .A2( u2_u5_u3_n141 ) , .A1( u2_u5_u3_n169 ) );
  OAI222_X1 u2_u5_u3_U32 (.C2( u2_u5_u3_n107 ) , .A2( u2_u5_u3_n108 ) , .B1( u2_u5_u3_n135 ) , .ZN( u2_u5_u3_n138 ) , .B2( u2_u5_u3_n146 ) , .C1( u2_u5_u3_n154 ) , .A1( u2_u5_u3_n164 ) );
  NOR4_X1 u2_u5_u3_U33 (.A4( u2_u5_u3_n157 ) , .A3( u2_u5_u3_n158 ) , .A2( u2_u5_u3_n159 ) , .A1( u2_u5_u3_n160 ) , .ZN( u2_u5_u3_n161 ) );
  AOI21_X1 u2_u5_u3_U34 (.B2( u2_u5_u3_n152 ) , .B1( u2_u5_u3_n153 ) , .ZN( u2_u5_u3_n158 ) , .A( u2_u5_u3_n164 ) );
  AOI21_X1 u2_u5_u3_U35 (.A( u2_u5_u3_n154 ) , .B2( u2_u5_u3_n155 ) , .B1( u2_u5_u3_n156 ) , .ZN( u2_u5_u3_n157 ) );
  AOI21_X1 u2_u5_u3_U36 (.A( u2_u5_u3_n149 ) , .B2( u2_u5_u3_n150 ) , .B1( u2_u5_u3_n151 ) , .ZN( u2_u5_u3_n159 ) );
  AOI211_X1 u2_u5_u3_U37 (.ZN( u2_u5_u3_n109 ) , .A( u2_u5_u3_n119 ) , .C2( u2_u5_u3_n129 ) , .B( u2_u5_u3_n138 ) , .C1( u2_u5_u3_n141 ) );
  AOI211_X1 u2_u5_u3_U38 (.B( u2_u5_u3_n119 ) , .A( u2_u5_u3_n120 ) , .C2( u2_u5_u3_n121 ) , .ZN( u2_u5_u3_n122 ) , .C1( u2_u5_u3_n179 ) );
  INV_X1 u2_u5_u3_U39 (.A( u2_u5_u3_n156 ) , .ZN( u2_u5_u3_n179 ) );
  INV_X1 u2_u5_u3_U4 (.A( u2_u5_u3_n140 ) , .ZN( u2_u5_u3_n182 ) );
  OAI22_X1 u2_u5_u3_U40 (.B1( u2_u5_u3_n118 ) , .ZN( u2_u5_u3_n120 ) , .A1( u2_u5_u3_n135 ) , .B2( u2_u5_u3_n154 ) , .A2( u2_u5_u3_n178 ) );
  AND3_X1 u2_u5_u3_U41 (.ZN( u2_u5_u3_n118 ) , .A2( u2_u5_u3_n124 ) , .A1( u2_u5_u3_n144 ) , .A3( u2_u5_u3_n152 ) );
  INV_X1 u2_u5_u3_U42 (.A( u2_u5_u3_n121 ) , .ZN( u2_u5_u3_n164 ) );
  NAND2_X1 u2_u5_u3_U43 (.ZN( u2_u5_u3_n133 ) , .A1( u2_u5_u3_n154 ) , .A2( u2_u5_u3_n164 ) );
  OAI211_X1 u2_u5_u3_U44 (.B( u2_u5_u3_n127 ) , .ZN( u2_u5_u3_n139 ) , .C1( u2_u5_u3_n150 ) , .C2( u2_u5_u3_n154 ) , .A( u2_u5_u3_n184 ) );
  INV_X1 u2_u5_u3_U45 (.A( u2_u5_u3_n125 ) , .ZN( u2_u5_u3_n184 ) );
  AOI221_X1 u2_u5_u3_U46 (.A( u2_u5_u3_n126 ) , .ZN( u2_u5_u3_n127 ) , .C2( u2_u5_u3_n132 ) , .C1( u2_u5_u3_n169 ) , .B2( u2_u5_u3_n170 ) , .B1( u2_u5_u3_n174 ) );
  OAI22_X1 u2_u5_u3_U47 (.A1( u2_u5_u3_n124 ) , .ZN( u2_u5_u3_n125 ) , .B2( u2_u5_u3_n145 ) , .A2( u2_u5_u3_n165 ) , .B1( u2_u5_u3_n167 ) );
  NOR2_X1 u2_u5_u3_U48 (.A1( u2_u5_u3_n113 ) , .ZN( u2_u5_u3_n131 ) , .A2( u2_u5_u3_n154 ) );
  NAND2_X1 u2_u5_u3_U49 (.A1( u2_u5_u3_n103 ) , .ZN( u2_u5_u3_n150 ) , .A2( u2_u5_u3_n99 ) );
  INV_X1 u2_u5_u3_U5 (.A( u2_u5_u3_n117 ) , .ZN( u2_u5_u3_n178 ) );
  NAND2_X1 u2_u5_u3_U50 (.A2( u2_u5_u3_n102 ) , .ZN( u2_u5_u3_n155 ) , .A1( u2_u5_u3_n97 ) );
  INV_X1 u2_u5_u3_U51 (.A( u2_u5_u3_n141 ) , .ZN( u2_u5_u3_n167 ) );
  AOI21_X1 u2_u5_u3_U52 (.B2( u2_u5_u3_n114 ) , .B1( u2_u5_u3_n146 ) , .A( u2_u5_u3_n154 ) , .ZN( u2_u5_u3_n94 ) );
  AOI21_X1 u2_u5_u3_U53 (.ZN( u2_u5_u3_n110 ) , .B2( u2_u5_u3_n142 ) , .B1( u2_u5_u3_n186 ) , .A( u2_u5_u3_n95 ) );
  INV_X1 u2_u5_u3_U54 (.A( u2_u5_u3_n145 ) , .ZN( u2_u5_u3_n186 ) );
  AOI21_X1 u2_u5_u3_U55 (.B1( u2_u5_u3_n124 ) , .A( u2_u5_u3_n149 ) , .B2( u2_u5_u3_n155 ) , .ZN( u2_u5_u3_n95 ) );
  INV_X1 u2_u5_u3_U56 (.A( u2_u5_u3_n149 ) , .ZN( u2_u5_u3_n169 ) );
  NAND2_X1 u2_u5_u3_U57 (.ZN( u2_u5_u3_n124 ) , .A1( u2_u5_u3_n96 ) , .A2( u2_u5_u3_n97 ) );
  NAND2_X1 u2_u5_u3_U58 (.A2( u2_u5_u3_n100 ) , .ZN( u2_u5_u3_n146 ) , .A1( u2_u5_u3_n96 ) );
  NAND2_X1 u2_u5_u3_U59 (.A1( u2_u5_u3_n101 ) , .ZN( u2_u5_u3_n145 ) , .A2( u2_u5_u3_n99 ) );
  AOI221_X1 u2_u5_u3_U6 (.A( u2_u5_u3_n131 ) , .C2( u2_u5_u3_n132 ) , .C1( u2_u5_u3_n133 ) , .ZN( u2_u5_u3_n134 ) , .B1( u2_u5_u3_n143 ) , .B2( u2_u5_u3_n177 ) );
  NAND2_X1 u2_u5_u3_U60 (.A1( u2_u5_u3_n100 ) , .ZN( u2_u5_u3_n156 ) , .A2( u2_u5_u3_n99 ) );
  NAND2_X1 u2_u5_u3_U61 (.A2( u2_u5_u3_n101 ) , .A1( u2_u5_u3_n104 ) , .ZN( u2_u5_u3_n148 ) );
  NAND2_X1 u2_u5_u3_U62 (.A1( u2_u5_u3_n100 ) , .A2( u2_u5_u3_n102 ) , .ZN( u2_u5_u3_n128 ) );
  NAND2_X1 u2_u5_u3_U63 (.A2( u2_u5_u3_n101 ) , .A1( u2_u5_u3_n102 ) , .ZN( u2_u5_u3_n152 ) );
  NAND2_X1 u2_u5_u3_U64 (.A2( u2_u5_u3_n101 ) , .ZN( u2_u5_u3_n114 ) , .A1( u2_u5_u3_n96 ) );
  NAND2_X1 u2_u5_u3_U65 (.ZN( u2_u5_u3_n107 ) , .A1( u2_u5_u3_n97 ) , .A2( u2_u5_u3_n99 ) );
  NAND2_X1 u2_u5_u3_U66 (.A2( u2_u5_u3_n100 ) , .A1( u2_u5_u3_n104 ) , .ZN( u2_u5_u3_n113 ) );
  NAND2_X1 u2_u5_u3_U67 (.A1( u2_u5_u3_n104 ) , .ZN( u2_u5_u3_n153 ) , .A2( u2_u5_u3_n97 ) );
  NAND2_X1 u2_u5_u3_U68 (.A2( u2_u5_u3_n103 ) , .A1( u2_u5_u3_n104 ) , .ZN( u2_u5_u3_n130 ) );
  NAND2_X1 u2_u5_u3_U69 (.A2( u2_u5_u3_n103 ) , .ZN( u2_u5_u3_n144 ) , .A1( u2_u5_u3_n96 ) );
  OAI22_X1 u2_u5_u3_U7 (.B2( u2_u5_u3_n147 ) , .A2( u2_u5_u3_n148 ) , .ZN( u2_u5_u3_n160 ) , .B1( u2_u5_u3_n165 ) , .A1( u2_u5_u3_n168 ) );
  NAND2_X1 u2_u5_u3_U70 (.A1( u2_u5_u3_n102 ) , .A2( u2_u5_u3_n103 ) , .ZN( u2_u5_u3_n108 ) );
  NOR2_X1 u2_u5_u3_U71 (.A2( u2_u5_X_19 ) , .A1( u2_u5_X_20 ) , .ZN( u2_u5_u3_n99 ) );
  NOR2_X1 u2_u5_u3_U72 (.A2( u2_u5_X_21 ) , .A1( u2_u5_X_24 ) , .ZN( u2_u5_u3_n103 ) );
  NOR2_X1 u2_u5_u3_U73 (.A2( u2_u5_X_24 ) , .A1( u2_u5_u3_n171 ) , .ZN( u2_u5_u3_n97 ) );
  NOR2_X1 u2_u5_u3_U74 (.A2( u2_u5_X_23 ) , .ZN( u2_u5_u3_n141 ) , .A1( u2_u5_u3_n166 ) );
  NOR2_X1 u2_u5_u3_U75 (.A2( u2_u5_X_19 ) , .A1( u2_u5_u3_n172 ) , .ZN( u2_u5_u3_n96 ) );
  NAND2_X1 u2_u5_u3_U76 (.A1( u2_u5_X_22 ) , .A2( u2_u5_X_23 ) , .ZN( u2_u5_u3_n154 ) );
  NAND2_X1 u2_u5_u3_U77 (.A1( u2_u5_X_23 ) , .ZN( u2_u5_u3_n149 ) , .A2( u2_u5_u3_n166 ) );
  NOR2_X1 u2_u5_u3_U78 (.A2( u2_u5_X_22 ) , .A1( u2_u5_X_23 ) , .ZN( u2_u5_u3_n121 ) );
  AND2_X1 u2_u5_u3_U79 (.A1( u2_u5_X_24 ) , .ZN( u2_u5_u3_n101 ) , .A2( u2_u5_u3_n171 ) );
  AND3_X1 u2_u5_u3_U8 (.A3( u2_u5_u3_n144 ) , .A2( u2_u5_u3_n145 ) , .A1( u2_u5_u3_n146 ) , .ZN( u2_u5_u3_n147 ) );
  AND2_X1 u2_u5_u3_U80 (.A1( u2_u5_X_19 ) , .ZN( u2_u5_u3_n102 ) , .A2( u2_u5_u3_n172 ) );
  AND2_X1 u2_u5_u3_U81 (.A1( u2_u5_X_21 ) , .A2( u2_u5_X_24 ) , .ZN( u2_u5_u3_n100 ) );
  AND2_X1 u2_u5_u3_U82 (.A2( u2_u5_X_19 ) , .A1( u2_u5_X_20 ) , .ZN( u2_u5_u3_n104 ) );
  INV_X1 u2_u5_u3_U83 (.A( u2_u5_X_22 ) , .ZN( u2_u5_u3_n166 ) );
  INV_X1 u2_u5_u3_U84 (.A( u2_u5_X_21 ) , .ZN( u2_u5_u3_n171 ) );
  INV_X1 u2_u5_u3_U85 (.A( u2_u5_X_20 ) , .ZN( u2_u5_u3_n172 ) );
  NAND4_X1 u2_u5_u3_U86 (.ZN( u2_out5_26 ) , .A4( u2_u5_u3_n109 ) , .A3( u2_u5_u3_n110 ) , .A2( u2_u5_u3_n111 ) , .A1( u2_u5_u3_n173 ) );
  INV_X1 u2_u5_u3_U87 (.ZN( u2_u5_u3_n173 ) , .A( u2_u5_u3_n94 ) );
  OAI21_X1 u2_u5_u3_U88 (.ZN( u2_u5_u3_n111 ) , .B2( u2_u5_u3_n117 ) , .A( u2_u5_u3_n133 ) , .B1( u2_u5_u3_n176 ) );
  NAND4_X1 u2_u5_u3_U89 (.ZN( u2_out5_20 ) , .A4( u2_u5_u3_n122 ) , .A3( u2_u5_u3_n123 ) , .A1( u2_u5_u3_n175 ) , .A2( u2_u5_u3_n180 ) );
  INV_X1 u2_u5_u3_U9 (.A( u2_u5_u3_n143 ) , .ZN( u2_u5_u3_n168 ) );
  INV_X1 u2_u5_u3_U90 (.A( u2_u5_u3_n126 ) , .ZN( u2_u5_u3_n180 ) );
  INV_X1 u2_u5_u3_U91 (.A( u2_u5_u3_n112 ) , .ZN( u2_u5_u3_n175 ) );
  NAND4_X1 u2_u5_u3_U92 (.ZN( u2_out5_1 ) , .A4( u2_u5_u3_n161 ) , .A3( u2_u5_u3_n162 ) , .A2( u2_u5_u3_n163 ) , .A1( u2_u5_u3_n185 ) );
  NAND2_X1 u2_u5_u3_U93 (.ZN( u2_u5_u3_n163 ) , .A2( u2_u5_u3_n170 ) , .A1( u2_u5_u3_n176 ) );
  AOI22_X1 u2_u5_u3_U94 (.B2( u2_u5_u3_n140 ) , .B1( u2_u5_u3_n141 ) , .A2( u2_u5_u3_n142 ) , .ZN( u2_u5_u3_n162 ) , .A1( u2_u5_u3_n177 ) );
  OR4_X1 u2_u5_u3_U95 (.ZN( u2_out5_10 ) , .A4( u2_u5_u3_n136 ) , .A3( u2_u5_u3_n137 ) , .A1( u2_u5_u3_n138 ) , .A2( u2_u5_u3_n139 ) );
  OAI222_X1 u2_u5_u3_U96 (.C1( u2_u5_u3_n128 ) , .ZN( u2_u5_u3_n137 ) , .B1( u2_u5_u3_n148 ) , .A2( u2_u5_u3_n150 ) , .B2( u2_u5_u3_n154 ) , .C2( u2_u5_u3_n164 ) , .A1( u2_u5_u3_n167 ) );
  OAI221_X1 u2_u5_u3_U97 (.A( u2_u5_u3_n134 ) , .B2( u2_u5_u3_n135 ) , .ZN( u2_u5_u3_n136 ) , .C1( u2_u5_u3_n149 ) , .B1( u2_u5_u3_n151 ) , .C2( u2_u5_u3_n183 ) );
  NAND3_X1 u2_u5_u3_U98 (.A1( u2_u5_u3_n114 ) , .ZN( u2_u5_u3_n115 ) , .A2( u2_u5_u3_n145 ) , .A3( u2_u5_u3_n153 ) );
  NAND3_X1 u2_u5_u3_U99 (.ZN( u2_u5_u3_n129 ) , .A2( u2_u5_u3_n144 ) , .A1( u2_u5_u3_n153 ) , .A3( u2_u5_u3_n182 ) );
  OAI22_X1 u2_u5_u4_U10 (.B2( u2_u5_u4_n135 ) , .ZN( u2_u5_u4_n137 ) , .B1( u2_u5_u4_n153 ) , .A1( u2_u5_u4_n155 ) , .A2( u2_u5_u4_n171 ) );
  AND3_X1 u2_u5_u4_U11 (.A2( u2_u5_u4_n134 ) , .ZN( u2_u5_u4_n135 ) , .A3( u2_u5_u4_n145 ) , .A1( u2_u5_u4_n157 ) );
  NAND2_X1 u2_u5_u4_U12 (.ZN( u2_u5_u4_n132 ) , .A2( u2_u5_u4_n170 ) , .A1( u2_u5_u4_n173 ) );
  AOI21_X1 u2_u5_u4_U13 (.B2( u2_u5_u4_n160 ) , .B1( u2_u5_u4_n161 ) , .ZN( u2_u5_u4_n162 ) , .A( u2_u5_u4_n170 ) );
  AOI21_X1 u2_u5_u4_U14 (.ZN( u2_u5_u4_n107 ) , .B2( u2_u5_u4_n143 ) , .A( u2_u5_u4_n174 ) , .B1( u2_u5_u4_n184 ) );
  AOI21_X1 u2_u5_u4_U15 (.B2( u2_u5_u4_n158 ) , .B1( u2_u5_u4_n159 ) , .ZN( u2_u5_u4_n163 ) , .A( u2_u5_u4_n174 ) );
  AOI21_X1 u2_u5_u4_U16 (.A( u2_u5_u4_n153 ) , .B2( u2_u5_u4_n154 ) , .B1( u2_u5_u4_n155 ) , .ZN( u2_u5_u4_n165 ) );
  AOI21_X1 u2_u5_u4_U17 (.A( u2_u5_u4_n156 ) , .B2( u2_u5_u4_n157 ) , .ZN( u2_u5_u4_n164 ) , .B1( u2_u5_u4_n184 ) );
  INV_X1 u2_u5_u4_U18 (.A( u2_u5_u4_n138 ) , .ZN( u2_u5_u4_n170 ) );
  AND2_X1 u2_u5_u4_U19 (.A2( u2_u5_u4_n120 ) , .ZN( u2_u5_u4_n155 ) , .A1( u2_u5_u4_n160 ) );
  INV_X1 u2_u5_u4_U20 (.A( u2_u5_u4_n156 ) , .ZN( u2_u5_u4_n175 ) );
  NAND2_X1 u2_u5_u4_U21 (.A2( u2_u5_u4_n118 ) , .ZN( u2_u5_u4_n131 ) , .A1( u2_u5_u4_n147 ) );
  NAND2_X1 u2_u5_u4_U22 (.A1( u2_u5_u4_n119 ) , .A2( u2_u5_u4_n120 ) , .ZN( u2_u5_u4_n130 ) );
  NAND2_X1 u2_u5_u4_U23 (.ZN( u2_u5_u4_n117 ) , .A2( u2_u5_u4_n118 ) , .A1( u2_u5_u4_n148 ) );
  NAND2_X1 u2_u5_u4_U24 (.ZN( u2_u5_u4_n129 ) , .A1( u2_u5_u4_n134 ) , .A2( u2_u5_u4_n148 ) );
  AND3_X1 u2_u5_u4_U25 (.A1( u2_u5_u4_n119 ) , .A2( u2_u5_u4_n143 ) , .A3( u2_u5_u4_n154 ) , .ZN( u2_u5_u4_n161 ) );
  AND2_X1 u2_u5_u4_U26 (.A1( u2_u5_u4_n145 ) , .A2( u2_u5_u4_n147 ) , .ZN( u2_u5_u4_n159 ) );
  OR3_X1 u2_u5_u4_U27 (.A3( u2_u5_u4_n114 ) , .A2( u2_u5_u4_n115 ) , .A1( u2_u5_u4_n116 ) , .ZN( u2_u5_u4_n136 ) );
  AOI21_X1 u2_u5_u4_U28 (.A( u2_u5_u4_n113 ) , .ZN( u2_u5_u4_n116 ) , .B2( u2_u5_u4_n173 ) , .B1( u2_u5_u4_n174 ) );
  AOI21_X1 u2_u5_u4_U29 (.ZN( u2_u5_u4_n115 ) , .B2( u2_u5_u4_n145 ) , .B1( u2_u5_u4_n146 ) , .A( u2_u5_u4_n156 ) );
  NOR2_X1 u2_u5_u4_U3 (.ZN( u2_u5_u4_n121 ) , .A1( u2_u5_u4_n181 ) , .A2( u2_u5_u4_n182 ) );
  OAI22_X1 u2_u5_u4_U30 (.ZN( u2_u5_u4_n114 ) , .A2( u2_u5_u4_n121 ) , .B1( u2_u5_u4_n160 ) , .B2( u2_u5_u4_n170 ) , .A1( u2_u5_u4_n171 ) );
  INV_X1 u2_u5_u4_U31 (.A( u2_u5_u4_n158 ) , .ZN( u2_u5_u4_n182 ) );
  INV_X1 u2_u5_u4_U32 (.ZN( u2_u5_u4_n181 ) , .A( u2_u5_u4_n96 ) );
  INV_X1 u2_u5_u4_U33 (.A( u2_u5_u4_n144 ) , .ZN( u2_u5_u4_n179 ) );
  INV_X1 u2_u5_u4_U34 (.A( u2_u5_u4_n157 ) , .ZN( u2_u5_u4_n178 ) );
  NAND2_X1 u2_u5_u4_U35 (.A2( u2_u5_u4_n154 ) , .A1( u2_u5_u4_n96 ) , .ZN( u2_u5_u4_n97 ) );
  INV_X1 u2_u5_u4_U36 (.ZN( u2_u5_u4_n186 ) , .A( u2_u5_u4_n95 ) );
  OAI221_X1 u2_u5_u4_U37 (.C1( u2_u5_u4_n134 ) , .B1( u2_u5_u4_n158 ) , .B2( u2_u5_u4_n171 ) , .C2( u2_u5_u4_n173 ) , .A( u2_u5_u4_n94 ) , .ZN( u2_u5_u4_n95 ) );
  AOI222_X1 u2_u5_u4_U38 (.B2( u2_u5_u4_n132 ) , .A1( u2_u5_u4_n138 ) , .C2( u2_u5_u4_n175 ) , .A2( u2_u5_u4_n179 ) , .C1( u2_u5_u4_n181 ) , .B1( u2_u5_u4_n185 ) , .ZN( u2_u5_u4_n94 ) );
  INV_X1 u2_u5_u4_U39 (.A( u2_u5_u4_n113 ) , .ZN( u2_u5_u4_n185 ) );
  INV_X1 u2_u5_u4_U4 (.A( u2_u5_u4_n117 ) , .ZN( u2_u5_u4_n184 ) );
  INV_X1 u2_u5_u4_U40 (.A( u2_u5_u4_n143 ) , .ZN( u2_u5_u4_n183 ) );
  NOR2_X1 u2_u5_u4_U41 (.ZN( u2_u5_u4_n138 ) , .A1( u2_u5_u4_n168 ) , .A2( u2_u5_u4_n169 ) );
  NOR2_X1 u2_u5_u4_U42 (.A1( u2_u5_u4_n150 ) , .A2( u2_u5_u4_n152 ) , .ZN( u2_u5_u4_n153 ) );
  NOR2_X1 u2_u5_u4_U43 (.A2( u2_u5_u4_n128 ) , .A1( u2_u5_u4_n138 ) , .ZN( u2_u5_u4_n156 ) );
  AOI22_X1 u2_u5_u4_U44 (.B2( u2_u5_u4_n122 ) , .A1( u2_u5_u4_n123 ) , .ZN( u2_u5_u4_n124 ) , .B1( u2_u5_u4_n128 ) , .A2( u2_u5_u4_n172 ) );
  INV_X1 u2_u5_u4_U45 (.A( u2_u5_u4_n153 ) , .ZN( u2_u5_u4_n172 ) );
  NAND2_X1 u2_u5_u4_U46 (.A2( u2_u5_u4_n120 ) , .ZN( u2_u5_u4_n123 ) , .A1( u2_u5_u4_n161 ) );
  AOI22_X1 u2_u5_u4_U47 (.B2( u2_u5_u4_n132 ) , .A2( u2_u5_u4_n133 ) , .ZN( u2_u5_u4_n140 ) , .A1( u2_u5_u4_n150 ) , .B1( u2_u5_u4_n179 ) );
  NAND2_X1 u2_u5_u4_U48 (.ZN( u2_u5_u4_n133 ) , .A2( u2_u5_u4_n146 ) , .A1( u2_u5_u4_n154 ) );
  NAND2_X1 u2_u5_u4_U49 (.A1( u2_u5_u4_n103 ) , .ZN( u2_u5_u4_n154 ) , .A2( u2_u5_u4_n98 ) );
  NOR4_X1 u2_u5_u4_U5 (.A4( u2_u5_u4_n106 ) , .A3( u2_u5_u4_n107 ) , .A2( u2_u5_u4_n108 ) , .A1( u2_u5_u4_n109 ) , .ZN( u2_u5_u4_n110 ) );
  NAND2_X1 u2_u5_u4_U50 (.A1( u2_u5_u4_n101 ) , .ZN( u2_u5_u4_n158 ) , .A2( u2_u5_u4_n99 ) );
  AOI21_X1 u2_u5_u4_U51 (.ZN( u2_u5_u4_n127 ) , .A( u2_u5_u4_n136 ) , .B2( u2_u5_u4_n150 ) , .B1( u2_u5_u4_n180 ) );
  INV_X1 u2_u5_u4_U52 (.A( u2_u5_u4_n160 ) , .ZN( u2_u5_u4_n180 ) );
  NAND2_X1 u2_u5_u4_U53 (.A2( u2_u5_u4_n104 ) , .A1( u2_u5_u4_n105 ) , .ZN( u2_u5_u4_n146 ) );
  NAND2_X1 u2_u5_u4_U54 (.A2( u2_u5_u4_n101 ) , .A1( u2_u5_u4_n102 ) , .ZN( u2_u5_u4_n160 ) );
  NAND2_X1 u2_u5_u4_U55 (.ZN( u2_u5_u4_n134 ) , .A1( u2_u5_u4_n98 ) , .A2( u2_u5_u4_n99 ) );
  NAND2_X1 u2_u5_u4_U56 (.A1( u2_u5_u4_n103 ) , .A2( u2_u5_u4_n104 ) , .ZN( u2_u5_u4_n143 ) );
  NAND2_X1 u2_u5_u4_U57 (.A2( u2_u5_u4_n105 ) , .ZN( u2_u5_u4_n145 ) , .A1( u2_u5_u4_n98 ) );
  NAND2_X1 u2_u5_u4_U58 (.A1( u2_u5_u4_n100 ) , .A2( u2_u5_u4_n105 ) , .ZN( u2_u5_u4_n120 ) );
  NAND2_X1 u2_u5_u4_U59 (.A1( u2_u5_u4_n102 ) , .A2( u2_u5_u4_n104 ) , .ZN( u2_u5_u4_n148 ) );
  AOI21_X1 u2_u5_u4_U6 (.ZN( u2_u5_u4_n106 ) , .B2( u2_u5_u4_n146 ) , .B1( u2_u5_u4_n158 ) , .A( u2_u5_u4_n170 ) );
  NAND2_X1 u2_u5_u4_U60 (.A2( u2_u5_u4_n100 ) , .A1( u2_u5_u4_n103 ) , .ZN( u2_u5_u4_n157 ) );
  INV_X1 u2_u5_u4_U61 (.A( u2_u5_u4_n150 ) , .ZN( u2_u5_u4_n173 ) );
  INV_X1 u2_u5_u4_U62 (.A( u2_u5_u4_n152 ) , .ZN( u2_u5_u4_n171 ) );
  NAND2_X1 u2_u5_u4_U63 (.A1( u2_u5_u4_n100 ) , .ZN( u2_u5_u4_n118 ) , .A2( u2_u5_u4_n99 ) );
  NAND2_X1 u2_u5_u4_U64 (.A2( u2_u5_u4_n100 ) , .A1( u2_u5_u4_n102 ) , .ZN( u2_u5_u4_n144 ) );
  NAND2_X1 u2_u5_u4_U65 (.A2( u2_u5_u4_n101 ) , .A1( u2_u5_u4_n105 ) , .ZN( u2_u5_u4_n96 ) );
  INV_X1 u2_u5_u4_U66 (.A( u2_u5_u4_n128 ) , .ZN( u2_u5_u4_n174 ) );
  NAND2_X1 u2_u5_u4_U67 (.A2( u2_u5_u4_n102 ) , .ZN( u2_u5_u4_n119 ) , .A1( u2_u5_u4_n98 ) );
  NAND2_X1 u2_u5_u4_U68 (.A2( u2_u5_u4_n101 ) , .A1( u2_u5_u4_n103 ) , .ZN( u2_u5_u4_n147 ) );
  NAND2_X1 u2_u5_u4_U69 (.A2( u2_u5_u4_n104 ) , .ZN( u2_u5_u4_n113 ) , .A1( u2_u5_u4_n99 ) );
  AOI21_X1 u2_u5_u4_U7 (.ZN( u2_u5_u4_n108 ) , .B2( u2_u5_u4_n134 ) , .B1( u2_u5_u4_n155 ) , .A( u2_u5_u4_n156 ) );
  NOR2_X1 u2_u5_u4_U70 (.A2( u2_u5_X_28 ) , .ZN( u2_u5_u4_n150 ) , .A1( u2_u5_u4_n168 ) );
  NOR2_X1 u2_u5_u4_U71 (.A2( u2_u5_X_29 ) , .ZN( u2_u5_u4_n152 ) , .A1( u2_u5_u4_n169 ) );
  NOR2_X1 u2_u5_u4_U72 (.A2( u2_u5_X_30 ) , .ZN( u2_u5_u4_n105 ) , .A1( u2_u5_u4_n176 ) );
  NOR2_X1 u2_u5_u4_U73 (.A2( u2_u5_X_26 ) , .ZN( u2_u5_u4_n100 ) , .A1( u2_u5_u4_n177 ) );
  NOR2_X1 u2_u5_u4_U74 (.A2( u2_u5_X_28 ) , .A1( u2_u5_X_29 ) , .ZN( u2_u5_u4_n128 ) );
  NOR2_X1 u2_u5_u4_U75 (.A2( u2_u5_X_27 ) , .A1( u2_u5_X_30 ) , .ZN( u2_u5_u4_n102 ) );
  NOR2_X1 u2_u5_u4_U76 (.A2( u2_u5_X_25 ) , .A1( u2_u5_X_26 ) , .ZN( u2_u5_u4_n98 ) );
  AND2_X1 u2_u5_u4_U77 (.A2( u2_u5_X_25 ) , .A1( u2_u5_X_26 ) , .ZN( u2_u5_u4_n104 ) );
  AND2_X1 u2_u5_u4_U78 (.A1( u2_u5_X_30 ) , .A2( u2_u5_u4_n176 ) , .ZN( u2_u5_u4_n99 ) );
  AND2_X1 u2_u5_u4_U79 (.A1( u2_u5_X_26 ) , .ZN( u2_u5_u4_n101 ) , .A2( u2_u5_u4_n177 ) );
  AOI21_X1 u2_u5_u4_U8 (.ZN( u2_u5_u4_n109 ) , .A( u2_u5_u4_n153 ) , .B1( u2_u5_u4_n159 ) , .B2( u2_u5_u4_n184 ) );
  AND2_X1 u2_u5_u4_U80 (.A1( u2_u5_X_27 ) , .A2( u2_u5_X_30 ) , .ZN( u2_u5_u4_n103 ) );
  INV_X1 u2_u5_u4_U81 (.A( u2_u5_X_28 ) , .ZN( u2_u5_u4_n169 ) );
  INV_X1 u2_u5_u4_U82 (.A( u2_u5_X_29 ) , .ZN( u2_u5_u4_n168 ) );
  INV_X1 u2_u5_u4_U83 (.A( u2_u5_X_25 ) , .ZN( u2_u5_u4_n177 ) );
  INV_X1 u2_u5_u4_U84 (.A( u2_u5_X_27 ) , .ZN( u2_u5_u4_n176 ) );
  NAND4_X1 u2_u5_u4_U85 (.ZN( u2_out5_25 ) , .A4( u2_u5_u4_n139 ) , .A3( u2_u5_u4_n140 ) , .A2( u2_u5_u4_n141 ) , .A1( u2_u5_u4_n142 ) );
  OAI21_X1 u2_u5_u4_U86 (.A( u2_u5_u4_n128 ) , .B2( u2_u5_u4_n129 ) , .B1( u2_u5_u4_n130 ) , .ZN( u2_u5_u4_n142 ) );
  OAI21_X1 u2_u5_u4_U87 (.B2( u2_u5_u4_n131 ) , .ZN( u2_u5_u4_n141 ) , .A( u2_u5_u4_n175 ) , .B1( u2_u5_u4_n183 ) );
  NAND4_X1 u2_u5_u4_U88 (.ZN( u2_out5_14 ) , .A4( u2_u5_u4_n124 ) , .A3( u2_u5_u4_n125 ) , .A2( u2_u5_u4_n126 ) , .A1( u2_u5_u4_n127 ) );
  AOI22_X1 u2_u5_u4_U89 (.B2( u2_u5_u4_n117 ) , .ZN( u2_u5_u4_n126 ) , .A1( u2_u5_u4_n129 ) , .B1( u2_u5_u4_n152 ) , .A2( u2_u5_u4_n175 ) );
  AOI211_X1 u2_u5_u4_U9 (.B( u2_u5_u4_n136 ) , .A( u2_u5_u4_n137 ) , .C2( u2_u5_u4_n138 ) , .ZN( u2_u5_u4_n139 ) , .C1( u2_u5_u4_n182 ) );
  AOI22_X1 u2_u5_u4_U90 (.ZN( u2_u5_u4_n125 ) , .B2( u2_u5_u4_n131 ) , .A2( u2_u5_u4_n132 ) , .B1( u2_u5_u4_n138 ) , .A1( u2_u5_u4_n178 ) );
  NAND4_X1 u2_u5_u4_U91 (.ZN( u2_out5_8 ) , .A4( u2_u5_u4_n110 ) , .A3( u2_u5_u4_n111 ) , .A2( u2_u5_u4_n112 ) , .A1( u2_u5_u4_n186 ) );
  NAND2_X1 u2_u5_u4_U92 (.ZN( u2_u5_u4_n112 ) , .A2( u2_u5_u4_n130 ) , .A1( u2_u5_u4_n150 ) );
  AOI22_X1 u2_u5_u4_U93 (.ZN( u2_u5_u4_n111 ) , .B2( u2_u5_u4_n132 ) , .A1( u2_u5_u4_n152 ) , .B1( u2_u5_u4_n178 ) , .A2( u2_u5_u4_n97 ) );
  AOI22_X1 u2_u5_u4_U94 (.B2( u2_u5_u4_n149 ) , .B1( u2_u5_u4_n150 ) , .A2( u2_u5_u4_n151 ) , .A1( u2_u5_u4_n152 ) , .ZN( u2_u5_u4_n167 ) );
  NOR4_X1 u2_u5_u4_U95 (.A4( u2_u5_u4_n162 ) , .A3( u2_u5_u4_n163 ) , .A2( u2_u5_u4_n164 ) , .A1( u2_u5_u4_n165 ) , .ZN( u2_u5_u4_n166 ) );
  NAND3_X1 u2_u5_u4_U96 (.ZN( u2_out5_3 ) , .A3( u2_u5_u4_n166 ) , .A1( u2_u5_u4_n167 ) , .A2( u2_u5_u4_n186 ) );
  NAND3_X1 u2_u5_u4_U97 (.A3( u2_u5_u4_n146 ) , .A2( u2_u5_u4_n147 ) , .A1( u2_u5_u4_n148 ) , .ZN( u2_u5_u4_n149 ) );
  NAND3_X1 u2_u5_u4_U98 (.A3( u2_u5_u4_n143 ) , .A2( u2_u5_u4_n144 ) , .A1( u2_u5_u4_n145 ) , .ZN( u2_u5_u4_n151 ) );
  NAND3_X1 u2_u5_u4_U99 (.A3( u2_u5_u4_n121 ) , .ZN( u2_u5_u4_n122 ) , .A2( u2_u5_u4_n144 ) , .A1( u2_u5_u4_n154 ) );
  XOR2_X1 u2_u6_U1 (.B( u2_K7_9 ) , .A( u2_R5_6 ) , .Z( u2_u6_X_9 ) );
  XOR2_X1 u2_u6_U10 (.B( u2_K7_45 ) , .A( u2_R5_30 ) , .Z( u2_u6_X_45 ) );
  XOR2_X1 u2_u6_U11 (.B( u2_K7_44 ) , .A( u2_R5_29 ) , .Z( u2_u6_X_44 ) );
  XOR2_X1 u2_u6_U12 (.B( u2_K7_43 ) , .A( u2_R5_28 ) , .Z( u2_u6_X_43 ) );
  XOR2_X1 u2_u6_U13 (.B( u2_K7_42 ) , .A( u2_R5_29 ) , .Z( u2_u6_X_42 ) );
  XOR2_X1 u2_u6_U14 (.B( u2_K7_41 ) , .A( u2_R5_28 ) , .Z( u2_u6_X_41 ) );
  XOR2_X1 u2_u6_U15 (.B( u2_K7_40 ) , .A( u2_R5_27 ) , .Z( u2_u6_X_40 ) );
  XOR2_X1 u2_u6_U16 (.B( u2_K7_3 ) , .A( u2_R5_2 ) , .Z( u2_u6_X_3 ) );
  XOR2_X1 u2_u6_U17 (.B( u2_K7_39 ) , .A( u2_R5_26 ) , .Z( u2_u6_X_39 ) );
  XOR2_X1 u2_u6_U18 (.B( u2_K7_38 ) , .A( u2_R5_25 ) , .Z( u2_u6_X_38 ) );
  XOR2_X1 u2_u6_U19 (.B( u2_K7_37 ) , .A( u2_R5_24 ) , .Z( u2_u6_X_37 ) );
  XOR2_X1 u2_u6_U2 (.B( u2_K7_8 ) , .A( u2_R5_5 ) , .Z( u2_u6_X_8 ) );
  XOR2_X1 u2_u6_U26 (.B( u2_K7_30 ) , .A( u2_R5_21 ) , .Z( u2_u6_X_30 ) );
  XOR2_X1 u2_u6_U27 (.B( u2_K7_2 ) , .A( u2_R5_1 ) , .Z( u2_u6_X_2 ) );
  XOR2_X1 u2_u6_U28 (.B( u2_K7_29 ) , .A( u2_R5_20 ) , .Z( u2_u6_X_29 ) );
  XOR2_X1 u2_u6_U29 (.B( u2_K7_28 ) , .A( u2_R5_19 ) , .Z( u2_u6_X_28 ) );
  XOR2_X1 u2_u6_U3 (.B( u2_K7_7 ) , .A( u2_R5_4 ) , .Z( u2_u6_X_7 ) );
  XOR2_X1 u2_u6_U30 (.B( u2_K7_27 ) , .A( u2_R5_18 ) , .Z( u2_u6_X_27 ) );
  XOR2_X1 u2_u6_U31 (.B( u2_K7_26 ) , .A( u2_R5_17 ) , .Z( u2_u6_X_26 ) );
  XOR2_X1 u2_u6_U32 (.B( u2_K7_25 ) , .A( u2_R5_16 ) , .Z( u2_u6_X_25 ) );
  XOR2_X1 u2_u6_U33 (.B( u2_K7_24 ) , .A( u2_R5_17 ) , .Z( u2_u6_X_24 ) );
  XOR2_X1 u2_u6_U34 (.B( u2_K7_23 ) , .A( u2_R5_16 ) , .Z( u2_u6_X_23 ) );
  XOR2_X1 u2_u6_U35 (.B( u2_K7_22 ) , .A( u2_R5_15 ) , .Z( u2_u6_X_22 ) );
  XOR2_X1 u2_u6_U36 (.B( u2_K7_21 ) , .A( u2_R5_14 ) , .Z( u2_u6_X_21 ) );
  XOR2_X1 u2_u6_U37 (.B( u2_K7_20 ) , .A( u2_R5_13 ) , .Z( u2_u6_X_20 ) );
  XOR2_X1 u2_u6_U38 (.B( u2_K7_1 ) , .A( u2_R5_32 ) , .Z( u2_u6_X_1 ) );
  XOR2_X1 u2_u6_U39 (.B( u2_K7_19 ) , .A( u2_R5_12 ) , .Z( u2_u6_X_19 ) );
  XOR2_X1 u2_u6_U4 (.B( u2_K7_6 ) , .A( u2_R5_5 ) , .Z( u2_u6_X_6 ) );
  XOR2_X1 u2_u6_U40 (.B( u2_K7_18 ) , .A( u2_R5_13 ) , .Z( u2_u6_X_18 ) );
  XOR2_X1 u2_u6_U41 (.B( u2_K7_17 ) , .A( u2_R5_12 ) , .Z( u2_u6_X_17 ) );
  XOR2_X1 u2_u6_U42 (.B( u2_K7_16 ) , .A( u2_R5_11 ) , .Z( u2_u6_X_16 ) );
  XOR2_X1 u2_u6_U43 (.B( u2_K7_15 ) , .A( u2_R5_10 ) , .Z( u2_u6_X_15 ) );
  XOR2_X1 u2_u6_U44 (.B( u2_K7_14 ) , .A( u2_R5_9 ) , .Z( u2_u6_X_14 ) );
  XOR2_X1 u2_u6_U45 (.B( u2_K7_13 ) , .A( u2_R5_8 ) , .Z( u2_u6_X_13 ) );
  XOR2_X1 u2_u6_U46 (.B( u2_K7_12 ) , .A( u2_R5_9 ) , .Z( u2_u6_X_12 ) );
  XOR2_X1 u2_u6_U47 (.B( u2_K7_11 ) , .A( u2_R5_8 ) , .Z( u2_u6_X_11 ) );
  XOR2_X1 u2_u6_U48 (.B( u2_K7_10 ) , .A( u2_R5_7 ) , .Z( u2_u6_X_10 ) );
  XOR2_X1 u2_u6_U5 (.B( u2_K7_5 ) , .A( u2_R5_4 ) , .Z( u2_u6_X_5 ) );
  XOR2_X1 u2_u6_U6 (.B( u2_K7_4 ) , .A( u2_R5_3 ) , .Z( u2_u6_X_4 ) );
  XOR2_X1 u2_u6_U7 (.B( u2_K7_48 ) , .A( u2_R5_1 ) , .Z( u2_u6_X_48 ) );
  XOR2_X1 u2_u6_U8 (.B( u2_K7_47 ) , .A( u2_R5_32 ) , .Z( u2_u6_X_47 ) );
  XOR2_X1 u2_u6_U9 (.B( u2_K7_46 ) , .A( u2_R5_31 ) , .Z( u2_u6_X_46 ) );
  AND3_X1 u2_u6_u0_U10 (.A2( u2_u6_u0_n112 ) , .ZN( u2_u6_u0_n127 ) , .A3( u2_u6_u0_n130 ) , .A1( u2_u6_u0_n148 ) );
  NAND2_X1 u2_u6_u0_U11 (.ZN( u2_u6_u0_n113 ) , .A1( u2_u6_u0_n139 ) , .A2( u2_u6_u0_n149 ) );
  AND2_X1 u2_u6_u0_U12 (.ZN( u2_u6_u0_n107 ) , .A1( u2_u6_u0_n130 ) , .A2( u2_u6_u0_n140 ) );
  AND2_X1 u2_u6_u0_U13 (.A2( u2_u6_u0_n129 ) , .A1( u2_u6_u0_n130 ) , .ZN( u2_u6_u0_n151 ) );
  AND2_X1 u2_u6_u0_U14 (.A1( u2_u6_u0_n108 ) , .A2( u2_u6_u0_n125 ) , .ZN( u2_u6_u0_n145 ) );
  INV_X1 u2_u6_u0_U15 (.A( u2_u6_u0_n143 ) , .ZN( u2_u6_u0_n173 ) );
  NOR2_X1 u2_u6_u0_U16 (.A2( u2_u6_u0_n136 ) , .ZN( u2_u6_u0_n147 ) , .A1( u2_u6_u0_n160 ) );
  NOR2_X1 u2_u6_u0_U17 (.A1( u2_u6_u0_n163 ) , .A2( u2_u6_u0_n164 ) , .ZN( u2_u6_u0_n95 ) );
  AOI21_X1 u2_u6_u0_U18 (.B1( u2_u6_u0_n103 ) , .ZN( u2_u6_u0_n132 ) , .A( u2_u6_u0_n165 ) , .B2( u2_u6_u0_n93 ) );
  INV_X1 u2_u6_u0_U19 (.A( u2_u6_u0_n142 ) , .ZN( u2_u6_u0_n165 ) );
  OAI22_X1 u2_u6_u0_U20 (.B1( u2_u6_u0_n125 ) , .ZN( u2_u6_u0_n126 ) , .A1( u2_u6_u0_n138 ) , .A2( u2_u6_u0_n146 ) , .B2( u2_u6_u0_n147 ) );
  OAI22_X1 u2_u6_u0_U21 (.B1( u2_u6_u0_n131 ) , .A1( u2_u6_u0_n144 ) , .B2( u2_u6_u0_n147 ) , .A2( u2_u6_u0_n90 ) , .ZN( u2_u6_u0_n91 ) );
  AND3_X1 u2_u6_u0_U22 (.A3( u2_u6_u0_n121 ) , .A2( u2_u6_u0_n125 ) , .A1( u2_u6_u0_n148 ) , .ZN( u2_u6_u0_n90 ) );
  NAND2_X1 u2_u6_u0_U23 (.A1( u2_u6_u0_n100 ) , .A2( u2_u6_u0_n103 ) , .ZN( u2_u6_u0_n125 ) );
  INV_X1 u2_u6_u0_U24 (.A( u2_u6_u0_n136 ) , .ZN( u2_u6_u0_n161 ) );
  AOI22_X1 u2_u6_u0_U25 (.B2( u2_u6_u0_n109 ) , .A2( u2_u6_u0_n110 ) , .ZN( u2_u6_u0_n111 ) , .B1( u2_u6_u0_n118 ) , .A1( u2_u6_u0_n160 ) );
  NAND2_X1 u2_u6_u0_U26 (.A1( u2_u6_u0_n100 ) , .ZN( u2_u6_u0_n129 ) , .A2( u2_u6_u0_n95 ) );
  INV_X1 u2_u6_u0_U27 (.A( u2_u6_u0_n118 ) , .ZN( u2_u6_u0_n158 ) );
  AOI21_X1 u2_u6_u0_U28 (.ZN( u2_u6_u0_n104 ) , .B1( u2_u6_u0_n107 ) , .B2( u2_u6_u0_n141 ) , .A( u2_u6_u0_n144 ) );
  AOI21_X1 u2_u6_u0_U29 (.B1( u2_u6_u0_n127 ) , .B2( u2_u6_u0_n129 ) , .A( u2_u6_u0_n138 ) , .ZN( u2_u6_u0_n96 ) );
  INV_X1 u2_u6_u0_U3 (.A( u2_u6_u0_n113 ) , .ZN( u2_u6_u0_n166 ) );
  AOI21_X1 u2_u6_u0_U30 (.ZN( u2_u6_u0_n116 ) , .B2( u2_u6_u0_n142 ) , .A( u2_u6_u0_n144 ) , .B1( u2_u6_u0_n166 ) );
  NOR2_X1 u2_u6_u0_U31 (.A1( u2_u6_u0_n120 ) , .ZN( u2_u6_u0_n143 ) , .A2( u2_u6_u0_n167 ) );
  OAI221_X1 u2_u6_u0_U32 (.C1( u2_u6_u0_n112 ) , .ZN( u2_u6_u0_n120 ) , .B1( u2_u6_u0_n138 ) , .B2( u2_u6_u0_n141 ) , .C2( u2_u6_u0_n147 ) , .A( u2_u6_u0_n172 ) );
  AOI211_X1 u2_u6_u0_U33 (.B( u2_u6_u0_n115 ) , .A( u2_u6_u0_n116 ) , .C2( u2_u6_u0_n117 ) , .C1( u2_u6_u0_n118 ) , .ZN( u2_u6_u0_n119 ) );
  NAND2_X1 u2_u6_u0_U34 (.A2( u2_u6_u0_n100 ) , .A1( u2_u6_u0_n101 ) , .ZN( u2_u6_u0_n139 ) );
  NAND2_X1 u2_u6_u0_U35 (.A2( u2_u6_u0_n100 ) , .ZN( u2_u6_u0_n131 ) , .A1( u2_u6_u0_n92 ) );
  NAND2_X1 u2_u6_u0_U36 (.A1( u2_u6_u0_n101 ) , .A2( u2_u6_u0_n102 ) , .ZN( u2_u6_u0_n150 ) );
  INV_X1 u2_u6_u0_U37 (.A( u2_u6_u0_n138 ) , .ZN( u2_u6_u0_n160 ) );
  NAND2_X1 u2_u6_u0_U38 (.A1( u2_u6_u0_n102 ) , .ZN( u2_u6_u0_n128 ) , .A2( u2_u6_u0_n95 ) );
  NAND2_X1 u2_u6_u0_U39 (.ZN( u2_u6_u0_n148 ) , .A1( u2_u6_u0_n93 ) , .A2( u2_u6_u0_n95 ) );
  AOI21_X1 u2_u6_u0_U4 (.B1( u2_u6_u0_n114 ) , .ZN( u2_u6_u0_n115 ) , .B2( u2_u6_u0_n129 ) , .A( u2_u6_u0_n161 ) );
  NAND2_X1 u2_u6_u0_U40 (.A2( u2_u6_u0_n102 ) , .A1( u2_u6_u0_n103 ) , .ZN( u2_u6_u0_n149 ) );
  NAND2_X1 u2_u6_u0_U41 (.A2( u2_u6_u0_n102 ) , .ZN( u2_u6_u0_n114 ) , .A1( u2_u6_u0_n92 ) );
  NAND2_X1 u2_u6_u0_U42 (.A2( u2_u6_u0_n101 ) , .ZN( u2_u6_u0_n121 ) , .A1( u2_u6_u0_n93 ) );
  NAND2_X1 u2_u6_u0_U43 (.ZN( u2_u6_u0_n112 ) , .A2( u2_u6_u0_n92 ) , .A1( u2_u6_u0_n93 ) );
  INV_X1 u2_u6_u0_U44 (.ZN( u2_u6_u0_n172 ) , .A( u2_u6_u0_n88 ) );
  OAI222_X1 u2_u6_u0_U45 (.C1( u2_u6_u0_n108 ) , .A1( u2_u6_u0_n125 ) , .B2( u2_u6_u0_n128 ) , .B1( u2_u6_u0_n144 ) , .A2( u2_u6_u0_n158 ) , .C2( u2_u6_u0_n161 ) , .ZN( u2_u6_u0_n88 ) );
  OR3_X1 u2_u6_u0_U46 (.A3( u2_u6_u0_n152 ) , .A2( u2_u6_u0_n153 ) , .A1( u2_u6_u0_n154 ) , .ZN( u2_u6_u0_n155 ) );
  AOI21_X1 u2_u6_u0_U47 (.A( u2_u6_u0_n144 ) , .B2( u2_u6_u0_n145 ) , .B1( u2_u6_u0_n146 ) , .ZN( u2_u6_u0_n154 ) );
  AOI21_X1 u2_u6_u0_U48 (.B2( u2_u6_u0_n150 ) , .B1( u2_u6_u0_n151 ) , .ZN( u2_u6_u0_n152 ) , .A( u2_u6_u0_n158 ) );
  AOI21_X1 u2_u6_u0_U49 (.A( u2_u6_u0_n147 ) , .B2( u2_u6_u0_n148 ) , .B1( u2_u6_u0_n149 ) , .ZN( u2_u6_u0_n153 ) );
  AOI21_X1 u2_u6_u0_U5 (.B2( u2_u6_u0_n131 ) , .ZN( u2_u6_u0_n134 ) , .B1( u2_u6_u0_n151 ) , .A( u2_u6_u0_n158 ) );
  INV_X1 u2_u6_u0_U50 (.ZN( u2_u6_u0_n171 ) , .A( u2_u6_u0_n99 ) );
  OAI211_X1 u2_u6_u0_U51 (.C2( u2_u6_u0_n140 ) , .C1( u2_u6_u0_n161 ) , .A( u2_u6_u0_n169 ) , .B( u2_u6_u0_n98 ) , .ZN( u2_u6_u0_n99 ) );
  INV_X1 u2_u6_u0_U52 (.ZN( u2_u6_u0_n169 ) , .A( u2_u6_u0_n91 ) );
  AOI211_X1 u2_u6_u0_U53 (.C1( u2_u6_u0_n118 ) , .A( u2_u6_u0_n123 ) , .B( u2_u6_u0_n96 ) , .C2( u2_u6_u0_n97 ) , .ZN( u2_u6_u0_n98 ) );
  NOR2_X1 u2_u6_u0_U54 (.A2( u2_u6_X_4 ) , .A1( u2_u6_X_5 ) , .ZN( u2_u6_u0_n118 ) );
  NOR2_X1 u2_u6_u0_U55 (.A2( u2_u6_X_2 ) , .ZN( u2_u6_u0_n103 ) , .A1( u2_u6_u0_n164 ) );
  NOR2_X1 u2_u6_u0_U56 (.A2( u2_u6_X_1 ) , .A1( u2_u6_X_2 ) , .ZN( u2_u6_u0_n92 ) );
  NOR2_X1 u2_u6_u0_U57 (.A2( u2_u6_X_1 ) , .ZN( u2_u6_u0_n101 ) , .A1( u2_u6_u0_n163 ) );
  NAND2_X1 u2_u6_u0_U58 (.A2( u2_u6_X_4 ) , .A1( u2_u6_X_5 ) , .ZN( u2_u6_u0_n144 ) );
  NOR2_X1 u2_u6_u0_U59 (.A2( u2_u6_X_5 ) , .ZN( u2_u6_u0_n136 ) , .A1( u2_u6_u0_n159 ) );
  NOR2_X1 u2_u6_u0_U6 (.A1( u2_u6_u0_n108 ) , .ZN( u2_u6_u0_n123 ) , .A2( u2_u6_u0_n158 ) );
  NAND2_X1 u2_u6_u0_U60 (.A1( u2_u6_X_5 ) , .ZN( u2_u6_u0_n138 ) , .A2( u2_u6_u0_n159 ) );
  INV_X1 u2_u6_u0_U61 (.A( u2_u6_X_4 ) , .ZN( u2_u6_u0_n159 ) );
  INV_X1 u2_u6_u0_U62 (.A( u2_u6_X_1 ) , .ZN( u2_u6_u0_n164 ) );
  INV_X1 u2_u6_u0_U63 (.A( u2_u6_X_2 ) , .ZN( u2_u6_u0_n163 ) );
  INV_X1 u2_u6_u0_U64 (.A( u2_u6_X_3 ) , .ZN( u2_u6_u0_n162 ) );
  INV_X1 u2_u6_u0_U65 (.A( u2_u6_u0_n126 ) , .ZN( u2_u6_u0_n168 ) );
  AOI211_X1 u2_u6_u0_U66 (.B( u2_u6_u0_n133 ) , .A( u2_u6_u0_n134 ) , .C2( u2_u6_u0_n135 ) , .C1( u2_u6_u0_n136 ) , .ZN( u2_u6_u0_n137 ) );
  OR4_X1 u2_u6_u0_U67 (.ZN( u2_out6_17 ) , .A4( u2_u6_u0_n122 ) , .A2( u2_u6_u0_n123 ) , .A1( u2_u6_u0_n124 ) , .A3( u2_u6_u0_n170 ) );
  AOI21_X1 u2_u6_u0_U68 (.B2( u2_u6_u0_n107 ) , .ZN( u2_u6_u0_n124 ) , .B1( u2_u6_u0_n128 ) , .A( u2_u6_u0_n161 ) );
  INV_X1 u2_u6_u0_U69 (.A( u2_u6_u0_n111 ) , .ZN( u2_u6_u0_n170 ) );
  OAI21_X1 u2_u6_u0_U7 (.B1( u2_u6_u0_n150 ) , .B2( u2_u6_u0_n158 ) , .A( u2_u6_u0_n172 ) , .ZN( u2_u6_u0_n89 ) );
  OR4_X1 u2_u6_u0_U70 (.ZN( u2_out6_31 ) , .A4( u2_u6_u0_n155 ) , .A2( u2_u6_u0_n156 ) , .A1( u2_u6_u0_n157 ) , .A3( u2_u6_u0_n173 ) );
  AOI21_X1 u2_u6_u0_U71 (.A( u2_u6_u0_n138 ) , .B2( u2_u6_u0_n139 ) , .B1( u2_u6_u0_n140 ) , .ZN( u2_u6_u0_n157 ) );
  AOI21_X1 u2_u6_u0_U72 (.B2( u2_u6_u0_n141 ) , .B1( u2_u6_u0_n142 ) , .ZN( u2_u6_u0_n156 ) , .A( u2_u6_u0_n161 ) );
  INV_X1 u2_u6_u0_U73 (.ZN( u2_u6_u0_n174 ) , .A( u2_u6_u0_n89 ) );
  AOI211_X1 u2_u6_u0_U74 (.B( u2_u6_u0_n104 ) , .A( u2_u6_u0_n105 ) , .ZN( u2_u6_u0_n106 ) , .C2( u2_u6_u0_n113 ) , .C1( u2_u6_u0_n160 ) );
  AND2_X1 u2_u6_u0_U75 (.A1( u2_u6_X_6 ) , .A2( u2_u6_u0_n162 ) , .ZN( u2_u6_u0_n93 ) );
  NOR2_X1 u2_u6_u0_U76 (.A2( u2_u6_X_3 ) , .A1( u2_u6_X_6 ) , .ZN( u2_u6_u0_n94 ) );
  NOR2_X1 u2_u6_u0_U77 (.A2( u2_u6_X_6 ) , .ZN( u2_u6_u0_n100 ) , .A1( u2_u6_u0_n162 ) );
  AND2_X1 u2_u6_u0_U78 (.A2( u2_u6_X_3 ) , .A1( u2_u6_X_6 ) , .ZN( u2_u6_u0_n102 ) );
  OAI221_X1 u2_u6_u0_U79 (.C1( u2_u6_u0_n121 ) , .ZN( u2_u6_u0_n122 ) , .B2( u2_u6_u0_n127 ) , .A( u2_u6_u0_n143 ) , .B1( u2_u6_u0_n144 ) , .C2( u2_u6_u0_n147 ) );
  AND2_X1 u2_u6_u0_U8 (.A1( u2_u6_u0_n114 ) , .A2( u2_u6_u0_n121 ) , .ZN( u2_u6_u0_n146 ) );
  AOI21_X1 u2_u6_u0_U80 (.B1( u2_u6_u0_n132 ) , .ZN( u2_u6_u0_n133 ) , .A( u2_u6_u0_n144 ) , .B2( u2_u6_u0_n166 ) );
  OAI22_X1 u2_u6_u0_U81 (.ZN( u2_u6_u0_n105 ) , .A2( u2_u6_u0_n132 ) , .B1( u2_u6_u0_n146 ) , .A1( u2_u6_u0_n147 ) , .B2( u2_u6_u0_n161 ) );
  NAND2_X1 u2_u6_u0_U82 (.ZN( u2_u6_u0_n110 ) , .A2( u2_u6_u0_n132 ) , .A1( u2_u6_u0_n145 ) );
  INV_X1 u2_u6_u0_U83 (.A( u2_u6_u0_n119 ) , .ZN( u2_u6_u0_n167 ) );
  NAND2_X1 u2_u6_u0_U84 (.A2( u2_u6_u0_n103 ) , .ZN( u2_u6_u0_n140 ) , .A1( u2_u6_u0_n94 ) );
  NAND2_X1 u2_u6_u0_U85 (.A1( u2_u6_u0_n101 ) , .ZN( u2_u6_u0_n130 ) , .A2( u2_u6_u0_n94 ) );
  NAND2_X1 u2_u6_u0_U86 (.ZN( u2_u6_u0_n108 ) , .A1( u2_u6_u0_n92 ) , .A2( u2_u6_u0_n94 ) );
  NAND2_X1 u2_u6_u0_U87 (.ZN( u2_u6_u0_n142 ) , .A1( u2_u6_u0_n94 ) , .A2( u2_u6_u0_n95 ) );
  NAND3_X1 u2_u6_u0_U88 (.ZN( u2_out6_23 ) , .A3( u2_u6_u0_n137 ) , .A1( u2_u6_u0_n168 ) , .A2( u2_u6_u0_n171 ) );
  NAND3_X1 u2_u6_u0_U89 (.A3( u2_u6_u0_n127 ) , .A2( u2_u6_u0_n128 ) , .ZN( u2_u6_u0_n135 ) , .A1( u2_u6_u0_n150 ) );
  AND2_X1 u2_u6_u0_U9 (.A1( u2_u6_u0_n131 ) , .ZN( u2_u6_u0_n141 ) , .A2( u2_u6_u0_n150 ) );
  NAND3_X1 u2_u6_u0_U90 (.ZN( u2_u6_u0_n117 ) , .A3( u2_u6_u0_n132 ) , .A2( u2_u6_u0_n139 ) , .A1( u2_u6_u0_n148 ) );
  NAND3_X1 u2_u6_u0_U91 (.ZN( u2_u6_u0_n109 ) , .A2( u2_u6_u0_n114 ) , .A3( u2_u6_u0_n140 ) , .A1( u2_u6_u0_n149 ) );
  NAND3_X1 u2_u6_u0_U92 (.ZN( u2_out6_9 ) , .A3( u2_u6_u0_n106 ) , .A2( u2_u6_u0_n171 ) , .A1( u2_u6_u0_n174 ) );
  NAND3_X1 u2_u6_u0_U93 (.A2( u2_u6_u0_n128 ) , .A1( u2_u6_u0_n132 ) , .A3( u2_u6_u0_n146 ) , .ZN( u2_u6_u0_n97 ) );
  AOI21_X1 u2_u6_u1_U10 (.B2( u2_u6_u1_n155 ) , .B1( u2_u6_u1_n156 ) , .ZN( u2_u6_u1_n157 ) , .A( u2_u6_u1_n174 ) );
  NAND3_X1 u2_u6_u1_U100 (.ZN( u2_u6_u1_n113 ) , .A1( u2_u6_u1_n120 ) , .A3( u2_u6_u1_n133 ) , .A2( u2_u6_u1_n155 ) );
  NAND2_X1 u2_u6_u1_U11 (.ZN( u2_u6_u1_n140 ) , .A2( u2_u6_u1_n150 ) , .A1( u2_u6_u1_n155 ) );
  NAND2_X1 u2_u6_u1_U12 (.A1( u2_u6_u1_n131 ) , .ZN( u2_u6_u1_n147 ) , .A2( u2_u6_u1_n153 ) );
  INV_X1 u2_u6_u1_U13 (.A( u2_u6_u1_n139 ) , .ZN( u2_u6_u1_n174 ) );
  OR4_X1 u2_u6_u1_U14 (.A4( u2_u6_u1_n106 ) , .A3( u2_u6_u1_n107 ) , .ZN( u2_u6_u1_n108 ) , .A1( u2_u6_u1_n117 ) , .A2( u2_u6_u1_n184 ) );
  AOI21_X1 u2_u6_u1_U15 (.ZN( u2_u6_u1_n106 ) , .A( u2_u6_u1_n112 ) , .B1( u2_u6_u1_n154 ) , .B2( u2_u6_u1_n156 ) );
  AOI21_X1 u2_u6_u1_U16 (.ZN( u2_u6_u1_n107 ) , .B1( u2_u6_u1_n134 ) , .B2( u2_u6_u1_n149 ) , .A( u2_u6_u1_n174 ) );
  INV_X1 u2_u6_u1_U17 (.A( u2_u6_u1_n101 ) , .ZN( u2_u6_u1_n184 ) );
  INV_X1 u2_u6_u1_U18 (.A( u2_u6_u1_n112 ) , .ZN( u2_u6_u1_n171 ) );
  NAND2_X1 u2_u6_u1_U19 (.ZN( u2_u6_u1_n141 ) , .A1( u2_u6_u1_n153 ) , .A2( u2_u6_u1_n156 ) );
  AND2_X1 u2_u6_u1_U20 (.A1( u2_u6_u1_n123 ) , .ZN( u2_u6_u1_n134 ) , .A2( u2_u6_u1_n161 ) );
  NAND2_X1 u2_u6_u1_U21 (.A2( u2_u6_u1_n115 ) , .A1( u2_u6_u1_n116 ) , .ZN( u2_u6_u1_n148 ) );
  NAND2_X1 u2_u6_u1_U22 (.A2( u2_u6_u1_n133 ) , .A1( u2_u6_u1_n135 ) , .ZN( u2_u6_u1_n159 ) );
  NAND2_X1 u2_u6_u1_U23 (.A2( u2_u6_u1_n115 ) , .A1( u2_u6_u1_n120 ) , .ZN( u2_u6_u1_n132 ) );
  INV_X1 u2_u6_u1_U24 (.A( u2_u6_u1_n154 ) , .ZN( u2_u6_u1_n178 ) );
  AOI22_X1 u2_u6_u1_U25 (.B2( u2_u6_u1_n113 ) , .A2( u2_u6_u1_n114 ) , .ZN( u2_u6_u1_n125 ) , .A1( u2_u6_u1_n171 ) , .B1( u2_u6_u1_n173 ) );
  NAND2_X1 u2_u6_u1_U26 (.ZN( u2_u6_u1_n114 ) , .A1( u2_u6_u1_n134 ) , .A2( u2_u6_u1_n156 ) );
  INV_X1 u2_u6_u1_U27 (.A( u2_u6_u1_n151 ) , .ZN( u2_u6_u1_n183 ) );
  AND2_X1 u2_u6_u1_U28 (.A1( u2_u6_u1_n129 ) , .A2( u2_u6_u1_n133 ) , .ZN( u2_u6_u1_n149 ) );
  INV_X1 u2_u6_u1_U29 (.A( u2_u6_u1_n131 ) , .ZN( u2_u6_u1_n180 ) );
  INV_X1 u2_u6_u1_U3 (.A( u2_u6_u1_n159 ) , .ZN( u2_u6_u1_n182 ) );
  AOI221_X1 u2_u6_u1_U30 (.B1( u2_u6_u1_n140 ) , .ZN( u2_u6_u1_n167 ) , .B2( u2_u6_u1_n172 ) , .C2( u2_u6_u1_n175 ) , .C1( u2_u6_u1_n178 ) , .A( u2_u6_u1_n188 ) );
  INV_X1 u2_u6_u1_U31 (.ZN( u2_u6_u1_n188 ) , .A( u2_u6_u1_n97 ) );
  AOI211_X1 u2_u6_u1_U32 (.A( u2_u6_u1_n118 ) , .C1( u2_u6_u1_n132 ) , .C2( u2_u6_u1_n139 ) , .B( u2_u6_u1_n96 ) , .ZN( u2_u6_u1_n97 ) );
  AOI21_X1 u2_u6_u1_U33 (.B2( u2_u6_u1_n121 ) , .B1( u2_u6_u1_n135 ) , .A( u2_u6_u1_n152 ) , .ZN( u2_u6_u1_n96 ) );
  OAI221_X1 u2_u6_u1_U34 (.A( u2_u6_u1_n119 ) , .C2( u2_u6_u1_n129 ) , .ZN( u2_u6_u1_n138 ) , .B2( u2_u6_u1_n152 ) , .C1( u2_u6_u1_n174 ) , .B1( u2_u6_u1_n187 ) );
  INV_X1 u2_u6_u1_U35 (.A( u2_u6_u1_n148 ) , .ZN( u2_u6_u1_n187 ) );
  AOI211_X1 u2_u6_u1_U36 (.B( u2_u6_u1_n117 ) , .A( u2_u6_u1_n118 ) , .ZN( u2_u6_u1_n119 ) , .C2( u2_u6_u1_n146 ) , .C1( u2_u6_u1_n159 ) );
  NOR2_X1 u2_u6_u1_U37 (.A1( u2_u6_u1_n168 ) , .A2( u2_u6_u1_n176 ) , .ZN( u2_u6_u1_n98 ) );
  AOI211_X1 u2_u6_u1_U38 (.B( u2_u6_u1_n162 ) , .A( u2_u6_u1_n163 ) , .C2( u2_u6_u1_n164 ) , .ZN( u2_u6_u1_n165 ) , .C1( u2_u6_u1_n171 ) );
  AOI21_X1 u2_u6_u1_U39 (.A( u2_u6_u1_n160 ) , .B2( u2_u6_u1_n161 ) , .ZN( u2_u6_u1_n162 ) , .B1( u2_u6_u1_n182 ) );
  AOI221_X1 u2_u6_u1_U4 (.A( u2_u6_u1_n138 ) , .C2( u2_u6_u1_n139 ) , .C1( u2_u6_u1_n140 ) , .B2( u2_u6_u1_n141 ) , .ZN( u2_u6_u1_n142 ) , .B1( u2_u6_u1_n175 ) );
  OR2_X1 u2_u6_u1_U40 (.A2( u2_u6_u1_n157 ) , .A1( u2_u6_u1_n158 ) , .ZN( u2_u6_u1_n163 ) );
  NAND2_X1 u2_u6_u1_U41 (.A1( u2_u6_u1_n128 ) , .ZN( u2_u6_u1_n146 ) , .A2( u2_u6_u1_n160 ) );
  NAND2_X1 u2_u6_u1_U42 (.A2( u2_u6_u1_n112 ) , .ZN( u2_u6_u1_n139 ) , .A1( u2_u6_u1_n152 ) );
  NAND2_X1 u2_u6_u1_U43 (.A1( u2_u6_u1_n105 ) , .ZN( u2_u6_u1_n156 ) , .A2( u2_u6_u1_n99 ) );
  NOR2_X1 u2_u6_u1_U44 (.ZN( u2_u6_u1_n117 ) , .A1( u2_u6_u1_n121 ) , .A2( u2_u6_u1_n160 ) );
  OAI21_X1 u2_u6_u1_U45 (.B2( u2_u6_u1_n123 ) , .ZN( u2_u6_u1_n145 ) , .B1( u2_u6_u1_n160 ) , .A( u2_u6_u1_n185 ) );
  INV_X1 u2_u6_u1_U46 (.A( u2_u6_u1_n122 ) , .ZN( u2_u6_u1_n185 ) );
  AOI21_X1 u2_u6_u1_U47 (.B2( u2_u6_u1_n120 ) , .B1( u2_u6_u1_n121 ) , .ZN( u2_u6_u1_n122 ) , .A( u2_u6_u1_n128 ) );
  AOI21_X1 u2_u6_u1_U48 (.A( u2_u6_u1_n128 ) , .B2( u2_u6_u1_n129 ) , .ZN( u2_u6_u1_n130 ) , .B1( u2_u6_u1_n150 ) );
  NAND2_X1 u2_u6_u1_U49 (.ZN( u2_u6_u1_n112 ) , .A1( u2_u6_u1_n169 ) , .A2( u2_u6_u1_n170 ) );
  AOI211_X1 u2_u6_u1_U5 (.ZN( u2_u6_u1_n124 ) , .A( u2_u6_u1_n138 ) , .C2( u2_u6_u1_n139 ) , .B( u2_u6_u1_n145 ) , .C1( u2_u6_u1_n147 ) );
  NAND2_X1 u2_u6_u1_U50 (.ZN( u2_u6_u1_n129 ) , .A2( u2_u6_u1_n95 ) , .A1( u2_u6_u1_n98 ) );
  NAND2_X1 u2_u6_u1_U51 (.A1( u2_u6_u1_n102 ) , .ZN( u2_u6_u1_n154 ) , .A2( u2_u6_u1_n99 ) );
  NAND2_X1 u2_u6_u1_U52 (.A2( u2_u6_u1_n100 ) , .ZN( u2_u6_u1_n135 ) , .A1( u2_u6_u1_n99 ) );
  AOI21_X1 u2_u6_u1_U53 (.A( u2_u6_u1_n152 ) , .B2( u2_u6_u1_n153 ) , .B1( u2_u6_u1_n154 ) , .ZN( u2_u6_u1_n158 ) );
  INV_X1 u2_u6_u1_U54 (.A( u2_u6_u1_n160 ) , .ZN( u2_u6_u1_n175 ) );
  NAND2_X1 u2_u6_u1_U55 (.A1( u2_u6_u1_n100 ) , .ZN( u2_u6_u1_n116 ) , .A2( u2_u6_u1_n95 ) );
  NAND2_X1 u2_u6_u1_U56 (.A1( u2_u6_u1_n102 ) , .ZN( u2_u6_u1_n131 ) , .A2( u2_u6_u1_n95 ) );
  NAND2_X1 u2_u6_u1_U57 (.A2( u2_u6_u1_n104 ) , .ZN( u2_u6_u1_n121 ) , .A1( u2_u6_u1_n98 ) );
  NAND2_X1 u2_u6_u1_U58 (.A1( u2_u6_u1_n103 ) , .ZN( u2_u6_u1_n153 ) , .A2( u2_u6_u1_n98 ) );
  NAND2_X1 u2_u6_u1_U59 (.A2( u2_u6_u1_n104 ) , .A1( u2_u6_u1_n105 ) , .ZN( u2_u6_u1_n133 ) );
  AOI22_X1 u2_u6_u1_U6 (.B2( u2_u6_u1_n136 ) , .A2( u2_u6_u1_n137 ) , .ZN( u2_u6_u1_n143 ) , .A1( u2_u6_u1_n171 ) , .B1( u2_u6_u1_n173 ) );
  NAND2_X1 u2_u6_u1_U60 (.ZN( u2_u6_u1_n150 ) , .A2( u2_u6_u1_n98 ) , .A1( u2_u6_u1_n99 ) );
  NAND2_X1 u2_u6_u1_U61 (.A1( u2_u6_u1_n105 ) , .ZN( u2_u6_u1_n155 ) , .A2( u2_u6_u1_n95 ) );
  OAI21_X1 u2_u6_u1_U62 (.ZN( u2_u6_u1_n109 ) , .B1( u2_u6_u1_n129 ) , .B2( u2_u6_u1_n160 ) , .A( u2_u6_u1_n167 ) );
  NAND2_X1 u2_u6_u1_U63 (.A2( u2_u6_u1_n100 ) , .A1( u2_u6_u1_n103 ) , .ZN( u2_u6_u1_n120 ) );
  NAND2_X1 u2_u6_u1_U64 (.A1( u2_u6_u1_n102 ) , .A2( u2_u6_u1_n104 ) , .ZN( u2_u6_u1_n115 ) );
  NAND2_X1 u2_u6_u1_U65 (.A2( u2_u6_u1_n100 ) , .A1( u2_u6_u1_n104 ) , .ZN( u2_u6_u1_n151 ) );
  NAND2_X1 u2_u6_u1_U66 (.A2( u2_u6_u1_n103 ) , .A1( u2_u6_u1_n105 ) , .ZN( u2_u6_u1_n161 ) );
  INV_X1 u2_u6_u1_U67 (.A( u2_u6_u1_n152 ) , .ZN( u2_u6_u1_n173 ) );
  INV_X1 u2_u6_u1_U68 (.A( u2_u6_u1_n128 ) , .ZN( u2_u6_u1_n172 ) );
  NAND2_X1 u2_u6_u1_U69 (.A2( u2_u6_u1_n102 ) , .A1( u2_u6_u1_n103 ) , .ZN( u2_u6_u1_n123 ) );
  INV_X1 u2_u6_u1_U7 (.A( u2_u6_u1_n147 ) , .ZN( u2_u6_u1_n181 ) );
  NOR2_X1 u2_u6_u1_U70 (.A2( u2_u6_X_7 ) , .A1( u2_u6_X_8 ) , .ZN( u2_u6_u1_n95 ) );
  NOR2_X1 u2_u6_u1_U71 (.A1( u2_u6_X_12 ) , .A2( u2_u6_X_9 ) , .ZN( u2_u6_u1_n100 ) );
  NOR2_X1 u2_u6_u1_U72 (.A2( u2_u6_X_8 ) , .A1( u2_u6_u1_n177 ) , .ZN( u2_u6_u1_n99 ) );
  NOR2_X1 u2_u6_u1_U73 (.A2( u2_u6_X_12 ) , .ZN( u2_u6_u1_n102 ) , .A1( u2_u6_u1_n176 ) );
  NOR2_X1 u2_u6_u1_U74 (.A2( u2_u6_X_9 ) , .ZN( u2_u6_u1_n105 ) , .A1( u2_u6_u1_n168 ) );
  NAND2_X1 u2_u6_u1_U75 (.A1( u2_u6_X_10 ) , .ZN( u2_u6_u1_n160 ) , .A2( u2_u6_u1_n169 ) );
  NAND2_X1 u2_u6_u1_U76 (.A2( u2_u6_X_10 ) , .A1( u2_u6_X_11 ) , .ZN( u2_u6_u1_n152 ) );
  NAND2_X1 u2_u6_u1_U77 (.A1( u2_u6_X_11 ) , .ZN( u2_u6_u1_n128 ) , .A2( u2_u6_u1_n170 ) );
  AND2_X1 u2_u6_u1_U78 (.A2( u2_u6_X_7 ) , .A1( u2_u6_X_8 ) , .ZN( u2_u6_u1_n104 ) );
  AND2_X1 u2_u6_u1_U79 (.A1( u2_u6_X_8 ) , .ZN( u2_u6_u1_n103 ) , .A2( u2_u6_u1_n177 ) );
  NOR2_X1 u2_u6_u1_U8 (.A1( u2_u6_u1_n112 ) , .A2( u2_u6_u1_n116 ) , .ZN( u2_u6_u1_n118 ) );
  INV_X1 u2_u6_u1_U80 (.A( u2_u6_X_10 ) , .ZN( u2_u6_u1_n170 ) );
  INV_X1 u2_u6_u1_U81 (.A( u2_u6_X_9 ) , .ZN( u2_u6_u1_n176 ) );
  INV_X1 u2_u6_u1_U82 (.A( u2_u6_X_11 ) , .ZN( u2_u6_u1_n169 ) );
  INV_X1 u2_u6_u1_U83 (.A( u2_u6_X_12 ) , .ZN( u2_u6_u1_n168 ) );
  INV_X1 u2_u6_u1_U84 (.A( u2_u6_X_7 ) , .ZN( u2_u6_u1_n177 ) );
  NAND4_X1 u2_u6_u1_U85 (.ZN( u2_out6_28 ) , .A4( u2_u6_u1_n124 ) , .A3( u2_u6_u1_n125 ) , .A2( u2_u6_u1_n126 ) , .A1( u2_u6_u1_n127 ) );
  OAI21_X1 u2_u6_u1_U86 (.ZN( u2_u6_u1_n127 ) , .B2( u2_u6_u1_n139 ) , .B1( u2_u6_u1_n175 ) , .A( u2_u6_u1_n183 ) );
  OAI21_X1 u2_u6_u1_U87 (.ZN( u2_u6_u1_n126 ) , .B2( u2_u6_u1_n140 ) , .A( u2_u6_u1_n146 ) , .B1( u2_u6_u1_n178 ) );
  NAND4_X1 u2_u6_u1_U88 (.ZN( u2_out6_18 ) , .A4( u2_u6_u1_n165 ) , .A3( u2_u6_u1_n166 ) , .A1( u2_u6_u1_n167 ) , .A2( u2_u6_u1_n186 ) );
  AOI22_X1 u2_u6_u1_U89 (.B2( u2_u6_u1_n146 ) , .B1( u2_u6_u1_n147 ) , .A2( u2_u6_u1_n148 ) , .ZN( u2_u6_u1_n166 ) , .A1( u2_u6_u1_n172 ) );
  OAI21_X1 u2_u6_u1_U9 (.ZN( u2_u6_u1_n101 ) , .B1( u2_u6_u1_n141 ) , .A( u2_u6_u1_n146 ) , .B2( u2_u6_u1_n183 ) );
  INV_X1 u2_u6_u1_U90 (.A( u2_u6_u1_n145 ) , .ZN( u2_u6_u1_n186 ) );
  NAND4_X1 u2_u6_u1_U91 (.ZN( u2_out6_2 ) , .A4( u2_u6_u1_n142 ) , .A3( u2_u6_u1_n143 ) , .A2( u2_u6_u1_n144 ) , .A1( u2_u6_u1_n179 ) );
  OAI21_X1 u2_u6_u1_U92 (.B2( u2_u6_u1_n132 ) , .ZN( u2_u6_u1_n144 ) , .A( u2_u6_u1_n146 ) , .B1( u2_u6_u1_n180 ) );
  INV_X1 u2_u6_u1_U93 (.A( u2_u6_u1_n130 ) , .ZN( u2_u6_u1_n179 ) );
  OR4_X1 u2_u6_u1_U94 (.ZN( u2_out6_13 ) , .A4( u2_u6_u1_n108 ) , .A3( u2_u6_u1_n109 ) , .A2( u2_u6_u1_n110 ) , .A1( u2_u6_u1_n111 ) );
  AOI21_X1 u2_u6_u1_U95 (.ZN( u2_u6_u1_n111 ) , .A( u2_u6_u1_n128 ) , .B2( u2_u6_u1_n131 ) , .B1( u2_u6_u1_n135 ) );
  AOI21_X1 u2_u6_u1_U96 (.ZN( u2_u6_u1_n110 ) , .A( u2_u6_u1_n116 ) , .B1( u2_u6_u1_n152 ) , .B2( u2_u6_u1_n160 ) );
  NAND3_X1 u2_u6_u1_U97 (.A3( u2_u6_u1_n149 ) , .A2( u2_u6_u1_n150 ) , .A1( u2_u6_u1_n151 ) , .ZN( u2_u6_u1_n164 ) );
  NAND3_X1 u2_u6_u1_U98 (.A3( u2_u6_u1_n134 ) , .A2( u2_u6_u1_n135 ) , .ZN( u2_u6_u1_n136 ) , .A1( u2_u6_u1_n151 ) );
  NAND3_X1 u2_u6_u1_U99 (.A1( u2_u6_u1_n133 ) , .ZN( u2_u6_u1_n137 ) , .A2( u2_u6_u1_n154 ) , .A3( u2_u6_u1_n181 ) );
  OAI22_X1 u2_u6_u2_U10 (.B1( u2_u6_u2_n151 ) , .A2( u2_u6_u2_n152 ) , .A1( u2_u6_u2_n153 ) , .ZN( u2_u6_u2_n160 ) , .B2( u2_u6_u2_n168 ) );
  NAND3_X1 u2_u6_u2_U100 (.A2( u2_u6_u2_n100 ) , .A1( u2_u6_u2_n104 ) , .A3( u2_u6_u2_n138 ) , .ZN( u2_u6_u2_n98 ) );
  NOR3_X1 u2_u6_u2_U11 (.A1( u2_u6_u2_n150 ) , .ZN( u2_u6_u2_n151 ) , .A3( u2_u6_u2_n175 ) , .A2( u2_u6_u2_n188 ) );
  AOI21_X1 u2_u6_u2_U12 (.B2( u2_u6_u2_n123 ) , .ZN( u2_u6_u2_n125 ) , .A( u2_u6_u2_n171 ) , .B1( u2_u6_u2_n184 ) );
  INV_X1 u2_u6_u2_U13 (.A( u2_u6_u2_n150 ) , .ZN( u2_u6_u2_n184 ) );
  AOI21_X1 u2_u6_u2_U14 (.ZN( u2_u6_u2_n144 ) , .B2( u2_u6_u2_n155 ) , .A( u2_u6_u2_n172 ) , .B1( u2_u6_u2_n185 ) );
  AOI21_X1 u2_u6_u2_U15 (.B2( u2_u6_u2_n143 ) , .ZN( u2_u6_u2_n145 ) , .B1( u2_u6_u2_n152 ) , .A( u2_u6_u2_n171 ) );
  INV_X1 u2_u6_u2_U16 (.A( u2_u6_u2_n156 ) , .ZN( u2_u6_u2_n171 ) );
  INV_X1 u2_u6_u2_U17 (.A( u2_u6_u2_n120 ) , .ZN( u2_u6_u2_n188 ) );
  NAND2_X1 u2_u6_u2_U18 (.A2( u2_u6_u2_n122 ) , .ZN( u2_u6_u2_n150 ) , .A1( u2_u6_u2_n152 ) );
  INV_X1 u2_u6_u2_U19 (.A( u2_u6_u2_n153 ) , .ZN( u2_u6_u2_n170 ) );
  INV_X1 u2_u6_u2_U20 (.A( u2_u6_u2_n137 ) , .ZN( u2_u6_u2_n173 ) );
  NAND2_X1 u2_u6_u2_U21 (.A1( u2_u6_u2_n132 ) , .A2( u2_u6_u2_n139 ) , .ZN( u2_u6_u2_n157 ) );
  INV_X1 u2_u6_u2_U22 (.A( u2_u6_u2_n113 ) , .ZN( u2_u6_u2_n178 ) );
  INV_X1 u2_u6_u2_U23 (.A( u2_u6_u2_n139 ) , .ZN( u2_u6_u2_n175 ) );
  INV_X1 u2_u6_u2_U24 (.A( u2_u6_u2_n155 ) , .ZN( u2_u6_u2_n181 ) );
  INV_X1 u2_u6_u2_U25 (.A( u2_u6_u2_n119 ) , .ZN( u2_u6_u2_n177 ) );
  INV_X1 u2_u6_u2_U26 (.A( u2_u6_u2_n116 ) , .ZN( u2_u6_u2_n180 ) );
  INV_X1 u2_u6_u2_U27 (.A( u2_u6_u2_n131 ) , .ZN( u2_u6_u2_n179 ) );
  INV_X1 u2_u6_u2_U28 (.A( u2_u6_u2_n154 ) , .ZN( u2_u6_u2_n176 ) );
  NAND2_X1 u2_u6_u2_U29 (.A2( u2_u6_u2_n116 ) , .A1( u2_u6_u2_n117 ) , .ZN( u2_u6_u2_n118 ) );
  NOR2_X1 u2_u6_u2_U3 (.ZN( u2_u6_u2_n121 ) , .A2( u2_u6_u2_n177 ) , .A1( u2_u6_u2_n180 ) );
  INV_X1 u2_u6_u2_U30 (.A( u2_u6_u2_n132 ) , .ZN( u2_u6_u2_n182 ) );
  INV_X1 u2_u6_u2_U31 (.A( u2_u6_u2_n158 ) , .ZN( u2_u6_u2_n183 ) );
  OAI21_X1 u2_u6_u2_U32 (.A( u2_u6_u2_n156 ) , .B1( u2_u6_u2_n157 ) , .ZN( u2_u6_u2_n158 ) , .B2( u2_u6_u2_n179 ) );
  NOR2_X1 u2_u6_u2_U33 (.ZN( u2_u6_u2_n156 ) , .A1( u2_u6_u2_n166 ) , .A2( u2_u6_u2_n169 ) );
  NOR2_X1 u2_u6_u2_U34 (.A2( u2_u6_u2_n114 ) , .ZN( u2_u6_u2_n137 ) , .A1( u2_u6_u2_n140 ) );
  NOR2_X1 u2_u6_u2_U35 (.A2( u2_u6_u2_n138 ) , .ZN( u2_u6_u2_n153 ) , .A1( u2_u6_u2_n156 ) );
  AOI211_X1 u2_u6_u2_U36 (.ZN( u2_u6_u2_n130 ) , .C1( u2_u6_u2_n138 ) , .C2( u2_u6_u2_n179 ) , .B( u2_u6_u2_n96 ) , .A( u2_u6_u2_n97 ) );
  OAI22_X1 u2_u6_u2_U37 (.B1( u2_u6_u2_n133 ) , .A2( u2_u6_u2_n137 ) , .A1( u2_u6_u2_n152 ) , .B2( u2_u6_u2_n168 ) , .ZN( u2_u6_u2_n97 ) );
  OAI221_X1 u2_u6_u2_U38 (.B1( u2_u6_u2_n113 ) , .C1( u2_u6_u2_n132 ) , .A( u2_u6_u2_n149 ) , .B2( u2_u6_u2_n171 ) , .C2( u2_u6_u2_n172 ) , .ZN( u2_u6_u2_n96 ) );
  OAI221_X1 u2_u6_u2_U39 (.A( u2_u6_u2_n115 ) , .C2( u2_u6_u2_n123 ) , .B2( u2_u6_u2_n143 ) , .B1( u2_u6_u2_n153 ) , .ZN( u2_u6_u2_n163 ) , .C1( u2_u6_u2_n168 ) );
  INV_X1 u2_u6_u2_U4 (.A( u2_u6_u2_n134 ) , .ZN( u2_u6_u2_n185 ) );
  OAI21_X1 u2_u6_u2_U40 (.A( u2_u6_u2_n114 ) , .ZN( u2_u6_u2_n115 ) , .B1( u2_u6_u2_n176 ) , .B2( u2_u6_u2_n178 ) );
  OAI221_X1 u2_u6_u2_U41 (.A( u2_u6_u2_n135 ) , .B2( u2_u6_u2_n136 ) , .B1( u2_u6_u2_n137 ) , .ZN( u2_u6_u2_n162 ) , .C2( u2_u6_u2_n167 ) , .C1( u2_u6_u2_n185 ) );
  AND3_X1 u2_u6_u2_U42 (.A3( u2_u6_u2_n131 ) , .A2( u2_u6_u2_n132 ) , .A1( u2_u6_u2_n133 ) , .ZN( u2_u6_u2_n136 ) );
  AOI22_X1 u2_u6_u2_U43 (.ZN( u2_u6_u2_n135 ) , .B1( u2_u6_u2_n140 ) , .A1( u2_u6_u2_n156 ) , .B2( u2_u6_u2_n180 ) , .A2( u2_u6_u2_n188 ) );
  AOI21_X1 u2_u6_u2_U44 (.ZN( u2_u6_u2_n149 ) , .B1( u2_u6_u2_n173 ) , .B2( u2_u6_u2_n188 ) , .A( u2_u6_u2_n95 ) );
  AND3_X1 u2_u6_u2_U45 (.A2( u2_u6_u2_n100 ) , .A1( u2_u6_u2_n104 ) , .A3( u2_u6_u2_n156 ) , .ZN( u2_u6_u2_n95 ) );
  OAI21_X1 u2_u6_u2_U46 (.A( u2_u6_u2_n141 ) , .B2( u2_u6_u2_n142 ) , .ZN( u2_u6_u2_n146 ) , .B1( u2_u6_u2_n153 ) );
  OAI21_X1 u2_u6_u2_U47 (.A( u2_u6_u2_n140 ) , .ZN( u2_u6_u2_n141 ) , .B1( u2_u6_u2_n176 ) , .B2( u2_u6_u2_n177 ) );
  NOR3_X1 u2_u6_u2_U48 (.ZN( u2_u6_u2_n142 ) , .A3( u2_u6_u2_n175 ) , .A2( u2_u6_u2_n178 ) , .A1( u2_u6_u2_n181 ) );
  OAI21_X1 u2_u6_u2_U49 (.A( u2_u6_u2_n101 ) , .B2( u2_u6_u2_n121 ) , .B1( u2_u6_u2_n153 ) , .ZN( u2_u6_u2_n164 ) );
  NOR4_X1 u2_u6_u2_U5 (.A4( u2_u6_u2_n124 ) , .A3( u2_u6_u2_n125 ) , .A2( u2_u6_u2_n126 ) , .A1( u2_u6_u2_n127 ) , .ZN( u2_u6_u2_n128 ) );
  NAND2_X1 u2_u6_u2_U50 (.A2( u2_u6_u2_n100 ) , .A1( u2_u6_u2_n107 ) , .ZN( u2_u6_u2_n155 ) );
  NAND2_X1 u2_u6_u2_U51 (.A2( u2_u6_u2_n105 ) , .A1( u2_u6_u2_n108 ) , .ZN( u2_u6_u2_n143 ) );
  NAND2_X1 u2_u6_u2_U52 (.A1( u2_u6_u2_n104 ) , .A2( u2_u6_u2_n106 ) , .ZN( u2_u6_u2_n152 ) );
  NAND2_X1 u2_u6_u2_U53 (.A1( u2_u6_u2_n100 ) , .A2( u2_u6_u2_n105 ) , .ZN( u2_u6_u2_n132 ) );
  INV_X1 u2_u6_u2_U54 (.A( u2_u6_u2_n140 ) , .ZN( u2_u6_u2_n168 ) );
  INV_X1 u2_u6_u2_U55 (.A( u2_u6_u2_n138 ) , .ZN( u2_u6_u2_n167 ) );
  INV_X1 u2_u6_u2_U56 (.ZN( u2_u6_u2_n187 ) , .A( u2_u6_u2_n99 ) );
  OAI21_X1 u2_u6_u2_U57 (.B1( u2_u6_u2_n137 ) , .B2( u2_u6_u2_n143 ) , .A( u2_u6_u2_n98 ) , .ZN( u2_u6_u2_n99 ) );
  NAND2_X1 u2_u6_u2_U58 (.A1( u2_u6_u2_n102 ) , .A2( u2_u6_u2_n106 ) , .ZN( u2_u6_u2_n113 ) );
  NAND2_X1 u2_u6_u2_U59 (.A1( u2_u6_u2_n106 ) , .A2( u2_u6_u2_n107 ) , .ZN( u2_u6_u2_n131 ) );
  AOI21_X1 u2_u6_u2_U6 (.B2( u2_u6_u2_n119 ) , .ZN( u2_u6_u2_n127 ) , .A( u2_u6_u2_n137 ) , .B1( u2_u6_u2_n155 ) );
  NAND2_X1 u2_u6_u2_U60 (.A1( u2_u6_u2_n103 ) , .A2( u2_u6_u2_n107 ) , .ZN( u2_u6_u2_n139 ) );
  NAND2_X1 u2_u6_u2_U61 (.A1( u2_u6_u2_n103 ) , .A2( u2_u6_u2_n105 ) , .ZN( u2_u6_u2_n133 ) );
  NAND2_X1 u2_u6_u2_U62 (.A1( u2_u6_u2_n102 ) , .A2( u2_u6_u2_n103 ) , .ZN( u2_u6_u2_n154 ) );
  NAND2_X1 u2_u6_u2_U63 (.A2( u2_u6_u2_n103 ) , .A1( u2_u6_u2_n104 ) , .ZN( u2_u6_u2_n119 ) );
  NAND2_X1 u2_u6_u2_U64 (.A2( u2_u6_u2_n107 ) , .A1( u2_u6_u2_n108 ) , .ZN( u2_u6_u2_n123 ) );
  NAND2_X1 u2_u6_u2_U65 (.A1( u2_u6_u2_n104 ) , .A2( u2_u6_u2_n108 ) , .ZN( u2_u6_u2_n122 ) );
  INV_X1 u2_u6_u2_U66 (.A( u2_u6_u2_n114 ) , .ZN( u2_u6_u2_n172 ) );
  NAND2_X1 u2_u6_u2_U67 (.A2( u2_u6_u2_n100 ) , .A1( u2_u6_u2_n102 ) , .ZN( u2_u6_u2_n116 ) );
  NAND2_X1 u2_u6_u2_U68 (.A1( u2_u6_u2_n102 ) , .A2( u2_u6_u2_n108 ) , .ZN( u2_u6_u2_n120 ) );
  NAND2_X1 u2_u6_u2_U69 (.A2( u2_u6_u2_n105 ) , .A1( u2_u6_u2_n106 ) , .ZN( u2_u6_u2_n117 ) );
  AOI21_X1 u2_u6_u2_U7 (.ZN( u2_u6_u2_n124 ) , .B1( u2_u6_u2_n131 ) , .B2( u2_u6_u2_n143 ) , .A( u2_u6_u2_n172 ) );
  NOR2_X1 u2_u6_u2_U70 (.A2( u2_u6_X_16 ) , .ZN( u2_u6_u2_n140 ) , .A1( u2_u6_u2_n166 ) );
  NOR2_X1 u2_u6_u2_U71 (.A2( u2_u6_X_13 ) , .A1( u2_u6_X_14 ) , .ZN( u2_u6_u2_n100 ) );
  NOR2_X1 u2_u6_u2_U72 (.A2( u2_u6_X_16 ) , .A1( u2_u6_X_17 ) , .ZN( u2_u6_u2_n138 ) );
  NOR2_X1 u2_u6_u2_U73 (.A2( u2_u6_X_15 ) , .A1( u2_u6_X_18 ) , .ZN( u2_u6_u2_n104 ) );
  NOR2_X1 u2_u6_u2_U74 (.A2( u2_u6_X_14 ) , .ZN( u2_u6_u2_n103 ) , .A1( u2_u6_u2_n174 ) );
  NOR2_X1 u2_u6_u2_U75 (.A2( u2_u6_X_15 ) , .ZN( u2_u6_u2_n102 ) , .A1( u2_u6_u2_n165 ) );
  NOR2_X1 u2_u6_u2_U76 (.A2( u2_u6_X_17 ) , .ZN( u2_u6_u2_n114 ) , .A1( u2_u6_u2_n169 ) );
  AND2_X1 u2_u6_u2_U77 (.A1( u2_u6_X_15 ) , .ZN( u2_u6_u2_n105 ) , .A2( u2_u6_u2_n165 ) );
  AND2_X1 u2_u6_u2_U78 (.A2( u2_u6_X_15 ) , .A1( u2_u6_X_18 ) , .ZN( u2_u6_u2_n107 ) );
  AND2_X1 u2_u6_u2_U79 (.A1( u2_u6_X_14 ) , .ZN( u2_u6_u2_n106 ) , .A2( u2_u6_u2_n174 ) );
  AOI21_X1 u2_u6_u2_U8 (.B2( u2_u6_u2_n120 ) , .B1( u2_u6_u2_n121 ) , .ZN( u2_u6_u2_n126 ) , .A( u2_u6_u2_n167 ) );
  AND2_X1 u2_u6_u2_U80 (.A1( u2_u6_X_13 ) , .A2( u2_u6_X_14 ) , .ZN( u2_u6_u2_n108 ) );
  INV_X1 u2_u6_u2_U81 (.A( u2_u6_X_16 ) , .ZN( u2_u6_u2_n169 ) );
  INV_X1 u2_u6_u2_U82 (.A( u2_u6_X_17 ) , .ZN( u2_u6_u2_n166 ) );
  INV_X1 u2_u6_u2_U83 (.A( u2_u6_X_13 ) , .ZN( u2_u6_u2_n174 ) );
  INV_X1 u2_u6_u2_U84 (.A( u2_u6_X_18 ) , .ZN( u2_u6_u2_n165 ) );
  NAND4_X1 u2_u6_u2_U85 (.ZN( u2_out6_30 ) , .A4( u2_u6_u2_n147 ) , .A3( u2_u6_u2_n148 ) , .A2( u2_u6_u2_n149 ) , .A1( u2_u6_u2_n187 ) );
  AOI21_X1 u2_u6_u2_U86 (.B2( u2_u6_u2_n138 ) , .ZN( u2_u6_u2_n148 ) , .A( u2_u6_u2_n162 ) , .B1( u2_u6_u2_n182 ) );
  NOR3_X1 u2_u6_u2_U87 (.A3( u2_u6_u2_n144 ) , .A2( u2_u6_u2_n145 ) , .A1( u2_u6_u2_n146 ) , .ZN( u2_u6_u2_n147 ) );
  NAND4_X1 u2_u6_u2_U88 (.ZN( u2_out6_24 ) , .A4( u2_u6_u2_n111 ) , .A3( u2_u6_u2_n112 ) , .A1( u2_u6_u2_n130 ) , .A2( u2_u6_u2_n187 ) );
  AOI221_X1 u2_u6_u2_U89 (.A( u2_u6_u2_n109 ) , .B1( u2_u6_u2_n110 ) , .ZN( u2_u6_u2_n111 ) , .C1( u2_u6_u2_n134 ) , .C2( u2_u6_u2_n170 ) , .B2( u2_u6_u2_n173 ) );
  OAI22_X1 u2_u6_u2_U9 (.ZN( u2_u6_u2_n109 ) , .A2( u2_u6_u2_n113 ) , .B2( u2_u6_u2_n133 ) , .B1( u2_u6_u2_n167 ) , .A1( u2_u6_u2_n168 ) );
  AOI21_X1 u2_u6_u2_U90 (.ZN( u2_u6_u2_n112 ) , .B2( u2_u6_u2_n156 ) , .A( u2_u6_u2_n164 ) , .B1( u2_u6_u2_n181 ) );
  NAND4_X1 u2_u6_u2_U91 (.ZN( u2_out6_16 ) , .A4( u2_u6_u2_n128 ) , .A3( u2_u6_u2_n129 ) , .A1( u2_u6_u2_n130 ) , .A2( u2_u6_u2_n186 ) );
  AOI22_X1 u2_u6_u2_U92 (.A2( u2_u6_u2_n118 ) , .ZN( u2_u6_u2_n129 ) , .A1( u2_u6_u2_n140 ) , .B1( u2_u6_u2_n157 ) , .B2( u2_u6_u2_n170 ) );
  INV_X1 u2_u6_u2_U93 (.A( u2_u6_u2_n163 ) , .ZN( u2_u6_u2_n186 ) );
  OR4_X1 u2_u6_u2_U94 (.ZN( u2_out6_6 ) , .A4( u2_u6_u2_n161 ) , .A3( u2_u6_u2_n162 ) , .A2( u2_u6_u2_n163 ) , .A1( u2_u6_u2_n164 ) );
  OR3_X1 u2_u6_u2_U95 (.A2( u2_u6_u2_n159 ) , .A1( u2_u6_u2_n160 ) , .ZN( u2_u6_u2_n161 ) , .A3( u2_u6_u2_n183 ) );
  AOI21_X1 u2_u6_u2_U96 (.B2( u2_u6_u2_n154 ) , .B1( u2_u6_u2_n155 ) , .ZN( u2_u6_u2_n159 ) , .A( u2_u6_u2_n167 ) );
  NAND3_X1 u2_u6_u2_U97 (.A2( u2_u6_u2_n117 ) , .A1( u2_u6_u2_n122 ) , .A3( u2_u6_u2_n123 ) , .ZN( u2_u6_u2_n134 ) );
  NAND3_X1 u2_u6_u2_U98 (.ZN( u2_u6_u2_n110 ) , .A2( u2_u6_u2_n131 ) , .A3( u2_u6_u2_n139 ) , .A1( u2_u6_u2_n154 ) );
  NAND3_X1 u2_u6_u2_U99 (.A2( u2_u6_u2_n100 ) , .ZN( u2_u6_u2_n101 ) , .A1( u2_u6_u2_n104 ) , .A3( u2_u6_u2_n114 ) );
  OAI22_X1 u2_u6_u3_U10 (.B1( u2_u6_u3_n113 ) , .A2( u2_u6_u3_n135 ) , .A1( u2_u6_u3_n150 ) , .B2( u2_u6_u3_n164 ) , .ZN( u2_u6_u3_n98 ) );
  OAI211_X1 u2_u6_u3_U11 (.B( u2_u6_u3_n106 ) , .ZN( u2_u6_u3_n119 ) , .C2( u2_u6_u3_n128 ) , .C1( u2_u6_u3_n167 ) , .A( u2_u6_u3_n181 ) );
  AOI221_X1 u2_u6_u3_U12 (.C1( u2_u6_u3_n105 ) , .ZN( u2_u6_u3_n106 ) , .A( u2_u6_u3_n131 ) , .B2( u2_u6_u3_n132 ) , .C2( u2_u6_u3_n133 ) , .B1( u2_u6_u3_n169 ) );
  INV_X1 u2_u6_u3_U13 (.ZN( u2_u6_u3_n181 ) , .A( u2_u6_u3_n98 ) );
  NAND2_X1 u2_u6_u3_U14 (.ZN( u2_u6_u3_n105 ) , .A2( u2_u6_u3_n130 ) , .A1( u2_u6_u3_n155 ) );
  NOR2_X1 u2_u6_u3_U15 (.ZN( u2_u6_u3_n126 ) , .A2( u2_u6_u3_n150 ) , .A1( u2_u6_u3_n164 ) );
  AOI21_X1 u2_u6_u3_U16 (.ZN( u2_u6_u3_n112 ) , .B2( u2_u6_u3_n146 ) , .B1( u2_u6_u3_n155 ) , .A( u2_u6_u3_n167 ) );
  NAND2_X1 u2_u6_u3_U17 (.A1( u2_u6_u3_n135 ) , .ZN( u2_u6_u3_n142 ) , .A2( u2_u6_u3_n164 ) );
  NAND2_X1 u2_u6_u3_U18 (.ZN( u2_u6_u3_n132 ) , .A2( u2_u6_u3_n152 ) , .A1( u2_u6_u3_n156 ) );
  AND2_X1 u2_u6_u3_U19 (.A2( u2_u6_u3_n113 ) , .A1( u2_u6_u3_n114 ) , .ZN( u2_u6_u3_n151 ) );
  INV_X1 u2_u6_u3_U20 (.A( u2_u6_u3_n133 ) , .ZN( u2_u6_u3_n165 ) );
  INV_X1 u2_u6_u3_U21 (.A( u2_u6_u3_n135 ) , .ZN( u2_u6_u3_n170 ) );
  NAND2_X1 u2_u6_u3_U22 (.A1( u2_u6_u3_n107 ) , .A2( u2_u6_u3_n108 ) , .ZN( u2_u6_u3_n140 ) );
  NAND2_X1 u2_u6_u3_U23 (.ZN( u2_u6_u3_n117 ) , .A1( u2_u6_u3_n124 ) , .A2( u2_u6_u3_n148 ) );
  NAND2_X1 u2_u6_u3_U24 (.ZN( u2_u6_u3_n143 ) , .A1( u2_u6_u3_n165 ) , .A2( u2_u6_u3_n167 ) );
  INV_X1 u2_u6_u3_U25 (.A( u2_u6_u3_n130 ) , .ZN( u2_u6_u3_n177 ) );
  INV_X1 u2_u6_u3_U26 (.A( u2_u6_u3_n128 ) , .ZN( u2_u6_u3_n176 ) );
  INV_X1 u2_u6_u3_U27 (.A( u2_u6_u3_n155 ) , .ZN( u2_u6_u3_n174 ) );
  AOI22_X1 u2_u6_u3_U28 (.B1( u2_u6_u3_n115 ) , .A2( u2_u6_u3_n116 ) , .ZN( u2_u6_u3_n123 ) , .B2( u2_u6_u3_n133 ) , .A1( u2_u6_u3_n169 ) );
  NAND2_X1 u2_u6_u3_U29 (.ZN( u2_u6_u3_n116 ) , .A2( u2_u6_u3_n151 ) , .A1( u2_u6_u3_n182 ) );
  INV_X1 u2_u6_u3_U3 (.A( u2_u6_u3_n129 ) , .ZN( u2_u6_u3_n183 ) );
  INV_X1 u2_u6_u3_U30 (.A( u2_u6_u3_n139 ) , .ZN( u2_u6_u3_n185 ) );
  NOR2_X1 u2_u6_u3_U31 (.ZN( u2_u6_u3_n135 ) , .A2( u2_u6_u3_n141 ) , .A1( u2_u6_u3_n169 ) );
  OAI222_X1 u2_u6_u3_U32 (.C2( u2_u6_u3_n107 ) , .A2( u2_u6_u3_n108 ) , .B1( u2_u6_u3_n135 ) , .ZN( u2_u6_u3_n138 ) , .B2( u2_u6_u3_n146 ) , .C1( u2_u6_u3_n154 ) , .A1( u2_u6_u3_n164 ) );
  NOR4_X1 u2_u6_u3_U33 (.A4( u2_u6_u3_n157 ) , .A3( u2_u6_u3_n158 ) , .A2( u2_u6_u3_n159 ) , .A1( u2_u6_u3_n160 ) , .ZN( u2_u6_u3_n161 ) );
  AOI21_X1 u2_u6_u3_U34 (.B2( u2_u6_u3_n152 ) , .B1( u2_u6_u3_n153 ) , .ZN( u2_u6_u3_n158 ) , .A( u2_u6_u3_n164 ) );
  AOI21_X1 u2_u6_u3_U35 (.A( u2_u6_u3_n154 ) , .B2( u2_u6_u3_n155 ) , .B1( u2_u6_u3_n156 ) , .ZN( u2_u6_u3_n157 ) );
  AOI21_X1 u2_u6_u3_U36 (.A( u2_u6_u3_n149 ) , .B2( u2_u6_u3_n150 ) , .B1( u2_u6_u3_n151 ) , .ZN( u2_u6_u3_n159 ) );
  AOI211_X1 u2_u6_u3_U37 (.ZN( u2_u6_u3_n109 ) , .A( u2_u6_u3_n119 ) , .C2( u2_u6_u3_n129 ) , .B( u2_u6_u3_n138 ) , .C1( u2_u6_u3_n141 ) );
  AOI211_X1 u2_u6_u3_U38 (.B( u2_u6_u3_n119 ) , .A( u2_u6_u3_n120 ) , .C2( u2_u6_u3_n121 ) , .ZN( u2_u6_u3_n122 ) , .C1( u2_u6_u3_n179 ) );
  INV_X1 u2_u6_u3_U39 (.A( u2_u6_u3_n156 ) , .ZN( u2_u6_u3_n179 ) );
  INV_X1 u2_u6_u3_U4 (.A( u2_u6_u3_n140 ) , .ZN( u2_u6_u3_n182 ) );
  OAI22_X1 u2_u6_u3_U40 (.B1( u2_u6_u3_n118 ) , .ZN( u2_u6_u3_n120 ) , .A1( u2_u6_u3_n135 ) , .B2( u2_u6_u3_n154 ) , .A2( u2_u6_u3_n178 ) );
  AND3_X1 u2_u6_u3_U41 (.ZN( u2_u6_u3_n118 ) , .A2( u2_u6_u3_n124 ) , .A1( u2_u6_u3_n144 ) , .A3( u2_u6_u3_n152 ) );
  INV_X1 u2_u6_u3_U42 (.A( u2_u6_u3_n121 ) , .ZN( u2_u6_u3_n164 ) );
  NAND2_X1 u2_u6_u3_U43 (.ZN( u2_u6_u3_n133 ) , .A1( u2_u6_u3_n154 ) , .A2( u2_u6_u3_n164 ) );
  OAI211_X1 u2_u6_u3_U44 (.B( u2_u6_u3_n127 ) , .ZN( u2_u6_u3_n139 ) , .C1( u2_u6_u3_n150 ) , .C2( u2_u6_u3_n154 ) , .A( u2_u6_u3_n184 ) );
  INV_X1 u2_u6_u3_U45 (.A( u2_u6_u3_n125 ) , .ZN( u2_u6_u3_n184 ) );
  AOI221_X1 u2_u6_u3_U46 (.A( u2_u6_u3_n126 ) , .ZN( u2_u6_u3_n127 ) , .C2( u2_u6_u3_n132 ) , .C1( u2_u6_u3_n169 ) , .B2( u2_u6_u3_n170 ) , .B1( u2_u6_u3_n174 ) );
  OAI22_X1 u2_u6_u3_U47 (.A1( u2_u6_u3_n124 ) , .ZN( u2_u6_u3_n125 ) , .B2( u2_u6_u3_n145 ) , .A2( u2_u6_u3_n165 ) , .B1( u2_u6_u3_n167 ) );
  NOR2_X1 u2_u6_u3_U48 (.A1( u2_u6_u3_n113 ) , .ZN( u2_u6_u3_n131 ) , .A2( u2_u6_u3_n154 ) );
  NAND2_X1 u2_u6_u3_U49 (.A1( u2_u6_u3_n103 ) , .ZN( u2_u6_u3_n150 ) , .A2( u2_u6_u3_n99 ) );
  INV_X1 u2_u6_u3_U5 (.A( u2_u6_u3_n117 ) , .ZN( u2_u6_u3_n178 ) );
  NAND2_X1 u2_u6_u3_U50 (.A2( u2_u6_u3_n102 ) , .ZN( u2_u6_u3_n155 ) , .A1( u2_u6_u3_n97 ) );
  INV_X1 u2_u6_u3_U51 (.A( u2_u6_u3_n141 ) , .ZN( u2_u6_u3_n167 ) );
  AOI21_X1 u2_u6_u3_U52 (.B2( u2_u6_u3_n114 ) , .B1( u2_u6_u3_n146 ) , .A( u2_u6_u3_n154 ) , .ZN( u2_u6_u3_n94 ) );
  AOI21_X1 u2_u6_u3_U53 (.ZN( u2_u6_u3_n110 ) , .B2( u2_u6_u3_n142 ) , .B1( u2_u6_u3_n186 ) , .A( u2_u6_u3_n95 ) );
  INV_X1 u2_u6_u3_U54 (.A( u2_u6_u3_n145 ) , .ZN( u2_u6_u3_n186 ) );
  AOI21_X1 u2_u6_u3_U55 (.B1( u2_u6_u3_n124 ) , .A( u2_u6_u3_n149 ) , .B2( u2_u6_u3_n155 ) , .ZN( u2_u6_u3_n95 ) );
  INV_X1 u2_u6_u3_U56 (.A( u2_u6_u3_n149 ) , .ZN( u2_u6_u3_n169 ) );
  NAND2_X1 u2_u6_u3_U57 (.ZN( u2_u6_u3_n124 ) , .A1( u2_u6_u3_n96 ) , .A2( u2_u6_u3_n97 ) );
  NAND2_X1 u2_u6_u3_U58 (.A2( u2_u6_u3_n100 ) , .ZN( u2_u6_u3_n146 ) , .A1( u2_u6_u3_n96 ) );
  NAND2_X1 u2_u6_u3_U59 (.A1( u2_u6_u3_n101 ) , .ZN( u2_u6_u3_n145 ) , .A2( u2_u6_u3_n99 ) );
  AOI221_X1 u2_u6_u3_U6 (.A( u2_u6_u3_n131 ) , .C2( u2_u6_u3_n132 ) , .C1( u2_u6_u3_n133 ) , .ZN( u2_u6_u3_n134 ) , .B1( u2_u6_u3_n143 ) , .B2( u2_u6_u3_n177 ) );
  NAND2_X1 u2_u6_u3_U60 (.A1( u2_u6_u3_n100 ) , .ZN( u2_u6_u3_n156 ) , .A2( u2_u6_u3_n99 ) );
  NAND2_X1 u2_u6_u3_U61 (.A2( u2_u6_u3_n101 ) , .A1( u2_u6_u3_n104 ) , .ZN( u2_u6_u3_n148 ) );
  NAND2_X1 u2_u6_u3_U62 (.A1( u2_u6_u3_n100 ) , .A2( u2_u6_u3_n102 ) , .ZN( u2_u6_u3_n128 ) );
  NAND2_X1 u2_u6_u3_U63 (.A2( u2_u6_u3_n101 ) , .A1( u2_u6_u3_n102 ) , .ZN( u2_u6_u3_n152 ) );
  NAND2_X1 u2_u6_u3_U64 (.A2( u2_u6_u3_n101 ) , .ZN( u2_u6_u3_n114 ) , .A1( u2_u6_u3_n96 ) );
  NAND2_X1 u2_u6_u3_U65 (.ZN( u2_u6_u3_n107 ) , .A1( u2_u6_u3_n97 ) , .A2( u2_u6_u3_n99 ) );
  NAND2_X1 u2_u6_u3_U66 (.A2( u2_u6_u3_n100 ) , .A1( u2_u6_u3_n104 ) , .ZN( u2_u6_u3_n113 ) );
  NAND2_X1 u2_u6_u3_U67 (.A1( u2_u6_u3_n104 ) , .ZN( u2_u6_u3_n153 ) , .A2( u2_u6_u3_n97 ) );
  NAND2_X1 u2_u6_u3_U68 (.A2( u2_u6_u3_n103 ) , .A1( u2_u6_u3_n104 ) , .ZN( u2_u6_u3_n130 ) );
  NAND2_X1 u2_u6_u3_U69 (.A2( u2_u6_u3_n103 ) , .ZN( u2_u6_u3_n144 ) , .A1( u2_u6_u3_n96 ) );
  OAI22_X1 u2_u6_u3_U7 (.B2( u2_u6_u3_n147 ) , .A2( u2_u6_u3_n148 ) , .ZN( u2_u6_u3_n160 ) , .B1( u2_u6_u3_n165 ) , .A1( u2_u6_u3_n168 ) );
  NAND2_X1 u2_u6_u3_U70 (.A1( u2_u6_u3_n102 ) , .A2( u2_u6_u3_n103 ) , .ZN( u2_u6_u3_n108 ) );
  NOR2_X1 u2_u6_u3_U71 (.A2( u2_u6_X_19 ) , .A1( u2_u6_X_20 ) , .ZN( u2_u6_u3_n99 ) );
  NOR2_X1 u2_u6_u3_U72 (.A2( u2_u6_X_21 ) , .A1( u2_u6_X_24 ) , .ZN( u2_u6_u3_n103 ) );
  NOR2_X1 u2_u6_u3_U73 (.A2( u2_u6_X_24 ) , .A1( u2_u6_u3_n171 ) , .ZN( u2_u6_u3_n97 ) );
  NOR2_X1 u2_u6_u3_U74 (.A2( u2_u6_X_23 ) , .ZN( u2_u6_u3_n141 ) , .A1( u2_u6_u3_n166 ) );
  NOR2_X1 u2_u6_u3_U75 (.A2( u2_u6_X_19 ) , .A1( u2_u6_u3_n172 ) , .ZN( u2_u6_u3_n96 ) );
  NAND2_X1 u2_u6_u3_U76 (.A1( u2_u6_X_22 ) , .A2( u2_u6_X_23 ) , .ZN( u2_u6_u3_n154 ) );
  NAND2_X1 u2_u6_u3_U77 (.A1( u2_u6_X_23 ) , .ZN( u2_u6_u3_n149 ) , .A2( u2_u6_u3_n166 ) );
  NOR2_X1 u2_u6_u3_U78 (.A2( u2_u6_X_22 ) , .A1( u2_u6_X_23 ) , .ZN( u2_u6_u3_n121 ) );
  AND2_X1 u2_u6_u3_U79 (.A1( u2_u6_X_24 ) , .ZN( u2_u6_u3_n101 ) , .A2( u2_u6_u3_n171 ) );
  AND3_X1 u2_u6_u3_U8 (.A3( u2_u6_u3_n144 ) , .A2( u2_u6_u3_n145 ) , .A1( u2_u6_u3_n146 ) , .ZN( u2_u6_u3_n147 ) );
  AND2_X1 u2_u6_u3_U80 (.A1( u2_u6_X_19 ) , .ZN( u2_u6_u3_n102 ) , .A2( u2_u6_u3_n172 ) );
  AND2_X1 u2_u6_u3_U81 (.A1( u2_u6_X_21 ) , .A2( u2_u6_X_24 ) , .ZN( u2_u6_u3_n100 ) );
  AND2_X1 u2_u6_u3_U82 (.A2( u2_u6_X_19 ) , .A1( u2_u6_X_20 ) , .ZN( u2_u6_u3_n104 ) );
  INV_X1 u2_u6_u3_U83 (.A( u2_u6_X_22 ) , .ZN( u2_u6_u3_n166 ) );
  INV_X1 u2_u6_u3_U84 (.A( u2_u6_X_21 ) , .ZN( u2_u6_u3_n171 ) );
  INV_X1 u2_u6_u3_U85 (.A( u2_u6_X_20 ) , .ZN( u2_u6_u3_n172 ) );
  NAND4_X1 u2_u6_u3_U86 (.ZN( u2_out6_26 ) , .A4( u2_u6_u3_n109 ) , .A3( u2_u6_u3_n110 ) , .A2( u2_u6_u3_n111 ) , .A1( u2_u6_u3_n173 ) );
  INV_X1 u2_u6_u3_U87 (.ZN( u2_u6_u3_n173 ) , .A( u2_u6_u3_n94 ) );
  OAI21_X1 u2_u6_u3_U88 (.ZN( u2_u6_u3_n111 ) , .B2( u2_u6_u3_n117 ) , .A( u2_u6_u3_n133 ) , .B1( u2_u6_u3_n176 ) );
  NAND4_X1 u2_u6_u3_U89 (.ZN( u2_out6_20 ) , .A4( u2_u6_u3_n122 ) , .A3( u2_u6_u3_n123 ) , .A1( u2_u6_u3_n175 ) , .A2( u2_u6_u3_n180 ) );
  INV_X1 u2_u6_u3_U9 (.A( u2_u6_u3_n143 ) , .ZN( u2_u6_u3_n168 ) );
  INV_X1 u2_u6_u3_U90 (.A( u2_u6_u3_n126 ) , .ZN( u2_u6_u3_n180 ) );
  INV_X1 u2_u6_u3_U91 (.A( u2_u6_u3_n112 ) , .ZN( u2_u6_u3_n175 ) );
  NAND4_X1 u2_u6_u3_U92 (.ZN( u2_out6_1 ) , .A4( u2_u6_u3_n161 ) , .A3( u2_u6_u3_n162 ) , .A2( u2_u6_u3_n163 ) , .A1( u2_u6_u3_n185 ) );
  NAND2_X1 u2_u6_u3_U93 (.ZN( u2_u6_u3_n163 ) , .A2( u2_u6_u3_n170 ) , .A1( u2_u6_u3_n176 ) );
  AOI22_X1 u2_u6_u3_U94 (.B2( u2_u6_u3_n140 ) , .B1( u2_u6_u3_n141 ) , .A2( u2_u6_u3_n142 ) , .ZN( u2_u6_u3_n162 ) , .A1( u2_u6_u3_n177 ) );
  OR4_X1 u2_u6_u3_U95 (.ZN( u2_out6_10 ) , .A4( u2_u6_u3_n136 ) , .A3( u2_u6_u3_n137 ) , .A1( u2_u6_u3_n138 ) , .A2( u2_u6_u3_n139 ) );
  OAI222_X1 u2_u6_u3_U96 (.C1( u2_u6_u3_n128 ) , .ZN( u2_u6_u3_n137 ) , .B1( u2_u6_u3_n148 ) , .A2( u2_u6_u3_n150 ) , .B2( u2_u6_u3_n154 ) , .C2( u2_u6_u3_n164 ) , .A1( u2_u6_u3_n167 ) );
  OAI221_X1 u2_u6_u3_U97 (.A( u2_u6_u3_n134 ) , .B2( u2_u6_u3_n135 ) , .ZN( u2_u6_u3_n136 ) , .C1( u2_u6_u3_n149 ) , .B1( u2_u6_u3_n151 ) , .C2( u2_u6_u3_n183 ) );
  NAND3_X1 u2_u6_u3_U98 (.A1( u2_u6_u3_n114 ) , .ZN( u2_u6_u3_n115 ) , .A2( u2_u6_u3_n145 ) , .A3( u2_u6_u3_n153 ) );
  NAND3_X1 u2_u6_u3_U99 (.ZN( u2_u6_u3_n129 ) , .A2( u2_u6_u3_n144 ) , .A1( u2_u6_u3_n153 ) , .A3( u2_u6_u3_n182 ) );
  OAI22_X1 u2_u6_u4_U10 (.B2( u2_u6_u4_n135 ) , .ZN( u2_u6_u4_n137 ) , .B1( u2_u6_u4_n153 ) , .A1( u2_u6_u4_n155 ) , .A2( u2_u6_u4_n171 ) );
  AND3_X1 u2_u6_u4_U11 (.A2( u2_u6_u4_n134 ) , .ZN( u2_u6_u4_n135 ) , .A3( u2_u6_u4_n145 ) , .A1( u2_u6_u4_n157 ) );
  NAND2_X1 u2_u6_u4_U12 (.ZN( u2_u6_u4_n132 ) , .A2( u2_u6_u4_n170 ) , .A1( u2_u6_u4_n173 ) );
  AOI21_X1 u2_u6_u4_U13 (.B2( u2_u6_u4_n160 ) , .B1( u2_u6_u4_n161 ) , .ZN( u2_u6_u4_n162 ) , .A( u2_u6_u4_n170 ) );
  AOI21_X1 u2_u6_u4_U14 (.ZN( u2_u6_u4_n107 ) , .B2( u2_u6_u4_n143 ) , .A( u2_u6_u4_n174 ) , .B1( u2_u6_u4_n184 ) );
  AOI21_X1 u2_u6_u4_U15 (.B2( u2_u6_u4_n158 ) , .B1( u2_u6_u4_n159 ) , .ZN( u2_u6_u4_n163 ) , .A( u2_u6_u4_n174 ) );
  AOI21_X1 u2_u6_u4_U16 (.A( u2_u6_u4_n153 ) , .B2( u2_u6_u4_n154 ) , .B1( u2_u6_u4_n155 ) , .ZN( u2_u6_u4_n165 ) );
  AOI21_X1 u2_u6_u4_U17 (.A( u2_u6_u4_n156 ) , .B2( u2_u6_u4_n157 ) , .ZN( u2_u6_u4_n164 ) , .B1( u2_u6_u4_n184 ) );
  INV_X1 u2_u6_u4_U18 (.A( u2_u6_u4_n138 ) , .ZN( u2_u6_u4_n170 ) );
  AND2_X1 u2_u6_u4_U19 (.A2( u2_u6_u4_n120 ) , .ZN( u2_u6_u4_n155 ) , .A1( u2_u6_u4_n160 ) );
  INV_X1 u2_u6_u4_U20 (.A( u2_u6_u4_n156 ) , .ZN( u2_u6_u4_n175 ) );
  NAND2_X1 u2_u6_u4_U21 (.A2( u2_u6_u4_n118 ) , .ZN( u2_u6_u4_n131 ) , .A1( u2_u6_u4_n147 ) );
  NAND2_X1 u2_u6_u4_U22 (.A1( u2_u6_u4_n119 ) , .A2( u2_u6_u4_n120 ) , .ZN( u2_u6_u4_n130 ) );
  NAND2_X1 u2_u6_u4_U23 (.ZN( u2_u6_u4_n117 ) , .A2( u2_u6_u4_n118 ) , .A1( u2_u6_u4_n148 ) );
  NAND2_X1 u2_u6_u4_U24 (.ZN( u2_u6_u4_n129 ) , .A1( u2_u6_u4_n134 ) , .A2( u2_u6_u4_n148 ) );
  AND3_X1 u2_u6_u4_U25 (.A1( u2_u6_u4_n119 ) , .A2( u2_u6_u4_n143 ) , .A3( u2_u6_u4_n154 ) , .ZN( u2_u6_u4_n161 ) );
  AND2_X1 u2_u6_u4_U26 (.A1( u2_u6_u4_n145 ) , .A2( u2_u6_u4_n147 ) , .ZN( u2_u6_u4_n159 ) );
  OR3_X1 u2_u6_u4_U27 (.A3( u2_u6_u4_n114 ) , .A2( u2_u6_u4_n115 ) , .A1( u2_u6_u4_n116 ) , .ZN( u2_u6_u4_n136 ) );
  AOI21_X1 u2_u6_u4_U28 (.A( u2_u6_u4_n113 ) , .ZN( u2_u6_u4_n116 ) , .B2( u2_u6_u4_n173 ) , .B1( u2_u6_u4_n174 ) );
  AOI21_X1 u2_u6_u4_U29 (.ZN( u2_u6_u4_n115 ) , .B2( u2_u6_u4_n145 ) , .B1( u2_u6_u4_n146 ) , .A( u2_u6_u4_n156 ) );
  NOR2_X1 u2_u6_u4_U3 (.ZN( u2_u6_u4_n121 ) , .A1( u2_u6_u4_n181 ) , .A2( u2_u6_u4_n182 ) );
  OAI22_X1 u2_u6_u4_U30 (.ZN( u2_u6_u4_n114 ) , .A2( u2_u6_u4_n121 ) , .B1( u2_u6_u4_n160 ) , .B2( u2_u6_u4_n170 ) , .A1( u2_u6_u4_n171 ) );
  INV_X1 u2_u6_u4_U31 (.A( u2_u6_u4_n158 ) , .ZN( u2_u6_u4_n182 ) );
  INV_X1 u2_u6_u4_U32 (.ZN( u2_u6_u4_n181 ) , .A( u2_u6_u4_n96 ) );
  INV_X1 u2_u6_u4_U33 (.A( u2_u6_u4_n144 ) , .ZN( u2_u6_u4_n179 ) );
  INV_X1 u2_u6_u4_U34 (.A( u2_u6_u4_n157 ) , .ZN( u2_u6_u4_n178 ) );
  NAND2_X1 u2_u6_u4_U35 (.A2( u2_u6_u4_n154 ) , .A1( u2_u6_u4_n96 ) , .ZN( u2_u6_u4_n97 ) );
  INV_X1 u2_u6_u4_U36 (.ZN( u2_u6_u4_n186 ) , .A( u2_u6_u4_n95 ) );
  OAI221_X1 u2_u6_u4_U37 (.C1( u2_u6_u4_n134 ) , .B1( u2_u6_u4_n158 ) , .B2( u2_u6_u4_n171 ) , .C2( u2_u6_u4_n173 ) , .A( u2_u6_u4_n94 ) , .ZN( u2_u6_u4_n95 ) );
  AOI222_X1 u2_u6_u4_U38 (.B2( u2_u6_u4_n132 ) , .A1( u2_u6_u4_n138 ) , .C2( u2_u6_u4_n175 ) , .A2( u2_u6_u4_n179 ) , .C1( u2_u6_u4_n181 ) , .B1( u2_u6_u4_n185 ) , .ZN( u2_u6_u4_n94 ) );
  INV_X1 u2_u6_u4_U39 (.A( u2_u6_u4_n113 ) , .ZN( u2_u6_u4_n185 ) );
  INV_X1 u2_u6_u4_U4 (.A( u2_u6_u4_n117 ) , .ZN( u2_u6_u4_n184 ) );
  INV_X1 u2_u6_u4_U40 (.A( u2_u6_u4_n143 ) , .ZN( u2_u6_u4_n183 ) );
  NOR2_X1 u2_u6_u4_U41 (.ZN( u2_u6_u4_n138 ) , .A1( u2_u6_u4_n168 ) , .A2( u2_u6_u4_n169 ) );
  NOR2_X1 u2_u6_u4_U42 (.A1( u2_u6_u4_n150 ) , .A2( u2_u6_u4_n152 ) , .ZN( u2_u6_u4_n153 ) );
  NOR2_X1 u2_u6_u4_U43 (.A2( u2_u6_u4_n128 ) , .A1( u2_u6_u4_n138 ) , .ZN( u2_u6_u4_n156 ) );
  AOI22_X1 u2_u6_u4_U44 (.B2( u2_u6_u4_n122 ) , .A1( u2_u6_u4_n123 ) , .ZN( u2_u6_u4_n124 ) , .B1( u2_u6_u4_n128 ) , .A2( u2_u6_u4_n172 ) );
  INV_X1 u2_u6_u4_U45 (.A( u2_u6_u4_n153 ) , .ZN( u2_u6_u4_n172 ) );
  NAND2_X1 u2_u6_u4_U46 (.A2( u2_u6_u4_n120 ) , .ZN( u2_u6_u4_n123 ) , .A1( u2_u6_u4_n161 ) );
  AOI22_X1 u2_u6_u4_U47 (.B2( u2_u6_u4_n132 ) , .A2( u2_u6_u4_n133 ) , .ZN( u2_u6_u4_n140 ) , .A1( u2_u6_u4_n150 ) , .B1( u2_u6_u4_n179 ) );
  NAND2_X1 u2_u6_u4_U48 (.ZN( u2_u6_u4_n133 ) , .A2( u2_u6_u4_n146 ) , .A1( u2_u6_u4_n154 ) );
  NAND2_X1 u2_u6_u4_U49 (.A1( u2_u6_u4_n103 ) , .ZN( u2_u6_u4_n154 ) , .A2( u2_u6_u4_n98 ) );
  NOR4_X1 u2_u6_u4_U5 (.A4( u2_u6_u4_n106 ) , .A3( u2_u6_u4_n107 ) , .A2( u2_u6_u4_n108 ) , .A1( u2_u6_u4_n109 ) , .ZN( u2_u6_u4_n110 ) );
  NAND2_X1 u2_u6_u4_U50 (.A1( u2_u6_u4_n101 ) , .ZN( u2_u6_u4_n158 ) , .A2( u2_u6_u4_n99 ) );
  AOI21_X1 u2_u6_u4_U51 (.ZN( u2_u6_u4_n127 ) , .A( u2_u6_u4_n136 ) , .B2( u2_u6_u4_n150 ) , .B1( u2_u6_u4_n180 ) );
  INV_X1 u2_u6_u4_U52 (.A( u2_u6_u4_n160 ) , .ZN( u2_u6_u4_n180 ) );
  NAND2_X1 u2_u6_u4_U53 (.A2( u2_u6_u4_n104 ) , .A1( u2_u6_u4_n105 ) , .ZN( u2_u6_u4_n146 ) );
  NAND2_X1 u2_u6_u4_U54 (.A2( u2_u6_u4_n101 ) , .A1( u2_u6_u4_n102 ) , .ZN( u2_u6_u4_n160 ) );
  NAND2_X1 u2_u6_u4_U55 (.ZN( u2_u6_u4_n134 ) , .A1( u2_u6_u4_n98 ) , .A2( u2_u6_u4_n99 ) );
  NAND2_X1 u2_u6_u4_U56 (.A1( u2_u6_u4_n103 ) , .A2( u2_u6_u4_n104 ) , .ZN( u2_u6_u4_n143 ) );
  NAND2_X1 u2_u6_u4_U57 (.A2( u2_u6_u4_n105 ) , .ZN( u2_u6_u4_n145 ) , .A1( u2_u6_u4_n98 ) );
  NAND2_X1 u2_u6_u4_U58 (.A1( u2_u6_u4_n100 ) , .A2( u2_u6_u4_n105 ) , .ZN( u2_u6_u4_n120 ) );
  NAND2_X1 u2_u6_u4_U59 (.A1( u2_u6_u4_n102 ) , .A2( u2_u6_u4_n104 ) , .ZN( u2_u6_u4_n148 ) );
  AOI21_X1 u2_u6_u4_U6 (.ZN( u2_u6_u4_n106 ) , .B2( u2_u6_u4_n146 ) , .B1( u2_u6_u4_n158 ) , .A( u2_u6_u4_n170 ) );
  NAND2_X1 u2_u6_u4_U60 (.A2( u2_u6_u4_n100 ) , .A1( u2_u6_u4_n103 ) , .ZN( u2_u6_u4_n157 ) );
  INV_X1 u2_u6_u4_U61 (.A( u2_u6_u4_n150 ) , .ZN( u2_u6_u4_n173 ) );
  INV_X1 u2_u6_u4_U62 (.A( u2_u6_u4_n152 ) , .ZN( u2_u6_u4_n171 ) );
  NAND2_X1 u2_u6_u4_U63 (.A1( u2_u6_u4_n100 ) , .ZN( u2_u6_u4_n118 ) , .A2( u2_u6_u4_n99 ) );
  NAND2_X1 u2_u6_u4_U64 (.A2( u2_u6_u4_n100 ) , .A1( u2_u6_u4_n102 ) , .ZN( u2_u6_u4_n144 ) );
  NAND2_X1 u2_u6_u4_U65 (.A2( u2_u6_u4_n101 ) , .A1( u2_u6_u4_n105 ) , .ZN( u2_u6_u4_n96 ) );
  INV_X1 u2_u6_u4_U66 (.A( u2_u6_u4_n128 ) , .ZN( u2_u6_u4_n174 ) );
  NAND2_X1 u2_u6_u4_U67 (.A2( u2_u6_u4_n102 ) , .ZN( u2_u6_u4_n119 ) , .A1( u2_u6_u4_n98 ) );
  NAND2_X1 u2_u6_u4_U68 (.A2( u2_u6_u4_n101 ) , .A1( u2_u6_u4_n103 ) , .ZN( u2_u6_u4_n147 ) );
  NAND2_X1 u2_u6_u4_U69 (.A2( u2_u6_u4_n104 ) , .ZN( u2_u6_u4_n113 ) , .A1( u2_u6_u4_n99 ) );
  AOI21_X1 u2_u6_u4_U7 (.ZN( u2_u6_u4_n108 ) , .B2( u2_u6_u4_n134 ) , .B1( u2_u6_u4_n155 ) , .A( u2_u6_u4_n156 ) );
  NOR2_X1 u2_u6_u4_U70 (.A2( u2_u6_X_28 ) , .ZN( u2_u6_u4_n150 ) , .A1( u2_u6_u4_n168 ) );
  NOR2_X1 u2_u6_u4_U71 (.A2( u2_u6_X_29 ) , .ZN( u2_u6_u4_n152 ) , .A1( u2_u6_u4_n169 ) );
  NOR2_X1 u2_u6_u4_U72 (.A2( u2_u6_X_30 ) , .ZN( u2_u6_u4_n105 ) , .A1( u2_u6_u4_n176 ) );
  NOR2_X1 u2_u6_u4_U73 (.A2( u2_u6_X_26 ) , .ZN( u2_u6_u4_n100 ) , .A1( u2_u6_u4_n177 ) );
  NOR2_X1 u2_u6_u4_U74 (.A2( u2_u6_X_28 ) , .A1( u2_u6_X_29 ) , .ZN( u2_u6_u4_n128 ) );
  NOR2_X1 u2_u6_u4_U75 (.A2( u2_u6_X_27 ) , .A1( u2_u6_X_30 ) , .ZN( u2_u6_u4_n102 ) );
  NOR2_X1 u2_u6_u4_U76 (.A2( u2_u6_X_25 ) , .A1( u2_u6_X_26 ) , .ZN( u2_u6_u4_n98 ) );
  AND2_X1 u2_u6_u4_U77 (.A2( u2_u6_X_25 ) , .A1( u2_u6_X_26 ) , .ZN( u2_u6_u4_n104 ) );
  AND2_X1 u2_u6_u4_U78 (.A1( u2_u6_X_30 ) , .A2( u2_u6_u4_n176 ) , .ZN( u2_u6_u4_n99 ) );
  AND2_X1 u2_u6_u4_U79 (.A1( u2_u6_X_26 ) , .ZN( u2_u6_u4_n101 ) , .A2( u2_u6_u4_n177 ) );
  AOI21_X1 u2_u6_u4_U8 (.ZN( u2_u6_u4_n109 ) , .A( u2_u6_u4_n153 ) , .B1( u2_u6_u4_n159 ) , .B2( u2_u6_u4_n184 ) );
  AND2_X1 u2_u6_u4_U80 (.A1( u2_u6_X_27 ) , .A2( u2_u6_X_30 ) , .ZN( u2_u6_u4_n103 ) );
  INV_X1 u2_u6_u4_U81 (.A( u2_u6_X_28 ) , .ZN( u2_u6_u4_n169 ) );
  INV_X1 u2_u6_u4_U82 (.A( u2_u6_X_29 ) , .ZN( u2_u6_u4_n168 ) );
  INV_X1 u2_u6_u4_U83 (.A( u2_u6_X_25 ) , .ZN( u2_u6_u4_n177 ) );
  INV_X1 u2_u6_u4_U84 (.A( u2_u6_X_27 ) , .ZN( u2_u6_u4_n176 ) );
  NAND4_X1 u2_u6_u4_U85 (.ZN( u2_out6_25 ) , .A4( u2_u6_u4_n139 ) , .A3( u2_u6_u4_n140 ) , .A2( u2_u6_u4_n141 ) , .A1( u2_u6_u4_n142 ) );
  OAI21_X1 u2_u6_u4_U86 (.B2( u2_u6_u4_n131 ) , .ZN( u2_u6_u4_n141 ) , .A( u2_u6_u4_n175 ) , .B1( u2_u6_u4_n183 ) );
  OAI21_X1 u2_u6_u4_U87 (.A( u2_u6_u4_n128 ) , .B2( u2_u6_u4_n129 ) , .B1( u2_u6_u4_n130 ) , .ZN( u2_u6_u4_n142 ) );
  NAND4_X1 u2_u6_u4_U88 (.ZN( u2_out6_14 ) , .A4( u2_u6_u4_n124 ) , .A3( u2_u6_u4_n125 ) , .A2( u2_u6_u4_n126 ) , .A1( u2_u6_u4_n127 ) );
  AOI22_X1 u2_u6_u4_U89 (.B2( u2_u6_u4_n117 ) , .ZN( u2_u6_u4_n126 ) , .A1( u2_u6_u4_n129 ) , .B1( u2_u6_u4_n152 ) , .A2( u2_u6_u4_n175 ) );
  AOI211_X1 u2_u6_u4_U9 (.B( u2_u6_u4_n136 ) , .A( u2_u6_u4_n137 ) , .C2( u2_u6_u4_n138 ) , .ZN( u2_u6_u4_n139 ) , .C1( u2_u6_u4_n182 ) );
  AOI22_X1 u2_u6_u4_U90 (.ZN( u2_u6_u4_n125 ) , .B2( u2_u6_u4_n131 ) , .A2( u2_u6_u4_n132 ) , .B1( u2_u6_u4_n138 ) , .A1( u2_u6_u4_n178 ) );
  NAND4_X1 u2_u6_u4_U91 (.ZN( u2_out6_8 ) , .A4( u2_u6_u4_n110 ) , .A3( u2_u6_u4_n111 ) , .A2( u2_u6_u4_n112 ) , .A1( u2_u6_u4_n186 ) );
  NAND2_X1 u2_u6_u4_U92 (.ZN( u2_u6_u4_n112 ) , .A2( u2_u6_u4_n130 ) , .A1( u2_u6_u4_n150 ) );
  AOI22_X1 u2_u6_u4_U93 (.ZN( u2_u6_u4_n111 ) , .B2( u2_u6_u4_n132 ) , .A1( u2_u6_u4_n152 ) , .B1( u2_u6_u4_n178 ) , .A2( u2_u6_u4_n97 ) );
  AOI22_X1 u2_u6_u4_U94 (.B2( u2_u6_u4_n149 ) , .B1( u2_u6_u4_n150 ) , .A2( u2_u6_u4_n151 ) , .A1( u2_u6_u4_n152 ) , .ZN( u2_u6_u4_n167 ) );
  NOR4_X1 u2_u6_u4_U95 (.A4( u2_u6_u4_n162 ) , .A3( u2_u6_u4_n163 ) , .A2( u2_u6_u4_n164 ) , .A1( u2_u6_u4_n165 ) , .ZN( u2_u6_u4_n166 ) );
  NAND3_X1 u2_u6_u4_U96 (.ZN( u2_out6_3 ) , .A3( u2_u6_u4_n166 ) , .A1( u2_u6_u4_n167 ) , .A2( u2_u6_u4_n186 ) );
  NAND3_X1 u2_u6_u4_U97 (.A3( u2_u6_u4_n146 ) , .A2( u2_u6_u4_n147 ) , .A1( u2_u6_u4_n148 ) , .ZN( u2_u6_u4_n149 ) );
  NAND3_X1 u2_u6_u4_U98 (.A3( u2_u6_u4_n143 ) , .A2( u2_u6_u4_n144 ) , .A1( u2_u6_u4_n145 ) , .ZN( u2_u6_u4_n151 ) );
  NAND3_X1 u2_u6_u4_U99 (.A3( u2_u6_u4_n121 ) , .ZN( u2_u6_u4_n122 ) , .A2( u2_u6_u4_n144 ) , .A1( u2_u6_u4_n154 ) );
  AOI21_X1 u2_u6_u6_U10 (.ZN( u2_u6_u6_n106 ) , .A( u2_u6_u6_n142 ) , .B2( u2_u6_u6_n159 ) , .B1( u2_u6_u6_n164 ) );
  INV_X1 u2_u6_u6_U11 (.A( u2_u6_u6_n155 ) , .ZN( u2_u6_u6_n161 ) );
  INV_X1 u2_u6_u6_U12 (.A( u2_u6_u6_n128 ) , .ZN( u2_u6_u6_n164 ) );
  NAND2_X1 u2_u6_u6_U13 (.ZN( u2_u6_u6_n110 ) , .A1( u2_u6_u6_n122 ) , .A2( u2_u6_u6_n129 ) );
  NAND2_X1 u2_u6_u6_U14 (.ZN( u2_u6_u6_n124 ) , .A2( u2_u6_u6_n146 ) , .A1( u2_u6_u6_n148 ) );
  INV_X1 u2_u6_u6_U15 (.A( u2_u6_u6_n132 ) , .ZN( u2_u6_u6_n171 ) );
  AND2_X1 u2_u6_u6_U16 (.A1( u2_u6_u6_n100 ) , .ZN( u2_u6_u6_n130 ) , .A2( u2_u6_u6_n147 ) );
  INV_X1 u2_u6_u6_U17 (.A( u2_u6_u6_n127 ) , .ZN( u2_u6_u6_n173 ) );
  INV_X1 u2_u6_u6_U18 (.A( u2_u6_u6_n121 ) , .ZN( u2_u6_u6_n167 ) );
  INV_X1 u2_u6_u6_U19 (.A( u2_u6_u6_n100 ) , .ZN( u2_u6_u6_n169 ) );
  INV_X1 u2_u6_u6_U20 (.A( u2_u6_u6_n123 ) , .ZN( u2_u6_u6_n170 ) );
  INV_X1 u2_u6_u6_U21 (.A( u2_u6_u6_n113 ) , .ZN( u2_u6_u6_n168 ) );
  AND2_X1 u2_u6_u6_U22 (.A1( u2_u6_u6_n107 ) , .A2( u2_u6_u6_n119 ) , .ZN( u2_u6_u6_n133 ) );
  AND2_X1 u2_u6_u6_U23 (.A2( u2_u6_u6_n121 ) , .A1( u2_u6_u6_n122 ) , .ZN( u2_u6_u6_n131 ) );
  AND3_X1 u2_u6_u6_U24 (.ZN( u2_u6_u6_n120 ) , .A2( u2_u6_u6_n127 ) , .A1( u2_u6_u6_n132 ) , .A3( u2_u6_u6_n145 ) );
  INV_X1 u2_u6_u6_U25 (.A( u2_u6_u6_n146 ) , .ZN( u2_u6_u6_n163 ) );
  AOI222_X1 u2_u6_u6_U26 (.ZN( u2_u6_u6_n114 ) , .A1( u2_u6_u6_n118 ) , .A2( u2_u6_u6_n126 ) , .B2( u2_u6_u6_n151 ) , .C2( u2_u6_u6_n159 ) , .C1( u2_u6_u6_n168 ) , .B1( u2_u6_u6_n169 ) );
  NOR2_X1 u2_u6_u6_U27 (.A1( u2_u6_u6_n162 ) , .A2( u2_u6_u6_n165 ) , .ZN( u2_u6_u6_n98 ) );
  AOI211_X1 u2_u6_u6_U28 (.B( u2_u6_u6_n149 ) , .A( u2_u6_u6_n150 ) , .C2( u2_u6_u6_n151 ) , .C1( u2_u6_u6_n152 ) , .ZN( u2_u6_u6_n153 ) );
  AOI21_X1 u2_u6_u6_U29 (.B2( u2_u6_u6_n147 ) , .B1( u2_u6_u6_n148 ) , .ZN( u2_u6_u6_n149 ) , .A( u2_u6_u6_n158 ) );
  INV_X1 u2_u6_u6_U3 (.A( u2_u6_u6_n110 ) , .ZN( u2_u6_u6_n166 ) );
  AOI21_X1 u2_u6_u6_U30 (.A( u2_u6_u6_n144 ) , .B2( u2_u6_u6_n145 ) , .B1( u2_u6_u6_n146 ) , .ZN( u2_u6_u6_n150 ) );
  NAND2_X1 u2_u6_u6_U31 (.A2( u2_u6_u6_n143 ) , .ZN( u2_u6_u6_n152 ) , .A1( u2_u6_u6_n166 ) );
  NAND2_X1 u2_u6_u6_U32 (.A1( u2_u6_u6_n144 ) , .ZN( u2_u6_u6_n151 ) , .A2( u2_u6_u6_n158 ) );
  NAND2_X1 u2_u6_u6_U33 (.ZN( u2_u6_u6_n132 ) , .A1( u2_u6_u6_n91 ) , .A2( u2_u6_u6_n97 ) );
  AOI22_X1 u2_u6_u6_U34 (.B2( u2_u6_u6_n110 ) , .B1( u2_u6_u6_n111 ) , .A1( u2_u6_u6_n112 ) , .ZN( u2_u6_u6_n115 ) , .A2( u2_u6_u6_n161 ) );
  NAND4_X1 u2_u6_u6_U35 (.A3( u2_u6_u6_n109 ) , .ZN( u2_u6_u6_n112 ) , .A4( u2_u6_u6_n132 ) , .A2( u2_u6_u6_n147 ) , .A1( u2_u6_u6_n166 ) );
  NOR2_X1 u2_u6_u6_U36 (.ZN( u2_u6_u6_n109 ) , .A1( u2_u6_u6_n170 ) , .A2( u2_u6_u6_n173 ) );
  NOR2_X1 u2_u6_u6_U37 (.A2( u2_u6_u6_n126 ) , .ZN( u2_u6_u6_n155 ) , .A1( u2_u6_u6_n160 ) );
  NAND2_X1 u2_u6_u6_U38 (.ZN( u2_u6_u6_n146 ) , .A2( u2_u6_u6_n94 ) , .A1( u2_u6_u6_n99 ) );
  AOI211_X1 u2_u6_u6_U39 (.B( u2_u6_u6_n134 ) , .A( u2_u6_u6_n135 ) , .C1( u2_u6_u6_n136 ) , .ZN( u2_u6_u6_n137 ) , .C2( u2_u6_u6_n151 ) );
  AOI22_X1 u2_u6_u6_U4 (.B2( u2_u6_u6_n101 ) , .A1( u2_u6_u6_n102 ) , .ZN( u2_u6_u6_n103 ) , .B1( u2_u6_u6_n160 ) , .A2( u2_u6_u6_n161 ) );
  NAND4_X1 u2_u6_u6_U40 (.A4( u2_u6_u6_n127 ) , .A3( u2_u6_u6_n128 ) , .A2( u2_u6_u6_n129 ) , .A1( u2_u6_u6_n130 ) , .ZN( u2_u6_u6_n136 ) );
  AOI21_X1 u2_u6_u6_U41 (.B2( u2_u6_u6_n132 ) , .B1( u2_u6_u6_n133 ) , .ZN( u2_u6_u6_n134 ) , .A( u2_u6_u6_n158 ) );
  AOI21_X1 u2_u6_u6_U42 (.B1( u2_u6_u6_n131 ) , .ZN( u2_u6_u6_n135 ) , .A( u2_u6_u6_n144 ) , .B2( u2_u6_u6_n146 ) );
  INV_X1 u2_u6_u6_U43 (.A( u2_u6_u6_n111 ) , .ZN( u2_u6_u6_n158 ) );
  NAND2_X1 u2_u6_u6_U44 (.ZN( u2_u6_u6_n127 ) , .A1( u2_u6_u6_n91 ) , .A2( u2_u6_u6_n92 ) );
  NAND2_X1 u2_u6_u6_U45 (.ZN( u2_u6_u6_n129 ) , .A2( u2_u6_u6_n95 ) , .A1( u2_u6_u6_n96 ) );
  INV_X1 u2_u6_u6_U46 (.A( u2_u6_u6_n144 ) , .ZN( u2_u6_u6_n159 ) );
  NAND2_X1 u2_u6_u6_U47 (.ZN( u2_u6_u6_n145 ) , .A2( u2_u6_u6_n97 ) , .A1( u2_u6_u6_n98 ) );
  NAND2_X1 u2_u6_u6_U48 (.ZN( u2_u6_u6_n148 ) , .A2( u2_u6_u6_n92 ) , .A1( u2_u6_u6_n94 ) );
  NAND2_X1 u2_u6_u6_U49 (.ZN( u2_u6_u6_n108 ) , .A2( u2_u6_u6_n139 ) , .A1( u2_u6_u6_n144 ) );
  NOR2_X1 u2_u6_u6_U5 (.A1( u2_u6_u6_n118 ) , .ZN( u2_u6_u6_n143 ) , .A2( u2_u6_u6_n168 ) );
  NAND2_X1 u2_u6_u6_U50 (.ZN( u2_u6_u6_n121 ) , .A2( u2_u6_u6_n95 ) , .A1( u2_u6_u6_n97 ) );
  NAND2_X1 u2_u6_u6_U51 (.ZN( u2_u6_u6_n107 ) , .A2( u2_u6_u6_n92 ) , .A1( u2_u6_u6_n95 ) );
  AND2_X1 u2_u6_u6_U52 (.ZN( u2_u6_u6_n118 ) , .A2( u2_u6_u6_n91 ) , .A1( u2_u6_u6_n99 ) );
  NAND2_X1 u2_u6_u6_U53 (.ZN( u2_u6_u6_n147 ) , .A2( u2_u6_u6_n98 ) , .A1( u2_u6_u6_n99 ) );
  NAND2_X1 u2_u6_u6_U54 (.ZN( u2_u6_u6_n128 ) , .A1( u2_u6_u6_n94 ) , .A2( u2_u6_u6_n96 ) );
  NAND2_X1 u2_u6_u6_U55 (.ZN( u2_u6_u6_n119 ) , .A2( u2_u6_u6_n95 ) , .A1( u2_u6_u6_n99 ) );
  NAND2_X1 u2_u6_u6_U56 (.ZN( u2_u6_u6_n123 ) , .A2( u2_u6_u6_n91 ) , .A1( u2_u6_u6_n96 ) );
  NAND2_X1 u2_u6_u6_U57 (.ZN( u2_u6_u6_n100 ) , .A2( u2_u6_u6_n92 ) , .A1( u2_u6_u6_n98 ) );
  NAND2_X1 u2_u6_u6_U58 (.ZN( u2_u6_u6_n122 ) , .A1( u2_u6_u6_n94 ) , .A2( u2_u6_u6_n97 ) );
  INV_X1 u2_u6_u6_U59 (.A( u2_u6_u6_n139 ) , .ZN( u2_u6_u6_n160 ) );
  AOI21_X1 u2_u6_u6_U6 (.B1( u2_u6_u6_n107 ) , .B2( u2_u6_u6_n132 ) , .A( u2_u6_u6_n158 ) , .ZN( u2_u6_u6_n88 ) );
  NAND2_X1 u2_u6_u6_U60 (.ZN( u2_u6_u6_n113 ) , .A1( u2_u6_u6_n96 ) , .A2( u2_u6_u6_n98 ) );
  NOR2_X1 u2_u6_u6_U61 (.A2( u2_u6_X_40 ) , .A1( u2_u6_X_41 ) , .ZN( u2_u6_u6_n126 ) );
  NOR2_X1 u2_u6_u6_U62 (.A2( u2_u6_X_39 ) , .A1( u2_u6_X_42 ) , .ZN( u2_u6_u6_n92 ) );
  NOR2_X1 u2_u6_u6_U63 (.A2( u2_u6_X_39 ) , .A1( u2_u6_u6_n156 ) , .ZN( u2_u6_u6_n97 ) );
  NOR2_X1 u2_u6_u6_U64 (.A2( u2_u6_X_38 ) , .A1( u2_u6_u6_n165 ) , .ZN( u2_u6_u6_n95 ) );
  NOR2_X1 u2_u6_u6_U65 (.A2( u2_u6_X_41 ) , .ZN( u2_u6_u6_n111 ) , .A1( u2_u6_u6_n157 ) );
  NOR2_X1 u2_u6_u6_U66 (.A2( u2_u6_X_37 ) , .A1( u2_u6_u6_n162 ) , .ZN( u2_u6_u6_n94 ) );
  NOR2_X1 u2_u6_u6_U67 (.A2( u2_u6_X_37 ) , .A1( u2_u6_X_38 ) , .ZN( u2_u6_u6_n91 ) );
  NAND2_X1 u2_u6_u6_U68 (.A1( u2_u6_X_41 ) , .ZN( u2_u6_u6_n144 ) , .A2( u2_u6_u6_n157 ) );
  NAND2_X1 u2_u6_u6_U69 (.A2( u2_u6_X_40 ) , .A1( u2_u6_X_41 ) , .ZN( u2_u6_u6_n139 ) );
  OAI21_X1 u2_u6_u6_U7 (.A( u2_u6_u6_n159 ) , .B1( u2_u6_u6_n169 ) , .B2( u2_u6_u6_n173 ) , .ZN( u2_u6_u6_n90 ) );
  AND2_X1 u2_u6_u6_U70 (.A1( u2_u6_X_39 ) , .A2( u2_u6_u6_n156 ) , .ZN( u2_u6_u6_n96 ) );
  AND2_X1 u2_u6_u6_U71 (.A1( u2_u6_X_39 ) , .A2( u2_u6_X_42 ) , .ZN( u2_u6_u6_n99 ) );
  INV_X1 u2_u6_u6_U72 (.A( u2_u6_X_40 ) , .ZN( u2_u6_u6_n157 ) );
  INV_X1 u2_u6_u6_U73 (.A( u2_u6_X_37 ) , .ZN( u2_u6_u6_n165 ) );
  INV_X1 u2_u6_u6_U74 (.A( u2_u6_X_38 ) , .ZN( u2_u6_u6_n162 ) );
  INV_X1 u2_u6_u6_U75 (.A( u2_u6_X_42 ) , .ZN( u2_u6_u6_n156 ) );
  NAND4_X1 u2_u6_u6_U76 (.ZN( u2_out6_32 ) , .A4( u2_u6_u6_n103 ) , .A3( u2_u6_u6_n104 ) , .A2( u2_u6_u6_n105 ) , .A1( u2_u6_u6_n106 ) );
  AOI22_X1 u2_u6_u6_U77 (.ZN( u2_u6_u6_n104 ) , .A1( u2_u6_u6_n111 ) , .B1( u2_u6_u6_n124 ) , .B2( u2_u6_u6_n151 ) , .A2( u2_u6_u6_n93 ) );
  AOI22_X1 u2_u6_u6_U78 (.ZN( u2_u6_u6_n105 ) , .A2( u2_u6_u6_n108 ) , .A1( u2_u6_u6_n118 ) , .B2( u2_u6_u6_n126 ) , .B1( u2_u6_u6_n171 ) );
  NAND4_X1 u2_u6_u6_U79 (.ZN( u2_out6_12 ) , .A4( u2_u6_u6_n114 ) , .A3( u2_u6_u6_n115 ) , .A2( u2_u6_u6_n116 ) , .A1( u2_u6_u6_n117 ) );
  INV_X1 u2_u6_u6_U8 (.ZN( u2_u6_u6_n172 ) , .A( u2_u6_u6_n88 ) );
  OAI22_X1 u2_u6_u6_U80 (.B2( u2_u6_u6_n111 ) , .ZN( u2_u6_u6_n116 ) , .B1( u2_u6_u6_n126 ) , .A2( u2_u6_u6_n164 ) , .A1( u2_u6_u6_n167 ) );
  OAI21_X1 u2_u6_u6_U81 (.A( u2_u6_u6_n108 ) , .ZN( u2_u6_u6_n117 ) , .B2( u2_u6_u6_n141 ) , .B1( u2_u6_u6_n163 ) );
  OAI211_X1 u2_u6_u6_U82 (.ZN( u2_out6_22 ) , .B( u2_u6_u6_n137 ) , .A( u2_u6_u6_n138 ) , .C2( u2_u6_u6_n139 ) , .C1( u2_u6_u6_n140 ) );
  AOI22_X1 u2_u6_u6_U83 (.B1( u2_u6_u6_n124 ) , .A2( u2_u6_u6_n125 ) , .A1( u2_u6_u6_n126 ) , .ZN( u2_u6_u6_n138 ) , .B2( u2_u6_u6_n161 ) );
  AND4_X1 u2_u6_u6_U84 (.A3( u2_u6_u6_n119 ) , .A1( u2_u6_u6_n120 ) , .A4( u2_u6_u6_n129 ) , .ZN( u2_u6_u6_n140 ) , .A2( u2_u6_u6_n143 ) );
  OAI211_X1 u2_u6_u6_U85 (.ZN( u2_out6_7 ) , .B( u2_u6_u6_n153 ) , .C2( u2_u6_u6_n154 ) , .C1( u2_u6_u6_n155 ) , .A( u2_u6_u6_n174 ) );
  NOR3_X1 u2_u6_u6_U86 (.A1( u2_u6_u6_n141 ) , .ZN( u2_u6_u6_n154 ) , .A3( u2_u6_u6_n164 ) , .A2( u2_u6_u6_n171 ) );
  INV_X1 u2_u6_u6_U87 (.A( u2_u6_u6_n142 ) , .ZN( u2_u6_u6_n174 ) );
  NAND3_X1 u2_u6_u6_U88 (.A2( u2_u6_u6_n123 ) , .ZN( u2_u6_u6_n125 ) , .A1( u2_u6_u6_n130 ) , .A3( u2_u6_u6_n131 ) );
  NAND3_X1 u2_u6_u6_U89 (.A3( u2_u6_u6_n133 ) , .ZN( u2_u6_u6_n141 ) , .A1( u2_u6_u6_n145 ) , .A2( u2_u6_u6_n148 ) );
  AOI22_X1 u2_u6_u6_U9 (.A2( u2_u6_u6_n151 ) , .B2( u2_u6_u6_n161 ) , .A1( u2_u6_u6_n167 ) , .B1( u2_u6_u6_n170 ) , .ZN( u2_u6_u6_n89 ) );
  NAND3_X1 u2_u6_u6_U90 (.ZN( u2_u6_u6_n101 ) , .A3( u2_u6_u6_n107 ) , .A2( u2_u6_u6_n121 ) , .A1( u2_u6_u6_n127 ) );
  NAND3_X1 u2_u6_u6_U91 (.ZN( u2_u6_u6_n102 ) , .A3( u2_u6_u6_n130 ) , .A2( u2_u6_u6_n145 ) , .A1( u2_u6_u6_n166 ) );
  NAND3_X1 u2_u6_u6_U92 (.A3( u2_u6_u6_n113 ) , .A1( u2_u6_u6_n119 ) , .A2( u2_u6_u6_n123 ) , .ZN( u2_u6_u6_n93 ) );
  NAND3_X1 u2_u6_u6_U93 (.ZN( u2_u6_u6_n142 ) , .A2( u2_u6_u6_n172 ) , .A3( u2_u6_u6_n89 ) , .A1( u2_u6_u6_n90 ) );
  AND3_X1 u2_u6_u7_U10 (.A3( u2_u6_u7_n110 ) , .A2( u2_u6_u7_n127 ) , .A1( u2_u6_u7_n132 ) , .ZN( u2_u6_u7_n92 ) );
  OAI21_X1 u2_u6_u7_U11 (.A( u2_u6_u7_n161 ) , .B1( u2_u6_u7_n168 ) , .B2( u2_u6_u7_n173 ) , .ZN( u2_u6_u7_n91 ) );
  AOI211_X1 u2_u6_u7_U12 (.A( u2_u6_u7_n117 ) , .ZN( u2_u6_u7_n118 ) , .C2( u2_u6_u7_n126 ) , .C1( u2_u6_u7_n177 ) , .B( u2_u6_u7_n180 ) );
  OAI22_X1 u2_u6_u7_U13 (.B1( u2_u6_u7_n115 ) , .ZN( u2_u6_u7_n117 ) , .A2( u2_u6_u7_n133 ) , .A1( u2_u6_u7_n137 ) , .B2( u2_u6_u7_n162 ) );
  INV_X1 u2_u6_u7_U14 (.A( u2_u6_u7_n116 ) , .ZN( u2_u6_u7_n180 ) );
  NOR3_X1 u2_u6_u7_U15 (.ZN( u2_u6_u7_n115 ) , .A3( u2_u6_u7_n145 ) , .A2( u2_u6_u7_n168 ) , .A1( u2_u6_u7_n169 ) );
  OAI211_X1 u2_u6_u7_U16 (.B( u2_u6_u7_n122 ) , .A( u2_u6_u7_n123 ) , .C2( u2_u6_u7_n124 ) , .ZN( u2_u6_u7_n154 ) , .C1( u2_u6_u7_n162 ) );
  AOI222_X1 u2_u6_u7_U17 (.ZN( u2_u6_u7_n122 ) , .C2( u2_u6_u7_n126 ) , .C1( u2_u6_u7_n145 ) , .B1( u2_u6_u7_n161 ) , .A2( u2_u6_u7_n165 ) , .B2( u2_u6_u7_n170 ) , .A1( u2_u6_u7_n176 ) );
  INV_X1 u2_u6_u7_U18 (.A( u2_u6_u7_n133 ) , .ZN( u2_u6_u7_n176 ) );
  NOR3_X1 u2_u6_u7_U19 (.A2( u2_u6_u7_n134 ) , .A1( u2_u6_u7_n135 ) , .ZN( u2_u6_u7_n136 ) , .A3( u2_u6_u7_n171 ) );
  NOR2_X1 u2_u6_u7_U20 (.A1( u2_u6_u7_n130 ) , .A2( u2_u6_u7_n134 ) , .ZN( u2_u6_u7_n153 ) );
  INV_X1 u2_u6_u7_U21 (.A( u2_u6_u7_n101 ) , .ZN( u2_u6_u7_n165 ) );
  NOR2_X1 u2_u6_u7_U22 (.ZN( u2_u6_u7_n111 ) , .A2( u2_u6_u7_n134 ) , .A1( u2_u6_u7_n169 ) );
  AOI21_X1 u2_u6_u7_U23 (.ZN( u2_u6_u7_n104 ) , .B2( u2_u6_u7_n112 ) , .B1( u2_u6_u7_n127 ) , .A( u2_u6_u7_n164 ) );
  AOI21_X1 u2_u6_u7_U24 (.ZN( u2_u6_u7_n106 ) , .B1( u2_u6_u7_n133 ) , .B2( u2_u6_u7_n146 ) , .A( u2_u6_u7_n162 ) );
  AOI21_X1 u2_u6_u7_U25 (.A( u2_u6_u7_n101 ) , .ZN( u2_u6_u7_n107 ) , .B2( u2_u6_u7_n128 ) , .B1( u2_u6_u7_n175 ) );
  INV_X1 u2_u6_u7_U26 (.A( u2_u6_u7_n138 ) , .ZN( u2_u6_u7_n171 ) );
  INV_X1 u2_u6_u7_U27 (.A( u2_u6_u7_n131 ) , .ZN( u2_u6_u7_n177 ) );
  INV_X1 u2_u6_u7_U28 (.A( u2_u6_u7_n110 ) , .ZN( u2_u6_u7_n174 ) );
  NAND2_X1 u2_u6_u7_U29 (.A1( u2_u6_u7_n129 ) , .A2( u2_u6_u7_n132 ) , .ZN( u2_u6_u7_n149 ) );
  OAI21_X1 u2_u6_u7_U3 (.ZN( u2_u6_u7_n159 ) , .A( u2_u6_u7_n165 ) , .B2( u2_u6_u7_n171 ) , .B1( u2_u6_u7_n174 ) );
  NAND2_X1 u2_u6_u7_U30 (.A1( u2_u6_u7_n113 ) , .A2( u2_u6_u7_n124 ) , .ZN( u2_u6_u7_n130 ) );
  INV_X1 u2_u6_u7_U31 (.A( u2_u6_u7_n112 ) , .ZN( u2_u6_u7_n173 ) );
  INV_X1 u2_u6_u7_U32 (.A( u2_u6_u7_n128 ) , .ZN( u2_u6_u7_n168 ) );
  INV_X1 u2_u6_u7_U33 (.A( u2_u6_u7_n148 ) , .ZN( u2_u6_u7_n169 ) );
  INV_X1 u2_u6_u7_U34 (.A( u2_u6_u7_n127 ) , .ZN( u2_u6_u7_n179 ) );
  NOR2_X1 u2_u6_u7_U35 (.ZN( u2_u6_u7_n101 ) , .A2( u2_u6_u7_n150 ) , .A1( u2_u6_u7_n156 ) );
  AOI211_X1 u2_u6_u7_U36 (.B( u2_u6_u7_n154 ) , .A( u2_u6_u7_n155 ) , .C1( u2_u6_u7_n156 ) , .ZN( u2_u6_u7_n157 ) , .C2( u2_u6_u7_n172 ) );
  INV_X1 u2_u6_u7_U37 (.A( u2_u6_u7_n153 ) , .ZN( u2_u6_u7_n172 ) );
  AOI211_X1 u2_u6_u7_U38 (.B( u2_u6_u7_n139 ) , .A( u2_u6_u7_n140 ) , .C2( u2_u6_u7_n141 ) , .ZN( u2_u6_u7_n142 ) , .C1( u2_u6_u7_n156 ) );
  NAND4_X1 u2_u6_u7_U39 (.A3( u2_u6_u7_n127 ) , .A2( u2_u6_u7_n128 ) , .A1( u2_u6_u7_n129 ) , .ZN( u2_u6_u7_n141 ) , .A4( u2_u6_u7_n147 ) );
  INV_X1 u2_u6_u7_U4 (.A( u2_u6_u7_n111 ) , .ZN( u2_u6_u7_n170 ) );
  AOI21_X1 u2_u6_u7_U40 (.A( u2_u6_u7_n137 ) , .B1( u2_u6_u7_n138 ) , .ZN( u2_u6_u7_n139 ) , .B2( u2_u6_u7_n146 ) );
  OAI22_X1 u2_u6_u7_U41 (.B1( u2_u6_u7_n136 ) , .ZN( u2_u6_u7_n140 ) , .A1( u2_u6_u7_n153 ) , .B2( u2_u6_u7_n162 ) , .A2( u2_u6_u7_n164 ) );
  AOI21_X1 u2_u6_u7_U42 (.ZN( u2_u6_u7_n123 ) , .B1( u2_u6_u7_n165 ) , .B2( u2_u6_u7_n177 ) , .A( u2_u6_u7_n97 ) );
  AOI21_X1 u2_u6_u7_U43 (.B2( u2_u6_u7_n113 ) , .B1( u2_u6_u7_n124 ) , .A( u2_u6_u7_n125 ) , .ZN( u2_u6_u7_n97 ) );
  INV_X1 u2_u6_u7_U44 (.A( u2_u6_u7_n125 ) , .ZN( u2_u6_u7_n161 ) );
  INV_X1 u2_u6_u7_U45 (.A( u2_u6_u7_n152 ) , .ZN( u2_u6_u7_n162 ) );
  AOI22_X1 u2_u6_u7_U46 (.A2( u2_u6_u7_n114 ) , .ZN( u2_u6_u7_n119 ) , .B1( u2_u6_u7_n130 ) , .A1( u2_u6_u7_n156 ) , .B2( u2_u6_u7_n165 ) );
  NAND2_X1 u2_u6_u7_U47 (.A2( u2_u6_u7_n112 ) , .ZN( u2_u6_u7_n114 ) , .A1( u2_u6_u7_n175 ) );
  AND2_X1 u2_u6_u7_U48 (.ZN( u2_u6_u7_n145 ) , .A2( u2_u6_u7_n98 ) , .A1( u2_u6_u7_n99 ) );
  NOR2_X1 u2_u6_u7_U49 (.ZN( u2_u6_u7_n137 ) , .A1( u2_u6_u7_n150 ) , .A2( u2_u6_u7_n161 ) );
  INV_X1 u2_u6_u7_U5 (.A( u2_u6_u7_n149 ) , .ZN( u2_u6_u7_n175 ) );
  AOI21_X1 u2_u6_u7_U50 (.ZN( u2_u6_u7_n105 ) , .B2( u2_u6_u7_n110 ) , .A( u2_u6_u7_n125 ) , .B1( u2_u6_u7_n147 ) );
  NAND2_X1 u2_u6_u7_U51 (.ZN( u2_u6_u7_n146 ) , .A1( u2_u6_u7_n95 ) , .A2( u2_u6_u7_n98 ) );
  NAND2_X1 u2_u6_u7_U52 (.A2( u2_u6_u7_n103 ) , .ZN( u2_u6_u7_n147 ) , .A1( u2_u6_u7_n93 ) );
  NAND2_X1 u2_u6_u7_U53 (.A1( u2_u6_u7_n103 ) , .ZN( u2_u6_u7_n127 ) , .A2( u2_u6_u7_n99 ) );
  OR2_X1 u2_u6_u7_U54 (.ZN( u2_u6_u7_n126 ) , .A2( u2_u6_u7_n152 ) , .A1( u2_u6_u7_n156 ) );
  NAND2_X1 u2_u6_u7_U55 (.A2( u2_u6_u7_n102 ) , .A1( u2_u6_u7_n103 ) , .ZN( u2_u6_u7_n133 ) );
  NAND2_X1 u2_u6_u7_U56 (.ZN( u2_u6_u7_n112 ) , .A2( u2_u6_u7_n96 ) , .A1( u2_u6_u7_n99 ) );
  NAND2_X1 u2_u6_u7_U57 (.A2( u2_u6_u7_n102 ) , .ZN( u2_u6_u7_n128 ) , .A1( u2_u6_u7_n98 ) );
  NAND2_X1 u2_u6_u7_U58 (.A1( u2_u6_u7_n100 ) , .ZN( u2_u6_u7_n113 ) , .A2( u2_u6_u7_n93 ) );
  NAND2_X1 u2_u6_u7_U59 (.A2( u2_u6_u7_n102 ) , .ZN( u2_u6_u7_n124 ) , .A1( u2_u6_u7_n96 ) );
  INV_X1 u2_u6_u7_U6 (.A( u2_u6_u7_n154 ) , .ZN( u2_u6_u7_n178 ) );
  NAND2_X1 u2_u6_u7_U60 (.ZN( u2_u6_u7_n110 ) , .A1( u2_u6_u7_n95 ) , .A2( u2_u6_u7_n96 ) );
  INV_X1 u2_u6_u7_U61 (.A( u2_u6_u7_n150 ) , .ZN( u2_u6_u7_n164 ) );
  AND2_X1 u2_u6_u7_U62 (.ZN( u2_u6_u7_n134 ) , .A1( u2_u6_u7_n93 ) , .A2( u2_u6_u7_n98 ) );
  NAND2_X1 u2_u6_u7_U63 (.A1( u2_u6_u7_n100 ) , .A2( u2_u6_u7_n102 ) , .ZN( u2_u6_u7_n129 ) );
  NAND2_X1 u2_u6_u7_U64 (.A2( u2_u6_u7_n103 ) , .ZN( u2_u6_u7_n131 ) , .A1( u2_u6_u7_n95 ) );
  NAND2_X1 u2_u6_u7_U65 (.A1( u2_u6_u7_n100 ) , .ZN( u2_u6_u7_n138 ) , .A2( u2_u6_u7_n99 ) );
  NAND2_X1 u2_u6_u7_U66 (.ZN( u2_u6_u7_n132 ) , .A1( u2_u6_u7_n93 ) , .A2( u2_u6_u7_n96 ) );
  NAND2_X1 u2_u6_u7_U67 (.A1( u2_u6_u7_n100 ) , .ZN( u2_u6_u7_n148 ) , .A2( u2_u6_u7_n95 ) );
  NOR2_X1 u2_u6_u7_U68 (.A2( u2_u6_X_47 ) , .ZN( u2_u6_u7_n150 ) , .A1( u2_u6_u7_n163 ) );
  NOR2_X1 u2_u6_u7_U69 (.A2( u2_u6_X_43 ) , .A1( u2_u6_X_44 ) , .ZN( u2_u6_u7_n103 ) );
  AOI211_X1 u2_u6_u7_U7 (.ZN( u2_u6_u7_n116 ) , .A( u2_u6_u7_n155 ) , .C1( u2_u6_u7_n161 ) , .C2( u2_u6_u7_n171 ) , .B( u2_u6_u7_n94 ) );
  NOR2_X1 u2_u6_u7_U70 (.A2( u2_u6_X_48 ) , .A1( u2_u6_u7_n166 ) , .ZN( u2_u6_u7_n95 ) );
  NOR2_X1 u2_u6_u7_U71 (.A2( u2_u6_X_45 ) , .A1( u2_u6_X_48 ) , .ZN( u2_u6_u7_n99 ) );
  NOR2_X1 u2_u6_u7_U72 (.A2( u2_u6_X_44 ) , .A1( u2_u6_u7_n167 ) , .ZN( u2_u6_u7_n98 ) );
  NOR2_X1 u2_u6_u7_U73 (.A2( u2_u6_X_46 ) , .A1( u2_u6_X_47 ) , .ZN( u2_u6_u7_n152 ) );
  AND2_X1 u2_u6_u7_U74 (.A1( u2_u6_X_47 ) , .ZN( u2_u6_u7_n156 ) , .A2( u2_u6_u7_n163 ) );
  NAND2_X1 u2_u6_u7_U75 (.A2( u2_u6_X_46 ) , .A1( u2_u6_X_47 ) , .ZN( u2_u6_u7_n125 ) );
  AND2_X1 u2_u6_u7_U76 (.A2( u2_u6_X_45 ) , .A1( u2_u6_X_48 ) , .ZN( u2_u6_u7_n102 ) );
  AND2_X1 u2_u6_u7_U77 (.A2( u2_u6_X_43 ) , .A1( u2_u6_X_44 ) , .ZN( u2_u6_u7_n96 ) );
  AND2_X1 u2_u6_u7_U78 (.A1( u2_u6_X_44 ) , .ZN( u2_u6_u7_n100 ) , .A2( u2_u6_u7_n167 ) );
  AND2_X1 u2_u6_u7_U79 (.A1( u2_u6_X_48 ) , .A2( u2_u6_u7_n166 ) , .ZN( u2_u6_u7_n93 ) );
  OAI222_X1 u2_u6_u7_U8 (.C2( u2_u6_u7_n101 ) , .B2( u2_u6_u7_n111 ) , .A1( u2_u6_u7_n113 ) , .C1( u2_u6_u7_n146 ) , .A2( u2_u6_u7_n162 ) , .B1( u2_u6_u7_n164 ) , .ZN( u2_u6_u7_n94 ) );
  INV_X1 u2_u6_u7_U80 (.A( u2_u6_X_46 ) , .ZN( u2_u6_u7_n163 ) );
  INV_X1 u2_u6_u7_U81 (.A( u2_u6_X_43 ) , .ZN( u2_u6_u7_n167 ) );
  INV_X1 u2_u6_u7_U82 (.A( u2_u6_X_45 ) , .ZN( u2_u6_u7_n166 ) );
  NAND4_X1 u2_u6_u7_U83 (.ZN( u2_out6_5 ) , .A4( u2_u6_u7_n108 ) , .A3( u2_u6_u7_n109 ) , .A1( u2_u6_u7_n116 ) , .A2( u2_u6_u7_n123 ) );
  AOI22_X1 u2_u6_u7_U84 (.ZN( u2_u6_u7_n109 ) , .A2( u2_u6_u7_n126 ) , .B2( u2_u6_u7_n145 ) , .B1( u2_u6_u7_n156 ) , .A1( u2_u6_u7_n171 ) );
  NOR4_X1 u2_u6_u7_U85 (.A4( u2_u6_u7_n104 ) , .A3( u2_u6_u7_n105 ) , .A2( u2_u6_u7_n106 ) , .A1( u2_u6_u7_n107 ) , .ZN( u2_u6_u7_n108 ) );
  NAND4_X1 u2_u6_u7_U86 (.ZN( u2_out6_27 ) , .A4( u2_u6_u7_n118 ) , .A3( u2_u6_u7_n119 ) , .A2( u2_u6_u7_n120 ) , .A1( u2_u6_u7_n121 ) );
  OAI21_X1 u2_u6_u7_U87 (.ZN( u2_u6_u7_n121 ) , .B2( u2_u6_u7_n145 ) , .A( u2_u6_u7_n150 ) , .B1( u2_u6_u7_n174 ) );
  OAI21_X1 u2_u6_u7_U88 (.ZN( u2_u6_u7_n120 ) , .A( u2_u6_u7_n161 ) , .B2( u2_u6_u7_n170 ) , .B1( u2_u6_u7_n179 ) );
  NAND4_X1 u2_u6_u7_U89 (.ZN( u2_out6_21 ) , .A4( u2_u6_u7_n157 ) , .A3( u2_u6_u7_n158 ) , .A2( u2_u6_u7_n159 ) , .A1( u2_u6_u7_n160 ) );
  OAI221_X1 u2_u6_u7_U9 (.C1( u2_u6_u7_n101 ) , .C2( u2_u6_u7_n147 ) , .ZN( u2_u6_u7_n155 ) , .B2( u2_u6_u7_n162 ) , .A( u2_u6_u7_n91 ) , .B1( u2_u6_u7_n92 ) );
  OAI21_X1 u2_u6_u7_U90 (.B1( u2_u6_u7_n145 ) , .ZN( u2_u6_u7_n160 ) , .A( u2_u6_u7_n161 ) , .B2( u2_u6_u7_n177 ) );
  AOI22_X1 u2_u6_u7_U91 (.B2( u2_u6_u7_n149 ) , .B1( u2_u6_u7_n150 ) , .A2( u2_u6_u7_n151 ) , .A1( u2_u6_u7_n152 ) , .ZN( u2_u6_u7_n158 ) );
  NAND4_X1 u2_u6_u7_U92 (.ZN( u2_out6_15 ) , .A4( u2_u6_u7_n142 ) , .A3( u2_u6_u7_n143 ) , .A2( u2_u6_u7_n144 ) , .A1( u2_u6_u7_n178 ) );
  OR2_X1 u2_u6_u7_U93 (.A2( u2_u6_u7_n125 ) , .A1( u2_u6_u7_n129 ) , .ZN( u2_u6_u7_n144 ) );
  AOI22_X1 u2_u6_u7_U94 (.A2( u2_u6_u7_n126 ) , .ZN( u2_u6_u7_n143 ) , .B2( u2_u6_u7_n165 ) , .B1( u2_u6_u7_n173 ) , .A1( u2_u6_u7_n174 ) );
  NAND3_X1 u2_u6_u7_U95 (.A3( u2_u6_u7_n146 ) , .A2( u2_u6_u7_n147 ) , .A1( u2_u6_u7_n148 ) , .ZN( u2_u6_u7_n151 ) );
  NAND3_X1 u2_u6_u7_U96 (.A3( u2_u6_u7_n131 ) , .A2( u2_u6_u7_n132 ) , .A1( u2_u6_u7_n133 ) , .ZN( u2_u6_u7_n135 ) );
  XOR2_X1 u2_u7_U10 (.B( u2_K8_45 ) , .A( u2_R6_30 ) , .Z( u2_u7_X_45 ) );
  XOR2_X1 u2_u7_U11 (.B( u2_K8_44 ) , .A( u2_R6_29 ) , .Z( u2_u7_X_44 ) );
  XOR2_X1 u2_u7_U12 (.B( u2_K8_43 ) , .A( u2_R6_28 ) , .Z( u2_u7_X_43 ) );
  XOR2_X1 u2_u7_U13 (.B( u2_K8_42 ) , .A( u2_R6_29 ) , .Z( u2_u7_X_42 ) );
  XOR2_X1 u2_u7_U14 (.B( u2_K8_41 ) , .A( u2_R6_28 ) , .Z( u2_u7_X_41 ) );
  XOR2_X1 u2_u7_U15 (.B( u2_K8_40 ) , .A( u2_R6_27 ) , .Z( u2_u7_X_40 ) );
  XOR2_X1 u2_u7_U17 (.B( u2_K8_39 ) , .A( u2_R6_26 ) , .Z( u2_u7_X_39 ) );
  XOR2_X1 u2_u7_U18 (.B( u2_K8_38 ) , .A( u2_R6_25 ) , .Z( u2_u7_X_38 ) );
  XOR2_X1 u2_u7_U19 (.B( u2_K8_37 ) , .A( u2_R6_24 ) , .Z( u2_u7_X_37 ) );
  XOR2_X1 u2_u7_U7 (.B( u2_K8_48 ) , .A( u2_R6_1 ) , .Z( u2_u7_X_48 ) );
  XOR2_X1 u2_u7_U8 (.B( u2_K8_47 ) , .A( u2_R6_32 ) , .Z( u2_u7_X_47 ) );
  XOR2_X1 u2_u7_U9 (.B( u2_K8_46 ) , .A( u2_R6_31 ) , .Z( u2_u7_X_46 ) );
  INV_X1 u2_u7_u6_U10 (.ZN( u2_u7_u6_n172 ) , .A( u2_u7_u6_n88 ) );
  OAI21_X1 u2_u7_u6_U11 (.A( u2_u7_u6_n159 ) , .B1( u2_u7_u6_n169 ) , .B2( u2_u7_u6_n173 ) , .ZN( u2_u7_u6_n90 ) );
  AOI22_X1 u2_u7_u6_U12 (.A2( u2_u7_u6_n151 ) , .B2( u2_u7_u6_n161 ) , .A1( u2_u7_u6_n167 ) , .B1( u2_u7_u6_n170 ) , .ZN( u2_u7_u6_n89 ) );
  AOI21_X1 u2_u7_u6_U13 (.ZN( u2_u7_u6_n106 ) , .A( u2_u7_u6_n142 ) , .B2( u2_u7_u6_n159 ) , .B1( u2_u7_u6_n164 ) );
  INV_X1 u2_u7_u6_U14 (.A( u2_u7_u6_n155 ) , .ZN( u2_u7_u6_n161 ) );
  INV_X1 u2_u7_u6_U15 (.A( u2_u7_u6_n128 ) , .ZN( u2_u7_u6_n164 ) );
  NAND2_X1 u2_u7_u6_U16 (.ZN( u2_u7_u6_n110 ) , .A1( u2_u7_u6_n122 ) , .A2( u2_u7_u6_n129 ) );
  NAND2_X1 u2_u7_u6_U17 (.ZN( u2_u7_u6_n124 ) , .A2( u2_u7_u6_n146 ) , .A1( u2_u7_u6_n148 ) );
  INV_X1 u2_u7_u6_U18 (.A( u2_u7_u6_n132 ) , .ZN( u2_u7_u6_n171 ) );
  AND2_X1 u2_u7_u6_U19 (.A1( u2_u7_u6_n100 ) , .ZN( u2_u7_u6_n130 ) , .A2( u2_u7_u6_n147 ) );
  INV_X1 u2_u7_u6_U20 (.A( u2_u7_u6_n127 ) , .ZN( u2_u7_u6_n173 ) );
  INV_X1 u2_u7_u6_U21 (.A( u2_u7_u6_n121 ) , .ZN( u2_u7_u6_n167 ) );
  INV_X1 u2_u7_u6_U22 (.A( u2_u7_u6_n100 ) , .ZN( u2_u7_u6_n169 ) );
  INV_X1 u2_u7_u6_U23 (.A( u2_u7_u6_n123 ) , .ZN( u2_u7_u6_n170 ) );
  INV_X1 u2_u7_u6_U24 (.A( u2_u7_u6_n113 ) , .ZN( u2_u7_u6_n168 ) );
  AND2_X1 u2_u7_u6_U25 (.A1( u2_u7_u6_n107 ) , .A2( u2_u7_u6_n119 ) , .ZN( u2_u7_u6_n133 ) );
  AND2_X1 u2_u7_u6_U26 (.A2( u2_u7_u6_n121 ) , .A1( u2_u7_u6_n122 ) , .ZN( u2_u7_u6_n131 ) );
  AND3_X1 u2_u7_u6_U27 (.ZN( u2_u7_u6_n120 ) , .A2( u2_u7_u6_n127 ) , .A1( u2_u7_u6_n132 ) , .A3( u2_u7_u6_n145 ) );
  INV_X1 u2_u7_u6_U28 (.A( u2_u7_u6_n146 ) , .ZN( u2_u7_u6_n163 ) );
  AOI222_X1 u2_u7_u6_U29 (.ZN( u2_u7_u6_n114 ) , .A1( u2_u7_u6_n118 ) , .A2( u2_u7_u6_n126 ) , .B2( u2_u7_u6_n151 ) , .C2( u2_u7_u6_n159 ) , .C1( u2_u7_u6_n168 ) , .B1( u2_u7_u6_n169 ) );
  INV_X1 u2_u7_u6_U3 (.A( u2_u7_u6_n110 ) , .ZN( u2_u7_u6_n166 ) );
  NOR2_X1 u2_u7_u6_U30 (.A1( u2_u7_u6_n162 ) , .A2( u2_u7_u6_n165 ) , .ZN( u2_u7_u6_n98 ) );
  NAND2_X1 u2_u7_u6_U31 (.A1( u2_u7_u6_n144 ) , .ZN( u2_u7_u6_n151 ) , .A2( u2_u7_u6_n158 ) );
  NAND2_X1 u2_u7_u6_U32 (.ZN( u2_u7_u6_n132 ) , .A1( u2_u7_u6_n91 ) , .A2( u2_u7_u6_n97 ) );
  AOI22_X1 u2_u7_u6_U33 (.B2( u2_u7_u6_n110 ) , .B1( u2_u7_u6_n111 ) , .A1( u2_u7_u6_n112 ) , .ZN( u2_u7_u6_n115 ) , .A2( u2_u7_u6_n161 ) );
  NAND4_X1 u2_u7_u6_U34 (.A3( u2_u7_u6_n109 ) , .ZN( u2_u7_u6_n112 ) , .A4( u2_u7_u6_n132 ) , .A2( u2_u7_u6_n147 ) , .A1( u2_u7_u6_n166 ) );
  NOR2_X1 u2_u7_u6_U35 (.ZN( u2_u7_u6_n109 ) , .A1( u2_u7_u6_n170 ) , .A2( u2_u7_u6_n173 ) );
  NOR2_X1 u2_u7_u6_U36 (.A2( u2_u7_u6_n126 ) , .ZN( u2_u7_u6_n155 ) , .A1( u2_u7_u6_n160 ) );
  NAND2_X1 u2_u7_u6_U37 (.ZN( u2_u7_u6_n146 ) , .A2( u2_u7_u6_n94 ) , .A1( u2_u7_u6_n99 ) );
  AOI21_X1 u2_u7_u6_U38 (.A( u2_u7_u6_n144 ) , .B2( u2_u7_u6_n145 ) , .B1( u2_u7_u6_n146 ) , .ZN( u2_u7_u6_n150 ) );
  AOI211_X1 u2_u7_u6_U39 (.B( u2_u7_u6_n134 ) , .A( u2_u7_u6_n135 ) , .C1( u2_u7_u6_n136 ) , .ZN( u2_u7_u6_n137 ) , .C2( u2_u7_u6_n151 ) );
  INV_X1 u2_u7_u6_U4 (.A( u2_u7_u6_n142 ) , .ZN( u2_u7_u6_n174 ) );
  NAND4_X1 u2_u7_u6_U40 (.A4( u2_u7_u6_n127 ) , .A3( u2_u7_u6_n128 ) , .A2( u2_u7_u6_n129 ) , .A1( u2_u7_u6_n130 ) , .ZN( u2_u7_u6_n136 ) );
  AOI21_X1 u2_u7_u6_U41 (.B2( u2_u7_u6_n132 ) , .B1( u2_u7_u6_n133 ) , .ZN( u2_u7_u6_n134 ) , .A( u2_u7_u6_n158 ) );
  AOI21_X1 u2_u7_u6_U42 (.B1( u2_u7_u6_n131 ) , .ZN( u2_u7_u6_n135 ) , .A( u2_u7_u6_n144 ) , .B2( u2_u7_u6_n146 ) );
  INV_X1 u2_u7_u6_U43 (.A( u2_u7_u6_n111 ) , .ZN( u2_u7_u6_n158 ) );
  NAND2_X1 u2_u7_u6_U44 (.ZN( u2_u7_u6_n127 ) , .A1( u2_u7_u6_n91 ) , .A2( u2_u7_u6_n92 ) );
  NAND2_X1 u2_u7_u6_U45 (.ZN( u2_u7_u6_n129 ) , .A2( u2_u7_u6_n95 ) , .A1( u2_u7_u6_n96 ) );
  INV_X1 u2_u7_u6_U46 (.A( u2_u7_u6_n144 ) , .ZN( u2_u7_u6_n159 ) );
  NAND2_X1 u2_u7_u6_U47 (.ZN( u2_u7_u6_n145 ) , .A2( u2_u7_u6_n97 ) , .A1( u2_u7_u6_n98 ) );
  NAND2_X1 u2_u7_u6_U48 (.ZN( u2_u7_u6_n148 ) , .A2( u2_u7_u6_n92 ) , .A1( u2_u7_u6_n94 ) );
  NAND2_X1 u2_u7_u6_U49 (.ZN( u2_u7_u6_n108 ) , .A2( u2_u7_u6_n139 ) , .A1( u2_u7_u6_n144 ) );
  NAND2_X1 u2_u7_u6_U5 (.A2( u2_u7_u6_n143 ) , .ZN( u2_u7_u6_n152 ) , .A1( u2_u7_u6_n166 ) );
  NAND2_X1 u2_u7_u6_U50 (.ZN( u2_u7_u6_n121 ) , .A2( u2_u7_u6_n95 ) , .A1( u2_u7_u6_n97 ) );
  NAND2_X1 u2_u7_u6_U51 (.ZN( u2_u7_u6_n107 ) , .A2( u2_u7_u6_n92 ) , .A1( u2_u7_u6_n95 ) );
  AND2_X1 u2_u7_u6_U52 (.ZN( u2_u7_u6_n118 ) , .A2( u2_u7_u6_n91 ) , .A1( u2_u7_u6_n99 ) );
  NAND2_X1 u2_u7_u6_U53 (.ZN( u2_u7_u6_n147 ) , .A2( u2_u7_u6_n98 ) , .A1( u2_u7_u6_n99 ) );
  NAND2_X1 u2_u7_u6_U54 (.ZN( u2_u7_u6_n128 ) , .A1( u2_u7_u6_n94 ) , .A2( u2_u7_u6_n96 ) );
  NAND2_X1 u2_u7_u6_U55 (.ZN( u2_u7_u6_n119 ) , .A2( u2_u7_u6_n95 ) , .A1( u2_u7_u6_n99 ) );
  NAND2_X1 u2_u7_u6_U56 (.ZN( u2_u7_u6_n123 ) , .A2( u2_u7_u6_n91 ) , .A1( u2_u7_u6_n96 ) );
  NAND2_X1 u2_u7_u6_U57 (.ZN( u2_u7_u6_n100 ) , .A2( u2_u7_u6_n92 ) , .A1( u2_u7_u6_n98 ) );
  NAND2_X1 u2_u7_u6_U58 (.ZN( u2_u7_u6_n122 ) , .A1( u2_u7_u6_n94 ) , .A2( u2_u7_u6_n97 ) );
  INV_X1 u2_u7_u6_U59 (.A( u2_u7_u6_n139 ) , .ZN( u2_u7_u6_n160 ) );
  AOI22_X1 u2_u7_u6_U6 (.B2( u2_u7_u6_n101 ) , .A1( u2_u7_u6_n102 ) , .ZN( u2_u7_u6_n103 ) , .B1( u2_u7_u6_n160 ) , .A2( u2_u7_u6_n161 ) );
  NAND2_X1 u2_u7_u6_U60 (.ZN( u2_u7_u6_n113 ) , .A1( u2_u7_u6_n96 ) , .A2( u2_u7_u6_n98 ) );
  NOR2_X1 u2_u7_u6_U61 (.A2( u2_u7_X_40 ) , .A1( u2_u7_X_41 ) , .ZN( u2_u7_u6_n126 ) );
  NOR2_X1 u2_u7_u6_U62 (.A2( u2_u7_X_39 ) , .A1( u2_u7_X_42 ) , .ZN( u2_u7_u6_n92 ) );
  NOR2_X1 u2_u7_u6_U63 (.A2( u2_u7_X_39 ) , .A1( u2_u7_u6_n156 ) , .ZN( u2_u7_u6_n97 ) );
  NOR2_X1 u2_u7_u6_U64 (.A2( u2_u7_X_38 ) , .A1( u2_u7_u6_n165 ) , .ZN( u2_u7_u6_n95 ) );
  NOR2_X1 u2_u7_u6_U65 (.A2( u2_u7_X_41 ) , .ZN( u2_u7_u6_n111 ) , .A1( u2_u7_u6_n157 ) );
  NOR2_X1 u2_u7_u6_U66 (.A2( u2_u7_X_37 ) , .A1( u2_u7_u6_n162 ) , .ZN( u2_u7_u6_n94 ) );
  NOR2_X1 u2_u7_u6_U67 (.A2( u2_u7_X_37 ) , .A1( u2_u7_X_38 ) , .ZN( u2_u7_u6_n91 ) );
  NAND2_X1 u2_u7_u6_U68 (.A1( u2_u7_X_41 ) , .ZN( u2_u7_u6_n144 ) , .A2( u2_u7_u6_n157 ) );
  NAND2_X1 u2_u7_u6_U69 (.A2( u2_u7_X_40 ) , .A1( u2_u7_X_41 ) , .ZN( u2_u7_u6_n139 ) );
  NOR2_X1 u2_u7_u6_U7 (.A1( u2_u7_u6_n118 ) , .ZN( u2_u7_u6_n143 ) , .A2( u2_u7_u6_n168 ) );
  AND2_X1 u2_u7_u6_U70 (.A1( u2_u7_X_39 ) , .A2( u2_u7_u6_n156 ) , .ZN( u2_u7_u6_n96 ) );
  AND2_X1 u2_u7_u6_U71 (.A1( u2_u7_X_39 ) , .A2( u2_u7_X_42 ) , .ZN( u2_u7_u6_n99 ) );
  INV_X1 u2_u7_u6_U72 (.A( u2_u7_X_40 ) , .ZN( u2_u7_u6_n157 ) );
  INV_X1 u2_u7_u6_U73 (.A( u2_u7_X_37 ) , .ZN( u2_u7_u6_n165 ) );
  INV_X1 u2_u7_u6_U74 (.A( u2_u7_X_38 ) , .ZN( u2_u7_u6_n162 ) );
  INV_X1 u2_u7_u6_U75 (.A( u2_u7_X_42 ) , .ZN( u2_u7_u6_n156 ) );
  NAND4_X1 u2_u7_u6_U76 (.ZN( u2_out7_12 ) , .A4( u2_u7_u6_n114 ) , .A3( u2_u7_u6_n115 ) , .A2( u2_u7_u6_n116 ) , .A1( u2_u7_u6_n117 ) );
  OAI22_X1 u2_u7_u6_U77 (.B2( u2_u7_u6_n111 ) , .ZN( u2_u7_u6_n116 ) , .B1( u2_u7_u6_n126 ) , .A2( u2_u7_u6_n164 ) , .A1( u2_u7_u6_n167 ) );
  OAI21_X1 u2_u7_u6_U78 (.A( u2_u7_u6_n108 ) , .ZN( u2_u7_u6_n117 ) , .B2( u2_u7_u6_n141 ) , .B1( u2_u7_u6_n163 ) );
  NAND4_X1 u2_u7_u6_U79 (.ZN( u2_out7_32 ) , .A4( u2_u7_u6_n103 ) , .A3( u2_u7_u6_n104 ) , .A2( u2_u7_u6_n105 ) , .A1( u2_u7_u6_n106 ) );
  AOI21_X1 u2_u7_u6_U8 (.B1( u2_u7_u6_n107 ) , .B2( u2_u7_u6_n132 ) , .A( u2_u7_u6_n158 ) , .ZN( u2_u7_u6_n88 ) );
  AOI22_X1 u2_u7_u6_U80 (.ZN( u2_u7_u6_n105 ) , .A2( u2_u7_u6_n108 ) , .A1( u2_u7_u6_n118 ) , .B2( u2_u7_u6_n126 ) , .B1( u2_u7_u6_n171 ) );
  AOI22_X1 u2_u7_u6_U81 (.ZN( u2_u7_u6_n104 ) , .A1( u2_u7_u6_n111 ) , .B1( u2_u7_u6_n124 ) , .B2( u2_u7_u6_n151 ) , .A2( u2_u7_u6_n93 ) );
  OAI211_X1 u2_u7_u6_U82 (.ZN( u2_out7_22 ) , .B( u2_u7_u6_n137 ) , .A( u2_u7_u6_n138 ) , .C2( u2_u7_u6_n139 ) , .C1( u2_u7_u6_n140 ) );
  AOI22_X1 u2_u7_u6_U83 (.B1( u2_u7_u6_n124 ) , .A2( u2_u7_u6_n125 ) , .A1( u2_u7_u6_n126 ) , .ZN( u2_u7_u6_n138 ) , .B2( u2_u7_u6_n161 ) );
  AND4_X1 u2_u7_u6_U84 (.A3( u2_u7_u6_n119 ) , .A1( u2_u7_u6_n120 ) , .A4( u2_u7_u6_n129 ) , .ZN( u2_u7_u6_n140 ) , .A2( u2_u7_u6_n143 ) );
  OAI211_X1 u2_u7_u6_U85 (.ZN( u2_out7_7 ) , .B( u2_u7_u6_n153 ) , .C2( u2_u7_u6_n154 ) , .C1( u2_u7_u6_n155 ) , .A( u2_u7_u6_n174 ) );
  NOR3_X1 u2_u7_u6_U86 (.A1( u2_u7_u6_n141 ) , .ZN( u2_u7_u6_n154 ) , .A3( u2_u7_u6_n164 ) , .A2( u2_u7_u6_n171 ) );
  AOI211_X1 u2_u7_u6_U87 (.B( u2_u7_u6_n149 ) , .A( u2_u7_u6_n150 ) , .C2( u2_u7_u6_n151 ) , .C1( u2_u7_u6_n152 ) , .ZN( u2_u7_u6_n153 ) );
  NAND3_X1 u2_u7_u6_U88 (.A2( u2_u7_u6_n123 ) , .ZN( u2_u7_u6_n125 ) , .A1( u2_u7_u6_n130 ) , .A3( u2_u7_u6_n131 ) );
  NAND3_X1 u2_u7_u6_U89 (.A3( u2_u7_u6_n133 ) , .ZN( u2_u7_u6_n141 ) , .A1( u2_u7_u6_n145 ) , .A2( u2_u7_u6_n148 ) );
  AOI21_X1 u2_u7_u6_U9 (.B2( u2_u7_u6_n147 ) , .B1( u2_u7_u6_n148 ) , .ZN( u2_u7_u6_n149 ) , .A( u2_u7_u6_n158 ) );
  NAND3_X1 u2_u7_u6_U90 (.ZN( u2_u7_u6_n101 ) , .A3( u2_u7_u6_n107 ) , .A2( u2_u7_u6_n121 ) , .A1( u2_u7_u6_n127 ) );
  NAND3_X1 u2_u7_u6_U91 (.ZN( u2_u7_u6_n102 ) , .A3( u2_u7_u6_n130 ) , .A2( u2_u7_u6_n145 ) , .A1( u2_u7_u6_n166 ) );
  NAND3_X1 u2_u7_u6_U92 (.A3( u2_u7_u6_n113 ) , .A1( u2_u7_u6_n119 ) , .A2( u2_u7_u6_n123 ) , .ZN( u2_u7_u6_n93 ) );
  NAND3_X1 u2_u7_u6_U93 (.ZN( u2_u7_u6_n142 ) , .A2( u2_u7_u6_n172 ) , .A3( u2_u7_u6_n89 ) , .A1( u2_u7_u6_n90 ) );
  OAI21_X1 u2_u7_u7_U10 (.A( u2_u7_u7_n161 ) , .B1( u2_u7_u7_n168 ) , .B2( u2_u7_u7_n173 ) , .ZN( u2_u7_u7_n91 ) );
  AOI211_X1 u2_u7_u7_U11 (.A( u2_u7_u7_n117 ) , .ZN( u2_u7_u7_n118 ) , .C2( u2_u7_u7_n126 ) , .C1( u2_u7_u7_n177 ) , .B( u2_u7_u7_n180 ) );
  OAI22_X1 u2_u7_u7_U12 (.B1( u2_u7_u7_n115 ) , .ZN( u2_u7_u7_n117 ) , .A2( u2_u7_u7_n133 ) , .A1( u2_u7_u7_n137 ) , .B2( u2_u7_u7_n162 ) );
  INV_X1 u2_u7_u7_U13 (.A( u2_u7_u7_n116 ) , .ZN( u2_u7_u7_n180 ) );
  NOR3_X1 u2_u7_u7_U14 (.ZN( u2_u7_u7_n115 ) , .A3( u2_u7_u7_n145 ) , .A2( u2_u7_u7_n168 ) , .A1( u2_u7_u7_n169 ) );
  INV_X1 u2_u7_u7_U15 (.A( u2_u7_u7_n133 ) , .ZN( u2_u7_u7_n176 ) );
  NOR3_X1 u2_u7_u7_U16 (.A2( u2_u7_u7_n134 ) , .A1( u2_u7_u7_n135 ) , .ZN( u2_u7_u7_n136 ) , .A3( u2_u7_u7_n171 ) );
  NOR2_X1 u2_u7_u7_U17 (.A1( u2_u7_u7_n130 ) , .A2( u2_u7_u7_n134 ) , .ZN( u2_u7_u7_n153 ) );
  AOI21_X1 u2_u7_u7_U18 (.ZN( u2_u7_u7_n104 ) , .B2( u2_u7_u7_n112 ) , .B1( u2_u7_u7_n127 ) , .A( u2_u7_u7_n164 ) );
  AOI21_X1 u2_u7_u7_U19 (.ZN( u2_u7_u7_n106 ) , .B1( u2_u7_u7_n133 ) , .B2( u2_u7_u7_n146 ) , .A( u2_u7_u7_n162 ) );
  AOI21_X1 u2_u7_u7_U20 (.A( u2_u7_u7_n101 ) , .ZN( u2_u7_u7_n107 ) , .B2( u2_u7_u7_n128 ) , .B1( u2_u7_u7_n175 ) );
  INV_X1 u2_u7_u7_U21 (.A( u2_u7_u7_n101 ) , .ZN( u2_u7_u7_n165 ) );
  NOR2_X1 u2_u7_u7_U22 (.ZN( u2_u7_u7_n111 ) , .A2( u2_u7_u7_n134 ) , .A1( u2_u7_u7_n169 ) );
  INV_X1 u2_u7_u7_U23 (.A( u2_u7_u7_n138 ) , .ZN( u2_u7_u7_n171 ) );
  INV_X1 u2_u7_u7_U24 (.A( u2_u7_u7_n131 ) , .ZN( u2_u7_u7_n177 ) );
  INV_X1 u2_u7_u7_U25 (.A( u2_u7_u7_n110 ) , .ZN( u2_u7_u7_n174 ) );
  NAND2_X1 u2_u7_u7_U26 (.A1( u2_u7_u7_n129 ) , .A2( u2_u7_u7_n132 ) , .ZN( u2_u7_u7_n149 ) );
  NAND2_X1 u2_u7_u7_U27 (.A1( u2_u7_u7_n113 ) , .A2( u2_u7_u7_n124 ) , .ZN( u2_u7_u7_n130 ) );
  INV_X1 u2_u7_u7_U28 (.A( u2_u7_u7_n112 ) , .ZN( u2_u7_u7_n173 ) );
  INV_X1 u2_u7_u7_U29 (.A( u2_u7_u7_n128 ) , .ZN( u2_u7_u7_n168 ) );
  OAI21_X1 u2_u7_u7_U3 (.ZN( u2_u7_u7_n159 ) , .A( u2_u7_u7_n165 ) , .B2( u2_u7_u7_n171 ) , .B1( u2_u7_u7_n174 ) );
  INV_X1 u2_u7_u7_U30 (.A( u2_u7_u7_n148 ) , .ZN( u2_u7_u7_n169 ) );
  INV_X1 u2_u7_u7_U31 (.A( u2_u7_u7_n127 ) , .ZN( u2_u7_u7_n179 ) );
  NOR2_X1 u2_u7_u7_U32 (.ZN( u2_u7_u7_n101 ) , .A2( u2_u7_u7_n150 ) , .A1( u2_u7_u7_n156 ) );
  AOI211_X1 u2_u7_u7_U33 (.B( u2_u7_u7_n139 ) , .A( u2_u7_u7_n140 ) , .C2( u2_u7_u7_n141 ) , .ZN( u2_u7_u7_n142 ) , .C1( u2_u7_u7_n156 ) );
  NAND4_X1 u2_u7_u7_U34 (.A3( u2_u7_u7_n127 ) , .A2( u2_u7_u7_n128 ) , .A1( u2_u7_u7_n129 ) , .ZN( u2_u7_u7_n141 ) , .A4( u2_u7_u7_n147 ) );
  AOI21_X1 u2_u7_u7_U35 (.A( u2_u7_u7_n137 ) , .B1( u2_u7_u7_n138 ) , .ZN( u2_u7_u7_n139 ) , .B2( u2_u7_u7_n146 ) );
  OAI22_X1 u2_u7_u7_U36 (.B1( u2_u7_u7_n136 ) , .ZN( u2_u7_u7_n140 ) , .A1( u2_u7_u7_n153 ) , .B2( u2_u7_u7_n162 ) , .A2( u2_u7_u7_n164 ) );
  INV_X1 u2_u7_u7_U37 (.A( u2_u7_u7_n125 ) , .ZN( u2_u7_u7_n161 ) );
  AOI21_X1 u2_u7_u7_U38 (.ZN( u2_u7_u7_n123 ) , .B1( u2_u7_u7_n165 ) , .B2( u2_u7_u7_n177 ) , .A( u2_u7_u7_n97 ) );
  AOI21_X1 u2_u7_u7_U39 (.B2( u2_u7_u7_n113 ) , .B1( u2_u7_u7_n124 ) , .A( u2_u7_u7_n125 ) , .ZN( u2_u7_u7_n97 ) );
  INV_X1 u2_u7_u7_U4 (.A( u2_u7_u7_n149 ) , .ZN( u2_u7_u7_n175 ) );
  INV_X1 u2_u7_u7_U40 (.A( u2_u7_u7_n152 ) , .ZN( u2_u7_u7_n162 ) );
  AOI22_X1 u2_u7_u7_U41 (.A2( u2_u7_u7_n114 ) , .ZN( u2_u7_u7_n119 ) , .B1( u2_u7_u7_n130 ) , .A1( u2_u7_u7_n156 ) , .B2( u2_u7_u7_n165 ) );
  NAND2_X1 u2_u7_u7_U42 (.A2( u2_u7_u7_n112 ) , .ZN( u2_u7_u7_n114 ) , .A1( u2_u7_u7_n175 ) );
  NOR2_X1 u2_u7_u7_U43 (.ZN( u2_u7_u7_n137 ) , .A1( u2_u7_u7_n150 ) , .A2( u2_u7_u7_n161 ) );
  AND2_X1 u2_u7_u7_U44 (.ZN( u2_u7_u7_n145 ) , .A2( u2_u7_u7_n98 ) , .A1( u2_u7_u7_n99 ) );
  AOI21_X1 u2_u7_u7_U45 (.ZN( u2_u7_u7_n105 ) , .B2( u2_u7_u7_n110 ) , .A( u2_u7_u7_n125 ) , .B1( u2_u7_u7_n147 ) );
  NAND2_X1 u2_u7_u7_U46 (.ZN( u2_u7_u7_n146 ) , .A1( u2_u7_u7_n95 ) , .A2( u2_u7_u7_n98 ) );
  NAND2_X1 u2_u7_u7_U47 (.A2( u2_u7_u7_n103 ) , .ZN( u2_u7_u7_n147 ) , .A1( u2_u7_u7_n93 ) );
  NAND2_X1 u2_u7_u7_U48 (.A1( u2_u7_u7_n103 ) , .ZN( u2_u7_u7_n127 ) , .A2( u2_u7_u7_n99 ) );
  NAND2_X1 u2_u7_u7_U49 (.A2( u2_u7_u7_n102 ) , .A1( u2_u7_u7_n103 ) , .ZN( u2_u7_u7_n133 ) );
  INV_X1 u2_u7_u7_U5 (.A( u2_u7_u7_n154 ) , .ZN( u2_u7_u7_n178 ) );
  OR2_X1 u2_u7_u7_U50 (.ZN( u2_u7_u7_n126 ) , .A2( u2_u7_u7_n152 ) , .A1( u2_u7_u7_n156 ) );
  NAND2_X1 u2_u7_u7_U51 (.ZN( u2_u7_u7_n112 ) , .A2( u2_u7_u7_n96 ) , .A1( u2_u7_u7_n99 ) );
  NAND2_X1 u2_u7_u7_U52 (.A2( u2_u7_u7_n102 ) , .ZN( u2_u7_u7_n128 ) , .A1( u2_u7_u7_n98 ) );
  NAND2_X1 u2_u7_u7_U53 (.A1( u2_u7_u7_n100 ) , .ZN( u2_u7_u7_n113 ) , .A2( u2_u7_u7_n93 ) );
  NAND2_X1 u2_u7_u7_U54 (.ZN( u2_u7_u7_n110 ) , .A1( u2_u7_u7_n95 ) , .A2( u2_u7_u7_n96 ) );
  INV_X1 u2_u7_u7_U55 (.A( u2_u7_u7_n150 ) , .ZN( u2_u7_u7_n164 ) );
  AND2_X1 u2_u7_u7_U56 (.ZN( u2_u7_u7_n134 ) , .A1( u2_u7_u7_n93 ) , .A2( u2_u7_u7_n98 ) );
  NAND2_X1 u2_u7_u7_U57 (.A2( u2_u7_u7_n102 ) , .ZN( u2_u7_u7_n124 ) , .A1( u2_u7_u7_n96 ) );
  NAND2_X1 u2_u7_u7_U58 (.A1( u2_u7_u7_n100 ) , .A2( u2_u7_u7_n102 ) , .ZN( u2_u7_u7_n129 ) );
  NAND2_X1 u2_u7_u7_U59 (.A2( u2_u7_u7_n103 ) , .ZN( u2_u7_u7_n131 ) , .A1( u2_u7_u7_n95 ) );
  AOI211_X1 u2_u7_u7_U6 (.ZN( u2_u7_u7_n116 ) , .A( u2_u7_u7_n155 ) , .C1( u2_u7_u7_n161 ) , .C2( u2_u7_u7_n171 ) , .B( u2_u7_u7_n94 ) );
  NAND2_X1 u2_u7_u7_U60 (.A1( u2_u7_u7_n100 ) , .ZN( u2_u7_u7_n138 ) , .A2( u2_u7_u7_n99 ) );
  NAND2_X1 u2_u7_u7_U61 (.ZN( u2_u7_u7_n132 ) , .A1( u2_u7_u7_n93 ) , .A2( u2_u7_u7_n96 ) );
  NAND2_X1 u2_u7_u7_U62 (.A1( u2_u7_u7_n100 ) , .ZN( u2_u7_u7_n148 ) , .A2( u2_u7_u7_n95 ) );
  AOI211_X1 u2_u7_u7_U63 (.B( u2_u7_u7_n154 ) , .A( u2_u7_u7_n155 ) , .C1( u2_u7_u7_n156 ) , .ZN( u2_u7_u7_n157 ) , .C2( u2_u7_u7_n172 ) );
  INV_X1 u2_u7_u7_U64 (.A( u2_u7_u7_n153 ) , .ZN( u2_u7_u7_n172 ) );
  NOR2_X1 u2_u7_u7_U65 (.A2( u2_u7_X_47 ) , .ZN( u2_u7_u7_n150 ) , .A1( u2_u7_u7_n163 ) );
  NOR2_X1 u2_u7_u7_U66 (.A2( u2_u7_X_43 ) , .A1( u2_u7_X_44 ) , .ZN( u2_u7_u7_n103 ) );
  NOR2_X1 u2_u7_u7_U67 (.A2( u2_u7_X_48 ) , .A1( u2_u7_u7_n166 ) , .ZN( u2_u7_u7_n95 ) );
  NOR2_X1 u2_u7_u7_U68 (.A2( u2_u7_X_45 ) , .A1( u2_u7_X_48 ) , .ZN( u2_u7_u7_n99 ) );
  NOR2_X1 u2_u7_u7_U69 (.A2( u2_u7_X_44 ) , .A1( u2_u7_u7_n167 ) , .ZN( u2_u7_u7_n98 ) );
  OAI222_X1 u2_u7_u7_U7 (.C2( u2_u7_u7_n101 ) , .B2( u2_u7_u7_n111 ) , .A1( u2_u7_u7_n113 ) , .C1( u2_u7_u7_n146 ) , .A2( u2_u7_u7_n162 ) , .B1( u2_u7_u7_n164 ) , .ZN( u2_u7_u7_n94 ) );
  NOR2_X1 u2_u7_u7_U70 (.A2( u2_u7_X_46 ) , .A1( u2_u7_X_47 ) , .ZN( u2_u7_u7_n152 ) );
  NAND2_X1 u2_u7_u7_U71 (.A2( u2_u7_X_46 ) , .A1( u2_u7_X_47 ) , .ZN( u2_u7_u7_n125 ) );
  AND2_X1 u2_u7_u7_U72 (.A1( u2_u7_X_47 ) , .ZN( u2_u7_u7_n156 ) , .A2( u2_u7_u7_n163 ) );
  AND2_X1 u2_u7_u7_U73 (.A2( u2_u7_X_45 ) , .A1( u2_u7_X_48 ) , .ZN( u2_u7_u7_n102 ) );
  AND2_X1 u2_u7_u7_U74 (.A2( u2_u7_X_43 ) , .A1( u2_u7_X_44 ) , .ZN( u2_u7_u7_n96 ) );
  AND2_X1 u2_u7_u7_U75 (.A1( u2_u7_X_44 ) , .ZN( u2_u7_u7_n100 ) , .A2( u2_u7_u7_n167 ) );
  AND2_X1 u2_u7_u7_U76 (.A1( u2_u7_X_48 ) , .A2( u2_u7_u7_n166 ) , .ZN( u2_u7_u7_n93 ) );
  INV_X1 u2_u7_u7_U77 (.A( u2_u7_X_46 ) , .ZN( u2_u7_u7_n163 ) );
  INV_X1 u2_u7_u7_U78 (.A( u2_u7_X_43 ) , .ZN( u2_u7_u7_n167 ) );
  INV_X1 u2_u7_u7_U79 (.A( u2_u7_X_45 ) , .ZN( u2_u7_u7_n166 ) );
  OAI221_X1 u2_u7_u7_U8 (.C1( u2_u7_u7_n101 ) , .C2( u2_u7_u7_n147 ) , .ZN( u2_u7_u7_n155 ) , .B2( u2_u7_u7_n162 ) , .A( u2_u7_u7_n91 ) , .B1( u2_u7_u7_n92 ) );
  NAND4_X1 u2_u7_u7_U80 (.ZN( u2_out7_5 ) , .A4( u2_u7_u7_n108 ) , .A3( u2_u7_u7_n109 ) , .A1( u2_u7_u7_n116 ) , .A2( u2_u7_u7_n123 ) );
  AOI22_X1 u2_u7_u7_U81 (.ZN( u2_u7_u7_n109 ) , .A2( u2_u7_u7_n126 ) , .B2( u2_u7_u7_n145 ) , .B1( u2_u7_u7_n156 ) , .A1( u2_u7_u7_n171 ) );
  NOR4_X1 u2_u7_u7_U82 (.A4( u2_u7_u7_n104 ) , .A3( u2_u7_u7_n105 ) , .A2( u2_u7_u7_n106 ) , .A1( u2_u7_u7_n107 ) , .ZN( u2_u7_u7_n108 ) );
  NAND4_X1 u2_u7_u7_U83 (.ZN( u2_out7_27 ) , .A4( u2_u7_u7_n118 ) , .A3( u2_u7_u7_n119 ) , .A2( u2_u7_u7_n120 ) , .A1( u2_u7_u7_n121 ) );
  OAI21_X1 u2_u7_u7_U84 (.ZN( u2_u7_u7_n121 ) , .B2( u2_u7_u7_n145 ) , .A( u2_u7_u7_n150 ) , .B1( u2_u7_u7_n174 ) );
  OAI21_X1 u2_u7_u7_U85 (.ZN( u2_u7_u7_n120 ) , .A( u2_u7_u7_n161 ) , .B2( u2_u7_u7_n170 ) , .B1( u2_u7_u7_n179 ) );
  NAND4_X1 u2_u7_u7_U86 (.ZN( u2_out7_21 ) , .A4( u2_u7_u7_n157 ) , .A3( u2_u7_u7_n158 ) , .A2( u2_u7_u7_n159 ) , .A1( u2_u7_u7_n160 ) );
  OAI21_X1 u2_u7_u7_U87 (.B1( u2_u7_u7_n145 ) , .ZN( u2_u7_u7_n160 ) , .A( u2_u7_u7_n161 ) , .B2( u2_u7_u7_n177 ) );
  AOI22_X1 u2_u7_u7_U88 (.B2( u2_u7_u7_n149 ) , .B1( u2_u7_u7_n150 ) , .A2( u2_u7_u7_n151 ) , .A1( u2_u7_u7_n152 ) , .ZN( u2_u7_u7_n158 ) );
  NAND4_X1 u2_u7_u7_U89 (.ZN( u2_out7_15 ) , .A4( u2_u7_u7_n142 ) , .A3( u2_u7_u7_n143 ) , .A2( u2_u7_u7_n144 ) , .A1( u2_u7_u7_n178 ) );
  AND3_X1 u2_u7_u7_U9 (.A3( u2_u7_u7_n110 ) , .A2( u2_u7_u7_n127 ) , .A1( u2_u7_u7_n132 ) , .ZN( u2_u7_u7_n92 ) );
  OR2_X1 u2_u7_u7_U90 (.A2( u2_u7_u7_n125 ) , .A1( u2_u7_u7_n129 ) , .ZN( u2_u7_u7_n144 ) );
  AOI22_X1 u2_u7_u7_U91 (.A2( u2_u7_u7_n126 ) , .ZN( u2_u7_u7_n143 ) , .B2( u2_u7_u7_n165 ) , .B1( u2_u7_u7_n173 ) , .A1( u2_u7_u7_n174 ) );
  OAI211_X1 u2_u7_u7_U92 (.B( u2_u7_u7_n122 ) , .A( u2_u7_u7_n123 ) , .C2( u2_u7_u7_n124 ) , .ZN( u2_u7_u7_n154 ) , .C1( u2_u7_u7_n162 ) );
  AOI222_X1 u2_u7_u7_U93 (.ZN( u2_u7_u7_n122 ) , .C2( u2_u7_u7_n126 ) , .C1( u2_u7_u7_n145 ) , .B1( u2_u7_u7_n161 ) , .A2( u2_u7_u7_n165 ) , .B2( u2_u7_u7_n170 ) , .A1( u2_u7_u7_n176 ) );
  INV_X1 u2_u7_u7_U94 (.A( u2_u7_u7_n111 ) , .ZN( u2_u7_u7_n170 ) );
  NAND3_X1 u2_u7_u7_U95 (.A3( u2_u7_u7_n146 ) , .A2( u2_u7_u7_n147 ) , .A1( u2_u7_u7_n148 ) , .ZN( u2_u7_u7_n151 ) );
  NAND3_X1 u2_u7_u7_U96 (.A3( u2_u7_u7_n131 ) , .A2( u2_u7_u7_n132 ) , .A1( u2_u7_u7_n133 ) , .ZN( u2_u7_u7_n135 ) );
  XOR2_X1 u2_u9_U1 (.B( u2_K10_9 ) , .A( u2_R8_6 ) , .Z( u2_u9_X_9 ) );
  XOR2_X1 u2_u9_U10 (.B( u2_K10_45 ) , .A( u2_R8_30 ) , .Z( u2_u9_X_45 ) );
  XOR2_X1 u2_u9_U11 (.B( u2_K10_44 ) , .A( u2_R8_29 ) , .Z( u2_u9_X_44 ) );
  XOR2_X1 u2_u9_U12 (.B( u2_K10_43 ) , .A( u2_R8_28 ) , .Z( u2_u9_X_43 ) );
  XOR2_X1 u2_u9_U16 (.B( u2_K10_3 ) , .A( u2_R8_2 ) , .Z( u2_u9_X_3 ) );
  XOR2_X1 u2_u9_U2 (.B( u2_K10_8 ) , .A( u2_R8_5 ) , .Z( u2_u9_X_8 ) );
  XOR2_X1 u2_u9_U27 (.B( u2_K10_2 ) , .A( u2_R8_1 ) , .Z( u2_u9_X_2 ) );
  XOR2_X1 u2_u9_U3 (.B( u2_K10_7 ) , .A( u2_R8_4 ) , .Z( u2_u9_X_7 ) );
  XOR2_X1 u2_u9_U38 (.B( u2_K10_1 ) , .A( u2_R8_32 ) , .Z( u2_u9_X_1 ) );
  XOR2_X1 u2_u9_U4 (.B( u2_K10_6 ) , .A( u2_R8_5 ) , .Z( u2_u9_X_6 ) );
  XOR2_X1 u2_u9_U40 (.B( u2_K10_18 ) , .A( u2_R8_13 ) , .Z( u2_u9_X_18 ) );
  XOR2_X1 u2_u9_U41 (.B( u2_K10_17 ) , .A( u2_R8_12 ) , .Z( u2_u9_X_17 ) );
  XOR2_X1 u2_u9_U42 (.B( u2_K10_16 ) , .A( u2_R8_11 ) , .Z( u2_u9_X_16 ) );
  XOR2_X1 u2_u9_U43 (.B( u2_K10_15 ) , .A( u2_R8_10 ) , .Z( u2_u9_X_15 ) );
  XOR2_X1 u2_u9_U44 (.B( u2_K10_14 ) , .A( u2_R8_9 ) , .Z( u2_u9_X_14 ) );
  XOR2_X1 u2_u9_U45 (.B( u2_K10_13 ) , .A( u2_R8_8 ) , .Z( u2_u9_X_13 ) );
  XOR2_X1 u2_u9_U46 (.B( u2_K10_12 ) , .A( u2_R8_9 ) , .Z( u2_u9_X_12 ) );
  XOR2_X1 u2_u9_U47 (.B( u2_K10_11 ) , .A( u2_R8_8 ) , .Z( u2_u9_X_11 ) );
  XOR2_X1 u2_u9_U48 (.B( u2_K10_10 ) , .A( u2_R8_7 ) , .Z( u2_u9_X_10 ) );
  XOR2_X1 u2_u9_U5 (.B( u2_K10_5 ) , .A( u2_R8_4 ) , .Z( u2_u9_X_5 ) );
  XOR2_X1 u2_u9_U6 (.B( u2_K10_4 ) , .A( u2_R8_3 ) , .Z( u2_u9_X_4 ) );
  XOR2_X1 u2_u9_U7 (.B( u2_K10_48 ) , .A( u2_R8_1 ) , .Z( u2_u9_X_48 ) );
  XOR2_X1 u2_u9_U8 (.B( u2_K10_47 ) , .A( u2_R8_32 ) , .Z( u2_u9_X_47 ) );
  XOR2_X1 u2_u9_U9 (.B( u2_K10_46 ) , .A( u2_R8_31 ) , .Z( u2_u9_X_46 ) );
  AND3_X1 u2_u9_u0_U10 (.A2( u2_u9_u0_n112 ) , .ZN( u2_u9_u0_n127 ) , .A3( u2_u9_u0_n130 ) , .A1( u2_u9_u0_n148 ) );
  NAND2_X1 u2_u9_u0_U11 (.ZN( u2_u9_u0_n113 ) , .A1( u2_u9_u0_n139 ) , .A2( u2_u9_u0_n149 ) );
  AND2_X1 u2_u9_u0_U12 (.ZN( u2_u9_u0_n107 ) , .A1( u2_u9_u0_n130 ) , .A2( u2_u9_u0_n140 ) );
  AND2_X1 u2_u9_u0_U13 (.A2( u2_u9_u0_n129 ) , .A1( u2_u9_u0_n130 ) , .ZN( u2_u9_u0_n151 ) );
  AND2_X1 u2_u9_u0_U14 (.A1( u2_u9_u0_n108 ) , .A2( u2_u9_u0_n125 ) , .ZN( u2_u9_u0_n145 ) );
  INV_X1 u2_u9_u0_U15 (.A( u2_u9_u0_n143 ) , .ZN( u2_u9_u0_n173 ) );
  NOR2_X1 u2_u9_u0_U16 (.A2( u2_u9_u0_n136 ) , .ZN( u2_u9_u0_n147 ) , .A1( u2_u9_u0_n160 ) );
  OAI221_X1 u2_u9_u0_U17 (.C1( u2_u9_u0_n112 ) , .ZN( u2_u9_u0_n120 ) , .B1( u2_u9_u0_n138 ) , .B2( u2_u9_u0_n141 ) , .C2( u2_u9_u0_n147 ) , .A( u2_u9_u0_n172 ) );
  AOI211_X1 u2_u9_u0_U18 (.B( u2_u9_u0_n115 ) , .A( u2_u9_u0_n116 ) , .C2( u2_u9_u0_n117 ) , .C1( u2_u9_u0_n118 ) , .ZN( u2_u9_u0_n119 ) );
  OAI22_X1 u2_u9_u0_U19 (.B1( u2_u9_u0_n125 ) , .ZN( u2_u9_u0_n126 ) , .A1( u2_u9_u0_n138 ) , .A2( u2_u9_u0_n146 ) , .B2( u2_u9_u0_n147 ) );
  OAI22_X1 u2_u9_u0_U20 (.B1( u2_u9_u0_n131 ) , .A1( u2_u9_u0_n144 ) , .B2( u2_u9_u0_n147 ) , .A2( u2_u9_u0_n90 ) , .ZN( u2_u9_u0_n91 ) );
  AND3_X1 u2_u9_u0_U21 (.A3( u2_u9_u0_n121 ) , .A2( u2_u9_u0_n125 ) , .A1( u2_u9_u0_n148 ) , .ZN( u2_u9_u0_n90 ) );
  NOR2_X1 u2_u9_u0_U22 (.A1( u2_u9_u0_n163 ) , .A2( u2_u9_u0_n164 ) , .ZN( u2_u9_u0_n95 ) );
  INV_X1 u2_u9_u0_U23 (.A( u2_u9_u0_n136 ) , .ZN( u2_u9_u0_n161 ) );
  AOI22_X1 u2_u9_u0_U24 (.B2( u2_u9_u0_n109 ) , .A2( u2_u9_u0_n110 ) , .ZN( u2_u9_u0_n111 ) , .B1( u2_u9_u0_n118 ) , .A1( u2_u9_u0_n160 ) );
  INV_X1 u2_u9_u0_U25 (.A( u2_u9_u0_n118 ) , .ZN( u2_u9_u0_n158 ) );
  AOI21_X1 u2_u9_u0_U26 (.ZN( u2_u9_u0_n104 ) , .B1( u2_u9_u0_n107 ) , .B2( u2_u9_u0_n141 ) , .A( u2_u9_u0_n144 ) );
  AOI21_X1 u2_u9_u0_U27 (.B1( u2_u9_u0_n127 ) , .B2( u2_u9_u0_n129 ) , .A( u2_u9_u0_n138 ) , .ZN( u2_u9_u0_n96 ) );
  AOI21_X1 u2_u9_u0_U28 (.ZN( u2_u9_u0_n116 ) , .B2( u2_u9_u0_n142 ) , .A( u2_u9_u0_n144 ) , .B1( u2_u9_u0_n166 ) );
  NAND2_X1 u2_u9_u0_U29 (.A1( u2_u9_u0_n100 ) , .A2( u2_u9_u0_n103 ) , .ZN( u2_u9_u0_n125 ) );
  INV_X1 u2_u9_u0_U3 (.A( u2_u9_u0_n113 ) , .ZN( u2_u9_u0_n166 ) );
  NAND2_X1 u2_u9_u0_U30 (.A2( u2_u9_u0_n103 ) , .ZN( u2_u9_u0_n140 ) , .A1( u2_u9_u0_n94 ) );
  NAND2_X1 u2_u9_u0_U31 (.A1( u2_u9_u0_n101 ) , .A2( u2_u9_u0_n102 ) , .ZN( u2_u9_u0_n150 ) );
  INV_X1 u2_u9_u0_U32 (.A( u2_u9_u0_n138 ) , .ZN( u2_u9_u0_n160 ) );
  NAND2_X1 u2_u9_u0_U33 (.A2( u2_u9_u0_n102 ) , .A1( u2_u9_u0_n103 ) , .ZN( u2_u9_u0_n149 ) );
  NAND2_X1 u2_u9_u0_U34 (.A2( u2_u9_u0_n100 ) , .A1( u2_u9_u0_n101 ) , .ZN( u2_u9_u0_n139 ) );
  NAND2_X1 u2_u9_u0_U35 (.A2( u2_u9_u0_n100 ) , .ZN( u2_u9_u0_n131 ) , .A1( u2_u9_u0_n92 ) );
  NAND2_X1 u2_u9_u0_U36 (.ZN( u2_u9_u0_n108 ) , .A1( u2_u9_u0_n92 ) , .A2( u2_u9_u0_n94 ) );
  NAND2_X1 u2_u9_u0_U37 (.A2( u2_u9_u0_n102 ) , .ZN( u2_u9_u0_n114 ) , .A1( u2_u9_u0_n92 ) );
  NAND2_X1 u2_u9_u0_U38 (.A1( u2_u9_u0_n101 ) , .ZN( u2_u9_u0_n130 ) , .A2( u2_u9_u0_n94 ) );
  NAND2_X1 u2_u9_u0_U39 (.A2( u2_u9_u0_n101 ) , .ZN( u2_u9_u0_n121 ) , .A1( u2_u9_u0_n93 ) );
  AOI21_X1 u2_u9_u0_U4 (.B1( u2_u9_u0_n114 ) , .ZN( u2_u9_u0_n115 ) , .B2( u2_u9_u0_n129 ) , .A( u2_u9_u0_n161 ) );
  INV_X1 u2_u9_u0_U40 (.ZN( u2_u9_u0_n172 ) , .A( u2_u9_u0_n88 ) );
  OAI222_X1 u2_u9_u0_U41 (.C1( u2_u9_u0_n108 ) , .A1( u2_u9_u0_n125 ) , .B2( u2_u9_u0_n128 ) , .B1( u2_u9_u0_n144 ) , .A2( u2_u9_u0_n158 ) , .C2( u2_u9_u0_n161 ) , .ZN( u2_u9_u0_n88 ) );
  NAND2_X1 u2_u9_u0_U42 (.ZN( u2_u9_u0_n112 ) , .A2( u2_u9_u0_n92 ) , .A1( u2_u9_u0_n93 ) );
  OR3_X1 u2_u9_u0_U43 (.A3( u2_u9_u0_n152 ) , .A2( u2_u9_u0_n153 ) , .A1( u2_u9_u0_n154 ) , .ZN( u2_u9_u0_n155 ) );
  AOI21_X1 u2_u9_u0_U44 (.A( u2_u9_u0_n144 ) , .B2( u2_u9_u0_n145 ) , .B1( u2_u9_u0_n146 ) , .ZN( u2_u9_u0_n154 ) );
  AOI21_X1 u2_u9_u0_U45 (.B2( u2_u9_u0_n150 ) , .B1( u2_u9_u0_n151 ) , .ZN( u2_u9_u0_n152 ) , .A( u2_u9_u0_n158 ) );
  AOI21_X1 u2_u9_u0_U46 (.A( u2_u9_u0_n147 ) , .B2( u2_u9_u0_n148 ) , .B1( u2_u9_u0_n149 ) , .ZN( u2_u9_u0_n153 ) );
  AOI21_X1 u2_u9_u0_U47 (.B1( u2_u9_u0_n103 ) , .ZN( u2_u9_u0_n132 ) , .A( u2_u9_u0_n165 ) , .B2( u2_u9_u0_n93 ) );
  INV_X1 u2_u9_u0_U48 (.A( u2_u9_u0_n142 ) , .ZN( u2_u9_u0_n165 ) );
  INV_X1 u2_u9_u0_U49 (.ZN( u2_u9_u0_n171 ) , .A( u2_u9_u0_n99 ) );
  AOI21_X1 u2_u9_u0_U5 (.B2( u2_u9_u0_n131 ) , .ZN( u2_u9_u0_n134 ) , .B1( u2_u9_u0_n151 ) , .A( u2_u9_u0_n158 ) );
  OAI211_X1 u2_u9_u0_U50 (.C2( u2_u9_u0_n140 ) , .C1( u2_u9_u0_n161 ) , .A( u2_u9_u0_n169 ) , .B( u2_u9_u0_n98 ) , .ZN( u2_u9_u0_n99 ) );
  INV_X1 u2_u9_u0_U51 (.ZN( u2_u9_u0_n169 ) , .A( u2_u9_u0_n91 ) );
  AOI211_X1 u2_u9_u0_U52 (.C1( u2_u9_u0_n118 ) , .A( u2_u9_u0_n123 ) , .B( u2_u9_u0_n96 ) , .C2( u2_u9_u0_n97 ) , .ZN( u2_u9_u0_n98 ) );
  NOR2_X1 u2_u9_u0_U53 (.A2( u2_u9_X_2 ) , .ZN( u2_u9_u0_n103 ) , .A1( u2_u9_u0_n164 ) );
  NOR2_X1 u2_u9_u0_U54 (.A2( u2_u9_X_4 ) , .A1( u2_u9_X_5 ) , .ZN( u2_u9_u0_n118 ) );
  NOR2_X1 u2_u9_u0_U55 (.A2( u2_u9_X_1 ) , .A1( u2_u9_X_2 ) , .ZN( u2_u9_u0_n92 ) );
  NOR2_X1 u2_u9_u0_U56 (.A2( u2_u9_X_1 ) , .ZN( u2_u9_u0_n101 ) , .A1( u2_u9_u0_n163 ) );
  NOR2_X1 u2_u9_u0_U57 (.A2( u2_u9_X_3 ) , .A1( u2_u9_X_6 ) , .ZN( u2_u9_u0_n94 ) );
  NOR2_X1 u2_u9_u0_U58 (.A2( u2_u9_X_6 ) , .ZN( u2_u9_u0_n100 ) , .A1( u2_u9_u0_n162 ) );
  NAND2_X1 u2_u9_u0_U59 (.A2( u2_u9_X_4 ) , .A1( u2_u9_X_5 ) , .ZN( u2_u9_u0_n144 ) );
  NOR2_X1 u2_u9_u0_U6 (.A1( u2_u9_u0_n108 ) , .ZN( u2_u9_u0_n123 ) , .A2( u2_u9_u0_n158 ) );
  NOR2_X1 u2_u9_u0_U60 (.A2( u2_u9_X_5 ) , .ZN( u2_u9_u0_n136 ) , .A1( u2_u9_u0_n159 ) );
  NAND2_X1 u2_u9_u0_U61 (.A1( u2_u9_X_5 ) , .ZN( u2_u9_u0_n138 ) , .A2( u2_u9_u0_n159 ) );
  AND2_X1 u2_u9_u0_U62 (.A2( u2_u9_X_3 ) , .A1( u2_u9_X_6 ) , .ZN( u2_u9_u0_n102 ) );
  AND2_X1 u2_u9_u0_U63 (.A1( u2_u9_X_6 ) , .A2( u2_u9_u0_n162 ) , .ZN( u2_u9_u0_n93 ) );
  INV_X1 u2_u9_u0_U64 (.A( u2_u9_X_4 ) , .ZN( u2_u9_u0_n159 ) );
  INV_X1 u2_u9_u0_U65 (.A( u2_u9_X_1 ) , .ZN( u2_u9_u0_n164 ) );
  INV_X1 u2_u9_u0_U66 (.A( u2_u9_X_2 ) , .ZN( u2_u9_u0_n163 ) );
  INV_X1 u2_u9_u0_U67 (.A( u2_u9_X_3 ) , .ZN( u2_u9_u0_n162 ) );
  INV_X1 u2_u9_u0_U68 (.A( u2_u9_u0_n126 ) , .ZN( u2_u9_u0_n168 ) );
  AOI211_X1 u2_u9_u0_U69 (.B( u2_u9_u0_n133 ) , .A( u2_u9_u0_n134 ) , .C2( u2_u9_u0_n135 ) , .C1( u2_u9_u0_n136 ) , .ZN( u2_u9_u0_n137 ) );
  OAI21_X1 u2_u9_u0_U7 (.B1( u2_u9_u0_n150 ) , .B2( u2_u9_u0_n158 ) , .A( u2_u9_u0_n172 ) , .ZN( u2_u9_u0_n89 ) );
  OR4_X1 u2_u9_u0_U70 (.ZN( u2_out9_17 ) , .A4( u2_u9_u0_n122 ) , .A2( u2_u9_u0_n123 ) , .A1( u2_u9_u0_n124 ) , .A3( u2_u9_u0_n170 ) );
  AOI21_X1 u2_u9_u0_U71 (.B2( u2_u9_u0_n107 ) , .ZN( u2_u9_u0_n124 ) , .B1( u2_u9_u0_n128 ) , .A( u2_u9_u0_n161 ) );
  INV_X1 u2_u9_u0_U72 (.A( u2_u9_u0_n111 ) , .ZN( u2_u9_u0_n170 ) );
  OR4_X1 u2_u9_u0_U73 (.ZN( u2_out9_31 ) , .A4( u2_u9_u0_n155 ) , .A2( u2_u9_u0_n156 ) , .A1( u2_u9_u0_n157 ) , .A3( u2_u9_u0_n173 ) );
  AOI21_X1 u2_u9_u0_U74 (.A( u2_u9_u0_n138 ) , .B2( u2_u9_u0_n139 ) , .B1( u2_u9_u0_n140 ) , .ZN( u2_u9_u0_n157 ) );
  AOI21_X1 u2_u9_u0_U75 (.B2( u2_u9_u0_n141 ) , .B1( u2_u9_u0_n142 ) , .ZN( u2_u9_u0_n156 ) , .A( u2_u9_u0_n161 ) );
  INV_X1 u2_u9_u0_U76 (.ZN( u2_u9_u0_n174 ) , .A( u2_u9_u0_n89 ) );
  AOI211_X1 u2_u9_u0_U77 (.B( u2_u9_u0_n104 ) , .A( u2_u9_u0_n105 ) , .ZN( u2_u9_u0_n106 ) , .C2( u2_u9_u0_n113 ) , .C1( u2_u9_u0_n160 ) );
  OAI221_X1 u2_u9_u0_U78 (.C1( u2_u9_u0_n121 ) , .ZN( u2_u9_u0_n122 ) , .B2( u2_u9_u0_n127 ) , .A( u2_u9_u0_n143 ) , .B1( u2_u9_u0_n144 ) , .C2( u2_u9_u0_n147 ) );
  NOR2_X1 u2_u9_u0_U79 (.A1( u2_u9_u0_n120 ) , .ZN( u2_u9_u0_n143 ) , .A2( u2_u9_u0_n167 ) );
  AND2_X1 u2_u9_u0_U8 (.A1( u2_u9_u0_n114 ) , .A2( u2_u9_u0_n121 ) , .ZN( u2_u9_u0_n146 ) );
  AOI21_X1 u2_u9_u0_U80 (.B1( u2_u9_u0_n132 ) , .ZN( u2_u9_u0_n133 ) , .A( u2_u9_u0_n144 ) , .B2( u2_u9_u0_n166 ) );
  OAI22_X1 u2_u9_u0_U81 (.ZN( u2_u9_u0_n105 ) , .A2( u2_u9_u0_n132 ) , .B1( u2_u9_u0_n146 ) , .A1( u2_u9_u0_n147 ) , .B2( u2_u9_u0_n161 ) );
  NAND2_X1 u2_u9_u0_U82 (.ZN( u2_u9_u0_n110 ) , .A2( u2_u9_u0_n132 ) , .A1( u2_u9_u0_n145 ) );
  INV_X1 u2_u9_u0_U83 (.A( u2_u9_u0_n119 ) , .ZN( u2_u9_u0_n167 ) );
  NAND2_X1 u2_u9_u0_U84 (.ZN( u2_u9_u0_n148 ) , .A1( u2_u9_u0_n93 ) , .A2( u2_u9_u0_n95 ) );
  NAND2_X1 u2_u9_u0_U85 (.A1( u2_u9_u0_n100 ) , .ZN( u2_u9_u0_n129 ) , .A2( u2_u9_u0_n95 ) );
  NAND2_X1 u2_u9_u0_U86 (.A1( u2_u9_u0_n102 ) , .ZN( u2_u9_u0_n128 ) , .A2( u2_u9_u0_n95 ) );
  NAND2_X1 u2_u9_u0_U87 (.ZN( u2_u9_u0_n142 ) , .A1( u2_u9_u0_n94 ) , .A2( u2_u9_u0_n95 ) );
  NAND3_X1 u2_u9_u0_U88 (.ZN( u2_out9_23 ) , .A3( u2_u9_u0_n137 ) , .A1( u2_u9_u0_n168 ) , .A2( u2_u9_u0_n171 ) );
  NAND3_X1 u2_u9_u0_U89 (.A3( u2_u9_u0_n127 ) , .A2( u2_u9_u0_n128 ) , .ZN( u2_u9_u0_n135 ) , .A1( u2_u9_u0_n150 ) );
  AND2_X1 u2_u9_u0_U9 (.A1( u2_u9_u0_n131 ) , .ZN( u2_u9_u0_n141 ) , .A2( u2_u9_u0_n150 ) );
  NAND3_X1 u2_u9_u0_U90 (.ZN( u2_u9_u0_n117 ) , .A3( u2_u9_u0_n132 ) , .A2( u2_u9_u0_n139 ) , .A1( u2_u9_u0_n148 ) );
  NAND3_X1 u2_u9_u0_U91 (.ZN( u2_u9_u0_n109 ) , .A2( u2_u9_u0_n114 ) , .A3( u2_u9_u0_n140 ) , .A1( u2_u9_u0_n149 ) );
  NAND3_X1 u2_u9_u0_U92 (.ZN( u2_out9_9 ) , .A3( u2_u9_u0_n106 ) , .A2( u2_u9_u0_n171 ) , .A1( u2_u9_u0_n174 ) );
  NAND3_X1 u2_u9_u0_U93 (.A2( u2_u9_u0_n128 ) , .A1( u2_u9_u0_n132 ) , .A3( u2_u9_u0_n146 ) , .ZN( u2_u9_u0_n97 ) );
  NOR2_X1 u2_u9_u1_U10 (.A1( u2_u9_u1_n112 ) , .A2( u2_u9_u1_n116 ) , .ZN( u2_u9_u1_n118 ) );
  NAND3_X1 u2_u9_u1_U100 (.ZN( u2_u9_u1_n113 ) , .A1( u2_u9_u1_n120 ) , .A3( u2_u9_u1_n133 ) , .A2( u2_u9_u1_n155 ) );
  OAI21_X1 u2_u9_u1_U11 (.ZN( u2_u9_u1_n101 ) , .B1( u2_u9_u1_n141 ) , .A( u2_u9_u1_n146 ) , .B2( u2_u9_u1_n183 ) );
  AOI21_X1 u2_u9_u1_U12 (.B2( u2_u9_u1_n155 ) , .B1( u2_u9_u1_n156 ) , .ZN( u2_u9_u1_n157 ) , .A( u2_u9_u1_n174 ) );
  NAND2_X1 u2_u9_u1_U13 (.ZN( u2_u9_u1_n140 ) , .A2( u2_u9_u1_n150 ) , .A1( u2_u9_u1_n155 ) );
  NAND2_X1 u2_u9_u1_U14 (.A1( u2_u9_u1_n131 ) , .ZN( u2_u9_u1_n147 ) , .A2( u2_u9_u1_n153 ) );
  INV_X1 u2_u9_u1_U15 (.A( u2_u9_u1_n139 ) , .ZN( u2_u9_u1_n174 ) );
  OR4_X1 u2_u9_u1_U16 (.A4( u2_u9_u1_n106 ) , .A3( u2_u9_u1_n107 ) , .ZN( u2_u9_u1_n108 ) , .A1( u2_u9_u1_n117 ) , .A2( u2_u9_u1_n184 ) );
  AOI21_X1 u2_u9_u1_U17 (.ZN( u2_u9_u1_n106 ) , .A( u2_u9_u1_n112 ) , .B1( u2_u9_u1_n154 ) , .B2( u2_u9_u1_n156 ) );
  AOI21_X1 u2_u9_u1_U18 (.ZN( u2_u9_u1_n107 ) , .B1( u2_u9_u1_n134 ) , .B2( u2_u9_u1_n149 ) , .A( u2_u9_u1_n174 ) );
  INV_X1 u2_u9_u1_U19 (.A( u2_u9_u1_n101 ) , .ZN( u2_u9_u1_n184 ) );
  INV_X1 u2_u9_u1_U20 (.A( u2_u9_u1_n112 ) , .ZN( u2_u9_u1_n171 ) );
  NAND2_X1 u2_u9_u1_U21 (.ZN( u2_u9_u1_n141 ) , .A1( u2_u9_u1_n153 ) , .A2( u2_u9_u1_n156 ) );
  AND2_X1 u2_u9_u1_U22 (.A1( u2_u9_u1_n123 ) , .ZN( u2_u9_u1_n134 ) , .A2( u2_u9_u1_n161 ) );
  NAND2_X1 u2_u9_u1_U23 (.A2( u2_u9_u1_n115 ) , .A1( u2_u9_u1_n116 ) , .ZN( u2_u9_u1_n148 ) );
  NAND2_X1 u2_u9_u1_U24 (.A2( u2_u9_u1_n133 ) , .A1( u2_u9_u1_n135 ) , .ZN( u2_u9_u1_n159 ) );
  NAND2_X1 u2_u9_u1_U25 (.A2( u2_u9_u1_n115 ) , .A1( u2_u9_u1_n120 ) , .ZN( u2_u9_u1_n132 ) );
  INV_X1 u2_u9_u1_U26 (.A( u2_u9_u1_n154 ) , .ZN( u2_u9_u1_n178 ) );
  INV_X1 u2_u9_u1_U27 (.A( u2_u9_u1_n151 ) , .ZN( u2_u9_u1_n183 ) );
  AND2_X1 u2_u9_u1_U28 (.A1( u2_u9_u1_n129 ) , .A2( u2_u9_u1_n133 ) , .ZN( u2_u9_u1_n149 ) );
  INV_X1 u2_u9_u1_U29 (.A( u2_u9_u1_n131 ) , .ZN( u2_u9_u1_n180 ) );
  INV_X1 u2_u9_u1_U3 (.A( u2_u9_u1_n159 ) , .ZN( u2_u9_u1_n182 ) );
  OAI221_X1 u2_u9_u1_U30 (.A( u2_u9_u1_n119 ) , .C2( u2_u9_u1_n129 ) , .ZN( u2_u9_u1_n138 ) , .B2( u2_u9_u1_n152 ) , .C1( u2_u9_u1_n174 ) , .B1( u2_u9_u1_n187 ) );
  INV_X1 u2_u9_u1_U31 (.A( u2_u9_u1_n148 ) , .ZN( u2_u9_u1_n187 ) );
  AOI211_X1 u2_u9_u1_U32 (.B( u2_u9_u1_n117 ) , .A( u2_u9_u1_n118 ) , .ZN( u2_u9_u1_n119 ) , .C2( u2_u9_u1_n146 ) , .C1( u2_u9_u1_n159 ) );
  NOR2_X1 u2_u9_u1_U33 (.A1( u2_u9_u1_n168 ) , .A2( u2_u9_u1_n176 ) , .ZN( u2_u9_u1_n98 ) );
  AOI211_X1 u2_u9_u1_U34 (.B( u2_u9_u1_n162 ) , .A( u2_u9_u1_n163 ) , .C2( u2_u9_u1_n164 ) , .ZN( u2_u9_u1_n165 ) , .C1( u2_u9_u1_n171 ) );
  AOI21_X1 u2_u9_u1_U35 (.A( u2_u9_u1_n160 ) , .B2( u2_u9_u1_n161 ) , .ZN( u2_u9_u1_n162 ) , .B1( u2_u9_u1_n182 ) );
  OR2_X1 u2_u9_u1_U36 (.A2( u2_u9_u1_n157 ) , .A1( u2_u9_u1_n158 ) , .ZN( u2_u9_u1_n163 ) );
  NAND2_X1 u2_u9_u1_U37 (.A1( u2_u9_u1_n128 ) , .ZN( u2_u9_u1_n146 ) , .A2( u2_u9_u1_n160 ) );
  NAND2_X1 u2_u9_u1_U38 (.A2( u2_u9_u1_n112 ) , .ZN( u2_u9_u1_n139 ) , .A1( u2_u9_u1_n152 ) );
  NAND2_X1 u2_u9_u1_U39 (.A1( u2_u9_u1_n105 ) , .ZN( u2_u9_u1_n156 ) , .A2( u2_u9_u1_n99 ) );
  AOI221_X1 u2_u9_u1_U4 (.A( u2_u9_u1_n138 ) , .C2( u2_u9_u1_n139 ) , .C1( u2_u9_u1_n140 ) , .B2( u2_u9_u1_n141 ) , .ZN( u2_u9_u1_n142 ) , .B1( u2_u9_u1_n175 ) );
  AOI221_X1 u2_u9_u1_U40 (.B1( u2_u9_u1_n140 ) , .ZN( u2_u9_u1_n167 ) , .B2( u2_u9_u1_n172 ) , .C2( u2_u9_u1_n175 ) , .C1( u2_u9_u1_n178 ) , .A( u2_u9_u1_n188 ) );
  INV_X1 u2_u9_u1_U41 (.ZN( u2_u9_u1_n188 ) , .A( u2_u9_u1_n97 ) );
  AOI211_X1 u2_u9_u1_U42 (.A( u2_u9_u1_n118 ) , .C1( u2_u9_u1_n132 ) , .C2( u2_u9_u1_n139 ) , .B( u2_u9_u1_n96 ) , .ZN( u2_u9_u1_n97 ) );
  AOI21_X1 u2_u9_u1_U43 (.B2( u2_u9_u1_n121 ) , .B1( u2_u9_u1_n135 ) , .A( u2_u9_u1_n152 ) , .ZN( u2_u9_u1_n96 ) );
  NOR2_X1 u2_u9_u1_U44 (.ZN( u2_u9_u1_n117 ) , .A1( u2_u9_u1_n121 ) , .A2( u2_u9_u1_n160 ) );
  OAI21_X1 u2_u9_u1_U45 (.B2( u2_u9_u1_n123 ) , .ZN( u2_u9_u1_n145 ) , .B1( u2_u9_u1_n160 ) , .A( u2_u9_u1_n185 ) );
  INV_X1 u2_u9_u1_U46 (.A( u2_u9_u1_n122 ) , .ZN( u2_u9_u1_n185 ) );
  AOI21_X1 u2_u9_u1_U47 (.B2( u2_u9_u1_n120 ) , .B1( u2_u9_u1_n121 ) , .ZN( u2_u9_u1_n122 ) , .A( u2_u9_u1_n128 ) );
  AOI21_X1 u2_u9_u1_U48 (.A( u2_u9_u1_n128 ) , .B2( u2_u9_u1_n129 ) , .ZN( u2_u9_u1_n130 ) , .B1( u2_u9_u1_n150 ) );
  NAND2_X1 u2_u9_u1_U49 (.ZN( u2_u9_u1_n112 ) , .A1( u2_u9_u1_n169 ) , .A2( u2_u9_u1_n170 ) );
  AOI211_X1 u2_u9_u1_U5 (.ZN( u2_u9_u1_n124 ) , .A( u2_u9_u1_n138 ) , .C2( u2_u9_u1_n139 ) , .B( u2_u9_u1_n145 ) , .C1( u2_u9_u1_n147 ) );
  NAND2_X1 u2_u9_u1_U50 (.ZN( u2_u9_u1_n129 ) , .A2( u2_u9_u1_n95 ) , .A1( u2_u9_u1_n98 ) );
  NAND2_X1 u2_u9_u1_U51 (.A1( u2_u9_u1_n102 ) , .ZN( u2_u9_u1_n154 ) , .A2( u2_u9_u1_n99 ) );
  NAND2_X1 u2_u9_u1_U52 (.A2( u2_u9_u1_n100 ) , .ZN( u2_u9_u1_n135 ) , .A1( u2_u9_u1_n99 ) );
  AOI21_X1 u2_u9_u1_U53 (.A( u2_u9_u1_n152 ) , .B2( u2_u9_u1_n153 ) , .B1( u2_u9_u1_n154 ) , .ZN( u2_u9_u1_n158 ) );
  INV_X1 u2_u9_u1_U54 (.A( u2_u9_u1_n160 ) , .ZN( u2_u9_u1_n175 ) );
  NAND2_X1 u2_u9_u1_U55 (.A1( u2_u9_u1_n100 ) , .ZN( u2_u9_u1_n116 ) , .A2( u2_u9_u1_n95 ) );
  NAND2_X1 u2_u9_u1_U56 (.A1( u2_u9_u1_n102 ) , .ZN( u2_u9_u1_n131 ) , .A2( u2_u9_u1_n95 ) );
  NAND2_X1 u2_u9_u1_U57 (.A2( u2_u9_u1_n104 ) , .ZN( u2_u9_u1_n121 ) , .A1( u2_u9_u1_n98 ) );
  NAND2_X1 u2_u9_u1_U58 (.A1( u2_u9_u1_n103 ) , .ZN( u2_u9_u1_n153 ) , .A2( u2_u9_u1_n98 ) );
  NAND2_X1 u2_u9_u1_U59 (.A2( u2_u9_u1_n104 ) , .A1( u2_u9_u1_n105 ) , .ZN( u2_u9_u1_n133 ) );
  AOI22_X1 u2_u9_u1_U6 (.B2( u2_u9_u1_n136 ) , .A2( u2_u9_u1_n137 ) , .ZN( u2_u9_u1_n143 ) , .A1( u2_u9_u1_n171 ) , .B1( u2_u9_u1_n173 ) );
  NAND2_X1 u2_u9_u1_U60 (.ZN( u2_u9_u1_n150 ) , .A2( u2_u9_u1_n98 ) , .A1( u2_u9_u1_n99 ) );
  NAND2_X1 u2_u9_u1_U61 (.A1( u2_u9_u1_n105 ) , .ZN( u2_u9_u1_n155 ) , .A2( u2_u9_u1_n95 ) );
  OAI21_X1 u2_u9_u1_U62 (.ZN( u2_u9_u1_n109 ) , .B1( u2_u9_u1_n129 ) , .B2( u2_u9_u1_n160 ) , .A( u2_u9_u1_n167 ) );
  NAND2_X1 u2_u9_u1_U63 (.A2( u2_u9_u1_n100 ) , .A1( u2_u9_u1_n103 ) , .ZN( u2_u9_u1_n120 ) );
  NAND2_X1 u2_u9_u1_U64 (.A1( u2_u9_u1_n102 ) , .A2( u2_u9_u1_n104 ) , .ZN( u2_u9_u1_n115 ) );
  NAND2_X1 u2_u9_u1_U65 (.A2( u2_u9_u1_n100 ) , .A1( u2_u9_u1_n104 ) , .ZN( u2_u9_u1_n151 ) );
  NAND2_X1 u2_u9_u1_U66 (.A2( u2_u9_u1_n103 ) , .A1( u2_u9_u1_n105 ) , .ZN( u2_u9_u1_n161 ) );
  INV_X1 u2_u9_u1_U67 (.A( u2_u9_u1_n152 ) , .ZN( u2_u9_u1_n173 ) );
  INV_X1 u2_u9_u1_U68 (.A( u2_u9_u1_n128 ) , .ZN( u2_u9_u1_n172 ) );
  NAND2_X1 u2_u9_u1_U69 (.A2( u2_u9_u1_n102 ) , .A1( u2_u9_u1_n103 ) , .ZN( u2_u9_u1_n123 ) );
  INV_X1 u2_u9_u1_U7 (.A( u2_u9_u1_n147 ) , .ZN( u2_u9_u1_n181 ) );
  NOR2_X1 u2_u9_u1_U70 (.A2( u2_u9_X_7 ) , .A1( u2_u9_X_8 ) , .ZN( u2_u9_u1_n95 ) );
  NOR2_X1 u2_u9_u1_U71 (.A1( u2_u9_X_12 ) , .A2( u2_u9_X_9 ) , .ZN( u2_u9_u1_n100 ) );
  NOR2_X1 u2_u9_u1_U72 (.A2( u2_u9_X_8 ) , .A1( u2_u9_u1_n177 ) , .ZN( u2_u9_u1_n99 ) );
  NOR2_X1 u2_u9_u1_U73 (.A2( u2_u9_X_12 ) , .ZN( u2_u9_u1_n102 ) , .A1( u2_u9_u1_n176 ) );
  NOR2_X1 u2_u9_u1_U74 (.A2( u2_u9_X_9 ) , .ZN( u2_u9_u1_n105 ) , .A1( u2_u9_u1_n168 ) );
  NAND2_X1 u2_u9_u1_U75 (.A1( u2_u9_X_10 ) , .ZN( u2_u9_u1_n160 ) , .A2( u2_u9_u1_n169 ) );
  NAND2_X1 u2_u9_u1_U76 (.A2( u2_u9_X_10 ) , .A1( u2_u9_X_11 ) , .ZN( u2_u9_u1_n152 ) );
  NAND2_X1 u2_u9_u1_U77 (.A1( u2_u9_X_11 ) , .ZN( u2_u9_u1_n128 ) , .A2( u2_u9_u1_n170 ) );
  AND2_X1 u2_u9_u1_U78 (.A2( u2_u9_X_7 ) , .A1( u2_u9_X_8 ) , .ZN( u2_u9_u1_n104 ) );
  AND2_X1 u2_u9_u1_U79 (.A1( u2_u9_X_8 ) , .ZN( u2_u9_u1_n103 ) , .A2( u2_u9_u1_n177 ) );
  AOI22_X1 u2_u9_u1_U8 (.B2( u2_u9_u1_n113 ) , .A2( u2_u9_u1_n114 ) , .ZN( u2_u9_u1_n125 ) , .A1( u2_u9_u1_n171 ) , .B1( u2_u9_u1_n173 ) );
  INV_X1 u2_u9_u1_U80 (.A( u2_u9_X_10 ) , .ZN( u2_u9_u1_n170 ) );
  INV_X1 u2_u9_u1_U81 (.A( u2_u9_X_9 ) , .ZN( u2_u9_u1_n176 ) );
  INV_X1 u2_u9_u1_U82 (.A( u2_u9_X_11 ) , .ZN( u2_u9_u1_n169 ) );
  INV_X1 u2_u9_u1_U83 (.A( u2_u9_X_12 ) , .ZN( u2_u9_u1_n168 ) );
  INV_X1 u2_u9_u1_U84 (.A( u2_u9_X_7 ) , .ZN( u2_u9_u1_n177 ) );
  NAND4_X1 u2_u9_u1_U85 (.ZN( u2_out9_28 ) , .A4( u2_u9_u1_n124 ) , .A3( u2_u9_u1_n125 ) , .A2( u2_u9_u1_n126 ) , .A1( u2_u9_u1_n127 ) );
  OAI21_X1 u2_u9_u1_U86 (.ZN( u2_u9_u1_n127 ) , .B2( u2_u9_u1_n139 ) , .B1( u2_u9_u1_n175 ) , .A( u2_u9_u1_n183 ) );
  OAI21_X1 u2_u9_u1_U87 (.ZN( u2_u9_u1_n126 ) , .B2( u2_u9_u1_n140 ) , .A( u2_u9_u1_n146 ) , .B1( u2_u9_u1_n178 ) );
  NAND4_X1 u2_u9_u1_U88 (.ZN( u2_out9_18 ) , .A4( u2_u9_u1_n165 ) , .A3( u2_u9_u1_n166 ) , .A1( u2_u9_u1_n167 ) , .A2( u2_u9_u1_n186 ) );
  AOI22_X1 u2_u9_u1_U89 (.B2( u2_u9_u1_n146 ) , .B1( u2_u9_u1_n147 ) , .A2( u2_u9_u1_n148 ) , .ZN( u2_u9_u1_n166 ) , .A1( u2_u9_u1_n172 ) );
  NAND2_X1 u2_u9_u1_U9 (.ZN( u2_u9_u1_n114 ) , .A1( u2_u9_u1_n134 ) , .A2( u2_u9_u1_n156 ) );
  INV_X1 u2_u9_u1_U90 (.A( u2_u9_u1_n145 ) , .ZN( u2_u9_u1_n186 ) );
  NAND4_X1 u2_u9_u1_U91 (.ZN( u2_out9_2 ) , .A4( u2_u9_u1_n142 ) , .A3( u2_u9_u1_n143 ) , .A2( u2_u9_u1_n144 ) , .A1( u2_u9_u1_n179 ) );
  OAI21_X1 u2_u9_u1_U92 (.B2( u2_u9_u1_n132 ) , .ZN( u2_u9_u1_n144 ) , .A( u2_u9_u1_n146 ) , .B1( u2_u9_u1_n180 ) );
  INV_X1 u2_u9_u1_U93 (.A( u2_u9_u1_n130 ) , .ZN( u2_u9_u1_n179 ) );
  OR4_X1 u2_u9_u1_U94 (.ZN( u2_out9_13 ) , .A4( u2_u9_u1_n108 ) , .A3( u2_u9_u1_n109 ) , .A2( u2_u9_u1_n110 ) , .A1( u2_u9_u1_n111 ) );
  AOI21_X1 u2_u9_u1_U95 (.ZN( u2_u9_u1_n110 ) , .A( u2_u9_u1_n116 ) , .B1( u2_u9_u1_n152 ) , .B2( u2_u9_u1_n160 ) );
  AOI21_X1 u2_u9_u1_U96 (.ZN( u2_u9_u1_n111 ) , .A( u2_u9_u1_n128 ) , .B2( u2_u9_u1_n131 ) , .B1( u2_u9_u1_n135 ) );
  NAND3_X1 u2_u9_u1_U97 (.A3( u2_u9_u1_n149 ) , .A2( u2_u9_u1_n150 ) , .A1( u2_u9_u1_n151 ) , .ZN( u2_u9_u1_n164 ) );
  NAND3_X1 u2_u9_u1_U98 (.A3( u2_u9_u1_n134 ) , .A2( u2_u9_u1_n135 ) , .ZN( u2_u9_u1_n136 ) , .A1( u2_u9_u1_n151 ) );
  NAND3_X1 u2_u9_u1_U99 (.A1( u2_u9_u1_n133 ) , .ZN( u2_u9_u1_n137 ) , .A2( u2_u9_u1_n154 ) , .A3( u2_u9_u1_n181 ) );
  OAI22_X1 u2_u9_u2_U10 (.B1( u2_u9_u2_n151 ) , .A2( u2_u9_u2_n152 ) , .A1( u2_u9_u2_n153 ) , .ZN( u2_u9_u2_n160 ) , .B2( u2_u9_u2_n168 ) );
  NAND3_X1 u2_u9_u2_U100 (.A2( u2_u9_u2_n100 ) , .A1( u2_u9_u2_n104 ) , .A3( u2_u9_u2_n138 ) , .ZN( u2_u9_u2_n98 ) );
  NOR3_X1 u2_u9_u2_U11 (.A1( u2_u9_u2_n150 ) , .ZN( u2_u9_u2_n151 ) , .A3( u2_u9_u2_n175 ) , .A2( u2_u9_u2_n188 ) );
  AOI21_X1 u2_u9_u2_U12 (.B2( u2_u9_u2_n123 ) , .ZN( u2_u9_u2_n125 ) , .A( u2_u9_u2_n171 ) , .B1( u2_u9_u2_n184 ) );
  INV_X1 u2_u9_u2_U13 (.A( u2_u9_u2_n150 ) , .ZN( u2_u9_u2_n184 ) );
  AOI21_X1 u2_u9_u2_U14 (.ZN( u2_u9_u2_n144 ) , .B2( u2_u9_u2_n155 ) , .A( u2_u9_u2_n172 ) , .B1( u2_u9_u2_n185 ) );
  AOI21_X1 u2_u9_u2_U15 (.B2( u2_u9_u2_n143 ) , .ZN( u2_u9_u2_n145 ) , .B1( u2_u9_u2_n152 ) , .A( u2_u9_u2_n171 ) );
  INV_X1 u2_u9_u2_U16 (.A( u2_u9_u2_n156 ) , .ZN( u2_u9_u2_n171 ) );
  INV_X1 u2_u9_u2_U17 (.A( u2_u9_u2_n120 ) , .ZN( u2_u9_u2_n188 ) );
  NAND2_X1 u2_u9_u2_U18 (.A2( u2_u9_u2_n122 ) , .ZN( u2_u9_u2_n150 ) , .A1( u2_u9_u2_n152 ) );
  INV_X1 u2_u9_u2_U19 (.A( u2_u9_u2_n153 ) , .ZN( u2_u9_u2_n170 ) );
  INV_X1 u2_u9_u2_U20 (.A( u2_u9_u2_n137 ) , .ZN( u2_u9_u2_n173 ) );
  NAND2_X1 u2_u9_u2_U21 (.A1( u2_u9_u2_n132 ) , .A2( u2_u9_u2_n139 ) , .ZN( u2_u9_u2_n157 ) );
  INV_X1 u2_u9_u2_U22 (.A( u2_u9_u2_n113 ) , .ZN( u2_u9_u2_n178 ) );
  INV_X1 u2_u9_u2_U23 (.A( u2_u9_u2_n139 ) , .ZN( u2_u9_u2_n175 ) );
  INV_X1 u2_u9_u2_U24 (.A( u2_u9_u2_n155 ) , .ZN( u2_u9_u2_n181 ) );
  INV_X1 u2_u9_u2_U25 (.A( u2_u9_u2_n119 ) , .ZN( u2_u9_u2_n177 ) );
  INV_X1 u2_u9_u2_U26 (.A( u2_u9_u2_n116 ) , .ZN( u2_u9_u2_n180 ) );
  INV_X1 u2_u9_u2_U27 (.A( u2_u9_u2_n131 ) , .ZN( u2_u9_u2_n179 ) );
  INV_X1 u2_u9_u2_U28 (.A( u2_u9_u2_n154 ) , .ZN( u2_u9_u2_n176 ) );
  NAND2_X1 u2_u9_u2_U29 (.A2( u2_u9_u2_n116 ) , .A1( u2_u9_u2_n117 ) , .ZN( u2_u9_u2_n118 ) );
  NOR2_X1 u2_u9_u2_U3 (.ZN( u2_u9_u2_n121 ) , .A2( u2_u9_u2_n177 ) , .A1( u2_u9_u2_n180 ) );
  INV_X1 u2_u9_u2_U30 (.A( u2_u9_u2_n132 ) , .ZN( u2_u9_u2_n182 ) );
  INV_X1 u2_u9_u2_U31 (.A( u2_u9_u2_n158 ) , .ZN( u2_u9_u2_n183 ) );
  OAI21_X1 u2_u9_u2_U32 (.A( u2_u9_u2_n156 ) , .B1( u2_u9_u2_n157 ) , .ZN( u2_u9_u2_n158 ) , .B2( u2_u9_u2_n179 ) );
  NOR2_X1 u2_u9_u2_U33 (.ZN( u2_u9_u2_n156 ) , .A1( u2_u9_u2_n166 ) , .A2( u2_u9_u2_n169 ) );
  NOR2_X1 u2_u9_u2_U34 (.A2( u2_u9_u2_n114 ) , .ZN( u2_u9_u2_n137 ) , .A1( u2_u9_u2_n140 ) );
  NOR2_X1 u2_u9_u2_U35 (.A2( u2_u9_u2_n138 ) , .ZN( u2_u9_u2_n153 ) , .A1( u2_u9_u2_n156 ) );
  AOI211_X1 u2_u9_u2_U36 (.ZN( u2_u9_u2_n130 ) , .C1( u2_u9_u2_n138 ) , .C2( u2_u9_u2_n179 ) , .B( u2_u9_u2_n96 ) , .A( u2_u9_u2_n97 ) );
  OAI22_X1 u2_u9_u2_U37 (.B1( u2_u9_u2_n133 ) , .A2( u2_u9_u2_n137 ) , .A1( u2_u9_u2_n152 ) , .B2( u2_u9_u2_n168 ) , .ZN( u2_u9_u2_n97 ) );
  OAI221_X1 u2_u9_u2_U38 (.B1( u2_u9_u2_n113 ) , .C1( u2_u9_u2_n132 ) , .A( u2_u9_u2_n149 ) , .B2( u2_u9_u2_n171 ) , .C2( u2_u9_u2_n172 ) , .ZN( u2_u9_u2_n96 ) );
  OAI221_X1 u2_u9_u2_U39 (.A( u2_u9_u2_n115 ) , .C2( u2_u9_u2_n123 ) , .B2( u2_u9_u2_n143 ) , .B1( u2_u9_u2_n153 ) , .ZN( u2_u9_u2_n163 ) , .C1( u2_u9_u2_n168 ) );
  INV_X1 u2_u9_u2_U4 (.A( u2_u9_u2_n134 ) , .ZN( u2_u9_u2_n185 ) );
  OAI21_X1 u2_u9_u2_U40 (.A( u2_u9_u2_n114 ) , .ZN( u2_u9_u2_n115 ) , .B1( u2_u9_u2_n176 ) , .B2( u2_u9_u2_n178 ) );
  OAI221_X1 u2_u9_u2_U41 (.A( u2_u9_u2_n135 ) , .B2( u2_u9_u2_n136 ) , .B1( u2_u9_u2_n137 ) , .ZN( u2_u9_u2_n162 ) , .C2( u2_u9_u2_n167 ) , .C1( u2_u9_u2_n185 ) );
  AND3_X1 u2_u9_u2_U42 (.A3( u2_u9_u2_n131 ) , .A2( u2_u9_u2_n132 ) , .A1( u2_u9_u2_n133 ) , .ZN( u2_u9_u2_n136 ) );
  AOI22_X1 u2_u9_u2_U43 (.ZN( u2_u9_u2_n135 ) , .B1( u2_u9_u2_n140 ) , .A1( u2_u9_u2_n156 ) , .B2( u2_u9_u2_n180 ) , .A2( u2_u9_u2_n188 ) );
  AOI21_X1 u2_u9_u2_U44 (.ZN( u2_u9_u2_n149 ) , .B1( u2_u9_u2_n173 ) , .B2( u2_u9_u2_n188 ) , .A( u2_u9_u2_n95 ) );
  AND3_X1 u2_u9_u2_U45 (.A2( u2_u9_u2_n100 ) , .A1( u2_u9_u2_n104 ) , .A3( u2_u9_u2_n156 ) , .ZN( u2_u9_u2_n95 ) );
  OAI21_X1 u2_u9_u2_U46 (.A( u2_u9_u2_n141 ) , .B2( u2_u9_u2_n142 ) , .ZN( u2_u9_u2_n146 ) , .B1( u2_u9_u2_n153 ) );
  OAI21_X1 u2_u9_u2_U47 (.A( u2_u9_u2_n140 ) , .ZN( u2_u9_u2_n141 ) , .B1( u2_u9_u2_n176 ) , .B2( u2_u9_u2_n177 ) );
  NOR3_X1 u2_u9_u2_U48 (.ZN( u2_u9_u2_n142 ) , .A3( u2_u9_u2_n175 ) , .A2( u2_u9_u2_n178 ) , .A1( u2_u9_u2_n181 ) );
  OAI21_X1 u2_u9_u2_U49 (.A( u2_u9_u2_n101 ) , .B2( u2_u9_u2_n121 ) , .B1( u2_u9_u2_n153 ) , .ZN( u2_u9_u2_n164 ) );
  NOR4_X1 u2_u9_u2_U5 (.A4( u2_u9_u2_n124 ) , .A3( u2_u9_u2_n125 ) , .A2( u2_u9_u2_n126 ) , .A1( u2_u9_u2_n127 ) , .ZN( u2_u9_u2_n128 ) );
  NAND2_X1 u2_u9_u2_U50 (.A2( u2_u9_u2_n100 ) , .A1( u2_u9_u2_n107 ) , .ZN( u2_u9_u2_n155 ) );
  NAND2_X1 u2_u9_u2_U51 (.A2( u2_u9_u2_n105 ) , .A1( u2_u9_u2_n108 ) , .ZN( u2_u9_u2_n143 ) );
  NAND2_X1 u2_u9_u2_U52 (.A1( u2_u9_u2_n104 ) , .A2( u2_u9_u2_n106 ) , .ZN( u2_u9_u2_n152 ) );
  NAND2_X1 u2_u9_u2_U53 (.A1( u2_u9_u2_n100 ) , .A2( u2_u9_u2_n105 ) , .ZN( u2_u9_u2_n132 ) );
  INV_X1 u2_u9_u2_U54 (.A( u2_u9_u2_n140 ) , .ZN( u2_u9_u2_n168 ) );
  INV_X1 u2_u9_u2_U55 (.A( u2_u9_u2_n138 ) , .ZN( u2_u9_u2_n167 ) );
  NAND2_X1 u2_u9_u2_U56 (.A1( u2_u9_u2_n102 ) , .A2( u2_u9_u2_n106 ) , .ZN( u2_u9_u2_n113 ) );
  NAND2_X1 u2_u9_u2_U57 (.A1( u2_u9_u2_n106 ) , .A2( u2_u9_u2_n107 ) , .ZN( u2_u9_u2_n131 ) );
  NAND2_X1 u2_u9_u2_U58 (.A1( u2_u9_u2_n103 ) , .A2( u2_u9_u2_n107 ) , .ZN( u2_u9_u2_n139 ) );
  NAND2_X1 u2_u9_u2_U59 (.A1( u2_u9_u2_n103 ) , .A2( u2_u9_u2_n105 ) , .ZN( u2_u9_u2_n133 ) );
  AOI21_X1 u2_u9_u2_U6 (.B2( u2_u9_u2_n119 ) , .ZN( u2_u9_u2_n127 ) , .A( u2_u9_u2_n137 ) , .B1( u2_u9_u2_n155 ) );
  NAND2_X1 u2_u9_u2_U60 (.A1( u2_u9_u2_n102 ) , .A2( u2_u9_u2_n103 ) , .ZN( u2_u9_u2_n154 ) );
  NAND2_X1 u2_u9_u2_U61 (.A2( u2_u9_u2_n103 ) , .A1( u2_u9_u2_n104 ) , .ZN( u2_u9_u2_n119 ) );
  NAND2_X1 u2_u9_u2_U62 (.A2( u2_u9_u2_n107 ) , .A1( u2_u9_u2_n108 ) , .ZN( u2_u9_u2_n123 ) );
  NAND2_X1 u2_u9_u2_U63 (.A1( u2_u9_u2_n104 ) , .A2( u2_u9_u2_n108 ) , .ZN( u2_u9_u2_n122 ) );
  INV_X1 u2_u9_u2_U64 (.A( u2_u9_u2_n114 ) , .ZN( u2_u9_u2_n172 ) );
  NAND2_X1 u2_u9_u2_U65 (.A2( u2_u9_u2_n100 ) , .A1( u2_u9_u2_n102 ) , .ZN( u2_u9_u2_n116 ) );
  NAND2_X1 u2_u9_u2_U66 (.A1( u2_u9_u2_n102 ) , .A2( u2_u9_u2_n108 ) , .ZN( u2_u9_u2_n120 ) );
  NAND2_X1 u2_u9_u2_U67 (.A2( u2_u9_u2_n105 ) , .A1( u2_u9_u2_n106 ) , .ZN( u2_u9_u2_n117 ) );
  INV_X1 u2_u9_u2_U68 (.ZN( u2_u9_u2_n187 ) , .A( u2_u9_u2_n99 ) );
  OAI21_X1 u2_u9_u2_U69 (.B1( u2_u9_u2_n137 ) , .B2( u2_u9_u2_n143 ) , .A( u2_u9_u2_n98 ) , .ZN( u2_u9_u2_n99 ) );
  AOI21_X1 u2_u9_u2_U7 (.ZN( u2_u9_u2_n124 ) , .B1( u2_u9_u2_n131 ) , .B2( u2_u9_u2_n143 ) , .A( u2_u9_u2_n172 ) );
  NOR2_X1 u2_u9_u2_U70 (.A2( u2_u9_X_16 ) , .ZN( u2_u9_u2_n140 ) , .A1( u2_u9_u2_n166 ) );
  NOR2_X1 u2_u9_u2_U71 (.A2( u2_u9_X_13 ) , .A1( u2_u9_X_14 ) , .ZN( u2_u9_u2_n100 ) );
  NOR2_X1 u2_u9_u2_U72 (.A2( u2_u9_X_16 ) , .A1( u2_u9_X_17 ) , .ZN( u2_u9_u2_n138 ) );
  NOR2_X1 u2_u9_u2_U73 (.A2( u2_u9_X_15 ) , .A1( u2_u9_X_18 ) , .ZN( u2_u9_u2_n104 ) );
  NOR2_X1 u2_u9_u2_U74 (.A2( u2_u9_X_14 ) , .ZN( u2_u9_u2_n103 ) , .A1( u2_u9_u2_n174 ) );
  NOR2_X1 u2_u9_u2_U75 (.A2( u2_u9_X_15 ) , .ZN( u2_u9_u2_n102 ) , .A1( u2_u9_u2_n165 ) );
  NOR2_X1 u2_u9_u2_U76 (.A2( u2_u9_X_17 ) , .ZN( u2_u9_u2_n114 ) , .A1( u2_u9_u2_n169 ) );
  AND2_X1 u2_u9_u2_U77 (.A1( u2_u9_X_15 ) , .ZN( u2_u9_u2_n105 ) , .A2( u2_u9_u2_n165 ) );
  AND2_X1 u2_u9_u2_U78 (.A2( u2_u9_X_15 ) , .A1( u2_u9_X_18 ) , .ZN( u2_u9_u2_n107 ) );
  AND2_X1 u2_u9_u2_U79 (.A1( u2_u9_X_14 ) , .ZN( u2_u9_u2_n106 ) , .A2( u2_u9_u2_n174 ) );
  AOI21_X1 u2_u9_u2_U8 (.B2( u2_u9_u2_n120 ) , .B1( u2_u9_u2_n121 ) , .ZN( u2_u9_u2_n126 ) , .A( u2_u9_u2_n167 ) );
  AND2_X1 u2_u9_u2_U80 (.A1( u2_u9_X_13 ) , .A2( u2_u9_X_14 ) , .ZN( u2_u9_u2_n108 ) );
  INV_X1 u2_u9_u2_U81 (.A( u2_u9_X_16 ) , .ZN( u2_u9_u2_n169 ) );
  INV_X1 u2_u9_u2_U82 (.A( u2_u9_X_17 ) , .ZN( u2_u9_u2_n166 ) );
  INV_X1 u2_u9_u2_U83 (.A( u2_u9_X_13 ) , .ZN( u2_u9_u2_n174 ) );
  INV_X1 u2_u9_u2_U84 (.A( u2_u9_X_18 ) , .ZN( u2_u9_u2_n165 ) );
  NAND4_X1 u2_u9_u2_U85 (.ZN( u2_out9_30 ) , .A4( u2_u9_u2_n147 ) , .A3( u2_u9_u2_n148 ) , .A2( u2_u9_u2_n149 ) , .A1( u2_u9_u2_n187 ) );
  AOI21_X1 u2_u9_u2_U86 (.B2( u2_u9_u2_n138 ) , .ZN( u2_u9_u2_n148 ) , .A( u2_u9_u2_n162 ) , .B1( u2_u9_u2_n182 ) );
  NOR3_X1 u2_u9_u2_U87 (.A3( u2_u9_u2_n144 ) , .A2( u2_u9_u2_n145 ) , .A1( u2_u9_u2_n146 ) , .ZN( u2_u9_u2_n147 ) );
  NAND4_X1 u2_u9_u2_U88 (.ZN( u2_out9_24 ) , .A4( u2_u9_u2_n111 ) , .A3( u2_u9_u2_n112 ) , .A1( u2_u9_u2_n130 ) , .A2( u2_u9_u2_n187 ) );
  AOI221_X1 u2_u9_u2_U89 (.A( u2_u9_u2_n109 ) , .B1( u2_u9_u2_n110 ) , .ZN( u2_u9_u2_n111 ) , .C1( u2_u9_u2_n134 ) , .C2( u2_u9_u2_n170 ) , .B2( u2_u9_u2_n173 ) );
  OAI22_X1 u2_u9_u2_U9 (.ZN( u2_u9_u2_n109 ) , .A2( u2_u9_u2_n113 ) , .B2( u2_u9_u2_n133 ) , .B1( u2_u9_u2_n167 ) , .A1( u2_u9_u2_n168 ) );
  AOI21_X1 u2_u9_u2_U90 (.ZN( u2_u9_u2_n112 ) , .B2( u2_u9_u2_n156 ) , .A( u2_u9_u2_n164 ) , .B1( u2_u9_u2_n181 ) );
  NAND4_X1 u2_u9_u2_U91 (.ZN( u2_out9_16 ) , .A4( u2_u9_u2_n128 ) , .A3( u2_u9_u2_n129 ) , .A1( u2_u9_u2_n130 ) , .A2( u2_u9_u2_n186 ) );
  AOI22_X1 u2_u9_u2_U92 (.A2( u2_u9_u2_n118 ) , .ZN( u2_u9_u2_n129 ) , .A1( u2_u9_u2_n140 ) , .B1( u2_u9_u2_n157 ) , .B2( u2_u9_u2_n170 ) );
  INV_X1 u2_u9_u2_U93 (.A( u2_u9_u2_n163 ) , .ZN( u2_u9_u2_n186 ) );
  OR4_X1 u2_u9_u2_U94 (.ZN( u2_out9_6 ) , .A4( u2_u9_u2_n161 ) , .A3( u2_u9_u2_n162 ) , .A2( u2_u9_u2_n163 ) , .A1( u2_u9_u2_n164 ) );
  OR3_X1 u2_u9_u2_U95 (.A2( u2_u9_u2_n159 ) , .A1( u2_u9_u2_n160 ) , .ZN( u2_u9_u2_n161 ) , .A3( u2_u9_u2_n183 ) );
  AOI21_X1 u2_u9_u2_U96 (.B2( u2_u9_u2_n154 ) , .B1( u2_u9_u2_n155 ) , .ZN( u2_u9_u2_n159 ) , .A( u2_u9_u2_n167 ) );
  NAND3_X1 u2_u9_u2_U97 (.A2( u2_u9_u2_n117 ) , .A1( u2_u9_u2_n122 ) , .A3( u2_u9_u2_n123 ) , .ZN( u2_u9_u2_n134 ) );
  NAND3_X1 u2_u9_u2_U98 (.ZN( u2_u9_u2_n110 ) , .A2( u2_u9_u2_n131 ) , .A3( u2_u9_u2_n139 ) , .A1( u2_u9_u2_n154 ) );
  NAND3_X1 u2_u9_u2_U99 (.A2( u2_u9_u2_n100 ) , .ZN( u2_u9_u2_n101 ) , .A1( u2_u9_u2_n104 ) , .A3( u2_u9_u2_n114 ) );
  AND3_X1 u2_u9_u7_U10 (.A3( u2_u9_u7_n110 ) , .A2( u2_u9_u7_n127 ) , .A1( u2_u9_u7_n132 ) , .ZN( u2_u9_u7_n92 ) );
  OAI21_X1 u2_u9_u7_U11 (.A( u2_u9_u7_n161 ) , .B1( u2_u9_u7_n168 ) , .B2( u2_u9_u7_n173 ) , .ZN( u2_u9_u7_n91 ) );
  AOI211_X1 u2_u9_u7_U12 (.A( u2_u9_u7_n117 ) , .ZN( u2_u9_u7_n118 ) , .C2( u2_u9_u7_n126 ) , .C1( u2_u9_u7_n177 ) , .B( u2_u9_u7_n180 ) );
  OAI22_X1 u2_u9_u7_U13 (.B1( u2_u9_u7_n115 ) , .ZN( u2_u9_u7_n117 ) , .A2( u2_u9_u7_n133 ) , .A1( u2_u9_u7_n137 ) , .B2( u2_u9_u7_n162 ) );
  INV_X1 u2_u9_u7_U14 (.A( u2_u9_u7_n116 ) , .ZN( u2_u9_u7_n180 ) );
  NOR3_X1 u2_u9_u7_U15 (.ZN( u2_u9_u7_n115 ) , .A3( u2_u9_u7_n145 ) , .A2( u2_u9_u7_n168 ) , .A1( u2_u9_u7_n169 ) );
  OAI211_X1 u2_u9_u7_U16 (.B( u2_u9_u7_n122 ) , .A( u2_u9_u7_n123 ) , .C2( u2_u9_u7_n124 ) , .ZN( u2_u9_u7_n154 ) , .C1( u2_u9_u7_n162 ) );
  AOI222_X1 u2_u9_u7_U17 (.ZN( u2_u9_u7_n122 ) , .C2( u2_u9_u7_n126 ) , .C1( u2_u9_u7_n145 ) , .B1( u2_u9_u7_n161 ) , .A2( u2_u9_u7_n165 ) , .B2( u2_u9_u7_n170 ) , .A1( u2_u9_u7_n176 ) );
  INV_X1 u2_u9_u7_U18 (.A( u2_u9_u7_n133 ) , .ZN( u2_u9_u7_n176 ) );
  NOR3_X1 u2_u9_u7_U19 (.A2( u2_u9_u7_n134 ) , .A1( u2_u9_u7_n135 ) , .ZN( u2_u9_u7_n136 ) , .A3( u2_u9_u7_n171 ) );
  NOR2_X1 u2_u9_u7_U20 (.A1( u2_u9_u7_n130 ) , .A2( u2_u9_u7_n134 ) , .ZN( u2_u9_u7_n153 ) );
  INV_X1 u2_u9_u7_U21 (.A( u2_u9_u7_n101 ) , .ZN( u2_u9_u7_n165 ) );
  NOR2_X1 u2_u9_u7_U22 (.ZN( u2_u9_u7_n111 ) , .A2( u2_u9_u7_n134 ) , .A1( u2_u9_u7_n169 ) );
  AOI21_X1 u2_u9_u7_U23 (.ZN( u2_u9_u7_n104 ) , .B2( u2_u9_u7_n112 ) , .B1( u2_u9_u7_n127 ) , .A( u2_u9_u7_n164 ) );
  AOI21_X1 u2_u9_u7_U24 (.ZN( u2_u9_u7_n106 ) , .B1( u2_u9_u7_n133 ) , .B2( u2_u9_u7_n146 ) , .A( u2_u9_u7_n162 ) );
  AOI21_X1 u2_u9_u7_U25 (.A( u2_u9_u7_n101 ) , .ZN( u2_u9_u7_n107 ) , .B2( u2_u9_u7_n128 ) , .B1( u2_u9_u7_n175 ) );
  INV_X1 u2_u9_u7_U26 (.A( u2_u9_u7_n138 ) , .ZN( u2_u9_u7_n171 ) );
  INV_X1 u2_u9_u7_U27 (.A( u2_u9_u7_n131 ) , .ZN( u2_u9_u7_n177 ) );
  INV_X1 u2_u9_u7_U28 (.A( u2_u9_u7_n110 ) , .ZN( u2_u9_u7_n174 ) );
  NAND2_X1 u2_u9_u7_U29 (.A1( u2_u9_u7_n129 ) , .A2( u2_u9_u7_n132 ) , .ZN( u2_u9_u7_n149 ) );
  OAI21_X1 u2_u9_u7_U3 (.ZN( u2_u9_u7_n159 ) , .A( u2_u9_u7_n165 ) , .B2( u2_u9_u7_n171 ) , .B1( u2_u9_u7_n174 ) );
  NAND2_X1 u2_u9_u7_U30 (.A1( u2_u9_u7_n113 ) , .A2( u2_u9_u7_n124 ) , .ZN( u2_u9_u7_n130 ) );
  INV_X1 u2_u9_u7_U31 (.A( u2_u9_u7_n112 ) , .ZN( u2_u9_u7_n173 ) );
  INV_X1 u2_u9_u7_U32 (.A( u2_u9_u7_n128 ) , .ZN( u2_u9_u7_n168 ) );
  INV_X1 u2_u9_u7_U33 (.A( u2_u9_u7_n148 ) , .ZN( u2_u9_u7_n169 ) );
  INV_X1 u2_u9_u7_U34 (.A( u2_u9_u7_n127 ) , .ZN( u2_u9_u7_n179 ) );
  NOR2_X1 u2_u9_u7_U35 (.ZN( u2_u9_u7_n101 ) , .A2( u2_u9_u7_n150 ) , .A1( u2_u9_u7_n156 ) );
  AOI211_X1 u2_u9_u7_U36 (.B( u2_u9_u7_n154 ) , .A( u2_u9_u7_n155 ) , .C1( u2_u9_u7_n156 ) , .ZN( u2_u9_u7_n157 ) , .C2( u2_u9_u7_n172 ) );
  INV_X1 u2_u9_u7_U37 (.A( u2_u9_u7_n153 ) , .ZN( u2_u9_u7_n172 ) );
  AOI211_X1 u2_u9_u7_U38 (.B( u2_u9_u7_n139 ) , .A( u2_u9_u7_n140 ) , .C2( u2_u9_u7_n141 ) , .ZN( u2_u9_u7_n142 ) , .C1( u2_u9_u7_n156 ) );
  NAND4_X1 u2_u9_u7_U39 (.A3( u2_u9_u7_n127 ) , .A2( u2_u9_u7_n128 ) , .A1( u2_u9_u7_n129 ) , .ZN( u2_u9_u7_n141 ) , .A4( u2_u9_u7_n147 ) );
  INV_X1 u2_u9_u7_U4 (.A( u2_u9_u7_n111 ) , .ZN( u2_u9_u7_n170 ) );
  AOI21_X1 u2_u9_u7_U40 (.A( u2_u9_u7_n137 ) , .B1( u2_u9_u7_n138 ) , .ZN( u2_u9_u7_n139 ) , .B2( u2_u9_u7_n146 ) );
  OAI22_X1 u2_u9_u7_U41 (.B1( u2_u9_u7_n136 ) , .ZN( u2_u9_u7_n140 ) , .A1( u2_u9_u7_n153 ) , .B2( u2_u9_u7_n162 ) , .A2( u2_u9_u7_n164 ) );
  AOI21_X1 u2_u9_u7_U42 (.ZN( u2_u9_u7_n123 ) , .B1( u2_u9_u7_n165 ) , .B2( u2_u9_u7_n177 ) , .A( u2_u9_u7_n97 ) );
  AOI21_X1 u2_u9_u7_U43 (.B2( u2_u9_u7_n113 ) , .B1( u2_u9_u7_n124 ) , .A( u2_u9_u7_n125 ) , .ZN( u2_u9_u7_n97 ) );
  INV_X1 u2_u9_u7_U44 (.A( u2_u9_u7_n125 ) , .ZN( u2_u9_u7_n161 ) );
  INV_X1 u2_u9_u7_U45 (.A( u2_u9_u7_n152 ) , .ZN( u2_u9_u7_n162 ) );
  AOI22_X1 u2_u9_u7_U46 (.A2( u2_u9_u7_n114 ) , .ZN( u2_u9_u7_n119 ) , .B1( u2_u9_u7_n130 ) , .A1( u2_u9_u7_n156 ) , .B2( u2_u9_u7_n165 ) );
  NAND2_X1 u2_u9_u7_U47 (.A2( u2_u9_u7_n112 ) , .ZN( u2_u9_u7_n114 ) , .A1( u2_u9_u7_n175 ) );
  AND2_X1 u2_u9_u7_U48 (.ZN( u2_u9_u7_n145 ) , .A2( u2_u9_u7_n98 ) , .A1( u2_u9_u7_n99 ) );
  NOR2_X1 u2_u9_u7_U49 (.ZN( u2_u9_u7_n137 ) , .A1( u2_u9_u7_n150 ) , .A2( u2_u9_u7_n161 ) );
  INV_X1 u2_u9_u7_U5 (.A( u2_u9_u7_n149 ) , .ZN( u2_u9_u7_n175 ) );
  AOI21_X1 u2_u9_u7_U50 (.ZN( u2_u9_u7_n105 ) , .B2( u2_u9_u7_n110 ) , .A( u2_u9_u7_n125 ) , .B1( u2_u9_u7_n147 ) );
  NAND2_X1 u2_u9_u7_U51 (.ZN( u2_u9_u7_n146 ) , .A1( u2_u9_u7_n95 ) , .A2( u2_u9_u7_n98 ) );
  NAND2_X1 u2_u9_u7_U52 (.A2( u2_u9_u7_n103 ) , .ZN( u2_u9_u7_n147 ) , .A1( u2_u9_u7_n93 ) );
  NAND2_X1 u2_u9_u7_U53 (.A1( u2_u9_u7_n103 ) , .ZN( u2_u9_u7_n127 ) , .A2( u2_u9_u7_n99 ) );
  OR2_X1 u2_u9_u7_U54 (.ZN( u2_u9_u7_n126 ) , .A2( u2_u9_u7_n152 ) , .A1( u2_u9_u7_n156 ) );
  NAND2_X1 u2_u9_u7_U55 (.A2( u2_u9_u7_n102 ) , .A1( u2_u9_u7_n103 ) , .ZN( u2_u9_u7_n133 ) );
  NAND2_X1 u2_u9_u7_U56 (.ZN( u2_u9_u7_n112 ) , .A2( u2_u9_u7_n96 ) , .A1( u2_u9_u7_n99 ) );
  NAND2_X1 u2_u9_u7_U57 (.A2( u2_u9_u7_n102 ) , .ZN( u2_u9_u7_n128 ) , .A1( u2_u9_u7_n98 ) );
  NAND2_X1 u2_u9_u7_U58 (.A1( u2_u9_u7_n100 ) , .ZN( u2_u9_u7_n113 ) , .A2( u2_u9_u7_n93 ) );
  NAND2_X1 u2_u9_u7_U59 (.A2( u2_u9_u7_n102 ) , .ZN( u2_u9_u7_n124 ) , .A1( u2_u9_u7_n96 ) );
  INV_X1 u2_u9_u7_U6 (.A( u2_u9_u7_n154 ) , .ZN( u2_u9_u7_n178 ) );
  NAND2_X1 u2_u9_u7_U60 (.ZN( u2_u9_u7_n110 ) , .A1( u2_u9_u7_n95 ) , .A2( u2_u9_u7_n96 ) );
  INV_X1 u2_u9_u7_U61 (.A( u2_u9_u7_n150 ) , .ZN( u2_u9_u7_n164 ) );
  AND2_X1 u2_u9_u7_U62 (.ZN( u2_u9_u7_n134 ) , .A1( u2_u9_u7_n93 ) , .A2( u2_u9_u7_n98 ) );
  NAND2_X1 u2_u9_u7_U63 (.A1( u2_u9_u7_n100 ) , .A2( u2_u9_u7_n102 ) , .ZN( u2_u9_u7_n129 ) );
  NAND2_X1 u2_u9_u7_U64 (.A2( u2_u9_u7_n103 ) , .ZN( u2_u9_u7_n131 ) , .A1( u2_u9_u7_n95 ) );
  NAND2_X1 u2_u9_u7_U65 (.A1( u2_u9_u7_n100 ) , .ZN( u2_u9_u7_n138 ) , .A2( u2_u9_u7_n99 ) );
  NAND2_X1 u2_u9_u7_U66 (.ZN( u2_u9_u7_n132 ) , .A1( u2_u9_u7_n93 ) , .A2( u2_u9_u7_n96 ) );
  NAND2_X1 u2_u9_u7_U67 (.A1( u2_u9_u7_n100 ) , .ZN( u2_u9_u7_n148 ) , .A2( u2_u9_u7_n95 ) );
  NOR2_X1 u2_u9_u7_U68 (.A2( u2_u9_X_47 ) , .ZN( u2_u9_u7_n150 ) , .A1( u2_u9_u7_n163 ) );
  NOR2_X1 u2_u9_u7_U69 (.A2( u2_u9_X_43 ) , .A1( u2_u9_X_44 ) , .ZN( u2_u9_u7_n103 ) );
  AOI211_X1 u2_u9_u7_U7 (.ZN( u2_u9_u7_n116 ) , .A( u2_u9_u7_n155 ) , .C1( u2_u9_u7_n161 ) , .C2( u2_u9_u7_n171 ) , .B( u2_u9_u7_n94 ) );
  NOR2_X1 u2_u9_u7_U70 (.A2( u2_u9_X_48 ) , .A1( u2_u9_u7_n166 ) , .ZN( u2_u9_u7_n95 ) );
  NOR2_X1 u2_u9_u7_U71 (.A2( u2_u9_X_45 ) , .A1( u2_u9_X_48 ) , .ZN( u2_u9_u7_n99 ) );
  NOR2_X1 u2_u9_u7_U72 (.A2( u2_u9_X_44 ) , .A1( u2_u9_u7_n167 ) , .ZN( u2_u9_u7_n98 ) );
  NOR2_X1 u2_u9_u7_U73 (.A2( u2_u9_X_46 ) , .A1( u2_u9_X_47 ) , .ZN( u2_u9_u7_n152 ) );
  AND2_X1 u2_u9_u7_U74 (.A1( u2_u9_X_47 ) , .ZN( u2_u9_u7_n156 ) , .A2( u2_u9_u7_n163 ) );
  NAND2_X1 u2_u9_u7_U75 (.A2( u2_u9_X_46 ) , .A1( u2_u9_X_47 ) , .ZN( u2_u9_u7_n125 ) );
  AND2_X1 u2_u9_u7_U76 (.A2( u2_u9_X_45 ) , .A1( u2_u9_X_48 ) , .ZN( u2_u9_u7_n102 ) );
  AND2_X1 u2_u9_u7_U77 (.A2( u2_u9_X_43 ) , .A1( u2_u9_X_44 ) , .ZN( u2_u9_u7_n96 ) );
  AND2_X1 u2_u9_u7_U78 (.A1( u2_u9_X_44 ) , .ZN( u2_u9_u7_n100 ) , .A2( u2_u9_u7_n167 ) );
  AND2_X1 u2_u9_u7_U79 (.A1( u2_u9_X_48 ) , .A2( u2_u9_u7_n166 ) , .ZN( u2_u9_u7_n93 ) );
  OAI222_X1 u2_u9_u7_U8 (.C2( u2_u9_u7_n101 ) , .B2( u2_u9_u7_n111 ) , .A1( u2_u9_u7_n113 ) , .C1( u2_u9_u7_n146 ) , .A2( u2_u9_u7_n162 ) , .B1( u2_u9_u7_n164 ) , .ZN( u2_u9_u7_n94 ) );
  INV_X1 u2_u9_u7_U80 (.A( u2_u9_X_46 ) , .ZN( u2_u9_u7_n163 ) );
  INV_X1 u2_u9_u7_U81 (.A( u2_u9_X_43 ) , .ZN( u2_u9_u7_n167 ) );
  INV_X1 u2_u9_u7_U82 (.A( u2_u9_X_45 ) , .ZN( u2_u9_u7_n166 ) );
  NAND4_X1 u2_u9_u7_U83 (.ZN( u2_out9_27 ) , .A4( u2_u9_u7_n118 ) , .A3( u2_u9_u7_n119 ) , .A2( u2_u9_u7_n120 ) , .A1( u2_u9_u7_n121 ) );
  OAI21_X1 u2_u9_u7_U84 (.ZN( u2_u9_u7_n121 ) , .B2( u2_u9_u7_n145 ) , .A( u2_u9_u7_n150 ) , .B1( u2_u9_u7_n174 ) );
  OAI21_X1 u2_u9_u7_U85 (.ZN( u2_u9_u7_n120 ) , .A( u2_u9_u7_n161 ) , .B2( u2_u9_u7_n170 ) , .B1( u2_u9_u7_n179 ) );
  NAND4_X1 u2_u9_u7_U86 (.ZN( u2_out9_21 ) , .A4( u2_u9_u7_n157 ) , .A3( u2_u9_u7_n158 ) , .A2( u2_u9_u7_n159 ) , .A1( u2_u9_u7_n160 ) );
  OAI21_X1 u2_u9_u7_U87 (.B1( u2_u9_u7_n145 ) , .ZN( u2_u9_u7_n160 ) , .A( u2_u9_u7_n161 ) , .B2( u2_u9_u7_n177 ) );
  AOI22_X1 u2_u9_u7_U88 (.B2( u2_u9_u7_n149 ) , .B1( u2_u9_u7_n150 ) , .A2( u2_u9_u7_n151 ) , .A1( u2_u9_u7_n152 ) , .ZN( u2_u9_u7_n158 ) );
  NAND4_X1 u2_u9_u7_U89 (.ZN( u2_out9_15 ) , .A4( u2_u9_u7_n142 ) , .A3( u2_u9_u7_n143 ) , .A2( u2_u9_u7_n144 ) , .A1( u2_u9_u7_n178 ) );
  OAI221_X1 u2_u9_u7_U9 (.C1( u2_u9_u7_n101 ) , .C2( u2_u9_u7_n147 ) , .ZN( u2_u9_u7_n155 ) , .B2( u2_u9_u7_n162 ) , .A( u2_u9_u7_n91 ) , .B1( u2_u9_u7_n92 ) );
  OR2_X1 u2_u9_u7_U90 (.A2( u2_u9_u7_n125 ) , .A1( u2_u9_u7_n129 ) , .ZN( u2_u9_u7_n144 ) );
  AOI22_X1 u2_u9_u7_U91 (.A2( u2_u9_u7_n126 ) , .ZN( u2_u9_u7_n143 ) , .B2( u2_u9_u7_n165 ) , .B1( u2_u9_u7_n173 ) , .A1( u2_u9_u7_n174 ) );
  NAND4_X1 u2_u9_u7_U92 (.ZN( u2_out9_5 ) , .A4( u2_u9_u7_n108 ) , .A3( u2_u9_u7_n109 ) , .A1( u2_u9_u7_n116 ) , .A2( u2_u9_u7_n123 ) );
  AOI22_X1 u2_u9_u7_U93 (.ZN( u2_u9_u7_n109 ) , .A2( u2_u9_u7_n126 ) , .B2( u2_u9_u7_n145 ) , .B1( u2_u9_u7_n156 ) , .A1( u2_u9_u7_n171 ) );
  NOR4_X1 u2_u9_u7_U94 (.A4( u2_u9_u7_n104 ) , .A3( u2_u9_u7_n105 ) , .A2( u2_u9_u7_n106 ) , .A1( u2_u9_u7_n107 ) , .ZN( u2_u9_u7_n108 ) );
  NAND3_X1 u2_u9_u7_U95 (.A3( u2_u9_u7_n146 ) , .A2( u2_u9_u7_n147 ) , .A1( u2_u9_u7_n148 ) , .ZN( u2_u9_u7_n151 ) );
  NAND3_X1 u2_u9_u7_U96 (.A3( u2_u9_u7_n131 ) , .A2( u2_u9_u7_n132 ) , .A1( u2_u9_u7_n133 ) , .ZN( u2_u9_u7_n135 ) );
  NAND2_X1 u2_uk_U1000 (.A1( u2_key_r_46 ) , .A2( u2_uk_n100 ) , .ZN( u2_uk_n969 ) );
  OAI21_X1 u2_uk_U1001 (.ZN( u2_K1_17 ) , .B1( u2_uk_n100 ) , .B2( u2_uk_n1153 ) , .A( u2_uk_n971 ) );
  NAND2_X1 u2_uk_U1002 (.A1( u2_key_r_10 ) , .A2( u2_uk_n27 ) , .ZN( u2_uk_n971 ) );
  OAI21_X1 u2_uk_U1003 (.ZN( u2_K12_7 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1720 ) , .A( u2_uk_n520 ) );
  NAND2_X1 u2_uk_U1008 (.A1( u2_key_r_50 ) , .A2( u2_uk_n31 ) , .ZN( u2_uk_n983 ) );
  OAI21_X1 u2_uk_U1015 (.ZN( u2_K8_46 ) , .A( u2_uk_n1115 ) , .B2( u2_uk_n1532 ) , .B1( u2_uk_n182 ) );
  NAND2_X1 u2_uk_U1016 (.A1( u2_uk_K_r6_37 ) , .ZN( u2_uk_n1115 ) , .A2( u2_uk_n155 ) );
  OAI21_X1 u2_uk_U1017 (.ZN( u2_K10_13 ) , .B1( u2_uk_n109 ) , .B2( u2_uk_n1605 ) , .A( u2_uk_n242 ) );
  NAND2_X1 u2_uk_U1018 (.A1( u2_uk_K_r8_48 ) , .A2( u2_uk_n10 ) , .ZN( u2_uk_n242 ) );
  OAI21_X1 u2_uk_U1025 (.ZN( u2_K4_28 ) , .A( u2_uk_n1029 ) , .B2( u2_uk_n1351 ) , .B1( u2_uk_n17 ) );
  NAND2_X1 u2_uk_U1026 (.A1( u2_uk_K_r2_21 ) , .ZN( u2_uk_n1029 ) , .A2( u2_uk_n99 ) );
  NAND2_X1 u2_uk_U1028 (.A1( u2_uk_K_r5_16 ) , .ZN( u2_uk_n1087 ) , .A2( u2_uk_n17 ) );
  OAI21_X1 u2_uk_U1033 (.ZN( u2_K15_32 ) , .B1( u2_uk_n109 ) , .B2( u2_uk_n1825 ) , .A( u2_uk_n941 ) );
  NAND2_X1 u2_uk_U1042 (.A1( u2_uk_K_r9_0 ) , .A2( u2_uk_n10 ) , .ZN( u2_uk_n366 ) );
  INV_X1 u2_uk_U1045 (.A( u2_key_r_6 ) , .ZN( u2_uk_n1146 ) );
  INV_X1 u2_uk_U1048 (.A( u2_key_r_26 ) , .ZN( u2_uk_n1161 ) );
  INV_X1 u2_uk_U1050 (.A( u2_key_r_47 ) , .ZN( u2_uk_n1179 ) );
  INV_X1 u2_uk_U1051 (.A( u2_key_r_34 ) , .ZN( u2_uk_n1168 ) );
  INV_X1 u2_uk_U1052 (.A( u2_key_r_27 ) , .ZN( u2_uk_n1162 ) );
  INV_X1 u2_uk_U1053 (.A( u2_key_r_24 ) , .ZN( u2_uk_n1159 ) );
  INV_X1 u2_uk_U1054 (.A( u2_key_r_20 ) , .ZN( u2_uk_n1155 ) );
  INV_X1 u2_uk_U1062 (.A( u2_key_r_19 ) , .ZN( u2_uk_n1154 ) );
  INV_X1 u2_uk_U1063 (.A( u2_key_r_4 ) , .ZN( u2_uk_n1145 ) );
  INV_X1 u2_uk_U1064 (.A( u2_key_r_17 ) , .ZN( u2_uk_n1153 ) );
  INV_X1 u2_uk_U1065 (.A( u2_key_r_53 ) , .ZN( u2_uk_n1184 ) );
  OAI21_X1 u2_uk_U1072 (.ZN( u2_K3_40 ) , .A( u2_uk_n1014 ) , .B2( u2_uk_n1300 ) , .B1( u2_uk_n230 ) );
  NAND2_X1 u2_uk_U1073 (.A1( u2_uk_K_r1_21 ) , .ZN( u2_uk_n1014 ) , .A2( u2_uk_n148 ) );
  OAI21_X1 u2_uk_U1074 (.ZN( u2_K16_39 ) , .B2( u2_uk_n1201 ) , .B1( u2_uk_n202 ) , .A( u2_uk_n960 ) );
  NAND2_X1 u2_uk_U1075 (.A1( u2_uk_K_r14_15 ) , .A2( u2_uk_n147 ) , .ZN( u2_uk_n960 ) );
  OAI21_X1 u2_uk_U1076 (.ZN( u2_K8_39 ) , .A( u2_uk_n1109 ) , .B2( u2_uk_n1526 ) , .B1( u2_uk_n202 ) );
  NAND2_X1 u2_uk_U1077 (.A1( u2_uk_K_r6_31 ) , .ZN( u2_uk_n1109 ) , .A2( u2_uk_n155 ) );
  INV_X1 u2_uk_U1080 (.A( u2_key_r_40 ) , .ZN( u2_uk_n1174 ) );
  INV_X1 u2_uk_U1084 (.ZN( u2_K1_11 ) , .A( u2_uk_n967 ) );
  INV_X1 u2_uk_U1086 (.ZN( u2_K1_18 ) , .A( u2_uk_n972 ) );
  OAI22_X1 u2_uk_U109 (.ZN( u2_K3_41 ) , .A2( u2_uk_n1283 ) , .B2( u2_uk_n1288 ) , .B1( u2_uk_n141 ) , .A1( u2_uk_n83 ) );
  INV_X1 u2_uk_U1090 (.ZN( u2_K7_6 ) , .A( u2_uk_n1095 ) );
  AOI22_X1 u2_uk_U1091 (.B2( u2_uk_K_r5_39 ) , .A2( u2_uk_K_r5_4 ) , .ZN( u2_uk_n1095 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n182 ) );
  INV_X1 u2_uk_U1100 (.ZN( u2_K1_20 ) , .A( u2_uk_n973 ) );
  AOI22_X1 u2_uk_U1101 (.B2( u2_key_r_48 ) , .A2( u2_key_r_55 ) , .A1( u2_uk_n202 ) , .B1( u2_uk_n63 ) , .ZN( u2_uk_n973 ) );
  INV_X1 u2_uk_U1114 (.ZN( u2_K5_20 ) , .A( u2_uk_n1043 ) );
  INV_X1 u2_uk_U1116 (.ZN( u2_K7_13 ) , .A( u2_uk_n1076 ) );
  AOI22_X1 u2_uk_U1117 (.B2( u2_uk_K_r5_26 ) , .A2( u2_uk_K_r5_48 ) , .ZN( u2_uk_n1076 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n145 ) );
  INV_X1 u2_uk_U1122 (.ZN( u2_K4_20 ) , .A( u2_uk_n1024 ) );
  INV_X1 u2_uk_U1132 (.ZN( u2_K10_12 ) , .A( u2_uk_n240 ) );
  INV_X1 u2_uk_U1139 (.ZN( u2_K8_43 ) , .A( u2_uk_n1113 ) );
  OAI21_X1 u2_uk_U1140 (.ZN( u2_K16_2 ) , .B2( u2_uk_n1190 ) , .B1( u2_uk_n31 ) , .A( u2_uk_n956 ) );
  INV_X1 u2_uk_U1145 (.ZN( u2_K12_1 ) , .A( u2_uk_n421 ) );
  OAI22_X1 u2_uk_U115 (.ZN( u2_K10_47 ) , .A2( u2_uk_n1594 ) , .B2( u2_uk_n1609 ) , .B1( u2_uk_n164 ) , .A1( u2_uk_n93 ) );
  OAI22_X1 u2_uk_U1150 (.ZN( u2_K1_23 ) , .B2( u2_uk_n1167 ) , .A2( u2_uk_n1174 ) , .A1( u2_uk_n118 ) , .B1( u2_uk_n238 ) );
  INV_X1 u2_uk_U1151 (.A( u2_key_r_33 ) , .ZN( u2_uk_n1167 ) );
  OAI22_X1 u2_uk_U116 (.ZN( u2_K8_47 ) , .B2( u2_uk_n1531 ) , .A2( u2_uk_n1537 ) , .B1( u2_uk_n17 ) , .A1( u2_uk_n223 ) );
  OAI22_X1 u2_uk_U117 (.ZN( u2_K7_47 ) , .A2( u2_uk_n1456 ) , .B2( u2_uk_n1470 ) , .A1( u2_uk_n164 ) , .B1( u2_uk_n31 ) );
  INV_X1 u2_uk_U12 (.A( u2_uk_n145 ) , .ZN( u2_uk_n83 ) );
  OAI22_X1 u2_uk_U125 (.ZN( u2_K4_15 ) , .B2( u2_uk_n1328 ) , .A2( u2_uk_n1356 ) , .A1( u2_uk_n182 ) , .B1( u2_uk_n63 ) );
  OAI21_X1 u2_uk_U126 (.ZN( u2_K5_15 ) , .A( u2_uk_n1042 ) , .B1( u2_uk_n110 ) , .B2( u2_uk_n1379 ) );
  INV_X1 u2_uk_U13 (.A( u2_uk_n182 ) , .ZN( u2_uk_n92 ) );
  OAI22_X1 u2_uk_U130 (.ZN( u2_K7_15 ) , .A2( u2_uk_n1454 ) , .A1( u2_uk_n148 ) , .B2( u2_uk_n1494 ) , .B1( u2_uk_n31 ) );
  INV_X1 u2_uk_U131 (.ZN( u2_K12_15 ) , .A( u2_uk_n409 ) );
  AOI22_X1 u2_uk_U132 (.B2( u2_uk_K_r10_25 ) , .A2( u2_uk_K_r10_34 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n222 ) , .ZN( u2_uk_n409 ) );
  OAI21_X1 u2_uk_U137 (.ZN( u2_K6_19 ) , .A( u2_uk_n1061 ) , .B2( u2_uk_n1414 ) , .B1( u2_uk_n63 ) );
  INV_X1 u2_uk_U14 (.A( u2_uk_n145 ) , .ZN( u2_uk_n94 ) );
  INV_X1 u2_uk_U15 (.A( u2_uk_n164 ) , .ZN( u2_uk_n93 ) );
  OAI22_X1 u2_uk_U153 (.ZN( u2_K7_19 ) , .B2( u2_uk_n1465 ) , .A2( u2_uk_n1475 ) , .A1( u2_uk_n209 ) , .B1( u2_uk_n31 ) );
  OAI21_X1 u2_uk_U154 (.ZN( u2_K3_19 ) , .A( u2_uk_n1007 ) , .B2( u2_uk_n1294 ) , .B1( u2_uk_n83 ) );
  OAI22_X1 u2_uk_U162 (.ZN( u2_K2_30 ) , .B1( u2_uk_n10 ) , .B2( u2_uk_n1230 ) , .A2( u2_uk_n1259 ) , .A1( u2_uk_n162 ) );
  OAI22_X1 u2_uk_U163 (.ZN( u2_K14_30 ) , .B1( u2_uk_n142 ) , .B2( u2_uk_n1781 ) , .A2( u2_uk_n1808 ) , .A1( u2_uk_n94 ) );
  OAI21_X1 u2_uk_U168 (.ZN( u2_K1_14 ) , .B1( u2_uk_n100 ) , .B2( u2_uk_n1160 ) , .A( u2_uk_n970 ) );
  INV_X1 u2_uk_U170 (.A( u2_key_r_25 ) , .ZN( u2_uk_n1160 ) );
  OAI21_X1 u2_uk_U173 (.ZN( u2_K16_30 ) , .B2( u2_uk_n1226 ) , .B1( u2_uk_n187 ) , .A( u2_uk_n957 ) );
  NAND2_X1 u2_uk_U174 (.A1( u2_uk_K_r14_45 ) , .A2( u2_uk_n148 ) , .ZN( u2_uk_n957 ) );
  OAI22_X1 u2_uk_U176 (.ZN( u2_K12_14 ) , .B2( u2_uk_n1688 ) , .A2( u2_uk_n1693 ) , .B1( u2_uk_n214 ) , .A1( u2_uk_n92 ) );
  OAI22_X1 u2_uk_U189 (.ZN( u2_K10_14 ) , .A1( u2_uk_n117 ) , .B2( u2_uk_n1600 ) , .A2( u2_uk_n1631 ) , .B1( u2_uk_n238 ) );
  INV_X1 u2_uk_U19 (.ZN( u2_uk_n100 ) , .A( u2_uk_n146 ) );
  INV_X1 u2_uk_U194 (.ZN( u2_K7_24 ) , .A( u2_uk_n1083 ) );
  AOI22_X1 u2_uk_U195 (.B2( u2_uk_K_r5_18 ) , .A2( u2_uk_K_r5_40 ) , .ZN( u2_uk_n1083 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n208 ) );
  OAI22_X1 u2_uk_U196 (.ZN( u2_K4_24 ) , .A1( u2_uk_n128 ) , .B2( u2_uk_n1322 ) , .A2( u2_uk_n1363 ) , .B1( u2_uk_n142 ) );
  INV_X1 u2_uk_U197 (.ZN( u2_K3_24 ) , .A( u2_uk_n1008 ) );
  AOI22_X1 u2_uk_U198 (.B2( u2_uk_K_r1_17 ) , .A2( u2_uk_K_r1_41 ) , .ZN( u2_uk_n1008 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n202 ) );
  OAI21_X1 u2_uk_U204 (.ZN( u2_K4_30 ) , .A( u2_uk_n1032 ) , .B2( u2_uk_n1345 ) , .B1( u2_uk_n187 ) );
  NAND2_X1 u2_uk_U205 (.A1( u2_uk_K_r2_28 ) , .ZN( u2_uk_n1032 ) , .A2( u2_uk_n148 ) );
  INV_X1 u2_uk_U206 (.ZN( u2_K15_30 ) , .A( u2_uk_n940 ) );
  AOI22_X1 u2_uk_U207 (.B2( u2_uk_K_r13_0 ) , .A2( u2_uk_K_r13_38 ) , .B1( u2_uk_n118 ) , .A1( u2_uk_n207 ) , .ZN( u2_uk_n940 ) );
  OAI22_X1 u2_uk_U208 (.ZN( u2_K3_14 ) , .B1( u2_uk_n10 ) , .B2( u2_uk_n1310 ) , .A2( u2_uk_n1317 ) , .A1( u2_uk_n202 ) );
  INV_X1 u2_uk_U209 (.ZN( u2_K4_31 ) , .A( u2_uk_n1033 ) );
  AOI22_X1 u2_uk_U210 (.B2( u2_uk_K_r2_31 ) , .A2( u2_uk_K_r2_49 ) , .B1( u2_uk_n10 ) , .ZN( u2_uk_n1033 ) , .A1( u2_uk_n188 ) );
  BUF_X1 u2_uk_U22 (.Z( u2_uk_n141 ) , .A( u2_uk_n223 ) );
  OAI22_X1 u2_uk_U228 (.ZN( u2_K3_31 ) , .B1( u2_uk_n110 ) , .B2( u2_uk_n1303 ) , .A2( u2_uk_n1309 ) , .A1( u2_uk_n213 ) );
  OAI22_X1 u2_uk_U235 (.ZN( u2_K14_31 ) , .B1( u2_uk_n142 ) , .B2( u2_uk_n1797 ) , .A2( u2_uk_n1803 ) , .A1( u2_uk_n94 ) );
  OAI22_X1 u2_uk_U242 (.ZN( u2_K16_48 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1200 ) , .A2( u2_uk_n1208 ) , .A1( u2_uk_n213 ) );
  BUF_X1 u2_uk_U25 (.Z( u2_uk_n142 ) , .A( u2_uk_n222 ) );
  OAI22_X1 u2_uk_U261 (.ZN( u2_K10_48 ) , .A1( u2_uk_n148 ) , .B2( u2_uk_n1610 ) , .A2( u2_uk_n1626 ) , .B1( u2_uk_n83 ) );
  OAI21_X1 u2_uk_U264 (.ZN( u2_K8_44 ) , .B1( u2_uk_n102 ) , .A( u2_uk_n1114 ) , .B2( u2_uk_n1538 ) );
  NAND2_X1 u2_uk_U265 (.A1( u2_uk_K_r6_0 ) , .ZN( u2_uk_n1114 ) , .A2( u2_uk_n31 ) );
  OAI22_X1 u2_uk_U266 (.ZN( u2_K8_48 ) , .A2( u2_uk_n1504 ) , .B2( u2_uk_n1511 ) , .B1( u2_uk_n217 ) , .A1( u2_uk_n92 ) );
  OAI22_X1 u2_uk_U267 (.ZN( u2_K7_44 ) , .A1( u2_uk_n118 ) , .B1( u2_uk_n142 ) , .B2( u2_uk_n1459 ) , .A2( u2_uk_n1480 ) );
  BUF_X1 u2_uk_U27 (.Z( u2_uk_n129 ) , .A( u2_uk_n220 ) );
  OAI21_X1 u2_uk_U272 (.ZN( u2_K3_44 ) , .A( u2_uk_n1015 ) , .B1( u2_uk_n109 ) , .B2( u2_uk_n1284 ) );
  NAND2_X1 u2_uk_U273 (.A1( u2_uk_K_r1_15 ) , .ZN( u2_uk_n1015 ) , .A2( u2_uk_n60 ) );
  OAI22_X1 u2_uk_U277 (.ZN( u2_K15_6 ) , .B1( u2_uk_n17 ) , .B2( u2_uk_n1834 ) , .A2( u2_uk_n1852 ) , .A1( u2_uk_n217 ) );
  BUF_X1 u2_uk_U28 (.Z( u2_uk_n146 ) , .A( u2_uk_n182 ) );
  OAI22_X1 u2_uk_U283 (.ZN( u2_K3_6 ) , .A2( u2_uk_n1282 ) , .B2( u2_uk_n1287 ) , .B1( u2_uk_n222 ) , .A1( u2_uk_n92 ) );
  OAI22_X1 u2_uk_U284 (.ZN( u2_K1_8 ) , .A2( u2_uk_n1146 ) , .B2( u2_uk_n1159 ) , .B1( u2_uk_n142 ) , .A1( u2_uk_n94 ) );
  INV_X1 u2_uk_U285 (.ZN( u2_K15_8 ) , .A( u2_uk_n946 ) );
  AOI22_X1 u2_uk_U286 (.B2( u2_uk_K_r13_13 ) , .A2( u2_uk_K_r13_17 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n141 ) , .ZN( u2_uk_n946 ) );
  INV_X1 u2_uk_U289 (.ZN( u2_K7_8 ) , .A( u2_uk_n1096 ) );
  OAI22_X1 u2_uk_U294 (.ZN( u2_K3_8 ) , .A2( u2_uk_n1280 ) , .B2( u2_uk_n1296 ) , .A1( u2_uk_n164 ) , .B1( u2_uk_n94 ) );
  INV_X1 u2_uk_U3 (.ZN( u2_uk_n10 ) , .A( u2_uk_n141 ) );
  BUF_X1 u2_uk_U30 (.Z( u2_uk_n161 ) , .A( u2_uk_n213 ) );
  INV_X1 u2_uk_U303 (.ZN( u2_K4_26 ) , .A( u2_uk_n1028 ) );
  INV_X1 u2_uk_U305 (.ZN( u2_K15_26 ) , .A( u2_uk_n939 ) );
  OAI21_X1 u2_uk_U307 (.ZN( u2_K6_26 ) , .A( u2_uk_n1064 ) , .B2( u2_uk_n1439 ) , .B1( u2_uk_n188 ) );
  NAND2_X1 u2_uk_U308 (.A1( u2_uk_K_r4_35 ) , .ZN( u2_uk_n1064 ) , .A2( u2_uk_n191 ) );
  NAND2_X1 u2_uk_U312 (.A1( u2_uk_K_r11_7 ) , .A2( u2_uk_n10 ) , .ZN( u2_uk_n656 ) );
  OAI22_X1 u2_uk_U314 (.ZN( u2_K2_26 ) , .B2( u2_uk_n1259 ) , .A2( u2_uk_n1265 ) , .B1( u2_uk_n17 ) , .A1( u2_uk_n203 ) );
  OAI22_X1 u2_uk_U316 (.ZN( u2_K14_26 ) , .B2( u2_uk_n1792 ) , .A2( u2_uk_n1809 ) , .A1( u2_uk_n191 ) , .B1( u2_uk_n63 ) );
  OAI21_X1 u2_uk_U326 (.ZN( u2_K3_46 ) , .A( u2_uk_n1017 ) , .B2( u2_uk_n1297 ) , .B1( u2_uk_n202 ) );
  NAND2_X1 u2_uk_U327 (.A1( u2_uk_K_r1_22 ) , .ZN( u2_uk_n1017 ) , .A2( u2_uk_n148 ) );
  BUF_X1 u2_uk_U33 (.Z( u2_uk_n182 ) , .A( u2_uk_n208 ) );
  NAND2_X1 u2_uk_U330 (.A1( u2_key_r_49 ) , .A2( u2_uk_n94 ) , .ZN( u2_uk_n988 ) );
  OAI22_X1 u2_uk_U331 (.ZN( u2_K15_4 ) , .B2( u2_uk_n1820 ) , .A2( u2_uk_n1850 ) , .B1( u2_uk_n208 ) , .A1( u2_uk_n99 ) );
  INV_X1 u2_uk_U338 (.ZN( u2_K12_4 ) , .A( u2_uk_n515 ) );
  AOI22_X1 u2_uk_U339 (.B2( u2_uk_K_r10_27 ) , .A2( u2_uk_K_r10_4 ) , .B1( u2_uk_n10 ) , .A1( u2_uk_n238 ) , .ZN( u2_uk_n515 ) );
  BUF_X1 u2_uk_U34 (.Z( u2_uk_n164 ) , .A( u2_uk_n208 ) );
  OAI22_X1 u2_uk_U342 (.ZN( u2_K3_4 ) , .B2( u2_uk_n1293 ) , .A2( u2_uk_n1301 ) , .A1( u2_uk_n213 ) , .B1( u2_uk_n93 ) );
  OAI21_X1 u2_uk_U344 (.ZN( u2_K1_4 ) , .B2( u2_uk_n1184 ) , .B1( u2_uk_n209 ) , .A( u2_uk_n990 ) );
  NAND2_X1 u2_uk_U345 (.A1( u2_key_r_3 ) , .A2( u2_uk_n207 ) , .ZN( u2_uk_n990 ) );
  INV_X1 u2_uk_U348 (.ZN( u2_K7_46 ) , .A( u2_uk_n1094 ) );
  BUF_X1 u2_uk_U35 (.A( u2_uk_n164 ) , .Z( u2_uk_n187 ) );
  OAI22_X1 u2_uk_U354 (.ZN( u2_K16_40 ) , .B2( u2_uk_n1188 ) , .A2( u2_uk_n1226 ) , .B1( u2_uk_n238 ) , .A1( u2_uk_n94 ) );
  OAI22_X1 u2_uk_U355 (.ZN( u2_K15_40 ) , .A1( u2_uk_n162 ) , .B1( u2_uk_n17 ) , .A2( u2_uk_n1817 ) , .B2( u2_uk_n1849 ) );
  OAI22_X1 u2_uk_U358 (.ZN( u2_K8_40 ) , .B2( u2_uk_n1525 ) , .A2( u2_uk_n1531 ) , .A1( u2_uk_n182 ) , .B1( u2_uk_n93 ) );
  OAI22_X1 u2_uk_U359 (.ZN( u2_K7_40 ) , .A2( u2_uk_n1452 ) , .B2( u2_uk_n1464 ) , .A1( u2_uk_n208 ) , .B1( u2_uk_n31 ) );
  OAI21_X1 u2_uk_U362 (.ZN( u2_K15_33 ) , .B1( u2_uk_n109 ) , .B2( u2_uk_n1840 ) , .A( u2_uk_n942 ) );
  OAI21_X1 u2_uk_U368 (.ZN( u2_K16_28 ) , .B1( u2_uk_n102 ) , .B2( u2_uk_n1189 ) , .A( u2_uk_n954 ) );
  BUF_X1 u2_uk_U37 (.Z( u2_uk_n213 ) , .A( u2_uk_n231 ) );
  OAI22_X1 u2_uk_U372 (.ZN( u2_K6_28 ) , .B2( u2_uk_n1420 ) , .A2( u2_uk_n1447 ) , .A1( u2_uk_n220 ) , .B1( u2_uk_n60 ) );
  BUF_X1 u2_uk_U38 (.Z( u2_uk_n208 ) , .A( u2_uk_n231 ) );
  OAI22_X1 u2_uk_U380 (.ZN( u2_K7_28 ) , .B2( u2_uk_n1471 ) , .A2( u2_uk_n1480 ) , .A1( u2_uk_n223 ) , .B1( u2_uk_n31 ) );
  OAI21_X1 u2_uk_U384 (.ZN( u2_K10_1 ) , .B1( u2_uk_n109 ) , .B2( u2_uk_n1600 ) , .A( u2_uk_n251 ) );
  OAI22_X1 u2_uk_U390 (.ZN( u2_K3_1 ) , .B2( u2_uk_n1285 ) , .A1( u2_uk_n129 ) , .A2( u2_uk_n1290 ) , .B1( u2_uk_n27 ) );
  OAI22_X1 u2_uk_U391 (.ZN( u2_K16_1 ) , .B2( u2_uk_n1218 ) , .A2( u2_uk_n1221 ) , .B1( u2_uk_n17 ) , .A1( u2_uk_n187 ) );
  OAI21_X1 u2_uk_U392 (.ZN( u2_K7_1 ) , .A( u2_uk_n1078 ) , .B2( u2_uk_n1462 ) , .B1( u2_uk_n208 ) );
  NAND2_X1 u2_uk_U393 (.A1( u2_uk_K_r5_10 ) , .ZN( u2_uk_n1078 ) , .A2( u2_uk_n129 ) );
  OAI21_X1 u2_uk_U396 (.ZN( u2_K10_16 ) , .B2( u2_uk_n1630 ) , .B1( u2_uk_n187 ) , .A( u2_uk_n250 ) );
  NAND2_X1 u2_uk_U397 (.A1( u2_uk_K_r8_32 ) , .A2( u2_uk_n230 ) , .ZN( u2_uk_n250 ) );
  INV_X1 u2_uk_U4 (.ZN( u2_uk_n118 ) , .A( u2_uk_n187 ) );
  OAI21_X1 u2_uk_U400 (.ZN( u2_K7_16 ) , .A( u2_uk_n1077 ) , .B1( u2_uk_n110 ) , .B2( u2_uk_n1496 ) );
  OAI22_X1 u2_uk_U403 (.ZN( u2_K4_16 ) , .B2( u2_uk_n1329 ) , .A2( u2_uk_n1333 ) , .A1( u2_uk_n207 ) , .B1( u2_uk_n99 ) );
  OAI21_X1 u2_uk_U407 (.ZN( u2_K15_9 ) , .B1( u2_uk_n109 ) , .B2( u2_uk_n1843 ) , .A( u2_uk_n947 ) );
  OAI22_X1 u2_uk_U412 (.ZN( u2_K12_9 ) , .A1( u2_uk_n100 ) , .B2( u2_uk_n1715 ) , .A2( u2_uk_n1722 ) , .B1( u2_uk_n222 ) );
  INV_X1 u2_uk_U418 (.ZN( u2_K8_37 ) , .A( u2_uk_n1108 ) );
  AOI22_X1 u2_uk_U419 (.B2( u2_uk_K_r6_14 ) , .A2( u2_uk_K_r6_7 ) , .ZN( u2_uk_n1108 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n162 ) );
  BUF_X1 u2_uk_U42 (.A( u2_uk_n182 ) , .Z( u2_uk_n202 ) );
  INV_X1 u2_uk_U420 (.ZN( u2_K10_9 ) , .A( u2_uk_n308 ) );
  AOI22_X1 u2_uk_U421 (.B2( u2_uk_K_r8_17 ) , .A2( u2_uk_K_r8_27 ) , .B1( u2_uk_n118 ) , .A1( u2_uk_n203 ) , .ZN( u2_uk_n308 ) );
  OAI22_X1 u2_uk_U426 (.ZN( u2_K7_9 ) , .B2( u2_uk_n1461 ) , .A2( u2_uk_n1468 ) , .A1( u2_uk_n231 ) , .B1( u2_uk_n31 ) );
  OAI21_X1 u2_uk_U428 (.ZN( u2_K3_9 ) , .A( u2_uk_n1019 ) , .B2( u2_uk_n1295 ) , .B1( u2_uk_n202 ) );
  NAND2_X1 u2_uk_U429 (.A1( u2_uk_K_r1_18 ) , .ZN( u2_uk_n1019 ) , .A2( u2_uk_n217 ) );
  BUF_X1 u2_uk_U43 (.A( u2_uk_n141 ) , .Z( u2_uk_n222 ) );
  INV_X1 u2_uk_U439 (.ZN( u2_K2_28 ) , .A( u2_uk_n998 ) );
  BUF_X1 u2_uk_U44 (.A( u2_uk_n182 ) , .Z( u2_uk_n220 ) );
  AOI22_X1 u2_uk_U440 (.B2( u2_uk_K_r0_15 ) , .A2( u2_uk_K_r0_49 ) , .A1( u2_uk_n102 ) , .B1( u2_uk_n208 ) , .ZN( u2_uk_n998 ) );
  INV_X1 u2_uk_U441 (.ZN( u2_K16_37 ) , .A( u2_uk_n959 ) );
  AOI22_X1 u2_uk_U442 (.B2( u2_uk_K_r14_2 ) , .A2( u2_uk_K_r14_50 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n213 ) , .ZN( u2_uk_n959 ) );
  OAI22_X1 u2_uk_U452 (.ZN( u2_K16_33 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1220 ) , .A2( u2_uk_n1225 ) , .A1( u2_uk_n129 ) );
  OAI22_X1 u2_uk_U453 (.ZN( u2_K14_33 ) , .A1( u2_uk_n155 ) , .B2( u2_uk_n1785 ) , .A2( u2_uk_n1803 ) , .B1( u2_uk_n83 ) );
  OAI22_X1 u2_uk_U459 (.ZN( u2_K3_33 ) , .A1( u2_uk_n128 ) , .B2( u2_uk_n1292 ) , .A2( u2_uk_n1309 ) , .B1( u2_uk_n145 ) );
  OAI22_X1 u2_uk_U460 (.ZN( u2_K15_37 ) , .A2( u2_uk_n1819 ) , .B2( u2_uk_n1846 ) , .A1( u2_uk_n223 ) , .B1( u2_uk_n99 ) );
  OAI22_X1 u2_uk_U471 (.ZN( u2_K3_37 ) , .B2( u2_uk_n1292 ) , .A2( u2_uk_n1298 ) , .A1( u2_uk_n202 ) , .B1( u2_uk_n92 ) );
  NAND2_X1 u2_uk_U474 (.A1( u2_uk_K_r8_21 ) , .A2( u2_uk_n11 ) , .ZN( u2_uk_n298 ) );
  OAI21_X1 u2_uk_U475 (.ZN( u2_K14_29 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1807 ) , .A( u2_uk_n689 ) );
  OAI21_X1 u2_uk_U478 (.ZN( u2_K6_29 ) , .A( u2_uk_n1065 ) , .B2( u2_uk_n1412 ) , .B1( u2_uk_n161 ) );
  NAND2_X1 u2_uk_U479 (.A1( u2_uk_K_r4_0 ) , .ZN( u2_uk_n1065 ) , .A2( u2_uk_n191 ) );
  INV_X1 u2_uk_U481 (.ZN( u2_K16_29 ) , .A( u2_uk_n955 ) );
  INV_X1 u2_uk_U483 (.ZN( u2_K4_29 ) , .A( u2_uk_n1030 ) );
  AOI22_X1 u2_uk_U484 (.B2( u2_uk_K_r2_31 ) , .A2( u2_uk_K_r2_36 ) , .ZN( u2_uk_n1030 ) , .B1( u2_uk_n191 ) , .A1( u2_uk_n83 ) );
  OAI22_X1 u2_uk_U487 (.ZN( u2_K2_29 ) , .A2( u2_uk_n1237 ) , .B2( u2_uk_n1252 ) , .A1( u2_uk_n161 ) , .B1( u2_uk_n27 ) );
  OAI22_X1 u2_uk_U493 (.ZN( u2_K7_29 ) , .B2( u2_uk_n1459 ) , .A2( u2_uk_n1490 ) , .A1( u2_uk_n238 ) , .B1( u2_uk_n31 ) );
  OAI21_X1 u2_uk_U497 (.ZN( u2_K10_2 ) , .B2( u2_uk_n1592 ) , .B1( u2_uk_n220 ) , .A( u2_uk_n286 ) );
  NAND2_X1 u2_uk_U498 (.A1( u2_uk_K_r8_41 ) , .A2( u2_uk_n230 ) , .ZN( u2_uk_n286 ) );
  INV_X1 u2_uk_U5 (.ZN( u2_uk_n117 ) , .A( u2_uk_n161 ) );
  OAI22_X1 u2_uk_U502 (.ZN( u2_K3_2 ) , .B2( u2_uk_n1301 ) , .A2( u2_uk_n1306 ) , .A1( u2_uk_n220 ) , .B1( u2_uk_n83 ) );
  OAI21_X1 u2_uk_U503 (.ZN( u2_K7_2 ) , .B1( u2_uk_n100 ) , .A( u2_uk_n1086 ) , .B2( u2_uk_n1454 ) );
  NAND2_X1 u2_uk_U504 (.A1( u2_uk_K_r5_41 ) , .ZN( u2_uk_n1086 ) , .A2( u2_uk_n63 ) );
  OAI21_X1 u2_uk_U507 (.ZN( u2_K1_12 ) , .B2( u2_uk_n1154 ) , .B1( u2_uk_n93 ) , .A( u2_uk_n968 ) );
  NAND2_X1 u2_uk_U508 (.A1( u2_key_r_12 ) , .A2( u2_uk_n10 ) , .ZN( u2_uk_n968 ) );
  OAI22_X1 u2_uk_U516 (.ZN( u2_K7_17 ) , .B2( u2_uk_n1458 ) , .A2( u2_uk_n1488 ) , .A1( u2_uk_n230 ) , .B1( u2_uk_n31 ) );
  OAI21_X1 u2_uk_U517 (.ZN( u2_K4_17 ) , .A( u2_uk_n1021 ) , .B2( u2_uk_n1339 ) , .B1( u2_uk_n187 ) );
  NAND2_X1 u2_uk_U518 (.A1( u2_uk_K_r2_27 ) , .ZN( u2_uk_n1021 ) , .A2( u2_uk_n155 ) );
  OAI22_X1 u2_uk_U519 (.ZN( u2_K3_17 ) , .B1( u2_uk_n10 ) , .B2( u2_uk_n1287 ) , .A2( u2_uk_n1310 ) , .A1( u2_uk_n202 ) );
  INV_X1 u2_uk_U52 (.ZN( u2_K16_34 ) , .A( u2_uk_n958 ) );
  OAI22_X1 u2_uk_U521 (.ZN( u2_K15_12 ) , .A1( u2_uk_n118 ) , .B1( u2_uk_n142 ) , .A2( u2_uk_n1815 ) , .B2( u2_uk_n1833 ) );
  OAI21_X1 u2_uk_U523 (.ZN( u2_K12_12 ) , .B2( u2_uk_n1689 ) , .B1( u2_uk_n31 ) , .A( u2_uk_n408 ) );
  INV_X1 u2_uk_U525 (.ZN( u2_K7_12 ) , .A( u2_uk_n1075 ) );
  AOI22_X1 u2_uk_U526 (.B2( u2_uk_K_r5_17 ) , .A2( u2_uk_K_r5_39 ) , .ZN( u2_uk_n1075 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n230 ) );
  OAI21_X1 u2_uk_U527 (.ZN( u2_K5_12 ) , .A( u2_uk_n1041 ) , .B2( u2_uk_n1375 ) , .B1( u2_uk_n163 ) );
  NAND2_X1 u2_uk_U528 (.A1( u2_uk_K_r3_11 ) , .ZN( u2_uk_n1041 ) , .A2( u2_uk_n155 ) );
  AOI22_X1 u2_uk_U53 (.B2( u2_uk_K_r14_2 ) , .A2( u2_uk_K_r14_9 ) , .A1( u2_uk_n117 ) , .B1( u2_uk_n238 ) , .ZN( u2_uk_n958 ) );
  OAI22_X1 u2_uk_U530 (.ZN( u2_K3_12 ) , .B1( u2_uk_n10 ) , .B2( u2_uk_n1306 ) , .A2( u2_uk_n1311 ) , .A1( u2_uk_n203 ) );
  INV_X1 u2_uk_U542 (.ZN( u2_K12_17 ) , .A( u2_uk_n415 ) );
  OAI22_X1 u2_uk_U548 (.ZN( u2_K15_36 ) , .B2( u2_uk_n1826 ) , .A2( u2_uk_n1840 ) , .A1( u2_uk_n222 ) , .B1( u2_uk_n92 ) );
  OAI22_X1 u2_uk_U549 (.ZN( u2_K14_36 ) , .A1( u2_uk_n141 ) , .B2( u2_uk_n1770 ) , .A2( u2_uk_n1808 ) , .B1( u2_uk_n63 ) );
  OAI22_X1 u2_uk_U551 (.ZN( u2_K3_36 ) , .B2( u2_uk_n1279 ) , .A1( u2_uk_n128 ) , .A2( u2_uk_n1314 ) , .B1( u2_uk_n145 ) );
  OAI22_X1 u2_uk_U563 (.ZN( u2_K16_36 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1203 ) , .A2( u2_uk_n1210 ) , .A1( u2_uk_n129 ) );
  INV_X1 u2_uk_U564 (.ZN( u2_K15_38 ) , .A( u2_uk_n943 ) );
  OAI21_X1 u2_uk_U571 (.ZN( u2_K15_10 ) , .B1( u2_uk_n109 ) , .B2( u2_uk_n1839 ) , .A( u2_uk_n934 ) );
  NAND2_X1 u2_uk_U572 (.A1( u2_uk_K_r13_55 ) , .A2( u2_uk_n11 ) , .ZN( u2_uk_n934 ) );
  INV_X1 u2_uk_U584 (.ZN( u2_K1_10 ) , .A( u2_uk_n966 ) );
  AOI22_X1 u2_uk_U585 (.B2( u2_key_r_41 ) , .A2( u2_key_r_48 ) , .B1( u2_uk_n118 ) , .A1( u2_uk_n161 ) , .ZN( u2_uk_n966 ) );
  OAI22_X1 u2_uk_U587 (.ZN( u2_K3_22 ) , .B2( u2_uk_n1281 ) , .A2( u2_uk_n1316 ) , .B1( u2_uk_n141 ) , .A1( u2_uk_n94 ) );
  OAI21_X1 u2_uk_U598 (.ZN( u2_K7_22 ) , .B1( u2_uk_n100 ) , .A( u2_uk_n1081 ) , .B2( u2_uk_n1468 ) );
  INV_X1 u2_uk_U600 (.ZN( u2_K5_22 ) , .A( u2_uk_n1044 ) );
  INV_X1 u2_uk_U602 (.ZN( u2_K1_22 ) , .A( u2_uk_n974 ) );
  AOI22_X1 u2_uk_U603 (.B2( u2_key_r_25 ) , .A2( u2_key_r_32 ) , .B1( u2_uk_n109 ) , .A1( u2_uk_n191 ) , .ZN( u2_uk_n974 ) );
  OAI22_X1 u2_uk_U604 (.ZN( u2_K16_35 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1208 ) , .A2( u2_uk_n1215 ) , .A1( u2_uk_n129 ) );
  NAND2_X1 u2_uk_U608 (.A1( u2_uk_K_r5_37 ) , .ZN( u2_uk_n1090 ) , .A2( u2_uk_n11 ) );
  INV_X1 u2_uk_U61 (.ZN( u2_K14_34 ) , .A( u2_uk_n692 ) );
  INV_X1 u2_uk_U612 (.ZN( u2_K14_35 ) , .A( u2_uk_n694 ) );
  AOI22_X1 u2_uk_U613 (.B2( u2_uk_K_r12_1 ) , .A2( u2_uk_K_r12_7 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n142 ) , .ZN( u2_uk_n694 ) );
  AOI22_X1 u2_uk_U62 (.B2( u2_uk_K_r12_30 ) , .A2( u2_uk_K_r12_36 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n213 ) , .ZN( u2_uk_n692 ) );
  OAI22_X1 u2_uk_U625 (.ZN( u2_K7_11 ) , .B2( u2_uk_n1458 ) , .A2( u2_uk_n1475 ) , .B1( u2_uk_n208 ) , .A1( u2_uk_n93 ) );
  OAI21_X1 u2_uk_U626 (.ZN( u2_K15_11 ) , .B2( u2_uk_n1850 ) , .B1( u2_uk_n231 ) , .A( u2_uk_n935 ) );
  NAND2_X1 u2_uk_U627 (.A1( u2_uk_K_r13_25 ) , .A2( u2_uk_n207 ) , .ZN( u2_uk_n935 ) );
  OAI22_X1 u2_uk_U639 (.ZN( u2_K3_11 ) , .A2( u2_uk_n1280 ) , .B2( u2_uk_n1285 ) , .B1( u2_uk_n141 ) , .A1( u2_uk_n99 ) );
  OAI21_X1 u2_uk_U646 (.ZN( u2_K12_6 ) , .B1( u2_uk_n162 ) , .B2( u2_uk_n1702 ) , .A( u2_uk_n518 ) );
  NAND2_X1 u2_uk_U647 (.A1( u2_uk_K_r10_10 ) , .A2( u2_uk_n148 ) , .ZN( u2_uk_n518 ) );
  OAI22_X1 u2_uk_U648 (.ZN( u2_K16_45 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1217 ) , .A2( u2_uk_n1220 ) , .A1( u2_uk_n238 ) );
  OAI22_X1 u2_uk_U658 (.ZN( u2_K1_7 ) , .B2( u2_uk_n1155 ) , .A2( u2_uk_n1162 ) , .B1( u2_uk_n142 ) , .A1( u2_uk_n94 ) );
  INV_X1 u2_uk_U661 (.ZN( u2_K16_43 ) , .A( u2_uk_n963 ) );
  AOI22_X1 u2_uk_U662 (.B2( u2_uk_K_r14_16 ) , .A2( u2_uk_K_r14_9 ) , .B1( u2_uk_n118 ) , .A1( u2_uk_n161 ) , .ZN( u2_uk_n963 ) );
  OAI21_X1 u2_uk_U67 (.ZN( u2_K3_34 ) , .A( u2_uk_n1011 ) , .B1( u2_uk_n110 ) , .B2( u2_uk_n1299 ) );
  OAI22_X1 u2_uk_U673 (.ZN( u2_K10_45 ) , .B2( u2_uk_n1598 ) , .A2( u2_uk_n1614 ) , .A1( u2_uk_n223 ) , .B1( u2_uk_n83 ) );
  OAI22_X1 u2_uk_U676 (.ZN( u2_K16_3 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1198 ) , .A2( u2_uk_n1206 ) , .A1( u2_uk_n191 ) );
  OAI22_X1 u2_uk_U679 (.ZN( u2_K10_7 ) , .B2( u2_uk_n1604 ) , .A2( u2_uk_n1624 ) , .A1( u2_uk_n188 ) , .B1( u2_uk_n83 ) );
  OAI21_X1 u2_uk_U682 (.ZN( u2_K3_3 ) , .A( u2_uk_n1013 ) , .B2( u2_uk_n1318 ) , .B1( u2_uk_n231 ) );
  NAND2_X1 u2_uk_U683 (.A1( u2_uk_K_r1_47 ) , .ZN( u2_uk_n1013 ) , .A2( u2_uk_n214 ) );
  OAI22_X1 u2_uk_U684 (.ZN( u2_K15_7 ) , .A1( u2_uk_n163 ) , .B1( u2_uk_n17 ) , .B2( u2_uk_n1823 ) , .A2( u2_uk_n1839 ) );
  OAI21_X1 u2_uk_U692 (.ZN( u2_K2_25 ) , .B1( u2_uk_n110 ) , .B2( u2_uk_n1264 ) , .A( u2_uk_n996 ) );
  OAI21_X1 u2_uk_U699 (.ZN( u2_K5_7 ) , .A( u2_uk_n1057 ) , .B2( u2_uk_n1405 ) , .B1( u2_uk_n214 ) );
  INV_X1 u2_uk_U7 (.ZN( u2_uk_n11 ) , .A( u2_uk_n141 ) );
  NAND2_X1 u2_uk_U700 (.A1( u2_uk_K_r3_19 ) , .ZN( u2_uk_n1057 ) , .A2( u2_uk_n217 ) );
  INV_X1 u2_uk_U701 (.ZN( u2_K7_25 ) , .A( u2_uk_n1084 ) );
  AOI22_X1 u2_uk_U702 (.B2( u2_uk_K_r5_31 ) , .A2( u2_uk_K_r5_7 ) , .A1( u2_uk_n10 ) , .ZN( u2_uk_n1084 ) , .B1( u2_uk_n217 ) );
  INV_X1 u2_uk_U705 (.ZN( u2_K4_25 ) , .A( u2_uk_n1027 ) );
  OAI21_X1 u2_uk_U707 (.ZN( u2_K15_25 ) , .B1( u2_uk_n146 ) , .B2( u2_uk_n1846 ) , .A( u2_uk_n938 ) );
  NAND2_X1 u2_uk_U708 (.A1( u2_uk_K_r13_22 ) , .A2( u2_uk_n214 ) , .ZN( u2_uk_n938 ) );
  OAI22_X1 u2_uk_U709 (.ZN( u2_K16_25 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1209 ) , .A2( u2_uk_n1216 ) , .A1( u2_uk_n208 ) );
  OAI21_X1 u2_uk_U711 (.ZN( u2_K1_2 ) , .B2( u2_uk_n1145 ) , .B1( u2_uk_n220 ) , .A( u2_uk_n978 ) );
  NAND2_X1 u2_uk_U712 (.A1( u2_key_r_11 ) , .A2( u2_uk_n191 ) , .ZN( u2_uk_n978 ) );
  OAI22_X1 u2_uk_U713 (.ZN( u2_K4_32 ) , .A1( u2_uk_n109 ) , .A2( u2_uk_n1326 ) , .B2( u2_uk_n1350 ) , .B1( u2_uk_n209 ) );
  OAI22_X1 u2_uk_U714 (.ZN( u2_K16_32 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1201 ) , .A2( u2_uk_n1209 ) , .A1( u2_uk_n202 ) );
  OAI22_X1 u2_uk_U723 (.ZN( u2_K14_32 ) , .A1( u2_uk_n155 ) , .B2( u2_uk_n1769 ) , .A2( u2_uk_n1807 ) , .B1( u2_uk_n83 ) );
  OAI22_X1 u2_uk_U727 (.ZN( u2_K15_42 ) , .B1( u2_uk_n161 ) , .B2( u2_uk_n1849 ) , .A2( u2_uk_n1855 ) , .A1( u2_uk_n31 ) );
  OAI21_X1 u2_uk_U732 (.ZN( u2_K8_42 ) , .A( u2_uk_n1112 ) , .B2( u2_uk_n1510 ) , .B1( u2_uk_n17 ) );
  OAI22_X1 u2_uk_U736 (.ZN( u2_K2_42 ) , .B2( u2_uk_n1266 ) , .A2( u2_uk_n1274 ) , .A1( u2_uk_n209 ) , .B1( u2_uk_n60 ) );
  INV_X1 u2_uk_U737 (.ZN( u2_K7_42 ) , .A( u2_uk_n1093 ) );
  OAI21_X1 u2_uk_U741 (.ZN( u2_K14_27 ) , .B1( u2_uk_n100 ) , .B2( u2_uk_n1809 ) , .A( u2_uk_n688 ) );
  NAND2_X1 u2_uk_U742 (.A1( u2_uk_K_r12_42 ) , .A2( u2_uk_n31 ) , .ZN( u2_uk_n688 ) );
  OAI22_X1 u2_uk_U747 (.ZN( u2_K16_27 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1195 ) , .A2( u2_uk_n1200 ) , .A1( u2_uk_n182 ) );
  OAI22_X1 u2_uk_U748 (.ZN( u2_K12_13 ) , .B2( u2_uk_n1689 ) , .A2( u2_uk_n1721 ) , .B1( u2_uk_n209 ) , .A1( u2_uk_n92 ) );
  OAI22_X1 u2_uk_U753 (.ZN( u2_K1_21 ) , .B2( u2_uk_n1153 ) , .A2( u2_uk_n1159 ) , .B1( u2_uk_n214 ) , .A1( u2_uk_n83 ) );
  INV_X1 u2_uk_U76 (.ZN( u2_K4_23 ) , .A( u2_uk_n1026 ) );
  OAI22_X1 u2_uk_U767 (.ZN( u2_K15_27 ) , .A2( u2_uk_n1817 ) , .B2( u2_uk_n1835 ) , .B1( u2_uk_n222 ) , .A1( u2_uk_n99 ) );
  INV_X1 u2_uk_U768 (.ZN( u2_K2_27 ) , .A( u2_uk_n997 ) );
  AOI22_X1 u2_uk_U77 (.B2( u2_uk_K_r2_18 ) , .A2( u2_uk_K_r2_55 ) , .ZN( u2_uk_n1026 ) , .B1( u2_uk_n191 ) , .A1( u2_uk_n83 ) );
  OAI22_X1 u2_uk_U775 (.ZN( u2_K4_13 ) , .A1( u2_uk_n102 ) , .A2( u2_uk_n1324 ) , .B2( u2_uk_n1328 ) , .B1( u2_uk_n230 ) );
  INV_X1 u2_uk_U778 (.ZN( u2_K6_21 ) , .A( u2_uk_n1062 ) );
  AOI22_X1 u2_uk_U779 (.B2( u2_uk_K_r4_11 ) , .A2( u2_uk_K_r4_5 ) , .ZN( u2_uk_n1062 ) , .B1( u2_uk_n118 ) , .A1( u2_uk_n217 ) );
  OAI21_X1 u2_uk_U782 (.ZN( u2_K7_21 ) , .A( u2_uk_n1080 ) , .B2( u2_uk_n1496 ) , .B1( u2_uk_n231 ) );
  NAND2_X1 u2_uk_U783 (.A1( u2_uk_K_r5_19 ) , .ZN( u2_uk_n1080 ) , .A2( u2_uk_n129 ) );
  INV_X1 u2_uk_U789 (.ZN( u2_K7_27 ) , .A( u2_uk_n1085 ) );
  AOI22_X1 u2_uk_U790 (.B2( u2_uk_K_r5_23 ) , .A2( u2_uk_K_r5_43 ) , .ZN( u2_uk_n1085 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n141 ) );
  OAI21_X1 u2_uk_U799 (.ZN( u2_K4_18 ) , .B1( u2_uk_n10 ) , .A( u2_uk_n1022 ) , .B2( u2_uk_n1348 ) );
  OAI21_X1 u2_uk_U80 (.ZN( u2_K16_41 ) , .B2( u2_uk_n1215 ) , .B1( u2_uk_n31 ) , .A( u2_uk_n961 ) );
  OAI22_X1 u2_uk_U802 (.ZN( u2_K7_18 ) , .A2( u2_uk_n1453 ) , .B2( u2_uk_n1466 ) , .A1( u2_uk_n223 ) , .B1( u2_uk_n31 ) );
  NAND2_X1 u2_uk_U806 (.A1( u2_uk_K_r6_46 ) , .ZN( u2_uk_n1102 ) , .A2( u2_uk_n17 ) );
  OAI22_X1 u2_uk_U810 (.ZN( u2_K10_18 ) , .A1( u2_uk_n110 ) , .A2( u2_uk_n1590 ) , .B2( u2_uk_n1604 ) , .B1( u2_uk_n208 ) );
  INV_X1 u2_uk_U826 (.ZN( u2_K7_20 ) , .A( u2_uk_n1079 ) );
  INV_X1 u2_uk_U831 (.ZN( u2_K12_3 ) , .A( u2_uk_n500 ) );
  OAI22_X1 u2_uk_U838 (.ZN( u2_K1_6 ) , .B2( u2_uk_n1168 ) , .A2( u2_uk_n1175 ) , .B1( u2_uk_n145 ) , .A1( u2_uk_n94 ) );
  INV_X1 u2_uk_U839 (.A( u2_key_r_41 ) , .ZN( u2_uk_n1175 ) );
  OAI22_X1 u2_uk_U844 (.ZN( u2_K1_1 ) , .A1( u2_uk_n11 ) , .B2( u2_uk_n1174 ) , .A2( u2_uk_n1179 ) , .B1( u2_uk_n182 ) );
  OAI22_X1 u2_uk_U845 (.ZN( u2_K3_18 ) , .B1( u2_uk_n10 ) , .B2( u2_uk_n1295 ) , .A2( u2_uk_n1302 ) , .A1( u2_uk_n220 ) );
  OAI22_X1 u2_uk_U847 (.ZN( u2_K10_5 ) , .B2( u2_uk_n1595 ) , .A2( u2_uk_n1612 ) , .A1( u2_uk_n231 ) , .B1( u2_uk_n83 ) );
  OAI22_X1 u2_uk_U859 (.ZN( u2_K12_10 ) , .B1( u2_uk_n10 ) , .B2( u2_uk_n1688 ) , .A2( u2_uk_n1709 ) , .A1( u2_uk_n207 ) );
  INV_X1 u2_uk_U86 (.ZN( u2_K2_41 ) , .A( u2_uk_n1001 ) );
  OAI22_X1 u2_uk_U860 (.ZN( u2_K12_11 ) , .A1( u2_uk_n146 ) , .A2( u2_uk_n1683 ) , .B2( u2_uk_n1709 ) , .B1( u2_uk_n63 ) );
  OAI22_X1 u2_uk_U861 (.ZN( u2_K7_10 ) , .B2( u2_uk_n1457 ) , .A2( u2_uk_n1487 ) , .A1( u2_uk_n209 ) , .B1( u2_uk_n60 ) );
  OAI22_X1 u2_uk_U863 (.ZN( u2_K3_10 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1286 ) , .A1( u2_uk_n129 ) , .A2( u2_uk_n1291 ) );
  OAI22_X1 u2_uk_U869 (.ZN( u2_K15_3 ) , .B1( u2_uk_n17 ) , .B2( u2_uk_n1822 ) , .A2( u2_uk_n1838 ) , .A1( u2_uk_n231 ) );
  OAI22_X1 u2_uk_U871 (.ZN( u2_K10_3 ) , .A1( u2_uk_n148 ) , .B2( u2_uk_n1603 ) , .A2( u2_uk_n1623 ) , .B1( u2_uk_n63 ) );
  OAI22_X1 u2_uk_U875 (.ZN( u2_K7_14 ) , .B2( u2_uk_n1462 ) , .A2( u2_uk_n1497 ) , .A1( u2_uk_n222 ) , .B1( u2_uk_n31 ) );
  OAI22_X1 u2_uk_U88 (.ZN( u2_K15_41 ) , .B1( u2_uk_n17 ) , .B2( u2_uk_n1835 ) , .A2( u2_uk_n1853 ) , .A1( u2_uk_n231 ) );
  OAI22_X1 u2_uk_U880 (.ZN( u2_K3_21 ) , .B1( u2_uk_n109 ) , .B2( u2_uk_n1291 ) , .A2( u2_uk_n1316 ) , .A1( u2_uk_n161 ) );
  OAI22_X1 u2_uk_U888 (.ZN( u2_K7_30 ) , .B2( u2_uk_n1460 ) , .A2( u2_uk_n1491 ) , .A1( u2_uk_n182 ) , .B1( u2_uk_n31 ) );
  OAI22_X1 u2_uk_U893 (.ZN( u2_K4_36 ) , .B1( u2_uk_n109 ) , .B2( u2_uk_n1346 ) , .A2( u2_uk_n1351 ) , .A1( u2_uk_n161 ) );
  OAI22_X1 u2_uk_U895 (.ZN( u2_K6_30 ) , .B2( u2_uk_n1408 ) , .A2( u2_uk_n1413 ) , .A1( u2_uk_n164 ) , .B1( u2_uk_n60 ) );
  OAI22_X1 u2_uk_U897 (.ZN( u2_K16_38 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1210 ) , .A2( u2_uk_n1217 ) , .A1( u2_uk_n161 ) );
  OAI22_X1 u2_uk_U898 (.ZN( u2_K8_38 ) , .B1( u2_uk_n118 ) , .B2( u2_uk_n1530 ) , .A2( u2_uk_n1536 ) , .A1( u2_uk_n163 ) );
  OAI22_X1 u2_uk_U899 (.ZN( u2_K7_39 ) , .B2( u2_uk_n1486 ) , .A2( u2_uk_n1493 ) , .A1( u2_uk_n161 ) , .B1( u2_uk_n31 ) );
  INV_X1 u2_uk_U9 (.A( u2_uk_n129 ) , .ZN( u2_uk_n31 ) );
  OAI22_X1 u2_uk_U90 (.ZN( u2_K7_41 ) , .A1( u2_uk_n118 ) , .A2( u2_uk_n1456 ) , .B2( u2_uk_n1486 ) , .B1( u2_uk_n208 ) );
  OAI22_X1 u2_uk_U903 (.ZN( u2_K3_38 ) , .B1( u2_uk_n128 ) , .A2( u2_uk_n1284 ) , .A1( u2_uk_n129 ) , .B2( u2_uk_n1300 ) );
  OAI22_X1 u2_uk_U904 (.ZN( u2_K3_39 ) , .B1( u2_uk_n118 ) , .B2( u2_uk_n1308 ) , .A2( u2_uk_n1312 ) , .A1( u2_uk_n202 ) );
  OAI22_X1 u2_uk_U905 (.ZN( u2_K2_39 ) , .B1( u2_uk_n11 ) , .A2( u2_uk_n1236 ) , .B2( u2_uk_n1251 ) , .A1( u2_uk_n164 ) );
  OAI22_X1 u2_uk_U910 (.ZN( u2_K12_16 ) , .A2( u2_uk_n1681 ) , .B2( u2_uk_n1693 ) , .B1( u2_uk_n209 ) , .A1( u2_uk_n92 ) );
  OAI22_X1 u2_uk_U916 (.ZN( u2_K12_18 ) , .A2( u2_uk_n1683 ) , .B2( u2_uk_n1721 ) , .B1( u2_uk_n231 ) , .A1( u2_uk_n92 ) );
  OAI22_X1 u2_uk_U922 (.ZN( u2_K16_46 ) , .B2( u2_uk_n1189 ) , .A2( u2_uk_n1223 ) , .B1( u2_uk_n217 ) , .A1( u2_uk_n94 ) );
  OAI22_X1 u2_uk_U933 (.ZN( u2_K10_8 ) , .A2( u2_uk_n1591 ) , .B2( u2_uk_n1605 ) , .B1( u2_uk_n161 ) , .A1( u2_uk_n93 ) );
  OAI22_X1 u2_uk_U937 (.ZN( u2_K4_19 ) , .B2( u2_uk_n1335 ) , .A2( u2_uk_n1347 ) , .B1( u2_uk_n223 ) , .A1( u2_uk_n63 ) );
  OAI22_X1 u2_uk_U945 (.ZN( u2_K2_38 ) , .B2( u2_uk_n1246 ) , .A2( u2_uk_n1265 ) , .B1( u2_uk_n129 ) , .A1( u2_uk_n92 ) );
  OAI22_X1 u2_uk_U947 (.ZN( u2_K2_37 ) , .A2( u2_uk_n1237 ) , .B2( u2_uk_n1264 ) , .B1( u2_uk_n129 ) , .A1( u2_uk_n93 ) );
  OAI22_X1 u2_uk_U967 (.ZN( u2_K1_3 ) , .B2( u2_uk_n1154 ) , .A2( u2_uk_n1161 ) , .A1( u2_uk_n118 ) , .B1( u2_uk_n207 ) );
  OAI21_X1 u2_uk_U977 (.ZN( u2_K7_23 ) , .B1( u2_uk_n100 ) , .A( u2_uk_n1082 ) , .B2( u2_uk_n1453 ) );
  OAI21_X1 u2_uk_U979 (.ZN( u2_K6_23 ) , .A( u2_uk_n1063 ) , .B1( u2_uk_n110 ) , .B2( u2_uk_n1442 ) );
  OAI22_X1 u2_uk_U98 (.ZN( u2_K12_5 ) , .A2( u2_uk_n1682 ) , .B2( u2_uk_n1708 ) , .A1( u2_uk_n202 ) , .B1( u2_uk_n94 ) );
  NAND2_X1 u2_uk_U982 (.A1( u2_uk_K_r1_7 ) , .ZN( u2_uk_n1012 ) , .A2( u2_uk_n92 ) );
  OAI21_X1 u2_uk_U987 (.ZN( u2_K16_4 ) , .B1( u2_uk_n100 ) , .B2( u2_uk_n1227 ) , .A( u2_uk_n965 ) );
  NAND2_X1 u2_uk_U988 (.A1( u2_uk_K_r14_3 ) , .A2( u2_uk_n92 ) , .ZN( u2_uk_n965 ) );
  OAI21_X1 u2_uk_U993 (.ZN( u2_K3_5 ) , .B1( u2_uk_n100 ) , .A( u2_uk_n1018 ) , .B2( u2_uk_n1302 ) );
  OAI21_X1 u2_uk_U997 (.ZN( u2_K3_45 ) , .A( u2_uk_n1016 ) , .B1( u2_uk_n102 ) , .B2( u2_uk_n1305 ) );
  NAND2_X1 u2_uk_U998 (.A1( u2_uk_K_r1_16 ) , .ZN( u2_uk_n1016 ) , .A2( u2_uk_n27 ) );
  OAI21_X1 u2_uk_U999 (.ZN( u2_K1_13 ) , .B1( u2_uk_n100 ) , .B2( u2_uk_n1184 ) , .A( u2_uk_n969 ) );
endmodule

