module des_des_die_9 ( n116, u0_K2_44, u0_K2_45, u0_K2_46, u0_K2_47, u0_K2_48, u0_K3_34, u0_L0_15, u0_L0_21, 
       u0_L0_27, u0_L0_5, u0_L13_1, u0_L13_10, u0_L13_20, u0_L13_26, u0_L1_11, u0_L1_14, u0_L1_19, 
       u0_L1_25, u0_L1_29, u0_L1_3, u0_L1_4, u0_L1_8, u0_L9_17, u0_L9_23, u0_L9_31, u0_L9_9, 
       u0_R0_1, u0_R0_28, u0_R0_29, u0_R0_30, u0_R0_31, u0_R0_32, u0_R13_12, u0_R13_13, u0_R13_14, 
       u0_R13_15, u0_R13_16, u0_R13_17, u0_R1_16, u0_R1_17, u0_R1_18, u0_R1_19, u0_R1_20, u0_R1_21, 
       u0_R1_22, u0_R1_23, u0_R1_24, u0_R1_25, u0_R9_1, u0_R9_2, u0_R9_3, u0_R9_32, u0_R9_4, 
       u0_R9_5, u0_uk_K_r0_2, u0_uk_K_r1_42, u0_uk_K_r1_44, u0_uk_K_r1_7, u0_uk_K_r9_19, u0_uk_K_r9_25, u0_uk_n109, u0_uk_n11, 
       u0_uk_n118, u0_uk_n129, u0_uk_n14, u0_uk_n141, u0_uk_n142, u0_uk_n148, u0_uk_n16, u0_uk_n163, u0_uk_n164, 
       u0_uk_n181, u0_uk_n183, u0_uk_n187, u0_uk_n188, u0_uk_n189, u0_uk_n191, u0_uk_n195, u0_uk_n200, u0_uk_n201, 
       u0_uk_n202, u0_uk_n209, u0_uk_n215, u0_uk_n219, u0_uk_n220, u0_uk_n222, u0_uk_n231, u0_uk_n238, u0_uk_n24, 
       u0_uk_n242, u0_uk_n25, u0_uk_n252, u0_uk_n30, u0_uk_n37, u0_uk_n38, u0_uk_n42, u0_uk_n43, u0_uk_n543, 
       u0_uk_n544, u0_uk_n545, u0_uk_n549, u0_uk_n555, u0_uk_n559, u0_uk_n560, u0_uk_n566, u0_uk_n570, u0_uk_n575, 
       u0_uk_n579, u0_uk_n580, u0_uk_n60, u0_uk_n612, u0_uk_n63, u0_uk_n7, u0_uk_n83, u0_uk_n92, u0_uk_n93, 
       u0_uk_n94, u1_FP_33, u1_FP_48, u1_FP_49, u1_FP_50, u1_FP_51, u1_FP_52, u1_FP_53, u1_FP_54, 
       u1_FP_55, u1_FP_56, u1_FP_57, u1_FP_58, u1_FP_59, u1_FP_60, u1_FP_61, u1_FP_62, u1_FP_63, 
       u1_FP_64, u1_L0_17, u1_L0_23, u1_L0_31, u1_L0_9, u1_L10_17, u1_L10_23, u1_L10_31, u1_L10_9, 
       u1_L13_1, u1_L13_10, u1_L13_13, u1_L13_14, u1_L13_16, u1_L13_17, u1_L13_18, u1_L13_2, u1_L13_20, 
       u1_L13_23, u1_L13_24, u1_L13_25, u1_L13_26, u1_L13_28, u1_L13_3, u1_L13_30, u1_L13_31, u1_L13_6, 
       u1_L13_8, u1_L13_9, u1_L14_11, u1_L14_12, u1_L14_14, u1_L14_15, u1_L14_19, u1_L14_21, u1_L14_22, 
       u1_L14_25, u1_L14_27, u1_L14_29, u1_L14_3, u1_L14_32, u1_L14_4, u1_L14_5, u1_L14_7, u1_L14_8, 
       u1_L2_11, u1_L2_12, u1_L2_19, u1_L2_22, u1_L2_29, u1_L2_32, u1_L2_4, u1_L2_7, u1_L3_14, 
       u1_L3_15, u1_L3_21, u1_L3_25, u1_L3_27, u1_L3_3, u1_L3_5, u1_L3_8, u1_L5_12, u1_L5_13, 
       u1_L5_15, u1_L5_16, u1_L5_18, u1_L5_2, u1_L5_21, u1_L5_22, u1_L5_24, u1_L5_27, u1_L5_28, 
       u1_L5_30, u1_L5_32, u1_L5_5, u1_L5_6, u1_L5_7, u1_L6_13, u1_L6_16, u1_L6_17, u1_L6_18, 
       u1_L6_2, u1_L6_23, u1_L6_24, u1_L6_28, u1_L6_30, u1_L6_31, u1_L6_6, u1_L6_9, u1_L7_15, 
       u1_L7_21, u1_L7_27, u1_L7_5, u1_L9_12, u1_L9_22, u1_L9_32, u1_L9_7, u1_R0_1, u1_R0_2, 
       u1_R0_3, u1_R0_32, u1_R0_4, u1_R0_5, u1_R10_1, u1_R10_2, u1_R10_3, u1_R10_32, u1_R10_4, 
       u1_R10_5, u1_R13_1, u1_R13_10, u1_R13_11, u1_R13_12, u1_R13_13, u1_R13_14, u1_R13_15, u1_R13_16, 
       u1_R13_17, u1_R13_18, u1_R13_19, u1_R13_2, u1_R13_20, u1_R13_21, u1_R13_3, u1_R13_32, u1_R13_4, 
       u1_R13_5, u1_R13_6, u1_R13_7, u1_R13_8, u1_R13_9, u1_R2_20, u1_R2_21, u1_R2_22, u1_R2_23, 
       u1_R2_24, u1_R2_25, u1_R2_26, u1_R2_27, u1_R2_28, u1_R2_29, u1_R3_1, u1_R3_16, u1_R3_17, 
       u1_R3_18, u1_R3_19, u1_R3_20, u1_R3_21, u1_R3_28, u1_R3_29, u1_R3_30, u1_R3_31, u1_R3_32, 
       u1_R5_1, u1_R5_10, u1_R5_11, u1_R5_12, u1_R5_13, u1_R5_24, u1_R5_25, u1_R5_26, u1_R5_27, 
       u1_R5_28, u1_R5_29, u1_R5_30, u1_R5_31, u1_R5_32, u1_R5_4, u1_R5_5, u1_R5_6, u1_R5_7, 
       u1_R5_8, u1_R5_9, u1_R6_1, u1_R6_10, u1_R6_11, u1_R6_12, u1_R6_13, u1_R6_2, u1_R6_3, 
       u1_R6_32, u1_R6_4, u1_R6_5, u1_R6_6, u1_R6_7, u1_R6_8, u1_R6_9, u1_R7_1, u1_R7_28, 
       u1_R7_29, u1_R7_30, u1_R7_31, u1_R7_32, u1_R9_24, u1_R9_25, u1_R9_26, u1_R9_27, u1_R9_28, 
       u1_R9_29, u1_uk_K_r10_10, u1_uk_K_r10_18, u1_uk_K_r10_27, u1_uk_K_r10_39, u1_uk_K_r10_4, u1_uk_K_r10_48, u1_uk_K_r13_0, u1_uk_K_r13_13, 
       u1_uk_K_r13_17, u1_uk_K_r13_19, u1_uk_K_r13_22, u1_uk_K_r13_25, u1_uk_K_r13_32, u1_uk_K_r13_38, u1_uk_K_r13_4, u1_uk_K_r13_44, u1_uk_K_r13_55, 
       u1_uk_K_r14_15, u1_uk_K_r14_16, u1_uk_K_r14_2, u1_uk_K_r14_23, u1_uk_K_r14_38, u1_uk_K_r14_42, u1_uk_K_r14_43, u1_uk_K_r14_45, u1_uk_K_r14_50, 
       u1_uk_K_r14_8, u1_uk_K_r14_9, u1_uk_K_r2_31, u1_uk_K_r2_49, u1_uk_K_r2_50, u1_uk_K_r3_15, u1_uk_K_r3_35, u1_uk_K_r3_38, u1_uk_K_r3_43, 
       u1_uk_K_r3_51, u1_uk_K_r5_1, u1_uk_K_r5_17, u1_uk_K_r5_23, u1_uk_K_r5_26, u1_uk_K_r5_31, u1_uk_K_r5_32, u1_uk_K_r5_36, u1_uk_K_r5_39, 
       u1_uk_K_r5_4, u1_uk_K_r5_48, u1_uk_K_r5_8, u1_uk_K_r6_10, u1_uk_K_r6_17, u1_uk_K_r6_19, u1_uk_K_r6_26, u1_uk_K_r6_27, u1_uk_K_r6_3, 
       u1_uk_K_r6_34, u1_uk_K_r6_46, u1_uk_K_r6_53, u1_uk_K_r6_55, u1_uk_K_r7_0, u1_uk_K_r7_16, u1_uk_K_r7_37, u1_uk_K_r7_9, u1_uk_K_r9_30, 
       u1_uk_K_r9_31, u1_uk_K_r9_38, u1_uk_K_r9_7, u1_uk_n102, u1_uk_n109, u1_uk_n11, u1_uk_n117, u1_uk_n118, u1_uk_n1218, 
       u1_uk_n1219, u1_uk_n1222, u1_uk_n1225, u1_uk_n1230, u1_uk_n1231, u1_uk_n1233, u1_uk_n1238, u1_uk_n1239, u1_uk_n1240, 
       u1_uk_n1241, u1_uk_n1245, u1_uk_n1246, u1_uk_n1247, u1_uk_n1250, u1_uk_n1253, u1_uk_n1255, u1_uk_n1256, u1_uk_n1268, 
       u1_uk_n1269, u1_uk_n1273, u1_uk_n1274, u1_uk_n1277, u1_uk_n1279, u1_uk_n1284, u1_uk_n129, u1_uk_n1297, u1_uk_n1300, 
       u1_uk_n1305, u1_uk_n1349, u1_uk_n1351, u1_uk_n1356, u1_uk_n1360, u1_uk_n1361, u1_uk_n1366, u1_uk_n1367, u1_uk_n1372, 
       u1_uk_n1375, u1_uk_n1376, u1_uk_n1380, u1_uk_n1381, u1_uk_n1382, u1_uk_n1383, u1_uk_n1390, u1_uk_n1394, u1_uk_n1395, 
       u1_uk_n1396, u1_uk_n1400, u1_uk_n1406, u1_uk_n1407, u1_uk_n1408, u1_uk_n141, u1_uk_n1413, u1_uk_n1414, u1_uk_n1419, 
       u1_uk_n142, u1_uk_n1425, u1_uk_n1426, u1_uk_n1431, u1_uk_n145, u1_uk_n146, u1_uk_n147, u1_uk_n148, u1_uk_n1482, 
       u1_uk_n1483, u1_uk_n1484, u1_uk_n1485, u1_uk_n1486, u1_uk_n1487, u1_uk_n1488, u1_uk_n1489, u1_uk_n1490, u1_uk_n1491, 
       u1_uk_n1492, u1_uk_n1494, u1_uk_n1496, u1_uk_n1498, u1_uk_n1499, u1_uk_n1500, u1_uk_n1501, u1_uk_n1505, u1_uk_n1507, 
       u1_uk_n1510, u1_uk_n1514, u1_uk_n1516, u1_uk_n1517, u1_uk_n1518, u1_uk_n1521, u1_uk_n1523, u1_uk_n1524, u1_uk_n1526, 
       u1_uk_n1527, u1_uk_n1530, u1_uk_n1531, u1_uk_n1532, u1_uk_n1536, u1_uk_n1537, u1_uk_n1538, u1_uk_n1544, u1_uk_n1545, 
       u1_uk_n1548, u1_uk_n1549, u1_uk_n155, u1_uk_n1551, u1_uk_n1552, u1_uk_n1557, u1_uk_n1558, u1_uk_n1559, u1_uk_n1564, 
       u1_uk_n1565, u1_uk_n1570, u1_uk_n1571, u1_uk_n1588, u1_uk_n1595, u1_uk_n1606, u1_uk_n1607, u1_uk_n161, u1_uk_n1612, 
       u1_uk_n1613, u1_uk_n1615, u1_uk_n162, u1_uk_n163, u1_uk_n1664, u1_uk_n1670, u1_uk_n1672, u1_uk_n1678, u1_uk_n1694, 
       u1_uk_n17, u1_uk_n1702, u1_uk_n1711, u1_uk_n1712, u1_uk_n1716, u1_uk_n1732, u1_uk_n1738, u1_uk_n182, u1_uk_n1844, 
       u1_uk_n1845, u1_uk_n1846, u1_uk_n1847, u1_uk_n1849, u1_uk_n1850, u1_uk_n1851, u1_uk_n1852, u1_uk_n1853, u1_uk_n1855, 
       u1_uk_n1858, u1_uk_n1859, u1_uk_n1862, u1_uk_n1863, u1_uk_n1864, u1_uk_n1865, u1_uk_n1867, u1_uk_n1868, u1_uk_n1869, 
       u1_uk_n1872, u1_uk_n1873, u1_uk_n1874, u1_uk_n1876, u1_uk_n188, u1_uk_n1880, u1_uk_n1881, u1_uk_n1882, u1_uk_n1883, 
       u1_uk_n1887, u1_uk_n191, u1_uk_n202, u1_uk_n208, u1_uk_n209, u1_uk_n213, u1_uk_n214, u1_uk_n217, u1_uk_n220, 
       u1_uk_n222, u1_uk_n223, u1_uk_n230, u1_uk_n231, u1_uk_n238, u1_uk_n240, u1_uk_n242, u1_uk_n250, u1_uk_n251, 
       u1_uk_n252, u1_uk_n257, u1_uk_n27, u1_uk_n271, u1_uk_n277, u1_uk_n279, u1_uk_n292, u1_uk_n31, u1_uk_n60, 
       u1_uk_n83, u1_uk_n93, u1_uk_n99, u2_L0_14, u2_L0_25, u2_L0_3, u2_L0_8, u2_R0_16, u2_R0_17, 
       u2_R0_18, u2_R0_19, u2_R0_20, u2_R0_21, u2_uk_K_r0_15, u2_uk_K_r0_49, u2_uk_n10, u2_uk_n102, u2_uk_n110, 
       u2_uk_n1230, u2_uk_n1237, u2_uk_n1252, u2_uk_n1259, u2_uk_n1264, u2_uk_n1265, u2_uk_n161, u2_uk_n162, u2_uk_n17, 
       u2_uk_n203, u2_uk_n208, u2_uk_n27, u2_uk_n996, u2_uk_n997, u0_N328, u0_N336, u0_N342, u0_N350, u0_N36, u0_N448, u0_N457, u0_N46, u0_N467, 
        u0_N473, u0_N52, u0_N58, u0_N66, u0_N67, u0_N71, u0_N74, u0_N77, u0_N82, 
        u0_N88, u0_N92, u1_FP_11, u1_FP_12, u1_FP_14, u1_FP_15, u1_FP_19, u1_FP_21, u1_FP_22, 
        u1_FP_25, u1_FP_27, u1_FP_29, u1_FP_3, u1_FP_32, u1_FP_4, u1_FP_5, u1_FP_7, u1_FP_8, 
        u1_N102, u1_N106, u1_N107, u1_N114, u1_N117, u1_N124, u1_N127, u1_N130, u1_N132, 
        u1_N135, u1_N141, u1_N142, u1_N148, u1_N152, u1_N154, u1_N193, u1_N196, u1_N197, 
        u1_N198, u1_N203, u1_N204, u1_N206, u1_N207, u1_N209, u1_N212, u1_N213, u1_N215, 
        u1_N218, u1_N219, u1_N221, u1_N223, u1_N225, u1_N229, u1_N232, u1_N236, u1_N239, 
        u1_N240, u1_N241, u1_N246, u1_N247, u1_N251, u1_N253, u1_N254, u1_N260, u1_N270, 
        u1_N276, u1_N282, u1_N326, u1_N331, u1_N341, u1_N351, u1_N360, u1_N368, u1_N374, 
        u1_N382, u1_N40, u1_N448, u1_N449, u1_N450, u1_N453, u1_N455, u1_N456, u1_N457, 
        u1_N460, u1_N461, u1_N463, u1_N464, u1_N465, u1_N467, u1_N470, u1_N471, u1_N472, 
        u1_N473, u1_N475, u1_N477, u1_N478, u1_N48, u1_N54, u1_N62, u1_N99, u1_uk_n100, 
        u1_uk_n110, u1_uk_n164, u1_uk_n187, u1_uk_n203, u1_uk_n207, u1_uk_n291, u1_uk_n294, u1_uk_n297, u1_uk_n298, 
        u1_uk_n63, u1_uk_n92, u1_uk_n94, u2_N34, u2_N39, u2_N45, u2_N56 );
  input n116, u0_K2_44, u0_K2_45, u0_K2_46, u0_K2_47, u0_K2_48, u0_K3_34, u0_L0_15, u0_L0_21, 
        u0_L0_27, u0_L0_5, u0_L13_1, u0_L13_10, u0_L13_20, u0_L13_26, u0_L1_11, u0_L1_14, u0_L1_19, 
        u0_L1_25, u0_L1_29, u0_L1_3, u0_L1_4, u0_L1_8, u0_L9_17, u0_L9_23, u0_L9_31, u0_L9_9, 
        u0_R0_1, u0_R0_28, u0_R0_29, u0_R0_30, u0_R0_31, u0_R0_32, u0_R13_12, u0_R13_13, u0_R13_14, 
        u0_R13_15, u0_R13_16, u0_R13_17, u0_R1_16, u0_R1_17, u0_R1_18, u0_R1_19, u0_R1_20, u0_R1_21, 
        u0_R1_22, u0_R1_23, u0_R1_24, u0_R1_25, u0_R9_1, u0_R9_2, u0_R9_3, u0_R9_32, u0_R9_4, 
        u0_R9_5, u0_uk_K_r0_2, u0_uk_K_r1_42, u0_uk_K_r1_44, u0_uk_K_r1_7, u0_uk_K_r9_19, u0_uk_K_r9_25, u0_uk_n109, u0_uk_n11, 
        u0_uk_n118, u0_uk_n129, u0_uk_n14, u0_uk_n141, u0_uk_n142, u0_uk_n148, u0_uk_n16, u0_uk_n163, u0_uk_n164, 
        u0_uk_n181, u0_uk_n183, u0_uk_n187, u0_uk_n188, u0_uk_n189, u0_uk_n191, u0_uk_n195, u0_uk_n200, u0_uk_n201, 
        u0_uk_n202, u0_uk_n209, u0_uk_n215, u0_uk_n219, u0_uk_n220, u0_uk_n222, u0_uk_n231, u0_uk_n238, u0_uk_n24, 
        u0_uk_n242, u0_uk_n25, u0_uk_n252, u0_uk_n30, u0_uk_n37, u0_uk_n38, u0_uk_n42, u0_uk_n43, u0_uk_n543, 
        u0_uk_n544, u0_uk_n545, u0_uk_n549, u0_uk_n555, u0_uk_n559, u0_uk_n560, u0_uk_n566, u0_uk_n570, u0_uk_n575, 
        u0_uk_n579, u0_uk_n580, u0_uk_n60, u0_uk_n612, u0_uk_n63, u0_uk_n7, u0_uk_n83, u0_uk_n92, u0_uk_n93, 
        u0_uk_n94, u1_FP_33, u1_FP_48, u1_FP_49, u1_FP_50, u1_FP_51, u1_FP_52, u1_FP_53, u1_FP_54, 
        u1_FP_55, u1_FP_56, u1_FP_57, u1_FP_58, u1_FP_59, u1_FP_60, u1_FP_61, u1_FP_62, u1_FP_63, 
        u1_FP_64, u1_L0_17, u1_L0_23, u1_L0_31, u1_L0_9, u1_L10_17, u1_L10_23, u1_L10_31, u1_L10_9, 
        u1_L13_1, u1_L13_10, u1_L13_13, u1_L13_14, u1_L13_16, u1_L13_17, u1_L13_18, u1_L13_2, u1_L13_20, 
        u1_L13_23, u1_L13_24, u1_L13_25, u1_L13_26, u1_L13_28, u1_L13_3, u1_L13_30, u1_L13_31, u1_L13_6, 
        u1_L13_8, u1_L13_9, u1_L14_11, u1_L14_12, u1_L14_14, u1_L14_15, u1_L14_19, u1_L14_21, u1_L14_22, 
        u1_L14_25, u1_L14_27, u1_L14_29, u1_L14_3, u1_L14_32, u1_L14_4, u1_L14_5, u1_L14_7, u1_L14_8, 
        u1_L2_11, u1_L2_12, u1_L2_19, u1_L2_22, u1_L2_29, u1_L2_32, u1_L2_4, u1_L2_7, u1_L3_14, 
        u1_L3_15, u1_L3_21, u1_L3_25, u1_L3_27, u1_L3_3, u1_L3_5, u1_L3_8, u1_L5_12, u1_L5_13, 
        u1_L5_15, u1_L5_16, u1_L5_18, u1_L5_2, u1_L5_21, u1_L5_22, u1_L5_24, u1_L5_27, u1_L5_28, 
        u1_L5_30, u1_L5_32, u1_L5_5, u1_L5_6, u1_L5_7, u1_L6_13, u1_L6_16, u1_L6_17, u1_L6_18, 
        u1_L6_2, u1_L6_23, u1_L6_24, u1_L6_28, u1_L6_30, u1_L6_31, u1_L6_6, u1_L6_9, u1_L7_15, 
        u1_L7_21, u1_L7_27, u1_L7_5, u1_L9_12, u1_L9_22, u1_L9_32, u1_L9_7, u1_R0_1, u1_R0_2, 
        u1_R0_3, u1_R0_32, u1_R0_4, u1_R0_5, u1_R10_1, u1_R10_2, u1_R10_3, u1_R10_32, u1_R10_4, 
        u1_R10_5, u1_R13_1, u1_R13_10, u1_R13_11, u1_R13_12, u1_R13_13, u1_R13_14, u1_R13_15, u1_R13_16, 
        u1_R13_17, u1_R13_18, u1_R13_19, u1_R13_2, u1_R13_20, u1_R13_21, u1_R13_3, u1_R13_32, u1_R13_4, 
        u1_R13_5, u1_R13_6, u1_R13_7, u1_R13_8, u1_R13_9, u1_R2_20, u1_R2_21, u1_R2_22, u1_R2_23, 
        u1_R2_24, u1_R2_25, u1_R2_26, u1_R2_27, u1_R2_28, u1_R2_29, u1_R3_1, u1_R3_16, u1_R3_17, 
        u1_R3_18, u1_R3_19, u1_R3_20, u1_R3_21, u1_R3_28, u1_R3_29, u1_R3_30, u1_R3_31, u1_R3_32, 
        u1_R5_1, u1_R5_10, u1_R5_11, u1_R5_12, u1_R5_13, u1_R5_24, u1_R5_25, u1_R5_26, u1_R5_27, 
        u1_R5_28, u1_R5_29, u1_R5_30, u1_R5_31, u1_R5_32, u1_R5_4, u1_R5_5, u1_R5_6, u1_R5_7, 
        u1_R5_8, u1_R5_9, u1_R6_1, u1_R6_10, u1_R6_11, u1_R6_12, u1_R6_13, u1_R6_2, u1_R6_3, 
        u1_R6_32, u1_R6_4, u1_R6_5, u1_R6_6, u1_R6_7, u1_R6_8, u1_R6_9, u1_R7_1, u1_R7_28, 
        u1_R7_29, u1_R7_30, u1_R7_31, u1_R7_32, u1_R9_24, u1_R9_25, u1_R9_26, u1_R9_27, u1_R9_28, 
        u1_R9_29, u1_uk_K_r10_10, u1_uk_K_r10_18, u1_uk_K_r10_27, u1_uk_K_r10_39, u1_uk_K_r10_4, u1_uk_K_r10_48, u1_uk_K_r13_0, u1_uk_K_r13_13, 
        u1_uk_K_r13_17, u1_uk_K_r13_19, u1_uk_K_r13_22, u1_uk_K_r13_25, u1_uk_K_r13_32, u1_uk_K_r13_38, u1_uk_K_r13_4, u1_uk_K_r13_44, u1_uk_K_r13_55, 
        u1_uk_K_r14_15, u1_uk_K_r14_16, u1_uk_K_r14_2, u1_uk_K_r14_23, u1_uk_K_r14_38, u1_uk_K_r14_42, u1_uk_K_r14_43, u1_uk_K_r14_45, u1_uk_K_r14_50, 
        u1_uk_K_r14_8, u1_uk_K_r14_9, u1_uk_K_r2_31, u1_uk_K_r2_49, u1_uk_K_r2_50, u1_uk_K_r3_15, u1_uk_K_r3_35, u1_uk_K_r3_38, u1_uk_K_r3_43, 
        u1_uk_K_r3_51, u1_uk_K_r5_1, u1_uk_K_r5_17, u1_uk_K_r5_23, u1_uk_K_r5_26, u1_uk_K_r5_31, u1_uk_K_r5_32, u1_uk_K_r5_36, u1_uk_K_r5_39, 
        u1_uk_K_r5_4, u1_uk_K_r5_48, u1_uk_K_r5_8, u1_uk_K_r6_10, u1_uk_K_r6_17, u1_uk_K_r6_19, u1_uk_K_r6_26, u1_uk_K_r6_27, u1_uk_K_r6_3, 
        u1_uk_K_r6_34, u1_uk_K_r6_46, u1_uk_K_r6_53, u1_uk_K_r6_55, u1_uk_K_r7_0, u1_uk_K_r7_16, u1_uk_K_r7_37, u1_uk_K_r7_9, u1_uk_K_r9_30, 
        u1_uk_K_r9_31, u1_uk_K_r9_38, u1_uk_K_r9_7, u1_uk_n102, u1_uk_n109, u1_uk_n11, u1_uk_n117, u1_uk_n118, u1_uk_n1218, 
        u1_uk_n1219, u1_uk_n1222, u1_uk_n1225, u1_uk_n1230, u1_uk_n1231, u1_uk_n1233, u1_uk_n1238, u1_uk_n1239, u1_uk_n1240, 
        u1_uk_n1241, u1_uk_n1245, u1_uk_n1246, u1_uk_n1247, u1_uk_n1250, u1_uk_n1253, u1_uk_n1255, u1_uk_n1256, u1_uk_n1268, 
        u1_uk_n1269, u1_uk_n1273, u1_uk_n1274, u1_uk_n1277, u1_uk_n1279, u1_uk_n1284, u1_uk_n129, u1_uk_n1297, u1_uk_n1300, 
        u1_uk_n1305, u1_uk_n1349, u1_uk_n1351, u1_uk_n1356, u1_uk_n1360, u1_uk_n1361, u1_uk_n1366, u1_uk_n1367, u1_uk_n1372, 
        u1_uk_n1375, u1_uk_n1376, u1_uk_n1380, u1_uk_n1381, u1_uk_n1382, u1_uk_n1383, u1_uk_n1390, u1_uk_n1394, u1_uk_n1395, 
        u1_uk_n1396, u1_uk_n1400, u1_uk_n1406, u1_uk_n1407, u1_uk_n1408, u1_uk_n141, u1_uk_n1413, u1_uk_n1414, u1_uk_n1419, 
        u1_uk_n142, u1_uk_n1425, u1_uk_n1426, u1_uk_n1431, u1_uk_n145, u1_uk_n146, u1_uk_n147, u1_uk_n148, u1_uk_n1482, 
        u1_uk_n1483, u1_uk_n1484, u1_uk_n1485, u1_uk_n1486, u1_uk_n1487, u1_uk_n1488, u1_uk_n1489, u1_uk_n1490, u1_uk_n1491, 
        u1_uk_n1492, u1_uk_n1494, u1_uk_n1496, u1_uk_n1498, u1_uk_n1499, u1_uk_n1500, u1_uk_n1501, u1_uk_n1505, u1_uk_n1507, 
        u1_uk_n1510, u1_uk_n1514, u1_uk_n1516, u1_uk_n1517, u1_uk_n1518, u1_uk_n1521, u1_uk_n1523, u1_uk_n1524, u1_uk_n1526, 
        u1_uk_n1527, u1_uk_n1530, u1_uk_n1531, u1_uk_n1532, u1_uk_n1536, u1_uk_n1537, u1_uk_n1538, u1_uk_n1544, u1_uk_n1545, 
        u1_uk_n1548, u1_uk_n1549, u1_uk_n155, u1_uk_n1551, u1_uk_n1552, u1_uk_n1557, u1_uk_n1558, u1_uk_n1559, u1_uk_n1564, 
        u1_uk_n1565, u1_uk_n1570, u1_uk_n1571, u1_uk_n1588, u1_uk_n1595, u1_uk_n1606, u1_uk_n1607, u1_uk_n161, u1_uk_n1612, 
        u1_uk_n1613, u1_uk_n1615, u1_uk_n162, u1_uk_n163, u1_uk_n1664, u1_uk_n1670, u1_uk_n1672, u1_uk_n1678, u1_uk_n1694, 
        u1_uk_n17, u1_uk_n1702, u1_uk_n1711, u1_uk_n1712, u1_uk_n1716, u1_uk_n1732, u1_uk_n1738, u1_uk_n182, u1_uk_n1844, 
        u1_uk_n1845, u1_uk_n1846, u1_uk_n1847, u1_uk_n1849, u1_uk_n1850, u1_uk_n1851, u1_uk_n1852, u1_uk_n1853, u1_uk_n1855, 
        u1_uk_n1858, u1_uk_n1859, u1_uk_n1862, u1_uk_n1863, u1_uk_n1864, u1_uk_n1865, u1_uk_n1867, u1_uk_n1868, u1_uk_n1869, 
        u1_uk_n1872, u1_uk_n1873, u1_uk_n1874, u1_uk_n1876, u1_uk_n188, u1_uk_n1880, u1_uk_n1881, u1_uk_n1882, u1_uk_n1883, 
        u1_uk_n1887, u1_uk_n191, u1_uk_n202, u1_uk_n208, u1_uk_n209, u1_uk_n213, u1_uk_n214, u1_uk_n217, u1_uk_n220, 
        u1_uk_n222, u1_uk_n223, u1_uk_n230, u1_uk_n231, u1_uk_n238, u1_uk_n240, u1_uk_n242, u1_uk_n250, u1_uk_n251, 
        u1_uk_n252, u1_uk_n257, u1_uk_n27, u1_uk_n271, u1_uk_n277, u1_uk_n279, u1_uk_n292, u1_uk_n31, u1_uk_n60, 
        u1_uk_n83, u1_uk_n93, u1_uk_n99, u2_L0_14, u2_L0_25, u2_L0_3, u2_L0_8, u2_R0_16, u2_R0_17, 
        u2_R0_18, u2_R0_19, u2_R0_20, u2_R0_21, u2_uk_K_r0_15, u2_uk_K_r0_49, u2_uk_n10, u2_uk_n102, u2_uk_n110, 
        u2_uk_n1230, u2_uk_n1237, u2_uk_n1252, u2_uk_n1259, u2_uk_n1264, u2_uk_n1265, u2_uk_n161, u2_uk_n162, u2_uk_n17, 
        u2_uk_n203, u2_uk_n208, u2_uk_n27, u2_uk_n996, u2_uk_n997;
  output u0_N328, u0_N336, u0_N342, u0_N350, u0_N36, u0_N448, u0_N457, u0_N46, u0_N467, 
        u0_N473, u0_N52, u0_N58, u0_N66, u0_N67, u0_N71, u0_N74, u0_N77, u0_N82, 
        u0_N88, u0_N92, u1_FP_11, u1_FP_12, u1_FP_14, u1_FP_15, u1_FP_19, u1_FP_21, u1_FP_22, 
        u1_FP_25, u1_FP_27, u1_FP_29, u1_FP_3, u1_FP_32, u1_FP_4, u1_FP_5, u1_FP_7, u1_FP_8, 
        u1_N102, u1_N106, u1_N107, u1_N114, u1_N117, u1_N124, u1_N127, u1_N130, u1_N132, 
        u1_N135, u1_N141, u1_N142, u1_N148, u1_N152, u1_N154, u1_N193, u1_N196, u1_N197, 
        u1_N198, u1_N203, u1_N204, u1_N206, u1_N207, u1_N209, u1_N212, u1_N213, u1_N215, 
        u1_N218, u1_N219, u1_N221, u1_N223, u1_N225, u1_N229, u1_N232, u1_N236, u1_N239, 
        u1_N240, u1_N241, u1_N246, u1_N247, u1_N251, u1_N253, u1_N254, u1_N260, u1_N270, 
        u1_N276, u1_N282, u1_N326, u1_N331, u1_N341, u1_N351, u1_N360, u1_N368, u1_N374, 
        u1_N382, u1_N40, u1_N448, u1_N449, u1_N450, u1_N453, u1_N455, u1_N456, u1_N457, 
        u1_N460, u1_N461, u1_N463, u1_N464, u1_N465, u1_N467, u1_N470, u1_N471, u1_N472, 
        u1_N473, u1_N475, u1_N477, u1_N478, u1_N48, u1_N54, u1_N62, u1_N99, u1_uk_n100, 
        u1_uk_n110, u1_uk_n164, u1_uk_n187, u1_uk_n203, u1_uk_n207, u1_uk_n291, u1_uk_n294, u1_uk_n297, u1_uk_n298, 
        u1_uk_n63, u1_uk_n92, u1_uk_n94, u2_N34, u2_N39, u2_N45, u2_N56;
  wire u0_K11_1, u0_K11_2, u0_K11_3, u0_K11_4, u0_K11_5, u0_K11_6, u0_K15_19, u0_K15_20, u0_K15_21, 
       u0_K15_22, u0_K15_23, u0_K15_24, u0_K2_43, u0_K3_25, u0_K3_26, u0_K3_27, u0_K3_28, u0_K3_29, 
       u0_K3_30, u0_K3_31, u0_K3_32, u0_K3_33, u0_K3_35, u0_K3_36, u0_out10_17, u0_out10_23, u0_out10_31, 
       u0_out10_9, u0_out14_1, u0_out14_10, u0_out14_20, u0_out14_26, u0_out1_15, u0_out1_21, u0_out1_27, u0_out1_5, 
       u0_out2_11, u0_out2_14, u0_out2_19, u0_out2_25, u0_out2_29, u0_out2_3, u0_out2_4, u0_out2_8, u0_u10_X_1, 
       u0_u10_X_2, u0_u10_X_3, u0_u10_X_4, u0_u10_X_5, u0_u10_X_6, u0_u10_u0_n100, u0_u10_u0_n101, u0_u10_u0_n102, u0_u10_u0_n103, 
       u0_u10_u0_n104, u0_u10_u0_n105, u0_u10_u0_n106, u0_u10_u0_n107, u0_u10_u0_n108, u0_u10_u0_n109, u0_u10_u0_n110, u0_u10_u0_n111, u0_u10_u0_n112, 
       u0_u10_u0_n113, u0_u10_u0_n114, u0_u10_u0_n115, u0_u10_u0_n116, u0_u10_u0_n117, u0_u10_u0_n118, u0_u10_u0_n119, u0_u10_u0_n120, u0_u10_u0_n121, 
       u0_u10_u0_n122, u0_u10_u0_n123, u0_u10_u0_n124, u0_u10_u0_n125, u0_u10_u0_n126, u0_u10_u0_n127, u0_u10_u0_n128, u0_u10_u0_n129, u0_u10_u0_n130, 
       u0_u10_u0_n131, u0_u10_u0_n132, u0_u10_u0_n133, u0_u10_u0_n134, u0_u10_u0_n135, u0_u10_u0_n136, u0_u10_u0_n137, u0_u10_u0_n138, u0_u10_u0_n139, 
       u0_u10_u0_n140, u0_u10_u0_n141, u0_u10_u0_n142, u0_u10_u0_n143, u0_u10_u0_n144, u0_u10_u0_n145, u0_u10_u0_n146, u0_u10_u0_n147, u0_u10_u0_n148, 
       u0_u10_u0_n149, u0_u10_u0_n150, u0_u10_u0_n151, u0_u10_u0_n152, u0_u10_u0_n153, u0_u10_u0_n154, u0_u10_u0_n155, u0_u10_u0_n156, u0_u10_u0_n157, 
       u0_u10_u0_n158, u0_u10_u0_n159, u0_u10_u0_n160, u0_u10_u0_n161, u0_u10_u0_n162, u0_u10_u0_n163, u0_u10_u0_n164, u0_u10_u0_n165, u0_u10_u0_n166, 
       u0_u10_u0_n167, u0_u10_u0_n168, u0_u10_u0_n169, u0_u10_u0_n170, u0_u10_u0_n171, u0_u10_u0_n172, u0_u10_u0_n173, u0_u10_u0_n174, u0_u10_u0_n88, 
       u0_u10_u0_n89, u0_u10_u0_n90, u0_u10_u0_n91, u0_u10_u0_n92, u0_u10_u0_n93, u0_u10_u0_n94, u0_u10_u0_n95, u0_u10_u0_n96, u0_u10_u0_n97, 
       u0_u10_u0_n98, u0_u10_u0_n99, u0_u14_X_19, u0_u14_X_20, u0_u14_X_21, u0_u14_X_22, u0_u14_X_23, u0_u14_X_24, u0_u14_u3_n100, 
       u0_u14_u3_n101, u0_u14_u3_n102, u0_u14_u3_n103, u0_u14_u3_n104, u0_u14_u3_n105, u0_u14_u3_n106, u0_u14_u3_n107, u0_u14_u3_n108, u0_u14_u3_n109, 
       u0_u14_u3_n110, u0_u14_u3_n111, u0_u14_u3_n112, u0_u14_u3_n113, u0_u14_u3_n114, u0_u14_u3_n115, u0_u14_u3_n116, u0_u14_u3_n117, u0_u14_u3_n118, 
       u0_u14_u3_n119, u0_u14_u3_n120, u0_u14_u3_n121, u0_u14_u3_n122, u0_u14_u3_n123, u0_u14_u3_n124, u0_u14_u3_n125, u0_u14_u3_n126, u0_u14_u3_n127, 
       u0_u14_u3_n128, u0_u14_u3_n129, u0_u14_u3_n130, u0_u14_u3_n131, u0_u14_u3_n132, u0_u14_u3_n133, u0_u14_u3_n134, u0_u14_u3_n135, u0_u14_u3_n136, 
       u0_u14_u3_n137, u0_u14_u3_n138, u0_u14_u3_n139, u0_u14_u3_n140, u0_u14_u3_n141, u0_u14_u3_n142, u0_u14_u3_n143, u0_u14_u3_n144, u0_u14_u3_n145, 
       u0_u14_u3_n146, u0_u14_u3_n147, u0_u14_u3_n148, u0_u14_u3_n149, u0_u14_u3_n150, u0_u14_u3_n151, u0_u14_u3_n152, u0_u14_u3_n153, u0_u14_u3_n154, 
       u0_u14_u3_n155, u0_u14_u3_n156, u0_u14_u3_n157, u0_u14_u3_n158, u0_u14_u3_n159, u0_u14_u3_n160, u0_u14_u3_n161, u0_u14_u3_n162, u0_u14_u3_n163, 
       u0_u14_u3_n164, u0_u14_u3_n165, u0_u14_u3_n166, u0_u14_u3_n167, u0_u14_u3_n168, u0_u14_u3_n169, u0_u14_u3_n170, u0_u14_u3_n171, u0_u14_u3_n172, 
       u0_u14_u3_n173, u0_u14_u3_n174, u0_u14_u3_n175, u0_u14_u3_n176, u0_u14_u3_n177, u0_u14_u3_n178, u0_u14_u3_n179, u0_u14_u3_n180, u0_u14_u3_n181, 
       u0_u14_u3_n182, u0_u14_u3_n183, u0_u14_u3_n184, u0_u14_u3_n185, u0_u14_u3_n186, u0_u14_u3_n94, u0_u14_u3_n95, u0_u14_u3_n96, u0_u14_u3_n97, 
       u0_u14_u3_n98, u0_u14_u3_n99, u0_u1_X_43, u0_u1_X_44, u0_u1_X_45, u0_u1_X_46, u0_u1_X_47, u0_u1_X_48, u0_u1_u7_n100, 
       u0_u1_u7_n101, u0_u1_u7_n102, u0_u1_u7_n103, u0_u1_u7_n104, u0_u1_u7_n105, u0_u1_u7_n106, u0_u1_u7_n107, u0_u1_u7_n108, u0_u1_u7_n109, 
       u0_u1_u7_n110, u0_u1_u7_n111, u0_u1_u7_n112, u0_u1_u7_n113, u0_u1_u7_n114, u0_u1_u7_n115, u0_u1_u7_n116, u0_u1_u7_n117, u0_u1_u7_n118, 
       u0_u1_u7_n119, u0_u1_u7_n120, u0_u1_u7_n121, u0_u1_u7_n122, u0_u1_u7_n123, u0_u1_u7_n124, u0_u1_u7_n125, u0_u1_u7_n126, u0_u1_u7_n127, 
       u0_u1_u7_n128, u0_u1_u7_n129, u0_u1_u7_n130, u0_u1_u7_n131, u0_u1_u7_n132, u0_u1_u7_n133, u0_u1_u7_n134, u0_u1_u7_n135, u0_u1_u7_n136, 
       u0_u1_u7_n137, u0_u1_u7_n138, u0_u1_u7_n139, u0_u1_u7_n140, u0_u1_u7_n141, u0_u1_u7_n142, u0_u1_u7_n143, u0_u1_u7_n144, u0_u1_u7_n145, 
       u0_u1_u7_n146, u0_u1_u7_n147, u0_u1_u7_n148, u0_u1_u7_n149, u0_u1_u7_n150, u0_u1_u7_n151, u0_u1_u7_n152, u0_u1_u7_n153, u0_u1_u7_n154, 
       u0_u1_u7_n155, u0_u1_u7_n156, u0_u1_u7_n157, u0_u1_u7_n158, u0_u1_u7_n159, u0_u1_u7_n160, u0_u1_u7_n161, u0_u1_u7_n162, u0_u1_u7_n163, 
       u0_u1_u7_n164, u0_u1_u7_n165, u0_u1_u7_n166, u0_u1_u7_n167, u0_u1_u7_n168, u0_u1_u7_n169, u0_u1_u7_n170, u0_u1_u7_n171, u0_u1_u7_n172, 
       u0_u1_u7_n173, u0_u1_u7_n174, u0_u1_u7_n175, u0_u1_u7_n176, u0_u1_u7_n177, u0_u1_u7_n178, u0_u1_u7_n179, u0_u1_u7_n180, u0_u1_u7_n91, 
       u0_u1_u7_n92, u0_u1_u7_n93, u0_u1_u7_n94, u0_u1_u7_n95, u0_u1_u7_n96, u0_u1_u7_n97, u0_u1_u7_n98, u0_u1_u7_n99, u0_u2_X_25, 
       u0_u2_X_26, u0_u2_X_27, u0_u2_X_28, u0_u2_X_29, u0_u2_X_30, u0_u2_X_31, u0_u2_X_32, u0_u2_X_33, u0_u2_X_34, 
       u0_u2_X_35, u0_u2_X_36, u0_u2_u4_n100, u0_u2_u4_n101, u0_u2_u4_n102, u0_u2_u4_n103, u0_u2_u4_n104, u0_u2_u4_n105, u0_u2_u4_n106, 
       u0_u2_u4_n107, u0_u2_u4_n108, u0_u2_u4_n109, u0_u2_u4_n110, u0_u2_u4_n111, u0_u2_u4_n112, u0_u2_u4_n113, u0_u2_u4_n114, u0_u2_u4_n115, 
       u0_u2_u4_n116, u0_u2_u4_n117, u0_u2_u4_n118, u0_u2_u4_n119, u0_u2_u4_n120, u0_u2_u4_n121, u0_u2_u4_n122, u0_u2_u4_n123, u0_u2_u4_n124, 
       u0_u2_u4_n125, u0_u2_u4_n126, u0_u2_u4_n127, u0_u2_u4_n128, u0_u2_u4_n129, u0_u2_u4_n130, u0_u2_u4_n131, u0_u2_u4_n132, u0_u2_u4_n133, 
       u0_u2_u4_n134, u0_u2_u4_n135, u0_u2_u4_n136, u0_u2_u4_n137, u0_u2_u4_n138, u0_u2_u4_n139, u0_u2_u4_n140, u0_u2_u4_n141, u0_u2_u4_n142, 
       u0_u2_u4_n143, u0_u2_u4_n144, u0_u2_u4_n145, u0_u2_u4_n146, u0_u2_u4_n147, u0_u2_u4_n148, u0_u2_u4_n149, u0_u2_u4_n150, u0_u2_u4_n151, 
       u0_u2_u4_n152, u0_u2_u4_n153, u0_u2_u4_n154, u0_u2_u4_n155, u0_u2_u4_n156, u0_u2_u4_n157, u0_u2_u4_n158, u0_u2_u4_n159, u0_u2_u4_n160, 
       u0_u2_u4_n161, u0_u2_u4_n162, u0_u2_u4_n163, u0_u2_u4_n164, u0_u2_u4_n165, u0_u2_u4_n166, u0_u2_u4_n167, u0_u2_u4_n168, u0_u2_u4_n169, 
       u0_u2_u4_n170, u0_u2_u4_n171, u0_u2_u4_n172, u0_u2_u4_n173, u0_u2_u4_n174, u0_u2_u4_n175, u0_u2_u4_n176, u0_u2_u4_n177, u0_u2_u4_n178, 
       u0_u2_u4_n179, u0_u2_u4_n180, u0_u2_u4_n181, u0_u2_u4_n182, u0_u2_u4_n183, u0_u2_u4_n184, u0_u2_u4_n185, u0_u2_u4_n186, u0_u2_u4_n94, 
       u0_u2_u4_n95, u0_u2_u4_n96, u0_u2_u4_n97, u0_u2_u4_n98, u0_u2_u4_n99, u0_u2_u5_n100, u0_u2_u5_n101, u0_u2_u5_n102, u0_u2_u5_n103, 
       u0_u2_u5_n104, u0_u2_u5_n105, u0_u2_u5_n106, u0_u2_u5_n107, u0_u2_u5_n108, u0_u2_u5_n109, u0_u2_u5_n110, u0_u2_u5_n111, u0_u2_u5_n112, 
       u0_u2_u5_n113, u0_u2_u5_n114, u0_u2_u5_n115, u0_u2_u5_n116, u0_u2_u5_n117, u0_u2_u5_n118, u0_u2_u5_n119, u0_u2_u5_n120, u0_u2_u5_n121, 
       u0_u2_u5_n122, u0_u2_u5_n123, u0_u2_u5_n124, u0_u2_u5_n125, u0_u2_u5_n126, u0_u2_u5_n127, u0_u2_u5_n128, u0_u2_u5_n129, u0_u2_u5_n130, 
       u0_u2_u5_n131, u0_u2_u5_n132, u0_u2_u5_n133, u0_u2_u5_n134, u0_u2_u5_n135, u0_u2_u5_n136, u0_u2_u5_n137, u0_u2_u5_n138, u0_u2_u5_n139, 
       u0_u2_u5_n140, u0_u2_u5_n141, u0_u2_u5_n142, u0_u2_u5_n143, u0_u2_u5_n144, u0_u2_u5_n145, u0_u2_u5_n146, u0_u2_u5_n147, u0_u2_u5_n148, 
       u0_u2_u5_n149, u0_u2_u5_n150, u0_u2_u5_n151, u0_u2_u5_n152, u0_u2_u5_n153, u0_u2_u5_n154, u0_u2_u5_n155, u0_u2_u5_n156, u0_u2_u5_n157, 
       u0_u2_u5_n158, u0_u2_u5_n159, u0_u2_u5_n160, u0_u2_u5_n161, u0_u2_u5_n162, u0_u2_u5_n163, u0_u2_u5_n164, u0_u2_u5_n165, u0_u2_u5_n166, 
       u0_u2_u5_n167, u0_u2_u5_n168, u0_u2_u5_n169, u0_u2_u5_n170, u0_u2_u5_n171, u0_u2_u5_n172, u0_u2_u5_n173, u0_u2_u5_n174, u0_u2_u5_n175, 
       u0_u2_u5_n176, u0_u2_u5_n177, u0_u2_u5_n178, u0_u2_u5_n179, u0_u2_u5_n180, u0_u2_u5_n181, u0_u2_u5_n182, u0_u2_u5_n183, u0_u2_u5_n184, 
       u0_u2_u5_n185, u0_u2_u5_n186, u0_u2_u5_n187, u0_u2_u5_n188, u0_u2_u5_n189, u0_u2_u5_n190, u0_u2_u5_n191, u0_u2_u5_n192, u0_u2_u5_n193, 
       u0_u2_u5_n194, u0_u2_u5_n195, u0_u2_u5_n196, u0_u2_u5_n99, u0_uk_n847, u0_uk_n849, u0_uk_n850, u0_uk_n857, u0_uk_n984, 
       u1_K11_37, u1_K11_38, u1_K11_39, u1_K11_40, u1_K11_41, u1_K11_42, u1_K12_1, u1_K12_2, u1_K12_3, 
       u1_K12_4, u1_K12_5, u1_K12_6, u1_K15_1, u1_K15_10, u1_K15_11, u1_K15_12, u1_K15_13, u1_K15_14, 
       u1_K15_15, u1_K15_16, u1_K15_17, u1_K15_18, u1_K15_19, u1_K15_2, u1_K15_20, u1_K15_21, u1_K15_22, 
       u1_K15_23, u1_K15_24, u1_K15_25, u1_K15_26, u1_K15_27, u1_K15_28, u1_K15_29, u1_K15_3, u1_K15_30, 
       u1_K15_4, u1_K15_5, u1_K15_6, u1_K15_7, u1_K15_8, u1_K15_9, u1_K16_25, u1_K16_26, u1_K16_27, 
       u1_K16_28, u1_K16_29, u1_K16_30, u1_K16_31, u1_K16_32, u1_K16_33, u1_K16_34, u1_K16_35, u1_K16_36, 
       u1_K16_37, u1_K16_38, u1_K16_39, u1_K16_40, u1_K16_41, u1_K16_42, u1_K16_43, u1_K16_44, u1_K16_45, 
       u1_K16_46, u1_K16_47, u1_K16_48, u1_K2_1, u1_K2_2, u1_K2_3, u1_K2_4, u1_K2_5, u1_K2_6, 
       u1_K4_31, u1_K4_32, u1_K4_33, u1_K4_34, u1_K4_35, u1_K4_36, u1_K4_37, u1_K4_38, u1_K4_39, 
       u1_K4_40, u1_K4_41, u1_K4_42, u1_K5_25, u1_K5_26, u1_K5_27, u1_K5_28, u1_K5_29, u1_K5_30, 
       u1_K5_43, u1_K5_44, u1_K5_45, u1_K5_46, u1_K5_47, u1_K5_48, u1_K7_10, u1_K7_11, u1_K7_12, 
       u1_K7_13, u1_K7_14, u1_K7_15, u1_K7_16, u1_K7_17, u1_K7_18, u1_K7_37, u1_K7_38, u1_K7_39, 
       u1_K7_40, u1_K7_41, u1_K7_42, u1_K7_43, u1_K7_44, u1_K7_45, u1_K7_46, u1_K7_47, u1_K7_48, 
       u1_K7_7, u1_K7_8, u1_K7_9, u1_K8_1, u1_K8_10, u1_K8_11, u1_K8_12, u1_K8_13, u1_K8_14, 
       u1_K8_15, u1_K8_16, u1_K8_17, u1_K8_18, u1_K8_2, u1_K8_3, u1_K8_4, u1_K8_5, u1_K8_6, 
       u1_K8_7, u1_K8_8, u1_K8_9, u1_K9_43, u1_K9_44, u1_K9_45, u1_K9_46, u1_K9_47, u1_K9_48, 
       u1_out10_12, u1_out10_22, u1_out10_32, u1_out10_7, u1_out11_17, u1_out11_23, u1_out11_31, u1_out11_9, u1_out14_1, 
       u1_out14_10, u1_out14_13, u1_out14_14, u1_out14_16, u1_out14_17, u1_out14_18, u1_out14_2, u1_out14_20, u1_out14_23, 
       u1_out14_24, u1_out14_25, u1_out14_26, u1_out14_28, u1_out14_3, u1_out14_30, u1_out14_31, u1_out14_6, u1_out14_8, 
       u1_out14_9, u1_out15_11, u1_out15_12, u1_out15_14, u1_out15_15, u1_out15_19, u1_out15_21, u1_out15_22, u1_out15_25, 
       u1_out15_27, u1_out15_29, u1_out15_3, u1_out15_32, u1_out15_4, u1_out15_5, u1_out15_7, u1_out15_8, u1_out1_17, 
       u1_out1_23, u1_out1_31, u1_out1_9, u1_out3_11, u1_out3_12, u1_out3_19, u1_out3_22, u1_out3_29, u1_out3_32, 
       u1_out3_4, u1_out3_7, u1_out4_14, u1_out4_15, u1_out4_21, u1_out4_25, u1_out4_27, u1_out4_3, u1_out4_5, 
       u1_out4_8, u1_out6_12, u1_out6_13, u1_out6_15, u1_out6_16, u1_out6_18, u1_out6_2, u1_out6_21, u1_out6_22, 
       u1_out6_24, u1_out6_27, u1_out6_28, u1_out6_30, u1_out6_32, u1_out6_5, u1_out6_6, u1_out6_7, u1_out7_13, 
       u1_out7_16, u1_out7_17, u1_out7_18, u1_out7_2, u1_out7_23, u1_out7_24, u1_out7_28, u1_out7_30, u1_out7_31, 
       u1_out7_6, u1_out7_9, u1_out8_15, u1_out8_21, u1_out8_27, u1_out8_5, u1_u10_X_37, u1_u10_X_38, u1_u10_X_39, 
       u1_u10_X_40, u1_u10_X_41, u1_u10_X_42, u1_u10_u6_n100, u1_u10_u6_n101, u1_u10_u6_n102, u1_u10_u6_n103, u1_u10_u6_n104, u1_u10_u6_n105, 
       u1_u10_u6_n106, u1_u10_u6_n107, u1_u10_u6_n108, u1_u10_u6_n109, u1_u10_u6_n110, u1_u10_u6_n111, u1_u10_u6_n112, u1_u10_u6_n113, u1_u10_u6_n114, 
       u1_u10_u6_n115, u1_u10_u6_n116, u1_u10_u6_n117, u1_u10_u6_n118, u1_u10_u6_n119, u1_u10_u6_n120, u1_u10_u6_n121, u1_u10_u6_n122, u1_u10_u6_n123, 
       u1_u10_u6_n124, u1_u10_u6_n125, u1_u10_u6_n126, u1_u10_u6_n127, u1_u10_u6_n128, u1_u10_u6_n129, u1_u10_u6_n130, u1_u10_u6_n131, u1_u10_u6_n132, 
       u1_u10_u6_n133, u1_u10_u6_n134, u1_u10_u6_n135, u1_u10_u6_n136, u1_u10_u6_n137, u1_u10_u6_n138, u1_u10_u6_n139, u1_u10_u6_n140, u1_u10_u6_n141, 
       u1_u10_u6_n142, u1_u10_u6_n143, u1_u10_u6_n144, u1_u10_u6_n145, u1_u10_u6_n146, u1_u10_u6_n147, u1_u10_u6_n148, u1_u10_u6_n149, u1_u10_u6_n150, 
       u1_u10_u6_n151, u1_u10_u6_n152, u1_u10_u6_n153, u1_u10_u6_n154, u1_u10_u6_n155, u1_u10_u6_n156, u1_u10_u6_n157, u1_u10_u6_n158, u1_u10_u6_n159, 
       u1_u10_u6_n160, u1_u10_u6_n161, u1_u10_u6_n162, u1_u10_u6_n163, u1_u10_u6_n164, u1_u10_u6_n165, u1_u10_u6_n166, u1_u10_u6_n167, u1_u10_u6_n168, 
       u1_u10_u6_n169, u1_u10_u6_n170, u1_u10_u6_n171, u1_u10_u6_n172, u1_u10_u6_n173, u1_u10_u6_n174, u1_u10_u6_n88, u1_u10_u6_n89, u1_u10_u6_n90, 
       u1_u10_u6_n91, u1_u10_u6_n92, u1_u10_u6_n93, u1_u10_u6_n94, u1_u10_u6_n95, u1_u10_u6_n96, u1_u10_u6_n97, u1_u10_u6_n98, u1_u10_u6_n99, 
       u1_u11_X_1, u1_u11_X_2, u1_u11_X_3, u1_u11_X_4, u1_u11_X_5, u1_u11_X_6, u1_u11_u0_n100, u1_u11_u0_n101, u1_u11_u0_n102, 
       u1_u11_u0_n103, u1_u11_u0_n104, u1_u11_u0_n105, u1_u11_u0_n106, u1_u11_u0_n107, u1_u11_u0_n108, u1_u11_u0_n109, u1_u11_u0_n110, u1_u11_u0_n111, 
       u1_u11_u0_n112, u1_u11_u0_n113, u1_u11_u0_n114, u1_u11_u0_n115, u1_u11_u0_n116, u1_u11_u0_n117, u1_u11_u0_n118, u1_u11_u0_n119, u1_u11_u0_n120, 
       u1_u11_u0_n121, u1_u11_u0_n122, u1_u11_u0_n123, u1_u11_u0_n124, u1_u11_u0_n125, u1_u11_u0_n126, u1_u11_u0_n127, u1_u11_u0_n128, u1_u11_u0_n129, 
       u1_u11_u0_n130, u1_u11_u0_n131, u1_u11_u0_n132, u1_u11_u0_n133, u1_u11_u0_n134, u1_u11_u0_n135, u1_u11_u0_n136, u1_u11_u0_n137, u1_u11_u0_n138, 
       u1_u11_u0_n139, u1_u11_u0_n140, u1_u11_u0_n141, u1_u11_u0_n142, u1_u11_u0_n143, u1_u11_u0_n144, u1_u11_u0_n145, u1_u11_u0_n146, u1_u11_u0_n147, 
       u1_u11_u0_n148, u1_u11_u0_n149, u1_u11_u0_n150, u1_u11_u0_n151, u1_u11_u0_n152, u1_u11_u0_n153, u1_u11_u0_n154, u1_u11_u0_n155, u1_u11_u0_n156, 
       u1_u11_u0_n157, u1_u11_u0_n158, u1_u11_u0_n159, u1_u11_u0_n160, u1_u11_u0_n161, u1_u11_u0_n162, u1_u11_u0_n163, u1_u11_u0_n164, u1_u11_u0_n165, 
       u1_u11_u0_n166, u1_u11_u0_n167, u1_u11_u0_n168, u1_u11_u0_n169, u1_u11_u0_n170, u1_u11_u0_n171, u1_u11_u0_n172, u1_u11_u0_n173, u1_u11_u0_n174, 
       u1_u11_u0_n88, u1_u11_u0_n89, u1_u11_u0_n90, u1_u11_u0_n91, u1_u11_u0_n92, u1_u11_u0_n93, u1_u11_u0_n94, u1_u11_u0_n95, u1_u11_u0_n96, 
       u1_u11_u0_n97, u1_u11_u0_n98, u1_u11_u0_n99, u1_u14_X_1, u1_u14_X_10, u1_u14_X_11, u1_u14_X_12, u1_u14_X_13, u1_u14_X_14, 
       u1_u14_X_15, u1_u14_X_16, u1_u14_X_17, u1_u14_X_18, u1_u14_X_19, u1_u14_X_2, u1_u14_X_20, u1_u14_X_21, u1_u14_X_22, 
       u1_u14_X_23, u1_u14_X_24, u1_u14_X_25, u1_u14_X_26, u1_u14_X_27, u1_u14_X_28, u1_u14_X_29, u1_u14_X_3, u1_u14_X_30, 
       u1_u14_X_4, u1_u14_X_5, u1_u14_X_6, u1_u14_X_7, u1_u14_X_8, u1_u14_X_9, u1_u14_u0_n100, u1_u14_u0_n101, u1_u14_u0_n102, 
       u1_u14_u0_n103, u1_u14_u0_n104, u1_u14_u0_n105, u1_u14_u0_n106, u1_u14_u0_n107, u1_u14_u0_n108, u1_u14_u0_n109, u1_u14_u0_n110, u1_u14_u0_n111, 
       u1_u14_u0_n112, u1_u14_u0_n113, u1_u14_u0_n114, u1_u14_u0_n115, u1_u14_u0_n116, u1_u14_u0_n117, u1_u14_u0_n118, u1_u14_u0_n119, u1_u14_u0_n120, 
       u1_u14_u0_n121, u1_u14_u0_n122, u1_u14_u0_n123, u1_u14_u0_n124, u1_u14_u0_n125, u1_u14_u0_n126, u1_u14_u0_n127, u1_u14_u0_n128, u1_u14_u0_n129, 
       u1_u14_u0_n130, u1_u14_u0_n131, u1_u14_u0_n132, u1_u14_u0_n133, u1_u14_u0_n134, u1_u14_u0_n135, u1_u14_u0_n136, u1_u14_u0_n137, u1_u14_u0_n138, 
       u1_u14_u0_n139, u1_u14_u0_n140, u1_u14_u0_n141, u1_u14_u0_n142, u1_u14_u0_n143, u1_u14_u0_n144, u1_u14_u0_n145, u1_u14_u0_n146, u1_u14_u0_n147, 
       u1_u14_u0_n148, u1_u14_u0_n149, u1_u14_u0_n150, u1_u14_u0_n151, u1_u14_u0_n152, u1_u14_u0_n153, u1_u14_u0_n154, u1_u14_u0_n155, u1_u14_u0_n156, 
       u1_u14_u0_n157, u1_u14_u0_n158, u1_u14_u0_n159, u1_u14_u0_n160, u1_u14_u0_n161, u1_u14_u0_n162, u1_u14_u0_n163, u1_u14_u0_n164, u1_u14_u0_n165, 
       u1_u14_u0_n166, u1_u14_u0_n167, u1_u14_u0_n168, u1_u14_u0_n169, u1_u14_u0_n170, u1_u14_u0_n171, u1_u14_u0_n172, u1_u14_u0_n173, u1_u14_u0_n174, 
       u1_u14_u0_n88, u1_u14_u0_n89, u1_u14_u0_n90, u1_u14_u0_n91, u1_u14_u0_n92, u1_u14_u0_n93, u1_u14_u0_n94, u1_u14_u0_n95, u1_u14_u0_n96, 
       u1_u14_u0_n97, u1_u14_u0_n98, u1_u14_u0_n99, u1_u14_u1_n100, u1_u14_u1_n101, u1_u14_u1_n102, u1_u14_u1_n103, u1_u14_u1_n104, u1_u14_u1_n105, 
       u1_u14_u1_n106, u1_u14_u1_n107, u1_u14_u1_n108, u1_u14_u1_n109, u1_u14_u1_n110, u1_u14_u1_n111, u1_u14_u1_n112, u1_u14_u1_n113, u1_u14_u1_n114, 
       u1_u14_u1_n115, u1_u14_u1_n116, u1_u14_u1_n117, u1_u14_u1_n118, u1_u14_u1_n119, u1_u14_u1_n120, u1_u14_u1_n121, u1_u14_u1_n122, u1_u14_u1_n123, 
       u1_u14_u1_n124, u1_u14_u1_n125, u1_u14_u1_n126, u1_u14_u1_n127, u1_u14_u1_n128, u1_u14_u1_n129, u1_u14_u1_n130, u1_u14_u1_n131, u1_u14_u1_n132, 
       u1_u14_u1_n133, u1_u14_u1_n134, u1_u14_u1_n135, u1_u14_u1_n136, u1_u14_u1_n137, u1_u14_u1_n138, u1_u14_u1_n139, u1_u14_u1_n140, u1_u14_u1_n141, 
       u1_u14_u1_n142, u1_u14_u1_n143, u1_u14_u1_n144, u1_u14_u1_n145, u1_u14_u1_n146, u1_u14_u1_n147, u1_u14_u1_n148, u1_u14_u1_n149, u1_u14_u1_n150, 
       u1_u14_u1_n151, u1_u14_u1_n152, u1_u14_u1_n153, u1_u14_u1_n154, u1_u14_u1_n155, u1_u14_u1_n156, u1_u14_u1_n157, u1_u14_u1_n158, u1_u14_u1_n159, 
       u1_u14_u1_n160, u1_u14_u1_n161, u1_u14_u1_n162, u1_u14_u1_n163, u1_u14_u1_n164, u1_u14_u1_n165, u1_u14_u1_n166, u1_u14_u1_n167, u1_u14_u1_n168, 
       u1_u14_u1_n169, u1_u14_u1_n170, u1_u14_u1_n171, u1_u14_u1_n172, u1_u14_u1_n173, u1_u14_u1_n174, u1_u14_u1_n175, u1_u14_u1_n176, u1_u14_u1_n177, 
       u1_u14_u1_n178, u1_u14_u1_n179, u1_u14_u1_n180, u1_u14_u1_n181, u1_u14_u1_n182, u1_u14_u1_n183, u1_u14_u1_n184, u1_u14_u1_n185, u1_u14_u1_n186, 
       u1_u14_u1_n187, u1_u14_u1_n188, u1_u14_u1_n95, u1_u14_u1_n96, u1_u14_u1_n97, u1_u14_u1_n98, u1_u14_u1_n99, u1_u14_u2_n100, u1_u14_u2_n101, 
       u1_u14_u2_n102, u1_u14_u2_n103, u1_u14_u2_n104, u1_u14_u2_n105, u1_u14_u2_n106, u1_u14_u2_n107, u1_u14_u2_n108, u1_u14_u2_n109, u1_u14_u2_n110, 
       u1_u14_u2_n111, u1_u14_u2_n112, u1_u14_u2_n113, u1_u14_u2_n114, u1_u14_u2_n115, u1_u14_u2_n116, u1_u14_u2_n117, u1_u14_u2_n118, u1_u14_u2_n119, 
       u1_u14_u2_n120, u1_u14_u2_n121, u1_u14_u2_n122, u1_u14_u2_n123, u1_u14_u2_n124, u1_u14_u2_n125, u1_u14_u2_n126, u1_u14_u2_n127, u1_u14_u2_n128, 
       u1_u14_u2_n129, u1_u14_u2_n130, u1_u14_u2_n131, u1_u14_u2_n132, u1_u14_u2_n133, u1_u14_u2_n134, u1_u14_u2_n135, u1_u14_u2_n136, u1_u14_u2_n137, 
       u1_u14_u2_n138, u1_u14_u2_n139, u1_u14_u2_n140, u1_u14_u2_n141, u1_u14_u2_n142, u1_u14_u2_n143, u1_u14_u2_n144, u1_u14_u2_n145, u1_u14_u2_n146, 
       u1_u14_u2_n147, u1_u14_u2_n148, u1_u14_u2_n149, u1_u14_u2_n150, u1_u14_u2_n151, u1_u14_u2_n152, u1_u14_u2_n153, u1_u14_u2_n154, u1_u14_u2_n155, 
       u1_u14_u2_n156, u1_u14_u2_n157, u1_u14_u2_n158, u1_u14_u2_n159, u1_u14_u2_n160, u1_u14_u2_n161, u1_u14_u2_n162, u1_u14_u2_n163, u1_u14_u2_n164, 
       u1_u14_u2_n165, u1_u14_u2_n166, u1_u14_u2_n167, u1_u14_u2_n168, u1_u14_u2_n169, u1_u14_u2_n170, u1_u14_u2_n171, u1_u14_u2_n172, u1_u14_u2_n173, 
       u1_u14_u2_n174, u1_u14_u2_n175, u1_u14_u2_n176, u1_u14_u2_n177, u1_u14_u2_n178, u1_u14_u2_n179, u1_u14_u2_n180, u1_u14_u2_n181, u1_u14_u2_n182, 
       u1_u14_u2_n183, u1_u14_u2_n184, u1_u14_u2_n185, u1_u14_u2_n186, u1_u14_u2_n187, u1_u14_u2_n188, u1_u14_u2_n95, u1_u14_u2_n96, u1_u14_u2_n97, 
       u1_u14_u2_n98, u1_u14_u2_n99, u1_u14_u3_n100, u1_u14_u3_n101, u1_u14_u3_n102, u1_u14_u3_n103, u1_u14_u3_n104, u1_u14_u3_n105, u1_u14_u3_n106, 
       u1_u14_u3_n107, u1_u14_u3_n108, u1_u14_u3_n109, u1_u14_u3_n110, u1_u14_u3_n111, u1_u14_u3_n112, u1_u14_u3_n113, u1_u14_u3_n114, u1_u14_u3_n115, 
       u1_u14_u3_n116, u1_u14_u3_n117, u1_u14_u3_n118, u1_u14_u3_n119, u1_u14_u3_n120, u1_u14_u3_n121, u1_u14_u3_n122, u1_u14_u3_n123, u1_u14_u3_n124, 
       u1_u14_u3_n125, u1_u14_u3_n126, u1_u14_u3_n127, u1_u14_u3_n128, u1_u14_u3_n129, u1_u14_u3_n130, u1_u14_u3_n131, u1_u14_u3_n132, u1_u14_u3_n133, 
       u1_u14_u3_n134, u1_u14_u3_n135, u1_u14_u3_n136, u1_u14_u3_n137, u1_u14_u3_n138, u1_u14_u3_n139, u1_u14_u3_n140, u1_u14_u3_n141, u1_u14_u3_n142, 
       u1_u14_u3_n143, u1_u14_u3_n144, u1_u14_u3_n145, u1_u14_u3_n146, u1_u14_u3_n147, u1_u14_u3_n148, u1_u14_u3_n149, u1_u14_u3_n150, u1_u14_u3_n151, 
       u1_u14_u3_n152, u1_u14_u3_n153, u1_u14_u3_n154, u1_u14_u3_n155, u1_u14_u3_n156, u1_u14_u3_n157, u1_u14_u3_n158, u1_u14_u3_n159, u1_u14_u3_n160, 
       u1_u14_u3_n161, u1_u14_u3_n162, u1_u14_u3_n163, u1_u14_u3_n164, u1_u14_u3_n165, u1_u14_u3_n166, u1_u14_u3_n167, u1_u14_u3_n168, u1_u14_u3_n169, 
       u1_u14_u3_n170, u1_u14_u3_n171, u1_u14_u3_n172, u1_u14_u3_n173, u1_u14_u3_n174, u1_u14_u3_n175, u1_u14_u3_n176, u1_u14_u3_n177, u1_u14_u3_n178, 
       u1_u14_u3_n179, u1_u14_u3_n180, u1_u14_u3_n181, u1_u14_u3_n182, u1_u14_u3_n183, u1_u14_u3_n184, u1_u14_u3_n185, u1_u14_u3_n186, u1_u14_u3_n94, 
       u1_u14_u3_n95, u1_u14_u3_n96, u1_u14_u3_n97, u1_u14_u3_n98, u1_u14_u3_n99, u1_u14_u4_n100, u1_u14_u4_n101, u1_u14_u4_n102, u1_u14_u4_n103, 
       u1_u14_u4_n104, u1_u14_u4_n105, u1_u14_u4_n106, u1_u14_u4_n107, u1_u14_u4_n108, u1_u14_u4_n109, u1_u14_u4_n110, u1_u14_u4_n111, u1_u14_u4_n112, 
       u1_u14_u4_n113, u1_u14_u4_n114, u1_u14_u4_n115, u1_u14_u4_n116, u1_u14_u4_n117, u1_u14_u4_n118, u1_u14_u4_n119, u1_u14_u4_n120, u1_u14_u4_n121, 
       u1_u14_u4_n122, u1_u14_u4_n123, u1_u14_u4_n124, u1_u14_u4_n125, u1_u14_u4_n126, u1_u14_u4_n127, u1_u14_u4_n128, u1_u14_u4_n129, u1_u14_u4_n130, 
       u1_u14_u4_n131, u1_u14_u4_n132, u1_u14_u4_n133, u1_u14_u4_n134, u1_u14_u4_n135, u1_u14_u4_n136, u1_u14_u4_n137, u1_u14_u4_n138, u1_u14_u4_n139, 
       u1_u14_u4_n140, u1_u14_u4_n141, u1_u14_u4_n142, u1_u14_u4_n143, u1_u14_u4_n144, u1_u14_u4_n145, u1_u14_u4_n146, u1_u14_u4_n147, u1_u14_u4_n148, 
       u1_u14_u4_n149, u1_u14_u4_n150, u1_u14_u4_n151, u1_u14_u4_n152, u1_u14_u4_n153, u1_u14_u4_n154, u1_u14_u4_n155, u1_u14_u4_n156, u1_u14_u4_n157, 
       u1_u14_u4_n158, u1_u14_u4_n159, u1_u14_u4_n160, u1_u14_u4_n161, u1_u14_u4_n162, u1_u14_u4_n163, u1_u14_u4_n164, u1_u14_u4_n165, u1_u14_u4_n166, 
       u1_u14_u4_n167, u1_u14_u4_n168, u1_u14_u4_n169, u1_u14_u4_n170, u1_u14_u4_n171, u1_u14_u4_n172, u1_u14_u4_n173, u1_u14_u4_n174, u1_u14_u4_n175, 
       u1_u14_u4_n176, u1_u14_u4_n177, u1_u14_u4_n178, u1_u14_u4_n179, u1_u14_u4_n180, u1_u14_u4_n181, u1_u14_u4_n182, u1_u14_u4_n183, u1_u14_u4_n184, 
       u1_u14_u4_n185, u1_u14_u4_n186, u1_u14_u4_n94, u1_u14_u4_n95, u1_u14_u4_n96, u1_u14_u4_n97, u1_u14_u4_n98, u1_u14_u4_n99, u1_u15_X_25, 
       u1_u15_X_26, u1_u15_X_27, u1_u15_X_28, u1_u15_X_29, u1_u15_X_30, u1_u15_X_31, u1_u15_X_32, u1_u15_X_33, u1_u15_X_34, 
       u1_u15_X_35, u1_u15_X_36, u1_u15_X_37, u1_u15_X_38, u1_u15_X_39, u1_u15_X_40, u1_u15_X_41, u1_u15_X_42, u1_u15_X_43, 
       u1_u15_X_44, u1_u15_X_45, u1_u15_X_46, u1_u15_X_47, u1_u15_X_48, u1_u15_u4_n100, u1_u15_u4_n101, u1_u15_u4_n102, u1_u15_u4_n103, 
       u1_u15_u4_n104, u1_u15_u4_n105, u1_u15_u4_n106, u1_u15_u4_n107, u1_u15_u4_n108, u1_u15_u4_n109, u1_u15_u4_n110, u1_u15_u4_n111, u1_u15_u4_n112, 
       u1_u15_u4_n113, u1_u15_u4_n114, u1_u15_u4_n115, u1_u15_u4_n116, u1_u15_u4_n117, u1_u15_u4_n118, u1_u15_u4_n119, u1_u15_u4_n120, u1_u15_u4_n121, 
       u1_u15_u4_n122, u1_u15_u4_n123, u1_u15_u4_n124, u1_u15_u4_n125, u1_u15_u4_n126, u1_u15_u4_n127, u1_u15_u4_n128, u1_u15_u4_n129, u1_u15_u4_n130, 
       u1_u15_u4_n131, u1_u15_u4_n132, u1_u15_u4_n133, u1_u15_u4_n134, u1_u15_u4_n135, u1_u15_u4_n136, u1_u15_u4_n137, u1_u15_u4_n138, u1_u15_u4_n139, 
       u1_u15_u4_n140, u1_u15_u4_n141, u1_u15_u4_n142, u1_u15_u4_n143, u1_u15_u4_n144, u1_u15_u4_n145, u1_u15_u4_n146, u1_u15_u4_n147, u1_u15_u4_n148, 
       u1_u15_u4_n149, u1_u15_u4_n150, u1_u15_u4_n151, u1_u15_u4_n152, u1_u15_u4_n153, u1_u15_u4_n154, u1_u15_u4_n155, u1_u15_u4_n156, u1_u15_u4_n157, 
       u1_u15_u4_n158, u1_u15_u4_n159, u1_u15_u4_n160, u1_u15_u4_n161, u1_u15_u4_n162, u1_u15_u4_n163, u1_u15_u4_n164, u1_u15_u4_n165, u1_u15_u4_n166, 
       u1_u15_u4_n167, u1_u15_u4_n168, u1_u15_u4_n169, u1_u15_u4_n170, u1_u15_u4_n171, u1_u15_u4_n172, u1_u15_u4_n173, u1_u15_u4_n174, u1_u15_u4_n175, 
       u1_u15_u4_n176, u1_u15_u4_n177, u1_u15_u4_n178, u1_u15_u4_n179, u1_u15_u4_n180, u1_u15_u4_n181, u1_u15_u4_n182, u1_u15_u4_n183, u1_u15_u4_n184, 
       u1_u15_u4_n185, u1_u15_u4_n186, u1_u15_u4_n94, u1_u15_u4_n95, u1_u15_u4_n96, u1_u15_u4_n97, u1_u15_u4_n98, u1_u15_u4_n99, u1_u15_u5_n100, 
       u1_u15_u5_n101, u1_u15_u5_n102, u1_u15_u5_n103, u1_u15_u5_n104, u1_u15_u5_n105, u1_u15_u5_n106, u1_u15_u5_n107, u1_u15_u5_n108, u1_u15_u5_n109, 
       u1_u15_u5_n110, u1_u15_u5_n111, u1_u15_u5_n112, u1_u15_u5_n113, u1_u15_u5_n114, u1_u15_u5_n115, u1_u15_u5_n116, u1_u15_u5_n117, u1_u15_u5_n118, 
       u1_u15_u5_n119, u1_u15_u5_n120, u1_u15_u5_n121, u1_u15_u5_n122, u1_u15_u5_n123, u1_u15_u5_n124, u1_u15_u5_n125, u1_u15_u5_n126, u1_u15_u5_n127, 
       u1_u15_u5_n128, u1_u15_u5_n129, u1_u15_u5_n130, u1_u15_u5_n131, u1_u15_u5_n132, u1_u15_u5_n133, u1_u15_u5_n134, u1_u15_u5_n135, u1_u15_u5_n136, 
       u1_u15_u5_n137, u1_u15_u5_n138, u1_u15_u5_n139, u1_u15_u5_n140, u1_u15_u5_n141, u1_u15_u5_n142, u1_u15_u5_n143, u1_u15_u5_n144, u1_u15_u5_n145, 
       u1_u15_u5_n146, u1_u15_u5_n147, u1_u15_u5_n148, u1_u15_u5_n149, u1_u15_u5_n150, u1_u15_u5_n151, u1_u15_u5_n152, u1_u15_u5_n153, u1_u15_u5_n154, 
       u1_u15_u5_n155, u1_u15_u5_n156, u1_u15_u5_n157, u1_u15_u5_n158, u1_u15_u5_n159, u1_u15_u5_n160, u1_u15_u5_n161, u1_u15_u5_n162, u1_u15_u5_n163, 
       u1_u15_u5_n164, u1_u15_u5_n165, u1_u15_u5_n166, u1_u15_u5_n167, u1_u15_u5_n168, u1_u15_u5_n169, u1_u15_u5_n170, u1_u15_u5_n171, u1_u15_u5_n172, 
       u1_u15_u5_n173, u1_u15_u5_n174, u1_u15_u5_n175, u1_u15_u5_n176, u1_u15_u5_n177, u1_u15_u5_n178, u1_u15_u5_n179, u1_u15_u5_n180, u1_u15_u5_n181, 
       u1_u15_u5_n182, u1_u15_u5_n183, u1_u15_u5_n184, u1_u15_u5_n185, u1_u15_u5_n186, u1_u15_u5_n187, u1_u15_u5_n188, u1_u15_u5_n189, u1_u15_u5_n190, 
       u1_u15_u5_n191, u1_u15_u5_n192, u1_u15_u5_n193, u1_u15_u5_n194, u1_u15_u5_n195, u1_u15_u5_n196, u1_u15_u5_n99, u1_u15_u6_n100, u1_u15_u6_n101, 
       u1_u15_u6_n102, u1_u15_u6_n103, u1_u15_u6_n104, u1_u15_u6_n105, u1_u15_u6_n106, u1_u15_u6_n107, u1_u15_u6_n108, u1_u15_u6_n109, u1_u15_u6_n110, 
       u1_u15_u6_n111, u1_u15_u6_n112, u1_u15_u6_n113, u1_u15_u6_n114, u1_u15_u6_n115, u1_u15_u6_n116, u1_u15_u6_n117, u1_u15_u6_n118, u1_u15_u6_n119, 
       u1_u15_u6_n120, u1_u15_u6_n121, u1_u15_u6_n122, u1_u15_u6_n123, u1_u15_u6_n124, u1_u15_u6_n125, u1_u15_u6_n126, u1_u15_u6_n127, u1_u15_u6_n128, 
       u1_u15_u6_n129, u1_u15_u6_n130, u1_u15_u6_n131, u1_u15_u6_n132, u1_u15_u6_n133, u1_u15_u6_n134, u1_u15_u6_n135, u1_u15_u6_n136, u1_u15_u6_n137, 
       u1_u15_u6_n138, u1_u15_u6_n139, u1_u15_u6_n140, u1_u15_u6_n141, u1_u15_u6_n142, u1_u15_u6_n143, u1_u15_u6_n144, u1_u15_u6_n145, u1_u15_u6_n146, 
       u1_u15_u6_n147, u1_u15_u6_n148, u1_u15_u6_n149, u1_u15_u6_n150, u1_u15_u6_n151, u1_u15_u6_n152, u1_u15_u6_n153, u1_u15_u6_n154, u1_u15_u6_n155, 
       u1_u15_u6_n156, u1_u15_u6_n157, u1_u15_u6_n158, u1_u15_u6_n159, u1_u15_u6_n160, u1_u15_u6_n161, u1_u15_u6_n162, u1_u15_u6_n163, u1_u15_u6_n164, 
       u1_u15_u6_n165, u1_u15_u6_n166, u1_u15_u6_n167, u1_u15_u6_n168, u1_u15_u6_n169, u1_u15_u6_n170, u1_u15_u6_n171, u1_u15_u6_n172, u1_u15_u6_n173, 
       u1_u15_u6_n174, u1_u15_u6_n88, u1_u15_u6_n89, u1_u15_u6_n90, u1_u15_u6_n91, u1_u15_u6_n92, u1_u15_u6_n93, u1_u15_u6_n94, u1_u15_u6_n95, 
       u1_u15_u6_n96, u1_u15_u6_n97, u1_u15_u6_n98, u1_u15_u6_n99, u1_u15_u7_n100, u1_u15_u7_n101, u1_u15_u7_n102, u1_u15_u7_n103, u1_u15_u7_n104, 
       u1_u15_u7_n105, u1_u15_u7_n106, u1_u15_u7_n107, u1_u15_u7_n108, u1_u15_u7_n109, u1_u15_u7_n110, u1_u15_u7_n111, u1_u15_u7_n112, u1_u15_u7_n113, 
       u1_u15_u7_n114, u1_u15_u7_n115, u1_u15_u7_n116, u1_u15_u7_n117, u1_u15_u7_n118, u1_u15_u7_n119, u1_u15_u7_n120, u1_u15_u7_n121, u1_u15_u7_n122, 
       u1_u15_u7_n123, u1_u15_u7_n124, u1_u15_u7_n125, u1_u15_u7_n126, u1_u15_u7_n127, u1_u15_u7_n128, u1_u15_u7_n129, u1_u15_u7_n130, u1_u15_u7_n131, 
       u1_u15_u7_n132, u1_u15_u7_n133, u1_u15_u7_n134, u1_u15_u7_n135, u1_u15_u7_n136, u1_u15_u7_n137, u1_u15_u7_n138, u1_u15_u7_n139, u1_u15_u7_n140, 
       u1_u15_u7_n141, u1_u15_u7_n142, u1_u15_u7_n143, u1_u15_u7_n144, u1_u15_u7_n145, u1_u15_u7_n146, u1_u15_u7_n147, u1_u15_u7_n148, u1_u15_u7_n149, 
       u1_u15_u7_n150, u1_u15_u7_n151, u1_u15_u7_n152, u1_u15_u7_n153, u1_u15_u7_n154, u1_u15_u7_n155, u1_u15_u7_n156, u1_u15_u7_n157, u1_u15_u7_n158, 
       u1_u15_u7_n159, u1_u15_u7_n160, u1_u15_u7_n161, u1_u15_u7_n162, u1_u15_u7_n163, u1_u15_u7_n164, u1_u15_u7_n165, u1_u15_u7_n166, u1_u15_u7_n167, 
       u1_u15_u7_n168, u1_u15_u7_n169, u1_u15_u7_n170, u1_u15_u7_n171, u1_u15_u7_n172, u1_u15_u7_n173, u1_u15_u7_n174, u1_u15_u7_n175, u1_u15_u7_n176, 
       u1_u15_u7_n177, u1_u15_u7_n178, u1_u15_u7_n179, u1_u15_u7_n180, u1_u15_u7_n91, u1_u15_u7_n92, u1_u15_u7_n93, u1_u15_u7_n94, u1_u15_u7_n95, 
       u1_u15_u7_n96, u1_u15_u7_n97, u1_u15_u7_n98, u1_u15_u7_n99, u1_u1_X_1, u1_u1_X_2, u1_u1_X_3, u1_u1_X_4, u1_u1_X_5, 
       u1_u1_X_6, u1_u1_u0_n100, u1_u1_u0_n101, u1_u1_u0_n102, u1_u1_u0_n103, u1_u1_u0_n104, u1_u1_u0_n105, u1_u1_u0_n106, u1_u1_u0_n107, 
       u1_u1_u0_n108, u1_u1_u0_n109, u1_u1_u0_n110, u1_u1_u0_n111, u1_u1_u0_n112, u1_u1_u0_n113, u1_u1_u0_n114, u1_u1_u0_n115, u1_u1_u0_n116, 
       u1_u1_u0_n117, u1_u1_u0_n118, u1_u1_u0_n119, u1_u1_u0_n120, u1_u1_u0_n121, u1_u1_u0_n122, u1_u1_u0_n123, u1_u1_u0_n124, u1_u1_u0_n125, 
       u1_u1_u0_n126, u1_u1_u0_n127, u1_u1_u0_n128, u1_u1_u0_n129, u1_u1_u0_n130, u1_u1_u0_n131, u1_u1_u0_n132, u1_u1_u0_n133, u1_u1_u0_n134, 
       u1_u1_u0_n135, u1_u1_u0_n136, u1_u1_u0_n137, u1_u1_u0_n138, u1_u1_u0_n139, u1_u1_u0_n140, u1_u1_u0_n141, u1_u1_u0_n142, u1_u1_u0_n143, 
       u1_u1_u0_n144, u1_u1_u0_n145, u1_u1_u0_n146, u1_u1_u0_n147, u1_u1_u0_n148, u1_u1_u0_n149, u1_u1_u0_n150, u1_u1_u0_n151, u1_u1_u0_n152, 
       u1_u1_u0_n153, u1_u1_u0_n154, u1_u1_u0_n155, u1_u1_u0_n156, u1_u1_u0_n157, u1_u1_u0_n158, u1_u1_u0_n159, u1_u1_u0_n160, u1_u1_u0_n161, 
       u1_u1_u0_n162, u1_u1_u0_n163, u1_u1_u0_n164, u1_u1_u0_n165, u1_u1_u0_n166, u1_u1_u0_n167, u1_u1_u0_n168, u1_u1_u0_n169, u1_u1_u0_n170, 
       u1_u1_u0_n171, u1_u1_u0_n172, u1_u1_u0_n173, u1_u1_u0_n174, u1_u1_u0_n88, u1_u1_u0_n89, u1_u1_u0_n90, u1_u1_u0_n91, u1_u1_u0_n92, 
       u1_u1_u0_n93, u1_u1_u0_n94, u1_u1_u0_n95, u1_u1_u0_n96, u1_u1_u0_n97, u1_u1_u0_n98, u1_u1_u0_n99, u1_u3_X_31, u1_u3_X_32, 
       u1_u3_X_33, u1_u3_X_34, u1_u3_X_35, u1_u3_X_36, u1_u3_X_37, u1_u3_X_38, u1_u3_X_39, u1_u3_X_40, u1_u3_X_41, 
       u1_u3_X_42, u1_u3_u5_n100, u1_u3_u5_n101, u1_u3_u5_n102, u1_u3_u5_n103, u1_u3_u5_n104, u1_u3_u5_n105, u1_u3_u5_n106, u1_u3_u5_n107, 
       u1_u3_u5_n108, u1_u3_u5_n109, u1_u3_u5_n110, u1_u3_u5_n111, u1_u3_u5_n112, u1_u3_u5_n113, u1_u3_u5_n114, u1_u3_u5_n115, u1_u3_u5_n116, 
       u1_u3_u5_n117, u1_u3_u5_n118, u1_u3_u5_n119, u1_u3_u5_n120, u1_u3_u5_n121, u1_u3_u5_n122, u1_u3_u5_n123, u1_u3_u5_n124, u1_u3_u5_n125, 
       u1_u3_u5_n126, u1_u3_u5_n127, u1_u3_u5_n128, u1_u3_u5_n129, u1_u3_u5_n130, u1_u3_u5_n131, u1_u3_u5_n132, u1_u3_u5_n133, u1_u3_u5_n134, 
       u1_u3_u5_n135, u1_u3_u5_n136, u1_u3_u5_n137, u1_u3_u5_n138, u1_u3_u5_n139, u1_u3_u5_n140, u1_u3_u5_n141, u1_u3_u5_n142, u1_u3_u5_n143, 
       u1_u3_u5_n144, u1_u3_u5_n145, u1_u3_u5_n146, u1_u3_u5_n147, u1_u3_u5_n148, u1_u3_u5_n149, u1_u3_u5_n150, u1_u3_u5_n151, u1_u3_u5_n152, 
       u1_u3_u5_n153, u1_u3_u5_n154, u1_u3_u5_n155, u1_u3_u5_n156, u1_u3_u5_n157, u1_u3_u5_n158, u1_u3_u5_n159, u1_u3_u5_n160, u1_u3_u5_n161, 
       u1_u3_u5_n162, u1_u3_u5_n163, u1_u3_u5_n164, u1_u3_u5_n165, u1_u3_u5_n166, u1_u3_u5_n167, u1_u3_u5_n168, u1_u3_u5_n169, u1_u3_u5_n170, 
       u1_u3_u5_n171, u1_u3_u5_n172, u1_u3_u5_n173, u1_u3_u5_n174, u1_u3_u5_n175, u1_u3_u5_n176, u1_u3_u5_n177, u1_u3_u5_n178, u1_u3_u5_n179, 
       u1_u3_u5_n180, u1_u3_u5_n181, u1_u3_u5_n182, u1_u3_u5_n183, u1_u3_u5_n184, u1_u3_u5_n185, u1_u3_u5_n186, u1_u3_u5_n187, u1_u3_u5_n188, 
       u1_u3_u5_n189, u1_u3_u5_n190, u1_u3_u5_n191, u1_u3_u5_n192, u1_u3_u5_n193, u1_u3_u5_n194, u1_u3_u5_n195, u1_u3_u5_n196, u1_u3_u5_n99, 
       u1_u3_u6_n100, u1_u3_u6_n101, u1_u3_u6_n102, u1_u3_u6_n103, u1_u3_u6_n104, u1_u3_u6_n105, u1_u3_u6_n106, u1_u3_u6_n107, u1_u3_u6_n108, 
       u1_u3_u6_n109, u1_u3_u6_n110, u1_u3_u6_n111, u1_u3_u6_n112, u1_u3_u6_n113, u1_u3_u6_n114, u1_u3_u6_n115, u1_u3_u6_n116, u1_u3_u6_n117, 
       u1_u3_u6_n118, u1_u3_u6_n119, u1_u3_u6_n120, u1_u3_u6_n121, u1_u3_u6_n122, u1_u3_u6_n123, u1_u3_u6_n124, u1_u3_u6_n125, u1_u3_u6_n126, 
       u1_u3_u6_n127, u1_u3_u6_n128, u1_u3_u6_n129, u1_u3_u6_n130, u1_u3_u6_n131, u1_u3_u6_n132, u1_u3_u6_n133, u1_u3_u6_n134, u1_u3_u6_n135, 
       u1_u3_u6_n136, u1_u3_u6_n137, u1_u3_u6_n138, u1_u3_u6_n139, u1_u3_u6_n140, u1_u3_u6_n141, u1_u3_u6_n142, u1_u3_u6_n143, u1_u3_u6_n144, 
       u1_u3_u6_n145, u1_u3_u6_n146, u1_u3_u6_n147, u1_u3_u6_n148, u1_u3_u6_n149, u1_u3_u6_n150, u1_u3_u6_n151, u1_u3_u6_n152, u1_u3_u6_n153, 
       u1_u3_u6_n154, u1_u3_u6_n155, u1_u3_u6_n156, u1_u3_u6_n157, u1_u3_u6_n158, u1_u3_u6_n159, u1_u3_u6_n160, u1_u3_u6_n161, u1_u3_u6_n162, 
       u1_u3_u6_n163, u1_u3_u6_n164, u1_u3_u6_n165, u1_u3_u6_n166, u1_u3_u6_n167, u1_u3_u6_n168, u1_u3_u6_n169, u1_u3_u6_n170, u1_u3_u6_n171, 
       u1_u3_u6_n172, u1_u3_u6_n173, u1_u3_u6_n174, u1_u3_u6_n88, u1_u3_u6_n89, u1_u3_u6_n90, u1_u3_u6_n91, u1_u3_u6_n92, u1_u3_u6_n93, 
       u1_u3_u6_n94, u1_u3_u6_n95, u1_u3_u6_n96, u1_u3_u6_n97, u1_u3_u6_n98, u1_u3_u6_n99, u1_u4_X_25, u1_u4_X_26, u1_u4_X_27, 
       u1_u4_X_28, u1_u4_X_29, u1_u4_X_30, u1_u4_X_43, u1_u4_X_44, u1_u4_X_45, u1_u4_X_46, u1_u4_X_47, u1_u4_X_48, 
       u1_u4_u4_n100, u1_u4_u4_n101, u1_u4_u4_n102, u1_u4_u4_n103, u1_u4_u4_n104, u1_u4_u4_n105, u1_u4_u4_n106, u1_u4_u4_n107, u1_u4_u4_n108, 
       u1_u4_u4_n109, u1_u4_u4_n110, u1_u4_u4_n111, u1_u4_u4_n112, u1_u4_u4_n113, u1_u4_u4_n114, u1_u4_u4_n115, u1_u4_u4_n116, u1_u4_u4_n117, 
       u1_u4_u4_n118, u1_u4_u4_n119, u1_u4_u4_n120, u1_u4_u4_n121, u1_u4_u4_n122, u1_u4_u4_n123, u1_u4_u4_n124, u1_u4_u4_n125, u1_u4_u4_n126, 
       u1_u4_u4_n127, u1_u4_u4_n128, u1_u4_u4_n129, u1_u4_u4_n130, u1_u4_u4_n131, u1_u4_u4_n132, u1_u4_u4_n133, u1_u4_u4_n134, u1_u4_u4_n135, 
       u1_u4_u4_n136, u1_u4_u4_n137, u1_u4_u4_n138, u1_u4_u4_n139, u1_u4_u4_n140, u1_u4_u4_n141, u1_u4_u4_n142, u1_u4_u4_n143, u1_u4_u4_n144, 
       u1_u4_u4_n145, u1_u4_u4_n146, u1_u4_u4_n147, u1_u4_u4_n148, u1_u4_u4_n149, u1_u4_u4_n150, u1_u4_u4_n151, u1_u4_u4_n152, u1_u4_u4_n153, 
       u1_u4_u4_n154, u1_u4_u4_n155, u1_u4_u4_n156, u1_u4_u4_n157, u1_u4_u4_n158, u1_u4_u4_n159, u1_u4_u4_n160, u1_u4_u4_n161, u1_u4_u4_n162, 
       u1_u4_u4_n163, u1_u4_u4_n164, u1_u4_u4_n165, u1_u4_u4_n166, u1_u4_u4_n167, u1_u4_u4_n168, u1_u4_u4_n169, u1_u4_u4_n170, u1_u4_u4_n171, 
       u1_u4_u4_n172, u1_u4_u4_n173, u1_u4_u4_n174, u1_u4_u4_n175, u1_u4_u4_n176, u1_u4_u4_n177, u1_u4_u4_n178, u1_u4_u4_n179, u1_u4_u4_n180, 
       u1_u4_u4_n181, u1_u4_u4_n182, u1_u4_u4_n183, u1_u4_u4_n184, u1_u4_u4_n185, u1_u4_u4_n186, u1_u4_u4_n94, u1_u4_u4_n95, u1_u4_u4_n96, 
       u1_u4_u4_n97, u1_u4_u4_n98, u1_u4_u4_n99, u1_u4_u7_n100, u1_u4_u7_n101, u1_u4_u7_n102, u1_u4_u7_n103, u1_u4_u7_n104, u1_u4_u7_n105, 
       u1_u4_u7_n106, u1_u4_u7_n107, u1_u4_u7_n108, u1_u4_u7_n109, u1_u4_u7_n110, u1_u4_u7_n111, u1_u4_u7_n112, u1_u4_u7_n113, u1_u4_u7_n114, 
       u1_u4_u7_n115, u1_u4_u7_n116, u1_u4_u7_n117, u1_u4_u7_n118, u1_u4_u7_n119, u1_u4_u7_n120, u1_u4_u7_n121, u1_u4_u7_n122, u1_u4_u7_n123, 
       u1_u4_u7_n124, u1_u4_u7_n125, u1_u4_u7_n126, u1_u4_u7_n127, u1_u4_u7_n128, u1_u4_u7_n129, u1_u4_u7_n130, u1_u4_u7_n131, u1_u4_u7_n132, 
       u1_u4_u7_n133, u1_u4_u7_n134, u1_u4_u7_n135, u1_u4_u7_n136, u1_u4_u7_n137, u1_u4_u7_n138, u1_u4_u7_n139, u1_u4_u7_n140, u1_u4_u7_n141, 
       u1_u4_u7_n142, u1_u4_u7_n143, u1_u4_u7_n144, u1_u4_u7_n145, u1_u4_u7_n146, u1_u4_u7_n147, u1_u4_u7_n148, u1_u4_u7_n149, u1_u4_u7_n150, 
       u1_u4_u7_n151, u1_u4_u7_n152, u1_u4_u7_n153, u1_u4_u7_n154, u1_u4_u7_n155, u1_u4_u7_n156, u1_u4_u7_n157, u1_u4_u7_n158, u1_u4_u7_n159, 
       u1_u4_u7_n160, u1_u4_u7_n161, u1_u4_u7_n162, u1_u4_u7_n163, u1_u4_u7_n164, u1_u4_u7_n165, u1_u4_u7_n166, u1_u4_u7_n167, u1_u4_u7_n168, 
       u1_u4_u7_n169, u1_u4_u7_n170, u1_u4_u7_n171, u1_u4_u7_n172, u1_u4_u7_n173, u1_u4_u7_n174, u1_u4_u7_n175, u1_u4_u7_n176, u1_u4_u7_n177, 
       u1_u4_u7_n178, u1_u4_u7_n179, u1_u4_u7_n180, u1_u4_u7_n91, u1_u4_u7_n92, u1_u4_u7_n93, u1_u4_u7_n94, u1_u4_u7_n95, u1_u4_u7_n96, 
       u1_u4_u7_n97, u1_u4_u7_n98, u1_u4_u7_n99, u1_u6_X_10, u1_u6_X_11, u1_u6_X_12, u1_u6_X_13, u1_u6_X_14, u1_u6_X_15, 
       u1_u6_X_16, u1_u6_X_17, u1_u6_X_18, u1_u6_X_37, u1_u6_X_38, u1_u6_X_39, u1_u6_X_40, u1_u6_X_41, u1_u6_X_42, 
       u1_u6_X_43, u1_u6_X_44, u1_u6_X_45, u1_u6_X_46, u1_u6_X_47, u1_u6_X_48, u1_u6_X_7, u1_u6_X_8, u1_u6_X_9, 
       u1_u6_u1_n100, u1_u6_u1_n101, u1_u6_u1_n102, u1_u6_u1_n103, u1_u6_u1_n104, u1_u6_u1_n105, u1_u6_u1_n106, u1_u6_u1_n107, u1_u6_u1_n108, 
       u1_u6_u1_n109, u1_u6_u1_n110, u1_u6_u1_n111, u1_u6_u1_n112, u1_u6_u1_n113, u1_u6_u1_n114, u1_u6_u1_n115, u1_u6_u1_n116, u1_u6_u1_n117, 
       u1_u6_u1_n118, u1_u6_u1_n119, u1_u6_u1_n120, u1_u6_u1_n121, u1_u6_u1_n122, u1_u6_u1_n123, u1_u6_u1_n124, u1_u6_u1_n125, u1_u6_u1_n126, 
       u1_u6_u1_n127, u1_u6_u1_n128, u1_u6_u1_n129, u1_u6_u1_n130, u1_u6_u1_n131, u1_u6_u1_n132, u1_u6_u1_n133, u1_u6_u1_n134, u1_u6_u1_n135, 
       u1_u6_u1_n136, u1_u6_u1_n137, u1_u6_u1_n138, u1_u6_u1_n139, u1_u6_u1_n140, u1_u6_u1_n141, u1_u6_u1_n142, u1_u6_u1_n143, u1_u6_u1_n144, 
       u1_u6_u1_n145, u1_u6_u1_n146, u1_u6_u1_n147, u1_u6_u1_n148, u1_u6_u1_n149, u1_u6_u1_n150, u1_u6_u1_n151, u1_u6_u1_n152, u1_u6_u1_n153, 
       u1_u6_u1_n154, u1_u6_u1_n155, u1_u6_u1_n156, u1_u6_u1_n157, u1_u6_u1_n158, u1_u6_u1_n159, u1_u6_u1_n160, u1_u6_u1_n161, u1_u6_u1_n162, 
       u1_u6_u1_n163, u1_u6_u1_n164, u1_u6_u1_n165, u1_u6_u1_n166, u1_u6_u1_n167, u1_u6_u1_n168, u1_u6_u1_n169, u1_u6_u1_n170, u1_u6_u1_n171, 
       u1_u6_u1_n172, u1_u6_u1_n173, u1_u6_u1_n174, u1_u6_u1_n175, u1_u6_u1_n176, u1_u6_u1_n177, u1_u6_u1_n178, u1_u6_u1_n179, u1_u6_u1_n180, 
       u1_u6_u1_n181, u1_u6_u1_n182, u1_u6_u1_n183, u1_u6_u1_n184, u1_u6_u1_n185, u1_u6_u1_n186, u1_u6_u1_n187, u1_u6_u1_n188, u1_u6_u1_n95, 
       u1_u6_u1_n96, u1_u6_u1_n97, u1_u6_u1_n98, u1_u6_u1_n99, u1_u6_u2_n100, u1_u6_u2_n101, u1_u6_u2_n102, u1_u6_u2_n103, u1_u6_u2_n104, 
       u1_u6_u2_n105, u1_u6_u2_n106, u1_u6_u2_n107, u1_u6_u2_n108, u1_u6_u2_n109, u1_u6_u2_n110, u1_u6_u2_n111, u1_u6_u2_n112, u1_u6_u2_n113, 
       u1_u6_u2_n114, u1_u6_u2_n115, u1_u6_u2_n116, u1_u6_u2_n117, u1_u6_u2_n118, u1_u6_u2_n119, u1_u6_u2_n120, u1_u6_u2_n121, u1_u6_u2_n122, 
       u1_u6_u2_n123, u1_u6_u2_n124, u1_u6_u2_n125, u1_u6_u2_n126, u1_u6_u2_n127, u1_u6_u2_n128, u1_u6_u2_n129, u1_u6_u2_n130, u1_u6_u2_n131, 
       u1_u6_u2_n132, u1_u6_u2_n133, u1_u6_u2_n134, u1_u6_u2_n135, u1_u6_u2_n136, u1_u6_u2_n137, u1_u6_u2_n138, u1_u6_u2_n139, u1_u6_u2_n140, 
       u1_u6_u2_n141, u1_u6_u2_n142, u1_u6_u2_n143, u1_u6_u2_n144, u1_u6_u2_n145, u1_u6_u2_n146, u1_u6_u2_n147, u1_u6_u2_n148, u1_u6_u2_n149, 
       u1_u6_u2_n150, u1_u6_u2_n151, u1_u6_u2_n152, u1_u6_u2_n153, u1_u6_u2_n154, u1_u6_u2_n155, u1_u6_u2_n156, u1_u6_u2_n157, u1_u6_u2_n158, 
       u1_u6_u2_n159, u1_u6_u2_n160, u1_u6_u2_n161, u1_u6_u2_n162, u1_u6_u2_n163, u1_u6_u2_n164, u1_u6_u2_n165, u1_u6_u2_n166, u1_u6_u2_n167, 
       u1_u6_u2_n168, u1_u6_u2_n169, u1_u6_u2_n170, u1_u6_u2_n171, u1_u6_u2_n172, u1_u6_u2_n173, u1_u6_u2_n174, u1_u6_u2_n175, u1_u6_u2_n176, 
       u1_u6_u2_n177, u1_u6_u2_n178, u1_u6_u2_n179, u1_u6_u2_n180, u1_u6_u2_n181, u1_u6_u2_n182, u1_u6_u2_n183, u1_u6_u2_n184, u1_u6_u2_n185, 
       u1_u6_u2_n186, u1_u6_u2_n187, u1_u6_u2_n188, u1_u6_u2_n95, u1_u6_u2_n96, u1_u6_u2_n97, u1_u6_u2_n98, u1_u6_u2_n99, u1_u6_u6_n100, 
       u1_u6_u6_n101, u1_u6_u6_n102, u1_u6_u6_n103, u1_u6_u6_n104, u1_u6_u6_n105, u1_u6_u6_n106, u1_u6_u6_n107, u1_u6_u6_n108, u1_u6_u6_n109, 
       u1_u6_u6_n110, u1_u6_u6_n111, u1_u6_u6_n112, u1_u6_u6_n113, u1_u6_u6_n114, u1_u6_u6_n115, u1_u6_u6_n116, u1_u6_u6_n117, u1_u6_u6_n118, 
       u1_u6_u6_n119, u1_u6_u6_n120, u1_u6_u6_n121, u1_u6_u6_n122, u1_u6_u6_n123, u1_u6_u6_n124, u1_u6_u6_n125, u1_u6_u6_n126, u1_u6_u6_n127, 
       u1_u6_u6_n128, u1_u6_u6_n129, u1_u6_u6_n130, u1_u6_u6_n131, u1_u6_u6_n132, u1_u6_u6_n133, u1_u6_u6_n134, u1_u6_u6_n135, u1_u6_u6_n136, 
       u1_u6_u6_n137, u1_u6_u6_n138, u1_u6_u6_n139, u1_u6_u6_n140, u1_u6_u6_n141, u1_u6_u6_n142, u1_u6_u6_n143, u1_u6_u6_n144, u1_u6_u6_n145, 
       u1_u6_u6_n146, u1_u6_u6_n147, u1_u6_u6_n148, u1_u6_u6_n149, u1_u6_u6_n150, u1_u6_u6_n151, u1_u6_u6_n152, u1_u6_u6_n153, u1_u6_u6_n154, 
       u1_u6_u6_n155, u1_u6_u6_n156, u1_u6_u6_n157, u1_u6_u6_n158, u1_u6_u6_n159, u1_u6_u6_n160, u1_u6_u6_n161, u1_u6_u6_n162, u1_u6_u6_n163, 
       u1_u6_u6_n164, u1_u6_u6_n165, u1_u6_u6_n166, u1_u6_u6_n167, u1_u6_u6_n168, u1_u6_u6_n169, u1_u6_u6_n170, u1_u6_u6_n171, u1_u6_u6_n172, 
       u1_u6_u6_n173, u1_u6_u6_n174, u1_u6_u6_n88, u1_u6_u6_n89, u1_u6_u6_n90, u1_u6_u6_n91, u1_u6_u6_n92, u1_u6_u6_n93, u1_u6_u6_n94, 
       u1_u6_u6_n95, u1_u6_u6_n96, u1_u6_u6_n97, u1_u6_u6_n98, u1_u6_u6_n99, u1_u6_u7_n100, u1_u6_u7_n101, u1_u6_u7_n102, u1_u6_u7_n103, 
       u1_u6_u7_n104, u1_u6_u7_n105, u1_u6_u7_n106, u1_u6_u7_n107, u1_u6_u7_n108, u1_u6_u7_n109, u1_u6_u7_n110, u1_u6_u7_n111, u1_u6_u7_n112, 
       u1_u6_u7_n113, u1_u6_u7_n114, u1_u6_u7_n115, u1_u6_u7_n116, u1_u6_u7_n117, u1_u6_u7_n118, u1_u6_u7_n119, u1_u6_u7_n120, u1_u6_u7_n121, 
       u1_u6_u7_n122, u1_u6_u7_n123, u1_u6_u7_n124, u1_u6_u7_n125, u1_u6_u7_n126, u1_u6_u7_n127, u1_u6_u7_n128, u1_u6_u7_n129, u1_u6_u7_n130, 
       u1_u6_u7_n131, u1_u6_u7_n132, u1_u6_u7_n133, u1_u6_u7_n134, u1_u6_u7_n135, u1_u6_u7_n136, u1_u6_u7_n137, u1_u6_u7_n138, u1_u6_u7_n139, 
       u1_u6_u7_n140, u1_u6_u7_n141, u1_u6_u7_n142, u1_u6_u7_n143, u1_u6_u7_n144, u1_u6_u7_n145, u1_u6_u7_n146, u1_u6_u7_n147, u1_u6_u7_n148, 
       u1_u6_u7_n149, u1_u6_u7_n150, u1_u6_u7_n151, u1_u6_u7_n152, u1_u6_u7_n153, u1_u6_u7_n154, u1_u6_u7_n155, u1_u6_u7_n156, u1_u6_u7_n157, 
       u1_u6_u7_n158, u1_u6_u7_n159, u1_u6_u7_n160, u1_u6_u7_n161, u1_u6_u7_n162, u1_u6_u7_n163, u1_u6_u7_n164, u1_u6_u7_n165, u1_u6_u7_n166, 
       u1_u6_u7_n167, u1_u6_u7_n168, u1_u6_u7_n169, u1_u6_u7_n170, u1_u6_u7_n171, u1_u6_u7_n172, u1_u6_u7_n173, u1_u6_u7_n174, u1_u6_u7_n175, 
       u1_u6_u7_n176, u1_u6_u7_n177, u1_u6_u7_n178, u1_u6_u7_n179, u1_u6_u7_n180, u1_u6_u7_n91, u1_u6_u7_n92, u1_u6_u7_n93, u1_u6_u7_n94, 
       u1_u6_u7_n95, u1_u6_u7_n96, u1_u6_u7_n97, u1_u6_u7_n98, u1_u6_u7_n99, u1_u7_X_1, u1_u7_X_10, u1_u7_X_11, u1_u7_X_12, 
       u1_u7_X_13, u1_u7_X_14, u1_u7_X_15, u1_u7_X_16, u1_u7_X_17, u1_u7_X_18, u1_u7_X_2, u1_u7_X_3, u1_u7_X_4, 
       u1_u7_X_5, u1_u7_X_6, u1_u7_X_7, u1_u7_X_8, u1_u7_X_9, u1_u7_u0_n100, u1_u7_u0_n101, u1_u7_u0_n102, u1_u7_u0_n103, 
       u1_u7_u0_n104, u1_u7_u0_n105, u1_u7_u0_n106, u1_u7_u0_n107, u1_u7_u0_n108, u1_u7_u0_n109, u1_u7_u0_n110, u1_u7_u0_n111, u1_u7_u0_n112, 
       u1_u7_u0_n113, u1_u7_u0_n114, u1_u7_u0_n115, u1_u7_u0_n116, u1_u7_u0_n117, u1_u7_u0_n118, u1_u7_u0_n119, u1_u7_u0_n120, u1_u7_u0_n121, 
       u1_u7_u0_n122, u1_u7_u0_n123, u1_u7_u0_n124, u1_u7_u0_n125, u1_u7_u0_n126, u1_u7_u0_n127, u1_u7_u0_n128, u1_u7_u0_n129, u1_u7_u0_n130, 
       u1_u7_u0_n131, u1_u7_u0_n132, u1_u7_u0_n133, u1_u7_u0_n134, u1_u7_u0_n135, u1_u7_u0_n136, u1_u7_u0_n137, u1_u7_u0_n138, u1_u7_u0_n139, 
       u1_u7_u0_n140, u1_u7_u0_n141, u1_u7_u0_n142, u1_u7_u0_n143, u1_u7_u0_n144, u1_u7_u0_n145, u1_u7_u0_n146, u1_u7_u0_n147, u1_u7_u0_n148, 
       u1_u7_u0_n149, u1_u7_u0_n150, u1_u7_u0_n151, u1_u7_u0_n152, u1_u7_u0_n153, u1_u7_u0_n154, u1_u7_u0_n155, u1_u7_u0_n156, u1_u7_u0_n157, 
       u1_u7_u0_n158, u1_u7_u0_n159, u1_u7_u0_n160, u1_u7_u0_n161, u1_u7_u0_n162, u1_u7_u0_n163, u1_u7_u0_n164, u1_u7_u0_n165, u1_u7_u0_n166, 
       u1_u7_u0_n167, u1_u7_u0_n168, u1_u7_u0_n169, u1_u7_u0_n170, u1_u7_u0_n171, u1_u7_u0_n172, u1_u7_u0_n173, u1_u7_u0_n174, u1_u7_u0_n88, 
       u1_u7_u0_n89, u1_u7_u0_n90, u1_u7_u0_n91, u1_u7_u0_n92, u1_u7_u0_n93, u1_u7_u0_n94, u1_u7_u0_n95, u1_u7_u0_n96, u1_u7_u0_n97, 
       u1_u7_u0_n98, u1_u7_u0_n99, u1_u7_u1_n100, u1_u7_u1_n101, u1_u7_u1_n102, u1_u7_u1_n103, u1_u7_u1_n104, u1_u7_u1_n105, u1_u7_u1_n106, 
       u1_u7_u1_n107, u1_u7_u1_n108, u1_u7_u1_n109, u1_u7_u1_n110, u1_u7_u1_n111, u1_u7_u1_n112, u1_u7_u1_n113, u1_u7_u1_n114, u1_u7_u1_n115, 
       u1_u7_u1_n116, u1_u7_u1_n117, u1_u7_u1_n118, u1_u7_u1_n119, u1_u7_u1_n120, u1_u7_u1_n121, u1_u7_u1_n122, u1_u7_u1_n123, u1_u7_u1_n124, 
       u1_u7_u1_n125, u1_u7_u1_n126, u1_u7_u1_n127, u1_u7_u1_n128, u1_u7_u1_n129, u1_u7_u1_n130, u1_u7_u1_n131, u1_u7_u1_n132, u1_u7_u1_n133, 
       u1_u7_u1_n134, u1_u7_u1_n135, u1_u7_u1_n136, u1_u7_u1_n137, u1_u7_u1_n138, u1_u7_u1_n139, u1_u7_u1_n140, u1_u7_u1_n141, u1_u7_u1_n142, 
       u1_u7_u1_n143, u1_u7_u1_n144, u1_u7_u1_n145, u1_u7_u1_n146, u1_u7_u1_n147, u1_u7_u1_n148, u1_u7_u1_n149, u1_u7_u1_n150, u1_u7_u1_n151, 
       u1_u7_u1_n152, u1_u7_u1_n153, u1_u7_u1_n154, u1_u7_u1_n155, u1_u7_u1_n156, u1_u7_u1_n157, u1_u7_u1_n158, u1_u7_u1_n159, u1_u7_u1_n160, 
       u1_u7_u1_n161, u1_u7_u1_n162, u1_u7_u1_n163, u1_u7_u1_n164, u1_u7_u1_n165, u1_u7_u1_n166, u1_u7_u1_n167, u1_u7_u1_n168, u1_u7_u1_n169, 
       u1_u7_u1_n170, u1_u7_u1_n171, u1_u7_u1_n172, u1_u7_u1_n173, u1_u7_u1_n174, u1_u7_u1_n175, u1_u7_u1_n176, u1_u7_u1_n177, u1_u7_u1_n178, 
       u1_u7_u1_n179, u1_u7_u1_n180, u1_u7_u1_n181, u1_u7_u1_n182, u1_u7_u1_n183, u1_u7_u1_n184, u1_u7_u1_n185, u1_u7_u1_n186, u1_u7_u1_n187, 
       u1_u7_u1_n188, u1_u7_u1_n95, u1_u7_u1_n96, u1_u7_u1_n97, u1_u7_u1_n98, u1_u7_u1_n99, u1_u7_u2_n100, u1_u7_u2_n101, u1_u7_u2_n102, 
       u1_u7_u2_n103, u1_u7_u2_n104, u1_u7_u2_n105, u1_u7_u2_n106, u1_u7_u2_n107, u1_u7_u2_n108, u1_u7_u2_n109, u1_u7_u2_n110, u1_u7_u2_n111, 
       u1_u7_u2_n112, u1_u7_u2_n113, u1_u7_u2_n114, u1_u7_u2_n115, u1_u7_u2_n116, u1_u7_u2_n117, u1_u7_u2_n118, u1_u7_u2_n119, u1_u7_u2_n120, 
       u1_u7_u2_n121, u1_u7_u2_n122, u1_u7_u2_n123, u1_u7_u2_n124, u1_u7_u2_n125, u1_u7_u2_n126, u1_u7_u2_n127, u1_u7_u2_n128, u1_u7_u2_n129, 
       u1_u7_u2_n130, u1_u7_u2_n131, u1_u7_u2_n132, u1_u7_u2_n133, u1_u7_u2_n134, u1_u7_u2_n135, u1_u7_u2_n136, u1_u7_u2_n137, u1_u7_u2_n138, 
       u1_u7_u2_n139, u1_u7_u2_n140, u1_u7_u2_n141, u1_u7_u2_n142, u1_u7_u2_n143, u1_u7_u2_n144, u1_u7_u2_n145, u1_u7_u2_n146, u1_u7_u2_n147, 
       u1_u7_u2_n148, u1_u7_u2_n149, u1_u7_u2_n150, u1_u7_u2_n151, u1_u7_u2_n152, u1_u7_u2_n153, u1_u7_u2_n154, u1_u7_u2_n155, u1_u7_u2_n156, 
       u1_u7_u2_n157, u1_u7_u2_n158, u1_u7_u2_n159, u1_u7_u2_n160, u1_u7_u2_n161, u1_u7_u2_n162, u1_u7_u2_n163, u1_u7_u2_n164, u1_u7_u2_n165, 
       u1_u7_u2_n166, u1_u7_u2_n167, u1_u7_u2_n168, u1_u7_u2_n169, u1_u7_u2_n170, u1_u7_u2_n171, u1_u7_u2_n172, u1_u7_u2_n173, u1_u7_u2_n174, 
       u1_u7_u2_n175, u1_u7_u2_n176, u1_u7_u2_n177, u1_u7_u2_n178, u1_u7_u2_n179, u1_u7_u2_n180, u1_u7_u2_n181, u1_u7_u2_n182, u1_u7_u2_n183, 
       u1_u7_u2_n184, u1_u7_u2_n185, u1_u7_u2_n186, u1_u7_u2_n187, u1_u7_u2_n188, u1_u7_u2_n95, u1_u7_u2_n96, u1_u7_u2_n97, u1_u7_u2_n98, 
       u1_u7_u2_n99, u1_u8_X_43, u1_u8_X_44, u1_u8_X_45, u1_u8_X_46, u1_u8_X_47, u1_u8_X_48, u1_u8_u7_n100, u1_u8_u7_n101, 
       u1_u8_u7_n102, u1_u8_u7_n103, u1_u8_u7_n104, u1_u8_u7_n105, u1_u8_u7_n106, u1_u8_u7_n107, u1_u8_u7_n108, u1_u8_u7_n109, u1_u8_u7_n110, 
       u1_u8_u7_n111, u1_u8_u7_n112, u1_u8_u7_n113, u1_u8_u7_n114, u1_u8_u7_n115, u1_u8_u7_n116, u1_u8_u7_n117, u1_u8_u7_n118, u1_u8_u7_n119, 
       u1_u8_u7_n120, u1_u8_u7_n121, u1_u8_u7_n122, u1_u8_u7_n123, u1_u8_u7_n124, u1_u8_u7_n125, u1_u8_u7_n126, u1_u8_u7_n127, u1_u8_u7_n128, 
       u1_u8_u7_n129, u1_u8_u7_n130, u1_u8_u7_n131, u1_u8_u7_n132, u1_u8_u7_n133, u1_u8_u7_n134, u1_u8_u7_n135, u1_u8_u7_n136, u1_u8_u7_n137, 
       u1_u8_u7_n138, u1_u8_u7_n139, u1_u8_u7_n140, u1_u8_u7_n141, u1_u8_u7_n142, u1_u8_u7_n143, u1_u8_u7_n144, u1_u8_u7_n145, u1_u8_u7_n146, 
       u1_u8_u7_n147, u1_u8_u7_n148, u1_u8_u7_n149, u1_u8_u7_n150, u1_u8_u7_n151, u1_u8_u7_n152, u1_u8_u7_n153, u1_u8_u7_n154, u1_u8_u7_n155, 
       u1_u8_u7_n156, u1_u8_u7_n157, u1_u8_u7_n158, u1_u8_u7_n159, u1_u8_u7_n160, u1_u8_u7_n161, u1_u8_u7_n162, u1_u8_u7_n163, u1_u8_u7_n164, 
       u1_u8_u7_n165, u1_u8_u7_n166, u1_u8_u7_n167, u1_u8_u7_n168, u1_u8_u7_n169, u1_u8_u7_n170, u1_u8_u7_n171, u1_u8_u7_n172, u1_u8_u7_n173, 
       u1_u8_u7_n174, u1_u8_u7_n175, u1_u8_u7_n176, u1_u8_u7_n177, u1_u8_u7_n178, u1_u8_u7_n179, u1_u8_u7_n180, u1_u8_u7_n91, u1_u8_u7_n92, 
       u1_u8_u7_n93, u1_u8_u7_n94, u1_u8_u7_n95, u1_u8_u7_n96, u1_u8_u7_n97, u1_u8_u7_n98, u1_u8_u7_n99, u1_uk_n1063, u1_uk_n1064, 
       u1_uk_n1075, u1_uk_n1076, u1_uk_n1083, u1_uk_n1084, u1_uk_n1105, u1_uk_n1106, u1_uk_n1107, u1_uk_n1122, u1_uk_n1123, 
       u1_uk_n1124, u1_uk_n1126, u1_uk_n1127, u1_uk_n1128, u1_uk_n1129, u1_uk_n1130, u1_uk_n1131, u1_uk_n1132, u1_uk_n1135, 
       u1_uk_n1140, u1_uk_n1146, u1_uk_n1168, u1_uk_n1169, u1_uk_n1170, u1_uk_n456, u1_uk_n460, u1_uk_n467, u1_uk_n515, 
       u1_uk_n601, u1_uk_n656, u1_uk_n662, u1_uk_n964, u1_uk_n965, u1_uk_n966, u1_uk_n967, u1_uk_n968, u1_uk_n969, 
       u1_uk_n970, u1_uk_n976, u1_uk_n977, u1_uk_n984, u1_uk_n985, u1_uk_n987, u1_uk_n988, u1_uk_n989, u1_uk_n990, 
       u1_uk_n991, u1_uk_n992, u1_uk_n993, u1_uk_n994, u2_K2_25, u2_K2_26, u2_K2_27, u2_K2_28, u2_K2_29, 
       u2_K2_30, u2_out1_14, u2_out1_25, u2_out1_3, u2_out1_8, u2_u1_X_25, u2_u1_X_26, u2_u1_X_27, u2_u1_X_28, 
       u2_u1_X_29, u2_u1_X_30, u2_u1_u4_n100, u2_u1_u4_n101, u2_u1_u4_n102, u2_u1_u4_n103, u2_u1_u4_n104, u2_u1_u4_n105, u2_u1_u4_n106, 
       u2_u1_u4_n107, u2_u1_u4_n108, u2_u1_u4_n109, u2_u1_u4_n110, u2_u1_u4_n111, u2_u1_u4_n112, u2_u1_u4_n113, u2_u1_u4_n114, u2_u1_u4_n115, 
       u2_u1_u4_n116, u2_u1_u4_n117, u2_u1_u4_n118, u2_u1_u4_n119, u2_u1_u4_n120, u2_u1_u4_n121, u2_u1_u4_n122, u2_u1_u4_n123, u2_u1_u4_n124, 
       u2_u1_u4_n125, u2_u1_u4_n126, u2_u1_u4_n127, u2_u1_u4_n128, u2_u1_u4_n129, u2_u1_u4_n130, u2_u1_u4_n131, u2_u1_u4_n132, u2_u1_u4_n133, 
       u2_u1_u4_n134, u2_u1_u4_n135, u2_u1_u4_n136, u2_u1_u4_n137, u2_u1_u4_n138, u2_u1_u4_n139, u2_u1_u4_n140, u2_u1_u4_n141, u2_u1_u4_n142, 
       u2_u1_u4_n143, u2_u1_u4_n144, u2_u1_u4_n145, u2_u1_u4_n146, u2_u1_u4_n147, u2_u1_u4_n148, u2_u1_u4_n149, u2_u1_u4_n150, u2_u1_u4_n151, 
       u2_u1_u4_n152, u2_u1_u4_n153, u2_u1_u4_n154, u2_u1_u4_n155, u2_u1_u4_n156, u2_u1_u4_n157, u2_u1_u4_n158, u2_u1_u4_n159, u2_u1_u4_n160, 
       u2_u1_u4_n161, u2_u1_u4_n162, u2_u1_u4_n163, u2_u1_u4_n164, u2_u1_u4_n165, u2_u1_u4_n166, u2_u1_u4_n167, u2_u1_u4_n168, u2_u1_u4_n169, 
       u2_u1_u4_n170, u2_u1_u4_n171, u2_u1_u4_n172, u2_u1_u4_n173, u2_u1_u4_n174, u2_u1_u4_n175, u2_u1_u4_n176, u2_u1_u4_n177, u2_u1_u4_n178, 
       u2_u1_u4_n179, u2_u1_u4_n180, u2_u1_u4_n181, u2_u1_u4_n182, u2_u1_u4_n183, u2_u1_u4_n184, u2_u1_u4_n185, u2_u1_u4_n186, u2_u1_u4_n94, 
       u2_u1_u4_n95, u2_u1_u4_n96, u2_u1_u4_n97, u2_u1_u4_n98, u2_u1_u4_n99,  u2_uk_n998;
  XOR2_X1 u0_U10 (.B( u0_L1_29 ) , .Z( u0_N92 ) , .A( u0_out2_29 ) );
  XOR2_X1 u0_U15 (.B( u0_L1_25 ) , .Z( u0_N88 ) , .A( u0_out2_25 ) );
  XOR2_X1 u0_U192 (.B( u0_L0_5 ) , .Z( u0_N36 ) , .A( u0_out1_5 ) );
  XOR2_X1 u0_U202 (.B( u0_L9_31 ) , .Z( u0_N350 ) , .A( u0_out10_31 ) );
  XOR2_X1 u0_U21 (.B( u0_L1_19 ) , .Z( u0_N82 ) , .A( u0_out2_19 ) );
  XOR2_X1 u0_U211 (.B( u0_L9_23 ) , .Z( u0_N342 ) , .A( u0_out10_23 ) );
  XOR2_X1 u0_U218 (.B( u0_L9_17 ) , .Z( u0_N336 ) , .A( u0_out10_17 ) );
  XOR2_X1 u0_U227 (.B( u0_L9_9 ) , .Z( u0_N328 ) , .A( u0_out10_9 ) );
  XOR2_X1 u0_U27 (.B( u0_L1_14 ) , .Z( u0_N77 ) , .A( u0_out2_14 ) );
  XOR2_X1 u0_U30 (.B( u0_L1_11 ) , .Z( u0_N74 ) , .A( u0_out2_11 ) );
  XOR2_X1 u0_U33 (.B( u0_L1_8 ) , .Z( u0_N71 ) , .A( u0_out2_8 ) );
  XOR2_X1 u0_U38 (.B( u0_L1_4 ) , .Z( u0_N67 ) , .A( u0_out2_4 ) );
  XOR2_X1 u0_U39 (.B( u0_L1_3 ) , .Z( u0_N66 ) , .A( u0_out2_3 ) );
  XOR2_X1 u0_U48 (.B( u0_L0_27 ) , .Z( u0_N58 ) , .A( u0_out1_27 ) );
  XOR2_X1 u0_U54 (.B( u0_L0_21 ) , .Z( u0_N52 ) , .A( u0_out1_21 ) );
  XOR2_X1 u0_U66 (.B( u0_L13_26 ) , .Z( u0_N473 ) , .A( u0_out14_26 ) );
  XOR2_X1 u0_U73 (.B( u0_L13_20 ) , .Z( u0_N467 ) , .A( u0_out14_20 ) );
  XOR2_X1 u0_U81 (.B( u0_L0_15 ) , .Z( u0_N46 ) , .A( u0_out1_15 ) );
  XOR2_X1 u0_U84 (.B( u0_L13_10 ) , .Z( u0_N457 ) , .A( u0_out14_10 ) );
  XOR2_X1 u0_U94 (.B( u0_L13_1 ) , .Z( u0_N448 ) , .A( u0_out14_1 ) );
  XOR2_X1 u0_u10_U16 (.B( u0_K11_3 ) , .A( u0_R9_2 ) , .Z( u0_u10_X_3 ) );
  XOR2_X1 u0_u10_U27 (.B( u0_K11_2 ) , .A( u0_R9_1 ) , .Z( u0_u10_X_2 ) );
  XOR2_X1 u0_u10_U38 (.B( u0_K11_1 ) , .A( u0_R9_32 ) , .Z( u0_u10_X_1 ) );
  XOR2_X1 u0_u10_U4 (.B( u0_K11_6 ) , .A( u0_R9_5 ) , .Z( u0_u10_X_6 ) );
  XOR2_X1 u0_u10_U5 (.B( u0_K11_5 ) , .A( u0_R9_4 ) , .Z( u0_u10_X_5 ) );
  XOR2_X1 u0_u10_U6 (.B( u0_K11_4 ) , .A( u0_R9_3 ) , .Z( u0_u10_X_4 ) );
  AND3_X1 u0_u10_u0_U10 (.A2( u0_u10_u0_n112 ) , .ZN( u0_u10_u0_n127 ) , .A3( u0_u10_u0_n130 ) , .A1( u0_u10_u0_n148 ) );
  NAND2_X1 u0_u10_u0_U11 (.ZN( u0_u10_u0_n113 ) , .A1( u0_u10_u0_n139 ) , .A2( u0_u10_u0_n149 ) );
  AND2_X1 u0_u10_u0_U12 (.ZN( u0_u10_u0_n107 ) , .A1( u0_u10_u0_n130 ) , .A2( u0_u10_u0_n140 ) );
  AND2_X1 u0_u10_u0_U13 (.A2( u0_u10_u0_n129 ) , .A1( u0_u10_u0_n130 ) , .ZN( u0_u10_u0_n151 ) );
  AND2_X1 u0_u10_u0_U14 (.A1( u0_u10_u0_n108 ) , .A2( u0_u10_u0_n125 ) , .ZN( u0_u10_u0_n145 ) );
  INV_X1 u0_u10_u0_U15 (.A( u0_u10_u0_n143 ) , .ZN( u0_u10_u0_n173 ) );
  NOR2_X1 u0_u10_u0_U16 (.A2( u0_u10_u0_n136 ) , .ZN( u0_u10_u0_n147 ) , .A1( u0_u10_u0_n160 ) );
  NOR2_X1 u0_u10_u0_U17 (.A1( u0_u10_u0_n163 ) , .A2( u0_u10_u0_n164 ) , .ZN( u0_u10_u0_n95 ) );
  AOI21_X1 u0_u10_u0_U18 (.B1( u0_u10_u0_n103 ) , .ZN( u0_u10_u0_n132 ) , .A( u0_u10_u0_n165 ) , .B2( u0_u10_u0_n93 ) );
  INV_X1 u0_u10_u0_U19 (.A( u0_u10_u0_n142 ) , .ZN( u0_u10_u0_n165 ) );
  OAI221_X1 u0_u10_u0_U20 (.C1( u0_u10_u0_n121 ) , .ZN( u0_u10_u0_n122 ) , .B2( u0_u10_u0_n127 ) , .A( u0_u10_u0_n143 ) , .B1( u0_u10_u0_n144 ) , .C2( u0_u10_u0_n147 ) );
  OAI22_X1 u0_u10_u0_U21 (.B1( u0_u10_u0_n125 ) , .ZN( u0_u10_u0_n126 ) , .A1( u0_u10_u0_n138 ) , .A2( u0_u10_u0_n146 ) , .B2( u0_u10_u0_n147 ) );
  OAI22_X1 u0_u10_u0_U22 (.B1( u0_u10_u0_n131 ) , .A1( u0_u10_u0_n144 ) , .B2( u0_u10_u0_n147 ) , .A2( u0_u10_u0_n90 ) , .ZN( u0_u10_u0_n91 ) );
  AND3_X1 u0_u10_u0_U23 (.A3( u0_u10_u0_n121 ) , .A2( u0_u10_u0_n125 ) , .A1( u0_u10_u0_n148 ) , .ZN( u0_u10_u0_n90 ) );
  INV_X1 u0_u10_u0_U24 (.A( u0_u10_u0_n136 ) , .ZN( u0_u10_u0_n161 ) );
  NOR2_X1 u0_u10_u0_U25 (.A1( u0_u10_u0_n120 ) , .ZN( u0_u10_u0_n143 ) , .A2( u0_u10_u0_n167 ) );
  OAI221_X1 u0_u10_u0_U26 (.C1( u0_u10_u0_n112 ) , .ZN( u0_u10_u0_n120 ) , .B1( u0_u10_u0_n138 ) , .B2( u0_u10_u0_n141 ) , .C2( u0_u10_u0_n147 ) , .A( u0_u10_u0_n172 ) );
  AOI22_X1 u0_u10_u0_U27 (.B2( u0_u10_u0_n109 ) , .A2( u0_u10_u0_n110 ) , .ZN( u0_u10_u0_n111 ) , .B1( u0_u10_u0_n118 ) , .A1( u0_u10_u0_n160 ) );
  INV_X1 u0_u10_u0_U28 (.A( u0_u10_u0_n118 ) , .ZN( u0_u10_u0_n158 ) );
  AOI21_X1 u0_u10_u0_U29 (.B1( u0_u10_u0_n132 ) , .ZN( u0_u10_u0_n133 ) , .A( u0_u10_u0_n144 ) , .B2( u0_u10_u0_n166 ) );
  INV_X1 u0_u10_u0_U3 (.A( u0_u10_u0_n113 ) , .ZN( u0_u10_u0_n166 ) );
  AOI21_X1 u0_u10_u0_U30 (.ZN( u0_u10_u0_n104 ) , .B1( u0_u10_u0_n107 ) , .B2( u0_u10_u0_n141 ) , .A( u0_u10_u0_n144 ) );
  AOI21_X1 u0_u10_u0_U31 (.B1( u0_u10_u0_n127 ) , .B2( u0_u10_u0_n129 ) , .A( u0_u10_u0_n138 ) , .ZN( u0_u10_u0_n96 ) );
  AOI21_X1 u0_u10_u0_U32 (.ZN( u0_u10_u0_n116 ) , .B2( u0_u10_u0_n142 ) , .A( u0_u10_u0_n144 ) , .B1( u0_u10_u0_n166 ) );
  NAND2_X1 u0_u10_u0_U33 (.A1( u0_u10_u0_n100 ) , .A2( u0_u10_u0_n103 ) , .ZN( u0_u10_u0_n125 ) );
  NAND2_X1 u0_u10_u0_U34 (.A2( u0_u10_u0_n103 ) , .ZN( u0_u10_u0_n140 ) , .A1( u0_u10_u0_n94 ) );
  NAND2_X1 u0_u10_u0_U35 (.A1( u0_u10_u0_n101 ) , .A2( u0_u10_u0_n102 ) , .ZN( u0_u10_u0_n150 ) );
  INV_X1 u0_u10_u0_U36 (.A( u0_u10_u0_n138 ) , .ZN( u0_u10_u0_n160 ) );
  NAND2_X1 u0_u10_u0_U37 (.ZN( u0_u10_u0_n142 ) , .A1( u0_u10_u0_n94 ) , .A2( u0_u10_u0_n95 ) );
  NAND2_X1 u0_u10_u0_U38 (.A1( u0_u10_u0_n102 ) , .ZN( u0_u10_u0_n128 ) , .A2( u0_u10_u0_n95 ) );
  NAND2_X1 u0_u10_u0_U39 (.A2( u0_u10_u0_n102 ) , .A1( u0_u10_u0_n103 ) , .ZN( u0_u10_u0_n149 ) );
  AOI21_X1 u0_u10_u0_U4 (.B2( u0_u10_u0_n131 ) , .ZN( u0_u10_u0_n134 ) , .B1( u0_u10_u0_n151 ) , .A( u0_u10_u0_n158 ) );
  NAND2_X1 u0_u10_u0_U40 (.A1( u0_u10_u0_n100 ) , .ZN( u0_u10_u0_n129 ) , .A2( u0_u10_u0_n95 ) );
  NAND2_X1 u0_u10_u0_U41 (.A2( u0_u10_u0_n100 ) , .A1( u0_u10_u0_n101 ) , .ZN( u0_u10_u0_n139 ) );
  NAND2_X1 u0_u10_u0_U42 (.A2( u0_u10_u0_n100 ) , .ZN( u0_u10_u0_n131 ) , .A1( u0_u10_u0_n92 ) );
  NAND2_X1 u0_u10_u0_U43 (.ZN( u0_u10_u0_n108 ) , .A1( u0_u10_u0_n92 ) , .A2( u0_u10_u0_n94 ) );
  NAND2_X1 u0_u10_u0_U44 (.ZN( u0_u10_u0_n148 ) , .A1( u0_u10_u0_n93 ) , .A2( u0_u10_u0_n95 ) );
  NAND2_X1 u0_u10_u0_U45 (.A2( u0_u10_u0_n102 ) , .ZN( u0_u10_u0_n114 ) , .A1( u0_u10_u0_n92 ) );
  NAND2_X1 u0_u10_u0_U46 (.A1( u0_u10_u0_n101 ) , .ZN( u0_u10_u0_n130 ) , .A2( u0_u10_u0_n94 ) );
  NAND2_X1 u0_u10_u0_U47 (.A2( u0_u10_u0_n101 ) , .ZN( u0_u10_u0_n121 ) , .A1( u0_u10_u0_n93 ) );
  INV_X1 u0_u10_u0_U48 (.ZN( u0_u10_u0_n172 ) , .A( u0_u10_u0_n88 ) );
  OAI222_X1 u0_u10_u0_U49 (.C1( u0_u10_u0_n108 ) , .A1( u0_u10_u0_n125 ) , .B2( u0_u10_u0_n128 ) , .B1( u0_u10_u0_n144 ) , .A2( u0_u10_u0_n158 ) , .C2( u0_u10_u0_n161 ) , .ZN( u0_u10_u0_n88 ) );
  NOR2_X1 u0_u10_u0_U5 (.A1( u0_u10_u0_n108 ) , .ZN( u0_u10_u0_n123 ) , .A2( u0_u10_u0_n158 ) );
  NAND2_X1 u0_u10_u0_U50 (.ZN( u0_u10_u0_n112 ) , .A2( u0_u10_u0_n92 ) , .A1( u0_u10_u0_n93 ) );
  OR3_X1 u0_u10_u0_U51 (.A3( u0_u10_u0_n152 ) , .A2( u0_u10_u0_n153 ) , .A1( u0_u10_u0_n154 ) , .ZN( u0_u10_u0_n155 ) );
  AOI21_X1 u0_u10_u0_U52 (.A( u0_u10_u0_n144 ) , .B2( u0_u10_u0_n145 ) , .B1( u0_u10_u0_n146 ) , .ZN( u0_u10_u0_n154 ) );
  AOI21_X1 u0_u10_u0_U53 (.B2( u0_u10_u0_n150 ) , .B1( u0_u10_u0_n151 ) , .ZN( u0_u10_u0_n152 ) , .A( u0_u10_u0_n158 ) );
  AOI21_X1 u0_u10_u0_U54 (.A( u0_u10_u0_n147 ) , .B2( u0_u10_u0_n148 ) , .B1( u0_u10_u0_n149 ) , .ZN( u0_u10_u0_n153 ) );
  INV_X1 u0_u10_u0_U55 (.ZN( u0_u10_u0_n171 ) , .A( u0_u10_u0_n99 ) );
  OAI211_X1 u0_u10_u0_U56 (.C2( u0_u10_u0_n140 ) , .C1( u0_u10_u0_n161 ) , .A( u0_u10_u0_n169 ) , .B( u0_u10_u0_n98 ) , .ZN( u0_u10_u0_n99 ) );
  INV_X1 u0_u10_u0_U57 (.ZN( u0_u10_u0_n169 ) , .A( u0_u10_u0_n91 ) );
  AOI211_X1 u0_u10_u0_U58 (.C1( u0_u10_u0_n118 ) , .A( u0_u10_u0_n123 ) , .B( u0_u10_u0_n96 ) , .C2( u0_u10_u0_n97 ) , .ZN( u0_u10_u0_n98 ) );
  NOR2_X1 u0_u10_u0_U59 (.A2( u0_u10_X_2 ) , .ZN( u0_u10_u0_n103 ) , .A1( u0_u10_u0_n164 ) );
  OAI21_X1 u0_u10_u0_U6 (.B1( u0_u10_u0_n150 ) , .B2( u0_u10_u0_n158 ) , .A( u0_u10_u0_n172 ) , .ZN( u0_u10_u0_n89 ) );
  NOR2_X1 u0_u10_u0_U60 (.A2( u0_u10_X_3 ) , .A1( u0_u10_X_6 ) , .ZN( u0_u10_u0_n94 ) );
  NOR2_X1 u0_u10_u0_U61 (.A2( u0_u10_X_6 ) , .ZN( u0_u10_u0_n100 ) , .A1( u0_u10_u0_n162 ) );
  NOR2_X1 u0_u10_u0_U62 (.A2( u0_u10_X_1 ) , .A1( u0_u10_X_2 ) , .ZN( u0_u10_u0_n92 ) );
  NOR2_X1 u0_u10_u0_U63 (.A2( u0_u10_X_1 ) , .ZN( u0_u10_u0_n101 ) , .A1( u0_u10_u0_n163 ) );
  NOR2_X1 u0_u10_u0_U64 (.A2( u0_u10_X_4 ) , .A1( u0_u10_X_5 ) , .ZN( u0_u10_u0_n118 ) );
  NAND2_X1 u0_u10_u0_U65 (.A2( u0_u10_X_4 ) , .A1( u0_u10_X_5 ) , .ZN( u0_u10_u0_n144 ) );
  NOR2_X1 u0_u10_u0_U66 (.A2( u0_u10_X_5 ) , .ZN( u0_u10_u0_n136 ) , .A1( u0_u10_u0_n159 ) );
  NAND2_X1 u0_u10_u0_U67 (.A1( u0_u10_X_5 ) , .ZN( u0_u10_u0_n138 ) , .A2( u0_u10_u0_n159 ) );
  AND2_X1 u0_u10_u0_U68 (.A2( u0_u10_X_3 ) , .A1( u0_u10_X_6 ) , .ZN( u0_u10_u0_n102 ) );
  AND2_X1 u0_u10_u0_U69 (.A1( u0_u10_X_6 ) , .A2( u0_u10_u0_n162 ) , .ZN( u0_u10_u0_n93 ) );
  AOI21_X1 u0_u10_u0_U7 (.B1( u0_u10_u0_n114 ) , .ZN( u0_u10_u0_n115 ) , .B2( u0_u10_u0_n129 ) , .A( u0_u10_u0_n161 ) );
  INV_X1 u0_u10_u0_U70 (.A( u0_u10_X_4 ) , .ZN( u0_u10_u0_n159 ) );
  INV_X1 u0_u10_u0_U71 (.A( u0_u10_X_1 ) , .ZN( u0_u10_u0_n164 ) );
  INV_X1 u0_u10_u0_U72 (.A( u0_u10_X_2 ) , .ZN( u0_u10_u0_n163 ) );
  INV_X1 u0_u10_u0_U73 (.A( u0_u10_X_3 ) , .ZN( u0_u10_u0_n162 ) );
  INV_X1 u0_u10_u0_U74 (.A( u0_u10_u0_n126 ) , .ZN( u0_u10_u0_n168 ) );
  AOI211_X1 u0_u10_u0_U75 (.B( u0_u10_u0_n133 ) , .A( u0_u10_u0_n134 ) , .C2( u0_u10_u0_n135 ) , .C1( u0_u10_u0_n136 ) , .ZN( u0_u10_u0_n137 ) );
  INV_X1 u0_u10_u0_U76 (.ZN( u0_u10_u0_n174 ) , .A( u0_u10_u0_n89 ) );
  AOI211_X1 u0_u10_u0_U77 (.B( u0_u10_u0_n104 ) , .A( u0_u10_u0_n105 ) , .ZN( u0_u10_u0_n106 ) , .C2( u0_u10_u0_n113 ) , .C1( u0_u10_u0_n160 ) );
  OR4_X1 u0_u10_u0_U78 (.ZN( u0_out10_31 ) , .A4( u0_u10_u0_n155 ) , .A2( u0_u10_u0_n156 ) , .A1( u0_u10_u0_n157 ) , .A3( u0_u10_u0_n173 ) );
  AOI21_X1 u0_u10_u0_U79 (.A( u0_u10_u0_n138 ) , .B2( u0_u10_u0_n139 ) , .B1( u0_u10_u0_n140 ) , .ZN( u0_u10_u0_n157 ) );
  AND2_X1 u0_u10_u0_U8 (.A1( u0_u10_u0_n114 ) , .A2( u0_u10_u0_n121 ) , .ZN( u0_u10_u0_n146 ) );
  AOI21_X1 u0_u10_u0_U80 (.B2( u0_u10_u0_n141 ) , .B1( u0_u10_u0_n142 ) , .ZN( u0_u10_u0_n156 ) , .A( u0_u10_u0_n161 ) );
  OR4_X1 u0_u10_u0_U81 (.ZN( u0_out10_17 ) , .A4( u0_u10_u0_n122 ) , .A2( u0_u10_u0_n123 ) , .A1( u0_u10_u0_n124 ) , .A3( u0_u10_u0_n170 ) );
  AOI21_X1 u0_u10_u0_U82 (.B2( u0_u10_u0_n107 ) , .ZN( u0_u10_u0_n124 ) , .B1( u0_u10_u0_n128 ) , .A( u0_u10_u0_n161 ) );
  INV_X1 u0_u10_u0_U83 (.A( u0_u10_u0_n111 ) , .ZN( u0_u10_u0_n170 ) );
  AOI211_X1 u0_u10_u0_U84 (.B( u0_u10_u0_n115 ) , .A( u0_u10_u0_n116 ) , .C2( u0_u10_u0_n117 ) , .C1( u0_u10_u0_n118 ) , .ZN( u0_u10_u0_n119 ) );
  INV_X1 u0_u10_u0_U85 (.A( u0_u10_u0_n119 ) , .ZN( u0_u10_u0_n167 ) );
  NAND2_X1 u0_u10_u0_U86 (.ZN( u0_u10_u0_n110 ) , .A2( u0_u10_u0_n132 ) , .A1( u0_u10_u0_n145 ) );
  OAI22_X1 u0_u10_u0_U87 (.ZN( u0_u10_u0_n105 ) , .A2( u0_u10_u0_n132 ) , .B1( u0_u10_u0_n146 ) , .A1( u0_u10_u0_n147 ) , .B2( u0_u10_u0_n161 ) );
  NAND3_X1 u0_u10_u0_U88 (.ZN( u0_out10_23 ) , .A3( u0_u10_u0_n137 ) , .A1( u0_u10_u0_n168 ) , .A2( u0_u10_u0_n171 ) );
  NAND3_X1 u0_u10_u0_U89 (.A3( u0_u10_u0_n127 ) , .A2( u0_u10_u0_n128 ) , .ZN( u0_u10_u0_n135 ) , .A1( u0_u10_u0_n150 ) );
  AND2_X1 u0_u10_u0_U9 (.A1( u0_u10_u0_n131 ) , .ZN( u0_u10_u0_n141 ) , .A2( u0_u10_u0_n150 ) );
  NAND3_X1 u0_u10_u0_U90 (.ZN( u0_u10_u0_n117 ) , .A3( u0_u10_u0_n132 ) , .A2( u0_u10_u0_n139 ) , .A1( u0_u10_u0_n148 ) );
  NAND3_X1 u0_u10_u0_U91 (.ZN( u0_u10_u0_n109 ) , .A2( u0_u10_u0_n114 ) , .A3( u0_u10_u0_n140 ) , .A1( u0_u10_u0_n149 ) );
  NAND3_X1 u0_u10_u0_U92 (.ZN( u0_out10_9 ) , .A3( u0_u10_u0_n106 ) , .A2( u0_u10_u0_n171 ) , .A1( u0_u10_u0_n174 ) );
  NAND3_X1 u0_u10_u0_U93 (.A2( u0_u10_u0_n128 ) , .A1( u0_u10_u0_n132 ) , .A3( u0_u10_u0_n146 ) , .ZN( u0_u10_u0_n97 ) );
  XOR2_X1 u0_u14_U33 (.B( u0_K15_24 ) , .A( u0_R13_17 ) , .Z( u0_u14_X_24 ) );
  XOR2_X1 u0_u14_U34 (.B( u0_K15_23 ) , .A( u0_R13_16 ) , .Z( u0_u14_X_23 ) );
  XOR2_X1 u0_u14_U35 (.B( u0_K15_22 ) , .A( u0_R13_15 ) , .Z( u0_u14_X_22 ) );
  XOR2_X1 u0_u14_U36 (.B( u0_K15_21 ) , .A( u0_R13_14 ) , .Z( u0_u14_X_21 ) );
  XOR2_X1 u0_u14_U37 (.B( u0_K15_20 ) , .A( u0_R13_13 ) , .Z( u0_u14_X_20 ) );
  XOR2_X1 u0_u14_U39 (.B( u0_K15_19 ) , .A( u0_R13_12 ) , .Z( u0_u14_X_19 ) );
  OAI22_X1 u0_u14_u3_U10 (.B1( u0_u14_u3_n113 ) , .A2( u0_u14_u3_n135 ) , .A1( u0_u14_u3_n150 ) , .B2( u0_u14_u3_n164 ) , .ZN( u0_u14_u3_n98 ) );
  OAI211_X1 u0_u14_u3_U11 (.B( u0_u14_u3_n106 ) , .ZN( u0_u14_u3_n119 ) , .C2( u0_u14_u3_n128 ) , .C1( u0_u14_u3_n167 ) , .A( u0_u14_u3_n181 ) );
  AOI221_X1 u0_u14_u3_U12 (.C1( u0_u14_u3_n105 ) , .ZN( u0_u14_u3_n106 ) , .A( u0_u14_u3_n131 ) , .B2( u0_u14_u3_n132 ) , .C2( u0_u14_u3_n133 ) , .B1( u0_u14_u3_n169 ) );
  INV_X1 u0_u14_u3_U13 (.ZN( u0_u14_u3_n181 ) , .A( u0_u14_u3_n98 ) );
  NAND2_X1 u0_u14_u3_U14 (.ZN( u0_u14_u3_n105 ) , .A2( u0_u14_u3_n130 ) , .A1( u0_u14_u3_n155 ) );
  AOI22_X1 u0_u14_u3_U15 (.B1( u0_u14_u3_n115 ) , .A2( u0_u14_u3_n116 ) , .ZN( u0_u14_u3_n123 ) , .B2( u0_u14_u3_n133 ) , .A1( u0_u14_u3_n169 ) );
  NAND2_X1 u0_u14_u3_U16 (.ZN( u0_u14_u3_n116 ) , .A2( u0_u14_u3_n151 ) , .A1( u0_u14_u3_n182 ) );
  NOR2_X1 u0_u14_u3_U17 (.ZN( u0_u14_u3_n126 ) , .A2( u0_u14_u3_n150 ) , .A1( u0_u14_u3_n164 ) );
  AOI21_X1 u0_u14_u3_U18 (.ZN( u0_u14_u3_n112 ) , .B2( u0_u14_u3_n146 ) , .B1( u0_u14_u3_n155 ) , .A( u0_u14_u3_n167 ) );
  NAND2_X1 u0_u14_u3_U19 (.A1( u0_u14_u3_n135 ) , .ZN( u0_u14_u3_n142 ) , .A2( u0_u14_u3_n164 ) );
  NAND2_X1 u0_u14_u3_U20 (.ZN( u0_u14_u3_n132 ) , .A2( u0_u14_u3_n152 ) , .A1( u0_u14_u3_n156 ) );
  AND2_X1 u0_u14_u3_U21 (.A2( u0_u14_u3_n113 ) , .A1( u0_u14_u3_n114 ) , .ZN( u0_u14_u3_n151 ) );
  INV_X1 u0_u14_u3_U22 (.A( u0_u14_u3_n133 ) , .ZN( u0_u14_u3_n165 ) );
  INV_X1 u0_u14_u3_U23 (.A( u0_u14_u3_n135 ) , .ZN( u0_u14_u3_n170 ) );
  NAND2_X1 u0_u14_u3_U24 (.A1( u0_u14_u3_n107 ) , .A2( u0_u14_u3_n108 ) , .ZN( u0_u14_u3_n140 ) );
  NAND2_X1 u0_u14_u3_U25 (.ZN( u0_u14_u3_n117 ) , .A1( u0_u14_u3_n124 ) , .A2( u0_u14_u3_n148 ) );
  NAND2_X1 u0_u14_u3_U26 (.ZN( u0_u14_u3_n143 ) , .A1( u0_u14_u3_n165 ) , .A2( u0_u14_u3_n167 ) );
  INV_X1 u0_u14_u3_U27 (.A( u0_u14_u3_n130 ) , .ZN( u0_u14_u3_n177 ) );
  INV_X1 u0_u14_u3_U28 (.A( u0_u14_u3_n128 ) , .ZN( u0_u14_u3_n176 ) );
  INV_X1 u0_u14_u3_U29 (.A( u0_u14_u3_n155 ) , .ZN( u0_u14_u3_n174 ) );
  INV_X1 u0_u14_u3_U3 (.A( u0_u14_u3_n129 ) , .ZN( u0_u14_u3_n183 ) );
  INV_X1 u0_u14_u3_U30 (.A( u0_u14_u3_n139 ) , .ZN( u0_u14_u3_n185 ) );
  NOR2_X1 u0_u14_u3_U31 (.ZN( u0_u14_u3_n135 ) , .A2( u0_u14_u3_n141 ) , .A1( u0_u14_u3_n169 ) );
  OAI222_X1 u0_u14_u3_U32 (.C2( u0_u14_u3_n107 ) , .A2( u0_u14_u3_n108 ) , .B1( u0_u14_u3_n135 ) , .ZN( u0_u14_u3_n138 ) , .B2( u0_u14_u3_n146 ) , .C1( u0_u14_u3_n154 ) , .A1( u0_u14_u3_n164 ) );
  NOR4_X1 u0_u14_u3_U33 (.A4( u0_u14_u3_n157 ) , .A3( u0_u14_u3_n158 ) , .A2( u0_u14_u3_n159 ) , .A1( u0_u14_u3_n160 ) , .ZN( u0_u14_u3_n161 ) );
  AOI21_X1 u0_u14_u3_U34 (.B2( u0_u14_u3_n152 ) , .B1( u0_u14_u3_n153 ) , .ZN( u0_u14_u3_n158 ) , .A( u0_u14_u3_n164 ) );
  AOI21_X1 u0_u14_u3_U35 (.A( u0_u14_u3_n154 ) , .B2( u0_u14_u3_n155 ) , .B1( u0_u14_u3_n156 ) , .ZN( u0_u14_u3_n157 ) );
  AOI21_X1 u0_u14_u3_U36 (.A( u0_u14_u3_n149 ) , .B2( u0_u14_u3_n150 ) , .B1( u0_u14_u3_n151 ) , .ZN( u0_u14_u3_n159 ) );
  AOI211_X1 u0_u14_u3_U37 (.ZN( u0_u14_u3_n109 ) , .A( u0_u14_u3_n119 ) , .C2( u0_u14_u3_n129 ) , .B( u0_u14_u3_n138 ) , .C1( u0_u14_u3_n141 ) );
  AOI211_X1 u0_u14_u3_U38 (.B( u0_u14_u3_n119 ) , .A( u0_u14_u3_n120 ) , .C2( u0_u14_u3_n121 ) , .ZN( u0_u14_u3_n122 ) , .C1( u0_u14_u3_n179 ) );
  INV_X1 u0_u14_u3_U39 (.A( u0_u14_u3_n156 ) , .ZN( u0_u14_u3_n179 ) );
  INV_X1 u0_u14_u3_U4 (.A( u0_u14_u3_n140 ) , .ZN( u0_u14_u3_n182 ) );
  OAI22_X1 u0_u14_u3_U40 (.B1( u0_u14_u3_n118 ) , .ZN( u0_u14_u3_n120 ) , .A1( u0_u14_u3_n135 ) , .B2( u0_u14_u3_n154 ) , .A2( u0_u14_u3_n178 ) );
  AND3_X1 u0_u14_u3_U41 (.ZN( u0_u14_u3_n118 ) , .A2( u0_u14_u3_n124 ) , .A1( u0_u14_u3_n144 ) , .A3( u0_u14_u3_n152 ) );
  INV_X1 u0_u14_u3_U42 (.A( u0_u14_u3_n121 ) , .ZN( u0_u14_u3_n164 ) );
  NAND2_X1 u0_u14_u3_U43 (.ZN( u0_u14_u3_n133 ) , .A1( u0_u14_u3_n154 ) , .A2( u0_u14_u3_n164 ) );
  OAI211_X1 u0_u14_u3_U44 (.B( u0_u14_u3_n127 ) , .ZN( u0_u14_u3_n139 ) , .C1( u0_u14_u3_n150 ) , .C2( u0_u14_u3_n154 ) , .A( u0_u14_u3_n184 ) );
  INV_X1 u0_u14_u3_U45 (.A( u0_u14_u3_n125 ) , .ZN( u0_u14_u3_n184 ) );
  AOI221_X1 u0_u14_u3_U46 (.A( u0_u14_u3_n126 ) , .ZN( u0_u14_u3_n127 ) , .C2( u0_u14_u3_n132 ) , .C1( u0_u14_u3_n169 ) , .B2( u0_u14_u3_n170 ) , .B1( u0_u14_u3_n174 ) );
  OAI22_X1 u0_u14_u3_U47 (.A1( u0_u14_u3_n124 ) , .ZN( u0_u14_u3_n125 ) , .B2( u0_u14_u3_n145 ) , .A2( u0_u14_u3_n165 ) , .B1( u0_u14_u3_n167 ) );
  NOR2_X1 u0_u14_u3_U48 (.A1( u0_u14_u3_n113 ) , .ZN( u0_u14_u3_n131 ) , .A2( u0_u14_u3_n154 ) );
  NAND2_X1 u0_u14_u3_U49 (.A1( u0_u14_u3_n103 ) , .ZN( u0_u14_u3_n150 ) , .A2( u0_u14_u3_n99 ) );
  INV_X1 u0_u14_u3_U5 (.A( u0_u14_u3_n117 ) , .ZN( u0_u14_u3_n178 ) );
  NAND2_X1 u0_u14_u3_U50 (.A2( u0_u14_u3_n102 ) , .ZN( u0_u14_u3_n155 ) , .A1( u0_u14_u3_n97 ) );
  INV_X1 u0_u14_u3_U51 (.A( u0_u14_u3_n141 ) , .ZN( u0_u14_u3_n167 ) );
  AOI21_X1 u0_u14_u3_U52 (.B2( u0_u14_u3_n114 ) , .B1( u0_u14_u3_n146 ) , .A( u0_u14_u3_n154 ) , .ZN( u0_u14_u3_n94 ) );
  AOI21_X1 u0_u14_u3_U53 (.ZN( u0_u14_u3_n110 ) , .B2( u0_u14_u3_n142 ) , .B1( u0_u14_u3_n186 ) , .A( u0_u14_u3_n95 ) );
  INV_X1 u0_u14_u3_U54 (.A( u0_u14_u3_n145 ) , .ZN( u0_u14_u3_n186 ) );
  AOI21_X1 u0_u14_u3_U55 (.B1( u0_u14_u3_n124 ) , .A( u0_u14_u3_n149 ) , .B2( u0_u14_u3_n155 ) , .ZN( u0_u14_u3_n95 ) );
  INV_X1 u0_u14_u3_U56 (.A( u0_u14_u3_n149 ) , .ZN( u0_u14_u3_n169 ) );
  NAND2_X1 u0_u14_u3_U57 (.ZN( u0_u14_u3_n124 ) , .A1( u0_u14_u3_n96 ) , .A2( u0_u14_u3_n97 ) );
  NAND2_X1 u0_u14_u3_U58 (.A2( u0_u14_u3_n100 ) , .ZN( u0_u14_u3_n146 ) , .A1( u0_u14_u3_n96 ) );
  NAND2_X1 u0_u14_u3_U59 (.A1( u0_u14_u3_n101 ) , .ZN( u0_u14_u3_n145 ) , .A2( u0_u14_u3_n99 ) );
  AOI221_X1 u0_u14_u3_U6 (.A( u0_u14_u3_n131 ) , .C2( u0_u14_u3_n132 ) , .C1( u0_u14_u3_n133 ) , .ZN( u0_u14_u3_n134 ) , .B1( u0_u14_u3_n143 ) , .B2( u0_u14_u3_n177 ) );
  NAND2_X1 u0_u14_u3_U60 (.A1( u0_u14_u3_n100 ) , .ZN( u0_u14_u3_n156 ) , .A2( u0_u14_u3_n99 ) );
  NAND2_X1 u0_u14_u3_U61 (.A2( u0_u14_u3_n101 ) , .A1( u0_u14_u3_n104 ) , .ZN( u0_u14_u3_n148 ) );
  NAND2_X1 u0_u14_u3_U62 (.A1( u0_u14_u3_n100 ) , .A2( u0_u14_u3_n102 ) , .ZN( u0_u14_u3_n128 ) );
  NAND2_X1 u0_u14_u3_U63 (.A2( u0_u14_u3_n101 ) , .A1( u0_u14_u3_n102 ) , .ZN( u0_u14_u3_n152 ) );
  NAND2_X1 u0_u14_u3_U64 (.A2( u0_u14_u3_n101 ) , .ZN( u0_u14_u3_n114 ) , .A1( u0_u14_u3_n96 ) );
  NAND2_X1 u0_u14_u3_U65 (.ZN( u0_u14_u3_n107 ) , .A1( u0_u14_u3_n97 ) , .A2( u0_u14_u3_n99 ) );
  NAND2_X1 u0_u14_u3_U66 (.A2( u0_u14_u3_n100 ) , .A1( u0_u14_u3_n104 ) , .ZN( u0_u14_u3_n113 ) );
  NAND2_X1 u0_u14_u3_U67 (.A1( u0_u14_u3_n104 ) , .ZN( u0_u14_u3_n153 ) , .A2( u0_u14_u3_n97 ) );
  NAND2_X1 u0_u14_u3_U68 (.A2( u0_u14_u3_n103 ) , .A1( u0_u14_u3_n104 ) , .ZN( u0_u14_u3_n130 ) );
  NAND2_X1 u0_u14_u3_U69 (.A2( u0_u14_u3_n103 ) , .ZN( u0_u14_u3_n144 ) , .A1( u0_u14_u3_n96 ) );
  OAI22_X1 u0_u14_u3_U7 (.B2( u0_u14_u3_n147 ) , .A2( u0_u14_u3_n148 ) , .ZN( u0_u14_u3_n160 ) , .B1( u0_u14_u3_n165 ) , .A1( u0_u14_u3_n168 ) );
  NAND2_X1 u0_u14_u3_U70 (.A1( u0_u14_u3_n102 ) , .A2( u0_u14_u3_n103 ) , .ZN( u0_u14_u3_n108 ) );
  NOR2_X1 u0_u14_u3_U71 (.A2( u0_u14_X_19 ) , .A1( u0_u14_X_20 ) , .ZN( u0_u14_u3_n99 ) );
  NOR2_X1 u0_u14_u3_U72 (.A2( u0_u14_X_21 ) , .A1( u0_u14_X_24 ) , .ZN( u0_u14_u3_n103 ) );
  NOR2_X1 u0_u14_u3_U73 (.A2( u0_u14_X_24 ) , .A1( u0_u14_u3_n171 ) , .ZN( u0_u14_u3_n97 ) );
  NOR2_X1 u0_u14_u3_U74 (.A2( u0_u14_X_23 ) , .ZN( u0_u14_u3_n141 ) , .A1( u0_u14_u3_n166 ) );
  NOR2_X1 u0_u14_u3_U75 (.A2( u0_u14_X_19 ) , .A1( u0_u14_u3_n172 ) , .ZN( u0_u14_u3_n96 ) );
  NAND2_X1 u0_u14_u3_U76 (.A1( u0_u14_X_22 ) , .A2( u0_u14_X_23 ) , .ZN( u0_u14_u3_n154 ) );
  NAND2_X1 u0_u14_u3_U77 (.A1( u0_u14_X_23 ) , .ZN( u0_u14_u3_n149 ) , .A2( u0_u14_u3_n166 ) );
  NOR2_X1 u0_u14_u3_U78 (.A2( u0_u14_X_22 ) , .A1( u0_u14_X_23 ) , .ZN( u0_u14_u3_n121 ) );
  AND2_X1 u0_u14_u3_U79 (.A1( u0_u14_X_24 ) , .ZN( u0_u14_u3_n101 ) , .A2( u0_u14_u3_n171 ) );
  AND3_X1 u0_u14_u3_U8 (.A3( u0_u14_u3_n144 ) , .A2( u0_u14_u3_n145 ) , .A1( u0_u14_u3_n146 ) , .ZN( u0_u14_u3_n147 ) );
  AND2_X1 u0_u14_u3_U80 (.A1( u0_u14_X_19 ) , .ZN( u0_u14_u3_n102 ) , .A2( u0_u14_u3_n172 ) );
  AND2_X1 u0_u14_u3_U81 (.A1( u0_u14_X_21 ) , .A2( u0_u14_X_24 ) , .ZN( u0_u14_u3_n100 ) );
  AND2_X1 u0_u14_u3_U82 (.A2( u0_u14_X_19 ) , .A1( u0_u14_X_20 ) , .ZN( u0_u14_u3_n104 ) );
  INV_X1 u0_u14_u3_U83 (.A( u0_u14_X_22 ) , .ZN( u0_u14_u3_n166 ) );
  INV_X1 u0_u14_u3_U84 (.A( u0_u14_X_21 ) , .ZN( u0_u14_u3_n171 ) );
  INV_X1 u0_u14_u3_U85 (.A( u0_u14_X_20 ) , .ZN( u0_u14_u3_n172 ) );
  NAND4_X1 u0_u14_u3_U86 (.ZN( u0_out14_26 ) , .A4( u0_u14_u3_n109 ) , .A3( u0_u14_u3_n110 ) , .A2( u0_u14_u3_n111 ) , .A1( u0_u14_u3_n173 ) );
  INV_X1 u0_u14_u3_U87 (.ZN( u0_u14_u3_n173 ) , .A( u0_u14_u3_n94 ) );
  OAI21_X1 u0_u14_u3_U88 (.ZN( u0_u14_u3_n111 ) , .B2( u0_u14_u3_n117 ) , .A( u0_u14_u3_n133 ) , .B1( u0_u14_u3_n176 ) );
  NAND4_X1 u0_u14_u3_U89 (.ZN( u0_out14_20 ) , .A4( u0_u14_u3_n122 ) , .A3( u0_u14_u3_n123 ) , .A1( u0_u14_u3_n175 ) , .A2( u0_u14_u3_n180 ) );
  INV_X1 u0_u14_u3_U9 (.A( u0_u14_u3_n143 ) , .ZN( u0_u14_u3_n168 ) );
  INV_X1 u0_u14_u3_U90 (.A( u0_u14_u3_n126 ) , .ZN( u0_u14_u3_n180 ) );
  INV_X1 u0_u14_u3_U91 (.A( u0_u14_u3_n112 ) , .ZN( u0_u14_u3_n175 ) );
  NAND4_X1 u0_u14_u3_U92 (.ZN( u0_out14_1 ) , .A4( u0_u14_u3_n161 ) , .A3( u0_u14_u3_n162 ) , .A2( u0_u14_u3_n163 ) , .A1( u0_u14_u3_n185 ) );
  NAND2_X1 u0_u14_u3_U93 (.ZN( u0_u14_u3_n163 ) , .A2( u0_u14_u3_n170 ) , .A1( u0_u14_u3_n176 ) );
  AOI22_X1 u0_u14_u3_U94 (.B2( u0_u14_u3_n140 ) , .B1( u0_u14_u3_n141 ) , .A2( u0_u14_u3_n142 ) , .ZN( u0_u14_u3_n162 ) , .A1( u0_u14_u3_n177 ) );
  OR4_X1 u0_u14_u3_U95 (.ZN( u0_out14_10 ) , .A4( u0_u14_u3_n136 ) , .A3( u0_u14_u3_n137 ) , .A1( u0_u14_u3_n138 ) , .A2( u0_u14_u3_n139 ) );
  OAI222_X1 u0_u14_u3_U96 (.C1( u0_u14_u3_n128 ) , .ZN( u0_u14_u3_n137 ) , .B1( u0_u14_u3_n148 ) , .A2( u0_u14_u3_n150 ) , .B2( u0_u14_u3_n154 ) , .C2( u0_u14_u3_n164 ) , .A1( u0_u14_u3_n167 ) );
  OAI221_X1 u0_u14_u3_U97 (.A( u0_u14_u3_n134 ) , .B2( u0_u14_u3_n135 ) , .ZN( u0_u14_u3_n136 ) , .C1( u0_u14_u3_n149 ) , .B1( u0_u14_u3_n151 ) , .C2( u0_u14_u3_n183 ) );
  NAND3_X1 u0_u14_u3_U98 (.A1( u0_u14_u3_n114 ) , .ZN( u0_u14_u3_n115 ) , .A2( u0_u14_u3_n145 ) , .A3( u0_u14_u3_n153 ) );
  NAND3_X1 u0_u14_u3_U99 (.ZN( u0_u14_u3_n129 ) , .A2( u0_u14_u3_n144 ) , .A1( u0_u14_u3_n153 ) , .A3( u0_u14_u3_n182 ) );
  XOR2_X1 u0_u1_U10 (.B( u0_K2_45 ) , .A( u0_R0_30 ) , .Z( u0_u1_X_45 ) );
  XOR2_X1 u0_u1_U11 (.B( u0_K2_44 ) , .A( u0_R0_29 ) , .Z( u0_u1_X_44 ) );
  XOR2_X1 u0_u1_U12 (.B( u0_K2_43 ) , .A( u0_R0_28 ) , .Z( u0_u1_X_43 ) );
  XOR2_X1 u0_u1_U7 (.B( u0_K2_48 ) , .A( u0_R0_1 ) , .Z( u0_u1_X_48 ) );
  XOR2_X1 u0_u1_U8 (.B( u0_K2_47 ) , .A( u0_R0_32 ) , .Z( u0_u1_X_47 ) );
  XOR2_X1 u0_u1_U9 (.B( u0_K2_46 ) , .A( u0_R0_31 ) , .Z( u0_u1_X_46 ) );
  AND3_X1 u0_u1_u7_U10 (.A3( u0_u1_u7_n110 ) , .A2( u0_u1_u7_n127 ) , .A1( u0_u1_u7_n132 ) , .ZN( u0_u1_u7_n92 ) );
  OAI21_X1 u0_u1_u7_U11 (.A( u0_u1_u7_n161 ) , .B1( u0_u1_u7_n168 ) , .B2( u0_u1_u7_n173 ) , .ZN( u0_u1_u7_n91 ) );
  AOI211_X1 u0_u1_u7_U12 (.A( u0_u1_u7_n117 ) , .ZN( u0_u1_u7_n118 ) , .C2( u0_u1_u7_n126 ) , .C1( u0_u1_u7_n177 ) , .B( u0_u1_u7_n180 ) );
  OAI22_X1 u0_u1_u7_U13 (.B1( u0_u1_u7_n115 ) , .ZN( u0_u1_u7_n117 ) , .A2( u0_u1_u7_n133 ) , .A1( u0_u1_u7_n137 ) , .B2( u0_u1_u7_n162 ) );
  INV_X1 u0_u1_u7_U14 (.A( u0_u1_u7_n116 ) , .ZN( u0_u1_u7_n180 ) );
  NOR3_X1 u0_u1_u7_U15 (.ZN( u0_u1_u7_n115 ) , .A3( u0_u1_u7_n145 ) , .A2( u0_u1_u7_n168 ) , .A1( u0_u1_u7_n169 ) );
  OAI211_X1 u0_u1_u7_U16 (.B( u0_u1_u7_n122 ) , .A( u0_u1_u7_n123 ) , .C2( u0_u1_u7_n124 ) , .ZN( u0_u1_u7_n154 ) , .C1( u0_u1_u7_n162 ) );
  AOI222_X1 u0_u1_u7_U17 (.ZN( u0_u1_u7_n122 ) , .C2( u0_u1_u7_n126 ) , .C1( u0_u1_u7_n145 ) , .B1( u0_u1_u7_n161 ) , .A2( u0_u1_u7_n165 ) , .B2( u0_u1_u7_n170 ) , .A1( u0_u1_u7_n176 ) );
  INV_X1 u0_u1_u7_U18 (.A( u0_u1_u7_n133 ) , .ZN( u0_u1_u7_n176 ) );
  NOR3_X1 u0_u1_u7_U19 (.A2( u0_u1_u7_n134 ) , .A1( u0_u1_u7_n135 ) , .ZN( u0_u1_u7_n136 ) , .A3( u0_u1_u7_n171 ) );
  NOR2_X1 u0_u1_u7_U20 (.A1( u0_u1_u7_n130 ) , .A2( u0_u1_u7_n134 ) , .ZN( u0_u1_u7_n153 ) );
  INV_X1 u0_u1_u7_U21 (.A( u0_u1_u7_n101 ) , .ZN( u0_u1_u7_n165 ) );
  NOR2_X1 u0_u1_u7_U22 (.ZN( u0_u1_u7_n111 ) , .A2( u0_u1_u7_n134 ) , .A1( u0_u1_u7_n169 ) );
  AOI21_X1 u0_u1_u7_U23 (.ZN( u0_u1_u7_n104 ) , .B2( u0_u1_u7_n112 ) , .B1( u0_u1_u7_n127 ) , .A( u0_u1_u7_n164 ) );
  AOI21_X1 u0_u1_u7_U24 (.ZN( u0_u1_u7_n106 ) , .B1( u0_u1_u7_n133 ) , .B2( u0_u1_u7_n146 ) , .A( u0_u1_u7_n162 ) );
  AOI21_X1 u0_u1_u7_U25 (.A( u0_u1_u7_n101 ) , .ZN( u0_u1_u7_n107 ) , .B2( u0_u1_u7_n128 ) , .B1( u0_u1_u7_n175 ) );
  INV_X1 u0_u1_u7_U26 (.A( u0_u1_u7_n138 ) , .ZN( u0_u1_u7_n171 ) );
  INV_X1 u0_u1_u7_U27 (.A( u0_u1_u7_n131 ) , .ZN( u0_u1_u7_n177 ) );
  INV_X1 u0_u1_u7_U28 (.A( u0_u1_u7_n110 ) , .ZN( u0_u1_u7_n174 ) );
  NAND2_X1 u0_u1_u7_U29 (.A1( u0_u1_u7_n129 ) , .A2( u0_u1_u7_n132 ) , .ZN( u0_u1_u7_n149 ) );
  OAI21_X1 u0_u1_u7_U3 (.ZN( u0_u1_u7_n159 ) , .A( u0_u1_u7_n165 ) , .B2( u0_u1_u7_n171 ) , .B1( u0_u1_u7_n174 ) );
  NAND2_X1 u0_u1_u7_U30 (.A1( u0_u1_u7_n113 ) , .A2( u0_u1_u7_n124 ) , .ZN( u0_u1_u7_n130 ) );
  INV_X1 u0_u1_u7_U31 (.A( u0_u1_u7_n112 ) , .ZN( u0_u1_u7_n173 ) );
  INV_X1 u0_u1_u7_U32 (.A( u0_u1_u7_n128 ) , .ZN( u0_u1_u7_n168 ) );
  INV_X1 u0_u1_u7_U33 (.A( u0_u1_u7_n148 ) , .ZN( u0_u1_u7_n169 ) );
  INV_X1 u0_u1_u7_U34 (.A( u0_u1_u7_n127 ) , .ZN( u0_u1_u7_n179 ) );
  NOR2_X1 u0_u1_u7_U35 (.ZN( u0_u1_u7_n101 ) , .A2( u0_u1_u7_n150 ) , .A1( u0_u1_u7_n156 ) );
  AOI211_X1 u0_u1_u7_U36 (.B( u0_u1_u7_n154 ) , .A( u0_u1_u7_n155 ) , .C1( u0_u1_u7_n156 ) , .ZN( u0_u1_u7_n157 ) , .C2( u0_u1_u7_n172 ) );
  INV_X1 u0_u1_u7_U37 (.A( u0_u1_u7_n153 ) , .ZN( u0_u1_u7_n172 ) );
  AOI211_X1 u0_u1_u7_U38 (.B( u0_u1_u7_n139 ) , .A( u0_u1_u7_n140 ) , .C2( u0_u1_u7_n141 ) , .ZN( u0_u1_u7_n142 ) , .C1( u0_u1_u7_n156 ) );
  NAND4_X1 u0_u1_u7_U39 (.A3( u0_u1_u7_n127 ) , .A2( u0_u1_u7_n128 ) , .A1( u0_u1_u7_n129 ) , .ZN( u0_u1_u7_n141 ) , .A4( u0_u1_u7_n147 ) );
  INV_X1 u0_u1_u7_U4 (.A( u0_u1_u7_n111 ) , .ZN( u0_u1_u7_n170 ) );
  AOI21_X1 u0_u1_u7_U40 (.A( u0_u1_u7_n137 ) , .B1( u0_u1_u7_n138 ) , .ZN( u0_u1_u7_n139 ) , .B2( u0_u1_u7_n146 ) );
  OAI22_X1 u0_u1_u7_U41 (.B1( u0_u1_u7_n136 ) , .ZN( u0_u1_u7_n140 ) , .A1( u0_u1_u7_n153 ) , .B2( u0_u1_u7_n162 ) , .A2( u0_u1_u7_n164 ) );
  AOI21_X1 u0_u1_u7_U42 (.ZN( u0_u1_u7_n123 ) , .B1( u0_u1_u7_n165 ) , .B2( u0_u1_u7_n177 ) , .A( u0_u1_u7_n97 ) );
  AOI21_X1 u0_u1_u7_U43 (.B2( u0_u1_u7_n113 ) , .B1( u0_u1_u7_n124 ) , .A( u0_u1_u7_n125 ) , .ZN( u0_u1_u7_n97 ) );
  INV_X1 u0_u1_u7_U44 (.A( u0_u1_u7_n125 ) , .ZN( u0_u1_u7_n161 ) );
  INV_X1 u0_u1_u7_U45 (.A( u0_u1_u7_n152 ) , .ZN( u0_u1_u7_n162 ) );
  AOI22_X1 u0_u1_u7_U46 (.A2( u0_u1_u7_n114 ) , .ZN( u0_u1_u7_n119 ) , .B1( u0_u1_u7_n130 ) , .A1( u0_u1_u7_n156 ) , .B2( u0_u1_u7_n165 ) );
  NAND2_X1 u0_u1_u7_U47 (.A2( u0_u1_u7_n112 ) , .ZN( u0_u1_u7_n114 ) , .A1( u0_u1_u7_n175 ) );
  AND2_X1 u0_u1_u7_U48 (.ZN( u0_u1_u7_n145 ) , .A2( u0_u1_u7_n98 ) , .A1( u0_u1_u7_n99 ) );
  NOR2_X1 u0_u1_u7_U49 (.ZN( u0_u1_u7_n137 ) , .A1( u0_u1_u7_n150 ) , .A2( u0_u1_u7_n161 ) );
  INV_X1 u0_u1_u7_U5 (.A( u0_u1_u7_n149 ) , .ZN( u0_u1_u7_n175 ) );
  AOI21_X1 u0_u1_u7_U50 (.ZN( u0_u1_u7_n105 ) , .B2( u0_u1_u7_n110 ) , .A( u0_u1_u7_n125 ) , .B1( u0_u1_u7_n147 ) );
  NAND2_X1 u0_u1_u7_U51 (.ZN( u0_u1_u7_n146 ) , .A1( u0_u1_u7_n95 ) , .A2( u0_u1_u7_n98 ) );
  NAND2_X1 u0_u1_u7_U52 (.A2( u0_u1_u7_n103 ) , .ZN( u0_u1_u7_n147 ) , .A1( u0_u1_u7_n93 ) );
  NAND2_X1 u0_u1_u7_U53 (.A1( u0_u1_u7_n103 ) , .ZN( u0_u1_u7_n127 ) , .A2( u0_u1_u7_n99 ) );
  OR2_X1 u0_u1_u7_U54 (.ZN( u0_u1_u7_n126 ) , .A2( u0_u1_u7_n152 ) , .A1( u0_u1_u7_n156 ) );
  NAND2_X1 u0_u1_u7_U55 (.A2( u0_u1_u7_n102 ) , .A1( u0_u1_u7_n103 ) , .ZN( u0_u1_u7_n133 ) );
  NAND2_X1 u0_u1_u7_U56 (.ZN( u0_u1_u7_n112 ) , .A2( u0_u1_u7_n96 ) , .A1( u0_u1_u7_n99 ) );
  NAND2_X1 u0_u1_u7_U57 (.A2( u0_u1_u7_n102 ) , .ZN( u0_u1_u7_n128 ) , .A1( u0_u1_u7_n98 ) );
  NAND2_X1 u0_u1_u7_U58 (.A1( u0_u1_u7_n100 ) , .ZN( u0_u1_u7_n113 ) , .A2( u0_u1_u7_n93 ) );
  NAND2_X1 u0_u1_u7_U59 (.A2( u0_u1_u7_n102 ) , .ZN( u0_u1_u7_n124 ) , .A1( u0_u1_u7_n96 ) );
  INV_X1 u0_u1_u7_U6 (.A( u0_u1_u7_n154 ) , .ZN( u0_u1_u7_n178 ) );
  NAND2_X1 u0_u1_u7_U60 (.ZN( u0_u1_u7_n110 ) , .A1( u0_u1_u7_n95 ) , .A2( u0_u1_u7_n96 ) );
  INV_X1 u0_u1_u7_U61 (.A( u0_u1_u7_n150 ) , .ZN( u0_u1_u7_n164 ) );
  AND2_X1 u0_u1_u7_U62 (.ZN( u0_u1_u7_n134 ) , .A1( u0_u1_u7_n93 ) , .A2( u0_u1_u7_n98 ) );
  NAND2_X1 u0_u1_u7_U63 (.A1( u0_u1_u7_n100 ) , .A2( u0_u1_u7_n102 ) , .ZN( u0_u1_u7_n129 ) );
  NAND2_X1 u0_u1_u7_U64 (.A2( u0_u1_u7_n103 ) , .ZN( u0_u1_u7_n131 ) , .A1( u0_u1_u7_n95 ) );
  NAND2_X1 u0_u1_u7_U65 (.A1( u0_u1_u7_n100 ) , .ZN( u0_u1_u7_n138 ) , .A2( u0_u1_u7_n99 ) );
  NAND2_X1 u0_u1_u7_U66 (.ZN( u0_u1_u7_n132 ) , .A1( u0_u1_u7_n93 ) , .A2( u0_u1_u7_n96 ) );
  NAND2_X1 u0_u1_u7_U67 (.A1( u0_u1_u7_n100 ) , .ZN( u0_u1_u7_n148 ) , .A2( u0_u1_u7_n95 ) );
  NOR2_X1 u0_u1_u7_U68 (.A2( u0_u1_X_47 ) , .ZN( u0_u1_u7_n150 ) , .A1( u0_u1_u7_n163 ) );
  NOR2_X1 u0_u1_u7_U69 (.A2( u0_u1_X_43 ) , .A1( u0_u1_X_44 ) , .ZN( u0_u1_u7_n103 ) );
  AOI211_X1 u0_u1_u7_U7 (.ZN( u0_u1_u7_n116 ) , .A( u0_u1_u7_n155 ) , .C1( u0_u1_u7_n161 ) , .C2( u0_u1_u7_n171 ) , .B( u0_u1_u7_n94 ) );
  NOR2_X1 u0_u1_u7_U70 (.A2( u0_u1_X_48 ) , .A1( u0_u1_u7_n166 ) , .ZN( u0_u1_u7_n95 ) );
  NOR2_X1 u0_u1_u7_U71 (.A2( u0_u1_X_45 ) , .A1( u0_u1_X_48 ) , .ZN( u0_u1_u7_n99 ) );
  NOR2_X1 u0_u1_u7_U72 (.A2( u0_u1_X_44 ) , .A1( u0_u1_u7_n167 ) , .ZN( u0_u1_u7_n98 ) );
  NOR2_X1 u0_u1_u7_U73 (.A2( u0_u1_X_46 ) , .A1( u0_u1_X_47 ) , .ZN( u0_u1_u7_n152 ) );
  AND2_X1 u0_u1_u7_U74 (.A1( u0_u1_X_47 ) , .ZN( u0_u1_u7_n156 ) , .A2( u0_u1_u7_n163 ) );
  NAND2_X1 u0_u1_u7_U75 (.A2( u0_u1_X_46 ) , .A1( u0_u1_X_47 ) , .ZN( u0_u1_u7_n125 ) );
  AND2_X1 u0_u1_u7_U76 (.A2( u0_u1_X_45 ) , .A1( u0_u1_X_48 ) , .ZN( u0_u1_u7_n102 ) );
  AND2_X1 u0_u1_u7_U77 (.A2( u0_u1_X_43 ) , .A1( u0_u1_X_44 ) , .ZN( u0_u1_u7_n96 ) );
  AND2_X1 u0_u1_u7_U78 (.A1( u0_u1_X_44 ) , .ZN( u0_u1_u7_n100 ) , .A2( u0_u1_u7_n167 ) );
  AND2_X1 u0_u1_u7_U79 (.A1( u0_u1_X_48 ) , .A2( u0_u1_u7_n166 ) , .ZN( u0_u1_u7_n93 ) );
  OAI222_X1 u0_u1_u7_U8 (.C2( u0_u1_u7_n101 ) , .B2( u0_u1_u7_n111 ) , .A1( u0_u1_u7_n113 ) , .C1( u0_u1_u7_n146 ) , .A2( u0_u1_u7_n162 ) , .B1( u0_u1_u7_n164 ) , .ZN( u0_u1_u7_n94 ) );
  INV_X1 u0_u1_u7_U80 (.A( u0_u1_X_46 ) , .ZN( u0_u1_u7_n163 ) );
  INV_X1 u0_u1_u7_U81 (.A( u0_u1_X_43 ) , .ZN( u0_u1_u7_n167 ) );
  INV_X1 u0_u1_u7_U82 (.A( u0_u1_X_45 ) , .ZN( u0_u1_u7_n166 ) );
  NAND4_X1 u0_u1_u7_U83 (.ZN( u0_out1_27 ) , .A4( u0_u1_u7_n118 ) , .A3( u0_u1_u7_n119 ) , .A2( u0_u1_u7_n120 ) , .A1( u0_u1_u7_n121 ) );
  OAI21_X1 u0_u1_u7_U84 (.ZN( u0_u1_u7_n121 ) , .B2( u0_u1_u7_n145 ) , .A( u0_u1_u7_n150 ) , .B1( u0_u1_u7_n174 ) );
  OAI21_X1 u0_u1_u7_U85 (.ZN( u0_u1_u7_n120 ) , .A( u0_u1_u7_n161 ) , .B2( u0_u1_u7_n170 ) , .B1( u0_u1_u7_n179 ) );
  NAND4_X1 u0_u1_u7_U86 (.ZN( u0_out1_15 ) , .A4( u0_u1_u7_n142 ) , .A3( u0_u1_u7_n143 ) , .A2( u0_u1_u7_n144 ) , .A1( u0_u1_u7_n178 ) );
  OR2_X1 u0_u1_u7_U87 (.A2( u0_u1_u7_n125 ) , .A1( u0_u1_u7_n129 ) , .ZN( u0_u1_u7_n144 ) );
  AOI22_X1 u0_u1_u7_U88 (.A2( u0_u1_u7_n126 ) , .ZN( u0_u1_u7_n143 ) , .B2( u0_u1_u7_n165 ) , .B1( u0_u1_u7_n173 ) , .A1( u0_u1_u7_n174 ) );
  NAND4_X1 u0_u1_u7_U89 (.ZN( u0_out1_5 ) , .A4( u0_u1_u7_n108 ) , .A3( u0_u1_u7_n109 ) , .A1( u0_u1_u7_n116 ) , .A2( u0_u1_u7_n123 ) );
  OAI221_X1 u0_u1_u7_U9 (.C1( u0_u1_u7_n101 ) , .C2( u0_u1_u7_n147 ) , .ZN( u0_u1_u7_n155 ) , .B2( u0_u1_u7_n162 ) , .A( u0_u1_u7_n91 ) , .B1( u0_u1_u7_n92 ) );
  AOI22_X1 u0_u1_u7_U90 (.ZN( u0_u1_u7_n109 ) , .A2( u0_u1_u7_n126 ) , .B2( u0_u1_u7_n145 ) , .B1( u0_u1_u7_n156 ) , .A1( u0_u1_u7_n171 ) );
  NOR4_X1 u0_u1_u7_U91 (.A4( u0_u1_u7_n104 ) , .A3( u0_u1_u7_n105 ) , .A2( u0_u1_u7_n106 ) , .A1( u0_u1_u7_n107 ) , .ZN( u0_u1_u7_n108 ) );
  NAND4_X1 u0_u1_u7_U92 (.ZN( u0_out1_21 ) , .A4( u0_u1_u7_n157 ) , .A3( u0_u1_u7_n158 ) , .A2( u0_u1_u7_n159 ) , .A1( u0_u1_u7_n160 ) );
  OAI21_X1 u0_u1_u7_U93 (.B1( u0_u1_u7_n145 ) , .ZN( u0_u1_u7_n160 ) , .A( u0_u1_u7_n161 ) , .B2( u0_u1_u7_n177 ) );
  AOI22_X1 u0_u1_u7_U94 (.B2( u0_u1_u7_n149 ) , .B1( u0_u1_u7_n150 ) , .A2( u0_u1_u7_n151 ) , .A1( u0_u1_u7_n152 ) , .ZN( u0_u1_u7_n158 ) );
  NAND3_X1 u0_u1_u7_U95 (.A3( u0_u1_u7_n146 ) , .A2( u0_u1_u7_n147 ) , .A1( u0_u1_u7_n148 ) , .ZN( u0_u1_u7_n151 ) );
  NAND3_X1 u0_u1_u7_U96 (.A3( u0_u1_u7_n131 ) , .A2( u0_u1_u7_n132 ) , .A1( u0_u1_u7_n133 ) , .ZN( u0_u1_u7_n135 ) );
  XOR2_X1 u0_u2_U20 (.B( u0_K3_36 ) , .A( u0_R1_25 ) , .Z( u0_u2_X_36 ) );
  XOR2_X1 u0_u2_U21 (.B( u0_K3_35 ) , .A( u0_R1_24 ) , .Z( u0_u2_X_35 ) );
  XOR2_X1 u0_u2_U22 (.B( u0_K3_34 ) , .A( u0_R1_23 ) , .Z( u0_u2_X_34 ) );
  XOR2_X1 u0_u2_U23 (.B( u0_K3_33 ) , .A( u0_R1_22 ) , .Z( u0_u2_X_33 ) );
  XOR2_X1 u0_u2_U24 (.B( u0_K3_32 ) , .A( u0_R1_21 ) , .Z( u0_u2_X_32 ) );
  XOR2_X1 u0_u2_U25 (.B( u0_K3_31 ) , .A( u0_R1_20 ) , .Z( u0_u2_X_31 ) );
  XOR2_X1 u0_u2_U26 (.B( u0_K3_30 ) , .A( u0_R1_21 ) , .Z( u0_u2_X_30 ) );
  XOR2_X1 u0_u2_U28 (.B( u0_K3_29 ) , .A( u0_R1_20 ) , .Z( u0_u2_X_29 ) );
  XOR2_X1 u0_u2_U29 (.B( u0_K3_28 ) , .A( u0_R1_19 ) , .Z( u0_u2_X_28 ) );
  XOR2_X1 u0_u2_U30 (.B( u0_K3_27 ) , .A( u0_R1_18 ) , .Z( u0_u2_X_27 ) );
  XOR2_X1 u0_u2_U31 (.B( u0_K3_26 ) , .A( u0_R1_17 ) , .Z( u0_u2_X_26 ) );
  XOR2_X1 u0_u2_U32 (.B( u0_K3_25 ) , .A( u0_R1_16 ) , .Z( u0_u2_X_25 ) );
  OAI22_X1 u0_u2_u4_U10 (.B2( u0_u2_u4_n135 ) , .ZN( u0_u2_u4_n137 ) , .B1( u0_u2_u4_n153 ) , .A1( u0_u2_u4_n155 ) , .A2( u0_u2_u4_n171 ) );
  AND3_X1 u0_u2_u4_U11 (.A2( u0_u2_u4_n134 ) , .ZN( u0_u2_u4_n135 ) , .A3( u0_u2_u4_n145 ) , .A1( u0_u2_u4_n157 ) );
  NAND2_X1 u0_u2_u4_U12 (.ZN( u0_u2_u4_n132 ) , .A2( u0_u2_u4_n170 ) , .A1( u0_u2_u4_n173 ) );
  AOI21_X1 u0_u2_u4_U13 (.B2( u0_u2_u4_n160 ) , .B1( u0_u2_u4_n161 ) , .ZN( u0_u2_u4_n162 ) , .A( u0_u2_u4_n170 ) );
  AOI21_X1 u0_u2_u4_U14 (.ZN( u0_u2_u4_n107 ) , .B2( u0_u2_u4_n143 ) , .A( u0_u2_u4_n174 ) , .B1( u0_u2_u4_n184 ) );
  AOI21_X1 u0_u2_u4_U15 (.B2( u0_u2_u4_n158 ) , .B1( u0_u2_u4_n159 ) , .ZN( u0_u2_u4_n163 ) , .A( u0_u2_u4_n174 ) );
  AOI21_X1 u0_u2_u4_U16 (.A( u0_u2_u4_n153 ) , .B2( u0_u2_u4_n154 ) , .B1( u0_u2_u4_n155 ) , .ZN( u0_u2_u4_n165 ) );
  AOI21_X1 u0_u2_u4_U17 (.A( u0_u2_u4_n156 ) , .B2( u0_u2_u4_n157 ) , .ZN( u0_u2_u4_n164 ) , .B1( u0_u2_u4_n184 ) );
  INV_X1 u0_u2_u4_U18 (.A( u0_u2_u4_n138 ) , .ZN( u0_u2_u4_n170 ) );
  AND2_X1 u0_u2_u4_U19 (.A2( u0_u2_u4_n120 ) , .ZN( u0_u2_u4_n155 ) , .A1( u0_u2_u4_n160 ) );
  INV_X1 u0_u2_u4_U20 (.A( u0_u2_u4_n156 ) , .ZN( u0_u2_u4_n175 ) );
  NAND2_X1 u0_u2_u4_U21 (.A2( u0_u2_u4_n118 ) , .ZN( u0_u2_u4_n131 ) , .A1( u0_u2_u4_n147 ) );
  NAND2_X1 u0_u2_u4_U22 (.A1( u0_u2_u4_n119 ) , .A2( u0_u2_u4_n120 ) , .ZN( u0_u2_u4_n130 ) );
  NAND2_X1 u0_u2_u4_U23 (.ZN( u0_u2_u4_n117 ) , .A2( u0_u2_u4_n118 ) , .A1( u0_u2_u4_n148 ) );
  NAND2_X1 u0_u2_u4_U24 (.ZN( u0_u2_u4_n129 ) , .A1( u0_u2_u4_n134 ) , .A2( u0_u2_u4_n148 ) );
  AND3_X1 u0_u2_u4_U25 (.A1( u0_u2_u4_n119 ) , .A2( u0_u2_u4_n143 ) , .A3( u0_u2_u4_n154 ) , .ZN( u0_u2_u4_n161 ) );
  AND2_X1 u0_u2_u4_U26 (.A1( u0_u2_u4_n145 ) , .A2( u0_u2_u4_n147 ) , .ZN( u0_u2_u4_n159 ) );
  OR3_X1 u0_u2_u4_U27 (.A3( u0_u2_u4_n114 ) , .A2( u0_u2_u4_n115 ) , .A1( u0_u2_u4_n116 ) , .ZN( u0_u2_u4_n136 ) );
  AOI21_X1 u0_u2_u4_U28 (.A( u0_u2_u4_n113 ) , .ZN( u0_u2_u4_n116 ) , .B2( u0_u2_u4_n173 ) , .B1( u0_u2_u4_n174 ) );
  AOI21_X1 u0_u2_u4_U29 (.ZN( u0_u2_u4_n115 ) , .B2( u0_u2_u4_n145 ) , .B1( u0_u2_u4_n146 ) , .A( u0_u2_u4_n156 ) );
  NOR2_X1 u0_u2_u4_U3 (.ZN( u0_u2_u4_n121 ) , .A1( u0_u2_u4_n181 ) , .A2( u0_u2_u4_n182 ) );
  OAI22_X1 u0_u2_u4_U30 (.ZN( u0_u2_u4_n114 ) , .A2( u0_u2_u4_n121 ) , .B1( u0_u2_u4_n160 ) , .B2( u0_u2_u4_n170 ) , .A1( u0_u2_u4_n171 ) );
  INV_X1 u0_u2_u4_U31 (.A( u0_u2_u4_n158 ) , .ZN( u0_u2_u4_n182 ) );
  INV_X1 u0_u2_u4_U32 (.ZN( u0_u2_u4_n181 ) , .A( u0_u2_u4_n96 ) );
  INV_X1 u0_u2_u4_U33 (.A( u0_u2_u4_n144 ) , .ZN( u0_u2_u4_n179 ) );
  INV_X1 u0_u2_u4_U34 (.A( u0_u2_u4_n157 ) , .ZN( u0_u2_u4_n178 ) );
  NAND2_X1 u0_u2_u4_U35 (.A2( u0_u2_u4_n154 ) , .A1( u0_u2_u4_n96 ) , .ZN( u0_u2_u4_n97 ) );
  INV_X1 u0_u2_u4_U36 (.ZN( u0_u2_u4_n186 ) , .A( u0_u2_u4_n95 ) );
  OAI221_X1 u0_u2_u4_U37 (.C1( u0_u2_u4_n134 ) , .B1( u0_u2_u4_n158 ) , .B2( u0_u2_u4_n171 ) , .C2( u0_u2_u4_n173 ) , .A( u0_u2_u4_n94 ) , .ZN( u0_u2_u4_n95 ) );
  AOI222_X1 u0_u2_u4_U38 (.B2( u0_u2_u4_n132 ) , .A1( u0_u2_u4_n138 ) , .C2( u0_u2_u4_n175 ) , .A2( u0_u2_u4_n179 ) , .C1( u0_u2_u4_n181 ) , .B1( u0_u2_u4_n185 ) , .ZN( u0_u2_u4_n94 ) );
  INV_X1 u0_u2_u4_U39 (.A( u0_u2_u4_n113 ) , .ZN( u0_u2_u4_n185 ) );
  INV_X1 u0_u2_u4_U4 (.A( u0_u2_u4_n117 ) , .ZN( u0_u2_u4_n184 ) );
  INV_X1 u0_u2_u4_U40 (.A( u0_u2_u4_n143 ) , .ZN( u0_u2_u4_n183 ) );
  NOR2_X1 u0_u2_u4_U41 (.ZN( u0_u2_u4_n138 ) , .A1( u0_u2_u4_n168 ) , .A2( u0_u2_u4_n169 ) );
  NOR2_X1 u0_u2_u4_U42 (.A1( u0_u2_u4_n150 ) , .A2( u0_u2_u4_n152 ) , .ZN( u0_u2_u4_n153 ) );
  NOR2_X1 u0_u2_u4_U43 (.A2( u0_u2_u4_n128 ) , .A1( u0_u2_u4_n138 ) , .ZN( u0_u2_u4_n156 ) );
  AOI22_X1 u0_u2_u4_U44 (.B2( u0_u2_u4_n122 ) , .A1( u0_u2_u4_n123 ) , .ZN( u0_u2_u4_n124 ) , .B1( u0_u2_u4_n128 ) , .A2( u0_u2_u4_n172 ) );
  INV_X1 u0_u2_u4_U45 (.A( u0_u2_u4_n153 ) , .ZN( u0_u2_u4_n172 ) );
  NAND2_X1 u0_u2_u4_U46 (.A2( u0_u2_u4_n120 ) , .ZN( u0_u2_u4_n123 ) , .A1( u0_u2_u4_n161 ) );
  AOI22_X1 u0_u2_u4_U47 (.B2( u0_u2_u4_n132 ) , .A2( u0_u2_u4_n133 ) , .ZN( u0_u2_u4_n140 ) , .A1( u0_u2_u4_n150 ) , .B1( u0_u2_u4_n179 ) );
  NAND2_X1 u0_u2_u4_U48 (.ZN( u0_u2_u4_n133 ) , .A2( u0_u2_u4_n146 ) , .A1( u0_u2_u4_n154 ) );
  NAND2_X1 u0_u2_u4_U49 (.A1( u0_u2_u4_n103 ) , .ZN( u0_u2_u4_n154 ) , .A2( u0_u2_u4_n98 ) );
  NOR4_X1 u0_u2_u4_U5 (.A4( u0_u2_u4_n106 ) , .A3( u0_u2_u4_n107 ) , .A2( u0_u2_u4_n108 ) , .A1( u0_u2_u4_n109 ) , .ZN( u0_u2_u4_n110 ) );
  NAND2_X1 u0_u2_u4_U50 (.A1( u0_u2_u4_n101 ) , .ZN( u0_u2_u4_n158 ) , .A2( u0_u2_u4_n99 ) );
  AOI21_X1 u0_u2_u4_U51 (.ZN( u0_u2_u4_n127 ) , .A( u0_u2_u4_n136 ) , .B2( u0_u2_u4_n150 ) , .B1( u0_u2_u4_n180 ) );
  INV_X1 u0_u2_u4_U52 (.A( u0_u2_u4_n160 ) , .ZN( u0_u2_u4_n180 ) );
  NAND2_X1 u0_u2_u4_U53 (.A2( u0_u2_u4_n104 ) , .A1( u0_u2_u4_n105 ) , .ZN( u0_u2_u4_n146 ) );
  NAND2_X1 u0_u2_u4_U54 (.A2( u0_u2_u4_n101 ) , .A1( u0_u2_u4_n102 ) , .ZN( u0_u2_u4_n160 ) );
  NAND2_X1 u0_u2_u4_U55 (.ZN( u0_u2_u4_n134 ) , .A1( u0_u2_u4_n98 ) , .A2( u0_u2_u4_n99 ) );
  NAND2_X1 u0_u2_u4_U56 (.A1( u0_u2_u4_n103 ) , .A2( u0_u2_u4_n104 ) , .ZN( u0_u2_u4_n143 ) );
  NAND2_X1 u0_u2_u4_U57 (.A2( u0_u2_u4_n105 ) , .ZN( u0_u2_u4_n145 ) , .A1( u0_u2_u4_n98 ) );
  NAND2_X1 u0_u2_u4_U58 (.A1( u0_u2_u4_n100 ) , .A2( u0_u2_u4_n105 ) , .ZN( u0_u2_u4_n120 ) );
  NAND2_X1 u0_u2_u4_U59 (.A1( u0_u2_u4_n102 ) , .A2( u0_u2_u4_n104 ) , .ZN( u0_u2_u4_n148 ) );
  AOI21_X1 u0_u2_u4_U6 (.ZN( u0_u2_u4_n106 ) , .B2( u0_u2_u4_n146 ) , .B1( u0_u2_u4_n158 ) , .A( u0_u2_u4_n170 ) );
  NAND2_X1 u0_u2_u4_U60 (.A2( u0_u2_u4_n100 ) , .A1( u0_u2_u4_n103 ) , .ZN( u0_u2_u4_n157 ) );
  INV_X1 u0_u2_u4_U61 (.A( u0_u2_u4_n150 ) , .ZN( u0_u2_u4_n173 ) );
  INV_X1 u0_u2_u4_U62 (.A( u0_u2_u4_n152 ) , .ZN( u0_u2_u4_n171 ) );
  NAND2_X1 u0_u2_u4_U63 (.A1( u0_u2_u4_n100 ) , .ZN( u0_u2_u4_n118 ) , .A2( u0_u2_u4_n99 ) );
  NAND2_X1 u0_u2_u4_U64 (.A2( u0_u2_u4_n100 ) , .A1( u0_u2_u4_n102 ) , .ZN( u0_u2_u4_n144 ) );
  NAND2_X1 u0_u2_u4_U65 (.A2( u0_u2_u4_n101 ) , .A1( u0_u2_u4_n105 ) , .ZN( u0_u2_u4_n96 ) );
  INV_X1 u0_u2_u4_U66 (.A( u0_u2_u4_n128 ) , .ZN( u0_u2_u4_n174 ) );
  NAND2_X1 u0_u2_u4_U67 (.A2( u0_u2_u4_n102 ) , .ZN( u0_u2_u4_n119 ) , .A1( u0_u2_u4_n98 ) );
  NAND2_X1 u0_u2_u4_U68 (.A2( u0_u2_u4_n101 ) , .A1( u0_u2_u4_n103 ) , .ZN( u0_u2_u4_n147 ) );
  NAND2_X1 u0_u2_u4_U69 (.A2( u0_u2_u4_n104 ) , .ZN( u0_u2_u4_n113 ) , .A1( u0_u2_u4_n99 ) );
  AOI21_X1 u0_u2_u4_U7 (.ZN( u0_u2_u4_n108 ) , .B2( u0_u2_u4_n134 ) , .B1( u0_u2_u4_n155 ) , .A( u0_u2_u4_n156 ) );
  NOR2_X1 u0_u2_u4_U70 (.A2( u0_u2_X_28 ) , .ZN( u0_u2_u4_n150 ) , .A1( u0_u2_u4_n168 ) );
  NOR2_X1 u0_u2_u4_U71 (.A2( u0_u2_X_29 ) , .ZN( u0_u2_u4_n152 ) , .A1( u0_u2_u4_n169 ) );
  NOR2_X1 u0_u2_u4_U72 (.A2( u0_u2_X_30 ) , .ZN( u0_u2_u4_n105 ) , .A1( u0_u2_u4_n176 ) );
  NOR2_X1 u0_u2_u4_U73 (.A2( u0_u2_X_26 ) , .ZN( u0_u2_u4_n100 ) , .A1( u0_u2_u4_n177 ) );
  NOR2_X1 u0_u2_u4_U74 (.A2( u0_u2_X_28 ) , .A1( u0_u2_X_29 ) , .ZN( u0_u2_u4_n128 ) );
  NOR2_X1 u0_u2_u4_U75 (.A2( u0_u2_X_27 ) , .A1( u0_u2_X_30 ) , .ZN( u0_u2_u4_n102 ) );
  NOR2_X1 u0_u2_u4_U76 (.A2( u0_u2_X_25 ) , .A1( u0_u2_X_26 ) , .ZN( u0_u2_u4_n98 ) );
  AND2_X1 u0_u2_u4_U77 (.A2( u0_u2_X_25 ) , .A1( u0_u2_X_26 ) , .ZN( u0_u2_u4_n104 ) );
  AND2_X1 u0_u2_u4_U78 (.A1( u0_u2_X_30 ) , .A2( u0_u2_u4_n176 ) , .ZN( u0_u2_u4_n99 ) );
  AND2_X1 u0_u2_u4_U79 (.A1( u0_u2_X_26 ) , .ZN( u0_u2_u4_n101 ) , .A2( u0_u2_u4_n177 ) );
  AOI21_X1 u0_u2_u4_U8 (.ZN( u0_u2_u4_n109 ) , .A( u0_u2_u4_n153 ) , .B1( u0_u2_u4_n159 ) , .B2( u0_u2_u4_n184 ) );
  AND2_X1 u0_u2_u4_U80 (.A1( u0_u2_X_27 ) , .A2( u0_u2_X_30 ) , .ZN( u0_u2_u4_n103 ) );
  INV_X1 u0_u2_u4_U81 (.A( u0_u2_X_28 ) , .ZN( u0_u2_u4_n169 ) );
  INV_X1 u0_u2_u4_U82 (.A( u0_u2_X_29 ) , .ZN( u0_u2_u4_n168 ) );
  INV_X1 u0_u2_u4_U83 (.A( u0_u2_X_25 ) , .ZN( u0_u2_u4_n177 ) );
  INV_X1 u0_u2_u4_U84 (.A( u0_u2_X_27 ) , .ZN( u0_u2_u4_n176 ) );
  NAND4_X1 u0_u2_u4_U85 (.ZN( u0_out2_25 ) , .A4( u0_u2_u4_n139 ) , .A3( u0_u2_u4_n140 ) , .A2( u0_u2_u4_n141 ) , .A1( u0_u2_u4_n142 ) );
  OAI21_X1 u0_u2_u4_U86 (.A( u0_u2_u4_n128 ) , .B2( u0_u2_u4_n129 ) , .B1( u0_u2_u4_n130 ) , .ZN( u0_u2_u4_n142 ) );
  OAI21_X1 u0_u2_u4_U87 (.B2( u0_u2_u4_n131 ) , .ZN( u0_u2_u4_n141 ) , .A( u0_u2_u4_n175 ) , .B1( u0_u2_u4_n183 ) );
  NAND4_X1 u0_u2_u4_U88 (.ZN( u0_out2_14 ) , .A4( u0_u2_u4_n124 ) , .A3( u0_u2_u4_n125 ) , .A2( u0_u2_u4_n126 ) , .A1( u0_u2_u4_n127 ) );
  AOI22_X1 u0_u2_u4_U89 (.B2( u0_u2_u4_n117 ) , .ZN( u0_u2_u4_n126 ) , .A1( u0_u2_u4_n129 ) , .B1( u0_u2_u4_n152 ) , .A2( u0_u2_u4_n175 ) );
  AOI211_X1 u0_u2_u4_U9 (.B( u0_u2_u4_n136 ) , .A( u0_u2_u4_n137 ) , .C2( u0_u2_u4_n138 ) , .ZN( u0_u2_u4_n139 ) , .C1( u0_u2_u4_n182 ) );
  AOI22_X1 u0_u2_u4_U90 (.ZN( u0_u2_u4_n125 ) , .B2( u0_u2_u4_n131 ) , .A2( u0_u2_u4_n132 ) , .B1( u0_u2_u4_n138 ) , .A1( u0_u2_u4_n178 ) );
  NAND4_X1 u0_u2_u4_U91 (.ZN( u0_out2_8 ) , .A4( u0_u2_u4_n110 ) , .A3( u0_u2_u4_n111 ) , .A2( u0_u2_u4_n112 ) , .A1( u0_u2_u4_n186 ) );
  NAND2_X1 u0_u2_u4_U92 (.ZN( u0_u2_u4_n112 ) , .A2( u0_u2_u4_n130 ) , .A1( u0_u2_u4_n150 ) );
  AOI22_X1 u0_u2_u4_U93 (.ZN( u0_u2_u4_n111 ) , .B2( u0_u2_u4_n132 ) , .A1( u0_u2_u4_n152 ) , .B1( u0_u2_u4_n178 ) , .A2( u0_u2_u4_n97 ) );
  AOI22_X1 u0_u2_u4_U94 (.B2( u0_u2_u4_n149 ) , .B1( u0_u2_u4_n150 ) , .A2( u0_u2_u4_n151 ) , .A1( u0_u2_u4_n152 ) , .ZN( u0_u2_u4_n167 ) );
  NOR4_X1 u0_u2_u4_U95 (.A4( u0_u2_u4_n162 ) , .A3( u0_u2_u4_n163 ) , .A2( u0_u2_u4_n164 ) , .A1( u0_u2_u4_n165 ) , .ZN( u0_u2_u4_n166 ) );
  NAND3_X1 u0_u2_u4_U96 (.ZN( u0_out2_3 ) , .A3( u0_u2_u4_n166 ) , .A1( u0_u2_u4_n167 ) , .A2( u0_u2_u4_n186 ) );
  NAND3_X1 u0_u2_u4_U97 (.A3( u0_u2_u4_n146 ) , .A2( u0_u2_u4_n147 ) , .A1( u0_u2_u4_n148 ) , .ZN( u0_u2_u4_n149 ) );
  NAND3_X1 u0_u2_u4_U98 (.A3( u0_u2_u4_n143 ) , .A2( u0_u2_u4_n144 ) , .A1( u0_u2_u4_n145 ) , .ZN( u0_u2_u4_n151 ) );
  NAND3_X1 u0_u2_u4_U99 (.A3( u0_u2_u4_n121 ) , .ZN( u0_u2_u4_n122 ) , .A2( u0_u2_u4_n144 ) , .A1( u0_u2_u4_n154 ) );
  INV_X1 u0_u2_u5_U10 (.A( u0_u2_u5_n121 ) , .ZN( u0_u2_u5_n177 ) );
  AOI222_X1 u0_u2_u5_U100 (.ZN( u0_u2_u5_n113 ) , .A1( u0_u2_u5_n131 ) , .C1( u0_u2_u5_n148 ) , .B2( u0_u2_u5_n174 ) , .C2( u0_u2_u5_n178 ) , .A2( u0_u2_u5_n179 ) , .B1( u0_u2_u5_n99 ) );
  NAND4_X1 u0_u2_u5_U101 (.ZN( u0_out2_29 ) , .A4( u0_u2_u5_n129 ) , .A3( u0_u2_u5_n130 ) , .A2( u0_u2_u5_n168 ) , .A1( u0_u2_u5_n196 ) );
  AOI221_X1 u0_u2_u5_U102 (.A( u0_u2_u5_n128 ) , .ZN( u0_u2_u5_n129 ) , .C2( u0_u2_u5_n132 ) , .B2( u0_u2_u5_n159 ) , .B1( u0_u2_u5_n176 ) , .C1( u0_u2_u5_n184 ) );
  AOI222_X1 u0_u2_u5_U103 (.ZN( u0_u2_u5_n130 ) , .A2( u0_u2_u5_n146 ) , .B1( u0_u2_u5_n147 ) , .C2( u0_u2_u5_n175 ) , .B2( u0_u2_u5_n179 ) , .A1( u0_u2_u5_n188 ) , .C1( u0_u2_u5_n194 ) );
  NAND3_X1 u0_u2_u5_U104 (.A2( u0_u2_u5_n154 ) , .A3( u0_u2_u5_n158 ) , .A1( u0_u2_u5_n161 ) , .ZN( u0_u2_u5_n99 ) );
  NOR2_X1 u0_u2_u5_U11 (.ZN( u0_u2_u5_n160 ) , .A2( u0_u2_u5_n173 ) , .A1( u0_u2_u5_n177 ) );
  INV_X1 u0_u2_u5_U12 (.A( u0_u2_u5_n150 ) , .ZN( u0_u2_u5_n174 ) );
  AOI21_X1 u0_u2_u5_U13 (.A( u0_u2_u5_n160 ) , .B2( u0_u2_u5_n161 ) , .ZN( u0_u2_u5_n162 ) , .B1( u0_u2_u5_n192 ) );
  INV_X1 u0_u2_u5_U14 (.A( u0_u2_u5_n159 ) , .ZN( u0_u2_u5_n192 ) );
  AOI21_X1 u0_u2_u5_U15 (.A( u0_u2_u5_n156 ) , .B2( u0_u2_u5_n157 ) , .B1( u0_u2_u5_n158 ) , .ZN( u0_u2_u5_n163 ) );
  AOI21_X1 u0_u2_u5_U16 (.B2( u0_u2_u5_n139 ) , .B1( u0_u2_u5_n140 ) , .ZN( u0_u2_u5_n141 ) , .A( u0_u2_u5_n150 ) );
  OAI21_X1 u0_u2_u5_U17 (.A( u0_u2_u5_n133 ) , .B2( u0_u2_u5_n134 ) , .B1( u0_u2_u5_n135 ) , .ZN( u0_u2_u5_n142 ) );
  OAI21_X1 u0_u2_u5_U18 (.ZN( u0_u2_u5_n133 ) , .B2( u0_u2_u5_n147 ) , .A( u0_u2_u5_n173 ) , .B1( u0_u2_u5_n188 ) );
  NAND2_X1 u0_u2_u5_U19 (.A2( u0_u2_u5_n119 ) , .A1( u0_u2_u5_n123 ) , .ZN( u0_u2_u5_n137 ) );
  INV_X1 u0_u2_u5_U20 (.A( u0_u2_u5_n155 ) , .ZN( u0_u2_u5_n194 ) );
  NAND2_X1 u0_u2_u5_U21 (.A1( u0_u2_u5_n121 ) , .ZN( u0_u2_u5_n132 ) , .A2( u0_u2_u5_n172 ) );
  NAND2_X1 u0_u2_u5_U22 (.A2( u0_u2_u5_n122 ) , .ZN( u0_u2_u5_n136 ) , .A1( u0_u2_u5_n154 ) );
  NAND2_X1 u0_u2_u5_U23 (.A2( u0_u2_u5_n119 ) , .A1( u0_u2_u5_n120 ) , .ZN( u0_u2_u5_n159 ) );
  INV_X1 u0_u2_u5_U24 (.A( u0_u2_u5_n156 ) , .ZN( u0_u2_u5_n175 ) );
  INV_X1 u0_u2_u5_U25 (.A( u0_u2_u5_n158 ) , .ZN( u0_u2_u5_n188 ) );
  INV_X1 u0_u2_u5_U26 (.A( u0_u2_u5_n152 ) , .ZN( u0_u2_u5_n179 ) );
  INV_X1 u0_u2_u5_U27 (.A( u0_u2_u5_n140 ) , .ZN( u0_u2_u5_n182 ) );
  INV_X1 u0_u2_u5_U28 (.A( u0_u2_u5_n151 ) , .ZN( u0_u2_u5_n183 ) );
  INV_X1 u0_u2_u5_U29 (.A( u0_u2_u5_n123 ) , .ZN( u0_u2_u5_n185 ) );
  NOR2_X1 u0_u2_u5_U3 (.ZN( u0_u2_u5_n134 ) , .A1( u0_u2_u5_n183 ) , .A2( u0_u2_u5_n190 ) );
  INV_X1 u0_u2_u5_U30 (.A( u0_u2_u5_n161 ) , .ZN( u0_u2_u5_n184 ) );
  INV_X1 u0_u2_u5_U31 (.A( u0_u2_u5_n139 ) , .ZN( u0_u2_u5_n189 ) );
  INV_X1 u0_u2_u5_U32 (.A( u0_u2_u5_n157 ) , .ZN( u0_u2_u5_n190 ) );
  INV_X1 u0_u2_u5_U33 (.A( u0_u2_u5_n120 ) , .ZN( u0_u2_u5_n193 ) );
  NAND2_X1 u0_u2_u5_U34 (.ZN( u0_u2_u5_n111 ) , .A1( u0_u2_u5_n140 ) , .A2( u0_u2_u5_n155 ) );
  INV_X1 u0_u2_u5_U35 (.A( u0_u2_u5_n117 ) , .ZN( u0_u2_u5_n196 ) );
  OAI221_X1 u0_u2_u5_U36 (.A( u0_u2_u5_n116 ) , .ZN( u0_u2_u5_n117 ) , .B2( u0_u2_u5_n119 ) , .C1( u0_u2_u5_n153 ) , .C2( u0_u2_u5_n158 ) , .B1( u0_u2_u5_n172 ) );
  AOI222_X1 u0_u2_u5_U37 (.ZN( u0_u2_u5_n116 ) , .B2( u0_u2_u5_n145 ) , .C1( u0_u2_u5_n148 ) , .A2( u0_u2_u5_n174 ) , .C2( u0_u2_u5_n177 ) , .B1( u0_u2_u5_n187 ) , .A1( u0_u2_u5_n193 ) );
  INV_X1 u0_u2_u5_U38 (.A( u0_u2_u5_n115 ) , .ZN( u0_u2_u5_n187 ) );
  NOR2_X1 u0_u2_u5_U39 (.ZN( u0_u2_u5_n100 ) , .A1( u0_u2_u5_n170 ) , .A2( u0_u2_u5_n180 ) );
  INV_X1 u0_u2_u5_U4 (.A( u0_u2_u5_n138 ) , .ZN( u0_u2_u5_n191 ) );
  AOI22_X1 u0_u2_u5_U40 (.B2( u0_u2_u5_n131 ) , .A2( u0_u2_u5_n146 ) , .ZN( u0_u2_u5_n169 ) , .B1( u0_u2_u5_n174 ) , .A1( u0_u2_u5_n185 ) );
  NOR2_X1 u0_u2_u5_U41 (.A1( u0_u2_u5_n146 ) , .ZN( u0_u2_u5_n150 ) , .A2( u0_u2_u5_n173 ) );
  AOI21_X1 u0_u2_u5_U42 (.A( u0_u2_u5_n118 ) , .B2( u0_u2_u5_n145 ) , .ZN( u0_u2_u5_n168 ) , .B1( u0_u2_u5_n186 ) );
  INV_X1 u0_u2_u5_U43 (.A( u0_u2_u5_n122 ) , .ZN( u0_u2_u5_n186 ) );
  NOR2_X1 u0_u2_u5_U44 (.A1( u0_u2_u5_n146 ) , .ZN( u0_u2_u5_n152 ) , .A2( u0_u2_u5_n176 ) );
  NOR2_X1 u0_u2_u5_U45 (.A1( u0_u2_u5_n115 ) , .ZN( u0_u2_u5_n118 ) , .A2( u0_u2_u5_n153 ) );
  NOR2_X1 u0_u2_u5_U46 (.A2( u0_u2_u5_n145 ) , .ZN( u0_u2_u5_n156 ) , .A1( u0_u2_u5_n174 ) );
  NOR2_X1 u0_u2_u5_U47 (.ZN( u0_u2_u5_n121 ) , .A2( u0_u2_u5_n145 ) , .A1( u0_u2_u5_n176 ) );
  AOI22_X1 u0_u2_u5_U48 (.ZN( u0_u2_u5_n114 ) , .A2( u0_u2_u5_n137 ) , .A1( u0_u2_u5_n145 ) , .B2( u0_u2_u5_n175 ) , .B1( u0_u2_u5_n193 ) );
  AOI21_X1 u0_u2_u5_U49 (.A( u0_u2_u5_n153 ) , .B2( u0_u2_u5_n154 ) , .B1( u0_u2_u5_n155 ) , .ZN( u0_u2_u5_n164 ) );
  OAI21_X1 u0_u2_u5_U5 (.B2( u0_u2_u5_n136 ) , .B1( u0_u2_u5_n137 ) , .ZN( u0_u2_u5_n138 ) , .A( u0_u2_u5_n177 ) );
  AOI21_X1 u0_u2_u5_U50 (.ZN( u0_u2_u5_n110 ) , .B1( u0_u2_u5_n122 ) , .B2( u0_u2_u5_n139 ) , .A( u0_u2_u5_n153 ) );
  INV_X1 u0_u2_u5_U51 (.A( u0_u2_u5_n153 ) , .ZN( u0_u2_u5_n176 ) );
  INV_X1 u0_u2_u5_U52 (.A( u0_u2_u5_n126 ) , .ZN( u0_u2_u5_n173 ) );
  AND2_X1 u0_u2_u5_U53 (.A2( u0_u2_u5_n104 ) , .A1( u0_u2_u5_n107 ) , .ZN( u0_u2_u5_n147 ) );
  AND2_X1 u0_u2_u5_U54 (.A2( u0_u2_u5_n104 ) , .A1( u0_u2_u5_n108 ) , .ZN( u0_u2_u5_n148 ) );
  NAND2_X1 u0_u2_u5_U55 (.A1( u0_u2_u5_n105 ) , .A2( u0_u2_u5_n106 ) , .ZN( u0_u2_u5_n158 ) );
  NAND2_X1 u0_u2_u5_U56 (.A2( u0_u2_u5_n108 ) , .A1( u0_u2_u5_n109 ) , .ZN( u0_u2_u5_n139 ) );
  NAND2_X1 u0_u2_u5_U57 (.A1( u0_u2_u5_n106 ) , .A2( u0_u2_u5_n108 ) , .ZN( u0_u2_u5_n119 ) );
  OAI211_X1 u0_u2_u5_U58 (.B( u0_u2_u5_n124 ) , .A( u0_u2_u5_n125 ) , .C2( u0_u2_u5_n126 ) , .C1( u0_u2_u5_n127 ) , .ZN( u0_u2_u5_n128 ) );
  NOR3_X1 u0_u2_u5_U59 (.ZN( u0_u2_u5_n127 ) , .A1( u0_u2_u5_n136 ) , .A3( u0_u2_u5_n148 ) , .A2( u0_u2_u5_n182 ) );
  INV_X1 u0_u2_u5_U6 (.A( u0_u2_u5_n135 ) , .ZN( u0_u2_u5_n178 ) );
  OAI21_X1 u0_u2_u5_U60 (.ZN( u0_u2_u5_n124 ) , .A( u0_u2_u5_n177 ) , .B2( u0_u2_u5_n183 ) , .B1( u0_u2_u5_n189 ) );
  OAI21_X1 u0_u2_u5_U61 (.ZN( u0_u2_u5_n125 ) , .A( u0_u2_u5_n174 ) , .B2( u0_u2_u5_n185 ) , .B1( u0_u2_u5_n190 ) );
  NAND2_X1 u0_u2_u5_U62 (.A2( u0_u2_u5_n103 ) , .A1( u0_u2_u5_n105 ) , .ZN( u0_u2_u5_n140 ) );
  NAND2_X1 u0_u2_u5_U63 (.A2( u0_u2_u5_n104 ) , .A1( u0_u2_u5_n105 ) , .ZN( u0_u2_u5_n155 ) );
  NAND2_X1 u0_u2_u5_U64 (.A2( u0_u2_u5_n106 ) , .A1( u0_u2_u5_n107 ) , .ZN( u0_u2_u5_n122 ) );
  NAND2_X1 u0_u2_u5_U65 (.A2( u0_u2_u5_n100 ) , .A1( u0_u2_u5_n106 ) , .ZN( u0_u2_u5_n115 ) );
  NAND2_X1 u0_u2_u5_U66 (.A2( u0_u2_u5_n100 ) , .A1( u0_u2_u5_n103 ) , .ZN( u0_u2_u5_n161 ) );
  NAND2_X1 u0_u2_u5_U67 (.A1( u0_u2_u5_n105 ) , .A2( u0_u2_u5_n109 ) , .ZN( u0_u2_u5_n154 ) );
  INV_X1 u0_u2_u5_U68 (.A( u0_u2_u5_n146 ) , .ZN( u0_u2_u5_n172 ) );
  NAND2_X1 u0_u2_u5_U69 (.A1( u0_u2_u5_n103 ) , .A2( u0_u2_u5_n108 ) , .ZN( u0_u2_u5_n123 ) );
  OAI22_X1 u0_u2_u5_U7 (.B2( u0_u2_u5_n149 ) , .B1( u0_u2_u5_n150 ) , .A2( u0_u2_u5_n151 ) , .A1( u0_u2_u5_n152 ) , .ZN( u0_u2_u5_n165 ) );
  NAND2_X1 u0_u2_u5_U70 (.A2( u0_u2_u5_n103 ) , .A1( u0_u2_u5_n107 ) , .ZN( u0_u2_u5_n151 ) );
  NAND2_X1 u0_u2_u5_U71 (.A2( u0_u2_u5_n107 ) , .A1( u0_u2_u5_n109 ) , .ZN( u0_u2_u5_n120 ) );
  NAND2_X1 u0_u2_u5_U72 (.A2( u0_u2_u5_n100 ) , .A1( u0_u2_u5_n109 ) , .ZN( u0_u2_u5_n157 ) );
  AND2_X1 u0_u2_u5_U73 (.A2( u0_u2_u5_n100 ) , .A1( u0_u2_u5_n104 ) , .ZN( u0_u2_u5_n131 ) );
  INV_X1 u0_u2_u5_U74 (.A( u0_u2_u5_n102 ) , .ZN( u0_u2_u5_n195 ) );
  OAI221_X1 u0_u2_u5_U75 (.A( u0_u2_u5_n101 ) , .ZN( u0_u2_u5_n102 ) , .C2( u0_u2_u5_n115 ) , .C1( u0_u2_u5_n126 ) , .B1( u0_u2_u5_n134 ) , .B2( u0_u2_u5_n160 ) );
  OAI21_X1 u0_u2_u5_U76 (.ZN( u0_u2_u5_n101 ) , .B1( u0_u2_u5_n137 ) , .A( u0_u2_u5_n146 ) , .B2( u0_u2_u5_n147 ) );
  NOR2_X1 u0_u2_u5_U77 (.A2( u0_u2_X_34 ) , .A1( u0_u2_X_35 ) , .ZN( u0_u2_u5_n145 ) );
  NOR2_X1 u0_u2_u5_U78 (.A2( u0_u2_X_34 ) , .ZN( u0_u2_u5_n146 ) , .A1( u0_u2_u5_n171 ) );
  NOR2_X1 u0_u2_u5_U79 (.A2( u0_u2_X_31 ) , .A1( u0_u2_X_32 ) , .ZN( u0_u2_u5_n103 ) );
  NOR3_X1 u0_u2_u5_U8 (.A2( u0_u2_u5_n147 ) , .A1( u0_u2_u5_n148 ) , .ZN( u0_u2_u5_n149 ) , .A3( u0_u2_u5_n194 ) );
  NOR2_X1 u0_u2_u5_U80 (.A2( u0_u2_X_36 ) , .ZN( u0_u2_u5_n105 ) , .A1( u0_u2_u5_n180 ) );
  NOR2_X1 u0_u2_u5_U81 (.A2( u0_u2_X_33 ) , .ZN( u0_u2_u5_n108 ) , .A1( u0_u2_u5_n170 ) );
  NOR2_X1 u0_u2_u5_U82 (.A2( u0_u2_X_33 ) , .A1( u0_u2_X_36 ) , .ZN( u0_u2_u5_n107 ) );
  NOR2_X1 u0_u2_u5_U83 (.A2( u0_u2_X_31 ) , .ZN( u0_u2_u5_n104 ) , .A1( u0_u2_u5_n181 ) );
  NAND2_X1 u0_u2_u5_U84 (.A2( u0_u2_X_34 ) , .A1( u0_u2_X_35 ) , .ZN( u0_u2_u5_n153 ) );
  NAND2_X1 u0_u2_u5_U85 (.A1( u0_u2_X_34 ) , .ZN( u0_u2_u5_n126 ) , .A2( u0_u2_u5_n171 ) );
  AND2_X1 u0_u2_u5_U86 (.A1( u0_u2_X_31 ) , .A2( u0_u2_X_32 ) , .ZN( u0_u2_u5_n106 ) );
  AND2_X1 u0_u2_u5_U87 (.A1( u0_u2_X_31 ) , .ZN( u0_u2_u5_n109 ) , .A2( u0_u2_u5_n181 ) );
  INV_X1 u0_u2_u5_U88 (.A( u0_u2_X_33 ) , .ZN( u0_u2_u5_n180 ) );
  INV_X1 u0_u2_u5_U89 (.A( u0_u2_X_35 ) , .ZN( u0_u2_u5_n171 ) );
  NOR2_X1 u0_u2_u5_U9 (.ZN( u0_u2_u5_n135 ) , .A1( u0_u2_u5_n173 ) , .A2( u0_u2_u5_n176 ) );
  INV_X1 u0_u2_u5_U90 (.A( u0_u2_X_36 ) , .ZN( u0_u2_u5_n170 ) );
  INV_X1 u0_u2_u5_U91 (.A( u0_u2_X_32 ) , .ZN( u0_u2_u5_n181 ) );
  NAND4_X1 u0_u2_u5_U92 (.ZN( u0_out2_19 ) , .A4( u0_u2_u5_n166 ) , .A3( u0_u2_u5_n167 ) , .A2( u0_u2_u5_n168 ) , .A1( u0_u2_u5_n169 ) );
  AOI22_X1 u0_u2_u5_U93 (.B2( u0_u2_u5_n145 ) , .A2( u0_u2_u5_n146 ) , .ZN( u0_u2_u5_n167 ) , .B1( u0_u2_u5_n182 ) , .A1( u0_u2_u5_n189 ) );
  NOR4_X1 u0_u2_u5_U94 (.A4( u0_u2_u5_n162 ) , .A3( u0_u2_u5_n163 ) , .A2( u0_u2_u5_n164 ) , .A1( u0_u2_u5_n165 ) , .ZN( u0_u2_u5_n166 ) );
  NAND4_X1 u0_u2_u5_U95 (.ZN( u0_out2_11 ) , .A4( u0_u2_u5_n143 ) , .A3( u0_u2_u5_n144 ) , .A2( u0_u2_u5_n169 ) , .A1( u0_u2_u5_n196 ) );
  AOI22_X1 u0_u2_u5_U96 (.A2( u0_u2_u5_n132 ) , .ZN( u0_u2_u5_n144 ) , .B2( u0_u2_u5_n145 ) , .B1( u0_u2_u5_n184 ) , .A1( u0_u2_u5_n194 ) );
  NOR3_X1 u0_u2_u5_U97 (.A3( u0_u2_u5_n141 ) , .A1( u0_u2_u5_n142 ) , .ZN( u0_u2_u5_n143 ) , .A2( u0_u2_u5_n191 ) );
  NAND4_X1 u0_u2_u5_U98 (.ZN( u0_out2_4 ) , .A4( u0_u2_u5_n112 ) , .A2( u0_u2_u5_n113 ) , .A1( u0_u2_u5_n114 ) , .A3( u0_u2_u5_n195 ) );
  AOI211_X1 u0_u2_u5_U99 (.A( u0_u2_u5_n110 ) , .C1( u0_u2_u5_n111 ) , .ZN( u0_u2_u5_n112 ) , .B( u0_u2_u5_n118 ) , .C2( u0_u2_u5_n177 ) );
  OAI22_X1 u0_uk_U200 (.ZN( u0_K15_24 ) , .A1( u0_uk_n109 ) , .B1( u0_uk_n188 ) , .B2( u0_uk_n24 ) , .A2( u0_uk_n42 ) );
  OAI22_X1 u0_uk_U229 (.ZN( u0_K3_31 ) , .A1( u0_uk_n191 ) , .A2( u0_uk_n549 ) , .B2( u0_uk_n555 ) , .B1( u0_uk_n63 ) );
  OAI22_X1 u0_uk_U319 (.ZN( u0_K3_26 ) , .A1( u0_uk_n109 ) , .B1( u0_uk_n242 ) , .A2( u0_uk_n543 ) , .B2( u0_uk_n559 ) );
  OAI22_X1 u0_uk_U332 (.ZN( u0_K11_4 ) , .A1( u0_uk_n118 ) , .A2( u0_uk_n189 ) , .B2( u0_uk_n195 ) , .B1( u0_uk_n202 ) );
  OAI22_X1 u0_uk_U378 (.ZN( u0_K3_28 ) , .A1( u0_uk_n209 ) , .A2( u0_uk_n555 ) , .B2( u0_uk_n560 ) , .B1( u0_uk_n63 ) );
  OAI22_X1 u0_uk_U388 (.ZN( u0_K11_1 ) , .A2( u0_uk_n183 ) , .B2( u0_uk_n200 ) , .A1( u0_uk_n238 ) , .B1( u0_uk_n93 ) );
  OAI22_X1 u0_uk_U450 (.ZN( u0_K3_33 ) , .A1( u0_uk_n118 ) , .B1( u0_uk_n231 ) , .A2( u0_uk_n549 ) , .B2( u0_uk_n566 ) );
  OAI21_X1 u0_uk_U479 (.ZN( u0_K3_29 ) , .B1( u0_uk_n252 ) , .B2( u0_uk_n545 ) , .A( u0_uk_n849 ) );
  NAND2_X1 u0_uk_U480 (.A1( u0_uk_K_r1_44 ) , .A2( u0_uk_n220 ) , .ZN( u0_uk_n849 ) );
  OAI22_X1 u0_uk_U490 (.ZN( u0_K11_2 ) , .A1( u0_uk_n109 ) , .A2( u0_uk_n181 ) , .B2( u0_uk_n215 ) , .B1( u0_uk_n222 ) );
  OAI22_X1 u0_uk_U547 (.ZN( u0_K3_36 ) , .B1( u0_uk_n231 ) , .A2( u0_uk_n544 ) , .B2( u0_uk_n579 ) , .A1( u0_uk_n94 ) );
  OAI21_X1 u0_uk_U653 (.ZN( u0_K2_43 ) , .B1( u0_uk_n129 ) , .B2( u0_uk_n612 ) , .A( u0_uk_n857 ) );
  NAND2_X1 u0_uk_U654 (.A1( u0_uk_K_r0_2 ) , .A2( u0_uk_n63 ) , .ZN( u0_uk_n857 ) );
  OAI22_X1 u0_uk_U655 (.ZN( u0_K11_3 ) , .A2( u0_uk_n201 ) , .B2( u0_uk_n219 ) , .A1( u0_uk_n222 ) , .B1( u0_uk_n93 ) );
  OAI22_X1 u0_uk_U722 (.ZN( u0_K3_32 ) , .A1( u0_uk_n118 ) , .B1( u0_uk_n148 ) , .A2( u0_uk_n545 ) , .B2( u0_uk_n580 ) );
  OAI22_X1 u0_uk_U768 (.ZN( u0_K15_21 ) , .A1( u0_uk_n164 ) , .B2( u0_uk_n38 ) , .A2( u0_uk_n42 ) , .B1( u0_uk_n92 ) );
  OAI21_X1 u0_uk_U778 (.ZN( u0_K3_27 ) , .B1( u0_uk_n252 ) , .B2( u0_uk_n543 ) , .A( u0_uk_n850 ) );
  NAND2_X1 u0_uk_U779 (.A1( u0_uk_K_r1_42 ) , .A2( u0_uk_n220 ) , .ZN( u0_uk_n850 ) );
  OAI22_X1 u0_uk_U823 (.ZN( u0_K15_20 ) , .B2( u0_uk_n14 ) , .A1( u0_uk_n164 ) , .A2( u0_uk_n43 ) , .B1( u0_uk_n92 ) );
  OAI22_X1 u0_uk_U871 (.ZN( u0_K15_22 ) , .A2( u0_uk_n16 ) , .A1( u0_uk_n188 ) , .B2( u0_uk_n30 ) , .B1( u0_uk_n83 ) );
  OAI22_X1 u0_uk_U873 (.ZN( u0_K15_23 ) , .A1( u0_uk_n187 ) , .B2( u0_uk_n25 ) , .A2( u0_uk_n7 ) , .B1( u0_uk_n83 ) );
  OAI22_X1 u0_uk_U890 (.ZN( u0_K3_30 ) , .A1( u0_uk_n209 ) , .A2( u0_uk_n544 ) , .B2( u0_uk_n570 ) , .B1( u0_uk_n63 ) );
  OAI22_X1 u0_uk_U919 (.ZN( u0_K3_25 ) , .A1( u0_uk_n191 ) , .A2( u0_uk_n575 ) , .B2( u0_uk_n579 ) , .B1( u0_uk_n63 ) );
  INV_X1 u0_uk_U92 (.ZN( u0_K11_5 ) , .A( u0_uk_n984 ) );
  AOI22_X1 u0_uk_U93 (.B2( u0_uk_K_r9_19 ) , .A2( u0_uk_K_r9_25 ) , .B1( u0_uk_n142 ) , .A1( u0_uk_n220 ) , .ZN( u0_uk_n984 ) );
  OAI22_X1 u0_uk_U935 (.ZN( u0_K11_6 ) , .B1( u0_uk_n163 ) , .A2( u0_uk_n183 ) , .B2( u0_uk_n189 ) , .A1( u0_uk_n94 ) );
  OAI22_X1 u0_uk_U962 (.ZN( u0_K15_19 ) , .A1( u0_uk_n141 ) , .B1( u0_uk_n188 ) , .B2( u0_uk_n37 ) , .A2( u0_uk_n7 ) );
  OAI21_X1 u0_uk_U998 (.ZN( u0_K3_35 ) , .B2( u0_uk_n580 ) , .B1( u0_uk_n60 ) , .A( u0_uk_n847 ) );
  NAND2_X1 u0_uk_U999 (.A1( u0_uk_K_r1_7 ) , .A2( u0_uk_n11 ) , .ZN( u0_uk_n847 ) );
  XOR2_X1 u1_U147 (.B( u1_L0_9 ) , .Z( u1_N40 ) , .A( u1_out1_9 ) );
  XOR2_X1 u1_U167 (.B( u1_L10_31 ) , .Z( u1_N382 ) , .A( u1_out11_31 ) );
  XOR2_X1 u1_U176 (.B( u1_L10_23 ) , .Z( u1_N374 ) , .A( u1_out11_23 ) );
  XOR2_X1 u1_U183 (.B( u1_L10_17 ) , .Z( u1_N368 ) , .A( u1_out11_17 ) );
  XOR2_X1 u1_U191 (.B( u1_L10_9 ) , .Z( u1_N360 ) , .A( u1_out11_9 ) );
  XOR2_X1 u1_U201 (.B( u1_L9_32 ) , .Z( u1_N351 ) , .A( u1_out10_32 ) );
  XOR2_X1 u1_U212 (.B( u1_L9_22 ) , .Z( u1_N341 ) , .A( u1_out10_22 ) );
  XOR2_X1 u1_U223 (.B( u1_L9_12 ) , .Z( u1_N331 ) , .A( u1_out10_12 ) );
  XOR2_X1 u1_U229 (.B( u1_L9_7 ) , .Z( u1_N326 ) , .A( u1_out10_7 ) );
  XOR2_X1 u1_U278 (.B( u1_L7_27 ) , .Z( u1_N282 ) , .A( u1_out8_27 ) );
  XOR2_X1 u1_U285 (.B( u1_L7_21 ) , .Z( u1_N276 ) , .A( u1_out8_21 ) );
  XOR2_X1 u1_U291 (.B( u1_L7_15 ) , .Z( u1_N270 ) , .A( u1_out8_15 ) );
  XOR2_X1 u1_U3 (.B( u1_L2_4 ) , .Z( u1_N99 ) , .A( u1_out3_4 ) );
  XOR2_X1 u1_U302 (.B( u1_L7_5 ) , .Z( u1_N260 ) , .A( u1_out8_5 ) );
  XOR2_X1 u1_U309 (.B( u1_L6_31 ) , .Z( u1_N254 ) , .A( u1_out7_31 ) );
  XOR2_X1 u1_U310 (.B( u1_L6_30 ) , .Z( u1_N253 ) , .A( u1_out7_30 ) );
  XOR2_X1 u1_U312 (.B( u1_L6_28 ) , .Z( u1_N251 ) , .A( u1_out7_28 ) );
  XOR2_X1 u1_U317 (.B( u1_L6_24 ) , .Z( u1_N247 ) , .A( u1_out7_24 ) );
  XOR2_X1 u1_U318 (.B( u1_L6_23 ) , .Z( u1_N246 ) , .A( u1_out7_23 ) );
  XOR2_X1 u1_U323 (.B( u1_L6_18 ) , .Z( u1_N241 ) , .A( u1_out7_18 ) );
  XOR2_X1 u1_U324 (.B( u1_L6_17 ) , .Z( u1_N240 ) , .A( u1_out7_17 ) );
  XOR2_X1 u1_U326 (.B( u1_L6_16 ) , .Z( u1_N239 ) , .A( u1_out7_16 ) );
  XOR2_X1 u1_U329 (.B( u1_L6_13 ) , .Z( u1_N236 ) , .A( u1_out7_13 ) );
  XOR2_X1 u1_U333 (.B( u1_L6_9 ) , .Z( u1_N232 ) , .A( u1_out7_9 ) );
  XOR2_X1 u1_U337 (.B( u1_L6_6 ) , .Z( u1_N229 ) , .A( u1_out7_6 ) );
  XOR2_X1 u1_U341 (.B( u1_L6_2 ) , .Z( u1_N225 ) , .A( u1_out7_2 ) );
  XOR2_X1 u1_U343 (.B( u1_L5_32 ) , .Z( u1_N223 ) , .A( u1_out6_32 ) );
  XOR2_X1 u1_U345 (.B( u1_L5_30 ) , .Z( u1_N221 ) , .A( u1_out6_30 ) );
  XOR2_X1 u1_U348 (.B( u1_L5_28 ) , .Z( u1_N219 ) , .A( u1_out6_28 ) );
  XOR2_X1 u1_U349 (.B( u1_L5_27 ) , .Z( u1_N218 ) , .A( u1_out6_27 ) );
  XOR2_X1 u1_U352 (.B( u1_L5_24 ) , .Z( u1_N215 ) , .A( u1_out6_24 ) );
  XOR2_X1 u1_U354 (.B( u1_L5_22 ) , .Z( u1_N213 ) , .A( u1_out6_22 ) );
  XOR2_X1 u1_U355 (.B( u1_L5_21 ) , .Z( u1_N212 ) , .A( u1_out6_21 ) );
  XOR2_X1 u1_U359 (.B( u1_L5_18 ) , .Z( u1_N209 ) , .A( u1_out6_18 ) );
  XOR2_X1 u1_U361 (.B( u1_L5_16 ) , .Z( u1_N207 ) , .A( u1_out6_16 ) );
  XOR2_X1 u1_U362 (.B( u1_L5_15 ) , .Z( u1_N206 ) , .A( u1_out6_15 ) );
  XOR2_X1 u1_U364 (.B( u1_L5_13 ) , .Z( u1_N204 ) , .A( u1_out6_13 ) );
  XOR2_X1 u1_U365 (.B( u1_L5_12 ) , .Z( u1_N203 ) , .A( u1_out6_12 ) );
  XOR2_X1 u1_U372 (.B( u1_L5_7 ) , .Z( u1_N198 ) , .A( u1_out6_7 ) );
  XOR2_X1 u1_U373 (.B( u1_L5_6 ) , .Z( u1_N197 ) , .A( u1_out6_6 ) );
  XOR2_X1 u1_U374 (.B( u1_L5_5 ) , .Z( u1_N196 ) , .A( u1_out6_5 ) );
  XOR2_X1 u1_U377 (.B( u1_L5_2 ) , .Z( u1_N193 ) , .A( u1_out6_2 ) );
  XOR2_X1 u1_U420 (.B( u1_L3_27 ) , .Z( u1_N154 ) , .A( u1_out4_27 ) );
  XOR2_X1 u1_U422 (.B( u1_L3_25 ) , .Z( u1_N152 ) , .A( u1_out4_25 ) );
  XOR2_X1 u1_U427 (.B( u1_L3_21 ) , .Z( u1_N148 ) , .A( u1_out4_21 ) );
  XOR2_X1 u1_U43 (.B( u1_L0_31 ) , .Z( u1_N62 ) , .A( u1_out1_31 ) );
  XOR2_X1 u1_U433 (.B( u1_L3_15 ) , .Z( u1_N142 ) , .A( u1_out4_15 ) );
  XOR2_X1 u1_U434 (.B( u1_L3_14 ) , .Z( u1_N141 ) , .A( u1_out4_14 ) );
  XOR2_X1 u1_U441 (.B( u1_L3_8 ) , .Z( u1_N135 ) , .A( u1_out4_8 ) );
  XOR2_X1 u1_U444 (.B( u1_L3_5 ) , .Z( u1_N132 ) , .A( u1_out4_5 ) );
  XOR2_X1 u1_U446 (.B( u1_L3_3 ) , .Z( u1_N130 ) , .A( u1_out4_3 ) );
  XOR2_X1 u1_U450 (.B( u1_L2_32 ) , .Z( u1_N127 ) , .A( u1_out3_32 ) );
  XOR2_X1 u1_U453 (.B( u1_L2_29 ) , .Z( u1_N124 ) , .A( u1_out3_29 ) );
  XOR2_X1 u1_U461 (.B( u1_L2_22 ) , .Z( u1_N117 ) , .A( u1_out3_22 ) );
  XOR2_X1 u1_U464 (.B( u1_L2_19 ) , .Z( u1_N114 ) , .A( u1_out3_19 ) );
  XOR2_X1 u1_U472 (.B( u1_L2_12 ) , .Z( u1_N107 ) , .A( u1_out3_12 ) );
  XOR2_X1 u1_U473 (.B( u1_L2_11 ) , .Z( u1_N106 ) , .A( u1_out3_11 ) );
  XOR2_X1 u1_U477 (.B( u1_L2_7 ) , .Z( u1_N102 ) , .A( u1_out3_7 ) );
  XOR2_X1 u1_U484 (.Z( u1_FP_8 ) , .B( u1_L14_8 ) , .A( u1_out15_8 ) );
  XOR2_X1 u1_U485 (.Z( u1_FP_7 ) , .B( u1_L14_7 ) , .A( u1_out15_7 ) );
  XOR2_X1 u1_U487 (.Z( u1_FP_5 ) , .B( u1_L14_5 ) , .A( u1_out15_5 ) );
  XOR2_X1 u1_U488 (.Z( u1_FP_4 ) , .B( u1_L14_4 ) , .A( u1_out15_4 ) );
  XOR2_X1 u1_U489 (.Z( u1_FP_3 ) , .B( u1_L14_3 ) , .A( u1_out15_3 ) );
  XOR2_X1 u1_U490 (.Z( u1_FP_32 ) , .B( u1_L14_32 ) , .A( u1_out15_32 ) );
  XOR2_X1 u1_U494 (.Z( u1_FP_29 ) , .B( u1_L14_29 ) , .A( u1_out15_29 ) );
  XOR2_X1 u1_U496 (.Z( u1_FP_27 ) , .B( u1_L14_27 ) , .A( u1_out15_27 ) );
  XOR2_X1 u1_U498 (.Z( u1_FP_25 ) , .B( u1_L14_25 ) , .A( u1_out15_25 ) );
  XOR2_X1 u1_U501 (.Z( u1_FP_22 ) , .B( u1_L14_22 ) , .A( u1_out15_22 ) );
  XOR2_X1 u1_U502 (.Z( u1_FP_21 ) , .B( u1_L14_21 ) , .A( u1_out15_21 ) );
  XOR2_X1 u1_U505 (.Z( u1_FP_19 ) , .B( u1_L14_19 ) , .A( u1_out15_19 ) );
  XOR2_X1 u1_U509 (.Z( u1_FP_15 ) , .B( u1_L14_15 ) , .A( u1_out15_15 ) );
  XOR2_X1 u1_U510 (.Z( u1_FP_14 ) , .B( u1_L14_14 ) , .A( u1_out15_14 ) );
  XOR2_X1 u1_U512 (.Z( u1_FP_12 ) , .B( u1_L14_12 ) , .A( u1_out15_12 ) );
  XOR2_X1 u1_U513 (.Z( u1_FP_11 ) , .B( u1_L14_11 ) , .A( u1_out15_11 ) );
  XOR2_X1 u1_U52 (.B( u1_L0_23 ) , .Z( u1_N54 ) , .A( u1_out1_23 ) );
  XOR2_X1 u1_U59 (.B( u1_L0_17 ) , .Z( u1_N48 ) , .A( u1_out1_17 ) );
  XOR2_X1 u1_U61 (.B( u1_L13_31 ) , .Z( u1_N478 ) , .A( u1_out14_31 ) );
  XOR2_X1 u1_U62 (.B( u1_L13_30 ) , .Z( u1_N477 ) , .A( u1_out14_30 ) );
  XOR2_X1 u1_U64 (.B( u1_L13_28 ) , .Z( u1_N475 ) , .A( u1_out14_28 ) );
  XOR2_X1 u1_U66 (.B( u1_L13_26 ) , .Z( u1_N473 ) , .A( u1_out14_26 ) );
  XOR2_X1 u1_U67 (.B( u1_L13_25 ) , .Z( u1_N472 ) , .A( u1_out14_25 ) );
  XOR2_X1 u1_U68 (.B( u1_L13_24 ) , .Z( u1_N471 ) , .A( u1_out14_24 ) );
  XOR2_X1 u1_U69 (.B( u1_L13_23 ) , .Z( u1_N470 ) , .A( u1_out14_23 ) );
  XOR2_X1 u1_U73 (.B( u1_L13_20 ) , .Z( u1_N467 ) , .A( u1_out14_20 ) );
  XOR2_X1 u1_U75 (.B( u1_L13_18 ) , .Z( u1_N465 ) , .A( u1_out14_18 ) );
  XOR2_X1 u1_U76 (.B( u1_L13_17 ) , .Z( u1_N464 ) , .A( u1_out14_17 ) );
  XOR2_X1 u1_U77 (.B( u1_L13_16 ) , .Z( u1_N463 ) , .A( u1_out14_16 ) );
  XOR2_X1 u1_U79 (.B( u1_L13_14 ) , .Z( u1_N461 ) , .A( u1_out14_14 ) );
  XOR2_X1 u1_U80 (.B( u1_L13_13 ) , .Z( u1_N460 ) , .A( u1_out14_13 ) );
  XOR2_X1 u1_U84 (.B( u1_L13_10 ) , .Z( u1_N457 ) , .A( u1_out14_10 ) );
  XOR2_X1 u1_U85 (.B( u1_L13_9 ) , .Z( u1_N456 ) , .A( u1_out14_9 ) );
  XOR2_X1 u1_U86 (.B( u1_L13_8 ) , .Z( u1_N455 ) , .A( u1_out14_8 ) );
  XOR2_X1 u1_U88 (.B( u1_L13_6 ) , .Z( u1_N453 ) , .A( u1_out14_6 ) );
  XOR2_X1 u1_U91 (.B( u1_L13_3 ) , .Z( u1_N450 ) , .A( u1_out14_3 ) );
  XOR2_X1 u1_U93 (.B( u1_L13_2 ) , .Z( u1_N449 ) , .A( u1_out14_2 ) );
  XOR2_X1 u1_U94 (.B( u1_L13_1 ) , .Z( u1_N448 ) , .A( u1_out14_1 ) );
  XOR2_X1 u1_u10_U13 (.B( u1_K11_42 ) , .A( u1_R9_29 ) , .Z( u1_u10_X_42 ) );
  XOR2_X1 u1_u10_U14 (.B( u1_K11_41 ) , .A( u1_R9_28 ) , .Z( u1_u10_X_41 ) );
  XOR2_X1 u1_u10_U15 (.B( u1_K11_40 ) , .A( u1_R9_27 ) , .Z( u1_u10_X_40 ) );
  XOR2_X1 u1_u10_U17 (.B( u1_K11_39 ) , .A( u1_R9_26 ) , .Z( u1_u10_X_39 ) );
  XOR2_X1 u1_u10_U18 (.B( u1_K11_38 ) , .A( u1_R9_25 ) , .Z( u1_u10_X_38 ) );
  XOR2_X1 u1_u10_U19 (.B( u1_K11_37 ) , .A( u1_R9_24 ) , .Z( u1_u10_X_37 ) );
  AOI22_X1 u1_u10_u6_U10 (.A2( u1_u10_u6_n151 ) , .B2( u1_u10_u6_n161 ) , .A1( u1_u10_u6_n167 ) , .B1( u1_u10_u6_n170 ) , .ZN( u1_u10_u6_n89 ) );
  AOI21_X1 u1_u10_u6_U11 (.B1( u1_u10_u6_n107 ) , .B2( u1_u10_u6_n132 ) , .A( u1_u10_u6_n158 ) , .ZN( u1_u10_u6_n88 ) );
  AOI21_X1 u1_u10_u6_U12 (.B2( u1_u10_u6_n147 ) , .B1( u1_u10_u6_n148 ) , .ZN( u1_u10_u6_n149 ) , .A( u1_u10_u6_n158 ) );
  AOI21_X1 u1_u10_u6_U13 (.ZN( u1_u10_u6_n106 ) , .A( u1_u10_u6_n142 ) , .B2( u1_u10_u6_n159 ) , .B1( u1_u10_u6_n164 ) );
  INV_X1 u1_u10_u6_U14 (.A( u1_u10_u6_n155 ) , .ZN( u1_u10_u6_n161 ) );
  INV_X1 u1_u10_u6_U15 (.A( u1_u10_u6_n128 ) , .ZN( u1_u10_u6_n164 ) );
  NAND2_X1 u1_u10_u6_U16 (.ZN( u1_u10_u6_n110 ) , .A1( u1_u10_u6_n122 ) , .A2( u1_u10_u6_n129 ) );
  NAND2_X1 u1_u10_u6_U17 (.ZN( u1_u10_u6_n124 ) , .A2( u1_u10_u6_n146 ) , .A1( u1_u10_u6_n148 ) );
  INV_X1 u1_u10_u6_U18 (.A( u1_u10_u6_n132 ) , .ZN( u1_u10_u6_n171 ) );
  AND2_X1 u1_u10_u6_U19 (.A1( u1_u10_u6_n100 ) , .ZN( u1_u10_u6_n130 ) , .A2( u1_u10_u6_n147 ) );
  INV_X1 u1_u10_u6_U20 (.A( u1_u10_u6_n127 ) , .ZN( u1_u10_u6_n173 ) );
  INV_X1 u1_u10_u6_U21 (.A( u1_u10_u6_n121 ) , .ZN( u1_u10_u6_n167 ) );
  INV_X1 u1_u10_u6_U22 (.A( u1_u10_u6_n100 ) , .ZN( u1_u10_u6_n169 ) );
  INV_X1 u1_u10_u6_U23 (.A( u1_u10_u6_n123 ) , .ZN( u1_u10_u6_n170 ) );
  INV_X1 u1_u10_u6_U24 (.A( u1_u10_u6_n113 ) , .ZN( u1_u10_u6_n168 ) );
  AND2_X1 u1_u10_u6_U25 (.A1( u1_u10_u6_n107 ) , .A2( u1_u10_u6_n119 ) , .ZN( u1_u10_u6_n133 ) );
  AND2_X1 u1_u10_u6_U26 (.A2( u1_u10_u6_n121 ) , .A1( u1_u10_u6_n122 ) , .ZN( u1_u10_u6_n131 ) );
  AND3_X1 u1_u10_u6_U27 (.ZN( u1_u10_u6_n120 ) , .A2( u1_u10_u6_n127 ) , .A1( u1_u10_u6_n132 ) , .A3( u1_u10_u6_n145 ) );
  INV_X1 u1_u10_u6_U28 (.A( u1_u10_u6_n146 ) , .ZN( u1_u10_u6_n163 ) );
  AOI222_X1 u1_u10_u6_U29 (.ZN( u1_u10_u6_n114 ) , .A1( u1_u10_u6_n118 ) , .A2( u1_u10_u6_n126 ) , .B2( u1_u10_u6_n151 ) , .C2( u1_u10_u6_n159 ) , .C1( u1_u10_u6_n168 ) , .B1( u1_u10_u6_n169 ) );
  INV_X1 u1_u10_u6_U3 (.A( u1_u10_u6_n110 ) , .ZN( u1_u10_u6_n166 ) );
  NOR2_X1 u1_u10_u6_U30 (.A1( u1_u10_u6_n162 ) , .A2( u1_u10_u6_n165 ) , .ZN( u1_u10_u6_n98 ) );
  AOI211_X1 u1_u10_u6_U31 (.B( u1_u10_u6_n134 ) , .A( u1_u10_u6_n135 ) , .C1( u1_u10_u6_n136 ) , .ZN( u1_u10_u6_n137 ) , .C2( u1_u10_u6_n151 ) );
  NAND4_X1 u1_u10_u6_U32 (.A4( u1_u10_u6_n127 ) , .A3( u1_u10_u6_n128 ) , .A2( u1_u10_u6_n129 ) , .A1( u1_u10_u6_n130 ) , .ZN( u1_u10_u6_n136 ) );
  AOI21_X1 u1_u10_u6_U33 (.B2( u1_u10_u6_n132 ) , .B1( u1_u10_u6_n133 ) , .ZN( u1_u10_u6_n134 ) , .A( u1_u10_u6_n158 ) );
  AOI21_X1 u1_u10_u6_U34 (.B1( u1_u10_u6_n131 ) , .ZN( u1_u10_u6_n135 ) , .A( u1_u10_u6_n144 ) , .B2( u1_u10_u6_n146 ) );
  NAND2_X1 u1_u10_u6_U35 (.A1( u1_u10_u6_n144 ) , .ZN( u1_u10_u6_n151 ) , .A2( u1_u10_u6_n158 ) );
  NAND2_X1 u1_u10_u6_U36 (.ZN( u1_u10_u6_n132 ) , .A1( u1_u10_u6_n91 ) , .A2( u1_u10_u6_n97 ) );
  AOI22_X1 u1_u10_u6_U37 (.B2( u1_u10_u6_n110 ) , .B1( u1_u10_u6_n111 ) , .A1( u1_u10_u6_n112 ) , .ZN( u1_u10_u6_n115 ) , .A2( u1_u10_u6_n161 ) );
  NAND4_X1 u1_u10_u6_U38 (.A3( u1_u10_u6_n109 ) , .ZN( u1_u10_u6_n112 ) , .A4( u1_u10_u6_n132 ) , .A2( u1_u10_u6_n147 ) , .A1( u1_u10_u6_n166 ) );
  NOR2_X1 u1_u10_u6_U39 (.ZN( u1_u10_u6_n109 ) , .A1( u1_u10_u6_n170 ) , .A2( u1_u10_u6_n173 ) );
  INV_X1 u1_u10_u6_U4 (.A( u1_u10_u6_n142 ) , .ZN( u1_u10_u6_n174 ) );
  NOR2_X1 u1_u10_u6_U40 (.A2( u1_u10_u6_n126 ) , .ZN( u1_u10_u6_n155 ) , .A1( u1_u10_u6_n160 ) );
  NAND2_X1 u1_u10_u6_U41 (.ZN( u1_u10_u6_n146 ) , .A2( u1_u10_u6_n94 ) , .A1( u1_u10_u6_n99 ) );
  AOI21_X1 u1_u10_u6_U42 (.A( u1_u10_u6_n144 ) , .B2( u1_u10_u6_n145 ) , .B1( u1_u10_u6_n146 ) , .ZN( u1_u10_u6_n150 ) );
  INV_X1 u1_u10_u6_U43 (.A( u1_u10_u6_n111 ) , .ZN( u1_u10_u6_n158 ) );
  NAND2_X1 u1_u10_u6_U44 (.ZN( u1_u10_u6_n127 ) , .A1( u1_u10_u6_n91 ) , .A2( u1_u10_u6_n92 ) );
  NAND2_X1 u1_u10_u6_U45 (.ZN( u1_u10_u6_n129 ) , .A2( u1_u10_u6_n95 ) , .A1( u1_u10_u6_n96 ) );
  INV_X1 u1_u10_u6_U46 (.A( u1_u10_u6_n144 ) , .ZN( u1_u10_u6_n159 ) );
  NAND2_X1 u1_u10_u6_U47 (.ZN( u1_u10_u6_n145 ) , .A2( u1_u10_u6_n97 ) , .A1( u1_u10_u6_n98 ) );
  NAND2_X1 u1_u10_u6_U48 (.ZN( u1_u10_u6_n148 ) , .A2( u1_u10_u6_n92 ) , .A1( u1_u10_u6_n94 ) );
  NAND2_X1 u1_u10_u6_U49 (.ZN( u1_u10_u6_n108 ) , .A2( u1_u10_u6_n139 ) , .A1( u1_u10_u6_n144 ) );
  NAND2_X1 u1_u10_u6_U5 (.A2( u1_u10_u6_n143 ) , .ZN( u1_u10_u6_n152 ) , .A1( u1_u10_u6_n166 ) );
  NAND2_X1 u1_u10_u6_U50 (.ZN( u1_u10_u6_n121 ) , .A2( u1_u10_u6_n95 ) , .A1( u1_u10_u6_n97 ) );
  NAND2_X1 u1_u10_u6_U51 (.ZN( u1_u10_u6_n107 ) , .A2( u1_u10_u6_n92 ) , .A1( u1_u10_u6_n95 ) );
  AND2_X1 u1_u10_u6_U52 (.ZN( u1_u10_u6_n118 ) , .A2( u1_u10_u6_n91 ) , .A1( u1_u10_u6_n99 ) );
  NAND2_X1 u1_u10_u6_U53 (.ZN( u1_u10_u6_n147 ) , .A2( u1_u10_u6_n98 ) , .A1( u1_u10_u6_n99 ) );
  NAND2_X1 u1_u10_u6_U54 (.ZN( u1_u10_u6_n128 ) , .A1( u1_u10_u6_n94 ) , .A2( u1_u10_u6_n96 ) );
  NAND2_X1 u1_u10_u6_U55 (.ZN( u1_u10_u6_n119 ) , .A2( u1_u10_u6_n95 ) , .A1( u1_u10_u6_n99 ) );
  NAND2_X1 u1_u10_u6_U56 (.ZN( u1_u10_u6_n123 ) , .A2( u1_u10_u6_n91 ) , .A1( u1_u10_u6_n96 ) );
  NAND2_X1 u1_u10_u6_U57 (.ZN( u1_u10_u6_n100 ) , .A2( u1_u10_u6_n92 ) , .A1( u1_u10_u6_n98 ) );
  NAND2_X1 u1_u10_u6_U58 (.ZN( u1_u10_u6_n122 ) , .A1( u1_u10_u6_n94 ) , .A2( u1_u10_u6_n97 ) );
  INV_X1 u1_u10_u6_U59 (.A( u1_u10_u6_n139 ) , .ZN( u1_u10_u6_n160 ) );
  AOI22_X1 u1_u10_u6_U6 (.B2( u1_u10_u6_n101 ) , .A1( u1_u10_u6_n102 ) , .ZN( u1_u10_u6_n103 ) , .B1( u1_u10_u6_n160 ) , .A2( u1_u10_u6_n161 ) );
  NAND2_X1 u1_u10_u6_U60 (.ZN( u1_u10_u6_n113 ) , .A1( u1_u10_u6_n96 ) , .A2( u1_u10_u6_n98 ) );
  NOR2_X1 u1_u10_u6_U61 (.A2( u1_u10_X_40 ) , .A1( u1_u10_X_41 ) , .ZN( u1_u10_u6_n126 ) );
  NOR2_X1 u1_u10_u6_U62 (.A2( u1_u10_X_39 ) , .A1( u1_u10_X_42 ) , .ZN( u1_u10_u6_n92 ) );
  NOR2_X1 u1_u10_u6_U63 (.A2( u1_u10_X_39 ) , .A1( u1_u10_u6_n156 ) , .ZN( u1_u10_u6_n97 ) );
  NOR2_X1 u1_u10_u6_U64 (.A2( u1_u10_X_38 ) , .A1( u1_u10_u6_n165 ) , .ZN( u1_u10_u6_n95 ) );
  NOR2_X1 u1_u10_u6_U65 (.A2( u1_u10_X_41 ) , .ZN( u1_u10_u6_n111 ) , .A1( u1_u10_u6_n157 ) );
  NOR2_X1 u1_u10_u6_U66 (.A2( u1_u10_X_37 ) , .A1( u1_u10_u6_n162 ) , .ZN( u1_u10_u6_n94 ) );
  NOR2_X1 u1_u10_u6_U67 (.A2( u1_u10_X_37 ) , .A1( u1_u10_X_38 ) , .ZN( u1_u10_u6_n91 ) );
  NAND2_X1 u1_u10_u6_U68 (.A1( u1_u10_X_41 ) , .ZN( u1_u10_u6_n144 ) , .A2( u1_u10_u6_n157 ) );
  NAND2_X1 u1_u10_u6_U69 (.A2( u1_u10_X_40 ) , .A1( u1_u10_X_41 ) , .ZN( u1_u10_u6_n139 ) );
  NOR2_X1 u1_u10_u6_U7 (.A1( u1_u10_u6_n118 ) , .ZN( u1_u10_u6_n143 ) , .A2( u1_u10_u6_n168 ) );
  AND2_X1 u1_u10_u6_U70 (.A1( u1_u10_X_39 ) , .A2( u1_u10_u6_n156 ) , .ZN( u1_u10_u6_n96 ) );
  AND2_X1 u1_u10_u6_U71 (.A1( u1_u10_X_39 ) , .A2( u1_u10_X_42 ) , .ZN( u1_u10_u6_n99 ) );
  INV_X1 u1_u10_u6_U72 (.A( u1_u10_X_40 ) , .ZN( u1_u10_u6_n157 ) );
  INV_X1 u1_u10_u6_U73 (.A( u1_u10_X_37 ) , .ZN( u1_u10_u6_n165 ) );
  INV_X1 u1_u10_u6_U74 (.A( u1_u10_X_38 ) , .ZN( u1_u10_u6_n162 ) );
  INV_X1 u1_u10_u6_U75 (.A( u1_u10_X_42 ) , .ZN( u1_u10_u6_n156 ) );
  NAND4_X1 u1_u10_u6_U76 (.ZN( u1_out10_32 ) , .A4( u1_u10_u6_n103 ) , .A3( u1_u10_u6_n104 ) , .A2( u1_u10_u6_n105 ) , .A1( u1_u10_u6_n106 ) );
  AOI22_X1 u1_u10_u6_U77 (.ZN( u1_u10_u6_n105 ) , .A2( u1_u10_u6_n108 ) , .A1( u1_u10_u6_n118 ) , .B2( u1_u10_u6_n126 ) , .B1( u1_u10_u6_n171 ) );
  AOI22_X1 u1_u10_u6_U78 (.ZN( u1_u10_u6_n104 ) , .A1( u1_u10_u6_n111 ) , .B1( u1_u10_u6_n124 ) , .B2( u1_u10_u6_n151 ) , .A2( u1_u10_u6_n93 ) );
  NAND4_X1 u1_u10_u6_U79 (.ZN( u1_out10_12 ) , .A4( u1_u10_u6_n114 ) , .A3( u1_u10_u6_n115 ) , .A2( u1_u10_u6_n116 ) , .A1( u1_u10_u6_n117 ) );
  INV_X1 u1_u10_u6_U8 (.ZN( u1_u10_u6_n172 ) , .A( u1_u10_u6_n88 ) );
  OAI22_X1 u1_u10_u6_U80 (.B2( u1_u10_u6_n111 ) , .ZN( u1_u10_u6_n116 ) , .B1( u1_u10_u6_n126 ) , .A2( u1_u10_u6_n164 ) , .A1( u1_u10_u6_n167 ) );
  OAI21_X1 u1_u10_u6_U81 (.A( u1_u10_u6_n108 ) , .ZN( u1_u10_u6_n117 ) , .B2( u1_u10_u6_n141 ) , .B1( u1_u10_u6_n163 ) );
  OAI211_X1 u1_u10_u6_U82 (.ZN( u1_out10_7 ) , .B( u1_u10_u6_n153 ) , .C2( u1_u10_u6_n154 ) , .C1( u1_u10_u6_n155 ) , .A( u1_u10_u6_n174 ) );
  NOR3_X1 u1_u10_u6_U83 (.A1( u1_u10_u6_n141 ) , .ZN( u1_u10_u6_n154 ) , .A3( u1_u10_u6_n164 ) , .A2( u1_u10_u6_n171 ) );
  AOI211_X1 u1_u10_u6_U84 (.B( u1_u10_u6_n149 ) , .A( u1_u10_u6_n150 ) , .C2( u1_u10_u6_n151 ) , .C1( u1_u10_u6_n152 ) , .ZN( u1_u10_u6_n153 ) );
  OAI211_X1 u1_u10_u6_U85 (.ZN( u1_out10_22 ) , .B( u1_u10_u6_n137 ) , .A( u1_u10_u6_n138 ) , .C2( u1_u10_u6_n139 ) , .C1( u1_u10_u6_n140 ) );
  AOI22_X1 u1_u10_u6_U86 (.B1( u1_u10_u6_n124 ) , .A2( u1_u10_u6_n125 ) , .A1( u1_u10_u6_n126 ) , .ZN( u1_u10_u6_n138 ) , .B2( u1_u10_u6_n161 ) );
  AND4_X1 u1_u10_u6_U87 (.A3( u1_u10_u6_n119 ) , .A1( u1_u10_u6_n120 ) , .A4( u1_u10_u6_n129 ) , .ZN( u1_u10_u6_n140 ) , .A2( u1_u10_u6_n143 ) );
  NAND3_X1 u1_u10_u6_U88 (.A2( u1_u10_u6_n123 ) , .ZN( u1_u10_u6_n125 ) , .A1( u1_u10_u6_n130 ) , .A3( u1_u10_u6_n131 ) );
  NAND3_X1 u1_u10_u6_U89 (.A3( u1_u10_u6_n133 ) , .ZN( u1_u10_u6_n141 ) , .A1( u1_u10_u6_n145 ) , .A2( u1_u10_u6_n148 ) );
  OAI21_X1 u1_u10_u6_U9 (.A( u1_u10_u6_n159 ) , .B1( u1_u10_u6_n169 ) , .B2( u1_u10_u6_n173 ) , .ZN( u1_u10_u6_n90 ) );
  NAND3_X1 u1_u10_u6_U90 (.ZN( u1_u10_u6_n101 ) , .A3( u1_u10_u6_n107 ) , .A2( u1_u10_u6_n121 ) , .A1( u1_u10_u6_n127 ) );
  NAND3_X1 u1_u10_u6_U91 (.ZN( u1_u10_u6_n102 ) , .A3( u1_u10_u6_n130 ) , .A2( u1_u10_u6_n145 ) , .A1( u1_u10_u6_n166 ) );
  NAND3_X1 u1_u10_u6_U92 (.A3( u1_u10_u6_n113 ) , .A1( u1_u10_u6_n119 ) , .A2( u1_u10_u6_n123 ) , .ZN( u1_u10_u6_n93 ) );
  NAND3_X1 u1_u10_u6_U93 (.ZN( u1_u10_u6_n142 ) , .A2( u1_u10_u6_n172 ) , .A3( u1_u10_u6_n89 ) , .A1( u1_u10_u6_n90 ) );
  XOR2_X1 u1_u11_U16 (.B( u1_K12_3 ) , .A( u1_R10_2 ) , .Z( u1_u11_X_3 ) );
  XOR2_X1 u1_u11_U27 (.B( u1_K12_2 ) , .A( u1_R10_1 ) , .Z( u1_u11_X_2 ) );
  XOR2_X1 u1_u11_U38 (.B( u1_K12_1 ) , .A( u1_R10_32 ) , .Z( u1_u11_X_1 ) );
  XOR2_X1 u1_u11_U4 (.B( u1_K12_6 ) , .A( u1_R10_5 ) , .Z( u1_u11_X_6 ) );
  XOR2_X1 u1_u11_U5 (.B( u1_K12_5 ) , .A( u1_R10_4 ) , .Z( u1_u11_X_5 ) );
  XOR2_X1 u1_u11_U6 (.B( u1_K12_4 ) , .A( u1_R10_3 ) , .Z( u1_u11_X_4 ) );
  NAND2_X1 u1_u11_u0_U10 (.ZN( u1_u11_u0_n113 ) , .A1( u1_u11_u0_n139 ) , .A2( u1_u11_u0_n149 ) );
  AND3_X1 u1_u11_u0_U11 (.A2( u1_u11_u0_n112 ) , .ZN( u1_u11_u0_n127 ) , .A3( u1_u11_u0_n130 ) , .A1( u1_u11_u0_n148 ) );
  AND2_X1 u1_u11_u0_U12 (.ZN( u1_u11_u0_n107 ) , .A1( u1_u11_u0_n130 ) , .A2( u1_u11_u0_n140 ) );
  AND2_X1 u1_u11_u0_U13 (.A2( u1_u11_u0_n129 ) , .A1( u1_u11_u0_n130 ) , .ZN( u1_u11_u0_n151 ) );
  AND2_X1 u1_u11_u0_U14 (.A1( u1_u11_u0_n108 ) , .A2( u1_u11_u0_n125 ) , .ZN( u1_u11_u0_n145 ) );
  INV_X1 u1_u11_u0_U15 (.A( u1_u11_u0_n143 ) , .ZN( u1_u11_u0_n173 ) );
  NOR2_X1 u1_u11_u0_U16 (.A2( u1_u11_u0_n136 ) , .ZN( u1_u11_u0_n147 ) , .A1( u1_u11_u0_n160 ) );
  OAI22_X1 u1_u11_u0_U17 (.B1( u1_u11_u0_n131 ) , .A1( u1_u11_u0_n144 ) , .B2( u1_u11_u0_n147 ) , .A2( u1_u11_u0_n90 ) , .ZN( u1_u11_u0_n91 ) );
  AND3_X1 u1_u11_u0_U18 (.A3( u1_u11_u0_n121 ) , .A2( u1_u11_u0_n125 ) , .A1( u1_u11_u0_n148 ) , .ZN( u1_u11_u0_n90 ) );
  OAI22_X1 u1_u11_u0_U19 (.B1( u1_u11_u0_n125 ) , .ZN( u1_u11_u0_n126 ) , .A1( u1_u11_u0_n138 ) , .A2( u1_u11_u0_n146 ) , .B2( u1_u11_u0_n147 ) );
  NOR2_X1 u1_u11_u0_U20 (.A1( u1_u11_u0_n163 ) , .A2( u1_u11_u0_n164 ) , .ZN( u1_u11_u0_n95 ) );
  NAND2_X1 u1_u11_u0_U21 (.A1( u1_u11_u0_n101 ) , .A2( u1_u11_u0_n102 ) , .ZN( u1_u11_u0_n150 ) );
  AOI22_X1 u1_u11_u0_U22 (.B2( u1_u11_u0_n109 ) , .A2( u1_u11_u0_n110 ) , .ZN( u1_u11_u0_n111 ) , .B1( u1_u11_u0_n118 ) , .A1( u1_u11_u0_n160 ) );
  INV_X1 u1_u11_u0_U23 (.A( u1_u11_u0_n136 ) , .ZN( u1_u11_u0_n161 ) );
  INV_X1 u1_u11_u0_U24 (.A( u1_u11_u0_n118 ) , .ZN( u1_u11_u0_n158 ) );
  NAND2_X1 u1_u11_u0_U25 (.A2( u1_u11_u0_n100 ) , .A1( u1_u11_u0_n101 ) , .ZN( u1_u11_u0_n139 ) );
  NAND2_X1 u1_u11_u0_U26 (.A2( u1_u11_u0_n100 ) , .ZN( u1_u11_u0_n131 ) , .A1( u1_u11_u0_n92 ) );
  NAND2_X1 u1_u11_u0_U27 (.ZN( u1_u11_u0_n108 ) , .A1( u1_u11_u0_n92 ) , .A2( u1_u11_u0_n94 ) );
  AOI21_X1 u1_u11_u0_U28 (.ZN( u1_u11_u0_n104 ) , .B1( u1_u11_u0_n107 ) , .B2( u1_u11_u0_n141 ) , .A( u1_u11_u0_n144 ) );
  AOI21_X1 u1_u11_u0_U29 (.B1( u1_u11_u0_n127 ) , .B2( u1_u11_u0_n129 ) , .A( u1_u11_u0_n138 ) , .ZN( u1_u11_u0_n96 ) );
  INV_X1 u1_u11_u0_U3 (.A( u1_u11_u0_n113 ) , .ZN( u1_u11_u0_n166 ) );
  NAND2_X1 u1_u11_u0_U30 (.A2( u1_u11_u0_n102 ) , .ZN( u1_u11_u0_n114 ) , .A1( u1_u11_u0_n92 ) );
  NAND2_X1 u1_u11_u0_U31 (.A1( u1_u11_u0_n101 ) , .ZN( u1_u11_u0_n130 ) , .A2( u1_u11_u0_n94 ) );
  NOR2_X1 u1_u11_u0_U32 (.A1( u1_u11_u0_n120 ) , .ZN( u1_u11_u0_n143 ) , .A2( u1_u11_u0_n167 ) );
  OAI221_X1 u1_u11_u0_U33 (.C1( u1_u11_u0_n112 ) , .ZN( u1_u11_u0_n120 ) , .B1( u1_u11_u0_n138 ) , .B2( u1_u11_u0_n141 ) , .C2( u1_u11_u0_n147 ) , .A( u1_u11_u0_n172 ) );
  AOI211_X1 u1_u11_u0_U34 (.B( u1_u11_u0_n115 ) , .A( u1_u11_u0_n116 ) , .C2( u1_u11_u0_n117 ) , .C1( u1_u11_u0_n118 ) , .ZN( u1_u11_u0_n119 ) );
  NAND2_X1 u1_u11_u0_U35 (.A1( u1_u11_u0_n100 ) , .A2( u1_u11_u0_n103 ) , .ZN( u1_u11_u0_n125 ) );
  NAND2_X1 u1_u11_u0_U36 (.A2( u1_u11_u0_n103 ) , .ZN( u1_u11_u0_n140 ) , .A1( u1_u11_u0_n94 ) );
  INV_X1 u1_u11_u0_U37 (.A( u1_u11_u0_n138 ) , .ZN( u1_u11_u0_n160 ) );
  NAND2_X1 u1_u11_u0_U38 (.A2( u1_u11_u0_n102 ) , .A1( u1_u11_u0_n103 ) , .ZN( u1_u11_u0_n149 ) );
  NAND2_X1 u1_u11_u0_U39 (.A2( u1_u11_u0_n101 ) , .ZN( u1_u11_u0_n121 ) , .A1( u1_u11_u0_n93 ) );
  AOI21_X1 u1_u11_u0_U4 (.B1( u1_u11_u0_n114 ) , .ZN( u1_u11_u0_n115 ) , .B2( u1_u11_u0_n129 ) , .A( u1_u11_u0_n161 ) );
  NAND2_X1 u1_u11_u0_U40 (.ZN( u1_u11_u0_n112 ) , .A2( u1_u11_u0_n92 ) , .A1( u1_u11_u0_n93 ) );
  INV_X1 u1_u11_u0_U41 (.ZN( u1_u11_u0_n172 ) , .A( u1_u11_u0_n88 ) );
  OAI222_X1 u1_u11_u0_U42 (.C1( u1_u11_u0_n108 ) , .A1( u1_u11_u0_n125 ) , .B2( u1_u11_u0_n128 ) , .B1( u1_u11_u0_n144 ) , .A2( u1_u11_u0_n158 ) , .C2( u1_u11_u0_n161 ) , .ZN( u1_u11_u0_n88 ) );
  AOI21_X1 u1_u11_u0_U43 (.B1( u1_u11_u0_n103 ) , .ZN( u1_u11_u0_n132 ) , .A( u1_u11_u0_n165 ) , .B2( u1_u11_u0_n93 ) );
  OR3_X1 u1_u11_u0_U44 (.A3( u1_u11_u0_n152 ) , .A2( u1_u11_u0_n153 ) , .A1( u1_u11_u0_n154 ) , .ZN( u1_u11_u0_n155 ) );
  AOI21_X1 u1_u11_u0_U45 (.A( u1_u11_u0_n144 ) , .B2( u1_u11_u0_n145 ) , .B1( u1_u11_u0_n146 ) , .ZN( u1_u11_u0_n154 ) );
  AOI21_X1 u1_u11_u0_U46 (.B2( u1_u11_u0_n150 ) , .B1( u1_u11_u0_n151 ) , .ZN( u1_u11_u0_n152 ) , .A( u1_u11_u0_n158 ) );
  AOI21_X1 u1_u11_u0_U47 (.A( u1_u11_u0_n147 ) , .B2( u1_u11_u0_n148 ) , .B1( u1_u11_u0_n149 ) , .ZN( u1_u11_u0_n153 ) );
  INV_X1 u1_u11_u0_U48 (.ZN( u1_u11_u0_n171 ) , .A( u1_u11_u0_n99 ) );
  OAI211_X1 u1_u11_u0_U49 (.C2( u1_u11_u0_n140 ) , .C1( u1_u11_u0_n161 ) , .A( u1_u11_u0_n169 ) , .B( u1_u11_u0_n98 ) , .ZN( u1_u11_u0_n99 ) );
  AOI21_X1 u1_u11_u0_U5 (.B2( u1_u11_u0_n131 ) , .ZN( u1_u11_u0_n134 ) , .B1( u1_u11_u0_n151 ) , .A( u1_u11_u0_n158 ) );
  AOI211_X1 u1_u11_u0_U50 (.C1( u1_u11_u0_n118 ) , .A( u1_u11_u0_n123 ) , .B( u1_u11_u0_n96 ) , .C2( u1_u11_u0_n97 ) , .ZN( u1_u11_u0_n98 ) );
  INV_X1 u1_u11_u0_U51 (.ZN( u1_u11_u0_n169 ) , .A( u1_u11_u0_n91 ) );
  NOR2_X1 u1_u11_u0_U52 (.A2( u1_u11_X_2 ) , .ZN( u1_u11_u0_n103 ) , .A1( u1_u11_u0_n164 ) );
  NOR2_X1 u1_u11_u0_U53 (.A2( u1_u11_X_4 ) , .A1( u1_u11_X_5 ) , .ZN( u1_u11_u0_n118 ) );
  NOR2_X1 u1_u11_u0_U54 (.A2( u1_u11_X_3 ) , .A1( u1_u11_X_6 ) , .ZN( u1_u11_u0_n94 ) );
  NOR2_X1 u1_u11_u0_U55 (.A2( u1_u11_X_6 ) , .ZN( u1_u11_u0_n100 ) , .A1( u1_u11_u0_n162 ) );
  NAND2_X1 u1_u11_u0_U56 (.A2( u1_u11_X_4 ) , .A1( u1_u11_X_5 ) , .ZN( u1_u11_u0_n144 ) );
  NOR2_X1 u1_u11_u0_U57 (.A2( u1_u11_X_5 ) , .ZN( u1_u11_u0_n136 ) , .A1( u1_u11_u0_n159 ) );
  NAND2_X1 u1_u11_u0_U58 (.A1( u1_u11_X_5 ) , .ZN( u1_u11_u0_n138 ) , .A2( u1_u11_u0_n159 ) );
  AND2_X1 u1_u11_u0_U59 (.A2( u1_u11_X_3 ) , .A1( u1_u11_X_6 ) , .ZN( u1_u11_u0_n102 ) );
  NOR2_X1 u1_u11_u0_U6 (.A1( u1_u11_u0_n108 ) , .ZN( u1_u11_u0_n123 ) , .A2( u1_u11_u0_n158 ) );
  AND2_X1 u1_u11_u0_U60 (.A1( u1_u11_X_6 ) , .A2( u1_u11_u0_n162 ) , .ZN( u1_u11_u0_n93 ) );
  INV_X1 u1_u11_u0_U61 (.A( u1_u11_X_4 ) , .ZN( u1_u11_u0_n159 ) );
  INV_X1 u1_u11_u0_U62 (.A( u1_u11_X_3 ) , .ZN( u1_u11_u0_n162 ) );
  INV_X1 u1_u11_u0_U63 (.A( u1_u11_X_2 ) , .ZN( u1_u11_u0_n163 ) );
  AOI211_X1 u1_u11_u0_U64 (.B( u1_u11_u0_n133 ) , .A( u1_u11_u0_n134 ) , .C2( u1_u11_u0_n135 ) , .C1( u1_u11_u0_n136 ) , .ZN( u1_u11_u0_n137 ) );
  INV_X1 u1_u11_u0_U65 (.A( u1_u11_u0_n126 ) , .ZN( u1_u11_u0_n168 ) );
  OR4_X1 u1_u11_u0_U66 (.ZN( u1_out11_17 ) , .A4( u1_u11_u0_n122 ) , .A2( u1_u11_u0_n123 ) , .A1( u1_u11_u0_n124 ) , .A3( u1_u11_u0_n170 ) );
  AOI21_X1 u1_u11_u0_U67 (.B2( u1_u11_u0_n107 ) , .ZN( u1_u11_u0_n124 ) , .B1( u1_u11_u0_n128 ) , .A( u1_u11_u0_n161 ) );
  INV_X1 u1_u11_u0_U68 (.A( u1_u11_u0_n111 ) , .ZN( u1_u11_u0_n170 ) );
  OR4_X1 u1_u11_u0_U69 (.ZN( u1_out11_31 ) , .A4( u1_u11_u0_n155 ) , .A2( u1_u11_u0_n156 ) , .A1( u1_u11_u0_n157 ) , .A3( u1_u11_u0_n173 ) );
  OAI21_X1 u1_u11_u0_U7 (.B1( u1_u11_u0_n150 ) , .B2( u1_u11_u0_n158 ) , .A( u1_u11_u0_n172 ) , .ZN( u1_u11_u0_n89 ) );
  AOI21_X1 u1_u11_u0_U70 (.A( u1_u11_u0_n138 ) , .B2( u1_u11_u0_n139 ) , .B1( u1_u11_u0_n140 ) , .ZN( u1_u11_u0_n157 ) );
  INV_X1 u1_u11_u0_U71 (.ZN( u1_u11_u0_n174 ) , .A( u1_u11_u0_n89 ) );
  AOI211_X1 u1_u11_u0_U72 (.B( u1_u11_u0_n104 ) , .A( u1_u11_u0_n105 ) , .ZN( u1_u11_u0_n106 ) , .C2( u1_u11_u0_n113 ) , .C1( u1_u11_u0_n160 ) );
  AOI21_X1 u1_u11_u0_U73 (.B2( u1_u11_u0_n141 ) , .B1( u1_u11_u0_n142 ) , .ZN( u1_u11_u0_n156 ) , .A( u1_u11_u0_n161 ) );
  AOI21_X1 u1_u11_u0_U74 (.ZN( u1_u11_u0_n116 ) , .B2( u1_u11_u0_n142 ) , .A( u1_u11_u0_n144 ) , .B1( u1_u11_u0_n166 ) );
  INV_X1 u1_u11_u0_U75 (.A( u1_u11_u0_n142 ) , .ZN( u1_u11_u0_n165 ) );
  NOR2_X1 u1_u11_u0_U76 (.A2( u1_u11_X_1 ) , .A1( u1_u11_X_2 ) , .ZN( u1_u11_u0_n92 ) );
  NOR2_X1 u1_u11_u0_U77 (.A2( u1_u11_X_1 ) , .ZN( u1_u11_u0_n101 ) , .A1( u1_u11_u0_n163 ) );
  INV_X1 u1_u11_u0_U78 (.A( u1_u11_X_1 ) , .ZN( u1_u11_u0_n164 ) );
  OAI221_X1 u1_u11_u0_U79 (.C1( u1_u11_u0_n121 ) , .ZN( u1_u11_u0_n122 ) , .B2( u1_u11_u0_n127 ) , .A( u1_u11_u0_n143 ) , .B1( u1_u11_u0_n144 ) , .C2( u1_u11_u0_n147 ) );
  AND2_X1 u1_u11_u0_U8 (.A1( u1_u11_u0_n114 ) , .A2( u1_u11_u0_n121 ) , .ZN( u1_u11_u0_n146 ) );
  AOI21_X1 u1_u11_u0_U80 (.B1( u1_u11_u0_n132 ) , .ZN( u1_u11_u0_n133 ) , .A( u1_u11_u0_n144 ) , .B2( u1_u11_u0_n166 ) );
  OAI22_X1 u1_u11_u0_U81 (.ZN( u1_u11_u0_n105 ) , .A2( u1_u11_u0_n132 ) , .B1( u1_u11_u0_n146 ) , .A1( u1_u11_u0_n147 ) , .B2( u1_u11_u0_n161 ) );
  NAND2_X1 u1_u11_u0_U82 (.ZN( u1_u11_u0_n110 ) , .A2( u1_u11_u0_n132 ) , .A1( u1_u11_u0_n145 ) );
  INV_X1 u1_u11_u0_U83 (.A( u1_u11_u0_n119 ) , .ZN( u1_u11_u0_n167 ) );
  NAND2_X1 u1_u11_u0_U84 (.ZN( u1_u11_u0_n148 ) , .A1( u1_u11_u0_n93 ) , .A2( u1_u11_u0_n95 ) );
  NAND2_X1 u1_u11_u0_U85 (.A1( u1_u11_u0_n100 ) , .ZN( u1_u11_u0_n129 ) , .A2( u1_u11_u0_n95 ) );
  NAND2_X1 u1_u11_u0_U86 (.A1( u1_u11_u0_n102 ) , .ZN( u1_u11_u0_n128 ) , .A2( u1_u11_u0_n95 ) );
  NAND2_X1 u1_u11_u0_U87 (.ZN( u1_u11_u0_n142 ) , .A1( u1_u11_u0_n94 ) , .A2( u1_u11_u0_n95 ) );
  NAND3_X1 u1_u11_u0_U88 (.ZN( u1_out11_23 ) , .A3( u1_u11_u0_n137 ) , .A1( u1_u11_u0_n168 ) , .A2( u1_u11_u0_n171 ) );
  NAND3_X1 u1_u11_u0_U89 (.A3( u1_u11_u0_n127 ) , .A2( u1_u11_u0_n128 ) , .ZN( u1_u11_u0_n135 ) , .A1( u1_u11_u0_n150 ) );
  AND2_X1 u1_u11_u0_U9 (.A1( u1_u11_u0_n131 ) , .ZN( u1_u11_u0_n141 ) , .A2( u1_u11_u0_n150 ) );
  NAND3_X1 u1_u11_u0_U90 (.ZN( u1_u11_u0_n117 ) , .A3( u1_u11_u0_n132 ) , .A2( u1_u11_u0_n139 ) , .A1( u1_u11_u0_n148 ) );
  NAND3_X1 u1_u11_u0_U91 (.ZN( u1_u11_u0_n109 ) , .A2( u1_u11_u0_n114 ) , .A3( u1_u11_u0_n140 ) , .A1( u1_u11_u0_n149 ) );
  NAND3_X1 u1_u11_u0_U92 (.ZN( u1_out11_9 ) , .A3( u1_u11_u0_n106 ) , .A2( u1_u11_u0_n171 ) , .A1( u1_u11_u0_n174 ) );
  NAND3_X1 u1_u11_u0_U93 (.A2( u1_u11_u0_n128 ) , .A1( u1_u11_u0_n132 ) , .A3( u1_u11_u0_n146 ) , .ZN( u1_u11_u0_n97 ) );
  XOR2_X1 u1_u14_U1 (.B( u1_K15_9 ) , .A( u1_R13_6 ) , .Z( u1_u14_X_9 ) );
  XOR2_X1 u1_u14_U16 (.B( u1_K15_3 ) , .A( u1_R13_2 ) , .Z( u1_u14_X_3 ) );
  XOR2_X1 u1_u14_U2 (.B( u1_K15_8 ) , .A( u1_R13_5 ) , .Z( u1_u14_X_8 ) );
  XOR2_X1 u1_u14_U26 (.B( u1_K15_30 ) , .A( u1_R13_21 ) , .Z( u1_u14_X_30 ) );
  XOR2_X1 u1_u14_U27 (.B( u1_K15_2 ) , .A( u1_R13_1 ) , .Z( u1_u14_X_2 ) );
  XOR2_X1 u1_u14_U28 (.B( u1_K15_29 ) , .A( u1_R13_20 ) , .Z( u1_u14_X_29 ) );
  XOR2_X1 u1_u14_U29 (.B( u1_K15_28 ) , .A( u1_R13_19 ) , .Z( u1_u14_X_28 ) );
  XOR2_X1 u1_u14_U3 (.B( u1_K15_7 ) , .A( u1_R13_4 ) , .Z( u1_u14_X_7 ) );
  XOR2_X1 u1_u14_U30 (.B( u1_K15_27 ) , .A( u1_R13_18 ) , .Z( u1_u14_X_27 ) );
  XOR2_X1 u1_u14_U31 (.B( u1_K15_26 ) , .A( u1_R13_17 ) , .Z( u1_u14_X_26 ) );
  XOR2_X1 u1_u14_U32 (.B( u1_K15_25 ) , .A( u1_R13_16 ) , .Z( u1_u14_X_25 ) );
  XOR2_X1 u1_u14_U33 (.B( u1_K15_24 ) , .A( u1_R13_17 ) , .Z( u1_u14_X_24 ) );
  XOR2_X1 u1_u14_U34 (.B( u1_K15_23 ) , .A( u1_R13_16 ) , .Z( u1_u14_X_23 ) );
  XOR2_X1 u1_u14_U35 (.B( u1_K15_22 ) , .A( u1_R13_15 ) , .Z( u1_u14_X_22 ) );
  XOR2_X1 u1_u14_U36 (.B( u1_K15_21 ) , .A( u1_R13_14 ) , .Z( u1_u14_X_21 ) );
  XOR2_X1 u1_u14_U37 (.B( u1_K15_20 ) , .A( u1_R13_13 ) , .Z( u1_u14_X_20 ) );
  XOR2_X1 u1_u14_U38 (.B( u1_K15_1 ) , .A( u1_R13_32 ) , .Z( u1_u14_X_1 ) );
  XOR2_X1 u1_u14_U39 (.B( u1_K15_19 ) , .A( u1_R13_12 ) , .Z( u1_u14_X_19 ) );
  XOR2_X1 u1_u14_U4 (.B( u1_K15_6 ) , .A( u1_R13_5 ) , .Z( u1_u14_X_6 ) );
  XOR2_X1 u1_u14_U40 (.B( u1_K15_18 ) , .A( u1_R13_13 ) , .Z( u1_u14_X_18 ) );
  XOR2_X1 u1_u14_U41 (.B( u1_K15_17 ) , .A( u1_R13_12 ) , .Z( u1_u14_X_17 ) );
  XOR2_X1 u1_u14_U42 (.B( u1_K15_16 ) , .A( u1_R13_11 ) , .Z( u1_u14_X_16 ) );
  XOR2_X1 u1_u14_U43 (.B( u1_K15_15 ) , .A( u1_R13_10 ) , .Z( u1_u14_X_15 ) );
  XOR2_X1 u1_u14_U44 (.B( u1_K15_14 ) , .A( u1_R13_9 ) , .Z( u1_u14_X_14 ) );
  XOR2_X1 u1_u14_U45 (.B( u1_K15_13 ) , .A( u1_R13_8 ) , .Z( u1_u14_X_13 ) );
  XOR2_X1 u1_u14_U46 (.B( u1_K15_12 ) , .A( u1_R13_9 ) , .Z( u1_u14_X_12 ) );
  XOR2_X1 u1_u14_U47 (.B( u1_K15_11 ) , .A( u1_R13_8 ) , .Z( u1_u14_X_11 ) );
  XOR2_X1 u1_u14_U48 (.B( u1_K15_10 ) , .A( u1_R13_7 ) , .Z( u1_u14_X_10 ) );
  XOR2_X1 u1_u14_U5 (.B( u1_K15_5 ) , .A( u1_R13_4 ) , .Z( u1_u14_X_5 ) );
  XOR2_X1 u1_u14_U6 (.B( u1_K15_4 ) , .A( u1_R13_3 ) , .Z( u1_u14_X_4 ) );
  AND3_X1 u1_u14_u0_U10 (.A2( u1_u14_u0_n112 ) , .ZN( u1_u14_u0_n127 ) , .A3( u1_u14_u0_n130 ) , .A1( u1_u14_u0_n148 ) );
  NAND2_X1 u1_u14_u0_U11 (.ZN( u1_u14_u0_n113 ) , .A1( u1_u14_u0_n139 ) , .A2( u1_u14_u0_n149 ) );
  AND2_X1 u1_u14_u0_U12 (.ZN( u1_u14_u0_n107 ) , .A1( u1_u14_u0_n130 ) , .A2( u1_u14_u0_n140 ) );
  AND2_X1 u1_u14_u0_U13 (.A2( u1_u14_u0_n129 ) , .A1( u1_u14_u0_n130 ) , .ZN( u1_u14_u0_n151 ) );
  AND2_X1 u1_u14_u0_U14 (.A1( u1_u14_u0_n108 ) , .A2( u1_u14_u0_n125 ) , .ZN( u1_u14_u0_n145 ) );
  INV_X1 u1_u14_u0_U15 (.A( u1_u14_u0_n143 ) , .ZN( u1_u14_u0_n173 ) );
  NOR2_X1 u1_u14_u0_U16 (.A2( u1_u14_u0_n136 ) , .ZN( u1_u14_u0_n147 ) , .A1( u1_u14_u0_n160 ) );
  NOR2_X1 u1_u14_u0_U17 (.A1( u1_u14_u0_n163 ) , .A2( u1_u14_u0_n164 ) , .ZN( u1_u14_u0_n95 ) );
  AOI21_X1 u1_u14_u0_U18 (.B1( u1_u14_u0_n103 ) , .ZN( u1_u14_u0_n132 ) , .A( u1_u14_u0_n165 ) , .B2( u1_u14_u0_n93 ) );
  INV_X1 u1_u14_u0_U19 (.A( u1_u14_u0_n142 ) , .ZN( u1_u14_u0_n165 ) );
  OAI221_X1 u1_u14_u0_U20 (.C1( u1_u14_u0_n121 ) , .ZN( u1_u14_u0_n122 ) , .B2( u1_u14_u0_n127 ) , .A( u1_u14_u0_n143 ) , .B1( u1_u14_u0_n144 ) , .C2( u1_u14_u0_n147 ) );
  OAI22_X1 u1_u14_u0_U21 (.B1( u1_u14_u0_n125 ) , .ZN( u1_u14_u0_n126 ) , .A1( u1_u14_u0_n138 ) , .A2( u1_u14_u0_n146 ) , .B2( u1_u14_u0_n147 ) );
  OAI22_X1 u1_u14_u0_U22 (.B1( u1_u14_u0_n131 ) , .A1( u1_u14_u0_n144 ) , .B2( u1_u14_u0_n147 ) , .A2( u1_u14_u0_n90 ) , .ZN( u1_u14_u0_n91 ) );
  AND3_X1 u1_u14_u0_U23 (.A3( u1_u14_u0_n121 ) , .A2( u1_u14_u0_n125 ) , .A1( u1_u14_u0_n148 ) , .ZN( u1_u14_u0_n90 ) );
  NAND2_X1 u1_u14_u0_U24 (.A1( u1_u14_u0_n100 ) , .A2( u1_u14_u0_n103 ) , .ZN( u1_u14_u0_n125 ) );
  INV_X1 u1_u14_u0_U25 (.A( u1_u14_u0_n136 ) , .ZN( u1_u14_u0_n161 ) );
  NOR2_X1 u1_u14_u0_U26 (.A1( u1_u14_u0_n120 ) , .ZN( u1_u14_u0_n143 ) , .A2( u1_u14_u0_n167 ) );
  OAI221_X1 u1_u14_u0_U27 (.C1( u1_u14_u0_n112 ) , .ZN( u1_u14_u0_n120 ) , .B1( u1_u14_u0_n138 ) , .B2( u1_u14_u0_n141 ) , .C2( u1_u14_u0_n147 ) , .A( u1_u14_u0_n172 ) );
  AOI211_X1 u1_u14_u0_U28 (.B( u1_u14_u0_n115 ) , .A( u1_u14_u0_n116 ) , .C2( u1_u14_u0_n117 ) , .C1( u1_u14_u0_n118 ) , .ZN( u1_u14_u0_n119 ) );
  AOI22_X1 u1_u14_u0_U29 (.B2( u1_u14_u0_n109 ) , .A2( u1_u14_u0_n110 ) , .ZN( u1_u14_u0_n111 ) , .B1( u1_u14_u0_n118 ) , .A1( u1_u14_u0_n160 ) );
  INV_X1 u1_u14_u0_U3 (.A( u1_u14_u0_n113 ) , .ZN( u1_u14_u0_n166 ) );
  NAND2_X1 u1_u14_u0_U30 (.A1( u1_u14_u0_n100 ) , .ZN( u1_u14_u0_n129 ) , .A2( u1_u14_u0_n95 ) );
  INV_X1 u1_u14_u0_U31 (.A( u1_u14_u0_n118 ) , .ZN( u1_u14_u0_n158 ) );
  AOI21_X1 u1_u14_u0_U32 (.ZN( u1_u14_u0_n104 ) , .B1( u1_u14_u0_n107 ) , .B2( u1_u14_u0_n141 ) , .A( u1_u14_u0_n144 ) );
  AOI21_X1 u1_u14_u0_U33 (.B1( u1_u14_u0_n127 ) , .B2( u1_u14_u0_n129 ) , .A( u1_u14_u0_n138 ) , .ZN( u1_u14_u0_n96 ) );
  AOI21_X1 u1_u14_u0_U34 (.ZN( u1_u14_u0_n116 ) , .B2( u1_u14_u0_n142 ) , .A( u1_u14_u0_n144 ) , .B1( u1_u14_u0_n166 ) );
  NAND2_X1 u1_u14_u0_U35 (.A2( u1_u14_u0_n100 ) , .A1( u1_u14_u0_n101 ) , .ZN( u1_u14_u0_n139 ) );
  NAND2_X1 u1_u14_u0_U36 (.A2( u1_u14_u0_n100 ) , .ZN( u1_u14_u0_n131 ) , .A1( u1_u14_u0_n92 ) );
  NAND2_X1 u1_u14_u0_U37 (.A1( u1_u14_u0_n101 ) , .A2( u1_u14_u0_n102 ) , .ZN( u1_u14_u0_n150 ) );
  INV_X1 u1_u14_u0_U38 (.A( u1_u14_u0_n138 ) , .ZN( u1_u14_u0_n160 ) );
  NAND2_X1 u1_u14_u0_U39 (.A1( u1_u14_u0_n102 ) , .ZN( u1_u14_u0_n128 ) , .A2( u1_u14_u0_n95 ) );
  AOI21_X1 u1_u14_u0_U4 (.B1( u1_u14_u0_n114 ) , .ZN( u1_u14_u0_n115 ) , .B2( u1_u14_u0_n129 ) , .A( u1_u14_u0_n161 ) );
  NAND2_X1 u1_u14_u0_U40 (.ZN( u1_u14_u0_n148 ) , .A1( u1_u14_u0_n93 ) , .A2( u1_u14_u0_n95 ) );
  NAND2_X1 u1_u14_u0_U41 (.A2( u1_u14_u0_n102 ) , .A1( u1_u14_u0_n103 ) , .ZN( u1_u14_u0_n149 ) );
  NAND2_X1 u1_u14_u0_U42 (.A2( u1_u14_u0_n102 ) , .ZN( u1_u14_u0_n114 ) , .A1( u1_u14_u0_n92 ) );
  NAND2_X1 u1_u14_u0_U43 (.A2( u1_u14_u0_n101 ) , .ZN( u1_u14_u0_n121 ) , .A1( u1_u14_u0_n93 ) );
  INV_X1 u1_u14_u0_U44 (.ZN( u1_u14_u0_n172 ) , .A( u1_u14_u0_n88 ) );
  OAI222_X1 u1_u14_u0_U45 (.C1( u1_u14_u0_n108 ) , .A1( u1_u14_u0_n125 ) , .B2( u1_u14_u0_n128 ) , .B1( u1_u14_u0_n144 ) , .A2( u1_u14_u0_n158 ) , .C2( u1_u14_u0_n161 ) , .ZN( u1_u14_u0_n88 ) );
  NAND2_X1 u1_u14_u0_U46 (.ZN( u1_u14_u0_n112 ) , .A2( u1_u14_u0_n92 ) , .A1( u1_u14_u0_n93 ) );
  OR3_X1 u1_u14_u0_U47 (.A3( u1_u14_u0_n152 ) , .A2( u1_u14_u0_n153 ) , .A1( u1_u14_u0_n154 ) , .ZN( u1_u14_u0_n155 ) );
  AOI21_X1 u1_u14_u0_U48 (.B2( u1_u14_u0_n150 ) , .B1( u1_u14_u0_n151 ) , .ZN( u1_u14_u0_n152 ) , .A( u1_u14_u0_n158 ) );
  AOI21_X1 u1_u14_u0_U49 (.A( u1_u14_u0_n144 ) , .B2( u1_u14_u0_n145 ) , .B1( u1_u14_u0_n146 ) , .ZN( u1_u14_u0_n154 ) );
  AOI21_X1 u1_u14_u0_U5 (.B2( u1_u14_u0_n131 ) , .ZN( u1_u14_u0_n134 ) , .B1( u1_u14_u0_n151 ) , .A( u1_u14_u0_n158 ) );
  AOI21_X1 u1_u14_u0_U50 (.A( u1_u14_u0_n147 ) , .B2( u1_u14_u0_n148 ) , .B1( u1_u14_u0_n149 ) , .ZN( u1_u14_u0_n153 ) );
  INV_X1 u1_u14_u0_U51 (.ZN( u1_u14_u0_n171 ) , .A( u1_u14_u0_n99 ) );
  OAI211_X1 u1_u14_u0_U52 (.C2( u1_u14_u0_n140 ) , .C1( u1_u14_u0_n161 ) , .A( u1_u14_u0_n169 ) , .B( u1_u14_u0_n98 ) , .ZN( u1_u14_u0_n99 ) );
  AOI211_X1 u1_u14_u0_U53 (.C1( u1_u14_u0_n118 ) , .A( u1_u14_u0_n123 ) , .B( u1_u14_u0_n96 ) , .C2( u1_u14_u0_n97 ) , .ZN( u1_u14_u0_n98 ) );
  INV_X1 u1_u14_u0_U54 (.ZN( u1_u14_u0_n169 ) , .A( u1_u14_u0_n91 ) );
  NOR2_X1 u1_u14_u0_U55 (.A2( u1_u14_X_4 ) , .A1( u1_u14_X_5 ) , .ZN( u1_u14_u0_n118 ) );
  NOR2_X1 u1_u14_u0_U56 (.A2( u1_u14_X_2 ) , .ZN( u1_u14_u0_n103 ) , .A1( u1_u14_u0_n164 ) );
  NOR2_X1 u1_u14_u0_U57 (.A2( u1_u14_X_1 ) , .A1( u1_u14_X_2 ) , .ZN( u1_u14_u0_n92 ) );
  NOR2_X1 u1_u14_u0_U58 (.A2( u1_u14_X_1 ) , .ZN( u1_u14_u0_n101 ) , .A1( u1_u14_u0_n163 ) );
  NAND2_X1 u1_u14_u0_U59 (.A2( u1_u14_X_4 ) , .A1( u1_u14_X_5 ) , .ZN( u1_u14_u0_n144 ) );
  NOR2_X1 u1_u14_u0_U6 (.A1( u1_u14_u0_n108 ) , .ZN( u1_u14_u0_n123 ) , .A2( u1_u14_u0_n158 ) );
  NOR2_X1 u1_u14_u0_U60 (.A2( u1_u14_X_5 ) , .ZN( u1_u14_u0_n136 ) , .A1( u1_u14_u0_n159 ) );
  NAND2_X1 u1_u14_u0_U61 (.A1( u1_u14_X_5 ) , .ZN( u1_u14_u0_n138 ) , .A2( u1_u14_u0_n159 ) );
  AND2_X1 u1_u14_u0_U62 (.A2( u1_u14_X_3 ) , .A1( u1_u14_X_6 ) , .ZN( u1_u14_u0_n102 ) );
  AND2_X1 u1_u14_u0_U63 (.A1( u1_u14_X_6 ) , .A2( u1_u14_u0_n162 ) , .ZN( u1_u14_u0_n93 ) );
  INV_X1 u1_u14_u0_U64 (.A( u1_u14_X_4 ) , .ZN( u1_u14_u0_n159 ) );
  INV_X1 u1_u14_u0_U65 (.A( u1_u14_X_1 ) , .ZN( u1_u14_u0_n164 ) );
  INV_X1 u1_u14_u0_U66 (.A( u1_u14_X_2 ) , .ZN( u1_u14_u0_n163 ) );
  INV_X1 u1_u14_u0_U67 (.A( u1_u14_X_3 ) , .ZN( u1_u14_u0_n162 ) );
  INV_X1 u1_u14_u0_U68 (.A( u1_u14_u0_n126 ) , .ZN( u1_u14_u0_n168 ) );
  AOI211_X1 u1_u14_u0_U69 (.B( u1_u14_u0_n133 ) , .A( u1_u14_u0_n134 ) , .C2( u1_u14_u0_n135 ) , .C1( u1_u14_u0_n136 ) , .ZN( u1_u14_u0_n137 ) );
  OAI21_X1 u1_u14_u0_U7 (.B1( u1_u14_u0_n150 ) , .B2( u1_u14_u0_n158 ) , .A( u1_u14_u0_n172 ) , .ZN( u1_u14_u0_n89 ) );
  INV_X1 u1_u14_u0_U70 (.ZN( u1_u14_u0_n174 ) , .A( u1_u14_u0_n89 ) );
  AOI211_X1 u1_u14_u0_U71 (.B( u1_u14_u0_n104 ) , .A( u1_u14_u0_n105 ) , .ZN( u1_u14_u0_n106 ) , .C2( u1_u14_u0_n113 ) , .C1( u1_u14_u0_n160 ) );
  OR4_X1 u1_u14_u0_U72 (.ZN( u1_out14_17 ) , .A4( u1_u14_u0_n122 ) , .A2( u1_u14_u0_n123 ) , .A1( u1_u14_u0_n124 ) , .A3( u1_u14_u0_n170 ) );
  AOI21_X1 u1_u14_u0_U73 (.B2( u1_u14_u0_n107 ) , .ZN( u1_u14_u0_n124 ) , .B1( u1_u14_u0_n128 ) , .A( u1_u14_u0_n161 ) );
  INV_X1 u1_u14_u0_U74 (.A( u1_u14_u0_n111 ) , .ZN( u1_u14_u0_n170 ) );
  OR4_X1 u1_u14_u0_U75 (.ZN( u1_out14_31 ) , .A4( u1_u14_u0_n155 ) , .A2( u1_u14_u0_n156 ) , .A1( u1_u14_u0_n157 ) , .A3( u1_u14_u0_n173 ) );
  AOI21_X1 u1_u14_u0_U76 (.A( u1_u14_u0_n138 ) , .B2( u1_u14_u0_n139 ) , .B1( u1_u14_u0_n140 ) , .ZN( u1_u14_u0_n157 ) );
  AOI21_X1 u1_u14_u0_U77 (.B2( u1_u14_u0_n141 ) , .B1( u1_u14_u0_n142 ) , .ZN( u1_u14_u0_n156 ) , .A( u1_u14_u0_n161 ) );
  AOI21_X1 u1_u14_u0_U78 (.B1( u1_u14_u0_n132 ) , .ZN( u1_u14_u0_n133 ) , .A( u1_u14_u0_n144 ) , .B2( u1_u14_u0_n166 ) );
  OAI22_X1 u1_u14_u0_U79 (.ZN( u1_u14_u0_n105 ) , .A2( u1_u14_u0_n132 ) , .B1( u1_u14_u0_n146 ) , .A1( u1_u14_u0_n147 ) , .B2( u1_u14_u0_n161 ) );
  AND2_X1 u1_u14_u0_U8 (.A1( u1_u14_u0_n114 ) , .A2( u1_u14_u0_n121 ) , .ZN( u1_u14_u0_n146 ) );
  NAND2_X1 u1_u14_u0_U80 (.ZN( u1_u14_u0_n110 ) , .A2( u1_u14_u0_n132 ) , .A1( u1_u14_u0_n145 ) );
  INV_X1 u1_u14_u0_U81 (.A( u1_u14_u0_n119 ) , .ZN( u1_u14_u0_n167 ) );
  NAND2_X1 u1_u14_u0_U82 (.A2( u1_u14_u0_n103 ) , .ZN( u1_u14_u0_n140 ) , .A1( u1_u14_u0_n94 ) );
  NAND2_X1 u1_u14_u0_U83 (.A1( u1_u14_u0_n101 ) , .ZN( u1_u14_u0_n130 ) , .A2( u1_u14_u0_n94 ) );
  NAND2_X1 u1_u14_u0_U84 (.ZN( u1_u14_u0_n108 ) , .A1( u1_u14_u0_n92 ) , .A2( u1_u14_u0_n94 ) );
  NAND2_X1 u1_u14_u0_U85 (.ZN( u1_u14_u0_n142 ) , .A1( u1_u14_u0_n94 ) , .A2( u1_u14_u0_n95 ) );
  NOR2_X1 u1_u14_u0_U86 (.A2( u1_u14_X_6 ) , .ZN( u1_u14_u0_n100 ) , .A1( u1_u14_u0_n162 ) );
  NOR2_X1 u1_u14_u0_U87 (.A2( u1_u14_X_3 ) , .A1( u1_u14_X_6 ) , .ZN( u1_u14_u0_n94 ) );
  NAND3_X1 u1_u14_u0_U88 (.ZN( u1_out14_23 ) , .A3( u1_u14_u0_n137 ) , .A1( u1_u14_u0_n168 ) , .A2( u1_u14_u0_n171 ) );
  NAND3_X1 u1_u14_u0_U89 (.A3( u1_u14_u0_n127 ) , .A2( u1_u14_u0_n128 ) , .ZN( u1_u14_u0_n135 ) , .A1( u1_u14_u0_n150 ) );
  AND2_X1 u1_u14_u0_U9 (.A1( u1_u14_u0_n131 ) , .ZN( u1_u14_u0_n141 ) , .A2( u1_u14_u0_n150 ) );
  NAND3_X1 u1_u14_u0_U90 (.ZN( u1_u14_u0_n117 ) , .A3( u1_u14_u0_n132 ) , .A2( u1_u14_u0_n139 ) , .A1( u1_u14_u0_n148 ) );
  NAND3_X1 u1_u14_u0_U91 (.ZN( u1_u14_u0_n109 ) , .A2( u1_u14_u0_n114 ) , .A3( u1_u14_u0_n140 ) , .A1( u1_u14_u0_n149 ) );
  NAND3_X1 u1_u14_u0_U92 (.ZN( u1_out14_9 ) , .A3( u1_u14_u0_n106 ) , .A2( u1_u14_u0_n171 ) , .A1( u1_u14_u0_n174 ) );
  NAND3_X1 u1_u14_u0_U93 (.A2( u1_u14_u0_n128 ) , .A1( u1_u14_u0_n132 ) , .A3( u1_u14_u0_n146 ) , .ZN( u1_u14_u0_n97 ) );
  AOI21_X1 u1_u14_u1_U10 (.ZN( u1_u14_u1_n106 ) , .A( u1_u14_u1_n112 ) , .B1( u1_u14_u1_n154 ) , .B2( u1_u14_u1_n156 ) );
  NAND3_X1 u1_u14_u1_U100 (.ZN( u1_u14_u1_n113 ) , .A1( u1_u14_u1_n120 ) , .A3( u1_u14_u1_n133 ) , .A2( u1_u14_u1_n155 ) );
  INV_X1 u1_u14_u1_U11 (.A( u1_u14_u1_n101 ) , .ZN( u1_u14_u1_n184 ) );
  AOI21_X1 u1_u14_u1_U12 (.ZN( u1_u14_u1_n107 ) , .B1( u1_u14_u1_n134 ) , .B2( u1_u14_u1_n149 ) , .A( u1_u14_u1_n174 ) );
  NAND2_X1 u1_u14_u1_U13 (.ZN( u1_u14_u1_n140 ) , .A2( u1_u14_u1_n150 ) , .A1( u1_u14_u1_n155 ) );
  NAND2_X1 u1_u14_u1_U14 (.A1( u1_u14_u1_n131 ) , .ZN( u1_u14_u1_n147 ) , .A2( u1_u14_u1_n153 ) );
  AOI22_X1 u1_u14_u1_U15 (.B2( u1_u14_u1_n136 ) , .A2( u1_u14_u1_n137 ) , .ZN( u1_u14_u1_n143 ) , .A1( u1_u14_u1_n171 ) , .B1( u1_u14_u1_n173 ) );
  INV_X1 u1_u14_u1_U16 (.A( u1_u14_u1_n147 ) , .ZN( u1_u14_u1_n181 ) );
  INV_X1 u1_u14_u1_U17 (.A( u1_u14_u1_n139 ) , .ZN( u1_u14_u1_n174 ) );
  INV_X1 u1_u14_u1_U18 (.A( u1_u14_u1_n112 ) , .ZN( u1_u14_u1_n171 ) );
  NAND2_X1 u1_u14_u1_U19 (.ZN( u1_u14_u1_n141 ) , .A1( u1_u14_u1_n153 ) , .A2( u1_u14_u1_n156 ) );
  AND2_X1 u1_u14_u1_U20 (.A1( u1_u14_u1_n123 ) , .ZN( u1_u14_u1_n134 ) , .A2( u1_u14_u1_n161 ) );
  NAND2_X1 u1_u14_u1_U21 (.A2( u1_u14_u1_n115 ) , .A1( u1_u14_u1_n116 ) , .ZN( u1_u14_u1_n148 ) );
  NAND2_X1 u1_u14_u1_U22 (.A2( u1_u14_u1_n133 ) , .A1( u1_u14_u1_n135 ) , .ZN( u1_u14_u1_n159 ) );
  NAND2_X1 u1_u14_u1_U23 (.A2( u1_u14_u1_n115 ) , .A1( u1_u14_u1_n120 ) , .ZN( u1_u14_u1_n132 ) );
  INV_X1 u1_u14_u1_U24 (.A( u1_u14_u1_n154 ) , .ZN( u1_u14_u1_n178 ) );
  AOI22_X1 u1_u14_u1_U25 (.B2( u1_u14_u1_n113 ) , .A2( u1_u14_u1_n114 ) , .ZN( u1_u14_u1_n125 ) , .A1( u1_u14_u1_n171 ) , .B1( u1_u14_u1_n173 ) );
  NAND2_X1 u1_u14_u1_U26 (.ZN( u1_u14_u1_n114 ) , .A1( u1_u14_u1_n134 ) , .A2( u1_u14_u1_n156 ) );
  INV_X1 u1_u14_u1_U27 (.A( u1_u14_u1_n151 ) , .ZN( u1_u14_u1_n183 ) );
  AND2_X1 u1_u14_u1_U28 (.A1( u1_u14_u1_n129 ) , .A2( u1_u14_u1_n133 ) , .ZN( u1_u14_u1_n149 ) );
  INV_X1 u1_u14_u1_U29 (.A( u1_u14_u1_n131 ) , .ZN( u1_u14_u1_n180 ) );
  INV_X1 u1_u14_u1_U3 (.A( u1_u14_u1_n159 ) , .ZN( u1_u14_u1_n182 ) );
  AOI221_X1 u1_u14_u1_U30 (.B1( u1_u14_u1_n140 ) , .ZN( u1_u14_u1_n167 ) , .B2( u1_u14_u1_n172 ) , .C2( u1_u14_u1_n175 ) , .C1( u1_u14_u1_n178 ) , .A( u1_u14_u1_n188 ) );
  INV_X1 u1_u14_u1_U31 (.ZN( u1_u14_u1_n188 ) , .A( u1_u14_u1_n97 ) );
  AOI211_X1 u1_u14_u1_U32 (.A( u1_u14_u1_n118 ) , .C1( u1_u14_u1_n132 ) , .C2( u1_u14_u1_n139 ) , .B( u1_u14_u1_n96 ) , .ZN( u1_u14_u1_n97 ) );
  AOI21_X1 u1_u14_u1_U33 (.B2( u1_u14_u1_n121 ) , .B1( u1_u14_u1_n135 ) , .A( u1_u14_u1_n152 ) , .ZN( u1_u14_u1_n96 ) );
  OAI221_X1 u1_u14_u1_U34 (.A( u1_u14_u1_n119 ) , .C2( u1_u14_u1_n129 ) , .ZN( u1_u14_u1_n138 ) , .B2( u1_u14_u1_n152 ) , .C1( u1_u14_u1_n174 ) , .B1( u1_u14_u1_n187 ) );
  INV_X1 u1_u14_u1_U35 (.A( u1_u14_u1_n148 ) , .ZN( u1_u14_u1_n187 ) );
  AOI211_X1 u1_u14_u1_U36 (.B( u1_u14_u1_n117 ) , .A( u1_u14_u1_n118 ) , .ZN( u1_u14_u1_n119 ) , .C2( u1_u14_u1_n146 ) , .C1( u1_u14_u1_n159 ) );
  NOR2_X1 u1_u14_u1_U37 (.A1( u1_u14_u1_n168 ) , .A2( u1_u14_u1_n176 ) , .ZN( u1_u14_u1_n98 ) );
  AOI211_X1 u1_u14_u1_U38 (.B( u1_u14_u1_n162 ) , .A( u1_u14_u1_n163 ) , .C2( u1_u14_u1_n164 ) , .ZN( u1_u14_u1_n165 ) , .C1( u1_u14_u1_n171 ) );
  AOI21_X1 u1_u14_u1_U39 (.A( u1_u14_u1_n160 ) , .B2( u1_u14_u1_n161 ) , .ZN( u1_u14_u1_n162 ) , .B1( u1_u14_u1_n182 ) );
  AOI221_X1 u1_u14_u1_U4 (.A( u1_u14_u1_n138 ) , .C2( u1_u14_u1_n139 ) , .C1( u1_u14_u1_n140 ) , .B2( u1_u14_u1_n141 ) , .ZN( u1_u14_u1_n142 ) , .B1( u1_u14_u1_n175 ) );
  OR2_X1 u1_u14_u1_U40 (.A2( u1_u14_u1_n157 ) , .A1( u1_u14_u1_n158 ) , .ZN( u1_u14_u1_n163 ) );
  OAI21_X1 u1_u14_u1_U41 (.B2( u1_u14_u1_n123 ) , .ZN( u1_u14_u1_n145 ) , .B1( u1_u14_u1_n160 ) , .A( u1_u14_u1_n185 ) );
  INV_X1 u1_u14_u1_U42 (.A( u1_u14_u1_n122 ) , .ZN( u1_u14_u1_n185 ) );
  AOI21_X1 u1_u14_u1_U43 (.B2( u1_u14_u1_n120 ) , .B1( u1_u14_u1_n121 ) , .ZN( u1_u14_u1_n122 ) , .A( u1_u14_u1_n128 ) );
  NAND2_X1 u1_u14_u1_U44 (.A1( u1_u14_u1_n128 ) , .ZN( u1_u14_u1_n146 ) , .A2( u1_u14_u1_n160 ) );
  NAND2_X1 u1_u14_u1_U45 (.A2( u1_u14_u1_n112 ) , .ZN( u1_u14_u1_n139 ) , .A1( u1_u14_u1_n152 ) );
  NAND2_X1 u1_u14_u1_U46 (.A1( u1_u14_u1_n105 ) , .ZN( u1_u14_u1_n156 ) , .A2( u1_u14_u1_n99 ) );
  NOR2_X1 u1_u14_u1_U47 (.ZN( u1_u14_u1_n117 ) , .A1( u1_u14_u1_n121 ) , .A2( u1_u14_u1_n160 ) );
  AOI21_X1 u1_u14_u1_U48 (.A( u1_u14_u1_n128 ) , .B2( u1_u14_u1_n129 ) , .ZN( u1_u14_u1_n130 ) , .B1( u1_u14_u1_n150 ) );
  NAND2_X1 u1_u14_u1_U49 (.ZN( u1_u14_u1_n112 ) , .A1( u1_u14_u1_n169 ) , .A2( u1_u14_u1_n170 ) );
  AOI211_X1 u1_u14_u1_U5 (.ZN( u1_u14_u1_n124 ) , .A( u1_u14_u1_n138 ) , .C2( u1_u14_u1_n139 ) , .B( u1_u14_u1_n145 ) , .C1( u1_u14_u1_n147 ) );
  NAND2_X1 u1_u14_u1_U50 (.ZN( u1_u14_u1_n129 ) , .A2( u1_u14_u1_n95 ) , .A1( u1_u14_u1_n98 ) );
  NAND2_X1 u1_u14_u1_U51 (.A1( u1_u14_u1_n102 ) , .ZN( u1_u14_u1_n154 ) , .A2( u1_u14_u1_n99 ) );
  NAND2_X1 u1_u14_u1_U52 (.A2( u1_u14_u1_n100 ) , .ZN( u1_u14_u1_n135 ) , .A1( u1_u14_u1_n99 ) );
  AOI21_X1 u1_u14_u1_U53 (.A( u1_u14_u1_n152 ) , .B2( u1_u14_u1_n153 ) , .B1( u1_u14_u1_n154 ) , .ZN( u1_u14_u1_n158 ) );
  INV_X1 u1_u14_u1_U54 (.A( u1_u14_u1_n160 ) , .ZN( u1_u14_u1_n175 ) );
  NAND2_X1 u1_u14_u1_U55 (.A1( u1_u14_u1_n100 ) , .ZN( u1_u14_u1_n116 ) , .A2( u1_u14_u1_n95 ) );
  NAND2_X1 u1_u14_u1_U56 (.A1( u1_u14_u1_n102 ) , .ZN( u1_u14_u1_n131 ) , .A2( u1_u14_u1_n95 ) );
  NAND2_X1 u1_u14_u1_U57 (.A2( u1_u14_u1_n104 ) , .ZN( u1_u14_u1_n121 ) , .A1( u1_u14_u1_n98 ) );
  NAND2_X1 u1_u14_u1_U58 (.A1( u1_u14_u1_n103 ) , .ZN( u1_u14_u1_n153 ) , .A2( u1_u14_u1_n98 ) );
  NAND2_X1 u1_u14_u1_U59 (.A2( u1_u14_u1_n104 ) , .A1( u1_u14_u1_n105 ) , .ZN( u1_u14_u1_n133 ) );
  NOR2_X1 u1_u14_u1_U6 (.A1( u1_u14_u1_n112 ) , .A2( u1_u14_u1_n116 ) , .ZN( u1_u14_u1_n118 ) );
  NAND2_X1 u1_u14_u1_U60 (.ZN( u1_u14_u1_n150 ) , .A2( u1_u14_u1_n98 ) , .A1( u1_u14_u1_n99 ) );
  NAND2_X1 u1_u14_u1_U61 (.A1( u1_u14_u1_n105 ) , .ZN( u1_u14_u1_n155 ) , .A2( u1_u14_u1_n95 ) );
  OAI21_X1 u1_u14_u1_U62 (.ZN( u1_u14_u1_n109 ) , .B1( u1_u14_u1_n129 ) , .B2( u1_u14_u1_n160 ) , .A( u1_u14_u1_n167 ) );
  NAND2_X1 u1_u14_u1_U63 (.A2( u1_u14_u1_n100 ) , .A1( u1_u14_u1_n103 ) , .ZN( u1_u14_u1_n120 ) );
  NAND2_X1 u1_u14_u1_U64 (.A1( u1_u14_u1_n102 ) , .A2( u1_u14_u1_n104 ) , .ZN( u1_u14_u1_n115 ) );
  NAND2_X1 u1_u14_u1_U65 (.A2( u1_u14_u1_n100 ) , .A1( u1_u14_u1_n104 ) , .ZN( u1_u14_u1_n151 ) );
  NAND2_X1 u1_u14_u1_U66 (.A2( u1_u14_u1_n103 ) , .A1( u1_u14_u1_n105 ) , .ZN( u1_u14_u1_n161 ) );
  INV_X1 u1_u14_u1_U67 (.A( u1_u14_u1_n152 ) , .ZN( u1_u14_u1_n173 ) );
  INV_X1 u1_u14_u1_U68 (.A( u1_u14_u1_n128 ) , .ZN( u1_u14_u1_n172 ) );
  NAND2_X1 u1_u14_u1_U69 (.A2( u1_u14_u1_n102 ) , .A1( u1_u14_u1_n103 ) , .ZN( u1_u14_u1_n123 ) );
  OAI21_X1 u1_u14_u1_U7 (.ZN( u1_u14_u1_n101 ) , .B1( u1_u14_u1_n141 ) , .A( u1_u14_u1_n146 ) , .B2( u1_u14_u1_n183 ) );
  NOR2_X1 u1_u14_u1_U70 (.A2( u1_u14_X_7 ) , .A1( u1_u14_X_8 ) , .ZN( u1_u14_u1_n95 ) );
  NOR2_X1 u1_u14_u1_U71 (.A1( u1_u14_X_12 ) , .A2( u1_u14_X_9 ) , .ZN( u1_u14_u1_n100 ) );
  NOR2_X1 u1_u14_u1_U72 (.A2( u1_u14_X_8 ) , .A1( u1_u14_u1_n177 ) , .ZN( u1_u14_u1_n99 ) );
  NOR2_X1 u1_u14_u1_U73 (.A2( u1_u14_X_12 ) , .ZN( u1_u14_u1_n102 ) , .A1( u1_u14_u1_n176 ) );
  NOR2_X1 u1_u14_u1_U74 (.A2( u1_u14_X_9 ) , .ZN( u1_u14_u1_n105 ) , .A1( u1_u14_u1_n168 ) );
  NAND2_X1 u1_u14_u1_U75 (.A1( u1_u14_X_10 ) , .ZN( u1_u14_u1_n160 ) , .A2( u1_u14_u1_n169 ) );
  NAND2_X1 u1_u14_u1_U76 (.A2( u1_u14_X_10 ) , .A1( u1_u14_X_11 ) , .ZN( u1_u14_u1_n152 ) );
  NAND2_X1 u1_u14_u1_U77 (.A1( u1_u14_X_11 ) , .ZN( u1_u14_u1_n128 ) , .A2( u1_u14_u1_n170 ) );
  AND2_X1 u1_u14_u1_U78 (.A2( u1_u14_X_7 ) , .A1( u1_u14_X_8 ) , .ZN( u1_u14_u1_n104 ) );
  AND2_X1 u1_u14_u1_U79 (.A1( u1_u14_X_8 ) , .ZN( u1_u14_u1_n103 ) , .A2( u1_u14_u1_n177 ) );
  AOI21_X1 u1_u14_u1_U8 (.B2( u1_u14_u1_n155 ) , .B1( u1_u14_u1_n156 ) , .ZN( u1_u14_u1_n157 ) , .A( u1_u14_u1_n174 ) );
  INV_X1 u1_u14_u1_U80 (.A( u1_u14_X_10 ) , .ZN( u1_u14_u1_n170 ) );
  INV_X1 u1_u14_u1_U81 (.A( u1_u14_X_9 ) , .ZN( u1_u14_u1_n176 ) );
  INV_X1 u1_u14_u1_U82 (.A( u1_u14_X_11 ) , .ZN( u1_u14_u1_n169 ) );
  INV_X1 u1_u14_u1_U83 (.A( u1_u14_X_12 ) , .ZN( u1_u14_u1_n168 ) );
  INV_X1 u1_u14_u1_U84 (.A( u1_u14_X_7 ) , .ZN( u1_u14_u1_n177 ) );
  NAND4_X1 u1_u14_u1_U85 (.ZN( u1_out14_18 ) , .A4( u1_u14_u1_n165 ) , .A3( u1_u14_u1_n166 ) , .A1( u1_u14_u1_n167 ) , .A2( u1_u14_u1_n186 ) );
  AOI22_X1 u1_u14_u1_U86 (.B2( u1_u14_u1_n146 ) , .B1( u1_u14_u1_n147 ) , .A2( u1_u14_u1_n148 ) , .ZN( u1_u14_u1_n166 ) , .A1( u1_u14_u1_n172 ) );
  INV_X1 u1_u14_u1_U87 (.A( u1_u14_u1_n145 ) , .ZN( u1_u14_u1_n186 ) );
  OR4_X1 u1_u14_u1_U88 (.ZN( u1_out14_13 ) , .A4( u1_u14_u1_n108 ) , .A3( u1_u14_u1_n109 ) , .A2( u1_u14_u1_n110 ) , .A1( u1_u14_u1_n111 ) );
  AOI21_X1 u1_u14_u1_U89 (.ZN( u1_u14_u1_n111 ) , .A( u1_u14_u1_n128 ) , .B2( u1_u14_u1_n131 ) , .B1( u1_u14_u1_n135 ) );
  OR4_X1 u1_u14_u1_U9 (.A4( u1_u14_u1_n106 ) , .A3( u1_u14_u1_n107 ) , .ZN( u1_u14_u1_n108 ) , .A1( u1_u14_u1_n117 ) , .A2( u1_u14_u1_n184 ) );
  AOI21_X1 u1_u14_u1_U90 (.ZN( u1_u14_u1_n110 ) , .A( u1_u14_u1_n116 ) , .B1( u1_u14_u1_n152 ) , .B2( u1_u14_u1_n160 ) );
  NAND4_X1 u1_u14_u1_U91 (.ZN( u1_out14_2 ) , .A4( u1_u14_u1_n142 ) , .A3( u1_u14_u1_n143 ) , .A2( u1_u14_u1_n144 ) , .A1( u1_u14_u1_n179 ) );
  OAI21_X1 u1_u14_u1_U92 (.B2( u1_u14_u1_n132 ) , .ZN( u1_u14_u1_n144 ) , .A( u1_u14_u1_n146 ) , .B1( u1_u14_u1_n180 ) );
  INV_X1 u1_u14_u1_U93 (.A( u1_u14_u1_n130 ) , .ZN( u1_u14_u1_n179 ) );
  NAND4_X1 u1_u14_u1_U94 (.ZN( u1_out14_28 ) , .A4( u1_u14_u1_n124 ) , .A3( u1_u14_u1_n125 ) , .A2( u1_u14_u1_n126 ) , .A1( u1_u14_u1_n127 ) );
  OAI21_X1 u1_u14_u1_U95 (.ZN( u1_u14_u1_n127 ) , .B2( u1_u14_u1_n139 ) , .B1( u1_u14_u1_n175 ) , .A( u1_u14_u1_n183 ) );
  OAI21_X1 u1_u14_u1_U96 (.ZN( u1_u14_u1_n126 ) , .B2( u1_u14_u1_n140 ) , .A( u1_u14_u1_n146 ) , .B1( u1_u14_u1_n178 ) );
  NAND3_X1 u1_u14_u1_U97 (.A3( u1_u14_u1_n149 ) , .A2( u1_u14_u1_n150 ) , .A1( u1_u14_u1_n151 ) , .ZN( u1_u14_u1_n164 ) );
  NAND3_X1 u1_u14_u1_U98 (.A3( u1_u14_u1_n134 ) , .A2( u1_u14_u1_n135 ) , .ZN( u1_u14_u1_n136 ) , .A1( u1_u14_u1_n151 ) );
  NAND3_X1 u1_u14_u1_U99 (.A1( u1_u14_u1_n133 ) , .ZN( u1_u14_u1_n137 ) , .A2( u1_u14_u1_n154 ) , .A3( u1_u14_u1_n181 ) );
  OAI22_X1 u1_u14_u2_U10 (.ZN( u1_u14_u2_n109 ) , .A2( u1_u14_u2_n113 ) , .B2( u1_u14_u2_n133 ) , .B1( u1_u14_u2_n167 ) , .A1( u1_u14_u2_n168 ) );
  NAND3_X1 u1_u14_u2_U100 (.A2( u1_u14_u2_n100 ) , .A1( u1_u14_u2_n104 ) , .A3( u1_u14_u2_n138 ) , .ZN( u1_u14_u2_n98 ) );
  OAI22_X1 u1_u14_u2_U11 (.B1( u1_u14_u2_n151 ) , .A2( u1_u14_u2_n152 ) , .A1( u1_u14_u2_n153 ) , .ZN( u1_u14_u2_n160 ) , .B2( u1_u14_u2_n168 ) );
  NOR3_X1 u1_u14_u2_U12 (.A1( u1_u14_u2_n150 ) , .ZN( u1_u14_u2_n151 ) , .A3( u1_u14_u2_n175 ) , .A2( u1_u14_u2_n188 ) );
  AOI21_X1 u1_u14_u2_U13 (.ZN( u1_u14_u2_n144 ) , .B2( u1_u14_u2_n155 ) , .A( u1_u14_u2_n172 ) , .B1( u1_u14_u2_n185 ) );
  AOI21_X1 u1_u14_u2_U14 (.B2( u1_u14_u2_n143 ) , .ZN( u1_u14_u2_n145 ) , .B1( u1_u14_u2_n152 ) , .A( u1_u14_u2_n171 ) );
  AOI21_X1 u1_u14_u2_U15 (.B2( u1_u14_u2_n120 ) , .B1( u1_u14_u2_n121 ) , .ZN( u1_u14_u2_n126 ) , .A( u1_u14_u2_n167 ) );
  INV_X1 u1_u14_u2_U16 (.A( u1_u14_u2_n156 ) , .ZN( u1_u14_u2_n171 ) );
  INV_X1 u1_u14_u2_U17 (.A( u1_u14_u2_n120 ) , .ZN( u1_u14_u2_n188 ) );
  NAND2_X1 u1_u14_u2_U18 (.A2( u1_u14_u2_n122 ) , .ZN( u1_u14_u2_n150 ) , .A1( u1_u14_u2_n152 ) );
  INV_X1 u1_u14_u2_U19 (.A( u1_u14_u2_n153 ) , .ZN( u1_u14_u2_n170 ) );
  INV_X1 u1_u14_u2_U20 (.A( u1_u14_u2_n137 ) , .ZN( u1_u14_u2_n173 ) );
  NAND2_X1 u1_u14_u2_U21 (.A1( u1_u14_u2_n132 ) , .A2( u1_u14_u2_n139 ) , .ZN( u1_u14_u2_n157 ) );
  INV_X1 u1_u14_u2_U22 (.A( u1_u14_u2_n113 ) , .ZN( u1_u14_u2_n178 ) );
  INV_X1 u1_u14_u2_U23 (.A( u1_u14_u2_n139 ) , .ZN( u1_u14_u2_n175 ) );
  INV_X1 u1_u14_u2_U24 (.A( u1_u14_u2_n155 ) , .ZN( u1_u14_u2_n181 ) );
  INV_X1 u1_u14_u2_U25 (.A( u1_u14_u2_n119 ) , .ZN( u1_u14_u2_n177 ) );
  INV_X1 u1_u14_u2_U26 (.A( u1_u14_u2_n116 ) , .ZN( u1_u14_u2_n180 ) );
  INV_X1 u1_u14_u2_U27 (.A( u1_u14_u2_n131 ) , .ZN( u1_u14_u2_n179 ) );
  INV_X1 u1_u14_u2_U28 (.A( u1_u14_u2_n154 ) , .ZN( u1_u14_u2_n176 ) );
  NAND2_X1 u1_u14_u2_U29 (.A2( u1_u14_u2_n116 ) , .A1( u1_u14_u2_n117 ) , .ZN( u1_u14_u2_n118 ) );
  NOR2_X1 u1_u14_u2_U3 (.ZN( u1_u14_u2_n121 ) , .A2( u1_u14_u2_n177 ) , .A1( u1_u14_u2_n180 ) );
  INV_X1 u1_u14_u2_U30 (.A( u1_u14_u2_n132 ) , .ZN( u1_u14_u2_n182 ) );
  INV_X1 u1_u14_u2_U31 (.A( u1_u14_u2_n158 ) , .ZN( u1_u14_u2_n183 ) );
  OAI21_X1 u1_u14_u2_U32 (.A( u1_u14_u2_n156 ) , .B1( u1_u14_u2_n157 ) , .ZN( u1_u14_u2_n158 ) , .B2( u1_u14_u2_n179 ) );
  NOR2_X1 u1_u14_u2_U33 (.ZN( u1_u14_u2_n156 ) , .A1( u1_u14_u2_n166 ) , .A2( u1_u14_u2_n169 ) );
  NOR2_X1 u1_u14_u2_U34 (.A2( u1_u14_u2_n114 ) , .ZN( u1_u14_u2_n137 ) , .A1( u1_u14_u2_n140 ) );
  NOR2_X1 u1_u14_u2_U35 (.A2( u1_u14_u2_n138 ) , .ZN( u1_u14_u2_n153 ) , .A1( u1_u14_u2_n156 ) );
  AOI211_X1 u1_u14_u2_U36 (.ZN( u1_u14_u2_n130 ) , .C1( u1_u14_u2_n138 ) , .C2( u1_u14_u2_n179 ) , .B( u1_u14_u2_n96 ) , .A( u1_u14_u2_n97 ) );
  OAI22_X1 u1_u14_u2_U37 (.B1( u1_u14_u2_n133 ) , .A2( u1_u14_u2_n137 ) , .A1( u1_u14_u2_n152 ) , .B2( u1_u14_u2_n168 ) , .ZN( u1_u14_u2_n97 ) );
  OAI221_X1 u1_u14_u2_U38 (.B1( u1_u14_u2_n113 ) , .C1( u1_u14_u2_n132 ) , .A( u1_u14_u2_n149 ) , .B2( u1_u14_u2_n171 ) , .C2( u1_u14_u2_n172 ) , .ZN( u1_u14_u2_n96 ) );
  OAI221_X1 u1_u14_u2_U39 (.A( u1_u14_u2_n115 ) , .C2( u1_u14_u2_n123 ) , .B2( u1_u14_u2_n143 ) , .B1( u1_u14_u2_n153 ) , .ZN( u1_u14_u2_n163 ) , .C1( u1_u14_u2_n168 ) );
  INV_X1 u1_u14_u2_U4 (.A( u1_u14_u2_n134 ) , .ZN( u1_u14_u2_n185 ) );
  OAI21_X1 u1_u14_u2_U40 (.A( u1_u14_u2_n114 ) , .ZN( u1_u14_u2_n115 ) , .B1( u1_u14_u2_n176 ) , .B2( u1_u14_u2_n178 ) );
  OAI221_X1 u1_u14_u2_U41 (.A( u1_u14_u2_n135 ) , .B2( u1_u14_u2_n136 ) , .B1( u1_u14_u2_n137 ) , .ZN( u1_u14_u2_n162 ) , .C2( u1_u14_u2_n167 ) , .C1( u1_u14_u2_n185 ) );
  AND3_X1 u1_u14_u2_U42 (.A3( u1_u14_u2_n131 ) , .A2( u1_u14_u2_n132 ) , .A1( u1_u14_u2_n133 ) , .ZN( u1_u14_u2_n136 ) );
  AOI22_X1 u1_u14_u2_U43 (.ZN( u1_u14_u2_n135 ) , .B1( u1_u14_u2_n140 ) , .A1( u1_u14_u2_n156 ) , .B2( u1_u14_u2_n180 ) , .A2( u1_u14_u2_n188 ) );
  AOI21_X1 u1_u14_u2_U44 (.ZN( u1_u14_u2_n149 ) , .B1( u1_u14_u2_n173 ) , .B2( u1_u14_u2_n188 ) , .A( u1_u14_u2_n95 ) );
  AND3_X1 u1_u14_u2_U45 (.A2( u1_u14_u2_n100 ) , .A1( u1_u14_u2_n104 ) , .A3( u1_u14_u2_n156 ) , .ZN( u1_u14_u2_n95 ) );
  OAI21_X1 u1_u14_u2_U46 (.A( u1_u14_u2_n101 ) , .B2( u1_u14_u2_n121 ) , .B1( u1_u14_u2_n153 ) , .ZN( u1_u14_u2_n164 ) );
  NAND2_X1 u1_u14_u2_U47 (.A2( u1_u14_u2_n100 ) , .A1( u1_u14_u2_n107 ) , .ZN( u1_u14_u2_n155 ) );
  NAND2_X1 u1_u14_u2_U48 (.A2( u1_u14_u2_n105 ) , .A1( u1_u14_u2_n108 ) , .ZN( u1_u14_u2_n143 ) );
  NAND2_X1 u1_u14_u2_U49 (.A1( u1_u14_u2_n104 ) , .A2( u1_u14_u2_n106 ) , .ZN( u1_u14_u2_n152 ) );
  INV_X1 u1_u14_u2_U5 (.A( u1_u14_u2_n150 ) , .ZN( u1_u14_u2_n184 ) );
  NAND2_X1 u1_u14_u2_U50 (.A1( u1_u14_u2_n100 ) , .A2( u1_u14_u2_n105 ) , .ZN( u1_u14_u2_n132 ) );
  INV_X1 u1_u14_u2_U51 (.A( u1_u14_u2_n140 ) , .ZN( u1_u14_u2_n168 ) );
  INV_X1 u1_u14_u2_U52 (.A( u1_u14_u2_n138 ) , .ZN( u1_u14_u2_n167 ) );
  OAI21_X1 u1_u14_u2_U53 (.A( u1_u14_u2_n141 ) , .B2( u1_u14_u2_n142 ) , .ZN( u1_u14_u2_n146 ) , .B1( u1_u14_u2_n153 ) );
  OAI21_X1 u1_u14_u2_U54 (.A( u1_u14_u2_n140 ) , .ZN( u1_u14_u2_n141 ) , .B1( u1_u14_u2_n176 ) , .B2( u1_u14_u2_n177 ) );
  NOR3_X1 u1_u14_u2_U55 (.ZN( u1_u14_u2_n142 ) , .A3( u1_u14_u2_n175 ) , .A2( u1_u14_u2_n178 ) , .A1( u1_u14_u2_n181 ) );
  INV_X1 u1_u14_u2_U56 (.ZN( u1_u14_u2_n187 ) , .A( u1_u14_u2_n99 ) );
  OAI21_X1 u1_u14_u2_U57 (.B1( u1_u14_u2_n137 ) , .B2( u1_u14_u2_n143 ) , .A( u1_u14_u2_n98 ) , .ZN( u1_u14_u2_n99 ) );
  NAND2_X1 u1_u14_u2_U58 (.A1( u1_u14_u2_n102 ) , .A2( u1_u14_u2_n106 ) , .ZN( u1_u14_u2_n113 ) );
  NAND2_X1 u1_u14_u2_U59 (.A1( u1_u14_u2_n106 ) , .A2( u1_u14_u2_n107 ) , .ZN( u1_u14_u2_n131 ) );
  NOR4_X1 u1_u14_u2_U6 (.A4( u1_u14_u2_n124 ) , .A3( u1_u14_u2_n125 ) , .A2( u1_u14_u2_n126 ) , .A1( u1_u14_u2_n127 ) , .ZN( u1_u14_u2_n128 ) );
  NAND2_X1 u1_u14_u2_U60 (.A1( u1_u14_u2_n103 ) , .A2( u1_u14_u2_n107 ) , .ZN( u1_u14_u2_n139 ) );
  NAND2_X1 u1_u14_u2_U61 (.A1( u1_u14_u2_n103 ) , .A2( u1_u14_u2_n105 ) , .ZN( u1_u14_u2_n133 ) );
  NAND2_X1 u1_u14_u2_U62 (.A1( u1_u14_u2_n102 ) , .A2( u1_u14_u2_n103 ) , .ZN( u1_u14_u2_n154 ) );
  NAND2_X1 u1_u14_u2_U63 (.A2( u1_u14_u2_n103 ) , .A1( u1_u14_u2_n104 ) , .ZN( u1_u14_u2_n119 ) );
  NAND2_X1 u1_u14_u2_U64 (.A2( u1_u14_u2_n107 ) , .A1( u1_u14_u2_n108 ) , .ZN( u1_u14_u2_n123 ) );
  NAND2_X1 u1_u14_u2_U65 (.A1( u1_u14_u2_n104 ) , .A2( u1_u14_u2_n108 ) , .ZN( u1_u14_u2_n122 ) );
  INV_X1 u1_u14_u2_U66 (.A( u1_u14_u2_n114 ) , .ZN( u1_u14_u2_n172 ) );
  NAND2_X1 u1_u14_u2_U67 (.A2( u1_u14_u2_n100 ) , .A1( u1_u14_u2_n102 ) , .ZN( u1_u14_u2_n116 ) );
  NAND2_X1 u1_u14_u2_U68 (.A1( u1_u14_u2_n102 ) , .A2( u1_u14_u2_n108 ) , .ZN( u1_u14_u2_n120 ) );
  NAND2_X1 u1_u14_u2_U69 (.A2( u1_u14_u2_n105 ) , .A1( u1_u14_u2_n106 ) , .ZN( u1_u14_u2_n117 ) );
  AOI21_X1 u1_u14_u2_U7 (.B2( u1_u14_u2_n119 ) , .ZN( u1_u14_u2_n127 ) , .A( u1_u14_u2_n137 ) , .B1( u1_u14_u2_n155 ) );
  NOR2_X1 u1_u14_u2_U70 (.A2( u1_u14_X_16 ) , .ZN( u1_u14_u2_n140 ) , .A1( u1_u14_u2_n166 ) );
  NOR2_X1 u1_u14_u2_U71 (.A2( u1_u14_X_13 ) , .A1( u1_u14_X_14 ) , .ZN( u1_u14_u2_n100 ) );
  NOR2_X1 u1_u14_u2_U72 (.A2( u1_u14_X_16 ) , .A1( u1_u14_X_17 ) , .ZN( u1_u14_u2_n138 ) );
  NOR2_X1 u1_u14_u2_U73 (.A2( u1_u14_X_15 ) , .A1( u1_u14_X_18 ) , .ZN( u1_u14_u2_n104 ) );
  NOR2_X1 u1_u14_u2_U74 (.A2( u1_u14_X_14 ) , .ZN( u1_u14_u2_n103 ) , .A1( u1_u14_u2_n174 ) );
  NOR2_X1 u1_u14_u2_U75 (.A2( u1_u14_X_15 ) , .ZN( u1_u14_u2_n102 ) , .A1( u1_u14_u2_n165 ) );
  NOR2_X1 u1_u14_u2_U76 (.A2( u1_u14_X_17 ) , .ZN( u1_u14_u2_n114 ) , .A1( u1_u14_u2_n169 ) );
  AND2_X1 u1_u14_u2_U77 (.A1( u1_u14_X_15 ) , .ZN( u1_u14_u2_n105 ) , .A2( u1_u14_u2_n165 ) );
  AND2_X1 u1_u14_u2_U78 (.A2( u1_u14_X_15 ) , .A1( u1_u14_X_18 ) , .ZN( u1_u14_u2_n107 ) );
  AND2_X1 u1_u14_u2_U79 (.A1( u1_u14_X_14 ) , .ZN( u1_u14_u2_n106 ) , .A2( u1_u14_u2_n174 ) );
  AOI21_X1 u1_u14_u2_U8 (.ZN( u1_u14_u2_n124 ) , .B1( u1_u14_u2_n131 ) , .B2( u1_u14_u2_n143 ) , .A( u1_u14_u2_n172 ) );
  AND2_X1 u1_u14_u2_U80 (.A1( u1_u14_X_13 ) , .A2( u1_u14_X_14 ) , .ZN( u1_u14_u2_n108 ) );
  INV_X1 u1_u14_u2_U81 (.A( u1_u14_X_16 ) , .ZN( u1_u14_u2_n169 ) );
  INV_X1 u1_u14_u2_U82 (.A( u1_u14_X_17 ) , .ZN( u1_u14_u2_n166 ) );
  INV_X1 u1_u14_u2_U83 (.A( u1_u14_X_13 ) , .ZN( u1_u14_u2_n174 ) );
  INV_X1 u1_u14_u2_U84 (.A( u1_u14_X_18 ) , .ZN( u1_u14_u2_n165 ) );
  NAND4_X1 u1_u14_u2_U85 (.ZN( u1_out14_30 ) , .A4( u1_u14_u2_n147 ) , .A3( u1_u14_u2_n148 ) , .A2( u1_u14_u2_n149 ) , .A1( u1_u14_u2_n187 ) );
  NOR3_X1 u1_u14_u2_U86 (.A3( u1_u14_u2_n144 ) , .A2( u1_u14_u2_n145 ) , .A1( u1_u14_u2_n146 ) , .ZN( u1_u14_u2_n147 ) );
  AOI21_X1 u1_u14_u2_U87 (.B2( u1_u14_u2_n138 ) , .ZN( u1_u14_u2_n148 ) , .A( u1_u14_u2_n162 ) , .B1( u1_u14_u2_n182 ) );
  NAND4_X1 u1_u14_u2_U88 (.ZN( u1_out14_24 ) , .A4( u1_u14_u2_n111 ) , .A3( u1_u14_u2_n112 ) , .A1( u1_u14_u2_n130 ) , .A2( u1_u14_u2_n187 ) );
  AOI221_X1 u1_u14_u2_U89 (.A( u1_u14_u2_n109 ) , .B1( u1_u14_u2_n110 ) , .ZN( u1_u14_u2_n111 ) , .C1( u1_u14_u2_n134 ) , .C2( u1_u14_u2_n170 ) , .B2( u1_u14_u2_n173 ) );
  AOI21_X1 u1_u14_u2_U9 (.B2( u1_u14_u2_n123 ) , .ZN( u1_u14_u2_n125 ) , .A( u1_u14_u2_n171 ) , .B1( u1_u14_u2_n184 ) );
  AOI21_X1 u1_u14_u2_U90 (.ZN( u1_u14_u2_n112 ) , .B2( u1_u14_u2_n156 ) , .A( u1_u14_u2_n164 ) , .B1( u1_u14_u2_n181 ) );
  NAND4_X1 u1_u14_u2_U91 (.ZN( u1_out14_16 ) , .A4( u1_u14_u2_n128 ) , .A3( u1_u14_u2_n129 ) , .A1( u1_u14_u2_n130 ) , .A2( u1_u14_u2_n186 ) );
  AOI22_X1 u1_u14_u2_U92 (.A2( u1_u14_u2_n118 ) , .ZN( u1_u14_u2_n129 ) , .A1( u1_u14_u2_n140 ) , .B1( u1_u14_u2_n157 ) , .B2( u1_u14_u2_n170 ) );
  INV_X1 u1_u14_u2_U93 (.A( u1_u14_u2_n163 ) , .ZN( u1_u14_u2_n186 ) );
  OR4_X1 u1_u14_u2_U94 (.ZN( u1_out14_6 ) , .A4( u1_u14_u2_n161 ) , .A3( u1_u14_u2_n162 ) , .A2( u1_u14_u2_n163 ) , .A1( u1_u14_u2_n164 ) );
  OR3_X1 u1_u14_u2_U95 (.A2( u1_u14_u2_n159 ) , .A1( u1_u14_u2_n160 ) , .ZN( u1_u14_u2_n161 ) , .A3( u1_u14_u2_n183 ) );
  AOI21_X1 u1_u14_u2_U96 (.B2( u1_u14_u2_n154 ) , .B1( u1_u14_u2_n155 ) , .ZN( u1_u14_u2_n159 ) , .A( u1_u14_u2_n167 ) );
  NAND3_X1 u1_u14_u2_U97 (.A2( u1_u14_u2_n117 ) , .A1( u1_u14_u2_n122 ) , .A3( u1_u14_u2_n123 ) , .ZN( u1_u14_u2_n134 ) );
  NAND3_X1 u1_u14_u2_U98 (.ZN( u1_u14_u2_n110 ) , .A2( u1_u14_u2_n131 ) , .A3( u1_u14_u2_n139 ) , .A1( u1_u14_u2_n154 ) );
  NAND3_X1 u1_u14_u2_U99 (.A2( u1_u14_u2_n100 ) , .ZN( u1_u14_u2_n101 ) , .A1( u1_u14_u2_n104 ) , .A3( u1_u14_u2_n114 ) );
  OAI22_X1 u1_u14_u3_U10 (.B1( u1_u14_u3_n113 ) , .A2( u1_u14_u3_n135 ) , .A1( u1_u14_u3_n150 ) , .B2( u1_u14_u3_n164 ) , .ZN( u1_u14_u3_n98 ) );
  OAI211_X1 u1_u14_u3_U11 (.B( u1_u14_u3_n106 ) , .ZN( u1_u14_u3_n119 ) , .C2( u1_u14_u3_n128 ) , .C1( u1_u14_u3_n167 ) , .A( u1_u14_u3_n181 ) );
  AOI221_X1 u1_u14_u3_U12 (.C1( u1_u14_u3_n105 ) , .ZN( u1_u14_u3_n106 ) , .A( u1_u14_u3_n131 ) , .B2( u1_u14_u3_n132 ) , .C2( u1_u14_u3_n133 ) , .B1( u1_u14_u3_n169 ) );
  INV_X1 u1_u14_u3_U13 (.ZN( u1_u14_u3_n181 ) , .A( u1_u14_u3_n98 ) );
  NAND2_X1 u1_u14_u3_U14 (.ZN( u1_u14_u3_n105 ) , .A2( u1_u14_u3_n130 ) , .A1( u1_u14_u3_n155 ) );
  AOI22_X1 u1_u14_u3_U15 (.B1( u1_u14_u3_n115 ) , .A2( u1_u14_u3_n116 ) , .ZN( u1_u14_u3_n123 ) , .B2( u1_u14_u3_n133 ) , .A1( u1_u14_u3_n169 ) );
  NAND2_X1 u1_u14_u3_U16 (.ZN( u1_u14_u3_n116 ) , .A2( u1_u14_u3_n151 ) , .A1( u1_u14_u3_n182 ) );
  NOR2_X1 u1_u14_u3_U17 (.ZN( u1_u14_u3_n126 ) , .A2( u1_u14_u3_n150 ) , .A1( u1_u14_u3_n164 ) );
  AOI21_X1 u1_u14_u3_U18 (.ZN( u1_u14_u3_n112 ) , .B2( u1_u14_u3_n146 ) , .B1( u1_u14_u3_n155 ) , .A( u1_u14_u3_n167 ) );
  NAND2_X1 u1_u14_u3_U19 (.A1( u1_u14_u3_n135 ) , .ZN( u1_u14_u3_n142 ) , .A2( u1_u14_u3_n164 ) );
  NAND2_X1 u1_u14_u3_U20 (.ZN( u1_u14_u3_n132 ) , .A2( u1_u14_u3_n152 ) , .A1( u1_u14_u3_n156 ) );
  AND2_X1 u1_u14_u3_U21 (.A2( u1_u14_u3_n113 ) , .A1( u1_u14_u3_n114 ) , .ZN( u1_u14_u3_n151 ) );
  INV_X1 u1_u14_u3_U22 (.A( u1_u14_u3_n133 ) , .ZN( u1_u14_u3_n165 ) );
  INV_X1 u1_u14_u3_U23 (.A( u1_u14_u3_n135 ) , .ZN( u1_u14_u3_n170 ) );
  NAND2_X1 u1_u14_u3_U24 (.A1( u1_u14_u3_n107 ) , .A2( u1_u14_u3_n108 ) , .ZN( u1_u14_u3_n140 ) );
  NAND2_X1 u1_u14_u3_U25 (.ZN( u1_u14_u3_n117 ) , .A1( u1_u14_u3_n124 ) , .A2( u1_u14_u3_n148 ) );
  NAND2_X1 u1_u14_u3_U26 (.ZN( u1_u14_u3_n143 ) , .A1( u1_u14_u3_n165 ) , .A2( u1_u14_u3_n167 ) );
  INV_X1 u1_u14_u3_U27 (.A( u1_u14_u3_n130 ) , .ZN( u1_u14_u3_n177 ) );
  INV_X1 u1_u14_u3_U28 (.A( u1_u14_u3_n128 ) , .ZN( u1_u14_u3_n176 ) );
  INV_X1 u1_u14_u3_U29 (.A( u1_u14_u3_n155 ) , .ZN( u1_u14_u3_n174 ) );
  INV_X1 u1_u14_u3_U3 (.A( u1_u14_u3_n129 ) , .ZN( u1_u14_u3_n183 ) );
  INV_X1 u1_u14_u3_U30 (.A( u1_u14_u3_n139 ) , .ZN( u1_u14_u3_n185 ) );
  NOR2_X1 u1_u14_u3_U31 (.ZN( u1_u14_u3_n135 ) , .A2( u1_u14_u3_n141 ) , .A1( u1_u14_u3_n169 ) );
  OAI222_X1 u1_u14_u3_U32 (.C2( u1_u14_u3_n107 ) , .A2( u1_u14_u3_n108 ) , .B1( u1_u14_u3_n135 ) , .ZN( u1_u14_u3_n138 ) , .B2( u1_u14_u3_n146 ) , .C1( u1_u14_u3_n154 ) , .A1( u1_u14_u3_n164 ) );
  NOR4_X1 u1_u14_u3_U33 (.A4( u1_u14_u3_n157 ) , .A3( u1_u14_u3_n158 ) , .A2( u1_u14_u3_n159 ) , .A1( u1_u14_u3_n160 ) , .ZN( u1_u14_u3_n161 ) );
  AOI21_X1 u1_u14_u3_U34 (.B2( u1_u14_u3_n152 ) , .B1( u1_u14_u3_n153 ) , .ZN( u1_u14_u3_n158 ) , .A( u1_u14_u3_n164 ) );
  AOI21_X1 u1_u14_u3_U35 (.A( u1_u14_u3_n154 ) , .B2( u1_u14_u3_n155 ) , .B1( u1_u14_u3_n156 ) , .ZN( u1_u14_u3_n157 ) );
  AOI21_X1 u1_u14_u3_U36 (.A( u1_u14_u3_n149 ) , .B2( u1_u14_u3_n150 ) , .B1( u1_u14_u3_n151 ) , .ZN( u1_u14_u3_n159 ) );
  AOI211_X1 u1_u14_u3_U37 (.ZN( u1_u14_u3_n109 ) , .A( u1_u14_u3_n119 ) , .C2( u1_u14_u3_n129 ) , .B( u1_u14_u3_n138 ) , .C1( u1_u14_u3_n141 ) );
  AOI211_X1 u1_u14_u3_U38 (.B( u1_u14_u3_n119 ) , .A( u1_u14_u3_n120 ) , .C2( u1_u14_u3_n121 ) , .ZN( u1_u14_u3_n122 ) , .C1( u1_u14_u3_n179 ) );
  INV_X1 u1_u14_u3_U39 (.A( u1_u14_u3_n156 ) , .ZN( u1_u14_u3_n179 ) );
  INV_X1 u1_u14_u3_U4 (.A( u1_u14_u3_n140 ) , .ZN( u1_u14_u3_n182 ) );
  OAI22_X1 u1_u14_u3_U40 (.B1( u1_u14_u3_n118 ) , .ZN( u1_u14_u3_n120 ) , .A1( u1_u14_u3_n135 ) , .B2( u1_u14_u3_n154 ) , .A2( u1_u14_u3_n178 ) );
  AND3_X1 u1_u14_u3_U41 (.ZN( u1_u14_u3_n118 ) , .A2( u1_u14_u3_n124 ) , .A1( u1_u14_u3_n144 ) , .A3( u1_u14_u3_n152 ) );
  INV_X1 u1_u14_u3_U42 (.A( u1_u14_u3_n121 ) , .ZN( u1_u14_u3_n164 ) );
  NAND2_X1 u1_u14_u3_U43 (.ZN( u1_u14_u3_n133 ) , .A1( u1_u14_u3_n154 ) , .A2( u1_u14_u3_n164 ) );
  OAI211_X1 u1_u14_u3_U44 (.B( u1_u14_u3_n127 ) , .ZN( u1_u14_u3_n139 ) , .C1( u1_u14_u3_n150 ) , .C2( u1_u14_u3_n154 ) , .A( u1_u14_u3_n184 ) );
  INV_X1 u1_u14_u3_U45 (.A( u1_u14_u3_n125 ) , .ZN( u1_u14_u3_n184 ) );
  AOI221_X1 u1_u14_u3_U46 (.A( u1_u14_u3_n126 ) , .ZN( u1_u14_u3_n127 ) , .C2( u1_u14_u3_n132 ) , .C1( u1_u14_u3_n169 ) , .B2( u1_u14_u3_n170 ) , .B1( u1_u14_u3_n174 ) );
  OAI22_X1 u1_u14_u3_U47 (.A1( u1_u14_u3_n124 ) , .ZN( u1_u14_u3_n125 ) , .B2( u1_u14_u3_n145 ) , .A2( u1_u14_u3_n165 ) , .B1( u1_u14_u3_n167 ) );
  NOR2_X1 u1_u14_u3_U48 (.A1( u1_u14_u3_n113 ) , .ZN( u1_u14_u3_n131 ) , .A2( u1_u14_u3_n154 ) );
  NAND2_X1 u1_u14_u3_U49 (.A1( u1_u14_u3_n103 ) , .ZN( u1_u14_u3_n150 ) , .A2( u1_u14_u3_n99 ) );
  INV_X1 u1_u14_u3_U5 (.A( u1_u14_u3_n117 ) , .ZN( u1_u14_u3_n178 ) );
  NAND2_X1 u1_u14_u3_U50 (.A2( u1_u14_u3_n102 ) , .ZN( u1_u14_u3_n155 ) , .A1( u1_u14_u3_n97 ) );
  INV_X1 u1_u14_u3_U51 (.A( u1_u14_u3_n141 ) , .ZN( u1_u14_u3_n167 ) );
  AOI21_X1 u1_u14_u3_U52 (.B2( u1_u14_u3_n114 ) , .B1( u1_u14_u3_n146 ) , .A( u1_u14_u3_n154 ) , .ZN( u1_u14_u3_n94 ) );
  AOI21_X1 u1_u14_u3_U53 (.ZN( u1_u14_u3_n110 ) , .B2( u1_u14_u3_n142 ) , .B1( u1_u14_u3_n186 ) , .A( u1_u14_u3_n95 ) );
  INV_X1 u1_u14_u3_U54 (.A( u1_u14_u3_n145 ) , .ZN( u1_u14_u3_n186 ) );
  AOI21_X1 u1_u14_u3_U55 (.B1( u1_u14_u3_n124 ) , .A( u1_u14_u3_n149 ) , .B2( u1_u14_u3_n155 ) , .ZN( u1_u14_u3_n95 ) );
  INV_X1 u1_u14_u3_U56 (.A( u1_u14_u3_n149 ) , .ZN( u1_u14_u3_n169 ) );
  NAND2_X1 u1_u14_u3_U57 (.ZN( u1_u14_u3_n124 ) , .A1( u1_u14_u3_n96 ) , .A2( u1_u14_u3_n97 ) );
  NAND2_X1 u1_u14_u3_U58 (.A2( u1_u14_u3_n100 ) , .ZN( u1_u14_u3_n146 ) , .A1( u1_u14_u3_n96 ) );
  NAND2_X1 u1_u14_u3_U59 (.A1( u1_u14_u3_n101 ) , .ZN( u1_u14_u3_n145 ) , .A2( u1_u14_u3_n99 ) );
  AOI221_X1 u1_u14_u3_U6 (.A( u1_u14_u3_n131 ) , .C2( u1_u14_u3_n132 ) , .C1( u1_u14_u3_n133 ) , .ZN( u1_u14_u3_n134 ) , .B1( u1_u14_u3_n143 ) , .B2( u1_u14_u3_n177 ) );
  NAND2_X1 u1_u14_u3_U60 (.A1( u1_u14_u3_n100 ) , .ZN( u1_u14_u3_n156 ) , .A2( u1_u14_u3_n99 ) );
  NAND2_X1 u1_u14_u3_U61 (.A2( u1_u14_u3_n101 ) , .A1( u1_u14_u3_n104 ) , .ZN( u1_u14_u3_n148 ) );
  NAND2_X1 u1_u14_u3_U62 (.A1( u1_u14_u3_n100 ) , .A2( u1_u14_u3_n102 ) , .ZN( u1_u14_u3_n128 ) );
  NAND2_X1 u1_u14_u3_U63 (.A2( u1_u14_u3_n101 ) , .A1( u1_u14_u3_n102 ) , .ZN( u1_u14_u3_n152 ) );
  NAND2_X1 u1_u14_u3_U64 (.A2( u1_u14_u3_n101 ) , .ZN( u1_u14_u3_n114 ) , .A1( u1_u14_u3_n96 ) );
  NAND2_X1 u1_u14_u3_U65 (.ZN( u1_u14_u3_n107 ) , .A1( u1_u14_u3_n97 ) , .A2( u1_u14_u3_n99 ) );
  NAND2_X1 u1_u14_u3_U66 (.A2( u1_u14_u3_n100 ) , .A1( u1_u14_u3_n104 ) , .ZN( u1_u14_u3_n113 ) );
  NAND2_X1 u1_u14_u3_U67 (.A1( u1_u14_u3_n104 ) , .ZN( u1_u14_u3_n153 ) , .A2( u1_u14_u3_n97 ) );
  NAND2_X1 u1_u14_u3_U68 (.A2( u1_u14_u3_n103 ) , .A1( u1_u14_u3_n104 ) , .ZN( u1_u14_u3_n130 ) );
  NAND2_X1 u1_u14_u3_U69 (.A2( u1_u14_u3_n103 ) , .ZN( u1_u14_u3_n144 ) , .A1( u1_u14_u3_n96 ) );
  OAI22_X1 u1_u14_u3_U7 (.B2( u1_u14_u3_n147 ) , .A2( u1_u14_u3_n148 ) , .ZN( u1_u14_u3_n160 ) , .B1( u1_u14_u3_n165 ) , .A1( u1_u14_u3_n168 ) );
  NAND2_X1 u1_u14_u3_U70 (.A1( u1_u14_u3_n102 ) , .A2( u1_u14_u3_n103 ) , .ZN( u1_u14_u3_n108 ) );
  NOR2_X1 u1_u14_u3_U71 (.A2( u1_u14_X_19 ) , .A1( u1_u14_X_20 ) , .ZN( u1_u14_u3_n99 ) );
  NOR2_X1 u1_u14_u3_U72 (.A2( u1_u14_X_21 ) , .A1( u1_u14_X_24 ) , .ZN( u1_u14_u3_n103 ) );
  NOR2_X1 u1_u14_u3_U73 (.A2( u1_u14_X_24 ) , .A1( u1_u14_u3_n171 ) , .ZN( u1_u14_u3_n97 ) );
  NOR2_X1 u1_u14_u3_U74 (.A2( u1_u14_X_23 ) , .ZN( u1_u14_u3_n141 ) , .A1( u1_u14_u3_n166 ) );
  NOR2_X1 u1_u14_u3_U75 (.A2( u1_u14_X_19 ) , .A1( u1_u14_u3_n172 ) , .ZN( u1_u14_u3_n96 ) );
  NAND2_X1 u1_u14_u3_U76 (.A1( u1_u14_X_22 ) , .A2( u1_u14_X_23 ) , .ZN( u1_u14_u3_n154 ) );
  NAND2_X1 u1_u14_u3_U77 (.A1( u1_u14_X_23 ) , .ZN( u1_u14_u3_n149 ) , .A2( u1_u14_u3_n166 ) );
  NOR2_X1 u1_u14_u3_U78 (.A2( u1_u14_X_22 ) , .A1( u1_u14_X_23 ) , .ZN( u1_u14_u3_n121 ) );
  AND2_X1 u1_u14_u3_U79 (.A1( u1_u14_X_24 ) , .ZN( u1_u14_u3_n101 ) , .A2( u1_u14_u3_n171 ) );
  AND3_X1 u1_u14_u3_U8 (.A3( u1_u14_u3_n144 ) , .A2( u1_u14_u3_n145 ) , .A1( u1_u14_u3_n146 ) , .ZN( u1_u14_u3_n147 ) );
  AND2_X1 u1_u14_u3_U80 (.A1( u1_u14_X_19 ) , .ZN( u1_u14_u3_n102 ) , .A2( u1_u14_u3_n172 ) );
  AND2_X1 u1_u14_u3_U81 (.A1( u1_u14_X_21 ) , .A2( u1_u14_X_24 ) , .ZN( u1_u14_u3_n100 ) );
  AND2_X1 u1_u14_u3_U82 (.A2( u1_u14_X_19 ) , .A1( u1_u14_X_20 ) , .ZN( u1_u14_u3_n104 ) );
  INV_X1 u1_u14_u3_U83 (.A( u1_u14_X_22 ) , .ZN( u1_u14_u3_n166 ) );
  INV_X1 u1_u14_u3_U84 (.A( u1_u14_X_21 ) , .ZN( u1_u14_u3_n171 ) );
  INV_X1 u1_u14_u3_U85 (.A( u1_u14_X_20 ) , .ZN( u1_u14_u3_n172 ) );
  NAND4_X1 u1_u14_u3_U86 (.ZN( u1_out14_26 ) , .A4( u1_u14_u3_n109 ) , .A3( u1_u14_u3_n110 ) , .A2( u1_u14_u3_n111 ) , .A1( u1_u14_u3_n173 ) );
  INV_X1 u1_u14_u3_U87 (.ZN( u1_u14_u3_n173 ) , .A( u1_u14_u3_n94 ) );
  OAI21_X1 u1_u14_u3_U88 (.ZN( u1_u14_u3_n111 ) , .B2( u1_u14_u3_n117 ) , .A( u1_u14_u3_n133 ) , .B1( u1_u14_u3_n176 ) );
  NAND4_X1 u1_u14_u3_U89 (.ZN( u1_out14_20 ) , .A4( u1_u14_u3_n122 ) , .A3( u1_u14_u3_n123 ) , .A1( u1_u14_u3_n175 ) , .A2( u1_u14_u3_n180 ) );
  INV_X1 u1_u14_u3_U9 (.A( u1_u14_u3_n143 ) , .ZN( u1_u14_u3_n168 ) );
  INV_X1 u1_u14_u3_U90 (.A( u1_u14_u3_n126 ) , .ZN( u1_u14_u3_n180 ) );
  INV_X1 u1_u14_u3_U91 (.A( u1_u14_u3_n112 ) , .ZN( u1_u14_u3_n175 ) );
  NAND4_X1 u1_u14_u3_U92 (.ZN( u1_out14_1 ) , .A4( u1_u14_u3_n161 ) , .A3( u1_u14_u3_n162 ) , .A2( u1_u14_u3_n163 ) , .A1( u1_u14_u3_n185 ) );
  NAND2_X1 u1_u14_u3_U93 (.ZN( u1_u14_u3_n163 ) , .A2( u1_u14_u3_n170 ) , .A1( u1_u14_u3_n176 ) );
  AOI22_X1 u1_u14_u3_U94 (.B2( u1_u14_u3_n140 ) , .B1( u1_u14_u3_n141 ) , .A2( u1_u14_u3_n142 ) , .ZN( u1_u14_u3_n162 ) , .A1( u1_u14_u3_n177 ) );
  OR4_X1 u1_u14_u3_U95 (.ZN( u1_out14_10 ) , .A4( u1_u14_u3_n136 ) , .A3( u1_u14_u3_n137 ) , .A1( u1_u14_u3_n138 ) , .A2( u1_u14_u3_n139 ) );
  OAI222_X1 u1_u14_u3_U96 (.C1( u1_u14_u3_n128 ) , .ZN( u1_u14_u3_n137 ) , .B1( u1_u14_u3_n148 ) , .A2( u1_u14_u3_n150 ) , .B2( u1_u14_u3_n154 ) , .C2( u1_u14_u3_n164 ) , .A1( u1_u14_u3_n167 ) );
  OAI221_X1 u1_u14_u3_U97 (.A( u1_u14_u3_n134 ) , .B2( u1_u14_u3_n135 ) , .ZN( u1_u14_u3_n136 ) , .C1( u1_u14_u3_n149 ) , .B1( u1_u14_u3_n151 ) , .C2( u1_u14_u3_n183 ) );
  NAND3_X1 u1_u14_u3_U98 (.A1( u1_u14_u3_n114 ) , .ZN( u1_u14_u3_n115 ) , .A2( u1_u14_u3_n145 ) , .A3( u1_u14_u3_n153 ) );
  NAND3_X1 u1_u14_u3_U99 (.ZN( u1_u14_u3_n129 ) , .A2( u1_u14_u3_n144 ) , .A1( u1_u14_u3_n153 ) , .A3( u1_u14_u3_n182 ) );
  OAI22_X1 u1_u14_u4_U10 (.B2( u1_u14_u4_n135 ) , .ZN( u1_u14_u4_n137 ) , .B1( u1_u14_u4_n153 ) , .A1( u1_u14_u4_n155 ) , .A2( u1_u14_u4_n171 ) );
  AND3_X1 u1_u14_u4_U11 (.A2( u1_u14_u4_n134 ) , .ZN( u1_u14_u4_n135 ) , .A3( u1_u14_u4_n145 ) , .A1( u1_u14_u4_n157 ) );
  NAND2_X1 u1_u14_u4_U12 (.ZN( u1_u14_u4_n132 ) , .A2( u1_u14_u4_n170 ) , .A1( u1_u14_u4_n173 ) );
  AOI21_X1 u1_u14_u4_U13 (.B2( u1_u14_u4_n160 ) , .B1( u1_u14_u4_n161 ) , .ZN( u1_u14_u4_n162 ) , .A( u1_u14_u4_n170 ) );
  AOI21_X1 u1_u14_u4_U14 (.ZN( u1_u14_u4_n107 ) , .B2( u1_u14_u4_n143 ) , .A( u1_u14_u4_n174 ) , .B1( u1_u14_u4_n184 ) );
  AOI21_X1 u1_u14_u4_U15 (.B2( u1_u14_u4_n158 ) , .B1( u1_u14_u4_n159 ) , .ZN( u1_u14_u4_n163 ) , .A( u1_u14_u4_n174 ) );
  AOI21_X1 u1_u14_u4_U16 (.A( u1_u14_u4_n153 ) , .B2( u1_u14_u4_n154 ) , .B1( u1_u14_u4_n155 ) , .ZN( u1_u14_u4_n165 ) );
  AOI21_X1 u1_u14_u4_U17 (.A( u1_u14_u4_n156 ) , .B2( u1_u14_u4_n157 ) , .ZN( u1_u14_u4_n164 ) , .B1( u1_u14_u4_n184 ) );
  INV_X1 u1_u14_u4_U18 (.A( u1_u14_u4_n138 ) , .ZN( u1_u14_u4_n170 ) );
  AND2_X1 u1_u14_u4_U19 (.A2( u1_u14_u4_n120 ) , .ZN( u1_u14_u4_n155 ) , .A1( u1_u14_u4_n160 ) );
  INV_X1 u1_u14_u4_U20 (.A( u1_u14_u4_n156 ) , .ZN( u1_u14_u4_n175 ) );
  NAND2_X1 u1_u14_u4_U21 (.A2( u1_u14_u4_n118 ) , .ZN( u1_u14_u4_n131 ) , .A1( u1_u14_u4_n147 ) );
  NAND2_X1 u1_u14_u4_U22 (.A1( u1_u14_u4_n119 ) , .A2( u1_u14_u4_n120 ) , .ZN( u1_u14_u4_n130 ) );
  NAND2_X1 u1_u14_u4_U23 (.ZN( u1_u14_u4_n117 ) , .A2( u1_u14_u4_n118 ) , .A1( u1_u14_u4_n148 ) );
  NAND2_X1 u1_u14_u4_U24 (.ZN( u1_u14_u4_n129 ) , .A1( u1_u14_u4_n134 ) , .A2( u1_u14_u4_n148 ) );
  AND3_X1 u1_u14_u4_U25 (.A1( u1_u14_u4_n119 ) , .A2( u1_u14_u4_n143 ) , .A3( u1_u14_u4_n154 ) , .ZN( u1_u14_u4_n161 ) );
  AND2_X1 u1_u14_u4_U26 (.A1( u1_u14_u4_n145 ) , .A2( u1_u14_u4_n147 ) , .ZN( u1_u14_u4_n159 ) );
  OR3_X1 u1_u14_u4_U27 (.A3( u1_u14_u4_n114 ) , .A2( u1_u14_u4_n115 ) , .A1( u1_u14_u4_n116 ) , .ZN( u1_u14_u4_n136 ) );
  AOI21_X1 u1_u14_u4_U28 (.A( u1_u14_u4_n113 ) , .ZN( u1_u14_u4_n116 ) , .B2( u1_u14_u4_n173 ) , .B1( u1_u14_u4_n174 ) );
  AOI21_X1 u1_u14_u4_U29 (.ZN( u1_u14_u4_n115 ) , .B2( u1_u14_u4_n145 ) , .B1( u1_u14_u4_n146 ) , .A( u1_u14_u4_n156 ) );
  NOR2_X1 u1_u14_u4_U3 (.ZN( u1_u14_u4_n121 ) , .A1( u1_u14_u4_n181 ) , .A2( u1_u14_u4_n182 ) );
  OAI22_X1 u1_u14_u4_U30 (.ZN( u1_u14_u4_n114 ) , .A2( u1_u14_u4_n121 ) , .B1( u1_u14_u4_n160 ) , .B2( u1_u14_u4_n170 ) , .A1( u1_u14_u4_n171 ) );
  INV_X1 u1_u14_u4_U31 (.A( u1_u14_u4_n158 ) , .ZN( u1_u14_u4_n182 ) );
  INV_X1 u1_u14_u4_U32 (.ZN( u1_u14_u4_n181 ) , .A( u1_u14_u4_n96 ) );
  INV_X1 u1_u14_u4_U33 (.A( u1_u14_u4_n144 ) , .ZN( u1_u14_u4_n179 ) );
  INV_X1 u1_u14_u4_U34 (.A( u1_u14_u4_n157 ) , .ZN( u1_u14_u4_n178 ) );
  NAND2_X1 u1_u14_u4_U35 (.A2( u1_u14_u4_n154 ) , .A1( u1_u14_u4_n96 ) , .ZN( u1_u14_u4_n97 ) );
  INV_X1 u1_u14_u4_U36 (.ZN( u1_u14_u4_n186 ) , .A( u1_u14_u4_n95 ) );
  OAI221_X1 u1_u14_u4_U37 (.C1( u1_u14_u4_n134 ) , .B1( u1_u14_u4_n158 ) , .B2( u1_u14_u4_n171 ) , .C2( u1_u14_u4_n173 ) , .A( u1_u14_u4_n94 ) , .ZN( u1_u14_u4_n95 ) );
  AOI222_X1 u1_u14_u4_U38 (.B2( u1_u14_u4_n132 ) , .A1( u1_u14_u4_n138 ) , .C2( u1_u14_u4_n175 ) , .A2( u1_u14_u4_n179 ) , .C1( u1_u14_u4_n181 ) , .B1( u1_u14_u4_n185 ) , .ZN( u1_u14_u4_n94 ) );
  INV_X1 u1_u14_u4_U39 (.A( u1_u14_u4_n113 ) , .ZN( u1_u14_u4_n185 ) );
  INV_X1 u1_u14_u4_U4 (.A( u1_u14_u4_n117 ) , .ZN( u1_u14_u4_n184 ) );
  INV_X1 u1_u14_u4_U40 (.A( u1_u14_u4_n143 ) , .ZN( u1_u14_u4_n183 ) );
  NOR2_X1 u1_u14_u4_U41 (.ZN( u1_u14_u4_n138 ) , .A1( u1_u14_u4_n168 ) , .A2( u1_u14_u4_n169 ) );
  NOR2_X1 u1_u14_u4_U42 (.A1( u1_u14_u4_n150 ) , .A2( u1_u14_u4_n152 ) , .ZN( u1_u14_u4_n153 ) );
  NOR2_X1 u1_u14_u4_U43 (.A2( u1_u14_u4_n128 ) , .A1( u1_u14_u4_n138 ) , .ZN( u1_u14_u4_n156 ) );
  AOI22_X1 u1_u14_u4_U44 (.B2( u1_u14_u4_n122 ) , .A1( u1_u14_u4_n123 ) , .ZN( u1_u14_u4_n124 ) , .B1( u1_u14_u4_n128 ) , .A2( u1_u14_u4_n172 ) );
  INV_X1 u1_u14_u4_U45 (.A( u1_u14_u4_n153 ) , .ZN( u1_u14_u4_n172 ) );
  NAND2_X1 u1_u14_u4_U46 (.A2( u1_u14_u4_n120 ) , .ZN( u1_u14_u4_n123 ) , .A1( u1_u14_u4_n161 ) );
  AOI22_X1 u1_u14_u4_U47 (.B2( u1_u14_u4_n132 ) , .A2( u1_u14_u4_n133 ) , .ZN( u1_u14_u4_n140 ) , .A1( u1_u14_u4_n150 ) , .B1( u1_u14_u4_n179 ) );
  NAND2_X1 u1_u14_u4_U48 (.ZN( u1_u14_u4_n133 ) , .A2( u1_u14_u4_n146 ) , .A1( u1_u14_u4_n154 ) );
  NAND2_X1 u1_u14_u4_U49 (.A1( u1_u14_u4_n103 ) , .ZN( u1_u14_u4_n154 ) , .A2( u1_u14_u4_n98 ) );
  NOR4_X1 u1_u14_u4_U5 (.A4( u1_u14_u4_n106 ) , .A3( u1_u14_u4_n107 ) , .A2( u1_u14_u4_n108 ) , .A1( u1_u14_u4_n109 ) , .ZN( u1_u14_u4_n110 ) );
  NAND2_X1 u1_u14_u4_U50 (.A1( u1_u14_u4_n101 ) , .ZN( u1_u14_u4_n158 ) , .A2( u1_u14_u4_n99 ) );
  AOI21_X1 u1_u14_u4_U51 (.ZN( u1_u14_u4_n127 ) , .A( u1_u14_u4_n136 ) , .B2( u1_u14_u4_n150 ) , .B1( u1_u14_u4_n180 ) );
  INV_X1 u1_u14_u4_U52 (.A( u1_u14_u4_n160 ) , .ZN( u1_u14_u4_n180 ) );
  NAND2_X1 u1_u14_u4_U53 (.A2( u1_u14_u4_n104 ) , .A1( u1_u14_u4_n105 ) , .ZN( u1_u14_u4_n146 ) );
  NAND2_X1 u1_u14_u4_U54 (.A2( u1_u14_u4_n101 ) , .A1( u1_u14_u4_n102 ) , .ZN( u1_u14_u4_n160 ) );
  NAND2_X1 u1_u14_u4_U55 (.ZN( u1_u14_u4_n134 ) , .A1( u1_u14_u4_n98 ) , .A2( u1_u14_u4_n99 ) );
  NAND2_X1 u1_u14_u4_U56 (.A1( u1_u14_u4_n103 ) , .A2( u1_u14_u4_n104 ) , .ZN( u1_u14_u4_n143 ) );
  NAND2_X1 u1_u14_u4_U57 (.A2( u1_u14_u4_n105 ) , .ZN( u1_u14_u4_n145 ) , .A1( u1_u14_u4_n98 ) );
  NAND2_X1 u1_u14_u4_U58 (.A1( u1_u14_u4_n100 ) , .A2( u1_u14_u4_n105 ) , .ZN( u1_u14_u4_n120 ) );
  NAND2_X1 u1_u14_u4_U59 (.A1( u1_u14_u4_n102 ) , .A2( u1_u14_u4_n104 ) , .ZN( u1_u14_u4_n148 ) );
  AOI21_X1 u1_u14_u4_U6 (.ZN( u1_u14_u4_n106 ) , .B2( u1_u14_u4_n146 ) , .B1( u1_u14_u4_n158 ) , .A( u1_u14_u4_n170 ) );
  NAND2_X1 u1_u14_u4_U60 (.A2( u1_u14_u4_n100 ) , .A1( u1_u14_u4_n103 ) , .ZN( u1_u14_u4_n157 ) );
  INV_X1 u1_u14_u4_U61 (.A( u1_u14_u4_n150 ) , .ZN( u1_u14_u4_n173 ) );
  INV_X1 u1_u14_u4_U62 (.A( u1_u14_u4_n152 ) , .ZN( u1_u14_u4_n171 ) );
  NAND2_X1 u1_u14_u4_U63 (.A1( u1_u14_u4_n100 ) , .ZN( u1_u14_u4_n118 ) , .A2( u1_u14_u4_n99 ) );
  NAND2_X1 u1_u14_u4_U64 (.A2( u1_u14_u4_n100 ) , .A1( u1_u14_u4_n102 ) , .ZN( u1_u14_u4_n144 ) );
  NAND2_X1 u1_u14_u4_U65 (.A2( u1_u14_u4_n101 ) , .A1( u1_u14_u4_n105 ) , .ZN( u1_u14_u4_n96 ) );
  INV_X1 u1_u14_u4_U66 (.A( u1_u14_u4_n128 ) , .ZN( u1_u14_u4_n174 ) );
  NAND2_X1 u1_u14_u4_U67 (.A2( u1_u14_u4_n102 ) , .ZN( u1_u14_u4_n119 ) , .A1( u1_u14_u4_n98 ) );
  NAND2_X1 u1_u14_u4_U68 (.A2( u1_u14_u4_n101 ) , .A1( u1_u14_u4_n103 ) , .ZN( u1_u14_u4_n147 ) );
  NAND2_X1 u1_u14_u4_U69 (.A2( u1_u14_u4_n104 ) , .ZN( u1_u14_u4_n113 ) , .A1( u1_u14_u4_n99 ) );
  AOI21_X1 u1_u14_u4_U7 (.ZN( u1_u14_u4_n108 ) , .B2( u1_u14_u4_n134 ) , .B1( u1_u14_u4_n155 ) , .A( u1_u14_u4_n156 ) );
  NOR2_X1 u1_u14_u4_U70 (.A2( u1_u14_X_28 ) , .ZN( u1_u14_u4_n150 ) , .A1( u1_u14_u4_n168 ) );
  NOR2_X1 u1_u14_u4_U71 (.A2( u1_u14_X_29 ) , .ZN( u1_u14_u4_n152 ) , .A1( u1_u14_u4_n169 ) );
  NOR2_X1 u1_u14_u4_U72 (.A2( u1_u14_X_30 ) , .ZN( u1_u14_u4_n105 ) , .A1( u1_u14_u4_n176 ) );
  NOR2_X1 u1_u14_u4_U73 (.A2( u1_u14_X_26 ) , .ZN( u1_u14_u4_n100 ) , .A1( u1_u14_u4_n177 ) );
  NOR2_X1 u1_u14_u4_U74 (.A2( u1_u14_X_28 ) , .A1( u1_u14_X_29 ) , .ZN( u1_u14_u4_n128 ) );
  NOR2_X1 u1_u14_u4_U75 (.A2( u1_u14_X_27 ) , .A1( u1_u14_X_30 ) , .ZN( u1_u14_u4_n102 ) );
  NOR2_X1 u1_u14_u4_U76 (.A2( u1_u14_X_25 ) , .A1( u1_u14_X_26 ) , .ZN( u1_u14_u4_n98 ) );
  AND2_X1 u1_u14_u4_U77 (.A2( u1_u14_X_25 ) , .A1( u1_u14_X_26 ) , .ZN( u1_u14_u4_n104 ) );
  AND2_X1 u1_u14_u4_U78 (.A1( u1_u14_X_30 ) , .A2( u1_u14_u4_n176 ) , .ZN( u1_u14_u4_n99 ) );
  AND2_X1 u1_u14_u4_U79 (.A1( u1_u14_X_26 ) , .ZN( u1_u14_u4_n101 ) , .A2( u1_u14_u4_n177 ) );
  AOI21_X1 u1_u14_u4_U8 (.ZN( u1_u14_u4_n109 ) , .A( u1_u14_u4_n153 ) , .B1( u1_u14_u4_n159 ) , .B2( u1_u14_u4_n184 ) );
  AND2_X1 u1_u14_u4_U80 (.A1( u1_u14_X_27 ) , .A2( u1_u14_X_30 ) , .ZN( u1_u14_u4_n103 ) );
  INV_X1 u1_u14_u4_U81 (.A( u1_u14_X_28 ) , .ZN( u1_u14_u4_n169 ) );
  INV_X1 u1_u14_u4_U82 (.A( u1_u14_X_29 ) , .ZN( u1_u14_u4_n168 ) );
  INV_X1 u1_u14_u4_U83 (.A( u1_u14_X_25 ) , .ZN( u1_u14_u4_n177 ) );
  INV_X1 u1_u14_u4_U84 (.A( u1_u14_X_27 ) , .ZN( u1_u14_u4_n176 ) );
  NAND4_X1 u1_u14_u4_U85 (.ZN( u1_out14_25 ) , .A4( u1_u14_u4_n139 ) , .A3( u1_u14_u4_n140 ) , .A2( u1_u14_u4_n141 ) , .A1( u1_u14_u4_n142 ) );
  OAI21_X1 u1_u14_u4_U86 (.A( u1_u14_u4_n128 ) , .B2( u1_u14_u4_n129 ) , .B1( u1_u14_u4_n130 ) , .ZN( u1_u14_u4_n142 ) );
  OAI21_X1 u1_u14_u4_U87 (.B2( u1_u14_u4_n131 ) , .ZN( u1_u14_u4_n141 ) , .A( u1_u14_u4_n175 ) , .B1( u1_u14_u4_n183 ) );
  NAND4_X1 u1_u14_u4_U88 (.ZN( u1_out14_14 ) , .A4( u1_u14_u4_n124 ) , .A3( u1_u14_u4_n125 ) , .A2( u1_u14_u4_n126 ) , .A1( u1_u14_u4_n127 ) );
  AOI22_X1 u1_u14_u4_U89 (.B2( u1_u14_u4_n117 ) , .ZN( u1_u14_u4_n126 ) , .A1( u1_u14_u4_n129 ) , .B1( u1_u14_u4_n152 ) , .A2( u1_u14_u4_n175 ) );
  AOI211_X1 u1_u14_u4_U9 (.B( u1_u14_u4_n136 ) , .A( u1_u14_u4_n137 ) , .C2( u1_u14_u4_n138 ) , .ZN( u1_u14_u4_n139 ) , .C1( u1_u14_u4_n182 ) );
  AOI22_X1 u1_u14_u4_U90 (.ZN( u1_u14_u4_n125 ) , .B2( u1_u14_u4_n131 ) , .A2( u1_u14_u4_n132 ) , .B1( u1_u14_u4_n138 ) , .A1( u1_u14_u4_n178 ) );
  NAND4_X1 u1_u14_u4_U91 (.ZN( u1_out14_8 ) , .A4( u1_u14_u4_n110 ) , .A3( u1_u14_u4_n111 ) , .A2( u1_u14_u4_n112 ) , .A1( u1_u14_u4_n186 ) );
  NAND2_X1 u1_u14_u4_U92 (.ZN( u1_u14_u4_n112 ) , .A2( u1_u14_u4_n130 ) , .A1( u1_u14_u4_n150 ) );
  AOI22_X1 u1_u14_u4_U93 (.ZN( u1_u14_u4_n111 ) , .B2( u1_u14_u4_n132 ) , .A1( u1_u14_u4_n152 ) , .B1( u1_u14_u4_n178 ) , .A2( u1_u14_u4_n97 ) );
  AOI22_X1 u1_u14_u4_U94 (.B2( u1_u14_u4_n149 ) , .B1( u1_u14_u4_n150 ) , .A2( u1_u14_u4_n151 ) , .A1( u1_u14_u4_n152 ) , .ZN( u1_u14_u4_n167 ) );
  NOR4_X1 u1_u14_u4_U95 (.A4( u1_u14_u4_n162 ) , .A3( u1_u14_u4_n163 ) , .A2( u1_u14_u4_n164 ) , .A1( u1_u14_u4_n165 ) , .ZN( u1_u14_u4_n166 ) );
  NAND3_X1 u1_u14_u4_U96 (.ZN( u1_out14_3 ) , .A3( u1_u14_u4_n166 ) , .A1( u1_u14_u4_n167 ) , .A2( u1_u14_u4_n186 ) );
  NAND3_X1 u1_u14_u4_U97 (.A3( u1_u14_u4_n146 ) , .A2( u1_u14_u4_n147 ) , .A1( u1_u14_u4_n148 ) , .ZN( u1_u14_u4_n149 ) );
  NAND3_X1 u1_u14_u4_U98 (.A3( u1_u14_u4_n143 ) , .A2( u1_u14_u4_n144 ) , .A1( u1_u14_u4_n145 ) , .ZN( u1_u14_u4_n151 ) );
  NAND3_X1 u1_u14_u4_U99 (.A3( u1_u14_u4_n121 ) , .ZN( u1_u14_u4_n122 ) , .A2( u1_u14_u4_n144 ) , .A1( u1_u14_u4_n154 ) );
  XOR2_X1 u1_u15_U10 (.A( u1_FP_62 ) , .B( u1_K16_45 ) , .Z( u1_u15_X_45 ) );
  XOR2_X1 u1_u15_U11 (.A( u1_FP_61 ) , .B( u1_K16_44 ) , .Z( u1_u15_X_44 ) );
  XOR2_X1 u1_u15_U12 (.A( u1_FP_60 ) , .B( u1_K16_43 ) , .Z( u1_u15_X_43 ) );
  XOR2_X1 u1_u15_U13 (.A( u1_FP_61 ) , .B( u1_K16_42 ) , .Z( u1_u15_X_42 ) );
  XOR2_X1 u1_u15_U14 (.A( u1_FP_60 ) , .B( u1_K16_41 ) , .Z( u1_u15_X_41 ) );
  XOR2_X1 u1_u15_U15 (.A( u1_FP_59 ) , .B( u1_K16_40 ) , .Z( u1_u15_X_40 ) );
  XOR2_X1 u1_u15_U17 (.A( u1_FP_58 ) , .B( u1_K16_39 ) , .Z( u1_u15_X_39 ) );
  XOR2_X1 u1_u15_U18 (.A( u1_FP_57 ) , .B( u1_K16_38 ) , .Z( u1_u15_X_38 ) );
  XOR2_X1 u1_u15_U19 (.A( u1_FP_56 ) , .B( u1_K16_37 ) , .Z( u1_u15_X_37 ) );
  XOR2_X1 u1_u15_U20 (.A( u1_FP_57 ) , .B( u1_K16_36 ) , .Z( u1_u15_X_36 ) );
  XOR2_X1 u1_u15_U21 (.A( u1_FP_56 ) , .B( u1_K16_35 ) , .Z( u1_u15_X_35 ) );
  XOR2_X1 u1_u15_U22 (.A( u1_FP_55 ) , .B( u1_K16_34 ) , .Z( u1_u15_X_34 ) );
  XOR2_X1 u1_u15_U23 (.A( u1_FP_54 ) , .B( u1_K16_33 ) , .Z( u1_u15_X_33 ) );
  XOR2_X1 u1_u15_U24 (.A( u1_FP_53 ) , .B( u1_K16_32 ) , .Z( u1_u15_X_32 ) );
  XOR2_X1 u1_u15_U25 (.A( u1_FP_52 ) , .B( u1_K16_31 ) , .Z( u1_u15_X_31 ) );
  XOR2_X1 u1_u15_U26 (.A( u1_FP_53 ) , .B( u1_K16_30 ) , .Z( u1_u15_X_30 ) );
  XOR2_X1 u1_u15_U28 (.A( u1_FP_52 ) , .B( u1_K16_29 ) , .Z( u1_u15_X_29 ) );
  XOR2_X1 u1_u15_U29 (.A( u1_FP_51 ) , .B( u1_K16_28 ) , .Z( u1_u15_X_28 ) );
  XOR2_X1 u1_u15_U30 (.A( u1_FP_50 ) , .B( u1_K16_27 ) , .Z( u1_u15_X_27 ) );
  XOR2_X1 u1_u15_U31 (.A( u1_FP_49 ) , .B( u1_K16_26 ) , .Z( u1_u15_X_26 ) );
  XOR2_X1 u1_u15_U32 (.A( u1_FP_48 ) , .B( u1_K16_25 ) , .Z( u1_u15_X_25 ) );
  XOR2_X1 u1_u15_U7 (.A( u1_FP_33 ) , .B( u1_K16_48 ) , .Z( u1_u15_X_48 ) );
  XOR2_X1 u1_u15_U8 (.A( u1_FP_64 ) , .B( u1_K16_47 ) , .Z( u1_u15_X_47 ) );
  XOR2_X1 u1_u15_U9 (.A( u1_FP_63 ) , .B( u1_K16_46 ) , .Z( u1_u15_X_46 ) );
  OAI22_X1 u1_u15_u4_U10 (.B2( u1_u15_u4_n135 ) , .ZN( u1_u15_u4_n137 ) , .B1( u1_u15_u4_n153 ) , .A1( u1_u15_u4_n155 ) , .A2( u1_u15_u4_n171 ) );
  AND3_X1 u1_u15_u4_U11 (.A2( u1_u15_u4_n134 ) , .ZN( u1_u15_u4_n135 ) , .A3( u1_u15_u4_n145 ) , .A1( u1_u15_u4_n157 ) );
  NAND2_X1 u1_u15_u4_U12 (.ZN( u1_u15_u4_n132 ) , .A2( u1_u15_u4_n170 ) , .A1( u1_u15_u4_n173 ) );
  AOI21_X1 u1_u15_u4_U13 (.B2( u1_u15_u4_n160 ) , .B1( u1_u15_u4_n161 ) , .ZN( u1_u15_u4_n162 ) , .A( u1_u15_u4_n170 ) );
  AOI21_X1 u1_u15_u4_U14 (.ZN( u1_u15_u4_n107 ) , .B2( u1_u15_u4_n143 ) , .A( u1_u15_u4_n174 ) , .B1( u1_u15_u4_n184 ) );
  AOI21_X1 u1_u15_u4_U15 (.B2( u1_u15_u4_n158 ) , .B1( u1_u15_u4_n159 ) , .ZN( u1_u15_u4_n163 ) , .A( u1_u15_u4_n174 ) );
  AOI21_X1 u1_u15_u4_U16 (.A( u1_u15_u4_n153 ) , .B2( u1_u15_u4_n154 ) , .B1( u1_u15_u4_n155 ) , .ZN( u1_u15_u4_n165 ) );
  AOI21_X1 u1_u15_u4_U17 (.A( u1_u15_u4_n156 ) , .B2( u1_u15_u4_n157 ) , .ZN( u1_u15_u4_n164 ) , .B1( u1_u15_u4_n184 ) );
  INV_X1 u1_u15_u4_U18 (.A( u1_u15_u4_n138 ) , .ZN( u1_u15_u4_n170 ) );
  AND2_X1 u1_u15_u4_U19 (.A2( u1_u15_u4_n120 ) , .ZN( u1_u15_u4_n155 ) , .A1( u1_u15_u4_n160 ) );
  INV_X1 u1_u15_u4_U20 (.A( u1_u15_u4_n156 ) , .ZN( u1_u15_u4_n175 ) );
  NAND2_X1 u1_u15_u4_U21 (.A2( u1_u15_u4_n118 ) , .ZN( u1_u15_u4_n131 ) , .A1( u1_u15_u4_n147 ) );
  NAND2_X1 u1_u15_u4_U22 (.A1( u1_u15_u4_n119 ) , .A2( u1_u15_u4_n120 ) , .ZN( u1_u15_u4_n130 ) );
  NAND2_X1 u1_u15_u4_U23 (.ZN( u1_u15_u4_n117 ) , .A2( u1_u15_u4_n118 ) , .A1( u1_u15_u4_n148 ) );
  NAND2_X1 u1_u15_u4_U24 (.ZN( u1_u15_u4_n129 ) , .A1( u1_u15_u4_n134 ) , .A2( u1_u15_u4_n148 ) );
  AND3_X1 u1_u15_u4_U25 (.A1( u1_u15_u4_n119 ) , .A2( u1_u15_u4_n143 ) , .A3( u1_u15_u4_n154 ) , .ZN( u1_u15_u4_n161 ) );
  AND2_X1 u1_u15_u4_U26 (.A1( u1_u15_u4_n145 ) , .A2( u1_u15_u4_n147 ) , .ZN( u1_u15_u4_n159 ) );
  OR3_X1 u1_u15_u4_U27 (.A3( u1_u15_u4_n114 ) , .A2( u1_u15_u4_n115 ) , .A1( u1_u15_u4_n116 ) , .ZN( u1_u15_u4_n136 ) );
  AOI21_X1 u1_u15_u4_U28 (.A( u1_u15_u4_n113 ) , .ZN( u1_u15_u4_n116 ) , .B2( u1_u15_u4_n173 ) , .B1( u1_u15_u4_n174 ) );
  AOI21_X1 u1_u15_u4_U29 (.ZN( u1_u15_u4_n115 ) , .B2( u1_u15_u4_n145 ) , .B1( u1_u15_u4_n146 ) , .A( u1_u15_u4_n156 ) );
  NOR2_X1 u1_u15_u4_U3 (.ZN( u1_u15_u4_n121 ) , .A1( u1_u15_u4_n181 ) , .A2( u1_u15_u4_n182 ) );
  OAI22_X1 u1_u15_u4_U30 (.ZN( u1_u15_u4_n114 ) , .A2( u1_u15_u4_n121 ) , .B1( u1_u15_u4_n160 ) , .B2( u1_u15_u4_n170 ) , .A1( u1_u15_u4_n171 ) );
  INV_X1 u1_u15_u4_U31 (.A( u1_u15_u4_n158 ) , .ZN( u1_u15_u4_n182 ) );
  INV_X1 u1_u15_u4_U32 (.ZN( u1_u15_u4_n181 ) , .A( u1_u15_u4_n96 ) );
  INV_X1 u1_u15_u4_U33 (.A( u1_u15_u4_n144 ) , .ZN( u1_u15_u4_n179 ) );
  INV_X1 u1_u15_u4_U34 (.A( u1_u15_u4_n157 ) , .ZN( u1_u15_u4_n178 ) );
  NAND2_X1 u1_u15_u4_U35 (.A2( u1_u15_u4_n154 ) , .A1( u1_u15_u4_n96 ) , .ZN( u1_u15_u4_n97 ) );
  INV_X1 u1_u15_u4_U36 (.ZN( u1_u15_u4_n186 ) , .A( u1_u15_u4_n95 ) );
  OAI221_X1 u1_u15_u4_U37 (.C1( u1_u15_u4_n134 ) , .B1( u1_u15_u4_n158 ) , .B2( u1_u15_u4_n171 ) , .C2( u1_u15_u4_n173 ) , .A( u1_u15_u4_n94 ) , .ZN( u1_u15_u4_n95 ) );
  AOI222_X1 u1_u15_u4_U38 (.B2( u1_u15_u4_n132 ) , .A1( u1_u15_u4_n138 ) , .C2( u1_u15_u4_n175 ) , .A2( u1_u15_u4_n179 ) , .C1( u1_u15_u4_n181 ) , .B1( u1_u15_u4_n185 ) , .ZN( u1_u15_u4_n94 ) );
  INV_X1 u1_u15_u4_U39 (.A( u1_u15_u4_n113 ) , .ZN( u1_u15_u4_n185 ) );
  INV_X1 u1_u15_u4_U4 (.A( u1_u15_u4_n117 ) , .ZN( u1_u15_u4_n184 ) );
  INV_X1 u1_u15_u4_U40 (.A( u1_u15_u4_n143 ) , .ZN( u1_u15_u4_n183 ) );
  NOR2_X1 u1_u15_u4_U41 (.ZN( u1_u15_u4_n138 ) , .A1( u1_u15_u4_n168 ) , .A2( u1_u15_u4_n169 ) );
  NOR2_X1 u1_u15_u4_U42 (.A1( u1_u15_u4_n150 ) , .A2( u1_u15_u4_n152 ) , .ZN( u1_u15_u4_n153 ) );
  NOR2_X1 u1_u15_u4_U43 (.A2( u1_u15_u4_n128 ) , .A1( u1_u15_u4_n138 ) , .ZN( u1_u15_u4_n156 ) );
  AOI22_X1 u1_u15_u4_U44 (.B2( u1_u15_u4_n122 ) , .A1( u1_u15_u4_n123 ) , .ZN( u1_u15_u4_n124 ) , .B1( u1_u15_u4_n128 ) , .A2( u1_u15_u4_n172 ) );
  NAND2_X1 u1_u15_u4_U45 (.A2( u1_u15_u4_n120 ) , .ZN( u1_u15_u4_n123 ) , .A1( u1_u15_u4_n161 ) );
  INV_X1 u1_u15_u4_U46 (.A( u1_u15_u4_n153 ) , .ZN( u1_u15_u4_n172 ) );
  AOI22_X1 u1_u15_u4_U47 (.B2( u1_u15_u4_n132 ) , .A2( u1_u15_u4_n133 ) , .ZN( u1_u15_u4_n140 ) , .A1( u1_u15_u4_n150 ) , .B1( u1_u15_u4_n179 ) );
  NAND2_X1 u1_u15_u4_U48 (.ZN( u1_u15_u4_n133 ) , .A2( u1_u15_u4_n146 ) , .A1( u1_u15_u4_n154 ) );
  NAND2_X1 u1_u15_u4_U49 (.A1( u1_u15_u4_n103 ) , .ZN( u1_u15_u4_n154 ) , .A2( u1_u15_u4_n98 ) );
  NOR4_X1 u1_u15_u4_U5 (.A4( u1_u15_u4_n106 ) , .A3( u1_u15_u4_n107 ) , .A2( u1_u15_u4_n108 ) , .A1( u1_u15_u4_n109 ) , .ZN( u1_u15_u4_n110 ) );
  NAND2_X1 u1_u15_u4_U50 (.A1( u1_u15_u4_n101 ) , .ZN( u1_u15_u4_n158 ) , .A2( u1_u15_u4_n99 ) );
  AOI21_X1 u1_u15_u4_U51 (.ZN( u1_u15_u4_n127 ) , .A( u1_u15_u4_n136 ) , .B2( u1_u15_u4_n150 ) , .B1( u1_u15_u4_n180 ) );
  INV_X1 u1_u15_u4_U52 (.A( u1_u15_u4_n160 ) , .ZN( u1_u15_u4_n180 ) );
  NAND2_X1 u1_u15_u4_U53 (.A2( u1_u15_u4_n104 ) , .A1( u1_u15_u4_n105 ) , .ZN( u1_u15_u4_n146 ) );
  NAND2_X1 u1_u15_u4_U54 (.A2( u1_u15_u4_n101 ) , .A1( u1_u15_u4_n102 ) , .ZN( u1_u15_u4_n160 ) );
  NAND2_X1 u1_u15_u4_U55 (.ZN( u1_u15_u4_n134 ) , .A1( u1_u15_u4_n98 ) , .A2( u1_u15_u4_n99 ) );
  NAND2_X1 u1_u15_u4_U56 (.A1( u1_u15_u4_n103 ) , .A2( u1_u15_u4_n104 ) , .ZN( u1_u15_u4_n143 ) );
  NAND2_X1 u1_u15_u4_U57 (.A2( u1_u15_u4_n105 ) , .ZN( u1_u15_u4_n145 ) , .A1( u1_u15_u4_n98 ) );
  NAND2_X1 u1_u15_u4_U58 (.A1( u1_u15_u4_n100 ) , .A2( u1_u15_u4_n105 ) , .ZN( u1_u15_u4_n120 ) );
  NAND2_X1 u1_u15_u4_U59 (.A1( u1_u15_u4_n102 ) , .A2( u1_u15_u4_n104 ) , .ZN( u1_u15_u4_n148 ) );
  AOI21_X1 u1_u15_u4_U6 (.ZN( u1_u15_u4_n106 ) , .B2( u1_u15_u4_n146 ) , .B1( u1_u15_u4_n158 ) , .A( u1_u15_u4_n170 ) );
  NAND2_X1 u1_u15_u4_U60 (.A2( u1_u15_u4_n100 ) , .A1( u1_u15_u4_n103 ) , .ZN( u1_u15_u4_n157 ) );
  INV_X1 u1_u15_u4_U61 (.A( u1_u15_u4_n150 ) , .ZN( u1_u15_u4_n173 ) );
  INV_X1 u1_u15_u4_U62 (.A( u1_u15_u4_n152 ) , .ZN( u1_u15_u4_n171 ) );
  NAND2_X1 u1_u15_u4_U63 (.A1( u1_u15_u4_n100 ) , .ZN( u1_u15_u4_n118 ) , .A2( u1_u15_u4_n99 ) );
  NAND2_X1 u1_u15_u4_U64 (.A2( u1_u15_u4_n100 ) , .A1( u1_u15_u4_n102 ) , .ZN( u1_u15_u4_n144 ) );
  NAND2_X1 u1_u15_u4_U65 (.A2( u1_u15_u4_n101 ) , .A1( u1_u15_u4_n105 ) , .ZN( u1_u15_u4_n96 ) );
  INV_X1 u1_u15_u4_U66 (.A( u1_u15_u4_n128 ) , .ZN( u1_u15_u4_n174 ) );
  NAND2_X1 u1_u15_u4_U67 (.A2( u1_u15_u4_n102 ) , .ZN( u1_u15_u4_n119 ) , .A1( u1_u15_u4_n98 ) );
  NAND2_X1 u1_u15_u4_U68 (.A2( u1_u15_u4_n101 ) , .A1( u1_u15_u4_n103 ) , .ZN( u1_u15_u4_n147 ) );
  NAND2_X1 u1_u15_u4_U69 (.A2( u1_u15_u4_n104 ) , .ZN( u1_u15_u4_n113 ) , .A1( u1_u15_u4_n99 ) );
  AOI21_X1 u1_u15_u4_U7 (.ZN( u1_u15_u4_n108 ) , .B2( u1_u15_u4_n134 ) , .B1( u1_u15_u4_n155 ) , .A( u1_u15_u4_n156 ) );
  NOR2_X1 u1_u15_u4_U70 (.A2( u1_u15_X_28 ) , .ZN( u1_u15_u4_n150 ) , .A1( u1_u15_u4_n168 ) );
  NOR2_X1 u1_u15_u4_U71 (.A2( u1_u15_X_29 ) , .ZN( u1_u15_u4_n152 ) , .A1( u1_u15_u4_n169 ) );
  NOR2_X1 u1_u15_u4_U72 (.A2( u1_u15_X_26 ) , .ZN( u1_u15_u4_n100 ) , .A1( u1_u15_u4_n177 ) );
  NOR2_X1 u1_u15_u4_U73 (.A2( u1_u15_X_30 ) , .ZN( u1_u15_u4_n105 ) , .A1( u1_u15_u4_n176 ) );
  NOR2_X1 u1_u15_u4_U74 (.A2( u1_u15_X_28 ) , .A1( u1_u15_X_29 ) , .ZN( u1_u15_u4_n128 ) );
  NOR2_X1 u1_u15_u4_U75 (.A2( u1_u15_X_25 ) , .A1( u1_u15_X_26 ) , .ZN( u1_u15_u4_n98 ) );
  NOR2_X1 u1_u15_u4_U76 (.A2( u1_u15_X_27 ) , .A1( u1_u15_X_30 ) , .ZN( u1_u15_u4_n102 ) );
  AND2_X1 u1_u15_u4_U77 (.A2( u1_u15_X_25 ) , .A1( u1_u15_X_26 ) , .ZN( u1_u15_u4_n104 ) );
  AND2_X1 u1_u15_u4_U78 (.A1( u1_u15_X_30 ) , .A2( u1_u15_u4_n176 ) , .ZN( u1_u15_u4_n99 ) );
  AND2_X1 u1_u15_u4_U79 (.A1( u1_u15_X_26 ) , .ZN( u1_u15_u4_n101 ) , .A2( u1_u15_u4_n177 ) );
  AOI21_X1 u1_u15_u4_U8 (.ZN( u1_u15_u4_n109 ) , .A( u1_u15_u4_n153 ) , .B1( u1_u15_u4_n159 ) , .B2( u1_u15_u4_n184 ) );
  AND2_X1 u1_u15_u4_U80 (.A1( u1_u15_X_27 ) , .A2( u1_u15_X_30 ) , .ZN( u1_u15_u4_n103 ) );
  INV_X1 u1_u15_u4_U81 (.A( u1_u15_X_28 ) , .ZN( u1_u15_u4_n169 ) );
  INV_X1 u1_u15_u4_U82 (.A( u1_u15_X_29 ) , .ZN( u1_u15_u4_n168 ) );
  INV_X1 u1_u15_u4_U83 (.A( u1_u15_X_25 ) , .ZN( u1_u15_u4_n177 ) );
  INV_X1 u1_u15_u4_U84 (.A( u1_u15_X_27 ) , .ZN( u1_u15_u4_n176 ) );
  NAND4_X1 u1_u15_u4_U85 (.ZN( u1_out15_25 ) , .A4( u1_u15_u4_n139 ) , .A3( u1_u15_u4_n140 ) , .A2( u1_u15_u4_n141 ) , .A1( u1_u15_u4_n142 ) );
  OAI21_X1 u1_u15_u4_U86 (.A( u1_u15_u4_n128 ) , .B2( u1_u15_u4_n129 ) , .B1( u1_u15_u4_n130 ) , .ZN( u1_u15_u4_n142 ) );
  OAI21_X1 u1_u15_u4_U87 (.B2( u1_u15_u4_n131 ) , .ZN( u1_u15_u4_n141 ) , .A( u1_u15_u4_n175 ) , .B1( u1_u15_u4_n183 ) );
  NAND4_X1 u1_u15_u4_U88 (.ZN( u1_out15_14 ) , .A4( u1_u15_u4_n124 ) , .A3( u1_u15_u4_n125 ) , .A2( u1_u15_u4_n126 ) , .A1( u1_u15_u4_n127 ) );
  AOI22_X1 u1_u15_u4_U89 (.B2( u1_u15_u4_n117 ) , .ZN( u1_u15_u4_n126 ) , .A1( u1_u15_u4_n129 ) , .B1( u1_u15_u4_n152 ) , .A2( u1_u15_u4_n175 ) );
  AOI211_X1 u1_u15_u4_U9 (.B( u1_u15_u4_n136 ) , .A( u1_u15_u4_n137 ) , .C2( u1_u15_u4_n138 ) , .ZN( u1_u15_u4_n139 ) , .C1( u1_u15_u4_n182 ) );
  AOI22_X1 u1_u15_u4_U90 (.ZN( u1_u15_u4_n125 ) , .B2( u1_u15_u4_n131 ) , .A2( u1_u15_u4_n132 ) , .B1( u1_u15_u4_n138 ) , .A1( u1_u15_u4_n178 ) );
  AOI22_X1 u1_u15_u4_U91 (.B2( u1_u15_u4_n149 ) , .B1( u1_u15_u4_n150 ) , .A2( u1_u15_u4_n151 ) , .A1( u1_u15_u4_n152 ) , .ZN( u1_u15_u4_n167 ) );
  NOR4_X1 u1_u15_u4_U92 (.A4( u1_u15_u4_n162 ) , .A3( u1_u15_u4_n163 ) , .A2( u1_u15_u4_n164 ) , .A1( u1_u15_u4_n165 ) , .ZN( u1_u15_u4_n166 ) );
  NAND4_X1 u1_u15_u4_U93 (.ZN( u1_out15_8 ) , .A4( u1_u15_u4_n110 ) , .A3( u1_u15_u4_n111 ) , .A2( u1_u15_u4_n112 ) , .A1( u1_u15_u4_n186 ) );
  NAND2_X1 u1_u15_u4_U94 (.ZN( u1_u15_u4_n112 ) , .A2( u1_u15_u4_n130 ) , .A1( u1_u15_u4_n150 ) );
  AOI22_X1 u1_u15_u4_U95 (.ZN( u1_u15_u4_n111 ) , .B2( u1_u15_u4_n132 ) , .A1( u1_u15_u4_n152 ) , .B1( u1_u15_u4_n178 ) , .A2( u1_u15_u4_n97 ) );
  NAND3_X1 u1_u15_u4_U96 (.ZN( u1_out15_3 ) , .A3( u1_u15_u4_n166 ) , .A1( u1_u15_u4_n167 ) , .A2( u1_u15_u4_n186 ) );
  NAND3_X1 u1_u15_u4_U97 (.A3( u1_u15_u4_n146 ) , .A2( u1_u15_u4_n147 ) , .A1( u1_u15_u4_n148 ) , .ZN( u1_u15_u4_n149 ) );
  NAND3_X1 u1_u15_u4_U98 (.A3( u1_u15_u4_n143 ) , .A2( u1_u15_u4_n144 ) , .A1( u1_u15_u4_n145 ) , .ZN( u1_u15_u4_n151 ) );
  NAND3_X1 u1_u15_u4_U99 (.A3( u1_u15_u4_n121 ) , .ZN( u1_u15_u4_n122 ) , .A2( u1_u15_u4_n144 ) , .A1( u1_u15_u4_n154 ) );
  INV_X1 u1_u15_u5_U10 (.A( u1_u15_u5_n121 ) , .ZN( u1_u15_u5_n177 ) );
  AOI222_X1 u1_u15_u5_U100 (.ZN( u1_u15_u5_n113 ) , .A1( u1_u15_u5_n131 ) , .C1( u1_u15_u5_n148 ) , .B2( u1_u15_u5_n174 ) , .C2( u1_u15_u5_n178 ) , .A2( u1_u15_u5_n179 ) , .B1( u1_u15_u5_n99 ) );
  NAND4_X1 u1_u15_u5_U101 (.ZN( u1_out15_29 ) , .A4( u1_u15_u5_n129 ) , .A3( u1_u15_u5_n130 ) , .A2( u1_u15_u5_n168 ) , .A1( u1_u15_u5_n196 ) );
  AOI221_X1 u1_u15_u5_U102 (.A( u1_u15_u5_n128 ) , .ZN( u1_u15_u5_n129 ) , .C2( u1_u15_u5_n132 ) , .B2( u1_u15_u5_n159 ) , .B1( u1_u15_u5_n176 ) , .C1( u1_u15_u5_n184 ) );
  AOI222_X1 u1_u15_u5_U103 (.ZN( u1_u15_u5_n130 ) , .A2( u1_u15_u5_n146 ) , .B1( u1_u15_u5_n147 ) , .C2( u1_u15_u5_n175 ) , .B2( u1_u15_u5_n179 ) , .A1( u1_u15_u5_n188 ) , .C1( u1_u15_u5_n194 ) );
  NAND3_X1 u1_u15_u5_U104 (.A2( u1_u15_u5_n154 ) , .A3( u1_u15_u5_n158 ) , .A1( u1_u15_u5_n161 ) , .ZN( u1_u15_u5_n99 ) );
  NOR2_X1 u1_u15_u5_U11 (.ZN( u1_u15_u5_n160 ) , .A2( u1_u15_u5_n173 ) , .A1( u1_u15_u5_n177 ) );
  INV_X1 u1_u15_u5_U12 (.A( u1_u15_u5_n150 ) , .ZN( u1_u15_u5_n174 ) );
  AOI21_X1 u1_u15_u5_U13 (.A( u1_u15_u5_n160 ) , .B2( u1_u15_u5_n161 ) , .ZN( u1_u15_u5_n162 ) , .B1( u1_u15_u5_n192 ) );
  INV_X1 u1_u15_u5_U14 (.A( u1_u15_u5_n159 ) , .ZN( u1_u15_u5_n192 ) );
  AOI21_X1 u1_u15_u5_U15 (.A( u1_u15_u5_n156 ) , .B2( u1_u15_u5_n157 ) , .B1( u1_u15_u5_n158 ) , .ZN( u1_u15_u5_n163 ) );
  AOI21_X1 u1_u15_u5_U16 (.B2( u1_u15_u5_n139 ) , .B1( u1_u15_u5_n140 ) , .ZN( u1_u15_u5_n141 ) , .A( u1_u15_u5_n150 ) );
  OAI21_X1 u1_u15_u5_U17 (.A( u1_u15_u5_n133 ) , .B2( u1_u15_u5_n134 ) , .B1( u1_u15_u5_n135 ) , .ZN( u1_u15_u5_n142 ) );
  OAI21_X1 u1_u15_u5_U18 (.ZN( u1_u15_u5_n133 ) , .B2( u1_u15_u5_n147 ) , .A( u1_u15_u5_n173 ) , .B1( u1_u15_u5_n188 ) );
  NAND2_X1 u1_u15_u5_U19 (.A2( u1_u15_u5_n119 ) , .A1( u1_u15_u5_n123 ) , .ZN( u1_u15_u5_n137 ) );
  INV_X1 u1_u15_u5_U20 (.A( u1_u15_u5_n155 ) , .ZN( u1_u15_u5_n194 ) );
  NAND2_X1 u1_u15_u5_U21 (.A1( u1_u15_u5_n121 ) , .ZN( u1_u15_u5_n132 ) , .A2( u1_u15_u5_n172 ) );
  NAND2_X1 u1_u15_u5_U22 (.A2( u1_u15_u5_n122 ) , .ZN( u1_u15_u5_n136 ) , .A1( u1_u15_u5_n154 ) );
  NAND2_X1 u1_u15_u5_U23 (.A2( u1_u15_u5_n119 ) , .A1( u1_u15_u5_n120 ) , .ZN( u1_u15_u5_n159 ) );
  INV_X1 u1_u15_u5_U24 (.A( u1_u15_u5_n156 ) , .ZN( u1_u15_u5_n175 ) );
  INV_X1 u1_u15_u5_U25 (.A( u1_u15_u5_n158 ) , .ZN( u1_u15_u5_n188 ) );
  INV_X1 u1_u15_u5_U26 (.A( u1_u15_u5_n152 ) , .ZN( u1_u15_u5_n179 ) );
  INV_X1 u1_u15_u5_U27 (.A( u1_u15_u5_n140 ) , .ZN( u1_u15_u5_n182 ) );
  INV_X1 u1_u15_u5_U28 (.A( u1_u15_u5_n151 ) , .ZN( u1_u15_u5_n183 ) );
  INV_X1 u1_u15_u5_U29 (.A( u1_u15_u5_n123 ) , .ZN( u1_u15_u5_n185 ) );
  NOR2_X1 u1_u15_u5_U3 (.ZN( u1_u15_u5_n134 ) , .A1( u1_u15_u5_n183 ) , .A2( u1_u15_u5_n190 ) );
  INV_X1 u1_u15_u5_U30 (.A( u1_u15_u5_n161 ) , .ZN( u1_u15_u5_n184 ) );
  INV_X1 u1_u15_u5_U31 (.A( u1_u15_u5_n139 ) , .ZN( u1_u15_u5_n189 ) );
  INV_X1 u1_u15_u5_U32 (.A( u1_u15_u5_n157 ) , .ZN( u1_u15_u5_n190 ) );
  INV_X1 u1_u15_u5_U33 (.A( u1_u15_u5_n120 ) , .ZN( u1_u15_u5_n193 ) );
  NAND2_X1 u1_u15_u5_U34 (.ZN( u1_u15_u5_n111 ) , .A1( u1_u15_u5_n140 ) , .A2( u1_u15_u5_n155 ) );
  NOR2_X1 u1_u15_u5_U35 (.ZN( u1_u15_u5_n100 ) , .A1( u1_u15_u5_n170 ) , .A2( u1_u15_u5_n180 ) );
  INV_X1 u1_u15_u5_U36 (.A( u1_u15_u5_n117 ) , .ZN( u1_u15_u5_n196 ) );
  OAI221_X1 u1_u15_u5_U37 (.A( u1_u15_u5_n116 ) , .ZN( u1_u15_u5_n117 ) , .B2( u1_u15_u5_n119 ) , .C1( u1_u15_u5_n153 ) , .C2( u1_u15_u5_n158 ) , .B1( u1_u15_u5_n172 ) );
  AOI222_X1 u1_u15_u5_U38 (.ZN( u1_u15_u5_n116 ) , .B2( u1_u15_u5_n145 ) , .C1( u1_u15_u5_n148 ) , .A2( u1_u15_u5_n174 ) , .C2( u1_u15_u5_n177 ) , .B1( u1_u15_u5_n187 ) , .A1( u1_u15_u5_n193 ) );
  INV_X1 u1_u15_u5_U39 (.A( u1_u15_u5_n115 ) , .ZN( u1_u15_u5_n187 ) );
  INV_X1 u1_u15_u5_U4 (.A( u1_u15_u5_n138 ) , .ZN( u1_u15_u5_n191 ) );
  AOI22_X1 u1_u15_u5_U40 (.B2( u1_u15_u5_n131 ) , .A2( u1_u15_u5_n146 ) , .ZN( u1_u15_u5_n169 ) , .B1( u1_u15_u5_n174 ) , .A1( u1_u15_u5_n185 ) );
  NOR2_X1 u1_u15_u5_U41 (.A1( u1_u15_u5_n146 ) , .ZN( u1_u15_u5_n150 ) , .A2( u1_u15_u5_n173 ) );
  AOI21_X1 u1_u15_u5_U42 (.A( u1_u15_u5_n118 ) , .B2( u1_u15_u5_n145 ) , .ZN( u1_u15_u5_n168 ) , .B1( u1_u15_u5_n186 ) );
  INV_X1 u1_u15_u5_U43 (.A( u1_u15_u5_n122 ) , .ZN( u1_u15_u5_n186 ) );
  NOR2_X1 u1_u15_u5_U44 (.A1( u1_u15_u5_n146 ) , .ZN( u1_u15_u5_n152 ) , .A2( u1_u15_u5_n176 ) );
  NOR2_X1 u1_u15_u5_U45 (.A1( u1_u15_u5_n115 ) , .ZN( u1_u15_u5_n118 ) , .A2( u1_u15_u5_n153 ) );
  NOR2_X1 u1_u15_u5_U46 (.A2( u1_u15_u5_n145 ) , .ZN( u1_u15_u5_n156 ) , .A1( u1_u15_u5_n174 ) );
  NOR2_X1 u1_u15_u5_U47 (.ZN( u1_u15_u5_n121 ) , .A2( u1_u15_u5_n145 ) , .A1( u1_u15_u5_n176 ) );
  AOI22_X1 u1_u15_u5_U48 (.ZN( u1_u15_u5_n114 ) , .A2( u1_u15_u5_n137 ) , .A1( u1_u15_u5_n145 ) , .B2( u1_u15_u5_n175 ) , .B1( u1_u15_u5_n193 ) );
  OAI211_X1 u1_u15_u5_U49 (.B( u1_u15_u5_n124 ) , .A( u1_u15_u5_n125 ) , .C2( u1_u15_u5_n126 ) , .C1( u1_u15_u5_n127 ) , .ZN( u1_u15_u5_n128 ) );
  OAI21_X1 u1_u15_u5_U5 (.B2( u1_u15_u5_n136 ) , .B1( u1_u15_u5_n137 ) , .ZN( u1_u15_u5_n138 ) , .A( u1_u15_u5_n177 ) );
  NOR3_X1 u1_u15_u5_U50 (.ZN( u1_u15_u5_n127 ) , .A1( u1_u15_u5_n136 ) , .A3( u1_u15_u5_n148 ) , .A2( u1_u15_u5_n182 ) );
  OAI21_X1 u1_u15_u5_U51 (.ZN( u1_u15_u5_n124 ) , .A( u1_u15_u5_n177 ) , .B2( u1_u15_u5_n183 ) , .B1( u1_u15_u5_n189 ) );
  OAI21_X1 u1_u15_u5_U52 (.ZN( u1_u15_u5_n125 ) , .A( u1_u15_u5_n174 ) , .B2( u1_u15_u5_n185 ) , .B1( u1_u15_u5_n190 ) );
  AOI21_X1 u1_u15_u5_U53 (.A( u1_u15_u5_n153 ) , .B2( u1_u15_u5_n154 ) , .B1( u1_u15_u5_n155 ) , .ZN( u1_u15_u5_n164 ) );
  AOI21_X1 u1_u15_u5_U54 (.ZN( u1_u15_u5_n110 ) , .B1( u1_u15_u5_n122 ) , .B2( u1_u15_u5_n139 ) , .A( u1_u15_u5_n153 ) );
  INV_X1 u1_u15_u5_U55 (.A( u1_u15_u5_n153 ) , .ZN( u1_u15_u5_n176 ) );
  INV_X1 u1_u15_u5_U56 (.A( u1_u15_u5_n126 ) , .ZN( u1_u15_u5_n173 ) );
  AND2_X1 u1_u15_u5_U57 (.A2( u1_u15_u5_n104 ) , .A1( u1_u15_u5_n107 ) , .ZN( u1_u15_u5_n147 ) );
  AND2_X1 u1_u15_u5_U58 (.A2( u1_u15_u5_n104 ) , .A1( u1_u15_u5_n108 ) , .ZN( u1_u15_u5_n148 ) );
  NAND2_X1 u1_u15_u5_U59 (.A1( u1_u15_u5_n105 ) , .A2( u1_u15_u5_n106 ) , .ZN( u1_u15_u5_n158 ) );
  INV_X1 u1_u15_u5_U6 (.A( u1_u15_u5_n135 ) , .ZN( u1_u15_u5_n178 ) );
  NAND2_X1 u1_u15_u5_U60 (.A2( u1_u15_u5_n108 ) , .A1( u1_u15_u5_n109 ) , .ZN( u1_u15_u5_n139 ) );
  NAND2_X1 u1_u15_u5_U61 (.A1( u1_u15_u5_n106 ) , .A2( u1_u15_u5_n108 ) , .ZN( u1_u15_u5_n119 ) );
  NAND2_X1 u1_u15_u5_U62 (.A2( u1_u15_u5_n103 ) , .A1( u1_u15_u5_n105 ) , .ZN( u1_u15_u5_n140 ) );
  NAND2_X1 u1_u15_u5_U63 (.A2( u1_u15_u5_n104 ) , .A1( u1_u15_u5_n105 ) , .ZN( u1_u15_u5_n155 ) );
  NAND2_X1 u1_u15_u5_U64 (.A2( u1_u15_u5_n106 ) , .A1( u1_u15_u5_n107 ) , .ZN( u1_u15_u5_n122 ) );
  NAND2_X1 u1_u15_u5_U65 (.A2( u1_u15_u5_n100 ) , .A1( u1_u15_u5_n106 ) , .ZN( u1_u15_u5_n115 ) );
  NAND2_X1 u1_u15_u5_U66 (.A2( u1_u15_u5_n100 ) , .A1( u1_u15_u5_n103 ) , .ZN( u1_u15_u5_n161 ) );
  NAND2_X1 u1_u15_u5_U67 (.A1( u1_u15_u5_n105 ) , .A2( u1_u15_u5_n109 ) , .ZN( u1_u15_u5_n154 ) );
  INV_X1 u1_u15_u5_U68 (.A( u1_u15_u5_n146 ) , .ZN( u1_u15_u5_n172 ) );
  NAND2_X1 u1_u15_u5_U69 (.A1( u1_u15_u5_n103 ) , .A2( u1_u15_u5_n108 ) , .ZN( u1_u15_u5_n123 ) );
  OAI22_X1 u1_u15_u5_U7 (.B2( u1_u15_u5_n149 ) , .B1( u1_u15_u5_n150 ) , .A2( u1_u15_u5_n151 ) , .A1( u1_u15_u5_n152 ) , .ZN( u1_u15_u5_n165 ) );
  NAND2_X1 u1_u15_u5_U70 (.A2( u1_u15_u5_n103 ) , .A1( u1_u15_u5_n107 ) , .ZN( u1_u15_u5_n151 ) );
  NAND2_X1 u1_u15_u5_U71 (.A2( u1_u15_u5_n107 ) , .A1( u1_u15_u5_n109 ) , .ZN( u1_u15_u5_n120 ) );
  NAND2_X1 u1_u15_u5_U72 (.A2( u1_u15_u5_n100 ) , .A1( u1_u15_u5_n109 ) , .ZN( u1_u15_u5_n157 ) );
  AND2_X1 u1_u15_u5_U73 (.A2( u1_u15_u5_n100 ) , .A1( u1_u15_u5_n104 ) , .ZN( u1_u15_u5_n131 ) );
  INV_X1 u1_u15_u5_U74 (.A( u1_u15_u5_n102 ) , .ZN( u1_u15_u5_n195 ) );
  OAI221_X1 u1_u15_u5_U75 (.A( u1_u15_u5_n101 ) , .ZN( u1_u15_u5_n102 ) , .C2( u1_u15_u5_n115 ) , .C1( u1_u15_u5_n126 ) , .B1( u1_u15_u5_n134 ) , .B2( u1_u15_u5_n160 ) );
  OAI21_X1 u1_u15_u5_U76 (.ZN( u1_u15_u5_n101 ) , .B1( u1_u15_u5_n137 ) , .A( u1_u15_u5_n146 ) , .B2( u1_u15_u5_n147 ) );
  NOR2_X1 u1_u15_u5_U77 (.A2( u1_u15_X_34 ) , .A1( u1_u15_X_35 ) , .ZN( u1_u15_u5_n145 ) );
  NOR2_X1 u1_u15_u5_U78 (.A2( u1_u15_X_34 ) , .ZN( u1_u15_u5_n146 ) , .A1( u1_u15_u5_n171 ) );
  NOR2_X1 u1_u15_u5_U79 (.A2( u1_u15_X_31 ) , .A1( u1_u15_X_32 ) , .ZN( u1_u15_u5_n103 ) );
  NOR3_X1 u1_u15_u5_U8 (.A2( u1_u15_u5_n147 ) , .A1( u1_u15_u5_n148 ) , .ZN( u1_u15_u5_n149 ) , .A3( u1_u15_u5_n194 ) );
  NOR2_X1 u1_u15_u5_U80 (.A2( u1_u15_X_36 ) , .ZN( u1_u15_u5_n105 ) , .A1( u1_u15_u5_n180 ) );
  NOR2_X1 u1_u15_u5_U81 (.A2( u1_u15_X_33 ) , .ZN( u1_u15_u5_n108 ) , .A1( u1_u15_u5_n170 ) );
  NOR2_X1 u1_u15_u5_U82 (.A2( u1_u15_X_33 ) , .A1( u1_u15_X_36 ) , .ZN( u1_u15_u5_n107 ) );
  NOR2_X1 u1_u15_u5_U83 (.A2( u1_u15_X_31 ) , .ZN( u1_u15_u5_n104 ) , .A1( u1_u15_u5_n181 ) );
  NAND2_X1 u1_u15_u5_U84 (.A2( u1_u15_X_34 ) , .A1( u1_u15_X_35 ) , .ZN( u1_u15_u5_n153 ) );
  NAND2_X1 u1_u15_u5_U85 (.A1( u1_u15_X_34 ) , .ZN( u1_u15_u5_n126 ) , .A2( u1_u15_u5_n171 ) );
  AND2_X1 u1_u15_u5_U86 (.A1( u1_u15_X_31 ) , .A2( u1_u15_X_32 ) , .ZN( u1_u15_u5_n106 ) );
  AND2_X1 u1_u15_u5_U87 (.A1( u1_u15_X_31 ) , .ZN( u1_u15_u5_n109 ) , .A2( u1_u15_u5_n181 ) );
  INV_X1 u1_u15_u5_U88 (.A( u1_u15_X_33 ) , .ZN( u1_u15_u5_n180 ) );
  INV_X1 u1_u15_u5_U89 (.A( u1_u15_X_35 ) , .ZN( u1_u15_u5_n171 ) );
  NOR2_X1 u1_u15_u5_U9 (.ZN( u1_u15_u5_n135 ) , .A1( u1_u15_u5_n173 ) , .A2( u1_u15_u5_n176 ) );
  INV_X1 u1_u15_u5_U90 (.A( u1_u15_X_36 ) , .ZN( u1_u15_u5_n170 ) );
  INV_X1 u1_u15_u5_U91 (.A( u1_u15_X_32 ) , .ZN( u1_u15_u5_n181 ) );
  NAND4_X1 u1_u15_u5_U92 (.ZN( u1_out15_19 ) , .A4( u1_u15_u5_n166 ) , .A3( u1_u15_u5_n167 ) , .A2( u1_u15_u5_n168 ) , .A1( u1_u15_u5_n169 ) );
  AOI22_X1 u1_u15_u5_U93 (.B2( u1_u15_u5_n145 ) , .A2( u1_u15_u5_n146 ) , .ZN( u1_u15_u5_n167 ) , .B1( u1_u15_u5_n182 ) , .A1( u1_u15_u5_n189 ) );
  NOR4_X1 u1_u15_u5_U94 (.A4( u1_u15_u5_n162 ) , .A3( u1_u15_u5_n163 ) , .A2( u1_u15_u5_n164 ) , .A1( u1_u15_u5_n165 ) , .ZN( u1_u15_u5_n166 ) );
  NAND4_X1 u1_u15_u5_U95 (.ZN( u1_out15_11 ) , .A4( u1_u15_u5_n143 ) , .A3( u1_u15_u5_n144 ) , .A2( u1_u15_u5_n169 ) , .A1( u1_u15_u5_n196 ) );
  AOI22_X1 u1_u15_u5_U96 (.A2( u1_u15_u5_n132 ) , .ZN( u1_u15_u5_n144 ) , .B2( u1_u15_u5_n145 ) , .B1( u1_u15_u5_n184 ) , .A1( u1_u15_u5_n194 ) );
  NOR3_X1 u1_u15_u5_U97 (.A3( u1_u15_u5_n141 ) , .A1( u1_u15_u5_n142 ) , .ZN( u1_u15_u5_n143 ) , .A2( u1_u15_u5_n191 ) );
  NAND4_X1 u1_u15_u5_U98 (.ZN( u1_out15_4 ) , .A4( u1_u15_u5_n112 ) , .A2( u1_u15_u5_n113 ) , .A1( u1_u15_u5_n114 ) , .A3( u1_u15_u5_n195 ) );
  AOI211_X1 u1_u15_u5_U99 (.A( u1_u15_u5_n110 ) , .C1( u1_u15_u5_n111 ) , .ZN( u1_u15_u5_n112 ) , .B( u1_u15_u5_n118 ) , .C2( u1_u15_u5_n177 ) );
  INV_X1 u1_u15_u6_U10 (.ZN( u1_u15_u6_n172 ) , .A( u1_u15_u6_n88 ) );
  OAI21_X1 u1_u15_u6_U11 (.A( u1_u15_u6_n159 ) , .B1( u1_u15_u6_n169 ) , .B2( u1_u15_u6_n173 ) , .ZN( u1_u15_u6_n90 ) );
  AOI22_X1 u1_u15_u6_U12 (.A2( u1_u15_u6_n151 ) , .B2( u1_u15_u6_n161 ) , .A1( u1_u15_u6_n167 ) , .B1( u1_u15_u6_n170 ) , .ZN( u1_u15_u6_n89 ) );
  AOI21_X1 u1_u15_u6_U13 (.ZN( u1_u15_u6_n106 ) , .A( u1_u15_u6_n142 ) , .B2( u1_u15_u6_n159 ) , .B1( u1_u15_u6_n164 ) );
  INV_X1 u1_u15_u6_U14 (.A( u1_u15_u6_n155 ) , .ZN( u1_u15_u6_n161 ) );
  INV_X1 u1_u15_u6_U15 (.A( u1_u15_u6_n128 ) , .ZN( u1_u15_u6_n164 ) );
  NAND2_X1 u1_u15_u6_U16 (.ZN( u1_u15_u6_n110 ) , .A1( u1_u15_u6_n122 ) , .A2( u1_u15_u6_n129 ) );
  NAND2_X1 u1_u15_u6_U17 (.ZN( u1_u15_u6_n124 ) , .A2( u1_u15_u6_n146 ) , .A1( u1_u15_u6_n148 ) );
  INV_X1 u1_u15_u6_U18 (.A( u1_u15_u6_n132 ) , .ZN( u1_u15_u6_n171 ) );
  AND2_X1 u1_u15_u6_U19 (.A1( u1_u15_u6_n100 ) , .ZN( u1_u15_u6_n130 ) , .A2( u1_u15_u6_n147 ) );
  INV_X1 u1_u15_u6_U20 (.A( u1_u15_u6_n127 ) , .ZN( u1_u15_u6_n173 ) );
  INV_X1 u1_u15_u6_U21 (.A( u1_u15_u6_n121 ) , .ZN( u1_u15_u6_n167 ) );
  INV_X1 u1_u15_u6_U22 (.A( u1_u15_u6_n100 ) , .ZN( u1_u15_u6_n169 ) );
  INV_X1 u1_u15_u6_U23 (.A( u1_u15_u6_n123 ) , .ZN( u1_u15_u6_n170 ) );
  INV_X1 u1_u15_u6_U24 (.A( u1_u15_u6_n113 ) , .ZN( u1_u15_u6_n168 ) );
  AND2_X1 u1_u15_u6_U25 (.A1( u1_u15_u6_n107 ) , .A2( u1_u15_u6_n119 ) , .ZN( u1_u15_u6_n133 ) );
  AND2_X1 u1_u15_u6_U26 (.A2( u1_u15_u6_n121 ) , .A1( u1_u15_u6_n122 ) , .ZN( u1_u15_u6_n131 ) );
  AND3_X1 u1_u15_u6_U27 (.ZN( u1_u15_u6_n120 ) , .A2( u1_u15_u6_n127 ) , .A1( u1_u15_u6_n132 ) , .A3( u1_u15_u6_n145 ) );
  INV_X1 u1_u15_u6_U28 (.A( u1_u15_u6_n146 ) , .ZN( u1_u15_u6_n163 ) );
  AOI222_X1 u1_u15_u6_U29 (.ZN( u1_u15_u6_n114 ) , .A1( u1_u15_u6_n118 ) , .A2( u1_u15_u6_n126 ) , .B2( u1_u15_u6_n151 ) , .C2( u1_u15_u6_n159 ) , .C1( u1_u15_u6_n168 ) , .B1( u1_u15_u6_n169 ) );
  INV_X1 u1_u15_u6_U3 (.A( u1_u15_u6_n110 ) , .ZN( u1_u15_u6_n166 ) );
  NOR2_X1 u1_u15_u6_U30 (.A1( u1_u15_u6_n162 ) , .A2( u1_u15_u6_n165 ) , .ZN( u1_u15_u6_n98 ) );
  NAND2_X1 u1_u15_u6_U31 (.A1( u1_u15_u6_n144 ) , .ZN( u1_u15_u6_n151 ) , .A2( u1_u15_u6_n158 ) );
  NAND2_X1 u1_u15_u6_U32 (.ZN( u1_u15_u6_n132 ) , .A1( u1_u15_u6_n91 ) , .A2( u1_u15_u6_n97 ) );
  AOI22_X1 u1_u15_u6_U33 (.B2( u1_u15_u6_n110 ) , .B1( u1_u15_u6_n111 ) , .A1( u1_u15_u6_n112 ) , .ZN( u1_u15_u6_n115 ) , .A2( u1_u15_u6_n161 ) );
  NAND4_X1 u1_u15_u6_U34 (.A3( u1_u15_u6_n109 ) , .ZN( u1_u15_u6_n112 ) , .A4( u1_u15_u6_n132 ) , .A2( u1_u15_u6_n147 ) , .A1( u1_u15_u6_n166 ) );
  NOR2_X1 u1_u15_u6_U35 (.ZN( u1_u15_u6_n109 ) , .A1( u1_u15_u6_n170 ) , .A2( u1_u15_u6_n173 ) );
  NOR2_X1 u1_u15_u6_U36 (.A2( u1_u15_u6_n126 ) , .ZN( u1_u15_u6_n155 ) , .A1( u1_u15_u6_n160 ) );
  NAND2_X1 u1_u15_u6_U37 (.ZN( u1_u15_u6_n146 ) , .A2( u1_u15_u6_n94 ) , .A1( u1_u15_u6_n99 ) );
  AOI21_X1 u1_u15_u6_U38 (.A( u1_u15_u6_n144 ) , .B2( u1_u15_u6_n145 ) , .B1( u1_u15_u6_n146 ) , .ZN( u1_u15_u6_n150 ) );
  AOI211_X1 u1_u15_u6_U39 (.B( u1_u15_u6_n134 ) , .A( u1_u15_u6_n135 ) , .C1( u1_u15_u6_n136 ) , .ZN( u1_u15_u6_n137 ) , .C2( u1_u15_u6_n151 ) );
  INV_X1 u1_u15_u6_U4 (.A( u1_u15_u6_n142 ) , .ZN( u1_u15_u6_n174 ) );
  NAND4_X1 u1_u15_u6_U40 (.A4( u1_u15_u6_n127 ) , .A3( u1_u15_u6_n128 ) , .A2( u1_u15_u6_n129 ) , .A1( u1_u15_u6_n130 ) , .ZN( u1_u15_u6_n136 ) );
  AOI21_X1 u1_u15_u6_U41 (.B2( u1_u15_u6_n132 ) , .B1( u1_u15_u6_n133 ) , .ZN( u1_u15_u6_n134 ) , .A( u1_u15_u6_n158 ) );
  AOI21_X1 u1_u15_u6_U42 (.B1( u1_u15_u6_n131 ) , .ZN( u1_u15_u6_n135 ) , .A( u1_u15_u6_n144 ) , .B2( u1_u15_u6_n146 ) );
  INV_X1 u1_u15_u6_U43 (.A( u1_u15_u6_n111 ) , .ZN( u1_u15_u6_n158 ) );
  NAND2_X1 u1_u15_u6_U44 (.ZN( u1_u15_u6_n127 ) , .A1( u1_u15_u6_n91 ) , .A2( u1_u15_u6_n92 ) );
  NAND2_X1 u1_u15_u6_U45 (.ZN( u1_u15_u6_n129 ) , .A2( u1_u15_u6_n95 ) , .A1( u1_u15_u6_n96 ) );
  INV_X1 u1_u15_u6_U46 (.A( u1_u15_u6_n144 ) , .ZN( u1_u15_u6_n159 ) );
  NAND2_X1 u1_u15_u6_U47 (.ZN( u1_u15_u6_n145 ) , .A2( u1_u15_u6_n97 ) , .A1( u1_u15_u6_n98 ) );
  NAND2_X1 u1_u15_u6_U48 (.ZN( u1_u15_u6_n148 ) , .A2( u1_u15_u6_n92 ) , .A1( u1_u15_u6_n94 ) );
  NAND2_X1 u1_u15_u6_U49 (.ZN( u1_u15_u6_n108 ) , .A2( u1_u15_u6_n139 ) , .A1( u1_u15_u6_n144 ) );
  NAND2_X1 u1_u15_u6_U5 (.A2( u1_u15_u6_n143 ) , .ZN( u1_u15_u6_n152 ) , .A1( u1_u15_u6_n166 ) );
  NAND2_X1 u1_u15_u6_U50 (.ZN( u1_u15_u6_n121 ) , .A2( u1_u15_u6_n95 ) , .A1( u1_u15_u6_n97 ) );
  NAND2_X1 u1_u15_u6_U51 (.ZN( u1_u15_u6_n107 ) , .A2( u1_u15_u6_n92 ) , .A1( u1_u15_u6_n95 ) );
  AND2_X1 u1_u15_u6_U52 (.ZN( u1_u15_u6_n118 ) , .A2( u1_u15_u6_n91 ) , .A1( u1_u15_u6_n99 ) );
  NAND2_X1 u1_u15_u6_U53 (.ZN( u1_u15_u6_n147 ) , .A2( u1_u15_u6_n98 ) , .A1( u1_u15_u6_n99 ) );
  NAND2_X1 u1_u15_u6_U54 (.ZN( u1_u15_u6_n128 ) , .A1( u1_u15_u6_n94 ) , .A2( u1_u15_u6_n96 ) );
  NAND2_X1 u1_u15_u6_U55 (.ZN( u1_u15_u6_n119 ) , .A2( u1_u15_u6_n95 ) , .A1( u1_u15_u6_n99 ) );
  NAND2_X1 u1_u15_u6_U56 (.ZN( u1_u15_u6_n123 ) , .A2( u1_u15_u6_n91 ) , .A1( u1_u15_u6_n96 ) );
  NAND2_X1 u1_u15_u6_U57 (.ZN( u1_u15_u6_n100 ) , .A2( u1_u15_u6_n92 ) , .A1( u1_u15_u6_n98 ) );
  NAND2_X1 u1_u15_u6_U58 (.ZN( u1_u15_u6_n122 ) , .A1( u1_u15_u6_n94 ) , .A2( u1_u15_u6_n97 ) );
  INV_X1 u1_u15_u6_U59 (.A( u1_u15_u6_n139 ) , .ZN( u1_u15_u6_n160 ) );
  AOI22_X1 u1_u15_u6_U6 (.B2( u1_u15_u6_n101 ) , .A1( u1_u15_u6_n102 ) , .ZN( u1_u15_u6_n103 ) , .B1( u1_u15_u6_n160 ) , .A2( u1_u15_u6_n161 ) );
  NAND2_X1 u1_u15_u6_U60 (.ZN( u1_u15_u6_n113 ) , .A1( u1_u15_u6_n96 ) , .A2( u1_u15_u6_n98 ) );
  NOR2_X1 u1_u15_u6_U61 (.A2( u1_u15_X_40 ) , .A1( u1_u15_X_41 ) , .ZN( u1_u15_u6_n126 ) );
  NOR2_X1 u1_u15_u6_U62 (.A2( u1_u15_X_39 ) , .A1( u1_u15_X_42 ) , .ZN( u1_u15_u6_n92 ) );
  NOR2_X1 u1_u15_u6_U63 (.A2( u1_u15_X_39 ) , .A1( u1_u15_u6_n156 ) , .ZN( u1_u15_u6_n97 ) );
  NOR2_X1 u1_u15_u6_U64 (.A2( u1_u15_X_38 ) , .A1( u1_u15_u6_n165 ) , .ZN( u1_u15_u6_n95 ) );
  NOR2_X1 u1_u15_u6_U65 (.A2( u1_u15_X_41 ) , .ZN( u1_u15_u6_n111 ) , .A1( u1_u15_u6_n157 ) );
  NOR2_X1 u1_u15_u6_U66 (.A2( u1_u15_X_37 ) , .A1( u1_u15_u6_n162 ) , .ZN( u1_u15_u6_n94 ) );
  NOR2_X1 u1_u15_u6_U67 (.A2( u1_u15_X_37 ) , .A1( u1_u15_X_38 ) , .ZN( u1_u15_u6_n91 ) );
  NAND2_X1 u1_u15_u6_U68 (.A1( u1_u15_X_41 ) , .ZN( u1_u15_u6_n144 ) , .A2( u1_u15_u6_n157 ) );
  NAND2_X1 u1_u15_u6_U69 (.A2( u1_u15_X_40 ) , .A1( u1_u15_X_41 ) , .ZN( u1_u15_u6_n139 ) );
  NOR2_X1 u1_u15_u6_U7 (.A1( u1_u15_u6_n118 ) , .ZN( u1_u15_u6_n143 ) , .A2( u1_u15_u6_n168 ) );
  AND2_X1 u1_u15_u6_U70 (.A1( u1_u15_X_39 ) , .A2( u1_u15_u6_n156 ) , .ZN( u1_u15_u6_n96 ) );
  AND2_X1 u1_u15_u6_U71 (.A1( u1_u15_X_39 ) , .A2( u1_u15_X_42 ) , .ZN( u1_u15_u6_n99 ) );
  INV_X1 u1_u15_u6_U72 (.A( u1_u15_X_40 ) , .ZN( u1_u15_u6_n157 ) );
  INV_X1 u1_u15_u6_U73 (.A( u1_u15_X_37 ) , .ZN( u1_u15_u6_n165 ) );
  INV_X1 u1_u15_u6_U74 (.A( u1_u15_X_38 ) , .ZN( u1_u15_u6_n162 ) );
  INV_X1 u1_u15_u6_U75 (.A( u1_u15_X_42 ) , .ZN( u1_u15_u6_n156 ) );
  NAND4_X1 u1_u15_u6_U76 (.ZN( u1_out15_12 ) , .A4( u1_u15_u6_n114 ) , .A3( u1_u15_u6_n115 ) , .A2( u1_u15_u6_n116 ) , .A1( u1_u15_u6_n117 ) );
  OAI22_X1 u1_u15_u6_U77 (.B2( u1_u15_u6_n111 ) , .ZN( u1_u15_u6_n116 ) , .B1( u1_u15_u6_n126 ) , .A2( u1_u15_u6_n164 ) , .A1( u1_u15_u6_n167 ) );
  OAI21_X1 u1_u15_u6_U78 (.A( u1_u15_u6_n108 ) , .ZN( u1_u15_u6_n117 ) , .B2( u1_u15_u6_n141 ) , .B1( u1_u15_u6_n163 ) );
  NAND4_X1 u1_u15_u6_U79 (.ZN( u1_out15_32 ) , .A4( u1_u15_u6_n103 ) , .A3( u1_u15_u6_n104 ) , .A2( u1_u15_u6_n105 ) , .A1( u1_u15_u6_n106 ) );
  AOI21_X1 u1_u15_u6_U8 (.B1( u1_u15_u6_n107 ) , .B2( u1_u15_u6_n132 ) , .A( u1_u15_u6_n158 ) , .ZN( u1_u15_u6_n88 ) );
  AOI22_X1 u1_u15_u6_U80 (.ZN( u1_u15_u6_n105 ) , .A2( u1_u15_u6_n108 ) , .A1( u1_u15_u6_n118 ) , .B2( u1_u15_u6_n126 ) , .B1( u1_u15_u6_n171 ) );
  AOI22_X1 u1_u15_u6_U81 (.ZN( u1_u15_u6_n104 ) , .A1( u1_u15_u6_n111 ) , .B1( u1_u15_u6_n124 ) , .B2( u1_u15_u6_n151 ) , .A2( u1_u15_u6_n93 ) );
  OAI211_X1 u1_u15_u6_U82 (.ZN( u1_out15_7 ) , .B( u1_u15_u6_n153 ) , .C2( u1_u15_u6_n154 ) , .C1( u1_u15_u6_n155 ) , .A( u1_u15_u6_n174 ) );
  NOR3_X1 u1_u15_u6_U83 (.A1( u1_u15_u6_n141 ) , .ZN( u1_u15_u6_n154 ) , .A3( u1_u15_u6_n164 ) , .A2( u1_u15_u6_n171 ) );
  AOI211_X1 u1_u15_u6_U84 (.B( u1_u15_u6_n149 ) , .A( u1_u15_u6_n150 ) , .C2( u1_u15_u6_n151 ) , .C1( u1_u15_u6_n152 ) , .ZN( u1_u15_u6_n153 ) );
  OAI211_X1 u1_u15_u6_U85 (.ZN( u1_out15_22 ) , .B( u1_u15_u6_n137 ) , .A( u1_u15_u6_n138 ) , .C2( u1_u15_u6_n139 ) , .C1( u1_u15_u6_n140 ) );
  AOI22_X1 u1_u15_u6_U86 (.B1( u1_u15_u6_n124 ) , .A2( u1_u15_u6_n125 ) , .A1( u1_u15_u6_n126 ) , .ZN( u1_u15_u6_n138 ) , .B2( u1_u15_u6_n161 ) );
  AND4_X1 u1_u15_u6_U87 (.A3( u1_u15_u6_n119 ) , .A1( u1_u15_u6_n120 ) , .A4( u1_u15_u6_n129 ) , .ZN( u1_u15_u6_n140 ) , .A2( u1_u15_u6_n143 ) );
  NAND3_X1 u1_u15_u6_U88 (.A2( u1_u15_u6_n123 ) , .ZN( u1_u15_u6_n125 ) , .A1( u1_u15_u6_n130 ) , .A3( u1_u15_u6_n131 ) );
  NAND3_X1 u1_u15_u6_U89 (.A3( u1_u15_u6_n133 ) , .ZN( u1_u15_u6_n141 ) , .A1( u1_u15_u6_n145 ) , .A2( u1_u15_u6_n148 ) );
  AOI21_X1 u1_u15_u6_U9 (.B2( u1_u15_u6_n147 ) , .B1( u1_u15_u6_n148 ) , .ZN( u1_u15_u6_n149 ) , .A( u1_u15_u6_n158 ) );
  NAND3_X1 u1_u15_u6_U90 (.ZN( u1_u15_u6_n101 ) , .A3( u1_u15_u6_n107 ) , .A2( u1_u15_u6_n121 ) , .A1( u1_u15_u6_n127 ) );
  NAND3_X1 u1_u15_u6_U91 (.ZN( u1_u15_u6_n102 ) , .A3( u1_u15_u6_n130 ) , .A2( u1_u15_u6_n145 ) , .A1( u1_u15_u6_n166 ) );
  NAND3_X1 u1_u15_u6_U92 (.A3( u1_u15_u6_n113 ) , .A1( u1_u15_u6_n119 ) , .A2( u1_u15_u6_n123 ) , .ZN( u1_u15_u6_n93 ) );
  NAND3_X1 u1_u15_u6_U93 (.ZN( u1_u15_u6_n142 ) , .A2( u1_u15_u6_n172 ) , .A3( u1_u15_u6_n89 ) , .A1( u1_u15_u6_n90 ) );
  OAI21_X1 u1_u15_u7_U10 (.A( u1_u15_u7_n161 ) , .B1( u1_u15_u7_n168 ) , .B2( u1_u15_u7_n173 ) , .ZN( u1_u15_u7_n91 ) );
  AOI211_X1 u1_u15_u7_U11 (.A( u1_u15_u7_n117 ) , .ZN( u1_u15_u7_n118 ) , .C2( u1_u15_u7_n126 ) , .C1( u1_u15_u7_n177 ) , .B( u1_u15_u7_n180 ) );
  OAI22_X1 u1_u15_u7_U12 (.B1( u1_u15_u7_n115 ) , .ZN( u1_u15_u7_n117 ) , .A2( u1_u15_u7_n133 ) , .A1( u1_u15_u7_n137 ) , .B2( u1_u15_u7_n162 ) );
  INV_X1 u1_u15_u7_U13 (.A( u1_u15_u7_n116 ) , .ZN( u1_u15_u7_n180 ) );
  NOR3_X1 u1_u15_u7_U14 (.ZN( u1_u15_u7_n115 ) , .A3( u1_u15_u7_n145 ) , .A2( u1_u15_u7_n168 ) , .A1( u1_u15_u7_n169 ) );
  OAI211_X1 u1_u15_u7_U15 (.B( u1_u15_u7_n122 ) , .A( u1_u15_u7_n123 ) , .C2( u1_u15_u7_n124 ) , .ZN( u1_u15_u7_n154 ) , .C1( u1_u15_u7_n162 ) );
  AOI222_X1 u1_u15_u7_U16 (.ZN( u1_u15_u7_n122 ) , .C2( u1_u15_u7_n126 ) , .C1( u1_u15_u7_n145 ) , .B1( u1_u15_u7_n161 ) , .A2( u1_u15_u7_n165 ) , .B2( u1_u15_u7_n170 ) , .A1( u1_u15_u7_n176 ) );
  INV_X1 u1_u15_u7_U17 (.A( u1_u15_u7_n133 ) , .ZN( u1_u15_u7_n176 ) );
  NOR3_X1 u1_u15_u7_U18 (.A2( u1_u15_u7_n134 ) , .A1( u1_u15_u7_n135 ) , .ZN( u1_u15_u7_n136 ) , .A3( u1_u15_u7_n171 ) );
  NOR2_X1 u1_u15_u7_U19 (.A1( u1_u15_u7_n130 ) , .A2( u1_u15_u7_n134 ) , .ZN( u1_u15_u7_n153 ) );
  INV_X1 u1_u15_u7_U20 (.A( u1_u15_u7_n101 ) , .ZN( u1_u15_u7_n165 ) );
  NOR2_X1 u1_u15_u7_U21 (.ZN( u1_u15_u7_n111 ) , .A2( u1_u15_u7_n134 ) , .A1( u1_u15_u7_n169 ) );
  AOI21_X1 u1_u15_u7_U22 (.ZN( u1_u15_u7_n104 ) , .B2( u1_u15_u7_n112 ) , .B1( u1_u15_u7_n127 ) , .A( u1_u15_u7_n164 ) );
  AOI21_X1 u1_u15_u7_U23 (.ZN( u1_u15_u7_n106 ) , .B1( u1_u15_u7_n133 ) , .B2( u1_u15_u7_n146 ) , .A( u1_u15_u7_n162 ) );
  AOI21_X1 u1_u15_u7_U24 (.A( u1_u15_u7_n101 ) , .ZN( u1_u15_u7_n107 ) , .B2( u1_u15_u7_n128 ) , .B1( u1_u15_u7_n175 ) );
  INV_X1 u1_u15_u7_U25 (.A( u1_u15_u7_n138 ) , .ZN( u1_u15_u7_n171 ) );
  INV_X1 u1_u15_u7_U26 (.A( u1_u15_u7_n131 ) , .ZN( u1_u15_u7_n177 ) );
  INV_X1 u1_u15_u7_U27 (.A( u1_u15_u7_n110 ) , .ZN( u1_u15_u7_n174 ) );
  NAND2_X1 u1_u15_u7_U28 (.A1( u1_u15_u7_n129 ) , .A2( u1_u15_u7_n132 ) , .ZN( u1_u15_u7_n149 ) );
  NAND2_X1 u1_u15_u7_U29 (.A1( u1_u15_u7_n113 ) , .A2( u1_u15_u7_n124 ) , .ZN( u1_u15_u7_n130 ) );
  INV_X1 u1_u15_u7_U3 (.A( u1_u15_u7_n111 ) , .ZN( u1_u15_u7_n170 ) );
  INV_X1 u1_u15_u7_U30 (.A( u1_u15_u7_n112 ) , .ZN( u1_u15_u7_n173 ) );
  INV_X1 u1_u15_u7_U31 (.A( u1_u15_u7_n128 ) , .ZN( u1_u15_u7_n168 ) );
  INV_X1 u1_u15_u7_U32 (.A( u1_u15_u7_n148 ) , .ZN( u1_u15_u7_n169 ) );
  INV_X1 u1_u15_u7_U33 (.A( u1_u15_u7_n127 ) , .ZN( u1_u15_u7_n179 ) );
  NOR2_X1 u1_u15_u7_U34 (.ZN( u1_u15_u7_n101 ) , .A2( u1_u15_u7_n150 ) , .A1( u1_u15_u7_n156 ) );
  AOI211_X1 u1_u15_u7_U35 (.B( u1_u15_u7_n154 ) , .A( u1_u15_u7_n155 ) , .C1( u1_u15_u7_n156 ) , .ZN( u1_u15_u7_n157 ) , .C2( u1_u15_u7_n172 ) );
  INV_X1 u1_u15_u7_U36 (.A( u1_u15_u7_n153 ) , .ZN( u1_u15_u7_n172 ) );
  AOI211_X1 u1_u15_u7_U37 (.B( u1_u15_u7_n139 ) , .A( u1_u15_u7_n140 ) , .C2( u1_u15_u7_n141 ) , .ZN( u1_u15_u7_n142 ) , .C1( u1_u15_u7_n156 ) );
  NAND4_X1 u1_u15_u7_U38 (.A3( u1_u15_u7_n127 ) , .A2( u1_u15_u7_n128 ) , .A1( u1_u15_u7_n129 ) , .ZN( u1_u15_u7_n141 ) , .A4( u1_u15_u7_n147 ) );
  AOI21_X1 u1_u15_u7_U39 (.A( u1_u15_u7_n137 ) , .B1( u1_u15_u7_n138 ) , .ZN( u1_u15_u7_n139 ) , .B2( u1_u15_u7_n146 ) );
  INV_X1 u1_u15_u7_U4 (.A( u1_u15_u7_n149 ) , .ZN( u1_u15_u7_n175 ) );
  OAI22_X1 u1_u15_u7_U40 (.B1( u1_u15_u7_n136 ) , .ZN( u1_u15_u7_n140 ) , .A1( u1_u15_u7_n153 ) , .B2( u1_u15_u7_n162 ) , .A2( u1_u15_u7_n164 ) );
  AOI21_X1 u1_u15_u7_U41 (.ZN( u1_u15_u7_n123 ) , .B1( u1_u15_u7_n165 ) , .B2( u1_u15_u7_n177 ) , .A( u1_u15_u7_n97 ) );
  AOI21_X1 u1_u15_u7_U42 (.B2( u1_u15_u7_n113 ) , .B1( u1_u15_u7_n124 ) , .A( u1_u15_u7_n125 ) , .ZN( u1_u15_u7_n97 ) );
  INV_X1 u1_u15_u7_U43 (.A( u1_u15_u7_n125 ) , .ZN( u1_u15_u7_n161 ) );
  INV_X1 u1_u15_u7_U44 (.A( u1_u15_u7_n152 ) , .ZN( u1_u15_u7_n162 ) );
  AOI22_X1 u1_u15_u7_U45 (.A2( u1_u15_u7_n114 ) , .ZN( u1_u15_u7_n119 ) , .B1( u1_u15_u7_n130 ) , .A1( u1_u15_u7_n156 ) , .B2( u1_u15_u7_n165 ) );
  NAND2_X1 u1_u15_u7_U46 (.A2( u1_u15_u7_n112 ) , .ZN( u1_u15_u7_n114 ) , .A1( u1_u15_u7_n175 ) );
  AOI22_X1 u1_u15_u7_U47 (.B2( u1_u15_u7_n149 ) , .B1( u1_u15_u7_n150 ) , .A2( u1_u15_u7_n151 ) , .A1( u1_u15_u7_n152 ) , .ZN( u1_u15_u7_n158 ) );
  AND2_X1 u1_u15_u7_U48 (.ZN( u1_u15_u7_n145 ) , .A2( u1_u15_u7_n98 ) , .A1( u1_u15_u7_n99 ) );
  NOR2_X1 u1_u15_u7_U49 (.ZN( u1_u15_u7_n137 ) , .A1( u1_u15_u7_n150 ) , .A2( u1_u15_u7_n161 ) );
  INV_X1 u1_u15_u7_U5 (.A( u1_u15_u7_n154 ) , .ZN( u1_u15_u7_n178 ) );
  AOI21_X1 u1_u15_u7_U50 (.ZN( u1_u15_u7_n105 ) , .B2( u1_u15_u7_n110 ) , .A( u1_u15_u7_n125 ) , .B1( u1_u15_u7_n147 ) );
  NAND2_X1 u1_u15_u7_U51 (.ZN( u1_u15_u7_n146 ) , .A1( u1_u15_u7_n95 ) , .A2( u1_u15_u7_n98 ) );
  NAND2_X1 u1_u15_u7_U52 (.A2( u1_u15_u7_n103 ) , .ZN( u1_u15_u7_n147 ) , .A1( u1_u15_u7_n93 ) );
  NAND2_X1 u1_u15_u7_U53 (.A1( u1_u15_u7_n103 ) , .ZN( u1_u15_u7_n127 ) , .A2( u1_u15_u7_n99 ) );
  OR2_X1 u1_u15_u7_U54 (.ZN( u1_u15_u7_n126 ) , .A2( u1_u15_u7_n152 ) , .A1( u1_u15_u7_n156 ) );
  NAND2_X1 u1_u15_u7_U55 (.A2( u1_u15_u7_n102 ) , .A1( u1_u15_u7_n103 ) , .ZN( u1_u15_u7_n133 ) );
  NAND2_X1 u1_u15_u7_U56 (.ZN( u1_u15_u7_n112 ) , .A2( u1_u15_u7_n96 ) , .A1( u1_u15_u7_n99 ) );
  NAND2_X1 u1_u15_u7_U57 (.A2( u1_u15_u7_n102 ) , .ZN( u1_u15_u7_n128 ) , .A1( u1_u15_u7_n98 ) );
  NAND2_X1 u1_u15_u7_U58 (.A1( u1_u15_u7_n100 ) , .ZN( u1_u15_u7_n113 ) , .A2( u1_u15_u7_n93 ) );
  NAND2_X1 u1_u15_u7_U59 (.A2( u1_u15_u7_n102 ) , .ZN( u1_u15_u7_n124 ) , .A1( u1_u15_u7_n96 ) );
  AOI211_X1 u1_u15_u7_U6 (.ZN( u1_u15_u7_n116 ) , .A( u1_u15_u7_n155 ) , .C1( u1_u15_u7_n161 ) , .C2( u1_u15_u7_n171 ) , .B( u1_u15_u7_n94 ) );
  NAND2_X1 u1_u15_u7_U60 (.ZN( u1_u15_u7_n110 ) , .A1( u1_u15_u7_n95 ) , .A2( u1_u15_u7_n96 ) );
  INV_X1 u1_u15_u7_U61 (.A( u1_u15_u7_n150 ) , .ZN( u1_u15_u7_n164 ) );
  AND2_X1 u1_u15_u7_U62 (.ZN( u1_u15_u7_n134 ) , .A1( u1_u15_u7_n93 ) , .A2( u1_u15_u7_n98 ) );
  NAND2_X1 u1_u15_u7_U63 (.A1( u1_u15_u7_n100 ) , .A2( u1_u15_u7_n102 ) , .ZN( u1_u15_u7_n129 ) );
  NAND2_X1 u1_u15_u7_U64 (.A2( u1_u15_u7_n103 ) , .ZN( u1_u15_u7_n131 ) , .A1( u1_u15_u7_n95 ) );
  NAND2_X1 u1_u15_u7_U65 (.A1( u1_u15_u7_n100 ) , .ZN( u1_u15_u7_n138 ) , .A2( u1_u15_u7_n99 ) );
  NAND2_X1 u1_u15_u7_U66 (.ZN( u1_u15_u7_n132 ) , .A1( u1_u15_u7_n93 ) , .A2( u1_u15_u7_n96 ) );
  NAND2_X1 u1_u15_u7_U67 (.A1( u1_u15_u7_n100 ) , .ZN( u1_u15_u7_n148 ) , .A2( u1_u15_u7_n95 ) );
  NOR2_X1 u1_u15_u7_U68 (.A2( u1_u15_X_47 ) , .ZN( u1_u15_u7_n150 ) , .A1( u1_u15_u7_n163 ) );
  NOR2_X1 u1_u15_u7_U69 (.A2( u1_u15_X_43 ) , .A1( u1_u15_X_44 ) , .ZN( u1_u15_u7_n103 ) );
  OAI222_X1 u1_u15_u7_U7 (.C2( u1_u15_u7_n101 ) , .B2( u1_u15_u7_n111 ) , .A1( u1_u15_u7_n113 ) , .C1( u1_u15_u7_n146 ) , .A2( u1_u15_u7_n162 ) , .B1( u1_u15_u7_n164 ) , .ZN( u1_u15_u7_n94 ) );
  NOR2_X1 u1_u15_u7_U70 (.A2( u1_u15_X_48 ) , .A1( u1_u15_u7_n166 ) , .ZN( u1_u15_u7_n95 ) );
  NOR2_X1 u1_u15_u7_U71 (.A2( u1_u15_X_45 ) , .A1( u1_u15_X_48 ) , .ZN( u1_u15_u7_n99 ) );
  NOR2_X1 u1_u15_u7_U72 (.A2( u1_u15_X_44 ) , .A1( u1_u15_u7_n167 ) , .ZN( u1_u15_u7_n98 ) );
  NOR2_X1 u1_u15_u7_U73 (.A2( u1_u15_X_46 ) , .A1( u1_u15_X_47 ) , .ZN( u1_u15_u7_n152 ) );
  AND2_X1 u1_u15_u7_U74 (.A1( u1_u15_X_47 ) , .ZN( u1_u15_u7_n156 ) , .A2( u1_u15_u7_n163 ) );
  NAND2_X1 u1_u15_u7_U75 (.A2( u1_u15_X_46 ) , .A1( u1_u15_X_47 ) , .ZN( u1_u15_u7_n125 ) );
  AND2_X1 u1_u15_u7_U76 (.A2( u1_u15_X_45 ) , .A1( u1_u15_X_48 ) , .ZN( u1_u15_u7_n102 ) );
  AND2_X1 u1_u15_u7_U77 (.A2( u1_u15_X_43 ) , .A1( u1_u15_X_44 ) , .ZN( u1_u15_u7_n96 ) );
  AND2_X1 u1_u15_u7_U78 (.A1( u1_u15_X_44 ) , .ZN( u1_u15_u7_n100 ) , .A2( u1_u15_u7_n167 ) );
  AND2_X1 u1_u15_u7_U79 (.A1( u1_u15_X_48 ) , .A2( u1_u15_u7_n166 ) , .ZN( u1_u15_u7_n93 ) );
  OAI221_X1 u1_u15_u7_U8 (.C1( u1_u15_u7_n101 ) , .C2( u1_u15_u7_n147 ) , .ZN( u1_u15_u7_n155 ) , .B2( u1_u15_u7_n162 ) , .A( u1_u15_u7_n91 ) , .B1( u1_u15_u7_n92 ) );
  INV_X1 u1_u15_u7_U80 (.A( u1_u15_X_46 ) , .ZN( u1_u15_u7_n163 ) );
  INV_X1 u1_u15_u7_U81 (.A( u1_u15_X_45 ) , .ZN( u1_u15_u7_n166 ) );
  INV_X1 u1_u15_u7_U82 (.A( u1_u15_X_43 ) , .ZN( u1_u15_u7_n167 ) );
  NAND4_X1 u1_u15_u7_U83 (.ZN( u1_out15_5 ) , .A4( u1_u15_u7_n108 ) , .A3( u1_u15_u7_n109 ) , .A1( u1_u15_u7_n116 ) , .A2( u1_u15_u7_n123 ) );
  AOI22_X1 u1_u15_u7_U84 (.ZN( u1_u15_u7_n109 ) , .A2( u1_u15_u7_n126 ) , .B2( u1_u15_u7_n145 ) , .B1( u1_u15_u7_n156 ) , .A1( u1_u15_u7_n171 ) );
  NOR4_X1 u1_u15_u7_U85 (.A4( u1_u15_u7_n104 ) , .A3( u1_u15_u7_n105 ) , .A2( u1_u15_u7_n106 ) , .A1( u1_u15_u7_n107 ) , .ZN( u1_u15_u7_n108 ) );
  NAND4_X1 u1_u15_u7_U86 (.ZN( u1_out15_27 ) , .A4( u1_u15_u7_n118 ) , .A3( u1_u15_u7_n119 ) , .A2( u1_u15_u7_n120 ) , .A1( u1_u15_u7_n121 ) );
  OAI21_X1 u1_u15_u7_U87 (.ZN( u1_u15_u7_n121 ) , .B2( u1_u15_u7_n145 ) , .A( u1_u15_u7_n150 ) , .B1( u1_u15_u7_n174 ) );
  OAI21_X1 u1_u15_u7_U88 (.ZN( u1_u15_u7_n120 ) , .A( u1_u15_u7_n161 ) , .B2( u1_u15_u7_n170 ) , .B1( u1_u15_u7_n179 ) );
  NAND4_X1 u1_u15_u7_U89 (.ZN( u1_out15_21 ) , .A4( u1_u15_u7_n157 ) , .A3( u1_u15_u7_n158 ) , .A2( u1_u15_u7_n159 ) , .A1( u1_u15_u7_n160 ) );
  AND3_X1 u1_u15_u7_U9 (.A3( u1_u15_u7_n110 ) , .A2( u1_u15_u7_n127 ) , .A1( u1_u15_u7_n132 ) , .ZN( u1_u15_u7_n92 ) );
  OAI21_X1 u1_u15_u7_U90 (.B1( u1_u15_u7_n145 ) , .ZN( u1_u15_u7_n160 ) , .A( u1_u15_u7_n161 ) , .B2( u1_u15_u7_n177 ) );
  OAI21_X1 u1_u15_u7_U91 (.ZN( u1_u15_u7_n159 ) , .A( u1_u15_u7_n165 ) , .B2( u1_u15_u7_n171 ) , .B1( u1_u15_u7_n174 ) );
  NAND4_X1 u1_u15_u7_U92 (.ZN( u1_out15_15 ) , .A4( u1_u15_u7_n142 ) , .A3( u1_u15_u7_n143 ) , .A2( u1_u15_u7_n144 ) , .A1( u1_u15_u7_n178 ) );
  OR2_X1 u1_u15_u7_U93 (.A2( u1_u15_u7_n125 ) , .A1( u1_u15_u7_n129 ) , .ZN( u1_u15_u7_n144 ) );
  AOI22_X1 u1_u15_u7_U94 (.A2( u1_u15_u7_n126 ) , .ZN( u1_u15_u7_n143 ) , .B2( u1_u15_u7_n165 ) , .B1( u1_u15_u7_n173 ) , .A1( u1_u15_u7_n174 ) );
  NAND3_X1 u1_u15_u7_U95 (.A3( u1_u15_u7_n146 ) , .A2( u1_u15_u7_n147 ) , .A1( u1_u15_u7_n148 ) , .ZN( u1_u15_u7_n151 ) );
  NAND3_X1 u1_u15_u7_U96 (.A3( u1_u15_u7_n131 ) , .A2( u1_u15_u7_n132 ) , .A1( u1_u15_u7_n133 ) , .ZN( u1_u15_u7_n135 ) );
  XOR2_X1 u1_u1_U16 (.B( u1_K2_3 ) , .A( u1_R0_2 ) , .Z( u1_u1_X_3 ) );
  XOR2_X1 u1_u1_U27 (.B( u1_K2_2 ) , .A( u1_R0_1 ) , .Z( u1_u1_X_2 ) );
  XOR2_X1 u1_u1_U38 (.B( u1_K2_1 ) , .A( u1_R0_32 ) , .Z( u1_u1_X_1 ) );
  XOR2_X1 u1_u1_U4 (.B( u1_K2_6 ) , .A( u1_R0_5 ) , .Z( u1_u1_X_6 ) );
  XOR2_X1 u1_u1_U5 (.B( u1_K2_5 ) , .A( u1_R0_4 ) , .Z( u1_u1_X_5 ) );
  XOR2_X1 u1_u1_U6 (.B( u1_K2_4 ) , .A( u1_R0_3 ) , .Z( u1_u1_X_4 ) );
  AND3_X1 u1_u1_u0_U10 (.A2( u1_u1_u0_n112 ) , .ZN( u1_u1_u0_n127 ) , .A3( u1_u1_u0_n130 ) , .A1( u1_u1_u0_n148 ) );
  NAND2_X1 u1_u1_u0_U11 (.ZN( u1_u1_u0_n113 ) , .A1( u1_u1_u0_n139 ) , .A2( u1_u1_u0_n149 ) );
  AND2_X1 u1_u1_u0_U12 (.ZN( u1_u1_u0_n107 ) , .A1( u1_u1_u0_n130 ) , .A2( u1_u1_u0_n140 ) );
  AND2_X1 u1_u1_u0_U13 (.A2( u1_u1_u0_n129 ) , .A1( u1_u1_u0_n130 ) , .ZN( u1_u1_u0_n151 ) );
  AND2_X1 u1_u1_u0_U14 (.A1( u1_u1_u0_n108 ) , .A2( u1_u1_u0_n125 ) , .ZN( u1_u1_u0_n145 ) );
  INV_X1 u1_u1_u0_U15 (.A( u1_u1_u0_n143 ) , .ZN( u1_u1_u0_n173 ) );
  NOR2_X1 u1_u1_u0_U16 (.A2( u1_u1_u0_n136 ) , .ZN( u1_u1_u0_n147 ) , .A1( u1_u1_u0_n160 ) );
  NOR2_X1 u1_u1_u0_U17 (.A1( u1_u1_u0_n163 ) , .A2( u1_u1_u0_n164 ) , .ZN( u1_u1_u0_n95 ) );
  AOI21_X1 u1_u1_u0_U18 (.B1( u1_u1_u0_n103 ) , .ZN( u1_u1_u0_n132 ) , .A( u1_u1_u0_n165 ) , .B2( u1_u1_u0_n93 ) );
  INV_X1 u1_u1_u0_U19 (.A( u1_u1_u0_n142 ) , .ZN( u1_u1_u0_n165 ) );
  OAI221_X1 u1_u1_u0_U20 (.C1( u1_u1_u0_n121 ) , .ZN( u1_u1_u0_n122 ) , .B2( u1_u1_u0_n127 ) , .A( u1_u1_u0_n143 ) , .B1( u1_u1_u0_n144 ) , .C2( u1_u1_u0_n147 ) );
  OAI22_X1 u1_u1_u0_U21 (.B1( u1_u1_u0_n125 ) , .ZN( u1_u1_u0_n126 ) , .A1( u1_u1_u0_n138 ) , .A2( u1_u1_u0_n146 ) , .B2( u1_u1_u0_n147 ) );
  OAI22_X1 u1_u1_u0_U22 (.B1( u1_u1_u0_n131 ) , .A1( u1_u1_u0_n144 ) , .B2( u1_u1_u0_n147 ) , .A2( u1_u1_u0_n90 ) , .ZN( u1_u1_u0_n91 ) );
  AND3_X1 u1_u1_u0_U23 (.A3( u1_u1_u0_n121 ) , .A2( u1_u1_u0_n125 ) , .A1( u1_u1_u0_n148 ) , .ZN( u1_u1_u0_n90 ) );
  INV_X1 u1_u1_u0_U24 (.A( u1_u1_u0_n136 ) , .ZN( u1_u1_u0_n161 ) );
  NOR2_X1 u1_u1_u0_U25 (.A1( u1_u1_u0_n120 ) , .ZN( u1_u1_u0_n143 ) , .A2( u1_u1_u0_n167 ) );
  OAI221_X1 u1_u1_u0_U26 (.C1( u1_u1_u0_n112 ) , .ZN( u1_u1_u0_n120 ) , .B1( u1_u1_u0_n138 ) , .B2( u1_u1_u0_n141 ) , .C2( u1_u1_u0_n147 ) , .A( u1_u1_u0_n172 ) );
  AOI211_X1 u1_u1_u0_U27 (.B( u1_u1_u0_n115 ) , .A( u1_u1_u0_n116 ) , .C2( u1_u1_u0_n117 ) , .C1( u1_u1_u0_n118 ) , .ZN( u1_u1_u0_n119 ) );
  AOI22_X1 u1_u1_u0_U28 (.B2( u1_u1_u0_n109 ) , .A2( u1_u1_u0_n110 ) , .ZN( u1_u1_u0_n111 ) , .B1( u1_u1_u0_n118 ) , .A1( u1_u1_u0_n160 ) );
  INV_X1 u1_u1_u0_U29 (.A( u1_u1_u0_n118 ) , .ZN( u1_u1_u0_n158 ) );
  INV_X1 u1_u1_u0_U3 (.A( u1_u1_u0_n113 ) , .ZN( u1_u1_u0_n166 ) );
  AOI21_X1 u1_u1_u0_U30 (.ZN( u1_u1_u0_n104 ) , .B1( u1_u1_u0_n107 ) , .B2( u1_u1_u0_n141 ) , .A( u1_u1_u0_n144 ) );
  AOI21_X1 u1_u1_u0_U31 (.B1( u1_u1_u0_n127 ) , .B2( u1_u1_u0_n129 ) , .A( u1_u1_u0_n138 ) , .ZN( u1_u1_u0_n96 ) );
  AOI21_X1 u1_u1_u0_U32 (.ZN( u1_u1_u0_n116 ) , .B2( u1_u1_u0_n142 ) , .A( u1_u1_u0_n144 ) , .B1( u1_u1_u0_n166 ) );
  NAND2_X1 u1_u1_u0_U33 (.A1( u1_u1_u0_n100 ) , .A2( u1_u1_u0_n103 ) , .ZN( u1_u1_u0_n125 ) );
  NAND2_X1 u1_u1_u0_U34 (.A2( u1_u1_u0_n103 ) , .ZN( u1_u1_u0_n140 ) , .A1( u1_u1_u0_n94 ) );
  NAND2_X1 u1_u1_u0_U35 (.A1( u1_u1_u0_n101 ) , .A2( u1_u1_u0_n102 ) , .ZN( u1_u1_u0_n150 ) );
  INV_X1 u1_u1_u0_U36 (.A( u1_u1_u0_n138 ) , .ZN( u1_u1_u0_n160 ) );
  NAND2_X1 u1_u1_u0_U37 (.ZN( u1_u1_u0_n142 ) , .A1( u1_u1_u0_n94 ) , .A2( u1_u1_u0_n95 ) );
  NAND2_X1 u1_u1_u0_U38 (.A1( u1_u1_u0_n102 ) , .ZN( u1_u1_u0_n128 ) , .A2( u1_u1_u0_n95 ) );
  NAND2_X1 u1_u1_u0_U39 (.A2( u1_u1_u0_n102 ) , .A1( u1_u1_u0_n103 ) , .ZN( u1_u1_u0_n149 ) );
  AOI21_X1 u1_u1_u0_U4 (.B1( u1_u1_u0_n114 ) , .ZN( u1_u1_u0_n115 ) , .B2( u1_u1_u0_n129 ) , .A( u1_u1_u0_n161 ) );
  NAND2_X1 u1_u1_u0_U40 (.A1( u1_u1_u0_n100 ) , .ZN( u1_u1_u0_n129 ) , .A2( u1_u1_u0_n95 ) );
  NAND2_X1 u1_u1_u0_U41 (.A2( u1_u1_u0_n100 ) , .A1( u1_u1_u0_n101 ) , .ZN( u1_u1_u0_n139 ) );
  NAND2_X1 u1_u1_u0_U42 (.A2( u1_u1_u0_n100 ) , .ZN( u1_u1_u0_n131 ) , .A1( u1_u1_u0_n92 ) );
  NAND2_X1 u1_u1_u0_U43 (.ZN( u1_u1_u0_n108 ) , .A1( u1_u1_u0_n92 ) , .A2( u1_u1_u0_n94 ) );
  NAND2_X1 u1_u1_u0_U44 (.ZN( u1_u1_u0_n148 ) , .A1( u1_u1_u0_n93 ) , .A2( u1_u1_u0_n95 ) );
  NAND2_X1 u1_u1_u0_U45 (.A2( u1_u1_u0_n102 ) , .ZN( u1_u1_u0_n114 ) , .A1( u1_u1_u0_n92 ) );
  NAND2_X1 u1_u1_u0_U46 (.A1( u1_u1_u0_n101 ) , .ZN( u1_u1_u0_n130 ) , .A2( u1_u1_u0_n94 ) );
  NAND2_X1 u1_u1_u0_U47 (.A2( u1_u1_u0_n101 ) , .ZN( u1_u1_u0_n121 ) , .A1( u1_u1_u0_n93 ) );
  INV_X1 u1_u1_u0_U48 (.ZN( u1_u1_u0_n172 ) , .A( u1_u1_u0_n88 ) );
  OAI222_X1 u1_u1_u0_U49 (.C1( u1_u1_u0_n108 ) , .A1( u1_u1_u0_n125 ) , .B2( u1_u1_u0_n128 ) , .B1( u1_u1_u0_n144 ) , .A2( u1_u1_u0_n158 ) , .C2( u1_u1_u0_n161 ) , .ZN( u1_u1_u0_n88 ) );
  AOI21_X1 u1_u1_u0_U5 (.B2( u1_u1_u0_n131 ) , .ZN( u1_u1_u0_n134 ) , .B1( u1_u1_u0_n151 ) , .A( u1_u1_u0_n158 ) );
  NAND2_X1 u1_u1_u0_U50 (.ZN( u1_u1_u0_n112 ) , .A2( u1_u1_u0_n92 ) , .A1( u1_u1_u0_n93 ) );
  OR3_X1 u1_u1_u0_U51 (.A3( u1_u1_u0_n152 ) , .A2( u1_u1_u0_n153 ) , .A1( u1_u1_u0_n154 ) , .ZN( u1_u1_u0_n155 ) );
  AOI21_X1 u1_u1_u0_U52 (.B2( u1_u1_u0_n150 ) , .B1( u1_u1_u0_n151 ) , .ZN( u1_u1_u0_n152 ) , .A( u1_u1_u0_n158 ) );
  AOI21_X1 u1_u1_u0_U53 (.A( u1_u1_u0_n144 ) , .B2( u1_u1_u0_n145 ) , .B1( u1_u1_u0_n146 ) , .ZN( u1_u1_u0_n154 ) );
  AOI21_X1 u1_u1_u0_U54 (.A( u1_u1_u0_n147 ) , .B2( u1_u1_u0_n148 ) , .B1( u1_u1_u0_n149 ) , .ZN( u1_u1_u0_n153 ) );
  INV_X1 u1_u1_u0_U55 (.ZN( u1_u1_u0_n171 ) , .A( u1_u1_u0_n99 ) );
  OAI211_X1 u1_u1_u0_U56 (.C2( u1_u1_u0_n140 ) , .C1( u1_u1_u0_n161 ) , .A( u1_u1_u0_n169 ) , .B( u1_u1_u0_n98 ) , .ZN( u1_u1_u0_n99 ) );
  INV_X1 u1_u1_u0_U57 (.ZN( u1_u1_u0_n169 ) , .A( u1_u1_u0_n91 ) );
  AOI211_X1 u1_u1_u0_U58 (.C1( u1_u1_u0_n118 ) , .A( u1_u1_u0_n123 ) , .B( u1_u1_u0_n96 ) , .C2( u1_u1_u0_n97 ) , .ZN( u1_u1_u0_n98 ) );
  NOR2_X1 u1_u1_u0_U59 (.A2( u1_u1_X_2 ) , .ZN( u1_u1_u0_n103 ) , .A1( u1_u1_u0_n164 ) );
  NOR2_X1 u1_u1_u0_U6 (.A1( u1_u1_u0_n108 ) , .ZN( u1_u1_u0_n123 ) , .A2( u1_u1_u0_n158 ) );
  NOR2_X1 u1_u1_u0_U60 (.A2( u1_u1_X_3 ) , .A1( u1_u1_X_6 ) , .ZN( u1_u1_u0_n94 ) );
  NOR2_X1 u1_u1_u0_U61 (.A2( u1_u1_X_6 ) , .ZN( u1_u1_u0_n100 ) , .A1( u1_u1_u0_n162 ) );
  NOR2_X1 u1_u1_u0_U62 (.A2( u1_u1_X_4 ) , .A1( u1_u1_X_5 ) , .ZN( u1_u1_u0_n118 ) );
  NOR2_X1 u1_u1_u0_U63 (.A2( u1_u1_X_1 ) , .A1( u1_u1_X_2 ) , .ZN( u1_u1_u0_n92 ) );
  NOR2_X1 u1_u1_u0_U64 (.A2( u1_u1_X_1 ) , .ZN( u1_u1_u0_n101 ) , .A1( u1_u1_u0_n163 ) );
  NAND2_X1 u1_u1_u0_U65 (.A2( u1_u1_X_4 ) , .A1( u1_u1_X_5 ) , .ZN( u1_u1_u0_n144 ) );
  NOR2_X1 u1_u1_u0_U66 (.A2( u1_u1_X_5 ) , .ZN( u1_u1_u0_n136 ) , .A1( u1_u1_u0_n159 ) );
  NAND2_X1 u1_u1_u0_U67 (.A1( u1_u1_X_5 ) , .ZN( u1_u1_u0_n138 ) , .A2( u1_u1_u0_n159 ) );
  AND2_X1 u1_u1_u0_U68 (.A2( u1_u1_X_3 ) , .A1( u1_u1_X_6 ) , .ZN( u1_u1_u0_n102 ) );
  AND2_X1 u1_u1_u0_U69 (.A1( u1_u1_X_6 ) , .A2( u1_u1_u0_n162 ) , .ZN( u1_u1_u0_n93 ) );
  OAI21_X1 u1_u1_u0_U7 (.B1( u1_u1_u0_n150 ) , .B2( u1_u1_u0_n158 ) , .A( u1_u1_u0_n172 ) , .ZN( u1_u1_u0_n89 ) );
  INV_X1 u1_u1_u0_U70 (.A( u1_u1_X_4 ) , .ZN( u1_u1_u0_n159 ) );
  INV_X1 u1_u1_u0_U71 (.A( u1_u1_X_1 ) , .ZN( u1_u1_u0_n164 ) );
  INV_X1 u1_u1_u0_U72 (.A( u1_u1_X_2 ) , .ZN( u1_u1_u0_n163 ) );
  INV_X1 u1_u1_u0_U73 (.A( u1_u1_X_3 ) , .ZN( u1_u1_u0_n162 ) );
  INV_X1 u1_u1_u0_U74 (.A( u1_u1_u0_n126 ) , .ZN( u1_u1_u0_n168 ) );
  AOI211_X1 u1_u1_u0_U75 (.B( u1_u1_u0_n133 ) , .A( u1_u1_u0_n134 ) , .C2( u1_u1_u0_n135 ) , .C1( u1_u1_u0_n136 ) , .ZN( u1_u1_u0_n137 ) );
  INV_X1 u1_u1_u0_U76 (.ZN( u1_u1_u0_n174 ) , .A( u1_u1_u0_n89 ) );
  AOI211_X1 u1_u1_u0_U77 (.B( u1_u1_u0_n104 ) , .A( u1_u1_u0_n105 ) , .ZN( u1_u1_u0_n106 ) , .C2( u1_u1_u0_n113 ) , .C1( u1_u1_u0_n160 ) );
  OR4_X1 u1_u1_u0_U78 (.ZN( u1_out1_17 ) , .A4( u1_u1_u0_n122 ) , .A2( u1_u1_u0_n123 ) , .A1( u1_u1_u0_n124 ) , .A3( u1_u1_u0_n170 ) );
  AOI21_X1 u1_u1_u0_U79 (.B2( u1_u1_u0_n107 ) , .ZN( u1_u1_u0_n124 ) , .B1( u1_u1_u0_n128 ) , .A( u1_u1_u0_n161 ) );
  AND2_X1 u1_u1_u0_U8 (.A1( u1_u1_u0_n114 ) , .A2( u1_u1_u0_n121 ) , .ZN( u1_u1_u0_n146 ) );
  INV_X1 u1_u1_u0_U80 (.A( u1_u1_u0_n111 ) , .ZN( u1_u1_u0_n170 ) );
  OR4_X1 u1_u1_u0_U81 (.ZN( u1_out1_31 ) , .A4( u1_u1_u0_n155 ) , .A2( u1_u1_u0_n156 ) , .A1( u1_u1_u0_n157 ) , .A3( u1_u1_u0_n173 ) );
  AOI21_X1 u1_u1_u0_U82 (.A( u1_u1_u0_n138 ) , .B2( u1_u1_u0_n139 ) , .B1( u1_u1_u0_n140 ) , .ZN( u1_u1_u0_n157 ) );
  AOI21_X1 u1_u1_u0_U83 (.B2( u1_u1_u0_n141 ) , .B1( u1_u1_u0_n142 ) , .ZN( u1_u1_u0_n156 ) , .A( u1_u1_u0_n161 ) );
  AOI21_X1 u1_u1_u0_U84 (.B1( u1_u1_u0_n132 ) , .ZN( u1_u1_u0_n133 ) , .A( u1_u1_u0_n144 ) , .B2( u1_u1_u0_n166 ) );
  OAI22_X1 u1_u1_u0_U85 (.ZN( u1_u1_u0_n105 ) , .A2( u1_u1_u0_n132 ) , .B1( u1_u1_u0_n146 ) , .A1( u1_u1_u0_n147 ) , .B2( u1_u1_u0_n161 ) );
  NAND2_X1 u1_u1_u0_U86 (.ZN( u1_u1_u0_n110 ) , .A2( u1_u1_u0_n132 ) , .A1( u1_u1_u0_n145 ) );
  INV_X1 u1_u1_u0_U87 (.A( u1_u1_u0_n119 ) , .ZN( u1_u1_u0_n167 ) );
  NAND3_X1 u1_u1_u0_U88 (.ZN( u1_out1_23 ) , .A3( u1_u1_u0_n137 ) , .A1( u1_u1_u0_n168 ) , .A2( u1_u1_u0_n171 ) );
  NAND3_X1 u1_u1_u0_U89 (.A3( u1_u1_u0_n127 ) , .A2( u1_u1_u0_n128 ) , .ZN( u1_u1_u0_n135 ) , .A1( u1_u1_u0_n150 ) );
  AND2_X1 u1_u1_u0_U9 (.A1( u1_u1_u0_n131 ) , .ZN( u1_u1_u0_n141 ) , .A2( u1_u1_u0_n150 ) );
  NAND3_X1 u1_u1_u0_U90 (.ZN( u1_u1_u0_n117 ) , .A3( u1_u1_u0_n132 ) , .A2( u1_u1_u0_n139 ) , .A1( u1_u1_u0_n148 ) );
  NAND3_X1 u1_u1_u0_U91 (.ZN( u1_u1_u0_n109 ) , .A2( u1_u1_u0_n114 ) , .A3( u1_u1_u0_n140 ) , .A1( u1_u1_u0_n149 ) );
  NAND3_X1 u1_u1_u0_U92 (.ZN( u1_out1_9 ) , .A3( u1_u1_u0_n106 ) , .A2( u1_u1_u0_n171 ) , .A1( u1_u1_u0_n174 ) );
  NAND3_X1 u1_u1_u0_U93 (.A2( u1_u1_u0_n128 ) , .A1( u1_u1_u0_n132 ) , .A3( u1_u1_u0_n146 ) , .ZN( u1_u1_u0_n97 ) );
  XOR2_X1 u1_u3_U13 (.B( u1_K4_42 ) , .A( u1_R2_29 ) , .Z( u1_u3_X_42 ) );
  XOR2_X1 u1_u3_U14 (.B( u1_K4_41 ) , .A( u1_R2_28 ) , .Z( u1_u3_X_41 ) );
  XOR2_X1 u1_u3_U15 (.B( u1_K4_40 ) , .A( u1_R2_27 ) , .Z( u1_u3_X_40 ) );
  XOR2_X1 u1_u3_U17 (.B( u1_K4_39 ) , .A( u1_R2_26 ) , .Z( u1_u3_X_39 ) );
  XOR2_X1 u1_u3_U18 (.B( u1_K4_38 ) , .A( u1_R2_25 ) , .Z( u1_u3_X_38 ) );
  XOR2_X1 u1_u3_U19 (.B( u1_K4_37 ) , .A( u1_R2_24 ) , .Z( u1_u3_X_37 ) );
  XOR2_X1 u1_u3_U20 (.B( u1_K4_36 ) , .A( u1_R2_25 ) , .Z( u1_u3_X_36 ) );
  XOR2_X1 u1_u3_U21 (.B( u1_K4_35 ) , .A( u1_R2_24 ) , .Z( u1_u3_X_35 ) );
  XOR2_X1 u1_u3_U22 (.B( u1_K4_34 ) , .A( u1_R2_23 ) , .Z( u1_u3_X_34 ) );
  XOR2_X1 u1_u3_U23 (.B( u1_K4_33 ) , .A( u1_R2_22 ) , .Z( u1_u3_X_33 ) );
  XOR2_X1 u1_u3_U24 (.B( u1_K4_32 ) , .A( u1_R2_21 ) , .Z( u1_u3_X_32 ) );
  XOR2_X1 u1_u3_U25 (.B( u1_K4_31 ) , .A( u1_R2_20 ) , .Z( u1_u3_X_31 ) );
  INV_X1 u1_u3_u5_U10 (.A( u1_u3_u5_n121 ) , .ZN( u1_u3_u5_n177 ) );
  NOR3_X1 u1_u3_u5_U100 (.A3( u1_u3_u5_n141 ) , .A1( u1_u3_u5_n142 ) , .ZN( u1_u3_u5_n143 ) , .A2( u1_u3_u5_n191 ) );
  NAND4_X1 u1_u3_u5_U101 (.ZN( u1_out3_4 ) , .A4( u1_u3_u5_n112 ) , .A2( u1_u3_u5_n113 ) , .A1( u1_u3_u5_n114 ) , .A3( u1_u3_u5_n195 ) );
  AOI211_X1 u1_u3_u5_U102 (.A( u1_u3_u5_n110 ) , .C1( u1_u3_u5_n111 ) , .ZN( u1_u3_u5_n112 ) , .B( u1_u3_u5_n118 ) , .C2( u1_u3_u5_n177 ) );
  AOI222_X1 u1_u3_u5_U103 (.ZN( u1_u3_u5_n113 ) , .A1( u1_u3_u5_n131 ) , .C1( u1_u3_u5_n148 ) , .B2( u1_u3_u5_n174 ) , .C2( u1_u3_u5_n178 ) , .A2( u1_u3_u5_n179 ) , .B1( u1_u3_u5_n99 ) );
  NAND3_X1 u1_u3_u5_U104 (.A2( u1_u3_u5_n154 ) , .A3( u1_u3_u5_n158 ) , .A1( u1_u3_u5_n161 ) , .ZN( u1_u3_u5_n99 ) );
  NOR2_X1 u1_u3_u5_U11 (.ZN( u1_u3_u5_n160 ) , .A2( u1_u3_u5_n173 ) , .A1( u1_u3_u5_n177 ) );
  INV_X1 u1_u3_u5_U12 (.A( u1_u3_u5_n150 ) , .ZN( u1_u3_u5_n174 ) );
  AOI21_X1 u1_u3_u5_U13 (.A( u1_u3_u5_n160 ) , .B2( u1_u3_u5_n161 ) , .ZN( u1_u3_u5_n162 ) , .B1( u1_u3_u5_n192 ) );
  INV_X1 u1_u3_u5_U14 (.A( u1_u3_u5_n159 ) , .ZN( u1_u3_u5_n192 ) );
  AOI21_X1 u1_u3_u5_U15 (.A( u1_u3_u5_n156 ) , .B2( u1_u3_u5_n157 ) , .B1( u1_u3_u5_n158 ) , .ZN( u1_u3_u5_n163 ) );
  AOI21_X1 u1_u3_u5_U16 (.B2( u1_u3_u5_n139 ) , .B1( u1_u3_u5_n140 ) , .ZN( u1_u3_u5_n141 ) , .A( u1_u3_u5_n150 ) );
  OAI21_X1 u1_u3_u5_U17 (.A( u1_u3_u5_n133 ) , .B2( u1_u3_u5_n134 ) , .B1( u1_u3_u5_n135 ) , .ZN( u1_u3_u5_n142 ) );
  OAI21_X1 u1_u3_u5_U18 (.ZN( u1_u3_u5_n133 ) , .B2( u1_u3_u5_n147 ) , .A( u1_u3_u5_n173 ) , .B1( u1_u3_u5_n188 ) );
  NAND2_X1 u1_u3_u5_U19 (.A2( u1_u3_u5_n119 ) , .A1( u1_u3_u5_n123 ) , .ZN( u1_u3_u5_n137 ) );
  INV_X1 u1_u3_u5_U20 (.A( u1_u3_u5_n155 ) , .ZN( u1_u3_u5_n194 ) );
  NAND2_X1 u1_u3_u5_U21 (.A1( u1_u3_u5_n121 ) , .ZN( u1_u3_u5_n132 ) , .A2( u1_u3_u5_n172 ) );
  NAND2_X1 u1_u3_u5_U22 (.A2( u1_u3_u5_n122 ) , .ZN( u1_u3_u5_n136 ) , .A1( u1_u3_u5_n154 ) );
  NAND2_X1 u1_u3_u5_U23 (.A2( u1_u3_u5_n119 ) , .A1( u1_u3_u5_n120 ) , .ZN( u1_u3_u5_n159 ) );
  INV_X1 u1_u3_u5_U24 (.A( u1_u3_u5_n156 ) , .ZN( u1_u3_u5_n175 ) );
  INV_X1 u1_u3_u5_U25 (.A( u1_u3_u5_n158 ) , .ZN( u1_u3_u5_n188 ) );
  INV_X1 u1_u3_u5_U26 (.A( u1_u3_u5_n152 ) , .ZN( u1_u3_u5_n179 ) );
  INV_X1 u1_u3_u5_U27 (.A( u1_u3_u5_n140 ) , .ZN( u1_u3_u5_n182 ) );
  INV_X1 u1_u3_u5_U28 (.A( u1_u3_u5_n151 ) , .ZN( u1_u3_u5_n183 ) );
  INV_X1 u1_u3_u5_U29 (.A( u1_u3_u5_n123 ) , .ZN( u1_u3_u5_n185 ) );
  NOR2_X1 u1_u3_u5_U3 (.ZN( u1_u3_u5_n134 ) , .A1( u1_u3_u5_n183 ) , .A2( u1_u3_u5_n190 ) );
  INV_X1 u1_u3_u5_U30 (.A( u1_u3_u5_n161 ) , .ZN( u1_u3_u5_n184 ) );
  INV_X1 u1_u3_u5_U31 (.A( u1_u3_u5_n139 ) , .ZN( u1_u3_u5_n189 ) );
  INV_X1 u1_u3_u5_U32 (.A( u1_u3_u5_n157 ) , .ZN( u1_u3_u5_n190 ) );
  INV_X1 u1_u3_u5_U33 (.A( u1_u3_u5_n120 ) , .ZN( u1_u3_u5_n193 ) );
  NAND2_X1 u1_u3_u5_U34 (.ZN( u1_u3_u5_n111 ) , .A1( u1_u3_u5_n140 ) , .A2( u1_u3_u5_n155 ) );
  INV_X1 u1_u3_u5_U35 (.A( u1_u3_u5_n117 ) , .ZN( u1_u3_u5_n196 ) );
  OAI221_X1 u1_u3_u5_U36 (.A( u1_u3_u5_n116 ) , .ZN( u1_u3_u5_n117 ) , .B2( u1_u3_u5_n119 ) , .C1( u1_u3_u5_n153 ) , .C2( u1_u3_u5_n158 ) , .B1( u1_u3_u5_n172 ) );
  AOI222_X1 u1_u3_u5_U37 (.ZN( u1_u3_u5_n116 ) , .B2( u1_u3_u5_n145 ) , .C1( u1_u3_u5_n148 ) , .A2( u1_u3_u5_n174 ) , .C2( u1_u3_u5_n177 ) , .B1( u1_u3_u5_n187 ) , .A1( u1_u3_u5_n193 ) );
  INV_X1 u1_u3_u5_U38 (.A( u1_u3_u5_n115 ) , .ZN( u1_u3_u5_n187 ) );
  NOR2_X1 u1_u3_u5_U39 (.ZN( u1_u3_u5_n100 ) , .A1( u1_u3_u5_n170 ) , .A2( u1_u3_u5_n180 ) );
  INV_X1 u1_u3_u5_U4 (.A( u1_u3_u5_n138 ) , .ZN( u1_u3_u5_n191 ) );
  AOI22_X1 u1_u3_u5_U40 (.B2( u1_u3_u5_n131 ) , .A2( u1_u3_u5_n146 ) , .ZN( u1_u3_u5_n169 ) , .B1( u1_u3_u5_n174 ) , .A1( u1_u3_u5_n185 ) );
  NOR2_X1 u1_u3_u5_U41 (.A1( u1_u3_u5_n146 ) , .ZN( u1_u3_u5_n150 ) , .A2( u1_u3_u5_n173 ) );
  AOI21_X1 u1_u3_u5_U42 (.A( u1_u3_u5_n118 ) , .B2( u1_u3_u5_n145 ) , .ZN( u1_u3_u5_n168 ) , .B1( u1_u3_u5_n186 ) );
  INV_X1 u1_u3_u5_U43 (.A( u1_u3_u5_n122 ) , .ZN( u1_u3_u5_n186 ) );
  NOR2_X1 u1_u3_u5_U44 (.A1( u1_u3_u5_n146 ) , .ZN( u1_u3_u5_n152 ) , .A2( u1_u3_u5_n176 ) );
  NOR2_X1 u1_u3_u5_U45 (.A1( u1_u3_u5_n115 ) , .ZN( u1_u3_u5_n118 ) , .A2( u1_u3_u5_n153 ) );
  NOR2_X1 u1_u3_u5_U46 (.A2( u1_u3_u5_n145 ) , .ZN( u1_u3_u5_n156 ) , .A1( u1_u3_u5_n174 ) );
  NOR2_X1 u1_u3_u5_U47 (.ZN( u1_u3_u5_n121 ) , .A2( u1_u3_u5_n145 ) , .A1( u1_u3_u5_n176 ) );
  AOI22_X1 u1_u3_u5_U48 (.ZN( u1_u3_u5_n114 ) , .A2( u1_u3_u5_n137 ) , .A1( u1_u3_u5_n145 ) , .B2( u1_u3_u5_n175 ) , .B1( u1_u3_u5_n193 ) );
  OAI211_X1 u1_u3_u5_U49 (.B( u1_u3_u5_n124 ) , .A( u1_u3_u5_n125 ) , .C2( u1_u3_u5_n126 ) , .C1( u1_u3_u5_n127 ) , .ZN( u1_u3_u5_n128 ) );
  OAI21_X1 u1_u3_u5_U5 (.B2( u1_u3_u5_n136 ) , .B1( u1_u3_u5_n137 ) , .ZN( u1_u3_u5_n138 ) , .A( u1_u3_u5_n177 ) );
  NOR3_X1 u1_u3_u5_U50 (.ZN( u1_u3_u5_n127 ) , .A1( u1_u3_u5_n136 ) , .A3( u1_u3_u5_n148 ) , .A2( u1_u3_u5_n182 ) );
  OAI21_X1 u1_u3_u5_U51 (.ZN( u1_u3_u5_n124 ) , .A( u1_u3_u5_n177 ) , .B2( u1_u3_u5_n183 ) , .B1( u1_u3_u5_n189 ) );
  OAI21_X1 u1_u3_u5_U52 (.ZN( u1_u3_u5_n125 ) , .A( u1_u3_u5_n174 ) , .B2( u1_u3_u5_n185 ) , .B1( u1_u3_u5_n190 ) );
  AOI21_X1 u1_u3_u5_U53 (.A( u1_u3_u5_n153 ) , .B2( u1_u3_u5_n154 ) , .B1( u1_u3_u5_n155 ) , .ZN( u1_u3_u5_n164 ) );
  AOI21_X1 u1_u3_u5_U54 (.ZN( u1_u3_u5_n110 ) , .B1( u1_u3_u5_n122 ) , .B2( u1_u3_u5_n139 ) , .A( u1_u3_u5_n153 ) );
  INV_X1 u1_u3_u5_U55 (.A( u1_u3_u5_n153 ) , .ZN( u1_u3_u5_n176 ) );
  INV_X1 u1_u3_u5_U56 (.A( u1_u3_u5_n126 ) , .ZN( u1_u3_u5_n173 ) );
  AND2_X1 u1_u3_u5_U57 (.A2( u1_u3_u5_n104 ) , .A1( u1_u3_u5_n107 ) , .ZN( u1_u3_u5_n147 ) );
  AND2_X1 u1_u3_u5_U58 (.A2( u1_u3_u5_n104 ) , .A1( u1_u3_u5_n108 ) , .ZN( u1_u3_u5_n148 ) );
  NAND2_X1 u1_u3_u5_U59 (.A1( u1_u3_u5_n105 ) , .A2( u1_u3_u5_n106 ) , .ZN( u1_u3_u5_n158 ) );
  INV_X1 u1_u3_u5_U6 (.A( u1_u3_u5_n135 ) , .ZN( u1_u3_u5_n178 ) );
  NAND2_X1 u1_u3_u5_U60 (.A2( u1_u3_u5_n108 ) , .A1( u1_u3_u5_n109 ) , .ZN( u1_u3_u5_n139 ) );
  NAND2_X1 u1_u3_u5_U61 (.A1( u1_u3_u5_n106 ) , .A2( u1_u3_u5_n108 ) , .ZN( u1_u3_u5_n119 ) );
  NAND2_X1 u1_u3_u5_U62 (.A2( u1_u3_u5_n103 ) , .A1( u1_u3_u5_n105 ) , .ZN( u1_u3_u5_n140 ) );
  NAND2_X1 u1_u3_u5_U63 (.A2( u1_u3_u5_n104 ) , .A1( u1_u3_u5_n105 ) , .ZN( u1_u3_u5_n155 ) );
  NAND2_X1 u1_u3_u5_U64 (.A2( u1_u3_u5_n106 ) , .A1( u1_u3_u5_n107 ) , .ZN( u1_u3_u5_n122 ) );
  NAND2_X1 u1_u3_u5_U65 (.A2( u1_u3_u5_n100 ) , .A1( u1_u3_u5_n106 ) , .ZN( u1_u3_u5_n115 ) );
  NAND2_X1 u1_u3_u5_U66 (.A2( u1_u3_u5_n100 ) , .A1( u1_u3_u5_n103 ) , .ZN( u1_u3_u5_n161 ) );
  NAND2_X1 u1_u3_u5_U67 (.A1( u1_u3_u5_n105 ) , .A2( u1_u3_u5_n109 ) , .ZN( u1_u3_u5_n154 ) );
  INV_X1 u1_u3_u5_U68 (.A( u1_u3_u5_n146 ) , .ZN( u1_u3_u5_n172 ) );
  NAND2_X1 u1_u3_u5_U69 (.A1( u1_u3_u5_n103 ) , .A2( u1_u3_u5_n108 ) , .ZN( u1_u3_u5_n123 ) );
  OAI22_X1 u1_u3_u5_U7 (.B2( u1_u3_u5_n149 ) , .B1( u1_u3_u5_n150 ) , .A2( u1_u3_u5_n151 ) , .A1( u1_u3_u5_n152 ) , .ZN( u1_u3_u5_n165 ) );
  NAND2_X1 u1_u3_u5_U70 (.A2( u1_u3_u5_n103 ) , .A1( u1_u3_u5_n107 ) , .ZN( u1_u3_u5_n151 ) );
  NAND2_X1 u1_u3_u5_U71 (.A2( u1_u3_u5_n107 ) , .A1( u1_u3_u5_n109 ) , .ZN( u1_u3_u5_n120 ) );
  NAND2_X1 u1_u3_u5_U72 (.A2( u1_u3_u5_n100 ) , .A1( u1_u3_u5_n109 ) , .ZN( u1_u3_u5_n157 ) );
  AND2_X1 u1_u3_u5_U73 (.A2( u1_u3_u5_n100 ) , .A1( u1_u3_u5_n104 ) , .ZN( u1_u3_u5_n131 ) );
  INV_X1 u1_u3_u5_U74 (.A( u1_u3_u5_n102 ) , .ZN( u1_u3_u5_n195 ) );
  OAI221_X1 u1_u3_u5_U75 (.A( u1_u3_u5_n101 ) , .ZN( u1_u3_u5_n102 ) , .C2( u1_u3_u5_n115 ) , .C1( u1_u3_u5_n126 ) , .B1( u1_u3_u5_n134 ) , .B2( u1_u3_u5_n160 ) );
  OAI21_X1 u1_u3_u5_U76 (.ZN( u1_u3_u5_n101 ) , .B1( u1_u3_u5_n137 ) , .A( u1_u3_u5_n146 ) , .B2( u1_u3_u5_n147 ) );
  NOR2_X1 u1_u3_u5_U77 (.A2( u1_u3_X_34 ) , .A1( u1_u3_X_35 ) , .ZN( u1_u3_u5_n145 ) );
  NOR2_X1 u1_u3_u5_U78 (.A2( u1_u3_X_34 ) , .ZN( u1_u3_u5_n146 ) , .A1( u1_u3_u5_n171 ) );
  NOR2_X1 u1_u3_u5_U79 (.A2( u1_u3_X_31 ) , .A1( u1_u3_X_32 ) , .ZN( u1_u3_u5_n103 ) );
  NOR3_X1 u1_u3_u5_U8 (.A2( u1_u3_u5_n147 ) , .A1( u1_u3_u5_n148 ) , .ZN( u1_u3_u5_n149 ) , .A3( u1_u3_u5_n194 ) );
  NOR2_X1 u1_u3_u5_U80 (.A2( u1_u3_X_36 ) , .ZN( u1_u3_u5_n105 ) , .A1( u1_u3_u5_n180 ) );
  NOR2_X1 u1_u3_u5_U81 (.A2( u1_u3_X_33 ) , .ZN( u1_u3_u5_n108 ) , .A1( u1_u3_u5_n170 ) );
  NOR2_X1 u1_u3_u5_U82 (.A2( u1_u3_X_33 ) , .A1( u1_u3_X_36 ) , .ZN( u1_u3_u5_n107 ) );
  NOR2_X1 u1_u3_u5_U83 (.A2( u1_u3_X_31 ) , .ZN( u1_u3_u5_n104 ) , .A1( u1_u3_u5_n181 ) );
  NAND2_X1 u1_u3_u5_U84 (.A2( u1_u3_X_34 ) , .A1( u1_u3_X_35 ) , .ZN( u1_u3_u5_n153 ) );
  NAND2_X1 u1_u3_u5_U85 (.A1( u1_u3_X_34 ) , .ZN( u1_u3_u5_n126 ) , .A2( u1_u3_u5_n171 ) );
  AND2_X1 u1_u3_u5_U86 (.A1( u1_u3_X_31 ) , .A2( u1_u3_X_32 ) , .ZN( u1_u3_u5_n106 ) );
  AND2_X1 u1_u3_u5_U87 (.A1( u1_u3_X_31 ) , .ZN( u1_u3_u5_n109 ) , .A2( u1_u3_u5_n181 ) );
  INV_X1 u1_u3_u5_U88 (.A( u1_u3_X_33 ) , .ZN( u1_u3_u5_n180 ) );
  INV_X1 u1_u3_u5_U89 (.A( u1_u3_X_35 ) , .ZN( u1_u3_u5_n171 ) );
  NOR2_X1 u1_u3_u5_U9 (.ZN( u1_u3_u5_n135 ) , .A1( u1_u3_u5_n173 ) , .A2( u1_u3_u5_n176 ) );
  INV_X1 u1_u3_u5_U90 (.A( u1_u3_X_36 ) , .ZN( u1_u3_u5_n170 ) );
  INV_X1 u1_u3_u5_U91 (.A( u1_u3_X_32 ) , .ZN( u1_u3_u5_n181 ) );
  NAND4_X1 u1_u3_u5_U92 (.ZN( u1_out3_29 ) , .A4( u1_u3_u5_n129 ) , .A3( u1_u3_u5_n130 ) , .A2( u1_u3_u5_n168 ) , .A1( u1_u3_u5_n196 ) );
  AOI221_X1 u1_u3_u5_U93 (.A( u1_u3_u5_n128 ) , .ZN( u1_u3_u5_n129 ) , .C2( u1_u3_u5_n132 ) , .B2( u1_u3_u5_n159 ) , .B1( u1_u3_u5_n176 ) , .C1( u1_u3_u5_n184 ) );
  AOI222_X1 u1_u3_u5_U94 (.ZN( u1_u3_u5_n130 ) , .A2( u1_u3_u5_n146 ) , .B1( u1_u3_u5_n147 ) , .C2( u1_u3_u5_n175 ) , .B2( u1_u3_u5_n179 ) , .A1( u1_u3_u5_n188 ) , .C1( u1_u3_u5_n194 ) );
  NAND4_X1 u1_u3_u5_U95 (.ZN( u1_out3_19 ) , .A4( u1_u3_u5_n166 ) , .A3( u1_u3_u5_n167 ) , .A2( u1_u3_u5_n168 ) , .A1( u1_u3_u5_n169 ) );
  AOI22_X1 u1_u3_u5_U96 (.B2( u1_u3_u5_n145 ) , .A2( u1_u3_u5_n146 ) , .ZN( u1_u3_u5_n167 ) , .B1( u1_u3_u5_n182 ) , .A1( u1_u3_u5_n189 ) );
  NOR4_X1 u1_u3_u5_U97 (.A4( u1_u3_u5_n162 ) , .A3( u1_u3_u5_n163 ) , .A2( u1_u3_u5_n164 ) , .A1( u1_u3_u5_n165 ) , .ZN( u1_u3_u5_n166 ) );
  NAND4_X1 u1_u3_u5_U98 (.ZN( u1_out3_11 ) , .A4( u1_u3_u5_n143 ) , .A3( u1_u3_u5_n144 ) , .A2( u1_u3_u5_n169 ) , .A1( u1_u3_u5_n196 ) );
  AOI22_X1 u1_u3_u5_U99 (.A2( u1_u3_u5_n132 ) , .ZN( u1_u3_u5_n144 ) , .B2( u1_u3_u5_n145 ) , .B1( u1_u3_u5_n184 ) , .A1( u1_u3_u5_n194 ) );
  INV_X1 u1_u3_u6_U10 (.ZN( u1_u3_u6_n172 ) , .A( u1_u3_u6_n88 ) );
  OAI21_X1 u1_u3_u6_U11 (.A( u1_u3_u6_n159 ) , .B1( u1_u3_u6_n169 ) , .B2( u1_u3_u6_n173 ) , .ZN( u1_u3_u6_n90 ) );
  AOI22_X1 u1_u3_u6_U12 (.A2( u1_u3_u6_n151 ) , .B2( u1_u3_u6_n161 ) , .A1( u1_u3_u6_n167 ) , .B1( u1_u3_u6_n170 ) , .ZN( u1_u3_u6_n89 ) );
  AOI21_X1 u1_u3_u6_U13 (.ZN( u1_u3_u6_n106 ) , .A( u1_u3_u6_n142 ) , .B2( u1_u3_u6_n159 ) , .B1( u1_u3_u6_n164 ) );
  INV_X1 u1_u3_u6_U14 (.A( u1_u3_u6_n155 ) , .ZN( u1_u3_u6_n161 ) );
  INV_X1 u1_u3_u6_U15 (.A( u1_u3_u6_n128 ) , .ZN( u1_u3_u6_n164 ) );
  NAND2_X1 u1_u3_u6_U16 (.ZN( u1_u3_u6_n110 ) , .A1( u1_u3_u6_n122 ) , .A2( u1_u3_u6_n129 ) );
  NAND2_X1 u1_u3_u6_U17 (.ZN( u1_u3_u6_n124 ) , .A2( u1_u3_u6_n146 ) , .A1( u1_u3_u6_n148 ) );
  INV_X1 u1_u3_u6_U18 (.A( u1_u3_u6_n132 ) , .ZN( u1_u3_u6_n171 ) );
  AND2_X1 u1_u3_u6_U19 (.A1( u1_u3_u6_n100 ) , .ZN( u1_u3_u6_n130 ) , .A2( u1_u3_u6_n147 ) );
  INV_X1 u1_u3_u6_U20 (.A( u1_u3_u6_n127 ) , .ZN( u1_u3_u6_n173 ) );
  INV_X1 u1_u3_u6_U21 (.A( u1_u3_u6_n121 ) , .ZN( u1_u3_u6_n167 ) );
  INV_X1 u1_u3_u6_U22 (.A( u1_u3_u6_n100 ) , .ZN( u1_u3_u6_n169 ) );
  INV_X1 u1_u3_u6_U23 (.A( u1_u3_u6_n123 ) , .ZN( u1_u3_u6_n170 ) );
  INV_X1 u1_u3_u6_U24 (.A( u1_u3_u6_n113 ) , .ZN( u1_u3_u6_n168 ) );
  AND2_X1 u1_u3_u6_U25 (.A1( u1_u3_u6_n107 ) , .A2( u1_u3_u6_n119 ) , .ZN( u1_u3_u6_n133 ) );
  AND2_X1 u1_u3_u6_U26 (.A2( u1_u3_u6_n121 ) , .A1( u1_u3_u6_n122 ) , .ZN( u1_u3_u6_n131 ) );
  AND3_X1 u1_u3_u6_U27 (.ZN( u1_u3_u6_n120 ) , .A2( u1_u3_u6_n127 ) , .A1( u1_u3_u6_n132 ) , .A3( u1_u3_u6_n145 ) );
  INV_X1 u1_u3_u6_U28 (.A( u1_u3_u6_n146 ) , .ZN( u1_u3_u6_n163 ) );
  AOI222_X1 u1_u3_u6_U29 (.ZN( u1_u3_u6_n114 ) , .A1( u1_u3_u6_n118 ) , .A2( u1_u3_u6_n126 ) , .B2( u1_u3_u6_n151 ) , .C2( u1_u3_u6_n159 ) , .C1( u1_u3_u6_n168 ) , .B1( u1_u3_u6_n169 ) );
  INV_X1 u1_u3_u6_U3 (.A( u1_u3_u6_n110 ) , .ZN( u1_u3_u6_n166 ) );
  NOR2_X1 u1_u3_u6_U30 (.A1( u1_u3_u6_n162 ) , .A2( u1_u3_u6_n165 ) , .ZN( u1_u3_u6_n98 ) );
  NAND2_X1 u1_u3_u6_U31 (.A1( u1_u3_u6_n144 ) , .ZN( u1_u3_u6_n151 ) , .A2( u1_u3_u6_n158 ) );
  NAND2_X1 u1_u3_u6_U32 (.ZN( u1_u3_u6_n132 ) , .A1( u1_u3_u6_n91 ) , .A2( u1_u3_u6_n97 ) );
  AOI22_X1 u1_u3_u6_U33 (.B2( u1_u3_u6_n110 ) , .B1( u1_u3_u6_n111 ) , .A1( u1_u3_u6_n112 ) , .ZN( u1_u3_u6_n115 ) , .A2( u1_u3_u6_n161 ) );
  NAND4_X1 u1_u3_u6_U34 (.A3( u1_u3_u6_n109 ) , .ZN( u1_u3_u6_n112 ) , .A4( u1_u3_u6_n132 ) , .A2( u1_u3_u6_n147 ) , .A1( u1_u3_u6_n166 ) );
  NOR2_X1 u1_u3_u6_U35 (.ZN( u1_u3_u6_n109 ) , .A1( u1_u3_u6_n170 ) , .A2( u1_u3_u6_n173 ) );
  NOR2_X1 u1_u3_u6_U36 (.A2( u1_u3_u6_n126 ) , .ZN( u1_u3_u6_n155 ) , .A1( u1_u3_u6_n160 ) );
  NAND2_X1 u1_u3_u6_U37 (.ZN( u1_u3_u6_n146 ) , .A2( u1_u3_u6_n94 ) , .A1( u1_u3_u6_n99 ) );
  AOI21_X1 u1_u3_u6_U38 (.A( u1_u3_u6_n144 ) , .B2( u1_u3_u6_n145 ) , .B1( u1_u3_u6_n146 ) , .ZN( u1_u3_u6_n150 ) );
  AOI211_X1 u1_u3_u6_U39 (.B( u1_u3_u6_n134 ) , .A( u1_u3_u6_n135 ) , .C1( u1_u3_u6_n136 ) , .ZN( u1_u3_u6_n137 ) , .C2( u1_u3_u6_n151 ) );
  INV_X1 u1_u3_u6_U4 (.A( u1_u3_u6_n142 ) , .ZN( u1_u3_u6_n174 ) );
  AOI21_X1 u1_u3_u6_U40 (.B2( u1_u3_u6_n132 ) , .B1( u1_u3_u6_n133 ) , .ZN( u1_u3_u6_n134 ) , .A( u1_u3_u6_n158 ) );
  NAND4_X1 u1_u3_u6_U41 (.A4( u1_u3_u6_n127 ) , .A3( u1_u3_u6_n128 ) , .A2( u1_u3_u6_n129 ) , .A1( u1_u3_u6_n130 ) , .ZN( u1_u3_u6_n136 ) );
  AOI21_X1 u1_u3_u6_U42 (.B1( u1_u3_u6_n131 ) , .ZN( u1_u3_u6_n135 ) , .A( u1_u3_u6_n144 ) , .B2( u1_u3_u6_n146 ) );
  INV_X1 u1_u3_u6_U43 (.A( u1_u3_u6_n111 ) , .ZN( u1_u3_u6_n158 ) );
  NAND2_X1 u1_u3_u6_U44 (.ZN( u1_u3_u6_n127 ) , .A1( u1_u3_u6_n91 ) , .A2( u1_u3_u6_n92 ) );
  NAND2_X1 u1_u3_u6_U45 (.ZN( u1_u3_u6_n129 ) , .A2( u1_u3_u6_n95 ) , .A1( u1_u3_u6_n96 ) );
  INV_X1 u1_u3_u6_U46 (.A( u1_u3_u6_n144 ) , .ZN( u1_u3_u6_n159 ) );
  NAND2_X1 u1_u3_u6_U47 (.ZN( u1_u3_u6_n145 ) , .A2( u1_u3_u6_n97 ) , .A1( u1_u3_u6_n98 ) );
  NAND2_X1 u1_u3_u6_U48 (.ZN( u1_u3_u6_n148 ) , .A2( u1_u3_u6_n92 ) , .A1( u1_u3_u6_n94 ) );
  NAND2_X1 u1_u3_u6_U49 (.ZN( u1_u3_u6_n108 ) , .A2( u1_u3_u6_n139 ) , .A1( u1_u3_u6_n144 ) );
  NAND2_X1 u1_u3_u6_U5 (.A2( u1_u3_u6_n143 ) , .ZN( u1_u3_u6_n152 ) , .A1( u1_u3_u6_n166 ) );
  NAND2_X1 u1_u3_u6_U50 (.ZN( u1_u3_u6_n121 ) , .A2( u1_u3_u6_n95 ) , .A1( u1_u3_u6_n97 ) );
  NAND2_X1 u1_u3_u6_U51 (.ZN( u1_u3_u6_n107 ) , .A2( u1_u3_u6_n92 ) , .A1( u1_u3_u6_n95 ) );
  AND2_X1 u1_u3_u6_U52 (.ZN( u1_u3_u6_n118 ) , .A2( u1_u3_u6_n91 ) , .A1( u1_u3_u6_n99 ) );
  NAND2_X1 u1_u3_u6_U53 (.ZN( u1_u3_u6_n147 ) , .A2( u1_u3_u6_n98 ) , .A1( u1_u3_u6_n99 ) );
  NAND2_X1 u1_u3_u6_U54 (.ZN( u1_u3_u6_n128 ) , .A1( u1_u3_u6_n94 ) , .A2( u1_u3_u6_n96 ) );
  NAND2_X1 u1_u3_u6_U55 (.ZN( u1_u3_u6_n119 ) , .A2( u1_u3_u6_n95 ) , .A1( u1_u3_u6_n99 ) );
  NAND2_X1 u1_u3_u6_U56 (.ZN( u1_u3_u6_n123 ) , .A2( u1_u3_u6_n91 ) , .A1( u1_u3_u6_n96 ) );
  NAND2_X1 u1_u3_u6_U57 (.ZN( u1_u3_u6_n100 ) , .A2( u1_u3_u6_n92 ) , .A1( u1_u3_u6_n98 ) );
  NAND2_X1 u1_u3_u6_U58 (.ZN( u1_u3_u6_n122 ) , .A1( u1_u3_u6_n94 ) , .A2( u1_u3_u6_n97 ) );
  INV_X1 u1_u3_u6_U59 (.A( u1_u3_u6_n139 ) , .ZN( u1_u3_u6_n160 ) );
  AOI22_X1 u1_u3_u6_U6 (.B2( u1_u3_u6_n101 ) , .A1( u1_u3_u6_n102 ) , .ZN( u1_u3_u6_n103 ) , .B1( u1_u3_u6_n160 ) , .A2( u1_u3_u6_n161 ) );
  NAND2_X1 u1_u3_u6_U60 (.ZN( u1_u3_u6_n113 ) , .A1( u1_u3_u6_n96 ) , .A2( u1_u3_u6_n98 ) );
  NOR2_X1 u1_u3_u6_U61 (.A2( u1_u3_X_40 ) , .A1( u1_u3_X_41 ) , .ZN( u1_u3_u6_n126 ) );
  NOR2_X1 u1_u3_u6_U62 (.A2( u1_u3_X_39 ) , .A1( u1_u3_X_42 ) , .ZN( u1_u3_u6_n92 ) );
  NOR2_X1 u1_u3_u6_U63 (.A2( u1_u3_X_39 ) , .A1( u1_u3_u6_n156 ) , .ZN( u1_u3_u6_n97 ) );
  NOR2_X1 u1_u3_u6_U64 (.A2( u1_u3_X_38 ) , .A1( u1_u3_u6_n165 ) , .ZN( u1_u3_u6_n95 ) );
  NOR2_X1 u1_u3_u6_U65 (.A2( u1_u3_X_41 ) , .ZN( u1_u3_u6_n111 ) , .A1( u1_u3_u6_n157 ) );
  NOR2_X1 u1_u3_u6_U66 (.A2( u1_u3_X_37 ) , .A1( u1_u3_u6_n162 ) , .ZN( u1_u3_u6_n94 ) );
  NOR2_X1 u1_u3_u6_U67 (.A2( u1_u3_X_37 ) , .A1( u1_u3_X_38 ) , .ZN( u1_u3_u6_n91 ) );
  NAND2_X1 u1_u3_u6_U68 (.A1( u1_u3_X_41 ) , .ZN( u1_u3_u6_n144 ) , .A2( u1_u3_u6_n157 ) );
  NAND2_X1 u1_u3_u6_U69 (.A2( u1_u3_X_40 ) , .A1( u1_u3_X_41 ) , .ZN( u1_u3_u6_n139 ) );
  NOR2_X1 u1_u3_u6_U7 (.A1( u1_u3_u6_n118 ) , .ZN( u1_u3_u6_n143 ) , .A2( u1_u3_u6_n168 ) );
  AND2_X1 u1_u3_u6_U70 (.A1( u1_u3_X_39 ) , .A2( u1_u3_u6_n156 ) , .ZN( u1_u3_u6_n96 ) );
  AND2_X1 u1_u3_u6_U71 (.A1( u1_u3_X_39 ) , .A2( u1_u3_X_42 ) , .ZN( u1_u3_u6_n99 ) );
  INV_X1 u1_u3_u6_U72 (.A( u1_u3_X_40 ) , .ZN( u1_u3_u6_n157 ) );
  INV_X1 u1_u3_u6_U73 (.A( u1_u3_X_37 ) , .ZN( u1_u3_u6_n165 ) );
  INV_X1 u1_u3_u6_U74 (.A( u1_u3_X_38 ) , .ZN( u1_u3_u6_n162 ) );
  INV_X1 u1_u3_u6_U75 (.A( u1_u3_X_42 ) , .ZN( u1_u3_u6_n156 ) );
  NAND4_X1 u1_u3_u6_U76 (.ZN( u1_out3_32 ) , .A4( u1_u3_u6_n103 ) , .A3( u1_u3_u6_n104 ) , .A2( u1_u3_u6_n105 ) , .A1( u1_u3_u6_n106 ) );
  AOI22_X1 u1_u3_u6_U77 (.ZN( u1_u3_u6_n105 ) , .A2( u1_u3_u6_n108 ) , .A1( u1_u3_u6_n118 ) , .B2( u1_u3_u6_n126 ) , .B1( u1_u3_u6_n171 ) );
  AOI22_X1 u1_u3_u6_U78 (.ZN( u1_u3_u6_n104 ) , .A1( u1_u3_u6_n111 ) , .B1( u1_u3_u6_n124 ) , .B2( u1_u3_u6_n151 ) , .A2( u1_u3_u6_n93 ) );
  NAND4_X1 u1_u3_u6_U79 (.ZN( u1_out3_12 ) , .A4( u1_u3_u6_n114 ) , .A3( u1_u3_u6_n115 ) , .A2( u1_u3_u6_n116 ) , .A1( u1_u3_u6_n117 ) );
  AOI21_X1 u1_u3_u6_U8 (.B1( u1_u3_u6_n107 ) , .B2( u1_u3_u6_n132 ) , .A( u1_u3_u6_n158 ) , .ZN( u1_u3_u6_n88 ) );
  OAI22_X1 u1_u3_u6_U80 (.B2( u1_u3_u6_n111 ) , .ZN( u1_u3_u6_n116 ) , .B1( u1_u3_u6_n126 ) , .A2( u1_u3_u6_n164 ) , .A1( u1_u3_u6_n167 ) );
  OAI21_X1 u1_u3_u6_U81 (.A( u1_u3_u6_n108 ) , .ZN( u1_u3_u6_n117 ) , .B2( u1_u3_u6_n141 ) , .B1( u1_u3_u6_n163 ) );
  OAI211_X1 u1_u3_u6_U82 (.ZN( u1_out3_22 ) , .B( u1_u3_u6_n137 ) , .A( u1_u3_u6_n138 ) , .C2( u1_u3_u6_n139 ) , .C1( u1_u3_u6_n140 ) );
  AOI22_X1 u1_u3_u6_U83 (.B1( u1_u3_u6_n124 ) , .A2( u1_u3_u6_n125 ) , .A1( u1_u3_u6_n126 ) , .ZN( u1_u3_u6_n138 ) , .B2( u1_u3_u6_n161 ) );
  AND4_X1 u1_u3_u6_U84 (.A3( u1_u3_u6_n119 ) , .A1( u1_u3_u6_n120 ) , .A4( u1_u3_u6_n129 ) , .ZN( u1_u3_u6_n140 ) , .A2( u1_u3_u6_n143 ) );
  OAI211_X1 u1_u3_u6_U85 (.ZN( u1_out3_7 ) , .B( u1_u3_u6_n153 ) , .C2( u1_u3_u6_n154 ) , .C1( u1_u3_u6_n155 ) , .A( u1_u3_u6_n174 ) );
  NOR3_X1 u1_u3_u6_U86 (.A1( u1_u3_u6_n141 ) , .ZN( u1_u3_u6_n154 ) , .A3( u1_u3_u6_n164 ) , .A2( u1_u3_u6_n171 ) );
  AOI211_X1 u1_u3_u6_U87 (.B( u1_u3_u6_n149 ) , .A( u1_u3_u6_n150 ) , .C2( u1_u3_u6_n151 ) , .C1( u1_u3_u6_n152 ) , .ZN( u1_u3_u6_n153 ) );
  NAND3_X1 u1_u3_u6_U88 (.A2( u1_u3_u6_n123 ) , .ZN( u1_u3_u6_n125 ) , .A1( u1_u3_u6_n130 ) , .A3( u1_u3_u6_n131 ) );
  NAND3_X1 u1_u3_u6_U89 (.A3( u1_u3_u6_n133 ) , .ZN( u1_u3_u6_n141 ) , .A1( u1_u3_u6_n145 ) , .A2( u1_u3_u6_n148 ) );
  AOI21_X1 u1_u3_u6_U9 (.B2( u1_u3_u6_n147 ) , .B1( u1_u3_u6_n148 ) , .ZN( u1_u3_u6_n149 ) , .A( u1_u3_u6_n158 ) );
  NAND3_X1 u1_u3_u6_U90 (.ZN( u1_u3_u6_n101 ) , .A3( u1_u3_u6_n107 ) , .A2( u1_u3_u6_n121 ) , .A1( u1_u3_u6_n127 ) );
  NAND3_X1 u1_u3_u6_U91 (.ZN( u1_u3_u6_n102 ) , .A3( u1_u3_u6_n130 ) , .A2( u1_u3_u6_n145 ) , .A1( u1_u3_u6_n166 ) );
  NAND3_X1 u1_u3_u6_U92 (.A3( u1_u3_u6_n113 ) , .A1( u1_u3_u6_n119 ) , .A2( u1_u3_u6_n123 ) , .ZN( u1_u3_u6_n93 ) );
  NAND3_X1 u1_u3_u6_U93 (.ZN( u1_u3_u6_n142 ) , .A2( u1_u3_u6_n172 ) , .A3( u1_u3_u6_n89 ) , .A1( u1_u3_u6_n90 ) );
  XOR2_X1 u1_u4_U10 (.B( u1_K5_45 ) , .A( u1_R3_30 ) , .Z( u1_u4_X_45 ) );
  XOR2_X1 u1_u4_U11 (.B( u1_K5_44 ) , .A( u1_R3_29 ) , .Z( u1_u4_X_44 ) );
  XOR2_X1 u1_u4_U12 (.B( u1_K5_43 ) , .A( u1_R3_28 ) , .Z( u1_u4_X_43 ) );
  XOR2_X1 u1_u4_U26 (.B( u1_K5_30 ) , .A( u1_R3_21 ) , .Z( u1_u4_X_30 ) );
  XOR2_X1 u1_u4_U28 (.B( u1_K5_29 ) , .A( u1_R3_20 ) , .Z( u1_u4_X_29 ) );
  XOR2_X1 u1_u4_U29 (.B( u1_K5_28 ) , .A( u1_R3_19 ) , .Z( u1_u4_X_28 ) );
  XOR2_X1 u1_u4_U30 (.B( u1_K5_27 ) , .A( u1_R3_18 ) , .Z( u1_u4_X_27 ) );
  XOR2_X1 u1_u4_U31 (.B( u1_K5_26 ) , .A( u1_R3_17 ) , .Z( u1_u4_X_26 ) );
  XOR2_X1 u1_u4_U32 (.B( u1_K5_25 ) , .A( u1_R3_16 ) , .Z( u1_u4_X_25 ) );
  XOR2_X1 u1_u4_U7 (.B( u1_K5_48 ) , .A( u1_R3_1 ) , .Z( u1_u4_X_48 ) );
  XOR2_X1 u1_u4_U8 (.B( u1_K5_47 ) , .A( u1_R3_32 ) , .Z( u1_u4_X_47 ) );
  XOR2_X1 u1_u4_U9 (.B( u1_K5_46 ) , .A( u1_R3_31 ) , .Z( u1_u4_X_46 ) );
  OAI22_X1 u1_u4_u4_U10 (.B2( u1_u4_u4_n135 ) , .ZN( u1_u4_u4_n137 ) , .B1( u1_u4_u4_n153 ) , .A1( u1_u4_u4_n155 ) , .A2( u1_u4_u4_n171 ) );
  AND3_X1 u1_u4_u4_U11 (.A2( u1_u4_u4_n134 ) , .ZN( u1_u4_u4_n135 ) , .A3( u1_u4_u4_n145 ) , .A1( u1_u4_u4_n157 ) );
  NAND2_X1 u1_u4_u4_U12 (.ZN( u1_u4_u4_n132 ) , .A2( u1_u4_u4_n170 ) , .A1( u1_u4_u4_n173 ) );
  AOI21_X1 u1_u4_u4_U13 (.B2( u1_u4_u4_n160 ) , .B1( u1_u4_u4_n161 ) , .ZN( u1_u4_u4_n162 ) , .A( u1_u4_u4_n170 ) );
  AOI21_X1 u1_u4_u4_U14 (.ZN( u1_u4_u4_n107 ) , .B2( u1_u4_u4_n143 ) , .A( u1_u4_u4_n174 ) , .B1( u1_u4_u4_n184 ) );
  AOI21_X1 u1_u4_u4_U15 (.B2( u1_u4_u4_n158 ) , .B1( u1_u4_u4_n159 ) , .ZN( u1_u4_u4_n163 ) , .A( u1_u4_u4_n174 ) );
  AOI21_X1 u1_u4_u4_U16 (.A( u1_u4_u4_n153 ) , .B2( u1_u4_u4_n154 ) , .B1( u1_u4_u4_n155 ) , .ZN( u1_u4_u4_n165 ) );
  AOI21_X1 u1_u4_u4_U17 (.A( u1_u4_u4_n156 ) , .B2( u1_u4_u4_n157 ) , .ZN( u1_u4_u4_n164 ) , .B1( u1_u4_u4_n184 ) );
  INV_X1 u1_u4_u4_U18 (.A( u1_u4_u4_n138 ) , .ZN( u1_u4_u4_n170 ) );
  AND2_X1 u1_u4_u4_U19 (.A2( u1_u4_u4_n120 ) , .ZN( u1_u4_u4_n155 ) , .A1( u1_u4_u4_n160 ) );
  INV_X1 u1_u4_u4_U20 (.A( u1_u4_u4_n156 ) , .ZN( u1_u4_u4_n175 ) );
  NAND2_X1 u1_u4_u4_U21 (.A2( u1_u4_u4_n118 ) , .ZN( u1_u4_u4_n131 ) , .A1( u1_u4_u4_n147 ) );
  NAND2_X1 u1_u4_u4_U22 (.A1( u1_u4_u4_n119 ) , .A2( u1_u4_u4_n120 ) , .ZN( u1_u4_u4_n130 ) );
  NAND2_X1 u1_u4_u4_U23 (.ZN( u1_u4_u4_n117 ) , .A2( u1_u4_u4_n118 ) , .A1( u1_u4_u4_n148 ) );
  NAND2_X1 u1_u4_u4_U24 (.ZN( u1_u4_u4_n129 ) , .A1( u1_u4_u4_n134 ) , .A2( u1_u4_u4_n148 ) );
  AND3_X1 u1_u4_u4_U25 (.A1( u1_u4_u4_n119 ) , .A2( u1_u4_u4_n143 ) , .A3( u1_u4_u4_n154 ) , .ZN( u1_u4_u4_n161 ) );
  AND2_X1 u1_u4_u4_U26 (.A1( u1_u4_u4_n145 ) , .A2( u1_u4_u4_n147 ) , .ZN( u1_u4_u4_n159 ) );
  OR3_X1 u1_u4_u4_U27 (.A3( u1_u4_u4_n114 ) , .A2( u1_u4_u4_n115 ) , .A1( u1_u4_u4_n116 ) , .ZN( u1_u4_u4_n136 ) );
  AOI21_X1 u1_u4_u4_U28 (.A( u1_u4_u4_n113 ) , .ZN( u1_u4_u4_n116 ) , .B2( u1_u4_u4_n173 ) , .B1( u1_u4_u4_n174 ) );
  AOI21_X1 u1_u4_u4_U29 (.ZN( u1_u4_u4_n115 ) , .B2( u1_u4_u4_n145 ) , .B1( u1_u4_u4_n146 ) , .A( u1_u4_u4_n156 ) );
  NOR2_X1 u1_u4_u4_U3 (.ZN( u1_u4_u4_n121 ) , .A1( u1_u4_u4_n181 ) , .A2( u1_u4_u4_n182 ) );
  OAI22_X1 u1_u4_u4_U30 (.ZN( u1_u4_u4_n114 ) , .A2( u1_u4_u4_n121 ) , .B1( u1_u4_u4_n160 ) , .B2( u1_u4_u4_n170 ) , .A1( u1_u4_u4_n171 ) );
  INV_X1 u1_u4_u4_U31 (.A( u1_u4_u4_n158 ) , .ZN( u1_u4_u4_n182 ) );
  INV_X1 u1_u4_u4_U32 (.ZN( u1_u4_u4_n181 ) , .A( u1_u4_u4_n96 ) );
  INV_X1 u1_u4_u4_U33 (.A( u1_u4_u4_n144 ) , .ZN( u1_u4_u4_n179 ) );
  INV_X1 u1_u4_u4_U34 (.A( u1_u4_u4_n157 ) , .ZN( u1_u4_u4_n178 ) );
  NAND2_X1 u1_u4_u4_U35 (.A2( u1_u4_u4_n154 ) , .A1( u1_u4_u4_n96 ) , .ZN( u1_u4_u4_n97 ) );
  INV_X1 u1_u4_u4_U36 (.ZN( u1_u4_u4_n186 ) , .A( u1_u4_u4_n95 ) );
  OAI221_X1 u1_u4_u4_U37 (.C1( u1_u4_u4_n134 ) , .B1( u1_u4_u4_n158 ) , .B2( u1_u4_u4_n171 ) , .C2( u1_u4_u4_n173 ) , .A( u1_u4_u4_n94 ) , .ZN( u1_u4_u4_n95 ) );
  AOI222_X1 u1_u4_u4_U38 (.B2( u1_u4_u4_n132 ) , .A1( u1_u4_u4_n138 ) , .C2( u1_u4_u4_n175 ) , .A2( u1_u4_u4_n179 ) , .C1( u1_u4_u4_n181 ) , .B1( u1_u4_u4_n185 ) , .ZN( u1_u4_u4_n94 ) );
  INV_X1 u1_u4_u4_U39 (.A( u1_u4_u4_n113 ) , .ZN( u1_u4_u4_n185 ) );
  INV_X1 u1_u4_u4_U4 (.A( u1_u4_u4_n117 ) , .ZN( u1_u4_u4_n184 ) );
  INV_X1 u1_u4_u4_U40 (.A( u1_u4_u4_n143 ) , .ZN( u1_u4_u4_n183 ) );
  NOR2_X1 u1_u4_u4_U41 (.ZN( u1_u4_u4_n138 ) , .A1( u1_u4_u4_n168 ) , .A2( u1_u4_u4_n169 ) );
  NOR2_X1 u1_u4_u4_U42 (.A1( u1_u4_u4_n150 ) , .A2( u1_u4_u4_n152 ) , .ZN( u1_u4_u4_n153 ) );
  NOR2_X1 u1_u4_u4_U43 (.A2( u1_u4_u4_n128 ) , .A1( u1_u4_u4_n138 ) , .ZN( u1_u4_u4_n156 ) );
  AOI22_X1 u1_u4_u4_U44 (.B2( u1_u4_u4_n122 ) , .A1( u1_u4_u4_n123 ) , .ZN( u1_u4_u4_n124 ) , .B1( u1_u4_u4_n128 ) , .A2( u1_u4_u4_n172 ) );
  INV_X1 u1_u4_u4_U45 (.A( u1_u4_u4_n153 ) , .ZN( u1_u4_u4_n172 ) );
  NAND2_X1 u1_u4_u4_U46 (.A2( u1_u4_u4_n120 ) , .ZN( u1_u4_u4_n123 ) , .A1( u1_u4_u4_n161 ) );
  AOI22_X1 u1_u4_u4_U47 (.B2( u1_u4_u4_n132 ) , .A2( u1_u4_u4_n133 ) , .ZN( u1_u4_u4_n140 ) , .A1( u1_u4_u4_n150 ) , .B1( u1_u4_u4_n179 ) );
  NAND2_X1 u1_u4_u4_U48 (.ZN( u1_u4_u4_n133 ) , .A2( u1_u4_u4_n146 ) , .A1( u1_u4_u4_n154 ) );
  NAND2_X1 u1_u4_u4_U49 (.A1( u1_u4_u4_n103 ) , .ZN( u1_u4_u4_n154 ) , .A2( u1_u4_u4_n98 ) );
  NOR4_X1 u1_u4_u4_U5 (.A4( u1_u4_u4_n106 ) , .A3( u1_u4_u4_n107 ) , .A2( u1_u4_u4_n108 ) , .A1( u1_u4_u4_n109 ) , .ZN( u1_u4_u4_n110 ) );
  NAND2_X1 u1_u4_u4_U50 (.A1( u1_u4_u4_n101 ) , .ZN( u1_u4_u4_n158 ) , .A2( u1_u4_u4_n99 ) );
  AOI21_X1 u1_u4_u4_U51 (.ZN( u1_u4_u4_n127 ) , .A( u1_u4_u4_n136 ) , .B2( u1_u4_u4_n150 ) , .B1( u1_u4_u4_n180 ) );
  INV_X1 u1_u4_u4_U52 (.A( u1_u4_u4_n160 ) , .ZN( u1_u4_u4_n180 ) );
  NAND2_X1 u1_u4_u4_U53 (.A2( u1_u4_u4_n104 ) , .A1( u1_u4_u4_n105 ) , .ZN( u1_u4_u4_n146 ) );
  NAND2_X1 u1_u4_u4_U54 (.A2( u1_u4_u4_n101 ) , .A1( u1_u4_u4_n102 ) , .ZN( u1_u4_u4_n160 ) );
  NAND2_X1 u1_u4_u4_U55 (.ZN( u1_u4_u4_n134 ) , .A1( u1_u4_u4_n98 ) , .A2( u1_u4_u4_n99 ) );
  NAND2_X1 u1_u4_u4_U56 (.A1( u1_u4_u4_n103 ) , .A2( u1_u4_u4_n104 ) , .ZN( u1_u4_u4_n143 ) );
  NAND2_X1 u1_u4_u4_U57 (.A2( u1_u4_u4_n105 ) , .ZN( u1_u4_u4_n145 ) , .A1( u1_u4_u4_n98 ) );
  NAND2_X1 u1_u4_u4_U58 (.A1( u1_u4_u4_n100 ) , .A2( u1_u4_u4_n105 ) , .ZN( u1_u4_u4_n120 ) );
  NAND2_X1 u1_u4_u4_U59 (.A1( u1_u4_u4_n102 ) , .A2( u1_u4_u4_n104 ) , .ZN( u1_u4_u4_n148 ) );
  AOI21_X1 u1_u4_u4_U6 (.ZN( u1_u4_u4_n106 ) , .B2( u1_u4_u4_n146 ) , .B1( u1_u4_u4_n158 ) , .A( u1_u4_u4_n170 ) );
  NAND2_X1 u1_u4_u4_U60 (.A2( u1_u4_u4_n100 ) , .A1( u1_u4_u4_n103 ) , .ZN( u1_u4_u4_n157 ) );
  INV_X1 u1_u4_u4_U61 (.A( u1_u4_u4_n150 ) , .ZN( u1_u4_u4_n173 ) );
  INV_X1 u1_u4_u4_U62 (.A( u1_u4_u4_n152 ) , .ZN( u1_u4_u4_n171 ) );
  NAND2_X1 u1_u4_u4_U63 (.A1( u1_u4_u4_n100 ) , .ZN( u1_u4_u4_n118 ) , .A2( u1_u4_u4_n99 ) );
  NAND2_X1 u1_u4_u4_U64 (.A2( u1_u4_u4_n100 ) , .A1( u1_u4_u4_n102 ) , .ZN( u1_u4_u4_n144 ) );
  NAND2_X1 u1_u4_u4_U65 (.A2( u1_u4_u4_n101 ) , .A1( u1_u4_u4_n105 ) , .ZN( u1_u4_u4_n96 ) );
  INV_X1 u1_u4_u4_U66 (.A( u1_u4_u4_n128 ) , .ZN( u1_u4_u4_n174 ) );
  NAND2_X1 u1_u4_u4_U67 (.A2( u1_u4_u4_n102 ) , .ZN( u1_u4_u4_n119 ) , .A1( u1_u4_u4_n98 ) );
  NAND2_X1 u1_u4_u4_U68 (.A2( u1_u4_u4_n101 ) , .A1( u1_u4_u4_n103 ) , .ZN( u1_u4_u4_n147 ) );
  NAND2_X1 u1_u4_u4_U69 (.A2( u1_u4_u4_n104 ) , .ZN( u1_u4_u4_n113 ) , .A1( u1_u4_u4_n99 ) );
  AOI21_X1 u1_u4_u4_U7 (.ZN( u1_u4_u4_n108 ) , .B2( u1_u4_u4_n134 ) , .B1( u1_u4_u4_n155 ) , .A( u1_u4_u4_n156 ) );
  NOR2_X1 u1_u4_u4_U70 (.A2( u1_u4_X_28 ) , .ZN( u1_u4_u4_n150 ) , .A1( u1_u4_u4_n168 ) );
  NOR2_X1 u1_u4_u4_U71 (.A2( u1_u4_X_29 ) , .ZN( u1_u4_u4_n152 ) , .A1( u1_u4_u4_n169 ) );
  NOR2_X1 u1_u4_u4_U72 (.A2( u1_u4_X_30 ) , .ZN( u1_u4_u4_n105 ) , .A1( u1_u4_u4_n176 ) );
  NOR2_X1 u1_u4_u4_U73 (.A2( u1_u4_X_26 ) , .ZN( u1_u4_u4_n100 ) , .A1( u1_u4_u4_n177 ) );
  NOR2_X1 u1_u4_u4_U74 (.A2( u1_u4_X_28 ) , .A1( u1_u4_X_29 ) , .ZN( u1_u4_u4_n128 ) );
  NOR2_X1 u1_u4_u4_U75 (.A2( u1_u4_X_27 ) , .A1( u1_u4_X_30 ) , .ZN( u1_u4_u4_n102 ) );
  NOR2_X1 u1_u4_u4_U76 (.A2( u1_u4_X_25 ) , .A1( u1_u4_X_26 ) , .ZN( u1_u4_u4_n98 ) );
  AND2_X1 u1_u4_u4_U77 (.A2( u1_u4_X_25 ) , .A1( u1_u4_X_26 ) , .ZN( u1_u4_u4_n104 ) );
  AND2_X1 u1_u4_u4_U78 (.A1( u1_u4_X_30 ) , .A2( u1_u4_u4_n176 ) , .ZN( u1_u4_u4_n99 ) );
  AND2_X1 u1_u4_u4_U79 (.A1( u1_u4_X_26 ) , .ZN( u1_u4_u4_n101 ) , .A2( u1_u4_u4_n177 ) );
  AOI21_X1 u1_u4_u4_U8 (.ZN( u1_u4_u4_n109 ) , .A( u1_u4_u4_n153 ) , .B1( u1_u4_u4_n159 ) , .B2( u1_u4_u4_n184 ) );
  AND2_X1 u1_u4_u4_U80 (.A1( u1_u4_X_27 ) , .A2( u1_u4_X_30 ) , .ZN( u1_u4_u4_n103 ) );
  INV_X1 u1_u4_u4_U81 (.A( u1_u4_X_28 ) , .ZN( u1_u4_u4_n169 ) );
  INV_X1 u1_u4_u4_U82 (.A( u1_u4_X_29 ) , .ZN( u1_u4_u4_n168 ) );
  INV_X1 u1_u4_u4_U83 (.A( u1_u4_X_25 ) , .ZN( u1_u4_u4_n177 ) );
  INV_X1 u1_u4_u4_U84 (.A( u1_u4_X_27 ) , .ZN( u1_u4_u4_n176 ) );
  NAND4_X1 u1_u4_u4_U85 (.ZN( u1_out4_25 ) , .A4( u1_u4_u4_n139 ) , .A3( u1_u4_u4_n140 ) , .A2( u1_u4_u4_n141 ) , .A1( u1_u4_u4_n142 ) );
  OAI21_X1 u1_u4_u4_U86 (.B2( u1_u4_u4_n131 ) , .ZN( u1_u4_u4_n141 ) , .A( u1_u4_u4_n175 ) , .B1( u1_u4_u4_n183 ) );
  OAI21_X1 u1_u4_u4_U87 (.A( u1_u4_u4_n128 ) , .B2( u1_u4_u4_n129 ) , .B1( u1_u4_u4_n130 ) , .ZN( u1_u4_u4_n142 ) );
  NAND4_X1 u1_u4_u4_U88 (.ZN( u1_out4_14 ) , .A4( u1_u4_u4_n124 ) , .A3( u1_u4_u4_n125 ) , .A2( u1_u4_u4_n126 ) , .A1( u1_u4_u4_n127 ) );
  AOI22_X1 u1_u4_u4_U89 (.B2( u1_u4_u4_n117 ) , .ZN( u1_u4_u4_n126 ) , .A1( u1_u4_u4_n129 ) , .B1( u1_u4_u4_n152 ) , .A2( u1_u4_u4_n175 ) );
  AOI211_X1 u1_u4_u4_U9 (.B( u1_u4_u4_n136 ) , .A( u1_u4_u4_n137 ) , .C2( u1_u4_u4_n138 ) , .ZN( u1_u4_u4_n139 ) , .C1( u1_u4_u4_n182 ) );
  AOI22_X1 u1_u4_u4_U90 (.ZN( u1_u4_u4_n125 ) , .B2( u1_u4_u4_n131 ) , .A2( u1_u4_u4_n132 ) , .B1( u1_u4_u4_n138 ) , .A1( u1_u4_u4_n178 ) );
  NAND4_X1 u1_u4_u4_U91 (.ZN( u1_out4_8 ) , .A4( u1_u4_u4_n110 ) , .A3( u1_u4_u4_n111 ) , .A2( u1_u4_u4_n112 ) , .A1( u1_u4_u4_n186 ) );
  NAND2_X1 u1_u4_u4_U92 (.ZN( u1_u4_u4_n112 ) , .A2( u1_u4_u4_n130 ) , .A1( u1_u4_u4_n150 ) );
  AOI22_X1 u1_u4_u4_U93 (.ZN( u1_u4_u4_n111 ) , .B2( u1_u4_u4_n132 ) , .A1( u1_u4_u4_n152 ) , .B1( u1_u4_u4_n178 ) , .A2( u1_u4_u4_n97 ) );
  AOI22_X1 u1_u4_u4_U94 (.B2( u1_u4_u4_n149 ) , .B1( u1_u4_u4_n150 ) , .A2( u1_u4_u4_n151 ) , .A1( u1_u4_u4_n152 ) , .ZN( u1_u4_u4_n167 ) );
  NOR4_X1 u1_u4_u4_U95 (.A4( u1_u4_u4_n162 ) , .A3( u1_u4_u4_n163 ) , .A2( u1_u4_u4_n164 ) , .A1( u1_u4_u4_n165 ) , .ZN( u1_u4_u4_n166 ) );
  NAND3_X1 u1_u4_u4_U96 (.ZN( u1_out4_3 ) , .A3( u1_u4_u4_n166 ) , .A1( u1_u4_u4_n167 ) , .A2( u1_u4_u4_n186 ) );
  NAND3_X1 u1_u4_u4_U97 (.A3( u1_u4_u4_n146 ) , .A2( u1_u4_u4_n147 ) , .A1( u1_u4_u4_n148 ) , .ZN( u1_u4_u4_n149 ) );
  NAND3_X1 u1_u4_u4_U98 (.A3( u1_u4_u4_n143 ) , .A2( u1_u4_u4_n144 ) , .A1( u1_u4_u4_n145 ) , .ZN( u1_u4_u4_n151 ) );
  NAND3_X1 u1_u4_u4_U99 (.A3( u1_u4_u4_n121 ) , .ZN( u1_u4_u4_n122 ) , .A2( u1_u4_u4_n144 ) , .A1( u1_u4_u4_n154 ) );
  AND3_X1 u1_u4_u7_U10 (.A3( u1_u4_u7_n110 ) , .A2( u1_u4_u7_n127 ) , .A1( u1_u4_u7_n132 ) , .ZN( u1_u4_u7_n92 ) );
  OAI21_X1 u1_u4_u7_U11 (.A( u1_u4_u7_n161 ) , .B1( u1_u4_u7_n168 ) , .B2( u1_u4_u7_n173 ) , .ZN( u1_u4_u7_n91 ) );
  AOI211_X1 u1_u4_u7_U12 (.A( u1_u4_u7_n117 ) , .ZN( u1_u4_u7_n118 ) , .C2( u1_u4_u7_n126 ) , .C1( u1_u4_u7_n177 ) , .B( u1_u4_u7_n180 ) );
  OAI22_X1 u1_u4_u7_U13 (.B1( u1_u4_u7_n115 ) , .ZN( u1_u4_u7_n117 ) , .A2( u1_u4_u7_n133 ) , .A1( u1_u4_u7_n137 ) , .B2( u1_u4_u7_n162 ) );
  INV_X1 u1_u4_u7_U14 (.A( u1_u4_u7_n116 ) , .ZN( u1_u4_u7_n180 ) );
  NOR3_X1 u1_u4_u7_U15 (.ZN( u1_u4_u7_n115 ) , .A3( u1_u4_u7_n145 ) , .A2( u1_u4_u7_n168 ) , .A1( u1_u4_u7_n169 ) );
  NOR3_X1 u1_u4_u7_U16 (.A2( u1_u4_u7_n134 ) , .A1( u1_u4_u7_n135 ) , .ZN( u1_u4_u7_n136 ) , .A3( u1_u4_u7_n171 ) );
  NOR2_X1 u1_u4_u7_U17 (.A1( u1_u4_u7_n130 ) , .A2( u1_u4_u7_n134 ) , .ZN( u1_u4_u7_n153 ) );
  NOR2_X1 u1_u4_u7_U18 (.ZN( u1_u4_u7_n111 ) , .A2( u1_u4_u7_n134 ) , .A1( u1_u4_u7_n169 ) );
  AOI21_X1 u1_u4_u7_U19 (.ZN( u1_u4_u7_n104 ) , .B2( u1_u4_u7_n112 ) , .B1( u1_u4_u7_n127 ) , .A( u1_u4_u7_n164 ) );
  AOI21_X1 u1_u4_u7_U20 (.ZN( u1_u4_u7_n106 ) , .B1( u1_u4_u7_n133 ) , .B2( u1_u4_u7_n146 ) , .A( u1_u4_u7_n162 ) );
  AOI21_X1 u1_u4_u7_U21 (.A( u1_u4_u7_n101 ) , .ZN( u1_u4_u7_n107 ) , .B2( u1_u4_u7_n128 ) , .B1( u1_u4_u7_n175 ) );
  INV_X1 u1_u4_u7_U22 (.A( u1_u4_u7_n101 ) , .ZN( u1_u4_u7_n165 ) );
  INV_X1 u1_u4_u7_U23 (.A( u1_u4_u7_n138 ) , .ZN( u1_u4_u7_n171 ) );
  INV_X1 u1_u4_u7_U24 (.A( u1_u4_u7_n131 ) , .ZN( u1_u4_u7_n177 ) );
  INV_X1 u1_u4_u7_U25 (.A( u1_u4_u7_n110 ) , .ZN( u1_u4_u7_n174 ) );
  NAND2_X1 u1_u4_u7_U26 (.A1( u1_u4_u7_n129 ) , .A2( u1_u4_u7_n132 ) , .ZN( u1_u4_u7_n149 ) );
  NAND2_X1 u1_u4_u7_U27 (.A1( u1_u4_u7_n113 ) , .A2( u1_u4_u7_n124 ) , .ZN( u1_u4_u7_n130 ) );
  INV_X1 u1_u4_u7_U28 (.A( u1_u4_u7_n128 ) , .ZN( u1_u4_u7_n168 ) );
  INV_X1 u1_u4_u7_U29 (.A( u1_u4_u7_n148 ) , .ZN( u1_u4_u7_n169 ) );
  INV_X1 u1_u4_u7_U3 (.A( u1_u4_u7_n149 ) , .ZN( u1_u4_u7_n175 ) );
  INV_X1 u1_u4_u7_U30 (.A( u1_u4_u7_n112 ) , .ZN( u1_u4_u7_n173 ) );
  INV_X1 u1_u4_u7_U31 (.A( u1_u4_u7_n127 ) , .ZN( u1_u4_u7_n179 ) );
  NOR2_X1 u1_u4_u7_U32 (.ZN( u1_u4_u7_n101 ) , .A2( u1_u4_u7_n150 ) , .A1( u1_u4_u7_n156 ) );
  AOI211_X1 u1_u4_u7_U33 (.B( u1_u4_u7_n154 ) , .A( u1_u4_u7_n155 ) , .C1( u1_u4_u7_n156 ) , .ZN( u1_u4_u7_n157 ) , .C2( u1_u4_u7_n172 ) );
  INV_X1 u1_u4_u7_U34 (.A( u1_u4_u7_n153 ) , .ZN( u1_u4_u7_n172 ) );
  AOI211_X1 u1_u4_u7_U35 (.B( u1_u4_u7_n139 ) , .A( u1_u4_u7_n140 ) , .C2( u1_u4_u7_n141 ) , .ZN( u1_u4_u7_n142 ) , .C1( u1_u4_u7_n156 ) );
  NAND4_X1 u1_u4_u7_U36 (.A3( u1_u4_u7_n127 ) , .A2( u1_u4_u7_n128 ) , .A1( u1_u4_u7_n129 ) , .ZN( u1_u4_u7_n141 ) , .A4( u1_u4_u7_n147 ) );
  AOI21_X1 u1_u4_u7_U37 (.A( u1_u4_u7_n137 ) , .B1( u1_u4_u7_n138 ) , .ZN( u1_u4_u7_n139 ) , .B2( u1_u4_u7_n146 ) );
  OAI22_X1 u1_u4_u7_U38 (.B1( u1_u4_u7_n136 ) , .ZN( u1_u4_u7_n140 ) , .A1( u1_u4_u7_n153 ) , .B2( u1_u4_u7_n162 ) , .A2( u1_u4_u7_n164 ) );
  INV_X1 u1_u4_u7_U39 (.A( u1_u4_u7_n125 ) , .ZN( u1_u4_u7_n161 ) );
  INV_X1 u1_u4_u7_U4 (.A( u1_u4_u7_n154 ) , .ZN( u1_u4_u7_n178 ) );
  AOI21_X1 u1_u4_u7_U40 (.ZN( u1_u4_u7_n123 ) , .B1( u1_u4_u7_n165 ) , .B2( u1_u4_u7_n177 ) , .A( u1_u4_u7_n97 ) );
  AOI21_X1 u1_u4_u7_U41 (.B2( u1_u4_u7_n113 ) , .B1( u1_u4_u7_n124 ) , .A( u1_u4_u7_n125 ) , .ZN( u1_u4_u7_n97 ) );
  INV_X1 u1_u4_u7_U42 (.A( u1_u4_u7_n152 ) , .ZN( u1_u4_u7_n162 ) );
  AOI22_X1 u1_u4_u7_U43 (.A2( u1_u4_u7_n114 ) , .ZN( u1_u4_u7_n119 ) , .B1( u1_u4_u7_n130 ) , .A1( u1_u4_u7_n156 ) , .B2( u1_u4_u7_n165 ) );
  NAND2_X1 u1_u4_u7_U44 (.A2( u1_u4_u7_n112 ) , .ZN( u1_u4_u7_n114 ) , .A1( u1_u4_u7_n175 ) );
  AOI22_X1 u1_u4_u7_U45 (.B2( u1_u4_u7_n149 ) , .B1( u1_u4_u7_n150 ) , .A2( u1_u4_u7_n151 ) , .A1( u1_u4_u7_n152 ) , .ZN( u1_u4_u7_n158 ) );
  NOR2_X1 u1_u4_u7_U46 (.ZN( u1_u4_u7_n137 ) , .A1( u1_u4_u7_n150 ) , .A2( u1_u4_u7_n161 ) );
  AND2_X1 u1_u4_u7_U47 (.ZN( u1_u4_u7_n145 ) , .A2( u1_u4_u7_n98 ) , .A1( u1_u4_u7_n99 ) );
  AOI21_X1 u1_u4_u7_U48 (.ZN( u1_u4_u7_n105 ) , .B2( u1_u4_u7_n110 ) , .A( u1_u4_u7_n125 ) , .B1( u1_u4_u7_n147 ) );
  NAND2_X1 u1_u4_u7_U49 (.ZN( u1_u4_u7_n146 ) , .A1( u1_u4_u7_n95 ) , .A2( u1_u4_u7_n98 ) );
  INV_X1 u1_u4_u7_U5 (.A( u1_u4_u7_n111 ) , .ZN( u1_u4_u7_n170 ) );
  NAND2_X1 u1_u4_u7_U50 (.A2( u1_u4_u7_n103 ) , .ZN( u1_u4_u7_n147 ) , .A1( u1_u4_u7_n93 ) );
  NAND2_X1 u1_u4_u7_U51 (.A1( u1_u4_u7_n103 ) , .ZN( u1_u4_u7_n127 ) , .A2( u1_u4_u7_n99 ) );
  NAND2_X1 u1_u4_u7_U52 (.A2( u1_u4_u7_n102 ) , .A1( u1_u4_u7_n103 ) , .ZN( u1_u4_u7_n133 ) );
  OR2_X1 u1_u4_u7_U53 (.ZN( u1_u4_u7_n126 ) , .A2( u1_u4_u7_n152 ) , .A1( u1_u4_u7_n156 ) );
  NAND2_X1 u1_u4_u7_U54 (.ZN( u1_u4_u7_n112 ) , .A2( u1_u4_u7_n96 ) , .A1( u1_u4_u7_n99 ) );
  NAND2_X1 u1_u4_u7_U55 (.A2( u1_u4_u7_n102 ) , .ZN( u1_u4_u7_n128 ) , .A1( u1_u4_u7_n98 ) );
  INV_X1 u1_u4_u7_U56 (.A( u1_u4_u7_n150 ) , .ZN( u1_u4_u7_n164 ) );
  AND2_X1 u1_u4_u7_U57 (.ZN( u1_u4_u7_n134 ) , .A1( u1_u4_u7_n93 ) , .A2( u1_u4_u7_n98 ) );
  NAND2_X1 u1_u4_u7_U58 (.ZN( u1_u4_u7_n110 ) , .A1( u1_u4_u7_n95 ) , .A2( u1_u4_u7_n96 ) );
  NAND2_X1 u1_u4_u7_U59 (.A2( u1_u4_u7_n102 ) , .ZN( u1_u4_u7_n124 ) , .A1( u1_u4_u7_n96 ) );
  AOI211_X1 u1_u4_u7_U6 (.ZN( u1_u4_u7_n116 ) , .A( u1_u4_u7_n155 ) , .C1( u1_u4_u7_n161 ) , .C2( u1_u4_u7_n171 ) , .B( u1_u4_u7_n94 ) );
  NAND2_X1 u1_u4_u7_U60 (.ZN( u1_u4_u7_n132 ) , .A1( u1_u4_u7_n93 ) , .A2( u1_u4_u7_n96 ) );
  NAND2_X1 u1_u4_u7_U61 (.A2( u1_u4_u7_n103 ) , .ZN( u1_u4_u7_n131 ) , .A1( u1_u4_u7_n95 ) );
  NOR2_X1 u1_u4_u7_U62 (.A2( u1_u4_X_47 ) , .ZN( u1_u4_u7_n150 ) , .A1( u1_u4_u7_n163 ) );
  NOR2_X1 u1_u4_u7_U63 (.A2( u1_u4_X_43 ) , .A1( u1_u4_X_44 ) , .ZN( u1_u4_u7_n103 ) );
  NOR2_X1 u1_u4_u7_U64 (.A2( u1_u4_X_48 ) , .A1( u1_u4_u7_n166 ) , .ZN( u1_u4_u7_n95 ) );
  NOR2_X1 u1_u4_u7_U65 (.A2( u1_u4_X_44 ) , .A1( u1_u4_u7_n167 ) , .ZN( u1_u4_u7_n98 ) );
  NOR2_X1 u1_u4_u7_U66 (.A2( u1_u4_X_45 ) , .A1( u1_u4_X_48 ) , .ZN( u1_u4_u7_n99 ) );
  NOR2_X1 u1_u4_u7_U67 (.A2( u1_u4_X_46 ) , .A1( u1_u4_X_47 ) , .ZN( u1_u4_u7_n152 ) );
  AND2_X1 u1_u4_u7_U68 (.A1( u1_u4_X_47 ) , .ZN( u1_u4_u7_n156 ) , .A2( u1_u4_u7_n163 ) );
  NAND2_X1 u1_u4_u7_U69 (.A2( u1_u4_X_46 ) , .A1( u1_u4_X_47 ) , .ZN( u1_u4_u7_n125 ) );
  OAI222_X1 u1_u4_u7_U7 (.C2( u1_u4_u7_n101 ) , .B2( u1_u4_u7_n111 ) , .A1( u1_u4_u7_n113 ) , .C1( u1_u4_u7_n146 ) , .A2( u1_u4_u7_n162 ) , .B1( u1_u4_u7_n164 ) , .ZN( u1_u4_u7_n94 ) );
  AND2_X1 u1_u4_u7_U70 (.A2( u1_u4_X_43 ) , .A1( u1_u4_X_44 ) , .ZN( u1_u4_u7_n96 ) );
  AND2_X1 u1_u4_u7_U71 (.A2( u1_u4_X_45 ) , .A1( u1_u4_X_48 ) , .ZN( u1_u4_u7_n102 ) );
  AND2_X1 u1_u4_u7_U72 (.A1( u1_u4_X_48 ) , .A2( u1_u4_u7_n166 ) , .ZN( u1_u4_u7_n93 ) );
  INV_X1 u1_u4_u7_U73 (.A( u1_u4_X_46 ) , .ZN( u1_u4_u7_n163 ) );
  AND2_X1 u1_u4_u7_U74 (.A1( u1_u4_X_44 ) , .ZN( u1_u4_u7_n100 ) , .A2( u1_u4_u7_n167 ) );
  INV_X1 u1_u4_u7_U75 (.A( u1_u4_X_45 ) , .ZN( u1_u4_u7_n166 ) );
  INV_X1 u1_u4_u7_U76 (.A( u1_u4_X_43 ) , .ZN( u1_u4_u7_n167 ) );
  NAND4_X1 u1_u4_u7_U77 (.ZN( u1_out4_5 ) , .A4( u1_u4_u7_n108 ) , .A3( u1_u4_u7_n109 ) , .A1( u1_u4_u7_n116 ) , .A2( u1_u4_u7_n123 ) );
  AOI22_X1 u1_u4_u7_U78 (.ZN( u1_u4_u7_n109 ) , .A2( u1_u4_u7_n126 ) , .B2( u1_u4_u7_n145 ) , .B1( u1_u4_u7_n156 ) , .A1( u1_u4_u7_n171 ) );
  NOR4_X1 u1_u4_u7_U79 (.A4( u1_u4_u7_n104 ) , .A3( u1_u4_u7_n105 ) , .A2( u1_u4_u7_n106 ) , .A1( u1_u4_u7_n107 ) , .ZN( u1_u4_u7_n108 ) );
  INV_X1 u1_u4_u7_U8 (.A( u1_u4_u7_n133 ) , .ZN( u1_u4_u7_n176 ) );
  NAND4_X1 u1_u4_u7_U80 (.ZN( u1_out4_27 ) , .A4( u1_u4_u7_n118 ) , .A3( u1_u4_u7_n119 ) , .A2( u1_u4_u7_n120 ) , .A1( u1_u4_u7_n121 ) );
  OAI21_X1 u1_u4_u7_U81 (.ZN( u1_u4_u7_n121 ) , .B2( u1_u4_u7_n145 ) , .A( u1_u4_u7_n150 ) , .B1( u1_u4_u7_n174 ) );
  OAI21_X1 u1_u4_u7_U82 (.ZN( u1_u4_u7_n120 ) , .A( u1_u4_u7_n161 ) , .B2( u1_u4_u7_n170 ) , .B1( u1_u4_u7_n179 ) );
  NAND4_X1 u1_u4_u7_U83 (.ZN( u1_out4_21 ) , .A4( u1_u4_u7_n157 ) , .A3( u1_u4_u7_n158 ) , .A2( u1_u4_u7_n159 ) , .A1( u1_u4_u7_n160 ) );
  OAI21_X1 u1_u4_u7_U84 (.B1( u1_u4_u7_n145 ) , .ZN( u1_u4_u7_n160 ) , .A( u1_u4_u7_n161 ) , .B2( u1_u4_u7_n177 ) );
  OAI21_X1 u1_u4_u7_U85 (.ZN( u1_u4_u7_n159 ) , .A( u1_u4_u7_n165 ) , .B2( u1_u4_u7_n171 ) , .B1( u1_u4_u7_n174 ) );
  NAND4_X1 u1_u4_u7_U86 (.ZN( u1_out4_15 ) , .A4( u1_u4_u7_n142 ) , .A3( u1_u4_u7_n143 ) , .A2( u1_u4_u7_n144 ) , .A1( u1_u4_u7_n178 ) );
  OR2_X1 u1_u4_u7_U87 (.A2( u1_u4_u7_n125 ) , .A1( u1_u4_u7_n129 ) , .ZN( u1_u4_u7_n144 ) );
  AOI22_X1 u1_u4_u7_U88 (.A2( u1_u4_u7_n126 ) , .ZN( u1_u4_u7_n143 ) , .B2( u1_u4_u7_n165 ) , .B1( u1_u4_u7_n173 ) , .A1( u1_u4_u7_n174 ) );
  NAND2_X1 u1_u4_u7_U89 (.A1( u1_u4_u7_n100 ) , .ZN( u1_u4_u7_n148 ) , .A2( u1_u4_u7_n95 ) );
  OAI221_X1 u1_u4_u7_U9 (.C1( u1_u4_u7_n101 ) , .C2( u1_u4_u7_n147 ) , .ZN( u1_u4_u7_n155 ) , .B2( u1_u4_u7_n162 ) , .A( u1_u4_u7_n91 ) , .B1( u1_u4_u7_n92 ) );
  NAND2_X1 u1_u4_u7_U90 (.A1( u1_u4_u7_n100 ) , .ZN( u1_u4_u7_n113 ) , .A2( u1_u4_u7_n93 ) );
  NAND2_X1 u1_u4_u7_U91 (.A1( u1_u4_u7_n100 ) , .ZN( u1_u4_u7_n138 ) , .A2( u1_u4_u7_n99 ) );
  NAND2_X1 u1_u4_u7_U92 (.A1( u1_u4_u7_n100 ) , .A2( u1_u4_u7_n102 ) , .ZN( u1_u4_u7_n129 ) );
  OAI211_X1 u1_u4_u7_U93 (.B( u1_u4_u7_n122 ) , .A( u1_u4_u7_n123 ) , .C2( u1_u4_u7_n124 ) , .ZN( u1_u4_u7_n154 ) , .C1( u1_u4_u7_n162 ) );
  AOI222_X1 u1_u4_u7_U94 (.ZN( u1_u4_u7_n122 ) , .C2( u1_u4_u7_n126 ) , .C1( u1_u4_u7_n145 ) , .B1( u1_u4_u7_n161 ) , .A2( u1_u4_u7_n165 ) , .B2( u1_u4_u7_n170 ) , .A1( u1_u4_u7_n176 ) );
  NAND3_X1 u1_u4_u7_U95 (.A3( u1_u4_u7_n146 ) , .A2( u1_u4_u7_n147 ) , .A1( u1_u4_u7_n148 ) , .ZN( u1_u4_u7_n151 ) );
  NAND3_X1 u1_u4_u7_U96 (.A3( u1_u4_u7_n131 ) , .A2( u1_u4_u7_n132 ) , .A1( u1_u4_u7_n133 ) , .ZN( u1_u4_u7_n135 ) );
  XOR2_X1 u1_u6_U1 (.B( u1_K7_9 ) , .A( u1_R5_6 ) , .Z( u1_u6_X_9 ) );
  XOR2_X1 u1_u6_U10 (.B( u1_K7_45 ) , .A( u1_R5_30 ) , .Z( u1_u6_X_45 ) );
  XOR2_X1 u1_u6_U11 (.B( u1_K7_44 ) , .A( u1_R5_29 ) , .Z( u1_u6_X_44 ) );
  XOR2_X1 u1_u6_U12 (.B( u1_K7_43 ) , .A( u1_R5_28 ) , .Z( u1_u6_X_43 ) );
  XOR2_X1 u1_u6_U13 (.B( u1_K7_42 ) , .A( u1_R5_29 ) , .Z( u1_u6_X_42 ) );
  XOR2_X1 u1_u6_U14 (.B( u1_K7_41 ) , .A( u1_R5_28 ) , .Z( u1_u6_X_41 ) );
  XOR2_X1 u1_u6_U15 (.B( u1_K7_40 ) , .A( u1_R5_27 ) , .Z( u1_u6_X_40 ) );
  XOR2_X1 u1_u6_U17 (.B( u1_K7_39 ) , .A( u1_R5_26 ) , .Z( u1_u6_X_39 ) );
  XOR2_X1 u1_u6_U18 (.B( u1_K7_38 ) , .A( u1_R5_25 ) , .Z( u1_u6_X_38 ) );
  XOR2_X1 u1_u6_U19 (.B( u1_K7_37 ) , .A( u1_R5_24 ) , .Z( u1_u6_X_37 ) );
  XOR2_X1 u1_u6_U2 (.B( u1_K7_8 ) , .A( u1_R5_5 ) , .Z( u1_u6_X_8 ) );
  XOR2_X1 u1_u6_U3 (.B( u1_K7_7 ) , .A( u1_R5_4 ) , .Z( u1_u6_X_7 ) );
  XOR2_X1 u1_u6_U40 (.B( u1_K7_18 ) , .A( u1_R5_13 ) , .Z( u1_u6_X_18 ) );
  XOR2_X1 u1_u6_U41 (.B( u1_K7_17 ) , .A( u1_R5_12 ) , .Z( u1_u6_X_17 ) );
  XOR2_X1 u1_u6_U42 (.B( u1_K7_16 ) , .A( u1_R5_11 ) , .Z( u1_u6_X_16 ) );
  XOR2_X1 u1_u6_U43 (.B( u1_K7_15 ) , .A( u1_R5_10 ) , .Z( u1_u6_X_15 ) );
  XOR2_X1 u1_u6_U44 (.B( u1_K7_14 ) , .A( u1_R5_9 ) , .Z( u1_u6_X_14 ) );
  XOR2_X1 u1_u6_U45 (.B( u1_K7_13 ) , .A( u1_R5_8 ) , .Z( u1_u6_X_13 ) );
  XOR2_X1 u1_u6_U46 (.B( u1_K7_12 ) , .A( u1_R5_9 ) , .Z( u1_u6_X_12 ) );
  XOR2_X1 u1_u6_U47 (.B( u1_K7_11 ) , .A( u1_R5_8 ) , .Z( u1_u6_X_11 ) );
  XOR2_X1 u1_u6_U48 (.B( u1_K7_10 ) , .A( u1_R5_7 ) , .Z( u1_u6_X_10 ) );
  XOR2_X1 u1_u6_U7 (.B( u1_K7_48 ) , .A( u1_R5_1 ) , .Z( u1_u6_X_48 ) );
  XOR2_X1 u1_u6_U8 (.B( u1_K7_47 ) , .A( u1_R5_32 ) , .Z( u1_u6_X_47 ) );
  XOR2_X1 u1_u6_U9 (.B( u1_K7_46 ) , .A( u1_R5_31 ) , .Z( u1_u6_X_46 ) );
  NOR2_X1 u1_u6_u1_U10 (.A1( u1_u6_u1_n112 ) , .A2( u1_u6_u1_n116 ) , .ZN( u1_u6_u1_n118 ) );
  NAND3_X1 u1_u6_u1_U100 (.ZN( u1_u6_u1_n113 ) , .A1( u1_u6_u1_n120 ) , .A3( u1_u6_u1_n133 ) , .A2( u1_u6_u1_n155 ) );
  OAI21_X1 u1_u6_u1_U11 (.ZN( u1_u6_u1_n101 ) , .B1( u1_u6_u1_n141 ) , .A( u1_u6_u1_n146 ) , .B2( u1_u6_u1_n183 ) );
  AOI21_X1 u1_u6_u1_U12 (.B2( u1_u6_u1_n155 ) , .B1( u1_u6_u1_n156 ) , .ZN( u1_u6_u1_n157 ) , .A( u1_u6_u1_n174 ) );
  NAND2_X1 u1_u6_u1_U13 (.ZN( u1_u6_u1_n140 ) , .A2( u1_u6_u1_n150 ) , .A1( u1_u6_u1_n155 ) );
  NAND2_X1 u1_u6_u1_U14 (.A1( u1_u6_u1_n131 ) , .ZN( u1_u6_u1_n147 ) , .A2( u1_u6_u1_n153 ) );
  INV_X1 u1_u6_u1_U15 (.A( u1_u6_u1_n139 ) , .ZN( u1_u6_u1_n174 ) );
  OR4_X1 u1_u6_u1_U16 (.A4( u1_u6_u1_n106 ) , .A3( u1_u6_u1_n107 ) , .ZN( u1_u6_u1_n108 ) , .A1( u1_u6_u1_n117 ) , .A2( u1_u6_u1_n184 ) );
  AOI21_X1 u1_u6_u1_U17 (.ZN( u1_u6_u1_n106 ) , .A( u1_u6_u1_n112 ) , .B1( u1_u6_u1_n154 ) , .B2( u1_u6_u1_n156 ) );
  AOI21_X1 u1_u6_u1_U18 (.ZN( u1_u6_u1_n107 ) , .B1( u1_u6_u1_n134 ) , .B2( u1_u6_u1_n149 ) , .A( u1_u6_u1_n174 ) );
  INV_X1 u1_u6_u1_U19 (.A( u1_u6_u1_n101 ) , .ZN( u1_u6_u1_n184 ) );
  INV_X1 u1_u6_u1_U20 (.A( u1_u6_u1_n112 ) , .ZN( u1_u6_u1_n171 ) );
  NAND2_X1 u1_u6_u1_U21 (.ZN( u1_u6_u1_n141 ) , .A1( u1_u6_u1_n153 ) , .A2( u1_u6_u1_n156 ) );
  AND2_X1 u1_u6_u1_U22 (.A1( u1_u6_u1_n123 ) , .ZN( u1_u6_u1_n134 ) , .A2( u1_u6_u1_n161 ) );
  NAND2_X1 u1_u6_u1_U23 (.A2( u1_u6_u1_n115 ) , .A1( u1_u6_u1_n116 ) , .ZN( u1_u6_u1_n148 ) );
  NAND2_X1 u1_u6_u1_U24 (.A2( u1_u6_u1_n133 ) , .A1( u1_u6_u1_n135 ) , .ZN( u1_u6_u1_n159 ) );
  NAND2_X1 u1_u6_u1_U25 (.A2( u1_u6_u1_n115 ) , .A1( u1_u6_u1_n120 ) , .ZN( u1_u6_u1_n132 ) );
  INV_X1 u1_u6_u1_U26 (.A( u1_u6_u1_n154 ) , .ZN( u1_u6_u1_n178 ) );
  INV_X1 u1_u6_u1_U27 (.A( u1_u6_u1_n151 ) , .ZN( u1_u6_u1_n183 ) );
  AND2_X1 u1_u6_u1_U28 (.A1( u1_u6_u1_n129 ) , .A2( u1_u6_u1_n133 ) , .ZN( u1_u6_u1_n149 ) );
  INV_X1 u1_u6_u1_U29 (.A( u1_u6_u1_n131 ) , .ZN( u1_u6_u1_n180 ) );
  INV_X1 u1_u6_u1_U3 (.A( u1_u6_u1_n159 ) , .ZN( u1_u6_u1_n182 ) );
  AOI221_X1 u1_u6_u1_U30 (.B1( u1_u6_u1_n140 ) , .ZN( u1_u6_u1_n167 ) , .B2( u1_u6_u1_n172 ) , .C2( u1_u6_u1_n175 ) , .C1( u1_u6_u1_n178 ) , .A( u1_u6_u1_n188 ) );
  INV_X1 u1_u6_u1_U31 (.ZN( u1_u6_u1_n188 ) , .A( u1_u6_u1_n97 ) );
  AOI211_X1 u1_u6_u1_U32 (.A( u1_u6_u1_n118 ) , .C1( u1_u6_u1_n132 ) , .C2( u1_u6_u1_n139 ) , .B( u1_u6_u1_n96 ) , .ZN( u1_u6_u1_n97 ) );
  AOI21_X1 u1_u6_u1_U33 (.B2( u1_u6_u1_n121 ) , .B1( u1_u6_u1_n135 ) , .A( u1_u6_u1_n152 ) , .ZN( u1_u6_u1_n96 ) );
  OAI221_X1 u1_u6_u1_U34 (.A( u1_u6_u1_n119 ) , .C2( u1_u6_u1_n129 ) , .ZN( u1_u6_u1_n138 ) , .B2( u1_u6_u1_n152 ) , .C1( u1_u6_u1_n174 ) , .B1( u1_u6_u1_n187 ) );
  INV_X1 u1_u6_u1_U35 (.A( u1_u6_u1_n148 ) , .ZN( u1_u6_u1_n187 ) );
  AOI211_X1 u1_u6_u1_U36 (.B( u1_u6_u1_n117 ) , .A( u1_u6_u1_n118 ) , .ZN( u1_u6_u1_n119 ) , .C2( u1_u6_u1_n146 ) , .C1( u1_u6_u1_n159 ) );
  NOR2_X1 u1_u6_u1_U37 (.A1( u1_u6_u1_n168 ) , .A2( u1_u6_u1_n176 ) , .ZN( u1_u6_u1_n98 ) );
  AOI211_X1 u1_u6_u1_U38 (.B( u1_u6_u1_n162 ) , .A( u1_u6_u1_n163 ) , .C2( u1_u6_u1_n164 ) , .ZN( u1_u6_u1_n165 ) , .C1( u1_u6_u1_n171 ) );
  AOI21_X1 u1_u6_u1_U39 (.A( u1_u6_u1_n160 ) , .B2( u1_u6_u1_n161 ) , .ZN( u1_u6_u1_n162 ) , .B1( u1_u6_u1_n182 ) );
  AOI221_X1 u1_u6_u1_U4 (.A( u1_u6_u1_n138 ) , .C2( u1_u6_u1_n139 ) , .C1( u1_u6_u1_n140 ) , .B2( u1_u6_u1_n141 ) , .ZN( u1_u6_u1_n142 ) , .B1( u1_u6_u1_n175 ) );
  OR2_X1 u1_u6_u1_U40 (.A2( u1_u6_u1_n157 ) , .A1( u1_u6_u1_n158 ) , .ZN( u1_u6_u1_n163 ) );
  NAND2_X1 u1_u6_u1_U41 (.A1( u1_u6_u1_n128 ) , .ZN( u1_u6_u1_n146 ) , .A2( u1_u6_u1_n160 ) );
  NAND2_X1 u1_u6_u1_U42 (.A2( u1_u6_u1_n112 ) , .ZN( u1_u6_u1_n139 ) , .A1( u1_u6_u1_n152 ) );
  NAND2_X1 u1_u6_u1_U43 (.A1( u1_u6_u1_n105 ) , .ZN( u1_u6_u1_n156 ) , .A2( u1_u6_u1_n99 ) );
  NOR2_X1 u1_u6_u1_U44 (.ZN( u1_u6_u1_n117 ) , .A1( u1_u6_u1_n121 ) , .A2( u1_u6_u1_n160 ) );
  OAI21_X1 u1_u6_u1_U45 (.B2( u1_u6_u1_n123 ) , .ZN( u1_u6_u1_n145 ) , .B1( u1_u6_u1_n160 ) , .A( u1_u6_u1_n185 ) );
  INV_X1 u1_u6_u1_U46 (.A( u1_u6_u1_n122 ) , .ZN( u1_u6_u1_n185 ) );
  AOI21_X1 u1_u6_u1_U47 (.B2( u1_u6_u1_n120 ) , .B1( u1_u6_u1_n121 ) , .ZN( u1_u6_u1_n122 ) , .A( u1_u6_u1_n128 ) );
  AOI21_X1 u1_u6_u1_U48 (.A( u1_u6_u1_n128 ) , .B2( u1_u6_u1_n129 ) , .ZN( u1_u6_u1_n130 ) , .B1( u1_u6_u1_n150 ) );
  NAND2_X1 u1_u6_u1_U49 (.ZN( u1_u6_u1_n112 ) , .A1( u1_u6_u1_n169 ) , .A2( u1_u6_u1_n170 ) );
  AOI211_X1 u1_u6_u1_U5 (.ZN( u1_u6_u1_n124 ) , .A( u1_u6_u1_n138 ) , .C2( u1_u6_u1_n139 ) , .B( u1_u6_u1_n145 ) , .C1( u1_u6_u1_n147 ) );
  NAND2_X1 u1_u6_u1_U50 (.ZN( u1_u6_u1_n129 ) , .A2( u1_u6_u1_n95 ) , .A1( u1_u6_u1_n98 ) );
  NAND2_X1 u1_u6_u1_U51 (.A1( u1_u6_u1_n102 ) , .ZN( u1_u6_u1_n154 ) , .A2( u1_u6_u1_n99 ) );
  NAND2_X1 u1_u6_u1_U52 (.A2( u1_u6_u1_n100 ) , .ZN( u1_u6_u1_n135 ) , .A1( u1_u6_u1_n99 ) );
  AOI21_X1 u1_u6_u1_U53 (.A( u1_u6_u1_n152 ) , .B2( u1_u6_u1_n153 ) , .B1( u1_u6_u1_n154 ) , .ZN( u1_u6_u1_n158 ) );
  INV_X1 u1_u6_u1_U54 (.A( u1_u6_u1_n160 ) , .ZN( u1_u6_u1_n175 ) );
  NAND2_X1 u1_u6_u1_U55 (.A1( u1_u6_u1_n100 ) , .ZN( u1_u6_u1_n116 ) , .A2( u1_u6_u1_n95 ) );
  NAND2_X1 u1_u6_u1_U56 (.A1( u1_u6_u1_n102 ) , .ZN( u1_u6_u1_n131 ) , .A2( u1_u6_u1_n95 ) );
  NAND2_X1 u1_u6_u1_U57 (.A2( u1_u6_u1_n104 ) , .ZN( u1_u6_u1_n121 ) , .A1( u1_u6_u1_n98 ) );
  NAND2_X1 u1_u6_u1_U58 (.A1( u1_u6_u1_n103 ) , .ZN( u1_u6_u1_n153 ) , .A2( u1_u6_u1_n98 ) );
  NAND2_X1 u1_u6_u1_U59 (.A2( u1_u6_u1_n104 ) , .A1( u1_u6_u1_n105 ) , .ZN( u1_u6_u1_n133 ) );
  AOI22_X1 u1_u6_u1_U6 (.B2( u1_u6_u1_n113 ) , .A2( u1_u6_u1_n114 ) , .ZN( u1_u6_u1_n125 ) , .A1( u1_u6_u1_n171 ) , .B1( u1_u6_u1_n173 ) );
  NAND2_X1 u1_u6_u1_U60 (.ZN( u1_u6_u1_n150 ) , .A2( u1_u6_u1_n98 ) , .A1( u1_u6_u1_n99 ) );
  NAND2_X1 u1_u6_u1_U61 (.A1( u1_u6_u1_n105 ) , .ZN( u1_u6_u1_n155 ) , .A2( u1_u6_u1_n95 ) );
  OAI21_X1 u1_u6_u1_U62 (.ZN( u1_u6_u1_n109 ) , .B1( u1_u6_u1_n129 ) , .B2( u1_u6_u1_n160 ) , .A( u1_u6_u1_n167 ) );
  NAND2_X1 u1_u6_u1_U63 (.A2( u1_u6_u1_n100 ) , .A1( u1_u6_u1_n103 ) , .ZN( u1_u6_u1_n120 ) );
  NAND2_X1 u1_u6_u1_U64 (.A1( u1_u6_u1_n102 ) , .A2( u1_u6_u1_n104 ) , .ZN( u1_u6_u1_n115 ) );
  NAND2_X1 u1_u6_u1_U65 (.A2( u1_u6_u1_n100 ) , .A1( u1_u6_u1_n104 ) , .ZN( u1_u6_u1_n151 ) );
  NAND2_X1 u1_u6_u1_U66 (.A2( u1_u6_u1_n103 ) , .A1( u1_u6_u1_n105 ) , .ZN( u1_u6_u1_n161 ) );
  INV_X1 u1_u6_u1_U67 (.A( u1_u6_u1_n152 ) , .ZN( u1_u6_u1_n173 ) );
  INV_X1 u1_u6_u1_U68 (.A( u1_u6_u1_n128 ) , .ZN( u1_u6_u1_n172 ) );
  NAND2_X1 u1_u6_u1_U69 (.A2( u1_u6_u1_n102 ) , .A1( u1_u6_u1_n103 ) , .ZN( u1_u6_u1_n123 ) );
  NAND2_X1 u1_u6_u1_U7 (.ZN( u1_u6_u1_n114 ) , .A1( u1_u6_u1_n134 ) , .A2( u1_u6_u1_n156 ) );
  NOR2_X1 u1_u6_u1_U70 (.A2( u1_u6_X_7 ) , .A1( u1_u6_X_8 ) , .ZN( u1_u6_u1_n95 ) );
  NOR2_X1 u1_u6_u1_U71 (.A1( u1_u6_X_12 ) , .A2( u1_u6_X_9 ) , .ZN( u1_u6_u1_n100 ) );
  NOR2_X1 u1_u6_u1_U72 (.A2( u1_u6_X_8 ) , .A1( u1_u6_u1_n177 ) , .ZN( u1_u6_u1_n99 ) );
  NOR2_X1 u1_u6_u1_U73 (.A2( u1_u6_X_12 ) , .ZN( u1_u6_u1_n102 ) , .A1( u1_u6_u1_n176 ) );
  NOR2_X1 u1_u6_u1_U74 (.A2( u1_u6_X_9 ) , .ZN( u1_u6_u1_n105 ) , .A1( u1_u6_u1_n168 ) );
  NAND2_X1 u1_u6_u1_U75 (.A1( u1_u6_X_10 ) , .ZN( u1_u6_u1_n160 ) , .A2( u1_u6_u1_n169 ) );
  NAND2_X1 u1_u6_u1_U76 (.A2( u1_u6_X_10 ) , .A1( u1_u6_X_11 ) , .ZN( u1_u6_u1_n152 ) );
  NAND2_X1 u1_u6_u1_U77 (.A1( u1_u6_X_11 ) , .ZN( u1_u6_u1_n128 ) , .A2( u1_u6_u1_n170 ) );
  AND2_X1 u1_u6_u1_U78 (.A2( u1_u6_X_7 ) , .A1( u1_u6_X_8 ) , .ZN( u1_u6_u1_n104 ) );
  AND2_X1 u1_u6_u1_U79 (.A1( u1_u6_X_8 ) , .ZN( u1_u6_u1_n103 ) , .A2( u1_u6_u1_n177 ) );
  AOI22_X1 u1_u6_u1_U8 (.B2( u1_u6_u1_n136 ) , .A2( u1_u6_u1_n137 ) , .ZN( u1_u6_u1_n143 ) , .A1( u1_u6_u1_n171 ) , .B1( u1_u6_u1_n173 ) );
  INV_X1 u1_u6_u1_U80 (.A( u1_u6_X_10 ) , .ZN( u1_u6_u1_n170 ) );
  INV_X1 u1_u6_u1_U81 (.A( u1_u6_X_9 ) , .ZN( u1_u6_u1_n176 ) );
  INV_X1 u1_u6_u1_U82 (.A( u1_u6_X_11 ) , .ZN( u1_u6_u1_n169 ) );
  INV_X1 u1_u6_u1_U83 (.A( u1_u6_X_12 ) , .ZN( u1_u6_u1_n168 ) );
  INV_X1 u1_u6_u1_U84 (.A( u1_u6_X_7 ) , .ZN( u1_u6_u1_n177 ) );
  NAND4_X1 u1_u6_u1_U85 (.ZN( u1_out6_18 ) , .A4( u1_u6_u1_n165 ) , .A3( u1_u6_u1_n166 ) , .A1( u1_u6_u1_n167 ) , .A2( u1_u6_u1_n186 ) );
  AOI22_X1 u1_u6_u1_U86 (.B2( u1_u6_u1_n146 ) , .B1( u1_u6_u1_n147 ) , .A2( u1_u6_u1_n148 ) , .ZN( u1_u6_u1_n166 ) , .A1( u1_u6_u1_n172 ) );
  INV_X1 u1_u6_u1_U87 (.A( u1_u6_u1_n145 ) , .ZN( u1_u6_u1_n186 ) );
  NAND4_X1 u1_u6_u1_U88 (.ZN( u1_out6_2 ) , .A4( u1_u6_u1_n142 ) , .A3( u1_u6_u1_n143 ) , .A2( u1_u6_u1_n144 ) , .A1( u1_u6_u1_n179 ) );
  OAI21_X1 u1_u6_u1_U89 (.B2( u1_u6_u1_n132 ) , .ZN( u1_u6_u1_n144 ) , .A( u1_u6_u1_n146 ) , .B1( u1_u6_u1_n180 ) );
  INV_X1 u1_u6_u1_U9 (.A( u1_u6_u1_n147 ) , .ZN( u1_u6_u1_n181 ) );
  INV_X1 u1_u6_u1_U90 (.A( u1_u6_u1_n130 ) , .ZN( u1_u6_u1_n179 ) );
  NAND4_X1 u1_u6_u1_U91 (.ZN( u1_out6_28 ) , .A4( u1_u6_u1_n124 ) , .A3( u1_u6_u1_n125 ) , .A2( u1_u6_u1_n126 ) , .A1( u1_u6_u1_n127 ) );
  OAI21_X1 u1_u6_u1_U92 (.ZN( u1_u6_u1_n127 ) , .B2( u1_u6_u1_n139 ) , .B1( u1_u6_u1_n175 ) , .A( u1_u6_u1_n183 ) );
  OAI21_X1 u1_u6_u1_U93 (.ZN( u1_u6_u1_n126 ) , .B2( u1_u6_u1_n140 ) , .A( u1_u6_u1_n146 ) , .B1( u1_u6_u1_n178 ) );
  OR4_X1 u1_u6_u1_U94 (.ZN( u1_out6_13 ) , .A4( u1_u6_u1_n108 ) , .A3( u1_u6_u1_n109 ) , .A2( u1_u6_u1_n110 ) , .A1( u1_u6_u1_n111 ) );
  AOI21_X1 u1_u6_u1_U95 (.ZN( u1_u6_u1_n111 ) , .A( u1_u6_u1_n128 ) , .B2( u1_u6_u1_n131 ) , .B1( u1_u6_u1_n135 ) );
  AOI21_X1 u1_u6_u1_U96 (.ZN( u1_u6_u1_n110 ) , .A( u1_u6_u1_n116 ) , .B1( u1_u6_u1_n152 ) , .B2( u1_u6_u1_n160 ) );
  NAND3_X1 u1_u6_u1_U97 (.A3( u1_u6_u1_n149 ) , .A2( u1_u6_u1_n150 ) , .A1( u1_u6_u1_n151 ) , .ZN( u1_u6_u1_n164 ) );
  NAND3_X1 u1_u6_u1_U98 (.A3( u1_u6_u1_n134 ) , .A2( u1_u6_u1_n135 ) , .ZN( u1_u6_u1_n136 ) , .A1( u1_u6_u1_n151 ) );
  NAND3_X1 u1_u6_u1_U99 (.A1( u1_u6_u1_n133 ) , .ZN( u1_u6_u1_n137 ) , .A2( u1_u6_u1_n154 ) , .A3( u1_u6_u1_n181 ) );
  OAI22_X1 u1_u6_u2_U10 (.B1( u1_u6_u2_n151 ) , .A2( u1_u6_u2_n152 ) , .A1( u1_u6_u2_n153 ) , .ZN( u1_u6_u2_n160 ) , .B2( u1_u6_u2_n168 ) );
  NAND3_X1 u1_u6_u2_U100 (.A2( u1_u6_u2_n100 ) , .A1( u1_u6_u2_n104 ) , .A3( u1_u6_u2_n138 ) , .ZN( u1_u6_u2_n98 ) );
  NOR3_X1 u1_u6_u2_U11 (.A1( u1_u6_u2_n150 ) , .ZN( u1_u6_u2_n151 ) , .A3( u1_u6_u2_n175 ) , .A2( u1_u6_u2_n188 ) );
  AOI21_X1 u1_u6_u2_U12 (.B2( u1_u6_u2_n123 ) , .ZN( u1_u6_u2_n125 ) , .A( u1_u6_u2_n171 ) , .B1( u1_u6_u2_n184 ) );
  INV_X1 u1_u6_u2_U13 (.A( u1_u6_u2_n150 ) , .ZN( u1_u6_u2_n184 ) );
  AOI21_X1 u1_u6_u2_U14 (.ZN( u1_u6_u2_n144 ) , .B2( u1_u6_u2_n155 ) , .A( u1_u6_u2_n172 ) , .B1( u1_u6_u2_n185 ) );
  AOI21_X1 u1_u6_u2_U15 (.B2( u1_u6_u2_n143 ) , .ZN( u1_u6_u2_n145 ) , .B1( u1_u6_u2_n152 ) , .A( u1_u6_u2_n171 ) );
  INV_X1 u1_u6_u2_U16 (.A( u1_u6_u2_n156 ) , .ZN( u1_u6_u2_n171 ) );
  INV_X1 u1_u6_u2_U17 (.A( u1_u6_u2_n120 ) , .ZN( u1_u6_u2_n188 ) );
  NAND2_X1 u1_u6_u2_U18 (.A2( u1_u6_u2_n122 ) , .ZN( u1_u6_u2_n150 ) , .A1( u1_u6_u2_n152 ) );
  INV_X1 u1_u6_u2_U19 (.A( u1_u6_u2_n153 ) , .ZN( u1_u6_u2_n170 ) );
  INV_X1 u1_u6_u2_U20 (.A( u1_u6_u2_n137 ) , .ZN( u1_u6_u2_n173 ) );
  NAND2_X1 u1_u6_u2_U21 (.A1( u1_u6_u2_n132 ) , .A2( u1_u6_u2_n139 ) , .ZN( u1_u6_u2_n157 ) );
  INV_X1 u1_u6_u2_U22 (.A( u1_u6_u2_n113 ) , .ZN( u1_u6_u2_n178 ) );
  INV_X1 u1_u6_u2_U23 (.A( u1_u6_u2_n139 ) , .ZN( u1_u6_u2_n175 ) );
  INV_X1 u1_u6_u2_U24 (.A( u1_u6_u2_n155 ) , .ZN( u1_u6_u2_n181 ) );
  INV_X1 u1_u6_u2_U25 (.A( u1_u6_u2_n119 ) , .ZN( u1_u6_u2_n177 ) );
  INV_X1 u1_u6_u2_U26 (.A( u1_u6_u2_n116 ) , .ZN( u1_u6_u2_n180 ) );
  INV_X1 u1_u6_u2_U27 (.A( u1_u6_u2_n131 ) , .ZN( u1_u6_u2_n179 ) );
  INV_X1 u1_u6_u2_U28 (.A( u1_u6_u2_n154 ) , .ZN( u1_u6_u2_n176 ) );
  NAND2_X1 u1_u6_u2_U29 (.A2( u1_u6_u2_n116 ) , .A1( u1_u6_u2_n117 ) , .ZN( u1_u6_u2_n118 ) );
  NOR2_X1 u1_u6_u2_U3 (.ZN( u1_u6_u2_n121 ) , .A2( u1_u6_u2_n177 ) , .A1( u1_u6_u2_n180 ) );
  INV_X1 u1_u6_u2_U30 (.A( u1_u6_u2_n132 ) , .ZN( u1_u6_u2_n182 ) );
  INV_X1 u1_u6_u2_U31 (.A( u1_u6_u2_n158 ) , .ZN( u1_u6_u2_n183 ) );
  OAI21_X1 u1_u6_u2_U32 (.A( u1_u6_u2_n156 ) , .B1( u1_u6_u2_n157 ) , .ZN( u1_u6_u2_n158 ) , .B2( u1_u6_u2_n179 ) );
  NOR2_X1 u1_u6_u2_U33 (.ZN( u1_u6_u2_n156 ) , .A1( u1_u6_u2_n166 ) , .A2( u1_u6_u2_n169 ) );
  NOR2_X1 u1_u6_u2_U34 (.A2( u1_u6_u2_n114 ) , .ZN( u1_u6_u2_n137 ) , .A1( u1_u6_u2_n140 ) );
  NOR2_X1 u1_u6_u2_U35 (.A2( u1_u6_u2_n138 ) , .ZN( u1_u6_u2_n153 ) , .A1( u1_u6_u2_n156 ) );
  AOI211_X1 u1_u6_u2_U36 (.ZN( u1_u6_u2_n130 ) , .C1( u1_u6_u2_n138 ) , .C2( u1_u6_u2_n179 ) , .B( u1_u6_u2_n96 ) , .A( u1_u6_u2_n97 ) );
  OAI22_X1 u1_u6_u2_U37 (.B1( u1_u6_u2_n133 ) , .A2( u1_u6_u2_n137 ) , .A1( u1_u6_u2_n152 ) , .B2( u1_u6_u2_n168 ) , .ZN( u1_u6_u2_n97 ) );
  OAI221_X1 u1_u6_u2_U38 (.B1( u1_u6_u2_n113 ) , .C1( u1_u6_u2_n132 ) , .A( u1_u6_u2_n149 ) , .B2( u1_u6_u2_n171 ) , .C2( u1_u6_u2_n172 ) , .ZN( u1_u6_u2_n96 ) );
  OAI221_X1 u1_u6_u2_U39 (.A( u1_u6_u2_n115 ) , .C2( u1_u6_u2_n123 ) , .B2( u1_u6_u2_n143 ) , .B1( u1_u6_u2_n153 ) , .ZN( u1_u6_u2_n163 ) , .C1( u1_u6_u2_n168 ) );
  INV_X1 u1_u6_u2_U4 (.A( u1_u6_u2_n134 ) , .ZN( u1_u6_u2_n185 ) );
  OAI21_X1 u1_u6_u2_U40 (.A( u1_u6_u2_n114 ) , .ZN( u1_u6_u2_n115 ) , .B1( u1_u6_u2_n176 ) , .B2( u1_u6_u2_n178 ) );
  OAI221_X1 u1_u6_u2_U41 (.A( u1_u6_u2_n135 ) , .B2( u1_u6_u2_n136 ) , .B1( u1_u6_u2_n137 ) , .ZN( u1_u6_u2_n162 ) , .C2( u1_u6_u2_n167 ) , .C1( u1_u6_u2_n185 ) );
  AND3_X1 u1_u6_u2_U42 (.A3( u1_u6_u2_n131 ) , .A2( u1_u6_u2_n132 ) , .A1( u1_u6_u2_n133 ) , .ZN( u1_u6_u2_n136 ) );
  AOI22_X1 u1_u6_u2_U43 (.ZN( u1_u6_u2_n135 ) , .B1( u1_u6_u2_n140 ) , .A1( u1_u6_u2_n156 ) , .B2( u1_u6_u2_n180 ) , .A2( u1_u6_u2_n188 ) );
  AOI21_X1 u1_u6_u2_U44 (.ZN( u1_u6_u2_n149 ) , .B1( u1_u6_u2_n173 ) , .B2( u1_u6_u2_n188 ) , .A( u1_u6_u2_n95 ) );
  AND3_X1 u1_u6_u2_U45 (.A2( u1_u6_u2_n100 ) , .A1( u1_u6_u2_n104 ) , .A3( u1_u6_u2_n156 ) , .ZN( u1_u6_u2_n95 ) );
  OAI21_X1 u1_u6_u2_U46 (.A( u1_u6_u2_n101 ) , .B2( u1_u6_u2_n121 ) , .B1( u1_u6_u2_n153 ) , .ZN( u1_u6_u2_n164 ) );
  NAND2_X1 u1_u6_u2_U47 (.A2( u1_u6_u2_n100 ) , .A1( u1_u6_u2_n107 ) , .ZN( u1_u6_u2_n155 ) );
  NAND2_X1 u1_u6_u2_U48 (.A2( u1_u6_u2_n105 ) , .A1( u1_u6_u2_n108 ) , .ZN( u1_u6_u2_n143 ) );
  NAND2_X1 u1_u6_u2_U49 (.A1( u1_u6_u2_n104 ) , .A2( u1_u6_u2_n106 ) , .ZN( u1_u6_u2_n152 ) );
  NOR4_X1 u1_u6_u2_U5 (.A4( u1_u6_u2_n124 ) , .A3( u1_u6_u2_n125 ) , .A2( u1_u6_u2_n126 ) , .A1( u1_u6_u2_n127 ) , .ZN( u1_u6_u2_n128 ) );
  NAND2_X1 u1_u6_u2_U50 (.A1( u1_u6_u2_n100 ) , .A2( u1_u6_u2_n105 ) , .ZN( u1_u6_u2_n132 ) );
  INV_X1 u1_u6_u2_U51 (.A( u1_u6_u2_n140 ) , .ZN( u1_u6_u2_n168 ) );
  INV_X1 u1_u6_u2_U52 (.A( u1_u6_u2_n138 ) , .ZN( u1_u6_u2_n167 ) );
  OAI21_X1 u1_u6_u2_U53 (.A( u1_u6_u2_n141 ) , .B2( u1_u6_u2_n142 ) , .ZN( u1_u6_u2_n146 ) , .B1( u1_u6_u2_n153 ) );
  OAI21_X1 u1_u6_u2_U54 (.A( u1_u6_u2_n140 ) , .ZN( u1_u6_u2_n141 ) , .B1( u1_u6_u2_n176 ) , .B2( u1_u6_u2_n177 ) );
  NOR3_X1 u1_u6_u2_U55 (.ZN( u1_u6_u2_n142 ) , .A3( u1_u6_u2_n175 ) , .A2( u1_u6_u2_n178 ) , .A1( u1_u6_u2_n181 ) );
  NAND2_X1 u1_u6_u2_U56 (.A1( u1_u6_u2_n102 ) , .A2( u1_u6_u2_n106 ) , .ZN( u1_u6_u2_n113 ) );
  NAND2_X1 u1_u6_u2_U57 (.A1( u1_u6_u2_n106 ) , .A2( u1_u6_u2_n107 ) , .ZN( u1_u6_u2_n131 ) );
  NAND2_X1 u1_u6_u2_U58 (.A1( u1_u6_u2_n103 ) , .A2( u1_u6_u2_n107 ) , .ZN( u1_u6_u2_n139 ) );
  NAND2_X1 u1_u6_u2_U59 (.A1( u1_u6_u2_n103 ) , .A2( u1_u6_u2_n105 ) , .ZN( u1_u6_u2_n133 ) );
  AOI21_X1 u1_u6_u2_U6 (.B2( u1_u6_u2_n119 ) , .ZN( u1_u6_u2_n127 ) , .A( u1_u6_u2_n137 ) , .B1( u1_u6_u2_n155 ) );
  NAND2_X1 u1_u6_u2_U60 (.A1( u1_u6_u2_n102 ) , .A2( u1_u6_u2_n103 ) , .ZN( u1_u6_u2_n154 ) );
  NAND2_X1 u1_u6_u2_U61 (.A2( u1_u6_u2_n103 ) , .A1( u1_u6_u2_n104 ) , .ZN( u1_u6_u2_n119 ) );
  NAND2_X1 u1_u6_u2_U62 (.A2( u1_u6_u2_n107 ) , .A1( u1_u6_u2_n108 ) , .ZN( u1_u6_u2_n123 ) );
  NAND2_X1 u1_u6_u2_U63 (.A1( u1_u6_u2_n104 ) , .A2( u1_u6_u2_n108 ) , .ZN( u1_u6_u2_n122 ) );
  INV_X1 u1_u6_u2_U64 (.A( u1_u6_u2_n114 ) , .ZN( u1_u6_u2_n172 ) );
  NAND2_X1 u1_u6_u2_U65 (.A2( u1_u6_u2_n100 ) , .A1( u1_u6_u2_n102 ) , .ZN( u1_u6_u2_n116 ) );
  NAND2_X1 u1_u6_u2_U66 (.A1( u1_u6_u2_n102 ) , .A2( u1_u6_u2_n108 ) , .ZN( u1_u6_u2_n120 ) );
  NAND2_X1 u1_u6_u2_U67 (.A2( u1_u6_u2_n105 ) , .A1( u1_u6_u2_n106 ) , .ZN( u1_u6_u2_n117 ) );
  INV_X1 u1_u6_u2_U68 (.ZN( u1_u6_u2_n187 ) , .A( u1_u6_u2_n99 ) );
  OAI21_X1 u1_u6_u2_U69 (.B1( u1_u6_u2_n137 ) , .B2( u1_u6_u2_n143 ) , .A( u1_u6_u2_n98 ) , .ZN( u1_u6_u2_n99 ) );
  AOI21_X1 u1_u6_u2_U7 (.ZN( u1_u6_u2_n124 ) , .B1( u1_u6_u2_n131 ) , .B2( u1_u6_u2_n143 ) , .A( u1_u6_u2_n172 ) );
  NOR2_X1 u1_u6_u2_U70 (.A2( u1_u6_X_16 ) , .ZN( u1_u6_u2_n140 ) , .A1( u1_u6_u2_n166 ) );
  NOR2_X1 u1_u6_u2_U71 (.A2( u1_u6_X_13 ) , .A1( u1_u6_X_14 ) , .ZN( u1_u6_u2_n100 ) );
  NOR2_X1 u1_u6_u2_U72 (.A2( u1_u6_X_16 ) , .A1( u1_u6_X_17 ) , .ZN( u1_u6_u2_n138 ) );
  NOR2_X1 u1_u6_u2_U73 (.A2( u1_u6_X_15 ) , .A1( u1_u6_X_18 ) , .ZN( u1_u6_u2_n104 ) );
  NOR2_X1 u1_u6_u2_U74 (.A2( u1_u6_X_14 ) , .ZN( u1_u6_u2_n103 ) , .A1( u1_u6_u2_n174 ) );
  NOR2_X1 u1_u6_u2_U75 (.A2( u1_u6_X_15 ) , .ZN( u1_u6_u2_n102 ) , .A1( u1_u6_u2_n165 ) );
  NOR2_X1 u1_u6_u2_U76 (.A2( u1_u6_X_17 ) , .ZN( u1_u6_u2_n114 ) , .A1( u1_u6_u2_n169 ) );
  AND2_X1 u1_u6_u2_U77 (.A1( u1_u6_X_15 ) , .ZN( u1_u6_u2_n105 ) , .A2( u1_u6_u2_n165 ) );
  AND2_X1 u1_u6_u2_U78 (.A2( u1_u6_X_15 ) , .A1( u1_u6_X_18 ) , .ZN( u1_u6_u2_n107 ) );
  AND2_X1 u1_u6_u2_U79 (.A1( u1_u6_X_14 ) , .ZN( u1_u6_u2_n106 ) , .A2( u1_u6_u2_n174 ) );
  AOI21_X1 u1_u6_u2_U8 (.B2( u1_u6_u2_n120 ) , .B1( u1_u6_u2_n121 ) , .ZN( u1_u6_u2_n126 ) , .A( u1_u6_u2_n167 ) );
  AND2_X1 u1_u6_u2_U80 (.A1( u1_u6_X_13 ) , .A2( u1_u6_X_14 ) , .ZN( u1_u6_u2_n108 ) );
  INV_X1 u1_u6_u2_U81 (.A( u1_u6_X_16 ) , .ZN( u1_u6_u2_n169 ) );
  INV_X1 u1_u6_u2_U82 (.A( u1_u6_X_17 ) , .ZN( u1_u6_u2_n166 ) );
  INV_X1 u1_u6_u2_U83 (.A( u1_u6_X_13 ) , .ZN( u1_u6_u2_n174 ) );
  INV_X1 u1_u6_u2_U84 (.A( u1_u6_X_18 ) , .ZN( u1_u6_u2_n165 ) );
  NAND4_X1 u1_u6_u2_U85 (.ZN( u1_out6_16 ) , .A4( u1_u6_u2_n128 ) , .A3( u1_u6_u2_n129 ) , .A1( u1_u6_u2_n130 ) , .A2( u1_u6_u2_n186 ) );
  AOI22_X1 u1_u6_u2_U86 (.A2( u1_u6_u2_n118 ) , .ZN( u1_u6_u2_n129 ) , .A1( u1_u6_u2_n140 ) , .B1( u1_u6_u2_n157 ) , .B2( u1_u6_u2_n170 ) );
  INV_X1 u1_u6_u2_U87 (.A( u1_u6_u2_n163 ) , .ZN( u1_u6_u2_n186 ) );
  NAND4_X1 u1_u6_u2_U88 (.ZN( u1_out6_24 ) , .A4( u1_u6_u2_n111 ) , .A3( u1_u6_u2_n112 ) , .A1( u1_u6_u2_n130 ) , .A2( u1_u6_u2_n187 ) );
  AOI221_X1 u1_u6_u2_U89 (.A( u1_u6_u2_n109 ) , .B1( u1_u6_u2_n110 ) , .ZN( u1_u6_u2_n111 ) , .C1( u1_u6_u2_n134 ) , .C2( u1_u6_u2_n170 ) , .B2( u1_u6_u2_n173 ) );
  OAI22_X1 u1_u6_u2_U9 (.ZN( u1_u6_u2_n109 ) , .A2( u1_u6_u2_n113 ) , .B2( u1_u6_u2_n133 ) , .B1( u1_u6_u2_n167 ) , .A1( u1_u6_u2_n168 ) );
  AOI21_X1 u1_u6_u2_U90 (.ZN( u1_u6_u2_n112 ) , .B2( u1_u6_u2_n156 ) , .A( u1_u6_u2_n164 ) , .B1( u1_u6_u2_n181 ) );
  NAND4_X1 u1_u6_u2_U91 (.ZN( u1_out6_30 ) , .A4( u1_u6_u2_n147 ) , .A3( u1_u6_u2_n148 ) , .A2( u1_u6_u2_n149 ) , .A1( u1_u6_u2_n187 ) );
  AOI21_X1 u1_u6_u2_U92 (.B2( u1_u6_u2_n138 ) , .ZN( u1_u6_u2_n148 ) , .A( u1_u6_u2_n162 ) , .B1( u1_u6_u2_n182 ) );
  NOR3_X1 u1_u6_u2_U93 (.A3( u1_u6_u2_n144 ) , .A2( u1_u6_u2_n145 ) , .A1( u1_u6_u2_n146 ) , .ZN( u1_u6_u2_n147 ) );
  OR4_X1 u1_u6_u2_U94 (.ZN( u1_out6_6 ) , .A4( u1_u6_u2_n161 ) , .A3( u1_u6_u2_n162 ) , .A2( u1_u6_u2_n163 ) , .A1( u1_u6_u2_n164 ) );
  OR3_X1 u1_u6_u2_U95 (.A2( u1_u6_u2_n159 ) , .A1( u1_u6_u2_n160 ) , .ZN( u1_u6_u2_n161 ) , .A3( u1_u6_u2_n183 ) );
  AOI21_X1 u1_u6_u2_U96 (.B2( u1_u6_u2_n154 ) , .B1( u1_u6_u2_n155 ) , .ZN( u1_u6_u2_n159 ) , .A( u1_u6_u2_n167 ) );
  NAND3_X1 u1_u6_u2_U97 (.A2( u1_u6_u2_n117 ) , .A1( u1_u6_u2_n122 ) , .A3( u1_u6_u2_n123 ) , .ZN( u1_u6_u2_n134 ) );
  NAND3_X1 u1_u6_u2_U98 (.ZN( u1_u6_u2_n110 ) , .A2( u1_u6_u2_n131 ) , .A3( u1_u6_u2_n139 ) , .A1( u1_u6_u2_n154 ) );
  NAND3_X1 u1_u6_u2_U99 (.A2( u1_u6_u2_n100 ) , .ZN( u1_u6_u2_n101 ) , .A1( u1_u6_u2_n104 ) , .A3( u1_u6_u2_n114 ) );
  AOI21_X1 u1_u6_u6_U10 (.ZN( u1_u6_u6_n106 ) , .A( u1_u6_u6_n142 ) , .B2( u1_u6_u6_n159 ) , .B1( u1_u6_u6_n164 ) );
  INV_X1 u1_u6_u6_U11 (.A( u1_u6_u6_n155 ) , .ZN( u1_u6_u6_n161 ) );
  INV_X1 u1_u6_u6_U12 (.A( u1_u6_u6_n128 ) , .ZN( u1_u6_u6_n164 ) );
  NAND2_X1 u1_u6_u6_U13 (.ZN( u1_u6_u6_n110 ) , .A1( u1_u6_u6_n122 ) , .A2( u1_u6_u6_n129 ) );
  NAND2_X1 u1_u6_u6_U14 (.ZN( u1_u6_u6_n124 ) , .A2( u1_u6_u6_n146 ) , .A1( u1_u6_u6_n148 ) );
  INV_X1 u1_u6_u6_U15 (.A( u1_u6_u6_n132 ) , .ZN( u1_u6_u6_n171 ) );
  AND2_X1 u1_u6_u6_U16 (.A1( u1_u6_u6_n100 ) , .ZN( u1_u6_u6_n130 ) , .A2( u1_u6_u6_n147 ) );
  INV_X1 u1_u6_u6_U17 (.A( u1_u6_u6_n127 ) , .ZN( u1_u6_u6_n173 ) );
  INV_X1 u1_u6_u6_U18 (.A( u1_u6_u6_n121 ) , .ZN( u1_u6_u6_n167 ) );
  INV_X1 u1_u6_u6_U19 (.A( u1_u6_u6_n100 ) , .ZN( u1_u6_u6_n169 ) );
  INV_X1 u1_u6_u6_U20 (.A( u1_u6_u6_n123 ) , .ZN( u1_u6_u6_n170 ) );
  INV_X1 u1_u6_u6_U21 (.A( u1_u6_u6_n113 ) , .ZN( u1_u6_u6_n168 ) );
  AND2_X1 u1_u6_u6_U22 (.A1( u1_u6_u6_n107 ) , .A2( u1_u6_u6_n119 ) , .ZN( u1_u6_u6_n133 ) );
  AND2_X1 u1_u6_u6_U23 (.A2( u1_u6_u6_n121 ) , .A1( u1_u6_u6_n122 ) , .ZN( u1_u6_u6_n131 ) );
  AND3_X1 u1_u6_u6_U24 (.ZN( u1_u6_u6_n120 ) , .A2( u1_u6_u6_n127 ) , .A1( u1_u6_u6_n132 ) , .A3( u1_u6_u6_n145 ) );
  INV_X1 u1_u6_u6_U25 (.A( u1_u6_u6_n146 ) , .ZN( u1_u6_u6_n163 ) );
  AOI222_X1 u1_u6_u6_U26 (.ZN( u1_u6_u6_n114 ) , .A1( u1_u6_u6_n118 ) , .A2( u1_u6_u6_n126 ) , .B2( u1_u6_u6_n151 ) , .C2( u1_u6_u6_n159 ) , .C1( u1_u6_u6_n168 ) , .B1( u1_u6_u6_n169 ) );
  NOR2_X1 u1_u6_u6_U27 (.A1( u1_u6_u6_n162 ) , .A2( u1_u6_u6_n165 ) , .ZN( u1_u6_u6_n98 ) );
  AOI211_X1 u1_u6_u6_U28 (.B( u1_u6_u6_n149 ) , .A( u1_u6_u6_n150 ) , .C2( u1_u6_u6_n151 ) , .C1( u1_u6_u6_n152 ) , .ZN( u1_u6_u6_n153 ) );
  AOI21_X1 u1_u6_u6_U29 (.B2( u1_u6_u6_n147 ) , .B1( u1_u6_u6_n148 ) , .ZN( u1_u6_u6_n149 ) , .A( u1_u6_u6_n158 ) );
  INV_X1 u1_u6_u6_U3 (.A( u1_u6_u6_n110 ) , .ZN( u1_u6_u6_n166 ) );
  AOI21_X1 u1_u6_u6_U30 (.A( u1_u6_u6_n144 ) , .B2( u1_u6_u6_n145 ) , .B1( u1_u6_u6_n146 ) , .ZN( u1_u6_u6_n150 ) );
  NAND2_X1 u1_u6_u6_U31 (.A2( u1_u6_u6_n143 ) , .ZN( u1_u6_u6_n152 ) , .A1( u1_u6_u6_n166 ) );
  NAND2_X1 u1_u6_u6_U32 (.A1( u1_u6_u6_n144 ) , .ZN( u1_u6_u6_n151 ) , .A2( u1_u6_u6_n158 ) );
  NAND2_X1 u1_u6_u6_U33 (.ZN( u1_u6_u6_n132 ) , .A1( u1_u6_u6_n91 ) , .A2( u1_u6_u6_n97 ) );
  AOI22_X1 u1_u6_u6_U34 (.B2( u1_u6_u6_n110 ) , .B1( u1_u6_u6_n111 ) , .A1( u1_u6_u6_n112 ) , .ZN( u1_u6_u6_n115 ) , .A2( u1_u6_u6_n161 ) );
  NAND4_X1 u1_u6_u6_U35 (.A3( u1_u6_u6_n109 ) , .ZN( u1_u6_u6_n112 ) , .A4( u1_u6_u6_n132 ) , .A2( u1_u6_u6_n147 ) , .A1( u1_u6_u6_n166 ) );
  NOR2_X1 u1_u6_u6_U36 (.ZN( u1_u6_u6_n109 ) , .A1( u1_u6_u6_n170 ) , .A2( u1_u6_u6_n173 ) );
  NOR2_X1 u1_u6_u6_U37 (.A2( u1_u6_u6_n126 ) , .ZN( u1_u6_u6_n155 ) , .A1( u1_u6_u6_n160 ) );
  NAND2_X1 u1_u6_u6_U38 (.ZN( u1_u6_u6_n146 ) , .A2( u1_u6_u6_n94 ) , .A1( u1_u6_u6_n99 ) );
  AOI211_X1 u1_u6_u6_U39 (.B( u1_u6_u6_n134 ) , .A( u1_u6_u6_n135 ) , .C1( u1_u6_u6_n136 ) , .ZN( u1_u6_u6_n137 ) , .C2( u1_u6_u6_n151 ) );
  AOI22_X1 u1_u6_u6_U4 (.B2( u1_u6_u6_n101 ) , .A1( u1_u6_u6_n102 ) , .ZN( u1_u6_u6_n103 ) , .B1( u1_u6_u6_n160 ) , .A2( u1_u6_u6_n161 ) );
  NAND4_X1 u1_u6_u6_U40 (.A4( u1_u6_u6_n127 ) , .A3( u1_u6_u6_n128 ) , .A2( u1_u6_u6_n129 ) , .A1( u1_u6_u6_n130 ) , .ZN( u1_u6_u6_n136 ) );
  AOI21_X1 u1_u6_u6_U41 (.B2( u1_u6_u6_n132 ) , .B1( u1_u6_u6_n133 ) , .ZN( u1_u6_u6_n134 ) , .A( u1_u6_u6_n158 ) );
  AOI21_X1 u1_u6_u6_U42 (.B1( u1_u6_u6_n131 ) , .ZN( u1_u6_u6_n135 ) , .A( u1_u6_u6_n144 ) , .B2( u1_u6_u6_n146 ) );
  INV_X1 u1_u6_u6_U43 (.A( u1_u6_u6_n111 ) , .ZN( u1_u6_u6_n158 ) );
  NAND2_X1 u1_u6_u6_U44 (.ZN( u1_u6_u6_n127 ) , .A1( u1_u6_u6_n91 ) , .A2( u1_u6_u6_n92 ) );
  NAND2_X1 u1_u6_u6_U45 (.ZN( u1_u6_u6_n129 ) , .A2( u1_u6_u6_n95 ) , .A1( u1_u6_u6_n96 ) );
  INV_X1 u1_u6_u6_U46 (.A( u1_u6_u6_n144 ) , .ZN( u1_u6_u6_n159 ) );
  NAND2_X1 u1_u6_u6_U47 (.ZN( u1_u6_u6_n145 ) , .A2( u1_u6_u6_n97 ) , .A1( u1_u6_u6_n98 ) );
  NAND2_X1 u1_u6_u6_U48 (.ZN( u1_u6_u6_n148 ) , .A2( u1_u6_u6_n92 ) , .A1( u1_u6_u6_n94 ) );
  NAND2_X1 u1_u6_u6_U49 (.ZN( u1_u6_u6_n108 ) , .A2( u1_u6_u6_n139 ) , .A1( u1_u6_u6_n144 ) );
  NOR2_X1 u1_u6_u6_U5 (.A1( u1_u6_u6_n118 ) , .ZN( u1_u6_u6_n143 ) , .A2( u1_u6_u6_n168 ) );
  NAND2_X1 u1_u6_u6_U50 (.ZN( u1_u6_u6_n121 ) , .A2( u1_u6_u6_n95 ) , .A1( u1_u6_u6_n97 ) );
  NAND2_X1 u1_u6_u6_U51 (.ZN( u1_u6_u6_n107 ) , .A2( u1_u6_u6_n92 ) , .A1( u1_u6_u6_n95 ) );
  AND2_X1 u1_u6_u6_U52 (.ZN( u1_u6_u6_n118 ) , .A2( u1_u6_u6_n91 ) , .A1( u1_u6_u6_n99 ) );
  NAND2_X1 u1_u6_u6_U53 (.ZN( u1_u6_u6_n147 ) , .A2( u1_u6_u6_n98 ) , .A1( u1_u6_u6_n99 ) );
  NAND2_X1 u1_u6_u6_U54 (.ZN( u1_u6_u6_n128 ) , .A1( u1_u6_u6_n94 ) , .A2( u1_u6_u6_n96 ) );
  NAND2_X1 u1_u6_u6_U55 (.ZN( u1_u6_u6_n119 ) , .A2( u1_u6_u6_n95 ) , .A1( u1_u6_u6_n99 ) );
  NAND2_X1 u1_u6_u6_U56 (.ZN( u1_u6_u6_n123 ) , .A2( u1_u6_u6_n91 ) , .A1( u1_u6_u6_n96 ) );
  NAND2_X1 u1_u6_u6_U57 (.ZN( u1_u6_u6_n100 ) , .A2( u1_u6_u6_n92 ) , .A1( u1_u6_u6_n98 ) );
  NAND2_X1 u1_u6_u6_U58 (.ZN( u1_u6_u6_n122 ) , .A1( u1_u6_u6_n94 ) , .A2( u1_u6_u6_n97 ) );
  INV_X1 u1_u6_u6_U59 (.A( u1_u6_u6_n139 ) , .ZN( u1_u6_u6_n160 ) );
  AOI21_X1 u1_u6_u6_U6 (.B1( u1_u6_u6_n107 ) , .B2( u1_u6_u6_n132 ) , .A( u1_u6_u6_n158 ) , .ZN( u1_u6_u6_n88 ) );
  NAND2_X1 u1_u6_u6_U60 (.ZN( u1_u6_u6_n113 ) , .A1( u1_u6_u6_n96 ) , .A2( u1_u6_u6_n98 ) );
  NOR2_X1 u1_u6_u6_U61 (.A2( u1_u6_X_40 ) , .A1( u1_u6_X_41 ) , .ZN( u1_u6_u6_n126 ) );
  NOR2_X1 u1_u6_u6_U62 (.A2( u1_u6_X_39 ) , .A1( u1_u6_X_42 ) , .ZN( u1_u6_u6_n92 ) );
  NOR2_X1 u1_u6_u6_U63 (.A2( u1_u6_X_39 ) , .A1( u1_u6_u6_n156 ) , .ZN( u1_u6_u6_n97 ) );
  NOR2_X1 u1_u6_u6_U64 (.A2( u1_u6_X_38 ) , .A1( u1_u6_u6_n165 ) , .ZN( u1_u6_u6_n95 ) );
  NOR2_X1 u1_u6_u6_U65 (.A2( u1_u6_X_41 ) , .ZN( u1_u6_u6_n111 ) , .A1( u1_u6_u6_n157 ) );
  NOR2_X1 u1_u6_u6_U66 (.A2( u1_u6_X_37 ) , .A1( u1_u6_u6_n162 ) , .ZN( u1_u6_u6_n94 ) );
  NOR2_X1 u1_u6_u6_U67 (.A2( u1_u6_X_37 ) , .A1( u1_u6_X_38 ) , .ZN( u1_u6_u6_n91 ) );
  NAND2_X1 u1_u6_u6_U68 (.A1( u1_u6_X_41 ) , .ZN( u1_u6_u6_n144 ) , .A2( u1_u6_u6_n157 ) );
  NAND2_X1 u1_u6_u6_U69 (.A2( u1_u6_X_40 ) , .A1( u1_u6_X_41 ) , .ZN( u1_u6_u6_n139 ) );
  OAI21_X1 u1_u6_u6_U7 (.A( u1_u6_u6_n159 ) , .B1( u1_u6_u6_n169 ) , .B2( u1_u6_u6_n173 ) , .ZN( u1_u6_u6_n90 ) );
  AND2_X1 u1_u6_u6_U70 (.A1( u1_u6_X_39 ) , .A2( u1_u6_u6_n156 ) , .ZN( u1_u6_u6_n96 ) );
  AND2_X1 u1_u6_u6_U71 (.A1( u1_u6_X_39 ) , .A2( u1_u6_X_42 ) , .ZN( u1_u6_u6_n99 ) );
  INV_X1 u1_u6_u6_U72 (.A( u1_u6_X_40 ) , .ZN( u1_u6_u6_n157 ) );
  INV_X1 u1_u6_u6_U73 (.A( u1_u6_X_37 ) , .ZN( u1_u6_u6_n165 ) );
  INV_X1 u1_u6_u6_U74 (.A( u1_u6_X_38 ) , .ZN( u1_u6_u6_n162 ) );
  INV_X1 u1_u6_u6_U75 (.A( u1_u6_X_42 ) , .ZN( u1_u6_u6_n156 ) );
  NAND4_X1 u1_u6_u6_U76 (.ZN( u1_out6_12 ) , .A4( u1_u6_u6_n114 ) , .A3( u1_u6_u6_n115 ) , .A2( u1_u6_u6_n116 ) , .A1( u1_u6_u6_n117 ) );
  OAI22_X1 u1_u6_u6_U77 (.B2( u1_u6_u6_n111 ) , .ZN( u1_u6_u6_n116 ) , .B1( u1_u6_u6_n126 ) , .A2( u1_u6_u6_n164 ) , .A1( u1_u6_u6_n167 ) );
  OAI21_X1 u1_u6_u6_U78 (.A( u1_u6_u6_n108 ) , .ZN( u1_u6_u6_n117 ) , .B2( u1_u6_u6_n141 ) , .B1( u1_u6_u6_n163 ) );
  NAND4_X1 u1_u6_u6_U79 (.ZN( u1_out6_32 ) , .A4( u1_u6_u6_n103 ) , .A3( u1_u6_u6_n104 ) , .A2( u1_u6_u6_n105 ) , .A1( u1_u6_u6_n106 ) );
  INV_X1 u1_u6_u6_U8 (.ZN( u1_u6_u6_n172 ) , .A( u1_u6_u6_n88 ) );
  AOI22_X1 u1_u6_u6_U80 (.ZN( u1_u6_u6_n104 ) , .A1( u1_u6_u6_n111 ) , .B1( u1_u6_u6_n124 ) , .B2( u1_u6_u6_n151 ) , .A2( u1_u6_u6_n93 ) );
  AOI22_X1 u1_u6_u6_U81 (.ZN( u1_u6_u6_n105 ) , .A2( u1_u6_u6_n108 ) , .A1( u1_u6_u6_n118 ) , .B2( u1_u6_u6_n126 ) , .B1( u1_u6_u6_n171 ) );
  OAI211_X1 u1_u6_u6_U82 (.ZN( u1_out6_22 ) , .B( u1_u6_u6_n137 ) , .A( u1_u6_u6_n138 ) , .C2( u1_u6_u6_n139 ) , .C1( u1_u6_u6_n140 ) );
  AOI22_X1 u1_u6_u6_U83 (.B1( u1_u6_u6_n124 ) , .A2( u1_u6_u6_n125 ) , .A1( u1_u6_u6_n126 ) , .ZN( u1_u6_u6_n138 ) , .B2( u1_u6_u6_n161 ) );
  AND4_X1 u1_u6_u6_U84 (.A3( u1_u6_u6_n119 ) , .A1( u1_u6_u6_n120 ) , .A4( u1_u6_u6_n129 ) , .ZN( u1_u6_u6_n140 ) , .A2( u1_u6_u6_n143 ) );
  OAI211_X1 u1_u6_u6_U85 (.ZN( u1_out6_7 ) , .B( u1_u6_u6_n153 ) , .C2( u1_u6_u6_n154 ) , .C1( u1_u6_u6_n155 ) , .A( u1_u6_u6_n174 ) );
  NOR3_X1 u1_u6_u6_U86 (.A1( u1_u6_u6_n141 ) , .ZN( u1_u6_u6_n154 ) , .A3( u1_u6_u6_n164 ) , .A2( u1_u6_u6_n171 ) );
  INV_X1 u1_u6_u6_U87 (.A( u1_u6_u6_n142 ) , .ZN( u1_u6_u6_n174 ) );
  NAND3_X1 u1_u6_u6_U88 (.A2( u1_u6_u6_n123 ) , .ZN( u1_u6_u6_n125 ) , .A1( u1_u6_u6_n130 ) , .A3( u1_u6_u6_n131 ) );
  NAND3_X1 u1_u6_u6_U89 (.A3( u1_u6_u6_n133 ) , .ZN( u1_u6_u6_n141 ) , .A1( u1_u6_u6_n145 ) , .A2( u1_u6_u6_n148 ) );
  AOI22_X1 u1_u6_u6_U9 (.A2( u1_u6_u6_n151 ) , .B2( u1_u6_u6_n161 ) , .A1( u1_u6_u6_n167 ) , .B1( u1_u6_u6_n170 ) , .ZN( u1_u6_u6_n89 ) );
  NAND3_X1 u1_u6_u6_U90 (.ZN( u1_u6_u6_n101 ) , .A3( u1_u6_u6_n107 ) , .A2( u1_u6_u6_n121 ) , .A1( u1_u6_u6_n127 ) );
  NAND3_X1 u1_u6_u6_U91 (.ZN( u1_u6_u6_n102 ) , .A3( u1_u6_u6_n130 ) , .A2( u1_u6_u6_n145 ) , .A1( u1_u6_u6_n166 ) );
  NAND3_X1 u1_u6_u6_U92 (.A3( u1_u6_u6_n113 ) , .A1( u1_u6_u6_n119 ) , .A2( u1_u6_u6_n123 ) , .ZN( u1_u6_u6_n93 ) );
  NAND3_X1 u1_u6_u6_U93 (.ZN( u1_u6_u6_n142 ) , .A2( u1_u6_u6_n172 ) , .A3( u1_u6_u6_n89 ) , .A1( u1_u6_u6_n90 ) );
  AND3_X1 u1_u6_u7_U10 (.A3( u1_u6_u7_n110 ) , .A2( u1_u6_u7_n127 ) , .A1( u1_u6_u7_n132 ) , .ZN( u1_u6_u7_n92 ) );
  OAI21_X1 u1_u6_u7_U11 (.A( u1_u6_u7_n161 ) , .B1( u1_u6_u7_n168 ) , .B2( u1_u6_u7_n173 ) , .ZN( u1_u6_u7_n91 ) );
  AOI211_X1 u1_u6_u7_U12 (.A( u1_u6_u7_n117 ) , .ZN( u1_u6_u7_n118 ) , .C2( u1_u6_u7_n126 ) , .C1( u1_u6_u7_n177 ) , .B( u1_u6_u7_n180 ) );
  OAI22_X1 u1_u6_u7_U13 (.B1( u1_u6_u7_n115 ) , .ZN( u1_u6_u7_n117 ) , .A2( u1_u6_u7_n133 ) , .A1( u1_u6_u7_n137 ) , .B2( u1_u6_u7_n162 ) );
  INV_X1 u1_u6_u7_U14 (.A( u1_u6_u7_n116 ) , .ZN( u1_u6_u7_n180 ) );
  NOR3_X1 u1_u6_u7_U15 (.ZN( u1_u6_u7_n115 ) , .A3( u1_u6_u7_n145 ) , .A2( u1_u6_u7_n168 ) , .A1( u1_u6_u7_n169 ) );
  OAI211_X1 u1_u6_u7_U16 (.B( u1_u6_u7_n122 ) , .A( u1_u6_u7_n123 ) , .C2( u1_u6_u7_n124 ) , .ZN( u1_u6_u7_n154 ) , .C1( u1_u6_u7_n162 ) );
  AOI222_X1 u1_u6_u7_U17 (.ZN( u1_u6_u7_n122 ) , .C2( u1_u6_u7_n126 ) , .C1( u1_u6_u7_n145 ) , .B1( u1_u6_u7_n161 ) , .A2( u1_u6_u7_n165 ) , .B2( u1_u6_u7_n170 ) , .A1( u1_u6_u7_n176 ) );
  INV_X1 u1_u6_u7_U18 (.A( u1_u6_u7_n133 ) , .ZN( u1_u6_u7_n176 ) );
  NOR3_X1 u1_u6_u7_U19 (.A2( u1_u6_u7_n134 ) , .A1( u1_u6_u7_n135 ) , .ZN( u1_u6_u7_n136 ) , .A3( u1_u6_u7_n171 ) );
  NOR2_X1 u1_u6_u7_U20 (.A1( u1_u6_u7_n130 ) , .A2( u1_u6_u7_n134 ) , .ZN( u1_u6_u7_n153 ) );
  INV_X1 u1_u6_u7_U21 (.A( u1_u6_u7_n101 ) , .ZN( u1_u6_u7_n165 ) );
  NOR2_X1 u1_u6_u7_U22 (.ZN( u1_u6_u7_n111 ) , .A2( u1_u6_u7_n134 ) , .A1( u1_u6_u7_n169 ) );
  AOI21_X1 u1_u6_u7_U23 (.ZN( u1_u6_u7_n104 ) , .B2( u1_u6_u7_n112 ) , .B1( u1_u6_u7_n127 ) , .A( u1_u6_u7_n164 ) );
  AOI21_X1 u1_u6_u7_U24 (.ZN( u1_u6_u7_n106 ) , .B1( u1_u6_u7_n133 ) , .B2( u1_u6_u7_n146 ) , .A( u1_u6_u7_n162 ) );
  AOI21_X1 u1_u6_u7_U25 (.A( u1_u6_u7_n101 ) , .ZN( u1_u6_u7_n107 ) , .B2( u1_u6_u7_n128 ) , .B1( u1_u6_u7_n175 ) );
  INV_X1 u1_u6_u7_U26 (.A( u1_u6_u7_n138 ) , .ZN( u1_u6_u7_n171 ) );
  INV_X1 u1_u6_u7_U27 (.A( u1_u6_u7_n131 ) , .ZN( u1_u6_u7_n177 ) );
  INV_X1 u1_u6_u7_U28 (.A( u1_u6_u7_n110 ) , .ZN( u1_u6_u7_n174 ) );
  NAND2_X1 u1_u6_u7_U29 (.A1( u1_u6_u7_n129 ) , .A2( u1_u6_u7_n132 ) , .ZN( u1_u6_u7_n149 ) );
  OAI21_X1 u1_u6_u7_U3 (.ZN( u1_u6_u7_n159 ) , .A( u1_u6_u7_n165 ) , .B2( u1_u6_u7_n171 ) , .B1( u1_u6_u7_n174 ) );
  NAND2_X1 u1_u6_u7_U30 (.A1( u1_u6_u7_n113 ) , .A2( u1_u6_u7_n124 ) , .ZN( u1_u6_u7_n130 ) );
  INV_X1 u1_u6_u7_U31 (.A( u1_u6_u7_n112 ) , .ZN( u1_u6_u7_n173 ) );
  INV_X1 u1_u6_u7_U32 (.A( u1_u6_u7_n128 ) , .ZN( u1_u6_u7_n168 ) );
  INV_X1 u1_u6_u7_U33 (.A( u1_u6_u7_n148 ) , .ZN( u1_u6_u7_n169 ) );
  INV_X1 u1_u6_u7_U34 (.A( u1_u6_u7_n127 ) , .ZN( u1_u6_u7_n179 ) );
  NOR2_X1 u1_u6_u7_U35 (.ZN( u1_u6_u7_n101 ) , .A2( u1_u6_u7_n150 ) , .A1( u1_u6_u7_n156 ) );
  AOI211_X1 u1_u6_u7_U36 (.B( u1_u6_u7_n154 ) , .A( u1_u6_u7_n155 ) , .C1( u1_u6_u7_n156 ) , .ZN( u1_u6_u7_n157 ) , .C2( u1_u6_u7_n172 ) );
  INV_X1 u1_u6_u7_U37 (.A( u1_u6_u7_n153 ) , .ZN( u1_u6_u7_n172 ) );
  AOI211_X1 u1_u6_u7_U38 (.B( u1_u6_u7_n139 ) , .A( u1_u6_u7_n140 ) , .C2( u1_u6_u7_n141 ) , .ZN( u1_u6_u7_n142 ) , .C1( u1_u6_u7_n156 ) );
  NAND4_X1 u1_u6_u7_U39 (.A3( u1_u6_u7_n127 ) , .A2( u1_u6_u7_n128 ) , .A1( u1_u6_u7_n129 ) , .ZN( u1_u6_u7_n141 ) , .A4( u1_u6_u7_n147 ) );
  INV_X1 u1_u6_u7_U4 (.A( u1_u6_u7_n111 ) , .ZN( u1_u6_u7_n170 ) );
  AOI21_X1 u1_u6_u7_U40 (.A( u1_u6_u7_n137 ) , .B1( u1_u6_u7_n138 ) , .ZN( u1_u6_u7_n139 ) , .B2( u1_u6_u7_n146 ) );
  OAI22_X1 u1_u6_u7_U41 (.B1( u1_u6_u7_n136 ) , .ZN( u1_u6_u7_n140 ) , .A1( u1_u6_u7_n153 ) , .B2( u1_u6_u7_n162 ) , .A2( u1_u6_u7_n164 ) );
  AOI21_X1 u1_u6_u7_U42 (.ZN( u1_u6_u7_n123 ) , .B1( u1_u6_u7_n165 ) , .B2( u1_u6_u7_n177 ) , .A( u1_u6_u7_n97 ) );
  AOI21_X1 u1_u6_u7_U43 (.B2( u1_u6_u7_n113 ) , .B1( u1_u6_u7_n124 ) , .A( u1_u6_u7_n125 ) , .ZN( u1_u6_u7_n97 ) );
  INV_X1 u1_u6_u7_U44 (.A( u1_u6_u7_n125 ) , .ZN( u1_u6_u7_n161 ) );
  INV_X1 u1_u6_u7_U45 (.A( u1_u6_u7_n152 ) , .ZN( u1_u6_u7_n162 ) );
  AOI22_X1 u1_u6_u7_U46 (.A2( u1_u6_u7_n114 ) , .ZN( u1_u6_u7_n119 ) , .B1( u1_u6_u7_n130 ) , .A1( u1_u6_u7_n156 ) , .B2( u1_u6_u7_n165 ) );
  NAND2_X1 u1_u6_u7_U47 (.A2( u1_u6_u7_n112 ) , .ZN( u1_u6_u7_n114 ) , .A1( u1_u6_u7_n175 ) );
  AND2_X1 u1_u6_u7_U48 (.ZN( u1_u6_u7_n145 ) , .A2( u1_u6_u7_n98 ) , .A1( u1_u6_u7_n99 ) );
  NOR2_X1 u1_u6_u7_U49 (.ZN( u1_u6_u7_n137 ) , .A1( u1_u6_u7_n150 ) , .A2( u1_u6_u7_n161 ) );
  INV_X1 u1_u6_u7_U5 (.A( u1_u6_u7_n149 ) , .ZN( u1_u6_u7_n175 ) );
  AOI21_X1 u1_u6_u7_U50 (.ZN( u1_u6_u7_n105 ) , .B2( u1_u6_u7_n110 ) , .A( u1_u6_u7_n125 ) , .B1( u1_u6_u7_n147 ) );
  NAND2_X1 u1_u6_u7_U51 (.ZN( u1_u6_u7_n146 ) , .A1( u1_u6_u7_n95 ) , .A2( u1_u6_u7_n98 ) );
  NAND2_X1 u1_u6_u7_U52 (.A2( u1_u6_u7_n103 ) , .ZN( u1_u6_u7_n147 ) , .A1( u1_u6_u7_n93 ) );
  NAND2_X1 u1_u6_u7_U53 (.A1( u1_u6_u7_n103 ) , .ZN( u1_u6_u7_n127 ) , .A2( u1_u6_u7_n99 ) );
  OR2_X1 u1_u6_u7_U54 (.ZN( u1_u6_u7_n126 ) , .A2( u1_u6_u7_n152 ) , .A1( u1_u6_u7_n156 ) );
  NAND2_X1 u1_u6_u7_U55 (.A2( u1_u6_u7_n102 ) , .A1( u1_u6_u7_n103 ) , .ZN( u1_u6_u7_n133 ) );
  NAND2_X1 u1_u6_u7_U56 (.ZN( u1_u6_u7_n112 ) , .A2( u1_u6_u7_n96 ) , .A1( u1_u6_u7_n99 ) );
  NAND2_X1 u1_u6_u7_U57 (.A2( u1_u6_u7_n102 ) , .ZN( u1_u6_u7_n128 ) , .A1( u1_u6_u7_n98 ) );
  NAND2_X1 u1_u6_u7_U58 (.A1( u1_u6_u7_n100 ) , .ZN( u1_u6_u7_n113 ) , .A2( u1_u6_u7_n93 ) );
  NAND2_X1 u1_u6_u7_U59 (.A2( u1_u6_u7_n102 ) , .ZN( u1_u6_u7_n124 ) , .A1( u1_u6_u7_n96 ) );
  INV_X1 u1_u6_u7_U6 (.A( u1_u6_u7_n154 ) , .ZN( u1_u6_u7_n178 ) );
  NAND2_X1 u1_u6_u7_U60 (.ZN( u1_u6_u7_n110 ) , .A1( u1_u6_u7_n95 ) , .A2( u1_u6_u7_n96 ) );
  INV_X1 u1_u6_u7_U61 (.A( u1_u6_u7_n150 ) , .ZN( u1_u6_u7_n164 ) );
  AND2_X1 u1_u6_u7_U62 (.ZN( u1_u6_u7_n134 ) , .A1( u1_u6_u7_n93 ) , .A2( u1_u6_u7_n98 ) );
  NAND2_X1 u1_u6_u7_U63 (.A1( u1_u6_u7_n100 ) , .A2( u1_u6_u7_n102 ) , .ZN( u1_u6_u7_n129 ) );
  NAND2_X1 u1_u6_u7_U64 (.A2( u1_u6_u7_n103 ) , .ZN( u1_u6_u7_n131 ) , .A1( u1_u6_u7_n95 ) );
  NAND2_X1 u1_u6_u7_U65 (.A1( u1_u6_u7_n100 ) , .ZN( u1_u6_u7_n138 ) , .A2( u1_u6_u7_n99 ) );
  NAND2_X1 u1_u6_u7_U66 (.ZN( u1_u6_u7_n132 ) , .A1( u1_u6_u7_n93 ) , .A2( u1_u6_u7_n96 ) );
  NAND2_X1 u1_u6_u7_U67 (.A1( u1_u6_u7_n100 ) , .ZN( u1_u6_u7_n148 ) , .A2( u1_u6_u7_n95 ) );
  NOR2_X1 u1_u6_u7_U68 (.A2( u1_u6_X_47 ) , .ZN( u1_u6_u7_n150 ) , .A1( u1_u6_u7_n163 ) );
  NOR2_X1 u1_u6_u7_U69 (.A2( u1_u6_X_43 ) , .A1( u1_u6_X_44 ) , .ZN( u1_u6_u7_n103 ) );
  AOI211_X1 u1_u6_u7_U7 (.ZN( u1_u6_u7_n116 ) , .A( u1_u6_u7_n155 ) , .C1( u1_u6_u7_n161 ) , .C2( u1_u6_u7_n171 ) , .B( u1_u6_u7_n94 ) );
  NOR2_X1 u1_u6_u7_U70 (.A2( u1_u6_X_48 ) , .A1( u1_u6_u7_n166 ) , .ZN( u1_u6_u7_n95 ) );
  NOR2_X1 u1_u6_u7_U71 (.A2( u1_u6_X_45 ) , .A1( u1_u6_X_48 ) , .ZN( u1_u6_u7_n99 ) );
  NOR2_X1 u1_u6_u7_U72 (.A2( u1_u6_X_44 ) , .A1( u1_u6_u7_n167 ) , .ZN( u1_u6_u7_n98 ) );
  NOR2_X1 u1_u6_u7_U73 (.A2( u1_u6_X_46 ) , .A1( u1_u6_X_47 ) , .ZN( u1_u6_u7_n152 ) );
  AND2_X1 u1_u6_u7_U74 (.A1( u1_u6_X_47 ) , .ZN( u1_u6_u7_n156 ) , .A2( u1_u6_u7_n163 ) );
  NAND2_X1 u1_u6_u7_U75 (.A2( u1_u6_X_46 ) , .A1( u1_u6_X_47 ) , .ZN( u1_u6_u7_n125 ) );
  AND2_X1 u1_u6_u7_U76 (.A2( u1_u6_X_45 ) , .A1( u1_u6_X_48 ) , .ZN( u1_u6_u7_n102 ) );
  AND2_X1 u1_u6_u7_U77 (.A2( u1_u6_X_43 ) , .A1( u1_u6_X_44 ) , .ZN( u1_u6_u7_n96 ) );
  AND2_X1 u1_u6_u7_U78 (.A1( u1_u6_X_44 ) , .ZN( u1_u6_u7_n100 ) , .A2( u1_u6_u7_n167 ) );
  AND2_X1 u1_u6_u7_U79 (.A1( u1_u6_X_48 ) , .A2( u1_u6_u7_n166 ) , .ZN( u1_u6_u7_n93 ) );
  OAI222_X1 u1_u6_u7_U8 (.C2( u1_u6_u7_n101 ) , .B2( u1_u6_u7_n111 ) , .A1( u1_u6_u7_n113 ) , .C1( u1_u6_u7_n146 ) , .A2( u1_u6_u7_n162 ) , .B1( u1_u6_u7_n164 ) , .ZN( u1_u6_u7_n94 ) );
  INV_X1 u1_u6_u7_U80 (.A( u1_u6_X_46 ) , .ZN( u1_u6_u7_n163 ) );
  INV_X1 u1_u6_u7_U81 (.A( u1_u6_X_43 ) , .ZN( u1_u6_u7_n167 ) );
  INV_X1 u1_u6_u7_U82 (.A( u1_u6_X_45 ) , .ZN( u1_u6_u7_n166 ) );
  NAND4_X1 u1_u6_u7_U83 (.ZN( u1_out6_5 ) , .A4( u1_u6_u7_n108 ) , .A3( u1_u6_u7_n109 ) , .A1( u1_u6_u7_n116 ) , .A2( u1_u6_u7_n123 ) );
  AOI22_X1 u1_u6_u7_U84 (.ZN( u1_u6_u7_n109 ) , .A2( u1_u6_u7_n126 ) , .B2( u1_u6_u7_n145 ) , .B1( u1_u6_u7_n156 ) , .A1( u1_u6_u7_n171 ) );
  NOR4_X1 u1_u6_u7_U85 (.A4( u1_u6_u7_n104 ) , .A3( u1_u6_u7_n105 ) , .A2( u1_u6_u7_n106 ) , .A1( u1_u6_u7_n107 ) , .ZN( u1_u6_u7_n108 ) );
  NAND4_X1 u1_u6_u7_U86 (.ZN( u1_out6_21 ) , .A4( u1_u6_u7_n157 ) , .A3( u1_u6_u7_n158 ) , .A2( u1_u6_u7_n159 ) , .A1( u1_u6_u7_n160 ) );
  OAI21_X1 u1_u6_u7_U87 (.B1( u1_u6_u7_n145 ) , .ZN( u1_u6_u7_n160 ) , .A( u1_u6_u7_n161 ) , .B2( u1_u6_u7_n177 ) );
  AOI22_X1 u1_u6_u7_U88 (.B2( u1_u6_u7_n149 ) , .B1( u1_u6_u7_n150 ) , .A2( u1_u6_u7_n151 ) , .A1( u1_u6_u7_n152 ) , .ZN( u1_u6_u7_n158 ) );
  NAND4_X1 u1_u6_u7_U89 (.ZN( u1_out6_15 ) , .A4( u1_u6_u7_n142 ) , .A3( u1_u6_u7_n143 ) , .A2( u1_u6_u7_n144 ) , .A1( u1_u6_u7_n178 ) );
  OAI221_X1 u1_u6_u7_U9 (.C1( u1_u6_u7_n101 ) , .C2( u1_u6_u7_n147 ) , .ZN( u1_u6_u7_n155 ) , .B2( u1_u6_u7_n162 ) , .A( u1_u6_u7_n91 ) , .B1( u1_u6_u7_n92 ) );
  OR2_X1 u1_u6_u7_U90 (.A2( u1_u6_u7_n125 ) , .A1( u1_u6_u7_n129 ) , .ZN( u1_u6_u7_n144 ) );
  AOI22_X1 u1_u6_u7_U91 (.A2( u1_u6_u7_n126 ) , .ZN( u1_u6_u7_n143 ) , .B2( u1_u6_u7_n165 ) , .B1( u1_u6_u7_n173 ) , .A1( u1_u6_u7_n174 ) );
  NAND4_X1 u1_u6_u7_U92 (.ZN( u1_out6_27 ) , .A4( u1_u6_u7_n118 ) , .A3( u1_u6_u7_n119 ) , .A2( u1_u6_u7_n120 ) , .A1( u1_u6_u7_n121 ) );
  OAI21_X1 u1_u6_u7_U93 (.ZN( u1_u6_u7_n121 ) , .B2( u1_u6_u7_n145 ) , .A( u1_u6_u7_n150 ) , .B1( u1_u6_u7_n174 ) );
  OAI21_X1 u1_u6_u7_U94 (.ZN( u1_u6_u7_n120 ) , .A( u1_u6_u7_n161 ) , .B2( u1_u6_u7_n170 ) , .B1( u1_u6_u7_n179 ) );
  NAND3_X1 u1_u6_u7_U95 (.A3( u1_u6_u7_n146 ) , .A2( u1_u6_u7_n147 ) , .A1( u1_u6_u7_n148 ) , .ZN( u1_u6_u7_n151 ) );
  NAND3_X1 u1_u6_u7_U96 (.A3( u1_u6_u7_n131 ) , .A2( u1_u6_u7_n132 ) , .A1( u1_u6_u7_n133 ) , .ZN( u1_u6_u7_n135 ) );
  XOR2_X1 u1_u7_U1 (.B( u1_K8_9 ) , .A( u1_R6_6 ) , .Z( u1_u7_X_9 ) );
  XOR2_X1 u1_u7_U16 (.B( u1_K8_3 ) , .A( u1_R6_2 ) , .Z( u1_u7_X_3 ) );
  XOR2_X1 u1_u7_U2 (.B( u1_K8_8 ) , .A( u1_R6_5 ) , .Z( u1_u7_X_8 ) );
  XOR2_X1 u1_u7_U27 (.B( u1_K8_2 ) , .A( u1_R6_1 ) , .Z( u1_u7_X_2 ) );
  XOR2_X1 u1_u7_U3 (.B( u1_K8_7 ) , .A( u1_R6_4 ) , .Z( u1_u7_X_7 ) );
  XOR2_X1 u1_u7_U38 (.B( u1_K8_1 ) , .A( u1_R6_32 ) , .Z( u1_u7_X_1 ) );
  XOR2_X1 u1_u7_U4 (.B( u1_K8_6 ) , .A( u1_R6_5 ) , .Z( u1_u7_X_6 ) );
  XOR2_X1 u1_u7_U40 (.B( u1_K8_18 ) , .A( u1_R6_13 ) , .Z( u1_u7_X_18 ) );
  XOR2_X1 u1_u7_U41 (.B( u1_K8_17 ) , .A( u1_R6_12 ) , .Z( u1_u7_X_17 ) );
  XOR2_X1 u1_u7_U42 (.B( u1_K8_16 ) , .A( u1_R6_11 ) , .Z( u1_u7_X_16 ) );
  XOR2_X1 u1_u7_U43 (.B( u1_K8_15 ) , .A( u1_R6_10 ) , .Z( u1_u7_X_15 ) );
  XOR2_X1 u1_u7_U44 (.B( u1_K8_14 ) , .A( u1_R6_9 ) , .Z( u1_u7_X_14 ) );
  XOR2_X1 u1_u7_U45 (.B( u1_K8_13 ) , .A( u1_R6_8 ) , .Z( u1_u7_X_13 ) );
  XOR2_X1 u1_u7_U46 (.B( u1_K8_12 ) , .A( u1_R6_9 ) , .Z( u1_u7_X_12 ) );
  XOR2_X1 u1_u7_U47 (.B( u1_K8_11 ) , .A( u1_R6_8 ) , .Z( u1_u7_X_11 ) );
  XOR2_X1 u1_u7_U48 (.B( u1_K8_10 ) , .A( u1_R6_7 ) , .Z( u1_u7_X_10 ) );
  XOR2_X1 u1_u7_U5 (.B( u1_K8_5 ) , .A( u1_R6_4 ) , .Z( u1_u7_X_5 ) );
  XOR2_X1 u1_u7_U6 (.B( u1_K8_4 ) , .A( u1_R6_3 ) , .Z( u1_u7_X_4 ) );
  AND3_X1 u1_u7_u0_U10 (.A2( u1_u7_u0_n112 ) , .ZN( u1_u7_u0_n127 ) , .A3( u1_u7_u0_n130 ) , .A1( u1_u7_u0_n148 ) );
  NAND2_X1 u1_u7_u0_U11 (.ZN( u1_u7_u0_n113 ) , .A1( u1_u7_u0_n139 ) , .A2( u1_u7_u0_n149 ) );
  AND2_X1 u1_u7_u0_U12 (.ZN( u1_u7_u0_n107 ) , .A1( u1_u7_u0_n130 ) , .A2( u1_u7_u0_n140 ) );
  AND2_X1 u1_u7_u0_U13 (.A2( u1_u7_u0_n129 ) , .A1( u1_u7_u0_n130 ) , .ZN( u1_u7_u0_n151 ) );
  AND2_X1 u1_u7_u0_U14 (.A1( u1_u7_u0_n108 ) , .A2( u1_u7_u0_n125 ) , .ZN( u1_u7_u0_n145 ) );
  INV_X1 u1_u7_u0_U15 (.A( u1_u7_u0_n143 ) , .ZN( u1_u7_u0_n173 ) );
  NOR2_X1 u1_u7_u0_U16 (.A2( u1_u7_u0_n136 ) , .ZN( u1_u7_u0_n147 ) , .A1( u1_u7_u0_n160 ) );
  NOR2_X1 u1_u7_u0_U17 (.A1( u1_u7_u0_n163 ) , .A2( u1_u7_u0_n164 ) , .ZN( u1_u7_u0_n95 ) );
  AOI21_X1 u1_u7_u0_U18 (.B1( u1_u7_u0_n103 ) , .ZN( u1_u7_u0_n132 ) , .A( u1_u7_u0_n165 ) , .B2( u1_u7_u0_n93 ) );
  INV_X1 u1_u7_u0_U19 (.A( u1_u7_u0_n142 ) , .ZN( u1_u7_u0_n165 ) );
  OAI22_X1 u1_u7_u0_U20 (.B1( u1_u7_u0_n125 ) , .ZN( u1_u7_u0_n126 ) , .A1( u1_u7_u0_n138 ) , .A2( u1_u7_u0_n146 ) , .B2( u1_u7_u0_n147 ) );
  OAI22_X1 u1_u7_u0_U21 (.B1( u1_u7_u0_n131 ) , .A1( u1_u7_u0_n144 ) , .B2( u1_u7_u0_n147 ) , .A2( u1_u7_u0_n90 ) , .ZN( u1_u7_u0_n91 ) );
  AND3_X1 u1_u7_u0_U22 (.A3( u1_u7_u0_n121 ) , .A2( u1_u7_u0_n125 ) , .A1( u1_u7_u0_n148 ) , .ZN( u1_u7_u0_n90 ) );
  INV_X1 u1_u7_u0_U23 (.A( u1_u7_u0_n136 ) , .ZN( u1_u7_u0_n161 ) );
  AOI22_X1 u1_u7_u0_U24 (.B2( u1_u7_u0_n109 ) , .A2( u1_u7_u0_n110 ) , .ZN( u1_u7_u0_n111 ) , .B1( u1_u7_u0_n118 ) , .A1( u1_u7_u0_n160 ) );
  INV_X1 u1_u7_u0_U25 (.A( u1_u7_u0_n118 ) , .ZN( u1_u7_u0_n158 ) );
  AOI21_X1 u1_u7_u0_U26 (.ZN( u1_u7_u0_n104 ) , .B1( u1_u7_u0_n107 ) , .B2( u1_u7_u0_n141 ) , .A( u1_u7_u0_n144 ) );
  AOI21_X1 u1_u7_u0_U27 (.B1( u1_u7_u0_n127 ) , .B2( u1_u7_u0_n129 ) , .A( u1_u7_u0_n138 ) , .ZN( u1_u7_u0_n96 ) );
  AOI21_X1 u1_u7_u0_U28 (.ZN( u1_u7_u0_n116 ) , .B2( u1_u7_u0_n142 ) , .A( u1_u7_u0_n144 ) , .B1( u1_u7_u0_n166 ) );
  NOR2_X1 u1_u7_u0_U29 (.A1( u1_u7_u0_n120 ) , .ZN( u1_u7_u0_n143 ) , .A2( u1_u7_u0_n167 ) );
  INV_X1 u1_u7_u0_U3 (.A( u1_u7_u0_n113 ) , .ZN( u1_u7_u0_n166 ) );
  OAI221_X1 u1_u7_u0_U30 (.C1( u1_u7_u0_n112 ) , .ZN( u1_u7_u0_n120 ) , .B1( u1_u7_u0_n138 ) , .B2( u1_u7_u0_n141 ) , .C2( u1_u7_u0_n147 ) , .A( u1_u7_u0_n172 ) );
  AOI211_X1 u1_u7_u0_U31 (.B( u1_u7_u0_n115 ) , .A( u1_u7_u0_n116 ) , .C2( u1_u7_u0_n117 ) , .C1( u1_u7_u0_n118 ) , .ZN( u1_u7_u0_n119 ) );
  NAND2_X1 u1_u7_u0_U32 (.A1( u1_u7_u0_n100 ) , .A2( u1_u7_u0_n103 ) , .ZN( u1_u7_u0_n125 ) );
  NAND2_X1 u1_u7_u0_U33 (.A1( u1_u7_u0_n101 ) , .A2( u1_u7_u0_n102 ) , .ZN( u1_u7_u0_n150 ) );
  INV_X1 u1_u7_u0_U34 (.A( u1_u7_u0_n138 ) , .ZN( u1_u7_u0_n160 ) );
  NAND2_X1 u1_u7_u0_U35 (.A1( u1_u7_u0_n102 ) , .ZN( u1_u7_u0_n128 ) , .A2( u1_u7_u0_n95 ) );
  NAND2_X1 u1_u7_u0_U36 (.A1( u1_u7_u0_n100 ) , .ZN( u1_u7_u0_n129 ) , .A2( u1_u7_u0_n95 ) );
  NAND2_X1 u1_u7_u0_U37 (.A2( u1_u7_u0_n100 ) , .ZN( u1_u7_u0_n131 ) , .A1( u1_u7_u0_n92 ) );
  NAND2_X1 u1_u7_u0_U38 (.A2( u1_u7_u0_n100 ) , .A1( u1_u7_u0_n101 ) , .ZN( u1_u7_u0_n139 ) );
  NAND2_X1 u1_u7_u0_U39 (.ZN( u1_u7_u0_n148 ) , .A1( u1_u7_u0_n93 ) , .A2( u1_u7_u0_n95 ) );
  AOI21_X1 u1_u7_u0_U4 (.B1( u1_u7_u0_n114 ) , .ZN( u1_u7_u0_n115 ) , .B2( u1_u7_u0_n129 ) , .A( u1_u7_u0_n161 ) );
  NAND2_X1 u1_u7_u0_U40 (.A2( u1_u7_u0_n102 ) , .A1( u1_u7_u0_n103 ) , .ZN( u1_u7_u0_n149 ) );
  NAND2_X1 u1_u7_u0_U41 (.A2( u1_u7_u0_n102 ) , .ZN( u1_u7_u0_n114 ) , .A1( u1_u7_u0_n92 ) );
  NAND2_X1 u1_u7_u0_U42 (.A2( u1_u7_u0_n101 ) , .ZN( u1_u7_u0_n121 ) , .A1( u1_u7_u0_n93 ) );
  INV_X1 u1_u7_u0_U43 (.ZN( u1_u7_u0_n172 ) , .A( u1_u7_u0_n88 ) );
  OAI222_X1 u1_u7_u0_U44 (.C1( u1_u7_u0_n108 ) , .A1( u1_u7_u0_n125 ) , .B2( u1_u7_u0_n128 ) , .B1( u1_u7_u0_n144 ) , .A2( u1_u7_u0_n158 ) , .C2( u1_u7_u0_n161 ) , .ZN( u1_u7_u0_n88 ) );
  NAND2_X1 u1_u7_u0_U45 (.ZN( u1_u7_u0_n112 ) , .A2( u1_u7_u0_n92 ) , .A1( u1_u7_u0_n93 ) );
  OR3_X1 u1_u7_u0_U46 (.A3( u1_u7_u0_n152 ) , .A2( u1_u7_u0_n153 ) , .A1( u1_u7_u0_n154 ) , .ZN( u1_u7_u0_n155 ) );
  AOI21_X1 u1_u7_u0_U47 (.A( u1_u7_u0_n144 ) , .B2( u1_u7_u0_n145 ) , .B1( u1_u7_u0_n146 ) , .ZN( u1_u7_u0_n154 ) );
  AOI21_X1 u1_u7_u0_U48 (.B2( u1_u7_u0_n150 ) , .B1( u1_u7_u0_n151 ) , .ZN( u1_u7_u0_n152 ) , .A( u1_u7_u0_n158 ) );
  AOI21_X1 u1_u7_u0_U49 (.A( u1_u7_u0_n147 ) , .B2( u1_u7_u0_n148 ) , .B1( u1_u7_u0_n149 ) , .ZN( u1_u7_u0_n153 ) );
  AOI21_X1 u1_u7_u0_U5 (.B2( u1_u7_u0_n131 ) , .ZN( u1_u7_u0_n134 ) , .B1( u1_u7_u0_n151 ) , .A( u1_u7_u0_n158 ) );
  INV_X1 u1_u7_u0_U50 (.ZN( u1_u7_u0_n171 ) , .A( u1_u7_u0_n99 ) );
  OAI211_X1 u1_u7_u0_U51 (.C2( u1_u7_u0_n140 ) , .C1( u1_u7_u0_n161 ) , .A( u1_u7_u0_n169 ) , .B( u1_u7_u0_n98 ) , .ZN( u1_u7_u0_n99 ) );
  INV_X1 u1_u7_u0_U52 (.ZN( u1_u7_u0_n169 ) , .A( u1_u7_u0_n91 ) );
  AOI211_X1 u1_u7_u0_U53 (.C1( u1_u7_u0_n118 ) , .A( u1_u7_u0_n123 ) , .B( u1_u7_u0_n96 ) , .C2( u1_u7_u0_n97 ) , .ZN( u1_u7_u0_n98 ) );
  NOR2_X1 u1_u7_u0_U54 (.A2( u1_u7_X_6 ) , .ZN( u1_u7_u0_n100 ) , .A1( u1_u7_u0_n162 ) );
  NOR2_X1 u1_u7_u0_U55 (.A2( u1_u7_X_4 ) , .A1( u1_u7_X_5 ) , .ZN( u1_u7_u0_n118 ) );
  NOR2_X1 u1_u7_u0_U56 (.A2( u1_u7_X_2 ) , .ZN( u1_u7_u0_n103 ) , .A1( u1_u7_u0_n164 ) );
  NOR2_X1 u1_u7_u0_U57 (.A2( u1_u7_X_1 ) , .A1( u1_u7_X_2 ) , .ZN( u1_u7_u0_n92 ) );
  NOR2_X1 u1_u7_u0_U58 (.A2( u1_u7_X_1 ) , .ZN( u1_u7_u0_n101 ) , .A1( u1_u7_u0_n163 ) );
  NAND2_X1 u1_u7_u0_U59 (.A2( u1_u7_X_4 ) , .A1( u1_u7_X_5 ) , .ZN( u1_u7_u0_n144 ) );
  NOR2_X1 u1_u7_u0_U6 (.A1( u1_u7_u0_n108 ) , .ZN( u1_u7_u0_n123 ) , .A2( u1_u7_u0_n158 ) );
  NOR2_X1 u1_u7_u0_U60 (.A2( u1_u7_X_5 ) , .ZN( u1_u7_u0_n136 ) , .A1( u1_u7_u0_n159 ) );
  NAND2_X1 u1_u7_u0_U61 (.A1( u1_u7_X_5 ) , .ZN( u1_u7_u0_n138 ) , .A2( u1_u7_u0_n159 ) );
  NOR2_X1 u1_u7_u0_U62 (.A2( u1_u7_X_3 ) , .A1( u1_u7_X_6 ) , .ZN( u1_u7_u0_n94 ) );
  AND2_X1 u1_u7_u0_U63 (.A2( u1_u7_X_3 ) , .A1( u1_u7_X_6 ) , .ZN( u1_u7_u0_n102 ) );
  AND2_X1 u1_u7_u0_U64 (.A1( u1_u7_X_6 ) , .A2( u1_u7_u0_n162 ) , .ZN( u1_u7_u0_n93 ) );
  INV_X1 u1_u7_u0_U65 (.A( u1_u7_X_4 ) , .ZN( u1_u7_u0_n159 ) );
  INV_X1 u1_u7_u0_U66 (.A( u1_u7_X_1 ) , .ZN( u1_u7_u0_n164 ) );
  INV_X1 u1_u7_u0_U67 (.A( u1_u7_X_2 ) , .ZN( u1_u7_u0_n163 ) );
  INV_X1 u1_u7_u0_U68 (.A( u1_u7_X_3 ) , .ZN( u1_u7_u0_n162 ) );
  INV_X1 u1_u7_u0_U69 (.A( u1_u7_u0_n126 ) , .ZN( u1_u7_u0_n168 ) );
  OAI21_X1 u1_u7_u0_U7 (.B1( u1_u7_u0_n150 ) , .B2( u1_u7_u0_n158 ) , .A( u1_u7_u0_n172 ) , .ZN( u1_u7_u0_n89 ) );
  AOI211_X1 u1_u7_u0_U70 (.B( u1_u7_u0_n133 ) , .A( u1_u7_u0_n134 ) , .C2( u1_u7_u0_n135 ) , .C1( u1_u7_u0_n136 ) , .ZN( u1_u7_u0_n137 ) );
  OR4_X1 u1_u7_u0_U71 (.ZN( u1_out7_17 ) , .A1( u1_u7_u0_n122 ) , .A2( u1_u7_u0_n123 ) , .A4( u1_u7_u0_n124 ) , .A3( u1_u7_u0_n170 ) );
  AOI21_X1 u1_u7_u0_U72 (.B2( u1_u7_u0_n107 ) , .ZN( u1_u7_u0_n124 ) , .B1( u1_u7_u0_n128 ) , .A( u1_u7_u0_n161 ) );
  INV_X1 u1_u7_u0_U73 (.A( u1_u7_u0_n111 ) , .ZN( u1_u7_u0_n170 ) );
  OR4_X1 u1_u7_u0_U74 (.ZN( u1_out7_31 ) , .A4( u1_u7_u0_n155 ) , .A2( u1_u7_u0_n156 ) , .A1( u1_u7_u0_n157 ) , .A3( u1_u7_u0_n173 ) );
  AOI21_X1 u1_u7_u0_U75 (.A( u1_u7_u0_n138 ) , .B2( u1_u7_u0_n139 ) , .B1( u1_u7_u0_n140 ) , .ZN( u1_u7_u0_n157 ) );
  AOI21_X1 u1_u7_u0_U76 (.B2( u1_u7_u0_n141 ) , .B1( u1_u7_u0_n142 ) , .ZN( u1_u7_u0_n156 ) , .A( u1_u7_u0_n161 ) );
  INV_X1 u1_u7_u0_U77 (.ZN( u1_u7_u0_n174 ) , .A( u1_u7_u0_n89 ) );
  AOI211_X1 u1_u7_u0_U78 (.B( u1_u7_u0_n104 ) , .A( u1_u7_u0_n105 ) , .ZN( u1_u7_u0_n106 ) , .C2( u1_u7_u0_n113 ) , .C1( u1_u7_u0_n160 ) );
  OAI221_X1 u1_u7_u0_U79 (.C1( u1_u7_u0_n121 ) , .ZN( u1_u7_u0_n122 ) , .B2( u1_u7_u0_n127 ) , .A( u1_u7_u0_n143 ) , .B1( u1_u7_u0_n144 ) , .C2( u1_u7_u0_n147 ) );
  AND2_X1 u1_u7_u0_U8 (.A1( u1_u7_u0_n114 ) , .A2( u1_u7_u0_n121 ) , .ZN( u1_u7_u0_n146 ) );
  AOI21_X1 u1_u7_u0_U80 (.B1( u1_u7_u0_n132 ) , .ZN( u1_u7_u0_n133 ) , .A( u1_u7_u0_n144 ) , .B2( u1_u7_u0_n166 ) );
  OAI22_X1 u1_u7_u0_U81 (.ZN( u1_u7_u0_n105 ) , .A2( u1_u7_u0_n132 ) , .B1( u1_u7_u0_n146 ) , .A1( u1_u7_u0_n147 ) , .B2( u1_u7_u0_n161 ) );
  NAND2_X1 u1_u7_u0_U82 (.ZN( u1_u7_u0_n110 ) , .A2( u1_u7_u0_n132 ) , .A1( u1_u7_u0_n145 ) );
  INV_X1 u1_u7_u0_U83 (.A( u1_u7_u0_n119 ) , .ZN( u1_u7_u0_n167 ) );
  NAND2_X1 u1_u7_u0_U84 (.A2( u1_u7_u0_n103 ) , .ZN( u1_u7_u0_n140 ) , .A1( u1_u7_u0_n94 ) );
  NAND2_X1 u1_u7_u0_U85 (.A1( u1_u7_u0_n101 ) , .ZN( u1_u7_u0_n130 ) , .A2( u1_u7_u0_n94 ) );
  NAND2_X1 u1_u7_u0_U86 (.ZN( u1_u7_u0_n108 ) , .A1( u1_u7_u0_n92 ) , .A2( u1_u7_u0_n94 ) );
  NAND2_X1 u1_u7_u0_U87 (.ZN( u1_u7_u0_n142 ) , .A1( u1_u7_u0_n94 ) , .A2( u1_u7_u0_n95 ) );
  NAND3_X1 u1_u7_u0_U88 (.ZN( u1_out7_23 ) , .A3( u1_u7_u0_n137 ) , .A1( u1_u7_u0_n168 ) , .A2( u1_u7_u0_n171 ) );
  NAND3_X1 u1_u7_u0_U89 (.A3( u1_u7_u0_n127 ) , .A2( u1_u7_u0_n128 ) , .ZN( u1_u7_u0_n135 ) , .A1( u1_u7_u0_n150 ) );
  AND2_X1 u1_u7_u0_U9 (.A1( u1_u7_u0_n131 ) , .ZN( u1_u7_u0_n141 ) , .A2( u1_u7_u0_n150 ) );
  NAND3_X1 u1_u7_u0_U90 (.ZN( u1_u7_u0_n117 ) , .A3( u1_u7_u0_n132 ) , .A2( u1_u7_u0_n139 ) , .A1( u1_u7_u0_n148 ) );
  NAND3_X1 u1_u7_u0_U91 (.ZN( u1_u7_u0_n109 ) , .A2( u1_u7_u0_n114 ) , .A3( u1_u7_u0_n140 ) , .A1( u1_u7_u0_n149 ) );
  NAND3_X1 u1_u7_u0_U92 (.ZN( u1_out7_9 ) , .A3( u1_u7_u0_n106 ) , .A2( u1_u7_u0_n171 ) , .A1( u1_u7_u0_n174 ) );
  NAND3_X1 u1_u7_u0_U93 (.A2( u1_u7_u0_n128 ) , .A1( u1_u7_u0_n132 ) , .A3( u1_u7_u0_n146 ) , .ZN( u1_u7_u0_n97 ) );
  AOI21_X1 u1_u7_u1_U10 (.B2( u1_u7_u1_n155 ) , .B1( u1_u7_u1_n156 ) , .ZN( u1_u7_u1_n157 ) , .A( u1_u7_u1_n174 ) );
  NAND3_X1 u1_u7_u1_U100 (.ZN( u1_u7_u1_n113 ) , .A1( u1_u7_u1_n120 ) , .A3( u1_u7_u1_n133 ) , .A2( u1_u7_u1_n155 ) );
  NAND2_X1 u1_u7_u1_U11 (.ZN( u1_u7_u1_n140 ) , .A2( u1_u7_u1_n150 ) , .A1( u1_u7_u1_n155 ) );
  NAND2_X1 u1_u7_u1_U12 (.A1( u1_u7_u1_n131 ) , .ZN( u1_u7_u1_n147 ) , .A2( u1_u7_u1_n153 ) );
  AOI22_X1 u1_u7_u1_U13 (.B2( u1_u7_u1_n136 ) , .A2( u1_u7_u1_n137 ) , .ZN( u1_u7_u1_n143 ) , .A1( u1_u7_u1_n171 ) , .B1( u1_u7_u1_n173 ) );
  INV_X1 u1_u7_u1_U14 (.A( u1_u7_u1_n147 ) , .ZN( u1_u7_u1_n181 ) );
  INV_X1 u1_u7_u1_U15 (.A( u1_u7_u1_n139 ) , .ZN( u1_u7_u1_n174 ) );
  OR4_X1 u1_u7_u1_U16 (.A4( u1_u7_u1_n106 ) , .A3( u1_u7_u1_n107 ) , .ZN( u1_u7_u1_n108 ) , .A1( u1_u7_u1_n117 ) , .A2( u1_u7_u1_n184 ) );
  AOI21_X1 u1_u7_u1_U17 (.ZN( u1_u7_u1_n106 ) , .A( u1_u7_u1_n112 ) , .B1( u1_u7_u1_n154 ) , .B2( u1_u7_u1_n156 ) );
  AOI21_X1 u1_u7_u1_U18 (.ZN( u1_u7_u1_n107 ) , .B1( u1_u7_u1_n134 ) , .B2( u1_u7_u1_n149 ) , .A( u1_u7_u1_n174 ) );
  INV_X1 u1_u7_u1_U19 (.A( u1_u7_u1_n101 ) , .ZN( u1_u7_u1_n184 ) );
  INV_X1 u1_u7_u1_U20 (.A( u1_u7_u1_n112 ) , .ZN( u1_u7_u1_n171 ) );
  NAND2_X1 u1_u7_u1_U21 (.ZN( u1_u7_u1_n141 ) , .A1( u1_u7_u1_n153 ) , .A2( u1_u7_u1_n156 ) );
  AND2_X1 u1_u7_u1_U22 (.A1( u1_u7_u1_n123 ) , .ZN( u1_u7_u1_n134 ) , .A2( u1_u7_u1_n161 ) );
  NAND2_X1 u1_u7_u1_U23 (.A2( u1_u7_u1_n115 ) , .A1( u1_u7_u1_n116 ) , .ZN( u1_u7_u1_n148 ) );
  NAND2_X1 u1_u7_u1_U24 (.A2( u1_u7_u1_n133 ) , .A1( u1_u7_u1_n135 ) , .ZN( u1_u7_u1_n159 ) );
  NAND2_X1 u1_u7_u1_U25 (.A2( u1_u7_u1_n115 ) , .A1( u1_u7_u1_n120 ) , .ZN( u1_u7_u1_n132 ) );
  INV_X1 u1_u7_u1_U26 (.A( u1_u7_u1_n154 ) , .ZN( u1_u7_u1_n178 ) );
  INV_X1 u1_u7_u1_U27 (.A( u1_u7_u1_n151 ) , .ZN( u1_u7_u1_n183 ) );
  AND2_X1 u1_u7_u1_U28 (.A1( u1_u7_u1_n129 ) , .A2( u1_u7_u1_n133 ) , .ZN( u1_u7_u1_n149 ) );
  INV_X1 u1_u7_u1_U29 (.A( u1_u7_u1_n131 ) , .ZN( u1_u7_u1_n180 ) );
  INV_X1 u1_u7_u1_U3 (.A( u1_u7_u1_n159 ) , .ZN( u1_u7_u1_n182 ) );
  OAI221_X1 u1_u7_u1_U30 (.A( u1_u7_u1_n119 ) , .C2( u1_u7_u1_n129 ) , .ZN( u1_u7_u1_n138 ) , .B2( u1_u7_u1_n152 ) , .C1( u1_u7_u1_n174 ) , .B1( u1_u7_u1_n187 ) );
  INV_X1 u1_u7_u1_U31 (.A( u1_u7_u1_n148 ) , .ZN( u1_u7_u1_n187 ) );
  AOI211_X1 u1_u7_u1_U32 (.B( u1_u7_u1_n117 ) , .A( u1_u7_u1_n118 ) , .ZN( u1_u7_u1_n119 ) , .C2( u1_u7_u1_n146 ) , .C1( u1_u7_u1_n159 ) );
  NOR2_X1 u1_u7_u1_U33 (.A1( u1_u7_u1_n168 ) , .A2( u1_u7_u1_n176 ) , .ZN( u1_u7_u1_n98 ) );
  AOI211_X1 u1_u7_u1_U34 (.B( u1_u7_u1_n162 ) , .A( u1_u7_u1_n163 ) , .C2( u1_u7_u1_n164 ) , .ZN( u1_u7_u1_n165 ) , .C1( u1_u7_u1_n171 ) );
  AOI21_X1 u1_u7_u1_U35 (.A( u1_u7_u1_n160 ) , .B2( u1_u7_u1_n161 ) , .ZN( u1_u7_u1_n162 ) , .B1( u1_u7_u1_n182 ) );
  OR2_X1 u1_u7_u1_U36 (.A2( u1_u7_u1_n157 ) , .A1( u1_u7_u1_n158 ) , .ZN( u1_u7_u1_n163 ) );
  NAND2_X1 u1_u7_u1_U37 (.A1( u1_u7_u1_n128 ) , .ZN( u1_u7_u1_n146 ) , .A2( u1_u7_u1_n160 ) );
  NAND2_X1 u1_u7_u1_U38 (.A2( u1_u7_u1_n112 ) , .ZN( u1_u7_u1_n139 ) , .A1( u1_u7_u1_n152 ) );
  NAND2_X1 u1_u7_u1_U39 (.A1( u1_u7_u1_n105 ) , .ZN( u1_u7_u1_n156 ) , .A2( u1_u7_u1_n99 ) );
  AOI221_X1 u1_u7_u1_U4 (.A( u1_u7_u1_n138 ) , .C2( u1_u7_u1_n139 ) , .C1( u1_u7_u1_n140 ) , .B2( u1_u7_u1_n141 ) , .ZN( u1_u7_u1_n142 ) , .B1( u1_u7_u1_n175 ) );
  AOI221_X1 u1_u7_u1_U40 (.B1( u1_u7_u1_n140 ) , .ZN( u1_u7_u1_n167 ) , .B2( u1_u7_u1_n172 ) , .C2( u1_u7_u1_n175 ) , .C1( u1_u7_u1_n178 ) , .A( u1_u7_u1_n188 ) );
  INV_X1 u1_u7_u1_U41 (.ZN( u1_u7_u1_n188 ) , .A( u1_u7_u1_n97 ) );
  AOI211_X1 u1_u7_u1_U42 (.A( u1_u7_u1_n118 ) , .C1( u1_u7_u1_n132 ) , .C2( u1_u7_u1_n139 ) , .B( u1_u7_u1_n96 ) , .ZN( u1_u7_u1_n97 ) );
  AOI21_X1 u1_u7_u1_U43 (.B2( u1_u7_u1_n121 ) , .B1( u1_u7_u1_n135 ) , .A( u1_u7_u1_n152 ) , .ZN( u1_u7_u1_n96 ) );
  NOR2_X1 u1_u7_u1_U44 (.ZN( u1_u7_u1_n117 ) , .A1( u1_u7_u1_n121 ) , .A2( u1_u7_u1_n160 ) );
  OAI21_X1 u1_u7_u1_U45 (.B2( u1_u7_u1_n123 ) , .ZN( u1_u7_u1_n145 ) , .B1( u1_u7_u1_n160 ) , .A( u1_u7_u1_n185 ) );
  INV_X1 u1_u7_u1_U46 (.A( u1_u7_u1_n122 ) , .ZN( u1_u7_u1_n185 ) );
  AOI21_X1 u1_u7_u1_U47 (.B2( u1_u7_u1_n120 ) , .B1( u1_u7_u1_n121 ) , .ZN( u1_u7_u1_n122 ) , .A( u1_u7_u1_n128 ) );
  AOI21_X1 u1_u7_u1_U48 (.A( u1_u7_u1_n128 ) , .B2( u1_u7_u1_n129 ) , .ZN( u1_u7_u1_n130 ) , .B1( u1_u7_u1_n150 ) );
  NAND2_X1 u1_u7_u1_U49 (.ZN( u1_u7_u1_n112 ) , .A1( u1_u7_u1_n169 ) , .A2( u1_u7_u1_n170 ) );
  AOI211_X1 u1_u7_u1_U5 (.ZN( u1_u7_u1_n124 ) , .A( u1_u7_u1_n138 ) , .C2( u1_u7_u1_n139 ) , .B( u1_u7_u1_n145 ) , .C1( u1_u7_u1_n147 ) );
  NAND2_X1 u1_u7_u1_U50 (.ZN( u1_u7_u1_n129 ) , .A2( u1_u7_u1_n95 ) , .A1( u1_u7_u1_n98 ) );
  NAND2_X1 u1_u7_u1_U51 (.A1( u1_u7_u1_n102 ) , .ZN( u1_u7_u1_n154 ) , .A2( u1_u7_u1_n99 ) );
  NAND2_X1 u1_u7_u1_U52 (.A2( u1_u7_u1_n100 ) , .ZN( u1_u7_u1_n135 ) , .A1( u1_u7_u1_n99 ) );
  AOI21_X1 u1_u7_u1_U53 (.A( u1_u7_u1_n152 ) , .B2( u1_u7_u1_n153 ) , .B1( u1_u7_u1_n154 ) , .ZN( u1_u7_u1_n158 ) );
  INV_X1 u1_u7_u1_U54 (.A( u1_u7_u1_n160 ) , .ZN( u1_u7_u1_n175 ) );
  NAND2_X1 u1_u7_u1_U55 (.A1( u1_u7_u1_n100 ) , .ZN( u1_u7_u1_n116 ) , .A2( u1_u7_u1_n95 ) );
  NAND2_X1 u1_u7_u1_U56 (.A1( u1_u7_u1_n102 ) , .ZN( u1_u7_u1_n131 ) , .A2( u1_u7_u1_n95 ) );
  NAND2_X1 u1_u7_u1_U57 (.A2( u1_u7_u1_n104 ) , .ZN( u1_u7_u1_n121 ) , .A1( u1_u7_u1_n98 ) );
  NAND2_X1 u1_u7_u1_U58 (.A1( u1_u7_u1_n103 ) , .ZN( u1_u7_u1_n153 ) , .A2( u1_u7_u1_n98 ) );
  NAND2_X1 u1_u7_u1_U59 (.A2( u1_u7_u1_n104 ) , .A1( u1_u7_u1_n105 ) , .ZN( u1_u7_u1_n133 ) );
  AOI22_X1 u1_u7_u1_U6 (.B2( u1_u7_u1_n113 ) , .A2( u1_u7_u1_n114 ) , .ZN( u1_u7_u1_n125 ) , .A1( u1_u7_u1_n171 ) , .B1( u1_u7_u1_n173 ) );
  NAND2_X1 u1_u7_u1_U60 (.ZN( u1_u7_u1_n150 ) , .A2( u1_u7_u1_n98 ) , .A1( u1_u7_u1_n99 ) );
  NAND2_X1 u1_u7_u1_U61 (.A1( u1_u7_u1_n105 ) , .ZN( u1_u7_u1_n155 ) , .A2( u1_u7_u1_n95 ) );
  OAI21_X1 u1_u7_u1_U62 (.ZN( u1_u7_u1_n109 ) , .B1( u1_u7_u1_n129 ) , .B2( u1_u7_u1_n160 ) , .A( u1_u7_u1_n167 ) );
  NAND2_X1 u1_u7_u1_U63 (.A2( u1_u7_u1_n100 ) , .A1( u1_u7_u1_n103 ) , .ZN( u1_u7_u1_n120 ) );
  NAND2_X1 u1_u7_u1_U64 (.A1( u1_u7_u1_n102 ) , .A2( u1_u7_u1_n104 ) , .ZN( u1_u7_u1_n115 ) );
  NAND2_X1 u1_u7_u1_U65 (.A2( u1_u7_u1_n100 ) , .A1( u1_u7_u1_n104 ) , .ZN( u1_u7_u1_n151 ) );
  NAND2_X1 u1_u7_u1_U66 (.A2( u1_u7_u1_n103 ) , .A1( u1_u7_u1_n105 ) , .ZN( u1_u7_u1_n161 ) );
  INV_X1 u1_u7_u1_U67 (.A( u1_u7_u1_n152 ) , .ZN( u1_u7_u1_n173 ) );
  INV_X1 u1_u7_u1_U68 (.A( u1_u7_u1_n128 ) , .ZN( u1_u7_u1_n172 ) );
  NAND2_X1 u1_u7_u1_U69 (.A2( u1_u7_u1_n102 ) , .A1( u1_u7_u1_n103 ) , .ZN( u1_u7_u1_n123 ) );
  NAND2_X1 u1_u7_u1_U7 (.ZN( u1_u7_u1_n114 ) , .A1( u1_u7_u1_n134 ) , .A2( u1_u7_u1_n156 ) );
  NOR2_X1 u1_u7_u1_U70 (.A2( u1_u7_X_7 ) , .A1( u1_u7_X_8 ) , .ZN( u1_u7_u1_n95 ) );
  NOR2_X1 u1_u7_u1_U71 (.A1( u1_u7_X_12 ) , .A2( u1_u7_X_9 ) , .ZN( u1_u7_u1_n100 ) );
  NOR2_X1 u1_u7_u1_U72 (.A2( u1_u7_X_8 ) , .A1( u1_u7_u1_n177 ) , .ZN( u1_u7_u1_n99 ) );
  NOR2_X1 u1_u7_u1_U73 (.A2( u1_u7_X_12 ) , .ZN( u1_u7_u1_n102 ) , .A1( u1_u7_u1_n176 ) );
  NOR2_X1 u1_u7_u1_U74 (.A2( u1_u7_X_9 ) , .ZN( u1_u7_u1_n105 ) , .A1( u1_u7_u1_n168 ) );
  NAND2_X1 u1_u7_u1_U75 (.A1( u1_u7_X_10 ) , .ZN( u1_u7_u1_n160 ) , .A2( u1_u7_u1_n169 ) );
  NAND2_X1 u1_u7_u1_U76 (.A2( u1_u7_X_10 ) , .A1( u1_u7_X_11 ) , .ZN( u1_u7_u1_n152 ) );
  NAND2_X1 u1_u7_u1_U77 (.A1( u1_u7_X_11 ) , .ZN( u1_u7_u1_n128 ) , .A2( u1_u7_u1_n170 ) );
  AND2_X1 u1_u7_u1_U78 (.A2( u1_u7_X_7 ) , .A1( u1_u7_X_8 ) , .ZN( u1_u7_u1_n104 ) );
  AND2_X1 u1_u7_u1_U79 (.A1( u1_u7_X_8 ) , .ZN( u1_u7_u1_n103 ) , .A2( u1_u7_u1_n177 ) );
  NOR2_X1 u1_u7_u1_U8 (.A1( u1_u7_u1_n112 ) , .A2( u1_u7_u1_n116 ) , .ZN( u1_u7_u1_n118 ) );
  INV_X1 u1_u7_u1_U80 (.A( u1_u7_X_10 ) , .ZN( u1_u7_u1_n170 ) );
  INV_X1 u1_u7_u1_U81 (.A( u1_u7_X_9 ) , .ZN( u1_u7_u1_n176 ) );
  INV_X1 u1_u7_u1_U82 (.A( u1_u7_X_11 ) , .ZN( u1_u7_u1_n169 ) );
  INV_X1 u1_u7_u1_U83 (.A( u1_u7_X_12 ) , .ZN( u1_u7_u1_n168 ) );
  INV_X1 u1_u7_u1_U84 (.A( u1_u7_X_7 ) , .ZN( u1_u7_u1_n177 ) );
  NAND4_X1 u1_u7_u1_U85 (.ZN( u1_out7_18 ) , .A4( u1_u7_u1_n165 ) , .A3( u1_u7_u1_n166 ) , .A1( u1_u7_u1_n167 ) , .A2( u1_u7_u1_n186 ) );
  AOI22_X1 u1_u7_u1_U86 (.B2( u1_u7_u1_n146 ) , .B1( u1_u7_u1_n147 ) , .A2( u1_u7_u1_n148 ) , .ZN( u1_u7_u1_n166 ) , .A1( u1_u7_u1_n172 ) );
  INV_X1 u1_u7_u1_U87 (.A( u1_u7_u1_n145 ) , .ZN( u1_u7_u1_n186 ) );
  NAND4_X1 u1_u7_u1_U88 (.ZN( u1_out7_2 ) , .A4( u1_u7_u1_n142 ) , .A3( u1_u7_u1_n143 ) , .A2( u1_u7_u1_n144 ) , .A1( u1_u7_u1_n179 ) );
  OAI21_X1 u1_u7_u1_U89 (.B2( u1_u7_u1_n132 ) , .ZN( u1_u7_u1_n144 ) , .A( u1_u7_u1_n146 ) , .B1( u1_u7_u1_n180 ) );
  OAI21_X1 u1_u7_u1_U9 (.ZN( u1_u7_u1_n101 ) , .B1( u1_u7_u1_n141 ) , .A( u1_u7_u1_n146 ) , .B2( u1_u7_u1_n183 ) );
  INV_X1 u1_u7_u1_U90 (.A( u1_u7_u1_n130 ) , .ZN( u1_u7_u1_n179 ) );
  NAND4_X1 u1_u7_u1_U91 (.ZN( u1_out7_28 ) , .A4( u1_u7_u1_n124 ) , .A3( u1_u7_u1_n125 ) , .A2( u1_u7_u1_n126 ) , .A1( u1_u7_u1_n127 ) );
  OAI21_X1 u1_u7_u1_U92 (.ZN( u1_u7_u1_n127 ) , .B2( u1_u7_u1_n139 ) , .B1( u1_u7_u1_n175 ) , .A( u1_u7_u1_n183 ) );
  OAI21_X1 u1_u7_u1_U93 (.ZN( u1_u7_u1_n126 ) , .B2( u1_u7_u1_n140 ) , .A( u1_u7_u1_n146 ) , .B1( u1_u7_u1_n178 ) );
  OR4_X1 u1_u7_u1_U94 (.ZN( u1_out7_13 ) , .A4( u1_u7_u1_n108 ) , .A3( u1_u7_u1_n109 ) , .A2( u1_u7_u1_n110 ) , .A1( u1_u7_u1_n111 ) );
  AOI21_X1 u1_u7_u1_U95 (.ZN( u1_u7_u1_n111 ) , .A( u1_u7_u1_n128 ) , .B2( u1_u7_u1_n131 ) , .B1( u1_u7_u1_n135 ) );
  AOI21_X1 u1_u7_u1_U96 (.ZN( u1_u7_u1_n110 ) , .A( u1_u7_u1_n116 ) , .B1( u1_u7_u1_n152 ) , .B2( u1_u7_u1_n160 ) );
  NAND3_X1 u1_u7_u1_U97 (.A3( u1_u7_u1_n149 ) , .A2( u1_u7_u1_n150 ) , .A1( u1_u7_u1_n151 ) , .ZN( u1_u7_u1_n164 ) );
  NAND3_X1 u1_u7_u1_U98 (.A3( u1_u7_u1_n134 ) , .A2( u1_u7_u1_n135 ) , .ZN( u1_u7_u1_n136 ) , .A1( u1_u7_u1_n151 ) );
  NAND3_X1 u1_u7_u1_U99 (.A1( u1_u7_u1_n133 ) , .ZN( u1_u7_u1_n137 ) , .A2( u1_u7_u1_n154 ) , .A3( u1_u7_u1_n181 ) );
  OAI22_X1 u1_u7_u2_U10 (.ZN( u1_u7_u2_n109 ) , .A2( u1_u7_u2_n113 ) , .B2( u1_u7_u2_n133 ) , .B1( u1_u7_u2_n167 ) , .A1( u1_u7_u2_n168 ) );
  NAND3_X1 u1_u7_u2_U100 (.A2( u1_u7_u2_n100 ) , .A1( u1_u7_u2_n104 ) , .A3( u1_u7_u2_n138 ) , .ZN( u1_u7_u2_n98 ) );
  OAI22_X1 u1_u7_u2_U11 (.B1( u1_u7_u2_n151 ) , .A2( u1_u7_u2_n152 ) , .A1( u1_u7_u2_n153 ) , .ZN( u1_u7_u2_n160 ) , .B2( u1_u7_u2_n168 ) );
  NOR3_X1 u1_u7_u2_U12 (.A1( u1_u7_u2_n150 ) , .ZN( u1_u7_u2_n151 ) , .A3( u1_u7_u2_n175 ) , .A2( u1_u7_u2_n188 ) );
  AOI21_X1 u1_u7_u2_U13 (.ZN( u1_u7_u2_n144 ) , .B2( u1_u7_u2_n155 ) , .A( u1_u7_u2_n172 ) , .B1( u1_u7_u2_n185 ) );
  AOI21_X1 u1_u7_u2_U14 (.B2( u1_u7_u2_n143 ) , .ZN( u1_u7_u2_n145 ) , .B1( u1_u7_u2_n152 ) , .A( u1_u7_u2_n171 ) );
  AOI21_X1 u1_u7_u2_U15 (.B2( u1_u7_u2_n120 ) , .B1( u1_u7_u2_n121 ) , .ZN( u1_u7_u2_n126 ) , .A( u1_u7_u2_n167 ) );
  INV_X1 u1_u7_u2_U16 (.A( u1_u7_u2_n156 ) , .ZN( u1_u7_u2_n171 ) );
  INV_X1 u1_u7_u2_U17 (.A( u1_u7_u2_n120 ) , .ZN( u1_u7_u2_n188 ) );
  NAND2_X1 u1_u7_u2_U18 (.A2( u1_u7_u2_n122 ) , .ZN( u1_u7_u2_n150 ) , .A1( u1_u7_u2_n152 ) );
  INV_X1 u1_u7_u2_U19 (.A( u1_u7_u2_n153 ) , .ZN( u1_u7_u2_n170 ) );
  INV_X1 u1_u7_u2_U20 (.A( u1_u7_u2_n137 ) , .ZN( u1_u7_u2_n173 ) );
  NAND2_X1 u1_u7_u2_U21 (.A1( u1_u7_u2_n132 ) , .A2( u1_u7_u2_n139 ) , .ZN( u1_u7_u2_n157 ) );
  INV_X1 u1_u7_u2_U22 (.A( u1_u7_u2_n113 ) , .ZN( u1_u7_u2_n178 ) );
  INV_X1 u1_u7_u2_U23 (.A( u1_u7_u2_n139 ) , .ZN( u1_u7_u2_n175 ) );
  INV_X1 u1_u7_u2_U24 (.A( u1_u7_u2_n155 ) , .ZN( u1_u7_u2_n181 ) );
  INV_X1 u1_u7_u2_U25 (.A( u1_u7_u2_n119 ) , .ZN( u1_u7_u2_n177 ) );
  INV_X1 u1_u7_u2_U26 (.A( u1_u7_u2_n116 ) , .ZN( u1_u7_u2_n180 ) );
  INV_X1 u1_u7_u2_U27 (.A( u1_u7_u2_n131 ) , .ZN( u1_u7_u2_n179 ) );
  INV_X1 u1_u7_u2_U28 (.A( u1_u7_u2_n154 ) , .ZN( u1_u7_u2_n176 ) );
  NAND2_X1 u1_u7_u2_U29 (.A2( u1_u7_u2_n116 ) , .A1( u1_u7_u2_n117 ) , .ZN( u1_u7_u2_n118 ) );
  NOR2_X1 u1_u7_u2_U3 (.ZN( u1_u7_u2_n121 ) , .A2( u1_u7_u2_n177 ) , .A1( u1_u7_u2_n180 ) );
  INV_X1 u1_u7_u2_U30 (.A( u1_u7_u2_n132 ) , .ZN( u1_u7_u2_n182 ) );
  INV_X1 u1_u7_u2_U31 (.A( u1_u7_u2_n158 ) , .ZN( u1_u7_u2_n183 ) );
  OAI21_X1 u1_u7_u2_U32 (.A( u1_u7_u2_n156 ) , .B1( u1_u7_u2_n157 ) , .ZN( u1_u7_u2_n158 ) , .B2( u1_u7_u2_n179 ) );
  NOR2_X1 u1_u7_u2_U33 (.ZN( u1_u7_u2_n156 ) , .A1( u1_u7_u2_n166 ) , .A2( u1_u7_u2_n169 ) );
  NOR2_X1 u1_u7_u2_U34 (.A2( u1_u7_u2_n114 ) , .ZN( u1_u7_u2_n137 ) , .A1( u1_u7_u2_n140 ) );
  NOR2_X1 u1_u7_u2_U35 (.A2( u1_u7_u2_n138 ) , .ZN( u1_u7_u2_n153 ) , .A1( u1_u7_u2_n156 ) );
  AOI211_X1 u1_u7_u2_U36 (.ZN( u1_u7_u2_n130 ) , .C1( u1_u7_u2_n138 ) , .C2( u1_u7_u2_n179 ) , .B( u1_u7_u2_n96 ) , .A( u1_u7_u2_n97 ) );
  OAI22_X1 u1_u7_u2_U37 (.B1( u1_u7_u2_n133 ) , .A2( u1_u7_u2_n137 ) , .A1( u1_u7_u2_n152 ) , .B2( u1_u7_u2_n168 ) , .ZN( u1_u7_u2_n97 ) );
  OAI221_X1 u1_u7_u2_U38 (.B1( u1_u7_u2_n113 ) , .C1( u1_u7_u2_n132 ) , .A( u1_u7_u2_n149 ) , .B2( u1_u7_u2_n171 ) , .C2( u1_u7_u2_n172 ) , .ZN( u1_u7_u2_n96 ) );
  OAI221_X1 u1_u7_u2_U39 (.A( u1_u7_u2_n115 ) , .C2( u1_u7_u2_n123 ) , .B2( u1_u7_u2_n143 ) , .B1( u1_u7_u2_n153 ) , .ZN( u1_u7_u2_n163 ) , .C1( u1_u7_u2_n168 ) );
  INV_X1 u1_u7_u2_U4 (.A( u1_u7_u2_n134 ) , .ZN( u1_u7_u2_n185 ) );
  OAI21_X1 u1_u7_u2_U40 (.A( u1_u7_u2_n114 ) , .ZN( u1_u7_u2_n115 ) , .B1( u1_u7_u2_n176 ) , .B2( u1_u7_u2_n178 ) );
  OAI221_X1 u1_u7_u2_U41 (.A( u1_u7_u2_n135 ) , .B2( u1_u7_u2_n136 ) , .B1( u1_u7_u2_n137 ) , .ZN( u1_u7_u2_n162 ) , .C2( u1_u7_u2_n167 ) , .C1( u1_u7_u2_n185 ) );
  AND3_X1 u1_u7_u2_U42 (.A3( u1_u7_u2_n131 ) , .A2( u1_u7_u2_n132 ) , .A1( u1_u7_u2_n133 ) , .ZN( u1_u7_u2_n136 ) );
  AOI22_X1 u1_u7_u2_U43 (.ZN( u1_u7_u2_n135 ) , .B1( u1_u7_u2_n140 ) , .A1( u1_u7_u2_n156 ) , .B2( u1_u7_u2_n180 ) , .A2( u1_u7_u2_n188 ) );
  AOI21_X1 u1_u7_u2_U44 (.ZN( u1_u7_u2_n149 ) , .B1( u1_u7_u2_n173 ) , .B2( u1_u7_u2_n188 ) , .A( u1_u7_u2_n95 ) );
  AND3_X1 u1_u7_u2_U45 (.A2( u1_u7_u2_n100 ) , .A1( u1_u7_u2_n104 ) , .A3( u1_u7_u2_n156 ) , .ZN( u1_u7_u2_n95 ) );
  OAI21_X1 u1_u7_u2_U46 (.A( u1_u7_u2_n101 ) , .B2( u1_u7_u2_n121 ) , .B1( u1_u7_u2_n153 ) , .ZN( u1_u7_u2_n164 ) );
  NAND2_X1 u1_u7_u2_U47 (.A2( u1_u7_u2_n100 ) , .A1( u1_u7_u2_n107 ) , .ZN( u1_u7_u2_n155 ) );
  NAND2_X1 u1_u7_u2_U48 (.A2( u1_u7_u2_n105 ) , .A1( u1_u7_u2_n108 ) , .ZN( u1_u7_u2_n143 ) );
  NAND2_X1 u1_u7_u2_U49 (.A1( u1_u7_u2_n104 ) , .A2( u1_u7_u2_n106 ) , .ZN( u1_u7_u2_n152 ) );
  INV_X1 u1_u7_u2_U5 (.A( u1_u7_u2_n150 ) , .ZN( u1_u7_u2_n184 ) );
  NAND2_X1 u1_u7_u2_U50 (.A1( u1_u7_u2_n100 ) , .A2( u1_u7_u2_n105 ) , .ZN( u1_u7_u2_n132 ) );
  INV_X1 u1_u7_u2_U51 (.A( u1_u7_u2_n140 ) , .ZN( u1_u7_u2_n168 ) );
  INV_X1 u1_u7_u2_U52 (.A( u1_u7_u2_n138 ) , .ZN( u1_u7_u2_n167 ) );
  OAI21_X1 u1_u7_u2_U53 (.A( u1_u7_u2_n141 ) , .B2( u1_u7_u2_n142 ) , .ZN( u1_u7_u2_n146 ) , .B1( u1_u7_u2_n153 ) );
  OAI21_X1 u1_u7_u2_U54 (.A( u1_u7_u2_n140 ) , .ZN( u1_u7_u2_n141 ) , .B1( u1_u7_u2_n176 ) , .B2( u1_u7_u2_n177 ) );
  NOR3_X1 u1_u7_u2_U55 (.ZN( u1_u7_u2_n142 ) , .A3( u1_u7_u2_n175 ) , .A2( u1_u7_u2_n178 ) , .A1( u1_u7_u2_n181 ) );
  INV_X1 u1_u7_u2_U56 (.ZN( u1_u7_u2_n187 ) , .A( u1_u7_u2_n99 ) );
  OAI21_X1 u1_u7_u2_U57 (.B1( u1_u7_u2_n137 ) , .B2( u1_u7_u2_n143 ) , .A( u1_u7_u2_n98 ) , .ZN( u1_u7_u2_n99 ) );
  NAND2_X1 u1_u7_u2_U58 (.A1( u1_u7_u2_n102 ) , .A2( u1_u7_u2_n106 ) , .ZN( u1_u7_u2_n113 ) );
  NAND2_X1 u1_u7_u2_U59 (.A1( u1_u7_u2_n106 ) , .A2( u1_u7_u2_n107 ) , .ZN( u1_u7_u2_n131 ) );
  NOR4_X1 u1_u7_u2_U6 (.A4( u1_u7_u2_n124 ) , .A3( u1_u7_u2_n125 ) , .A2( u1_u7_u2_n126 ) , .A1( u1_u7_u2_n127 ) , .ZN( u1_u7_u2_n128 ) );
  NAND2_X1 u1_u7_u2_U60 (.A1( u1_u7_u2_n103 ) , .A2( u1_u7_u2_n107 ) , .ZN( u1_u7_u2_n139 ) );
  NAND2_X1 u1_u7_u2_U61 (.A1( u1_u7_u2_n103 ) , .A2( u1_u7_u2_n105 ) , .ZN( u1_u7_u2_n133 ) );
  NAND2_X1 u1_u7_u2_U62 (.A1( u1_u7_u2_n102 ) , .A2( u1_u7_u2_n103 ) , .ZN( u1_u7_u2_n154 ) );
  NAND2_X1 u1_u7_u2_U63 (.A2( u1_u7_u2_n103 ) , .A1( u1_u7_u2_n104 ) , .ZN( u1_u7_u2_n119 ) );
  NAND2_X1 u1_u7_u2_U64 (.A2( u1_u7_u2_n107 ) , .A1( u1_u7_u2_n108 ) , .ZN( u1_u7_u2_n123 ) );
  NAND2_X1 u1_u7_u2_U65 (.A1( u1_u7_u2_n104 ) , .A2( u1_u7_u2_n108 ) , .ZN( u1_u7_u2_n122 ) );
  INV_X1 u1_u7_u2_U66 (.A( u1_u7_u2_n114 ) , .ZN( u1_u7_u2_n172 ) );
  NAND2_X1 u1_u7_u2_U67 (.A2( u1_u7_u2_n100 ) , .A1( u1_u7_u2_n102 ) , .ZN( u1_u7_u2_n116 ) );
  NAND2_X1 u1_u7_u2_U68 (.A1( u1_u7_u2_n102 ) , .A2( u1_u7_u2_n108 ) , .ZN( u1_u7_u2_n120 ) );
  NAND2_X1 u1_u7_u2_U69 (.A2( u1_u7_u2_n105 ) , .A1( u1_u7_u2_n106 ) , .ZN( u1_u7_u2_n117 ) );
  AOI21_X1 u1_u7_u2_U7 (.B2( u1_u7_u2_n119 ) , .ZN( u1_u7_u2_n127 ) , .A( u1_u7_u2_n137 ) , .B1( u1_u7_u2_n155 ) );
  NOR2_X1 u1_u7_u2_U70 (.A2( u1_u7_X_16 ) , .ZN( u1_u7_u2_n140 ) , .A1( u1_u7_u2_n166 ) );
  NOR2_X1 u1_u7_u2_U71 (.A2( u1_u7_X_13 ) , .A1( u1_u7_X_14 ) , .ZN( u1_u7_u2_n100 ) );
  NOR2_X1 u1_u7_u2_U72 (.A2( u1_u7_X_16 ) , .A1( u1_u7_X_17 ) , .ZN( u1_u7_u2_n138 ) );
  NOR2_X1 u1_u7_u2_U73 (.A2( u1_u7_X_15 ) , .A1( u1_u7_X_18 ) , .ZN( u1_u7_u2_n104 ) );
  NOR2_X1 u1_u7_u2_U74 (.A2( u1_u7_X_14 ) , .ZN( u1_u7_u2_n103 ) , .A1( u1_u7_u2_n174 ) );
  NOR2_X1 u1_u7_u2_U75 (.A2( u1_u7_X_15 ) , .ZN( u1_u7_u2_n102 ) , .A1( u1_u7_u2_n165 ) );
  NOR2_X1 u1_u7_u2_U76 (.A2( u1_u7_X_17 ) , .ZN( u1_u7_u2_n114 ) , .A1( u1_u7_u2_n169 ) );
  AND2_X1 u1_u7_u2_U77 (.A1( u1_u7_X_15 ) , .ZN( u1_u7_u2_n105 ) , .A2( u1_u7_u2_n165 ) );
  AND2_X1 u1_u7_u2_U78 (.A2( u1_u7_X_15 ) , .A1( u1_u7_X_18 ) , .ZN( u1_u7_u2_n107 ) );
  AND2_X1 u1_u7_u2_U79 (.A1( u1_u7_X_14 ) , .ZN( u1_u7_u2_n106 ) , .A2( u1_u7_u2_n174 ) );
  AOI21_X1 u1_u7_u2_U8 (.ZN( u1_u7_u2_n124 ) , .B1( u1_u7_u2_n131 ) , .B2( u1_u7_u2_n143 ) , .A( u1_u7_u2_n172 ) );
  AND2_X1 u1_u7_u2_U80 (.A1( u1_u7_X_13 ) , .A2( u1_u7_X_14 ) , .ZN( u1_u7_u2_n108 ) );
  INV_X1 u1_u7_u2_U81 (.A( u1_u7_X_16 ) , .ZN( u1_u7_u2_n169 ) );
  INV_X1 u1_u7_u2_U82 (.A( u1_u7_X_17 ) , .ZN( u1_u7_u2_n166 ) );
  INV_X1 u1_u7_u2_U83 (.A( u1_u7_X_13 ) , .ZN( u1_u7_u2_n174 ) );
  INV_X1 u1_u7_u2_U84 (.A( u1_u7_X_18 ) , .ZN( u1_u7_u2_n165 ) );
  NAND4_X1 u1_u7_u2_U85 (.ZN( u1_out7_24 ) , .A4( u1_u7_u2_n111 ) , .A3( u1_u7_u2_n112 ) , .A1( u1_u7_u2_n130 ) , .A2( u1_u7_u2_n187 ) );
  AOI221_X1 u1_u7_u2_U86 (.A( u1_u7_u2_n109 ) , .B1( u1_u7_u2_n110 ) , .ZN( u1_u7_u2_n111 ) , .C1( u1_u7_u2_n134 ) , .C2( u1_u7_u2_n170 ) , .B2( u1_u7_u2_n173 ) );
  AOI21_X1 u1_u7_u2_U87 (.ZN( u1_u7_u2_n112 ) , .B2( u1_u7_u2_n156 ) , .A( u1_u7_u2_n164 ) , .B1( u1_u7_u2_n181 ) );
  NAND4_X1 u1_u7_u2_U88 (.ZN( u1_out7_30 ) , .A4( u1_u7_u2_n147 ) , .A3( u1_u7_u2_n148 ) , .A2( u1_u7_u2_n149 ) , .A1( u1_u7_u2_n187 ) );
  NOR3_X1 u1_u7_u2_U89 (.A3( u1_u7_u2_n144 ) , .A2( u1_u7_u2_n145 ) , .A1( u1_u7_u2_n146 ) , .ZN( u1_u7_u2_n147 ) );
  AOI21_X1 u1_u7_u2_U9 (.B2( u1_u7_u2_n123 ) , .ZN( u1_u7_u2_n125 ) , .A( u1_u7_u2_n171 ) , .B1( u1_u7_u2_n184 ) );
  AOI21_X1 u1_u7_u2_U90 (.B2( u1_u7_u2_n138 ) , .ZN( u1_u7_u2_n148 ) , .A( u1_u7_u2_n162 ) , .B1( u1_u7_u2_n182 ) );
  NAND4_X1 u1_u7_u2_U91 (.ZN( u1_out7_16 ) , .A4( u1_u7_u2_n128 ) , .A3( u1_u7_u2_n129 ) , .A1( u1_u7_u2_n130 ) , .A2( u1_u7_u2_n186 ) );
  AOI22_X1 u1_u7_u2_U92 (.A2( u1_u7_u2_n118 ) , .ZN( u1_u7_u2_n129 ) , .A1( u1_u7_u2_n140 ) , .B1( u1_u7_u2_n157 ) , .B2( u1_u7_u2_n170 ) );
  INV_X1 u1_u7_u2_U93 (.A( u1_u7_u2_n163 ) , .ZN( u1_u7_u2_n186 ) );
  OR4_X1 u1_u7_u2_U94 (.ZN( u1_out7_6 ) , .A4( u1_u7_u2_n161 ) , .A3( u1_u7_u2_n162 ) , .A2( u1_u7_u2_n163 ) , .A1( u1_u7_u2_n164 ) );
  OR3_X1 u1_u7_u2_U95 (.A2( u1_u7_u2_n159 ) , .A1( u1_u7_u2_n160 ) , .ZN( u1_u7_u2_n161 ) , .A3( u1_u7_u2_n183 ) );
  AOI21_X1 u1_u7_u2_U96 (.B2( u1_u7_u2_n154 ) , .B1( u1_u7_u2_n155 ) , .ZN( u1_u7_u2_n159 ) , .A( u1_u7_u2_n167 ) );
  NAND3_X1 u1_u7_u2_U97 (.A2( u1_u7_u2_n117 ) , .A1( u1_u7_u2_n122 ) , .A3( u1_u7_u2_n123 ) , .ZN( u1_u7_u2_n134 ) );
  NAND3_X1 u1_u7_u2_U98 (.ZN( u1_u7_u2_n110 ) , .A2( u1_u7_u2_n131 ) , .A3( u1_u7_u2_n139 ) , .A1( u1_u7_u2_n154 ) );
  NAND3_X1 u1_u7_u2_U99 (.A2( u1_u7_u2_n100 ) , .ZN( u1_u7_u2_n101 ) , .A1( u1_u7_u2_n104 ) , .A3( u1_u7_u2_n114 ) );
  XOR2_X1 u1_u8_U10 (.B( u1_K9_45 ) , .A( u1_R7_30 ) , .Z( u1_u8_X_45 ) );
  XOR2_X1 u1_u8_U11 (.B( u1_K9_44 ) , .A( u1_R7_29 ) , .Z( u1_u8_X_44 ) );
  XOR2_X1 u1_u8_U12 (.B( u1_K9_43 ) , .A( u1_R7_28 ) , .Z( u1_u8_X_43 ) );
  XOR2_X1 u1_u8_U7 (.B( u1_K9_48 ) , .A( u1_R7_1 ) , .Z( u1_u8_X_48 ) );
  XOR2_X1 u1_u8_U8 (.B( u1_K9_47 ) , .A( u1_R7_32 ) , .Z( u1_u8_X_47 ) );
  XOR2_X1 u1_u8_U9 (.B( u1_K9_46 ) , .A( u1_R7_31 ) , .Z( u1_u8_X_46 ) );
  AND3_X1 u1_u8_u7_U10 (.A3( u1_u8_u7_n110 ) , .A2( u1_u8_u7_n127 ) , .A1( u1_u8_u7_n132 ) , .ZN( u1_u8_u7_n92 ) );
  OAI21_X1 u1_u8_u7_U11 (.A( u1_u8_u7_n161 ) , .B1( u1_u8_u7_n168 ) , .B2( u1_u8_u7_n173 ) , .ZN( u1_u8_u7_n91 ) );
  AOI211_X1 u1_u8_u7_U12 (.A( u1_u8_u7_n117 ) , .ZN( u1_u8_u7_n118 ) , .C2( u1_u8_u7_n126 ) , .C1( u1_u8_u7_n177 ) , .B( u1_u8_u7_n180 ) );
  OAI22_X1 u1_u8_u7_U13 (.B1( u1_u8_u7_n115 ) , .ZN( u1_u8_u7_n117 ) , .A2( u1_u8_u7_n133 ) , .A1( u1_u8_u7_n137 ) , .B2( u1_u8_u7_n162 ) );
  INV_X1 u1_u8_u7_U14 (.A( u1_u8_u7_n116 ) , .ZN( u1_u8_u7_n180 ) );
  NOR3_X1 u1_u8_u7_U15 (.ZN( u1_u8_u7_n115 ) , .A3( u1_u8_u7_n145 ) , .A2( u1_u8_u7_n168 ) , .A1( u1_u8_u7_n169 ) );
  OAI211_X1 u1_u8_u7_U16 (.B( u1_u8_u7_n122 ) , .A( u1_u8_u7_n123 ) , .C2( u1_u8_u7_n124 ) , .ZN( u1_u8_u7_n154 ) , .C1( u1_u8_u7_n162 ) );
  AOI222_X1 u1_u8_u7_U17 (.ZN( u1_u8_u7_n122 ) , .C2( u1_u8_u7_n126 ) , .C1( u1_u8_u7_n145 ) , .B1( u1_u8_u7_n161 ) , .A2( u1_u8_u7_n165 ) , .B2( u1_u8_u7_n170 ) , .A1( u1_u8_u7_n176 ) );
  INV_X1 u1_u8_u7_U18 (.A( u1_u8_u7_n133 ) , .ZN( u1_u8_u7_n176 ) );
  NOR3_X1 u1_u8_u7_U19 (.A2( u1_u8_u7_n134 ) , .A1( u1_u8_u7_n135 ) , .ZN( u1_u8_u7_n136 ) , .A3( u1_u8_u7_n171 ) );
  NOR2_X1 u1_u8_u7_U20 (.A1( u1_u8_u7_n130 ) , .A2( u1_u8_u7_n134 ) , .ZN( u1_u8_u7_n153 ) );
  INV_X1 u1_u8_u7_U21 (.A( u1_u8_u7_n101 ) , .ZN( u1_u8_u7_n165 ) );
  NOR2_X1 u1_u8_u7_U22 (.ZN( u1_u8_u7_n111 ) , .A2( u1_u8_u7_n134 ) , .A1( u1_u8_u7_n169 ) );
  AOI21_X1 u1_u8_u7_U23 (.ZN( u1_u8_u7_n104 ) , .B2( u1_u8_u7_n112 ) , .B1( u1_u8_u7_n127 ) , .A( u1_u8_u7_n164 ) );
  AOI21_X1 u1_u8_u7_U24 (.ZN( u1_u8_u7_n106 ) , .B1( u1_u8_u7_n133 ) , .B2( u1_u8_u7_n146 ) , .A( u1_u8_u7_n162 ) );
  AOI21_X1 u1_u8_u7_U25 (.A( u1_u8_u7_n101 ) , .ZN( u1_u8_u7_n107 ) , .B2( u1_u8_u7_n128 ) , .B1( u1_u8_u7_n175 ) );
  INV_X1 u1_u8_u7_U26 (.A( u1_u8_u7_n138 ) , .ZN( u1_u8_u7_n171 ) );
  INV_X1 u1_u8_u7_U27 (.A( u1_u8_u7_n131 ) , .ZN( u1_u8_u7_n177 ) );
  INV_X1 u1_u8_u7_U28 (.A( u1_u8_u7_n110 ) , .ZN( u1_u8_u7_n174 ) );
  NAND2_X1 u1_u8_u7_U29 (.A1( u1_u8_u7_n129 ) , .A2( u1_u8_u7_n132 ) , .ZN( u1_u8_u7_n149 ) );
  OAI21_X1 u1_u8_u7_U3 (.ZN( u1_u8_u7_n159 ) , .A( u1_u8_u7_n165 ) , .B2( u1_u8_u7_n171 ) , .B1( u1_u8_u7_n174 ) );
  NAND2_X1 u1_u8_u7_U30 (.A1( u1_u8_u7_n113 ) , .A2( u1_u8_u7_n124 ) , .ZN( u1_u8_u7_n130 ) );
  INV_X1 u1_u8_u7_U31 (.A( u1_u8_u7_n112 ) , .ZN( u1_u8_u7_n173 ) );
  INV_X1 u1_u8_u7_U32 (.A( u1_u8_u7_n128 ) , .ZN( u1_u8_u7_n168 ) );
  INV_X1 u1_u8_u7_U33 (.A( u1_u8_u7_n148 ) , .ZN( u1_u8_u7_n169 ) );
  INV_X1 u1_u8_u7_U34 (.A( u1_u8_u7_n127 ) , .ZN( u1_u8_u7_n179 ) );
  NOR2_X1 u1_u8_u7_U35 (.ZN( u1_u8_u7_n101 ) , .A2( u1_u8_u7_n150 ) , .A1( u1_u8_u7_n156 ) );
  AOI211_X1 u1_u8_u7_U36 (.B( u1_u8_u7_n154 ) , .A( u1_u8_u7_n155 ) , .C1( u1_u8_u7_n156 ) , .ZN( u1_u8_u7_n157 ) , .C2( u1_u8_u7_n172 ) );
  INV_X1 u1_u8_u7_U37 (.A( u1_u8_u7_n153 ) , .ZN( u1_u8_u7_n172 ) );
  AOI211_X1 u1_u8_u7_U38 (.B( u1_u8_u7_n139 ) , .A( u1_u8_u7_n140 ) , .C2( u1_u8_u7_n141 ) , .ZN( u1_u8_u7_n142 ) , .C1( u1_u8_u7_n156 ) );
  NAND4_X1 u1_u8_u7_U39 (.A3( u1_u8_u7_n127 ) , .A2( u1_u8_u7_n128 ) , .A1( u1_u8_u7_n129 ) , .ZN( u1_u8_u7_n141 ) , .A4( u1_u8_u7_n147 ) );
  INV_X1 u1_u8_u7_U4 (.A( u1_u8_u7_n111 ) , .ZN( u1_u8_u7_n170 ) );
  AOI21_X1 u1_u8_u7_U40 (.A( u1_u8_u7_n137 ) , .B1( u1_u8_u7_n138 ) , .ZN( u1_u8_u7_n139 ) , .B2( u1_u8_u7_n146 ) );
  OAI22_X1 u1_u8_u7_U41 (.B1( u1_u8_u7_n136 ) , .ZN( u1_u8_u7_n140 ) , .A1( u1_u8_u7_n153 ) , .B2( u1_u8_u7_n162 ) , .A2( u1_u8_u7_n164 ) );
  AOI21_X1 u1_u8_u7_U42 (.ZN( u1_u8_u7_n123 ) , .B1( u1_u8_u7_n165 ) , .B2( u1_u8_u7_n177 ) , .A( u1_u8_u7_n97 ) );
  AOI21_X1 u1_u8_u7_U43 (.B2( u1_u8_u7_n113 ) , .B1( u1_u8_u7_n124 ) , .A( u1_u8_u7_n125 ) , .ZN( u1_u8_u7_n97 ) );
  INV_X1 u1_u8_u7_U44 (.A( u1_u8_u7_n125 ) , .ZN( u1_u8_u7_n161 ) );
  INV_X1 u1_u8_u7_U45 (.A( u1_u8_u7_n152 ) , .ZN( u1_u8_u7_n162 ) );
  AOI22_X1 u1_u8_u7_U46 (.A2( u1_u8_u7_n114 ) , .ZN( u1_u8_u7_n119 ) , .B1( u1_u8_u7_n130 ) , .A1( u1_u8_u7_n156 ) , .B2( u1_u8_u7_n165 ) );
  NAND2_X1 u1_u8_u7_U47 (.A2( u1_u8_u7_n112 ) , .ZN( u1_u8_u7_n114 ) , .A1( u1_u8_u7_n175 ) );
  AND2_X1 u1_u8_u7_U48 (.ZN( u1_u8_u7_n145 ) , .A2( u1_u8_u7_n98 ) , .A1( u1_u8_u7_n99 ) );
  NOR2_X1 u1_u8_u7_U49 (.ZN( u1_u8_u7_n137 ) , .A1( u1_u8_u7_n150 ) , .A2( u1_u8_u7_n161 ) );
  INV_X1 u1_u8_u7_U5 (.A( u1_u8_u7_n149 ) , .ZN( u1_u8_u7_n175 ) );
  AOI21_X1 u1_u8_u7_U50 (.ZN( u1_u8_u7_n105 ) , .B2( u1_u8_u7_n110 ) , .A( u1_u8_u7_n125 ) , .B1( u1_u8_u7_n147 ) );
  NAND2_X1 u1_u8_u7_U51 (.ZN( u1_u8_u7_n146 ) , .A1( u1_u8_u7_n95 ) , .A2( u1_u8_u7_n98 ) );
  NAND2_X1 u1_u8_u7_U52 (.A2( u1_u8_u7_n103 ) , .ZN( u1_u8_u7_n147 ) , .A1( u1_u8_u7_n93 ) );
  NAND2_X1 u1_u8_u7_U53 (.A1( u1_u8_u7_n103 ) , .ZN( u1_u8_u7_n127 ) , .A2( u1_u8_u7_n99 ) );
  OR2_X1 u1_u8_u7_U54 (.ZN( u1_u8_u7_n126 ) , .A2( u1_u8_u7_n152 ) , .A1( u1_u8_u7_n156 ) );
  NAND2_X1 u1_u8_u7_U55 (.A2( u1_u8_u7_n102 ) , .A1( u1_u8_u7_n103 ) , .ZN( u1_u8_u7_n133 ) );
  NAND2_X1 u1_u8_u7_U56 (.ZN( u1_u8_u7_n112 ) , .A2( u1_u8_u7_n96 ) , .A1( u1_u8_u7_n99 ) );
  NAND2_X1 u1_u8_u7_U57 (.A2( u1_u8_u7_n102 ) , .ZN( u1_u8_u7_n128 ) , .A1( u1_u8_u7_n98 ) );
  NAND2_X1 u1_u8_u7_U58 (.A1( u1_u8_u7_n100 ) , .ZN( u1_u8_u7_n113 ) , .A2( u1_u8_u7_n93 ) );
  NAND2_X1 u1_u8_u7_U59 (.A2( u1_u8_u7_n102 ) , .ZN( u1_u8_u7_n124 ) , .A1( u1_u8_u7_n96 ) );
  INV_X1 u1_u8_u7_U6 (.A( u1_u8_u7_n154 ) , .ZN( u1_u8_u7_n178 ) );
  NAND2_X1 u1_u8_u7_U60 (.ZN( u1_u8_u7_n110 ) , .A1( u1_u8_u7_n95 ) , .A2( u1_u8_u7_n96 ) );
  INV_X1 u1_u8_u7_U61 (.A( u1_u8_u7_n150 ) , .ZN( u1_u8_u7_n164 ) );
  AND2_X1 u1_u8_u7_U62 (.ZN( u1_u8_u7_n134 ) , .A1( u1_u8_u7_n93 ) , .A2( u1_u8_u7_n98 ) );
  NAND2_X1 u1_u8_u7_U63 (.A1( u1_u8_u7_n100 ) , .A2( u1_u8_u7_n102 ) , .ZN( u1_u8_u7_n129 ) );
  NAND2_X1 u1_u8_u7_U64 (.A2( u1_u8_u7_n103 ) , .ZN( u1_u8_u7_n131 ) , .A1( u1_u8_u7_n95 ) );
  NAND2_X1 u1_u8_u7_U65 (.A1( u1_u8_u7_n100 ) , .ZN( u1_u8_u7_n138 ) , .A2( u1_u8_u7_n99 ) );
  NAND2_X1 u1_u8_u7_U66 (.ZN( u1_u8_u7_n132 ) , .A1( u1_u8_u7_n93 ) , .A2( u1_u8_u7_n96 ) );
  NAND2_X1 u1_u8_u7_U67 (.A1( u1_u8_u7_n100 ) , .ZN( u1_u8_u7_n148 ) , .A2( u1_u8_u7_n95 ) );
  NOR2_X1 u1_u8_u7_U68 (.A2( u1_u8_X_47 ) , .ZN( u1_u8_u7_n150 ) , .A1( u1_u8_u7_n163 ) );
  NOR2_X1 u1_u8_u7_U69 (.A2( u1_u8_X_43 ) , .A1( u1_u8_X_44 ) , .ZN( u1_u8_u7_n103 ) );
  AOI211_X1 u1_u8_u7_U7 (.ZN( u1_u8_u7_n116 ) , .A( u1_u8_u7_n155 ) , .C1( u1_u8_u7_n161 ) , .C2( u1_u8_u7_n171 ) , .B( u1_u8_u7_n94 ) );
  NOR2_X1 u1_u8_u7_U70 (.A2( u1_u8_X_48 ) , .A1( u1_u8_u7_n166 ) , .ZN( u1_u8_u7_n95 ) );
  NOR2_X1 u1_u8_u7_U71 (.A2( u1_u8_X_45 ) , .A1( u1_u8_X_48 ) , .ZN( u1_u8_u7_n99 ) );
  NOR2_X1 u1_u8_u7_U72 (.A2( u1_u8_X_44 ) , .A1( u1_u8_u7_n167 ) , .ZN( u1_u8_u7_n98 ) );
  NOR2_X1 u1_u8_u7_U73 (.A2( u1_u8_X_46 ) , .A1( u1_u8_X_47 ) , .ZN( u1_u8_u7_n152 ) );
  AND2_X1 u1_u8_u7_U74 (.A1( u1_u8_X_47 ) , .ZN( u1_u8_u7_n156 ) , .A2( u1_u8_u7_n163 ) );
  NAND2_X1 u1_u8_u7_U75 (.A2( u1_u8_X_46 ) , .A1( u1_u8_X_47 ) , .ZN( u1_u8_u7_n125 ) );
  AND2_X1 u1_u8_u7_U76 (.A2( u1_u8_X_45 ) , .A1( u1_u8_X_48 ) , .ZN( u1_u8_u7_n102 ) );
  AND2_X1 u1_u8_u7_U77 (.A2( u1_u8_X_43 ) , .A1( u1_u8_X_44 ) , .ZN( u1_u8_u7_n96 ) );
  AND2_X1 u1_u8_u7_U78 (.A1( u1_u8_X_44 ) , .ZN( u1_u8_u7_n100 ) , .A2( u1_u8_u7_n167 ) );
  AND2_X1 u1_u8_u7_U79 (.A1( u1_u8_X_48 ) , .A2( u1_u8_u7_n166 ) , .ZN( u1_u8_u7_n93 ) );
  OAI222_X1 u1_u8_u7_U8 (.C2( u1_u8_u7_n101 ) , .B2( u1_u8_u7_n111 ) , .A1( u1_u8_u7_n113 ) , .C1( u1_u8_u7_n146 ) , .A2( u1_u8_u7_n162 ) , .B1( u1_u8_u7_n164 ) , .ZN( u1_u8_u7_n94 ) );
  INV_X1 u1_u8_u7_U80 (.A( u1_u8_X_46 ) , .ZN( u1_u8_u7_n163 ) );
  INV_X1 u1_u8_u7_U81 (.A( u1_u8_X_43 ) , .ZN( u1_u8_u7_n167 ) );
  INV_X1 u1_u8_u7_U82 (.A( u1_u8_X_45 ) , .ZN( u1_u8_u7_n166 ) );
  NAND4_X1 u1_u8_u7_U83 (.ZN( u1_out8_5 ) , .A4( u1_u8_u7_n108 ) , .A3( u1_u8_u7_n109 ) , .A1( u1_u8_u7_n116 ) , .A2( u1_u8_u7_n123 ) );
  AOI22_X1 u1_u8_u7_U84 (.ZN( u1_u8_u7_n109 ) , .A2( u1_u8_u7_n126 ) , .B2( u1_u8_u7_n145 ) , .B1( u1_u8_u7_n156 ) , .A1( u1_u8_u7_n171 ) );
  NOR4_X1 u1_u8_u7_U85 (.A4( u1_u8_u7_n104 ) , .A3( u1_u8_u7_n105 ) , .A2( u1_u8_u7_n106 ) , .A1( u1_u8_u7_n107 ) , .ZN( u1_u8_u7_n108 ) );
  NAND4_X1 u1_u8_u7_U86 (.ZN( u1_out8_27 ) , .A4( u1_u8_u7_n118 ) , .A3( u1_u8_u7_n119 ) , .A2( u1_u8_u7_n120 ) , .A1( u1_u8_u7_n121 ) );
  OAI21_X1 u1_u8_u7_U87 (.ZN( u1_u8_u7_n121 ) , .B2( u1_u8_u7_n145 ) , .A( u1_u8_u7_n150 ) , .B1( u1_u8_u7_n174 ) );
  OAI21_X1 u1_u8_u7_U88 (.ZN( u1_u8_u7_n120 ) , .A( u1_u8_u7_n161 ) , .B2( u1_u8_u7_n170 ) , .B1( u1_u8_u7_n179 ) );
  NAND4_X1 u1_u8_u7_U89 (.ZN( u1_out8_21 ) , .A4( u1_u8_u7_n157 ) , .A3( u1_u8_u7_n158 ) , .A2( u1_u8_u7_n159 ) , .A1( u1_u8_u7_n160 ) );
  OAI221_X1 u1_u8_u7_U9 (.C1( u1_u8_u7_n101 ) , .C2( u1_u8_u7_n147 ) , .ZN( u1_u8_u7_n155 ) , .B2( u1_u8_u7_n162 ) , .A( u1_u8_u7_n91 ) , .B1( u1_u8_u7_n92 ) );
  OAI21_X1 u1_u8_u7_U90 (.B1( u1_u8_u7_n145 ) , .ZN( u1_u8_u7_n160 ) , .A( u1_u8_u7_n161 ) , .B2( u1_u8_u7_n177 ) );
  AOI22_X1 u1_u8_u7_U91 (.B2( u1_u8_u7_n149 ) , .B1( u1_u8_u7_n150 ) , .A2( u1_u8_u7_n151 ) , .A1( u1_u8_u7_n152 ) , .ZN( u1_u8_u7_n158 ) );
  NAND4_X1 u1_u8_u7_U92 (.ZN( u1_out8_15 ) , .A4( u1_u8_u7_n142 ) , .A3( u1_u8_u7_n143 ) , .A2( u1_u8_u7_n144 ) , .A1( u1_u8_u7_n178 ) );
  OR2_X1 u1_u8_u7_U93 (.A2( u1_u8_u7_n125 ) , .A1( u1_u8_u7_n129 ) , .ZN( u1_u8_u7_n144 ) );
  AOI22_X1 u1_u8_u7_U94 (.A2( u1_u8_u7_n126 ) , .ZN( u1_u8_u7_n143 ) , .B2( u1_u8_u7_n165 ) , .B1( u1_u8_u7_n173 ) , .A1( u1_u8_u7_n174 ) );
  NAND3_X1 u1_u8_u7_U95 (.A3( u1_u8_u7_n146 ) , .A2( u1_u8_u7_n147 ) , .A1( u1_u8_u7_n148 ) , .ZN( u1_u8_u7_n151 ) );
  NAND3_X1 u1_u8_u7_U96 (.A3( u1_u8_u7_n131 ) , .A2( u1_u8_u7_n132 ) , .A1( u1_u8_u7_n133 ) , .ZN( u1_u8_u7_n135 ) );
  OAI21_X1 u1_uk_U1008 (.ZN( u1_K8_4 ) , .A( u1_uk_n1146 ) , .B2( u1_uk_n1537 ) , .B1( u1_uk_n17 ) );
  NAND2_X1 u1_uk_U1009 (.A1( u1_uk_K_r6_19 ) , .ZN( u1_uk_n1146 ) , .A2( u1_uk_n27 ) );
  OAI21_X1 u1_uk_U1016 (.ZN( u1_K5_45 ) , .A( u1_uk_n1084 ) , .B2( u1_uk_n1400 ) , .B1( u1_uk_n99 ) );
  NAND2_X1 u1_uk_U1017 (.A1( u1_uk_K_r3_43 ) , .ZN( u1_uk_n1084 ) , .A2( u1_uk_n11 ) );
  OAI22_X1 u1_uk_U103 (.ZN( u1_K7_41 ) , .A2( u1_uk_n1486 ) , .B2( u1_uk_n1516 ) , .A1( u1_uk_n187 ) , .B1( u1_uk_n292 ) );
  OAI21_X1 u1_uk_U1032 (.ZN( u1_K9_44 ) , .A( u1_uk_n1168 ) , .B2( u1_uk_n1615 ) , .B1( u1_uk_n223 ) );
  NAND2_X1 u1_uk_U1033 (.A1( u1_uk_K_r7_0 ) , .ZN( u1_uk_n1168 ) , .A2( u1_uk_n207 ) );
  OAI21_X1 u1_uk_U1034 (.ZN( u1_K12_6 ) , .B2( u1_uk_n1732 ) , .B1( u1_uk_n230 ) , .A( u1_uk_n662 ) );
  NAND2_X1 u1_uk_U1035 (.A1( u1_uk_K_r10_10 ) , .A2( u1_uk_n251 ) , .ZN( u1_uk_n662 ) );
  OAI22_X1 u1_uk_U104 (.ZN( u1_K4_41 ) , .B2( u1_uk_n1349 ) , .A2( u1_uk_n1366 ) , .A1( u1_uk_n141 ) , .B1( u1_uk_n298 ) );
  OAI21_X1 u1_uk_U1042 (.ZN( u1_K16_41 ) , .B2( u1_uk_n1245 ) , .B1( u1_uk_n155 ) , .A( u1_uk_n991 ) );
  NAND2_X1 u1_uk_U1043 (.A1( u1_uk_K_r14_42 ) , .A2( u1_uk_n141 ) , .ZN( u1_uk_n991 ) );
  OAI21_X1 u1_uk_U1048 (.ZN( u1_K16_28 ) , .B2( u1_uk_n1219 ) , .A( u1_uk_n984 ) , .B1( u1_uk_n99 ) );
  NAND2_X1 u1_uk_U1049 (.A1( u1_uk_K_r14_8 ) , .A2( u1_uk_n11 ) , .ZN( u1_uk_n984 ) );
  OAI21_X1 u1_uk_U1062 (.ZN( u1_K15_14 ) , .B1( u1_uk_n102 ) , .B2( u1_uk_n1851 ) , .A( u1_uk_n966 ) );
  NAND2_X1 u1_uk_U1063 (.A1( u1_uk_K_r13_32 ) , .A2( u1_uk_n27 ) , .ZN( u1_uk_n966 ) );
  OAI21_X1 u1_uk_U1068 (.ZN( u1_K16_42 ) , .B2( u1_uk_n1241 ) , .B1( u1_uk_n155 ) , .A( u1_uk_n992 ) );
  NAND2_X1 u1_uk_U1069 (.A1( u1_uk_K_r14_38 ) , .A2( u1_uk_n31 ) , .ZN( u1_uk_n992 ) );
  OAI21_X1 u1_uk_U1072 (.ZN( u1_K7_38 ) , .A( u1_uk_n1122 ) , .B1( u1_uk_n148 ) , .B2( u1_uk_n1499 ) );
  NAND2_X1 u1_uk_U1073 (.A1( u1_uk_K_r5_8 ) , .ZN( u1_uk_n1122 ) , .A2( u1_uk_n17 ) );
  OAI21_X1 u1_uk_U1076 (.ZN( u1_K4_38 ) , .A( u1_uk_n1064 ) , .B2( u1_uk_n1383 ) , .B1( u1_uk_n92 ) );
  NAND2_X1 u1_uk_U1077 (.A1( u1_uk_K_r2_50 ) , .ZN( u1_uk_n1064 ) , .A2( u1_uk_n155 ) );
  OAI22_X1 u1_uk_U109 (.ZN( u1_K15_5 ) , .A1( u1_uk_n147 ) , .B2( u1_uk_n1859 ) , .A2( u1_uk_n1862 ) , .B1( u1_uk_n217 ) );
  INV_X1 u1_uk_U11 (.A( u1_uk_n298 ) , .ZN( u1_uk_n92 ) );
  OAI21_X1 u1_uk_U1105 (.ZN( u1_K8_14 ) , .A( u1_uk_n1129 ) , .B2( u1_uk_n1559 ) , .B1( u1_uk_n203 ) );
  NAND2_X1 u1_uk_U1106 (.A1( u1_uk_K_r6_34 ) , .ZN( u1_uk_n1129 ) , .A2( u1_uk_n291 ) );
  OAI21_X1 u1_uk_U1111 (.ZN( u1_K16_39 ) , .B2( u1_uk_n1231 ) , .B1( u1_uk_n291 ) , .A( u1_uk_n990 ) );
  NAND2_X1 u1_uk_U1112 (.A1( u1_uk_K_r14_15 ) , .A2( u1_uk_n214 ) , .ZN( u1_uk_n990 ) );
  INV_X1 u1_uk_U1133 (.ZN( u1_K8_12 ) , .A( u1_uk_n1128 ) );
  AOI22_X1 u1_uk_U1134 (.B2( u1_uk_K_r6_3 ) , .A2( u1_uk_K_r6_53 ) , .ZN( u1_uk_n1128 ) , .B1( u1_uk_n164 ) , .A1( u1_uk_n220 ) );
  OAI22_X1 u1_uk_U114 (.ZN( u1_K12_5 ) , .A2( u1_uk_n1712 ) , .B2( u1_uk_n1738 ) , .A1( u1_uk_n213 ) , .B1( u1_uk_n99 ) );
  INV_X1 u1_uk_U1149 (.ZN( u1_K7_13 ) , .A( u1_uk_n1106 ) );
  AOI22_X1 u1_uk_U1150 (.B2( u1_uk_K_r5_26 ) , .A2( u1_uk_K_r5_48 ) , .ZN( u1_uk_n1106 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n217 ) );
  INV_X1 u1_uk_U1159 (.ZN( u1_K8_15 ) , .A( u1_uk_n1130 ) );
  AOI22_X1 u1_uk_U1160 (.B2( u1_uk_K_r6_10 ) , .A2( u1_uk_K_r6_17 ) , .A1( u1_uk_n110 ) , .ZN( u1_uk_n1130 ) , .B1( u1_uk_n207 ) );
  INV_X1 u1_uk_U1169 (.ZN( u1_K12_1 ) , .A( u1_uk_n515 ) );
  OAI22_X1 u1_uk_U118 (.ZN( u1_K2_5 ) , .B2( u1_uk_n1274 ) , .A2( u1_uk_n1277 ) , .A1( u1_uk_n291 ) , .B1( u1_uk_n31 ) );
  OAI22_X1 u1_uk_U123 (.ZN( u1_K16_47 ) , .B2( u1_uk_n1218 ) , .A2( u1_uk_n1222 ) , .A1( u1_uk_n240 ) , .B1( u1_uk_n60 ) );
  OAI22_X1 u1_uk_U130 (.ZN( u1_K7_47 ) , .A2( u1_uk_n1486 ) , .B2( u1_uk_n1500 ) , .A1( u1_uk_n222 ) , .B1( u1_uk_n92 ) );
  OAI22_X1 u1_uk_U133 (.ZN( u1_K5_47 ) , .B2( u1_uk_n1395 ) , .A2( u1_uk_n1419 ) , .A1( u1_uk_n208 ) , .B1( u1_uk_n93 ) );
  INV_X1 u1_uk_U14 (.ZN( u1_uk_n100 ) , .A( u1_uk_n213 ) );
  OAI22_X1 u1_uk_U143 (.ZN( u1_K7_15 ) , .A2( u1_uk_n1484 ) , .B2( u1_uk_n1524 ) , .A1( u1_uk_n252 ) , .B1( u1_uk_n92 ) );
  OAI21_X1 u1_uk_U157 (.ZN( u1_K15_15 ) , .B2( u1_uk_n1873 ) , .B1( u1_uk_n222 ) , .A( u1_uk_n967 ) );
  NAND2_X1 u1_uk_U158 (.A1( u1_uk_K_r13_19 ) , .A2( u1_uk_n294 ) , .ZN( u1_uk_n967 ) );
  INV_X1 u1_uk_U17 (.ZN( u1_uk_n110 ) , .A( u1_uk_n209 ) );
  OAI22_X1 u1_uk_U174 (.ZN( u1_K5_30 ) , .B2( u1_uk_n1408 ) , .A2( u1_uk_n1425 ) , .A1( u1_uk_n147 ) , .B1( u1_uk_n297 ) );
  OAI21_X1 u1_uk_U186 (.ZN( u1_K16_30 ) , .B2( u1_uk_n1256 ) , .B1( u1_uk_n222 ) , .A( u1_uk_n987 ) );
  NAND2_X1 u1_uk_U187 (.A1( u1_uk_K_r14_45 ) , .A2( u1_uk_n279 ) , .ZN( u1_uk_n987 ) );
  OAI22_X1 u1_uk_U208 (.ZN( u1_K15_24 ) , .A1( u1_uk_n146 ) , .A2( u1_uk_n1846 ) , .B2( u1_uk_n1864 ) , .B1( u1_uk_n238 ) );
  INV_X1 u1_uk_U215 (.ZN( u1_K15_30 ) , .A( u1_uk_n970 ) );
  AOI22_X1 u1_uk_U216 (.B2( u1_uk_K_r13_0 ) , .A2( u1_uk_K_r13_38 ) , .B1( u1_uk_n164 ) , .A1( u1_uk_n240 ) , .ZN( u1_uk_n970 ) );
  INV_X1 u1_uk_U218 (.ZN( u1_K4_31 ) , .A( u1_uk_n1063 ) );
  AOI22_X1 u1_uk_U219 (.B2( u1_uk_K_r2_31 ) , .A2( u1_uk_K_r2_49 ) , .ZN( u1_uk_n1063 ) , .B1( u1_uk_n147 ) , .A1( u1_uk_n257 ) );
  OAI22_X1 u1_uk_U222 (.ZN( u1_K16_31 ) , .A2( u1_uk_n1222 ) , .B2( u1_uk_n1225 ) , .A1( u1_uk_n141 ) , .B1( u1_uk_n257 ) );
  INV_X1 u1_uk_U229 (.ZN( u1_K11_39 ) , .A( u1_uk_n460 ) );
  AOI22_X1 u1_uk_U230 (.B2( u1_uk_K_r9_30 ) , .A2( u1_uk_K_r9_7 ) , .B1( u1_uk_n182 ) , .A1( u1_uk_n292 ) , .ZN( u1_uk_n460 ) );
  OAI22_X1 u1_uk_U251 (.ZN( u1_K16_48 ) , .B2( u1_uk_n1230 ) , .A2( u1_uk_n1238 ) , .A1( u1_uk_n213 ) , .B1( u1_uk_n60 ) );
  OAI21_X1 u1_uk_U252 (.ZN( u1_K16_44 ) , .B2( u1_uk_n1246 ) , .B1( u1_uk_n155 ) , .A( u1_uk_n994 ) );
  NAND2_X1 u1_uk_U253 (.A1( u1_uk_K_r14_43 ) , .A2( u1_uk_n94 ) , .ZN( u1_uk_n994 ) );
  OAI22_X1 u1_uk_U257 (.ZN( u1_K5_44 ) , .B2( u1_uk_n1419 ) , .A2( u1_uk_n1425 ) , .A1( u1_uk_n252 ) , .B1( u1_uk_n93 ) );
  OAI22_X1 u1_uk_U258 (.ZN( u1_K5_48 ) , .B2( u1_uk_n1407 ) , .A2( u1_uk_n1414 ) , .A1( u1_uk_n209 ) , .B1( u1_uk_n93 ) );
  INV_X1 u1_uk_U276 (.ZN( u1_K9_48 ) , .A( u1_uk_n1170 ) );
  AOI22_X1 u1_uk_U277 (.B2( u1_uk_K_r7_16 ) , .A2( u1_uk_K_r7_9 ) , .A1( u1_uk_n110 ) , .ZN( u1_uk_n1170 ) , .B1( u1_uk_n251 ) );
  OAI22_X1 u1_uk_U278 (.ZN( u1_K7_44 ) , .A1( u1_uk_n141 ) , .B2( u1_uk_n1489 ) , .A2( u1_uk_n1510 ) , .B1( u1_uk_n214 ) );
  OAI22_X1 u1_uk_U279 (.ZN( u1_K7_48 ) , .A1( u1_uk_n141 ) , .B2( u1_uk_n1501 ) , .A2( u1_uk_n1521 ) , .B1( u1_uk_n291 ) );
  OAI22_X1 u1_uk_U289 (.ZN( u1_K8_6 ) , .B2( u1_uk_n1544 ) , .A2( u1_uk_n1549 ) , .A1( u1_uk_n207 ) , .B1( u1_uk_n92 ) );
  OAI22_X1 u1_uk_U297 (.ZN( u1_K2_6 ) , .B2( u1_uk_n1279 ) , .A2( u1_uk_n1300 ) , .A1( u1_uk_n146 ) , .B1( u1_uk_n188 ) );
  INV_X1 u1_uk_U299 (.ZN( u1_K15_8 ) , .A( u1_uk_n976 ) );
  AOI22_X1 u1_uk_U300 (.B2( u1_uk_K_r13_13 ) , .A2( u1_uk_K_r13_17 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n231 ) , .ZN( u1_uk_n976 ) );
  OAI22_X1 u1_uk_U302 (.ZN( u1_K8_8 ) , .B2( u1_uk_n1558 ) , .A2( u1_uk_n1564 ) , .A1( u1_uk_n220 ) , .B1( u1_uk_n94 ) );
  INV_X1 u1_uk_U303 (.ZN( u1_K7_8 ) , .A( u1_uk_n1126 ) );
  AOI22_X1 u1_uk_U304 (.B2( u1_uk_K_r5_26 ) , .A2( u1_uk_K_r5_4 ) , .A1( u1_uk_n110 ) , .ZN( u1_uk_n1126 ) , .B1( u1_uk_n223 ) );
  INV_X1 u1_uk_U319 (.ZN( u1_K15_26 ) , .A( u1_uk_n969 ) );
  AOI22_X1 u1_uk_U320 (.B2( u1_uk_K_r13_38 ) , .A2( u1_uk_K_r13_44 ) , .B1( u1_uk_n162 ) , .A1( u1_uk_n291 ) , .ZN( u1_uk_n969 ) );
  OAI22_X1 u1_uk_U327 (.ZN( u1_K5_26 ) , .A2( u1_uk_n1396 ) , .B2( u1_uk_n1406 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n252 ) );
  OAI22_X1 u1_uk_U329 (.ZN( u1_K16_26 ) , .B2( u1_uk_n1241 ) , .A2( u1_uk_n1255 ) , .A1( u1_uk_n145 ) , .B1( u1_uk_n279 ) );
  OAI22_X1 u1_uk_U335 (.ZN( u1_K5_46 ) , .B2( u1_uk_n1394 ) , .A1( u1_uk_n141 ) , .A2( u1_uk_n1431 ) , .B1( u1_uk_n240 ) );
  OAI22_X1 u1_uk_U346 (.ZN( u1_K15_4 ) , .A1( u1_uk_n145 ) , .B2( u1_uk_n1850 ) , .A2( u1_uk_n1880 ) , .B1( u1_uk_n257 ) );
  INV_X1 u1_uk_U35 (.ZN( u1_uk_n187 ) , .A( u1_uk_n213 ) );
  OAI22_X1 u1_uk_U356 (.ZN( u1_K2_4 ) , .B2( u1_uk_n1268 ) , .A2( u1_uk_n1297 ) , .A1( u1_uk_n250 ) , .B1( u1_uk_n31 ) );
  OAI22_X1 u1_uk_U358 (.ZN( u1_K16_40 ) , .A1( u1_uk_n110 ) , .B2( u1_uk_n1218 ) , .A2( u1_uk_n1256 ) , .B1( u1_uk_n257 ) );
  INV_X1 u1_uk_U359 (.ZN( u1_K12_4 ) , .A( u1_uk_n656 ) );
  AOI22_X1 u1_uk_U360 (.B2( u1_uk_K_r10_27 ) , .A2( u1_uk_K_r10_4 ) , .A1( u1_uk_n298 ) , .B1( u1_uk_n31 ) , .ZN( u1_uk_n656 ) );
  OAI21_X1 u1_uk_U367 (.ZN( u1_K9_46 ) , .B1( u1_uk_n11 ) , .A( u1_uk_n1169 ) , .B2( u1_uk_n1607 ) );
  NAND2_X1 u1_uk_U368 (.A1( u1_uk_K_r7_37 ) , .ZN( u1_uk_n1169 ) , .A2( u1_uk_n31 ) );
  INV_X1 u1_uk_U369 (.ZN( u1_K7_46 ) , .A( u1_uk_n1124 ) );
  AOI22_X1 u1_uk_U370 (.B2( u1_uk_K_r5_23 ) , .A2( u1_uk_K_r5_31 ) , .A1( u1_uk_n110 ) , .ZN( u1_uk_n1124 ) , .B1( u1_uk_n208 ) );
  OAI22_X1 u1_uk_U373 (.ZN( u1_K11_40 ) , .B1( u1_uk_n102 ) , .A2( u1_uk_n1664 ) , .B2( u1_uk_n1672 ) , .A1( u1_uk_n250 ) );
  OAI22_X1 u1_uk_U375 (.ZN( u1_K7_40 ) , .A2( u1_uk_n1482 ) , .B2( u1_uk_n1494 ) , .A1( u1_uk_n188 ) , .B1( u1_uk_n92 ) );
  OAI22_X1 u1_uk_U376 (.ZN( u1_K4_40 ) , .B1( u1_uk_n118 ) , .B2( u1_uk_n1372 ) , .A2( u1_uk_n1382 ) , .A1( u1_uk_n214 ) );
  OAI22_X1 u1_uk_U390 (.ZN( u1_K15_28 ) , .A1( u1_uk_n148 ) , .B2( u1_uk_n1855 ) , .A2( u1_uk_n1883 ) , .B1( u1_uk_n209 ) );
  OAI22_X1 u1_uk_U395 (.ZN( u1_K5_28 ) , .B2( u1_uk_n1396 ) , .A2( u1_uk_n1400 ) , .B1( u1_uk_n148 ) , .A1( u1_uk_n223 ) );
  OAI22_X1 u1_uk_U399 (.ZN( u1_K2_1 ) , .B2( u1_uk_n1284 ) , .A2( u1_uk_n1305 ) , .A1( u1_uk_n142 ) , .B1( u1_uk_n230 ) );
  INV_X1 u1_uk_U4 (.ZN( u1_uk_n164 ) , .A( u1_uk_n203 ) );
  OAI22_X1 u1_uk_U408 (.ZN( u1_K8_16 ) , .B2( u1_uk_n1536 ) , .A2( u1_uk_n1544 ) , .A1( u1_uk_n202 ) , .B1( u1_uk_n94 ) );
  OAI21_X1 u1_uk_U409 (.ZN( u1_K7_16 ) , .A( u1_uk_n1107 ) , .B2( u1_uk_n1526 ) , .B1( u1_uk_n161 ) );
  BUF_X1 u1_uk_U41 (.Z( u1_uk_n203 ) , .A( u1_uk_n291 ) );
  NAND2_X1 u1_uk_U410 (.A1( u1_uk_K_r5_32 ) , .A2( u1_uk_n11 ) , .ZN( u1_uk_n1107 ) );
  OAI21_X1 u1_uk_U416 (.ZN( u1_K15_9 ) , .B1( u1_uk_n155 ) , .B2( u1_uk_n1873 ) , .A( u1_uk_n977 ) );
  NAND2_X1 u1_uk_U417 (.A1( u1_uk_K_r13_4 ) , .A2( u1_uk_n63 ) , .ZN( u1_uk_n977 ) );
  OAI22_X1 u1_uk_U423 (.ZN( u1_K8_9 ) , .A1( u1_uk_n109 ) , .A2( u1_uk_n1532 ) , .B2( u1_uk_n1538 ) , .B1( u1_uk_n251 ) );
  OAI22_X1 u1_uk_U433 (.ZN( u1_K15_16 ) , .B1( u1_uk_n100 ) , .B2( u1_uk_n1859 ) , .A2( u1_uk_n1874 ) , .A1( u1_uk_n207 ) );
  OAI22_X1 u1_uk_U440 (.ZN( u1_K4_37 ) , .B2( u1_uk_n1361 ) , .A2( u1_uk_n1375 ) , .A1( u1_uk_n163 ) , .B1( u1_uk_n209 ) );
  OAI22_X1 u1_uk_U451 (.ZN( u1_K7_9 ) , .B2( u1_uk_n1491 ) , .A2( u1_uk_n1498 ) , .A1( u1_uk_n297 ) , .B1( u1_uk_n92 ) );
  OAI22_X1 u1_uk_U452 (.ZN( u1_K15_1 ) , .B2( u1_uk_n1868 ) , .A2( u1_uk_n1887 ) , .A1( u1_uk_n271 ) , .B1( u1_uk_n99 ) );
  INV_X1 u1_uk_U453 (.ZN( u1_K16_37 ) , .A( u1_uk_n989 ) );
  AOI22_X1 u1_uk_U454 (.B2( u1_uk_K_r14_2 ) , .A2( u1_uk_K_r14_50 ) , .B1( u1_uk_n163 ) , .A1( u1_uk_n213 ) , .ZN( u1_uk_n989 ) );
  OAI22_X1 u1_uk_U455 (.ZN( u1_K16_33 ) , .B2( u1_uk_n1250 ) , .A2( u1_uk_n1255 ) , .A1( u1_uk_n188 ) , .B1( u1_uk_n63 ) );
  OAI22_X1 u1_uk_U469 (.ZN( u1_K4_33 ) , .B1( u1_uk_n117 ) , .B2( u1_uk_n1349 ) , .A2( u1_uk_n1356 ) , .A1( u1_uk_n250 ) );
  OAI21_X1 u1_uk_U473 (.ZN( u1_K11_37 ) , .B2( u1_uk_n1694 ) , .A( u1_uk_n456 ) , .B1( u1_uk_n92 ) );
  NAND2_X1 u1_uk_U474 (.A1( u1_uk_K_r9_38 ) , .ZN( u1_uk_n456 ) , .A2( u1_uk_n63 ) );
  OAI22_X1 u1_uk_U491 (.ZN( u1_K15_29 ) , .A1( u1_uk_n148 ) , .A2( u1_uk_n1849 ) , .B2( u1_uk_n1867 ) , .B1( u1_uk_n298 ) );
  OAI22_X1 u1_uk_U494 (.ZN( u1_K5_29 ) , .B2( u1_uk_n1407 ) , .A1( u1_uk_n142 ) , .A2( u1_uk_n1426 ) , .B1( u1_uk_n277 ) );
  INV_X1 u1_uk_U495 (.ZN( u1_K16_29 ) , .A( u1_uk_n985 ) );
  AOI22_X1 u1_uk_U496 (.B2( u1_uk_K_r14_16 ) , .A2( u1_uk_K_r14_23 ) , .A1( u1_uk_n110 ) , .B1( u1_uk_n277 ) , .ZN( u1_uk_n985 ) );
  OAI22_X1 u1_uk_U508 (.ZN( u1_K2_2 ) , .B2( u1_uk_n1273 ) , .A2( u1_uk_n1305 ) , .A1( u1_uk_n271 ) , .B1( u1_uk_n92 ) );
  OAI21_X1 u1_uk_U509 (.ZN( u1_K8_2 ) , .A( u1_uk_n1135 ) , .B2( u1_uk_n1545 ) , .B1( u1_uk_n155 ) );
  BUF_X1 u1_uk_U51 (.Z( u1_uk_n207 ) , .A( u1_uk_n291 ) );
  NAND2_X1 u1_uk_U510 (.A1( u1_uk_K_r6_27 ) , .ZN( u1_uk_n1135 ) , .A2( u1_uk_n27 ) );
  OAI21_X1 u1_uk_U523 (.ZN( u1_K8_17 ) , .A( u1_uk_n1131 ) , .B2( u1_uk_n1552 ) , .B1( u1_uk_n298 ) );
  NAND2_X1 u1_uk_U524 (.A1( u1_uk_K_r6_26 ) , .ZN( u1_uk_n1131 ) , .A2( u1_uk_n242 ) );
  OAI22_X1 u1_uk_U525 (.ZN( u1_K7_17 ) , .B2( u1_uk_n1488 ) , .A2( u1_uk_n1518 ) , .A1( u1_uk_n188 ) , .B1( u1_uk_n92 ) );
  OAI22_X1 u1_uk_U529 (.ZN( u1_K15_12 ) , .A1( u1_uk_n147 ) , .A2( u1_uk_n1845 ) , .B2( u1_uk_n1863 ) , .B1( u1_uk_n240 ) );
  OAI22_X1 u1_uk_U533 (.ZN( u1_K15_2 ) , .A1( u1_uk_n148 ) , .B2( u1_uk_n1858 ) , .A2( u1_uk_n1887 ) , .B1( u1_uk_n213 ) );
  INV_X1 u1_uk_U538 (.ZN( u1_K7_12 ) , .A( u1_uk_n1105 ) );
  AOI22_X1 u1_uk_U539 (.B2( u1_uk_K_r5_17 ) , .A2( u1_uk_K_r5_39 ) , .ZN( u1_uk_n1105 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n242 ) );
  OAI22_X1 u1_uk_U551 (.ZN( u1_K15_17 ) , .A1( u1_uk_n117 ) , .A2( u1_uk_n1844 ) , .B2( u1_uk_n1862 ) , .B1( u1_uk_n242 ) );
  OAI22_X1 u1_uk_U562 (.ZN( u1_K16_36 ) , .B2( u1_uk_n1233 ) , .A2( u1_uk_n1240 ) , .A1( u1_uk_n202 ) , .B1( u1_uk_n63 ) );
  OAI22_X1 u1_uk_U564 (.ZN( u1_K11_38 ) , .B2( u1_uk_n1670 ) , .A2( u1_uk_n1678 ) , .A1( u1_uk_n182 ) , .B1( u1_uk_n294 ) );
  BUF_X1 u1_uk_U58 (.Z( u1_uk_n291 ) , .A( u1_uk_n294 ) );
  OAI21_X1 u1_uk_U580 (.ZN( u1_K15_10 ) , .B2( u1_uk_n1869 ) , .B1( u1_uk_n94 ) , .A( u1_uk_n964 ) );
  NAND2_X1 u1_uk_U581 (.A1( u1_uk_K_r13_55 ) , .A2( u1_uk_n92 ) , .ZN( u1_uk_n964 ) );
  OAI22_X1 u1_uk_U589 (.ZN( u1_K8_10 ) , .B2( u1_uk_n1549 ) , .A2( u1_uk_n1551 ) , .A1( u1_uk_n277 ) , .B1( u1_uk_n92 ) );
  OAI22_X1 u1_uk_U612 (.ZN( u1_K16_35 ) , .B2( u1_uk_n1238 ) , .A2( u1_uk_n1245 ) , .A1( u1_uk_n238 ) , .B1( u1_uk_n63 ) );
  OAI22_X1 u1_uk_U629 (.ZN( u1_K4_35 ) , .B2( u1_uk_n1361 ) , .A2( u1_uk_n1390 ) , .B1( u1_uk_n142 ) , .A1( u1_uk_n271 ) );
  OAI21_X1 u1_uk_U635 (.ZN( u1_K15_11 ) , .B2( u1_uk_n1880 ) , .B1( u1_uk_n250 ) , .A( u1_uk_n965 ) );
  NAND2_X1 u1_uk_U636 (.A1( u1_uk_K_r13_25 ) , .A2( u1_uk_n230 ) , .ZN( u1_uk_n965 ) );
  BUF_X1 u1_uk_U64 (.Z( u1_uk_n294 ) , .A( u1_uk_n298 ) );
  OAI21_X1 u1_uk_U645 (.ZN( u1_K8_11 ) , .A( u1_uk_n1127 ) , .B2( u1_uk_n1565 ) , .B1( u1_uk_n94 ) );
  NAND2_X1 u1_uk_U646 (.A1( u1_uk_K_r6_55 ) , .ZN( u1_uk_n1127 ) , .A2( u1_uk_n147 ) );
  OAI22_X1 u1_uk_U647 (.ZN( u1_K7_11 ) , .A1( u1_uk_n129 ) , .B2( u1_uk_n1488 ) , .A2( u1_uk_n1505 ) , .B1( u1_uk_n203 ) );
  BUF_X1 u1_uk_U65 (.Z( u1_uk_n297 ) , .A( u1_uk_n298 ) );
  OAI22_X1 u1_uk_U652 (.ZN( u1_K16_45 ) , .B2( u1_uk_n1247 ) , .A2( u1_uk_n1250 ) , .A1( u1_uk_n294 ) , .B1( u1_uk_n63 ) );
  INV_X1 u1_uk_U66 (.A( n116 ) , .ZN( u1_uk_n298 ) );
  INV_X1 u1_uk_U665 (.ZN( u1_K16_43 ) , .A( u1_uk_n993 ) );
  AOI22_X1 u1_uk_U666 (.B2( u1_uk_K_r14_16 ) , .A2( u1_uk_K_r14_9 ) , .B1( u1_uk_n164 ) , .A1( u1_uk_n220 ) , .ZN( u1_uk_n993 ) );
  INV_X1 u1_uk_U667 (.ZN( u1_K5_43 ) , .A( u1_uk_n1083 ) );
  AOI22_X1 u1_uk_U668 (.B2( u1_uk_K_r3_15 ) , .A2( u1_uk_K_r3_38 ) , .ZN( u1_uk_n1083 ) , .B1( u1_uk_n163 ) , .A1( u1_uk_n217 ) );
  INV_X1 u1_uk_U67 (.ZN( u1_K16_34 ) , .A( u1_uk_n988 ) );
  OAI22_X1 u1_uk_U678 (.ZN( u1_K9_43 ) , .A1( u1_uk_n11 ) , .B2( u1_uk_n1588 ) , .A2( u1_uk_n1595 ) , .B1( u1_uk_n297 ) );
  OAI22_X1 u1_uk_U679 (.ZN( u1_K9_45 ) , .B2( u1_uk_n1571 ) , .A2( u1_uk_n1612 ) , .A1( u1_uk_n191 ) , .B1( u1_uk_n93 ) );
  AOI22_X1 u1_uk_U68 (.A1( n116 ) , .B2( u1_uk_K_r14_2 ) , .A2( u1_uk_K_r14_9 ) , .B1( u1_uk_n213 ) , .ZN( u1_uk_n988 ) );
  OAI22_X1 u1_uk_U680 (.ZN( u1_K7_43 ) , .A1( u1_uk_n141 ) , .A2( u1_uk_n1485 ) , .B2( u1_uk_n1514 ) , .B1( u1_uk_n207 ) );
  OAI21_X1 u1_uk_U688 (.ZN( u1_K15_25 ) , .B2( u1_uk_n1876 ) , .B1( u1_uk_n223 ) , .A( u1_uk_n968 ) );
  NAND2_X1 u1_uk_U689 (.A1( u1_uk_K_r13_22 ) , .A2( u1_uk_n213 ) , .ZN( u1_uk_n968 ) );
  OAI22_X1 u1_uk_U694 (.ZN( u1_K16_25 ) , .B2( u1_uk_n1239 ) , .A2( u1_uk_n1246 ) , .A1( u1_uk_n294 ) , .B1( u1_uk_n63 ) );
  OAI22_X1 u1_uk_U701 (.ZN( u1_K15_7 ) , .B2( u1_uk_n1853 ) , .A2( u1_uk_n1869 ) , .A1( u1_uk_n191 ) , .B1( u1_uk_n83 ) );
  INV_X1 u1_uk_U703 (.ZN( u1_K12_3 ) , .A( u1_uk_n601 ) );
  AOI22_X1 u1_uk_U704 (.B2( u1_uk_K_r10_18 ) , .A2( u1_uk_K_r10_27 ) , .B1( u1_uk_n129 ) , .A1( u1_uk_n231 ) , .ZN( u1_uk_n601 ) );
  INV_X1 u1_uk_U705 (.ZN( u1_K8_3 ) , .A( u1_uk_n1140 ) );
  AOI22_X1 u1_uk_U706 (.B2( u1_uk_K_r6_10 ) , .A2( u1_uk_K_r6_3 ) , .ZN( u1_uk_n1140 ) , .B1( u1_uk_n163 ) , .A1( u1_uk_n294 ) );
  OAI22_X1 u1_uk_U717 (.ZN( u1_K12_2 ) , .B1( u1_uk_n100 ) , .A2( u1_uk_n1711 ) , .B2( u1_uk_n1716 ) , .A1( u1_uk_n271 ) );
  OAI22_X1 u1_uk_U722 (.ZN( u1_K4_32 ) , .A1( u1_uk_n110 ) , .A2( u1_uk_n1356 ) , .B2( u1_uk_n1380 ) , .B1( u1_uk_n242 ) );
  OAI22_X1 u1_uk_U723 (.ZN( u1_K16_32 ) , .B2( u1_uk_n1231 ) , .A2( u1_uk_n1239 ) , .A1( u1_uk_n292 ) , .B1( u1_uk_n63 ) );
  OAI22_X1 u1_uk_U735 (.ZN( u1_K11_42 ) , .A1( u1_uk_n164 ) , .B2( u1_uk_n1694 ) , .A2( u1_uk_n1702 ) , .B1( u1_uk_n220 ) );
  OAI22_X1 u1_uk_U737 (.ZN( u1_K4_42 ) , .B2( u1_uk_n1360 ) , .A2( u1_uk_n1367 ) , .B1( u1_uk_n141 ) , .A1( u1_uk_n251 ) );
  INV_X1 u1_uk_U744 (.ZN( u1_K7_42 ) , .A( u1_uk_n1123 ) );
  AOI22_X1 u1_uk_U745 (.B2( u1_uk_K_r5_1 ) , .A2( u1_uk_K_r5_36 ) , .A1( u1_uk_n110 ) , .ZN( u1_uk_n1123 ) , .B1( u1_uk_n297 ) );
  OAI22_X1 u1_uk_U754 (.ZN( u1_K16_27 ) , .B2( u1_uk_n1225 ) , .A2( u1_uk_n1230 ) , .A1( u1_uk_n240 ) , .B1( u1_uk_n63 ) );
  OAI22_X1 u1_uk_U757 (.ZN( u1_K8_13 ) , .A1( u1_uk_n129 ) , .A2( u1_uk_n1531 ) , .B2( u1_uk_n1537 ) , .B1( u1_uk_n252 ) );
  OAI22_X1 u1_uk_U774 (.ZN( u1_K15_21 ) , .B1( u1_uk_n100 ) , .A2( u1_uk_n1846 ) , .B2( u1_uk_n1850 ) , .A1( u1_uk_n223 ) );
  OAI22_X1 u1_uk_U777 (.ZN( u1_K15_27 ) , .A1( u1_uk_n148 ) , .A2( u1_uk_n1847 ) , .B2( u1_uk_n1865 ) , .B1( u1_uk_n214 ) );
  INV_X1 u1_uk_U790 (.ZN( u1_K5_27 ) , .A( u1_uk_n1076 ) );
  AOI22_X1 u1_uk_U791 (.B2( u1_uk_K_r3_15 ) , .A2( u1_uk_K_r3_51 ) , .ZN( u1_uk_n1076 ) , .B1( u1_uk_n240 ) , .A1( u1_uk_n83 ) );
  INV_X1 u1_uk_U8 (.A( u1_uk_n203 ) , .ZN( u1_uk_n63 ) );
  OAI22_X1 u1_uk_U81 (.ZN( u1_K4_34 ) , .A1( u1_uk_n117 ) , .B2( u1_uk_n1366 ) , .A2( u1_uk_n1382 ) , .B1( u1_uk_n202 ) );
  OAI22_X1 u1_uk_U817 (.ZN( u1_K7_18 ) , .A2( u1_uk_n1483 ) , .B2( u1_uk_n1496 ) , .A1( u1_uk_n230 ) , .B1( u1_uk_n92 ) );
  OAI21_X1 u1_uk_U818 (.ZN( u1_K8_18 ) , .A( u1_uk_n1132 ) , .B1( u1_uk_n155 ) , .B2( u1_uk_n1557 ) );
  NAND2_X1 u1_uk_U819 (.A1( u1_uk_K_r6_46 ) , .ZN( u1_uk_n1132 ) , .A2( u1_uk_n146 ) );
  OAI22_X1 u1_uk_U824 (.ZN( u1_K15_18 ) , .A1( u1_uk_n109 ) , .B2( u1_uk_n1852 ) , .A2( u1_uk_n1882 ) , .B1( u1_uk_n242 ) );
  OAI22_X1 u1_uk_U829 (.ZN( u1_K15_20 ) , .B1( u1_uk_n100 ) , .A2( u1_uk_n1845 ) , .B2( u1_uk_n1874 ) , .A1( u1_uk_n298 ) );
  OAI22_X1 u1_uk_U845 (.ZN( u1_K15_6 ) , .B2( u1_uk_n1864 ) , .A2( u1_uk_n1882 ) , .A1( u1_uk_n257 ) , .B1( u1_uk_n83 ) );
  OAI22_X1 u1_uk_U850 (.ZN( u1_K15_3 ) , .B2( u1_uk_n1852 ) , .A2( u1_uk_n1868 ) , .A1( u1_uk_n217 ) , .B1( u1_uk_n83 ) );
  AOI22_X1 u1_uk_U864 (.B2( u1_uk_K_r10_39 ) , .A2( u1_uk_K_r10_48 ) , .B1( u1_uk_n155 ) , .A1( u1_uk_n213 ) , .ZN( u1_uk_n515 ) );
  OAI22_X1 u1_uk_U870 (.ZN( u1_K15_22 ) , .B2( u1_uk_n1858 ) , .A2( u1_uk_n1872 ) , .A1( u1_uk_n209 ) , .B1( u1_uk_n99 ) );
  OAI22_X1 u1_uk_U872 (.ZN( u1_K15_23 ) , .B2( u1_uk_n1863 ) , .A2( u1_uk_n1881 ) , .A1( u1_uk_n251 ) , .B1( u1_uk_n99 ) );
  OAI22_X1 u1_uk_U878 (.ZN( u1_K8_5 ) , .B1( u1_uk_n102 ) , .B2( u1_uk_n1564 ) , .A2( u1_uk_n1570 ) , .A1( u1_uk_n294 ) );
  OAI22_X1 u1_uk_U882 (.ZN( u1_K7_10 ) , .B1( u1_uk_n147 ) , .B2( u1_uk_n1487 ) , .A2( u1_uk_n1517 ) , .A1( u1_uk_n202 ) );
  OAI22_X1 u1_uk_U890 (.ZN( u1_K8_1 ) , .B1( u1_uk_n146 ) , .A2( u1_uk_n1532 ) , .B2( u1_uk_n1548 ) , .A1( u1_uk_n214 ) );
  OAI22_X1 u1_uk_U897 (.ZN( u1_K7_14 ) , .B2( u1_uk_n1492 ) , .A2( u1_uk_n1527 ) , .A1( u1_uk_n202 ) , .B1( u1_uk_n92 ) );
  INV_X1 u1_uk_U9 (.A( u1_uk_n209 ) , .ZN( u1_uk_n94 ) );
  OAI22_X1 u1_uk_U901 (.ZN( u1_K15_13 ) , .B1( u1_uk_n100 ) , .A2( u1_uk_n1844 ) , .B2( u1_uk_n1872 ) , .A1( u1_uk_n294 ) );
  OAI22_X1 u1_uk_U915 (.ZN( u1_K4_36 ) , .B2( u1_uk_n1376 ) , .A2( u1_uk_n1381 ) , .B1( u1_uk_n163 ) , .A1( u1_uk_n238 ) );
  OAI22_X1 u1_uk_U919 (.ZN( u1_K16_38 ) , .B2( u1_uk_n1240 ) , .A2( u1_uk_n1247 ) , .A1( u1_uk_n222 ) , .B1( u1_uk_n63 ) );
  OAI22_X1 u1_uk_U921 (.ZN( u1_K7_39 ) , .B2( u1_uk_n1516 ) , .A2( u1_uk_n1523 ) , .A1( u1_uk_n203 ) , .B1( u1_uk_n92 ) );
  OAI22_X1 u1_uk_U924 (.ZN( u1_K4_39 ) , .B2( u1_uk_n1351 ) , .A2( u1_uk_n1372 ) , .B1( u1_uk_n182 ) , .A1( u1_uk_n257 ) );
  OAI22_X1 u1_uk_U930 (.ZN( u1_K9_47 ) , .B2( u1_uk_n1606 ) , .A2( u1_uk_n1613 ) , .A1( u1_uk_n163 ) , .B1( u1_uk_n209 ) );
  OAI22_X1 u1_uk_U944 (.ZN( u1_K16_46 ) , .B2( u1_uk_n1219 ) , .A2( u1_uk_n1253 ) , .A1( u1_uk_n161 ) , .B1( u1_uk_n208 ) );
  OAI21_X1 u1_uk_U95 (.ZN( u1_K11_41 ) , .B2( u1_uk_n1702 ) , .B1( u1_uk_n217 ) , .A( u1_uk_n467 ) );
  NAND2_X1 u1_uk_U96 (.A1( u1_uk_K_r9_31 ) , .A2( u1_uk_n203 ) , .ZN( u1_uk_n467 ) );
  OAI22_X1 u1_uk_U962 (.ZN( u1_K15_19 ) , .A1( u1_uk_n163 ) , .B2( u1_uk_n1851 ) , .A2( u1_uk_n1881 ) , .B1( u1_uk_n222 ) );
  OAI22_X1 u1_uk_U969 (.ZN( u1_K7_37 ) , .A1( u1_uk_n141 ) , .B2( u1_uk_n1499 ) , .A2( u1_uk_n1523 ) , .B1( u1_uk_n250 ) );
  OAI22_X1 u1_uk_U976 (.ZN( u1_K7_45 ) , .A1( u1_uk_n141 ) , .B2( u1_uk_n1490 ) , .A2( u1_uk_n1507 ) , .B1( u1_uk_n214 ) );
  OAI22_X1 u1_uk_U980 (.ZN( u1_K2_3 ) , .B2( u1_uk_n1269 ) , .A2( u1_uk_n1284 ) , .A1( u1_uk_n164 ) , .B1( u1_uk_n213 ) );
  OAI22_X1 u1_uk_U983 (.ZN( u1_K8_7 ) , .A2( u1_uk_n1530 ) , .B2( u1_uk_n1536 ) , .A1( u1_uk_n155 ) , .B1( u1_uk_n230 ) );
  OAI22_X1 u1_uk_U984 (.ZN( u1_K7_7 ) , .A1( u1_uk_n141 ) , .B2( u1_uk_n1496 ) , .A2( u1_uk_n1518 ) , .B1( u1_uk_n291 ) );
  OAI21_X1 u1_uk_U994 (.ZN( u1_K5_25 ) , .A( u1_uk_n1075 ) , .B2( u1_uk_n1413 ) , .B1( u1_uk_n162 ) );
  NAND2_X1 u1_uk_U995 (.A1( u1_uk_K_r3_35 ) , .ZN( u1_uk_n1075 ) , .A2( u1_uk_n63 ) );
  XOR2_X1 u2_U159 (.B( u2_L0_8 ) , .Z( u2_N39 ) , .A( u2_out1_8 ) );
  XOR2_X1 u2_U214 (.B( u2_L0_3 ) , .Z( u2_N34 ) , .A( u2_out1_3 ) );
  XOR2_X1 u2_U50 (.B( u2_L0_25 ) , .Z( u2_N56 ) , .A( u2_out1_25 ) );
  XOR2_X1 u2_U92 (.B( u2_L0_14 ) , .Z( u2_N45 ) , .A( u2_out1_14 ) );
  XOR2_X1 u2_u1_U26 (.B( u2_K2_30 ) , .A( u2_R0_21 ) , .Z( u2_u1_X_30 ) );
  XOR2_X1 u2_u1_U28 (.B( u2_K2_29 ) , .A( u2_R0_20 ) , .Z( u2_u1_X_29 ) );
  XOR2_X1 u2_u1_U29 (.B( u2_K2_28 ) , .A( u2_R0_19 ) , .Z( u2_u1_X_28 ) );
  XOR2_X1 u2_u1_U30 (.B( u2_K2_27 ) , .A( u2_R0_18 ) , .Z( u2_u1_X_27 ) );
  XOR2_X1 u2_u1_U31 (.B( u2_K2_26 ) , .A( u2_R0_17 ) , .Z( u2_u1_X_26 ) );
  XOR2_X1 u2_u1_U32 (.B( u2_K2_25 ) , .A( u2_R0_16 ) , .Z( u2_u1_X_25 ) );
  OAI22_X1 u2_u1_u4_U10 (.B2( u2_u1_u4_n135 ) , .ZN( u2_u1_u4_n137 ) , .B1( u2_u1_u4_n153 ) , .A1( u2_u1_u4_n155 ) , .A2( u2_u1_u4_n171 ) );
  AND3_X1 u2_u1_u4_U11 (.A2( u2_u1_u4_n134 ) , .ZN( u2_u1_u4_n135 ) , .A3( u2_u1_u4_n145 ) , .A1( u2_u1_u4_n157 ) );
  NAND2_X1 u2_u1_u4_U12 (.ZN( u2_u1_u4_n132 ) , .A2( u2_u1_u4_n170 ) , .A1( u2_u1_u4_n173 ) );
  AOI21_X1 u2_u1_u4_U13 (.B2( u2_u1_u4_n160 ) , .B1( u2_u1_u4_n161 ) , .ZN( u2_u1_u4_n162 ) , .A( u2_u1_u4_n170 ) );
  AOI21_X1 u2_u1_u4_U14 (.ZN( u2_u1_u4_n107 ) , .B2( u2_u1_u4_n143 ) , .A( u2_u1_u4_n174 ) , .B1( u2_u1_u4_n184 ) );
  AOI21_X1 u2_u1_u4_U15 (.B2( u2_u1_u4_n158 ) , .B1( u2_u1_u4_n159 ) , .ZN( u2_u1_u4_n163 ) , .A( u2_u1_u4_n174 ) );
  AOI21_X1 u2_u1_u4_U16 (.A( u2_u1_u4_n153 ) , .B2( u2_u1_u4_n154 ) , .B1( u2_u1_u4_n155 ) , .ZN( u2_u1_u4_n165 ) );
  AOI21_X1 u2_u1_u4_U17 (.A( u2_u1_u4_n156 ) , .B2( u2_u1_u4_n157 ) , .ZN( u2_u1_u4_n164 ) , .B1( u2_u1_u4_n184 ) );
  INV_X1 u2_u1_u4_U18 (.A( u2_u1_u4_n138 ) , .ZN( u2_u1_u4_n170 ) );
  AND2_X1 u2_u1_u4_U19 (.A2( u2_u1_u4_n120 ) , .ZN( u2_u1_u4_n155 ) , .A1( u2_u1_u4_n160 ) );
  INV_X1 u2_u1_u4_U20 (.A( u2_u1_u4_n156 ) , .ZN( u2_u1_u4_n175 ) );
  NAND2_X1 u2_u1_u4_U21 (.A2( u2_u1_u4_n118 ) , .ZN( u2_u1_u4_n131 ) , .A1( u2_u1_u4_n147 ) );
  NAND2_X1 u2_u1_u4_U22 (.A1( u2_u1_u4_n119 ) , .A2( u2_u1_u4_n120 ) , .ZN( u2_u1_u4_n130 ) );
  NAND2_X1 u2_u1_u4_U23 (.ZN( u2_u1_u4_n117 ) , .A2( u2_u1_u4_n118 ) , .A1( u2_u1_u4_n148 ) );
  NAND2_X1 u2_u1_u4_U24 (.ZN( u2_u1_u4_n129 ) , .A1( u2_u1_u4_n134 ) , .A2( u2_u1_u4_n148 ) );
  AND3_X1 u2_u1_u4_U25 (.A1( u2_u1_u4_n119 ) , .A2( u2_u1_u4_n143 ) , .A3( u2_u1_u4_n154 ) , .ZN( u2_u1_u4_n161 ) );
  AND2_X1 u2_u1_u4_U26 (.A1( u2_u1_u4_n145 ) , .A2( u2_u1_u4_n147 ) , .ZN( u2_u1_u4_n159 ) );
  OR3_X1 u2_u1_u4_U27 (.A3( u2_u1_u4_n114 ) , .A2( u2_u1_u4_n115 ) , .A1( u2_u1_u4_n116 ) , .ZN( u2_u1_u4_n136 ) );
  AOI21_X1 u2_u1_u4_U28 (.A( u2_u1_u4_n113 ) , .ZN( u2_u1_u4_n116 ) , .B2( u2_u1_u4_n173 ) , .B1( u2_u1_u4_n174 ) );
  AOI21_X1 u2_u1_u4_U29 (.ZN( u2_u1_u4_n115 ) , .B2( u2_u1_u4_n145 ) , .B1( u2_u1_u4_n146 ) , .A( u2_u1_u4_n156 ) );
  NOR2_X1 u2_u1_u4_U3 (.ZN( u2_u1_u4_n121 ) , .A1( u2_u1_u4_n181 ) , .A2( u2_u1_u4_n182 ) );
  OAI22_X1 u2_u1_u4_U30 (.ZN( u2_u1_u4_n114 ) , .A2( u2_u1_u4_n121 ) , .B1( u2_u1_u4_n160 ) , .B2( u2_u1_u4_n170 ) , .A1( u2_u1_u4_n171 ) );
  INV_X1 u2_u1_u4_U31 (.A( u2_u1_u4_n158 ) , .ZN( u2_u1_u4_n182 ) );
  INV_X1 u2_u1_u4_U32 (.ZN( u2_u1_u4_n181 ) , .A( u2_u1_u4_n96 ) );
  INV_X1 u2_u1_u4_U33 (.A( u2_u1_u4_n144 ) , .ZN( u2_u1_u4_n179 ) );
  INV_X1 u2_u1_u4_U34 (.A( u2_u1_u4_n157 ) , .ZN( u2_u1_u4_n178 ) );
  NAND2_X1 u2_u1_u4_U35 (.A2( u2_u1_u4_n154 ) , .A1( u2_u1_u4_n96 ) , .ZN( u2_u1_u4_n97 ) );
  INV_X1 u2_u1_u4_U36 (.ZN( u2_u1_u4_n186 ) , .A( u2_u1_u4_n95 ) );
  OAI221_X1 u2_u1_u4_U37 (.C1( u2_u1_u4_n134 ) , .B1( u2_u1_u4_n158 ) , .B2( u2_u1_u4_n171 ) , .C2( u2_u1_u4_n173 ) , .A( u2_u1_u4_n94 ) , .ZN( u2_u1_u4_n95 ) );
  AOI222_X1 u2_u1_u4_U38 (.B2( u2_u1_u4_n132 ) , .A1( u2_u1_u4_n138 ) , .C2( u2_u1_u4_n175 ) , .A2( u2_u1_u4_n179 ) , .C1( u2_u1_u4_n181 ) , .B1( u2_u1_u4_n185 ) , .ZN( u2_u1_u4_n94 ) );
  INV_X1 u2_u1_u4_U39 (.A( u2_u1_u4_n113 ) , .ZN( u2_u1_u4_n185 ) );
  INV_X1 u2_u1_u4_U4 (.A( u2_u1_u4_n117 ) , .ZN( u2_u1_u4_n184 ) );
  INV_X1 u2_u1_u4_U40 (.A( u2_u1_u4_n143 ) , .ZN( u2_u1_u4_n183 ) );
  NOR2_X1 u2_u1_u4_U41 (.ZN( u2_u1_u4_n138 ) , .A1( u2_u1_u4_n168 ) , .A2( u2_u1_u4_n169 ) );
  NOR2_X1 u2_u1_u4_U42 (.A1( u2_u1_u4_n150 ) , .A2( u2_u1_u4_n152 ) , .ZN( u2_u1_u4_n153 ) );
  NOR2_X1 u2_u1_u4_U43 (.A2( u2_u1_u4_n128 ) , .A1( u2_u1_u4_n138 ) , .ZN( u2_u1_u4_n156 ) );
  AOI22_X1 u2_u1_u4_U44 (.B2( u2_u1_u4_n122 ) , .A1( u2_u1_u4_n123 ) , .ZN( u2_u1_u4_n124 ) , .B1( u2_u1_u4_n128 ) , .A2( u2_u1_u4_n172 ) );
  NAND2_X1 u2_u1_u4_U45 (.A2( u2_u1_u4_n120 ) , .ZN( u2_u1_u4_n123 ) , .A1( u2_u1_u4_n161 ) );
  INV_X1 u2_u1_u4_U46 (.A( u2_u1_u4_n153 ) , .ZN( u2_u1_u4_n172 ) );
  AOI22_X1 u2_u1_u4_U47 (.B2( u2_u1_u4_n132 ) , .A2( u2_u1_u4_n133 ) , .ZN( u2_u1_u4_n140 ) , .A1( u2_u1_u4_n150 ) , .B1( u2_u1_u4_n179 ) );
  NAND2_X1 u2_u1_u4_U48 (.ZN( u2_u1_u4_n133 ) , .A2( u2_u1_u4_n146 ) , .A1( u2_u1_u4_n154 ) );
  NAND2_X1 u2_u1_u4_U49 (.A1( u2_u1_u4_n103 ) , .ZN( u2_u1_u4_n154 ) , .A2( u2_u1_u4_n98 ) );
  NOR4_X1 u2_u1_u4_U5 (.A4( u2_u1_u4_n106 ) , .A3( u2_u1_u4_n107 ) , .A2( u2_u1_u4_n108 ) , .A1( u2_u1_u4_n109 ) , .ZN( u2_u1_u4_n110 ) );
  NAND2_X1 u2_u1_u4_U50 (.A1( u2_u1_u4_n101 ) , .ZN( u2_u1_u4_n158 ) , .A2( u2_u1_u4_n99 ) );
  AOI21_X1 u2_u1_u4_U51 (.ZN( u2_u1_u4_n127 ) , .A( u2_u1_u4_n136 ) , .B2( u2_u1_u4_n150 ) , .B1( u2_u1_u4_n180 ) );
  INV_X1 u2_u1_u4_U52 (.A( u2_u1_u4_n160 ) , .ZN( u2_u1_u4_n180 ) );
  NAND2_X1 u2_u1_u4_U53 (.A2( u2_u1_u4_n104 ) , .A1( u2_u1_u4_n105 ) , .ZN( u2_u1_u4_n146 ) );
  NAND2_X1 u2_u1_u4_U54 (.A2( u2_u1_u4_n101 ) , .A1( u2_u1_u4_n102 ) , .ZN( u2_u1_u4_n160 ) );
  NAND2_X1 u2_u1_u4_U55 (.ZN( u2_u1_u4_n134 ) , .A1( u2_u1_u4_n98 ) , .A2( u2_u1_u4_n99 ) );
  NAND2_X1 u2_u1_u4_U56 (.A1( u2_u1_u4_n103 ) , .A2( u2_u1_u4_n104 ) , .ZN( u2_u1_u4_n143 ) );
  NAND2_X1 u2_u1_u4_U57 (.A2( u2_u1_u4_n105 ) , .ZN( u2_u1_u4_n145 ) , .A1( u2_u1_u4_n98 ) );
  NAND2_X1 u2_u1_u4_U58 (.A1( u2_u1_u4_n100 ) , .A2( u2_u1_u4_n105 ) , .ZN( u2_u1_u4_n120 ) );
  NAND2_X1 u2_u1_u4_U59 (.A1( u2_u1_u4_n102 ) , .A2( u2_u1_u4_n104 ) , .ZN( u2_u1_u4_n148 ) );
  AOI21_X1 u2_u1_u4_U6 (.ZN( u2_u1_u4_n106 ) , .B2( u2_u1_u4_n146 ) , .B1( u2_u1_u4_n158 ) , .A( u2_u1_u4_n170 ) );
  NAND2_X1 u2_u1_u4_U60 (.A2( u2_u1_u4_n100 ) , .A1( u2_u1_u4_n103 ) , .ZN( u2_u1_u4_n157 ) );
  INV_X1 u2_u1_u4_U61 (.A( u2_u1_u4_n150 ) , .ZN( u2_u1_u4_n173 ) );
  INV_X1 u2_u1_u4_U62 (.A( u2_u1_u4_n152 ) , .ZN( u2_u1_u4_n171 ) );
  NAND2_X1 u2_u1_u4_U63 (.A1( u2_u1_u4_n100 ) , .ZN( u2_u1_u4_n118 ) , .A2( u2_u1_u4_n99 ) );
  NAND2_X1 u2_u1_u4_U64 (.A2( u2_u1_u4_n100 ) , .A1( u2_u1_u4_n102 ) , .ZN( u2_u1_u4_n144 ) );
  NAND2_X1 u2_u1_u4_U65 (.A2( u2_u1_u4_n101 ) , .A1( u2_u1_u4_n105 ) , .ZN( u2_u1_u4_n96 ) );
  INV_X1 u2_u1_u4_U66 (.A( u2_u1_u4_n128 ) , .ZN( u2_u1_u4_n174 ) );
  NAND2_X1 u2_u1_u4_U67 (.A2( u2_u1_u4_n102 ) , .ZN( u2_u1_u4_n119 ) , .A1( u2_u1_u4_n98 ) );
  NAND2_X1 u2_u1_u4_U68 (.A2( u2_u1_u4_n101 ) , .A1( u2_u1_u4_n103 ) , .ZN( u2_u1_u4_n147 ) );
  NAND2_X1 u2_u1_u4_U69 (.A2( u2_u1_u4_n104 ) , .ZN( u2_u1_u4_n113 ) , .A1( u2_u1_u4_n99 ) );
  AOI21_X1 u2_u1_u4_U7 (.ZN( u2_u1_u4_n108 ) , .B2( u2_u1_u4_n134 ) , .B1( u2_u1_u4_n155 ) , .A( u2_u1_u4_n156 ) );
  NOR2_X1 u2_u1_u4_U70 (.A2( u2_u1_X_28 ) , .ZN( u2_u1_u4_n150 ) , .A1( u2_u1_u4_n168 ) );
  NOR2_X1 u2_u1_u4_U71 (.A2( u2_u1_X_29 ) , .ZN( u2_u1_u4_n152 ) , .A1( u2_u1_u4_n169 ) );
  NOR2_X1 u2_u1_u4_U72 (.A2( u2_u1_X_30 ) , .ZN( u2_u1_u4_n105 ) , .A1( u2_u1_u4_n176 ) );
  NOR2_X1 u2_u1_u4_U73 (.A2( u2_u1_X_26 ) , .ZN( u2_u1_u4_n100 ) , .A1( u2_u1_u4_n177 ) );
  NOR2_X1 u2_u1_u4_U74 (.A2( u2_u1_X_28 ) , .A1( u2_u1_X_29 ) , .ZN( u2_u1_u4_n128 ) );
  NOR2_X1 u2_u1_u4_U75 (.A2( u2_u1_X_27 ) , .A1( u2_u1_X_30 ) , .ZN( u2_u1_u4_n102 ) );
  NOR2_X1 u2_u1_u4_U76 (.A2( u2_u1_X_25 ) , .A1( u2_u1_X_26 ) , .ZN( u2_u1_u4_n98 ) );
  AND2_X1 u2_u1_u4_U77 (.A2( u2_u1_X_25 ) , .A1( u2_u1_X_26 ) , .ZN( u2_u1_u4_n104 ) );
  AND2_X1 u2_u1_u4_U78 (.A1( u2_u1_X_30 ) , .A2( u2_u1_u4_n176 ) , .ZN( u2_u1_u4_n99 ) );
  AND2_X1 u2_u1_u4_U79 (.A1( u2_u1_X_26 ) , .ZN( u2_u1_u4_n101 ) , .A2( u2_u1_u4_n177 ) );
  AOI21_X1 u2_u1_u4_U8 (.ZN( u2_u1_u4_n109 ) , .A( u2_u1_u4_n153 ) , .B1( u2_u1_u4_n159 ) , .B2( u2_u1_u4_n184 ) );
  AND2_X1 u2_u1_u4_U80 (.A1( u2_u1_X_27 ) , .A2( u2_u1_X_30 ) , .ZN( u2_u1_u4_n103 ) );
  INV_X1 u2_u1_u4_U81 (.A( u2_u1_X_28 ) , .ZN( u2_u1_u4_n169 ) );
  INV_X1 u2_u1_u4_U82 (.A( u2_u1_X_29 ) , .ZN( u2_u1_u4_n168 ) );
  INV_X1 u2_u1_u4_U83 (.A( u2_u1_X_25 ) , .ZN( u2_u1_u4_n177 ) );
  INV_X1 u2_u1_u4_U84 (.A( u2_u1_X_27 ) , .ZN( u2_u1_u4_n176 ) );
  NAND4_X1 u2_u1_u4_U85 (.ZN( u2_out1_25 ) , .A4( u2_u1_u4_n139 ) , .A3( u2_u1_u4_n140 ) , .A2( u2_u1_u4_n141 ) , .A1( u2_u1_u4_n142 ) );
  OAI21_X1 u2_u1_u4_U86 (.A( u2_u1_u4_n128 ) , .B2( u2_u1_u4_n129 ) , .B1( u2_u1_u4_n130 ) , .ZN( u2_u1_u4_n142 ) );
  OAI21_X1 u2_u1_u4_U87 (.B2( u2_u1_u4_n131 ) , .ZN( u2_u1_u4_n141 ) , .A( u2_u1_u4_n175 ) , .B1( u2_u1_u4_n183 ) );
  NAND4_X1 u2_u1_u4_U88 (.ZN( u2_out1_14 ) , .A4( u2_u1_u4_n124 ) , .A3( u2_u1_u4_n125 ) , .A2( u2_u1_u4_n126 ) , .A1( u2_u1_u4_n127 ) );
  AOI22_X1 u2_u1_u4_U89 (.B2( u2_u1_u4_n117 ) , .ZN( u2_u1_u4_n126 ) , .A1( u2_u1_u4_n129 ) , .B1( u2_u1_u4_n152 ) , .A2( u2_u1_u4_n175 ) );
  AOI211_X1 u2_u1_u4_U9 (.B( u2_u1_u4_n136 ) , .A( u2_u1_u4_n137 ) , .C2( u2_u1_u4_n138 ) , .ZN( u2_u1_u4_n139 ) , .C1( u2_u1_u4_n182 ) );
  AOI22_X1 u2_u1_u4_U90 (.ZN( u2_u1_u4_n125 ) , .B2( u2_u1_u4_n131 ) , .A2( u2_u1_u4_n132 ) , .B1( u2_u1_u4_n138 ) , .A1( u2_u1_u4_n178 ) );
  NAND4_X1 u2_u1_u4_U91 (.ZN( u2_out1_8 ) , .A4( u2_u1_u4_n110 ) , .A3( u2_u1_u4_n111 ) , .A2( u2_u1_u4_n112 ) , .A1( u2_u1_u4_n186 ) );
  NAND2_X1 u2_u1_u4_U92 (.ZN( u2_u1_u4_n112 ) , .A2( u2_u1_u4_n130 ) , .A1( u2_u1_u4_n150 ) );
  AOI22_X1 u2_u1_u4_U93 (.ZN( u2_u1_u4_n111 ) , .B2( u2_u1_u4_n132 ) , .A1( u2_u1_u4_n152 ) , .B1( u2_u1_u4_n178 ) , .A2( u2_u1_u4_n97 ) );
  AOI22_X1 u2_u1_u4_U94 (.B2( u2_u1_u4_n149 ) , .B1( u2_u1_u4_n150 ) , .A2( u2_u1_u4_n151 ) , .A1( u2_u1_u4_n152 ) , .ZN( u2_u1_u4_n167 ) );
  NOR4_X1 u2_u1_u4_U95 (.A4( u2_u1_u4_n162 ) , .A3( u2_u1_u4_n163 ) , .A2( u2_u1_u4_n164 ) , .A1( u2_u1_u4_n165 ) , .ZN( u2_u1_u4_n166 ) );
  NAND3_X1 u2_u1_u4_U96 (.ZN( u2_out1_3 ) , .A3( u2_u1_u4_n166 ) , .A1( u2_u1_u4_n167 ) , .A2( u2_u1_u4_n186 ) );
  NAND3_X1 u2_u1_u4_U97 (.A3( u2_u1_u4_n146 ) , .A2( u2_u1_u4_n147 ) , .A1( u2_u1_u4_n148 ) , .ZN( u2_u1_u4_n149 ) );
  NAND3_X1 u2_u1_u4_U98 (.A3( u2_u1_u4_n143 ) , .A2( u2_u1_u4_n144 ) , .A1( u2_u1_u4_n145 ) , .ZN( u2_u1_u4_n151 ) );
  NAND3_X1 u2_u1_u4_U99 (.A3( u2_u1_u4_n121 ) , .ZN( u2_u1_u4_n122 ) , .A2( u2_u1_u4_n144 ) , .A1( u2_u1_u4_n154 ) );
  OAI22_X1 u2_uk_U162 (.ZN( u2_K2_30 ) , .B1( u2_uk_n10 ) , .B2( u2_uk_n1230 ) , .A2( u2_uk_n1259 ) , .A1( u2_uk_n162 ) );
  OAI22_X1 u2_uk_U314 (.ZN( u2_K2_26 ) , .B2( u2_uk_n1259 ) , .A2( u2_uk_n1265 ) , .B1( u2_uk_n17 ) , .A1( u2_uk_n203 ) );
  INV_X1 u2_uk_U439 (.ZN( u2_K2_28 ) , .A( u2_uk_n998 ) );
  AOI22_X1 u2_uk_U440 (.B2( u2_uk_K_r0_15 ) , .A2( u2_uk_K_r0_49 ) , .A1( u2_uk_n102 ) , .B1( u2_uk_n208 ) , .ZN( u2_uk_n998 ) );
  OAI22_X1 u2_uk_U487 (.ZN( u2_K2_29 ) , .A2( u2_uk_n1237 ) , .B2( u2_uk_n1252 ) , .A1( u2_uk_n161 ) , .B1( u2_uk_n27 ) );
  OAI21_X1 u2_uk_U692 (.ZN( u2_K2_25 ) , .B1( u2_uk_n110 ) , .B2( u2_uk_n1264 ) , .A( u2_uk_n996 ) );
  INV_X1 u2_uk_U768 (.ZN( u2_K2_27 ) , .A( u2_uk_n997 ) );
endmodule

