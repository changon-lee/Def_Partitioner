module des_des_die_0 ( clk, decrypt, desIn, key1, key2, key3, desOut, u0_FP_1, u0_FP_10, 
       u0_FP_11, u0_FP_12, u0_FP_13, u0_FP_14, u0_FP_15, u0_FP_16, u0_FP_17, u0_FP_18, u0_FP_19, 
       u0_FP_2, u0_FP_20, u0_FP_21, u0_FP_22, u0_FP_23, u0_FP_24, u0_FP_25, u0_FP_26, u0_FP_27, 
       u0_FP_28, u0_FP_29, u0_FP_3, u0_FP_30, u0_FP_31, u0_FP_32, u0_FP_4, u0_FP_5, u0_FP_6, 
       u0_FP_7, u0_FP_8, u0_FP_9, u0_N0, u0_N1, u0_N10, u0_N100, u0_N101, u0_N102, 
       u0_N103, u0_N104, u0_N105, u0_N106, u0_N107, u0_N108, u0_N109, u0_N11, u0_N110, 
       u0_N111, u0_N112, u0_N113, u0_N114, u0_N115, u0_N116, u0_N117, u0_N118, u0_N119, 
       u0_N12, u0_N120, u0_N121, u0_N122, u0_N123, u0_N124, u0_N125, u0_N126, u0_N127, 
       u0_N128, u0_N129, u0_N13, u0_N130, u0_N131, u0_N132, u0_N133, u0_N134, u0_N135, 
       u0_N136, u0_N137, u0_N138, u0_N139, u0_N14, u0_N140, u0_N141, u0_N142, u0_N143, 
       u0_N144, u0_N145, u0_N146, u0_N147, u0_N148, u0_N149, u0_N15, u0_N150, u0_N151, 
       u0_N152, u0_N153, u0_N154, u0_N155, u0_N156, u0_N157, u0_N158, u0_N159, u0_N16, 
       u0_N160, u0_N161, u0_N162, u0_N163, u0_N164, u0_N165, u0_N166, u0_N167, u0_N168, 
       u0_N169, u0_N17, u0_N170, u0_N171, u0_N172, u0_N173, u0_N174, u0_N175, u0_N176, 
       u0_N177, u0_N178, u0_N179, u0_N18, u0_N180, u0_N181, u0_N182, u0_N183, u0_N184, 
       u0_N185, u0_N186, u0_N187, u0_N188, u0_N189, u0_N19, u0_N190, u0_N191, u0_N192, 
       u0_N193, u0_N194, u0_N195, u0_N196, u0_N197, u0_N198, u0_N199, u0_N2, u0_N20, 
       u0_N200, u0_N201, u0_N202, u0_N203, u0_N204, u0_N205, u0_N206, u0_N207, u0_N208, 
       u0_N209, u0_N21, u0_N210, u0_N211, u0_N212, u0_N213, u0_N214, u0_N215, u0_N216, 
       u0_N217, u0_N218, u0_N219, u0_N22, u0_N220, u0_N221, u0_N222, u0_N223, u0_N224, 
       u0_N225, u0_N226, u0_N227, u0_N228, u0_N229, u0_N23, u0_N230, u0_N231, u0_N232, 
       u0_N233, u0_N234, u0_N235, u0_N236, u0_N237, u0_N238, u0_N239, u0_N24, u0_N240, 
       u0_N241, u0_N242, u0_N243, u0_N244, u0_N245, u0_N246, u0_N247, u0_N248, u0_N249, 
       u0_N25, u0_N250, u0_N251, u0_N252, u0_N253, u0_N254, u0_N255, u0_N256, u0_N257, 
       u0_N258, u0_N259, u0_N26, u0_N260, u0_N261, u0_N262, u0_N263, u0_N264, u0_N265, 
       u0_N266, u0_N267, u0_N268, u0_N269, u0_N27, u0_N270, u0_N271, u0_N272, u0_N273, 
       u0_N274, u0_N275, u0_N276, u0_N277, u0_N278, u0_N279, u0_N28, u0_N280, u0_N281, 
       u0_N282, u0_N283, u0_N284, u0_N285, u0_N286, u0_N287, u0_N288, u0_N289, u0_N29, 
       u0_N290, u0_N291, u0_N292, u0_N293, u0_N294, u0_N295, u0_N296, u0_N297, u0_N298, 
       u0_N299, u0_N3, u0_N30, u0_N300, u0_N301, u0_N302, u0_N303, u0_N304, u0_N305, 
       u0_N306, u0_N307, u0_N308, u0_N309, u0_N31, u0_N310, u0_N311, u0_N312, u0_N313, 
       u0_N314, u0_N315, u0_N316, u0_N317, u0_N318, u0_N319, u0_N32, u0_N320, u0_N321, 
       u0_N322, u0_N323, u0_N324, u0_N325, u0_N326, u0_N327, u0_N328, u0_N329, u0_N33, 
       u0_N330, u0_N331, u0_N332, u0_N333, u0_N334, u0_N335, u0_N336, u0_N337, u0_N338, 
       u0_N339, u0_N34, u0_N340, u0_N341, u0_N342, u0_N343, u0_N344, u0_N345, u0_N346, 
       u0_N347, u0_N348, u0_N349, u0_N35, u0_N350, u0_N351, u0_N352, u0_N353, u0_N354, 
       u0_N355, u0_N356, u0_N357, u0_N358, u0_N359, u0_N36, u0_N360, u0_N361, u0_N362, 
       u0_N363, u0_N364, u0_N365, u0_N366, u0_N367, u0_N368, u0_N369, u0_N37, u0_N370, 
       u0_N371, u0_N372, u0_N373, u0_N374, u0_N375, u0_N376, u0_N377, u0_N378, u0_N379, 
       u0_N38, u0_N380, u0_N381, u0_N382, u0_N383, u0_N384, u0_N385, u0_N386, u0_N387, 
       u0_N388, u0_N389, u0_N39, u0_N390, u0_N391, u0_N392, u0_N393, u0_N394, u0_N395, 
       u0_N396, u0_N397, u0_N398, u0_N399, u0_N4, u0_N40, u0_N400, u0_N401, u0_N402, 
       u0_N403, u0_N404, u0_N405, u0_N406, u0_N407, u0_N408, u0_N409, u0_N41, u0_N410, 
       u0_N411, u0_N412, u0_N413, u0_N414, u0_N415, u0_N416, u0_N417, u0_N418, u0_N419, 
       u0_N42, u0_N420, u0_N421, u0_N422, u0_N423, u0_N424, u0_N425, u0_N426, u0_N427, 
       u0_N428, u0_N429, u0_N43, u0_N430, u0_N431, u0_N432, u0_N433, u0_N434, u0_N435, 
       u0_N436, u0_N437, u0_N438, u0_N439, u0_N44, u0_N440, u0_N441, u0_N442, u0_N443, 
       u0_N444, u0_N445, u0_N446, u0_N447, u0_N448, u0_N449, u0_N45, u0_N450, u0_N451, 
       u0_N452, u0_N453, u0_N454, u0_N455, u0_N456, u0_N457, u0_N458, u0_N459, u0_N46, 
       u0_N460, u0_N461, u0_N462, u0_N463, u0_N464, u0_N465, u0_N466, u0_N467, u0_N468, 
       u0_N469, u0_N47, u0_N470, u0_N471, u0_N472, u0_N473, u0_N474, u0_N475, u0_N476, 
       u0_N477, u0_N478, u0_N479, u0_N48, u0_N49, u0_N5, u0_N50, u0_N51, u0_N52, 
       u0_N53, u0_N54, u0_N55, u0_N56, u0_N57, u0_N58, u0_N59, u0_N6, u0_N60, 
       u0_N61, u0_N62, u0_N63, u0_N64, u0_N65, u0_N66, u0_N67, u0_N68, u0_N69, 
       u0_N7, u0_N70, u0_N71, u0_N72, u0_N73, u0_N74, u0_N75, u0_N76, u0_N77, 
       u0_N78, u0_N79, u0_N8, u0_N80, u0_N81, u0_N82, u0_N83, u0_N84, u0_N85, 
       u0_N86, u0_N87, u0_N88, u0_N89, u0_N9, u0_N90, u0_N91, u0_N92, u0_N93, 
       u0_N94, u0_N95, u0_N96, u0_N97, u0_N98, u0_N99, u0_uk_n1010, u0_uk_n1016, u0_uk_n147, 
       u0_uk_n148, u0_uk_n155, u0_uk_n161, u0_uk_n162, u0_uk_n163, u0_uk_n164, u0_uk_n182, u0_uk_n187, u0_uk_n188, 
       u0_uk_n191, u0_uk_n202, u0_uk_n203, u0_uk_n207, u0_uk_n208, u0_uk_n209, u0_uk_n213, u0_uk_n214, u0_uk_n217, 
       u0_uk_n220, u0_uk_n222, u0_uk_n223, u0_uk_n230, u0_uk_n231, u0_uk_n238, u0_uk_n240, u0_uk_n242, u0_uk_n250, 
       u0_uk_n251, u0_uk_n252, u0_uk_n674, u0_uk_n675, u0_uk_n680, u0_uk_n684, u0_uk_n687, u0_uk_n690, u0_uk_n691, 
       u0_uk_n696, u0_uk_n697, u0_uk_n698, u0_uk_n705, u0_uk_n707, u0_uk_n711, u0_uk_n715, u0_uk_n756, u0_uk_n762, 
       u0_uk_n773, u0_uk_n777, u0_uk_n778, u0_uk_n790, u0_uk_n798, u0_uk_n804, u0_uk_n823, u0_uk_n841, u0_uk_n848, 
       u0_uk_n856, u0_uk_n863, u0_uk_n867, u0_uk_n871, u0_uk_n880, u0_uk_n888, u0_uk_n889, u0_uk_n890, u0_uk_n894, 
       u0_uk_n906, u0_uk_n926, u0_uk_n936, u0_uk_n942, u0_uk_n945, u0_uk_n961, u0_uk_n969, u0_uk_n989, u0_uk_n998, 
       u1_FP_1, u1_FP_10, u1_FP_11, u1_FP_12, u1_FP_13, u1_FP_14, u1_FP_15, u1_FP_16, u1_FP_17, 
       u1_FP_18, u1_FP_19, u1_FP_2, u1_FP_20, u1_FP_21, u1_FP_22, u1_FP_23, u1_FP_24, u1_FP_25, 
       u1_FP_26, u1_FP_27, u1_FP_28, u1_FP_29, u1_FP_3, u1_FP_30, u1_FP_31, u1_FP_32, u1_FP_4, 
       u1_FP_5, u1_FP_6, u1_FP_7, u1_FP_8, u1_FP_9, u1_N0, u1_N1, u1_N10, u1_N100, 
       u1_N101, u1_N102, u1_N103, u1_N104, u1_N105, u1_N106, u1_N107, u1_N108, u1_N109, 
       u1_N11, u1_N110, u1_N111, u1_N112, u1_N113, u1_N114, u1_N115, u1_N116, u1_N117, 
       u1_N118, u1_N119, u1_N12, u1_N120, u1_N121, u1_N122, u1_N123, u1_N124, u1_N125, 
       u1_N126, u1_N127, u1_N128, u1_N129, u1_N13, u1_N130, u1_N131, u1_N132, u1_N133, 
       u1_N134, u1_N135, u1_N136, u1_N137, u1_N138, u1_N139, u1_N14, u1_N140, u1_N141, 
       u1_N142, u1_N143, u1_N144, u1_N145, u1_N146, u1_N147, u1_N148, u1_N149, u1_N15, 
       u1_N150, u1_N151, u1_N152, u1_N153, u1_N154, u1_N155, u1_N156, u1_N157, u1_N158, 
       u1_N159, u1_N16, u1_N160, u1_N161, u1_N162, u1_N163, u1_N164, u1_N165, u1_N166, 
       u1_N167, u1_N168, u1_N169, u1_N17, u1_N170, u1_N171, u1_N172, u1_N173, u1_N174, 
       u1_N175, u1_N176, u1_N177, u1_N178, u1_N179, u1_N18, u1_N180, u1_N181, u1_N182, 
       u1_N183, u1_N184, u1_N185, u1_N186, u1_N187, u1_N188, u1_N189, u1_N19, u1_N190, 
       u1_N191, u1_N192, u1_N193, u1_N194, u1_N195, u1_N196, u1_N197, u1_N198, u1_N199, 
       u1_N2, u1_N20, u1_N200, u1_N201, u1_N202, u1_N203, u1_N204, u1_N205, u1_N206, 
       u1_N207, u1_N208, u1_N209, u1_N21, u1_N210, u1_N211, u1_N212, u1_N213, u1_N214, 
       u1_N215, u1_N216, u1_N217, u1_N218, u1_N219, u1_N22, u1_N220, u1_N221, u1_N222, 
       u1_N223, u1_N224, u1_N225, u1_N226, u1_N227, u1_N228, u1_N229, u1_N23, u1_N230, 
       u1_N231, u1_N232, u1_N233, u1_N234, u1_N235, u1_N236, u1_N237, u1_N238, u1_N239, 
       u1_N24, u1_N240, u1_N241, u1_N242, u1_N243, u1_N244, u1_N245, u1_N246, u1_N247, 
       u1_N248, u1_N249, u1_N25, u1_N250, u1_N251, u1_N252, u1_N253, u1_N254, u1_N255, 
       u1_N256, u1_N257, u1_N258, u1_N259, u1_N26, u1_N260, u1_N261, u1_N262, u1_N263, 
       u1_N264, u1_N265, u1_N266, u1_N267, u1_N268, u1_N269, u1_N27, u1_N270, u1_N271, 
       u1_N272, u1_N273, u1_N274, u1_N275, u1_N276, u1_N277, u1_N278, u1_N279, u1_N28, 
       u1_N280, u1_N281, u1_N282, u1_N283, u1_N284, u1_N285, u1_N286, u1_N287, u1_N288, 
       u1_N289, u1_N29, u1_N290, u1_N291, u1_N292, u1_N293, u1_N294, u1_N295, u1_N296, 
       u1_N297, u1_N298, u1_N299, u1_N3, u1_N30, u1_N300, u1_N301, u1_N302, u1_N303, 
       u1_N304, u1_N305, u1_N306, u1_N307, u1_N308, u1_N309, u1_N31, u1_N310, u1_N311, 
       u1_N312, u1_N313, u1_N314, u1_N315, u1_N316, u1_N317, u1_N318, u1_N319, u1_N32, 
       u1_N320, u1_N321, u1_N322, u1_N323, u1_N324, u1_N325, u1_N326, u1_N327, u1_N328, 
       u1_N329, u1_N33, u1_N330, u1_N331, u1_N332, u1_N333, u1_N334, u1_N335, u1_N336, 
       u1_N337, u1_N338, u1_N339, u1_N34, u1_N340, u1_N341, u1_N342, u1_N343, u1_N344, 
       u1_N345, u1_N346, u1_N347, u1_N348, u1_N349, u1_N35, u1_N350, u1_N351, u1_N352, 
       u1_N353, u1_N354, u1_N355, u1_N356, u1_N357, u1_N358, u1_N359, u1_N36, u1_N360, 
       u1_N361, u1_N362, u1_N363, u1_N364, u1_N365, u1_N366, u1_N367, u1_N368, u1_N369, 
       u1_N37, u1_N370, u1_N371, u1_N372, u1_N373, u1_N374, u1_N375, u1_N376, u1_N377, 
       u1_N378, u1_N379, u1_N38, u1_N380, u1_N381, u1_N382, u1_N383, u1_N384, u1_N385, 
       u1_N386, u1_N387, u1_N388, u1_N389, u1_N39, u1_N390, u1_N391, u1_N392, u1_N393, 
       u1_N394, u1_N395, u1_N396, u1_N397, u1_N398, u1_N399, u1_N4, u1_N40, u1_N400, 
       u1_N401, u1_N402, u1_N403, u1_N404, u1_N405, u1_N406, u1_N407, u1_N408, u1_N409, 
       u1_N41, u1_N410, u1_N411, u1_N412, u1_N413, u1_N414, u1_N415, u1_N416, u1_N417, 
       u1_N418, u1_N419, u1_N42, u1_N420, u1_N421, u1_N422, u1_N423, u1_N424, u1_N425, 
       u1_N426, u1_N427, u1_N428, u1_N429, u1_N43, u1_N430, u1_N431, u1_N432, u1_N433, 
       u1_N434, u1_N435, u1_N436, u1_N437, u1_N438, u1_N439, u1_N44, u1_N440, u1_N441, 
       u1_N442, u1_N443, u1_N444, u1_N445, u1_N446, u1_N447, u1_N448, u1_N449, u1_N45, 
       u1_N450, u1_N451, u1_N452, u1_N453, u1_N454, u1_N455, u1_N456, u1_N457, u1_N458, 
       u1_N459, u1_N46, u1_N460, u1_N461, u1_N462, u1_N463, u1_N464, u1_N465, u1_N466, 
       u1_N467, u1_N468, u1_N469, u1_N47, u1_N470, u1_N471, u1_N472, u1_N473, u1_N474, 
       u1_N475, u1_N476, u1_N477, u1_N478, u1_N479, u1_N48, u1_N49, u1_N5, u1_N50, 
       u1_N51, u1_N52, u1_N53, u1_N54, u1_N55, u1_N56, u1_N57, u1_N58, u1_N59, 
       u1_N6, u1_N60, u1_N61, u1_N62, u1_N63, u1_N64, u1_N65, u1_N66, u1_N67, 
       u1_N68, u1_N69, u1_N7, u1_N70, u1_N71, u1_N72, u1_N73, u1_N74, u1_N75, 
       u1_N76, u1_N77, u1_N78, u1_N79, u1_N8, u1_N80, u1_N81, u1_N82, u1_N83, 
       u1_N84, u1_N85, u1_N86, u1_N87, u1_N88, u1_N89, u1_N9, u1_N90, u1_N91, 
       u1_N92, u1_N93, u1_N94, u1_N95, u1_N96, u1_N97, u1_N98, u1_N99, u2_FP_1, 
       u2_FP_10, u2_FP_11, u2_FP_12, u2_FP_13, u2_FP_14, u2_FP_15, u2_FP_16, u2_FP_17, u2_FP_18, 
       u2_FP_19, u2_FP_2, u2_FP_20, u2_FP_21, u2_FP_22, u2_FP_23, u2_FP_24, u2_FP_25, u2_FP_26, 
       u2_FP_27, u2_FP_28, u2_FP_29, u2_FP_3, u2_FP_30, u2_FP_31, u2_FP_32, u2_FP_4, u2_FP_5, 
       u2_FP_6, u2_FP_7, u2_FP_8, u2_FP_9, u2_N0, u2_N1, u2_N10, u2_N100, u2_N101, 
       u2_N102, u2_N103, u2_N104, u2_N105, u2_N106, u2_N107, u2_N108, u2_N109, u2_N11, 
       u2_N110, u2_N111, u2_N112, u2_N113, u2_N114, u2_N115, u2_N116, u2_N117, u2_N118, 
       u2_N119, u2_N12, u2_N120, u2_N121, u2_N122, u2_N123, u2_N124, u2_N125, u2_N126, 
       u2_N127, u2_N128, u2_N129, u2_N13, u2_N130, u2_N131, u2_N132, u2_N133, u2_N134, 
       u2_N135, u2_N136, u2_N137, u2_N138, u2_N139, u2_N14, u2_N140, u2_N141, u2_N142, 
       u2_N143, u2_N144, u2_N145, u2_N146, u2_N147, u2_N148, u2_N149, u2_N15, u2_N150, 
       u2_N151, u2_N152, u2_N153, u2_N154, u2_N155, u2_N156, u2_N157, u2_N158, u2_N159, 
       u2_N16, u2_N160, u2_N161, u2_N162, u2_N163, u2_N164, u2_N165, u2_N166, u2_N167, 
       u2_N168, u2_N169, u2_N17, u2_N170, u2_N171, u2_N172, u2_N173, u2_N174, u2_N175, 
       u2_N176, u2_N177, u2_N178, u2_N179, u2_N18, u2_N180, u2_N181, u2_N182, u2_N183, 
       u2_N184, u2_N185, u2_N186, u2_N187, u2_N188, u2_N189, u2_N19, u2_N190, u2_N191, 
       u2_N192, u2_N193, u2_N194, u2_N195, u2_N196, u2_N197, u2_N198, u2_N199, u2_N2, 
       u2_N20, u2_N200, u2_N201, u2_N202, u2_N203, u2_N204, u2_N205, u2_N206, u2_N207, 
       u2_N208, u2_N209, u2_N21, u2_N210, u2_N211, u2_N212, u2_N213, u2_N214, u2_N215, 
       u2_N216, u2_N217, u2_N218, u2_N219, u2_N22, u2_N220, u2_N221, u2_N222, u2_N223, 
       u2_N224, u2_N225, u2_N226, u2_N227, u2_N228, u2_N229, u2_N23, u2_N230, u2_N231, 
       u2_N232, u2_N233, u2_N234, u2_N235, u2_N236, u2_N237, u2_N238, u2_N239, u2_N24, 
       u2_N240, u2_N241, u2_N242, u2_N243, u2_N244, u2_N245, u2_N246, u2_N247, u2_N248, 
       u2_N249, u2_N25, u2_N250, u2_N251, u2_N252, u2_N253, u2_N254, u2_N255, u2_N256, 
       u2_N257, u2_N258, u2_N259, u2_N26, u2_N260, u2_N261, u2_N262, u2_N263, u2_N264, 
       u2_N265, u2_N266, u2_N267, u2_N268, u2_N269, u2_N27, u2_N270, u2_N271, u2_N272, 
       u2_N273, u2_N274, u2_N275, u2_N276, u2_N277, u2_N278, u2_N279, u2_N28, u2_N280, 
       u2_N281, u2_N282, u2_N283, u2_N284, u2_N285, u2_N286, u2_N287, u2_N288, u2_N289, 
       u2_N29, u2_N290, u2_N291, u2_N292, u2_N293, u2_N294, u2_N295, u2_N296, u2_N297, 
       u2_N298, u2_N299, u2_N3, u2_N30, u2_N300, u2_N301, u2_N302, u2_N303, u2_N304, 
       u2_N305, u2_N306, u2_N307, u2_N308, u2_N309, u2_N31, u2_N310, u2_N311, u2_N312, 
       u2_N313, u2_N314, u2_N315, u2_N316, u2_N317, u2_N318, u2_N319, u2_N32, u2_N320, 
       u2_N321, u2_N322, u2_N323, u2_N324, u2_N325, u2_N326, u2_N327, u2_N328, u2_N329, 
       u2_N33, u2_N330, u2_N331, u2_N332, u2_N333, u2_N334, u2_N335, u2_N336, u2_N337, 
       u2_N338, u2_N339, u2_N34, u2_N340, u2_N341, u2_N342, u2_N343, u2_N344, u2_N345, 
       u2_N346, u2_N347, u2_N348, u2_N349, u2_N35, u2_N350, u2_N351, u2_N352, u2_N353, 
       u2_N354, u2_N355, u2_N356, u2_N357, u2_N358, u2_N359, u2_N36, u2_N360, u2_N361, 
       u2_N362, u2_N363, u2_N364, u2_N365, u2_N366, u2_N367, u2_N368, u2_N369, u2_N37, 
       u2_N370, u2_N371, u2_N372, u2_N373, u2_N374, u2_N375, u2_N376, u2_N377, u2_N378, 
       u2_N379, u2_N38, u2_N380, u2_N381, u2_N382, u2_N383, u2_N384, u2_N385, u2_N386, 
       u2_N387, u2_N388, u2_N389, u2_N39, u2_N390, u2_N391, u2_N392, u2_N393, u2_N394, 
       u2_N395, u2_N396, u2_N397, u2_N398, u2_N399, u2_N4, u2_N40, u2_N400, u2_N401, 
       u2_N402, u2_N403, u2_N404, u2_N405, u2_N406, u2_N407, u2_N408, u2_N409, u2_N41, 
       u2_N410, u2_N411, u2_N412, u2_N413, u2_N414, u2_N415, u2_N416, u2_N417, u2_N418, 
       u2_N419, u2_N42, u2_N420, u2_N421, u2_N422, u2_N423, u2_N424, u2_N425, u2_N426, 
       u2_N427, u2_N428, u2_N429, u2_N43, u2_N430, u2_N431, u2_N432, u2_N433, u2_N434, 
       u2_N435, u2_N436, u2_N437, u2_N438, u2_N439, u2_N44, u2_N440, u2_N441, u2_N442, 
       u2_N443, u2_N444, u2_N445, u2_N446, u2_N447, u2_N448, u2_N449, u2_N45, u2_N450, 
       u2_N451, u2_N452, u2_N453, u2_N454, u2_N455, u2_N456, u2_N457, u2_N458, u2_N459, 
       u2_N46, u2_N460, u2_N461, u2_N462, u2_N463, u2_N464, u2_N465, u2_N466, u2_N467, 
       u2_N468, u2_N469, u2_N47, u2_N470, u2_N471, u2_N472, u2_N473, u2_N474, u2_N475, 
       u2_N476, u2_N477, u2_N478, u2_N479, u2_N48, u2_N49, u2_N5, u2_N50, u2_N51, 
       u2_N52, u2_N53, u2_N54, u2_N55, u2_N56, u2_N57, u2_N58, u2_N59, u2_N6, 
       u2_N60, u2_N61, u2_N62, u2_N63, u2_N64, u2_N65, u2_N66, u2_N67, u2_N68, 
       u2_N69, u2_N7, u2_N70, u2_N71, u2_N72, u2_N73, u2_N74, u2_N75, u2_N76, 
       u2_N77, u2_N78, u2_N79, u2_N8, u2_N80, u2_N81, u2_N82, u2_N83, u2_N84, 
       u2_N85, u2_N86, u2_N87, u2_N88, u2_N89, u2_N9, u2_N90, u2_N91, u2_N92, 
       u2_N93, u2_N94, u2_N95, u2_N96, u2_N97, u2_N98, u2_N99, u2_uk_n1012, u2_uk_n1034, 
       u2_uk_n1039, u2_uk_n1056, u2_uk_n1087, u2_uk_n1090, u2_uk_n1102, u2_uk_n1142, u2_uk_n1143, u2_uk_n1144, u2_uk_n1145, 
       u2_uk_n1146, u2_uk_n1148, u2_uk_n1149, u2_uk_n1150, u2_uk_n1152, u2_uk_n1155, u2_uk_n1161, u2_uk_n1162, u2_uk_n1167, 
       u2_uk_n1168, u2_uk_n1171, u2_uk_n1178, u2_uk_n1179, u2_uk_n1183, u2_uk_n1185, u2_uk_n129, u2_uk_n141, u2_uk_n142, 
       u2_uk_n145, u2_uk_n146, u2_uk_n147, u2_uk_n148, u2_uk_n155, u2_uk_n161, u2_uk_n162, u2_uk_n163, u2_uk_n164, 
       u2_uk_n182, u2_uk_n187, u2_uk_n188, u2_uk_n191, u2_uk_n202, u2_uk_n203, u2_uk_n207, u2_uk_n208, u2_uk_n209, 
       u2_uk_n213, u2_uk_n214, u2_uk_n217, u2_uk_n220, u2_uk_n222, u2_uk_n223, u2_uk_n230, u2_uk_n231, u2_uk_n298, 
       u2_uk_n346, u2_uk_n366, u2_uk_n395, u2_uk_n605, u2_uk_n656, u2_uk_n672, u2_uk_n983, u2_uk_n988, n116, u0_FP_33, u0_FP_34, u0_FP_35, u0_FP_36, u0_FP_37, u0_FP_38, u0_FP_39, u0_FP_40, 
        u0_FP_41, u0_FP_42, u0_FP_43, u0_FP_44, u0_FP_45, u0_FP_46, u0_FP_47, u0_FP_48, u0_FP_49, 
        u0_FP_50, u0_FP_51, u0_FP_52, u0_FP_53, u0_FP_54, u0_FP_55, u0_FP_56, u0_FP_57, u0_FP_58, 
        u0_FP_59, u0_FP_60, u0_FP_61, u0_FP_62, u0_FP_63, u0_FP_64, u0_K10_10, u0_K10_13, u0_K10_14, 
        u0_K10_18, u0_K10_19, u0_K10_20, u0_K10_25, u0_K10_27, u0_K10_32, u0_K10_34, u0_K10_36, u0_K10_41, 
        u0_K11_21, u0_K11_37, u0_K11_48, u0_K12_19, u0_K12_22, u0_K12_34, u0_K12_35, u0_K12_36, u0_K12_39, 
        u0_K12_40, u0_K12_48, u0_K12_7, u0_K12_9, u0_K13_30, u0_K13_36, u0_K13_39, u0_K13_40, u0_K13_42, 
        u0_K13_45, u0_K13_46, u0_K13_48, u0_K14_10, u0_K14_12, u0_K14_13, u0_K14_14, u0_K14_15, u0_K14_18, 
        u0_K14_21, u0_K14_24, u0_K14_27, u0_K14_4, u0_K14_42, u0_K14_46, u0_K14_9, u0_K15_18, u0_K15_47, 
        u0_K16_18, u0_K16_19, u0_K16_22, u0_K16_24, u0_K16_26, u0_K16_38, u0_K16_4, u0_K16_8, u0_K1_13, 
        u0_K1_14, u0_K1_15, u0_K1_16, u0_K1_17, u0_K1_23, u0_K1_30, u0_K1_31, u0_K1_45, u0_K1_46, 
        u0_K2_11, u0_K2_12, u0_K2_25, u0_K2_30, u0_K2_34, u0_K2_35, u0_K2_4, u0_K2_44, u0_K2_45, 
        u0_K2_46, u0_K2_47, u0_K2_48, u0_K2_5, u0_K2_6, u0_K2_8, u0_K3_10, u0_K3_12, u0_K3_14, 
        u0_K3_15, u0_K3_17, u0_K3_18, u0_K3_19, u0_K3_23, u0_K3_34, u0_K3_5, u0_K4_24, u0_K4_27, 
        u0_K4_28, u0_K4_35, u0_K4_43, u0_K4_48, u0_K4_6, u0_K5_1, u0_K5_13, u0_K5_14, u0_K5_15, 
        u0_K5_16, u0_K5_18, u0_K5_19, u0_K5_23, u0_K5_24, u0_K5_26, u0_K5_28, u0_K5_3, u0_K5_31, 
        u0_K5_32, u0_K5_34, u0_K5_38, u0_K5_4, u0_K5_41, u0_K5_44, u0_K5_47, u0_K5_48, u0_K5_9, 
        u0_K6_11, u0_K6_13, u0_K6_16, u0_K6_19, u0_K6_20, u0_K6_22, u0_K6_23, u0_K6_24, u0_K6_27, 
        u0_K6_41, u0_K7_2, u0_K7_22, u0_K7_23, u0_K8_1, u0_K8_11, u0_K8_19, u0_K8_28, u0_K8_33, 
        u0_K8_36, u0_K8_45, u0_K9_14, u0_K9_15, u0_K9_32, u0_K9_39, u0_K9_4, u0_K9_40, u0_K9_45, 
        u0_K9_6, u0_L0_1, u0_L0_10, u0_L0_11, u0_L0_12, u0_L0_13, u0_L0_14, u0_L0_15, u0_L0_16, 
        u0_L0_17, u0_L0_18, u0_L0_19, u0_L0_2, u0_L0_20, u0_L0_21, u0_L0_22, u0_L0_23, u0_L0_24, 
        u0_L0_25, u0_L0_26, u0_L0_27, u0_L0_28, u0_L0_29, u0_L0_3, u0_L0_30, u0_L0_31, u0_L0_32, 
        u0_L0_4, u0_L0_5, u0_L0_6, u0_L0_7, u0_L0_8, u0_L0_9, u0_L10_1, u0_L10_10, u0_L10_11, 
        u0_L10_12, u0_L10_13, u0_L10_14, u0_L10_15, u0_L10_16, u0_L10_17, u0_L10_18, u0_L10_19, u0_L10_2, 
        u0_L10_20, u0_L10_21, u0_L10_22, u0_L10_23, u0_L10_24, u0_L10_25, u0_L10_26, u0_L10_27, u0_L10_28, 
        u0_L10_29, u0_L10_3, u0_L10_30, u0_L10_31, u0_L10_32, u0_L10_4, u0_L10_5, u0_L10_6, u0_L10_7, 
        u0_L10_8, u0_L10_9, u0_L11_1, u0_L11_10, u0_L11_11, u0_L11_12, u0_L11_13, u0_L11_14, u0_L11_15, 
        u0_L11_16, u0_L11_17, u0_L11_18, u0_L11_19, u0_L11_2, u0_L11_20, u0_L11_21, u0_L11_22, u0_L11_23, 
        u0_L11_24, u0_L11_25, u0_L11_26, u0_L11_27, u0_L11_28, u0_L11_29, u0_L11_3, u0_L11_30, u0_L11_31, 
        u0_L11_32, u0_L11_4, u0_L11_5, u0_L11_6, u0_L11_7, u0_L11_8, u0_L11_9, u0_L12_1, u0_L12_10, 
        u0_L12_11, u0_L12_12, u0_L12_13, u0_L12_14, u0_L12_15, u0_L12_16, u0_L12_17, u0_L12_18, u0_L12_19, 
        u0_L12_2, u0_L12_20, u0_L12_21, u0_L12_22, u0_L12_23, u0_L12_24, u0_L12_25, u0_L12_26, u0_L12_27, 
        u0_L12_28, u0_L12_29, u0_L12_3, u0_L12_30, u0_L12_31, u0_L12_32, u0_L12_4, u0_L12_5, u0_L12_6, 
        u0_L12_7, u0_L12_8, u0_L12_9, u0_L13_1, u0_L13_10, u0_L13_11, u0_L13_12, u0_L13_13, u0_L13_14, 
        u0_L13_15, u0_L13_16, u0_L13_17, u0_L13_18, u0_L13_19, u0_L13_2, u0_L13_20, u0_L13_21, u0_L13_22, 
        u0_L13_23, u0_L13_24, u0_L13_25, u0_L13_26, u0_L13_27, u0_L13_28, u0_L13_29, u0_L13_3, u0_L13_30, 
        u0_L13_31, u0_L13_32, u0_L13_4, u0_L13_5, u0_L13_6, u0_L13_7, u0_L13_8, u0_L13_9, u0_L14_1, 
        u0_L14_10, u0_L14_11, u0_L14_12, u0_L14_13, u0_L14_14, u0_L14_15, u0_L14_16, u0_L14_17, u0_L14_18, 
        u0_L14_19, u0_L14_2, u0_L14_20, u0_L14_21, u0_L14_22, u0_L14_23, u0_L14_24, u0_L14_25, u0_L14_26, 
        u0_L14_27, u0_L14_28, u0_L14_29, u0_L14_3, u0_L14_30, u0_L14_31, u0_L14_32, u0_L14_4, u0_L14_5, 
        u0_L14_6, u0_L14_7, u0_L14_8, u0_L14_9, u0_L1_1, u0_L1_10, u0_L1_11, u0_L1_12, u0_L1_13, 
        u0_L1_14, u0_L1_15, u0_L1_16, u0_L1_17, u0_L1_18, u0_L1_19, u0_L1_2, u0_L1_20, u0_L1_21, 
        u0_L1_22, u0_L1_23, u0_L1_24, u0_L1_25, u0_L1_26, u0_L1_27, u0_L1_28, u0_L1_29, u0_L1_3, 
        u0_L1_30, u0_L1_31, u0_L1_32, u0_L1_4, u0_L1_5, u0_L1_6, u0_L1_7, u0_L1_8, u0_L1_9, 
        u0_L2_1, u0_L2_10, u0_L2_11, u0_L2_12, u0_L2_13, u0_L2_14, u0_L2_15, u0_L2_16, u0_L2_17, 
        u0_L2_18, u0_L2_19, u0_L2_2, u0_L2_20, u0_L2_21, u0_L2_22, u0_L2_23, u0_L2_24, u0_L2_25, 
        u0_L2_26, u0_L2_27, u0_L2_28, u0_L2_29, u0_L2_3, u0_L2_30, u0_L2_31, u0_L2_32, u0_L2_4, 
        u0_L2_5, u0_L2_6, u0_L2_7, u0_L2_8, u0_L2_9, u0_L3_1, u0_L3_10, u0_L3_11, u0_L3_12, 
        u0_L3_13, u0_L3_14, u0_L3_15, u0_L3_16, u0_L3_17, u0_L3_18, u0_L3_19, u0_L3_2, u0_L3_20, 
        u0_L3_21, u0_L3_22, u0_L3_23, u0_L3_24, u0_L3_25, u0_L3_26, u0_L3_27, u0_L3_28, u0_L3_29, 
        u0_L3_3, u0_L3_30, u0_L3_31, u0_L3_32, u0_L3_4, u0_L3_5, u0_L3_6, u0_L3_7, u0_L3_8, 
        u0_L3_9, u0_L4_1, u0_L4_10, u0_L4_11, u0_L4_12, u0_L4_13, u0_L4_14, u0_L4_15, u0_L4_16, 
        u0_L4_17, u0_L4_18, u0_L4_19, u0_L4_2, u0_L4_20, u0_L4_21, u0_L4_22, u0_L4_23, u0_L4_24, 
        u0_L4_25, u0_L4_26, u0_L4_27, u0_L4_28, u0_L4_29, u0_L4_3, u0_L4_30, u0_L4_31, u0_L4_32, 
        u0_L4_4, u0_L4_5, u0_L4_6, u0_L4_7, u0_L4_8, u0_L4_9, u0_L5_1, u0_L5_10, u0_L5_11, 
        u0_L5_12, u0_L5_13, u0_L5_14, u0_L5_15, u0_L5_16, u0_L5_17, u0_L5_18, u0_L5_19, u0_L5_2, 
        u0_L5_20, u0_L5_21, u0_L5_22, u0_L5_23, u0_L5_24, u0_L5_25, u0_L5_26, u0_L5_27, u0_L5_28, 
        u0_L5_29, u0_L5_3, u0_L5_30, u0_L5_31, u0_L5_32, u0_L5_4, u0_L5_5, u0_L5_6, u0_L5_7, 
        u0_L5_8, u0_L5_9, u0_L6_1, u0_L6_10, u0_L6_11, u0_L6_12, u0_L6_13, u0_L6_14, u0_L6_15, 
        u0_L6_16, u0_L6_17, u0_L6_18, u0_L6_19, u0_L6_2, u0_L6_20, u0_L6_21, u0_L6_22, u0_L6_23, 
        u0_L6_24, u0_L6_25, u0_L6_26, u0_L6_27, u0_L6_28, u0_L6_29, u0_L6_3, u0_L6_30, u0_L6_31, 
        u0_L6_32, u0_L6_4, u0_L6_5, u0_L6_6, u0_L6_7, u0_L6_8, u0_L6_9, u0_L7_1, u0_L7_10, 
        u0_L7_11, u0_L7_12, u0_L7_13, u0_L7_14, u0_L7_15, u0_L7_16, u0_L7_17, u0_L7_18, u0_L7_19, 
        u0_L7_2, u0_L7_20, u0_L7_21, u0_L7_22, u0_L7_23, u0_L7_24, u0_L7_25, u0_L7_26, u0_L7_27, 
        u0_L7_28, u0_L7_29, u0_L7_3, u0_L7_30, u0_L7_31, u0_L7_32, u0_L7_4, u0_L7_5, u0_L7_6, 
        u0_L7_7, u0_L7_8, u0_L7_9, u0_L8_1, u0_L8_10, u0_L8_11, u0_L8_12, u0_L8_13, u0_L8_14, 
        u0_L8_15, u0_L8_16, u0_L8_17, u0_L8_18, u0_L8_19, u0_L8_2, u0_L8_20, u0_L8_21, u0_L8_22, 
        u0_L8_23, u0_L8_24, u0_L8_25, u0_L8_26, u0_L8_27, u0_L8_28, u0_L8_29, u0_L8_3, u0_L8_30, 
        u0_L8_31, u0_L8_32, u0_L8_4, u0_L8_5, u0_L8_6, u0_L8_7, u0_L8_8, u0_L8_9, u0_L9_1, 
        u0_L9_10, u0_L9_11, u0_L9_12, u0_L9_13, u0_L9_14, u0_L9_15, u0_L9_16, u0_L9_17, u0_L9_18, 
        u0_L9_19, u0_L9_2, u0_L9_20, u0_L9_21, u0_L9_22, u0_L9_23, u0_L9_24, u0_L9_25, u0_L9_26, 
        u0_L9_27, u0_L9_28, u0_L9_29, u0_L9_3, u0_L9_30, u0_L9_31, u0_L9_32, u0_L9_4, u0_L9_5, 
        u0_L9_6, u0_L9_7, u0_L9_8, u0_L9_9, u0_R0_1, u0_R0_10, u0_R0_11, u0_R0_12, u0_R0_13, 
        u0_R0_14, u0_R0_15, u0_R0_16, u0_R0_17, u0_R0_18, u0_R0_19, u0_R0_2, u0_R0_20, u0_R0_21, 
        u0_R0_22, u0_R0_23, u0_R0_24, u0_R0_25, u0_R0_26, u0_R0_27, u0_R0_28, u0_R0_29, u0_R0_3, 
        u0_R0_30, u0_R0_31, u0_R0_32, u0_R0_4, u0_R0_5, u0_R0_6, u0_R0_7, u0_R0_8, u0_R0_9, 
        u0_R10_1, u0_R10_10, u0_R10_11, u0_R10_12, u0_R10_13, u0_R10_14, u0_R10_15, u0_R10_16, u0_R10_17, 
        u0_R10_18, u0_R10_19, u0_R10_2, u0_R10_20, u0_R10_21, u0_R10_22, u0_R10_23, u0_R10_24, u0_R10_25, 
        u0_R10_26, u0_R10_27, u0_R10_28, u0_R10_29, u0_R10_3, u0_R10_30, u0_R10_31, u0_R10_32, u0_R10_4, 
        u0_R10_5, u0_R10_6, u0_R10_7, u0_R10_8, u0_R10_9, u0_R11_1, u0_R11_10, u0_R11_11, u0_R11_12, 
        u0_R11_13, u0_R11_14, u0_R11_15, u0_R11_16, u0_R11_17, u0_R11_18, u0_R11_19, u0_R11_2, u0_R11_20, 
        u0_R11_21, u0_R11_22, u0_R11_23, u0_R11_24, u0_R11_25, u0_R11_26, u0_R11_27, u0_R11_28, u0_R11_29, 
        u0_R11_3, u0_R11_30, u0_R11_31, u0_R11_32, u0_R11_4, u0_R11_5, u0_R11_6, u0_R11_7, u0_R11_8, 
        u0_R11_9, u0_R12_1, u0_R12_10, u0_R12_11, u0_R12_12, u0_R12_13, u0_R12_14, u0_R12_15, u0_R12_16, 
        u0_R12_17, u0_R12_18, u0_R12_19, u0_R12_2, u0_R12_20, u0_R12_21, u0_R12_22, u0_R12_23, u0_R12_24, 
        u0_R12_25, u0_R12_26, u0_R12_27, u0_R12_28, u0_R12_29, u0_R12_3, u0_R12_30, u0_R12_31, u0_R12_32, 
        u0_R12_4, u0_R12_5, u0_R12_6, u0_R12_7, u0_R12_8, u0_R12_9, u0_R13_1, u0_R13_10, u0_R13_11, 
        u0_R13_12, u0_R13_13, u0_R13_14, u0_R13_15, u0_R13_16, u0_R13_17, u0_R13_18, u0_R13_19, u0_R13_2, 
        u0_R13_20, u0_R13_21, u0_R13_22, u0_R13_23, u0_R13_24, u0_R13_25, u0_R13_26, u0_R13_27, u0_R13_28, 
        u0_R13_29, u0_R13_3, u0_R13_30, u0_R13_31, u0_R13_32, u0_R13_4, u0_R13_5, u0_R13_6, u0_R13_7, 
        u0_R13_8, u0_R13_9, u0_R1_1, u0_R1_10, u0_R1_11, u0_R1_12, u0_R1_13, u0_R1_14, u0_R1_15, 
        u0_R1_16, u0_R1_17, u0_R1_18, u0_R1_19, u0_R1_2, u0_R1_20, u0_R1_21, u0_R1_22, u0_R1_23, 
        u0_R1_24, u0_R1_25, u0_R1_26, u0_R1_27, u0_R1_28, u0_R1_29, u0_R1_3, u0_R1_30, u0_R1_31, 
        u0_R1_32, u0_R1_4, u0_R1_5, u0_R1_6, u0_R1_7, u0_R1_8, u0_R1_9, u0_R2_1, u0_R2_10, 
        u0_R2_11, u0_R2_12, u0_R2_13, u0_R2_14, u0_R2_15, u0_R2_16, u0_R2_17, u0_R2_18, u0_R2_19, 
        u0_R2_2, u0_R2_20, u0_R2_21, u0_R2_22, u0_R2_23, u0_R2_24, u0_R2_25, u0_R2_26, u0_R2_27, 
        u0_R2_28, u0_R2_29, u0_R2_3, u0_R2_30, u0_R2_31, u0_R2_32, u0_R2_4, u0_R2_5, u0_R2_6, 
        u0_R2_7, u0_R2_8, u0_R2_9, u0_R3_1, u0_R3_10, u0_R3_11, u0_R3_12, u0_R3_13, u0_R3_14, 
        u0_R3_15, u0_R3_16, u0_R3_17, u0_R3_18, u0_R3_19, u0_R3_2, u0_R3_20, u0_R3_21, u0_R3_22, 
        u0_R3_23, u0_R3_24, u0_R3_25, u0_R3_26, u0_R3_27, u0_R3_28, u0_R3_29, u0_R3_3, u0_R3_30, 
        u0_R3_31, u0_R3_32, u0_R3_4, u0_R3_5, u0_R3_6, u0_R3_7, u0_R3_8, u0_R3_9, u0_R4_1, 
        u0_R4_10, u0_R4_11, u0_R4_12, u0_R4_13, u0_R4_14, u0_R4_15, u0_R4_16, u0_R4_17, u0_R4_18, 
        u0_R4_19, u0_R4_2, u0_R4_20, u0_R4_21, u0_R4_22, u0_R4_23, u0_R4_24, u0_R4_25, u0_R4_26, 
        u0_R4_27, u0_R4_28, u0_R4_29, u0_R4_3, u0_R4_30, u0_R4_31, u0_R4_32, u0_R4_4, u0_R4_5, 
        u0_R4_6, u0_R4_7, u0_R4_8, u0_R4_9, u0_R5_1, u0_R5_10, u0_R5_11, u0_R5_12, u0_R5_13, 
        u0_R5_14, u0_R5_15, u0_R5_16, u0_R5_17, u0_R5_18, u0_R5_19, u0_R5_2, u0_R5_20, u0_R5_21, 
        u0_R5_22, u0_R5_23, u0_R5_24, u0_R5_25, u0_R5_26, u0_R5_27, u0_R5_28, u0_R5_29, u0_R5_3, 
        u0_R5_30, u0_R5_31, u0_R5_32, u0_R5_4, u0_R5_5, u0_R5_6, u0_R5_7, u0_R5_8, u0_R5_9, 
        u0_R6_1, u0_R6_10, u0_R6_11, u0_R6_12, u0_R6_13, u0_R6_14, u0_R6_15, u0_R6_16, u0_R6_17, 
        u0_R6_18, u0_R6_19, u0_R6_2, u0_R6_20, u0_R6_21, u0_R6_22, u0_R6_23, u0_R6_24, u0_R6_25, 
        u0_R6_26, u0_R6_27, u0_R6_28, u0_R6_29, u0_R6_3, u0_R6_30, u0_R6_31, u0_R6_32, u0_R6_4, 
        u0_R6_5, u0_R6_6, u0_R6_7, u0_R6_8, u0_R6_9, u0_R7_1, u0_R7_10, u0_R7_11, u0_R7_12, 
        u0_R7_13, u0_R7_14, u0_R7_15, u0_R7_16, u0_R7_17, u0_R7_18, u0_R7_19, u0_R7_2, u0_R7_20, 
        u0_R7_21, u0_R7_22, u0_R7_23, u0_R7_24, u0_R7_25, u0_R7_26, u0_R7_27, u0_R7_28, u0_R7_29, 
        u0_R7_3, u0_R7_30, u0_R7_31, u0_R7_32, u0_R7_4, u0_R7_5, u0_R7_6, u0_R7_7, u0_R7_8, 
        u0_R7_9, u0_R8_1, u0_R8_10, u0_R8_11, u0_R8_12, u0_R8_13, u0_R8_14, u0_R8_15, u0_R8_16, 
        u0_R8_17, u0_R8_18, u0_R8_19, u0_R8_2, u0_R8_20, u0_R8_21, u0_R8_22, u0_R8_23, u0_R8_24, 
        u0_R8_25, u0_R8_26, u0_R8_27, u0_R8_28, u0_R8_29, u0_R8_3, u0_R8_30, u0_R8_31, u0_R8_32, 
        u0_R8_4, u0_R8_5, u0_R8_6, u0_R8_7, u0_R8_8, u0_R8_9, u0_R9_1, u0_R9_10, u0_R9_11, 
        u0_R9_12, u0_R9_13, u0_R9_14, u0_R9_15, u0_R9_16, u0_R9_17, u0_R9_18, u0_R9_19, u0_R9_2, 
        u0_R9_20, u0_R9_21, u0_R9_22, u0_R9_23, u0_R9_24, u0_R9_25, u0_R9_26, u0_R9_27, u0_R9_28, 
        u0_R9_29, u0_R9_3, u0_R9_30, u0_R9_31, u0_R9_32, u0_R9_4, u0_R9_5, u0_R9_6, u0_R9_7, 
        u0_R9_8, u0_R9_9, u0_desIn_r_0, u0_desIn_r_1, u0_desIn_r_10, u0_desIn_r_11, u0_desIn_r_12, u0_desIn_r_13, u0_desIn_r_14, 
        u0_desIn_r_15, u0_desIn_r_16, u0_desIn_r_17, u0_desIn_r_18, u0_desIn_r_19, u0_desIn_r_2, u0_desIn_r_20, u0_desIn_r_21, u0_desIn_r_22, 
        u0_desIn_r_23, u0_desIn_r_24, u0_desIn_r_25, u0_desIn_r_26, u0_desIn_r_27, u0_desIn_r_28, u0_desIn_r_29, u0_desIn_r_3, u0_desIn_r_30, 
        u0_desIn_r_31, u0_desIn_r_32, u0_desIn_r_33, u0_desIn_r_34, u0_desIn_r_35, u0_desIn_r_36, u0_desIn_r_37, u0_desIn_r_38, u0_desIn_r_39, 
        u0_desIn_r_4, u0_desIn_r_40, u0_desIn_r_41, u0_desIn_r_42, u0_desIn_r_43, u0_desIn_r_44, u0_desIn_r_45, u0_desIn_r_46, u0_desIn_r_47, 
        u0_desIn_r_48, u0_desIn_r_49, u0_desIn_r_5, u0_desIn_r_50, u0_desIn_r_51, u0_desIn_r_52, u0_desIn_r_53, u0_desIn_r_54, u0_desIn_r_55, 
        u0_desIn_r_56, u0_desIn_r_57, u0_desIn_r_58, u0_desIn_r_59, u0_desIn_r_6, u0_desIn_r_60, u0_desIn_r_61, u0_desIn_r_62, u0_desIn_r_63, 
        u0_desIn_r_7, u0_desIn_r_8, u0_desIn_r_9, u0_key_r_0, u0_key_r_1, u0_key_r_10, u0_key_r_11, u0_key_r_12, u0_key_r_13, 
        u0_key_r_14, u0_key_r_16, u0_key_r_17, u0_key_r_18, u0_key_r_19, u0_key_r_2, u0_key_r_20, u0_key_r_21, u0_key_r_22, 
        u0_key_r_23, u0_key_r_24, u0_key_r_25, u0_key_r_26, u0_key_r_27, u0_key_r_28, u0_key_r_29, u0_key_r_3, u0_key_r_30, 
        u0_key_r_31, u0_key_r_32, u0_key_r_33, u0_key_r_34, u0_key_r_35, u0_key_r_36, u0_key_r_37, u0_key_r_38, u0_key_r_39, 
        u0_key_r_4, u0_key_r_40, u0_key_r_41, u0_key_r_42, u0_key_r_43, u0_key_r_44, u0_key_r_45, u0_key_r_46, u0_key_r_47, 
        u0_key_r_48, u0_key_r_49, u0_key_r_5, u0_key_r_50, u0_key_r_51, u0_key_r_52, u0_key_r_53, u0_key_r_54, u0_key_r_55, 
        u0_key_r_6, u0_key_r_7, u0_key_r_8, u0_key_r_9, u0_uk_K_r0_11, u0_uk_K_r0_15, u0_uk_K_r0_19, u0_uk_K_r0_2, u0_uk_K_r0_22, 
        u0_uk_K_r0_25, u0_uk_K_r0_28, u0_uk_K_r0_31, u0_uk_K_r0_32, u0_uk_K_r0_34, u0_uk_K_r0_36, u0_uk_K_r0_47, u0_uk_K_r0_49, u0_uk_K_r0_52, 
        u0_uk_K_r0_55, u0_uk_K_r0_7, u0_uk_K_r10_10, u0_uk_K_r10_14, u0_uk_K_r10_16, u0_uk_K_r10_18, u0_uk_K_r10_19, u0_uk_K_r10_23, u0_uk_K_r10_25, 
        u0_uk_K_r10_27, u0_uk_K_r10_28, u0_uk_K_r10_32, u0_uk_K_r10_34, u0_uk_K_r10_37, u0_uk_K_r10_39, u0_uk_K_r10_41, u0_uk_K_r10_42, u0_uk_K_r10_43, 
        u0_uk_K_r10_44, u0_uk_K_r10_47, u0_uk_K_r10_48, u0_uk_K_r10_9, u0_uk_K_r11_10, u0_uk_K_r11_11, u0_uk_K_r11_17, u0_uk_K_r11_19, u0_uk_K_r11_20, 
        u0_uk_K_r11_21, u0_uk_K_r11_24, u0_uk_K_r11_25, u0_uk_K_r11_26, u0_uk_K_r11_27, u0_uk_K_r11_28, u0_uk_K_r11_29, u0_uk_K_r11_33, u0_uk_K_r11_34, 
        u0_uk_K_r11_39, u0_uk_K_r11_4, u0_uk_K_r11_46, u0_uk_K_r11_47, u0_uk_K_r11_48, u0_uk_K_r11_53, u0_uk_K_r11_54, u0_uk_K_r11_6, u0_uk_K_r11_8, 
        u0_uk_K_r12_1, u0_uk_K_r12_10, u0_uk_K_r12_15, u0_uk_K_r12_16, u0_uk_K_r12_18, u0_uk_K_r12_21, u0_uk_K_r12_25, u0_uk_K_r12_30, u0_uk_K_r12_33, 
        u0_uk_K_r12_36, u0_uk_K_r12_42, u0_uk_K_r12_44, u0_uk_K_r12_47, u0_uk_K_r12_7, u0_uk_K_r13_0, u0_uk_K_r13_13, u0_uk_K_r13_17, u0_uk_K_r13_19, 
        u0_uk_K_r13_2, u0_uk_K_r13_22, u0_uk_K_r13_23, u0_uk_K_r13_25, u0_uk_K_r13_32, u0_uk_K_r13_35, u0_uk_K_r13_38, u0_uk_K_r13_4, u0_uk_K_r13_44, 
        u0_uk_K_r13_55, u0_uk_K_r14_10, u0_uk_K_r14_11, u0_uk_K_r14_12, u0_uk_K_r14_15, u0_uk_K_r14_16, u0_uk_K_r14_18, u0_uk_K_r14_2, u0_uk_K_r14_3, 
        u0_uk_K_r14_39, u0_uk_K_r14_43, u0_uk_K_r14_45, u0_uk_K_r14_46, u0_uk_K_r14_5, u0_uk_K_r14_50, u0_uk_K_r14_8, u0_uk_K_r14_9, u0_uk_K_r1_10, 
        u0_uk_K_r1_15, u0_uk_K_r1_16, u0_uk_K_r1_17, u0_uk_K_r1_18, u0_uk_K_r1_21, u0_uk_K_r1_22, u0_uk_K_r1_36, u0_uk_K_r1_41, u0_uk_K_r1_42, 
        u0_uk_K_r1_44, u0_uk_K_r1_47, u0_uk_K_r1_7, u0_uk_K_r2_13, u0_uk_K_r2_16, u0_uk_K_r2_18, u0_uk_K_r2_20, u0_uk_K_r2_25, u0_uk_K_r2_26, 
        u0_uk_K_r2_27, u0_uk_K_r2_28, u0_uk_K_r2_29, u0_uk_K_r2_31, u0_uk_K_r2_33, u0_uk_K_r2_36, u0_uk_K_r2_4, u0_uk_K_r2_41, u0_uk_K_r2_46, 
        u0_uk_K_r2_50, u0_uk_K_r2_53, u0_uk_K_r2_55, u0_uk_K_r2_7, u0_uk_K_r3_10, u0_uk_K_r3_11, u0_uk_K_r3_14, u0_uk_K_r3_15, u0_uk_K_r3_16, 
        u0_uk_K_r3_19, u0_uk_K_r3_24, u0_uk_K_r3_29, u0_uk_K_r3_35, u0_uk_K_r3_38, u0_uk_K_r3_4, u0_uk_K_r3_47, u0_uk_K_r3_52, u0_uk_K_r3_9, 
        u0_uk_K_r4_0, u0_uk_K_r4_11, u0_uk_K_r4_23, u0_uk_K_r4_3, u0_uk_K_r4_31, u0_uk_K_r4_33, u0_uk_K_r4_35, u0_uk_K_r4_38, u0_uk_K_r4_4, 
        u0_uk_K_r4_41, u0_uk_K_r4_47, u0_uk_K_r4_48, u0_uk_K_r4_49, u0_uk_K_r4_5, u0_uk_K_r4_54, u0_uk_K_r4_55, u0_uk_K_r5_0, u0_uk_K_r5_1, 
        u0_uk_K_r5_10, u0_uk_K_r5_13, u0_uk_K_r5_16, u0_uk_K_r5_17, u0_uk_K_r5_18, u0_uk_K_r5_19, u0_uk_K_r5_21, u0_uk_K_r5_23, u0_uk_K_r5_26, 
        u0_uk_K_r5_32, u0_uk_K_r5_37, u0_uk_K_r5_39, u0_uk_K_r5_4, u0_uk_K_r5_40, u0_uk_K_r5_41, u0_uk_K_r5_43, u0_uk_K_r5_48, u0_uk_K_r5_5, 
        u0_uk_K_r5_51, u0_uk_K_r5_8, u0_uk_K_r6_0, u0_uk_K_r6_10, u0_uk_K_r6_14, u0_uk_K_r6_19, u0_uk_K_r6_21, u0_uk_K_r6_22, u0_uk_K_r6_26, 
        u0_uk_K_r6_27, u0_uk_K_r6_29, u0_uk_K_r6_3, u0_uk_K_r6_31, u0_uk_K_r6_34, u0_uk_K_r6_37, u0_uk_K_r6_46, u0_uk_K_r6_51, u0_uk_K_r6_53, 
        u0_uk_K_r6_55, u0_uk_K_r6_7, u0_uk_K_r7_0, u0_uk_K_r7_1, u0_uk_K_r7_13, u0_uk_K_r7_15, u0_uk_K_r7_2, u0_uk_K_r7_20, u0_uk_K_r7_22, 
        u0_uk_K_r7_23, u0_uk_K_r7_24, u0_uk_K_r7_25, u0_uk_K_r7_26, u0_uk_K_r7_27, u0_uk_K_r7_30, u0_uk_K_r7_32, u0_uk_K_r7_39, u0_uk_K_r7_48, 
        u0_uk_K_r7_55, u0_uk_K_r7_6, u0_uk_K_r7_8, u0_uk_K_r7_9, u0_uk_K_r8_13, u0_uk_K_r8_16, u0_uk_K_r8_17, u0_uk_K_r8_2, u0_uk_K_r8_21, 
        u0_uk_K_r8_22, u0_uk_K_r8_27, u0_uk_K_r8_28, u0_uk_K_r8_32, u0_uk_K_r8_37, u0_uk_K_r8_40, u0_uk_K_r8_41, u0_uk_K_r8_43, u0_uk_K_r8_44, 
        u0_uk_K_r8_52, u0_uk_K_r8_8, u0_uk_K_r9_0, u0_uk_K_r9_1, u0_uk_K_r9_10, u0_uk_K_r9_12, u0_uk_K_r9_13, u0_uk_K_r9_15, u0_uk_K_r9_18, 
        u0_uk_K_r9_19, u0_uk_K_r9_22, u0_uk_K_r9_23, u0_uk_K_r9_25, u0_uk_K_r9_27, u0_uk_K_r9_30, u0_uk_K_r9_31, u0_uk_K_r9_33, u0_uk_K_r9_35, 
        u0_uk_K_r9_38, u0_uk_K_r9_45, u0_uk_K_r9_48, u0_uk_K_r9_49, u0_uk_K_r9_5, u0_uk_K_r9_6, u0_uk_K_r9_7, u0_uk_K_r9_9, u0_uk_n1, 
        u0_uk_n1001, u0_uk_n1002, u0_uk_n1004, u0_uk_n1009, u0_uk_n101, u0_uk_n1012, u0_uk_n1019, u0_uk_n1020, u0_uk_n1021, 
        u0_uk_n1024, u0_uk_n103, u0_uk_n104, u0_uk_n105, u0_uk_n106, u0_uk_n107, u0_uk_n108, u0_uk_n111, u0_uk_n112, 
        u0_uk_n113, u0_uk_n115, u0_uk_n116, u0_uk_n119, u0_uk_n12, u0_uk_n120, u0_uk_n121, u0_uk_n122, u0_uk_n123, 
        u0_uk_n124, u0_uk_n126, u0_uk_n127, u0_uk_n13, u0_uk_n130, u0_uk_n131, u0_uk_n132, u0_uk_n134, u0_uk_n135, 
        u0_uk_n136, u0_uk_n137, u0_uk_n139, u0_uk_n14, u0_uk_n140, u0_uk_n143, u0_uk_n144, u0_uk_n149, u0_uk_n15, 
        u0_uk_n150, u0_uk_n151, u0_uk_n152, u0_uk_n153, u0_uk_n154, u0_uk_n156, u0_uk_n157, u0_uk_n159, u0_uk_n16, 
        u0_uk_n165, u0_uk_n166, u0_uk_n167, u0_uk_n168, u0_uk_n169, u0_uk_n170, u0_uk_n171, u0_uk_n172, u0_uk_n173, 
        u0_uk_n174, u0_uk_n175, u0_uk_n176, u0_uk_n177, u0_uk_n178, u0_uk_n179, u0_uk_n18, u0_uk_n180, u0_uk_n181, 
        u0_uk_n183, u0_uk_n184, u0_uk_n185, u0_uk_n186, u0_uk_n189, u0_uk_n19, u0_uk_n190, u0_uk_n192, u0_uk_n193, 
        u0_uk_n194, u0_uk_n195, u0_uk_n196, u0_uk_n197, u0_uk_n198, u0_uk_n199, u0_uk_n20, u0_uk_n200, u0_uk_n201, 
        u0_uk_n204, u0_uk_n205, u0_uk_n206, u0_uk_n21, u0_uk_n210, u0_uk_n211, u0_uk_n212, u0_uk_n215, u0_uk_n216, 
        u0_uk_n218, u0_uk_n219, u0_uk_n22, u0_uk_n221, u0_uk_n224, u0_uk_n225, u0_uk_n226, u0_uk_n227, u0_uk_n228, 
        u0_uk_n229, u0_uk_n23, u0_uk_n232, u0_uk_n233, u0_uk_n234, u0_uk_n235, u0_uk_n237, u0_uk_n239, u0_uk_n24, 
        u0_uk_n241, u0_uk_n243, u0_uk_n244, u0_uk_n245, u0_uk_n246, u0_uk_n247, u0_uk_n248, u0_uk_n249, u0_uk_n25, 
        u0_uk_n253, u0_uk_n254, u0_uk_n255, u0_uk_n256, u0_uk_n257, u0_uk_n258, u0_uk_n259, u0_uk_n26, u0_uk_n260, 
        u0_uk_n261, u0_uk_n262, u0_uk_n263, u0_uk_n264, u0_uk_n265, u0_uk_n266, u0_uk_n267, u0_uk_n268, u0_uk_n269, 
        u0_uk_n272, u0_uk_n273, u0_uk_n274, u0_uk_n275, u0_uk_n276, u0_uk_n278, u0_uk_n28, u0_uk_n280, u0_uk_n281, 
        u0_uk_n282, u0_uk_n283, u0_uk_n285, u0_uk_n288, u0_uk_n289, u0_uk_n29, u0_uk_n290, u0_uk_n293, u0_uk_n296, 
        u0_uk_n3, u0_uk_n30, u0_uk_n300, u0_uk_n303, u0_uk_n304, u0_uk_n307, u0_uk_n309, u0_uk_n310, u0_uk_n311, 
        u0_uk_n314, u0_uk_n315, u0_uk_n316, u0_uk_n318, u0_uk_n32, u0_uk_n320, u0_uk_n321, u0_uk_n322, u0_uk_n323, 
        u0_uk_n324, u0_uk_n325, u0_uk_n326, u0_uk_n327, u0_uk_n328, u0_uk_n329, u0_uk_n33, u0_uk_n330, u0_uk_n331, 
        u0_uk_n332, u0_uk_n333, u0_uk_n336, u0_uk_n337, u0_uk_n339, u0_uk_n34, u0_uk_n340, u0_uk_n341, u0_uk_n343, 
        u0_uk_n344, u0_uk_n345, u0_uk_n347, u0_uk_n348, u0_uk_n35, u0_uk_n350, u0_uk_n351, u0_uk_n352, u0_uk_n354, 
        u0_uk_n355, u0_uk_n356, u0_uk_n357, u0_uk_n358, u0_uk_n359, u0_uk_n36, u0_uk_n361, u0_uk_n362, u0_uk_n364, 
        u0_uk_n365, u0_uk_n367, u0_uk_n368, u0_uk_n37, u0_uk_n370, u0_uk_n371, u0_uk_n372, u0_uk_n374, u0_uk_n378, 
        u0_uk_n38, u0_uk_n380, u0_uk_n381, u0_uk_n383, u0_uk_n384, u0_uk_n387, u0_uk_n388, u0_uk_n389, u0_uk_n39, 
        u0_uk_n390, u0_uk_n392, u0_uk_n393, u0_uk_n394, u0_uk_n396, u0_uk_n397, u0_uk_n398, u0_uk_n399, u0_uk_n4, 
        u0_uk_n40, u0_uk_n400, u0_uk_n401, u0_uk_n402, u0_uk_n403, u0_uk_n404, u0_uk_n405, u0_uk_n406, u0_uk_n41, 
        u0_uk_n410, u0_uk_n411, u0_uk_n412, u0_uk_n413, u0_uk_n414, u0_uk_n417, u0_uk_n418, u0_uk_n419, u0_uk_n42, 
        u0_uk_n420, u0_uk_n423, u0_uk_n424, u0_uk_n425, u0_uk_n426, u0_uk_n427, u0_uk_n428, u0_uk_n429, u0_uk_n43, 
        u0_uk_n430, u0_uk_n432, u0_uk_n433, u0_uk_n434, u0_uk_n435, u0_uk_n436, u0_uk_n438, u0_uk_n439, u0_uk_n44, 
        u0_uk_n440, u0_uk_n441, u0_uk_n442, u0_uk_n445, u0_uk_n446, u0_uk_n447, u0_uk_n448, u0_uk_n45, u0_uk_n450, 
        u0_uk_n451, u0_uk_n453, u0_uk_n455, u0_uk_n457, u0_uk_n458, u0_uk_n459, u0_uk_n46, u0_uk_n462, u0_uk_n463, 
        u0_uk_n464, u0_uk_n465, u0_uk_n466, u0_uk_n471, u0_uk_n473, u0_uk_n475, u0_uk_n476, u0_uk_n479, u0_uk_n48, 
        u0_uk_n480, u0_uk_n481, u0_uk_n482, u0_uk_n483, u0_uk_n484, u0_uk_n485, u0_uk_n486, u0_uk_n488, u0_uk_n489, 
        u0_uk_n49, u0_uk_n490, u0_uk_n491, u0_uk_n493, u0_uk_n494, u0_uk_n497, u0_uk_n498, u0_uk_n499, u0_uk_n5, 
        u0_uk_n50, u0_uk_n502, u0_uk_n505, u0_uk_n506, u0_uk_n507, u0_uk_n508, u0_uk_n51, u0_uk_n510, u0_uk_n511, 
        u0_uk_n512, u0_uk_n513, u0_uk_n514, u0_uk_n516, u0_uk_n517, u0_uk_n519, u0_uk_n52, u0_uk_n521, u0_uk_n522, 
        u0_uk_n523, u0_uk_n525, u0_uk_n527, u0_uk_n528, u0_uk_n529, u0_uk_n53, u0_uk_n530, u0_uk_n531, u0_uk_n532, 
        u0_uk_n534, u0_uk_n535, u0_uk_n536, u0_uk_n537, u0_uk_n538, u0_uk_n539, u0_uk_n54, u0_uk_n540, u0_uk_n542, 
        u0_uk_n543, u0_uk_n544, u0_uk_n545, u0_uk_n546, u0_uk_n547, u0_uk_n549, u0_uk_n55, u0_uk_n550, u0_uk_n552, 
        u0_uk_n553, u0_uk_n554, u0_uk_n555, u0_uk_n557, u0_uk_n558, u0_uk_n559, u0_uk_n56, u0_uk_n560, u0_uk_n561, 
        u0_uk_n562, u0_uk_n563, u0_uk_n564, u0_uk_n565, u0_uk_n566, u0_uk_n567, u0_uk_n568, u0_uk_n569, u0_uk_n57, 
        u0_uk_n570, u0_uk_n571, u0_uk_n573, u0_uk_n574, u0_uk_n575, u0_uk_n576, u0_uk_n577, u0_uk_n578, u0_uk_n579, 
        u0_uk_n58, u0_uk_n580, u0_uk_n581, u0_uk_n583, u0_uk_n584, u0_uk_n588, u0_uk_n589, u0_uk_n59, u0_uk_n592, 
        u0_uk_n593, u0_uk_n594, u0_uk_n596, u0_uk_n597, u0_uk_n598, u0_uk_n599, u0_uk_n6, u0_uk_n600, u0_uk_n604, 
        u0_uk_n606, u0_uk_n607, u0_uk_n609, u0_uk_n61, u0_uk_n610, u0_uk_n611, u0_uk_n612, u0_uk_n613, u0_uk_n614, 
        u0_uk_n615, u0_uk_n616, u0_uk_n619, u0_uk_n62, u0_uk_n620, u0_uk_n621, u0_uk_n622, u0_uk_n623, u0_uk_n624, 
        u0_uk_n625, u0_uk_n626, u0_uk_n627, u0_uk_n628, u0_uk_n629, u0_uk_n630, u0_uk_n631, u0_uk_n632, u0_uk_n633, 
        u0_uk_n635, u0_uk_n636, u0_uk_n637, u0_uk_n638, u0_uk_n639, u0_uk_n64, u0_uk_n640, u0_uk_n641, u0_uk_n642, 
        u0_uk_n643, u0_uk_n644, u0_uk_n645, u0_uk_n646, u0_uk_n647, u0_uk_n648, u0_uk_n649, u0_uk_n65, u0_uk_n650, 
        u0_uk_n651, u0_uk_n652, u0_uk_n653, u0_uk_n654, u0_uk_n655, u0_uk_n657, u0_uk_n658, u0_uk_n659, u0_uk_n66, 
        u0_uk_n660, u0_uk_n661, u0_uk_n663, u0_uk_n664, u0_uk_n666, u0_uk_n667, u0_uk_n668, u0_uk_n669, u0_uk_n67, 
        u0_uk_n670, u0_uk_n68, u0_uk_n69, u0_uk_n7, u0_uk_n719, u0_uk_n72, u0_uk_n720, u0_uk_n725, u0_uk_n726, 
        u0_uk_n728, u0_uk_n73, u0_uk_n731, u0_uk_n732, u0_uk_n735, u0_uk_n736, u0_uk_n739, u0_uk_n740, u0_uk_n746, 
        u0_uk_n748, u0_uk_n75, u0_uk_n755, u0_uk_n759, u0_uk_n763, u0_uk_n765, u0_uk_n766, u0_uk_n77, u0_uk_n770, 
        u0_uk_n775, u0_uk_n78, u0_uk_n780, u0_uk_n785, u0_uk_n786, u0_uk_n79, u0_uk_n793, u0_uk_n799, u0_uk_n8, 
        u0_uk_n80, u0_uk_n805, u0_uk_n81, u0_uk_n810, u0_uk_n813, u0_uk_n815, u0_uk_n82, u0_uk_n826, u0_uk_n832, 
        u0_uk_n834, u0_uk_n839, u0_uk_n84, u0_uk_n85, u0_uk_n853, u0_uk_n855, u0_uk_n86, u0_uk_n87, u0_uk_n875, 
        u0_uk_n878, u0_uk_n88, u0_uk_n89, u0_uk_n897, u0_uk_n898, u0_uk_n9, u0_uk_n90, u0_uk_n904, u0_uk_n91, 
        u0_uk_n916, u0_uk_n917, u0_uk_n918, u0_uk_n939, u0_uk_n948, u0_uk_n95, u0_uk_n950, u0_uk_n96, u0_uk_n960, 
        u0_uk_n963, u0_uk_n97, u0_uk_n98, u0_uk_n981, u0_uk_n990, u0_uk_n999, u1_FP_33, u1_FP_34, u1_FP_35, 
        u1_FP_36, u1_FP_37, u1_FP_38, u1_FP_39, u1_FP_40, u1_FP_41, u1_FP_42, u1_FP_43, u1_FP_44, 
        u1_FP_45, u1_FP_46, u1_FP_47, u1_FP_48, u1_FP_49, u1_FP_50, u1_FP_51, u1_FP_52, u1_FP_53, 
        u1_FP_54, u1_FP_55, u1_FP_56, u1_FP_57, u1_FP_58, u1_FP_59, u1_FP_60, u1_FP_61, u1_FP_62, 
        u1_FP_63, u1_FP_64, u1_L0_1, u1_L0_10, u1_L0_11, u1_L0_12, u1_L0_13, u1_L0_14, u1_L0_15, 
        u1_L0_16, u1_L0_17, u1_L0_18, u1_L0_19, u1_L0_2, u1_L0_20, u1_L0_21, u1_L0_22, u1_L0_23, 
        u1_L0_24, u1_L0_25, u1_L0_26, u1_L0_27, u1_L0_28, u1_L0_29, u1_L0_3, u1_L0_30, u1_L0_31, 
        u1_L0_32, u1_L0_4, u1_L0_5, u1_L0_6, u1_L0_7, u1_L0_8, u1_L0_9, u1_L10_1, u1_L10_10, 
        u1_L10_11, u1_L10_12, u1_L10_13, u1_L10_14, u1_L10_15, u1_L10_16, u1_L10_17, u1_L10_18, u1_L10_19, 
        u1_L10_2, u1_L10_20, u1_L10_21, u1_L10_22, u1_L10_23, u1_L10_24, u1_L10_25, u1_L10_26, u1_L10_27, 
        u1_L10_28, u1_L10_29, u1_L10_3, u1_L10_30, u1_L10_31, u1_L10_32, u1_L10_4, u1_L10_5, u1_L10_6, 
        u1_L10_7, u1_L10_8, u1_L10_9, u1_L11_1, u1_L11_10, u1_L11_11, u1_L11_12, u1_L11_13, u1_L11_14, 
        u1_L11_15, u1_L11_16, u1_L11_17, u1_L11_18, u1_L11_19, u1_L11_2, u1_L11_20, u1_L11_21, u1_L11_22, 
        u1_L11_23, u1_L11_24, u1_L11_25, u1_L11_26, u1_L11_27, u1_L11_28, u1_L11_29, u1_L11_3, u1_L11_30, 
        u1_L11_31, u1_L11_32, u1_L11_4, u1_L11_5, u1_L11_6, u1_L11_7, u1_L11_8, u1_L11_9, u1_L12_1, 
        u1_L12_10, u1_L12_11, u1_L12_12, u1_L12_13, u1_L12_14, u1_L12_15, u1_L12_16, u1_L12_17, u1_L12_18, 
        u1_L12_19, u1_L12_2, u1_L12_20, u1_L12_21, u1_L12_22, u1_L12_23, u1_L12_24, u1_L12_25, u1_L12_26, 
        u1_L12_27, u1_L12_28, u1_L12_29, u1_L12_3, u1_L12_30, u1_L12_31, u1_L12_32, u1_L12_4, u1_L12_5, 
        u1_L12_6, u1_L12_7, u1_L12_8, u1_L12_9, u1_L13_1, u1_L13_10, u1_L13_11, u1_L13_12, u1_L13_13, 
        u1_L13_14, u1_L13_15, u1_L13_16, u1_L13_17, u1_L13_18, u1_L13_19, u1_L13_2, u1_L13_20, u1_L13_21, 
        u1_L13_22, u1_L13_23, u1_L13_24, u1_L13_25, u1_L13_26, u1_L13_27, u1_L13_28, u1_L13_29, u1_L13_3, 
        u1_L13_30, u1_L13_31, u1_L13_32, u1_L13_4, u1_L13_5, u1_L13_6, u1_L13_7, u1_L13_8, u1_L13_9, 
        u1_L14_1, u1_L14_10, u1_L14_11, u1_L14_12, u1_L14_13, u1_L14_14, u1_L14_15, u1_L14_16, u1_L14_17, 
        u1_L14_18, u1_L14_19, u1_L14_2, u1_L14_20, u1_L14_21, u1_L14_22, u1_L14_23, u1_L14_24, u1_L14_25, 
        u1_L14_26, u1_L14_27, u1_L14_28, u1_L14_29, u1_L14_3, u1_L14_30, u1_L14_31, u1_L14_32, u1_L14_4, 
        u1_L14_5, u1_L14_6, u1_L14_7, u1_L14_8, u1_L14_9, u1_L1_1, u1_L1_10, u1_L1_11, u1_L1_12, 
        u1_L1_13, u1_L1_14, u1_L1_15, u1_L1_16, u1_L1_17, u1_L1_18, u1_L1_19, u1_L1_2, u1_L1_20, 
        u1_L1_21, u1_L1_22, u1_L1_23, u1_L1_24, u1_L1_25, u1_L1_26, u1_L1_27, u1_L1_28, u1_L1_29, 
        u1_L1_3, u1_L1_30, u1_L1_31, u1_L1_32, u1_L1_4, u1_L1_5, u1_L1_6, u1_L1_7, u1_L1_8, 
        u1_L1_9, u1_L2_1, u1_L2_10, u1_L2_11, u1_L2_12, u1_L2_13, u1_L2_14, u1_L2_15, u1_L2_16, 
        u1_L2_17, u1_L2_18, u1_L2_19, u1_L2_2, u1_L2_20, u1_L2_21, u1_L2_22, u1_L2_23, u1_L2_24, 
        u1_L2_25, u1_L2_26, u1_L2_27, u1_L2_28, u1_L2_29, u1_L2_3, u1_L2_30, u1_L2_31, u1_L2_32, 
        u1_L2_4, u1_L2_5, u1_L2_6, u1_L2_7, u1_L2_8, u1_L2_9, u1_L3_1, u1_L3_10, u1_L3_11, 
        u1_L3_12, u1_L3_13, u1_L3_14, u1_L3_15, u1_L3_16, u1_L3_17, u1_L3_18, u1_L3_19, u1_L3_2, 
        u1_L3_20, u1_L3_21, u1_L3_22, u1_L3_23, u1_L3_24, u1_L3_25, u1_L3_26, u1_L3_27, u1_L3_28, 
        u1_L3_29, u1_L3_3, u1_L3_30, u1_L3_31, u1_L3_32, u1_L3_4, u1_L3_5, u1_L3_6, u1_L3_7, 
        u1_L3_8, u1_L3_9, u1_L4_1, u1_L4_10, u1_L4_11, u1_L4_12, u1_L4_13, u1_L4_14, u1_L4_15, 
        u1_L4_16, u1_L4_17, u1_L4_18, u1_L4_19, u1_L4_2, u1_L4_20, u1_L4_21, u1_L4_22, u1_L4_23, 
        u1_L4_24, u1_L4_25, u1_L4_26, u1_L4_27, u1_L4_28, u1_L4_29, u1_L4_3, u1_L4_30, u1_L4_31, 
        u1_L4_32, u1_L4_4, u1_L4_5, u1_L4_6, u1_L4_7, u1_L4_8, u1_L4_9, u1_L5_1, u1_L5_10, 
        u1_L5_11, u1_L5_12, u1_L5_13, u1_L5_14, u1_L5_15, u1_L5_16, u1_L5_17, u1_L5_18, u1_L5_19, 
        u1_L5_2, u1_L5_20, u1_L5_21, u1_L5_22, u1_L5_23, u1_L5_24, u1_L5_25, u1_L5_26, u1_L5_27, 
        u1_L5_28, u1_L5_29, u1_L5_3, u1_L5_30, u1_L5_31, u1_L5_32, u1_L5_4, u1_L5_5, u1_L5_6, 
        u1_L5_7, u1_L5_8, u1_L5_9, u1_L6_1, u1_L6_10, u1_L6_11, u1_L6_12, u1_L6_13, u1_L6_14, 
        u1_L6_15, u1_L6_16, u1_L6_17, u1_L6_18, u1_L6_19, u1_L6_2, u1_L6_20, u1_L6_21, u1_L6_22, 
        u1_L6_23, u1_L6_24, u1_L6_25, u1_L6_26, u1_L6_27, u1_L6_28, u1_L6_29, u1_L6_3, u1_L6_30, 
        u1_L6_31, u1_L6_32, u1_L6_4, u1_L6_5, u1_L6_6, u1_L6_7, u1_L6_8, u1_L6_9, u1_L7_1, 
        u1_L7_10, u1_L7_11, u1_L7_12, u1_L7_13, u1_L7_14, u1_L7_15, u1_L7_16, u1_L7_17, u1_L7_18, 
        u1_L7_19, u1_L7_2, u1_L7_20, u1_L7_21, u1_L7_22, u1_L7_23, u1_L7_24, u1_L7_25, u1_L7_26, 
        u1_L7_27, u1_L7_28, u1_L7_29, u1_L7_3, u1_L7_30, u1_L7_31, u1_L7_32, u1_L7_4, u1_L7_5, 
        u1_L7_6, u1_L7_7, u1_L7_8, u1_L7_9, u1_L8_1, u1_L8_10, u1_L8_11, u1_L8_12, u1_L8_13, 
        u1_L8_14, u1_L8_15, u1_L8_16, u1_L8_17, u1_L8_18, u1_L8_19, u1_L8_2, u1_L8_20, u1_L8_21, 
        u1_L8_22, u1_L8_23, u1_L8_24, u1_L8_25, u1_L8_26, u1_L8_27, u1_L8_28, u1_L8_29, u1_L8_3, 
        u1_L8_30, u1_L8_31, u1_L8_32, u1_L8_4, u1_L8_5, u1_L8_6, u1_L8_7, u1_L8_8, u1_L8_9, 
        u1_L9_1, u1_L9_10, u1_L9_11, u1_L9_12, u1_L9_13, u1_L9_14, u1_L9_15, u1_L9_16, u1_L9_17, 
        u1_L9_18, u1_L9_19, u1_L9_2, u1_L9_20, u1_L9_21, u1_L9_22, u1_L9_23, u1_L9_24, u1_L9_25, 
        u1_L9_26, u1_L9_27, u1_L9_28, u1_L9_29, u1_L9_3, u1_L9_30, u1_L9_31, u1_L9_32, u1_L9_4, 
        u1_L9_5, u1_L9_6, u1_L9_7, u1_L9_8, u1_L9_9, u1_R0_1, u1_R0_10, u1_R0_11, u1_R0_12, 
        u1_R0_13, u1_R0_14, u1_R0_15, u1_R0_16, u1_R0_17, u1_R0_18, u1_R0_19, u1_R0_2, u1_R0_20, 
        u1_R0_21, u1_R0_22, u1_R0_23, u1_R0_24, u1_R0_25, u1_R0_26, u1_R0_27, u1_R0_28, u1_R0_29, 
        u1_R0_3, u1_R0_30, u1_R0_31, u1_R0_32, u1_R0_4, u1_R0_5, u1_R0_6, u1_R0_7, u1_R0_8, 
        u1_R0_9, u1_R10_1, u1_R10_10, u1_R10_11, u1_R10_12, u1_R10_13, u1_R10_14, u1_R10_15, u1_R10_16, 
        u1_R10_17, u1_R10_18, u1_R10_19, u1_R10_2, u1_R10_20, u1_R10_21, u1_R10_22, u1_R10_23, u1_R10_24, 
        u1_R10_25, u1_R10_26, u1_R10_27, u1_R10_28, u1_R10_29, u1_R10_3, u1_R10_30, u1_R10_31, u1_R10_32, 
        u1_R10_4, u1_R10_5, u1_R10_6, u1_R10_7, u1_R10_8, u1_R10_9, u1_R11_1, u1_R11_10, u1_R11_11, 
        u1_R11_12, u1_R11_13, u1_R11_14, u1_R11_15, u1_R11_16, u1_R11_17, u1_R11_18, u1_R11_19, u1_R11_2, 
        u1_R11_20, u1_R11_21, u1_R11_22, u1_R11_23, u1_R11_24, u1_R11_25, u1_R11_26, u1_R11_27, u1_R11_28, 
        u1_R11_29, u1_R11_3, u1_R11_30, u1_R11_31, u1_R11_32, u1_R11_4, u1_R11_5, u1_R11_6, u1_R11_7, 
        u1_R11_8, u1_R11_9, u1_R12_1, u1_R12_10, u1_R12_11, u1_R12_12, u1_R12_13, u1_R12_14, u1_R12_15, 
        u1_R12_16, u1_R12_17, u1_R12_18, u1_R12_19, u1_R12_2, u1_R12_20, u1_R12_21, u1_R12_22, u1_R12_23, 
        u1_R12_24, u1_R12_25, u1_R12_26, u1_R12_27, u1_R12_28, u1_R12_29, u1_R12_3, u1_R12_30, u1_R12_31, 
        u1_R12_32, u1_R12_4, u1_R12_5, u1_R12_6, u1_R12_7, u1_R12_8, u1_R12_9, u1_R13_1, u1_R13_10, 
        u1_R13_11, u1_R13_12, u1_R13_13, u1_R13_14, u1_R13_15, u1_R13_16, u1_R13_17, u1_R13_18, u1_R13_19, 
        u1_R13_2, u1_R13_20, u1_R13_21, u1_R13_22, u1_R13_23, u1_R13_24, u1_R13_25, u1_R13_26, u1_R13_27, 
        u1_R13_28, u1_R13_29, u1_R13_3, u1_R13_30, u1_R13_31, u1_R13_32, u1_R13_4, u1_R13_5, u1_R13_6, 
        u1_R13_7, u1_R13_8, u1_R13_9, u1_R1_1, u1_R1_10, u1_R1_11, u1_R1_12, u1_R1_13, u1_R1_14, 
        u1_R1_15, u1_R1_16, u1_R1_17, u1_R1_18, u1_R1_19, u1_R1_2, u1_R1_20, u1_R1_21, u1_R1_22, 
        u1_R1_23, u1_R1_24, u1_R1_25, u1_R1_26, u1_R1_27, u1_R1_28, u1_R1_29, u1_R1_3, u1_R1_30, 
        u1_R1_31, u1_R1_32, u1_R1_4, u1_R1_5, u1_R1_6, u1_R1_7, u1_R1_8, u1_R1_9, u1_R2_1, 
        u1_R2_10, u1_R2_11, u1_R2_12, u1_R2_13, u1_R2_14, u1_R2_15, u1_R2_16, u1_R2_17, u1_R2_18, 
        u1_R2_19, u1_R2_2, u1_R2_20, u1_R2_21, u1_R2_22, u1_R2_23, u1_R2_24, u1_R2_25, u1_R2_26, 
        u1_R2_27, u1_R2_28, u1_R2_29, u1_R2_3, u1_R2_30, u1_R2_31, u1_R2_32, u1_R2_4, u1_R2_5, 
        u1_R2_6, u1_R2_7, u1_R2_8, u1_R2_9, u1_R3_1, u1_R3_10, u1_R3_11, u1_R3_12, u1_R3_13, 
        u1_R3_14, u1_R3_15, u1_R3_16, u1_R3_17, u1_R3_18, u1_R3_19, u1_R3_2, u1_R3_20, u1_R3_21, 
        u1_R3_22, u1_R3_23, u1_R3_24, u1_R3_25, u1_R3_26, u1_R3_27, u1_R3_28, u1_R3_29, u1_R3_3, 
        u1_R3_30, u1_R3_31, u1_R3_32, u1_R3_4, u1_R3_5, u1_R3_6, u1_R3_7, u1_R3_8, u1_R3_9, 
        u1_R4_1, u1_R4_10, u1_R4_11, u1_R4_12, u1_R4_13, u1_R4_14, u1_R4_15, u1_R4_16, u1_R4_17, 
        u1_R4_18, u1_R4_19, u1_R4_2, u1_R4_20, u1_R4_21, u1_R4_22, u1_R4_23, u1_R4_24, u1_R4_25, 
        u1_R4_26, u1_R4_27, u1_R4_28, u1_R4_29, u1_R4_3, u1_R4_30, u1_R4_31, u1_R4_32, u1_R4_4, 
        u1_R4_5, u1_R4_6, u1_R4_7, u1_R4_8, u1_R4_9, u1_R5_1, u1_R5_10, u1_R5_11, u1_R5_12, 
        u1_R5_13, u1_R5_14, u1_R5_15, u1_R5_16, u1_R5_17, u1_R5_18, u1_R5_19, u1_R5_2, u1_R5_20, 
        u1_R5_21, u1_R5_22, u1_R5_23, u1_R5_24, u1_R5_25, u1_R5_26, u1_R5_27, u1_R5_28, u1_R5_29, 
        u1_R5_3, u1_R5_30, u1_R5_31, u1_R5_32, u1_R5_4, u1_R5_5, u1_R5_6, u1_R5_7, u1_R5_8, 
        u1_R5_9, u1_R6_1, u1_R6_10, u1_R6_11, u1_R6_12, u1_R6_13, u1_R6_14, u1_R6_15, u1_R6_16, 
        u1_R6_17, u1_R6_18, u1_R6_19, u1_R6_2, u1_R6_20, u1_R6_21, u1_R6_22, u1_R6_23, u1_R6_24, 
        u1_R6_25, u1_R6_26, u1_R6_27, u1_R6_28, u1_R6_29, u1_R6_3, u1_R6_30, u1_R6_31, u1_R6_32, 
        u1_R6_4, u1_R6_5, u1_R6_6, u1_R6_7, u1_R6_8, u1_R6_9, u1_R7_1, u1_R7_10, u1_R7_11, 
        u1_R7_12, u1_R7_13, u1_R7_14, u1_R7_15, u1_R7_16, u1_R7_17, u1_R7_18, u1_R7_19, u1_R7_2, 
        u1_R7_20, u1_R7_21, u1_R7_22, u1_R7_23, u1_R7_24, u1_R7_25, u1_R7_26, u1_R7_27, u1_R7_28, 
        u1_R7_29, u1_R7_3, u1_R7_30, u1_R7_31, u1_R7_32, u1_R7_4, u1_R7_5, u1_R7_6, u1_R7_7, 
        u1_R7_8, u1_R7_9, u1_R8_1, u1_R8_10, u1_R8_11, u1_R8_12, u1_R8_13, u1_R8_14, u1_R8_15, 
        u1_R8_16, u1_R8_17, u1_R8_18, u1_R8_19, u1_R8_2, u1_R8_20, u1_R8_21, u1_R8_22, u1_R8_23, 
        u1_R8_24, u1_R8_25, u1_R8_26, u1_R8_27, u1_R8_28, u1_R8_29, u1_R8_3, u1_R8_30, u1_R8_31, 
        u1_R8_32, u1_R8_4, u1_R8_5, u1_R8_6, u1_R8_7, u1_R8_8, u1_R8_9, u1_R9_1, u1_R9_10, 
        u1_R9_11, u1_R9_12, u1_R9_13, u1_R9_14, u1_R9_15, u1_R9_16, u1_R9_17, u1_R9_18, u1_R9_19, 
        u1_R9_2, u1_R9_20, u1_R9_21, u1_R9_22, u1_R9_23, u1_R9_24, u1_R9_25, u1_R9_26, u1_R9_27, 
        u1_R9_28, u1_R9_29, u1_R9_3, u1_R9_30, u1_R9_31, u1_R9_32, u1_R9_4, u1_R9_5, u1_R9_6, 
        u1_R9_7, u1_R9_8, u1_R9_9, u1_desIn_r_0, u1_desIn_r_1, u1_desIn_r_10, u1_desIn_r_11, u1_desIn_r_12, u1_desIn_r_13, 
        u1_desIn_r_14, u1_desIn_r_15, u1_desIn_r_16, u1_desIn_r_17, u1_desIn_r_18, u1_desIn_r_19, u1_desIn_r_2, u1_desIn_r_20, u1_desIn_r_21, 
        u1_desIn_r_22, u1_desIn_r_23, u1_desIn_r_24, u1_desIn_r_25, u1_desIn_r_26, u1_desIn_r_27, u1_desIn_r_28, u1_desIn_r_29, u1_desIn_r_3, 
        u1_desIn_r_30, u1_desIn_r_31, u1_desIn_r_32, u1_desIn_r_33, u1_desIn_r_34, u1_desIn_r_35, u1_desIn_r_36, u1_desIn_r_37, u1_desIn_r_38, 
        u1_desIn_r_39, u1_desIn_r_4, u1_desIn_r_40, u1_desIn_r_41, u1_desIn_r_42, u1_desIn_r_43, u1_desIn_r_44, u1_desIn_r_45, u1_desIn_r_46, 
        u1_desIn_r_47, u1_desIn_r_48, u1_desIn_r_49, u1_desIn_r_5, u1_desIn_r_50, u1_desIn_r_51, u1_desIn_r_52, u1_desIn_r_53, u1_desIn_r_54, 
        u1_desIn_r_55, u1_desIn_r_56, u1_desIn_r_57, u1_desIn_r_58, u1_desIn_r_59, u1_desIn_r_6, u1_desIn_r_60, u1_desIn_r_61, u1_desIn_r_62, 
        u1_desIn_r_63, u1_desIn_r_7, u1_desIn_r_8, u1_desIn_r_9, u1_key_r_0, u1_key_r_1, u1_key_r_10, u1_key_r_11, u1_key_r_12, 
        u1_key_r_13, u1_key_r_14, u1_key_r_15, u1_key_r_16, u1_key_r_17, u1_key_r_18, u1_key_r_19, u1_key_r_2, u1_key_r_20, 
        u1_key_r_21, u1_key_r_22, u1_key_r_23, u1_key_r_24, u1_key_r_25, u1_key_r_26, u1_key_r_27, u1_key_r_28, u1_key_r_29, 
        u1_key_r_3, u1_key_r_30, u1_key_r_31, u1_key_r_32, u1_key_r_33, u1_key_r_34, u1_key_r_35, u1_key_r_36, u1_key_r_37, 
        u1_key_r_38, u1_key_r_39, u1_key_r_4, u1_key_r_40, u1_key_r_41, u1_key_r_42, u1_key_r_43, u1_key_r_44, u1_key_r_45, 
        u1_key_r_46, u1_key_r_47, u1_key_r_48, u1_key_r_49, u1_key_r_5, u1_key_r_50, u1_key_r_51, u1_key_r_52, u1_key_r_53, 
        u1_key_r_54, u1_key_r_55, u1_key_r_6, u1_key_r_7, u1_key_r_8, u1_key_r_9, u1_uk_K_r0_11, u1_uk_K_r0_13, u1_uk_K_r0_15, 
        u1_uk_K_r0_17, u1_uk_K_r0_19, u1_uk_K_r0_2, u1_uk_K_r0_22, u1_uk_K_r0_25, u1_uk_K_r0_28, u1_uk_K_r0_31, u1_uk_K_r0_32, u1_uk_K_r0_34, 
        u1_uk_K_r0_36, u1_uk_K_r0_47, u1_uk_K_r0_49, u1_uk_K_r0_52, u1_uk_K_r0_55, u1_uk_K_r0_7, u1_uk_K_r10_10, u1_uk_K_r10_11, u1_uk_K_r10_14, 
        u1_uk_K_r10_16, u1_uk_K_r10_18, u1_uk_K_r10_19, u1_uk_K_r10_23, u1_uk_K_r10_25, u1_uk_K_r10_27, u1_uk_K_r10_28, u1_uk_K_r10_32, u1_uk_K_r10_34, 
        u1_uk_K_r10_37, u1_uk_K_r10_39, u1_uk_K_r10_4, u1_uk_K_r10_41, u1_uk_K_r10_42, u1_uk_K_r10_43, u1_uk_K_r10_44, u1_uk_K_r10_47, u1_uk_K_r10_48, 
        u1_uk_K_r10_49, u1_uk_K_r10_52, u1_uk_K_r10_9, u1_uk_K_r11_10, u1_uk_K_r11_11, u1_uk_K_r11_17, u1_uk_K_r11_19, u1_uk_K_r11_20, u1_uk_K_r11_21, 
        u1_uk_K_r11_24, u1_uk_K_r11_25, u1_uk_K_r11_26, u1_uk_K_r11_27, u1_uk_K_r11_28, u1_uk_K_r11_29, u1_uk_K_r11_33, u1_uk_K_r11_34, u1_uk_K_r11_39, 
        u1_uk_K_r11_4, u1_uk_K_r11_46, u1_uk_K_r11_47, u1_uk_K_r11_48, u1_uk_K_r11_5, u1_uk_K_r11_53, u1_uk_K_r11_54, u1_uk_K_r11_6, u1_uk_K_r11_7, 
        u1_uk_K_r11_8, u1_uk_K_r12_1, u1_uk_K_r12_10, u1_uk_K_r12_15, u1_uk_K_r12_16, u1_uk_K_r12_18, u1_uk_K_r12_21, u1_uk_K_r12_22, u1_uk_K_r12_25, 
        u1_uk_K_r12_30, u1_uk_K_r12_33, u1_uk_K_r12_36, u1_uk_K_r12_41, u1_uk_K_r12_42, u1_uk_K_r12_44, u1_uk_K_r12_47, u1_uk_K_r12_7, u1_uk_K_r13_0, 
        u1_uk_K_r13_13, u1_uk_K_r13_17, u1_uk_K_r13_19, u1_uk_K_r13_2, u1_uk_K_r13_22, u1_uk_K_r13_23, u1_uk_K_r13_25, u1_uk_K_r13_31, u1_uk_K_r13_32, 
        u1_uk_K_r13_35, u1_uk_K_r13_36, u1_uk_K_r13_38, u1_uk_K_r13_4, u1_uk_K_r13_44, u1_uk_K_r13_55, u1_uk_K_r14_10, u1_uk_K_r14_11, u1_uk_K_r14_12, 
        u1_uk_K_r14_15, u1_uk_K_r14_16, u1_uk_K_r14_18, u1_uk_K_r14_2, u1_uk_K_r14_23, u1_uk_K_r14_3, u1_uk_K_r14_38, u1_uk_K_r14_39, u1_uk_K_r14_42, 
        u1_uk_K_r14_43, u1_uk_K_r14_45, u1_uk_K_r14_46, u1_uk_K_r14_5, u1_uk_K_r14_50, u1_uk_K_r14_8, u1_uk_K_r14_9, u1_uk_K_r1_10, u1_uk_K_r1_15, 
        u1_uk_K_r1_16, u1_uk_K_r1_17, u1_uk_K_r1_18, u1_uk_K_r1_21, u1_uk_K_r1_22, u1_uk_K_r1_33, u1_uk_K_r1_36, u1_uk_K_r1_41, u1_uk_K_r1_42, 
        u1_uk_K_r1_44, u1_uk_K_r1_47, u1_uk_K_r1_6, u1_uk_K_r1_7, u1_uk_K_r2_13, u1_uk_K_r2_16, u1_uk_K_r2_18, u1_uk_K_r2_20, u1_uk_K_r2_21, 
        u1_uk_K_r2_24, u1_uk_K_r2_25, u1_uk_K_r2_26, u1_uk_K_r2_27, u1_uk_K_r2_28, u1_uk_K_r2_29, u1_uk_K_r2_31, u1_uk_K_r2_33, u1_uk_K_r2_36, 
        u1_uk_K_r2_4, u1_uk_K_r2_41, u1_uk_K_r2_46, u1_uk_K_r2_47, u1_uk_K_r2_49, u1_uk_K_r2_50, u1_uk_K_r2_53, u1_uk_K_r2_55, u1_uk_K_r2_6, 
        u1_uk_K_r2_7, u1_uk_K_r3_10, u1_uk_K_r3_11, u1_uk_K_r3_14, u1_uk_K_r3_15, u1_uk_K_r3_16, u1_uk_K_r3_19, u1_uk_K_r3_24, u1_uk_K_r3_29, 
        u1_uk_K_r3_33, u1_uk_K_r3_34, u1_uk_K_r3_35, u1_uk_K_r3_38, u1_uk_K_r3_4, u1_uk_K_r3_43, u1_uk_K_r3_44, u1_uk_K_r3_47, u1_uk_K_r3_51, 
        u1_uk_K_r3_52, u1_uk_K_r3_9, u1_uk_K_r4_0, u1_uk_K_r4_11, u1_uk_K_r4_17, u1_uk_K_r4_18, u1_uk_K_r4_23, u1_uk_K_r4_27, u1_uk_K_r4_3, 
        u1_uk_K_r4_31, u1_uk_K_r4_33, u1_uk_K_r4_35, u1_uk_K_r4_38, u1_uk_K_r4_4, u1_uk_K_r4_41, u1_uk_K_r4_47, u1_uk_K_r4_48, u1_uk_K_r4_49, 
        u1_uk_K_r4_5, u1_uk_K_r4_54, u1_uk_K_r4_55, u1_uk_K_r5_0, u1_uk_K_r5_1, u1_uk_K_r5_10, u1_uk_K_r5_13, u1_uk_K_r5_16, u1_uk_K_r5_17, 
        u1_uk_K_r5_18, u1_uk_K_r5_19, u1_uk_K_r5_21, u1_uk_K_r5_23, u1_uk_K_r5_26, u1_uk_K_r5_31, u1_uk_K_r5_32, u1_uk_K_r5_35, u1_uk_K_r5_36, 
        u1_uk_K_r5_37, u1_uk_K_r5_39, u1_uk_K_r5_4, u1_uk_K_r5_40, u1_uk_K_r5_41, u1_uk_K_r5_43, u1_uk_K_r5_48, u1_uk_K_r5_5, u1_uk_K_r5_51, 
        u1_uk_K_r5_53, u1_uk_K_r5_7, u1_uk_K_r5_8, u1_uk_K_r6_0, u1_uk_K_r6_10, u1_uk_K_r6_14, u1_uk_K_r6_17, u1_uk_K_r6_19, u1_uk_K_r6_21, 
        u1_uk_K_r6_22, u1_uk_K_r6_26, u1_uk_K_r6_27, u1_uk_K_r6_28, u1_uk_K_r6_29, u1_uk_K_r6_3, u1_uk_K_r6_30, u1_uk_K_r6_31, u1_uk_K_r6_34, 
        u1_uk_K_r6_35, u1_uk_K_r6_37, u1_uk_K_r6_46, u1_uk_K_r6_51, u1_uk_K_r6_53, u1_uk_K_r6_55, u1_uk_K_r6_7, u1_uk_K_r7_0, u1_uk_K_r7_1, 
        u1_uk_K_r7_13, u1_uk_K_r7_15, u1_uk_K_r7_16, u1_uk_K_r7_2, u1_uk_K_r7_20, u1_uk_K_r7_22, u1_uk_K_r7_23, u1_uk_K_r7_24, u1_uk_K_r7_25, 
        u1_uk_K_r7_26, u1_uk_K_r7_27, u1_uk_K_r7_29, u1_uk_K_r7_30, u1_uk_K_r7_31, u1_uk_K_r7_32, u1_uk_K_r7_34, u1_uk_K_r7_37, u1_uk_K_r7_39, 
        u1_uk_K_r7_41, u1_uk_K_r7_46, u1_uk_K_r7_48, u1_uk_K_r7_5, u1_uk_K_r7_53, u1_uk_K_r7_55, u1_uk_K_r7_6, u1_uk_K_r7_7, u1_uk_K_r7_8, 
        u1_uk_K_r7_9, u1_uk_K_r8_10, u1_uk_K_r8_13, u1_uk_K_r8_16, u1_uk_K_r8_17, u1_uk_K_r8_19, u1_uk_K_r8_2, u1_uk_K_r8_21, u1_uk_K_r8_22, 
        u1_uk_K_r8_27, u1_uk_K_r8_28, u1_uk_K_r8_32, u1_uk_K_r8_37, u1_uk_K_r8_39, u1_uk_K_r8_40, u1_uk_K_r8_41, u1_uk_K_r8_42, u1_uk_K_r8_43, 
        u1_uk_K_r8_44, u1_uk_K_r8_48, u1_uk_K_r8_5, u1_uk_K_r8_51, u1_uk_K_r8_52, u1_uk_K_r8_8, u1_uk_K_r9_0, u1_uk_K_r9_1, u1_uk_K_r9_10, 
        u1_uk_K_r9_12, u1_uk_K_r9_13, u1_uk_K_r9_15, u1_uk_K_r9_18, u1_uk_K_r9_19, u1_uk_K_r9_22, u1_uk_K_r9_23, u1_uk_K_r9_25, u1_uk_K_r9_27, 
        u1_uk_K_r9_30, u1_uk_K_r9_31, u1_uk_K_r9_33, u1_uk_K_r9_35, u1_uk_K_r9_38, u1_uk_K_r9_4, u1_uk_K_r9_45, u1_uk_K_r9_48, u1_uk_K_r9_49, 
        u1_uk_K_r9_5, u1_uk_K_r9_54, u1_uk_K_r9_55, u1_uk_K_r9_6, u1_uk_K_r9_7, u1_uk_K_r9_9, u1_uk_n1218, u1_uk_n1219, u1_uk_n1220, 
        u1_uk_n1221, u1_uk_n1222, u1_uk_n1224, u1_uk_n1225, u1_uk_n1227, u1_uk_n1228, u1_uk_n1229, u1_uk_n1230, u1_uk_n1231, 
        u1_uk_n1233, u1_uk_n1234, u1_uk_n1235, u1_uk_n1236, u1_uk_n1237, u1_uk_n1238, u1_uk_n1239, u1_uk_n1240, u1_uk_n1241, 
        u1_uk_n1242, u1_uk_n1243, u1_uk_n1244, u1_uk_n1245, u1_uk_n1246, u1_uk_n1247, u1_uk_n1248, u1_uk_n1249, u1_uk_n1250, 
        u1_uk_n1251, u1_uk_n1252, u1_uk_n1253, u1_uk_n1255, u1_uk_n1256, u1_uk_n1257, u1_uk_n1258, u1_uk_n1259, u1_uk_n1260, 
        u1_uk_n1261, u1_uk_n1262, u1_uk_n1263, u1_uk_n1264, u1_uk_n1265, u1_uk_n1266, u1_uk_n1267, u1_uk_n1268, u1_uk_n1269, 
        u1_uk_n1270, u1_uk_n1271, u1_uk_n1272, u1_uk_n1273, u1_uk_n1274, u1_uk_n1275, u1_uk_n1276, u1_uk_n1277, u1_uk_n1278, 
        u1_uk_n1279, u1_uk_n1281, u1_uk_n1282, u1_uk_n1284, u1_uk_n1286, u1_uk_n1288, u1_uk_n1289, u1_uk_n1290, u1_uk_n1291, 
        u1_uk_n1292, u1_uk_n1293, u1_uk_n1294, u1_uk_n1295, u1_uk_n1296, u1_uk_n1297, u1_uk_n1299, u1_uk_n1300, u1_uk_n1303, 
        u1_uk_n1304, u1_uk_n1305, u1_uk_n1307, u1_uk_n1308, u1_uk_n1309, u1_uk_n1310, u1_uk_n1311, u1_uk_n1312, u1_uk_n1313, 
        u1_uk_n1314, u1_uk_n1315, u1_uk_n1316, u1_uk_n1317, u1_uk_n1318, u1_uk_n1319, u1_uk_n1320, u1_uk_n1321, u1_uk_n1322, 
        u1_uk_n1323, u1_uk_n1324, u1_uk_n1325, u1_uk_n1326, u1_uk_n1327, u1_uk_n1328, u1_uk_n1329, u1_uk_n1330, u1_uk_n1331, 
        u1_uk_n1332, u1_uk_n1333, u1_uk_n1334, u1_uk_n1335, u1_uk_n1336, u1_uk_n1338, u1_uk_n1339, u1_uk_n1340, u1_uk_n1341, 
        u1_uk_n1342, u1_uk_n1343, u1_uk_n1344, u1_uk_n1345, u1_uk_n1346, u1_uk_n1347, u1_uk_n1348, u1_uk_n1349, u1_uk_n1350, 
        u1_uk_n1351, u1_uk_n1352, u1_uk_n1353, u1_uk_n1354, u1_uk_n1355, u1_uk_n1356, u1_uk_n1357, u1_uk_n1358, u1_uk_n1359, 
        u1_uk_n1360, u1_uk_n1361, u1_uk_n1363, u1_uk_n1365, u1_uk_n1366, u1_uk_n1367, u1_uk_n1369, u1_uk_n1371, u1_uk_n1372, 
        u1_uk_n1374, u1_uk_n1375, u1_uk_n1376, u1_uk_n1377, u1_uk_n1378, u1_uk_n1380, u1_uk_n1381, u1_uk_n1382, u1_uk_n1383, 
        u1_uk_n1386, u1_uk_n1389, u1_uk_n1390, u1_uk_n1391, u1_uk_n1393, u1_uk_n1394, u1_uk_n1395, u1_uk_n1396, u1_uk_n1397, 
        u1_uk_n1398, u1_uk_n1399, u1_uk_n1400, u1_uk_n1401, u1_uk_n1402, u1_uk_n1403, u1_uk_n1404, u1_uk_n1405, u1_uk_n1406, 
        u1_uk_n1407, u1_uk_n1408, u1_uk_n1409, u1_uk_n1410, u1_uk_n1411, u1_uk_n1412, u1_uk_n1413, u1_uk_n1414, u1_uk_n1415, 
        u1_uk_n1417, u1_uk_n1418, u1_uk_n1419, u1_uk_n1422, u1_uk_n1423, u1_uk_n1424, u1_uk_n1425, u1_uk_n1426, u1_uk_n1427, 
        u1_uk_n1429, u1_uk_n1430, u1_uk_n1431, u1_uk_n1433, u1_uk_n1435, u1_uk_n1436, u1_uk_n1437, u1_uk_n1438, u1_uk_n1439, 
        u1_uk_n1440, u1_uk_n1441, u1_uk_n1442, u1_uk_n1443, u1_uk_n1444, u1_uk_n1446, u1_uk_n1447, u1_uk_n1448, u1_uk_n1449, 
        u1_uk_n1450, u1_uk_n1452, u1_uk_n1453, u1_uk_n1454, u1_uk_n1455, u1_uk_n1456, u1_uk_n1457, u1_uk_n1458, u1_uk_n1459, 
        u1_uk_n1460, u1_uk_n1461, u1_uk_n1462, u1_uk_n1463, u1_uk_n1464, u1_uk_n1465, u1_uk_n1466, u1_uk_n1468, u1_uk_n1469, 
        u1_uk_n1470, u1_uk_n1471, u1_uk_n1472, u1_uk_n1474, u1_uk_n1475, u1_uk_n1476, u1_uk_n1477, u1_uk_n1478, u1_uk_n1482, 
        u1_uk_n1483, u1_uk_n1484, u1_uk_n1485, u1_uk_n1486, u1_uk_n1487, u1_uk_n1488, u1_uk_n1489, u1_uk_n1490, u1_uk_n1491, 
        u1_uk_n1492, u1_uk_n1494, u1_uk_n1495, u1_uk_n1496, u1_uk_n1498, u1_uk_n1499, u1_uk_n1500, u1_uk_n1501, u1_uk_n1504, 
        u1_uk_n1505, u1_uk_n1507, u1_uk_n1508, u1_uk_n1510, u1_uk_n1514, u1_uk_n1516, u1_uk_n1517, u1_uk_n1518, u1_uk_n1520, 
        u1_uk_n1521, u1_uk_n1523, u1_uk_n1524, u1_uk_n1526, u1_uk_n1527, u1_uk_n1528, u1_uk_n1529, u1_uk_n1530, u1_uk_n1531, 
        u1_uk_n1532, u1_uk_n1533, u1_uk_n1534, u1_uk_n1536, u1_uk_n1537, u1_uk_n1538, u1_uk_n1540, u1_uk_n1541, u1_uk_n1543, 
        u1_uk_n1544, u1_uk_n1545, u1_uk_n1547, u1_uk_n1548, u1_uk_n1549, u1_uk_n1551, u1_uk_n1552, u1_uk_n1554, u1_uk_n1555, 
        u1_uk_n1556, u1_uk_n1557, u1_uk_n1558, u1_uk_n1559, u1_uk_n1560, u1_uk_n1561, u1_uk_n1562, u1_uk_n1563, u1_uk_n1564, 
        u1_uk_n1565, u1_uk_n1566, u1_uk_n1567, u1_uk_n1568, u1_uk_n1570, u1_uk_n1571, u1_uk_n1572, u1_uk_n1573, u1_uk_n1574, 
        u1_uk_n1577, u1_uk_n1578, u1_uk_n1579, u1_uk_n1581, u1_uk_n1584, u1_uk_n1585, u1_uk_n1586, u1_uk_n1588, u1_uk_n1592, 
        u1_uk_n1593, u1_uk_n1595, u1_uk_n1598, u1_uk_n1599, u1_uk_n1600, u1_uk_n1601, u1_uk_n1603, u1_uk_n1604, u1_uk_n1605, 
        u1_uk_n1606, u1_uk_n1607, u1_uk_n1608, u1_uk_n1610, u1_uk_n1612, u1_uk_n1613, u1_uk_n1614, u1_uk_n1615, u1_uk_n1616, 
        u1_uk_n1618, u1_uk_n1619, u1_uk_n1620, u1_uk_n1621, u1_uk_n1622, u1_uk_n1623, u1_uk_n1624, u1_uk_n1625, u1_uk_n1626, 
        u1_uk_n1627, u1_uk_n1628, u1_uk_n1629, u1_uk_n1630, u1_uk_n1632, u1_uk_n1633, u1_uk_n1634, u1_uk_n1635, u1_uk_n1639, 
        u1_uk_n1640, u1_uk_n1641, u1_uk_n1642, u1_uk_n1643, u1_uk_n1644, u1_uk_n1645, u1_uk_n1647, u1_uk_n1649, u1_uk_n1651, 
        u1_uk_n1652, u1_uk_n1653, u1_uk_n1654, u1_uk_n1655, u1_uk_n1656, u1_uk_n1659, u1_uk_n1660, u1_uk_n1661, u1_uk_n1662, 
        u1_uk_n1663, u1_uk_n1664, u1_uk_n1667, u1_uk_n1669, u1_uk_n1670, u1_uk_n1672, u1_uk_n1673, u1_uk_n1676, u1_uk_n1677, 
        u1_uk_n1678, u1_uk_n1682, u1_uk_n1683, u1_uk_n1684, u1_uk_n1687, u1_uk_n1688, u1_uk_n1689, u1_uk_n1690, u1_uk_n1691, 
        u1_uk_n1692, u1_uk_n1693, u1_uk_n1694, u1_uk_n1695, u1_uk_n1696, u1_uk_n1698, u1_uk_n1699, u1_uk_n1702, u1_uk_n1703, 
        u1_uk_n1704, u1_uk_n1705, u1_uk_n1707, u1_uk_n1708, u1_uk_n1709, u1_uk_n1710, u1_uk_n1711, u1_uk_n1712, u1_uk_n1713, 
        u1_uk_n1714, u1_uk_n1715, u1_uk_n1716, u1_uk_n1717, u1_uk_n1718, u1_uk_n1719, u1_uk_n1720, u1_uk_n1721, u1_uk_n1722, 
        u1_uk_n1723, u1_uk_n1728, u1_uk_n1729, u1_uk_n1730, u1_uk_n1731, u1_uk_n1732, u1_uk_n1734, u1_uk_n1735, u1_uk_n1736, 
        u1_uk_n1737, u1_uk_n1738, u1_uk_n1739, u1_uk_n1744, u1_uk_n1745, u1_uk_n1748, u1_uk_n1749, u1_uk_n1750, u1_uk_n1751, 
        u1_uk_n1752, u1_uk_n1753, u1_uk_n1754, u1_uk_n1755, u1_uk_n1756, u1_uk_n1757, u1_uk_n1758, u1_uk_n1761, u1_uk_n1762, 
        u1_uk_n1763, u1_uk_n1764, u1_uk_n1765, u1_uk_n1766, u1_uk_n1767, u1_uk_n1768, u1_uk_n1769, u1_uk_n1772, u1_uk_n1773, 
        u1_uk_n1774, u1_uk_n1775, u1_uk_n1776, u1_uk_n1777, u1_uk_n1780, u1_uk_n1781, u1_uk_n1782, u1_uk_n1783, u1_uk_n1784, 
        u1_uk_n1785, u1_uk_n1787, u1_uk_n1790, u1_uk_n1791, u1_uk_n1792, u1_uk_n1793, u1_uk_n1797, u1_uk_n1798, u1_uk_n1799, 
        u1_uk_n1800, u1_uk_n1801, u1_uk_n1802, u1_uk_n1803, u1_uk_n1804, u1_uk_n1806, u1_uk_n1807, u1_uk_n1808, u1_uk_n1809, 
        u1_uk_n1810, u1_uk_n1811, u1_uk_n1812, u1_uk_n1813, u1_uk_n1814, u1_uk_n1815, u1_uk_n1816, u1_uk_n1817, u1_uk_n1818, 
        u1_uk_n1819, u1_uk_n1820, u1_uk_n1821, u1_uk_n1822, u1_uk_n1823, u1_uk_n1824, u1_uk_n1826, u1_uk_n1827, u1_uk_n1829, 
        u1_uk_n1830, u1_uk_n1831, u1_uk_n1832, u1_uk_n1833, u1_uk_n1834, u1_uk_n1835, u1_uk_n1836, u1_uk_n1837, u1_uk_n1838, 
        u1_uk_n1839, u1_uk_n1840, u1_uk_n1841, u1_uk_n1842, u1_uk_n1843, u1_uk_n1844, u1_uk_n1845, u1_uk_n1846, u1_uk_n1847, 
        u1_uk_n1848, u1_uk_n1849, u1_uk_n1850, u1_uk_n1851, u1_uk_n1852, u1_uk_n1853, u1_uk_n1854, u1_uk_n1855, u1_uk_n1856, 
        u1_uk_n1858, u1_uk_n1859, u1_uk_n1860, u1_uk_n1862, u1_uk_n1863, u1_uk_n1864, u1_uk_n1865, u1_uk_n1866, u1_uk_n1867, 
        u1_uk_n1868, u1_uk_n1869, u1_uk_n1870, u1_uk_n1872, u1_uk_n1873, u1_uk_n1874, u1_uk_n1875, u1_uk_n1876, u1_uk_n1879, 
        u1_uk_n1880, u1_uk_n1881, u1_uk_n1882, u1_uk_n1883, u1_uk_n1884, u1_uk_n1885, u1_uk_n1886, u1_uk_n1887, u2_FP_33, 
        u2_FP_34, u2_FP_35, u2_FP_36, u2_FP_37, u2_FP_38, u2_FP_39, u2_FP_40, u2_FP_41, u2_FP_42, 
        u2_FP_43, u2_FP_44, u2_FP_45, u2_FP_46, u2_FP_47, u2_FP_48, u2_FP_49, u2_FP_50, u2_FP_51, 
        u2_FP_52, u2_FP_53, u2_FP_54, u2_FP_55, u2_FP_56, u2_FP_57, u2_FP_58, u2_FP_59, u2_FP_60, 
        u2_FP_61, u2_FP_62, u2_FP_63, u2_FP_64, u2_K10_10, u2_K10_11, u2_K10_15, u2_K10_17, u2_K10_25, 
        u2_K10_26, u2_K10_30, u2_K10_32, u2_K10_34, u2_K10_36, u2_K10_4, u2_K10_42, u2_K10_43, u2_K10_44, 
        u2_K10_46, u2_K10_6, u2_K11_11, u2_K11_13, u2_K11_16, u2_K11_18, u2_K11_21, u2_K11_29, u2_K11_38, 
        u2_K11_4, u2_K11_42, u2_K11_45, u2_K11_48, u2_K11_6, u2_K11_7, u2_K11_9, u2_K12_2, u2_K12_20, 
        u2_K12_22, u2_K12_24, u2_K12_25, u2_K12_26, u2_K12_27, u2_K12_29, u2_K12_34, u2_K12_37, u2_K12_41, 
        u2_K12_46, u2_K12_47, u2_K12_8, u2_K13_14, u2_K13_20, u2_K13_26, u2_K13_3, u2_K13_31, u2_K13_32, 
        u2_K13_34, u2_K13_37, u2_K13_40, u2_K13_42, u2_K13_44, u2_K13_45, u2_K13_46, u2_K13_47, u2_K13_8, 
        u2_K14_10, u2_K14_11, u2_K14_12, u2_K14_13, u2_K14_14, u2_K14_16, u2_K14_17, u2_K14_18, u2_K14_21, 
        u2_K14_25, u2_K14_28, u2_K14_3, u2_K14_39, u2_K14_42, u2_K14_6, u2_K14_8, u2_K15_1, u2_K15_13, 
        u2_K15_16, u2_K15_18, u2_K15_2, u2_K15_20, u2_K15_21, u2_K15_23, u2_K15_28, u2_K15_29, u2_K15_31, 
        u2_K15_34, u2_K15_35, u2_K15_39, u2_K15_5, u2_K16_26, u2_K16_31, u2_K16_42, u2_K16_44, u2_K16_47, 
        u2_K16_5, u2_K16_6, u2_K16_8, u2_K16_9, u2_K1_15, u2_K1_16, u2_K1_19, u2_K1_24, u2_K1_28, 
        u2_K1_37, u2_K1_40, u2_K1_43, u2_K1_45, u2_K1_46, u2_K1_5, u2_K1_9, u2_K2_1, u2_K2_16, 
        u2_K2_18, u2_K2_20, u2_K2_34, u2_K2_35, u2_K2_36, u2_K2_40, u2_K2_43, u2_K2_44, u2_K2_45, 
        u2_K2_46, u2_K2_47, u2_K2_48, u2_K3_13, u2_K3_15, u2_K3_16, u2_K3_20, u2_K3_23, u2_K3_30, 
        u2_K3_32, u2_K3_35, u2_K3_42, u2_K3_43, u2_K3_47, u2_K3_48, u2_K3_7, u2_K4_14, u2_K4_21, 
        u2_K4_22, u2_K4_27, u2_K4_33, u2_K4_34, u2_K4_35, u2_K4_38, u2_K4_39, u2_K4_42, u2_K4_6, 
        u2_K4_7, u2_K5_1, u2_K5_10, u2_K5_11, u2_K5_13, u2_K5_14, u2_K5_16, u2_K5_17, u2_K5_18, 
        u2_K5_19, u2_K5_21, u2_K5_23, u2_K5_24, u2_K5_25, u2_K5_26, u2_K5_28, u2_K5_3, u2_K5_31, 
        u2_K5_32, u2_K5_34, u2_K5_38, u2_K5_41, u2_K5_44, u2_K5_47, u2_K5_48, u2_K5_5, u2_K5_6, 
        u2_K5_8, u2_K5_9, u2_K6_1, u2_K6_11, u2_K6_13, u2_K6_14, u2_K6_15, u2_K6_16, u2_K6_20, 
        u2_K6_22, u2_K6_24, u2_K6_25, u2_K6_27, u2_K6_3, u2_K6_32, u2_K6_34, u2_K6_36, u2_K6_40, 
        u2_K7_26, u2_K7_3, u2_K7_31, u2_K7_33, u2_K7_35, u2_K7_37, u2_K7_38, u2_K7_4, u2_K7_43, 
        u2_K7_45, u2_K7_48, u2_K7_5, u2_K7_7, u2_K8_18, u2_K8_24, u2_K8_26, u2_K8_31, u2_K8_41, 
        u2_K8_45, u2_K8_5, u2_K8_8, u2_K9_15, u2_K9_23, u2_K9_25, u2_K9_28, u2_K9_29, u2_K9_3, 
        u2_K9_32, u2_K9_36, u2_K9_38, u2_K9_40, u2_K9_45, u2_K9_5, u2_L0_1, u2_L0_10, u2_L0_11, 
        u2_L0_12, u2_L0_13, u2_L0_14, u2_L0_15, u2_L0_16, u2_L0_17, u2_L0_18, u2_L0_19, u2_L0_2, 
        u2_L0_20, u2_L0_21, u2_L0_22, u2_L0_23, u2_L0_24, u2_L0_25, u2_L0_26, u2_L0_27, u2_L0_28, 
        u2_L0_29, u2_L0_3, u2_L0_30, u2_L0_31, u2_L0_32, u2_L0_4, u2_L0_5, u2_L0_6, u2_L0_7, 
        u2_L0_8, u2_L0_9, u2_L10_1, u2_L10_10, u2_L10_11, u2_L10_12, u2_L10_13, u2_L10_14, u2_L10_15, 
        u2_L10_16, u2_L10_17, u2_L10_18, u2_L10_19, u2_L10_2, u2_L10_20, u2_L10_21, u2_L10_22, u2_L10_23, 
        u2_L10_24, u2_L10_25, u2_L10_26, u2_L10_27, u2_L10_28, u2_L10_29, u2_L10_3, u2_L10_30, u2_L10_31, 
        u2_L10_32, u2_L10_4, u2_L10_5, u2_L10_6, u2_L10_7, u2_L10_8, u2_L10_9, u2_L11_1, u2_L11_10, 
        u2_L11_11, u2_L11_12, u2_L11_13, u2_L11_14, u2_L11_15, u2_L11_16, u2_L11_17, u2_L11_18, u2_L11_19, 
        u2_L11_2, u2_L11_20, u2_L11_21, u2_L11_22, u2_L11_23, u2_L11_24, u2_L11_25, u2_L11_26, u2_L11_27, 
        u2_L11_28, u2_L11_29, u2_L11_3, u2_L11_30, u2_L11_31, u2_L11_32, u2_L11_4, u2_L11_5, u2_L11_6, 
        u2_L11_7, u2_L11_8, u2_L11_9, u2_L12_1, u2_L12_10, u2_L12_11, u2_L12_12, u2_L12_13, u2_L12_14, 
        u2_L12_15, u2_L12_16, u2_L12_17, u2_L12_18, u2_L12_19, u2_L12_2, u2_L12_20, u2_L12_21, u2_L12_22, 
        u2_L12_23, u2_L12_24, u2_L12_25, u2_L12_26, u2_L12_27, u2_L12_28, u2_L12_29, u2_L12_3, u2_L12_30, 
        u2_L12_31, u2_L12_32, u2_L12_4, u2_L12_5, u2_L12_6, u2_L12_7, u2_L12_8, u2_L12_9, u2_L13_1, 
        u2_L13_10, u2_L13_11, u2_L13_12, u2_L13_13, u2_L13_14, u2_L13_15, u2_L13_16, u2_L13_17, u2_L13_18, 
        u2_L13_19, u2_L13_2, u2_L13_20, u2_L13_21, u2_L13_22, u2_L13_23, u2_L13_24, u2_L13_25, u2_L13_26, 
        u2_L13_27, u2_L13_28, u2_L13_29, u2_L13_3, u2_L13_30, u2_L13_31, u2_L13_32, u2_L13_4, u2_L13_5, 
        u2_L13_6, u2_L13_7, u2_L13_8, u2_L13_9, u2_L14_1, u2_L14_10, u2_L14_11, u2_L14_12, u2_L14_13, 
        u2_L14_14, u2_L14_15, u2_L14_16, u2_L14_17, u2_L14_18, u2_L14_19, u2_L14_2, u2_L14_20, u2_L14_21, 
        u2_L14_22, u2_L14_23, u2_L14_24, u2_L14_25, u2_L14_26, u2_L14_27, u2_L14_28, u2_L14_29, u2_L14_3, 
        u2_L14_30, u2_L14_31, u2_L14_32, u2_L14_4, u2_L14_5, u2_L14_6, u2_L14_7, u2_L14_8, u2_L14_9, 
        u2_L1_1, u2_L1_10, u2_L1_11, u2_L1_12, u2_L1_13, u2_L1_14, u2_L1_15, u2_L1_16, u2_L1_17, 
        u2_L1_18, u2_L1_19, u2_L1_2, u2_L1_20, u2_L1_21, u2_L1_22, u2_L1_23, u2_L1_24, u2_L1_25, 
        u2_L1_26, u2_L1_27, u2_L1_28, u2_L1_29, u2_L1_3, u2_L1_30, u2_L1_31, u2_L1_32, u2_L1_4, 
        u2_L1_5, u2_L1_6, u2_L1_7, u2_L1_8, u2_L1_9, u2_L2_1, u2_L2_10, u2_L2_11, u2_L2_12, 
        u2_L2_13, u2_L2_14, u2_L2_15, u2_L2_16, u2_L2_17, u2_L2_18, u2_L2_19, u2_L2_2, u2_L2_20, 
        u2_L2_21, u2_L2_22, u2_L2_23, u2_L2_24, u2_L2_25, u2_L2_26, u2_L2_27, u2_L2_28, u2_L2_29, 
        u2_L2_3, u2_L2_30, u2_L2_31, u2_L2_32, u2_L2_4, u2_L2_5, u2_L2_6, u2_L2_7, u2_L2_8, 
        u2_L2_9, u2_L3_1, u2_L3_10, u2_L3_11, u2_L3_12, u2_L3_13, u2_L3_14, u2_L3_15, u2_L3_16, 
        u2_L3_17, u2_L3_18, u2_L3_19, u2_L3_2, u2_L3_20, u2_L3_21, u2_L3_22, u2_L3_23, u2_L3_24, 
        u2_L3_25, u2_L3_26, u2_L3_27, u2_L3_28, u2_L3_29, u2_L3_3, u2_L3_30, u2_L3_31, u2_L3_32, 
        u2_L3_4, u2_L3_5, u2_L3_6, u2_L3_7, u2_L3_8, u2_L3_9, u2_L4_1, u2_L4_10, u2_L4_11, 
        u2_L4_12, u2_L4_13, u2_L4_14, u2_L4_15, u2_L4_16, u2_L4_17, u2_L4_18, u2_L4_19, u2_L4_2, 
        u2_L4_20, u2_L4_21, u2_L4_22, u2_L4_23, u2_L4_24, u2_L4_25, u2_L4_26, u2_L4_27, u2_L4_28, 
        u2_L4_29, u2_L4_3, u2_L4_30, u2_L4_31, u2_L4_32, u2_L4_4, u2_L4_5, u2_L4_6, u2_L4_7, 
        u2_L4_8, u2_L4_9, u2_L5_1, u2_L5_10, u2_L5_11, u2_L5_12, u2_L5_13, u2_L5_14, u2_L5_15, 
        u2_L5_16, u2_L5_17, u2_L5_18, u2_L5_19, u2_L5_2, u2_L5_20, u2_L5_21, u2_L5_22, u2_L5_23, 
        u2_L5_24, u2_L5_25, u2_L5_26, u2_L5_27, u2_L5_28, u2_L5_29, u2_L5_3, u2_L5_30, u2_L5_31, 
        u2_L5_32, u2_L5_4, u2_L5_5, u2_L5_6, u2_L5_7, u2_L5_8, u2_L5_9, u2_L6_1, u2_L6_10, 
        u2_L6_11, u2_L6_12, u2_L6_13, u2_L6_14, u2_L6_15, u2_L6_16, u2_L6_17, u2_L6_18, u2_L6_19, 
        u2_L6_2, u2_L6_20, u2_L6_21, u2_L6_22, u2_L6_23, u2_L6_24, u2_L6_25, u2_L6_26, u2_L6_27, 
        u2_L6_28, u2_L6_29, u2_L6_3, u2_L6_30, u2_L6_31, u2_L6_32, u2_L6_4, u2_L6_5, u2_L6_6, 
        u2_L6_7, u2_L6_8, u2_L6_9, u2_L7_1, u2_L7_10, u2_L7_11, u2_L7_12, u2_L7_13, u2_L7_14, 
        u2_L7_15, u2_L7_16, u2_L7_17, u2_L7_18, u2_L7_19, u2_L7_2, u2_L7_20, u2_L7_21, u2_L7_22, 
        u2_L7_23, u2_L7_24, u2_L7_25, u2_L7_26, u2_L7_27, u2_L7_28, u2_L7_29, u2_L7_3, u2_L7_30, 
        u2_L7_31, u2_L7_32, u2_L7_4, u2_L7_5, u2_L7_6, u2_L7_7, u2_L7_8, u2_L7_9, u2_L8_1, 
        u2_L8_10, u2_L8_11, u2_L8_12, u2_L8_13, u2_L8_14, u2_L8_15, u2_L8_16, u2_L8_17, u2_L8_18, 
        u2_L8_19, u2_L8_2, u2_L8_20, u2_L8_21, u2_L8_22, u2_L8_23, u2_L8_24, u2_L8_25, u2_L8_26, 
        u2_L8_27, u2_L8_28, u2_L8_29, u2_L8_3, u2_L8_30, u2_L8_31, u2_L8_32, u2_L8_4, u2_L8_5, 
        u2_L8_6, u2_L8_7, u2_L8_8, u2_L8_9, u2_L9_1, u2_L9_10, u2_L9_11, u2_L9_12, u2_L9_13, 
        u2_L9_14, u2_L9_15, u2_L9_16, u2_L9_17, u2_L9_18, u2_L9_19, u2_L9_2, u2_L9_20, u2_L9_21, 
        u2_L9_22, u2_L9_23, u2_L9_24, u2_L9_25, u2_L9_26, u2_L9_27, u2_L9_28, u2_L9_29, u2_L9_3, 
        u2_L9_30, u2_L9_31, u2_L9_32, u2_L9_4, u2_L9_5, u2_L9_6, u2_L9_7, u2_L9_8, u2_L9_9, 
        u2_R0_1, u2_R0_10, u2_R0_11, u2_R0_12, u2_R0_13, u2_R0_14, u2_R0_15, u2_R0_16, u2_R0_17, 
        u2_R0_18, u2_R0_19, u2_R0_2, u2_R0_20, u2_R0_21, u2_R0_22, u2_R0_23, u2_R0_24, u2_R0_25, 
        u2_R0_26, u2_R0_27, u2_R0_28, u2_R0_29, u2_R0_3, u2_R0_30, u2_R0_31, u2_R0_32, u2_R0_4, 
        u2_R0_5, u2_R0_6, u2_R0_7, u2_R0_8, u2_R0_9, u2_R10_1, u2_R10_10, u2_R10_11, u2_R10_12, 
        u2_R10_13, u2_R10_14, u2_R10_15, u2_R10_16, u2_R10_17, u2_R10_18, u2_R10_19, u2_R10_2, u2_R10_20, 
        u2_R10_21, u2_R10_22, u2_R10_23, u2_R10_24, u2_R10_25, u2_R10_26, u2_R10_27, u2_R10_28, u2_R10_29, 
        u2_R10_3, u2_R10_30, u2_R10_31, u2_R10_32, u2_R10_4, u2_R10_5, u2_R10_6, u2_R10_7, u2_R10_8, 
        u2_R10_9, u2_R11_1, u2_R11_10, u2_R11_11, u2_R11_12, u2_R11_13, u2_R11_14, u2_R11_15, u2_R11_16, 
        u2_R11_17, u2_R11_18, u2_R11_19, u2_R11_2, u2_R11_20, u2_R11_21, u2_R11_22, u2_R11_23, u2_R11_24, 
        u2_R11_25, u2_R11_26, u2_R11_27, u2_R11_28, u2_R11_29, u2_R11_3, u2_R11_30, u2_R11_31, u2_R11_32, 
        u2_R11_4, u2_R11_5, u2_R11_6, u2_R11_7, u2_R11_8, u2_R11_9, u2_R12_1, u2_R12_10, u2_R12_11, 
        u2_R12_12, u2_R12_13, u2_R12_14, u2_R12_15, u2_R12_16, u2_R12_17, u2_R12_18, u2_R12_19, u2_R12_2, 
        u2_R12_20, u2_R12_21, u2_R12_22, u2_R12_23, u2_R12_24, u2_R12_25, u2_R12_26, u2_R12_27, u2_R12_28, 
        u2_R12_29, u2_R12_3, u2_R12_30, u2_R12_31, u2_R12_32, u2_R12_4, u2_R12_5, u2_R12_6, u2_R12_7, 
        u2_R12_8, u2_R12_9, u2_R13_1, u2_R13_10, u2_R13_11, u2_R13_12, u2_R13_13, u2_R13_14, u2_R13_15, 
        u2_R13_16, u2_R13_17, u2_R13_18, u2_R13_19, u2_R13_2, u2_R13_20, u2_R13_21, u2_R13_22, u2_R13_23, 
        u2_R13_24, u2_R13_25, u2_R13_26, u2_R13_27, u2_R13_28, u2_R13_29, u2_R13_3, u2_R13_30, u2_R13_31, 
        u2_R13_32, u2_R13_4, u2_R13_5, u2_R13_6, u2_R13_7, u2_R13_8, u2_R13_9, u2_R1_1, u2_R1_10, 
        u2_R1_11, u2_R1_12, u2_R1_13, u2_R1_14, u2_R1_15, u2_R1_16, u2_R1_17, u2_R1_18, u2_R1_19, 
        u2_R1_2, u2_R1_20, u2_R1_21, u2_R1_22, u2_R1_23, u2_R1_24, u2_R1_25, u2_R1_26, u2_R1_27, 
        u2_R1_28, u2_R1_29, u2_R1_3, u2_R1_30, u2_R1_31, u2_R1_32, u2_R1_4, u2_R1_5, u2_R1_6, 
        u2_R1_7, u2_R1_8, u2_R1_9, u2_R2_1, u2_R2_10, u2_R2_11, u2_R2_12, u2_R2_13, u2_R2_14, 
        u2_R2_15, u2_R2_16, u2_R2_17, u2_R2_18, u2_R2_19, u2_R2_2, u2_R2_20, u2_R2_21, u2_R2_22, 
        u2_R2_23, u2_R2_24, u2_R2_25, u2_R2_26, u2_R2_27, u2_R2_28, u2_R2_29, u2_R2_3, u2_R2_30, 
        u2_R2_31, u2_R2_32, u2_R2_4, u2_R2_5, u2_R2_6, u2_R2_7, u2_R2_8, u2_R2_9, u2_R3_1, 
        u2_R3_10, u2_R3_11, u2_R3_12, u2_R3_13, u2_R3_14, u2_R3_15, u2_R3_16, u2_R3_17, u2_R3_18, 
        u2_R3_19, u2_R3_2, u2_R3_20, u2_R3_21, u2_R3_22, u2_R3_23, u2_R3_24, u2_R3_25, u2_R3_26, 
        u2_R3_27, u2_R3_28, u2_R3_29, u2_R3_3, u2_R3_30, u2_R3_31, u2_R3_32, u2_R3_4, u2_R3_5, 
        u2_R3_6, u2_R3_7, u2_R3_8, u2_R3_9, u2_R4_1, u2_R4_10, u2_R4_11, u2_R4_12, u2_R4_13, 
        u2_R4_14, u2_R4_15, u2_R4_16, u2_R4_17, u2_R4_18, u2_R4_19, u2_R4_2, u2_R4_20, u2_R4_21, 
        u2_R4_22, u2_R4_23, u2_R4_24, u2_R4_25, u2_R4_26, u2_R4_27, u2_R4_28, u2_R4_29, u2_R4_3, 
        u2_R4_30, u2_R4_31, u2_R4_32, u2_R4_4, u2_R4_5, u2_R4_6, u2_R4_7, u2_R4_8, u2_R4_9, 
        u2_R5_1, u2_R5_10, u2_R5_11, u2_R5_12, u2_R5_13, u2_R5_14, u2_R5_15, u2_R5_16, u2_R5_17, 
        u2_R5_18, u2_R5_19, u2_R5_2, u2_R5_20, u2_R5_21, u2_R5_22, u2_R5_23, u2_R5_24, u2_R5_25, 
        u2_R5_26, u2_R5_27, u2_R5_28, u2_R5_29, u2_R5_3, u2_R5_30, u2_R5_31, u2_R5_32, u2_R5_4, 
        u2_R5_5, u2_R5_6, u2_R5_7, u2_R5_8, u2_R5_9, u2_R6_1, u2_R6_10, u2_R6_11, u2_R6_12, 
        u2_R6_13, u2_R6_14, u2_R6_15, u2_R6_16, u2_R6_17, u2_R6_18, u2_R6_19, u2_R6_2, u2_R6_20, 
        u2_R6_21, u2_R6_22, u2_R6_23, u2_R6_24, u2_R6_25, u2_R6_26, u2_R6_27, u2_R6_28, u2_R6_29, 
        u2_R6_3, u2_R6_30, u2_R6_31, u2_R6_32, u2_R6_4, u2_R6_5, u2_R6_6, u2_R6_7, u2_R6_8, 
        u2_R6_9, u2_R7_1, u2_R7_10, u2_R7_11, u2_R7_12, u2_R7_13, u2_R7_14, u2_R7_15, u2_R7_16, 
        u2_R7_17, u2_R7_18, u2_R7_19, u2_R7_2, u2_R7_20, u2_R7_21, u2_R7_22, u2_R7_23, u2_R7_24, 
        u2_R7_25, u2_R7_26, u2_R7_27, u2_R7_28, u2_R7_29, u2_R7_3, u2_R7_30, u2_R7_31, u2_R7_32, 
        u2_R7_4, u2_R7_5, u2_R7_6, u2_R7_7, u2_R7_8, u2_R7_9, u2_R8_1, u2_R8_10, u2_R8_11, 
        u2_R8_12, u2_R8_13, u2_R8_14, u2_R8_15, u2_R8_16, u2_R8_17, u2_R8_18, u2_R8_19, u2_R8_2, 
        u2_R8_20, u2_R8_21, u2_R8_22, u2_R8_23, u2_R8_24, u2_R8_25, u2_R8_26, u2_R8_27, u2_R8_28, 
        u2_R8_29, u2_R8_3, u2_R8_30, u2_R8_31, u2_R8_32, u2_R8_4, u2_R8_5, u2_R8_6, u2_R8_7, 
        u2_R8_8, u2_R8_9, u2_R9_1, u2_R9_10, u2_R9_11, u2_R9_12, u2_R9_13, u2_R9_14, u2_R9_15, 
        u2_R9_16, u2_R9_17, u2_R9_18, u2_R9_19, u2_R9_2, u2_R9_20, u2_R9_21, u2_R9_22, u2_R9_23, 
        u2_R9_24, u2_R9_25, u2_R9_26, u2_R9_27, u2_R9_28, u2_R9_29, u2_R9_3, u2_R9_30, u2_R9_31, 
        u2_R9_32, u2_R9_4, u2_R9_5, u2_R9_6, u2_R9_7, u2_R9_8, u2_R9_9, u2_desIn_r_0, u2_desIn_r_1, 
        u2_desIn_r_10, u2_desIn_r_11, u2_desIn_r_12, u2_desIn_r_13, u2_desIn_r_14, u2_desIn_r_15, u2_desIn_r_16, u2_desIn_r_17, u2_desIn_r_18, 
        u2_desIn_r_19, u2_desIn_r_2, u2_desIn_r_20, u2_desIn_r_21, u2_desIn_r_22, u2_desIn_r_23, u2_desIn_r_24, u2_desIn_r_25, u2_desIn_r_26, 
        u2_desIn_r_27, u2_desIn_r_28, u2_desIn_r_29, u2_desIn_r_3, u2_desIn_r_30, u2_desIn_r_31, u2_desIn_r_32, u2_desIn_r_33, u2_desIn_r_34, 
        u2_desIn_r_35, u2_desIn_r_36, u2_desIn_r_37, u2_desIn_r_38, u2_desIn_r_39, u2_desIn_r_4, u2_desIn_r_40, u2_desIn_r_41, u2_desIn_r_42, 
        u2_desIn_r_43, u2_desIn_r_44, u2_desIn_r_45, u2_desIn_r_46, u2_desIn_r_47, u2_desIn_r_48, u2_desIn_r_49, u2_desIn_r_5, u2_desIn_r_50, 
        u2_desIn_r_51, u2_desIn_r_52, u2_desIn_r_53, u2_desIn_r_54, u2_desIn_r_55, u2_desIn_r_56, u2_desIn_r_57, u2_desIn_r_58, u2_desIn_r_59, 
        u2_desIn_r_6, u2_desIn_r_60, u2_desIn_r_61, u2_desIn_r_62, u2_desIn_r_63, u2_desIn_r_7, u2_desIn_r_8, u2_desIn_r_9, u2_key_r_0, 
        u2_key_r_1, u2_key_r_10, u2_key_r_11, u2_key_r_12, u2_key_r_13, u2_key_r_14, u2_key_r_16, u2_key_r_17, u2_key_r_19, 
        u2_key_r_2, u2_key_r_20, u2_key_r_21, u2_key_r_22, u2_key_r_23, u2_key_r_24, u2_key_r_25, u2_key_r_26, u2_key_r_27, 
        u2_key_r_28, u2_key_r_29, u2_key_r_3, u2_key_r_30, u2_key_r_31, u2_key_r_32, u2_key_r_33, u2_key_r_34, u2_key_r_35, 
        u2_key_r_36, u2_key_r_37, u2_key_r_4, u2_key_r_40, u2_key_r_41, u2_key_r_42, u2_key_r_43, u2_key_r_44, u2_key_r_46, 
        u2_key_r_47, u2_key_r_48, u2_key_r_49, u2_key_r_50, u2_key_r_51, u2_key_r_52, u2_key_r_53, u2_key_r_54, u2_key_r_55, 
        u2_key_r_6, u2_key_r_7, u2_key_r_8, u2_key_r_9, u2_uk_K_r0_11, u2_uk_K_r0_13, u2_uk_K_r0_15, u2_uk_K_r0_17, u2_uk_K_r0_25, 
        u2_uk_K_r0_31, u2_uk_K_r0_32, u2_uk_K_r0_34, u2_uk_K_r0_36, u2_uk_K_r0_47, u2_uk_K_r0_49, u2_uk_K_r0_55, u2_uk_K_r10_10, u2_uk_K_r10_16, 
        u2_uk_K_r10_25, u2_uk_K_r10_27, u2_uk_K_r10_32, u2_uk_K_r10_34, u2_uk_K_r10_4, u2_uk_K_r10_41, u2_uk_K_r10_43, u2_uk_K_r10_44, u2_uk_K_r10_49, 
        u2_uk_K_r11_10, u2_uk_K_r11_11, u2_uk_K_r11_19, u2_uk_K_r11_20, u2_uk_K_r11_21, u2_uk_K_r11_24, u2_uk_K_r11_25, u2_uk_K_r11_26, u2_uk_K_r11_27, 
        u2_uk_K_r11_28, u2_uk_K_r11_29, u2_uk_K_r11_33, u2_uk_K_r11_39, u2_uk_K_r11_4, u2_uk_K_r11_47, u2_uk_K_r11_48, u2_uk_K_r11_53, u2_uk_K_r11_6, 
        u2_uk_K_r11_7, u2_uk_K_r12_1, u2_uk_K_r12_10, u2_uk_K_r12_15, u2_uk_K_r12_16, u2_uk_K_r12_25, u2_uk_K_r12_30, u2_uk_K_r12_33, u2_uk_K_r12_36, 
        u2_uk_K_r12_41, u2_uk_K_r12_42, u2_uk_K_r12_7, u2_uk_K_r13_0, u2_uk_K_r13_13, u2_uk_K_r13_17, u2_uk_K_r13_19, u2_uk_K_r13_22, u2_uk_K_r13_25, 
        u2_uk_K_r13_32, u2_uk_K_r13_38, u2_uk_K_r13_55, u2_uk_K_r14_10, u2_uk_K_r14_12, u2_uk_K_r14_15, u2_uk_K_r14_16, u2_uk_K_r14_18, u2_uk_K_r14_2, 
        u2_uk_K_r14_3, u2_uk_K_r14_45, u2_uk_K_r14_46, u2_uk_K_r14_5, u2_uk_K_r14_50, u2_uk_K_r14_9, u2_uk_K_r1_15, u2_uk_K_r1_16, u2_uk_K_r1_17, 
        u2_uk_K_r1_18, u2_uk_K_r1_21, u2_uk_K_r1_22, u2_uk_K_r1_41, u2_uk_K_r1_42, u2_uk_K_r1_44, u2_uk_K_r1_47, u2_uk_K_r1_7, u2_uk_K_r2_13, 
        u2_uk_K_r2_18, u2_uk_K_r2_21, u2_uk_K_r2_24, u2_uk_K_r2_25, u2_uk_K_r2_26, u2_uk_K_r2_27, u2_uk_K_r2_28, u2_uk_K_r2_31, u2_uk_K_r2_36, 
        u2_uk_K_r2_49, u2_uk_K_r2_50, u2_uk_K_r2_55, u2_uk_K_r2_6, u2_uk_K_r3_10, u2_uk_K_r3_11, u2_uk_K_r3_14, u2_uk_K_r3_15, u2_uk_K_r3_16, 
        u2_uk_K_r3_19, u2_uk_K_r3_29, u2_uk_K_r3_38, u2_uk_K_r3_4, u2_uk_K_r3_43, u2_uk_K_r3_52, u2_uk_K_r3_9, u2_uk_K_r4_0, u2_uk_K_r4_11, 
        u2_uk_K_r4_17, u2_uk_K_r4_3, u2_uk_K_r4_33, u2_uk_K_r4_35, u2_uk_K_r4_38, u2_uk_K_r4_4, u2_uk_K_r4_41, u2_uk_K_r4_47, u2_uk_K_r4_5, 
        u2_uk_K_r4_54, u2_uk_K_r4_55, u2_uk_K_r5_0, u2_uk_K_r5_1, u2_uk_K_r5_10, u2_uk_K_r5_16, u2_uk_K_r5_17, u2_uk_K_r5_18, u2_uk_K_r5_19, 
        u2_uk_K_r5_21, u2_uk_K_r5_23, u2_uk_K_r5_26, u2_uk_K_r5_31, u2_uk_K_r5_37, u2_uk_K_r5_39, u2_uk_K_r5_4, u2_uk_K_r5_40, u2_uk_K_r5_41, 
        u2_uk_K_r5_43, u2_uk_K_r5_48, u2_uk_K_r5_51, u2_uk_K_r5_7, u2_uk_K_r6_0, u2_uk_K_r6_10, u2_uk_K_r6_14, u2_uk_K_r6_26, u2_uk_K_r6_29, 
        u2_uk_K_r6_3, u2_uk_K_r6_31, u2_uk_K_r6_34, u2_uk_K_r6_37, u2_uk_K_r6_46, u2_uk_K_r6_51, u2_uk_K_r6_53, u2_uk_K_r6_7, u2_uk_K_r7_0, 
        u2_uk_K_r7_13, u2_uk_K_r7_16, u2_uk_K_r7_2, u2_uk_K_r7_20, u2_uk_K_r7_23, u2_uk_K_r7_25, u2_uk_K_r7_26, u2_uk_K_r7_31, u2_uk_K_r7_32, 
        u2_uk_K_r7_37, u2_uk_K_r7_39, u2_uk_K_r7_41, u2_uk_K_r7_46, u2_uk_K_r7_48, u2_uk_K_r7_55, u2_uk_K_r7_9, u2_uk_K_r8_13, u2_uk_K_r8_16, 
        u2_uk_K_r8_17, u2_uk_K_r8_19, u2_uk_K_r8_2, u2_uk_K_r8_21, u2_uk_K_r8_22, u2_uk_K_r8_27, u2_uk_K_r8_28, u2_uk_K_r8_32, u2_uk_K_r8_37, 
        u2_uk_K_r8_40, u2_uk_K_r8_41, u2_uk_K_r8_42, u2_uk_K_r8_43, u2_uk_K_r8_44, u2_uk_K_r8_48, u2_uk_K_r8_52, u2_uk_K_r8_8, u2_uk_K_r9_0, 
        u2_uk_K_r9_1, u2_uk_K_r9_10, u2_uk_K_r9_12, u2_uk_K_r9_13, u2_uk_K_r9_15, u2_uk_K_r9_18, u2_uk_K_r9_19, u2_uk_K_r9_23, u2_uk_K_r9_25, 
        u2_uk_K_r9_27, u2_uk_K_r9_31, u2_uk_K_r9_33, u2_uk_K_r9_4, u2_uk_K_r9_45, u2_uk_K_r9_48, u2_uk_K_r9_49, u2_uk_K_r9_5, u2_uk_K_r9_54, 
        u2_uk_K_r9_55, u2_uk_K_r9_9, u2_uk_n1001, u2_uk_n1007, u2_uk_n1011, u2_uk_n1018, u2_uk_n1022, u2_uk_n1024, u2_uk_n1027, 
        u2_uk_n1028, u2_uk_n1031, u2_uk_n1035, u2_uk_n1036, u2_uk_n1038, u2_uk_n1040, u2_uk_n1042, u2_uk_n1043, u2_uk_n1044, 
        u2_uk_n1046, u2_uk_n1049, u2_uk_n1061, u2_uk_n1063, u2_uk_n1069, u2_uk_n1070, u2_uk_n1073, u2_uk_n1074, u2_uk_n1077, 
        u2_uk_n1079, u2_uk_n1081, u2_uk_n1082, u2_uk_n1089, u2_uk_n1093, u2_uk_n1094, u2_uk_n1096, u2_uk_n1097, u2_uk_n1100, 
        u2_uk_n1104, u2_uk_n1105, u2_uk_n1107, u2_uk_n1112, u2_uk_n1113, u2_uk_n1116, u2_uk_n1119, u2_uk_n1120, u2_uk_n1121, 
        u2_uk_n1125, u2_uk_n1128, u2_uk_n1130, u2_uk_n1131, u2_uk_n1132, u2_uk_n1134, u2_uk_n1136, u2_uk_n1137, u2_uk_n1140, 
        u2_uk_n1141, u2_uk_n1188, u2_uk_n1189, u2_uk_n1190, u2_uk_n1194, u2_uk_n1195, u2_uk_n1197, u2_uk_n1198, u2_uk_n1199, 
        u2_uk_n1200, u2_uk_n1201, u2_uk_n1203, u2_uk_n1204, u2_uk_n1205, u2_uk_n1206, u2_uk_n1207, u2_uk_n1208, u2_uk_n1209, 
        u2_uk_n1210, u2_uk_n1212, u2_uk_n1213, u2_uk_n1214, u2_uk_n1215, u2_uk_n1216, u2_uk_n1217, u2_uk_n1218, u2_uk_n1219, 
        u2_uk_n1220, u2_uk_n1221, u2_uk_n1222, u2_uk_n1223, u2_uk_n1225, u2_uk_n1226, u2_uk_n1227, u2_uk_n1228, u2_uk_n1229, 
        u2_uk_n1230, u2_uk_n1231, u2_uk_n1232, u2_uk_n1233, u2_uk_n1234, u2_uk_n1236, u2_uk_n1237, u2_uk_n1238, u2_uk_n1239, 
        u2_uk_n1240, u2_uk_n1243, u2_uk_n1244, u2_uk_n1245, u2_uk_n1246, u2_uk_n1247, u2_uk_n1248, u2_uk_n1249, u2_uk_n1251, 
        u2_uk_n1252, u2_uk_n1254, u2_uk_n1258, u2_uk_n1259, u2_uk_n1260, u2_uk_n1261, u2_uk_n1264, u2_uk_n1265, u2_uk_n1266, 
        u2_uk_n1267, u2_uk_n1269, u2_uk_n1270, u2_uk_n1274, u2_uk_n1275, u2_uk_n1279, u2_uk_n1280, u2_uk_n1281, u2_uk_n1282, 
        u2_uk_n1283, u2_uk_n1284, u2_uk_n1285, u2_uk_n1286, u2_uk_n1287, u2_uk_n1288, u2_uk_n1290, u2_uk_n1291, u2_uk_n1292, 
        u2_uk_n1293, u2_uk_n1294, u2_uk_n1295, u2_uk_n1296, u2_uk_n1297, u2_uk_n1298, u2_uk_n1299, u2_uk_n1300, u2_uk_n1301, 
        u2_uk_n1302, u2_uk_n1303, u2_uk_n1305, u2_uk_n1306, u2_uk_n1308, u2_uk_n1309, u2_uk_n1310, u2_uk_n1311, u2_uk_n1312, 
        u2_uk_n1313, u2_uk_n1314, u2_uk_n1315, u2_uk_n1316, u2_uk_n1317, u2_uk_n1318, u2_uk_n1319, u2_uk_n1320, u2_uk_n1321, 
        u2_uk_n1322, u2_uk_n1323, u2_uk_n1324, u2_uk_n1325, u2_uk_n1326, u2_uk_n1328, u2_uk_n1329, u2_uk_n1330, u2_uk_n1331, 
        u2_uk_n1333, u2_uk_n1335, u2_uk_n1336, u2_uk_n1337, u2_uk_n1339, u2_uk_n1341, u2_uk_n1342, u2_uk_n1344, u2_uk_n1345, 
        u2_uk_n1346, u2_uk_n1347, u2_uk_n1348, u2_uk_n1350, u2_uk_n1351, u2_uk_n1352, u2_uk_n1353, u2_uk_n1356, u2_uk_n1359, 
        u2_uk_n1360, u2_uk_n1361, u2_uk_n1363, u2_uk_n1364, u2_uk_n1365, u2_uk_n1367, u2_uk_n1370, u2_uk_n1372, u2_uk_n1375, 
        u2_uk_n1376, u2_uk_n1377, u2_uk_n1378, u2_uk_n1379, u2_uk_n1381, u2_uk_n1382, u2_uk_n1383, u2_uk_n1395, u2_uk_n1396, 
        u2_uk_n1400, u2_uk_n1401, u2_uk_n1403, u2_uk_n1405, u2_uk_n1408, u2_uk_n1410, u2_uk_n1411, u2_uk_n1412, u2_uk_n1413, 
        u2_uk_n1414, u2_uk_n1416, u2_uk_n1418, u2_uk_n1419, u2_uk_n1420, u2_uk_n1422, u2_uk_n1424, u2_uk_n1425, u2_uk_n1426, 
        u2_uk_n1428, u2_uk_n1429, u2_uk_n1430, u2_uk_n1433, u2_uk_n1435, u2_uk_n1438, u2_uk_n1439, u2_uk_n1440, u2_uk_n1441, 
        u2_uk_n1442, u2_uk_n1444, u2_uk_n1445, u2_uk_n1446, u2_uk_n1447, u2_uk_n1448, u2_uk_n1452, u2_uk_n1453, u2_uk_n1454, 
        u2_uk_n1456, u2_uk_n1457, u2_uk_n1458, u2_uk_n1459, u2_uk_n1460, u2_uk_n1461, u2_uk_n1462, u2_uk_n1464, u2_uk_n1465, 
        u2_uk_n1466, u2_uk_n1468, u2_uk_n1470, u2_uk_n1471, u2_uk_n1475, u2_uk_n1480, u2_uk_n1486, u2_uk_n1487, u2_uk_n1488, 
        u2_uk_n1490, u2_uk_n1491, u2_uk_n1493, u2_uk_n1494, u2_uk_n1496, u2_uk_n1497, u2_uk_n1498, u2_uk_n1499, u2_uk_n1500, 
        u2_uk_n1501, u2_uk_n1502, u2_uk_n1503, u2_uk_n1504, u2_uk_n1506, u2_uk_n1507, u2_uk_n1508, u2_uk_n1510, u2_uk_n1511, 
        u2_uk_n1513, u2_uk_n1514, u2_uk_n1515, u2_uk_n1517, u2_uk_n1518, u2_uk_n1519, u2_uk_n1521, u2_uk_n1522, u2_uk_n1524, 
        u2_uk_n1525, u2_uk_n1526, u2_uk_n1527, u2_uk_n1528, u2_uk_n1529, u2_uk_n1530, u2_uk_n1531, u2_uk_n1532, u2_uk_n1533, 
        u2_uk_n1535, u2_uk_n1536, u2_uk_n1537, u2_uk_n1538, u2_uk_n1542, u2_uk_n1543, u2_uk_n1544, u2_uk_n1548, u2_uk_n1549, 
        u2_uk_n1551, u2_uk_n1555, u2_uk_n1556, u2_uk_n1558, u2_uk_n1563, u2_uk_n1565, u2_uk_n1568, u2_uk_n1570, u2_uk_n1571, 
        u2_uk_n1573, u2_uk_n1574, u2_uk_n1576, u2_uk_n1577, u2_uk_n1580, u2_uk_n1583, u2_uk_n1585, u2_uk_n1586, u2_uk_n1590, 
        u2_uk_n1591, u2_uk_n1592, u2_uk_n1594, u2_uk_n1595, u2_uk_n1597, u2_uk_n1598, u2_uk_n1599, u2_uk_n1600, u2_uk_n1602, 
        u2_uk_n1603, u2_uk_n1604, u2_uk_n1605, u2_uk_n1609, u2_uk_n1610, u2_uk_n1612, u2_uk_n1613, u2_uk_n1614, u2_uk_n1615, 
        u2_uk_n1617, u2_uk_n1622, u2_uk_n1623, u2_uk_n1624, u2_uk_n1625, u2_uk_n1626, u2_uk_n1629, u2_uk_n1630, u2_uk_n1631, 
        u2_uk_n1632, u2_uk_n1633, u2_uk_n1634, u2_uk_n1639, u2_uk_n1640, u2_uk_n1642, u2_uk_n1643, u2_uk_n1646, u2_uk_n1647, 
        u2_uk_n1652, u2_uk_n1653, u2_uk_n1654, u2_uk_n1657, u2_uk_n1658, u2_uk_n1659, u2_uk_n1660, u2_uk_n1661, u2_uk_n1664, 
        u2_uk_n1665, u2_uk_n1666, u2_uk_n1668, u2_uk_n1672, u2_uk_n1673, u2_uk_n1674, u2_uk_n1675, u2_uk_n1677, u2_uk_n1678, 
        u2_uk_n1680, u2_uk_n1681, u2_uk_n1682, u2_uk_n1683, u2_uk_n1684, u2_uk_n1685, u2_uk_n1687, u2_uk_n1688, u2_uk_n1689, 
        u2_uk_n1690, u2_uk_n1691, u2_uk_n1693, u2_uk_n1698, u2_uk_n1699, u2_uk_n1700, u2_uk_n1702, u2_uk_n1705, u2_uk_n1707, 
        u2_uk_n1708, u2_uk_n1709, u2_uk_n1715, u2_uk_n1718, u2_uk_n1720, u2_uk_n1721, u2_uk_n1722, u2_uk_n1723, u2_uk_n1724, 
        u2_uk_n1725, u2_uk_n1726, u2_uk_n1727, u2_uk_n1728, u2_uk_n1731, u2_uk_n1732, u2_uk_n1734, u2_uk_n1735, u2_uk_n1736, 
        u2_uk_n1737, u2_uk_n1738, u2_uk_n1742, u2_uk_n1743, u2_uk_n1744, u2_uk_n1745, u2_uk_n1746, u2_uk_n1747, u2_uk_n1750, 
        u2_uk_n1753, u2_uk_n1755, u2_uk_n1760, u2_uk_n1761, u2_uk_n1762, u2_uk_n1763, u2_uk_n1767, u2_uk_n1768, u2_uk_n1769, 
        u2_uk_n1770, u2_uk_n1772, u2_uk_n1773, u2_uk_n1776, u2_uk_n1777, u2_uk_n1778, u2_uk_n1779, u2_uk_n1781, u2_uk_n1782, 
        u2_uk_n1783, u2_uk_n1785, u2_uk_n1786, u2_uk_n1788, u2_uk_n1789, u2_uk_n1790, u2_uk_n1791, u2_uk_n1792, u2_uk_n1793, 
        u2_uk_n1794, u2_uk_n1796, u2_uk_n1797, u2_uk_n1799, u2_uk_n1800, u2_uk_n1801, u2_uk_n1802, u2_uk_n1803, u2_uk_n1805, 
        u2_uk_n1806, u2_uk_n1807, u2_uk_n1808, u2_uk_n1809, u2_uk_n1810, u2_uk_n1811, u2_uk_n1814, u2_uk_n1815, u2_uk_n1816, 
        u2_uk_n1817, u2_uk_n1818, u2_uk_n1819, u2_uk_n1820, u2_uk_n1821, u2_uk_n1822, u2_uk_n1823, u2_uk_n1824, u2_uk_n1825, 
        u2_uk_n1826, u2_uk_n1828, u2_uk_n1832, u2_uk_n1833, u2_uk_n1834, u2_uk_n1835, u2_uk_n1836, u2_uk_n1837, u2_uk_n1838, 
        u2_uk_n1839, u2_uk_n1840, u2_uk_n1842, u2_uk_n1843, u2_uk_n1845, u2_uk_n1846, u2_uk_n1849, u2_uk_n1850, u2_uk_n1851, 
        u2_uk_n1852, u2_uk_n1853, u2_uk_n1854, u2_uk_n1855, u2_uk_n1856, u2_uk_n238, u2_uk_n240, u2_uk_n251, u2_uk_n257, 
        u2_uk_n299, u2_uk_n313, u2_uk_n319, u2_uk_n363, u2_uk_n373, u2_uk_n376, u2_uk_n377, u2_uk_n379, u2_uk_n385, 
        u2_uk_n408, u2_uk_n415, u2_uk_n421, u2_uk_n443, u2_uk_n456, u2_uk_n467, u2_uk_n468, u2_uk_n472, u2_uk_n500, 
        u2_uk_n503, u2_uk_n504, u2_uk_n520, u2_uk_n526, u2_uk_n551, u2_uk_n586, u2_uk_n608, u2_uk_n665, u2_uk_n677, 
        u2_uk_n682, u2_uk_n689, u2_uk_n702, u2_uk_n931, u2_uk_n933, u2_uk_n939, u2_uk_n941, u2_uk_n942, u2_uk_n943, 
        u2_uk_n944, u2_uk_n945, u2_uk_n947, u2_uk_n948, u2_uk_n954, u2_uk_n955, u2_uk_n956, u2_uk_n961, u2_uk_n967, 
        u2_uk_n970, u2_uk_n972, u2_uk_n979, u2_uk_n984, u2_uk_n986, u2_uk_n994, u2_uk_n996, u2_uk_n997 );
  input clk;
  input decrypt;
  input [63:0] desIn;
  input [55:0] key1;
  input [55:0] key2;
  input [55:0] key3;
  output [63:0] desOut;
  input u0_FP_1, u0_FP_10, u0_FP_11, u0_FP_12, u0_FP_13, u0_FP_14, u0_FP_15, u0_FP_16, u0_FP_17, 
        u0_FP_18, u0_FP_19, u0_FP_2, u0_FP_20, u0_FP_21, u0_FP_22, u0_FP_23, u0_FP_24, u0_FP_25, 
        u0_FP_26, u0_FP_27, u0_FP_28, u0_FP_29, u0_FP_3, u0_FP_30, u0_FP_31, u0_FP_32, u0_FP_4, 
        u0_FP_5, u0_FP_6, u0_FP_7, u0_FP_8, u0_FP_9, u0_N0, u0_N1, u0_N10, u0_N100, 
        u0_N101, u0_N102, u0_N103, u0_N104, u0_N105, u0_N106, u0_N107, u0_N108, u0_N109, 
        u0_N11, u0_N110, u0_N111, u0_N112, u0_N113, u0_N114, u0_N115, u0_N116, u0_N117, 
        u0_N118, u0_N119, u0_N12, u0_N120, u0_N121, u0_N122, u0_N123, u0_N124, u0_N125, 
        u0_N126, u0_N127, u0_N128, u0_N129, u0_N13, u0_N130, u0_N131, u0_N132, u0_N133, 
        u0_N134, u0_N135, u0_N136, u0_N137, u0_N138, u0_N139, u0_N14, u0_N140, u0_N141, 
        u0_N142, u0_N143, u0_N144, u0_N145, u0_N146, u0_N147, u0_N148, u0_N149, u0_N15, 
        u0_N150, u0_N151, u0_N152, u0_N153, u0_N154, u0_N155, u0_N156, u0_N157, u0_N158, 
        u0_N159, u0_N16, u0_N160, u0_N161, u0_N162, u0_N163, u0_N164, u0_N165, u0_N166, 
        u0_N167, u0_N168, u0_N169, u0_N17, u0_N170, u0_N171, u0_N172, u0_N173, u0_N174, 
        u0_N175, u0_N176, u0_N177, u0_N178, u0_N179, u0_N18, u0_N180, u0_N181, u0_N182, 
        u0_N183, u0_N184, u0_N185, u0_N186, u0_N187, u0_N188, u0_N189, u0_N19, u0_N190, 
        u0_N191, u0_N192, u0_N193, u0_N194, u0_N195, u0_N196, u0_N197, u0_N198, u0_N199, 
        u0_N2, u0_N20, u0_N200, u0_N201, u0_N202, u0_N203, u0_N204, u0_N205, u0_N206, 
        u0_N207, u0_N208, u0_N209, u0_N21, u0_N210, u0_N211, u0_N212, u0_N213, u0_N214, 
        u0_N215, u0_N216, u0_N217, u0_N218, u0_N219, u0_N22, u0_N220, u0_N221, u0_N222, 
        u0_N223, u0_N224, u0_N225, u0_N226, u0_N227, u0_N228, u0_N229, u0_N23, u0_N230, 
        u0_N231, u0_N232, u0_N233, u0_N234, u0_N235, u0_N236, u0_N237, u0_N238, u0_N239, 
        u0_N24, u0_N240, u0_N241, u0_N242, u0_N243, u0_N244, u0_N245, u0_N246, u0_N247, 
        u0_N248, u0_N249, u0_N25, u0_N250, u0_N251, u0_N252, u0_N253, u0_N254, u0_N255, 
        u0_N256, u0_N257, u0_N258, u0_N259, u0_N26, u0_N260, u0_N261, u0_N262, u0_N263, 
        u0_N264, u0_N265, u0_N266, u0_N267, u0_N268, u0_N269, u0_N27, u0_N270, u0_N271, 
        u0_N272, u0_N273, u0_N274, u0_N275, u0_N276, u0_N277, u0_N278, u0_N279, u0_N28, 
        u0_N280, u0_N281, u0_N282, u0_N283, u0_N284, u0_N285, u0_N286, u0_N287, u0_N288, 
        u0_N289, u0_N29, u0_N290, u0_N291, u0_N292, u0_N293, u0_N294, u0_N295, u0_N296, 
        u0_N297, u0_N298, u0_N299, u0_N3, u0_N30, u0_N300, u0_N301, u0_N302, u0_N303, 
        u0_N304, u0_N305, u0_N306, u0_N307, u0_N308, u0_N309, u0_N31, u0_N310, u0_N311, 
        u0_N312, u0_N313, u0_N314, u0_N315, u0_N316, u0_N317, u0_N318, u0_N319, u0_N32, 
        u0_N320, u0_N321, u0_N322, u0_N323, u0_N324, u0_N325, u0_N326, u0_N327, u0_N328, 
        u0_N329, u0_N33, u0_N330, u0_N331, u0_N332, u0_N333, u0_N334, u0_N335, u0_N336, 
        u0_N337, u0_N338, u0_N339, u0_N34, u0_N340, u0_N341, u0_N342, u0_N343, u0_N344, 
        u0_N345, u0_N346, u0_N347, u0_N348, u0_N349, u0_N35, u0_N350, u0_N351, u0_N352, 
        u0_N353, u0_N354, u0_N355, u0_N356, u0_N357, u0_N358, u0_N359, u0_N36, u0_N360, 
        u0_N361, u0_N362, u0_N363, u0_N364, u0_N365, u0_N366, u0_N367, u0_N368, u0_N369, 
        u0_N37, u0_N370, u0_N371, u0_N372, u0_N373, u0_N374, u0_N375, u0_N376, u0_N377, 
        u0_N378, u0_N379, u0_N38, u0_N380, u0_N381, u0_N382, u0_N383, u0_N384, u0_N385, 
        u0_N386, u0_N387, u0_N388, u0_N389, u0_N39, u0_N390, u0_N391, u0_N392, u0_N393, 
        u0_N394, u0_N395, u0_N396, u0_N397, u0_N398, u0_N399, u0_N4, u0_N40, u0_N400, 
        u0_N401, u0_N402, u0_N403, u0_N404, u0_N405, u0_N406, u0_N407, u0_N408, u0_N409, 
        u0_N41, u0_N410, u0_N411, u0_N412, u0_N413, u0_N414, u0_N415, u0_N416, u0_N417, 
        u0_N418, u0_N419, u0_N42, u0_N420, u0_N421, u0_N422, u0_N423, u0_N424, u0_N425, 
        u0_N426, u0_N427, u0_N428, u0_N429, u0_N43, u0_N430, u0_N431, u0_N432, u0_N433, 
        u0_N434, u0_N435, u0_N436, u0_N437, u0_N438, u0_N439, u0_N44, u0_N440, u0_N441, 
        u0_N442, u0_N443, u0_N444, u0_N445, u0_N446, u0_N447, u0_N448, u0_N449, u0_N45, 
        u0_N450, u0_N451, u0_N452, u0_N453, u0_N454, u0_N455, u0_N456, u0_N457, u0_N458, 
        u0_N459, u0_N46, u0_N460, u0_N461, u0_N462, u0_N463, u0_N464, u0_N465, u0_N466, 
        u0_N467, u0_N468, u0_N469, u0_N47, u0_N470, u0_N471, u0_N472, u0_N473, u0_N474, 
        u0_N475, u0_N476, u0_N477, u0_N478, u0_N479, u0_N48, u0_N49, u0_N5, u0_N50, 
        u0_N51, u0_N52, u0_N53, u0_N54, u0_N55, u0_N56, u0_N57, u0_N58, u0_N59, 
        u0_N6, u0_N60, u0_N61, u0_N62, u0_N63, u0_N64, u0_N65, u0_N66, u0_N67, 
        u0_N68, u0_N69, u0_N7, u0_N70, u0_N71, u0_N72, u0_N73, u0_N74, u0_N75, 
        u0_N76, u0_N77, u0_N78, u0_N79, u0_N8, u0_N80, u0_N81, u0_N82, u0_N83, 
        u0_N84, u0_N85, u0_N86, u0_N87, u0_N88, u0_N89, u0_N9, u0_N90, u0_N91, 
        u0_N92, u0_N93, u0_N94, u0_N95, u0_N96, u0_N97, u0_N98, u0_N99, u0_uk_n1010, 
        u0_uk_n1016, u0_uk_n147, u0_uk_n148, u0_uk_n155, u0_uk_n161, u0_uk_n162, u0_uk_n163, u0_uk_n164, u0_uk_n182, 
        u0_uk_n187, u0_uk_n188, u0_uk_n191, u0_uk_n202, u0_uk_n203, u0_uk_n207, u0_uk_n208, u0_uk_n209, u0_uk_n213, 
        u0_uk_n214, u0_uk_n217, u0_uk_n220, u0_uk_n222, u0_uk_n223, u0_uk_n230, u0_uk_n231, u0_uk_n238, u0_uk_n240, 
        u0_uk_n242, u0_uk_n250, u0_uk_n251, u0_uk_n252, u0_uk_n674, u0_uk_n675, u0_uk_n680, u0_uk_n684, u0_uk_n687, 
        u0_uk_n690, u0_uk_n691, u0_uk_n696, u0_uk_n697, u0_uk_n698, u0_uk_n705, u0_uk_n707, u0_uk_n711, u0_uk_n715, 
        u0_uk_n756, u0_uk_n762, u0_uk_n773, u0_uk_n777, u0_uk_n778, u0_uk_n790, u0_uk_n798, u0_uk_n804, u0_uk_n823, 
        u0_uk_n841, u0_uk_n848, u0_uk_n856, u0_uk_n863, u0_uk_n867, u0_uk_n871, u0_uk_n880, u0_uk_n888, u0_uk_n889, 
        u0_uk_n890, u0_uk_n894, u0_uk_n906, u0_uk_n926, u0_uk_n936, u0_uk_n942, u0_uk_n945, u0_uk_n961, u0_uk_n969, 
        u0_uk_n989, u0_uk_n998, u1_FP_1, u1_FP_10, u1_FP_11, u1_FP_12, u1_FP_13, u1_FP_14, u1_FP_15, 
        u1_FP_16, u1_FP_17, u1_FP_18, u1_FP_19, u1_FP_2, u1_FP_20, u1_FP_21, u1_FP_22, u1_FP_23, 
        u1_FP_24, u1_FP_25, u1_FP_26, u1_FP_27, u1_FP_28, u1_FP_29, u1_FP_3, u1_FP_30, u1_FP_31, 
        u1_FP_32, u1_FP_4, u1_FP_5, u1_FP_6, u1_FP_7, u1_FP_8, u1_FP_9, u1_N0, u1_N1, 
        u1_N10, u1_N100, u1_N101, u1_N102, u1_N103, u1_N104, u1_N105, u1_N106, u1_N107, 
        u1_N108, u1_N109, u1_N11, u1_N110, u1_N111, u1_N112, u1_N113, u1_N114, u1_N115, 
        u1_N116, u1_N117, u1_N118, u1_N119, u1_N12, u1_N120, u1_N121, u1_N122, u1_N123, 
        u1_N124, u1_N125, u1_N126, u1_N127, u1_N128, u1_N129, u1_N13, u1_N130, u1_N131, 
        u1_N132, u1_N133, u1_N134, u1_N135, u1_N136, u1_N137, u1_N138, u1_N139, u1_N14, 
        u1_N140, u1_N141, u1_N142, u1_N143, u1_N144, u1_N145, u1_N146, u1_N147, u1_N148, 
        u1_N149, u1_N15, u1_N150, u1_N151, u1_N152, u1_N153, u1_N154, u1_N155, u1_N156, 
        u1_N157, u1_N158, u1_N159, u1_N16, u1_N160, u1_N161, u1_N162, u1_N163, u1_N164, 
        u1_N165, u1_N166, u1_N167, u1_N168, u1_N169, u1_N17, u1_N170, u1_N171, u1_N172, 
        u1_N173, u1_N174, u1_N175, u1_N176, u1_N177, u1_N178, u1_N179, u1_N18, u1_N180, 
        u1_N181, u1_N182, u1_N183, u1_N184, u1_N185, u1_N186, u1_N187, u1_N188, u1_N189, 
        u1_N19, u1_N190, u1_N191, u1_N192, u1_N193, u1_N194, u1_N195, u1_N196, u1_N197, 
        u1_N198, u1_N199, u1_N2, u1_N20, u1_N200, u1_N201, u1_N202, u1_N203, u1_N204, 
        u1_N205, u1_N206, u1_N207, u1_N208, u1_N209, u1_N21, u1_N210, u1_N211, u1_N212, 
        u1_N213, u1_N214, u1_N215, u1_N216, u1_N217, u1_N218, u1_N219, u1_N22, u1_N220, 
        u1_N221, u1_N222, u1_N223, u1_N224, u1_N225, u1_N226, u1_N227, u1_N228, u1_N229, 
        u1_N23, u1_N230, u1_N231, u1_N232, u1_N233, u1_N234, u1_N235, u1_N236, u1_N237, 
        u1_N238, u1_N239, u1_N24, u1_N240, u1_N241, u1_N242, u1_N243, u1_N244, u1_N245, 
        u1_N246, u1_N247, u1_N248, u1_N249, u1_N25, u1_N250, u1_N251, u1_N252, u1_N253, 
        u1_N254, u1_N255, u1_N256, u1_N257, u1_N258, u1_N259, u1_N26, u1_N260, u1_N261, 
        u1_N262, u1_N263, u1_N264, u1_N265, u1_N266, u1_N267, u1_N268, u1_N269, u1_N27, 
        u1_N270, u1_N271, u1_N272, u1_N273, u1_N274, u1_N275, u1_N276, u1_N277, u1_N278, 
        u1_N279, u1_N28, u1_N280, u1_N281, u1_N282, u1_N283, u1_N284, u1_N285, u1_N286, 
        u1_N287, u1_N288, u1_N289, u1_N29, u1_N290, u1_N291, u1_N292, u1_N293, u1_N294, 
        u1_N295, u1_N296, u1_N297, u1_N298, u1_N299, u1_N3, u1_N30, u1_N300, u1_N301, 
        u1_N302, u1_N303, u1_N304, u1_N305, u1_N306, u1_N307, u1_N308, u1_N309, u1_N31, 
        u1_N310, u1_N311, u1_N312, u1_N313, u1_N314, u1_N315, u1_N316, u1_N317, u1_N318, 
        u1_N319, u1_N32, u1_N320, u1_N321, u1_N322, u1_N323, u1_N324, u1_N325, u1_N326, 
        u1_N327, u1_N328, u1_N329, u1_N33, u1_N330, u1_N331, u1_N332, u1_N333, u1_N334, 
        u1_N335, u1_N336, u1_N337, u1_N338, u1_N339, u1_N34, u1_N340, u1_N341, u1_N342, 
        u1_N343, u1_N344, u1_N345, u1_N346, u1_N347, u1_N348, u1_N349, u1_N35, u1_N350, 
        u1_N351, u1_N352, u1_N353, u1_N354, u1_N355, u1_N356, u1_N357, u1_N358, u1_N359, 
        u1_N36, u1_N360, u1_N361, u1_N362, u1_N363, u1_N364, u1_N365, u1_N366, u1_N367, 
        u1_N368, u1_N369, u1_N37, u1_N370, u1_N371, u1_N372, u1_N373, u1_N374, u1_N375, 
        u1_N376, u1_N377, u1_N378, u1_N379, u1_N38, u1_N380, u1_N381, u1_N382, u1_N383, 
        u1_N384, u1_N385, u1_N386, u1_N387, u1_N388, u1_N389, u1_N39, u1_N390, u1_N391, 
        u1_N392, u1_N393, u1_N394, u1_N395, u1_N396, u1_N397, u1_N398, u1_N399, u1_N4, 
        u1_N40, u1_N400, u1_N401, u1_N402, u1_N403, u1_N404, u1_N405, u1_N406, u1_N407, 
        u1_N408, u1_N409, u1_N41, u1_N410, u1_N411, u1_N412, u1_N413, u1_N414, u1_N415, 
        u1_N416, u1_N417, u1_N418, u1_N419, u1_N42, u1_N420, u1_N421, u1_N422, u1_N423, 
        u1_N424, u1_N425, u1_N426, u1_N427, u1_N428, u1_N429, u1_N43, u1_N430, u1_N431, 
        u1_N432, u1_N433, u1_N434, u1_N435, u1_N436, u1_N437, u1_N438, u1_N439, u1_N44, 
        u1_N440, u1_N441, u1_N442, u1_N443, u1_N444, u1_N445, u1_N446, u1_N447, u1_N448, 
        u1_N449, u1_N45, u1_N450, u1_N451, u1_N452, u1_N453, u1_N454, u1_N455, u1_N456, 
        u1_N457, u1_N458, u1_N459, u1_N46, u1_N460, u1_N461, u1_N462, u1_N463, u1_N464, 
        u1_N465, u1_N466, u1_N467, u1_N468, u1_N469, u1_N47, u1_N470, u1_N471, u1_N472, 
        u1_N473, u1_N474, u1_N475, u1_N476, u1_N477, u1_N478, u1_N479, u1_N48, u1_N49, 
        u1_N5, u1_N50, u1_N51, u1_N52, u1_N53, u1_N54, u1_N55, u1_N56, u1_N57, 
        u1_N58, u1_N59, u1_N6, u1_N60, u1_N61, u1_N62, u1_N63, u1_N64, u1_N65, 
        u1_N66, u1_N67, u1_N68, u1_N69, u1_N7, u1_N70, u1_N71, u1_N72, u1_N73, 
        u1_N74, u1_N75, u1_N76, u1_N77, u1_N78, u1_N79, u1_N8, u1_N80, u1_N81, 
        u1_N82, u1_N83, u1_N84, u1_N85, u1_N86, u1_N87, u1_N88, u1_N89, u1_N9, 
        u1_N90, u1_N91, u1_N92, u1_N93, u1_N94, u1_N95, u1_N96, u1_N97, u1_N98, 
        u1_N99, u2_FP_1, u2_FP_10, u2_FP_11, u2_FP_12, u2_FP_13, u2_FP_14, u2_FP_15, u2_FP_16, 
        u2_FP_17, u2_FP_18, u2_FP_19, u2_FP_2, u2_FP_20, u2_FP_21, u2_FP_22, u2_FP_23, u2_FP_24, 
        u2_FP_25, u2_FP_26, u2_FP_27, u2_FP_28, u2_FP_29, u2_FP_3, u2_FP_30, u2_FP_31, u2_FP_32, 
        u2_FP_4, u2_FP_5, u2_FP_6, u2_FP_7, u2_FP_8, u2_FP_9, u2_N0, u2_N1, u2_N10, 
        u2_N100, u2_N101, u2_N102, u2_N103, u2_N104, u2_N105, u2_N106, u2_N107, u2_N108, 
        u2_N109, u2_N11, u2_N110, u2_N111, u2_N112, u2_N113, u2_N114, u2_N115, u2_N116, 
        u2_N117, u2_N118, u2_N119, u2_N12, u2_N120, u2_N121, u2_N122, u2_N123, u2_N124, 
        u2_N125, u2_N126, u2_N127, u2_N128, u2_N129, u2_N13, u2_N130, u2_N131, u2_N132, 
        u2_N133, u2_N134, u2_N135, u2_N136, u2_N137, u2_N138, u2_N139, u2_N14, u2_N140, 
        u2_N141, u2_N142, u2_N143, u2_N144, u2_N145, u2_N146, u2_N147, u2_N148, u2_N149, 
        u2_N15, u2_N150, u2_N151, u2_N152, u2_N153, u2_N154, u2_N155, u2_N156, u2_N157, 
        u2_N158, u2_N159, u2_N16, u2_N160, u2_N161, u2_N162, u2_N163, u2_N164, u2_N165, 
        u2_N166, u2_N167, u2_N168, u2_N169, u2_N17, u2_N170, u2_N171, u2_N172, u2_N173, 
        u2_N174, u2_N175, u2_N176, u2_N177, u2_N178, u2_N179, u2_N18, u2_N180, u2_N181, 
        u2_N182, u2_N183, u2_N184, u2_N185, u2_N186, u2_N187, u2_N188, u2_N189, u2_N19, 
        u2_N190, u2_N191, u2_N192, u2_N193, u2_N194, u2_N195, u2_N196, u2_N197, u2_N198, 
        u2_N199, u2_N2, u2_N20, u2_N200, u2_N201, u2_N202, u2_N203, u2_N204, u2_N205, 
        u2_N206, u2_N207, u2_N208, u2_N209, u2_N21, u2_N210, u2_N211, u2_N212, u2_N213, 
        u2_N214, u2_N215, u2_N216, u2_N217, u2_N218, u2_N219, u2_N22, u2_N220, u2_N221, 
        u2_N222, u2_N223, u2_N224, u2_N225, u2_N226, u2_N227, u2_N228, u2_N229, u2_N23, 
        u2_N230, u2_N231, u2_N232, u2_N233, u2_N234, u2_N235, u2_N236, u2_N237, u2_N238, 
        u2_N239, u2_N24, u2_N240, u2_N241, u2_N242, u2_N243, u2_N244, u2_N245, u2_N246, 
        u2_N247, u2_N248, u2_N249, u2_N25, u2_N250, u2_N251, u2_N252, u2_N253, u2_N254, 
        u2_N255, u2_N256, u2_N257, u2_N258, u2_N259, u2_N26, u2_N260, u2_N261, u2_N262, 
        u2_N263, u2_N264, u2_N265, u2_N266, u2_N267, u2_N268, u2_N269, u2_N27, u2_N270, 
        u2_N271, u2_N272, u2_N273, u2_N274, u2_N275, u2_N276, u2_N277, u2_N278, u2_N279, 
        u2_N28, u2_N280, u2_N281, u2_N282, u2_N283, u2_N284, u2_N285, u2_N286, u2_N287, 
        u2_N288, u2_N289, u2_N29, u2_N290, u2_N291, u2_N292, u2_N293, u2_N294, u2_N295, 
        u2_N296, u2_N297, u2_N298, u2_N299, u2_N3, u2_N30, u2_N300, u2_N301, u2_N302, 
        u2_N303, u2_N304, u2_N305, u2_N306, u2_N307, u2_N308, u2_N309, u2_N31, u2_N310, 
        u2_N311, u2_N312, u2_N313, u2_N314, u2_N315, u2_N316, u2_N317, u2_N318, u2_N319, 
        u2_N32, u2_N320, u2_N321, u2_N322, u2_N323, u2_N324, u2_N325, u2_N326, u2_N327, 
        u2_N328, u2_N329, u2_N33, u2_N330, u2_N331, u2_N332, u2_N333, u2_N334, u2_N335, 
        u2_N336, u2_N337, u2_N338, u2_N339, u2_N34, u2_N340, u2_N341, u2_N342, u2_N343, 
        u2_N344, u2_N345, u2_N346, u2_N347, u2_N348, u2_N349, u2_N35, u2_N350, u2_N351, 
        u2_N352, u2_N353, u2_N354, u2_N355, u2_N356, u2_N357, u2_N358, u2_N359, u2_N36, 
        u2_N360, u2_N361, u2_N362, u2_N363, u2_N364, u2_N365, u2_N366, u2_N367, u2_N368, 
        u2_N369, u2_N37, u2_N370, u2_N371, u2_N372, u2_N373, u2_N374, u2_N375, u2_N376, 
        u2_N377, u2_N378, u2_N379, u2_N38, u2_N380, u2_N381, u2_N382, u2_N383, u2_N384, 
        u2_N385, u2_N386, u2_N387, u2_N388, u2_N389, u2_N39, u2_N390, u2_N391, u2_N392, 
        u2_N393, u2_N394, u2_N395, u2_N396, u2_N397, u2_N398, u2_N399, u2_N4, u2_N40, 
        u2_N400, u2_N401, u2_N402, u2_N403, u2_N404, u2_N405, u2_N406, u2_N407, u2_N408, 
        u2_N409, u2_N41, u2_N410, u2_N411, u2_N412, u2_N413, u2_N414, u2_N415, u2_N416, 
        u2_N417, u2_N418, u2_N419, u2_N42, u2_N420, u2_N421, u2_N422, u2_N423, u2_N424, 
        u2_N425, u2_N426, u2_N427, u2_N428, u2_N429, u2_N43, u2_N430, u2_N431, u2_N432, 
        u2_N433, u2_N434, u2_N435, u2_N436, u2_N437, u2_N438, u2_N439, u2_N44, u2_N440, 
        u2_N441, u2_N442, u2_N443, u2_N444, u2_N445, u2_N446, u2_N447, u2_N448, u2_N449, 
        u2_N45, u2_N450, u2_N451, u2_N452, u2_N453, u2_N454, u2_N455, u2_N456, u2_N457, 
        u2_N458, u2_N459, u2_N46, u2_N460, u2_N461, u2_N462, u2_N463, u2_N464, u2_N465, 
        u2_N466, u2_N467, u2_N468, u2_N469, u2_N47, u2_N470, u2_N471, u2_N472, u2_N473, 
        u2_N474, u2_N475, u2_N476, u2_N477, u2_N478, u2_N479, u2_N48, u2_N49, u2_N5, 
        u2_N50, u2_N51, u2_N52, u2_N53, u2_N54, u2_N55, u2_N56, u2_N57, u2_N58, 
        u2_N59, u2_N6, u2_N60, u2_N61, u2_N62, u2_N63, u2_N64, u2_N65, u2_N66, 
        u2_N67, u2_N68, u2_N69, u2_N7, u2_N70, u2_N71, u2_N72, u2_N73, u2_N74, 
        u2_N75, u2_N76, u2_N77, u2_N78, u2_N79, u2_N8, u2_N80, u2_N81, u2_N82, 
        u2_N83, u2_N84, u2_N85, u2_N86, u2_N87, u2_N88, u2_N89, u2_N9, u2_N90, 
        u2_N91, u2_N92, u2_N93, u2_N94, u2_N95, u2_N96, u2_N97, u2_N98, u2_N99, 
        u2_uk_n1012, u2_uk_n1034, u2_uk_n1039, u2_uk_n1056, u2_uk_n1087, u2_uk_n1090, u2_uk_n1102, u2_uk_n1142, u2_uk_n1143, 
        u2_uk_n1144, u2_uk_n1145, u2_uk_n1146, u2_uk_n1148, u2_uk_n1149, u2_uk_n1150, u2_uk_n1152, u2_uk_n1155, u2_uk_n1161, 
        u2_uk_n1162, u2_uk_n1167, u2_uk_n1168, u2_uk_n1171, u2_uk_n1178, u2_uk_n1179, u2_uk_n1183, u2_uk_n1185, u2_uk_n129, 
        u2_uk_n141, u2_uk_n142, u2_uk_n145, u2_uk_n146, u2_uk_n147, u2_uk_n148, u2_uk_n155, u2_uk_n161, u2_uk_n162, 
        u2_uk_n163, u2_uk_n164, u2_uk_n182, u2_uk_n187, u2_uk_n188, u2_uk_n191, u2_uk_n202, u2_uk_n203, u2_uk_n207, 
        u2_uk_n208, u2_uk_n209, u2_uk_n213, u2_uk_n214, u2_uk_n217, u2_uk_n220, u2_uk_n222, u2_uk_n223, u2_uk_n230, 
        u2_uk_n231, u2_uk_n298, u2_uk_n346, u2_uk_n366, u2_uk_n395, u2_uk_n605, u2_uk_n656, u2_uk_n672, u2_uk_n983, 
        u2_uk_n988;
  output n116, u0_FP_33, u0_FP_34, u0_FP_35, u0_FP_36, u0_FP_37, u0_FP_38, u0_FP_39, u0_FP_40, 
        u0_FP_41, u0_FP_42, u0_FP_43, u0_FP_44, u0_FP_45, u0_FP_46, u0_FP_47, u0_FP_48, u0_FP_49, 
        u0_FP_50, u0_FP_51, u0_FP_52, u0_FP_53, u0_FP_54, u0_FP_55, u0_FP_56, u0_FP_57, u0_FP_58, 
        u0_FP_59, u0_FP_60, u0_FP_61, u0_FP_62, u0_FP_63, u0_FP_64, u0_K10_10, u0_K10_13, u0_K10_14, 
        u0_K10_18, u0_K10_19, u0_K10_20, u0_K10_25, u0_K10_27, u0_K10_32, u0_K10_34, u0_K10_36, u0_K10_41, 
        u0_K11_21, u0_K11_37, u0_K11_48, u0_K12_19, u0_K12_22, u0_K12_34, u0_K12_35, u0_K12_36, u0_K12_39, 
        u0_K12_40, u0_K12_48, u0_K12_7, u0_K12_9, u0_K13_30, u0_K13_36, u0_K13_39, u0_K13_40, u0_K13_42, 
        u0_K13_45, u0_K13_46, u0_K13_48, u0_K14_10, u0_K14_12, u0_K14_13, u0_K14_14, u0_K14_15, u0_K14_18, 
        u0_K14_21, u0_K14_24, u0_K14_27, u0_K14_4, u0_K14_42, u0_K14_46, u0_K14_9, u0_K15_18, u0_K15_47, 
        u0_K16_18, u0_K16_19, u0_K16_22, u0_K16_24, u0_K16_26, u0_K16_38, u0_K16_4, u0_K16_8, u0_K1_13, 
        u0_K1_14, u0_K1_15, u0_K1_16, u0_K1_17, u0_K1_23, u0_K1_30, u0_K1_31, u0_K1_45, u0_K1_46, 
        u0_K2_11, u0_K2_12, u0_K2_25, u0_K2_30, u0_K2_34, u0_K2_35, u0_K2_4, u0_K2_44, u0_K2_45, 
        u0_K2_46, u0_K2_47, u0_K2_48, u0_K2_5, u0_K2_6, u0_K2_8, u0_K3_10, u0_K3_12, u0_K3_14, 
        u0_K3_15, u0_K3_17, u0_K3_18, u0_K3_19, u0_K3_23, u0_K3_34, u0_K3_5, u0_K4_24, u0_K4_27, 
        u0_K4_28, u0_K4_35, u0_K4_43, u0_K4_48, u0_K4_6, u0_K5_1, u0_K5_13, u0_K5_14, u0_K5_15, 
        u0_K5_16, u0_K5_18, u0_K5_19, u0_K5_23, u0_K5_24, u0_K5_26, u0_K5_28, u0_K5_3, u0_K5_31, 
        u0_K5_32, u0_K5_34, u0_K5_38, u0_K5_4, u0_K5_41, u0_K5_44, u0_K5_47, u0_K5_48, u0_K5_9, 
        u0_K6_11, u0_K6_13, u0_K6_16, u0_K6_19, u0_K6_20, u0_K6_22, u0_K6_23, u0_K6_24, u0_K6_27, 
        u0_K6_41, u0_K7_2, u0_K7_22, u0_K7_23, u0_K8_1, u0_K8_11, u0_K8_19, u0_K8_28, u0_K8_33, 
        u0_K8_36, u0_K8_45, u0_K9_14, u0_K9_15, u0_K9_32, u0_K9_39, u0_K9_4, u0_K9_40, u0_K9_45, 
        u0_K9_6, u0_L0_1, u0_L0_10, u0_L0_11, u0_L0_12, u0_L0_13, u0_L0_14, u0_L0_15, u0_L0_16, 
        u0_L0_17, u0_L0_18, u0_L0_19, u0_L0_2, u0_L0_20, u0_L0_21, u0_L0_22, u0_L0_23, u0_L0_24, 
        u0_L0_25, u0_L0_26, u0_L0_27, u0_L0_28, u0_L0_29, u0_L0_3, u0_L0_30, u0_L0_31, u0_L0_32, 
        u0_L0_4, u0_L0_5, u0_L0_6, u0_L0_7, u0_L0_8, u0_L0_9, u0_L10_1, u0_L10_10, u0_L10_11, 
        u0_L10_12, u0_L10_13, u0_L10_14, u0_L10_15, u0_L10_16, u0_L10_17, u0_L10_18, u0_L10_19, u0_L10_2, 
        u0_L10_20, u0_L10_21, u0_L10_22, u0_L10_23, u0_L10_24, u0_L10_25, u0_L10_26, u0_L10_27, u0_L10_28, 
        u0_L10_29, u0_L10_3, u0_L10_30, u0_L10_31, u0_L10_32, u0_L10_4, u0_L10_5, u0_L10_6, u0_L10_7, 
        u0_L10_8, u0_L10_9, u0_L11_1, u0_L11_10, u0_L11_11, u0_L11_12, u0_L11_13, u0_L11_14, u0_L11_15, 
        u0_L11_16, u0_L11_17, u0_L11_18, u0_L11_19, u0_L11_2, u0_L11_20, u0_L11_21, u0_L11_22, u0_L11_23, 
        u0_L11_24, u0_L11_25, u0_L11_26, u0_L11_27, u0_L11_28, u0_L11_29, u0_L11_3, u0_L11_30, u0_L11_31, 
        u0_L11_32, u0_L11_4, u0_L11_5, u0_L11_6, u0_L11_7, u0_L11_8, u0_L11_9, u0_L12_1, u0_L12_10, 
        u0_L12_11, u0_L12_12, u0_L12_13, u0_L12_14, u0_L12_15, u0_L12_16, u0_L12_17, u0_L12_18, u0_L12_19, 
        u0_L12_2, u0_L12_20, u0_L12_21, u0_L12_22, u0_L12_23, u0_L12_24, u0_L12_25, u0_L12_26, u0_L12_27, 
        u0_L12_28, u0_L12_29, u0_L12_3, u0_L12_30, u0_L12_31, u0_L12_32, u0_L12_4, u0_L12_5, u0_L12_6, 
        u0_L12_7, u0_L12_8, u0_L12_9, u0_L13_1, u0_L13_10, u0_L13_11, u0_L13_12, u0_L13_13, u0_L13_14, 
        u0_L13_15, u0_L13_16, u0_L13_17, u0_L13_18, u0_L13_19, u0_L13_2, u0_L13_20, u0_L13_21, u0_L13_22, 
        u0_L13_23, u0_L13_24, u0_L13_25, u0_L13_26, u0_L13_27, u0_L13_28, u0_L13_29, u0_L13_3, u0_L13_30, 
        u0_L13_31, u0_L13_32, u0_L13_4, u0_L13_5, u0_L13_6, u0_L13_7, u0_L13_8, u0_L13_9, u0_L14_1, 
        u0_L14_10, u0_L14_11, u0_L14_12, u0_L14_13, u0_L14_14, u0_L14_15, u0_L14_16, u0_L14_17, u0_L14_18, 
        u0_L14_19, u0_L14_2, u0_L14_20, u0_L14_21, u0_L14_22, u0_L14_23, u0_L14_24, u0_L14_25, u0_L14_26, 
        u0_L14_27, u0_L14_28, u0_L14_29, u0_L14_3, u0_L14_30, u0_L14_31, u0_L14_32, u0_L14_4, u0_L14_5, 
        u0_L14_6, u0_L14_7, u0_L14_8, u0_L14_9, u0_L1_1, u0_L1_10, u0_L1_11, u0_L1_12, u0_L1_13, 
        u0_L1_14, u0_L1_15, u0_L1_16, u0_L1_17, u0_L1_18, u0_L1_19, u0_L1_2, u0_L1_20, u0_L1_21, 
        u0_L1_22, u0_L1_23, u0_L1_24, u0_L1_25, u0_L1_26, u0_L1_27, u0_L1_28, u0_L1_29, u0_L1_3, 
        u0_L1_30, u0_L1_31, u0_L1_32, u0_L1_4, u0_L1_5, u0_L1_6, u0_L1_7, u0_L1_8, u0_L1_9, 
        u0_L2_1, u0_L2_10, u0_L2_11, u0_L2_12, u0_L2_13, u0_L2_14, u0_L2_15, u0_L2_16, u0_L2_17, 
        u0_L2_18, u0_L2_19, u0_L2_2, u0_L2_20, u0_L2_21, u0_L2_22, u0_L2_23, u0_L2_24, u0_L2_25, 
        u0_L2_26, u0_L2_27, u0_L2_28, u0_L2_29, u0_L2_3, u0_L2_30, u0_L2_31, u0_L2_32, u0_L2_4, 
        u0_L2_5, u0_L2_6, u0_L2_7, u0_L2_8, u0_L2_9, u0_L3_1, u0_L3_10, u0_L3_11, u0_L3_12, 
        u0_L3_13, u0_L3_14, u0_L3_15, u0_L3_16, u0_L3_17, u0_L3_18, u0_L3_19, u0_L3_2, u0_L3_20, 
        u0_L3_21, u0_L3_22, u0_L3_23, u0_L3_24, u0_L3_25, u0_L3_26, u0_L3_27, u0_L3_28, u0_L3_29, 
        u0_L3_3, u0_L3_30, u0_L3_31, u0_L3_32, u0_L3_4, u0_L3_5, u0_L3_6, u0_L3_7, u0_L3_8, 
        u0_L3_9, u0_L4_1, u0_L4_10, u0_L4_11, u0_L4_12, u0_L4_13, u0_L4_14, u0_L4_15, u0_L4_16, 
        u0_L4_17, u0_L4_18, u0_L4_19, u0_L4_2, u0_L4_20, u0_L4_21, u0_L4_22, u0_L4_23, u0_L4_24, 
        u0_L4_25, u0_L4_26, u0_L4_27, u0_L4_28, u0_L4_29, u0_L4_3, u0_L4_30, u0_L4_31, u0_L4_32, 
        u0_L4_4, u0_L4_5, u0_L4_6, u0_L4_7, u0_L4_8, u0_L4_9, u0_L5_1, u0_L5_10, u0_L5_11, 
        u0_L5_12, u0_L5_13, u0_L5_14, u0_L5_15, u0_L5_16, u0_L5_17, u0_L5_18, u0_L5_19, u0_L5_2, 
        u0_L5_20, u0_L5_21, u0_L5_22, u0_L5_23, u0_L5_24, u0_L5_25, u0_L5_26, u0_L5_27, u0_L5_28, 
        u0_L5_29, u0_L5_3, u0_L5_30, u0_L5_31, u0_L5_32, u0_L5_4, u0_L5_5, u0_L5_6, u0_L5_7, 
        u0_L5_8, u0_L5_9, u0_L6_1, u0_L6_10, u0_L6_11, u0_L6_12, u0_L6_13, u0_L6_14, u0_L6_15, 
        u0_L6_16, u0_L6_17, u0_L6_18, u0_L6_19, u0_L6_2, u0_L6_20, u0_L6_21, u0_L6_22, u0_L6_23, 
        u0_L6_24, u0_L6_25, u0_L6_26, u0_L6_27, u0_L6_28, u0_L6_29, u0_L6_3, u0_L6_30, u0_L6_31, 
        u0_L6_32, u0_L6_4, u0_L6_5, u0_L6_6, u0_L6_7, u0_L6_8, u0_L6_9, u0_L7_1, u0_L7_10, 
        u0_L7_11, u0_L7_12, u0_L7_13, u0_L7_14, u0_L7_15, u0_L7_16, u0_L7_17, u0_L7_18, u0_L7_19, 
        u0_L7_2, u0_L7_20, u0_L7_21, u0_L7_22, u0_L7_23, u0_L7_24, u0_L7_25, u0_L7_26, u0_L7_27, 
        u0_L7_28, u0_L7_29, u0_L7_3, u0_L7_30, u0_L7_31, u0_L7_32, u0_L7_4, u0_L7_5, u0_L7_6, 
        u0_L7_7, u0_L7_8, u0_L7_9, u0_L8_1, u0_L8_10, u0_L8_11, u0_L8_12, u0_L8_13, u0_L8_14, 
        u0_L8_15, u0_L8_16, u0_L8_17, u0_L8_18, u0_L8_19, u0_L8_2, u0_L8_20, u0_L8_21, u0_L8_22, 
        u0_L8_23, u0_L8_24, u0_L8_25, u0_L8_26, u0_L8_27, u0_L8_28, u0_L8_29, u0_L8_3, u0_L8_30, 
        u0_L8_31, u0_L8_32, u0_L8_4, u0_L8_5, u0_L8_6, u0_L8_7, u0_L8_8, u0_L8_9, u0_L9_1, 
        u0_L9_10, u0_L9_11, u0_L9_12, u0_L9_13, u0_L9_14, u0_L9_15, u0_L9_16, u0_L9_17, u0_L9_18, 
        u0_L9_19, u0_L9_2, u0_L9_20, u0_L9_21, u0_L9_22, u0_L9_23, u0_L9_24, u0_L9_25, u0_L9_26, 
        u0_L9_27, u0_L9_28, u0_L9_29, u0_L9_3, u0_L9_30, u0_L9_31, u0_L9_32, u0_L9_4, u0_L9_5, 
        u0_L9_6, u0_L9_7, u0_L9_8, u0_L9_9, u0_R0_1, u0_R0_10, u0_R0_11, u0_R0_12, u0_R0_13, 
        u0_R0_14, u0_R0_15, u0_R0_16, u0_R0_17, u0_R0_18, u0_R0_19, u0_R0_2, u0_R0_20, u0_R0_21, 
        u0_R0_22, u0_R0_23, u0_R0_24, u0_R0_25, u0_R0_26, u0_R0_27, u0_R0_28, u0_R0_29, u0_R0_3, 
        u0_R0_30, u0_R0_31, u0_R0_32, u0_R0_4, u0_R0_5, u0_R0_6, u0_R0_7, u0_R0_8, u0_R0_9, 
        u0_R10_1, u0_R10_10, u0_R10_11, u0_R10_12, u0_R10_13, u0_R10_14, u0_R10_15, u0_R10_16, u0_R10_17, 
        u0_R10_18, u0_R10_19, u0_R10_2, u0_R10_20, u0_R10_21, u0_R10_22, u0_R10_23, u0_R10_24, u0_R10_25, 
        u0_R10_26, u0_R10_27, u0_R10_28, u0_R10_29, u0_R10_3, u0_R10_30, u0_R10_31, u0_R10_32, u0_R10_4, 
        u0_R10_5, u0_R10_6, u0_R10_7, u0_R10_8, u0_R10_9, u0_R11_1, u0_R11_10, u0_R11_11, u0_R11_12, 
        u0_R11_13, u0_R11_14, u0_R11_15, u0_R11_16, u0_R11_17, u0_R11_18, u0_R11_19, u0_R11_2, u0_R11_20, 
        u0_R11_21, u0_R11_22, u0_R11_23, u0_R11_24, u0_R11_25, u0_R11_26, u0_R11_27, u0_R11_28, u0_R11_29, 
        u0_R11_3, u0_R11_30, u0_R11_31, u0_R11_32, u0_R11_4, u0_R11_5, u0_R11_6, u0_R11_7, u0_R11_8, 
        u0_R11_9, u0_R12_1, u0_R12_10, u0_R12_11, u0_R12_12, u0_R12_13, u0_R12_14, u0_R12_15, u0_R12_16, 
        u0_R12_17, u0_R12_18, u0_R12_19, u0_R12_2, u0_R12_20, u0_R12_21, u0_R12_22, u0_R12_23, u0_R12_24, 
        u0_R12_25, u0_R12_26, u0_R12_27, u0_R12_28, u0_R12_29, u0_R12_3, u0_R12_30, u0_R12_31, u0_R12_32, 
        u0_R12_4, u0_R12_5, u0_R12_6, u0_R12_7, u0_R12_8, u0_R12_9, u0_R13_1, u0_R13_10, u0_R13_11, 
        u0_R13_12, u0_R13_13, u0_R13_14, u0_R13_15, u0_R13_16, u0_R13_17, u0_R13_18, u0_R13_19, u0_R13_2, 
        u0_R13_20, u0_R13_21, u0_R13_22, u0_R13_23, u0_R13_24, u0_R13_25, u0_R13_26, u0_R13_27, u0_R13_28, 
        u0_R13_29, u0_R13_3, u0_R13_30, u0_R13_31, u0_R13_32, u0_R13_4, u0_R13_5, u0_R13_6, u0_R13_7, 
        u0_R13_8, u0_R13_9, u0_R1_1, u0_R1_10, u0_R1_11, u0_R1_12, u0_R1_13, u0_R1_14, u0_R1_15, 
        u0_R1_16, u0_R1_17, u0_R1_18, u0_R1_19, u0_R1_2, u0_R1_20, u0_R1_21, u0_R1_22, u0_R1_23, 
        u0_R1_24, u0_R1_25, u0_R1_26, u0_R1_27, u0_R1_28, u0_R1_29, u0_R1_3, u0_R1_30, u0_R1_31, 
        u0_R1_32, u0_R1_4, u0_R1_5, u0_R1_6, u0_R1_7, u0_R1_8, u0_R1_9, u0_R2_1, u0_R2_10, 
        u0_R2_11, u0_R2_12, u0_R2_13, u0_R2_14, u0_R2_15, u0_R2_16, u0_R2_17, u0_R2_18, u0_R2_19, 
        u0_R2_2, u0_R2_20, u0_R2_21, u0_R2_22, u0_R2_23, u0_R2_24, u0_R2_25, u0_R2_26, u0_R2_27, 
        u0_R2_28, u0_R2_29, u0_R2_3, u0_R2_30, u0_R2_31, u0_R2_32, u0_R2_4, u0_R2_5, u0_R2_6, 
        u0_R2_7, u0_R2_8, u0_R2_9, u0_R3_1, u0_R3_10, u0_R3_11, u0_R3_12, u0_R3_13, u0_R3_14, 
        u0_R3_15, u0_R3_16, u0_R3_17, u0_R3_18, u0_R3_19, u0_R3_2, u0_R3_20, u0_R3_21, u0_R3_22, 
        u0_R3_23, u0_R3_24, u0_R3_25, u0_R3_26, u0_R3_27, u0_R3_28, u0_R3_29, u0_R3_3, u0_R3_30, 
        u0_R3_31, u0_R3_32, u0_R3_4, u0_R3_5, u0_R3_6, u0_R3_7, u0_R3_8, u0_R3_9, u0_R4_1, 
        u0_R4_10, u0_R4_11, u0_R4_12, u0_R4_13, u0_R4_14, u0_R4_15, u0_R4_16, u0_R4_17, u0_R4_18, 
        u0_R4_19, u0_R4_2, u0_R4_20, u0_R4_21, u0_R4_22, u0_R4_23, u0_R4_24, u0_R4_25, u0_R4_26, 
        u0_R4_27, u0_R4_28, u0_R4_29, u0_R4_3, u0_R4_30, u0_R4_31, u0_R4_32, u0_R4_4, u0_R4_5, 
        u0_R4_6, u0_R4_7, u0_R4_8, u0_R4_9, u0_R5_1, u0_R5_10, u0_R5_11, u0_R5_12, u0_R5_13, 
        u0_R5_14, u0_R5_15, u0_R5_16, u0_R5_17, u0_R5_18, u0_R5_19, u0_R5_2, u0_R5_20, u0_R5_21, 
        u0_R5_22, u0_R5_23, u0_R5_24, u0_R5_25, u0_R5_26, u0_R5_27, u0_R5_28, u0_R5_29, u0_R5_3, 
        u0_R5_30, u0_R5_31, u0_R5_32, u0_R5_4, u0_R5_5, u0_R5_6, u0_R5_7, u0_R5_8, u0_R5_9, 
        u0_R6_1, u0_R6_10, u0_R6_11, u0_R6_12, u0_R6_13, u0_R6_14, u0_R6_15, u0_R6_16, u0_R6_17, 
        u0_R6_18, u0_R6_19, u0_R6_2, u0_R6_20, u0_R6_21, u0_R6_22, u0_R6_23, u0_R6_24, u0_R6_25, 
        u0_R6_26, u0_R6_27, u0_R6_28, u0_R6_29, u0_R6_3, u0_R6_30, u0_R6_31, u0_R6_32, u0_R6_4, 
        u0_R6_5, u0_R6_6, u0_R6_7, u0_R6_8, u0_R6_9, u0_R7_1, u0_R7_10, u0_R7_11, u0_R7_12, 
        u0_R7_13, u0_R7_14, u0_R7_15, u0_R7_16, u0_R7_17, u0_R7_18, u0_R7_19, u0_R7_2, u0_R7_20, 
        u0_R7_21, u0_R7_22, u0_R7_23, u0_R7_24, u0_R7_25, u0_R7_26, u0_R7_27, u0_R7_28, u0_R7_29, 
        u0_R7_3, u0_R7_30, u0_R7_31, u0_R7_32, u0_R7_4, u0_R7_5, u0_R7_6, u0_R7_7, u0_R7_8, 
        u0_R7_9, u0_R8_1, u0_R8_10, u0_R8_11, u0_R8_12, u0_R8_13, u0_R8_14, u0_R8_15, u0_R8_16, 
        u0_R8_17, u0_R8_18, u0_R8_19, u0_R8_2, u0_R8_20, u0_R8_21, u0_R8_22, u0_R8_23, u0_R8_24, 
        u0_R8_25, u0_R8_26, u0_R8_27, u0_R8_28, u0_R8_29, u0_R8_3, u0_R8_30, u0_R8_31, u0_R8_32, 
        u0_R8_4, u0_R8_5, u0_R8_6, u0_R8_7, u0_R8_8, u0_R8_9, u0_R9_1, u0_R9_10, u0_R9_11, 
        u0_R9_12, u0_R9_13, u0_R9_14, u0_R9_15, u0_R9_16, u0_R9_17, u0_R9_18, u0_R9_19, u0_R9_2, 
        u0_R9_20, u0_R9_21, u0_R9_22, u0_R9_23, u0_R9_24, u0_R9_25, u0_R9_26, u0_R9_27, u0_R9_28, 
        u0_R9_29, u0_R9_3, u0_R9_30, u0_R9_31, u0_R9_32, u0_R9_4, u0_R9_5, u0_R9_6, u0_R9_7, 
        u0_R9_8, u0_R9_9, u0_desIn_r_0, u0_desIn_r_1, u0_desIn_r_10, u0_desIn_r_11, u0_desIn_r_12, u0_desIn_r_13, u0_desIn_r_14, 
        u0_desIn_r_15, u0_desIn_r_16, u0_desIn_r_17, u0_desIn_r_18, u0_desIn_r_19, u0_desIn_r_2, u0_desIn_r_20, u0_desIn_r_21, u0_desIn_r_22, 
        u0_desIn_r_23, u0_desIn_r_24, u0_desIn_r_25, u0_desIn_r_26, u0_desIn_r_27, u0_desIn_r_28, u0_desIn_r_29, u0_desIn_r_3, u0_desIn_r_30, 
        u0_desIn_r_31, u0_desIn_r_32, u0_desIn_r_33, u0_desIn_r_34, u0_desIn_r_35, u0_desIn_r_36, u0_desIn_r_37, u0_desIn_r_38, u0_desIn_r_39, 
        u0_desIn_r_4, u0_desIn_r_40, u0_desIn_r_41, u0_desIn_r_42, u0_desIn_r_43, u0_desIn_r_44, u0_desIn_r_45, u0_desIn_r_46, u0_desIn_r_47, 
        u0_desIn_r_48, u0_desIn_r_49, u0_desIn_r_5, u0_desIn_r_50, u0_desIn_r_51, u0_desIn_r_52, u0_desIn_r_53, u0_desIn_r_54, u0_desIn_r_55, 
        u0_desIn_r_56, u0_desIn_r_57, u0_desIn_r_58, u0_desIn_r_59, u0_desIn_r_6, u0_desIn_r_60, u0_desIn_r_61, u0_desIn_r_62, u0_desIn_r_63, 
        u0_desIn_r_7, u0_desIn_r_8, u0_desIn_r_9, u0_key_r_0, u0_key_r_1, u0_key_r_10, u0_key_r_11, u0_key_r_12, u0_key_r_13, 
        u0_key_r_14, u0_key_r_16, u0_key_r_17, u0_key_r_18, u0_key_r_19, u0_key_r_2, u0_key_r_20, u0_key_r_21, u0_key_r_22, 
        u0_key_r_23, u0_key_r_24, u0_key_r_25, u0_key_r_26, u0_key_r_27, u0_key_r_28, u0_key_r_29, u0_key_r_3, u0_key_r_30, 
        u0_key_r_31, u0_key_r_32, u0_key_r_33, u0_key_r_34, u0_key_r_35, u0_key_r_36, u0_key_r_37, u0_key_r_38, u0_key_r_39, 
        u0_key_r_4, u0_key_r_40, u0_key_r_41, u0_key_r_42, u0_key_r_43, u0_key_r_44, u0_key_r_45, u0_key_r_46, u0_key_r_47, 
        u0_key_r_48, u0_key_r_49, u0_key_r_5, u0_key_r_50, u0_key_r_51, u0_key_r_52, u0_key_r_53, u0_key_r_54, u0_key_r_55, 
        u0_key_r_6, u0_key_r_7, u0_key_r_8, u0_key_r_9, u0_uk_K_r0_11, u0_uk_K_r0_15, u0_uk_K_r0_19, u0_uk_K_r0_2, u0_uk_K_r0_22, 
        u0_uk_K_r0_25, u0_uk_K_r0_28, u0_uk_K_r0_31, u0_uk_K_r0_32, u0_uk_K_r0_34, u0_uk_K_r0_36, u0_uk_K_r0_47, u0_uk_K_r0_49, u0_uk_K_r0_52, 
        u0_uk_K_r0_55, u0_uk_K_r0_7, u0_uk_K_r10_10, u0_uk_K_r10_14, u0_uk_K_r10_16, u0_uk_K_r10_18, u0_uk_K_r10_19, u0_uk_K_r10_23, u0_uk_K_r10_25, 
        u0_uk_K_r10_27, u0_uk_K_r10_28, u0_uk_K_r10_32, u0_uk_K_r10_34, u0_uk_K_r10_37, u0_uk_K_r10_39, u0_uk_K_r10_41, u0_uk_K_r10_42, u0_uk_K_r10_43, 
        u0_uk_K_r10_44, u0_uk_K_r10_47, u0_uk_K_r10_48, u0_uk_K_r10_9, u0_uk_K_r11_10, u0_uk_K_r11_11, u0_uk_K_r11_17, u0_uk_K_r11_19, u0_uk_K_r11_20, 
        u0_uk_K_r11_21, u0_uk_K_r11_24, u0_uk_K_r11_25, u0_uk_K_r11_26, u0_uk_K_r11_27, u0_uk_K_r11_28, u0_uk_K_r11_29, u0_uk_K_r11_33, u0_uk_K_r11_34, 
        u0_uk_K_r11_39, u0_uk_K_r11_4, u0_uk_K_r11_46, u0_uk_K_r11_47, u0_uk_K_r11_48, u0_uk_K_r11_53, u0_uk_K_r11_54, u0_uk_K_r11_6, u0_uk_K_r11_8, 
        u0_uk_K_r12_1, u0_uk_K_r12_10, u0_uk_K_r12_15, u0_uk_K_r12_16, u0_uk_K_r12_18, u0_uk_K_r12_21, u0_uk_K_r12_25, u0_uk_K_r12_30, u0_uk_K_r12_33, 
        u0_uk_K_r12_36, u0_uk_K_r12_42, u0_uk_K_r12_44, u0_uk_K_r12_47, u0_uk_K_r12_7, u0_uk_K_r13_0, u0_uk_K_r13_13, u0_uk_K_r13_17, u0_uk_K_r13_19, 
        u0_uk_K_r13_2, u0_uk_K_r13_22, u0_uk_K_r13_23, u0_uk_K_r13_25, u0_uk_K_r13_32, u0_uk_K_r13_35, u0_uk_K_r13_38, u0_uk_K_r13_4, u0_uk_K_r13_44, 
        u0_uk_K_r13_55, u0_uk_K_r14_10, u0_uk_K_r14_11, u0_uk_K_r14_12, u0_uk_K_r14_15, u0_uk_K_r14_16, u0_uk_K_r14_18, u0_uk_K_r14_2, u0_uk_K_r14_3, 
        u0_uk_K_r14_39, u0_uk_K_r14_43, u0_uk_K_r14_45, u0_uk_K_r14_46, u0_uk_K_r14_5, u0_uk_K_r14_50, u0_uk_K_r14_8, u0_uk_K_r14_9, u0_uk_K_r1_10, 
        u0_uk_K_r1_15, u0_uk_K_r1_16, u0_uk_K_r1_17, u0_uk_K_r1_18, u0_uk_K_r1_21, u0_uk_K_r1_22, u0_uk_K_r1_36, u0_uk_K_r1_41, u0_uk_K_r1_42, 
        u0_uk_K_r1_44, u0_uk_K_r1_47, u0_uk_K_r1_7, u0_uk_K_r2_13, u0_uk_K_r2_16, u0_uk_K_r2_18, u0_uk_K_r2_20, u0_uk_K_r2_25, u0_uk_K_r2_26, 
        u0_uk_K_r2_27, u0_uk_K_r2_28, u0_uk_K_r2_29, u0_uk_K_r2_31, u0_uk_K_r2_33, u0_uk_K_r2_36, u0_uk_K_r2_4, u0_uk_K_r2_41, u0_uk_K_r2_46, 
        u0_uk_K_r2_50, u0_uk_K_r2_53, u0_uk_K_r2_55, u0_uk_K_r2_7, u0_uk_K_r3_10, u0_uk_K_r3_11, u0_uk_K_r3_14, u0_uk_K_r3_15, u0_uk_K_r3_16, 
        u0_uk_K_r3_19, u0_uk_K_r3_24, u0_uk_K_r3_29, u0_uk_K_r3_35, u0_uk_K_r3_38, u0_uk_K_r3_4, u0_uk_K_r3_47, u0_uk_K_r3_52, u0_uk_K_r3_9, 
        u0_uk_K_r4_0, u0_uk_K_r4_11, u0_uk_K_r4_23, u0_uk_K_r4_3, u0_uk_K_r4_31, u0_uk_K_r4_33, u0_uk_K_r4_35, u0_uk_K_r4_38, u0_uk_K_r4_4, 
        u0_uk_K_r4_41, u0_uk_K_r4_47, u0_uk_K_r4_48, u0_uk_K_r4_49, u0_uk_K_r4_5, u0_uk_K_r4_54, u0_uk_K_r4_55, u0_uk_K_r5_0, u0_uk_K_r5_1, 
        u0_uk_K_r5_10, u0_uk_K_r5_13, u0_uk_K_r5_16, u0_uk_K_r5_17, u0_uk_K_r5_18, u0_uk_K_r5_19, u0_uk_K_r5_21, u0_uk_K_r5_23, u0_uk_K_r5_26, 
        u0_uk_K_r5_32, u0_uk_K_r5_37, u0_uk_K_r5_39, u0_uk_K_r5_4, u0_uk_K_r5_40, u0_uk_K_r5_41, u0_uk_K_r5_43, u0_uk_K_r5_48, u0_uk_K_r5_5, 
        u0_uk_K_r5_51, u0_uk_K_r5_8, u0_uk_K_r6_0, u0_uk_K_r6_10, u0_uk_K_r6_14, u0_uk_K_r6_19, u0_uk_K_r6_21, u0_uk_K_r6_22, u0_uk_K_r6_26, 
        u0_uk_K_r6_27, u0_uk_K_r6_29, u0_uk_K_r6_3, u0_uk_K_r6_31, u0_uk_K_r6_34, u0_uk_K_r6_37, u0_uk_K_r6_46, u0_uk_K_r6_51, u0_uk_K_r6_53, 
        u0_uk_K_r6_55, u0_uk_K_r6_7, u0_uk_K_r7_0, u0_uk_K_r7_1, u0_uk_K_r7_13, u0_uk_K_r7_15, u0_uk_K_r7_2, u0_uk_K_r7_20, u0_uk_K_r7_22, 
        u0_uk_K_r7_23, u0_uk_K_r7_24, u0_uk_K_r7_25, u0_uk_K_r7_26, u0_uk_K_r7_27, u0_uk_K_r7_30, u0_uk_K_r7_32, u0_uk_K_r7_39, u0_uk_K_r7_48, 
        u0_uk_K_r7_55, u0_uk_K_r7_6, u0_uk_K_r7_8, u0_uk_K_r7_9, u0_uk_K_r8_13, u0_uk_K_r8_16, u0_uk_K_r8_17, u0_uk_K_r8_2, u0_uk_K_r8_21, 
        u0_uk_K_r8_22, u0_uk_K_r8_27, u0_uk_K_r8_28, u0_uk_K_r8_32, u0_uk_K_r8_37, u0_uk_K_r8_40, u0_uk_K_r8_41, u0_uk_K_r8_43, u0_uk_K_r8_44, 
        u0_uk_K_r8_52, u0_uk_K_r8_8, u0_uk_K_r9_0, u0_uk_K_r9_1, u0_uk_K_r9_10, u0_uk_K_r9_12, u0_uk_K_r9_13, u0_uk_K_r9_15, u0_uk_K_r9_18, 
        u0_uk_K_r9_19, u0_uk_K_r9_22, u0_uk_K_r9_23, u0_uk_K_r9_25, u0_uk_K_r9_27, u0_uk_K_r9_30, u0_uk_K_r9_31, u0_uk_K_r9_33, u0_uk_K_r9_35, 
        u0_uk_K_r9_38, u0_uk_K_r9_45, u0_uk_K_r9_48, u0_uk_K_r9_49, u0_uk_K_r9_5, u0_uk_K_r9_6, u0_uk_K_r9_7, u0_uk_K_r9_9, u0_uk_n1, 
        u0_uk_n1001, u0_uk_n1002, u0_uk_n1004, u0_uk_n1009, u0_uk_n101, u0_uk_n1012, u0_uk_n1019, u0_uk_n1020, u0_uk_n1021, 
        u0_uk_n1024, u0_uk_n103, u0_uk_n104, u0_uk_n105, u0_uk_n106, u0_uk_n107, u0_uk_n108, u0_uk_n111, u0_uk_n112, 
        u0_uk_n113, u0_uk_n115, u0_uk_n116, u0_uk_n119, u0_uk_n12, u0_uk_n120, u0_uk_n121, u0_uk_n122, u0_uk_n123, 
        u0_uk_n124, u0_uk_n126, u0_uk_n127, u0_uk_n13, u0_uk_n130, u0_uk_n131, u0_uk_n132, u0_uk_n134, u0_uk_n135, 
        u0_uk_n136, u0_uk_n137, u0_uk_n139, u0_uk_n14, u0_uk_n140, u0_uk_n143, u0_uk_n144, u0_uk_n149, u0_uk_n15, 
        u0_uk_n150, u0_uk_n151, u0_uk_n152, u0_uk_n153, u0_uk_n154, u0_uk_n156, u0_uk_n157, u0_uk_n159, u0_uk_n16, 
        u0_uk_n165, u0_uk_n166, u0_uk_n167, u0_uk_n168, u0_uk_n169, u0_uk_n170, u0_uk_n171, u0_uk_n172, u0_uk_n173, 
        u0_uk_n174, u0_uk_n175, u0_uk_n176, u0_uk_n177, u0_uk_n178, u0_uk_n179, u0_uk_n18, u0_uk_n180, u0_uk_n181, 
        u0_uk_n183, u0_uk_n184, u0_uk_n185, u0_uk_n186, u0_uk_n189, u0_uk_n19, u0_uk_n190, u0_uk_n192, u0_uk_n193, 
        u0_uk_n194, u0_uk_n195, u0_uk_n196, u0_uk_n197, u0_uk_n198, u0_uk_n199, u0_uk_n20, u0_uk_n200, u0_uk_n201, 
        u0_uk_n204, u0_uk_n205, u0_uk_n206, u0_uk_n21, u0_uk_n210, u0_uk_n211, u0_uk_n212, u0_uk_n215, u0_uk_n216, 
        u0_uk_n218, u0_uk_n219, u0_uk_n22, u0_uk_n221, u0_uk_n224, u0_uk_n225, u0_uk_n226, u0_uk_n227, u0_uk_n228, 
        u0_uk_n229, u0_uk_n23, u0_uk_n232, u0_uk_n233, u0_uk_n234, u0_uk_n235, u0_uk_n237, u0_uk_n239, u0_uk_n24, 
        u0_uk_n241, u0_uk_n243, u0_uk_n244, u0_uk_n245, u0_uk_n246, u0_uk_n247, u0_uk_n248, u0_uk_n249, u0_uk_n25, 
        u0_uk_n253, u0_uk_n254, u0_uk_n255, u0_uk_n256, u0_uk_n257, u0_uk_n258, u0_uk_n259, u0_uk_n26, u0_uk_n260, 
        u0_uk_n261, u0_uk_n262, u0_uk_n263, u0_uk_n264, u0_uk_n265, u0_uk_n266, u0_uk_n267, u0_uk_n268, u0_uk_n269, 
        u0_uk_n272, u0_uk_n273, u0_uk_n274, u0_uk_n275, u0_uk_n276, u0_uk_n278, u0_uk_n28, u0_uk_n280, u0_uk_n281, 
        u0_uk_n282, u0_uk_n283, u0_uk_n285, u0_uk_n288, u0_uk_n289, u0_uk_n29, u0_uk_n290, u0_uk_n293, u0_uk_n296, 
        u0_uk_n3, u0_uk_n30, u0_uk_n300, u0_uk_n303, u0_uk_n304, u0_uk_n307, u0_uk_n309, u0_uk_n310, u0_uk_n311, 
        u0_uk_n314, u0_uk_n315, u0_uk_n316, u0_uk_n318, u0_uk_n32, u0_uk_n320, u0_uk_n321, u0_uk_n322, u0_uk_n323, 
        u0_uk_n324, u0_uk_n325, u0_uk_n326, u0_uk_n327, u0_uk_n328, u0_uk_n329, u0_uk_n33, u0_uk_n330, u0_uk_n331, 
        u0_uk_n332, u0_uk_n333, u0_uk_n336, u0_uk_n337, u0_uk_n339, u0_uk_n34, u0_uk_n340, u0_uk_n341, u0_uk_n343, 
        u0_uk_n344, u0_uk_n345, u0_uk_n347, u0_uk_n348, u0_uk_n35, u0_uk_n350, u0_uk_n351, u0_uk_n352, u0_uk_n354, 
        u0_uk_n355, u0_uk_n356, u0_uk_n357, u0_uk_n358, u0_uk_n359, u0_uk_n36, u0_uk_n361, u0_uk_n362, u0_uk_n364, 
        u0_uk_n365, u0_uk_n367, u0_uk_n368, u0_uk_n37, u0_uk_n370, u0_uk_n371, u0_uk_n372, u0_uk_n374, u0_uk_n378, 
        u0_uk_n38, u0_uk_n380, u0_uk_n381, u0_uk_n383, u0_uk_n384, u0_uk_n387, u0_uk_n388, u0_uk_n389, u0_uk_n39, 
        u0_uk_n390, u0_uk_n392, u0_uk_n393, u0_uk_n394, u0_uk_n396, u0_uk_n397, u0_uk_n398, u0_uk_n399, u0_uk_n4, 
        u0_uk_n40, u0_uk_n400, u0_uk_n401, u0_uk_n402, u0_uk_n403, u0_uk_n404, u0_uk_n405, u0_uk_n406, u0_uk_n41, 
        u0_uk_n410, u0_uk_n411, u0_uk_n412, u0_uk_n413, u0_uk_n414, u0_uk_n417, u0_uk_n418, u0_uk_n419, u0_uk_n42, 
        u0_uk_n420, u0_uk_n423, u0_uk_n424, u0_uk_n425, u0_uk_n426, u0_uk_n427, u0_uk_n428, u0_uk_n429, u0_uk_n43, 
        u0_uk_n430, u0_uk_n432, u0_uk_n433, u0_uk_n434, u0_uk_n435, u0_uk_n436, u0_uk_n438, u0_uk_n439, u0_uk_n44, 
        u0_uk_n440, u0_uk_n441, u0_uk_n442, u0_uk_n445, u0_uk_n446, u0_uk_n447, u0_uk_n448, u0_uk_n45, u0_uk_n450, 
        u0_uk_n451, u0_uk_n453, u0_uk_n455, u0_uk_n457, u0_uk_n458, u0_uk_n459, u0_uk_n46, u0_uk_n462, u0_uk_n463, 
        u0_uk_n464, u0_uk_n465, u0_uk_n466, u0_uk_n471, u0_uk_n473, u0_uk_n475, u0_uk_n476, u0_uk_n479, u0_uk_n48, 
        u0_uk_n480, u0_uk_n481, u0_uk_n482, u0_uk_n483, u0_uk_n484, u0_uk_n485, u0_uk_n486, u0_uk_n488, u0_uk_n489, 
        u0_uk_n49, u0_uk_n490, u0_uk_n491, u0_uk_n493, u0_uk_n494, u0_uk_n497, u0_uk_n498, u0_uk_n499, u0_uk_n5, 
        u0_uk_n50, u0_uk_n502, u0_uk_n505, u0_uk_n506, u0_uk_n507, u0_uk_n508, u0_uk_n51, u0_uk_n510, u0_uk_n511, 
        u0_uk_n512, u0_uk_n513, u0_uk_n514, u0_uk_n516, u0_uk_n517, u0_uk_n519, u0_uk_n52, u0_uk_n521, u0_uk_n522, 
        u0_uk_n523, u0_uk_n525, u0_uk_n527, u0_uk_n528, u0_uk_n529, u0_uk_n53, u0_uk_n530, u0_uk_n531, u0_uk_n532, 
        u0_uk_n534, u0_uk_n535, u0_uk_n536, u0_uk_n537, u0_uk_n538, u0_uk_n539, u0_uk_n54, u0_uk_n540, u0_uk_n542, 
        u0_uk_n543, u0_uk_n544, u0_uk_n545, u0_uk_n546, u0_uk_n547, u0_uk_n549, u0_uk_n55, u0_uk_n550, u0_uk_n552, 
        u0_uk_n553, u0_uk_n554, u0_uk_n555, u0_uk_n557, u0_uk_n558, u0_uk_n559, u0_uk_n56, u0_uk_n560, u0_uk_n561, 
        u0_uk_n562, u0_uk_n563, u0_uk_n564, u0_uk_n565, u0_uk_n566, u0_uk_n567, u0_uk_n568, u0_uk_n569, u0_uk_n57, 
        u0_uk_n570, u0_uk_n571, u0_uk_n573, u0_uk_n574, u0_uk_n575, u0_uk_n576, u0_uk_n577, u0_uk_n578, u0_uk_n579, 
        u0_uk_n58, u0_uk_n580, u0_uk_n581, u0_uk_n583, u0_uk_n584, u0_uk_n588, u0_uk_n589, u0_uk_n59, u0_uk_n592, 
        u0_uk_n593, u0_uk_n594, u0_uk_n596, u0_uk_n597, u0_uk_n598, u0_uk_n599, u0_uk_n6, u0_uk_n600, u0_uk_n604, 
        u0_uk_n606, u0_uk_n607, u0_uk_n609, u0_uk_n61, u0_uk_n610, u0_uk_n611, u0_uk_n612, u0_uk_n613, u0_uk_n614, 
        u0_uk_n615, u0_uk_n616, u0_uk_n619, u0_uk_n62, u0_uk_n620, u0_uk_n621, u0_uk_n622, u0_uk_n623, u0_uk_n624, 
        u0_uk_n625, u0_uk_n626, u0_uk_n627, u0_uk_n628, u0_uk_n629, u0_uk_n630, u0_uk_n631, u0_uk_n632, u0_uk_n633, 
        u0_uk_n635, u0_uk_n636, u0_uk_n637, u0_uk_n638, u0_uk_n639, u0_uk_n64, u0_uk_n640, u0_uk_n641, u0_uk_n642, 
        u0_uk_n643, u0_uk_n644, u0_uk_n645, u0_uk_n646, u0_uk_n647, u0_uk_n648, u0_uk_n649, u0_uk_n65, u0_uk_n650, 
        u0_uk_n651, u0_uk_n652, u0_uk_n653, u0_uk_n654, u0_uk_n655, u0_uk_n657, u0_uk_n658, u0_uk_n659, u0_uk_n66, 
        u0_uk_n660, u0_uk_n661, u0_uk_n663, u0_uk_n664, u0_uk_n666, u0_uk_n667, u0_uk_n668, u0_uk_n669, u0_uk_n67, 
        u0_uk_n670, u0_uk_n68, u0_uk_n69, u0_uk_n7, u0_uk_n719, u0_uk_n72, u0_uk_n720, u0_uk_n725, u0_uk_n726, 
        u0_uk_n728, u0_uk_n73, u0_uk_n731, u0_uk_n732, u0_uk_n735, u0_uk_n736, u0_uk_n739, u0_uk_n740, u0_uk_n746, 
        u0_uk_n748, u0_uk_n75, u0_uk_n755, u0_uk_n759, u0_uk_n763, u0_uk_n765, u0_uk_n766, u0_uk_n77, u0_uk_n770, 
        u0_uk_n775, u0_uk_n78, u0_uk_n780, u0_uk_n785, u0_uk_n786, u0_uk_n79, u0_uk_n793, u0_uk_n799, u0_uk_n8, 
        u0_uk_n80, u0_uk_n805, u0_uk_n81, u0_uk_n810, u0_uk_n813, u0_uk_n815, u0_uk_n82, u0_uk_n826, u0_uk_n832, 
        u0_uk_n834, u0_uk_n839, u0_uk_n84, u0_uk_n85, u0_uk_n853, u0_uk_n855, u0_uk_n86, u0_uk_n87, u0_uk_n875, 
        u0_uk_n878, u0_uk_n88, u0_uk_n89, u0_uk_n897, u0_uk_n898, u0_uk_n9, u0_uk_n90, u0_uk_n904, u0_uk_n91, 
        u0_uk_n916, u0_uk_n917, u0_uk_n918, u0_uk_n939, u0_uk_n948, u0_uk_n95, u0_uk_n950, u0_uk_n96, u0_uk_n960, 
        u0_uk_n963, u0_uk_n97, u0_uk_n98, u0_uk_n981, u0_uk_n990, u0_uk_n999, u1_FP_33, u1_FP_34, u1_FP_35, 
        u1_FP_36, u1_FP_37, u1_FP_38, u1_FP_39, u1_FP_40, u1_FP_41, u1_FP_42, u1_FP_43, u1_FP_44, 
        u1_FP_45, u1_FP_46, u1_FP_47, u1_FP_48, u1_FP_49, u1_FP_50, u1_FP_51, u1_FP_52, u1_FP_53, 
        u1_FP_54, u1_FP_55, u1_FP_56, u1_FP_57, u1_FP_58, u1_FP_59, u1_FP_60, u1_FP_61, u1_FP_62, 
        u1_FP_63, u1_FP_64, u1_L0_1, u1_L0_10, u1_L0_11, u1_L0_12, u1_L0_13, u1_L0_14, u1_L0_15, 
        u1_L0_16, u1_L0_17, u1_L0_18, u1_L0_19, u1_L0_2, u1_L0_20, u1_L0_21, u1_L0_22, u1_L0_23, 
        u1_L0_24, u1_L0_25, u1_L0_26, u1_L0_27, u1_L0_28, u1_L0_29, u1_L0_3, u1_L0_30, u1_L0_31, 
        u1_L0_32, u1_L0_4, u1_L0_5, u1_L0_6, u1_L0_7, u1_L0_8, u1_L0_9, u1_L10_1, u1_L10_10, 
        u1_L10_11, u1_L10_12, u1_L10_13, u1_L10_14, u1_L10_15, u1_L10_16, u1_L10_17, u1_L10_18, u1_L10_19, 
        u1_L10_2, u1_L10_20, u1_L10_21, u1_L10_22, u1_L10_23, u1_L10_24, u1_L10_25, u1_L10_26, u1_L10_27, 
        u1_L10_28, u1_L10_29, u1_L10_3, u1_L10_30, u1_L10_31, u1_L10_32, u1_L10_4, u1_L10_5, u1_L10_6, 
        u1_L10_7, u1_L10_8, u1_L10_9, u1_L11_1, u1_L11_10, u1_L11_11, u1_L11_12, u1_L11_13, u1_L11_14, 
        u1_L11_15, u1_L11_16, u1_L11_17, u1_L11_18, u1_L11_19, u1_L11_2, u1_L11_20, u1_L11_21, u1_L11_22, 
        u1_L11_23, u1_L11_24, u1_L11_25, u1_L11_26, u1_L11_27, u1_L11_28, u1_L11_29, u1_L11_3, u1_L11_30, 
        u1_L11_31, u1_L11_32, u1_L11_4, u1_L11_5, u1_L11_6, u1_L11_7, u1_L11_8, u1_L11_9, u1_L12_1, 
        u1_L12_10, u1_L12_11, u1_L12_12, u1_L12_13, u1_L12_14, u1_L12_15, u1_L12_16, u1_L12_17, u1_L12_18, 
        u1_L12_19, u1_L12_2, u1_L12_20, u1_L12_21, u1_L12_22, u1_L12_23, u1_L12_24, u1_L12_25, u1_L12_26, 
        u1_L12_27, u1_L12_28, u1_L12_29, u1_L12_3, u1_L12_30, u1_L12_31, u1_L12_32, u1_L12_4, u1_L12_5, 
        u1_L12_6, u1_L12_7, u1_L12_8, u1_L12_9, u1_L13_1, u1_L13_10, u1_L13_11, u1_L13_12, u1_L13_13, 
        u1_L13_14, u1_L13_15, u1_L13_16, u1_L13_17, u1_L13_18, u1_L13_19, u1_L13_2, u1_L13_20, u1_L13_21, 
        u1_L13_22, u1_L13_23, u1_L13_24, u1_L13_25, u1_L13_26, u1_L13_27, u1_L13_28, u1_L13_29, u1_L13_3, 
        u1_L13_30, u1_L13_31, u1_L13_32, u1_L13_4, u1_L13_5, u1_L13_6, u1_L13_7, u1_L13_8, u1_L13_9, 
        u1_L14_1, u1_L14_10, u1_L14_11, u1_L14_12, u1_L14_13, u1_L14_14, u1_L14_15, u1_L14_16, u1_L14_17, 
        u1_L14_18, u1_L14_19, u1_L14_2, u1_L14_20, u1_L14_21, u1_L14_22, u1_L14_23, u1_L14_24, u1_L14_25, 
        u1_L14_26, u1_L14_27, u1_L14_28, u1_L14_29, u1_L14_3, u1_L14_30, u1_L14_31, u1_L14_32, u1_L14_4, 
        u1_L14_5, u1_L14_6, u1_L14_7, u1_L14_8, u1_L14_9, u1_L1_1, u1_L1_10, u1_L1_11, u1_L1_12, 
        u1_L1_13, u1_L1_14, u1_L1_15, u1_L1_16, u1_L1_17, u1_L1_18, u1_L1_19, u1_L1_2, u1_L1_20, 
        u1_L1_21, u1_L1_22, u1_L1_23, u1_L1_24, u1_L1_25, u1_L1_26, u1_L1_27, u1_L1_28, u1_L1_29, 
        u1_L1_3, u1_L1_30, u1_L1_31, u1_L1_32, u1_L1_4, u1_L1_5, u1_L1_6, u1_L1_7, u1_L1_8, 
        u1_L1_9, u1_L2_1, u1_L2_10, u1_L2_11, u1_L2_12, u1_L2_13, u1_L2_14, u1_L2_15, u1_L2_16, 
        u1_L2_17, u1_L2_18, u1_L2_19, u1_L2_2, u1_L2_20, u1_L2_21, u1_L2_22, u1_L2_23, u1_L2_24, 
        u1_L2_25, u1_L2_26, u1_L2_27, u1_L2_28, u1_L2_29, u1_L2_3, u1_L2_30, u1_L2_31, u1_L2_32, 
        u1_L2_4, u1_L2_5, u1_L2_6, u1_L2_7, u1_L2_8, u1_L2_9, u1_L3_1, u1_L3_10, u1_L3_11, 
        u1_L3_12, u1_L3_13, u1_L3_14, u1_L3_15, u1_L3_16, u1_L3_17, u1_L3_18, u1_L3_19, u1_L3_2, 
        u1_L3_20, u1_L3_21, u1_L3_22, u1_L3_23, u1_L3_24, u1_L3_25, u1_L3_26, u1_L3_27, u1_L3_28, 
        u1_L3_29, u1_L3_3, u1_L3_30, u1_L3_31, u1_L3_32, u1_L3_4, u1_L3_5, u1_L3_6, u1_L3_7, 
        u1_L3_8, u1_L3_9, u1_L4_1, u1_L4_10, u1_L4_11, u1_L4_12, u1_L4_13, u1_L4_14, u1_L4_15, 
        u1_L4_16, u1_L4_17, u1_L4_18, u1_L4_19, u1_L4_2, u1_L4_20, u1_L4_21, u1_L4_22, u1_L4_23, 
        u1_L4_24, u1_L4_25, u1_L4_26, u1_L4_27, u1_L4_28, u1_L4_29, u1_L4_3, u1_L4_30, u1_L4_31, 
        u1_L4_32, u1_L4_4, u1_L4_5, u1_L4_6, u1_L4_7, u1_L4_8, u1_L4_9, u1_L5_1, u1_L5_10, 
        u1_L5_11, u1_L5_12, u1_L5_13, u1_L5_14, u1_L5_15, u1_L5_16, u1_L5_17, u1_L5_18, u1_L5_19, 
        u1_L5_2, u1_L5_20, u1_L5_21, u1_L5_22, u1_L5_23, u1_L5_24, u1_L5_25, u1_L5_26, u1_L5_27, 
        u1_L5_28, u1_L5_29, u1_L5_3, u1_L5_30, u1_L5_31, u1_L5_32, u1_L5_4, u1_L5_5, u1_L5_6, 
        u1_L5_7, u1_L5_8, u1_L5_9, u1_L6_1, u1_L6_10, u1_L6_11, u1_L6_12, u1_L6_13, u1_L6_14, 
        u1_L6_15, u1_L6_16, u1_L6_17, u1_L6_18, u1_L6_19, u1_L6_2, u1_L6_20, u1_L6_21, u1_L6_22, 
        u1_L6_23, u1_L6_24, u1_L6_25, u1_L6_26, u1_L6_27, u1_L6_28, u1_L6_29, u1_L6_3, u1_L6_30, 
        u1_L6_31, u1_L6_32, u1_L6_4, u1_L6_5, u1_L6_6, u1_L6_7, u1_L6_8, u1_L6_9, u1_L7_1, 
        u1_L7_10, u1_L7_11, u1_L7_12, u1_L7_13, u1_L7_14, u1_L7_15, u1_L7_16, u1_L7_17, u1_L7_18, 
        u1_L7_19, u1_L7_2, u1_L7_20, u1_L7_21, u1_L7_22, u1_L7_23, u1_L7_24, u1_L7_25, u1_L7_26, 
        u1_L7_27, u1_L7_28, u1_L7_29, u1_L7_3, u1_L7_30, u1_L7_31, u1_L7_32, u1_L7_4, u1_L7_5, 
        u1_L7_6, u1_L7_7, u1_L7_8, u1_L7_9, u1_L8_1, u1_L8_10, u1_L8_11, u1_L8_12, u1_L8_13, 
        u1_L8_14, u1_L8_15, u1_L8_16, u1_L8_17, u1_L8_18, u1_L8_19, u1_L8_2, u1_L8_20, u1_L8_21, 
        u1_L8_22, u1_L8_23, u1_L8_24, u1_L8_25, u1_L8_26, u1_L8_27, u1_L8_28, u1_L8_29, u1_L8_3, 
        u1_L8_30, u1_L8_31, u1_L8_32, u1_L8_4, u1_L8_5, u1_L8_6, u1_L8_7, u1_L8_8, u1_L8_9, 
        u1_L9_1, u1_L9_10, u1_L9_11, u1_L9_12, u1_L9_13, u1_L9_14, u1_L9_15, u1_L9_16, u1_L9_17, 
        u1_L9_18, u1_L9_19, u1_L9_2, u1_L9_20, u1_L9_21, u1_L9_22, u1_L9_23, u1_L9_24, u1_L9_25, 
        u1_L9_26, u1_L9_27, u1_L9_28, u1_L9_29, u1_L9_3, u1_L9_30, u1_L9_31, u1_L9_32, u1_L9_4, 
        u1_L9_5, u1_L9_6, u1_L9_7, u1_L9_8, u1_L9_9, u1_R0_1, u1_R0_10, u1_R0_11, u1_R0_12, 
        u1_R0_13, u1_R0_14, u1_R0_15, u1_R0_16, u1_R0_17, u1_R0_18, u1_R0_19, u1_R0_2, u1_R0_20, 
        u1_R0_21, u1_R0_22, u1_R0_23, u1_R0_24, u1_R0_25, u1_R0_26, u1_R0_27, u1_R0_28, u1_R0_29, 
        u1_R0_3, u1_R0_30, u1_R0_31, u1_R0_32, u1_R0_4, u1_R0_5, u1_R0_6, u1_R0_7, u1_R0_8, 
        u1_R0_9, u1_R10_1, u1_R10_10, u1_R10_11, u1_R10_12, u1_R10_13, u1_R10_14, u1_R10_15, u1_R10_16, 
        u1_R10_17, u1_R10_18, u1_R10_19, u1_R10_2, u1_R10_20, u1_R10_21, u1_R10_22, u1_R10_23, u1_R10_24, 
        u1_R10_25, u1_R10_26, u1_R10_27, u1_R10_28, u1_R10_29, u1_R10_3, u1_R10_30, u1_R10_31, u1_R10_32, 
        u1_R10_4, u1_R10_5, u1_R10_6, u1_R10_7, u1_R10_8, u1_R10_9, u1_R11_1, u1_R11_10, u1_R11_11, 
        u1_R11_12, u1_R11_13, u1_R11_14, u1_R11_15, u1_R11_16, u1_R11_17, u1_R11_18, u1_R11_19, u1_R11_2, 
        u1_R11_20, u1_R11_21, u1_R11_22, u1_R11_23, u1_R11_24, u1_R11_25, u1_R11_26, u1_R11_27, u1_R11_28, 
        u1_R11_29, u1_R11_3, u1_R11_30, u1_R11_31, u1_R11_32, u1_R11_4, u1_R11_5, u1_R11_6, u1_R11_7, 
        u1_R11_8, u1_R11_9, u1_R12_1, u1_R12_10, u1_R12_11, u1_R12_12, u1_R12_13, u1_R12_14, u1_R12_15, 
        u1_R12_16, u1_R12_17, u1_R12_18, u1_R12_19, u1_R12_2, u1_R12_20, u1_R12_21, u1_R12_22, u1_R12_23, 
        u1_R12_24, u1_R12_25, u1_R12_26, u1_R12_27, u1_R12_28, u1_R12_29, u1_R12_3, u1_R12_30, u1_R12_31, 
        u1_R12_32, u1_R12_4, u1_R12_5, u1_R12_6, u1_R12_7, u1_R12_8, u1_R12_9, u1_R13_1, u1_R13_10, 
        u1_R13_11, u1_R13_12, u1_R13_13, u1_R13_14, u1_R13_15, u1_R13_16, u1_R13_17, u1_R13_18, u1_R13_19, 
        u1_R13_2, u1_R13_20, u1_R13_21, u1_R13_22, u1_R13_23, u1_R13_24, u1_R13_25, u1_R13_26, u1_R13_27, 
        u1_R13_28, u1_R13_29, u1_R13_3, u1_R13_30, u1_R13_31, u1_R13_32, u1_R13_4, u1_R13_5, u1_R13_6, 
        u1_R13_7, u1_R13_8, u1_R13_9, u1_R1_1, u1_R1_10, u1_R1_11, u1_R1_12, u1_R1_13, u1_R1_14, 
        u1_R1_15, u1_R1_16, u1_R1_17, u1_R1_18, u1_R1_19, u1_R1_2, u1_R1_20, u1_R1_21, u1_R1_22, 
        u1_R1_23, u1_R1_24, u1_R1_25, u1_R1_26, u1_R1_27, u1_R1_28, u1_R1_29, u1_R1_3, u1_R1_30, 
        u1_R1_31, u1_R1_32, u1_R1_4, u1_R1_5, u1_R1_6, u1_R1_7, u1_R1_8, u1_R1_9, u1_R2_1, 
        u1_R2_10, u1_R2_11, u1_R2_12, u1_R2_13, u1_R2_14, u1_R2_15, u1_R2_16, u1_R2_17, u1_R2_18, 
        u1_R2_19, u1_R2_2, u1_R2_20, u1_R2_21, u1_R2_22, u1_R2_23, u1_R2_24, u1_R2_25, u1_R2_26, 
        u1_R2_27, u1_R2_28, u1_R2_29, u1_R2_3, u1_R2_30, u1_R2_31, u1_R2_32, u1_R2_4, u1_R2_5, 
        u1_R2_6, u1_R2_7, u1_R2_8, u1_R2_9, u1_R3_1, u1_R3_10, u1_R3_11, u1_R3_12, u1_R3_13, 
        u1_R3_14, u1_R3_15, u1_R3_16, u1_R3_17, u1_R3_18, u1_R3_19, u1_R3_2, u1_R3_20, u1_R3_21, 
        u1_R3_22, u1_R3_23, u1_R3_24, u1_R3_25, u1_R3_26, u1_R3_27, u1_R3_28, u1_R3_29, u1_R3_3, 
        u1_R3_30, u1_R3_31, u1_R3_32, u1_R3_4, u1_R3_5, u1_R3_6, u1_R3_7, u1_R3_8, u1_R3_9, 
        u1_R4_1, u1_R4_10, u1_R4_11, u1_R4_12, u1_R4_13, u1_R4_14, u1_R4_15, u1_R4_16, u1_R4_17, 
        u1_R4_18, u1_R4_19, u1_R4_2, u1_R4_20, u1_R4_21, u1_R4_22, u1_R4_23, u1_R4_24, u1_R4_25, 
        u1_R4_26, u1_R4_27, u1_R4_28, u1_R4_29, u1_R4_3, u1_R4_30, u1_R4_31, u1_R4_32, u1_R4_4, 
        u1_R4_5, u1_R4_6, u1_R4_7, u1_R4_8, u1_R4_9, u1_R5_1, u1_R5_10, u1_R5_11, u1_R5_12, 
        u1_R5_13, u1_R5_14, u1_R5_15, u1_R5_16, u1_R5_17, u1_R5_18, u1_R5_19, u1_R5_2, u1_R5_20, 
        u1_R5_21, u1_R5_22, u1_R5_23, u1_R5_24, u1_R5_25, u1_R5_26, u1_R5_27, u1_R5_28, u1_R5_29, 
        u1_R5_3, u1_R5_30, u1_R5_31, u1_R5_32, u1_R5_4, u1_R5_5, u1_R5_6, u1_R5_7, u1_R5_8, 
        u1_R5_9, u1_R6_1, u1_R6_10, u1_R6_11, u1_R6_12, u1_R6_13, u1_R6_14, u1_R6_15, u1_R6_16, 
        u1_R6_17, u1_R6_18, u1_R6_19, u1_R6_2, u1_R6_20, u1_R6_21, u1_R6_22, u1_R6_23, u1_R6_24, 
        u1_R6_25, u1_R6_26, u1_R6_27, u1_R6_28, u1_R6_29, u1_R6_3, u1_R6_30, u1_R6_31, u1_R6_32, 
        u1_R6_4, u1_R6_5, u1_R6_6, u1_R6_7, u1_R6_8, u1_R6_9, u1_R7_1, u1_R7_10, u1_R7_11, 
        u1_R7_12, u1_R7_13, u1_R7_14, u1_R7_15, u1_R7_16, u1_R7_17, u1_R7_18, u1_R7_19, u1_R7_2, 
        u1_R7_20, u1_R7_21, u1_R7_22, u1_R7_23, u1_R7_24, u1_R7_25, u1_R7_26, u1_R7_27, u1_R7_28, 
        u1_R7_29, u1_R7_3, u1_R7_30, u1_R7_31, u1_R7_32, u1_R7_4, u1_R7_5, u1_R7_6, u1_R7_7, 
        u1_R7_8, u1_R7_9, u1_R8_1, u1_R8_10, u1_R8_11, u1_R8_12, u1_R8_13, u1_R8_14, u1_R8_15, 
        u1_R8_16, u1_R8_17, u1_R8_18, u1_R8_19, u1_R8_2, u1_R8_20, u1_R8_21, u1_R8_22, u1_R8_23, 
        u1_R8_24, u1_R8_25, u1_R8_26, u1_R8_27, u1_R8_28, u1_R8_29, u1_R8_3, u1_R8_30, u1_R8_31, 
        u1_R8_32, u1_R8_4, u1_R8_5, u1_R8_6, u1_R8_7, u1_R8_8, u1_R8_9, u1_R9_1, u1_R9_10, 
        u1_R9_11, u1_R9_12, u1_R9_13, u1_R9_14, u1_R9_15, u1_R9_16, u1_R9_17, u1_R9_18, u1_R9_19, 
        u1_R9_2, u1_R9_20, u1_R9_21, u1_R9_22, u1_R9_23, u1_R9_24, u1_R9_25, u1_R9_26, u1_R9_27, 
        u1_R9_28, u1_R9_29, u1_R9_3, u1_R9_30, u1_R9_31, u1_R9_32, u1_R9_4, u1_R9_5, u1_R9_6, 
        u1_R9_7, u1_R9_8, u1_R9_9, u1_desIn_r_0, u1_desIn_r_1, u1_desIn_r_10, u1_desIn_r_11, u1_desIn_r_12, u1_desIn_r_13, 
        u1_desIn_r_14, u1_desIn_r_15, u1_desIn_r_16, u1_desIn_r_17, u1_desIn_r_18, u1_desIn_r_19, u1_desIn_r_2, u1_desIn_r_20, u1_desIn_r_21, 
        u1_desIn_r_22, u1_desIn_r_23, u1_desIn_r_24, u1_desIn_r_25, u1_desIn_r_26, u1_desIn_r_27, u1_desIn_r_28, u1_desIn_r_29, u1_desIn_r_3, 
        u1_desIn_r_30, u1_desIn_r_31, u1_desIn_r_32, u1_desIn_r_33, u1_desIn_r_34, u1_desIn_r_35, u1_desIn_r_36, u1_desIn_r_37, u1_desIn_r_38, 
        u1_desIn_r_39, u1_desIn_r_4, u1_desIn_r_40, u1_desIn_r_41, u1_desIn_r_42, u1_desIn_r_43, u1_desIn_r_44, u1_desIn_r_45, u1_desIn_r_46, 
        u1_desIn_r_47, u1_desIn_r_48, u1_desIn_r_49, u1_desIn_r_5, u1_desIn_r_50, u1_desIn_r_51, u1_desIn_r_52, u1_desIn_r_53, u1_desIn_r_54, 
        u1_desIn_r_55, u1_desIn_r_56, u1_desIn_r_57, u1_desIn_r_58, u1_desIn_r_59, u1_desIn_r_6, u1_desIn_r_60, u1_desIn_r_61, u1_desIn_r_62, 
        u1_desIn_r_63, u1_desIn_r_7, u1_desIn_r_8, u1_desIn_r_9, u1_key_r_0, u1_key_r_1, u1_key_r_10, u1_key_r_11, u1_key_r_12, 
        u1_key_r_13, u1_key_r_14, u1_key_r_15, u1_key_r_16, u1_key_r_17, u1_key_r_18, u1_key_r_19, u1_key_r_2, u1_key_r_20, 
        u1_key_r_21, u1_key_r_22, u1_key_r_23, u1_key_r_24, u1_key_r_25, u1_key_r_26, u1_key_r_27, u1_key_r_28, u1_key_r_29, 
        u1_key_r_3, u1_key_r_30, u1_key_r_31, u1_key_r_32, u1_key_r_33, u1_key_r_34, u1_key_r_35, u1_key_r_36, u1_key_r_37, 
        u1_key_r_38, u1_key_r_39, u1_key_r_4, u1_key_r_40, u1_key_r_41, u1_key_r_42, u1_key_r_43, u1_key_r_44, u1_key_r_45, 
        u1_key_r_46, u1_key_r_47, u1_key_r_48, u1_key_r_49, u1_key_r_5, u1_key_r_50, u1_key_r_51, u1_key_r_52, u1_key_r_53, 
        u1_key_r_54, u1_key_r_55, u1_key_r_6, u1_key_r_7, u1_key_r_8, u1_key_r_9, u1_uk_K_r0_11, u1_uk_K_r0_13, u1_uk_K_r0_15, 
        u1_uk_K_r0_17, u1_uk_K_r0_19, u1_uk_K_r0_2, u1_uk_K_r0_22, u1_uk_K_r0_25, u1_uk_K_r0_28, u1_uk_K_r0_31, u1_uk_K_r0_32, u1_uk_K_r0_34, 
        u1_uk_K_r0_36, u1_uk_K_r0_47, u1_uk_K_r0_49, u1_uk_K_r0_52, u1_uk_K_r0_55, u1_uk_K_r0_7, u1_uk_K_r10_10, u1_uk_K_r10_11, u1_uk_K_r10_14, 
        u1_uk_K_r10_16, u1_uk_K_r10_18, u1_uk_K_r10_19, u1_uk_K_r10_23, u1_uk_K_r10_25, u1_uk_K_r10_27, u1_uk_K_r10_28, u1_uk_K_r10_32, u1_uk_K_r10_34, 
        u1_uk_K_r10_37, u1_uk_K_r10_39, u1_uk_K_r10_4, u1_uk_K_r10_41, u1_uk_K_r10_42, u1_uk_K_r10_43, u1_uk_K_r10_44, u1_uk_K_r10_47, u1_uk_K_r10_48, 
        u1_uk_K_r10_49, u1_uk_K_r10_52, u1_uk_K_r10_9, u1_uk_K_r11_10, u1_uk_K_r11_11, u1_uk_K_r11_17, u1_uk_K_r11_19, u1_uk_K_r11_20, u1_uk_K_r11_21, 
        u1_uk_K_r11_24, u1_uk_K_r11_25, u1_uk_K_r11_26, u1_uk_K_r11_27, u1_uk_K_r11_28, u1_uk_K_r11_29, u1_uk_K_r11_33, u1_uk_K_r11_34, u1_uk_K_r11_39, 
        u1_uk_K_r11_4, u1_uk_K_r11_46, u1_uk_K_r11_47, u1_uk_K_r11_48, u1_uk_K_r11_5, u1_uk_K_r11_53, u1_uk_K_r11_54, u1_uk_K_r11_6, u1_uk_K_r11_7, 
        u1_uk_K_r11_8, u1_uk_K_r12_1, u1_uk_K_r12_10, u1_uk_K_r12_15, u1_uk_K_r12_16, u1_uk_K_r12_18, u1_uk_K_r12_21, u1_uk_K_r12_22, u1_uk_K_r12_25, 
        u1_uk_K_r12_30, u1_uk_K_r12_33, u1_uk_K_r12_36, u1_uk_K_r12_41, u1_uk_K_r12_42, u1_uk_K_r12_44, u1_uk_K_r12_47, u1_uk_K_r12_7, u1_uk_K_r13_0, 
        u1_uk_K_r13_13, u1_uk_K_r13_17, u1_uk_K_r13_19, u1_uk_K_r13_2, u1_uk_K_r13_22, u1_uk_K_r13_23, u1_uk_K_r13_25, u1_uk_K_r13_31, u1_uk_K_r13_32, 
        u1_uk_K_r13_35, u1_uk_K_r13_36, u1_uk_K_r13_38, u1_uk_K_r13_4, u1_uk_K_r13_44, u1_uk_K_r13_55, u1_uk_K_r14_10, u1_uk_K_r14_11, u1_uk_K_r14_12, 
        u1_uk_K_r14_15, u1_uk_K_r14_16, u1_uk_K_r14_18, u1_uk_K_r14_2, u1_uk_K_r14_23, u1_uk_K_r14_3, u1_uk_K_r14_38, u1_uk_K_r14_39, u1_uk_K_r14_42, 
        u1_uk_K_r14_43, u1_uk_K_r14_45, u1_uk_K_r14_46, u1_uk_K_r14_5, u1_uk_K_r14_50, u1_uk_K_r14_8, u1_uk_K_r14_9, u1_uk_K_r1_10, u1_uk_K_r1_15, 
        u1_uk_K_r1_16, u1_uk_K_r1_17, u1_uk_K_r1_18, u1_uk_K_r1_21, u1_uk_K_r1_22, u1_uk_K_r1_33, u1_uk_K_r1_36, u1_uk_K_r1_41, u1_uk_K_r1_42, 
        u1_uk_K_r1_44, u1_uk_K_r1_47, u1_uk_K_r1_6, u1_uk_K_r1_7, u1_uk_K_r2_13, u1_uk_K_r2_16, u1_uk_K_r2_18, u1_uk_K_r2_20, u1_uk_K_r2_21, 
        u1_uk_K_r2_24, u1_uk_K_r2_25, u1_uk_K_r2_26, u1_uk_K_r2_27, u1_uk_K_r2_28, u1_uk_K_r2_29, u1_uk_K_r2_31, u1_uk_K_r2_33, u1_uk_K_r2_36, 
        u1_uk_K_r2_4, u1_uk_K_r2_41, u1_uk_K_r2_46, u1_uk_K_r2_47, u1_uk_K_r2_49, u1_uk_K_r2_50, u1_uk_K_r2_53, u1_uk_K_r2_55, u1_uk_K_r2_6, 
        u1_uk_K_r2_7, u1_uk_K_r3_10, u1_uk_K_r3_11, u1_uk_K_r3_14, u1_uk_K_r3_15, u1_uk_K_r3_16, u1_uk_K_r3_19, u1_uk_K_r3_24, u1_uk_K_r3_29, 
        u1_uk_K_r3_33, u1_uk_K_r3_34, u1_uk_K_r3_35, u1_uk_K_r3_38, u1_uk_K_r3_4, u1_uk_K_r3_43, u1_uk_K_r3_44, u1_uk_K_r3_47, u1_uk_K_r3_51, 
        u1_uk_K_r3_52, u1_uk_K_r3_9, u1_uk_K_r4_0, u1_uk_K_r4_11, u1_uk_K_r4_17, u1_uk_K_r4_18, u1_uk_K_r4_23, u1_uk_K_r4_27, u1_uk_K_r4_3, 
        u1_uk_K_r4_31, u1_uk_K_r4_33, u1_uk_K_r4_35, u1_uk_K_r4_38, u1_uk_K_r4_4, u1_uk_K_r4_41, u1_uk_K_r4_47, u1_uk_K_r4_48, u1_uk_K_r4_49, 
        u1_uk_K_r4_5, u1_uk_K_r4_54, u1_uk_K_r4_55, u1_uk_K_r5_0, u1_uk_K_r5_1, u1_uk_K_r5_10, u1_uk_K_r5_13, u1_uk_K_r5_16, u1_uk_K_r5_17, 
        u1_uk_K_r5_18, u1_uk_K_r5_19, u1_uk_K_r5_21, u1_uk_K_r5_23, u1_uk_K_r5_26, u1_uk_K_r5_31, u1_uk_K_r5_32, u1_uk_K_r5_35, u1_uk_K_r5_36, 
        u1_uk_K_r5_37, u1_uk_K_r5_39, u1_uk_K_r5_4, u1_uk_K_r5_40, u1_uk_K_r5_41, u1_uk_K_r5_43, u1_uk_K_r5_48, u1_uk_K_r5_5, u1_uk_K_r5_51, 
        u1_uk_K_r5_53, u1_uk_K_r5_7, u1_uk_K_r5_8, u1_uk_K_r6_0, u1_uk_K_r6_10, u1_uk_K_r6_14, u1_uk_K_r6_17, u1_uk_K_r6_19, u1_uk_K_r6_21, 
        u1_uk_K_r6_22, u1_uk_K_r6_26, u1_uk_K_r6_27, u1_uk_K_r6_28, u1_uk_K_r6_29, u1_uk_K_r6_3, u1_uk_K_r6_30, u1_uk_K_r6_31, u1_uk_K_r6_34, 
        u1_uk_K_r6_35, u1_uk_K_r6_37, u1_uk_K_r6_46, u1_uk_K_r6_51, u1_uk_K_r6_53, u1_uk_K_r6_55, u1_uk_K_r6_7, u1_uk_K_r7_0, u1_uk_K_r7_1, 
        u1_uk_K_r7_13, u1_uk_K_r7_15, u1_uk_K_r7_16, u1_uk_K_r7_2, u1_uk_K_r7_20, u1_uk_K_r7_22, u1_uk_K_r7_23, u1_uk_K_r7_24, u1_uk_K_r7_25, 
        u1_uk_K_r7_26, u1_uk_K_r7_27, u1_uk_K_r7_29, u1_uk_K_r7_30, u1_uk_K_r7_31, u1_uk_K_r7_32, u1_uk_K_r7_34, u1_uk_K_r7_37, u1_uk_K_r7_39, 
        u1_uk_K_r7_41, u1_uk_K_r7_46, u1_uk_K_r7_48, u1_uk_K_r7_5, u1_uk_K_r7_53, u1_uk_K_r7_55, u1_uk_K_r7_6, u1_uk_K_r7_7, u1_uk_K_r7_8, 
        u1_uk_K_r7_9, u1_uk_K_r8_10, u1_uk_K_r8_13, u1_uk_K_r8_16, u1_uk_K_r8_17, u1_uk_K_r8_19, u1_uk_K_r8_2, u1_uk_K_r8_21, u1_uk_K_r8_22, 
        u1_uk_K_r8_27, u1_uk_K_r8_28, u1_uk_K_r8_32, u1_uk_K_r8_37, u1_uk_K_r8_39, u1_uk_K_r8_40, u1_uk_K_r8_41, u1_uk_K_r8_42, u1_uk_K_r8_43, 
        u1_uk_K_r8_44, u1_uk_K_r8_48, u1_uk_K_r8_5, u1_uk_K_r8_51, u1_uk_K_r8_52, u1_uk_K_r8_8, u1_uk_K_r9_0, u1_uk_K_r9_1, u1_uk_K_r9_10, 
        u1_uk_K_r9_12, u1_uk_K_r9_13, u1_uk_K_r9_15, u1_uk_K_r9_18, u1_uk_K_r9_19, u1_uk_K_r9_22, u1_uk_K_r9_23, u1_uk_K_r9_25, u1_uk_K_r9_27, 
        u1_uk_K_r9_30, u1_uk_K_r9_31, u1_uk_K_r9_33, u1_uk_K_r9_35, u1_uk_K_r9_38, u1_uk_K_r9_4, u1_uk_K_r9_45, u1_uk_K_r9_48, u1_uk_K_r9_49, 
        u1_uk_K_r9_5, u1_uk_K_r9_54, u1_uk_K_r9_55, u1_uk_K_r9_6, u1_uk_K_r9_7, u1_uk_K_r9_9, u1_uk_n1218, u1_uk_n1219, u1_uk_n1220, 
        u1_uk_n1221, u1_uk_n1222, u1_uk_n1224, u1_uk_n1225, u1_uk_n1227, u1_uk_n1228, u1_uk_n1229, u1_uk_n1230, u1_uk_n1231, 
        u1_uk_n1233, u1_uk_n1234, u1_uk_n1235, u1_uk_n1236, u1_uk_n1237, u1_uk_n1238, u1_uk_n1239, u1_uk_n1240, u1_uk_n1241, 
        u1_uk_n1242, u1_uk_n1243, u1_uk_n1244, u1_uk_n1245, u1_uk_n1246, u1_uk_n1247, u1_uk_n1248, u1_uk_n1249, u1_uk_n1250, 
        u1_uk_n1251, u1_uk_n1252, u1_uk_n1253, u1_uk_n1255, u1_uk_n1256, u1_uk_n1257, u1_uk_n1258, u1_uk_n1259, u1_uk_n1260, 
        u1_uk_n1261, u1_uk_n1262, u1_uk_n1263, u1_uk_n1264, u1_uk_n1265, u1_uk_n1266, u1_uk_n1267, u1_uk_n1268, u1_uk_n1269, 
        u1_uk_n1270, u1_uk_n1271, u1_uk_n1272, u1_uk_n1273, u1_uk_n1274, u1_uk_n1275, u1_uk_n1276, u1_uk_n1277, u1_uk_n1278, 
        u1_uk_n1279, u1_uk_n1281, u1_uk_n1282, u1_uk_n1284, u1_uk_n1286, u1_uk_n1288, u1_uk_n1289, u1_uk_n1290, u1_uk_n1291, 
        u1_uk_n1292, u1_uk_n1293, u1_uk_n1294, u1_uk_n1295, u1_uk_n1296, u1_uk_n1297, u1_uk_n1299, u1_uk_n1300, u1_uk_n1303, 
        u1_uk_n1304, u1_uk_n1305, u1_uk_n1307, u1_uk_n1308, u1_uk_n1309, u1_uk_n1310, u1_uk_n1311, u1_uk_n1312, u1_uk_n1313, 
        u1_uk_n1314, u1_uk_n1315, u1_uk_n1316, u1_uk_n1317, u1_uk_n1318, u1_uk_n1319, u1_uk_n1320, u1_uk_n1321, u1_uk_n1322, 
        u1_uk_n1323, u1_uk_n1324, u1_uk_n1325, u1_uk_n1326, u1_uk_n1327, u1_uk_n1328, u1_uk_n1329, u1_uk_n1330, u1_uk_n1331, 
        u1_uk_n1332, u1_uk_n1333, u1_uk_n1334, u1_uk_n1335, u1_uk_n1336, u1_uk_n1338, u1_uk_n1339, u1_uk_n1340, u1_uk_n1341, 
        u1_uk_n1342, u1_uk_n1343, u1_uk_n1344, u1_uk_n1345, u1_uk_n1346, u1_uk_n1347, u1_uk_n1348, u1_uk_n1349, u1_uk_n1350, 
        u1_uk_n1351, u1_uk_n1352, u1_uk_n1353, u1_uk_n1354, u1_uk_n1355, u1_uk_n1356, u1_uk_n1357, u1_uk_n1358, u1_uk_n1359, 
        u1_uk_n1360, u1_uk_n1361, u1_uk_n1363, u1_uk_n1365, u1_uk_n1366, u1_uk_n1367, u1_uk_n1369, u1_uk_n1371, u1_uk_n1372, 
        u1_uk_n1374, u1_uk_n1375, u1_uk_n1376, u1_uk_n1377, u1_uk_n1378, u1_uk_n1380, u1_uk_n1381, u1_uk_n1382, u1_uk_n1383, 
        u1_uk_n1386, u1_uk_n1389, u1_uk_n1390, u1_uk_n1391, u1_uk_n1393, u1_uk_n1394, u1_uk_n1395, u1_uk_n1396, u1_uk_n1397, 
        u1_uk_n1398, u1_uk_n1399, u1_uk_n1400, u1_uk_n1401, u1_uk_n1402, u1_uk_n1403, u1_uk_n1404, u1_uk_n1405, u1_uk_n1406, 
        u1_uk_n1407, u1_uk_n1408, u1_uk_n1409, u1_uk_n1410, u1_uk_n1411, u1_uk_n1412, u1_uk_n1413, u1_uk_n1414, u1_uk_n1415, 
        u1_uk_n1417, u1_uk_n1418, u1_uk_n1419, u1_uk_n1422, u1_uk_n1423, u1_uk_n1424, u1_uk_n1425, u1_uk_n1426, u1_uk_n1427, 
        u1_uk_n1429, u1_uk_n1430, u1_uk_n1431, u1_uk_n1433, u1_uk_n1435, u1_uk_n1436, u1_uk_n1437, u1_uk_n1438, u1_uk_n1439, 
        u1_uk_n1440, u1_uk_n1441, u1_uk_n1442, u1_uk_n1443, u1_uk_n1444, u1_uk_n1446, u1_uk_n1447, u1_uk_n1448, u1_uk_n1449, 
        u1_uk_n1450, u1_uk_n1452, u1_uk_n1453, u1_uk_n1454, u1_uk_n1455, u1_uk_n1456, u1_uk_n1457, u1_uk_n1458, u1_uk_n1459, 
        u1_uk_n1460, u1_uk_n1461, u1_uk_n1462, u1_uk_n1463, u1_uk_n1464, u1_uk_n1465, u1_uk_n1466, u1_uk_n1468, u1_uk_n1469, 
        u1_uk_n1470, u1_uk_n1471, u1_uk_n1472, u1_uk_n1474, u1_uk_n1475, u1_uk_n1476, u1_uk_n1477, u1_uk_n1478, u1_uk_n1482, 
        u1_uk_n1483, u1_uk_n1484, u1_uk_n1485, u1_uk_n1486, u1_uk_n1487, u1_uk_n1488, u1_uk_n1489, u1_uk_n1490, u1_uk_n1491, 
        u1_uk_n1492, u1_uk_n1494, u1_uk_n1495, u1_uk_n1496, u1_uk_n1498, u1_uk_n1499, u1_uk_n1500, u1_uk_n1501, u1_uk_n1504, 
        u1_uk_n1505, u1_uk_n1507, u1_uk_n1508, u1_uk_n1510, u1_uk_n1514, u1_uk_n1516, u1_uk_n1517, u1_uk_n1518, u1_uk_n1520, 
        u1_uk_n1521, u1_uk_n1523, u1_uk_n1524, u1_uk_n1526, u1_uk_n1527, u1_uk_n1528, u1_uk_n1529, u1_uk_n1530, u1_uk_n1531, 
        u1_uk_n1532, u1_uk_n1533, u1_uk_n1534, u1_uk_n1536, u1_uk_n1537, u1_uk_n1538, u1_uk_n1540, u1_uk_n1541, u1_uk_n1543, 
        u1_uk_n1544, u1_uk_n1545, u1_uk_n1547, u1_uk_n1548, u1_uk_n1549, u1_uk_n1551, u1_uk_n1552, u1_uk_n1554, u1_uk_n1555, 
        u1_uk_n1556, u1_uk_n1557, u1_uk_n1558, u1_uk_n1559, u1_uk_n1560, u1_uk_n1561, u1_uk_n1562, u1_uk_n1563, u1_uk_n1564, 
        u1_uk_n1565, u1_uk_n1566, u1_uk_n1567, u1_uk_n1568, u1_uk_n1570, u1_uk_n1571, u1_uk_n1572, u1_uk_n1573, u1_uk_n1574, 
        u1_uk_n1577, u1_uk_n1578, u1_uk_n1579, u1_uk_n1581, u1_uk_n1584, u1_uk_n1585, u1_uk_n1586, u1_uk_n1588, u1_uk_n1592, 
        u1_uk_n1593, u1_uk_n1595, u1_uk_n1598, u1_uk_n1599, u1_uk_n1600, u1_uk_n1601, u1_uk_n1603, u1_uk_n1604, u1_uk_n1605, 
        u1_uk_n1606, u1_uk_n1607, u1_uk_n1608, u1_uk_n1610, u1_uk_n1612, u1_uk_n1613, u1_uk_n1614, u1_uk_n1615, u1_uk_n1616, 
        u1_uk_n1618, u1_uk_n1619, u1_uk_n1620, u1_uk_n1621, u1_uk_n1622, u1_uk_n1623, u1_uk_n1624, u1_uk_n1625, u1_uk_n1626, 
        u1_uk_n1627, u1_uk_n1628, u1_uk_n1629, u1_uk_n1630, u1_uk_n1632, u1_uk_n1633, u1_uk_n1634, u1_uk_n1635, u1_uk_n1639, 
        u1_uk_n1640, u1_uk_n1641, u1_uk_n1642, u1_uk_n1643, u1_uk_n1644, u1_uk_n1645, u1_uk_n1647, u1_uk_n1649, u1_uk_n1651, 
        u1_uk_n1652, u1_uk_n1653, u1_uk_n1654, u1_uk_n1655, u1_uk_n1656, u1_uk_n1659, u1_uk_n1660, u1_uk_n1661, u1_uk_n1662, 
        u1_uk_n1663, u1_uk_n1664, u1_uk_n1667, u1_uk_n1669, u1_uk_n1670, u1_uk_n1672, u1_uk_n1673, u1_uk_n1676, u1_uk_n1677, 
        u1_uk_n1678, u1_uk_n1682, u1_uk_n1683, u1_uk_n1684, u1_uk_n1687, u1_uk_n1688, u1_uk_n1689, u1_uk_n1690, u1_uk_n1691, 
        u1_uk_n1692, u1_uk_n1693, u1_uk_n1694, u1_uk_n1695, u1_uk_n1696, u1_uk_n1698, u1_uk_n1699, u1_uk_n1702, u1_uk_n1703, 
        u1_uk_n1704, u1_uk_n1705, u1_uk_n1707, u1_uk_n1708, u1_uk_n1709, u1_uk_n1710, u1_uk_n1711, u1_uk_n1712, u1_uk_n1713, 
        u1_uk_n1714, u1_uk_n1715, u1_uk_n1716, u1_uk_n1717, u1_uk_n1718, u1_uk_n1719, u1_uk_n1720, u1_uk_n1721, u1_uk_n1722, 
        u1_uk_n1723, u1_uk_n1728, u1_uk_n1729, u1_uk_n1730, u1_uk_n1731, u1_uk_n1732, u1_uk_n1734, u1_uk_n1735, u1_uk_n1736, 
        u1_uk_n1737, u1_uk_n1738, u1_uk_n1739, u1_uk_n1744, u1_uk_n1745, u1_uk_n1748, u1_uk_n1749, u1_uk_n1750, u1_uk_n1751, 
        u1_uk_n1752, u1_uk_n1753, u1_uk_n1754, u1_uk_n1755, u1_uk_n1756, u1_uk_n1757, u1_uk_n1758, u1_uk_n1761, u1_uk_n1762, 
        u1_uk_n1763, u1_uk_n1764, u1_uk_n1765, u1_uk_n1766, u1_uk_n1767, u1_uk_n1768, u1_uk_n1769, u1_uk_n1772, u1_uk_n1773, 
        u1_uk_n1774, u1_uk_n1775, u1_uk_n1776, u1_uk_n1777, u1_uk_n1780, u1_uk_n1781, u1_uk_n1782, u1_uk_n1783, u1_uk_n1784, 
        u1_uk_n1785, u1_uk_n1787, u1_uk_n1790, u1_uk_n1791, u1_uk_n1792, u1_uk_n1793, u1_uk_n1797, u1_uk_n1798, u1_uk_n1799, 
        u1_uk_n1800, u1_uk_n1801, u1_uk_n1802, u1_uk_n1803, u1_uk_n1804, u1_uk_n1806, u1_uk_n1807, u1_uk_n1808, u1_uk_n1809, 
        u1_uk_n1810, u1_uk_n1811, u1_uk_n1812, u1_uk_n1813, u1_uk_n1814, u1_uk_n1815, u1_uk_n1816, u1_uk_n1817, u1_uk_n1818, 
        u1_uk_n1819, u1_uk_n1820, u1_uk_n1821, u1_uk_n1822, u1_uk_n1823, u1_uk_n1824, u1_uk_n1826, u1_uk_n1827, u1_uk_n1829, 
        u1_uk_n1830, u1_uk_n1831, u1_uk_n1832, u1_uk_n1833, u1_uk_n1834, u1_uk_n1835, u1_uk_n1836, u1_uk_n1837, u1_uk_n1838, 
        u1_uk_n1839, u1_uk_n1840, u1_uk_n1841, u1_uk_n1842, u1_uk_n1843, u1_uk_n1844, u1_uk_n1845, u1_uk_n1846, u1_uk_n1847, 
        u1_uk_n1848, u1_uk_n1849, u1_uk_n1850, u1_uk_n1851, u1_uk_n1852, u1_uk_n1853, u1_uk_n1854, u1_uk_n1855, u1_uk_n1856, 
        u1_uk_n1858, u1_uk_n1859, u1_uk_n1860, u1_uk_n1862, u1_uk_n1863, u1_uk_n1864, u1_uk_n1865, u1_uk_n1866, u1_uk_n1867, 
        u1_uk_n1868, u1_uk_n1869, u1_uk_n1870, u1_uk_n1872, u1_uk_n1873, u1_uk_n1874, u1_uk_n1875, u1_uk_n1876, u1_uk_n1879, 
        u1_uk_n1880, u1_uk_n1881, u1_uk_n1882, u1_uk_n1883, u1_uk_n1884, u1_uk_n1885, u1_uk_n1886, u1_uk_n1887, u2_FP_33, 
        u2_FP_34, u2_FP_35, u2_FP_36, u2_FP_37, u2_FP_38, u2_FP_39, u2_FP_40, u2_FP_41, u2_FP_42, 
        u2_FP_43, u2_FP_44, u2_FP_45, u2_FP_46, u2_FP_47, u2_FP_48, u2_FP_49, u2_FP_50, u2_FP_51, 
        u2_FP_52, u2_FP_53, u2_FP_54, u2_FP_55, u2_FP_56, u2_FP_57, u2_FP_58, u2_FP_59, u2_FP_60, 
        u2_FP_61, u2_FP_62, u2_FP_63, u2_FP_64, u2_K10_10, u2_K10_11, u2_K10_15, u2_K10_17, u2_K10_25, 
        u2_K10_26, u2_K10_30, u2_K10_32, u2_K10_34, u2_K10_36, u2_K10_4, u2_K10_42, u2_K10_43, u2_K10_44, 
        u2_K10_46, u2_K10_6, u2_K11_11, u2_K11_13, u2_K11_16, u2_K11_18, u2_K11_21, u2_K11_29, u2_K11_38, 
        u2_K11_4, u2_K11_42, u2_K11_45, u2_K11_48, u2_K11_6, u2_K11_7, u2_K11_9, u2_K12_2, u2_K12_20, 
        u2_K12_22, u2_K12_24, u2_K12_25, u2_K12_26, u2_K12_27, u2_K12_29, u2_K12_34, u2_K12_37, u2_K12_41, 
        u2_K12_46, u2_K12_47, u2_K12_8, u2_K13_14, u2_K13_20, u2_K13_26, u2_K13_3, u2_K13_31, u2_K13_32, 
        u2_K13_34, u2_K13_37, u2_K13_40, u2_K13_42, u2_K13_44, u2_K13_45, u2_K13_46, u2_K13_47, u2_K13_8, 
        u2_K14_10, u2_K14_11, u2_K14_12, u2_K14_13, u2_K14_14, u2_K14_16, u2_K14_17, u2_K14_18, u2_K14_21, 
        u2_K14_25, u2_K14_28, u2_K14_3, u2_K14_39, u2_K14_42, u2_K14_6, u2_K14_8, u2_K15_1, u2_K15_13, 
        u2_K15_16, u2_K15_18, u2_K15_2, u2_K15_20, u2_K15_21, u2_K15_23, u2_K15_28, u2_K15_29, u2_K15_31, 
        u2_K15_34, u2_K15_35, u2_K15_39, u2_K15_5, u2_K16_26, u2_K16_31, u2_K16_42, u2_K16_44, u2_K16_47, 
        u2_K16_5, u2_K16_6, u2_K16_8, u2_K16_9, u2_K1_15, u2_K1_16, u2_K1_19, u2_K1_24, u2_K1_28, 
        u2_K1_37, u2_K1_40, u2_K1_43, u2_K1_45, u2_K1_46, u2_K1_5, u2_K1_9, u2_K2_1, u2_K2_16, 
        u2_K2_18, u2_K2_20, u2_K2_34, u2_K2_35, u2_K2_36, u2_K2_40, u2_K2_43, u2_K2_44, u2_K2_45, 
        u2_K2_46, u2_K2_47, u2_K2_48, u2_K3_13, u2_K3_15, u2_K3_16, u2_K3_20, u2_K3_23, u2_K3_30, 
        u2_K3_32, u2_K3_35, u2_K3_42, u2_K3_43, u2_K3_47, u2_K3_48, u2_K3_7, u2_K4_14, u2_K4_21, 
        u2_K4_22, u2_K4_27, u2_K4_33, u2_K4_34, u2_K4_35, u2_K4_38, u2_K4_39, u2_K4_42, u2_K4_6, 
        u2_K4_7, u2_K5_1, u2_K5_10, u2_K5_11, u2_K5_13, u2_K5_14, u2_K5_16, u2_K5_17, u2_K5_18, 
        u2_K5_19, u2_K5_21, u2_K5_23, u2_K5_24, u2_K5_25, u2_K5_26, u2_K5_28, u2_K5_3, u2_K5_31, 
        u2_K5_32, u2_K5_34, u2_K5_38, u2_K5_41, u2_K5_44, u2_K5_47, u2_K5_48, u2_K5_5, u2_K5_6, 
        u2_K5_8, u2_K5_9, u2_K6_1, u2_K6_11, u2_K6_13, u2_K6_14, u2_K6_15, u2_K6_16, u2_K6_20, 
        u2_K6_22, u2_K6_24, u2_K6_25, u2_K6_27, u2_K6_3, u2_K6_32, u2_K6_34, u2_K6_36, u2_K6_40, 
        u2_K7_26, u2_K7_3, u2_K7_31, u2_K7_33, u2_K7_35, u2_K7_37, u2_K7_38, u2_K7_4, u2_K7_43, 
        u2_K7_45, u2_K7_48, u2_K7_5, u2_K7_7, u2_K8_18, u2_K8_24, u2_K8_26, u2_K8_31, u2_K8_41, 
        u2_K8_45, u2_K8_5, u2_K8_8, u2_K9_15, u2_K9_23, u2_K9_25, u2_K9_28, u2_K9_29, u2_K9_3, 
        u2_K9_32, u2_K9_36, u2_K9_38, u2_K9_40, u2_K9_45, u2_K9_5, u2_L0_1, u2_L0_10, u2_L0_11, 
        u2_L0_12, u2_L0_13, u2_L0_14, u2_L0_15, u2_L0_16, u2_L0_17, u2_L0_18, u2_L0_19, u2_L0_2, 
        u2_L0_20, u2_L0_21, u2_L0_22, u2_L0_23, u2_L0_24, u2_L0_25, u2_L0_26, u2_L0_27, u2_L0_28, 
        u2_L0_29, u2_L0_3, u2_L0_30, u2_L0_31, u2_L0_32, u2_L0_4, u2_L0_5, u2_L0_6, u2_L0_7, 
        u2_L0_8, u2_L0_9, u2_L10_1, u2_L10_10, u2_L10_11, u2_L10_12, u2_L10_13, u2_L10_14, u2_L10_15, 
        u2_L10_16, u2_L10_17, u2_L10_18, u2_L10_19, u2_L10_2, u2_L10_20, u2_L10_21, u2_L10_22, u2_L10_23, 
        u2_L10_24, u2_L10_25, u2_L10_26, u2_L10_27, u2_L10_28, u2_L10_29, u2_L10_3, u2_L10_30, u2_L10_31, 
        u2_L10_32, u2_L10_4, u2_L10_5, u2_L10_6, u2_L10_7, u2_L10_8, u2_L10_9, u2_L11_1, u2_L11_10, 
        u2_L11_11, u2_L11_12, u2_L11_13, u2_L11_14, u2_L11_15, u2_L11_16, u2_L11_17, u2_L11_18, u2_L11_19, 
        u2_L11_2, u2_L11_20, u2_L11_21, u2_L11_22, u2_L11_23, u2_L11_24, u2_L11_25, u2_L11_26, u2_L11_27, 
        u2_L11_28, u2_L11_29, u2_L11_3, u2_L11_30, u2_L11_31, u2_L11_32, u2_L11_4, u2_L11_5, u2_L11_6, 
        u2_L11_7, u2_L11_8, u2_L11_9, u2_L12_1, u2_L12_10, u2_L12_11, u2_L12_12, u2_L12_13, u2_L12_14, 
        u2_L12_15, u2_L12_16, u2_L12_17, u2_L12_18, u2_L12_19, u2_L12_2, u2_L12_20, u2_L12_21, u2_L12_22, 
        u2_L12_23, u2_L12_24, u2_L12_25, u2_L12_26, u2_L12_27, u2_L12_28, u2_L12_29, u2_L12_3, u2_L12_30, 
        u2_L12_31, u2_L12_32, u2_L12_4, u2_L12_5, u2_L12_6, u2_L12_7, u2_L12_8, u2_L12_9, u2_L13_1, 
        u2_L13_10, u2_L13_11, u2_L13_12, u2_L13_13, u2_L13_14, u2_L13_15, u2_L13_16, u2_L13_17, u2_L13_18, 
        u2_L13_19, u2_L13_2, u2_L13_20, u2_L13_21, u2_L13_22, u2_L13_23, u2_L13_24, u2_L13_25, u2_L13_26, 
        u2_L13_27, u2_L13_28, u2_L13_29, u2_L13_3, u2_L13_30, u2_L13_31, u2_L13_32, u2_L13_4, u2_L13_5, 
        u2_L13_6, u2_L13_7, u2_L13_8, u2_L13_9, u2_L14_1, u2_L14_10, u2_L14_11, u2_L14_12, u2_L14_13, 
        u2_L14_14, u2_L14_15, u2_L14_16, u2_L14_17, u2_L14_18, u2_L14_19, u2_L14_2, u2_L14_20, u2_L14_21, 
        u2_L14_22, u2_L14_23, u2_L14_24, u2_L14_25, u2_L14_26, u2_L14_27, u2_L14_28, u2_L14_29, u2_L14_3, 
        u2_L14_30, u2_L14_31, u2_L14_32, u2_L14_4, u2_L14_5, u2_L14_6, u2_L14_7, u2_L14_8, u2_L14_9, 
        u2_L1_1, u2_L1_10, u2_L1_11, u2_L1_12, u2_L1_13, u2_L1_14, u2_L1_15, u2_L1_16, u2_L1_17, 
        u2_L1_18, u2_L1_19, u2_L1_2, u2_L1_20, u2_L1_21, u2_L1_22, u2_L1_23, u2_L1_24, u2_L1_25, 
        u2_L1_26, u2_L1_27, u2_L1_28, u2_L1_29, u2_L1_3, u2_L1_30, u2_L1_31, u2_L1_32, u2_L1_4, 
        u2_L1_5, u2_L1_6, u2_L1_7, u2_L1_8, u2_L1_9, u2_L2_1, u2_L2_10, u2_L2_11, u2_L2_12, 
        u2_L2_13, u2_L2_14, u2_L2_15, u2_L2_16, u2_L2_17, u2_L2_18, u2_L2_19, u2_L2_2, u2_L2_20, 
        u2_L2_21, u2_L2_22, u2_L2_23, u2_L2_24, u2_L2_25, u2_L2_26, u2_L2_27, u2_L2_28, u2_L2_29, 
        u2_L2_3, u2_L2_30, u2_L2_31, u2_L2_32, u2_L2_4, u2_L2_5, u2_L2_6, u2_L2_7, u2_L2_8, 
        u2_L2_9, u2_L3_1, u2_L3_10, u2_L3_11, u2_L3_12, u2_L3_13, u2_L3_14, u2_L3_15, u2_L3_16, 
        u2_L3_17, u2_L3_18, u2_L3_19, u2_L3_2, u2_L3_20, u2_L3_21, u2_L3_22, u2_L3_23, u2_L3_24, 
        u2_L3_25, u2_L3_26, u2_L3_27, u2_L3_28, u2_L3_29, u2_L3_3, u2_L3_30, u2_L3_31, u2_L3_32, 
        u2_L3_4, u2_L3_5, u2_L3_6, u2_L3_7, u2_L3_8, u2_L3_9, u2_L4_1, u2_L4_10, u2_L4_11, 
        u2_L4_12, u2_L4_13, u2_L4_14, u2_L4_15, u2_L4_16, u2_L4_17, u2_L4_18, u2_L4_19, u2_L4_2, 
        u2_L4_20, u2_L4_21, u2_L4_22, u2_L4_23, u2_L4_24, u2_L4_25, u2_L4_26, u2_L4_27, u2_L4_28, 
        u2_L4_29, u2_L4_3, u2_L4_30, u2_L4_31, u2_L4_32, u2_L4_4, u2_L4_5, u2_L4_6, u2_L4_7, 
        u2_L4_8, u2_L4_9, u2_L5_1, u2_L5_10, u2_L5_11, u2_L5_12, u2_L5_13, u2_L5_14, u2_L5_15, 
        u2_L5_16, u2_L5_17, u2_L5_18, u2_L5_19, u2_L5_2, u2_L5_20, u2_L5_21, u2_L5_22, u2_L5_23, 
        u2_L5_24, u2_L5_25, u2_L5_26, u2_L5_27, u2_L5_28, u2_L5_29, u2_L5_3, u2_L5_30, u2_L5_31, 
        u2_L5_32, u2_L5_4, u2_L5_5, u2_L5_6, u2_L5_7, u2_L5_8, u2_L5_9, u2_L6_1, u2_L6_10, 
        u2_L6_11, u2_L6_12, u2_L6_13, u2_L6_14, u2_L6_15, u2_L6_16, u2_L6_17, u2_L6_18, u2_L6_19, 
        u2_L6_2, u2_L6_20, u2_L6_21, u2_L6_22, u2_L6_23, u2_L6_24, u2_L6_25, u2_L6_26, u2_L6_27, 
        u2_L6_28, u2_L6_29, u2_L6_3, u2_L6_30, u2_L6_31, u2_L6_32, u2_L6_4, u2_L6_5, u2_L6_6, 
        u2_L6_7, u2_L6_8, u2_L6_9, u2_L7_1, u2_L7_10, u2_L7_11, u2_L7_12, u2_L7_13, u2_L7_14, 
        u2_L7_15, u2_L7_16, u2_L7_17, u2_L7_18, u2_L7_19, u2_L7_2, u2_L7_20, u2_L7_21, u2_L7_22, 
        u2_L7_23, u2_L7_24, u2_L7_25, u2_L7_26, u2_L7_27, u2_L7_28, u2_L7_29, u2_L7_3, u2_L7_30, 
        u2_L7_31, u2_L7_32, u2_L7_4, u2_L7_5, u2_L7_6, u2_L7_7, u2_L7_8, u2_L7_9, u2_L8_1, 
        u2_L8_10, u2_L8_11, u2_L8_12, u2_L8_13, u2_L8_14, u2_L8_15, u2_L8_16, u2_L8_17, u2_L8_18, 
        u2_L8_19, u2_L8_2, u2_L8_20, u2_L8_21, u2_L8_22, u2_L8_23, u2_L8_24, u2_L8_25, u2_L8_26, 
        u2_L8_27, u2_L8_28, u2_L8_29, u2_L8_3, u2_L8_30, u2_L8_31, u2_L8_32, u2_L8_4, u2_L8_5, 
        u2_L8_6, u2_L8_7, u2_L8_8, u2_L8_9, u2_L9_1, u2_L9_10, u2_L9_11, u2_L9_12, u2_L9_13, 
        u2_L9_14, u2_L9_15, u2_L9_16, u2_L9_17, u2_L9_18, u2_L9_19, u2_L9_2, u2_L9_20, u2_L9_21, 
        u2_L9_22, u2_L9_23, u2_L9_24, u2_L9_25, u2_L9_26, u2_L9_27, u2_L9_28, u2_L9_29, u2_L9_3, 
        u2_L9_30, u2_L9_31, u2_L9_32, u2_L9_4, u2_L9_5, u2_L9_6, u2_L9_7, u2_L9_8, u2_L9_9, 
        u2_R0_1, u2_R0_10, u2_R0_11, u2_R0_12, u2_R0_13, u2_R0_14, u2_R0_15, u2_R0_16, u2_R0_17, 
        u2_R0_18, u2_R0_19, u2_R0_2, u2_R0_20, u2_R0_21, u2_R0_22, u2_R0_23, u2_R0_24, u2_R0_25, 
        u2_R0_26, u2_R0_27, u2_R0_28, u2_R0_29, u2_R0_3, u2_R0_30, u2_R0_31, u2_R0_32, u2_R0_4, 
        u2_R0_5, u2_R0_6, u2_R0_7, u2_R0_8, u2_R0_9, u2_R10_1, u2_R10_10, u2_R10_11, u2_R10_12, 
        u2_R10_13, u2_R10_14, u2_R10_15, u2_R10_16, u2_R10_17, u2_R10_18, u2_R10_19, u2_R10_2, u2_R10_20, 
        u2_R10_21, u2_R10_22, u2_R10_23, u2_R10_24, u2_R10_25, u2_R10_26, u2_R10_27, u2_R10_28, u2_R10_29, 
        u2_R10_3, u2_R10_30, u2_R10_31, u2_R10_32, u2_R10_4, u2_R10_5, u2_R10_6, u2_R10_7, u2_R10_8, 
        u2_R10_9, u2_R11_1, u2_R11_10, u2_R11_11, u2_R11_12, u2_R11_13, u2_R11_14, u2_R11_15, u2_R11_16, 
        u2_R11_17, u2_R11_18, u2_R11_19, u2_R11_2, u2_R11_20, u2_R11_21, u2_R11_22, u2_R11_23, u2_R11_24, 
        u2_R11_25, u2_R11_26, u2_R11_27, u2_R11_28, u2_R11_29, u2_R11_3, u2_R11_30, u2_R11_31, u2_R11_32, 
        u2_R11_4, u2_R11_5, u2_R11_6, u2_R11_7, u2_R11_8, u2_R11_9, u2_R12_1, u2_R12_10, u2_R12_11, 
        u2_R12_12, u2_R12_13, u2_R12_14, u2_R12_15, u2_R12_16, u2_R12_17, u2_R12_18, u2_R12_19, u2_R12_2, 
        u2_R12_20, u2_R12_21, u2_R12_22, u2_R12_23, u2_R12_24, u2_R12_25, u2_R12_26, u2_R12_27, u2_R12_28, 
        u2_R12_29, u2_R12_3, u2_R12_30, u2_R12_31, u2_R12_32, u2_R12_4, u2_R12_5, u2_R12_6, u2_R12_7, 
        u2_R12_8, u2_R12_9, u2_R13_1, u2_R13_10, u2_R13_11, u2_R13_12, u2_R13_13, u2_R13_14, u2_R13_15, 
        u2_R13_16, u2_R13_17, u2_R13_18, u2_R13_19, u2_R13_2, u2_R13_20, u2_R13_21, u2_R13_22, u2_R13_23, 
        u2_R13_24, u2_R13_25, u2_R13_26, u2_R13_27, u2_R13_28, u2_R13_29, u2_R13_3, u2_R13_30, u2_R13_31, 
        u2_R13_32, u2_R13_4, u2_R13_5, u2_R13_6, u2_R13_7, u2_R13_8, u2_R13_9, u2_R1_1, u2_R1_10, 
        u2_R1_11, u2_R1_12, u2_R1_13, u2_R1_14, u2_R1_15, u2_R1_16, u2_R1_17, u2_R1_18, u2_R1_19, 
        u2_R1_2, u2_R1_20, u2_R1_21, u2_R1_22, u2_R1_23, u2_R1_24, u2_R1_25, u2_R1_26, u2_R1_27, 
        u2_R1_28, u2_R1_29, u2_R1_3, u2_R1_30, u2_R1_31, u2_R1_32, u2_R1_4, u2_R1_5, u2_R1_6, 
        u2_R1_7, u2_R1_8, u2_R1_9, u2_R2_1, u2_R2_10, u2_R2_11, u2_R2_12, u2_R2_13, u2_R2_14, 
        u2_R2_15, u2_R2_16, u2_R2_17, u2_R2_18, u2_R2_19, u2_R2_2, u2_R2_20, u2_R2_21, u2_R2_22, 
        u2_R2_23, u2_R2_24, u2_R2_25, u2_R2_26, u2_R2_27, u2_R2_28, u2_R2_29, u2_R2_3, u2_R2_30, 
        u2_R2_31, u2_R2_32, u2_R2_4, u2_R2_5, u2_R2_6, u2_R2_7, u2_R2_8, u2_R2_9, u2_R3_1, 
        u2_R3_10, u2_R3_11, u2_R3_12, u2_R3_13, u2_R3_14, u2_R3_15, u2_R3_16, u2_R3_17, u2_R3_18, 
        u2_R3_19, u2_R3_2, u2_R3_20, u2_R3_21, u2_R3_22, u2_R3_23, u2_R3_24, u2_R3_25, u2_R3_26, 
        u2_R3_27, u2_R3_28, u2_R3_29, u2_R3_3, u2_R3_30, u2_R3_31, u2_R3_32, u2_R3_4, u2_R3_5, 
        u2_R3_6, u2_R3_7, u2_R3_8, u2_R3_9, u2_R4_1, u2_R4_10, u2_R4_11, u2_R4_12, u2_R4_13, 
        u2_R4_14, u2_R4_15, u2_R4_16, u2_R4_17, u2_R4_18, u2_R4_19, u2_R4_2, u2_R4_20, u2_R4_21, 
        u2_R4_22, u2_R4_23, u2_R4_24, u2_R4_25, u2_R4_26, u2_R4_27, u2_R4_28, u2_R4_29, u2_R4_3, 
        u2_R4_30, u2_R4_31, u2_R4_32, u2_R4_4, u2_R4_5, u2_R4_6, u2_R4_7, u2_R4_8, u2_R4_9, 
        u2_R5_1, u2_R5_10, u2_R5_11, u2_R5_12, u2_R5_13, u2_R5_14, u2_R5_15, u2_R5_16, u2_R5_17, 
        u2_R5_18, u2_R5_19, u2_R5_2, u2_R5_20, u2_R5_21, u2_R5_22, u2_R5_23, u2_R5_24, u2_R5_25, 
        u2_R5_26, u2_R5_27, u2_R5_28, u2_R5_29, u2_R5_3, u2_R5_30, u2_R5_31, u2_R5_32, u2_R5_4, 
        u2_R5_5, u2_R5_6, u2_R5_7, u2_R5_8, u2_R5_9, u2_R6_1, u2_R6_10, u2_R6_11, u2_R6_12, 
        u2_R6_13, u2_R6_14, u2_R6_15, u2_R6_16, u2_R6_17, u2_R6_18, u2_R6_19, u2_R6_2, u2_R6_20, 
        u2_R6_21, u2_R6_22, u2_R6_23, u2_R6_24, u2_R6_25, u2_R6_26, u2_R6_27, u2_R6_28, u2_R6_29, 
        u2_R6_3, u2_R6_30, u2_R6_31, u2_R6_32, u2_R6_4, u2_R6_5, u2_R6_6, u2_R6_7, u2_R6_8, 
        u2_R6_9, u2_R7_1, u2_R7_10, u2_R7_11, u2_R7_12, u2_R7_13, u2_R7_14, u2_R7_15, u2_R7_16, 
        u2_R7_17, u2_R7_18, u2_R7_19, u2_R7_2, u2_R7_20, u2_R7_21, u2_R7_22, u2_R7_23, u2_R7_24, 
        u2_R7_25, u2_R7_26, u2_R7_27, u2_R7_28, u2_R7_29, u2_R7_3, u2_R7_30, u2_R7_31, u2_R7_32, 
        u2_R7_4, u2_R7_5, u2_R7_6, u2_R7_7, u2_R7_8, u2_R7_9, u2_R8_1, u2_R8_10, u2_R8_11, 
        u2_R8_12, u2_R8_13, u2_R8_14, u2_R8_15, u2_R8_16, u2_R8_17, u2_R8_18, u2_R8_19, u2_R8_2, 
        u2_R8_20, u2_R8_21, u2_R8_22, u2_R8_23, u2_R8_24, u2_R8_25, u2_R8_26, u2_R8_27, u2_R8_28, 
        u2_R8_29, u2_R8_3, u2_R8_30, u2_R8_31, u2_R8_32, u2_R8_4, u2_R8_5, u2_R8_6, u2_R8_7, 
        u2_R8_8, u2_R8_9, u2_R9_1, u2_R9_10, u2_R9_11, u2_R9_12, u2_R9_13, u2_R9_14, u2_R9_15, 
        u2_R9_16, u2_R9_17, u2_R9_18, u2_R9_19, u2_R9_2, u2_R9_20, u2_R9_21, u2_R9_22, u2_R9_23, 
        u2_R9_24, u2_R9_25, u2_R9_26, u2_R9_27, u2_R9_28, u2_R9_29, u2_R9_3, u2_R9_30, u2_R9_31, 
        u2_R9_32, u2_R9_4, u2_R9_5, u2_R9_6, u2_R9_7, u2_R9_8, u2_R9_9, u2_desIn_r_0, u2_desIn_r_1, 
        u2_desIn_r_10, u2_desIn_r_11, u2_desIn_r_12, u2_desIn_r_13, u2_desIn_r_14, u2_desIn_r_15, u2_desIn_r_16, u2_desIn_r_17, u2_desIn_r_18, 
        u2_desIn_r_19, u2_desIn_r_2, u2_desIn_r_20, u2_desIn_r_21, u2_desIn_r_22, u2_desIn_r_23, u2_desIn_r_24, u2_desIn_r_25, u2_desIn_r_26, 
        u2_desIn_r_27, u2_desIn_r_28, u2_desIn_r_29, u2_desIn_r_3, u2_desIn_r_30, u2_desIn_r_31, u2_desIn_r_32, u2_desIn_r_33, u2_desIn_r_34, 
        u2_desIn_r_35, u2_desIn_r_36, u2_desIn_r_37, u2_desIn_r_38, u2_desIn_r_39, u2_desIn_r_4, u2_desIn_r_40, u2_desIn_r_41, u2_desIn_r_42, 
        u2_desIn_r_43, u2_desIn_r_44, u2_desIn_r_45, u2_desIn_r_46, u2_desIn_r_47, u2_desIn_r_48, u2_desIn_r_49, u2_desIn_r_5, u2_desIn_r_50, 
        u2_desIn_r_51, u2_desIn_r_52, u2_desIn_r_53, u2_desIn_r_54, u2_desIn_r_55, u2_desIn_r_56, u2_desIn_r_57, u2_desIn_r_58, u2_desIn_r_59, 
        u2_desIn_r_6, u2_desIn_r_60, u2_desIn_r_61, u2_desIn_r_62, u2_desIn_r_63, u2_desIn_r_7, u2_desIn_r_8, u2_desIn_r_9, u2_key_r_0, 
        u2_key_r_1, u2_key_r_10, u2_key_r_11, u2_key_r_12, u2_key_r_13, u2_key_r_14, u2_key_r_16, u2_key_r_17, u2_key_r_19, 
        u2_key_r_2, u2_key_r_20, u2_key_r_21, u2_key_r_22, u2_key_r_23, u2_key_r_24, u2_key_r_25, u2_key_r_26, u2_key_r_27, 
        u2_key_r_28, u2_key_r_29, u2_key_r_3, u2_key_r_30, u2_key_r_31, u2_key_r_32, u2_key_r_33, u2_key_r_34, u2_key_r_35, 
        u2_key_r_36, u2_key_r_37, u2_key_r_4, u2_key_r_40, u2_key_r_41, u2_key_r_42, u2_key_r_43, u2_key_r_44, u2_key_r_46, 
        u2_key_r_47, u2_key_r_48, u2_key_r_49, u2_key_r_50, u2_key_r_51, u2_key_r_52, u2_key_r_53, u2_key_r_54, u2_key_r_55, 
        u2_key_r_6, u2_key_r_7, u2_key_r_8, u2_key_r_9, u2_uk_K_r0_11, u2_uk_K_r0_13, u2_uk_K_r0_15, u2_uk_K_r0_17, u2_uk_K_r0_25, 
        u2_uk_K_r0_31, u2_uk_K_r0_32, u2_uk_K_r0_34, u2_uk_K_r0_36, u2_uk_K_r0_47, u2_uk_K_r0_49, u2_uk_K_r0_55, u2_uk_K_r10_10, u2_uk_K_r10_16, 
        u2_uk_K_r10_25, u2_uk_K_r10_27, u2_uk_K_r10_32, u2_uk_K_r10_34, u2_uk_K_r10_4, u2_uk_K_r10_41, u2_uk_K_r10_43, u2_uk_K_r10_44, u2_uk_K_r10_49, 
        u2_uk_K_r11_10, u2_uk_K_r11_11, u2_uk_K_r11_19, u2_uk_K_r11_20, u2_uk_K_r11_21, u2_uk_K_r11_24, u2_uk_K_r11_25, u2_uk_K_r11_26, u2_uk_K_r11_27, 
        u2_uk_K_r11_28, u2_uk_K_r11_29, u2_uk_K_r11_33, u2_uk_K_r11_39, u2_uk_K_r11_4, u2_uk_K_r11_47, u2_uk_K_r11_48, u2_uk_K_r11_53, u2_uk_K_r11_6, 
        u2_uk_K_r11_7, u2_uk_K_r12_1, u2_uk_K_r12_10, u2_uk_K_r12_15, u2_uk_K_r12_16, u2_uk_K_r12_25, u2_uk_K_r12_30, u2_uk_K_r12_33, u2_uk_K_r12_36, 
        u2_uk_K_r12_41, u2_uk_K_r12_42, u2_uk_K_r12_7, u2_uk_K_r13_0, u2_uk_K_r13_13, u2_uk_K_r13_17, u2_uk_K_r13_19, u2_uk_K_r13_22, u2_uk_K_r13_25, 
        u2_uk_K_r13_32, u2_uk_K_r13_38, u2_uk_K_r13_55, u2_uk_K_r14_10, u2_uk_K_r14_12, u2_uk_K_r14_15, u2_uk_K_r14_16, u2_uk_K_r14_18, u2_uk_K_r14_2, 
        u2_uk_K_r14_3, u2_uk_K_r14_45, u2_uk_K_r14_46, u2_uk_K_r14_5, u2_uk_K_r14_50, u2_uk_K_r14_9, u2_uk_K_r1_15, u2_uk_K_r1_16, u2_uk_K_r1_17, 
        u2_uk_K_r1_18, u2_uk_K_r1_21, u2_uk_K_r1_22, u2_uk_K_r1_41, u2_uk_K_r1_42, u2_uk_K_r1_44, u2_uk_K_r1_47, u2_uk_K_r1_7, u2_uk_K_r2_13, 
        u2_uk_K_r2_18, u2_uk_K_r2_21, u2_uk_K_r2_24, u2_uk_K_r2_25, u2_uk_K_r2_26, u2_uk_K_r2_27, u2_uk_K_r2_28, u2_uk_K_r2_31, u2_uk_K_r2_36, 
        u2_uk_K_r2_49, u2_uk_K_r2_50, u2_uk_K_r2_55, u2_uk_K_r2_6, u2_uk_K_r3_10, u2_uk_K_r3_11, u2_uk_K_r3_14, u2_uk_K_r3_15, u2_uk_K_r3_16, 
        u2_uk_K_r3_19, u2_uk_K_r3_29, u2_uk_K_r3_38, u2_uk_K_r3_4, u2_uk_K_r3_43, u2_uk_K_r3_52, u2_uk_K_r3_9, u2_uk_K_r4_0, u2_uk_K_r4_11, 
        u2_uk_K_r4_17, u2_uk_K_r4_3, u2_uk_K_r4_33, u2_uk_K_r4_35, u2_uk_K_r4_38, u2_uk_K_r4_4, u2_uk_K_r4_41, u2_uk_K_r4_47, u2_uk_K_r4_5, 
        u2_uk_K_r4_54, u2_uk_K_r4_55, u2_uk_K_r5_0, u2_uk_K_r5_1, u2_uk_K_r5_10, u2_uk_K_r5_16, u2_uk_K_r5_17, u2_uk_K_r5_18, u2_uk_K_r5_19, 
        u2_uk_K_r5_21, u2_uk_K_r5_23, u2_uk_K_r5_26, u2_uk_K_r5_31, u2_uk_K_r5_37, u2_uk_K_r5_39, u2_uk_K_r5_4, u2_uk_K_r5_40, u2_uk_K_r5_41, 
        u2_uk_K_r5_43, u2_uk_K_r5_48, u2_uk_K_r5_51, u2_uk_K_r5_7, u2_uk_K_r6_0, u2_uk_K_r6_10, u2_uk_K_r6_14, u2_uk_K_r6_26, u2_uk_K_r6_29, 
        u2_uk_K_r6_3, u2_uk_K_r6_31, u2_uk_K_r6_34, u2_uk_K_r6_37, u2_uk_K_r6_46, u2_uk_K_r6_51, u2_uk_K_r6_53, u2_uk_K_r6_7, u2_uk_K_r7_0, 
        u2_uk_K_r7_13, u2_uk_K_r7_16, u2_uk_K_r7_2, u2_uk_K_r7_20, u2_uk_K_r7_23, u2_uk_K_r7_25, u2_uk_K_r7_26, u2_uk_K_r7_31, u2_uk_K_r7_32, 
        u2_uk_K_r7_37, u2_uk_K_r7_39, u2_uk_K_r7_41, u2_uk_K_r7_46, u2_uk_K_r7_48, u2_uk_K_r7_55, u2_uk_K_r7_9, u2_uk_K_r8_13, u2_uk_K_r8_16, 
        u2_uk_K_r8_17, u2_uk_K_r8_19, u2_uk_K_r8_2, u2_uk_K_r8_21, u2_uk_K_r8_22, u2_uk_K_r8_27, u2_uk_K_r8_28, u2_uk_K_r8_32, u2_uk_K_r8_37, 
        u2_uk_K_r8_40, u2_uk_K_r8_41, u2_uk_K_r8_42, u2_uk_K_r8_43, u2_uk_K_r8_44, u2_uk_K_r8_48, u2_uk_K_r8_52, u2_uk_K_r8_8, u2_uk_K_r9_0, 
        u2_uk_K_r9_1, u2_uk_K_r9_10, u2_uk_K_r9_12, u2_uk_K_r9_13, u2_uk_K_r9_15, u2_uk_K_r9_18, u2_uk_K_r9_19, u2_uk_K_r9_23, u2_uk_K_r9_25, 
        u2_uk_K_r9_27, u2_uk_K_r9_31, u2_uk_K_r9_33, u2_uk_K_r9_4, u2_uk_K_r9_45, u2_uk_K_r9_48, u2_uk_K_r9_49, u2_uk_K_r9_5, u2_uk_K_r9_54, 
        u2_uk_K_r9_55, u2_uk_K_r9_9, u2_uk_n1001, u2_uk_n1007, u2_uk_n1011, u2_uk_n1018, u2_uk_n1022, u2_uk_n1024, u2_uk_n1027, 
        u2_uk_n1028, u2_uk_n1031, u2_uk_n1035, u2_uk_n1036, u2_uk_n1038, u2_uk_n1040, u2_uk_n1042, u2_uk_n1043, u2_uk_n1044, 
        u2_uk_n1046, u2_uk_n1049, u2_uk_n1061, u2_uk_n1063, u2_uk_n1069, u2_uk_n1070, u2_uk_n1073, u2_uk_n1074, u2_uk_n1077, 
        u2_uk_n1079, u2_uk_n1081, u2_uk_n1082, u2_uk_n1089, u2_uk_n1093, u2_uk_n1094, u2_uk_n1096, u2_uk_n1097, u2_uk_n1100, 
        u2_uk_n1104, u2_uk_n1105, u2_uk_n1107, u2_uk_n1112, u2_uk_n1113, u2_uk_n1116, u2_uk_n1119, u2_uk_n1120, u2_uk_n1121, 
        u2_uk_n1125, u2_uk_n1128, u2_uk_n1130, u2_uk_n1131, u2_uk_n1132, u2_uk_n1134, u2_uk_n1136, u2_uk_n1137, u2_uk_n1140, 
        u2_uk_n1141, u2_uk_n1188, u2_uk_n1189, u2_uk_n1190, u2_uk_n1194, u2_uk_n1195, u2_uk_n1197, u2_uk_n1198, u2_uk_n1199, 
        u2_uk_n1200, u2_uk_n1201, u2_uk_n1203, u2_uk_n1204, u2_uk_n1205, u2_uk_n1206, u2_uk_n1207, u2_uk_n1208, u2_uk_n1209, 
        u2_uk_n1210, u2_uk_n1212, u2_uk_n1213, u2_uk_n1214, u2_uk_n1215, u2_uk_n1216, u2_uk_n1217, u2_uk_n1218, u2_uk_n1219, 
        u2_uk_n1220, u2_uk_n1221, u2_uk_n1222, u2_uk_n1223, u2_uk_n1225, u2_uk_n1226, u2_uk_n1227, u2_uk_n1228, u2_uk_n1229, 
        u2_uk_n1230, u2_uk_n1231, u2_uk_n1232, u2_uk_n1233, u2_uk_n1234, u2_uk_n1236, u2_uk_n1237, u2_uk_n1238, u2_uk_n1239, 
        u2_uk_n1240, u2_uk_n1243, u2_uk_n1244, u2_uk_n1245, u2_uk_n1246, u2_uk_n1247, u2_uk_n1248, u2_uk_n1249, u2_uk_n1251, 
        u2_uk_n1252, u2_uk_n1254, u2_uk_n1258, u2_uk_n1259, u2_uk_n1260, u2_uk_n1261, u2_uk_n1264, u2_uk_n1265, u2_uk_n1266, 
        u2_uk_n1267, u2_uk_n1269, u2_uk_n1270, u2_uk_n1274, u2_uk_n1275, u2_uk_n1279, u2_uk_n1280, u2_uk_n1281, u2_uk_n1282, 
        u2_uk_n1283, u2_uk_n1284, u2_uk_n1285, u2_uk_n1286, u2_uk_n1287, u2_uk_n1288, u2_uk_n1290, u2_uk_n1291, u2_uk_n1292, 
        u2_uk_n1293, u2_uk_n1294, u2_uk_n1295, u2_uk_n1296, u2_uk_n1297, u2_uk_n1298, u2_uk_n1299, u2_uk_n1300, u2_uk_n1301, 
        u2_uk_n1302, u2_uk_n1303, u2_uk_n1305, u2_uk_n1306, u2_uk_n1308, u2_uk_n1309, u2_uk_n1310, u2_uk_n1311, u2_uk_n1312, 
        u2_uk_n1313, u2_uk_n1314, u2_uk_n1315, u2_uk_n1316, u2_uk_n1317, u2_uk_n1318, u2_uk_n1319, u2_uk_n1320, u2_uk_n1321, 
        u2_uk_n1322, u2_uk_n1323, u2_uk_n1324, u2_uk_n1325, u2_uk_n1326, u2_uk_n1328, u2_uk_n1329, u2_uk_n1330, u2_uk_n1331, 
        u2_uk_n1333, u2_uk_n1335, u2_uk_n1336, u2_uk_n1337, u2_uk_n1339, u2_uk_n1341, u2_uk_n1342, u2_uk_n1344, u2_uk_n1345, 
        u2_uk_n1346, u2_uk_n1347, u2_uk_n1348, u2_uk_n1350, u2_uk_n1351, u2_uk_n1352, u2_uk_n1353, u2_uk_n1356, u2_uk_n1359, 
        u2_uk_n1360, u2_uk_n1361, u2_uk_n1363, u2_uk_n1364, u2_uk_n1365, u2_uk_n1367, u2_uk_n1370, u2_uk_n1372, u2_uk_n1375, 
        u2_uk_n1376, u2_uk_n1377, u2_uk_n1378, u2_uk_n1379, u2_uk_n1381, u2_uk_n1382, u2_uk_n1383, u2_uk_n1395, u2_uk_n1396, 
        u2_uk_n1400, u2_uk_n1401, u2_uk_n1403, u2_uk_n1405, u2_uk_n1408, u2_uk_n1410, u2_uk_n1411, u2_uk_n1412, u2_uk_n1413, 
        u2_uk_n1414, u2_uk_n1416, u2_uk_n1418, u2_uk_n1419, u2_uk_n1420, u2_uk_n1422, u2_uk_n1424, u2_uk_n1425, u2_uk_n1426, 
        u2_uk_n1428, u2_uk_n1429, u2_uk_n1430, u2_uk_n1433, u2_uk_n1435, u2_uk_n1438, u2_uk_n1439, u2_uk_n1440, u2_uk_n1441, 
        u2_uk_n1442, u2_uk_n1444, u2_uk_n1445, u2_uk_n1446, u2_uk_n1447, u2_uk_n1448, u2_uk_n1452, u2_uk_n1453, u2_uk_n1454, 
        u2_uk_n1456, u2_uk_n1457, u2_uk_n1458, u2_uk_n1459, u2_uk_n1460, u2_uk_n1461, u2_uk_n1462, u2_uk_n1464, u2_uk_n1465, 
        u2_uk_n1466, u2_uk_n1468, u2_uk_n1470, u2_uk_n1471, u2_uk_n1475, u2_uk_n1480, u2_uk_n1486, u2_uk_n1487, u2_uk_n1488, 
        u2_uk_n1490, u2_uk_n1491, u2_uk_n1493, u2_uk_n1494, u2_uk_n1496, u2_uk_n1497, u2_uk_n1498, u2_uk_n1499, u2_uk_n1500, 
        u2_uk_n1501, u2_uk_n1502, u2_uk_n1503, u2_uk_n1504, u2_uk_n1506, u2_uk_n1507, u2_uk_n1508, u2_uk_n1510, u2_uk_n1511, 
        u2_uk_n1513, u2_uk_n1514, u2_uk_n1515, u2_uk_n1517, u2_uk_n1518, u2_uk_n1519, u2_uk_n1521, u2_uk_n1522, u2_uk_n1524, 
        u2_uk_n1525, u2_uk_n1526, u2_uk_n1527, u2_uk_n1528, u2_uk_n1529, u2_uk_n1530, u2_uk_n1531, u2_uk_n1532, u2_uk_n1533, 
        u2_uk_n1535, u2_uk_n1536, u2_uk_n1537, u2_uk_n1538, u2_uk_n1542, u2_uk_n1543, u2_uk_n1544, u2_uk_n1548, u2_uk_n1549, 
        u2_uk_n1551, u2_uk_n1555, u2_uk_n1556, u2_uk_n1558, u2_uk_n1563, u2_uk_n1565, u2_uk_n1568, u2_uk_n1570, u2_uk_n1571, 
        u2_uk_n1573, u2_uk_n1574, u2_uk_n1576, u2_uk_n1577, u2_uk_n1580, u2_uk_n1583, u2_uk_n1585, u2_uk_n1586, u2_uk_n1590, 
        u2_uk_n1591, u2_uk_n1592, u2_uk_n1594, u2_uk_n1595, u2_uk_n1597, u2_uk_n1598, u2_uk_n1599, u2_uk_n1600, u2_uk_n1602, 
        u2_uk_n1603, u2_uk_n1604, u2_uk_n1605, u2_uk_n1609, u2_uk_n1610, u2_uk_n1612, u2_uk_n1613, u2_uk_n1614, u2_uk_n1615, 
        u2_uk_n1617, u2_uk_n1622, u2_uk_n1623, u2_uk_n1624, u2_uk_n1625, u2_uk_n1626, u2_uk_n1629, u2_uk_n1630, u2_uk_n1631, 
        u2_uk_n1632, u2_uk_n1633, u2_uk_n1634, u2_uk_n1639, u2_uk_n1640, u2_uk_n1642, u2_uk_n1643, u2_uk_n1646, u2_uk_n1647, 
        u2_uk_n1652, u2_uk_n1653, u2_uk_n1654, u2_uk_n1657, u2_uk_n1658, u2_uk_n1659, u2_uk_n1660, u2_uk_n1661, u2_uk_n1664, 
        u2_uk_n1665, u2_uk_n1666, u2_uk_n1668, u2_uk_n1672, u2_uk_n1673, u2_uk_n1674, u2_uk_n1675, u2_uk_n1677, u2_uk_n1678, 
        u2_uk_n1680, u2_uk_n1681, u2_uk_n1682, u2_uk_n1683, u2_uk_n1684, u2_uk_n1685, u2_uk_n1687, u2_uk_n1688, u2_uk_n1689, 
        u2_uk_n1690, u2_uk_n1691, u2_uk_n1693, u2_uk_n1698, u2_uk_n1699, u2_uk_n1700, u2_uk_n1702, u2_uk_n1705, u2_uk_n1707, 
        u2_uk_n1708, u2_uk_n1709, u2_uk_n1715, u2_uk_n1718, u2_uk_n1720, u2_uk_n1721, u2_uk_n1722, u2_uk_n1723, u2_uk_n1724, 
        u2_uk_n1725, u2_uk_n1726, u2_uk_n1727, u2_uk_n1728, u2_uk_n1731, u2_uk_n1732, u2_uk_n1734, u2_uk_n1735, u2_uk_n1736, 
        u2_uk_n1737, u2_uk_n1738, u2_uk_n1742, u2_uk_n1743, u2_uk_n1744, u2_uk_n1745, u2_uk_n1746, u2_uk_n1747, u2_uk_n1750, 
        u2_uk_n1753, u2_uk_n1755, u2_uk_n1760, u2_uk_n1761, u2_uk_n1762, u2_uk_n1763, u2_uk_n1767, u2_uk_n1768, u2_uk_n1769, 
        u2_uk_n1770, u2_uk_n1772, u2_uk_n1773, u2_uk_n1776, u2_uk_n1777, u2_uk_n1778, u2_uk_n1779, u2_uk_n1781, u2_uk_n1782, 
        u2_uk_n1783, u2_uk_n1785, u2_uk_n1786, u2_uk_n1788, u2_uk_n1789, u2_uk_n1790, u2_uk_n1791, u2_uk_n1792, u2_uk_n1793, 
        u2_uk_n1794, u2_uk_n1796, u2_uk_n1797, u2_uk_n1799, u2_uk_n1800, u2_uk_n1801, u2_uk_n1802, u2_uk_n1803, u2_uk_n1805, 
        u2_uk_n1806, u2_uk_n1807, u2_uk_n1808, u2_uk_n1809, u2_uk_n1810, u2_uk_n1811, u2_uk_n1814, u2_uk_n1815, u2_uk_n1816, 
        u2_uk_n1817, u2_uk_n1818, u2_uk_n1819, u2_uk_n1820, u2_uk_n1821, u2_uk_n1822, u2_uk_n1823, u2_uk_n1824, u2_uk_n1825, 
        u2_uk_n1826, u2_uk_n1828, u2_uk_n1832, u2_uk_n1833, u2_uk_n1834, u2_uk_n1835, u2_uk_n1836, u2_uk_n1837, u2_uk_n1838, 
        u2_uk_n1839, u2_uk_n1840, u2_uk_n1842, u2_uk_n1843, u2_uk_n1845, u2_uk_n1846, u2_uk_n1849, u2_uk_n1850, u2_uk_n1851, 
        u2_uk_n1852, u2_uk_n1853, u2_uk_n1854, u2_uk_n1855, u2_uk_n1856, u2_uk_n238, u2_uk_n240, u2_uk_n251, u2_uk_n257, 
        u2_uk_n299, u2_uk_n313, u2_uk_n319, u2_uk_n363, u2_uk_n373, u2_uk_n376, u2_uk_n377, u2_uk_n379, u2_uk_n385, 
        u2_uk_n408, u2_uk_n415, u2_uk_n421, u2_uk_n443, u2_uk_n456, u2_uk_n467, u2_uk_n468, u2_uk_n472, u2_uk_n500, 
        u2_uk_n503, u2_uk_n504, u2_uk_n520, u2_uk_n526, u2_uk_n551, u2_uk_n586, u2_uk_n608, u2_uk_n665, u2_uk_n677, 
        u2_uk_n682, u2_uk_n689, u2_uk_n702, u2_uk_n931, u2_uk_n933, u2_uk_n939, u2_uk_n941, u2_uk_n942, u2_uk_n943, 
        u2_uk_n944, u2_uk_n945, u2_uk_n947, u2_uk_n948, u2_uk_n954, u2_uk_n955, u2_uk_n956, u2_uk_n961, u2_uk_n967, 
        u2_uk_n970, u2_uk_n972, u2_uk_n979, u2_uk_n984, u2_uk_n986, u2_uk_n994, u2_uk_n996, u2_uk_n997;
  wire key_a_0, key_a_1, key_a_10, key_a_11, key_a_12, key_a_13, key_a_14, key_a_15, key_a_16, 
       key_a_17, key_a_18, key_a_19, key_a_2, key_a_20, key_a_21, key_a_22, key_a_23, key_a_24, 
       key_a_25, key_a_26, key_a_27, key_a_28, key_a_29, key_a_3, key_a_30, key_a_31, key_a_32, 
       key_a_33, key_a_34, key_a_35, key_a_36, key_a_37, key_a_38, key_a_39, key_a_4, key_a_40, 
       key_a_41, key_a_42, key_a_43, key_a_44, key_a_45, key_a_46, key_a_47, key_a_48, key_a_49, 
       key_a_5, key_a_50, key_a_51, key_a_52, key_a_53, key_a_54, key_a_55, key_a_6, key_a_7, 
       key_a_8, key_a_9, key_b_r_0_0, key_b_r_0_1, key_b_r_0_10, key_b_r_0_11, key_b_r_0_12, key_b_r_0_13, key_b_r_0_14, 
       key_b_r_0_15, key_b_r_0_16, key_b_r_0_17, key_b_r_0_18, key_b_r_0_19, key_b_r_0_2, key_b_r_0_20, key_b_r_0_21, key_b_r_0_22, 
       key_b_r_0_23, key_b_r_0_24, key_b_r_0_25, key_b_r_0_26, key_b_r_0_27, key_b_r_0_28, key_b_r_0_29, key_b_r_0_3, key_b_r_0_30, 
       key_b_r_0_31, key_b_r_0_32, key_b_r_0_33, key_b_r_0_34, key_b_r_0_35, key_b_r_0_36, key_b_r_0_37, key_b_r_0_38, key_b_r_0_39, 
       key_b_r_0_4, key_b_r_0_40, key_b_r_0_41, key_b_r_0_42, key_b_r_0_43, key_b_r_0_44, key_b_r_0_45, key_b_r_0_46, key_b_r_0_47, 
       key_b_r_0_48, key_b_r_0_49, key_b_r_0_5, key_b_r_0_50, key_b_r_0_51, key_b_r_0_52, key_b_r_0_53, key_b_r_0_54, key_b_r_0_55, 
       key_b_r_0_6, key_b_r_0_7, key_b_r_0_8, key_b_r_0_9, key_b_r_10_0, key_b_r_10_1, key_b_r_10_10, key_b_r_10_11, key_b_r_10_12, 
       key_b_r_10_13, key_b_r_10_14, key_b_r_10_15, key_b_r_10_16, key_b_r_10_17, key_b_r_10_18, key_b_r_10_19, key_b_r_10_2, key_b_r_10_20, 
       key_b_r_10_21, key_b_r_10_22, key_b_r_10_23, key_b_r_10_24, key_b_r_10_25, key_b_r_10_26, key_b_r_10_27, key_b_r_10_28, key_b_r_10_29, 
       key_b_r_10_3, key_b_r_10_30, key_b_r_10_31, key_b_r_10_32, key_b_r_10_33, key_b_r_10_34, key_b_r_10_35, key_b_r_10_36, key_b_r_10_37, 
       key_b_r_10_38, key_b_r_10_39, key_b_r_10_4, key_b_r_10_40, key_b_r_10_41, key_b_r_10_42, key_b_r_10_43, key_b_r_10_44, key_b_r_10_45, 
       key_b_r_10_46, key_b_r_10_47, key_b_r_10_48, key_b_r_10_49, key_b_r_10_5, key_b_r_10_50, key_b_r_10_51, key_b_r_10_52, key_b_r_10_53, 
       key_b_r_10_54, key_b_r_10_55, key_b_r_10_6, key_b_r_10_7, key_b_r_10_8, key_b_r_10_9, key_b_r_11_0, key_b_r_11_1, key_b_r_11_10, 
       key_b_r_11_11, key_b_r_11_12, key_b_r_11_13, key_b_r_11_14, key_b_r_11_15, key_b_r_11_16, key_b_r_11_17, key_b_r_11_18, key_b_r_11_19, 
       key_b_r_11_2, key_b_r_11_20, key_b_r_11_21, key_b_r_11_22, key_b_r_11_23, key_b_r_11_24, key_b_r_11_25, key_b_r_11_26, key_b_r_11_27, 
       key_b_r_11_28, key_b_r_11_29, key_b_r_11_3, key_b_r_11_30, key_b_r_11_31, key_b_r_11_32, key_b_r_11_33, key_b_r_11_34, key_b_r_11_35, 
       key_b_r_11_36, key_b_r_11_37, key_b_r_11_38, key_b_r_11_39, key_b_r_11_4, key_b_r_11_40, key_b_r_11_41, key_b_r_11_42, key_b_r_11_43, 
       key_b_r_11_44, key_b_r_11_45, key_b_r_11_46, key_b_r_11_47, key_b_r_11_48, key_b_r_11_49, key_b_r_11_5, key_b_r_11_50, key_b_r_11_51, 
       key_b_r_11_52, key_b_r_11_53, key_b_r_11_54, key_b_r_11_55, key_b_r_11_6, key_b_r_11_7, key_b_r_11_8, key_b_r_11_9, key_b_r_12_0, 
       key_b_r_12_1, key_b_r_12_10, key_b_r_12_11, key_b_r_12_12, key_b_r_12_13, key_b_r_12_14, key_b_r_12_15, key_b_r_12_16, key_b_r_12_17, 
       key_b_r_12_18, key_b_r_12_19, key_b_r_12_2, key_b_r_12_20, key_b_r_12_21, key_b_r_12_22, key_b_r_12_23, key_b_r_12_24, key_b_r_12_25, 
       key_b_r_12_26, key_b_r_12_27, key_b_r_12_28, key_b_r_12_29, key_b_r_12_3, key_b_r_12_30, key_b_r_12_31, key_b_r_12_32, key_b_r_12_33, 
       key_b_r_12_34, key_b_r_12_35, key_b_r_12_36, key_b_r_12_37, key_b_r_12_38, key_b_r_12_39, key_b_r_12_4, key_b_r_12_40, key_b_r_12_41, 
       key_b_r_12_42, key_b_r_12_43, key_b_r_12_44, key_b_r_12_45, key_b_r_12_46, key_b_r_12_47, key_b_r_12_48, key_b_r_12_49, key_b_r_12_5, 
       key_b_r_12_50, key_b_r_12_51, key_b_r_12_52, key_b_r_12_53, key_b_r_12_54, key_b_r_12_55, key_b_r_12_6, key_b_r_12_7, key_b_r_12_8, 
       key_b_r_12_9, key_b_r_13_0, key_b_r_13_1, key_b_r_13_10, key_b_r_13_11, key_b_r_13_12, key_b_r_13_13, key_b_r_13_14, key_b_r_13_15, 
       key_b_r_13_16, key_b_r_13_17, key_b_r_13_18, key_b_r_13_19, key_b_r_13_2, key_b_r_13_20, key_b_r_13_21, key_b_r_13_22, key_b_r_13_23, 
       key_b_r_13_24, key_b_r_13_25, key_b_r_13_26, key_b_r_13_27, key_b_r_13_28, key_b_r_13_29, key_b_r_13_3, key_b_r_13_30, key_b_r_13_31, 
       key_b_r_13_32, key_b_r_13_33, key_b_r_13_34, key_b_r_13_35, key_b_r_13_36, key_b_r_13_37, key_b_r_13_38, key_b_r_13_39, key_b_r_13_4, 
       key_b_r_13_40, key_b_r_13_41, key_b_r_13_42, key_b_r_13_43, key_b_r_13_44, key_b_r_13_45, key_b_r_13_46, key_b_r_13_47, key_b_r_13_48, 
       key_b_r_13_49, key_b_r_13_5, key_b_r_13_50, key_b_r_13_51, key_b_r_13_52, key_b_r_13_53, key_b_r_13_54, key_b_r_13_55, key_b_r_13_6, 
       key_b_r_13_7, key_b_r_13_8, key_b_r_13_9, key_b_r_14_0, key_b_r_14_1, key_b_r_14_10, key_b_r_14_11, key_b_r_14_12, key_b_r_14_13, 
       key_b_r_14_14, key_b_r_14_15, key_b_r_14_16, key_b_r_14_17, key_b_r_14_18, key_b_r_14_19, key_b_r_14_2, key_b_r_14_20, key_b_r_14_21, 
       key_b_r_14_22, key_b_r_14_23, key_b_r_14_24, key_b_r_14_25, key_b_r_14_26, key_b_r_14_27, key_b_r_14_28, key_b_r_14_29, key_b_r_14_3, 
       key_b_r_14_30, key_b_r_14_31, key_b_r_14_32, key_b_r_14_33, key_b_r_14_34, key_b_r_14_35, key_b_r_14_36, key_b_r_14_37, key_b_r_14_38, 
       key_b_r_14_39, key_b_r_14_4, key_b_r_14_40, key_b_r_14_41, key_b_r_14_42, key_b_r_14_43, key_b_r_14_44, key_b_r_14_45, key_b_r_14_46, 
       key_b_r_14_47, key_b_r_14_48, key_b_r_14_49, key_b_r_14_5, key_b_r_14_50, key_b_r_14_51, key_b_r_14_52, key_b_r_14_53, key_b_r_14_54, 
       key_b_r_14_55, key_b_r_14_6, key_b_r_14_7, key_b_r_14_8, key_b_r_14_9, key_b_r_15_0, key_b_r_15_1, key_b_r_15_10, key_b_r_15_11, 
       key_b_r_15_12, key_b_r_15_13, key_b_r_15_14, key_b_r_15_15, key_b_r_15_16, key_b_r_15_17, key_b_r_15_18, key_b_r_15_19, key_b_r_15_2, 
       key_b_r_15_20, key_b_r_15_21, key_b_r_15_22, key_b_r_15_23, key_b_r_15_24, key_b_r_15_25, key_b_r_15_26, key_b_r_15_27, key_b_r_15_28, 
       key_b_r_15_29, key_b_r_15_3, key_b_r_15_30, key_b_r_15_31, key_b_r_15_32, key_b_r_15_33, key_b_r_15_34, key_b_r_15_35, key_b_r_15_36, 
       key_b_r_15_37, key_b_r_15_38, key_b_r_15_39, key_b_r_15_4, key_b_r_15_40, key_b_r_15_41, key_b_r_15_42, key_b_r_15_43, key_b_r_15_44, 
       key_b_r_15_45, key_b_r_15_46, key_b_r_15_47, key_b_r_15_48, key_b_r_15_49, key_b_r_15_5, key_b_r_15_50, key_b_r_15_51, key_b_r_15_52, 
       key_b_r_15_53, key_b_r_15_54, key_b_r_15_55, key_b_r_15_6, key_b_r_15_7, key_b_r_15_8, key_b_r_15_9, key_b_r_16_0, key_b_r_16_1, 
       key_b_r_16_10, key_b_r_16_11, key_b_r_16_12, key_b_r_16_13, key_b_r_16_14, key_b_r_16_15, key_b_r_16_16, key_b_r_16_17, key_b_r_16_18, 
       key_b_r_16_19, key_b_r_16_2, key_b_r_16_20, key_b_r_16_21, key_b_r_16_22, key_b_r_16_23, key_b_r_16_24, key_b_r_16_25, key_b_r_16_26, 
       key_b_r_16_27, key_b_r_16_28, key_b_r_16_29, key_b_r_16_3, key_b_r_16_30, key_b_r_16_31, key_b_r_16_32, key_b_r_16_33, key_b_r_16_34, 
       key_b_r_16_35, key_b_r_16_36, key_b_r_16_37, key_b_r_16_38, key_b_r_16_39, key_b_r_16_4, key_b_r_16_40, key_b_r_16_41, key_b_r_16_42, 
       key_b_r_16_43, key_b_r_16_44, key_b_r_16_45, key_b_r_16_46, key_b_r_16_47, key_b_r_16_48, key_b_r_16_49, key_b_r_16_5, key_b_r_16_50, 
       key_b_r_16_51, key_b_r_16_52, key_b_r_16_53, key_b_r_16_54, key_b_r_16_55, key_b_r_16_6, key_b_r_16_7, key_b_r_16_8, key_b_r_16_9, 
       key_b_r_1_0, key_b_r_1_1, key_b_r_1_10, key_b_r_1_11, key_b_r_1_12, key_b_r_1_13, key_b_r_1_14, key_b_r_1_15, key_b_r_1_16, 
       key_b_r_1_17, key_b_r_1_18, key_b_r_1_19, key_b_r_1_2, key_b_r_1_20, key_b_r_1_21, key_b_r_1_22, key_b_r_1_23, key_b_r_1_24, 
       key_b_r_1_25, key_b_r_1_26, key_b_r_1_27, key_b_r_1_28, key_b_r_1_29, key_b_r_1_3, key_b_r_1_30, key_b_r_1_31, key_b_r_1_32, 
       key_b_r_1_33, key_b_r_1_34, key_b_r_1_35, key_b_r_1_36, key_b_r_1_37, key_b_r_1_38, key_b_r_1_39, key_b_r_1_4, key_b_r_1_40, 
       key_b_r_1_41, key_b_r_1_42, key_b_r_1_43, key_b_r_1_44, key_b_r_1_45, key_b_r_1_46, key_b_r_1_47, key_b_r_1_48, key_b_r_1_49, 
       key_b_r_1_5, key_b_r_1_50, key_b_r_1_51, key_b_r_1_52, key_b_r_1_53, key_b_r_1_54, key_b_r_1_55, key_b_r_1_6, key_b_r_1_7, 
       key_b_r_1_8, key_b_r_1_9, key_b_r_2_0, key_b_r_2_1, key_b_r_2_10, key_b_r_2_11, key_b_r_2_12, key_b_r_2_13, key_b_r_2_14, 
       key_b_r_2_15, key_b_r_2_16, key_b_r_2_17, key_b_r_2_18, key_b_r_2_19, key_b_r_2_2, key_b_r_2_20, key_b_r_2_21, key_b_r_2_22, 
       key_b_r_2_23, key_b_r_2_24, key_b_r_2_25, key_b_r_2_26, key_b_r_2_27, key_b_r_2_28, key_b_r_2_29, key_b_r_2_3, key_b_r_2_30, 
       key_b_r_2_31, key_b_r_2_32, key_b_r_2_33, key_b_r_2_34, key_b_r_2_35, key_b_r_2_36, key_b_r_2_37, key_b_r_2_38, key_b_r_2_39, 
       key_b_r_2_4, key_b_r_2_40, key_b_r_2_41, key_b_r_2_42, key_b_r_2_43, key_b_r_2_44, key_b_r_2_45, key_b_r_2_46, key_b_r_2_47, 
       key_b_r_2_48, key_b_r_2_49, key_b_r_2_5, key_b_r_2_50, key_b_r_2_51, key_b_r_2_52, key_b_r_2_53, key_b_r_2_54, key_b_r_2_55, 
       key_b_r_2_6, key_b_r_2_7, key_b_r_2_8, key_b_r_2_9, key_b_r_3_0, key_b_r_3_1, key_b_r_3_10, key_b_r_3_11, key_b_r_3_12, 
       key_b_r_3_13, key_b_r_3_14, key_b_r_3_15, key_b_r_3_16, key_b_r_3_17, key_b_r_3_18, key_b_r_3_19, key_b_r_3_2, key_b_r_3_20, 
       key_b_r_3_21, key_b_r_3_22, key_b_r_3_23, key_b_r_3_24, key_b_r_3_25, key_b_r_3_26, key_b_r_3_27, key_b_r_3_28, key_b_r_3_29, 
       key_b_r_3_3, key_b_r_3_30, key_b_r_3_31, key_b_r_3_32, key_b_r_3_33, key_b_r_3_34, key_b_r_3_35, key_b_r_3_36, key_b_r_3_37, 
       key_b_r_3_38, key_b_r_3_39, key_b_r_3_4, key_b_r_3_40, key_b_r_3_41, key_b_r_3_42, key_b_r_3_43, key_b_r_3_44, key_b_r_3_45, 
       key_b_r_3_46, key_b_r_3_47, key_b_r_3_48, key_b_r_3_49, key_b_r_3_5, key_b_r_3_50, key_b_r_3_51, key_b_r_3_52, key_b_r_3_53, 
       key_b_r_3_54, key_b_r_3_55, key_b_r_3_6, key_b_r_3_7, key_b_r_3_8, key_b_r_3_9, key_b_r_4_0, key_b_r_4_1, key_b_r_4_10, 
       key_b_r_4_11, key_b_r_4_12, key_b_r_4_13, key_b_r_4_14, key_b_r_4_15, key_b_r_4_16, key_b_r_4_17, key_b_r_4_18, key_b_r_4_19, 
       key_b_r_4_2, key_b_r_4_20, key_b_r_4_21, key_b_r_4_22, key_b_r_4_23, key_b_r_4_24, key_b_r_4_25, key_b_r_4_26, key_b_r_4_27, 
       key_b_r_4_28, key_b_r_4_29, key_b_r_4_3, key_b_r_4_30, key_b_r_4_31, key_b_r_4_32, key_b_r_4_33, key_b_r_4_34, key_b_r_4_35, 
       key_b_r_4_36, key_b_r_4_37, key_b_r_4_38, key_b_r_4_39, key_b_r_4_4, key_b_r_4_40, key_b_r_4_41, key_b_r_4_42, key_b_r_4_43, 
       key_b_r_4_44, key_b_r_4_45, key_b_r_4_46, key_b_r_4_47, key_b_r_4_48, key_b_r_4_49, key_b_r_4_5, key_b_r_4_50, key_b_r_4_51, 
       key_b_r_4_52, key_b_r_4_53, key_b_r_4_54, key_b_r_4_55, key_b_r_4_6, key_b_r_4_7, key_b_r_4_8, key_b_r_4_9, key_b_r_5_0, 
       key_b_r_5_1, key_b_r_5_10, key_b_r_5_11, key_b_r_5_12, key_b_r_5_13, key_b_r_5_14, key_b_r_5_15, key_b_r_5_16, key_b_r_5_17, 
       key_b_r_5_18, key_b_r_5_19, key_b_r_5_2, key_b_r_5_20, key_b_r_5_21, key_b_r_5_22, key_b_r_5_23, key_b_r_5_24, key_b_r_5_25, 
       key_b_r_5_26, key_b_r_5_27, key_b_r_5_28, key_b_r_5_29, key_b_r_5_3, key_b_r_5_30, key_b_r_5_31, key_b_r_5_32, key_b_r_5_33, 
       key_b_r_5_34, key_b_r_5_35, key_b_r_5_36, key_b_r_5_37, key_b_r_5_38, key_b_r_5_39, key_b_r_5_4, key_b_r_5_40, key_b_r_5_41, 
       key_b_r_5_42, key_b_r_5_43, key_b_r_5_44, key_b_r_5_45, key_b_r_5_46, key_b_r_5_47, key_b_r_5_48, key_b_r_5_49, key_b_r_5_5, 
       key_b_r_5_50, key_b_r_5_51, key_b_r_5_52, key_b_r_5_53, key_b_r_5_54, key_b_r_5_55, key_b_r_5_6, key_b_r_5_7, key_b_r_5_8, 
       key_b_r_5_9, key_b_r_6_0, key_b_r_6_1, key_b_r_6_10, key_b_r_6_11, key_b_r_6_12, key_b_r_6_13, key_b_r_6_14, key_b_r_6_15, 
       key_b_r_6_16, key_b_r_6_17, key_b_r_6_18, key_b_r_6_19, key_b_r_6_2, key_b_r_6_20, key_b_r_6_21, key_b_r_6_22, key_b_r_6_23, 
       key_b_r_6_24, key_b_r_6_25, key_b_r_6_26, key_b_r_6_27, key_b_r_6_28, key_b_r_6_29, key_b_r_6_3, key_b_r_6_30, key_b_r_6_31, 
       key_b_r_6_32, key_b_r_6_33, key_b_r_6_34, key_b_r_6_35, key_b_r_6_36, key_b_r_6_37, key_b_r_6_38, key_b_r_6_39, key_b_r_6_4, 
       key_b_r_6_40, key_b_r_6_41, key_b_r_6_42, key_b_r_6_43, key_b_r_6_44, key_b_r_6_45, key_b_r_6_46, key_b_r_6_47, key_b_r_6_48, 
       key_b_r_6_49, key_b_r_6_5, key_b_r_6_50, key_b_r_6_51, key_b_r_6_52, key_b_r_6_53, key_b_r_6_54, key_b_r_6_55, key_b_r_6_6, 
       key_b_r_6_7, key_b_r_6_8, key_b_r_6_9, key_b_r_7_0, key_b_r_7_1, key_b_r_7_10, key_b_r_7_11, key_b_r_7_12, key_b_r_7_13, 
       key_b_r_7_14, key_b_r_7_15, key_b_r_7_16, key_b_r_7_17, key_b_r_7_18, key_b_r_7_19, key_b_r_7_2, key_b_r_7_20, key_b_r_7_21, 
       key_b_r_7_22, key_b_r_7_23, key_b_r_7_24, key_b_r_7_25, key_b_r_7_26, key_b_r_7_27, key_b_r_7_28, key_b_r_7_29, key_b_r_7_3, 
       key_b_r_7_30, key_b_r_7_31, key_b_r_7_32, key_b_r_7_33, key_b_r_7_34, key_b_r_7_35, key_b_r_7_36, key_b_r_7_37, key_b_r_7_38, 
       key_b_r_7_39, key_b_r_7_4, key_b_r_7_40, key_b_r_7_41, key_b_r_7_42, key_b_r_7_43, key_b_r_7_44, key_b_r_7_45, key_b_r_7_46, 
       key_b_r_7_47, key_b_r_7_48, key_b_r_7_49, key_b_r_7_5, key_b_r_7_50, key_b_r_7_51, key_b_r_7_52, key_b_r_7_53, key_b_r_7_54, 
       key_b_r_7_55, key_b_r_7_6, key_b_r_7_7, key_b_r_7_8, key_b_r_7_9, key_b_r_8_0, key_b_r_8_1, key_b_r_8_10, key_b_r_8_11, 
       key_b_r_8_12, key_b_r_8_13, key_b_r_8_14, key_b_r_8_15, key_b_r_8_16, key_b_r_8_17, key_b_r_8_18, key_b_r_8_19, key_b_r_8_2, 
       key_b_r_8_20, key_b_r_8_21, key_b_r_8_22, key_b_r_8_23, key_b_r_8_24, key_b_r_8_25, key_b_r_8_26, key_b_r_8_27, key_b_r_8_28, 
       key_b_r_8_29, key_b_r_8_3, key_b_r_8_30, key_b_r_8_31, key_b_r_8_32, key_b_r_8_33, key_b_r_8_34, key_b_r_8_35, key_b_r_8_36, 
       key_b_r_8_37, key_b_r_8_38, key_b_r_8_39, key_b_r_8_4, key_b_r_8_40, key_b_r_8_41, key_b_r_8_42, key_b_r_8_43, key_b_r_8_44, 
       key_b_r_8_45, key_b_r_8_46, key_b_r_8_47, key_b_r_8_48, key_b_r_8_49, key_b_r_8_5, key_b_r_8_50, key_b_r_8_51, key_b_r_8_52, 
       key_b_r_8_53, key_b_r_8_54, key_b_r_8_55, key_b_r_8_6, key_b_r_8_7, key_b_r_8_8, key_b_r_8_9, key_b_r_9_0, key_b_r_9_1, 
       key_b_r_9_10, key_b_r_9_11, key_b_r_9_12, key_b_r_9_13, key_b_r_9_14, key_b_r_9_15, key_b_r_9_16, key_b_r_9_17, key_b_r_9_18, 
       key_b_r_9_19, key_b_r_9_2, key_b_r_9_20, key_b_r_9_21, key_b_r_9_22, key_b_r_9_23, key_b_r_9_24, key_b_r_9_25, key_b_r_9_26, 
       key_b_r_9_27, key_b_r_9_28, key_b_r_9_29, key_b_r_9_3, key_b_r_9_30, key_b_r_9_31, key_b_r_9_32, key_b_r_9_33, key_b_r_9_34, 
       key_b_r_9_35, key_b_r_9_36, key_b_r_9_37, key_b_r_9_38, key_b_r_9_39, key_b_r_9_4, key_b_r_9_40, key_b_r_9_41, key_b_r_9_42, 
       key_b_r_9_43, key_b_r_9_44, key_b_r_9_45, key_b_r_9_46, key_b_r_9_47, key_b_r_9_48, key_b_r_9_49, key_b_r_9_5, key_b_r_9_50, 
       key_b_r_9_51, key_b_r_9_52, key_b_r_9_53, key_b_r_9_54, key_b_r_9_55, key_b_r_9_6, key_b_r_9_7, key_b_r_9_8, key_b_r_9_9, 
       key_c_r_0_0, key_c_r_0_1, key_c_r_0_10, key_c_r_0_11, key_c_r_0_12, key_c_r_0_13, key_c_r_0_14, key_c_r_0_15, key_c_r_0_16, 
       key_c_r_0_17, key_c_r_0_18, key_c_r_0_19, key_c_r_0_2, key_c_r_0_20, key_c_r_0_21, key_c_r_0_22, key_c_r_0_23, key_c_r_0_24, 
       key_c_r_0_25, key_c_r_0_26, key_c_r_0_27, key_c_r_0_28, key_c_r_0_29, key_c_r_0_3, key_c_r_0_30, key_c_r_0_31, key_c_r_0_32, 
       key_c_r_0_33, key_c_r_0_34, key_c_r_0_35, key_c_r_0_36, key_c_r_0_37, key_c_r_0_38, key_c_r_0_39, key_c_r_0_4, key_c_r_0_40, 
       key_c_r_0_41, key_c_r_0_42, key_c_r_0_43, key_c_r_0_44, key_c_r_0_45, key_c_r_0_46, key_c_r_0_47, key_c_r_0_48, key_c_r_0_49, 
       key_c_r_0_5, key_c_r_0_50, key_c_r_0_51, key_c_r_0_52, key_c_r_0_53, key_c_r_0_54, key_c_r_0_55, key_c_r_0_6, key_c_r_0_7, 
       key_c_r_0_8, key_c_r_0_9, key_c_r_10_0, key_c_r_10_1, key_c_r_10_10, key_c_r_10_11, key_c_r_10_12, key_c_r_10_13, key_c_r_10_14, 
       key_c_r_10_15, key_c_r_10_16, key_c_r_10_17, key_c_r_10_18, key_c_r_10_19, key_c_r_10_2, key_c_r_10_20, key_c_r_10_21, key_c_r_10_22, 
       key_c_r_10_23, key_c_r_10_24, key_c_r_10_25, key_c_r_10_26, key_c_r_10_27, key_c_r_10_28, key_c_r_10_29, key_c_r_10_3, key_c_r_10_30, 
       key_c_r_10_31, key_c_r_10_32, key_c_r_10_33, key_c_r_10_34, key_c_r_10_35, key_c_r_10_36, key_c_r_10_37, key_c_r_10_38, key_c_r_10_39, 
       key_c_r_10_4, key_c_r_10_40, key_c_r_10_41, key_c_r_10_42, key_c_r_10_43, key_c_r_10_44, key_c_r_10_45, key_c_r_10_46, key_c_r_10_47, 
       key_c_r_10_48, key_c_r_10_49, key_c_r_10_5, key_c_r_10_50, key_c_r_10_51, key_c_r_10_52, key_c_r_10_53, key_c_r_10_54, key_c_r_10_55, 
       key_c_r_10_6, key_c_r_10_7, key_c_r_10_8, key_c_r_10_9, key_c_r_11_0, key_c_r_11_1, key_c_r_11_10, key_c_r_11_11, key_c_r_11_12, 
       key_c_r_11_13, key_c_r_11_14, key_c_r_11_15, key_c_r_11_16, key_c_r_11_17, key_c_r_11_18, key_c_r_11_19, key_c_r_11_2, key_c_r_11_20, 
       key_c_r_11_21, key_c_r_11_22, key_c_r_11_23, key_c_r_11_24, key_c_r_11_25, key_c_r_11_26, key_c_r_11_27, key_c_r_11_28, key_c_r_11_29, 
       key_c_r_11_3, key_c_r_11_30, key_c_r_11_31, key_c_r_11_32, key_c_r_11_33, key_c_r_11_34, key_c_r_11_35, key_c_r_11_36, key_c_r_11_37, 
       key_c_r_11_38, key_c_r_11_39, key_c_r_11_4, key_c_r_11_40, key_c_r_11_41, key_c_r_11_42, key_c_r_11_43, key_c_r_11_44, key_c_r_11_45, 
       key_c_r_11_46, key_c_r_11_47, key_c_r_11_48, key_c_r_11_49, key_c_r_11_5, key_c_r_11_50, key_c_r_11_51, key_c_r_11_52, key_c_r_11_53, 
       key_c_r_11_54, key_c_r_11_55, key_c_r_11_6, key_c_r_11_7, key_c_r_11_8, key_c_r_11_9, key_c_r_12_0, key_c_r_12_1, key_c_r_12_10, 
       key_c_r_12_11, key_c_r_12_12, key_c_r_12_13, key_c_r_12_14, key_c_r_12_15, key_c_r_12_16, key_c_r_12_17, key_c_r_12_18, key_c_r_12_19, 
       key_c_r_12_2, key_c_r_12_20, key_c_r_12_21, key_c_r_12_22, key_c_r_12_23, key_c_r_12_24, key_c_r_12_25, key_c_r_12_26, key_c_r_12_27, 
       key_c_r_12_28, key_c_r_12_29, key_c_r_12_3, key_c_r_12_30, key_c_r_12_31, key_c_r_12_32, key_c_r_12_33, key_c_r_12_34, key_c_r_12_35, 
       key_c_r_12_36, key_c_r_12_37, key_c_r_12_38, key_c_r_12_39, key_c_r_12_4, key_c_r_12_40, key_c_r_12_41, key_c_r_12_42, key_c_r_12_43, 
       key_c_r_12_44, key_c_r_12_45, key_c_r_12_46, key_c_r_12_47, key_c_r_12_48, key_c_r_12_49, key_c_r_12_5, key_c_r_12_50, key_c_r_12_51, 
       key_c_r_12_52, key_c_r_12_53, key_c_r_12_54, key_c_r_12_55, key_c_r_12_6, key_c_r_12_7, key_c_r_12_8, key_c_r_12_9, key_c_r_13_0, 
       key_c_r_13_1, key_c_r_13_10, key_c_r_13_11, key_c_r_13_12, key_c_r_13_13, key_c_r_13_14, key_c_r_13_15, key_c_r_13_16, key_c_r_13_17, 
       key_c_r_13_18, key_c_r_13_19, key_c_r_13_2, key_c_r_13_20, key_c_r_13_21, key_c_r_13_22, key_c_r_13_23, key_c_r_13_24, key_c_r_13_25, 
       key_c_r_13_26, key_c_r_13_27, key_c_r_13_28, key_c_r_13_29, key_c_r_13_3, key_c_r_13_30, key_c_r_13_31, key_c_r_13_32, key_c_r_13_33, 
       key_c_r_13_34, key_c_r_13_35, key_c_r_13_36, key_c_r_13_37, key_c_r_13_38, key_c_r_13_39, key_c_r_13_4, key_c_r_13_40, key_c_r_13_41, 
       key_c_r_13_42, key_c_r_13_43, key_c_r_13_44, key_c_r_13_45, key_c_r_13_46, key_c_r_13_47, key_c_r_13_48, key_c_r_13_49, key_c_r_13_5, 
       key_c_r_13_50, key_c_r_13_51, key_c_r_13_52, key_c_r_13_53, key_c_r_13_54, key_c_r_13_55, key_c_r_13_6, key_c_r_13_7, key_c_r_13_8, 
       key_c_r_13_9, key_c_r_14_0, key_c_r_14_1, key_c_r_14_10, key_c_r_14_11, key_c_r_14_12, key_c_r_14_13, key_c_r_14_14, key_c_r_14_15, 
       key_c_r_14_16, key_c_r_14_17, key_c_r_14_18, key_c_r_14_19, key_c_r_14_2, key_c_r_14_20, key_c_r_14_21, key_c_r_14_22, key_c_r_14_23, 
       key_c_r_14_24, key_c_r_14_25, key_c_r_14_26, key_c_r_14_27, key_c_r_14_28, key_c_r_14_29, key_c_r_14_3, key_c_r_14_30, key_c_r_14_31, 
       key_c_r_14_32, key_c_r_14_33, key_c_r_14_34, key_c_r_14_35, key_c_r_14_36, key_c_r_14_37, key_c_r_14_38, key_c_r_14_39, key_c_r_14_4, 
       key_c_r_14_40, key_c_r_14_41, key_c_r_14_42, key_c_r_14_43, key_c_r_14_44, key_c_r_14_45, key_c_r_14_46, key_c_r_14_47, key_c_r_14_48, 
       key_c_r_14_49, key_c_r_14_5, key_c_r_14_50, key_c_r_14_51, key_c_r_14_52, key_c_r_14_53, key_c_r_14_54, key_c_r_14_55, key_c_r_14_6, 
       key_c_r_14_7, key_c_r_14_8, key_c_r_14_9, key_c_r_15_0, key_c_r_15_1, key_c_r_15_10, key_c_r_15_11, key_c_r_15_12, key_c_r_15_13, 
       key_c_r_15_14, key_c_r_15_15, key_c_r_15_16, key_c_r_15_17, key_c_r_15_18, key_c_r_15_19, key_c_r_15_2, key_c_r_15_20, key_c_r_15_21, 
       key_c_r_15_22, key_c_r_15_23, key_c_r_15_24, key_c_r_15_25, key_c_r_15_26, key_c_r_15_27, key_c_r_15_28, key_c_r_15_29, key_c_r_15_3, 
       key_c_r_15_30, key_c_r_15_31, key_c_r_15_32, key_c_r_15_33, key_c_r_15_34, key_c_r_15_35, key_c_r_15_36, key_c_r_15_37, key_c_r_15_38, 
       key_c_r_15_39, key_c_r_15_4, key_c_r_15_40, key_c_r_15_41, key_c_r_15_42, key_c_r_15_43, key_c_r_15_44, key_c_r_15_45, key_c_r_15_46, 
       key_c_r_15_47, key_c_r_15_48, key_c_r_15_49, key_c_r_15_5, key_c_r_15_50, key_c_r_15_51, key_c_r_15_52, key_c_r_15_53, key_c_r_15_54, 
       key_c_r_15_55, key_c_r_15_6, key_c_r_15_7, key_c_r_15_8, key_c_r_15_9, key_c_r_16_0, key_c_r_16_1, key_c_r_16_10, key_c_r_16_11, 
       key_c_r_16_12, key_c_r_16_13, key_c_r_16_14, key_c_r_16_15, key_c_r_16_16, key_c_r_16_17, key_c_r_16_18, key_c_r_16_19, key_c_r_16_2, 
       key_c_r_16_20, key_c_r_16_21, key_c_r_16_22, key_c_r_16_23, key_c_r_16_24, key_c_r_16_25, key_c_r_16_26, key_c_r_16_27, key_c_r_16_28, 
       key_c_r_16_29, key_c_r_16_3, key_c_r_16_30, key_c_r_16_31, key_c_r_16_32, key_c_r_16_33, key_c_r_16_34, key_c_r_16_35, key_c_r_16_36, 
       key_c_r_16_37, key_c_r_16_38, key_c_r_16_39, key_c_r_16_4, key_c_r_16_40, key_c_r_16_41, key_c_r_16_42, key_c_r_16_43, key_c_r_16_44, 
       key_c_r_16_45, key_c_r_16_46, key_c_r_16_47, key_c_r_16_48, key_c_r_16_49, key_c_r_16_5, key_c_r_16_50, key_c_r_16_51, key_c_r_16_52, 
       key_c_r_16_53, key_c_r_16_54, key_c_r_16_55, key_c_r_16_6, key_c_r_16_7, key_c_r_16_8, key_c_r_16_9, key_c_r_17_0, key_c_r_17_1, 
       key_c_r_17_10, key_c_r_17_11, key_c_r_17_12, key_c_r_17_13, key_c_r_17_14, key_c_r_17_15, key_c_r_17_16, key_c_r_17_17, key_c_r_17_18, 
       key_c_r_17_19, key_c_r_17_2, key_c_r_17_20, key_c_r_17_21, key_c_r_17_22, key_c_r_17_23, key_c_r_17_24, key_c_r_17_25, key_c_r_17_26, 
       key_c_r_17_27, key_c_r_17_28, key_c_r_17_29, key_c_r_17_3, key_c_r_17_30, key_c_r_17_31, key_c_r_17_32, key_c_r_17_33, key_c_r_17_34, 
       key_c_r_17_35, key_c_r_17_36, key_c_r_17_37, key_c_r_17_38, key_c_r_17_39, key_c_r_17_4, key_c_r_17_40, key_c_r_17_41, key_c_r_17_42, 
       key_c_r_17_43, key_c_r_17_44, key_c_r_17_45, key_c_r_17_46, key_c_r_17_47, key_c_r_17_48, key_c_r_17_49, key_c_r_17_5, key_c_r_17_50, 
       key_c_r_17_51, key_c_r_17_52, key_c_r_17_53, key_c_r_17_54, key_c_r_17_55, key_c_r_17_6, key_c_r_17_7, key_c_r_17_8, key_c_r_17_9, 
       key_c_r_18_0, key_c_r_18_1, key_c_r_18_10, key_c_r_18_11, key_c_r_18_12, key_c_r_18_13, key_c_r_18_14, key_c_r_18_15, key_c_r_18_16, 
       key_c_r_18_17, key_c_r_18_18, key_c_r_18_19, key_c_r_18_2, key_c_r_18_20, key_c_r_18_21, key_c_r_18_22, key_c_r_18_23, key_c_r_18_24, 
       key_c_r_18_25, key_c_r_18_26, key_c_r_18_27, key_c_r_18_28, key_c_r_18_29, key_c_r_18_3, key_c_r_18_30, key_c_r_18_31, key_c_r_18_32, 
       key_c_r_18_33, key_c_r_18_34, key_c_r_18_35, key_c_r_18_36, key_c_r_18_37, key_c_r_18_38, key_c_r_18_39, key_c_r_18_4, key_c_r_18_40, 
       key_c_r_18_41, key_c_r_18_42, key_c_r_18_43, key_c_r_18_44, key_c_r_18_45, key_c_r_18_46, key_c_r_18_47, key_c_r_18_48, key_c_r_18_49, 
       key_c_r_18_5, key_c_r_18_50, key_c_r_18_51, key_c_r_18_52, key_c_r_18_53, key_c_r_18_54, key_c_r_18_55, key_c_r_18_6, key_c_r_18_7, 
       key_c_r_18_8, key_c_r_18_9, key_c_r_19_0, key_c_r_19_1, key_c_r_19_10, key_c_r_19_11, key_c_r_19_12, key_c_r_19_13, key_c_r_19_14, 
       key_c_r_19_15, key_c_r_19_16, key_c_r_19_17, key_c_r_19_18, key_c_r_19_19, key_c_r_19_2, key_c_r_19_20, key_c_r_19_21, key_c_r_19_22, 
       key_c_r_19_23, key_c_r_19_24, key_c_r_19_25, key_c_r_19_26, key_c_r_19_27, key_c_r_19_28, key_c_r_19_29, key_c_r_19_3, key_c_r_19_30, 
       key_c_r_19_31, key_c_r_19_32, key_c_r_19_33, key_c_r_19_34, key_c_r_19_35, key_c_r_19_36, key_c_r_19_37, key_c_r_19_38, key_c_r_19_39, 
       key_c_r_19_4, key_c_r_19_40, key_c_r_19_41, key_c_r_19_42, key_c_r_19_43, key_c_r_19_44, key_c_r_19_45, key_c_r_19_46, key_c_r_19_47, 
       key_c_r_19_48, key_c_r_19_49, key_c_r_19_5, key_c_r_19_50, key_c_r_19_51, key_c_r_19_52, key_c_r_19_53, key_c_r_19_54, key_c_r_19_55, 
       key_c_r_19_6, key_c_r_19_7, key_c_r_19_8, key_c_r_19_9, key_c_r_1_0, key_c_r_1_1, key_c_r_1_10, key_c_r_1_11, key_c_r_1_12, 
       key_c_r_1_13, key_c_r_1_14, key_c_r_1_15, key_c_r_1_16, key_c_r_1_17, key_c_r_1_18, key_c_r_1_19, key_c_r_1_2, key_c_r_1_20, 
       key_c_r_1_21, key_c_r_1_22, key_c_r_1_23, key_c_r_1_24, key_c_r_1_25, key_c_r_1_26, key_c_r_1_27, key_c_r_1_28, key_c_r_1_29, 
       key_c_r_1_3, key_c_r_1_30, key_c_r_1_31, key_c_r_1_32, key_c_r_1_33, key_c_r_1_34, key_c_r_1_35, key_c_r_1_36, key_c_r_1_37, 
       key_c_r_1_38, key_c_r_1_39, key_c_r_1_4, key_c_r_1_40, key_c_r_1_41, key_c_r_1_42, key_c_r_1_43, key_c_r_1_44, key_c_r_1_45, 
       key_c_r_1_46, key_c_r_1_47, key_c_r_1_48, key_c_r_1_49, key_c_r_1_5, key_c_r_1_50, key_c_r_1_51, key_c_r_1_52, key_c_r_1_53, 
       key_c_r_1_54, key_c_r_1_55, key_c_r_1_6, key_c_r_1_7, key_c_r_1_8, key_c_r_1_9, key_c_r_20_0, key_c_r_20_1, key_c_r_20_10, 
       key_c_r_20_11, key_c_r_20_12, key_c_r_20_13, key_c_r_20_14, key_c_r_20_15, key_c_r_20_16, key_c_r_20_17, key_c_r_20_18, key_c_r_20_19, 
       key_c_r_20_2, key_c_r_20_20, key_c_r_20_21, key_c_r_20_22, key_c_r_20_23, key_c_r_20_24, key_c_r_20_25, key_c_r_20_26, key_c_r_20_27, 
       key_c_r_20_28, key_c_r_20_29, key_c_r_20_3, key_c_r_20_30, key_c_r_20_31, key_c_r_20_32, key_c_r_20_33, key_c_r_20_34, key_c_r_20_35, 
       key_c_r_20_36, key_c_r_20_37, key_c_r_20_38, key_c_r_20_39, key_c_r_20_4, key_c_r_20_40, key_c_r_20_41, key_c_r_20_42, key_c_r_20_43, 
       key_c_r_20_44, key_c_r_20_45, key_c_r_20_46, key_c_r_20_47, key_c_r_20_48, key_c_r_20_49, key_c_r_20_5, key_c_r_20_50, key_c_r_20_51, 
       key_c_r_20_52, key_c_r_20_53, key_c_r_20_54, key_c_r_20_55, key_c_r_20_6, key_c_r_20_7, key_c_r_20_8, key_c_r_20_9, key_c_r_21_0, 
       key_c_r_21_1, key_c_r_21_10, key_c_r_21_11, key_c_r_21_12, key_c_r_21_13, key_c_r_21_14, key_c_r_21_15, key_c_r_21_16, key_c_r_21_17, 
       key_c_r_21_18, key_c_r_21_19, key_c_r_21_2, key_c_r_21_20, key_c_r_21_21, key_c_r_21_22, key_c_r_21_23, key_c_r_21_24, key_c_r_21_25, 
       key_c_r_21_26, key_c_r_21_27, key_c_r_21_28, key_c_r_21_29, key_c_r_21_3, key_c_r_21_30, key_c_r_21_31, key_c_r_21_32, key_c_r_21_33, 
       key_c_r_21_34, key_c_r_21_35, key_c_r_21_36, key_c_r_21_37, key_c_r_21_38, key_c_r_21_39, key_c_r_21_4, key_c_r_21_40, key_c_r_21_41, 
       key_c_r_21_42, key_c_r_21_43, key_c_r_21_44, key_c_r_21_45, key_c_r_21_46, key_c_r_21_47, key_c_r_21_48, key_c_r_21_49, key_c_r_21_5, 
       key_c_r_21_50, key_c_r_21_51, key_c_r_21_52, key_c_r_21_53, key_c_r_21_54, key_c_r_21_55, key_c_r_21_6, key_c_r_21_7, key_c_r_21_8, 
       key_c_r_21_9, key_c_r_22_0, key_c_r_22_1, key_c_r_22_10, key_c_r_22_11, key_c_r_22_12, key_c_r_22_13, key_c_r_22_14, key_c_r_22_15, 
       key_c_r_22_16, key_c_r_22_17, key_c_r_22_18, key_c_r_22_19, key_c_r_22_2, key_c_r_22_20, key_c_r_22_21, key_c_r_22_22, key_c_r_22_23, 
       key_c_r_22_24, key_c_r_22_25, key_c_r_22_26, key_c_r_22_27, key_c_r_22_28, key_c_r_22_29, key_c_r_22_3, key_c_r_22_30, key_c_r_22_31, 
       key_c_r_22_32, key_c_r_22_33, key_c_r_22_34, key_c_r_22_35, key_c_r_22_36, key_c_r_22_37, key_c_r_22_38, key_c_r_22_39, key_c_r_22_4, 
       key_c_r_22_40, key_c_r_22_41, key_c_r_22_42, key_c_r_22_43, key_c_r_22_44, key_c_r_22_45, key_c_r_22_46, key_c_r_22_47, key_c_r_22_48, 
       key_c_r_22_49, key_c_r_22_5, key_c_r_22_50, key_c_r_22_51, key_c_r_22_52, key_c_r_22_53, key_c_r_22_54, key_c_r_22_55, key_c_r_22_6, 
       key_c_r_22_7, key_c_r_22_8, key_c_r_22_9, key_c_r_23_0, key_c_r_23_1, key_c_r_23_10, key_c_r_23_11, key_c_r_23_12, key_c_r_23_13, 
       key_c_r_23_14, key_c_r_23_15, key_c_r_23_16, key_c_r_23_17, key_c_r_23_18, key_c_r_23_19, key_c_r_23_2, key_c_r_23_20, key_c_r_23_21, 
       key_c_r_23_22, key_c_r_23_23, key_c_r_23_24, key_c_r_23_25, key_c_r_23_26, key_c_r_23_27, key_c_r_23_28, key_c_r_23_29, key_c_r_23_3, 
       key_c_r_23_30, key_c_r_23_31, key_c_r_23_32, key_c_r_23_33, key_c_r_23_34, key_c_r_23_35, key_c_r_23_36, key_c_r_23_37, key_c_r_23_38, 
       key_c_r_23_39, key_c_r_23_4, key_c_r_23_40, key_c_r_23_41, key_c_r_23_42, key_c_r_23_43, key_c_r_23_44, key_c_r_23_45, key_c_r_23_46, 
       key_c_r_23_47, key_c_r_23_48, key_c_r_23_49, key_c_r_23_5, key_c_r_23_50, key_c_r_23_51, key_c_r_23_52, key_c_r_23_53, key_c_r_23_54, 
       key_c_r_23_55, key_c_r_23_6, key_c_r_23_7, key_c_r_23_8, key_c_r_23_9, key_c_r_24_0, key_c_r_24_1, key_c_r_24_10, key_c_r_24_11, 
       key_c_r_24_12, key_c_r_24_13, key_c_r_24_14, key_c_r_24_15, key_c_r_24_16, key_c_r_24_17, key_c_r_24_18, key_c_r_24_19, key_c_r_24_2, 
       key_c_r_24_20, key_c_r_24_21, key_c_r_24_22, key_c_r_24_23, key_c_r_24_24, key_c_r_24_25, key_c_r_24_26, key_c_r_24_27, key_c_r_24_28, 
       key_c_r_24_29, key_c_r_24_3, key_c_r_24_30, key_c_r_24_31, key_c_r_24_32, key_c_r_24_33, key_c_r_24_34, key_c_r_24_35, key_c_r_24_36, 
       key_c_r_24_37, key_c_r_24_38, key_c_r_24_39, key_c_r_24_4, key_c_r_24_40, key_c_r_24_41, key_c_r_24_42, key_c_r_24_43, key_c_r_24_44, 
       key_c_r_24_45, key_c_r_24_46, key_c_r_24_47, key_c_r_24_48, key_c_r_24_49, key_c_r_24_5, key_c_r_24_50, key_c_r_24_51, key_c_r_24_52, 
       key_c_r_24_53, key_c_r_24_54, key_c_r_24_55, key_c_r_24_6, key_c_r_24_7, key_c_r_24_8, key_c_r_24_9, key_c_r_25_0, key_c_r_25_1, 
       key_c_r_25_10, key_c_r_25_11, key_c_r_25_12, key_c_r_25_13, key_c_r_25_14, key_c_r_25_15, key_c_r_25_16, key_c_r_25_17, key_c_r_25_18, 
       key_c_r_25_19, key_c_r_25_2, key_c_r_25_20, key_c_r_25_21, key_c_r_25_22, key_c_r_25_23, key_c_r_25_24, key_c_r_25_25, key_c_r_25_26, 
       key_c_r_25_27, key_c_r_25_28, key_c_r_25_29, key_c_r_25_3, key_c_r_25_30, key_c_r_25_31, key_c_r_25_32, key_c_r_25_33, key_c_r_25_34, 
       key_c_r_25_35, key_c_r_25_36, key_c_r_25_37, key_c_r_25_38, key_c_r_25_39, key_c_r_25_4, key_c_r_25_40, key_c_r_25_41, key_c_r_25_42, 
       key_c_r_25_43, key_c_r_25_44, key_c_r_25_45, key_c_r_25_46, key_c_r_25_47, key_c_r_25_48, key_c_r_25_49, key_c_r_25_5, key_c_r_25_50, 
       key_c_r_25_51, key_c_r_25_52, key_c_r_25_53, key_c_r_25_54, key_c_r_25_55, key_c_r_25_6, key_c_r_25_7, key_c_r_25_8, key_c_r_25_9, 
       key_c_r_26_0, key_c_r_26_1, key_c_r_26_10, key_c_r_26_11, key_c_r_26_12, key_c_r_26_13, key_c_r_26_14, key_c_r_26_15, key_c_r_26_16, 
       key_c_r_26_17, key_c_r_26_18, key_c_r_26_19, key_c_r_26_2, key_c_r_26_20, key_c_r_26_21, key_c_r_26_22, key_c_r_26_23, key_c_r_26_24, 
       key_c_r_26_25, key_c_r_26_26, key_c_r_26_27, key_c_r_26_28, key_c_r_26_29, key_c_r_26_3, key_c_r_26_30, key_c_r_26_31, key_c_r_26_32, 
       key_c_r_26_33, key_c_r_26_34, key_c_r_26_35, key_c_r_26_36, key_c_r_26_37, key_c_r_26_38, key_c_r_26_39, key_c_r_26_4, key_c_r_26_40, 
       key_c_r_26_41, key_c_r_26_42, key_c_r_26_43, key_c_r_26_44, key_c_r_26_45, key_c_r_26_46, key_c_r_26_47, key_c_r_26_48, key_c_r_26_49, 
       key_c_r_26_5, key_c_r_26_50, key_c_r_26_51, key_c_r_26_52, key_c_r_26_53, key_c_r_26_54, key_c_r_26_55, key_c_r_26_6, key_c_r_26_7, 
       key_c_r_26_8, key_c_r_26_9, key_c_r_27_0, key_c_r_27_1, key_c_r_27_10, key_c_r_27_11, key_c_r_27_12, key_c_r_27_13, key_c_r_27_14, 
       key_c_r_27_15, key_c_r_27_16, key_c_r_27_17, key_c_r_27_18, key_c_r_27_19, key_c_r_27_2, key_c_r_27_20, key_c_r_27_21, key_c_r_27_22, 
       key_c_r_27_23, key_c_r_27_24, key_c_r_27_25, key_c_r_27_26, key_c_r_27_27, key_c_r_27_28, key_c_r_27_29, key_c_r_27_3, key_c_r_27_30, 
       key_c_r_27_31, key_c_r_27_32, key_c_r_27_33, key_c_r_27_34, key_c_r_27_35, key_c_r_27_36, key_c_r_27_37, key_c_r_27_38, key_c_r_27_39, 
       key_c_r_27_4, key_c_r_27_40, key_c_r_27_41, key_c_r_27_42, key_c_r_27_43, key_c_r_27_44, key_c_r_27_45, key_c_r_27_46, key_c_r_27_47, 
       key_c_r_27_48, key_c_r_27_49, key_c_r_27_5, key_c_r_27_50, key_c_r_27_51, key_c_r_27_52, key_c_r_27_53, key_c_r_27_54, key_c_r_27_55, 
       key_c_r_27_6, key_c_r_27_7, key_c_r_27_8, key_c_r_27_9, key_c_r_28_0, key_c_r_28_1, key_c_r_28_10, key_c_r_28_11, key_c_r_28_12, 
       key_c_r_28_13, key_c_r_28_14, key_c_r_28_15, key_c_r_28_16, key_c_r_28_17, key_c_r_28_18, key_c_r_28_19, key_c_r_28_2, key_c_r_28_20, 
       key_c_r_28_21, key_c_r_28_22, key_c_r_28_23, key_c_r_28_24, key_c_r_28_25, key_c_r_28_26, key_c_r_28_27, key_c_r_28_28, key_c_r_28_29, 
       key_c_r_28_3, key_c_r_28_30, key_c_r_28_31, key_c_r_28_32, key_c_r_28_33, key_c_r_28_34, key_c_r_28_35, key_c_r_28_36, key_c_r_28_37, 
       key_c_r_28_38, key_c_r_28_39, key_c_r_28_4, key_c_r_28_40, key_c_r_28_41, key_c_r_28_42, key_c_r_28_43, key_c_r_28_44, key_c_r_28_45, 
       key_c_r_28_46, key_c_r_28_47, key_c_r_28_48, key_c_r_28_49, key_c_r_28_5, key_c_r_28_50, key_c_r_28_51, key_c_r_28_52, key_c_r_28_53, 
       key_c_r_28_54, key_c_r_28_55, key_c_r_28_6, key_c_r_28_7, key_c_r_28_8, key_c_r_28_9, key_c_r_29_0, key_c_r_29_1, key_c_r_29_10, 
       key_c_r_29_11, key_c_r_29_12, key_c_r_29_13, key_c_r_29_14, key_c_r_29_15, key_c_r_29_16, key_c_r_29_17, key_c_r_29_18, key_c_r_29_19, 
       key_c_r_29_2, key_c_r_29_20, key_c_r_29_21, key_c_r_29_22, key_c_r_29_23, key_c_r_29_24, key_c_r_29_25, key_c_r_29_26, key_c_r_29_27, 
       key_c_r_29_28, key_c_r_29_29, key_c_r_29_3, key_c_r_29_30, key_c_r_29_31, key_c_r_29_32, key_c_r_29_33, key_c_r_29_34, key_c_r_29_35, 
       key_c_r_29_36, key_c_r_29_37, key_c_r_29_38, key_c_r_29_39, key_c_r_29_4, key_c_r_29_40, key_c_r_29_41, key_c_r_29_42, key_c_r_29_43, 
       key_c_r_29_44, key_c_r_29_45, key_c_r_29_46, key_c_r_29_47, key_c_r_29_48, key_c_r_29_49, key_c_r_29_5, key_c_r_29_50, key_c_r_29_51, 
       key_c_r_29_52, key_c_r_29_53, key_c_r_29_54, key_c_r_29_55, key_c_r_29_6, key_c_r_29_7, key_c_r_29_8, key_c_r_29_9, key_c_r_2_0, 
       key_c_r_2_1, key_c_r_2_10, key_c_r_2_11, key_c_r_2_12, key_c_r_2_13, key_c_r_2_14, key_c_r_2_15, key_c_r_2_16, key_c_r_2_17, 
       key_c_r_2_18, key_c_r_2_19, key_c_r_2_2, key_c_r_2_20, key_c_r_2_21, key_c_r_2_22, key_c_r_2_23, key_c_r_2_24, key_c_r_2_25, 
       key_c_r_2_26, key_c_r_2_27, key_c_r_2_28, key_c_r_2_29, key_c_r_2_3, key_c_r_2_30, key_c_r_2_31, key_c_r_2_32, key_c_r_2_33, 
       key_c_r_2_34, key_c_r_2_35, key_c_r_2_36, key_c_r_2_37, key_c_r_2_38, key_c_r_2_39, key_c_r_2_4, key_c_r_2_40, key_c_r_2_41, 
       key_c_r_2_42, key_c_r_2_43, key_c_r_2_44, key_c_r_2_45, key_c_r_2_46, key_c_r_2_47, key_c_r_2_48, key_c_r_2_49, key_c_r_2_5, 
       key_c_r_2_50, key_c_r_2_51, key_c_r_2_52, key_c_r_2_53, key_c_r_2_54, key_c_r_2_55, key_c_r_2_6, key_c_r_2_7, key_c_r_2_8, 
       key_c_r_2_9, key_c_r_30_0, key_c_r_30_1, key_c_r_30_10, key_c_r_30_11, key_c_r_30_12, key_c_r_30_13, key_c_r_30_14, key_c_r_30_15, 
       key_c_r_30_16, key_c_r_30_17, key_c_r_30_18, key_c_r_30_19, key_c_r_30_2, key_c_r_30_20, key_c_r_30_21, key_c_r_30_22, key_c_r_30_23, 
       key_c_r_30_24, key_c_r_30_25, key_c_r_30_26, key_c_r_30_27, key_c_r_30_28, key_c_r_30_29, key_c_r_30_3, key_c_r_30_30, key_c_r_30_31, 
       key_c_r_30_32, key_c_r_30_33, key_c_r_30_34, key_c_r_30_35, key_c_r_30_36, key_c_r_30_37, key_c_r_30_38, key_c_r_30_39, key_c_r_30_4, 
       key_c_r_30_40, key_c_r_30_41, key_c_r_30_42, key_c_r_30_43, key_c_r_30_44, key_c_r_30_45, key_c_r_30_46, key_c_r_30_47, key_c_r_30_48, 
       key_c_r_30_49, key_c_r_30_5, key_c_r_30_50, key_c_r_30_51, key_c_r_30_52, key_c_r_30_53, key_c_r_30_54, key_c_r_30_55, key_c_r_30_6, 
       key_c_r_30_7, key_c_r_30_8, key_c_r_30_9, key_c_r_31_0, key_c_r_31_1, key_c_r_31_10, key_c_r_31_11, key_c_r_31_12, key_c_r_31_13, 
       key_c_r_31_14, key_c_r_31_15, key_c_r_31_16, key_c_r_31_17, key_c_r_31_18, key_c_r_31_19, key_c_r_31_2, key_c_r_31_20, key_c_r_31_21, 
       key_c_r_31_22, key_c_r_31_23, key_c_r_31_24, key_c_r_31_25, key_c_r_31_26, key_c_r_31_27, key_c_r_31_28, key_c_r_31_29, key_c_r_31_3, 
       key_c_r_31_30, key_c_r_31_31, key_c_r_31_32, key_c_r_31_33, key_c_r_31_34, key_c_r_31_35, key_c_r_31_36, key_c_r_31_37, key_c_r_31_38, 
       key_c_r_31_39, key_c_r_31_4, key_c_r_31_40, key_c_r_31_41, key_c_r_31_42, key_c_r_31_43, key_c_r_31_44, key_c_r_31_45, key_c_r_31_46, 
       key_c_r_31_47, key_c_r_31_48, key_c_r_31_49, key_c_r_31_5, key_c_r_31_50, key_c_r_31_51, key_c_r_31_52, key_c_r_31_53, key_c_r_31_54, 
       key_c_r_31_55, key_c_r_31_6, key_c_r_31_7, key_c_r_31_8, key_c_r_31_9, key_c_r_32_0, key_c_r_32_1, key_c_r_32_10, key_c_r_32_11, 
       key_c_r_32_12, key_c_r_32_13, key_c_r_32_14, key_c_r_32_15, key_c_r_32_16, key_c_r_32_17, key_c_r_32_18, key_c_r_32_19, key_c_r_32_2, 
       key_c_r_32_20, key_c_r_32_21, key_c_r_32_22, key_c_r_32_23, key_c_r_32_24, key_c_r_32_25, key_c_r_32_26, key_c_r_32_27, key_c_r_32_28, 
       key_c_r_32_29, key_c_r_32_3, key_c_r_32_30, key_c_r_32_31, key_c_r_32_32, key_c_r_32_33, key_c_r_32_34, key_c_r_32_35, key_c_r_32_36, 
       key_c_r_32_37, key_c_r_32_38, key_c_r_32_39, key_c_r_32_4, key_c_r_32_40, key_c_r_32_41, key_c_r_32_42, key_c_r_32_43, key_c_r_32_44, 
       key_c_r_32_45, key_c_r_32_46, key_c_r_32_47, key_c_r_32_48, key_c_r_32_49, key_c_r_32_5, key_c_r_32_50, key_c_r_32_51, key_c_r_32_52, 
       key_c_r_32_53, key_c_r_32_54, key_c_r_32_55, key_c_r_32_6, key_c_r_32_7, key_c_r_32_8, key_c_r_32_9, key_c_r_33_0, key_c_r_33_1, 
       key_c_r_33_10, key_c_r_33_11, key_c_r_33_12, key_c_r_33_13, key_c_r_33_14, key_c_r_33_15, key_c_r_33_16, key_c_r_33_17, key_c_r_33_18, 
       key_c_r_33_19, key_c_r_33_2, key_c_r_33_20, key_c_r_33_21, key_c_r_33_22, key_c_r_33_23, key_c_r_33_24, key_c_r_33_25, key_c_r_33_26, 
       key_c_r_33_27, key_c_r_33_28, key_c_r_33_29, key_c_r_33_3, key_c_r_33_30, key_c_r_33_31, key_c_r_33_32, key_c_r_33_33, key_c_r_33_34, 
       key_c_r_33_35, key_c_r_33_36, key_c_r_33_37, key_c_r_33_38, key_c_r_33_39, key_c_r_33_4, key_c_r_33_40, key_c_r_33_41, key_c_r_33_42, 
       key_c_r_33_43, key_c_r_33_44, key_c_r_33_45, key_c_r_33_46, key_c_r_33_47, key_c_r_33_48, key_c_r_33_49, key_c_r_33_5, key_c_r_33_50, 
       key_c_r_33_51, key_c_r_33_52, key_c_r_33_53, key_c_r_33_54, key_c_r_33_55, key_c_r_33_6, key_c_r_33_7, key_c_r_33_8, key_c_r_33_9, 
       key_c_r_3_0, key_c_r_3_1, key_c_r_3_10, key_c_r_3_11, key_c_r_3_12, key_c_r_3_13, key_c_r_3_14, key_c_r_3_15, key_c_r_3_16, 
       key_c_r_3_17, key_c_r_3_18, key_c_r_3_19, key_c_r_3_2, key_c_r_3_20, key_c_r_3_21, key_c_r_3_22, key_c_r_3_23, key_c_r_3_24, 
       key_c_r_3_25, key_c_r_3_26, key_c_r_3_27, key_c_r_3_28, key_c_r_3_29, key_c_r_3_3, key_c_r_3_30, key_c_r_3_31, key_c_r_3_32, 
       key_c_r_3_33, key_c_r_3_34, key_c_r_3_35, key_c_r_3_36, key_c_r_3_37, key_c_r_3_38, key_c_r_3_39, key_c_r_3_4, key_c_r_3_40, 
       key_c_r_3_41, key_c_r_3_42, key_c_r_3_43, key_c_r_3_44, key_c_r_3_45, key_c_r_3_46, key_c_r_3_47, key_c_r_3_48, key_c_r_3_49, 
       key_c_r_3_5, key_c_r_3_50, key_c_r_3_51, key_c_r_3_52, key_c_r_3_53, key_c_r_3_54, key_c_r_3_55, key_c_r_3_6, key_c_r_3_7, 
       key_c_r_3_8, key_c_r_3_9, key_c_r_4_0, key_c_r_4_1, key_c_r_4_10, key_c_r_4_11, key_c_r_4_12, key_c_r_4_13, key_c_r_4_14, 
       key_c_r_4_15, key_c_r_4_16, key_c_r_4_17, key_c_r_4_18, key_c_r_4_19, key_c_r_4_2, key_c_r_4_20, key_c_r_4_21, key_c_r_4_22, 
       key_c_r_4_23, key_c_r_4_24, key_c_r_4_25, key_c_r_4_26, key_c_r_4_27, key_c_r_4_28, key_c_r_4_29, key_c_r_4_3, key_c_r_4_30, 
       key_c_r_4_31, key_c_r_4_32, key_c_r_4_33, key_c_r_4_34, key_c_r_4_35, key_c_r_4_36, key_c_r_4_37, key_c_r_4_38, key_c_r_4_39, 
       key_c_r_4_4, key_c_r_4_40, key_c_r_4_41, key_c_r_4_42, key_c_r_4_43, key_c_r_4_44, key_c_r_4_45, key_c_r_4_46, key_c_r_4_47, 
       key_c_r_4_48, key_c_r_4_49, key_c_r_4_5, key_c_r_4_50, key_c_r_4_51, key_c_r_4_52, key_c_r_4_53, key_c_r_4_54, key_c_r_4_55, 
       key_c_r_4_6, key_c_r_4_7, key_c_r_4_8, key_c_r_4_9, key_c_r_5_0, key_c_r_5_1, key_c_r_5_10, key_c_r_5_11, key_c_r_5_12, 
       key_c_r_5_13, key_c_r_5_14, key_c_r_5_15, key_c_r_5_16, key_c_r_5_17, key_c_r_5_18, key_c_r_5_19, key_c_r_5_2, key_c_r_5_20, 
       key_c_r_5_21, key_c_r_5_22, key_c_r_5_23, key_c_r_5_24, key_c_r_5_25, key_c_r_5_26, key_c_r_5_27, key_c_r_5_28, key_c_r_5_29, 
       key_c_r_5_3, key_c_r_5_30, key_c_r_5_31, key_c_r_5_32, key_c_r_5_33, key_c_r_5_34, key_c_r_5_35, key_c_r_5_36, key_c_r_5_37, 
       key_c_r_5_38, key_c_r_5_39, key_c_r_5_4, key_c_r_5_40, key_c_r_5_41, key_c_r_5_42, key_c_r_5_43, key_c_r_5_44, key_c_r_5_45, 
       key_c_r_5_46, key_c_r_5_47, key_c_r_5_48, key_c_r_5_49, key_c_r_5_5, key_c_r_5_50, key_c_r_5_51, key_c_r_5_52, key_c_r_5_53, 
       key_c_r_5_54, key_c_r_5_55, key_c_r_5_6, key_c_r_5_7, key_c_r_5_8, key_c_r_5_9, key_c_r_6_0, key_c_r_6_1, key_c_r_6_10, 
       key_c_r_6_11, key_c_r_6_12, key_c_r_6_13, key_c_r_6_14, key_c_r_6_15, key_c_r_6_16, key_c_r_6_17, key_c_r_6_18, key_c_r_6_19, 
       key_c_r_6_2, key_c_r_6_20, key_c_r_6_21, key_c_r_6_22, key_c_r_6_23, key_c_r_6_24, key_c_r_6_25, key_c_r_6_26, key_c_r_6_27, 
       key_c_r_6_28, key_c_r_6_29, key_c_r_6_3, key_c_r_6_30, key_c_r_6_31, key_c_r_6_32, key_c_r_6_33, key_c_r_6_34, key_c_r_6_35, 
       key_c_r_6_36, key_c_r_6_37, key_c_r_6_38, key_c_r_6_39, key_c_r_6_4, key_c_r_6_40, key_c_r_6_41, key_c_r_6_42, key_c_r_6_43, 
       key_c_r_6_44, key_c_r_6_45, key_c_r_6_46, key_c_r_6_47, key_c_r_6_48, key_c_r_6_49, key_c_r_6_5, key_c_r_6_50, key_c_r_6_51, 
       key_c_r_6_52, key_c_r_6_53, key_c_r_6_54, key_c_r_6_55, key_c_r_6_6, key_c_r_6_7, key_c_r_6_8, key_c_r_6_9, key_c_r_7_0, 
       key_c_r_7_1, key_c_r_7_10, key_c_r_7_11, key_c_r_7_12, key_c_r_7_13, key_c_r_7_14, key_c_r_7_15, key_c_r_7_16, key_c_r_7_17, 
       key_c_r_7_18, key_c_r_7_19, key_c_r_7_2, key_c_r_7_20, key_c_r_7_21, key_c_r_7_22, key_c_r_7_23, key_c_r_7_24, key_c_r_7_25, 
       key_c_r_7_26, key_c_r_7_27, key_c_r_7_28, key_c_r_7_29, key_c_r_7_3, key_c_r_7_30, key_c_r_7_31, key_c_r_7_32, key_c_r_7_33, 
       key_c_r_7_34, key_c_r_7_35, key_c_r_7_36, key_c_r_7_37, key_c_r_7_38, key_c_r_7_39, key_c_r_7_4, key_c_r_7_40, key_c_r_7_41, 
       key_c_r_7_42, key_c_r_7_43, key_c_r_7_44, key_c_r_7_45, key_c_r_7_46, key_c_r_7_47, key_c_r_7_48, key_c_r_7_49, key_c_r_7_5, 
       key_c_r_7_50, key_c_r_7_51, key_c_r_7_52, key_c_r_7_53, key_c_r_7_54, key_c_r_7_55, key_c_r_7_6, key_c_r_7_7, key_c_r_7_8, 
       key_c_r_7_9, key_c_r_8_0, key_c_r_8_1, key_c_r_8_10, key_c_r_8_11, key_c_r_8_12, key_c_r_8_13, key_c_r_8_14, key_c_r_8_15, 
       key_c_r_8_16, key_c_r_8_17, key_c_r_8_18, key_c_r_8_19, key_c_r_8_2, key_c_r_8_20, key_c_r_8_21, key_c_r_8_22, key_c_r_8_23, 
       key_c_r_8_24, key_c_r_8_25, key_c_r_8_26, key_c_r_8_27, key_c_r_8_28, key_c_r_8_29, key_c_r_8_3, key_c_r_8_30, key_c_r_8_31, 
       key_c_r_8_32, key_c_r_8_33, key_c_r_8_34, key_c_r_8_35, key_c_r_8_36, key_c_r_8_37, key_c_r_8_38, key_c_r_8_39, key_c_r_8_4, 
       key_c_r_8_40, key_c_r_8_41, key_c_r_8_42, key_c_r_8_43, key_c_r_8_44, key_c_r_8_45, key_c_r_8_46, key_c_r_8_47, key_c_r_8_48, 
       key_c_r_8_49, key_c_r_8_5, key_c_r_8_50, key_c_r_8_51, key_c_r_8_52, key_c_r_8_53, key_c_r_8_54, key_c_r_8_55, key_c_r_8_6, 
       key_c_r_8_7, key_c_r_8_8, key_c_r_8_9, key_c_r_9_0, key_c_r_9_1, key_c_r_9_10, key_c_r_9_11, key_c_r_9_12, key_c_r_9_13, 
       key_c_r_9_14, key_c_r_9_15, key_c_r_9_16, key_c_r_9_17, key_c_r_9_18, key_c_r_9_19, key_c_r_9_2, key_c_r_9_20, key_c_r_9_21, 
       key_c_r_9_22, key_c_r_9_23, key_c_r_9_24, key_c_r_9_25, key_c_r_9_26, key_c_r_9_27, key_c_r_9_28, key_c_r_9_29, key_c_r_9_3, 
       key_c_r_9_30, key_c_r_9_31, key_c_r_9_32, key_c_r_9_33, key_c_r_9_34, key_c_r_9_35, key_c_r_9_36, key_c_r_9_37, key_c_r_9_38, 
       key_c_r_9_39, key_c_r_9_4, key_c_r_9_40, key_c_r_9_41, key_c_r_9_42, key_c_r_9_43, key_c_r_9_44, key_c_r_9_45, key_c_r_9_46, 
       key_c_r_9_47, key_c_r_9_48, key_c_r_9_49, key_c_r_9_5, key_c_r_9_50, key_c_r_9_51, key_c_r_9_52, key_c_r_9_53, key_c_r_9_54, 
       key_c_r_9_55, key_c_r_9_6, key_c_r_9_7, key_c_r_9_8, key_c_r_9_9, n1, n10, n100, n101, 
       n102, n103, n104, n105, n106, n107, n108, n109, n11, 
       n110, n111, n112, n114, n115, n12, n13, n14, n15, 
       n16, n17, n18, n19, n2, n20, n21, n22, n23, 
       n24, n25, n26, n27, n28, n29, n3, n30, n31, 
       n32, n33, n34, n35, n36, n37, n38, n39, n4, 
       n40, n41, n42, n43, n44, n45, n46, n47, n48, 
       n49, n5, n50, n51, n52, n53, n54, n55, n56, 
       n57, n58, n59, n6, n60, n61, n62, n63, n64, 
       n65, n66, n67, n68, n69, n7, n70, n71, n72, 
       n73, n74, n75, n76, n77, n78, n79, n8, n80, 
       n81, n82, n83, n84, n85, n86, n87, n88, n89, 
       n9, n90, n91, n92, n93, n94, n95, n96, n97, 
       n98, n99, stage1_out_0, stage1_out_1, stage1_out_10, stage1_out_11, stage1_out_12, stage1_out_13, stage1_out_14, 
       stage1_out_15, stage1_out_16, stage1_out_17, stage1_out_18, stage1_out_19, stage1_out_2, stage1_out_20, stage1_out_21, stage1_out_22, 
       stage1_out_23, stage1_out_24, stage1_out_25, stage1_out_26, stage1_out_27, stage1_out_28, stage1_out_29, stage1_out_3, stage1_out_30, 
       stage1_out_31, stage1_out_32, stage1_out_33, stage1_out_34, stage1_out_35, stage1_out_36, stage1_out_37, stage1_out_38, stage1_out_39, 
       stage1_out_4, stage1_out_40, stage1_out_41, stage1_out_42, stage1_out_43, stage1_out_44, stage1_out_45, stage1_out_46, stage1_out_47, 
       stage1_out_48, stage1_out_49, stage1_out_5, stage1_out_50, stage1_out_51, stage1_out_52, stage1_out_53, stage1_out_54, stage1_out_55, 
       stage1_out_56, stage1_out_57, stage1_out_58, stage1_out_59, stage1_out_6, stage1_out_60, stage1_out_61, stage1_out_62, stage1_out_63, 
       stage1_out_7, stage1_out_8, stage1_out_9, stage2_out_0, stage2_out_1, stage2_out_10, stage2_out_11, stage2_out_12, stage2_out_13, 
       stage2_out_14, stage2_out_15, stage2_out_16, stage2_out_17, stage2_out_18, stage2_out_19, stage2_out_2, stage2_out_20, stage2_out_21, 
       stage2_out_22, stage2_out_23, stage2_out_24, stage2_out_25, stage2_out_26, stage2_out_27, stage2_out_28, stage2_out_29, stage2_out_3, 
       stage2_out_30, stage2_out_31, stage2_out_32, stage2_out_33, stage2_out_34, stage2_out_35, stage2_out_36, stage2_out_37, stage2_out_38, 
       stage2_out_39, stage2_out_4, stage2_out_40, stage2_out_41, stage2_out_42, stage2_out_43, stage2_out_44, stage2_out_45, stage2_out_46, 
       stage2_out_47, stage2_out_48, stage2_out_49, stage2_out_5, stage2_out_50, stage2_out_51, stage2_out_52, stage2_out_53, stage2_out_54, 
       stage2_out_55, stage2_out_56, stage2_out_57, stage2_out_58, stage2_out_59, stage2_out_6, stage2_out_60, stage2_out_61, stage2_out_62, 
       stage2_out_63, stage2_out_7, stage2_out_8, stage2_out_9, u0_key_r_15, u0_uk_K_r0_0, u0_uk_K_r0_1, u0_uk_K_r0_10, u0_uk_K_r0_12, 
       u0_uk_K_r0_13, u0_uk_K_r0_14, u0_uk_K_r0_16, u0_uk_K_r0_17, u0_uk_K_r0_18, u0_uk_K_r0_20, u0_uk_K_r0_21, u0_uk_K_r0_23, u0_uk_K_r0_24, 
       u0_uk_K_r0_26, u0_uk_K_r0_27, u0_uk_K_r0_29, u0_uk_K_r0_3, u0_uk_K_r0_30, u0_uk_K_r0_33, u0_uk_K_r0_35, u0_uk_K_r0_37, u0_uk_K_r0_38, 
       u0_uk_K_r0_39, u0_uk_K_r0_4, u0_uk_K_r0_40, u0_uk_K_r0_41, u0_uk_K_r0_42, u0_uk_K_r0_43, u0_uk_K_r0_44, u0_uk_K_r0_45, u0_uk_K_r0_46, 
       u0_uk_K_r0_48, u0_uk_K_r0_5, u0_uk_K_r0_50, u0_uk_K_r0_51, u0_uk_K_r0_53, u0_uk_K_r0_54, u0_uk_K_r0_6, u0_uk_K_r0_8, u0_uk_K_r0_9, 
       u0_uk_K_r10_0, u0_uk_K_r10_1, u0_uk_K_r10_11, u0_uk_K_r10_12, u0_uk_K_r10_13, u0_uk_K_r10_15, u0_uk_K_r10_17, u0_uk_K_r10_2, u0_uk_K_r10_20, 
       u0_uk_K_r10_21, u0_uk_K_r10_22, u0_uk_K_r10_24, u0_uk_K_r10_26, u0_uk_K_r10_29, u0_uk_K_r10_3, u0_uk_K_r10_30, u0_uk_K_r10_31, u0_uk_K_r10_33, 
       u0_uk_K_r10_35, u0_uk_K_r10_36, u0_uk_K_r10_38, u0_uk_K_r10_4, u0_uk_K_r10_40, u0_uk_K_r10_45, u0_uk_K_r10_46, u0_uk_K_r10_49, u0_uk_K_r10_5, 
       u0_uk_K_r10_50, u0_uk_K_r10_51, u0_uk_K_r10_52, u0_uk_K_r10_53, u0_uk_K_r10_54, u0_uk_K_r10_55, u0_uk_K_r10_6, u0_uk_K_r10_7, u0_uk_K_r10_8, 
       u0_uk_K_r11_0, u0_uk_K_r11_1, u0_uk_K_r11_12, u0_uk_K_r11_13, u0_uk_K_r11_14, u0_uk_K_r11_15, u0_uk_K_r11_16, u0_uk_K_r11_18, u0_uk_K_r11_2, 
       u0_uk_K_r11_22, u0_uk_K_r11_23, u0_uk_K_r11_3, u0_uk_K_r11_30, u0_uk_K_r11_31, u0_uk_K_r11_32, u0_uk_K_r11_35, u0_uk_K_r11_36, u0_uk_K_r11_37, 
       u0_uk_K_r11_38, u0_uk_K_r11_40, u0_uk_K_r11_41, u0_uk_K_r11_42, u0_uk_K_r11_43, u0_uk_K_r11_44, u0_uk_K_r11_45, u0_uk_K_r11_49, u0_uk_K_r11_5, 
       u0_uk_K_r11_50, u0_uk_K_r11_51, u0_uk_K_r11_52, u0_uk_K_r11_55, u0_uk_K_r11_7, u0_uk_K_r11_9, u0_uk_K_r12_0, u0_uk_K_r12_11, u0_uk_K_r12_12, 
       u0_uk_K_r12_13, u0_uk_K_r12_14, u0_uk_K_r12_17, u0_uk_K_r12_19, u0_uk_K_r12_2, u0_uk_K_r12_20, u0_uk_K_r12_22, u0_uk_K_r12_23, u0_uk_K_r12_24, 
       u0_uk_K_r12_26, u0_uk_K_r12_27, u0_uk_K_r12_28, u0_uk_K_r12_29, u0_uk_K_r12_3, u0_uk_K_r12_31, u0_uk_K_r12_32, u0_uk_K_r12_34, u0_uk_K_r12_35, 
       u0_uk_K_r12_37, u0_uk_K_r12_38, u0_uk_K_r12_39, u0_uk_K_r12_4, u0_uk_K_r12_40, u0_uk_K_r12_41, u0_uk_K_r12_43, u0_uk_K_r12_45, u0_uk_K_r12_46, 
       u0_uk_K_r12_48, u0_uk_K_r12_49, u0_uk_K_r12_5, u0_uk_K_r12_50, u0_uk_K_r12_51, u0_uk_K_r12_52, u0_uk_K_r12_53, u0_uk_K_r12_54, u0_uk_K_r12_55, 
       u0_uk_K_r12_6, u0_uk_K_r12_8, u0_uk_K_r12_9, u0_uk_K_r13_1, u0_uk_K_r13_10, u0_uk_K_r13_11, u0_uk_K_r13_12, u0_uk_K_r13_14, u0_uk_K_r13_15, 
       u0_uk_K_r13_16, u0_uk_K_r13_18, u0_uk_K_r13_20, u0_uk_K_r13_21, u0_uk_K_r13_24, u0_uk_K_r13_26, u0_uk_K_r13_27, u0_uk_K_r13_28, u0_uk_K_r13_29, 
       u0_uk_K_r13_3, u0_uk_K_r13_30, u0_uk_K_r13_31, u0_uk_K_r13_33, u0_uk_K_r13_34, u0_uk_K_r13_36, u0_uk_K_r13_37, u0_uk_K_r13_39, u0_uk_K_r13_40, 
       u0_uk_K_r13_41, u0_uk_K_r13_42, u0_uk_K_r13_43, u0_uk_K_r13_45, u0_uk_K_r13_46, u0_uk_K_r13_47, u0_uk_K_r13_48, u0_uk_K_r13_49, u0_uk_K_r13_5, 
       u0_uk_K_r13_50, u0_uk_K_r13_51, u0_uk_K_r13_52, u0_uk_K_r13_53, u0_uk_K_r13_54, u0_uk_K_r13_6, u0_uk_K_r13_7, u0_uk_K_r13_8, u0_uk_K_r13_9, 
       u0_uk_K_r14_23, u0_uk_K_r14_38, u0_uk_K_r14_42, u0_uk_K_r1_0, u0_uk_K_r1_1, u0_uk_K_r1_11, u0_uk_K_r1_12, u0_uk_K_r1_13, u0_uk_K_r1_14, 
       u0_uk_K_r1_19, u0_uk_K_r1_2, u0_uk_K_r1_20, u0_uk_K_r1_23, u0_uk_K_r1_24, u0_uk_K_r1_25, u0_uk_K_r1_26, u0_uk_K_r1_27, u0_uk_K_r1_28, 
       u0_uk_K_r1_29, u0_uk_K_r1_3, u0_uk_K_r1_30, u0_uk_K_r1_31, u0_uk_K_r1_32, u0_uk_K_r1_33, u0_uk_K_r1_34, u0_uk_K_r1_35, u0_uk_K_r1_37, 
       u0_uk_K_r1_38, u0_uk_K_r1_39, u0_uk_K_r1_4, u0_uk_K_r1_40, u0_uk_K_r1_43, u0_uk_K_r1_45, u0_uk_K_r1_46, u0_uk_K_r1_48, u0_uk_K_r1_49, 
       u0_uk_K_r1_5, u0_uk_K_r1_50, u0_uk_K_r1_51, u0_uk_K_r1_52, u0_uk_K_r1_53, u0_uk_K_r1_54, u0_uk_K_r1_55, u0_uk_K_r1_6, u0_uk_K_r1_8, 
       u0_uk_K_r1_9, u0_uk_K_r2_0, u0_uk_K_r2_1, u0_uk_K_r2_10, u0_uk_K_r2_11, u0_uk_K_r2_12, u0_uk_K_r2_14, u0_uk_K_r2_15, u0_uk_K_r2_17, 
       u0_uk_K_r2_19, u0_uk_K_r2_2, u0_uk_K_r2_21, u0_uk_K_r2_22, u0_uk_K_r2_23, u0_uk_K_r2_24, u0_uk_K_r2_3, u0_uk_K_r2_30, u0_uk_K_r2_32, 
       u0_uk_K_r2_34, u0_uk_K_r2_35, u0_uk_K_r2_37, u0_uk_K_r2_38, u0_uk_K_r2_39, u0_uk_K_r2_40, u0_uk_K_r2_42, u0_uk_K_r2_43, u0_uk_K_r2_44, 
       u0_uk_K_r2_45, u0_uk_K_r2_47, u0_uk_K_r2_48, u0_uk_K_r2_49, u0_uk_K_r2_5, u0_uk_K_r2_51, u0_uk_K_r2_52, u0_uk_K_r2_54, u0_uk_K_r2_6, 
       u0_uk_K_r2_8, u0_uk_K_r2_9, u0_uk_K_r3_0, u0_uk_K_r3_1, u0_uk_K_r3_12, u0_uk_K_r3_13, u0_uk_K_r3_17, u0_uk_K_r3_18, u0_uk_K_r3_2, 
       u0_uk_K_r3_20, u0_uk_K_r3_21, u0_uk_K_r3_22, u0_uk_K_r3_23, u0_uk_K_r3_25, u0_uk_K_r3_26, u0_uk_K_r3_27, u0_uk_K_r3_28, u0_uk_K_r3_3, 
       u0_uk_K_r3_30, u0_uk_K_r3_31, u0_uk_K_r3_32, u0_uk_K_r3_33, u0_uk_K_r3_34, u0_uk_K_r3_36, u0_uk_K_r3_37, u0_uk_K_r3_39, u0_uk_K_r3_40, 
       u0_uk_K_r3_41, u0_uk_K_r3_42, u0_uk_K_r3_43, u0_uk_K_r3_44, u0_uk_K_r3_45, u0_uk_K_r3_46, u0_uk_K_r3_48, u0_uk_K_r3_49, u0_uk_K_r3_5, 
       u0_uk_K_r3_50, u0_uk_K_r3_51, u0_uk_K_r3_53, u0_uk_K_r3_54, u0_uk_K_r3_55, u0_uk_K_r3_6, u0_uk_K_r3_7, u0_uk_K_r3_8, u0_uk_K_r4_1, 
       u0_uk_K_r4_10, u0_uk_K_r4_12, u0_uk_K_r4_13, u0_uk_K_r4_14, u0_uk_K_r4_15, u0_uk_K_r4_16, u0_uk_K_r4_17, u0_uk_K_r4_18, u0_uk_K_r4_19, 
       u0_uk_K_r4_2, u0_uk_K_r4_20, u0_uk_K_r4_21, u0_uk_K_r4_22, u0_uk_K_r4_24, u0_uk_K_r4_25, u0_uk_K_r4_26, u0_uk_K_r4_27, u0_uk_K_r4_28, 
       u0_uk_K_r4_29, u0_uk_K_r4_30, u0_uk_K_r4_32, u0_uk_K_r4_34, u0_uk_K_r4_36, u0_uk_K_r4_37, u0_uk_K_r4_39, u0_uk_K_r4_40, u0_uk_K_r4_42, 
       u0_uk_K_r4_43, u0_uk_K_r4_44, u0_uk_K_r4_45, u0_uk_K_r4_46, u0_uk_K_r4_50, u0_uk_K_r4_51, u0_uk_K_r4_52, u0_uk_K_r4_53, u0_uk_K_r4_6, 
       u0_uk_K_r4_7, u0_uk_K_r4_8, u0_uk_K_r4_9, u0_uk_K_r5_11, u0_uk_K_r5_12, u0_uk_K_r5_14, u0_uk_K_r5_15, u0_uk_K_r5_2, u0_uk_K_r5_20, 
       u0_uk_K_r5_22, u0_uk_K_r5_24, u0_uk_K_r5_25, u0_uk_K_r5_27, u0_uk_K_r5_28, u0_uk_K_r5_29, u0_uk_K_r5_3, u0_uk_K_r5_30, u0_uk_K_r5_31, 
       u0_uk_K_r5_33, u0_uk_K_r5_34, u0_uk_K_r5_35, u0_uk_K_r5_36, u0_uk_K_r5_38, u0_uk_K_r5_42, u0_uk_K_r5_44, u0_uk_K_r5_45, u0_uk_K_r5_46, 
       u0_uk_K_r5_47, u0_uk_K_r5_49, u0_uk_K_r5_50, u0_uk_K_r5_52, u0_uk_K_r5_53, u0_uk_K_r5_54, u0_uk_K_r5_55, u0_uk_K_r5_6, u0_uk_K_r5_7, 
       u0_uk_K_r5_9, u0_uk_K_r6_1, u0_uk_K_r6_11, u0_uk_K_r6_12, u0_uk_K_r6_13, u0_uk_K_r6_15, u0_uk_K_r6_16, u0_uk_K_r6_17, u0_uk_K_r6_18, 
       u0_uk_K_r6_2, u0_uk_K_r6_20, u0_uk_K_r6_23, u0_uk_K_r6_24, u0_uk_K_r6_25, u0_uk_K_r6_28, u0_uk_K_r6_30, u0_uk_K_r6_32, u0_uk_K_r6_33, 
       u0_uk_K_r6_35, u0_uk_K_r6_36, u0_uk_K_r6_38, u0_uk_K_r6_39, u0_uk_K_r6_4, u0_uk_K_r6_40, u0_uk_K_r6_41, u0_uk_K_r6_42, u0_uk_K_r6_43, 
       u0_uk_K_r6_44, u0_uk_K_r6_45, u0_uk_K_r6_47, u0_uk_K_r6_48, u0_uk_K_r6_49, u0_uk_K_r6_5, u0_uk_K_r6_50, u0_uk_K_r6_52, u0_uk_K_r6_54, 
       u0_uk_K_r6_6, u0_uk_K_r6_8, u0_uk_K_r6_9, u0_uk_K_r7_10, u0_uk_K_r7_11, u0_uk_K_r7_12, u0_uk_K_r7_14, u0_uk_K_r7_16, u0_uk_K_r7_17, 
       u0_uk_K_r7_18, u0_uk_K_r7_19, u0_uk_K_r7_21, u0_uk_K_r7_28, u0_uk_K_r7_29, u0_uk_K_r7_3, u0_uk_K_r7_31, u0_uk_K_r7_33, u0_uk_K_r7_34, 
       u0_uk_K_r7_35, u0_uk_K_r7_36, u0_uk_K_r7_37, u0_uk_K_r7_38, u0_uk_K_r7_4, u0_uk_K_r7_40, u0_uk_K_r7_41, u0_uk_K_r7_42, u0_uk_K_r7_43, 
       u0_uk_K_r7_44, u0_uk_K_r7_45, u0_uk_K_r7_46, u0_uk_K_r7_47, u0_uk_K_r7_49, u0_uk_K_r7_5, u0_uk_K_r7_50, u0_uk_K_r7_51, u0_uk_K_r7_52, 
       u0_uk_K_r7_53, u0_uk_K_r7_54, u0_uk_K_r7_7, u0_uk_K_r8_0, u0_uk_K_r8_1, u0_uk_K_r8_10, u0_uk_K_r8_11, u0_uk_K_r8_12, u0_uk_K_r8_14, 
       u0_uk_K_r8_15, u0_uk_K_r8_18, u0_uk_K_r8_19, u0_uk_K_r8_20, u0_uk_K_r8_23, u0_uk_K_r8_24, u0_uk_K_r8_25, u0_uk_K_r8_26, u0_uk_K_r8_29, 
       u0_uk_K_r8_3, u0_uk_K_r8_30, u0_uk_K_r8_31, u0_uk_K_r8_33, u0_uk_K_r8_34, u0_uk_K_r8_35, u0_uk_K_r8_36, u0_uk_K_r8_38, u0_uk_K_r8_39, 
       u0_uk_K_r8_4, u0_uk_K_r8_42, u0_uk_K_r8_45, u0_uk_K_r8_46, u0_uk_K_r8_47, u0_uk_K_r8_48, u0_uk_K_r8_49, u0_uk_K_r8_5, u0_uk_K_r8_50, 
       u0_uk_K_r8_51, u0_uk_K_r8_53, u0_uk_K_r8_54, u0_uk_K_r8_55, u0_uk_K_r8_6, u0_uk_K_r8_7, u0_uk_K_r8_9, u0_uk_K_r9_11, u0_uk_K_r9_14, 
       u0_uk_K_r9_16, u0_uk_K_r9_17, u0_uk_K_r9_2, u0_uk_K_r9_20, u0_uk_K_r9_21, u0_uk_K_r9_24, u0_uk_K_r9_26, u0_uk_K_r9_28, u0_uk_K_r9_29, 
       u0_uk_K_r9_3, u0_uk_K_r9_32, u0_uk_K_r9_34, u0_uk_K_r9_36, u0_uk_K_r9_37, u0_uk_K_r9_39, u0_uk_K_r9_4, u0_uk_K_r9_40, u0_uk_K_r9_41, 
       u0_uk_K_r9_42, u0_uk_K_r9_43, u0_uk_K_r9_44, u0_uk_K_r9_46, u0_uk_K_r9_47, u0_uk_K_r9_50, u0_uk_K_r9_51, u0_uk_K_r9_52, u0_uk_K_r9_53, 
       u0_uk_K_r9_54, u0_uk_K_r9_55, u0_uk_K_r9_8, u0_uk_n1013, u0_uk_n1023, u0_uk_n114, u0_uk_n125, u0_uk_n133, u0_uk_n138, 
       u0_uk_n158, u0_uk_n160, u0_uk_n2, u0_uk_n236, u0_uk_n270, u0_uk_n284, u0_uk_n287, u0_uk_n295, u0_uk_n302, 
       u0_uk_n317, u0_uk_n334, u0_uk_n360, u0_uk_n416, u0_uk_n422, u0_uk_n431, u0_uk_n444, u0_uk_n449, u0_uk_n452, 
       u0_uk_n461, u0_uk_n469, u0_uk_n47, u0_uk_n470, u0_uk_n474, u0_uk_n477, u0_uk_n478, u0_uk_n487, u0_uk_n492, 
       u0_uk_n495, u0_uk_n533, u0_uk_n541, u0_uk_n548, u0_uk_n556, u0_uk_n572, u0_uk_n585, u0_uk_n591, u0_uk_n595, 
       u0_uk_n602, u0_uk_n617, u0_uk_n618, u0_uk_n70, u0_uk_n71, u0_uk_n724, u0_uk_n738, u0_uk_n74, u0_uk_n76, 
       u0_uk_n796, u0_uk_n812, u0_uk_n817, u0_uk_n820, u0_uk_n830, u0_uk_n852, u0_uk_n854, u0_uk_n928, u0_uk_n937, 
       u0_uk_n967, u0_uk_n970, u1_uk_K_r0_0, u1_uk_K_r0_1, u1_uk_K_r0_10, u1_uk_K_r0_12, u1_uk_K_r0_14, u1_uk_K_r0_16, u1_uk_K_r0_18, 
       u1_uk_K_r0_20, u1_uk_K_r0_21, u1_uk_K_r0_23, u1_uk_K_r0_24, u1_uk_K_r0_26, u1_uk_K_r0_27, u1_uk_K_r0_29, u1_uk_K_r0_3, u1_uk_K_r0_30, 
       u1_uk_K_r0_33, u1_uk_K_r0_35, u1_uk_K_r0_37, u1_uk_K_r0_38, u1_uk_K_r0_39, u1_uk_K_r0_4, u1_uk_K_r0_40, u1_uk_K_r0_41, u1_uk_K_r0_42, 
       u1_uk_K_r0_43, u1_uk_K_r0_44, u1_uk_K_r0_45, u1_uk_K_r0_46, u1_uk_K_r0_48, u1_uk_K_r0_5, u1_uk_K_r0_50, u1_uk_K_r0_51, u1_uk_K_r0_53, 
       u1_uk_K_r0_54, u1_uk_K_r0_6, u1_uk_K_r0_8, u1_uk_K_r0_9, u1_uk_K_r10_0, u1_uk_K_r10_1, u1_uk_K_r10_12, u1_uk_K_r10_13, u1_uk_K_r10_15, 
       u1_uk_K_r10_17, u1_uk_K_r10_2, u1_uk_K_r10_20, u1_uk_K_r10_21, u1_uk_K_r10_22, u1_uk_K_r10_24, u1_uk_K_r10_26, u1_uk_K_r10_29, u1_uk_K_r10_3, 
       u1_uk_K_r10_30, u1_uk_K_r10_31, u1_uk_K_r10_33, u1_uk_K_r10_35, u1_uk_K_r10_36, u1_uk_K_r10_38, u1_uk_K_r10_40, u1_uk_K_r10_45, u1_uk_K_r10_46, 
       u1_uk_K_r10_5, u1_uk_K_r10_50, u1_uk_K_r10_51, u1_uk_K_r10_53, u1_uk_K_r10_54, u1_uk_K_r10_55, u1_uk_K_r10_6, u1_uk_K_r10_7, u1_uk_K_r10_8, 
       u1_uk_K_r11_0, u1_uk_K_r11_1, u1_uk_K_r11_12, u1_uk_K_r11_13, u1_uk_K_r11_14, u1_uk_K_r11_15, u1_uk_K_r11_16, u1_uk_K_r11_18, u1_uk_K_r11_2, 
       u1_uk_K_r11_22, u1_uk_K_r11_23, u1_uk_K_r11_3, u1_uk_K_r11_30, u1_uk_K_r11_31, u1_uk_K_r11_32, u1_uk_K_r11_35, u1_uk_K_r11_36, u1_uk_K_r11_37, 
       u1_uk_K_r11_38, u1_uk_K_r11_40, u1_uk_K_r11_41, u1_uk_K_r11_42, u1_uk_K_r11_43, u1_uk_K_r11_44, u1_uk_K_r11_45, u1_uk_K_r11_49, u1_uk_K_r11_50, 
       u1_uk_K_r11_51, u1_uk_K_r11_52, u1_uk_K_r11_55, u1_uk_K_r11_9, u1_uk_K_r12_0, u1_uk_K_r12_11, u1_uk_K_r12_12, u1_uk_K_r12_13, u1_uk_K_r12_14, 
       u1_uk_K_r12_17, u1_uk_K_r12_19, u1_uk_K_r12_2, u1_uk_K_r12_20, u1_uk_K_r12_23, u1_uk_K_r12_24, u1_uk_K_r12_26, u1_uk_K_r12_27, u1_uk_K_r12_28, 
       u1_uk_K_r12_29, u1_uk_K_r12_3, u1_uk_K_r12_31, u1_uk_K_r12_32, u1_uk_K_r12_34, u1_uk_K_r12_35, u1_uk_K_r12_37, u1_uk_K_r12_38, u1_uk_K_r12_39, 
       u1_uk_K_r12_4, u1_uk_K_r12_40, u1_uk_K_r12_43, u1_uk_K_r12_45, u1_uk_K_r12_46, u1_uk_K_r12_48, u1_uk_K_r12_49, u1_uk_K_r12_5, u1_uk_K_r12_50, 
       u1_uk_K_r12_51, u1_uk_K_r12_52, u1_uk_K_r12_53, u1_uk_K_r12_54, u1_uk_K_r12_55, u1_uk_K_r12_6, u1_uk_K_r12_8, u1_uk_K_r12_9, u1_uk_K_r13_1, 
       u1_uk_K_r13_10, u1_uk_K_r13_11, u1_uk_K_r13_12, u1_uk_K_r13_14, u1_uk_K_r13_15, u1_uk_K_r13_16, u1_uk_K_r13_18, u1_uk_K_r13_20, u1_uk_K_r13_21, 
       u1_uk_K_r13_24, u1_uk_K_r13_26, u1_uk_K_r13_27, u1_uk_K_r13_28, u1_uk_K_r13_29, u1_uk_K_r13_3, u1_uk_K_r13_30, u1_uk_K_r13_33, u1_uk_K_r13_34, 
       u1_uk_K_r13_37, u1_uk_K_r13_39, u1_uk_K_r13_40, u1_uk_K_r13_41, u1_uk_K_r13_42, u1_uk_K_r13_43, u1_uk_K_r13_45, u1_uk_K_r13_46, u1_uk_K_r13_47, 
       u1_uk_K_r13_48, u1_uk_K_r13_49, u1_uk_K_r13_5, u1_uk_K_r13_50, u1_uk_K_r13_51, u1_uk_K_r13_52, u1_uk_K_r13_53, u1_uk_K_r13_54, u1_uk_K_r13_6, 
       u1_uk_K_r13_7, u1_uk_K_r13_8, u1_uk_K_r13_9, u1_uk_K_r1_0, u1_uk_K_r1_1, u1_uk_K_r1_11, u1_uk_K_r1_12, u1_uk_K_r1_13, u1_uk_K_r1_14, 
       u1_uk_K_r1_19, u1_uk_K_r1_2, u1_uk_K_r1_20, u1_uk_K_r1_23, u1_uk_K_r1_24, u1_uk_K_r1_25, u1_uk_K_r1_26, u1_uk_K_r1_27, u1_uk_K_r1_28, 
       u1_uk_K_r1_29, u1_uk_K_r1_3, u1_uk_K_r1_30, u1_uk_K_r1_31, u1_uk_K_r1_32, u1_uk_K_r1_34, u1_uk_K_r1_35, u1_uk_K_r1_37, u1_uk_K_r1_38, 
       u1_uk_K_r1_39, u1_uk_K_r1_4, u1_uk_K_r1_40, u1_uk_K_r1_43, u1_uk_K_r1_45, u1_uk_K_r1_46, u1_uk_K_r1_48, u1_uk_K_r1_49, u1_uk_K_r1_5, 
       u1_uk_K_r1_50, u1_uk_K_r1_51, u1_uk_K_r1_52, u1_uk_K_r1_53, u1_uk_K_r1_54, u1_uk_K_r1_55, u1_uk_K_r1_8, u1_uk_K_r1_9, u1_uk_K_r2_0, 
       u1_uk_K_r2_1, u1_uk_K_r2_10, u1_uk_K_r2_11, u1_uk_K_r2_12, u1_uk_K_r2_14, u1_uk_K_r2_15, u1_uk_K_r2_17, u1_uk_K_r2_19, u1_uk_K_r2_2, 
       u1_uk_K_r2_22, u1_uk_K_r2_23, u1_uk_K_r2_3, u1_uk_K_r2_30, u1_uk_K_r2_32, u1_uk_K_r2_34, u1_uk_K_r2_35, u1_uk_K_r2_37, u1_uk_K_r2_38, 
       u1_uk_K_r2_39, u1_uk_K_r2_40, u1_uk_K_r2_42, u1_uk_K_r2_43, u1_uk_K_r2_44, u1_uk_K_r2_45, u1_uk_K_r2_48, u1_uk_K_r2_5, u1_uk_K_r2_51, 
       u1_uk_K_r2_52, u1_uk_K_r2_54, u1_uk_K_r2_8, u1_uk_K_r2_9, u1_uk_K_r3_0, u1_uk_K_r3_1, u1_uk_K_r3_12, u1_uk_K_r3_13, u1_uk_K_r3_17, 
       u1_uk_K_r3_18, u1_uk_K_r3_2, u1_uk_K_r3_20, u1_uk_K_r3_21, u1_uk_K_r3_22, u1_uk_K_r3_23, u1_uk_K_r3_25, u1_uk_K_r3_26, u1_uk_K_r3_27, 
       u1_uk_K_r3_28, u1_uk_K_r3_3, u1_uk_K_r3_30, u1_uk_K_r3_31, u1_uk_K_r3_32, u1_uk_K_r3_36, u1_uk_K_r3_37, u1_uk_K_r3_39, u1_uk_K_r3_40, 
       u1_uk_K_r3_41, u1_uk_K_r3_42, u1_uk_K_r3_45, u1_uk_K_r3_46, u1_uk_K_r3_48, u1_uk_K_r3_49, u1_uk_K_r3_5, u1_uk_K_r3_50, u1_uk_K_r3_53, 
       u1_uk_K_r3_54, u1_uk_K_r3_55, u1_uk_K_r3_6, u1_uk_K_r3_7, u1_uk_K_r3_8, u1_uk_K_r4_1, u1_uk_K_r4_10, u1_uk_K_r4_12, u1_uk_K_r4_13, 
       u1_uk_K_r4_14, u1_uk_K_r4_15, u1_uk_K_r4_16, u1_uk_K_r4_19, u1_uk_K_r4_2, u1_uk_K_r4_20, u1_uk_K_r4_21, u1_uk_K_r4_22, u1_uk_K_r4_24, 
       u1_uk_K_r4_25, u1_uk_K_r4_26, u1_uk_K_r4_28, u1_uk_K_r4_29, u1_uk_K_r4_30, u1_uk_K_r4_32, u1_uk_K_r4_34, u1_uk_K_r4_36, u1_uk_K_r4_37, 
       u1_uk_K_r4_39, u1_uk_K_r4_40, u1_uk_K_r4_42, u1_uk_K_r4_43, u1_uk_K_r4_44, u1_uk_K_r4_45, u1_uk_K_r4_46, u1_uk_K_r4_50, u1_uk_K_r4_51, 
       u1_uk_K_r4_52, u1_uk_K_r4_53, u1_uk_K_r4_6, u1_uk_K_r4_7, u1_uk_K_r4_8, u1_uk_K_r4_9, u1_uk_K_r5_11, u1_uk_K_r5_12, u1_uk_K_r5_14, 
       u1_uk_K_r5_15, u1_uk_K_r5_2, u1_uk_K_r5_20, u1_uk_K_r5_22, u1_uk_K_r5_24, u1_uk_K_r5_25, u1_uk_K_r5_27, u1_uk_K_r5_28, u1_uk_K_r5_29, 
       u1_uk_K_r5_3, u1_uk_K_r5_30, u1_uk_K_r5_33, u1_uk_K_r5_34, u1_uk_K_r5_38, u1_uk_K_r5_42, u1_uk_K_r5_44, u1_uk_K_r5_45, u1_uk_K_r5_46, 
       u1_uk_K_r5_47, u1_uk_K_r5_49, u1_uk_K_r5_50, u1_uk_K_r5_52, u1_uk_K_r5_54, u1_uk_K_r5_55, u1_uk_K_r5_6, u1_uk_K_r5_9, u1_uk_K_r6_1, 
       u1_uk_K_r6_11, u1_uk_K_r6_12, u1_uk_K_r6_13, u1_uk_K_r6_15, u1_uk_K_r6_16, u1_uk_K_r6_18, u1_uk_K_r6_2, u1_uk_K_r6_20, u1_uk_K_r6_23, 
       u1_uk_K_r6_24, u1_uk_K_r6_25, u1_uk_K_r6_32, u1_uk_K_r6_33, u1_uk_K_r6_36, u1_uk_K_r6_38, u1_uk_K_r6_39, u1_uk_K_r6_4, u1_uk_K_r6_40, 
       u1_uk_K_r6_41, u1_uk_K_r6_42, u1_uk_K_r6_43, u1_uk_K_r6_44, u1_uk_K_r6_45, u1_uk_K_r6_47, u1_uk_K_r6_48, u1_uk_K_r6_49, u1_uk_K_r6_5, 
       u1_uk_K_r6_50, u1_uk_K_r6_52, u1_uk_K_r6_54, u1_uk_K_r6_6, u1_uk_K_r6_8, u1_uk_K_r6_9, u1_uk_K_r7_10, u1_uk_K_r7_11, u1_uk_K_r7_12, 
       u1_uk_K_r7_14, u1_uk_K_r7_17, u1_uk_K_r7_18, u1_uk_K_r7_19, u1_uk_K_r7_21, u1_uk_K_r7_28, u1_uk_K_r7_3, u1_uk_K_r7_33, u1_uk_K_r7_35, 
       u1_uk_K_r7_36, u1_uk_K_r7_38, u1_uk_K_r7_4, u1_uk_K_r7_40, u1_uk_K_r7_42, u1_uk_K_r7_43, u1_uk_K_r7_44, u1_uk_K_r7_45, u1_uk_K_r7_47, 
       u1_uk_K_r7_49, u1_uk_K_r7_50, u1_uk_K_r7_51, u1_uk_K_r7_52, u1_uk_K_r7_54, u1_uk_K_r8_0, u1_uk_K_r8_1, u1_uk_K_r8_11, u1_uk_K_r8_12, 
       u1_uk_K_r8_14, u1_uk_K_r8_15, u1_uk_K_r8_18, u1_uk_K_r8_20, u1_uk_K_r8_23, u1_uk_K_r8_24, u1_uk_K_r8_25, u1_uk_K_r8_26, u1_uk_K_r8_29, 
       u1_uk_K_r8_3, u1_uk_K_r8_30, u1_uk_K_r8_31, u1_uk_K_r8_33, u1_uk_K_r8_34, u1_uk_K_r8_35, u1_uk_K_r8_36, u1_uk_K_r8_38, u1_uk_K_r8_4, 
       u1_uk_K_r8_45, u1_uk_K_r8_46, u1_uk_K_r8_47, u1_uk_K_r8_49, u1_uk_K_r8_50, u1_uk_K_r8_53, u1_uk_K_r8_54, u1_uk_K_r8_55, u1_uk_K_r8_6, 
       u1_uk_K_r8_7, u1_uk_K_r8_9, u1_uk_K_r9_11, u1_uk_K_r9_14, u1_uk_K_r9_16, u1_uk_K_r9_17, u1_uk_K_r9_2, u1_uk_K_r9_20, u1_uk_K_r9_21, 
       u1_uk_K_r9_24, u1_uk_K_r9_26, u1_uk_K_r9_28, u1_uk_K_r9_29, u1_uk_K_r9_3, u1_uk_K_r9_32, u1_uk_K_r9_34, u1_uk_K_r9_36, u1_uk_K_r9_37, 
       u1_uk_K_r9_39, u1_uk_K_r9_40, u1_uk_K_r9_41, u1_uk_K_r9_42, u1_uk_K_r9_43, u1_uk_K_r9_44, u1_uk_K_r9_46, u1_uk_K_r9_47, u1_uk_K_r9_50, 
       u1_uk_K_r9_51, u1_uk_K_r9_52, u1_uk_K_r9_53, u1_uk_K_r9_8, u2_key_r_15, u2_key_r_18, u2_key_r_38, u2_key_r_39, u2_key_r_45, 
       u2_key_r_5, u2_uk_K_r0_0, u2_uk_K_r0_1, u2_uk_K_r0_10, u2_uk_K_r0_12, u2_uk_K_r0_14, u2_uk_K_r0_16, u2_uk_K_r0_18, u2_uk_K_r0_19, 
       u2_uk_K_r0_2, u2_uk_K_r0_20, u2_uk_K_r0_21, u2_uk_K_r0_22, u2_uk_K_r0_23, u2_uk_K_r0_24, u2_uk_K_r0_26, u2_uk_K_r0_27, u2_uk_K_r0_28, 
       u2_uk_K_r0_29, u2_uk_K_r0_3, u2_uk_K_r0_30, u2_uk_K_r0_33, u2_uk_K_r0_35, u2_uk_K_r0_37, u2_uk_K_r0_38, u2_uk_K_r0_39, u2_uk_K_r0_4, 
       u2_uk_K_r0_40, u2_uk_K_r0_41, u2_uk_K_r0_42, u2_uk_K_r0_43, u2_uk_K_r0_44, u2_uk_K_r0_45, u2_uk_K_r0_46, u2_uk_K_r0_48, u2_uk_K_r0_5, 
       u2_uk_K_r0_50, u2_uk_K_r0_51, u2_uk_K_r0_52, u2_uk_K_r0_53, u2_uk_K_r0_54, u2_uk_K_r0_6, u2_uk_K_r0_7, u2_uk_K_r0_8, u2_uk_K_r0_9, 
       u2_uk_K_r10_0, u2_uk_K_r10_1, u2_uk_K_r10_11, u2_uk_K_r10_12, u2_uk_K_r10_13, u2_uk_K_r10_14, u2_uk_K_r10_15, u2_uk_K_r10_17, u2_uk_K_r10_18, 
       u2_uk_K_r10_19, u2_uk_K_r10_2, u2_uk_K_r10_20, u2_uk_K_r10_21, u2_uk_K_r10_22, u2_uk_K_r10_23, u2_uk_K_r10_24, u2_uk_K_r10_26, u2_uk_K_r10_28, 
       u2_uk_K_r10_29, u2_uk_K_r10_3, u2_uk_K_r10_30, u2_uk_K_r10_31, u2_uk_K_r10_33, u2_uk_K_r10_35, u2_uk_K_r10_36, u2_uk_K_r10_37, u2_uk_K_r10_38, 
       u2_uk_K_r10_39, u2_uk_K_r10_40, u2_uk_K_r10_42, u2_uk_K_r10_45, u2_uk_K_r10_46, u2_uk_K_r10_47, u2_uk_K_r10_48, u2_uk_K_r10_5, u2_uk_K_r10_50, 
       u2_uk_K_r10_51, u2_uk_K_r10_52, u2_uk_K_r10_53, u2_uk_K_r10_54, u2_uk_K_r10_55, u2_uk_K_r10_6, u2_uk_K_r10_7, u2_uk_K_r10_8, u2_uk_K_r10_9, 
       u2_uk_K_r11_0, u2_uk_K_r11_1, u2_uk_K_r11_12, u2_uk_K_r11_13, u2_uk_K_r11_14, u2_uk_K_r11_15, u2_uk_K_r11_16, u2_uk_K_r11_17, u2_uk_K_r11_18, 
       u2_uk_K_r11_2, u2_uk_K_r11_22, u2_uk_K_r11_23, u2_uk_K_r11_3, u2_uk_K_r11_30, u2_uk_K_r11_31, u2_uk_K_r11_32, u2_uk_K_r11_34, u2_uk_K_r11_35, 
       u2_uk_K_r11_36, u2_uk_K_r11_37, u2_uk_K_r11_38, u2_uk_K_r11_40, u2_uk_K_r11_41, u2_uk_K_r11_42, u2_uk_K_r11_43, u2_uk_K_r11_44, u2_uk_K_r11_45, 
       u2_uk_K_r11_46, u2_uk_K_r11_49, u2_uk_K_r11_5, u2_uk_K_r11_50, u2_uk_K_r11_51, u2_uk_K_r11_52, u2_uk_K_r11_54, u2_uk_K_r11_55, u2_uk_K_r11_8, 
       u2_uk_K_r11_9, u2_uk_K_r12_0, u2_uk_K_r12_11, u2_uk_K_r12_12, u2_uk_K_r12_13, u2_uk_K_r12_14, u2_uk_K_r12_17, u2_uk_K_r12_18, u2_uk_K_r12_19, 
       u2_uk_K_r12_2, u2_uk_K_r12_20, u2_uk_K_r12_21, u2_uk_K_r12_22, u2_uk_K_r12_23, u2_uk_K_r12_24, u2_uk_K_r12_26, u2_uk_K_r12_27, u2_uk_K_r12_28, 
       u2_uk_K_r12_29, u2_uk_K_r12_3, u2_uk_K_r12_31, u2_uk_K_r12_32, u2_uk_K_r12_34, u2_uk_K_r12_35, u2_uk_K_r12_37, u2_uk_K_r12_38, u2_uk_K_r12_39, 
       u2_uk_K_r12_4, u2_uk_K_r12_40, u2_uk_K_r12_43, u2_uk_K_r12_44, u2_uk_K_r12_45, u2_uk_K_r12_46, u2_uk_K_r12_47, u2_uk_K_r12_48, u2_uk_K_r12_49, 
       u2_uk_K_r12_5, u2_uk_K_r12_50, u2_uk_K_r12_51, u2_uk_K_r12_52, u2_uk_K_r12_53, u2_uk_K_r12_54, u2_uk_K_r12_55, u2_uk_K_r12_6, u2_uk_K_r12_8, 
       u2_uk_K_r12_9, u2_uk_K_r13_1, u2_uk_K_r13_10, u2_uk_K_r13_11, u2_uk_K_r13_12, u2_uk_K_r13_14, u2_uk_K_r13_15, u2_uk_K_r13_16, u2_uk_K_r13_18, 
       u2_uk_K_r13_2, u2_uk_K_r13_20, u2_uk_K_r13_21, u2_uk_K_r13_23, u2_uk_K_r13_24, u2_uk_K_r13_26, u2_uk_K_r13_27, u2_uk_K_r13_28, u2_uk_K_r13_29, 
       u2_uk_K_r13_3, u2_uk_K_r13_30, u2_uk_K_r13_31, u2_uk_K_r13_33, u2_uk_K_r13_34, u2_uk_K_r13_35, u2_uk_K_r13_36, u2_uk_K_r13_37, u2_uk_K_r13_39, 
       u2_uk_K_r13_4, u2_uk_K_r13_40, u2_uk_K_r13_41, u2_uk_K_r13_42, u2_uk_K_r13_43, u2_uk_K_r13_44, u2_uk_K_r13_45, u2_uk_K_r13_46, u2_uk_K_r13_47, 
       u2_uk_K_r13_48, u2_uk_K_r13_49, u2_uk_K_r13_5, u2_uk_K_r13_50, u2_uk_K_r13_51, u2_uk_K_r13_52, u2_uk_K_r13_53, u2_uk_K_r13_54, u2_uk_K_r13_6, 
       u2_uk_K_r13_7, u2_uk_K_r13_8, u2_uk_K_r13_9, u2_uk_K_r14_11, u2_uk_K_r14_23, u2_uk_K_r14_38, u2_uk_K_r14_39, u2_uk_K_r14_42, u2_uk_K_r14_43, 
       u2_uk_K_r14_8, u2_uk_K_r1_0, u2_uk_K_r1_1, u2_uk_K_r1_10, u2_uk_K_r1_11, u2_uk_K_r1_12, u2_uk_K_r1_13, u2_uk_K_r1_14, u2_uk_K_r1_19, 
       u2_uk_K_r1_2, u2_uk_K_r1_20, u2_uk_K_r1_23, u2_uk_K_r1_24, u2_uk_K_r1_25, u2_uk_K_r1_26, u2_uk_K_r1_27, u2_uk_K_r1_28, u2_uk_K_r1_29, 
       u2_uk_K_r1_3, u2_uk_K_r1_30, u2_uk_K_r1_31, u2_uk_K_r1_32, u2_uk_K_r1_33, u2_uk_K_r1_34, u2_uk_K_r1_35, u2_uk_K_r1_36, u2_uk_K_r1_37, 
       u2_uk_K_r1_38, u2_uk_K_r1_39, u2_uk_K_r1_4, u2_uk_K_r1_40, u2_uk_K_r1_43, u2_uk_K_r1_45, u2_uk_K_r1_46, u2_uk_K_r1_48, u2_uk_K_r1_49, 
       u2_uk_K_r1_5, u2_uk_K_r1_50, u2_uk_K_r1_51, u2_uk_K_r1_52, u2_uk_K_r1_53, u2_uk_K_r1_54, u2_uk_K_r1_55, u2_uk_K_r1_6, u2_uk_K_r1_8, 
       u2_uk_K_r1_9, u2_uk_K_r2_0, u2_uk_K_r2_1, u2_uk_K_r2_10, u2_uk_K_r2_11, u2_uk_K_r2_12, u2_uk_K_r2_14, u2_uk_K_r2_15, u2_uk_K_r2_16, 
       u2_uk_K_r2_17, u2_uk_K_r2_19, u2_uk_K_r2_2, u2_uk_K_r2_20, u2_uk_K_r2_22, u2_uk_K_r2_23, u2_uk_K_r2_29, u2_uk_K_r2_3, u2_uk_K_r2_30, 
       u2_uk_K_r2_32, u2_uk_K_r2_33, u2_uk_K_r2_34, u2_uk_K_r2_35, u2_uk_K_r2_37, u2_uk_K_r2_38, u2_uk_K_r2_39, u2_uk_K_r2_4, u2_uk_K_r2_40, 
       u2_uk_K_r2_41, u2_uk_K_r2_42, u2_uk_K_r2_43, u2_uk_K_r2_44, u2_uk_K_r2_45, u2_uk_K_r2_46, u2_uk_K_r2_47, u2_uk_K_r2_48, u2_uk_K_r2_5, 
       u2_uk_K_r2_51, u2_uk_K_r2_52, u2_uk_K_r2_53, u2_uk_K_r2_54, u2_uk_K_r2_7, u2_uk_K_r2_8, u2_uk_K_r2_9, u2_uk_K_r3_0, u2_uk_K_r3_1, 
       u2_uk_K_r3_12, u2_uk_K_r3_13, u2_uk_K_r3_17, u2_uk_K_r3_18, u2_uk_K_r3_2, u2_uk_K_r3_20, u2_uk_K_r3_21, u2_uk_K_r3_22, u2_uk_K_r3_23, 
       u2_uk_K_r3_24, u2_uk_K_r3_25, u2_uk_K_r3_26, u2_uk_K_r3_27, u2_uk_K_r3_28, u2_uk_K_r3_3, u2_uk_K_r3_30, u2_uk_K_r3_31, u2_uk_K_r3_32, 
       u2_uk_K_r3_33, u2_uk_K_r3_34, u2_uk_K_r3_35, u2_uk_K_r3_36, u2_uk_K_r3_37, u2_uk_K_r3_39, u2_uk_K_r3_40, u2_uk_K_r3_41, u2_uk_K_r3_42, 
       u2_uk_K_r3_44, u2_uk_K_r3_45, u2_uk_K_r3_46, u2_uk_K_r3_47, u2_uk_K_r3_48, u2_uk_K_r3_49, u2_uk_K_r3_5, u2_uk_K_r3_50, u2_uk_K_r3_51, 
       u2_uk_K_r3_53, u2_uk_K_r3_54, u2_uk_K_r3_55, u2_uk_K_r3_6, u2_uk_K_r3_7, u2_uk_K_r3_8, u2_uk_K_r4_1, u2_uk_K_r4_10, u2_uk_K_r4_12, 
       u2_uk_K_r4_13, u2_uk_K_r4_14, u2_uk_K_r4_15, u2_uk_K_r4_16, u2_uk_K_r4_18, u2_uk_K_r4_19, u2_uk_K_r4_2, u2_uk_K_r4_20, u2_uk_K_r4_21, 
       u2_uk_K_r4_22, u2_uk_K_r4_23, u2_uk_K_r4_24, u2_uk_K_r4_25, u2_uk_K_r4_26, u2_uk_K_r4_27, u2_uk_K_r4_28, u2_uk_K_r4_29, u2_uk_K_r4_30, 
       u2_uk_K_r4_31, u2_uk_K_r4_32, u2_uk_K_r4_34, u2_uk_K_r4_36, u2_uk_K_r4_37, u2_uk_K_r4_39, u2_uk_K_r4_40, u2_uk_K_r4_42, u2_uk_K_r4_43, 
       u2_uk_K_r4_44, u2_uk_K_r4_45, u2_uk_K_r4_46, u2_uk_K_r4_48, u2_uk_K_r4_49, u2_uk_K_r4_50, u2_uk_K_r4_51, u2_uk_K_r4_52, u2_uk_K_r4_53, 
       u2_uk_K_r4_6, u2_uk_K_r4_7, u2_uk_K_r4_8, u2_uk_K_r4_9, u2_uk_K_r5_11, u2_uk_K_r5_12, u2_uk_K_r5_13, u2_uk_K_r5_14, u2_uk_K_r5_15, 
       u2_uk_K_r5_2, u2_uk_K_r5_20, u2_uk_K_r5_22, u2_uk_K_r5_24, u2_uk_K_r5_25, u2_uk_K_r5_27, u2_uk_K_r5_28, u2_uk_K_r5_29, u2_uk_K_r5_3, 
       u2_uk_K_r5_30, u2_uk_K_r5_32, u2_uk_K_r5_33, u2_uk_K_r5_34, u2_uk_K_r5_35, u2_uk_K_r5_36, u2_uk_K_r5_38, u2_uk_K_r5_42, u2_uk_K_r5_44, 
       u2_uk_K_r5_45, u2_uk_K_r5_46, u2_uk_K_r5_47, u2_uk_K_r5_49, u2_uk_K_r5_5, u2_uk_K_r5_50, u2_uk_K_r5_52, u2_uk_K_r5_53, u2_uk_K_r5_54, 
       u2_uk_K_r5_55, u2_uk_K_r5_6, u2_uk_K_r5_8, u2_uk_K_r5_9, u2_uk_K_r6_1, u2_uk_K_r6_11, u2_uk_K_r6_12, u2_uk_K_r6_13, u2_uk_K_r6_15, 
       u2_uk_K_r6_16, u2_uk_K_r6_17, u2_uk_K_r6_18, u2_uk_K_r6_19, u2_uk_K_r6_2, u2_uk_K_r6_20, u2_uk_K_r6_21, u2_uk_K_r6_22, u2_uk_K_r6_23, 
       u2_uk_K_r6_24, u2_uk_K_r6_25, u2_uk_K_r6_27, u2_uk_K_r6_28, u2_uk_K_r6_30, u2_uk_K_r6_32, u2_uk_K_r6_33, u2_uk_K_r6_35, u2_uk_K_r6_36, 
       u2_uk_K_r6_38, u2_uk_K_r6_39, u2_uk_K_r6_4, u2_uk_K_r6_40, u2_uk_K_r6_41, u2_uk_K_r6_42, u2_uk_K_r6_43, u2_uk_K_r6_44, u2_uk_K_r6_45, 
       u2_uk_K_r6_47, u2_uk_K_r6_48, u2_uk_K_r6_49, u2_uk_K_r6_5, u2_uk_K_r6_50, u2_uk_K_r6_52, u2_uk_K_r6_54, u2_uk_K_r6_55, u2_uk_K_r6_6, 
       u2_uk_K_r6_8, u2_uk_K_r6_9, u2_uk_K_r7_1, u2_uk_K_r7_10, u2_uk_K_r7_11, u2_uk_K_r7_12, u2_uk_K_r7_14, u2_uk_K_r7_15, u2_uk_K_r7_17, 
       u2_uk_K_r7_18, u2_uk_K_r7_19, u2_uk_K_r7_21, u2_uk_K_r7_22, u2_uk_K_r7_24, u2_uk_K_r7_27, u2_uk_K_r7_28, u2_uk_K_r7_29, u2_uk_K_r7_3, 
       u2_uk_K_r7_30, u2_uk_K_r7_33, u2_uk_K_r7_34, u2_uk_K_r7_35, u2_uk_K_r7_36, u2_uk_K_r7_38, u2_uk_K_r7_4, u2_uk_K_r7_40, u2_uk_K_r7_42, 
       u2_uk_K_r7_43, u2_uk_K_r7_44, u2_uk_K_r7_45, u2_uk_K_r7_47, u2_uk_K_r7_49, u2_uk_K_r7_5, u2_uk_K_r7_50, u2_uk_K_r7_51, u2_uk_K_r7_52, 
       u2_uk_K_r7_53, u2_uk_K_r7_54, u2_uk_K_r7_6, u2_uk_K_r7_7, u2_uk_K_r7_8, u2_uk_K_r8_0, u2_uk_K_r8_1, u2_uk_K_r8_10, u2_uk_K_r8_11, 
       u2_uk_K_r8_12, u2_uk_K_r8_14, u2_uk_K_r8_15, u2_uk_K_r8_18, u2_uk_K_r8_20, u2_uk_K_r8_23, u2_uk_K_r8_24, u2_uk_K_r8_25, u2_uk_K_r8_26, 
       u2_uk_K_r8_29, u2_uk_K_r8_3, u2_uk_K_r8_30, u2_uk_K_r8_31, u2_uk_K_r8_33, u2_uk_K_r8_34, u2_uk_K_r8_35, u2_uk_K_r8_36, u2_uk_K_r8_38, 
       u2_uk_K_r8_39, u2_uk_K_r8_4, u2_uk_K_r8_45, u2_uk_K_r8_46, u2_uk_K_r8_47, u2_uk_K_r8_49, u2_uk_K_r8_5, u2_uk_K_r8_50, u2_uk_K_r8_51, 
       u2_uk_K_r8_53, u2_uk_K_r8_54, u2_uk_K_r8_55, u2_uk_K_r8_6, u2_uk_K_r8_7, u2_uk_K_r8_9, u2_uk_K_r9_11, u2_uk_K_r9_14, u2_uk_K_r9_16, 
       u2_uk_K_r9_17, u2_uk_K_r9_2, u2_uk_K_r9_20, u2_uk_K_r9_21, u2_uk_K_r9_22, u2_uk_K_r9_24, u2_uk_K_r9_26, u2_uk_K_r9_28, u2_uk_K_r9_29, 
       u2_uk_K_r9_3, u2_uk_K_r9_30, u2_uk_K_r9_32, u2_uk_K_r9_34, u2_uk_K_r9_35, u2_uk_K_r9_36, u2_uk_K_r9_37, u2_uk_K_r9_38, u2_uk_K_r9_39, 
       u2_uk_K_r9_40, u2_uk_K_r9_41, u2_uk_K_r9_42, u2_uk_K_r9_43, u2_uk_K_r9_44, u2_uk_K_r9_46, u2_uk_K_r9_47, u2_uk_K_r9_50, u2_uk_K_r9_51, 
       u2_uk_K_r9_52, u2_uk_K_r9_53, u2_uk_K_r9_6, u2_uk_K_r9_7, u2_uk_K_r9_8, u2_uk_n1002, u2_uk_n1003, u2_uk_n1006, u2_uk_n1025, 
       u2_uk_n1045, u2_uk_n1047, u2_uk_n1067, u2_uk_n1092, u2_uk_n1111, u2_uk_n1191, u2_uk_n1192, u2_uk_n1211, u2_uk_n1235, 
       u2_uk_n1241, u2_uk_n1242, u2_uk_n1256, u2_uk_n1262, u2_uk_n1263, u2_uk_n1273, u2_uk_n1277, u2_uk_n1278, u2_uk_n1289, 
       u2_uk_n1304, u2_uk_n1327, u2_uk_n1366, u2_uk_n1368, u2_uk_n1369, u2_uk_n1371, u2_uk_n1373, u2_uk_n1374, u2_uk_n1380, 
       u2_uk_n1384, u2_uk_n1385, u2_uk_n1387, u2_uk_n1388, u2_uk_n1389, u2_uk_n1392, u2_uk_n1393, u2_uk_n1394, u2_uk_n1397, 
       u2_uk_n1399, u2_uk_n1406, u2_uk_n1407, u2_uk_n1409, u2_uk_n1417, u2_uk_n1423, u2_uk_n1427, u2_uk_n1431, u2_uk_n1432, 
       u2_uk_n1434, u2_uk_n1436, u2_uk_n1455, u2_uk_n1469, u2_uk_n1474, u2_uk_n1477, u2_uk_n1478, u2_uk_n1484, u2_uk_n1534, 
       u2_uk_n1540, u2_uk_n1541, u2_uk_n1547, u2_uk_n1554, u2_uk_n1562, u2_uk_n1569, u2_uk_n1575, u2_uk_n1578, u2_uk_n1582, 
       u2_uk_n1584, u2_uk_n1588, u2_uk_n1589, u2_uk_n1593, u2_uk_n1596, u2_uk_n1611, u2_uk_n1619, u2_uk_n1621, u2_uk_n1637, 
       u2_uk_n1648, u2_uk_n1662, u2_uk_n1663, u2_uk_n1669, u2_uk_n1679, u2_uk_n1686, u2_uk_n1692, u2_uk_n1701, u2_uk_n1704, 
       u2_uk_n1706, u2_uk_n1714, u2_uk_n1719, u2_uk_n1733, u2_uk_n1739, u2_uk_n1751, u2_uk_n1752, u2_uk_n1754, u2_uk_n1757, 
       u2_uk_n1771, u2_uk_n1774, u2_uk_n1780, u2_uk_n1784, u2_uk_n1787, u2_uk_n1804, u2_uk_n1812, u2_uk_n1813, u2_uk_n1829, 
       u2_uk_n1830, u2_uk_n1844, u2_uk_n1857, u2_uk_n292, u2_uk_n437, u2_uk_n695, u2_uk_n962,  u2_uk_n964;
  OAI22_X1 U172 (.B1( decrypt ) , .ZN( key_a_0 ) , .A2( n112 ) , .A1( n115 ) , .B2( n56 ) );
  INV_X1 U173 (.A( key1[0] ) , .ZN( n56 ) );
  INV_X1 U174 (.A( key3[0] ) , .ZN( n112 ) );
  OAI22_X1 U175 (.B1( decrypt ) , .ZN( key_a_10 ) , .A2( n102 ) , .A1( n114 ) , .B2( n46 ) );
  INV_X1 U176 (.A( key1[10] ) , .ZN( n46 ) );
  INV_X1 U177 (.A( key3[10] ) , .ZN( n102 ) );
  OAI22_X1 U178 (.B1( decrypt ) , .ZN( key_a_11 ) , .A2( n101 ) , .A1( n116 ) , .B2( n45 ) );
  INV_X1 U179 (.A( key1[11] ) , .ZN( n45 ) );
  INV_X1 U180 (.A( key3[11] ) , .ZN( n101 ) );
  OAI22_X1 U181 (.B1( decrypt ) , .ZN( key_a_12 ) , .A2( n100 ) , .A1( n116 ) , .B2( n44 ) );
  INV_X1 U182 (.A( key1[12] ) , .ZN( n44 ) );
  INV_X1 U183 (.A( key3[12] ) , .ZN( n100 ) );
  OAI22_X1 U184 (.B1( decrypt ) , .ZN( key_a_13 ) , .A1( n116 ) , .B2( n43 ) , .A2( n99 ) );
  INV_X1 U185 (.A( key1[13] ) , .ZN( n43 ) );
  INV_X1 U186 (.A( key3[13] ) , .ZN( n99 ) );
  OAI22_X1 U187 (.B1( decrypt ) , .ZN( key_a_14 ) , .A1( n116 ) , .B2( n42 ) , .A2( n98 ) );
  INV_X1 U188 (.A( key1[14] ) , .ZN( n42 ) );
  INV_X1 U189 (.A( key3[14] ) , .ZN( n98 ) );
  OAI22_X1 U190 (.B1( decrypt ) , .ZN( key_a_1 ) , .A2( n111 ) , .A1( n116 ) , .B2( n55 ) );
  INV_X1 U191 (.A( key1[1] ) , .ZN( n55 ) );
  INV_X1 U192 (.A( key3[1] ) , .ZN( n111 ) );
  OAI22_X1 U193 (.B1( decrypt ) , .ZN( key_a_2 ) , .A2( n110 ) , .A1( n115 ) , .B2( n54 ) );
  INV_X1 U194 (.A( key1[2] ) , .ZN( n54 ) );
  INV_X1 U195 (.A( key3[2] ) , .ZN( n110 ) );
  OAI22_X1 U196 (.B1( decrypt ) , .ZN( key_a_3 ) , .A2( n109 ) , .A1( n114 ) , .B2( n53 ) );
  INV_X1 U197 (.A( key1[3] ) , .ZN( n53 ) );
  INV_X1 U198 (.A( key3[3] ) , .ZN( n109 ) );
  OAI22_X1 U199 (.B1( decrypt ) , .ZN( key_a_4 ) , .A2( n108 ) , .A1( n114 ) , .B2( n52 ) );
  INV_X1 U200 (.A( key1[4] ) , .ZN( n52 ) );
  INV_X1 U201 (.A( key3[4] ) , .ZN( n108 ) );
  OAI22_X1 U202 (.B1( decrypt ) , .ZN( key_a_9 ) , .A2( n103 ) , .A1( n115 ) , .B2( n47 ) );
  INV_X1 U203 (.A( key1[9] ) , .ZN( n47 ) );
  INV_X1 U204 (.A( key3[9] ) , .ZN( n103 ) );
  OAI22_X1 U205 (.B1( decrypt ) , .ZN( key_a_15 ) , .A1( n116 ) , .B2( n41 ) , .A2( n97 ) );
  INV_X1 U206 (.A( key1[15] ) , .ZN( n41 ) );
  INV_X1 U207 (.A( key3[15] ) , .ZN( n97 ) );
  OAI22_X1 U208 (.B1( decrypt ) , .ZN( key_a_16 ) , .A1( n116 ) , .B2( n40 ) , .A2( n96 ) );
  INV_X1 U209 (.A( key1[16] ) , .ZN( n40 ) );
  INV_X1 U210 (.A( key3[16] ) , .ZN( n96 ) );
  OAI22_X1 U211 (.B1( decrypt ) , .ZN( key_a_17 ) , .A1( n116 ) , .B2( n39 ) , .A2( n95 ) );
  INV_X1 U212 (.A( key1[17] ) , .ZN( n39 ) );
  INV_X1 U213 (.A( key3[17] ) , .ZN( n95 ) );
  OAI22_X1 U214 (.B1( decrypt ) , .ZN( key_a_18 ) , .A1( n116 ) , .B2( n38 ) , .A2( n94 ) );
  INV_X1 U215 (.A( key1[18] ) , .ZN( n38 ) );
  INV_X1 U216 (.A( key3[18] ) , .ZN( n94 ) );
  OAI22_X1 U217 (.B1( decrypt ) , .ZN( key_a_19 ) , .A1( n116 ) , .B2( n37 ) , .A2( n93 ) );
  INV_X1 U218 (.A( key1[19] ) , .ZN( n37 ) );
  INV_X1 U219 (.A( key3[19] ) , .ZN( n93 ) );
  OAI22_X1 U220 (.B1( decrypt ) , .ZN( key_a_20 ) , .A1( n116 ) , .B2( n36 ) , .A2( n92 ) );
  INV_X1 U221 (.A( key1[20] ) , .ZN( n36 ) );
  INV_X1 U222 (.A( key3[20] ) , .ZN( n92 ) );
  OAI22_X1 U223 (.B1( decrypt ) , .ZN( key_a_21 ) , .A1( n116 ) , .B2( n35 ) , .A2( n91 ) );
  INV_X1 U224 (.A( key1[21] ) , .ZN( n35 ) );
  INV_X1 U225 (.A( key3[21] ) , .ZN( n91 ) );
  OAI22_X1 U226 (.B1( decrypt ) , .ZN( key_a_22 ) , .A1( n116 ) , .B2( n34 ) , .A2( n90 ) );
  INV_X1 U227 (.A( key1[22] ) , .ZN( n34 ) );
  INV_X1 U228 (.A( key3[22] ) , .ZN( n90 ) );
  OAI22_X1 U229 (.B1( decrypt ) , .ZN( key_a_23 ) , .A1( n116 ) , .B2( n33 ) , .A2( n89 ) );
  INV_X1 U230 (.A( key1[23] ) , .ZN( n33 ) );
  INV_X1 U231 (.A( key3[23] ) , .ZN( n89 ) );
  OAI22_X1 U232 (.B1( decrypt ) , .ZN( key_a_24 ) , .A1( n116 ) , .B2( n32 ) , .A2( n88 ) );
  INV_X1 U233 (.A( key1[24] ) , .ZN( n32 ) );
  INV_X1 U234 (.A( key3[24] ) , .ZN( n88 ) );
  OAI22_X1 U235 (.B1( decrypt ) , .ZN( key_a_25 ) , .A1( n116 ) , .B2( n31 ) , .A2( n87 ) );
  INV_X1 U236 (.A( key1[25] ) , .ZN( n31 ) );
  INV_X1 U237 (.A( key3[25] ) , .ZN( n87 ) );
  OAI22_X1 U238 (.B1( decrypt ) , .ZN( key_a_26 ) , .A1( n115 ) , .B2( n30 ) , .A2( n86 ) );
  INV_X1 U239 (.A( key1[26] ) , .ZN( n30 ) );
  INV_X1 U240 (.A( key3[26] ) , .ZN( n86 ) );
  OAI22_X1 U241 (.B1( decrypt ) , .ZN( key_a_27 ) , .A1( n115 ) , .B2( n29 ) , .A2( n85 ) );
  INV_X1 U242 (.A( key1[27] ) , .ZN( n29 ) );
  INV_X1 U243 (.A( key3[27] ) , .ZN( n85 ) );
  OAI22_X1 U244 (.B1( decrypt ) , .ZN( key_a_28 ) , .A1( n115 ) , .B2( n28 ) , .A2( n84 ) );
  INV_X1 U245 (.A( key1[28] ) , .ZN( n28 ) );
  INV_X1 U246 (.A( key3[28] ) , .ZN( n84 ) );
  OAI22_X1 U247 (.B1( decrypt ) , .ZN( key_a_29 ) , .A1( n115 ) , .B2( n27 ) , .A2( n83 ) );
  INV_X1 U248 (.A( key1[29] ) , .ZN( n27 ) );
  INV_X1 U249 (.A( key3[29] ) , .ZN( n83 ) );
  OAI22_X1 U250 (.B1( decrypt ) , .ZN( key_a_30 ) , .A1( n115 ) , .B2( n26 ) , .A2( n82 ) );
  INV_X1 U251 (.A( key1[30] ) , .ZN( n26 ) );
  INV_X1 U252 (.A( key3[30] ) , .ZN( n82 ) );
  OAI22_X1 U253 (.B1( decrypt ) , .ZN( key_a_31 ) , .A1( n115 ) , .B2( n25 ) , .A2( n81 ) );
  INV_X1 U254 (.A( key1[31] ) , .ZN( n25 ) );
  INV_X1 U255 (.A( key3[31] ) , .ZN( n81 ) );
  OAI22_X1 U256 (.B1( decrypt ) , .ZN( key_a_32 ) , .A1( n115 ) , .B2( n24 ) , .A2( n80 ) );
  INV_X1 U257 (.A( key1[32] ) , .ZN( n24 ) );
  INV_X1 U258 (.A( key3[32] ) , .ZN( n80 ) );
  OAI22_X1 U259 (.B1( decrypt ) , .ZN( key_a_33 ) , .A1( n115 ) , .B2( n23 ) , .A2( n79 ) );
  INV_X1 U260 (.A( key1[33] ) , .ZN( n23 ) );
  INV_X1 U261 (.A( key3[33] ) , .ZN( n79 ) );
  OAI22_X1 U262 (.B1( decrypt ) , .ZN( key_a_34 ) , .A1( n115 ) , .B2( n22 ) , .A2( n78 ) );
  INV_X1 U263 (.A( key1[34] ) , .ZN( n22 ) );
  INV_X1 U264 (.A( key3[34] ) , .ZN( n78 ) );
  OAI22_X1 U265 (.B1( decrypt ) , .ZN( key_a_35 ) , .A1( n115 ) , .B2( n21 ) , .A2( n77 ) );
  INV_X1 U266 (.A( key1[35] ) , .ZN( n21 ) );
  INV_X1 U267 (.A( key3[35] ) , .ZN( n77 ) );
  OAI22_X1 U268 (.B1( decrypt ) , .ZN( key_a_36 ) , .A1( n115 ) , .B2( n20 ) , .A2( n76 ) );
  INV_X1 U269 (.A( key1[36] ) , .ZN( n20 ) );
  INV_X1 U270 (.A( key3[36] ) , .ZN( n76 ) );
  OAI22_X1 U271 (.B1( decrypt ) , .ZN( key_a_37 ) , .A1( n115 ) , .B2( n19 ) , .A2( n75 ) );
  INV_X1 U272 (.A( key1[37] ) , .ZN( n19 ) );
  INV_X1 U273 (.A( key3[37] ) , .ZN( n75 ) );
  OAI22_X1 U274 (.B1( decrypt ) , .ZN( key_a_38 ) , .A1( n115 ) , .B2( n18 ) , .A2( n74 ) );
  INV_X1 U275 (.A( key1[38] ) , .ZN( n18 ) );
  INV_X1 U276 (.A( key3[38] ) , .ZN( n74 ) );
  OAI22_X1 U277 (.B1( decrypt ) , .ZN( key_a_39 ) , .A1( n115 ) , .B2( n17 ) , .A2( n73 ) );
  INV_X1 U278 (.A( key1[39] ) , .ZN( n17 ) );
  INV_X1 U279 (.A( key3[39] ) , .ZN( n73 ) );
  OAI22_X1 U280 (.B1( decrypt ) , .ZN( key_a_40 ) , .A1( n114 ) , .B2( n16 ) , .A2( n72 ) );
  INV_X1 U281 (.A( key1[40] ) , .ZN( n16 ) );
  INV_X1 U282 (.A( key3[40] ) , .ZN( n72 ) );
  OAI22_X1 U283 (.B1( decrypt ) , .ZN( key_a_41 ) , .A1( n114 ) , .B2( n15 ) , .A2( n71 ) );
  INV_X1 U284 (.A( key1[41] ) , .ZN( n15 ) );
  INV_X1 U285 (.A( key3[41] ) , .ZN( n71 ) );
  OAI22_X1 U286 (.B1( decrypt ) , .ZN( key_a_42 ) , .A1( n114 ) , .B2( n14 ) , .A2( n70 ) );
  INV_X1 U287 (.A( key1[42] ) , .ZN( n14 ) );
  INV_X1 U288 (.A( key3[42] ) , .ZN( n70 ) );
  OAI22_X1 U289 (.B1( decrypt ) , .ZN( key_a_43 ) , .A1( n114 ) , .B2( n13 ) , .A2( n69 ) );
  INV_X1 U290 (.A( key1[43] ) , .ZN( n13 ) );
  INV_X1 U291 (.A( key3[43] ) , .ZN( n69 ) );
  OAI22_X1 U292 (.B1( decrypt ) , .ZN( key_a_44 ) , .A1( n114 ) , .B2( n12 ) , .A2( n68 ) );
  INV_X1 U293 (.A( key1[44] ) , .ZN( n12 ) );
  INV_X1 U294 (.A( key3[44] ) , .ZN( n68 ) );
  OAI22_X1 U295 (.B1( decrypt ) , .ZN( key_a_45 ) , .B2( n11 ) , .A1( n114 ) , .A2( n67 ) );
  INV_X1 U296 (.A( key1[45] ) , .ZN( n11 ) );
  INV_X1 U297 (.A( key3[45] ) , .ZN( n67 ) );
  OAI22_X1 U298 (.B1( decrypt ) , .ZN( key_a_46 ) , .B2( n10 ) , .A1( n114 ) , .A2( n66 ) );
  INV_X1 U299 (.A( key1[46] ) , .ZN( n10 ) );
  INV_X1 U300 (.A( key3[46] ) , .ZN( n66 ) );
  OAI22_X1 U301 (.B1( decrypt ) , .ZN( key_a_47 ) , .A1( n114 ) , .A2( n65 ) , .B2( n9 ) );
  INV_X1 U302 (.A( key1[47] ) , .ZN( n9 ) );
  INV_X1 U303 (.A( key3[47] ) , .ZN( n65 ) );
  OAI22_X1 U304 (.B1( decrypt ) , .ZN( key_a_48 ) , .A1( n114 ) , .A2( n64 ) , .B2( n8 ) );
  INV_X1 U305 (.A( key1[48] ) , .ZN( n8 ) );
  INV_X1 U306 (.A( key3[48] ) , .ZN( n64 ) );
  OAI22_X1 U307 (.B1( decrypt ) , .ZN( key_a_49 ) , .A1( n114 ) , .A2( n63 ) , .B2( n7 ) );
  INV_X1 U308 (.A( key1[49] ) , .ZN( n7 ) );
  INV_X1 U309 (.A( key3[49] ) , .ZN( n63 ) );
  OAI22_X1 U310 (.B1( decrypt ) , .ZN( key_a_50 ) , .A1( n114 ) , .B2( n6 ) , .A2( n62 ) );
  INV_X1 U311 (.A( key1[50] ) , .ZN( n6 ) );
  INV_X1 U312 (.A( key3[50] ) , .ZN( n62 ) );
  OAI22_X1 U313 (.B1( decrypt ) , .ZN( key_a_51 ) , .A1( n114 ) , .B2( n5 ) , .A2( n61 ) );
  INV_X1 U314 (.A( key1[51] ) , .ZN( n5 ) );
  INV_X1 U315 (.A( key3[51] ) , .ZN( n61 ) );
  OAI22_X1 U316 (.B1( decrypt ) , .ZN( key_a_5 ) , .A2( n107 ) , .A1( n114 ) , .B2( n51 ) );
  INV_X1 U317 (.A( key1[5] ) , .ZN( n51 ) );
  INV_X1 U318 (.A( key3[5] ) , .ZN( n107 ) );
  OAI22_X1 U319 (.B1( decrypt ) , .ZN( key_a_6 ) , .A2( n106 ) , .A1( n114 ) , .B2( n50 ) );
  INV_X1 U320 (.A( key1[6] ) , .ZN( n50 ) );
  INV_X1 U321 (.A( key3[6] ) , .ZN( n106 ) );
  OAI22_X1 U322 (.B1( decrypt ) , .ZN( key_a_7 ) , .A2( n105 ) , .A1( n116 ) , .B2( n49 ) );
  INV_X1 U323 (.A( key1[7] ) , .ZN( n49 ) );
  INV_X1 U324 (.A( key3[7] ) , .ZN( n105 ) );
  OAI22_X1 U325 (.B1( decrypt ) , .ZN( key_a_8 ) , .A2( n104 ) , .A1( n115 ) , .B2( n48 ) );
  INV_X1 U326 (.A( key1[8] ) , .ZN( n48 ) );
  INV_X1 U327 (.A( key3[8] ) , .ZN( n104 ) );
  OAI22_X1 U328 (.B1( decrypt ) , .ZN( key_a_52 ) , .A1( n114 ) , .B2( n4 ) , .A2( n60 ) );
  INV_X1 U329 (.A( key1[52] ) , .ZN( n4 ) );
  INV_X1 U330 (.A( key3[52] ) , .ZN( n60 ) );
  OAI22_X1 U331 (.B1( decrypt ) , .ZN( key_a_53 ) , .A1( n114 ) , .B2( n3 ) , .A2( n59 ) );
  INV_X1 U332 (.A( key1[53] ) , .ZN( n3 ) );
  INV_X1 U333 (.A( key3[53] ) , .ZN( n59 ) );
  OAI22_X1 U334 (.B1( decrypt ) , .ZN( key_a_54 ) , .A1( n114 ) , .B2( n2 ) , .A2( n58 ) );
  INV_X1 U335 (.A( key1[54] ) , .ZN( n2 ) );
  INV_X1 U336 (.A( key3[54] ) , .ZN( n58 ) );
  OAI22_X1 U337 (.B1( decrypt ) , .ZN( key_a_55 ) , .B2( n1 ) , .A1( n116 ) , .A2( n57 ) );
  INV_X1 U338 (.A( key1[55] ) , .ZN( n1 ) );
  INV_X1 U339 (.A( key3[55] ) , .ZN( n57 ) );
  INV_X1 U340 (.A( decrypt ) , .ZN( n116 ) );
  INV_X1 U341 (.A( decrypt ) , .ZN( n115 ) );
  INV_X1 U342 (.A( decrypt ) , .ZN( n114 ) );
  DFF_X1 key_b_r_reg_0_0 (.CK( clk ) , .D( key2[0] ) , .Q( key_b_r_0_0 ) );
  DFF_X1 key_b_r_reg_0_1 (.CK( clk ) , .D( key2[1] ) , .Q( key_b_r_0_1 ) );
  DFF_X1 key_b_r_reg_0_10 (.CK( clk ) , .D( key2[10] ) , .Q( key_b_r_0_10 ) );
  DFF_X1 key_b_r_reg_0_11 (.CK( clk ) , .D( key2[11] ) , .Q( key_b_r_0_11 ) );
  DFF_X1 key_b_r_reg_0_12 (.CK( clk ) , .D( key2[12] ) , .Q( key_b_r_0_12 ) );
  DFF_X1 key_b_r_reg_0_13 (.CK( clk ) , .D( key2[13] ) , .Q( key_b_r_0_13 ) );
  DFF_X1 key_b_r_reg_0_14 (.CK( clk ) , .D( key2[14] ) , .Q( key_b_r_0_14 ) );
  DFF_X1 key_b_r_reg_0_15 (.CK( clk ) , .D( key2[15] ) , .Q( key_b_r_0_15 ) );
  DFF_X1 key_b_r_reg_0_16 (.CK( clk ) , .D( key2[16] ) , .Q( key_b_r_0_16 ) );
  DFF_X1 key_b_r_reg_0_17 (.CK( clk ) , .D( key2[17] ) , .Q( key_b_r_0_17 ) );
  DFF_X1 key_b_r_reg_0_18 (.CK( clk ) , .D( key2[18] ) , .Q( key_b_r_0_18 ) );
  DFF_X1 key_b_r_reg_0_19 (.CK( clk ) , .D( key2[19] ) , .Q( key_b_r_0_19 ) );
  DFF_X1 key_b_r_reg_0_2 (.CK( clk ) , .D( key2[2] ) , .Q( key_b_r_0_2 ) );
  DFF_X1 key_b_r_reg_0_20 (.CK( clk ) , .D( key2[20] ) , .Q( key_b_r_0_20 ) );
  DFF_X1 key_b_r_reg_0_21 (.CK( clk ) , .D( key2[21] ) , .Q( key_b_r_0_21 ) );
  DFF_X1 key_b_r_reg_0_22 (.CK( clk ) , .D( key2[22] ) , .Q( key_b_r_0_22 ) );
  DFF_X1 key_b_r_reg_0_23 (.CK( clk ) , .D( key2[23] ) , .Q( key_b_r_0_23 ) );
  DFF_X1 key_b_r_reg_0_24 (.CK( clk ) , .D( key2[24] ) , .Q( key_b_r_0_24 ) );
  DFF_X1 key_b_r_reg_0_25 (.CK( clk ) , .D( key2[25] ) , .Q( key_b_r_0_25 ) );
  DFF_X1 key_b_r_reg_0_26 (.CK( clk ) , .D( key2[26] ) , .Q( key_b_r_0_26 ) );
  DFF_X1 key_b_r_reg_0_27 (.CK( clk ) , .D( key2[27] ) , .Q( key_b_r_0_27 ) );
  DFF_X1 key_b_r_reg_0_28 (.CK( clk ) , .D( key2[28] ) , .Q( key_b_r_0_28 ) );
  DFF_X1 key_b_r_reg_0_29 (.CK( clk ) , .D( key2[29] ) , .Q( key_b_r_0_29 ) );
  DFF_X1 key_b_r_reg_0_3 (.CK( clk ) , .D( key2[3] ) , .Q( key_b_r_0_3 ) );
  DFF_X1 key_b_r_reg_0_30 (.CK( clk ) , .D( key2[30] ) , .Q( key_b_r_0_30 ) );
  DFF_X1 key_b_r_reg_0_31 (.CK( clk ) , .D( key2[31] ) , .Q( key_b_r_0_31 ) );
  DFF_X1 key_b_r_reg_0_32 (.CK( clk ) , .D( key2[32] ) , .Q( key_b_r_0_32 ) );
  DFF_X1 key_b_r_reg_0_33 (.CK( clk ) , .D( key2[33] ) , .Q( key_b_r_0_33 ) );
  DFF_X1 key_b_r_reg_0_34 (.CK( clk ) , .D( key2[34] ) , .Q( key_b_r_0_34 ) );
  DFF_X1 key_b_r_reg_0_35 (.CK( clk ) , .D( key2[35] ) , .Q( key_b_r_0_35 ) );
  DFF_X1 key_b_r_reg_0_36 (.CK( clk ) , .D( key2[36] ) , .Q( key_b_r_0_36 ) );
  DFF_X1 key_b_r_reg_0_37 (.CK( clk ) , .D( key2[37] ) , .Q( key_b_r_0_37 ) );
  DFF_X1 key_b_r_reg_0_38 (.CK( clk ) , .D( key2[38] ) , .Q( key_b_r_0_38 ) );
  DFF_X1 key_b_r_reg_0_39 (.CK( clk ) , .D( key2[39] ) , .Q( key_b_r_0_39 ) );
  DFF_X1 key_b_r_reg_0_4 (.CK( clk ) , .D( key2[4] ) , .Q( key_b_r_0_4 ) );
  DFF_X1 key_b_r_reg_0_40 (.CK( clk ) , .D( key2[40] ) , .Q( key_b_r_0_40 ) );
  DFF_X1 key_b_r_reg_0_41 (.CK( clk ) , .D( key2[41] ) , .Q( key_b_r_0_41 ) );
  DFF_X1 key_b_r_reg_0_42 (.CK( clk ) , .D( key2[42] ) , .Q( key_b_r_0_42 ) );
  DFF_X1 key_b_r_reg_0_43 (.CK( clk ) , .D( key2[43] ) , .Q( key_b_r_0_43 ) );
  DFF_X1 key_b_r_reg_0_44 (.CK( clk ) , .D( key2[44] ) , .Q( key_b_r_0_44 ) );
  DFF_X1 key_b_r_reg_0_45 (.CK( clk ) , .D( key2[45] ) , .Q( key_b_r_0_45 ) );
  DFF_X1 key_b_r_reg_0_46 (.CK( clk ) , .D( key2[46] ) , .Q( key_b_r_0_46 ) );
  DFF_X1 key_b_r_reg_0_47 (.CK( clk ) , .D( key2[47] ) , .Q( key_b_r_0_47 ) );
  DFF_X1 key_b_r_reg_0_48 (.CK( clk ) , .D( key2[48] ) , .Q( key_b_r_0_48 ) );
  DFF_X1 key_b_r_reg_0_49 (.CK( clk ) , .D( key2[49] ) , .Q( key_b_r_0_49 ) );
  DFF_X1 key_b_r_reg_0_5 (.CK( clk ) , .D( key2[5] ) , .Q( key_b_r_0_5 ) );
  DFF_X1 key_b_r_reg_0_50 (.CK( clk ) , .D( key2[50] ) , .Q( key_b_r_0_50 ) );
  DFF_X1 key_b_r_reg_0_51 (.CK( clk ) , .D( key2[51] ) , .Q( key_b_r_0_51 ) );
  DFF_X1 key_b_r_reg_0_52 (.CK( clk ) , .D( key2[52] ) , .Q( key_b_r_0_52 ) );
  DFF_X1 key_b_r_reg_0_53 (.CK( clk ) , .D( key2[53] ) , .Q( key_b_r_0_53 ) );
  DFF_X1 key_b_r_reg_0_54 (.CK( clk ) , .D( key2[54] ) , .Q( key_b_r_0_54 ) );
  DFF_X1 key_b_r_reg_0_55 (.CK( clk ) , .D( key2[55] ) , .Q( key_b_r_0_55 ) );
  DFF_X1 key_b_r_reg_0_6 (.CK( clk ) , .D( key2[6] ) , .Q( key_b_r_0_6 ) );
  DFF_X1 key_b_r_reg_0_7 (.CK( clk ) , .D( key2[7] ) , .Q( key_b_r_0_7 ) );
  DFF_X1 key_b_r_reg_0_8 (.CK( clk ) , .D( key2[8] ) , .Q( key_b_r_0_8 ) );
  DFF_X1 key_b_r_reg_0_9 (.CK( clk ) , .D( key2[9] ) , .Q( key_b_r_0_9 ) );
  DFF_X1 key_b_r_reg_10_0 (.CK( clk ) , .Q( key_b_r_10_0 ) , .D( key_b_r_9_0 ) );
  DFF_X1 key_b_r_reg_10_1 (.CK( clk ) , .Q( key_b_r_10_1 ) , .D( key_b_r_9_1 ) );
  DFF_X1 key_b_r_reg_10_10 (.CK( clk ) , .Q( key_b_r_10_10 ) , .D( key_b_r_9_10 ) );
  DFF_X1 key_b_r_reg_10_11 (.CK( clk ) , .Q( key_b_r_10_11 ) , .D( key_b_r_9_11 ) );
  DFF_X1 key_b_r_reg_10_12 (.CK( clk ) , .Q( key_b_r_10_12 ) , .D( key_b_r_9_12 ) );
  DFF_X1 key_b_r_reg_10_13 (.CK( clk ) , .Q( key_b_r_10_13 ) , .D( key_b_r_9_13 ) );
  DFF_X1 key_b_r_reg_10_14 (.CK( clk ) , .Q( key_b_r_10_14 ) , .D( key_b_r_9_14 ) );
  DFF_X1 key_b_r_reg_10_15 (.CK( clk ) , .Q( key_b_r_10_15 ) , .D( key_b_r_9_15 ) );
  DFF_X1 key_b_r_reg_10_16 (.CK( clk ) , .Q( key_b_r_10_16 ) , .D( key_b_r_9_16 ) );
  DFF_X1 key_b_r_reg_10_17 (.CK( clk ) , .Q( key_b_r_10_17 ) , .D( key_b_r_9_17 ) );
  DFF_X1 key_b_r_reg_10_18 (.CK( clk ) , .Q( key_b_r_10_18 ) , .D( key_b_r_9_18 ) );
  DFF_X1 key_b_r_reg_10_19 (.CK( clk ) , .Q( key_b_r_10_19 ) , .D( key_b_r_9_19 ) );
  DFF_X1 key_b_r_reg_10_2 (.CK( clk ) , .Q( key_b_r_10_2 ) , .D( key_b_r_9_2 ) );
  DFF_X1 key_b_r_reg_10_20 (.CK( clk ) , .Q( key_b_r_10_20 ) , .D( key_b_r_9_20 ) );
  DFF_X1 key_b_r_reg_10_21 (.CK( clk ) , .Q( key_b_r_10_21 ) , .D( key_b_r_9_21 ) );
  DFF_X1 key_b_r_reg_10_22 (.CK( clk ) , .Q( key_b_r_10_22 ) , .D( key_b_r_9_22 ) );
  DFF_X1 key_b_r_reg_10_23 (.CK( clk ) , .Q( key_b_r_10_23 ) , .D( key_b_r_9_23 ) );
  DFF_X1 key_b_r_reg_10_24 (.CK( clk ) , .Q( key_b_r_10_24 ) , .D( key_b_r_9_24 ) );
  DFF_X1 key_b_r_reg_10_25 (.CK( clk ) , .Q( key_b_r_10_25 ) , .D( key_b_r_9_25 ) );
  DFF_X1 key_b_r_reg_10_26 (.CK( clk ) , .Q( key_b_r_10_26 ) , .D( key_b_r_9_26 ) );
  DFF_X1 key_b_r_reg_10_27 (.CK( clk ) , .Q( key_b_r_10_27 ) , .D( key_b_r_9_27 ) );
  DFF_X1 key_b_r_reg_10_28 (.CK( clk ) , .Q( key_b_r_10_28 ) , .D( key_b_r_9_28 ) );
  DFF_X1 key_b_r_reg_10_29 (.CK( clk ) , .Q( key_b_r_10_29 ) , .D( key_b_r_9_29 ) );
  DFF_X1 key_b_r_reg_10_3 (.CK( clk ) , .Q( key_b_r_10_3 ) , .D( key_b_r_9_3 ) );
  DFF_X1 key_b_r_reg_10_30 (.CK( clk ) , .Q( key_b_r_10_30 ) , .D( key_b_r_9_30 ) );
  DFF_X1 key_b_r_reg_10_31 (.CK( clk ) , .Q( key_b_r_10_31 ) , .D( key_b_r_9_31 ) );
  DFF_X1 key_b_r_reg_10_32 (.CK( clk ) , .Q( key_b_r_10_32 ) , .D( key_b_r_9_32 ) );
  DFF_X1 key_b_r_reg_10_33 (.CK( clk ) , .Q( key_b_r_10_33 ) , .D( key_b_r_9_33 ) );
  DFF_X1 key_b_r_reg_10_34 (.CK( clk ) , .Q( key_b_r_10_34 ) , .D( key_b_r_9_34 ) );
  DFF_X1 key_b_r_reg_10_35 (.CK( clk ) , .Q( key_b_r_10_35 ) , .D( key_b_r_9_35 ) );
  DFF_X1 key_b_r_reg_10_36 (.CK( clk ) , .Q( key_b_r_10_36 ) , .D( key_b_r_9_36 ) );
  DFF_X1 key_b_r_reg_10_37 (.CK( clk ) , .Q( key_b_r_10_37 ) , .D( key_b_r_9_37 ) );
  DFF_X1 key_b_r_reg_10_38 (.CK( clk ) , .Q( key_b_r_10_38 ) , .D( key_b_r_9_38 ) );
  DFF_X1 key_b_r_reg_10_39 (.CK( clk ) , .Q( key_b_r_10_39 ) , .D( key_b_r_9_39 ) );
  DFF_X1 key_b_r_reg_10_4 (.CK( clk ) , .Q( key_b_r_10_4 ) , .D( key_b_r_9_4 ) );
  DFF_X1 key_b_r_reg_10_40 (.CK( clk ) , .Q( key_b_r_10_40 ) , .D( key_b_r_9_40 ) );
  DFF_X1 key_b_r_reg_10_41 (.CK( clk ) , .Q( key_b_r_10_41 ) , .D( key_b_r_9_41 ) );
  DFF_X1 key_b_r_reg_10_42 (.CK( clk ) , .Q( key_b_r_10_42 ) , .D( key_b_r_9_42 ) );
  DFF_X1 key_b_r_reg_10_43 (.CK( clk ) , .Q( key_b_r_10_43 ) , .D( key_b_r_9_43 ) );
  DFF_X1 key_b_r_reg_10_44 (.CK( clk ) , .Q( key_b_r_10_44 ) , .D( key_b_r_9_44 ) );
  DFF_X1 key_b_r_reg_10_45 (.CK( clk ) , .Q( key_b_r_10_45 ) , .D( key_b_r_9_45 ) );
  DFF_X1 key_b_r_reg_10_46 (.CK( clk ) , .Q( key_b_r_10_46 ) , .D( key_b_r_9_46 ) );
  DFF_X1 key_b_r_reg_10_47 (.CK( clk ) , .Q( key_b_r_10_47 ) , .D( key_b_r_9_47 ) );
  DFF_X1 key_b_r_reg_10_48 (.CK( clk ) , .Q( key_b_r_10_48 ) , .D( key_b_r_9_48 ) );
  DFF_X1 key_b_r_reg_10_49 (.CK( clk ) , .Q( key_b_r_10_49 ) , .D( key_b_r_9_49 ) );
  DFF_X1 key_b_r_reg_10_5 (.CK( clk ) , .Q( key_b_r_10_5 ) , .D( key_b_r_9_5 ) );
  DFF_X1 key_b_r_reg_10_50 (.CK( clk ) , .Q( key_b_r_10_50 ) , .D( key_b_r_9_50 ) );
  DFF_X1 key_b_r_reg_10_51 (.CK( clk ) , .Q( key_b_r_10_51 ) , .D( key_b_r_9_51 ) );
  DFF_X1 key_b_r_reg_10_52 (.CK( clk ) , .Q( key_b_r_10_52 ) , .D( key_b_r_9_52 ) );
  DFF_X1 key_b_r_reg_10_53 (.CK( clk ) , .Q( key_b_r_10_53 ) , .D( key_b_r_9_53 ) );
  DFF_X1 key_b_r_reg_10_54 (.CK( clk ) , .Q( key_b_r_10_54 ) , .D( key_b_r_9_54 ) );
  DFF_X1 key_b_r_reg_10_55 (.CK( clk ) , .Q( key_b_r_10_55 ) , .D( key_b_r_9_55 ) );
  DFF_X1 key_b_r_reg_10_6 (.CK( clk ) , .Q( key_b_r_10_6 ) , .D( key_b_r_9_6 ) );
  DFF_X1 key_b_r_reg_10_7 (.CK( clk ) , .Q( key_b_r_10_7 ) , .D( key_b_r_9_7 ) );
  DFF_X1 key_b_r_reg_10_8 (.CK( clk ) , .Q( key_b_r_10_8 ) , .D( key_b_r_9_8 ) );
  DFF_X1 key_b_r_reg_10_9 (.CK( clk ) , .Q( key_b_r_10_9 ) , .D( key_b_r_9_9 ) );
  DFF_X1 key_b_r_reg_11_0 (.CK( clk ) , .D( key_b_r_10_0 ) , .Q( key_b_r_11_0 ) );
  DFF_X1 key_b_r_reg_11_1 (.CK( clk ) , .D( key_b_r_10_1 ) , .Q( key_b_r_11_1 ) );
  DFF_X1 key_b_r_reg_11_10 (.CK( clk ) , .D( key_b_r_10_10 ) , .Q( key_b_r_11_10 ) );
  DFF_X1 key_b_r_reg_11_11 (.CK( clk ) , .D( key_b_r_10_11 ) , .Q( key_b_r_11_11 ) );
  DFF_X1 key_b_r_reg_11_12 (.CK( clk ) , .D( key_b_r_10_12 ) , .Q( key_b_r_11_12 ) );
  DFF_X1 key_b_r_reg_11_13 (.CK( clk ) , .D( key_b_r_10_13 ) , .Q( key_b_r_11_13 ) );
  DFF_X1 key_b_r_reg_11_14 (.CK( clk ) , .D( key_b_r_10_14 ) , .Q( key_b_r_11_14 ) );
  DFF_X1 key_b_r_reg_11_15 (.CK( clk ) , .D( key_b_r_10_15 ) , .Q( key_b_r_11_15 ) );
  DFF_X1 key_b_r_reg_11_16 (.CK( clk ) , .D( key_b_r_10_16 ) , .Q( key_b_r_11_16 ) );
  DFF_X1 key_b_r_reg_11_17 (.CK( clk ) , .D( key_b_r_10_17 ) , .Q( key_b_r_11_17 ) );
  DFF_X1 key_b_r_reg_11_18 (.CK( clk ) , .D( key_b_r_10_18 ) , .Q( key_b_r_11_18 ) );
  DFF_X1 key_b_r_reg_11_19 (.CK( clk ) , .D( key_b_r_10_19 ) , .Q( key_b_r_11_19 ) );
  DFF_X1 key_b_r_reg_11_2 (.CK( clk ) , .D( key_b_r_10_2 ) , .Q( key_b_r_11_2 ) );
  DFF_X1 key_b_r_reg_11_20 (.CK( clk ) , .D( key_b_r_10_20 ) , .Q( key_b_r_11_20 ) );
  DFF_X1 key_b_r_reg_11_21 (.CK( clk ) , .D( key_b_r_10_21 ) , .Q( key_b_r_11_21 ) );
  DFF_X1 key_b_r_reg_11_22 (.CK( clk ) , .D( key_b_r_10_22 ) , .Q( key_b_r_11_22 ) );
  DFF_X1 key_b_r_reg_11_23 (.CK( clk ) , .D( key_b_r_10_23 ) , .Q( key_b_r_11_23 ) );
  DFF_X1 key_b_r_reg_11_24 (.CK( clk ) , .D( key_b_r_10_24 ) , .Q( key_b_r_11_24 ) );
  DFF_X1 key_b_r_reg_11_25 (.CK( clk ) , .D( key_b_r_10_25 ) , .Q( key_b_r_11_25 ) );
  DFF_X1 key_b_r_reg_11_26 (.CK( clk ) , .D( key_b_r_10_26 ) , .Q( key_b_r_11_26 ) );
  DFF_X1 key_b_r_reg_11_27 (.CK( clk ) , .D( key_b_r_10_27 ) , .Q( key_b_r_11_27 ) );
  DFF_X1 key_b_r_reg_11_28 (.CK( clk ) , .D( key_b_r_10_28 ) , .Q( key_b_r_11_28 ) );
  DFF_X1 key_b_r_reg_11_29 (.CK( clk ) , .D( key_b_r_10_29 ) , .Q( key_b_r_11_29 ) );
  DFF_X1 key_b_r_reg_11_3 (.CK( clk ) , .D( key_b_r_10_3 ) , .Q( key_b_r_11_3 ) );
  DFF_X1 key_b_r_reg_11_30 (.CK( clk ) , .D( key_b_r_10_30 ) , .Q( key_b_r_11_30 ) );
  DFF_X1 key_b_r_reg_11_31 (.CK( clk ) , .D( key_b_r_10_31 ) , .Q( key_b_r_11_31 ) );
  DFF_X1 key_b_r_reg_11_32 (.CK( clk ) , .D( key_b_r_10_32 ) , .Q( key_b_r_11_32 ) );
  DFF_X1 key_b_r_reg_11_33 (.CK( clk ) , .D( key_b_r_10_33 ) , .Q( key_b_r_11_33 ) );
  DFF_X1 key_b_r_reg_11_34 (.CK( clk ) , .D( key_b_r_10_34 ) , .Q( key_b_r_11_34 ) );
  DFF_X1 key_b_r_reg_11_35 (.CK( clk ) , .D( key_b_r_10_35 ) , .Q( key_b_r_11_35 ) );
  DFF_X1 key_b_r_reg_11_36 (.CK( clk ) , .D( key_b_r_10_36 ) , .Q( key_b_r_11_36 ) );
  DFF_X1 key_b_r_reg_11_37 (.CK( clk ) , .D( key_b_r_10_37 ) , .Q( key_b_r_11_37 ) );
  DFF_X1 key_b_r_reg_11_38 (.CK( clk ) , .D( key_b_r_10_38 ) , .Q( key_b_r_11_38 ) );
  DFF_X1 key_b_r_reg_11_39 (.CK( clk ) , .D( key_b_r_10_39 ) , .Q( key_b_r_11_39 ) );
  DFF_X1 key_b_r_reg_11_4 (.CK( clk ) , .D( key_b_r_10_4 ) , .Q( key_b_r_11_4 ) );
  DFF_X1 key_b_r_reg_11_40 (.CK( clk ) , .D( key_b_r_10_40 ) , .Q( key_b_r_11_40 ) );
  DFF_X1 key_b_r_reg_11_41 (.CK( clk ) , .D( key_b_r_10_41 ) , .Q( key_b_r_11_41 ) );
  DFF_X1 key_b_r_reg_11_42 (.CK( clk ) , .D( key_b_r_10_42 ) , .Q( key_b_r_11_42 ) );
  DFF_X1 key_b_r_reg_11_43 (.CK( clk ) , .D( key_b_r_10_43 ) , .Q( key_b_r_11_43 ) );
  DFF_X1 key_b_r_reg_11_44 (.CK( clk ) , .D( key_b_r_10_44 ) , .Q( key_b_r_11_44 ) );
  DFF_X1 key_b_r_reg_11_45 (.CK( clk ) , .D( key_b_r_10_45 ) , .Q( key_b_r_11_45 ) );
  DFF_X1 key_b_r_reg_11_46 (.CK( clk ) , .D( key_b_r_10_46 ) , .Q( key_b_r_11_46 ) );
  DFF_X1 key_b_r_reg_11_47 (.CK( clk ) , .D( key_b_r_10_47 ) , .Q( key_b_r_11_47 ) );
  DFF_X1 key_b_r_reg_11_48 (.CK( clk ) , .D( key_b_r_10_48 ) , .Q( key_b_r_11_48 ) );
  DFF_X1 key_b_r_reg_11_49 (.CK( clk ) , .D( key_b_r_10_49 ) , .Q( key_b_r_11_49 ) );
  DFF_X1 key_b_r_reg_11_5 (.CK( clk ) , .D( key_b_r_10_5 ) , .Q( key_b_r_11_5 ) );
  DFF_X1 key_b_r_reg_11_50 (.CK( clk ) , .D( key_b_r_10_50 ) , .Q( key_b_r_11_50 ) );
  DFF_X1 key_b_r_reg_11_51 (.CK( clk ) , .D( key_b_r_10_51 ) , .Q( key_b_r_11_51 ) );
  DFF_X1 key_b_r_reg_11_52 (.CK( clk ) , .D( key_b_r_10_52 ) , .Q( key_b_r_11_52 ) );
  DFF_X1 key_b_r_reg_11_53 (.CK( clk ) , .D( key_b_r_10_53 ) , .Q( key_b_r_11_53 ) );
  DFF_X1 key_b_r_reg_11_54 (.CK( clk ) , .D( key_b_r_10_54 ) , .Q( key_b_r_11_54 ) );
  DFF_X1 key_b_r_reg_11_55 (.CK( clk ) , .D( key_b_r_10_55 ) , .Q( key_b_r_11_55 ) );
  DFF_X1 key_b_r_reg_11_6 (.CK( clk ) , .D( key_b_r_10_6 ) , .Q( key_b_r_11_6 ) );
  DFF_X1 key_b_r_reg_11_7 (.CK( clk ) , .D( key_b_r_10_7 ) , .Q( key_b_r_11_7 ) );
  DFF_X1 key_b_r_reg_11_8 (.CK( clk ) , .D( key_b_r_10_8 ) , .Q( key_b_r_11_8 ) );
  DFF_X1 key_b_r_reg_11_9 (.CK( clk ) , .D( key_b_r_10_9 ) , .Q( key_b_r_11_9 ) );
  DFF_X1 key_b_r_reg_12_0 (.CK( clk ) , .D( key_b_r_11_0 ) , .Q( key_b_r_12_0 ) );
  DFF_X1 key_b_r_reg_12_1 (.CK( clk ) , .D( key_b_r_11_1 ) , .Q( key_b_r_12_1 ) );
  DFF_X1 key_b_r_reg_12_10 (.CK( clk ) , .D( key_b_r_11_10 ) , .Q( key_b_r_12_10 ) );
  DFF_X1 key_b_r_reg_12_11 (.CK( clk ) , .D( key_b_r_11_11 ) , .Q( key_b_r_12_11 ) );
  DFF_X1 key_b_r_reg_12_12 (.CK( clk ) , .D( key_b_r_11_12 ) , .Q( key_b_r_12_12 ) );
  DFF_X1 key_b_r_reg_12_13 (.CK( clk ) , .D( key_b_r_11_13 ) , .Q( key_b_r_12_13 ) );
  DFF_X1 key_b_r_reg_12_14 (.CK( clk ) , .D( key_b_r_11_14 ) , .Q( key_b_r_12_14 ) );
  DFF_X1 key_b_r_reg_12_15 (.CK( clk ) , .D( key_b_r_11_15 ) , .Q( key_b_r_12_15 ) );
  DFF_X1 key_b_r_reg_12_16 (.CK( clk ) , .D( key_b_r_11_16 ) , .Q( key_b_r_12_16 ) );
  DFF_X1 key_b_r_reg_12_17 (.CK( clk ) , .D( key_b_r_11_17 ) , .Q( key_b_r_12_17 ) );
  DFF_X1 key_b_r_reg_12_18 (.CK( clk ) , .D( key_b_r_11_18 ) , .Q( key_b_r_12_18 ) );
  DFF_X1 key_b_r_reg_12_19 (.CK( clk ) , .D( key_b_r_11_19 ) , .Q( key_b_r_12_19 ) );
  DFF_X1 key_b_r_reg_12_2 (.CK( clk ) , .D( key_b_r_11_2 ) , .Q( key_b_r_12_2 ) );
  DFF_X1 key_b_r_reg_12_20 (.CK( clk ) , .D( key_b_r_11_20 ) , .Q( key_b_r_12_20 ) );
  DFF_X1 key_b_r_reg_12_21 (.CK( clk ) , .D( key_b_r_11_21 ) , .Q( key_b_r_12_21 ) );
  DFF_X1 key_b_r_reg_12_22 (.CK( clk ) , .D( key_b_r_11_22 ) , .Q( key_b_r_12_22 ) );
  DFF_X1 key_b_r_reg_12_23 (.CK( clk ) , .D( key_b_r_11_23 ) , .Q( key_b_r_12_23 ) );
  DFF_X1 key_b_r_reg_12_24 (.CK( clk ) , .D( key_b_r_11_24 ) , .Q( key_b_r_12_24 ) );
  DFF_X1 key_b_r_reg_12_25 (.CK( clk ) , .D( key_b_r_11_25 ) , .Q( key_b_r_12_25 ) );
  DFF_X1 key_b_r_reg_12_26 (.CK( clk ) , .D( key_b_r_11_26 ) , .Q( key_b_r_12_26 ) );
  DFF_X1 key_b_r_reg_12_27 (.CK( clk ) , .D( key_b_r_11_27 ) , .Q( key_b_r_12_27 ) );
  DFF_X1 key_b_r_reg_12_28 (.CK( clk ) , .D( key_b_r_11_28 ) , .Q( key_b_r_12_28 ) );
  DFF_X1 key_b_r_reg_12_29 (.CK( clk ) , .D( key_b_r_11_29 ) , .Q( key_b_r_12_29 ) );
  DFF_X1 key_b_r_reg_12_3 (.CK( clk ) , .D( key_b_r_11_3 ) , .Q( key_b_r_12_3 ) );
  DFF_X1 key_b_r_reg_12_30 (.CK( clk ) , .D( key_b_r_11_30 ) , .Q( key_b_r_12_30 ) );
  DFF_X1 key_b_r_reg_12_31 (.CK( clk ) , .D( key_b_r_11_31 ) , .Q( key_b_r_12_31 ) );
  DFF_X1 key_b_r_reg_12_32 (.CK( clk ) , .D( key_b_r_11_32 ) , .Q( key_b_r_12_32 ) );
  DFF_X1 key_b_r_reg_12_33 (.CK( clk ) , .D( key_b_r_11_33 ) , .Q( key_b_r_12_33 ) );
  DFF_X1 key_b_r_reg_12_34 (.CK( clk ) , .D( key_b_r_11_34 ) , .Q( key_b_r_12_34 ) );
  DFF_X1 key_b_r_reg_12_35 (.CK( clk ) , .D( key_b_r_11_35 ) , .Q( key_b_r_12_35 ) );
  DFF_X1 key_b_r_reg_12_36 (.CK( clk ) , .D( key_b_r_11_36 ) , .Q( key_b_r_12_36 ) );
  DFF_X1 key_b_r_reg_12_37 (.CK( clk ) , .D( key_b_r_11_37 ) , .Q( key_b_r_12_37 ) );
  DFF_X1 key_b_r_reg_12_38 (.CK( clk ) , .D( key_b_r_11_38 ) , .Q( key_b_r_12_38 ) );
  DFF_X1 key_b_r_reg_12_39 (.CK( clk ) , .D( key_b_r_11_39 ) , .Q( key_b_r_12_39 ) );
  DFF_X1 key_b_r_reg_12_4 (.CK( clk ) , .D( key_b_r_11_4 ) , .Q( key_b_r_12_4 ) );
  DFF_X1 key_b_r_reg_12_40 (.CK( clk ) , .D( key_b_r_11_40 ) , .Q( key_b_r_12_40 ) );
  DFF_X1 key_b_r_reg_12_41 (.CK( clk ) , .D( key_b_r_11_41 ) , .Q( key_b_r_12_41 ) );
  DFF_X1 key_b_r_reg_12_42 (.CK( clk ) , .D( key_b_r_11_42 ) , .Q( key_b_r_12_42 ) );
  DFF_X1 key_b_r_reg_12_43 (.CK( clk ) , .D( key_b_r_11_43 ) , .Q( key_b_r_12_43 ) );
  DFF_X1 key_b_r_reg_12_44 (.CK( clk ) , .D( key_b_r_11_44 ) , .Q( key_b_r_12_44 ) );
  DFF_X1 key_b_r_reg_12_45 (.CK( clk ) , .D( key_b_r_11_45 ) , .Q( key_b_r_12_45 ) );
  DFF_X1 key_b_r_reg_12_46 (.CK( clk ) , .D( key_b_r_11_46 ) , .Q( key_b_r_12_46 ) );
  DFF_X1 key_b_r_reg_12_47 (.CK( clk ) , .D( key_b_r_11_47 ) , .Q( key_b_r_12_47 ) );
  DFF_X1 key_b_r_reg_12_48 (.CK( clk ) , .D( key_b_r_11_48 ) , .Q( key_b_r_12_48 ) );
  DFF_X1 key_b_r_reg_12_49 (.CK( clk ) , .D( key_b_r_11_49 ) , .Q( key_b_r_12_49 ) );
  DFF_X1 key_b_r_reg_12_5 (.CK( clk ) , .D( key_b_r_11_5 ) , .Q( key_b_r_12_5 ) );
  DFF_X1 key_b_r_reg_12_50 (.CK( clk ) , .D( key_b_r_11_50 ) , .Q( key_b_r_12_50 ) );
  DFF_X1 key_b_r_reg_12_51 (.CK( clk ) , .D( key_b_r_11_51 ) , .Q( key_b_r_12_51 ) );
  DFF_X1 key_b_r_reg_12_52 (.CK( clk ) , .D( key_b_r_11_52 ) , .Q( key_b_r_12_52 ) );
  DFF_X1 key_b_r_reg_12_53 (.CK( clk ) , .D( key_b_r_11_53 ) , .Q( key_b_r_12_53 ) );
  DFF_X1 key_b_r_reg_12_54 (.CK( clk ) , .D( key_b_r_11_54 ) , .Q( key_b_r_12_54 ) );
  DFF_X1 key_b_r_reg_12_55 (.CK( clk ) , .D( key_b_r_11_55 ) , .Q( key_b_r_12_55 ) );
  DFF_X1 key_b_r_reg_12_6 (.CK( clk ) , .D( key_b_r_11_6 ) , .Q( key_b_r_12_6 ) );
  DFF_X1 key_b_r_reg_12_7 (.CK( clk ) , .D( key_b_r_11_7 ) , .Q( key_b_r_12_7 ) );
  DFF_X1 key_b_r_reg_12_8 (.CK( clk ) , .D( key_b_r_11_8 ) , .Q( key_b_r_12_8 ) );
  DFF_X1 key_b_r_reg_12_9 (.CK( clk ) , .D( key_b_r_11_9 ) , .Q( key_b_r_12_9 ) );
  DFF_X1 key_b_r_reg_13_0 (.CK( clk ) , .D( key_b_r_12_0 ) , .Q( key_b_r_13_0 ) );
  DFF_X1 key_b_r_reg_13_1 (.CK( clk ) , .D( key_b_r_12_1 ) , .Q( key_b_r_13_1 ) );
  DFF_X1 key_b_r_reg_13_10 (.CK( clk ) , .D( key_b_r_12_10 ) , .Q( key_b_r_13_10 ) );
  DFF_X1 key_b_r_reg_13_11 (.CK( clk ) , .D( key_b_r_12_11 ) , .Q( key_b_r_13_11 ) );
  DFF_X1 key_b_r_reg_13_12 (.CK( clk ) , .D( key_b_r_12_12 ) , .Q( key_b_r_13_12 ) );
  DFF_X1 key_b_r_reg_13_13 (.CK( clk ) , .D( key_b_r_12_13 ) , .Q( key_b_r_13_13 ) );
  DFF_X1 key_b_r_reg_13_14 (.CK( clk ) , .D( key_b_r_12_14 ) , .Q( key_b_r_13_14 ) );
  DFF_X1 key_b_r_reg_13_15 (.CK( clk ) , .D( key_b_r_12_15 ) , .Q( key_b_r_13_15 ) );
  DFF_X1 key_b_r_reg_13_16 (.CK( clk ) , .D( key_b_r_12_16 ) , .Q( key_b_r_13_16 ) );
  DFF_X1 key_b_r_reg_13_17 (.CK( clk ) , .D( key_b_r_12_17 ) , .Q( key_b_r_13_17 ) );
  DFF_X1 key_b_r_reg_13_18 (.CK( clk ) , .D( key_b_r_12_18 ) , .Q( key_b_r_13_18 ) );
  DFF_X1 key_b_r_reg_13_19 (.CK( clk ) , .D( key_b_r_12_19 ) , .Q( key_b_r_13_19 ) );
  DFF_X1 key_b_r_reg_13_2 (.CK( clk ) , .D( key_b_r_12_2 ) , .Q( key_b_r_13_2 ) );
  DFF_X1 key_b_r_reg_13_20 (.CK( clk ) , .D( key_b_r_12_20 ) , .Q( key_b_r_13_20 ) );
  DFF_X1 key_b_r_reg_13_21 (.CK( clk ) , .D( key_b_r_12_21 ) , .Q( key_b_r_13_21 ) );
  DFF_X1 key_b_r_reg_13_22 (.CK( clk ) , .D( key_b_r_12_22 ) , .Q( key_b_r_13_22 ) );
  DFF_X1 key_b_r_reg_13_23 (.CK( clk ) , .D( key_b_r_12_23 ) , .Q( key_b_r_13_23 ) );
  DFF_X1 key_b_r_reg_13_24 (.CK( clk ) , .D( key_b_r_12_24 ) , .Q( key_b_r_13_24 ) );
  DFF_X1 key_b_r_reg_13_25 (.CK( clk ) , .D( key_b_r_12_25 ) , .Q( key_b_r_13_25 ) );
  DFF_X1 key_b_r_reg_13_26 (.CK( clk ) , .D( key_b_r_12_26 ) , .Q( key_b_r_13_26 ) );
  DFF_X1 key_b_r_reg_13_27 (.CK( clk ) , .D( key_b_r_12_27 ) , .Q( key_b_r_13_27 ) );
  DFF_X1 key_b_r_reg_13_28 (.CK( clk ) , .D( key_b_r_12_28 ) , .Q( key_b_r_13_28 ) );
  DFF_X1 key_b_r_reg_13_29 (.CK( clk ) , .D( key_b_r_12_29 ) , .Q( key_b_r_13_29 ) );
  DFF_X1 key_b_r_reg_13_3 (.CK( clk ) , .D( key_b_r_12_3 ) , .Q( key_b_r_13_3 ) );
  DFF_X1 key_b_r_reg_13_30 (.CK( clk ) , .D( key_b_r_12_30 ) , .Q( key_b_r_13_30 ) );
  DFF_X1 key_b_r_reg_13_31 (.CK( clk ) , .D( key_b_r_12_31 ) , .Q( key_b_r_13_31 ) );
  DFF_X1 key_b_r_reg_13_32 (.CK( clk ) , .D( key_b_r_12_32 ) , .Q( key_b_r_13_32 ) );
  DFF_X1 key_b_r_reg_13_33 (.CK( clk ) , .D( key_b_r_12_33 ) , .Q( key_b_r_13_33 ) );
  DFF_X1 key_b_r_reg_13_34 (.CK( clk ) , .D( key_b_r_12_34 ) , .Q( key_b_r_13_34 ) );
  DFF_X1 key_b_r_reg_13_35 (.CK( clk ) , .D( key_b_r_12_35 ) , .Q( key_b_r_13_35 ) );
  DFF_X1 key_b_r_reg_13_36 (.CK( clk ) , .D( key_b_r_12_36 ) , .Q( key_b_r_13_36 ) );
  DFF_X1 key_b_r_reg_13_37 (.CK( clk ) , .D( key_b_r_12_37 ) , .Q( key_b_r_13_37 ) );
  DFF_X1 key_b_r_reg_13_38 (.CK( clk ) , .D( key_b_r_12_38 ) , .Q( key_b_r_13_38 ) );
  DFF_X1 key_b_r_reg_13_39 (.CK( clk ) , .D( key_b_r_12_39 ) , .Q( key_b_r_13_39 ) );
  DFF_X1 key_b_r_reg_13_4 (.CK( clk ) , .D( key_b_r_12_4 ) , .Q( key_b_r_13_4 ) );
  DFF_X1 key_b_r_reg_13_40 (.CK( clk ) , .D( key_b_r_12_40 ) , .Q( key_b_r_13_40 ) );
  DFF_X1 key_b_r_reg_13_41 (.CK( clk ) , .D( key_b_r_12_41 ) , .Q( key_b_r_13_41 ) );
  DFF_X1 key_b_r_reg_13_42 (.CK( clk ) , .D( key_b_r_12_42 ) , .Q( key_b_r_13_42 ) );
  DFF_X1 key_b_r_reg_13_43 (.CK( clk ) , .D( key_b_r_12_43 ) , .Q( key_b_r_13_43 ) );
  DFF_X1 key_b_r_reg_13_44 (.CK( clk ) , .D( key_b_r_12_44 ) , .Q( key_b_r_13_44 ) );
  DFF_X1 key_b_r_reg_13_45 (.CK( clk ) , .D( key_b_r_12_45 ) , .Q( key_b_r_13_45 ) );
  DFF_X1 key_b_r_reg_13_46 (.CK( clk ) , .D( key_b_r_12_46 ) , .Q( key_b_r_13_46 ) );
  DFF_X1 key_b_r_reg_13_47 (.CK( clk ) , .D( key_b_r_12_47 ) , .Q( key_b_r_13_47 ) );
  DFF_X1 key_b_r_reg_13_48 (.CK( clk ) , .D( key_b_r_12_48 ) , .Q( key_b_r_13_48 ) );
  DFF_X1 key_b_r_reg_13_49 (.CK( clk ) , .D( key_b_r_12_49 ) , .Q( key_b_r_13_49 ) );
  DFF_X1 key_b_r_reg_13_5 (.CK( clk ) , .D( key_b_r_12_5 ) , .Q( key_b_r_13_5 ) );
  DFF_X1 key_b_r_reg_13_50 (.CK( clk ) , .D( key_b_r_12_50 ) , .Q( key_b_r_13_50 ) );
  DFF_X1 key_b_r_reg_13_51 (.CK( clk ) , .D( key_b_r_12_51 ) , .Q( key_b_r_13_51 ) );
  DFF_X1 key_b_r_reg_13_52 (.CK( clk ) , .D( key_b_r_12_52 ) , .Q( key_b_r_13_52 ) );
  DFF_X1 key_b_r_reg_13_53 (.CK( clk ) , .D( key_b_r_12_53 ) , .Q( key_b_r_13_53 ) );
  DFF_X1 key_b_r_reg_13_54 (.CK( clk ) , .D( key_b_r_12_54 ) , .Q( key_b_r_13_54 ) );
  DFF_X1 key_b_r_reg_13_55 (.CK( clk ) , .D( key_b_r_12_55 ) , .Q( key_b_r_13_55 ) );
  DFF_X1 key_b_r_reg_13_6 (.CK( clk ) , .D( key_b_r_12_6 ) , .Q( key_b_r_13_6 ) );
  DFF_X1 key_b_r_reg_13_7 (.CK( clk ) , .D( key_b_r_12_7 ) , .Q( key_b_r_13_7 ) );
  DFF_X1 key_b_r_reg_13_8 (.CK( clk ) , .D( key_b_r_12_8 ) , .Q( key_b_r_13_8 ) );
  DFF_X1 key_b_r_reg_13_9 (.CK( clk ) , .D( key_b_r_12_9 ) , .Q( key_b_r_13_9 ) );
  DFF_X1 key_b_r_reg_14_0 (.CK( clk ) , .D( key_b_r_13_0 ) , .Q( key_b_r_14_0 ) );
  DFF_X1 key_b_r_reg_14_1 (.CK( clk ) , .D( key_b_r_13_1 ) , .Q( key_b_r_14_1 ) );
  DFF_X1 key_b_r_reg_14_10 (.CK( clk ) , .D( key_b_r_13_10 ) , .Q( key_b_r_14_10 ) );
  DFF_X1 key_b_r_reg_14_11 (.CK( clk ) , .D( key_b_r_13_11 ) , .Q( key_b_r_14_11 ) );
  DFF_X1 key_b_r_reg_14_12 (.CK( clk ) , .D( key_b_r_13_12 ) , .Q( key_b_r_14_12 ) );
  DFF_X1 key_b_r_reg_14_13 (.CK( clk ) , .D( key_b_r_13_13 ) , .Q( key_b_r_14_13 ) );
  DFF_X1 key_b_r_reg_14_14 (.CK( clk ) , .D( key_b_r_13_14 ) , .Q( key_b_r_14_14 ) );
  DFF_X1 key_b_r_reg_14_15 (.CK( clk ) , .D( key_b_r_13_15 ) , .Q( key_b_r_14_15 ) );
  DFF_X1 key_b_r_reg_14_16 (.CK( clk ) , .D( key_b_r_13_16 ) , .Q( key_b_r_14_16 ) );
  DFF_X1 key_b_r_reg_14_17 (.CK( clk ) , .D( key_b_r_13_17 ) , .Q( key_b_r_14_17 ) );
  DFF_X1 key_b_r_reg_14_18 (.CK( clk ) , .D( key_b_r_13_18 ) , .Q( key_b_r_14_18 ) );
  DFF_X1 key_b_r_reg_14_19 (.CK( clk ) , .D( key_b_r_13_19 ) , .Q( key_b_r_14_19 ) );
  DFF_X1 key_b_r_reg_14_2 (.CK( clk ) , .D( key_b_r_13_2 ) , .Q( key_b_r_14_2 ) );
  DFF_X1 key_b_r_reg_14_20 (.CK( clk ) , .D( key_b_r_13_20 ) , .Q( key_b_r_14_20 ) );
  DFF_X1 key_b_r_reg_14_21 (.CK( clk ) , .D( key_b_r_13_21 ) , .Q( key_b_r_14_21 ) );
  DFF_X1 key_b_r_reg_14_22 (.CK( clk ) , .D( key_b_r_13_22 ) , .Q( key_b_r_14_22 ) );
  DFF_X1 key_b_r_reg_14_23 (.CK( clk ) , .D( key_b_r_13_23 ) , .Q( key_b_r_14_23 ) );
  DFF_X1 key_b_r_reg_14_24 (.CK( clk ) , .D( key_b_r_13_24 ) , .Q( key_b_r_14_24 ) );
  DFF_X1 key_b_r_reg_14_25 (.CK( clk ) , .D( key_b_r_13_25 ) , .Q( key_b_r_14_25 ) );
  DFF_X1 key_b_r_reg_14_26 (.CK( clk ) , .D( key_b_r_13_26 ) , .Q( key_b_r_14_26 ) );
  DFF_X1 key_b_r_reg_14_27 (.CK( clk ) , .D( key_b_r_13_27 ) , .Q( key_b_r_14_27 ) );
  DFF_X1 key_b_r_reg_14_28 (.CK( clk ) , .D( key_b_r_13_28 ) , .Q( key_b_r_14_28 ) );
  DFF_X1 key_b_r_reg_14_29 (.CK( clk ) , .D( key_b_r_13_29 ) , .Q( key_b_r_14_29 ) );
  DFF_X1 key_b_r_reg_14_3 (.CK( clk ) , .D( key_b_r_13_3 ) , .Q( key_b_r_14_3 ) );
  DFF_X1 key_b_r_reg_14_30 (.CK( clk ) , .D( key_b_r_13_30 ) , .Q( key_b_r_14_30 ) );
  DFF_X1 key_b_r_reg_14_31 (.CK( clk ) , .D( key_b_r_13_31 ) , .Q( key_b_r_14_31 ) );
  DFF_X1 key_b_r_reg_14_32 (.CK( clk ) , .D( key_b_r_13_32 ) , .Q( key_b_r_14_32 ) );
  DFF_X1 key_b_r_reg_14_33 (.CK( clk ) , .D( key_b_r_13_33 ) , .Q( key_b_r_14_33 ) );
  DFF_X1 key_b_r_reg_14_34 (.CK( clk ) , .D( key_b_r_13_34 ) , .Q( key_b_r_14_34 ) );
  DFF_X1 key_b_r_reg_14_35 (.CK( clk ) , .D( key_b_r_13_35 ) , .Q( key_b_r_14_35 ) );
  DFF_X1 key_b_r_reg_14_36 (.CK( clk ) , .D( key_b_r_13_36 ) , .Q( key_b_r_14_36 ) );
  DFF_X1 key_b_r_reg_14_37 (.CK( clk ) , .D( key_b_r_13_37 ) , .Q( key_b_r_14_37 ) );
  DFF_X1 key_b_r_reg_14_38 (.CK( clk ) , .D( key_b_r_13_38 ) , .Q( key_b_r_14_38 ) );
  DFF_X1 key_b_r_reg_14_39 (.CK( clk ) , .D( key_b_r_13_39 ) , .Q( key_b_r_14_39 ) );
  DFF_X1 key_b_r_reg_14_4 (.CK( clk ) , .D( key_b_r_13_4 ) , .Q( key_b_r_14_4 ) );
  DFF_X1 key_b_r_reg_14_40 (.CK( clk ) , .D( key_b_r_13_40 ) , .Q( key_b_r_14_40 ) );
  DFF_X1 key_b_r_reg_14_41 (.CK( clk ) , .D( key_b_r_13_41 ) , .Q( key_b_r_14_41 ) );
  DFF_X1 key_b_r_reg_14_42 (.CK( clk ) , .D( key_b_r_13_42 ) , .Q( key_b_r_14_42 ) );
  DFF_X1 key_b_r_reg_14_43 (.CK( clk ) , .D( key_b_r_13_43 ) , .Q( key_b_r_14_43 ) );
  DFF_X1 key_b_r_reg_14_44 (.CK( clk ) , .D( key_b_r_13_44 ) , .Q( key_b_r_14_44 ) );
  DFF_X1 key_b_r_reg_14_45 (.CK( clk ) , .D( key_b_r_13_45 ) , .Q( key_b_r_14_45 ) );
  DFF_X1 key_b_r_reg_14_46 (.CK( clk ) , .D( key_b_r_13_46 ) , .Q( key_b_r_14_46 ) );
  DFF_X1 key_b_r_reg_14_47 (.CK( clk ) , .D( key_b_r_13_47 ) , .Q( key_b_r_14_47 ) );
  DFF_X1 key_b_r_reg_14_48 (.CK( clk ) , .D( key_b_r_13_48 ) , .Q( key_b_r_14_48 ) );
  DFF_X1 key_b_r_reg_14_49 (.CK( clk ) , .D( key_b_r_13_49 ) , .Q( key_b_r_14_49 ) );
  DFF_X1 key_b_r_reg_14_5 (.CK( clk ) , .D( key_b_r_13_5 ) , .Q( key_b_r_14_5 ) );
  DFF_X1 key_b_r_reg_14_50 (.CK( clk ) , .D( key_b_r_13_50 ) , .Q( key_b_r_14_50 ) );
  DFF_X1 key_b_r_reg_14_51 (.CK( clk ) , .D( key_b_r_13_51 ) , .Q( key_b_r_14_51 ) );
  DFF_X1 key_b_r_reg_14_52 (.CK( clk ) , .D( key_b_r_13_52 ) , .Q( key_b_r_14_52 ) );
  DFF_X1 key_b_r_reg_14_53 (.CK( clk ) , .D( key_b_r_13_53 ) , .Q( key_b_r_14_53 ) );
  DFF_X1 key_b_r_reg_14_54 (.CK( clk ) , .D( key_b_r_13_54 ) , .Q( key_b_r_14_54 ) );
  DFF_X1 key_b_r_reg_14_55 (.CK( clk ) , .D( key_b_r_13_55 ) , .Q( key_b_r_14_55 ) );
  DFF_X1 key_b_r_reg_14_6 (.CK( clk ) , .D( key_b_r_13_6 ) , .Q( key_b_r_14_6 ) );
  DFF_X1 key_b_r_reg_14_7 (.CK( clk ) , .D( key_b_r_13_7 ) , .Q( key_b_r_14_7 ) );
  DFF_X1 key_b_r_reg_14_8 (.CK( clk ) , .D( key_b_r_13_8 ) , .Q( key_b_r_14_8 ) );
  DFF_X1 key_b_r_reg_14_9 (.CK( clk ) , .D( key_b_r_13_9 ) , .Q( key_b_r_14_9 ) );
  DFF_X1 key_b_r_reg_15_0 (.CK( clk ) , .D( key_b_r_14_0 ) , .Q( key_b_r_15_0 ) );
  DFF_X1 key_b_r_reg_15_1 (.CK( clk ) , .D( key_b_r_14_1 ) , .Q( key_b_r_15_1 ) );
  DFF_X1 key_b_r_reg_15_10 (.CK( clk ) , .D( key_b_r_14_10 ) , .Q( key_b_r_15_10 ) );
  DFF_X1 key_b_r_reg_15_11 (.CK( clk ) , .D( key_b_r_14_11 ) , .Q( key_b_r_15_11 ) );
  DFF_X1 key_b_r_reg_15_12 (.CK( clk ) , .D( key_b_r_14_12 ) , .Q( key_b_r_15_12 ) );
  DFF_X1 key_b_r_reg_15_13 (.CK( clk ) , .D( key_b_r_14_13 ) , .Q( key_b_r_15_13 ) );
  DFF_X1 key_b_r_reg_15_14 (.CK( clk ) , .D( key_b_r_14_14 ) , .Q( key_b_r_15_14 ) );
  DFF_X1 key_b_r_reg_15_15 (.CK( clk ) , .D( key_b_r_14_15 ) , .Q( key_b_r_15_15 ) );
  DFF_X1 key_b_r_reg_15_16 (.CK( clk ) , .D( key_b_r_14_16 ) , .Q( key_b_r_15_16 ) );
  DFF_X1 key_b_r_reg_15_17 (.CK( clk ) , .D( key_b_r_14_17 ) , .Q( key_b_r_15_17 ) );
  DFF_X1 key_b_r_reg_15_18 (.CK( clk ) , .D( key_b_r_14_18 ) , .Q( key_b_r_15_18 ) );
  DFF_X1 key_b_r_reg_15_19 (.CK( clk ) , .D( key_b_r_14_19 ) , .Q( key_b_r_15_19 ) );
  DFF_X1 key_b_r_reg_15_2 (.CK( clk ) , .D( key_b_r_14_2 ) , .Q( key_b_r_15_2 ) );
  DFF_X1 key_b_r_reg_15_20 (.CK( clk ) , .D( key_b_r_14_20 ) , .Q( key_b_r_15_20 ) );
  DFF_X1 key_b_r_reg_15_21 (.CK( clk ) , .D( key_b_r_14_21 ) , .Q( key_b_r_15_21 ) );
  DFF_X1 key_b_r_reg_15_22 (.CK( clk ) , .D( key_b_r_14_22 ) , .Q( key_b_r_15_22 ) );
  DFF_X1 key_b_r_reg_15_23 (.CK( clk ) , .D( key_b_r_14_23 ) , .Q( key_b_r_15_23 ) );
  DFF_X1 key_b_r_reg_15_24 (.CK( clk ) , .D( key_b_r_14_24 ) , .Q( key_b_r_15_24 ) );
  DFF_X1 key_b_r_reg_15_25 (.CK( clk ) , .D( key_b_r_14_25 ) , .Q( key_b_r_15_25 ) );
  DFF_X1 key_b_r_reg_15_26 (.CK( clk ) , .D( key_b_r_14_26 ) , .Q( key_b_r_15_26 ) );
  DFF_X1 key_b_r_reg_15_27 (.CK( clk ) , .D( key_b_r_14_27 ) , .Q( key_b_r_15_27 ) );
  DFF_X1 key_b_r_reg_15_28 (.CK( clk ) , .D( key_b_r_14_28 ) , .Q( key_b_r_15_28 ) );
  DFF_X1 key_b_r_reg_15_29 (.CK( clk ) , .D( key_b_r_14_29 ) , .Q( key_b_r_15_29 ) );
  DFF_X1 key_b_r_reg_15_3 (.CK( clk ) , .D( key_b_r_14_3 ) , .Q( key_b_r_15_3 ) );
  DFF_X1 key_b_r_reg_15_30 (.CK( clk ) , .D( key_b_r_14_30 ) , .Q( key_b_r_15_30 ) );
  DFF_X1 key_b_r_reg_15_31 (.CK( clk ) , .D( key_b_r_14_31 ) , .Q( key_b_r_15_31 ) );
  DFF_X1 key_b_r_reg_15_32 (.CK( clk ) , .D( key_b_r_14_32 ) , .Q( key_b_r_15_32 ) );
  DFF_X1 key_b_r_reg_15_33 (.CK( clk ) , .D( key_b_r_14_33 ) , .Q( key_b_r_15_33 ) );
  DFF_X1 key_b_r_reg_15_34 (.CK( clk ) , .D( key_b_r_14_34 ) , .Q( key_b_r_15_34 ) );
  DFF_X1 key_b_r_reg_15_35 (.CK( clk ) , .D( key_b_r_14_35 ) , .Q( key_b_r_15_35 ) );
  DFF_X1 key_b_r_reg_15_36 (.CK( clk ) , .D( key_b_r_14_36 ) , .Q( key_b_r_15_36 ) );
  DFF_X1 key_b_r_reg_15_37 (.CK( clk ) , .D( key_b_r_14_37 ) , .Q( key_b_r_15_37 ) );
  DFF_X1 key_b_r_reg_15_38 (.CK( clk ) , .D( key_b_r_14_38 ) , .Q( key_b_r_15_38 ) );
  DFF_X1 key_b_r_reg_15_39 (.CK( clk ) , .D( key_b_r_14_39 ) , .Q( key_b_r_15_39 ) );
  DFF_X1 key_b_r_reg_15_4 (.CK( clk ) , .D( key_b_r_14_4 ) , .Q( key_b_r_15_4 ) );
  DFF_X1 key_b_r_reg_15_40 (.CK( clk ) , .D( key_b_r_14_40 ) , .Q( key_b_r_15_40 ) );
  DFF_X1 key_b_r_reg_15_41 (.CK( clk ) , .D( key_b_r_14_41 ) , .Q( key_b_r_15_41 ) );
  DFF_X1 key_b_r_reg_15_42 (.CK( clk ) , .D( key_b_r_14_42 ) , .Q( key_b_r_15_42 ) );
  DFF_X1 key_b_r_reg_15_43 (.CK( clk ) , .D( key_b_r_14_43 ) , .Q( key_b_r_15_43 ) );
  DFF_X1 key_b_r_reg_15_44 (.CK( clk ) , .D( key_b_r_14_44 ) , .Q( key_b_r_15_44 ) );
  DFF_X1 key_b_r_reg_15_45 (.CK( clk ) , .D( key_b_r_14_45 ) , .Q( key_b_r_15_45 ) );
  DFF_X1 key_b_r_reg_15_46 (.CK( clk ) , .D( key_b_r_14_46 ) , .Q( key_b_r_15_46 ) );
  DFF_X1 key_b_r_reg_15_47 (.CK( clk ) , .D( key_b_r_14_47 ) , .Q( key_b_r_15_47 ) );
  DFF_X1 key_b_r_reg_15_48 (.CK( clk ) , .D( key_b_r_14_48 ) , .Q( key_b_r_15_48 ) );
  DFF_X1 key_b_r_reg_15_49 (.CK( clk ) , .D( key_b_r_14_49 ) , .Q( key_b_r_15_49 ) );
  DFF_X1 key_b_r_reg_15_5 (.CK( clk ) , .D( key_b_r_14_5 ) , .Q( key_b_r_15_5 ) );
  DFF_X1 key_b_r_reg_15_50 (.CK( clk ) , .D( key_b_r_14_50 ) , .Q( key_b_r_15_50 ) );
  DFF_X1 key_b_r_reg_15_51 (.CK( clk ) , .D( key_b_r_14_51 ) , .Q( key_b_r_15_51 ) );
  DFF_X1 key_b_r_reg_15_52 (.CK( clk ) , .D( key_b_r_14_52 ) , .Q( key_b_r_15_52 ) );
  DFF_X1 key_b_r_reg_15_53 (.CK( clk ) , .D( key_b_r_14_53 ) , .Q( key_b_r_15_53 ) );
  DFF_X1 key_b_r_reg_15_54 (.CK( clk ) , .D( key_b_r_14_54 ) , .Q( key_b_r_15_54 ) );
  DFF_X1 key_b_r_reg_15_55 (.CK( clk ) , .D( key_b_r_14_55 ) , .Q( key_b_r_15_55 ) );
  DFF_X1 key_b_r_reg_15_6 (.CK( clk ) , .D( key_b_r_14_6 ) , .Q( key_b_r_15_6 ) );
  DFF_X1 key_b_r_reg_15_7 (.CK( clk ) , .D( key_b_r_14_7 ) , .Q( key_b_r_15_7 ) );
  DFF_X1 key_b_r_reg_15_8 (.CK( clk ) , .D( key_b_r_14_8 ) , .Q( key_b_r_15_8 ) );
  DFF_X1 key_b_r_reg_15_9 (.CK( clk ) , .D( key_b_r_14_9 ) , .Q( key_b_r_15_9 ) );
  DFF_X1 key_b_r_reg_16_0 (.CK( clk ) , .D( key_b_r_15_0 ) , .Q( key_b_r_16_0 ) );
  DFF_X1 key_b_r_reg_16_1 (.CK( clk ) , .D( key_b_r_15_1 ) , .Q( key_b_r_16_1 ) );
  DFF_X1 key_b_r_reg_16_10 (.CK( clk ) , .D( key_b_r_15_10 ) , .Q( key_b_r_16_10 ) );
  DFF_X1 key_b_r_reg_16_11 (.CK( clk ) , .D( key_b_r_15_11 ) , .Q( key_b_r_16_11 ) );
  DFF_X1 key_b_r_reg_16_12 (.CK( clk ) , .D( key_b_r_15_12 ) , .Q( key_b_r_16_12 ) );
  DFF_X1 key_b_r_reg_16_13 (.CK( clk ) , .D( key_b_r_15_13 ) , .Q( key_b_r_16_13 ) );
  DFF_X1 key_b_r_reg_16_14 (.CK( clk ) , .D( key_b_r_15_14 ) , .Q( key_b_r_16_14 ) );
  DFF_X1 key_b_r_reg_16_15 (.CK( clk ) , .D( key_b_r_15_15 ) , .Q( key_b_r_16_15 ) );
  DFF_X1 key_b_r_reg_16_16 (.CK( clk ) , .D( key_b_r_15_16 ) , .Q( key_b_r_16_16 ) );
  DFF_X1 key_b_r_reg_16_17 (.CK( clk ) , .D( key_b_r_15_17 ) , .Q( key_b_r_16_17 ) );
  DFF_X1 key_b_r_reg_16_18 (.CK( clk ) , .D( key_b_r_15_18 ) , .Q( key_b_r_16_18 ) );
  DFF_X1 key_b_r_reg_16_19 (.CK( clk ) , .D( key_b_r_15_19 ) , .Q( key_b_r_16_19 ) );
  DFF_X1 key_b_r_reg_16_2 (.CK( clk ) , .D( key_b_r_15_2 ) , .Q( key_b_r_16_2 ) );
  DFF_X1 key_b_r_reg_16_20 (.CK( clk ) , .D( key_b_r_15_20 ) , .Q( key_b_r_16_20 ) );
  DFF_X1 key_b_r_reg_16_21 (.CK( clk ) , .D( key_b_r_15_21 ) , .Q( key_b_r_16_21 ) );
  DFF_X1 key_b_r_reg_16_22 (.CK( clk ) , .D( key_b_r_15_22 ) , .Q( key_b_r_16_22 ) );
  DFF_X1 key_b_r_reg_16_23 (.CK( clk ) , .D( key_b_r_15_23 ) , .Q( key_b_r_16_23 ) );
  DFF_X1 key_b_r_reg_16_24 (.CK( clk ) , .D( key_b_r_15_24 ) , .Q( key_b_r_16_24 ) );
  DFF_X1 key_b_r_reg_16_25 (.CK( clk ) , .D( key_b_r_15_25 ) , .Q( key_b_r_16_25 ) );
  DFF_X1 key_b_r_reg_16_26 (.CK( clk ) , .D( key_b_r_15_26 ) , .Q( key_b_r_16_26 ) );
  DFF_X1 key_b_r_reg_16_27 (.CK( clk ) , .D( key_b_r_15_27 ) , .Q( key_b_r_16_27 ) );
  DFF_X1 key_b_r_reg_16_28 (.CK( clk ) , .D( key_b_r_15_28 ) , .Q( key_b_r_16_28 ) );
  DFF_X1 key_b_r_reg_16_29 (.CK( clk ) , .D( key_b_r_15_29 ) , .Q( key_b_r_16_29 ) );
  DFF_X1 key_b_r_reg_16_3 (.CK( clk ) , .D( key_b_r_15_3 ) , .Q( key_b_r_16_3 ) );
  DFF_X1 key_b_r_reg_16_30 (.CK( clk ) , .D( key_b_r_15_30 ) , .Q( key_b_r_16_30 ) );
  DFF_X1 key_b_r_reg_16_31 (.CK( clk ) , .D( key_b_r_15_31 ) , .Q( key_b_r_16_31 ) );
  DFF_X1 key_b_r_reg_16_32 (.CK( clk ) , .D( key_b_r_15_32 ) , .Q( key_b_r_16_32 ) );
  DFF_X1 key_b_r_reg_16_33 (.CK( clk ) , .D( key_b_r_15_33 ) , .Q( key_b_r_16_33 ) );
  DFF_X1 key_b_r_reg_16_34 (.CK( clk ) , .D( key_b_r_15_34 ) , .Q( key_b_r_16_34 ) );
  DFF_X1 key_b_r_reg_16_35 (.CK( clk ) , .D( key_b_r_15_35 ) , .Q( key_b_r_16_35 ) );
  DFF_X1 key_b_r_reg_16_36 (.CK( clk ) , .D( key_b_r_15_36 ) , .Q( key_b_r_16_36 ) );
  DFF_X1 key_b_r_reg_16_37 (.CK( clk ) , .D( key_b_r_15_37 ) , .Q( key_b_r_16_37 ) );
  DFF_X1 key_b_r_reg_16_38 (.CK( clk ) , .D( key_b_r_15_38 ) , .Q( key_b_r_16_38 ) );
  DFF_X1 key_b_r_reg_16_39 (.CK( clk ) , .D( key_b_r_15_39 ) , .Q( key_b_r_16_39 ) );
  DFF_X1 key_b_r_reg_16_4 (.CK( clk ) , .D( key_b_r_15_4 ) , .Q( key_b_r_16_4 ) );
  DFF_X1 key_b_r_reg_16_40 (.CK( clk ) , .D( key_b_r_15_40 ) , .Q( key_b_r_16_40 ) );
  DFF_X1 key_b_r_reg_16_41 (.CK( clk ) , .D( key_b_r_15_41 ) , .Q( key_b_r_16_41 ) );
  DFF_X1 key_b_r_reg_16_42 (.CK( clk ) , .D( key_b_r_15_42 ) , .Q( key_b_r_16_42 ) );
  DFF_X1 key_b_r_reg_16_43 (.CK( clk ) , .D( key_b_r_15_43 ) , .Q( key_b_r_16_43 ) );
  DFF_X1 key_b_r_reg_16_44 (.CK( clk ) , .D( key_b_r_15_44 ) , .Q( key_b_r_16_44 ) );
  DFF_X1 key_b_r_reg_16_45 (.CK( clk ) , .D( key_b_r_15_45 ) , .Q( key_b_r_16_45 ) );
  DFF_X1 key_b_r_reg_16_46 (.CK( clk ) , .D( key_b_r_15_46 ) , .Q( key_b_r_16_46 ) );
  DFF_X1 key_b_r_reg_16_47 (.CK( clk ) , .D( key_b_r_15_47 ) , .Q( key_b_r_16_47 ) );
  DFF_X1 key_b_r_reg_16_48 (.CK( clk ) , .D( key_b_r_15_48 ) , .Q( key_b_r_16_48 ) );
  DFF_X1 key_b_r_reg_16_49 (.CK( clk ) , .D( key_b_r_15_49 ) , .Q( key_b_r_16_49 ) );
  DFF_X1 key_b_r_reg_16_5 (.CK( clk ) , .D( key_b_r_15_5 ) , .Q( key_b_r_16_5 ) );
  DFF_X1 key_b_r_reg_16_50 (.CK( clk ) , .D( key_b_r_15_50 ) , .Q( key_b_r_16_50 ) );
  DFF_X1 key_b_r_reg_16_51 (.CK( clk ) , .D( key_b_r_15_51 ) , .Q( key_b_r_16_51 ) );
  DFF_X1 key_b_r_reg_16_52 (.CK( clk ) , .D( key_b_r_15_52 ) , .Q( key_b_r_16_52 ) );
  DFF_X1 key_b_r_reg_16_53 (.CK( clk ) , .D( key_b_r_15_53 ) , .Q( key_b_r_16_53 ) );
  DFF_X1 key_b_r_reg_16_54 (.CK( clk ) , .D( key_b_r_15_54 ) , .Q( key_b_r_16_54 ) );
  DFF_X1 key_b_r_reg_16_55 (.CK( clk ) , .D( key_b_r_15_55 ) , .Q( key_b_r_16_55 ) );
  DFF_X1 key_b_r_reg_16_6 (.CK( clk ) , .D( key_b_r_15_6 ) , .Q( key_b_r_16_6 ) );
  DFF_X1 key_b_r_reg_16_7 (.CK( clk ) , .D( key_b_r_15_7 ) , .Q( key_b_r_16_7 ) );
  DFF_X1 key_b_r_reg_16_8 (.CK( clk ) , .D( key_b_r_15_8 ) , .Q( key_b_r_16_8 ) );
  DFF_X1 key_b_r_reg_16_9 (.CK( clk ) , .D( key_b_r_15_9 ) , .Q( key_b_r_16_9 ) );
  DFF_X1 key_b_r_reg_1_0 (.CK( clk ) , .D( key_b_r_0_0 ) , .Q( key_b_r_1_0 ) );
  DFF_X1 key_b_r_reg_1_1 (.CK( clk ) , .D( key_b_r_0_1 ) , .Q( key_b_r_1_1 ) );
  DFF_X1 key_b_r_reg_1_10 (.CK( clk ) , .D( key_b_r_0_10 ) , .Q( key_b_r_1_10 ) );
  DFF_X1 key_b_r_reg_1_11 (.CK( clk ) , .D( key_b_r_0_11 ) , .Q( key_b_r_1_11 ) );
  DFF_X1 key_b_r_reg_1_12 (.CK( clk ) , .D( key_b_r_0_12 ) , .Q( key_b_r_1_12 ) );
  DFF_X1 key_b_r_reg_1_13 (.CK( clk ) , .D( key_b_r_0_13 ) , .Q( key_b_r_1_13 ) );
  DFF_X1 key_b_r_reg_1_14 (.CK( clk ) , .D( key_b_r_0_14 ) , .Q( key_b_r_1_14 ) );
  DFF_X1 key_b_r_reg_1_15 (.CK( clk ) , .D( key_b_r_0_15 ) , .Q( key_b_r_1_15 ) );
  DFF_X1 key_b_r_reg_1_16 (.CK( clk ) , .D( key_b_r_0_16 ) , .Q( key_b_r_1_16 ) );
  DFF_X1 key_b_r_reg_1_17 (.CK( clk ) , .D( key_b_r_0_17 ) , .Q( key_b_r_1_17 ) );
  DFF_X1 key_b_r_reg_1_18 (.CK( clk ) , .D( key_b_r_0_18 ) , .Q( key_b_r_1_18 ) );
  DFF_X1 key_b_r_reg_1_19 (.CK( clk ) , .D( key_b_r_0_19 ) , .Q( key_b_r_1_19 ) );
  DFF_X1 key_b_r_reg_1_2 (.CK( clk ) , .D( key_b_r_0_2 ) , .Q( key_b_r_1_2 ) );
  DFF_X1 key_b_r_reg_1_20 (.CK( clk ) , .D( key_b_r_0_20 ) , .Q( key_b_r_1_20 ) );
  DFF_X1 key_b_r_reg_1_21 (.CK( clk ) , .D( key_b_r_0_21 ) , .Q( key_b_r_1_21 ) );
  DFF_X1 key_b_r_reg_1_22 (.CK( clk ) , .D( key_b_r_0_22 ) , .Q( key_b_r_1_22 ) );
  DFF_X1 key_b_r_reg_1_23 (.CK( clk ) , .D( key_b_r_0_23 ) , .Q( key_b_r_1_23 ) );
  DFF_X1 key_b_r_reg_1_24 (.CK( clk ) , .D( key_b_r_0_24 ) , .Q( key_b_r_1_24 ) );
  DFF_X1 key_b_r_reg_1_25 (.CK( clk ) , .D( key_b_r_0_25 ) , .Q( key_b_r_1_25 ) );
  DFF_X1 key_b_r_reg_1_26 (.CK( clk ) , .D( key_b_r_0_26 ) , .Q( key_b_r_1_26 ) );
  DFF_X1 key_b_r_reg_1_27 (.CK( clk ) , .D( key_b_r_0_27 ) , .Q( key_b_r_1_27 ) );
  DFF_X1 key_b_r_reg_1_28 (.CK( clk ) , .D( key_b_r_0_28 ) , .Q( key_b_r_1_28 ) );
  DFF_X1 key_b_r_reg_1_29 (.CK( clk ) , .D( key_b_r_0_29 ) , .Q( key_b_r_1_29 ) );
  DFF_X1 key_b_r_reg_1_3 (.CK( clk ) , .D( key_b_r_0_3 ) , .Q( key_b_r_1_3 ) );
  DFF_X1 key_b_r_reg_1_30 (.CK( clk ) , .D( key_b_r_0_30 ) , .Q( key_b_r_1_30 ) );
  DFF_X1 key_b_r_reg_1_31 (.CK( clk ) , .D( key_b_r_0_31 ) , .Q( key_b_r_1_31 ) );
  DFF_X1 key_b_r_reg_1_32 (.CK( clk ) , .D( key_b_r_0_32 ) , .Q( key_b_r_1_32 ) );
  DFF_X1 key_b_r_reg_1_33 (.CK( clk ) , .D( key_b_r_0_33 ) , .Q( key_b_r_1_33 ) );
  DFF_X1 key_b_r_reg_1_34 (.CK( clk ) , .D( key_b_r_0_34 ) , .Q( key_b_r_1_34 ) );
  DFF_X1 key_b_r_reg_1_35 (.CK( clk ) , .D( key_b_r_0_35 ) , .Q( key_b_r_1_35 ) );
  DFF_X1 key_b_r_reg_1_36 (.CK( clk ) , .D( key_b_r_0_36 ) , .Q( key_b_r_1_36 ) );
  DFF_X1 key_b_r_reg_1_37 (.CK( clk ) , .D( key_b_r_0_37 ) , .Q( key_b_r_1_37 ) );
  DFF_X1 key_b_r_reg_1_38 (.CK( clk ) , .D( key_b_r_0_38 ) , .Q( key_b_r_1_38 ) );
  DFF_X1 key_b_r_reg_1_39 (.CK( clk ) , .D( key_b_r_0_39 ) , .Q( key_b_r_1_39 ) );
  DFF_X1 key_b_r_reg_1_4 (.CK( clk ) , .D( key_b_r_0_4 ) , .Q( key_b_r_1_4 ) );
  DFF_X1 key_b_r_reg_1_40 (.CK( clk ) , .D( key_b_r_0_40 ) , .Q( key_b_r_1_40 ) );
  DFF_X1 key_b_r_reg_1_41 (.CK( clk ) , .D( key_b_r_0_41 ) , .Q( key_b_r_1_41 ) );
  DFF_X1 key_b_r_reg_1_42 (.CK( clk ) , .D( key_b_r_0_42 ) , .Q( key_b_r_1_42 ) );
  DFF_X1 key_b_r_reg_1_43 (.CK( clk ) , .D( key_b_r_0_43 ) , .Q( key_b_r_1_43 ) );
  DFF_X1 key_b_r_reg_1_44 (.CK( clk ) , .D( key_b_r_0_44 ) , .Q( key_b_r_1_44 ) );
  DFF_X1 key_b_r_reg_1_45 (.CK( clk ) , .D( key_b_r_0_45 ) , .Q( key_b_r_1_45 ) );
  DFF_X1 key_b_r_reg_1_46 (.CK( clk ) , .D( key_b_r_0_46 ) , .Q( key_b_r_1_46 ) );
  DFF_X1 key_b_r_reg_1_47 (.CK( clk ) , .D( key_b_r_0_47 ) , .Q( key_b_r_1_47 ) );
  DFF_X1 key_b_r_reg_1_48 (.CK( clk ) , .D( key_b_r_0_48 ) , .Q( key_b_r_1_48 ) );
  DFF_X1 key_b_r_reg_1_49 (.CK( clk ) , .D( key_b_r_0_49 ) , .Q( key_b_r_1_49 ) );
  DFF_X1 key_b_r_reg_1_5 (.CK( clk ) , .D( key_b_r_0_5 ) , .Q( key_b_r_1_5 ) );
  DFF_X1 key_b_r_reg_1_50 (.CK( clk ) , .D( key_b_r_0_50 ) , .Q( key_b_r_1_50 ) );
  DFF_X1 key_b_r_reg_1_51 (.CK( clk ) , .D( key_b_r_0_51 ) , .Q( key_b_r_1_51 ) );
  DFF_X1 key_b_r_reg_1_52 (.CK( clk ) , .D( key_b_r_0_52 ) , .Q( key_b_r_1_52 ) );
  DFF_X1 key_b_r_reg_1_53 (.CK( clk ) , .D( key_b_r_0_53 ) , .Q( key_b_r_1_53 ) );
  DFF_X1 key_b_r_reg_1_54 (.CK( clk ) , .D( key_b_r_0_54 ) , .Q( key_b_r_1_54 ) );
  DFF_X1 key_b_r_reg_1_55 (.CK( clk ) , .D( key_b_r_0_55 ) , .Q( key_b_r_1_55 ) );
  DFF_X1 key_b_r_reg_1_6 (.CK( clk ) , .D( key_b_r_0_6 ) , .Q( key_b_r_1_6 ) );
  DFF_X1 key_b_r_reg_1_7 (.CK( clk ) , .D( key_b_r_0_7 ) , .Q( key_b_r_1_7 ) );
  DFF_X1 key_b_r_reg_1_8 (.CK( clk ) , .D( key_b_r_0_8 ) , .Q( key_b_r_1_8 ) );
  DFF_X1 key_b_r_reg_1_9 (.CK( clk ) , .D( key_b_r_0_9 ) , .Q( key_b_r_1_9 ) );
  DFF_X1 key_b_r_reg_2_0 (.CK( clk ) , .D( key_b_r_1_0 ) , .Q( key_b_r_2_0 ) );
  DFF_X1 key_b_r_reg_2_1 (.CK( clk ) , .D( key_b_r_1_1 ) , .Q( key_b_r_2_1 ) );
  DFF_X1 key_b_r_reg_2_10 (.CK( clk ) , .D( key_b_r_1_10 ) , .Q( key_b_r_2_10 ) );
  DFF_X1 key_b_r_reg_2_11 (.CK( clk ) , .D( key_b_r_1_11 ) , .Q( key_b_r_2_11 ) );
  DFF_X1 key_b_r_reg_2_12 (.CK( clk ) , .D( key_b_r_1_12 ) , .Q( key_b_r_2_12 ) );
  DFF_X1 key_b_r_reg_2_13 (.CK( clk ) , .D( key_b_r_1_13 ) , .Q( key_b_r_2_13 ) );
  DFF_X1 key_b_r_reg_2_14 (.CK( clk ) , .D( key_b_r_1_14 ) , .Q( key_b_r_2_14 ) );
  DFF_X1 key_b_r_reg_2_15 (.CK( clk ) , .D( key_b_r_1_15 ) , .Q( key_b_r_2_15 ) );
  DFF_X1 key_b_r_reg_2_16 (.CK( clk ) , .D( key_b_r_1_16 ) , .Q( key_b_r_2_16 ) );
  DFF_X1 key_b_r_reg_2_17 (.CK( clk ) , .D( key_b_r_1_17 ) , .Q( key_b_r_2_17 ) );
  DFF_X1 key_b_r_reg_2_18 (.CK( clk ) , .D( key_b_r_1_18 ) , .Q( key_b_r_2_18 ) );
  DFF_X1 key_b_r_reg_2_19 (.CK( clk ) , .D( key_b_r_1_19 ) , .Q( key_b_r_2_19 ) );
  DFF_X1 key_b_r_reg_2_2 (.CK( clk ) , .D( key_b_r_1_2 ) , .Q( key_b_r_2_2 ) );
  DFF_X1 key_b_r_reg_2_20 (.CK( clk ) , .D( key_b_r_1_20 ) , .Q( key_b_r_2_20 ) );
  DFF_X1 key_b_r_reg_2_21 (.CK( clk ) , .D( key_b_r_1_21 ) , .Q( key_b_r_2_21 ) );
  DFF_X1 key_b_r_reg_2_22 (.CK( clk ) , .D( key_b_r_1_22 ) , .Q( key_b_r_2_22 ) );
  DFF_X1 key_b_r_reg_2_23 (.CK( clk ) , .D( key_b_r_1_23 ) , .Q( key_b_r_2_23 ) );
  DFF_X1 key_b_r_reg_2_24 (.CK( clk ) , .D( key_b_r_1_24 ) , .Q( key_b_r_2_24 ) );
  DFF_X1 key_b_r_reg_2_25 (.CK( clk ) , .D( key_b_r_1_25 ) , .Q( key_b_r_2_25 ) );
  DFF_X1 key_b_r_reg_2_26 (.CK( clk ) , .D( key_b_r_1_26 ) , .Q( key_b_r_2_26 ) );
  DFF_X1 key_b_r_reg_2_27 (.CK( clk ) , .D( key_b_r_1_27 ) , .Q( key_b_r_2_27 ) );
  DFF_X1 key_b_r_reg_2_28 (.CK( clk ) , .D( key_b_r_1_28 ) , .Q( key_b_r_2_28 ) );
  DFF_X1 key_b_r_reg_2_29 (.CK( clk ) , .D( key_b_r_1_29 ) , .Q( key_b_r_2_29 ) );
  DFF_X1 key_b_r_reg_2_3 (.CK( clk ) , .D( key_b_r_1_3 ) , .Q( key_b_r_2_3 ) );
  DFF_X1 key_b_r_reg_2_30 (.CK( clk ) , .D( key_b_r_1_30 ) , .Q( key_b_r_2_30 ) );
  DFF_X1 key_b_r_reg_2_31 (.CK( clk ) , .D( key_b_r_1_31 ) , .Q( key_b_r_2_31 ) );
  DFF_X1 key_b_r_reg_2_32 (.CK( clk ) , .D( key_b_r_1_32 ) , .Q( key_b_r_2_32 ) );
  DFF_X1 key_b_r_reg_2_33 (.CK( clk ) , .D( key_b_r_1_33 ) , .Q( key_b_r_2_33 ) );
  DFF_X1 key_b_r_reg_2_34 (.CK( clk ) , .D( key_b_r_1_34 ) , .Q( key_b_r_2_34 ) );
  DFF_X1 key_b_r_reg_2_35 (.CK( clk ) , .D( key_b_r_1_35 ) , .Q( key_b_r_2_35 ) );
  DFF_X1 key_b_r_reg_2_36 (.CK( clk ) , .D( key_b_r_1_36 ) , .Q( key_b_r_2_36 ) );
  DFF_X1 key_b_r_reg_2_37 (.CK( clk ) , .D( key_b_r_1_37 ) , .Q( key_b_r_2_37 ) );
  DFF_X1 key_b_r_reg_2_38 (.CK( clk ) , .D( key_b_r_1_38 ) , .Q( key_b_r_2_38 ) );
  DFF_X1 key_b_r_reg_2_39 (.CK( clk ) , .D( key_b_r_1_39 ) , .Q( key_b_r_2_39 ) );
  DFF_X1 key_b_r_reg_2_4 (.CK( clk ) , .D( key_b_r_1_4 ) , .Q( key_b_r_2_4 ) );
  DFF_X1 key_b_r_reg_2_40 (.CK( clk ) , .D( key_b_r_1_40 ) , .Q( key_b_r_2_40 ) );
  DFF_X1 key_b_r_reg_2_41 (.CK( clk ) , .D( key_b_r_1_41 ) , .Q( key_b_r_2_41 ) );
  DFF_X1 key_b_r_reg_2_42 (.CK( clk ) , .D( key_b_r_1_42 ) , .Q( key_b_r_2_42 ) );
  DFF_X1 key_b_r_reg_2_43 (.CK( clk ) , .D( key_b_r_1_43 ) , .Q( key_b_r_2_43 ) );
  DFF_X1 key_b_r_reg_2_44 (.CK( clk ) , .D( key_b_r_1_44 ) , .Q( key_b_r_2_44 ) );
  DFF_X1 key_b_r_reg_2_45 (.CK( clk ) , .D( key_b_r_1_45 ) , .Q( key_b_r_2_45 ) );
  DFF_X1 key_b_r_reg_2_46 (.CK( clk ) , .D( key_b_r_1_46 ) , .Q( key_b_r_2_46 ) );
  DFF_X1 key_b_r_reg_2_47 (.CK( clk ) , .D( key_b_r_1_47 ) , .Q( key_b_r_2_47 ) );
  DFF_X1 key_b_r_reg_2_48 (.CK( clk ) , .D( key_b_r_1_48 ) , .Q( key_b_r_2_48 ) );
  DFF_X1 key_b_r_reg_2_49 (.CK( clk ) , .D( key_b_r_1_49 ) , .Q( key_b_r_2_49 ) );
  DFF_X1 key_b_r_reg_2_5 (.CK( clk ) , .D( key_b_r_1_5 ) , .Q( key_b_r_2_5 ) );
  DFF_X1 key_b_r_reg_2_50 (.CK( clk ) , .D( key_b_r_1_50 ) , .Q( key_b_r_2_50 ) );
  DFF_X1 key_b_r_reg_2_51 (.CK( clk ) , .D( key_b_r_1_51 ) , .Q( key_b_r_2_51 ) );
  DFF_X1 key_b_r_reg_2_52 (.CK( clk ) , .D( key_b_r_1_52 ) , .Q( key_b_r_2_52 ) );
  DFF_X1 key_b_r_reg_2_53 (.CK( clk ) , .D( key_b_r_1_53 ) , .Q( key_b_r_2_53 ) );
  DFF_X1 key_b_r_reg_2_54 (.CK( clk ) , .D( key_b_r_1_54 ) , .Q( key_b_r_2_54 ) );
  DFF_X1 key_b_r_reg_2_55 (.CK( clk ) , .D( key_b_r_1_55 ) , .Q( key_b_r_2_55 ) );
  DFF_X1 key_b_r_reg_2_6 (.CK( clk ) , .D( key_b_r_1_6 ) , .Q( key_b_r_2_6 ) );
  DFF_X1 key_b_r_reg_2_7 (.CK( clk ) , .D( key_b_r_1_7 ) , .Q( key_b_r_2_7 ) );
  DFF_X1 key_b_r_reg_2_8 (.CK( clk ) , .D( key_b_r_1_8 ) , .Q( key_b_r_2_8 ) );
  DFF_X1 key_b_r_reg_2_9 (.CK( clk ) , .D( key_b_r_1_9 ) , .Q( key_b_r_2_9 ) );
  DFF_X1 key_b_r_reg_3_0 (.CK( clk ) , .D( key_b_r_2_0 ) , .Q( key_b_r_3_0 ) );
  DFF_X1 key_b_r_reg_3_1 (.CK( clk ) , .D( key_b_r_2_1 ) , .Q( key_b_r_3_1 ) );
  DFF_X1 key_b_r_reg_3_10 (.CK( clk ) , .D( key_b_r_2_10 ) , .Q( key_b_r_3_10 ) );
  DFF_X1 key_b_r_reg_3_11 (.CK( clk ) , .D( key_b_r_2_11 ) , .Q( key_b_r_3_11 ) );
  DFF_X1 key_b_r_reg_3_12 (.CK( clk ) , .D( key_b_r_2_12 ) , .Q( key_b_r_3_12 ) );
  DFF_X1 key_b_r_reg_3_13 (.CK( clk ) , .D( key_b_r_2_13 ) , .Q( key_b_r_3_13 ) );
  DFF_X1 key_b_r_reg_3_14 (.CK( clk ) , .D( key_b_r_2_14 ) , .Q( key_b_r_3_14 ) );
  DFF_X1 key_b_r_reg_3_15 (.CK( clk ) , .D( key_b_r_2_15 ) , .Q( key_b_r_3_15 ) );
  DFF_X1 key_b_r_reg_3_16 (.CK( clk ) , .D( key_b_r_2_16 ) , .Q( key_b_r_3_16 ) );
  DFF_X1 key_b_r_reg_3_17 (.CK( clk ) , .D( key_b_r_2_17 ) , .Q( key_b_r_3_17 ) );
  DFF_X1 key_b_r_reg_3_18 (.CK( clk ) , .D( key_b_r_2_18 ) , .Q( key_b_r_3_18 ) );
  DFF_X1 key_b_r_reg_3_19 (.CK( clk ) , .D( key_b_r_2_19 ) , .Q( key_b_r_3_19 ) );
  DFF_X1 key_b_r_reg_3_2 (.CK( clk ) , .D( key_b_r_2_2 ) , .Q( key_b_r_3_2 ) );
  DFF_X1 key_b_r_reg_3_20 (.CK( clk ) , .D( key_b_r_2_20 ) , .Q( key_b_r_3_20 ) );
  DFF_X1 key_b_r_reg_3_21 (.CK( clk ) , .D( key_b_r_2_21 ) , .Q( key_b_r_3_21 ) );
  DFF_X1 key_b_r_reg_3_22 (.CK( clk ) , .D( key_b_r_2_22 ) , .Q( key_b_r_3_22 ) );
  DFF_X1 key_b_r_reg_3_23 (.CK( clk ) , .D( key_b_r_2_23 ) , .Q( key_b_r_3_23 ) );
  DFF_X1 key_b_r_reg_3_24 (.CK( clk ) , .D( key_b_r_2_24 ) , .Q( key_b_r_3_24 ) );
  DFF_X1 key_b_r_reg_3_25 (.CK( clk ) , .D( key_b_r_2_25 ) , .Q( key_b_r_3_25 ) );
  DFF_X1 key_b_r_reg_3_26 (.CK( clk ) , .D( key_b_r_2_26 ) , .Q( key_b_r_3_26 ) );
  DFF_X1 key_b_r_reg_3_27 (.CK( clk ) , .D( key_b_r_2_27 ) , .Q( key_b_r_3_27 ) );
  DFF_X1 key_b_r_reg_3_28 (.CK( clk ) , .D( key_b_r_2_28 ) , .Q( key_b_r_3_28 ) );
  DFF_X1 key_b_r_reg_3_29 (.CK( clk ) , .D( key_b_r_2_29 ) , .Q( key_b_r_3_29 ) );
  DFF_X1 key_b_r_reg_3_3 (.CK( clk ) , .D( key_b_r_2_3 ) , .Q( key_b_r_3_3 ) );
  DFF_X1 key_b_r_reg_3_30 (.CK( clk ) , .D( key_b_r_2_30 ) , .Q( key_b_r_3_30 ) );
  DFF_X1 key_b_r_reg_3_31 (.CK( clk ) , .D( key_b_r_2_31 ) , .Q( key_b_r_3_31 ) );
  DFF_X1 key_b_r_reg_3_32 (.CK( clk ) , .D( key_b_r_2_32 ) , .Q( key_b_r_3_32 ) );
  DFF_X1 key_b_r_reg_3_33 (.CK( clk ) , .D( key_b_r_2_33 ) , .Q( key_b_r_3_33 ) );
  DFF_X1 key_b_r_reg_3_34 (.CK( clk ) , .D( key_b_r_2_34 ) , .Q( key_b_r_3_34 ) );
  DFF_X1 key_b_r_reg_3_35 (.CK( clk ) , .D( key_b_r_2_35 ) , .Q( key_b_r_3_35 ) );
  DFF_X1 key_b_r_reg_3_36 (.CK( clk ) , .D( key_b_r_2_36 ) , .Q( key_b_r_3_36 ) );
  DFF_X1 key_b_r_reg_3_37 (.CK( clk ) , .D( key_b_r_2_37 ) , .Q( key_b_r_3_37 ) );
  DFF_X1 key_b_r_reg_3_38 (.CK( clk ) , .D( key_b_r_2_38 ) , .Q( key_b_r_3_38 ) );
  DFF_X1 key_b_r_reg_3_39 (.CK( clk ) , .D( key_b_r_2_39 ) , .Q( key_b_r_3_39 ) );
  DFF_X1 key_b_r_reg_3_4 (.CK( clk ) , .D( key_b_r_2_4 ) , .Q( key_b_r_3_4 ) );
  DFF_X1 key_b_r_reg_3_40 (.CK( clk ) , .D( key_b_r_2_40 ) , .Q( key_b_r_3_40 ) );
  DFF_X1 key_b_r_reg_3_41 (.CK( clk ) , .D( key_b_r_2_41 ) , .Q( key_b_r_3_41 ) );
  DFF_X1 key_b_r_reg_3_42 (.CK( clk ) , .D( key_b_r_2_42 ) , .Q( key_b_r_3_42 ) );
  DFF_X1 key_b_r_reg_3_43 (.CK( clk ) , .D( key_b_r_2_43 ) , .Q( key_b_r_3_43 ) );
  DFF_X1 key_b_r_reg_3_44 (.CK( clk ) , .D( key_b_r_2_44 ) , .Q( key_b_r_3_44 ) );
  DFF_X1 key_b_r_reg_3_45 (.CK( clk ) , .D( key_b_r_2_45 ) , .Q( key_b_r_3_45 ) );
  DFF_X1 key_b_r_reg_3_46 (.CK( clk ) , .D( key_b_r_2_46 ) , .Q( key_b_r_3_46 ) );
  DFF_X1 key_b_r_reg_3_47 (.CK( clk ) , .D( key_b_r_2_47 ) , .Q( key_b_r_3_47 ) );
  DFF_X1 key_b_r_reg_3_48 (.CK( clk ) , .D( key_b_r_2_48 ) , .Q( key_b_r_3_48 ) );
  DFF_X1 key_b_r_reg_3_49 (.CK( clk ) , .D( key_b_r_2_49 ) , .Q( key_b_r_3_49 ) );
  DFF_X1 key_b_r_reg_3_5 (.CK( clk ) , .D( key_b_r_2_5 ) , .Q( key_b_r_3_5 ) );
  DFF_X1 key_b_r_reg_3_50 (.CK( clk ) , .D( key_b_r_2_50 ) , .Q( key_b_r_3_50 ) );
  DFF_X1 key_b_r_reg_3_51 (.CK( clk ) , .D( key_b_r_2_51 ) , .Q( key_b_r_3_51 ) );
  DFF_X1 key_b_r_reg_3_52 (.CK( clk ) , .D( key_b_r_2_52 ) , .Q( key_b_r_3_52 ) );
  DFF_X1 key_b_r_reg_3_53 (.CK( clk ) , .D( key_b_r_2_53 ) , .Q( key_b_r_3_53 ) );
  DFF_X1 key_b_r_reg_3_54 (.CK( clk ) , .D( key_b_r_2_54 ) , .Q( key_b_r_3_54 ) );
  DFF_X1 key_b_r_reg_3_55 (.CK( clk ) , .D( key_b_r_2_55 ) , .Q( key_b_r_3_55 ) );
  DFF_X1 key_b_r_reg_3_6 (.CK( clk ) , .D( key_b_r_2_6 ) , .Q( key_b_r_3_6 ) );
  DFF_X1 key_b_r_reg_3_7 (.CK( clk ) , .D( key_b_r_2_7 ) , .Q( key_b_r_3_7 ) );
  DFF_X1 key_b_r_reg_3_8 (.CK( clk ) , .D( key_b_r_2_8 ) , .Q( key_b_r_3_8 ) );
  DFF_X1 key_b_r_reg_3_9 (.CK( clk ) , .D( key_b_r_2_9 ) , .Q( key_b_r_3_9 ) );
  DFF_X1 key_b_r_reg_4_0 (.CK( clk ) , .D( key_b_r_3_0 ) , .Q( key_b_r_4_0 ) );
  DFF_X1 key_b_r_reg_4_1 (.CK( clk ) , .D( key_b_r_3_1 ) , .Q( key_b_r_4_1 ) );
  DFF_X1 key_b_r_reg_4_10 (.CK( clk ) , .D( key_b_r_3_10 ) , .Q( key_b_r_4_10 ) );
  DFF_X1 key_b_r_reg_4_11 (.CK( clk ) , .D( key_b_r_3_11 ) , .Q( key_b_r_4_11 ) );
  DFF_X1 key_b_r_reg_4_12 (.CK( clk ) , .D( key_b_r_3_12 ) , .Q( key_b_r_4_12 ) );
  DFF_X1 key_b_r_reg_4_13 (.CK( clk ) , .D( key_b_r_3_13 ) , .Q( key_b_r_4_13 ) );
  DFF_X1 key_b_r_reg_4_14 (.CK( clk ) , .D( key_b_r_3_14 ) , .Q( key_b_r_4_14 ) );
  DFF_X1 key_b_r_reg_4_15 (.CK( clk ) , .D( key_b_r_3_15 ) , .Q( key_b_r_4_15 ) );
  DFF_X1 key_b_r_reg_4_16 (.CK( clk ) , .D( key_b_r_3_16 ) , .Q( key_b_r_4_16 ) );
  DFF_X1 key_b_r_reg_4_17 (.CK( clk ) , .D( key_b_r_3_17 ) , .Q( key_b_r_4_17 ) );
  DFF_X1 key_b_r_reg_4_18 (.CK( clk ) , .D( key_b_r_3_18 ) , .Q( key_b_r_4_18 ) );
  DFF_X1 key_b_r_reg_4_19 (.CK( clk ) , .D( key_b_r_3_19 ) , .Q( key_b_r_4_19 ) );
  DFF_X1 key_b_r_reg_4_2 (.CK( clk ) , .D( key_b_r_3_2 ) , .Q( key_b_r_4_2 ) );
  DFF_X1 key_b_r_reg_4_20 (.CK( clk ) , .D( key_b_r_3_20 ) , .Q( key_b_r_4_20 ) );
  DFF_X1 key_b_r_reg_4_21 (.CK( clk ) , .D( key_b_r_3_21 ) , .Q( key_b_r_4_21 ) );
  DFF_X1 key_b_r_reg_4_22 (.CK( clk ) , .D( key_b_r_3_22 ) , .Q( key_b_r_4_22 ) );
  DFF_X1 key_b_r_reg_4_23 (.CK( clk ) , .D( key_b_r_3_23 ) , .Q( key_b_r_4_23 ) );
  DFF_X1 key_b_r_reg_4_24 (.CK( clk ) , .D( key_b_r_3_24 ) , .Q( key_b_r_4_24 ) );
  DFF_X1 key_b_r_reg_4_25 (.CK( clk ) , .D( key_b_r_3_25 ) , .Q( key_b_r_4_25 ) );
  DFF_X1 key_b_r_reg_4_26 (.CK( clk ) , .D( key_b_r_3_26 ) , .Q( key_b_r_4_26 ) );
  DFF_X1 key_b_r_reg_4_27 (.CK( clk ) , .D( key_b_r_3_27 ) , .Q( key_b_r_4_27 ) );
  DFF_X1 key_b_r_reg_4_28 (.CK( clk ) , .D( key_b_r_3_28 ) , .Q( key_b_r_4_28 ) );
  DFF_X1 key_b_r_reg_4_29 (.CK( clk ) , .D( key_b_r_3_29 ) , .Q( key_b_r_4_29 ) );
  DFF_X1 key_b_r_reg_4_3 (.CK( clk ) , .D( key_b_r_3_3 ) , .Q( key_b_r_4_3 ) );
  DFF_X1 key_b_r_reg_4_30 (.CK( clk ) , .D( key_b_r_3_30 ) , .Q( key_b_r_4_30 ) );
  DFF_X1 key_b_r_reg_4_31 (.CK( clk ) , .D( key_b_r_3_31 ) , .Q( key_b_r_4_31 ) );
  DFF_X1 key_b_r_reg_4_32 (.CK( clk ) , .D( key_b_r_3_32 ) , .Q( key_b_r_4_32 ) );
  DFF_X1 key_b_r_reg_4_33 (.CK( clk ) , .D( key_b_r_3_33 ) , .Q( key_b_r_4_33 ) );
  DFF_X1 key_b_r_reg_4_34 (.CK( clk ) , .D( key_b_r_3_34 ) , .Q( key_b_r_4_34 ) );
  DFF_X1 key_b_r_reg_4_35 (.CK( clk ) , .D( key_b_r_3_35 ) , .Q( key_b_r_4_35 ) );
  DFF_X1 key_b_r_reg_4_36 (.CK( clk ) , .D( key_b_r_3_36 ) , .Q( key_b_r_4_36 ) );
  DFF_X1 key_b_r_reg_4_37 (.CK( clk ) , .D( key_b_r_3_37 ) , .Q( key_b_r_4_37 ) );
  DFF_X1 key_b_r_reg_4_38 (.CK( clk ) , .D( key_b_r_3_38 ) , .Q( key_b_r_4_38 ) );
  DFF_X1 key_b_r_reg_4_39 (.CK( clk ) , .D( key_b_r_3_39 ) , .Q( key_b_r_4_39 ) );
  DFF_X1 key_b_r_reg_4_4 (.CK( clk ) , .D( key_b_r_3_4 ) , .Q( key_b_r_4_4 ) );
  DFF_X1 key_b_r_reg_4_40 (.CK( clk ) , .D( key_b_r_3_40 ) , .Q( key_b_r_4_40 ) );
  DFF_X1 key_b_r_reg_4_41 (.CK( clk ) , .D( key_b_r_3_41 ) , .Q( key_b_r_4_41 ) );
  DFF_X1 key_b_r_reg_4_42 (.CK( clk ) , .D( key_b_r_3_42 ) , .Q( key_b_r_4_42 ) );
  DFF_X1 key_b_r_reg_4_43 (.CK( clk ) , .D( key_b_r_3_43 ) , .Q( key_b_r_4_43 ) );
  DFF_X1 key_b_r_reg_4_44 (.CK( clk ) , .D( key_b_r_3_44 ) , .Q( key_b_r_4_44 ) );
  DFF_X1 key_b_r_reg_4_45 (.CK( clk ) , .D( key_b_r_3_45 ) , .Q( key_b_r_4_45 ) );
  DFF_X1 key_b_r_reg_4_46 (.CK( clk ) , .D( key_b_r_3_46 ) , .Q( key_b_r_4_46 ) );
  DFF_X1 key_b_r_reg_4_47 (.CK( clk ) , .D( key_b_r_3_47 ) , .Q( key_b_r_4_47 ) );
  DFF_X1 key_b_r_reg_4_48 (.CK( clk ) , .D( key_b_r_3_48 ) , .Q( key_b_r_4_48 ) );
  DFF_X1 key_b_r_reg_4_49 (.CK( clk ) , .D( key_b_r_3_49 ) , .Q( key_b_r_4_49 ) );
  DFF_X1 key_b_r_reg_4_5 (.CK( clk ) , .D( key_b_r_3_5 ) , .Q( key_b_r_4_5 ) );
  DFF_X1 key_b_r_reg_4_50 (.CK( clk ) , .D( key_b_r_3_50 ) , .Q( key_b_r_4_50 ) );
  DFF_X1 key_b_r_reg_4_51 (.CK( clk ) , .D( key_b_r_3_51 ) , .Q( key_b_r_4_51 ) );
  DFF_X1 key_b_r_reg_4_52 (.CK( clk ) , .D( key_b_r_3_52 ) , .Q( key_b_r_4_52 ) );
  DFF_X1 key_b_r_reg_4_53 (.CK( clk ) , .D( key_b_r_3_53 ) , .Q( key_b_r_4_53 ) );
  DFF_X1 key_b_r_reg_4_54 (.CK( clk ) , .D( key_b_r_3_54 ) , .Q( key_b_r_4_54 ) );
  DFF_X1 key_b_r_reg_4_55 (.CK( clk ) , .D( key_b_r_3_55 ) , .Q( key_b_r_4_55 ) );
  DFF_X1 key_b_r_reg_4_6 (.CK( clk ) , .D( key_b_r_3_6 ) , .Q( key_b_r_4_6 ) );
  DFF_X1 key_b_r_reg_4_7 (.CK( clk ) , .D( key_b_r_3_7 ) , .Q( key_b_r_4_7 ) );
  DFF_X1 key_b_r_reg_4_8 (.CK( clk ) , .D( key_b_r_3_8 ) , .Q( key_b_r_4_8 ) );
  DFF_X1 key_b_r_reg_4_9 (.CK( clk ) , .D( key_b_r_3_9 ) , .Q( key_b_r_4_9 ) );
  DFF_X1 key_b_r_reg_5_0 (.CK( clk ) , .D( key_b_r_4_0 ) , .Q( key_b_r_5_0 ) );
  DFF_X1 key_b_r_reg_5_1 (.CK( clk ) , .D( key_b_r_4_1 ) , .Q( key_b_r_5_1 ) );
  DFF_X1 key_b_r_reg_5_10 (.CK( clk ) , .D( key_b_r_4_10 ) , .Q( key_b_r_5_10 ) );
  DFF_X1 key_b_r_reg_5_11 (.CK( clk ) , .D( key_b_r_4_11 ) , .Q( key_b_r_5_11 ) );
  DFF_X1 key_b_r_reg_5_12 (.CK( clk ) , .D( key_b_r_4_12 ) , .Q( key_b_r_5_12 ) );
  DFF_X1 key_b_r_reg_5_13 (.CK( clk ) , .D( key_b_r_4_13 ) , .Q( key_b_r_5_13 ) );
  DFF_X1 key_b_r_reg_5_14 (.CK( clk ) , .D( key_b_r_4_14 ) , .Q( key_b_r_5_14 ) );
  DFF_X1 key_b_r_reg_5_15 (.CK( clk ) , .D( key_b_r_4_15 ) , .Q( key_b_r_5_15 ) );
  DFF_X1 key_b_r_reg_5_16 (.CK( clk ) , .D( key_b_r_4_16 ) , .Q( key_b_r_5_16 ) );
  DFF_X1 key_b_r_reg_5_17 (.CK( clk ) , .D( key_b_r_4_17 ) , .Q( key_b_r_5_17 ) );
  DFF_X1 key_b_r_reg_5_18 (.CK( clk ) , .D( key_b_r_4_18 ) , .Q( key_b_r_5_18 ) );
  DFF_X1 key_b_r_reg_5_19 (.CK( clk ) , .D( key_b_r_4_19 ) , .Q( key_b_r_5_19 ) );
  DFF_X1 key_b_r_reg_5_2 (.CK( clk ) , .D( key_b_r_4_2 ) , .Q( key_b_r_5_2 ) );
  DFF_X1 key_b_r_reg_5_20 (.CK( clk ) , .D( key_b_r_4_20 ) , .Q( key_b_r_5_20 ) );
  DFF_X1 key_b_r_reg_5_21 (.CK( clk ) , .D( key_b_r_4_21 ) , .Q( key_b_r_5_21 ) );
  DFF_X1 key_b_r_reg_5_22 (.CK( clk ) , .D( key_b_r_4_22 ) , .Q( key_b_r_5_22 ) );
  DFF_X1 key_b_r_reg_5_23 (.CK( clk ) , .D( key_b_r_4_23 ) , .Q( key_b_r_5_23 ) );
  DFF_X1 key_b_r_reg_5_24 (.CK( clk ) , .D( key_b_r_4_24 ) , .Q( key_b_r_5_24 ) );
  DFF_X1 key_b_r_reg_5_25 (.CK( clk ) , .D( key_b_r_4_25 ) , .Q( key_b_r_5_25 ) );
  DFF_X1 key_b_r_reg_5_26 (.CK( clk ) , .D( key_b_r_4_26 ) , .Q( key_b_r_5_26 ) );
  DFF_X1 key_b_r_reg_5_27 (.CK( clk ) , .D( key_b_r_4_27 ) , .Q( key_b_r_5_27 ) );
  DFF_X1 key_b_r_reg_5_28 (.CK( clk ) , .D( key_b_r_4_28 ) , .Q( key_b_r_5_28 ) );
  DFF_X1 key_b_r_reg_5_29 (.CK( clk ) , .D( key_b_r_4_29 ) , .Q( key_b_r_5_29 ) );
  DFF_X1 key_b_r_reg_5_3 (.CK( clk ) , .D( key_b_r_4_3 ) , .Q( key_b_r_5_3 ) );
  DFF_X1 key_b_r_reg_5_30 (.CK( clk ) , .D( key_b_r_4_30 ) , .Q( key_b_r_5_30 ) );
  DFF_X1 key_b_r_reg_5_31 (.CK( clk ) , .D( key_b_r_4_31 ) , .Q( key_b_r_5_31 ) );
  DFF_X1 key_b_r_reg_5_32 (.CK( clk ) , .D( key_b_r_4_32 ) , .Q( key_b_r_5_32 ) );
  DFF_X1 key_b_r_reg_5_33 (.CK( clk ) , .D( key_b_r_4_33 ) , .Q( key_b_r_5_33 ) );
  DFF_X1 key_b_r_reg_5_34 (.CK( clk ) , .D( key_b_r_4_34 ) , .Q( key_b_r_5_34 ) );
  DFF_X1 key_b_r_reg_5_35 (.CK( clk ) , .D( key_b_r_4_35 ) , .Q( key_b_r_5_35 ) );
  DFF_X1 key_b_r_reg_5_36 (.CK( clk ) , .D( key_b_r_4_36 ) , .Q( key_b_r_5_36 ) );
  DFF_X1 key_b_r_reg_5_37 (.CK( clk ) , .D( key_b_r_4_37 ) , .Q( key_b_r_5_37 ) );
  DFF_X1 key_b_r_reg_5_38 (.CK( clk ) , .D( key_b_r_4_38 ) , .Q( key_b_r_5_38 ) );
  DFF_X1 key_b_r_reg_5_39 (.CK( clk ) , .D( key_b_r_4_39 ) , .Q( key_b_r_5_39 ) );
  DFF_X1 key_b_r_reg_5_4 (.CK( clk ) , .D( key_b_r_4_4 ) , .Q( key_b_r_5_4 ) );
  DFF_X1 key_b_r_reg_5_40 (.CK( clk ) , .D( key_b_r_4_40 ) , .Q( key_b_r_5_40 ) );
  DFF_X1 key_b_r_reg_5_41 (.CK( clk ) , .D( key_b_r_4_41 ) , .Q( key_b_r_5_41 ) );
  DFF_X1 key_b_r_reg_5_42 (.CK( clk ) , .D( key_b_r_4_42 ) , .Q( key_b_r_5_42 ) );
  DFF_X1 key_b_r_reg_5_43 (.CK( clk ) , .D( key_b_r_4_43 ) , .Q( key_b_r_5_43 ) );
  DFF_X1 key_b_r_reg_5_44 (.CK( clk ) , .D( key_b_r_4_44 ) , .Q( key_b_r_5_44 ) );
  DFF_X1 key_b_r_reg_5_45 (.CK( clk ) , .D( key_b_r_4_45 ) , .Q( key_b_r_5_45 ) );
  DFF_X1 key_b_r_reg_5_46 (.CK( clk ) , .D( key_b_r_4_46 ) , .Q( key_b_r_5_46 ) );
  DFF_X1 key_b_r_reg_5_47 (.CK( clk ) , .D( key_b_r_4_47 ) , .Q( key_b_r_5_47 ) );
  DFF_X1 key_b_r_reg_5_48 (.CK( clk ) , .D( key_b_r_4_48 ) , .Q( key_b_r_5_48 ) );
  DFF_X1 key_b_r_reg_5_49 (.CK( clk ) , .D( key_b_r_4_49 ) , .Q( key_b_r_5_49 ) );
  DFF_X1 key_b_r_reg_5_5 (.CK( clk ) , .D( key_b_r_4_5 ) , .Q( key_b_r_5_5 ) );
  DFF_X1 key_b_r_reg_5_50 (.CK( clk ) , .D( key_b_r_4_50 ) , .Q( key_b_r_5_50 ) );
  DFF_X1 key_b_r_reg_5_51 (.CK( clk ) , .D( key_b_r_4_51 ) , .Q( key_b_r_5_51 ) );
  DFF_X1 key_b_r_reg_5_52 (.CK( clk ) , .D( key_b_r_4_52 ) , .Q( key_b_r_5_52 ) );
  DFF_X1 key_b_r_reg_5_53 (.CK( clk ) , .D( key_b_r_4_53 ) , .Q( key_b_r_5_53 ) );
  DFF_X1 key_b_r_reg_5_54 (.CK( clk ) , .D( key_b_r_4_54 ) , .Q( key_b_r_5_54 ) );
  DFF_X1 key_b_r_reg_5_55 (.CK( clk ) , .D( key_b_r_4_55 ) , .Q( key_b_r_5_55 ) );
  DFF_X1 key_b_r_reg_5_6 (.CK( clk ) , .D( key_b_r_4_6 ) , .Q( key_b_r_5_6 ) );
  DFF_X1 key_b_r_reg_5_7 (.CK( clk ) , .D( key_b_r_4_7 ) , .Q( key_b_r_5_7 ) );
  DFF_X1 key_b_r_reg_5_8 (.CK( clk ) , .D( key_b_r_4_8 ) , .Q( key_b_r_5_8 ) );
  DFF_X1 key_b_r_reg_5_9 (.CK( clk ) , .D( key_b_r_4_9 ) , .Q( key_b_r_5_9 ) );
  DFF_X1 key_b_r_reg_6_0 (.CK( clk ) , .D( key_b_r_5_0 ) , .Q( key_b_r_6_0 ) );
  DFF_X1 key_b_r_reg_6_1 (.CK( clk ) , .D( key_b_r_5_1 ) , .Q( key_b_r_6_1 ) );
  DFF_X1 key_b_r_reg_6_10 (.CK( clk ) , .D( key_b_r_5_10 ) , .Q( key_b_r_6_10 ) );
  DFF_X1 key_b_r_reg_6_11 (.CK( clk ) , .D( key_b_r_5_11 ) , .Q( key_b_r_6_11 ) );
  DFF_X1 key_b_r_reg_6_12 (.CK( clk ) , .D( key_b_r_5_12 ) , .Q( key_b_r_6_12 ) );
  DFF_X1 key_b_r_reg_6_13 (.CK( clk ) , .D( key_b_r_5_13 ) , .Q( key_b_r_6_13 ) );
  DFF_X1 key_b_r_reg_6_14 (.CK( clk ) , .D( key_b_r_5_14 ) , .Q( key_b_r_6_14 ) );
  DFF_X1 key_b_r_reg_6_15 (.CK( clk ) , .D( key_b_r_5_15 ) , .Q( key_b_r_6_15 ) );
  DFF_X1 key_b_r_reg_6_16 (.CK( clk ) , .D( key_b_r_5_16 ) , .Q( key_b_r_6_16 ) );
  DFF_X1 key_b_r_reg_6_17 (.CK( clk ) , .D( key_b_r_5_17 ) , .Q( key_b_r_6_17 ) );
  DFF_X1 key_b_r_reg_6_18 (.CK( clk ) , .D( key_b_r_5_18 ) , .Q( key_b_r_6_18 ) );
  DFF_X1 key_b_r_reg_6_19 (.CK( clk ) , .D( key_b_r_5_19 ) , .Q( key_b_r_6_19 ) );
  DFF_X1 key_b_r_reg_6_2 (.CK( clk ) , .D( key_b_r_5_2 ) , .Q( key_b_r_6_2 ) );
  DFF_X1 key_b_r_reg_6_20 (.CK( clk ) , .D( key_b_r_5_20 ) , .Q( key_b_r_6_20 ) );
  DFF_X1 key_b_r_reg_6_21 (.CK( clk ) , .D( key_b_r_5_21 ) , .Q( key_b_r_6_21 ) );
  DFF_X1 key_b_r_reg_6_22 (.CK( clk ) , .D( key_b_r_5_22 ) , .Q( key_b_r_6_22 ) );
  DFF_X1 key_b_r_reg_6_23 (.CK( clk ) , .D( key_b_r_5_23 ) , .Q( key_b_r_6_23 ) );
  DFF_X1 key_b_r_reg_6_24 (.CK( clk ) , .D( key_b_r_5_24 ) , .Q( key_b_r_6_24 ) );
  DFF_X1 key_b_r_reg_6_25 (.CK( clk ) , .D( key_b_r_5_25 ) , .Q( key_b_r_6_25 ) );
  DFF_X1 key_b_r_reg_6_26 (.CK( clk ) , .D( key_b_r_5_26 ) , .Q( key_b_r_6_26 ) );
  DFF_X1 key_b_r_reg_6_27 (.CK( clk ) , .D( key_b_r_5_27 ) , .Q( key_b_r_6_27 ) );
  DFF_X1 key_b_r_reg_6_28 (.CK( clk ) , .D( key_b_r_5_28 ) , .Q( key_b_r_6_28 ) );
  DFF_X1 key_b_r_reg_6_29 (.CK( clk ) , .D( key_b_r_5_29 ) , .Q( key_b_r_6_29 ) );
  DFF_X1 key_b_r_reg_6_3 (.CK( clk ) , .D( key_b_r_5_3 ) , .Q( key_b_r_6_3 ) );
  DFF_X1 key_b_r_reg_6_30 (.CK( clk ) , .D( key_b_r_5_30 ) , .Q( key_b_r_6_30 ) );
  DFF_X1 key_b_r_reg_6_31 (.CK( clk ) , .D( key_b_r_5_31 ) , .Q( key_b_r_6_31 ) );
  DFF_X1 key_b_r_reg_6_32 (.CK( clk ) , .D( key_b_r_5_32 ) , .Q( key_b_r_6_32 ) );
  DFF_X1 key_b_r_reg_6_33 (.CK( clk ) , .D( key_b_r_5_33 ) , .Q( key_b_r_6_33 ) );
  DFF_X1 key_b_r_reg_6_34 (.CK( clk ) , .D( key_b_r_5_34 ) , .Q( key_b_r_6_34 ) );
  DFF_X1 key_b_r_reg_6_35 (.CK( clk ) , .D( key_b_r_5_35 ) , .Q( key_b_r_6_35 ) );
  DFF_X1 key_b_r_reg_6_36 (.CK( clk ) , .D( key_b_r_5_36 ) , .Q( key_b_r_6_36 ) );
  DFF_X1 key_b_r_reg_6_37 (.CK( clk ) , .D( key_b_r_5_37 ) , .Q( key_b_r_6_37 ) );
  DFF_X1 key_b_r_reg_6_38 (.CK( clk ) , .D( key_b_r_5_38 ) , .Q( key_b_r_6_38 ) );
  DFF_X1 key_b_r_reg_6_39 (.CK( clk ) , .D( key_b_r_5_39 ) , .Q( key_b_r_6_39 ) );
  DFF_X1 key_b_r_reg_6_4 (.CK( clk ) , .D( key_b_r_5_4 ) , .Q( key_b_r_6_4 ) );
  DFF_X1 key_b_r_reg_6_40 (.CK( clk ) , .D( key_b_r_5_40 ) , .Q( key_b_r_6_40 ) );
  DFF_X1 key_b_r_reg_6_41 (.CK( clk ) , .D( key_b_r_5_41 ) , .Q( key_b_r_6_41 ) );
  DFF_X1 key_b_r_reg_6_42 (.CK( clk ) , .D( key_b_r_5_42 ) , .Q( key_b_r_6_42 ) );
  DFF_X1 key_b_r_reg_6_43 (.CK( clk ) , .D( key_b_r_5_43 ) , .Q( key_b_r_6_43 ) );
  DFF_X1 key_b_r_reg_6_44 (.CK( clk ) , .D( key_b_r_5_44 ) , .Q( key_b_r_6_44 ) );
  DFF_X1 key_b_r_reg_6_45 (.CK( clk ) , .D( key_b_r_5_45 ) , .Q( key_b_r_6_45 ) );
  DFF_X1 key_b_r_reg_6_46 (.CK( clk ) , .D( key_b_r_5_46 ) , .Q( key_b_r_6_46 ) );
  DFF_X1 key_b_r_reg_6_47 (.CK( clk ) , .D( key_b_r_5_47 ) , .Q( key_b_r_6_47 ) );
  DFF_X1 key_b_r_reg_6_48 (.CK( clk ) , .D( key_b_r_5_48 ) , .Q( key_b_r_6_48 ) );
  DFF_X1 key_b_r_reg_6_49 (.CK( clk ) , .D( key_b_r_5_49 ) , .Q( key_b_r_6_49 ) );
  DFF_X1 key_b_r_reg_6_5 (.CK( clk ) , .D( key_b_r_5_5 ) , .Q( key_b_r_6_5 ) );
  DFF_X1 key_b_r_reg_6_50 (.CK( clk ) , .D( key_b_r_5_50 ) , .Q( key_b_r_6_50 ) );
  DFF_X1 key_b_r_reg_6_51 (.CK( clk ) , .D( key_b_r_5_51 ) , .Q( key_b_r_6_51 ) );
  DFF_X1 key_b_r_reg_6_52 (.CK( clk ) , .D( key_b_r_5_52 ) , .Q( key_b_r_6_52 ) );
  DFF_X1 key_b_r_reg_6_53 (.CK( clk ) , .D( key_b_r_5_53 ) , .Q( key_b_r_6_53 ) );
  DFF_X1 key_b_r_reg_6_54 (.CK( clk ) , .D( key_b_r_5_54 ) , .Q( key_b_r_6_54 ) );
  DFF_X1 key_b_r_reg_6_55 (.CK( clk ) , .D( key_b_r_5_55 ) , .Q( key_b_r_6_55 ) );
  DFF_X1 key_b_r_reg_6_6 (.CK( clk ) , .D( key_b_r_5_6 ) , .Q( key_b_r_6_6 ) );
  DFF_X1 key_b_r_reg_6_7 (.CK( clk ) , .D( key_b_r_5_7 ) , .Q( key_b_r_6_7 ) );
  DFF_X1 key_b_r_reg_6_8 (.CK( clk ) , .D( key_b_r_5_8 ) , .Q( key_b_r_6_8 ) );
  DFF_X1 key_b_r_reg_6_9 (.CK( clk ) , .D( key_b_r_5_9 ) , .Q( key_b_r_6_9 ) );
  DFF_X1 key_b_r_reg_7_0 (.CK( clk ) , .D( key_b_r_6_0 ) , .Q( key_b_r_7_0 ) );
  DFF_X1 key_b_r_reg_7_1 (.CK( clk ) , .D( key_b_r_6_1 ) , .Q( key_b_r_7_1 ) );
  DFF_X1 key_b_r_reg_7_10 (.CK( clk ) , .D( key_b_r_6_10 ) , .Q( key_b_r_7_10 ) );
  DFF_X1 key_b_r_reg_7_11 (.CK( clk ) , .D( key_b_r_6_11 ) , .Q( key_b_r_7_11 ) );
  DFF_X1 key_b_r_reg_7_12 (.CK( clk ) , .D( key_b_r_6_12 ) , .Q( key_b_r_7_12 ) );
  DFF_X1 key_b_r_reg_7_13 (.CK( clk ) , .D( key_b_r_6_13 ) , .Q( key_b_r_7_13 ) );
  DFF_X1 key_b_r_reg_7_14 (.CK( clk ) , .D( key_b_r_6_14 ) , .Q( key_b_r_7_14 ) );
  DFF_X1 key_b_r_reg_7_15 (.CK( clk ) , .D( key_b_r_6_15 ) , .Q( key_b_r_7_15 ) );
  DFF_X1 key_b_r_reg_7_16 (.CK( clk ) , .D( key_b_r_6_16 ) , .Q( key_b_r_7_16 ) );
  DFF_X1 key_b_r_reg_7_17 (.CK( clk ) , .D( key_b_r_6_17 ) , .Q( key_b_r_7_17 ) );
  DFF_X1 key_b_r_reg_7_18 (.CK( clk ) , .D( key_b_r_6_18 ) , .Q( key_b_r_7_18 ) );
  DFF_X1 key_b_r_reg_7_19 (.CK( clk ) , .D( key_b_r_6_19 ) , .Q( key_b_r_7_19 ) );
  DFF_X1 key_b_r_reg_7_2 (.CK( clk ) , .D( key_b_r_6_2 ) , .Q( key_b_r_7_2 ) );
  DFF_X1 key_b_r_reg_7_20 (.CK( clk ) , .D( key_b_r_6_20 ) , .Q( key_b_r_7_20 ) );
  DFF_X1 key_b_r_reg_7_21 (.CK( clk ) , .D( key_b_r_6_21 ) , .Q( key_b_r_7_21 ) );
  DFF_X1 key_b_r_reg_7_22 (.CK( clk ) , .D( key_b_r_6_22 ) , .Q( key_b_r_7_22 ) );
  DFF_X1 key_b_r_reg_7_23 (.CK( clk ) , .D( key_b_r_6_23 ) , .Q( key_b_r_7_23 ) );
  DFF_X1 key_b_r_reg_7_24 (.CK( clk ) , .D( key_b_r_6_24 ) , .Q( key_b_r_7_24 ) );
  DFF_X1 key_b_r_reg_7_25 (.CK( clk ) , .D( key_b_r_6_25 ) , .Q( key_b_r_7_25 ) );
  DFF_X1 key_b_r_reg_7_26 (.CK( clk ) , .D( key_b_r_6_26 ) , .Q( key_b_r_7_26 ) );
  DFF_X1 key_b_r_reg_7_27 (.CK( clk ) , .D( key_b_r_6_27 ) , .Q( key_b_r_7_27 ) );
  DFF_X1 key_b_r_reg_7_28 (.CK( clk ) , .D( key_b_r_6_28 ) , .Q( key_b_r_7_28 ) );
  DFF_X1 key_b_r_reg_7_29 (.CK( clk ) , .D( key_b_r_6_29 ) , .Q( key_b_r_7_29 ) );
  DFF_X1 key_b_r_reg_7_3 (.CK( clk ) , .D( key_b_r_6_3 ) , .Q( key_b_r_7_3 ) );
  DFF_X1 key_b_r_reg_7_30 (.CK( clk ) , .D( key_b_r_6_30 ) , .Q( key_b_r_7_30 ) );
  DFF_X1 key_b_r_reg_7_31 (.CK( clk ) , .D( key_b_r_6_31 ) , .Q( key_b_r_7_31 ) );
  DFF_X1 key_b_r_reg_7_32 (.CK( clk ) , .D( key_b_r_6_32 ) , .Q( key_b_r_7_32 ) );
  DFF_X1 key_b_r_reg_7_33 (.CK( clk ) , .D( key_b_r_6_33 ) , .Q( key_b_r_7_33 ) );
  DFF_X1 key_b_r_reg_7_34 (.CK( clk ) , .D( key_b_r_6_34 ) , .Q( key_b_r_7_34 ) );
  DFF_X1 key_b_r_reg_7_35 (.CK( clk ) , .D( key_b_r_6_35 ) , .Q( key_b_r_7_35 ) );
  DFF_X1 key_b_r_reg_7_36 (.CK( clk ) , .D( key_b_r_6_36 ) , .Q( key_b_r_7_36 ) );
  DFF_X1 key_b_r_reg_7_37 (.CK( clk ) , .D( key_b_r_6_37 ) , .Q( key_b_r_7_37 ) );
  DFF_X1 key_b_r_reg_7_38 (.CK( clk ) , .D( key_b_r_6_38 ) , .Q( key_b_r_7_38 ) );
  DFF_X1 key_b_r_reg_7_39 (.CK( clk ) , .D( key_b_r_6_39 ) , .Q( key_b_r_7_39 ) );
  DFF_X1 key_b_r_reg_7_4 (.CK( clk ) , .D( key_b_r_6_4 ) , .Q( key_b_r_7_4 ) );
  DFF_X1 key_b_r_reg_7_40 (.CK( clk ) , .D( key_b_r_6_40 ) , .Q( key_b_r_7_40 ) );
  DFF_X1 key_b_r_reg_7_41 (.CK( clk ) , .D( key_b_r_6_41 ) , .Q( key_b_r_7_41 ) );
  DFF_X1 key_b_r_reg_7_42 (.CK( clk ) , .D( key_b_r_6_42 ) , .Q( key_b_r_7_42 ) );
  DFF_X1 key_b_r_reg_7_43 (.CK( clk ) , .D( key_b_r_6_43 ) , .Q( key_b_r_7_43 ) );
  DFF_X1 key_b_r_reg_7_44 (.CK( clk ) , .D( key_b_r_6_44 ) , .Q( key_b_r_7_44 ) );
  DFF_X1 key_b_r_reg_7_45 (.CK( clk ) , .D( key_b_r_6_45 ) , .Q( key_b_r_7_45 ) );
  DFF_X1 key_b_r_reg_7_46 (.CK( clk ) , .D( key_b_r_6_46 ) , .Q( key_b_r_7_46 ) );
  DFF_X1 key_b_r_reg_7_47 (.CK( clk ) , .D( key_b_r_6_47 ) , .Q( key_b_r_7_47 ) );
  DFF_X1 key_b_r_reg_7_48 (.CK( clk ) , .D( key_b_r_6_48 ) , .Q( key_b_r_7_48 ) );
  DFF_X1 key_b_r_reg_7_49 (.CK( clk ) , .D( key_b_r_6_49 ) , .Q( key_b_r_7_49 ) );
  DFF_X1 key_b_r_reg_7_5 (.CK( clk ) , .D( key_b_r_6_5 ) , .Q( key_b_r_7_5 ) );
  DFF_X1 key_b_r_reg_7_50 (.CK( clk ) , .D( key_b_r_6_50 ) , .Q( key_b_r_7_50 ) );
  DFF_X1 key_b_r_reg_7_51 (.CK( clk ) , .D( key_b_r_6_51 ) , .Q( key_b_r_7_51 ) );
  DFF_X1 key_b_r_reg_7_52 (.CK( clk ) , .D( key_b_r_6_52 ) , .Q( key_b_r_7_52 ) );
  DFF_X1 key_b_r_reg_7_53 (.CK( clk ) , .D( key_b_r_6_53 ) , .Q( key_b_r_7_53 ) );
  DFF_X1 key_b_r_reg_7_54 (.CK( clk ) , .D( key_b_r_6_54 ) , .Q( key_b_r_7_54 ) );
  DFF_X1 key_b_r_reg_7_55 (.CK( clk ) , .D( key_b_r_6_55 ) , .Q( key_b_r_7_55 ) );
  DFF_X1 key_b_r_reg_7_6 (.CK( clk ) , .D( key_b_r_6_6 ) , .Q( key_b_r_7_6 ) );
  DFF_X1 key_b_r_reg_7_7 (.CK( clk ) , .D( key_b_r_6_7 ) , .Q( key_b_r_7_7 ) );
  DFF_X1 key_b_r_reg_7_8 (.CK( clk ) , .D( key_b_r_6_8 ) , .Q( key_b_r_7_8 ) );
  DFF_X1 key_b_r_reg_7_9 (.CK( clk ) , .D( key_b_r_6_9 ) , .Q( key_b_r_7_9 ) );
  DFF_X1 key_b_r_reg_8_0 (.CK( clk ) , .D( key_b_r_7_0 ) , .Q( key_b_r_8_0 ) );
  DFF_X1 key_b_r_reg_8_1 (.CK( clk ) , .D( key_b_r_7_1 ) , .Q( key_b_r_8_1 ) );
  DFF_X1 key_b_r_reg_8_10 (.CK( clk ) , .D( key_b_r_7_10 ) , .Q( key_b_r_8_10 ) );
  DFF_X1 key_b_r_reg_8_11 (.CK( clk ) , .D( key_b_r_7_11 ) , .Q( key_b_r_8_11 ) );
  DFF_X1 key_b_r_reg_8_12 (.CK( clk ) , .D( key_b_r_7_12 ) , .Q( key_b_r_8_12 ) );
  DFF_X1 key_b_r_reg_8_13 (.CK( clk ) , .D( key_b_r_7_13 ) , .Q( key_b_r_8_13 ) );
  DFF_X1 key_b_r_reg_8_14 (.CK( clk ) , .D( key_b_r_7_14 ) , .Q( key_b_r_8_14 ) );
  DFF_X1 key_b_r_reg_8_15 (.CK( clk ) , .D( key_b_r_7_15 ) , .Q( key_b_r_8_15 ) );
  DFF_X1 key_b_r_reg_8_16 (.CK( clk ) , .D( key_b_r_7_16 ) , .Q( key_b_r_8_16 ) );
  DFF_X1 key_b_r_reg_8_17 (.CK( clk ) , .D( key_b_r_7_17 ) , .Q( key_b_r_8_17 ) );
  DFF_X1 key_b_r_reg_8_18 (.CK( clk ) , .D( key_b_r_7_18 ) , .Q( key_b_r_8_18 ) );
  DFF_X1 key_b_r_reg_8_19 (.CK( clk ) , .D( key_b_r_7_19 ) , .Q( key_b_r_8_19 ) );
  DFF_X1 key_b_r_reg_8_2 (.CK( clk ) , .D( key_b_r_7_2 ) , .Q( key_b_r_8_2 ) );
  DFF_X1 key_b_r_reg_8_20 (.CK( clk ) , .D( key_b_r_7_20 ) , .Q( key_b_r_8_20 ) );
  DFF_X1 key_b_r_reg_8_21 (.CK( clk ) , .D( key_b_r_7_21 ) , .Q( key_b_r_8_21 ) );
  DFF_X1 key_b_r_reg_8_22 (.CK( clk ) , .D( key_b_r_7_22 ) , .Q( key_b_r_8_22 ) );
  DFF_X1 key_b_r_reg_8_23 (.CK( clk ) , .D( key_b_r_7_23 ) , .Q( key_b_r_8_23 ) );
  DFF_X1 key_b_r_reg_8_24 (.CK( clk ) , .D( key_b_r_7_24 ) , .Q( key_b_r_8_24 ) );
  DFF_X1 key_b_r_reg_8_25 (.CK( clk ) , .D( key_b_r_7_25 ) , .Q( key_b_r_8_25 ) );
  DFF_X1 key_b_r_reg_8_26 (.CK( clk ) , .D( key_b_r_7_26 ) , .Q( key_b_r_8_26 ) );
  DFF_X1 key_b_r_reg_8_27 (.CK( clk ) , .D( key_b_r_7_27 ) , .Q( key_b_r_8_27 ) );
  DFF_X1 key_b_r_reg_8_28 (.CK( clk ) , .D( key_b_r_7_28 ) , .Q( key_b_r_8_28 ) );
  DFF_X1 key_b_r_reg_8_29 (.CK( clk ) , .D( key_b_r_7_29 ) , .Q( key_b_r_8_29 ) );
  DFF_X1 key_b_r_reg_8_3 (.CK( clk ) , .D( key_b_r_7_3 ) , .Q( key_b_r_8_3 ) );
  DFF_X1 key_b_r_reg_8_30 (.CK( clk ) , .D( key_b_r_7_30 ) , .Q( key_b_r_8_30 ) );
  DFF_X1 key_b_r_reg_8_31 (.CK( clk ) , .D( key_b_r_7_31 ) , .Q( key_b_r_8_31 ) );
  DFF_X1 key_b_r_reg_8_32 (.CK( clk ) , .D( key_b_r_7_32 ) , .Q( key_b_r_8_32 ) );
  DFF_X1 key_b_r_reg_8_33 (.CK( clk ) , .D( key_b_r_7_33 ) , .Q( key_b_r_8_33 ) );
  DFF_X1 key_b_r_reg_8_34 (.CK( clk ) , .D( key_b_r_7_34 ) , .Q( key_b_r_8_34 ) );
  DFF_X1 key_b_r_reg_8_35 (.CK( clk ) , .D( key_b_r_7_35 ) , .Q( key_b_r_8_35 ) );
  DFF_X1 key_b_r_reg_8_36 (.CK( clk ) , .D( key_b_r_7_36 ) , .Q( key_b_r_8_36 ) );
  DFF_X1 key_b_r_reg_8_37 (.CK( clk ) , .D( key_b_r_7_37 ) , .Q( key_b_r_8_37 ) );
  DFF_X1 key_b_r_reg_8_38 (.CK( clk ) , .D( key_b_r_7_38 ) , .Q( key_b_r_8_38 ) );
  DFF_X1 key_b_r_reg_8_39 (.CK( clk ) , .D( key_b_r_7_39 ) , .Q( key_b_r_8_39 ) );
  DFF_X1 key_b_r_reg_8_4 (.CK( clk ) , .D( key_b_r_7_4 ) , .Q( key_b_r_8_4 ) );
  DFF_X1 key_b_r_reg_8_40 (.CK( clk ) , .D( key_b_r_7_40 ) , .Q( key_b_r_8_40 ) );
  DFF_X1 key_b_r_reg_8_41 (.CK( clk ) , .D( key_b_r_7_41 ) , .Q( key_b_r_8_41 ) );
  DFF_X1 key_b_r_reg_8_42 (.CK( clk ) , .D( key_b_r_7_42 ) , .Q( key_b_r_8_42 ) );
  DFF_X1 key_b_r_reg_8_43 (.CK( clk ) , .D( key_b_r_7_43 ) , .Q( key_b_r_8_43 ) );
  DFF_X1 key_b_r_reg_8_44 (.CK( clk ) , .D( key_b_r_7_44 ) , .Q( key_b_r_8_44 ) );
  DFF_X1 key_b_r_reg_8_45 (.CK( clk ) , .D( key_b_r_7_45 ) , .Q( key_b_r_8_45 ) );
  DFF_X1 key_b_r_reg_8_46 (.CK( clk ) , .D( key_b_r_7_46 ) , .Q( key_b_r_8_46 ) );
  DFF_X1 key_b_r_reg_8_47 (.CK( clk ) , .D( key_b_r_7_47 ) , .Q( key_b_r_8_47 ) );
  DFF_X1 key_b_r_reg_8_48 (.CK( clk ) , .D( key_b_r_7_48 ) , .Q( key_b_r_8_48 ) );
  DFF_X1 key_b_r_reg_8_49 (.CK( clk ) , .D( key_b_r_7_49 ) , .Q( key_b_r_8_49 ) );
  DFF_X1 key_b_r_reg_8_5 (.CK( clk ) , .D( key_b_r_7_5 ) , .Q( key_b_r_8_5 ) );
  DFF_X1 key_b_r_reg_8_50 (.CK( clk ) , .D( key_b_r_7_50 ) , .Q( key_b_r_8_50 ) );
  DFF_X1 key_b_r_reg_8_51 (.CK( clk ) , .D( key_b_r_7_51 ) , .Q( key_b_r_8_51 ) );
  DFF_X1 key_b_r_reg_8_52 (.CK( clk ) , .D( key_b_r_7_52 ) , .Q( key_b_r_8_52 ) );
  DFF_X1 key_b_r_reg_8_53 (.CK( clk ) , .D( key_b_r_7_53 ) , .Q( key_b_r_8_53 ) );
  DFF_X1 key_b_r_reg_8_54 (.CK( clk ) , .D( key_b_r_7_54 ) , .Q( key_b_r_8_54 ) );
  DFF_X1 key_b_r_reg_8_55 (.CK( clk ) , .D( key_b_r_7_55 ) , .Q( key_b_r_8_55 ) );
  DFF_X1 key_b_r_reg_8_6 (.CK( clk ) , .D( key_b_r_7_6 ) , .Q( key_b_r_8_6 ) );
  DFF_X1 key_b_r_reg_8_7 (.CK( clk ) , .D( key_b_r_7_7 ) , .Q( key_b_r_8_7 ) );
  DFF_X1 key_b_r_reg_8_8 (.CK( clk ) , .D( key_b_r_7_8 ) , .Q( key_b_r_8_8 ) );
  DFF_X1 key_b_r_reg_8_9 (.CK( clk ) , .D( key_b_r_7_9 ) , .Q( key_b_r_8_9 ) );
  DFF_X1 key_b_r_reg_9_0 (.CK( clk ) , .D( key_b_r_8_0 ) , .Q( key_b_r_9_0 ) );
  DFF_X1 key_b_r_reg_9_1 (.CK( clk ) , .D( key_b_r_8_1 ) , .Q( key_b_r_9_1 ) );
  DFF_X1 key_b_r_reg_9_10 (.CK( clk ) , .D( key_b_r_8_10 ) , .Q( key_b_r_9_10 ) );
  DFF_X1 key_b_r_reg_9_11 (.CK( clk ) , .D( key_b_r_8_11 ) , .Q( key_b_r_9_11 ) );
  DFF_X1 key_b_r_reg_9_12 (.CK( clk ) , .D( key_b_r_8_12 ) , .Q( key_b_r_9_12 ) );
  DFF_X1 key_b_r_reg_9_13 (.CK( clk ) , .D( key_b_r_8_13 ) , .Q( key_b_r_9_13 ) );
  DFF_X1 key_b_r_reg_9_14 (.CK( clk ) , .D( key_b_r_8_14 ) , .Q( key_b_r_9_14 ) );
  DFF_X1 key_b_r_reg_9_15 (.CK( clk ) , .D( key_b_r_8_15 ) , .Q( key_b_r_9_15 ) );
  DFF_X1 key_b_r_reg_9_16 (.CK( clk ) , .D( key_b_r_8_16 ) , .Q( key_b_r_9_16 ) );
  DFF_X1 key_b_r_reg_9_17 (.CK( clk ) , .D( key_b_r_8_17 ) , .Q( key_b_r_9_17 ) );
  DFF_X1 key_b_r_reg_9_18 (.CK( clk ) , .D( key_b_r_8_18 ) , .Q( key_b_r_9_18 ) );
  DFF_X1 key_b_r_reg_9_19 (.CK( clk ) , .D( key_b_r_8_19 ) , .Q( key_b_r_9_19 ) );
  DFF_X1 key_b_r_reg_9_2 (.CK( clk ) , .D( key_b_r_8_2 ) , .Q( key_b_r_9_2 ) );
  DFF_X1 key_b_r_reg_9_20 (.CK( clk ) , .D( key_b_r_8_20 ) , .Q( key_b_r_9_20 ) );
  DFF_X1 key_b_r_reg_9_21 (.CK( clk ) , .D( key_b_r_8_21 ) , .Q( key_b_r_9_21 ) );
  DFF_X1 key_b_r_reg_9_22 (.CK( clk ) , .D( key_b_r_8_22 ) , .Q( key_b_r_9_22 ) );
  DFF_X1 key_b_r_reg_9_23 (.CK( clk ) , .D( key_b_r_8_23 ) , .Q( key_b_r_9_23 ) );
  DFF_X1 key_b_r_reg_9_24 (.CK( clk ) , .D( key_b_r_8_24 ) , .Q( key_b_r_9_24 ) );
  DFF_X1 key_b_r_reg_9_25 (.CK( clk ) , .D( key_b_r_8_25 ) , .Q( key_b_r_9_25 ) );
  DFF_X1 key_b_r_reg_9_26 (.CK( clk ) , .D( key_b_r_8_26 ) , .Q( key_b_r_9_26 ) );
  DFF_X1 key_b_r_reg_9_27 (.CK( clk ) , .D( key_b_r_8_27 ) , .Q( key_b_r_9_27 ) );
  DFF_X1 key_b_r_reg_9_28 (.CK( clk ) , .D( key_b_r_8_28 ) , .Q( key_b_r_9_28 ) );
  DFF_X1 key_b_r_reg_9_29 (.CK( clk ) , .D( key_b_r_8_29 ) , .Q( key_b_r_9_29 ) );
  DFF_X1 key_b_r_reg_9_3 (.CK( clk ) , .D( key_b_r_8_3 ) , .Q( key_b_r_9_3 ) );
  DFF_X1 key_b_r_reg_9_30 (.CK( clk ) , .D( key_b_r_8_30 ) , .Q( key_b_r_9_30 ) );
  DFF_X1 key_b_r_reg_9_31 (.CK( clk ) , .D( key_b_r_8_31 ) , .Q( key_b_r_9_31 ) );
  DFF_X1 key_b_r_reg_9_32 (.CK( clk ) , .D( key_b_r_8_32 ) , .Q( key_b_r_9_32 ) );
  DFF_X1 key_b_r_reg_9_33 (.CK( clk ) , .D( key_b_r_8_33 ) , .Q( key_b_r_9_33 ) );
  DFF_X1 key_b_r_reg_9_34 (.CK( clk ) , .D( key_b_r_8_34 ) , .Q( key_b_r_9_34 ) );
  DFF_X1 key_b_r_reg_9_35 (.CK( clk ) , .D( key_b_r_8_35 ) , .Q( key_b_r_9_35 ) );
  DFF_X1 key_b_r_reg_9_36 (.CK( clk ) , .D( key_b_r_8_36 ) , .Q( key_b_r_9_36 ) );
  DFF_X1 key_b_r_reg_9_37 (.CK( clk ) , .D( key_b_r_8_37 ) , .Q( key_b_r_9_37 ) );
  DFF_X1 key_b_r_reg_9_38 (.CK( clk ) , .D( key_b_r_8_38 ) , .Q( key_b_r_9_38 ) );
  DFF_X1 key_b_r_reg_9_39 (.CK( clk ) , .D( key_b_r_8_39 ) , .Q( key_b_r_9_39 ) );
  DFF_X1 key_b_r_reg_9_4 (.CK( clk ) , .D( key_b_r_8_4 ) , .Q( key_b_r_9_4 ) );
  DFF_X1 key_b_r_reg_9_40 (.CK( clk ) , .D( key_b_r_8_40 ) , .Q( key_b_r_9_40 ) );
  DFF_X1 key_b_r_reg_9_41 (.CK( clk ) , .D( key_b_r_8_41 ) , .Q( key_b_r_9_41 ) );
  DFF_X1 key_b_r_reg_9_42 (.CK( clk ) , .D( key_b_r_8_42 ) , .Q( key_b_r_9_42 ) );
  DFF_X1 key_b_r_reg_9_43 (.CK( clk ) , .D( key_b_r_8_43 ) , .Q( key_b_r_9_43 ) );
  DFF_X1 key_b_r_reg_9_44 (.CK( clk ) , .D( key_b_r_8_44 ) , .Q( key_b_r_9_44 ) );
  DFF_X1 key_b_r_reg_9_45 (.CK( clk ) , .D( key_b_r_8_45 ) , .Q( key_b_r_9_45 ) );
  DFF_X1 key_b_r_reg_9_46 (.CK( clk ) , .D( key_b_r_8_46 ) , .Q( key_b_r_9_46 ) );
  DFF_X1 key_b_r_reg_9_47 (.CK( clk ) , .D( key_b_r_8_47 ) , .Q( key_b_r_9_47 ) );
  DFF_X1 key_b_r_reg_9_48 (.CK( clk ) , .D( key_b_r_8_48 ) , .Q( key_b_r_9_48 ) );
  DFF_X1 key_b_r_reg_9_49 (.CK( clk ) , .D( key_b_r_8_49 ) , .Q( key_b_r_9_49 ) );
  DFF_X1 key_b_r_reg_9_5 (.CK( clk ) , .D( key_b_r_8_5 ) , .Q( key_b_r_9_5 ) );
  DFF_X1 key_b_r_reg_9_50 (.CK( clk ) , .D( key_b_r_8_50 ) , .Q( key_b_r_9_50 ) );
  DFF_X1 key_b_r_reg_9_51 (.CK( clk ) , .D( key_b_r_8_51 ) , .Q( key_b_r_9_51 ) );
  DFF_X1 key_b_r_reg_9_52 (.CK( clk ) , .D( key_b_r_8_52 ) , .Q( key_b_r_9_52 ) );
  DFF_X1 key_b_r_reg_9_53 (.CK( clk ) , .D( key_b_r_8_53 ) , .Q( key_b_r_9_53 ) );
  DFF_X1 key_b_r_reg_9_54 (.CK( clk ) , .D( key_b_r_8_54 ) , .Q( key_b_r_9_54 ) );
  DFF_X1 key_b_r_reg_9_55 (.CK( clk ) , .D( key_b_r_8_55 ) , .Q( key_b_r_9_55 ) );
  DFF_X1 key_b_r_reg_9_6 (.CK( clk ) , .D( key_b_r_8_6 ) , .Q( key_b_r_9_6 ) );
  DFF_X1 key_b_r_reg_9_7 (.CK( clk ) , .D( key_b_r_8_7 ) , .Q( key_b_r_9_7 ) );
  DFF_X1 key_b_r_reg_9_8 (.CK( clk ) , .D( key_b_r_8_8 ) , .Q( key_b_r_9_8 ) );
  DFF_X1 key_b_r_reg_9_9 (.CK( clk ) , .D( key_b_r_8_9 ) , .Q( key_b_r_9_9 ) );
  SDFF_X1 key_c_r_reg_0_0 (.CK( clk ) , .SE( decrypt ) , .SI( key1[0] ) , .D( key3[0] ) , .Q( key_c_r_0_0 ) );
  SDFF_X1 key_c_r_reg_0_1 (.CK( clk ) , .SE( decrypt ) , .SI( key1[1] ) , .D( key3[1] ) , .Q( key_c_r_0_1 ) );
  SDFF_X1 key_c_r_reg_0_10 (.CK( clk ) , .SE( decrypt ) , .SI( key1[10] ) , .D( key3[10] ) , .Q( key_c_r_0_10 ) );
  SDFF_X1 key_c_r_reg_0_11 (.CK( clk ) , .SE( decrypt ) , .SI( key1[11] ) , .D( key3[11] ) , .Q( key_c_r_0_11 ) );
  SDFF_X1 key_c_r_reg_0_12 (.CK( clk ) , .SE( decrypt ) , .SI( key1[12] ) , .D( key3[12] ) , .Q( key_c_r_0_12 ) );
  SDFF_X1 key_c_r_reg_0_13 (.CK( clk ) , .SE( decrypt ) , .SI( key1[13] ) , .D( key3[13] ) , .Q( key_c_r_0_13 ) );
  SDFF_X1 key_c_r_reg_0_14 (.CK( clk ) , .SE( decrypt ) , .SI( key1[14] ) , .D( key3[14] ) , .Q( key_c_r_0_14 ) );
  SDFF_X1 key_c_r_reg_0_15 (.CK( clk ) , .SE( decrypt ) , .SI( key1[15] ) , .D( key3[15] ) , .Q( key_c_r_0_15 ) );
  SDFF_X1 key_c_r_reg_0_16 (.CK( clk ) , .SE( decrypt ) , .SI( key1[16] ) , .D( key3[16] ) , .Q( key_c_r_0_16 ) );
  SDFF_X1 key_c_r_reg_0_17 (.CK( clk ) , .SE( decrypt ) , .SI( key1[17] ) , .D( key3[17] ) , .Q( key_c_r_0_17 ) );
  SDFF_X1 key_c_r_reg_0_18 (.CK( clk ) , .SE( decrypt ) , .SI( key1[18] ) , .D( key3[18] ) , .Q( key_c_r_0_18 ) );
  SDFF_X1 key_c_r_reg_0_19 (.CK( clk ) , .SE( decrypt ) , .SI( key1[19] ) , .D( key3[19] ) , .Q( key_c_r_0_19 ) );
  SDFF_X1 key_c_r_reg_0_2 (.CK( clk ) , .SE( decrypt ) , .SI( key1[2] ) , .D( key3[2] ) , .Q( key_c_r_0_2 ) );
  SDFF_X1 key_c_r_reg_0_20 (.CK( clk ) , .SE( decrypt ) , .SI( key1[20] ) , .D( key3[20] ) , .Q( key_c_r_0_20 ) );
  SDFF_X1 key_c_r_reg_0_21 (.CK( clk ) , .SE( decrypt ) , .SI( key1[21] ) , .D( key3[21] ) , .Q( key_c_r_0_21 ) );
  SDFF_X1 key_c_r_reg_0_22 (.CK( clk ) , .SE( decrypt ) , .SI( key1[22] ) , .D( key3[22] ) , .Q( key_c_r_0_22 ) );
  SDFF_X1 key_c_r_reg_0_23 (.CK( clk ) , .SE( decrypt ) , .SI( key1[23] ) , .D( key3[23] ) , .Q( key_c_r_0_23 ) );
  SDFF_X1 key_c_r_reg_0_24 (.CK( clk ) , .SE( decrypt ) , .SI( key1[24] ) , .D( key3[24] ) , .Q( key_c_r_0_24 ) );
  SDFF_X1 key_c_r_reg_0_25 (.CK( clk ) , .SE( decrypt ) , .SI( key1[25] ) , .D( key3[25] ) , .Q( key_c_r_0_25 ) );
  SDFF_X1 key_c_r_reg_0_26 (.CK( clk ) , .SE( decrypt ) , .SI( key1[26] ) , .D( key3[26] ) , .Q( key_c_r_0_26 ) );
  SDFF_X1 key_c_r_reg_0_27 (.CK( clk ) , .SE( decrypt ) , .SI( key1[27] ) , .D( key3[27] ) , .Q( key_c_r_0_27 ) );
  SDFF_X1 key_c_r_reg_0_28 (.CK( clk ) , .SE( decrypt ) , .SI( key1[28] ) , .D( key3[28] ) , .Q( key_c_r_0_28 ) );
  SDFF_X1 key_c_r_reg_0_29 (.CK( clk ) , .SE( decrypt ) , .SI( key1[29] ) , .D( key3[29] ) , .Q( key_c_r_0_29 ) );
  SDFF_X1 key_c_r_reg_0_3 (.CK( clk ) , .SE( decrypt ) , .SI( key1[3] ) , .D( key3[3] ) , .Q( key_c_r_0_3 ) );
  SDFF_X1 key_c_r_reg_0_30 (.CK( clk ) , .SE( decrypt ) , .SI( key1[30] ) , .D( key3[30] ) , .Q( key_c_r_0_30 ) );
  SDFF_X1 key_c_r_reg_0_31 (.CK( clk ) , .SE( decrypt ) , .SI( key1[31] ) , .D( key3[31] ) , .Q( key_c_r_0_31 ) );
  SDFF_X1 key_c_r_reg_0_32 (.CK( clk ) , .SE( decrypt ) , .SI( key1[32] ) , .D( key3[32] ) , .Q( key_c_r_0_32 ) );
  SDFF_X1 key_c_r_reg_0_33 (.CK( clk ) , .SE( decrypt ) , .SI( key1[33] ) , .D( key3[33] ) , .Q( key_c_r_0_33 ) );
  SDFF_X1 key_c_r_reg_0_34 (.CK( clk ) , .SE( decrypt ) , .SI( key1[34] ) , .D( key3[34] ) , .Q( key_c_r_0_34 ) );
  SDFF_X1 key_c_r_reg_0_35 (.CK( clk ) , .SE( decrypt ) , .SI( key1[35] ) , .D( key3[35] ) , .Q( key_c_r_0_35 ) );
  SDFF_X1 key_c_r_reg_0_36 (.CK( clk ) , .SE( decrypt ) , .SI( key1[36] ) , .D( key3[36] ) , .Q( key_c_r_0_36 ) );
  SDFF_X1 key_c_r_reg_0_37 (.CK( clk ) , .SE( decrypt ) , .SI( key1[37] ) , .D( key3[37] ) , .Q( key_c_r_0_37 ) );
  SDFF_X1 key_c_r_reg_0_38 (.CK( clk ) , .SE( decrypt ) , .SI( key1[38] ) , .D( key3[38] ) , .Q( key_c_r_0_38 ) );
  SDFF_X1 key_c_r_reg_0_39 (.CK( clk ) , .SE( decrypt ) , .SI( key1[39] ) , .D( key3[39] ) , .Q( key_c_r_0_39 ) );
  SDFF_X1 key_c_r_reg_0_4 (.CK( clk ) , .SE( decrypt ) , .SI( key1[4] ) , .D( key3[4] ) , .Q( key_c_r_0_4 ) );
  SDFF_X1 key_c_r_reg_0_40 (.CK( clk ) , .SE( decrypt ) , .SI( key1[40] ) , .D( key3[40] ) , .Q( key_c_r_0_40 ) );
  SDFF_X1 key_c_r_reg_0_41 (.CK( clk ) , .SE( decrypt ) , .SI( key1[41] ) , .D( key3[41] ) , .Q( key_c_r_0_41 ) );
  SDFF_X1 key_c_r_reg_0_42 (.CK( clk ) , .SE( decrypt ) , .SI( key1[42] ) , .D( key3[42] ) , .Q( key_c_r_0_42 ) );
  SDFF_X1 key_c_r_reg_0_43 (.CK( clk ) , .SE( decrypt ) , .SI( key1[43] ) , .D( key3[43] ) , .Q( key_c_r_0_43 ) );
  SDFF_X1 key_c_r_reg_0_44 (.CK( clk ) , .SE( decrypt ) , .SI( key1[44] ) , .D( key3[44] ) , .Q( key_c_r_0_44 ) );
  SDFF_X1 key_c_r_reg_0_45 (.CK( clk ) , .SE( decrypt ) , .SI( key1[45] ) , .D( key3[45] ) , .Q( key_c_r_0_45 ) );
  SDFF_X1 key_c_r_reg_0_46 (.CK( clk ) , .SE( decrypt ) , .SI( key1[46] ) , .D( key3[46] ) , .Q( key_c_r_0_46 ) );
  SDFF_X1 key_c_r_reg_0_47 (.CK( clk ) , .SE( decrypt ) , .SI( key1[47] ) , .D( key3[47] ) , .Q( key_c_r_0_47 ) );
  SDFF_X1 key_c_r_reg_0_48 (.CK( clk ) , .SE( decrypt ) , .SI( key1[48] ) , .D( key3[48] ) , .Q( key_c_r_0_48 ) );
  SDFF_X1 key_c_r_reg_0_49 (.CK( clk ) , .SE( decrypt ) , .SI( key1[49] ) , .D( key3[49] ) , .Q( key_c_r_0_49 ) );
  SDFF_X1 key_c_r_reg_0_5 (.CK( clk ) , .SE( decrypt ) , .SI( key1[5] ) , .D( key3[5] ) , .Q( key_c_r_0_5 ) );
  SDFF_X1 key_c_r_reg_0_50 (.CK( clk ) , .SE( decrypt ) , .SI( key1[50] ) , .D( key3[50] ) , .Q( key_c_r_0_50 ) );
  SDFF_X1 key_c_r_reg_0_51 (.CK( clk ) , .SE( decrypt ) , .SI( key1[51] ) , .D( key3[51] ) , .Q( key_c_r_0_51 ) );
  SDFF_X1 key_c_r_reg_0_52 (.CK( clk ) , .SE( decrypt ) , .SI( key1[52] ) , .D( key3[52] ) , .Q( key_c_r_0_52 ) );
  SDFF_X1 key_c_r_reg_0_53 (.CK( clk ) , .SE( decrypt ) , .SI( key1[53] ) , .D( key3[53] ) , .Q( key_c_r_0_53 ) );
  SDFF_X1 key_c_r_reg_0_54 (.CK( clk ) , .SE( decrypt ) , .SI( key1[54] ) , .D( key3[54] ) , .Q( key_c_r_0_54 ) );
  SDFF_X1 key_c_r_reg_0_55 (.CK( clk ) , .SE( decrypt ) , .SI( key1[55] ) , .D( key3[55] ) , .Q( key_c_r_0_55 ) );
  SDFF_X1 key_c_r_reg_0_6 (.CK( clk ) , .SE( decrypt ) , .SI( key1[6] ) , .D( key3[6] ) , .Q( key_c_r_0_6 ) );
  SDFF_X1 key_c_r_reg_0_7 (.CK( clk ) , .SE( decrypt ) , .SI( key1[7] ) , .D( key3[7] ) , .Q( key_c_r_0_7 ) );
  SDFF_X1 key_c_r_reg_0_8 (.CK( clk ) , .SE( decrypt ) , .SI( key1[8] ) , .D( key3[8] ) , .Q( key_c_r_0_8 ) );
  SDFF_X1 key_c_r_reg_0_9 (.CK( clk ) , .SE( decrypt ) , .SI( key1[9] ) , .D( key3[9] ) , .Q( key_c_r_0_9 ) );
  DFF_X1 key_c_r_reg_10_0 (.CK( clk ) , .Q( key_c_r_10_0 ) , .D( key_c_r_9_0 ) );
  DFF_X1 key_c_r_reg_10_1 (.CK( clk ) , .Q( key_c_r_10_1 ) , .D( key_c_r_9_1 ) );
  DFF_X1 key_c_r_reg_10_10 (.CK( clk ) , .Q( key_c_r_10_10 ) , .D( key_c_r_9_10 ) );
  DFF_X1 key_c_r_reg_10_11 (.CK( clk ) , .Q( key_c_r_10_11 ) , .D( key_c_r_9_11 ) );
  DFF_X1 key_c_r_reg_10_12 (.CK( clk ) , .Q( key_c_r_10_12 ) , .D( key_c_r_9_12 ) );
  DFF_X1 key_c_r_reg_10_13 (.CK( clk ) , .Q( key_c_r_10_13 ) , .D( key_c_r_9_13 ) );
  DFF_X1 key_c_r_reg_10_14 (.CK( clk ) , .Q( key_c_r_10_14 ) , .D( key_c_r_9_14 ) );
  DFF_X1 key_c_r_reg_10_15 (.CK( clk ) , .Q( key_c_r_10_15 ) , .D( key_c_r_9_15 ) );
  DFF_X1 key_c_r_reg_10_16 (.CK( clk ) , .Q( key_c_r_10_16 ) , .D( key_c_r_9_16 ) );
  DFF_X1 key_c_r_reg_10_17 (.CK( clk ) , .Q( key_c_r_10_17 ) , .D( key_c_r_9_17 ) );
  DFF_X1 key_c_r_reg_10_18 (.CK( clk ) , .Q( key_c_r_10_18 ) , .D( key_c_r_9_18 ) );
  DFF_X1 key_c_r_reg_10_19 (.CK( clk ) , .Q( key_c_r_10_19 ) , .D( key_c_r_9_19 ) );
  DFF_X1 key_c_r_reg_10_2 (.CK( clk ) , .Q( key_c_r_10_2 ) , .D( key_c_r_9_2 ) );
  DFF_X1 key_c_r_reg_10_20 (.CK( clk ) , .Q( key_c_r_10_20 ) , .D( key_c_r_9_20 ) );
  DFF_X1 key_c_r_reg_10_21 (.CK( clk ) , .Q( key_c_r_10_21 ) , .D( key_c_r_9_21 ) );
  DFF_X1 key_c_r_reg_10_22 (.CK( clk ) , .Q( key_c_r_10_22 ) , .D( key_c_r_9_22 ) );
  DFF_X1 key_c_r_reg_10_23 (.CK( clk ) , .Q( key_c_r_10_23 ) , .D( key_c_r_9_23 ) );
  DFF_X1 key_c_r_reg_10_24 (.CK( clk ) , .Q( key_c_r_10_24 ) , .D( key_c_r_9_24 ) );
  DFF_X1 key_c_r_reg_10_25 (.CK( clk ) , .Q( key_c_r_10_25 ) , .D( key_c_r_9_25 ) );
  DFF_X1 key_c_r_reg_10_26 (.CK( clk ) , .Q( key_c_r_10_26 ) , .D( key_c_r_9_26 ) );
  DFF_X1 key_c_r_reg_10_27 (.CK( clk ) , .Q( key_c_r_10_27 ) , .D( key_c_r_9_27 ) );
  DFF_X1 key_c_r_reg_10_28 (.CK( clk ) , .Q( key_c_r_10_28 ) , .D( key_c_r_9_28 ) );
  DFF_X1 key_c_r_reg_10_29 (.CK( clk ) , .Q( key_c_r_10_29 ) , .D( key_c_r_9_29 ) );
  DFF_X1 key_c_r_reg_10_3 (.CK( clk ) , .Q( key_c_r_10_3 ) , .D( key_c_r_9_3 ) );
  DFF_X1 key_c_r_reg_10_30 (.CK( clk ) , .Q( key_c_r_10_30 ) , .D( key_c_r_9_30 ) );
  DFF_X1 key_c_r_reg_10_31 (.CK( clk ) , .Q( key_c_r_10_31 ) , .D( key_c_r_9_31 ) );
  DFF_X1 key_c_r_reg_10_32 (.CK( clk ) , .Q( key_c_r_10_32 ) , .D( key_c_r_9_32 ) );
  DFF_X1 key_c_r_reg_10_33 (.CK( clk ) , .Q( key_c_r_10_33 ) , .D( key_c_r_9_33 ) );
  DFF_X1 key_c_r_reg_10_34 (.CK( clk ) , .Q( key_c_r_10_34 ) , .D( key_c_r_9_34 ) );
  DFF_X1 key_c_r_reg_10_35 (.CK( clk ) , .Q( key_c_r_10_35 ) , .D( key_c_r_9_35 ) );
  DFF_X1 key_c_r_reg_10_36 (.CK( clk ) , .Q( key_c_r_10_36 ) , .D( key_c_r_9_36 ) );
  DFF_X1 key_c_r_reg_10_37 (.CK( clk ) , .Q( key_c_r_10_37 ) , .D( key_c_r_9_37 ) );
  DFF_X1 key_c_r_reg_10_38 (.CK( clk ) , .Q( key_c_r_10_38 ) , .D( key_c_r_9_38 ) );
  DFF_X1 key_c_r_reg_10_39 (.CK( clk ) , .Q( key_c_r_10_39 ) , .D( key_c_r_9_39 ) );
  DFF_X1 key_c_r_reg_10_4 (.CK( clk ) , .Q( key_c_r_10_4 ) , .D( key_c_r_9_4 ) );
  DFF_X1 key_c_r_reg_10_40 (.CK( clk ) , .Q( key_c_r_10_40 ) , .D( key_c_r_9_40 ) );
  DFF_X1 key_c_r_reg_10_41 (.CK( clk ) , .Q( key_c_r_10_41 ) , .D( key_c_r_9_41 ) );
  DFF_X1 key_c_r_reg_10_42 (.CK( clk ) , .Q( key_c_r_10_42 ) , .D( key_c_r_9_42 ) );
  DFF_X1 key_c_r_reg_10_43 (.CK( clk ) , .Q( key_c_r_10_43 ) , .D( key_c_r_9_43 ) );
  DFF_X1 key_c_r_reg_10_44 (.CK( clk ) , .Q( key_c_r_10_44 ) , .D( key_c_r_9_44 ) );
  DFF_X1 key_c_r_reg_10_45 (.CK( clk ) , .Q( key_c_r_10_45 ) , .D( key_c_r_9_45 ) );
  DFF_X1 key_c_r_reg_10_46 (.CK( clk ) , .Q( key_c_r_10_46 ) , .D( key_c_r_9_46 ) );
  DFF_X1 key_c_r_reg_10_47 (.CK( clk ) , .Q( key_c_r_10_47 ) , .D( key_c_r_9_47 ) );
  DFF_X1 key_c_r_reg_10_48 (.CK( clk ) , .Q( key_c_r_10_48 ) , .D( key_c_r_9_48 ) );
  DFF_X1 key_c_r_reg_10_49 (.CK( clk ) , .Q( key_c_r_10_49 ) , .D( key_c_r_9_49 ) );
  DFF_X1 key_c_r_reg_10_5 (.CK( clk ) , .Q( key_c_r_10_5 ) , .D( key_c_r_9_5 ) );
  DFF_X1 key_c_r_reg_10_50 (.CK( clk ) , .Q( key_c_r_10_50 ) , .D( key_c_r_9_50 ) );
  DFF_X1 key_c_r_reg_10_51 (.CK( clk ) , .Q( key_c_r_10_51 ) , .D( key_c_r_9_51 ) );
  DFF_X1 key_c_r_reg_10_52 (.CK( clk ) , .Q( key_c_r_10_52 ) , .D( key_c_r_9_52 ) );
  DFF_X1 key_c_r_reg_10_53 (.CK( clk ) , .Q( key_c_r_10_53 ) , .D( key_c_r_9_53 ) );
  DFF_X1 key_c_r_reg_10_54 (.CK( clk ) , .Q( key_c_r_10_54 ) , .D( key_c_r_9_54 ) );
  DFF_X1 key_c_r_reg_10_55 (.CK( clk ) , .Q( key_c_r_10_55 ) , .D( key_c_r_9_55 ) );
  DFF_X1 key_c_r_reg_10_6 (.CK( clk ) , .Q( key_c_r_10_6 ) , .D( key_c_r_9_6 ) );
  DFF_X1 key_c_r_reg_10_7 (.CK( clk ) , .Q( key_c_r_10_7 ) , .D( key_c_r_9_7 ) );
  DFF_X1 key_c_r_reg_10_8 (.CK( clk ) , .Q( key_c_r_10_8 ) , .D( key_c_r_9_8 ) );
  DFF_X1 key_c_r_reg_10_9 (.CK( clk ) , .Q( key_c_r_10_9 ) , .D( key_c_r_9_9 ) );
  DFF_X1 key_c_r_reg_11_0 (.CK( clk ) , .D( key_c_r_10_0 ) , .Q( key_c_r_11_0 ) );
  DFF_X1 key_c_r_reg_11_1 (.CK( clk ) , .D( key_c_r_10_1 ) , .Q( key_c_r_11_1 ) );
  DFF_X1 key_c_r_reg_11_10 (.CK( clk ) , .D( key_c_r_10_10 ) , .Q( key_c_r_11_10 ) );
  DFF_X1 key_c_r_reg_11_11 (.CK( clk ) , .D( key_c_r_10_11 ) , .Q( key_c_r_11_11 ) );
  DFF_X1 key_c_r_reg_11_12 (.CK( clk ) , .D( key_c_r_10_12 ) , .Q( key_c_r_11_12 ) );
  DFF_X1 key_c_r_reg_11_13 (.CK( clk ) , .D( key_c_r_10_13 ) , .Q( key_c_r_11_13 ) );
  DFF_X1 key_c_r_reg_11_14 (.CK( clk ) , .D( key_c_r_10_14 ) , .Q( key_c_r_11_14 ) );
  DFF_X1 key_c_r_reg_11_15 (.CK( clk ) , .D( key_c_r_10_15 ) , .Q( key_c_r_11_15 ) );
  DFF_X1 key_c_r_reg_11_16 (.CK( clk ) , .D( key_c_r_10_16 ) , .Q( key_c_r_11_16 ) );
  DFF_X1 key_c_r_reg_11_17 (.CK( clk ) , .D( key_c_r_10_17 ) , .Q( key_c_r_11_17 ) );
  DFF_X1 key_c_r_reg_11_18 (.CK( clk ) , .D( key_c_r_10_18 ) , .Q( key_c_r_11_18 ) );
  DFF_X1 key_c_r_reg_11_19 (.CK( clk ) , .D( key_c_r_10_19 ) , .Q( key_c_r_11_19 ) );
  DFF_X1 key_c_r_reg_11_2 (.CK( clk ) , .D( key_c_r_10_2 ) , .Q( key_c_r_11_2 ) );
  DFF_X1 key_c_r_reg_11_20 (.CK( clk ) , .D( key_c_r_10_20 ) , .Q( key_c_r_11_20 ) );
  DFF_X1 key_c_r_reg_11_21 (.CK( clk ) , .D( key_c_r_10_21 ) , .Q( key_c_r_11_21 ) );
  DFF_X1 key_c_r_reg_11_22 (.CK( clk ) , .D( key_c_r_10_22 ) , .Q( key_c_r_11_22 ) );
  DFF_X1 key_c_r_reg_11_23 (.CK( clk ) , .D( key_c_r_10_23 ) , .Q( key_c_r_11_23 ) );
  DFF_X1 key_c_r_reg_11_24 (.CK( clk ) , .D( key_c_r_10_24 ) , .Q( key_c_r_11_24 ) );
  DFF_X1 key_c_r_reg_11_25 (.CK( clk ) , .D( key_c_r_10_25 ) , .Q( key_c_r_11_25 ) );
  DFF_X1 key_c_r_reg_11_26 (.CK( clk ) , .D( key_c_r_10_26 ) , .Q( key_c_r_11_26 ) );
  DFF_X1 key_c_r_reg_11_27 (.CK( clk ) , .D( key_c_r_10_27 ) , .Q( key_c_r_11_27 ) );
  DFF_X1 key_c_r_reg_11_28 (.CK( clk ) , .D( key_c_r_10_28 ) , .Q( key_c_r_11_28 ) );
  DFF_X1 key_c_r_reg_11_29 (.CK( clk ) , .D( key_c_r_10_29 ) , .Q( key_c_r_11_29 ) );
  DFF_X1 key_c_r_reg_11_3 (.CK( clk ) , .D( key_c_r_10_3 ) , .Q( key_c_r_11_3 ) );
  DFF_X1 key_c_r_reg_11_30 (.CK( clk ) , .D( key_c_r_10_30 ) , .Q( key_c_r_11_30 ) );
  DFF_X1 key_c_r_reg_11_31 (.CK( clk ) , .D( key_c_r_10_31 ) , .Q( key_c_r_11_31 ) );
  DFF_X1 key_c_r_reg_11_32 (.CK( clk ) , .D( key_c_r_10_32 ) , .Q( key_c_r_11_32 ) );
  DFF_X1 key_c_r_reg_11_33 (.CK( clk ) , .D( key_c_r_10_33 ) , .Q( key_c_r_11_33 ) );
  DFF_X1 key_c_r_reg_11_34 (.CK( clk ) , .D( key_c_r_10_34 ) , .Q( key_c_r_11_34 ) );
  DFF_X1 key_c_r_reg_11_35 (.CK( clk ) , .D( key_c_r_10_35 ) , .Q( key_c_r_11_35 ) );
  DFF_X1 key_c_r_reg_11_36 (.CK( clk ) , .D( key_c_r_10_36 ) , .Q( key_c_r_11_36 ) );
  DFF_X1 key_c_r_reg_11_37 (.CK( clk ) , .D( key_c_r_10_37 ) , .Q( key_c_r_11_37 ) );
  DFF_X1 key_c_r_reg_11_38 (.CK( clk ) , .D( key_c_r_10_38 ) , .Q( key_c_r_11_38 ) );
  DFF_X1 key_c_r_reg_11_39 (.CK( clk ) , .D( key_c_r_10_39 ) , .Q( key_c_r_11_39 ) );
  DFF_X1 key_c_r_reg_11_4 (.CK( clk ) , .D( key_c_r_10_4 ) , .Q( key_c_r_11_4 ) );
  DFF_X1 key_c_r_reg_11_40 (.CK( clk ) , .D( key_c_r_10_40 ) , .Q( key_c_r_11_40 ) );
  DFF_X1 key_c_r_reg_11_41 (.CK( clk ) , .D( key_c_r_10_41 ) , .Q( key_c_r_11_41 ) );
  DFF_X1 key_c_r_reg_11_42 (.CK( clk ) , .D( key_c_r_10_42 ) , .Q( key_c_r_11_42 ) );
  DFF_X1 key_c_r_reg_11_43 (.CK( clk ) , .D( key_c_r_10_43 ) , .Q( key_c_r_11_43 ) );
  DFF_X1 key_c_r_reg_11_44 (.CK( clk ) , .D( key_c_r_10_44 ) , .Q( key_c_r_11_44 ) );
  DFF_X1 key_c_r_reg_11_45 (.CK( clk ) , .D( key_c_r_10_45 ) , .Q( key_c_r_11_45 ) );
  DFF_X1 key_c_r_reg_11_46 (.CK( clk ) , .D( key_c_r_10_46 ) , .Q( key_c_r_11_46 ) );
  DFF_X1 key_c_r_reg_11_47 (.CK( clk ) , .D( key_c_r_10_47 ) , .Q( key_c_r_11_47 ) );
  DFF_X1 key_c_r_reg_11_48 (.CK( clk ) , .D( key_c_r_10_48 ) , .Q( key_c_r_11_48 ) );
  DFF_X1 key_c_r_reg_11_49 (.CK( clk ) , .D( key_c_r_10_49 ) , .Q( key_c_r_11_49 ) );
  DFF_X1 key_c_r_reg_11_5 (.CK( clk ) , .D( key_c_r_10_5 ) , .Q( key_c_r_11_5 ) );
  DFF_X1 key_c_r_reg_11_50 (.CK( clk ) , .D( key_c_r_10_50 ) , .Q( key_c_r_11_50 ) );
  DFF_X1 key_c_r_reg_11_51 (.CK( clk ) , .D( key_c_r_10_51 ) , .Q( key_c_r_11_51 ) );
  DFF_X1 key_c_r_reg_11_52 (.CK( clk ) , .D( key_c_r_10_52 ) , .Q( key_c_r_11_52 ) );
  DFF_X1 key_c_r_reg_11_53 (.CK( clk ) , .D( key_c_r_10_53 ) , .Q( key_c_r_11_53 ) );
  DFF_X1 key_c_r_reg_11_54 (.CK( clk ) , .D( key_c_r_10_54 ) , .Q( key_c_r_11_54 ) );
  DFF_X1 key_c_r_reg_11_55 (.CK( clk ) , .D( key_c_r_10_55 ) , .Q( key_c_r_11_55 ) );
  DFF_X1 key_c_r_reg_11_6 (.CK( clk ) , .D( key_c_r_10_6 ) , .Q( key_c_r_11_6 ) );
  DFF_X1 key_c_r_reg_11_7 (.CK( clk ) , .D( key_c_r_10_7 ) , .Q( key_c_r_11_7 ) );
  DFF_X1 key_c_r_reg_11_8 (.CK( clk ) , .D( key_c_r_10_8 ) , .Q( key_c_r_11_8 ) );
  DFF_X1 key_c_r_reg_11_9 (.CK( clk ) , .D( key_c_r_10_9 ) , .Q( key_c_r_11_9 ) );
  DFF_X1 key_c_r_reg_12_0 (.CK( clk ) , .D( key_c_r_11_0 ) , .Q( key_c_r_12_0 ) );
  DFF_X1 key_c_r_reg_12_1 (.CK( clk ) , .D( key_c_r_11_1 ) , .Q( key_c_r_12_1 ) );
  DFF_X1 key_c_r_reg_12_10 (.CK( clk ) , .D( key_c_r_11_10 ) , .Q( key_c_r_12_10 ) );
  DFF_X1 key_c_r_reg_12_11 (.CK( clk ) , .D( key_c_r_11_11 ) , .Q( key_c_r_12_11 ) );
  DFF_X1 key_c_r_reg_12_12 (.CK( clk ) , .D( key_c_r_11_12 ) , .Q( key_c_r_12_12 ) );
  DFF_X1 key_c_r_reg_12_13 (.CK( clk ) , .D( key_c_r_11_13 ) , .Q( key_c_r_12_13 ) );
  DFF_X1 key_c_r_reg_12_14 (.CK( clk ) , .D( key_c_r_11_14 ) , .Q( key_c_r_12_14 ) );
  DFF_X1 key_c_r_reg_12_15 (.CK( clk ) , .D( key_c_r_11_15 ) , .Q( key_c_r_12_15 ) );
  DFF_X1 key_c_r_reg_12_16 (.CK( clk ) , .D( key_c_r_11_16 ) , .Q( key_c_r_12_16 ) );
  DFF_X1 key_c_r_reg_12_17 (.CK( clk ) , .D( key_c_r_11_17 ) , .Q( key_c_r_12_17 ) );
  DFF_X1 key_c_r_reg_12_18 (.CK( clk ) , .D( key_c_r_11_18 ) , .Q( key_c_r_12_18 ) );
  DFF_X1 key_c_r_reg_12_19 (.CK( clk ) , .D( key_c_r_11_19 ) , .Q( key_c_r_12_19 ) );
  DFF_X1 key_c_r_reg_12_2 (.CK( clk ) , .D( key_c_r_11_2 ) , .Q( key_c_r_12_2 ) );
  DFF_X1 key_c_r_reg_12_20 (.CK( clk ) , .D( key_c_r_11_20 ) , .Q( key_c_r_12_20 ) );
  DFF_X1 key_c_r_reg_12_21 (.CK( clk ) , .D( key_c_r_11_21 ) , .Q( key_c_r_12_21 ) );
  DFF_X1 key_c_r_reg_12_22 (.CK( clk ) , .D( key_c_r_11_22 ) , .Q( key_c_r_12_22 ) );
  DFF_X1 key_c_r_reg_12_23 (.CK( clk ) , .D( key_c_r_11_23 ) , .Q( key_c_r_12_23 ) );
  DFF_X1 key_c_r_reg_12_24 (.CK( clk ) , .D( key_c_r_11_24 ) , .Q( key_c_r_12_24 ) );
  DFF_X1 key_c_r_reg_12_25 (.CK( clk ) , .D( key_c_r_11_25 ) , .Q( key_c_r_12_25 ) );
  DFF_X1 key_c_r_reg_12_26 (.CK( clk ) , .D( key_c_r_11_26 ) , .Q( key_c_r_12_26 ) );
  DFF_X1 key_c_r_reg_12_27 (.CK( clk ) , .D( key_c_r_11_27 ) , .Q( key_c_r_12_27 ) );
  DFF_X1 key_c_r_reg_12_28 (.CK( clk ) , .D( key_c_r_11_28 ) , .Q( key_c_r_12_28 ) );
  DFF_X1 key_c_r_reg_12_29 (.CK( clk ) , .D( key_c_r_11_29 ) , .Q( key_c_r_12_29 ) );
  DFF_X1 key_c_r_reg_12_3 (.CK( clk ) , .D( key_c_r_11_3 ) , .Q( key_c_r_12_3 ) );
  DFF_X1 key_c_r_reg_12_30 (.CK( clk ) , .D( key_c_r_11_30 ) , .Q( key_c_r_12_30 ) );
  DFF_X1 key_c_r_reg_12_31 (.CK( clk ) , .D( key_c_r_11_31 ) , .Q( key_c_r_12_31 ) );
  DFF_X1 key_c_r_reg_12_32 (.CK( clk ) , .D( key_c_r_11_32 ) , .Q( key_c_r_12_32 ) );
  DFF_X1 key_c_r_reg_12_33 (.CK( clk ) , .D( key_c_r_11_33 ) , .Q( key_c_r_12_33 ) );
  DFF_X1 key_c_r_reg_12_34 (.CK( clk ) , .D( key_c_r_11_34 ) , .Q( key_c_r_12_34 ) );
  DFF_X1 key_c_r_reg_12_35 (.CK( clk ) , .D( key_c_r_11_35 ) , .Q( key_c_r_12_35 ) );
  DFF_X1 key_c_r_reg_12_36 (.CK( clk ) , .D( key_c_r_11_36 ) , .Q( key_c_r_12_36 ) );
  DFF_X1 key_c_r_reg_12_37 (.CK( clk ) , .D( key_c_r_11_37 ) , .Q( key_c_r_12_37 ) );
  DFF_X1 key_c_r_reg_12_38 (.CK( clk ) , .D( key_c_r_11_38 ) , .Q( key_c_r_12_38 ) );
  DFF_X1 key_c_r_reg_12_39 (.CK( clk ) , .D( key_c_r_11_39 ) , .Q( key_c_r_12_39 ) );
  DFF_X1 key_c_r_reg_12_4 (.CK( clk ) , .D( key_c_r_11_4 ) , .Q( key_c_r_12_4 ) );
  DFF_X1 key_c_r_reg_12_40 (.CK( clk ) , .D( key_c_r_11_40 ) , .Q( key_c_r_12_40 ) );
  DFF_X1 key_c_r_reg_12_41 (.CK( clk ) , .D( key_c_r_11_41 ) , .Q( key_c_r_12_41 ) );
  DFF_X1 key_c_r_reg_12_42 (.CK( clk ) , .D( key_c_r_11_42 ) , .Q( key_c_r_12_42 ) );
  DFF_X1 key_c_r_reg_12_43 (.CK( clk ) , .D( key_c_r_11_43 ) , .Q( key_c_r_12_43 ) );
  DFF_X1 key_c_r_reg_12_44 (.CK( clk ) , .D( key_c_r_11_44 ) , .Q( key_c_r_12_44 ) );
  DFF_X1 key_c_r_reg_12_45 (.CK( clk ) , .D( key_c_r_11_45 ) , .Q( key_c_r_12_45 ) );
  DFF_X1 key_c_r_reg_12_46 (.CK( clk ) , .D( key_c_r_11_46 ) , .Q( key_c_r_12_46 ) );
  DFF_X1 key_c_r_reg_12_47 (.CK( clk ) , .D( key_c_r_11_47 ) , .Q( key_c_r_12_47 ) );
  DFF_X1 key_c_r_reg_12_48 (.CK( clk ) , .D( key_c_r_11_48 ) , .Q( key_c_r_12_48 ) );
  DFF_X1 key_c_r_reg_12_49 (.CK( clk ) , .D( key_c_r_11_49 ) , .Q( key_c_r_12_49 ) );
  DFF_X1 key_c_r_reg_12_5 (.CK( clk ) , .D( key_c_r_11_5 ) , .Q( key_c_r_12_5 ) );
  DFF_X1 key_c_r_reg_12_50 (.CK( clk ) , .D( key_c_r_11_50 ) , .Q( key_c_r_12_50 ) );
  DFF_X1 key_c_r_reg_12_51 (.CK( clk ) , .D( key_c_r_11_51 ) , .Q( key_c_r_12_51 ) );
  DFF_X1 key_c_r_reg_12_52 (.CK( clk ) , .D( key_c_r_11_52 ) , .Q( key_c_r_12_52 ) );
  DFF_X1 key_c_r_reg_12_53 (.CK( clk ) , .D( key_c_r_11_53 ) , .Q( key_c_r_12_53 ) );
  DFF_X1 key_c_r_reg_12_54 (.CK( clk ) , .D( key_c_r_11_54 ) , .Q( key_c_r_12_54 ) );
  DFF_X1 key_c_r_reg_12_55 (.CK( clk ) , .D( key_c_r_11_55 ) , .Q( key_c_r_12_55 ) );
  DFF_X1 key_c_r_reg_12_6 (.CK( clk ) , .D( key_c_r_11_6 ) , .Q( key_c_r_12_6 ) );
  DFF_X1 key_c_r_reg_12_7 (.CK( clk ) , .D( key_c_r_11_7 ) , .Q( key_c_r_12_7 ) );
  DFF_X1 key_c_r_reg_12_8 (.CK( clk ) , .D( key_c_r_11_8 ) , .Q( key_c_r_12_8 ) );
  DFF_X1 key_c_r_reg_12_9 (.CK( clk ) , .D( key_c_r_11_9 ) , .Q( key_c_r_12_9 ) );
  DFF_X1 key_c_r_reg_13_0 (.CK( clk ) , .D( key_c_r_12_0 ) , .Q( key_c_r_13_0 ) );
  DFF_X1 key_c_r_reg_13_1 (.CK( clk ) , .D( key_c_r_12_1 ) , .Q( key_c_r_13_1 ) );
  DFF_X1 key_c_r_reg_13_10 (.CK( clk ) , .D( key_c_r_12_10 ) , .Q( key_c_r_13_10 ) );
  DFF_X1 key_c_r_reg_13_11 (.CK( clk ) , .D( key_c_r_12_11 ) , .Q( key_c_r_13_11 ) );
  DFF_X1 key_c_r_reg_13_12 (.CK( clk ) , .D( key_c_r_12_12 ) , .Q( key_c_r_13_12 ) );
  DFF_X1 key_c_r_reg_13_13 (.CK( clk ) , .D( key_c_r_12_13 ) , .Q( key_c_r_13_13 ) );
  DFF_X1 key_c_r_reg_13_14 (.CK( clk ) , .D( key_c_r_12_14 ) , .Q( key_c_r_13_14 ) );
  DFF_X1 key_c_r_reg_13_15 (.CK( clk ) , .D( key_c_r_12_15 ) , .Q( key_c_r_13_15 ) );
  DFF_X1 key_c_r_reg_13_16 (.CK( clk ) , .D( key_c_r_12_16 ) , .Q( key_c_r_13_16 ) );
  DFF_X1 key_c_r_reg_13_17 (.CK( clk ) , .D( key_c_r_12_17 ) , .Q( key_c_r_13_17 ) );
  DFF_X1 key_c_r_reg_13_18 (.CK( clk ) , .D( key_c_r_12_18 ) , .Q( key_c_r_13_18 ) );
  DFF_X1 key_c_r_reg_13_19 (.CK( clk ) , .D( key_c_r_12_19 ) , .Q( key_c_r_13_19 ) );
  DFF_X1 key_c_r_reg_13_2 (.CK( clk ) , .D( key_c_r_12_2 ) , .Q( key_c_r_13_2 ) );
  DFF_X1 key_c_r_reg_13_20 (.CK( clk ) , .D( key_c_r_12_20 ) , .Q( key_c_r_13_20 ) );
  DFF_X1 key_c_r_reg_13_21 (.CK( clk ) , .D( key_c_r_12_21 ) , .Q( key_c_r_13_21 ) );
  DFF_X1 key_c_r_reg_13_22 (.CK( clk ) , .D( key_c_r_12_22 ) , .Q( key_c_r_13_22 ) );
  DFF_X1 key_c_r_reg_13_23 (.CK( clk ) , .D( key_c_r_12_23 ) , .Q( key_c_r_13_23 ) );
  DFF_X1 key_c_r_reg_13_24 (.CK( clk ) , .D( key_c_r_12_24 ) , .Q( key_c_r_13_24 ) );
  DFF_X1 key_c_r_reg_13_25 (.CK( clk ) , .D( key_c_r_12_25 ) , .Q( key_c_r_13_25 ) );
  DFF_X1 key_c_r_reg_13_26 (.CK( clk ) , .D( key_c_r_12_26 ) , .Q( key_c_r_13_26 ) );
  DFF_X1 key_c_r_reg_13_27 (.CK( clk ) , .D( key_c_r_12_27 ) , .Q( key_c_r_13_27 ) );
  DFF_X1 key_c_r_reg_13_28 (.CK( clk ) , .D( key_c_r_12_28 ) , .Q( key_c_r_13_28 ) );
  DFF_X1 key_c_r_reg_13_29 (.CK( clk ) , .D( key_c_r_12_29 ) , .Q( key_c_r_13_29 ) );
  DFF_X1 key_c_r_reg_13_3 (.CK( clk ) , .D( key_c_r_12_3 ) , .Q( key_c_r_13_3 ) );
  DFF_X1 key_c_r_reg_13_30 (.CK( clk ) , .D( key_c_r_12_30 ) , .Q( key_c_r_13_30 ) );
  DFF_X1 key_c_r_reg_13_31 (.CK( clk ) , .D( key_c_r_12_31 ) , .Q( key_c_r_13_31 ) );
  DFF_X1 key_c_r_reg_13_32 (.CK( clk ) , .D( key_c_r_12_32 ) , .Q( key_c_r_13_32 ) );
  DFF_X1 key_c_r_reg_13_33 (.CK( clk ) , .D( key_c_r_12_33 ) , .Q( key_c_r_13_33 ) );
  DFF_X1 key_c_r_reg_13_34 (.CK( clk ) , .D( key_c_r_12_34 ) , .Q( key_c_r_13_34 ) );
  DFF_X1 key_c_r_reg_13_35 (.CK( clk ) , .D( key_c_r_12_35 ) , .Q( key_c_r_13_35 ) );
  DFF_X1 key_c_r_reg_13_36 (.CK( clk ) , .D( key_c_r_12_36 ) , .Q( key_c_r_13_36 ) );
  DFF_X1 key_c_r_reg_13_37 (.CK( clk ) , .D( key_c_r_12_37 ) , .Q( key_c_r_13_37 ) );
  DFF_X1 key_c_r_reg_13_38 (.CK( clk ) , .D( key_c_r_12_38 ) , .Q( key_c_r_13_38 ) );
  DFF_X1 key_c_r_reg_13_39 (.CK( clk ) , .D( key_c_r_12_39 ) , .Q( key_c_r_13_39 ) );
  DFF_X1 key_c_r_reg_13_4 (.CK( clk ) , .D( key_c_r_12_4 ) , .Q( key_c_r_13_4 ) );
  DFF_X1 key_c_r_reg_13_40 (.CK( clk ) , .D( key_c_r_12_40 ) , .Q( key_c_r_13_40 ) );
  DFF_X1 key_c_r_reg_13_41 (.CK( clk ) , .D( key_c_r_12_41 ) , .Q( key_c_r_13_41 ) );
  DFF_X1 key_c_r_reg_13_42 (.CK( clk ) , .D( key_c_r_12_42 ) , .Q( key_c_r_13_42 ) );
  DFF_X1 key_c_r_reg_13_43 (.CK( clk ) , .D( key_c_r_12_43 ) , .Q( key_c_r_13_43 ) );
  DFF_X1 key_c_r_reg_13_44 (.CK( clk ) , .D( key_c_r_12_44 ) , .Q( key_c_r_13_44 ) );
  DFF_X1 key_c_r_reg_13_45 (.CK( clk ) , .D( key_c_r_12_45 ) , .Q( key_c_r_13_45 ) );
  DFF_X1 key_c_r_reg_13_46 (.CK( clk ) , .D( key_c_r_12_46 ) , .Q( key_c_r_13_46 ) );
  DFF_X1 key_c_r_reg_13_47 (.CK( clk ) , .D( key_c_r_12_47 ) , .Q( key_c_r_13_47 ) );
  DFF_X1 key_c_r_reg_13_48 (.CK( clk ) , .D( key_c_r_12_48 ) , .Q( key_c_r_13_48 ) );
  DFF_X1 key_c_r_reg_13_49 (.CK( clk ) , .D( key_c_r_12_49 ) , .Q( key_c_r_13_49 ) );
  DFF_X1 key_c_r_reg_13_5 (.CK( clk ) , .D( key_c_r_12_5 ) , .Q( key_c_r_13_5 ) );
  DFF_X1 key_c_r_reg_13_50 (.CK( clk ) , .D( key_c_r_12_50 ) , .Q( key_c_r_13_50 ) );
  DFF_X1 key_c_r_reg_13_51 (.CK( clk ) , .D( key_c_r_12_51 ) , .Q( key_c_r_13_51 ) );
  DFF_X1 key_c_r_reg_13_52 (.CK( clk ) , .D( key_c_r_12_52 ) , .Q( key_c_r_13_52 ) );
  DFF_X1 key_c_r_reg_13_53 (.CK( clk ) , .D( key_c_r_12_53 ) , .Q( key_c_r_13_53 ) );
  DFF_X1 key_c_r_reg_13_54 (.CK( clk ) , .D( key_c_r_12_54 ) , .Q( key_c_r_13_54 ) );
  DFF_X1 key_c_r_reg_13_55 (.CK( clk ) , .D( key_c_r_12_55 ) , .Q( key_c_r_13_55 ) );
  DFF_X1 key_c_r_reg_13_6 (.CK( clk ) , .D( key_c_r_12_6 ) , .Q( key_c_r_13_6 ) );
  DFF_X1 key_c_r_reg_13_7 (.CK( clk ) , .D( key_c_r_12_7 ) , .Q( key_c_r_13_7 ) );
  DFF_X1 key_c_r_reg_13_8 (.CK( clk ) , .D( key_c_r_12_8 ) , .Q( key_c_r_13_8 ) );
  DFF_X1 key_c_r_reg_13_9 (.CK( clk ) , .D( key_c_r_12_9 ) , .Q( key_c_r_13_9 ) );
  DFF_X1 key_c_r_reg_14_0 (.CK( clk ) , .D( key_c_r_13_0 ) , .Q( key_c_r_14_0 ) );
  DFF_X1 key_c_r_reg_14_1 (.CK( clk ) , .D( key_c_r_13_1 ) , .Q( key_c_r_14_1 ) );
  DFF_X1 key_c_r_reg_14_10 (.CK( clk ) , .D( key_c_r_13_10 ) , .Q( key_c_r_14_10 ) );
  DFF_X1 key_c_r_reg_14_11 (.CK( clk ) , .D( key_c_r_13_11 ) , .Q( key_c_r_14_11 ) );
  DFF_X1 key_c_r_reg_14_12 (.CK( clk ) , .D( key_c_r_13_12 ) , .Q( key_c_r_14_12 ) );
  DFF_X1 key_c_r_reg_14_13 (.CK( clk ) , .D( key_c_r_13_13 ) , .Q( key_c_r_14_13 ) );
  DFF_X1 key_c_r_reg_14_14 (.CK( clk ) , .D( key_c_r_13_14 ) , .Q( key_c_r_14_14 ) );
  DFF_X1 key_c_r_reg_14_15 (.CK( clk ) , .D( key_c_r_13_15 ) , .Q( key_c_r_14_15 ) );
  DFF_X1 key_c_r_reg_14_16 (.CK( clk ) , .D( key_c_r_13_16 ) , .Q( key_c_r_14_16 ) );
  DFF_X1 key_c_r_reg_14_17 (.CK( clk ) , .D( key_c_r_13_17 ) , .Q( key_c_r_14_17 ) );
  DFF_X1 key_c_r_reg_14_18 (.CK( clk ) , .D( key_c_r_13_18 ) , .Q( key_c_r_14_18 ) );
  DFF_X1 key_c_r_reg_14_19 (.CK( clk ) , .D( key_c_r_13_19 ) , .Q( key_c_r_14_19 ) );
  DFF_X1 key_c_r_reg_14_2 (.CK( clk ) , .D( key_c_r_13_2 ) , .Q( key_c_r_14_2 ) );
  DFF_X1 key_c_r_reg_14_20 (.CK( clk ) , .D( key_c_r_13_20 ) , .Q( key_c_r_14_20 ) );
  DFF_X1 key_c_r_reg_14_21 (.CK( clk ) , .D( key_c_r_13_21 ) , .Q( key_c_r_14_21 ) );
  DFF_X1 key_c_r_reg_14_22 (.CK( clk ) , .D( key_c_r_13_22 ) , .Q( key_c_r_14_22 ) );
  DFF_X1 key_c_r_reg_14_23 (.CK( clk ) , .D( key_c_r_13_23 ) , .Q( key_c_r_14_23 ) );
  DFF_X1 key_c_r_reg_14_24 (.CK( clk ) , .D( key_c_r_13_24 ) , .Q( key_c_r_14_24 ) );
  DFF_X1 key_c_r_reg_14_25 (.CK( clk ) , .D( key_c_r_13_25 ) , .Q( key_c_r_14_25 ) );
  DFF_X1 key_c_r_reg_14_26 (.CK( clk ) , .D( key_c_r_13_26 ) , .Q( key_c_r_14_26 ) );
  DFF_X1 key_c_r_reg_14_27 (.CK( clk ) , .D( key_c_r_13_27 ) , .Q( key_c_r_14_27 ) );
  DFF_X1 key_c_r_reg_14_28 (.CK( clk ) , .D( key_c_r_13_28 ) , .Q( key_c_r_14_28 ) );
  DFF_X1 key_c_r_reg_14_29 (.CK( clk ) , .D( key_c_r_13_29 ) , .Q( key_c_r_14_29 ) );
  DFF_X1 key_c_r_reg_14_3 (.CK( clk ) , .D( key_c_r_13_3 ) , .Q( key_c_r_14_3 ) );
  DFF_X1 key_c_r_reg_14_30 (.CK( clk ) , .D( key_c_r_13_30 ) , .Q( key_c_r_14_30 ) );
  DFF_X1 key_c_r_reg_14_31 (.CK( clk ) , .D( key_c_r_13_31 ) , .Q( key_c_r_14_31 ) );
  DFF_X1 key_c_r_reg_14_32 (.CK( clk ) , .D( key_c_r_13_32 ) , .Q( key_c_r_14_32 ) );
  DFF_X1 key_c_r_reg_14_33 (.CK( clk ) , .D( key_c_r_13_33 ) , .Q( key_c_r_14_33 ) );
  DFF_X1 key_c_r_reg_14_34 (.CK( clk ) , .D( key_c_r_13_34 ) , .Q( key_c_r_14_34 ) );
  DFF_X1 key_c_r_reg_14_35 (.CK( clk ) , .D( key_c_r_13_35 ) , .Q( key_c_r_14_35 ) );
  DFF_X1 key_c_r_reg_14_36 (.CK( clk ) , .D( key_c_r_13_36 ) , .Q( key_c_r_14_36 ) );
  DFF_X1 key_c_r_reg_14_37 (.CK( clk ) , .D( key_c_r_13_37 ) , .Q( key_c_r_14_37 ) );
  DFF_X1 key_c_r_reg_14_38 (.CK( clk ) , .D( key_c_r_13_38 ) , .Q( key_c_r_14_38 ) );
  DFF_X1 key_c_r_reg_14_39 (.CK( clk ) , .D( key_c_r_13_39 ) , .Q( key_c_r_14_39 ) );
  DFF_X1 key_c_r_reg_14_4 (.CK( clk ) , .D( key_c_r_13_4 ) , .Q( key_c_r_14_4 ) );
  DFF_X1 key_c_r_reg_14_40 (.CK( clk ) , .D( key_c_r_13_40 ) , .Q( key_c_r_14_40 ) );
  DFF_X1 key_c_r_reg_14_41 (.CK( clk ) , .D( key_c_r_13_41 ) , .Q( key_c_r_14_41 ) );
  DFF_X1 key_c_r_reg_14_42 (.CK( clk ) , .D( key_c_r_13_42 ) , .Q( key_c_r_14_42 ) );
  DFF_X1 key_c_r_reg_14_43 (.CK( clk ) , .D( key_c_r_13_43 ) , .Q( key_c_r_14_43 ) );
  DFF_X1 key_c_r_reg_14_44 (.CK( clk ) , .D( key_c_r_13_44 ) , .Q( key_c_r_14_44 ) );
  DFF_X1 key_c_r_reg_14_45 (.CK( clk ) , .D( key_c_r_13_45 ) , .Q( key_c_r_14_45 ) );
  DFF_X1 key_c_r_reg_14_46 (.CK( clk ) , .D( key_c_r_13_46 ) , .Q( key_c_r_14_46 ) );
  DFF_X1 key_c_r_reg_14_47 (.CK( clk ) , .D( key_c_r_13_47 ) , .Q( key_c_r_14_47 ) );
  DFF_X1 key_c_r_reg_14_48 (.CK( clk ) , .D( key_c_r_13_48 ) , .Q( key_c_r_14_48 ) );
  DFF_X1 key_c_r_reg_14_49 (.CK( clk ) , .D( key_c_r_13_49 ) , .Q( key_c_r_14_49 ) );
  DFF_X1 key_c_r_reg_14_5 (.CK( clk ) , .D( key_c_r_13_5 ) , .Q( key_c_r_14_5 ) );
  DFF_X1 key_c_r_reg_14_50 (.CK( clk ) , .D( key_c_r_13_50 ) , .Q( key_c_r_14_50 ) );
  DFF_X1 key_c_r_reg_14_51 (.CK( clk ) , .D( key_c_r_13_51 ) , .Q( key_c_r_14_51 ) );
  DFF_X1 key_c_r_reg_14_52 (.CK( clk ) , .D( key_c_r_13_52 ) , .Q( key_c_r_14_52 ) );
  DFF_X1 key_c_r_reg_14_53 (.CK( clk ) , .D( key_c_r_13_53 ) , .Q( key_c_r_14_53 ) );
  DFF_X1 key_c_r_reg_14_54 (.CK( clk ) , .D( key_c_r_13_54 ) , .Q( key_c_r_14_54 ) );
  DFF_X1 key_c_r_reg_14_55 (.CK( clk ) , .D( key_c_r_13_55 ) , .Q( key_c_r_14_55 ) );
  DFF_X1 key_c_r_reg_14_6 (.CK( clk ) , .D( key_c_r_13_6 ) , .Q( key_c_r_14_6 ) );
  DFF_X1 key_c_r_reg_14_7 (.CK( clk ) , .D( key_c_r_13_7 ) , .Q( key_c_r_14_7 ) );
  DFF_X1 key_c_r_reg_14_8 (.CK( clk ) , .D( key_c_r_13_8 ) , .Q( key_c_r_14_8 ) );
  DFF_X1 key_c_r_reg_14_9 (.CK( clk ) , .D( key_c_r_13_9 ) , .Q( key_c_r_14_9 ) );
  DFF_X1 key_c_r_reg_15_0 (.CK( clk ) , .D( key_c_r_14_0 ) , .Q( key_c_r_15_0 ) );
  DFF_X1 key_c_r_reg_15_1 (.CK( clk ) , .D( key_c_r_14_1 ) , .Q( key_c_r_15_1 ) );
  DFF_X1 key_c_r_reg_15_10 (.CK( clk ) , .D( key_c_r_14_10 ) , .Q( key_c_r_15_10 ) );
  DFF_X1 key_c_r_reg_15_11 (.CK( clk ) , .D( key_c_r_14_11 ) , .Q( key_c_r_15_11 ) );
  DFF_X1 key_c_r_reg_15_12 (.CK( clk ) , .D( key_c_r_14_12 ) , .Q( key_c_r_15_12 ) );
  DFF_X1 key_c_r_reg_15_13 (.CK( clk ) , .D( key_c_r_14_13 ) , .Q( key_c_r_15_13 ) );
  DFF_X1 key_c_r_reg_15_14 (.CK( clk ) , .D( key_c_r_14_14 ) , .Q( key_c_r_15_14 ) );
  DFF_X1 key_c_r_reg_15_15 (.CK( clk ) , .D( key_c_r_14_15 ) , .Q( key_c_r_15_15 ) );
  DFF_X1 key_c_r_reg_15_16 (.CK( clk ) , .D( key_c_r_14_16 ) , .Q( key_c_r_15_16 ) );
  DFF_X1 key_c_r_reg_15_17 (.CK( clk ) , .D( key_c_r_14_17 ) , .Q( key_c_r_15_17 ) );
  DFF_X1 key_c_r_reg_15_18 (.CK( clk ) , .D( key_c_r_14_18 ) , .Q( key_c_r_15_18 ) );
  DFF_X1 key_c_r_reg_15_19 (.CK( clk ) , .D( key_c_r_14_19 ) , .Q( key_c_r_15_19 ) );
  DFF_X1 key_c_r_reg_15_2 (.CK( clk ) , .D( key_c_r_14_2 ) , .Q( key_c_r_15_2 ) );
  DFF_X1 key_c_r_reg_15_20 (.CK( clk ) , .D( key_c_r_14_20 ) , .Q( key_c_r_15_20 ) );
  DFF_X1 key_c_r_reg_15_21 (.CK( clk ) , .D( key_c_r_14_21 ) , .Q( key_c_r_15_21 ) );
  DFF_X1 key_c_r_reg_15_22 (.CK( clk ) , .D( key_c_r_14_22 ) , .Q( key_c_r_15_22 ) );
  DFF_X1 key_c_r_reg_15_23 (.CK( clk ) , .D( key_c_r_14_23 ) , .Q( key_c_r_15_23 ) );
  DFF_X1 key_c_r_reg_15_24 (.CK( clk ) , .D( key_c_r_14_24 ) , .Q( key_c_r_15_24 ) );
  DFF_X1 key_c_r_reg_15_25 (.CK( clk ) , .D( key_c_r_14_25 ) , .Q( key_c_r_15_25 ) );
  DFF_X1 key_c_r_reg_15_26 (.CK( clk ) , .D( key_c_r_14_26 ) , .Q( key_c_r_15_26 ) );
  DFF_X1 key_c_r_reg_15_27 (.CK( clk ) , .D( key_c_r_14_27 ) , .Q( key_c_r_15_27 ) );
  DFF_X1 key_c_r_reg_15_28 (.CK( clk ) , .D( key_c_r_14_28 ) , .Q( key_c_r_15_28 ) );
  DFF_X1 key_c_r_reg_15_29 (.CK( clk ) , .D( key_c_r_14_29 ) , .Q( key_c_r_15_29 ) );
  DFF_X1 key_c_r_reg_15_3 (.CK( clk ) , .D( key_c_r_14_3 ) , .Q( key_c_r_15_3 ) );
  DFF_X1 key_c_r_reg_15_30 (.CK( clk ) , .D( key_c_r_14_30 ) , .Q( key_c_r_15_30 ) );
  DFF_X1 key_c_r_reg_15_31 (.CK( clk ) , .D( key_c_r_14_31 ) , .Q( key_c_r_15_31 ) );
  DFF_X1 key_c_r_reg_15_32 (.CK( clk ) , .D( key_c_r_14_32 ) , .Q( key_c_r_15_32 ) );
  DFF_X1 key_c_r_reg_15_33 (.CK( clk ) , .D( key_c_r_14_33 ) , .Q( key_c_r_15_33 ) );
  DFF_X1 key_c_r_reg_15_34 (.CK( clk ) , .D( key_c_r_14_34 ) , .Q( key_c_r_15_34 ) );
  DFF_X1 key_c_r_reg_15_35 (.CK( clk ) , .D( key_c_r_14_35 ) , .Q( key_c_r_15_35 ) );
  DFF_X1 key_c_r_reg_15_36 (.CK( clk ) , .D( key_c_r_14_36 ) , .Q( key_c_r_15_36 ) );
  DFF_X1 key_c_r_reg_15_37 (.CK( clk ) , .D( key_c_r_14_37 ) , .Q( key_c_r_15_37 ) );
  DFF_X1 key_c_r_reg_15_38 (.CK( clk ) , .D( key_c_r_14_38 ) , .Q( key_c_r_15_38 ) );
  DFF_X1 key_c_r_reg_15_39 (.CK( clk ) , .D( key_c_r_14_39 ) , .Q( key_c_r_15_39 ) );
  DFF_X1 key_c_r_reg_15_4 (.CK( clk ) , .D( key_c_r_14_4 ) , .Q( key_c_r_15_4 ) );
  DFF_X1 key_c_r_reg_15_40 (.CK( clk ) , .D( key_c_r_14_40 ) , .Q( key_c_r_15_40 ) );
  DFF_X1 key_c_r_reg_15_41 (.CK( clk ) , .D( key_c_r_14_41 ) , .Q( key_c_r_15_41 ) );
  DFF_X1 key_c_r_reg_15_42 (.CK( clk ) , .D( key_c_r_14_42 ) , .Q( key_c_r_15_42 ) );
  DFF_X1 key_c_r_reg_15_43 (.CK( clk ) , .D( key_c_r_14_43 ) , .Q( key_c_r_15_43 ) );
  DFF_X1 key_c_r_reg_15_44 (.CK( clk ) , .D( key_c_r_14_44 ) , .Q( key_c_r_15_44 ) );
  DFF_X1 key_c_r_reg_15_45 (.CK( clk ) , .D( key_c_r_14_45 ) , .Q( key_c_r_15_45 ) );
  DFF_X1 key_c_r_reg_15_46 (.CK( clk ) , .D( key_c_r_14_46 ) , .Q( key_c_r_15_46 ) );
  DFF_X1 key_c_r_reg_15_47 (.CK( clk ) , .D( key_c_r_14_47 ) , .Q( key_c_r_15_47 ) );
  DFF_X1 key_c_r_reg_15_48 (.CK( clk ) , .D( key_c_r_14_48 ) , .Q( key_c_r_15_48 ) );
  DFF_X1 key_c_r_reg_15_49 (.CK( clk ) , .D( key_c_r_14_49 ) , .Q( key_c_r_15_49 ) );
  DFF_X1 key_c_r_reg_15_5 (.CK( clk ) , .D( key_c_r_14_5 ) , .Q( key_c_r_15_5 ) );
  DFF_X1 key_c_r_reg_15_50 (.CK( clk ) , .D( key_c_r_14_50 ) , .Q( key_c_r_15_50 ) );
  DFF_X1 key_c_r_reg_15_51 (.CK( clk ) , .D( key_c_r_14_51 ) , .Q( key_c_r_15_51 ) );
  DFF_X1 key_c_r_reg_15_52 (.CK( clk ) , .D( key_c_r_14_52 ) , .Q( key_c_r_15_52 ) );
  DFF_X1 key_c_r_reg_15_53 (.CK( clk ) , .D( key_c_r_14_53 ) , .Q( key_c_r_15_53 ) );
  DFF_X1 key_c_r_reg_15_54 (.CK( clk ) , .D( key_c_r_14_54 ) , .Q( key_c_r_15_54 ) );
  DFF_X1 key_c_r_reg_15_55 (.CK( clk ) , .D( key_c_r_14_55 ) , .Q( key_c_r_15_55 ) );
  DFF_X1 key_c_r_reg_15_6 (.CK( clk ) , .D( key_c_r_14_6 ) , .Q( key_c_r_15_6 ) );
  DFF_X1 key_c_r_reg_15_7 (.CK( clk ) , .D( key_c_r_14_7 ) , .Q( key_c_r_15_7 ) );
  DFF_X1 key_c_r_reg_15_8 (.CK( clk ) , .D( key_c_r_14_8 ) , .Q( key_c_r_15_8 ) );
  DFF_X1 key_c_r_reg_15_9 (.CK( clk ) , .D( key_c_r_14_9 ) , .Q( key_c_r_15_9 ) );
  DFF_X1 key_c_r_reg_16_0 (.CK( clk ) , .D( key_c_r_15_0 ) , .Q( key_c_r_16_0 ) );
  DFF_X1 key_c_r_reg_16_1 (.CK( clk ) , .D( key_c_r_15_1 ) , .Q( key_c_r_16_1 ) );
  DFF_X1 key_c_r_reg_16_10 (.CK( clk ) , .D( key_c_r_15_10 ) , .Q( key_c_r_16_10 ) );
  DFF_X1 key_c_r_reg_16_11 (.CK( clk ) , .D( key_c_r_15_11 ) , .Q( key_c_r_16_11 ) );
  DFF_X1 key_c_r_reg_16_12 (.CK( clk ) , .D( key_c_r_15_12 ) , .Q( key_c_r_16_12 ) );
  DFF_X1 key_c_r_reg_16_13 (.CK( clk ) , .D( key_c_r_15_13 ) , .Q( key_c_r_16_13 ) );
  DFF_X1 key_c_r_reg_16_14 (.CK( clk ) , .D( key_c_r_15_14 ) , .Q( key_c_r_16_14 ) );
  DFF_X1 key_c_r_reg_16_15 (.CK( clk ) , .D( key_c_r_15_15 ) , .Q( key_c_r_16_15 ) );
  DFF_X1 key_c_r_reg_16_16 (.CK( clk ) , .D( key_c_r_15_16 ) , .Q( key_c_r_16_16 ) );
  DFF_X1 key_c_r_reg_16_17 (.CK( clk ) , .D( key_c_r_15_17 ) , .Q( key_c_r_16_17 ) );
  DFF_X1 key_c_r_reg_16_18 (.CK( clk ) , .D( key_c_r_15_18 ) , .Q( key_c_r_16_18 ) );
  DFF_X1 key_c_r_reg_16_19 (.CK( clk ) , .D( key_c_r_15_19 ) , .Q( key_c_r_16_19 ) );
  DFF_X1 key_c_r_reg_16_2 (.CK( clk ) , .D( key_c_r_15_2 ) , .Q( key_c_r_16_2 ) );
  DFF_X1 key_c_r_reg_16_20 (.CK( clk ) , .D( key_c_r_15_20 ) , .Q( key_c_r_16_20 ) );
  DFF_X1 key_c_r_reg_16_21 (.CK( clk ) , .D( key_c_r_15_21 ) , .Q( key_c_r_16_21 ) );
  DFF_X1 key_c_r_reg_16_22 (.CK( clk ) , .D( key_c_r_15_22 ) , .Q( key_c_r_16_22 ) );
  DFF_X1 key_c_r_reg_16_23 (.CK( clk ) , .D( key_c_r_15_23 ) , .Q( key_c_r_16_23 ) );
  DFF_X1 key_c_r_reg_16_24 (.CK( clk ) , .D( key_c_r_15_24 ) , .Q( key_c_r_16_24 ) );
  DFF_X1 key_c_r_reg_16_25 (.CK( clk ) , .D( key_c_r_15_25 ) , .Q( key_c_r_16_25 ) );
  DFF_X1 key_c_r_reg_16_26 (.CK( clk ) , .D( key_c_r_15_26 ) , .Q( key_c_r_16_26 ) );
  DFF_X1 key_c_r_reg_16_27 (.CK( clk ) , .D( key_c_r_15_27 ) , .Q( key_c_r_16_27 ) );
  DFF_X1 key_c_r_reg_16_28 (.CK( clk ) , .D( key_c_r_15_28 ) , .Q( key_c_r_16_28 ) );
  DFF_X1 key_c_r_reg_16_29 (.CK( clk ) , .D( key_c_r_15_29 ) , .Q( key_c_r_16_29 ) );
  DFF_X1 key_c_r_reg_16_3 (.CK( clk ) , .D( key_c_r_15_3 ) , .Q( key_c_r_16_3 ) );
  DFF_X1 key_c_r_reg_16_30 (.CK( clk ) , .D( key_c_r_15_30 ) , .Q( key_c_r_16_30 ) );
  DFF_X1 key_c_r_reg_16_31 (.CK( clk ) , .D( key_c_r_15_31 ) , .Q( key_c_r_16_31 ) );
  DFF_X1 key_c_r_reg_16_32 (.CK( clk ) , .D( key_c_r_15_32 ) , .Q( key_c_r_16_32 ) );
  DFF_X1 key_c_r_reg_16_33 (.CK( clk ) , .D( key_c_r_15_33 ) , .Q( key_c_r_16_33 ) );
  DFF_X1 key_c_r_reg_16_34 (.CK( clk ) , .D( key_c_r_15_34 ) , .Q( key_c_r_16_34 ) );
  DFF_X1 key_c_r_reg_16_35 (.CK( clk ) , .D( key_c_r_15_35 ) , .Q( key_c_r_16_35 ) );
  DFF_X1 key_c_r_reg_16_36 (.CK( clk ) , .D( key_c_r_15_36 ) , .Q( key_c_r_16_36 ) );
  DFF_X1 key_c_r_reg_16_37 (.CK( clk ) , .D( key_c_r_15_37 ) , .Q( key_c_r_16_37 ) );
  DFF_X1 key_c_r_reg_16_38 (.CK( clk ) , .D( key_c_r_15_38 ) , .Q( key_c_r_16_38 ) );
  DFF_X1 key_c_r_reg_16_39 (.CK( clk ) , .D( key_c_r_15_39 ) , .Q( key_c_r_16_39 ) );
  DFF_X1 key_c_r_reg_16_4 (.CK( clk ) , .D( key_c_r_15_4 ) , .Q( key_c_r_16_4 ) );
  DFF_X1 key_c_r_reg_16_40 (.CK( clk ) , .D( key_c_r_15_40 ) , .Q( key_c_r_16_40 ) );
  DFF_X1 key_c_r_reg_16_41 (.CK( clk ) , .D( key_c_r_15_41 ) , .Q( key_c_r_16_41 ) );
  DFF_X1 key_c_r_reg_16_42 (.CK( clk ) , .D( key_c_r_15_42 ) , .Q( key_c_r_16_42 ) );
  DFF_X1 key_c_r_reg_16_43 (.CK( clk ) , .D( key_c_r_15_43 ) , .Q( key_c_r_16_43 ) );
  DFF_X1 key_c_r_reg_16_44 (.CK( clk ) , .D( key_c_r_15_44 ) , .Q( key_c_r_16_44 ) );
  DFF_X1 key_c_r_reg_16_45 (.CK( clk ) , .D( key_c_r_15_45 ) , .Q( key_c_r_16_45 ) );
  DFF_X1 key_c_r_reg_16_46 (.CK( clk ) , .D( key_c_r_15_46 ) , .Q( key_c_r_16_46 ) );
  DFF_X1 key_c_r_reg_16_47 (.CK( clk ) , .D( key_c_r_15_47 ) , .Q( key_c_r_16_47 ) );
  DFF_X1 key_c_r_reg_16_48 (.CK( clk ) , .D( key_c_r_15_48 ) , .Q( key_c_r_16_48 ) );
  DFF_X1 key_c_r_reg_16_49 (.CK( clk ) , .D( key_c_r_15_49 ) , .Q( key_c_r_16_49 ) );
  DFF_X1 key_c_r_reg_16_5 (.CK( clk ) , .D( key_c_r_15_5 ) , .Q( key_c_r_16_5 ) );
  DFF_X1 key_c_r_reg_16_50 (.CK( clk ) , .D( key_c_r_15_50 ) , .Q( key_c_r_16_50 ) );
  DFF_X1 key_c_r_reg_16_51 (.CK( clk ) , .D( key_c_r_15_51 ) , .Q( key_c_r_16_51 ) );
  DFF_X1 key_c_r_reg_16_52 (.CK( clk ) , .D( key_c_r_15_52 ) , .Q( key_c_r_16_52 ) );
  DFF_X1 key_c_r_reg_16_53 (.CK( clk ) , .D( key_c_r_15_53 ) , .Q( key_c_r_16_53 ) );
  DFF_X1 key_c_r_reg_16_54 (.CK( clk ) , .D( key_c_r_15_54 ) , .Q( key_c_r_16_54 ) );
  DFF_X1 key_c_r_reg_16_55 (.CK( clk ) , .D( key_c_r_15_55 ) , .Q( key_c_r_16_55 ) );
  DFF_X1 key_c_r_reg_16_6 (.CK( clk ) , .D( key_c_r_15_6 ) , .Q( key_c_r_16_6 ) );
  DFF_X1 key_c_r_reg_16_7 (.CK( clk ) , .D( key_c_r_15_7 ) , .Q( key_c_r_16_7 ) );
  DFF_X1 key_c_r_reg_16_8 (.CK( clk ) , .D( key_c_r_15_8 ) , .Q( key_c_r_16_8 ) );
  DFF_X1 key_c_r_reg_16_9 (.CK( clk ) , .D( key_c_r_15_9 ) , .Q( key_c_r_16_9 ) );
  DFF_X1 key_c_r_reg_17_0 (.CK( clk ) , .D( key_c_r_16_0 ) , .Q( key_c_r_17_0 ) );
  DFF_X1 key_c_r_reg_17_1 (.CK( clk ) , .D( key_c_r_16_1 ) , .Q( key_c_r_17_1 ) );
  DFF_X1 key_c_r_reg_17_10 (.CK( clk ) , .D( key_c_r_16_10 ) , .Q( key_c_r_17_10 ) );
  DFF_X1 key_c_r_reg_17_11 (.CK( clk ) , .D( key_c_r_16_11 ) , .Q( key_c_r_17_11 ) );
  DFF_X1 key_c_r_reg_17_12 (.CK( clk ) , .D( key_c_r_16_12 ) , .Q( key_c_r_17_12 ) );
  DFF_X1 key_c_r_reg_17_13 (.CK( clk ) , .D( key_c_r_16_13 ) , .Q( key_c_r_17_13 ) );
  DFF_X1 key_c_r_reg_17_14 (.CK( clk ) , .D( key_c_r_16_14 ) , .Q( key_c_r_17_14 ) );
  DFF_X1 key_c_r_reg_17_15 (.CK( clk ) , .D( key_c_r_16_15 ) , .Q( key_c_r_17_15 ) );
  DFF_X1 key_c_r_reg_17_16 (.CK( clk ) , .D( key_c_r_16_16 ) , .Q( key_c_r_17_16 ) );
  DFF_X1 key_c_r_reg_17_17 (.CK( clk ) , .D( key_c_r_16_17 ) , .Q( key_c_r_17_17 ) );
  DFF_X1 key_c_r_reg_17_18 (.CK( clk ) , .D( key_c_r_16_18 ) , .Q( key_c_r_17_18 ) );
  DFF_X1 key_c_r_reg_17_19 (.CK( clk ) , .D( key_c_r_16_19 ) , .Q( key_c_r_17_19 ) );
  DFF_X1 key_c_r_reg_17_2 (.CK( clk ) , .D( key_c_r_16_2 ) , .Q( key_c_r_17_2 ) );
  DFF_X1 key_c_r_reg_17_20 (.CK( clk ) , .D( key_c_r_16_20 ) , .Q( key_c_r_17_20 ) );
  DFF_X1 key_c_r_reg_17_21 (.CK( clk ) , .D( key_c_r_16_21 ) , .Q( key_c_r_17_21 ) );
  DFF_X1 key_c_r_reg_17_22 (.CK( clk ) , .D( key_c_r_16_22 ) , .Q( key_c_r_17_22 ) );
  DFF_X1 key_c_r_reg_17_23 (.CK( clk ) , .D( key_c_r_16_23 ) , .Q( key_c_r_17_23 ) );
  DFF_X1 key_c_r_reg_17_24 (.CK( clk ) , .D( key_c_r_16_24 ) , .Q( key_c_r_17_24 ) );
  DFF_X1 key_c_r_reg_17_25 (.CK( clk ) , .D( key_c_r_16_25 ) , .Q( key_c_r_17_25 ) );
  DFF_X1 key_c_r_reg_17_26 (.CK( clk ) , .D( key_c_r_16_26 ) , .Q( key_c_r_17_26 ) );
  DFF_X1 key_c_r_reg_17_27 (.CK( clk ) , .D( key_c_r_16_27 ) , .Q( key_c_r_17_27 ) );
  DFF_X1 key_c_r_reg_17_28 (.CK( clk ) , .D( key_c_r_16_28 ) , .Q( key_c_r_17_28 ) );
  DFF_X1 key_c_r_reg_17_29 (.CK( clk ) , .D( key_c_r_16_29 ) , .Q( key_c_r_17_29 ) );
  DFF_X1 key_c_r_reg_17_3 (.CK( clk ) , .D( key_c_r_16_3 ) , .Q( key_c_r_17_3 ) );
  DFF_X1 key_c_r_reg_17_30 (.CK( clk ) , .D( key_c_r_16_30 ) , .Q( key_c_r_17_30 ) );
  DFF_X1 key_c_r_reg_17_31 (.CK( clk ) , .D( key_c_r_16_31 ) , .Q( key_c_r_17_31 ) );
  DFF_X1 key_c_r_reg_17_32 (.CK( clk ) , .D( key_c_r_16_32 ) , .Q( key_c_r_17_32 ) );
  DFF_X1 key_c_r_reg_17_33 (.CK( clk ) , .D( key_c_r_16_33 ) , .Q( key_c_r_17_33 ) );
  DFF_X1 key_c_r_reg_17_34 (.CK( clk ) , .D( key_c_r_16_34 ) , .Q( key_c_r_17_34 ) );
  DFF_X1 key_c_r_reg_17_35 (.CK( clk ) , .D( key_c_r_16_35 ) , .Q( key_c_r_17_35 ) );
  DFF_X1 key_c_r_reg_17_36 (.CK( clk ) , .D( key_c_r_16_36 ) , .Q( key_c_r_17_36 ) );
  DFF_X1 key_c_r_reg_17_37 (.CK( clk ) , .D( key_c_r_16_37 ) , .Q( key_c_r_17_37 ) );
  DFF_X1 key_c_r_reg_17_38 (.CK( clk ) , .D( key_c_r_16_38 ) , .Q( key_c_r_17_38 ) );
  DFF_X1 key_c_r_reg_17_39 (.CK( clk ) , .D( key_c_r_16_39 ) , .Q( key_c_r_17_39 ) );
  DFF_X1 key_c_r_reg_17_4 (.CK( clk ) , .D( key_c_r_16_4 ) , .Q( key_c_r_17_4 ) );
  DFF_X1 key_c_r_reg_17_40 (.CK( clk ) , .D( key_c_r_16_40 ) , .Q( key_c_r_17_40 ) );
  DFF_X1 key_c_r_reg_17_41 (.CK( clk ) , .D( key_c_r_16_41 ) , .Q( key_c_r_17_41 ) );
  DFF_X1 key_c_r_reg_17_42 (.CK( clk ) , .D( key_c_r_16_42 ) , .Q( key_c_r_17_42 ) );
  DFF_X1 key_c_r_reg_17_43 (.CK( clk ) , .D( key_c_r_16_43 ) , .Q( key_c_r_17_43 ) );
  DFF_X1 key_c_r_reg_17_44 (.CK( clk ) , .D( key_c_r_16_44 ) , .Q( key_c_r_17_44 ) );
  DFF_X1 key_c_r_reg_17_45 (.CK( clk ) , .D( key_c_r_16_45 ) , .Q( key_c_r_17_45 ) );
  DFF_X1 key_c_r_reg_17_46 (.CK( clk ) , .D( key_c_r_16_46 ) , .Q( key_c_r_17_46 ) );
  DFF_X1 key_c_r_reg_17_47 (.CK( clk ) , .D( key_c_r_16_47 ) , .Q( key_c_r_17_47 ) );
  DFF_X1 key_c_r_reg_17_48 (.CK( clk ) , .D( key_c_r_16_48 ) , .Q( key_c_r_17_48 ) );
  DFF_X1 key_c_r_reg_17_49 (.CK( clk ) , .D( key_c_r_16_49 ) , .Q( key_c_r_17_49 ) );
  DFF_X1 key_c_r_reg_17_5 (.CK( clk ) , .D( key_c_r_16_5 ) , .Q( key_c_r_17_5 ) );
  DFF_X1 key_c_r_reg_17_50 (.CK( clk ) , .D( key_c_r_16_50 ) , .Q( key_c_r_17_50 ) );
  DFF_X1 key_c_r_reg_17_51 (.CK( clk ) , .D( key_c_r_16_51 ) , .Q( key_c_r_17_51 ) );
  DFF_X1 key_c_r_reg_17_52 (.CK( clk ) , .D( key_c_r_16_52 ) , .Q( key_c_r_17_52 ) );
  DFF_X1 key_c_r_reg_17_53 (.CK( clk ) , .D( key_c_r_16_53 ) , .Q( key_c_r_17_53 ) );
  DFF_X1 key_c_r_reg_17_54 (.CK( clk ) , .D( key_c_r_16_54 ) , .Q( key_c_r_17_54 ) );
  DFF_X1 key_c_r_reg_17_55 (.CK( clk ) , .D( key_c_r_16_55 ) , .Q( key_c_r_17_55 ) );
  DFF_X1 key_c_r_reg_17_6 (.CK( clk ) , .D( key_c_r_16_6 ) , .Q( key_c_r_17_6 ) );
  DFF_X1 key_c_r_reg_17_7 (.CK( clk ) , .D( key_c_r_16_7 ) , .Q( key_c_r_17_7 ) );
  DFF_X1 key_c_r_reg_17_8 (.CK( clk ) , .D( key_c_r_16_8 ) , .Q( key_c_r_17_8 ) );
  DFF_X1 key_c_r_reg_17_9 (.CK( clk ) , .D( key_c_r_16_9 ) , .Q( key_c_r_17_9 ) );
  DFF_X1 key_c_r_reg_18_0 (.CK( clk ) , .D( key_c_r_17_0 ) , .Q( key_c_r_18_0 ) );
  DFF_X1 key_c_r_reg_18_1 (.CK( clk ) , .D( key_c_r_17_1 ) , .Q( key_c_r_18_1 ) );
  DFF_X1 key_c_r_reg_18_10 (.CK( clk ) , .D( key_c_r_17_10 ) , .Q( key_c_r_18_10 ) );
  DFF_X1 key_c_r_reg_18_11 (.CK( clk ) , .D( key_c_r_17_11 ) , .Q( key_c_r_18_11 ) );
  DFF_X1 key_c_r_reg_18_12 (.CK( clk ) , .D( key_c_r_17_12 ) , .Q( key_c_r_18_12 ) );
  DFF_X1 key_c_r_reg_18_13 (.CK( clk ) , .D( key_c_r_17_13 ) , .Q( key_c_r_18_13 ) );
  DFF_X1 key_c_r_reg_18_14 (.CK( clk ) , .D( key_c_r_17_14 ) , .Q( key_c_r_18_14 ) );
  DFF_X1 key_c_r_reg_18_15 (.CK( clk ) , .D( key_c_r_17_15 ) , .Q( key_c_r_18_15 ) );
  DFF_X1 key_c_r_reg_18_16 (.CK( clk ) , .D( key_c_r_17_16 ) , .Q( key_c_r_18_16 ) );
  DFF_X1 key_c_r_reg_18_17 (.CK( clk ) , .D( key_c_r_17_17 ) , .Q( key_c_r_18_17 ) );
  DFF_X1 key_c_r_reg_18_18 (.CK( clk ) , .D( key_c_r_17_18 ) , .Q( key_c_r_18_18 ) );
  DFF_X1 key_c_r_reg_18_19 (.CK( clk ) , .D( key_c_r_17_19 ) , .Q( key_c_r_18_19 ) );
  DFF_X1 key_c_r_reg_18_2 (.CK( clk ) , .D( key_c_r_17_2 ) , .Q( key_c_r_18_2 ) );
  DFF_X1 key_c_r_reg_18_20 (.CK( clk ) , .D( key_c_r_17_20 ) , .Q( key_c_r_18_20 ) );
  DFF_X1 key_c_r_reg_18_21 (.CK( clk ) , .D( key_c_r_17_21 ) , .Q( key_c_r_18_21 ) );
  DFF_X1 key_c_r_reg_18_22 (.CK( clk ) , .D( key_c_r_17_22 ) , .Q( key_c_r_18_22 ) );
  DFF_X1 key_c_r_reg_18_23 (.CK( clk ) , .D( key_c_r_17_23 ) , .Q( key_c_r_18_23 ) );
  DFF_X1 key_c_r_reg_18_24 (.CK( clk ) , .D( key_c_r_17_24 ) , .Q( key_c_r_18_24 ) );
  DFF_X1 key_c_r_reg_18_25 (.CK( clk ) , .D( key_c_r_17_25 ) , .Q( key_c_r_18_25 ) );
  DFF_X1 key_c_r_reg_18_26 (.CK( clk ) , .D( key_c_r_17_26 ) , .Q( key_c_r_18_26 ) );
  DFF_X1 key_c_r_reg_18_27 (.CK( clk ) , .D( key_c_r_17_27 ) , .Q( key_c_r_18_27 ) );
  DFF_X1 key_c_r_reg_18_28 (.CK( clk ) , .D( key_c_r_17_28 ) , .Q( key_c_r_18_28 ) );
  DFF_X1 key_c_r_reg_18_29 (.CK( clk ) , .D( key_c_r_17_29 ) , .Q( key_c_r_18_29 ) );
  DFF_X1 key_c_r_reg_18_3 (.CK( clk ) , .D( key_c_r_17_3 ) , .Q( key_c_r_18_3 ) );
  DFF_X1 key_c_r_reg_18_30 (.CK( clk ) , .D( key_c_r_17_30 ) , .Q( key_c_r_18_30 ) );
  DFF_X1 key_c_r_reg_18_31 (.CK( clk ) , .D( key_c_r_17_31 ) , .Q( key_c_r_18_31 ) );
  DFF_X1 key_c_r_reg_18_32 (.CK( clk ) , .D( key_c_r_17_32 ) , .Q( key_c_r_18_32 ) );
  DFF_X1 key_c_r_reg_18_33 (.CK( clk ) , .D( key_c_r_17_33 ) , .Q( key_c_r_18_33 ) );
  DFF_X1 key_c_r_reg_18_34 (.CK( clk ) , .D( key_c_r_17_34 ) , .Q( key_c_r_18_34 ) );
  DFF_X1 key_c_r_reg_18_35 (.CK( clk ) , .D( key_c_r_17_35 ) , .Q( key_c_r_18_35 ) );
  DFF_X1 key_c_r_reg_18_36 (.CK( clk ) , .D( key_c_r_17_36 ) , .Q( key_c_r_18_36 ) );
  DFF_X1 key_c_r_reg_18_37 (.CK( clk ) , .D( key_c_r_17_37 ) , .Q( key_c_r_18_37 ) );
  DFF_X1 key_c_r_reg_18_38 (.CK( clk ) , .D( key_c_r_17_38 ) , .Q( key_c_r_18_38 ) );
  DFF_X1 key_c_r_reg_18_39 (.CK( clk ) , .D( key_c_r_17_39 ) , .Q( key_c_r_18_39 ) );
  DFF_X1 key_c_r_reg_18_4 (.CK( clk ) , .D( key_c_r_17_4 ) , .Q( key_c_r_18_4 ) );
  DFF_X1 key_c_r_reg_18_40 (.CK( clk ) , .D( key_c_r_17_40 ) , .Q( key_c_r_18_40 ) );
  DFF_X1 key_c_r_reg_18_41 (.CK( clk ) , .D( key_c_r_17_41 ) , .Q( key_c_r_18_41 ) );
  DFF_X1 key_c_r_reg_18_42 (.CK( clk ) , .D( key_c_r_17_42 ) , .Q( key_c_r_18_42 ) );
  DFF_X1 key_c_r_reg_18_43 (.CK( clk ) , .D( key_c_r_17_43 ) , .Q( key_c_r_18_43 ) );
  DFF_X1 key_c_r_reg_18_44 (.CK( clk ) , .D( key_c_r_17_44 ) , .Q( key_c_r_18_44 ) );
  DFF_X1 key_c_r_reg_18_45 (.CK( clk ) , .D( key_c_r_17_45 ) , .Q( key_c_r_18_45 ) );
  DFF_X1 key_c_r_reg_18_46 (.CK( clk ) , .D( key_c_r_17_46 ) , .Q( key_c_r_18_46 ) );
  DFF_X1 key_c_r_reg_18_47 (.CK( clk ) , .D( key_c_r_17_47 ) , .Q( key_c_r_18_47 ) );
  DFF_X1 key_c_r_reg_18_48 (.CK( clk ) , .D( key_c_r_17_48 ) , .Q( key_c_r_18_48 ) );
  DFF_X1 key_c_r_reg_18_49 (.CK( clk ) , .D( key_c_r_17_49 ) , .Q( key_c_r_18_49 ) );
  DFF_X1 key_c_r_reg_18_5 (.CK( clk ) , .D( key_c_r_17_5 ) , .Q( key_c_r_18_5 ) );
  DFF_X1 key_c_r_reg_18_50 (.CK( clk ) , .D( key_c_r_17_50 ) , .Q( key_c_r_18_50 ) );
  DFF_X1 key_c_r_reg_18_51 (.CK( clk ) , .D( key_c_r_17_51 ) , .Q( key_c_r_18_51 ) );
  DFF_X1 key_c_r_reg_18_52 (.CK( clk ) , .D( key_c_r_17_52 ) , .Q( key_c_r_18_52 ) );
  DFF_X1 key_c_r_reg_18_53 (.CK( clk ) , .D( key_c_r_17_53 ) , .Q( key_c_r_18_53 ) );
  DFF_X1 key_c_r_reg_18_54 (.CK( clk ) , .D( key_c_r_17_54 ) , .Q( key_c_r_18_54 ) );
  DFF_X1 key_c_r_reg_18_55 (.CK( clk ) , .D( key_c_r_17_55 ) , .Q( key_c_r_18_55 ) );
  DFF_X1 key_c_r_reg_18_6 (.CK( clk ) , .D( key_c_r_17_6 ) , .Q( key_c_r_18_6 ) );
  DFF_X1 key_c_r_reg_18_7 (.CK( clk ) , .D( key_c_r_17_7 ) , .Q( key_c_r_18_7 ) );
  DFF_X1 key_c_r_reg_18_8 (.CK( clk ) , .D( key_c_r_17_8 ) , .Q( key_c_r_18_8 ) );
  DFF_X1 key_c_r_reg_18_9 (.CK( clk ) , .D( key_c_r_17_9 ) , .Q( key_c_r_18_9 ) );
  DFF_X1 key_c_r_reg_19_0 (.CK( clk ) , .D( key_c_r_18_0 ) , .Q( key_c_r_19_0 ) );
  DFF_X1 key_c_r_reg_19_1 (.CK( clk ) , .D( key_c_r_18_1 ) , .Q( key_c_r_19_1 ) );
  DFF_X1 key_c_r_reg_19_10 (.CK( clk ) , .D( key_c_r_18_10 ) , .Q( key_c_r_19_10 ) );
  DFF_X1 key_c_r_reg_19_11 (.CK( clk ) , .D( key_c_r_18_11 ) , .Q( key_c_r_19_11 ) );
  DFF_X1 key_c_r_reg_19_12 (.CK( clk ) , .D( key_c_r_18_12 ) , .Q( key_c_r_19_12 ) );
  DFF_X1 key_c_r_reg_19_13 (.CK( clk ) , .D( key_c_r_18_13 ) , .Q( key_c_r_19_13 ) );
  DFF_X1 key_c_r_reg_19_14 (.CK( clk ) , .D( key_c_r_18_14 ) , .Q( key_c_r_19_14 ) );
  DFF_X1 key_c_r_reg_19_15 (.CK( clk ) , .D( key_c_r_18_15 ) , .Q( key_c_r_19_15 ) );
  DFF_X1 key_c_r_reg_19_16 (.CK( clk ) , .D( key_c_r_18_16 ) , .Q( key_c_r_19_16 ) );
  DFF_X1 key_c_r_reg_19_17 (.CK( clk ) , .D( key_c_r_18_17 ) , .Q( key_c_r_19_17 ) );
  DFF_X1 key_c_r_reg_19_18 (.CK( clk ) , .D( key_c_r_18_18 ) , .Q( key_c_r_19_18 ) );
  DFF_X1 key_c_r_reg_19_19 (.CK( clk ) , .D( key_c_r_18_19 ) , .Q( key_c_r_19_19 ) );
  DFF_X1 key_c_r_reg_19_2 (.CK( clk ) , .D( key_c_r_18_2 ) , .Q( key_c_r_19_2 ) );
  DFF_X1 key_c_r_reg_19_20 (.CK( clk ) , .D( key_c_r_18_20 ) , .Q( key_c_r_19_20 ) );
  DFF_X1 key_c_r_reg_19_21 (.CK( clk ) , .D( key_c_r_18_21 ) , .Q( key_c_r_19_21 ) );
  DFF_X1 key_c_r_reg_19_22 (.CK( clk ) , .D( key_c_r_18_22 ) , .Q( key_c_r_19_22 ) );
  DFF_X1 key_c_r_reg_19_23 (.CK( clk ) , .D( key_c_r_18_23 ) , .Q( key_c_r_19_23 ) );
  DFF_X1 key_c_r_reg_19_24 (.CK( clk ) , .D( key_c_r_18_24 ) , .Q( key_c_r_19_24 ) );
  DFF_X1 key_c_r_reg_19_25 (.CK( clk ) , .D( key_c_r_18_25 ) , .Q( key_c_r_19_25 ) );
  DFF_X1 key_c_r_reg_19_26 (.CK( clk ) , .D( key_c_r_18_26 ) , .Q( key_c_r_19_26 ) );
  DFF_X1 key_c_r_reg_19_27 (.CK( clk ) , .D( key_c_r_18_27 ) , .Q( key_c_r_19_27 ) );
  DFF_X1 key_c_r_reg_19_28 (.CK( clk ) , .D( key_c_r_18_28 ) , .Q( key_c_r_19_28 ) );
  DFF_X1 key_c_r_reg_19_29 (.CK( clk ) , .D( key_c_r_18_29 ) , .Q( key_c_r_19_29 ) );
  DFF_X1 key_c_r_reg_19_3 (.CK( clk ) , .D( key_c_r_18_3 ) , .Q( key_c_r_19_3 ) );
  DFF_X1 key_c_r_reg_19_30 (.CK( clk ) , .D( key_c_r_18_30 ) , .Q( key_c_r_19_30 ) );
  DFF_X1 key_c_r_reg_19_31 (.CK( clk ) , .D( key_c_r_18_31 ) , .Q( key_c_r_19_31 ) );
  DFF_X1 key_c_r_reg_19_32 (.CK( clk ) , .D( key_c_r_18_32 ) , .Q( key_c_r_19_32 ) );
  DFF_X1 key_c_r_reg_19_33 (.CK( clk ) , .D( key_c_r_18_33 ) , .Q( key_c_r_19_33 ) );
  DFF_X1 key_c_r_reg_19_34 (.CK( clk ) , .D( key_c_r_18_34 ) , .Q( key_c_r_19_34 ) );
  DFF_X1 key_c_r_reg_19_35 (.CK( clk ) , .D( key_c_r_18_35 ) , .Q( key_c_r_19_35 ) );
  DFF_X1 key_c_r_reg_19_36 (.CK( clk ) , .D( key_c_r_18_36 ) , .Q( key_c_r_19_36 ) );
  DFF_X1 key_c_r_reg_19_37 (.CK( clk ) , .D( key_c_r_18_37 ) , .Q( key_c_r_19_37 ) );
  DFF_X1 key_c_r_reg_19_38 (.CK( clk ) , .D( key_c_r_18_38 ) , .Q( key_c_r_19_38 ) );
  DFF_X1 key_c_r_reg_19_39 (.CK( clk ) , .D( key_c_r_18_39 ) , .Q( key_c_r_19_39 ) );
  DFF_X1 key_c_r_reg_19_4 (.CK( clk ) , .D( key_c_r_18_4 ) , .Q( key_c_r_19_4 ) );
  DFF_X1 key_c_r_reg_19_40 (.CK( clk ) , .D( key_c_r_18_40 ) , .Q( key_c_r_19_40 ) );
  DFF_X1 key_c_r_reg_19_41 (.CK( clk ) , .D( key_c_r_18_41 ) , .Q( key_c_r_19_41 ) );
  DFF_X1 key_c_r_reg_19_42 (.CK( clk ) , .D( key_c_r_18_42 ) , .Q( key_c_r_19_42 ) );
  DFF_X1 key_c_r_reg_19_43 (.CK( clk ) , .D( key_c_r_18_43 ) , .Q( key_c_r_19_43 ) );
  DFF_X1 key_c_r_reg_19_44 (.CK( clk ) , .D( key_c_r_18_44 ) , .Q( key_c_r_19_44 ) );
  DFF_X1 key_c_r_reg_19_45 (.CK( clk ) , .D( key_c_r_18_45 ) , .Q( key_c_r_19_45 ) );
  DFF_X1 key_c_r_reg_19_46 (.CK( clk ) , .D( key_c_r_18_46 ) , .Q( key_c_r_19_46 ) );
  DFF_X1 key_c_r_reg_19_47 (.CK( clk ) , .D( key_c_r_18_47 ) , .Q( key_c_r_19_47 ) );
  DFF_X1 key_c_r_reg_19_48 (.CK( clk ) , .D( key_c_r_18_48 ) , .Q( key_c_r_19_48 ) );
  DFF_X1 key_c_r_reg_19_49 (.CK( clk ) , .D( key_c_r_18_49 ) , .Q( key_c_r_19_49 ) );
  DFF_X1 key_c_r_reg_19_5 (.CK( clk ) , .D( key_c_r_18_5 ) , .Q( key_c_r_19_5 ) );
  DFF_X1 key_c_r_reg_19_50 (.CK( clk ) , .D( key_c_r_18_50 ) , .Q( key_c_r_19_50 ) );
  DFF_X1 key_c_r_reg_19_51 (.CK( clk ) , .D( key_c_r_18_51 ) , .Q( key_c_r_19_51 ) );
  DFF_X1 key_c_r_reg_19_52 (.CK( clk ) , .D( key_c_r_18_52 ) , .Q( key_c_r_19_52 ) );
  DFF_X1 key_c_r_reg_19_53 (.CK( clk ) , .D( key_c_r_18_53 ) , .Q( key_c_r_19_53 ) );
  DFF_X1 key_c_r_reg_19_54 (.CK( clk ) , .D( key_c_r_18_54 ) , .Q( key_c_r_19_54 ) );
  DFF_X1 key_c_r_reg_19_55 (.CK( clk ) , .D( key_c_r_18_55 ) , .Q( key_c_r_19_55 ) );
  DFF_X1 key_c_r_reg_19_6 (.CK( clk ) , .D( key_c_r_18_6 ) , .Q( key_c_r_19_6 ) );
  DFF_X1 key_c_r_reg_19_7 (.CK( clk ) , .D( key_c_r_18_7 ) , .Q( key_c_r_19_7 ) );
  DFF_X1 key_c_r_reg_19_8 (.CK( clk ) , .D( key_c_r_18_8 ) , .Q( key_c_r_19_8 ) );
  DFF_X1 key_c_r_reg_19_9 (.CK( clk ) , .D( key_c_r_18_9 ) , .Q( key_c_r_19_9 ) );
  DFF_X1 key_c_r_reg_1_0 (.CK( clk ) , .D( key_c_r_0_0 ) , .Q( key_c_r_1_0 ) );
  DFF_X1 key_c_r_reg_1_1 (.CK( clk ) , .D( key_c_r_0_1 ) , .Q( key_c_r_1_1 ) );
  DFF_X1 key_c_r_reg_1_10 (.CK( clk ) , .D( key_c_r_0_10 ) , .Q( key_c_r_1_10 ) );
  DFF_X1 key_c_r_reg_1_11 (.CK( clk ) , .D( key_c_r_0_11 ) , .Q( key_c_r_1_11 ) );
  DFF_X1 key_c_r_reg_1_12 (.CK( clk ) , .D( key_c_r_0_12 ) , .Q( key_c_r_1_12 ) );
  DFF_X1 key_c_r_reg_1_13 (.CK( clk ) , .D( key_c_r_0_13 ) , .Q( key_c_r_1_13 ) );
  DFF_X1 key_c_r_reg_1_14 (.CK( clk ) , .D( key_c_r_0_14 ) , .Q( key_c_r_1_14 ) );
  DFF_X1 key_c_r_reg_1_15 (.CK( clk ) , .D( key_c_r_0_15 ) , .Q( key_c_r_1_15 ) );
  DFF_X1 key_c_r_reg_1_16 (.CK( clk ) , .D( key_c_r_0_16 ) , .Q( key_c_r_1_16 ) );
  DFF_X1 key_c_r_reg_1_17 (.CK( clk ) , .D( key_c_r_0_17 ) , .Q( key_c_r_1_17 ) );
  DFF_X1 key_c_r_reg_1_18 (.CK( clk ) , .D( key_c_r_0_18 ) , .Q( key_c_r_1_18 ) );
  DFF_X1 key_c_r_reg_1_19 (.CK( clk ) , .D( key_c_r_0_19 ) , .Q( key_c_r_1_19 ) );
  DFF_X1 key_c_r_reg_1_2 (.CK( clk ) , .D( key_c_r_0_2 ) , .Q( key_c_r_1_2 ) );
  DFF_X1 key_c_r_reg_1_20 (.CK( clk ) , .D( key_c_r_0_20 ) , .Q( key_c_r_1_20 ) );
  DFF_X1 key_c_r_reg_1_21 (.CK( clk ) , .D( key_c_r_0_21 ) , .Q( key_c_r_1_21 ) );
  DFF_X1 key_c_r_reg_1_22 (.CK( clk ) , .D( key_c_r_0_22 ) , .Q( key_c_r_1_22 ) );
  DFF_X1 key_c_r_reg_1_23 (.CK( clk ) , .D( key_c_r_0_23 ) , .Q( key_c_r_1_23 ) );
  DFF_X1 key_c_r_reg_1_24 (.CK( clk ) , .D( key_c_r_0_24 ) , .Q( key_c_r_1_24 ) );
  DFF_X1 key_c_r_reg_1_25 (.CK( clk ) , .D( key_c_r_0_25 ) , .Q( key_c_r_1_25 ) );
  DFF_X1 key_c_r_reg_1_26 (.CK( clk ) , .D( key_c_r_0_26 ) , .Q( key_c_r_1_26 ) );
  DFF_X1 key_c_r_reg_1_27 (.CK( clk ) , .D( key_c_r_0_27 ) , .Q( key_c_r_1_27 ) );
  DFF_X1 key_c_r_reg_1_28 (.CK( clk ) , .D( key_c_r_0_28 ) , .Q( key_c_r_1_28 ) );
  DFF_X1 key_c_r_reg_1_29 (.CK( clk ) , .D( key_c_r_0_29 ) , .Q( key_c_r_1_29 ) );
  DFF_X1 key_c_r_reg_1_3 (.CK( clk ) , .D( key_c_r_0_3 ) , .Q( key_c_r_1_3 ) );
  DFF_X1 key_c_r_reg_1_30 (.CK( clk ) , .D( key_c_r_0_30 ) , .Q( key_c_r_1_30 ) );
  DFF_X1 key_c_r_reg_1_31 (.CK( clk ) , .D( key_c_r_0_31 ) , .Q( key_c_r_1_31 ) );
  DFF_X1 key_c_r_reg_1_32 (.CK( clk ) , .D( key_c_r_0_32 ) , .Q( key_c_r_1_32 ) );
  DFF_X1 key_c_r_reg_1_33 (.CK( clk ) , .D( key_c_r_0_33 ) , .Q( key_c_r_1_33 ) );
  DFF_X1 key_c_r_reg_1_34 (.CK( clk ) , .D( key_c_r_0_34 ) , .Q( key_c_r_1_34 ) );
  DFF_X1 key_c_r_reg_1_35 (.CK( clk ) , .D( key_c_r_0_35 ) , .Q( key_c_r_1_35 ) );
  DFF_X1 key_c_r_reg_1_36 (.CK( clk ) , .D( key_c_r_0_36 ) , .Q( key_c_r_1_36 ) );
  DFF_X1 key_c_r_reg_1_37 (.CK( clk ) , .D( key_c_r_0_37 ) , .Q( key_c_r_1_37 ) );
  DFF_X1 key_c_r_reg_1_38 (.CK( clk ) , .D( key_c_r_0_38 ) , .Q( key_c_r_1_38 ) );
  DFF_X1 key_c_r_reg_1_39 (.CK( clk ) , .D( key_c_r_0_39 ) , .Q( key_c_r_1_39 ) );
  DFF_X1 key_c_r_reg_1_4 (.CK( clk ) , .D( key_c_r_0_4 ) , .Q( key_c_r_1_4 ) );
  DFF_X1 key_c_r_reg_1_40 (.CK( clk ) , .D( key_c_r_0_40 ) , .Q( key_c_r_1_40 ) );
  DFF_X1 key_c_r_reg_1_41 (.CK( clk ) , .D( key_c_r_0_41 ) , .Q( key_c_r_1_41 ) );
  DFF_X1 key_c_r_reg_1_42 (.CK( clk ) , .D( key_c_r_0_42 ) , .Q( key_c_r_1_42 ) );
  DFF_X1 key_c_r_reg_1_43 (.CK( clk ) , .D( key_c_r_0_43 ) , .Q( key_c_r_1_43 ) );
  DFF_X1 key_c_r_reg_1_44 (.CK( clk ) , .D( key_c_r_0_44 ) , .Q( key_c_r_1_44 ) );
  DFF_X1 key_c_r_reg_1_45 (.CK( clk ) , .D( key_c_r_0_45 ) , .Q( key_c_r_1_45 ) );
  DFF_X1 key_c_r_reg_1_46 (.CK( clk ) , .D( key_c_r_0_46 ) , .Q( key_c_r_1_46 ) );
  DFF_X1 key_c_r_reg_1_47 (.CK( clk ) , .D( key_c_r_0_47 ) , .Q( key_c_r_1_47 ) );
  DFF_X1 key_c_r_reg_1_48 (.CK( clk ) , .D( key_c_r_0_48 ) , .Q( key_c_r_1_48 ) );
  DFF_X1 key_c_r_reg_1_49 (.CK( clk ) , .D( key_c_r_0_49 ) , .Q( key_c_r_1_49 ) );
  DFF_X1 key_c_r_reg_1_5 (.CK( clk ) , .D( key_c_r_0_5 ) , .Q( key_c_r_1_5 ) );
  DFF_X1 key_c_r_reg_1_50 (.CK( clk ) , .D( key_c_r_0_50 ) , .Q( key_c_r_1_50 ) );
  DFF_X1 key_c_r_reg_1_51 (.CK( clk ) , .D( key_c_r_0_51 ) , .Q( key_c_r_1_51 ) );
  DFF_X1 key_c_r_reg_1_52 (.CK( clk ) , .D( key_c_r_0_52 ) , .Q( key_c_r_1_52 ) );
  DFF_X1 key_c_r_reg_1_53 (.CK( clk ) , .D( key_c_r_0_53 ) , .Q( key_c_r_1_53 ) );
  DFF_X1 key_c_r_reg_1_54 (.CK( clk ) , .D( key_c_r_0_54 ) , .Q( key_c_r_1_54 ) );
  DFF_X1 key_c_r_reg_1_55 (.CK( clk ) , .D( key_c_r_0_55 ) , .Q( key_c_r_1_55 ) );
  DFF_X1 key_c_r_reg_1_6 (.CK( clk ) , .D( key_c_r_0_6 ) , .Q( key_c_r_1_6 ) );
  DFF_X1 key_c_r_reg_1_7 (.CK( clk ) , .D( key_c_r_0_7 ) , .Q( key_c_r_1_7 ) );
  DFF_X1 key_c_r_reg_1_8 (.CK( clk ) , .D( key_c_r_0_8 ) , .Q( key_c_r_1_8 ) );
  DFF_X1 key_c_r_reg_1_9 (.CK( clk ) , .D( key_c_r_0_9 ) , .Q( key_c_r_1_9 ) );
  DFF_X1 key_c_r_reg_20_0 (.CK( clk ) , .D( key_c_r_19_0 ) , .Q( key_c_r_20_0 ) );
  DFF_X1 key_c_r_reg_20_1 (.CK( clk ) , .D( key_c_r_19_1 ) , .Q( key_c_r_20_1 ) );
  DFF_X1 key_c_r_reg_20_10 (.CK( clk ) , .D( key_c_r_19_10 ) , .Q( key_c_r_20_10 ) );
  DFF_X1 key_c_r_reg_20_11 (.CK( clk ) , .D( key_c_r_19_11 ) , .Q( key_c_r_20_11 ) );
  DFF_X1 key_c_r_reg_20_12 (.CK( clk ) , .D( key_c_r_19_12 ) , .Q( key_c_r_20_12 ) );
  DFF_X1 key_c_r_reg_20_13 (.CK( clk ) , .D( key_c_r_19_13 ) , .Q( key_c_r_20_13 ) );
  DFF_X1 key_c_r_reg_20_14 (.CK( clk ) , .D( key_c_r_19_14 ) , .Q( key_c_r_20_14 ) );
  DFF_X1 key_c_r_reg_20_15 (.CK( clk ) , .D( key_c_r_19_15 ) , .Q( key_c_r_20_15 ) );
  DFF_X1 key_c_r_reg_20_16 (.CK( clk ) , .D( key_c_r_19_16 ) , .Q( key_c_r_20_16 ) );
  DFF_X1 key_c_r_reg_20_17 (.CK( clk ) , .D( key_c_r_19_17 ) , .Q( key_c_r_20_17 ) );
  DFF_X1 key_c_r_reg_20_18 (.CK( clk ) , .D( key_c_r_19_18 ) , .Q( key_c_r_20_18 ) );
  DFF_X1 key_c_r_reg_20_19 (.CK( clk ) , .D( key_c_r_19_19 ) , .Q( key_c_r_20_19 ) );
  DFF_X1 key_c_r_reg_20_2 (.CK( clk ) , .D( key_c_r_19_2 ) , .Q( key_c_r_20_2 ) );
  DFF_X1 key_c_r_reg_20_20 (.CK( clk ) , .D( key_c_r_19_20 ) , .Q( key_c_r_20_20 ) );
  DFF_X1 key_c_r_reg_20_21 (.CK( clk ) , .D( key_c_r_19_21 ) , .Q( key_c_r_20_21 ) );
  DFF_X1 key_c_r_reg_20_22 (.CK( clk ) , .D( key_c_r_19_22 ) , .Q( key_c_r_20_22 ) );
  DFF_X1 key_c_r_reg_20_23 (.CK( clk ) , .D( key_c_r_19_23 ) , .Q( key_c_r_20_23 ) );
  DFF_X1 key_c_r_reg_20_24 (.CK( clk ) , .D( key_c_r_19_24 ) , .Q( key_c_r_20_24 ) );
  DFF_X1 key_c_r_reg_20_25 (.CK( clk ) , .D( key_c_r_19_25 ) , .Q( key_c_r_20_25 ) );
  DFF_X1 key_c_r_reg_20_26 (.CK( clk ) , .D( key_c_r_19_26 ) , .Q( key_c_r_20_26 ) );
  DFF_X1 key_c_r_reg_20_27 (.CK( clk ) , .D( key_c_r_19_27 ) , .Q( key_c_r_20_27 ) );
  DFF_X1 key_c_r_reg_20_28 (.CK( clk ) , .D( key_c_r_19_28 ) , .Q( key_c_r_20_28 ) );
  DFF_X1 key_c_r_reg_20_29 (.CK( clk ) , .D( key_c_r_19_29 ) , .Q( key_c_r_20_29 ) );
  DFF_X1 key_c_r_reg_20_3 (.CK( clk ) , .D( key_c_r_19_3 ) , .Q( key_c_r_20_3 ) );
  DFF_X1 key_c_r_reg_20_30 (.CK( clk ) , .D( key_c_r_19_30 ) , .Q( key_c_r_20_30 ) );
  DFF_X1 key_c_r_reg_20_31 (.CK( clk ) , .D( key_c_r_19_31 ) , .Q( key_c_r_20_31 ) );
  DFF_X1 key_c_r_reg_20_32 (.CK( clk ) , .D( key_c_r_19_32 ) , .Q( key_c_r_20_32 ) );
  DFF_X1 key_c_r_reg_20_33 (.CK( clk ) , .D( key_c_r_19_33 ) , .Q( key_c_r_20_33 ) );
  DFF_X1 key_c_r_reg_20_34 (.CK( clk ) , .D( key_c_r_19_34 ) , .Q( key_c_r_20_34 ) );
  DFF_X1 key_c_r_reg_20_35 (.CK( clk ) , .D( key_c_r_19_35 ) , .Q( key_c_r_20_35 ) );
  DFF_X1 key_c_r_reg_20_36 (.CK( clk ) , .D( key_c_r_19_36 ) , .Q( key_c_r_20_36 ) );
  DFF_X1 key_c_r_reg_20_37 (.CK( clk ) , .D( key_c_r_19_37 ) , .Q( key_c_r_20_37 ) );
  DFF_X1 key_c_r_reg_20_38 (.CK( clk ) , .D( key_c_r_19_38 ) , .Q( key_c_r_20_38 ) );
  DFF_X1 key_c_r_reg_20_39 (.CK( clk ) , .D( key_c_r_19_39 ) , .Q( key_c_r_20_39 ) );
  DFF_X1 key_c_r_reg_20_4 (.CK( clk ) , .D( key_c_r_19_4 ) , .Q( key_c_r_20_4 ) );
  DFF_X1 key_c_r_reg_20_40 (.CK( clk ) , .D( key_c_r_19_40 ) , .Q( key_c_r_20_40 ) );
  DFF_X1 key_c_r_reg_20_41 (.CK( clk ) , .D( key_c_r_19_41 ) , .Q( key_c_r_20_41 ) );
  DFF_X1 key_c_r_reg_20_42 (.CK( clk ) , .D( key_c_r_19_42 ) , .Q( key_c_r_20_42 ) );
  DFF_X1 key_c_r_reg_20_43 (.CK( clk ) , .D( key_c_r_19_43 ) , .Q( key_c_r_20_43 ) );
  DFF_X1 key_c_r_reg_20_44 (.CK( clk ) , .D( key_c_r_19_44 ) , .Q( key_c_r_20_44 ) );
  DFF_X1 key_c_r_reg_20_45 (.CK( clk ) , .D( key_c_r_19_45 ) , .Q( key_c_r_20_45 ) );
  DFF_X1 key_c_r_reg_20_46 (.CK( clk ) , .D( key_c_r_19_46 ) , .Q( key_c_r_20_46 ) );
  DFF_X1 key_c_r_reg_20_47 (.CK( clk ) , .D( key_c_r_19_47 ) , .Q( key_c_r_20_47 ) );
  DFF_X1 key_c_r_reg_20_48 (.CK( clk ) , .D( key_c_r_19_48 ) , .Q( key_c_r_20_48 ) );
  DFF_X1 key_c_r_reg_20_49 (.CK( clk ) , .D( key_c_r_19_49 ) , .Q( key_c_r_20_49 ) );
  DFF_X1 key_c_r_reg_20_5 (.CK( clk ) , .D( key_c_r_19_5 ) , .Q( key_c_r_20_5 ) );
  DFF_X1 key_c_r_reg_20_50 (.CK( clk ) , .D( key_c_r_19_50 ) , .Q( key_c_r_20_50 ) );
  DFF_X1 key_c_r_reg_20_51 (.CK( clk ) , .D( key_c_r_19_51 ) , .Q( key_c_r_20_51 ) );
  DFF_X1 key_c_r_reg_20_52 (.CK( clk ) , .D( key_c_r_19_52 ) , .Q( key_c_r_20_52 ) );
  DFF_X1 key_c_r_reg_20_53 (.CK( clk ) , .D( key_c_r_19_53 ) , .Q( key_c_r_20_53 ) );
  DFF_X1 key_c_r_reg_20_54 (.CK( clk ) , .D( key_c_r_19_54 ) , .Q( key_c_r_20_54 ) );
  DFF_X1 key_c_r_reg_20_55 (.CK( clk ) , .D( key_c_r_19_55 ) , .Q( key_c_r_20_55 ) );
  DFF_X1 key_c_r_reg_20_6 (.CK( clk ) , .D( key_c_r_19_6 ) , .Q( key_c_r_20_6 ) );
  DFF_X1 key_c_r_reg_20_7 (.CK( clk ) , .D( key_c_r_19_7 ) , .Q( key_c_r_20_7 ) );
  DFF_X1 key_c_r_reg_20_8 (.CK( clk ) , .D( key_c_r_19_8 ) , .Q( key_c_r_20_8 ) );
  DFF_X1 key_c_r_reg_20_9 (.CK( clk ) , .D( key_c_r_19_9 ) , .Q( key_c_r_20_9 ) );
  DFF_X1 key_c_r_reg_21_0 (.CK( clk ) , .D( key_c_r_20_0 ) , .Q( key_c_r_21_0 ) );
  DFF_X1 key_c_r_reg_21_1 (.CK( clk ) , .D( key_c_r_20_1 ) , .Q( key_c_r_21_1 ) );
  DFF_X1 key_c_r_reg_21_10 (.CK( clk ) , .D( key_c_r_20_10 ) , .Q( key_c_r_21_10 ) );
  DFF_X1 key_c_r_reg_21_11 (.CK( clk ) , .D( key_c_r_20_11 ) , .Q( key_c_r_21_11 ) );
  DFF_X1 key_c_r_reg_21_12 (.CK( clk ) , .D( key_c_r_20_12 ) , .Q( key_c_r_21_12 ) );
  DFF_X1 key_c_r_reg_21_13 (.CK( clk ) , .D( key_c_r_20_13 ) , .Q( key_c_r_21_13 ) );
  DFF_X1 key_c_r_reg_21_14 (.CK( clk ) , .D( key_c_r_20_14 ) , .Q( key_c_r_21_14 ) );
  DFF_X1 key_c_r_reg_21_15 (.CK( clk ) , .D( key_c_r_20_15 ) , .Q( key_c_r_21_15 ) );
  DFF_X1 key_c_r_reg_21_16 (.CK( clk ) , .D( key_c_r_20_16 ) , .Q( key_c_r_21_16 ) );
  DFF_X1 key_c_r_reg_21_17 (.CK( clk ) , .D( key_c_r_20_17 ) , .Q( key_c_r_21_17 ) );
  DFF_X1 key_c_r_reg_21_18 (.CK( clk ) , .D( key_c_r_20_18 ) , .Q( key_c_r_21_18 ) );
  DFF_X1 key_c_r_reg_21_19 (.CK( clk ) , .D( key_c_r_20_19 ) , .Q( key_c_r_21_19 ) );
  DFF_X1 key_c_r_reg_21_2 (.CK( clk ) , .D( key_c_r_20_2 ) , .Q( key_c_r_21_2 ) );
  DFF_X1 key_c_r_reg_21_20 (.CK( clk ) , .D( key_c_r_20_20 ) , .Q( key_c_r_21_20 ) );
  DFF_X1 key_c_r_reg_21_21 (.CK( clk ) , .D( key_c_r_20_21 ) , .Q( key_c_r_21_21 ) );
  DFF_X1 key_c_r_reg_21_22 (.CK( clk ) , .D( key_c_r_20_22 ) , .Q( key_c_r_21_22 ) );
  DFF_X1 key_c_r_reg_21_23 (.CK( clk ) , .D( key_c_r_20_23 ) , .Q( key_c_r_21_23 ) );
  DFF_X1 key_c_r_reg_21_24 (.CK( clk ) , .D( key_c_r_20_24 ) , .Q( key_c_r_21_24 ) );
  DFF_X1 key_c_r_reg_21_25 (.CK( clk ) , .D( key_c_r_20_25 ) , .Q( key_c_r_21_25 ) );
  DFF_X1 key_c_r_reg_21_26 (.CK( clk ) , .D( key_c_r_20_26 ) , .Q( key_c_r_21_26 ) );
  DFF_X1 key_c_r_reg_21_27 (.CK( clk ) , .D( key_c_r_20_27 ) , .Q( key_c_r_21_27 ) );
  DFF_X1 key_c_r_reg_21_28 (.CK( clk ) , .D( key_c_r_20_28 ) , .Q( key_c_r_21_28 ) );
  DFF_X1 key_c_r_reg_21_29 (.CK( clk ) , .D( key_c_r_20_29 ) , .Q( key_c_r_21_29 ) );
  DFF_X1 key_c_r_reg_21_3 (.CK( clk ) , .D( key_c_r_20_3 ) , .Q( key_c_r_21_3 ) );
  DFF_X1 key_c_r_reg_21_30 (.CK( clk ) , .D( key_c_r_20_30 ) , .Q( key_c_r_21_30 ) );
  DFF_X1 key_c_r_reg_21_31 (.CK( clk ) , .D( key_c_r_20_31 ) , .Q( key_c_r_21_31 ) );
  DFF_X1 key_c_r_reg_21_32 (.CK( clk ) , .D( key_c_r_20_32 ) , .Q( key_c_r_21_32 ) );
  DFF_X1 key_c_r_reg_21_33 (.CK( clk ) , .D( key_c_r_20_33 ) , .Q( key_c_r_21_33 ) );
  DFF_X1 key_c_r_reg_21_34 (.CK( clk ) , .D( key_c_r_20_34 ) , .Q( key_c_r_21_34 ) );
  DFF_X1 key_c_r_reg_21_35 (.CK( clk ) , .D( key_c_r_20_35 ) , .Q( key_c_r_21_35 ) );
  DFF_X1 key_c_r_reg_21_36 (.CK( clk ) , .D( key_c_r_20_36 ) , .Q( key_c_r_21_36 ) );
  DFF_X1 key_c_r_reg_21_37 (.CK( clk ) , .D( key_c_r_20_37 ) , .Q( key_c_r_21_37 ) );
  DFF_X1 key_c_r_reg_21_38 (.CK( clk ) , .D( key_c_r_20_38 ) , .Q( key_c_r_21_38 ) );
  DFF_X1 key_c_r_reg_21_39 (.CK( clk ) , .D( key_c_r_20_39 ) , .Q( key_c_r_21_39 ) );
  DFF_X1 key_c_r_reg_21_4 (.CK( clk ) , .D( key_c_r_20_4 ) , .Q( key_c_r_21_4 ) );
  DFF_X1 key_c_r_reg_21_40 (.CK( clk ) , .D( key_c_r_20_40 ) , .Q( key_c_r_21_40 ) );
  DFF_X1 key_c_r_reg_21_41 (.CK( clk ) , .D( key_c_r_20_41 ) , .Q( key_c_r_21_41 ) );
  DFF_X1 key_c_r_reg_21_42 (.CK( clk ) , .D( key_c_r_20_42 ) , .Q( key_c_r_21_42 ) );
  DFF_X1 key_c_r_reg_21_43 (.CK( clk ) , .D( key_c_r_20_43 ) , .Q( key_c_r_21_43 ) );
  DFF_X1 key_c_r_reg_21_44 (.CK( clk ) , .D( key_c_r_20_44 ) , .Q( key_c_r_21_44 ) );
  DFF_X1 key_c_r_reg_21_45 (.CK( clk ) , .D( key_c_r_20_45 ) , .Q( key_c_r_21_45 ) );
  DFF_X1 key_c_r_reg_21_46 (.CK( clk ) , .D( key_c_r_20_46 ) , .Q( key_c_r_21_46 ) );
  DFF_X1 key_c_r_reg_21_47 (.CK( clk ) , .D( key_c_r_20_47 ) , .Q( key_c_r_21_47 ) );
  DFF_X1 key_c_r_reg_21_48 (.CK( clk ) , .D( key_c_r_20_48 ) , .Q( key_c_r_21_48 ) );
  DFF_X1 key_c_r_reg_21_49 (.CK( clk ) , .D( key_c_r_20_49 ) , .Q( key_c_r_21_49 ) );
  DFF_X1 key_c_r_reg_21_5 (.CK( clk ) , .D( key_c_r_20_5 ) , .Q( key_c_r_21_5 ) );
  DFF_X1 key_c_r_reg_21_50 (.CK( clk ) , .D( key_c_r_20_50 ) , .Q( key_c_r_21_50 ) );
  DFF_X1 key_c_r_reg_21_51 (.CK( clk ) , .D( key_c_r_20_51 ) , .Q( key_c_r_21_51 ) );
  DFF_X1 key_c_r_reg_21_52 (.CK( clk ) , .D( key_c_r_20_52 ) , .Q( key_c_r_21_52 ) );
  DFF_X1 key_c_r_reg_21_53 (.CK( clk ) , .D( key_c_r_20_53 ) , .Q( key_c_r_21_53 ) );
  DFF_X1 key_c_r_reg_21_54 (.CK( clk ) , .D( key_c_r_20_54 ) , .Q( key_c_r_21_54 ) );
  DFF_X1 key_c_r_reg_21_55 (.CK( clk ) , .D( key_c_r_20_55 ) , .Q( key_c_r_21_55 ) );
  DFF_X1 key_c_r_reg_21_6 (.CK( clk ) , .D( key_c_r_20_6 ) , .Q( key_c_r_21_6 ) );
  DFF_X1 key_c_r_reg_21_7 (.CK( clk ) , .D( key_c_r_20_7 ) , .Q( key_c_r_21_7 ) );
  DFF_X1 key_c_r_reg_21_8 (.CK( clk ) , .D( key_c_r_20_8 ) , .Q( key_c_r_21_8 ) );
  DFF_X1 key_c_r_reg_21_9 (.CK( clk ) , .D( key_c_r_20_9 ) , .Q( key_c_r_21_9 ) );
  DFF_X1 key_c_r_reg_22_0 (.CK( clk ) , .D( key_c_r_21_0 ) , .Q( key_c_r_22_0 ) );
  DFF_X1 key_c_r_reg_22_1 (.CK( clk ) , .D( key_c_r_21_1 ) , .Q( key_c_r_22_1 ) );
  DFF_X1 key_c_r_reg_22_10 (.CK( clk ) , .D( key_c_r_21_10 ) , .Q( key_c_r_22_10 ) );
  DFF_X1 key_c_r_reg_22_11 (.CK( clk ) , .D( key_c_r_21_11 ) , .Q( key_c_r_22_11 ) );
  DFF_X1 key_c_r_reg_22_12 (.CK( clk ) , .D( key_c_r_21_12 ) , .Q( key_c_r_22_12 ) );
  DFF_X1 key_c_r_reg_22_13 (.CK( clk ) , .D( key_c_r_21_13 ) , .Q( key_c_r_22_13 ) );
  DFF_X1 key_c_r_reg_22_14 (.CK( clk ) , .D( key_c_r_21_14 ) , .Q( key_c_r_22_14 ) );
  DFF_X1 key_c_r_reg_22_15 (.CK( clk ) , .D( key_c_r_21_15 ) , .Q( key_c_r_22_15 ) );
  DFF_X1 key_c_r_reg_22_16 (.CK( clk ) , .D( key_c_r_21_16 ) , .Q( key_c_r_22_16 ) );
  DFF_X1 key_c_r_reg_22_17 (.CK( clk ) , .D( key_c_r_21_17 ) , .Q( key_c_r_22_17 ) );
  DFF_X1 key_c_r_reg_22_18 (.CK( clk ) , .D( key_c_r_21_18 ) , .Q( key_c_r_22_18 ) );
  DFF_X1 key_c_r_reg_22_19 (.CK( clk ) , .D( key_c_r_21_19 ) , .Q( key_c_r_22_19 ) );
  DFF_X1 key_c_r_reg_22_2 (.CK( clk ) , .D( key_c_r_21_2 ) , .Q( key_c_r_22_2 ) );
  DFF_X1 key_c_r_reg_22_20 (.CK( clk ) , .D( key_c_r_21_20 ) , .Q( key_c_r_22_20 ) );
  DFF_X1 key_c_r_reg_22_21 (.CK( clk ) , .D( key_c_r_21_21 ) , .Q( key_c_r_22_21 ) );
  DFF_X1 key_c_r_reg_22_22 (.CK( clk ) , .D( key_c_r_21_22 ) , .Q( key_c_r_22_22 ) );
  DFF_X1 key_c_r_reg_22_23 (.CK( clk ) , .D( key_c_r_21_23 ) , .Q( key_c_r_22_23 ) );
  DFF_X1 key_c_r_reg_22_24 (.CK( clk ) , .D( key_c_r_21_24 ) , .Q( key_c_r_22_24 ) );
  DFF_X1 key_c_r_reg_22_25 (.CK( clk ) , .D( key_c_r_21_25 ) , .Q( key_c_r_22_25 ) );
  DFF_X1 key_c_r_reg_22_26 (.CK( clk ) , .D( key_c_r_21_26 ) , .Q( key_c_r_22_26 ) );
  DFF_X1 key_c_r_reg_22_27 (.CK( clk ) , .D( key_c_r_21_27 ) , .Q( key_c_r_22_27 ) );
  DFF_X1 key_c_r_reg_22_28 (.CK( clk ) , .D( key_c_r_21_28 ) , .Q( key_c_r_22_28 ) );
  DFF_X1 key_c_r_reg_22_29 (.CK( clk ) , .D( key_c_r_21_29 ) , .Q( key_c_r_22_29 ) );
  DFF_X1 key_c_r_reg_22_3 (.CK( clk ) , .D( key_c_r_21_3 ) , .Q( key_c_r_22_3 ) );
  DFF_X1 key_c_r_reg_22_30 (.CK( clk ) , .D( key_c_r_21_30 ) , .Q( key_c_r_22_30 ) );
  DFF_X1 key_c_r_reg_22_31 (.CK( clk ) , .D( key_c_r_21_31 ) , .Q( key_c_r_22_31 ) );
  DFF_X1 key_c_r_reg_22_32 (.CK( clk ) , .D( key_c_r_21_32 ) , .Q( key_c_r_22_32 ) );
  DFF_X1 key_c_r_reg_22_33 (.CK( clk ) , .D( key_c_r_21_33 ) , .Q( key_c_r_22_33 ) );
  DFF_X1 key_c_r_reg_22_34 (.CK( clk ) , .D( key_c_r_21_34 ) , .Q( key_c_r_22_34 ) );
  DFF_X1 key_c_r_reg_22_35 (.CK( clk ) , .D( key_c_r_21_35 ) , .Q( key_c_r_22_35 ) );
  DFF_X1 key_c_r_reg_22_36 (.CK( clk ) , .D( key_c_r_21_36 ) , .Q( key_c_r_22_36 ) );
  DFF_X1 key_c_r_reg_22_37 (.CK( clk ) , .D( key_c_r_21_37 ) , .Q( key_c_r_22_37 ) );
  DFF_X1 key_c_r_reg_22_38 (.CK( clk ) , .D( key_c_r_21_38 ) , .Q( key_c_r_22_38 ) );
  DFF_X1 key_c_r_reg_22_39 (.CK( clk ) , .D( key_c_r_21_39 ) , .Q( key_c_r_22_39 ) );
  DFF_X1 key_c_r_reg_22_4 (.CK( clk ) , .D( key_c_r_21_4 ) , .Q( key_c_r_22_4 ) );
  DFF_X1 key_c_r_reg_22_40 (.CK( clk ) , .D( key_c_r_21_40 ) , .Q( key_c_r_22_40 ) );
  DFF_X1 key_c_r_reg_22_41 (.CK( clk ) , .D( key_c_r_21_41 ) , .Q( key_c_r_22_41 ) );
  DFF_X1 key_c_r_reg_22_42 (.CK( clk ) , .D( key_c_r_21_42 ) , .Q( key_c_r_22_42 ) );
  DFF_X1 key_c_r_reg_22_43 (.CK( clk ) , .D( key_c_r_21_43 ) , .Q( key_c_r_22_43 ) );
  DFF_X1 key_c_r_reg_22_44 (.CK( clk ) , .D( key_c_r_21_44 ) , .Q( key_c_r_22_44 ) );
  DFF_X1 key_c_r_reg_22_45 (.CK( clk ) , .D( key_c_r_21_45 ) , .Q( key_c_r_22_45 ) );
  DFF_X1 key_c_r_reg_22_46 (.CK( clk ) , .D( key_c_r_21_46 ) , .Q( key_c_r_22_46 ) );
  DFF_X1 key_c_r_reg_22_47 (.CK( clk ) , .D( key_c_r_21_47 ) , .Q( key_c_r_22_47 ) );
  DFF_X1 key_c_r_reg_22_48 (.CK( clk ) , .D( key_c_r_21_48 ) , .Q( key_c_r_22_48 ) );
  DFF_X1 key_c_r_reg_22_49 (.CK( clk ) , .D( key_c_r_21_49 ) , .Q( key_c_r_22_49 ) );
  DFF_X1 key_c_r_reg_22_5 (.CK( clk ) , .D( key_c_r_21_5 ) , .Q( key_c_r_22_5 ) );
  DFF_X1 key_c_r_reg_22_50 (.CK( clk ) , .D( key_c_r_21_50 ) , .Q( key_c_r_22_50 ) );
  DFF_X1 key_c_r_reg_22_51 (.CK( clk ) , .D( key_c_r_21_51 ) , .Q( key_c_r_22_51 ) );
  DFF_X1 key_c_r_reg_22_52 (.CK( clk ) , .D( key_c_r_21_52 ) , .Q( key_c_r_22_52 ) );
  DFF_X1 key_c_r_reg_22_53 (.CK( clk ) , .D( key_c_r_21_53 ) , .Q( key_c_r_22_53 ) );
  DFF_X1 key_c_r_reg_22_54 (.CK( clk ) , .D( key_c_r_21_54 ) , .Q( key_c_r_22_54 ) );
  DFF_X1 key_c_r_reg_22_55 (.CK( clk ) , .D( key_c_r_21_55 ) , .Q( key_c_r_22_55 ) );
  DFF_X1 key_c_r_reg_22_6 (.CK( clk ) , .D( key_c_r_21_6 ) , .Q( key_c_r_22_6 ) );
  DFF_X1 key_c_r_reg_22_7 (.CK( clk ) , .D( key_c_r_21_7 ) , .Q( key_c_r_22_7 ) );
  DFF_X1 key_c_r_reg_22_8 (.CK( clk ) , .D( key_c_r_21_8 ) , .Q( key_c_r_22_8 ) );
  DFF_X1 key_c_r_reg_22_9 (.CK( clk ) , .D( key_c_r_21_9 ) , .Q( key_c_r_22_9 ) );
  DFF_X1 key_c_r_reg_23_0 (.CK( clk ) , .D( key_c_r_22_0 ) , .Q( key_c_r_23_0 ) );
  DFF_X1 key_c_r_reg_23_1 (.CK( clk ) , .D( key_c_r_22_1 ) , .Q( key_c_r_23_1 ) );
  DFF_X1 key_c_r_reg_23_10 (.CK( clk ) , .D( key_c_r_22_10 ) , .Q( key_c_r_23_10 ) );
  DFF_X1 key_c_r_reg_23_11 (.CK( clk ) , .D( key_c_r_22_11 ) , .Q( key_c_r_23_11 ) );
  DFF_X1 key_c_r_reg_23_12 (.CK( clk ) , .D( key_c_r_22_12 ) , .Q( key_c_r_23_12 ) );
  DFF_X1 key_c_r_reg_23_13 (.CK( clk ) , .D( key_c_r_22_13 ) , .Q( key_c_r_23_13 ) );
  DFF_X1 key_c_r_reg_23_14 (.CK( clk ) , .D( key_c_r_22_14 ) , .Q( key_c_r_23_14 ) );
  DFF_X1 key_c_r_reg_23_15 (.CK( clk ) , .D( key_c_r_22_15 ) , .Q( key_c_r_23_15 ) );
  DFF_X1 key_c_r_reg_23_16 (.CK( clk ) , .D( key_c_r_22_16 ) , .Q( key_c_r_23_16 ) );
  DFF_X1 key_c_r_reg_23_17 (.CK( clk ) , .D( key_c_r_22_17 ) , .Q( key_c_r_23_17 ) );
  DFF_X1 key_c_r_reg_23_18 (.CK( clk ) , .D( key_c_r_22_18 ) , .Q( key_c_r_23_18 ) );
  DFF_X1 key_c_r_reg_23_19 (.CK( clk ) , .D( key_c_r_22_19 ) , .Q( key_c_r_23_19 ) );
  DFF_X1 key_c_r_reg_23_2 (.CK( clk ) , .D( key_c_r_22_2 ) , .Q( key_c_r_23_2 ) );
  DFF_X1 key_c_r_reg_23_20 (.CK( clk ) , .D( key_c_r_22_20 ) , .Q( key_c_r_23_20 ) );
  DFF_X1 key_c_r_reg_23_21 (.CK( clk ) , .D( key_c_r_22_21 ) , .Q( key_c_r_23_21 ) );
  DFF_X1 key_c_r_reg_23_22 (.CK( clk ) , .D( key_c_r_22_22 ) , .Q( key_c_r_23_22 ) );
  DFF_X1 key_c_r_reg_23_23 (.CK( clk ) , .D( key_c_r_22_23 ) , .Q( key_c_r_23_23 ) );
  DFF_X1 key_c_r_reg_23_24 (.CK( clk ) , .D( key_c_r_22_24 ) , .Q( key_c_r_23_24 ) );
  DFF_X1 key_c_r_reg_23_25 (.CK( clk ) , .D( key_c_r_22_25 ) , .Q( key_c_r_23_25 ) );
  DFF_X1 key_c_r_reg_23_26 (.CK( clk ) , .D( key_c_r_22_26 ) , .Q( key_c_r_23_26 ) );
  DFF_X1 key_c_r_reg_23_27 (.CK( clk ) , .D( key_c_r_22_27 ) , .Q( key_c_r_23_27 ) );
  DFF_X1 key_c_r_reg_23_28 (.CK( clk ) , .D( key_c_r_22_28 ) , .Q( key_c_r_23_28 ) );
  DFF_X1 key_c_r_reg_23_29 (.CK( clk ) , .D( key_c_r_22_29 ) , .Q( key_c_r_23_29 ) );
  DFF_X1 key_c_r_reg_23_3 (.CK( clk ) , .D( key_c_r_22_3 ) , .Q( key_c_r_23_3 ) );
  DFF_X1 key_c_r_reg_23_30 (.CK( clk ) , .D( key_c_r_22_30 ) , .Q( key_c_r_23_30 ) );
  DFF_X1 key_c_r_reg_23_31 (.CK( clk ) , .D( key_c_r_22_31 ) , .Q( key_c_r_23_31 ) );
  DFF_X1 key_c_r_reg_23_32 (.CK( clk ) , .D( key_c_r_22_32 ) , .Q( key_c_r_23_32 ) );
  DFF_X1 key_c_r_reg_23_33 (.CK( clk ) , .D( key_c_r_22_33 ) , .Q( key_c_r_23_33 ) );
  DFF_X1 key_c_r_reg_23_34 (.CK( clk ) , .D( key_c_r_22_34 ) , .Q( key_c_r_23_34 ) );
  DFF_X1 key_c_r_reg_23_35 (.CK( clk ) , .D( key_c_r_22_35 ) , .Q( key_c_r_23_35 ) );
  DFF_X1 key_c_r_reg_23_36 (.CK( clk ) , .D( key_c_r_22_36 ) , .Q( key_c_r_23_36 ) );
  DFF_X1 key_c_r_reg_23_37 (.CK( clk ) , .D( key_c_r_22_37 ) , .Q( key_c_r_23_37 ) );
  DFF_X1 key_c_r_reg_23_38 (.CK( clk ) , .D( key_c_r_22_38 ) , .Q( key_c_r_23_38 ) );
  DFF_X1 key_c_r_reg_23_39 (.CK( clk ) , .D( key_c_r_22_39 ) , .Q( key_c_r_23_39 ) );
  DFF_X1 key_c_r_reg_23_4 (.CK( clk ) , .D( key_c_r_22_4 ) , .Q( key_c_r_23_4 ) );
  DFF_X1 key_c_r_reg_23_40 (.CK( clk ) , .D( key_c_r_22_40 ) , .Q( key_c_r_23_40 ) );
  DFF_X1 key_c_r_reg_23_41 (.CK( clk ) , .D( key_c_r_22_41 ) , .Q( key_c_r_23_41 ) );
  DFF_X1 key_c_r_reg_23_42 (.CK( clk ) , .D( key_c_r_22_42 ) , .Q( key_c_r_23_42 ) );
  DFF_X1 key_c_r_reg_23_43 (.CK( clk ) , .D( key_c_r_22_43 ) , .Q( key_c_r_23_43 ) );
  DFF_X1 key_c_r_reg_23_44 (.CK( clk ) , .D( key_c_r_22_44 ) , .Q( key_c_r_23_44 ) );
  DFF_X1 key_c_r_reg_23_45 (.CK( clk ) , .D( key_c_r_22_45 ) , .Q( key_c_r_23_45 ) );
  DFF_X1 key_c_r_reg_23_46 (.CK( clk ) , .D( key_c_r_22_46 ) , .Q( key_c_r_23_46 ) );
  DFF_X1 key_c_r_reg_23_47 (.CK( clk ) , .D( key_c_r_22_47 ) , .Q( key_c_r_23_47 ) );
  DFF_X1 key_c_r_reg_23_48 (.CK( clk ) , .D( key_c_r_22_48 ) , .Q( key_c_r_23_48 ) );
  DFF_X1 key_c_r_reg_23_49 (.CK( clk ) , .D( key_c_r_22_49 ) , .Q( key_c_r_23_49 ) );
  DFF_X1 key_c_r_reg_23_5 (.CK( clk ) , .D( key_c_r_22_5 ) , .Q( key_c_r_23_5 ) );
  DFF_X1 key_c_r_reg_23_50 (.CK( clk ) , .D( key_c_r_22_50 ) , .Q( key_c_r_23_50 ) );
  DFF_X1 key_c_r_reg_23_51 (.CK( clk ) , .D( key_c_r_22_51 ) , .Q( key_c_r_23_51 ) );
  DFF_X1 key_c_r_reg_23_52 (.CK( clk ) , .D( key_c_r_22_52 ) , .Q( key_c_r_23_52 ) );
  DFF_X1 key_c_r_reg_23_53 (.CK( clk ) , .D( key_c_r_22_53 ) , .Q( key_c_r_23_53 ) );
  DFF_X1 key_c_r_reg_23_54 (.CK( clk ) , .D( key_c_r_22_54 ) , .Q( key_c_r_23_54 ) );
  DFF_X1 key_c_r_reg_23_55 (.CK( clk ) , .D( key_c_r_22_55 ) , .Q( key_c_r_23_55 ) );
  DFF_X1 key_c_r_reg_23_6 (.CK( clk ) , .D( key_c_r_22_6 ) , .Q( key_c_r_23_6 ) );
  DFF_X1 key_c_r_reg_23_7 (.CK( clk ) , .D( key_c_r_22_7 ) , .Q( key_c_r_23_7 ) );
  DFF_X1 key_c_r_reg_23_8 (.CK( clk ) , .D( key_c_r_22_8 ) , .Q( key_c_r_23_8 ) );
  DFF_X1 key_c_r_reg_23_9 (.CK( clk ) , .D( key_c_r_22_9 ) , .Q( key_c_r_23_9 ) );
  DFF_X1 key_c_r_reg_24_0 (.CK( clk ) , .D( key_c_r_23_0 ) , .Q( key_c_r_24_0 ) );
  DFF_X1 key_c_r_reg_24_1 (.CK( clk ) , .D( key_c_r_23_1 ) , .Q( key_c_r_24_1 ) );
  DFF_X1 key_c_r_reg_24_10 (.CK( clk ) , .D( key_c_r_23_10 ) , .Q( key_c_r_24_10 ) );
  DFF_X1 key_c_r_reg_24_11 (.CK( clk ) , .D( key_c_r_23_11 ) , .Q( key_c_r_24_11 ) );
  DFF_X1 key_c_r_reg_24_12 (.CK( clk ) , .D( key_c_r_23_12 ) , .Q( key_c_r_24_12 ) );
  DFF_X1 key_c_r_reg_24_13 (.CK( clk ) , .D( key_c_r_23_13 ) , .Q( key_c_r_24_13 ) );
  DFF_X1 key_c_r_reg_24_14 (.CK( clk ) , .D( key_c_r_23_14 ) , .Q( key_c_r_24_14 ) );
  DFF_X1 key_c_r_reg_24_15 (.CK( clk ) , .D( key_c_r_23_15 ) , .Q( key_c_r_24_15 ) );
  DFF_X1 key_c_r_reg_24_16 (.CK( clk ) , .D( key_c_r_23_16 ) , .Q( key_c_r_24_16 ) );
  DFF_X1 key_c_r_reg_24_17 (.CK( clk ) , .D( key_c_r_23_17 ) , .Q( key_c_r_24_17 ) );
  DFF_X1 key_c_r_reg_24_18 (.CK( clk ) , .D( key_c_r_23_18 ) , .Q( key_c_r_24_18 ) );
  DFF_X1 key_c_r_reg_24_19 (.CK( clk ) , .D( key_c_r_23_19 ) , .Q( key_c_r_24_19 ) );
  DFF_X1 key_c_r_reg_24_2 (.CK( clk ) , .D( key_c_r_23_2 ) , .Q( key_c_r_24_2 ) );
  DFF_X1 key_c_r_reg_24_20 (.CK( clk ) , .D( key_c_r_23_20 ) , .Q( key_c_r_24_20 ) );
  DFF_X1 key_c_r_reg_24_21 (.CK( clk ) , .D( key_c_r_23_21 ) , .Q( key_c_r_24_21 ) );
  DFF_X1 key_c_r_reg_24_22 (.CK( clk ) , .D( key_c_r_23_22 ) , .Q( key_c_r_24_22 ) );
  DFF_X1 key_c_r_reg_24_23 (.CK( clk ) , .D( key_c_r_23_23 ) , .Q( key_c_r_24_23 ) );
  DFF_X1 key_c_r_reg_24_24 (.CK( clk ) , .D( key_c_r_23_24 ) , .Q( key_c_r_24_24 ) );
  DFF_X1 key_c_r_reg_24_25 (.CK( clk ) , .D( key_c_r_23_25 ) , .Q( key_c_r_24_25 ) );
  DFF_X1 key_c_r_reg_24_26 (.CK( clk ) , .D( key_c_r_23_26 ) , .Q( key_c_r_24_26 ) );
  DFF_X1 key_c_r_reg_24_27 (.CK( clk ) , .D( key_c_r_23_27 ) , .Q( key_c_r_24_27 ) );
  DFF_X1 key_c_r_reg_24_28 (.CK( clk ) , .D( key_c_r_23_28 ) , .Q( key_c_r_24_28 ) );
  DFF_X1 key_c_r_reg_24_29 (.CK( clk ) , .D( key_c_r_23_29 ) , .Q( key_c_r_24_29 ) );
  DFF_X1 key_c_r_reg_24_3 (.CK( clk ) , .D( key_c_r_23_3 ) , .Q( key_c_r_24_3 ) );
  DFF_X1 key_c_r_reg_24_30 (.CK( clk ) , .D( key_c_r_23_30 ) , .Q( key_c_r_24_30 ) );
  DFF_X1 key_c_r_reg_24_31 (.CK( clk ) , .D( key_c_r_23_31 ) , .Q( key_c_r_24_31 ) );
  DFF_X1 key_c_r_reg_24_32 (.CK( clk ) , .D( key_c_r_23_32 ) , .Q( key_c_r_24_32 ) );
  DFF_X1 key_c_r_reg_24_33 (.CK( clk ) , .D( key_c_r_23_33 ) , .Q( key_c_r_24_33 ) );
  DFF_X1 key_c_r_reg_24_34 (.CK( clk ) , .D( key_c_r_23_34 ) , .Q( key_c_r_24_34 ) );
  DFF_X1 key_c_r_reg_24_35 (.CK( clk ) , .D( key_c_r_23_35 ) , .Q( key_c_r_24_35 ) );
  DFF_X1 key_c_r_reg_24_36 (.CK( clk ) , .D( key_c_r_23_36 ) , .Q( key_c_r_24_36 ) );
  DFF_X1 key_c_r_reg_24_37 (.CK( clk ) , .D( key_c_r_23_37 ) , .Q( key_c_r_24_37 ) );
  DFF_X1 key_c_r_reg_24_38 (.CK( clk ) , .D( key_c_r_23_38 ) , .Q( key_c_r_24_38 ) );
  DFF_X1 key_c_r_reg_24_39 (.CK( clk ) , .D( key_c_r_23_39 ) , .Q( key_c_r_24_39 ) );
  DFF_X1 key_c_r_reg_24_4 (.CK( clk ) , .D( key_c_r_23_4 ) , .Q( key_c_r_24_4 ) );
  DFF_X1 key_c_r_reg_24_40 (.CK( clk ) , .D( key_c_r_23_40 ) , .Q( key_c_r_24_40 ) );
  DFF_X1 key_c_r_reg_24_41 (.CK( clk ) , .D( key_c_r_23_41 ) , .Q( key_c_r_24_41 ) );
  DFF_X1 key_c_r_reg_24_42 (.CK( clk ) , .D( key_c_r_23_42 ) , .Q( key_c_r_24_42 ) );
  DFF_X1 key_c_r_reg_24_43 (.CK( clk ) , .D( key_c_r_23_43 ) , .Q( key_c_r_24_43 ) );
  DFF_X1 key_c_r_reg_24_44 (.CK( clk ) , .D( key_c_r_23_44 ) , .Q( key_c_r_24_44 ) );
  DFF_X1 key_c_r_reg_24_45 (.CK( clk ) , .D( key_c_r_23_45 ) , .Q( key_c_r_24_45 ) );
  DFF_X1 key_c_r_reg_24_46 (.CK( clk ) , .D( key_c_r_23_46 ) , .Q( key_c_r_24_46 ) );
  DFF_X1 key_c_r_reg_24_47 (.CK( clk ) , .D( key_c_r_23_47 ) , .Q( key_c_r_24_47 ) );
  DFF_X1 key_c_r_reg_24_48 (.CK( clk ) , .D( key_c_r_23_48 ) , .Q( key_c_r_24_48 ) );
  DFF_X1 key_c_r_reg_24_49 (.CK( clk ) , .D( key_c_r_23_49 ) , .Q( key_c_r_24_49 ) );
  DFF_X1 key_c_r_reg_24_5 (.CK( clk ) , .D( key_c_r_23_5 ) , .Q( key_c_r_24_5 ) );
  DFF_X1 key_c_r_reg_24_50 (.CK( clk ) , .D( key_c_r_23_50 ) , .Q( key_c_r_24_50 ) );
  DFF_X1 key_c_r_reg_24_51 (.CK( clk ) , .D( key_c_r_23_51 ) , .Q( key_c_r_24_51 ) );
  DFF_X1 key_c_r_reg_24_52 (.CK( clk ) , .D( key_c_r_23_52 ) , .Q( key_c_r_24_52 ) );
  DFF_X1 key_c_r_reg_24_53 (.CK( clk ) , .D( key_c_r_23_53 ) , .Q( key_c_r_24_53 ) );
  DFF_X1 key_c_r_reg_24_54 (.CK( clk ) , .D( key_c_r_23_54 ) , .Q( key_c_r_24_54 ) );
  DFF_X1 key_c_r_reg_24_55 (.CK( clk ) , .D( key_c_r_23_55 ) , .Q( key_c_r_24_55 ) );
  DFF_X1 key_c_r_reg_24_6 (.CK( clk ) , .D( key_c_r_23_6 ) , .Q( key_c_r_24_6 ) );
  DFF_X1 key_c_r_reg_24_7 (.CK( clk ) , .D( key_c_r_23_7 ) , .Q( key_c_r_24_7 ) );
  DFF_X1 key_c_r_reg_24_8 (.CK( clk ) , .D( key_c_r_23_8 ) , .Q( key_c_r_24_8 ) );
  DFF_X1 key_c_r_reg_24_9 (.CK( clk ) , .D( key_c_r_23_9 ) , .Q( key_c_r_24_9 ) );
  DFF_X1 key_c_r_reg_25_0 (.CK( clk ) , .D( key_c_r_24_0 ) , .Q( key_c_r_25_0 ) );
  DFF_X1 key_c_r_reg_25_1 (.CK( clk ) , .D( key_c_r_24_1 ) , .Q( key_c_r_25_1 ) );
  DFF_X1 key_c_r_reg_25_10 (.CK( clk ) , .D( key_c_r_24_10 ) , .Q( key_c_r_25_10 ) );
  DFF_X1 key_c_r_reg_25_11 (.CK( clk ) , .D( key_c_r_24_11 ) , .Q( key_c_r_25_11 ) );
  DFF_X1 key_c_r_reg_25_12 (.CK( clk ) , .D( key_c_r_24_12 ) , .Q( key_c_r_25_12 ) );
  DFF_X1 key_c_r_reg_25_13 (.CK( clk ) , .D( key_c_r_24_13 ) , .Q( key_c_r_25_13 ) );
  DFF_X1 key_c_r_reg_25_14 (.CK( clk ) , .D( key_c_r_24_14 ) , .Q( key_c_r_25_14 ) );
  DFF_X1 key_c_r_reg_25_15 (.CK( clk ) , .D( key_c_r_24_15 ) , .Q( key_c_r_25_15 ) );
  DFF_X1 key_c_r_reg_25_16 (.CK( clk ) , .D( key_c_r_24_16 ) , .Q( key_c_r_25_16 ) );
  DFF_X1 key_c_r_reg_25_17 (.CK( clk ) , .D( key_c_r_24_17 ) , .Q( key_c_r_25_17 ) );
  DFF_X1 key_c_r_reg_25_18 (.CK( clk ) , .D( key_c_r_24_18 ) , .Q( key_c_r_25_18 ) );
  DFF_X1 key_c_r_reg_25_19 (.CK( clk ) , .D( key_c_r_24_19 ) , .Q( key_c_r_25_19 ) );
  DFF_X1 key_c_r_reg_25_2 (.CK( clk ) , .D( key_c_r_24_2 ) , .Q( key_c_r_25_2 ) );
  DFF_X1 key_c_r_reg_25_20 (.CK( clk ) , .D( key_c_r_24_20 ) , .Q( key_c_r_25_20 ) );
  DFF_X1 key_c_r_reg_25_21 (.CK( clk ) , .D( key_c_r_24_21 ) , .Q( key_c_r_25_21 ) );
  DFF_X1 key_c_r_reg_25_22 (.CK( clk ) , .D( key_c_r_24_22 ) , .Q( key_c_r_25_22 ) );
  DFF_X1 key_c_r_reg_25_23 (.CK( clk ) , .D( key_c_r_24_23 ) , .Q( key_c_r_25_23 ) );
  DFF_X1 key_c_r_reg_25_24 (.CK( clk ) , .D( key_c_r_24_24 ) , .Q( key_c_r_25_24 ) );
  DFF_X1 key_c_r_reg_25_25 (.CK( clk ) , .D( key_c_r_24_25 ) , .Q( key_c_r_25_25 ) );
  DFF_X1 key_c_r_reg_25_26 (.CK( clk ) , .D( key_c_r_24_26 ) , .Q( key_c_r_25_26 ) );
  DFF_X1 key_c_r_reg_25_27 (.CK( clk ) , .D( key_c_r_24_27 ) , .Q( key_c_r_25_27 ) );
  DFF_X1 key_c_r_reg_25_28 (.CK( clk ) , .D( key_c_r_24_28 ) , .Q( key_c_r_25_28 ) );
  DFF_X1 key_c_r_reg_25_29 (.CK( clk ) , .D( key_c_r_24_29 ) , .Q( key_c_r_25_29 ) );
  DFF_X1 key_c_r_reg_25_3 (.CK( clk ) , .D( key_c_r_24_3 ) , .Q( key_c_r_25_3 ) );
  DFF_X1 key_c_r_reg_25_30 (.CK( clk ) , .D( key_c_r_24_30 ) , .Q( key_c_r_25_30 ) );
  DFF_X1 key_c_r_reg_25_31 (.CK( clk ) , .D( key_c_r_24_31 ) , .Q( key_c_r_25_31 ) );
  DFF_X1 key_c_r_reg_25_32 (.CK( clk ) , .D( key_c_r_24_32 ) , .Q( key_c_r_25_32 ) );
  DFF_X1 key_c_r_reg_25_33 (.CK( clk ) , .D( key_c_r_24_33 ) , .Q( key_c_r_25_33 ) );
  DFF_X1 key_c_r_reg_25_34 (.CK( clk ) , .D( key_c_r_24_34 ) , .Q( key_c_r_25_34 ) );
  DFF_X1 key_c_r_reg_25_35 (.CK( clk ) , .D( key_c_r_24_35 ) , .Q( key_c_r_25_35 ) );
  DFF_X1 key_c_r_reg_25_36 (.CK( clk ) , .D( key_c_r_24_36 ) , .Q( key_c_r_25_36 ) );
  DFF_X1 key_c_r_reg_25_37 (.CK( clk ) , .D( key_c_r_24_37 ) , .Q( key_c_r_25_37 ) );
  DFF_X1 key_c_r_reg_25_38 (.CK( clk ) , .D( key_c_r_24_38 ) , .Q( key_c_r_25_38 ) );
  DFF_X1 key_c_r_reg_25_39 (.CK( clk ) , .D( key_c_r_24_39 ) , .Q( key_c_r_25_39 ) );
  DFF_X1 key_c_r_reg_25_4 (.CK( clk ) , .D( key_c_r_24_4 ) , .Q( key_c_r_25_4 ) );
  DFF_X1 key_c_r_reg_25_40 (.CK( clk ) , .D( key_c_r_24_40 ) , .Q( key_c_r_25_40 ) );
  DFF_X1 key_c_r_reg_25_41 (.CK( clk ) , .D( key_c_r_24_41 ) , .Q( key_c_r_25_41 ) );
  DFF_X1 key_c_r_reg_25_42 (.CK( clk ) , .D( key_c_r_24_42 ) , .Q( key_c_r_25_42 ) );
  DFF_X1 key_c_r_reg_25_43 (.CK( clk ) , .D( key_c_r_24_43 ) , .Q( key_c_r_25_43 ) );
  DFF_X1 key_c_r_reg_25_44 (.CK( clk ) , .D( key_c_r_24_44 ) , .Q( key_c_r_25_44 ) );
  DFF_X1 key_c_r_reg_25_45 (.CK( clk ) , .D( key_c_r_24_45 ) , .Q( key_c_r_25_45 ) );
  DFF_X1 key_c_r_reg_25_46 (.CK( clk ) , .D( key_c_r_24_46 ) , .Q( key_c_r_25_46 ) );
  DFF_X1 key_c_r_reg_25_47 (.CK( clk ) , .D( key_c_r_24_47 ) , .Q( key_c_r_25_47 ) );
  DFF_X1 key_c_r_reg_25_48 (.CK( clk ) , .D( key_c_r_24_48 ) , .Q( key_c_r_25_48 ) );
  DFF_X1 key_c_r_reg_25_49 (.CK( clk ) , .D( key_c_r_24_49 ) , .Q( key_c_r_25_49 ) );
  DFF_X1 key_c_r_reg_25_5 (.CK( clk ) , .D( key_c_r_24_5 ) , .Q( key_c_r_25_5 ) );
  DFF_X1 key_c_r_reg_25_50 (.CK( clk ) , .D( key_c_r_24_50 ) , .Q( key_c_r_25_50 ) );
  DFF_X1 key_c_r_reg_25_51 (.CK( clk ) , .D( key_c_r_24_51 ) , .Q( key_c_r_25_51 ) );
  DFF_X1 key_c_r_reg_25_52 (.CK( clk ) , .D( key_c_r_24_52 ) , .Q( key_c_r_25_52 ) );
  DFF_X1 key_c_r_reg_25_53 (.CK( clk ) , .D( key_c_r_24_53 ) , .Q( key_c_r_25_53 ) );
  DFF_X1 key_c_r_reg_25_54 (.CK( clk ) , .D( key_c_r_24_54 ) , .Q( key_c_r_25_54 ) );
  DFF_X1 key_c_r_reg_25_55 (.CK( clk ) , .D( key_c_r_24_55 ) , .Q( key_c_r_25_55 ) );
  DFF_X1 key_c_r_reg_25_6 (.CK( clk ) , .D( key_c_r_24_6 ) , .Q( key_c_r_25_6 ) );
  DFF_X1 key_c_r_reg_25_7 (.CK( clk ) , .D( key_c_r_24_7 ) , .Q( key_c_r_25_7 ) );
  DFF_X1 key_c_r_reg_25_8 (.CK( clk ) , .D( key_c_r_24_8 ) , .Q( key_c_r_25_8 ) );
  DFF_X1 key_c_r_reg_25_9 (.CK( clk ) , .D( key_c_r_24_9 ) , .Q( key_c_r_25_9 ) );
  DFF_X1 key_c_r_reg_26_0 (.CK( clk ) , .D( key_c_r_25_0 ) , .Q( key_c_r_26_0 ) );
  DFF_X1 key_c_r_reg_26_1 (.CK( clk ) , .D( key_c_r_25_1 ) , .Q( key_c_r_26_1 ) );
  DFF_X1 key_c_r_reg_26_10 (.CK( clk ) , .D( key_c_r_25_10 ) , .Q( key_c_r_26_10 ) );
  DFF_X1 key_c_r_reg_26_11 (.CK( clk ) , .D( key_c_r_25_11 ) , .Q( key_c_r_26_11 ) );
  DFF_X1 key_c_r_reg_26_12 (.CK( clk ) , .D( key_c_r_25_12 ) , .Q( key_c_r_26_12 ) );
  DFF_X1 key_c_r_reg_26_13 (.CK( clk ) , .D( key_c_r_25_13 ) , .Q( key_c_r_26_13 ) );
  DFF_X1 key_c_r_reg_26_14 (.CK( clk ) , .D( key_c_r_25_14 ) , .Q( key_c_r_26_14 ) );
  DFF_X1 key_c_r_reg_26_15 (.CK( clk ) , .D( key_c_r_25_15 ) , .Q( key_c_r_26_15 ) );
  DFF_X1 key_c_r_reg_26_16 (.CK( clk ) , .D( key_c_r_25_16 ) , .Q( key_c_r_26_16 ) );
  DFF_X1 key_c_r_reg_26_17 (.CK( clk ) , .D( key_c_r_25_17 ) , .Q( key_c_r_26_17 ) );
  DFF_X1 key_c_r_reg_26_18 (.CK( clk ) , .D( key_c_r_25_18 ) , .Q( key_c_r_26_18 ) );
  DFF_X1 key_c_r_reg_26_19 (.CK( clk ) , .D( key_c_r_25_19 ) , .Q( key_c_r_26_19 ) );
  DFF_X1 key_c_r_reg_26_2 (.CK( clk ) , .D( key_c_r_25_2 ) , .Q( key_c_r_26_2 ) );
  DFF_X1 key_c_r_reg_26_20 (.CK( clk ) , .D( key_c_r_25_20 ) , .Q( key_c_r_26_20 ) );
  DFF_X1 key_c_r_reg_26_21 (.CK( clk ) , .D( key_c_r_25_21 ) , .Q( key_c_r_26_21 ) );
  DFF_X1 key_c_r_reg_26_22 (.CK( clk ) , .D( key_c_r_25_22 ) , .Q( key_c_r_26_22 ) );
  DFF_X1 key_c_r_reg_26_23 (.CK( clk ) , .D( key_c_r_25_23 ) , .Q( key_c_r_26_23 ) );
  DFF_X1 key_c_r_reg_26_24 (.CK( clk ) , .D( key_c_r_25_24 ) , .Q( key_c_r_26_24 ) );
  DFF_X1 key_c_r_reg_26_25 (.CK( clk ) , .D( key_c_r_25_25 ) , .Q( key_c_r_26_25 ) );
  DFF_X1 key_c_r_reg_26_26 (.CK( clk ) , .D( key_c_r_25_26 ) , .Q( key_c_r_26_26 ) );
  DFF_X1 key_c_r_reg_26_27 (.CK( clk ) , .D( key_c_r_25_27 ) , .Q( key_c_r_26_27 ) );
  DFF_X1 key_c_r_reg_26_28 (.CK( clk ) , .D( key_c_r_25_28 ) , .Q( key_c_r_26_28 ) );
  DFF_X1 key_c_r_reg_26_29 (.CK( clk ) , .D( key_c_r_25_29 ) , .Q( key_c_r_26_29 ) );
  DFF_X1 key_c_r_reg_26_3 (.CK( clk ) , .D( key_c_r_25_3 ) , .Q( key_c_r_26_3 ) );
  DFF_X1 key_c_r_reg_26_30 (.CK( clk ) , .D( key_c_r_25_30 ) , .Q( key_c_r_26_30 ) );
  DFF_X1 key_c_r_reg_26_31 (.CK( clk ) , .D( key_c_r_25_31 ) , .Q( key_c_r_26_31 ) );
  DFF_X1 key_c_r_reg_26_32 (.CK( clk ) , .D( key_c_r_25_32 ) , .Q( key_c_r_26_32 ) );
  DFF_X1 key_c_r_reg_26_33 (.CK( clk ) , .D( key_c_r_25_33 ) , .Q( key_c_r_26_33 ) );
  DFF_X1 key_c_r_reg_26_34 (.CK( clk ) , .D( key_c_r_25_34 ) , .Q( key_c_r_26_34 ) );
  DFF_X1 key_c_r_reg_26_35 (.CK( clk ) , .D( key_c_r_25_35 ) , .Q( key_c_r_26_35 ) );
  DFF_X1 key_c_r_reg_26_36 (.CK( clk ) , .D( key_c_r_25_36 ) , .Q( key_c_r_26_36 ) );
  DFF_X1 key_c_r_reg_26_37 (.CK( clk ) , .D( key_c_r_25_37 ) , .Q( key_c_r_26_37 ) );
  DFF_X1 key_c_r_reg_26_38 (.CK( clk ) , .D( key_c_r_25_38 ) , .Q( key_c_r_26_38 ) );
  DFF_X1 key_c_r_reg_26_39 (.CK( clk ) , .D( key_c_r_25_39 ) , .Q( key_c_r_26_39 ) );
  DFF_X1 key_c_r_reg_26_4 (.CK( clk ) , .D( key_c_r_25_4 ) , .Q( key_c_r_26_4 ) );
  DFF_X1 key_c_r_reg_26_40 (.CK( clk ) , .D( key_c_r_25_40 ) , .Q( key_c_r_26_40 ) );
  DFF_X1 key_c_r_reg_26_41 (.CK( clk ) , .D( key_c_r_25_41 ) , .Q( key_c_r_26_41 ) );
  DFF_X1 key_c_r_reg_26_42 (.CK( clk ) , .D( key_c_r_25_42 ) , .Q( key_c_r_26_42 ) );
  DFF_X1 key_c_r_reg_26_43 (.CK( clk ) , .D( key_c_r_25_43 ) , .Q( key_c_r_26_43 ) );
  DFF_X1 key_c_r_reg_26_44 (.CK( clk ) , .D( key_c_r_25_44 ) , .Q( key_c_r_26_44 ) );
  DFF_X1 key_c_r_reg_26_45 (.CK( clk ) , .D( key_c_r_25_45 ) , .Q( key_c_r_26_45 ) );
  DFF_X1 key_c_r_reg_26_46 (.CK( clk ) , .D( key_c_r_25_46 ) , .Q( key_c_r_26_46 ) );
  DFF_X1 key_c_r_reg_26_47 (.CK( clk ) , .D( key_c_r_25_47 ) , .Q( key_c_r_26_47 ) );
  DFF_X1 key_c_r_reg_26_48 (.CK( clk ) , .D( key_c_r_25_48 ) , .Q( key_c_r_26_48 ) );
  DFF_X1 key_c_r_reg_26_49 (.CK( clk ) , .D( key_c_r_25_49 ) , .Q( key_c_r_26_49 ) );
  DFF_X1 key_c_r_reg_26_5 (.CK( clk ) , .D( key_c_r_25_5 ) , .Q( key_c_r_26_5 ) );
  DFF_X1 key_c_r_reg_26_50 (.CK( clk ) , .D( key_c_r_25_50 ) , .Q( key_c_r_26_50 ) );
  DFF_X1 key_c_r_reg_26_51 (.CK( clk ) , .D( key_c_r_25_51 ) , .Q( key_c_r_26_51 ) );
  DFF_X1 key_c_r_reg_26_52 (.CK( clk ) , .D( key_c_r_25_52 ) , .Q( key_c_r_26_52 ) );
  DFF_X1 key_c_r_reg_26_53 (.CK( clk ) , .D( key_c_r_25_53 ) , .Q( key_c_r_26_53 ) );
  DFF_X1 key_c_r_reg_26_54 (.CK( clk ) , .D( key_c_r_25_54 ) , .Q( key_c_r_26_54 ) );
  DFF_X1 key_c_r_reg_26_55 (.CK( clk ) , .D( key_c_r_25_55 ) , .Q( key_c_r_26_55 ) );
  DFF_X1 key_c_r_reg_26_6 (.CK( clk ) , .D( key_c_r_25_6 ) , .Q( key_c_r_26_6 ) );
  DFF_X1 key_c_r_reg_26_7 (.CK( clk ) , .D( key_c_r_25_7 ) , .Q( key_c_r_26_7 ) );
  DFF_X1 key_c_r_reg_26_8 (.CK( clk ) , .D( key_c_r_25_8 ) , .Q( key_c_r_26_8 ) );
  DFF_X1 key_c_r_reg_26_9 (.CK( clk ) , .D( key_c_r_25_9 ) , .Q( key_c_r_26_9 ) );
  DFF_X1 key_c_r_reg_27_0 (.CK( clk ) , .D( key_c_r_26_0 ) , .Q( key_c_r_27_0 ) );
  DFF_X1 key_c_r_reg_27_1 (.CK( clk ) , .D( key_c_r_26_1 ) , .Q( key_c_r_27_1 ) );
  DFF_X1 key_c_r_reg_27_10 (.CK( clk ) , .D( key_c_r_26_10 ) , .Q( key_c_r_27_10 ) );
  DFF_X1 key_c_r_reg_27_11 (.CK( clk ) , .D( key_c_r_26_11 ) , .Q( key_c_r_27_11 ) );
  DFF_X1 key_c_r_reg_27_12 (.CK( clk ) , .D( key_c_r_26_12 ) , .Q( key_c_r_27_12 ) );
  DFF_X1 key_c_r_reg_27_13 (.CK( clk ) , .D( key_c_r_26_13 ) , .Q( key_c_r_27_13 ) );
  DFF_X1 key_c_r_reg_27_14 (.CK( clk ) , .D( key_c_r_26_14 ) , .Q( key_c_r_27_14 ) );
  DFF_X1 key_c_r_reg_27_15 (.CK( clk ) , .D( key_c_r_26_15 ) , .Q( key_c_r_27_15 ) );
  DFF_X1 key_c_r_reg_27_16 (.CK( clk ) , .D( key_c_r_26_16 ) , .Q( key_c_r_27_16 ) );
  DFF_X1 key_c_r_reg_27_17 (.CK( clk ) , .D( key_c_r_26_17 ) , .Q( key_c_r_27_17 ) );
  DFF_X1 key_c_r_reg_27_18 (.CK( clk ) , .D( key_c_r_26_18 ) , .Q( key_c_r_27_18 ) );
  DFF_X1 key_c_r_reg_27_19 (.CK( clk ) , .D( key_c_r_26_19 ) , .Q( key_c_r_27_19 ) );
  DFF_X1 key_c_r_reg_27_2 (.CK( clk ) , .D( key_c_r_26_2 ) , .Q( key_c_r_27_2 ) );
  DFF_X1 key_c_r_reg_27_20 (.CK( clk ) , .D( key_c_r_26_20 ) , .Q( key_c_r_27_20 ) );
  DFF_X1 key_c_r_reg_27_21 (.CK( clk ) , .D( key_c_r_26_21 ) , .Q( key_c_r_27_21 ) );
  DFF_X1 key_c_r_reg_27_22 (.CK( clk ) , .D( key_c_r_26_22 ) , .Q( key_c_r_27_22 ) );
  DFF_X1 key_c_r_reg_27_23 (.CK( clk ) , .D( key_c_r_26_23 ) , .Q( key_c_r_27_23 ) );
  DFF_X1 key_c_r_reg_27_24 (.CK( clk ) , .D( key_c_r_26_24 ) , .Q( key_c_r_27_24 ) );
  DFF_X1 key_c_r_reg_27_25 (.CK( clk ) , .D( key_c_r_26_25 ) , .Q( key_c_r_27_25 ) );
  DFF_X1 key_c_r_reg_27_26 (.CK( clk ) , .D( key_c_r_26_26 ) , .Q( key_c_r_27_26 ) );
  DFF_X1 key_c_r_reg_27_27 (.CK( clk ) , .D( key_c_r_26_27 ) , .Q( key_c_r_27_27 ) );
  DFF_X1 key_c_r_reg_27_28 (.CK( clk ) , .D( key_c_r_26_28 ) , .Q( key_c_r_27_28 ) );
  DFF_X1 key_c_r_reg_27_29 (.CK( clk ) , .D( key_c_r_26_29 ) , .Q( key_c_r_27_29 ) );
  DFF_X1 key_c_r_reg_27_3 (.CK( clk ) , .D( key_c_r_26_3 ) , .Q( key_c_r_27_3 ) );
  DFF_X1 key_c_r_reg_27_30 (.CK( clk ) , .D( key_c_r_26_30 ) , .Q( key_c_r_27_30 ) );
  DFF_X1 key_c_r_reg_27_31 (.CK( clk ) , .D( key_c_r_26_31 ) , .Q( key_c_r_27_31 ) );
  DFF_X1 key_c_r_reg_27_32 (.CK( clk ) , .D( key_c_r_26_32 ) , .Q( key_c_r_27_32 ) );
  DFF_X1 key_c_r_reg_27_33 (.CK( clk ) , .D( key_c_r_26_33 ) , .Q( key_c_r_27_33 ) );
  DFF_X1 key_c_r_reg_27_34 (.CK( clk ) , .D( key_c_r_26_34 ) , .Q( key_c_r_27_34 ) );
  DFF_X1 key_c_r_reg_27_35 (.CK( clk ) , .D( key_c_r_26_35 ) , .Q( key_c_r_27_35 ) );
  DFF_X1 key_c_r_reg_27_36 (.CK( clk ) , .D( key_c_r_26_36 ) , .Q( key_c_r_27_36 ) );
  DFF_X1 key_c_r_reg_27_37 (.CK( clk ) , .D( key_c_r_26_37 ) , .Q( key_c_r_27_37 ) );
  DFF_X1 key_c_r_reg_27_38 (.CK( clk ) , .D( key_c_r_26_38 ) , .Q( key_c_r_27_38 ) );
  DFF_X1 key_c_r_reg_27_39 (.CK( clk ) , .D( key_c_r_26_39 ) , .Q( key_c_r_27_39 ) );
  DFF_X1 key_c_r_reg_27_4 (.CK( clk ) , .D( key_c_r_26_4 ) , .Q( key_c_r_27_4 ) );
  DFF_X1 key_c_r_reg_27_40 (.CK( clk ) , .D( key_c_r_26_40 ) , .Q( key_c_r_27_40 ) );
  DFF_X1 key_c_r_reg_27_41 (.CK( clk ) , .D( key_c_r_26_41 ) , .Q( key_c_r_27_41 ) );
  DFF_X1 key_c_r_reg_27_42 (.CK( clk ) , .D( key_c_r_26_42 ) , .Q( key_c_r_27_42 ) );
  DFF_X1 key_c_r_reg_27_43 (.CK( clk ) , .D( key_c_r_26_43 ) , .Q( key_c_r_27_43 ) );
  DFF_X1 key_c_r_reg_27_44 (.CK( clk ) , .D( key_c_r_26_44 ) , .Q( key_c_r_27_44 ) );
  DFF_X1 key_c_r_reg_27_45 (.CK( clk ) , .D( key_c_r_26_45 ) , .Q( key_c_r_27_45 ) );
  DFF_X1 key_c_r_reg_27_46 (.CK( clk ) , .D( key_c_r_26_46 ) , .Q( key_c_r_27_46 ) );
  DFF_X1 key_c_r_reg_27_47 (.CK( clk ) , .D( key_c_r_26_47 ) , .Q( key_c_r_27_47 ) );
  DFF_X1 key_c_r_reg_27_48 (.CK( clk ) , .D( key_c_r_26_48 ) , .Q( key_c_r_27_48 ) );
  DFF_X1 key_c_r_reg_27_49 (.CK( clk ) , .D( key_c_r_26_49 ) , .Q( key_c_r_27_49 ) );
  DFF_X1 key_c_r_reg_27_5 (.CK( clk ) , .D( key_c_r_26_5 ) , .Q( key_c_r_27_5 ) );
  DFF_X1 key_c_r_reg_27_50 (.CK( clk ) , .D( key_c_r_26_50 ) , .Q( key_c_r_27_50 ) );
  DFF_X1 key_c_r_reg_27_51 (.CK( clk ) , .D( key_c_r_26_51 ) , .Q( key_c_r_27_51 ) );
  DFF_X1 key_c_r_reg_27_52 (.CK( clk ) , .D( key_c_r_26_52 ) , .Q( key_c_r_27_52 ) );
  DFF_X1 key_c_r_reg_27_53 (.CK( clk ) , .D( key_c_r_26_53 ) , .Q( key_c_r_27_53 ) );
  DFF_X1 key_c_r_reg_27_54 (.CK( clk ) , .D( key_c_r_26_54 ) , .Q( key_c_r_27_54 ) );
  DFF_X1 key_c_r_reg_27_55 (.CK( clk ) , .D( key_c_r_26_55 ) , .Q( key_c_r_27_55 ) );
  DFF_X1 key_c_r_reg_27_6 (.CK( clk ) , .D( key_c_r_26_6 ) , .Q( key_c_r_27_6 ) );
  DFF_X1 key_c_r_reg_27_7 (.CK( clk ) , .D( key_c_r_26_7 ) , .Q( key_c_r_27_7 ) );
  DFF_X1 key_c_r_reg_27_8 (.CK( clk ) , .D( key_c_r_26_8 ) , .Q( key_c_r_27_8 ) );
  DFF_X1 key_c_r_reg_27_9 (.CK( clk ) , .D( key_c_r_26_9 ) , .Q( key_c_r_27_9 ) );
  DFF_X1 key_c_r_reg_28_0 (.CK( clk ) , .D( key_c_r_27_0 ) , .Q( key_c_r_28_0 ) );
  DFF_X1 key_c_r_reg_28_1 (.CK( clk ) , .D( key_c_r_27_1 ) , .Q( key_c_r_28_1 ) );
  DFF_X1 key_c_r_reg_28_10 (.CK( clk ) , .D( key_c_r_27_10 ) , .Q( key_c_r_28_10 ) );
  DFF_X1 key_c_r_reg_28_11 (.CK( clk ) , .D( key_c_r_27_11 ) , .Q( key_c_r_28_11 ) );
  DFF_X1 key_c_r_reg_28_12 (.CK( clk ) , .D( key_c_r_27_12 ) , .Q( key_c_r_28_12 ) );
  DFF_X1 key_c_r_reg_28_13 (.CK( clk ) , .D( key_c_r_27_13 ) , .Q( key_c_r_28_13 ) );
  DFF_X1 key_c_r_reg_28_14 (.CK( clk ) , .D( key_c_r_27_14 ) , .Q( key_c_r_28_14 ) );
  DFF_X1 key_c_r_reg_28_15 (.CK( clk ) , .D( key_c_r_27_15 ) , .Q( key_c_r_28_15 ) );
  DFF_X1 key_c_r_reg_28_16 (.CK( clk ) , .D( key_c_r_27_16 ) , .Q( key_c_r_28_16 ) );
  DFF_X1 key_c_r_reg_28_17 (.CK( clk ) , .D( key_c_r_27_17 ) , .Q( key_c_r_28_17 ) );
  DFF_X1 key_c_r_reg_28_18 (.CK( clk ) , .D( key_c_r_27_18 ) , .Q( key_c_r_28_18 ) );
  DFF_X1 key_c_r_reg_28_19 (.CK( clk ) , .D( key_c_r_27_19 ) , .Q( key_c_r_28_19 ) );
  DFF_X1 key_c_r_reg_28_2 (.CK( clk ) , .D( key_c_r_27_2 ) , .Q( key_c_r_28_2 ) );
  DFF_X1 key_c_r_reg_28_20 (.CK( clk ) , .D( key_c_r_27_20 ) , .Q( key_c_r_28_20 ) );
  DFF_X1 key_c_r_reg_28_21 (.CK( clk ) , .D( key_c_r_27_21 ) , .Q( key_c_r_28_21 ) );
  DFF_X1 key_c_r_reg_28_22 (.CK( clk ) , .D( key_c_r_27_22 ) , .Q( key_c_r_28_22 ) );
  DFF_X1 key_c_r_reg_28_23 (.CK( clk ) , .D( key_c_r_27_23 ) , .Q( key_c_r_28_23 ) );
  DFF_X1 key_c_r_reg_28_24 (.CK( clk ) , .D( key_c_r_27_24 ) , .Q( key_c_r_28_24 ) );
  DFF_X1 key_c_r_reg_28_25 (.CK( clk ) , .D( key_c_r_27_25 ) , .Q( key_c_r_28_25 ) );
  DFF_X1 key_c_r_reg_28_26 (.CK( clk ) , .D( key_c_r_27_26 ) , .Q( key_c_r_28_26 ) );
  DFF_X1 key_c_r_reg_28_27 (.CK( clk ) , .D( key_c_r_27_27 ) , .Q( key_c_r_28_27 ) );
  DFF_X1 key_c_r_reg_28_28 (.CK( clk ) , .D( key_c_r_27_28 ) , .Q( key_c_r_28_28 ) );
  DFF_X1 key_c_r_reg_28_29 (.CK( clk ) , .D( key_c_r_27_29 ) , .Q( key_c_r_28_29 ) );
  DFF_X1 key_c_r_reg_28_3 (.CK( clk ) , .D( key_c_r_27_3 ) , .Q( key_c_r_28_3 ) );
  DFF_X1 key_c_r_reg_28_30 (.CK( clk ) , .D( key_c_r_27_30 ) , .Q( key_c_r_28_30 ) );
  DFF_X1 key_c_r_reg_28_31 (.CK( clk ) , .D( key_c_r_27_31 ) , .Q( key_c_r_28_31 ) );
  DFF_X1 key_c_r_reg_28_32 (.CK( clk ) , .D( key_c_r_27_32 ) , .Q( key_c_r_28_32 ) );
  DFF_X1 key_c_r_reg_28_33 (.CK( clk ) , .D( key_c_r_27_33 ) , .Q( key_c_r_28_33 ) );
  DFF_X1 key_c_r_reg_28_34 (.CK( clk ) , .D( key_c_r_27_34 ) , .Q( key_c_r_28_34 ) );
  DFF_X1 key_c_r_reg_28_35 (.CK( clk ) , .D( key_c_r_27_35 ) , .Q( key_c_r_28_35 ) );
  DFF_X1 key_c_r_reg_28_36 (.CK( clk ) , .D( key_c_r_27_36 ) , .Q( key_c_r_28_36 ) );
  DFF_X1 key_c_r_reg_28_37 (.CK( clk ) , .D( key_c_r_27_37 ) , .Q( key_c_r_28_37 ) );
  DFF_X1 key_c_r_reg_28_38 (.CK( clk ) , .D( key_c_r_27_38 ) , .Q( key_c_r_28_38 ) );
  DFF_X1 key_c_r_reg_28_39 (.CK( clk ) , .D( key_c_r_27_39 ) , .Q( key_c_r_28_39 ) );
  DFF_X1 key_c_r_reg_28_4 (.CK( clk ) , .D( key_c_r_27_4 ) , .Q( key_c_r_28_4 ) );
  DFF_X1 key_c_r_reg_28_40 (.CK( clk ) , .D( key_c_r_27_40 ) , .Q( key_c_r_28_40 ) );
  DFF_X1 key_c_r_reg_28_41 (.CK( clk ) , .D( key_c_r_27_41 ) , .Q( key_c_r_28_41 ) );
  DFF_X1 key_c_r_reg_28_42 (.CK( clk ) , .D( key_c_r_27_42 ) , .Q( key_c_r_28_42 ) );
  DFF_X1 key_c_r_reg_28_43 (.CK( clk ) , .D( key_c_r_27_43 ) , .Q( key_c_r_28_43 ) );
  DFF_X1 key_c_r_reg_28_44 (.CK( clk ) , .D( key_c_r_27_44 ) , .Q( key_c_r_28_44 ) );
  DFF_X1 key_c_r_reg_28_45 (.CK( clk ) , .D( key_c_r_27_45 ) , .Q( key_c_r_28_45 ) );
  DFF_X1 key_c_r_reg_28_46 (.CK( clk ) , .D( key_c_r_27_46 ) , .Q( key_c_r_28_46 ) );
  DFF_X1 key_c_r_reg_28_47 (.CK( clk ) , .D( key_c_r_27_47 ) , .Q( key_c_r_28_47 ) );
  DFF_X1 key_c_r_reg_28_48 (.CK( clk ) , .D( key_c_r_27_48 ) , .Q( key_c_r_28_48 ) );
  DFF_X1 key_c_r_reg_28_49 (.CK( clk ) , .D( key_c_r_27_49 ) , .Q( key_c_r_28_49 ) );
  DFF_X1 key_c_r_reg_28_5 (.CK( clk ) , .D( key_c_r_27_5 ) , .Q( key_c_r_28_5 ) );
  DFF_X1 key_c_r_reg_28_50 (.CK( clk ) , .D( key_c_r_27_50 ) , .Q( key_c_r_28_50 ) );
  DFF_X1 key_c_r_reg_28_51 (.CK( clk ) , .D( key_c_r_27_51 ) , .Q( key_c_r_28_51 ) );
  DFF_X1 key_c_r_reg_28_52 (.CK( clk ) , .D( key_c_r_27_52 ) , .Q( key_c_r_28_52 ) );
  DFF_X1 key_c_r_reg_28_53 (.CK( clk ) , .D( key_c_r_27_53 ) , .Q( key_c_r_28_53 ) );
  DFF_X1 key_c_r_reg_28_54 (.CK( clk ) , .D( key_c_r_27_54 ) , .Q( key_c_r_28_54 ) );
  DFF_X1 key_c_r_reg_28_55 (.CK( clk ) , .D( key_c_r_27_55 ) , .Q( key_c_r_28_55 ) );
  DFF_X1 key_c_r_reg_28_6 (.CK( clk ) , .D( key_c_r_27_6 ) , .Q( key_c_r_28_6 ) );
  DFF_X1 key_c_r_reg_28_7 (.CK( clk ) , .D( key_c_r_27_7 ) , .Q( key_c_r_28_7 ) );
  DFF_X1 key_c_r_reg_28_8 (.CK( clk ) , .D( key_c_r_27_8 ) , .Q( key_c_r_28_8 ) );
  DFF_X1 key_c_r_reg_28_9 (.CK( clk ) , .D( key_c_r_27_9 ) , .Q( key_c_r_28_9 ) );
  DFF_X1 key_c_r_reg_29_0 (.CK( clk ) , .D( key_c_r_28_0 ) , .Q( key_c_r_29_0 ) );
  DFF_X1 key_c_r_reg_29_1 (.CK( clk ) , .D( key_c_r_28_1 ) , .Q( key_c_r_29_1 ) );
  DFF_X1 key_c_r_reg_29_10 (.CK( clk ) , .D( key_c_r_28_10 ) , .Q( key_c_r_29_10 ) );
  DFF_X1 key_c_r_reg_29_11 (.CK( clk ) , .D( key_c_r_28_11 ) , .Q( key_c_r_29_11 ) );
  DFF_X1 key_c_r_reg_29_12 (.CK( clk ) , .D( key_c_r_28_12 ) , .Q( key_c_r_29_12 ) );
  DFF_X1 key_c_r_reg_29_13 (.CK( clk ) , .D( key_c_r_28_13 ) , .Q( key_c_r_29_13 ) );
  DFF_X1 key_c_r_reg_29_14 (.CK( clk ) , .D( key_c_r_28_14 ) , .Q( key_c_r_29_14 ) );
  DFF_X1 key_c_r_reg_29_15 (.CK( clk ) , .D( key_c_r_28_15 ) , .Q( key_c_r_29_15 ) );
  DFF_X1 key_c_r_reg_29_16 (.CK( clk ) , .D( key_c_r_28_16 ) , .Q( key_c_r_29_16 ) );
  DFF_X1 key_c_r_reg_29_17 (.CK( clk ) , .D( key_c_r_28_17 ) , .Q( key_c_r_29_17 ) );
  DFF_X1 key_c_r_reg_29_18 (.CK( clk ) , .D( key_c_r_28_18 ) , .Q( key_c_r_29_18 ) );
  DFF_X1 key_c_r_reg_29_19 (.CK( clk ) , .D( key_c_r_28_19 ) , .Q( key_c_r_29_19 ) );
  DFF_X1 key_c_r_reg_29_2 (.CK( clk ) , .D( key_c_r_28_2 ) , .Q( key_c_r_29_2 ) );
  DFF_X1 key_c_r_reg_29_20 (.CK( clk ) , .D( key_c_r_28_20 ) , .Q( key_c_r_29_20 ) );
  DFF_X1 key_c_r_reg_29_21 (.CK( clk ) , .D( key_c_r_28_21 ) , .Q( key_c_r_29_21 ) );
  DFF_X1 key_c_r_reg_29_22 (.CK( clk ) , .D( key_c_r_28_22 ) , .Q( key_c_r_29_22 ) );
  DFF_X1 key_c_r_reg_29_23 (.CK( clk ) , .D( key_c_r_28_23 ) , .Q( key_c_r_29_23 ) );
  DFF_X1 key_c_r_reg_29_24 (.CK( clk ) , .D( key_c_r_28_24 ) , .Q( key_c_r_29_24 ) );
  DFF_X1 key_c_r_reg_29_25 (.CK( clk ) , .D( key_c_r_28_25 ) , .Q( key_c_r_29_25 ) );
  DFF_X1 key_c_r_reg_29_26 (.CK( clk ) , .D( key_c_r_28_26 ) , .Q( key_c_r_29_26 ) );
  DFF_X1 key_c_r_reg_29_27 (.CK( clk ) , .D( key_c_r_28_27 ) , .Q( key_c_r_29_27 ) );
  DFF_X1 key_c_r_reg_29_28 (.CK( clk ) , .D( key_c_r_28_28 ) , .Q( key_c_r_29_28 ) );
  DFF_X1 key_c_r_reg_29_29 (.CK( clk ) , .D( key_c_r_28_29 ) , .Q( key_c_r_29_29 ) );
  DFF_X1 key_c_r_reg_29_3 (.CK( clk ) , .D( key_c_r_28_3 ) , .Q( key_c_r_29_3 ) );
  DFF_X1 key_c_r_reg_29_30 (.CK( clk ) , .D( key_c_r_28_30 ) , .Q( key_c_r_29_30 ) );
  DFF_X1 key_c_r_reg_29_31 (.CK( clk ) , .D( key_c_r_28_31 ) , .Q( key_c_r_29_31 ) );
  DFF_X1 key_c_r_reg_29_32 (.CK( clk ) , .D( key_c_r_28_32 ) , .Q( key_c_r_29_32 ) );
  DFF_X1 key_c_r_reg_29_33 (.CK( clk ) , .D( key_c_r_28_33 ) , .Q( key_c_r_29_33 ) );
  DFF_X1 key_c_r_reg_29_34 (.CK( clk ) , .D( key_c_r_28_34 ) , .Q( key_c_r_29_34 ) );
  DFF_X1 key_c_r_reg_29_35 (.CK( clk ) , .D( key_c_r_28_35 ) , .Q( key_c_r_29_35 ) );
  DFF_X1 key_c_r_reg_29_36 (.CK( clk ) , .D( key_c_r_28_36 ) , .Q( key_c_r_29_36 ) );
  DFF_X1 key_c_r_reg_29_37 (.CK( clk ) , .D( key_c_r_28_37 ) , .Q( key_c_r_29_37 ) );
  DFF_X1 key_c_r_reg_29_38 (.CK( clk ) , .D( key_c_r_28_38 ) , .Q( key_c_r_29_38 ) );
  DFF_X1 key_c_r_reg_29_39 (.CK( clk ) , .D( key_c_r_28_39 ) , .Q( key_c_r_29_39 ) );
  DFF_X1 key_c_r_reg_29_4 (.CK( clk ) , .D( key_c_r_28_4 ) , .Q( key_c_r_29_4 ) );
  DFF_X1 key_c_r_reg_29_40 (.CK( clk ) , .D( key_c_r_28_40 ) , .Q( key_c_r_29_40 ) );
  DFF_X1 key_c_r_reg_29_41 (.CK( clk ) , .D( key_c_r_28_41 ) , .Q( key_c_r_29_41 ) );
  DFF_X1 key_c_r_reg_29_42 (.CK( clk ) , .D( key_c_r_28_42 ) , .Q( key_c_r_29_42 ) );
  DFF_X1 key_c_r_reg_29_43 (.CK( clk ) , .D( key_c_r_28_43 ) , .Q( key_c_r_29_43 ) );
  DFF_X1 key_c_r_reg_29_44 (.CK( clk ) , .D( key_c_r_28_44 ) , .Q( key_c_r_29_44 ) );
  DFF_X1 key_c_r_reg_29_45 (.CK( clk ) , .D( key_c_r_28_45 ) , .Q( key_c_r_29_45 ) );
  DFF_X1 key_c_r_reg_29_46 (.CK( clk ) , .D( key_c_r_28_46 ) , .Q( key_c_r_29_46 ) );
  DFF_X1 key_c_r_reg_29_47 (.CK( clk ) , .D( key_c_r_28_47 ) , .Q( key_c_r_29_47 ) );
  DFF_X1 key_c_r_reg_29_48 (.CK( clk ) , .D( key_c_r_28_48 ) , .Q( key_c_r_29_48 ) );
  DFF_X1 key_c_r_reg_29_49 (.CK( clk ) , .D( key_c_r_28_49 ) , .Q( key_c_r_29_49 ) );
  DFF_X1 key_c_r_reg_29_5 (.CK( clk ) , .D( key_c_r_28_5 ) , .Q( key_c_r_29_5 ) );
  DFF_X1 key_c_r_reg_29_50 (.CK( clk ) , .D( key_c_r_28_50 ) , .Q( key_c_r_29_50 ) );
  DFF_X1 key_c_r_reg_29_51 (.CK( clk ) , .D( key_c_r_28_51 ) , .Q( key_c_r_29_51 ) );
  DFF_X1 key_c_r_reg_29_52 (.CK( clk ) , .D( key_c_r_28_52 ) , .Q( key_c_r_29_52 ) );
  DFF_X1 key_c_r_reg_29_53 (.CK( clk ) , .D( key_c_r_28_53 ) , .Q( key_c_r_29_53 ) );
  DFF_X1 key_c_r_reg_29_54 (.CK( clk ) , .D( key_c_r_28_54 ) , .Q( key_c_r_29_54 ) );
  DFF_X1 key_c_r_reg_29_55 (.CK( clk ) , .D( key_c_r_28_55 ) , .Q( key_c_r_29_55 ) );
  DFF_X1 key_c_r_reg_29_6 (.CK( clk ) , .D( key_c_r_28_6 ) , .Q( key_c_r_29_6 ) );
  DFF_X1 key_c_r_reg_29_7 (.CK( clk ) , .D( key_c_r_28_7 ) , .Q( key_c_r_29_7 ) );
  DFF_X1 key_c_r_reg_29_8 (.CK( clk ) , .D( key_c_r_28_8 ) , .Q( key_c_r_29_8 ) );
  DFF_X1 key_c_r_reg_29_9 (.CK( clk ) , .D( key_c_r_28_9 ) , .Q( key_c_r_29_9 ) );
  DFF_X1 key_c_r_reg_2_0 (.CK( clk ) , .D( key_c_r_1_0 ) , .Q( key_c_r_2_0 ) );
  DFF_X1 key_c_r_reg_2_1 (.CK( clk ) , .D( key_c_r_1_1 ) , .Q( key_c_r_2_1 ) );
  DFF_X1 key_c_r_reg_2_10 (.CK( clk ) , .D( key_c_r_1_10 ) , .Q( key_c_r_2_10 ) );
  DFF_X1 key_c_r_reg_2_11 (.CK( clk ) , .D( key_c_r_1_11 ) , .Q( key_c_r_2_11 ) );
  DFF_X1 key_c_r_reg_2_12 (.CK( clk ) , .D( key_c_r_1_12 ) , .Q( key_c_r_2_12 ) );
  DFF_X1 key_c_r_reg_2_13 (.CK( clk ) , .D( key_c_r_1_13 ) , .Q( key_c_r_2_13 ) );
  DFF_X1 key_c_r_reg_2_14 (.CK( clk ) , .D( key_c_r_1_14 ) , .Q( key_c_r_2_14 ) );
  DFF_X1 key_c_r_reg_2_15 (.CK( clk ) , .D( key_c_r_1_15 ) , .Q( key_c_r_2_15 ) );
  DFF_X1 key_c_r_reg_2_16 (.CK( clk ) , .D( key_c_r_1_16 ) , .Q( key_c_r_2_16 ) );
  DFF_X1 key_c_r_reg_2_17 (.CK( clk ) , .D( key_c_r_1_17 ) , .Q( key_c_r_2_17 ) );
  DFF_X1 key_c_r_reg_2_18 (.CK( clk ) , .D( key_c_r_1_18 ) , .Q( key_c_r_2_18 ) );
  DFF_X1 key_c_r_reg_2_19 (.CK( clk ) , .D( key_c_r_1_19 ) , .Q( key_c_r_2_19 ) );
  DFF_X1 key_c_r_reg_2_2 (.CK( clk ) , .D( key_c_r_1_2 ) , .Q( key_c_r_2_2 ) );
  DFF_X1 key_c_r_reg_2_20 (.CK( clk ) , .D( key_c_r_1_20 ) , .Q( key_c_r_2_20 ) );
  DFF_X1 key_c_r_reg_2_21 (.CK( clk ) , .D( key_c_r_1_21 ) , .Q( key_c_r_2_21 ) );
  DFF_X1 key_c_r_reg_2_22 (.CK( clk ) , .D( key_c_r_1_22 ) , .Q( key_c_r_2_22 ) );
  DFF_X1 key_c_r_reg_2_23 (.CK( clk ) , .D( key_c_r_1_23 ) , .Q( key_c_r_2_23 ) );
  DFF_X1 key_c_r_reg_2_24 (.CK( clk ) , .D( key_c_r_1_24 ) , .Q( key_c_r_2_24 ) );
  DFF_X1 key_c_r_reg_2_25 (.CK( clk ) , .D( key_c_r_1_25 ) , .Q( key_c_r_2_25 ) );
  DFF_X1 key_c_r_reg_2_26 (.CK( clk ) , .D( key_c_r_1_26 ) , .Q( key_c_r_2_26 ) );
  DFF_X1 key_c_r_reg_2_27 (.CK( clk ) , .D( key_c_r_1_27 ) , .Q( key_c_r_2_27 ) );
  DFF_X1 key_c_r_reg_2_28 (.CK( clk ) , .D( key_c_r_1_28 ) , .Q( key_c_r_2_28 ) );
  DFF_X1 key_c_r_reg_2_29 (.CK( clk ) , .D( key_c_r_1_29 ) , .Q( key_c_r_2_29 ) );
  DFF_X1 key_c_r_reg_2_3 (.CK( clk ) , .D( key_c_r_1_3 ) , .Q( key_c_r_2_3 ) );
  DFF_X1 key_c_r_reg_2_30 (.CK( clk ) , .D( key_c_r_1_30 ) , .Q( key_c_r_2_30 ) );
  DFF_X1 key_c_r_reg_2_31 (.CK( clk ) , .D( key_c_r_1_31 ) , .Q( key_c_r_2_31 ) );
  DFF_X1 key_c_r_reg_2_32 (.CK( clk ) , .D( key_c_r_1_32 ) , .Q( key_c_r_2_32 ) );
  DFF_X1 key_c_r_reg_2_33 (.CK( clk ) , .D( key_c_r_1_33 ) , .Q( key_c_r_2_33 ) );
  DFF_X1 key_c_r_reg_2_34 (.CK( clk ) , .D( key_c_r_1_34 ) , .Q( key_c_r_2_34 ) );
  DFF_X1 key_c_r_reg_2_35 (.CK( clk ) , .D( key_c_r_1_35 ) , .Q( key_c_r_2_35 ) );
  DFF_X1 key_c_r_reg_2_36 (.CK( clk ) , .D( key_c_r_1_36 ) , .Q( key_c_r_2_36 ) );
  DFF_X1 key_c_r_reg_2_37 (.CK( clk ) , .D( key_c_r_1_37 ) , .Q( key_c_r_2_37 ) );
  DFF_X1 key_c_r_reg_2_38 (.CK( clk ) , .D( key_c_r_1_38 ) , .Q( key_c_r_2_38 ) );
  DFF_X1 key_c_r_reg_2_39 (.CK( clk ) , .D( key_c_r_1_39 ) , .Q( key_c_r_2_39 ) );
  DFF_X1 key_c_r_reg_2_4 (.CK( clk ) , .D( key_c_r_1_4 ) , .Q( key_c_r_2_4 ) );
  DFF_X1 key_c_r_reg_2_40 (.CK( clk ) , .D( key_c_r_1_40 ) , .Q( key_c_r_2_40 ) );
  DFF_X1 key_c_r_reg_2_41 (.CK( clk ) , .D( key_c_r_1_41 ) , .Q( key_c_r_2_41 ) );
  DFF_X1 key_c_r_reg_2_42 (.CK( clk ) , .D( key_c_r_1_42 ) , .Q( key_c_r_2_42 ) );
  DFF_X1 key_c_r_reg_2_43 (.CK( clk ) , .D( key_c_r_1_43 ) , .Q( key_c_r_2_43 ) );
  DFF_X1 key_c_r_reg_2_44 (.CK( clk ) , .D( key_c_r_1_44 ) , .Q( key_c_r_2_44 ) );
  DFF_X1 key_c_r_reg_2_45 (.CK( clk ) , .D( key_c_r_1_45 ) , .Q( key_c_r_2_45 ) );
  DFF_X1 key_c_r_reg_2_46 (.CK( clk ) , .D( key_c_r_1_46 ) , .Q( key_c_r_2_46 ) );
  DFF_X1 key_c_r_reg_2_47 (.CK( clk ) , .D( key_c_r_1_47 ) , .Q( key_c_r_2_47 ) );
  DFF_X1 key_c_r_reg_2_48 (.CK( clk ) , .D( key_c_r_1_48 ) , .Q( key_c_r_2_48 ) );
  DFF_X1 key_c_r_reg_2_49 (.CK( clk ) , .D( key_c_r_1_49 ) , .Q( key_c_r_2_49 ) );
  DFF_X1 key_c_r_reg_2_5 (.CK( clk ) , .D( key_c_r_1_5 ) , .Q( key_c_r_2_5 ) );
  DFF_X1 key_c_r_reg_2_50 (.CK( clk ) , .D( key_c_r_1_50 ) , .Q( key_c_r_2_50 ) );
  DFF_X1 key_c_r_reg_2_51 (.CK( clk ) , .D( key_c_r_1_51 ) , .Q( key_c_r_2_51 ) );
  DFF_X1 key_c_r_reg_2_52 (.CK( clk ) , .D( key_c_r_1_52 ) , .Q( key_c_r_2_52 ) );
  DFF_X1 key_c_r_reg_2_53 (.CK( clk ) , .D( key_c_r_1_53 ) , .Q( key_c_r_2_53 ) );
  DFF_X1 key_c_r_reg_2_54 (.CK( clk ) , .D( key_c_r_1_54 ) , .Q( key_c_r_2_54 ) );
  DFF_X1 key_c_r_reg_2_55 (.CK( clk ) , .D( key_c_r_1_55 ) , .Q( key_c_r_2_55 ) );
  DFF_X1 key_c_r_reg_2_6 (.CK( clk ) , .D( key_c_r_1_6 ) , .Q( key_c_r_2_6 ) );
  DFF_X1 key_c_r_reg_2_7 (.CK( clk ) , .D( key_c_r_1_7 ) , .Q( key_c_r_2_7 ) );
  DFF_X1 key_c_r_reg_2_8 (.CK( clk ) , .D( key_c_r_1_8 ) , .Q( key_c_r_2_8 ) );
  DFF_X1 key_c_r_reg_2_9 (.CK( clk ) , .D( key_c_r_1_9 ) , .Q( key_c_r_2_9 ) );
  DFF_X1 key_c_r_reg_30_0 (.CK( clk ) , .D( key_c_r_29_0 ) , .Q( key_c_r_30_0 ) );
  DFF_X1 key_c_r_reg_30_1 (.CK( clk ) , .D( key_c_r_29_1 ) , .Q( key_c_r_30_1 ) );
  DFF_X1 key_c_r_reg_30_10 (.CK( clk ) , .D( key_c_r_29_10 ) , .Q( key_c_r_30_10 ) );
  DFF_X1 key_c_r_reg_30_11 (.CK( clk ) , .D( key_c_r_29_11 ) , .Q( key_c_r_30_11 ) );
  DFF_X1 key_c_r_reg_30_12 (.CK( clk ) , .D( key_c_r_29_12 ) , .Q( key_c_r_30_12 ) );
  DFF_X1 key_c_r_reg_30_13 (.CK( clk ) , .D( key_c_r_29_13 ) , .Q( key_c_r_30_13 ) );
  DFF_X1 key_c_r_reg_30_14 (.CK( clk ) , .D( key_c_r_29_14 ) , .Q( key_c_r_30_14 ) );
  DFF_X1 key_c_r_reg_30_15 (.CK( clk ) , .D( key_c_r_29_15 ) , .Q( key_c_r_30_15 ) );
  DFF_X1 key_c_r_reg_30_16 (.CK( clk ) , .D( key_c_r_29_16 ) , .Q( key_c_r_30_16 ) );
  DFF_X1 key_c_r_reg_30_17 (.CK( clk ) , .D( key_c_r_29_17 ) , .Q( key_c_r_30_17 ) );
  DFF_X1 key_c_r_reg_30_18 (.CK( clk ) , .D( key_c_r_29_18 ) , .Q( key_c_r_30_18 ) );
  DFF_X1 key_c_r_reg_30_19 (.CK( clk ) , .D( key_c_r_29_19 ) , .Q( key_c_r_30_19 ) );
  DFF_X1 key_c_r_reg_30_2 (.CK( clk ) , .D( key_c_r_29_2 ) , .Q( key_c_r_30_2 ) );
  DFF_X1 key_c_r_reg_30_20 (.CK( clk ) , .D( key_c_r_29_20 ) , .Q( key_c_r_30_20 ) );
  DFF_X1 key_c_r_reg_30_21 (.CK( clk ) , .D( key_c_r_29_21 ) , .Q( key_c_r_30_21 ) );
  DFF_X1 key_c_r_reg_30_22 (.CK( clk ) , .D( key_c_r_29_22 ) , .Q( key_c_r_30_22 ) );
  DFF_X1 key_c_r_reg_30_23 (.CK( clk ) , .D( key_c_r_29_23 ) , .Q( key_c_r_30_23 ) );
  DFF_X1 key_c_r_reg_30_24 (.CK( clk ) , .D( key_c_r_29_24 ) , .Q( key_c_r_30_24 ) );
  DFF_X1 key_c_r_reg_30_25 (.CK( clk ) , .D( key_c_r_29_25 ) , .Q( key_c_r_30_25 ) );
  DFF_X1 key_c_r_reg_30_26 (.CK( clk ) , .D( key_c_r_29_26 ) , .Q( key_c_r_30_26 ) );
  DFF_X1 key_c_r_reg_30_27 (.CK( clk ) , .D( key_c_r_29_27 ) , .Q( key_c_r_30_27 ) );
  DFF_X1 key_c_r_reg_30_28 (.CK( clk ) , .D( key_c_r_29_28 ) , .Q( key_c_r_30_28 ) );
  DFF_X1 key_c_r_reg_30_29 (.CK( clk ) , .D( key_c_r_29_29 ) , .Q( key_c_r_30_29 ) );
  DFF_X1 key_c_r_reg_30_3 (.CK( clk ) , .D( key_c_r_29_3 ) , .Q( key_c_r_30_3 ) );
  DFF_X1 key_c_r_reg_30_30 (.CK( clk ) , .D( key_c_r_29_30 ) , .Q( key_c_r_30_30 ) );
  DFF_X1 key_c_r_reg_30_31 (.CK( clk ) , .D( key_c_r_29_31 ) , .Q( key_c_r_30_31 ) );
  DFF_X1 key_c_r_reg_30_32 (.CK( clk ) , .D( key_c_r_29_32 ) , .Q( key_c_r_30_32 ) );
  DFF_X1 key_c_r_reg_30_33 (.CK( clk ) , .D( key_c_r_29_33 ) , .Q( key_c_r_30_33 ) );
  DFF_X1 key_c_r_reg_30_34 (.CK( clk ) , .D( key_c_r_29_34 ) , .Q( key_c_r_30_34 ) );
  DFF_X1 key_c_r_reg_30_35 (.CK( clk ) , .D( key_c_r_29_35 ) , .Q( key_c_r_30_35 ) );
  DFF_X1 key_c_r_reg_30_36 (.CK( clk ) , .D( key_c_r_29_36 ) , .Q( key_c_r_30_36 ) );
  DFF_X1 key_c_r_reg_30_37 (.CK( clk ) , .D( key_c_r_29_37 ) , .Q( key_c_r_30_37 ) );
  DFF_X1 key_c_r_reg_30_38 (.CK( clk ) , .D( key_c_r_29_38 ) , .Q( key_c_r_30_38 ) );
  DFF_X1 key_c_r_reg_30_39 (.CK( clk ) , .D( key_c_r_29_39 ) , .Q( key_c_r_30_39 ) );
  DFF_X1 key_c_r_reg_30_4 (.CK( clk ) , .D( key_c_r_29_4 ) , .Q( key_c_r_30_4 ) );
  DFF_X1 key_c_r_reg_30_40 (.CK( clk ) , .D( key_c_r_29_40 ) , .Q( key_c_r_30_40 ) );
  DFF_X1 key_c_r_reg_30_41 (.CK( clk ) , .D( key_c_r_29_41 ) , .Q( key_c_r_30_41 ) );
  DFF_X1 key_c_r_reg_30_42 (.CK( clk ) , .D( key_c_r_29_42 ) , .Q( key_c_r_30_42 ) );
  DFF_X1 key_c_r_reg_30_43 (.CK( clk ) , .D( key_c_r_29_43 ) , .Q( key_c_r_30_43 ) );
  DFF_X1 key_c_r_reg_30_44 (.CK( clk ) , .D( key_c_r_29_44 ) , .Q( key_c_r_30_44 ) );
  DFF_X1 key_c_r_reg_30_45 (.CK( clk ) , .D( key_c_r_29_45 ) , .Q( key_c_r_30_45 ) );
  DFF_X1 key_c_r_reg_30_46 (.CK( clk ) , .D( key_c_r_29_46 ) , .Q( key_c_r_30_46 ) );
  DFF_X1 key_c_r_reg_30_47 (.CK( clk ) , .D( key_c_r_29_47 ) , .Q( key_c_r_30_47 ) );
  DFF_X1 key_c_r_reg_30_48 (.CK( clk ) , .D( key_c_r_29_48 ) , .Q( key_c_r_30_48 ) );
  DFF_X1 key_c_r_reg_30_49 (.CK( clk ) , .D( key_c_r_29_49 ) , .Q( key_c_r_30_49 ) );
  DFF_X1 key_c_r_reg_30_5 (.CK( clk ) , .D( key_c_r_29_5 ) , .Q( key_c_r_30_5 ) );
  DFF_X1 key_c_r_reg_30_50 (.CK( clk ) , .D( key_c_r_29_50 ) , .Q( key_c_r_30_50 ) );
  DFF_X1 key_c_r_reg_30_51 (.CK( clk ) , .D( key_c_r_29_51 ) , .Q( key_c_r_30_51 ) );
  DFF_X1 key_c_r_reg_30_52 (.CK( clk ) , .D( key_c_r_29_52 ) , .Q( key_c_r_30_52 ) );
  DFF_X1 key_c_r_reg_30_53 (.CK( clk ) , .D( key_c_r_29_53 ) , .Q( key_c_r_30_53 ) );
  DFF_X1 key_c_r_reg_30_54 (.CK( clk ) , .D( key_c_r_29_54 ) , .Q( key_c_r_30_54 ) );
  DFF_X1 key_c_r_reg_30_55 (.CK( clk ) , .D( key_c_r_29_55 ) , .Q( key_c_r_30_55 ) );
  DFF_X1 key_c_r_reg_30_6 (.CK( clk ) , .D( key_c_r_29_6 ) , .Q( key_c_r_30_6 ) );
  DFF_X1 key_c_r_reg_30_7 (.CK( clk ) , .D( key_c_r_29_7 ) , .Q( key_c_r_30_7 ) );
  DFF_X1 key_c_r_reg_30_8 (.CK( clk ) , .D( key_c_r_29_8 ) , .Q( key_c_r_30_8 ) );
  DFF_X1 key_c_r_reg_30_9 (.CK( clk ) , .D( key_c_r_29_9 ) , .Q( key_c_r_30_9 ) );
  DFF_X1 key_c_r_reg_31_0 (.CK( clk ) , .D( key_c_r_30_0 ) , .Q( key_c_r_31_0 ) );
  DFF_X1 key_c_r_reg_31_1 (.CK( clk ) , .D( key_c_r_30_1 ) , .Q( key_c_r_31_1 ) );
  DFF_X1 key_c_r_reg_31_10 (.CK( clk ) , .D( key_c_r_30_10 ) , .Q( key_c_r_31_10 ) );
  DFF_X1 key_c_r_reg_31_11 (.CK( clk ) , .D( key_c_r_30_11 ) , .Q( key_c_r_31_11 ) );
  DFF_X1 key_c_r_reg_31_12 (.CK( clk ) , .D( key_c_r_30_12 ) , .Q( key_c_r_31_12 ) );
  DFF_X1 key_c_r_reg_31_13 (.CK( clk ) , .D( key_c_r_30_13 ) , .Q( key_c_r_31_13 ) );
  DFF_X1 key_c_r_reg_31_14 (.CK( clk ) , .D( key_c_r_30_14 ) , .Q( key_c_r_31_14 ) );
  DFF_X1 key_c_r_reg_31_15 (.CK( clk ) , .D( key_c_r_30_15 ) , .Q( key_c_r_31_15 ) );
  DFF_X1 key_c_r_reg_31_16 (.CK( clk ) , .D( key_c_r_30_16 ) , .Q( key_c_r_31_16 ) );
  DFF_X1 key_c_r_reg_31_17 (.CK( clk ) , .D( key_c_r_30_17 ) , .Q( key_c_r_31_17 ) );
  DFF_X1 key_c_r_reg_31_18 (.CK( clk ) , .D( key_c_r_30_18 ) , .Q( key_c_r_31_18 ) );
  DFF_X1 key_c_r_reg_31_19 (.CK( clk ) , .D( key_c_r_30_19 ) , .Q( key_c_r_31_19 ) );
  DFF_X1 key_c_r_reg_31_2 (.CK( clk ) , .D( key_c_r_30_2 ) , .Q( key_c_r_31_2 ) );
  DFF_X1 key_c_r_reg_31_20 (.CK( clk ) , .D( key_c_r_30_20 ) , .Q( key_c_r_31_20 ) );
  DFF_X1 key_c_r_reg_31_21 (.CK( clk ) , .D( key_c_r_30_21 ) , .Q( key_c_r_31_21 ) );
  DFF_X1 key_c_r_reg_31_22 (.CK( clk ) , .D( key_c_r_30_22 ) , .Q( key_c_r_31_22 ) );
  DFF_X1 key_c_r_reg_31_23 (.CK( clk ) , .D( key_c_r_30_23 ) , .Q( key_c_r_31_23 ) );
  DFF_X1 key_c_r_reg_31_24 (.CK( clk ) , .D( key_c_r_30_24 ) , .Q( key_c_r_31_24 ) );
  DFF_X1 key_c_r_reg_31_25 (.CK( clk ) , .D( key_c_r_30_25 ) , .Q( key_c_r_31_25 ) );
  DFF_X1 key_c_r_reg_31_26 (.CK( clk ) , .D( key_c_r_30_26 ) , .Q( key_c_r_31_26 ) );
  DFF_X1 key_c_r_reg_31_27 (.CK( clk ) , .D( key_c_r_30_27 ) , .Q( key_c_r_31_27 ) );
  DFF_X1 key_c_r_reg_31_28 (.CK( clk ) , .D( key_c_r_30_28 ) , .Q( key_c_r_31_28 ) );
  DFF_X1 key_c_r_reg_31_29 (.CK( clk ) , .D( key_c_r_30_29 ) , .Q( key_c_r_31_29 ) );
  DFF_X1 key_c_r_reg_31_3 (.CK( clk ) , .D( key_c_r_30_3 ) , .Q( key_c_r_31_3 ) );
  DFF_X1 key_c_r_reg_31_30 (.CK( clk ) , .D( key_c_r_30_30 ) , .Q( key_c_r_31_30 ) );
  DFF_X1 key_c_r_reg_31_31 (.CK( clk ) , .D( key_c_r_30_31 ) , .Q( key_c_r_31_31 ) );
  DFF_X1 key_c_r_reg_31_32 (.CK( clk ) , .D( key_c_r_30_32 ) , .Q( key_c_r_31_32 ) );
  DFF_X1 key_c_r_reg_31_33 (.CK( clk ) , .D( key_c_r_30_33 ) , .Q( key_c_r_31_33 ) );
  DFF_X1 key_c_r_reg_31_34 (.CK( clk ) , .D( key_c_r_30_34 ) , .Q( key_c_r_31_34 ) );
  DFF_X1 key_c_r_reg_31_35 (.CK( clk ) , .D( key_c_r_30_35 ) , .Q( key_c_r_31_35 ) );
  DFF_X1 key_c_r_reg_31_36 (.CK( clk ) , .D( key_c_r_30_36 ) , .Q( key_c_r_31_36 ) );
  DFF_X1 key_c_r_reg_31_37 (.CK( clk ) , .D( key_c_r_30_37 ) , .Q( key_c_r_31_37 ) );
  DFF_X1 key_c_r_reg_31_38 (.CK( clk ) , .D( key_c_r_30_38 ) , .Q( key_c_r_31_38 ) );
  DFF_X1 key_c_r_reg_31_39 (.CK( clk ) , .D( key_c_r_30_39 ) , .Q( key_c_r_31_39 ) );
  DFF_X1 key_c_r_reg_31_4 (.CK( clk ) , .D( key_c_r_30_4 ) , .Q( key_c_r_31_4 ) );
  DFF_X1 key_c_r_reg_31_40 (.CK( clk ) , .D( key_c_r_30_40 ) , .Q( key_c_r_31_40 ) );
  DFF_X1 key_c_r_reg_31_41 (.CK( clk ) , .D( key_c_r_30_41 ) , .Q( key_c_r_31_41 ) );
  DFF_X1 key_c_r_reg_31_42 (.CK( clk ) , .D( key_c_r_30_42 ) , .Q( key_c_r_31_42 ) );
  DFF_X1 key_c_r_reg_31_43 (.CK( clk ) , .D( key_c_r_30_43 ) , .Q( key_c_r_31_43 ) );
  DFF_X1 key_c_r_reg_31_44 (.CK( clk ) , .D( key_c_r_30_44 ) , .Q( key_c_r_31_44 ) );
  DFF_X1 key_c_r_reg_31_45 (.CK( clk ) , .D( key_c_r_30_45 ) , .Q( key_c_r_31_45 ) );
  DFF_X1 key_c_r_reg_31_46 (.CK( clk ) , .D( key_c_r_30_46 ) , .Q( key_c_r_31_46 ) );
  DFF_X1 key_c_r_reg_31_47 (.CK( clk ) , .D( key_c_r_30_47 ) , .Q( key_c_r_31_47 ) );
  DFF_X1 key_c_r_reg_31_48 (.CK( clk ) , .D( key_c_r_30_48 ) , .Q( key_c_r_31_48 ) );
  DFF_X1 key_c_r_reg_31_49 (.CK( clk ) , .D( key_c_r_30_49 ) , .Q( key_c_r_31_49 ) );
  DFF_X1 key_c_r_reg_31_5 (.CK( clk ) , .D( key_c_r_30_5 ) , .Q( key_c_r_31_5 ) );
  DFF_X1 key_c_r_reg_31_50 (.CK( clk ) , .D( key_c_r_30_50 ) , .Q( key_c_r_31_50 ) );
  DFF_X1 key_c_r_reg_31_51 (.CK( clk ) , .D( key_c_r_30_51 ) , .Q( key_c_r_31_51 ) );
  DFF_X1 key_c_r_reg_31_52 (.CK( clk ) , .D( key_c_r_30_52 ) , .Q( key_c_r_31_52 ) );
  DFF_X1 key_c_r_reg_31_53 (.CK( clk ) , .D( key_c_r_30_53 ) , .Q( key_c_r_31_53 ) );
  DFF_X1 key_c_r_reg_31_54 (.CK( clk ) , .D( key_c_r_30_54 ) , .Q( key_c_r_31_54 ) );
  DFF_X1 key_c_r_reg_31_55 (.CK( clk ) , .D( key_c_r_30_55 ) , .Q( key_c_r_31_55 ) );
  DFF_X1 key_c_r_reg_31_6 (.CK( clk ) , .D( key_c_r_30_6 ) , .Q( key_c_r_31_6 ) );
  DFF_X1 key_c_r_reg_31_7 (.CK( clk ) , .D( key_c_r_30_7 ) , .Q( key_c_r_31_7 ) );
  DFF_X1 key_c_r_reg_31_8 (.CK( clk ) , .D( key_c_r_30_8 ) , .Q( key_c_r_31_8 ) );
  DFF_X1 key_c_r_reg_31_9 (.CK( clk ) , .D( key_c_r_30_9 ) , .Q( key_c_r_31_9 ) );
  DFF_X1 key_c_r_reg_32_0 (.CK( clk ) , .D( key_c_r_31_0 ) , .Q( key_c_r_32_0 ) );
  DFF_X1 key_c_r_reg_32_1 (.CK( clk ) , .D( key_c_r_31_1 ) , .Q( key_c_r_32_1 ) );
  DFF_X1 key_c_r_reg_32_10 (.CK( clk ) , .D( key_c_r_31_10 ) , .Q( key_c_r_32_10 ) );
  DFF_X1 key_c_r_reg_32_11 (.CK( clk ) , .D( key_c_r_31_11 ) , .Q( key_c_r_32_11 ) );
  DFF_X1 key_c_r_reg_32_12 (.CK( clk ) , .D( key_c_r_31_12 ) , .Q( key_c_r_32_12 ) );
  DFF_X1 key_c_r_reg_32_13 (.CK( clk ) , .D( key_c_r_31_13 ) , .Q( key_c_r_32_13 ) );
  DFF_X1 key_c_r_reg_32_14 (.CK( clk ) , .D( key_c_r_31_14 ) , .Q( key_c_r_32_14 ) );
  DFF_X1 key_c_r_reg_32_15 (.CK( clk ) , .D( key_c_r_31_15 ) , .Q( key_c_r_32_15 ) );
  DFF_X1 key_c_r_reg_32_16 (.CK( clk ) , .D( key_c_r_31_16 ) , .Q( key_c_r_32_16 ) );
  DFF_X1 key_c_r_reg_32_17 (.CK( clk ) , .D( key_c_r_31_17 ) , .Q( key_c_r_32_17 ) );
  DFF_X1 key_c_r_reg_32_18 (.CK( clk ) , .D( key_c_r_31_18 ) , .Q( key_c_r_32_18 ) );
  DFF_X1 key_c_r_reg_32_19 (.CK( clk ) , .D( key_c_r_31_19 ) , .Q( key_c_r_32_19 ) );
  DFF_X1 key_c_r_reg_32_2 (.CK( clk ) , .D( key_c_r_31_2 ) , .Q( key_c_r_32_2 ) );
  DFF_X1 key_c_r_reg_32_20 (.CK( clk ) , .D( key_c_r_31_20 ) , .Q( key_c_r_32_20 ) );
  DFF_X1 key_c_r_reg_32_21 (.CK( clk ) , .D( key_c_r_31_21 ) , .Q( key_c_r_32_21 ) );
  DFF_X1 key_c_r_reg_32_22 (.CK( clk ) , .D( key_c_r_31_22 ) , .Q( key_c_r_32_22 ) );
  DFF_X1 key_c_r_reg_32_23 (.CK( clk ) , .D( key_c_r_31_23 ) , .Q( key_c_r_32_23 ) );
  DFF_X1 key_c_r_reg_32_24 (.CK( clk ) , .D( key_c_r_31_24 ) , .Q( key_c_r_32_24 ) );
  DFF_X1 key_c_r_reg_32_25 (.CK( clk ) , .D( key_c_r_31_25 ) , .Q( key_c_r_32_25 ) );
  DFF_X1 key_c_r_reg_32_26 (.CK( clk ) , .D( key_c_r_31_26 ) , .Q( key_c_r_32_26 ) );
  DFF_X1 key_c_r_reg_32_27 (.CK( clk ) , .D( key_c_r_31_27 ) , .Q( key_c_r_32_27 ) );
  DFF_X1 key_c_r_reg_32_28 (.CK( clk ) , .D( key_c_r_31_28 ) , .Q( key_c_r_32_28 ) );
  DFF_X1 key_c_r_reg_32_29 (.CK( clk ) , .D( key_c_r_31_29 ) , .Q( key_c_r_32_29 ) );
  DFF_X1 key_c_r_reg_32_3 (.CK( clk ) , .D( key_c_r_31_3 ) , .Q( key_c_r_32_3 ) );
  DFF_X1 key_c_r_reg_32_30 (.CK( clk ) , .D( key_c_r_31_30 ) , .Q( key_c_r_32_30 ) );
  DFF_X1 key_c_r_reg_32_31 (.CK( clk ) , .D( key_c_r_31_31 ) , .Q( key_c_r_32_31 ) );
  DFF_X1 key_c_r_reg_32_32 (.CK( clk ) , .D( key_c_r_31_32 ) , .Q( key_c_r_32_32 ) );
  DFF_X1 key_c_r_reg_32_33 (.CK( clk ) , .D( key_c_r_31_33 ) , .Q( key_c_r_32_33 ) );
  DFF_X1 key_c_r_reg_32_34 (.CK( clk ) , .D( key_c_r_31_34 ) , .Q( key_c_r_32_34 ) );
  DFF_X1 key_c_r_reg_32_35 (.CK( clk ) , .D( key_c_r_31_35 ) , .Q( key_c_r_32_35 ) );
  DFF_X1 key_c_r_reg_32_36 (.CK( clk ) , .D( key_c_r_31_36 ) , .Q( key_c_r_32_36 ) );
  DFF_X1 key_c_r_reg_32_37 (.CK( clk ) , .D( key_c_r_31_37 ) , .Q( key_c_r_32_37 ) );
  DFF_X1 key_c_r_reg_32_38 (.CK( clk ) , .D( key_c_r_31_38 ) , .Q( key_c_r_32_38 ) );
  DFF_X1 key_c_r_reg_32_39 (.CK( clk ) , .D( key_c_r_31_39 ) , .Q( key_c_r_32_39 ) );
  DFF_X1 key_c_r_reg_32_4 (.CK( clk ) , .D( key_c_r_31_4 ) , .Q( key_c_r_32_4 ) );
  DFF_X1 key_c_r_reg_32_40 (.CK( clk ) , .D( key_c_r_31_40 ) , .Q( key_c_r_32_40 ) );
  DFF_X1 key_c_r_reg_32_41 (.CK( clk ) , .D( key_c_r_31_41 ) , .Q( key_c_r_32_41 ) );
  DFF_X1 key_c_r_reg_32_42 (.CK( clk ) , .D( key_c_r_31_42 ) , .Q( key_c_r_32_42 ) );
  DFF_X1 key_c_r_reg_32_43 (.CK( clk ) , .D( key_c_r_31_43 ) , .Q( key_c_r_32_43 ) );
  DFF_X1 key_c_r_reg_32_44 (.CK( clk ) , .D( key_c_r_31_44 ) , .Q( key_c_r_32_44 ) );
  DFF_X1 key_c_r_reg_32_45 (.CK( clk ) , .D( key_c_r_31_45 ) , .Q( key_c_r_32_45 ) );
  DFF_X1 key_c_r_reg_32_46 (.CK( clk ) , .D( key_c_r_31_46 ) , .Q( key_c_r_32_46 ) );
  DFF_X1 key_c_r_reg_32_47 (.CK( clk ) , .D( key_c_r_31_47 ) , .Q( key_c_r_32_47 ) );
  DFF_X1 key_c_r_reg_32_48 (.CK( clk ) , .D( key_c_r_31_48 ) , .Q( key_c_r_32_48 ) );
  DFF_X1 key_c_r_reg_32_49 (.CK( clk ) , .D( key_c_r_31_49 ) , .Q( key_c_r_32_49 ) );
  DFF_X1 key_c_r_reg_32_5 (.CK( clk ) , .D( key_c_r_31_5 ) , .Q( key_c_r_32_5 ) );
  DFF_X1 key_c_r_reg_32_50 (.CK( clk ) , .D( key_c_r_31_50 ) , .Q( key_c_r_32_50 ) );
  DFF_X1 key_c_r_reg_32_51 (.CK( clk ) , .D( key_c_r_31_51 ) , .Q( key_c_r_32_51 ) );
  DFF_X1 key_c_r_reg_32_52 (.CK( clk ) , .D( key_c_r_31_52 ) , .Q( key_c_r_32_52 ) );
  DFF_X1 key_c_r_reg_32_53 (.CK( clk ) , .D( key_c_r_31_53 ) , .Q( key_c_r_32_53 ) );
  DFF_X1 key_c_r_reg_32_54 (.CK( clk ) , .D( key_c_r_31_54 ) , .Q( key_c_r_32_54 ) );
  DFF_X1 key_c_r_reg_32_55 (.CK( clk ) , .D( key_c_r_31_55 ) , .Q( key_c_r_32_55 ) );
  DFF_X1 key_c_r_reg_32_6 (.CK( clk ) , .D( key_c_r_31_6 ) , .Q( key_c_r_32_6 ) );
  DFF_X1 key_c_r_reg_32_7 (.CK( clk ) , .D( key_c_r_31_7 ) , .Q( key_c_r_32_7 ) );
  DFF_X1 key_c_r_reg_32_8 (.CK( clk ) , .D( key_c_r_31_8 ) , .Q( key_c_r_32_8 ) );
  DFF_X1 key_c_r_reg_32_9 (.CK( clk ) , .D( key_c_r_31_9 ) , .Q( key_c_r_32_9 ) );
  DFF_X1 key_c_r_reg_33_0 (.CK( clk ) , .D( key_c_r_32_0 ) , .Q( key_c_r_33_0 ) );
  DFF_X1 key_c_r_reg_33_1 (.CK( clk ) , .D( key_c_r_32_1 ) , .Q( key_c_r_33_1 ) );
  DFF_X1 key_c_r_reg_33_10 (.CK( clk ) , .D( key_c_r_32_10 ) , .Q( key_c_r_33_10 ) );
  DFF_X1 key_c_r_reg_33_11 (.CK( clk ) , .D( key_c_r_32_11 ) , .Q( key_c_r_33_11 ) );
  DFF_X1 key_c_r_reg_33_12 (.CK( clk ) , .D( key_c_r_32_12 ) , .Q( key_c_r_33_12 ) );
  DFF_X1 key_c_r_reg_33_13 (.CK( clk ) , .D( key_c_r_32_13 ) , .Q( key_c_r_33_13 ) );
  DFF_X1 key_c_r_reg_33_14 (.CK( clk ) , .D( key_c_r_32_14 ) , .Q( key_c_r_33_14 ) );
  DFF_X1 key_c_r_reg_33_15 (.CK( clk ) , .D( key_c_r_32_15 ) , .Q( key_c_r_33_15 ) );
  DFF_X1 key_c_r_reg_33_16 (.CK( clk ) , .D( key_c_r_32_16 ) , .Q( key_c_r_33_16 ) );
  DFF_X1 key_c_r_reg_33_17 (.CK( clk ) , .D( key_c_r_32_17 ) , .Q( key_c_r_33_17 ) );
  DFF_X1 key_c_r_reg_33_18 (.CK( clk ) , .D( key_c_r_32_18 ) , .Q( key_c_r_33_18 ) );
  DFF_X1 key_c_r_reg_33_19 (.CK( clk ) , .D( key_c_r_32_19 ) , .Q( key_c_r_33_19 ) );
  DFF_X1 key_c_r_reg_33_2 (.CK( clk ) , .D( key_c_r_32_2 ) , .Q( key_c_r_33_2 ) );
  DFF_X1 key_c_r_reg_33_20 (.CK( clk ) , .D( key_c_r_32_20 ) , .Q( key_c_r_33_20 ) );
  DFF_X1 key_c_r_reg_33_21 (.CK( clk ) , .D( key_c_r_32_21 ) , .Q( key_c_r_33_21 ) );
  DFF_X1 key_c_r_reg_33_22 (.CK( clk ) , .D( key_c_r_32_22 ) , .Q( key_c_r_33_22 ) );
  DFF_X1 key_c_r_reg_33_23 (.CK( clk ) , .D( key_c_r_32_23 ) , .Q( key_c_r_33_23 ) );
  DFF_X1 key_c_r_reg_33_24 (.CK( clk ) , .D( key_c_r_32_24 ) , .Q( key_c_r_33_24 ) );
  DFF_X1 key_c_r_reg_33_25 (.CK( clk ) , .D( key_c_r_32_25 ) , .Q( key_c_r_33_25 ) );
  DFF_X1 key_c_r_reg_33_26 (.CK( clk ) , .D( key_c_r_32_26 ) , .Q( key_c_r_33_26 ) );
  DFF_X1 key_c_r_reg_33_27 (.CK( clk ) , .D( key_c_r_32_27 ) , .Q( key_c_r_33_27 ) );
  DFF_X1 key_c_r_reg_33_28 (.CK( clk ) , .D( key_c_r_32_28 ) , .Q( key_c_r_33_28 ) );
  DFF_X1 key_c_r_reg_33_29 (.CK( clk ) , .D( key_c_r_32_29 ) , .Q( key_c_r_33_29 ) );
  DFF_X1 key_c_r_reg_33_3 (.CK( clk ) , .D( key_c_r_32_3 ) , .Q( key_c_r_33_3 ) );
  DFF_X1 key_c_r_reg_33_30 (.CK( clk ) , .D( key_c_r_32_30 ) , .Q( key_c_r_33_30 ) );
  DFF_X1 key_c_r_reg_33_31 (.CK( clk ) , .D( key_c_r_32_31 ) , .Q( key_c_r_33_31 ) );
  DFF_X1 key_c_r_reg_33_32 (.CK( clk ) , .D( key_c_r_32_32 ) , .Q( key_c_r_33_32 ) );
  DFF_X1 key_c_r_reg_33_33 (.CK( clk ) , .D( key_c_r_32_33 ) , .Q( key_c_r_33_33 ) );
  DFF_X1 key_c_r_reg_33_34 (.CK( clk ) , .D( key_c_r_32_34 ) , .Q( key_c_r_33_34 ) );
  DFF_X1 key_c_r_reg_33_35 (.CK( clk ) , .D( key_c_r_32_35 ) , .Q( key_c_r_33_35 ) );
  DFF_X1 key_c_r_reg_33_36 (.CK( clk ) , .D( key_c_r_32_36 ) , .Q( key_c_r_33_36 ) );
  DFF_X1 key_c_r_reg_33_37 (.CK( clk ) , .D( key_c_r_32_37 ) , .Q( key_c_r_33_37 ) );
  DFF_X1 key_c_r_reg_33_38 (.CK( clk ) , .D( key_c_r_32_38 ) , .Q( key_c_r_33_38 ) );
  DFF_X1 key_c_r_reg_33_39 (.CK( clk ) , .D( key_c_r_32_39 ) , .Q( key_c_r_33_39 ) );
  DFF_X1 key_c_r_reg_33_4 (.CK( clk ) , .D( key_c_r_32_4 ) , .Q( key_c_r_33_4 ) );
  DFF_X1 key_c_r_reg_33_40 (.CK( clk ) , .D( key_c_r_32_40 ) , .Q( key_c_r_33_40 ) );
  DFF_X1 key_c_r_reg_33_41 (.CK( clk ) , .D( key_c_r_32_41 ) , .Q( key_c_r_33_41 ) );
  DFF_X1 key_c_r_reg_33_42 (.CK( clk ) , .D( key_c_r_32_42 ) , .Q( key_c_r_33_42 ) );
  DFF_X1 key_c_r_reg_33_43 (.CK( clk ) , .D( key_c_r_32_43 ) , .Q( key_c_r_33_43 ) );
  DFF_X1 key_c_r_reg_33_44 (.CK( clk ) , .D( key_c_r_32_44 ) , .Q( key_c_r_33_44 ) );
  DFF_X1 key_c_r_reg_33_45 (.CK( clk ) , .D( key_c_r_32_45 ) , .Q( key_c_r_33_45 ) );
  DFF_X1 key_c_r_reg_33_46 (.CK( clk ) , .D( key_c_r_32_46 ) , .Q( key_c_r_33_46 ) );
  DFF_X1 key_c_r_reg_33_47 (.CK( clk ) , .D( key_c_r_32_47 ) , .Q( key_c_r_33_47 ) );
  DFF_X1 key_c_r_reg_33_48 (.CK( clk ) , .D( key_c_r_32_48 ) , .Q( key_c_r_33_48 ) );
  DFF_X1 key_c_r_reg_33_49 (.CK( clk ) , .D( key_c_r_32_49 ) , .Q( key_c_r_33_49 ) );
  DFF_X1 key_c_r_reg_33_5 (.CK( clk ) , .D( key_c_r_32_5 ) , .Q( key_c_r_33_5 ) );
  DFF_X1 key_c_r_reg_33_50 (.CK( clk ) , .D( key_c_r_32_50 ) , .Q( key_c_r_33_50 ) );
  DFF_X1 key_c_r_reg_33_51 (.CK( clk ) , .D( key_c_r_32_51 ) , .Q( key_c_r_33_51 ) );
  DFF_X1 key_c_r_reg_33_52 (.CK( clk ) , .D( key_c_r_32_52 ) , .Q( key_c_r_33_52 ) );
  DFF_X1 key_c_r_reg_33_53 (.CK( clk ) , .D( key_c_r_32_53 ) , .Q( key_c_r_33_53 ) );
  DFF_X1 key_c_r_reg_33_54 (.CK( clk ) , .D( key_c_r_32_54 ) , .Q( key_c_r_33_54 ) );
  DFF_X1 key_c_r_reg_33_55 (.CK( clk ) , .D( key_c_r_32_55 ) , .Q( key_c_r_33_55 ) );
  DFF_X1 key_c_r_reg_33_6 (.CK( clk ) , .D( key_c_r_32_6 ) , .Q( key_c_r_33_6 ) );
  DFF_X1 key_c_r_reg_33_7 (.CK( clk ) , .D( key_c_r_32_7 ) , .Q( key_c_r_33_7 ) );
  DFF_X1 key_c_r_reg_33_8 (.CK( clk ) , .D( key_c_r_32_8 ) , .Q( key_c_r_33_8 ) );
  DFF_X1 key_c_r_reg_33_9 (.CK( clk ) , .D( key_c_r_32_9 ) , .Q( key_c_r_33_9 ) );
  DFF_X1 key_c_r_reg_3_0 (.CK( clk ) , .D( key_c_r_2_0 ) , .Q( key_c_r_3_0 ) );
  DFF_X1 key_c_r_reg_3_1 (.CK( clk ) , .D( key_c_r_2_1 ) , .Q( key_c_r_3_1 ) );
  DFF_X1 key_c_r_reg_3_10 (.CK( clk ) , .D( key_c_r_2_10 ) , .Q( key_c_r_3_10 ) );
  DFF_X1 key_c_r_reg_3_11 (.CK( clk ) , .D( key_c_r_2_11 ) , .Q( key_c_r_3_11 ) );
  DFF_X1 key_c_r_reg_3_12 (.CK( clk ) , .D( key_c_r_2_12 ) , .Q( key_c_r_3_12 ) );
  DFF_X1 key_c_r_reg_3_13 (.CK( clk ) , .D( key_c_r_2_13 ) , .Q( key_c_r_3_13 ) );
  DFF_X1 key_c_r_reg_3_14 (.CK( clk ) , .D( key_c_r_2_14 ) , .Q( key_c_r_3_14 ) );
  DFF_X1 key_c_r_reg_3_15 (.CK( clk ) , .D( key_c_r_2_15 ) , .Q( key_c_r_3_15 ) );
  DFF_X1 key_c_r_reg_3_16 (.CK( clk ) , .D( key_c_r_2_16 ) , .Q( key_c_r_3_16 ) );
  DFF_X1 key_c_r_reg_3_17 (.CK( clk ) , .D( key_c_r_2_17 ) , .Q( key_c_r_3_17 ) );
  DFF_X1 key_c_r_reg_3_18 (.CK( clk ) , .D( key_c_r_2_18 ) , .Q( key_c_r_3_18 ) );
  DFF_X1 key_c_r_reg_3_19 (.CK( clk ) , .D( key_c_r_2_19 ) , .Q( key_c_r_3_19 ) );
  DFF_X1 key_c_r_reg_3_2 (.CK( clk ) , .D( key_c_r_2_2 ) , .Q( key_c_r_3_2 ) );
  DFF_X1 key_c_r_reg_3_20 (.CK( clk ) , .D( key_c_r_2_20 ) , .Q( key_c_r_3_20 ) );
  DFF_X1 key_c_r_reg_3_21 (.CK( clk ) , .D( key_c_r_2_21 ) , .Q( key_c_r_3_21 ) );
  DFF_X1 key_c_r_reg_3_22 (.CK( clk ) , .D( key_c_r_2_22 ) , .Q( key_c_r_3_22 ) );
  DFF_X1 key_c_r_reg_3_23 (.CK( clk ) , .D( key_c_r_2_23 ) , .Q( key_c_r_3_23 ) );
  DFF_X1 key_c_r_reg_3_24 (.CK( clk ) , .D( key_c_r_2_24 ) , .Q( key_c_r_3_24 ) );
  DFF_X1 key_c_r_reg_3_25 (.CK( clk ) , .D( key_c_r_2_25 ) , .Q( key_c_r_3_25 ) );
  DFF_X1 key_c_r_reg_3_26 (.CK( clk ) , .D( key_c_r_2_26 ) , .Q( key_c_r_3_26 ) );
  DFF_X1 key_c_r_reg_3_27 (.CK( clk ) , .D( key_c_r_2_27 ) , .Q( key_c_r_3_27 ) );
  DFF_X1 key_c_r_reg_3_28 (.CK( clk ) , .D( key_c_r_2_28 ) , .Q( key_c_r_3_28 ) );
  DFF_X1 key_c_r_reg_3_29 (.CK( clk ) , .D( key_c_r_2_29 ) , .Q( key_c_r_3_29 ) );
  DFF_X1 key_c_r_reg_3_3 (.CK( clk ) , .D( key_c_r_2_3 ) , .Q( key_c_r_3_3 ) );
  DFF_X1 key_c_r_reg_3_30 (.CK( clk ) , .D( key_c_r_2_30 ) , .Q( key_c_r_3_30 ) );
  DFF_X1 key_c_r_reg_3_31 (.CK( clk ) , .D( key_c_r_2_31 ) , .Q( key_c_r_3_31 ) );
  DFF_X1 key_c_r_reg_3_32 (.CK( clk ) , .D( key_c_r_2_32 ) , .Q( key_c_r_3_32 ) );
  DFF_X1 key_c_r_reg_3_33 (.CK( clk ) , .D( key_c_r_2_33 ) , .Q( key_c_r_3_33 ) );
  DFF_X1 key_c_r_reg_3_34 (.CK( clk ) , .D( key_c_r_2_34 ) , .Q( key_c_r_3_34 ) );
  DFF_X1 key_c_r_reg_3_35 (.CK( clk ) , .D( key_c_r_2_35 ) , .Q( key_c_r_3_35 ) );
  DFF_X1 key_c_r_reg_3_36 (.CK( clk ) , .D( key_c_r_2_36 ) , .Q( key_c_r_3_36 ) );
  DFF_X1 key_c_r_reg_3_37 (.CK( clk ) , .D( key_c_r_2_37 ) , .Q( key_c_r_3_37 ) );
  DFF_X1 key_c_r_reg_3_38 (.CK( clk ) , .D( key_c_r_2_38 ) , .Q( key_c_r_3_38 ) );
  DFF_X1 key_c_r_reg_3_39 (.CK( clk ) , .D( key_c_r_2_39 ) , .Q( key_c_r_3_39 ) );
  DFF_X1 key_c_r_reg_3_4 (.CK( clk ) , .D( key_c_r_2_4 ) , .Q( key_c_r_3_4 ) );
  DFF_X1 key_c_r_reg_3_40 (.CK( clk ) , .D( key_c_r_2_40 ) , .Q( key_c_r_3_40 ) );
  DFF_X1 key_c_r_reg_3_41 (.CK( clk ) , .D( key_c_r_2_41 ) , .Q( key_c_r_3_41 ) );
  DFF_X1 key_c_r_reg_3_42 (.CK( clk ) , .D( key_c_r_2_42 ) , .Q( key_c_r_3_42 ) );
  DFF_X1 key_c_r_reg_3_43 (.CK( clk ) , .D( key_c_r_2_43 ) , .Q( key_c_r_3_43 ) );
  DFF_X1 key_c_r_reg_3_44 (.CK( clk ) , .D( key_c_r_2_44 ) , .Q( key_c_r_3_44 ) );
  DFF_X1 key_c_r_reg_3_45 (.CK( clk ) , .D( key_c_r_2_45 ) , .Q( key_c_r_3_45 ) );
  DFF_X1 key_c_r_reg_3_46 (.CK( clk ) , .D( key_c_r_2_46 ) , .Q( key_c_r_3_46 ) );
  DFF_X1 key_c_r_reg_3_47 (.CK( clk ) , .D( key_c_r_2_47 ) , .Q( key_c_r_3_47 ) );
  DFF_X1 key_c_r_reg_3_48 (.CK( clk ) , .D( key_c_r_2_48 ) , .Q( key_c_r_3_48 ) );
  DFF_X1 key_c_r_reg_3_49 (.CK( clk ) , .D( key_c_r_2_49 ) , .Q( key_c_r_3_49 ) );
  DFF_X1 key_c_r_reg_3_5 (.CK( clk ) , .D( key_c_r_2_5 ) , .Q( key_c_r_3_5 ) );
  DFF_X1 key_c_r_reg_3_50 (.CK( clk ) , .D( key_c_r_2_50 ) , .Q( key_c_r_3_50 ) );
  DFF_X1 key_c_r_reg_3_51 (.CK( clk ) , .D( key_c_r_2_51 ) , .Q( key_c_r_3_51 ) );
  DFF_X1 key_c_r_reg_3_52 (.CK( clk ) , .D( key_c_r_2_52 ) , .Q( key_c_r_3_52 ) );
  DFF_X1 key_c_r_reg_3_53 (.CK( clk ) , .D( key_c_r_2_53 ) , .Q( key_c_r_3_53 ) );
  DFF_X1 key_c_r_reg_3_54 (.CK( clk ) , .D( key_c_r_2_54 ) , .Q( key_c_r_3_54 ) );
  DFF_X1 key_c_r_reg_3_55 (.CK( clk ) , .D( key_c_r_2_55 ) , .Q( key_c_r_3_55 ) );
  DFF_X1 key_c_r_reg_3_6 (.CK( clk ) , .D( key_c_r_2_6 ) , .Q( key_c_r_3_6 ) );
  DFF_X1 key_c_r_reg_3_7 (.CK( clk ) , .D( key_c_r_2_7 ) , .Q( key_c_r_3_7 ) );
  DFF_X1 key_c_r_reg_3_8 (.CK( clk ) , .D( key_c_r_2_8 ) , .Q( key_c_r_3_8 ) );
  DFF_X1 key_c_r_reg_3_9 (.CK( clk ) , .D( key_c_r_2_9 ) , .Q( key_c_r_3_9 ) );
  DFF_X1 key_c_r_reg_4_0 (.CK( clk ) , .D( key_c_r_3_0 ) , .Q( key_c_r_4_0 ) );
  DFF_X1 key_c_r_reg_4_1 (.CK( clk ) , .D( key_c_r_3_1 ) , .Q( key_c_r_4_1 ) );
  DFF_X1 key_c_r_reg_4_10 (.CK( clk ) , .D( key_c_r_3_10 ) , .Q( key_c_r_4_10 ) );
  DFF_X1 key_c_r_reg_4_11 (.CK( clk ) , .D( key_c_r_3_11 ) , .Q( key_c_r_4_11 ) );
  DFF_X1 key_c_r_reg_4_12 (.CK( clk ) , .D( key_c_r_3_12 ) , .Q( key_c_r_4_12 ) );
  DFF_X1 key_c_r_reg_4_13 (.CK( clk ) , .D( key_c_r_3_13 ) , .Q( key_c_r_4_13 ) );
  DFF_X1 key_c_r_reg_4_14 (.CK( clk ) , .D( key_c_r_3_14 ) , .Q( key_c_r_4_14 ) );
  DFF_X1 key_c_r_reg_4_15 (.CK( clk ) , .D( key_c_r_3_15 ) , .Q( key_c_r_4_15 ) );
  DFF_X1 key_c_r_reg_4_16 (.CK( clk ) , .D( key_c_r_3_16 ) , .Q( key_c_r_4_16 ) );
  DFF_X1 key_c_r_reg_4_17 (.CK( clk ) , .D( key_c_r_3_17 ) , .Q( key_c_r_4_17 ) );
  DFF_X1 key_c_r_reg_4_18 (.CK( clk ) , .D( key_c_r_3_18 ) , .Q( key_c_r_4_18 ) );
  DFF_X1 key_c_r_reg_4_19 (.CK( clk ) , .D( key_c_r_3_19 ) , .Q( key_c_r_4_19 ) );
  DFF_X1 key_c_r_reg_4_2 (.CK( clk ) , .D( key_c_r_3_2 ) , .Q( key_c_r_4_2 ) );
  DFF_X1 key_c_r_reg_4_20 (.CK( clk ) , .D( key_c_r_3_20 ) , .Q( key_c_r_4_20 ) );
  DFF_X1 key_c_r_reg_4_21 (.CK( clk ) , .D( key_c_r_3_21 ) , .Q( key_c_r_4_21 ) );
  DFF_X1 key_c_r_reg_4_22 (.CK( clk ) , .D( key_c_r_3_22 ) , .Q( key_c_r_4_22 ) );
  DFF_X1 key_c_r_reg_4_23 (.CK( clk ) , .D( key_c_r_3_23 ) , .Q( key_c_r_4_23 ) );
  DFF_X1 key_c_r_reg_4_24 (.CK( clk ) , .D( key_c_r_3_24 ) , .Q( key_c_r_4_24 ) );
  DFF_X1 key_c_r_reg_4_25 (.CK( clk ) , .D( key_c_r_3_25 ) , .Q( key_c_r_4_25 ) );
  DFF_X1 key_c_r_reg_4_26 (.CK( clk ) , .D( key_c_r_3_26 ) , .Q( key_c_r_4_26 ) );
  DFF_X1 key_c_r_reg_4_27 (.CK( clk ) , .D( key_c_r_3_27 ) , .Q( key_c_r_4_27 ) );
  DFF_X1 key_c_r_reg_4_28 (.CK( clk ) , .D( key_c_r_3_28 ) , .Q( key_c_r_4_28 ) );
  DFF_X1 key_c_r_reg_4_29 (.CK( clk ) , .D( key_c_r_3_29 ) , .Q( key_c_r_4_29 ) );
  DFF_X1 key_c_r_reg_4_3 (.CK( clk ) , .D( key_c_r_3_3 ) , .Q( key_c_r_4_3 ) );
  DFF_X1 key_c_r_reg_4_30 (.CK( clk ) , .D( key_c_r_3_30 ) , .Q( key_c_r_4_30 ) );
  DFF_X1 key_c_r_reg_4_31 (.CK( clk ) , .D( key_c_r_3_31 ) , .Q( key_c_r_4_31 ) );
  DFF_X1 key_c_r_reg_4_32 (.CK( clk ) , .D( key_c_r_3_32 ) , .Q( key_c_r_4_32 ) );
  DFF_X1 key_c_r_reg_4_33 (.CK( clk ) , .D( key_c_r_3_33 ) , .Q( key_c_r_4_33 ) );
  DFF_X1 key_c_r_reg_4_34 (.CK( clk ) , .D( key_c_r_3_34 ) , .Q( key_c_r_4_34 ) );
  DFF_X1 key_c_r_reg_4_35 (.CK( clk ) , .D( key_c_r_3_35 ) , .Q( key_c_r_4_35 ) );
  DFF_X1 key_c_r_reg_4_36 (.CK( clk ) , .D( key_c_r_3_36 ) , .Q( key_c_r_4_36 ) );
  DFF_X1 key_c_r_reg_4_37 (.CK( clk ) , .D( key_c_r_3_37 ) , .Q( key_c_r_4_37 ) );
  DFF_X1 key_c_r_reg_4_38 (.CK( clk ) , .D( key_c_r_3_38 ) , .Q( key_c_r_4_38 ) );
  DFF_X1 key_c_r_reg_4_39 (.CK( clk ) , .D( key_c_r_3_39 ) , .Q( key_c_r_4_39 ) );
  DFF_X1 key_c_r_reg_4_4 (.CK( clk ) , .D( key_c_r_3_4 ) , .Q( key_c_r_4_4 ) );
  DFF_X1 key_c_r_reg_4_40 (.CK( clk ) , .D( key_c_r_3_40 ) , .Q( key_c_r_4_40 ) );
  DFF_X1 key_c_r_reg_4_41 (.CK( clk ) , .D( key_c_r_3_41 ) , .Q( key_c_r_4_41 ) );
  DFF_X1 key_c_r_reg_4_42 (.CK( clk ) , .D( key_c_r_3_42 ) , .Q( key_c_r_4_42 ) );
  DFF_X1 key_c_r_reg_4_43 (.CK( clk ) , .D( key_c_r_3_43 ) , .Q( key_c_r_4_43 ) );
  DFF_X1 key_c_r_reg_4_44 (.CK( clk ) , .D( key_c_r_3_44 ) , .Q( key_c_r_4_44 ) );
  DFF_X1 key_c_r_reg_4_45 (.CK( clk ) , .D( key_c_r_3_45 ) , .Q( key_c_r_4_45 ) );
  DFF_X1 key_c_r_reg_4_46 (.CK( clk ) , .D( key_c_r_3_46 ) , .Q( key_c_r_4_46 ) );
  DFF_X1 key_c_r_reg_4_47 (.CK( clk ) , .D( key_c_r_3_47 ) , .Q( key_c_r_4_47 ) );
  DFF_X1 key_c_r_reg_4_48 (.CK( clk ) , .D( key_c_r_3_48 ) , .Q( key_c_r_4_48 ) );
  DFF_X1 key_c_r_reg_4_49 (.CK( clk ) , .D( key_c_r_3_49 ) , .Q( key_c_r_4_49 ) );
  DFF_X1 key_c_r_reg_4_5 (.CK( clk ) , .D( key_c_r_3_5 ) , .Q( key_c_r_4_5 ) );
  DFF_X1 key_c_r_reg_4_50 (.CK( clk ) , .D( key_c_r_3_50 ) , .Q( key_c_r_4_50 ) );
  DFF_X1 key_c_r_reg_4_51 (.CK( clk ) , .D( key_c_r_3_51 ) , .Q( key_c_r_4_51 ) );
  DFF_X1 key_c_r_reg_4_52 (.CK( clk ) , .D( key_c_r_3_52 ) , .Q( key_c_r_4_52 ) );
  DFF_X1 key_c_r_reg_4_53 (.CK( clk ) , .D( key_c_r_3_53 ) , .Q( key_c_r_4_53 ) );
  DFF_X1 key_c_r_reg_4_54 (.CK( clk ) , .D( key_c_r_3_54 ) , .Q( key_c_r_4_54 ) );
  DFF_X1 key_c_r_reg_4_55 (.CK( clk ) , .D( key_c_r_3_55 ) , .Q( key_c_r_4_55 ) );
  DFF_X1 key_c_r_reg_4_6 (.CK( clk ) , .D( key_c_r_3_6 ) , .Q( key_c_r_4_6 ) );
  DFF_X1 key_c_r_reg_4_7 (.CK( clk ) , .D( key_c_r_3_7 ) , .Q( key_c_r_4_7 ) );
  DFF_X1 key_c_r_reg_4_8 (.CK( clk ) , .D( key_c_r_3_8 ) , .Q( key_c_r_4_8 ) );
  DFF_X1 key_c_r_reg_4_9 (.CK( clk ) , .D( key_c_r_3_9 ) , .Q( key_c_r_4_9 ) );
  DFF_X1 key_c_r_reg_5_0 (.CK( clk ) , .D( key_c_r_4_0 ) , .Q( key_c_r_5_0 ) );
  DFF_X1 key_c_r_reg_5_1 (.CK( clk ) , .D( key_c_r_4_1 ) , .Q( key_c_r_5_1 ) );
  DFF_X1 key_c_r_reg_5_10 (.CK( clk ) , .D( key_c_r_4_10 ) , .Q( key_c_r_5_10 ) );
  DFF_X1 key_c_r_reg_5_11 (.CK( clk ) , .D( key_c_r_4_11 ) , .Q( key_c_r_5_11 ) );
  DFF_X1 key_c_r_reg_5_12 (.CK( clk ) , .D( key_c_r_4_12 ) , .Q( key_c_r_5_12 ) );
  DFF_X1 key_c_r_reg_5_13 (.CK( clk ) , .D( key_c_r_4_13 ) , .Q( key_c_r_5_13 ) );
  DFF_X1 key_c_r_reg_5_14 (.CK( clk ) , .D( key_c_r_4_14 ) , .Q( key_c_r_5_14 ) );
  DFF_X1 key_c_r_reg_5_15 (.CK( clk ) , .D( key_c_r_4_15 ) , .Q( key_c_r_5_15 ) );
  DFF_X1 key_c_r_reg_5_16 (.CK( clk ) , .D( key_c_r_4_16 ) , .Q( key_c_r_5_16 ) );
  DFF_X1 key_c_r_reg_5_17 (.CK( clk ) , .D( key_c_r_4_17 ) , .Q( key_c_r_5_17 ) );
  DFF_X1 key_c_r_reg_5_18 (.CK( clk ) , .D( key_c_r_4_18 ) , .Q( key_c_r_5_18 ) );
  DFF_X1 key_c_r_reg_5_19 (.CK( clk ) , .D( key_c_r_4_19 ) , .Q( key_c_r_5_19 ) );
  DFF_X1 key_c_r_reg_5_2 (.CK( clk ) , .D( key_c_r_4_2 ) , .Q( key_c_r_5_2 ) );
  DFF_X1 key_c_r_reg_5_20 (.CK( clk ) , .D( key_c_r_4_20 ) , .Q( key_c_r_5_20 ) );
  DFF_X1 key_c_r_reg_5_21 (.CK( clk ) , .D( key_c_r_4_21 ) , .Q( key_c_r_5_21 ) );
  DFF_X1 key_c_r_reg_5_22 (.CK( clk ) , .D( key_c_r_4_22 ) , .Q( key_c_r_5_22 ) );
  DFF_X1 key_c_r_reg_5_23 (.CK( clk ) , .D( key_c_r_4_23 ) , .Q( key_c_r_5_23 ) );
  DFF_X1 key_c_r_reg_5_24 (.CK( clk ) , .D( key_c_r_4_24 ) , .Q( key_c_r_5_24 ) );
  DFF_X1 key_c_r_reg_5_25 (.CK( clk ) , .D( key_c_r_4_25 ) , .Q( key_c_r_5_25 ) );
  DFF_X1 key_c_r_reg_5_26 (.CK( clk ) , .D( key_c_r_4_26 ) , .Q( key_c_r_5_26 ) );
  DFF_X1 key_c_r_reg_5_27 (.CK( clk ) , .D( key_c_r_4_27 ) , .Q( key_c_r_5_27 ) );
  DFF_X1 key_c_r_reg_5_28 (.CK( clk ) , .D( key_c_r_4_28 ) , .Q( key_c_r_5_28 ) );
  DFF_X1 key_c_r_reg_5_29 (.CK( clk ) , .D( key_c_r_4_29 ) , .Q( key_c_r_5_29 ) );
  DFF_X1 key_c_r_reg_5_3 (.CK( clk ) , .D( key_c_r_4_3 ) , .Q( key_c_r_5_3 ) );
  DFF_X1 key_c_r_reg_5_30 (.CK( clk ) , .D( key_c_r_4_30 ) , .Q( key_c_r_5_30 ) );
  DFF_X1 key_c_r_reg_5_31 (.CK( clk ) , .D( key_c_r_4_31 ) , .Q( key_c_r_5_31 ) );
  DFF_X1 key_c_r_reg_5_32 (.CK( clk ) , .D( key_c_r_4_32 ) , .Q( key_c_r_5_32 ) );
  DFF_X1 key_c_r_reg_5_33 (.CK( clk ) , .D( key_c_r_4_33 ) , .Q( key_c_r_5_33 ) );
  DFF_X1 key_c_r_reg_5_34 (.CK( clk ) , .D( key_c_r_4_34 ) , .Q( key_c_r_5_34 ) );
  DFF_X1 key_c_r_reg_5_35 (.CK( clk ) , .D( key_c_r_4_35 ) , .Q( key_c_r_5_35 ) );
  DFF_X1 key_c_r_reg_5_36 (.CK( clk ) , .D( key_c_r_4_36 ) , .Q( key_c_r_5_36 ) );
  DFF_X1 key_c_r_reg_5_37 (.CK( clk ) , .D( key_c_r_4_37 ) , .Q( key_c_r_5_37 ) );
  DFF_X1 key_c_r_reg_5_38 (.CK( clk ) , .D( key_c_r_4_38 ) , .Q( key_c_r_5_38 ) );
  DFF_X1 key_c_r_reg_5_39 (.CK( clk ) , .D( key_c_r_4_39 ) , .Q( key_c_r_5_39 ) );
  DFF_X1 key_c_r_reg_5_4 (.CK( clk ) , .D( key_c_r_4_4 ) , .Q( key_c_r_5_4 ) );
  DFF_X1 key_c_r_reg_5_40 (.CK( clk ) , .D( key_c_r_4_40 ) , .Q( key_c_r_5_40 ) );
  DFF_X1 key_c_r_reg_5_41 (.CK( clk ) , .D( key_c_r_4_41 ) , .Q( key_c_r_5_41 ) );
  DFF_X1 key_c_r_reg_5_42 (.CK( clk ) , .D( key_c_r_4_42 ) , .Q( key_c_r_5_42 ) );
  DFF_X1 key_c_r_reg_5_43 (.CK( clk ) , .D( key_c_r_4_43 ) , .Q( key_c_r_5_43 ) );
  DFF_X1 key_c_r_reg_5_44 (.CK( clk ) , .D( key_c_r_4_44 ) , .Q( key_c_r_5_44 ) );
  DFF_X1 key_c_r_reg_5_45 (.CK( clk ) , .D( key_c_r_4_45 ) , .Q( key_c_r_5_45 ) );
  DFF_X1 key_c_r_reg_5_46 (.CK( clk ) , .D( key_c_r_4_46 ) , .Q( key_c_r_5_46 ) );
  DFF_X1 key_c_r_reg_5_47 (.CK( clk ) , .D( key_c_r_4_47 ) , .Q( key_c_r_5_47 ) );
  DFF_X1 key_c_r_reg_5_48 (.CK( clk ) , .D( key_c_r_4_48 ) , .Q( key_c_r_5_48 ) );
  DFF_X1 key_c_r_reg_5_49 (.CK( clk ) , .D( key_c_r_4_49 ) , .Q( key_c_r_5_49 ) );
  DFF_X1 key_c_r_reg_5_5 (.CK( clk ) , .D( key_c_r_4_5 ) , .Q( key_c_r_5_5 ) );
  DFF_X1 key_c_r_reg_5_50 (.CK( clk ) , .D( key_c_r_4_50 ) , .Q( key_c_r_5_50 ) );
  DFF_X1 key_c_r_reg_5_51 (.CK( clk ) , .D( key_c_r_4_51 ) , .Q( key_c_r_5_51 ) );
  DFF_X1 key_c_r_reg_5_52 (.CK( clk ) , .D( key_c_r_4_52 ) , .Q( key_c_r_5_52 ) );
  DFF_X1 key_c_r_reg_5_53 (.CK( clk ) , .D( key_c_r_4_53 ) , .Q( key_c_r_5_53 ) );
  DFF_X1 key_c_r_reg_5_54 (.CK( clk ) , .D( key_c_r_4_54 ) , .Q( key_c_r_5_54 ) );
  DFF_X1 key_c_r_reg_5_55 (.CK( clk ) , .D( key_c_r_4_55 ) , .Q( key_c_r_5_55 ) );
  DFF_X1 key_c_r_reg_5_6 (.CK( clk ) , .D( key_c_r_4_6 ) , .Q( key_c_r_5_6 ) );
  DFF_X1 key_c_r_reg_5_7 (.CK( clk ) , .D( key_c_r_4_7 ) , .Q( key_c_r_5_7 ) );
  DFF_X1 key_c_r_reg_5_8 (.CK( clk ) , .D( key_c_r_4_8 ) , .Q( key_c_r_5_8 ) );
  DFF_X1 key_c_r_reg_5_9 (.CK( clk ) , .D( key_c_r_4_9 ) , .Q( key_c_r_5_9 ) );
  DFF_X1 key_c_r_reg_6_0 (.CK( clk ) , .D( key_c_r_5_0 ) , .Q( key_c_r_6_0 ) );
  DFF_X1 key_c_r_reg_6_1 (.CK( clk ) , .D( key_c_r_5_1 ) , .Q( key_c_r_6_1 ) );
  DFF_X1 key_c_r_reg_6_10 (.CK( clk ) , .D( key_c_r_5_10 ) , .Q( key_c_r_6_10 ) );
  DFF_X1 key_c_r_reg_6_11 (.CK( clk ) , .D( key_c_r_5_11 ) , .Q( key_c_r_6_11 ) );
  DFF_X1 key_c_r_reg_6_12 (.CK( clk ) , .D( key_c_r_5_12 ) , .Q( key_c_r_6_12 ) );
  DFF_X1 key_c_r_reg_6_13 (.CK( clk ) , .D( key_c_r_5_13 ) , .Q( key_c_r_6_13 ) );
  DFF_X1 key_c_r_reg_6_14 (.CK( clk ) , .D( key_c_r_5_14 ) , .Q( key_c_r_6_14 ) );
  DFF_X1 key_c_r_reg_6_15 (.CK( clk ) , .D( key_c_r_5_15 ) , .Q( key_c_r_6_15 ) );
  DFF_X1 key_c_r_reg_6_16 (.CK( clk ) , .D( key_c_r_5_16 ) , .Q( key_c_r_6_16 ) );
  DFF_X1 key_c_r_reg_6_17 (.CK( clk ) , .D( key_c_r_5_17 ) , .Q( key_c_r_6_17 ) );
  DFF_X1 key_c_r_reg_6_18 (.CK( clk ) , .D( key_c_r_5_18 ) , .Q( key_c_r_6_18 ) );
  DFF_X1 key_c_r_reg_6_19 (.CK( clk ) , .D( key_c_r_5_19 ) , .Q( key_c_r_6_19 ) );
  DFF_X1 key_c_r_reg_6_2 (.CK( clk ) , .D( key_c_r_5_2 ) , .Q( key_c_r_6_2 ) );
  DFF_X1 key_c_r_reg_6_20 (.CK( clk ) , .D( key_c_r_5_20 ) , .Q( key_c_r_6_20 ) );
  DFF_X1 key_c_r_reg_6_21 (.CK( clk ) , .D( key_c_r_5_21 ) , .Q( key_c_r_6_21 ) );
  DFF_X1 key_c_r_reg_6_22 (.CK( clk ) , .D( key_c_r_5_22 ) , .Q( key_c_r_6_22 ) );
  DFF_X1 key_c_r_reg_6_23 (.CK( clk ) , .D( key_c_r_5_23 ) , .Q( key_c_r_6_23 ) );
  DFF_X1 key_c_r_reg_6_24 (.CK( clk ) , .D( key_c_r_5_24 ) , .Q( key_c_r_6_24 ) );
  DFF_X1 key_c_r_reg_6_25 (.CK( clk ) , .D( key_c_r_5_25 ) , .Q( key_c_r_6_25 ) );
  DFF_X1 key_c_r_reg_6_26 (.CK( clk ) , .D( key_c_r_5_26 ) , .Q( key_c_r_6_26 ) );
  DFF_X1 key_c_r_reg_6_27 (.CK( clk ) , .D( key_c_r_5_27 ) , .Q( key_c_r_6_27 ) );
  DFF_X1 key_c_r_reg_6_28 (.CK( clk ) , .D( key_c_r_5_28 ) , .Q( key_c_r_6_28 ) );
  DFF_X1 key_c_r_reg_6_29 (.CK( clk ) , .D( key_c_r_5_29 ) , .Q( key_c_r_6_29 ) );
  DFF_X1 key_c_r_reg_6_3 (.CK( clk ) , .D( key_c_r_5_3 ) , .Q( key_c_r_6_3 ) );
  DFF_X1 key_c_r_reg_6_30 (.CK( clk ) , .D( key_c_r_5_30 ) , .Q( key_c_r_6_30 ) );
  DFF_X1 key_c_r_reg_6_31 (.CK( clk ) , .D( key_c_r_5_31 ) , .Q( key_c_r_6_31 ) );
  DFF_X1 key_c_r_reg_6_32 (.CK( clk ) , .D( key_c_r_5_32 ) , .Q( key_c_r_6_32 ) );
  DFF_X1 key_c_r_reg_6_33 (.CK( clk ) , .D( key_c_r_5_33 ) , .Q( key_c_r_6_33 ) );
  DFF_X1 key_c_r_reg_6_34 (.CK( clk ) , .D( key_c_r_5_34 ) , .Q( key_c_r_6_34 ) );
  DFF_X1 key_c_r_reg_6_35 (.CK( clk ) , .D( key_c_r_5_35 ) , .Q( key_c_r_6_35 ) );
  DFF_X1 key_c_r_reg_6_36 (.CK( clk ) , .D( key_c_r_5_36 ) , .Q( key_c_r_6_36 ) );
  DFF_X1 key_c_r_reg_6_37 (.CK( clk ) , .D( key_c_r_5_37 ) , .Q( key_c_r_6_37 ) );
  DFF_X1 key_c_r_reg_6_38 (.CK( clk ) , .D( key_c_r_5_38 ) , .Q( key_c_r_6_38 ) );
  DFF_X1 key_c_r_reg_6_39 (.CK( clk ) , .D( key_c_r_5_39 ) , .Q( key_c_r_6_39 ) );
  DFF_X1 key_c_r_reg_6_4 (.CK( clk ) , .D( key_c_r_5_4 ) , .Q( key_c_r_6_4 ) );
  DFF_X1 key_c_r_reg_6_40 (.CK( clk ) , .D( key_c_r_5_40 ) , .Q( key_c_r_6_40 ) );
  DFF_X1 key_c_r_reg_6_41 (.CK( clk ) , .D( key_c_r_5_41 ) , .Q( key_c_r_6_41 ) );
  DFF_X1 key_c_r_reg_6_42 (.CK( clk ) , .D( key_c_r_5_42 ) , .Q( key_c_r_6_42 ) );
  DFF_X1 key_c_r_reg_6_43 (.CK( clk ) , .D( key_c_r_5_43 ) , .Q( key_c_r_6_43 ) );
  DFF_X1 key_c_r_reg_6_44 (.CK( clk ) , .D( key_c_r_5_44 ) , .Q( key_c_r_6_44 ) );
  DFF_X1 key_c_r_reg_6_45 (.CK( clk ) , .D( key_c_r_5_45 ) , .Q( key_c_r_6_45 ) );
  DFF_X1 key_c_r_reg_6_46 (.CK( clk ) , .D( key_c_r_5_46 ) , .Q( key_c_r_6_46 ) );
  DFF_X1 key_c_r_reg_6_47 (.CK( clk ) , .D( key_c_r_5_47 ) , .Q( key_c_r_6_47 ) );
  DFF_X1 key_c_r_reg_6_48 (.CK( clk ) , .D( key_c_r_5_48 ) , .Q( key_c_r_6_48 ) );
  DFF_X1 key_c_r_reg_6_49 (.CK( clk ) , .D( key_c_r_5_49 ) , .Q( key_c_r_6_49 ) );
  DFF_X1 key_c_r_reg_6_5 (.CK( clk ) , .D( key_c_r_5_5 ) , .Q( key_c_r_6_5 ) );
  DFF_X1 key_c_r_reg_6_50 (.CK( clk ) , .D( key_c_r_5_50 ) , .Q( key_c_r_6_50 ) );
  DFF_X1 key_c_r_reg_6_51 (.CK( clk ) , .D( key_c_r_5_51 ) , .Q( key_c_r_6_51 ) );
  DFF_X1 key_c_r_reg_6_52 (.CK( clk ) , .D( key_c_r_5_52 ) , .Q( key_c_r_6_52 ) );
  DFF_X1 key_c_r_reg_6_53 (.CK( clk ) , .D( key_c_r_5_53 ) , .Q( key_c_r_6_53 ) );
  DFF_X1 key_c_r_reg_6_54 (.CK( clk ) , .D( key_c_r_5_54 ) , .Q( key_c_r_6_54 ) );
  DFF_X1 key_c_r_reg_6_55 (.CK( clk ) , .D( key_c_r_5_55 ) , .Q( key_c_r_6_55 ) );
  DFF_X1 key_c_r_reg_6_6 (.CK( clk ) , .D( key_c_r_5_6 ) , .Q( key_c_r_6_6 ) );
  DFF_X1 key_c_r_reg_6_7 (.CK( clk ) , .D( key_c_r_5_7 ) , .Q( key_c_r_6_7 ) );
  DFF_X1 key_c_r_reg_6_8 (.CK( clk ) , .D( key_c_r_5_8 ) , .Q( key_c_r_6_8 ) );
  DFF_X1 key_c_r_reg_6_9 (.CK( clk ) , .D( key_c_r_5_9 ) , .Q( key_c_r_6_9 ) );
  DFF_X1 key_c_r_reg_7_0 (.CK( clk ) , .D( key_c_r_6_0 ) , .Q( key_c_r_7_0 ) );
  DFF_X1 key_c_r_reg_7_1 (.CK( clk ) , .D( key_c_r_6_1 ) , .Q( key_c_r_7_1 ) );
  DFF_X1 key_c_r_reg_7_10 (.CK( clk ) , .D( key_c_r_6_10 ) , .Q( key_c_r_7_10 ) );
  DFF_X1 key_c_r_reg_7_11 (.CK( clk ) , .D( key_c_r_6_11 ) , .Q( key_c_r_7_11 ) );
  DFF_X1 key_c_r_reg_7_12 (.CK( clk ) , .D( key_c_r_6_12 ) , .Q( key_c_r_7_12 ) );
  DFF_X1 key_c_r_reg_7_13 (.CK( clk ) , .D( key_c_r_6_13 ) , .Q( key_c_r_7_13 ) );
  DFF_X1 key_c_r_reg_7_14 (.CK( clk ) , .D( key_c_r_6_14 ) , .Q( key_c_r_7_14 ) );
  DFF_X1 key_c_r_reg_7_15 (.CK( clk ) , .D( key_c_r_6_15 ) , .Q( key_c_r_7_15 ) );
  DFF_X1 key_c_r_reg_7_16 (.CK( clk ) , .D( key_c_r_6_16 ) , .Q( key_c_r_7_16 ) );
  DFF_X1 key_c_r_reg_7_17 (.CK( clk ) , .D( key_c_r_6_17 ) , .Q( key_c_r_7_17 ) );
  DFF_X1 key_c_r_reg_7_18 (.CK( clk ) , .D( key_c_r_6_18 ) , .Q( key_c_r_7_18 ) );
  DFF_X1 key_c_r_reg_7_19 (.CK( clk ) , .D( key_c_r_6_19 ) , .Q( key_c_r_7_19 ) );
  DFF_X1 key_c_r_reg_7_2 (.CK( clk ) , .D( key_c_r_6_2 ) , .Q( key_c_r_7_2 ) );
  DFF_X1 key_c_r_reg_7_20 (.CK( clk ) , .D( key_c_r_6_20 ) , .Q( key_c_r_7_20 ) );
  DFF_X1 key_c_r_reg_7_21 (.CK( clk ) , .D( key_c_r_6_21 ) , .Q( key_c_r_7_21 ) );
  DFF_X1 key_c_r_reg_7_22 (.CK( clk ) , .D( key_c_r_6_22 ) , .Q( key_c_r_7_22 ) );
  DFF_X1 key_c_r_reg_7_23 (.CK( clk ) , .D( key_c_r_6_23 ) , .Q( key_c_r_7_23 ) );
  DFF_X1 key_c_r_reg_7_24 (.CK( clk ) , .D( key_c_r_6_24 ) , .Q( key_c_r_7_24 ) );
  DFF_X1 key_c_r_reg_7_25 (.CK( clk ) , .D( key_c_r_6_25 ) , .Q( key_c_r_7_25 ) );
  DFF_X1 key_c_r_reg_7_26 (.CK( clk ) , .D( key_c_r_6_26 ) , .Q( key_c_r_7_26 ) );
  DFF_X1 key_c_r_reg_7_27 (.CK( clk ) , .D( key_c_r_6_27 ) , .Q( key_c_r_7_27 ) );
  DFF_X1 key_c_r_reg_7_28 (.CK( clk ) , .D( key_c_r_6_28 ) , .Q( key_c_r_7_28 ) );
  DFF_X1 key_c_r_reg_7_29 (.CK( clk ) , .D( key_c_r_6_29 ) , .Q( key_c_r_7_29 ) );
  DFF_X1 key_c_r_reg_7_3 (.CK( clk ) , .D( key_c_r_6_3 ) , .Q( key_c_r_7_3 ) );
  DFF_X1 key_c_r_reg_7_30 (.CK( clk ) , .D( key_c_r_6_30 ) , .Q( key_c_r_7_30 ) );
  DFF_X1 key_c_r_reg_7_31 (.CK( clk ) , .D( key_c_r_6_31 ) , .Q( key_c_r_7_31 ) );
  DFF_X1 key_c_r_reg_7_32 (.CK( clk ) , .D( key_c_r_6_32 ) , .Q( key_c_r_7_32 ) );
  DFF_X1 key_c_r_reg_7_33 (.CK( clk ) , .D( key_c_r_6_33 ) , .Q( key_c_r_7_33 ) );
  DFF_X1 key_c_r_reg_7_34 (.CK( clk ) , .D( key_c_r_6_34 ) , .Q( key_c_r_7_34 ) );
  DFF_X1 key_c_r_reg_7_35 (.CK( clk ) , .D( key_c_r_6_35 ) , .Q( key_c_r_7_35 ) );
  DFF_X1 key_c_r_reg_7_36 (.CK( clk ) , .D( key_c_r_6_36 ) , .Q( key_c_r_7_36 ) );
  DFF_X1 key_c_r_reg_7_37 (.CK( clk ) , .D( key_c_r_6_37 ) , .Q( key_c_r_7_37 ) );
  DFF_X1 key_c_r_reg_7_38 (.CK( clk ) , .D( key_c_r_6_38 ) , .Q( key_c_r_7_38 ) );
  DFF_X1 key_c_r_reg_7_39 (.CK( clk ) , .D( key_c_r_6_39 ) , .Q( key_c_r_7_39 ) );
  DFF_X1 key_c_r_reg_7_4 (.CK( clk ) , .D( key_c_r_6_4 ) , .Q( key_c_r_7_4 ) );
  DFF_X1 key_c_r_reg_7_40 (.CK( clk ) , .D( key_c_r_6_40 ) , .Q( key_c_r_7_40 ) );
  DFF_X1 key_c_r_reg_7_41 (.CK( clk ) , .D( key_c_r_6_41 ) , .Q( key_c_r_7_41 ) );
  DFF_X1 key_c_r_reg_7_42 (.CK( clk ) , .D( key_c_r_6_42 ) , .Q( key_c_r_7_42 ) );
  DFF_X1 key_c_r_reg_7_43 (.CK( clk ) , .D( key_c_r_6_43 ) , .Q( key_c_r_7_43 ) );
  DFF_X1 key_c_r_reg_7_44 (.CK( clk ) , .D( key_c_r_6_44 ) , .Q( key_c_r_7_44 ) );
  DFF_X1 key_c_r_reg_7_45 (.CK( clk ) , .D( key_c_r_6_45 ) , .Q( key_c_r_7_45 ) );
  DFF_X1 key_c_r_reg_7_46 (.CK( clk ) , .D( key_c_r_6_46 ) , .Q( key_c_r_7_46 ) );
  DFF_X1 key_c_r_reg_7_47 (.CK( clk ) , .D( key_c_r_6_47 ) , .Q( key_c_r_7_47 ) );
  DFF_X1 key_c_r_reg_7_48 (.CK( clk ) , .D( key_c_r_6_48 ) , .Q( key_c_r_7_48 ) );
  DFF_X1 key_c_r_reg_7_49 (.CK( clk ) , .D( key_c_r_6_49 ) , .Q( key_c_r_7_49 ) );
  DFF_X1 key_c_r_reg_7_5 (.CK( clk ) , .D( key_c_r_6_5 ) , .Q( key_c_r_7_5 ) );
  DFF_X1 key_c_r_reg_7_50 (.CK( clk ) , .D( key_c_r_6_50 ) , .Q( key_c_r_7_50 ) );
  DFF_X1 key_c_r_reg_7_51 (.CK( clk ) , .D( key_c_r_6_51 ) , .Q( key_c_r_7_51 ) );
  DFF_X1 key_c_r_reg_7_52 (.CK( clk ) , .D( key_c_r_6_52 ) , .Q( key_c_r_7_52 ) );
  DFF_X1 key_c_r_reg_7_53 (.CK( clk ) , .D( key_c_r_6_53 ) , .Q( key_c_r_7_53 ) );
  DFF_X1 key_c_r_reg_7_54 (.CK( clk ) , .D( key_c_r_6_54 ) , .Q( key_c_r_7_54 ) );
  DFF_X1 key_c_r_reg_7_55 (.CK( clk ) , .D( key_c_r_6_55 ) , .Q( key_c_r_7_55 ) );
  DFF_X1 key_c_r_reg_7_6 (.CK( clk ) , .D( key_c_r_6_6 ) , .Q( key_c_r_7_6 ) );
  DFF_X1 key_c_r_reg_7_7 (.CK( clk ) , .D( key_c_r_6_7 ) , .Q( key_c_r_7_7 ) );
  DFF_X1 key_c_r_reg_7_8 (.CK( clk ) , .D( key_c_r_6_8 ) , .Q( key_c_r_7_8 ) );
  DFF_X1 key_c_r_reg_7_9 (.CK( clk ) , .D( key_c_r_6_9 ) , .Q( key_c_r_7_9 ) );
  DFF_X1 key_c_r_reg_8_0 (.CK( clk ) , .D( key_c_r_7_0 ) , .Q( key_c_r_8_0 ) );
  DFF_X1 key_c_r_reg_8_1 (.CK( clk ) , .D( key_c_r_7_1 ) , .Q( key_c_r_8_1 ) );
  DFF_X1 key_c_r_reg_8_10 (.CK( clk ) , .D( key_c_r_7_10 ) , .Q( key_c_r_8_10 ) );
  DFF_X1 key_c_r_reg_8_11 (.CK( clk ) , .D( key_c_r_7_11 ) , .Q( key_c_r_8_11 ) );
  DFF_X1 key_c_r_reg_8_12 (.CK( clk ) , .D( key_c_r_7_12 ) , .Q( key_c_r_8_12 ) );
  DFF_X1 key_c_r_reg_8_13 (.CK( clk ) , .D( key_c_r_7_13 ) , .Q( key_c_r_8_13 ) );
  DFF_X1 key_c_r_reg_8_14 (.CK( clk ) , .D( key_c_r_7_14 ) , .Q( key_c_r_8_14 ) );
  DFF_X1 key_c_r_reg_8_15 (.CK( clk ) , .D( key_c_r_7_15 ) , .Q( key_c_r_8_15 ) );
  DFF_X1 key_c_r_reg_8_16 (.CK( clk ) , .D( key_c_r_7_16 ) , .Q( key_c_r_8_16 ) );
  DFF_X1 key_c_r_reg_8_17 (.CK( clk ) , .D( key_c_r_7_17 ) , .Q( key_c_r_8_17 ) );
  DFF_X1 key_c_r_reg_8_18 (.CK( clk ) , .D( key_c_r_7_18 ) , .Q( key_c_r_8_18 ) );
  DFF_X1 key_c_r_reg_8_19 (.CK( clk ) , .D( key_c_r_7_19 ) , .Q( key_c_r_8_19 ) );
  DFF_X1 key_c_r_reg_8_2 (.CK( clk ) , .D( key_c_r_7_2 ) , .Q( key_c_r_8_2 ) );
  DFF_X1 key_c_r_reg_8_20 (.CK( clk ) , .D( key_c_r_7_20 ) , .Q( key_c_r_8_20 ) );
  DFF_X1 key_c_r_reg_8_21 (.CK( clk ) , .D( key_c_r_7_21 ) , .Q( key_c_r_8_21 ) );
  DFF_X1 key_c_r_reg_8_22 (.CK( clk ) , .D( key_c_r_7_22 ) , .Q( key_c_r_8_22 ) );
  DFF_X1 key_c_r_reg_8_23 (.CK( clk ) , .D( key_c_r_7_23 ) , .Q( key_c_r_8_23 ) );
  DFF_X1 key_c_r_reg_8_24 (.CK( clk ) , .D( key_c_r_7_24 ) , .Q( key_c_r_8_24 ) );
  DFF_X1 key_c_r_reg_8_25 (.CK( clk ) , .D( key_c_r_7_25 ) , .Q( key_c_r_8_25 ) );
  DFF_X1 key_c_r_reg_8_26 (.CK( clk ) , .D( key_c_r_7_26 ) , .Q( key_c_r_8_26 ) );
  DFF_X1 key_c_r_reg_8_27 (.CK( clk ) , .D( key_c_r_7_27 ) , .Q( key_c_r_8_27 ) );
  DFF_X1 key_c_r_reg_8_28 (.CK( clk ) , .D( key_c_r_7_28 ) , .Q( key_c_r_8_28 ) );
  DFF_X1 key_c_r_reg_8_29 (.CK( clk ) , .D( key_c_r_7_29 ) , .Q( key_c_r_8_29 ) );
  DFF_X1 key_c_r_reg_8_3 (.CK( clk ) , .D( key_c_r_7_3 ) , .Q( key_c_r_8_3 ) );
  DFF_X1 key_c_r_reg_8_30 (.CK( clk ) , .D( key_c_r_7_30 ) , .Q( key_c_r_8_30 ) );
  DFF_X1 key_c_r_reg_8_31 (.CK( clk ) , .D( key_c_r_7_31 ) , .Q( key_c_r_8_31 ) );
  DFF_X1 key_c_r_reg_8_32 (.CK( clk ) , .D( key_c_r_7_32 ) , .Q( key_c_r_8_32 ) );
  DFF_X1 key_c_r_reg_8_33 (.CK( clk ) , .D( key_c_r_7_33 ) , .Q( key_c_r_8_33 ) );
  DFF_X1 key_c_r_reg_8_34 (.CK( clk ) , .D( key_c_r_7_34 ) , .Q( key_c_r_8_34 ) );
  DFF_X1 key_c_r_reg_8_35 (.CK( clk ) , .D( key_c_r_7_35 ) , .Q( key_c_r_8_35 ) );
  DFF_X1 key_c_r_reg_8_36 (.CK( clk ) , .D( key_c_r_7_36 ) , .Q( key_c_r_8_36 ) );
  DFF_X1 key_c_r_reg_8_37 (.CK( clk ) , .D( key_c_r_7_37 ) , .Q( key_c_r_8_37 ) );
  DFF_X1 key_c_r_reg_8_38 (.CK( clk ) , .D( key_c_r_7_38 ) , .Q( key_c_r_8_38 ) );
  DFF_X1 key_c_r_reg_8_39 (.CK( clk ) , .D( key_c_r_7_39 ) , .Q( key_c_r_8_39 ) );
  DFF_X1 key_c_r_reg_8_4 (.CK( clk ) , .D( key_c_r_7_4 ) , .Q( key_c_r_8_4 ) );
  DFF_X1 key_c_r_reg_8_40 (.CK( clk ) , .D( key_c_r_7_40 ) , .Q( key_c_r_8_40 ) );
  DFF_X1 key_c_r_reg_8_41 (.CK( clk ) , .D( key_c_r_7_41 ) , .Q( key_c_r_8_41 ) );
  DFF_X1 key_c_r_reg_8_42 (.CK( clk ) , .D( key_c_r_7_42 ) , .Q( key_c_r_8_42 ) );
  DFF_X1 key_c_r_reg_8_43 (.CK( clk ) , .D( key_c_r_7_43 ) , .Q( key_c_r_8_43 ) );
  DFF_X1 key_c_r_reg_8_44 (.CK( clk ) , .D( key_c_r_7_44 ) , .Q( key_c_r_8_44 ) );
  DFF_X1 key_c_r_reg_8_45 (.CK( clk ) , .D( key_c_r_7_45 ) , .Q( key_c_r_8_45 ) );
  DFF_X1 key_c_r_reg_8_46 (.CK( clk ) , .D( key_c_r_7_46 ) , .Q( key_c_r_8_46 ) );
  DFF_X1 key_c_r_reg_8_47 (.CK( clk ) , .D( key_c_r_7_47 ) , .Q( key_c_r_8_47 ) );
  DFF_X1 key_c_r_reg_8_48 (.CK( clk ) , .D( key_c_r_7_48 ) , .Q( key_c_r_8_48 ) );
  DFF_X1 key_c_r_reg_8_49 (.CK( clk ) , .D( key_c_r_7_49 ) , .Q( key_c_r_8_49 ) );
  DFF_X1 key_c_r_reg_8_5 (.CK( clk ) , .D( key_c_r_7_5 ) , .Q( key_c_r_8_5 ) );
  DFF_X1 key_c_r_reg_8_50 (.CK( clk ) , .D( key_c_r_7_50 ) , .Q( key_c_r_8_50 ) );
  DFF_X1 key_c_r_reg_8_51 (.CK( clk ) , .D( key_c_r_7_51 ) , .Q( key_c_r_8_51 ) );
  DFF_X1 key_c_r_reg_8_52 (.CK( clk ) , .D( key_c_r_7_52 ) , .Q( key_c_r_8_52 ) );
  DFF_X1 key_c_r_reg_8_53 (.CK( clk ) , .D( key_c_r_7_53 ) , .Q( key_c_r_8_53 ) );
  DFF_X1 key_c_r_reg_8_54 (.CK( clk ) , .D( key_c_r_7_54 ) , .Q( key_c_r_8_54 ) );
  DFF_X1 key_c_r_reg_8_55 (.CK( clk ) , .D( key_c_r_7_55 ) , .Q( key_c_r_8_55 ) );
  DFF_X1 key_c_r_reg_8_6 (.CK( clk ) , .D( key_c_r_7_6 ) , .Q( key_c_r_8_6 ) );
  DFF_X1 key_c_r_reg_8_7 (.CK( clk ) , .D( key_c_r_7_7 ) , .Q( key_c_r_8_7 ) );
  DFF_X1 key_c_r_reg_8_8 (.CK( clk ) , .D( key_c_r_7_8 ) , .Q( key_c_r_8_8 ) );
  DFF_X1 key_c_r_reg_8_9 (.CK( clk ) , .D( key_c_r_7_9 ) , .Q( key_c_r_8_9 ) );
  DFF_X1 key_c_r_reg_9_0 (.CK( clk ) , .D( key_c_r_8_0 ) , .Q( key_c_r_9_0 ) );
  DFF_X1 key_c_r_reg_9_1 (.CK( clk ) , .D( key_c_r_8_1 ) , .Q( key_c_r_9_1 ) );
  DFF_X1 key_c_r_reg_9_10 (.CK( clk ) , .D( key_c_r_8_10 ) , .Q( key_c_r_9_10 ) );
  DFF_X1 key_c_r_reg_9_11 (.CK( clk ) , .D( key_c_r_8_11 ) , .Q( key_c_r_9_11 ) );
  DFF_X1 key_c_r_reg_9_12 (.CK( clk ) , .D( key_c_r_8_12 ) , .Q( key_c_r_9_12 ) );
  DFF_X1 key_c_r_reg_9_13 (.CK( clk ) , .D( key_c_r_8_13 ) , .Q( key_c_r_9_13 ) );
  DFF_X1 key_c_r_reg_9_14 (.CK( clk ) , .D( key_c_r_8_14 ) , .Q( key_c_r_9_14 ) );
  DFF_X1 key_c_r_reg_9_15 (.CK( clk ) , .D( key_c_r_8_15 ) , .Q( key_c_r_9_15 ) );
  DFF_X1 key_c_r_reg_9_16 (.CK( clk ) , .D( key_c_r_8_16 ) , .Q( key_c_r_9_16 ) );
  DFF_X1 key_c_r_reg_9_17 (.CK( clk ) , .D( key_c_r_8_17 ) , .Q( key_c_r_9_17 ) );
  DFF_X1 key_c_r_reg_9_18 (.CK( clk ) , .D( key_c_r_8_18 ) , .Q( key_c_r_9_18 ) );
  DFF_X1 key_c_r_reg_9_19 (.CK( clk ) , .D( key_c_r_8_19 ) , .Q( key_c_r_9_19 ) );
  DFF_X1 key_c_r_reg_9_2 (.CK( clk ) , .D( key_c_r_8_2 ) , .Q( key_c_r_9_2 ) );
  DFF_X1 key_c_r_reg_9_20 (.CK( clk ) , .D( key_c_r_8_20 ) , .Q( key_c_r_9_20 ) );
  DFF_X1 key_c_r_reg_9_21 (.CK( clk ) , .D( key_c_r_8_21 ) , .Q( key_c_r_9_21 ) );
  DFF_X1 key_c_r_reg_9_22 (.CK( clk ) , .D( key_c_r_8_22 ) , .Q( key_c_r_9_22 ) );
  DFF_X1 key_c_r_reg_9_23 (.CK( clk ) , .D( key_c_r_8_23 ) , .Q( key_c_r_9_23 ) );
  DFF_X1 key_c_r_reg_9_24 (.CK( clk ) , .D( key_c_r_8_24 ) , .Q( key_c_r_9_24 ) );
  DFF_X1 key_c_r_reg_9_25 (.CK( clk ) , .D( key_c_r_8_25 ) , .Q( key_c_r_9_25 ) );
  DFF_X1 key_c_r_reg_9_26 (.CK( clk ) , .D( key_c_r_8_26 ) , .Q( key_c_r_9_26 ) );
  DFF_X1 key_c_r_reg_9_27 (.CK( clk ) , .D( key_c_r_8_27 ) , .Q( key_c_r_9_27 ) );
  DFF_X1 key_c_r_reg_9_28 (.CK( clk ) , .D( key_c_r_8_28 ) , .Q( key_c_r_9_28 ) );
  DFF_X1 key_c_r_reg_9_29 (.CK( clk ) , .D( key_c_r_8_29 ) , .Q( key_c_r_9_29 ) );
  DFF_X1 key_c_r_reg_9_3 (.CK( clk ) , .D( key_c_r_8_3 ) , .Q( key_c_r_9_3 ) );
  DFF_X1 key_c_r_reg_9_30 (.CK( clk ) , .D( key_c_r_8_30 ) , .Q( key_c_r_9_30 ) );
  DFF_X1 key_c_r_reg_9_31 (.CK( clk ) , .D( key_c_r_8_31 ) , .Q( key_c_r_9_31 ) );
  DFF_X1 key_c_r_reg_9_32 (.CK( clk ) , .D( key_c_r_8_32 ) , .Q( key_c_r_9_32 ) );
  DFF_X1 key_c_r_reg_9_33 (.CK( clk ) , .D( key_c_r_8_33 ) , .Q( key_c_r_9_33 ) );
  DFF_X1 key_c_r_reg_9_34 (.CK( clk ) , .D( key_c_r_8_34 ) , .Q( key_c_r_9_34 ) );
  DFF_X1 key_c_r_reg_9_35 (.CK( clk ) , .D( key_c_r_8_35 ) , .Q( key_c_r_9_35 ) );
  DFF_X1 key_c_r_reg_9_36 (.CK( clk ) , .D( key_c_r_8_36 ) , .Q( key_c_r_9_36 ) );
  DFF_X1 key_c_r_reg_9_37 (.CK( clk ) , .D( key_c_r_8_37 ) , .Q( key_c_r_9_37 ) );
  DFF_X1 key_c_r_reg_9_38 (.CK( clk ) , .D( key_c_r_8_38 ) , .Q( key_c_r_9_38 ) );
  DFF_X1 key_c_r_reg_9_39 (.CK( clk ) , .D( key_c_r_8_39 ) , .Q( key_c_r_9_39 ) );
  DFF_X1 key_c_r_reg_9_4 (.CK( clk ) , .D( key_c_r_8_4 ) , .Q( key_c_r_9_4 ) );
  DFF_X1 key_c_r_reg_9_40 (.CK( clk ) , .D( key_c_r_8_40 ) , .Q( key_c_r_9_40 ) );
  DFF_X1 key_c_r_reg_9_41 (.CK( clk ) , .D( key_c_r_8_41 ) , .Q( key_c_r_9_41 ) );
  DFF_X1 key_c_r_reg_9_42 (.CK( clk ) , .D( key_c_r_8_42 ) , .Q( key_c_r_9_42 ) );
  DFF_X1 key_c_r_reg_9_43 (.CK( clk ) , .D( key_c_r_8_43 ) , .Q( key_c_r_9_43 ) );
  DFF_X1 key_c_r_reg_9_44 (.CK( clk ) , .D( key_c_r_8_44 ) , .Q( key_c_r_9_44 ) );
  DFF_X1 key_c_r_reg_9_45 (.CK( clk ) , .D( key_c_r_8_45 ) , .Q( key_c_r_9_45 ) );
  DFF_X1 key_c_r_reg_9_46 (.CK( clk ) , .D( key_c_r_8_46 ) , .Q( key_c_r_9_46 ) );
  DFF_X1 key_c_r_reg_9_47 (.CK( clk ) , .D( key_c_r_8_47 ) , .Q( key_c_r_9_47 ) );
  DFF_X1 key_c_r_reg_9_48 (.CK( clk ) , .D( key_c_r_8_48 ) , .Q( key_c_r_9_48 ) );
  DFF_X1 key_c_r_reg_9_49 (.CK( clk ) , .D( key_c_r_8_49 ) , .Q( key_c_r_9_49 ) );
  DFF_X1 key_c_r_reg_9_5 (.CK( clk ) , .D( key_c_r_8_5 ) , .Q( key_c_r_9_5 ) );
  DFF_X1 key_c_r_reg_9_50 (.CK( clk ) , .D( key_c_r_8_50 ) , .Q( key_c_r_9_50 ) );
  DFF_X1 key_c_r_reg_9_51 (.CK( clk ) , .D( key_c_r_8_51 ) , .Q( key_c_r_9_51 ) );
  DFF_X1 key_c_r_reg_9_52 (.CK( clk ) , .D( key_c_r_8_52 ) , .Q( key_c_r_9_52 ) );
  DFF_X1 key_c_r_reg_9_53 (.CK( clk ) , .D( key_c_r_8_53 ) , .Q( key_c_r_9_53 ) );
  DFF_X1 key_c_r_reg_9_54 (.CK( clk ) , .D( key_c_r_8_54 ) , .Q( key_c_r_9_54 ) );
  DFF_X1 key_c_r_reg_9_55 (.CK( clk ) , .D( key_c_r_8_55 ) , .Q( key_c_r_9_55 ) );
  DFF_X1 key_c_r_reg_9_6 (.CK( clk ) , .D( key_c_r_8_6 ) , .Q( key_c_r_9_6 ) );
  DFF_X1 key_c_r_reg_9_7 (.CK( clk ) , .D( key_c_r_8_7 ) , .Q( key_c_r_9_7 ) );
  DFF_X1 key_c_r_reg_9_8 (.CK( clk ) , .D( key_c_r_8_8 ) , .Q( key_c_r_9_8 ) );
  DFF_X1 key_c_r_reg_9_9 (.CK( clk ) , .D( key_c_r_8_9 ) , .Q( key_c_r_9_9 ) );
  DFF_X1 u0_L0_reg_1 (.CK( clk ) , .Q( u0_L0_1 ) , .D( u0_desIn_r_7 ) );
  DFF_X1 u0_L0_reg_10 (.CK( clk ) , .Q( u0_L0_10 ) , .D( u0_desIn_r_13 ) );
  DFF_X1 u0_L0_reg_11 (.CK( clk ) , .Q( u0_L0_11 ) , .D( u0_desIn_r_21 ) );
  DFF_X1 u0_L0_reg_12 (.CK( clk ) , .Q( u0_L0_12 ) , .D( u0_desIn_r_29 ) );
  DFF_X1 u0_L0_reg_13 (.CK( clk ) , .Q( u0_L0_13 ) , .D( u0_desIn_r_37 ) );
  DFF_X1 u0_L0_reg_14 (.CK( clk ) , .Q( u0_L0_14 ) , .D( u0_desIn_r_45 ) );
  DFF_X1 u0_L0_reg_15 (.CK( clk ) , .Q( u0_L0_15 ) , .D( u0_desIn_r_53 ) );
  DFF_X1 u0_L0_reg_16 (.CK( clk ) , .Q( u0_L0_16 ) , .D( u0_desIn_r_61 ) );
  DFF_X1 u0_L0_reg_17 (.CK( clk ) , .Q( u0_L0_17 ) , .D( u0_desIn_r_3 ) );
  DFF_X1 u0_L0_reg_18 (.CK( clk ) , .Q( u0_L0_18 ) , .D( u0_desIn_r_11 ) );
  DFF_X1 u0_L0_reg_19 (.CK( clk ) , .Q( u0_L0_19 ) , .D( u0_desIn_r_19 ) );
  DFF_X1 u0_L0_reg_2 (.CK( clk ) , .Q( u0_L0_2 ) , .D( u0_desIn_r_15 ) );
  DFF_X1 u0_L0_reg_20 (.CK( clk ) , .Q( u0_L0_20 ) , .D( u0_desIn_r_27 ) );
  DFF_X1 u0_L0_reg_21 (.CK( clk ) , .Q( u0_L0_21 ) , .D( u0_desIn_r_35 ) );
  DFF_X1 u0_L0_reg_22 (.CK( clk ) , .Q( u0_L0_22 ) , .D( u0_desIn_r_43 ) );
  DFF_X1 u0_L0_reg_23 (.CK( clk ) , .Q( u0_L0_23 ) , .D( u0_desIn_r_51 ) );
  DFF_X1 u0_L0_reg_24 (.CK( clk ) , .Q( u0_L0_24 ) , .D( u0_desIn_r_59 ) );
  DFF_X1 u0_L0_reg_25 (.CK( clk ) , .Q( u0_L0_25 ) , .D( u0_desIn_r_1 ) );
  DFF_X1 u0_L0_reg_26 (.CK( clk ) , .Q( u0_L0_26 ) , .D( u0_desIn_r_9 ) );
  DFF_X1 u0_L0_reg_27 (.CK( clk ) , .Q( u0_L0_27 ) , .D( u0_desIn_r_17 ) );
  DFF_X1 u0_L0_reg_28 (.CK( clk ) , .Q( u0_L0_28 ) , .D( u0_desIn_r_25 ) );
  DFF_X1 u0_L0_reg_29 (.CK( clk ) , .Q( u0_L0_29 ) , .D( u0_desIn_r_33 ) );
  DFF_X1 u0_L0_reg_3 (.CK( clk ) , .Q( u0_L0_3 ) , .D( u0_desIn_r_23 ) );
  DFF_X1 u0_L0_reg_30 (.CK( clk ) , .Q( u0_L0_30 ) , .D( u0_desIn_r_41 ) );
  DFF_X1 u0_L0_reg_31 (.CK( clk ) , .Q( u0_L0_31 ) , .D( u0_desIn_r_49 ) );
  DFF_X1 u0_L0_reg_32 (.CK( clk ) , .Q( u0_L0_32 ) , .D( u0_desIn_r_57 ) );
  DFF_X1 u0_L0_reg_4 (.CK( clk ) , .Q( u0_L0_4 ) , .D( u0_desIn_r_31 ) );
  DFF_X1 u0_L0_reg_5 (.CK( clk ) , .Q( u0_L0_5 ) , .D( u0_desIn_r_39 ) );
  DFF_X1 u0_L0_reg_6 (.CK( clk ) , .Q( u0_L0_6 ) , .D( u0_desIn_r_47 ) );
  DFF_X1 u0_L0_reg_7 (.CK( clk ) , .Q( u0_L0_7 ) , .D( u0_desIn_r_55 ) );
  DFF_X1 u0_L0_reg_8 (.CK( clk ) , .Q( u0_L0_8 ) , .D( u0_desIn_r_63 ) );
  DFF_X1 u0_L0_reg_9 (.CK( clk ) , .Q( u0_L0_9 ) , .D( u0_desIn_r_5 ) );
  DFF_X1 u0_L10_reg_1 (.CK( clk ) , .Q( u0_L10_1 ) , .D( u0_R9_1 ) );
  DFF_X1 u0_L10_reg_10 (.CK( clk ) , .Q( u0_L10_10 ) , .D( u0_R9_10 ) );
  DFF_X1 u0_L10_reg_11 (.CK( clk ) , .Q( u0_L10_11 ) , .D( u0_R9_11 ) );
  DFF_X1 u0_L10_reg_12 (.CK( clk ) , .Q( u0_L10_12 ) , .D( u0_R9_12 ) );
  DFF_X1 u0_L10_reg_13 (.CK( clk ) , .Q( u0_L10_13 ) , .D( u0_R9_13 ) );
  DFF_X1 u0_L10_reg_14 (.CK( clk ) , .Q( u0_L10_14 ) , .D( u0_R9_14 ) );
  DFF_X1 u0_L10_reg_15 (.CK( clk ) , .Q( u0_L10_15 ) , .D( u0_R9_15 ) );
  DFF_X1 u0_L10_reg_16 (.CK( clk ) , .Q( u0_L10_16 ) , .D( u0_R9_16 ) );
  DFF_X1 u0_L10_reg_17 (.CK( clk ) , .Q( u0_L10_17 ) , .D( u0_R9_17 ) );
  DFF_X1 u0_L10_reg_18 (.CK( clk ) , .Q( u0_L10_18 ) , .D( u0_R9_18 ) );
  DFF_X1 u0_L10_reg_19 (.CK( clk ) , .Q( u0_L10_19 ) , .D( u0_R9_19 ) );
  DFF_X1 u0_L10_reg_2 (.CK( clk ) , .Q( u0_L10_2 ) , .D( u0_R9_2 ) );
  DFF_X1 u0_L10_reg_20 (.CK( clk ) , .Q( u0_L10_20 ) , .D( u0_R9_20 ) );
  DFF_X1 u0_L10_reg_21 (.CK( clk ) , .Q( u0_L10_21 ) , .D( u0_R9_21 ) );
  DFF_X1 u0_L10_reg_22 (.CK( clk ) , .Q( u0_L10_22 ) , .D( u0_R9_22 ) );
  DFF_X1 u0_L10_reg_23 (.CK( clk ) , .Q( u0_L10_23 ) , .D( u0_R9_23 ) );
  DFF_X1 u0_L10_reg_24 (.CK( clk ) , .Q( u0_L10_24 ) , .D( u0_R9_24 ) );
  DFF_X1 u0_L10_reg_25 (.CK( clk ) , .Q( u0_L10_25 ) , .D( u0_R9_25 ) );
  DFF_X1 u0_L10_reg_26 (.CK( clk ) , .Q( u0_L10_26 ) , .D( u0_R9_26 ) );
  DFF_X1 u0_L10_reg_27 (.CK( clk ) , .Q( u0_L10_27 ) , .D( u0_R9_27 ) );
  DFF_X1 u0_L10_reg_28 (.CK( clk ) , .Q( u0_L10_28 ) , .D( u0_R9_28 ) );
  DFF_X1 u0_L10_reg_29 (.CK( clk ) , .Q( u0_L10_29 ) , .D( u0_R9_29 ) );
  DFF_X1 u0_L10_reg_3 (.CK( clk ) , .Q( u0_L10_3 ) , .D( u0_R9_3 ) );
  DFF_X1 u0_L10_reg_30 (.CK( clk ) , .Q( u0_L10_30 ) , .D( u0_R9_30 ) );
  DFF_X1 u0_L10_reg_31 (.CK( clk ) , .Q( u0_L10_31 ) , .D( u0_R9_31 ) );
  DFF_X1 u0_L10_reg_32 (.CK( clk ) , .Q( u0_L10_32 ) , .D( u0_R9_32 ) );
  DFF_X1 u0_L10_reg_4 (.CK( clk ) , .Q( u0_L10_4 ) , .D( u0_R9_4 ) );
  DFF_X1 u0_L10_reg_5 (.CK( clk ) , .Q( u0_L10_5 ) , .D( u0_R9_5 ) );
  DFF_X1 u0_L10_reg_6 (.CK( clk ) , .Q( u0_L10_6 ) , .D( u0_R9_6 ) );
  DFF_X1 u0_L10_reg_7 (.CK( clk ) , .Q( u0_L10_7 ) , .D( u0_R9_7 ) );
  DFF_X1 u0_L10_reg_8 (.CK( clk ) , .Q( u0_L10_8 ) , .D( u0_R9_8 ) );
  DFF_X1 u0_L10_reg_9 (.CK( clk ) , .Q( u0_L10_9 ) , .D( u0_R9_9 ) );
  DFF_X1 u0_L11_reg_1 (.CK( clk ) , .Q( u0_L11_1 ) , .D( u0_R10_1 ) );
  DFF_X1 u0_L11_reg_10 (.CK( clk ) , .Q( u0_L11_10 ) , .D( u0_R10_10 ) );
  DFF_X1 u0_L11_reg_11 (.CK( clk ) , .Q( u0_L11_11 ) , .D( u0_R10_11 ) );
  DFF_X1 u0_L11_reg_12 (.CK( clk ) , .Q( u0_L11_12 ) , .D( u0_R10_12 ) );
  DFF_X1 u0_L11_reg_13 (.CK( clk ) , .Q( u0_L11_13 ) , .D( u0_R10_13 ) );
  DFF_X1 u0_L11_reg_14 (.CK( clk ) , .Q( u0_L11_14 ) , .D( u0_R10_14 ) );
  DFF_X1 u0_L11_reg_15 (.CK( clk ) , .Q( u0_L11_15 ) , .D( u0_R10_15 ) );
  DFF_X1 u0_L11_reg_16 (.CK( clk ) , .Q( u0_L11_16 ) , .D( u0_R10_16 ) );
  DFF_X1 u0_L11_reg_17 (.CK( clk ) , .Q( u0_L11_17 ) , .D( u0_R10_17 ) );
  DFF_X1 u0_L11_reg_18 (.CK( clk ) , .Q( u0_L11_18 ) , .D( u0_R10_18 ) );
  DFF_X1 u0_L11_reg_19 (.CK( clk ) , .Q( u0_L11_19 ) , .D( u0_R10_19 ) );
  DFF_X1 u0_L11_reg_2 (.CK( clk ) , .Q( u0_L11_2 ) , .D( u0_R10_2 ) );
  DFF_X1 u0_L11_reg_20 (.CK( clk ) , .Q( u0_L11_20 ) , .D( u0_R10_20 ) );
  DFF_X1 u0_L11_reg_21 (.CK( clk ) , .Q( u0_L11_21 ) , .D( u0_R10_21 ) );
  DFF_X1 u0_L11_reg_22 (.CK( clk ) , .Q( u0_L11_22 ) , .D( u0_R10_22 ) );
  DFF_X1 u0_L11_reg_23 (.CK( clk ) , .Q( u0_L11_23 ) , .D( u0_R10_23 ) );
  DFF_X1 u0_L11_reg_24 (.CK( clk ) , .Q( u0_L11_24 ) , .D( u0_R10_24 ) );
  DFF_X1 u0_L11_reg_25 (.CK( clk ) , .Q( u0_L11_25 ) , .D( u0_R10_25 ) );
  DFF_X1 u0_L11_reg_26 (.CK( clk ) , .Q( u0_L11_26 ) , .D( u0_R10_26 ) );
  DFF_X1 u0_L11_reg_27 (.CK( clk ) , .Q( u0_L11_27 ) , .D( u0_R10_27 ) );
  DFF_X1 u0_L11_reg_28 (.CK( clk ) , .Q( u0_L11_28 ) , .D( u0_R10_28 ) );
  DFF_X1 u0_L11_reg_29 (.CK( clk ) , .Q( u0_L11_29 ) , .D( u0_R10_29 ) );
  DFF_X1 u0_L11_reg_3 (.CK( clk ) , .Q( u0_L11_3 ) , .D( u0_R10_3 ) );
  DFF_X1 u0_L11_reg_30 (.CK( clk ) , .Q( u0_L11_30 ) , .D( u0_R10_30 ) );
  DFF_X1 u0_L11_reg_31 (.CK( clk ) , .Q( u0_L11_31 ) , .D( u0_R10_31 ) );
  DFF_X1 u0_L11_reg_32 (.CK( clk ) , .Q( u0_L11_32 ) , .D( u0_R10_32 ) );
  DFF_X1 u0_L11_reg_4 (.CK( clk ) , .Q( u0_L11_4 ) , .D( u0_R10_4 ) );
  DFF_X1 u0_L11_reg_5 (.CK( clk ) , .Q( u0_L11_5 ) , .D( u0_R10_5 ) );
  DFF_X1 u0_L11_reg_6 (.CK( clk ) , .Q( u0_L11_6 ) , .D( u0_R10_6 ) );
  DFF_X1 u0_L11_reg_7 (.CK( clk ) , .Q( u0_L11_7 ) , .D( u0_R10_7 ) );
  DFF_X1 u0_L11_reg_8 (.CK( clk ) , .Q( u0_L11_8 ) , .D( u0_R10_8 ) );
  DFF_X1 u0_L11_reg_9 (.CK( clk ) , .Q( u0_L11_9 ) , .D( u0_R10_9 ) );
  DFF_X1 u0_L12_reg_1 (.CK( clk ) , .Q( u0_L12_1 ) , .D( u0_R11_1 ) );
  DFF_X1 u0_L12_reg_10 (.CK( clk ) , .Q( u0_L12_10 ) , .D( u0_R11_10 ) );
  DFF_X1 u0_L12_reg_11 (.CK( clk ) , .Q( u0_L12_11 ) , .D( u0_R11_11 ) );
  DFF_X1 u0_L12_reg_12 (.CK( clk ) , .Q( u0_L12_12 ) , .D( u0_R11_12 ) );
  DFF_X1 u0_L12_reg_13 (.CK( clk ) , .Q( u0_L12_13 ) , .D( u0_R11_13 ) );
  DFF_X1 u0_L12_reg_14 (.CK( clk ) , .Q( u0_L12_14 ) , .D( u0_R11_14 ) );
  DFF_X1 u0_L12_reg_15 (.CK( clk ) , .Q( u0_L12_15 ) , .D( u0_R11_15 ) );
  DFF_X1 u0_L12_reg_16 (.CK( clk ) , .Q( u0_L12_16 ) , .D( u0_R11_16 ) );
  DFF_X1 u0_L12_reg_17 (.CK( clk ) , .Q( u0_L12_17 ) , .D( u0_R11_17 ) );
  DFF_X1 u0_L12_reg_18 (.CK( clk ) , .Q( u0_L12_18 ) , .D( u0_R11_18 ) );
  DFF_X1 u0_L12_reg_19 (.CK( clk ) , .Q( u0_L12_19 ) , .D( u0_R11_19 ) );
  DFF_X1 u0_L12_reg_2 (.CK( clk ) , .Q( u0_L12_2 ) , .D( u0_R11_2 ) );
  DFF_X1 u0_L12_reg_20 (.CK( clk ) , .Q( u0_L12_20 ) , .D( u0_R11_20 ) );
  DFF_X1 u0_L12_reg_21 (.CK( clk ) , .Q( u0_L12_21 ) , .D( u0_R11_21 ) );
  DFF_X1 u0_L12_reg_22 (.CK( clk ) , .Q( u0_L12_22 ) , .D( u0_R11_22 ) );
  DFF_X1 u0_L12_reg_23 (.CK( clk ) , .Q( u0_L12_23 ) , .D( u0_R11_23 ) );
  DFF_X1 u0_L12_reg_24 (.CK( clk ) , .Q( u0_L12_24 ) , .D( u0_R11_24 ) );
  DFF_X1 u0_L12_reg_25 (.CK( clk ) , .Q( u0_L12_25 ) , .D( u0_R11_25 ) );
  DFF_X1 u0_L12_reg_26 (.CK( clk ) , .Q( u0_L12_26 ) , .D( u0_R11_26 ) );
  DFF_X1 u0_L12_reg_27 (.CK( clk ) , .Q( u0_L12_27 ) , .D( u0_R11_27 ) );
  DFF_X1 u0_L12_reg_28 (.CK( clk ) , .Q( u0_L12_28 ) , .D( u0_R11_28 ) );
  DFF_X1 u0_L12_reg_29 (.CK( clk ) , .Q( u0_L12_29 ) , .D( u0_R11_29 ) );
  DFF_X1 u0_L12_reg_3 (.CK( clk ) , .Q( u0_L12_3 ) , .D( u0_R11_3 ) );
  DFF_X1 u0_L12_reg_30 (.CK( clk ) , .Q( u0_L12_30 ) , .D( u0_R11_30 ) );
  DFF_X1 u0_L12_reg_31 (.CK( clk ) , .Q( u0_L12_31 ) , .D( u0_R11_31 ) );
  DFF_X1 u0_L12_reg_32 (.CK( clk ) , .Q( u0_L12_32 ) , .D( u0_R11_32 ) );
  DFF_X1 u0_L12_reg_4 (.CK( clk ) , .Q( u0_L12_4 ) , .D( u0_R11_4 ) );
  DFF_X1 u0_L12_reg_5 (.CK( clk ) , .Q( u0_L12_5 ) , .D( u0_R11_5 ) );
  DFF_X1 u0_L12_reg_6 (.CK( clk ) , .Q( u0_L12_6 ) , .D( u0_R11_6 ) );
  DFF_X1 u0_L12_reg_7 (.CK( clk ) , .Q( u0_L12_7 ) , .D( u0_R11_7 ) );
  DFF_X1 u0_L12_reg_8 (.CK( clk ) , .Q( u0_L12_8 ) , .D( u0_R11_8 ) );
  DFF_X1 u0_L12_reg_9 (.CK( clk ) , .Q( u0_L12_9 ) , .D( u0_R11_9 ) );
  DFF_X1 u0_L13_reg_1 (.CK( clk ) , .Q( u0_L13_1 ) , .D( u0_R12_1 ) );
  DFF_X1 u0_L13_reg_10 (.CK( clk ) , .Q( u0_L13_10 ) , .D( u0_R12_10 ) );
  DFF_X1 u0_L13_reg_11 (.CK( clk ) , .Q( u0_L13_11 ) , .D( u0_R12_11 ) );
  DFF_X1 u0_L13_reg_12 (.CK( clk ) , .Q( u0_L13_12 ) , .D( u0_R12_12 ) );
  DFF_X1 u0_L13_reg_13 (.CK( clk ) , .Q( u0_L13_13 ) , .D( u0_R12_13 ) );
  DFF_X1 u0_L13_reg_14 (.CK( clk ) , .Q( u0_L13_14 ) , .D( u0_R12_14 ) );
  DFF_X1 u0_L13_reg_15 (.CK( clk ) , .Q( u0_L13_15 ) , .D( u0_R12_15 ) );
  DFF_X1 u0_L13_reg_16 (.CK( clk ) , .Q( u0_L13_16 ) , .D( u0_R12_16 ) );
  DFF_X1 u0_L13_reg_17 (.CK( clk ) , .Q( u0_L13_17 ) , .D( u0_R12_17 ) );
  DFF_X1 u0_L13_reg_18 (.CK( clk ) , .Q( u0_L13_18 ) , .D( u0_R12_18 ) );
  DFF_X1 u0_L13_reg_19 (.CK( clk ) , .Q( u0_L13_19 ) , .D( u0_R12_19 ) );
  DFF_X1 u0_L13_reg_2 (.CK( clk ) , .Q( u0_L13_2 ) , .D( u0_R12_2 ) );
  DFF_X1 u0_L13_reg_20 (.CK( clk ) , .Q( u0_L13_20 ) , .D( u0_R12_20 ) );
  DFF_X1 u0_L13_reg_21 (.CK( clk ) , .Q( u0_L13_21 ) , .D( u0_R12_21 ) );
  DFF_X1 u0_L13_reg_22 (.CK( clk ) , .Q( u0_L13_22 ) , .D( u0_R12_22 ) );
  DFF_X1 u0_L13_reg_23 (.CK( clk ) , .Q( u0_L13_23 ) , .D( u0_R12_23 ) );
  DFF_X1 u0_L13_reg_24 (.CK( clk ) , .Q( u0_L13_24 ) , .D( u0_R12_24 ) );
  DFF_X1 u0_L13_reg_25 (.CK( clk ) , .Q( u0_L13_25 ) , .D( u0_R12_25 ) );
  DFF_X1 u0_L13_reg_26 (.CK( clk ) , .Q( u0_L13_26 ) , .D( u0_R12_26 ) );
  DFF_X1 u0_L13_reg_27 (.CK( clk ) , .Q( u0_L13_27 ) , .D( u0_R12_27 ) );
  DFF_X1 u0_L13_reg_28 (.CK( clk ) , .Q( u0_L13_28 ) , .D( u0_R12_28 ) );
  DFF_X1 u0_L13_reg_29 (.CK( clk ) , .Q( u0_L13_29 ) , .D( u0_R12_29 ) );
  DFF_X1 u0_L13_reg_3 (.CK( clk ) , .Q( u0_L13_3 ) , .D( u0_R12_3 ) );
  DFF_X1 u0_L13_reg_30 (.CK( clk ) , .Q( u0_L13_30 ) , .D( u0_R12_30 ) );
  DFF_X1 u0_L13_reg_31 (.CK( clk ) , .Q( u0_L13_31 ) , .D( u0_R12_31 ) );
  DFF_X1 u0_L13_reg_32 (.CK( clk ) , .Q( u0_L13_32 ) , .D( u0_R12_32 ) );
  DFF_X1 u0_L13_reg_4 (.CK( clk ) , .Q( u0_L13_4 ) , .D( u0_R12_4 ) );
  DFF_X1 u0_L13_reg_5 (.CK( clk ) , .Q( u0_L13_5 ) , .D( u0_R12_5 ) );
  DFF_X1 u0_L13_reg_6 (.CK( clk ) , .Q( u0_L13_6 ) , .D( u0_R12_6 ) );
  DFF_X1 u0_L13_reg_7 (.CK( clk ) , .Q( u0_L13_7 ) , .D( u0_R12_7 ) );
  DFF_X1 u0_L13_reg_8 (.CK( clk ) , .Q( u0_L13_8 ) , .D( u0_R12_8 ) );
  DFF_X1 u0_L13_reg_9 (.CK( clk ) , .Q( u0_L13_9 ) , .D( u0_R12_9 ) );
  DFF_X1 u0_L14_reg_1 (.CK( clk ) , .Q( u0_L14_1 ) , .D( u0_R13_1 ) );
  DFF_X1 u0_L14_reg_10 (.CK( clk ) , .Q( u0_L14_10 ) , .D( u0_R13_10 ) );
  DFF_X1 u0_L14_reg_11 (.CK( clk ) , .Q( u0_L14_11 ) , .D( u0_R13_11 ) );
  DFF_X1 u0_L14_reg_12 (.CK( clk ) , .Q( u0_L14_12 ) , .D( u0_R13_12 ) );
  DFF_X1 u0_L14_reg_13 (.CK( clk ) , .Q( u0_L14_13 ) , .D( u0_R13_13 ) );
  DFF_X1 u0_L14_reg_14 (.CK( clk ) , .Q( u0_L14_14 ) , .D( u0_R13_14 ) );
  DFF_X1 u0_L14_reg_15 (.CK( clk ) , .Q( u0_L14_15 ) , .D( u0_R13_15 ) );
  DFF_X1 u0_L14_reg_16 (.CK( clk ) , .Q( u0_L14_16 ) , .D( u0_R13_16 ) );
  DFF_X1 u0_L14_reg_17 (.CK( clk ) , .Q( u0_L14_17 ) , .D( u0_R13_17 ) );
  DFF_X1 u0_L14_reg_18 (.CK( clk ) , .Q( u0_L14_18 ) , .D( u0_R13_18 ) );
  DFF_X1 u0_L14_reg_19 (.CK( clk ) , .Q( u0_L14_19 ) , .D( u0_R13_19 ) );
  DFF_X1 u0_L14_reg_2 (.CK( clk ) , .Q( u0_L14_2 ) , .D( u0_R13_2 ) );
  DFF_X1 u0_L14_reg_20 (.CK( clk ) , .Q( u0_L14_20 ) , .D( u0_R13_20 ) );
  DFF_X1 u0_L14_reg_21 (.CK( clk ) , .Q( u0_L14_21 ) , .D( u0_R13_21 ) );
  DFF_X1 u0_L14_reg_22 (.CK( clk ) , .Q( u0_L14_22 ) , .D( u0_R13_22 ) );
  DFF_X1 u0_L14_reg_23 (.CK( clk ) , .Q( u0_L14_23 ) , .D( u0_R13_23 ) );
  DFF_X1 u0_L14_reg_24 (.CK( clk ) , .Q( u0_L14_24 ) , .D( u0_R13_24 ) );
  DFF_X1 u0_L14_reg_25 (.CK( clk ) , .Q( u0_L14_25 ) , .D( u0_R13_25 ) );
  DFF_X1 u0_L14_reg_26 (.CK( clk ) , .Q( u0_L14_26 ) , .D( u0_R13_26 ) );
  DFF_X1 u0_L14_reg_27 (.CK( clk ) , .Q( u0_L14_27 ) , .D( u0_R13_27 ) );
  DFF_X1 u0_L14_reg_28 (.CK( clk ) , .Q( u0_L14_28 ) , .D( u0_R13_28 ) );
  DFF_X1 u0_L14_reg_29 (.CK( clk ) , .Q( u0_L14_29 ) , .D( u0_R13_29 ) );
  DFF_X1 u0_L14_reg_3 (.CK( clk ) , .Q( u0_L14_3 ) , .D( u0_R13_3 ) );
  DFF_X1 u0_L14_reg_30 (.CK( clk ) , .Q( u0_L14_30 ) , .D( u0_R13_30 ) );
  DFF_X1 u0_L14_reg_31 (.CK( clk ) , .Q( u0_L14_31 ) , .D( u0_R13_31 ) );
  DFF_X1 u0_L14_reg_32 (.CK( clk ) , .Q( u0_L14_32 ) , .D( u0_R13_32 ) );
  DFF_X1 u0_L14_reg_4 (.CK( clk ) , .Q( u0_L14_4 ) , .D( u0_R13_4 ) );
  DFF_X1 u0_L14_reg_5 (.CK( clk ) , .Q( u0_L14_5 ) , .D( u0_R13_5 ) );
  DFF_X1 u0_L14_reg_6 (.CK( clk ) , .Q( u0_L14_6 ) , .D( u0_R13_6 ) );
  DFF_X1 u0_L14_reg_7 (.CK( clk ) , .Q( u0_L14_7 ) , .D( u0_R13_7 ) );
  DFF_X1 u0_L14_reg_8 (.CK( clk ) , .Q( u0_L14_8 ) , .D( u0_R13_8 ) );
  DFF_X1 u0_L14_reg_9 (.CK( clk ) , .Q( u0_L14_9 ) , .D( u0_R13_9 ) );
  DFF_X1 u0_L1_reg_1 (.CK( clk ) , .Q( u0_L1_1 ) , .D( u0_R0_1 ) );
  DFF_X1 u0_L1_reg_10 (.CK( clk ) , .Q( u0_L1_10 ) , .D( u0_R0_10 ) );
  DFF_X1 u0_L1_reg_11 (.CK( clk ) , .Q( u0_L1_11 ) , .D( u0_R0_11 ) );
  DFF_X1 u0_L1_reg_12 (.CK( clk ) , .Q( u0_L1_12 ) , .D( u0_R0_12 ) );
  DFF_X1 u0_L1_reg_13 (.CK( clk ) , .Q( u0_L1_13 ) , .D( u0_R0_13 ) );
  DFF_X1 u0_L1_reg_14 (.CK( clk ) , .Q( u0_L1_14 ) , .D( u0_R0_14 ) );
  DFF_X1 u0_L1_reg_15 (.CK( clk ) , .Q( u0_L1_15 ) , .D( u0_R0_15 ) );
  DFF_X1 u0_L1_reg_16 (.CK( clk ) , .Q( u0_L1_16 ) , .D( u0_R0_16 ) );
  DFF_X1 u0_L1_reg_17 (.CK( clk ) , .Q( u0_L1_17 ) , .D( u0_R0_17 ) );
  DFF_X1 u0_L1_reg_18 (.CK( clk ) , .Q( u0_L1_18 ) , .D( u0_R0_18 ) );
  DFF_X1 u0_L1_reg_19 (.CK( clk ) , .Q( u0_L1_19 ) , .D( u0_R0_19 ) );
  DFF_X1 u0_L1_reg_2 (.CK( clk ) , .Q( u0_L1_2 ) , .D( u0_R0_2 ) );
  DFF_X1 u0_L1_reg_20 (.CK( clk ) , .Q( u0_L1_20 ) , .D( u0_R0_20 ) );
  DFF_X1 u0_L1_reg_21 (.CK( clk ) , .Q( u0_L1_21 ) , .D( u0_R0_21 ) );
  DFF_X1 u0_L1_reg_22 (.CK( clk ) , .Q( u0_L1_22 ) , .D( u0_R0_22 ) );
  DFF_X1 u0_L1_reg_23 (.CK( clk ) , .Q( u0_L1_23 ) , .D( u0_R0_23 ) );
  DFF_X1 u0_L1_reg_24 (.CK( clk ) , .Q( u0_L1_24 ) , .D( u0_R0_24 ) );
  DFF_X1 u0_L1_reg_25 (.CK( clk ) , .Q( u0_L1_25 ) , .D( u0_R0_25 ) );
  DFF_X1 u0_L1_reg_26 (.CK( clk ) , .Q( u0_L1_26 ) , .D( u0_R0_26 ) );
  DFF_X1 u0_L1_reg_27 (.CK( clk ) , .Q( u0_L1_27 ) , .D( u0_R0_27 ) );
  DFF_X1 u0_L1_reg_28 (.CK( clk ) , .Q( u0_L1_28 ) , .D( u0_R0_28 ) );
  DFF_X1 u0_L1_reg_29 (.CK( clk ) , .Q( u0_L1_29 ) , .D( u0_R0_29 ) );
  DFF_X1 u0_L1_reg_3 (.CK( clk ) , .Q( u0_L1_3 ) , .D( u0_R0_3 ) );
  DFF_X1 u0_L1_reg_30 (.CK( clk ) , .Q( u0_L1_30 ) , .D( u0_R0_30 ) );
  DFF_X1 u0_L1_reg_31 (.CK( clk ) , .Q( u0_L1_31 ) , .D( u0_R0_31 ) );
  DFF_X1 u0_L1_reg_32 (.CK( clk ) , .Q( u0_L1_32 ) , .D( u0_R0_32 ) );
  DFF_X1 u0_L1_reg_4 (.CK( clk ) , .Q( u0_L1_4 ) , .D( u0_R0_4 ) );
  DFF_X1 u0_L1_reg_5 (.CK( clk ) , .Q( u0_L1_5 ) , .D( u0_R0_5 ) );
  DFF_X1 u0_L1_reg_6 (.CK( clk ) , .Q( u0_L1_6 ) , .D( u0_R0_6 ) );
  DFF_X1 u0_L1_reg_7 (.CK( clk ) , .Q( u0_L1_7 ) , .D( u0_R0_7 ) );
  DFF_X1 u0_L1_reg_8 (.CK( clk ) , .Q( u0_L1_8 ) , .D( u0_R0_8 ) );
  DFF_X1 u0_L1_reg_9 (.CK( clk ) , .Q( u0_L1_9 ) , .D( u0_R0_9 ) );
  DFF_X1 u0_L2_reg_1 (.CK( clk ) , .Q( u0_L2_1 ) , .D( u0_R1_1 ) );
  DFF_X1 u0_L2_reg_10 (.CK( clk ) , .Q( u0_L2_10 ) , .D( u0_R1_10 ) );
  DFF_X1 u0_L2_reg_11 (.CK( clk ) , .Q( u0_L2_11 ) , .D( u0_R1_11 ) );
  DFF_X1 u0_L2_reg_12 (.CK( clk ) , .Q( u0_L2_12 ) , .D( u0_R1_12 ) );
  DFF_X1 u0_L2_reg_13 (.CK( clk ) , .Q( u0_L2_13 ) , .D( u0_R1_13 ) );
  DFF_X1 u0_L2_reg_14 (.CK( clk ) , .Q( u0_L2_14 ) , .D( u0_R1_14 ) );
  DFF_X1 u0_L2_reg_15 (.CK( clk ) , .Q( u0_L2_15 ) , .D( u0_R1_15 ) );
  DFF_X1 u0_L2_reg_16 (.CK( clk ) , .Q( u0_L2_16 ) , .D( u0_R1_16 ) );
  DFF_X1 u0_L2_reg_17 (.CK( clk ) , .Q( u0_L2_17 ) , .D( u0_R1_17 ) );
  DFF_X1 u0_L2_reg_18 (.CK( clk ) , .Q( u0_L2_18 ) , .D( u0_R1_18 ) );
  DFF_X1 u0_L2_reg_19 (.CK( clk ) , .Q( u0_L2_19 ) , .D( u0_R1_19 ) );
  DFF_X1 u0_L2_reg_2 (.CK( clk ) , .Q( u0_L2_2 ) , .D( u0_R1_2 ) );
  DFF_X1 u0_L2_reg_20 (.CK( clk ) , .Q( u0_L2_20 ) , .D( u0_R1_20 ) );
  DFF_X1 u0_L2_reg_21 (.CK( clk ) , .Q( u0_L2_21 ) , .D( u0_R1_21 ) );
  DFF_X1 u0_L2_reg_22 (.CK( clk ) , .Q( u0_L2_22 ) , .D( u0_R1_22 ) );
  DFF_X1 u0_L2_reg_23 (.CK( clk ) , .Q( u0_L2_23 ) , .D( u0_R1_23 ) );
  DFF_X1 u0_L2_reg_24 (.CK( clk ) , .Q( u0_L2_24 ) , .D( u0_R1_24 ) );
  DFF_X1 u0_L2_reg_25 (.CK( clk ) , .Q( u0_L2_25 ) , .D( u0_R1_25 ) );
  DFF_X1 u0_L2_reg_26 (.CK( clk ) , .Q( u0_L2_26 ) , .D( u0_R1_26 ) );
  DFF_X1 u0_L2_reg_27 (.CK( clk ) , .Q( u0_L2_27 ) , .D( u0_R1_27 ) );
  DFF_X1 u0_L2_reg_28 (.CK( clk ) , .Q( u0_L2_28 ) , .D( u0_R1_28 ) );
  DFF_X1 u0_L2_reg_29 (.CK( clk ) , .Q( u0_L2_29 ) , .D( u0_R1_29 ) );
  DFF_X1 u0_L2_reg_3 (.CK( clk ) , .Q( u0_L2_3 ) , .D( u0_R1_3 ) );
  DFF_X1 u0_L2_reg_30 (.CK( clk ) , .Q( u0_L2_30 ) , .D( u0_R1_30 ) );
  DFF_X1 u0_L2_reg_31 (.CK( clk ) , .Q( u0_L2_31 ) , .D( u0_R1_31 ) );
  DFF_X1 u0_L2_reg_32 (.CK( clk ) , .Q( u0_L2_32 ) , .D( u0_R1_32 ) );
  DFF_X1 u0_L2_reg_4 (.CK( clk ) , .Q( u0_L2_4 ) , .D( u0_R1_4 ) );
  DFF_X1 u0_L2_reg_5 (.CK( clk ) , .Q( u0_L2_5 ) , .D( u0_R1_5 ) );
  DFF_X1 u0_L2_reg_6 (.CK( clk ) , .Q( u0_L2_6 ) , .D( u0_R1_6 ) );
  DFF_X1 u0_L2_reg_7 (.CK( clk ) , .Q( u0_L2_7 ) , .D( u0_R1_7 ) );
  DFF_X1 u0_L2_reg_8 (.CK( clk ) , .Q( u0_L2_8 ) , .D( u0_R1_8 ) );
  DFF_X1 u0_L2_reg_9 (.CK( clk ) , .Q( u0_L2_9 ) , .D( u0_R1_9 ) );
  DFF_X1 u0_L3_reg_1 (.CK( clk ) , .Q( u0_L3_1 ) , .D( u0_R2_1 ) );
  DFF_X1 u0_L3_reg_10 (.CK( clk ) , .Q( u0_L3_10 ) , .D( u0_R2_10 ) );
  DFF_X1 u0_L3_reg_11 (.CK( clk ) , .Q( u0_L3_11 ) , .D( u0_R2_11 ) );
  DFF_X1 u0_L3_reg_12 (.CK( clk ) , .Q( u0_L3_12 ) , .D( u0_R2_12 ) );
  DFF_X1 u0_L3_reg_13 (.CK( clk ) , .Q( u0_L3_13 ) , .D( u0_R2_13 ) );
  DFF_X1 u0_L3_reg_14 (.CK( clk ) , .Q( u0_L3_14 ) , .D( u0_R2_14 ) );
  DFF_X1 u0_L3_reg_15 (.CK( clk ) , .Q( u0_L3_15 ) , .D( u0_R2_15 ) );
  DFF_X1 u0_L3_reg_16 (.CK( clk ) , .Q( u0_L3_16 ) , .D( u0_R2_16 ) );
  DFF_X1 u0_L3_reg_17 (.CK( clk ) , .Q( u0_L3_17 ) , .D( u0_R2_17 ) );
  DFF_X1 u0_L3_reg_18 (.CK( clk ) , .Q( u0_L3_18 ) , .D( u0_R2_18 ) );
  DFF_X1 u0_L3_reg_19 (.CK( clk ) , .Q( u0_L3_19 ) , .D( u0_R2_19 ) );
  DFF_X1 u0_L3_reg_2 (.CK( clk ) , .Q( u0_L3_2 ) , .D( u0_R2_2 ) );
  DFF_X1 u0_L3_reg_20 (.CK( clk ) , .Q( u0_L3_20 ) , .D( u0_R2_20 ) );
  DFF_X1 u0_L3_reg_21 (.CK( clk ) , .Q( u0_L3_21 ) , .D( u0_R2_21 ) );
  DFF_X1 u0_L3_reg_22 (.CK( clk ) , .Q( u0_L3_22 ) , .D( u0_R2_22 ) );
  DFF_X1 u0_L3_reg_23 (.CK( clk ) , .Q( u0_L3_23 ) , .D( u0_R2_23 ) );
  DFF_X1 u0_L3_reg_24 (.CK( clk ) , .Q( u0_L3_24 ) , .D( u0_R2_24 ) );
  DFF_X1 u0_L3_reg_25 (.CK( clk ) , .Q( u0_L3_25 ) , .D( u0_R2_25 ) );
  DFF_X1 u0_L3_reg_26 (.CK( clk ) , .Q( u0_L3_26 ) , .D( u0_R2_26 ) );
  DFF_X1 u0_L3_reg_27 (.CK( clk ) , .Q( u0_L3_27 ) , .D( u0_R2_27 ) );
  DFF_X1 u0_L3_reg_28 (.CK( clk ) , .Q( u0_L3_28 ) , .D( u0_R2_28 ) );
  DFF_X1 u0_L3_reg_29 (.CK( clk ) , .Q( u0_L3_29 ) , .D( u0_R2_29 ) );
  DFF_X1 u0_L3_reg_3 (.CK( clk ) , .Q( u0_L3_3 ) , .D( u0_R2_3 ) );
  DFF_X1 u0_L3_reg_30 (.CK( clk ) , .Q( u0_L3_30 ) , .D( u0_R2_30 ) );
  DFF_X1 u0_L3_reg_31 (.CK( clk ) , .Q( u0_L3_31 ) , .D( u0_R2_31 ) );
  DFF_X1 u0_L3_reg_32 (.CK( clk ) , .Q( u0_L3_32 ) , .D( u0_R2_32 ) );
  DFF_X1 u0_L3_reg_4 (.CK( clk ) , .Q( u0_L3_4 ) , .D( u0_R2_4 ) );
  DFF_X1 u0_L3_reg_5 (.CK( clk ) , .Q( u0_L3_5 ) , .D( u0_R2_5 ) );
  DFF_X1 u0_L3_reg_6 (.CK( clk ) , .Q( u0_L3_6 ) , .D( u0_R2_6 ) );
  DFF_X1 u0_L3_reg_7 (.CK( clk ) , .Q( u0_L3_7 ) , .D( u0_R2_7 ) );
  DFF_X1 u0_L3_reg_8 (.CK( clk ) , .Q( u0_L3_8 ) , .D( u0_R2_8 ) );
  DFF_X1 u0_L3_reg_9 (.CK( clk ) , .Q( u0_L3_9 ) , .D( u0_R2_9 ) );
  DFF_X1 u0_L4_reg_1 (.CK( clk ) , .Q( u0_L4_1 ) , .D( u0_R3_1 ) );
  DFF_X1 u0_L4_reg_10 (.CK( clk ) , .Q( u0_L4_10 ) , .D( u0_R3_10 ) );
  DFF_X1 u0_L4_reg_11 (.CK( clk ) , .Q( u0_L4_11 ) , .D( u0_R3_11 ) );
  DFF_X1 u0_L4_reg_12 (.CK( clk ) , .Q( u0_L4_12 ) , .D( u0_R3_12 ) );
  DFF_X1 u0_L4_reg_13 (.CK( clk ) , .Q( u0_L4_13 ) , .D( u0_R3_13 ) );
  DFF_X1 u0_L4_reg_14 (.CK( clk ) , .Q( u0_L4_14 ) , .D( u0_R3_14 ) );
  DFF_X1 u0_L4_reg_15 (.CK( clk ) , .Q( u0_L4_15 ) , .D( u0_R3_15 ) );
  DFF_X1 u0_L4_reg_16 (.CK( clk ) , .Q( u0_L4_16 ) , .D( u0_R3_16 ) );
  DFF_X1 u0_L4_reg_17 (.CK( clk ) , .Q( u0_L4_17 ) , .D( u0_R3_17 ) );
  DFF_X1 u0_L4_reg_18 (.CK( clk ) , .Q( u0_L4_18 ) , .D( u0_R3_18 ) );
  DFF_X1 u0_L4_reg_19 (.CK( clk ) , .Q( u0_L4_19 ) , .D( u0_R3_19 ) );
  DFF_X1 u0_L4_reg_2 (.CK( clk ) , .Q( u0_L4_2 ) , .D( u0_R3_2 ) );
  DFF_X1 u0_L4_reg_20 (.CK( clk ) , .Q( u0_L4_20 ) , .D( u0_R3_20 ) );
  DFF_X1 u0_L4_reg_21 (.CK( clk ) , .Q( u0_L4_21 ) , .D( u0_R3_21 ) );
  DFF_X1 u0_L4_reg_22 (.CK( clk ) , .Q( u0_L4_22 ) , .D( u0_R3_22 ) );
  DFF_X1 u0_L4_reg_23 (.CK( clk ) , .Q( u0_L4_23 ) , .D( u0_R3_23 ) );
  DFF_X1 u0_L4_reg_24 (.CK( clk ) , .Q( u0_L4_24 ) , .D( u0_R3_24 ) );
  DFF_X1 u0_L4_reg_25 (.CK( clk ) , .Q( u0_L4_25 ) , .D( u0_R3_25 ) );
  DFF_X1 u0_L4_reg_26 (.CK( clk ) , .Q( u0_L4_26 ) , .D( u0_R3_26 ) );
  DFF_X1 u0_L4_reg_27 (.CK( clk ) , .Q( u0_L4_27 ) , .D( u0_R3_27 ) );
  DFF_X1 u0_L4_reg_28 (.CK( clk ) , .Q( u0_L4_28 ) , .D( u0_R3_28 ) );
  DFF_X1 u0_L4_reg_29 (.CK( clk ) , .Q( u0_L4_29 ) , .D( u0_R3_29 ) );
  DFF_X1 u0_L4_reg_3 (.CK( clk ) , .Q( u0_L4_3 ) , .D( u0_R3_3 ) );
  DFF_X1 u0_L4_reg_30 (.CK( clk ) , .Q( u0_L4_30 ) , .D( u0_R3_30 ) );
  DFF_X1 u0_L4_reg_31 (.CK( clk ) , .Q( u0_L4_31 ) , .D( u0_R3_31 ) );
  DFF_X1 u0_L4_reg_32 (.CK( clk ) , .Q( u0_L4_32 ) , .D( u0_R3_32 ) );
  DFF_X1 u0_L4_reg_4 (.CK( clk ) , .Q( u0_L4_4 ) , .D( u0_R3_4 ) );
  DFF_X1 u0_L4_reg_5 (.CK( clk ) , .Q( u0_L4_5 ) , .D( u0_R3_5 ) );
  DFF_X1 u0_L4_reg_6 (.CK( clk ) , .Q( u0_L4_6 ) , .D( u0_R3_6 ) );
  DFF_X1 u0_L4_reg_7 (.CK( clk ) , .Q( u0_L4_7 ) , .D( u0_R3_7 ) );
  DFF_X1 u0_L4_reg_8 (.CK( clk ) , .Q( u0_L4_8 ) , .D( u0_R3_8 ) );
  DFF_X1 u0_L4_reg_9 (.CK( clk ) , .Q( u0_L4_9 ) , .D( u0_R3_9 ) );
  DFF_X1 u0_L5_reg_1 (.CK( clk ) , .Q( u0_L5_1 ) , .D( u0_R4_1 ) );
  DFF_X1 u0_L5_reg_10 (.CK( clk ) , .Q( u0_L5_10 ) , .D( u0_R4_10 ) );
  DFF_X1 u0_L5_reg_11 (.CK( clk ) , .Q( u0_L5_11 ) , .D( u0_R4_11 ) );
  DFF_X1 u0_L5_reg_12 (.CK( clk ) , .Q( u0_L5_12 ) , .D( u0_R4_12 ) );
  DFF_X1 u0_L5_reg_13 (.CK( clk ) , .Q( u0_L5_13 ) , .D( u0_R4_13 ) );
  DFF_X1 u0_L5_reg_14 (.CK( clk ) , .Q( u0_L5_14 ) , .D( u0_R4_14 ) );
  DFF_X1 u0_L5_reg_15 (.CK( clk ) , .Q( u0_L5_15 ) , .D( u0_R4_15 ) );
  DFF_X1 u0_L5_reg_16 (.CK( clk ) , .Q( u0_L5_16 ) , .D( u0_R4_16 ) );
  DFF_X1 u0_L5_reg_17 (.CK( clk ) , .Q( u0_L5_17 ) , .D( u0_R4_17 ) );
  DFF_X1 u0_L5_reg_18 (.CK( clk ) , .Q( u0_L5_18 ) , .D( u0_R4_18 ) );
  DFF_X1 u0_L5_reg_19 (.CK( clk ) , .Q( u0_L5_19 ) , .D( u0_R4_19 ) );
  DFF_X1 u0_L5_reg_2 (.CK( clk ) , .Q( u0_L5_2 ) , .D( u0_R4_2 ) );
  DFF_X1 u0_L5_reg_20 (.CK( clk ) , .Q( u0_L5_20 ) , .D( u0_R4_20 ) );
  DFF_X1 u0_L5_reg_21 (.CK( clk ) , .Q( u0_L5_21 ) , .D( u0_R4_21 ) );
  DFF_X1 u0_L5_reg_22 (.CK( clk ) , .Q( u0_L5_22 ) , .D( u0_R4_22 ) );
  DFF_X1 u0_L5_reg_23 (.CK( clk ) , .Q( u0_L5_23 ) , .D( u0_R4_23 ) );
  DFF_X1 u0_L5_reg_24 (.CK( clk ) , .Q( u0_L5_24 ) , .D( u0_R4_24 ) );
  DFF_X1 u0_L5_reg_25 (.CK( clk ) , .Q( u0_L5_25 ) , .D( u0_R4_25 ) );
  DFF_X1 u0_L5_reg_26 (.CK( clk ) , .Q( u0_L5_26 ) , .D( u0_R4_26 ) );
  DFF_X1 u0_L5_reg_27 (.CK( clk ) , .Q( u0_L5_27 ) , .D( u0_R4_27 ) );
  DFF_X1 u0_L5_reg_28 (.CK( clk ) , .Q( u0_L5_28 ) , .D( u0_R4_28 ) );
  DFF_X1 u0_L5_reg_29 (.CK( clk ) , .Q( u0_L5_29 ) , .D( u0_R4_29 ) );
  DFF_X1 u0_L5_reg_3 (.CK( clk ) , .Q( u0_L5_3 ) , .D( u0_R4_3 ) );
  DFF_X1 u0_L5_reg_30 (.CK( clk ) , .Q( u0_L5_30 ) , .D( u0_R4_30 ) );
  DFF_X1 u0_L5_reg_31 (.CK( clk ) , .Q( u0_L5_31 ) , .D( u0_R4_31 ) );
  DFF_X1 u0_L5_reg_32 (.CK( clk ) , .Q( u0_L5_32 ) , .D( u0_R4_32 ) );
  DFF_X1 u0_L5_reg_4 (.CK( clk ) , .Q( u0_L5_4 ) , .D( u0_R4_4 ) );
  DFF_X1 u0_L5_reg_5 (.CK( clk ) , .Q( u0_L5_5 ) , .D( u0_R4_5 ) );
  DFF_X1 u0_L5_reg_6 (.CK( clk ) , .Q( u0_L5_6 ) , .D( u0_R4_6 ) );
  DFF_X1 u0_L5_reg_7 (.CK( clk ) , .Q( u0_L5_7 ) , .D( u0_R4_7 ) );
  DFF_X1 u0_L5_reg_8 (.CK( clk ) , .Q( u0_L5_8 ) , .D( u0_R4_8 ) );
  DFF_X1 u0_L5_reg_9 (.CK( clk ) , .Q( u0_L5_9 ) , .D( u0_R4_9 ) );
  DFF_X1 u0_L6_reg_1 (.CK( clk ) , .Q( u0_L6_1 ) , .D( u0_R5_1 ) );
  DFF_X1 u0_L6_reg_10 (.CK( clk ) , .Q( u0_L6_10 ) , .D( u0_R5_10 ) );
  DFF_X1 u0_L6_reg_11 (.CK( clk ) , .Q( u0_L6_11 ) , .D( u0_R5_11 ) );
  DFF_X1 u0_L6_reg_12 (.CK( clk ) , .Q( u0_L6_12 ) , .D( u0_R5_12 ) );
  DFF_X1 u0_L6_reg_13 (.CK( clk ) , .Q( u0_L6_13 ) , .D( u0_R5_13 ) );
  DFF_X1 u0_L6_reg_14 (.CK( clk ) , .Q( u0_L6_14 ) , .D( u0_R5_14 ) );
  DFF_X1 u0_L6_reg_15 (.CK( clk ) , .Q( u0_L6_15 ) , .D( u0_R5_15 ) );
  DFF_X1 u0_L6_reg_16 (.CK( clk ) , .Q( u0_L6_16 ) , .D( u0_R5_16 ) );
  DFF_X1 u0_L6_reg_17 (.CK( clk ) , .Q( u0_L6_17 ) , .D( u0_R5_17 ) );
  DFF_X1 u0_L6_reg_18 (.CK( clk ) , .Q( u0_L6_18 ) , .D( u0_R5_18 ) );
  DFF_X1 u0_L6_reg_19 (.CK( clk ) , .Q( u0_L6_19 ) , .D( u0_R5_19 ) );
  DFF_X1 u0_L6_reg_2 (.CK( clk ) , .Q( u0_L6_2 ) , .D( u0_R5_2 ) );
  DFF_X1 u0_L6_reg_20 (.CK( clk ) , .Q( u0_L6_20 ) , .D( u0_R5_20 ) );
  DFF_X1 u0_L6_reg_21 (.CK( clk ) , .Q( u0_L6_21 ) , .D( u0_R5_21 ) );
  DFF_X1 u0_L6_reg_22 (.CK( clk ) , .Q( u0_L6_22 ) , .D( u0_R5_22 ) );
  DFF_X1 u0_L6_reg_23 (.CK( clk ) , .Q( u0_L6_23 ) , .D( u0_R5_23 ) );
  DFF_X1 u0_L6_reg_24 (.CK( clk ) , .Q( u0_L6_24 ) , .D( u0_R5_24 ) );
  DFF_X1 u0_L6_reg_25 (.CK( clk ) , .Q( u0_L6_25 ) , .D( u0_R5_25 ) );
  DFF_X1 u0_L6_reg_26 (.CK( clk ) , .Q( u0_L6_26 ) , .D( u0_R5_26 ) );
  DFF_X1 u0_L6_reg_27 (.CK( clk ) , .Q( u0_L6_27 ) , .D( u0_R5_27 ) );
  DFF_X1 u0_L6_reg_28 (.CK( clk ) , .Q( u0_L6_28 ) , .D( u0_R5_28 ) );
  DFF_X1 u0_L6_reg_29 (.CK( clk ) , .Q( u0_L6_29 ) , .D( u0_R5_29 ) );
  DFF_X1 u0_L6_reg_3 (.CK( clk ) , .Q( u0_L6_3 ) , .D( u0_R5_3 ) );
  DFF_X1 u0_L6_reg_30 (.CK( clk ) , .Q( u0_L6_30 ) , .D( u0_R5_30 ) );
  DFF_X1 u0_L6_reg_31 (.CK( clk ) , .Q( u0_L6_31 ) , .D( u0_R5_31 ) );
  DFF_X1 u0_L6_reg_32 (.CK( clk ) , .Q( u0_L6_32 ) , .D( u0_R5_32 ) );
  DFF_X1 u0_L6_reg_4 (.CK( clk ) , .Q( u0_L6_4 ) , .D( u0_R5_4 ) );
  DFF_X1 u0_L6_reg_5 (.CK( clk ) , .Q( u0_L6_5 ) , .D( u0_R5_5 ) );
  DFF_X1 u0_L6_reg_6 (.CK( clk ) , .Q( u0_L6_6 ) , .D( u0_R5_6 ) );
  DFF_X1 u0_L6_reg_7 (.CK( clk ) , .Q( u0_L6_7 ) , .D( u0_R5_7 ) );
  DFF_X1 u0_L6_reg_8 (.CK( clk ) , .Q( u0_L6_8 ) , .D( u0_R5_8 ) );
  DFF_X1 u0_L6_reg_9 (.CK( clk ) , .Q( u0_L6_9 ) , .D( u0_R5_9 ) );
  DFF_X1 u0_L7_reg_1 (.CK( clk ) , .Q( u0_L7_1 ) , .D( u0_R6_1 ) );
  DFF_X1 u0_L7_reg_10 (.CK( clk ) , .Q( u0_L7_10 ) , .D( u0_R6_10 ) );
  DFF_X1 u0_L7_reg_11 (.CK( clk ) , .Q( u0_L7_11 ) , .D( u0_R6_11 ) );
  DFF_X1 u0_L7_reg_12 (.CK( clk ) , .Q( u0_L7_12 ) , .D( u0_R6_12 ) );
  DFF_X1 u0_L7_reg_13 (.CK( clk ) , .Q( u0_L7_13 ) , .D( u0_R6_13 ) );
  DFF_X1 u0_L7_reg_14 (.CK( clk ) , .Q( u0_L7_14 ) , .D( u0_R6_14 ) );
  DFF_X1 u0_L7_reg_15 (.CK( clk ) , .Q( u0_L7_15 ) , .D( u0_R6_15 ) );
  DFF_X1 u0_L7_reg_16 (.CK( clk ) , .Q( u0_L7_16 ) , .D( u0_R6_16 ) );
  DFF_X1 u0_L7_reg_17 (.CK( clk ) , .Q( u0_L7_17 ) , .D( u0_R6_17 ) );
  DFF_X1 u0_L7_reg_18 (.CK( clk ) , .Q( u0_L7_18 ) , .D( u0_R6_18 ) );
  DFF_X1 u0_L7_reg_19 (.CK( clk ) , .Q( u0_L7_19 ) , .D( u0_R6_19 ) );
  DFF_X1 u0_L7_reg_2 (.CK( clk ) , .Q( u0_L7_2 ) , .D( u0_R6_2 ) );
  DFF_X1 u0_L7_reg_20 (.CK( clk ) , .Q( u0_L7_20 ) , .D( u0_R6_20 ) );
  DFF_X1 u0_L7_reg_21 (.CK( clk ) , .Q( u0_L7_21 ) , .D( u0_R6_21 ) );
  DFF_X1 u0_L7_reg_22 (.CK( clk ) , .Q( u0_L7_22 ) , .D( u0_R6_22 ) );
  DFF_X1 u0_L7_reg_23 (.CK( clk ) , .Q( u0_L7_23 ) , .D( u0_R6_23 ) );
  DFF_X1 u0_L7_reg_24 (.CK( clk ) , .Q( u0_L7_24 ) , .D( u0_R6_24 ) );
  DFF_X1 u0_L7_reg_25 (.CK( clk ) , .Q( u0_L7_25 ) , .D( u0_R6_25 ) );
  DFF_X1 u0_L7_reg_26 (.CK( clk ) , .Q( u0_L7_26 ) , .D( u0_R6_26 ) );
  DFF_X1 u0_L7_reg_27 (.CK( clk ) , .Q( u0_L7_27 ) , .D( u0_R6_27 ) );
  DFF_X1 u0_L7_reg_28 (.CK( clk ) , .Q( u0_L7_28 ) , .D( u0_R6_28 ) );
  DFF_X1 u0_L7_reg_29 (.CK( clk ) , .Q( u0_L7_29 ) , .D( u0_R6_29 ) );
  DFF_X1 u0_L7_reg_3 (.CK( clk ) , .Q( u0_L7_3 ) , .D( u0_R6_3 ) );
  DFF_X1 u0_L7_reg_30 (.CK( clk ) , .Q( u0_L7_30 ) , .D( u0_R6_30 ) );
  DFF_X1 u0_L7_reg_31 (.CK( clk ) , .Q( u0_L7_31 ) , .D( u0_R6_31 ) );
  DFF_X1 u0_L7_reg_32 (.CK( clk ) , .Q( u0_L7_32 ) , .D( u0_R6_32 ) );
  DFF_X1 u0_L7_reg_4 (.CK( clk ) , .Q( u0_L7_4 ) , .D( u0_R6_4 ) );
  DFF_X1 u0_L7_reg_5 (.CK( clk ) , .Q( u0_L7_5 ) , .D( u0_R6_5 ) );
  DFF_X1 u0_L7_reg_6 (.CK( clk ) , .Q( u0_L7_6 ) , .D( u0_R6_6 ) );
  DFF_X1 u0_L7_reg_7 (.CK( clk ) , .Q( u0_L7_7 ) , .D( u0_R6_7 ) );
  DFF_X1 u0_L7_reg_8 (.CK( clk ) , .Q( u0_L7_8 ) , .D( u0_R6_8 ) );
  DFF_X1 u0_L7_reg_9 (.CK( clk ) , .Q( u0_L7_9 ) , .D( u0_R6_9 ) );
  DFF_X1 u0_L8_reg_1 (.CK( clk ) , .Q( u0_L8_1 ) , .D( u0_R7_1 ) );
  DFF_X1 u0_L8_reg_10 (.CK( clk ) , .Q( u0_L8_10 ) , .D( u0_R7_10 ) );
  DFF_X1 u0_L8_reg_11 (.CK( clk ) , .Q( u0_L8_11 ) , .D( u0_R7_11 ) );
  DFF_X1 u0_L8_reg_12 (.CK( clk ) , .Q( u0_L8_12 ) , .D( u0_R7_12 ) );
  DFF_X1 u0_L8_reg_13 (.CK( clk ) , .Q( u0_L8_13 ) , .D( u0_R7_13 ) );
  DFF_X1 u0_L8_reg_14 (.CK( clk ) , .Q( u0_L8_14 ) , .D( u0_R7_14 ) );
  DFF_X1 u0_L8_reg_15 (.CK( clk ) , .Q( u0_L8_15 ) , .D( u0_R7_15 ) );
  DFF_X1 u0_L8_reg_16 (.CK( clk ) , .Q( u0_L8_16 ) , .D( u0_R7_16 ) );
  DFF_X1 u0_L8_reg_17 (.CK( clk ) , .Q( u0_L8_17 ) , .D( u0_R7_17 ) );
  DFF_X1 u0_L8_reg_18 (.CK( clk ) , .Q( u0_L8_18 ) , .D( u0_R7_18 ) );
  DFF_X1 u0_L8_reg_19 (.CK( clk ) , .Q( u0_L8_19 ) , .D( u0_R7_19 ) );
  DFF_X1 u0_L8_reg_2 (.CK( clk ) , .Q( u0_L8_2 ) , .D( u0_R7_2 ) );
  DFF_X1 u0_L8_reg_20 (.CK( clk ) , .Q( u0_L8_20 ) , .D( u0_R7_20 ) );
  DFF_X1 u0_L8_reg_21 (.CK( clk ) , .Q( u0_L8_21 ) , .D( u0_R7_21 ) );
  DFF_X1 u0_L8_reg_22 (.CK( clk ) , .Q( u0_L8_22 ) , .D( u0_R7_22 ) );
  DFF_X1 u0_L8_reg_23 (.CK( clk ) , .Q( u0_L8_23 ) , .D( u0_R7_23 ) );
  DFF_X1 u0_L8_reg_24 (.CK( clk ) , .Q( u0_L8_24 ) , .D( u0_R7_24 ) );
  DFF_X1 u0_L8_reg_25 (.CK( clk ) , .Q( u0_L8_25 ) , .D( u0_R7_25 ) );
  DFF_X1 u0_L8_reg_26 (.CK( clk ) , .Q( u0_L8_26 ) , .D( u0_R7_26 ) );
  DFF_X1 u0_L8_reg_27 (.CK( clk ) , .Q( u0_L8_27 ) , .D( u0_R7_27 ) );
  DFF_X1 u0_L8_reg_28 (.CK( clk ) , .Q( u0_L8_28 ) , .D( u0_R7_28 ) );
  DFF_X1 u0_L8_reg_29 (.CK( clk ) , .Q( u0_L8_29 ) , .D( u0_R7_29 ) );
  DFF_X1 u0_L8_reg_3 (.CK( clk ) , .Q( u0_L8_3 ) , .D( u0_R7_3 ) );
  DFF_X1 u0_L8_reg_30 (.CK( clk ) , .Q( u0_L8_30 ) , .D( u0_R7_30 ) );
  DFF_X1 u0_L8_reg_31 (.CK( clk ) , .Q( u0_L8_31 ) , .D( u0_R7_31 ) );
  DFF_X1 u0_L8_reg_32 (.CK( clk ) , .Q( u0_L8_32 ) , .D( u0_R7_32 ) );
  DFF_X1 u0_L8_reg_4 (.CK( clk ) , .Q( u0_L8_4 ) , .D( u0_R7_4 ) );
  DFF_X1 u0_L8_reg_5 (.CK( clk ) , .Q( u0_L8_5 ) , .D( u0_R7_5 ) );
  DFF_X1 u0_L8_reg_6 (.CK( clk ) , .Q( u0_L8_6 ) , .D( u0_R7_6 ) );
  DFF_X1 u0_L8_reg_7 (.CK( clk ) , .Q( u0_L8_7 ) , .D( u0_R7_7 ) );
  DFF_X1 u0_L8_reg_8 (.CK( clk ) , .Q( u0_L8_8 ) , .D( u0_R7_8 ) );
  DFF_X1 u0_L8_reg_9 (.CK( clk ) , .Q( u0_L8_9 ) , .D( u0_R7_9 ) );
  DFF_X1 u0_L9_reg_1 (.CK( clk ) , .Q( u0_L9_1 ) , .D( u0_R8_1 ) );
  DFF_X1 u0_L9_reg_10 (.CK( clk ) , .Q( u0_L9_10 ) , .D( u0_R8_10 ) );
  DFF_X1 u0_L9_reg_11 (.CK( clk ) , .Q( u0_L9_11 ) , .D( u0_R8_11 ) );
  DFF_X1 u0_L9_reg_12 (.CK( clk ) , .Q( u0_L9_12 ) , .D( u0_R8_12 ) );
  DFF_X1 u0_L9_reg_13 (.CK( clk ) , .Q( u0_L9_13 ) , .D( u0_R8_13 ) );
  DFF_X1 u0_L9_reg_14 (.CK( clk ) , .Q( u0_L9_14 ) , .D( u0_R8_14 ) );
  DFF_X1 u0_L9_reg_15 (.CK( clk ) , .Q( u0_L9_15 ) , .D( u0_R8_15 ) );
  DFF_X1 u0_L9_reg_16 (.CK( clk ) , .Q( u0_L9_16 ) , .D( u0_R8_16 ) );
  DFF_X1 u0_L9_reg_17 (.CK( clk ) , .Q( u0_L9_17 ) , .D( u0_R8_17 ) );
  DFF_X1 u0_L9_reg_18 (.CK( clk ) , .Q( u0_L9_18 ) , .D( u0_R8_18 ) );
  DFF_X1 u0_L9_reg_19 (.CK( clk ) , .Q( u0_L9_19 ) , .D( u0_R8_19 ) );
  DFF_X1 u0_L9_reg_2 (.CK( clk ) , .Q( u0_L9_2 ) , .D( u0_R8_2 ) );
  DFF_X1 u0_L9_reg_20 (.CK( clk ) , .Q( u0_L9_20 ) , .D( u0_R8_20 ) );
  DFF_X1 u0_L9_reg_21 (.CK( clk ) , .Q( u0_L9_21 ) , .D( u0_R8_21 ) );
  DFF_X1 u0_L9_reg_22 (.CK( clk ) , .Q( u0_L9_22 ) , .D( u0_R8_22 ) );
  DFF_X1 u0_L9_reg_23 (.CK( clk ) , .Q( u0_L9_23 ) , .D( u0_R8_23 ) );
  DFF_X1 u0_L9_reg_24 (.CK( clk ) , .Q( u0_L9_24 ) , .D( u0_R8_24 ) );
  DFF_X1 u0_L9_reg_25 (.CK( clk ) , .Q( u0_L9_25 ) , .D( u0_R8_25 ) );
  DFF_X1 u0_L9_reg_26 (.CK( clk ) , .Q( u0_L9_26 ) , .D( u0_R8_26 ) );
  DFF_X1 u0_L9_reg_27 (.CK( clk ) , .Q( u0_L9_27 ) , .D( u0_R8_27 ) );
  DFF_X1 u0_L9_reg_28 (.CK( clk ) , .Q( u0_L9_28 ) , .D( u0_R8_28 ) );
  DFF_X1 u0_L9_reg_29 (.CK( clk ) , .Q( u0_L9_29 ) , .D( u0_R8_29 ) );
  DFF_X1 u0_L9_reg_3 (.CK( clk ) , .Q( u0_L9_3 ) , .D( u0_R8_3 ) );
  DFF_X1 u0_L9_reg_30 (.CK( clk ) , .Q( u0_L9_30 ) , .D( u0_R8_30 ) );
  DFF_X1 u0_L9_reg_31 (.CK( clk ) , .Q( u0_L9_31 ) , .D( u0_R8_31 ) );
  DFF_X1 u0_L9_reg_32 (.CK( clk ) , .Q( u0_L9_32 ) , .D( u0_R8_32 ) );
  DFF_X1 u0_L9_reg_4 (.CK( clk ) , .Q( u0_L9_4 ) , .D( u0_R8_4 ) );
  DFF_X1 u0_L9_reg_5 (.CK( clk ) , .Q( u0_L9_5 ) , .D( u0_R8_5 ) );
  DFF_X1 u0_L9_reg_6 (.CK( clk ) , .Q( u0_L9_6 ) , .D( u0_R8_6 ) );
  DFF_X1 u0_L9_reg_7 (.CK( clk ) , .Q( u0_L9_7 ) , .D( u0_R8_7 ) );
  DFF_X1 u0_L9_reg_8 (.CK( clk ) , .Q( u0_L9_8 ) , .D( u0_R8_8 ) );
  DFF_X1 u0_L9_reg_9 (.CK( clk ) , .Q( u0_L9_9 ) , .D( u0_R8_9 ) );
  DFF_X1 u0_R0_reg_1 (.CK( clk ) , .D( u0_N0 ) , .Q( u0_R0_1 ) );
  DFF_X1 u0_R0_reg_10 (.CK( clk ) , .D( u0_N9 ) , .Q( u0_R0_10 ) );
  DFF_X1 u0_R0_reg_11 (.CK( clk ) , .D( u0_N10 ) , .Q( u0_R0_11 ) );
  DFF_X1 u0_R0_reg_12 (.CK( clk ) , .D( u0_N11 ) , .Q( u0_R0_12 ) );
  DFF_X1 u0_R0_reg_13 (.CK( clk ) , .D( u0_N12 ) , .Q( u0_R0_13 ) );
  DFF_X1 u0_R0_reg_14 (.CK( clk ) , .D( u0_N13 ) , .Q( u0_R0_14 ) );
  DFF_X1 u0_R0_reg_15 (.CK( clk ) , .D( u0_N14 ) , .Q( u0_R0_15 ) );
  DFF_X1 u0_R0_reg_16 (.CK( clk ) , .D( u0_N15 ) , .Q( u0_R0_16 ) );
  DFF_X1 u0_R0_reg_17 (.CK( clk ) , .D( u0_N16 ) , .Q( u0_R0_17 ) );
  DFF_X1 u0_R0_reg_18 (.CK( clk ) , .D( u0_N17 ) , .Q( u0_R0_18 ) );
  DFF_X1 u0_R0_reg_19 (.CK( clk ) , .D( u0_N18 ) , .Q( u0_R0_19 ) );
  DFF_X1 u0_R0_reg_2 (.CK( clk ) , .D( u0_N1 ) , .Q( u0_R0_2 ) );
  DFF_X1 u0_R0_reg_20 (.CK( clk ) , .D( u0_N19 ) , .Q( u0_R0_20 ) );
  DFF_X1 u0_R0_reg_21 (.CK( clk ) , .D( u0_N20 ) , .Q( u0_R0_21 ) );
  DFF_X1 u0_R0_reg_22 (.CK( clk ) , .D( u0_N21 ) , .Q( u0_R0_22 ) );
  DFF_X1 u0_R0_reg_23 (.CK( clk ) , .D( u0_N22 ) , .Q( u0_R0_23 ) );
  DFF_X1 u0_R0_reg_24 (.CK( clk ) , .D( u0_N23 ) , .Q( u0_R0_24 ) );
  DFF_X1 u0_R0_reg_25 (.CK( clk ) , .D( u0_N24 ) , .Q( u0_R0_25 ) );
  DFF_X1 u0_R0_reg_26 (.CK( clk ) , .D( u0_N25 ) , .Q( u0_R0_26 ) );
  DFF_X1 u0_R0_reg_27 (.CK( clk ) , .D( u0_N26 ) , .Q( u0_R0_27 ) );
  DFF_X1 u0_R0_reg_28 (.CK( clk ) , .D( u0_N27 ) , .Q( u0_R0_28 ) );
  DFF_X1 u0_R0_reg_29 (.CK( clk ) , .D( u0_N28 ) , .Q( u0_R0_29 ) );
  DFF_X1 u0_R0_reg_3 (.CK( clk ) , .D( u0_N2 ) , .Q( u0_R0_3 ) );
  DFF_X1 u0_R0_reg_30 (.CK( clk ) , .D( u0_N29 ) , .Q( u0_R0_30 ) );
  DFF_X1 u0_R0_reg_31 (.CK( clk ) , .D( u0_N30 ) , .Q( u0_R0_31 ) );
  DFF_X1 u0_R0_reg_32 (.CK( clk ) , .D( u0_N31 ) , .Q( u0_R0_32 ) );
  DFF_X1 u0_R0_reg_4 (.CK( clk ) , .D( u0_N3 ) , .Q( u0_R0_4 ) );
  DFF_X1 u0_R0_reg_5 (.CK( clk ) , .D( u0_N4 ) , .Q( u0_R0_5 ) );
  DFF_X1 u0_R0_reg_6 (.CK( clk ) , .D( u0_N5 ) , .Q( u0_R0_6 ) );
  DFF_X1 u0_R0_reg_7 (.CK( clk ) , .D( u0_N6 ) , .Q( u0_R0_7 ) );
  DFF_X1 u0_R0_reg_8 (.CK( clk ) , .D( u0_N7 ) , .Q( u0_R0_8 ) );
  DFF_X1 u0_R0_reg_9 (.CK( clk ) , .D( u0_N8 ) , .Q( u0_R0_9 ) );
  DFF_X1 u0_R10_reg_1 (.CK( clk ) , .D( u0_N320 ) , .Q( u0_R10_1 ) );
  DFF_X1 u0_R10_reg_10 (.CK( clk ) , .D( u0_N329 ) , .Q( u0_R10_10 ) );
  DFF_X1 u0_R10_reg_11 (.CK( clk ) , .D( u0_N330 ) , .Q( u0_R10_11 ) );
  DFF_X1 u0_R10_reg_12 (.CK( clk ) , .D( u0_N331 ) , .Q( u0_R10_12 ) );
  DFF_X1 u0_R10_reg_13 (.CK( clk ) , .D( u0_N332 ) , .Q( u0_R10_13 ) );
  DFF_X1 u0_R10_reg_14 (.CK( clk ) , .D( u0_N333 ) , .Q( u0_R10_14 ) );
  DFF_X1 u0_R10_reg_15 (.CK( clk ) , .D( u0_N334 ) , .Q( u0_R10_15 ) );
  DFF_X1 u0_R10_reg_16 (.CK( clk ) , .D( u0_N335 ) , .Q( u0_R10_16 ) );
  DFF_X1 u0_R10_reg_17 (.CK( clk ) , .D( u0_N336 ) , .Q( u0_R10_17 ) );
  DFF_X1 u0_R10_reg_18 (.CK( clk ) , .D( u0_N337 ) , .Q( u0_R10_18 ) );
  DFF_X1 u0_R10_reg_19 (.CK( clk ) , .D( u0_N338 ) , .Q( u0_R10_19 ) );
  DFF_X1 u0_R10_reg_2 (.CK( clk ) , .D( u0_N321 ) , .Q( u0_R10_2 ) );
  DFF_X1 u0_R10_reg_20 (.CK( clk ) , .D( u0_N339 ) , .Q( u0_R10_20 ) );
  DFF_X1 u0_R10_reg_21 (.CK( clk ) , .D( u0_N340 ) , .Q( u0_R10_21 ) );
  DFF_X1 u0_R10_reg_22 (.CK( clk ) , .D( u0_N341 ) , .Q( u0_R10_22 ) );
  DFF_X1 u0_R10_reg_23 (.CK( clk ) , .D( u0_N342 ) , .Q( u0_R10_23 ) );
  DFF_X1 u0_R10_reg_24 (.CK( clk ) , .D( u0_N343 ) , .Q( u0_R10_24 ) );
  DFF_X1 u0_R10_reg_25 (.CK( clk ) , .D( u0_N344 ) , .Q( u0_R10_25 ) );
  DFF_X1 u0_R10_reg_26 (.CK( clk ) , .D( u0_N345 ) , .Q( u0_R10_26 ) );
  DFF_X1 u0_R10_reg_27 (.CK( clk ) , .D( u0_N346 ) , .Q( u0_R10_27 ) );
  DFF_X1 u0_R10_reg_28 (.CK( clk ) , .D( u0_N347 ) , .Q( u0_R10_28 ) );
  DFF_X1 u0_R10_reg_29 (.CK( clk ) , .D( u0_N348 ) , .Q( u0_R10_29 ) );
  DFF_X1 u0_R10_reg_3 (.CK( clk ) , .D( u0_N322 ) , .Q( u0_R10_3 ) );
  DFF_X1 u0_R10_reg_30 (.CK( clk ) , .D( u0_N349 ) , .Q( u0_R10_30 ) );
  DFF_X1 u0_R10_reg_31 (.CK( clk ) , .D( u0_N350 ) , .Q( u0_R10_31 ) );
  DFF_X1 u0_R10_reg_32 (.CK( clk ) , .D( u0_N351 ) , .Q( u0_R10_32 ) );
  DFF_X1 u0_R10_reg_4 (.CK( clk ) , .D( u0_N323 ) , .Q( u0_R10_4 ) );
  DFF_X1 u0_R10_reg_5 (.CK( clk ) , .D( u0_N324 ) , .Q( u0_R10_5 ) );
  DFF_X1 u0_R10_reg_6 (.CK( clk ) , .D( u0_N325 ) , .Q( u0_R10_6 ) );
  DFF_X1 u0_R10_reg_7 (.CK( clk ) , .D( u0_N326 ) , .Q( u0_R10_7 ) );
  DFF_X1 u0_R10_reg_8 (.CK( clk ) , .D( u0_N327 ) , .Q( u0_R10_8 ) );
  DFF_X1 u0_R10_reg_9 (.CK( clk ) , .D( u0_N328 ) , .Q( u0_R10_9 ) );
  DFF_X1 u0_R11_reg_1 (.CK( clk ) , .D( u0_N352 ) , .Q( u0_R11_1 ) );
  DFF_X1 u0_R11_reg_10 (.CK( clk ) , .D( u0_N361 ) , .Q( u0_R11_10 ) );
  DFF_X1 u0_R11_reg_11 (.CK( clk ) , .D( u0_N362 ) , .Q( u0_R11_11 ) );
  DFF_X1 u0_R11_reg_12 (.CK( clk ) , .D( u0_N363 ) , .Q( u0_R11_12 ) );
  DFF_X1 u0_R11_reg_13 (.CK( clk ) , .D( u0_N364 ) , .Q( u0_R11_13 ) );
  DFF_X1 u0_R11_reg_14 (.CK( clk ) , .D( u0_N365 ) , .Q( u0_R11_14 ) );
  DFF_X1 u0_R11_reg_15 (.CK( clk ) , .D( u0_N366 ) , .Q( u0_R11_15 ) );
  DFF_X1 u0_R11_reg_16 (.CK( clk ) , .D( u0_N367 ) , .Q( u0_R11_16 ) );
  DFF_X1 u0_R11_reg_17 (.CK( clk ) , .D( u0_N368 ) , .Q( u0_R11_17 ) );
  DFF_X1 u0_R11_reg_18 (.CK( clk ) , .D( u0_N369 ) , .Q( u0_R11_18 ) );
  DFF_X1 u0_R11_reg_19 (.CK( clk ) , .D( u0_N370 ) , .Q( u0_R11_19 ) );
  DFF_X1 u0_R11_reg_2 (.CK( clk ) , .D( u0_N353 ) , .Q( u0_R11_2 ) );
  DFF_X1 u0_R11_reg_20 (.CK( clk ) , .D( u0_N371 ) , .Q( u0_R11_20 ) );
  DFF_X1 u0_R11_reg_21 (.CK( clk ) , .D( u0_N372 ) , .Q( u0_R11_21 ) );
  DFF_X1 u0_R11_reg_22 (.CK( clk ) , .D( u0_N373 ) , .Q( u0_R11_22 ) );
  DFF_X1 u0_R11_reg_23 (.CK( clk ) , .D( u0_N374 ) , .Q( u0_R11_23 ) );
  DFF_X1 u0_R11_reg_24 (.CK( clk ) , .D( u0_N375 ) , .Q( u0_R11_24 ) );
  DFF_X1 u0_R11_reg_25 (.CK( clk ) , .D( u0_N376 ) , .Q( u0_R11_25 ) );
  DFF_X1 u0_R11_reg_26 (.CK( clk ) , .D( u0_N377 ) , .Q( u0_R11_26 ) );
  DFF_X1 u0_R11_reg_27 (.CK( clk ) , .D( u0_N378 ) , .Q( u0_R11_27 ) );
  DFF_X1 u0_R11_reg_28 (.CK( clk ) , .D( u0_N379 ) , .Q( u0_R11_28 ) );
  DFF_X1 u0_R11_reg_29 (.CK( clk ) , .D( u0_N380 ) , .Q( u0_R11_29 ) );
  DFF_X1 u0_R11_reg_3 (.CK( clk ) , .D( u0_N354 ) , .Q( u0_R11_3 ) );
  DFF_X1 u0_R11_reg_30 (.CK( clk ) , .D( u0_N381 ) , .Q( u0_R11_30 ) );
  DFF_X1 u0_R11_reg_31 (.CK( clk ) , .D( u0_N382 ) , .Q( u0_R11_31 ) );
  DFF_X1 u0_R11_reg_32 (.CK( clk ) , .D( u0_N383 ) , .Q( u0_R11_32 ) );
  DFF_X1 u0_R11_reg_4 (.CK( clk ) , .D( u0_N355 ) , .Q( u0_R11_4 ) );
  DFF_X1 u0_R11_reg_5 (.CK( clk ) , .D( u0_N356 ) , .Q( u0_R11_5 ) );
  DFF_X1 u0_R11_reg_6 (.CK( clk ) , .D( u0_N357 ) , .Q( u0_R11_6 ) );
  DFF_X1 u0_R11_reg_7 (.CK( clk ) , .D( u0_N358 ) , .Q( u0_R11_7 ) );
  DFF_X1 u0_R11_reg_8 (.CK( clk ) , .D( u0_N359 ) , .Q( u0_R11_8 ) );
  DFF_X1 u0_R11_reg_9 (.CK( clk ) , .D( u0_N360 ) , .Q( u0_R11_9 ) );
  DFF_X1 u0_R12_reg_1 (.CK( clk ) , .D( u0_N384 ) , .Q( u0_R12_1 ) );
  DFF_X1 u0_R12_reg_10 (.CK( clk ) , .D( u0_N393 ) , .Q( u0_R12_10 ) );
  DFF_X1 u0_R12_reg_11 (.CK( clk ) , .D( u0_N394 ) , .Q( u0_R12_11 ) );
  DFF_X1 u0_R12_reg_12 (.CK( clk ) , .D( u0_N395 ) , .Q( u0_R12_12 ) );
  DFF_X1 u0_R12_reg_13 (.CK( clk ) , .D( u0_N396 ) , .Q( u0_R12_13 ) );
  DFF_X1 u0_R12_reg_14 (.CK( clk ) , .D( u0_N397 ) , .Q( u0_R12_14 ) );
  DFF_X1 u0_R12_reg_15 (.CK( clk ) , .D( u0_N398 ) , .Q( u0_R12_15 ) );
  DFF_X1 u0_R12_reg_16 (.CK( clk ) , .D( u0_N399 ) , .Q( u0_R12_16 ) );
  DFF_X1 u0_R12_reg_17 (.CK( clk ) , .D( u0_N400 ) , .Q( u0_R12_17 ) );
  DFF_X1 u0_R12_reg_18 (.CK( clk ) , .D( u0_N401 ) , .Q( u0_R12_18 ) );
  DFF_X1 u0_R12_reg_19 (.CK( clk ) , .D( u0_N402 ) , .Q( u0_R12_19 ) );
  DFF_X1 u0_R12_reg_2 (.CK( clk ) , .D( u0_N385 ) , .Q( u0_R12_2 ) );
  DFF_X1 u0_R12_reg_20 (.CK( clk ) , .D( u0_N403 ) , .Q( u0_R12_20 ) );
  DFF_X1 u0_R12_reg_21 (.CK( clk ) , .D( u0_N404 ) , .Q( u0_R12_21 ) );
  DFF_X1 u0_R12_reg_22 (.CK( clk ) , .D( u0_N405 ) , .Q( u0_R12_22 ) );
  DFF_X1 u0_R12_reg_23 (.CK( clk ) , .D( u0_N406 ) , .Q( u0_R12_23 ) );
  DFF_X1 u0_R12_reg_24 (.CK( clk ) , .D( u0_N407 ) , .Q( u0_R12_24 ) );
  DFF_X1 u0_R12_reg_25 (.CK( clk ) , .D( u0_N408 ) , .Q( u0_R12_25 ) );
  DFF_X1 u0_R12_reg_26 (.CK( clk ) , .D( u0_N409 ) , .Q( u0_R12_26 ) );
  DFF_X1 u0_R12_reg_27 (.CK( clk ) , .D( u0_N410 ) , .Q( u0_R12_27 ) );
  DFF_X1 u0_R12_reg_28 (.CK( clk ) , .D( u0_N411 ) , .Q( u0_R12_28 ) );
  DFF_X1 u0_R12_reg_29 (.CK( clk ) , .D( u0_N412 ) , .Q( u0_R12_29 ) );
  DFF_X1 u0_R12_reg_3 (.CK( clk ) , .D( u0_N386 ) , .Q( u0_R12_3 ) );
  DFF_X1 u0_R12_reg_30 (.CK( clk ) , .D( u0_N413 ) , .Q( u0_R12_30 ) );
  DFF_X1 u0_R12_reg_31 (.CK( clk ) , .D( u0_N414 ) , .Q( u0_R12_31 ) );
  DFF_X1 u0_R12_reg_32 (.CK( clk ) , .D( u0_N415 ) , .Q( u0_R12_32 ) );
  DFF_X1 u0_R12_reg_4 (.CK( clk ) , .D( u0_N387 ) , .Q( u0_R12_4 ) );
  DFF_X1 u0_R12_reg_5 (.CK( clk ) , .D( u0_N388 ) , .Q( u0_R12_5 ) );
  DFF_X1 u0_R12_reg_6 (.CK( clk ) , .D( u0_N389 ) , .Q( u0_R12_6 ) );
  DFF_X1 u0_R12_reg_7 (.CK( clk ) , .D( u0_N390 ) , .Q( u0_R12_7 ) );
  DFF_X1 u0_R12_reg_8 (.CK( clk ) , .D( u0_N391 ) , .Q( u0_R12_8 ) );
  DFF_X1 u0_R12_reg_9 (.CK( clk ) , .D( u0_N392 ) , .Q( u0_R12_9 ) );
  DFF_X1 u0_R13_reg_1 (.CK( clk ) , .D( u0_N416 ) , .Q( u0_R13_1 ) );
  DFF_X1 u0_R13_reg_10 (.CK( clk ) , .D( u0_N425 ) , .Q( u0_R13_10 ) );
  DFF_X1 u0_R13_reg_11 (.CK( clk ) , .D( u0_N426 ) , .Q( u0_R13_11 ) );
  DFF_X1 u0_R13_reg_12 (.CK( clk ) , .D( u0_N427 ) , .Q( u0_R13_12 ) );
  DFF_X1 u0_R13_reg_13 (.CK( clk ) , .D( u0_N428 ) , .Q( u0_R13_13 ) );
  DFF_X1 u0_R13_reg_14 (.CK( clk ) , .D( u0_N429 ) , .Q( u0_R13_14 ) );
  DFF_X1 u0_R13_reg_15 (.CK( clk ) , .D( u0_N430 ) , .Q( u0_R13_15 ) );
  DFF_X1 u0_R13_reg_16 (.CK( clk ) , .D( u0_N431 ) , .Q( u0_R13_16 ) );
  DFF_X1 u0_R13_reg_17 (.CK( clk ) , .D( u0_N432 ) , .Q( u0_R13_17 ) );
  DFF_X1 u0_R13_reg_18 (.CK( clk ) , .D( u0_N433 ) , .Q( u0_R13_18 ) );
  DFF_X1 u0_R13_reg_19 (.CK( clk ) , .D( u0_N434 ) , .Q( u0_R13_19 ) );
  DFF_X1 u0_R13_reg_2 (.CK( clk ) , .D( u0_N417 ) , .Q( u0_R13_2 ) );
  DFF_X1 u0_R13_reg_20 (.CK( clk ) , .D( u0_N435 ) , .Q( u0_R13_20 ) );
  DFF_X1 u0_R13_reg_21 (.CK( clk ) , .D( u0_N436 ) , .Q( u0_R13_21 ) );
  DFF_X1 u0_R13_reg_22 (.CK( clk ) , .D( u0_N437 ) , .Q( u0_R13_22 ) );
  DFF_X1 u0_R13_reg_23 (.CK( clk ) , .D( u0_N438 ) , .Q( u0_R13_23 ) );
  DFF_X1 u0_R13_reg_24 (.CK( clk ) , .D( u0_N439 ) , .Q( u0_R13_24 ) );
  DFF_X1 u0_R13_reg_25 (.CK( clk ) , .D( u0_N440 ) , .Q( u0_R13_25 ) );
  DFF_X1 u0_R13_reg_26 (.CK( clk ) , .D( u0_N441 ) , .Q( u0_R13_26 ) );
  DFF_X1 u0_R13_reg_27 (.CK( clk ) , .D( u0_N442 ) , .Q( u0_R13_27 ) );
  DFF_X1 u0_R13_reg_28 (.CK( clk ) , .D( u0_N443 ) , .Q( u0_R13_28 ) );
  DFF_X1 u0_R13_reg_29 (.CK( clk ) , .D( u0_N444 ) , .Q( u0_R13_29 ) );
  DFF_X1 u0_R13_reg_3 (.CK( clk ) , .D( u0_N418 ) , .Q( u0_R13_3 ) );
  DFF_X1 u0_R13_reg_30 (.CK( clk ) , .D( u0_N445 ) , .Q( u0_R13_30 ) );
  DFF_X1 u0_R13_reg_31 (.CK( clk ) , .D( u0_N446 ) , .Q( u0_R13_31 ) );
  DFF_X1 u0_R13_reg_32 (.CK( clk ) , .D( u0_N447 ) , .Q( u0_R13_32 ) );
  DFF_X1 u0_R13_reg_4 (.CK( clk ) , .D( u0_N419 ) , .Q( u0_R13_4 ) );
  DFF_X1 u0_R13_reg_5 (.CK( clk ) , .D( u0_N420 ) , .Q( u0_R13_5 ) );
  DFF_X1 u0_R13_reg_6 (.CK( clk ) , .D( u0_N421 ) , .Q( u0_R13_6 ) );
  DFF_X1 u0_R13_reg_7 (.CK( clk ) , .D( u0_N422 ) , .Q( u0_R13_7 ) );
  DFF_X1 u0_R13_reg_8 (.CK( clk ) , .D( u0_N423 ) , .Q( u0_R13_8 ) );
  DFF_X1 u0_R13_reg_9 (.CK( clk ) , .D( u0_N424 ) , .Q( u0_R13_9 ) );
  DFF_X1 u0_R14_reg_1 (.CK( clk ) , .Q( u0_FP_33 ) , .D( u0_N448 ) );
  DFF_X1 u0_R14_reg_10 (.CK( clk ) , .Q( u0_FP_42 ) , .D( u0_N457 ) );
  DFF_X1 u0_R14_reg_11 (.CK( clk ) , .Q( u0_FP_43 ) , .D( u0_N458 ) );
  DFF_X1 u0_R14_reg_12 (.CK( clk ) , .Q( u0_FP_44 ) , .D( u0_N459 ) );
  DFF_X1 u0_R14_reg_13 (.CK( clk ) , .Q( u0_FP_45 ) , .D( u0_N460 ) );
  DFF_X1 u0_R14_reg_14 (.CK( clk ) , .Q( u0_FP_46 ) , .D( u0_N461 ) );
  DFF_X1 u0_R14_reg_15 (.CK( clk ) , .Q( u0_FP_47 ) , .D( u0_N462 ) );
  DFF_X1 u0_R14_reg_16 (.CK( clk ) , .Q( u0_FP_48 ) , .D( u0_N463 ) );
  DFF_X1 u0_R14_reg_17 (.CK( clk ) , .Q( u0_FP_49 ) , .D( u0_N464 ) );
  DFF_X1 u0_R14_reg_18 (.CK( clk ) , .Q( u0_FP_50 ) , .D( u0_N465 ) );
  DFF_X1 u0_R14_reg_19 (.CK( clk ) , .Q( u0_FP_51 ) , .D( u0_N466 ) );
  DFF_X1 u0_R14_reg_2 (.CK( clk ) , .Q( u0_FP_34 ) , .D( u0_N449 ) );
  DFF_X1 u0_R14_reg_20 (.CK( clk ) , .Q( u0_FP_52 ) , .D( u0_N467 ) );
  DFF_X1 u0_R14_reg_21 (.CK( clk ) , .Q( u0_FP_53 ) , .D( u0_N468 ) );
  DFF_X1 u0_R14_reg_22 (.CK( clk ) , .Q( u0_FP_54 ) , .D( u0_N469 ) );
  DFF_X1 u0_R14_reg_23 (.CK( clk ) , .Q( u0_FP_55 ) , .D( u0_N470 ) );
  DFF_X1 u0_R14_reg_24 (.CK( clk ) , .Q( u0_FP_56 ) , .D( u0_N471 ) );
  DFF_X1 u0_R14_reg_25 (.CK( clk ) , .Q( u0_FP_57 ) , .D( u0_N472 ) );
  DFF_X1 u0_R14_reg_26 (.CK( clk ) , .Q( u0_FP_58 ) , .D( u0_N473 ) );
  DFF_X1 u0_R14_reg_27 (.CK( clk ) , .Q( u0_FP_59 ) , .D( u0_N474 ) );
  DFF_X1 u0_R14_reg_28 (.CK( clk ) , .Q( u0_FP_60 ) , .D( u0_N475 ) );
  DFF_X1 u0_R14_reg_29 (.CK( clk ) , .Q( u0_FP_61 ) , .D( u0_N476 ) );
  DFF_X1 u0_R14_reg_3 (.CK( clk ) , .Q( u0_FP_35 ) , .D( u0_N450 ) );
  DFF_X1 u0_R14_reg_30 (.CK( clk ) , .Q( u0_FP_62 ) , .D( u0_N477 ) );
  DFF_X1 u0_R14_reg_31 (.CK( clk ) , .Q( u0_FP_63 ) , .D( u0_N478 ) );
  DFF_X1 u0_R14_reg_32 (.CK( clk ) , .Q( u0_FP_64 ) , .D( u0_N479 ) );
  DFF_X1 u0_R14_reg_4 (.CK( clk ) , .Q( u0_FP_36 ) , .D( u0_N451 ) );
  DFF_X1 u0_R14_reg_5 (.CK( clk ) , .Q( u0_FP_37 ) , .D( u0_N452 ) );
  DFF_X1 u0_R14_reg_6 (.CK( clk ) , .Q( u0_FP_38 ) , .D( u0_N453 ) );
  DFF_X1 u0_R14_reg_7 (.CK( clk ) , .Q( u0_FP_39 ) , .D( u0_N454 ) );
  DFF_X1 u0_R14_reg_8 (.CK( clk ) , .Q( u0_FP_40 ) , .D( u0_N455 ) );
  DFF_X1 u0_R14_reg_9 (.CK( clk ) , .Q( u0_FP_41 ) , .D( u0_N456 ) );
  DFF_X1 u0_R1_reg_1 (.CK( clk ) , .D( u0_N32 ) , .Q( u0_R1_1 ) );
  DFF_X1 u0_R1_reg_10 (.CK( clk ) , .D( u0_N41 ) , .Q( u0_R1_10 ) );
  DFF_X1 u0_R1_reg_11 (.CK( clk ) , .D( u0_N42 ) , .Q( u0_R1_11 ) );
  DFF_X1 u0_R1_reg_12 (.CK( clk ) , .D( u0_N43 ) , .Q( u0_R1_12 ) );
  DFF_X1 u0_R1_reg_13 (.CK( clk ) , .D( u0_N44 ) , .Q( u0_R1_13 ) );
  DFF_X1 u0_R1_reg_14 (.CK( clk ) , .D( u0_N45 ) , .Q( u0_R1_14 ) );
  DFF_X1 u0_R1_reg_15 (.CK( clk ) , .D( u0_N46 ) , .Q( u0_R1_15 ) );
  DFF_X1 u0_R1_reg_16 (.CK( clk ) , .D( u0_N47 ) , .Q( u0_R1_16 ) );
  DFF_X1 u0_R1_reg_17 (.CK( clk ) , .D( u0_N48 ) , .Q( u0_R1_17 ) );
  DFF_X1 u0_R1_reg_18 (.CK( clk ) , .D( u0_N49 ) , .Q( u0_R1_18 ) );
  DFF_X1 u0_R1_reg_19 (.CK( clk ) , .D( u0_N50 ) , .Q( u0_R1_19 ) );
  DFF_X1 u0_R1_reg_2 (.CK( clk ) , .D( u0_N33 ) , .Q( u0_R1_2 ) );
  DFF_X1 u0_R1_reg_20 (.CK( clk ) , .D( u0_N51 ) , .Q( u0_R1_20 ) );
  DFF_X1 u0_R1_reg_21 (.CK( clk ) , .D( u0_N52 ) , .Q( u0_R1_21 ) );
  DFF_X1 u0_R1_reg_22 (.CK( clk ) , .D( u0_N53 ) , .Q( u0_R1_22 ) );
  DFF_X1 u0_R1_reg_23 (.CK( clk ) , .D( u0_N54 ) , .Q( u0_R1_23 ) );
  DFF_X1 u0_R1_reg_24 (.CK( clk ) , .D( u0_N55 ) , .Q( u0_R1_24 ) );
  DFF_X1 u0_R1_reg_25 (.CK( clk ) , .D( u0_N56 ) , .Q( u0_R1_25 ) );
  DFF_X1 u0_R1_reg_26 (.CK( clk ) , .D( u0_N57 ) , .Q( u0_R1_26 ) );
  DFF_X1 u0_R1_reg_27 (.CK( clk ) , .D( u0_N58 ) , .Q( u0_R1_27 ) );
  DFF_X1 u0_R1_reg_28 (.CK( clk ) , .D( u0_N59 ) , .Q( u0_R1_28 ) );
  DFF_X1 u0_R1_reg_29 (.CK( clk ) , .D( u0_N60 ) , .Q( u0_R1_29 ) );
  DFF_X1 u0_R1_reg_3 (.CK( clk ) , .D( u0_N34 ) , .Q( u0_R1_3 ) );
  DFF_X1 u0_R1_reg_30 (.CK( clk ) , .D( u0_N61 ) , .Q( u0_R1_30 ) );
  DFF_X1 u0_R1_reg_31 (.CK( clk ) , .D( u0_N62 ) , .Q( u0_R1_31 ) );
  DFF_X1 u0_R1_reg_32 (.CK( clk ) , .D( u0_N63 ) , .Q( u0_R1_32 ) );
  DFF_X1 u0_R1_reg_4 (.CK( clk ) , .D( u0_N35 ) , .Q( u0_R1_4 ) );
  DFF_X1 u0_R1_reg_5 (.CK( clk ) , .D( u0_N36 ) , .Q( u0_R1_5 ) );
  DFF_X1 u0_R1_reg_6 (.CK( clk ) , .D( u0_N37 ) , .Q( u0_R1_6 ) );
  DFF_X1 u0_R1_reg_7 (.CK( clk ) , .D( u0_N38 ) , .Q( u0_R1_7 ) );
  DFF_X1 u0_R1_reg_8 (.CK( clk ) , .D( u0_N39 ) , .Q( u0_R1_8 ) );
  DFF_X1 u0_R1_reg_9 (.CK( clk ) , .D( u0_N40 ) , .Q( u0_R1_9 ) );
  DFF_X1 u0_R2_reg_1 (.CK( clk ) , .D( u0_N64 ) , .Q( u0_R2_1 ) );
  DFF_X1 u0_R2_reg_10 (.CK( clk ) , .D( u0_N73 ) , .Q( u0_R2_10 ) );
  DFF_X1 u0_R2_reg_11 (.CK( clk ) , .D( u0_N74 ) , .Q( u0_R2_11 ) );
  DFF_X1 u0_R2_reg_12 (.CK( clk ) , .D( u0_N75 ) , .Q( u0_R2_12 ) );
  DFF_X1 u0_R2_reg_13 (.CK( clk ) , .D( u0_N76 ) , .Q( u0_R2_13 ) );
  DFF_X1 u0_R2_reg_14 (.CK( clk ) , .D( u0_N77 ) , .Q( u0_R2_14 ) );
  DFF_X1 u0_R2_reg_15 (.CK( clk ) , .D( u0_N78 ) , .Q( u0_R2_15 ) );
  DFF_X1 u0_R2_reg_16 (.CK( clk ) , .D( u0_N79 ) , .Q( u0_R2_16 ) );
  DFF_X1 u0_R2_reg_17 (.CK( clk ) , .D( u0_N80 ) , .Q( u0_R2_17 ) );
  DFF_X1 u0_R2_reg_18 (.CK( clk ) , .D( u0_N81 ) , .Q( u0_R2_18 ) );
  DFF_X1 u0_R2_reg_19 (.CK( clk ) , .D( u0_N82 ) , .Q( u0_R2_19 ) );
  DFF_X1 u0_R2_reg_2 (.CK( clk ) , .D( u0_N65 ) , .Q( u0_R2_2 ) );
  DFF_X1 u0_R2_reg_20 (.CK( clk ) , .D( u0_N83 ) , .Q( u0_R2_20 ) );
  DFF_X1 u0_R2_reg_21 (.CK( clk ) , .D( u0_N84 ) , .Q( u0_R2_21 ) );
  DFF_X1 u0_R2_reg_22 (.CK( clk ) , .D( u0_N85 ) , .Q( u0_R2_22 ) );
  DFF_X1 u0_R2_reg_23 (.CK( clk ) , .D( u0_N86 ) , .Q( u0_R2_23 ) );
  DFF_X1 u0_R2_reg_24 (.CK( clk ) , .D( u0_N87 ) , .Q( u0_R2_24 ) );
  DFF_X1 u0_R2_reg_25 (.CK( clk ) , .D( u0_N88 ) , .Q( u0_R2_25 ) );
  DFF_X1 u0_R2_reg_26 (.CK( clk ) , .D( u0_N89 ) , .Q( u0_R2_26 ) );
  DFF_X1 u0_R2_reg_27 (.CK( clk ) , .D( u0_N90 ) , .Q( u0_R2_27 ) );
  DFF_X1 u0_R2_reg_28 (.CK( clk ) , .D( u0_N91 ) , .Q( u0_R2_28 ) );
  DFF_X1 u0_R2_reg_29 (.CK( clk ) , .D( u0_N92 ) , .Q( u0_R2_29 ) );
  DFF_X1 u0_R2_reg_3 (.CK( clk ) , .D( u0_N66 ) , .Q( u0_R2_3 ) );
  DFF_X1 u0_R2_reg_30 (.CK( clk ) , .D( u0_N93 ) , .Q( u0_R2_30 ) );
  DFF_X1 u0_R2_reg_31 (.CK( clk ) , .D( u0_N94 ) , .Q( u0_R2_31 ) );
  DFF_X1 u0_R2_reg_32 (.CK( clk ) , .D( u0_N95 ) , .Q( u0_R2_32 ) );
  DFF_X1 u0_R2_reg_4 (.CK( clk ) , .D( u0_N67 ) , .Q( u0_R2_4 ) );
  DFF_X1 u0_R2_reg_5 (.CK( clk ) , .D( u0_N68 ) , .Q( u0_R2_5 ) );
  DFF_X1 u0_R2_reg_6 (.CK( clk ) , .D( u0_N69 ) , .Q( u0_R2_6 ) );
  DFF_X1 u0_R2_reg_7 (.CK( clk ) , .D( u0_N70 ) , .Q( u0_R2_7 ) );
  DFF_X1 u0_R2_reg_8 (.CK( clk ) , .D( u0_N71 ) , .Q( u0_R2_8 ) );
  DFF_X1 u0_R2_reg_9 (.CK( clk ) , .D( u0_N72 ) , .Q( u0_R2_9 ) );
  DFF_X1 u0_R3_reg_1 (.CK( clk ) , .D( u0_N96 ) , .Q( u0_R3_1 ) );
  DFF_X1 u0_R3_reg_10 (.CK( clk ) , .D( u0_N105 ) , .Q( u0_R3_10 ) );
  DFF_X1 u0_R3_reg_11 (.CK( clk ) , .D( u0_N106 ) , .Q( u0_R3_11 ) );
  DFF_X1 u0_R3_reg_12 (.CK( clk ) , .D( u0_N107 ) , .Q( u0_R3_12 ) );
  DFF_X1 u0_R3_reg_13 (.CK( clk ) , .D( u0_N108 ) , .Q( u0_R3_13 ) );
  DFF_X1 u0_R3_reg_14 (.CK( clk ) , .D( u0_N109 ) , .Q( u0_R3_14 ) );
  DFF_X1 u0_R3_reg_15 (.CK( clk ) , .D( u0_N110 ) , .Q( u0_R3_15 ) );
  DFF_X1 u0_R3_reg_16 (.CK( clk ) , .D( u0_N111 ) , .Q( u0_R3_16 ) );
  DFF_X1 u0_R3_reg_17 (.CK( clk ) , .D( u0_N112 ) , .Q( u0_R3_17 ) );
  DFF_X1 u0_R3_reg_18 (.CK( clk ) , .D( u0_N113 ) , .Q( u0_R3_18 ) );
  DFF_X1 u0_R3_reg_19 (.CK( clk ) , .D( u0_N114 ) , .Q( u0_R3_19 ) );
  DFF_X1 u0_R3_reg_2 (.CK( clk ) , .D( u0_N97 ) , .Q( u0_R3_2 ) );
  DFF_X1 u0_R3_reg_20 (.CK( clk ) , .D( u0_N115 ) , .Q( u0_R3_20 ) );
  DFF_X1 u0_R3_reg_21 (.CK( clk ) , .D( u0_N116 ) , .Q( u0_R3_21 ) );
  DFF_X1 u0_R3_reg_22 (.CK( clk ) , .D( u0_N117 ) , .Q( u0_R3_22 ) );
  DFF_X1 u0_R3_reg_23 (.CK( clk ) , .D( u0_N118 ) , .Q( u0_R3_23 ) );
  DFF_X1 u0_R3_reg_24 (.CK( clk ) , .D( u0_N119 ) , .Q( u0_R3_24 ) );
  DFF_X1 u0_R3_reg_25 (.CK( clk ) , .D( u0_N120 ) , .Q( u0_R3_25 ) );
  DFF_X1 u0_R3_reg_26 (.CK( clk ) , .D( u0_N121 ) , .Q( u0_R3_26 ) );
  DFF_X1 u0_R3_reg_27 (.CK( clk ) , .D( u0_N122 ) , .Q( u0_R3_27 ) );
  DFF_X1 u0_R3_reg_28 (.CK( clk ) , .D( u0_N123 ) , .Q( u0_R3_28 ) );
  DFF_X1 u0_R3_reg_29 (.CK( clk ) , .D( u0_N124 ) , .Q( u0_R3_29 ) );
  DFF_X1 u0_R3_reg_3 (.CK( clk ) , .D( u0_N98 ) , .Q( u0_R3_3 ) );
  DFF_X1 u0_R3_reg_30 (.CK( clk ) , .D( u0_N125 ) , .Q( u0_R3_30 ) );
  DFF_X1 u0_R3_reg_31 (.CK( clk ) , .D( u0_N126 ) , .Q( u0_R3_31 ) );
  DFF_X1 u0_R3_reg_32 (.CK( clk ) , .D( u0_N127 ) , .Q( u0_R3_32 ) );
  DFF_X1 u0_R3_reg_4 (.CK( clk ) , .D( u0_N99 ) , .Q( u0_R3_4 ) );
  DFF_X1 u0_R3_reg_5 (.CK( clk ) , .D( u0_N100 ) , .Q( u0_R3_5 ) );
  DFF_X1 u0_R3_reg_6 (.CK( clk ) , .D( u0_N101 ) , .Q( u0_R3_6 ) );
  DFF_X1 u0_R3_reg_7 (.CK( clk ) , .D( u0_N102 ) , .Q( u0_R3_7 ) );
  DFF_X1 u0_R3_reg_8 (.CK( clk ) , .D( u0_N103 ) , .Q( u0_R3_8 ) );
  DFF_X1 u0_R3_reg_9 (.CK( clk ) , .D( u0_N104 ) , .Q( u0_R3_9 ) );
  DFF_X1 u0_R4_reg_1 (.CK( clk ) , .D( u0_N128 ) , .Q( u0_R4_1 ) );
  DFF_X1 u0_R4_reg_10 (.CK( clk ) , .D( u0_N137 ) , .Q( u0_R4_10 ) );
  DFF_X1 u0_R4_reg_11 (.CK( clk ) , .D( u0_N138 ) , .Q( u0_R4_11 ) );
  DFF_X1 u0_R4_reg_12 (.CK( clk ) , .D( u0_N139 ) , .Q( u0_R4_12 ) );
  DFF_X1 u0_R4_reg_13 (.CK( clk ) , .D( u0_N140 ) , .Q( u0_R4_13 ) );
  DFF_X1 u0_R4_reg_14 (.CK( clk ) , .D( u0_N141 ) , .Q( u0_R4_14 ) );
  DFF_X1 u0_R4_reg_15 (.CK( clk ) , .D( u0_N142 ) , .Q( u0_R4_15 ) );
  DFF_X1 u0_R4_reg_16 (.CK( clk ) , .D( u0_N143 ) , .Q( u0_R4_16 ) );
  DFF_X1 u0_R4_reg_17 (.CK( clk ) , .D( u0_N144 ) , .Q( u0_R4_17 ) );
  DFF_X1 u0_R4_reg_18 (.CK( clk ) , .D( u0_N145 ) , .Q( u0_R4_18 ) );
  DFF_X1 u0_R4_reg_19 (.CK( clk ) , .D( u0_N146 ) , .Q( u0_R4_19 ) );
  DFF_X1 u0_R4_reg_2 (.CK( clk ) , .D( u0_N129 ) , .Q( u0_R4_2 ) );
  DFF_X1 u0_R4_reg_20 (.CK( clk ) , .D( u0_N147 ) , .Q( u0_R4_20 ) );
  DFF_X1 u0_R4_reg_21 (.CK( clk ) , .D( u0_N148 ) , .Q( u0_R4_21 ) );
  DFF_X1 u0_R4_reg_22 (.CK( clk ) , .D( u0_N149 ) , .Q( u0_R4_22 ) );
  DFF_X1 u0_R4_reg_23 (.CK( clk ) , .D( u0_N150 ) , .Q( u0_R4_23 ) );
  DFF_X1 u0_R4_reg_24 (.CK( clk ) , .D( u0_N151 ) , .Q( u0_R4_24 ) );
  DFF_X1 u0_R4_reg_25 (.CK( clk ) , .D( u0_N152 ) , .Q( u0_R4_25 ) );
  DFF_X1 u0_R4_reg_26 (.CK( clk ) , .D( u0_N153 ) , .Q( u0_R4_26 ) );
  DFF_X1 u0_R4_reg_27 (.CK( clk ) , .D( u0_N154 ) , .Q( u0_R4_27 ) );
  DFF_X1 u0_R4_reg_28 (.CK( clk ) , .D( u0_N155 ) , .Q( u0_R4_28 ) );
  DFF_X1 u0_R4_reg_29 (.CK( clk ) , .D( u0_N156 ) , .Q( u0_R4_29 ) );
  DFF_X1 u0_R4_reg_3 (.CK( clk ) , .D( u0_N130 ) , .Q( u0_R4_3 ) );
  DFF_X1 u0_R4_reg_30 (.CK( clk ) , .D( u0_N157 ) , .Q( u0_R4_30 ) );
  DFF_X1 u0_R4_reg_31 (.CK( clk ) , .D( u0_N158 ) , .Q( u0_R4_31 ) );
  DFF_X1 u0_R4_reg_32 (.CK( clk ) , .D( u0_N159 ) , .Q( u0_R4_32 ) );
  DFF_X1 u0_R4_reg_4 (.CK( clk ) , .D( u0_N131 ) , .Q( u0_R4_4 ) );
  DFF_X1 u0_R4_reg_5 (.CK( clk ) , .D( u0_N132 ) , .Q( u0_R4_5 ) );
  DFF_X1 u0_R4_reg_6 (.CK( clk ) , .D( u0_N133 ) , .Q( u0_R4_6 ) );
  DFF_X1 u0_R4_reg_7 (.CK( clk ) , .D( u0_N134 ) , .Q( u0_R4_7 ) );
  DFF_X1 u0_R4_reg_8 (.CK( clk ) , .D( u0_N135 ) , .Q( u0_R4_8 ) );
  DFF_X1 u0_R4_reg_9 (.CK( clk ) , .D( u0_N136 ) , .Q( u0_R4_9 ) );
  DFF_X1 u0_R5_reg_1 (.CK( clk ) , .D( u0_N160 ) , .Q( u0_R5_1 ) );
  DFF_X1 u0_R5_reg_10 (.CK( clk ) , .D( u0_N169 ) , .Q( u0_R5_10 ) );
  DFF_X1 u0_R5_reg_11 (.CK( clk ) , .D( u0_N170 ) , .Q( u0_R5_11 ) );
  DFF_X1 u0_R5_reg_12 (.CK( clk ) , .D( u0_N171 ) , .Q( u0_R5_12 ) );
  DFF_X1 u0_R5_reg_13 (.CK( clk ) , .D( u0_N172 ) , .Q( u0_R5_13 ) );
  DFF_X1 u0_R5_reg_14 (.CK( clk ) , .D( u0_N173 ) , .Q( u0_R5_14 ) );
  DFF_X1 u0_R5_reg_15 (.CK( clk ) , .D( u0_N174 ) , .Q( u0_R5_15 ) );
  DFF_X1 u0_R5_reg_16 (.CK( clk ) , .D( u0_N175 ) , .Q( u0_R5_16 ) );
  DFF_X1 u0_R5_reg_17 (.CK( clk ) , .D( u0_N176 ) , .Q( u0_R5_17 ) );
  DFF_X1 u0_R5_reg_18 (.CK( clk ) , .D( u0_N177 ) , .Q( u0_R5_18 ) );
  DFF_X1 u0_R5_reg_19 (.CK( clk ) , .D( u0_N178 ) , .Q( u0_R5_19 ) );
  DFF_X1 u0_R5_reg_2 (.CK( clk ) , .D( u0_N161 ) , .Q( u0_R5_2 ) );
  DFF_X1 u0_R5_reg_20 (.CK( clk ) , .D( u0_N179 ) , .Q( u0_R5_20 ) );
  DFF_X1 u0_R5_reg_21 (.CK( clk ) , .D( u0_N180 ) , .Q( u0_R5_21 ) );
  DFF_X1 u0_R5_reg_22 (.CK( clk ) , .D( u0_N181 ) , .Q( u0_R5_22 ) );
  DFF_X1 u0_R5_reg_23 (.CK( clk ) , .D( u0_N182 ) , .Q( u0_R5_23 ) );
  DFF_X1 u0_R5_reg_24 (.CK( clk ) , .D( u0_N183 ) , .Q( u0_R5_24 ) );
  DFF_X1 u0_R5_reg_25 (.CK( clk ) , .D( u0_N184 ) , .Q( u0_R5_25 ) );
  DFF_X1 u0_R5_reg_26 (.CK( clk ) , .D( u0_N185 ) , .Q( u0_R5_26 ) );
  DFF_X1 u0_R5_reg_27 (.CK( clk ) , .D( u0_N186 ) , .Q( u0_R5_27 ) );
  DFF_X1 u0_R5_reg_28 (.CK( clk ) , .D( u0_N187 ) , .Q( u0_R5_28 ) );
  DFF_X1 u0_R5_reg_29 (.CK( clk ) , .D( u0_N188 ) , .Q( u0_R5_29 ) );
  DFF_X1 u0_R5_reg_3 (.CK( clk ) , .D( u0_N162 ) , .Q( u0_R5_3 ) );
  DFF_X1 u0_R5_reg_30 (.CK( clk ) , .D( u0_N189 ) , .Q( u0_R5_30 ) );
  DFF_X1 u0_R5_reg_31 (.CK( clk ) , .D( u0_N190 ) , .Q( u0_R5_31 ) );
  DFF_X1 u0_R5_reg_32 (.CK( clk ) , .D( u0_N191 ) , .Q( u0_R5_32 ) );
  DFF_X1 u0_R5_reg_4 (.CK( clk ) , .D( u0_N163 ) , .Q( u0_R5_4 ) );
  DFF_X1 u0_R5_reg_5 (.CK( clk ) , .D( u0_N164 ) , .Q( u0_R5_5 ) );
  DFF_X1 u0_R5_reg_6 (.CK( clk ) , .D( u0_N165 ) , .Q( u0_R5_6 ) );
  DFF_X1 u0_R5_reg_7 (.CK( clk ) , .D( u0_N166 ) , .Q( u0_R5_7 ) );
  DFF_X1 u0_R5_reg_8 (.CK( clk ) , .D( u0_N167 ) , .Q( u0_R5_8 ) );
  DFF_X1 u0_R5_reg_9 (.CK( clk ) , .D( u0_N168 ) , .Q( u0_R5_9 ) );
  DFF_X1 u0_R6_reg_1 (.CK( clk ) , .D( u0_N192 ) , .Q( u0_R6_1 ) );
  DFF_X1 u0_R6_reg_10 (.CK( clk ) , .D( u0_N201 ) , .Q( u0_R6_10 ) );
  DFF_X1 u0_R6_reg_11 (.CK( clk ) , .D( u0_N202 ) , .Q( u0_R6_11 ) );
  DFF_X1 u0_R6_reg_12 (.CK( clk ) , .D( u0_N203 ) , .Q( u0_R6_12 ) );
  DFF_X1 u0_R6_reg_13 (.CK( clk ) , .D( u0_N204 ) , .Q( u0_R6_13 ) );
  DFF_X1 u0_R6_reg_14 (.CK( clk ) , .D( u0_N205 ) , .Q( u0_R6_14 ) );
  DFF_X1 u0_R6_reg_15 (.CK( clk ) , .D( u0_N206 ) , .Q( u0_R6_15 ) );
  DFF_X1 u0_R6_reg_16 (.CK( clk ) , .D( u0_N207 ) , .Q( u0_R6_16 ) );
  DFF_X1 u0_R6_reg_17 (.CK( clk ) , .D( u0_N208 ) , .Q( u0_R6_17 ) );
  DFF_X1 u0_R6_reg_18 (.CK( clk ) , .D( u0_N209 ) , .Q( u0_R6_18 ) );
  DFF_X1 u0_R6_reg_19 (.CK( clk ) , .D( u0_N210 ) , .Q( u0_R6_19 ) );
  DFF_X1 u0_R6_reg_2 (.CK( clk ) , .D( u0_N193 ) , .Q( u0_R6_2 ) );
  DFF_X1 u0_R6_reg_20 (.CK( clk ) , .D( u0_N211 ) , .Q( u0_R6_20 ) );
  DFF_X1 u0_R6_reg_21 (.CK( clk ) , .D( u0_N212 ) , .Q( u0_R6_21 ) );
  DFF_X1 u0_R6_reg_22 (.CK( clk ) , .D( u0_N213 ) , .Q( u0_R6_22 ) );
  DFF_X1 u0_R6_reg_23 (.CK( clk ) , .D( u0_N214 ) , .Q( u0_R6_23 ) );
  DFF_X1 u0_R6_reg_24 (.CK( clk ) , .D( u0_N215 ) , .Q( u0_R6_24 ) );
  DFF_X1 u0_R6_reg_25 (.CK( clk ) , .D( u0_N216 ) , .Q( u0_R6_25 ) );
  DFF_X1 u0_R6_reg_26 (.CK( clk ) , .D( u0_N217 ) , .Q( u0_R6_26 ) );
  DFF_X1 u0_R6_reg_27 (.CK( clk ) , .D( u0_N218 ) , .Q( u0_R6_27 ) );
  DFF_X1 u0_R6_reg_28 (.CK( clk ) , .D( u0_N219 ) , .Q( u0_R6_28 ) );
  DFF_X1 u0_R6_reg_29 (.CK( clk ) , .D( u0_N220 ) , .Q( u0_R6_29 ) );
  DFF_X1 u0_R6_reg_3 (.CK( clk ) , .D( u0_N194 ) , .Q( u0_R6_3 ) );
  DFF_X1 u0_R6_reg_30 (.CK( clk ) , .D( u0_N221 ) , .Q( u0_R6_30 ) );
  DFF_X1 u0_R6_reg_31 (.CK( clk ) , .D( u0_N222 ) , .Q( u0_R6_31 ) );
  DFF_X1 u0_R6_reg_32 (.CK( clk ) , .D( u0_N223 ) , .Q( u0_R6_32 ) );
  DFF_X1 u0_R6_reg_4 (.CK( clk ) , .D( u0_N195 ) , .Q( u0_R6_4 ) );
  DFF_X1 u0_R6_reg_5 (.CK( clk ) , .D( u0_N196 ) , .Q( u0_R6_5 ) );
  DFF_X1 u0_R6_reg_6 (.CK( clk ) , .D( u0_N197 ) , .Q( u0_R6_6 ) );
  DFF_X1 u0_R6_reg_7 (.CK( clk ) , .D( u0_N198 ) , .Q( u0_R6_7 ) );
  DFF_X1 u0_R6_reg_8 (.CK( clk ) , .D( u0_N199 ) , .Q( u0_R6_8 ) );
  DFF_X1 u0_R6_reg_9 (.CK( clk ) , .D( u0_N200 ) , .Q( u0_R6_9 ) );
  DFF_X1 u0_R7_reg_1 (.CK( clk ) , .D( u0_N224 ) , .Q( u0_R7_1 ) );
  DFF_X1 u0_R7_reg_10 (.CK( clk ) , .D( u0_N233 ) , .Q( u0_R7_10 ) );
  DFF_X1 u0_R7_reg_11 (.CK( clk ) , .D( u0_N234 ) , .Q( u0_R7_11 ) );
  DFF_X1 u0_R7_reg_12 (.CK( clk ) , .D( u0_N235 ) , .Q( u0_R7_12 ) );
  DFF_X1 u0_R7_reg_13 (.CK( clk ) , .D( u0_N236 ) , .Q( u0_R7_13 ) );
  DFF_X1 u0_R7_reg_14 (.CK( clk ) , .D( u0_N237 ) , .Q( u0_R7_14 ) );
  DFF_X1 u0_R7_reg_15 (.CK( clk ) , .D( u0_N238 ) , .Q( u0_R7_15 ) );
  DFF_X1 u0_R7_reg_16 (.CK( clk ) , .D( u0_N239 ) , .Q( u0_R7_16 ) );
  DFF_X1 u0_R7_reg_17 (.CK( clk ) , .D( u0_N240 ) , .Q( u0_R7_17 ) );
  DFF_X1 u0_R7_reg_18 (.CK( clk ) , .D( u0_N241 ) , .Q( u0_R7_18 ) );
  DFF_X1 u0_R7_reg_19 (.CK( clk ) , .D( u0_N242 ) , .Q( u0_R7_19 ) );
  DFF_X1 u0_R7_reg_2 (.CK( clk ) , .D( u0_N225 ) , .Q( u0_R7_2 ) );
  DFF_X1 u0_R7_reg_20 (.CK( clk ) , .D( u0_N243 ) , .Q( u0_R7_20 ) );
  DFF_X1 u0_R7_reg_21 (.CK( clk ) , .D( u0_N244 ) , .Q( u0_R7_21 ) );
  DFF_X1 u0_R7_reg_22 (.CK( clk ) , .D( u0_N245 ) , .Q( u0_R7_22 ) );
  DFF_X1 u0_R7_reg_23 (.CK( clk ) , .D( u0_N246 ) , .Q( u0_R7_23 ) );
  DFF_X1 u0_R7_reg_24 (.CK( clk ) , .D( u0_N247 ) , .Q( u0_R7_24 ) );
  DFF_X1 u0_R7_reg_25 (.CK( clk ) , .D( u0_N248 ) , .Q( u0_R7_25 ) );
  DFF_X1 u0_R7_reg_26 (.CK( clk ) , .D( u0_N249 ) , .Q( u0_R7_26 ) );
  DFF_X1 u0_R7_reg_27 (.CK( clk ) , .D( u0_N250 ) , .Q( u0_R7_27 ) );
  DFF_X1 u0_R7_reg_28 (.CK( clk ) , .D( u0_N251 ) , .Q( u0_R7_28 ) );
  DFF_X1 u0_R7_reg_29 (.CK( clk ) , .D( u0_N252 ) , .Q( u0_R7_29 ) );
  DFF_X1 u0_R7_reg_3 (.CK( clk ) , .D( u0_N226 ) , .Q( u0_R7_3 ) );
  DFF_X1 u0_R7_reg_30 (.CK( clk ) , .D( u0_N253 ) , .Q( u0_R7_30 ) );
  DFF_X1 u0_R7_reg_31 (.CK( clk ) , .D( u0_N254 ) , .Q( u0_R7_31 ) );
  DFF_X1 u0_R7_reg_32 (.CK( clk ) , .D( u0_N255 ) , .Q( u0_R7_32 ) );
  DFF_X1 u0_R7_reg_4 (.CK( clk ) , .D( u0_N227 ) , .Q( u0_R7_4 ) );
  DFF_X1 u0_R7_reg_5 (.CK( clk ) , .D( u0_N228 ) , .Q( u0_R7_5 ) );
  DFF_X1 u0_R7_reg_6 (.CK( clk ) , .D( u0_N229 ) , .Q( u0_R7_6 ) );
  DFF_X1 u0_R7_reg_7 (.CK( clk ) , .D( u0_N230 ) , .Q( u0_R7_7 ) );
  DFF_X1 u0_R7_reg_8 (.CK( clk ) , .D( u0_N231 ) , .Q( u0_R7_8 ) );
  DFF_X1 u0_R7_reg_9 (.CK( clk ) , .D( u0_N232 ) , .Q( u0_R7_9 ) );
  DFF_X1 u0_R8_reg_1 (.CK( clk ) , .D( u0_N256 ) , .Q( u0_R8_1 ) );
  DFF_X1 u0_R8_reg_10 (.CK( clk ) , .D( u0_N265 ) , .Q( u0_R8_10 ) );
  DFF_X1 u0_R8_reg_11 (.CK( clk ) , .D( u0_N266 ) , .Q( u0_R8_11 ) );
  DFF_X1 u0_R8_reg_12 (.CK( clk ) , .D( u0_N267 ) , .Q( u0_R8_12 ) );
  DFF_X1 u0_R8_reg_13 (.CK( clk ) , .D( u0_N268 ) , .Q( u0_R8_13 ) );
  DFF_X1 u0_R8_reg_14 (.CK( clk ) , .D( u0_N269 ) , .Q( u0_R8_14 ) );
  DFF_X1 u0_R8_reg_15 (.CK( clk ) , .D( u0_N270 ) , .Q( u0_R8_15 ) );
  DFF_X1 u0_R8_reg_16 (.CK( clk ) , .D( u0_N271 ) , .Q( u0_R8_16 ) );
  DFF_X1 u0_R8_reg_17 (.CK( clk ) , .D( u0_N272 ) , .Q( u0_R8_17 ) );
  DFF_X1 u0_R8_reg_18 (.CK( clk ) , .D( u0_N273 ) , .Q( u0_R8_18 ) );
  DFF_X1 u0_R8_reg_19 (.CK( clk ) , .D( u0_N274 ) , .Q( u0_R8_19 ) );
  DFF_X1 u0_R8_reg_2 (.CK( clk ) , .D( u0_N257 ) , .Q( u0_R8_2 ) );
  DFF_X1 u0_R8_reg_20 (.CK( clk ) , .D( u0_N275 ) , .Q( u0_R8_20 ) );
  DFF_X1 u0_R8_reg_21 (.CK( clk ) , .D( u0_N276 ) , .Q( u0_R8_21 ) );
  DFF_X1 u0_R8_reg_22 (.CK( clk ) , .D( u0_N277 ) , .Q( u0_R8_22 ) );
  DFF_X1 u0_R8_reg_23 (.CK( clk ) , .D( u0_N278 ) , .Q( u0_R8_23 ) );
  DFF_X1 u0_R8_reg_24 (.CK( clk ) , .D( u0_N279 ) , .Q( u0_R8_24 ) );
  DFF_X1 u0_R8_reg_25 (.CK( clk ) , .D( u0_N280 ) , .Q( u0_R8_25 ) );
  DFF_X1 u0_R8_reg_26 (.CK( clk ) , .D( u0_N281 ) , .Q( u0_R8_26 ) );
  DFF_X1 u0_R8_reg_27 (.CK( clk ) , .D( u0_N282 ) , .Q( u0_R8_27 ) );
  DFF_X1 u0_R8_reg_28 (.CK( clk ) , .D( u0_N283 ) , .Q( u0_R8_28 ) );
  DFF_X1 u0_R8_reg_29 (.CK( clk ) , .D( u0_N284 ) , .Q( u0_R8_29 ) );
  DFF_X1 u0_R8_reg_3 (.CK( clk ) , .D( u0_N258 ) , .Q( u0_R8_3 ) );
  DFF_X1 u0_R8_reg_30 (.CK( clk ) , .D( u0_N285 ) , .Q( u0_R8_30 ) );
  DFF_X1 u0_R8_reg_31 (.CK( clk ) , .D( u0_N286 ) , .Q( u0_R8_31 ) );
  DFF_X1 u0_R8_reg_32 (.CK( clk ) , .D( u0_N287 ) , .Q( u0_R8_32 ) );
  DFF_X1 u0_R8_reg_4 (.CK( clk ) , .D( u0_N259 ) , .Q( u0_R8_4 ) );
  DFF_X1 u0_R8_reg_5 (.CK( clk ) , .D( u0_N260 ) , .Q( u0_R8_5 ) );
  DFF_X1 u0_R8_reg_6 (.CK( clk ) , .D( u0_N261 ) , .Q( u0_R8_6 ) );
  DFF_X1 u0_R8_reg_7 (.CK( clk ) , .D( u0_N262 ) , .Q( u0_R8_7 ) );
  DFF_X1 u0_R8_reg_8 (.CK( clk ) , .D( u0_N263 ) , .Q( u0_R8_8 ) );
  DFF_X1 u0_R8_reg_9 (.CK( clk ) , .D( u0_N264 ) , .Q( u0_R8_9 ) );
  DFF_X1 u0_R9_reg_1 (.CK( clk ) , .D( u0_N288 ) , .Q( u0_R9_1 ) );
  DFF_X1 u0_R9_reg_10 (.CK( clk ) , .D( u0_N297 ) , .Q( u0_R9_10 ) );
  DFF_X1 u0_R9_reg_11 (.CK( clk ) , .D( u0_N298 ) , .Q( u0_R9_11 ) );
  DFF_X1 u0_R9_reg_12 (.CK( clk ) , .D( u0_N299 ) , .Q( u0_R9_12 ) );
  DFF_X1 u0_R9_reg_13 (.CK( clk ) , .D( u0_N300 ) , .Q( u0_R9_13 ) );
  DFF_X1 u0_R9_reg_14 (.CK( clk ) , .D( u0_N301 ) , .Q( u0_R9_14 ) );
  DFF_X1 u0_R9_reg_15 (.CK( clk ) , .D( u0_N302 ) , .Q( u0_R9_15 ) );
  DFF_X1 u0_R9_reg_16 (.CK( clk ) , .D( u0_N303 ) , .Q( u0_R9_16 ) );
  DFF_X1 u0_R9_reg_17 (.CK( clk ) , .D( u0_N304 ) , .Q( u0_R9_17 ) );
  DFF_X1 u0_R9_reg_18 (.CK( clk ) , .D( u0_N305 ) , .Q( u0_R9_18 ) );
  DFF_X1 u0_R9_reg_19 (.CK( clk ) , .D( u0_N306 ) , .Q( u0_R9_19 ) );
  DFF_X1 u0_R9_reg_2 (.CK( clk ) , .D( u0_N289 ) , .Q( u0_R9_2 ) );
  DFF_X1 u0_R9_reg_20 (.CK( clk ) , .D( u0_N307 ) , .Q( u0_R9_20 ) );
  DFF_X1 u0_R9_reg_21 (.CK( clk ) , .D( u0_N308 ) , .Q( u0_R9_21 ) );
  DFF_X1 u0_R9_reg_22 (.CK( clk ) , .D( u0_N309 ) , .Q( u0_R9_22 ) );
  DFF_X1 u0_R9_reg_23 (.CK( clk ) , .D( u0_N310 ) , .Q( u0_R9_23 ) );
  DFF_X1 u0_R9_reg_24 (.CK( clk ) , .D( u0_N311 ) , .Q( u0_R9_24 ) );
  DFF_X1 u0_R9_reg_25 (.CK( clk ) , .D( u0_N312 ) , .Q( u0_R9_25 ) );
  DFF_X1 u0_R9_reg_26 (.CK( clk ) , .D( u0_N313 ) , .Q( u0_R9_26 ) );
  DFF_X1 u0_R9_reg_27 (.CK( clk ) , .D( u0_N314 ) , .Q( u0_R9_27 ) );
  DFF_X1 u0_R9_reg_28 (.CK( clk ) , .D( u0_N315 ) , .Q( u0_R9_28 ) );
  DFF_X1 u0_R9_reg_29 (.CK( clk ) , .D( u0_N316 ) , .Q( u0_R9_29 ) );
  DFF_X1 u0_R9_reg_3 (.CK( clk ) , .D( u0_N290 ) , .Q( u0_R9_3 ) );
  DFF_X1 u0_R9_reg_30 (.CK( clk ) , .D( u0_N317 ) , .Q( u0_R9_30 ) );
  DFF_X1 u0_R9_reg_31 (.CK( clk ) , .D( u0_N318 ) , .Q( u0_R9_31 ) );
  DFF_X1 u0_R9_reg_32 (.CK( clk ) , .D( u0_N319 ) , .Q( u0_R9_32 ) );
  DFF_X1 u0_R9_reg_4 (.CK( clk ) , .D( u0_N291 ) , .Q( u0_R9_4 ) );
  DFF_X1 u0_R9_reg_5 (.CK( clk ) , .D( u0_N292 ) , .Q( u0_R9_5 ) );
  DFF_X1 u0_R9_reg_6 (.CK( clk ) , .D( u0_N293 ) , .Q( u0_R9_6 ) );
  DFF_X1 u0_R9_reg_7 (.CK( clk ) , .D( u0_N294 ) , .Q( u0_R9_7 ) );
  DFF_X1 u0_R9_reg_8 (.CK( clk ) , .D( u0_N295 ) , .Q( u0_R9_8 ) );
  DFF_X1 u0_R9_reg_9 (.CK( clk ) , .D( u0_N296 ) , .Q( u0_R9_9 ) );
  DFF_X1 u0_desIn_r_reg_0 (.CK( clk ) , .D( desIn[0] ) , .Q( u0_desIn_r_0 ) );
  DFF_X1 u0_desIn_r_reg_1 (.CK( clk ) , .D( desIn[1] ) , .Q( u0_desIn_r_1 ) );
  DFF_X1 u0_desIn_r_reg_10 (.CK( clk ) , .D( desIn[10] ) , .Q( u0_desIn_r_10 ) );
  DFF_X1 u0_desIn_r_reg_11 (.CK( clk ) , .D( desIn[11] ) , .Q( u0_desIn_r_11 ) );
  DFF_X1 u0_desIn_r_reg_12 (.CK( clk ) , .D( desIn[12] ) , .Q( u0_desIn_r_12 ) );
  DFF_X1 u0_desIn_r_reg_13 (.CK( clk ) , .D( desIn[13] ) , .Q( u0_desIn_r_13 ) );
  DFF_X1 u0_desIn_r_reg_14 (.CK( clk ) , .D( desIn[14] ) , .Q( u0_desIn_r_14 ) );
  DFF_X1 u0_desIn_r_reg_15 (.CK( clk ) , .D( desIn[15] ) , .Q( u0_desIn_r_15 ) );
  DFF_X1 u0_desIn_r_reg_16 (.CK( clk ) , .D( desIn[16] ) , .Q( u0_desIn_r_16 ) );
  DFF_X1 u0_desIn_r_reg_17 (.CK( clk ) , .D( desIn[17] ) , .Q( u0_desIn_r_17 ) );
  DFF_X1 u0_desIn_r_reg_18 (.CK( clk ) , .D( desIn[18] ) , .Q( u0_desIn_r_18 ) );
  DFF_X1 u0_desIn_r_reg_19 (.CK( clk ) , .D( desIn[19] ) , .Q( u0_desIn_r_19 ) );
  DFF_X1 u0_desIn_r_reg_2 (.CK( clk ) , .D( desIn[2] ) , .Q( u0_desIn_r_2 ) );
  DFF_X1 u0_desIn_r_reg_20 (.CK( clk ) , .D( desIn[20] ) , .Q( u0_desIn_r_20 ) );
  DFF_X1 u0_desIn_r_reg_21 (.CK( clk ) , .D( desIn[21] ) , .Q( u0_desIn_r_21 ) );
  DFF_X1 u0_desIn_r_reg_22 (.CK( clk ) , .D( desIn[22] ) , .Q( u0_desIn_r_22 ) );
  DFF_X1 u0_desIn_r_reg_23 (.CK( clk ) , .D( desIn[23] ) , .Q( u0_desIn_r_23 ) );
  DFF_X1 u0_desIn_r_reg_24 (.CK( clk ) , .D( desIn[24] ) , .Q( u0_desIn_r_24 ) );
  DFF_X1 u0_desIn_r_reg_25 (.CK( clk ) , .D( desIn[25] ) , .Q( u0_desIn_r_25 ) );
  DFF_X1 u0_desIn_r_reg_26 (.CK( clk ) , .D( desIn[26] ) , .Q( u0_desIn_r_26 ) );
  DFF_X1 u0_desIn_r_reg_27 (.CK( clk ) , .D( desIn[27] ) , .Q( u0_desIn_r_27 ) );
  DFF_X1 u0_desIn_r_reg_28 (.CK( clk ) , .D( desIn[28] ) , .Q( u0_desIn_r_28 ) );
  DFF_X1 u0_desIn_r_reg_29 (.CK( clk ) , .D( desIn[29] ) , .Q( u0_desIn_r_29 ) );
  DFF_X1 u0_desIn_r_reg_3 (.CK( clk ) , .D( desIn[3] ) , .Q( u0_desIn_r_3 ) );
  DFF_X1 u0_desIn_r_reg_30 (.CK( clk ) , .D( desIn[30] ) , .Q( u0_desIn_r_30 ) );
  DFF_X1 u0_desIn_r_reg_31 (.CK( clk ) , .D( desIn[31] ) , .Q( u0_desIn_r_31 ) );
  DFF_X1 u0_desIn_r_reg_32 (.CK( clk ) , .D( desIn[32] ) , .Q( u0_desIn_r_32 ) );
  DFF_X1 u0_desIn_r_reg_33 (.CK( clk ) , .D( desIn[33] ) , .Q( u0_desIn_r_33 ) );
  DFF_X1 u0_desIn_r_reg_34 (.CK( clk ) , .D( desIn[34] ) , .Q( u0_desIn_r_34 ) );
  DFF_X1 u0_desIn_r_reg_35 (.CK( clk ) , .D( desIn[35] ) , .Q( u0_desIn_r_35 ) );
  DFF_X1 u0_desIn_r_reg_36 (.CK( clk ) , .D( desIn[36] ) , .Q( u0_desIn_r_36 ) );
  DFF_X1 u0_desIn_r_reg_37 (.CK( clk ) , .D( desIn[37] ) , .Q( u0_desIn_r_37 ) );
  DFF_X1 u0_desIn_r_reg_38 (.CK( clk ) , .D( desIn[38] ) , .Q( u0_desIn_r_38 ) );
  DFF_X1 u0_desIn_r_reg_39 (.CK( clk ) , .D( desIn[39] ) , .Q( u0_desIn_r_39 ) );
  DFF_X1 u0_desIn_r_reg_4 (.CK( clk ) , .D( desIn[4] ) , .Q( u0_desIn_r_4 ) );
  DFF_X1 u0_desIn_r_reg_40 (.CK( clk ) , .D( desIn[40] ) , .Q( u0_desIn_r_40 ) );
  DFF_X1 u0_desIn_r_reg_41 (.CK( clk ) , .D( desIn[41] ) , .Q( u0_desIn_r_41 ) );
  DFF_X1 u0_desIn_r_reg_42 (.CK( clk ) , .D( desIn[42] ) , .Q( u0_desIn_r_42 ) );
  DFF_X1 u0_desIn_r_reg_43 (.CK( clk ) , .D( desIn[43] ) , .Q( u0_desIn_r_43 ) );
  DFF_X1 u0_desIn_r_reg_44 (.CK( clk ) , .D( desIn[44] ) , .Q( u0_desIn_r_44 ) );
  DFF_X1 u0_desIn_r_reg_45 (.CK( clk ) , .D( desIn[45] ) , .Q( u0_desIn_r_45 ) );
  DFF_X1 u0_desIn_r_reg_46 (.CK( clk ) , .D( desIn[46] ) , .Q( u0_desIn_r_46 ) );
  DFF_X1 u0_desIn_r_reg_47 (.CK( clk ) , .D( desIn[47] ) , .Q( u0_desIn_r_47 ) );
  DFF_X1 u0_desIn_r_reg_48 (.CK( clk ) , .D( desIn[48] ) , .Q( u0_desIn_r_48 ) );
  DFF_X1 u0_desIn_r_reg_49 (.CK( clk ) , .D( desIn[49] ) , .Q( u0_desIn_r_49 ) );
  DFF_X1 u0_desIn_r_reg_5 (.CK( clk ) , .D( desIn[5] ) , .Q( u0_desIn_r_5 ) );
  DFF_X1 u0_desIn_r_reg_50 (.CK( clk ) , .D( desIn[50] ) , .Q( u0_desIn_r_50 ) );
  DFF_X1 u0_desIn_r_reg_51 (.CK( clk ) , .D( desIn[51] ) , .Q( u0_desIn_r_51 ) );
  DFF_X1 u0_desIn_r_reg_52 (.CK( clk ) , .D( desIn[52] ) , .Q( u0_desIn_r_52 ) );
  DFF_X1 u0_desIn_r_reg_53 (.CK( clk ) , .D( desIn[53] ) , .Q( u0_desIn_r_53 ) );
  DFF_X1 u0_desIn_r_reg_54 (.CK( clk ) , .D( desIn[54] ) , .Q( u0_desIn_r_54 ) );
  DFF_X1 u0_desIn_r_reg_55 (.CK( clk ) , .D( desIn[55] ) , .Q( u0_desIn_r_55 ) );
  DFF_X1 u0_desIn_r_reg_56 (.CK( clk ) , .D( desIn[56] ) , .Q( u0_desIn_r_56 ) );
  DFF_X1 u0_desIn_r_reg_57 (.CK( clk ) , .D( desIn[57] ) , .Q( u0_desIn_r_57 ) );
  DFF_X1 u0_desIn_r_reg_58 (.CK( clk ) , .D( desIn[58] ) , .Q( u0_desIn_r_58 ) );
  DFF_X1 u0_desIn_r_reg_59 (.CK( clk ) , .D( desIn[59] ) , .Q( u0_desIn_r_59 ) );
  DFF_X1 u0_desIn_r_reg_6 (.CK( clk ) , .D( desIn[6] ) , .Q( u0_desIn_r_6 ) );
  DFF_X1 u0_desIn_r_reg_60 (.CK( clk ) , .D( desIn[60] ) , .Q( u0_desIn_r_60 ) );
  DFF_X1 u0_desIn_r_reg_61 (.CK( clk ) , .D( desIn[61] ) , .Q( u0_desIn_r_61 ) );
  DFF_X1 u0_desIn_r_reg_62 (.CK( clk ) , .D( desIn[62] ) , .Q( u0_desIn_r_62 ) );
  DFF_X1 u0_desIn_r_reg_63 (.CK( clk ) , .D( desIn[63] ) , .Q( u0_desIn_r_63 ) );
  DFF_X1 u0_desIn_r_reg_7 (.CK( clk ) , .D( desIn[7] ) , .Q( u0_desIn_r_7 ) );
  DFF_X1 u0_desIn_r_reg_8 (.CK( clk ) , .D( desIn[8] ) , .Q( u0_desIn_r_8 ) );
  DFF_X1 u0_desIn_r_reg_9 (.CK( clk ) , .D( desIn[9] ) , .Q( u0_desIn_r_9 ) );
  DFF_X1 u0_desOut_reg_0 (.CK( clk ) , .Q( stage1_out_0 ) , .D( u0_FP_25 ) );
  DFF_X1 u0_desOut_reg_1 (.CK( clk ) , .Q( stage1_out_1 ) , .D( u0_FP_57 ) );
  DFF_X1 u0_desOut_reg_10 (.CK( clk ) , .Q( stage1_out_10 ) , .D( u0_FP_18 ) );
  DFF_X1 u0_desOut_reg_11 (.CK( clk ) , .Q( stage1_out_11 ) , .D( u0_FP_50 ) );
  DFF_X1 u0_desOut_reg_12 (.CK( clk ) , .Q( stage1_out_12 ) , .D( u0_FP_10 ) );
  DFF_X1 u0_desOut_reg_13 (.CK( clk ) , .Q( stage1_out_13 ) , .D( u0_FP_42 ) );
  DFF_X1 u0_desOut_reg_14 (.CK( clk ) , .Q( stage1_out_14 ) , .D( u0_FP_2 ) );
  DFF_X1 u0_desOut_reg_15 (.CK( clk ) , .Q( stage1_out_15 ) , .D( u0_FP_34 ) );
  DFF_X1 u0_desOut_reg_16 (.CK( clk ) , .Q( stage1_out_16 ) , .D( u0_FP_27 ) );
  DFF_X1 u0_desOut_reg_17 (.CK( clk ) , .Q( stage1_out_17 ) , .D( u0_FP_59 ) );
  DFF_X1 u0_desOut_reg_18 (.CK( clk ) , .Q( stage1_out_18 ) , .D( u0_FP_19 ) );
  DFF_X1 u0_desOut_reg_19 (.CK( clk ) , .Q( stage1_out_19 ) , .D( u0_FP_51 ) );
  DFF_X1 u0_desOut_reg_2 (.CK( clk ) , .Q( stage1_out_2 ) , .D( u0_FP_17 ) );
  DFF_X1 u0_desOut_reg_20 (.CK( clk ) , .Q( stage1_out_20 ) , .D( u0_FP_11 ) );
  DFF_X1 u0_desOut_reg_21 (.CK( clk ) , .Q( stage1_out_21 ) , .D( u0_FP_43 ) );
  DFF_X1 u0_desOut_reg_22 (.CK( clk ) , .Q( stage1_out_22 ) , .D( u0_FP_3 ) );
  DFF_X1 u0_desOut_reg_23 (.CK( clk ) , .Q( stage1_out_23 ) , .D( u0_FP_35 ) );
  DFF_X1 u0_desOut_reg_24 (.CK( clk ) , .Q( stage1_out_24 ) , .D( u0_FP_28 ) );
  DFF_X1 u0_desOut_reg_25 (.CK( clk ) , .Q( stage1_out_25 ) , .D( u0_FP_60 ) );
  DFF_X1 u0_desOut_reg_26 (.CK( clk ) , .Q( stage1_out_26 ) , .D( u0_FP_20 ) );
  DFF_X1 u0_desOut_reg_27 (.CK( clk ) , .Q( stage1_out_27 ) , .D( u0_FP_52 ) );
  DFF_X1 u0_desOut_reg_28 (.CK( clk ) , .Q( stage1_out_28 ) , .D( u0_FP_12 ) );
  DFF_X1 u0_desOut_reg_29 (.CK( clk ) , .Q( stage1_out_29 ) , .D( u0_FP_44 ) );
  DFF_X1 u0_desOut_reg_3 (.CK( clk ) , .Q( stage1_out_3 ) , .D( u0_FP_49 ) );
  DFF_X1 u0_desOut_reg_30 (.CK( clk ) , .Q( stage1_out_30 ) , .D( u0_FP_4 ) );
  DFF_X1 u0_desOut_reg_31 (.CK( clk ) , .Q( stage1_out_31 ) , .D( u0_FP_36 ) );
  DFF_X1 u0_desOut_reg_32 (.CK( clk ) , .Q( stage1_out_32 ) , .D( u0_FP_29 ) );
  DFF_X1 u0_desOut_reg_33 (.CK( clk ) , .Q( stage1_out_33 ) , .D( u0_FP_61 ) );
  DFF_X1 u0_desOut_reg_34 (.CK( clk ) , .Q( stage1_out_34 ) , .D( u0_FP_21 ) );
  DFF_X1 u0_desOut_reg_35 (.CK( clk ) , .Q( stage1_out_35 ) , .D( u0_FP_53 ) );
  DFF_X1 u0_desOut_reg_36 (.CK( clk ) , .Q( stage1_out_36 ) , .D( u0_FP_13 ) );
  DFF_X1 u0_desOut_reg_37 (.CK( clk ) , .Q( stage1_out_37 ) , .D( u0_FP_45 ) );
  DFF_X1 u0_desOut_reg_38 (.CK( clk ) , .Q( stage1_out_38 ) , .D( u0_FP_5 ) );
  DFF_X1 u0_desOut_reg_39 (.CK( clk ) , .Q( stage1_out_39 ) , .D( u0_FP_37 ) );
  DFF_X1 u0_desOut_reg_4 (.CK( clk ) , .Q( stage1_out_4 ) , .D( u0_FP_9 ) );
  DFF_X1 u0_desOut_reg_40 (.CK( clk ) , .Q( stage1_out_40 ) , .D( u0_FP_30 ) );
  DFF_X1 u0_desOut_reg_41 (.CK( clk ) , .Q( stage1_out_41 ) , .D( u0_FP_62 ) );
  DFF_X1 u0_desOut_reg_42 (.CK( clk ) , .Q( stage1_out_42 ) , .D( u0_FP_22 ) );
  DFF_X1 u0_desOut_reg_43 (.CK( clk ) , .Q( stage1_out_43 ) , .D( u0_FP_54 ) );
  DFF_X1 u0_desOut_reg_44 (.CK( clk ) , .Q( stage1_out_44 ) , .D( u0_FP_14 ) );
  DFF_X1 u0_desOut_reg_45 (.CK( clk ) , .Q( stage1_out_45 ) , .D( u0_FP_46 ) );
  DFF_X1 u0_desOut_reg_46 (.CK( clk ) , .Q( stage1_out_46 ) , .D( u0_FP_6 ) );
  DFF_X1 u0_desOut_reg_47 (.CK( clk ) , .Q( stage1_out_47 ) , .D( u0_FP_38 ) );
  DFF_X1 u0_desOut_reg_48 (.CK( clk ) , .Q( stage1_out_48 ) , .D( u0_FP_31 ) );
  DFF_X1 u0_desOut_reg_49 (.CK( clk ) , .Q( stage1_out_49 ) , .D( u0_FP_63 ) );
  DFF_X1 u0_desOut_reg_5 (.CK( clk ) , .Q( stage1_out_5 ) , .D( u0_FP_41 ) );
  DFF_X1 u0_desOut_reg_50 (.CK( clk ) , .Q( stage1_out_50 ) , .D( u0_FP_23 ) );
  DFF_X1 u0_desOut_reg_51 (.CK( clk ) , .Q( stage1_out_51 ) , .D( u0_FP_55 ) );
  DFF_X1 u0_desOut_reg_52 (.CK( clk ) , .Q( stage1_out_52 ) , .D( u0_FP_15 ) );
  DFF_X1 u0_desOut_reg_53 (.CK( clk ) , .Q( stage1_out_53 ) , .D( u0_FP_47 ) );
  DFF_X1 u0_desOut_reg_54 (.CK( clk ) , .Q( stage1_out_54 ) , .D( u0_FP_7 ) );
  DFF_X1 u0_desOut_reg_55 (.CK( clk ) , .Q( stage1_out_55 ) , .D( u0_FP_39 ) );
  DFF_X1 u0_desOut_reg_56 (.CK( clk ) , .Q( stage1_out_56 ) , .D( u0_FP_32 ) );
  DFF_X1 u0_desOut_reg_57 (.CK( clk ) , .Q( stage1_out_57 ) , .D( u0_FP_64 ) );
  DFF_X1 u0_desOut_reg_58 (.CK( clk ) , .Q( stage1_out_58 ) , .D( u0_FP_24 ) );
  DFF_X1 u0_desOut_reg_59 (.CK( clk ) , .Q( stage1_out_59 ) , .D( u0_FP_56 ) );
  DFF_X1 u0_desOut_reg_6 (.CK( clk ) , .Q( stage1_out_6 ) , .D( u0_FP_1 ) );
  DFF_X1 u0_desOut_reg_60 (.CK( clk ) , .Q( stage1_out_60 ) , .D( u0_FP_16 ) );
  DFF_X1 u0_desOut_reg_61 (.CK( clk ) , .Q( stage1_out_61 ) , .D( u0_FP_48 ) );
  DFF_X1 u0_desOut_reg_62 (.CK( clk ) , .Q( stage1_out_62 ) , .D( u0_FP_8 ) );
  DFF_X1 u0_desOut_reg_63 (.CK( clk ) , .Q( stage1_out_63 ) , .D( u0_FP_40 ) );
  DFF_X1 u0_desOut_reg_7 (.CK( clk ) , .Q( stage1_out_7 ) , .D( u0_FP_33 ) );
  DFF_X1 u0_desOut_reg_8 (.CK( clk ) , .Q( stage1_out_8 ) , .D( u0_FP_26 ) );
  DFF_X1 u0_desOut_reg_9 (.CK( clk ) , .Q( stage1_out_9 ) , .D( u0_FP_58 ) );
  DFF_X1 u0_key_r_reg_0 (.CK( clk ) , .D( key_a_0 ) , .Q( u0_key_r_0 ) );
  DFF_X1 u0_key_r_reg_1 (.CK( clk ) , .D( key_a_1 ) , .Q( u0_key_r_1 ) );
  DFF_X1 u0_key_r_reg_10 (.CK( clk ) , .D( key_a_10 ) , .Q( u0_key_r_10 ) );
  DFF_X1 u0_key_r_reg_11 (.CK( clk ) , .D( key_a_11 ) , .Q( u0_key_r_11 ) );
  DFF_X1 u0_key_r_reg_12 (.CK( clk ) , .D( key_a_12 ) , .Q( u0_key_r_12 ) );
  DFF_X1 u0_key_r_reg_13 (.CK( clk ) , .D( key_a_13 ) , .Q( u0_key_r_13 ) );
  DFF_X1 u0_key_r_reg_14 (.CK( clk ) , .D( key_a_14 ) , .Q( u0_key_r_14 ) );
  DFF_X1 u0_key_r_reg_15 (.CK( clk ) , .D( key_a_15 ) , .Q( u0_key_r_15 ) );
  DFF_X1 u0_key_r_reg_16 (.CK( clk ) , .D( key_a_16 ) , .Q( u0_key_r_16 ) );
  DFF_X1 u0_key_r_reg_17 (.CK( clk ) , .D( key_a_17 ) , .Q( u0_key_r_17 ) );
  DFF_X1 u0_key_r_reg_18 (.CK( clk ) , .D( key_a_18 ) , .Q( u0_key_r_18 ) );
  DFF_X1 u0_key_r_reg_19 (.CK( clk ) , .D( key_a_19 ) , .Q( u0_key_r_19 ) );
  DFF_X1 u0_key_r_reg_2 (.CK( clk ) , .D( key_a_2 ) , .Q( u0_key_r_2 ) );
  DFF_X1 u0_key_r_reg_20 (.CK( clk ) , .D( key_a_20 ) , .Q( u0_key_r_20 ) );
  DFF_X1 u0_key_r_reg_21 (.CK( clk ) , .D( key_a_21 ) , .Q( u0_key_r_21 ) );
  DFF_X1 u0_key_r_reg_22 (.CK( clk ) , .D( key_a_22 ) , .Q( u0_key_r_22 ) );
  DFF_X1 u0_key_r_reg_23 (.CK( clk ) , .D( key_a_23 ) , .Q( u0_key_r_23 ) );
  DFF_X1 u0_key_r_reg_24 (.CK( clk ) , .D( key_a_24 ) , .Q( u0_key_r_24 ) );
  DFF_X1 u0_key_r_reg_25 (.CK( clk ) , .D( key_a_25 ) , .Q( u0_key_r_25 ) );
  DFF_X1 u0_key_r_reg_26 (.CK( clk ) , .D( key_a_26 ) , .Q( u0_key_r_26 ) );
  DFF_X1 u0_key_r_reg_27 (.CK( clk ) , .D( key_a_27 ) , .Q( u0_key_r_27 ) );
  DFF_X1 u0_key_r_reg_28 (.CK( clk ) , .D( key_a_28 ) , .Q( u0_key_r_28 ) );
  DFF_X1 u0_key_r_reg_29 (.CK( clk ) , .D( key_a_29 ) , .Q( u0_key_r_29 ) );
  DFF_X1 u0_key_r_reg_3 (.CK( clk ) , .D( key_a_3 ) , .Q( u0_key_r_3 ) );
  DFF_X1 u0_key_r_reg_30 (.CK( clk ) , .D( key_a_30 ) , .Q( u0_key_r_30 ) );
  DFF_X1 u0_key_r_reg_31 (.CK( clk ) , .D( key_a_31 ) , .Q( u0_key_r_31 ) );
  DFF_X1 u0_key_r_reg_32 (.CK( clk ) , .D( key_a_32 ) , .Q( u0_key_r_32 ) );
  DFF_X1 u0_key_r_reg_33 (.CK( clk ) , .D( key_a_33 ) , .Q( u0_key_r_33 ) );
  DFF_X1 u0_key_r_reg_34 (.CK( clk ) , .D( key_a_34 ) , .Q( u0_key_r_34 ) );
  DFF_X1 u0_key_r_reg_35 (.CK( clk ) , .D( key_a_35 ) , .Q( u0_key_r_35 ) );
  DFF_X1 u0_key_r_reg_36 (.CK( clk ) , .D( key_a_36 ) , .Q( u0_key_r_36 ) );
  DFF_X1 u0_key_r_reg_37 (.CK( clk ) , .D( key_a_37 ) , .Q( u0_key_r_37 ) );
  DFF_X1 u0_key_r_reg_38 (.CK( clk ) , .D( key_a_38 ) , .Q( u0_key_r_38 ) );
  DFF_X1 u0_key_r_reg_39 (.CK( clk ) , .D( key_a_39 ) , .Q( u0_key_r_39 ) );
  DFF_X1 u0_key_r_reg_4 (.CK( clk ) , .D( key_a_4 ) , .Q( u0_key_r_4 ) );
  DFF_X1 u0_key_r_reg_40 (.CK( clk ) , .D( key_a_40 ) , .Q( u0_key_r_40 ) );
  DFF_X1 u0_key_r_reg_41 (.CK( clk ) , .D( key_a_41 ) , .Q( u0_key_r_41 ) );
  DFF_X1 u0_key_r_reg_42 (.CK( clk ) , .D( key_a_42 ) , .Q( u0_key_r_42 ) );
  DFF_X1 u0_key_r_reg_43 (.CK( clk ) , .D( key_a_43 ) , .Q( u0_key_r_43 ) );
  DFF_X1 u0_key_r_reg_44 (.CK( clk ) , .D( key_a_44 ) , .Q( u0_key_r_44 ) );
  DFF_X1 u0_key_r_reg_45 (.CK( clk ) , .D( key_a_45 ) , .Q( u0_key_r_45 ) );
  DFF_X1 u0_key_r_reg_46 (.CK( clk ) , .D( key_a_46 ) , .Q( u0_key_r_46 ) );
  DFF_X1 u0_key_r_reg_47 (.CK( clk ) , .D( key_a_47 ) , .Q( u0_key_r_47 ) );
  DFF_X1 u0_key_r_reg_48 (.CK( clk ) , .D( key_a_48 ) , .Q( u0_key_r_48 ) );
  DFF_X1 u0_key_r_reg_49 (.CK( clk ) , .D( key_a_49 ) , .Q( u0_key_r_49 ) );
  DFF_X1 u0_key_r_reg_5 (.CK( clk ) , .D( key_a_5 ) , .Q( u0_key_r_5 ) );
  DFF_X1 u0_key_r_reg_50 (.CK( clk ) , .D( key_a_50 ) , .Q( u0_key_r_50 ) );
  DFF_X1 u0_key_r_reg_51 (.CK( clk ) , .D( key_a_51 ) , .Q( u0_key_r_51 ) );
  DFF_X1 u0_key_r_reg_52 (.CK( clk ) , .D( key_a_52 ) , .Q( u0_key_r_52 ) );
  DFF_X1 u0_key_r_reg_53 (.CK( clk ) , .D( key_a_53 ) , .Q( u0_key_r_53 ) );
  DFF_X1 u0_key_r_reg_54 (.CK( clk ) , .D( key_a_54 ) , .Q( u0_key_r_54 ) );
  DFF_X1 u0_key_r_reg_55 (.CK( clk ) , .D( key_a_55 ) , .Q( u0_key_r_55 ) );
  DFF_X1 u0_key_r_reg_6 (.CK( clk ) , .D( key_a_6 ) , .Q( u0_key_r_6 ) );
  DFF_X1 u0_key_r_reg_7 (.CK( clk ) , .D( key_a_7 ) , .Q( u0_key_r_7 ) );
  DFF_X1 u0_key_r_reg_8 (.CK( clk ) , .D( key_a_8 ) , .Q( u0_key_r_8 ) );
  DFF_X1 u0_key_r_reg_9 (.CK( clk ) , .D( key_a_9 ) , .Q( u0_key_r_9 ) );
  DFF_X1 u0_uk_K_r0_reg_0 (.CK( clk ) , .D( u0_key_r_0 ) , .Q( u0_uk_K_r0_0 ) , .QN( u0_uk_n628 ) );
  DFF_X1 u0_uk_K_r0_reg_1 (.CK( clk ) , .D( u0_key_r_1 ) , .Q( u0_uk_K_r0_1 ) );
  DFF_X1 u0_uk_K_r0_reg_10 (.CK( clk ) , .D( u0_key_r_10 ) , .Q( u0_uk_K_r0_10 ) , .QN( u0_uk_n620 ) );
  DFF_X1 u0_uk_K_r0_reg_11 (.CK( clk ) , .D( u0_key_r_11 ) , .Q( u0_uk_K_r0_11 ) );
  DFF_X1 u0_uk_K_r0_reg_12 (.CK( clk ) , .D( u0_key_r_12 ) , .Q( u0_uk_K_r0_12 ) , .QN( u0_uk_n619 ) );
  DFF_X1 u0_uk_K_r0_reg_13 (.CK( clk ) , .D( u0_key_r_13 ) , .Q( u0_uk_K_r0_13 ) , .QN( u0_uk_n618 ) );
  DFF_X1 u0_uk_K_r0_reg_14 (.CK( clk ) , .D( u0_key_r_14 ) , .Q( u0_uk_K_r0_14 ) , .QN( u0_uk_n617 ) );
  DFF_X1 u0_uk_K_r0_reg_15 (.CK( clk ) , .D( u0_key_r_15 ) , .Q( u0_uk_K_r0_15 ) );
  DFF_X1 u0_uk_K_r0_reg_16 (.CK( clk ) , .D( u0_key_r_16 ) , .Q( u0_uk_K_r0_16 ) , .QN( u0_uk_n616 ) );
  DFF_X1 u0_uk_K_r0_reg_17 (.CK( clk ) , .D( u0_key_r_17 ) , .Q( u0_uk_K_r0_17 ) );
  DFF_X1 u0_uk_K_r0_reg_18 (.CK( clk ) , .D( u0_key_r_18 ) , .Q( u0_uk_K_r0_18 ) , .QN( u0_uk_n615 ) );
  DFF_X1 u0_uk_K_r0_reg_19 (.CK( clk ) , .D( u0_key_r_19 ) , .Q( u0_uk_K_r0_19 ) );
  DFF_X1 u0_uk_K_r0_reg_2 (.CK( clk ) , .D( u0_key_r_2 ) , .Q( u0_uk_K_r0_2 ) );
  DFF_X1 u0_uk_K_r0_reg_20 (.CK( clk ) , .D( u0_key_r_20 ) , .Q( u0_uk_K_r0_20 ) , .QN( u0_uk_n614 ) );
  DFF_X1 u0_uk_K_r0_reg_21 (.CK( clk ) , .D( u0_key_r_21 ) , .Q( u0_uk_K_r0_21 ) , .QN( u0_uk_n613 ) );
  DFF_X1 u0_uk_K_r0_reg_22 (.CK( clk ) , .D( u0_key_r_22 ) , .Q( u0_uk_K_r0_22 ) );
  DFF_X1 u0_uk_K_r0_reg_23 (.CK( clk ) , .D( u0_key_r_23 ) , .Q( u0_uk_K_r0_23 ) , .QN( u0_uk_n612 ) );
  DFF_X1 u0_uk_K_r0_reg_24 (.CK( clk ) , .D( u0_key_r_24 ) , .Q( u0_uk_K_r0_24 ) , .QN( u0_uk_n611 ) );
  DFF_X1 u0_uk_K_r0_reg_25 (.CK( clk ) , .D( u0_key_r_25 ) , .Q( u0_uk_K_r0_25 ) );
  DFF_X1 u0_uk_K_r0_reg_26 (.CK( clk ) , .D( u0_key_r_26 ) , .Q( u0_uk_K_r0_26 ) , .QN( u0_uk_n610 ) );
  DFF_X1 u0_uk_K_r0_reg_27 (.CK( clk ) , .D( u0_key_r_27 ) , .Q( u0_uk_K_r0_27 ) , .QN( u0_uk_n609 ) );
  DFF_X1 u0_uk_K_r0_reg_28 (.CK( clk ) , .D( u0_key_r_28 ) , .Q( u0_uk_K_r0_28 ) );
  DFF_X1 u0_uk_K_r0_reg_29 (.CK( clk ) , .D( u0_key_r_29 ) , .Q( u0_uk_K_r0_29 ) , .QN( u0_uk_n607 ) );
  DFF_X1 u0_uk_K_r0_reg_3 (.CK( clk ) , .D( u0_key_r_3 ) , .Q( u0_uk_K_r0_3 ) , .QN( u0_uk_n627 ) );
  DFF_X1 u0_uk_K_r0_reg_30 (.CK( clk ) , .D( u0_key_r_30 ) , .Q( u0_uk_K_r0_30 ) , .QN( u0_uk_n606 ) );
  DFF_X1 u0_uk_K_r0_reg_31 (.CK( clk ) , .D( u0_key_r_31 ) , .Q( u0_uk_K_r0_31 ) );
  DFF_X1 u0_uk_K_r0_reg_32 (.CK( clk ) , .D( u0_key_r_32 ) , .Q( u0_uk_K_r0_32 ) );
  DFF_X1 u0_uk_K_r0_reg_33 (.CK( clk ) , .D( u0_key_r_33 ) , .Q( u0_uk_K_r0_33 ) , .QN( u0_uk_n604 ) );
  DFF_X1 u0_uk_K_r0_reg_34 (.CK( clk ) , .D( u0_key_r_34 ) , .Q( u0_uk_K_r0_34 ) );
  DFF_X1 u0_uk_K_r0_reg_35 (.CK( clk ) , .D( u0_key_r_35 ) , .Q( u0_uk_K_r0_35 ) , .QN( u0_uk_n602 ) );
  DFF_X1 u0_uk_K_r0_reg_36 (.CK( clk ) , .D( u0_key_r_36 ) , .Q( u0_uk_K_r0_36 ) );
  DFF_X1 u0_uk_K_r0_reg_37 (.CK( clk ) , .D( u0_key_r_37 ) , .Q( u0_uk_K_r0_37 ) , .QN( u0_uk_n600 ) );
  DFF_X1 u0_uk_K_r0_reg_38 (.CK( clk ) , .D( u0_key_r_38 ) , .Q( u0_uk_K_r0_38 ) , .QN( u0_uk_n599 ) );
  DFF_X1 u0_uk_K_r0_reg_39 (.CK( clk ) , .D( u0_key_r_39 ) , .Q( u0_uk_K_r0_39 ) , .QN( u0_uk_n598 ) );
  DFF_X1 u0_uk_K_r0_reg_4 (.CK( clk ) , .D( u0_key_r_4 ) , .Q( u0_uk_K_r0_4 ) , .QN( u0_uk_n626 ) );
  DFF_X1 u0_uk_K_r0_reg_40 (.CK( clk ) , .D( u0_key_r_40 ) , .Q( u0_uk_K_r0_40 ) , .QN( u0_uk_n597 ) );
  DFF_X1 u0_uk_K_r0_reg_41 (.CK( clk ) , .D( u0_key_r_41 ) , .Q( u0_uk_K_r0_41 ) , .QN( u0_uk_n596 ) );
  DFF_X1 u0_uk_K_r0_reg_42 (.CK( clk ) , .D( u0_key_r_42 ) , .Q( u0_uk_K_r0_42 ) , .QN( u0_uk_n595 ) );
  DFF_X1 u0_uk_K_r0_reg_43 (.CK( clk ) , .D( u0_key_r_43 ) , .Q( u0_uk_K_r0_43 ) , .QN( u0_uk_n594 ) );
  DFF_X1 u0_uk_K_r0_reg_44 (.CK( clk ) , .D( u0_key_r_44 ) , .Q( u0_uk_K_r0_44 ) , .QN( u0_uk_n593 ) );
  DFF_X1 u0_uk_K_r0_reg_45 (.CK( clk ) , .D( u0_key_r_45 ) , .Q( u0_uk_K_r0_45 ) , .QN( u0_uk_n592 ) );
  DFF_X1 u0_uk_K_r0_reg_46 (.CK( clk ) , .D( u0_key_r_46 ) , .Q( u0_uk_K_r0_46 ) , .QN( u0_uk_n591 ) );
  DFF_X1 u0_uk_K_r0_reg_47 (.CK( clk ) , .D( u0_key_r_47 ) , .Q( u0_uk_K_r0_47 ) , .QN( u0_uk_n589 ) );
  DFF_X1 u0_uk_K_r0_reg_48 (.CK( clk ) , .D( u0_key_r_48 ) , .Q( u0_uk_K_r0_48 ) , .QN( u0_uk_n588 ) );
  DFF_X1 u0_uk_K_r0_reg_49 (.CK( clk ) , .D( u0_key_r_49 ) , .Q( u0_uk_K_r0_49 ) );
  DFF_X1 u0_uk_K_r0_reg_5 (.CK( clk ) , .D( u0_key_r_5 ) , .Q( u0_uk_K_r0_5 ) , .QN( u0_uk_n625 ) );
  DFF_X1 u0_uk_K_r0_reg_50 (.CK( clk ) , .D( u0_key_r_50 ) , .Q( u0_uk_K_r0_50 ) , .QN( u0_uk_n585 ) );
  DFF_X1 u0_uk_K_r0_reg_51 (.CK( clk ) , .D( u0_key_r_51 ) , .Q( u0_uk_K_r0_51 ) , .QN( u0_uk_n584 ) );
  DFF_X1 u0_uk_K_r0_reg_52 (.CK( clk ) , .D( u0_key_r_52 ) , .Q( u0_uk_K_r0_52 ) );
  DFF_X1 u0_uk_K_r0_reg_53 (.CK( clk ) , .D( u0_key_r_53 ) , .Q( u0_uk_K_r0_53 ) );
  DFF_X1 u0_uk_K_r0_reg_54 (.CK( clk ) , .D( u0_key_r_54 ) , .Q( u0_uk_K_r0_54 ) , .QN( u0_uk_n583 ) );
  DFF_X1 u0_uk_K_r0_reg_55 (.CK( clk ) , .D( u0_key_r_55 ) , .Q( u0_uk_K_r0_55 ) );
  DFF_X1 u0_uk_K_r0_reg_6 (.CK( clk ) , .D( u0_key_r_6 ) , .Q( u0_uk_K_r0_6 ) , .QN( u0_uk_n624 ) );
  DFF_X1 u0_uk_K_r0_reg_7 (.CK( clk ) , .D( u0_key_r_7 ) , .Q( u0_uk_K_r0_7 ) , .QN( u0_uk_n623 ) );
  DFF_X1 u0_uk_K_r0_reg_8 (.CK( clk ) , .D( u0_key_r_8 ) , .Q( u0_uk_K_r0_8 ) , .QN( u0_uk_n622 ) );
  DFF_X1 u0_uk_K_r0_reg_9 (.CK( clk ) , .D( u0_key_r_9 ) , .Q( u0_uk_K_r0_9 ) , .QN( u0_uk_n621 ) );
  DFF_X1 u0_uk_K_r10_reg_0 (.CK( clk ) , .Q( u0_uk_K_r10_0 ) , .D( u0_uk_K_r9_0 ) , .QN( u0_uk_n180 ) );
  DFF_X1 u0_uk_K_r10_reg_1 (.CK( clk ) , .Q( u0_uk_K_r10_1 ) , .D( u0_uk_K_r9_1 ) , .QN( u0_uk_n179 ) );
  DFF_X1 u0_uk_K_r10_reg_10 (.CK( clk ) , .Q( u0_uk_K_r10_10 ) , .D( u0_uk_K_r9_10 ) );
  DFF_X1 u0_uk_K_r10_reg_11 (.CK( clk ) , .Q( u0_uk_K_r10_11 ) , .D( u0_uk_K_r9_11 ) );
  DFF_X1 u0_uk_K_r10_reg_12 (.CK( clk ) , .Q( u0_uk_K_r10_12 ) , .D( u0_uk_K_r9_12 ) , .QN( u0_uk_n172 ) );
  DFF_X1 u0_uk_K_r10_reg_13 (.CK( clk ) , .Q( u0_uk_K_r10_13 ) , .D( u0_uk_K_r9_13 ) );
  DFF_X1 u0_uk_K_r10_reg_14 (.CK( clk ) , .Q( u0_uk_K_r10_14 ) , .D( u0_uk_K_r9_14 ) );
  DFF_X1 u0_uk_K_r10_reg_15 (.CK( clk ) , .Q( u0_uk_K_r10_15 ) , .D( u0_uk_K_r9_15 ) , .QN( u0_uk_n171 ) );
  DFF_X1 u0_uk_K_r10_reg_16 (.CK( clk ) , .Q( u0_uk_K_r10_16 ) , .D( u0_uk_K_r9_16 ) );
  DFF_X1 u0_uk_K_r10_reg_17 (.CK( clk ) , .Q( u0_uk_K_r10_17 ) , .D( u0_uk_K_r9_17 ) , .QN( u0_uk_n170 ) );
  DFF_X1 u0_uk_K_r10_reg_18 (.CK( clk ) , .Q( u0_uk_K_r10_18 ) , .D( u0_uk_K_r9_18 ) );
  DFF_X1 u0_uk_K_r10_reg_19 (.CK( clk ) , .Q( u0_uk_K_r10_19 ) , .D( u0_uk_K_r9_19 ) );
  DFF_X1 u0_uk_K_r10_reg_2 (.CK( clk ) , .Q( u0_uk_K_r10_2 ) , .D( u0_uk_K_r9_2 ) , .QN( u0_uk_n178 ) );
  DFF_X1 u0_uk_K_r10_reg_20 (.CK( clk ) , .Q( u0_uk_K_r10_20 ) , .D( u0_uk_K_r9_20 ) , .QN( u0_uk_n169 ) );
  DFF_X1 u0_uk_K_r10_reg_21 (.CK( clk ) , .Q( u0_uk_K_r10_21 ) , .D( u0_uk_K_r9_21 ) , .QN( u0_uk_n168 ) );
  DFF_X1 u0_uk_K_r10_reg_22 (.CK( clk ) , .Q( u0_uk_K_r10_22 ) , .D( u0_uk_K_r9_22 ) , .QN( u0_uk_n167 ) );
  DFF_X1 u0_uk_K_r10_reg_23 (.CK( clk ) , .Q( u0_uk_K_r10_23 ) , .D( u0_uk_K_r9_23 ) );
  DFF_X1 u0_uk_K_r10_reg_24 (.CK( clk ) , .Q( u0_uk_K_r10_24 ) , .D( u0_uk_K_r9_24 ) , .QN( u0_uk_n166 ) );
  DFF_X1 u0_uk_K_r10_reg_25 (.CK( clk ) , .Q( u0_uk_K_r10_25 ) , .D( u0_uk_K_r9_25 ) );
  DFF_X1 u0_uk_K_r10_reg_26 (.CK( clk ) , .Q( u0_uk_K_r10_26 ) , .D( u0_uk_K_r9_26 ) , .QN( u0_uk_n165 ) );
  DFF_X1 u0_uk_K_r10_reg_27 (.CK( clk ) , .Q( u0_uk_K_r10_27 ) , .D( u0_uk_K_r9_27 ) );
  DFF_X1 u0_uk_K_r10_reg_28 (.CK( clk ) , .Q( u0_uk_K_r10_28 ) , .D( u0_uk_K_r9_28 ) );
  DFF_X1 u0_uk_K_r10_reg_29 (.CK( clk ) , .Q( u0_uk_K_r10_29 ) , .D( u0_uk_K_r9_29 ) , .QN( u0_uk_n160 ) );
  DFF_X1 u0_uk_K_r10_reg_3 (.CK( clk ) , .Q( u0_uk_K_r10_3 ) , .D( u0_uk_K_r9_3 ) , .QN( u0_uk_n177 ) );
  DFF_X1 u0_uk_K_r10_reg_30 (.CK( clk ) , .Q( u0_uk_K_r10_30 ) , .D( u0_uk_K_r9_30 ) , .QN( u0_uk_n159 ) );
  DFF_X1 u0_uk_K_r10_reg_31 (.CK( clk ) , .Q( u0_uk_K_r10_31 ) , .D( u0_uk_K_r9_31 ) , .QN( u0_uk_n158 ) );
  DFF_X1 u0_uk_K_r10_reg_32 (.CK( clk ) , .Q( u0_uk_K_r10_32 ) , .D( u0_uk_K_r9_32 ) , .QN( u0_uk_n157 ) );
  DFF_X1 u0_uk_K_r10_reg_33 (.CK( clk ) , .Q( u0_uk_K_r10_33 ) , .D( u0_uk_K_r9_33 ) , .QN( u0_uk_n156 ) );
  DFF_X1 u0_uk_K_r10_reg_34 (.CK( clk ) , .Q( u0_uk_K_r10_34 ) , .D( u0_uk_K_r9_34 ) );
  DFF_X1 u0_uk_K_r10_reg_35 (.CK( clk ) , .Q( u0_uk_K_r10_35 ) , .D( u0_uk_K_r9_35 ) , .QN( u0_uk_n154 ) );
  DFF_X1 u0_uk_K_r10_reg_36 (.CK( clk ) , .Q( u0_uk_K_r10_36 ) , .D( u0_uk_K_r9_36 ) , .QN( u0_uk_n153 ) );
  DFF_X1 u0_uk_K_r10_reg_37 (.CK( clk ) , .Q( u0_uk_K_r10_37 ) , .D( u0_uk_K_r9_37 ) , .QN( u0_uk_n152 ) );
  DFF_X1 u0_uk_K_r10_reg_38 (.CK( clk ) , .Q( u0_uk_K_r10_38 ) , .D( u0_uk_K_r9_38 ) , .QN( u0_uk_n151 ) );
  DFF_X1 u0_uk_K_r10_reg_39 (.CK( clk ) , .Q( u0_uk_K_r10_39 ) , .D( u0_uk_K_r9_39 ) , .QN( u0_uk_n150 ) );
  DFF_X1 u0_uk_K_r10_reg_4 (.CK( clk ) , .Q( u0_uk_K_r10_4 ) , .D( u0_uk_K_r9_4 ) );
  DFF_X1 u0_uk_K_r10_reg_40 (.CK( clk ) , .Q( u0_uk_K_r10_40 ) , .D( u0_uk_K_r9_40 ) , .QN( u0_uk_n149 ) );
  DFF_X1 u0_uk_K_r10_reg_41 (.CK( clk ) , .Q( u0_uk_K_r10_41 ) , .D( u0_uk_K_r9_41 ) );
  DFF_X1 u0_uk_K_r10_reg_42 (.CK( clk ) , .Q( u0_uk_K_r10_42 ) , .D( u0_uk_K_r9_42 ) );
  DFF_X1 u0_uk_K_r10_reg_43 (.CK( clk ) , .Q( u0_uk_K_r10_43 ) , .D( u0_uk_K_r9_43 ) );
  DFF_X1 u0_uk_K_r10_reg_44 (.CK( clk ) , .Q( u0_uk_K_r10_44 ) , .D( u0_uk_K_r9_44 ) );
  DFF_X1 u0_uk_K_r10_reg_45 (.CK( clk ) , .Q( u0_uk_K_r10_45 ) , .D( u0_uk_K_r9_45 ) , .QN( u0_uk_n144 ) );
  DFF_X1 u0_uk_K_r10_reg_46 (.CK( clk ) , .Q( u0_uk_K_r10_46 ) , .D( u0_uk_K_r9_46 ) , .QN( u0_uk_n143 ) );
  DFF_X1 u0_uk_K_r10_reg_47 (.CK( clk ) , .Q( u0_uk_K_r10_47 ) , .D( u0_uk_K_r9_47 ) );
  DFF_X1 u0_uk_K_r10_reg_48 (.CK( clk ) , .Q( u0_uk_K_r10_48 ) , .D( u0_uk_K_r9_48 ) );
  DFF_X1 u0_uk_K_r10_reg_49 (.CK( clk ) , .Q( u0_uk_K_r10_49 ) , .D( u0_uk_K_r9_49 ) );
  DFF_X1 u0_uk_K_r10_reg_5 (.CK( clk ) , .Q( u0_uk_K_r10_5 ) , .D( u0_uk_K_r9_5 ) , .QN( u0_uk_n176 ) );
  DFF_X1 u0_uk_K_r10_reg_50 (.CK( clk ) , .Q( u0_uk_K_r10_50 ) , .D( u0_uk_K_r9_50 ) , .QN( u0_uk_n140 ) );
  DFF_X1 u0_uk_K_r10_reg_51 (.CK( clk ) , .Q( u0_uk_K_r10_51 ) , .D( u0_uk_K_r9_51 ) , .QN( u0_uk_n139 ) );
  DFF_X1 u0_uk_K_r10_reg_52 (.CK( clk ) , .Q( u0_uk_K_r10_52 ) , .D( u0_uk_K_r9_52 ) );
  DFF_X1 u0_uk_K_r10_reg_53 (.CK( clk ) , .Q( u0_uk_K_r10_53 ) , .D( u0_uk_K_r9_53 ) , .QN( u0_uk_n138 ) );
  DFF_X1 u0_uk_K_r10_reg_54 (.CK( clk ) , .Q( u0_uk_K_r10_54 ) , .D( u0_uk_K_r9_54 ) , .QN( u0_uk_n137 ) );
  DFF_X1 u0_uk_K_r10_reg_55 (.CK( clk ) , .Q( u0_uk_K_r10_55 ) , .D( u0_uk_K_r9_55 ) , .QN( u0_uk_n136 ) );
  DFF_X1 u0_uk_K_r10_reg_6 (.CK( clk ) , .Q( u0_uk_K_r10_6 ) , .D( u0_uk_K_r9_6 ) , .QN( u0_uk_n175 ) );
  DFF_X1 u0_uk_K_r10_reg_7 (.CK( clk ) , .Q( u0_uk_K_r10_7 ) , .D( u0_uk_K_r9_7 ) , .QN( u0_uk_n174 ) );
  DFF_X1 u0_uk_K_r10_reg_8 (.CK( clk ) , .Q( u0_uk_K_r10_8 ) , .D( u0_uk_K_r9_8 ) , .QN( u0_uk_n173 ) );
  DFF_X1 u0_uk_K_r10_reg_9 (.CK( clk ) , .Q( u0_uk_K_r10_9 ) , .D( u0_uk_K_r9_9 ) );
  DFF_X1 u0_uk_K_r11_reg_0 (.CK( clk ) , .D( u0_uk_K_r10_0 ) , .Q( u0_uk_K_r11_0 ) , .QN( u0_uk_n135 ) );
  DFF_X1 u0_uk_K_r11_reg_1 (.CK( clk ) , .D( u0_uk_K_r10_1 ) , .Q( u0_uk_K_r11_1 ) , .QN( u0_uk_n134 ) );
  DFF_X1 u0_uk_K_r11_reg_10 (.CK( clk ) , .D( u0_uk_K_r10_10 ) , .Q( u0_uk_K_r11_10 ) );
  DFF_X1 u0_uk_K_r11_reg_11 (.CK( clk ) , .D( u0_uk_K_r10_11 ) , .Q( u0_uk_K_r11_11 ) );
  DFF_X1 u0_uk_K_r11_reg_12 (.CK( clk ) , .D( u0_uk_K_r10_12 ) , .Q( u0_uk_K_r11_12 ) , .QN( u0_uk_n127 ) );
  DFF_X1 u0_uk_K_r11_reg_13 (.CK( clk ) , .D( u0_uk_K_r10_13 ) , .Q( u0_uk_K_r11_13 ) , .QN( u0_uk_n126 ) );
  DFF_X1 u0_uk_K_r11_reg_14 (.CK( clk ) , .D( u0_uk_K_r10_14 ) , .Q( u0_uk_K_r11_14 ) , .QN( u0_uk_n125 ) );
  DFF_X1 u0_uk_K_r11_reg_15 (.CK( clk ) , .D( u0_uk_K_r10_15 ) , .Q( u0_uk_K_r11_15 ) , .QN( u0_uk_n124 ) );
  DFF_X1 u0_uk_K_r11_reg_16 (.CK( clk ) , .D( u0_uk_K_r10_16 ) , .Q( u0_uk_K_r11_16 ) , .QN( u0_uk_n123 ) );
  DFF_X1 u0_uk_K_r11_reg_17 (.CK( clk ) , .D( u0_uk_K_r10_17 ) , .Q( u0_uk_K_r11_17 ) , .QN( u0_uk_n122 ) );
  DFF_X1 u0_uk_K_r11_reg_18 (.CK( clk ) , .D( u0_uk_K_r10_18 ) , .Q( u0_uk_K_r11_18 ) , .QN( u0_uk_n121 ) );
  DFF_X1 u0_uk_K_r11_reg_19 (.CK( clk ) , .D( u0_uk_K_r10_19 ) , .Q( u0_uk_K_r11_19 ) );
  DFF_X1 u0_uk_K_r11_reg_2 (.CK( clk ) , .D( u0_uk_K_r10_2 ) , .Q( u0_uk_K_r11_2 ) , .QN( u0_uk_n133 ) );
  DFF_X1 u0_uk_K_r11_reg_20 (.CK( clk ) , .D( u0_uk_K_r10_20 ) , .Q( u0_uk_K_r11_20 ) );
  DFF_X1 u0_uk_K_r11_reg_21 (.CK( clk ) , .D( u0_uk_K_r10_21 ) , .Q( u0_uk_K_r11_21 ) );
  DFF_X1 u0_uk_K_r11_reg_22 (.CK( clk ) , .D( u0_uk_K_r10_22 ) , .Q( u0_uk_K_r11_22 ) , .QN( u0_uk_n120 ) );
  DFF_X1 u0_uk_K_r11_reg_23 (.CK( clk ) , .D( u0_uk_K_r10_23 ) , .Q( u0_uk_K_r11_23 ) , .QN( u0_uk_n119 ) );
  DFF_X1 u0_uk_K_r11_reg_24 (.CK( clk ) , .D( u0_uk_K_r10_24 ) , .Q( u0_uk_K_r11_24 ) );
  DFF_X1 u0_uk_K_r11_reg_25 (.CK( clk ) , .D( u0_uk_K_r10_25 ) , .Q( u0_uk_K_r11_25 ) );
  DFF_X1 u0_uk_K_r11_reg_26 (.CK( clk ) , .D( u0_uk_K_r10_26 ) , .Q( u0_uk_K_r11_26 ) );
  DFF_X1 u0_uk_K_r11_reg_27 (.CK( clk ) , .D( u0_uk_K_r10_27 ) , .Q( u0_uk_K_r11_27 ) );
  DFF_X1 u0_uk_K_r11_reg_28 (.CK( clk ) , .D( u0_uk_K_r10_28 ) , .Q( u0_uk_K_r11_28 ) );
  DFF_X1 u0_uk_K_r11_reg_29 (.CK( clk ) , .D( u0_uk_K_r10_29 ) , .Q( u0_uk_K_r11_29 ) );
  DFF_X1 u0_uk_K_r11_reg_3 (.CK( clk ) , .D( u0_uk_K_r10_3 ) , .Q( u0_uk_K_r11_3 ) , .QN( u0_uk_n132 ) );
  DFF_X1 u0_uk_K_r11_reg_30 (.CK( clk ) , .D( u0_uk_K_r10_30 ) , .Q( u0_uk_K_r11_30 ) );
  DFF_X1 u0_uk_K_r11_reg_31 (.CK( clk ) , .D( u0_uk_K_r10_31 ) , .Q( u0_uk_K_r11_31 ) , .QN( u0_uk_n116 ) );
  DFF_X1 u0_uk_K_r11_reg_32 (.CK( clk ) , .D( u0_uk_K_r10_32 ) , .Q( u0_uk_K_r11_32 ) , .QN( u0_uk_n115 ) );
  DFF_X1 u0_uk_K_r11_reg_33 (.CK( clk ) , .D( u0_uk_K_r10_33 ) , .Q( u0_uk_K_r11_33 ) );
  DFF_X1 u0_uk_K_r11_reg_34 (.CK( clk ) , .D( u0_uk_K_r10_34 ) , .Q( u0_uk_K_r11_34 ) );
  DFF_X1 u0_uk_K_r11_reg_35 (.CK( clk ) , .D( u0_uk_K_r10_35 ) , .Q( u0_uk_K_r11_35 ) , .QN( u0_uk_n114 ) );
  DFF_X1 u0_uk_K_r11_reg_36 (.CK( clk ) , .D( u0_uk_K_r10_36 ) , .Q( u0_uk_K_r11_36 ) , .QN( u0_uk_n113 ) );
  DFF_X1 u0_uk_K_r11_reg_37 (.CK( clk ) , .D( u0_uk_K_r10_37 ) , .Q( u0_uk_K_r11_37 ) , .QN( u0_uk_n112 ) );
  DFF_X1 u0_uk_K_r11_reg_38 (.CK( clk ) , .D( u0_uk_K_r10_38 ) , .Q( u0_uk_K_r11_38 ) , .QN( u0_uk_n111 ) );
  DFF_X1 u0_uk_K_r11_reg_39 (.CK( clk ) , .D( u0_uk_K_r10_39 ) , .Q( u0_uk_K_r11_39 ) );
  DFF_X1 u0_uk_K_r11_reg_4 (.CK( clk ) , .D( u0_uk_K_r10_4 ) , .Q( u0_uk_K_r11_4 ) );
  DFF_X1 u0_uk_K_r11_reg_40 (.CK( clk ) , .D( u0_uk_K_r10_40 ) , .Q( u0_uk_K_r11_40 ) , .QN( u0_uk_n108 ) );
  DFF_X1 u0_uk_K_r11_reg_41 (.CK( clk ) , .D( u0_uk_K_r10_41 ) , .Q( u0_uk_K_r11_41 ) , .QN( u0_uk_n107 ) );
  DFF_X1 u0_uk_K_r11_reg_42 (.CK( clk ) , .D( u0_uk_K_r10_42 ) , .Q( u0_uk_K_r11_42 ) , .QN( u0_uk_n106 ) );
  DFF_X1 u0_uk_K_r11_reg_43 (.CK( clk ) , .D( u0_uk_K_r10_43 ) , .Q( u0_uk_K_r11_43 ) , .QN( u0_uk_n105 ) );
  DFF_X1 u0_uk_K_r11_reg_44 (.CK( clk ) , .D( u0_uk_K_r10_44 ) , .Q( u0_uk_K_r11_44 ) , .QN( u0_uk_n104 ) );
  DFF_X1 u0_uk_K_r11_reg_45 (.CK( clk ) , .D( u0_uk_K_r10_45 ) , .Q( u0_uk_K_r11_45 ) , .QN( u0_uk_n103 ) );
  DFF_X1 u0_uk_K_r11_reg_46 (.CK( clk ) , .D( u0_uk_K_r10_46 ) , .Q( u0_uk_K_r11_46 ) , .QN( u0_uk_n101 ) );
  DFF_X1 u0_uk_K_r11_reg_47 (.CK( clk ) , .D( u0_uk_K_r10_47 ) , .Q( u0_uk_K_r11_47 ) );
  DFF_X1 u0_uk_K_r11_reg_48 (.CK( clk ) , .D( u0_uk_K_r10_48 ) , .Q( u0_uk_K_r11_48 ) );
  DFF_X1 u0_uk_K_r11_reg_49 (.CK( clk ) , .D( u0_uk_K_r10_49 ) , .Q( u0_uk_K_r11_49 ) , .QN( u0_uk_n98 ) );
  DFF_X1 u0_uk_K_r11_reg_5 (.CK( clk ) , .D( u0_uk_K_r10_5 ) , .Q( u0_uk_K_r11_5 ) , .QN( u0_uk_n131 ) );
  DFF_X1 u0_uk_K_r11_reg_50 (.CK( clk ) , .D( u0_uk_K_r10_50 ) , .Q( u0_uk_K_r11_50 ) , .QN( u0_uk_n97 ) );
  DFF_X1 u0_uk_K_r11_reg_51 (.CK( clk ) , .D( u0_uk_K_r10_51 ) , .Q( u0_uk_K_r11_51 ) , .QN( u0_uk_n96 ) );
  DFF_X1 u0_uk_K_r11_reg_52 (.CK( clk ) , .D( u0_uk_K_r10_52 ) , .Q( u0_uk_K_r11_52 ) , .QN( u0_uk_n95 ) );
  DFF_X1 u0_uk_K_r11_reg_53 (.CK( clk ) , .D( u0_uk_K_r10_53 ) , .Q( u0_uk_K_r11_53 ) );
  DFF_X1 u0_uk_K_r11_reg_54 (.CK( clk ) , .D( u0_uk_K_r10_54 ) , .Q( u0_uk_K_r11_54 ) );
  DFF_X1 u0_uk_K_r11_reg_55 (.CK( clk ) , .D( u0_uk_K_r10_55 ) , .Q( u0_uk_K_r11_55 ) , .QN( u0_uk_n91 ) );
  DFF_X1 u0_uk_K_r11_reg_6 (.CK( clk ) , .D( u0_uk_K_r10_6 ) , .Q( u0_uk_K_r11_6 ) );
  DFF_X1 u0_uk_K_r11_reg_7 (.CK( clk ) , .D( u0_uk_K_r10_7 ) , .Q( u0_uk_K_r11_7 ) );
  DFF_X1 u0_uk_K_r11_reg_8 (.CK( clk ) , .D( u0_uk_K_r10_8 ) , .Q( u0_uk_K_r11_8 ) );
  DFF_X1 u0_uk_K_r11_reg_9 (.CK( clk ) , .D( u0_uk_K_r10_9 ) , .Q( u0_uk_K_r11_9 ) , .QN( u0_uk_n130 ) );
  DFF_X1 u0_uk_K_r12_reg_0 (.CK( clk ) , .D( u0_uk_K_r11_0 ) , .Q( u0_uk_K_r12_0 ) , .QN( u0_uk_n90 ) );
  DFF_X1 u0_uk_K_r12_reg_1 (.CK( clk ) , .D( u0_uk_K_r11_1 ) , .Q( u0_uk_K_r12_1 ) , .QN( u0_uk_n89 ) );
  DFF_X1 u0_uk_K_r12_reg_10 (.CK( clk ) , .D( u0_uk_K_r11_10 ) , .Q( u0_uk_K_r12_10 ) );
  DFF_X1 u0_uk_K_r12_reg_11 (.CK( clk ) , .D( u0_uk_K_r11_11 ) , .Q( u0_uk_K_r12_11 ) , .QN( u0_uk_n80 ) );
  DFF_X1 u0_uk_K_r12_reg_12 (.CK( clk ) , .D( u0_uk_K_r11_12 ) , .Q( u0_uk_K_r12_12 ) , .QN( u0_uk_n79 ) );
  DFF_X1 u0_uk_K_r12_reg_13 (.CK( clk ) , .D( u0_uk_K_r11_13 ) , .Q( u0_uk_K_r12_13 ) , .QN( u0_uk_n78 ) );
  DFF_X1 u0_uk_K_r12_reg_14 (.CK( clk ) , .D( u0_uk_K_r11_14 ) , .Q( u0_uk_K_r12_14 ) , .QN( u0_uk_n77 ) );
  DFF_X1 u0_uk_K_r12_reg_15 (.CK( clk ) , .D( u0_uk_K_r11_15 ) , .Q( u0_uk_K_r12_15 ) );
  DFF_X1 u0_uk_K_r12_reg_16 (.CK( clk ) , .D( u0_uk_K_r11_16 ) , .Q( u0_uk_K_r12_16 ) );
  DFF_X1 u0_uk_K_r12_reg_17 (.CK( clk ) , .D( u0_uk_K_r11_17 ) , .Q( u0_uk_K_r12_17 ) , .QN( u0_uk_n76 ) );
  DFF_X1 u0_uk_K_r12_reg_18 (.CK( clk ) , .D( u0_uk_K_r11_18 ) , .Q( u0_uk_K_r12_18 ) );
  DFF_X1 u0_uk_K_r12_reg_19 (.CK( clk ) , .D( u0_uk_K_r11_19 ) , .Q( u0_uk_K_r12_19 ) , .QN( u0_uk_n75 ) );
  DFF_X1 u0_uk_K_r12_reg_2 (.CK( clk ) , .D( u0_uk_K_r11_2 ) , .Q( u0_uk_K_r12_2 ) , .QN( u0_uk_n88 ) );
  DFF_X1 u0_uk_K_r12_reg_20 (.CK( clk ) , .D( u0_uk_K_r11_20 ) , .Q( u0_uk_K_r12_20 ) , .QN( u0_uk_n74 ) );
  DFF_X1 u0_uk_K_r12_reg_21 (.CK( clk ) , .D( u0_uk_K_r11_21 ) , .Q( u0_uk_K_r12_21 ) );
  DFF_X1 u0_uk_K_r12_reg_22 (.CK( clk ) , .D( u0_uk_K_r11_22 ) , .Q( u0_uk_K_r12_22 ) );
  DFF_X1 u0_uk_K_r12_reg_23 (.CK( clk ) , .D( u0_uk_K_r11_23 ) , .Q( u0_uk_K_r12_23 ) , .QN( u0_uk_n73 ) );
  DFF_X1 u0_uk_K_r12_reg_24 (.CK( clk ) , .D( u0_uk_K_r11_24 ) , .Q( u0_uk_K_r12_24 ) , .QN( u0_uk_n72 ) );
  DFF_X1 u0_uk_K_r12_reg_25 (.CK( clk ) , .D( u0_uk_K_r11_25 ) , .Q( u0_uk_K_r12_25 ) , .QN( u0_uk_n71 ) );
  DFF_X1 u0_uk_K_r12_reg_26 (.CK( clk ) , .D( u0_uk_K_r11_26 ) , .Q( u0_uk_K_r12_26 ) , .QN( u0_uk_n70 ) );
  DFF_X1 u0_uk_K_r12_reg_27 (.CK( clk ) , .D( u0_uk_K_r11_27 ) , .Q( u0_uk_K_r12_27 ) , .QN( u0_uk_n69 ) );
  DFF_X1 u0_uk_K_r12_reg_28 (.CK( clk ) , .D( u0_uk_K_r11_28 ) , .Q( u0_uk_K_r12_28 ) , .QN( u0_uk_n68 ) );
  DFF_X1 u0_uk_K_r12_reg_29 (.CK( clk ) , .D( u0_uk_K_r11_29 ) , .Q( u0_uk_K_r12_29 ) , .QN( u0_uk_n67 ) );
  DFF_X1 u0_uk_K_r12_reg_3 (.CK( clk ) , .D( u0_uk_K_r11_3 ) , .Q( u0_uk_K_r12_3 ) , .QN( u0_uk_n87 ) );
  DFF_X1 u0_uk_K_r12_reg_30 (.CK( clk ) , .D( u0_uk_K_r11_30 ) , .Q( u0_uk_K_r12_30 ) , .QN( u0_uk_n66 ) );
  DFF_X1 u0_uk_K_r12_reg_31 (.CK( clk ) , .D( u0_uk_K_r11_31 ) , .Q( u0_uk_K_r12_31 ) , .QN( u0_uk_n65 ) );
  DFF_X1 u0_uk_K_r12_reg_32 (.CK( clk ) , .D( u0_uk_K_r11_32 ) , .Q( u0_uk_K_r12_32 ) , .QN( u0_uk_n64 ) );
  DFF_X1 u0_uk_K_r12_reg_33 (.CK( clk ) , .D( u0_uk_K_r11_33 ) , .Q( u0_uk_K_r12_33 ) );
  DFF_X1 u0_uk_K_r12_reg_34 (.CK( clk ) , .D( u0_uk_K_r11_34 ) , .Q( u0_uk_K_r12_34 ) , .QN( u0_uk_n62 ) );
  DFF_X1 u0_uk_K_r12_reg_35 (.CK( clk ) , .D( u0_uk_K_r11_35 ) , .Q( u0_uk_K_r12_35 ) , .QN( u0_uk_n61 ) );
  DFF_X1 u0_uk_K_r12_reg_36 (.CK( clk ) , .D( u0_uk_K_r11_36 ) , .Q( u0_uk_K_r12_36 ) );
  DFF_X1 u0_uk_K_r12_reg_37 (.CK( clk ) , .D( u0_uk_K_r11_37 ) , .Q( u0_uk_K_r12_37 ) , .QN( u0_uk_n59 ) );
  DFF_X1 u0_uk_K_r12_reg_38 (.CK( clk ) , .D( u0_uk_K_r11_38 ) , .Q( u0_uk_K_r12_38 ) , .QN( u0_uk_n58 ) );
  DFF_X1 u0_uk_K_r12_reg_39 (.CK( clk ) , .D( u0_uk_K_r11_39 ) , .Q( u0_uk_K_r12_39 ) );
  DFF_X1 u0_uk_K_r12_reg_4 (.CK( clk ) , .D( u0_uk_K_r11_4 ) , .Q( u0_uk_K_r12_4 ) , .QN( u0_uk_n86 ) );
  DFF_X1 u0_uk_K_r12_reg_40 (.CK( clk ) , .D( u0_uk_K_r11_40 ) , .Q( u0_uk_K_r12_40 ) , .QN( u0_uk_n57 ) );
  DFF_X1 u0_uk_K_r12_reg_41 (.CK( clk ) , .D( u0_uk_K_r11_41 ) , .Q( u0_uk_K_r12_41 ) );
  DFF_X1 u0_uk_K_r12_reg_42 (.CK( clk ) , .D( u0_uk_K_r11_42 ) , .Q( u0_uk_K_r12_42 ) );
  DFF_X1 u0_uk_K_r12_reg_43 (.CK( clk ) , .D( u0_uk_K_r11_43 ) , .Q( u0_uk_K_r12_43 ) , .QN( u0_uk_n56 ) );
  DFF_X1 u0_uk_K_r12_reg_44 (.CK( clk ) , .D( u0_uk_K_r11_44 ) , .Q( u0_uk_K_r12_44 ) );
  DFF_X1 u0_uk_K_r12_reg_45 (.CK( clk ) , .D( u0_uk_K_r11_45 ) , .Q( u0_uk_K_r12_45 ) , .QN( u0_uk_n55 ) );
  DFF_X1 u0_uk_K_r12_reg_46 (.CK( clk ) , .D( u0_uk_K_r11_46 ) , .Q( u0_uk_K_r12_46 ) , .QN( u0_uk_n54 ) );
  DFF_X1 u0_uk_K_r12_reg_47 (.CK( clk ) , .D( u0_uk_K_r11_47 ) , .Q( u0_uk_K_r12_47 ) );
  DFF_X1 u0_uk_K_r12_reg_48 (.CK( clk ) , .D( u0_uk_K_r11_48 ) , .Q( u0_uk_K_r12_48 ) , .QN( u0_uk_n53 ) );
  DFF_X1 u0_uk_K_r12_reg_49 (.CK( clk ) , .D( u0_uk_K_r11_49 ) , .Q( u0_uk_K_r12_49 ) , .QN( u0_uk_n52 ) );
  DFF_X1 u0_uk_K_r12_reg_5 (.CK( clk ) , .D( u0_uk_K_r11_5 ) , .Q( u0_uk_K_r12_5 ) , .QN( u0_uk_n85 ) );
  DFF_X1 u0_uk_K_r12_reg_50 (.CK( clk ) , .D( u0_uk_K_r11_50 ) , .Q( u0_uk_K_r12_50 ) , .QN( u0_uk_n51 ) );
  DFF_X1 u0_uk_K_r12_reg_51 (.CK( clk ) , .D( u0_uk_K_r11_51 ) , .Q( u0_uk_K_r12_51 ) , .QN( u0_uk_n50 ) );
  DFF_X1 u0_uk_K_r12_reg_52 (.CK( clk ) , .D( u0_uk_K_r11_52 ) , .Q( u0_uk_K_r12_52 ) , .QN( u0_uk_n49 ) );
  DFF_X1 u0_uk_K_r12_reg_53 (.CK( clk ) , .D( u0_uk_K_r11_53 ) , .Q( u0_uk_K_r12_53 ) , .QN( u0_uk_n48 ) );
  DFF_X1 u0_uk_K_r12_reg_54 (.CK( clk ) , .D( u0_uk_K_r11_54 ) , .Q( u0_uk_K_r12_54 ) , .QN( u0_uk_n47 ) );
  DFF_X1 u0_uk_K_r12_reg_55 (.CK( clk ) , .D( u0_uk_K_r11_55 ) , .Q( u0_uk_K_r12_55 ) , .QN( u0_uk_n46 ) );
  DFF_X1 u0_uk_K_r12_reg_6 (.CK( clk ) , .D( u0_uk_K_r11_6 ) , .Q( u0_uk_K_r12_6 ) , .QN( u0_uk_n84 ) );
  DFF_X1 u0_uk_K_r12_reg_7 (.CK( clk ) , .D( u0_uk_K_r11_7 ) , .Q( u0_uk_K_r12_7 ) );
  DFF_X1 u0_uk_K_r12_reg_8 (.CK( clk ) , .D( u0_uk_K_r11_8 ) , .Q( u0_uk_K_r12_8 ) , .QN( u0_uk_n82 ) );
  DFF_X1 u0_uk_K_r12_reg_9 (.CK( clk ) , .D( u0_uk_K_r11_9 ) , .Q( u0_uk_K_r12_9 ) , .QN( u0_uk_n81 ) );
  DFF_X1 u0_uk_K_r13_reg_0 (.CK( clk ) , .D( u0_uk_K_r12_0 ) , .Q( u0_uk_K_r13_0 ) , .QN( u0_uk_n45 ) );
  DFF_X1 u0_uk_K_r13_reg_1 (.CK( clk ) , .D( u0_uk_K_r12_1 ) , .Q( u0_uk_K_r13_1 ) );
  DFF_X1 u0_uk_K_r13_reg_10 (.CK( clk ) , .D( u0_uk_K_r12_10 ) , .Q( u0_uk_K_r13_10 ) , .QN( u0_uk_n38 ) );
  DFF_X1 u0_uk_K_r13_reg_11 (.CK( clk ) , .D( u0_uk_K_r12_11 ) , .Q( u0_uk_K_r13_11 ) , .QN( u0_uk_n37 ) );
  DFF_X1 u0_uk_K_r13_reg_12 (.CK( clk ) , .D( u0_uk_K_r12_12 ) , .Q( u0_uk_K_r13_12 ) , .QN( u0_uk_n36 ) );
  DFF_X1 u0_uk_K_r13_reg_13 (.CK( clk ) , .D( u0_uk_K_r12_13 ) , .Q( u0_uk_K_r13_13 ) , .QN( u0_uk_n35 ) );
  DFF_X1 u0_uk_K_r13_reg_14 (.CK( clk ) , .D( u0_uk_K_r12_14 ) , .Q( u0_uk_K_r13_14 ) , .QN( u0_uk_n34 ) );
  DFF_X1 u0_uk_K_r13_reg_15 (.CK( clk ) , .D( u0_uk_K_r12_15 ) , .Q( u0_uk_K_r13_15 ) , .QN( u0_uk_n33 ) );
  DFF_X1 u0_uk_K_r13_reg_16 (.CK( clk ) , .D( u0_uk_K_r12_16 ) , .Q( u0_uk_K_r13_16 ) , .QN( u0_uk_n32 ) );
  DFF_X1 u0_uk_K_r13_reg_17 (.CK( clk ) , .D( u0_uk_K_r12_17 ) , .Q( u0_uk_K_r13_17 ) );
  DFF_X1 u0_uk_K_r13_reg_18 (.CK( clk ) , .D( u0_uk_K_r12_18 ) , .Q( u0_uk_K_r13_18 ) , .QN( u0_uk_n30 ) );
  DFF_X1 u0_uk_K_r13_reg_19 (.CK( clk ) , .D( u0_uk_K_r12_19 ) , .Q( u0_uk_K_r13_19 ) );
  DFF_X1 u0_uk_K_r13_reg_2 (.CK( clk ) , .D( u0_uk_K_r12_2 ) , .Q( u0_uk_K_r13_2 ) );
  DFF_X1 u0_uk_K_r13_reg_20 (.CK( clk ) , .D( u0_uk_K_r12_20 ) , .Q( u0_uk_K_r13_20 ) , .QN( u0_uk_n29 ) );
  DFF_X1 u0_uk_K_r13_reg_21 (.CK( clk ) , .D( u0_uk_K_r12_21 ) , .Q( u0_uk_K_r13_21 ) , .QN( u0_uk_n28 ) );
  DFF_X1 u0_uk_K_r13_reg_22 (.CK( clk ) , .D( u0_uk_K_r12_22 ) , .Q( u0_uk_K_r13_22 ) );
  DFF_X1 u0_uk_K_r13_reg_23 (.CK( clk ) , .D( u0_uk_K_r12_23 ) , .Q( u0_uk_K_r13_23 ) );
  DFF_X1 u0_uk_K_r13_reg_24 (.CK( clk ) , .D( u0_uk_K_r12_24 ) , .Q( u0_uk_K_r13_24 ) , .QN( u0_uk_n26 ) );
  DFF_X1 u0_uk_K_r13_reg_25 (.CK( clk ) , .D( u0_uk_K_r12_25 ) , .Q( u0_uk_K_r13_25 ) );
  DFF_X1 u0_uk_K_r13_reg_26 (.CK( clk ) , .D( u0_uk_K_r12_26 ) , .Q( u0_uk_K_r13_26 ) , .QN( u0_uk_n25 ) );
  DFF_X1 u0_uk_K_r13_reg_27 (.CK( clk ) , .D( u0_uk_K_r12_27 ) , .Q( u0_uk_K_r13_27 ) , .QN( u0_uk_n24 ) );
  DFF_X1 u0_uk_K_r13_reg_28 (.CK( clk ) , .D( u0_uk_K_r12_28 ) , .Q( u0_uk_K_r13_28 ) , .QN( u0_uk_n23 ) );
  DFF_X1 u0_uk_K_r13_reg_29 (.CK( clk ) , .D( u0_uk_K_r12_29 ) , .Q( u0_uk_K_r13_29 ) , .QN( u0_uk_n22 ) );
  DFF_X1 u0_uk_K_r13_reg_3 (.CK( clk ) , .D( u0_uk_K_r12_3 ) , .Q( u0_uk_K_r13_3 ) , .QN( u0_uk_n44 ) );
  DFF_X1 u0_uk_K_r13_reg_30 (.CK( clk ) , .D( u0_uk_K_r12_30 ) , .Q( u0_uk_K_r13_30 ) , .QN( u0_uk_n21 ) );
  DFF_X1 u0_uk_K_r13_reg_31 (.CK( clk ) , .D( u0_uk_K_r12_31 ) , .Q( u0_uk_K_r13_31 ) );
  DFF_X1 u0_uk_K_r13_reg_32 (.CK( clk ) , .D( u0_uk_K_r12_32 ) , .Q( u0_uk_K_r13_32 ) );
  DFF_X1 u0_uk_K_r13_reg_33 (.CK( clk ) , .D( u0_uk_K_r12_33 ) , .Q( u0_uk_K_r13_33 ) , .QN( u0_uk_n20 ) );
  DFF_X1 u0_uk_K_r13_reg_34 (.CK( clk ) , .D( u0_uk_K_r12_34 ) , .Q( u0_uk_K_r13_34 ) , .QN( u0_uk_n19 ) );
  DFF_X1 u0_uk_K_r13_reg_35 (.CK( clk ) , .D( u0_uk_K_r12_35 ) , .Q( u0_uk_K_r13_35 ) );
  DFF_X1 u0_uk_K_r13_reg_36 (.CK( clk ) , .D( u0_uk_K_r12_36 ) , .Q( u0_uk_K_r13_36 ) );
  DFF_X1 u0_uk_K_r13_reg_37 (.CK( clk ) , .D( u0_uk_K_r12_37 ) , .Q( u0_uk_K_r13_37 ) , .QN( u0_uk_n18 ) );
  DFF_X1 u0_uk_K_r13_reg_38 (.CK( clk ) , .D( u0_uk_K_r12_38 ) , .Q( u0_uk_K_r13_38 ) );
  DFF_X1 u0_uk_K_r13_reg_39 (.CK( clk ) , .D( u0_uk_K_r12_39 ) , .Q( u0_uk_K_r13_39 ) , .QN( u0_uk_n16 ) );
  DFF_X1 u0_uk_K_r13_reg_4 (.CK( clk ) , .D( u0_uk_K_r12_4 ) , .Q( u0_uk_K_r13_4 ) );
  DFF_X1 u0_uk_K_r13_reg_40 (.CK( clk ) , .D( u0_uk_K_r12_40 ) , .Q( u0_uk_K_r13_40 ) , .QN( u0_uk_n15 ) );
  DFF_X1 u0_uk_K_r13_reg_41 (.CK( clk ) , .D( u0_uk_K_r12_41 ) , .Q( u0_uk_K_r13_41 ) , .QN( u0_uk_n14 ) );
  DFF_X1 u0_uk_K_r13_reg_42 (.CK( clk ) , .D( u0_uk_K_r12_42 ) , .Q( u0_uk_K_r13_42 ) , .QN( u0_uk_n13 ) );
  DFF_X1 u0_uk_K_r13_reg_43 (.CK( clk ) , .D( u0_uk_K_r12_43 ) , .Q( u0_uk_K_r13_43 ) , .QN( u0_uk_n12 ) );
  DFF_X1 u0_uk_K_r13_reg_44 (.CK( clk ) , .D( u0_uk_K_r12_44 ) , .Q( u0_uk_K_r13_44 ) );
  DFF_X1 u0_uk_K_r13_reg_45 (.CK( clk ) , .D( u0_uk_K_r12_45 ) , .Q( u0_uk_K_r13_45 ) , .QN( u0_uk_n9 ) );
  DFF_X1 u0_uk_K_r13_reg_46 (.CK( clk ) , .D( u0_uk_K_r12_46 ) , .Q( u0_uk_K_r13_46 ) , .QN( u0_uk_n8 ) );
  DFF_X1 u0_uk_K_r13_reg_47 (.CK( clk ) , .D( u0_uk_K_r12_47 ) , .Q( u0_uk_K_r13_47 ) , .QN( u0_uk_n7 ) );
  DFF_X1 u0_uk_K_r13_reg_48 (.CK( clk ) , .D( u0_uk_K_r12_48 ) , .Q( u0_uk_K_r13_48 ) , .QN( u0_uk_n6 ) );
  DFF_X1 u0_uk_K_r13_reg_49 (.CK( clk ) , .D( u0_uk_K_r12_49 ) , .Q( u0_uk_K_r13_49 ) , .QN( u0_uk_n5 ) );
  DFF_X1 u0_uk_K_r13_reg_5 (.CK( clk ) , .D( u0_uk_K_r12_5 ) , .Q( u0_uk_K_r13_5 ) , .QN( u0_uk_n43 ) );
  DFF_X1 u0_uk_K_r13_reg_50 (.CK( clk ) , .D( u0_uk_K_r12_50 ) , .Q( u0_uk_K_r13_50 ) , .QN( u0_uk_n4 ) );
  DFF_X1 u0_uk_K_r13_reg_51 (.CK( clk ) , .D( u0_uk_K_r12_51 ) , .Q( u0_uk_K_r13_51 ) , .QN( u0_uk_n3 ) );
  DFF_X1 u0_uk_K_r13_reg_52 (.CK( clk ) , .D( u0_uk_K_r12_52 ) , .Q( u0_uk_K_r13_52 ) , .QN( u0_uk_n2 ) );
  DFF_X1 u0_uk_K_r13_reg_53 (.CK( clk ) , .D( u0_uk_K_r12_53 ) , .Q( u0_uk_K_r13_53 ) );
  DFF_X1 u0_uk_K_r13_reg_54 (.CK( clk ) , .D( u0_uk_K_r12_54 ) , .Q( u0_uk_K_r13_54 ) , .QN( u0_uk_n1 ) );
  DFF_X1 u0_uk_K_r13_reg_55 (.CK( clk ) , .D( u0_uk_K_r12_55 ) , .Q( u0_uk_K_r13_55 ) );
  DFF_X1 u0_uk_K_r13_reg_6 (.CK( clk ) , .D( u0_uk_K_r12_6 ) , .Q( u0_uk_K_r13_6 ) , .QN( u0_uk_n42 ) );
  DFF_X1 u0_uk_K_r13_reg_7 (.CK( clk ) , .D( u0_uk_K_r12_7 ) , .Q( u0_uk_K_r13_7 ) , .QN( u0_uk_n41 ) );
  DFF_X1 u0_uk_K_r13_reg_8 (.CK( clk ) , .D( u0_uk_K_r12_8 ) , .Q( u0_uk_K_r13_8 ) , .QN( u0_uk_n40 ) );
  DFF_X1 u0_uk_K_r13_reg_9 (.CK( clk ) , .D( u0_uk_K_r12_9 ) , .Q( u0_uk_K_r13_9 ) , .QN( u0_uk_n39 ) );
  DFF_X1 u0_uk_K_r14_reg_0 (.CK( clk ) , .D( u0_uk_K_r13_0 ) , .QN( u0_uk_n670 ) );
  DFF_X1 u0_uk_K_r14_reg_1 (.CK( clk ) , .D( u0_uk_K_r13_1 ) , .QN( u0_uk_n669 ) );
  DFF_X1 u0_uk_K_r14_reg_10 (.CK( clk ) , .D( u0_uk_K_r13_10 ) , .Q( u0_uk_K_r14_10 ) );
  DFF_X1 u0_uk_K_r14_reg_11 (.CK( clk ) , .D( u0_uk_K_r13_11 ) , .Q( u0_uk_K_r14_11 ) );
  DFF_X1 u0_uk_K_r14_reg_12 (.CK( clk ) , .D( u0_uk_K_r13_12 ) , .Q( u0_uk_K_r14_12 ) );
  DFF_X1 u0_uk_K_r14_reg_13 (.CK( clk ) , .D( u0_uk_K_r13_13 ) , .QN( u0_uk_n664 ) );
  DFF_X1 u0_uk_K_r14_reg_14 (.CK( clk ) , .D( u0_uk_K_r13_14 ) , .QN( u0_uk_n663 ) );
  DFF_X1 u0_uk_K_r14_reg_15 (.CK( clk ) , .D( u0_uk_K_r13_15 ) , .Q( u0_uk_K_r14_15 ) );
  DFF_X1 u0_uk_K_r14_reg_16 (.CK( clk ) , .D( u0_uk_K_r13_16 ) , .Q( u0_uk_K_r14_16 ) );
  DFF_X1 u0_uk_K_r14_reg_17 (.CK( clk ) , .D( u0_uk_K_r13_17 ) , .QN( u0_uk_n661 ) );
  DFF_X1 u0_uk_K_r14_reg_18 (.CK( clk ) , .D( u0_uk_K_r13_18 ) , .Q( u0_uk_K_r14_18 ) );
  DFF_X1 u0_uk_K_r14_reg_19 (.CK( clk ) , .D( u0_uk_K_r13_19 ) , .QN( u0_uk_n660 ) );
  DFF_X1 u0_uk_K_r14_reg_2 (.CK( clk ) , .D( u0_uk_K_r13_2 ) , .Q( u0_uk_K_r14_2 ) );
  DFF_X1 u0_uk_K_r14_reg_20 (.CK( clk ) , .D( u0_uk_K_r13_20 ) , .QN( u0_uk_n659 ) );
  DFF_X1 u0_uk_K_r14_reg_21 (.CK( clk ) , .D( u0_uk_K_r13_21 ) , .QN( u0_uk_n658 ) );
  DFF_X1 u0_uk_K_r14_reg_22 (.CK( clk ) , .D( u0_uk_K_r13_22 ) , .QN( u0_uk_n657 ) );
  DFF_X1 u0_uk_K_r14_reg_23 (.CK( clk ) , .D( u0_uk_K_r13_23 ) , .Q( u0_uk_K_r14_23 ) , .QN( u0_uk_n655 ) );
  DFF_X1 u0_uk_K_r14_reg_24 (.CK( clk ) , .D( u0_uk_K_r13_24 ) , .QN( u0_uk_n654 ) );
  DFF_X1 u0_uk_K_r14_reg_25 (.CK( clk ) , .D( u0_uk_K_r13_25 ) , .QN( u0_uk_n653 ) );
  DFF_X1 u0_uk_K_r14_reg_26 (.CK( clk ) , .D( u0_uk_K_r13_26 ) , .QN( u0_uk_n652 ) );
  DFF_X1 u0_uk_K_r14_reg_27 (.CK( clk ) , .D( u0_uk_K_r13_27 ) , .QN( u0_uk_n651 ) );
  DFF_X1 u0_uk_K_r14_reg_28 (.CK( clk ) , .D( u0_uk_K_r13_28 ) , .QN( u0_uk_n650 ) );
  DFF_X1 u0_uk_K_r14_reg_29 (.CK( clk ) , .D( u0_uk_K_r13_29 ) , .QN( u0_uk_n649 ) );
  DFF_X1 u0_uk_K_r14_reg_3 (.CK( clk ) , .D( u0_uk_K_r13_3 ) , .Q( u0_uk_K_r14_3 ) );
  DFF_X1 u0_uk_K_r14_reg_30 (.CK( clk ) , .D( u0_uk_K_r13_30 ) , .QN( u0_uk_n648 ) );
  DFF_X1 u0_uk_K_r14_reg_31 (.CK( clk ) , .D( u0_uk_K_r13_31 ) , .QN( u0_uk_n647 ) );
  DFF_X1 u0_uk_K_r14_reg_32 (.CK( clk ) , .D( u0_uk_K_r13_32 ) , .QN( u0_uk_n646 ) );
  DFF_X1 u0_uk_K_r14_reg_33 (.CK( clk ) , .D( u0_uk_K_r13_33 ) , .QN( u0_uk_n645 ) );
  DFF_X1 u0_uk_K_r14_reg_34 (.CK( clk ) , .D( u0_uk_K_r13_34 ) , .QN( u0_uk_n644 ) );
  DFF_X1 u0_uk_K_r14_reg_35 (.CK( clk ) , .D( u0_uk_K_r13_35 ) , .QN( u0_uk_n643 ) );
  DFF_X1 u0_uk_K_r14_reg_36 (.CK( clk ) , .D( u0_uk_K_r13_36 ) , .QN( u0_uk_n642 ) );
  DFF_X1 u0_uk_K_r14_reg_37 (.CK( clk ) , .D( u0_uk_K_r13_37 ) , .QN( u0_uk_n641 ) );
  DFF_X1 u0_uk_K_r14_reg_38 (.CK( clk ) , .D( u0_uk_K_r13_38 ) , .Q( u0_uk_K_r14_38 ) );
  DFF_X1 u0_uk_K_r14_reg_39 (.CK( clk ) , .D( u0_uk_K_r13_39 ) , .Q( u0_uk_K_r14_39 ) );
  DFF_X1 u0_uk_K_r14_reg_4 (.CK( clk ) , .D( u0_uk_K_r13_4 ) , .QN( u0_uk_n668 ) );
  DFF_X1 u0_uk_K_r14_reg_40 (.CK( clk ) , .D( u0_uk_K_r13_40 ) , .QN( u0_uk_n640 ) );
  DFF_X1 u0_uk_K_r14_reg_41 (.CK( clk ) , .D( u0_uk_K_r13_41 ) , .QN( u0_uk_n639 ) );
  DFF_X1 u0_uk_K_r14_reg_42 (.CK( clk ) , .D( u0_uk_K_r13_42 ) , .Q( u0_uk_K_r14_42 ) );
  DFF_X1 u0_uk_K_r14_reg_43 (.CK( clk ) , .D( u0_uk_K_r13_43 ) , .Q( u0_uk_K_r14_43 ) );
  DFF_X1 u0_uk_K_r14_reg_44 (.CK( clk ) , .D( u0_uk_K_r13_44 ) , .QN( u0_uk_n638 ) );
  DFF_X1 u0_uk_K_r14_reg_45 (.CK( clk ) , .D( u0_uk_K_r13_45 ) , .Q( u0_uk_K_r14_45 ) );
  DFF_X1 u0_uk_K_r14_reg_46 (.CK( clk ) , .D( u0_uk_K_r13_46 ) , .Q( u0_uk_K_r14_46 ) );
  DFF_X1 u0_uk_K_r14_reg_47 (.CK( clk ) , .D( u0_uk_K_r13_47 ) , .QN( u0_uk_n637 ) );
  DFF_X1 u0_uk_K_r14_reg_48 (.CK( clk ) , .D( u0_uk_K_r13_48 ) , .QN( u0_uk_n636 ) );
  DFF_X1 u0_uk_K_r14_reg_49 (.CK( clk ) , .D( u0_uk_K_r13_49 ) , .QN( u0_uk_n635 ) );
  DFF_X1 u0_uk_K_r14_reg_5 (.CK( clk ) , .D( u0_uk_K_r13_5 ) , .Q( u0_uk_K_r14_5 ) );
  DFF_X1 u0_uk_K_r14_reg_50 (.CK( clk ) , .D( u0_uk_K_r13_50 ) , .Q( u0_uk_K_r14_50 ) );
  DFF_X1 u0_uk_K_r14_reg_51 (.CK( clk ) , .D( u0_uk_K_r13_51 ) , .QN( u0_uk_n633 ) );
  DFF_X1 u0_uk_K_r14_reg_52 (.CK( clk ) , .D( u0_uk_K_r13_52 ) , .QN( u0_uk_n632 ) );
  DFF_X1 u0_uk_K_r14_reg_53 (.CK( clk ) , .D( u0_uk_K_r13_53 ) , .QN( u0_uk_n631 ) );
  DFF_X1 u0_uk_K_r14_reg_54 (.CK( clk ) , .D( u0_uk_K_r13_54 ) , .QN( u0_uk_n630 ) );
  DFF_X1 u0_uk_K_r14_reg_55 (.CK( clk ) , .D( u0_uk_K_r13_55 ) , .QN( u0_uk_n629 ) );
  DFF_X1 u0_uk_K_r14_reg_6 (.CK( clk ) , .D( u0_uk_K_r13_6 ) , .QN( u0_uk_n667 ) );
  DFF_X1 u0_uk_K_r14_reg_7 (.CK( clk ) , .D( u0_uk_K_r13_7 ) , .QN( u0_uk_n666 ) );
  DFF_X1 u0_uk_K_r14_reg_8 (.CK( clk ) , .D( u0_uk_K_r13_8 ) , .Q( u0_uk_K_r14_8 ) );
  DFF_X1 u0_uk_K_r14_reg_9 (.CK( clk ) , .D( u0_uk_K_r13_9 ) , .Q( u0_uk_K_r14_9 ) );
  DFF_X1 u0_uk_K_r1_reg_0 (.CK( clk ) , .D( u0_uk_K_r0_0 ) , .Q( u0_uk_K_r1_0 ) , .QN( u0_uk_n581 ) );
  DFF_X1 u0_uk_K_r1_reg_1 (.CK( clk ) , .D( u0_uk_K_r0_1 ) , .Q( u0_uk_K_r1_1 ) , .QN( u0_uk_n580 ) );
  DFF_X1 u0_uk_K_r1_reg_10 (.CK( clk ) , .D( u0_uk_K_r0_10 ) , .Q( u0_uk_K_r1_10 ) );
  DFF_X1 u0_uk_K_r1_reg_11 (.CK( clk ) , .D( u0_uk_K_r0_11 ) , .Q( u0_uk_K_r1_11 ) , .QN( u0_uk_n573 ) );
  DFF_X1 u0_uk_K_r1_reg_12 (.CK( clk ) , .D( u0_uk_K_r0_12 ) , .Q( u0_uk_K_r1_12 ) , .QN( u0_uk_n572 ) );
  DFF_X1 u0_uk_K_r1_reg_13 (.CK( clk ) , .D( u0_uk_K_r0_13 ) , .Q( u0_uk_K_r1_13 ) , .QN( u0_uk_n571 ) );
  DFF_X1 u0_uk_K_r1_reg_14 (.CK( clk ) , .D( u0_uk_K_r0_14 ) , .Q( u0_uk_K_r1_14 ) , .QN( u0_uk_n570 ) );
  DFF_X1 u0_uk_K_r1_reg_15 (.CK( clk ) , .D( u0_uk_K_r0_15 ) , .Q( u0_uk_K_r1_15 ) );
  DFF_X1 u0_uk_K_r1_reg_16 (.CK( clk ) , .D( u0_uk_K_r0_16 ) , .Q( u0_uk_K_r1_16 ) );
  DFF_X1 u0_uk_K_r1_reg_17 (.CK( clk ) , .D( u0_uk_K_r0_17 ) , .Q( u0_uk_K_r1_17 ) , .QN( u0_uk_n569 ) );
  DFF_X1 u0_uk_K_r1_reg_18 (.CK( clk ) , .D( u0_uk_K_r0_18 ) , .Q( u0_uk_K_r1_18 ) );
  DFF_X1 u0_uk_K_r1_reg_19 (.CK( clk ) , .D( u0_uk_K_r0_19 ) , .Q( u0_uk_K_r1_19 ) , .QN( u0_uk_n568 ) );
  DFF_X1 u0_uk_K_r1_reg_2 (.CK( clk ) , .D( u0_uk_K_r0_2 ) , .Q( u0_uk_K_r1_2 ) , .QN( u0_uk_n579 ) );
  DFF_X1 u0_uk_K_r1_reg_20 (.CK( clk ) , .D( u0_uk_K_r0_20 ) , .Q( u0_uk_K_r1_20 ) , .QN( u0_uk_n567 ) );
  DFF_X1 u0_uk_K_r1_reg_21 (.CK( clk ) , .D( u0_uk_K_r0_21 ) , .Q( u0_uk_K_r1_21 ) );
  DFF_X1 u0_uk_K_r1_reg_22 (.CK( clk ) , .D( u0_uk_K_r0_22 ) , .Q( u0_uk_K_r1_22 ) );
  DFF_X1 u0_uk_K_r1_reg_23 (.CK( clk ) , .D( u0_uk_K_r0_23 ) , .Q( u0_uk_K_r1_23 ) , .QN( u0_uk_n566 ) );
  DFF_X1 u0_uk_K_r1_reg_24 (.CK( clk ) , .D( u0_uk_K_r0_24 ) , .Q( u0_uk_K_r1_24 ) , .QN( u0_uk_n565 ) );
  DFF_X1 u0_uk_K_r1_reg_25 (.CK( clk ) , .D( u0_uk_K_r0_25 ) , .Q( u0_uk_K_r1_25 ) , .QN( u0_uk_n564 ) );
  DFF_X1 u0_uk_K_r1_reg_26 (.CK( clk ) , .D( u0_uk_K_r0_26 ) , .Q( u0_uk_K_r1_26 ) , .QN( u0_uk_n563 ) );
  DFF_X1 u0_uk_K_r1_reg_27 (.CK( clk ) , .D( u0_uk_K_r0_27 ) , .Q( u0_uk_K_r1_27 ) , .QN( u0_uk_n562 ) );
  DFF_X1 u0_uk_K_r1_reg_28 (.CK( clk ) , .D( u0_uk_K_r0_28 ) , .Q( u0_uk_K_r1_28 ) , .QN( u0_uk_n561 ) );
  DFF_X1 u0_uk_K_r1_reg_29 (.CK( clk ) , .D( u0_uk_K_r0_29 ) , .Q( u0_uk_K_r1_29 ) , .QN( u0_uk_n560 ) );
  DFF_X1 u0_uk_K_r1_reg_3 (.CK( clk ) , .D( u0_uk_K_r0_3 ) , .Q( u0_uk_K_r1_3 ) , .QN( u0_uk_n578 ) );
  DFF_X1 u0_uk_K_r1_reg_30 (.CK( clk ) , .D( u0_uk_K_r0_30 ) , .Q( u0_uk_K_r1_30 ) , .QN( u0_uk_n559 ) );
  DFF_X1 u0_uk_K_r1_reg_31 (.CK( clk ) , .D( u0_uk_K_r0_31 ) , .Q( u0_uk_K_r1_31 ) , .QN( u0_uk_n558 ) );
  DFF_X1 u0_uk_K_r1_reg_32 (.CK( clk ) , .D( u0_uk_K_r0_32 ) , .Q( u0_uk_K_r1_32 ) , .QN( u0_uk_n557 ) );
  DFF_X1 u0_uk_K_r1_reg_33 (.CK( clk ) , .D( u0_uk_K_r0_33 ) , .Q( u0_uk_K_r1_33 ) );
  DFF_X1 u0_uk_K_r1_reg_34 (.CK( clk ) , .D( u0_uk_K_r0_34 ) , .Q( u0_uk_K_r1_34 ) , .QN( u0_uk_n556 ) );
  DFF_X1 u0_uk_K_r1_reg_35 (.CK( clk ) , .D( u0_uk_K_r0_35 ) , .Q( u0_uk_K_r1_35 ) , .QN( u0_uk_n555 ) );
  DFF_X1 u0_uk_K_r1_reg_36 (.CK( clk ) , .D( u0_uk_K_r0_36 ) , .Q( u0_uk_K_r1_36 ) );
  DFF_X1 u0_uk_K_r1_reg_37 (.CK( clk ) , .D( u0_uk_K_r0_37 ) , .Q( u0_uk_K_r1_37 ) , .QN( u0_uk_n554 ) );
  DFF_X1 u0_uk_K_r1_reg_38 (.CK( clk ) , .D( u0_uk_K_r0_38 ) , .Q( u0_uk_K_r1_38 ) , .QN( u0_uk_n553 ) );
  DFF_X1 u0_uk_K_r1_reg_39 (.CK( clk ) , .D( u0_uk_K_r0_39 ) , .Q( u0_uk_K_r1_39 ) );
  DFF_X1 u0_uk_K_r1_reg_4 (.CK( clk ) , .D( u0_uk_K_r0_4 ) , .Q( u0_uk_K_r1_4 ) , .QN( u0_uk_n577 ) );
  DFF_X1 u0_uk_K_r1_reg_40 (.CK( clk ) , .D( u0_uk_K_r0_40 ) , .Q( u0_uk_K_r1_40 ) , .QN( u0_uk_n552 ) );
  DFF_X1 u0_uk_K_r1_reg_41 (.CK( clk ) , .D( u0_uk_K_r0_41 ) , .Q( u0_uk_K_r1_41 ) );
  DFF_X1 u0_uk_K_r1_reg_42 (.CK( clk ) , .D( u0_uk_K_r0_42 ) , .Q( u0_uk_K_r1_42 ) );
  DFF_X1 u0_uk_K_r1_reg_43 (.CK( clk ) , .D( u0_uk_K_r0_43 ) , .Q( u0_uk_K_r1_43 ) , .QN( u0_uk_n550 ) );
  DFF_X1 u0_uk_K_r1_reg_44 (.CK( clk ) , .D( u0_uk_K_r0_44 ) , .Q( u0_uk_K_r1_44 ) );
  DFF_X1 u0_uk_K_r1_reg_45 (.CK( clk ) , .D( u0_uk_K_r0_45 ) , .Q( u0_uk_K_r1_45 ) , .QN( u0_uk_n549 ) );
  DFF_X1 u0_uk_K_r1_reg_46 (.CK( clk ) , .D( u0_uk_K_r0_46 ) , .Q( u0_uk_K_r1_46 ) , .QN( u0_uk_n548 ) );
  DFF_X1 u0_uk_K_r1_reg_47 (.CK( clk ) , .D( u0_uk_K_r0_47 ) , .Q( u0_uk_K_r1_47 ) );
  DFF_X1 u0_uk_K_r1_reg_48 (.CK( clk ) , .D( u0_uk_K_r0_48 ) , .Q( u0_uk_K_r1_48 ) , .QN( u0_uk_n547 ) );
  DFF_X1 u0_uk_K_r1_reg_49 (.CK( clk ) , .D( u0_uk_K_r0_49 ) , .Q( u0_uk_K_r1_49 ) , .QN( u0_uk_n546 ) );
  DFF_X1 u0_uk_K_r1_reg_5 (.CK( clk ) , .D( u0_uk_K_r0_5 ) , .Q( u0_uk_K_r1_5 ) , .QN( u0_uk_n576 ) );
  DFF_X1 u0_uk_K_r1_reg_50 (.CK( clk ) , .D( u0_uk_K_r0_50 ) , .Q( u0_uk_K_r1_50 ) , .QN( u0_uk_n545 ) );
  DFF_X1 u0_uk_K_r1_reg_51 (.CK( clk ) , .D( u0_uk_K_r0_51 ) , .Q( u0_uk_K_r1_51 ) , .QN( u0_uk_n544 ) );
  DFF_X1 u0_uk_K_r1_reg_52 (.CK( clk ) , .D( u0_uk_K_r0_52 ) , .Q( u0_uk_K_r1_52 ) , .QN( u0_uk_n543 ) );
  DFF_X1 u0_uk_K_r1_reg_53 (.CK( clk ) , .D( u0_uk_K_r0_53 ) , .Q( u0_uk_K_r1_53 ) , .QN( u0_uk_n542 ) );
  DFF_X1 u0_uk_K_r1_reg_54 (.CK( clk ) , .D( u0_uk_K_r0_54 ) , .Q( u0_uk_K_r1_54 ) , .QN( u0_uk_n541 ) );
  DFF_X1 u0_uk_K_r1_reg_55 (.CK( clk ) , .D( u0_uk_K_r0_55 ) , .Q( u0_uk_K_r1_55 ) , .QN( u0_uk_n540 ) );
  DFF_X1 u0_uk_K_r1_reg_6 (.CK( clk ) , .D( u0_uk_K_r0_6 ) , .Q( u0_uk_K_r1_6 ) );
  DFF_X1 u0_uk_K_r1_reg_7 (.CK( clk ) , .D( u0_uk_K_r0_7 ) , .Q( u0_uk_K_r1_7 ) );
  DFF_X1 u0_uk_K_r1_reg_8 (.CK( clk ) , .D( u0_uk_K_r0_8 ) , .Q( u0_uk_K_r1_8 ) , .QN( u0_uk_n575 ) );
  DFF_X1 u0_uk_K_r1_reg_9 (.CK( clk ) , .D( u0_uk_K_r0_9 ) , .Q( u0_uk_K_r1_9 ) , .QN( u0_uk_n574 ) );
  DFF_X1 u0_uk_K_r2_reg_0 (.CK( clk ) , .D( u0_uk_K_r1_0 ) , .Q( u0_uk_K_r2_0 ) , .QN( u0_uk_n539 ) );
  DFF_X1 u0_uk_K_r2_reg_1 (.CK( clk ) , .D( u0_uk_K_r1_1 ) , .Q( u0_uk_K_r2_1 ) , .QN( u0_uk_n538 ) );
  DFF_X1 u0_uk_K_r2_reg_10 (.CK( clk ) , .D( u0_uk_K_r1_10 ) , .Q( u0_uk_K_r2_10 ) , .QN( u0_uk_n531 ) );
  DFF_X1 u0_uk_K_r2_reg_11 (.CK( clk ) , .D( u0_uk_K_r1_11 ) , .Q( u0_uk_K_r2_11 ) , .QN( u0_uk_n530 ) );
  DFF_X1 u0_uk_K_r2_reg_12 (.CK( clk ) , .D( u0_uk_K_r1_12 ) , .Q( u0_uk_K_r2_12 ) , .QN( u0_uk_n529 ) );
  DFF_X1 u0_uk_K_r2_reg_13 (.CK( clk ) , .D( u0_uk_K_r1_13 ) , .Q( u0_uk_K_r2_13 ) );
  DFF_X1 u0_uk_K_r2_reg_14 (.CK( clk ) , .D( u0_uk_K_r1_14 ) , .Q( u0_uk_K_r2_14 ) , .QN( u0_uk_n528 ) );
  DFF_X1 u0_uk_K_r2_reg_15 (.CK( clk ) , .D( u0_uk_K_r1_15 ) , .Q( u0_uk_K_r2_15 ) , .QN( u0_uk_n527 ) );
  DFF_X1 u0_uk_K_r2_reg_16 (.CK( clk ) , .D( u0_uk_K_r1_16 ) , .Q( u0_uk_K_r2_16 ) );
  DFF_X1 u0_uk_K_r2_reg_17 (.CK( clk ) , .D( u0_uk_K_r1_17 ) , .Q( u0_uk_K_r2_17 ) , .QN( u0_uk_n525 ) );
  DFF_X1 u0_uk_K_r2_reg_18 (.CK( clk ) , .D( u0_uk_K_r1_18 ) , .Q( u0_uk_K_r2_18 ) );
  DFF_X1 u0_uk_K_r2_reg_19 (.CK( clk ) , .D( u0_uk_K_r1_19 ) , .Q( u0_uk_K_r2_19 ) , .QN( u0_uk_n523 ) );
  DFF_X1 u0_uk_K_r2_reg_2 (.CK( clk ) , .D( u0_uk_K_r1_2 ) , .Q( u0_uk_K_r2_2 ) , .QN( u0_uk_n537 ) );
  DFF_X1 u0_uk_K_r2_reg_20 (.CK( clk ) , .D( u0_uk_K_r1_20 ) , .Q( u0_uk_K_r2_20 ) );
  DFF_X1 u0_uk_K_r2_reg_21 (.CK( clk ) , .D( u0_uk_K_r1_21 ) , .Q( u0_uk_K_r2_21 ) );
  DFF_X1 u0_uk_K_r2_reg_22 (.CK( clk ) , .D( u0_uk_K_r1_22 ) , .Q( u0_uk_K_r2_22 ) , .QN( u0_uk_n522 ) );
  DFF_X1 u0_uk_K_r2_reg_23 (.CK( clk ) , .D( u0_uk_K_r1_23 ) , .Q( u0_uk_K_r2_23 ) , .QN( u0_uk_n521 ) );
  DFF_X1 u0_uk_K_r2_reg_24 (.CK( clk ) , .D( u0_uk_K_r1_24 ) , .Q( u0_uk_K_r2_24 ) );
  DFF_X1 u0_uk_K_r2_reg_25 (.CK( clk ) , .D( u0_uk_K_r1_25 ) , .Q( u0_uk_K_r2_25 ) );
  DFF_X1 u0_uk_K_r2_reg_26 (.CK( clk ) , .D( u0_uk_K_r1_26 ) , .Q( u0_uk_K_r2_26 ) );
  DFF_X1 u0_uk_K_r2_reg_27 (.CK( clk ) , .D( u0_uk_K_r1_27 ) , .Q( u0_uk_K_r2_27 ) );
  DFF_X1 u0_uk_K_r2_reg_28 (.CK( clk ) , .D( u0_uk_K_r1_28 ) , .Q( u0_uk_K_r2_28 ) );
  DFF_X1 u0_uk_K_r2_reg_29 (.CK( clk ) , .D( u0_uk_K_r1_29 ) , .Q( u0_uk_K_r2_29 ) );
  DFF_X1 u0_uk_K_r2_reg_3 (.CK( clk ) , .D( u0_uk_K_r1_3 ) , .Q( u0_uk_K_r2_3 ) , .QN( u0_uk_n536 ) );
  DFF_X1 u0_uk_K_r2_reg_30 (.CK( clk ) , .D( u0_uk_K_r1_30 ) , .Q( u0_uk_K_r2_30 ) );
  DFF_X1 u0_uk_K_r2_reg_31 (.CK( clk ) , .D( u0_uk_K_r1_31 ) , .Q( u0_uk_K_r2_31 ) );
  DFF_X1 u0_uk_K_r2_reg_32 (.CK( clk ) , .D( u0_uk_K_r1_32 ) , .Q( u0_uk_K_r2_32 ) , .QN( u0_uk_n519 ) );
  DFF_X1 u0_uk_K_r2_reg_33 (.CK( clk ) , .D( u0_uk_K_r1_33 ) , .Q( u0_uk_K_r2_33 ) );
  DFF_X1 u0_uk_K_r2_reg_34 (.CK( clk ) , .D( u0_uk_K_r1_34 ) , .Q( u0_uk_K_r2_34 ) , .QN( u0_uk_n517 ) );
  DFF_X1 u0_uk_K_r2_reg_35 (.CK( clk ) , .D( u0_uk_K_r1_35 ) , .Q( u0_uk_K_r2_35 ) , .QN( u0_uk_n516 ) );
  DFF_X1 u0_uk_K_r2_reg_36 (.CK( clk ) , .D( u0_uk_K_r1_36 ) , .Q( u0_uk_K_r2_36 ) , .QN( u0_uk_n514 ) );
  DFF_X1 u0_uk_K_r2_reg_37 (.CK( clk ) , .D( u0_uk_K_r1_37 ) , .Q( u0_uk_K_r2_37 ) , .QN( u0_uk_n513 ) );
  DFF_X1 u0_uk_K_r2_reg_38 (.CK( clk ) , .D( u0_uk_K_r1_38 ) , .Q( u0_uk_K_r2_38 ) , .QN( u0_uk_n512 ) );
  DFF_X1 u0_uk_K_r2_reg_39 (.CK( clk ) , .D( u0_uk_K_r1_39 ) , .Q( u0_uk_K_r2_39 ) , .QN( u0_uk_n511 ) );
  DFF_X1 u0_uk_K_r2_reg_4 (.CK( clk ) , .D( u0_uk_K_r1_4 ) , .Q( u0_uk_K_r2_4 ) );
  DFF_X1 u0_uk_K_r2_reg_40 (.CK( clk ) , .D( u0_uk_K_r1_40 ) , .Q( u0_uk_K_r2_40 ) , .QN( u0_uk_n510 ) );
  DFF_X1 u0_uk_K_r2_reg_41 (.CK( clk ) , .D( u0_uk_K_r1_41 ) , .Q( u0_uk_K_r2_41 ) );
  DFF_X1 u0_uk_K_r2_reg_42 (.CK( clk ) , .D( u0_uk_K_r1_42 ) , .Q( u0_uk_K_r2_42 ) , .QN( u0_uk_n508 ) );
  DFF_X1 u0_uk_K_r2_reg_43 (.CK( clk ) , .D( u0_uk_K_r1_43 ) , .Q( u0_uk_K_r2_43 ) , .QN( u0_uk_n507 ) );
  DFF_X1 u0_uk_K_r2_reg_44 (.CK( clk ) , .D( u0_uk_K_r1_44 ) , .Q( u0_uk_K_r2_44 ) , .QN( u0_uk_n506 ) );
  DFF_X1 u0_uk_K_r2_reg_45 (.CK( clk ) , .D( u0_uk_K_r1_45 ) , .Q( u0_uk_K_r2_45 ) , .QN( u0_uk_n505 ) );
  DFF_X1 u0_uk_K_r2_reg_46 (.CK( clk ) , .D( u0_uk_K_r1_46 ) , .Q( u0_uk_K_r2_46 ) );
  DFF_X1 u0_uk_K_r2_reg_47 (.CK( clk ) , .D( u0_uk_K_r1_47 ) , .Q( u0_uk_K_r2_47 ) );
  DFF_X1 u0_uk_K_r2_reg_48 (.CK( clk ) , .D( u0_uk_K_r1_48 ) , .Q( u0_uk_K_r2_48 ) , .QN( u0_uk_n502 ) );
  DFF_X1 u0_uk_K_r2_reg_49 (.CK( clk ) , .D( u0_uk_K_r1_49 ) , .Q( u0_uk_K_r2_49 ) );
  DFF_X1 u0_uk_K_r2_reg_5 (.CK( clk ) , .D( u0_uk_K_r1_5 ) , .Q( u0_uk_K_r2_5 ) , .QN( u0_uk_n535 ) );
  DFF_X1 u0_uk_K_r2_reg_50 (.CK( clk ) , .D( u0_uk_K_r1_50 ) , .Q( u0_uk_K_r2_50 ) );
  DFF_X1 u0_uk_K_r2_reg_51 (.CK( clk ) , .D( u0_uk_K_r1_51 ) , .Q( u0_uk_K_r2_51 ) , .QN( u0_uk_n499 ) );
  DFF_X1 u0_uk_K_r2_reg_52 (.CK( clk ) , .D( u0_uk_K_r1_52 ) , .Q( u0_uk_K_r2_52 ) , .QN( u0_uk_n498 ) );
  DFF_X1 u0_uk_K_r2_reg_53 (.CK( clk ) , .D( u0_uk_K_r1_53 ) , .Q( u0_uk_K_r2_53 ) );
  DFF_X1 u0_uk_K_r2_reg_54 (.CK( clk ) , .D( u0_uk_K_r1_54 ) , .Q( u0_uk_K_r2_54 ) , .QN( u0_uk_n497 ) );
  DFF_X1 u0_uk_K_r2_reg_55 (.CK( clk ) , .D( u0_uk_K_r1_55 ) , .Q( u0_uk_K_r2_55 ) , .QN( u0_uk_n495 ) );
  DFF_X1 u0_uk_K_r2_reg_6 (.CK( clk ) , .D( u0_uk_K_r1_6 ) , .Q( u0_uk_K_r2_6 ) , .QN( u0_uk_n534 ) );
  DFF_X1 u0_uk_K_r2_reg_7 (.CK( clk ) , .D( u0_uk_K_r1_7 ) , .Q( u0_uk_K_r2_7 ) );
  DFF_X1 u0_uk_K_r2_reg_8 (.CK( clk ) , .D( u0_uk_K_r1_8 ) , .Q( u0_uk_K_r2_8 ) , .QN( u0_uk_n533 ) );
  DFF_X1 u0_uk_K_r2_reg_9 (.CK( clk ) , .D( u0_uk_K_r1_9 ) , .Q( u0_uk_K_r2_9 ) , .QN( u0_uk_n532 ) );
  DFF_X1 u0_uk_K_r3_reg_0 (.CK( clk ) , .D( u0_uk_K_r2_0 ) , .Q( u0_uk_K_r3_0 ) , .QN( u0_uk_n494 ) );
  DFF_X1 u0_uk_K_r3_reg_1 (.CK( clk ) , .D( u0_uk_K_r2_1 ) , .Q( u0_uk_K_r3_1 ) , .QN( u0_uk_n493 ) );
  DFF_X1 u0_uk_K_r3_reg_10 (.CK( clk ) , .D( u0_uk_K_r2_10 ) , .Q( u0_uk_K_r3_10 ) );
  DFF_X1 u0_uk_K_r3_reg_11 (.CK( clk ) , .D( u0_uk_K_r2_11 ) , .Q( u0_uk_K_r3_11 ) );
  DFF_X1 u0_uk_K_r3_reg_12 (.CK( clk ) , .D( u0_uk_K_r2_12 ) , .Q( u0_uk_K_r3_12 ) , .QN( u0_uk_n486 ) );
  DFF_X1 u0_uk_K_r3_reg_13 (.CK( clk ) , .D( u0_uk_K_r2_13 ) , .Q( u0_uk_K_r3_13 ) );
  DFF_X1 u0_uk_K_r3_reg_14 (.CK( clk ) , .D( u0_uk_K_r2_14 ) , .Q( u0_uk_K_r3_14 ) );
  DFF_X1 u0_uk_K_r3_reg_15 (.CK( clk ) , .D( u0_uk_K_r2_15 ) , .Q( u0_uk_K_r3_15 ) );
  DFF_X1 u0_uk_K_r3_reg_16 (.CK( clk ) , .D( u0_uk_K_r2_16 ) , .Q( u0_uk_K_r3_16 ) );
  DFF_X1 u0_uk_K_r3_reg_17 (.CK( clk ) , .D( u0_uk_K_r2_17 ) , .Q( u0_uk_K_r3_17 ) , .QN( u0_uk_n485 ) );
  DFF_X1 u0_uk_K_r3_reg_18 (.CK( clk ) , .D( u0_uk_K_r2_18 ) , .Q( u0_uk_K_r3_18 ) , .QN( u0_uk_n484 ) );
  DFF_X1 u0_uk_K_r3_reg_19 (.CK( clk ) , .D( u0_uk_K_r2_19 ) , .Q( u0_uk_K_r3_19 ) );
  DFF_X1 u0_uk_K_r3_reg_2 (.CK( clk ) , .D( u0_uk_K_r2_2 ) , .Q( u0_uk_K_r3_2 ) , .QN( u0_uk_n492 ) );
  DFF_X1 u0_uk_K_r3_reg_20 (.CK( clk ) , .D( u0_uk_K_r2_20 ) , .Q( u0_uk_K_r3_20 ) , .QN( u0_uk_n483 ) );
  DFF_X1 u0_uk_K_r3_reg_21 (.CK( clk ) , .D( u0_uk_K_r2_21 ) , .Q( u0_uk_K_r3_21 ) , .QN( u0_uk_n482 ) );
  DFF_X1 u0_uk_K_r3_reg_22 (.CK( clk ) , .D( u0_uk_K_r2_22 ) , .Q( u0_uk_K_r3_22 ) , .QN( u0_uk_n481 ) );
  DFF_X1 u0_uk_K_r3_reg_23 (.CK( clk ) , .D( u0_uk_K_r2_23 ) , .Q( u0_uk_K_r3_23 ) , .QN( u0_uk_n480 ) );
  DFF_X1 u0_uk_K_r3_reg_24 (.CK( clk ) , .D( u0_uk_K_r2_24 ) , .Q( u0_uk_K_r3_24 ) );
  DFF_X1 u0_uk_K_r3_reg_25 (.CK( clk ) , .D( u0_uk_K_r2_25 ) , .Q( u0_uk_K_r3_25 ) , .QN( u0_uk_n479 ) );
  DFF_X1 u0_uk_K_r3_reg_26 (.CK( clk ) , .D( u0_uk_K_r2_26 ) , .Q( u0_uk_K_r3_26 ) , .QN( u0_uk_n478 ) );
  DFF_X1 u0_uk_K_r3_reg_27 (.CK( clk ) , .D( u0_uk_K_r2_27 ) , .Q( u0_uk_K_r3_27 ) , .QN( u0_uk_n477 ) );
  DFF_X1 u0_uk_K_r3_reg_28 (.CK( clk ) , .D( u0_uk_K_r2_28 ) , .Q( u0_uk_K_r3_28 ) , .QN( u0_uk_n476 ) );
  DFF_X1 u0_uk_K_r3_reg_29 (.CK( clk ) , .D( u0_uk_K_r2_29 ) , .Q( u0_uk_K_r3_29 ) );
  DFF_X1 u0_uk_K_r3_reg_3 (.CK( clk ) , .D( u0_uk_K_r2_3 ) , .Q( u0_uk_K_r3_3 ) , .QN( u0_uk_n491 ) );
  DFF_X1 u0_uk_K_r3_reg_30 (.CK( clk ) , .D( u0_uk_K_r2_30 ) , .Q( u0_uk_K_r3_30 ) , .QN( u0_uk_n475 ) );
  DFF_X1 u0_uk_K_r3_reg_31 (.CK( clk ) , .D( u0_uk_K_r2_31 ) , .Q( u0_uk_K_r3_31 ) , .QN( u0_uk_n474 ) );
  DFF_X1 u0_uk_K_r3_reg_32 (.CK( clk ) , .D( u0_uk_K_r2_32 ) , .Q( u0_uk_K_r3_32 ) , .QN( u0_uk_n473 ) );
  DFF_X1 u0_uk_K_r3_reg_33 (.CK( clk ) , .D( u0_uk_K_r2_33 ) , .Q( u0_uk_K_r3_33 ) , .QN( u0_uk_n471 ) );
  DFF_X1 u0_uk_K_r3_reg_34 (.CK( clk ) , .D( u0_uk_K_r2_34 ) , .Q( u0_uk_K_r3_34 ) );
  DFF_X1 u0_uk_K_r3_reg_35 (.CK( clk ) , .D( u0_uk_K_r2_35 ) , .Q( u0_uk_K_r3_35 ) );
  DFF_X1 u0_uk_K_r3_reg_36 (.CK( clk ) , .D( u0_uk_K_r2_36 ) , .Q( u0_uk_K_r3_36 ) , .QN( u0_uk_n470 ) );
  DFF_X1 u0_uk_K_r3_reg_37 (.CK( clk ) , .D( u0_uk_K_r2_37 ) , .Q( u0_uk_K_r3_37 ) , .QN( u0_uk_n469 ) );
  DFF_X1 u0_uk_K_r3_reg_38 (.CK( clk ) , .D( u0_uk_K_r2_38 ) , .Q( u0_uk_K_r3_38 ) );
  DFF_X1 u0_uk_K_r3_reg_39 (.CK( clk ) , .D( u0_uk_K_r2_39 ) , .Q( u0_uk_K_r3_39 ) , .QN( u0_uk_n466 ) );
  DFF_X1 u0_uk_K_r3_reg_4 (.CK( clk ) , .D( u0_uk_K_r2_4 ) , .Q( u0_uk_K_r3_4 ) );
  DFF_X1 u0_uk_K_r3_reg_40 (.CK( clk ) , .D( u0_uk_K_r2_40 ) , .Q( u0_uk_K_r3_40 ) , .QN( u0_uk_n465 ) );
  DFF_X1 u0_uk_K_r3_reg_41 (.CK( clk ) , .D( u0_uk_K_r2_41 ) , .Q( u0_uk_K_r3_41 ) , .QN( u0_uk_n464 ) );
  DFF_X1 u0_uk_K_r3_reg_42 (.CK( clk ) , .D( u0_uk_K_r2_42 ) , .Q( u0_uk_K_r3_42 ) , .QN( u0_uk_n463 ) );
  DFF_X1 u0_uk_K_r3_reg_43 (.CK( clk ) , .D( u0_uk_K_r2_43 ) , .Q( u0_uk_K_r3_43 ) );
  DFF_X1 u0_uk_K_r3_reg_44 (.CK( clk ) , .D( u0_uk_K_r2_44 ) , .Q( u0_uk_K_r3_44 ) );
  DFF_X1 u0_uk_K_r3_reg_45 (.CK( clk ) , .D( u0_uk_K_r2_45 ) , .Q( u0_uk_K_r3_45 ) , .QN( u0_uk_n462 ) );
  DFF_X1 u0_uk_K_r3_reg_46 (.CK( clk ) , .D( u0_uk_K_r2_46 ) , .Q( u0_uk_K_r3_46 ) , .QN( u0_uk_n461 ) );
  DFF_X1 u0_uk_K_r3_reg_47 (.CK( clk ) , .D( u0_uk_K_r2_47 ) , .Q( u0_uk_K_r3_47 ) );
  DFF_X1 u0_uk_K_r3_reg_48 (.CK( clk ) , .D( u0_uk_K_r2_48 ) , .Q( u0_uk_K_r3_48 ) , .QN( u0_uk_n459 ) );
  DFF_X1 u0_uk_K_r3_reg_49 (.CK( clk ) , .D( u0_uk_K_r2_49 ) , .Q( u0_uk_K_r3_49 ) , .QN( u0_uk_n458 ) );
  DFF_X1 u0_uk_K_r3_reg_5 (.CK( clk ) , .D( u0_uk_K_r2_5 ) , .Q( u0_uk_K_r3_5 ) , .QN( u0_uk_n490 ) );
  DFF_X1 u0_uk_K_r3_reg_50 (.CK( clk ) , .D( u0_uk_K_r2_50 ) , .Q( u0_uk_K_r3_50 ) , .QN( u0_uk_n457 ) );
  DFF_X1 u0_uk_K_r3_reg_51 (.CK( clk ) , .D( u0_uk_K_r2_51 ) , .Q( u0_uk_K_r3_51 ) , .QN( u0_uk_n455 ) );
  DFF_X1 u0_uk_K_r3_reg_52 (.CK( clk ) , .D( u0_uk_K_r2_52 ) , .Q( u0_uk_K_r3_52 ) );
  DFF_X1 u0_uk_K_r3_reg_53 (.CK( clk ) , .D( u0_uk_K_r2_53 ) , .Q( u0_uk_K_r3_53 ) , .QN( u0_uk_n453 ) );
  DFF_X1 u0_uk_K_r3_reg_54 (.CK( clk ) , .D( u0_uk_K_r2_54 ) , .Q( u0_uk_K_r3_54 ) , .QN( u0_uk_n452 ) );
  DFF_X1 u0_uk_K_r3_reg_55 (.CK( clk ) , .D( u0_uk_K_r2_55 ) , .Q( u0_uk_K_r3_55 ) , .QN( u0_uk_n451 ) );
  DFF_X1 u0_uk_K_r3_reg_6 (.CK( clk ) , .D( u0_uk_K_r2_6 ) , .Q( u0_uk_K_r3_6 ) , .QN( u0_uk_n489 ) );
  DFF_X1 u0_uk_K_r3_reg_7 (.CK( clk ) , .D( u0_uk_K_r2_7 ) , .Q( u0_uk_K_r3_7 ) , .QN( u0_uk_n488 ) );
  DFF_X1 u0_uk_K_r3_reg_8 (.CK( clk ) , .D( u0_uk_K_r2_8 ) , .Q( u0_uk_K_r3_8 ) , .QN( u0_uk_n487 ) );
  DFF_X1 u0_uk_K_r3_reg_9 (.CK( clk ) , .D( u0_uk_K_r2_9 ) , .Q( u0_uk_K_r3_9 ) );
  DFF_X1 u0_uk_K_r4_reg_0 (.CK( clk ) , .D( u0_uk_K_r3_0 ) , .Q( u0_uk_K_r4_0 ) );
  DFF_X1 u0_uk_K_r4_reg_1 (.CK( clk ) , .D( u0_uk_K_r3_1 ) , .Q( u0_uk_K_r4_1 ) , .QN( u0_uk_n450 ) );
  DFF_X1 u0_uk_K_r4_reg_10 (.CK( clk ) , .D( u0_uk_K_r3_10 ) , .Q( u0_uk_K_r4_10 ) , .QN( u0_uk_n444 ) );
  DFF_X1 u0_uk_K_r4_reg_11 (.CK( clk ) , .D( u0_uk_K_r3_11 ) , .Q( u0_uk_K_r4_11 ) );
  DFF_X1 u0_uk_K_r4_reg_12 (.CK( clk ) , .D( u0_uk_K_r3_12 ) , .Q( u0_uk_K_r4_12 ) , .QN( u0_uk_n442 ) );
  DFF_X1 u0_uk_K_r4_reg_13 (.CK( clk ) , .D( u0_uk_K_r3_13 ) , .Q( u0_uk_K_r4_13 ) , .QN( u0_uk_n441 ) );
  DFF_X1 u0_uk_K_r4_reg_14 (.CK( clk ) , .D( u0_uk_K_r3_14 ) , .Q( u0_uk_K_r4_14 ) , .QN( u0_uk_n440 ) );
  DFF_X1 u0_uk_K_r4_reg_15 (.CK( clk ) , .D( u0_uk_K_r3_15 ) , .Q( u0_uk_K_r4_15 ) , .QN( u0_uk_n439 ) );
  DFF_X1 u0_uk_K_r4_reg_16 (.CK( clk ) , .D( u0_uk_K_r3_16 ) , .Q( u0_uk_K_r4_16 ) , .QN( u0_uk_n438 ) );
  DFF_X1 u0_uk_K_r4_reg_17 (.CK( clk ) , .D( u0_uk_K_r3_17 ) , .Q( u0_uk_K_r4_17 ) );
  DFF_X1 u0_uk_K_r4_reg_18 (.CK( clk ) , .D( u0_uk_K_r3_18 ) , .Q( u0_uk_K_r4_18 ) );
  DFF_X1 u0_uk_K_r4_reg_19 (.CK( clk ) , .D( u0_uk_K_r3_19 ) , .Q( u0_uk_K_r4_19 ) , .QN( u0_uk_n436 ) );
  DFF_X1 u0_uk_K_r4_reg_2 (.CK( clk ) , .D( u0_uk_K_r3_2 ) , .Q( u0_uk_K_r4_2 ) );
  DFF_X1 u0_uk_K_r4_reg_20 (.CK( clk ) , .D( u0_uk_K_r3_20 ) , .Q( u0_uk_K_r4_20 ) , .QN( u0_uk_n435 ) );
  DFF_X1 u0_uk_K_r4_reg_21 (.CK( clk ) , .D( u0_uk_K_r3_21 ) , .Q( u0_uk_K_r4_21 ) , .QN( u0_uk_n434 ) );
  DFF_X1 u0_uk_K_r4_reg_22 (.CK( clk ) , .D( u0_uk_K_r3_22 ) , .Q( u0_uk_K_r4_22 ) , .QN( u0_uk_n433 ) );
  DFF_X1 u0_uk_K_r4_reg_23 (.CK( clk ) , .D( u0_uk_K_r3_23 ) , .Q( u0_uk_K_r4_23 ) );
  DFF_X1 u0_uk_K_r4_reg_24 (.CK( clk ) , .D( u0_uk_K_r3_24 ) , .Q( u0_uk_K_r4_24 ) );
  DFF_X1 u0_uk_K_r4_reg_25 (.CK( clk ) , .D( u0_uk_K_r3_25 ) , .Q( u0_uk_K_r4_25 ) , .QN( u0_uk_n432 ) );
  DFF_X1 u0_uk_K_r4_reg_26 (.CK( clk ) , .D( u0_uk_K_r3_26 ) , .Q( u0_uk_K_r4_26 ) , .QN( u0_uk_n431 ) );
  DFF_X1 u0_uk_K_r4_reg_27 (.CK( clk ) , .D( u0_uk_K_r3_27 ) , .Q( u0_uk_K_r4_27 ) );
  DFF_X1 u0_uk_K_r4_reg_28 (.CK( clk ) , .D( u0_uk_K_r3_28 ) , .Q( u0_uk_K_r4_28 ) , .QN( u0_uk_n430 ) );
  DFF_X1 u0_uk_K_r4_reg_29 (.CK( clk ) , .D( u0_uk_K_r3_29 ) , .Q( u0_uk_K_r4_29 ) , .QN( u0_uk_n429 ) );
  DFF_X1 u0_uk_K_r4_reg_3 (.CK( clk ) , .D( u0_uk_K_r3_3 ) , .Q( u0_uk_K_r4_3 ) );
  DFF_X1 u0_uk_K_r4_reg_30 (.CK( clk ) , .D( u0_uk_K_r3_30 ) , .Q( u0_uk_K_r4_30 ) , .QN( u0_uk_n428 ) );
  DFF_X1 u0_uk_K_r4_reg_31 (.CK( clk ) , .D( u0_uk_K_r3_31 ) , .Q( u0_uk_K_r4_31 ) );
  DFF_X1 u0_uk_K_r4_reg_32 (.CK( clk ) , .D( u0_uk_K_r3_32 ) , .Q( u0_uk_K_r4_32 ) , .QN( u0_uk_n427 ) );
  DFF_X1 u0_uk_K_r4_reg_33 (.CK( clk ) , .D( u0_uk_K_r3_33 ) , .Q( u0_uk_K_r4_33 ) );
  DFF_X1 u0_uk_K_r4_reg_34 (.CK( clk ) , .D( u0_uk_K_r3_34 ) , .Q( u0_uk_K_r4_34 ) , .QN( u0_uk_n426 ) );
  DFF_X1 u0_uk_K_r4_reg_35 (.CK( clk ) , .D( u0_uk_K_r3_35 ) , .Q( u0_uk_K_r4_35 ) );
  DFF_X1 u0_uk_K_r4_reg_36 (.CK( clk ) , .D( u0_uk_K_r3_36 ) , .Q( u0_uk_K_r4_36 ) , .QN( u0_uk_n425 ) );
  DFF_X1 u0_uk_K_r4_reg_37 (.CK( clk ) , .D( u0_uk_K_r3_37 ) , .Q( u0_uk_K_r4_37 ) , .QN( u0_uk_n424 ) );
  DFF_X1 u0_uk_K_r4_reg_38 (.CK( clk ) , .D( u0_uk_K_r3_38 ) , .Q( u0_uk_K_r4_38 ) );
  DFF_X1 u0_uk_K_r4_reg_39 (.CK( clk ) , .D( u0_uk_K_r3_39 ) , .Q( u0_uk_K_r4_39 ) , .QN( u0_uk_n423 ) );
  DFF_X1 u0_uk_K_r4_reg_4 (.CK( clk ) , .D( u0_uk_K_r3_4 ) , .Q( u0_uk_K_r4_4 ) , .QN( u0_uk_n449 ) );
  DFF_X1 u0_uk_K_r4_reg_40 (.CK( clk ) , .D( u0_uk_K_r3_40 ) , .Q( u0_uk_K_r4_40 ) , .QN( u0_uk_n422 ) );
  DFF_X1 u0_uk_K_r4_reg_41 (.CK( clk ) , .D( u0_uk_K_r3_41 ) , .Q( u0_uk_K_r4_41 ) );
  DFF_X1 u0_uk_K_r4_reg_42 (.CK( clk ) , .D( u0_uk_K_r3_42 ) , .Q( u0_uk_K_r4_42 ) , .QN( u0_uk_n420 ) );
  DFF_X1 u0_uk_K_r4_reg_43 (.CK( clk ) , .D( u0_uk_K_r3_43 ) , .Q( u0_uk_K_r4_43 ) , .QN( u0_uk_n419 ) );
  DFF_X1 u0_uk_K_r4_reg_44 (.CK( clk ) , .D( u0_uk_K_r3_44 ) , .Q( u0_uk_K_r4_44 ) , .QN( u0_uk_n418 ) );
  DFF_X1 u0_uk_K_r4_reg_45 (.CK( clk ) , .D( u0_uk_K_r3_45 ) , .Q( u0_uk_K_r4_45 ) , .QN( u0_uk_n417 ) );
  DFF_X1 u0_uk_K_r4_reg_46 (.CK( clk ) , .D( u0_uk_K_r3_46 ) , .Q( u0_uk_K_r4_46 ) , .QN( u0_uk_n416 ) );
  DFF_X1 u0_uk_K_r4_reg_47 (.CK( clk ) , .D( u0_uk_K_r3_47 ) , .Q( u0_uk_K_r4_47 ) , .QN( u0_uk_n414 ) );
  DFF_X1 u0_uk_K_r4_reg_48 (.CK( clk ) , .D( u0_uk_K_r3_48 ) , .Q( u0_uk_K_r4_48 ) );
  DFF_X1 u0_uk_K_r4_reg_49 (.CK( clk ) , .D( u0_uk_K_r3_49 ) , .Q( u0_uk_K_r4_49 ) );
  DFF_X1 u0_uk_K_r4_reg_5 (.CK( clk ) , .D( u0_uk_K_r3_5 ) , .Q( u0_uk_K_r4_5 ) );
  DFF_X1 u0_uk_K_r4_reg_50 (.CK( clk ) , .D( u0_uk_K_r3_50 ) , .Q( u0_uk_K_r4_50 ) , .QN( u0_uk_n413 ) );
  DFF_X1 u0_uk_K_r4_reg_51 (.CK( clk ) , .D( u0_uk_K_r3_51 ) , .Q( u0_uk_K_r4_51 ) , .QN( u0_uk_n412 ) );
  DFF_X1 u0_uk_K_r4_reg_52 (.CK( clk ) , .D( u0_uk_K_r3_52 ) , .Q( u0_uk_K_r4_52 ) , .QN( u0_uk_n411 ) );
  DFF_X1 u0_uk_K_r4_reg_53 (.CK( clk ) , .D( u0_uk_K_r3_53 ) , .Q( u0_uk_K_r4_53 ) , .QN( u0_uk_n410 ) );
  DFF_X1 u0_uk_K_r4_reg_54 (.CK( clk ) , .D( u0_uk_K_r3_54 ) , .Q( u0_uk_K_r4_54 ) );
  DFF_X1 u0_uk_K_r4_reg_55 (.CK( clk ) , .D( u0_uk_K_r3_55 ) , .Q( u0_uk_K_r4_55 ) );
  DFF_X1 u0_uk_K_r4_reg_6 (.CK( clk ) , .D( u0_uk_K_r3_6 ) , .Q( u0_uk_K_r4_6 ) , .QN( u0_uk_n448 ) );
  DFF_X1 u0_uk_K_r4_reg_7 (.CK( clk ) , .D( u0_uk_K_r3_7 ) , .Q( u0_uk_K_r4_7 ) , .QN( u0_uk_n447 ) );
  DFF_X1 u0_uk_K_r4_reg_8 (.CK( clk ) , .D( u0_uk_K_r3_8 ) , .Q( u0_uk_K_r4_8 ) , .QN( u0_uk_n446 ) );
  DFF_X1 u0_uk_K_r4_reg_9 (.CK( clk ) , .D( u0_uk_K_r3_9 ) , .Q( u0_uk_K_r4_9 ) , .QN( u0_uk_n445 ) );
  DFF_X1 u0_uk_K_r5_reg_0 (.CK( clk ) , .D( u0_uk_K_r4_0 ) , .Q( u0_uk_K_r5_0 ) );
  DFF_X1 u0_uk_K_r5_reg_1 (.CK( clk ) , .D( u0_uk_K_r4_1 ) , .Q( u0_uk_K_r5_1 ) );
  DFF_X1 u0_uk_K_r5_reg_10 (.CK( clk ) , .D( u0_uk_K_r4_10 ) , .Q( u0_uk_K_r5_10 ) );
  DFF_X1 u0_uk_K_r5_reg_11 (.CK( clk ) , .D( u0_uk_K_r4_11 ) , .Q( u0_uk_K_r5_11 ) , .QN( u0_uk_n401 ) );
  DFF_X1 u0_uk_K_r5_reg_12 (.CK( clk ) , .D( u0_uk_K_r4_12 ) , .Q( u0_uk_K_r5_12 ) , .QN( u0_uk_n400 ) );
  DFF_X1 u0_uk_K_r5_reg_13 (.CK( clk ) , .D( u0_uk_K_r4_13 ) , .Q( u0_uk_K_r5_13 ) );
  DFF_X1 u0_uk_K_r5_reg_14 (.CK( clk ) , .D( u0_uk_K_r4_14 ) , .Q( u0_uk_K_r5_14 ) , .QN( u0_uk_n399 ) );
  DFF_X1 u0_uk_K_r5_reg_15 (.CK( clk ) , .D( u0_uk_K_r4_15 ) , .Q( u0_uk_K_r5_15 ) , .QN( u0_uk_n398 ) );
  DFF_X1 u0_uk_K_r5_reg_16 (.CK( clk ) , .D( u0_uk_K_r4_16 ) , .Q( u0_uk_K_r5_16 ) );
  DFF_X1 u0_uk_K_r5_reg_17 (.CK( clk ) , .D( u0_uk_K_r4_17 ) , .Q( u0_uk_K_r5_17 ) , .QN( u0_uk_n397 ) );
  DFF_X1 u0_uk_K_r5_reg_18 (.CK( clk ) , .D( u0_uk_K_r4_18 ) , .Q( u0_uk_K_r5_18 ) );
  DFF_X1 u0_uk_K_r5_reg_19 (.CK( clk ) , .D( u0_uk_K_r4_19 ) , .Q( u0_uk_K_r5_19 ) );
  DFF_X1 u0_uk_K_r5_reg_2 (.CK( clk ) , .D( u0_uk_K_r4_2 ) , .Q( u0_uk_K_r5_2 ) , .QN( u0_uk_n406 ) );
  DFF_X1 u0_uk_K_r5_reg_20 (.CK( clk ) , .D( u0_uk_K_r4_20 ) , .Q( u0_uk_K_r5_20 ) , .QN( u0_uk_n396 ) );
  DFF_X1 u0_uk_K_r5_reg_21 (.CK( clk ) , .D( u0_uk_K_r4_21 ) , .Q( u0_uk_K_r5_21 ) );
  DFF_X1 u0_uk_K_r5_reg_22 (.CK( clk ) , .D( u0_uk_K_r4_22 ) , .Q( u0_uk_K_r5_22 ) , .QN( u0_uk_n394 ) );
  DFF_X1 u0_uk_K_r5_reg_23 (.CK( clk ) , .D( u0_uk_K_r4_23 ) , .Q( u0_uk_K_r5_23 ) );
  DFF_X1 u0_uk_K_r5_reg_24 (.CK( clk ) , .D( u0_uk_K_r4_24 ) , .Q( u0_uk_K_r5_24 ) , .QN( u0_uk_n393 ) );
  DFF_X1 u0_uk_K_r5_reg_25 (.CK( clk ) , .D( u0_uk_K_r4_25 ) , .Q( u0_uk_K_r5_25 ) , .QN( u0_uk_n392 ) );
  DFF_X1 u0_uk_K_r5_reg_26 (.CK( clk ) , .D( u0_uk_K_r4_26 ) , .Q( u0_uk_K_r5_26 ) );
  DFF_X1 u0_uk_K_r5_reg_27 (.CK( clk ) , .D( u0_uk_K_r4_27 ) , .Q( u0_uk_K_r5_27 ) , .QN( u0_uk_n390 ) );
  DFF_X1 u0_uk_K_r5_reg_28 (.CK( clk ) , .D( u0_uk_K_r4_28 ) , .Q( u0_uk_K_r5_28 ) , .QN( u0_uk_n389 ) );
  DFF_X1 u0_uk_K_r5_reg_29 (.CK( clk ) , .D( u0_uk_K_r4_29 ) , .Q( u0_uk_K_r5_29 ) , .QN( u0_uk_n388 ) );
  DFF_X1 u0_uk_K_r5_reg_3 (.CK( clk ) , .D( u0_uk_K_r4_3 ) , .Q( u0_uk_K_r5_3 ) , .QN( u0_uk_n405 ) );
  DFF_X1 u0_uk_K_r5_reg_30 (.CK( clk ) , .D( u0_uk_K_r4_30 ) , .Q( u0_uk_K_r5_30 ) , .QN( u0_uk_n387 ) );
  DFF_X1 u0_uk_K_r5_reg_31 (.CK( clk ) , .D( u0_uk_K_r4_31 ) , .Q( u0_uk_K_r5_31 ) );
  DFF_X1 u0_uk_K_r5_reg_32 (.CK( clk ) , .D( u0_uk_K_r4_32 ) , .Q( u0_uk_K_r5_32 ) );
  DFF_X1 u0_uk_K_r5_reg_33 (.CK( clk ) , .D( u0_uk_K_r4_33 ) , .Q( u0_uk_K_r5_33 ) , .QN( u0_uk_n384 ) );
  DFF_X1 u0_uk_K_r5_reg_34 (.CK( clk ) , .D( u0_uk_K_r4_34 ) , .Q( u0_uk_K_r5_34 ) , .QN( u0_uk_n383 ) );
  DFF_X1 u0_uk_K_r5_reg_35 (.CK( clk ) , .D( u0_uk_K_r4_35 ) , .Q( u0_uk_K_r5_35 ) , .QN( u0_uk_n381 ) );
  DFF_X1 u0_uk_K_r5_reg_36 (.CK( clk ) , .D( u0_uk_K_r4_36 ) , .Q( u0_uk_K_r5_36 ) , .QN( u0_uk_n380 ) );
  DFF_X1 u0_uk_K_r5_reg_37 (.CK( clk ) , .D( u0_uk_K_r4_37 ) , .Q( u0_uk_K_r5_37 ) );
  DFF_X1 u0_uk_K_r5_reg_38 (.CK( clk ) , .D( u0_uk_K_r4_38 ) , .Q( u0_uk_K_r5_38 ) , .QN( u0_uk_n378 ) );
  DFF_X1 u0_uk_K_r5_reg_39 (.CK( clk ) , .D( u0_uk_K_r4_39 ) , .Q( u0_uk_K_r5_39 ) );
  DFF_X1 u0_uk_K_r5_reg_4 (.CK( clk ) , .D( u0_uk_K_r4_4 ) , .Q( u0_uk_K_r5_4 ) );
  DFF_X1 u0_uk_K_r5_reg_40 (.CK( clk ) , .D( u0_uk_K_r4_40 ) , .Q( u0_uk_K_r5_40 ) );
  DFF_X1 u0_uk_K_r5_reg_41 (.CK( clk ) , .D( u0_uk_K_r4_41 ) , .Q( u0_uk_K_r5_41 ) );
  DFF_X1 u0_uk_K_r5_reg_42 (.CK( clk ) , .D( u0_uk_K_r4_42 ) , .Q( u0_uk_K_r5_42 ) , .QN( u0_uk_n374 ) );
  DFF_X1 u0_uk_K_r5_reg_43 (.CK( clk ) , .D( u0_uk_K_r4_43 ) , .Q( u0_uk_K_r5_43 ) );
  DFF_X1 u0_uk_K_r5_reg_44 (.CK( clk ) , .D( u0_uk_K_r4_44 ) , .Q( u0_uk_K_r5_44 ) , .QN( u0_uk_n372 ) );
  DFF_X1 u0_uk_K_r5_reg_45 (.CK( clk ) , .D( u0_uk_K_r4_45 ) , .Q( u0_uk_K_r5_45 ) );
  DFF_X1 u0_uk_K_r5_reg_46 (.CK( clk ) , .D( u0_uk_K_r4_46 ) , .Q( u0_uk_K_r5_46 ) , .QN( u0_uk_n371 ) );
  DFF_X1 u0_uk_K_r5_reg_47 (.CK( clk ) , .D( u0_uk_K_r4_47 ) , .Q( u0_uk_K_r5_47 ) , .QN( u0_uk_n370 ) );
  DFF_X1 u0_uk_K_r5_reg_48 (.CK( clk ) , .D( u0_uk_K_r4_48 ) , .Q( u0_uk_K_r5_48 ) );
  DFF_X1 u0_uk_K_r5_reg_49 (.CK( clk ) , .D( u0_uk_K_r4_49 ) , .Q( u0_uk_K_r5_49 ) , .QN( u0_uk_n368 ) );
  DFF_X1 u0_uk_K_r5_reg_5 (.CK( clk ) , .D( u0_uk_K_r4_5 ) , .Q( u0_uk_K_r5_5 ) );
  DFF_X1 u0_uk_K_r5_reg_50 (.CK( clk ) , .D( u0_uk_K_r4_50 ) , .Q( u0_uk_K_r5_50 ) , .QN( u0_uk_n367 ) );
  DFF_X1 u0_uk_K_r5_reg_51 (.CK( clk ) , .D( u0_uk_K_r4_51 ) , .Q( u0_uk_K_r5_51 ) );
  DFF_X1 u0_uk_K_r5_reg_52 (.CK( clk ) , .D( u0_uk_K_r4_52 ) , .Q( u0_uk_K_r5_52 ) , .QN( u0_uk_n365 ) );
  DFF_X1 u0_uk_K_r5_reg_53 (.CK( clk ) , .D( u0_uk_K_r4_53 ) , .Q( u0_uk_K_r5_53 ) , .QN( u0_uk_n364 ) );
  DFF_X1 u0_uk_K_r5_reg_54 (.CK( clk ) , .D( u0_uk_K_r4_54 ) , .Q( u0_uk_K_r5_54 ) , .QN( u0_uk_n362 ) );
  DFF_X1 u0_uk_K_r5_reg_55 (.CK( clk ) , .D( u0_uk_K_r4_55 ) , .Q( u0_uk_K_r5_55 ) , .QN( u0_uk_n361 ) );
  DFF_X1 u0_uk_K_r5_reg_6 (.CK( clk ) , .D( u0_uk_K_r4_6 ) , .Q( u0_uk_K_r5_6 ) , .QN( u0_uk_n404 ) );
  DFF_X1 u0_uk_K_r5_reg_7 (.CK( clk ) , .D( u0_uk_K_r4_7 ) , .Q( u0_uk_K_r5_7 ) , .QN( u0_uk_n403 ) );
  DFF_X1 u0_uk_K_r5_reg_8 (.CK( clk ) , .D( u0_uk_K_r4_8 ) , .Q( u0_uk_K_r5_8 ) );
  DFF_X1 u0_uk_K_r5_reg_9 (.CK( clk ) , .D( u0_uk_K_r4_9 ) , .Q( u0_uk_K_r5_9 ) , .QN( u0_uk_n402 ) );
  DFF_X1 u0_uk_K_r6_reg_0 (.CK( clk ) , .D( u0_uk_K_r5_0 ) , .Q( u0_uk_K_r6_0 ) );
  DFF_X1 u0_uk_K_r6_reg_1 (.CK( clk ) , .D( u0_uk_K_r5_1 ) , .Q( u0_uk_K_r6_1 ) , .QN( u0_uk_n360 ) );
  DFF_X1 u0_uk_K_r6_reg_10 (.CK( clk ) , .D( u0_uk_K_r5_10 ) , .Q( u0_uk_K_r6_10 ) );
  DFF_X1 u0_uk_K_r6_reg_11 (.CK( clk ) , .D( u0_uk_K_r5_11 ) , .Q( u0_uk_K_r6_11 ) , .QN( u0_uk_n352 ) );
  DFF_X1 u0_uk_K_r6_reg_12 (.CK( clk ) , .D( u0_uk_K_r5_12 ) , .Q( u0_uk_K_r6_12 ) , .QN( u0_uk_n351 ) );
  DFF_X1 u0_uk_K_r6_reg_13 (.CK( clk ) , .D( u0_uk_K_r5_13 ) , .Q( u0_uk_K_r6_13 ) , .QN( u0_uk_n350 ) );
  DFF_X1 u0_uk_K_r6_reg_14 (.CK( clk ) , .D( u0_uk_K_r5_14 ) , .Q( u0_uk_K_r6_14 ) );
  DFF_X1 u0_uk_K_r6_reg_15 (.CK( clk ) , .D( u0_uk_K_r5_15 ) , .Q( u0_uk_K_r6_15 ) , .QN( u0_uk_n348 ) );
  DFF_X1 u0_uk_K_r6_reg_16 (.CK( clk ) , .D( u0_uk_K_r5_16 ) , .Q( u0_uk_K_r6_16 ) , .QN( u0_uk_n347 ) );
  DFF_X1 u0_uk_K_r6_reg_17 (.CK( clk ) , .D( u0_uk_K_r5_17 ) , .Q( u0_uk_K_r6_17 ) , .QN( u0_uk_n345 ) );
  DFF_X1 u0_uk_K_r6_reg_18 (.CK( clk ) , .D( u0_uk_K_r5_18 ) , .Q( u0_uk_K_r6_18 ) , .QN( u0_uk_n344 ) );
  DFF_X1 u0_uk_K_r6_reg_19 (.CK( clk ) , .D( u0_uk_K_r5_19 ) , .Q( u0_uk_K_r6_19 ) );
  DFF_X1 u0_uk_K_r6_reg_2 (.CK( clk ) , .D( u0_uk_K_r5_2 ) , .Q( u0_uk_K_r6_2 ) , .QN( u0_uk_n359 ) );
  DFF_X1 u0_uk_K_r6_reg_20 (.CK( clk ) , .D( u0_uk_K_r5_20 ) , .Q( u0_uk_K_r6_20 ) , .QN( u0_uk_n343 ) );
  DFF_X1 u0_uk_K_r6_reg_21 (.CK( clk ) , .D( u0_uk_K_r5_21 ) , .Q( u0_uk_K_r6_21 ) );
  DFF_X1 u0_uk_K_r6_reg_22 (.CK( clk ) , .D( u0_uk_K_r5_22 ) , .Q( u0_uk_K_r6_22 ) );
  DFF_X1 u0_uk_K_r6_reg_23 (.CK( clk ) , .D( u0_uk_K_r5_23 ) , .Q( u0_uk_K_r6_23 ) , .QN( u0_uk_n341 ) );
  DFF_X1 u0_uk_K_r6_reg_24 (.CK( clk ) , .D( u0_uk_K_r5_24 ) , .Q( u0_uk_K_r6_24 ) , .QN( u0_uk_n340 ) );
  DFF_X1 u0_uk_K_r6_reg_25 (.CK( clk ) , .D( u0_uk_K_r5_25 ) , .Q( u0_uk_K_r6_25 ) , .QN( u0_uk_n339 ) );
  DFF_X1 u0_uk_K_r6_reg_26 (.CK( clk ) , .D( u0_uk_K_r5_26 ) , .Q( u0_uk_K_r6_26 ) );
  DFF_X1 u0_uk_K_r6_reg_27 (.CK( clk ) , .D( u0_uk_K_r5_27 ) , .Q( u0_uk_K_r6_27 ) );
  DFF_X1 u0_uk_K_r6_reg_28 (.CK( clk ) , .D( u0_uk_K_r5_28 ) , .Q( u0_uk_K_r6_28 ) );
  DFF_X1 u0_uk_K_r6_reg_29 (.CK( clk ) , .D( u0_uk_K_r5_29 ) , .Q( u0_uk_K_r6_29 ) );
  DFF_X1 u0_uk_K_r6_reg_3 (.CK( clk ) , .D( u0_uk_K_r5_3 ) , .Q( u0_uk_K_r6_3 ) );
  DFF_X1 u0_uk_K_r6_reg_30 (.CK( clk ) , .D( u0_uk_K_r5_30 ) , .Q( u0_uk_K_r6_30 ) );
  DFF_X1 u0_uk_K_r6_reg_31 (.CK( clk ) , .D( u0_uk_K_r5_31 ) , .Q( u0_uk_K_r6_31 ) );
  DFF_X1 u0_uk_K_r6_reg_32 (.CK( clk ) , .D( u0_uk_K_r5_32 ) , .Q( u0_uk_K_r6_32 ) , .QN( u0_uk_n337 ) );
  DFF_X1 u0_uk_K_r6_reg_33 (.CK( clk ) , .D( u0_uk_K_r5_33 ) , .Q( u0_uk_K_r6_33 ) , .QN( u0_uk_n336 ) );
  DFF_X1 u0_uk_K_r6_reg_34 (.CK( clk ) , .D( u0_uk_K_r5_34 ) , .Q( u0_uk_K_r6_34 ) );
  DFF_X1 u0_uk_K_r6_reg_35 (.CK( clk ) , .D( u0_uk_K_r5_35 ) , .Q( u0_uk_K_r6_35 ) , .QN( u0_uk_n334 ) );
  DFF_X1 u0_uk_K_r6_reg_36 (.CK( clk ) , .D( u0_uk_K_r5_36 ) , .Q( u0_uk_K_r6_36 ) , .QN( u0_uk_n333 ) );
  DFF_X1 u0_uk_K_r6_reg_37 (.CK( clk ) , .D( u0_uk_K_r5_37 ) , .Q( u0_uk_K_r6_37 ) );
  DFF_X1 u0_uk_K_r6_reg_38 (.CK( clk ) , .D( u0_uk_K_r5_38 ) , .Q( u0_uk_K_r6_38 ) , .QN( u0_uk_n332 ) );
  DFF_X1 u0_uk_K_r6_reg_39 (.CK( clk ) , .D( u0_uk_K_r5_39 ) , .Q( u0_uk_K_r6_39 ) , .QN( u0_uk_n331 ) );
  DFF_X1 u0_uk_K_r6_reg_4 (.CK( clk ) , .D( u0_uk_K_r5_4 ) , .Q( u0_uk_K_r6_4 ) , .QN( u0_uk_n358 ) );
  DFF_X1 u0_uk_K_r6_reg_40 (.CK( clk ) , .D( u0_uk_K_r5_40 ) , .Q( u0_uk_K_r6_40 ) , .QN( u0_uk_n330 ) );
  DFF_X1 u0_uk_K_r6_reg_41 (.CK( clk ) , .D( u0_uk_K_r5_41 ) , .Q( u0_uk_K_r6_41 ) , .QN( u0_uk_n329 ) );
  DFF_X1 u0_uk_K_r6_reg_42 (.CK( clk ) , .D( u0_uk_K_r5_42 ) , .Q( u0_uk_K_r6_42 ) , .QN( u0_uk_n328 ) );
  DFF_X1 u0_uk_K_r6_reg_43 (.CK( clk ) , .D( u0_uk_K_r5_43 ) , .Q( u0_uk_K_r6_43 ) , .QN( u0_uk_n327 ) );
  DFF_X1 u0_uk_K_r6_reg_44 (.CK( clk ) , .D( u0_uk_K_r5_44 ) , .Q( u0_uk_K_r6_44 ) , .QN( u0_uk_n326 ) );
  DFF_X1 u0_uk_K_r6_reg_45 (.CK( clk ) , .D( u0_uk_K_r5_45 ) , .Q( u0_uk_K_r6_45 ) , .QN( u0_uk_n325 ) );
  DFF_X1 u0_uk_K_r6_reg_46 (.CK( clk ) , .D( u0_uk_K_r5_46 ) , .Q( u0_uk_K_r6_46 ) );
  DFF_X1 u0_uk_K_r6_reg_47 (.CK( clk ) , .D( u0_uk_K_r5_47 ) , .Q( u0_uk_K_r6_47 ) , .QN( u0_uk_n324 ) );
  DFF_X1 u0_uk_K_r6_reg_48 (.CK( clk ) , .D( u0_uk_K_r5_48 ) , .Q( u0_uk_K_r6_48 ) , .QN( u0_uk_n323 ) );
  DFF_X1 u0_uk_K_r6_reg_49 (.CK( clk ) , .D( u0_uk_K_r5_49 ) , .Q( u0_uk_K_r6_49 ) , .QN( u0_uk_n322 ) );
  DFF_X1 u0_uk_K_r6_reg_5 (.CK( clk ) , .D( u0_uk_K_r5_5 ) , .Q( u0_uk_K_r6_5 ) , .QN( u0_uk_n357 ) );
  DFF_X1 u0_uk_K_r6_reg_50 (.CK( clk ) , .D( u0_uk_K_r5_50 ) , .Q( u0_uk_K_r6_50 ) , .QN( u0_uk_n321 ) );
  DFF_X1 u0_uk_K_r6_reg_51 (.CK( clk ) , .D( u0_uk_K_r5_51 ) , .Q( u0_uk_K_r6_51 ) );
  DFF_X1 u0_uk_K_r6_reg_52 (.CK( clk ) , .D( u0_uk_K_r5_52 ) , .Q( u0_uk_K_r6_52 ) , .QN( u0_uk_n320 ) );
  DFF_X1 u0_uk_K_r6_reg_53 (.CK( clk ) , .D( u0_uk_K_r5_53 ) , .Q( u0_uk_K_r6_53 ) );
  DFF_X1 u0_uk_K_r6_reg_54 (.CK( clk ) , .D( u0_uk_K_r5_54 ) , .Q( u0_uk_K_r6_54 ) , .QN( u0_uk_n318 ) );
  DFF_X1 u0_uk_K_r6_reg_55 (.CK( clk ) , .D( u0_uk_K_r5_55 ) , .Q( u0_uk_K_r6_55 ) );
  DFF_X1 u0_uk_K_r6_reg_6 (.CK( clk ) , .D( u0_uk_K_r5_6 ) , .Q( u0_uk_K_r6_6 ) , .QN( u0_uk_n356 ) );
  DFF_X1 u0_uk_K_r6_reg_7 (.CK( clk ) , .D( u0_uk_K_r5_7 ) , .Q( u0_uk_K_r6_7 ) );
  DFF_X1 u0_uk_K_r6_reg_8 (.CK( clk ) , .D( u0_uk_K_r5_8 ) , .Q( u0_uk_K_r6_8 ) , .QN( u0_uk_n355 ) );
  DFF_X1 u0_uk_K_r6_reg_9 (.CK( clk ) , .D( u0_uk_K_r5_9 ) , .Q( u0_uk_K_r6_9 ) , .QN( u0_uk_n354 ) );
  DFF_X1 u0_uk_K_r7_reg_0 (.CK( clk ) , .D( u0_uk_K_r6_0 ) , .Q( u0_uk_K_r7_0 ) );
  DFF_X1 u0_uk_K_r7_reg_1 (.CK( clk ) , .D( u0_uk_K_r6_1 ) , .Q( u0_uk_K_r7_1 ) , .QN( u0_uk_n317 ) );
  DFF_X1 u0_uk_K_r7_reg_10 (.CK( clk ) , .D( u0_uk_K_r6_10 ) , .Q( u0_uk_K_r7_10 ) , .QN( u0_uk_n311 ) );
  DFF_X1 u0_uk_K_r7_reg_11 (.CK( clk ) , .D( u0_uk_K_r6_11 ) , .Q( u0_uk_K_r7_11 ) , .QN( u0_uk_n310 ) );
  DFF_X1 u0_uk_K_r7_reg_12 (.CK( clk ) , .D( u0_uk_K_r6_12 ) , .Q( u0_uk_K_r7_12 ) , .QN( u0_uk_n309 ) );
  DFF_X1 u0_uk_K_r7_reg_13 (.CK( clk ) , .D( u0_uk_K_r6_13 ) , .Q( u0_uk_K_r7_13 ) );
  DFF_X1 u0_uk_K_r7_reg_14 (.CK( clk ) , .D( u0_uk_K_r6_14 ) , .Q( u0_uk_K_r7_14 ) , .QN( u0_uk_n307 ) );
  DFF_X1 u0_uk_K_r7_reg_15 (.CK( clk ) , .D( u0_uk_K_r6_15 ) , .Q( u0_uk_K_r7_15 ) );
  DFF_X1 u0_uk_K_r7_reg_16 (.CK( clk ) , .D( u0_uk_K_r6_16 ) , .Q( u0_uk_K_r7_16 ) );
  DFF_X1 u0_uk_K_r7_reg_17 (.CK( clk ) , .D( u0_uk_K_r6_17 ) , .Q( u0_uk_K_r7_17 ) , .QN( u0_uk_n304 ) );
  DFF_X1 u0_uk_K_r7_reg_18 (.CK( clk ) , .D( u0_uk_K_r6_18 ) , .Q( u0_uk_K_r7_18 ) , .QN( u0_uk_n303 ) );
  DFF_X1 u0_uk_K_r7_reg_19 (.CK( clk ) , .D( u0_uk_K_r6_19 ) , .Q( u0_uk_K_r7_19 ) , .QN( u0_uk_n302 ) );
  DFF_X1 u0_uk_K_r7_reg_2 (.CK( clk ) , .D( u0_uk_K_r6_2 ) , .Q( u0_uk_K_r7_2 ) , .QN( u0_uk_n316 ) );
  DFF_X1 u0_uk_K_r7_reg_20 (.CK( clk ) , .D( u0_uk_K_r6_20 ) , .Q( u0_uk_K_r7_20 ) );
  DFF_X1 u0_uk_K_r7_reg_21 (.CK( clk ) , .D( u0_uk_K_r6_21 ) , .Q( u0_uk_K_r7_21 ) , .QN( u0_uk_n300 ) );
  DFF_X1 u0_uk_K_r7_reg_22 (.CK( clk ) , .D( u0_uk_K_r6_22 ) , .Q( u0_uk_K_r7_22 ) );
  DFF_X1 u0_uk_K_r7_reg_23 (.CK( clk ) , .D( u0_uk_K_r6_23 ) , .Q( u0_uk_K_r7_23 ) );
  DFF_X1 u0_uk_K_r7_reg_24 (.CK( clk ) , .D( u0_uk_K_r6_24 ) , .Q( u0_uk_K_r7_24 ) , .QN( u0_uk_n296 ) );
  DFF_X1 u0_uk_K_r7_reg_25 (.CK( clk ) , .D( u0_uk_K_r6_25 ) , .Q( u0_uk_K_r7_25 ) , .QN( u0_uk_n295 ) );
  DFF_X1 u0_uk_K_r7_reg_26 (.CK( clk ) , .D( u0_uk_K_r6_26 ) , .Q( u0_uk_K_r7_26 ) );
  DFF_X1 u0_uk_K_r7_reg_27 (.CK( clk ) , .D( u0_uk_K_r6_27 ) , .Q( u0_uk_K_r7_27 ) );
  DFF_X1 u0_uk_K_r7_reg_28 (.CK( clk ) , .D( u0_uk_K_r6_28 ) , .Q( u0_uk_K_r7_28 ) , .QN( u0_uk_n293 ) );
  DFF_X1 u0_uk_K_r7_reg_29 (.CK( clk ) , .D( u0_uk_K_r6_29 ) , .Q( u0_uk_K_r7_29 ) );
  DFF_X1 u0_uk_K_r7_reg_3 (.CK( clk ) , .D( u0_uk_K_r6_3 ) , .Q( u0_uk_K_r7_3 ) , .QN( u0_uk_n315 ) );
  DFF_X1 u0_uk_K_r7_reg_30 (.CK( clk ) , .D( u0_uk_K_r6_30 ) , .Q( u0_uk_K_r7_30 ) );
  DFF_X1 u0_uk_K_r7_reg_31 (.CK( clk ) , .D( u0_uk_K_r6_31 ) , .Q( u0_uk_K_r7_31 ) );
  DFF_X1 u0_uk_K_r7_reg_32 (.CK( clk ) , .D( u0_uk_K_r6_32 ) , .Q( u0_uk_K_r7_32 ) );
  DFF_X1 u0_uk_K_r7_reg_33 (.CK( clk ) , .D( u0_uk_K_r6_33 ) , .Q( u0_uk_K_r7_33 ) , .QN( u0_uk_n290 ) );
  DFF_X1 u0_uk_K_r7_reg_34 (.CK( clk ) , .D( u0_uk_K_r6_34 ) , .Q( u0_uk_K_r7_34 ) );
  DFF_X1 u0_uk_K_r7_reg_35 (.CK( clk ) , .D( u0_uk_K_r6_35 ) , .Q( u0_uk_K_r7_35 ) , .QN( u0_uk_n289 ) );
  DFF_X1 u0_uk_K_r7_reg_36 (.CK( clk ) , .D( u0_uk_K_r6_36 ) , .Q( u0_uk_K_r7_36 ) , .QN( u0_uk_n288 ) );
  DFF_X1 u0_uk_K_r7_reg_37 (.CK( clk ) , .D( u0_uk_K_r6_37 ) , .Q( u0_uk_K_r7_37 ) );
  DFF_X1 u0_uk_K_r7_reg_38 (.CK( clk ) , .D( u0_uk_K_r6_38 ) , .Q( u0_uk_K_r7_38 ) , .QN( u0_uk_n287 ) );
  DFF_X1 u0_uk_K_r7_reg_39 (.CK( clk ) , .D( u0_uk_K_r6_39 ) , .Q( u0_uk_K_r7_39 ) );
  DFF_X1 u0_uk_K_r7_reg_4 (.CK( clk ) , .D( u0_uk_K_r6_4 ) , .Q( u0_uk_K_r7_4 ) , .QN( u0_uk_n314 ) );
  DFF_X1 u0_uk_K_r7_reg_40 (.CK( clk ) , .D( u0_uk_K_r6_40 ) , .Q( u0_uk_K_r7_40 ) , .QN( u0_uk_n285 ) );
  DFF_X1 u0_uk_K_r7_reg_41 (.CK( clk ) , .D( u0_uk_K_r6_41 ) , .Q( u0_uk_K_r7_41 ) , .QN( u0_uk_n284 ) );
  DFF_X1 u0_uk_K_r7_reg_42 (.CK( clk ) , .D( u0_uk_K_r6_42 ) , .Q( u0_uk_K_r7_42 ) , .QN( u0_uk_n283 ) );
  DFF_X1 u0_uk_K_r7_reg_43 (.CK( clk ) , .D( u0_uk_K_r6_43 ) , .Q( u0_uk_K_r7_43 ) , .QN( u0_uk_n282 ) );
  DFF_X1 u0_uk_K_r7_reg_44 (.CK( clk ) , .D( u0_uk_K_r6_44 ) , .Q( u0_uk_K_r7_44 ) , .QN( u0_uk_n281 ) );
  DFF_X1 u0_uk_K_r7_reg_45 (.CK( clk ) , .D( u0_uk_K_r6_45 ) , .Q( u0_uk_K_r7_45 ) , .QN( u0_uk_n280 ) );
  DFF_X1 u0_uk_K_r7_reg_46 (.CK( clk ) , .D( u0_uk_K_r6_46 ) , .Q( u0_uk_K_r7_46 ) );
  DFF_X1 u0_uk_K_r7_reg_47 (.CK( clk ) , .D( u0_uk_K_r6_47 ) , .Q( u0_uk_K_r7_47 ) , .QN( u0_uk_n278 ) );
  DFF_X1 u0_uk_K_r7_reg_48 (.CK( clk ) , .D( u0_uk_K_r6_48 ) , .Q( u0_uk_K_r7_48 ) );
  DFF_X1 u0_uk_K_r7_reg_49 (.CK( clk ) , .D( u0_uk_K_r6_49 ) , .Q( u0_uk_K_r7_49 ) , .QN( u0_uk_n276 ) );
  DFF_X1 u0_uk_K_r7_reg_5 (.CK( clk ) , .D( u0_uk_K_r6_5 ) , .Q( u0_uk_K_r7_5 ) );
  DFF_X1 u0_uk_K_r7_reg_50 (.CK( clk ) , .D( u0_uk_K_r6_50 ) , .Q( u0_uk_K_r7_50 ) , .QN( u0_uk_n275 ) );
  DFF_X1 u0_uk_K_r7_reg_51 (.CK( clk ) , .D( u0_uk_K_r6_51 ) , .Q( u0_uk_K_r7_51 ) , .QN( u0_uk_n274 ) );
  DFF_X1 u0_uk_K_r7_reg_52 (.CK( clk ) , .D( u0_uk_K_r6_52 ) , .Q( u0_uk_K_r7_52 ) , .QN( u0_uk_n273 ) );
  DFF_X1 u0_uk_K_r7_reg_53 (.CK( clk ) , .D( u0_uk_K_r6_53 ) , .Q( u0_uk_K_r7_53 ) );
  DFF_X1 u0_uk_K_r7_reg_54 (.CK( clk ) , .D( u0_uk_K_r6_54 ) , .Q( u0_uk_K_r7_54 ) , .QN( u0_uk_n272 ) );
  DFF_X1 u0_uk_K_r7_reg_55 (.CK( clk ) , .D( u0_uk_K_r6_55 ) , .Q( u0_uk_K_r7_55 ) );
  DFF_X1 u0_uk_K_r7_reg_6 (.CK( clk ) , .D( u0_uk_K_r6_6 ) , .Q( u0_uk_K_r7_6 ) );
  DFF_X1 u0_uk_K_r7_reg_7 (.CK( clk ) , .D( u0_uk_K_r6_7 ) , .Q( u0_uk_K_r7_7 ) );
  DFF_X1 u0_uk_K_r7_reg_8 (.CK( clk ) , .D( u0_uk_K_r6_8 ) , .Q( u0_uk_K_r7_8 ) );
  DFF_X1 u0_uk_K_r7_reg_9 (.CK( clk ) , .D( u0_uk_K_r6_9 ) , .Q( u0_uk_K_r7_9 ) );
  DFF_X1 u0_uk_K_r8_reg_0 (.CK( clk ) , .D( u0_uk_K_r7_0 ) , .Q( u0_uk_K_r8_0 ) , .QN( u0_uk_n270 ) );
  DFF_X1 u0_uk_K_r8_reg_1 (.CK( clk ) , .D( u0_uk_K_r7_1 ) , .Q( u0_uk_K_r8_1 ) , .QN( u0_uk_n269 ) );
  DFF_X1 u0_uk_K_r8_reg_10 (.CK( clk ) , .D( u0_uk_K_r7_10 ) , .Q( u0_uk_K_r8_10 ) );
  DFF_X1 u0_uk_K_r8_reg_11 (.CK( clk ) , .D( u0_uk_K_r7_11 ) , .Q( u0_uk_K_r8_11 ) , .QN( u0_uk_n263 ) );
  DFF_X1 u0_uk_K_r8_reg_12 (.CK( clk ) , .D( u0_uk_K_r7_12 ) , .Q( u0_uk_K_r8_12 ) , .QN( u0_uk_n262 ) );
  DFF_X1 u0_uk_K_r8_reg_13 (.CK( clk ) , .D( u0_uk_K_r7_13 ) , .Q( u0_uk_K_r8_13 ) );
  DFF_X1 u0_uk_K_r8_reg_14 (.CK( clk ) , .D( u0_uk_K_r7_14 ) , .Q( u0_uk_K_r8_14 ) , .QN( u0_uk_n261 ) );
  DFF_X1 u0_uk_K_r8_reg_15 (.CK( clk ) , .D( u0_uk_K_r7_15 ) , .Q( u0_uk_K_r8_15 ) , .QN( u0_uk_n260 ) );
  DFF_X1 u0_uk_K_r8_reg_16 (.CK( clk ) , .D( u0_uk_K_r7_16 ) , .Q( u0_uk_K_r8_16 ) );
  DFF_X1 u0_uk_K_r8_reg_17 (.CK( clk ) , .D( u0_uk_K_r7_17 ) , .Q( u0_uk_K_r8_17 ) );
  DFF_X1 u0_uk_K_r8_reg_18 (.CK( clk ) , .D( u0_uk_K_r7_18 ) , .Q( u0_uk_K_r8_18 ) , .QN( u0_uk_n259 ) );
  DFF_X1 u0_uk_K_r8_reg_19 (.CK( clk ) , .D( u0_uk_K_r7_19 ) , .Q( u0_uk_K_r8_19 ) );
  DFF_X1 u0_uk_K_r8_reg_2 (.CK( clk ) , .D( u0_uk_K_r7_2 ) , .Q( u0_uk_K_r8_2 ) );
  DFF_X1 u0_uk_K_r8_reg_20 (.CK( clk ) , .D( u0_uk_K_r7_20 ) , .Q( u0_uk_K_r8_20 ) , .QN( u0_uk_n258 ) );
  DFF_X1 u0_uk_K_r8_reg_21 (.CK( clk ) , .D( u0_uk_K_r7_21 ) , .Q( u0_uk_K_r8_21 ) );
  DFF_X1 u0_uk_K_r8_reg_22 (.CK( clk ) , .D( u0_uk_K_r7_22 ) , .Q( u0_uk_K_r8_22 ) );
  DFF_X1 u0_uk_K_r8_reg_23 (.CK( clk ) , .D( u0_uk_K_r7_23 ) , .Q( u0_uk_K_r8_23 ) , .QN( u0_uk_n256 ) );
  DFF_X1 u0_uk_K_r8_reg_24 (.CK( clk ) , .D( u0_uk_K_r7_24 ) , .Q( u0_uk_K_r8_24 ) , .QN( u0_uk_n255 ) );
  DFF_X1 u0_uk_K_r8_reg_25 (.CK( clk ) , .D( u0_uk_K_r7_25 ) , .Q( u0_uk_K_r8_25 ) , .QN( u0_uk_n254 ) );
  DFF_X1 u0_uk_K_r8_reg_26 (.CK( clk ) , .D( u0_uk_K_r7_26 ) , .Q( u0_uk_K_r8_26 ) , .QN( u0_uk_n253 ) );
  DFF_X1 u0_uk_K_r8_reg_27 (.CK( clk ) , .D( u0_uk_K_r7_27 ) , .Q( u0_uk_K_r8_27 ) );
  DFF_X1 u0_uk_K_r8_reg_28 (.CK( clk ) , .D( u0_uk_K_r7_28 ) , .Q( u0_uk_K_r8_28 ) );
  DFF_X1 u0_uk_K_r8_reg_29 (.CK( clk ) , .D( u0_uk_K_r7_29 ) , .Q( u0_uk_K_r8_29 ) , .QN( u0_uk_n249 ) );
  DFF_X1 u0_uk_K_r8_reg_3 (.CK( clk ) , .D( u0_uk_K_r7_3 ) , .Q( u0_uk_K_r8_3 ) , .QN( u0_uk_n268 ) );
  DFF_X1 u0_uk_K_r8_reg_30 (.CK( clk ) , .D( u0_uk_K_r7_30 ) , .Q( u0_uk_K_r8_30 ) , .QN( u0_uk_n248 ) );
  DFF_X1 u0_uk_K_r8_reg_31 (.CK( clk ) , .D( u0_uk_K_r7_31 ) , .Q( u0_uk_K_r8_31 ) , .QN( u0_uk_n247 ) );
  DFF_X1 u0_uk_K_r8_reg_32 (.CK( clk ) , .D( u0_uk_K_r7_32 ) , .Q( u0_uk_K_r8_32 ) );
  DFF_X1 u0_uk_K_r8_reg_33 (.CK( clk ) , .D( u0_uk_K_r7_33 ) , .Q( u0_uk_K_r8_33 ) , .QN( u0_uk_n246 ) );
  DFF_X1 u0_uk_K_r8_reg_34 (.CK( clk ) , .D( u0_uk_K_r7_34 ) , .Q( u0_uk_K_r8_34 ) , .QN( u0_uk_n245 ) );
  DFF_X1 u0_uk_K_r8_reg_35 (.CK( clk ) , .D( u0_uk_K_r7_35 ) , .Q( u0_uk_K_r8_35 ) , .QN( u0_uk_n244 ) );
  DFF_X1 u0_uk_K_r8_reg_36 (.CK( clk ) , .D( u0_uk_K_r7_36 ) , .Q( u0_uk_K_r8_36 ) , .QN( u0_uk_n243 ) );
  DFF_X1 u0_uk_K_r8_reg_37 (.CK( clk ) , .D( u0_uk_K_r7_37 ) , .Q( u0_uk_K_r8_37 ) );
  DFF_X1 u0_uk_K_r8_reg_38 (.CK( clk ) , .D( u0_uk_K_r7_38 ) , .Q( u0_uk_K_r8_38 ) , .QN( u0_uk_n241 ) );
  DFF_X1 u0_uk_K_r8_reg_39 (.CK( clk ) , .D( u0_uk_K_r7_39 ) , .Q( u0_uk_K_r8_39 ) , .QN( u0_uk_n239 ) );
  DFF_X1 u0_uk_K_r8_reg_4 (.CK( clk ) , .D( u0_uk_K_r7_4 ) , .Q( u0_uk_K_r8_4 ) , .QN( u0_uk_n267 ) );
  DFF_X1 u0_uk_K_r8_reg_40 (.CK( clk ) , .D( u0_uk_K_r7_40 ) , .Q( u0_uk_K_r8_40 ) );
  DFF_X1 u0_uk_K_r8_reg_41 (.CK( clk ) , .D( u0_uk_K_r7_41 ) , .Q( u0_uk_K_r8_41 ) );
  DFF_X1 u0_uk_K_r8_reg_42 (.CK( clk ) , .D( u0_uk_K_r7_42 ) , .Q( u0_uk_K_r8_42 ) , .QN( u0_uk_n237 ) );
  DFF_X1 u0_uk_K_r8_reg_43 (.CK( clk ) , .D( u0_uk_K_r7_43 ) , .Q( u0_uk_K_r8_43 ) );
  DFF_X1 u0_uk_K_r8_reg_44 (.CK( clk ) , .D( u0_uk_K_r7_44 ) , .Q( u0_uk_K_r8_44 ) , .QN( u0_uk_n236 ) );
  DFF_X1 u0_uk_K_r8_reg_45 (.CK( clk ) , .D( u0_uk_K_r7_45 ) , .Q( u0_uk_K_r8_45 ) );
  DFF_X1 u0_uk_K_r8_reg_46 (.CK( clk ) , .D( u0_uk_K_r7_46 ) , .Q( u0_uk_K_r8_46 ) , .QN( u0_uk_n235 ) );
  DFF_X1 u0_uk_K_r8_reg_47 (.CK( clk ) , .D( u0_uk_K_r7_47 ) , .Q( u0_uk_K_r8_47 ) , .QN( u0_uk_n234 ) );
  DFF_X1 u0_uk_K_r8_reg_48 (.CK( clk ) , .D( u0_uk_K_r7_48 ) , .Q( u0_uk_K_r8_48 ) );
  DFF_X1 u0_uk_K_r8_reg_49 (.CK( clk ) , .D( u0_uk_K_r7_49 ) , .Q( u0_uk_K_r8_49 ) , .QN( u0_uk_n233 ) );
  DFF_X1 u0_uk_K_r8_reg_5 (.CK( clk ) , .D( u0_uk_K_r7_5 ) , .Q( u0_uk_K_r8_5 ) );
  DFF_X1 u0_uk_K_r8_reg_50 (.CK( clk ) , .D( u0_uk_K_r7_50 ) , .Q( u0_uk_K_r8_50 ) , .QN( u0_uk_n232 ) );
  DFF_X1 u0_uk_K_r8_reg_51 (.CK( clk ) , .D( u0_uk_K_r7_51 ) , .Q( u0_uk_K_r8_51 ) );
  DFF_X1 u0_uk_K_r8_reg_52 (.CK( clk ) , .D( u0_uk_K_r7_52 ) , .Q( u0_uk_K_r8_52 ) );
  DFF_X1 u0_uk_K_r8_reg_53 (.CK( clk ) , .D( u0_uk_K_r7_53 ) , .Q( u0_uk_K_r8_53 ) , .QN( u0_uk_n229 ) );
  DFF_X1 u0_uk_K_r8_reg_54 (.CK( clk ) , .D( u0_uk_K_r7_54 ) , .Q( u0_uk_K_r8_54 ) , .QN( u0_uk_n228 ) );
  DFF_X1 u0_uk_K_r8_reg_55 (.CK( clk ) , .D( u0_uk_K_r7_55 ) , .Q( u0_uk_K_r8_55 ) , .QN( u0_uk_n227 ) );
  DFF_X1 u0_uk_K_r8_reg_6 (.CK( clk ) , .D( u0_uk_K_r7_6 ) , .Q( u0_uk_K_r8_6 ) , .QN( u0_uk_n266 ) );
  DFF_X1 u0_uk_K_r8_reg_7 (.CK( clk ) , .D( u0_uk_K_r7_7 ) , .Q( u0_uk_K_r8_7 ) , .QN( u0_uk_n265 ) );
  DFF_X1 u0_uk_K_r8_reg_8 (.CK( clk ) , .D( u0_uk_K_r7_8 ) , .Q( u0_uk_K_r8_8 ) );
  DFF_X1 u0_uk_K_r8_reg_9 (.CK( clk ) , .D( u0_uk_K_r7_9 ) , .Q( u0_uk_K_r8_9 ) , .QN( u0_uk_n264 ) );
  DFF_X1 u0_uk_K_r9_reg_0 (.CK( clk ) , .D( u0_uk_K_r8_0 ) , .Q( u0_uk_K_r9_0 ) );
  DFF_X1 u0_uk_K_r9_reg_1 (.CK( clk ) , .D( u0_uk_K_r8_1 ) , .Q( u0_uk_K_r9_1 ) , .QN( u0_uk_n226 ) );
  DFF_X1 u0_uk_K_r9_reg_10 (.CK( clk ) , .D( u0_uk_K_r8_10 ) , .Q( u0_uk_K_r9_10 ) );
  DFF_X1 u0_uk_K_r9_reg_11 (.CK( clk ) , .D( u0_uk_K_r8_11 ) , .Q( u0_uk_K_r9_11 ) , .QN( u0_uk_n221 ) );
  DFF_X1 u0_uk_K_r9_reg_12 (.CK( clk ) , .D( u0_uk_K_r8_12 ) , .Q( u0_uk_K_r9_12 ) );
  DFF_X1 u0_uk_K_r9_reg_13 (.CK( clk ) , .D( u0_uk_K_r8_13 ) , .Q( u0_uk_K_r9_13 ) , .QN( u0_uk_n219 ) );
  DFF_X1 u0_uk_K_r9_reg_14 (.CK( clk ) , .D( u0_uk_K_r8_14 ) , .Q( u0_uk_K_r9_14 ) , .QN( u0_uk_n218 ) );
  DFF_X1 u0_uk_K_r9_reg_15 (.CK( clk ) , .D( u0_uk_K_r8_15 ) , .Q( u0_uk_K_r9_15 ) );
  DFF_X1 u0_uk_K_r9_reg_16 (.CK( clk ) , .D( u0_uk_K_r8_16 ) , .Q( u0_uk_K_r9_16 ) , .QN( u0_uk_n216 ) );
  DFF_X1 u0_uk_K_r9_reg_17 (.CK( clk ) , .D( u0_uk_K_r8_17 ) , .Q( u0_uk_K_r9_17 ) , .QN( u0_uk_n215 ) );
  DFF_X1 u0_uk_K_r9_reg_18 (.CK( clk ) , .D( u0_uk_K_r8_18 ) , .Q( u0_uk_K_r9_18 ) );
  DFF_X1 u0_uk_K_r9_reg_19 (.CK( clk ) , .D( u0_uk_K_r8_19 ) , .Q( u0_uk_K_r9_19 ) );
  DFF_X1 u0_uk_K_r9_reg_2 (.CK( clk ) , .D( u0_uk_K_r8_2 ) , .Q( u0_uk_K_r9_2 ) );
  DFF_X1 u0_uk_K_r9_reg_20 (.CK( clk ) , .D( u0_uk_K_r8_20 ) , .Q( u0_uk_K_r9_20 ) , .QN( u0_uk_n212 ) );
  DFF_X1 u0_uk_K_r9_reg_21 (.CK( clk ) , .D( u0_uk_K_r8_21 ) , .Q( u0_uk_K_r9_21 ) , .QN( u0_uk_n211 ) );
  DFF_X1 u0_uk_K_r9_reg_22 (.CK( clk ) , .D( u0_uk_K_r8_22 ) , .Q( u0_uk_K_r9_22 ) , .QN( u0_uk_n210 ) );
  DFF_X1 u0_uk_K_r9_reg_23 (.CK( clk ) , .D( u0_uk_K_r8_23 ) , .Q( u0_uk_K_r9_23 ) );
  DFF_X1 u0_uk_K_r9_reg_24 (.CK( clk ) , .D( u0_uk_K_r8_24 ) , .Q( u0_uk_K_r9_24 ) );
  DFF_X1 u0_uk_K_r9_reg_25 (.CK( clk ) , .D( u0_uk_K_r8_25 ) , .Q( u0_uk_K_r9_25 ) );
  DFF_X1 u0_uk_K_r9_reg_26 (.CK( clk ) , .D( u0_uk_K_r8_26 ) , .Q( u0_uk_K_r9_26 ) , .QN( u0_uk_n206 ) );
  DFF_X1 u0_uk_K_r9_reg_27 (.CK( clk ) , .D( u0_uk_K_r8_27 ) , .Q( u0_uk_K_r9_27 ) );
  DFF_X1 u0_uk_K_r9_reg_28 (.CK( clk ) , .D( u0_uk_K_r8_28 ) , .Q( u0_uk_K_r9_28 ) , .QN( u0_uk_n205 ) );
  DFF_X1 u0_uk_K_r9_reg_29 (.CK( clk ) , .D( u0_uk_K_r8_29 ) , .Q( u0_uk_K_r9_29 ) , .QN( u0_uk_n204 ) );
  DFF_X1 u0_uk_K_r9_reg_3 (.CK( clk ) , .D( u0_uk_K_r8_3 ) , .Q( u0_uk_K_r9_3 ) , .QN( u0_uk_n225 ) );
  DFF_X1 u0_uk_K_r9_reg_30 (.CK( clk ) , .D( u0_uk_K_r8_30 ) , .Q( u0_uk_K_r9_30 ) );
  DFF_X1 u0_uk_K_r9_reg_31 (.CK( clk ) , .D( u0_uk_K_r8_31 ) , .Q( u0_uk_K_r9_31 ) );
  DFF_X1 u0_uk_K_r9_reg_32 (.CK( clk ) , .D( u0_uk_K_r8_32 ) , .Q( u0_uk_K_r9_32 ) , .QN( u0_uk_n201 ) );
  DFF_X1 u0_uk_K_r9_reg_33 (.CK( clk ) , .D( u0_uk_K_r8_33 ) , .Q( u0_uk_K_r9_33 ) );
  DFF_X1 u0_uk_K_r9_reg_34 (.CK( clk ) , .D( u0_uk_K_r8_34 ) , .Q( u0_uk_K_r9_34 ) , .QN( u0_uk_n200 ) );
  DFF_X1 u0_uk_K_r9_reg_35 (.CK( clk ) , .D( u0_uk_K_r8_35 ) , .Q( u0_uk_K_r9_35 ) );
  DFF_X1 u0_uk_K_r9_reg_36 (.CK( clk ) , .D( u0_uk_K_r8_36 ) , .Q( u0_uk_K_r9_36 ) , .QN( u0_uk_n199 ) );
  DFF_X1 u0_uk_K_r9_reg_37 (.CK( clk ) , .D( u0_uk_K_r8_37 ) , .Q( u0_uk_K_r9_37 ) , .QN( u0_uk_n198 ) );
  DFF_X1 u0_uk_K_r9_reg_38 (.CK( clk ) , .D( u0_uk_K_r8_38 ) , .Q( u0_uk_K_r9_38 ) );
  DFF_X1 u0_uk_K_r9_reg_39 (.CK( clk ) , .D( u0_uk_K_r8_39 ) , .Q( u0_uk_K_r9_39 ) , .QN( u0_uk_n197 ) );
  DFF_X1 u0_uk_K_r9_reg_4 (.CK( clk ) , .D( u0_uk_K_r8_4 ) , .Q( u0_uk_K_r9_4 ) );
  DFF_X1 u0_uk_K_r9_reg_40 (.CK( clk ) , .D( u0_uk_K_r8_40 ) , .Q( u0_uk_K_r9_40 ) , .QN( u0_uk_n196 ) );
  DFF_X1 u0_uk_K_r9_reg_41 (.CK( clk ) , .D( u0_uk_K_r8_41 ) , .Q( u0_uk_K_r9_41 ) , .QN( u0_uk_n195 ) );
  DFF_X1 u0_uk_K_r9_reg_42 (.CK( clk ) , .D( u0_uk_K_r8_42 ) , .Q( u0_uk_K_r9_42 ) , .QN( u0_uk_n194 ) );
  DFF_X1 u0_uk_K_r9_reg_43 (.CK( clk ) , .D( u0_uk_K_r8_43 ) , .Q( u0_uk_K_r9_43 ) , .QN( u0_uk_n193 ) );
  DFF_X1 u0_uk_K_r9_reg_44 (.CK( clk ) , .D( u0_uk_K_r8_44 ) , .Q( u0_uk_K_r9_44 ) , .QN( u0_uk_n192 ) );
  DFF_X1 u0_uk_K_r9_reg_45 (.CK( clk ) , .D( u0_uk_K_r8_45 ) , .Q( u0_uk_K_r9_45 ) );
  DFF_X1 u0_uk_K_r9_reg_46 (.CK( clk ) , .D( u0_uk_K_r8_46 ) , .Q( u0_uk_K_r9_46 ) , .QN( u0_uk_n190 ) );
  DFF_X1 u0_uk_K_r9_reg_47 (.CK( clk ) , .D( u0_uk_K_r8_47 ) , .Q( u0_uk_K_r9_47 ) , .QN( u0_uk_n189 ) );
  DFF_X1 u0_uk_K_r9_reg_48 (.CK( clk ) , .D( u0_uk_K_r8_48 ) , .Q( u0_uk_K_r9_48 ) );
  DFF_X1 u0_uk_K_r9_reg_49 (.CK( clk ) , .D( u0_uk_K_r8_49 ) , .Q( u0_uk_K_r9_49 ) );
  DFF_X1 u0_uk_K_r9_reg_5 (.CK( clk ) , .D( u0_uk_K_r8_5 ) , .Q( u0_uk_K_r9_5 ) );
  DFF_X1 u0_uk_K_r9_reg_50 (.CK( clk ) , .D( u0_uk_K_r8_50 ) , .Q( u0_uk_K_r9_50 ) , .QN( u0_uk_n186 ) );
  DFF_X1 u0_uk_K_r9_reg_51 (.CK( clk ) , .D( u0_uk_K_r8_51 ) , .Q( u0_uk_K_r9_51 ) , .QN( u0_uk_n185 ) );
  DFF_X1 u0_uk_K_r9_reg_52 (.CK( clk ) , .D( u0_uk_K_r8_52 ) , .Q( u0_uk_K_r9_52 ) , .QN( u0_uk_n184 ) );
  DFF_X1 u0_uk_K_r9_reg_53 (.CK( clk ) , .D( u0_uk_K_r8_53 ) , .Q( u0_uk_K_r9_53 ) , .QN( u0_uk_n183 ) );
  DFF_X1 u0_uk_K_r9_reg_54 (.CK( clk ) , .D( u0_uk_K_r8_54 ) , .Q( u0_uk_K_r9_54 ) );
  DFF_X1 u0_uk_K_r9_reg_55 (.CK( clk ) , .D( u0_uk_K_r8_55 ) , .Q( u0_uk_K_r9_55 ) , .QN( u0_uk_n181 ) );
  DFF_X1 u0_uk_K_r9_reg_6 (.CK( clk ) , .D( u0_uk_K_r8_6 ) , .Q( u0_uk_K_r9_6 ) );
  DFF_X1 u0_uk_K_r9_reg_7 (.CK( clk ) , .D( u0_uk_K_r8_7 ) , .Q( u0_uk_K_r9_7 ) );
  DFF_X1 u0_uk_K_r9_reg_8 (.CK( clk ) , .D( u0_uk_K_r8_8 ) , .Q( u0_uk_K_r9_8 ) , .QN( u0_uk_n224 ) );
  DFF_X1 u0_uk_K_r9_reg_9 (.CK( clk ) , .D( u0_uk_K_r8_9 ) , .Q( u0_uk_K_r9_9 ) );
  OAI21_X1 u0_uk_U1000 (.B1( decrypt ) , .ZN( u0_K14_46 ) , .B2( u0_uk_n68 ) , .A( u0_uk_n928 ) );
  NAND2_X1 u0_uk_U1001 (.A2( decrypt ) , .A1( u0_uk_K_r12_22 ) , .ZN( u0_uk_n928 ) );
  OAI21_X1 u0_uk_U1004 (.B1( decrypt ) , .ZN( u0_K3_5 ) , .B2( u0_uk_n556 ) , .A( u0_uk_n841 ) );
  OAI21_X1 u0_uk_U1008 (.B1( decrypt ) , .ZN( u0_K1_13 ) , .B2( u0_uk_n674 ) , .A( u0_uk_n890 ) );
  OAI21_X1 u0_uk_U1010 (.B1( decrypt ) , .ZN( u0_K1_17 ) , .B2( u0_uk_n705 ) , .A( u0_uk_n888 ) );
  NAND2_X1 u0_uk_U1013 (.A2( decrypt ) , .A1( u0_uk_K_r8_19 ) , .ZN( u0_uk_n1020 ) );
  OAI21_X1 u0_uk_U1016 (.B1( decrypt ) , .ZN( u0_K9_39 ) , .B2( u0_uk_n287 ) , .A( u0_uk_n724 ) );
  NAND2_X1 u0_uk_U1017 (.A2( decrypt ) , .A1( u0_uk_K_r7_31 ) , .ZN( u0_uk_n724 ) );
  OAI21_X1 u0_uk_U1018 (.B1( decrypt ) , .ZN( u0_K4_6 ) , .B2( u0_uk_n523 ) , .A( u0_uk_n820 ) );
  NAND2_X1 u0_uk_U1019 (.A2( decrypt ) , .A1( u0_uk_K_r2_24 ) , .ZN( u0_uk_n820 ) );
  OAI21_X1 u0_uk_U1026 (.B1( decrypt ) , .ZN( u0_K10_13 ) , .A( u0_uk_n1023 ) , .B2( u0_uk_n253 ) );
  NAND2_X1 u0_uk_U1027 (.A2( decrypt ) , .A1( u0_uk_K_r8_48 ) , .ZN( u0_uk_n1023 ) );
  OAI21_X1 u0_uk_U1028 (.B1( decrypt ) , .ZN( u0_K12_36 ) , .B2( u0_uk_n160 ) , .A( u0_uk_n970 ) );
  NAND2_X1 u0_uk_U1029 (.A2( decrypt ) , .A1( u0_uk_K_r10_52 ) , .ZN( u0_uk_n970 ) );
  NAND2_X1 u0_uk_U1031 (.A2( decrypt ) , .A1( u0_uk_K_r14_42 ) , .ZN( u0_uk_n898 ) );
  NAND2_X1 u0_uk_U1033 (.A2( decrypt ) , .A1( u0_uk_K_r6_30 ) , .ZN( u0_uk_n748 ) );
  OAI21_X1 u0_uk_U1034 (.B1( decrypt ) , .ZN( u0_K6_41 ) , .B2( u0_uk_n413 ) , .A( u0_uk_n790 ) );
  OAI21_X1 u0_uk_U1038 (.B1( decrypt ) , .ZN( u0_K8_28 ) , .B2( u0_uk_n326 ) , .A( u0_uk_n756 ) );
  OAI21_X1 u0_uk_U1046 (.B1( decrypt ) , .ZN( u0_K10_32 ) , .A( u0_uk_n1013 ) , .B2( u0_uk_n270 ) );
  NAND2_X1 u0_uk_U1047 (.A2( decrypt ) , .A1( u0_uk_K_r8_51 ) , .ZN( u0_uk_n1013 ) );
  OAI21_X1 u0_uk_U1048 (.B1( decrypt ) , .ZN( u0_K5_31 ) , .B2( u0_uk_n487 ) , .A( u0_uk_n812 ) );
  NAND2_X1 u0_uk_U1049 (.A2( decrypt ) , .A1( u0_uk_K_r3_44 ) , .ZN( u0_uk_n812 ) );
  NAND2_X1 u0_uk_U1051 (.A2( decrypt ) , .A1( u0_uk_K_r13_36 ) , .ZN( u0_uk_n918 ) );
  NAND2_X1 u0_uk_U1053 (.A2( decrypt ) , .A1( u0_uk_K_r14_38 ) , .ZN( u0_uk_n897 ) );
  OAI22_X1 u0_uk_U106 (.B1( decrypt ) , .ZN( u0_K2_5 ) , .A1( u0_uk_n209 ) , .A2( u0_uk_n611 ) , .B2( u0_uk_n614 ) );
  OAI21_X1 u0_uk_U1060 (.B1( decrypt ) , .ZN( u0_K14_24 ) , .B2( u0_uk_n76 ) , .A( u0_uk_n937 ) );
  NAND2_X1 u0_uk_U1061 (.A2( decrypt ) , .A1( u0_uk_K_r12_41 ) , .ZN( u0_uk_n937 ) );
  OAI22_X1 u0_uk_U108 (.B1( decrypt ) , .ZN( u0_K10_41 ) , .A1( u0_uk_n163 ) , .B2( u0_uk_n236 ) , .A2( u0_uk_n264 ) );
  AOI22_X1 u0_uk_U1118 (.B1( decrypt ) , .B2( u0_uk_K_r10_27 ) , .A2( u0_uk_K_r10_4 ) , .A1( u0_uk_n238 ) , .ZN( u0_uk_n963 ) );
  AOI22_X1 u0_uk_U1120 (.B1( decrypt ) , .B2( u0_uk_K_r0_13 ) , .A2( u0_uk_K_r0_34 ) , .A1( u0_uk_n222 ) , .ZN( u0_uk_n855 ) );
  AOI22_X1 u0_uk_U1140 (.A1( decrypt ) , .B2( u0_uk_K_r5_0 ) , .A2( u0_uk_K_r5_35 ) , .B1( u0_uk_n207 ) , .ZN( u0_uk_n770 ) );
  AOI22_X1 u0_uk_U1142 (.A1( decrypt ) , .B2( u0_uk_K_r8_17 ) , .A2( u0_uk_K_r8_39 ) , .ZN( u0_uk_n1024 ) , .B1( u0_uk_n203 ) );
  AOI22_X1 u0_uk_U1146 (.A1( decrypt ) , .B2( u0_uk_K_r6_10 ) , .A2( u0_uk_K_r6_17 ) , .B1( u0_uk_n163 ) , .ZN( u0_uk_n759 ) );
  AOI22_X1 u0_uk_U1148 (.A1( decrypt ) , .B2( u0_uk_K_r3_29 ) , .A2( u0_uk_K_r3_38 ) , .B1( u0_uk_n202 ) , .ZN( u0_uk_n810 ) );
  AOI22_X1 u0_uk_U1155 (.A1( decrypt ) , .B2( u0_uk_K_r4_17 ) , .A2( u0_uk_K_r4_55 ) , .B1( u0_uk_n207 ) , .ZN( u0_uk_n793 ) );
  OAI22_X1 u0_uk_U122 (.B1( decrypt ) , .ZN( u0_K5_47 ) , .A1( u0_uk_n238 ) , .A2( u0_uk_n469 ) , .B2( u0_uk_n493 ) );
  OAI21_X1 u0_uk_U124 (.B1( decrypt ) , .ZN( u0_K2_47 ) , .B2( u0_uk_n617 ) , .A( u0_uk_n856 ) );
  OAI22_X1 u0_uk_U126 (.A1( decrypt ) , .ZN( u0_K1_15 ) , .B1( u0_uk_n252 ) , .A2( u0_uk_n691 ) , .B2( u0_uk_n697 ) );
  OAI21_X1 u0_uk_U128 (.B1( decrypt ) , .ZN( u0_K5_15 ) , .B2( u0_uk_n479 ) , .A( u0_uk_n817 ) );
  NAND2_X1 u0_uk_U129 (.A2( decrypt ) , .A1( u0_uk_K_r3_34 ) , .ZN( u0_uk_n817 ) );
  OAI22_X1 u0_uk_U135 (.B1( decrypt ) , .ZN( u0_K3_15 ) , .A1( u0_uk_n191 ) , .B2( u0_uk_n541 ) , .A2( u0_uk_n576 ) );
  OAI22_X1 u0_uk_U138 (.A1( decrypt ) , .ZN( u0_K12_19 ) , .B2( u0_uk_n138 ) , .A2( u0_uk_n176 ) , .B1( u0_uk_n217 ) );
  OAI21_X1 u0_uk_U140 (.B1( decrypt ) , .ZN( u0_K6_19 ) , .B2( u0_uk_n444 ) , .A( u0_uk_n798 ) );
  AOI22_X1 u0_uk_U154 (.B2( decrypt ) , .B1( u0_uk_K_r7_13 ) , .A2( u0_uk_K_r7_20 ) , .A1( u0_uk_n238 ) , .ZN( u0_uk_n735 ) );
  OAI21_X1 u0_uk_U157 (.B1( decrypt ) , .ZN( u0_K3_19 ) , .B2( u0_uk_n564 ) , .A( u0_uk_n852 ) );
  NAND2_X1 u0_uk_U158 (.A2( decrypt ) , .A1( u0_uk_K_r1_33 ) , .ZN( u0_uk_n852 ) );
  OAI22_X1 u0_uk_U161 (.A1( decrypt ) , .ZN( u0_K14_15 ) , .B1( u0_uk_n148 ) , .B2( u0_uk_n47 ) , .A2( u0_uk_n85 ) );
  OAI22_X1 u0_uk_U162 (.B1( decrypt ) , .ZN( u0_K8_19 ) , .A1( u0_uk_n223 ) , .A2( u0_uk_n343 ) , .B2( u0_uk_n350 ) );
  OAI22_X1 u0_uk_U163 (.A1( decrypt ) , .ZN( u0_K10_19 ) , .B1( u0_uk_n188 ) , .A2( u0_uk_n245 ) , .B2( u0_uk_n255 ) );
  OAI22_X1 u0_uk_U165 (.B1( decrypt ) , .ZN( u0_K2_30 ) , .A1( u0_uk_n188 ) , .A2( u0_uk_n599 ) , .B2( u0_uk_n628 ) );
  OAI21_X1 u0_uk_U170 (.B1( decrypt ) , .ZN( u0_K1_14 ) , .B2( u0_uk_n698 ) , .A( u0_uk_n889 ) );
  AOI22_X1 u0_uk_U181 (.A1( decrypt ) , .B2( u0_uk_K_r9_12 ) , .A2( u0_uk_K_r9_6 ) , .ZN( u0_uk_n1002 ) , .B1( u0_uk_n163 ) );
  OAI21_X1 u0_uk_U184 (.B1( decrypt ) , .ZN( u0_K9_14 ) , .B2( u0_uk_n284 ) , .A( u0_uk_n738 ) );
  NAND2_X1 u0_uk_U185 (.A2( decrypt ) , .A1( u0_uk_K_r7_34 ) , .ZN( u0_uk_n738 ) );
  OAI22_X1 u0_uk_U192 (.A1( decrypt ) , .ZN( u0_K10_14 ) , .B1( u0_uk_n182 ) , .A2( u0_uk_n227 ) , .B2( u0_uk_n258 ) );
  OAI21_X1 u0_uk_U193 (.B1( decrypt ) , .ZN( u0_K13_30 ) , .B2( u0_uk_n112 ) , .A( u0_uk_n945 ) );
  OAI22_X1 u0_uk_U197 (.A1( decrypt ) , .ZN( u0_K4_24 ) , .B1( u0_uk_n148 ) , .A2( u0_uk_n495 ) , .B2( u0_uk_n536 ) );
  OAI21_X1 u0_uk_U201 (.B1( decrypt ) , .ZN( u0_K1_30 ) , .B2( u0_uk_n675 ) , .A( u0_uk_n880 ) );
  NAND2_X1 u0_uk_U204 (.A2( decrypt ) , .A1( u0_uk_K_r7_29 ) , .ZN( u0_uk_n728 ) );
  OAI22_X1 u0_uk_U209 (.B1( decrypt ) , .ZN( u0_K3_14 ) , .A1( u0_uk_n191 ) , .A2( u0_uk_n541 ) , .B2( u0_uk_n548 ) );
  AOI22_X1 u0_uk_U211 (.B1( decrypt ) , .B2( u0_uk_K_r2_31 ) , .A2( u0_uk_K_r2_49 ) , .A1( u0_uk_n242 ) , .ZN( u0_uk_n826 ) );
  OAI22_X1 u0_uk_U212 (.B1( decrypt ) , .ZN( u0_K1_31 ) , .A1( u0_uk_n187 ) , .B2( u0_uk_n707 ) , .A2( u0_uk_n711 ) );
  NAND2_X1 u0_uk_U232 (.A2( decrypt ) , .A1( u0_key_r_15 ) , .ZN( u0_uk_n875 ) );
  OAI22_X1 u0_uk_U238 (.A1( decrypt ) , .ZN( u0_K13_39 ) , .A2( u0_uk_n114 ) , .B2( u0_uk_n133 ) , .B1( u0_uk_n250 ) );
  OAI21_X1 u0_uk_U239 (.B1( decrypt ) , .ZN( u0_K12_39 ) , .B2( u0_uk_n168 ) , .A( u0_uk_n969 ) );
  OAI21_X1 u0_uk_U256 (.B1( decrypt ) , .ZN( u0_K13_48 ) , .B2( u0_uk_n103 ) , .A( u0_uk_n942 ) );
  OAI22_X1 u0_uk_U260 (.A1( decrypt ) , .ZN( u0_K12_48 ) , .B1( u0_uk_n148 ) , .A2( u0_uk_n158 ) , .B2( u0_uk_n167 ) );
  AOI22_X1 u0_uk_U265 (.A1( decrypt ) , .B2( u0_uk_K_r7_16 ) , .A2( u0_uk_K_r7_9 ) , .B1( u0_uk_n202 ) , .ZN( u0_uk_n719 ) );
  OAI22_X1 u0_uk_U270 (.B1( decrypt ) , .ZN( u0_K5_44 ) , .A1( u0_uk_n161 ) , .A2( u0_uk_n463 ) , .B2( u0_uk_n469 ) );
  OAI22_X1 u0_uk_U271 (.B1( decrypt ) , .ZN( u0_K5_48 ) , .A1( u0_uk_n240 ) , .A2( u0_uk_n474 ) , .B2( u0_uk_n481 ) );
  OAI22_X1 u0_uk_U276 (.A1( decrypt ) , .ZN( u0_K2_44 ) , .B1( u0_uk_n147 ) , .A2( u0_uk_n585 ) , .B2( u0_uk_n607 ) );
  NAND2_X1 u0_uk_U281 (.A2( decrypt ) , .A1( u0_uk_K_r4_18 ) , .ZN( u0_uk_n786 ) );
  OAI22_X1 u0_uk_U282 (.A1( decrypt ) , .ZN( u0_K2_6 ) , .B1( u0_uk_n161 ) , .A2( u0_uk_n588 ) , .B2( u0_uk_n609 ) );
  AOI22_X1 u0_uk_U289 (.A1( decrypt ) , .B2( u0_uk_K_r5_26 ) , .A2( u0_uk_K_r5_4 ) , .B1( u0_uk_n202 ) , .ZN( u0_uk_n763 ) );
  OAI21_X1 u0_uk_U294 (.B1( decrypt ) , .ZN( u0_K2_8 ) , .B2( u0_uk_n618 ) , .A( u0_uk_n854 ) );
  NAND2_X1 u0_uk_U295 (.A2( decrypt ) , .A1( u0_uk_K_r0_17 ) , .ZN( u0_uk_n854 ) );
  OAI22_X1 u0_uk_U299 (.B1( decrypt ) , .ZN( u0_K16_8 ) , .A1( u0_uk_n187 ) , .B2( u0_uk_n654 ) , .A2( u0_uk_n667 ) );
  AOI22_X1 u0_uk_U301 (.A1( decrypt ) , .B2( u0_uk_K_r7_15 ) , .A2( u0_uk_K_r7_8 ) , .B1( u0_uk_n217 ) , .ZN( u0_uk_n731 ) );
  NAND2_X1 u0_uk_U311 (.A2( decrypt ) , .A1( u0_uk_K_r11_7 ) , .ZN( u0_uk_n948 ) );
  OAI22_X1 u0_uk_U312 (.B1( decrypt ) , .ZN( u0_K5_26 ) , .A1( u0_uk_n242 ) , .B2( u0_uk_n482 ) , .A2( u0_uk_n492 ) );
  OAI22_X1 u0_uk_U314 (.A1( decrypt ) , .ZN( u0_K16_26 ) , .B1( u0_uk_n182 ) , .A2( u0_uk_n633 ) , .B2( u0_uk_n647 ) );
  OAI22_X1 u0_uk_U321 (.B1( decrypt ) , .ZN( u0_K13_46 ) , .A2( u0_uk_n113 ) , .B2( u0_uk_n125 ) , .A1( u0_uk_n230 ) );
  NAND2_X1 u0_uk_U324 (.A2( decrypt ) , .A1( u0_uk_K_r7_37 ) , .ZN( u0_uk_n720 ) );
  OAI22_X1 u0_uk_U329 (.A1( decrypt ) , .ZN( u0_K2_46 ) , .B1( u0_uk_n147 ) , .B2( u0_uk_n595 ) , .A2( u0_uk_n622 ) );
  OAI21_X1 u0_uk_U330 (.B1( decrypt ) , .ZN( u0_K1_46 ) , .B2( u0_uk_n715 ) , .A( u0_uk_n871 ) );
  AOI22_X1 u0_uk_U334 (.A1( decrypt ) , .B2( u0_uk_K_r5_23 ) , .A2( u0_uk_K_r5_31 ) , .B1( u0_uk_n202 ) , .ZN( u0_uk_n765 ) );
  OAI21_X1 u0_uk_U335 (.B1( decrypt ) , .ZN( u0_K16_4 ) , .B2( u0_uk_n631 ) , .A( u0_uk_n894 ) );
  OAI22_X1 u0_uk_U338 (.A1( decrypt ) , .ZN( u0_K14_4 ) , .B1( u0_uk_n231 ) , .A2( u0_uk_n64 ) , .B2( u0_uk_n72 ) );
  OAI21_X1 u0_uk_U343 (.B1( decrypt ) , .ZN( u0_K5_4 ) , .B2( u0_uk_n477 ) , .A( u0_uk_n804 ) );
  OAI22_X1 u0_uk_U348 (.B1( decrypt ) , .ZN( u0_K2_4 ) , .A1( u0_uk_n209 ) , .A2( u0_uk_n591 ) , .B2( u0_uk_n620 ) );
  OAI21_X1 u0_uk_U358 (.B1( decrypt ) , .ZN( u0_K12_40 ) , .B2( u0_uk_n159 ) , .A( u0_uk_n967 ) );
  NAND2_X1 u0_uk_U359 (.A2( decrypt ) , .A1( u0_uk_K_r10_49 ) , .ZN( u0_uk_n967 ) );
  OAI22_X1 u0_uk_U361 (.A1( decrypt ) , .ZN( u0_K13_40 ) , .A2( u0_uk_n104 ) , .B2( u0_uk_n114 ) , .B1( u0_uk_n147 ) );
  NAND2_X1 u0_uk_U368 (.A2( decrypt ) , .A1( u0_uk_K_r13_31 ) , .ZN( u0_uk_n917 ) );
  OAI21_X1 u0_uk_U376 (.B1( decrypt ) , .ZN( u0_K4_28 ) , .B2( u0_uk_n507 ) , .A( u0_uk_n830 ) );
  NAND2_X1 u0_uk_U377 (.A2( decrypt ) , .A1( u0_uk_K_r2_21 ) , .ZN( u0_uk_n830 ) );
  OAI22_X1 u0_uk_U386 (.B1( decrypt ) , .ZN( u0_K5_28 ) , .A1( u0_uk_n242 ) , .A2( u0_uk_n488 ) , .B2( u0_uk_n492 ) );
  OAI22_X1 u0_uk_U397 (.B1( decrypt ) , .ZN( u0_K6_16 ) , .A1( u0_uk_n213 ) , .A2( u0_uk_n416 ) , .B2( u0_uk_n422 ) );
  NAND2_X1 u0_uk_U399 (.A2( decrypt ) , .A1( u0_uk_K_r1_6 ) , .ZN( u0_uk_n853 ) );
  OAI22_X1 u0_uk_U400 (.A1( decrypt ) , .ZN( u0_K1_16 ) , .B1( u0_uk_n147 ) , .A2( u0_uk_n690 ) , .B2( u0_uk_n696 ) );
  OAI21_X1 u0_uk_U404 (.B1( decrypt ) , .ZN( u0_K14_9 ) , .B2( u0_uk_n70 ) , .A( u0_uk_n926 ) );
  OAI22_X1 u0_uk_U407 (.A1( decrypt ) , .ZN( u0_K12_9 ) , .A2( u0_uk_n136 ) , .B2( u0_uk_n143 ) , .B1( u0_uk_n148 ) );
  AOI22_X1 u0_uk_U413 (.A1( decrypt ) , .B2( u0_uk_K_r8_28 ) , .A2( u0_uk_K_r8_52 ) , .ZN( u0_uk_n1009 ) , .B1( u0_uk_n207 ) );
  AOI22_X1 u0_uk_U427 (.B1( decrypt ) , .B2( u0_key_r_44 ) , .A2( u0_key_r_51 ) , .A1( u0_uk_n222 ) , .ZN( u0_uk_n878 ) );
  OAI22_X1 u0_uk_U428 (.B1( decrypt ) , .ZN( u0_K5_1 ) , .A1( u0_uk_n148 ) , .A2( u0_uk_n459 ) , .B2( u0_uk_n466 ) );
  OAI22_X1 u0_uk_U435 (.B1( decrypt ) , .ZN( u0_K5_16 ) , .A1( u0_uk_n164 ) , .B2( u0_uk_n478 ) , .A2( u0_uk_n491 ) );
  AOI22_X1 u0_uk_U440 (.A1( decrypt ) , .B2( u0_uk_K_r8_22 ) , .A2( u0_uk_K_r8_42 ) , .ZN( u0_uk_n1012 ) , .B1( u0_uk_n207 ) );
  OAI22_X1 u0_uk_U446 (.B1( decrypt ) , .ZN( u0_K8_33 ) , .A1( u0_uk_n257 ) , .A2( u0_uk_n355 ) , .B2( u0_uk_n360 ) );
  OAI21_X1 u0_uk_U457 (.B1( decrypt ) , .ZN( u0_K11_37 ) , .B2( u0_uk_n194 ) , .A( u0_uk_n989 ) );
  NAND2_X1 u0_uk_U460 (.A2( decrypt ) , .A1( u0_uk_K_r7_7 ) , .ZN( u0_uk_n725 ) );
  AOI22_X1 u0_uk_U465 (.A1( decrypt ) , .B2( u0_uk_K_r4_3 ) , .A2( u0_uk_K_r4_41 ) , .B1( u0_uk_n207 ) , .ZN( u0_uk_n785 ) );
  OAI22_X1 u0_uk_U466 (.B1( decrypt ) , .ZN( u0_K5_9 ) , .A1( u0_uk_n223 ) , .A2( u0_uk_n451 ) , .B2( u0_uk_n461 ) );
  OAI21_X1 u0_uk_U470 (.B1( decrypt ) , .ZN( u0_K10_36 ) , .A( u0_uk_n1010 ) , .B2( u0_uk_n269 ) );
  NAND2_X1 u0_uk_U498 (.A2( decrypt ) , .A1( u0_uk_K_r7_53 ) , .ZN( u0_uk_n740 ) );
  AOI22_X1 u0_uk_U507 (.A1( decrypt ) , .B2( u0_uk_K_r6_28 ) , .A2( u0_uk_K_r6_35 ) , .B1( u0_uk_n208 ) , .ZN( u0_uk_n755 ) );
  AOI22_X1 u0_uk_U509 (.A1( decrypt ) , .B2( u0_uk_K_r9_4 ) , .A2( u0_uk_K_r9_55 ) , .ZN( u0_uk_n1001 ) , .B1( u0_uk_n217 ) );
  OAI22_X1 u0_uk_U515 (.B1( decrypt ) , .ZN( u0_K3_17 ) , .A1( u0_uk_n191 ) , .A2( u0_uk_n548 ) , .B2( u0_uk_n571 ) );
  OAI22_X1 u0_uk_U519 (.A1( decrypt ) , .ZN( u0_K14_12 ) , .B1( u0_uk_n238 ) , .A2( u0_uk_n53 ) , .B2( u0_uk_n57 ) );
  NAND2_X1 u0_uk_U521 (.A2( decrypt ) , .A1( u0_uk_K_r10_11 ) , .ZN( u0_uk_n981 ) );
  OAI22_X1 u0_uk_U527 (.B1( decrypt ) , .ZN( u0_K3_12 ) , .A1( u0_uk_n191 ) , .A2( u0_uk_n547 ) , .B2( u0_uk_n552 ) );
  OAI22_X1 u0_uk_U528 (.B1( decrypt ) , .ZN( u0_K2_12 ) , .A1( u0_uk_n164 ) , .B2( u0_uk_n610 ) , .A2( u0_uk_n625 ) );
  OAI22_X1 u0_uk_U546 (.A1( decrypt ) , .ZN( u0_K13_36 ) , .A2( u0_uk_n105 ) , .B2( u0_uk_n111 ) , .B1( u0_uk_n147 ) );
  AOI22_X1 u0_uk_U553 (.A1( decrypt ) , .B2( u0_uk_K_r14_16 ) , .A2( u0_uk_K_r14_23 ) , .B1( u0_uk_n217 ) , .ZN( u0_uk_n904 ) );
  AOI22_X1 u0_uk_U561 (.A1( decrypt ) , .B2( u0_uk_K_r9_15 ) , .A2( u0_uk_K_r9_7 ) , .B1( u0_uk_n217 ) , .ZN( u0_uk_n990 ) );
  AOI22_X1 u0_uk_U563 (.A1( decrypt ) , .B2( u0_uk_K_r13_23 ) , .A2( u0_uk_K_r13_44 ) , .B1( u0_uk_n203 ) , .ZN( u0_uk_n916 ) );
  OAI22_X1 u0_uk_U566 (.B1( decrypt ) , .ZN( u0_K8_36 ) , .A1( u0_uk_n223 ) , .A2( u0_uk_n328 ) , .B2( u0_uk_n334 ) );
  OAI22_X1 u0_uk_U568 (.B1( decrypt ) , .ZN( u0_K5_38 ) , .A1( u0_uk_n240 ) , .A2( u0_uk_n470 ) , .B2( u0_uk_n494 ) );
  OAI22_X1 u0_uk_U569 (.A1( decrypt ) , .ZN( u0_K10_10 ) , .B1( u0_uk_n188 ) , .A2( u0_uk_n235 ) , .B2( u0_uk_n263 ) );
  INV_X1 u0_uk_U57 (.A( decrypt ) , .ZN( u0_uk_n257 ) );
  OAI22_X1 u0_uk_U574 (.A1( decrypt ) , .ZN( u0_K14_10 ) , .B1( u0_uk_n148 ) , .A2( u0_uk_n74 ) , .B2( u0_uk_n79 ) );
  NAND2_X1 u0_uk_U576 (.A2( decrypt ) , .A1( u0_uk_K_r9_54 ) , .ZN( u0_uk_n1004 ) );
  AOI22_X1 u0_uk_U578 (.B1( decrypt ) , .B2( u0_uk_K_r11_26 ) , .A2( u0_uk_K_r11_6 ) , .A1( u0_uk_n238 ) , .ZN( u0_uk_n960 ) );
  AOI22_X1 u0_uk_U585 (.A1( decrypt ) , .B2( u0_uk_K_r2_26 ) , .A2( u0_uk_K_r2_6 ) , .B1( u0_uk_n163 ) , .ZN( u0_uk_n839 ) );
  OAI22_X1 u0_uk_U589 (.B1( decrypt ) , .ZN( u0_K16_22 ) , .A1( u0_uk_n187 ) , .A2( u0_uk_n646 ) , .B2( u0_uk_n653 ) );
  AOI22_X1 u0_uk_U595 (.B1( decrypt ) , .B2( u0_uk_K_r8_27 ) , .A2( u0_uk_K_r8_5 ) , .ZN( u0_uk_n1019 ) , .A1( u0_uk_n162 ) );
  AOI22_X1 u0_uk_U597 (.B1( decrypt ) , .B2( u0_uk_K_r7_41 ) , .A2( u0_uk_K_r7_48 ) , .A1( u0_uk_n240 ) , .ZN( u0_uk_n732 ) );
  AOI22_X1 u0_uk_U600 (.A1( decrypt ) , .B2( u0_uk_K_r3_24 ) , .A2( u0_uk_K_r3_33 ) , .B1( u0_uk_n163 ) , .ZN( u0_uk_n815 ) );
  OAI22_X1 u0_uk_U608 (.A1( decrypt ) , .ZN( u0_K2_35 ) , .B1( u0_uk_n182 ) , .A2( u0_uk_n595 ) , .B2( u0_uk_n613 ) );
  OAI22_X1 u0_uk_U610 (.A1( decrypt ) , .ZN( u0_K12_35 ) , .A2( u0_uk_n151 ) , .B2( u0_uk_n160 ) , .B1( u0_uk_n238 ) );
  AOI22_X1 u0_uk_U617 (.B1( decrypt ) , .B2( u0_uk_K_r7_16 ) , .A2( u0_uk_K_r7_23 ) , .A1( u0_uk_n191 ) , .ZN( u0_uk_n726 ) );
  OAI22_X1 u0_uk_U619 (.B1( decrypt ) , .ZN( u0_K4_35 ) , .A1( u0_uk_n182 ) , .A2( u0_uk_n498 ) , .B2( u0_uk_n527 ) );
  OAI21_X1 u0_uk_U631 (.B1( decrypt ) , .ZN( u0_K8_11 ) , .B2( u0_uk_n323 ) , .A( u0_uk_n762 ) );
  OAI21_X1 u0_uk_U635 (.B1( decrypt ) , .ZN( u0_K2_11 ) , .B2( u0_uk_n591 ) , .A( u0_uk_n867 ) );
  OAI22_X1 u0_uk_U639 (.B1( decrypt ) , .ZN( u0_K6_11 ) , .A1( u0_uk_n213 ) , .A2( u0_uk_n431 ) , .B2( u0_uk_n435 ) );
  OAI22_X1 u0_uk_U648 (.A1( decrypt ) , .ZN( u0_K1_45 ) , .B1( u0_uk_n231 ) , .A2( u0_uk_n680 ) , .B2( u0_uk_n687 ) );
  OAI22_X1 u0_uk_U67 (.A1( decrypt ) , .ZN( u0_K12_34 ) , .B1( u0_uk_n148 ) , .B2( u0_uk_n158 ) , .A2( u0_uk_n173 ) );
  OAI22_X1 u0_uk_U672 (.B1( decrypt ) , .ZN( u0_K9_45 ) , .A1( u0_uk_n257 ) , .A2( u0_uk_n276 ) , .B2( u0_uk_n317 ) );
  NAND2_X1 u0_uk_U674 (.A2( decrypt ) , .A1( u0_uk_K_r3_43 ) , .ZN( u0_uk_n805 ) );
  OAI21_X1 u0_uk_U675 (.B1( decrypt ) , .ZN( u0_K4_43 ) , .B2( u0_uk_n499 ) , .A( u0_uk_n823 ) );
  OAI21_X1 u0_uk_U680 (.B1( decrypt ) , .ZN( u0_K12_7 ) , .B2( u0_uk_n138 ) , .A( u0_uk_n961 ) );
  OAI21_X1 u0_uk_U692 (.B1( decrypt ) , .ZN( u0_K2_25 ) , .B2( u0_uk_n594 ) , .A( u0_uk_n863 ) );
  OAI22_X1 u0_uk_U696 (.A1( decrypt ) , .ZN( u0_K10_25 ) , .B1( u0_uk_n182 ) , .B2( u0_uk_n247 ) , .A2( u0_uk_n265 ) );
  AOI22_X1 u0_uk_U698 (.A1( decrypt ) , .B2( u0_uk_K_r6_21 ) , .A2( u0_uk_K_r6_28 ) , .B1( u0_uk_n217 ) , .ZN( u0_uk_n746 ) );
  AOI22_X1 u0_uk_U705 (.A1( decrypt ) , .B2( u0_uk_K_r11_10 ) , .A2( u0_uk_K_r11_5 ) , .B1( u0_uk_n207 ) , .ZN( u0_uk_n939 ) );
  AOI22_X1 u0_uk_U709 (.A1( decrypt ) , .B2( u0_uk_K_r5_31 ) , .A2( u0_uk_K_r5_7 ) , .B1( u0_uk_n207 ) , .ZN( u0_uk_n775 ) );
  OAI21_X1 u0_uk_U71 (.B1( decrypt ) , .ZN( u0_K3_34 ) , .B2( u0_uk_n559 ) , .A( u0_uk_n848 ) );
  AOI22_X1 u0_uk_U713 (.A1( decrypt ) , .B2( u0_uk_K_r2_16 ) , .A2( u0_uk_K_r2_49 ) , .B1( u0_uk_n203 ) , .ZN( u0_uk_n832 ) );
  OAI22_X1 u0_uk_U723 (.B1( decrypt ) , .ZN( u0_K5_32 ) , .A1( u0_uk_n251 ) , .A2( u0_uk_n476 ) , .B2( u0_uk_n480 ) );
  OAI22_X1 u0_uk_U725 (.A1( decrypt ) , .ZN( u0_K9_32 ) , .B1( u0_uk_n161 ) , .A2( u0_uk_n280 ) , .B2( u0_uk_n287 ) );
  OAI22_X1 u0_uk_U727 (.A1( decrypt ) , .ZN( u0_K14_42 ) , .B1( u0_uk_n147 ) , .A2( u0_uk_n59 ) , .B2( u0_uk_n90 ) );
  OAI22_X1 u0_uk_U728 (.A1( decrypt ) , .ZN( u0_K13_42 ) , .A2( u0_uk_n119 ) , .B2( u0_uk_n125 ) , .B1( u0_uk_n147 ) );
  OAI22_X1 u0_uk_U73 (.B1( decrypt ) , .ZN( u0_K2_34 ) , .A1( u0_uk_n188 ) , .A2( u0_uk_n585 ) , .B2( u0_uk_n616 ) );
  AOI22_X1 u0_uk_U737 (.A1( decrypt ) , .B2( u0_uk_K_r5_1 ) , .A2( u0_uk_K_r5_36 ) , .B1( u0_uk_n202 ) , .ZN( u0_uk_n766 ) );
  OAI21_X1 u0_uk_U744 (.B1( decrypt ) , .ZN( u0_K14_27 ) , .B2( u0_uk_n49 ) , .A( u0_uk_n936 ) );
  OAI21_X1 u0_uk_U747 (.B1( decrypt ) , .ZN( u0_K10_27 ) , .A( u0_uk_n1016 ) , .B2( u0_uk_n256 ) );
  OAI22_X1 u0_uk_U754 (.B1( decrypt ) , .ZN( u0_K6_13 ) , .A1( u0_uk_n238 ) , .A2( u0_uk_n422 ) , .B2( u0_uk_n426 ) );
  NAND2_X1 u0_uk_U758 (.A2( decrypt ) , .A1( u0_uk_K_r7_5 ) , .ZN( u0_uk_n739 ) );
  OAI22_X1 u0_uk_U761 (.A1( decrypt ) , .ZN( u0_K14_21 ) , .B1( u0_uk_n231 ) , .A2( u0_uk_n48 ) , .B2( u0_uk_n74 ) );
  OAI21_X1 u0_uk_U762 (.B1( decrypt ) , .ZN( u0_K11_21 ) , .B2( u0_uk_n221 ) , .A( u0_uk_n998 ) );
  OAI22_X1 u0_uk_U769 (.A1( decrypt ) , .ZN( u0_K14_13 ) , .B1( u0_uk_n148 ) , .A2( u0_uk_n71 ) , .B2( u0_uk_n76 ) );
  OAI22_X1 u0_uk_U770 (.B1( decrypt ) , .ZN( u0_K4_27 ) , .A1( u0_uk_n202 ) , .A2( u0_uk_n512 ) , .B2( u0_uk_n538 ) );
  OAI22_X1 u0_uk_U773 (.B1( decrypt ) , .ZN( u0_K6_27 ) , .A1( u0_uk_n162 ) , .A2( u0_uk_n424 ) , .B2( u0_uk_n429 ) );
  AOI22_X1 u0_uk_U775 (.A1( decrypt ) , .B2( u0_uk_K_r3_15 ) , .A2( u0_uk_K_r3_51 ) , .B1( u0_uk_n217 ) , .ZN( u0_uk_n813 ) );
  AOI22_X1 u0_uk_U783 (.B1( decrypt ) , .B2( u0_uk_K_r11_34 ) , .A2( u0_uk_K_r11_39 ) , .A1( u0_uk_n251 ) , .ZN( u0_uk_n950 ) );
  OAI21_X1 u0_uk_U80 (.B1( decrypt ) , .ZN( u0_K6_23 ) , .B2( u0_uk_n416 ) , .A( u0_uk_n796 ) );
  OAI22_X1 u0_uk_U806 (.B1( decrypt ) , .ZN( u0_K5_18 ) , .A1( u0_uk_n251 ) , .B2( u0_uk_n452 ) , .A2( u0_uk_n489 ) );
  NAND2_X1 u0_uk_U81 (.A2( decrypt ) , .A1( u0_uk_K_r4_27 ) , .ZN( u0_uk_n796 ) );
  OAI21_X1 u0_uk_U815 (.B1( decrypt ) , .ZN( u0_K16_18 ) , .B2( u0_uk_n629 ) , .A( u0_uk_n906 ) );
  OAI22_X1 u0_uk_U817 (.A1( decrypt ) , .ZN( u0_K10_18 ) , .B1( u0_uk_n230 ) , .B2( u0_uk_n254 ) , .A2( u0_uk_n268 ) );
  OAI22_X1 u0_uk_U818 (.A1( decrypt ) , .ZN( u0_K15_18 ) , .B1( u0_uk_n202 ) , .B2( u0_uk_n36 ) , .A2( u0_uk_n6 ) );
  OAI22_X1 u0_uk_U82 (.A1( decrypt ) , .ZN( u0_K3_23 ) , .B1( u0_uk_n242 ) , .B2( u0_uk_n572 ) , .A2( u0_uk_n577 ) );
  AOI22_X1 u0_uk_U826 (.B1( decrypt ) , .B2( u0_uk_K_r7_39 ) , .A2( u0_uk_K_r7_46 ) , .A1( u0_uk_n240 ) , .ZN( u0_uk_n736 ) );
  AOI22_X1 u0_uk_U828 (.A1( decrypt ) , .B2( u0_uk_K_r4_11 ) , .A2( u0_uk_K_r4_17 ) , .B1( u0_uk_n208 ) , .ZN( u0_uk_n799 ) );
  AOI22_X1 u0_uk_U830 (.A1( decrypt ) , .B2( u0_uk_K_r9_10 ) , .A2( u0_uk_K_r9_4 ) , .B1( u0_uk_n163 ) , .ZN( u0_uk_n999 ) );
  AOI22_X1 u0_uk_U834 (.A1( decrypt ) , .B2( u0_uk_K_r5_18 ) , .A2( u0_uk_K_r5_53 ) , .B1( u0_uk_n203 ) , .ZN( u0_uk_n780 ) );
  OAI22_X1 u0_uk_U837 (.A1( decrypt ) , .ZN( u0_K12_22 ) , .A2( u0_uk_n156 ) , .B2( u0_uk_n166 ) , .B1( u0_uk_n222 ) );
  NAND2_X1 u0_uk_U839 (.A2( decrypt ) , .A1( u0_uk_K_r2_47 ) , .ZN( u0_uk_n834 ) );
  OAI22_X1 u0_uk_U851 (.B1( decrypt ) , .ZN( u0_K5_3 ) , .A1( u0_uk_n230 ) , .A2( u0_uk_n477 ) , .B2( u0_uk_n484 ) );
  OAI21_X1 u0_uk_U862 (.B1( decrypt ) , .ZN( u0_K7_2 ) , .B2( u0_uk_n404 ) , .A( u0_uk_n773 ) );
  NAND2_X1 u0_uk_U865 (.A2( decrypt ) , .A1( u0_uk_K_r8_10 ) , .ZN( u0_uk_n1021 ) );
  OAI22_X1 u0_uk_U867 (.B1( decrypt ) , .ZN( u0_K3_18 ) , .A1( u0_uk_n191 ) , .A2( u0_uk_n556 ) , .B2( u0_uk_n563 ) );
  OAI22_X1 u0_uk_U870 (.B1( decrypt ) , .ZN( u0_K5_41 ) , .A1( u0_uk_n220 ) , .A2( u0_uk_n462 ) , .B2( u0_uk_n470 ) );
  OAI22_X1 u0_uk_U872 (.B1( decrypt ) , .ZN( u0_K6_22 ) , .A1( u0_uk_n257 ) , .A2( u0_uk_n436 ) , .B2( u0_uk_n441 ) );
  OAI22_X1 u0_uk_U875 (.B1( decrypt ) , .ZN( u0_K5_23 ) , .A1( u0_uk_n251 ) , .A2( u0_uk_n464 ) , .B2( u0_uk_n473 ) );
  OAI22_X1 u0_uk_U877 (.B1( decrypt ) , .ZN( u0_K5_34 ) , .A1( u0_uk_n240 ) , .B2( u0_uk_n474 ) , .A2( u0_uk_n487 ) );
  OAI22_X1 u0_uk_U885 (.B1( decrypt ) , .ZN( u0_K3_10 ) , .A1( u0_uk_n191 ) , .A2( u0_uk_n567 ) , .B2( u0_uk_n572 ) );
  OAI22_X1 u0_uk_U887 (.B1( decrypt ) , .ZN( u0_K13_45 ) , .B2( u0_uk_n133 ) , .A1( u0_uk_n230 ) , .A2( u0_uk_n95 ) );
  OAI22_X1 u0_uk_U892 (.B1( decrypt ) , .ZN( u0_K8_1 ) , .A1( u0_uk_n257 ) , .B2( u0_uk_n340 ) , .A2( u0_uk_n356 ) );
  OAI22_X1 u0_uk_U901 (.B1( decrypt ) , .ZN( u0_K6_24 ) , .A1( u0_uk_n213 ) , .A2( u0_uk_n427 ) , .B2( u0_uk_n431 ) );
  OAI22_X1 u0_uk_U905 (.B1( decrypt ) , .ZN( u0_K5_19 ) , .A1( u0_uk_n161 ) , .B2( u0_uk_n453 ) , .A2( u0_uk_n490 ) );
  OAI22_X1 u0_uk_U906 (.B1( decrypt ) , .ZN( u0_K5_24 ) , .A1( u0_uk_n202 ) , .A2( u0_uk_n461 ) , .B2( u0_uk_n486 ) );
  OAI22_X1 u0_uk_U910 (.B1( decrypt ) , .ZN( u0_K16_24 ) , .A1( u0_uk_n162 ) , .A2( u0_uk_n659 ) , .B2( u0_uk_n664 ) );
  OAI22_X1 u0_uk_U912 (.B1( decrypt ) , .ZN( u0_K5_13 ) , .A1( u0_uk_n240 ) , .A2( u0_uk_n452 ) , .B2( u0_uk_n483 ) );
  OAI22_X1 u0_uk_U913 (.B1( decrypt ) , .ZN( u0_K5_14 ) , .A1( u0_uk_n222 ) , .A2( u0_uk_n478 ) , .B2( u0_uk_n485 ) );
  OAI22_X1 u0_uk_U920 (.B1( decrypt ) , .ZN( u0_K16_38 ) , .A1( u0_uk_n155 ) , .A2( u0_uk_n641 ) , .B2( u0_uk_n648 ) );
  OAI22_X1 u0_uk_U934 (.A1( decrypt ) , .ZN( u0_K11_48 ) , .A2( u0_uk_n192 ) , .B2( u0_uk_n199 ) , .B1( u0_uk_n202 ) );
  OAI22_X1 u0_uk_U936 (.A1( decrypt ) , .ZN( u0_K9_6 ) , .B1( u0_uk_n155 ) , .A2( u0_uk_n295 ) , .B2( u0_uk_n303 ) );
  OAI22_X1 u0_uk_U943 (.A1( decrypt ) , .ZN( u0_K14_14 ) , .B1( u0_uk_n148 ) , .A2( u0_uk_n47 ) , .B2( u0_uk_n54 ) );
  OAI22_X1 u0_uk_U946 (.A1( decrypt ) , .ZN( u0_K15_47 ) , .A2( u0_uk_n2 ) , .B1( u0_uk_n214 ) , .B2( u0_uk_n34 ) );
  OAI22_X1 u0_uk_U949 (.A1( decrypt ) , .ZN( u0_K10_34 ) , .B1( u0_uk_n182 ) , .A2( u0_uk_n244 ) , .B2( u0_uk_n270 ) );
  OAI22_X1 u0_uk_U953 (.A1( decrypt ) , .ZN( u0_K9_4 ) , .B1( u0_uk_n155 ) , .A2( u0_uk_n302 ) , .B2( u0_uk_n309 ) );
  OAI22_X1 u0_uk_U954 (.A1( decrypt ) , .ZN( u0_K4_48 ) , .B1( u0_uk_n208 ) , .B2( u0_uk_n505 ) , .A2( u0_uk_n533 ) );
  OAI22_X1 u0_uk_U955 (.A1( decrypt ) , .ZN( u0_K2_48 ) , .B1( u0_uk_n182 ) , .A2( u0_uk_n602 ) , .B2( u0_uk_n617 ) );
  OAI22_X1 u0_uk_U958 (.A1( decrypt ) , .ZN( u0_K6_20 ) , .B1( u0_uk_n231 ) , .B2( u0_uk_n444 ) , .A2( u0_uk_n449 ) );
  OAI22_X1 u0_uk_U960 (.A1( decrypt ) , .ZN( u0_K14_18 ) , .B1( u0_uk_n230 ) , .A2( u0_uk_n62 ) , .B2( u0_uk_n70 ) );
  OAI22_X1 u0_uk_U961 (.A1( decrypt ) , .ZN( u0_K16_19 ) , .B1( u0_uk_n187 ) , .A2( u0_uk_n630 ) , .B2( u0_uk_n668 ) );
  OAI22_X1 u0_uk_U963 (.A1( decrypt ) , .ZN( u0_K10_20 ) , .B1( u0_uk_n182 ) , .A2( u0_uk_n229 ) , .B2( u0_uk_n259 ) );
  OAI22_X1 u0_uk_U971 (.A1( decrypt ) , .ZN( u0_K9_40 ) , .B1( u0_uk_n223 ) , .A2( u0_uk_n282 ) , .B2( u0_uk_n288 ) );
  OAI22_X1 u0_uk_U974 (.A1( decrypt ) , .ZN( u0_K8_45 ) , .B1( u0_uk_n213 ) , .A2( u0_uk_n322 ) , .B2( u0_uk_n360 ) );
  OAI22_X1 u0_uk_U979 (.A1( decrypt ) , .ZN( u0_K2_45 ) , .B1( u0_uk_n147 ) , .A2( u0_uk_n584 ) , .B2( u0_uk_n606 ) );
  OAI22_X1 u0_uk_U986 (.A1( decrypt ) , .ZN( u0_K9_15 ) , .B1( u0_uk_n240 ) , .A2( u0_uk_n304 ) , .B2( u0_uk_n311 ) );
  OAI22_X1 u0_uk_U990 (.A1( decrypt ) , .ZN( u0_K1_23 ) , .B1( u0_uk_n222 ) , .A2( u0_uk_n684 ) , .B2( u0_uk_n691 ) );
  OAI21_X1 u0_uk_U994 (.B1( decrypt ) , .ZN( u0_K7_22 ) , .B2( u0_uk_n390 ) , .A( u0_uk_n778 ) );
  OAI21_X1 u0_uk_U996 (.B1( decrypt ) , .ZN( u0_K7_23 ) , .B2( u0_uk_n405 ) , .A( u0_uk_n777 ) );
  DFF_X1 u1_L0_reg_1 (.CK( clk ) , .Q( u1_L0_1 ) , .D( u1_desIn_r_7 ) );
  DFF_X1 u1_L0_reg_10 (.CK( clk ) , .Q( u1_L0_10 ) , .D( u1_desIn_r_13 ) );
  DFF_X1 u1_L0_reg_11 (.CK( clk ) , .Q( u1_L0_11 ) , .D( u1_desIn_r_21 ) );
  DFF_X1 u1_L0_reg_12 (.CK( clk ) , .Q( u1_L0_12 ) , .D( u1_desIn_r_29 ) );
  DFF_X1 u1_L0_reg_13 (.CK( clk ) , .Q( u1_L0_13 ) , .D( u1_desIn_r_37 ) );
  DFF_X1 u1_L0_reg_14 (.CK( clk ) , .Q( u1_L0_14 ) , .D( u1_desIn_r_45 ) );
  DFF_X1 u1_L0_reg_15 (.CK( clk ) , .Q( u1_L0_15 ) , .D( u1_desIn_r_53 ) );
  DFF_X1 u1_L0_reg_16 (.CK( clk ) , .Q( u1_L0_16 ) , .D( u1_desIn_r_61 ) );
  DFF_X1 u1_L0_reg_17 (.CK( clk ) , .Q( u1_L0_17 ) , .D( u1_desIn_r_3 ) );
  DFF_X1 u1_L0_reg_18 (.CK( clk ) , .Q( u1_L0_18 ) , .D( u1_desIn_r_11 ) );
  DFF_X1 u1_L0_reg_19 (.CK( clk ) , .Q( u1_L0_19 ) , .D( u1_desIn_r_19 ) );
  DFF_X1 u1_L0_reg_2 (.CK( clk ) , .Q( u1_L0_2 ) , .D( u1_desIn_r_15 ) );
  DFF_X1 u1_L0_reg_20 (.CK( clk ) , .Q( u1_L0_20 ) , .D( u1_desIn_r_27 ) );
  DFF_X1 u1_L0_reg_21 (.CK( clk ) , .Q( u1_L0_21 ) , .D( u1_desIn_r_35 ) );
  DFF_X1 u1_L0_reg_22 (.CK( clk ) , .Q( u1_L0_22 ) , .D( u1_desIn_r_43 ) );
  DFF_X1 u1_L0_reg_23 (.CK( clk ) , .Q( u1_L0_23 ) , .D( u1_desIn_r_51 ) );
  DFF_X1 u1_L0_reg_24 (.CK( clk ) , .Q( u1_L0_24 ) , .D( u1_desIn_r_59 ) );
  DFF_X1 u1_L0_reg_25 (.CK( clk ) , .Q( u1_L0_25 ) , .D( u1_desIn_r_1 ) );
  DFF_X1 u1_L0_reg_26 (.CK( clk ) , .Q( u1_L0_26 ) , .D( u1_desIn_r_9 ) );
  DFF_X1 u1_L0_reg_27 (.CK( clk ) , .Q( u1_L0_27 ) , .D( u1_desIn_r_17 ) );
  DFF_X1 u1_L0_reg_28 (.CK( clk ) , .Q( u1_L0_28 ) , .D( u1_desIn_r_25 ) );
  DFF_X1 u1_L0_reg_29 (.CK( clk ) , .Q( u1_L0_29 ) , .D( u1_desIn_r_33 ) );
  DFF_X1 u1_L0_reg_3 (.CK( clk ) , .Q( u1_L0_3 ) , .D( u1_desIn_r_23 ) );
  DFF_X1 u1_L0_reg_30 (.CK( clk ) , .Q( u1_L0_30 ) , .D( u1_desIn_r_41 ) );
  DFF_X1 u1_L0_reg_31 (.CK( clk ) , .Q( u1_L0_31 ) , .D( u1_desIn_r_49 ) );
  DFF_X1 u1_L0_reg_32 (.CK( clk ) , .Q( u1_L0_32 ) , .D( u1_desIn_r_57 ) );
  DFF_X1 u1_L0_reg_4 (.CK( clk ) , .Q( u1_L0_4 ) , .D( u1_desIn_r_31 ) );
  DFF_X1 u1_L0_reg_5 (.CK( clk ) , .Q( u1_L0_5 ) , .D( u1_desIn_r_39 ) );
  DFF_X1 u1_L0_reg_6 (.CK( clk ) , .Q( u1_L0_6 ) , .D( u1_desIn_r_47 ) );
  DFF_X1 u1_L0_reg_7 (.CK( clk ) , .Q( u1_L0_7 ) , .D( u1_desIn_r_55 ) );
  DFF_X1 u1_L0_reg_8 (.CK( clk ) , .Q( u1_L0_8 ) , .D( u1_desIn_r_63 ) );
  DFF_X1 u1_L0_reg_9 (.CK( clk ) , .Q( u1_L0_9 ) , .D( u1_desIn_r_5 ) );
  DFF_X1 u1_L10_reg_1 (.CK( clk ) , .Q( u1_L10_1 ) , .D( u1_R9_1 ) );
  DFF_X1 u1_L10_reg_10 (.CK( clk ) , .Q( u1_L10_10 ) , .D( u1_R9_10 ) );
  DFF_X1 u1_L10_reg_11 (.CK( clk ) , .Q( u1_L10_11 ) , .D( u1_R9_11 ) );
  DFF_X1 u1_L10_reg_12 (.CK( clk ) , .Q( u1_L10_12 ) , .D( u1_R9_12 ) );
  DFF_X1 u1_L10_reg_13 (.CK( clk ) , .Q( u1_L10_13 ) , .D( u1_R9_13 ) );
  DFF_X1 u1_L10_reg_14 (.CK( clk ) , .Q( u1_L10_14 ) , .D( u1_R9_14 ) );
  DFF_X1 u1_L10_reg_15 (.CK( clk ) , .Q( u1_L10_15 ) , .D( u1_R9_15 ) );
  DFF_X1 u1_L10_reg_16 (.CK( clk ) , .Q( u1_L10_16 ) , .D( u1_R9_16 ) );
  DFF_X1 u1_L10_reg_17 (.CK( clk ) , .Q( u1_L10_17 ) , .D( u1_R9_17 ) );
  DFF_X1 u1_L10_reg_18 (.CK( clk ) , .Q( u1_L10_18 ) , .D( u1_R9_18 ) );
  DFF_X1 u1_L10_reg_19 (.CK( clk ) , .Q( u1_L10_19 ) , .D( u1_R9_19 ) );
  DFF_X1 u1_L10_reg_2 (.CK( clk ) , .Q( u1_L10_2 ) , .D( u1_R9_2 ) );
  DFF_X1 u1_L10_reg_20 (.CK( clk ) , .Q( u1_L10_20 ) , .D( u1_R9_20 ) );
  DFF_X1 u1_L10_reg_21 (.CK( clk ) , .Q( u1_L10_21 ) , .D( u1_R9_21 ) );
  DFF_X1 u1_L10_reg_22 (.CK( clk ) , .Q( u1_L10_22 ) , .D( u1_R9_22 ) );
  DFF_X1 u1_L10_reg_23 (.CK( clk ) , .Q( u1_L10_23 ) , .D( u1_R9_23 ) );
  DFF_X1 u1_L10_reg_24 (.CK( clk ) , .Q( u1_L10_24 ) , .D( u1_R9_24 ) );
  DFF_X1 u1_L10_reg_25 (.CK( clk ) , .Q( u1_L10_25 ) , .D( u1_R9_25 ) );
  DFF_X1 u1_L10_reg_26 (.CK( clk ) , .Q( u1_L10_26 ) , .D( u1_R9_26 ) );
  DFF_X1 u1_L10_reg_27 (.CK( clk ) , .Q( u1_L10_27 ) , .D( u1_R9_27 ) );
  DFF_X1 u1_L10_reg_28 (.CK( clk ) , .Q( u1_L10_28 ) , .D( u1_R9_28 ) );
  DFF_X1 u1_L10_reg_29 (.CK( clk ) , .Q( u1_L10_29 ) , .D( u1_R9_29 ) );
  DFF_X1 u1_L10_reg_3 (.CK( clk ) , .Q( u1_L10_3 ) , .D( u1_R9_3 ) );
  DFF_X1 u1_L10_reg_30 (.CK( clk ) , .Q( u1_L10_30 ) , .D( u1_R9_30 ) );
  DFF_X1 u1_L10_reg_31 (.CK( clk ) , .Q( u1_L10_31 ) , .D( u1_R9_31 ) );
  DFF_X1 u1_L10_reg_32 (.CK( clk ) , .Q( u1_L10_32 ) , .D( u1_R9_32 ) );
  DFF_X1 u1_L10_reg_4 (.CK( clk ) , .Q( u1_L10_4 ) , .D( u1_R9_4 ) );
  DFF_X1 u1_L10_reg_5 (.CK( clk ) , .Q( u1_L10_5 ) , .D( u1_R9_5 ) );
  DFF_X1 u1_L10_reg_6 (.CK( clk ) , .Q( u1_L10_6 ) , .D( u1_R9_6 ) );
  DFF_X1 u1_L10_reg_7 (.CK( clk ) , .Q( u1_L10_7 ) , .D( u1_R9_7 ) );
  DFF_X1 u1_L10_reg_8 (.CK( clk ) , .Q( u1_L10_8 ) , .D( u1_R9_8 ) );
  DFF_X1 u1_L10_reg_9 (.CK( clk ) , .Q( u1_L10_9 ) , .D( u1_R9_9 ) );
  DFF_X1 u1_L11_reg_1 (.CK( clk ) , .Q( u1_L11_1 ) , .D( u1_R10_1 ) );
  DFF_X1 u1_L11_reg_10 (.CK( clk ) , .Q( u1_L11_10 ) , .D( u1_R10_10 ) );
  DFF_X1 u1_L11_reg_11 (.CK( clk ) , .Q( u1_L11_11 ) , .D( u1_R10_11 ) );
  DFF_X1 u1_L11_reg_12 (.CK( clk ) , .Q( u1_L11_12 ) , .D( u1_R10_12 ) );
  DFF_X1 u1_L11_reg_13 (.CK( clk ) , .Q( u1_L11_13 ) , .D( u1_R10_13 ) );
  DFF_X1 u1_L11_reg_14 (.CK( clk ) , .Q( u1_L11_14 ) , .D( u1_R10_14 ) );
  DFF_X1 u1_L11_reg_15 (.CK( clk ) , .Q( u1_L11_15 ) , .D( u1_R10_15 ) );
  DFF_X1 u1_L11_reg_16 (.CK( clk ) , .Q( u1_L11_16 ) , .D( u1_R10_16 ) );
  DFF_X1 u1_L11_reg_17 (.CK( clk ) , .Q( u1_L11_17 ) , .D( u1_R10_17 ) );
  DFF_X1 u1_L11_reg_18 (.CK( clk ) , .Q( u1_L11_18 ) , .D( u1_R10_18 ) );
  DFF_X1 u1_L11_reg_19 (.CK( clk ) , .Q( u1_L11_19 ) , .D( u1_R10_19 ) );
  DFF_X1 u1_L11_reg_2 (.CK( clk ) , .Q( u1_L11_2 ) , .D( u1_R10_2 ) );
  DFF_X1 u1_L11_reg_20 (.CK( clk ) , .Q( u1_L11_20 ) , .D( u1_R10_20 ) );
  DFF_X1 u1_L11_reg_21 (.CK( clk ) , .Q( u1_L11_21 ) , .D( u1_R10_21 ) );
  DFF_X1 u1_L11_reg_22 (.CK( clk ) , .Q( u1_L11_22 ) , .D( u1_R10_22 ) );
  DFF_X1 u1_L11_reg_23 (.CK( clk ) , .Q( u1_L11_23 ) , .D( u1_R10_23 ) );
  DFF_X1 u1_L11_reg_24 (.CK( clk ) , .Q( u1_L11_24 ) , .D( u1_R10_24 ) );
  DFF_X1 u1_L11_reg_25 (.CK( clk ) , .Q( u1_L11_25 ) , .D( u1_R10_25 ) );
  DFF_X1 u1_L11_reg_26 (.CK( clk ) , .Q( u1_L11_26 ) , .D( u1_R10_26 ) );
  DFF_X1 u1_L11_reg_27 (.CK( clk ) , .Q( u1_L11_27 ) , .D( u1_R10_27 ) );
  DFF_X1 u1_L11_reg_28 (.CK( clk ) , .Q( u1_L11_28 ) , .D( u1_R10_28 ) );
  DFF_X1 u1_L11_reg_29 (.CK( clk ) , .Q( u1_L11_29 ) , .D( u1_R10_29 ) );
  DFF_X1 u1_L11_reg_3 (.CK( clk ) , .Q( u1_L11_3 ) , .D( u1_R10_3 ) );
  DFF_X1 u1_L11_reg_30 (.CK( clk ) , .Q( u1_L11_30 ) , .D( u1_R10_30 ) );
  DFF_X1 u1_L11_reg_31 (.CK( clk ) , .Q( u1_L11_31 ) , .D( u1_R10_31 ) );
  DFF_X1 u1_L11_reg_32 (.CK( clk ) , .Q( u1_L11_32 ) , .D( u1_R10_32 ) );
  DFF_X1 u1_L11_reg_4 (.CK( clk ) , .Q( u1_L11_4 ) , .D( u1_R10_4 ) );
  DFF_X1 u1_L11_reg_5 (.CK( clk ) , .Q( u1_L11_5 ) , .D( u1_R10_5 ) );
  DFF_X1 u1_L11_reg_6 (.CK( clk ) , .Q( u1_L11_6 ) , .D( u1_R10_6 ) );
  DFF_X1 u1_L11_reg_7 (.CK( clk ) , .Q( u1_L11_7 ) , .D( u1_R10_7 ) );
  DFF_X1 u1_L11_reg_8 (.CK( clk ) , .Q( u1_L11_8 ) , .D( u1_R10_8 ) );
  DFF_X1 u1_L11_reg_9 (.CK( clk ) , .Q( u1_L11_9 ) , .D( u1_R10_9 ) );
  DFF_X1 u1_L12_reg_1 (.CK( clk ) , .Q( u1_L12_1 ) , .D( u1_R11_1 ) );
  DFF_X1 u1_L12_reg_10 (.CK( clk ) , .Q( u1_L12_10 ) , .D( u1_R11_10 ) );
  DFF_X1 u1_L12_reg_11 (.CK( clk ) , .Q( u1_L12_11 ) , .D( u1_R11_11 ) );
  DFF_X1 u1_L12_reg_12 (.CK( clk ) , .Q( u1_L12_12 ) , .D( u1_R11_12 ) );
  DFF_X1 u1_L12_reg_13 (.CK( clk ) , .Q( u1_L12_13 ) , .D( u1_R11_13 ) );
  DFF_X1 u1_L12_reg_14 (.CK( clk ) , .Q( u1_L12_14 ) , .D( u1_R11_14 ) );
  DFF_X1 u1_L12_reg_15 (.CK( clk ) , .Q( u1_L12_15 ) , .D( u1_R11_15 ) );
  DFF_X1 u1_L12_reg_16 (.CK( clk ) , .Q( u1_L12_16 ) , .D( u1_R11_16 ) );
  DFF_X1 u1_L12_reg_17 (.CK( clk ) , .Q( u1_L12_17 ) , .D( u1_R11_17 ) );
  DFF_X1 u1_L12_reg_18 (.CK( clk ) , .Q( u1_L12_18 ) , .D( u1_R11_18 ) );
  DFF_X1 u1_L12_reg_19 (.CK( clk ) , .Q( u1_L12_19 ) , .D( u1_R11_19 ) );
  DFF_X1 u1_L12_reg_2 (.CK( clk ) , .Q( u1_L12_2 ) , .D( u1_R11_2 ) );
  DFF_X1 u1_L12_reg_20 (.CK( clk ) , .Q( u1_L12_20 ) , .D( u1_R11_20 ) );
  DFF_X1 u1_L12_reg_21 (.CK( clk ) , .Q( u1_L12_21 ) , .D( u1_R11_21 ) );
  DFF_X1 u1_L12_reg_22 (.CK( clk ) , .Q( u1_L12_22 ) , .D( u1_R11_22 ) );
  DFF_X1 u1_L12_reg_23 (.CK( clk ) , .Q( u1_L12_23 ) , .D( u1_R11_23 ) );
  DFF_X1 u1_L12_reg_24 (.CK( clk ) , .Q( u1_L12_24 ) , .D( u1_R11_24 ) );
  DFF_X1 u1_L12_reg_25 (.CK( clk ) , .Q( u1_L12_25 ) , .D( u1_R11_25 ) );
  DFF_X1 u1_L12_reg_26 (.CK( clk ) , .Q( u1_L12_26 ) , .D( u1_R11_26 ) );
  DFF_X1 u1_L12_reg_27 (.CK( clk ) , .Q( u1_L12_27 ) , .D( u1_R11_27 ) );
  DFF_X1 u1_L12_reg_28 (.CK( clk ) , .Q( u1_L12_28 ) , .D( u1_R11_28 ) );
  DFF_X1 u1_L12_reg_29 (.CK( clk ) , .Q( u1_L12_29 ) , .D( u1_R11_29 ) );
  DFF_X1 u1_L12_reg_3 (.CK( clk ) , .Q( u1_L12_3 ) , .D( u1_R11_3 ) );
  DFF_X1 u1_L12_reg_30 (.CK( clk ) , .Q( u1_L12_30 ) , .D( u1_R11_30 ) );
  DFF_X1 u1_L12_reg_31 (.CK( clk ) , .Q( u1_L12_31 ) , .D( u1_R11_31 ) );
  DFF_X1 u1_L12_reg_32 (.CK( clk ) , .Q( u1_L12_32 ) , .D( u1_R11_32 ) );
  DFF_X1 u1_L12_reg_4 (.CK( clk ) , .Q( u1_L12_4 ) , .D( u1_R11_4 ) );
  DFF_X1 u1_L12_reg_5 (.CK( clk ) , .Q( u1_L12_5 ) , .D( u1_R11_5 ) );
  DFF_X1 u1_L12_reg_6 (.CK( clk ) , .Q( u1_L12_6 ) , .D( u1_R11_6 ) );
  DFF_X1 u1_L12_reg_7 (.CK( clk ) , .Q( u1_L12_7 ) , .D( u1_R11_7 ) );
  DFF_X1 u1_L12_reg_8 (.CK( clk ) , .Q( u1_L12_8 ) , .D( u1_R11_8 ) );
  DFF_X1 u1_L12_reg_9 (.CK( clk ) , .Q( u1_L12_9 ) , .D( u1_R11_9 ) );
  DFF_X1 u1_L13_reg_1 (.CK( clk ) , .Q( u1_L13_1 ) , .D( u1_R12_1 ) );
  DFF_X1 u1_L13_reg_10 (.CK( clk ) , .Q( u1_L13_10 ) , .D( u1_R12_10 ) );
  DFF_X1 u1_L13_reg_11 (.CK( clk ) , .Q( u1_L13_11 ) , .D( u1_R12_11 ) );
  DFF_X1 u1_L13_reg_12 (.CK( clk ) , .Q( u1_L13_12 ) , .D( u1_R12_12 ) );
  DFF_X1 u1_L13_reg_13 (.CK( clk ) , .Q( u1_L13_13 ) , .D( u1_R12_13 ) );
  DFF_X1 u1_L13_reg_14 (.CK( clk ) , .Q( u1_L13_14 ) , .D( u1_R12_14 ) );
  DFF_X1 u1_L13_reg_15 (.CK( clk ) , .Q( u1_L13_15 ) , .D( u1_R12_15 ) );
  DFF_X1 u1_L13_reg_16 (.CK( clk ) , .Q( u1_L13_16 ) , .D( u1_R12_16 ) );
  DFF_X1 u1_L13_reg_17 (.CK( clk ) , .Q( u1_L13_17 ) , .D( u1_R12_17 ) );
  DFF_X1 u1_L13_reg_18 (.CK( clk ) , .Q( u1_L13_18 ) , .D( u1_R12_18 ) );
  DFF_X1 u1_L13_reg_19 (.CK( clk ) , .Q( u1_L13_19 ) , .D( u1_R12_19 ) );
  DFF_X1 u1_L13_reg_2 (.CK( clk ) , .Q( u1_L13_2 ) , .D( u1_R12_2 ) );
  DFF_X1 u1_L13_reg_20 (.CK( clk ) , .Q( u1_L13_20 ) , .D( u1_R12_20 ) );
  DFF_X1 u1_L13_reg_21 (.CK( clk ) , .Q( u1_L13_21 ) , .D( u1_R12_21 ) );
  DFF_X1 u1_L13_reg_22 (.CK( clk ) , .Q( u1_L13_22 ) , .D( u1_R12_22 ) );
  DFF_X1 u1_L13_reg_23 (.CK( clk ) , .Q( u1_L13_23 ) , .D( u1_R12_23 ) );
  DFF_X1 u1_L13_reg_24 (.CK( clk ) , .Q( u1_L13_24 ) , .D( u1_R12_24 ) );
  DFF_X1 u1_L13_reg_25 (.CK( clk ) , .Q( u1_L13_25 ) , .D( u1_R12_25 ) );
  DFF_X1 u1_L13_reg_26 (.CK( clk ) , .Q( u1_L13_26 ) , .D( u1_R12_26 ) );
  DFF_X1 u1_L13_reg_27 (.CK( clk ) , .Q( u1_L13_27 ) , .D( u1_R12_27 ) );
  DFF_X1 u1_L13_reg_28 (.CK( clk ) , .Q( u1_L13_28 ) , .D( u1_R12_28 ) );
  DFF_X1 u1_L13_reg_29 (.CK( clk ) , .Q( u1_L13_29 ) , .D( u1_R12_29 ) );
  DFF_X1 u1_L13_reg_3 (.CK( clk ) , .Q( u1_L13_3 ) , .D( u1_R12_3 ) );
  DFF_X1 u1_L13_reg_30 (.CK( clk ) , .Q( u1_L13_30 ) , .D( u1_R12_30 ) );
  DFF_X1 u1_L13_reg_31 (.CK( clk ) , .Q( u1_L13_31 ) , .D( u1_R12_31 ) );
  DFF_X1 u1_L13_reg_32 (.CK( clk ) , .Q( u1_L13_32 ) , .D( u1_R12_32 ) );
  DFF_X1 u1_L13_reg_4 (.CK( clk ) , .Q( u1_L13_4 ) , .D( u1_R12_4 ) );
  DFF_X1 u1_L13_reg_5 (.CK( clk ) , .Q( u1_L13_5 ) , .D( u1_R12_5 ) );
  DFF_X1 u1_L13_reg_6 (.CK( clk ) , .Q( u1_L13_6 ) , .D( u1_R12_6 ) );
  DFF_X1 u1_L13_reg_7 (.CK( clk ) , .Q( u1_L13_7 ) , .D( u1_R12_7 ) );
  DFF_X1 u1_L13_reg_8 (.CK( clk ) , .Q( u1_L13_8 ) , .D( u1_R12_8 ) );
  DFF_X1 u1_L13_reg_9 (.CK( clk ) , .Q( u1_L13_9 ) , .D( u1_R12_9 ) );
  DFF_X1 u1_L14_reg_1 (.CK( clk ) , .Q( u1_L14_1 ) , .D( u1_R13_1 ) );
  DFF_X1 u1_L14_reg_10 (.CK( clk ) , .Q( u1_L14_10 ) , .D( u1_R13_10 ) );
  DFF_X1 u1_L14_reg_11 (.CK( clk ) , .Q( u1_L14_11 ) , .D( u1_R13_11 ) );
  DFF_X1 u1_L14_reg_12 (.CK( clk ) , .Q( u1_L14_12 ) , .D( u1_R13_12 ) );
  DFF_X1 u1_L14_reg_13 (.CK( clk ) , .Q( u1_L14_13 ) , .D( u1_R13_13 ) );
  DFF_X1 u1_L14_reg_14 (.CK( clk ) , .Q( u1_L14_14 ) , .D( u1_R13_14 ) );
  DFF_X1 u1_L14_reg_15 (.CK( clk ) , .Q( u1_L14_15 ) , .D( u1_R13_15 ) );
  DFF_X1 u1_L14_reg_16 (.CK( clk ) , .Q( u1_L14_16 ) , .D( u1_R13_16 ) );
  DFF_X1 u1_L14_reg_17 (.CK( clk ) , .Q( u1_L14_17 ) , .D( u1_R13_17 ) );
  DFF_X1 u1_L14_reg_18 (.CK( clk ) , .Q( u1_L14_18 ) , .D( u1_R13_18 ) );
  DFF_X1 u1_L14_reg_19 (.CK( clk ) , .Q( u1_L14_19 ) , .D( u1_R13_19 ) );
  DFF_X1 u1_L14_reg_2 (.CK( clk ) , .Q( u1_L14_2 ) , .D( u1_R13_2 ) );
  DFF_X1 u1_L14_reg_20 (.CK( clk ) , .Q( u1_L14_20 ) , .D( u1_R13_20 ) );
  DFF_X1 u1_L14_reg_21 (.CK( clk ) , .Q( u1_L14_21 ) , .D( u1_R13_21 ) );
  DFF_X1 u1_L14_reg_22 (.CK( clk ) , .Q( u1_L14_22 ) , .D( u1_R13_22 ) );
  DFF_X1 u1_L14_reg_23 (.CK( clk ) , .Q( u1_L14_23 ) , .D( u1_R13_23 ) );
  DFF_X1 u1_L14_reg_24 (.CK( clk ) , .Q( u1_L14_24 ) , .D( u1_R13_24 ) );
  DFF_X1 u1_L14_reg_25 (.CK( clk ) , .Q( u1_L14_25 ) , .D( u1_R13_25 ) );
  DFF_X1 u1_L14_reg_26 (.CK( clk ) , .Q( u1_L14_26 ) , .D( u1_R13_26 ) );
  DFF_X1 u1_L14_reg_27 (.CK( clk ) , .Q( u1_L14_27 ) , .D( u1_R13_27 ) );
  DFF_X1 u1_L14_reg_28 (.CK( clk ) , .Q( u1_L14_28 ) , .D( u1_R13_28 ) );
  DFF_X1 u1_L14_reg_29 (.CK( clk ) , .Q( u1_L14_29 ) , .D( u1_R13_29 ) );
  DFF_X1 u1_L14_reg_3 (.CK( clk ) , .Q( u1_L14_3 ) , .D( u1_R13_3 ) );
  DFF_X1 u1_L14_reg_30 (.CK( clk ) , .Q( u1_L14_30 ) , .D( u1_R13_30 ) );
  DFF_X1 u1_L14_reg_31 (.CK( clk ) , .Q( u1_L14_31 ) , .D( u1_R13_31 ) );
  DFF_X1 u1_L14_reg_32 (.CK( clk ) , .Q( u1_L14_32 ) , .D( u1_R13_32 ) );
  DFF_X1 u1_L14_reg_4 (.CK( clk ) , .Q( u1_L14_4 ) , .D( u1_R13_4 ) );
  DFF_X1 u1_L14_reg_5 (.CK( clk ) , .Q( u1_L14_5 ) , .D( u1_R13_5 ) );
  DFF_X1 u1_L14_reg_6 (.CK( clk ) , .Q( u1_L14_6 ) , .D( u1_R13_6 ) );
  DFF_X1 u1_L14_reg_7 (.CK( clk ) , .Q( u1_L14_7 ) , .D( u1_R13_7 ) );
  DFF_X1 u1_L14_reg_8 (.CK( clk ) , .Q( u1_L14_8 ) , .D( u1_R13_8 ) );
  DFF_X1 u1_L14_reg_9 (.CK( clk ) , .Q( u1_L14_9 ) , .D( u1_R13_9 ) );
  DFF_X1 u1_L1_reg_1 (.CK( clk ) , .Q( u1_L1_1 ) , .D( u1_R0_1 ) );
  DFF_X1 u1_L1_reg_10 (.CK( clk ) , .Q( u1_L1_10 ) , .D( u1_R0_10 ) );
  DFF_X1 u1_L1_reg_11 (.CK( clk ) , .Q( u1_L1_11 ) , .D( u1_R0_11 ) );
  DFF_X1 u1_L1_reg_12 (.CK( clk ) , .Q( u1_L1_12 ) , .D( u1_R0_12 ) );
  DFF_X1 u1_L1_reg_13 (.CK( clk ) , .Q( u1_L1_13 ) , .D( u1_R0_13 ) );
  DFF_X1 u1_L1_reg_14 (.CK( clk ) , .Q( u1_L1_14 ) , .D( u1_R0_14 ) );
  DFF_X1 u1_L1_reg_15 (.CK( clk ) , .Q( u1_L1_15 ) , .D( u1_R0_15 ) );
  DFF_X1 u1_L1_reg_16 (.CK( clk ) , .Q( u1_L1_16 ) , .D( u1_R0_16 ) );
  DFF_X1 u1_L1_reg_17 (.CK( clk ) , .Q( u1_L1_17 ) , .D( u1_R0_17 ) );
  DFF_X1 u1_L1_reg_18 (.CK( clk ) , .Q( u1_L1_18 ) , .D( u1_R0_18 ) );
  DFF_X1 u1_L1_reg_19 (.CK( clk ) , .Q( u1_L1_19 ) , .D( u1_R0_19 ) );
  DFF_X1 u1_L1_reg_2 (.CK( clk ) , .Q( u1_L1_2 ) , .D( u1_R0_2 ) );
  DFF_X1 u1_L1_reg_20 (.CK( clk ) , .Q( u1_L1_20 ) , .D( u1_R0_20 ) );
  DFF_X1 u1_L1_reg_21 (.CK( clk ) , .Q( u1_L1_21 ) , .D( u1_R0_21 ) );
  DFF_X1 u1_L1_reg_22 (.CK( clk ) , .Q( u1_L1_22 ) , .D( u1_R0_22 ) );
  DFF_X1 u1_L1_reg_23 (.CK( clk ) , .Q( u1_L1_23 ) , .D( u1_R0_23 ) );
  DFF_X1 u1_L1_reg_24 (.CK( clk ) , .Q( u1_L1_24 ) , .D( u1_R0_24 ) );
  DFF_X1 u1_L1_reg_25 (.CK( clk ) , .Q( u1_L1_25 ) , .D( u1_R0_25 ) );
  DFF_X1 u1_L1_reg_26 (.CK( clk ) , .Q( u1_L1_26 ) , .D( u1_R0_26 ) );
  DFF_X1 u1_L1_reg_27 (.CK( clk ) , .Q( u1_L1_27 ) , .D( u1_R0_27 ) );
  DFF_X1 u1_L1_reg_28 (.CK( clk ) , .Q( u1_L1_28 ) , .D( u1_R0_28 ) );
  DFF_X1 u1_L1_reg_29 (.CK( clk ) , .Q( u1_L1_29 ) , .D( u1_R0_29 ) );
  DFF_X1 u1_L1_reg_3 (.CK( clk ) , .Q( u1_L1_3 ) , .D( u1_R0_3 ) );
  DFF_X1 u1_L1_reg_30 (.CK( clk ) , .Q( u1_L1_30 ) , .D( u1_R0_30 ) );
  DFF_X1 u1_L1_reg_31 (.CK( clk ) , .Q( u1_L1_31 ) , .D( u1_R0_31 ) );
  DFF_X1 u1_L1_reg_32 (.CK( clk ) , .Q( u1_L1_32 ) , .D( u1_R0_32 ) );
  DFF_X1 u1_L1_reg_4 (.CK( clk ) , .Q( u1_L1_4 ) , .D( u1_R0_4 ) );
  DFF_X1 u1_L1_reg_5 (.CK( clk ) , .Q( u1_L1_5 ) , .D( u1_R0_5 ) );
  DFF_X1 u1_L1_reg_6 (.CK( clk ) , .Q( u1_L1_6 ) , .D( u1_R0_6 ) );
  DFF_X1 u1_L1_reg_7 (.CK( clk ) , .Q( u1_L1_7 ) , .D( u1_R0_7 ) );
  DFF_X1 u1_L1_reg_8 (.CK( clk ) , .Q( u1_L1_8 ) , .D( u1_R0_8 ) );
  DFF_X1 u1_L1_reg_9 (.CK( clk ) , .Q( u1_L1_9 ) , .D( u1_R0_9 ) );
  DFF_X1 u1_L2_reg_1 (.CK( clk ) , .Q( u1_L2_1 ) , .D( u1_R1_1 ) );
  DFF_X1 u1_L2_reg_10 (.CK( clk ) , .Q( u1_L2_10 ) , .D( u1_R1_10 ) );
  DFF_X1 u1_L2_reg_11 (.CK( clk ) , .Q( u1_L2_11 ) , .D( u1_R1_11 ) );
  DFF_X1 u1_L2_reg_12 (.CK( clk ) , .Q( u1_L2_12 ) , .D( u1_R1_12 ) );
  DFF_X1 u1_L2_reg_13 (.CK( clk ) , .Q( u1_L2_13 ) , .D( u1_R1_13 ) );
  DFF_X1 u1_L2_reg_14 (.CK( clk ) , .Q( u1_L2_14 ) , .D( u1_R1_14 ) );
  DFF_X1 u1_L2_reg_15 (.CK( clk ) , .Q( u1_L2_15 ) , .D( u1_R1_15 ) );
  DFF_X1 u1_L2_reg_16 (.CK( clk ) , .Q( u1_L2_16 ) , .D( u1_R1_16 ) );
  DFF_X1 u1_L2_reg_17 (.CK( clk ) , .Q( u1_L2_17 ) , .D( u1_R1_17 ) );
  DFF_X1 u1_L2_reg_18 (.CK( clk ) , .Q( u1_L2_18 ) , .D( u1_R1_18 ) );
  DFF_X1 u1_L2_reg_19 (.CK( clk ) , .Q( u1_L2_19 ) , .D( u1_R1_19 ) );
  DFF_X1 u1_L2_reg_2 (.CK( clk ) , .Q( u1_L2_2 ) , .D( u1_R1_2 ) );
  DFF_X1 u1_L2_reg_20 (.CK( clk ) , .Q( u1_L2_20 ) , .D( u1_R1_20 ) );
  DFF_X1 u1_L2_reg_21 (.CK( clk ) , .Q( u1_L2_21 ) , .D( u1_R1_21 ) );
  DFF_X1 u1_L2_reg_22 (.CK( clk ) , .Q( u1_L2_22 ) , .D( u1_R1_22 ) );
  DFF_X1 u1_L2_reg_23 (.CK( clk ) , .Q( u1_L2_23 ) , .D( u1_R1_23 ) );
  DFF_X1 u1_L2_reg_24 (.CK( clk ) , .Q( u1_L2_24 ) , .D( u1_R1_24 ) );
  DFF_X1 u1_L2_reg_25 (.CK( clk ) , .Q( u1_L2_25 ) , .D( u1_R1_25 ) );
  DFF_X1 u1_L2_reg_26 (.CK( clk ) , .Q( u1_L2_26 ) , .D( u1_R1_26 ) );
  DFF_X1 u1_L2_reg_27 (.CK( clk ) , .Q( u1_L2_27 ) , .D( u1_R1_27 ) );
  DFF_X1 u1_L2_reg_28 (.CK( clk ) , .Q( u1_L2_28 ) , .D( u1_R1_28 ) );
  DFF_X1 u1_L2_reg_29 (.CK( clk ) , .Q( u1_L2_29 ) , .D( u1_R1_29 ) );
  DFF_X1 u1_L2_reg_3 (.CK( clk ) , .Q( u1_L2_3 ) , .D( u1_R1_3 ) );
  DFF_X1 u1_L2_reg_30 (.CK( clk ) , .Q( u1_L2_30 ) , .D( u1_R1_30 ) );
  DFF_X1 u1_L2_reg_31 (.CK( clk ) , .Q( u1_L2_31 ) , .D( u1_R1_31 ) );
  DFF_X1 u1_L2_reg_32 (.CK( clk ) , .Q( u1_L2_32 ) , .D( u1_R1_32 ) );
  DFF_X1 u1_L2_reg_4 (.CK( clk ) , .Q( u1_L2_4 ) , .D( u1_R1_4 ) );
  DFF_X1 u1_L2_reg_5 (.CK( clk ) , .Q( u1_L2_5 ) , .D( u1_R1_5 ) );
  DFF_X1 u1_L2_reg_6 (.CK( clk ) , .Q( u1_L2_6 ) , .D( u1_R1_6 ) );
  DFF_X1 u1_L2_reg_7 (.CK( clk ) , .Q( u1_L2_7 ) , .D( u1_R1_7 ) );
  DFF_X1 u1_L2_reg_8 (.CK( clk ) , .Q( u1_L2_8 ) , .D( u1_R1_8 ) );
  DFF_X1 u1_L2_reg_9 (.CK( clk ) , .Q( u1_L2_9 ) , .D( u1_R1_9 ) );
  DFF_X1 u1_L3_reg_1 (.CK( clk ) , .Q( u1_L3_1 ) , .D( u1_R2_1 ) );
  DFF_X1 u1_L3_reg_10 (.CK( clk ) , .Q( u1_L3_10 ) , .D( u1_R2_10 ) );
  DFF_X1 u1_L3_reg_11 (.CK( clk ) , .Q( u1_L3_11 ) , .D( u1_R2_11 ) );
  DFF_X1 u1_L3_reg_12 (.CK( clk ) , .Q( u1_L3_12 ) , .D( u1_R2_12 ) );
  DFF_X1 u1_L3_reg_13 (.CK( clk ) , .Q( u1_L3_13 ) , .D( u1_R2_13 ) );
  DFF_X1 u1_L3_reg_14 (.CK( clk ) , .Q( u1_L3_14 ) , .D( u1_R2_14 ) );
  DFF_X1 u1_L3_reg_15 (.CK( clk ) , .Q( u1_L3_15 ) , .D( u1_R2_15 ) );
  DFF_X1 u1_L3_reg_16 (.CK( clk ) , .Q( u1_L3_16 ) , .D( u1_R2_16 ) );
  DFF_X1 u1_L3_reg_17 (.CK( clk ) , .Q( u1_L3_17 ) , .D( u1_R2_17 ) );
  DFF_X1 u1_L3_reg_18 (.CK( clk ) , .Q( u1_L3_18 ) , .D( u1_R2_18 ) );
  DFF_X1 u1_L3_reg_19 (.CK( clk ) , .Q( u1_L3_19 ) , .D( u1_R2_19 ) );
  DFF_X1 u1_L3_reg_2 (.CK( clk ) , .Q( u1_L3_2 ) , .D( u1_R2_2 ) );
  DFF_X1 u1_L3_reg_20 (.CK( clk ) , .Q( u1_L3_20 ) , .D( u1_R2_20 ) );
  DFF_X1 u1_L3_reg_21 (.CK( clk ) , .Q( u1_L3_21 ) , .D( u1_R2_21 ) );
  DFF_X1 u1_L3_reg_22 (.CK( clk ) , .Q( u1_L3_22 ) , .D( u1_R2_22 ) );
  DFF_X1 u1_L3_reg_23 (.CK( clk ) , .Q( u1_L3_23 ) , .D( u1_R2_23 ) );
  DFF_X1 u1_L3_reg_24 (.CK( clk ) , .Q( u1_L3_24 ) , .D( u1_R2_24 ) );
  DFF_X1 u1_L3_reg_25 (.CK( clk ) , .Q( u1_L3_25 ) , .D( u1_R2_25 ) );
  DFF_X1 u1_L3_reg_26 (.CK( clk ) , .Q( u1_L3_26 ) , .D( u1_R2_26 ) );
  DFF_X1 u1_L3_reg_27 (.CK( clk ) , .Q( u1_L3_27 ) , .D( u1_R2_27 ) );
  DFF_X1 u1_L3_reg_28 (.CK( clk ) , .Q( u1_L3_28 ) , .D( u1_R2_28 ) );
  DFF_X1 u1_L3_reg_29 (.CK( clk ) , .Q( u1_L3_29 ) , .D( u1_R2_29 ) );
  DFF_X1 u1_L3_reg_3 (.CK( clk ) , .Q( u1_L3_3 ) , .D( u1_R2_3 ) );
  DFF_X1 u1_L3_reg_30 (.CK( clk ) , .Q( u1_L3_30 ) , .D( u1_R2_30 ) );
  DFF_X1 u1_L3_reg_31 (.CK( clk ) , .Q( u1_L3_31 ) , .D( u1_R2_31 ) );
  DFF_X1 u1_L3_reg_32 (.CK( clk ) , .Q( u1_L3_32 ) , .D( u1_R2_32 ) );
  DFF_X1 u1_L3_reg_4 (.CK( clk ) , .Q( u1_L3_4 ) , .D( u1_R2_4 ) );
  DFF_X1 u1_L3_reg_5 (.CK( clk ) , .Q( u1_L3_5 ) , .D( u1_R2_5 ) );
  DFF_X1 u1_L3_reg_6 (.CK( clk ) , .Q( u1_L3_6 ) , .D( u1_R2_6 ) );
  DFF_X1 u1_L3_reg_7 (.CK( clk ) , .Q( u1_L3_7 ) , .D( u1_R2_7 ) );
  DFF_X1 u1_L3_reg_8 (.CK( clk ) , .Q( u1_L3_8 ) , .D( u1_R2_8 ) );
  DFF_X1 u1_L3_reg_9 (.CK( clk ) , .Q( u1_L3_9 ) , .D( u1_R2_9 ) );
  DFF_X1 u1_L4_reg_1 (.CK( clk ) , .Q( u1_L4_1 ) , .D( u1_R3_1 ) );
  DFF_X1 u1_L4_reg_10 (.CK( clk ) , .Q( u1_L4_10 ) , .D( u1_R3_10 ) );
  DFF_X1 u1_L4_reg_11 (.CK( clk ) , .Q( u1_L4_11 ) , .D( u1_R3_11 ) );
  DFF_X1 u1_L4_reg_12 (.CK( clk ) , .Q( u1_L4_12 ) , .D( u1_R3_12 ) );
  DFF_X1 u1_L4_reg_13 (.CK( clk ) , .Q( u1_L4_13 ) , .D( u1_R3_13 ) );
  DFF_X1 u1_L4_reg_14 (.CK( clk ) , .Q( u1_L4_14 ) , .D( u1_R3_14 ) );
  DFF_X1 u1_L4_reg_15 (.CK( clk ) , .Q( u1_L4_15 ) , .D( u1_R3_15 ) );
  DFF_X1 u1_L4_reg_16 (.CK( clk ) , .Q( u1_L4_16 ) , .D( u1_R3_16 ) );
  DFF_X1 u1_L4_reg_17 (.CK( clk ) , .Q( u1_L4_17 ) , .D( u1_R3_17 ) );
  DFF_X1 u1_L4_reg_18 (.CK( clk ) , .Q( u1_L4_18 ) , .D( u1_R3_18 ) );
  DFF_X1 u1_L4_reg_19 (.CK( clk ) , .Q( u1_L4_19 ) , .D( u1_R3_19 ) );
  DFF_X1 u1_L4_reg_2 (.CK( clk ) , .Q( u1_L4_2 ) , .D( u1_R3_2 ) );
  DFF_X1 u1_L4_reg_20 (.CK( clk ) , .Q( u1_L4_20 ) , .D( u1_R3_20 ) );
  DFF_X1 u1_L4_reg_21 (.CK( clk ) , .Q( u1_L4_21 ) , .D( u1_R3_21 ) );
  DFF_X1 u1_L4_reg_22 (.CK( clk ) , .Q( u1_L4_22 ) , .D( u1_R3_22 ) );
  DFF_X1 u1_L4_reg_23 (.CK( clk ) , .Q( u1_L4_23 ) , .D( u1_R3_23 ) );
  DFF_X1 u1_L4_reg_24 (.CK( clk ) , .Q( u1_L4_24 ) , .D( u1_R3_24 ) );
  DFF_X1 u1_L4_reg_25 (.CK( clk ) , .Q( u1_L4_25 ) , .D( u1_R3_25 ) );
  DFF_X1 u1_L4_reg_26 (.CK( clk ) , .Q( u1_L4_26 ) , .D( u1_R3_26 ) );
  DFF_X1 u1_L4_reg_27 (.CK( clk ) , .Q( u1_L4_27 ) , .D( u1_R3_27 ) );
  DFF_X1 u1_L4_reg_28 (.CK( clk ) , .Q( u1_L4_28 ) , .D( u1_R3_28 ) );
  DFF_X1 u1_L4_reg_29 (.CK( clk ) , .Q( u1_L4_29 ) , .D( u1_R3_29 ) );
  DFF_X1 u1_L4_reg_3 (.CK( clk ) , .Q( u1_L4_3 ) , .D( u1_R3_3 ) );
  DFF_X1 u1_L4_reg_30 (.CK( clk ) , .Q( u1_L4_30 ) , .D( u1_R3_30 ) );
  DFF_X1 u1_L4_reg_31 (.CK( clk ) , .Q( u1_L4_31 ) , .D( u1_R3_31 ) );
  DFF_X1 u1_L4_reg_32 (.CK( clk ) , .Q( u1_L4_32 ) , .D( u1_R3_32 ) );
  DFF_X1 u1_L4_reg_4 (.CK( clk ) , .Q( u1_L4_4 ) , .D( u1_R3_4 ) );
  DFF_X1 u1_L4_reg_5 (.CK( clk ) , .Q( u1_L4_5 ) , .D( u1_R3_5 ) );
  DFF_X1 u1_L4_reg_6 (.CK( clk ) , .Q( u1_L4_6 ) , .D( u1_R3_6 ) );
  DFF_X1 u1_L4_reg_7 (.CK( clk ) , .Q( u1_L4_7 ) , .D( u1_R3_7 ) );
  DFF_X1 u1_L4_reg_8 (.CK( clk ) , .Q( u1_L4_8 ) , .D( u1_R3_8 ) );
  DFF_X1 u1_L4_reg_9 (.CK( clk ) , .Q( u1_L4_9 ) , .D( u1_R3_9 ) );
  DFF_X1 u1_L5_reg_1 (.CK( clk ) , .Q( u1_L5_1 ) , .D( u1_R4_1 ) );
  DFF_X1 u1_L5_reg_10 (.CK( clk ) , .Q( u1_L5_10 ) , .D( u1_R4_10 ) );
  DFF_X1 u1_L5_reg_11 (.CK( clk ) , .Q( u1_L5_11 ) , .D( u1_R4_11 ) );
  DFF_X1 u1_L5_reg_12 (.CK( clk ) , .Q( u1_L5_12 ) , .D( u1_R4_12 ) );
  DFF_X1 u1_L5_reg_13 (.CK( clk ) , .Q( u1_L5_13 ) , .D( u1_R4_13 ) );
  DFF_X1 u1_L5_reg_14 (.CK( clk ) , .Q( u1_L5_14 ) , .D( u1_R4_14 ) );
  DFF_X1 u1_L5_reg_15 (.CK( clk ) , .Q( u1_L5_15 ) , .D( u1_R4_15 ) );
  DFF_X1 u1_L5_reg_16 (.CK( clk ) , .Q( u1_L5_16 ) , .D( u1_R4_16 ) );
  DFF_X1 u1_L5_reg_17 (.CK( clk ) , .Q( u1_L5_17 ) , .D( u1_R4_17 ) );
  DFF_X1 u1_L5_reg_18 (.CK( clk ) , .Q( u1_L5_18 ) , .D( u1_R4_18 ) );
  DFF_X1 u1_L5_reg_19 (.CK( clk ) , .Q( u1_L5_19 ) , .D( u1_R4_19 ) );
  DFF_X1 u1_L5_reg_2 (.CK( clk ) , .Q( u1_L5_2 ) , .D( u1_R4_2 ) );
  DFF_X1 u1_L5_reg_20 (.CK( clk ) , .Q( u1_L5_20 ) , .D( u1_R4_20 ) );
  DFF_X1 u1_L5_reg_21 (.CK( clk ) , .Q( u1_L5_21 ) , .D( u1_R4_21 ) );
  DFF_X1 u1_L5_reg_22 (.CK( clk ) , .Q( u1_L5_22 ) , .D( u1_R4_22 ) );
  DFF_X1 u1_L5_reg_23 (.CK( clk ) , .Q( u1_L5_23 ) , .D( u1_R4_23 ) );
  DFF_X1 u1_L5_reg_24 (.CK( clk ) , .Q( u1_L5_24 ) , .D( u1_R4_24 ) );
  DFF_X1 u1_L5_reg_25 (.CK( clk ) , .Q( u1_L5_25 ) , .D( u1_R4_25 ) );
  DFF_X1 u1_L5_reg_26 (.CK( clk ) , .Q( u1_L5_26 ) , .D( u1_R4_26 ) );
  DFF_X1 u1_L5_reg_27 (.CK( clk ) , .Q( u1_L5_27 ) , .D( u1_R4_27 ) );
  DFF_X1 u1_L5_reg_28 (.CK( clk ) , .Q( u1_L5_28 ) , .D( u1_R4_28 ) );
  DFF_X1 u1_L5_reg_29 (.CK( clk ) , .Q( u1_L5_29 ) , .D( u1_R4_29 ) );
  DFF_X1 u1_L5_reg_3 (.CK( clk ) , .Q( u1_L5_3 ) , .D( u1_R4_3 ) );
  DFF_X1 u1_L5_reg_30 (.CK( clk ) , .Q( u1_L5_30 ) , .D( u1_R4_30 ) );
  DFF_X1 u1_L5_reg_31 (.CK( clk ) , .Q( u1_L5_31 ) , .D( u1_R4_31 ) );
  DFF_X1 u1_L5_reg_32 (.CK( clk ) , .Q( u1_L5_32 ) , .D( u1_R4_32 ) );
  DFF_X1 u1_L5_reg_4 (.CK( clk ) , .Q( u1_L5_4 ) , .D( u1_R4_4 ) );
  DFF_X1 u1_L5_reg_5 (.CK( clk ) , .Q( u1_L5_5 ) , .D( u1_R4_5 ) );
  DFF_X1 u1_L5_reg_6 (.CK( clk ) , .Q( u1_L5_6 ) , .D( u1_R4_6 ) );
  DFF_X1 u1_L5_reg_7 (.CK( clk ) , .Q( u1_L5_7 ) , .D( u1_R4_7 ) );
  DFF_X1 u1_L5_reg_8 (.CK( clk ) , .Q( u1_L5_8 ) , .D( u1_R4_8 ) );
  DFF_X1 u1_L5_reg_9 (.CK( clk ) , .Q( u1_L5_9 ) , .D( u1_R4_9 ) );
  DFF_X1 u1_L6_reg_1 (.CK( clk ) , .Q( u1_L6_1 ) , .D( u1_R5_1 ) );
  DFF_X1 u1_L6_reg_10 (.CK( clk ) , .Q( u1_L6_10 ) , .D( u1_R5_10 ) );
  DFF_X1 u1_L6_reg_11 (.CK( clk ) , .Q( u1_L6_11 ) , .D( u1_R5_11 ) );
  DFF_X1 u1_L6_reg_12 (.CK( clk ) , .Q( u1_L6_12 ) , .D( u1_R5_12 ) );
  DFF_X1 u1_L6_reg_13 (.CK( clk ) , .Q( u1_L6_13 ) , .D( u1_R5_13 ) );
  DFF_X1 u1_L6_reg_14 (.CK( clk ) , .Q( u1_L6_14 ) , .D( u1_R5_14 ) );
  DFF_X1 u1_L6_reg_15 (.CK( clk ) , .Q( u1_L6_15 ) , .D( u1_R5_15 ) );
  DFF_X1 u1_L6_reg_16 (.CK( clk ) , .Q( u1_L6_16 ) , .D( u1_R5_16 ) );
  DFF_X1 u1_L6_reg_17 (.CK( clk ) , .Q( u1_L6_17 ) , .D( u1_R5_17 ) );
  DFF_X1 u1_L6_reg_18 (.CK( clk ) , .Q( u1_L6_18 ) , .D( u1_R5_18 ) );
  DFF_X1 u1_L6_reg_19 (.CK( clk ) , .Q( u1_L6_19 ) , .D( u1_R5_19 ) );
  DFF_X1 u1_L6_reg_2 (.CK( clk ) , .Q( u1_L6_2 ) , .D( u1_R5_2 ) );
  DFF_X1 u1_L6_reg_20 (.CK( clk ) , .Q( u1_L6_20 ) , .D( u1_R5_20 ) );
  DFF_X1 u1_L6_reg_21 (.CK( clk ) , .Q( u1_L6_21 ) , .D( u1_R5_21 ) );
  DFF_X1 u1_L6_reg_22 (.CK( clk ) , .Q( u1_L6_22 ) , .D( u1_R5_22 ) );
  DFF_X1 u1_L6_reg_23 (.CK( clk ) , .Q( u1_L6_23 ) , .D( u1_R5_23 ) );
  DFF_X1 u1_L6_reg_24 (.CK( clk ) , .Q( u1_L6_24 ) , .D( u1_R5_24 ) );
  DFF_X1 u1_L6_reg_25 (.CK( clk ) , .Q( u1_L6_25 ) , .D( u1_R5_25 ) );
  DFF_X1 u1_L6_reg_26 (.CK( clk ) , .Q( u1_L6_26 ) , .D( u1_R5_26 ) );
  DFF_X1 u1_L6_reg_27 (.CK( clk ) , .Q( u1_L6_27 ) , .D( u1_R5_27 ) );
  DFF_X1 u1_L6_reg_28 (.CK( clk ) , .Q( u1_L6_28 ) , .D( u1_R5_28 ) );
  DFF_X1 u1_L6_reg_29 (.CK( clk ) , .Q( u1_L6_29 ) , .D( u1_R5_29 ) );
  DFF_X1 u1_L6_reg_3 (.CK( clk ) , .Q( u1_L6_3 ) , .D( u1_R5_3 ) );
  DFF_X1 u1_L6_reg_30 (.CK( clk ) , .Q( u1_L6_30 ) , .D( u1_R5_30 ) );
  DFF_X1 u1_L6_reg_31 (.CK( clk ) , .Q( u1_L6_31 ) , .D( u1_R5_31 ) );
  DFF_X1 u1_L6_reg_32 (.CK( clk ) , .Q( u1_L6_32 ) , .D( u1_R5_32 ) );
  DFF_X1 u1_L6_reg_4 (.CK( clk ) , .Q( u1_L6_4 ) , .D( u1_R5_4 ) );
  DFF_X1 u1_L6_reg_5 (.CK( clk ) , .Q( u1_L6_5 ) , .D( u1_R5_5 ) );
  DFF_X1 u1_L6_reg_6 (.CK( clk ) , .Q( u1_L6_6 ) , .D( u1_R5_6 ) );
  DFF_X1 u1_L6_reg_7 (.CK( clk ) , .Q( u1_L6_7 ) , .D( u1_R5_7 ) );
  DFF_X1 u1_L6_reg_8 (.CK( clk ) , .Q( u1_L6_8 ) , .D( u1_R5_8 ) );
  DFF_X1 u1_L6_reg_9 (.CK( clk ) , .Q( u1_L6_9 ) , .D( u1_R5_9 ) );
  DFF_X1 u1_L7_reg_1 (.CK( clk ) , .Q( u1_L7_1 ) , .D( u1_R6_1 ) );
  DFF_X1 u1_L7_reg_10 (.CK( clk ) , .Q( u1_L7_10 ) , .D( u1_R6_10 ) );
  DFF_X1 u1_L7_reg_11 (.CK( clk ) , .Q( u1_L7_11 ) , .D( u1_R6_11 ) );
  DFF_X1 u1_L7_reg_12 (.CK( clk ) , .Q( u1_L7_12 ) , .D( u1_R6_12 ) );
  DFF_X1 u1_L7_reg_13 (.CK( clk ) , .Q( u1_L7_13 ) , .D( u1_R6_13 ) );
  DFF_X1 u1_L7_reg_14 (.CK( clk ) , .Q( u1_L7_14 ) , .D( u1_R6_14 ) );
  DFF_X1 u1_L7_reg_15 (.CK( clk ) , .Q( u1_L7_15 ) , .D( u1_R6_15 ) );
  DFF_X1 u1_L7_reg_16 (.CK( clk ) , .Q( u1_L7_16 ) , .D( u1_R6_16 ) );
  DFF_X1 u1_L7_reg_17 (.CK( clk ) , .Q( u1_L7_17 ) , .D( u1_R6_17 ) );
  DFF_X1 u1_L7_reg_18 (.CK( clk ) , .Q( u1_L7_18 ) , .D( u1_R6_18 ) );
  DFF_X1 u1_L7_reg_19 (.CK( clk ) , .Q( u1_L7_19 ) , .D( u1_R6_19 ) );
  DFF_X1 u1_L7_reg_2 (.CK( clk ) , .Q( u1_L7_2 ) , .D( u1_R6_2 ) );
  DFF_X1 u1_L7_reg_20 (.CK( clk ) , .Q( u1_L7_20 ) , .D( u1_R6_20 ) );
  DFF_X1 u1_L7_reg_21 (.CK( clk ) , .Q( u1_L7_21 ) , .D( u1_R6_21 ) );
  DFF_X1 u1_L7_reg_22 (.CK( clk ) , .Q( u1_L7_22 ) , .D( u1_R6_22 ) );
  DFF_X1 u1_L7_reg_23 (.CK( clk ) , .Q( u1_L7_23 ) , .D( u1_R6_23 ) );
  DFF_X1 u1_L7_reg_24 (.CK( clk ) , .Q( u1_L7_24 ) , .D( u1_R6_24 ) );
  DFF_X1 u1_L7_reg_25 (.CK( clk ) , .Q( u1_L7_25 ) , .D( u1_R6_25 ) );
  DFF_X1 u1_L7_reg_26 (.CK( clk ) , .Q( u1_L7_26 ) , .D( u1_R6_26 ) );
  DFF_X1 u1_L7_reg_27 (.CK( clk ) , .Q( u1_L7_27 ) , .D( u1_R6_27 ) );
  DFF_X1 u1_L7_reg_28 (.CK( clk ) , .Q( u1_L7_28 ) , .D( u1_R6_28 ) );
  DFF_X1 u1_L7_reg_29 (.CK( clk ) , .Q( u1_L7_29 ) , .D( u1_R6_29 ) );
  DFF_X1 u1_L7_reg_3 (.CK( clk ) , .Q( u1_L7_3 ) , .D( u1_R6_3 ) );
  DFF_X1 u1_L7_reg_30 (.CK( clk ) , .Q( u1_L7_30 ) , .D( u1_R6_30 ) );
  DFF_X1 u1_L7_reg_31 (.CK( clk ) , .Q( u1_L7_31 ) , .D( u1_R6_31 ) );
  DFF_X1 u1_L7_reg_32 (.CK( clk ) , .Q( u1_L7_32 ) , .D( u1_R6_32 ) );
  DFF_X1 u1_L7_reg_4 (.CK( clk ) , .Q( u1_L7_4 ) , .D( u1_R6_4 ) );
  DFF_X1 u1_L7_reg_5 (.CK( clk ) , .Q( u1_L7_5 ) , .D( u1_R6_5 ) );
  DFF_X1 u1_L7_reg_6 (.CK( clk ) , .Q( u1_L7_6 ) , .D( u1_R6_6 ) );
  DFF_X1 u1_L7_reg_7 (.CK( clk ) , .Q( u1_L7_7 ) , .D( u1_R6_7 ) );
  DFF_X1 u1_L7_reg_8 (.CK( clk ) , .Q( u1_L7_8 ) , .D( u1_R6_8 ) );
  DFF_X1 u1_L7_reg_9 (.CK( clk ) , .Q( u1_L7_9 ) , .D( u1_R6_9 ) );
  DFF_X1 u1_L8_reg_1 (.CK( clk ) , .Q( u1_L8_1 ) , .D( u1_R7_1 ) );
  DFF_X1 u1_L8_reg_10 (.CK( clk ) , .Q( u1_L8_10 ) , .D( u1_R7_10 ) );
  DFF_X1 u1_L8_reg_11 (.CK( clk ) , .Q( u1_L8_11 ) , .D( u1_R7_11 ) );
  DFF_X1 u1_L8_reg_12 (.CK( clk ) , .Q( u1_L8_12 ) , .D( u1_R7_12 ) );
  DFF_X1 u1_L8_reg_13 (.CK( clk ) , .Q( u1_L8_13 ) , .D( u1_R7_13 ) );
  DFF_X1 u1_L8_reg_14 (.CK( clk ) , .Q( u1_L8_14 ) , .D( u1_R7_14 ) );
  DFF_X1 u1_L8_reg_15 (.CK( clk ) , .Q( u1_L8_15 ) , .D( u1_R7_15 ) );
  DFF_X1 u1_L8_reg_16 (.CK( clk ) , .Q( u1_L8_16 ) , .D( u1_R7_16 ) );
  DFF_X1 u1_L8_reg_17 (.CK( clk ) , .Q( u1_L8_17 ) , .D( u1_R7_17 ) );
  DFF_X1 u1_L8_reg_18 (.CK( clk ) , .Q( u1_L8_18 ) , .D( u1_R7_18 ) );
  DFF_X1 u1_L8_reg_19 (.CK( clk ) , .Q( u1_L8_19 ) , .D( u1_R7_19 ) );
  DFF_X1 u1_L8_reg_2 (.CK( clk ) , .Q( u1_L8_2 ) , .D( u1_R7_2 ) );
  DFF_X1 u1_L8_reg_20 (.CK( clk ) , .Q( u1_L8_20 ) , .D( u1_R7_20 ) );
  DFF_X1 u1_L8_reg_21 (.CK( clk ) , .Q( u1_L8_21 ) , .D( u1_R7_21 ) );
  DFF_X1 u1_L8_reg_22 (.CK( clk ) , .Q( u1_L8_22 ) , .D( u1_R7_22 ) );
  DFF_X1 u1_L8_reg_23 (.CK( clk ) , .Q( u1_L8_23 ) , .D( u1_R7_23 ) );
  DFF_X1 u1_L8_reg_24 (.CK( clk ) , .Q( u1_L8_24 ) , .D( u1_R7_24 ) );
  DFF_X1 u1_L8_reg_25 (.CK( clk ) , .Q( u1_L8_25 ) , .D( u1_R7_25 ) );
  DFF_X1 u1_L8_reg_26 (.CK( clk ) , .Q( u1_L8_26 ) , .D( u1_R7_26 ) );
  DFF_X1 u1_L8_reg_27 (.CK( clk ) , .Q( u1_L8_27 ) , .D( u1_R7_27 ) );
  DFF_X1 u1_L8_reg_28 (.CK( clk ) , .Q( u1_L8_28 ) , .D( u1_R7_28 ) );
  DFF_X1 u1_L8_reg_29 (.CK( clk ) , .Q( u1_L8_29 ) , .D( u1_R7_29 ) );
  DFF_X1 u1_L8_reg_3 (.CK( clk ) , .Q( u1_L8_3 ) , .D( u1_R7_3 ) );
  DFF_X1 u1_L8_reg_30 (.CK( clk ) , .Q( u1_L8_30 ) , .D( u1_R7_30 ) );
  DFF_X1 u1_L8_reg_31 (.CK( clk ) , .Q( u1_L8_31 ) , .D( u1_R7_31 ) );
  DFF_X1 u1_L8_reg_32 (.CK( clk ) , .Q( u1_L8_32 ) , .D( u1_R7_32 ) );
  DFF_X1 u1_L8_reg_4 (.CK( clk ) , .Q( u1_L8_4 ) , .D( u1_R7_4 ) );
  DFF_X1 u1_L8_reg_5 (.CK( clk ) , .Q( u1_L8_5 ) , .D( u1_R7_5 ) );
  DFF_X1 u1_L8_reg_6 (.CK( clk ) , .Q( u1_L8_6 ) , .D( u1_R7_6 ) );
  DFF_X1 u1_L8_reg_7 (.CK( clk ) , .Q( u1_L8_7 ) , .D( u1_R7_7 ) );
  DFF_X1 u1_L8_reg_8 (.CK( clk ) , .Q( u1_L8_8 ) , .D( u1_R7_8 ) );
  DFF_X1 u1_L8_reg_9 (.CK( clk ) , .Q( u1_L8_9 ) , .D( u1_R7_9 ) );
  DFF_X1 u1_L9_reg_1 (.CK( clk ) , .Q( u1_L9_1 ) , .D( u1_R8_1 ) );
  DFF_X1 u1_L9_reg_10 (.CK( clk ) , .Q( u1_L9_10 ) , .D( u1_R8_10 ) );
  DFF_X1 u1_L9_reg_11 (.CK( clk ) , .Q( u1_L9_11 ) , .D( u1_R8_11 ) );
  DFF_X1 u1_L9_reg_12 (.CK( clk ) , .Q( u1_L9_12 ) , .D( u1_R8_12 ) );
  DFF_X1 u1_L9_reg_13 (.CK( clk ) , .Q( u1_L9_13 ) , .D( u1_R8_13 ) );
  DFF_X1 u1_L9_reg_14 (.CK( clk ) , .Q( u1_L9_14 ) , .D( u1_R8_14 ) );
  DFF_X1 u1_L9_reg_15 (.CK( clk ) , .Q( u1_L9_15 ) , .D( u1_R8_15 ) );
  DFF_X1 u1_L9_reg_16 (.CK( clk ) , .Q( u1_L9_16 ) , .D( u1_R8_16 ) );
  DFF_X1 u1_L9_reg_17 (.CK( clk ) , .Q( u1_L9_17 ) , .D( u1_R8_17 ) );
  DFF_X1 u1_L9_reg_18 (.CK( clk ) , .Q( u1_L9_18 ) , .D( u1_R8_18 ) );
  DFF_X1 u1_L9_reg_19 (.CK( clk ) , .Q( u1_L9_19 ) , .D( u1_R8_19 ) );
  DFF_X1 u1_L9_reg_2 (.CK( clk ) , .Q( u1_L9_2 ) , .D( u1_R8_2 ) );
  DFF_X1 u1_L9_reg_20 (.CK( clk ) , .Q( u1_L9_20 ) , .D( u1_R8_20 ) );
  DFF_X1 u1_L9_reg_21 (.CK( clk ) , .Q( u1_L9_21 ) , .D( u1_R8_21 ) );
  DFF_X1 u1_L9_reg_22 (.CK( clk ) , .Q( u1_L9_22 ) , .D( u1_R8_22 ) );
  DFF_X1 u1_L9_reg_23 (.CK( clk ) , .Q( u1_L9_23 ) , .D( u1_R8_23 ) );
  DFF_X1 u1_L9_reg_24 (.CK( clk ) , .Q( u1_L9_24 ) , .D( u1_R8_24 ) );
  DFF_X1 u1_L9_reg_25 (.CK( clk ) , .Q( u1_L9_25 ) , .D( u1_R8_25 ) );
  DFF_X1 u1_L9_reg_26 (.CK( clk ) , .Q( u1_L9_26 ) , .D( u1_R8_26 ) );
  DFF_X1 u1_L9_reg_27 (.CK( clk ) , .Q( u1_L9_27 ) , .D( u1_R8_27 ) );
  DFF_X1 u1_L9_reg_28 (.CK( clk ) , .Q( u1_L9_28 ) , .D( u1_R8_28 ) );
  DFF_X1 u1_L9_reg_29 (.CK( clk ) , .Q( u1_L9_29 ) , .D( u1_R8_29 ) );
  DFF_X1 u1_L9_reg_3 (.CK( clk ) , .Q( u1_L9_3 ) , .D( u1_R8_3 ) );
  DFF_X1 u1_L9_reg_30 (.CK( clk ) , .Q( u1_L9_30 ) , .D( u1_R8_30 ) );
  DFF_X1 u1_L9_reg_31 (.CK( clk ) , .Q( u1_L9_31 ) , .D( u1_R8_31 ) );
  DFF_X1 u1_L9_reg_32 (.CK( clk ) , .Q( u1_L9_32 ) , .D( u1_R8_32 ) );
  DFF_X1 u1_L9_reg_4 (.CK( clk ) , .Q( u1_L9_4 ) , .D( u1_R8_4 ) );
  DFF_X1 u1_L9_reg_5 (.CK( clk ) , .Q( u1_L9_5 ) , .D( u1_R8_5 ) );
  DFF_X1 u1_L9_reg_6 (.CK( clk ) , .Q( u1_L9_6 ) , .D( u1_R8_6 ) );
  DFF_X1 u1_L9_reg_7 (.CK( clk ) , .Q( u1_L9_7 ) , .D( u1_R8_7 ) );
  DFF_X1 u1_L9_reg_8 (.CK( clk ) , .Q( u1_L9_8 ) , .D( u1_R8_8 ) );
  DFF_X1 u1_L9_reg_9 (.CK( clk ) , .Q( u1_L9_9 ) , .D( u1_R8_9 ) );
  DFF_X1 u1_R0_reg_1 (.CK( clk ) , .D( u1_N0 ) , .Q( u1_R0_1 ) );
  DFF_X1 u1_R0_reg_10 (.CK( clk ) , .D( u1_N9 ) , .Q( u1_R0_10 ) );
  DFF_X1 u1_R0_reg_11 (.CK( clk ) , .D( u1_N10 ) , .Q( u1_R0_11 ) );
  DFF_X1 u1_R0_reg_12 (.CK( clk ) , .D( u1_N11 ) , .Q( u1_R0_12 ) );
  DFF_X1 u1_R0_reg_13 (.CK( clk ) , .D( u1_N12 ) , .Q( u1_R0_13 ) );
  DFF_X1 u1_R0_reg_14 (.CK( clk ) , .D( u1_N13 ) , .Q( u1_R0_14 ) );
  DFF_X1 u1_R0_reg_15 (.CK( clk ) , .D( u1_N14 ) , .Q( u1_R0_15 ) );
  DFF_X1 u1_R0_reg_16 (.CK( clk ) , .D( u1_N15 ) , .Q( u1_R0_16 ) );
  DFF_X1 u1_R0_reg_17 (.CK( clk ) , .D( u1_N16 ) , .Q( u1_R0_17 ) );
  DFF_X1 u1_R0_reg_18 (.CK( clk ) , .D( u1_N17 ) , .Q( u1_R0_18 ) );
  DFF_X1 u1_R0_reg_19 (.CK( clk ) , .D( u1_N18 ) , .Q( u1_R0_19 ) );
  DFF_X1 u1_R0_reg_2 (.CK( clk ) , .D( u1_N1 ) , .Q( u1_R0_2 ) );
  DFF_X1 u1_R0_reg_20 (.CK( clk ) , .D( u1_N19 ) , .Q( u1_R0_20 ) );
  DFF_X1 u1_R0_reg_21 (.CK( clk ) , .D( u1_N20 ) , .Q( u1_R0_21 ) );
  DFF_X1 u1_R0_reg_22 (.CK( clk ) , .D( u1_N21 ) , .Q( u1_R0_22 ) );
  DFF_X1 u1_R0_reg_23 (.CK( clk ) , .D( u1_N22 ) , .Q( u1_R0_23 ) );
  DFF_X1 u1_R0_reg_24 (.CK( clk ) , .D( u1_N23 ) , .Q( u1_R0_24 ) );
  DFF_X1 u1_R0_reg_25 (.CK( clk ) , .D( u1_N24 ) , .Q( u1_R0_25 ) );
  DFF_X1 u1_R0_reg_26 (.CK( clk ) , .D( u1_N25 ) , .Q( u1_R0_26 ) );
  DFF_X1 u1_R0_reg_27 (.CK( clk ) , .D( u1_N26 ) , .Q( u1_R0_27 ) );
  DFF_X1 u1_R0_reg_28 (.CK( clk ) , .D( u1_N27 ) , .Q( u1_R0_28 ) );
  DFF_X1 u1_R0_reg_29 (.CK( clk ) , .D( u1_N28 ) , .Q( u1_R0_29 ) );
  DFF_X1 u1_R0_reg_3 (.CK( clk ) , .D( u1_N2 ) , .Q( u1_R0_3 ) );
  DFF_X1 u1_R0_reg_30 (.CK( clk ) , .D( u1_N29 ) , .Q( u1_R0_30 ) );
  DFF_X1 u1_R0_reg_31 (.CK( clk ) , .D( u1_N30 ) , .Q( u1_R0_31 ) );
  DFF_X1 u1_R0_reg_32 (.CK( clk ) , .D( u1_N31 ) , .Q( u1_R0_32 ) );
  DFF_X1 u1_R0_reg_4 (.CK( clk ) , .D( u1_N3 ) , .Q( u1_R0_4 ) );
  DFF_X1 u1_R0_reg_5 (.CK( clk ) , .D( u1_N4 ) , .Q( u1_R0_5 ) );
  DFF_X1 u1_R0_reg_6 (.CK( clk ) , .D( u1_N5 ) , .Q( u1_R0_6 ) );
  DFF_X1 u1_R0_reg_7 (.CK( clk ) , .D( u1_N6 ) , .Q( u1_R0_7 ) );
  DFF_X1 u1_R0_reg_8 (.CK( clk ) , .D( u1_N7 ) , .Q( u1_R0_8 ) );
  DFF_X1 u1_R0_reg_9 (.CK( clk ) , .D( u1_N8 ) , .Q( u1_R0_9 ) );
  DFF_X1 u1_R10_reg_1 (.CK( clk ) , .D( u1_N320 ) , .Q( u1_R10_1 ) );
  DFF_X1 u1_R10_reg_10 (.CK( clk ) , .D( u1_N329 ) , .Q( u1_R10_10 ) );
  DFF_X1 u1_R10_reg_11 (.CK( clk ) , .D( u1_N330 ) , .Q( u1_R10_11 ) );
  DFF_X1 u1_R10_reg_12 (.CK( clk ) , .D( u1_N331 ) , .Q( u1_R10_12 ) );
  DFF_X1 u1_R10_reg_13 (.CK( clk ) , .D( u1_N332 ) , .Q( u1_R10_13 ) );
  DFF_X1 u1_R10_reg_14 (.CK( clk ) , .D( u1_N333 ) , .Q( u1_R10_14 ) );
  DFF_X1 u1_R10_reg_15 (.CK( clk ) , .D( u1_N334 ) , .Q( u1_R10_15 ) );
  DFF_X1 u1_R10_reg_16 (.CK( clk ) , .D( u1_N335 ) , .Q( u1_R10_16 ) );
  DFF_X1 u1_R10_reg_17 (.CK( clk ) , .D( u1_N336 ) , .Q( u1_R10_17 ) );
  DFF_X1 u1_R10_reg_18 (.CK( clk ) , .D( u1_N337 ) , .Q( u1_R10_18 ) );
  DFF_X1 u1_R10_reg_19 (.CK( clk ) , .D( u1_N338 ) , .Q( u1_R10_19 ) );
  DFF_X1 u1_R10_reg_2 (.CK( clk ) , .D( u1_N321 ) , .Q( u1_R10_2 ) );
  DFF_X1 u1_R10_reg_20 (.CK( clk ) , .D( u1_N339 ) , .Q( u1_R10_20 ) );
  DFF_X1 u1_R10_reg_21 (.CK( clk ) , .D( u1_N340 ) , .Q( u1_R10_21 ) );
  DFF_X1 u1_R10_reg_22 (.CK( clk ) , .D( u1_N341 ) , .Q( u1_R10_22 ) );
  DFF_X1 u1_R10_reg_23 (.CK( clk ) , .D( u1_N342 ) , .Q( u1_R10_23 ) );
  DFF_X1 u1_R10_reg_24 (.CK( clk ) , .D( u1_N343 ) , .Q( u1_R10_24 ) );
  DFF_X1 u1_R10_reg_25 (.CK( clk ) , .D( u1_N344 ) , .Q( u1_R10_25 ) );
  DFF_X1 u1_R10_reg_26 (.CK( clk ) , .D( u1_N345 ) , .Q( u1_R10_26 ) );
  DFF_X1 u1_R10_reg_27 (.CK( clk ) , .D( u1_N346 ) , .Q( u1_R10_27 ) );
  DFF_X1 u1_R10_reg_28 (.CK( clk ) , .D( u1_N347 ) , .Q( u1_R10_28 ) );
  DFF_X1 u1_R10_reg_29 (.CK( clk ) , .D( u1_N348 ) , .Q( u1_R10_29 ) );
  DFF_X1 u1_R10_reg_3 (.CK( clk ) , .D( u1_N322 ) , .Q( u1_R10_3 ) );
  DFF_X1 u1_R10_reg_30 (.CK( clk ) , .D( u1_N349 ) , .Q( u1_R10_30 ) );
  DFF_X1 u1_R10_reg_31 (.CK( clk ) , .D( u1_N350 ) , .Q( u1_R10_31 ) );
  DFF_X1 u1_R10_reg_32 (.CK( clk ) , .D( u1_N351 ) , .Q( u1_R10_32 ) );
  DFF_X1 u1_R10_reg_4 (.CK( clk ) , .D( u1_N323 ) , .Q( u1_R10_4 ) );
  DFF_X1 u1_R10_reg_5 (.CK( clk ) , .D( u1_N324 ) , .Q( u1_R10_5 ) );
  DFF_X1 u1_R10_reg_6 (.CK( clk ) , .D( u1_N325 ) , .Q( u1_R10_6 ) );
  DFF_X1 u1_R10_reg_7 (.CK( clk ) , .D( u1_N326 ) , .Q( u1_R10_7 ) );
  DFF_X1 u1_R10_reg_8 (.CK( clk ) , .D( u1_N327 ) , .Q( u1_R10_8 ) );
  DFF_X1 u1_R10_reg_9 (.CK( clk ) , .D( u1_N328 ) , .Q( u1_R10_9 ) );
  DFF_X1 u1_R11_reg_1 (.CK( clk ) , .D( u1_N352 ) , .Q( u1_R11_1 ) );
  DFF_X1 u1_R11_reg_10 (.CK( clk ) , .D( u1_N361 ) , .Q( u1_R11_10 ) );
  DFF_X1 u1_R11_reg_11 (.CK( clk ) , .D( u1_N362 ) , .Q( u1_R11_11 ) );
  DFF_X1 u1_R11_reg_12 (.CK( clk ) , .D( u1_N363 ) , .Q( u1_R11_12 ) );
  DFF_X1 u1_R11_reg_13 (.CK( clk ) , .D( u1_N364 ) , .Q( u1_R11_13 ) );
  DFF_X1 u1_R11_reg_14 (.CK( clk ) , .D( u1_N365 ) , .Q( u1_R11_14 ) );
  DFF_X1 u1_R11_reg_15 (.CK( clk ) , .D( u1_N366 ) , .Q( u1_R11_15 ) );
  DFF_X1 u1_R11_reg_16 (.CK( clk ) , .D( u1_N367 ) , .Q( u1_R11_16 ) );
  DFF_X1 u1_R11_reg_17 (.CK( clk ) , .D( u1_N368 ) , .Q( u1_R11_17 ) );
  DFF_X1 u1_R11_reg_18 (.CK( clk ) , .D( u1_N369 ) , .Q( u1_R11_18 ) );
  DFF_X1 u1_R11_reg_19 (.CK( clk ) , .D( u1_N370 ) , .Q( u1_R11_19 ) );
  DFF_X1 u1_R11_reg_2 (.CK( clk ) , .D( u1_N353 ) , .Q( u1_R11_2 ) );
  DFF_X1 u1_R11_reg_20 (.CK( clk ) , .D( u1_N371 ) , .Q( u1_R11_20 ) );
  DFF_X1 u1_R11_reg_21 (.CK( clk ) , .D( u1_N372 ) , .Q( u1_R11_21 ) );
  DFF_X1 u1_R11_reg_22 (.CK( clk ) , .D( u1_N373 ) , .Q( u1_R11_22 ) );
  DFF_X1 u1_R11_reg_23 (.CK( clk ) , .D( u1_N374 ) , .Q( u1_R11_23 ) );
  DFF_X1 u1_R11_reg_24 (.CK( clk ) , .D( u1_N375 ) , .Q( u1_R11_24 ) );
  DFF_X1 u1_R11_reg_25 (.CK( clk ) , .D( u1_N376 ) , .Q( u1_R11_25 ) );
  DFF_X1 u1_R11_reg_26 (.CK( clk ) , .D( u1_N377 ) , .Q( u1_R11_26 ) );
  DFF_X1 u1_R11_reg_27 (.CK( clk ) , .D( u1_N378 ) , .Q( u1_R11_27 ) );
  DFF_X1 u1_R11_reg_28 (.CK( clk ) , .D( u1_N379 ) , .Q( u1_R11_28 ) );
  DFF_X1 u1_R11_reg_29 (.CK( clk ) , .D( u1_N380 ) , .Q( u1_R11_29 ) );
  DFF_X1 u1_R11_reg_3 (.CK( clk ) , .D( u1_N354 ) , .Q( u1_R11_3 ) );
  DFF_X1 u1_R11_reg_30 (.CK( clk ) , .D( u1_N381 ) , .Q( u1_R11_30 ) );
  DFF_X1 u1_R11_reg_31 (.CK( clk ) , .D( u1_N382 ) , .Q( u1_R11_31 ) );
  DFF_X1 u1_R11_reg_32 (.CK( clk ) , .D( u1_N383 ) , .Q( u1_R11_32 ) );
  DFF_X1 u1_R11_reg_4 (.CK( clk ) , .D( u1_N355 ) , .Q( u1_R11_4 ) );
  DFF_X1 u1_R11_reg_5 (.CK( clk ) , .D( u1_N356 ) , .Q( u1_R11_5 ) );
  DFF_X1 u1_R11_reg_6 (.CK( clk ) , .D( u1_N357 ) , .Q( u1_R11_6 ) );
  DFF_X1 u1_R11_reg_7 (.CK( clk ) , .D( u1_N358 ) , .Q( u1_R11_7 ) );
  DFF_X1 u1_R11_reg_8 (.CK( clk ) , .D( u1_N359 ) , .Q( u1_R11_8 ) );
  DFF_X1 u1_R11_reg_9 (.CK( clk ) , .D( u1_N360 ) , .Q( u1_R11_9 ) );
  DFF_X1 u1_R12_reg_1 (.CK( clk ) , .D( u1_N384 ) , .Q( u1_R12_1 ) );
  DFF_X1 u1_R12_reg_10 (.CK( clk ) , .D( u1_N393 ) , .Q( u1_R12_10 ) );
  DFF_X1 u1_R12_reg_11 (.CK( clk ) , .D( u1_N394 ) , .Q( u1_R12_11 ) );
  DFF_X1 u1_R12_reg_12 (.CK( clk ) , .D( u1_N395 ) , .Q( u1_R12_12 ) );
  DFF_X1 u1_R12_reg_13 (.CK( clk ) , .D( u1_N396 ) , .Q( u1_R12_13 ) );
  DFF_X1 u1_R12_reg_14 (.CK( clk ) , .D( u1_N397 ) , .Q( u1_R12_14 ) );
  DFF_X1 u1_R12_reg_15 (.CK( clk ) , .D( u1_N398 ) , .Q( u1_R12_15 ) );
  DFF_X1 u1_R12_reg_16 (.CK( clk ) , .D( u1_N399 ) , .Q( u1_R12_16 ) );
  DFF_X1 u1_R12_reg_17 (.CK( clk ) , .D( u1_N400 ) , .Q( u1_R12_17 ) );
  DFF_X1 u1_R12_reg_18 (.CK( clk ) , .D( u1_N401 ) , .Q( u1_R12_18 ) );
  DFF_X1 u1_R12_reg_19 (.CK( clk ) , .D( u1_N402 ) , .Q( u1_R12_19 ) );
  DFF_X1 u1_R12_reg_2 (.CK( clk ) , .D( u1_N385 ) , .Q( u1_R12_2 ) );
  DFF_X1 u1_R12_reg_20 (.CK( clk ) , .D( u1_N403 ) , .Q( u1_R12_20 ) );
  DFF_X1 u1_R12_reg_21 (.CK( clk ) , .D( u1_N404 ) , .Q( u1_R12_21 ) );
  DFF_X1 u1_R12_reg_22 (.CK( clk ) , .D( u1_N405 ) , .Q( u1_R12_22 ) );
  DFF_X1 u1_R12_reg_23 (.CK( clk ) , .D( u1_N406 ) , .Q( u1_R12_23 ) );
  DFF_X1 u1_R12_reg_24 (.CK( clk ) , .D( u1_N407 ) , .Q( u1_R12_24 ) );
  DFF_X1 u1_R12_reg_25 (.CK( clk ) , .D( u1_N408 ) , .Q( u1_R12_25 ) );
  DFF_X1 u1_R12_reg_26 (.CK( clk ) , .D( u1_N409 ) , .Q( u1_R12_26 ) );
  DFF_X1 u1_R12_reg_27 (.CK( clk ) , .D( u1_N410 ) , .Q( u1_R12_27 ) );
  DFF_X1 u1_R12_reg_28 (.CK( clk ) , .D( u1_N411 ) , .Q( u1_R12_28 ) );
  DFF_X1 u1_R12_reg_29 (.CK( clk ) , .D( u1_N412 ) , .Q( u1_R12_29 ) );
  DFF_X1 u1_R12_reg_3 (.CK( clk ) , .D( u1_N386 ) , .Q( u1_R12_3 ) );
  DFF_X1 u1_R12_reg_30 (.CK( clk ) , .D( u1_N413 ) , .Q( u1_R12_30 ) );
  DFF_X1 u1_R12_reg_31 (.CK( clk ) , .D( u1_N414 ) , .Q( u1_R12_31 ) );
  DFF_X1 u1_R12_reg_32 (.CK( clk ) , .D( u1_N415 ) , .Q( u1_R12_32 ) );
  DFF_X1 u1_R12_reg_4 (.CK( clk ) , .D( u1_N387 ) , .Q( u1_R12_4 ) );
  DFF_X1 u1_R12_reg_5 (.CK( clk ) , .D( u1_N388 ) , .Q( u1_R12_5 ) );
  DFF_X1 u1_R12_reg_6 (.CK( clk ) , .D( u1_N389 ) , .Q( u1_R12_6 ) );
  DFF_X1 u1_R12_reg_7 (.CK( clk ) , .D( u1_N390 ) , .Q( u1_R12_7 ) );
  DFF_X1 u1_R12_reg_8 (.CK( clk ) , .D( u1_N391 ) , .Q( u1_R12_8 ) );
  DFF_X1 u1_R12_reg_9 (.CK( clk ) , .D( u1_N392 ) , .Q( u1_R12_9 ) );
  DFF_X1 u1_R13_reg_1 (.CK( clk ) , .D( u1_N416 ) , .Q( u1_R13_1 ) );
  DFF_X1 u1_R13_reg_10 (.CK( clk ) , .D( u1_N425 ) , .Q( u1_R13_10 ) );
  DFF_X1 u1_R13_reg_11 (.CK( clk ) , .D( u1_N426 ) , .Q( u1_R13_11 ) );
  DFF_X1 u1_R13_reg_12 (.CK( clk ) , .D( u1_N427 ) , .Q( u1_R13_12 ) );
  DFF_X1 u1_R13_reg_13 (.CK( clk ) , .D( u1_N428 ) , .Q( u1_R13_13 ) );
  DFF_X1 u1_R13_reg_14 (.CK( clk ) , .D( u1_N429 ) , .Q( u1_R13_14 ) );
  DFF_X1 u1_R13_reg_15 (.CK( clk ) , .D( u1_N430 ) , .Q( u1_R13_15 ) );
  DFF_X1 u1_R13_reg_16 (.CK( clk ) , .D( u1_N431 ) , .Q( u1_R13_16 ) );
  DFF_X1 u1_R13_reg_17 (.CK( clk ) , .D( u1_N432 ) , .Q( u1_R13_17 ) );
  DFF_X1 u1_R13_reg_18 (.CK( clk ) , .D( u1_N433 ) , .Q( u1_R13_18 ) );
  DFF_X1 u1_R13_reg_19 (.CK( clk ) , .D( u1_N434 ) , .Q( u1_R13_19 ) );
  DFF_X1 u1_R13_reg_2 (.CK( clk ) , .D( u1_N417 ) , .Q( u1_R13_2 ) );
  DFF_X1 u1_R13_reg_20 (.CK( clk ) , .D( u1_N435 ) , .Q( u1_R13_20 ) );
  DFF_X1 u1_R13_reg_21 (.CK( clk ) , .D( u1_N436 ) , .Q( u1_R13_21 ) );
  DFF_X1 u1_R13_reg_22 (.CK( clk ) , .D( u1_N437 ) , .Q( u1_R13_22 ) );
  DFF_X1 u1_R13_reg_23 (.CK( clk ) , .D( u1_N438 ) , .Q( u1_R13_23 ) );
  DFF_X1 u1_R13_reg_24 (.CK( clk ) , .D( u1_N439 ) , .Q( u1_R13_24 ) );
  DFF_X1 u1_R13_reg_25 (.CK( clk ) , .D( u1_N440 ) , .Q( u1_R13_25 ) );
  DFF_X1 u1_R13_reg_26 (.CK( clk ) , .D( u1_N441 ) , .Q( u1_R13_26 ) );
  DFF_X1 u1_R13_reg_27 (.CK( clk ) , .D( u1_N442 ) , .Q( u1_R13_27 ) );
  DFF_X1 u1_R13_reg_28 (.CK( clk ) , .D( u1_N443 ) , .Q( u1_R13_28 ) );
  DFF_X1 u1_R13_reg_29 (.CK( clk ) , .D( u1_N444 ) , .Q( u1_R13_29 ) );
  DFF_X1 u1_R13_reg_3 (.CK( clk ) , .D( u1_N418 ) , .Q( u1_R13_3 ) );
  DFF_X1 u1_R13_reg_30 (.CK( clk ) , .D( u1_N445 ) , .Q( u1_R13_30 ) );
  DFF_X1 u1_R13_reg_31 (.CK( clk ) , .D( u1_N446 ) , .Q( u1_R13_31 ) );
  DFF_X1 u1_R13_reg_32 (.CK( clk ) , .D( u1_N447 ) , .Q( u1_R13_32 ) );
  DFF_X1 u1_R13_reg_4 (.CK( clk ) , .D( u1_N419 ) , .Q( u1_R13_4 ) );
  DFF_X1 u1_R13_reg_5 (.CK( clk ) , .D( u1_N420 ) , .Q( u1_R13_5 ) );
  DFF_X1 u1_R13_reg_6 (.CK( clk ) , .D( u1_N421 ) , .Q( u1_R13_6 ) );
  DFF_X1 u1_R13_reg_7 (.CK( clk ) , .D( u1_N422 ) , .Q( u1_R13_7 ) );
  DFF_X1 u1_R13_reg_8 (.CK( clk ) , .D( u1_N423 ) , .Q( u1_R13_8 ) );
  DFF_X1 u1_R13_reg_9 (.CK( clk ) , .D( u1_N424 ) , .Q( u1_R13_9 ) );
  DFF_X1 u1_R14_reg_1 (.CK( clk ) , .Q( u1_FP_33 ) , .D( u1_N448 ) );
  DFF_X1 u1_R14_reg_10 (.CK( clk ) , .Q( u1_FP_42 ) , .D( u1_N457 ) );
  DFF_X1 u1_R14_reg_11 (.CK( clk ) , .Q( u1_FP_43 ) , .D( u1_N458 ) );
  DFF_X1 u1_R14_reg_12 (.CK( clk ) , .Q( u1_FP_44 ) , .D( u1_N459 ) );
  DFF_X1 u1_R14_reg_13 (.CK( clk ) , .Q( u1_FP_45 ) , .D( u1_N460 ) );
  DFF_X1 u1_R14_reg_14 (.CK( clk ) , .Q( u1_FP_46 ) , .D( u1_N461 ) );
  DFF_X1 u1_R14_reg_15 (.CK( clk ) , .Q( u1_FP_47 ) , .D( u1_N462 ) );
  DFF_X1 u1_R14_reg_16 (.CK( clk ) , .Q( u1_FP_48 ) , .D( u1_N463 ) );
  DFF_X1 u1_R14_reg_17 (.CK( clk ) , .Q( u1_FP_49 ) , .D( u1_N464 ) );
  DFF_X1 u1_R14_reg_18 (.CK( clk ) , .Q( u1_FP_50 ) , .D( u1_N465 ) );
  DFF_X1 u1_R14_reg_19 (.CK( clk ) , .Q( u1_FP_51 ) , .D( u1_N466 ) );
  DFF_X1 u1_R14_reg_2 (.CK( clk ) , .Q( u1_FP_34 ) , .D( u1_N449 ) );
  DFF_X1 u1_R14_reg_20 (.CK( clk ) , .Q( u1_FP_52 ) , .D( u1_N467 ) );
  DFF_X1 u1_R14_reg_21 (.CK( clk ) , .Q( u1_FP_53 ) , .D( u1_N468 ) );
  DFF_X1 u1_R14_reg_22 (.CK( clk ) , .Q( u1_FP_54 ) , .D( u1_N469 ) );
  DFF_X1 u1_R14_reg_23 (.CK( clk ) , .Q( u1_FP_55 ) , .D( u1_N470 ) );
  DFF_X1 u1_R14_reg_24 (.CK( clk ) , .Q( u1_FP_56 ) , .D( u1_N471 ) );
  DFF_X1 u1_R14_reg_25 (.CK( clk ) , .Q( u1_FP_57 ) , .D( u1_N472 ) );
  DFF_X1 u1_R14_reg_26 (.CK( clk ) , .Q( u1_FP_58 ) , .D( u1_N473 ) );
  DFF_X1 u1_R14_reg_27 (.CK( clk ) , .Q( u1_FP_59 ) , .D( u1_N474 ) );
  DFF_X1 u1_R14_reg_28 (.CK( clk ) , .Q( u1_FP_60 ) , .D( u1_N475 ) );
  DFF_X1 u1_R14_reg_29 (.CK( clk ) , .Q( u1_FP_61 ) , .D( u1_N476 ) );
  DFF_X1 u1_R14_reg_3 (.CK( clk ) , .Q( u1_FP_35 ) , .D( u1_N450 ) );
  DFF_X1 u1_R14_reg_30 (.CK( clk ) , .Q( u1_FP_62 ) , .D( u1_N477 ) );
  DFF_X1 u1_R14_reg_31 (.CK( clk ) , .Q( u1_FP_63 ) , .D( u1_N478 ) );
  DFF_X1 u1_R14_reg_32 (.CK( clk ) , .Q( u1_FP_64 ) , .D( u1_N479 ) );
  DFF_X1 u1_R14_reg_4 (.CK( clk ) , .Q( u1_FP_36 ) , .D( u1_N451 ) );
  DFF_X1 u1_R14_reg_5 (.CK( clk ) , .Q( u1_FP_37 ) , .D( u1_N452 ) );
  DFF_X1 u1_R14_reg_6 (.CK( clk ) , .Q( u1_FP_38 ) , .D( u1_N453 ) );
  DFF_X1 u1_R14_reg_7 (.CK( clk ) , .Q( u1_FP_39 ) , .D( u1_N454 ) );
  DFF_X1 u1_R14_reg_8 (.CK( clk ) , .Q( u1_FP_40 ) , .D( u1_N455 ) );
  DFF_X1 u1_R14_reg_9 (.CK( clk ) , .Q( u1_FP_41 ) , .D( u1_N456 ) );
  DFF_X1 u1_R1_reg_1 (.CK( clk ) , .D( u1_N32 ) , .Q( u1_R1_1 ) );
  DFF_X1 u1_R1_reg_10 (.CK( clk ) , .D( u1_N41 ) , .Q( u1_R1_10 ) );
  DFF_X1 u1_R1_reg_11 (.CK( clk ) , .D( u1_N42 ) , .Q( u1_R1_11 ) );
  DFF_X1 u1_R1_reg_12 (.CK( clk ) , .D( u1_N43 ) , .Q( u1_R1_12 ) );
  DFF_X1 u1_R1_reg_13 (.CK( clk ) , .D( u1_N44 ) , .Q( u1_R1_13 ) );
  DFF_X1 u1_R1_reg_14 (.CK( clk ) , .D( u1_N45 ) , .Q( u1_R1_14 ) );
  DFF_X1 u1_R1_reg_15 (.CK( clk ) , .D( u1_N46 ) , .Q( u1_R1_15 ) );
  DFF_X1 u1_R1_reg_16 (.CK( clk ) , .D( u1_N47 ) , .Q( u1_R1_16 ) );
  DFF_X1 u1_R1_reg_17 (.CK( clk ) , .D( u1_N48 ) , .Q( u1_R1_17 ) );
  DFF_X1 u1_R1_reg_18 (.CK( clk ) , .D( u1_N49 ) , .Q( u1_R1_18 ) );
  DFF_X1 u1_R1_reg_19 (.CK( clk ) , .D( u1_N50 ) , .Q( u1_R1_19 ) );
  DFF_X1 u1_R1_reg_2 (.CK( clk ) , .D( u1_N33 ) , .Q( u1_R1_2 ) );
  DFF_X1 u1_R1_reg_20 (.CK( clk ) , .D( u1_N51 ) , .Q( u1_R1_20 ) );
  DFF_X1 u1_R1_reg_21 (.CK( clk ) , .D( u1_N52 ) , .Q( u1_R1_21 ) );
  DFF_X1 u1_R1_reg_22 (.CK( clk ) , .D( u1_N53 ) , .Q( u1_R1_22 ) );
  DFF_X1 u1_R1_reg_23 (.CK( clk ) , .D( u1_N54 ) , .Q( u1_R1_23 ) );
  DFF_X1 u1_R1_reg_24 (.CK( clk ) , .D( u1_N55 ) , .Q( u1_R1_24 ) );
  DFF_X1 u1_R1_reg_25 (.CK( clk ) , .D( u1_N56 ) , .Q( u1_R1_25 ) );
  DFF_X1 u1_R1_reg_26 (.CK( clk ) , .D( u1_N57 ) , .Q( u1_R1_26 ) );
  DFF_X1 u1_R1_reg_27 (.CK( clk ) , .D( u1_N58 ) , .Q( u1_R1_27 ) );
  DFF_X1 u1_R1_reg_28 (.CK( clk ) , .D( u1_N59 ) , .Q( u1_R1_28 ) );
  DFF_X1 u1_R1_reg_29 (.CK( clk ) , .D( u1_N60 ) , .Q( u1_R1_29 ) );
  DFF_X1 u1_R1_reg_3 (.CK( clk ) , .D( u1_N34 ) , .Q( u1_R1_3 ) );
  DFF_X1 u1_R1_reg_30 (.CK( clk ) , .D( u1_N61 ) , .Q( u1_R1_30 ) );
  DFF_X1 u1_R1_reg_31 (.CK( clk ) , .D( u1_N62 ) , .Q( u1_R1_31 ) );
  DFF_X1 u1_R1_reg_32 (.CK( clk ) , .D( u1_N63 ) , .Q( u1_R1_32 ) );
  DFF_X1 u1_R1_reg_4 (.CK( clk ) , .D( u1_N35 ) , .Q( u1_R1_4 ) );
  DFF_X1 u1_R1_reg_5 (.CK( clk ) , .D( u1_N36 ) , .Q( u1_R1_5 ) );
  DFF_X1 u1_R1_reg_6 (.CK( clk ) , .D( u1_N37 ) , .Q( u1_R1_6 ) );
  DFF_X1 u1_R1_reg_7 (.CK( clk ) , .D( u1_N38 ) , .Q( u1_R1_7 ) );
  DFF_X1 u1_R1_reg_8 (.CK( clk ) , .D( u1_N39 ) , .Q( u1_R1_8 ) );
  DFF_X1 u1_R1_reg_9 (.CK( clk ) , .D( u1_N40 ) , .Q( u1_R1_9 ) );
  DFF_X1 u1_R2_reg_1 (.CK( clk ) , .D( u1_N64 ) , .Q( u1_R2_1 ) );
  DFF_X1 u1_R2_reg_10 (.CK( clk ) , .D( u1_N73 ) , .Q( u1_R2_10 ) );
  DFF_X1 u1_R2_reg_11 (.CK( clk ) , .D( u1_N74 ) , .Q( u1_R2_11 ) );
  DFF_X1 u1_R2_reg_12 (.CK( clk ) , .D( u1_N75 ) , .Q( u1_R2_12 ) );
  DFF_X1 u1_R2_reg_13 (.CK( clk ) , .D( u1_N76 ) , .Q( u1_R2_13 ) );
  DFF_X1 u1_R2_reg_14 (.CK( clk ) , .D( u1_N77 ) , .Q( u1_R2_14 ) );
  DFF_X1 u1_R2_reg_15 (.CK( clk ) , .D( u1_N78 ) , .Q( u1_R2_15 ) );
  DFF_X1 u1_R2_reg_16 (.CK( clk ) , .D( u1_N79 ) , .Q( u1_R2_16 ) );
  DFF_X1 u1_R2_reg_17 (.CK( clk ) , .D( u1_N80 ) , .Q( u1_R2_17 ) );
  DFF_X1 u1_R2_reg_18 (.CK( clk ) , .D( u1_N81 ) , .Q( u1_R2_18 ) );
  DFF_X1 u1_R2_reg_19 (.CK( clk ) , .D( u1_N82 ) , .Q( u1_R2_19 ) );
  DFF_X1 u1_R2_reg_2 (.CK( clk ) , .D( u1_N65 ) , .Q( u1_R2_2 ) );
  DFF_X1 u1_R2_reg_20 (.CK( clk ) , .D( u1_N83 ) , .Q( u1_R2_20 ) );
  DFF_X1 u1_R2_reg_21 (.CK( clk ) , .D( u1_N84 ) , .Q( u1_R2_21 ) );
  DFF_X1 u1_R2_reg_22 (.CK( clk ) , .D( u1_N85 ) , .Q( u1_R2_22 ) );
  DFF_X1 u1_R2_reg_23 (.CK( clk ) , .D( u1_N86 ) , .Q( u1_R2_23 ) );
  DFF_X1 u1_R2_reg_24 (.CK( clk ) , .D( u1_N87 ) , .Q( u1_R2_24 ) );
  DFF_X1 u1_R2_reg_25 (.CK( clk ) , .D( u1_N88 ) , .Q( u1_R2_25 ) );
  DFF_X1 u1_R2_reg_26 (.CK( clk ) , .D( u1_N89 ) , .Q( u1_R2_26 ) );
  DFF_X1 u1_R2_reg_27 (.CK( clk ) , .D( u1_N90 ) , .Q( u1_R2_27 ) );
  DFF_X1 u1_R2_reg_28 (.CK( clk ) , .D( u1_N91 ) , .Q( u1_R2_28 ) );
  DFF_X1 u1_R2_reg_29 (.CK( clk ) , .D( u1_N92 ) , .Q( u1_R2_29 ) );
  DFF_X1 u1_R2_reg_3 (.CK( clk ) , .D( u1_N66 ) , .Q( u1_R2_3 ) );
  DFF_X1 u1_R2_reg_30 (.CK( clk ) , .D( u1_N93 ) , .Q( u1_R2_30 ) );
  DFF_X1 u1_R2_reg_31 (.CK( clk ) , .D( u1_N94 ) , .Q( u1_R2_31 ) );
  DFF_X1 u1_R2_reg_32 (.CK( clk ) , .D( u1_N95 ) , .Q( u1_R2_32 ) );
  DFF_X1 u1_R2_reg_4 (.CK( clk ) , .D( u1_N67 ) , .Q( u1_R2_4 ) );
  DFF_X1 u1_R2_reg_5 (.CK( clk ) , .D( u1_N68 ) , .Q( u1_R2_5 ) );
  DFF_X1 u1_R2_reg_6 (.CK( clk ) , .D( u1_N69 ) , .Q( u1_R2_6 ) );
  DFF_X1 u1_R2_reg_7 (.CK( clk ) , .D( u1_N70 ) , .Q( u1_R2_7 ) );
  DFF_X1 u1_R2_reg_8 (.CK( clk ) , .D( u1_N71 ) , .Q( u1_R2_8 ) );
  DFF_X1 u1_R2_reg_9 (.CK( clk ) , .D( u1_N72 ) , .Q( u1_R2_9 ) );
  DFF_X1 u1_R3_reg_1 (.CK( clk ) , .D( u1_N96 ) , .Q( u1_R3_1 ) );
  DFF_X1 u1_R3_reg_10 (.CK( clk ) , .D( u1_N105 ) , .Q( u1_R3_10 ) );
  DFF_X1 u1_R3_reg_11 (.CK( clk ) , .D( u1_N106 ) , .Q( u1_R3_11 ) );
  DFF_X1 u1_R3_reg_12 (.CK( clk ) , .D( u1_N107 ) , .Q( u1_R3_12 ) );
  DFF_X1 u1_R3_reg_13 (.CK( clk ) , .D( u1_N108 ) , .Q( u1_R3_13 ) );
  DFF_X1 u1_R3_reg_14 (.CK( clk ) , .D( u1_N109 ) , .Q( u1_R3_14 ) );
  DFF_X1 u1_R3_reg_15 (.CK( clk ) , .D( u1_N110 ) , .Q( u1_R3_15 ) );
  DFF_X1 u1_R3_reg_16 (.CK( clk ) , .D( u1_N111 ) , .Q( u1_R3_16 ) );
  DFF_X1 u1_R3_reg_17 (.CK( clk ) , .D( u1_N112 ) , .Q( u1_R3_17 ) );
  DFF_X1 u1_R3_reg_18 (.CK( clk ) , .D( u1_N113 ) , .Q( u1_R3_18 ) );
  DFF_X1 u1_R3_reg_19 (.CK( clk ) , .D( u1_N114 ) , .Q( u1_R3_19 ) );
  DFF_X1 u1_R3_reg_2 (.CK( clk ) , .D( u1_N97 ) , .Q( u1_R3_2 ) );
  DFF_X1 u1_R3_reg_20 (.CK( clk ) , .D( u1_N115 ) , .Q( u1_R3_20 ) );
  DFF_X1 u1_R3_reg_21 (.CK( clk ) , .D( u1_N116 ) , .Q( u1_R3_21 ) );
  DFF_X1 u1_R3_reg_22 (.CK( clk ) , .D( u1_N117 ) , .Q( u1_R3_22 ) );
  DFF_X1 u1_R3_reg_23 (.CK( clk ) , .D( u1_N118 ) , .Q( u1_R3_23 ) );
  DFF_X1 u1_R3_reg_24 (.CK( clk ) , .D( u1_N119 ) , .Q( u1_R3_24 ) );
  DFF_X1 u1_R3_reg_25 (.CK( clk ) , .D( u1_N120 ) , .Q( u1_R3_25 ) );
  DFF_X1 u1_R3_reg_26 (.CK( clk ) , .D( u1_N121 ) , .Q( u1_R3_26 ) );
  DFF_X1 u1_R3_reg_27 (.CK( clk ) , .D( u1_N122 ) , .Q( u1_R3_27 ) );
  DFF_X1 u1_R3_reg_28 (.CK( clk ) , .D( u1_N123 ) , .Q( u1_R3_28 ) );
  DFF_X1 u1_R3_reg_29 (.CK( clk ) , .D( u1_N124 ) , .Q( u1_R3_29 ) );
  DFF_X1 u1_R3_reg_3 (.CK( clk ) , .D( u1_N98 ) , .Q( u1_R3_3 ) );
  DFF_X1 u1_R3_reg_30 (.CK( clk ) , .D( u1_N125 ) , .Q( u1_R3_30 ) );
  DFF_X1 u1_R3_reg_31 (.CK( clk ) , .D( u1_N126 ) , .Q( u1_R3_31 ) );
  DFF_X1 u1_R3_reg_32 (.CK( clk ) , .D( u1_N127 ) , .Q( u1_R3_32 ) );
  DFF_X1 u1_R3_reg_4 (.CK( clk ) , .D( u1_N99 ) , .Q( u1_R3_4 ) );
  DFF_X1 u1_R3_reg_5 (.CK( clk ) , .D( u1_N100 ) , .Q( u1_R3_5 ) );
  DFF_X1 u1_R3_reg_6 (.CK( clk ) , .D( u1_N101 ) , .Q( u1_R3_6 ) );
  DFF_X1 u1_R3_reg_7 (.CK( clk ) , .D( u1_N102 ) , .Q( u1_R3_7 ) );
  DFF_X1 u1_R3_reg_8 (.CK( clk ) , .D( u1_N103 ) , .Q( u1_R3_8 ) );
  DFF_X1 u1_R3_reg_9 (.CK( clk ) , .D( u1_N104 ) , .Q( u1_R3_9 ) );
  DFF_X1 u1_R4_reg_1 (.CK( clk ) , .D( u1_N128 ) , .Q( u1_R4_1 ) );
  DFF_X1 u1_R4_reg_10 (.CK( clk ) , .D( u1_N137 ) , .Q( u1_R4_10 ) );
  DFF_X1 u1_R4_reg_11 (.CK( clk ) , .D( u1_N138 ) , .Q( u1_R4_11 ) );
  DFF_X1 u1_R4_reg_12 (.CK( clk ) , .D( u1_N139 ) , .Q( u1_R4_12 ) );
  DFF_X1 u1_R4_reg_13 (.CK( clk ) , .D( u1_N140 ) , .Q( u1_R4_13 ) );
  DFF_X1 u1_R4_reg_14 (.CK( clk ) , .D( u1_N141 ) , .Q( u1_R4_14 ) );
  DFF_X1 u1_R4_reg_15 (.CK( clk ) , .D( u1_N142 ) , .Q( u1_R4_15 ) );
  DFF_X1 u1_R4_reg_16 (.CK( clk ) , .D( u1_N143 ) , .Q( u1_R4_16 ) );
  DFF_X1 u1_R4_reg_17 (.CK( clk ) , .D( u1_N144 ) , .Q( u1_R4_17 ) );
  DFF_X1 u1_R4_reg_18 (.CK( clk ) , .D( u1_N145 ) , .Q( u1_R4_18 ) );
  DFF_X1 u1_R4_reg_19 (.CK( clk ) , .D( u1_N146 ) , .Q( u1_R4_19 ) );
  DFF_X1 u1_R4_reg_2 (.CK( clk ) , .D( u1_N129 ) , .Q( u1_R4_2 ) );
  DFF_X1 u1_R4_reg_20 (.CK( clk ) , .D( u1_N147 ) , .Q( u1_R4_20 ) );
  DFF_X1 u1_R4_reg_21 (.CK( clk ) , .D( u1_N148 ) , .Q( u1_R4_21 ) );
  DFF_X1 u1_R4_reg_22 (.CK( clk ) , .D( u1_N149 ) , .Q( u1_R4_22 ) );
  DFF_X1 u1_R4_reg_23 (.CK( clk ) , .D( u1_N150 ) , .Q( u1_R4_23 ) );
  DFF_X1 u1_R4_reg_24 (.CK( clk ) , .D( u1_N151 ) , .Q( u1_R4_24 ) );
  DFF_X1 u1_R4_reg_25 (.CK( clk ) , .D( u1_N152 ) , .Q( u1_R4_25 ) );
  DFF_X1 u1_R4_reg_26 (.CK( clk ) , .D( u1_N153 ) , .Q( u1_R4_26 ) );
  DFF_X1 u1_R4_reg_27 (.CK( clk ) , .D( u1_N154 ) , .Q( u1_R4_27 ) );
  DFF_X1 u1_R4_reg_28 (.CK( clk ) , .D( u1_N155 ) , .Q( u1_R4_28 ) );
  DFF_X1 u1_R4_reg_29 (.CK( clk ) , .D( u1_N156 ) , .Q( u1_R4_29 ) );
  DFF_X1 u1_R4_reg_3 (.CK( clk ) , .D( u1_N130 ) , .Q( u1_R4_3 ) );
  DFF_X1 u1_R4_reg_30 (.CK( clk ) , .D( u1_N157 ) , .Q( u1_R4_30 ) );
  DFF_X1 u1_R4_reg_31 (.CK( clk ) , .D( u1_N158 ) , .Q( u1_R4_31 ) );
  DFF_X1 u1_R4_reg_32 (.CK( clk ) , .D( u1_N159 ) , .Q( u1_R4_32 ) );
  DFF_X1 u1_R4_reg_4 (.CK( clk ) , .D( u1_N131 ) , .Q( u1_R4_4 ) );
  DFF_X1 u1_R4_reg_5 (.CK( clk ) , .D( u1_N132 ) , .Q( u1_R4_5 ) );
  DFF_X1 u1_R4_reg_6 (.CK( clk ) , .D( u1_N133 ) , .Q( u1_R4_6 ) );
  DFF_X1 u1_R4_reg_7 (.CK( clk ) , .D( u1_N134 ) , .Q( u1_R4_7 ) );
  DFF_X1 u1_R4_reg_8 (.CK( clk ) , .D( u1_N135 ) , .Q( u1_R4_8 ) );
  DFF_X1 u1_R4_reg_9 (.CK( clk ) , .D( u1_N136 ) , .Q( u1_R4_9 ) );
  DFF_X1 u1_R5_reg_1 (.CK( clk ) , .D( u1_N160 ) , .Q( u1_R5_1 ) );
  DFF_X1 u1_R5_reg_10 (.CK( clk ) , .D( u1_N169 ) , .Q( u1_R5_10 ) );
  DFF_X1 u1_R5_reg_11 (.CK( clk ) , .D( u1_N170 ) , .Q( u1_R5_11 ) );
  DFF_X1 u1_R5_reg_12 (.CK( clk ) , .D( u1_N171 ) , .Q( u1_R5_12 ) );
  DFF_X1 u1_R5_reg_13 (.CK( clk ) , .D( u1_N172 ) , .Q( u1_R5_13 ) );
  DFF_X1 u1_R5_reg_14 (.CK( clk ) , .D( u1_N173 ) , .Q( u1_R5_14 ) );
  DFF_X1 u1_R5_reg_15 (.CK( clk ) , .D( u1_N174 ) , .Q( u1_R5_15 ) );
  DFF_X1 u1_R5_reg_16 (.CK( clk ) , .D( u1_N175 ) , .Q( u1_R5_16 ) );
  DFF_X1 u1_R5_reg_17 (.CK( clk ) , .D( u1_N176 ) , .Q( u1_R5_17 ) );
  DFF_X1 u1_R5_reg_18 (.CK( clk ) , .D( u1_N177 ) , .Q( u1_R5_18 ) );
  DFF_X1 u1_R5_reg_19 (.CK( clk ) , .D( u1_N178 ) , .Q( u1_R5_19 ) );
  DFF_X1 u1_R5_reg_2 (.CK( clk ) , .D( u1_N161 ) , .Q( u1_R5_2 ) );
  DFF_X1 u1_R5_reg_20 (.CK( clk ) , .D( u1_N179 ) , .Q( u1_R5_20 ) );
  DFF_X1 u1_R5_reg_21 (.CK( clk ) , .D( u1_N180 ) , .Q( u1_R5_21 ) );
  DFF_X1 u1_R5_reg_22 (.CK( clk ) , .D( u1_N181 ) , .Q( u1_R5_22 ) );
  DFF_X1 u1_R5_reg_23 (.CK( clk ) , .D( u1_N182 ) , .Q( u1_R5_23 ) );
  DFF_X1 u1_R5_reg_24 (.CK( clk ) , .D( u1_N183 ) , .Q( u1_R5_24 ) );
  DFF_X1 u1_R5_reg_25 (.CK( clk ) , .D( u1_N184 ) , .Q( u1_R5_25 ) );
  DFF_X1 u1_R5_reg_26 (.CK( clk ) , .D( u1_N185 ) , .Q( u1_R5_26 ) );
  DFF_X1 u1_R5_reg_27 (.CK( clk ) , .D( u1_N186 ) , .Q( u1_R5_27 ) );
  DFF_X1 u1_R5_reg_28 (.CK( clk ) , .D( u1_N187 ) , .Q( u1_R5_28 ) );
  DFF_X1 u1_R5_reg_29 (.CK( clk ) , .D( u1_N188 ) , .Q( u1_R5_29 ) );
  DFF_X1 u1_R5_reg_3 (.CK( clk ) , .D( u1_N162 ) , .Q( u1_R5_3 ) );
  DFF_X1 u1_R5_reg_30 (.CK( clk ) , .D( u1_N189 ) , .Q( u1_R5_30 ) );
  DFF_X1 u1_R5_reg_31 (.CK( clk ) , .D( u1_N190 ) , .Q( u1_R5_31 ) );
  DFF_X1 u1_R5_reg_32 (.CK( clk ) , .D( u1_N191 ) , .Q( u1_R5_32 ) );
  DFF_X1 u1_R5_reg_4 (.CK( clk ) , .D( u1_N163 ) , .Q( u1_R5_4 ) );
  DFF_X1 u1_R5_reg_5 (.CK( clk ) , .D( u1_N164 ) , .Q( u1_R5_5 ) );
  DFF_X1 u1_R5_reg_6 (.CK( clk ) , .D( u1_N165 ) , .Q( u1_R5_6 ) );
  DFF_X1 u1_R5_reg_7 (.CK( clk ) , .D( u1_N166 ) , .Q( u1_R5_7 ) );
  DFF_X1 u1_R5_reg_8 (.CK( clk ) , .D( u1_N167 ) , .Q( u1_R5_8 ) );
  DFF_X1 u1_R5_reg_9 (.CK( clk ) , .D( u1_N168 ) , .Q( u1_R5_9 ) );
  DFF_X1 u1_R6_reg_1 (.CK( clk ) , .D( u1_N192 ) , .Q( u1_R6_1 ) );
  DFF_X1 u1_R6_reg_10 (.CK( clk ) , .D( u1_N201 ) , .Q( u1_R6_10 ) );
  DFF_X1 u1_R6_reg_11 (.CK( clk ) , .D( u1_N202 ) , .Q( u1_R6_11 ) );
  DFF_X1 u1_R6_reg_12 (.CK( clk ) , .D( u1_N203 ) , .Q( u1_R6_12 ) );
  DFF_X1 u1_R6_reg_13 (.CK( clk ) , .D( u1_N204 ) , .Q( u1_R6_13 ) );
  DFF_X1 u1_R6_reg_14 (.CK( clk ) , .D( u1_N205 ) , .Q( u1_R6_14 ) );
  DFF_X1 u1_R6_reg_15 (.CK( clk ) , .D( u1_N206 ) , .Q( u1_R6_15 ) );
  DFF_X1 u1_R6_reg_16 (.CK( clk ) , .D( u1_N207 ) , .Q( u1_R6_16 ) );
  DFF_X1 u1_R6_reg_17 (.CK( clk ) , .D( u1_N208 ) , .Q( u1_R6_17 ) );
  DFF_X1 u1_R6_reg_18 (.CK( clk ) , .D( u1_N209 ) , .Q( u1_R6_18 ) );
  DFF_X1 u1_R6_reg_19 (.CK( clk ) , .D( u1_N210 ) , .Q( u1_R6_19 ) );
  DFF_X1 u1_R6_reg_2 (.CK( clk ) , .D( u1_N193 ) , .Q( u1_R6_2 ) );
  DFF_X1 u1_R6_reg_20 (.CK( clk ) , .D( u1_N211 ) , .Q( u1_R6_20 ) );
  DFF_X1 u1_R6_reg_21 (.CK( clk ) , .D( u1_N212 ) , .Q( u1_R6_21 ) );
  DFF_X1 u1_R6_reg_22 (.CK( clk ) , .D( u1_N213 ) , .Q( u1_R6_22 ) );
  DFF_X1 u1_R6_reg_23 (.CK( clk ) , .D( u1_N214 ) , .Q( u1_R6_23 ) );
  DFF_X1 u1_R6_reg_24 (.CK( clk ) , .D( u1_N215 ) , .Q( u1_R6_24 ) );
  DFF_X1 u1_R6_reg_25 (.CK( clk ) , .D( u1_N216 ) , .Q( u1_R6_25 ) );
  DFF_X1 u1_R6_reg_26 (.CK( clk ) , .D( u1_N217 ) , .Q( u1_R6_26 ) );
  DFF_X1 u1_R6_reg_27 (.CK( clk ) , .D( u1_N218 ) , .Q( u1_R6_27 ) );
  DFF_X1 u1_R6_reg_28 (.CK( clk ) , .D( u1_N219 ) , .Q( u1_R6_28 ) );
  DFF_X1 u1_R6_reg_29 (.CK( clk ) , .D( u1_N220 ) , .Q( u1_R6_29 ) );
  DFF_X1 u1_R6_reg_3 (.CK( clk ) , .D( u1_N194 ) , .Q( u1_R6_3 ) );
  DFF_X1 u1_R6_reg_30 (.CK( clk ) , .D( u1_N221 ) , .Q( u1_R6_30 ) );
  DFF_X1 u1_R6_reg_31 (.CK( clk ) , .D( u1_N222 ) , .Q( u1_R6_31 ) );
  DFF_X1 u1_R6_reg_32 (.CK( clk ) , .D( u1_N223 ) , .Q( u1_R6_32 ) );
  DFF_X1 u1_R6_reg_4 (.CK( clk ) , .D( u1_N195 ) , .Q( u1_R6_4 ) );
  DFF_X1 u1_R6_reg_5 (.CK( clk ) , .D( u1_N196 ) , .Q( u1_R6_5 ) );
  DFF_X1 u1_R6_reg_6 (.CK( clk ) , .D( u1_N197 ) , .Q( u1_R6_6 ) );
  DFF_X1 u1_R6_reg_7 (.CK( clk ) , .D( u1_N198 ) , .Q( u1_R6_7 ) );
  DFF_X1 u1_R6_reg_8 (.CK( clk ) , .D( u1_N199 ) , .Q( u1_R6_8 ) );
  DFF_X1 u1_R6_reg_9 (.CK( clk ) , .D( u1_N200 ) , .Q( u1_R6_9 ) );
  DFF_X1 u1_R7_reg_1 (.CK( clk ) , .D( u1_N224 ) , .Q( u1_R7_1 ) );
  DFF_X1 u1_R7_reg_10 (.CK( clk ) , .D( u1_N233 ) , .Q( u1_R7_10 ) );
  DFF_X1 u1_R7_reg_11 (.CK( clk ) , .D( u1_N234 ) , .Q( u1_R7_11 ) );
  DFF_X1 u1_R7_reg_12 (.CK( clk ) , .D( u1_N235 ) , .Q( u1_R7_12 ) );
  DFF_X1 u1_R7_reg_13 (.CK( clk ) , .D( u1_N236 ) , .Q( u1_R7_13 ) );
  DFF_X1 u1_R7_reg_14 (.CK( clk ) , .D( u1_N237 ) , .Q( u1_R7_14 ) );
  DFF_X1 u1_R7_reg_15 (.CK( clk ) , .D( u1_N238 ) , .Q( u1_R7_15 ) );
  DFF_X1 u1_R7_reg_16 (.CK( clk ) , .D( u1_N239 ) , .Q( u1_R7_16 ) );
  DFF_X1 u1_R7_reg_17 (.CK( clk ) , .D( u1_N240 ) , .Q( u1_R7_17 ) );
  DFF_X1 u1_R7_reg_18 (.CK( clk ) , .D( u1_N241 ) , .Q( u1_R7_18 ) );
  DFF_X1 u1_R7_reg_19 (.CK( clk ) , .D( u1_N242 ) , .Q( u1_R7_19 ) );
  DFF_X1 u1_R7_reg_2 (.CK( clk ) , .D( u1_N225 ) , .Q( u1_R7_2 ) );
  DFF_X1 u1_R7_reg_20 (.CK( clk ) , .D( u1_N243 ) , .Q( u1_R7_20 ) );
  DFF_X1 u1_R7_reg_21 (.CK( clk ) , .D( u1_N244 ) , .Q( u1_R7_21 ) );
  DFF_X1 u1_R7_reg_22 (.CK( clk ) , .D( u1_N245 ) , .Q( u1_R7_22 ) );
  DFF_X1 u1_R7_reg_23 (.CK( clk ) , .D( u1_N246 ) , .Q( u1_R7_23 ) );
  DFF_X1 u1_R7_reg_24 (.CK( clk ) , .D( u1_N247 ) , .Q( u1_R7_24 ) );
  DFF_X1 u1_R7_reg_25 (.CK( clk ) , .D( u1_N248 ) , .Q( u1_R7_25 ) );
  DFF_X1 u1_R7_reg_26 (.CK( clk ) , .D( u1_N249 ) , .Q( u1_R7_26 ) );
  DFF_X1 u1_R7_reg_27 (.CK( clk ) , .D( u1_N250 ) , .Q( u1_R7_27 ) );
  DFF_X1 u1_R7_reg_28 (.CK( clk ) , .D( u1_N251 ) , .Q( u1_R7_28 ) );
  DFF_X1 u1_R7_reg_29 (.CK( clk ) , .D( u1_N252 ) , .Q( u1_R7_29 ) );
  DFF_X1 u1_R7_reg_3 (.CK( clk ) , .D( u1_N226 ) , .Q( u1_R7_3 ) );
  DFF_X1 u1_R7_reg_30 (.CK( clk ) , .D( u1_N253 ) , .Q( u1_R7_30 ) );
  DFF_X1 u1_R7_reg_31 (.CK( clk ) , .D( u1_N254 ) , .Q( u1_R7_31 ) );
  DFF_X1 u1_R7_reg_32 (.CK( clk ) , .D( u1_N255 ) , .Q( u1_R7_32 ) );
  DFF_X1 u1_R7_reg_4 (.CK( clk ) , .D( u1_N227 ) , .Q( u1_R7_4 ) );
  DFF_X1 u1_R7_reg_5 (.CK( clk ) , .D( u1_N228 ) , .Q( u1_R7_5 ) );
  DFF_X1 u1_R7_reg_6 (.CK( clk ) , .D( u1_N229 ) , .Q( u1_R7_6 ) );
  DFF_X1 u1_R7_reg_7 (.CK( clk ) , .D( u1_N230 ) , .Q( u1_R7_7 ) );
  DFF_X1 u1_R7_reg_8 (.CK( clk ) , .D( u1_N231 ) , .Q( u1_R7_8 ) );
  DFF_X1 u1_R7_reg_9 (.CK( clk ) , .D( u1_N232 ) , .Q( u1_R7_9 ) );
  DFF_X1 u1_R8_reg_1 (.CK( clk ) , .D( u1_N256 ) , .Q( u1_R8_1 ) );
  DFF_X1 u1_R8_reg_10 (.CK( clk ) , .D( u1_N265 ) , .Q( u1_R8_10 ) );
  DFF_X1 u1_R8_reg_11 (.CK( clk ) , .D( u1_N266 ) , .Q( u1_R8_11 ) );
  DFF_X1 u1_R8_reg_12 (.CK( clk ) , .D( u1_N267 ) , .Q( u1_R8_12 ) );
  DFF_X1 u1_R8_reg_13 (.CK( clk ) , .D( u1_N268 ) , .Q( u1_R8_13 ) );
  DFF_X1 u1_R8_reg_14 (.CK( clk ) , .D( u1_N269 ) , .Q( u1_R8_14 ) );
  DFF_X1 u1_R8_reg_15 (.CK( clk ) , .D( u1_N270 ) , .Q( u1_R8_15 ) );
  DFF_X1 u1_R8_reg_16 (.CK( clk ) , .D( u1_N271 ) , .Q( u1_R8_16 ) );
  DFF_X1 u1_R8_reg_17 (.CK( clk ) , .D( u1_N272 ) , .Q( u1_R8_17 ) );
  DFF_X1 u1_R8_reg_18 (.CK( clk ) , .D( u1_N273 ) , .Q( u1_R8_18 ) );
  DFF_X1 u1_R8_reg_19 (.CK( clk ) , .D( u1_N274 ) , .Q( u1_R8_19 ) );
  DFF_X1 u1_R8_reg_2 (.CK( clk ) , .D( u1_N257 ) , .Q( u1_R8_2 ) );
  DFF_X1 u1_R8_reg_20 (.CK( clk ) , .D( u1_N275 ) , .Q( u1_R8_20 ) );
  DFF_X1 u1_R8_reg_21 (.CK( clk ) , .D( u1_N276 ) , .Q( u1_R8_21 ) );
  DFF_X1 u1_R8_reg_22 (.CK( clk ) , .D( u1_N277 ) , .Q( u1_R8_22 ) );
  DFF_X1 u1_R8_reg_23 (.CK( clk ) , .D( u1_N278 ) , .Q( u1_R8_23 ) );
  DFF_X1 u1_R8_reg_24 (.CK( clk ) , .D( u1_N279 ) , .Q( u1_R8_24 ) );
  DFF_X1 u1_R8_reg_25 (.CK( clk ) , .D( u1_N280 ) , .Q( u1_R8_25 ) );
  DFF_X1 u1_R8_reg_26 (.CK( clk ) , .D( u1_N281 ) , .Q( u1_R8_26 ) );
  DFF_X1 u1_R8_reg_27 (.CK( clk ) , .D( u1_N282 ) , .Q( u1_R8_27 ) );
  DFF_X1 u1_R8_reg_28 (.CK( clk ) , .D( u1_N283 ) , .Q( u1_R8_28 ) );
  DFF_X1 u1_R8_reg_29 (.CK( clk ) , .D( u1_N284 ) , .Q( u1_R8_29 ) );
  DFF_X1 u1_R8_reg_3 (.CK( clk ) , .D( u1_N258 ) , .Q( u1_R8_3 ) );
  DFF_X1 u1_R8_reg_30 (.CK( clk ) , .D( u1_N285 ) , .Q( u1_R8_30 ) );
  DFF_X1 u1_R8_reg_31 (.CK( clk ) , .D( u1_N286 ) , .Q( u1_R8_31 ) );
  DFF_X1 u1_R8_reg_32 (.CK( clk ) , .D( u1_N287 ) , .Q( u1_R8_32 ) );
  DFF_X1 u1_R8_reg_4 (.CK( clk ) , .D( u1_N259 ) , .Q( u1_R8_4 ) );
  DFF_X1 u1_R8_reg_5 (.CK( clk ) , .D( u1_N260 ) , .Q( u1_R8_5 ) );
  DFF_X1 u1_R8_reg_6 (.CK( clk ) , .D( u1_N261 ) , .Q( u1_R8_6 ) );
  DFF_X1 u1_R8_reg_7 (.CK( clk ) , .D( u1_N262 ) , .Q( u1_R8_7 ) );
  DFF_X1 u1_R8_reg_8 (.CK( clk ) , .D( u1_N263 ) , .Q( u1_R8_8 ) );
  DFF_X1 u1_R8_reg_9 (.CK( clk ) , .D( u1_N264 ) , .Q( u1_R8_9 ) );
  DFF_X1 u1_R9_reg_1 (.CK( clk ) , .D( u1_N288 ) , .Q( u1_R9_1 ) );
  DFF_X1 u1_R9_reg_10 (.CK( clk ) , .D( u1_N297 ) , .Q( u1_R9_10 ) );
  DFF_X1 u1_R9_reg_11 (.CK( clk ) , .D( u1_N298 ) , .Q( u1_R9_11 ) );
  DFF_X1 u1_R9_reg_12 (.CK( clk ) , .D( u1_N299 ) , .Q( u1_R9_12 ) );
  DFF_X1 u1_R9_reg_13 (.CK( clk ) , .D( u1_N300 ) , .Q( u1_R9_13 ) );
  DFF_X1 u1_R9_reg_14 (.CK( clk ) , .D( u1_N301 ) , .Q( u1_R9_14 ) );
  DFF_X1 u1_R9_reg_15 (.CK( clk ) , .D( u1_N302 ) , .Q( u1_R9_15 ) );
  DFF_X1 u1_R9_reg_16 (.CK( clk ) , .D( u1_N303 ) , .Q( u1_R9_16 ) );
  DFF_X1 u1_R9_reg_17 (.CK( clk ) , .D( u1_N304 ) , .Q( u1_R9_17 ) );
  DFF_X1 u1_R9_reg_18 (.CK( clk ) , .D( u1_N305 ) , .Q( u1_R9_18 ) );
  DFF_X1 u1_R9_reg_19 (.CK( clk ) , .D( u1_N306 ) , .Q( u1_R9_19 ) );
  DFF_X1 u1_R9_reg_2 (.CK( clk ) , .D( u1_N289 ) , .Q( u1_R9_2 ) );
  DFF_X1 u1_R9_reg_20 (.CK( clk ) , .D( u1_N307 ) , .Q( u1_R9_20 ) );
  DFF_X1 u1_R9_reg_21 (.CK( clk ) , .D( u1_N308 ) , .Q( u1_R9_21 ) );
  DFF_X1 u1_R9_reg_22 (.CK( clk ) , .D( u1_N309 ) , .Q( u1_R9_22 ) );
  DFF_X1 u1_R9_reg_23 (.CK( clk ) , .D( u1_N310 ) , .Q( u1_R9_23 ) );
  DFF_X1 u1_R9_reg_24 (.CK( clk ) , .D( u1_N311 ) , .Q( u1_R9_24 ) );
  DFF_X1 u1_R9_reg_25 (.CK( clk ) , .D( u1_N312 ) , .Q( u1_R9_25 ) );
  DFF_X1 u1_R9_reg_26 (.CK( clk ) , .D( u1_N313 ) , .Q( u1_R9_26 ) );
  DFF_X1 u1_R9_reg_27 (.CK( clk ) , .D( u1_N314 ) , .Q( u1_R9_27 ) );
  DFF_X1 u1_R9_reg_28 (.CK( clk ) , .D( u1_N315 ) , .Q( u1_R9_28 ) );
  DFF_X1 u1_R9_reg_29 (.CK( clk ) , .D( u1_N316 ) , .Q( u1_R9_29 ) );
  DFF_X1 u1_R9_reg_3 (.CK( clk ) , .D( u1_N290 ) , .Q( u1_R9_3 ) );
  DFF_X1 u1_R9_reg_30 (.CK( clk ) , .D( u1_N317 ) , .Q( u1_R9_30 ) );
  DFF_X1 u1_R9_reg_31 (.CK( clk ) , .D( u1_N318 ) , .Q( u1_R9_31 ) );
  DFF_X1 u1_R9_reg_32 (.CK( clk ) , .D( u1_N319 ) , .Q( u1_R9_32 ) );
  DFF_X1 u1_R9_reg_4 (.CK( clk ) , .D( u1_N291 ) , .Q( u1_R9_4 ) );
  DFF_X1 u1_R9_reg_5 (.CK( clk ) , .D( u1_N292 ) , .Q( u1_R9_5 ) );
  DFF_X1 u1_R9_reg_6 (.CK( clk ) , .D( u1_N293 ) , .Q( u1_R9_6 ) );
  DFF_X1 u1_R9_reg_7 (.CK( clk ) , .D( u1_N294 ) , .Q( u1_R9_7 ) );
  DFF_X1 u1_R9_reg_8 (.CK( clk ) , .D( u1_N295 ) , .Q( u1_R9_8 ) );
  DFF_X1 u1_R9_reg_9 (.CK( clk ) , .D( u1_N296 ) , .Q( u1_R9_9 ) );
  DFF_X1 u1_desIn_r_reg_0 (.CK( clk ) , .D( stage1_out_0 ) , .Q( u1_desIn_r_0 ) );
  DFF_X1 u1_desIn_r_reg_1 (.CK( clk ) , .D( stage1_out_1 ) , .Q( u1_desIn_r_1 ) );
  DFF_X1 u1_desIn_r_reg_10 (.CK( clk ) , .D( stage1_out_10 ) , .Q( u1_desIn_r_10 ) );
  DFF_X1 u1_desIn_r_reg_11 (.CK( clk ) , .D( stage1_out_11 ) , .Q( u1_desIn_r_11 ) );
  DFF_X1 u1_desIn_r_reg_12 (.CK( clk ) , .D( stage1_out_12 ) , .Q( u1_desIn_r_12 ) );
  DFF_X1 u1_desIn_r_reg_13 (.CK( clk ) , .D( stage1_out_13 ) , .Q( u1_desIn_r_13 ) );
  DFF_X1 u1_desIn_r_reg_14 (.CK( clk ) , .D( stage1_out_14 ) , .Q( u1_desIn_r_14 ) );
  DFF_X1 u1_desIn_r_reg_15 (.CK( clk ) , .D( stage1_out_15 ) , .Q( u1_desIn_r_15 ) );
  DFF_X1 u1_desIn_r_reg_16 (.CK( clk ) , .D( stage1_out_16 ) , .Q( u1_desIn_r_16 ) );
  DFF_X1 u1_desIn_r_reg_17 (.CK( clk ) , .D( stage1_out_17 ) , .Q( u1_desIn_r_17 ) );
  DFF_X1 u1_desIn_r_reg_18 (.CK( clk ) , .D( stage1_out_18 ) , .Q( u1_desIn_r_18 ) );
  DFF_X1 u1_desIn_r_reg_19 (.CK( clk ) , .D( stage1_out_19 ) , .Q( u1_desIn_r_19 ) );
  DFF_X1 u1_desIn_r_reg_2 (.CK( clk ) , .D( stage1_out_2 ) , .Q( u1_desIn_r_2 ) );
  DFF_X1 u1_desIn_r_reg_20 (.CK( clk ) , .D( stage1_out_20 ) , .Q( u1_desIn_r_20 ) );
  DFF_X1 u1_desIn_r_reg_21 (.CK( clk ) , .D( stage1_out_21 ) , .Q( u1_desIn_r_21 ) );
  DFF_X1 u1_desIn_r_reg_22 (.CK( clk ) , .D( stage1_out_22 ) , .Q( u1_desIn_r_22 ) );
  DFF_X1 u1_desIn_r_reg_23 (.CK( clk ) , .D( stage1_out_23 ) , .Q( u1_desIn_r_23 ) );
  DFF_X1 u1_desIn_r_reg_24 (.CK( clk ) , .D( stage1_out_24 ) , .Q( u1_desIn_r_24 ) );
  DFF_X1 u1_desIn_r_reg_25 (.CK( clk ) , .D( stage1_out_25 ) , .Q( u1_desIn_r_25 ) );
  DFF_X1 u1_desIn_r_reg_26 (.CK( clk ) , .D( stage1_out_26 ) , .Q( u1_desIn_r_26 ) );
  DFF_X1 u1_desIn_r_reg_27 (.CK( clk ) , .D( stage1_out_27 ) , .Q( u1_desIn_r_27 ) );
  DFF_X1 u1_desIn_r_reg_28 (.CK( clk ) , .D( stage1_out_28 ) , .Q( u1_desIn_r_28 ) );
  DFF_X1 u1_desIn_r_reg_29 (.CK( clk ) , .D( stage1_out_29 ) , .Q( u1_desIn_r_29 ) );
  DFF_X1 u1_desIn_r_reg_3 (.CK( clk ) , .D( stage1_out_3 ) , .Q( u1_desIn_r_3 ) );
  DFF_X1 u1_desIn_r_reg_30 (.CK( clk ) , .D( stage1_out_30 ) , .Q( u1_desIn_r_30 ) );
  DFF_X1 u1_desIn_r_reg_31 (.CK( clk ) , .D( stage1_out_31 ) , .Q( u1_desIn_r_31 ) );
  DFF_X1 u1_desIn_r_reg_32 (.CK( clk ) , .D( stage1_out_32 ) , .Q( u1_desIn_r_32 ) );
  DFF_X1 u1_desIn_r_reg_33 (.CK( clk ) , .D( stage1_out_33 ) , .Q( u1_desIn_r_33 ) );
  DFF_X1 u1_desIn_r_reg_34 (.CK( clk ) , .D( stage1_out_34 ) , .Q( u1_desIn_r_34 ) );
  DFF_X1 u1_desIn_r_reg_35 (.CK( clk ) , .D( stage1_out_35 ) , .Q( u1_desIn_r_35 ) );
  DFF_X1 u1_desIn_r_reg_36 (.CK( clk ) , .D( stage1_out_36 ) , .Q( u1_desIn_r_36 ) );
  DFF_X1 u1_desIn_r_reg_37 (.CK( clk ) , .D( stage1_out_37 ) , .Q( u1_desIn_r_37 ) );
  DFF_X1 u1_desIn_r_reg_38 (.CK( clk ) , .D( stage1_out_38 ) , .Q( u1_desIn_r_38 ) );
  DFF_X1 u1_desIn_r_reg_39 (.CK( clk ) , .D( stage1_out_39 ) , .Q( u1_desIn_r_39 ) );
  DFF_X1 u1_desIn_r_reg_4 (.CK( clk ) , .D( stage1_out_4 ) , .Q( u1_desIn_r_4 ) );
  DFF_X1 u1_desIn_r_reg_40 (.CK( clk ) , .D( stage1_out_40 ) , .Q( u1_desIn_r_40 ) );
  DFF_X1 u1_desIn_r_reg_41 (.CK( clk ) , .D( stage1_out_41 ) , .Q( u1_desIn_r_41 ) );
  DFF_X1 u1_desIn_r_reg_42 (.CK( clk ) , .D( stage1_out_42 ) , .Q( u1_desIn_r_42 ) );
  DFF_X1 u1_desIn_r_reg_43 (.CK( clk ) , .D( stage1_out_43 ) , .Q( u1_desIn_r_43 ) );
  DFF_X1 u1_desIn_r_reg_44 (.CK( clk ) , .D( stage1_out_44 ) , .Q( u1_desIn_r_44 ) );
  DFF_X1 u1_desIn_r_reg_45 (.CK( clk ) , .D( stage1_out_45 ) , .Q( u1_desIn_r_45 ) );
  DFF_X1 u1_desIn_r_reg_46 (.CK( clk ) , .D( stage1_out_46 ) , .Q( u1_desIn_r_46 ) );
  DFF_X1 u1_desIn_r_reg_47 (.CK( clk ) , .D( stage1_out_47 ) , .Q( u1_desIn_r_47 ) );
  DFF_X1 u1_desIn_r_reg_48 (.CK( clk ) , .D( stage1_out_48 ) , .Q( u1_desIn_r_48 ) );
  DFF_X1 u1_desIn_r_reg_49 (.CK( clk ) , .D( stage1_out_49 ) , .Q( u1_desIn_r_49 ) );
  DFF_X1 u1_desIn_r_reg_5 (.CK( clk ) , .D( stage1_out_5 ) , .Q( u1_desIn_r_5 ) );
  DFF_X1 u1_desIn_r_reg_50 (.CK( clk ) , .D( stage1_out_50 ) , .Q( u1_desIn_r_50 ) );
  DFF_X1 u1_desIn_r_reg_51 (.CK( clk ) , .D( stage1_out_51 ) , .Q( u1_desIn_r_51 ) );
  DFF_X1 u1_desIn_r_reg_52 (.CK( clk ) , .D( stage1_out_52 ) , .Q( u1_desIn_r_52 ) );
  DFF_X1 u1_desIn_r_reg_53 (.CK( clk ) , .D( stage1_out_53 ) , .Q( u1_desIn_r_53 ) );
  DFF_X1 u1_desIn_r_reg_54 (.CK( clk ) , .D( stage1_out_54 ) , .Q( u1_desIn_r_54 ) );
  DFF_X1 u1_desIn_r_reg_55 (.CK( clk ) , .D( stage1_out_55 ) , .Q( u1_desIn_r_55 ) );
  DFF_X1 u1_desIn_r_reg_56 (.CK( clk ) , .D( stage1_out_56 ) , .Q( u1_desIn_r_56 ) );
  DFF_X1 u1_desIn_r_reg_57 (.CK( clk ) , .D( stage1_out_57 ) , .Q( u1_desIn_r_57 ) );
  DFF_X1 u1_desIn_r_reg_58 (.CK( clk ) , .D( stage1_out_58 ) , .Q( u1_desIn_r_58 ) );
  DFF_X1 u1_desIn_r_reg_59 (.CK( clk ) , .D( stage1_out_59 ) , .Q( u1_desIn_r_59 ) );
  DFF_X1 u1_desIn_r_reg_6 (.CK( clk ) , .D( stage1_out_6 ) , .Q( u1_desIn_r_6 ) );
  DFF_X1 u1_desIn_r_reg_60 (.CK( clk ) , .D( stage1_out_60 ) , .Q( u1_desIn_r_60 ) );
  DFF_X1 u1_desIn_r_reg_61 (.CK( clk ) , .D( stage1_out_61 ) , .Q( u1_desIn_r_61 ) );
  DFF_X1 u1_desIn_r_reg_62 (.CK( clk ) , .D( stage1_out_62 ) , .Q( u1_desIn_r_62 ) );
  DFF_X1 u1_desIn_r_reg_63 (.CK( clk ) , .D( stage1_out_63 ) , .Q( u1_desIn_r_63 ) );
  DFF_X1 u1_desIn_r_reg_7 (.CK( clk ) , .D( stage1_out_7 ) , .Q( u1_desIn_r_7 ) );
  DFF_X1 u1_desIn_r_reg_8 (.CK( clk ) , .D( stage1_out_8 ) , .Q( u1_desIn_r_8 ) );
  DFF_X1 u1_desIn_r_reg_9 (.CK( clk ) , .D( stage1_out_9 ) , .Q( u1_desIn_r_9 ) );
  DFF_X1 u1_desOut_reg_0 (.CK( clk ) , .Q( stage2_out_0 ) , .D( u1_FP_25 ) );
  DFF_X1 u1_desOut_reg_1 (.CK( clk ) , .Q( stage2_out_1 ) , .D( u1_FP_57 ) );
  DFF_X1 u1_desOut_reg_10 (.CK( clk ) , .Q( stage2_out_10 ) , .D( u1_FP_18 ) );
  DFF_X1 u1_desOut_reg_11 (.CK( clk ) , .Q( stage2_out_11 ) , .D( u1_FP_50 ) );
  DFF_X1 u1_desOut_reg_12 (.CK( clk ) , .Q( stage2_out_12 ) , .D( u1_FP_10 ) );
  DFF_X1 u1_desOut_reg_13 (.CK( clk ) , .Q( stage2_out_13 ) , .D( u1_FP_42 ) );
  DFF_X1 u1_desOut_reg_14 (.CK( clk ) , .Q( stage2_out_14 ) , .D( u1_FP_2 ) );
  DFF_X1 u1_desOut_reg_15 (.CK( clk ) , .Q( stage2_out_15 ) , .D( u1_FP_34 ) );
  DFF_X1 u1_desOut_reg_16 (.CK( clk ) , .Q( stage2_out_16 ) , .D( u1_FP_27 ) );
  DFF_X1 u1_desOut_reg_17 (.CK( clk ) , .Q( stage2_out_17 ) , .D( u1_FP_59 ) );
  DFF_X1 u1_desOut_reg_18 (.CK( clk ) , .Q( stage2_out_18 ) , .D( u1_FP_19 ) );
  DFF_X1 u1_desOut_reg_19 (.CK( clk ) , .Q( stage2_out_19 ) , .D( u1_FP_51 ) );
  DFF_X1 u1_desOut_reg_2 (.CK( clk ) , .Q( stage2_out_2 ) , .D( u1_FP_17 ) );
  DFF_X1 u1_desOut_reg_20 (.CK( clk ) , .Q( stage2_out_20 ) , .D( u1_FP_11 ) );
  DFF_X1 u1_desOut_reg_21 (.CK( clk ) , .Q( stage2_out_21 ) , .D( u1_FP_43 ) );
  DFF_X1 u1_desOut_reg_22 (.CK( clk ) , .Q( stage2_out_22 ) , .D( u1_FP_3 ) );
  DFF_X1 u1_desOut_reg_23 (.CK( clk ) , .Q( stage2_out_23 ) , .D( u1_FP_35 ) );
  DFF_X1 u1_desOut_reg_24 (.CK( clk ) , .Q( stage2_out_24 ) , .D( u1_FP_28 ) );
  DFF_X1 u1_desOut_reg_25 (.CK( clk ) , .Q( stage2_out_25 ) , .D( u1_FP_60 ) );
  DFF_X1 u1_desOut_reg_26 (.CK( clk ) , .Q( stage2_out_26 ) , .D( u1_FP_20 ) );
  DFF_X1 u1_desOut_reg_27 (.CK( clk ) , .Q( stage2_out_27 ) , .D( u1_FP_52 ) );
  DFF_X1 u1_desOut_reg_28 (.CK( clk ) , .Q( stage2_out_28 ) , .D( u1_FP_12 ) );
  DFF_X1 u1_desOut_reg_29 (.CK( clk ) , .Q( stage2_out_29 ) , .D( u1_FP_44 ) );
  DFF_X1 u1_desOut_reg_3 (.CK( clk ) , .Q( stage2_out_3 ) , .D( u1_FP_49 ) );
  DFF_X1 u1_desOut_reg_30 (.CK( clk ) , .Q( stage2_out_30 ) , .D( u1_FP_4 ) );
  DFF_X1 u1_desOut_reg_31 (.CK( clk ) , .Q( stage2_out_31 ) , .D( u1_FP_36 ) );
  DFF_X1 u1_desOut_reg_32 (.CK( clk ) , .Q( stage2_out_32 ) , .D( u1_FP_29 ) );
  DFF_X1 u1_desOut_reg_33 (.CK( clk ) , .Q( stage2_out_33 ) , .D( u1_FP_61 ) );
  DFF_X1 u1_desOut_reg_34 (.CK( clk ) , .Q( stage2_out_34 ) , .D( u1_FP_21 ) );
  DFF_X1 u1_desOut_reg_35 (.CK( clk ) , .Q( stage2_out_35 ) , .D( u1_FP_53 ) );
  DFF_X1 u1_desOut_reg_36 (.CK( clk ) , .Q( stage2_out_36 ) , .D( u1_FP_13 ) );
  DFF_X1 u1_desOut_reg_37 (.CK( clk ) , .Q( stage2_out_37 ) , .D( u1_FP_45 ) );
  DFF_X1 u1_desOut_reg_38 (.CK( clk ) , .Q( stage2_out_38 ) , .D( u1_FP_5 ) );
  DFF_X1 u1_desOut_reg_39 (.CK( clk ) , .Q( stage2_out_39 ) , .D( u1_FP_37 ) );
  DFF_X1 u1_desOut_reg_4 (.CK( clk ) , .Q( stage2_out_4 ) , .D( u1_FP_9 ) );
  DFF_X1 u1_desOut_reg_40 (.CK( clk ) , .Q( stage2_out_40 ) , .D( u1_FP_30 ) );
  DFF_X1 u1_desOut_reg_41 (.CK( clk ) , .Q( stage2_out_41 ) , .D( u1_FP_62 ) );
  DFF_X1 u1_desOut_reg_42 (.CK( clk ) , .Q( stage2_out_42 ) , .D( u1_FP_22 ) );
  DFF_X1 u1_desOut_reg_43 (.CK( clk ) , .Q( stage2_out_43 ) , .D( u1_FP_54 ) );
  DFF_X1 u1_desOut_reg_44 (.CK( clk ) , .Q( stage2_out_44 ) , .D( u1_FP_14 ) );
  DFF_X1 u1_desOut_reg_45 (.CK( clk ) , .Q( stage2_out_45 ) , .D( u1_FP_46 ) );
  DFF_X1 u1_desOut_reg_46 (.CK( clk ) , .Q( stage2_out_46 ) , .D( u1_FP_6 ) );
  DFF_X1 u1_desOut_reg_47 (.CK( clk ) , .Q( stage2_out_47 ) , .D( u1_FP_38 ) );
  DFF_X1 u1_desOut_reg_48 (.CK( clk ) , .Q( stage2_out_48 ) , .D( u1_FP_31 ) );
  DFF_X1 u1_desOut_reg_49 (.CK( clk ) , .Q( stage2_out_49 ) , .D( u1_FP_63 ) );
  DFF_X1 u1_desOut_reg_5 (.CK( clk ) , .Q( stage2_out_5 ) , .D( u1_FP_41 ) );
  DFF_X1 u1_desOut_reg_50 (.CK( clk ) , .Q( stage2_out_50 ) , .D( u1_FP_23 ) );
  DFF_X1 u1_desOut_reg_51 (.CK( clk ) , .Q( stage2_out_51 ) , .D( u1_FP_55 ) );
  DFF_X1 u1_desOut_reg_52 (.CK( clk ) , .Q( stage2_out_52 ) , .D( u1_FP_15 ) );
  DFF_X1 u1_desOut_reg_53 (.CK( clk ) , .Q( stage2_out_53 ) , .D( u1_FP_47 ) );
  DFF_X1 u1_desOut_reg_54 (.CK( clk ) , .Q( stage2_out_54 ) , .D( u1_FP_7 ) );
  DFF_X1 u1_desOut_reg_55 (.CK( clk ) , .Q( stage2_out_55 ) , .D( u1_FP_39 ) );
  DFF_X1 u1_desOut_reg_56 (.CK( clk ) , .Q( stage2_out_56 ) , .D( u1_FP_32 ) );
  DFF_X1 u1_desOut_reg_57 (.CK( clk ) , .Q( stage2_out_57 ) , .D( u1_FP_64 ) );
  DFF_X1 u1_desOut_reg_58 (.CK( clk ) , .Q( stage2_out_58 ) , .D( u1_FP_24 ) );
  DFF_X1 u1_desOut_reg_59 (.CK( clk ) , .Q( stage2_out_59 ) , .D( u1_FP_56 ) );
  DFF_X1 u1_desOut_reg_6 (.CK( clk ) , .Q( stage2_out_6 ) , .D( u1_FP_1 ) );
  DFF_X1 u1_desOut_reg_60 (.CK( clk ) , .Q( stage2_out_60 ) , .D( u1_FP_16 ) );
  DFF_X1 u1_desOut_reg_61 (.CK( clk ) , .Q( stage2_out_61 ) , .D( u1_FP_48 ) );
  DFF_X1 u1_desOut_reg_62 (.CK( clk ) , .Q( stage2_out_62 ) , .D( u1_FP_8 ) );
  DFF_X1 u1_desOut_reg_63 (.CK( clk ) , .Q( stage2_out_63 ) , .D( u1_FP_40 ) );
  DFF_X1 u1_desOut_reg_7 (.CK( clk ) , .Q( stage2_out_7 ) , .D( u1_FP_33 ) );
  DFF_X1 u1_desOut_reg_8 (.CK( clk ) , .Q( stage2_out_8 ) , .D( u1_FP_26 ) );
  DFF_X1 u1_desOut_reg_9 (.CK( clk ) , .Q( stage2_out_9 ) , .D( u1_FP_58 ) );
  DFF_X1 u1_key_r_reg_0 (.CK( clk ) , .D( key_b_r_16_0 ) , .Q( u1_key_r_0 ) );
  DFF_X1 u1_key_r_reg_1 (.CK( clk ) , .D( key_b_r_16_1 ) , .Q( u1_key_r_1 ) );
  DFF_X1 u1_key_r_reg_10 (.CK( clk ) , .D( key_b_r_16_10 ) , .Q( u1_key_r_10 ) );
  DFF_X1 u1_key_r_reg_11 (.CK( clk ) , .D( key_b_r_16_11 ) , .Q( u1_key_r_11 ) );
  DFF_X1 u1_key_r_reg_12 (.CK( clk ) , .D( key_b_r_16_12 ) , .Q( u1_key_r_12 ) );
  DFF_X1 u1_key_r_reg_13 (.CK( clk ) , .D( key_b_r_16_13 ) , .Q( u1_key_r_13 ) );
  DFF_X1 u1_key_r_reg_14 (.CK( clk ) , .D( key_b_r_16_14 ) , .Q( u1_key_r_14 ) );
  DFF_X1 u1_key_r_reg_15 (.CK( clk ) , .D( key_b_r_16_15 ) , .Q( u1_key_r_15 ) );
  DFF_X1 u1_key_r_reg_16 (.CK( clk ) , .D( key_b_r_16_16 ) , .Q( u1_key_r_16 ) );
  DFF_X1 u1_key_r_reg_17 (.CK( clk ) , .D( key_b_r_16_17 ) , .Q( u1_key_r_17 ) );
  DFF_X1 u1_key_r_reg_18 (.CK( clk ) , .D( key_b_r_16_18 ) , .Q( u1_key_r_18 ) );
  DFF_X1 u1_key_r_reg_19 (.CK( clk ) , .D( key_b_r_16_19 ) , .Q( u1_key_r_19 ) );
  DFF_X1 u1_key_r_reg_2 (.CK( clk ) , .D( key_b_r_16_2 ) , .Q( u1_key_r_2 ) );
  DFF_X1 u1_key_r_reg_20 (.CK( clk ) , .D( key_b_r_16_20 ) , .Q( u1_key_r_20 ) );
  DFF_X1 u1_key_r_reg_21 (.CK( clk ) , .D( key_b_r_16_21 ) , .Q( u1_key_r_21 ) );
  DFF_X1 u1_key_r_reg_22 (.CK( clk ) , .D( key_b_r_16_22 ) , .Q( u1_key_r_22 ) );
  DFF_X1 u1_key_r_reg_23 (.CK( clk ) , .D( key_b_r_16_23 ) , .Q( u1_key_r_23 ) );
  DFF_X1 u1_key_r_reg_24 (.CK( clk ) , .D( key_b_r_16_24 ) , .Q( u1_key_r_24 ) );
  DFF_X1 u1_key_r_reg_25 (.CK( clk ) , .D( key_b_r_16_25 ) , .Q( u1_key_r_25 ) );
  DFF_X1 u1_key_r_reg_26 (.CK( clk ) , .D( key_b_r_16_26 ) , .Q( u1_key_r_26 ) );
  DFF_X1 u1_key_r_reg_27 (.CK( clk ) , .D( key_b_r_16_27 ) , .Q( u1_key_r_27 ) );
  DFF_X1 u1_key_r_reg_28 (.CK( clk ) , .D( key_b_r_16_28 ) , .Q( u1_key_r_28 ) );
  DFF_X1 u1_key_r_reg_29 (.CK( clk ) , .D( key_b_r_16_29 ) , .Q( u1_key_r_29 ) );
  DFF_X1 u1_key_r_reg_3 (.CK( clk ) , .D( key_b_r_16_3 ) , .Q( u1_key_r_3 ) );
  DFF_X1 u1_key_r_reg_30 (.CK( clk ) , .D( key_b_r_16_30 ) , .Q( u1_key_r_30 ) );
  DFF_X1 u1_key_r_reg_31 (.CK( clk ) , .D( key_b_r_16_31 ) , .Q( u1_key_r_31 ) );
  DFF_X1 u1_key_r_reg_32 (.CK( clk ) , .D( key_b_r_16_32 ) , .Q( u1_key_r_32 ) );
  DFF_X1 u1_key_r_reg_33 (.CK( clk ) , .D( key_b_r_16_33 ) , .Q( u1_key_r_33 ) );
  DFF_X1 u1_key_r_reg_34 (.CK( clk ) , .D( key_b_r_16_34 ) , .Q( u1_key_r_34 ) );
  DFF_X1 u1_key_r_reg_35 (.CK( clk ) , .D( key_b_r_16_35 ) , .Q( u1_key_r_35 ) );
  DFF_X1 u1_key_r_reg_36 (.CK( clk ) , .D( key_b_r_16_36 ) , .Q( u1_key_r_36 ) );
  DFF_X1 u1_key_r_reg_37 (.CK( clk ) , .D( key_b_r_16_37 ) , .Q( u1_key_r_37 ) );
  DFF_X1 u1_key_r_reg_38 (.CK( clk ) , .D( key_b_r_16_38 ) , .Q( u1_key_r_38 ) );
  DFF_X1 u1_key_r_reg_39 (.CK( clk ) , .D( key_b_r_16_39 ) , .Q( u1_key_r_39 ) );
  DFF_X1 u1_key_r_reg_4 (.CK( clk ) , .D( key_b_r_16_4 ) , .Q( u1_key_r_4 ) );
  DFF_X1 u1_key_r_reg_40 (.CK( clk ) , .D( key_b_r_16_40 ) , .Q( u1_key_r_40 ) );
  DFF_X1 u1_key_r_reg_41 (.CK( clk ) , .D( key_b_r_16_41 ) , .Q( u1_key_r_41 ) );
  DFF_X1 u1_key_r_reg_42 (.CK( clk ) , .D( key_b_r_16_42 ) , .Q( u1_key_r_42 ) );
  DFF_X1 u1_key_r_reg_43 (.CK( clk ) , .D( key_b_r_16_43 ) , .Q( u1_key_r_43 ) );
  DFF_X1 u1_key_r_reg_44 (.CK( clk ) , .D( key_b_r_16_44 ) , .Q( u1_key_r_44 ) );
  DFF_X1 u1_key_r_reg_45 (.CK( clk ) , .D( key_b_r_16_45 ) , .Q( u1_key_r_45 ) );
  DFF_X1 u1_key_r_reg_46 (.CK( clk ) , .D( key_b_r_16_46 ) , .Q( u1_key_r_46 ) );
  DFF_X1 u1_key_r_reg_47 (.CK( clk ) , .D( key_b_r_16_47 ) , .Q( u1_key_r_47 ) );
  DFF_X1 u1_key_r_reg_48 (.CK( clk ) , .D( key_b_r_16_48 ) , .Q( u1_key_r_48 ) );
  DFF_X1 u1_key_r_reg_49 (.CK( clk ) , .D( key_b_r_16_49 ) , .Q( u1_key_r_49 ) );
  DFF_X1 u1_key_r_reg_5 (.CK( clk ) , .D( key_b_r_16_5 ) , .Q( u1_key_r_5 ) );
  DFF_X1 u1_key_r_reg_50 (.CK( clk ) , .D( key_b_r_16_50 ) , .Q( u1_key_r_50 ) );
  DFF_X1 u1_key_r_reg_51 (.CK( clk ) , .D( key_b_r_16_51 ) , .Q( u1_key_r_51 ) );
  DFF_X1 u1_key_r_reg_52 (.CK( clk ) , .D( key_b_r_16_52 ) , .Q( u1_key_r_52 ) );
  DFF_X1 u1_key_r_reg_53 (.CK( clk ) , .D( key_b_r_16_53 ) , .Q( u1_key_r_53 ) );
  DFF_X1 u1_key_r_reg_54 (.CK( clk ) , .D( key_b_r_16_54 ) , .Q( u1_key_r_54 ) );
  DFF_X1 u1_key_r_reg_55 (.CK( clk ) , .D( key_b_r_16_55 ) , .Q( u1_key_r_55 ) );
  DFF_X1 u1_key_r_reg_6 (.CK( clk ) , .D( key_b_r_16_6 ) , .Q( u1_key_r_6 ) );
  DFF_X1 u1_key_r_reg_7 (.CK( clk ) , .D( key_b_r_16_7 ) , .Q( u1_key_r_7 ) );
  DFF_X1 u1_key_r_reg_8 (.CK( clk ) , .D( key_b_r_16_8 ) , .Q( u1_key_r_8 ) );
  DFF_X1 u1_key_r_reg_9 (.CK( clk ) , .D( key_b_r_16_9 ) , .Q( u1_key_r_9 ) );
  DFF_X1 u1_uk_K_r0_reg_0 (.CK( clk ) , .D( u1_key_r_0 ) , .Q( u1_uk_K_r0_0 ) , .QN( u1_uk_n1260 ) );
  DFF_X1 u1_uk_K_r0_reg_1 (.CK( clk ) , .D( u1_key_r_1 ) , .Q( u1_uk_K_r0_1 ) );
  DFF_X1 u1_uk_K_r0_reg_10 (.CK( clk ) , .D( u1_key_r_10 ) , .Q( u1_uk_K_r0_10 ) , .QN( u1_uk_n1268 ) );
  DFF_X1 u1_uk_K_r0_reg_11 (.CK( clk ) , .D( u1_key_r_11 ) , .Q( u1_uk_K_r0_11 ) );
  DFF_X1 u1_uk_K_r0_reg_12 (.CK( clk ) , .D( u1_key_r_12 ) , .Q( u1_uk_K_r0_12 ) , .QN( u1_uk_n1269 ) );
  DFF_X1 u1_uk_K_r0_reg_13 (.CK( clk ) , .D( u1_key_r_13 ) , .Q( u1_uk_K_r0_13 ) , .QN( u1_uk_n1270 ) );
  DFF_X1 u1_uk_K_r0_reg_14 (.CK( clk ) , .D( u1_key_r_14 ) , .Q( u1_uk_K_r0_14 ) , .QN( u1_uk_n1271 ) );
  DFF_X1 u1_uk_K_r0_reg_15 (.CK( clk ) , .D( u1_key_r_15 ) , .Q( u1_uk_K_r0_15 ) );
  DFF_X1 u1_uk_K_r0_reg_16 (.CK( clk ) , .D( u1_key_r_16 ) , .Q( u1_uk_K_r0_16 ) , .QN( u1_uk_n1272 ) );
  DFF_X1 u1_uk_K_r0_reg_17 (.CK( clk ) , .D( u1_key_r_17 ) , .Q( u1_uk_K_r0_17 ) );
  DFF_X1 u1_uk_K_r0_reg_18 (.CK( clk ) , .D( u1_key_r_18 ) , .Q( u1_uk_K_r0_18 ) , .QN( u1_uk_n1273 ) );
  DFF_X1 u1_uk_K_r0_reg_19 (.CK( clk ) , .D( u1_key_r_19 ) , .Q( u1_uk_K_r0_19 ) );
  DFF_X1 u1_uk_K_r0_reg_2 (.CK( clk ) , .D( u1_key_r_2 ) , .Q( u1_uk_K_r0_2 ) );
  DFF_X1 u1_uk_K_r0_reg_20 (.CK( clk ) , .D( u1_key_r_20 ) , .Q( u1_uk_K_r0_20 ) , .QN( u1_uk_n1274 ) );
  DFF_X1 u1_uk_K_r0_reg_21 (.CK( clk ) , .D( u1_key_r_21 ) , .Q( u1_uk_K_r0_21 ) , .QN( u1_uk_n1275 ) );
  DFF_X1 u1_uk_K_r0_reg_22 (.CK( clk ) , .D( u1_key_r_22 ) , .Q( u1_uk_K_r0_22 ) );
  DFF_X1 u1_uk_K_r0_reg_23 (.CK( clk ) , .D( u1_key_r_23 ) , .Q( u1_uk_K_r0_23 ) , .QN( u1_uk_n1276 ) );
  DFF_X1 u1_uk_K_r0_reg_24 (.CK( clk ) , .D( u1_key_r_24 ) , .Q( u1_uk_K_r0_24 ) , .QN( u1_uk_n1277 ) );
  DFF_X1 u1_uk_K_r0_reg_25 (.CK( clk ) , .D( u1_key_r_25 ) , .Q( u1_uk_K_r0_25 ) );
  DFF_X1 u1_uk_K_r0_reg_26 (.CK( clk ) , .D( u1_key_r_26 ) , .Q( u1_uk_K_r0_26 ) , .QN( u1_uk_n1278 ) );
  DFF_X1 u1_uk_K_r0_reg_27 (.CK( clk ) , .D( u1_key_r_27 ) , .Q( u1_uk_K_r0_27 ) , .QN( u1_uk_n1279 ) );
  DFF_X1 u1_uk_K_r0_reg_28 (.CK( clk ) , .D( u1_key_r_28 ) , .Q( u1_uk_K_r0_28 ) );
  DFF_X1 u1_uk_K_r0_reg_29 (.CK( clk ) , .D( u1_key_r_29 ) , .Q( u1_uk_K_r0_29 ) , .QN( u1_uk_n1281 ) );
  DFF_X1 u1_uk_K_r0_reg_3 (.CK( clk ) , .D( u1_key_r_3 ) , .Q( u1_uk_K_r0_3 ) , .QN( u1_uk_n1261 ) );
  DFF_X1 u1_uk_K_r0_reg_30 (.CK( clk ) , .D( u1_key_r_30 ) , .Q( u1_uk_K_r0_30 ) , .QN( u1_uk_n1282 ) );
  DFF_X1 u1_uk_K_r0_reg_31 (.CK( clk ) , .D( u1_key_r_31 ) , .Q( u1_uk_K_r0_31 ) );
  DFF_X1 u1_uk_K_r0_reg_32 (.CK( clk ) , .D( u1_key_r_32 ) , .Q( u1_uk_K_r0_32 ) );
  DFF_X1 u1_uk_K_r0_reg_33 (.CK( clk ) , .D( u1_key_r_33 ) , .Q( u1_uk_K_r0_33 ) , .QN( u1_uk_n1284 ) );
  DFF_X1 u1_uk_K_r0_reg_34 (.CK( clk ) , .D( u1_key_r_34 ) , .Q( u1_uk_K_r0_34 ) );
  DFF_X1 u1_uk_K_r0_reg_35 (.CK( clk ) , .D( u1_key_r_35 ) , .Q( u1_uk_K_r0_35 ) , .QN( u1_uk_n1286 ) );
  DFF_X1 u1_uk_K_r0_reg_36 (.CK( clk ) , .D( u1_key_r_36 ) , .Q( u1_uk_K_r0_36 ) );
  DFF_X1 u1_uk_K_r0_reg_37 (.CK( clk ) , .D( u1_key_r_37 ) , .Q( u1_uk_K_r0_37 ) , .QN( u1_uk_n1288 ) );
  DFF_X1 u1_uk_K_r0_reg_38 (.CK( clk ) , .D( u1_key_r_38 ) , .Q( u1_uk_K_r0_38 ) , .QN( u1_uk_n1289 ) );
  DFF_X1 u1_uk_K_r0_reg_39 (.CK( clk ) , .D( u1_key_r_39 ) , .Q( u1_uk_K_r0_39 ) , .QN( u1_uk_n1290 ) );
  DFF_X1 u1_uk_K_r0_reg_4 (.CK( clk ) , .D( u1_key_r_4 ) , .Q( u1_uk_K_r0_4 ) , .QN( u1_uk_n1262 ) );
  DFF_X1 u1_uk_K_r0_reg_40 (.CK( clk ) , .D( u1_key_r_40 ) , .Q( u1_uk_K_r0_40 ) , .QN( u1_uk_n1291 ) );
  DFF_X1 u1_uk_K_r0_reg_41 (.CK( clk ) , .D( u1_key_r_41 ) , .Q( u1_uk_K_r0_41 ) , .QN( u1_uk_n1292 ) );
  DFF_X1 u1_uk_K_r0_reg_42 (.CK( clk ) , .D( u1_key_r_42 ) , .Q( u1_uk_K_r0_42 ) , .QN( u1_uk_n1293 ) );
  DFF_X1 u1_uk_K_r0_reg_43 (.CK( clk ) , .D( u1_key_r_43 ) , .Q( u1_uk_K_r0_43 ) , .QN( u1_uk_n1294 ) );
  DFF_X1 u1_uk_K_r0_reg_44 (.CK( clk ) , .D( u1_key_r_44 ) , .Q( u1_uk_K_r0_44 ) , .QN( u1_uk_n1295 ) );
  DFF_X1 u1_uk_K_r0_reg_45 (.CK( clk ) , .D( u1_key_r_45 ) , .Q( u1_uk_K_r0_45 ) , .QN( u1_uk_n1296 ) );
  DFF_X1 u1_uk_K_r0_reg_46 (.CK( clk ) , .D( u1_key_r_46 ) , .Q( u1_uk_K_r0_46 ) , .QN( u1_uk_n1297 ) );
  DFF_X1 u1_uk_K_r0_reg_47 (.CK( clk ) , .D( u1_key_r_47 ) , .Q( u1_uk_K_r0_47 ) , .QN( u1_uk_n1299 ) );
  DFF_X1 u1_uk_K_r0_reg_48 (.CK( clk ) , .D( u1_key_r_48 ) , .Q( u1_uk_K_r0_48 ) , .QN( u1_uk_n1300 ) );
  DFF_X1 u1_uk_K_r0_reg_49 (.CK( clk ) , .D( u1_key_r_49 ) , .Q( u1_uk_K_r0_49 ) );
  DFF_X1 u1_uk_K_r0_reg_5 (.CK( clk ) , .D( u1_key_r_5 ) , .Q( u1_uk_K_r0_5 ) , .QN( u1_uk_n1263 ) );
  DFF_X1 u1_uk_K_r0_reg_50 (.CK( clk ) , .D( u1_key_r_50 ) , .Q( u1_uk_K_r0_50 ) , .QN( u1_uk_n1303 ) );
  DFF_X1 u1_uk_K_r0_reg_51 (.CK( clk ) , .D( u1_key_r_51 ) , .Q( u1_uk_K_r0_51 ) , .QN( u1_uk_n1304 ) );
  DFF_X1 u1_uk_K_r0_reg_52 (.CK( clk ) , .D( u1_key_r_52 ) , .Q( u1_uk_K_r0_52 ) );
  DFF_X1 u1_uk_K_r0_reg_53 (.CK( clk ) , .D( u1_key_r_53 ) , .Q( u1_uk_K_r0_53 ) );
  DFF_X1 u1_uk_K_r0_reg_54 (.CK( clk ) , .D( u1_key_r_54 ) , .Q( u1_uk_K_r0_54 ) , .QN( u1_uk_n1305 ) );
  DFF_X1 u1_uk_K_r0_reg_55 (.CK( clk ) , .D( u1_key_r_55 ) , .Q( u1_uk_K_r0_55 ) );
  DFF_X1 u1_uk_K_r0_reg_6 (.CK( clk ) , .D( u1_key_r_6 ) , .Q( u1_uk_K_r0_6 ) , .QN( u1_uk_n1264 ) );
  DFF_X1 u1_uk_K_r0_reg_7 (.CK( clk ) , .D( u1_key_r_7 ) , .Q( u1_uk_K_r0_7 ) , .QN( u1_uk_n1265 ) );
  DFF_X1 u1_uk_K_r0_reg_8 (.CK( clk ) , .D( u1_key_r_8 ) , .Q( u1_uk_K_r0_8 ) , .QN( u1_uk_n1266 ) );
  DFF_X1 u1_uk_K_r0_reg_9 (.CK( clk ) , .D( u1_key_r_9 ) , .Q( u1_uk_K_r0_9 ) , .QN( u1_uk_n1267 ) );
  DFF_X1 u1_uk_K_r10_reg_0 (.CK( clk ) , .Q( u1_uk_K_r10_0 ) , .D( u1_uk_K_r9_0 ) , .QN( u1_uk_n1708 ) );
  DFF_X1 u1_uk_K_r10_reg_1 (.CK( clk ) , .Q( u1_uk_K_r10_1 ) , .D( u1_uk_K_r9_1 ) , .QN( u1_uk_n1709 ) );
  DFF_X1 u1_uk_K_r10_reg_10 (.CK( clk ) , .Q( u1_uk_K_r10_10 ) , .D( u1_uk_K_r9_10 ) );
  DFF_X1 u1_uk_K_r10_reg_11 (.CK( clk ) , .Q( u1_uk_K_r10_11 ) , .D( u1_uk_K_r9_11 ) );
  DFF_X1 u1_uk_K_r10_reg_12 (.CK( clk ) , .Q( u1_uk_K_r10_12 ) , .D( u1_uk_K_r9_12 ) , .QN( u1_uk_n1716 ) );
  DFF_X1 u1_uk_K_r10_reg_13 (.CK( clk ) , .Q( u1_uk_K_r10_13 ) , .D( u1_uk_K_r9_13 ) );
  DFF_X1 u1_uk_K_r10_reg_14 (.CK( clk ) , .Q( u1_uk_K_r10_14 ) , .D( u1_uk_K_r9_14 ) );
  DFF_X1 u1_uk_K_r10_reg_15 (.CK( clk ) , .Q( u1_uk_K_r10_15 ) , .D( u1_uk_K_r9_15 ) , .QN( u1_uk_n1717 ) );
  DFF_X1 u1_uk_K_r10_reg_16 (.CK( clk ) , .Q( u1_uk_K_r10_16 ) , .D( u1_uk_K_r9_16 ) );
  DFF_X1 u1_uk_K_r10_reg_17 (.CK( clk ) , .Q( u1_uk_K_r10_17 ) , .D( u1_uk_K_r9_17 ) , .QN( u1_uk_n1718 ) );
  DFF_X1 u1_uk_K_r10_reg_18 (.CK( clk ) , .Q( u1_uk_K_r10_18 ) , .D( u1_uk_K_r9_18 ) );
  DFF_X1 u1_uk_K_r10_reg_19 (.CK( clk ) , .Q( u1_uk_K_r10_19 ) , .D( u1_uk_K_r9_19 ) );
  DFF_X1 u1_uk_K_r10_reg_2 (.CK( clk ) , .Q( u1_uk_K_r10_2 ) , .D( u1_uk_K_r9_2 ) , .QN( u1_uk_n1710 ) );
  DFF_X1 u1_uk_K_r10_reg_20 (.CK( clk ) , .Q( u1_uk_K_r10_20 ) , .D( u1_uk_K_r9_20 ) , .QN( u1_uk_n1719 ) );
  DFF_X1 u1_uk_K_r10_reg_21 (.CK( clk ) , .Q( u1_uk_K_r10_21 ) , .D( u1_uk_K_r9_21 ) , .QN( u1_uk_n1720 ) );
  DFF_X1 u1_uk_K_r10_reg_22 (.CK( clk ) , .Q( u1_uk_K_r10_22 ) , .D( u1_uk_K_r9_22 ) , .QN( u1_uk_n1721 ) );
  DFF_X1 u1_uk_K_r10_reg_23 (.CK( clk ) , .Q( u1_uk_K_r10_23 ) , .D( u1_uk_K_r9_23 ) );
  DFF_X1 u1_uk_K_r10_reg_24 (.CK( clk ) , .Q( u1_uk_K_r10_24 ) , .D( u1_uk_K_r9_24 ) , .QN( u1_uk_n1722 ) );
  DFF_X1 u1_uk_K_r10_reg_25 (.CK( clk ) , .Q( u1_uk_K_r10_25 ) , .D( u1_uk_K_r9_25 ) );
  DFF_X1 u1_uk_K_r10_reg_26 (.CK( clk ) , .Q( u1_uk_K_r10_26 ) , .D( u1_uk_K_r9_26 ) , .QN( u1_uk_n1723 ) );
  DFF_X1 u1_uk_K_r10_reg_27 (.CK( clk ) , .Q( u1_uk_K_r10_27 ) , .D( u1_uk_K_r9_27 ) );
  DFF_X1 u1_uk_K_r10_reg_28 (.CK( clk ) , .Q( u1_uk_K_r10_28 ) , .D( u1_uk_K_r9_28 ) );
  DFF_X1 u1_uk_K_r10_reg_29 (.CK( clk ) , .Q( u1_uk_K_r10_29 ) , .D( u1_uk_K_r9_29 ) , .QN( u1_uk_n1728 ) );
  DFF_X1 u1_uk_K_r10_reg_3 (.CK( clk ) , .Q( u1_uk_K_r10_3 ) , .D( u1_uk_K_r9_3 ) , .QN( u1_uk_n1711 ) );
  DFF_X1 u1_uk_K_r10_reg_30 (.CK( clk ) , .Q( u1_uk_K_r10_30 ) , .D( u1_uk_K_r9_30 ) , .QN( u1_uk_n1729 ) );
  DFF_X1 u1_uk_K_r10_reg_31 (.CK( clk ) , .Q( u1_uk_K_r10_31 ) , .D( u1_uk_K_r9_31 ) , .QN( u1_uk_n1730 ) );
  DFF_X1 u1_uk_K_r10_reg_32 (.CK( clk ) , .Q( u1_uk_K_r10_32 ) , .D( u1_uk_K_r9_32 ) , .QN( u1_uk_n1731 ) );
  DFF_X1 u1_uk_K_r10_reg_33 (.CK( clk ) , .Q( u1_uk_K_r10_33 ) , .D( u1_uk_K_r9_33 ) , .QN( u1_uk_n1732 ) );
  DFF_X1 u1_uk_K_r10_reg_34 (.CK( clk ) , .Q( u1_uk_K_r10_34 ) , .D( u1_uk_K_r9_34 ) );
  DFF_X1 u1_uk_K_r10_reg_35 (.CK( clk ) , .Q( u1_uk_K_r10_35 ) , .D( u1_uk_K_r9_35 ) , .QN( u1_uk_n1734 ) );
  DFF_X1 u1_uk_K_r10_reg_36 (.CK( clk ) , .Q( u1_uk_K_r10_36 ) , .D( u1_uk_K_r9_36 ) , .QN( u1_uk_n1735 ) );
  DFF_X1 u1_uk_K_r10_reg_37 (.CK( clk ) , .Q( u1_uk_K_r10_37 ) , .D( u1_uk_K_r9_37 ) , .QN( u1_uk_n1736 ) );
  DFF_X1 u1_uk_K_r10_reg_38 (.CK( clk ) , .Q( u1_uk_K_r10_38 ) , .D( u1_uk_K_r9_38 ) , .QN( u1_uk_n1737 ) );
  DFF_X1 u1_uk_K_r10_reg_39 (.CK( clk ) , .Q( u1_uk_K_r10_39 ) , .D( u1_uk_K_r9_39 ) , .QN( u1_uk_n1738 ) );
  DFF_X1 u1_uk_K_r10_reg_4 (.CK( clk ) , .Q( u1_uk_K_r10_4 ) , .D( u1_uk_K_r9_4 ) );
  DFF_X1 u1_uk_K_r10_reg_40 (.CK( clk ) , .Q( u1_uk_K_r10_40 ) , .D( u1_uk_K_r9_40 ) , .QN( u1_uk_n1739 ) );
  DFF_X1 u1_uk_K_r10_reg_41 (.CK( clk ) , .Q( u1_uk_K_r10_41 ) , .D( u1_uk_K_r9_41 ) );
  DFF_X1 u1_uk_K_r10_reg_42 (.CK( clk ) , .Q( u1_uk_K_r10_42 ) , .D( u1_uk_K_r9_42 ) );
  DFF_X1 u1_uk_K_r10_reg_43 (.CK( clk ) , .Q( u1_uk_K_r10_43 ) , .D( u1_uk_K_r9_43 ) );
  DFF_X1 u1_uk_K_r10_reg_44 (.CK( clk ) , .Q( u1_uk_K_r10_44 ) , .D( u1_uk_K_r9_44 ) );
  DFF_X1 u1_uk_K_r10_reg_45 (.CK( clk ) , .Q( u1_uk_K_r10_45 ) , .D( u1_uk_K_r9_45 ) , .QN( u1_uk_n1744 ) );
  DFF_X1 u1_uk_K_r10_reg_46 (.CK( clk ) , .Q( u1_uk_K_r10_46 ) , .D( u1_uk_K_r9_46 ) , .QN( u1_uk_n1745 ) );
  DFF_X1 u1_uk_K_r10_reg_47 (.CK( clk ) , .Q( u1_uk_K_r10_47 ) , .D( u1_uk_K_r9_47 ) );
  DFF_X1 u1_uk_K_r10_reg_48 (.CK( clk ) , .Q( u1_uk_K_r10_48 ) , .D( u1_uk_K_r9_48 ) );
  DFF_X1 u1_uk_K_r10_reg_49 (.CK( clk ) , .Q( u1_uk_K_r10_49 ) , .D( u1_uk_K_r9_49 ) );
  DFF_X1 u1_uk_K_r10_reg_5 (.CK( clk ) , .Q( u1_uk_K_r10_5 ) , .D( u1_uk_K_r9_5 ) , .QN( u1_uk_n1712 ) );
  DFF_X1 u1_uk_K_r10_reg_50 (.CK( clk ) , .Q( u1_uk_K_r10_50 ) , .D( u1_uk_K_r9_50 ) , .QN( u1_uk_n1748 ) );
  DFF_X1 u1_uk_K_r10_reg_51 (.CK( clk ) , .Q( u1_uk_K_r10_51 ) , .D( u1_uk_K_r9_51 ) , .QN( u1_uk_n1749 ) );
  DFF_X1 u1_uk_K_r10_reg_52 (.CK( clk ) , .Q( u1_uk_K_r10_52 ) , .D( u1_uk_K_r9_52 ) );
  DFF_X1 u1_uk_K_r10_reg_53 (.CK( clk ) , .Q( u1_uk_K_r10_53 ) , .D( u1_uk_K_r9_53 ) , .QN( u1_uk_n1750 ) );
  DFF_X1 u1_uk_K_r10_reg_54 (.CK( clk ) , .Q( u1_uk_K_r10_54 ) , .D( u1_uk_K_r9_54 ) , .QN( u1_uk_n1751 ) );
  DFF_X1 u1_uk_K_r10_reg_55 (.CK( clk ) , .Q( u1_uk_K_r10_55 ) , .D( u1_uk_K_r9_55 ) , .QN( u1_uk_n1752 ) );
  DFF_X1 u1_uk_K_r10_reg_6 (.CK( clk ) , .Q( u1_uk_K_r10_6 ) , .D( u1_uk_K_r9_6 ) , .QN( u1_uk_n1713 ) );
  DFF_X1 u1_uk_K_r10_reg_7 (.CK( clk ) , .Q( u1_uk_K_r10_7 ) , .D( u1_uk_K_r9_7 ) , .QN( u1_uk_n1714 ) );
  DFF_X1 u1_uk_K_r10_reg_8 (.CK( clk ) , .Q( u1_uk_K_r10_8 ) , .D( u1_uk_K_r9_8 ) , .QN( u1_uk_n1715 ) );
  DFF_X1 u1_uk_K_r10_reg_9 (.CK( clk ) , .Q( u1_uk_K_r10_9 ) , .D( u1_uk_K_r9_9 ) );
  DFF_X1 u1_uk_K_r11_reg_0 (.CK( clk ) , .D( u1_uk_K_r10_0 ) , .Q( u1_uk_K_r11_0 ) , .QN( u1_uk_n1753 ) );
  DFF_X1 u1_uk_K_r11_reg_1 (.CK( clk ) , .D( u1_uk_K_r10_1 ) , .Q( u1_uk_K_r11_1 ) , .QN( u1_uk_n1754 ) );
  DFF_X1 u1_uk_K_r11_reg_10 (.CK( clk ) , .D( u1_uk_K_r10_10 ) , .Q( u1_uk_K_r11_10 ) );
  DFF_X1 u1_uk_K_r11_reg_11 (.CK( clk ) , .D( u1_uk_K_r10_11 ) , .Q( u1_uk_K_r11_11 ) );
  DFF_X1 u1_uk_K_r11_reg_12 (.CK( clk ) , .D( u1_uk_K_r10_12 ) , .Q( u1_uk_K_r11_12 ) , .QN( u1_uk_n1761 ) );
  DFF_X1 u1_uk_K_r11_reg_13 (.CK( clk ) , .D( u1_uk_K_r10_13 ) , .Q( u1_uk_K_r11_13 ) , .QN( u1_uk_n1762 ) );
  DFF_X1 u1_uk_K_r11_reg_14 (.CK( clk ) , .D( u1_uk_K_r10_14 ) , .Q( u1_uk_K_r11_14 ) , .QN( u1_uk_n1763 ) );
  DFF_X1 u1_uk_K_r11_reg_15 (.CK( clk ) , .D( u1_uk_K_r10_15 ) , .Q( u1_uk_K_r11_15 ) , .QN( u1_uk_n1764 ) );
  DFF_X1 u1_uk_K_r11_reg_16 (.CK( clk ) , .D( u1_uk_K_r10_16 ) , .Q( u1_uk_K_r11_16 ) , .QN( u1_uk_n1765 ) );
  DFF_X1 u1_uk_K_r11_reg_17 (.CK( clk ) , .D( u1_uk_K_r10_17 ) , .Q( u1_uk_K_r11_17 ) , .QN( u1_uk_n1766 ) );
  DFF_X1 u1_uk_K_r11_reg_18 (.CK( clk ) , .D( u1_uk_K_r10_18 ) , .Q( u1_uk_K_r11_18 ) , .QN( u1_uk_n1767 ) );
  DFF_X1 u1_uk_K_r11_reg_19 (.CK( clk ) , .D( u1_uk_K_r10_19 ) , .Q( u1_uk_K_r11_19 ) );
  DFF_X1 u1_uk_K_r11_reg_2 (.CK( clk ) , .D( u1_uk_K_r10_2 ) , .Q( u1_uk_K_r11_2 ) , .QN( u1_uk_n1755 ) );
  DFF_X1 u1_uk_K_r11_reg_20 (.CK( clk ) , .D( u1_uk_K_r10_20 ) , .Q( u1_uk_K_r11_20 ) );
  DFF_X1 u1_uk_K_r11_reg_21 (.CK( clk ) , .D( u1_uk_K_r10_21 ) , .Q( u1_uk_K_r11_21 ) );
  DFF_X1 u1_uk_K_r11_reg_22 (.CK( clk ) , .D( u1_uk_K_r10_22 ) , .Q( u1_uk_K_r11_22 ) , .QN( u1_uk_n1768 ) );
  DFF_X1 u1_uk_K_r11_reg_23 (.CK( clk ) , .D( u1_uk_K_r10_23 ) , .Q( u1_uk_K_r11_23 ) , .QN( u1_uk_n1769 ) );
  DFF_X1 u1_uk_K_r11_reg_24 (.CK( clk ) , .D( u1_uk_K_r10_24 ) , .Q( u1_uk_K_r11_24 ) );
  DFF_X1 u1_uk_K_r11_reg_25 (.CK( clk ) , .D( u1_uk_K_r10_25 ) , .Q( u1_uk_K_r11_25 ) );
  DFF_X1 u1_uk_K_r11_reg_26 (.CK( clk ) , .D( u1_uk_K_r10_26 ) , .Q( u1_uk_K_r11_26 ) );
  DFF_X1 u1_uk_K_r11_reg_27 (.CK( clk ) , .D( u1_uk_K_r10_27 ) , .Q( u1_uk_K_r11_27 ) );
  DFF_X1 u1_uk_K_r11_reg_28 (.CK( clk ) , .D( u1_uk_K_r10_28 ) , .Q( u1_uk_K_r11_28 ) );
  DFF_X1 u1_uk_K_r11_reg_29 (.CK( clk ) , .D( u1_uk_K_r10_29 ) , .Q( u1_uk_K_r11_29 ) );
  DFF_X1 u1_uk_K_r11_reg_3 (.CK( clk ) , .D( u1_uk_K_r10_3 ) , .Q( u1_uk_K_r11_3 ) , .QN( u1_uk_n1756 ) );
  DFF_X1 u1_uk_K_r11_reg_30 (.CK( clk ) , .D( u1_uk_K_r10_30 ) , .Q( u1_uk_K_r11_30 ) );
  DFF_X1 u1_uk_K_r11_reg_31 (.CK( clk ) , .D( u1_uk_K_r10_31 ) , .Q( u1_uk_K_r11_31 ) , .QN( u1_uk_n1772 ) );
  DFF_X1 u1_uk_K_r11_reg_32 (.CK( clk ) , .D( u1_uk_K_r10_32 ) , .Q( u1_uk_K_r11_32 ) , .QN( u1_uk_n1773 ) );
  DFF_X1 u1_uk_K_r11_reg_33 (.CK( clk ) , .D( u1_uk_K_r10_33 ) , .Q( u1_uk_K_r11_33 ) );
  DFF_X1 u1_uk_K_r11_reg_34 (.CK( clk ) , .D( u1_uk_K_r10_34 ) , .Q( u1_uk_K_r11_34 ) );
  DFF_X1 u1_uk_K_r11_reg_35 (.CK( clk ) , .D( u1_uk_K_r10_35 ) , .Q( u1_uk_K_r11_35 ) , .QN( u1_uk_n1774 ) );
  DFF_X1 u1_uk_K_r11_reg_36 (.CK( clk ) , .D( u1_uk_K_r10_36 ) , .Q( u1_uk_K_r11_36 ) , .QN( u1_uk_n1775 ) );
  DFF_X1 u1_uk_K_r11_reg_37 (.CK( clk ) , .D( u1_uk_K_r10_37 ) , .Q( u1_uk_K_r11_37 ) , .QN( u1_uk_n1776 ) );
  DFF_X1 u1_uk_K_r11_reg_38 (.CK( clk ) , .D( u1_uk_K_r10_38 ) , .Q( u1_uk_K_r11_38 ) , .QN( u1_uk_n1777 ) );
  DFF_X1 u1_uk_K_r11_reg_39 (.CK( clk ) , .D( u1_uk_K_r10_39 ) , .Q( u1_uk_K_r11_39 ) );
  DFF_X1 u1_uk_K_r11_reg_4 (.CK( clk ) , .D( u1_uk_K_r10_4 ) , .Q( u1_uk_K_r11_4 ) );
  DFF_X1 u1_uk_K_r11_reg_40 (.CK( clk ) , .D( u1_uk_K_r10_40 ) , .Q( u1_uk_K_r11_40 ) , .QN( u1_uk_n1780 ) );
  DFF_X1 u1_uk_K_r11_reg_41 (.CK( clk ) , .D( u1_uk_K_r10_41 ) , .Q( u1_uk_K_r11_41 ) , .QN( u1_uk_n1781 ) );
  DFF_X1 u1_uk_K_r11_reg_42 (.CK( clk ) , .D( u1_uk_K_r10_42 ) , .Q( u1_uk_K_r11_42 ) , .QN( u1_uk_n1782 ) );
  DFF_X1 u1_uk_K_r11_reg_43 (.CK( clk ) , .D( u1_uk_K_r10_43 ) , .Q( u1_uk_K_r11_43 ) , .QN( u1_uk_n1783 ) );
  DFF_X1 u1_uk_K_r11_reg_44 (.CK( clk ) , .D( u1_uk_K_r10_44 ) , .Q( u1_uk_K_r11_44 ) , .QN( u1_uk_n1784 ) );
  DFF_X1 u1_uk_K_r11_reg_45 (.CK( clk ) , .D( u1_uk_K_r10_45 ) , .Q( u1_uk_K_r11_45 ) , .QN( u1_uk_n1785 ) );
  DFF_X1 u1_uk_K_r11_reg_46 (.CK( clk ) , .D( u1_uk_K_r10_46 ) , .Q( u1_uk_K_r11_46 ) , .QN( u1_uk_n1787 ) );
  DFF_X1 u1_uk_K_r11_reg_47 (.CK( clk ) , .D( u1_uk_K_r10_47 ) , .Q( u1_uk_K_r11_47 ) );
  DFF_X1 u1_uk_K_r11_reg_48 (.CK( clk ) , .D( u1_uk_K_r10_48 ) , .Q( u1_uk_K_r11_48 ) );
  DFF_X1 u1_uk_K_r11_reg_49 (.CK( clk ) , .D( u1_uk_K_r10_49 ) , .Q( u1_uk_K_r11_49 ) , .QN( u1_uk_n1790 ) );
  DFF_X1 u1_uk_K_r11_reg_5 (.CK( clk ) , .D( u1_uk_K_r10_5 ) , .Q( u1_uk_K_r11_5 ) , .QN( u1_uk_n1757 ) );
  DFF_X1 u1_uk_K_r11_reg_50 (.CK( clk ) , .D( u1_uk_K_r10_50 ) , .Q( u1_uk_K_r11_50 ) , .QN( u1_uk_n1791 ) );
  DFF_X1 u1_uk_K_r11_reg_51 (.CK( clk ) , .D( u1_uk_K_r10_51 ) , .Q( u1_uk_K_r11_51 ) , .QN( u1_uk_n1792 ) );
  DFF_X1 u1_uk_K_r11_reg_52 (.CK( clk ) , .D( u1_uk_K_r10_52 ) , .Q( u1_uk_K_r11_52 ) , .QN( u1_uk_n1793 ) );
  DFF_X1 u1_uk_K_r11_reg_53 (.CK( clk ) , .D( u1_uk_K_r10_53 ) , .Q( u1_uk_K_r11_53 ) );
  DFF_X1 u1_uk_K_r11_reg_54 (.CK( clk ) , .D( u1_uk_K_r10_54 ) , .Q( u1_uk_K_r11_54 ) );
  DFF_X1 u1_uk_K_r11_reg_55 (.CK( clk ) , .D( u1_uk_K_r10_55 ) , .Q( u1_uk_K_r11_55 ) , .QN( u1_uk_n1797 ) );
  DFF_X1 u1_uk_K_r11_reg_6 (.CK( clk ) , .D( u1_uk_K_r10_6 ) , .Q( u1_uk_K_r11_6 ) );
  DFF_X1 u1_uk_K_r11_reg_7 (.CK( clk ) , .D( u1_uk_K_r10_7 ) , .Q( u1_uk_K_r11_7 ) );
  DFF_X1 u1_uk_K_r11_reg_8 (.CK( clk ) , .D( u1_uk_K_r10_8 ) , .Q( u1_uk_K_r11_8 ) );
  DFF_X1 u1_uk_K_r11_reg_9 (.CK( clk ) , .D( u1_uk_K_r10_9 ) , .Q( u1_uk_K_r11_9 ) , .QN( u1_uk_n1758 ) );
  DFF_X1 u1_uk_K_r12_reg_0 (.CK( clk ) , .D( u1_uk_K_r11_0 ) , .Q( u1_uk_K_r12_0 ) , .QN( u1_uk_n1798 ) );
  DFF_X1 u1_uk_K_r12_reg_1 (.CK( clk ) , .D( u1_uk_K_r11_1 ) , .Q( u1_uk_K_r12_1 ) , .QN( u1_uk_n1799 ) );
  DFF_X1 u1_uk_K_r12_reg_10 (.CK( clk ) , .D( u1_uk_K_r11_10 ) , .Q( u1_uk_K_r12_10 ) );
  DFF_X1 u1_uk_K_r12_reg_11 (.CK( clk ) , .D( u1_uk_K_r11_11 ) , .Q( u1_uk_K_r12_11 ) , .QN( u1_uk_n1808 ) );
  DFF_X1 u1_uk_K_r12_reg_12 (.CK( clk ) , .D( u1_uk_K_r11_12 ) , .Q( u1_uk_K_r12_12 ) , .QN( u1_uk_n1809 ) );
  DFF_X1 u1_uk_K_r12_reg_13 (.CK( clk ) , .D( u1_uk_K_r11_13 ) , .Q( u1_uk_K_r12_13 ) , .QN( u1_uk_n1810 ) );
  DFF_X1 u1_uk_K_r12_reg_14 (.CK( clk ) , .D( u1_uk_K_r11_14 ) , .Q( u1_uk_K_r12_14 ) , .QN( u1_uk_n1811 ) );
  DFF_X1 u1_uk_K_r12_reg_15 (.CK( clk ) , .D( u1_uk_K_r11_15 ) , .Q( u1_uk_K_r12_15 ) );
  DFF_X1 u1_uk_K_r12_reg_16 (.CK( clk ) , .D( u1_uk_K_r11_16 ) , .Q( u1_uk_K_r12_16 ) );
  DFF_X1 u1_uk_K_r12_reg_17 (.CK( clk ) , .D( u1_uk_K_r11_17 ) , .Q( u1_uk_K_r12_17 ) , .QN( u1_uk_n1812 ) );
  DFF_X1 u1_uk_K_r12_reg_18 (.CK( clk ) , .D( u1_uk_K_r11_18 ) , .Q( u1_uk_K_r12_18 ) );
  DFF_X1 u1_uk_K_r12_reg_19 (.CK( clk ) , .D( u1_uk_K_r11_19 ) , .Q( u1_uk_K_r12_19 ) , .QN( u1_uk_n1813 ) );
  DFF_X1 u1_uk_K_r12_reg_2 (.CK( clk ) , .D( u1_uk_K_r11_2 ) , .Q( u1_uk_K_r12_2 ) , .QN( u1_uk_n1800 ) );
  DFF_X1 u1_uk_K_r12_reg_20 (.CK( clk ) , .D( u1_uk_K_r11_20 ) , .Q( u1_uk_K_r12_20 ) , .QN( u1_uk_n1814 ) );
  DFF_X1 u1_uk_K_r12_reg_21 (.CK( clk ) , .D( u1_uk_K_r11_21 ) , .Q( u1_uk_K_r12_21 ) );
  DFF_X1 u1_uk_K_r12_reg_22 (.CK( clk ) , .D( u1_uk_K_r11_22 ) , .Q( u1_uk_K_r12_22 ) );
  DFF_X1 u1_uk_K_r12_reg_23 (.CK( clk ) , .D( u1_uk_K_r11_23 ) , .Q( u1_uk_K_r12_23 ) , .QN( u1_uk_n1815 ) );
  DFF_X1 u1_uk_K_r12_reg_24 (.CK( clk ) , .D( u1_uk_K_r11_24 ) , .Q( u1_uk_K_r12_24 ) , .QN( u1_uk_n1816 ) );
  DFF_X1 u1_uk_K_r12_reg_25 (.CK( clk ) , .D( u1_uk_K_r11_25 ) , .Q( u1_uk_K_r12_25 ) , .QN( u1_uk_n1817 ) );
  DFF_X1 u1_uk_K_r12_reg_26 (.CK( clk ) , .D( u1_uk_K_r11_26 ) , .Q( u1_uk_K_r12_26 ) , .QN( u1_uk_n1818 ) );
  DFF_X1 u1_uk_K_r12_reg_27 (.CK( clk ) , .D( u1_uk_K_r11_27 ) , .Q( u1_uk_K_r12_27 ) , .QN( u1_uk_n1819 ) );
  DFF_X1 u1_uk_K_r12_reg_28 (.CK( clk ) , .D( u1_uk_K_r11_28 ) , .Q( u1_uk_K_r12_28 ) , .QN( u1_uk_n1820 ) );
  DFF_X1 u1_uk_K_r12_reg_29 (.CK( clk ) , .D( u1_uk_K_r11_29 ) , .Q( u1_uk_K_r12_29 ) , .QN( u1_uk_n1821 ) );
  DFF_X1 u1_uk_K_r12_reg_3 (.CK( clk ) , .D( u1_uk_K_r11_3 ) , .Q( u1_uk_K_r12_3 ) , .QN( u1_uk_n1801 ) );
  DFF_X1 u1_uk_K_r12_reg_30 (.CK( clk ) , .D( u1_uk_K_r11_30 ) , .Q( u1_uk_K_r12_30 ) , .QN( u1_uk_n1822 ) );
  DFF_X1 u1_uk_K_r12_reg_31 (.CK( clk ) , .D( u1_uk_K_r11_31 ) , .Q( u1_uk_K_r12_31 ) , .QN( u1_uk_n1823 ) );
  DFF_X1 u1_uk_K_r12_reg_32 (.CK( clk ) , .D( u1_uk_K_r11_32 ) , .Q( u1_uk_K_r12_32 ) , .QN( u1_uk_n1824 ) );
  DFF_X1 u1_uk_K_r12_reg_33 (.CK( clk ) , .D( u1_uk_K_r11_33 ) , .Q( u1_uk_K_r12_33 ) );
  DFF_X1 u1_uk_K_r12_reg_34 (.CK( clk ) , .D( u1_uk_K_r11_34 ) , .Q( u1_uk_K_r12_34 ) , .QN( u1_uk_n1826 ) );
  DFF_X1 u1_uk_K_r12_reg_35 (.CK( clk ) , .D( u1_uk_K_r11_35 ) , .Q( u1_uk_K_r12_35 ) , .QN( u1_uk_n1827 ) );
  DFF_X1 u1_uk_K_r12_reg_36 (.CK( clk ) , .D( u1_uk_K_r11_36 ) , .Q( u1_uk_K_r12_36 ) );
  DFF_X1 u1_uk_K_r12_reg_37 (.CK( clk ) , .D( u1_uk_K_r11_37 ) , .Q( u1_uk_K_r12_37 ) , .QN( u1_uk_n1829 ) );
  DFF_X1 u1_uk_K_r12_reg_38 (.CK( clk ) , .D( u1_uk_K_r11_38 ) , .Q( u1_uk_K_r12_38 ) , .QN( u1_uk_n1830 ) );
  DFF_X1 u1_uk_K_r12_reg_39 (.CK( clk ) , .D( u1_uk_K_r11_39 ) , .Q( u1_uk_K_r12_39 ) );
  DFF_X1 u1_uk_K_r12_reg_4 (.CK( clk ) , .D( u1_uk_K_r11_4 ) , .Q( u1_uk_K_r12_4 ) , .QN( u1_uk_n1802 ) );
  DFF_X1 u1_uk_K_r12_reg_40 (.CK( clk ) , .D( u1_uk_K_r11_40 ) , .Q( u1_uk_K_r12_40 ) , .QN( u1_uk_n1831 ) );
  DFF_X1 u1_uk_K_r12_reg_41 (.CK( clk ) , .D( u1_uk_K_r11_41 ) , .Q( u1_uk_K_r12_41 ) );
  DFF_X1 u1_uk_K_r12_reg_42 (.CK( clk ) , .D( u1_uk_K_r11_42 ) , .Q( u1_uk_K_r12_42 ) );
  DFF_X1 u1_uk_K_r12_reg_43 (.CK( clk ) , .D( u1_uk_K_r11_43 ) , .Q( u1_uk_K_r12_43 ) , .QN( u1_uk_n1832 ) );
  DFF_X1 u1_uk_K_r12_reg_44 (.CK( clk ) , .D( u1_uk_K_r11_44 ) , .Q( u1_uk_K_r12_44 ) );
  DFF_X1 u1_uk_K_r12_reg_45 (.CK( clk ) , .D( u1_uk_K_r11_45 ) , .Q( u1_uk_K_r12_45 ) , .QN( u1_uk_n1833 ) );
  DFF_X1 u1_uk_K_r12_reg_46 (.CK( clk ) , .D( u1_uk_K_r11_46 ) , .Q( u1_uk_K_r12_46 ) , .QN( u1_uk_n1834 ) );
  DFF_X1 u1_uk_K_r12_reg_47 (.CK( clk ) , .D( u1_uk_K_r11_47 ) , .Q( u1_uk_K_r12_47 ) );
  DFF_X1 u1_uk_K_r12_reg_48 (.CK( clk ) , .D( u1_uk_K_r11_48 ) , .Q( u1_uk_K_r12_48 ) , .QN( u1_uk_n1835 ) );
  DFF_X1 u1_uk_K_r12_reg_49 (.CK( clk ) , .D( u1_uk_K_r11_49 ) , .Q( u1_uk_K_r12_49 ) , .QN( u1_uk_n1836 ) );
  DFF_X1 u1_uk_K_r12_reg_5 (.CK( clk ) , .D( u1_uk_K_r11_5 ) , .Q( u1_uk_K_r12_5 ) , .QN( u1_uk_n1803 ) );
  DFF_X1 u1_uk_K_r12_reg_50 (.CK( clk ) , .D( u1_uk_K_r11_50 ) , .Q( u1_uk_K_r12_50 ) , .QN( u1_uk_n1837 ) );
  DFF_X1 u1_uk_K_r12_reg_51 (.CK( clk ) , .D( u1_uk_K_r11_51 ) , .Q( u1_uk_K_r12_51 ) , .QN( u1_uk_n1838 ) );
  DFF_X1 u1_uk_K_r12_reg_52 (.CK( clk ) , .D( u1_uk_K_r11_52 ) , .Q( u1_uk_K_r12_52 ) , .QN( u1_uk_n1839 ) );
  DFF_X1 u1_uk_K_r12_reg_53 (.CK( clk ) , .D( u1_uk_K_r11_53 ) , .Q( u1_uk_K_r12_53 ) , .QN( u1_uk_n1840 ) );
  DFF_X1 u1_uk_K_r12_reg_54 (.CK( clk ) , .D( u1_uk_K_r11_54 ) , .Q( u1_uk_K_r12_54 ) , .QN( u1_uk_n1841 ) );
  DFF_X1 u1_uk_K_r12_reg_55 (.CK( clk ) , .D( u1_uk_K_r11_55 ) , .Q( u1_uk_K_r12_55 ) , .QN( u1_uk_n1842 ) );
  DFF_X1 u1_uk_K_r12_reg_6 (.CK( clk ) , .D( u1_uk_K_r11_6 ) , .Q( u1_uk_K_r12_6 ) , .QN( u1_uk_n1804 ) );
  DFF_X1 u1_uk_K_r12_reg_7 (.CK( clk ) , .D( u1_uk_K_r11_7 ) , .Q( u1_uk_K_r12_7 ) );
  DFF_X1 u1_uk_K_r12_reg_8 (.CK( clk ) , .D( u1_uk_K_r11_8 ) , .Q( u1_uk_K_r12_8 ) , .QN( u1_uk_n1806 ) );
  DFF_X1 u1_uk_K_r12_reg_9 (.CK( clk ) , .D( u1_uk_K_r11_9 ) , .Q( u1_uk_K_r12_9 ) , .QN( u1_uk_n1807 ) );
  DFF_X1 u1_uk_K_r13_reg_0 (.CK( clk ) , .D( u1_uk_K_r12_0 ) , .Q( u1_uk_K_r13_0 ) , .QN( u1_uk_n1843 ) );
  DFF_X1 u1_uk_K_r13_reg_1 (.CK( clk ) , .D( u1_uk_K_r12_1 ) , .Q( u1_uk_K_r13_1 ) );
  DFF_X1 u1_uk_K_r13_reg_10 (.CK( clk ) , .D( u1_uk_K_r12_10 ) , .Q( u1_uk_K_r13_10 ) , .QN( u1_uk_n1850 ) );
  DFF_X1 u1_uk_K_r13_reg_11 (.CK( clk ) , .D( u1_uk_K_r12_11 ) , .Q( u1_uk_K_r13_11 ) , .QN( u1_uk_n1851 ) );
  DFF_X1 u1_uk_K_r13_reg_12 (.CK( clk ) , .D( u1_uk_K_r12_12 ) , .Q( u1_uk_K_r13_12 ) , .QN( u1_uk_n1852 ) );
  DFF_X1 u1_uk_K_r13_reg_13 (.CK( clk ) , .D( u1_uk_K_r12_13 ) , .Q( u1_uk_K_r13_13 ) , .QN( u1_uk_n1853 ) );
  DFF_X1 u1_uk_K_r13_reg_14 (.CK( clk ) , .D( u1_uk_K_r12_14 ) , .Q( u1_uk_K_r13_14 ) , .QN( u1_uk_n1854 ) );
  DFF_X1 u1_uk_K_r13_reg_15 (.CK( clk ) , .D( u1_uk_K_r12_15 ) , .Q( u1_uk_K_r13_15 ) , .QN( u1_uk_n1855 ) );
  DFF_X1 u1_uk_K_r13_reg_16 (.CK( clk ) , .D( u1_uk_K_r12_16 ) , .Q( u1_uk_K_r13_16 ) , .QN( u1_uk_n1856 ) );
  DFF_X1 u1_uk_K_r13_reg_17 (.CK( clk ) , .D( u1_uk_K_r12_17 ) , .Q( u1_uk_K_r13_17 ) );
  DFF_X1 u1_uk_K_r13_reg_18 (.CK( clk ) , .D( u1_uk_K_r12_18 ) , .Q( u1_uk_K_r13_18 ) , .QN( u1_uk_n1858 ) );
  DFF_X1 u1_uk_K_r13_reg_19 (.CK( clk ) , .D( u1_uk_K_r12_19 ) , .Q( u1_uk_K_r13_19 ) );
  DFF_X1 u1_uk_K_r13_reg_2 (.CK( clk ) , .D( u1_uk_K_r12_2 ) , .Q( u1_uk_K_r13_2 ) );
  DFF_X1 u1_uk_K_r13_reg_20 (.CK( clk ) , .D( u1_uk_K_r12_20 ) , .Q( u1_uk_K_r13_20 ) , .QN( u1_uk_n1859 ) );
  DFF_X1 u1_uk_K_r13_reg_21 (.CK( clk ) , .D( u1_uk_K_r12_21 ) , .Q( u1_uk_K_r13_21 ) , .QN( u1_uk_n1860 ) );
  DFF_X1 u1_uk_K_r13_reg_22 (.CK( clk ) , .D( u1_uk_K_r12_22 ) , .Q( u1_uk_K_r13_22 ) );
  DFF_X1 u1_uk_K_r13_reg_23 (.CK( clk ) , .D( u1_uk_K_r12_23 ) , .Q( u1_uk_K_r13_23 ) );
  DFF_X1 u1_uk_K_r13_reg_24 (.CK( clk ) , .D( u1_uk_K_r12_24 ) , .Q( u1_uk_K_r13_24 ) , .QN( u1_uk_n1862 ) );
  DFF_X1 u1_uk_K_r13_reg_25 (.CK( clk ) , .D( u1_uk_K_r12_25 ) , .Q( u1_uk_K_r13_25 ) );
  DFF_X1 u1_uk_K_r13_reg_26 (.CK( clk ) , .D( u1_uk_K_r12_26 ) , .Q( u1_uk_K_r13_26 ) , .QN( u1_uk_n1863 ) );
  DFF_X1 u1_uk_K_r13_reg_27 (.CK( clk ) , .D( u1_uk_K_r12_27 ) , .Q( u1_uk_K_r13_27 ) , .QN( u1_uk_n1864 ) );
  DFF_X1 u1_uk_K_r13_reg_28 (.CK( clk ) , .D( u1_uk_K_r12_28 ) , .Q( u1_uk_K_r13_28 ) , .QN( u1_uk_n1865 ) );
  DFF_X1 u1_uk_K_r13_reg_29 (.CK( clk ) , .D( u1_uk_K_r12_29 ) , .Q( u1_uk_K_r13_29 ) , .QN( u1_uk_n1866 ) );
  DFF_X1 u1_uk_K_r13_reg_3 (.CK( clk ) , .D( u1_uk_K_r12_3 ) , .Q( u1_uk_K_r13_3 ) , .QN( u1_uk_n1844 ) );
  DFF_X1 u1_uk_K_r13_reg_30 (.CK( clk ) , .D( u1_uk_K_r12_30 ) , .Q( u1_uk_K_r13_30 ) , .QN( u1_uk_n1867 ) );
  DFF_X1 u1_uk_K_r13_reg_31 (.CK( clk ) , .D( u1_uk_K_r12_31 ) , .Q( u1_uk_K_r13_31 ) );
  DFF_X1 u1_uk_K_r13_reg_32 (.CK( clk ) , .D( u1_uk_K_r12_32 ) , .Q( u1_uk_K_r13_32 ) );
  DFF_X1 u1_uk_K_r13_reg_33 (.CK( clk ) , .D( u1_uk_K_r12_33 ) , .Q( u1_uk_K_r13_33 ) , .QN( u1_uk_n1868 ) );
  DFF_X1 u1_uk_K_r13_reg_34 (.CK( clk ) , .D( u1_uk_K_r12_34 ) , .Q( u1_uk_K_r13_34 ) , .QN( u1_uk_n1869 ) );
  DFF_X1 u1_uk_K_r13_reg_35 (.CK( clk ) , .D( u1_uk_K_r12_35 ) , .Q( u1_uk_K_r13_35 ) );
  DFF_X1 u1_uk_K_r13_reg_36 (.CK( clk ) , .D( u1_uk_K_r12_36 ) , .Q( u1_uk_K_r13_36 ) );
  DFF_X1 u1_uk_K_r13_reg_37 (.CK( clk ) , .D( u1_uk_K_r12_37 ) , .Q( u1_uk_K_r13_37 ) , .QN( u1_uk_n1870 ) );
  DFF_X1 u1_uk_K_r13_reg_38 (.CK( clk ) , .D( u1_uk_K_r12_38 ) , .Q( u1_uk_K_r13_38 ) );
  DFF_X1 u1_uk_K_r13_reg_39 (.CK( clk ) , .D( u1_uk_K_r12_39 ) , .Q( u1_uk_K_r13_39 ) , .QN( u1_uk_n1872 ) );
  DFF_X1 u1_uk_K_r13_reg_4 (.CK( clk ) , .D( u1_uk_K_r12_4 ) , .Q( u1_uk_K_r13_4 ) );
  DFF_X1 u1_uk_K_r13_reg_40 (.CK( clk ) , .D( u1_uk_K_r12_40 ) , .Q( u1_uk_K_r13_40 ) , .QN( u1_uk_n1873 ) );
  DFF_X1 u1_uk_K_r13_reg_41 (.CK( clk ) , .D( u1_uk_K_r12_41 ) , .Q( u1_uk_K_r13_41 ) , .QN( u1_uk_n1874 ) );
  DFF_X1 u1_uk_K_r13_reg_42 (.CK( clk ) , .D( u1_uk_K_r12_42 ) , .Q( u1_uk_K_r13_42 ) , .QN( u1_uk_n1875 ) );
  DFF_X1 u1_uk_K_r13_reg_43 (.CK( clk ) , .D( u1_uk_K_r12_43 ) , .Q( u1_uk_K_r13_43 ) , .QN( u1_uk_n1876 ) );
  DFF_X1 u1_uk_K_r13_reg_44 (.CK( clk ) , .D( u1_uk_K_r12_44 ) , .Q( u1_uk_K_r13_44 ) );
  DFF_X1 u1_uk_K_r13_reg_45 (.CK( clk ) , .D( u1_uk_K_r12_45 ) , .Q( u1_uk_K_r13_45 ) , .QN( u1_uk_n1879 ) );
  DFF_X1 u1_uk_K_r13_reg_46 (.CK( clk ) , .D( u1_uk_K_r12_46 ) , .Q( u1_uk_K_r13_46 ) , .QN( u1_uk_n1880 ) );
  DFF_X1 u1_uk_K_r13_reg_47 (.CK( clk ) , .D( u1_uk_K_r12_47 ) , .Q( u1_uk_K_r13_47 ) , .QN( u1_uk_n1881 ) );
  DFF_X1 u1_uk_K_r13_reg_48 (.CK( clk ) , .D( u1_uk_K_r12_48 ) , .Q( u1_uk_K_r13_48 ) , .QN( u1_uk_n1882 ) );
  DFF_X1 u1_uk_K_r13_reg_49 (.CK( clk ) , .D( u1_uk_K_r12_49 ) , .Q( u1_uk_K_r13_49 ) , .QN( u1_uk_n1883 ) );
  DFF_X1 u1_uk_K_r13_reg_5 (.CK( clk ) , .D( u1_uk_K_r12_5 ) , .Q( u1_uk_K_r13_5 ) , .QN( u1_uk_n1845 ) );
  DFF_X1 u1_uk_K_r13_reg_50 (.CK( clk ) , .D( u1_uk_K_r12_50 ) , .Q( u1_uk_K_r13_50 ) , .QN( u1_uk_n1884 ) );
  DFF_X1 u1_uk_K_r13_reg_51 (.CK( clk ) , .D( u1_uk_K_r12_51 ) , .Q( u1_uk_K_r13_51 ) , .QN( u1_uk_n1885 ) );
  DFF_X1 u1_uk_K_r13_reg_52 (.CK( clk ) , .D( u1_uk_K_r12_52 ) , .Q( u1_uk_K_r13_52 ) , .QN( u1_uk_n1886 ) );
  DFF_X1 u1_uk_K_r13_reg_53 (.CK( clk ) , .D( u1_uk_K_r12_53 ) , .Q( u1_uk_K_r13_53 ) );
  DFF_X1 u1_uk_K_r13_reg_54 (.CK( clk ) , .D( u1_uk_K_r12_54 ) , .Q( u1_uk_K_r13_54 ) , .QN( u1_uk_n1887 ) );
  DFF_X1 u1_uk_K_r13_reg_55 (.CK( clk ) , .D( u1_uk_K_r12_55 ) , .Q( u1_uk_K_r13_55 ) );
  DFF_X1 u1_uk_K_r13_reg_6 (.CK( clk ) , .D( u1_uk_K_r12_6 ) , .Q( u1_uk_K_r13_6 ) , .QN( u1_uk_n1846 ) );
  DFF_X1 u1_uk_K_r13_reg_7 (.CK( clk ) , .D( u1_uk_K_r12_7 ) , .Q( u1_uk_K_r13_7 ) , .QN( u1_uk_n1847 ) );
  DFF_X1 u1_uk_K_r13_reg_8 (.CK( clk ) , .D( u1_uk_K_r12_8 ) , .Q( u1_uk_K_r13_8 ) , .QN( u1_uk_n1848 ) );
  DFF_X1 u1_uk_K_r13_reg_9 (.CK( clk ) , .D( u1_uk_K_r12_9 ) , .Q( u1_uk_K_r13_9 ) , .QN( u1_uk_n1849 ) );
  DFF_X1 u1_uk_K_r14_reg_0 (.CK( clk ) , .D( u1_uk_K_r13_0 ) , .QN( u1_uk_n1218 ) );
  DFF_X1 u1_uk_K_r14_reg_1 (.CK( clk ) , .D( u1_uk_K_r13_1 ) , .QN( u1_uk_n1219 ) );
  DFF_X1 u1_uk_K_r14_reg_10 (.CK( clk ) , .D( u1_uk_K_r13_10 ) , .Q( u1_uk_K_r14_10 ) );
  DFF_X1 u1_uk_K_r14_reg_11 (.CK( clk ) , .D( u1_uk_K_r13_11 ) , .Q( u1_uk_K_r14_11 ) );
  DFF_X1 u1_uk_K_r14_reg_12 (.CK( clk ) , .D( u1_uk_K_r13_12 ) , .Q( u1_uk_K_r14_12 ) );
  DFF_X1 u1_uk_K_r14_reg_13 (.CK( clk ) , .D( u1_uk_K_r13_13 ) , .QN( u1_uk_n1224 ) );
  DFF_X1 u1_uk_K_r14_reg_14 (.CK( clk ) , .D( u1_uk_K_r13_14 ) , .QN( u1_uk_n1225 ) );
  DFF_X1 u1_uk_K_r14_reg_15 (.CK( clk ) , .D( u1_uk_K_r13_15 ) , .Q( u1_uk_K_r14_15 ) );
  DFF_X1 u1_uk_K_r14_reg_16 (.CK( clk ) , .D( u1_uk_K_r13_16 ) , .Q( u1_uk_K_r14_16 ) );
  DFF_X1 u1_uk_K_r14_reg_17 (.CK( clk ) , .D( u1_uk_K_r13_17 ) , .QN( u1_uk_n1227 ) );
  DFF_X1 u1_uk_K_r14_reg_18 (.CK( clk ) , .D( u1_uk_K_r13_18 ) , .Q( u1_uk_K_r14_18 ) );
  DFF_X1 u1_uk_K_r14_reg_19 (.CK( clk ) , .D( u1_uk_K_r13_19 ) , .QN( u1_uk_n1228 ) );
  DFF_X1 u1_uk_K_r14_reg_2 (.CK( clk ) , .D( u1_uk_K_r13_2 ) , .Q( u1_uk_K_r14_2 ) );
  DFF_X1 u1_uk_K_r14_reg_20 (.CK( clk ) , .D( u1_uk_K_r13_20 ) , .QN( u1_uk_n1229 ) );
  DFF_X1 u1_uk_K_r14_reg_21 (.CK( clk ) , .D( u1_uk_K_r13_21 ) , .QN( u1_uk_n1230 ) );
  DFF_X1 u1_uk_K_r14_reg_22 (.CK( clk ) , .D( u1_uk_K_r13_22 ) , .QN( u1_uk_n1231 ) );
  DFF_X1 u1_uk_K_r14_reg_23 (.CK( clk ) , .D( u1_uk_K_r13_23 ) , .Q( u1_uk_K_r14_23 ) , .QN( u1_uk_n1233 ) );
  DFF_X1 u1_uk_K_r14_reg_24 (.CK( clk ) , .D( u1_uk_K_r13_24 ) , .QN( u1_uk_n1234 ) );
  DFF_X1 u1_uk_K_r14_reg_25 (.CK( clk ) , .D( u1_uk_K_r13_25 ) , .QN( u1_uk_n1235 ) );
  DFF_X1 u1_uk_K_r14_reg_26 (.CK( clk ) , .D( u1_uk_K_r13_26 ) , .QN( u1_uk_n1236 ) );
  DFF_X1 u1_uk_K_r14_reg_27 (.CK( clk ) , .D( u1_uk_K_r13_27 ) , .QN( u1_uk_n1237 ) );
  DFF_X1 u1_uk_K_r14_reg_28 (.CK( clk ) , .D( u1_uk_K_r13_28 ) , .QN( u1_uk_n1238 ) );
  DFF_X1 u1_uk_K_r14_reg_29 (.CK( clk ) , .D( u1_uk_K_r13_29 ) , .QN( u1_uk_n1239 ) );
  DFF_X1 u1_uk_K_r14_reg_3 (.CK( clk ) , .D( u1_uk_K_r13_3 ) , .Q( u1_uk_K_r14_3 ) );
  DFF_X1 u1_uk_K_r14_reg_30 (.CK( clk ) , .D( u1_uk_K_r13_30 ) , .QN( u1_uk_n1240 ) );
  DFF_X1 u1_uk_K_r14_reg_31 (.CK( clk ) , .D( u1_uk_K_r13_31 ) , .QN( u1_uk_n1241 ) );
  DFF_X1 u1_uk_K_r14_reg_32 (.CK( clk ) , .D( u1_uk_K_r13_32 ) , .QN( u1_uk_n1242 ) );
  DFF_X1 u1_uk_K_r14_reg_33 (.CK( clk ) , .D( u1_uk_K_r13_33 ) , .QN( u1_uk_n1243 ) );
  DFF_X1 u1_uk_K_r14_reg_34 (.CK( clk ) , .D( u1_uk_K_r13_34 ) , .QN( u1_uk_n1244 ) );
  DFF_X1 u1_uk_K_r14_reg_35 (.CK( clk ) , .D( u1_uk_K_r13_35 ) , .QN( u1_uk_n1245 ) );
  DFF_X1 u1_uk_K_r14_reg_36 (.CK( clk ) , .D( u1_uk_K_r13_36 ) , .QN( u1_uk_n1246 ) );
  DFF_X1 u1_uk_K_r14_reg_37 (.CK( clk ) , .D( u1_uk_K_r13_37 ) , .QN( u1_uk_n1247 ) );
  DFF_X1 u1_uk_K_r14_reg_38 (.CK( clk ) , .D( u1_uk_K_r13_38 ) , .Q( u1_uk_K_r14_38 ) );
  DFF_X1 u1_uk_K_r14_reg_39 (.CK( clk ) , .D( u1_uk_K_r13_39 ) , .Q( u1_uk_K_r14_39 ) );
  DFF_X1 u1_uk_K_r14_reg_4 (.CK( clk ) , .D( u1_uk_K_r13_4 ) , .QN( u1_uk_n1220 ) );
  DFF_X1 u1_uk_K_r14_reg_40 (.CK( clk ) , .D( u1_uk_K_r13_40 ) , .QN( u1_uk_n1248 ) );
  DFF_X1 u1_uk_K_r14_reg_41 (.CK( clk ) , .D( u1_uk_K_r13_41 ) , .QN( u1_uk_n1249 ) );
  DFF_X1 u1_uk_K_r14_reg_42 (.CK( clk ) , .D( u1_uk_K_r13_42 ) , .Q( u1_uk_K_r14_42 ) );
  DFF_X1 u1_uk_K_r14_reg_43 (.CK( clk ) , .D( u1_uk_K_r13_43 ) , .Q( u1_uk_K_r14_43 ) );
  DFF_X1 u1_uk_K_r14_reg_44 (.CK( clk ) , .D( u1_uk_K_r13_44 ) , .QN( u1_uk_n1250 ) );
  DFF_X1 u1_uk_K_r14_reg_45 (.CK( clk ) , .D( u1_uk_K_r13_45 ) , .Q( u1_uk_K_r14_45 ) );
  DFF_X1 u1_uk_K_r14_reg_46 (.CK( clk ) , .D( u1_uk_K_r13_46 ) , .Q( u1_uk_K_r14_46 ) );
  DFF_X1 u1_uk_K_r14_reg_47 (.CK( clk ) , .D( u1_uk_K_r13_47 ) , .QN( u1_uk_n1251 ) );
  DFF_X1 u1_uk_K_r14_reg_48 (.CK( clk ) , .D( u1_uk_K_r13_48 ) , .QN( u1_uk_n1252 ) );
  DFF_X1 u1_uk_K_r14_reg_49 (.CK( clk ) , .D( u1_uk_K_r13_49 ) , .QN( u1_uk_n1253 ) );
  DFF_X1 u1_uk_K_r14_reg_5 (.CK( clk ) , .D( u1_uk_K_r13_5 ) , .Q( u1_uk_K_r14_5 ) );
  DFF_X1 u1_uk_K_r14_reg_50 (.CK( clk ) , .D( u1_uk_K_r13_50 ) , .Q( u1_uk_K_r14_50 ) );
  DFF_X1 u1_uk_K_r14_reg_51 (.CK( clk ) , .D( u1_uk_K_r13_51 ) , .QN( u1_uk_n1255 ) );
  DFF_X1 u1_uk_K_r14_reg_52 (.CK( clk ) , .D( u1_uk_K_r13_52 ) , .QN( u1_uk_n1256 ) );
  DFF_X1 u1_uk_K_r14_reg_53 (.CK( clk ) , .D( u1_uk_K_r13_53 ) , .QN( u1_uk_n1257 ) );
  DFF_X1 u1_uk_K_r14_reg_54 (.CK( clk ) , .D( u1_uk_K_r13_54 ) , .QN( u1_uk_n1258 ) );
  DFF_X1 u1_uk_K_r14_reg_55 (.CK( clk ) , .D( u1_uk_K_r13_55 ) , .QN( u1_uk_n1259 ) );
  DFF_X1 u1_uk_K_r14_reg_6 (.CK( clk ) , .D( u1_uk_K_r13_6 ) , .QN( u1_uk_n1221 ) );
  DFF_X1 u1_uk_K_r14_reg_7 (.CK( clk ) , .D( u1_uk_K_r13_7 ) , .QN( u1_uk_n1222 ) );
  DFF_X1 u1_uk_K_r14_reg_8 (.CK( clk ) , .D( u1_uk_K_r13_8 ) , .Q( u1_uk_K_r14_8 ) );
  DFF_X1 u1_uk_K_r14_reg_9 (.CK( clk ) , .D( u1_uk_K_r13_9 ) , .Q( u1_uk_K_r14_9 ) );
  DFF_X1 u1_uk_K_r1_reg_0 (.CK( clk ) , .D( u1_uk_K_r0_0 ) , .Q( u1_uk_K_r1_0 ) , .QN( u1_uk_n1307 ) );
  DFF_X1 u1_uk_K_r1_reg_1 (.CK( clk ) , .D( u1_uk_K_r0_1 ) , .Q( u1_uk_K_r1_1 ) , .QN( u1_uk_n1308 ) );
  DFF_X1 u1_uk_K_r1_reg_10 (.CK( clk ) , .D( u1_uk_K_r0_10 ) , .Q( u1_uk_K_r1_10 ) );
  DFF_X1 u1_uk_K_r1_reg_11 (.CK( clk ) , .D( u1_uk_K_r0_11 ) , .Q( u1_uk_K_r1_11 ) , .QN( u1_uk_n1315 ) );
  DFF_X1 u1_uk_K_r1_reg_12 (.CK( clk ) , .D( u1_uk_K_r0_12 ) , .Q( u1_uk_K_r1_12 ) , .QN( u1_uk_n1316 ) );
  DFF_X1 u1_uk_K_r1_reg_13 (.CK( clk ) , .D( u1_uk_K_r0_13 ) , .Q( u1_uk_K_r1_13 ) , .QN( u1_uk_n1317 ) );
  DFF_X1 u1_uk_K_r1_reg_14 (.CK( clk ) , .D( u1_uk_K_r0_14 ) , .Q( u1_uk_K_r1_14 ) , .QN( u1_uk_n1318 ) );
  DFF_X1 u1_uk_K_r1_reg_15 (.CK( clk ) , .D( u1_uk_K_r0_15 ) , .Q( u1_uk_K_r1_15 ) );
  DFF_X1 u1_uk_K_r1_reg_16 (.CK( clk ) , .D( u1_uk_K_r0_16 ) , .Q( u1_uk_K_r1_16 ) );
  DFF_X1 u1_uk_K_r1_reg_17 (.CK( clk ) , .D( u1_uk_K_r0_17 ) , .Q( u1_uk_K_r1_17 ) , .QN( u1_uk_n1319 ) );
  DFF_X1 u1_uk_K_r1_reg_18 (.CK( clk ) , .D( u1_uk_K_r0_18 ) , .Q( u1_uk_K_r1_18 ) );
  DFF_X1 u1_uk_K_r1_reg_19 (.CK( clk ) , .D( u1_uk_K_r0_19 ) , .Q( u1_uk_K_r1_19 ) , .QN( u1_uk_n1320 ) );
  DFF_X1 u1_uk_K_r1_reg_2 (.CK( clk ) , .D( u1_uk_K_r0_2 ) , .Q( u1_uk_K_r1_2 ) , .QN( u1_uk_n1309 ) );
  DFF_X1 u1_uk_K_r1_reg_20 (.CK( clk ) , .D( u1_uk_K_r0_20 ) , .Q( u1_uk_K_r1_20 ) , .QN( u1_uk_n1321 ) );
  DFF_X1 u1_uk_K_r1_reg_21 (.CK( clk ) , .D( u1_uk_K_r0_21 ) , .Q( u1_uk_K_r1_21 ) );
  DFF_X1 u1_uk_K_r1_reg_22 (.CK( clk ) , .D( u1_uk_K_r0_22 ) , .Q( u1_uk_K_r1_22 ) );
  DFF_X1 u1_uk_K_r1_reg_23 (.CK( clk ) , .D( u1_uk_K_r0_23 ) , .Q( u1_uk_K_r1_23 ) , .QN( u1_uk_n1322 ) );
  DFF_X1 u1_uk_K_r1_reg_24 (.CK( clk ) , .D( u1_uk_K_r0_24 ) , .Q( u1_uk_K_r1_24 ) , .QN( u1_uk_n1323 ) );
  DFF_X1 u1_uk_K_r1_reg_25 (.CK( clk ) , .D( u1_uk_K_r0_25 ) , .Q( u1_uk_K_r1_25 ) , .QN( u1_uk_n1324 ) );
  DFF_X1 u1_uk_K_r1_reg_26 (.CK( clk ) , .D( u1_uk_K_r0_26 ) , .Q( u1_uk_K_r1_26 ) , .QN( u1_uk_n1325 ) );
  DFF_X1 u1_uk_K_r1_reg_27 (.CK( clk ) , .D( u1_uk_K_r0_27 ) , .Q( u1_uk_K_r1_27 ) , .QN( u1_uk_n1326 ) );
  DFF_X1 u1_uk_K_r1_reg_28 (.CK( clk ) , .D( u1_uk_K_r0_28 ) , .Q( u1_uk_K_r1_28 ) , .QN( u1_uk_n1327 ) );
  DFF_X1 u1_uk_K_r1_reg_29 (.CK( clk ) , .D( u1_uk_K_r0_29 ) , .Q( u1_uk_K_r1_29 ) , .QN( u1_uk_n1328 ) );
  DFF_X1 u1_uk_K_r1_reg_3 (.CK( clk ) , .D( u1_uk_K_r0_3 ) , .Q( u1_uk_K_r1_3 ) , .QN( u1_uk_n1310 ) );
  DFF_X1 u1_uk_K_r1_reg_30 (.CK( clk ) , .D( u1_uk_K_r0_30 ) , .Q( u1_uk_K_r1_30 ) , .QN( u1_uk_n1329 ) );
  DFF_X1 u1_uk_K_r1_reg_31 (.CK( clk ) , .D( u1_uk_K_r0_31 ) , .Q( u1_uk_K_r1_31 ) , .QN( u1_uk_n1330 ) );
  DFF_X1 u1_uk_K_r1_reg_32 (.CK( clk ) , .D( u1_uk_K_r0_32 ) , .Q( u1_uk_K_r1_32 ) , .QN( u1_uk_n1331 ) );
  DFF_X1 u1_uk_K_r1_reg_33 (.CK( clk ) , .D( u1_uk_K_r0_33 ) , .Q( u1_uk_K_r1_33 ) );
  DFF_X1 u1_uk_K_r1_reg_34 (.CK( clk ) , .D( u1_uk_K_r0_34 ) , .Q( u1_uk_K_r1_34 ) , .QN( u1_uk_n1332 ) );
  DFF_X1 u1_uk_K_r1_reg_35 (.CK( clk ) , .D( u1_uk_K_r0_35 ) , .Q( u1_uk_K_r1_35 ) , .QN( u1_uk_n1333 ) );
  DFF_X1 u1_uk_K_r1_reg_36 (.CK( clk ) , .D( u1_uk_K_r0_36 ) , .Q( u1_uk_K_r1_36 ) );
  DFF_X1 u1_uk_K_r1_reg_37 (.CK( clk ) , .D( u1_uk_K_r0_37 ) , .Q( u1_uk_K_r1_37 ) , .QN( u1_uk_n1334 ) );
  DFF_X1 u1_uk_K_r1_reg_38 (.CK( clk ) , .D( u1_uk_K_r0_38 ) , .Q( u1_uk_K_r1_38 ) , .QN( u1_uk_n1335 ) );
  DFF_X1 u1_uk_K_r1_reg_39 (.CK( clk ) , .D( u1_uk_K_r0_39 ) , .Q( u1_uk_K_r1_39 ) );
  DFF_X1 u1_uk_K_r1_reg_4 (.CK( clk ) , .D( u1_uk_K_r0_4 ) , .Q( u1_uk_K_r1_4 ) , .QN( u1_uk_n1311 ) );
  DFF_X1 u1_uk_K_r1_reg_40 (.CK( clk ) , .D( u1_uk_K_r0_40 ) , .Q( u1_uk_K_r1_40 ) , .QN( u1_uk_n1336 ) );
  DFF_X1 u1_uk_K_r1_reg_41 (.CK( clk ) , .D( u1_uk_K_r0_41 ) , .Q( u1_uk_K_r1_41 ) );
  DFF_X1 u1_uk_K_r1_reg_42 (.CK( clk ) , .D( u1_uk_K_r0_42 ) , .Q( u1_uk_K_r1_42 ) );
  DFF_X1 u1_uk_K_r1_reg_43 (.CK( clk ) , .D( u1_uk_K_r0_43 ) , .Q( u1_uk_K_r1_43 ) , .QN( u1_uk_n1338 ) );
  DFF_X1 u1_uk_K_r1_reg_44 (.CK( clk ) , .D( u1_uk_K_r0_44 ) , .Q( u1_uk_K_r1_44 ) );
  DFF_X1 u1_uk_K_r1_reg_45 (.CK( clk ) , .D( u1_uk_K_r0_45 ) , .Q( u1_uk_K_r1_45 ) , .QN( u1_uk_n1339 ) );
  DFF_X1 u1_uk_K_r1_reg_46 (.CK( clk ) , .D( u1_uk_K_r0_46 ) , .Q( u1_uk_K_r1_46 ) , .QN( u1_uk_n1340 ) );
  DFF_X1 u1_uk_K_r1_reg_47 (.CK( clk ) , .D( u1_uk_K_r0_47 ) , .Q( u1_uk_K_r1_47 ) );
  DFF_X1 u1_uk_K_r1_reg_48 (.CK( clk ) , .D( u1_uk_K_r0_48 ) , .Q( u1_uk_K_r1_48 ) , .QN( u1_uk_n1341 ) );
  DFF_X1 u1_uk_K_r1_reg_49 (.CK( clk ) , .D( u1_uk_K_r0_49 ) , .Q( u1_uk_K_r1_49 ) , .QN( u1_uk_n1342 ) );
  DFF_X1 u1_uk_K_r1_reg_5 (.CK( clk ) , .D( u1_uk_K_r0_5 ) , .Q( u1_uk_K_r1_5 ) , .QN( u1_uk_n1312 ) );
  DFF_X1 u1_uk_K_r1_reg_50 (.CK( clk ) , .D( u1_uk_K_r0_50 ) , .Q( u1_uk_K_r1_50 ) , .QN( u1_uk_n1343 ) );
  DFF_X1 u1_uk_K_r1_reg_51 (.CK( clk ) , .D( u1_uk_K_r0_51 ) , .Q( u1_uk_K_r1_51 ) , .QN( u1_uk_n1344 ) );
  DFF_X1 u1_uk_K_r1_reg_52 (.CK( clk ) , .D( u1_uk_K_r0_52 ) , .Q( u1_uk_K_r1_52 ) , .QN( u1_uk_n1345 ) );
  DFF_X1 u1_uk_K_r1_reg_53 (.CK( clk ) , .D( u1_uk_K_r0_53 ) , .Q( u1_uk_K_r1_53 ) , .QN( u1_uk_n1346 ) );
  DFF_X1 u1_uk_K_r1_reg_54 (.CK( clk ) , .D( u1_uk_K_r0_54 ) , .Q( u1_uk_K_r1_54 ) , .QN( u1_uk_n1347 ) );
  DFF_X1 u1_uk_K_r1_reg_55 (.CK( clk ) , .D( u1_uk_K_r0_55 ) , .Q( u1_uk_K_r1_55 ) , .QN( u1_uk_n1348 ) );
  DFF_X1 u1_uk_K_r1_reg_6 (.CK( clk ) , .D( u1_uk_K_r0_6 ) , .Q( u1_uk_K_r1_6 ) );
  DFF_X1 u1_uk_K_r1_reg_7 (.CK( clk ) , .D( u1_uk_K_r0_7 ) , .Q( u1_uk_K_r1_7 ) );
  DFF_X1 u1_uk_K_r1_reg_8 (.CK( clk ) , .D( u1_uk_K_r0_8 ) , .Q( u1_uk_K_r1_8 ) , .QN( u1_uk_n1313 ) );
  DFF_X1 u1_uk_K_r1_reg_9 (.CK( clk ) , .D( u1_uk_K_r0_9 ) , .Q( u1_uk_K_r1_9 ) , .QN( u1_uk_n1314 ) );
  DFF_X1 u1_uk_K_r2_reg_0 (.CK( clk ) , .D( u1_uk_K_r1_0 ) , .Q( u1_uk_K_r2_0 ) , .QN( u1_uk_n1349 ) );
  DFF_X1 u1_uk_K_r2_reg_1 (.CK( clk ) , .D( u1_uk_K_r1_1 ) , .Q( u1_uk_K_r2_1 ) , .QN( u1_uk_n1350 ) );
  DFF_X1 u1_uk_K_r2_reg_10 (.CK( clk ) , .D( u1_uk_K_r1_10 ) , .Q( u1_uk_K_r2_10 ) , .QN( u1_uk_n1357 ) );
  DFF_X1 u1_uk_K_r2_reg_11 (.CK( clk ) , .D( u1_uk_K_r1_11 ) , .Q( u1_uk_K_r2_11 ) , .QN( u1_uk_n1358 ) );
  DFF_X1 u1_uk_K_r2_reg_12 (.CK( clk ) , .D( u1_uk_K_r1_12 ) , .Q( u1_uk_K_r2_12 ) , .QN( u1_uk_n1359 ) );
  DFF_X1 u1_uk_K_r2_reg_13 (.CK( clk ) , .D( u1_uk_K_r1_13 ) , .Q( u1_uk_K_r2_13 ) );
  DFF_X1 u1_uk_K_r2_reg_14 (.CK( clk ) , .D( u1_uk_K_r1_14 ) , .Q( u1_uk_K_r2_14 ) , .QN( u1_uk_n1360 ) );
  DFF_X1 u1_uk_K_r2_reg_15 (.CK( clk ) , .D( u1_uk_K_r1_15 ) , .Q( u1_uk_K_r2_15 ) , .QN( u1_uk_n1361 ) );
  DFF_X1 u1_uk_K_r2_reg_16 (.CK( clk ) , .D( u1_uk_K_r1_16 ) , .Q( u1_uk_K_r2_16 ) );
  DFF_X1 u1_uk_K_r2_reg_17 (.CK( clk ) , .D( u1_uk_K_r1_17 ) , .Q( u1_uk_K_r2_17 ) , .QN( u1_uk_n1363 ) );
  DFF_X1 u1_uk_K_r2_reg_18 (.CK( clk ) , .D( u1_uk_K_r1_18 ) , .Q( u1_uk_K_r2_18 ) );
  DFF_X1 u1_uk_K_r2_reg_19 (.CK( clk ) , .D( u1_uk_K_r1_19 ) , .Q( u1_uk_K_r2_19 ) , .QN( u1_uk_n1365 ) );
  DFF_X1 u1_uk_K_r2_reg_2 (.CK( clk ) , .D( u1_uk_K_r1_2 ) , .Q( u1_uk_K_r2_2 ) , .QN( u1_uk_n1351 ) );
  DFF_X1 u1_uk_K_r2_reg_20 (.CK( clk ) , .D( u1_uk_K_r1_20 ) , .Q( u1_uk_K_r2_20 ) );
  DFF_X1 u1_uk_K_r2_reg_21 (.CK( clk ) , .D( u1_uk_K_r1_21 ) , .Q( u1_uk_K_r2_21 ) );
  DFF_X1 u1_uk_K_r2_reg_22 (.CK( clk ) , .D( u1_uk_K_r1_22 ) , .Q( u1_uk_K_r2_22 ) , .QN( u1_uk_n1366 ) );
  DFF_X1 u1_uk_K_r2_reg_23 (.CK( clk ) , .D( u1_uk_K_r1_23 ) , .Q( u1_uk_K_r2_23 ) , .QN( u1_uk_n1367 ) );
  DFF_X1 u1_uk_K_r2_reg_24 (.CK( clk ) , .D( u1_uk_K_r1_24 ) , .Q( u1_uk_K_r2_24 ) );
  DFF_X1 u1_uk_K_r2_reg_25 (.CK( clk ) , .D( u1_uk_K_r1_25 ) , .Q( u1_uk_K_r2_25 ) );
  DFF_X1 u1_uk_K_r2_reg_26 (.CK( clk ) , .D( u1_uk_K_r1_26 ) , .Q( u1_uk_K_r2_26 ) );
  DFF_X1 u1_uk_K_r2_reg_27 (.CK( clk ) , .D( u1_uk_K_r1_27 ) , .Q( u1_uk_K_r2_27 ) );
  DFF_X1 u1_uk_K_r2_reg_28 (.CK( clk ) , .D( u1_uk_K_r1_28 ) , .Q( u1_uk_K_r2_28 ) );
  DFF_X1 u1_uk_K_r2_reg_29 (.CK( clk ) , .D( u1_uk_K_r1_29 ) , .Q( u1_uk_K_r2_29 ) );
  DFF_X1 u1_uk_K_r2_reg_3 (.CK( clk ) , .D( u1_uk_K_r1_3 ) , .Q( u1_uk_K_r2_3 ) , .QN( u1_uk_n1352 ) );
  DFF_X1 u1_uk_K_r2_reg_30 (.CK( clk ) , .D( u1_uk_K_r1_30 ) , .Q( u1_uk_K_r2_30 ) );
  DFF_X1 u1_uk_K_r2_reg_31 (.CK( clk ) , .D( u1_uk_K_r1_31 ) , .Q( u1_uk_K_r2_31 ) );
  DFF_X1 u1_uk_K_r2_reg_32 (.CK( clk ) , .D( u1_uk_K_r1_32 ) , .Q( u1_uk_K_r2_32 ) , .QN( u1_uk_n1369 ) );
  DFF_X1 u1_uk_K_r2_reg_33 (.CK( clk ) , .D( u1_uk_K_r1_33 ) , .Q( u1_uk_K_r2_33 ) );
  DFF_X1 u1_uk_K_r2_reg_34 (.CK( clk ) , .D( u1_uk_K_r1_34 ) , .Q( u1_uk_K_r2_34 ) , .QN( u1_uk_n1371 ) );
  DFF_X1 u1_uk_K_r2_reg_35 (.CK( clk ) , .D( u1_uk_K_r1_35 ) , .Q( u1_uk_K_r2_35 ) , .QN( u1_uk_n1372 ) );
  DFF_X1 u1_uk_K_r2_reg_36 (.CK( clk ) , .D( u1_uk_K_r1_36 ) , .Q( u1_uk_K_r2_36 ) , .QN( u1_uk_n1374 ) );
  DFF_X1 u1_uk_K_r2_reg_37 (.CK( clk ) , .D( u1_uk_K_r1_37 ) , .Q( u1_uk_K_r2_37 ) , .QN( u1_uk_n1375 ) );
  DFF_X1 u1_uk_K_r2_reg_38 (.CK( clk ) , .D( u1_uk_K_r1_38 ) , .Q( u1_uk_K_r2_38 ) , .QN( u1_uk_n1376 ) );
  DFF_X1 u1_uk_K_r2_reg_39 (.CK( clk ) , .D( u1_uk_K_r1_39 ) , .Q( u1_uk_K_r2_39 ) , .QN( u1_uk_n1377 ) );
  DFF_X1 u1_uk_K_r2_reg_4 (.CK( clk ) , .D( u1_uk_K_r1_4 ) , .Q( u1_uk_K_r2_4 ) );
  DFF_X1 u1_uk_K_r2_reg_40 (.CK( clk ) , .D( u1_uk_K_r1_40 ) , .Q( u1_uk_K_r2_40 ) , .QN( u1_uk_n1378 ) );
  DFF_X1 u1_uk_K_r2_reg_41 (.CK( clk ) , .D( u1_uk_K_r1_41 ) , .Q( u1_uk_K_r2_41 ) );
  DFF_X1 u1_uk_K_r2_reg_42 (.CK( clk ) , .D( u1_uk_K_r1_42 ) , .Q( u1_uk_K_r2_42 ) , .QN( u1_uk_n1380 ) );
  DFF_X1 u1_uk_K_r2_reg_43 (.CK( clk ) , .D( u1_uk_K_r1_43 ) , .Q( u1_uk_K_r2_43 ) , .QN( u1_uk_n1381 ) );
  DFF_X1 u1_uk_K_r2_reg_44 (.CK( clk ) , .D( u1_uk_K_r1_44 ) , .Q( u1_uk_K_r2_44 ) , .QN( u1_uk_n1382 ) );
  DFF_X1 u1_uk_K_r2_reg_45 (.CK( clk ) , .D( u1_uk_K_r1_45 ) , .Q( u1_uk_K_r2_45 ) , .QN( u1_uk_n1383 ) );
  DFF_X1 u1_uk_K_r2_reg_46 (.CK( clk ) , .D( u1_uk_K_r1_46 ) , .Q( u1_uk_K_r2_46 ) );
  DFF_X1 u1_uk_K_r2_reg_47 (.CK( clk ) , .D( u1_uk_K_r1_47 ) , .Q( u1_uk_K_r2_47 ) );
  DFF_X1 u1_uk_K_r2_reg_48 (.CK( clk ) , .D( u1_uk_K_r1_48 ) , .Q( u1_uk_K_r2_48 ) , .QN( u1_uk_n1386 ) );
  DFF_X1 u1_uk_K_r2_reg_49 (.CK( clk ) , .D( u1_uk_K_r1_49 ) , .Q( u1_uk_K_r2_49 ) );
  DFF_X1 u1_uk_K_r2_reg_5 (.CK( clk ) , .D( u1_uk_K_r1_5 ) , .Q( u1_uk_K_r2_5 ) , .QN( u1_uk_n1353 ) );
  DFF_X1 u1_uk_K_r2_reg_50 (.CK( clk ) , .D( u1_uk_K_r1_50 ) , .Q( u1_uk_K_r2_50 ) );
  DFF_X1 u1_uk_K_r2_reg_51 (.CK( clk ) , .D( u1_uk_K_r1_51 ) , .Q( u1_uk_K_r2_51 ) , .QN( u1_uk_n1389 ) );
  DFF_X1 u1_uk_K_r2_reg_52 (.CK( clk ) , .D( u1_uk_K_r1_52 ) , .Q( u1_uk_K_r2_52 ) , .QN( u1_uk_n1390 ) );
  DFF_X1 u1_uk_K_r2_reg_53 (.CK( clk ) , .D( u1_uk_K_r1_53 ) , .Q( u1_uk_K_r2_53 ) );
  DFF_X1 u1_uk_K_r2_reg_54 (.CK( clk ) , .D( u1_uk_K_r1_54 ) , .Q( u1_uk_K_r2_54 ) , .QN( u1_uk_n1391 ) );
  DFF_X1 u1_uk_K_r2_reg_55 (.CK( clk ) , .D( u1_uk_K_r1_55 ) , .Q( u1_uk_K_r2_55 ) , .QN( u1_uk_n1393 ) );
  DFF_X1 u1_uk_K_r2_reg_6 (.CK( clk ) , .D( u1_uk_K_r1_6 ) , .Q( u1_uk_K_r2_6 ) , .QN( u1_uk_n1354 ) );
  DFF_X1 u1_uk_K_r2_reg_7 (.CK( clk ) , .D( u1_uk_K_r1_7 ) , .Q( u1_uk_K_r2_7 ) );
  DFF_X1 u1_uk_K_r2_reg_8 (.CK( clk ) , .D( u1_uk_K_r1_8 ) , .Q( u1_uk_K_r2_8 ) , .QN( u1_uk_n1355 ) );
  DFF_X1 u1_uk_K_r2_reg_9 (.CK( clk ) , .D( u1_uk_K_r1_9 ) , .Q( u1_uk_K_r2_9 ) , .QN( u1_uk_n1356 ) );
  DFF_X1 u1_uk_K_r3_reg_0 (.CK( clk ) , .D( u1_uk_K_r2_0 ) , .Q( u1_uk_K_r3_0 ) , .QN( u1_uk_n1394 ) );
  DFF_X1 u1_uk_K_r3_reg_1 (.CK( clk ) , .D( u1_uk_K_r2_1 ) , .Q( u1_uk_K_r3_1 ) , .QN( u1_uk_n1395 ) );
  DFF_X1 u1_uk_K_r3_reg_10 (.CK( clk ) , .D( u1_uk_K_r2_10 ) , .Q( u1_uk_K_r3_10 ) );
  DFF_X1 u1_uk_K_r3_reg_11 (.CK( clk ) , .D( u1_uk_K_r2_11 ) , .Q( u1_uk_K_r3_11 ) );
  DFF_X1 u1_uk_K_r3_reg_12 (.CK( clk ) , .D( u1_uk_K_r2_12 ) , .Q( u1_uk_K_r3_12 ) , .QN( u1_uk_n1402 ) );
  DFF_X1 u1_uk_K_r3_reg_13 (.CK( clk ) , .D( u1_uk_K_r2_13 ) , .Q( u1_uk_K_r3_13 ) );
  DFF_X1 u1_uk_K_r3_reg_14 (.CK( clk ) , .D( u1_uk_K_r2_14 ) , .Q( u1_uk_K_r3_14 ) );
  DFF_X1 u1_uk_K_r3_reg_15 (.CK( clk ) , .D( u1_uk_K_r2_15 ) , .Q( u1_uk_K_r3_15 ) );
  DFF_X1 u1_uk_K_r3_reg_16 (.CK( clk ) , .D( u1_uk_K_r2_16 ) , .Q( u1_uk_K_r3_16 ) );
  DFF_X1 u1_uk_K_r3_reg_17 (.CK( clk ) , .D( u1_uk_K_r2_17 ) , .Q( u1_uk_K_r3_17 ) , .QN( u1_uk_n1403 ) );
  DFF_X1 u1_uk_K_r3_reg_18 (.CK( clk ) , .D( u1_uk_K_r2_18 ) , .Q( u1_uk_K_r3_18 ) , .QN( u1_uk_n1404 ) );
  DFF_X1 u1_uk_K_r3_reg_19 (.CK( clk ) , .D( u1_uk_K_r2_19 ) , .Q( u1_uk_K_r3_19 ) );
  DFF_X1 u1_uk_K_r3_reg_2 (.CK( clk ) , .D( u1_uk_K_r2_2 ) , .Q( u1_uk_K_r3_2 ) , .QN( u1_uk_n1396 ) );
  DFF_X1 u1_uk_K_r3_reg_20 (.CK( clk ) , .D( u1_uk_K_r2_20 ) , .Q( u1_uk_K_r3_20 ) , .QN( u1_uk_n1405 ) );
  DFF_X1 u1_uk_K_r3_reg_21 (.CK( clk ) , .D( u1_uk_K_r2_21 ) , .Q( u1_uk_K_r3_21 ) , .QN( u1_uk_n1406 ) );
  DFF_X1 u1_uk_K_r3_reg_22 (.CK( clk ) , .D( u1_uk_K_r2_22 ) , .Q( u1_uk_K_r3_22 ) , .QN( u1_uk_n1407 ) );
  DFF_X1 u1_uk_K_r3_reg_23 (.CK( clk ) , .D( u1_uk_K_r2_23 ) , .Q( u1_uk_K_r3_23 ) , .QN( u1_uk_n1408 ) );
  DFF_X1 u1_uk_K_r3_reg_24 (.CK( clk ) , .D( u1_uk_K_r2_24 ) , .Q( u1_uk_K_r3_24 ) );
  DFF_X1 u1_uk_K_r3_reg_25 (.CK( clk ) , .D( u1_uk_K_r2_25 ) , .Q( u1_uk_K_r3_25 ) , .QN( u1_uk_n1409 ) );
  DFF_X1 u1_uk_K_r3_reg_26 (.CK( clk ) , .D( u1_uk_K_r2_26 ) , .Q( u1_uk_K_r3_26 ) , .QN( u1_uk_n1410 ) );
  DFF_X1 u1_uk_K_r3_reg_27 (.CK( clk ) , .D( u1_uk_K_r2_27 ) , .Q( u1_uk_K_r3_27 ) , .QN( u1_uk_n1411 ) );
  DFF_X1 u1_uk_K_r3_reg_28 (.CK( clk ) , .D( u1_uk_K_r2_28 ) , .Q( u1_uk_K_r3_28 ) , .QN( u1_uk_n1412 ) );
  DFF_X1 u1_uk_K_r3_reg_29 (.CK( clk ) , .D( u1_uk_K_r2_29 ) , .Q( u1_uk_K_r3_29 ) );
  DFF_X1 u1_uk_K_r3_reg_3 (.CK( clk ) , .D( u1_uk_K_r2_3 ) , .Q( u1_uk_K_r3_3 ) , .QN( u1_uk_n1397 ) );
  DFF_X1 u1_uk_K_r3_reg_30 (.CK( clk ) , .D( u1_uk_K_r2_30 ) , .Q( u1_uk_K_r3_30 ) , .QN( u1_uk_n1413 ) );
  DFF_X1 u1_uk_K_r3_reg_31 (.CK( clk ) , .D( u1_uk_K_r2_31 ) , .Q( u1_uk_K_r3_31 ) , .QN( u1_uk_n1414 ) );
  DFF_X1 u1_uk_K_r3_reg_32 (.CK( clk ) , .D( u1_uk_K_r2_32 ) , .Q( u1_uk_K_r3_32 ) , .QN( u1_uk_n1415 ) );
  DFF_X1 u1_uk_K_r3_reg_33 (.CK( clk ) , .D( u1_uk_K_r2_33 ) , .Q( u1_uk_K_r3_33 ) , .QN( u1_uk_n1417 ) );
  DFF_X1 u1_uk_K_r3_reg_34 (.CK( clk ) , .D( u1_uk_K_r2_34 ) , .Q( u1_uk_K_r3_34 ) );
  DFF_X1 u1_uk_K_r3_reg_35 (.CK( clk ) , .D( u1_uk_K_r2_35 ) , .Q( u1_uk_K_r3_35 ) );
  DFF_X1 u1_uk_K_r3_reg_36 (.CK( clk ) , .D( u1_uk_K_r2_36 ) , .Q( u1_uk_K_r3_36 ) , .QN( u1_uk_n1418 ) );
  DFF_X1 u1_uk_K_r3_reg_37 (.CK( clk ) , .D( u1_uk_K_r2_37 ) , .Q( u1_uk_K_r3_37 ) , .QN( u1_uk_n1419 ) );
  DFF_X1 u1_uk_K_r3_reg_38 (.CK( clk ) , .D( u1_uk_K_r2_38 ) , .Q( u1_uk_K_r3_38 ) );
  DFF_X1 u1_uk_K_r3_reg_39 (.CK( clk ) , .D( u1_uk_K_r2_39 ) , .Q( u1_uk_K_r3_39 ) , .QN( u1_uk_n1422 ) );
  DFF_X1 u1_uk_K_r3_reg_4 (.CK( clk ) , .D( u1_uk_K_r2_4 ) , .Q( u1_uk_K_r3_4 ) );
  DFF_X1 u1_uk_K_r3_reg_40 (.CK( clk ) , .D( u1_uk_K_r2_40 ) , .Q( u1_uk_K_r3_40 ) , .QN( u1_uk_n1423 ) );
  DFF_X1 u1_uk_K_r3_reg_41 (.CK( clk ) , .D( u1_uk_K_r2_41 ) , .Q( u1_uk_K_r3_41 ) , .QN( u1_uk_n1424 ) );
  DFF_X1 u1_uk_K_r3_reg_42 (.CK( clk ) , .D( u1_uk_K_r2_42 ) , .Q( u1_uk_K_r3_42 ) , .QN( u1_uk_n1425 ) );
  DFF_X1 u1_uk_K_r3_reg_43 (.CK( clk ) , .D( u1_uk_K_r2_43 ) , .Q( u1_uk_K_r3_43 ) );
  DFF_X1 u1_uk_K_r3_reg_44 (.CK( clk ) , .D( u1_uk_K_r2_44 ) , .Q( u1_uk_K_r3_44 ) );
  DFF_X1 u1_uk_K_r3_reg_45 (.CK( clk ) , .D( u1_uk_K_r2_45 ) , .Q( u1_uk_K_r3_45 ) , .QN( u1_uk_n1426 ) );
  DFF_X1 u1_uk_K_r3_reg_46 (.CK( clk ) , .D( u1_uk_K_r2_46 ) , .Q( u1_uk_K_r3_46 ) , .QN( u1_uk_n1427 ) );
  DFF_X1 u1_uk_K_r3_reg_47 (.CK( clk ) , .D( u1_uk_K_r2_47 ) , .Q( u1_uk_K_r3_47 ) );
  DFF_X1 u1_uk_K_r3_reg_48 (.CK( clk ) , .D( u1_uk_K_r2_48 ) , .Q( u1_uk_K_r3_48 ) , .QN( u1_uk_n1429 ) );
  DFF_X1 u1_uk_K_r3_reg_49 (.CK( clk ) , .D( u1_uk_K_r2_49 ) , .Q( u1_uk_K_r3_49 ) , .QN( u1_uk_n1430 ) );
  DFF_X1 u1_uk_K_r3_reg_5 (.CK( clk ) , .D( u1_uk_K_r2_5 ) , .Q( u1_uk_K_r3_5 ) , .QN( u1_uk_n1398 ) );
  DFF_X1 u1_uk_K_r3_reg_50 (.CK( clk ) , .D( u1_uk_K_r2_50 ) , .Q( u1_uk_K_r3_50 ) , .QN( u1_uk_n1431 ) );
  DFF_X1 u1_uk_K_r3_reg_51 (.CK( clk ) , .D( u1_uk_K_r2_51 ) , .Q( u1_uk_K_r3_51 ) , .QN( u1_uk_n1433 ) );
  DFF_X1 u1_uk_K_r3_reg_52 (.CK( clk ) , .D( u1_uk_K_r2_52 ) , .Q( u1_uk_K_r3_52 ) );
  DFF_X1 u1_uk_K_r3_reg_53 (.CK( clk ) , .D( u1_uk_K_r2_53 ) , .Q( u1_uk_K_r3_53 ) , .QN( u1_uk_n1435 ) );
  DFF_X1 u1_uk_K_r3_reg_54 (.CK( clk ) , .D( u1_uk_K_r2_54 ) , .Q( u1_uk_K_r3_54 ) , .QN( u1_uk_n1436 ) );
  DFF_X1 u1_uk_K_r3_reg_55 (.CK( clk ) , .D( u1_uk_K_r2_55 ) , .Q( u1_uk_K_r3_55 ) , .QN( u1_uk_n1437 ) );
  DFF_X1 u1_uk_K_r3_reg_6 (.CK( clk ) , .D( u1_uk_K_r2_6 ) , .Q( u1_uk_K_r3_6 ) , .QN( u1_uk_n1399 ) );
  DFF_X1 u1_uk_K_r3_reg_7 (.CK( clk ) , .D( u1_uk_K_r2_7 ) , .Q( u1_uk_K_r3_7 ) , .QN( u1_uk_n1400 ) );
  DFF_X1 u1_uk_K_r3_reg_8 (.CK( clk ) , .D( u1_uk_K_r2_8 ) , .Q( u1_uk_K_r3_8 ) , .QN( u1_uk_n1401 ) );
  DFF_X1 u1_uk_K_r3_reg_9 (.CK( clk ) , .D( u1_uk_K_r2_9 ) , .Q( u1_uk_K_r3_9 ) );
  DFF_X1 u1_uk_K_r4_reg_0 (.CK( clk ) , .D( u1_uk_K_r3_0 ) , .Q( u1_uk_K_r4_0 ) );
  DFF_X1 u1_uk_K_r4_reg_1 (.CK( clk ) , .D( u1_uk_K_r3_1 ) , .Q( u1_uk_K_r4_1 ) , .QN( u1_uk_n1438 ) );
  DFF_X1 u1_uk_K_r4_reg_10 (.CK( clk ) , .D( u1_uk_K_r3_10 ) , .Q( u1_uk_K_r4_10 ) , .QN( u1_uk_n1444 ) );
  DFF_X1 u1_uk_K_r4_reg_11 (.CK( clk ) , .D( u1_uk_K_r3_11 ) , .Q( u1_uk_K_r4_11 ) );
  DFF_X1 u1_uk_K_r4_reg_12 (.CK( clk ) , .D( u1_uk_K_r3_12 ) , .Q( u1_uk_K_r4_12 ) , .QN( u1_uk_n1446 ) );
  DFF_X1 u1_uk_K_r4_reg_13 (.CK( clk ) , .D( u1_uk_K_r3_13 ) , .Q( u1_uk_K_r4_13 ) , .QN( u1_uk_n1447 ) );
  DFF_X1 u1_uk_K_r4_reg_14 (.CK( clk ) , .D( u1_uk_K_r3_14 ) , .Q( u1_uk_K_r4_14 ) , .QN( u1_uk_n1448 ) );
  DFF_X1 u1_uk_K_r4_reg_15 (.CK( clk ) , .D( u1_uk_K_r3_15 ) , .Q( u1_uk_K_r4_15 ) , .QN( u1_uk_n1449 ) );
  DFF_X1 u1_uk_K_r4_reg_16 (.CK( clk ) , .D( u1_uk_K_r3_16 ) , .Q( u1_uk_K_r4_16 ) , .QN( u1_uk_n1450 ) );
  DFF_X1 u1_uk_K_r4_reg_17 (.CK( clk ) , .D( u1_uk_K_r3_17 ) , .Q( u1_uk_K_r4_17 ) );
  DFF_X1 u1_uk_K_r4_reg_18 (.CK( clk ) , .D( u1_uk_K_r3_18 ) , .Q( u1_uk_K_r4_18 ) );
  DFF_X1 u1_uk_K_r4_reg_19 (.CK( clk ) , .D( u1_uk_K_r3_19 ) , .Q( u1_uk_K_r4_19 ) , .QN( u1_uk_n1452 ) );
  DFF_X1 u1_uk_K_r4_reg_2 (.CK( clk ) , .D( u1_uk_K_r3_2 ) , .Q( u1_uk_K_r4_2 ) );
  DFF_X1 u1_uk_K_r4_reg_20 (.CK( clk ) , .D( u1_uk_K_r3_20 ) , .Q( u1_uk_K_r4_20 ) , .QN( u1_uk_n1453 ) );
  DFF_X1 u1_uk_K_r4_reg_21 (.CK( clk ) , .D( u1_uk_K_r3_21 ) , .Q( u1_uk_K_r4_21 ) , .QN( u1_uk_n1454 ) );
  DFF_X1 u1_uk_K_r4_reg_22 (.CK( clk ) , .D( u1_uk_K_r3_22 ) , .Q( u1_uk_K_r4_22 ) , .QN( u1_uk_n1455 ) );
  DFF_X1 u1_uk_K_r4_reg_23 (.CK( clk ) , .D( u1_uk_K_r3_23 ) , .Q( u1_uk_K_r4_23 ) );
  DFF_X1 u1_uk_K_r4_reg_24 (.CK( clk ) , .D( u1_uk_K_r3_24 ) , .Q( u1_uk_K_r4_24 ) );
  DFF_X1 u1_uk_K_r4_reg_25 (.CK( clk ) , .D( u1_uk_K_r3_25 ) , .Q( u1_uk_K_r4_25 ) , .QN( u1_uk_n1456 ) );
  DFF_X1 u1_uk_K_r4_reg_26 (.CK( clk ) , .D( u1_uk_K_r3_26 ) , .Q( u1_uk_K_r4_26 ) , .QN( u1_uk_n1457 ) );
  DFF_X1 u1_uk_K_r4_reg_27 (.CK( clk ) , .D( u1_uk_K_r3_27 ) , .Q( u1_uk_K_r4_27 ) );
  DFF_X1 u1_uk_K_r4_reg_28 (.CK( clk ) , .D( u1_uk_K_r3_28 ) , .Q( u1_uk_K_r4_28 ) , .QN( u1_uk_n1458 ) );
  DFF_X1 u1_uk_K_r4_reg_29 (.CK( clk ) , .D( u1_uk_K_r3_29 ) , .Q( u1_uk_K_r4_29 ) , .QN( u1_uk_n1459 ) );
  DFF_X1 u1_uk_K_r4_reg_3 (.CK( clk ) , .D( u1_uk_K_r3_3 ) , .Q( u1_uk_K_r4_3 ) );
  DFF_X1 u1_uk_K_r4_reg_30 (.CK( clk ) , .D( u1_uk_K_r3_30 ) , .Q( u1_uk_K_r4_30 ) , .QN( u1_uk_n1460 ) );
  DFF_X1 u1_uk_K_r4_reg_31 (.CK( clk ) , .D( u1_uk_K_r3_31 ) , .Q( u1_uk_K_r4_31 ) );
  DFF_X1 u1_uk_K_r4_reg_32 (.CK( clk ) , .D( u1_uk_K_r3_32 ) , .Q( u1_uk_K_r4_32 ) , .QN( u1_uk_n1461 ) );
  DFF_X1 u1_uk_K_r4_reg_33 (.CK( clk ) , .D( u1_uk_K_r3_33 ) , .Q( u1_uk_K_r4_33 ) );
  DFF_X1 u1_uk_K_r4_reg_34 (.CK( clk ) , .D( u1_uk_K_r3_34 ) , .Q( u1_uk_K_r4_34 ) , .QN( u1_uk_n1462 ) );
  DFF_X1 u1_uk_K_r4_reg_35 (.CK( clk ) , .D( u1_uk_K_r3_35 ) , .Q( u1_uk_K_r4_35 ) );
  DFF_X1 u1_uk_K_r4_reg_36 (.CK( clk ) , .D( u1_uk_K_r3_36 ) , .Q( u1_uk_K_r4_36 ) , .QN( u1_uk_n1463 ) );
  DFF_X1 u1_uk_K_r4_reg_37 (.CK( clk ) , .D( u1_uk_K_r3_37 ) , .Q( u1_uk_K_r4_37 ) , .QN( u1_uk_n1464 ) );
  DFF_X1 u1_uk_K_r4_reg_38 (.CK( clk ) , .D( u1_uk_K_r3_38 ) , .Q( u1_uk_K_r4_38 ) );
  DFF_X1 u1_uk_K_r4_reg_39 (.CK( clk ) , .D( u1_uk_K_r3_39 ) , .Q( u1_uk_K_r4_39 ) , .QN( u1_uk_n1465 ) );
  DFF_X1 u1_uk_K_r4_reg_4 (.CK( clk ) , .D( u1_uk_K_r3_4 ) , .Q( u1_uk_K_r4_4 ) , .QN( u1_uk_n1439 ) );
  DFF_X1 u1_uk_K_r4_reg_40 (.CK( clk ) , .D( u1_uk_K_r3_40 ) , .Q( u1_uk_K_r4_40 ) , .QN( u1_uk_n1466 ) );
  DFF_X1 u1_uk_K_r4_reg_41 (.CK( clk ) , .D( u1_uk_K_r3_41 ) , .Q( u1_uk_K_r4_41 ) );
  DFF_X1 u1_uk_K_r4_reg_42 (.CK( clk ) , .D( u1_uk_K_r3_42 ) , .Q( u1_uk_K_r4_42 ) , .QN( u1_uk_n1468 ) );
  DFF_X1 u1_uk_K_r4_reg_43 (.CK( clk ) , .D( u1_uk_K_r3_43 ) , .Q( u1_uk_K_r4_43 ) , .QN( u1_uk_n1469 ) );
  DFF_X1 u1_uk_K_r4_reg_44 (.CK( clk ) , .D( u1_uk_K_r3_44 ) , .Q( u1_uk_K_r4_44 ) , .QN( u1_uk_n1470 ) );
  DFF_X1 u1_uk_K_r4_reg_45 (.CK( clk ) , .D( u1_uk_K_r3_45 ) , .Q( u1_uk_K_r4_45 ) , .QN( u1_uk_n1471 ) );
  DFF_X1 u1_uk_K_r4_reg_46 (.CK( clk ) , .D( u1_uk_K_r3_46 ) , .Q( u1_uk_K_r4_46 ) , .QN( u1_uk_n1472 ) );
  DFF_X1 u1_uk_K_r4_reg_47 (.CK( clk ) , .D( u1_uk_K_r3_47 ) , .Q( u1_uk_K_r4_47 ) , .QN( u1_uk_n1474 ) );
  DFF_X1 u1_uk_K_r4_reg_48 (.CK( clk ) , .D( u1_uk_K_r3_48 ) , .Q( u1_uk_K_r4_48 ) );
  DFF_X1 u1_uk_K_r4_reg_49 (.CK( clk ) , .D( u1_uk_K_r3_49 ) , .Q( u1_uk_K_r4_49 ) );
  DFF_X1 u1_uk_K_r4_reg_5 (.CK( clk ) , .D( u1_uk_K_r3_5 ) , .Q( u1_uk_K_r4_5 ) );
  DFF_X1 u1_uk_K_r4_reg_50 (.CK( clk ) , .D( u1_uk_K_r3_50 ) , .Q( u1_uk_K_r4_50 ) , .QN( u1_uk_n1475 ) );
  DFF_X1 u1_uk_K_r4_reg_51 (.CK( clk ) , .D( u1_uk_K_r3_51 ) , .Q( u1_uk_K_r4_51 ) , .QN( u1_uk_n1476 ) );
  DFF_X1 u1_uk_K_r4_reg_52 (.CK( clk ) , .D( u1_uk_K_r3_52 ) , .Q( u1_uk_K_r4_52 ) , .QN( u1_uk_n1477 ) );
  DFF_X1 u1_uk_K_r4_reg_53 (.CK( clk ) , .D( u1_uk_K_r3_53 ) , .Q( u1_uk_K_r4_53 ) , .QN( u1_uk_n1478 ) );
  DFF_X1 u1_uk_K_r4_reg_54 (.CK( clk ) , .D( u1_uk_K_r3_54 ) , .Q( u1_uk_K_r4_54 ) );
  DFF_X1 u1_uk_K_r4_reg_55 (.CK( clk ) , .D( u1_uk_K_r3_55 ) , .Q( u1_uk_K_r4_55 ) );
  DFF_X1 u1_uk_K_r4_reg_6 (.CK( clk ) , .D( u1_uk_K_r3_6 ) , .Q( u1_uk_K_r4_6 ) , .QN( u1_uk_n1440 ) );
  DFF_X1 u1_uk_K_r4_reg_7 (.CK( clk ) , .D( u1_uk_K_r3_7 ) , .Q( u1_uk_K_r4_7 ) , .QN( u1_uk_n1441 ) );
  DFF_X1 u1_uk_K_r4_reg_8 (.CK( clk ) , .D( u1_uk_K_r3_8 ) , .Q( u1_uk_K_r4_8 ) , .QN( u1_uk_n1442 ) );
  DFF_X1 u1_uk_K_r4_reg_9 (.CK( clk ) , .D( u1_uk_K_r3_9 ) , .Q( u1_uk_K_r4_9 ) , .QN( u1_uk_n1443 ) );
  DFF_X1 u1_uk_K_r5_reg_0 (.CK( clk ) , .D( u1_uk_K_r4_0 ) , .Q( u1_uk_K_r5_0 ) );
  DFF_X1 u1_uk_K_r5_reg_1 (.CK( clk ) , .D( u1_uk_K_r4_1 ) , .Q( u1_uk_K_r5_1 ) );
  DFF_X1 u1_uk_K_r5_reg_10 (.CK( clk ) , .D( u1_uk_K_r4_10 ) , .Q( u1_uk_K_r5_10 ) );
  DFF_X1 u1_uk_K_r5_reg_11 (.CK( clk ) , .D( u1_uk_K_r4_11 ) , .Q( u1_uk_K_r5_11 ) , .QN( u1_uk_n1487 ) );
  DFF_X1 u1_uk_K_r5_reg_12 (.CK( clk ) , .D( u1_uk_K_r4_12 ) , .Q( u1_uk_K_r5_12 ) , .QN( u1_uk_n1488 ) );
  DFF_X1 u1_uk_K_r5_reg_13 (.CK( clk ) , .D( u1_uk_K_r4_13 ) , .Q( u1_uk_K_r5_13 ) );
  DFF_X1 u1_uk_K_r5_reg_14 (.CK( clk ) , .D( u1_uk_K_r4_14 ) , .Q( u1_uk_K_r5_14 ) , .QN( u1_uk_n1489 ) );
  DFF_X1 u1_uk_K_r5_reg_15 (.CK( clk ) , .D( u1_uk_K_r4_15 ) , .Q( u1_uk_K_r5_15 ) , .QN( u1_uk_n1490 ) );
  DFF_X1 u1_uk_K_r5_reg_16 (.CK( clk ) , .D( u1_uk_K_r4_16 ) , .Q( u1_uk_K_r5_16 ) );
  DFF_X1 u1_uk_K_r5_reg_17 (.CK( clk ) , .D( u1_uk_K_r4_17 ) , .Q( u1_uk_K_r5_17 ) , .QN( u1_uk_n1491 ) );
  DFF_X1 u1_uk_K_r5_reg_18 (.CK( clk ) , .D( u1_uk_K_r4_18 ) , .Q( u1_uk_K_r5_18 ) );
  DFF_X1 u1_uk_K_r5_reg_19 (.CK( clk ) , .D( u1_uk_K_r4_19 ) , .Q( u1_uk_K_r5_19 ) );
  DFF_X1 u1_uk_K_r5_reg_2 (.CK( clk ) , .D( u1_uk_K_r4_2 ) , .Q( u1_uk_K_r5_2 ) , .QN( u1_uk_n1482 ) );
  DFF_X1 u1_uk_K_r5_reg_20 (.CK( clk ) , .D( u1_uk_K_r4_20 ) , .Q( u1_uk_K_r5_20 ) , .QN( u1_uk_n1492 ) );
  DFF_X1 u1_uk_K_r5_reg_21 (.CK( clk ) , .D( u1_uk_K_r4_21 ) , .Q( u1_uk_K_r5_21 ) );
  DFF_X1 u1_uk_K_r5_reg_22 (.CK( clk ) , .D( u1_uk_K_r4_22 ) , .Q( u1_uk_K_r5_22 ) , .QN( u1_uk_n1494 ) );
  DFF_X1 u1_uk_K_r5_reg_23 (.CK( clk ) , .D( u1_uk_K_r4_23 ) , .Q( u1_uk_K_r5_23 ) );
  DFF_X1 u1_uk_K_r5_reg_24 (.CK( clk ) , .D( u1_uk_K_r4_24 ) , .Q( u1_uk_K_r5_24 ) , .QN( u1_uk_n1495 ) );
  DFF_X1 u1_uk_K_r5_reg_25 (.CK( clk ) , .D( u1_uk_K_r4_25 ) , .Q( u1_uk_K_r5_25 ) , .QN( u1_uk_n1496 ) );
  DFF_X1 u1_uk_K_r5_reg_26 (.CK( clk ) , .D( u1_uk_K_r4_26 ) , .Q( u1_uk_K_r5_26 ) );
  DFF_X1 u1_uk_K_r5_reg_27 (.CK( clk ) , .D( u1_uk_K_r4_27 ) , .Q( u1_uk_K_r5_27 ) , .QN( u1_uk_n1498 ) );
  DFF_X1 u1_uk_K_r5_reg_28 (.CK( clk ) , .D( u1_uk_K_r4_28 ) , .Q( u1_uk_K_r5_28 ) , .QN( u1_uk_n1499 ) );
  DFF_X1 u1_uk_K_r5_reg_29 (.CK( clk ) , .D( u1_uk_K_r4_29 ) , .Q( u1_uk_K_r5_29 ) , .QN( u1_uk_n1500 ) );
  DFF_X1 u1_uk_K_r5_reg_3 (.CK( clk ) , .D( u1_uk_K_r4_3 ) , .Q( u1_uk_K_r5_3 ) , .QN( u1_uk_n1483 ) );
  DFF_X1 u1_uk_K_r5_reg_30 (.CK( clk ) , .D( u1_uk_K_r4_30 ) , .Q( u1_uk_K_r5_30 ) , .QN( u1_uk_n1501 ) );
  DFF_X1 u1_uk_K_r5_reg_31 (.CK( clk ) , .D( u1_uk_K_r4_31 ) , .Q( u1_uk_K_r5_31 ) );
  DFF_X1 u1_uk_K_r5_reg_32 (.CK( clk ) , .D( u1_uk_K_r4_32 ) , .Q( u1_uk_K_r5_32 ) );
  DFF_X1 u1_uk_K_r5_reg_33 (.CK( clk ) , .D( u1_uk_K_r4_33 ) , .Q( u1_uk_K_r5_33 ) , .QN( u1_uk_n1504 ) );
  DFF_X1 u1_uk_K_r5_reg_34 (.CK( clk ) , .D( u1_uk_K_r4_34 ) , .Q( u1_uk_K_r5_34 ) , .QN( u1_uk_n1505 ) );
  DFF_X1 u1_uk_K_r5_reg_35 (.CK( clk ) , .D( u1_uk_K_r4_35 ) , .Q( u1_uk_K_r5_35 ) , .QN( u1_uk_n1507 ) );
  DFF_X1 u1_uk_K_r5_reg_36 (.CK( clk ) , .D( u1_uk_K_r4_36 ) , .Q( u1_uk_K_r5_36 ) , .QN( u1_uk_n1508 ) );
  DFF_X1 u1_uk_K_r5_reg_37 (.CK( clk ) , .D( u1_uk_K_r4_37 ) , .Q( u1_uk_K_r5_37 ) );
  DFF_X1 u1_uk_K_r5_reg_38 (.CK( clk ) , .D( u1_uk_K_r4_38 ) , .Q( u1_uk_K_r5_38 ) , .QN( u1_uk_n1510 ) );
  DFF_X1 u1_uk_K_r5_reg_39 (.CK( clk ) , .D( u1_uk_K_r4_39 ) , .Q( u1_uk_K_r5_39 ) );
  DFF_X1 u1_uk_K_r5_reg_4 (.CK( clk ) , .D( u1_uk_K_r4_4 ) , .Q( u1_uk_K_r5_4 ) );
  DFF_X1 u1_uk_K_r5_reg_40 (.CK( clk ) , .D( u1_uk_K_r4_40 ) , .Q( u1_uk_K_r5_40 ) );
  DFF_X1 u1_uk_K_r5_reg_41 (.CK( clk ) , .D( u1_uk_K_r4_41 ) , .Q( u1_uk_K_r5_41 ) );
  DFF_X1 u1_uk_K_r5_reg_42 (.CK( clk ) , .D( u1_uk_K_r4_42 ) , .Q( u1_uk_K_r5_42 ) , .QN( u1_uk_n1514 ) );
  DFF_X1 u1_uk_K_r5_reg_43 (.CK( clk ) , .D( u1_uk_K_r4_43 ) , .Q( u1_uk_K_r5_43 ) );
  DFF_X1 u1_uk_K_r5_reg_44 (.CK( clk ) , .D( u1_uk_K_r4_44 ) , .Q( u1_uk_K_r5_44 ) , .QN( u1_uk_n1516 ) );
  DFF_X1 u1_uk_K_r5_reg_45 (.CK( clk ) , .D( u1_uk_K_r4_45 ) , .Q( u1_uk_K_r5_45 ) );
  DFF_X1 u1_uk_K_r5_reg_46 (.CK( clk ) , .D( u1_uk_K_r4_46 ) , .Q( u1_uk_K_r5_46 ) , .QN( u1_uk_n1517 ) );
  DFF_X1 u1_uk_K_r5_reg_47 (.CK( clk ) , .D( u1_uk_K_r4_47 ) , .Q( u1_uk_K_r5_47 ) , .QN( u1_uk_n1518 ) );
  DFF_X1 u1_uk_K_r5_reg_48 (.CK( clk ) , .D( u1_uk_K_r4_48 ) , .Q( u1_uk_K_r5_48 ) );
  DFF_X1 u1_uk_K_r5_reg_49 (.CK( clk ) , .D( u1_uk_K_r4_49 ) , .Q( u1_uk_K_r5_49 ) , .QN( u1_uk_n1520 ) );
  DFF_X1 u1_uk_K_r5_reg_5 (.CK( clk ) , .D( u1_uk_K_r4_5 ) , .Q( u1_uk_K_r5_5 ) );
  DFF_X1 u1_uk_K_r5_reg_50 (.CK( clk ) , .D( u1_uk_K_r4_50 ) , .Q( u1_uk_K_r5_50 ) , .QN( u1_uk_n1521 ) );
  DFF_X1 u1_uk_K_r5_reg_51 (.CK( clk ) , .D( u1_uk_K_r4_51 ) , .Q( u1_uk_K_r5_51 ) );
  DFF_X1 u1_uk_K_r5_reg_52 (.CK( clk ) , .D( u1_uk_K_r4_52 ) , .Q( u1_uk_K_r5_52 ) , .QN( u1_uk_n1523 ) );
  DFF_X1 u1_uk_K_r5_reg_53 (.CK( clk ) , .D( u1_uk_K_r4_53 ) , .Q( u1_uk_K_r5_53 ) , .QN( u1_uk_n1524 ) );
  DFF_X1 u1_uk_K_r5_reg_54 (.CK( clk ) , .D( u1_uk_K_r4_54 ) , .Q( u1_uk_K_r5_54 ) , .QN( u1_uk_n1526 ) );
  DFF_X1 u1_uk_K_r5_reg_55 (.CK( clk ) , .D( u1_uk_K_r4_55 ) , .Q( u1_uk_K_r5_55 ) , .QN( u1_uk_n1527 ) );
  DFF_X1 u1_uk_K_r5_reg_6 (.CK( clk ) , .D( u1_uk_K_r4_6 ) , .Q( u1_uk_K_r5_6 ) , .QN( u1_uk_n1484 ) );
  DFF_X1 u1_uk_K_r5_reg_7 (.CK( clk ) , .D( u1_uk_K_r4_7 ) , .Q( u1_uk_K_r5_7 ) , .QN( u1_uk_n1485 ) );
  DFF_X1 u1_uk_K_r5_reg_8 (.CK( clk ) , .D( u1_uk_K_r4_8 ) , .Q( u1_uk_K_r5_8 ) );
  DFF_X1 u1_uk_K_r5_reg_9 (.CK( clk ) , .D( u1_uk_K_r4_9 ) , .Q( u1_uk_K_r5_9 ) , .QN( u1_uk_n1486 ) );
  DFF_X1 u1_uk_K_r6_reg_0 (.CK( clk ) , .D( u1_uk_K_r5_0 ) , .Q( u1_uk_K_r6_0 ) );
  DFF_X1 u1_uk_K_r6_reg_1 (.CK( clk ) , .D( u1_uk_K_r5_1 ) , .Q( u1_uk_K_r6_1 ) , .QN( u1_uk_n1528 ) );
  DFF_X1 u1_uk_K_r6_reg_10 (.CK( clk ) , .D( u1_uk_K_r5_10 ) , .Q( u1_uk_K_r6_10 ) );
  DFF_X1 u1_uk_K_r6_reg_11 (.CK( clk ) , .D( u1_uk_K_r5_11 ) , .Q( u1_uk_K_r6_11 ) , .QN( u1_uk_n1536 ) );
  DFF_X1 u1_uk_K_r6_reg_12 (.CK( clk ) , .D( u1_uk_K_r5_12 ) , .Q( u1_uk_K_r6_12 ) , .QN( u1_uk_n1537 ) );
  DFF_X1 u1_uk_K_r6_reg_13 (.CK( clk ) , .D( u1_uk_K_r5_13 ) , .Q( u1_uk_K_r6_13 ) , .QN( u1_uk_n1538 ) );
  DFF_X1 u1_uk_K_r6_reg_14 (.CK( clk ) , .D( u1_uk_K_r5_14 ) , .Q( u1_uk_K_r6_14 ) );
  DFF_X1 u1_uk_K_r6_reg_15 (.CK( clk ) , .D( u1_uk_K_r5_15 ) , .Q( u1_uk_K_r6_15 ) , .QN( u1_uk_n1540 ) );
  DFF_X1 u1_uk_K_r6_reg_16 (.CK( clk ) , .D( u1_uk_K_r5_16 ) , .Q( u1_uk_K_r6_16 ) , .QN( u1_uk_n1541 ) );
  DFF_X1 u1_uk_K_r6_reg_17 (.CK( clk ) , .D( u1_uk_K_r5_17 ) , .Q( u1_uk_K_r6_17 ) , .QN( u1_uk_n1543 ) );
  DFF_X1 u1_uk_K_r6_reg_18 (.CK( clk ) , .D( u1_uk_K_r5_18 ) , .Q( u1_uk_K_r6_18 ) , .QN( u1_uk_n1544 ) );
  DFF_X1 u1_uk_K_r6_reg_19 (.CK( clk ) , .D( u1_uk_K_r5_19 ) , .Q( u1_uk_K_r6_19 ) );
  DFF_X1 u1_uk_K_r6_reg_2 (.CK( clk ) , .D( u1_uk_K_r5_2 ) , .Q( u1_uk_K_r6_2 ) , .QN( u1_uk_n1529 ) );
  DFF_X1 u1_uk_K_r6_reg_20 (.CK( clk ) , .D( u1_uk_K_r5_20 ) , .Q( u1_uk_K_r6_20 ) , .QN( u1_uk_n1545 ) );
  DFF_X1 u1_uk_K_r6_reg_21 (.CK( clk ) , .D( u1_uk_K_r5_21 ) , .Q( u1_uk_K_r6_21 ) );
  DFF_X1 u1_uk_K_r6_reg_22 (.CK( clk ) , .D( u1_uk_K_r5_22 ) , .Q( u1_uk_K_r6_22 ) );
  DFF_X1 u1_uk_K_r6_reg_23 (.CK( clk ) , .D( u1_uk_K_r5_23 ) , .Q( u1_uk_K_r6_23 ) , .QN( u1_uk_n1547 ) );
  DFF_X1 u1_uk_K_r6_reg_24 (.CK( clk ) , .D( u1_uk_K_r5_24 ) , .Q( u1_uk_K_r6_24 ) , .QN( u1_uk_n1548 ) );
  DFF_X1 u1_uk_K_r6_reg_25 (.CK( clk ) , .D( u1_uk_K_r5_25 ) , .Q( u1_uk_K_r6_25 ) , .QN( u1_uk_n1549 ) );
  DFF_X1 u1_uk_K_r6_reg_26 (.CK( clk ) , .D( u1_uk_K_r5_26 ) , .Q( u1_uk_K_r6_26 ) );
  DFF_X1 u1_uk_K_r6_reg_27 (.CK( clk ) , .D( u1_uk_K_r5_27 ) , .Q( u1_uk_K_r6_27 ) );
  DFF_X1 u1_uk_K_r6_reg_28 (.CK( clk ) , .D( u1_uk_K_r5_28 ) , .Q( u1_uk_K_r6_28 ) );
  DFF_X1 u1_uk_K_r6_reg_29 (.CK( clk ) , .D( u1_uk_K_r5_29 ) , .Q( u1_uk_K_r6_29 ) );
  DFF_X1 u1_uk_K_r6_reg_3 (.CK( clk ) , .D( u1_uk_K_r5_3 ) , .Q( u1_uk_K_r6_3 ) );
  DFF_X1 u1_uk_K_r6_reg_30 (.CK( clk ) , .D( u1_uk_K_r5_30 ) , .Q( u1_uk_K_r6_30 ) );
  DFF_X1 u1_uk_K_r6_reg_31 (.CK( clk ) , .D( u1_uk_K_r5_31 ) , .Q( u1_uk_K_r6_31 ) );
  DFF_X1 u1_uk_K_r6_reg_32 (.CK( clk ) , .D( u1_uk_K_r5_32 ) , .Q( u1_uk_K_r6_32 ) , .QN( u1_uk_n1551 ) );
  DFF_X1 u1_uk_K_r6_reg_33 (.CK( clk ) , .D( u1_uk_K_r5_33 ) , .Q( u1_uk_K_r6_33 ) , .QN( u1_uk_n1552 ) );
  DFF_X1 u1_uk_K_r6_reg_34 (.CK( clk ) , .D( u1_uk_K_r5_34 ) , .Q( u1_uk_K_r6_34 ) );
  DFF_X1 u1_uk_K_r6_reg_35 (.CK( clk ) , .D( u1_uk_K_r5_35 ) , .Q( u1_uk_K_r6_35 ) , .QN( u1_uk_n1554 ) );
  DFF_X1 u1_uk_K_r6_reg_36 (.CK( clk ) , .D( u1_uk_K_r5_36 ) , .Q( u1_uk_K_r6_36 ) , .QN( u1_uk_n1555 ) );
  DFF_X1 u1_uk_K_r6_reg_37 (.CK( clk ) , .D( u1_uk_K_r5_37 ) , .Q( u1_uk_K_r6_37 ) );
  DFF_X1 u1_uk_K_r6_reg_38 (.CK( clk ) , .D( u1_uk_K_r5_38 ) , .Q( u1_uk_K_r6_38 ) , .QN( u1_uk_n1556 ) );
  DFF_X1 u1_uk_K_r6_reg_39 (.CK( clk ) , .D( u1_uk_K_r5_39 ) , .Q( u1_uk_K_r6_39 ) , .QN( u1_uk_n1557 ) );
  DFF_X1 u1_uk_K_r6_reg_4 (.CK( clk ) , .D( u1_uk_K_r5_4 ) , .Q( u1_uk_K_r6_4 ) , .QN( u1_uk_n1530 ) );
  DFF_X1 u1_uk_K_r6_reg_40 (.CK( clk ) , .D( u1_uk_K_r5_40 ) , .Q( u1_uk_K_r6_40 ) , .QN( u1_uk_n1558 ) );
  DFF_X1 u1_uk_K_r6_reg_41 (.CK( clk ) , .D( u1_uk_K_r5_41 ) , .Q( u1_uk_K_r6_41 ) , .QN( u1_uk_n1559 ) );
  DFF_X1 u1_uk_K_r6_reg_42 (.CK( clk ) , .D( u1_uk_K_r5_42 ) , .Q( u1_uk_K_r6_42 ) , .QN( u1_uk_n1560 ) );
  DFF_X1 u1_uk_K_r6_reg_43 (.CK( clk ) , .D( u1_uk_K_r5_43 ) , .Q( u1_uk_K_r6_43 ) , .QN( u1_uk_n1561 ) );
  DFF_X1 u1_uk_K_r6_reg_44 (.CK( clk ) , .D( u1_uk_K_r5_44 ) , .Q( u1_uk_K_r6_44 ) , .QN( u1_uk_n1562 ) );
  DFF_X1 u1_uk_K_r6_reg_45 (.CK( clk ) , .D( u1_uk_K_r5_45 ) , .Q( u1_uk_K_r6_45 ) , .QN( u1_uk_n1563 ) );
  DFF_X1 u1_uk_K_r6_reg_46 (.CK( clk ) , .D( u1_uk_K_r5_46 ) , .Q( u1_uk_K_r6_46 ) );
  DFF_X1 u1_uk_K_r6_reg_47 (.CK( clk ) , .D( u1_uk_K_r5_47 ) , .Q( u1_uk_K_r6_47 ) , .QN( u1_uk_n1564 ) );
  DFF_X1 u1_uk_K_r6_reg_48 (.CK( clk ) , .D( u1_uk_K_r5_48 ) , .Q( u1_uk_K_r6_48 ) , .QN( u1_uk_n1565 ) );
  DFF_X1 u1_uk_K_r6_reg_49 (.CK( clk ) , .D( u1_uk_K_r5_49 ) , .Q( u1_uk_K_r6_49 ) , .QN( u1_uk_n1566 ) );
  DFF_X1 u1_uk_K_r6_reg_5 (.CK( clk ) , .D( u1_uk_K_r5_5 ) , .Q( u1_uk_K_r6_5 ) , .QN( u1_uk_n1531 ) );
  DFF_X1 u1_uk_K_r6_reg_50 (.CK( clk ) , .D( u1_uk_K_r5_50 ) , .Q( u1_uk_K_r6_50 ) , .QN( u1_uk_n1567 ) );
  DFF_X1 u1_uk_K_r6_reg_51 (.CK( clk ) , .D( u1_uk_K_r5_51 ) , .Q( u1_uk_K_r6_51 ) );
  DFF_X1 u1_uk_K_r6_reg_52 (.CK( clk ) , .D( u1_uk_K_r5_52 ) , .Q( u1_uk_K_r6_52 ) , .QN( u1_uk_n1568 ) );
  DFF_X1 u1_uk_K_r6_reg_53 (.CK( clk ) , .D( u1_uk_K_r5_53 ) , .Q( u1_uk_K_r6_53 ) );
  DFF_X1 u1_uk_K_r6_reg_54 (.CK( clk ) , .D( u1_uk_K_r5_54 ) , .Q( u1_uk_K_r6_54 ) , .QN( u1_uk_n1570 ) );
  DFF_X1 u1_uk_K_r6_reg_55 (.CK( clk ) , .D( u1_uk_K_r5_55 ) , .Q( u1_uk_K_r6_55 ) );
  DFF_X1 u1_uk_K_r6_reg_6 (.CK( clk ) , .D( u1_uk_K_r5_6 ) , .Q( u1_uk_K_r6_6 ) , .QN( u1_uk_n1532 ) );
  DFF_X1 u1_uk_K_r6_reg_7 (.CK( clk ) , .D( u1_uk_K_r5_7 ) , .Q( u1_uk_K_r6_7 ) );
  DFF_X1 u1_uk_K_r6_reg_8 (.CK( clk ) , .D( u1_uk_K_r5_8 ) , .Q( u1_uk_K_r6_8 ) , .QN( u1_uk_n1533 ) );
  DFF_X1 u1_uk_K_r6_reg_9 (.CK( clk ) , .D( u1_uk_K_r5_9 ) , .Q( u1_uk_K_r6_9 ) , .QN( u1_uk_n1534 ) );
  DFF_X1 u1_uk_K_r7_reg_0 (.CK( clk ) , .D( u1_uk_K_r6_0 ) , .Q( u1_uk_K_r7_0 ) );
  DFF_X1 u1_uk_K_r7_reg_1 (.CK( clk ) , .D( u1_uk_K_r6_1 ) , .Q( u1_uk_K_r7_1 ) , .QN( u1_uk_n1571 ) );
  DFF_X1 u1_uk_K_r7_reg_10 (.CK( clk ) , .D( u1_uk_K_r6_10 ) , .Q( u1_uk_K_r7_10 ) , .QN( u1_uk_n1577 ) );
  DFF_X1 u1_uk_K_r7_reg_11 (.CK( clk ) , .D( u1_uk_K_r6_11 ) , .Q( u1_uk_K_r7_11 ) , .QN( u1_uk_n1578 ) );
  DFF_X1 u1_uk_K_r7_reg_12 (.CK( clk ) , .D( u1_uk_K_r6_12 ) , .Q( u1_uk_K_r7_12 ) , .QN( u1_uk_n1579 ) );
  DFF_X1 u1_uk_K_r7_reg_13 (.CK( clk ) , .D( u1_uk_K_r6_13 ) , .Q( u1_uk_K_r7_13 ) );
  DFF_X1 u1_uk_K_r7_reg_14 (.CK( clk ) , .D( u1_uk_K_r6_14 ) , .Q( u1_uk_K_r7_14 ) , .QN( u1_uk_n1581 ) );
  DFF_X1 u1_uk_K_r7_reg_15 (.CK( clk ) , .D( u1_uk_K_r6_15 ) , .Q( u1_uk_K_r7_15 ) );
  DFF_X1 u1_uk_K_r7_reg_16 (.CK( clk ) , .D( u1_uk_K_r6_16 ) , .Q( u1_uk_K_r7_16 ) );
  DFF_X1 u1_uk_K_r7_reg_17 (.CK( clk ) , .D( u1_uk_K_r6_17 ) , .Q( u1_uk_K_r7_17 ) , .QN( u1_uk_n1584 ) );
  DFF_X1 u1_uk_K_r7_reg_18 (.CK( clk ) , .D( u1_uk_K_r6_18 ) , .Q( u1_uk_K_r7_18 ) , .QN( u1_uk_n1585 ) );
  DFF_X1 u1_uk_K_r7_reg_19 (.CK( clk ) , .D( u1_uk_K_r6_19 ) , .Q( u1_uk_K_r7_19 ) , .QN( u1_uk_n1586 ) );
  DFF_X1 u1_uk_K_r7_reg_2 (.CK( clk ) , .D( u1_uk_K_r6_2 ) , .Q( u1_uk_K_r7_2 ) , .QN( u1_uk_n1572 ) );
  DFF_X1 u1_uk_K_r7_reg_20 (.CK( clk ) , .D( u1_uk_K_r6_20 ) , .Q( u1_uk_K_r7_20 ) );
  DFF_X1 u1_uk_K_r7_reg_21 (.CK( clk ) , .D( u1_uk_K_r6_21 ) , .Q( u1_uk_K_r7_21 ) , .QN( u1_uk_n1588 ) );
  DFF_X1 u1_uk_K_r7_reg_22 (.CK( clk ) , .D( u1_uk_K_r6_22 ) , .Q( u1_uk_K_r7_22 ) );
  DFF_X1 u1_uk_K_r7_reg_23 (.CK( clk ) , .D( u1_uk_K_r6_23 ) , .Q( u1_uk_K_r7_23 ) );
  DFF_X1 u1_uk_K_r7_reg_24 (.CK( clk ) , .D( u1_uk_K_r6_24 ) , .Q( u1_uk_K_r7_24 ) , .QN( u1_uk_n1592 ) );
  DFF_X1 u1_uk_K_r7_reg_25 (.CK( clk ) , .D( u1_uk_K_r6_25 ) , .Q( u1_uk_K_r7_25 ) , .QN( u1_uk_n1593 ) );
  DFF_X1 u1_uk_K_r7_reg_26 (.CK( clk ) , .D( u1_uk_K_r6_26 ) , .Q( u1_uk_K_r7_26 ) );
  DFF_X1 u1_uk_K_r7_reg_27 (.CK( clk ) , .D( u1_uk_K_r6_27 ) , .Q( u1_uk_K_r7_27 ) );
  DFF_X1 u1_uk_K_r7_reg_28 (.CK( clk ) , .D( u1_uk_K_r6_28 ) , .Q( u1_uk_K_r7_28 ) , .QN( u1_uk_n1595 ) );
  DFF_X1 u1_uk_K_r7_reg_29 (.CK( clk ) , .D( u1_uk_K_r6_29 ) , .Q( u1_uk_K_r7_29 ) );
  DFF_X1 u1_uk_K_r7_reg_3 (.CK( clk ) , .D( u1_uk_K_r6_3 ) , .Q( u1_uk_K_r7_3 ) , .QN( u1_uk_n1573 ) );
  DFF_X1 u1_uk_K_r7_reg_30 (.CK( clk ) , .D( u1_uk_K_r6_30 ) , .Q( u1_uk_K_r7_30 ) );
  DFF_X1 u1_uk_K_r7_reg_31 (.CK( clk ) , .D( u1_uk_K_r6_31 ) , .Q( u1_uk_K_r7_31 ) );
  DFF_X1 u1_uk_K_r7_reg_32 (.CK( clk ) , .D( u1_uk_K_r6_32 ) , .Q( u1_uk_K_r7_32 ) );
  DFF_X1 u1_uk_K_r7_reg_33 (.CK( clk ) , .D( u1_uk_K_r6_33 ) , .Q( u1_uk_K_r7_33 ) , .QN( u1_uk_n1598 ) );
  DFF_X1 u1_uk_K_r7_reg_34 (.CK( clk ) , .D( u1_uk_K_r6_34 ) , .Q( u1_uk_K_r7_34 ) );
  DFF_X1 u1_uk_K_r7_reg_35 (.CK( clk ) , .D( u1_uk_K_r6_35 ) , .Q( u1_uk_K_r7_35 ) , .QN( u1_uk_n1599 ) );
  DFF_X1 u1_uk_K_r7_reg_36 (.CK( clk ) , .D( u1_uk_K_r6_36 ) , .Q( u1_uk_K_r7_36 ) , .QN( u1_uk_n1600 ) );
  DFF_X1 u1_uk_K_r7_reg_37 (.CK( clk ) , .D( u1_uk_K_r6_37 ) , .Q( u1_uk_K_r7_37 ) );
  DFF_X1 u1_uk_K_r7_reg_38 (.CK( clk ) , .D( u1_uk_K_r6_38 ) , .Q( u1_uk_K_r7_38 ) , .QN( u1_uk_n1601 ) );
  DFF_X1 u1_uk_K_r7_reg_39 (.CK( clk ) , .D( u1_uk_K_r6_39 ) , .Q( u1_uk_K_r7_39 ) );
  DFF_X1 u1_uk_K_r7_reg_4 (.CK( clk ) , .D( u1_uk_K_r6_4 ) , .Q( u1_uk_K_r7_4 ) , .QN( u1_uk_n1574 ) );
  DFF_X1 u1_uk_K_r7_reg_40 (.CK( clk ) , .D( u1_uk_K_r6_40 ) , .Q( u1_uk_K_r7_40 ) , .QN( u1_uk_n1603 ) );
  DFF_X1 u1_uk_K_r7_reg_41 (.CK( clk ) , .D( u1_uk_K_r6_41 ) , .Q( u1_uk_K_r7_41 ) , .QN( u1_uk_n1604 ) );
  DFF_X1 u1_uk_K_r7_reg_42 (.CK( clk ) , .D( u1_uk_K_r6_42 ) , .Q( u1_uk_K_r7_42 ) , .QN( u1_uk_n1605 ) );
  DFF_X1 u1_uk_K_r7_reg_43 (.CK( clk ) , .D( u1_uk_K_r6_43 ) , .Q( u1_uk_K_r7_43 ) , .QN( u1_uk_n1606 ) );
  DFF_X1 u1_uk_K_r7_reg_44 (.CK( clk ) , .D( u1_uk_K_r6_44 ) , .Q( u1_uk_K_r7_44 ) , .QN( u1_uk_n1607 ) );
  DFF_X1 u1_uk_K_r7_reg_45 (.CK( clk ) , .D( u1_uk_K_r6_45 ) , .Q( u1_uk_K_r7_45 ) , .QN( u1_uk_n1608 ) );
  DFF_X1 u1_uk_K_r7_reg_46 (.CK( clk ) , .D( u1_uk_K_r6_46 ) , .Q( u1_uk_K_r7_46 ) );
  DFF_X1 u1_uk_K_r7_reg_47 (.CK( clk ) , .D( u1_uk_K_r6_47 ) , .Q( u1_uk_K_r7_47 ) , .QN( u1_uk_n1610 ) );
  DFF_X1 u1_uk_K_r7_reg_48 (.CK( clk ) , .D( u1_uk_K_r6_48 ) , .Q( u1_uk_K_r7_48 ) );
  DFF_X1 u1_uk_K_r7_reg_49 (.CK( clk ) , .D( u1_uk_K_r6_49 ) , .Q( u1_uk_K_r7_49 ) , .QN( u1_uk_n1612 ) );
  DFF_X1 u1_uk_K_r7_reg_5 (.CK( clk ) , .D( u1_uk_K_r6_5 ) , .Q( u1_uk_K_r7_5 ) );
  DFF_X1 u1_uk_K_r7_reg_50 (.CK( clk ) , .D( u1_uk_K_r6_50 ) , .Q( u1_uk_K_r7_50 ) , .QN( u1_uk_n1613 ) );
  DFF_X1 u1_uk_K_r7_reg_51 (.CK( clk ) , .D( u1_uk_K_r6_51 ) , .Q( u1_uk_K_r7_51 ) , .QN( u1_uk_n1614 ) );
  DFF_X1 u1_uk_K_r7_reg_52 (.CK( clk ) , .D( u1_uk_K_r6_52 ) , .Q( u1_uk_K_r7_52 ) , .QN( u1_uk_n1615 ) );
  DFF_X1 u1_uk_K_r7_reg_53 (.CK( clk ) , .D( u1_uk_K_r6_53 ) , .Q( u1_uk_K_r7_53 ) );
  DFF_X1 u1_uk_K_r7_reg_54 (.CK( clk ) , .D( u1_uk_K_r6_54 ) , .Q( u1_uk_K_r7_54 ) , .QN( u1_uk_n1616 ) );
  DFF_X1 u1_uk_K_r7_reg_55 (.CK( clk ) , .D( u1_uk_K_r6_55 ) , .Q( u1_uk_K_r7_55 ) );
  DFF_X1 u1_uk_K_r7_reg_6 (.CK( clk ) , .D( u1_uk_K_r6_6 ) , .Q( u1_uk_K_r7_6 ) );
  DFF_X1 u1_uk_K_r7_reg_7 (.CK( clk ) , .D( u1_uk_K_r6_7 ) , .Q( u1_uk_K_r7_7 ) );
  DFF_X1 u1_uk_K_r7_reg_8 (.CK( clk ) , .D( u1_uk_K_r6_8 ) , .Q( u1_uk_K_r7_8 ) );
  DFF_X1 u1_uk_K_r7_reg_9 (.CK( clk ) , .D( u1_uk_K_r6_9 ) , .Q( u1_uk_K_r7_9 ) );
  DFF_X1 u1_uk_K_r8_reg_0 (.CK( clk ) , .D( u1_uk_K_r7_0 ) , .Q( u1_uk_K_r8_0 ) , .QN( u1_uk_n1618 ) );
  DFF_X1 u1_uk_K_r8_reg_1 (.CK( clk ) , .D( u1_uk_K_r7_1 ) , .Q( u1_uk_K_r8_1 ) , .QN( u1_uk_n1619 ) );
  DFF_X1 u1_uk_K_r8_reg_10 (.CK( clk ) , .D( u1_uk_K_r7_10 ) , .Q( u1_uk_K_r8_10 ) );
  DFF_X1 u1_uk_K_r8_reg_11 (.CK( clk ) , .D( u1_uk_K_r7_11 ) , .Q( u1_uk_K_r8_11 ) , .QN( u1_uk_n1625 ) );
  DFF_X1 u1_uk_K_r8_reg_12 (.CK( clk ) , .D( u1_uk_K_r7_12 ) , .Q( u1_uk_K_r8_12 ) , .QN( u1_uk_n1626 ) );
  DFF_X1 u1_uk_K_r8_reg_13 (.CK( clk ) , .D( u1_uk_K_r7_13 ) , .Q( u1_uk_K_r8_13 ) );
  DFF_X1 u1_uk_K_r8_reg_14 (.CK( clk ) , .D( u1_uk_K_r7_14 ) , .Q( u1_uk_K_r8_14 ) , .QN( u1_uk_n1627 ) );
  DFF_X1 u1_uk_K_r8_reg_15 (.CK( clk ) , .D( u1_uk_K_r7_15 ) , .Q( u1_uk_K_r8_15 ) , .QN( u1_uk_n1628 ) );
  DFF_X1 u1_uk_K_r8_reg_16 (.CK( clk ) , .D( u1_uk_K_r7_16 ) , .Q( u1_uk_K_r8_16 ) );
  DFF_X1 u1_uk_K_r8_reg_17 (.CK( clk ) , .D( u1_uk_K_r7_17 ) , .Q( u1_uk_K_r8_17 ) );
  DFF_X1 u1_uk_K_r8_reg_18 (.CK( clk ) , .D( u1_uk_K_r7_18 ) , .Q( u1_uk_K_r8_18 ) , .QN( u1_uk_n1629 ) );
  DFF_X1 u1_uk_K_r8_reg_19 (.CK( clk ) , .D( u1_uk_K_r7_19 ) , .Q( u1_uk_K_r8_19 ) );
  DFF_X1 u1_uk_K_r8_reg_2 (.CK( clk ) , .D( u1_uk_K_r7_2 ) , .Q( u1_uk_K_r8_2 ) );
  DFF_X1 u1_uk_K_r8_reg_20 (.CK( clk ) , .D( u1_uk_K_r7_20 ) , .Q( u1_uk_K_r8_20 ) , .QN( u1_uk_n1630 ) );
  DFF_X1 u1_uk_K_r8_reg_21 (.CK( clk ) , .D( u1_uk_K_r7_21 ) , .Q( u1_uk_K_r8_21 ) );
  DFF_X1 u1_uk_K_r8_reg_22 (.CK( clk ) , .D( u1_uk_K_r7_22 ) , .Q( u1_uk_K_r8_22 ) );
  DFF_X1 u1_uk_K_r8_reg_23 (.CK( clk ) , .D( u1_uk_K_r7_23 ) , .Q( u1_uk_K_r8_23 ) , .QN( u1_uk_n1632 ) );
  DFF_X1 u1_uk_K_r8_reg_24 (.CK( clk ) , .D( u1_uk_K_r7_24 ) , .Q( u1_uk_K_r8_24 ) , .QN( u1_uk_n1633 ) );
  DFF_X1 u1_uk_K_r8_reg_25 (.CK( clk ) , .D( u1_uk_K_r7_25 ) , .Q( u1_uk_K_r8_25 ) , .QN( u1_uk_n1634 ) );
  DFF_X1 u1_uk_K_r8_reg_26 (.CK( clk ) , .D( u1_uk_K_r7_26 ) , .Q( u1_uk_K_r8_26 ) , .QN( u1_uk_n1635 ) );
  DFF_X1 u1_uk_K_r8_reg_27 (.CK( clk ) , .D( u1_uk_K_r7_27 ) , .Q( u1_uk_K_r8_27 ) );
  DFF_X1 u1_uk_K_r8_reg_28 (.CK( clk ) , .D( u1_uk_K_r7_28 ) , .Q( u1_uk_K_r8_28 ) );
  DFF_X1 u1_uk_K_r8_reg_29 (.CK( clk ) , .D( u1_uk_K_r7_29 ) , .Q( u1_uk_K_r8_29 ) , .QN( u1_uk_n1639 ) );
  DFF_X1 u1_uk_K_r8_reg_3 (.CK( clk ) , .D( u1_uk_K_r7_3 ) , .Q( u1_uk_K_r8_3 ) , .QN( u1_uk_n1620 ) );
  DFF_X1 u1_uk_K_r8_reg_30 (.CK( clk ) , .D( u1_uk_K_r7_30 ) , .Q( u1_uk_K_r8_30 ) , .QN( u1_uk_n1640 ) );
  DFF_X1 u1_uk_K_r8_reg_31 (.CK( clk ) , .D( u1_uk_K_r7_31 ) , .Q( u1_uk_K_r8_31 ) , .QN( u1_uk_n1641 ) );
  DFF_X1 u1_uk_K_r8_reg_32 (.CK( clk ) , .D( u1_uk_K_r7_32 ) , .Q( u1_uk_K_r8_32 ) );
  DFF_X1 u1_uk_K_r8_reg_33 (.CK( clk ) , .D( u1_uk_K_r7_33 ) , .Q( u1_uk_K_r8_33 ) , .QN( u1_uk_n1642 ) );
  DFF_X1 u1_uk_K_r8_reg_34 (.CK( clk ) , .D( u1_uk_K_r7_34 ) , .Q( u1_uk_K_r8_34 ) , .QN( u1_uk_n1643 ) );
  DFF_X1 u1_uk_K_r8_reg_35 (.CK( clk ) , .D( u1_uk_K_r7_35 ) , .Q( u1_uk_K_r8_35 ) , .QN( u1_uk_n1644 ) );
  DFF_X1 u1_uk_K_r8_reg_36 (.CK( clk ) , .D( u1_uk_K_r7_36 ) , .Q( u1_uk_K_r8_36 ) , .QN( u1_uk_n1645 ) );
  DFF_X1 u1_uk_K_r8_reg_37 (.CK( clk ) , .D( u1_uk_K_r7_37 ) , .Q( u1_uk_K_r8_37 ) );
  DFF_X1 u1_uk_K_r8_reg_38 (.CK( clk ) , .D( u1_uk_K_r7_38 ) , .Q( u1_uk_K_r8_38 ) , .QN( u1_uk_n1647 ) );
  DFF_X1 u1_uk_K_r8_reg_39 (.CK( clk ) , .D( u1_uk_K_r7_39 ) , .Q( u1_uk_K_r8_39 ) , .QN( u1_uk_n1649 ) );
  DFF_X1 u1_uk_K_r8_reg_4 (.CK( clk ) , .D( u1_uk_K_r7_4 ) , .Q( u1_uk_K_r8_4 ) , .QN( u1_uk_n1621 ) );
  DFF_X1 u1_uk_K_r8_reg_40 (.CK( clk ) , .D( u1_uk_K_r7_40 ) , .Q( u1_uk_K_r8_40 ) );
  DFF_X1 u1_uk_K_r8_reg_41 (.CK( clk ) , .D( u1_uk_K_r7_41 ) , .Q( u1_uk_K_r8_41 ) );
  DFF_X1 u1_uk_K_r8_reg_42 (.CK( clk ) , .D( u1_uk_K_r7_42 ) , .Q( u1_uk_K_r8_42 ) , .QN( u1_uk_n1651 ) );
  DFF_X1 u1_uk_K_r8_reg_43 (.CK( clk ) , .D( u1_uk_K_r7_43 ) , .Q( u1_uk_K_r8_43 ) );
  DFF_X1 u1_uk_K_r8_reg_44 (.CK( clk ) , .D( u1_uk_K_r7_44 ) , .Q( u1_uk_K_r8_44 ) , .QN( u1_uk_n1652 ) );
  DFF_X1 u1_uk_K_r8_reg_45 (.CK( clk ) , .D( u1_uk_K_r7_45 ) , .Q( u1_uk_K_r8_45 ) );
  DFF_X1 u1_uk_K_r8_reg_46 (.CK( clk ) , .D( u1_uk_K_r7_46 ) , .Q( u1_uk_K_r8_46 ) , .QN( u1_uk_n1653 ) );
  DFF_X1 u1_uk_K_r8_reg_47 (.CK( clk ) , .D( u1_uk_K_r7_47 ) , .Q( u1_uk_K_r8_47 ) , .QN( u1_uk_n1654 ) );
  DFF_X1 u1_uk_K_r8_reg_48 (.CK( clk ) , .D( u1_uk_K_r7_48 ) , .Q( u1_uk_K_r8_48 ) );
  DFF_X1 u1_uk_K_r8_reg_49 (.CK( clk ) , .D( u1_uk_K_r7_49 ) , .Q( u1_uk_K_r8_49 ) , .QN( u1_uk_n1655 ) );
  DFF_X1 u1_uk_K_r8_reg_5 (.CK( clk ) , .D( u1_uk_K_r7_5 ) , .Q( u1_uk_K_r8_5 ) );
  DFF_X1 u1_uk_K_r8_reg_50 (.CK( clk ) , .D( u1_uk_K_r7_50 ) , .Q( u1_uk_K_r8_50 ) , .QN( u1_uk_n1656 ) );
  DFF_X1 u1_uk_K_r8_reg_51 (.CK( clk ) , .D( u1_uk_K_r7_51 ) , .Q( u1_uk_K_r8_51 ) );
  DFF_X1 u1_uk_K_r8_reg_52 (.CK( clk ) , .D( u1_uk_K_r7_52 ) , .Q( u1_uk_K_r8_52 ) );
  DFF_X1 u1_uk_K_r8_reg_53 (.CK( clk ) , .D( u1_uk_K_r7_53 ) , .Q( u1_uk_K_r8_53 ) , .QN( u1_uk_n1659 ) );
  DFF_X1 u1_uk_K_r8_reg_54 (.CK( clk ) , .D( u1_uk_K_r7_54 ) , .Q( u1_uk_K_r8_54 ) , .QN( u1_uk_n1660 ) );
  DFF_X1 u1_uk_K_r8_reg_55 (.CK( clk ) , .D( u1_uk_K_r7_55 ) , .Q( u1_uk_K_r8_55 ) , .QN( u1_uk_n1661 ) );
  DFF_X1 u1_uk_K_r8_reg_6 (.CK( clk ) , .D( u1_uk_K_r7_6 ) , .Q( u1_uk_K_r8_6 ) , .QN( u1_uk_n1622 ) );
  DFF_X1 u1_uk_K_r8_reg_7 (.CK( clk ) , .D( u1_uk_K_r7_7 ) , .Q( u1_uk_K_r8_7 ) , .QN( u1_uk_n1623 ) );
  DFF_X1 u1_uk_K_r8_reg_8 (.CK( clk ) , .D( u1_uk_K_r7_8 ) , .Q( u1_uk_K_r8_8 ) );
  DFF_X1 u1_uk_K_r8_reg_9 (.CK( clk ) , .D( u1_uk_K_r7_9 ) , .Q( u1_uk_K_r8_9 ) , .QN( u1_uk_n1624 ) );
  DFF_X1 u1_uk_K_r9_reg_0 (.CK( clk ) , .D( u1_uk_K_r8_0 ) , .Q( u1_uk_K_r9_0 ) );
  DFF_X1 u1_uk_K_r9_reg_1 (.CK( clk ) , .D( u1_uk_K_r8_1 ) , .Q( u1_uk_K_r9_1 ) , .QN( u1_uk_n1662 ) );
  DFF_X1 u1_uk_K_r9_reg_10 (.CK( clk ) , .D( u1_uk_K_r8_10 ) , .Q( u1_uk_K_r9_10 ) );
  DFF_X1 u1_uk_K_r9_reg_11 (.CK( clk ) , .D( u1_uk_K_r8_11 ) , .Q( u1_uk_K_r9_11 ) , .QN( u1_uk_n1667 ) );
  DFF_X1 u1_uk_K_r9_reg_12 (.CK( clk ) , .D( u1_uk_K_r8_12 ) , .Q( u1_uk_K_r9_12 ) );
  DFF_X1 u1_uk_K_r9_reg_13 (.CK( clk ) , .D( u1_uk_K_r8_13 ) , .Q( u1_uk_K_r9_13 ) , .QN( u1_uk_n1669 ) );
  DFF_X1 u1_uk_K_r9_reg_14 (.CK( clk ) , .D( u1_uk_K_r8_14 ) , .Q( u1_uk_K_r9_14 ) , .QN( u1_uk_n1670 ) );
  DFF_X1 u1_uk_K_r9_reg_15 (.CK( clk ) , .D( u1_uk_K_r8_15 ) , .Q( u1_uk_K_r9_15 ) );
  DFF_X1 u1_uk_K_r9_reg_16 (.CK( clk ) , .D( u1_uk_K_r8_16 ) , .Q( u1_uk_K_r9_16 ) , .QN( u1_uk_n1672 ) );
  DFF_X1 u1_uk_K_r9_reg_17 (.CK( clk ) , .D( u1_uk_K_r8_17 ) , .Q( u1_uk_K_r9_17 ) , .QN( u1_uk_n1673 ) );
  DFF_X1 u1_uk_K_r9_reg_18 (.CK( clk ) , .D( u1_uk_K_r8_18 ) , .Q( u1_uk_K_r9_18 ) );
  DFF_X1 u1_uk_K_r9_reg_19 (.CK( clk ) , .D( u1_uk_K_r8_19 ) , .Q( u1_uk_K_r9_19 ) );
  DFF_X1 u1_uk_K_r9_reg_2 (.CK( clk ) , .D( u1_uk_K_r8_2 ) , .Q( u1_uk_K_r9_2 ) );
  DFF_X1 u1_uk_K_r9_reg_20 (.CK( clk ) , .D( u1_uk_K_r8_20 ) , .Q( u1_uk_K_r9_20 ) , .QN( u1_uk_n1676 ) );
  DFF_X1 u1_uk_K_r9_reg_21 (.CK( clk ) , .D( u1_uk_K_r8_21 ) , .Q( u1_uk_K_r9_21 ) , .QN( u1_uk_n1677 ) );
  DFF_X1 u1_uk_K_r9_reg_22 (.CK( clk ) , .D( u1_uk_K_r8_22 ) , .Q( u1_uk_K_r9_22 ) , .QN( u1_uk_n1678 ) );
  DFF_X1 u1_uk_K_r9_reg_23 (.CK( clk ) , .D( u1_uk_K_r8_23 ) , .Q( u1_uk_K_r9_23 ) );
  DFF_X1 u1_uk_K_r9_reg_24 (.CK( clk ) , .D( u1_uk_K_r8_24 ) , .Q( u1_uk_K_r9_24 ) );
  DFF_X1 u1_uk_K_r9_reg_25 (.CK( clk ) , .D( u1_uk_K_r8_25 ) , .Q( u1_uk_K_r9_25 ) );
  DFF_X1 u1_uk_K_r9_reg_26 (.CK( clk ) , .D( u1_uk_K_r8_26 ) , .Q( u1_uk_K_r9_26 ) , .QN( u1_uk_n1682 ) );
  DFF_X1 u1_uk_K_r9_reg_27 (.CK( clk ) , .D( u1_uk_K_r8_27 ) , .Q( u1_uk_K_r9_27 ) );
  DFF_X1 u1_uk_K_r9_reg_28 (.CK( clk ) , .D( u1_uk_K_r8_28 ) , .Q( u1_uk_K_r9_28 ) , .QN( u1_uk_n1683 ) );
  DFF_X1 u1_uk_K_r9_reg_29 (.CK( clk ) , .D( u1_uk_K_r8_29 ) , .Q( u1_uk_K_r9_29 ) , .QN( u1_uk_n1684 ) );
  DFF_X1 u1_uk_K_r9_reg_3 (.CK( clk ) , .D( u1_uk_K_r8_3 ) , .Q( u1_uk_K_r9_3 ) , .QN( u1_uk_n1663 ) );
  DFF_X1 u1_uk_K_r9_reg_30 (.CK( clk ) , .D( u1_uk_K_r8_30 ) , .Q( u1_uk_K_r9_30 ) );
  DFF_X1 u1_uk_K_r9_reg_31 (.CK( clk ) , .D( u1_uk_K_r8_31 ) , .Q( u1_uk_K_r9_31 ) );
  DFF_X1 u1_uk_K_r9_reg_32 (.CK( clk ) , .D( u1_uk_K_r8_32 ) , .Q( u1_uk_K_r9_32 ) , .QN( u1_uk_n1687 ) );
  DFF_X1 u1_uk_K_r9_reg_33 (.CK( clk ) , .D( u1_uk_K_r8_33 ) , .Q( u1_uk_K_r9_33 ) );
  DFF_X1 u1_uk_K_r9_reg_34 (.CK( clk ) , .D( u1_uk_K_r8_34 ) , .Q( u1_uk_K_r9_34 ) , .QN( u1_uk_n1688 ) );
  DFF_X1 u1_uk_K_r9_reg_35 (.CK( clk ) , .D( u1_uk_K_r8_35 ) , .Q( u1_uk_K_r9_35 ) );
  DFF_X1 u1_uk_K_r9_reg_36 (.CK( clk ) , .D( u1_uk_K_r8_36 ) , .Q( u1_uk_K_r9_36 ) , .QN( u1_uk_n1689 ) );
  DFF_X1 u1_uk_K_r9_reg_37 (.CK( clk ) , .D( u1_uk_K_r8_37 ) , .Q( u1_uk_K_r9_37 ) , .QN( u1_uk_n1690 ) );
  DFF_X1 u1_uk_K_r9_reg_38 (.CK( clk ) , .D( u1_uk_K_r8_38 ) , .Q( u1_uk_K_r9_38 ) );
  DFF_X1 u1_uk_K_r9_reg_39 (.CK( clk ) , .D( u1_uk_K_r8_39 ) , .Q( u1_uk_K_r9_39 ) , .QN( u1_uk_n1691 ) );
  DFF_X1 u1_uk_K_r9_reg_4 (.CK( clk ) , .D( u1_uk_K_r8_4 ) , .Q( u1_uk_K_r9_4 ) );
  DFF_X1 u1_uk_K_r9_reg_40 (.CK( clk ) , .D( u1_uk_K_r8_40 ) , .Q( u1_uk_K_r9_40 ) , .QN( u1_uk_n1692 ) );
  DFF_X1 u1_uk_K_r9_reg_41 (.CK( clk ) , .D( u1_uk_K_r8_41 ) , .Q( u1_uk_K_r9_41 ) , .QN( u1_uk_n1693 ) );
  DFF_X1 u1_uk_K_r9_reg_42 (.CK( clk ) , .D( u1_uk_K_r8_42 ) , .Q( u1_uk_K_r9_42 ) , .QN( u1_uk_n1694 ) );
  DFF_X1 u1_uk_K_r9_reg_43 (.CK( clk ) , .D( u1_uk_K_r8_43 ) , .Q( u1_uk_K_r9_43 ) , .QN( u1_uk_n1695 ) );
  DFF_X1 u1_uk_K_r9_reg_44 (.CK( clk ) , .D( u1_uk_K_r8_44 ) , .Q( u1_uk_K_r9_44 ) , .QN( u1_uk_n1696 ) );
  DFF_X1 u1_uk_K_r9_reg_45 (.CK( clk ) , .D( u1_uk_K_r8_45 ) , .Q( u1_uk_K_r9_45 ) );
  DFF_X1 u1_uk_K_r9_reg_46 (.CK( clk ) , .D( u1_uk_K_r8_46 ) , .Q( u1_uk_K_r9_46 ) , .QN( u1_uk_n1698 ) );
  DFF_X1 u1_uk_K_r9_reg_47 (.CK( clk ) , .D( u1_uk_K_r8_47 ) , .Q( u1_uk_K_r9_47 ) , .QN( u1_uk_n1699 ) );
  DFF_X1 u1_uk_K_r9_reg_48 (.CK( clk ) , .D( u1_uk_K_r8_48 ) , .Q( u1_uk_K_r9_48 ) );
  DFF_X1 u1_uk_K_r9_reg_49 (.CK( clk ) , .D( u1_uk_K_r8_49 ) , .Q( u1_uk_K_r9_49 ) );
  DFF_X1 u1_uk_K_r9_reg_5 (.CK( clk ) , .D( u1_uk_K_r8_5 ) , .Q( u1_uk_K_r9_5 ) );
  DFF_X1 u1_uk_K_r9_reg_50 (.CK( clk ) , .D( u1_uk_K_r8_50 ) , .Q( u1_uk_K_r9_50 ) , .QN( u1_uk_n1702 ) );
  DFF_X1 u1_uk_K_r9_reg_51 (.CK( clk ) , .D( u1_uk_K_r8_51 ) , .Q( u1_uk_K_r9_51 ) , .QN( u1_uk_n1703 ) );
  DFF_X1 u1_uk_K_r9_reg_52 (.CK( clk ) , .D( u1_uk_K_r8_52 ) , .Q( u1_uk_K_r9_52 ) , .QN( u1_uk_n1704 ) );
  DFF_X1 u1_uk_K_r9_reg_53 (.CK( clk ) , .D( u1_uk_K_r8_53 ) , .Q( u1_uk_K_r9_53 ) , .QN( u1_uk_n1705 ) );
  DFF_X1 u1_uk_K_r9_reg_54 (.CK( clk ) , .D( u1_uk_K_r8_54 ) , .Q( u1_uk_K_r9_54 ) );
  DFF_X1 u1_uk_K_r9_reg_55 (.CK( clk ) , .D( u1_uk_K_r8_55 ) , .Q( u1_uk_K_r9_55 ) , .QN( u1_uk_n1707 ) );
  DFF_X1 u1_uk_K_r9_reg_6 (.CK( clk ) , .D( u1_uk_K_r8_6 ) , .Q( u1_uk_K_r9_6 ) );
  DFF_X1 u1_uk_K_r9_reg_7 (.CK( clk ) , .D( u1_uk_K_r8_7 ) , .Q( u1_uk_K_r9_7 ) );
  DFF_X1 u1_uk_K_r9_reg_8 (.CK( clk ) , .D( u1_uk_K_r8_8 ) , .Q( u1_uk_K_r9_8 ) , .QN( u1_uk_n1664 ) );
  DFF_X1 u1_uk_K_r9_reg_9 (.CK( clk ) , .D( u1_uk_K_r8_9 ) , .Q( u1_uk_K_r9_9 ) );
  DFF_X1 u2_L0_reg_1 (.CK( clk ) , .Q( u2_L0_1 ) , .D( u2_desIn_r_7 ) );
  DFF_X1 u2_L0_reg_10 (.CK( clk ) , .Q( u2_L0_10 ) , .D( u2_desIn_r_13 ) );
  DFF_X1 u2_L0_reg_11 (.CK( clk ) , .Q( u2_L0_11 ) , .D( u2_desIn_r_21 ) );
  DFF_X1 u2_L0_reg_12 (.CK( clk ) , .Q( u2_L0_12 ) , .D( u2_desIn_r_29 ) );
  DFF_X1 u2_L0_reg_13 (.CK( clk ) , .Q( u2_L0_13 ) , .D( u2_desIn_r_37 ) );
  DFF_X1 u2_L0_reg_14 (.CK( clk ) , .Q( u2_L0_14 ) , .D( u2_desIn_r_45 ) );
  DFF_X1 u2_L0_reg_15 (.CK( clk ) , .Q( u2_L0_15 ) , .D( u2_desIn_r_53 ) );
  DFF_X1 u2_L0_reg_16 (.CK( clk ) , .Q( u2_L0_16 ) , .D( u2_desIn_r_61 ) );
  DFF_X1 u2_L0_reg_17 (.CK( clk ) , .Q( u2_L0_17 ) , .D( u2_desIn_r_3 ) );
  DFF_X1 u2_L0_reg_18 (.CK( clk ) , .Q( u2_L0_18 ) , .D( u2_desIn_r_11 ) );
  DFF_X1 u2_L0_reg_19 (.CK( clk ) , .Q( u2_L0_19 ) , .D( u2_desIn_r_19 ) );
  DFF_X1 u2_L0_reg_2 (.CK( clk ) , .Q( u2_L0_2 ) , .D( u2_desIn_r_15 ) );
  DFF_X1 u2_L0_reg_20 (.CK( clk ) , .Q( u2_L0_20 ) , .D( u2_desIn_r_27 ) );
  DFF_X1 u2_L0_reg_21 (.CK( clk ) , .Q( u2_L0_21 ) , .D( u2_desIn_r_35 ) );
  DFF_X1 u2_L0_reg_22 (.CK( clk ) , .Q( u2_L0_22 ) , .D( u2_desIn_r_43 ) );
  DFF_X1 u2_L0_reg_23 (.CK( clk ) , .Q( u2_L0_23 ) , .D( u2_desIn_r_51 ) );
  DFF_X1 u2_L0_reg_24 (.CK( clk ) , .Q( u2_L0_24 ) , .D( u2_desIn_r_59 ) );
  DFF_X1 u2_L0_reg_25 (.CK( clk ) , .Q( u2_L0_25 ) , .D( u2_desIn_r_1 ) );
  DFF_X1 u2_L0_reg_26 (.CK( clk ) , .Q( u2_L0_26 ) , .D( u2_desIn_r_9 ) );
  DFF_X1 u2_L0_reg_27 (.CK( clk ) , .Q( u2_L0_27 ) , .D( u2_desIn_r_17 ) );
  DFF_X1 u2_L0_reg_28 (.CK( clk ) , .Q( u2_L0_28 ) , .D( u2_desIn_r_25 ) );
  DFF_X1 u2_L0_reg_29 (.CK( clk ) , .Q( u2_L0_29 ) , .D( u2_desIn_r_33 ) );
  DFF_X1 u2_L0_reg_3 (.CK( clk ) , .Q( u2_L0_3 ) , .D( u2_desIn_r_23 ) );
  DFF_X1 u2_L0_reg_30 (.CK( clk ) , .Q( u2_L0_30 ) , .D( u2_desIn_r_41 ) );
  DFF_X1 u2_L0_reg_31 (.CK( clk ) , .Q( u2_L0_31 ) , .D( u2_desIn_r_49 ) );
  DFF_X1 u2_L0_reg_32 (.CK( clk ) , .Q( u2_L0_32 ) , .D( u2_desIn_r_57 ) );
  DFF_X1 u2_L0_reg_4 (.CK( clk ) , .Q( u2_L0_4 ) , .D( u2_desIn_r_31 ) );
  DFF_X1 u2_L0_reg_5 (.CK( clk ) , .Q( u2_L0_5 ) , .D( u2_desIn_r_39 ) );
  DFF_X1 u2_L0_reg_6 (.CK( clk ) , .Q( u2_L0_6 ) , .D( u2_desIn_r_47 ) );
  DFF_X1 u2_L0_reg_7 (.CK( clk ) , .Q( u2_L0_7 ) , .D( u2_desIn_r_55 ) );
  DFF_X1 u2_L0_reg_8 (.CK( clk ) , .Q( u2_L0_8 ) , .D( u2_desIn_r_63 ) );
  DFF_X1 u2_L0_reg_9 (.CK( clk ) , .Q( u2_L0_9 ) , .D( u2_desIn_r_5 ) );
  DFF_X1 u2_L10_reg_1 (.CK( clk ) , .Q( u2_L10_1 ) , .D( u2_R9_1 ) );
  DFF_X1 u2_L10_reg_10 (.CK( clk ) , .Q( u2_L10_10 ) , .D( u2_R9_10 ) );
  DFF_X1 u2_L10_reg_11 (.CK( clk ) , .Q( u2_L10_11 ) , .D( u2_R9_11 ) );
  DFF_X1 u2_L10_reg_12 (.CK( clk ) , .Q( u2_L10_12 ) , .D( u2_R9_12 ) );
  DFF_X1 u2_L10_reg_13 (.CK( clk ) , .Q( u2_L10_13 ) , .D( u2_R9_13 ) );
  DFF_X1 u2_L10_reg_14 (.CK( clk ) , .Q( u2_L10_14 ) , .D( u2_R9_14 ) );
  DFF_X1 u2_L10_reg_15 (.CK( clk ) , .Q( u2_L10_15 ) , .D( u2_R9_15 ) );
  DFF_X1 u2_L10_reg_16 (.CK( clk ) , .Q( u2_L10_16 ) , .D( u2_R9_16 ) );
  DFF_X1 u2_L10_reg_17 (.CK( clk ) , .Q( u2_L10_17 ) , .D( u2_R9_17 ) );
  DFF_X1 u2_L10_reg_18 (.CK( clk ) , .Q( u2_L10_18 ) , .D( u2_R9_18 ) );
  DFF_X1 u2_L10_reg_19 (.CK( clk ) , .Q( u2_L10_19 ) , .D( u2_R9_19 ) );
  DFF_X1 u2_L10_reg_2 (.CK( clk ) , .Q( u2_L10_2 ) , .D( u2_R9_2 ) );
  DFF_X1 u2_L10_reg_20 (.CK( clk ) , .Q( u2_L10_20 ) , .D( u2_R9_20 ) );
  DFF_X1 u2_L10_reg_21 (.CK( clk ) , .Q( u2_L10_21 ) , .D( u2_R9_21 ) );
  DFF_X1 u2_L10_reg_22 (.CK( clk ) , .Q( u2_L10_22 ) , .D( u2_R9_22 ) );
  DFF_X1 u2_L10_reg_23 (.CK( clk ) , .Q( u2_L10_23 ) , .D( u2_R9_23 ) );
  DFF_X1 u2_L10_reg_24 (.CK( clk ) , .Q( u2_L10_24 ) , .D( u2_R9_24 ) );
  DFF_X1 u2_L10_reg_25 (.CK( clk ) , .Q( u2_L10_25 ) , .D( u2_R9_25 ) );
  DFF_X1 u2_L10_reg_26 (.CK( clk ) , .Q( u2_L10_26 ) , .D( u2_R9_26 ) );
  DFF_X1 u2_L10_reg_27 (.CK( clk ) , .Q( u2_L10_27 ) , .D( u2_R9_27 ) );
  DFF_X1 u2_L10_reg_28 (.CK( clk ) , .Q( u2_L10_28 ) , .D( u2_R9_28 ) );
  DFF_X1 u2_L10_reg_29 (.CK( clk ) , .Q( u2_L10_29 ) , .D( u2_R9_29 ) );
  DFF_X1 u2_L10_reg_3 (.CK( clk ) , .Q( u2_L10_3 ) , .D( u2_R9_3 ) );
  DFF_X1 u2_L10_reg_30 (.CK( clk ) , .Q( u2_L10_30 ) , .D( u2_R9_30 ) );
  DFF_X1 u2_L10_reg_31 (.CK( clk ) , .Q( u2_L10_31 ) , .D( u2_R9_31 ) );
  DFF_X1 u2_L10_reg_32 (.CK( clk ) , .Q( u2_L10_32 ) , .D( u2_R9_32 ) );
  DFF_X1 u2_L10_reg_4 (.CK( clk ) , .Q( u2_L10_4 ) , .D( u2_R9_4 ) );
  DFF_X1 u2_L10_reg_5 (.CK( clk ) , .Q( u2_L10_5 ) , .D( u2_R9_5 ) );
  DFF_X1 u2_L10_reg_6 (.CK( clk ) , .Q( u2_L10_6 ) , .D( u2_R9_6 ) );
  DFF_X1 u2_L10_reg_7 (.CK( clk ) , .Q( u2_L10_7 ) , .D( u2_R9_7 ) );
  DFF_X1 u2_L10_reg_8 (.CK( clk ) , .Q( u2_L10_8 ) , .D( u2_R9_8 ) );
  DFF_X1 u2_L10_reg_9 (.CK( clk ) , .Q( u2_L10_9 ) , .D( u2_R9_9 ) );
  DFF_X1 u2_L11_reg_1 (.CK( clk ) , .Q( u2_L11_1 ) , .D( u2_R10_1 ) );
  DFF_X1 u2_L11_reg_10 (.CK( clk ) , .Q( u2_L11_10 ) , .D( u2_R10_10 ) );
  DFF_X1 u2_L11_reg_11 (.CK( clk ) , .Q( u2_L11_11 ) , .D( u2_R10_11 ) );
  DFF_X1 u2_L11_reg_12 (.CK( clk ) , .Q( u2_L11_12 ) , .D( u2_R10_12 ) );
  DFF_X1 u2_L11_reg_13 (.CK( clk ) , .Q( u2_L11_13 ) , .D( u2_R10_13 ) );
  DFF_X1 u2_L11_reg_14 (.CK( clk ) , .Q( u2_L11_14 ) , .D( u2_R10_14 ) );
  DFF_X1 u2_L11_reg_15 (.CK( clk ) , .Q( u2_L11_15 ) , .D( u2_R10_15 ) );
  DFF_X1 u2_L11_reg_16 (.CK( clk ) , .Q( u2_L11_16 ) , .D( u2_R10_16 ) );
  DFF_X1 u2_L11_reg_17 (.CK( clk ) , .Q( u2_L11_17 ) , .D( u2_R10_17 ) );
  DFF_X1 u2_L11_reg_18 (.CK( clk ) , .Q( u2_L11_18 ) , .D( u2_R10_18 ) );
  DFF_X1 u2_L11_reg_19 (.CK( clk ) , .Q( u2_L11_19 ) , .D( u2_R10_19 ) );
  DFF_X1 u2_L11_reg_2 (.CK( clk ) , .Q( u2_L11_2 ) , .D( u2_R10_2 ) );
  DFF_X1 u2_L11_reg_20 (.CK( clk ) , .Q( u2_L11_20 ) , .D( u2_R10_20 ) );
  DFF_X1 u2_L11_reg_21 (.CK( clk ) , .Q( u2_L11_21 ) , .D( u2_R10_21 ) );
  DFF_X1 u2_L11_reg_22 (.CK( clk ) , .Q( u2_L11_22 ) , .D( u2_R10_22 ) );
  DFF_X1 u2_L11_reg_23 (.CK( clk ) , .Q( u2_L11_23 ) , .D( u2_R10_23 ) );
  DFF_X1 u2_L11_reg_24 (.CK( clk ) , .Q( u2_L11_24 ) , .D( u2_R10_24 ) );
  DFF_X1 u2_L11_reg_25 (.CK( clk ) , .Q( u2_L11_25 ) , .D( u2_R10_25 ) );
  DFF_X1 u2_L11_reg_26 (.CK( clk ) , .Q( u2_L11_26 ) , .D( u2_R10_26 ) );
  DFF_X1 u2_L11_reg_27 (.CK( clk ) , .Q( u2_L11_27 ) , .D( u2_R10_27 ) );
  DFF_X1 u2_L11_reg_28 (.CK( clk ) , .Q( u2_L11_28 ) , .D( u2_R10_28 ) );
  DFF_X1 u2_L11_reg_29 (.CK( clk ) , .Q( u2_L11_29 ) , .D( u2_R10_29 ) );
  DFF_X1 u2_L11_reg_3 (.CK( clk ) , .Q( u2_L11_3 ) , .D( u2_R10_3 ) );
  DFF_X1 u2_L11_reg_30 (.CK( clk ) , .Q( u2_L11_30 ) , .D( u2_R10_30 ) );
  DFF_X1 u2_L11_reg_31 (.CK( clk ) , .Q( u2_L11_31 ) , .D( u2_R10_31 ) );
  DFF_X1 u2_L11_reg_32 (.CK( clk ) , .Q( u2_L11_32 ) , .D( u2_R10_32 ) );
  DFF_X1 u2_L11_reg_4 (.CK( clk ) , .Q( u2_L11_4 ) , .D( u2_R10_4 ) );
  DFF_X1 u2_L11_reg_5 (.CK( clk ) , .Q( u2_L11_5 ) , .D( u2_R10_5 ) );
  DFF_X1 u2_L11_reg_6 (.CK( clk ) , .Q( u2_L11_6 ) , .D( u2_R10_6 ) );
  DFF_X1 u2_L11_reg_7 (.CK( clk ) , .Q( u2_L11_7 ) , .D( u2_R10_7 ) );
  DFF_X1 u2_L11_reg_8 (.CK( clk ) , .Q( u2_L11_8 ) , .D( u2_R10_8 ) );
  DFF_X1 u2_L11_reg_9 (.CK( clk ) , .Q( u2_L11_9 ) , .D( u2_R10_9 ) );
  DFF_X1 u2_L12_reg_1 (.CK( clk ) , .Q( u2_L12_1 ) , .D( u2_R11_1 ) );
  DFF_X1 u2_L12_reg_10 (.CK( clk ) , .Q( u2_L12_10 ) , .D( u2_R11_10 ) );
  DFF_X1 u2_L12_reg_11 (.CK( clk ) , .Q( u2_L12_11 ) , .D( u2_R11_11 ) );
  DFF_X1 u2_L12_reg_12 (.CK( clk ) , .Q( u2_L12_12 ) , .D( u2_R11_12 ) );
  DFF_X1 u2_L12_reg_13 (.CK( clk ) , .Q( u2_L12_13 ) , .D( u2_R11_13 ) );
  DFF_X1 u2_L12_reg_14 (.CK( clk ) , .Q( u2_L12_14 ) , .D( u2_R11_14 ) );
  DFF_X1 u2_L12_reg_15 (.CK( clk ) , .Q( u2_L12_15 ) , .D( u2_R11_15 ) );
  DFF_X1 u2_L12_reg_16 (.CK( clk ) , .Q( u2_L12_16 ) , .D( u2_R11_16 ) );
  DFF_X1 u2_L12_reg_17 (.CK( clk ) , .Q( u2_L12_17 ) , .D( u2_R11_17 ) );
  DFF_X1 u2_L12_reg_18 (.CK( clk ) , .Q( u2_L12_18 ) , .D( u2_R11_18 ) );
  DFF_X1 u2_L12_reg_19 (.CK( clk ) , .Q( u2_L12_19 ) , .D( u2_R11_19 ) );
  DFF_X1 u2_L12_reg_2 (.CK( clk ) , .Q( u2_L12_2 ) , .D( u2_R11_2 ) );
  DFF_X1 u2_L12_reg_20 (.CK( clk ) , .Q( u2_L12_20 ) , .D( u2_R11_20 ) );
  DFF_X1 u2_L12_reg_21 (.CK( clk ) , .Q( u2_L12_21 ) , .D( u2_R11_21 ) );
  DFF_X1 u2_L12_reg_22 (.CK( clk ) , .Q( u2_L12_22 ) , .D( u2_R11_22 ) );
  DFF_X1 u2_L12_reg_23 (.CK( clk ) , .Q( u2_L12_23 ) , .D( u2_R11_23 ) );
  DFF_X1 u2_L12_reg_24 (.CK( clk ) , .Q( u2_L12_24 ) , .D( u2_R11_24 ) );
  DFF_X1 u2_L12_reg_25 (.CK( clk ) , .Q( u2_L12_25 ) , .D( u2_R11_25 ) );
  DFF_X1 u2_L12_reg_26 (.CK( clk ) , .Q( u2_L12_26 ) , .D( u2_R11_26 ) );
  DFF_X1 u2_L12_reg_27 (.CK( clk ) , .Q( u2_L12_27 ) , .D( u2_R11_27 ) );
  DFF_X1 u2_L12_reg_28 (.CK( clk ) , .Q( u2_L12_28 ) , .D( u2_R11_28 ) );
  DFF_X1 u2_L12_reg_29 (.CK( clk ) , .Q( u2_L12_29 ) , .D( u2_R11_29 ) );
  DFF_X1 u2_L12_reg_3 (.CK( clk ) , .Q( u2_L12_3 ) , .D( u2_R11_3 ) );
  DFF_X1 u2_L12_reg_30 (.CK( clk ) , .Q( u2_L12_30 ) , .D( u2_R11_30 ) );
  DFF_X1 u2_L12_reg_31 (.CK( clk ) , .Q( u2_L12_31 ) , .D( u2_R11_31 ) );
  DFF_X1 u2_L12_reg_32 (.CK( clk ) , .Q( u2_L12_32 ) , .D( u2_R11_32 ) );
  DFF_X1 u2_L12_reg_4 (.CK( clk ) , .Q( u2_L12_4 ) , .D( u2_R11_4 ) );
  DFF_X1 u2_L12_reg_5 (.CK( clk ) , .Q( u2_L12_5 ) , .D( u2_R11_5 ) );
  DFF_X1 u2_L12_reg_6 (.CK( clk ) , .Q( u2_L12_6 ) , .D( u2_R11_6 ) );
  DFF_X1 u2_L12_reg_7 (.CK( clk ) , .Q( u2_L12_7 ) , .D( u2_R11_7 ) );
  DFF_X1 u2_L12_reg_8 (.CK( clk ) , .Q( u2_L12_8 ) , .D( u2_R11_8 ) );
  DFF_X1 u2_L12_reg_9 (.CK( clk ) , .Q( u2_L12_9 ) , .D( u2_R11_9 ) );
  DFF_X1 u2_L13_reg_1 (.CK( clk ) , .Q( u2_L13_1 ) , .D( u2_R12_1 ) );
  DFF_X1 u2_L13_reg_10 (.CK( clk ) , .Q( u2_L13_10 ) , .D( u2_R12_10 ) );
  DFF_X1 u2_L13_reg_11 (.CK( clk ) , .Q( u2_L13_11 ) , .D( u2_R12_11 ) );
  DFF_X1 u2_L13_reg_12 (.CK( clk ) , .Q( u2_L13_12 ) , .D( u2_R12_12 ) );
  DFF_X1 u2_L13_reg_13 (.CK( clk ) , .Q( u2_L13_13 ) , .D( u2_R12_13 ) );
  DFF_X1 u2_L13_reg_14 (.CK( clk ) , .Q( u2_L13_14 ) , .D( u2_R12_14 ) );
  DFF_X1 u2_L13_reg_15 (.CK( clk ) , .Q( u2_L13_15 ) , .D( u2_R12_15 ) );
  DFF_X1 u2_L13_reg_16 (.CK( clk ) , .Q( u2_L13_16 ) , .D( u2_R12_16 ) );
  DFF_X1 u2_L13_reg_17 (.CK( clk ) , .Q( u2_L13_17 ) , .D( u2_R12_17 ) );
  DFF_X1 u2_L13_reg_18 (.CK( clk ) , .Q( u2_L13_18 ) , .D( u2_R12_18 ) );
  DFF_X1 u2_L13_reg_19 (.CK( clk ) , .Q( u2_L13_19 ) , .D( u2_R12_19 ) );
  DFF_X1 u2_L13_reg_2 (.CK( clk ) , .Q( u2_L13_2 ) , .D( u2_R12_2 ) );
  DFF_X1 u2_L13_reg_20 (.CK( clk ) , .Q( u2_L13_20 ) , .D( u2_R12_20 ) );
  DFF_X1 u2_L13_reg_21 (.CK( clk ) , .Q( u2_L13_21 ) , .D( u2_R12_21 ) );
  DFF_X1 u2_L13_reg_22 (.CK( clk ) , .Q( u2_L13_22 ) , .D( u2_R12_22 ) );
  DFF_X1 u2_L13_reg_23 (.CK( clk ) , .Q( u2_L13_23 ) , .D( u2_R12_23 ) );
  DFF_X1 u2_L13_reg_24 (.CK( clk ) , .Q( u2_L13_24 ) , .D( u2_R12_24 ) );
  DFF_X1 u2_L13_reg_25 (.CK( clk ) , .Q( u2_L13_25 ) , .D( u2_R12_25 ) );
  DFF_X1 u2_L13_reg_26 (.CK( clk ) , .Q( u2_L13_26 ) , .D( u2_R12_26 ) );
  DFF_X1 u2_L13_reg_27 (.CK( clk ) , .Q( u2_L13_27 ) , .D( u2_R12_27 ) );
  DFF_X1 u2_L13_reg_28 (.CK( clk ) , .Q( u2_L13_28 ) , .D( u2_R12_28 ) );
  DFF_X1 u2_L13_reg_29 (.CK( clk ) , .Q( u2_L13_29 ) , .D( u2_R12_29 ) );
  DFF_X1 u2_L13_reg_3 (.CK( clk ) , .Q( u2_L13_3 ) , .D( u2_R12_3 ) );
  DFF_X1 u2_L13_reg_30 (.CK( clk ) , .Q( u2_L13_30 ) , .D( u2_R12_30 ) );
  DFF_X1 u2_L13_reg_31 (.CK( clk ) , .Q( u2_L13_31 ) , .D( u2_R12_31 ) );
  DFF_X1 u2_L13_reg_32 (.CK( clk ) , .Q( u2_L13_32 ) , .D( u2_R12_32 ) );
  DFF_X1 u2_L13_reg_4 (.CK( clk ) , .Q( u2_L13_4 ) , .D( u2_R12_4 ) );
  DFF_X1 u2_L13_reg_5 (.CK( clk ) , .Q( u2_L13_5 ) , .D( u2_R12_5 ) );
  DFF_X1 u2_L13_reg_6 (.CK( clk ) , .Q( u2_L13_6 ) , .D( u2_R12_6 ) );
  DFF_X1 u2_L13_reg_7 (.CK( clk ) , .Q( u2_L13_7 ) , .D( u2_R12_7 ) );
  DFF_X1 u2_L13_reg_8 (.CK( clk ) , .Q( u2_L13_8 ) , .D( u2_R12_8 ) );
  DFF_X1 u2_L13_reg_9 (.CK( clk ) , .Q( u2_L13_9 ) , .D( u2_R12_9 ) );
  DFF_X1 u2_L14_reg_1 (.CK( clk ) , .Q( u2_L14_1 ) , .D( u2_R13_1 ) );
  DFF_X1 u2_L14_reg_10 (.CK( clk ) , .Q( u2_L14_10 ) , .D( u2_R13_10 ) );
  DFF_X1 u2_L14_reg_11 (.CK( clk ) , .Q( u2_L14_11 ) , .D( u2_R13_11 ) );
  DFF_X1 u2_L14_reg_12 (.CK( clk ) , .Q( u2_L14_12 ) , .D( u2_R13_12 ) );
  DFF_X1 u2_L14_reg_13 (.CK( clk ) , .Q( u2_L14_13 ) , .D( u2_R13_13 ) );
  DFF_X1 u2_L14_reg_14 (.CK( clk ) , .Q( u2_L14_14 ) , .D( u2_R13_14 ) );
  DFF_X1 u2_L14_reg_15 (.CK( clk ) , .Q( u2_L14_15 ) , .D( u2_R13_15 ) );
  DFF_X1 u2_L14_reg_16 (.CK( clk ) , .Q( u2_L14_16 ) , .D( u2_R13_16 ) );
  DFF_X1 u2_L14_reg_17 (.CK( clk ) , .Q( u2_L14_17 ) , .D( u2_R13_17 ) );
  DFF_X1 u2_L14_reg_18 (.CK( clk ) , .Q( u2_L14_18 ) , .D( u2_R13_18 ) );
  DFF_X1 u2_L14_reg_19 (.CK( clk ) , .Q( u2_L14_19 ) , .D( u2_R13_19 ) );
  DFF_X1 u2_L14_reg_2 (.CK( clk ) , .Q( u2_L14_2 ) , .D( u2_R13_2 ) );
  DFF_X1 u2_L14_reg_20 (.CK( clk ) , .Q( u2_L14_20 ) , .D( u2_R13_20 ) );
  DFF_X1 u2_L14_reg_21 (.CK( clk ) , .Q( u2_L14_21 ) , .D( u2_R13_21 ) );
  DFF_X1 u2_L14_reg_22 (.CK( clk ) , .Q( u2_L14_22 ) , .D( u2_R13_22 ) );
  DFF_X1 u2_L14_reg_23 (.CK( clk ) , .Q( u2_L14_23 ) , .D( u2_R13_23 ) );
  DFF_X1 u2_L14_reg_24 (.CK( clk ) , .Q( u2_L14_24 ) , .D( u2_R13_24 ) );
  DFF_X1 u2_L14_reg_25 (.CK( clk ) , .Q( u2_L14_25 ) , .D( u2_R13_25 ) );
  DFF_X1 u2_L14_reg_26 (.CK( clk ) , .Q( u2_L14_26 ) , .D( u2_R13_26 ) );
  DFF_X1 u2_L14_reg_27 (.CK( clk ) , .Q( u2_L14_27 ) , .D( u2_R13_27 ) );
  DFF_X1 u2_L14_reg_28 (.CK( clk ) , .Q( u2_L14_28 ) , .D( u2_R13_28 ) );
  DFF_X1 u2_L14_reg_29 (.CK( clk ) , .Q( u2_L14_29 ) , .D( u2_R13_29 ) );
  DFF_X1 u2_L14_reg_3 (.CK( clk ) , .Q( u2_L14_3 ) , .D( u2_R13_3 ) );
  DFF_X1 u2_L14_reg_30 (.CK( clk ) , .Q( u2_L14_30 ) , .D( u2_R13_30 ) );
  DFF_X1 u2_L14_reg_31 (.CK( clk ) , .Q( u2_L14_31 ) , .D( u2_R13_31 ) );
  DFF_X1 u2_L14_reg_32 (.CK( clk ) , .Q( u2_L14_32 ) , .D( u2_R13_32 ) );
  DFF_X1 u2_L14_reg_4 (.CK( clk ) , .Q( u2_L14_4 ) , .D( u2_R13_4 ) );
  DFF_X1 u2_L14_reg_5 (.CK( clk ) , .Q( u2_L14_5 ) , .D( u2_R13_5 ) );
  DFF_X1 u2_L14_reg_6 (.CK( clk ) , .Q( u2_L14_6 ) , .D( u2_R13_6 ) );
  DFF_X1 u2_L14_reg_7 (.CK( clk ) , .Q( u2_L14_7 ) , .D( u2_R13_7 ) );
  DFF_X1 u2_L14_reg_8 (.CK( clk ) , .Q( u2_L14_8 ) , .D( u2_R13_8 ) );
  DFF_X1 u2_L14_reg_9 (.CK( clk ) , .Q( u2_L14_9 ) , .D( u2_R13_9 ) );
  DFF_X1 u2_L1_reg_1 (.CK( clk ) , .Q( u2_L1_1 ) , .D( u2_R0_1 ) );
  DFF_X1 u2_L1_reg_10 (.CK( clk ) , .Q( u2_L1_10 ) , .D( u2_R0_10 ) );
  DFF_X1 u2_L1_reg_11 (.CK( clk ) , .Q( u2_L1_11 ) , .D( u2_R0_11 ) );
  DFF_X1 u2_L1_reg_12 (.CK( clk ) , .Q( u2_L1_12 ) , .D( u2_R0_12 ) );
  DFF_X1 u2_L1_reg_13 (.CK( clk ) , .Q( u2_L1_13 ) , .D( u2_R0_13 ) );
  DFF_X1 u2_L1_reg_14 (.CK( clk ) , .Q( u2_L1_14 ) , .D( u2_R0_14 ) );
  DFF_X1 u2_L1_reg_15 (.CK( clk ) , .Q( u2_L1_15 ) , .D( u2_R0_15 ) );
  DFF_X1 u2_L1_reg_16 (.CK( clk ) , .Q( u2_L1_16 ) , .D( u2_R0_16 ) );
  DFF_X1 u2_L1_reg_17 (.CK( clk ) , .Q( u2_L1_17 ) , .D( u2_R0_17 ) );
  DFF_X1 u2_L1_reg_18 (.CK( clk ) , .Q( u2_L1_18 ) , .D( u2_R0_18 ) );
  DFF_X1 u2_L1_reg_19 (.CK( clk ) , .Q( u2_L1_19 ) , .D( u2_R0_19 ) );
  DFF_X1 u2_L1_reg_2 (.CK( clk ) , .Q( u2_L1_2 ) , .D( u2_R0_2 ) );
  DFF_X1 u2_L1_reg_20 (.CK( clk ) , .Q( u2_L1_20 ) , .D( u2_R0_20 ) );
  DFF_X1 u2_L1_reg_21 (.CK( clk ) , .Q( u2_L1_21 ) , .D( u2_R0_21 ) );
  DFF_X1 u2_L1_reg_22 (.CK( clk ) , .Q( u2_L1_22 ) , .D( u2_R0_22 ) );
  DFF_X1 u2_L1_reg_23 (.CK( clk ) , .Q( u2_L1_23 ) , .D( u2_R0_23 ) );
  DFF_X1 u2_L1_reg_24 (.CK( clk ) , .Q( u2_L1_24 ) , .D( u2_R0_24 ) );
  DFF_X1 u2_L1_reg_25 (.CK( clk ) , .Q( u2_L1_25 ) , .D( u2_R0_25 ) );
  DFF_X1 u2_L1_reg_26 (.CK( clk ) , .Q( u2_L1_26 ) , .D( u2_R0_26 ) );
  DFF_X1 u2_L1_reg_27 (.CK( clk ) , .Q( u2_L1_27 ) , .D( u2_R0_27 ) );
  DFF_X1 u2_L1_reg_28 (.CK( clk ) , .Q( u2_L1_28 ) , .D( u2_R0_28 ) );
  DFF_X1 u2_L1_reg_29 (.CK( clk ) , .Q( u2_L1_29 ) , .D( u2_R0_29 ) );
  DFF_X1 u2_L1_reg_3 (.CK( clk ) , .Q( u2_L1_3 ) , .D( u2_R0_3 ) );
  DFF_X1 u2_L1_reg_30 (.CK( clk ) , .Q( u2_L1_30 ) , .D( u2_R0_30 ) );
  DFF_X1 u2_L1_reg_31 (.CK( clk ) , .Q( u2_L1_31 ) , .D( u2_R0_31 ) );
  DFF_X1 u2_L1_reg_32 (.CK( clk ) , .Q( u2_L1_32 ) , .D( u2_R0_32 ) );
  DFF_X1 u2_L1_reg_4 (.CK( clk ) , .Q( u2_L1_4 ) , .D( u2_R0_4 ) );
  DFF_X1 u2_L1_reg_5 (.CK( clk ) , .Q( u2_L1_5 ) , .D( u2_R0_5 ) );
  DFF_X1 u2_L1_reg_6 (.CK( clk ) , .Q( u2_L1_6 ) , .D( u2_R0_6 ) );
  DFF_X1 u2_L1_reg_7 (.CK( clk ) , .Q( u2_L1_7 ) , .D( u2_R0_7 ) );
  DFF_X1 u2_L1_reg_8 (.CK( clk ) , .Q( u2_L1_8 ) , .D( u2_R0_8 ) );
  DFF_X1 u2_L1_reg_9 (.CK( clk ) , .Q( u2_L1_9 ) , .D( u2_R0_9 ) );
  DFF_X1 u2_L2_reg_1 (.CK( clk ) , .Q( u2_L2_1 ) , .D( u2_R1_1 ) );
  DFF_X1 u2_L2_reg_10 (.CK( clk ) , .Q( u2_L2_10 ) , .D( u2_R1_10 ) );
  DFF_X1 u2_L2_reg_11 (.CK( clk ) , .Q( u2_L2_11 ) , .D( u2_R1_11 ) );
  DFF_X1 u2_L2_reg_12 (.CK( clk ) , .Q( u2_L2_12 ) , .D( u2_R1_12 ) );
  DFF_X1 u2_L2_reg_13 (.CK( clk ) , .Q( u2_L2_13 ) , .D( u2_R1_13 ) );
  DFF_X1 u2_L2_reg_14 (.CK( clk ) , .Q( u2_L2_14 ) , .D( u2_R1_14 ) );
  DFF_X1 u2_L2_reg_15 (.CK( clk ) , .Q( u2_L2_15 ) , .D( u2_R1_15 ) );
  DFF_X1 u2_L2_reg_16 (.CK( clk ) , .Q( u2_L2_16 ) , .D( u2_R1_16 ) );
  DFF_X1 u2_L2_reg_17 (.CK( clk ) , .Q( u2_L2_17 ) , .D( u2_R1_17 ) );
  DFF_X1 u2_L2_reg_18 (.CK( clk ) , .Q( u2_L2_18 ) , .D( u2_R1_18 ) );
  DFF_X1 u2_L2_reg_19 (.CK( clk ) , .Q( u2_L2_19 ) , .D( u2_R1_19 ) );
  DFF_X1 u2_L2_reg_2 (.CK( clk ) , .Q( u2_L2_2 ) , .D( u2_R1_2 ) );
  DFF_X1 u2_L2_reg_20 (.CK( clk ) , .Q( u2_L2_20 ) , .D( u2_R1_20 ) );
  DFF_X1 u2_L2_reg_21 (.CK( clk ) , .Q( u2_L2_21 ) , .D( u2_R1_21 ) );
  DFF_X1 u2_L2_reg_22 (.CK( clk ) , .Q( u2_L2_22 ) , .D( u2_R1_22 ) );
  DFF_X1 u2_L2_reg_23 (.CK( clk ) , .Q( u2_L2_23 ) , .D( u2_R1_23 ) );
  DFF_X1 u2_L2_reg_24 (.CK( clk ) , .Q( u2_L2_24 ) , .D( u2_R1_24 ) );
  DFF_X1 u2_L2_reg_25 (.CK( clk ) , .Q( u2_L2_25 ) , .D( u2_R1_25 ) );
  DFF_X1 u2_L2_reg_26 (.CK( clk ) , .Q( u2_L2_26 ) , .D( u2_R1_26 ) );
  DFF_X1 u2_L2_reg_27 (.CK( clk ) , .Q( u2_L2_27 ) , .D( u2_R1_27 ) );
  DFF_X1 u2_L2_reg_28 (.CK( clk ) , .Q( u2_L2_28 ) , .D( u2_R1_28 ) );
  DFF_X1 u2_L2_reg_29 (.CK( clk ) , .Q( u2_L2_29 ) , .D( u2_R1_29 ) );
  DFF_X1 u2_L2_reg_3 (.CK( clk ) , .Q( u2_L2_3 ) , .D( u2_R1_3 ) );
  DFF_X1 u2_L2_reg_30 (.CK( clk ) , .Q( u2_L2_30 ) , .D( u2_R1_30 ) );
  DFF_X1 u2_L2_reg_31 (.CK( clk ) , .Q( u2_L2_31 ) , .D( u2_R1_31 ) );
  DFF_X1 u2_L2_reg_32 (.CK( clk ) , .Q( u2_L2_32 ) , .D( u2_R1_32 ) );
  DFF_X1 u2_L2_reg_4 (.CK( clk ) , .Q( u2_L2_4 ) , .D( u2_R1_4 ) );
  DFF_X1 u2_L2_reg_5 (.CK( clk ) , .Q( u2_L2_5 ) , .D( u2_R1_5 ) );
  DFF_X1 u2_L2_reg_6 (.CK( clk ) , .Q( u2_L2_6 ) , .D( u2_R1_6 ) );
  DFF_X1 u2_L2_reg_7 (.CK( clk ) , .Q( u2_L2_7 ) , .D( u2_R1_7 ) );
  DFF_X1 u2_L2_reg_8 (.CK( clk ) , .Q( u2_L2_8 ) , .D( u2_R1_8 ) );
  DFF_X1 u2_L2_reg_9 (.CK( clk ) , .Q( u2_L2_9 ) , .D( u2_R1_9 ) );
  DFF_X1 u2_L3_reg_1 (.CK( clk ) , .Q( u2_L3_1 ) , .D( u2_R2_1 ) );
  DFF_X1 u2_L3_reg_10 (.CK( clk ) , .Q( u2_L3_10 ) , .D( u2_R2_10 ) );
  DFF_X1 u2_L3_reg_11 (.CK( clk ) , .Q( u2_L3_11 ) , .D( u2_R2_11 ) );
  DFF_X1 u2_L3_reg_12 (.CK( clk ) , .Q( u2_L3_12 ) , .D( u2_R2_12 ) );
  DFF_X1 u2_L3_reg_13 (.CK( clk ) , .Q( u2_L3_13 ) , .D( u2_R2_13 ) );
  DFF_X1 u2_L3_reg_14 (.CK( clk ) , .Q( u2_L3_14 ) , .D( u2_R2_14 ) );
  DFF_X1 u2_L3_reg_15 (.CK( clk ) , .Q( u2_L3_15 ) , .D( u2_R2_15 ) );
  DFF_X1 u2_L3_reg_16 (.CK( clk ) , .Q( u2_L3_16 ) , .D( u2_R2_16 ) );
  DFF_X1 u2_L3_reg_17 (.CK( clk ) , .Q( u2_L3_17 ) , .D( u2_R2_17 ) );
  DFF_X1 u2_L3_reg_18 (.CK( clk ) , .Q( u2_L3_18 ) , .D( u2_R2_18 ) );
  DFF_X1 u2_L3_reg_19 (.CK( clk ) , .Q( u2_L3_19 ) , .D( u2_R2_19 ) );
  DFF_X1 u2_L3_reg_2 (.CK( clk ) , .Q( u2_L3_2 ) , .D( u2_R2_2 ) );
  DFF_X1 u2_L3_reg_20 (.CK( clk ) , .Q( u2_L3_20 ) , .D( u2_R2_20 ) );
  DFF_X1 u2_L3_reg_21 (.CK( clk ) , .Q( u2_L3_21 ) , .D( u2_R2_21 ) );
  DFF_X1 u2_L3_reg_22 (.CK( clk ) , .Q( u2_L3_22 ) , .D( u2_R2_22 ) );
  DFF_X1 u2_L3_reg_23 (.CK( clk ) , .Q( u2_L3_23 ) , .D( u2_R2_23 ) );
  DFF_X1 u2_L3_reg_24 (.CK( clk ) , .Q( u2_L3_24 ) , .D( u2_R2_24 ) );
  DFF_X1 u2_L3_reg_25 (.CK( clk ) , .Q( u2_L3_25 ) , .D( u2_R2_25 ) );
  DFF_X1 u2_L3_reg_26 (.CK( clk ) , .Q( u2_L3_26 ) , .D( u2_R2_26 ) );
  DFF_X1 u2_L3_reg_27 (.CK( clk ) , .Q( u2_L3_27 ) , .D( u2_R2_27 ) );
  DFF_X1 u2_L3_reg_28 (.CK( clk ) , .Q( u2_L3_28 ) , .D( u2_R2_28 ) );
  DFF_X1 u2_L3_reg_29 (.CK( clk ) , .Q( u2_L3_29 ) , .D( u2_R2_29 ) );
  DFF_X1 u2_L3_reg_3 (.CK( clk ) , .Q( u2_L3_3 ) , .D( u2_R2_3 ) );
  DFF_X1 u2_L3_reg_30 (.CK( clk ) , .Q( u2_L3_30 ) , .D( u2_R2_30 ) );
  DFF_X1 u2_L3_reg_31 (.CK( clk ) , .Q( u2_L3_31 ) , .D( u2_R2_31 ) );
  DFF_X1 u2_L3_reg_32 (.CK( clk ) , .Q( u2_L3_32 ) , .D( u2_R2_32 ) );
  DFF_X1 u2_L3_reg_4 (.CK( clk ) , .Q( u2_L3_4 ) , .D( u2_R2_4 ) );
  DFF_X1 u2_L3_reg_5 (.CK( clk ) , .Q( u2_L3_5 ) , .D( u2_R2_5 ) );
  DFF_X1 u2_L3_reg_6 (.CK( clk ) , .Q( u2_L3_6 ) , .D( u2_R2_6 ) );
  DFF_X1 u2_L3_reg_7 (.CK( clk ) , .Q( u2_L3_7 ) , .D( u2_R2_7 ) );
  DFF_X1 u2_L3_reg_8 (.CK( clk ) , .Q( u2_L3_8 ) , .D( u2_R2_8 ) );
  DFF_X1 u2_L3_reg_9 (.CK( clk ) , .Q( u2_L3_9 ) , .D( u2_R2_9 ) );
  DFF_X1 u2_L4_reg_1 (.CK( clk ) , .Q( u2_L4_1 ) , .D( u2_R3_1 ) );
  DFF_X1 u2_L4_reg_10 (.CK( clk ) , .Q( u2_L4_10 ) , .D( u2_R3_10 ) );
  DFF_X1 u2_L4_reg_11 (.CK( clk ) , .Q( u2_L4_11 ) , .D( u2_R3_11 ) );
  DFF_X1 u2_L4_reg_12 (.CK( clk ) , .Q( u2_L4_12 ) , .D( u2_R3_12 ) );
  DFF_X1 u2_L4_reg_13 (.CK( clk ) , .Q( u2_L4_13 ) , .D( u2_R3_13 ) );
  DFF_X1 u2_L4_reg_14 (.CK( clk ) , .Q( u2_L4_14 ) , .D( u2_R3_14 ) );
  DFF_X1 u2_L4_reg_15 (.CK( clk ) , .Q( u2_L4_15 ) , .D( u2_R3_15 ) );
  DFF_X1 u2_L4_reg_16 (.CK( clk ) , .Q( u2_L4_16 ) , .D( u2_R3_16 ) );
  DFF_X1 u2_L4_reg_17 (.CK( clk ) , .Q( u2_L4_17 ) , .D( u2_R3_17 ) );
  DFF_X1 u2_L4_reg_18 (.CK( clk ) , .Q( u2_L4_18 ) , .D( u2_R3_18 ) );
  DFF_X1 u2_L4_reg_19 (.CK( clk ) , .Q( u2_L4_19 ) , .D( u2_R3_19 ) );
  DFF_X1 u2_L4_reg_2 (.CK( clk ) , .Q( u2_L4_2 ) , .D( u2_R3_2 ) );
  DFF_X1 u2_L4_reg_20 (.CK( clk ) , .Q( u2_L4_20 ) , .D( u2_R3_20 ) );
  DFF_X1 u2_L4_reg_21 (.CK( clk ) , .Q( u2_L4_21 ) , .D( u2_R3_21 ) );
  DFF_X1 u2_L4_reg_22 (.CK( clk ) , .Q( u2_L4_22 ) , .D( u2_R3_22 ) );
  DFF_X1 u2_L4_reg_23 (.CK( clk ) , .Q( u2_L4_23 ) , .D( u2_R3_23 ) );
  DFF_X1 u2_L4_reg_24 (.CK( clk ) , .Q( u2_L4_24 ) , .D( u2_R3_24 ) );
  DFF_X1 u2_L4_reg_25 (.CK( clk ) , .Q( u2_L4_25 ) , .D( u2_R3_25 ) );
  DFF_X1 u2_L4_reg_26 (.CK( clk ) , .Q( u2_L4_26 ) , .D( u2_R3_26 ) );
  DFF_X1 u2_L4_reg_27 (.CK( clk ) , .Q( u2_L4_27 ) , .D( u2_R3_27 ) );
  DFF_X1 u2_L4_reg_28 (.CK( clk ) , .Q( u2_L4_28 ) , .D( u2_R3_28 ) );
  DFF_X1 u2_L4_reg_29 (.CK( clk ) , .Q( u2_L4_29 ) , .D( u2_R3_29 ) );
  DFF_X1 u2_L4_reg_3 (.CK( clk ) , .Q( u2_L4_3 ) , .D( u2_R3_3 ) );
  DFF_X1 u2_L4_reg_30 (.CK( clk ) , .Q( u2_L4_30 ) , .D( u2_R3_30 ) );
  DFF_X1 u2_L4_reg_31 (.CK( clk ) , .Q( u2_L4_31 ) , .D( u2_R3_31 ) );
  DFF_X1 u2_L4_reg_32 (.CK( clk ) , .Q( u2_L4_32 ) , .D( u2_R3_32 ) );
  DFF_X1 u2_L4_reg_4 (.CK( clk ) , .Q( u2_L4_4 ) , .D( u2_R3_4 ) );
  DFF_X1 u2_L4_reg_5 (.CK( clk ) , .Q( u2_L4_5 ) , .D( u2_R3_5 ) );
  DFF_X1 u2_L4_reg_6 (.CK( clk ) , .Q( u2_L4_6 ) , .D( u2_R3_6 ) );
  DFF_X1 u2_L4_reg_7 (.CK( clk ) , .Q( u2_L4_7 ) , .D( u2_R3_7 ) );
  DFF_X1 u2_L4_reg_8 (.CK( clk ) , .Q( u2_L4_8 ) , .D( u2_R3_8 ) );
  DFF_X1 u2_L4_reg_9 (.CK( clk ) , .Q( u2_L4_9 ) , .D( u2_R3_9 ) );
  DFF_X1 u2_L5_reg_1 (.CK( clk ) , .Q( u2_L5_1 ) , .D( u2_R4_1 ) );
  DFF_X1 u2_L5_reg_10 (.CK( clk ) , .Q( u2_L5_10 ) , .D( u2_R4_10 ) );
  DFF_X1 u2_L5_reg_11 (.CK( clk ) , .Q( u2_L5_11 ) , .D( u2_R4_11 ) );
  DFF_X1 u2_L5_reg_12 (.CK( clk ) , .Q( u2_L5_12 ) , .D( u2_R4_12 ) );
  DFF_X1 u2_L5_reg_13 (.CK( clk ) , .Q( u2_L5_13 ) , .D( u2_R4_13 ) );
  DFF_X1 u2_L5_reg_14 (.CK( clk ) , .Q( u2_L5_14 ) , .D( u2_R4_14 ) );
  DFF_X1 u2_L5_reg_15 (.CK( clk ) , .Q( u2_L5_15 ) , .D( u2_R4_15 ) );
  DFF_X1 u2_L5_reg_16 (.CK( clk ) , .Q( u2_L5_16 ) , .D( u2_R4_16 ) );
  DFF_X1 u2_L5_reg_17 (.CK( clk ) , .Q( u2_L5_17 ) , .D( u2_R4_17 ) );
  DFF_X1 u2_L5_reg_18 (.CK( clk ) , .Q( u2_L5_18 ) , .D( u2_R4_18 ) );
  DFF_X1 u2_L5_reg_19 (.CK( clk ) , .Q( u2_L5_19 ) , .D( u2_R4_19 ) );
  DFF_X1 u2_L5_reg_2 (.CK( clk ) , .Q( u2_L5_2 ) , .D( u2_R4_2 ) );
  DFF_X1 u2_L5_reg_20 (.CK( clk ) , .Q( u2_L5_20 ) , .D( u2_R4_20 ) );
  DFF_X1 u2_L5_reg_21 (.CK( clk ) , .Q( u2_L5_21 ) , .D( u2_R4_21 ) );
  DFF_X1 u2_L5_reg_22 (.CK( clk ) , .Q( u2_L5_22 ) , .D( u2_R4_22 ) );
  DFF_X1 u2_L5_reg_23 (.CK( clk ) , .Q( u2_L5_23 ) , .D( u2_R4_23 ) );
  DFF_X1 u2_L5_reg_24 (.CK( clk ) , .Q( u2_L5_24 ) , .D( u2_R4_24 ) );
  DFF_X1 u2_L5_reg_25 (.CK( clk ) , .Q( u2_L5_25 ) , .D( u2_R4_25 ) );
  DFF_X1 u2_L5_reg_26 (.CK( clk ) , .Q( u2_L5_26 ) , .D( u2_R4_26 ) );
  DFF_X1 u2_L5_reg_27 (.CK( clk ) , .Q( u2_L5_27 ) , .D( u2_R4_27 ) );
  DFF_X1 u2_L5_reg_28 (.CK( clk ) , .Q( u2_L5_28 ) , .D( u2_R4_28 ) );
  DFF_X1 u2_L5_reg_29 (.CK( clk ) , .Q( u2_L5_29 ) , .D( u2_R4_29 ) );
  DFF_X1 u2_L5_reg_3 (.CK( clk ) , .Q( u2_L5_3 ) , .D( u2_R4_3 ) );
  DFF_X1 u2_L5_reg_30 (.CK( clk ) , .Q( u2_L5_30 ) , .D( u2_R4_30 ) );
  DFF_X1 u2_L5_reg_31 (.CK( clk ) , .Q( u2_L5_31 ) , .D( u2_R4_31 ) );
  DFF_X1 u2_L5_reg_32 (.CK( clk ) , .Q( u2_L5_32 ) , .D( u2_R4_32 ) );
  DFF_X1 u2_L5_reg_4 (.CK( clk ) , .Q( u2_L5_4 ) , .D( u2_R4_4 ) );
  DFF_X1 u2_L5_reg_5 (.CK( clk ) , .Q( u2_L5_5 ) , .D( u2_R4_5 ) );
  DFF_X1 u2_L5_reg_6 (.CK( clk ) , .Q( u2_L5_6 ) , .D( u2_R4_6 ) );
  DFF_X1 u2_L5_reg_7 (.CK( clk ) , .Q( u2_L5_7 ) , .D( u2_R4_7 ) );
  DFF_X1 u2_L5_reg_8 (.CK( clk ) , .Q( u2_L5_8 ) , .D( u2_R4_8 ) );
  DFF_X1 u2_L5_reg_9 (.CK( clk ) , .Q( u2_L5_9 ) , .D( u2_R4_9 ) );
  DFF_X1 u2_L6_reg_1 (.CK( clk ) , .Q( u2_L6_1 ) , .D( u2_R5_1 ) );
  DFF_X1 u2_L6_reg_10 (.CK( clk ) , .Q( u2_L6_10 ) , .D( u2_R5_10 ) );
  DFF_X1 u2_L6_reg_11 (.CK( clk ) , .Q( u2_L6_11 ) , .D( u2_R5_11 ) );
  DFF_X1 u2_L6_reg_12 (.CK( clk ) , .Q( u2_L6_12 ) , .D( u2_R5_12 ) );
  DFF_X1 u2_L6_reg_13 (.CK( clk ) , .Q( u2_L6_13 ) , .D( u2_R5_13 ) );
  DFF_X1 u2_L6_reg_14 (.CK( clk ) , .Q( u2_L6_14 ) , .D( u2_R5_14 ) );
  DFF_X1 u2_L6_reg_15 (.CK( clk ) , .Q( u2_L6_15 ) , .D( u2_R5_15 ) );
  DFF_X1 u2_L6_reg_16 (.CK( clk ) , .Q( u2_L6_16 ) , .D( u2_R5_16 ) );
  DFF_X1 u2_L6_reg_17 (.CK( clk ) , .Q( u2_L6_17 ) , .D( u2_R5_17 ) );
  DFF_X1 u2_L6_reg_18 (.CK( clk ) , .Q( u2_L6_18 ) , .D( u2_R5_18 ) );
  DFF_X1 u2_L6_reg_19 (.CK( clk ) , .Q( u2_L6_19 ) , .D( u2_R5_19 ) );
  DFF_X1 u2_L6_reg_2 (.CK( clk ) , .Q( u2_L6_2 ) , .D( u2_R5_2 ) );
  DFF_X1 u2_L6_reg_20 (.CK( clk ) , .Q( u2_L6_20 ) , .D( u2_R5_20 ) );
  DFF_X1 u2_L6_reg_21 (.CK( clk ) , .Q( u2_L6_21 ) , .D( u2_R5_21 ) );
  DFF_X1 u2_L6_reg_22 (.CK( clk ) , .Q( u2_L6_22 ) , .D( u2_R5_22 ) );
  DFF_X1 u2_L6_reg_23 (.CK( clk ) , .Q( u2_L6_23 ) , .D( u2_R5_23 ) );
  DFF_X1 u2_L6_reg_24 (.CK( clk ) , .Q( u2_L6_24 ) , .D( u2_R5_24 ) );
  DFF_X1 u2_L6_reg_25 (.CK( clk ) , .Q( u2_L6_25 ) , .D( u2_R5_25 ) );
  DFF_X1 u2_L6_reg_26 (.CK( clk ) , .Q( u2_L6_26 ) , .D( u2_R5_26 ) );
  DFF_X1 u2_L6_reg_27 (.CK( clk ) , .Q( u2_L6_27 ) , .D( u2_R5_27 ) );
  DFF_X1 u2_L6_reg_28 (.CK( clk ) , .Q( u2_L6_28 ) , .D( u2_R5_28 ) );
  DFF_X1 u2_L6_reg_29 (.CK( clk ) , .Q( u2_L6_29 ) , .D( u2_R5_29 ) );
  DFF_X1 u2_L6_reg_3 (.CK( clk ) , .Q( u2_L6_3 ) , .D( u2_R5_3 ) );
  DFF_X1 u2_L6_reg_30 (.CK( clk ) , .Q( u2_L6_30 ) , .D( u2_R5_30 ) );
  DFF_X1 u2_L6_reg_31 (.CK( clk ) , .Q( u2_L6_31 ) , .D( u2_R5_31 ) );
  DFF_X1 u2_L6_reg_32 (.CK( clk ) , .Q( u2_L6_32 ) , .D( u2_R5_32 ) );
  DFF_X1 u2_L6_reg_4 (.CK( clk ) , .Q( u2_L6_4 ) , .D( u2_R5_4 ) );
  DFF_X1 u2_L6_reg_5 (.CK( clk ) , .Q( u2_L6_5 ) , .D( u2_R5_5 ) );
  DFF_X1 u2_L6_reg_6 (.CK( clk ) , .Q( u2_L6_6 ) , .D( u2_R5_6 ) );
  DFF_X1 u2_L6_reg_7 (.CK( clk ) , .Q( u2_L6_7 ) , .D( u2_R5_7 ) );
  DFF_X1 u2_L6_reg_8 (.CK( clk ) , .Q( u2_L6_8 ) , .D( u2_R5_8 ) );
  DFF_X1 u2_L6_reg_9 (.CK( clk ) , .Q( u2_L6_9 ) , .D( u2_R5_9 ) );
  DFF_X1 u2_L7_reg_1 (.CK( clk ) , .Q( u2_L7_1 ) , .D( u2_R6_1 ) );
  DFF_X1 u2_L7_reg_10 (.CK( clk ) , .Q( u2_L7_10 ) , .D( u2_R6_10 ) );
  DFF_X1 u2_L7_reg_11 (.CK( clk ) , .Q( u2_L7_11 ) , .D( u2_R6_11 ) );
  DFF_X1 u2_L7_reg_12 (.CK( clk ) , .Q( u2_L7_12 ) , .D( u2_R6_12 ) );
  DFF_X1 u2_L7_reg_13 (.CK( clk ) , .Q( u2_L7_13 ) , .D( u2_R6_13 ) );
  DFF_X1 u2_L7_reg_14 (.CK( clk ) , .Q( u2_L7_14 ) , .D( u2_R6_14 ) );
  DFF_X1 u2_L7_reg_15 (.CK( clk ) , .Q( u2_L7_15 ) , .D( u2_R6_15 ) );
  DFF_X1 u2_L7_reg_16 (.CK( clk ) , .Q( u2_L7_16 ) , .D( u2_R6_16 ) );
  DFF_X1 u2_L7_reg_17 (.CK( clk ) , .Q( u2_L7_17 ) , .D( u2_R6_17 ) );
  DFF_X1 u2_L7_reg_18 (.CK( clk ) , .Q( u2_L7_18 ) , .D( u2_R6_18 ) );
  DFF_X1 u2_L7_reg_19 (.CK( clk ) , .Q( u2_L7_19 ) , .D( u2_R6_19 ) );
  DFF_X1 u2_L7_reg_2 (.CK( clk ) , .Q( u2_L7_2 ) , .D( u2_R6_2 ) );
  DFF_X1 u2_L7_reg_20 (.CK( clk ) , .Q( u2_L7_20 ) , .D( u2_R6_20 ) );
  DFF_X1 u2_L7_reg_21 (.CK( clk ) , .Q( u2_L7_21 ) , .D( u2_R6_21 ) );
  DFF_X1 u2_L7_reg_22 (.CK( clk ) , .Q( u2_L7_22 ) , .D( u2_R6_22 ) );
  DFF_X1 u2_L7_reg_23 (.CK( clk ) , .Q( u2_L7_23 ) , .D( u2_R6_23 ) );
  DFF_X1 u2_L7_reg_24 (.CK( clk ) , .Q( u2_L7_24 ) , .D( u2_R6_24 ) );
  DFF_X1 u2_L7_reg_25 (.CK( clk ) , .Q( u2_L7_25 ) , .D( u2_R6_25 ) );
  DFF_X1 u2_L7_reg_26 (.CK( clk ) , .Q( u2_L7_26 ) , .D( u2_R6_26 ) );
  DFF_X1 u2_L7_reg_27 (.CK( clk ) , .Q( u2_L7_27 ) , .D( u2_R6_27 ) );
  DFF_X1 u2_L7_reg_28 (.CK( clk ) , .Q( u2_L7_28 ) , .D( u2_R6_28 ) );
  DFF_X1 u2_L7_reg_29 (.CK( clk ) , .Q( u2_L7_29 ) , .D( u2_R6_29 ) );
  DFF_X1 u2_L7_reg_3 (.CK( clk ) , .Q( u2_L7_3 ) , .D( u2_R6_3 ) );
  DFF_X1 u2_L7_reg_30 (.CK( clk ) , .Q( u2_L7_30 ) , .D( u2_R6_30 ) );
  DFF_X1 u2_L7_reg_31 (.CK( clk ) , .Q( u2_L7_31 ) , .D( u2_R6_31 ) );
  DFF_X1 u2_L7_reg_32 (.CK( clk ) , .Q( u2_L7_32 ) , .D( u2_R6_32 ) );
  DFF_X1 u2_L7_reg_4 (.CK( clk ) , .Q( u2_L7_4 ) , .D( u2_R6_4 ) );
  DFF_X1 u2_L7_reg_5 (.CK( clk ) , .Q( u2_L7_5 ) , .D( u2_R6_5 ) );
  DFF_X1 u2_L7_reg_6 (.CK( clk ) , .Q( u2_L7_6 ) , .D( u2_R6_6 ) );
  DFF_X1 u2_L7_reg_7 (.CK( clk ) , .Q( u2_L7_7 ) , .D( u2_R6_7 ) );
  DFF_X1 u2_L7_reg_8 (.CK( clk ) , .Q( u2_L7_8 ) , .D( u2_R6_8 ) );
  DFF_X1 u2_L7_reg_9 (.CK( clk ) , .Q( u2_L7_9 ) , .D( u2_R6_9 ) );
  DFF_X1 u2_L8_reg_1 (.CK( clk ) , .Q( u2_L8_1 ) , .D( u2_R7_1 ) );
  DFF_X1 u2_L8_reg_10 (.CK( clk ) , .Q( u2_L8_10 ) , .D( u2_R7_10 ) );
  DFF_X1 u2_L8_reg_11 (.CK( clk ) , .Q( u2_L8_11 ) , .D( u2_R7_11 ) );
  DFF_X1 u2_L8_reg_12 (.CK( clk ) , .Q( u2_L8_12 ) , .D( u2_R7_12 ) );
  DFF_X1 u2_L8_reg_13 (.CK( clk ) , .Q( u2_L8_13 ) , .D( u2_R7_13 ) );
  DFF_X1 u2_L8_reg_14 (.CK( clk ) , .Q( u2_L8_14 ) , .D( u2_R7_14 ) );
  DFF_X1 u2_L8_reg_15 (.CK( clk ) , .Q( u2_L8_15 ) , .D( u2_R7_15 ) );
  DFF_X1 u2_L8_reg_16 (.CK( clk ) , .Q( u2_L8_16 ) , .D( u2_R7_16 ) );
  DFF_X1 u2_L8_reg_17 (.CK( clk ) , .Q( u2_L8_17 ) , .D( u2_R7_17 ) );
  DFF_X1 u2_L8_reg_18 (.CK( clk ) , .Q( u2_L8_18 ) , .D( u2_R7_18 ) );
  DFF_X1 u2_L8_reg_19 (.CK( clk ) , .Q( u2_L8_19 ) , .D( u2_R7_19 ) );
  DFF_X1 u2_L8_reg_2 (.CK( clk ) , .Q( u2_L8_2 ) , .D( u2_R7_2 ) );
  DFF_X1 u2_L8_reg_20 (.CK( clk ) , .Q( u2_L8_20 ) , .D( u2_R7_20 ) );
  DFF_X1 u2_L8_reg_21 (.CK( clk ) , .Q( u2_L8_21 ) , .D( u2_R7_21 ) );
  DFF_X1 u2_L8_reg_22 (.CK( clk ) , .Q( u2_L8_22 ) , .D( u2_R7_22 ) );
  DFF_X1 u2_L8_reg_23 (.CK( clk ) , .Q( u2_L8_23 ) , .D( u2_R7_23 ) );
  DFF_X1 u2_L8_reg_24 (.CK( clk ) , .Q( u2_L8_24 ) , .D( u2_R7_24 ) );
  DFF_X1 u2_L8_reg_25 (.CK( clk ) , .Q( u2_L8_25 ) , .D( u2_R7_25 ) );
  DFF_X1 u2_L8_reg_26 (.CK( clk ) , .Q( u2_L8_26 ) , .D( u2_R7_26 ) );
  DFF_X1 u2_L8_reg_27 (.CK( clk ) , .Q( u2_L8_27 ) , .D( u2_R7_27 ) );
  DFF_X1 u2_L8_reg_28 (.CK( clk ) , .Q( u2_L8_28 ) , .D( u2_R7_28 ) );
  DFF_X1 u2_L8_reg_29 (.CK( clk ) , .Q( u2_L8_29 ) , .D( u2_R7_29 ) );
  DFF_X1 u2_L8_reg_3 (.CK( clk ) , .Q( u2_L8_3 ) , .D( u2_R7_3 ) );
  DFF_X1 u2_L8_reg_30 (.CK( clk ) , .Q( u2_L8_30 ) , .D( u2_R7_30 ) );
  DFF_X1 u2_L8_reg_31 (.CK( clk ) , .Q( u2_L8_31 ) , .D( u2_R7_31 ) );
  DFF_X1 u2_L8_reg_32 (.CK( clk ) , .Q( u2_L8_32 ) , .D( u2_R7_32 ) );
  DFF_X1 u2_L8_reg_4 (.CK( clk ) , .Q( u2_L8_4 ) , .D( u2_R7_4 ) );
  DFF_X1 u2_L8_reg_5 (.CK( clk ) , .Q( u2_L8_5 ) , .D( u2_R7_5 ) );
  DFF_X1 u2_L8_reg_6 (.CK( clk ) , .Q( u2_L8_6 ) , .D( u2_R7_6 ) );
  DFF_X1 u2_L8_reg_7 (.CK( clk ) , .Q( u2_L8_7 ) , .D( u2_R7_7 ) );
  DFF_X1 u2_L8_reg_8 (.CK( clk ) , .Q( u2_L8_8 ) , .D( u2_R7_8 ) );
  DFF_X1 u2_L8_reg_9 (.CK( clk ) , .Q( u2_L8_9 ) , .D( u2_R7_9 ) );
  DFF_X1 u2_L9_reg_1 (.CK( clk ) , .Q( u2_L9_1 ) , .D( u2_R8_1 ) );
  DFF_X1 u2_L9_reg_10 (.CK( clk ) , .Q( u2_L9_10 ) , .D( u2_R8_10 ) );
  DFF_X1 u2_L9_reg_11 (.CK( clk ) , .Q( u2_L9_11 ) , .D( u2_R8_11 ) );
  DFF_X1 u2_L9_reg_12 (.CK( clk ) , .Q( u2_L9_12 ) , .D( u2_R8_12 ) );
  DFF_X1 u2_L9_reg_13 (.CK( clk ) , .Q( u2_L9_13 ) , .D( u2_R8_13 ) );
  DFF_X1 u2_L9_reg_14 (.CK( clk ) , .Q( u2_L9_14 ) , .D( u2_R8_14 ) );
  DFF_X1 u2_L9_reg_15 (.CK( clk ) , .Q( u2_L9_15 ) , .D( u2_R8_15 ) );
  DFF_X1 u2_L9_reg_16 (.CK( clk ) , .Q( u2_L9_16 ) , .D( u2_R8_16 ) );
  DFF_X1 u2_L9_reg_17 (.CK( clk ) , .Q( u2_L9_17 ) , .D( u2_R8_17 ) );
  DFF_X1 u2_L9_reg_18 (.CK( clk ) , .Q( u2_L9_18 ) , .D( u2_R8_18 ) );
  DFF_X1 u2_L9_reg_19 (.CK( clk ) , .Q( u2_L9_19 ) , .D( u2_R8_19 ) );
  DFF_X1 u2_L9_reg_2 (.CK( clk ) , .Q( u2_L9_2 ) , .D( u2_R8_2 ) );
  DFF_X1 u2_L9_reg_20 (.CK( clk ) , .Q( u2_L9_20 ) , .D( u2_R8_20 ) );
  DFF_X1 u2_L9_reg_21 (.CK( clk ) , .Q( u2_L9_21 ) , .D( u2_R8_21 ) );
  DFF_X1 u2_L9_reg_22 (.CK( clk ) , .Q( u2_L9_22 ) , .D( u2_R8_22 ) );
  DFF_X1 u2_L9_reg_23 (.CK( clk ) , .Q( u2_L9_23 ) , .D( u2_R8_23 ) );
  DFF_X1 u2_L9_reg_24 (.CK( clk ) , .Q( u2_L9_24 ) , .D( u2_R8_24 ) );
  DFF_X1 u2_L9_reg_25 (.CK( clk ) , .Q( u2_L9_25 ) , .D( u2_R8_25 ) );
  DFF_X1 u2_L9_reg_26 (.CK( clk ) , .Q( u2_L9_26 ) , .D( u2_R8_26 ) );
  DFF_X1 u2_L9_reg_27 (.CK( clk ) , .Q( u2_L9_27 ) , .D( u2_R8_27 ) );
  DFF_X1 u2_L9_reg_28 (.CK( clk ) , .Q( u2_L9_28 ) , .D( u2_R8_28 ) );
  DFF_X1 u2_L9_reg_29 (.CK( clk ) , .Q( u2_L9_29 ) , .D( u2_R8_29 ) );
  DFF_X1 u2_L9_reg_3 (.CK( clk ) , .Q( u2_L9_3 ) , .D( u2_R8_3 ) );
  DFF_X1 u2_L9_reg_30 (.CK( clk ) , .Q( u2_L9_30 ) , .D( u2_R8_30 ) );
  DFF_X1 u2_L9_reg_31 (.CK( clk ) , .Q( u2_L9_31 ) , .D( u2_R8_31 ) );
  DFF_X1 u2_L9_reg_32 (.CK( clk ) , .Q( u2_L9_32 ) , .D( u2_R8_32 ) );
  DFF_X1 u2_L9_reg_4 (.CK( clk ) , .Q( u2_L9_4 ) , .D( u2_R8_4 ) );
  DFF_X1 u2_L9_reg_5 (.CK( clk ) , .Q( u2_L9_5 ) , .D( u2_R8_5 ) );
  DFF_X1 u2_L9_reg_6 (.CK( clk ) , .Q( u2_L9_6 ) , .D( u2_R8_6 ) );
  DFF_X1 u2_L9_reg_7 (.CK( clk ) , .Q( u2_L9_7 ) , .D( u2_R8_7 ) );
  DFF_X1 u2_L9_reg_8 (.CK( clk ) , .Q( u2_L9_8 ) , .D( u2_R8_8 ) );
  DFF_X1 u2_L9_reg_9 (.CK( clk ) , .Q( u2_L9_9 ) , .D( u2_R8_9 ) );
  DFF_X1 u2_R0_reg_1 (.CK( clk ) , .D( u2_N0 ) , .Q( u2_R0_1 ) );
  DFF_X1 u2_R0_reg_10 (.CK( clk ) , .D( u2_N9 ) , .Q( u2_R0_10 ) );
  DFF_X1 u2_R0_reg_11 (.CK( clk ) , .D( u2_N10 ) , .Q( u2_R0_11 ) );
  DFF_X1 u2_R0_reg_12 (.CK( clk ) , .D( u2_N11 ) , .Q( u2_R0_12 ) );
  DFF_X1 u2_R0_reg_13 (.CK( clk ) , .D( u2_N12 ) , .Q( u2_R0_13 ) );
  DFF_X1 u2_R0_reg_14 (.CK( clk ) , .D( u2_N13 ) , .Q( u2_R0_14 ) );
  DFF_X1 u2_R0_reg_15 (.CK( clk ) , .D( u2_N14 ) , .Q( u2_R0_15 ) );
  DFF_X1 u2_R0_reg_16 (.CK( clk ) , .D( u2_N15 ) , .Q( u2_R0_16 ) );
  DFF_X1 u2_R0_reg_17 (.CK( clk ) , .D( u2_N16 ) , .Q( u2_R0_17 ) );
  DFF_X1 u2_R0_reg_18 (.CK( clk ) , .D( u2_N17 ) , .Q( u2_R0_18 ) );
  DFF_X1 u2_R0_reg_19 (.CK( clk ) , .D( u2_N18 ) , .Q( u2_R0_19 ) );
  DFF_X1 u2_R0_reg_2 (.CK( clk ) , .D( u2_N1 ) , .Q( u2_R0_2 ) );
  DFF_X1 u2_R0_reg_20 (.CK( clk ) , .D( u2_N19 ) , .Q( u2_R0_20 ) );
  DFF_X1 u2_R0_reg_21 (.CK( clk ) , .D( u2_N20 ) , .Q( u2_R0_21 ) );
  DFF_X1 u2_R0_reg_22 (.CK( clk ) , .D( u2_N21 ) , .Q( u2_R0_22 ) );
  DFF_X1 u2_R0_reg_23 (.CK( clk ) , .D( u2_N22 ) , .Q( u2_R0_23 ) );
  DFF_X1 u2_R0_reg_24 (.CK( clk ) , .D( u2_N23 ) , .Q( u2_R0_24 ) );
  DFF_X1 u2_R0_reg_25 (.CK( clk ) , .D( u2_N24 ) , .Q( u2_R0_25 ) );
  DFF_X1 u2_R0_reg_26 (.CK( clk ) , .D( u2_N25 ) , .Q( u2_R0_26 ) );
  DFF_X1 u2_R0_reg_27 (.CK( clk ) , .D( u2_N26 ) , .Q( u2_R0_27 ) );
  DFF_X1 u2_R0_reg_28 (.CK( clk ) , .D( u2_N27 ) , .Q( u2_R0_28 ) );
  DFF_X1 u2_R0_reg_29 (.CK( clk ) , .D( u2_N28 ) , .Q( u2_R0_29 ) );
  DFF_X1 u2_R0_reg_3 (.CK( clk ) , .D( u2_N2 ) , .Q( u2_R0_3 ) );
  DFF_X1 u2_R0_reg_30 (.CK( clk ) , .D( u2_N29 ) , .Q( u2_R0_30 ) );
  DFF_X1 u2_R0_reg_31 (.CK( clk ) , .D( u2_N30 ) , .Q( u2_R0_31 ) );
  DFF_X1 u2_R0_reg_32 (.CK( clk ) , .D( u2_N31 ) , .Q( u2_R0_32 ) );
  DFF_X1 u2_R0_reg_4 (.CK( clk ) , .D( u2_N3 ) , .Q( u2_R0_4 ) );
  DFF_X1 u2_R0_reg_5 (.CK( clk ) , .D( u2_N4 ) , .Q( u2_R0_5 ) );
  DFF_X1 u2_R0_reg_6 (.CK( clk ) , .D( u2_N5 ) , .Q( u2_R0_6 ) );
  DFF_X1 u2_R0_reg_7 (.CK( clk ) , .D( u2_N6 ) , .Q( u2_R0_7 ) );
  DFF_X1 u2_R0_reg_8 (.CK( clk ) , .D( u2_N7 ) , .Q( u2_R0_8 ) );
  DFF_X1 u2_R0_reg_9 (.CK( clk ) , .D( u2_N8 ) , .Q( u2_R0_9 ) );
  DFF_X1 u2_R10_reg_1 (.CK( clk ) , .D( u2_N320 ) , .Q( u2_R10_1 ) );
  DFF_X1 u2_R10_reg_10 (.CK( clk ) , .D( u2_N329 ) , .Q( u2_R10_10 ) );
  DFF_X1 u2_R10_reg_11 (.CK( clk ) , .D( u2_N330 ) , .Q( u2_R10_11 ) );
  DFF_X1 u2_R10_reg_12 (.CK( clk ) , .D( u2_N331 ) , .Q( u2_R10_12 ) );
  DFF_X1 u2_R10_reg_13 (.CK( clk ) , .D( u2_N332 ) , .Q( u2_R10_13 ) );
  DFF_X1 u2_R10_reg_14 (.CK( clk ) , .D( u2_N333 ) , .Q( u2_R10_14 ) );
  DFF_X1 u2_R10_reg_15 (.CK( clk ) , .D( u2_N334 ) , .Q( u2_R10_15 ) );
  DFF_X1 u2_R10_reg_16 (.CK( clk ) , .D( u2_N335 ) , .Q( u2_R10_16 ) );
  DFF_X1 u2_R10_reg_17 (.CK( clk ) , .D( u2_N336 ) , .Q( u2_R10_17 ) );
  DFF_X1 u2_R10_reg_18 (.CK( clk ) , .D( u2_N337 ) , .Q( u2_R10_18 ) );
  DFF_X1 u2_R10_reg_19 (.CK( clk ) , .D( u2_N338 ) , .Q( u2_R10_19 ) );
  DFF_X1 u2_R10_reg_2 (.CK( clk ) , .D( u2_N321 ) , .Q( u2_R10_2 ) );
  DFF_X1 u2_R10_reg_20 (.CK( clk ) , .D( u2_N339 ) , .Q( u2_R10_20 ) );
  DFF_X1 u2_R10_reg_21 (.CK( clk ) , .D( u2_N340 ) , .Q( u2_R10_21 ) );
  DFF_X1 u2_R10_reg_22 (.CK( clk ) , .D( u2_N341 ) , .Q( u2_R10_22 ) );
  DFF_X1 u2_R10_reg_23 (.CK( clk ) , .D( u2_N342 ) , .Q( u2_R10_23 ) );
  DFF_X1 u2_R10_reg_24 (.CK( clk ) , .D( u2_N343 ) , .Q( u2_R10_24 ) );
  DFF_X1 u2_R10_reg_25 (.CK( clk ) , .D( u2_N344 ) , .Q( u2_R10_25 ) );
  DFF_X1 u2_R10_reg_26 (.CK( clk ) , .D( u2_N345 ) , .Q( u2_R10_26 ) );
  DFF_X1 u2_R10_reg_27 (.CK( clk ) , .D( u2_N346 ) , .Q( u2_R10_27 ) );
  DFF_X1 u2_R10_reg_28 (.CK( clk ) , .D( u2_N347 ) , .Q( u2_R10_28 ) );
  DFF_X1 u2_R10_reg_29 (.CK( clk ) , .D( u2_N348 ) , .Q( u2_R10_29 ) );
  DFF_X1 u2_R10_reg_3 (.CK( clk ) , .D( u2_N322 ) , .Q( u2_R10_3 ) );
  DFF_X1 u2_R10_reg_30 (.CK( clk ) , .D( u2_N349 ) , .Q( u2_R10_30 ) );
  DFF_X1 u2_R10_reg_31 (.CK( clk ) , .D( u2_N350 ) , .Q( u2_R10_31 ) );
  DFF_X1 u2_R10_reg_32 (.CK( clk ) , .D( u2_N351 ) , .Q( u2_R10_32 ) );
  DFF_X1 u2_R10_reg_4 (.CK( clk ) , .D( u2_N323 ) , .Q( u2_R10_4 ) );
  DFF_X1 u2_R10_reg_5 (.CK( clk ) , .D( u2_N324 ) , .Q( u2_R10_5 ) );
  DFF_X1 u2_R10_reg_6 (.CK( clk ) , .D( u2_N325 ) , .Q( u2_R10_6 ) );
  DFF_X1 u2_R10_reg_7 (.CK( clk ) , .D( u2_N326 ) , .Q( u2_R10_7 ) );
  DFF_X1 u2_R10_reg_8 (.CK( clk ) , .D( u2_N327 ) , .Q( u2_R10_8 ) );
  DFF_X1 u2_R10_reg_9 (.CK( clk ) , .D( u2_N328 ) , .Q( u2_R10_9 ) );
  DFF_X1 u2_R11_reg_1 (.CK( clk ) , .D( u2_N352 ) , .Q( u2_R11_1 ) );
  DFF_X1 u2_R11_reg_10 (.CK( clk ) , .D( u2_N361 ) , .Q( u2_R11_10 ) );
  DFF_X1 u2_R11_reg_11 (.CK( clk ) , .D( u2_N362 ) , .Q( u2_R11_11 ) );
  DFF_X1 u2_R11_reg_12 (.CK( clk ) , .D( u2_N363 ) , .Q( u2_R11_12 ) );
  DFF_X1 u2_R11_reg_13 (.CK( clk ) , .D( u2_N364 ) , .Q( u2_R11_13 ) );
  DFF_X1 u2_R11_reg_14 (.CK( clk ) , .D( u2_N365 ) , .Q( u2_R11_14 ) );
  DFF_X1 u2_R11_reg_15 (.CK( clk ) , .D( u2_N366 ) , .Q( u2_R11_15 ) );
  DFF_X1 u2_R11_reg_16 (.CK( clk ) , .D( u2_N367 ) , .Q( u2_R11_16 ) );
  DFF_X1 u2_R11_reg_17 (.CK( clk ) , .D( u2_N368 ) , .Q( u2_R11_17 ) );
  DFF_X1 u2_R11_reg_18 (.CK( clk ) , .D( u2_N369 ) , .Q( u2_R11_18 ) );
  DFF_X1 u2_R11_reg_19 (.CK( clk ) , .D( u2_N370 ) , .Q( u2_R11_19 ) );
  DFF_X1 u2_R11_reg_2 (.CK( clk ) , .D( u2_N353 ) , .Q( u2_R11_2 ) );
  DFF_X1 u2_R11_reg_20 (.CK( clk ) , .D( u2_N371 ) , .Q( u2_R11_20 ) );
  DFF_X1 u2_R11_reg_21 (.CK( clk ) , .D( u2_N372 ) , .Q( u2_R11_21 ) );
  DFF_X1 u2_R11_reg_22 (.CK( clk ) , .D( u2_N373 ) , .Q( u2_R11_22 ) );
  DFF_X1 u2_R11_reg_23 (.CK( clk ) , .D( u2_N374 ) , .Q( u2_R11_23 ) );
  DFF_X1 u2_R11_reg_24 (.CK( clk ) , .D( u2_N375 ) , .Q( u2_R11_24 ) );
  DFF_X1 u2_R11_reg_25 (.CK( clk ) , .D( u2_N376 ) , .Q( u2_R11_25 ) );
  DFF_X1 u2_R11_reg_26 (.CK( clk ) , .D( u2_N377 ) , .Q( u2_R11_26 ) );
  DFF_X1 u2_R11_reg_27 (.CK( clk ) , .D( u2_N378 ) , .Q( u2_R11_27 ) );
  DFF_X1 u2_R11_reg_28 (.CK( clk ) , .D( u2_N379 ) , .Q( u2_R11_28 ) );
  DFF_X1 u2_R11_reg_29 (.CK( clk ) , .D( u2_N380 ) , .Q( u2_R11_29 ) );
  DFF_X1 u2_R11_reg_3 (.CK( clk ) , .D( u2_N354 ) , .Q( u2_R11_3 ) );
  DFF_X1 u2_R11_reg_30 (.CK( clk ) , .D( u2_N381 ) , .Q( u2_R11_30 ) );
  DFF_X1 u2_R11_reg_31 (.CK( clk ) , .D( u2_N382 ) , .Q( u2_R11_31 ) );
  DFF_X1 u2_R11_reg_32 (.CK( clk ) , .D( u2_N383 ) , .Q( u2_R11_32 ) );
  DFF_X1 u2_R11_reg_4 (.CK( clk ) , .D( u2_N355 ) , .Q( u2_R11_4 ) );
  DFF_X1 u2_R11_reg_5 (.CK( clk ) , .D( u2_N356 ) , .Q( u2_R11_5 ) );
  DFF_X1 u2_R11_reg_6 (.CK( clk ) , .D( u2_N357 ) , .Q( u2_R11_6 ) );
  DFF_X1 u2_R11_reg_7 (.CK( clk ) , .D( u2_N358 ) , .Q( u2_R11_7 ) );
  DFF_X1 u2_R11_reg_8 (.CK( clk ) , .D( u2_N359 ) , .Q( u2_R11_8 ) );
  DFF_X1 u2_R11_reg_9 (.CK( clk ) , .D( u2_N360 ) , .Q( u2_R11_9 ) );
  DFF_X1 u2_R12_reg_1 (.CK( clk ) , .D( u2_N384 ) , .Q( u2_R12_1 ) );
  DFF_X1 u2_R12_reg_10 (.CK( clk ) , .D( u2_N393 ) , .Q( u2_R12_10 ) );
  DFF_X1 u2_R12_reg_11 (.CK( clk ) , .D( u2_N394 ) , .Q( u2_R12_11 ) );
  DFF_X1 u2_R12_reg_12 (.CK( clk ) , .D( u2_N395 ) , .Q( u2_R12_12 ) );
  DFF_X1 u2_R12_reg_13 (.CK( clk ) , .D( u2_N396 ) , .Q( u2_R12_13 ) );
  DFF_X1 u2_R12_reg_14 (.CK( clk ) , .D( u2_N397 ) , .Q( u2_R12_14 ) );
  DFF_X1 u2_R12_reg_15 (.CK( clk ) , .D( u2_N398 ) , .Q( u2_R12_15 ) );
  DFF_X1 u2_R12_reg_16 (.CK( clk ) , .D( u2_N399 ) , .Q( u2_R12_16 ) );
  DFF_X1 u2_R12_reg_17 (.CK( clk ) , .D( u2_N400 ) , .Q( u2_R12_17 ) );
  DFF_X1 u2_R12_reg_18 (.CK( clk ) , .D( u2_N401 ) , .Q( u2_R12_18 ) );
  DFF_X1 u2_R12_reg_19 (.CK( clk ) , .D( u2_N402 ) , .Q( u2_R12_19 ) );
  DFF_X1 u2_R12_reg_2 (.CK( clk ) , .D( u2_N385 ) , .Q( u2_R12_2 ) );
  DFF_X1 u2_R12_reg_20 (.CK( clk ) , .D( u2_N403 ) , .Q( u2_R12_20 ) );
  DFF_X1 u2_R12_reg_21 (.CK( clk ) , .D( u2_N404 ) , .Q( u2_R12_21 ) );
  DFF_X1 u2_R12_reg_22 (.CK( clk ) , .D( u2_N405 ) , .Q( u2_R12_22 ) );
  DFF_X1 u2_R12_reg_23 (.CK( clk ) , .D( u2_N406 ) , .Q( u2_R12_23 ) );
  DFF_X1 u2_R12_reg_24 (.CK( clk ) , .D( u2_N407 ) , .Q( u2_R12_24 ) );
  DFF_X1 u2_R12_reg_25 (.CK( clk ) , .D( u2_N408 ) , .Q( u2_R12_25 ) );
  DFF_X1 u2_R12_reg_26 (.CK( clk ) , .D( u2_N409 ) , .Q( u2_R12_26 ) );
  DFF_X1 u2_R12_reg_27 (.CK( clk ) , .D( u2_N410 ) , .Q( u2_R12_27 ) );
  DFF_X1 u2_R12_reg_28 (.CK( clk ) , .D( u2_N411 ) , .Q( u2_R12_28 ) );
  DFF_X1 u2_R12_reg_29 (.CK( clk ) , .D( u2_N412 ) , .Q( u2_R12_29 ) );
  DFF_X1 u2_R12_reg_3 (.CK( clk ) , .D( u2_N386 ) , .Q( u2_R12_3 ) );
  DFF_X1 u2_R12_reg_30 (.CK( clk ) , .D( u2_N413 ) , .Q( u2_R12_30 ) );
  DFF_X1 u2_R12_reg_31 (.CK( clk ) , .D( u2_N414 ) , .Q( u2_R12_31 ) );
  DFF_X1 u2_R12_reg_32 (.CK( clk ) , .D( u2_N415 ) , .Q( u2_R12_32 ) );
  DFF_X1 u2_R12_reg_4 (.CK( clk ) , .D( u2_N387 ) , .Q( u2_R12_4 ) );
  DFF_X1 u2_R12_reg_5 (.CK( clk ) , .D( u2_N388 ) , .Q( u2_R12_5 ) );
  DFF_X1 u2_R12_reg_6 (.CK( clk ) , .D( u2_N389 ) , .Q( u2_R12_6 ) );
  DFF_X1 u2_R12_reg_7 (.CK( clk ) , .D( u2_N390 ) , .Q( u2_R12_7 ) );
  DFF_X1 u2_R12_reg_8 (.CK( clk ) , .D( u2_N391 ) , .Q( u2_R12_8 ) );
  DFF_X1 u2_R12_reg_9 (.CK( clk ) , .D( u2_N392 ) , .Q( u2_R12_9 ) );
  DFF_X1 u2_R13_reg_1 (.CK( clk ) , .D( u2_N416 ) , .Q( u2_R13_1 ) );
  DFF_X1 u2_R13_reg_10 (.CK( clk ) , .D( u2_N425 ) , .Q( u2_R13_10 ) );
  DFF_X1 u2_R13_reg_11 (.CK( clk ) , .D( u2_N426 ) , .Q( u2_R13_11 ) );
  DFF_X1 u2_R13_reg_12 (.CK( clk ) , .D( u2_N427 ) , .Q( u2_R13_12 ) );
  DFF_X1 u2_R13_reg_13 (.CK( clk ) , .D( u2_N428 ) , .Q( u2_R13_13 ) );
  DFF_X1 u2_R13_reg_14 (.CK( clk ) , .D( u2_N429 ) , .Q( u2_R13_14 ) );
  DFF_X1 u2_R13_reg_15 (.CK( clk ) , .D( u2_N430 ) , .Q( u2_R13_15 ) );
  DFF_X1 u2_R13_reg_16 (.CK( clk ) , .D( u2_N431 ) , .Q( u2_R13_16 ) );
  DFF_X1 u2_R13_reg_17 (.CK( clk ) , .D( u2_N432 ) , .Q( u2_R13_17 ) );
  DFF_X1 u2_R13_reg_18 (.CK( clk ) , .D( u2_N433 ) , .Q( u2_R13_18 ) );
  DFF_X1 u2_R13_reg_19 (.CK( clk ) , .D( u2_N434 ) , .Q( u2_R13_19 ) );
  DFF_X1 u2_R13_reg_2 (.CK( clk ) , .D( u2_N417 ) , .Q( u2_R13_2 ) );
  DFF_X1 u2_R13_reg_20 (.CK( clk ) , .D( u2_N435 ) , .Q( u2_R13_20 ) );
  DFF_X1 u2_R13_reg_21 (.CK( clk ) , .D( u2_N436 ) , .Q( u2_R13_21 ) );
  DFF_X1 u2_R13_reg_22 (.CK( clk ) , .D( u2_N437 ) , .Q( u2_R13_22 ) );
  DFF_X1 u2_R13_reg_23 (.CK( clk ) , .D( u2_N438 ) , .Q( u2_R13_23 ) );
  DFF_X1 u2_R13_reg_24 (.CK( clk ) , .D( u2_N439 ) , .Q( u2_R13_24 ) );
  DFF_X1 u2_R13_reg_25 (.CK( clk ) , .D( u2_N440 ) , .Q( u2_R13_25 ) );
  DFF_X1 u2_R13_reg_26 (.CK( clk ) , .D( u2_N441 ) , .Q( u2_R13_26 ) );
  DFF_X1 u2_R13_reg_27 (.CK( clk ) , .D( u2_N442 ) , .Q( u2_R13_27 ) );
  DFF_X1 u2_R13_reg_28 (.CK( clk ) , .D( u2_N443 ) , .Q( u2_R13_28 ) );
  DFF_X1 u2_R13_reg_29 (.CK( clk ) , .D( u2_N444 ) , .Q( u2_R13_29 ) );
  DFF_X1 u2_R13_reg_3 (.CK( clk ) , .D( u2_N418 ) , .Q( u2_R13_3 ) );
  DFF_X1 u2_R13_reg_30 (.CK( clk ) , .D( u2_N445 ) , .Q( u2_R13_30 ) );
  DFF_X1 u2_R13_reg_31 (.CK( clk ) , .D( u2_N446 ) , .Q( u2_R13_31 ) );
  DFF_X1 u2_R13_reg_32 (.CK( clk ) , .D( u2_N447 ) , .Q( u2_R13_32 ) );
  DFF_X1 u2_R13_reg_4 (.CK( clk ) , .D( u2_N419 ) , .Q( u2_R13_4 ) );
  DFF_X1 u2_R13_reg_5 (.CK( clk ) , .D( u2_N420 ) , .Q( u2_R13_5 ) );
  DFF_X1 u2_R13_reg_6 (.CK( clk ) , .D( u2_N421 ) , .Q( u2_R13_6 ) );
  DFF_X1 u2_R13_reg_7 (.CK( clk ) , .D( u2_N422 ) , .Q( u2_R13_7 ) );
  DFF_X1 u2_R13_reg_8 (.CK( clk ) , .D( u2_N423 ) , .Q( u2_R13_8 ) );
  DFF_X1 u2_R13_reg_9 (.CK( clk ) , .D( u2_N424 ) , .Q( u2_R13_9 ) );
  DFF_X1 u2_R14_reg_1 (.CK( clk ) , .Q( u2_FP_33 ) , .D( u2_N448 ) );
  DFF_X1 u2_R14_reg_10 (.CK( clk ) , .Q( u2_FP_42 ) , .D( u2_N457 ) );
  DFF_X1 u2_R14_reg_11 (.CK( clk ) , .Q( u2_FP_43 ) , .D( u2_N458 ) );
  DFF_X1 u2_R14_reg_12 (.CK( clk ) , .Q( u2_FP_44 ) , .D( u2_N459 ) );
  DFF_X1 u2_R14_reg_13 (.CK( clk ) , .Q( u2_FP_45 ) , .D( u2_N460 ) );
  DFF_X1 u2_R14_reg_14 (.CK( clk ) , .Q( u2_FP_46 ) , .D( u2_N461 ) );
  DFF_X1 u2_R14_reg_15 (.CK( clk ) , .Q( u2_FP_47 ) , .D( u2_N462 ) );
  DFF_X1 u2_R14_reg_16 (.CK( clk ) , .Q( u2_FP_48 ) , .D( u2_N463 ) );
  DFF_X1 u2_R14_reg_17 (.CK( clk ) , .Q( u2_FP_49 ) , .D( u2_N464 ) );
  DFF_X1 u2_R14_reg_18 (.CK( clk ) , .Q( u2_FP_50 ) , .D( u2_N465 ) );
  DFF_X1 u2_R14_reg_19 (.CK( clk ) , .Q( u2_FP_51 ) , .D( u2_N466 ) );
  DFF_X1 u2_R14_reg_2 (.CK( clk ) , .Q( u2_FP_34 ) , .D( u2_N449 ) );
  DFF_X1 u2_R14_reg_20 (.CK( clk ) , .Q( u2_FP_52 ) , .D( u2_N467 ) );
  DFF_X1 u2_R14_reg_21 (.CK( clk ) , .Q( u2_FP_53 ) , .D( u2_N468 ) );
  DFF_X1 u2_R14_reg_22 (.CK( clk ) , .Q( u2_FP_54 ) , .D( u2_N469 ) );
  DFF_X1 u2_R14_reg_23 (.CK( clk ) , .Q( u2_FP_55 ) , .D( u2_N470 ) );
  DFF_X1 u2_R14_reg_24 (.CK( clk ) , .Q( u2_FP_56 ) , .D( u2_N471 ) );
  DFF_X1 u2_R14_reg_25 (.CK( clk ) , .Q( u2_FP_57 ) , .D( u2_N472 ) );
  DFF_X1 u2_R14_reg_26 (.CK( clk ) , .Q( u2_FP_58 ) , .D( u2_N473 ) );
  DFF_X1 u2_R14_reg_27 (.CK( clk ) , .Q( u2_FP_59 ) , .D( u2_N474 ) );
  DFF_X1 u2_R14_reg_28 (.CK( clk ) , .Q( u2_FP_60 ) , .D( u2_N475 ) );
  DFF_X1 u2_R14_reg_29 (.CK( clk ) , .Q( u2_FP_61 ) , .D( u2_N476 ) );
  DFF_X1 u2_R14_reg_3 (.CK( clk ) , .Q( u2_FP_35 ) , .D( u2_N450 ) );
  DFF_X1 u2_R14_reg_30 (.CK( clk ) , .Q( u2_FP_62 ) , .D( u2_N477 ) );
  DFF_X1 u2_R14_reg_31 (.CK( clk ) , .Q( u2_FP_63 ) , .D( u2_N478 ) );
  DFF_X1 u2_R14_reg_32 (.CK( clk ) , .Q( u2_FP_64 ) , .D( u2_N479 ) );
  DFF_X1 u2_R14_reg_4 (.CK( clk ) , .Q( u2_FP_36 ) , .D( u2_N451 ) );
  DFF_X1 u2_R14_reg_5 (.CK( clk ) , .Q( u2_FP_37 ) , .D( u2_N452 ) );
  DFF_X1 u2_R14_reg_6 (.CK( clk ) , .Q( u2_FP_38 ) , .D( u2_N453 ) );
  DFF_X1 u2_R14_reg_7 (.CK( clk ) , .Q( u2_FP_39 ) , .D( u2_N454 ) );
  DFF_X1 u2_R14_reg_8 (.CK( clk ) , .Q( u2_FP_40 ) , .D( u2_N455 ) );
  DFF_X1 u2_R14_reg_9 (.CK( clk ) , .Q( u2_FP_41 ) , .D( u2_N456 ) );
  DFF_X1 u2_R1_reg_1 (.CK( clk ) , .D( u2_N32 ) , .Q( u2_R1_1 ) );
  DFF_X1 u2_R1_reg_10 (.CK( clk ) , .D( u2_N41 ) , .Q( u2_R1_10 ) );
  DFF_X1 u2_R1_reg_11 (.CK( clk ) , .D( u2_N42 ) , .Q( u2_R1_11 ) );
  DFF_X1 u2_R1_reg_12 (.CK( clk ) , .D( u2_N43 ) , .Q( u2_R1_12 ) );
  DFF_X1 u2_R1_reg_13 (.CK( clk ) , .D( u2_N44 ) , .Q( u2_R1_13 ) );
  DFF_X1 u2_R1_reg_14 (.CK( clk ) , .D( u2_N45 ) , .Q( u2_R1_14 ) );
  DFF_X1 u2_R1_reg_15 (.CK( clk ) , .D( u2_N46 ) , .Q( u2_R1_15 ) );
  DFF_X1 u2_R1_reg_16 (.CK( clk ) , .D( u2_N47 ) , .Q( u2_R1_16 ) );
  DFF_X1 u2_R1_reg_17 (.CK( clk ) , .D( u2_N48 ) , .Q( u2_R1_17 ) );
  DFF_X1 u2_R1_reg_18 (.CK( clk ) , .D( u2_N49 ) , .Q( u2_R1_18 ) );
  DFF_X1 u2_R1_reg_19 (.CK( clk ) , .D( u2_N50 ) , .Q( u2_R1_19 ) );
  DFF_X1 u2_R1_reg_2 (.CK( clk ) , .D( u2_N33 ) , .Q( u2_R1_2 ) );
  DFF_X1 u2_R1_reg_20 (.CK( clk ) , .D( u2_N51 ) , .Q( u2_R1_20 ) );
  DFF_X1 u2_R1_reg_21 (.CK( clk ) , .D( u2_N52 ) , .Q( u2_R1_21 ) );
  DFF_X1 u2_R1_reg_22 (.CK( clk ) , .D( u2_N53 ) , .Q( u2_R1_22 ) );
  DFF_X1 u2_R1_reg_23 (.CK( clk ) , .D( u2_N54 ) , .Q( u2_R1_23 ) );
  DFF_X1 u2_R1_reg_24 (.CK( clk ) , .D( u2_N55 ) , .Q( u2_R1_24 ) );
  DFF_X1 u2_R1_reg_25 (.CK( clk ) , .D( u2_N56 ) , .Q( u2_R1_25 ) );
  DFF_X1 u2_R1_reg_26 (.CK( clk ) , .D( u2_N57 ) , .Q( u2_R1_26 ) );
  DFF_X1 u2_R1_reg_27 (.CK( clk ) , .D( u2_N58 ) , .Q( u2_R1_27 ) );
  DFF_X1 u2_R1_reg_28 (.CK( clk ) , .D( u2_N59 ) , .Q( u2_R1_28 ) );
  DFF_X1 u2_R1_reg_29 (.CK( clk ) , .D( u2_N60 ) , .Q( u2_R1_29 ) );
  DFF_X1 u2_R1_reg_3 (.CK( clk ) , .D( u2_N34 ) , .Q( u2_R1_3 ) );
  DFF_X1 u2_R1_reg_30 (.CK( clk ) , .D( u2_N61 ) , .Q( u2_R1_30 ) );
  DFF_X1 u2_R1_reg_31 (.CK( clk ) , .D( u2_N62 ) , .Q( u2_R1_31 ) );
  DFF_X1 u2_R1_reg_32 (.CK( clk ) , .D( u2_N63 ) , .Q( u2_R1_32 ) );
  DFF_X1 u2_R1_reg_4 (.CK( clk ) , .D( u2_N35 ) , .Q( u2_R1_4 ) );
  DFF_X1 u2_R1_reg_5 (.CK( clk ) , .D( u2_N36 ) , .Q( u2_R1_5 ) );
  DFF_X1 u2_R1_reg_6 (.CK( clk ) , .D( u2_N37 ) , .Q( u2_R1_6 ) );
  DFF_X1 u2_R1_reg_7 (.CK( clk ) , .D( u2_N38 ) , .Q( u2_R1_7 ) );
  DFF_X1 u2_R1_reg_8 (.CK( clk ) , .D( u2_N39 ) , .Q( u2_R1_8 ) );
  DFF_X1 u2_R1_reg_9 (.CK( clk ) , .D( u2_N40 ) , .Q( u2_R1_9 ) );
  DFF_X1 u2_R2_reg_1 (.CK( clk ) , .D( u2_N64 ) , .Q( u2_R2_1 ) );
  DFF_X1 u2_R2_reg_10 (.CK( clk ) , .D( u2_N73 ) , .Q( u2_R2_10 ) );
  DFF_X1 u2_R2_reg_11 (.CK( clk ) , .D( u2_N74 ) , .Q( u2_R2_11 ) );
  DFF_X1 u2_R2_reg_12 (.CK( clk ) , .D( u2_N75 ) , .Q( u2_R2_12 ) );
  DFF_X1 u2_R2_reg_13 (.CK( clk ) , .D( u2_N76 ) , .Q( u2_R2_13 ) );
  DFF_X1 u2_R2_reg_14 (.CK( clk ) , .D( u2_N77 ) , .Q( u2_R2_14 ) );
  DFF_X1 u2_R2_reg_15 (.CK( clk ) , .D( u2_N78 ) , .Q( u2_R2_15 ) );
  DFF_X1 u2_R2_reg_16 (.CK( clk ) , .D( u2_N79 ) , .Q( u2_R2_16 ) );
  DFF_X1 u2_R2_reg_17 (.CK( clk ) , .D( u2_N80 ) , .Q( u2_R2_17 ) );
  DFF_X1 u2_R2_reg_18 (.CK( clk ) , .D( u2_N81 ) , .Q( u2_R2_18 ) );
  DFF_X1 u2_R2_reg_19 (.CK( clk ) , .D( u2_N82 ) , .Q( u2_R2_19 ) );
  DFF_X1 u2_R2_reg_2 (.CK( clk ) , .D( u2_N65 ) , .Q( u2_R2_2 ) );
  DFF_X1 u2_R2_reg_20 (.CK( clk ) , .D( u2_N83 ) , .Q( u2_R2_20 ) );
  DFF_X1 u2_R2_reg_21 (.CK( clk ) , .D( u2_N84 ) , .Q( u2_R2_21 ) );
  DFF_X1 u2_R2_reg_22 (.CK( clk ) , .D( u2_N85 ) , .Q( u2_R2_22 ) );
  DFF_X1 u2_R2_reg_23 (.CK( clk ) , .D( u2_N86 ) , .Q( u2_R2_23 ) );
  DFF_X1 u2_R2_reg_24 (.CK( clk ) , .D( u2_N87 ) , .Q( u2_R2_24 ) );
  DFF_X1 u2_R2_reg_25 (.CK( clk ) , .D( u2_N88 ) , .Q( u2_R2_25 ) );
  DFF_X1 u2_R2_reg_26 (.CK( clk ) , .D( u2_N89 ) , .Q( u2_R2_26 ) );
  DFF_X1 u2_R2_reg_27 (.CK( clk ) , .D( u2_N90 ) , .Q( u2_R2_27 ) );
  DFF_X1 u2_R2_reg_28 (.CK( clk ) , .D( u2_N91 ) , .Q( u2_R2_28 ) );
  DFF_X1 u2_R2_reg_29 (.CK( clk ) , .D( u2_N92 ) , .Q( u2_R2_29 ) );
  DFF_X1 u2_R2_reg_3 (.CK( clk ) , .D( u2_N66 ) , .Q( u2_R2_3 ) );
  DFF_X1 u2_R2_reg_30 (.CK( clk ) , .D( u2_N93 ) , .Q( u2_R2_30 ) );
  DFF_X1 u2_R2_reg_31 (.CK( clk ) , .D( u2_N94 ) , .Q( u2_R2_31 ) );
  DFF_X1 u2_R2_reg_32 (.CK( clk ) , .D( u2_N95 ) , .Q( u2_R2_32 ) );
  DFF_X1 u2_R2_reg_4 (.CK( clk ) , .D( u2_N67 ) , .Q( u2_R2_4 ) );
  DFF_X1 u2_R2_reg_5 (.CK( clk ) , .D( u2_N68 ) , .Q( u2_R2_5 ) );
  DFF_X1 u2_R2_reg_6 (.CK( clk ) , .D( u2_N69 ) , .Q( u2_R2_6 ) );
  DFF_X1 u2_R2_reg_7 (.CK( clk ) , .D( u2_N70 ) , .Q( u2_R2_7 ) );
  DFF_X1 u2_R2_reg_8 (.CK( clk ) , .D( u2_N71 ) , .Q( u2_R2_8 ) );
  DFF_X1 u2_R2_reg_9 (.CK( clk ) , .D( u2_N72 ) , .Q( u2_R2_9 ) );
  DFF_X1 u2_R3_reg_1 (.CK( clk ) , .D( u2_N96 ) , .Q( u2_R3_1 ) );
  DFF_X1 u2_R3_reg_10 (.CK( clk ) , .D( u2_N105 ) , .Q( u2_R3_10 ) );
  DFF_X1 u2_R3_reg_11 (.CK( clk ) , .D( u2_N106 ) , .Q( u2_R3_11 ) );
  DFF_X1 u2_R3_reg_12 (.CK( clk ) , .D( u2_N107 ) , .Q( u2_R3_12 ) );
  DFF_X1 u2_R3_reg_13 (.CK( clk ) , .D( u2_N108 ) , .Q( u2_R3_13 ) );
  DFF_X1 u2_R3_reg_14 (.CK( clk ) , .D( u2_N109 ) , .Q( u2_R3_14 ) );
  DFF_X1 u2_R3_reg_15 (.CK( clk ) , .D( u2_N110 ) , .Q( u2_R3_15 ) );
  DFF_X1 u2_R3_reg_16 (.CK( clk ) , .D( u2_N111 ) , .Q( u2_R3_16 ) );
  DFF_X1 u2_R3_reg_17 (.CK( clk ) , .D( u2_N112 ) , .Q( u2_R3_17 ) );
  DFF_X1 u2_R3_reg_18 (.CK( clk ) , .D( u2_N113 ) , .Q( u2_R3_18 ) );
  DFF_X1 u2_R3_reg_19 (.CK( clk ) , .D( u2_N114 ) , .Q( u2_R3_19 ) );
  DFF_X1 u2_R3_reg_2 (.CK( clk ) , .D( u2_N97 ) , .Q( u2_R3_2 ) );
  DFF_X1 u2_R3_reg_20 (.CK( clk ) , .D( u2_N115 ) , .Q( u2_R3_20 ) );
  DFF_X1 u2_R3_reg_21 (.CK( clk ) , .D( u2_N116 ) , .Q( u2_R3_21 ) );
  DFF_X1 u2_R3_reg_22 (.CK( clk ) , .D( u2_N117 ) , .Q( u2_R3_22 ) );
  DFF_X1 u2_R3_reg_23 (.CK( clk ) , .D( u2_N118 ) , .Q( u2_R3_23 ) );
  DFF_X1 u2_R3_reg_24 (.CK( clk ) , .D( u2_N119 ) , .Q( u2_R3_24 ) );
  DFF_X1 u2_R3_reg_25 (.CK( clk ) , .D( u2_N120 ) , .Q( u2_R3_25 ) );
  DFF_X1 u2_R3_reg_26 (.CK( clk ) , .D( u2_N121 ) , .Q( u2_R3_26 ) );
  DFF_X1 u2_R3_reg_27 (.CK( clk ) , .D( u2_N122 ) , .Q( u2_R3_27 ) );
  DFF_X1 u2_R3_reg_28 (.CK( clk ) , .D( u2_N123 ) , .Q( u2_R3_28 ) );
  DFF_X1 u2_R3_reg_29 (.CK( clk ) , .D( u2_N124 ) , .Q( u2_R3_29 ) );
  DFF_X1 u2_R3_reg_3 (.CK( clk ) , .D( u2_N98 ) , .Q( u2_R3_3 ) );
  DFF_X1 u2_R3_reg_30 (.CK( clk ) , .D( u2_N125 ) , .Q( u2_R3_30 ) );
  DFF_X1 u2_R3_reg_31 (.CK( clk ) , .D( u2_N126 ) , .Q( u2_R3_31 ) );
  DFF_X1 u2_R3_reg_32 (.CK( clk ) , .D( u2_N127 ) , .Q( u2_R3_32 ) );
  DFF_X1 u2_R3_reg_4 (.CK( clk ) , .D( u2_N99 ) , .Q( u2_R3_4 ) );
  DFF_X1 u2_R3_reg_5 (.CK( clk ) , .D( u2_N100 ) , .Q( u2_R3_5 ) );
  DFF_X1 u2_R3_reg_6 (.CK( clk ) , .D( u2_N101 ) , .Q( u2_R3_6 ) );
  DFF_X1 u2_R3_reg_7 (.CK( clk ) , .D( u2_N102 ) , .Q( u2_R3_7 ) );
  DFF_X1 u2_R3_reg_8 (.CK( clk ) , .D( u2_N103 ) , .Q( u2_R3_8 ) );
  DFF_X1 u2_R3_reg_9 (.CK( clk ) , .D( u2_N104 ) , .Q( u2_R3_9 ) );
  DFF_X1 u2_R4_reg_1 (.CK( clk ) , .D( u2_N128 ) , .Q( u2_R4_1 ) );
  DFF_X1 u2_R4_reg_10 (.CK( clk ) , .D( u2_N137 ) , .Q( u2_R4_10 ) );
  DFF_X1 u2_R4_reg_11 (.CK( clk ) , .D( u2_N138 ) , .Q( u2_R4_11 ) );
  DFF_X1 u2_R4_reg_12 (.CK( clk ) , .D( u2_N139 ) , .Q( u2_R4_12 ) );
  DFF_X1 u2_R4_reg_13 (.CK( clk ) , .D( u2_N140 ) , .Q( u2_R4_13 ) );
  DFF_X1 u2_R4_reg_14 (.CK( clk ) , .D( u2_N141 ) , .Q( u2_R4_14 ) );
  DFF_X1 u2_R4_reg_15 (.CK( clk ) , .D( u2_N142 ) , .Q( u2_R4_15 ) );
  DFF_X1 u2_R4_reg_16 (.CK( clk ) , .D( u2_N143 ) , .Q( u2_R4_16 ) );
  DFF_X1 u2_R4_reg_17 (.CK( clk ) , .D( u2_N144 ) , .Q( u2_R4_17 ) );
  DFF_X1 u2_R4_reg_18 (.CK( clk ) , .D( u2_N145 ) , .Q( u2_R4_18 ) );
  DFF_X1 u2_R4_reg_19 (.CK( clk ) , .D( u2_N146 ) , .Q( u2_R4_19 ) );
  DFF_X1 u2_R4_reg_2 (.CK( clk ) , .D( u2_N129 ) , .Q( u2_R4_2 ) );
  DFF_X1 u2_R4_reg_20 (.CK( clk ) , .D( u2_N147 ) , .Q( u2_R4_20 ) );
  DFF_X1 u2_R4_reg_21 (.CK( clk ) , .D( u2_N148 ) , .Q( u2_R4_21 ) );
  DFF_X1 u2_R4_reg_22 (.CK( clk ) , .D( u2_N149 ) , .Q( u2_R4_22 ) );
  DFF_X1 u2_R4_reg_23 (.CK( clk ) , .D( u2_N150 ) , .Q( u2_R4_23 ) );
  DFF_X1 u2_R4_reg_24 (.CK( clk ) , .D( u2_N151 ) , .Q( u2_R4_24 ) );
  DFF_X1 u2_R4_reg_25 (.CK( clk ) , .D( u2_N152 ) , .Q( u2_R4_25 ) );
  DFF_X1 u2_R4_reg_26 (.CK( clk ) , .D( u2_N153 ) , .Q( u2_R4_26 ) );
  DFF_X1 u2_R4_reg_27 (.CK( clk ) , .D( u2_N154 ) , .Q( u2_R4_27 ) );
  DFF_X1 u2_R4_reg_28 (.CK( clk ) , .D( u2_N155 ) , .Q( u2_R4_28 ) );
  DFF_X1 u2_R4_reg_29 (.CK( clk ) , .D( u2_N156 ) , .Q( u2_R4_29 ) );
  DFF_X1 u2_R4_reg_3 (.CK( clk ) , .D( u2_N130 ) , .Q( u2_R4_3 ) );
  DFF_X1 u2_R4_reg_30 (.CK( clk ) , .D( u2_N157 ) , .Q( u2_R4_30 ) );
  DFF_X1 u2_R4_reg_31 (.CK( clk ) , .D( u2_N158 ) , .Q( u2_R4_31 ) );
  DFF_X1 u2_R4_reg_32 (.CK( clk ) , .D( u2_N159 ) , .Q( u2_R4_32 ) );
  DFF_X1 u2_R4_reg_4 (.CK( clk ) , .D( u2_N131 ) , .Q( u2_R4_4 ) );
  DFF_X1 u2_R4_reg_5 (.CK( clk ) , .D( u2_N132 ) , .Q( u2_R4_5 ) );
  DFF_X1 u2_R4_reg_6 (.CK( clk ) , .D( u2_N133 ) , .Q( u2_R4_6 ) );
  DFF_X1 u2_R4_reg_7 (.CK( clk ) , .D( u2_N134 ) , .Q( u2_R4_7 ) );
  DFF_X1 u2_R4_reg_8 (.CK( clk ) , .D( u2_N135 ) , .Q( u2_R4_8 ) );
  DFF_X1 u2_R4_reg_9 (.CK( clk ) , .D( u2_N136 ) , .Q( u2_R4_9 ) );
  DFF_X1 u2_R5_reg_1 (.CK( clk ) , .D( u2_N160 ) , .Q( u2_R5_1 ) );
  DFF_X1 u2_R5_reg_10 (.CK( clk ) , .D( u2_N169 ) , .Q( u2_R5_10 ) );
  DFF_X1 u2_R5_reg_11 (.CK( clk ) , .D( u2_N170 ) , .Q( u2_R5_11 ) );
  DFF_X1 u2_R5_reg_12 (.CK( clk ) , .D( u2_N171 ) , .Q( u2_R5_12 ) );
  DFF_X1 u2_R5_reg_13 (.CK( clk ) , .D( u2_N172 ) , .Q( u2_R5_13 ) );
  DFF_X1 u2_R5_reg_14 (.CK( clk ) , .D( u2_N173 ) , .Q( u2_R5_14 ) );
  DFF_X1 u2_R5_reg_15 (.CK( clk ) , .D( u2_N174 ) , .Q( u2_R5_15 ) );
  DFF_X1 u2_R5_reg_16 (.CK( clk ) , .D( u2_N175 ) , .Q( u2_R5_16 ) );
  DFF_X1 u2_R5_reg_17 (.CK( clk ) , .D( u2_N176 ) , .Q( u2_R5_17 ) );
  DFF_X1 u2_R5_reg_18 (.CK( clk ) , .D( u2_N177 ) , .Q( u2_R5_18 ) );
  DFF_X1 u2_R5_reg_19 (.CK( clk ) , .D( u2_N178 ) , .Q( u2_R5_19 ) );
  DFF_X1 u2_R5_reg_2 (.CK( clk ) , .D( u2_N161 ) , .Q( u2_R5_2 ) );
  DFF_X1 u2_R5_reg_20 (.CK( clk ) , .D( u2_N179 ) , .Q( u2_R5_20 ) );
  DFF_X1 u2_R5_reg_21 (.CK( clk ) , .D( u2_N180 ) , .Q( u2_R5_21 ) );
  DFF_X1 u2_R5_reg_22 (.CK( clk ) , .D( u2_N181 ) , .Q( u2_R5_22 ) );
  DFF_X1 u2_R5_reg_23 (.CK( clk ) , .D( u2_N182 ) , .Q( u2_R5_23 ) );
  DFF_X1 u2_R5_reg_24 (.CK( clk ) , .D( u2_N183 ) , .Q( u2_R5_24 ) );
  DFF_X1 u2_R5_reg_25 (.CK( clk ) , .D( u2_N184 ) , .Q( u2_R5_25 ) );
  DFF_X1 u2_R5_reg_26 (.CK( clk ) , .D( u2_N185 ) , .Q( u2_R5_26 ) );
  DFF_X1 u2_R5_reg_27 (.CK( clk ) , .D( u2_N186 ) , .Q( u2_R5_27 ) );
  DFF_X1 u2_R5_reg_28 (.CK( clk ) , .D( u2_N187 ) , .Q( u2_R5_28 ) );
  DFF_X1 u2_R5_reg_29 (.CK( clk ) , .D( u2_N188 ) , .Q( u2_R5_29 ) );
  DFF_X1 u2_R5_reg_3 (.CK( clk ) , .D( u2_N162 ) , .Q( u2_R5_3 ) );
  DFF_X1 u2_R5_reg_30 (.CK( clk ) , .D( u2_N189 ) , .Q( u2_R5_30 ) );
  DFF_X1 u2_R5_reg_31 (.CK( clk ) , .D( u2_N190 ) , .Q( u2_R5_31 ) );
  DFF_X1 u2_R5_reg_32 (.CK( clk ) , .D( u2_N191 ) , .Q( u2_R5_32 ) );
  DFF_X1 u2_R5_reg_4 (.CK( clk ) , .D( u2_N163 ) , .Q( u2_R5_4 ) );
  DFF_X1 u2_R5_reg_5 (.CK( clk ) , .D( u2_N164 ) , .Q( u2_R5_5 ) );
  DFF_X1 u2_R5_reg_6 (.CK( clk ) , .D( u2_N165 ) , .Q( u2_R5_6 ) );
  DFF_X1 u2_R5_reg_7 (.CK( clk ) , .D( u2_N166 ) , .Q( u2_R5_7 ) );
  DFF_X1 u2_R5_reg_8 (.CK( clk ) , .D( u2_N167 ) , .Q( u2_R5_8 ) );
  DFF_X1 u2_R5_reg_9 (.CK( clk ) , .D( u2_N168 ) , .Q( u2_R5_9 ) );
  DFF_X1 u2_R6_reg_1 (.CK( clk ) , .D( u2_N192 ) , .Q( u2_R6_1 ) );
  DFF_X1 u2_R6_reg_10 (.CK( clk ) , .D( u2_N201 ) , .Q( u2_R6_10 ) );
  DFF_X1 u2_R6_reg_11 (.CK( clk ) , .D( u2_N202 ) , .Q( u2_R6_11 ) );
  DFF_X1 u2_R6_reg_12 (.CK( clk ) , .D( u2_N203 ) , .Q( u2_R6_12 ) );
  DFF_X1 u2_R6_reg_13 (.CK( clk ) , .D( u2_N204 ) , .Q( u2_R6_13 ) );
  DFF_X1 u2_R6_reg_14 (.CK( clk ) , .D( u2_N205 ) , .Q( u2_R6_14 ) );
  DFF_X1 u2_R6_reg_15 (.CK( clk ) , .D( u2_N206 ) , .Q( u2_R6_15 ) );
  DFF_X1 u2_R6_reg_16 (.CK( clk ) , .D( u2_N207 ) , .Q( u2_R6_16 ) );
  DFF_X1 u2_R6_reg_17 (.CK( clk ) , .D( u2_N208 ) , .Q( u2_R6_17 ) );
  DFF_X1 u2_R6_reg_18 (.CK( clk ) , .D( u2_N209 ) , .Q( u2_R6_18 ) );
  DFF_X1 u2_R6_reg_19 (.CK( clk ) , .D( u2_N210 ) , .Q( u2_R6_19 ) );
  DFF_X1 u2_R6_reg_2 (.CK( clk ) , .D( u2_N193 ) , .Q( u2_R6_2 ) );
  DFF_X1 u2_R6_reg_20 (.CK( clk ) , .D( u2_N211 ) , .Q( u2_R6_20 ) );
  DFF_X1 u2_R6_reg_21 (.CK( clk ) , .D( u2_N212 ) , .Q( u2_R6_21 ) );
  DFF_X1 u2_R6_reg_22 (.CK( clk ) , .D( u2_N213 ) , .Q( u2_R6_22 ) );
  DFF_X1 u2_R6_reg_23 (.CK( clk ) , .D( u2_N214 ) , .Q( u2_R6_23 ) );
  DFF_X1 u2_R6_reg_24 (.CK( clk ) , .D( u2_N215 ) , .Q( u2_R6_24 ) );
  DFF_X1 u2_R6_reg_25 (.CK( clk ) , .D( u2_N216 ) , .Q( u2_R6_25 ) );
  DFF_X1 u2_R6_reg_26 (.CK( clk ) , .D( u2_N217 ) , .Q( u2_R6_26 ) );
  DFF_X1 u2_R6_reg_27 (.CK( clk ) , .D( u2_N218 ) , .Q( u2_R6_27 ) );
  DFF_X1 u2_R6_reg_28 (.CK( clk ) , .D( u2_N219 ) , .Q( u2_R6_28 ) );
  DFF_X1 u2_R6_reg_29 (.CK( clk ) , .D( u2_N220 ) , .Q( u2_R6_29 ) );
  DFF_X1 u2_R6_reg_3 (.CK( clk ) , .D( u2_N194 ) , .Q( u2_R6_3 ) );
  DFF_X1 u2_R6_reg_30 (.CK( clk ) , .D( u2_N221 ) , .Q( u2_R6_30 ) );
  DFF_X1 u2_R6_reg_31 (.CK( clk ) , .D( u2_N222 ) , .Q( u2_R6_31 ) );
  DFF_X1 u2_R6_reg_32 (.CK( clk ) , .D( u2_N223 ) , .Q( u2_R6_32 ) );
  DFF_X1 u2_R6_reg_4 (.CK( clk ) , .D( u2_N195 ) , .Q( u2_R6_4 ) );
  DFF_X1 u2_R6_reg_5 (.CK( clk ) , .D( u2_N196 ) , .Q( u2_R6_5 ) );
  DFF_X1 u2_R6_reg_6 (.CK( clk ) , .D( u2_N197 ) , .Q( u2_R6_6 ) );
  DFF_X1 u2_R6_reg_7 (.CK( clk ) , .D( u2_N198 ) , .Q( u2_R6_7 ) );
  DFF_X1 u2_R6_reg_8 (.CK( clk ) , .D( u2_N199 ) , .Q( u2_R6_8 ) );
  DFF_X1 u2_R6_reg_9 (.CK( clk ) , .D( u2_N200 ) , .Q( u2_R6_9 ) );
  DFF_X1 u2_R7_reg_1 (.CK( clk ) , .D( u2_N224 ) , .Q( u2_R7_1 ) );
  DFF_X1 u2_R7_reg_10 (.CK( clk ) , .D( u2_N233 ) , .Q( u2_R7_10 ) );
  DFF_X1 u2_R7_reg_11 (.CK( clk ) , .D( u2_N234 ) , .Q( u2_R7_11 ) );
  DFF_X1 u2_R7_reg_12 (.CK( clk ) , .D( u2_N235 ) , .Q( u2_R7_12 ) );
  DFF_X1 u2_R7_reg_13 (.CK( clk ) , .D( u2_N236 ) , .Q( u2_R7_13 ) );
  DFF_X1 u2_R7_reg_14 (.CK( clk ) , .D( u2_N237 ) , .Q( u2_R7_14 ) );
  DFF_X1 u2_R7_reg_15 (.CK( clk ) , .D( u2_N238 ) , .Q( u2_R7_15 ) );
  DFF_X1 u2_R7_reg_16 (.CK( clk ) , .D( u2_N239 ) , .Q( u2_R7_16 ) );
  DFF_X1 u2_R7_reg_17 (.CK( clk ) , .D( u2_N240 ) , .Q( u2_R7_17 ) );
  DFF_X1 u2_R7_reg_18 (.CK( clk ) , .D( u2_N241 ) , .Q( u2_R7_18 ) );
  DFF_X1 u2_R7_reg_19 (.CK( clk ) , .D( u2_N242 ) , .Q( u2_R7_19 ) );
  DFF_X1 u2_R7_reg_2 (.CK( clk ) , .D( u2_N225 ) , .Q( u2_R7_2 ) );
  DFF_X1 u2_R7_reg_20 (.CK( clk ) , .D( u2_N243 ) , .Q( u2_R7_20 ) );
  DFF_X1 u2_R7_reg_21 (.CK( clk ) , .D( u2_N244 ) , .Q( u2_R7_21 ) );
  DFF_X1 u2_R7_reg_22 (.CK( clk ) , .D( u2_N245 ) , .Q( u2_R7_22 ) );
  DFF_X1 u2_R7_reg_23 (.CK( clk ) , .D( u2_N246 ) , .Q( u2_R7_23 ) );
  DFF_X1 u2_R7_reg_24 (.CK( clk ) , .D( u2_N247 ) , .Q( u2_R7_24 ) );
  DFF_X1 u2_R7_reg_25 (.CK( clk ) , .D( u2_N248 ) , .Q( u2_R7_25 ) );
  DFF_X1 u2_R7_reg_26 (.CK( clk ) , .D( u2_N249 ) , .Q( u2_R7_26 ) );
  DFF_X1 u2_R7_reg_27 (.CK( clk ) , .D( u2_N250 ) , .Q( u2_R7_27 ) );
  DFF_X1 u2_R7_reg_28 (.CK( clk ) , .D( u2_N251 ) , .Q( u2_R7_28 ) );
  DFF_X1 u2_R7_reg_29 (.CK( clk ) , .D( u2_N252 ) , .Q( u2_R7_29 ) );
  DFF_X1 u2_R7_reg_3 (.CK( clk ) , .D( u2_N226 ) , .Q( u2_R7_3 ) );
  DFF_X1 u2_R7_reg_30 (.CK( clk ) , .D( u2_N253 ) , .Q( u2_R7_30 ) );
  DFF_X1 u2_R7_reg_31 (.CK( clk ) , .D( u2_N254 ) , .Q( u2_R7_31 ) );
  DFF_X1 u2_R7_reg_32 (.CK( clk ) , .D( u2_N255 ) , .Q( u2_R7_32 ) );
  DFF_X1 u2_R7_reg_4 (.CK( clk ) , .D( u2_N227 ) , .Q( u2_R7_4 ) );
  DFF_X1 u2_R7_reg_5 (.CK( clk ) , .D( u2_N228 ) , .Q( u2_R7_5 ) );
  DFF_X1 u2_R7_reg_6 (.CK( clk ) , .D( u2_N229 ) , .Q( u2_R7_6 ) );
  DFF_X1 u2_R7_reg_7 (.CK( clk ) , .D( u2_N230 ) , .Q( u2_R7_7 ) );
  DFF_X1 u2_R7_reg_8 (.CK( clk ) , .D( u2_N231 ) , .Q( u2_R7_8 ) );
  DFF_X1 u2_R7_reg_9 (.CK( clk ) , .D( u2_N232 ) , .Q( u2_R7_9 ) );
  DFF_X1 u2_R8_reg_1 (.CK( clk ) , .D( u2_N256 ) , .Q( u2_R8_1 ) );
  DFF_X1 u2_R8_reg_10 (.CK( clk ) , .D( u2_N265 ) , .Q( u2_R8_10 ) );
  DFF_X1 u2_R8_reg_11 (.CK( clk ) , .D( u2_N266 ) , .Q( u2_R8_11 ) );
  DFF_X1 u2_R8_reg_12 (.CK( clk ) , .D( u2_N267 ) , .Q( u2_R8_12 ) );
  DFF_X1 u2_R8_reg_13 (.CK( clk ) , .D( u2_N268 ) , .Q( u2_R8_13 ) );
  DFF_X1 u2_R8_reg_14 (.CK( clk ) , .D( u2_N269 ) , .Q( u2_R8_14 ) );
  DFF_X1 u2_R8_reg_15 (.CK( clk ) , .D( u2_N270 ) , .Q( u2_R8_15 ) );
  DFF_X1 u2_R8_reg_16 (.CK( clk ) , .D( u2_N271 ) , .Q( u2_R8_16 ) );
  DFF_X1 u2_R8_reg_17 (.CK( clk ) , .D( u2_N272 ) , .Q( u2_R8_17 ) );
  DFF_X1 u2_R8_reg_18 (.CK( clk ) , .D( u2_N273 ) , .Q( u2_R8_18 ) );
  DFF_X1 u2_R8_reg_19 (.CK( clk ) , .D( u2_N274 ) , .Q( u2_R8_19 ) );
  DFF_X1 u2_R8_reg_2 (.CK( clk ) , .D( u2_N257 ) , .Q( u2_R8_2 ) );
  DFF_X1 u2_R8_reg_20 (.CK( clk ) , .D( u2_N275 ) , .Q( u2_R8_20 ) );
  DFF_X1 u2_R8_reg_21 (.CK( clk ) , .D( u2_N276 ) , .Q( u2_R8_21 ) );
  DFF_X1 u2_R8_reg_22 (.CK( clk ) , .D( u2_N277 ) , .Q( u2_R8_22 ) );
  DFF_X1 u2_R8_reg_23 (.CK( clk ) , .D( u2_N278 ) , .Q( u2_R8_23 ) );
  DFF_X1 u2_R8_reg_24 (.CK( clk ) , .D( u2_N279 ) , .Q( u2_R8_24 ) );
  DFF_X1 u2_R8_reg_25 (.CK( clk ) , .D( u2_N280 ) , .Q( u2_R8_25 ) );
  DFF_X1 u2_R8_reg_26 (.CK( clk ) , .D( u2_N281 ) , .Q( u2_R8_26 ) );
  DFF_X1 u2_R8_reg_27 (.CK( clk ) , .D( u2_N282 ) , .Q( u2_R8_27 ) );
  DFF_X1 u2_R8_reg_28 (.CK( clk ) , .D( u2_N283 ) , .Q( u2_R8_28 ) );
  DFF_X1 u2_R8_reg_29 (.CK( clk ) , .D( u2_N284 ) , .Q( u2_R8_29 ) );
  DFF_X1 u2_R8_reg_3 (.CK( clk ) , .D( u2_N258 ) , .Q( u2_R8_3 ) );
  DFF_X1 u2_R8_reg_30 (.CK( clk ) , .D( u2_N285 ) , .Q( u2_R8_30 ) );
  DFF_X1 u2_R8_reg_31 (.CK( clk ) , .D( u2_N286 ) , .Q( u2_R8_31 ) );
  DFF_X1 u2_R8_reg_32 (.CK( clk ) , .D( u2_N287 ) , .Q( u2_R8_32 ) );
  DFF_X1 u2_R8_reg_4 (.CK( clk ) , .D( u2_N259 ) , .Q( u2_R8_4 ) );
  DFF_X1 u2_R8_reg_5 (.CK( clk ) , .D( u2_N260 ) , .Q( u2_R8_5 ) );
  DFF_X1 u2_R8_reg_6 (.CK( clk ) , .D( u2_N261 ) , .Q( u2_R8_6 ) );
  DFF_X1 u2_R8_reg_7 (.CK( clk ) , .D( u2_N262 ) , .Q( u2_R8_7 ) );
  DFF_X1 u2_R8_reg_8 (.CK( clk ) , .D( u2_N263 ) , .Q( u2_R8_8 ) );
  DFF_X1 u2_R8_reg_9 (.CK( clk ) , .D( u2_N264 ) , .Q( u2_R8_9 ) );
  DFF_X1 u2_R9_reg_1 (.CK( clk ) , .D( u2_N288 ) , .Q( u2_R9_1 ) );
  DFF_X1 u2_R9_reg_10 (.CK( clk ) , .D( u2_N297 ) , .Q( u2_R9_10 ) );
  DFF_X1 u2_R9_reg_11 (.CK( clk ) , .D( u2_N298 ) , .Q( u2_R9_11 ) );
  DFF_X1 u2_R9_reg_12 (.CK( clk ) , .D( u2_N299 ) , .Q( u2_R9_12 ) );
  DFF_X1 u2_R9_reg_13 (.CK( clk ) , .D( u2_N300 ) , .Q( u2_R9_13 ) );
  DFF_X1 u2_R9_reg_14 (.CK( clk ) , .D( u2_N301 ) , .Q( u2_R9_14 ) );
  DFF_X1 u2_R9_reg_15 (.CK( clk ) , .D( u2_N302 ) , .Q( u2_R9_15 ) );
  DFF_X1 u2_R9_reg_16 (.CK( clk ) , .D( u2_N303 ) , .Q( u2_R9_16 ) );
  DFF_X1 u2_R9_reg_17 (.CK( clk ) , .D( u2_N304 ) , .Q( u2_R9_17 ) );
  DFF_X1 u2_R9_reg_18 (.CK( clk ) , .D( u2_N305 ) , .Q( u2_R9_18 ) );
  DFF_X1 u2_R9_reg_19 (.CK( clk ) , .D( u2_N306 ) , .Q( u2_R9_19 ) );
  DFF_X1 u2_R9_reg_2 (.CK( clk ) , .D( u2_N289 ) , .Q( u2_R9_2 ) );
  DFF_X1 u2_R9_reg_20 (.CK( clk ) , .D( u2_N307 ) , .Q( u2_R9_20 ) );
  DFF_X1 u2_R9_reg_21 (.CK( clk ) , .D( u2_N308 ) , .Q( u2_R9_21 ) );
  DFF_X1 u2_R9_reg_22 (.CK( clk ) , .D( u2_N309 ) , .Q( u2_R9_22 ) );
  DFF_X1 u2_R9_reg_23 (.CK( clk ) , .D( u2_N310 ) , .Q( u2_R9_23 ) );
  DFF_X1 u2_R9_reg_24 (.CK( clk ) , .D( u2_N311 ) , .Q( u2_R9_24 ) );
  DFF_X1 u2_R9_reg_25 (.CK( clk ) , .D( u2_N312 ) , .Q( u2_R9_25 ) );
  DFF_X1 u2_R9_reg_26 (.CK( clk ) , .D( u2_N313 ) , .Q( u2_R9_26 ) );
  DFF_X1 u2_R9_reg_27 (.CK( clk ) , .D( u2_N314 ) , .Q( u2_R9_27 ) );
  DFF_X1 u2_R9_reg_28 (.CK( clk ) , .D( u2_N315 ) , .Q( u2_R9_28 ) );
  DFF_X1 u2_R9_reg_29 (.CK( clk ) , .D( u2_N316 ) , .Q( u2_R9_29 ) );
  DFF_X1 u2_R9_reg_3 (.CK( clk ) , .D( u2_N290 ) , .Q( u2_R9_3 ) );
  DFF_X1 u2_R9_reg_30 (.CK( clk ) , .D( u2_N317 ) , .Q( u2_R9_30 ) );
  DFF_X1 u2_R9_reg_31 (.CK( clk ) , .D( u2_N318 ) , .Q( u2_R9_31 ) );
  DFF_X1 u2_R9_reg_32 (.CK( clk ) , .D( u2_N319 ) , .Q( u2_R9_32 ) );
  DFF_X1 u2_R9_reg_4 (.CK( clk ) , .D( u2_N291 ) , .Q( u2_R9_4 ) );
  DFF_X1 u2_R9_reg_5 (.CK( clk ) , .D( u2_N292 ) , .Q( u2_R9_5 ) );
  DFF_X1 u2_R9_reg_6 (.CK( clk ) , .D( u2_N293 ) , .Q( u2_R9_6 ) );
  DFF_X1 u2_R9_reg_7 (.CK( clk ) , .D( u2_N294 ) , .Q( u2_R9_7 ) );
  DFF_X1 u2_R9_reg_8 (.CK( clk ) , .D( u2_N295 ) , .Q( u2_R9_8 ) );
  DFF_X1 u2_R9_reg_9 (.CK( clk ) , .D( u2_N296 ) , .Q( u2_R9_9 ) );
  DFF_X1 u2_desIn_r_reg_0 (.CK( clk ) , .D( stage2_out_0 ) , .Q( u2_desIn_r_0 ) );
  DFF_X1 u2_desIn_r_reg_1 (.CK( clk ) , .D( stage2_out_1 ) , .Q( u2_desIn_r_1 ) );
  DFF_X1 u2_desIn_r_reg_10 (.CK( clk ) , .D( stage2_out_10 ) , .Q( u2_desIn_r_10 ) );
  DFF_X1 u2_desIn_r_reg_11 (.CK( clk ) , .D( stage2_out_11 ) , .Q( u2_desIn_r_11 ) );
  DFF_X1 u2_desIn_r_reg_12 (.CK( clk ) , .D( stage2_out_12 ) , .Q( u2_desIn_r_12 ) );
  DFF_X1 u2_desIn_r_reg_13 (.CK( clk ) , .D( stage2_out_13 ) , .Q( u2_desIn_r_13 ) );
  DFF_X1 u2_desIn_r_reg_14 (.CK( clk ) , .D( stage2_out_14 ) , .Q( u2_desIn_r_14 ) );
  DFF_X1 u2_desIn_r_reg_15 (.CK( clk ) , .D( stage2_out_15 ) , .Q( u2_desIn_r_15 ) );
  DFF_X1 u2_desIn_r_reg_16 (.CK( clk ) , .D( stage2_out_16 ) , .Q( u2_desIn_r_16 ) );
  DFF_X1 u2_desIn_r_reg_17 (.CK( clk ) , .D( stage2_out_17 ) , .Q( u2_desIn_r_17 ) );
  DFF_X1 u2_desIn_r_reg_18 (.CK( clk ) , .D( stage2_out_18 ) , .Q( u2_desIn_r_18 ) );
  DFF_X1 u2_desIn_r_reg_19 (.CK( clk ) , .D( stage2_out_19 ) , .Q( u2_desIn_r_19 ) );
  DFF_X1 u2_desIn_r_reg_2 (.CK( clk ) , .D( stage2_out_2 ) , .Q( u2_desIn_r_2 ) );
  DFF_X1 u2_desIn_r_reg_20 (.CK( clk ) , .D( stage2_out_20 ) , .Q( u2_desIn_r_20 ) );
  DFF_X1 u2_desIn_r_reg_21 (.CK( clk ) , .D( stage2_out_21 ) , .Q( u2_desIn_r_21 ) );
  DFF_X1 u2_desIn_r_reg_22 (.CK( clk ) , .D( stage2_out_22 ) , .Q( u2_desIn_r_22 ) );
  DFF_X1 u2_desIn_r_reg_23 (.CK( clk ) , .D( stage2_out_23 ) , .Q( u2_desIn_r_23 ) );
  DFF_X1 u2_desIn_r_reg_24 (.CK( clk ) , .D( stage2_out_24 ) , .Q( u2_desIn_r_24 ) );
  DFF_X1 u2_desIn_r_reg_25 (.CK( clk ) , .D( stage2_out_25 ) , .Q( u2_desIn_r_25 ) );
  DFF_X1 u2_desIn_r_reg_26 (.CK( clk ) , .D( stage2_out_26 ) , .Q( u2_desIn_r_26 ) );
  DFF_X1 u2_desIn_r_reg_27 (.CK( clk ) , .D( stage2_out_27 ) , .Q( u2_desIn_r_27 ) );
  DFF_X1 u2_desIn_r_reg_28 (.CK( clk ) , .D( stage2_out_28 ) , .Q( u2_desIn_r_28 ) );
  DFF_X1 u2_desIn_r_reg_29 (.CK( clk ) , .D( stage2_out_29 ) , .Q( u2_desIn_r_29 ) );
  DFF_X1 u2_desIn_r_reg_3 (.CK( clk ) , .D( stage2_out_3 ) , .Q( u2_desIn_r_3 ) );
  DFF_X1 u2_desIn_r_reg_30 (.CK( clk ) , .D( stage2_out_30 ) , .Q( u2_desIn_r_30 ) );
  DFF_X1 u2_desIn_r_reg_31 (.CK( clk ) , .D( stage2_out_31 ) , .Q( u2_desIn_r_31 ) );
  DFF_X1 u2_desIn_r_reg_32 (.CK( clk ) , .D( stage2_out_32 ) , .Q( u2_desIn_r_32 ) );
  DFF_X1 u2_desIn_r_reg_33 (.CK( clk ) , .D( stage2_out_33 ) , .Q( u2_desIn_r_33 ) );
  DFF_X1 u2_desIn_r_reg_34 (.CK( clk ) , .D( stage2_out_34 ) , .Q( u2_desIn_r_34 ) );
  DFF_X1 u2_desIn_r_reg_35 (.CK( clk ) , .D( stage2_out_35 ) , .Q( u2_desIn_r_35 ) );
  DFF_X1 u2_desIn_r_reg_36 (.CK( clk ) , .D( stage2_out_36 ) , .Q( u2_desIn_r_36 ) );
  DFF_X1 u2_desIn_r_reg_37 (.CK( clk ) , .D( stage2_out_37 ) , .Q( u2_desIn_r_37 ) );
  DFF_X1 u2_desIn_r_reg_38 (.CK( clk ) , .D( stage2_out_38 ) , .Q( u2_desIn_r_38 ) );
  DFF_X1 u2_desIn_r_reg_39 (.CK( clk ) , .D( stage2_out_39 ) , .Q( u2_desIn_r_39 ) );
  DFF_X1 u2_desIn_r_reg_4 (.CK( clk ) , .D( stage2_out_4 ) , .Q( u2_desIn_r_4 ) );
  DFF_X1 u2_desIn_r_reg_40 (.CK( clk ) , .D( stage2_out_40 ) , .Q( u2_desIn_r_40 ) );
  DFF_X1 u2_desIn_r_reg_41 (.CK( clk ) , .D( stage2_out_41 ) , .Q( u2_desIn_r_41 ) );
  DFF_X1 u2_desIn_r_reg_42 (.CK( clk ) , .D( stage2_out_42 ) , .Q( u2_desIn_r_42 ) );
  DFF_X1 u2_desIn_r_reg_43 (.CK( clk ) , .D( stage2_out_43 ) , .Q( u2_desIn_r_43 ) );
  DFF_X1 u2_desIn_r_reg_44 (.CK( clk ) , .D( stage2_out_44 ) , .Q( u2_desIn_r_44 ) );
  DFF_X1 u2_desIn_r_reg_45 (.CK( clk ) , .D( stage2_out_45 ) , .Q( u2_desIn_r_45 ) );
  DFF_X1 u2_desIn_r_reg_46 (.CK( clk ) , .D( stage2_out_46 ) , .Q( u2_desIn_r_46 ) );
  DFF_X1 u2_desIn_r_reg_47 (.CK( clk ) , .D( stage2_out_47 ) , .Q( u2_desIn_r_47 ) );
  DFF_X1 u2_desIn_r_reg_48 (.CK( clk ) , .D( stage2_out_48 ) , .Q( u2_desIn_r_48 ) );
  DFF_X1 u2_desIn_r_reg_49 (.CK( clk ) , .D( stage2_out_49 ) , .Q( u2_desIn_r_49 ) );
  DFF_X1 u2_desIn_r_reg_5 (.CK( clk ) , .D( stage2_out_5 ) , .Q( u2_desIn_r_5 ) );
  DFF_X1 u2_desIn_r_reg_50 (.CK( clk ) , .D( stage2_out_50 ) , .Q( u2_desIn_r_50 ) );
  DFF_X1 u2_desIn_r_reg_51 (.CK( clk ) , .D( stage2_out_51 ) , .Q( u2_desIn_r_51 ) );
  DFF_X1 u2_desIn_r_reg_52 (.CK( clk ) , .D( stage2_out_52 ) , .Q( u2_desIn_r_52 ) );
  DFF_X1 u2_desIn_r_reg_53 (.CK( clk ) , .D( stage2_out_53 ) , .Q( u2_desIn_r_53 ) );
  DFF_X1 u2_desIn_r_reg_54 (.CK( clk ) , .D( stage2_out_54 ) , .Q( u2_desIn_r_54 ) );
  DFF_X1 u2_desIn_r_reg_55 (.CK( clk ) , .D( stage2_out_55 ) , .Q( u2_desIn_r_55 ) );
  DFF_X1 u2_desIn_r_reg_56 (.CK( clk ) , .D( stage2_out_56 ) , .Q( u2_desIn_r_56 ) );
  DFF_X1 u2_desIn_r_reg_57 (.CK( clk ) , .D( stage2_out_57 ) , .Q( u2_desIn_r_57 ) );
  DFF_X1 u2_desIn_r_reg_58 (.CK( clk ) , .D( stage2_out_58 ) , .Q( u2_desIn_r_58 ) );
  DFF_X1 u2_desIn_r_reg_59 (.CK( clk ) , .D( stage2_out_59 ) , .Q( u2_desIn_r_59 ) );
  DFF_X1 u2_desIn_r_reg_6 (.CK( clk ) , .D( stage2_out_6 ) , .Q( u2_desIn_r_6 ) );
  DFF_X1 u2_desIn_r_reg_60 (.CK( clk ) , .D( stage2_out_60 ) , .Q( u2_desIn_r_60 ) );
  DFF_X1 u2_desIn_r_reg_61 (.CK( clk ) , .D( stage2_out_61 ) , .Q( u2_desIn_r_61 ) );
  DFF_X1 u2_desIn_r_reg_62 (.CK( clk ) , .D( stage2_out_62 ) , .Q( u2_desIn_r_62 ) );
  DFF_X1 u2_desIn_r_reg_63 (.CK( clk ) , .D( stage2_out_63 ) , .Q( u2_desIn_r_63 ) );
  DFF_X1 u2_desIn_r_reg_7 (.CK( clk ) , .D( stage2_out_7 ) , .Q( u2_desIn_r_7 ) );
  DFF_X1 u2_desIn_r_reg_8 (.CK( clk ) , .D( stage2_out_8 ) , .Q( u2_desIn_r_8 ) );
  DFF_X1 u2_desIn_r_reg_9 (.CK( clk ) , .D( stage2_out_9 ) , .Q( u2_desIn_r_9 ) );
  DFF_X1 u2_desOut_reg_0 (.CK( clk ) , .Q( desOut[0] ) , .D( u2_FP_25 ) );
  DFF_X1 u2_desOut_reg_1 (.CK( clk ) , .Q( desOut[1] ) , .D( u2_FP_57 ) );
  DFF_X1 u2_desOut_reg_10 (.CK( clk ) , .Q( desOut[10] ) , .D( u2_FP_18 ) );
  DFF_X1 u2_desOut_reg_11 (.CK( clk ) , .Q( desOut[11] ) , .D( u2_FP_50 ) );
  DFF_X1 u2_desOut_reg_12 (.CK( clk ) , .Q( desOut[12] ) , .D( u2_FP_10 ) );
  DFF_X1 u2_desOut_reg_13 (.CK( clk ) , .Q( desOut[13] ) , .D( u2_FP_42 ) );
  DFF_X1 u2_desOut_reg_14 (.CK( clk ) , .Q( desOut[14] ) , .D( u2_FP_2 ) );
  DFF_X1 u2_desOut_reg_15 (.CK( clk ) , .Q( desOut[15] ) , .D( u2_FP_34 ) );
  DFF_X1 u2_desOut_reg_16 (.CK( clk ) , .Q( desOut[16] ) , .D( u2_FP_27 ) );
  DFF_X1 u2_desOut_reg_17 (.CK( clk ) , .Q( desOut[17] ) , .D( u2_FP_59 ) );
  DFF_X1 u2_desOut_reg_18 (.CK( clk ) , .Q( desOut[18] ) , .D( u2_FP_19 ) );
  DFF_X1 u2_desOut_reg_19 (.CK( clk ) , .Q( desOut[19] ) , .D( u2_FP_51 ) );
  DFF_X1 u2_desOut_reg_2 (.CK( clk ) , .Q( desOut[2] ) , .D( u2_FP_17 ) );
  DFF_X1 u2_desOut_reg_20 (.CK( clk ) , .Q( desOut[20] ) , .D( u2_FP_11 ) );
  DFF_X1 u2_desOut_reg_21 (.CK( clk ) , .Q( desOut[21] ) , .D( u2_FP_43 ) );
  DFF_X1 u2_desOut_reg_22 (.CK( clk ) , .Q( desOut[22] ) , .D( u2_FP_3 ) );
  DFF_X1 u2_desOut_reg_23 (.CK( clk ) , .Q( desOut[23] ) , .D( u2_FP_35 ) );
  DFF_X1 u2_desOut_reg_24 (.CK( clk ) , .Q( desOut[24] ) , .D( u2_FP_28 ) );
  DFF_X1 u2_desOut_reg_25 (.CK( clk ) , .Q( desOut[25] ) , .D( u2_FP_60 ) );
  DFF_X1 u2_desOut_reg_26 (.CK( clk ) , .Q( desOut[26] ) , .D( u2_FP_20 ) );
  DFF_X1 u2_desOut_reg_27 (.CK( clk ) , .Q( desOut[27] ) , .D( u2_FP_52 ) );
  DFF_X1 u2_desOut_reg_28 (.CK( clk ) , .Q( desOut[28] ) , .D( u2_FP_12 ) );
  DFF_X1 u2_desOut_reg_29 (.CK( clk ) , .Q( desOut[29] ) , .D( u2_FP_44 ) );
  DFF_X1 u2_desOut_reg_3 (.CK( clk ) , .Q( desOut[3] ) , .D( u2_FP_49 ) );
  DFF_X1 u2_desOut_reg_30 (.CK( clk ) , .Q( desOut[30] ) , .D( u2_FP_4 ) );
  DFF_X1 u2_desOut_reg_31 (.CK( clk ) , .Q( desOut[31] ) , .D( u2_FP_36 ) );
  DFF_X1 u2_desOut_reg_32 (.CK( clk ) , .Q( desOut[32] ) , .D( u2_FP_29 ) );
  DFF_X1 u2_desOut_reg_33 (.CK( clk ) , .Q( desOut[33] ) , .D( u2_FP_61 ) );
  DFF_X1 u2_desOut_reg_34 (.CK( clk ) , .Q( desOut[34] ) , .D( u2_FP_21 ) );
  DFF_X1 u2_desOut_reg_35 (.CK( clk ) , .Q( desOut[35] ) , .D( u2_FP_53 ) );
  DFF_X1 u2_desOut_reg_36 (.CK( clk ) , .Q( desOut[36] ) , .D( u2_FP_13 ) );
  DFF_X1 u2_desOut_reg_37 (.CK( clk ) , .Q( desOut[37] ) , .D( u2_FP_45 ) );
  DFF_X1 u2_desOut_reg_38 (.CK( clk ) , .Q( desOut[38] ) , .D( u2_FP_5 ) );
  DFF_X1 u2_desOut_reg_39 (.CK( clk ) , .Q( desOut[39] ) , .D( u2_FP_37 ) );
  DFF_X1 u2_desOut_reg_4 (.CK( clk ) , .Q( desOut[4] ) , .D( u2_FP_9 ) );
  DFF_X1 u2_desOut_reg_40 (.CK( clk ) , .Q( desOut[40] ) , .D( u2_FP_30 ) );
  DFF_X1 u2_desOut_reg_41 (.CK( clk ) , .Q( desOut[41] ) , .D( u2_FP_62 ) );
  DFF_X1 u2_desOut_reg_42 (.CK( clk ) , .Q( desOut[42] ) , .D( u2_FP_22 ) );
  DFF_X1 u2_desOut_reg_43 (.CK( clk ) , .Q( desOut[43] ) , .D( u2_FP_54 ) );
  DFF_X1 u2_desOut_reg_44 (.CK( clk ) , .Q( desOut[44] ) , .D( u2_FP_14 ) );
  DFF_X1 u2_desOut_reg_45 (.CK( clk ) , .Q( desOut[45] ) , .D( u2_FP_46 ) );
  DFF_X1 u2_desOut_reg_46 (.CK( clk ) , .Q( desOut[46] ) , .D( u2_FP_6 ) );
  DFF_X1 u2_desOut_reg_47 (.CK( clk ) , .Q( desOut[47] ) , .D( u2_FP_38 ) );
  DFF_X1 u2_desOut_reg_48 (.CK( clk ) , .Q( desOut[48] ) , .D( u2_FP_31 ) );
  DFF_X1 u2_desOut_reg_49 (.CK( clk ) , .Q( desOut[49] ) , .D( u2_FP_63 ) );
  DFF_X1 u2_desOut_reg_5 (.CK( clk ) , .Q( desOut[5] ) , .D( u2_FP_41 ) );
  DFF_X1 u2_desOut_reg_50 (.CK( clk ) , .Q( desOut[50] ) , .D( u2_FP_23 ) );
  DFF_X1 u2_desOut_reg_51 (.CK( clk ) , .Q( desOut[51] ) , .D( u2_FP_55 ) );
  DFF_X1 u2_desOut_reg_52 (.CK( clk ) , .Q( desOut[52] ) , .D( u2_FP_15 ) );
  DFF_X1 u2_desOut_reg_53 (.CK( clk ) , .Q( desOut[53] ) , .D( u2_FP_47 ) );
  DFF_X1 u2_desOut_reg_54 (.CK( clk ) , .Q( desOut[54] ) , .D( u2_FP_7 ) );
  DFF_X1 u2_desOut_reg_55 (.CK( clk ) , .Q( desOut[55] ) , .D( u2_FP_39 ) );
  DFF_X1 u2_desOut_reg_56 (.CK( clk ) , .Q( desOut[56] ) , .D( u2_FP_32 ) );
  DFF_X1 u2_desOut_reg_57 (.CK( clk ) , .Q( desOut[57] ) , .D( u2_FP_64 ) );
  DFF_X1 u2_desOut_reg_58 (.CK( clk ) , .Q( desOut[58] ) , .D( u2_FP_24 ) );
  DFF_X1 u2_desOut_reg_59 (.CK( clk ) , .Q( desOut[59] ) , .D( u2_FP_56 ) );
  DFF_X1 u2_desOut_reg_6 (.CK( clk ) , .Q( desOut[6] ) , .D( u2_FP_1 ) );
  DFF_X1 u2_desOut_reg_60 (.CK( clk ) , .Q( desOut[60] ) , .D( u2_FP_16 ) );
  DFF_X1 u2_desOut_reg_61 (.CK( clk ) , .Q( desOut[61] ) , .D( u2_FP_48 ) );
  DFF_X1 u2_desOut_reg_62 (.CK( clk ) , .Q( desOut[62] ) , .D( u2_FP_8 ) );
  DFF_X1 u2_desOut_reg_63 (.CK( clk ) , .Q( desOut[63] ) , .D( u2_FP_40 ) );
  DFF_X1 u2_desOut_reg_7 (.CK( clk ) , .Q( desOut[7] ) , .D( u2_FP_33 ) );
  DFF_X1 u2_desOut_reg_8 (.CK( clk ) , .Q( desOut[8] ) , .D( u2_FP_26 ) );
  DFF_X1 u2_desOut_reg_9 (.CK( clk ) , .Q( desOut[9] ) , .D( u2_FP_58 ) );
  DFF_X1 u2_key_r_reg_0 (.CK( clk ) , .D( key_c_r_33_0 ) , .Q( u2_key_r_0 ) );
  DFF_X1 u2_key_r_reg_1 (.CK( clk ) , .D( key_c_r_33_1 ) , .Q( u2_key_r_1 ) );
  DFF_X1 u2_key_r_reg_10 (.CK( clk ) , .D( key_c_r_33_10 ) , .Q( u2_key_r_10 ) );
  DFF_X1 u2_key_r_reg_11 (.CK( clk ) , .D( key_c_r_33_11 ) , .Q( u2_key_r_11 ) );
  DFF_X1 u2_key_r_reg_12 (.CK( clk ) , .D( key_c_r_33_12 ) , .Q( u2_key_r_12 ) );
  DFF_X1 u2_key_r_reg_13 (.CK( clk ) , .D( key_c_r_33_13 ) , .Q( u2_key_r_13 ) );
  DFF_X1 u2_key_r_reg_14 (.CK( clk ) , .D( key_c_r_33_14 ) , .Q( u2_key_r_14 ) );
  DFF_X1 u2_key_r_reg_15 (.CK( clk ) , .D( key_c_r_33_15 ) , .Q( u2_key_r_15 ) );
  DFF_X1 u2_key_r_reg_16 (.CK( clk ) , .D( key_c_r_33_16 ) , .Q( u2_key_r_16 ) );
  DFF_X1 u2_key_r_reg_17 (.CK( clk ) , .D( key_c_r_33_17 ) , .Q( u2_key_r_17 ) );
  DFF_X1 u2_key_r_reg_18 (.CK( clk ) , .D( key_c_r_33_18 ) , .Q( u2_key_r_18 ) );
  DFF_X1 u2_key_r_reg_19 (.CK( clk ) , .D( key_c_r_33_19 ) , .Q( u2_key_r_19 ) );
  DFF_X1 u2_key_r_reg_2 (.CK( clk ) , .D( key_c_r_33_2 ) , .Q( u2_key_r_2 ) );
  DFF_X1 u2_key_r_reg_20 (.CK( clk ) , .D( key_c_r_33_20 ) , .Q( u2_key_r_20 ) );
  DFF_X1 u2_key_r_reg_21 (.CK( clk ) , .D( key_c_r_33_21 ) , .Q( u2_key_r_21 ) );
  DFF_X1 u2_key_r_reg_22 (.CK( clk ) , .D( key_c_r_33_22 ) , .Q( u2_key_r_22 ) );
  DFF_X1 u2_key_r_reg_23 (.CK( clk ) , .D( key_c_r_33_23 ) , .Q( u2_key_r_23 ) );
  DFF_X1 u2_key_r_reg_24 (.CK( clk ) , .D( key_c_r_33_24 ) , .Q( u2_key_r_24 ) );
  DFF_X1 u2_key_r_reg_25 (.CK( clk ) , .D( key_c_r_33_25 ) , .Q( u2_key_r_25 ) );
  DFF_X1 u2_key_r_reg_26 (.CK( clk ) , .D( key_c_r_33_26 ) , .Q( u2_key_r_26 ) );
  DFF_X1 u2_key_r_reg_27 (.CK( clk ) , .D( key_c_r_33_27 ) , .Q( u2_key_r_27 ) );
  DFF_X1 u2_key_r_reg_28 (.CK( clk ) , .D( key_c_r_33_28 ) , .Q( u2_key_r_28 ) );
  DFF_X1 u2_key_r_reg_29 (.CK( clk ) , .D( key_c_r_33_29 ) , .Q( u2_key_r_29 ) );
  DFF_X1 u2_key_r_reg_3 (.CK( clk ) , .D( key_c_r_33_3 ) , .Q( u2_key_r_3 ) );
  DFF_X1 u2_key_r_reg_30 (.CK( clk ) , .D( key_c_r_33_30 ) , .Q( u2_key_r_30 ) );
  DFF_X1 u2_key_r_reg_31 (.CK( clk ) , .D( key_c_r_33_31 ) , .Q( u2_key_r_31 ) );
  DFF_X1 u2_key_r_reg_32 (.CK( clk ) , .D( key_c_r_33_32 ) , .Q( u2_key_r_32 ) );
  DFF_X1 u2_key_r_reg_33 (.CK( clk ) , .D( key_c_r_33_33 ) , .Q( u2_key_r_33 ) );
  DFF_X1 u2_key_r_reg_34 (.CK( clk ) , .D( key_c_r_33_34 ) , .Q( u2_key_r_34 ) );
  DFF_X1 u2_key_r_reg_35 (.CK( clk ) , .D( key_c_r_33_35 ) , .Q( u2_key_r_35 ) );
  DFF_X1 u2_key_r_reg_36 (.CK( clk ) , .D( key_c_r_33_36 ) , .Q( u2_key_r_36 ) );
  DFF_X1 u2_key_r_reg_37 (.CK( clk ) , .D( key_c_r_33_37 ) , .Q( u2_key_r_37 ) );
  DFF_X1 u2_key_r_reg_38 (.CK( clk ) , .D( key_c_r_33_38 ) , .Q( u2_key_r_38 ) );
  DFF_X1 u2_key_r_reg_39 (.CK( clk ) , .D( key_c_r_33_39 ) , .Q( u2_key_r_39 ) );
  DFF_X1 u2_key_r_reg_4 (.CK( clk ) , .D( key_c_r_33_4 ) , .Q( u2_key_r_4 ) );
  DFF_X1 u2_key_r_reg_40 (.CK( clk ) , .D( key_c_r_33_40 ) , .Q( u2_key_r_40 ) );
  DFF_X1 u2_key_r_reg_41 (.CK( clk ) , .D( key_c_r_33_41 ) , .Q( u2_key_r_41 ) );
  DFF_X1 u2_key_r_reg_42 (.CK( clk ) , .D( key_c_r_33_42 ) , .Q( u2_key_r_42 ) );
  DFF_X1 u2_key_r_reg_43 (.CK( clk ) , .D( key_c_r_33_43 ) , .Q( u2_key_r_43 ) );
  DFF_X1 u2_key_r_reg_44 (.CK( clk ) , .D( key_c_r_33_44 ) , .Q( u2_key_r_44 ) );
  DFF_X1 u2_key_r_reg_45 (.CK( clk ) , .D( key_c_r_33_45 ) , .Q( u2_key_r_45 ) );
  DFF_X1 u2_key_r_reg_46 (.CK( clk ) , .D( key_c_r_33_46 ) , .Q( u2_key_r_46 ) );
  DFF_X1 u2_key_r_reg_47 (.CK( clk ) , .D( key_c_r_33_47 ) , .Q( u2_key_r_47 ) );
  DFF_X1 u2_key_r_reg_48 (.CK( clk ) , .D( key_c_r_33_48 ) , .Q( u2_key_r_48 ) );
  DFF_X1 u2_key_r_reg_49 (.CK( clk ) , .D( key_c_r_33_49 ) , .Q( u2_key_r_49 ) );
  DFF_X1 u2_key_r_reg_5 (.CK( clk ) , .D( key_c_r_33_5 ) , .Q( u2_key_r_5 ) );
  DFF_X1 u2_key_r_reg_50 (.CK( clk ) , .D( key_c_r_33_50 ) , .Q( u2_key_r_50 ) );
  DFF_X1 u2_key_r_reg_51 (.CK( clk ) , .D( key_c_r_33_51 ) , .Q( u2_key_r_51 ) );
  DFF_X1 u2_key_r_reg_52 (.CK( clk ) , .D( key_c_r_33_52 ) , .Q( u2_key_r_52 ) );
  DFF_X1 u2_key_r_reg_53 (.CK( clk ) , .D( key_c_r_33_53 ) , .Q( u2_key_r_53 ) );
  DFF_X1 u2_key_r_reg_54 (.CK( clk ) , .D( key_c_r_33_54 ) , .Q( u2_key_r_54 ) );
  DFF_X1 u2_key_r_reg_55 (.CK( clk ) , .D( key_c_r_33_55 ) , .Q( u2_key_r_55 ) );
  DFF_X1 u2_key_r_reg_6 (.CK( clk ) , .D( key_c_r_33_6 ) , .Q( u2_key_r_6 ) );
  DFF_X1 u2_key_r_reg_7 (.CK( clk ) , .D( key_c_r_33_7 ) , .Q( u2_key_r_7 ) );
  DFF_X1 u2_key_r_reg_8 (.CK( clk ) , .D( key_c_r_33_8 ) , .Q( u2_key_r_8 ) );
  DFF_X1 u2_key_r_reg_9 (.CK( clk ) , .D( key_c_r_33_9 ) , .Q( u2_key_r_9 ) );
  DFF_X1 u2_uk_K_r0_reg_0 (.CK( clk ) , .D( u2_key_r_0 ) , .Q( u2_uk_K_r0_0 ) , .QN( u2_uk_n1230 ) );
  DFF_X1 u2_uk_K_r0_reg_1 (.CK( clk ) , .D( u2_key_r_1 ) , .Q( u2_uk_K_r0_1 ) );
  DFF_X1 u2_uk_K_r0_reg_10 (.CK( clk ) , .D( u2_key_r_10 ) , .Q( u2_uk_K_r0_10 ) , .QN( u2_uk_n1238 ) );
  DFF_X1 u2_uk_K_r0_reg_11 (.CK( clk ) , .D( u2_key_r_11 ) , .Q( u2_uk_K_r0_11 ) );
  DFF_X1 u2_uk_K_r0_reg_12 (.CK( clk ) , .D( u2_key_r_12 ) , .Q( u2_uk_K_r0_12 ) , .QN( u2_uk_n1239 ) );
  DFF_X1 u2_uk_K_r0_reg_13 (.CK( clk ) , .D( u2_key_r_13 ) , .Q( u2_uk_K_r0_13 ) , .QN( u2_uk_n1240 ) );
  DFF_X1 u2_uk_K_r0_reg_14 (.CK( clk ) , .D( u2_key_r_14 ) , .Q( u2_uk_K_r0_14 ) , .QN( u2_uk_n1241 ) );
  DFF_X1 u2_uk_K_r0_reg_15 (.CK( clk ) , .D( u2_key_r_15 ) , .Q( u2_uk_K_r0_15 ) );
  DFF_X1 u2_uk_K_r0_reg_16 (.CK( clk ) , .D( u2_key_r_16 ) , .Q( u2_uk_K_r0_16 ) , .QN( u2_uk_n1242 ) );
  DFF_X1 u2_uk_K_r0_reg_17 (.CK( clk ) , .D( u2_key_r_17 ) , .Q( u2_uk_K_r0_17 ) );
  DFF_X1 u2_uk_K_r0_reg_18 (.CK( clk ) , .D( u2_key_r_18 ) , .Q( u2_uk_K_r0_18 ) , .QN( u2_uk_n1243 ) );
  DFF_X1 u2_uk_K_r0_reg_19 (.CK( clk ) , .D( u2_key_r_19 ) , .Q( u2_uk_K_r0_19 ) );
  DFF_X1 u2_uk_K_r0_reg_2 (.CK( clk ) , .D( u2_key_r_2 ) , .Q( u2_uk_K_r0_2 ) );
  DFF_X1 u2_uk_K_r0_reg_20 (.CK( clk ) , .D( u2_key_r_20 ) , .Q( u2_uk_K_r0_20 ) , .QN( u2_uk_n1244 ) );
  DFF_X1 u2_uk_K_r0_reg_21 (.CK( clk ) , .D( u2_key_r_21 ) , .Q( u2_uk_K_r0_21 ) , .QN( u2_uk_n1245 ) );
  DFF_X1 u2_uk_K_r0_reg_22 (.CK( clk ) , .D( u2_key_r_22 ) , .Q( u2_uk_K_r0_22 ) );
  DFF_X1 u2_uk_K_r0_reg_23 (.CK( clk ) , .D( u2_key_r_23 ) , .Q( u2_uk_K_r0_23 ) , .QN( u2_uk_n1246 ) );
  DFF_X1 u2_uk_K_r0_reg_24 (.CK( clk ) , .D( u2_key_r_24 ) , .Q( u2_uk_K_r0_24 ) , .QN( u2_uk_n1247 ) );
  DFF_X1 u2_uk_K_r0_reg_25 (.CK( clk ) , .D( u2_key_r_25 ) , .Q( u2_uk_K_r0_25 ) );
  DFF_X1 u2_uk_K_r0_reg_26 (.CK( clk ) , .D( u2_key_r_26 ) , .Q( u2_uk_K_r0_26 ) , .QN( u2_uk_n1248 ) );
  DFF_X1 u2_uk_K_r0_reg_27 (.CK( clk ) , .D( u2_key_r_27 ) , .Q( u2_uk_K_r0_27 ) , .QN( u2_uk_n1249 ) );
  DFF_X1 u2_uk_K_r0_reg_28 (.CK( clk ) , .D( u2_key_r_28 ) , .Q( u2_uk_K_r0_28 ) );
  DFF_X1 u2_uk_K_r0_reg_29 (.CK( clk ) , .D( u2_key_r_29 ) , .Q( u2_uk_K_r0_29 ) , .QN( u2_uk_n1251 ) );
  DFF_X1 u2_uk_K_r0_reg_3 (.CK( clk ) , .D( u2_key_r_3 ) , .Q( u2_uk_K_r0_3 ) , .QN( u2_uk_n1231 ) );
  DFF_X1 u2_uk_K_r0_reg_30 (.CK( clk ) , .D( u2_key_r_30 ) , .Q( u2_uk_K_r0_30 ) , .QN( u2_uk_n1252 ) );
  DFF_X1 u2_uk_K_r0_reg_31 (.CK( clk ) , .D( u2_key_r_31 ) , .Q( u2_uk_K_r0_31 ) );
  DFF_X1 u2_uk_K_r0_reg_32 (.CK( clk ) , .D( u2_key_r_32 ) , .Q( u2_uk_K_r0_32 ) );
  DFF_X1 u2_uk_K_r0_reg_33 (.CK( clk ) , .D( u2_key_r_33 ) , .Q( u2_uk_K_r0_33 ) , .QN( u2_uk_n1254 ) );
  DFF_X1 u2_uk_K_r0_reg_34 (.CK( clk ) , .D( u2_key_r_34 ) , .Q( u2_uk_K_r0_34 ) );
  DFF_X1 u2_uk_K_r0_reg_35 (.CK( clk ) , .D( u2_key_r_35 ) , .Q( u2_uk_K_r0_35 ) , .QN( u2_uk_n1256 ) );
  DFF_X1 u2_uk_K_r0_reg_36 (.CK( clk ) , .D( u2_key_r_36 ) , .Q( u2_uk_K_r0_36 ) );
  DFF_X1 u2_uk_K_r0_reg_37 (.CK( clk ) , .D( u2_key_r_37 ) , .Q( u2_uk_K_r0_37 ) , .QN( u2_uk_n1258 ) );
  DFF_X1 u2_uk_K_r0_reg_38 (.CK( clk ) , .D( u2_key_r_38 ) , .Q( u2_uk_K_r0_38 ) , .QN( u2_uk_n1259 ) );
  DFF_X1 u2_uk_K_r0_reg_39 (.CK( clk ) , .D( u2_key_r_39 ) , .Q( u2_uk_K_r0_39 ) , .QN( u2_uk_n1260 ) );
  DFF_X1 u2_uk_K_r0_reg_4 (.CK( clk ) , .D( u2_key_r_4 ) , .Q( u2_uk_K_r0_4 ) , .QN( u2_uk_n1232 ) );
  DFF_X1 u2_uk_K_r0_reg_40 (.CK( clk ) , .D( u2_key_r_40 ) , .Q( u2_uk_K_r0_40 ) , .QN( u2_uk_n1261 ) );
  DFF_X1 u2_uk_K_r0_reg_41 (.CK( clk ) , .D( u2_key_r_41 ) , .Q( u2_uk_K_r0_41 ) , .QN( u2_uk_n1262 ) );
  DFF_X1 u2_uk_K_r0_reg_42 (.CK( clk ) , .D( u2_key_r_42 ) , .Q( u2_uk_K_r0_42 ) , .QN( u2_uk_n1263 ) );
  DFF_X1 u2_uk_K_r0_reg_43 (.CK( clk ) , .D( u2_key_r_43 ) , .Q( u2_uk_K_r0_43 ) , .QN( u2_uk_n1264 ) );
  DFF_X1 u2_uk_K_r0_reg_44 (.CK( clk ) , .D( u2_key_r_44 ) , .Q( u2_uk_K_r0_44 ) , .QN( u2_uk_n1265 ) );
  DFF_X1 u2_uk_K_r0_reg_45 (.CK( clk ) , .D( u2_key_r_45 ) , .Q( u2_uk_K_r0_45 ) , .QN( u2_uk_n1266 ) );
  DFF_X1 u2_uk_K_r0_reg_46 (.CK( clk ) , .D( u2_key_r_46 ) , .Q( u2_uk_K_r0_46 ) , .QN( u2_uk_n1267 ) );
  DFF_X1 u2_uk_K_r0_reg_47 (.CK( clk ) , .D( u2_key_r_47 ) , .Q( u2_uk_K_r0_47 ) , .QN( u2_uk_n1269 ) );
  DFF_X1 u2_uk_K_r0_reg_48 (.CK( clk ) , .D( u2_key_r_48 ) , .Q( u2_uk_K_r0_48 ) , .QN( u2_uk_n1270 ) );
  DFF_X1 u2_uk_K_r0_reg_49 (.CK( clk ) , .D( u2_key_r_49 ) , .Q( u2_uk_K_r0_49 ) );
  DFF_X1 u2_uk_K_r0_reg_5 (.CK( clk ) , .D( u2_key_r_5 ) , .Q( u2_uk_K_r0_5 ) , .QN( u2_uk_n1233 ) );
  DFF_X1 u2_uk_K_r0_reg_50 (.CK( clk ) , .D( u2_key_r_50 ) , .Q( u2_uk_K_r0_50 ) , .QN( u2_uk_n1273 ) );
  DFF_X1 u2_uk_K_r0_reg_51 (.CK( clk ) , .D( u2_key_r_51 ) , .Q( u2_uk_K_r0_51 ) , .QN( u2_uk_n1274 ) );
  DFF_X1 u2_uk_K_r0_reg_52 (.CK( clk ) , .D( u2_key_r_52 ) , .Q( u2_uk_K_r0_52 ) );
  DFF_X1 u2_uk_K_r0_reg_53 (.CK( clk ) , .D( u2_key_r_53 ) , .Q( u2_uk_K_r0_53 ) );
  DFF_X1 u2_uk_K_r0_reg_54 (.CK( clk ) , .D( u2_key_r_54 ) , .Q( u2_uk_K_r0_54 ) , .QN( u2_uk_n1275 ) );
  DFF_X1 u2_uk_K_r0_reg_55 (.CK( clk ) , .D( u2_key_r_55 ) , .Q( u2_uk_K_r0_55 ) );
  DFF_X1 u2_uk_K_r0_reg_6 (.CK( clk ) , .D( u2_key_r_6 ) , .Q( u2_uk_K_r0_6 ) , .QN( u2_uk_n1234 ) );
  DFF_X1 u2_uk_K_r0_reg_7 (.CK( clk ) , .D( u2_key_r_7 ) , .Q( u2_uk_K_r0_7 ) , .QN( u2_uk_n1235 ) );
  DFF_X1 u2_uk_K_r0_reg_8 (.CK( clk ) , .D( u2_key_r_8 ) , .Q( u2_uk_K_r0_8 ) , .QN( u2_uk_n1236 ) );
  DFF_X1 u2_uk_K_r0_reg_9 (.CK( clk ) , .D( u2_key_r_9 ) , .Q( u2_uk_K_r0_9 ) , .QN( u2_uk_n1237 ) );
  DFF_X1 u2_uk_K_r10_reg_0 (.CK( clk ) , .Q( u2_uk_K_r10_0 ) , .D( u2_uk_K_r9_0 ) , .QN( u2_uk_n1678 ) );
  DFF_X1 u2_uk_K_r10_reg_1 (.CK( clk ) , .Q( u2_uk_K_r10_1 ) , .D( u2_uk_K_r9_1 ) , .QN( u2_uk_n1679 ) );
  DFF_X1 u2_uk_K_r10_reg_10 (.CK( clk ) , .Q( u2_uk_K_r10_10 ) , .D( u2_uk_K_r9_10 ) );
  DFF_X1 u2_uk_K_r10_reg_11 (.CK( clk ) , .Q( u2_uk_K_r10_11 ) , .D( u2_uk_K_r9_11 ) );
  DFF_X1 u2_uk_K_r10_reg_12 (.CK( clk ) , .Q( u2_uk_K_r10_12 ) , .D( u2_uk_K_r9_12 ) , .QN( u2_uk_n1686 ) );
  DFF_X1 u2_uk_K_r10_reg_13 (.CK( clk ) , .Q( u2_uk_K_r10_13 ) , .D( u2_uk_K_r9_13 ) );
  DFF_X1 u2_uk_K_r10_reg_14 (.CK( clk ) , .Q( u2_uk_K_r10_14 ) , .D( u2_uk_K_r9_14 ) );
  DFF_X1 u2_uk_K_r10_reg_15 (.CK( clk ) , .Q( u2_uk_K_r10_15 ) , .D( u2_uk_K_r9_15 ) , .QN( u2_uk_n1687 ) );
  DFF_X1 u2_uk_K_r10_reg_16 (.CK( clk ) , .Q( u2_uk_K_r10_16 ) , .D( u2_uk_K_r9_16 ) );
  DFF_X1 u2_uk_K_r10_reg_17 (.CK( clk ) , .Q( u2_uk_K_r10_17 ) , .D( u2_uk_K_r9_17 ) , .QN( u2_uk_n1688 ) );
  DFF_X1 u2_uk_K_r10_reg_18 (.CK( clk ) , .Q( u2_uk_K_r10_18 ) , .D( u2_uk_K_r9_18 ) );
  DFF_X1 u2_uk_K_r10_reg_19 (.CK( clk ) , .Q( u2_uk_K_r10_19 ) , .D( u2_uk_K_r9_19 ) );
  DFF_X1 u2_uk_K_r10_reg_2 (.CK( clk ) , .Q( u2_uk_K_r10_2 ) , .D( u2_uk_K_r9_2 ) , .QN( u2_uk_n1680 ) );
  DFF_X1 u2_uk_K_r10_reg_20 (.CK( clk ) , .Q( u2_uk_K_r10_20 ) , .D( u2_uk_K_r9_20 ) , .QN( u2_uk_n1689 ) );
  DFF_X1 u2_uk_K_r10_reg_21 (.CK( clk ) , .Q( u2_uk_K_r10_21 ) , .D( u2_uk_K_r9_21 ) , .QN( u2_uk_n1690 ) );
  DFF_X1 u2_uk_K_r10_reg_22 (.CK( clk ) , .Q( u2_uk_K_r10_22 ) , .D( u2_uk_K_r9_22 ) , .QN( u2_uk_n1691 ) );
  DFF_X1 u2_uk_K_r10_reg_23 (.CK( clk ) , .Q( u2_uk_K_r10_23 ) , .D( u2_uk_K_r9_23 ) );
  DFF_X1 u2_uk_K_r10_reg_24 (.CK( clk ) , .Q( u2_uk_K_r10_24 ) , .D( u2_uk_K_r9_24 ) , .QN( u2_uk_n1692 ) );
  DFF_X1 u2_uk_K_r10_reg_25 (.CK( clk ) , .Q( u2_uk_K_r10_25 ) , .D( u2_uk_K_r9_25 ) );
  DFF_X1 u2_uk_K_r10_reg_26 (.CK( clk ) , .Q( u2_uk_K_r10_26 ) , .D( u2_uk_K_r9_26 ) , .QN( u2_uk_n1693 ) );
  DFF_X1 u2_uk_K_r10_reg_27 (.CK( clk ) , .Q( u2_uk_K_r10_27 ) , .D( u2_uk_K_r9_27 ) );
  DFF_X1 u2_uk_K_r10_reg_28 (.CK( clk ) , .Q( u2_uk_K_r10_28 ) , .D( u2_uk_K_r9_28 ) );
  DFF_X1 u2_uk_K_r10_reg_29 (.CK( clk ) , .Q( u2_uk_K_r10_29 ) , .D( u2_uk_K_r9_29 ) , .QN( u2_uk_n1698 ) );
  DFF_X1 u2_uk_K_r10_reg_3 (.CK( clk ) , .Q( u2_uk_K_r10_3 ) , .D( u2_uk_K_r9_3 ) , .QN( u2_uk_n1681 ) );
  DFF_X1 u2_uk_K_r10_reg_30 (.CK( clk ) , .Q( u2_uk_K_r10_30 ) , .D( u2_uk_K_r9_30 ) , .QN( u2_uk_n1699 ) );
  DFF_X1 u2_uk_K_r10_reg_31 (.CK( clk ) , .Q( u2_uk_K_r10_31 ) , .D( u2_uk_K_r9_31 ) , .QN( u2_uk_n1700 ) );
  DFF_X1 u2_uk_K_r10_reg_32 (.CK( clk ) , .Q( u2_uk_K_r10_32 ) , .D( u2_uk_K_r9_32 ) , .QN( u2_uk_n1701 ) );
  DFF_X1 u2_uk_K_r10_reg_33 (.CK( clk ) , .Q( u2_uk_K_r10_33 ) , .D( u2_uk_K_r9_33 ) , .QN( u2_uk_n1702 ) );
  DFF_X1 u2_uk_K_r10_reg_34 (.CK( clk ) , .Q( u2_uk_K_r10_34 ) , .D( u2_uk_K_r9_34 ) );
  DFF_X1 u2_uk_K_r10_reg_35 (.CK( clk ) , .Q( u2_uk_K_r10_35 ) , .D( u2_uk_K_r9_35 ) , .QN( u2_uk_n1704 ) );
  DFF_X1 u2_uk_K_r10_reg_36 (.CK( clk ) , .Q( u2_uk_K_r10_36 ) , .D( u2_uk_K_r9_36 ) , .QN( u2_uk_n1705 ) );
  DFF_X1 u2_uk_K_r10_reg_37 (.CK( clk ) , .Q( u2_uk_K_r10_37 ) , .D( u2_uk_K_r9_37 ) , .QN( u2_uk_n1706 ) );
  DFF_X1 u2_uk_K_r10_reg_38 (.CK( clk ) , .Q( u2_uk_K_r10_38 ) , .D( u2_uk_K_r9_38 ) , .QN( u2_uk_n1707 ) );
  DFF_X1 u2_uk_K_r10_reg_39 (.CK( clk ) , .Q( u2_uk_K_r10_39 ) , .D( u2_uk_K_r9_39 ) , .QN( u2_uk_n1708 ) );
  DFF_X1 u2_uk_K_r10_reg_4 (.CK( clk ) , .Q( u2_uk_K_r10_4 ) , .D( u2_uk_K_r9_4 ) );
  DFF_X1 u2_uk_K_r10_reg_40 (.CK( clk ) , .Q( u2_uk_K_r10_40 ) , .D( u2_uk_K_r9_40 ) , .QN( u2_uk_n1709 ) );
  DFF_X1 u2_uk_K_r10_reg_41 (.CK( clk ) , .Q( u2_uk_K_r10_41 ) , .D( u2_uk_K_r9_41 ) );
  DFF_X1 u2_uk_K_r10_reg_42 (.CK( clk ) , .Q( u2_uk_K_r10_42 ) , .D( u2_uk_K_r9_42 ) );
  DFF_X1 u2_uk_K_r10_reg_43 (.CK( clk ) , .Q( u2_uk_K_r10_43 ) , .D( u2_uk_K_r9_43 ) );
  DFF_X1 u2_uk_K_r10_reg_44 (.CK( clk ) , .Q( u2_uk_K_r10_44 ) , .D( u2_uk_K_r9_44 ) );
  DFF_X1 u2_uk_K_r10_reg_45 (.CK( clk ) , .Q( u2_uk_K_r10_45 ) , .D( u2_uk_K_r9_45 ) , .QN( u2_uk_n1714 ) );
  DFF_X1 u2_uk_K_r10_reg_46 (.CK( clk ) , .Q( u2_uk_K_r10_46 ) , .D( u2_uk_K_r9_46 ) , .QN( u2_uk_n1715 ) );
  DFF_X1 u2_uk_K_r10_reg_47 (.CK( clk ) , .Q( u2_uk_K_r10_47 ) , .D( u2_uk_K_r9_47 ) );
  DFF_X1 u2_uk_K_r10_reg_48 (.CK( clk ) , .Q( u2_uk_K_r10_48 ) , .D( u2_uk_K_r9_48 ) );
  DFF_X1 u2_uk_K_r10_reg_49 (.CK( clk ) , .Q( u2_uk_K_r10_49 ) , .D( u2_uk_K_r9_49 ) );
  DFF_X1 u2_uk_K_r10_reg_5 (.CK( clk ) , .Q( u2_uk_K_r10_5 ) , .D( u2_uk_K_r9_5 ) , .QN( u2_uk_n1682 ) );
  DFF_X1 u2_uk_K_r10_reg_50 (.CK( clk ) , .Q( u2_uk_K_r10_50 ) , .D( u2_uk_K_r9_50 ) , .QN( u2_uk_n1718 ) );
  DFF_X1 u2_uk_K_r10_reg_51 (.CK( clk ) , .Q( u2_uk_K_r10_51 ) , .D( u2_uk_K_r9_51 ) , .QN( u2_uk_n1719 ) );
  DFF_X1 u2_uk_K_r10_reg_52 (.CK( clk ) , .Q( u2_uk_K_r10_52 ) , .D( u2_uk_K_r9_52 ) );
  DFF_X1 u2_uk_K_r10_reg_53 (.CK( clk ) , .Q( u2_uk_K_r10_53 ) , .D( u2_uk_K_r9_53 ) , .QN( u2_uk_n1720 ) );
  DFF_X1 u2_uk_K_r10_reg_54 (.CK( clk ) , .Q( u2_uk_K_r10_54 ) , .D( u2_uk_K_r9_54 ) , .QN( u2_uk_n1721 ) );
  DFF_X1 u2_uk_K_r10_reg_55 (.CK( clk ) , .Q( u2_uk_K_r10_55 ) , .D( u2_uk_K_r9_55 ) , .QN( u2_uk_n1722 ) );
  DFF_X1 u2_uk_K_r10_reg_6 (.CK( clk ) , .Q( u2_uk_K_r10_6 ) , .D( u2_uk_K_r9_6 ) , .QN( u2_uk_n1683 ) );
  DFF_X1 u2_uk_K_r10_reg_7 (.CK( clk ) , .Q( u2_uk_K_r10_7 ) , .D( u2_uk_K_r9_7 ) , .QN( u2_uk_n1684 ) );
  DFF_X1 u2_uk_K_r10_reg_8 (.CK( clk ) , .Q( u2_uk_K_r10_8 ) , .D( u2_uk_K_r9_8 ) , .QN( u2_uk_n1685 ) );
  DFF_X1 u2_uk_K_r10_reg_9 (.CK( clk ) , .Q( u2_uk_K_r10_9 ) , .D( u2_uk_K_r9_9 ) );
  DFF_X1 u2_uk_K_r11_reg_0 (.CK( clk ) , .D( u2_uk_K_r10_0 ) , .Q( u2_uk_K_r11_0 ) , .QN( u2_uk_n1723 ) );
  DFF_X1 u2_uk_K_r11_reg_1 (.CK( clk ) , .D( u2_uk_K_r10_1 ) , .Q( u2_uk_K_r11_1 ) , .QN( u2_uk_n1724 ) );
  DFF_X1 u2_uk_K_r11_reg_10 (.CK( clk ) , .D( u2_uk_K_r10_10 ) , .Q( u2_uk_K_r11_10 ) );
  DFF_X1 u2_uk_K_r11_reg_11 (.CK( clk ) , .D( u2_uk_K_r10_11 ) , .Q( u2_uk_K_r11_11 ) );
  DFF_X1 u2_uk_K_r11_reg_12 (.CK( clk ) , .D( u2_uk_K_r10_12 ) , .Q( u2_uk_K_r11_12 ) , .QN( u2_uk_n1731 ) );
  DFF_X1 u2_uk_K_r11_reg_13 (.CK( clk ) , .D( u2_uk_K_r10_13 ) , .Q( u2_uk_K_r11_13 ) , .QN( u2_uk_n1732 ) );
  DFF_X1 u2_uk_K_r11_reg_14 (.CK( clk ) , .D( u2_uk_K_r10_14 ) , .Q( u2_uk_K_r11_14 ) , .QN( u2_uk_n1733 ) );
  DFF_X1 u2_uk_K_r11_reg_15 (.CK( clk ) , .D( u2_uk_K_r10_15 ) , .Q( u2_uk_K_r11_15 ) , .QN( u2_uk_n1734 ) );
  DFF_X1 u2_uk_K_r11_reg_16 (.CK( clk ) , .D( u2_uk_K_r10_16 ) , .Q( u2_uk_K_r11_16 ) , .QN( u2_uk_n1735 ) );
  DFF_X1 u2_uk_K_r11_reg_17 (.CK( clk ) , .D( u2_uk_K_r10_17 ) , .Q( u2_uk_K_r11_17 ) , .QN( u2_uk_n1736 ) );
  DFF_X1 u2_uk_K_r11_reg_18 (.CK( clk ) , .D( u2_uk_K_r10_18 ) , .Q( u2_uk_K_r11_18 ) , .QN( u2_uk_n1737 ) );
  DFF_X1 u2_uk_K_r11_reg_19 (.CK( clk ) , .D( u2_uk_K_r10_19 ) , .Q( u2_uk_K_r11_19 ) );
  DFF_X1 u2_uk_K_r11_reg_2 (.CK( clk ) , .D( u2_uk_K_r10_2 ) , .Q( u2_uk_K_r11_2 ) , .QN( u2_uk_n1725 ) );
  DFF_X1 u2_uk_K_r11_reg_20 (.CK( clk ) , .D( u2_uk_K_r10_20 ) , .Q( u2_uk_K_r11_20 ) );
  DFF_X1 u2_uk_K_r11_reg_21 (.CK( clk ) , .D( u2_uk_K_r10_21 ) , .Q( u2_uk_K_r11_21 ) );
  DFF_X1 u2_uk_K_r11_reg_22 (.CK( clk ) , .D( u2_uk_K_r10_22 ) , .Q( u2_uk_K_r11_22 ) , .QN( u2_uk_n1738 ) );
  DFF_X1 u2_uk_K_r11_reg_23 (.CK( clk ) , .D( u2_uk_K_r10_23 ) , .Q( u2_uk_K_r11_23 ) , .QN( u2_uk_n1739 ) );
  DFF_X1 u2_uk_K_r11_reg_24 (.CK( clk ) , .D( u2_uk_K_r10_24 ) , .Q( u2_uk_K_r11_24 ) );
  DFF_X1 u2_uk_K_r11_reg_25 (.CK( clk ) , .D( u2_uk_K_r10_25 ) , .Q( u2_uk_K_r11_25 ) );
  DFF_X1 u2_uk_K_r11_reg_26 (.CK( clk ) , .D( u2_uk_K_r10_26 ) , .Q( u2_uk_K_r11_26 ) );
  DFF_X1 u2_uk_K_r11_reg_27 (.CK( clk ) , .D( u2_uk_K_r10_27 ) , .Q( u2_uk_K_r11_27 ) );
  DFF_X1 u2_uk_K_r11_reg_28 (.CK( clk ) , .D( u2_uk_K_r10_28 ) , .Q( u2_uk_K_r11_28 ) );
  DFF_X1 u2_uk_K_r11_reg_29 (.CK( clk ) , .D( u2_uk_K_r10_29 ) , .Q( u2_uk_K_r11_29 ) );
  DFF_X1 u2_uk_K_r11_reg_3 (.CK( clk ) , .D( u2_uk_K_r10_3 ) , .Q( u2_uk_K_r11_3 ) , .QN( u2_uk_n1726 ) );
  DFF_X1 u2_uk_K_r11_reg_30 (.CK( clk ) , .D( u2_uk_K_r10_30 ) , .Q( u2_uk_K_r11_30 ) );
  DFF_X1 u2_uk_K_r11_reg_31 (.CK( clk ) , .D( u2_uk_K_r10_31 ) , .Q( u2_uk_K_r11_31 ) , .QN( u2_uk_n1742 ) );
  DFF_X1 u2_uk_K_r11_reg_32 (.CK( clk ) , .D( u2_uk_K_r10_32 ) , .Q( u2_uk_K_r11_32 ) , .QN( u2_uk_n1743 ) );
  DFF_X1 u2_uk_K_r11_reg_33 (.CK( clk ) , .D( u2_uk_K_r10_33 ) , .Q( u2_uk_K_r11_33 ) );
  DFF_X1 u2_uk_K_r11_reg_34 (.CK( clk ) , .D( u2_uk_K_r10_34 ) , .Q( u2_uk_K_r11_34 ) );
  DFF_X1 u2_uk_K_r11_reg_35 (.CK( clk ) , .D( u2_uk_K_r10_35 ) , .Q( u2_uk_K_r11_35 ) , .QN( u2_uk_n1744 ) );
  DFF_X1 u2_uk_K_r11_reg_36 (.CK( clk ) , .D( u2_uk_K_r10_36 ) , .Q( u2_uk_K_r11_36 ) , .QN( u2_uk_n1745 ) );
  DFF_X1 u2_uk_K_r11_reg_37 (.CK( clk ) , .D( u2_uk_K_r10_37 ) , .Q( u2_uk_K_r11_37 ) , .QN( u2_uk_n1746 ) );
  DFF_X1 u2_uk_K_r11_reg_38 (.CK( clk ) , .D( u2_uk_K_r10_38 ) , .Q( u2_uk_K_r11_38 ) , .QN( u2_uk_n1747 ) );
  DFF_X1 u2_uk_K_r11_reg_39 (.CK( clk ) , .D( u2_uk_K_r10_39 ) , .Q( u2_uk_K_r11_39 ) );
  DFF_X1 u2_uk_K_r11_reg_4 (.CK( clk ) , .D( u2_uk_K_r10_4 ) , .Q( u2_uk_K_r11_4 ) );
  DFF_X1 u2_uk_K_r11_reg_40 (.CK( clk ) , .D( u2_uk_K_r10_40 ) , .Q( u2_uk_K_r11_40 ) , .QN( u2_uk_n1750 ) );
  DFF_X1 u2_uk_K_r11_reg_41 (.CK( clk ) , .D( u2_uk_K_r10_41 ) , .Q( u2_uk_K_r11_41 ) , .QN( u2_uk_n1751 ) );
  DFF_X1 u2_uk_K_r11_reg_42 (.CK( clk ) , .D( u2_uk_K_r10_42 ) , .Q( u2_uk_K_r11_42 ) , .QN( u2_uk_n1752 ) );
  DFF_X1 u2_uk_K_r11_reg_43 (.CK( clk ) , .D( u2_uk_K_r10_43 ) , .Q( u2_uk_K_r11_43 ) , .QN( u2_uk_n1753 ) );
  DFF_X1 u2_uk_K_r11_reg_44 (.CK( clk ) , .D( u2_uk_K_r10_44 ) , .Q( u2_uk_K_r11_44 ) , .QN( u2_uk_n1754 ) );
  DFF_X1 u2_uk_K_r11_reg_45 (.CK( clk ) , .D( u2_uk_K_r10_45 ) , .Q( u2_uk_K_r11_45 ) , .QN( u2_uk_n1755 ) );
  DFF_X1 u2_uk_K_r11_reg_46 (.CK( clk ) , .D( u2_uk_K_r10_46 ) , .Q( u2_uk_K_r11_46 ) , .QN( u2_uk_n1757 ) );
  DFF_X1 u2_uk_K_r11_reg_47 (.CK( clk ) , .D( u2_uk_K_r10_47 ) , .Q( u2_uk_K_r11_47 ) );
  DFF_X1 u2_uk_K_r11_reg_48 (.CK( clk ) , .D( u2_uk_K_r10_48 ) , .Q( u2_uk_K_r11_48 ) );
  DFF_X1 u2_uk_K_r11_reg_49 (.CK( clk ) , .D( u2_uk_K_r10_49 ) , .Q( u2_uk_K_r11_49 ) , .QN( u2_uk_n1760 ) );
  DFF_X1 u2_uk_K_r11_reg_5 (.CK( clk ) , .D( u2_uk_K_r10_5 ) , .Q( u2_uk_K_r11_5 ) , .QN( u2_uk_n1727 ) );
  DFF_X1 u2_uk_K_r11_reg_50 (.CK( clk ) , .D( u2_uk_K_r10_50 ) , .Q( u2_uk_K_r11_50 ) , .QN( u2_uk_n1761 ) );
  DFF_X1 u2_uk_K_r11_reg_51 (.CK( clk ) , .D( u2_uk_K_r10_51 ) , .Q( u2_uk_K_r11_51 ) , .QN( u2_uk_n1762 ) );
  DFF_X1 u2_uk_K_r11_reg_52 (.CK( clk ) , .D( u2_uk_K_r10_52 ) , .Q( u2_uk_K_r11_52 ) , .QN( u2_uk_n1763 ) );
  DFF_X1 u2_uk_K_r11_reg_53 (.CK( clk ) , .D( u2_uk_K_r10_53 ) , .Q( u2_uk_K_r11_53 ) );
  DFF_X1 u2_uk_K_r11_reg_54 (.CK( clk ) , .D( u2_uk_K_r10_54 ) , .Q( u2_uk_K_r11_54 ) );
  DFF_X1 u2_uk_K_r11_reg_55 (.CK( clk ) , .D( u2_uk_K_r10_55 ) , .Q( u2_uk_K_r11_55 ) , .QN( u2_uk_n1767 ) );
  DFF_X1 u2_uk_K_r11_reg_6 (.CK( clk ) , .D( u2_uk_K_r10_6 ) , .Q( u2_uk_K_r11_6 ) );
  DFF_X1 u2_uk_K_r11_reg_7 (.CK( clk ) , .D( u2_uk_K_r10_7 ) , .Q( u2_uk_K_r11_7 ) );
  DFF_X1 u2_uk_K_r11_reg_8 (.CK( clk ) , .D( u2_uk_K_r10_8 ) , .Q( u2_uk_K_r11_8 ) );
  DFF_X1 u2_uk_K_r11_reg_9 (.CK( clk ) , .D( u2_uk_K_r10_9 ) , .Q( u2_uk_K_r11_9 ) , .QN( u2_uk_n1728 ) );
  DFF_X1 u2_uk_K_r12_reg_0 (.CK( clk ) , .D( u2_uk_K_r11_0 ) , .Q( u2_uk_K_r12_0 ) , .QN( u2_uk_n1768 ) );
  DFF_X1 u2_uk_K_r12_reg_1 (.CK( clk ) , .D( u2_uk_K_r11_1 ) , .Q( u2_uk_K_r12_1 ) , .QN( u2_uk_n1769 ) );
  DFF_X1 u2_uk_K_r12_reg_10 (.CK( clk ) , .D( u2_uk_K_r11_10 ) , .Q( u2_uk_K_r12_10 ) );
  DFF_X1 u2_uk_K_r12_reg_11 (.CK( clk ) , .D( u2_uk_K_r11_11 ) , .Q( u2_uk_K_r12_11 ) , .QN( u2_uk_n1778 ) );
  DFF_X1 u2_uk_K_r12_reg_12 (.CK( clk ) , .D( u2_uk_K_r11_12 ) , .Q( u2_uk_K_r12_12 ) , .QN( u2_uk_n1779 ) );
  DFF_X1 u2_uk_K_r12_reg_13 (.CK( clk ) , .D( u2_uk_K_r11_13 ) , .Q( u2_uk_K_r12_13 ) , .QN( u2_uk_n1780 ) );
  DFF_X1 u2_uk_K_r12_reg_14 (.CK( clk ) , .D( u2_uk_K_r11_14 ) , .Q( u2_uk_K_r12_14 ) , .QN( u2_uk_n1781 ) );
  DFF_X1 u2_uk_K_r12_reg_15 (.CK( clk ) , .D( u2_uk_K_r11_15 ) , .Q( u2_uk_K_r12_15 ) );
  DFF_X1 u2_uk_K_r12_reg_16 (.CK( clk ) , .D( u2_uk_K_r11_16 ) , .Q( u2_uk_K_r12_16 ) );
  DFF_X1 u2_uk_K_r12_reg_17 (.CK( clk ) , .D( u2_uk_K_r11_17 ) , .Q( u2_uk_K_r12_17 ) , .QN( u2_uk_n1782 ) );
  DFF_X1 u2_uk_K_r12_reg_18 (.CK( clk ) , .D( u2_uk_K_r11_18 ) , .Q( u2_uk_K_r12_18 ) );
  DFF_X1 u2_uk_K_r12_reg_19 (.CK( clk ) , .D( u2_uk_K_r11_19 ) , .Q( u2_uk_K_r12_19 ) , .QN( u2_uk_n1783 ) );
  DFF_X1 u2_uk_K_r12_reg_2 (.CK( clk ) , .D( u2_uk_K_r11_2 ) , .Q( u2_uk_K_r12_2 ) , .QN( u2_uk_n1770 ) );
  DFF_X1 u2_uk_K_r12_reg_20 (.CK( clk ) , .D( u2_uk_K_r11_20 ) , .Q( u2_uk_K_r12_20 ) , .QN( u2_uk_n1784 ) );
  DFF_X1 u2_uk_K_r12_reg_21 (.CK( clk ) , .D( u2_uk_K_r11_21 ) , .Q( u2_uk_K_r12_21 ) );
  DFF_X1 u2_uk_K_r12_reg_22 (.CK( clk ) , .D( u2_uk_K_r11_22 ) , .Q( u2_uk_K_r12_22 ) );
  DFF_X1 u2_uk_K_r12_reg_23 (.CK( clk ) , .D( u2_uk_K_r11_23 ) , .Q( u2_uk_K_r12_23 ) , .QN( u2_uk_n1785 ) );
  DFF_X1 u2_uk_K_r12_reg_24 (.CK( clk ) , .D( u2_uk_K_r11_24 ) , .Q( u2_uk_K_r12_24 ) , .QN( u2_uk_n1786 ) );
  DFF_X1 u2_uk_K_r12_reg_25 (.CK( clk ) , .D( u2_uk_K_r11_25 ) , .Q( u2_uk_K_r12_25 ) , .QN( u2_uk_n1787 ) );
  DFF_X1 u2_uk_K_r12_reg_26 (.CK( clk ) , .D( u2_uk_K_r11_26 ) , .Q( u2_uk_K_r12_26 ) , .QN( u2_uk_n1788 ) );
  DFF_X1 u2_uk_K_r12_reg_27 (.CK( clk ) , .D( u2_uk_K_r11_27 ) , .Q( u2_uk_K_r12_27 ) , .QN( u2_uk_n1789 ) );
  DFF_X1 u2_uk_K_r12_reg_28 (.CK( clk ) , .D( u2_uk_K_r11_28 ) , .Q( u2_uk_K_r12_28 ) , .QN( u2_uk_n1790 ) );
  DFF_X1 u2_uk_K_r12_reg_29 (.CK( clk ) , .D( u2_uk_K_r11_29 ) , .Q( u2_uk_K_r12_29 ) , .QN( u2_uk_n1791 ) );
  DFF_X1 u2_uk_K_r12_reg_3 (.CK( clk ) , .D( u2_uk_K_r11_3 ) , .Q( u2_uk_K_r12_3 ) , .QN( u2_uk_n1771 ) );
  DFF_X1 u2_uk_K_r12_reg_30 (.CK( clk ) , .D( u2_uk_K_r11_30 ) , .Q( u2_uk_K_r12_30 ) , .QN( u2_uk_n1792 ) );
  DFF_X1 u2_uk_K_r12_reg_31 (.CK( clk ) , .D( u2_uk_K_r11_31 ) , .Q( u2_uk_K_r12_31 ) , .QN( u2_uk_n1793 ) );
  DFF_X1 u2_uk_K_r12_reg_32 (.CK( clk ) , .D( u2_uk_K_r11_32 ) , .Q( u2_uk_K_r12_32 ) , .QN( u2_uk_n1794 ) );
  DFF_X1 u2_uk_K_r12_reg_33 (.CK( clk ) , .D( u2_uk_K_r11_33 ) , .Q( u2_uk_K_r12_33 ) );
  DFF_X1 u2_uk_K_r12_reg_34 (.CK( clk ) , .D( u2_uk_K_r11_34 ) , .Q( u2_uk_K_r12_34 ) , .QN( u2_uk_n1796 ) );
  DFF_X1 u2_uk_K_r12_reg_35 (.CK( clk ) , .D( u2_uk_K_r11_35 ) , .Q( u2_uk_K_r12_35 ) , .QN( u2_uk_n1797 ) );
  DFF_X1 u2_uk_K_r12_reg_36 (.CK( clk ) , .D( u2_uk_K_r11_36 ) , .Q( u2_uk_K_r12_36 ) );
  DFF_X1 u2_uk_K_r12_reg_37 (.CK( clk ) , .D( u2_uk_K_r11_37 ) , .Q( u2_uk_K_r12_37 ) , .QN( u2_uk_n1799 ) );
  DFF_X1 u2_uk_K_r12_reg_38 (.CK( clk ) , .D( u2_uk_K_r11_38 ) , .Q( u2_uk_K_r12_38 ) , .QN( u2_uk_n1800 ) );
  DFF_X1 u2_uk_K_r12_reg_39 (.CK( clk ) , .D( u2_uk_K_r11_39 ) , .Q( u2_uk_K_r12_39 ) );
  DFF_X1 u2_uk_K_r12_reg_4 (.CK( clk ) , .D( u2_uk_K_r11_4 ) , .Q( u2_uk_K_r12_4 ) , .QN( u2_uk_n1772 ) );
  DFF_X1 u2_uk_K_r12_reg_40 (.CK( clk ) , .D( u2_uk_K_r11_40 ) , .Q( u2_uk_K_r12_40 ) , .QN( u2_uk_n1801 ) );
  DFF_X1 u2_uk_K_r12_reg_41 (.CK( clk ) , .D( u2_uk_K_r11_41 ) , .Q( u2_uk_K_r12_41 ) );
  DFF_X1 u2_uk_K_r12_reg_42 (.CK( clk ) , .D( u2_uk_K_r11_42 ) , .Q( u2_uk_K_r12_42 ) );
  DFF_X1 u2_uk_K_r12_reg_43 (.CK( clk ) , .D( u2_uk_K_r11_43 ) , .Q( u2_uk_K_r12_43 ) , .QN( u2_uk_n1802 ) );
  DFF_X1 u2_uk_K_r12_reg_44 (.CK( clk ) , .D( u2_uk_K_r11_44 ) , .Q( u2_uk_K_r12_44 ) );
  DFF_X1 u2_uk_K_r12_reg_45 (.CK( clk ) , .D( u2_uk_K_r11_45 ) , .Q( u2_uk_K_r12_45 ) , .QN( u2_uk_n1803 ) );
  DFF_X1 u2_uk_K_r12_reg_46 (.CK( clk ) , .D( u2_uk_K_r11_46 ) , .Q( u2_uk_K_r12_46 ) , .QN( u2_uk_n1804 ) );
  DFF_X1 u2_uk_K_r12_reg_47 (.CK( clk ) , .D( u2_uk_K_r11_47 ) , .Q( u2_uk_K_r12_47 ) );
  DFF_X1 u2_uk_K_r12_reg_48 (.CK( clk ) , .D( u2_uk_K_r11_48 ) , .Q( u2_uk_K_r12_48 ) , .QN( u2_uk_n1805 ) );
  DFF_X1 u2_uk_K_r12_reg_49 (.CK( clk ) , .D( u2_uk_K_r11_49 ) , .Q( u2_uk_K_r12_49 ) , .QN( u2_uk_n1806 ) );
  DFF_X1 u2_uk_K_r12_reg_5 (.CK( clk ) , .D( u2_uk_K_r11_5 ) , .Q( u2_uk_K_r12_5 ) , .QN( u2_uk_n1773 ) );
  DFF_X1 u2_uk_K_r12_reg_50 (.CK( clk ) , .D( u2_uk_K_r11_50 ) , .Q( u2_uk_K_r12_50 ) , .QN( u2_uk_n1807 ) );
  DFF_X1 u2_uk_K_r12_reg_51 (.CK( clk ) , .D( u2_uk_K_r11_51 ) , .Q( u2_uk_K_r12_51 ) , .QN( u2_uk_n1808 ) );
  DFF_X1 u2_uk_K_r12_reg_52 (.CK( clk ) , .D( u2_uk_K_r11_52 ) , .Q( u2_uk_K_r12_52 ) , .QN( u2_uk_n1809 ) );
  DFF_X1 u2_uk_K_r12_reg_53 (.CK( clk ) , .D( u2_uk_K_r11_53 ) , .Q( u2_uk_K_r12_53 ) , .QN( u2_uk_n1810 ) );
  DFF_X1 u2_uk_K_r12_reg_54 (.CK( clk ) , .D( u2_uk_K_r11_54 ) , .Q( u2_uk_K_r12_54 ) , .QN( u2_uk_n1811 ) );
  DFF_X1 u2_uk_K_r12_reg_55 (.CK( clk ) , .D( u2_uk_K_r11_55 ) , .Q( u2_uk_K_r12_55 ) , .QN( u2_uk_n1812 ) );
  DFF_X1 u2_uk_K_r12_reg_6 (.CK( clk ) , .D( u2_uk_K_r11_6 ) , .Q( u2_uk_K_r12_6 ) , .QN( u2_uk_n1774 ) );
  DFF_X1 u2_uk_K_r12_reg_7 (.CK( clk ) , .D( u2_uk_K_r11_7 ) , .Q( u2_uk_K_r12_7 ) );
  DFF_X1 u2_uk_K_r12_reg_8 (.CK( clk ) , .D( u2_uk_K_r11_8 ) , .Q( u2_uk_K_r12_8 ) , .QN( u2_uk_n1776 ) );
  DFF_X1 u2_uk_K_r12_reg_9 (.CK( clk ) , .D( u2_uk_K_r11_9 ) , .Q( u2_uk_K_r12_9 ) , .QN( u2_uk_n1777 ) );
  DFF_X1 u2_uk_K_r13_reg_0 (.CK( clk ) , .D( u2_uk_K_r12_0 ) , .Q( u2_uk_K_r13_0 ) , .QN( u2_uk_n1813 ) );
  DFF_X1 u2_uk_K_r13_reg_1 (.CK( clk ) , .D( u2_uk_K_r12_1 ) , .Q( u2_uk_K_r13_1 ) );
  DFF_X1 u2_uk_K_r13_reg_10 (.CK( clk ) , .D( u2_uk_K_r12_10 ) , .Q( u2_uk_K_r13_10 ) , .QN( u2_uk_n1820 ) );
  DFF_X1 u2_uk_K_r13_reg_11 (.CK( clk ) , .D( u2_uk_K_r12_11 ) , .Q( u2_uk_K_r13_11 ) , .QN( u2_uk_n1821 ) );
  DFF_X1 u2_uk_K_r13_reg_12 (.CK( clk ) , .D( u2_uk_K_r12_12 ) , .Q( u2_uk_K_r13_12 ) , .QN( u2_uk_n1822 ) );
  DFF_X1 u2_uk_K_r13_reg_13 (.CK( clk ) , .D( u2_uk_K_r12_13 ) , .Q( u2_uk_K_r13_13 ) , .QN( u2_uk_n1823 ) );
  DFF_X1 u2_uk_K_r13_reg_14 (.CK( clk ) , .D( u2_uk_K_r12_14 ) , .Q( u2_uk_K_r13_14 ) , .QN( u2_uk_n1824 ) );
  DFF_X1 u2_uk_K_r13_reg_15 (.CK( clk ) , .D( u2_uk_K_r12_15 ) , .Q( u2_uk_K_r13_15 ) , .QN( u2_uk_n1825 ) );
  DFF_X1 u2_uk_K_r13_reg_16 (.CK( clk ) , .D( u2_uk_K_r12_16 ) , .Q( u2_uk_K_r13_16 ) , .QN( u2_uk_n1826 ) );
  DFF_X1 u2_uk_K_r13_reg_17 (.CK( clk ) , .D( u2_uk_K_r12_17 ) , .Q( u2_uk_K_r13_17 ) );
  DFF_X1 u2_uk_K_r13_reg_18 (.CK( clk ) , .D( u2_uk_K_r12_18 ) , .Q( u2_uk_K_r13_18 ) , .QN( u2_uk_n1828 ) );
  DFF_X1 u2_uk_K_r13_reg_19 (.CK( clk ) , .D( u2_uk_K_r12_19 ) , .Q( u2_uk_K_r13_19 ) );
  DFF_X1 u2_uk_K_r13_reg_2 (.CK( clk ) , .D( u2_uk_K_r12_2 ) , .Q( u2_uk_K_r13_2 ) );
  DFF_X1 u2_uk_K_r13_reg_20 (.CK( clk ) , .D( u2_uk_K_r12_20 ) , .Q( u2_uk_K_r13_20 ) , .QN( u2_uk_n1829 ) );
  DFF_X1 u2_uk_K_r13_reg_21 (.CK( clk ) , .D( u2_uk_K_r12_21 ) , .Q( u2_uk_K_r13_21 ) , .QN( u2_uk_n1830 ) );
  DFF_X1 u2_uk_K_r13_reg_22 (.CK( clk ) , .D( u2_uk_K_r12_22 ) , .Q( u2_uk_K_r13_22 ) );
  DFF_X1 u2_uk_K_r13_reg_23 (.CK( clk ) , .D( u2_uk_K_r12_23 ) , .Q( u2_uk_K_r13_23 ) );
  DFF_X1 u2_uk_K_r13_reg_24 (.CK( clk ) , .D( u2_uk_K_r12_24 ) , .Q( u2_uk_K_r13_24 ) , .QN( u2_uk_n1832 ) );
  DFF_X1 u2_uk_K_r13_reg_25 (.CK( clk ) , .D( u2_uk_K_r12_25 ) , .Q( u2_uk_K_r13_25 ) );
  DFF_X1 u2_uk_K_r13_reg_26 (.CK( clk ) , .D( u2_uk_K_r12_26 ) , .Q( u2_uk_K_r13_26 ) , .QN( u2_uk_n1833 ) );
  DFF_X1 u2_uk_K_r13_reg_27 (.CK( clk ) , .D( u2_uk_K_r12_27 ) , .Q( u2_uk_K_r13_27 ) , .QN( u2_uk_n1834 ) );
  DFF_X1 u2_uk_K_r13_reg_28 (.CK( clk ) , .D( u2_uk_K_r12_28 ) , .Q( u2_uk_K_r13_28 ) , .QN( u2_uk_n1835 ) );
  DFF_X1 u2_uk_K_r13_reg_29 (.CK( clk ) , .D( u2_uk_K_r12_29 ) , .Q( u2_uk_K_r13_29 ) , .QN( u2_uk_n1836 ) );
  DFF_X1 u2_uk_K_r13_reg_3 (.CK( clk ) , .D( u2_uk_K_r12_3 ) , .Q( u2_uk_K_r13_3 ) , .QN( u2_uk_n1814 ) );
  DFF_X1 u2_uk_K_r13_reg_30 (.CK( clk ) , .D( u2_uk_K_r12_30 ) , .Q( u2_uk_K_r13_30 ) , .QN( u2_uk_n1837 ) );
  DFF_X1 u2_uk_K_r13_reg_31 (.CK( clk ) , .D( u2_uk_K_r12_31 ) , .Q( u2_uk_K_r13_31 ) );
  DFF_X1 u2_uk_K_r13_reg_32 (.CK( clk ) , .D( u2_uk_K_r12_32 ) , .Q( u2_uk_K_r13_32 ) );
  DFF_X1 u2_uk_K_r13_reg_33 (.CK( clk ) , .D( u2_uk_K_r12_33 ) , .Q( u2_uk_K_r13_33 ) , .QN( u2_uk_n1838 ) );
  DFF_X1 u2_uk_K_r13_reg_34 (.CK( clk ) , .D( u2_uk_K_r12_34 ) , .Q( u2_uk_K_r13_34 ) , .QN( u2_uk_n1839 ) );
  DFF_X1 u2_uk_K_r13_reg_35 (.CK( clk ) , .D( u2_uk_K_r12_35 ) , .Q( u2_uk_K_r13_35 ) );
  DFF_X1 u2_uk_K_r13_reg_36 (.CK( clk ) , .D( u2_uk_K_r12_36 ) , .Q( u2_uk_K_r13_36 ) );
  DFF_X1 u2_uk_K_r13_reg_37 (.CK( clk ) , .D( u2_uk_K_r12_37 ) , .Q( u2_uk_K_r13_37 ) , .QN( u2_uk_n1840 ) );
  DFF_X1 u2_uk_K_r13_reg_38 (.CK( clk ) , .D( u2_uk_K_r12_38 ) , .Q( u2_uk_K_r13_38 ) );
  DFF_X1 u2_uk_K_r13_reg_39 (.CK( clk ) , .D( u2_uk_K_r12_39 ) , .Q( u2_uk_K_r13_39 ) , .QN( u2_uk_n1842 ) );
  DFF_X1 u2_uk_K_r13_reg_4 (.CK( clk ) , .D( u2_uk_K_r12_4 ) , .Q( u2_uk_K_r13_4 ) );
  DFF_X1 u2_uk_K_r13_reg_40 (.CK( clk ) , .D( u2_uk_K_r12_40 ) , .Q( u2_uk_K_r13_40 ) , .QN( u2_uk_n1843 ) );
  DFF_X1 u2_uk_K_r13_reg_41 (.CK( clk ) , .D( u2_uk_K_r12_41 ) , .Q( u2_uk_K_r13_41 ) , .QN( u2_uk_n1844 ) );
  DFF_X1 u2_uk_K_r13_reg_42 (.CK( clk ) , .D( u2_uk_K_r12_42 ) , .Q( u2_uk_K_r13_42 ) , .QN( u2_uk_n1845 ) );
  DFF_X1 u2_uk_K_r13_reg_43 (.CK( clk ) , .D( u2_uk_K_r12_43 ) , .Q( u2_uk_K_r13_43 ) , .QN( u2_uk_n1846 ) );
  DFF_X1 u2_uk_K_r13_reg_44 (.CK( clk ) , .D( u2_uk_K_r12_44 ) , .Q( u2_uk_K_r13_44 ) );
  DFF_X1 u2_uk_K_r13_reg_45 (.CK( clk ) , .D( u2_uk_K_r12_45 ) , .Q( u2_uk_K_r13_45 ) , .QN( u2_uk_n1849 ) );
  DFF_X1 u2_uk_K_r13_reg_46 (.CK( clk ) , .D( u2_uk_K_r12_46 ) , .Q( u2_uk_K_r13_46 ) , .QN( u2_uk_n1850 ) );
  DFF_X1 u2_uk_K_r13_reg_47 (.CK( clk ) , .D( u2_uk_K_r12_47 ) , .Q( u2_uk_K_r13_47 ) , .QN( u2_uk_n1851 ) );
  DFF_X1 u2_uk_K_r13_reg_48 (.CK( clk ) , .D( u2_uk_K_r12_48 ) , .Q( u2_uk_K_r13_48 ) , .QN( u2_uk_n1852 ) );
  DFF_X1 u2_uk_K_r13_reg_49 (.CK( clk ) , .D( u2_uk_K_r12_49 ) , .Q( u2_uk_K_r13_49 ) , .QN( u2_uk_n1853 ) );
  DFF_X1 u2_uk_K_r13_reg_5 (.CK( clk ) , .D( u2_uk_K_r12_5 ) , .Q( u2_uk_K_r13_5 ) , .QN( u2_uk_n1815 ) );
  DFF_X1 u2_uk_K_r13_reg_50 (.CK( clk ) , .D( u2_uk_K_r12_50 ) , .Q( u2_uk_K_r13_50 ) , .QN( u2_uk_n1854 ) );
  DFF_X1 u2_uk_K_r13_reg_51 (.CK( clk ) , .D( u2_uk_K_r12_51 ) , .Q( u2_uk_K_r13_51 ) , .QN( u2_uk_n1855 ) );
  DFF_X1 u2_uk_K_r13_reg_52 (.CK( clk ) , .D( u2_uk_K_r12_52 ) , .Q( u2_uk_K_r13_52 ) , .QN( u2_uk_n1856 ) );
  DFF_X1 u2_uk_K_r13_reg_53 (.CK( clk ) , .D( u2_uk_K_r12_53 ) , .Q( u2_uk_K_r13_53 ) );
  DFF_X1 u2_uk_K_r13_reg_54 (.CK( clk ) , .D( u2_uk_K_r12_54 ) , .Q( u2_uk_K_r13_54 ) , .QN( u2_uk_n1857 ) );
  DFF_X1 u2_uk_K_r13_reg_55 (.CK( clk ) , .D( u2_uk_K_r12_55 ) , .Q( u2_uk_K_r13_55 ) );
  DFF_X1 u2_uk_K_r13_reg_6 (.CK( clk ) , .D( u2_uk_K_r12_6 ) , .Q( u2_uk_K_r13_6 ) , .QN( u2_uk_n1816 ) );
  DFF_X1 u2_uk_K_r13_reg_7 (.CK( clk ) , .D( u2_uk_K_r12_7 ) , .Q( u2_uk_K_r13_7 ) , .QN( u2_uk_n1817 ) );
  DFF_X1 u2_uk_K_r13_reg_8 (.CK( clk ) , .D( u2_uk_K_r12_8 ) , .Q( u2_uk_K_r13_8 ) , .QN( u2_uk_n1818 ) );
  DFF_X1 u2_uk_K_r13_reg_9 (.CK( clk ) , .D( u2_uk_K_r12_9 ) , .Q( u2_uk_K_r13_9 ) , .QN( u2_uk_n1819 ) );
  DFF_X1 u2_uk_K_r14_reg_0 (.CK( clk ) , .D( u2_uk_K_r13_0 ) , .QN( u2_uk_n1188 ) );
  DFF_X1 u2_uk_K_r14_reg_1 (.CK( clk ) , .D( u2_uk_K_r13_1 ) , .QN( u2_uk_n1189 ) );
  DFF_X1 u2_uk_K_r14_reg_10 (.CK( clk ) , .D( u2_uk_K_r13_10 ) , .Q( u2_uk_K_r14_10 ) );
  DFF_X1 u2_uk_K_r14_reg_11 (.CK( clk ) , .D( u2_uk_K_r13_11 ) , .Q( u2_uk_K_r14_11 ) );
  DFF_X1 u2_uk_K_r14_reg_12 (.CK( clk ) , .D( u2_uk_K_r13_12 ) , .Q( u2_uk_K_r14_12 ) );
  DFF_X1 u2_uk_K_r14_reg_13 (.CK( clk ) , .D( u2_uk_K_r13_13 ) , .QN( u2_uk_n1194 ) );
  DFF_X1 u2_uk_K_r14_reg_14 (.CK( clk ) , .D( u2_uk_K_r13_14 ) , .QN( u2_uk_n1195 ) );
  DFF_X1 u2_uk_K_r14_reg_15 (.CK( clk ) , .D( u2_uk_K_r13_15 ) , .Q( u2_uk_K_r14_15 ) );
  DFF_X1 u2_uk_K_r14_reg_16 (.CK( clk ) , .D( u2_uk_K_r13_16 ) , .Q( u2_uk_K_r14_16 ) );
  DFF_X1 u2_uk_K_r14_reg_17 (.CK( clk ) , .D( u2_uk_K_r13_17 ) , .QN( u2_uk_n1197 ) );
  DFF_X1 u2_uk_K_r14_reg_18 (.CK( clk ) , .D( u2_uk_K_r13_18 ) , .Q( u2_uk_K_r14_18 ) );
  DFF_X1 u2_uk_K_r14_reg_19 (.CK( clk ) , .D( u2_uk_K_r13_19 ) , .QN( u2_uk_n1198 ) );
  DFF_X1 u2_uk_K_r14_reg_2 (.CK( clk ) , .D( u2_uk_K_r13_2 ) , .Q( u2_uk_K_r14_2 ) );
  DFF_X1 u2_uk_K_r14_reg_20 (.CK( clk ) , .D( u2_uk_K_r13_20 ) , .QN( u2_uk_n1199 ) );
  DFF_X1 u2_uk_K_r14_reg_21 (.CK( clk ) , .D( u2_uk_K_r13_21 ) , .QN( u2_uk_n1200 ) );
  DFF_X1 u2_uk_K_r14_reg_22 (.CK( clk ) , .D( u2_uk_K_r13_22 ) , .QN( u2_uk_n1201 ) );
  DFF_X1 u2_uk_K_r14_reg_23 (.CK( clk ) , .D( u2_uk_K_r13_23 ) , .Q( u2_uk_K_r14_23 ) , .QN( u2_uk_n1203 ) );
  DFF_X1 u2_uk_K_r14_reg_24 (.CK( clk ) , .D( u2_uk_K_r13_24 ) , .QN( u2_uk_n1204 ) );
  DFF_X1 u2_uk_K_r14_reg_25 (.CK( clk ) , .D( u2_uk_K_r13_25 ) , .QN( u2_uk_n1205 ) );
  DFF_X1 u2_uk_K_r14_reg_26 (.CK( clk ) , .D( u2_uk_K_r13_26 ) , .QN( u2_uk_n1206 ) );
  DFF_X1 u2_uk_K_r14_reg_27 (.CK( clk ) , .D( u2_uk_K_r13_27 ) , .QN( u2_uk_n1207 ) );
  DFF_X1 u2_uk_K_r14_reg_28 (.CK( clk ) , .D( u2_uk_K_r13_28 ) , .QN( u2_uk_n1208 ) );
  DFF_X1 u2_uk_K_r14_reg_29 (.CK( clk ) , .D( u2_uk_K_r13_29 ) , .QN( u2_uk_n1209 ) );
  DFF_X1 u2_uk_K_r14_reg_3 (.CK( clk ) , .D( u2_uk_K_r13_3 ) , .Q( u2_uk_K_r14_3 ) );
  DFF_X1 u2_uk_K_r14_reg_30 (.CK( clk ) , .D( u2_uk_K_r13_30 ) , .QN( u2_uk_n1210 ) );
  DFF_X1 u2_uk_K_r14_reg_31 (.CK( clk ) , .D( u2_uk_K_r13_31 ) , .QN( u2_uk_n1211 ) );
  DFF_X1 u2_uk_K_r14_reg_32 (.CK( clk ) , .D( u2_uk_K_r13_32 ) , .QN( u2_uk_n1212 ) );
  DFF_X1 u2_uk_K_r14_reg_33 (.CK( clk ) , .D( u2_uk_K_r13_33 ) , .QN( u2_uk_n1213 ) );
  DFF_X1 u2_uk_K_r14_reg_34 (.CK( clk ) , .D( u2_uk_K_r13_34 ) , .QN( u2_uk_n1214 ) );
  DFF_X1 u2_uk_K_r14_reg_35 (.CK( clk ) , .D( u2_uk_K_r13_35 ) , .QN( u2_uk_n1215 ) );
  DFF_X1 u2_uk_K_r14_reg_36 (.CK( clk ) , .D( u2_uk_K_r13_36 ) , .QN( u2_uk_n1216 ) );
  DFF_X1 u2_uk_K_r14_reg_37 (.CK( clk ) , .D( u2_uk_K_r13_37 ) , .QN( u2_uk_n1217 ) );
  DFF_X1 u2_uk_K_r14_reg_38 (.CK( clk ) , .D( u2_uk_K_r13_38 ) , .Q( u2_uk_K_r14_38 ) );
  DFF_X1 u2_uk_K_r14_reg_39 (.CK( clk ) , .D( u2_uk_K_r13_39 ) , .Q( u2_uk_K_r14_39 ) );
  DFF_X1 u2_uk_K_r14_reg_4 (.CK( clk ) , .D( u2_uk_K_r13_4 ) , .QN( u2_uk_n1190 ) );
  DFF_X1 u2_uk_K_r14_reg_40 (.CK( clk ) , .D( u2_uk_K_r13_40 ) , .QN( u2_uk_n1218 ) );
  DFF_X1 u2_uk_K_r14_reg_41 (.CK( clk ) , .D( u2_uk_K_r13_41 ) , .QN( u2_uk_n1219 ) );
  DFF_X1 u2_uk_K_r14_reg_42 (.CK( clk ) , .D( u2_uk_K_r13_42 ) , .Q( u2_uk_K_r14_42 ) );
  DFF_X1 u2_uk_K_r14_reg_43 (.CK( clk ) , .D( u2_uk_K_r13_43 ) , .Q( u2_uk_K_r14_43 ) );
  DFF_X1 u2_uk_K_r14_reg_44 (.CK( clk ) , .D( u2_uk_K_r13_44 ) , .QN( u2_uk_n1220 ) );
  DFF_X1 u2_uk_K_r14_reg_45 (.CK( clk ) , .D( u2_uk_K_r13_45 ) , .Q( u2_uk_K_r14_45 ) );
  DFF_X1 u2_uk_K_r14_reg_46 (.CK( clk ) , .D( u2_uk_K_r13_46 ) , .Q( u2_uk_K_r14_46 ) );
  DFF_X1 u2_uk_K_r14_reg_47 (.CK( clk ) , .D( u2_uk_K_r13_47 ) , .QN( u2_uk_n1221 ) );
  DFF_X1 u2_uk_K_r14_reg_48 (.CK( clk ) , .D( u2_uk_K_r13_48 ) , .QN( u2_uk_n1222 ) );
  DFF_X1 u2_uk_K_r14_reg_49 (.CK( clk ) , .D( u2_uk_K_r13_49 ) , .QN( u2_uk_n1223 ) );
  DFF_X1 u2_uk_K_r14_reg_5 (.CK( clk ) , .D( u2_uk_K_r13_5 ) , .Q( u2_uk_K_r14_5 ) );
  DFF_X1 u2_uk_K_r14_reg_50 (.CK( clk ) , .D( u2_uk_K_r13_50 ) , .Q( u2_uk_K_r14_50 ) );
  DFF_X1 u2_uk_K_r14_reg_51 (.CK( clk ) , .D( u2_uk_K_r13_51 ) , .QN( u2_uk_n1225 ) );
  DFF_X1 u2_uk_K_r14_reg_52 (.CK( clk ) , .D( u2_uk_K_r13_52 ) , .QN( u2_uk_n1226 ) );
  DFF_X1 u2_uk_K_r14_reg_53 (.CK( clk ) , .D( u2_uk_K_r13_53 ) , .QN( u2_uk_n1227 ) );
  DFF_X1 u2_uk_K_r14_reg_54 (.CK( clk ) , .D( u2_uk_K_r13_54 ) , .QN( u2_uk_n1228 ) );
  DFF_X1 u2_uk_K_r14_reg_55 (.CK( clk ) , .D( u2_uk_K_r13_55 ) , .QN( u2_uk_n1229 ) );
  DFF_X1 u2_uk_K_r14_reg_6 (.CK( clk ) , .D( u2_uk_K_r13_6 ) , .QN( u2_uk_n1191 ) );
  DFF_X1 u2_uk_K_r14_reg_7 (.CK( clk ) , .D( u2_uk_K_r13_7 ) , .QN( u2_uk_n1192 ) );
  DFF_X1 u2_uk_K_r14_reg_8 (.CK( clk ) , .D( u2_uk_K_r13_8 ) , .Q( u2_uk_K_r14_8 ) );
  DFF_X1 u2_uk_K_r14_reg_9 (.CK( clk ) , .D( u2_uk_K_r13_9 ) , .Q( u2_uk_K_r14_9 ) );
  DFF_X1 u2_uk_K_r1_reg_0 (.CK( clk ) , .D( u2_uk_K_r0_0 ) , .Q( u2_uk_K_r1_0 ) , .QN( u2_uk_n1277 ) );
  DFF_X1 u2_uk_K_r1_reg_1 (.CK( clk ) , .D( u2_uk_K_r0_1 ) , .Q( u2_uk_K_r1_1 ) , .QN( u2_uk_n1278 ) );
  DFF_X1 u2_uk_K_r1_reg_10 (.CK( clk ) , .D( u2_uk_K_r0_10 ) , .Q( u2_uk_K_r1_10 ) );
  DFF_X1 u2_uk_K_r1_reg_11 (.CK( clk ) , .D( u2_uk_K_r0_11 ) , .Q( u2_uk_K_r1_11 ) , .QN( u2_uk_n1285 ) );
  DFF_X1 u2_uk_K_r1_reg_12 (.CK( clk ) , .D( u2_uk_K_r0_12 ) , .Q( u2_uk_K_r1_12 ) , .QN( u2_uk_n1286 ) );
  DFF_X1 u2_uk_K_r1_reg_13 (.CK( clk ) , .D( u2_uk_K_r0_13 ) , .Q( u2_uk_K_r1_13 ) , .QN( u2_uk_n1287 ) );
  DFF_X1 u2_uk_K_r1_reg_14 (.CK( clk ) , .D( u2_uk_K_r0_14 ) , .Q( u2_uk_K_r1_14 ) , .QN( u2_uk_n1288 ) );
  DFF_X1 u2_uk_K_r1_reg_15 (.CK( clk ) , .D( u2_uk_K_r0_15 ) , .Q( u2_uk_K_r1_15 ) );
  DFF_X1 u2_uk_K_r1_reg_16 (.CK( clk ) , .D( u2_uk_K_r0_16 ) , .Q( u2_uk_K_r1_16 ) );
  DFF_X1 u2_uk_K_r1_reg_17 (.CK( clk ) , .D( u2_uk_K_r0_17 ) , .Q( u2_uk_K_r1_17 ) , .QN( u2_uk_n1289 ) );
  DFF_X1 u2_uk_K_r1_reg_18 (.CK( clk ) , .D( u2_uk_K_r0_18 ) , .Q( u2_uk_K_r1_18 ) );
  DFF_X1 u2_uk_K_r1_reg_19 (.CK( clk ) , .D( u2_uk_K_r0_19 ) , .Q( u2_uk_K_r1_19 ) , .QN( u2_uk_n1290 ) );
  DFF_X1 u2_uk_K_r1_reg_2 (.CK( clk ) , .D( u2_uk_K_r0_2 ) , .Q( u2_uk_K_r1_2 ) , .QN( u2_uk_n1279 ) );
  DFF_X1 u2_uk_K_r1_reg_20 (.CK( clk ) , .D( u2_uk_K_r0_20 ) , .Q( u2_uk_K_r1_20 ) , .QN( u2_uk_n1291 ) );
  DFF_X1 u2_uk_K_r1_reg_21 (.CK( clk ) , .D( u2_uk_K_r0_21 ) , .Q( u2_uk_K_r1_21 ) );
  DFF_X1 u2_uk_K_r1_reg_22 (.CK( clk ) , .D( u2_uk_K_r0_22 ) , .Q( u2_uk_K_r1_22 ) );
  DFF_X1 u2_uk_K_r1_reg_23 (.CK( clk ) , .D( u2_uk_K_r0_23 ) , .Q( u2_uk_K_r1_23 ) , .QN( u2_uk_n1292 ) );
  DFF_X1 u2_uk_K_r1_reg_24 (.CK( clk ) , .D( u2_uk_K_r0_24 ) , .Q( u2_uk_K_r1_24 ) , .QN( u2_uk_n1293 ) );
  DFF_X1 u2_uk_K_r1_reg_25 (.CK( clk ) , .D( u2_uk_K_r0_25 ) , .Q( u2_uk_K_r1_25 ) , .QN( u2_uk_n1294 ) );
  DFF_X1 u2_uk_K_r1_reg_26 (.CK( clk ) , .D( u2_uk_K_r0_26 ) , .Q( u2_uk_K_r1_26 ) , .QN( u2_uk_n1295 ) );
  DFF_X1 u2_uk_K_r1_reg_27 (.CK( clk ) , .D( u2_uk_K_r0_27 ) , .Q( u2_uk_K_r1_27 ) , .QN( u2_uk_n1296 ) );
  DFF_X1 u2_uk_K_r1_reg_28 (.CK( clk ) , .D( u2_uk_K_r0_28 ) , .Q( u2_uk_K_r1_28 ) , .QN( u2_uk_n1297 ) );
  DFF_X1 u2_uk_K_r1_reg_29 (.CK( clk ) , .D( u2_uk_K_r0_29 ) , .Q( u2_uk_K_r1_29 ) , .QN( u2_uk_n1298 ) );
  DFF_X1 u2_uk_K_r1_reg_3 (.CK( clk ) , .D( u2_uk_K_r0_3 ) , .Q( u2_uk_K_r1_3 ) , .QN( u2_uk_n1280 ) );
  DFF_X1 u2_uk_K_r1_reg_30 (.CK( clk ) , .D( u2_uk_K_r0_30 ) , .Q( u2_uk_K_r1_30 ) , .QN( u2_uk_n1299 ) );
  DFF_X1 u2_uk_K_r1_reg_31 (.CK( clk ) , .D( u2_uk_K_r0_31 ) , .Q( u2_uk_K_r1_31 ) , .QN( u2_uk_n1300 ) );
  DFF_X1 u2_uk_K_r1_reg_32 (.CK( clk ) , .D( u2_uk_K_r0_32 ) , .Q( u2_uk_K_r1_32 ) , .QN( u2_uk_n1301 ) );
  DFF_X1 u2_uk_K_r1_reg_33 (.CK( clk ) , .D( u2_uk_K_r0_33 ) , .Q( u2_uk_K_r1_33 ) );
  DFF_X1 u2_uk_K_r1_reg_34 (.CK( clk ) , .D( u2_uk_K_r0_34 ) , .Q( u2_uk_K_r1_34 ) , .QN( u2_uk_n1302 ) );
  DFF_X1 u2_uk_K_r1_reg_35 (.CK( clk ) , .D( u2_uk_K_r0_35 ) , .Q( u2_uk_K_r1_35 ) , .QN( u2_uk_n1303 ) );
  DFF_X1 u2_uk_K_r1_reg_36 (.CK( clk ) , .D( u2_uk_K_r0_36 ) , .Q( u2_uk_K_r1_36 ) );
  DFF_X1 u2_uk_K_r1_reg_37 (.CK( clk ) , .D( u2_uk_K_r0_37 ) , .Q( u2_uk_K_r1_37 ) , .QN( u2_uk_n1304 ) );
  DFF_X1 u2_uk_K_r1_reg_38 (.CK( clk ) , .D( u2_uk_K_r0_38 ) , .Q( u2_uk_K_r1_38 ) , .QN( u2_uk_n1305 ) );
  DFF_X1 u2_uk_K_r1_reg_39 (.CK( clk ) , .D( u2_uk_K_r0_39 ) , .Q( u2_uk_K_r1_39 ) );
  DFF_X1 u2_uk_K_r1_reg_4 (.CK( clk ) , .D( u2_uk_K_r0_4 ) , .Q( u2_uk_K_r1_4 ) , .QN( u2_uk_n1281 ) );
  DFF_X1 u2_uk_K_r1_reg_40 (.CK( clk ) , .D( u2_uk_K_r0_40 ) , .Q( u2_uk_K_r1_40 ) , .QN( u2_uk_n1306 ) );
  DFF_X1 u2_uk_K_r1_reg_41 (.CK( clk ) , .D( u2_uk_K_r0_41 ) , .Q( u2_uk_K_r1_41 ) );
  DFF_X1 u2_uk_K_r1_reg_42 (.CK( clk ) , .D( u2_uk_K_r0_42 ) , .Q( u2_uk_K_r1_42 ) );
  DFF_X1 u2_uk_K_r1_reg_43 (.CK( clk ) , .D( u2_uk_K_r0_43 ) , .Q( u2_uk_K_r1_43 ) , .QN( u2_uk_n1308 ) );
  DFF_X1 u2_uk_K_r1_reg_44 (.CK( clk ) , .D( u2_uk_K_r0_44 ) , .Q( u2_uk_K_r1_44 ) );
  DFF_X1 u2_uk_K_r1_reg_45 (.CK( clk ) , .D( u2_uk_K_r0_45 ) , .Q( u2_uk_K_r1_45 ) , .QN( u2_uk_n1309 ) );
  DFF_X1 u2_uk_K_r1_reg_46 (.CK( clk ) , .D( u2_uk_K_r0_46 ) , .Q( u2_uk_K_r1_46 ) , .QN( u2_uk_n1310 ) );
  DFF_X1 u2_uk_K_r1_reg_47 (.CK( clk ) , .D( u2_uk_K_r0_47 ) , .Q( u2_uk_K_r1_47 ) );
  DFF_X1 u2_uk_K_r1_reg_48 (.CK( clk ) , .D( u2_uk_K_r0_48 ) , .Q( u2_uk_K_r1_48 ) , .QN( u2_uk_n1311 ) );
  DFF_X1 u2_uk_K_r1_reg_49 (.CK( clk ) , .D( u2_uk_K_r0_49 ) , .Q( u2_uk_K_r1_49 ) , .QN( u2_uk_n1312 ) );
  DFF_X1 u2_uk_K_r1_reg_5 (.CK( clk ) , .D( u2_uk_K_r0_5 ) , .Q( u2_uk_K_r1_5 ) , .QN( u2_uk_n1282 ) );
  DFF_X1 u2_uk_K_r1_reg_50 (.CK( clk ) , .D( u2_uk_K_r0_50 ) , .Q( u2_uk_K_r1_50 ) , .QN( u2_uk_n1313 ) );
  DFF_X1 u2_uk_K_r1_reg_51 (.CK( clk ) , .D( u2_uk_K_r0_51 ) , .Q( u2_uk_K_r1_51 ) , .QN( u2_uk_n1314 ) );
  DFF_X1 u2_uk_K_r1_reg_52 (.CK( clk ) , .D( u2_uk_K_r0_52 ) , .Q( u2_uk_K_r1_52 ) , .QN( u2_uk_n1315 ) );
  DFF_X1 u2_uk_K_r1_reg_53 (.CK( clk ) , .D( u2_uk_K_r0_53 ) , .Q( u2_uk_K_r1_53 ) , .QN( u2_uk_n1316 ) );
  DFF_X1 u2_uk_K_r1_reg_54 (.CK( clk ) , .D( u2_uk_K_r0_54 ) , .Q( u2_uk_K_r1_54 ) , .QN( u2_uk_n1317 ) );
  DFF_X1 u2_uk_K_r1_reg_55 (.CK( clk ) , .D( u2_uk_K_r0_55 ) , .Q( u2_uk_K_r1_55 ) , .QN( u2_uk_n1318 ) );
  DFF_X1 u2_uk_K_r1_reg_6 (.CK( clk ) , .D( u2_uk_K_r0_6 ) , .Q( u2_uk_K_r1_6 ) );
  DFF_X1 u2_uk_K_r1_reg_7 (.CK( clk ) , .D( u2_uk_K_r0_7 ) , .Q( u2_uk_K_r1_7 ) );
  DFF_X1 u2_uk_K_r1_reg_8 (.CK( clk ) , .D( u2_uk_K_r0_8 ) , .Q( u2_uk_K_r1_8 ) , .QN( u2_uk_n1283 ) );
  DFF_X1 u2_uk_K_r1_reg_9 (.CK( clk ) , .D( u2_uk_K_r0_9 ) , .Q( u2_uk_K_r1_9 ) , .QN( u2_uk_n1284 ) );
  DFF_X1 u2_uk_K_r2_reg_0 (.CK( clk ) , .D( u2_uk_K_r1_0 ) , .Q( u2_uk_K_r2_0 ) , .QN( u2_uk_n1319 ) );
  DFF_X1 u2_uk_K_r2_reg_1 (.CK( clk ) , .D( u2_uk_K_r1_1 ) , .Q( u2_uk_K_r2_1 ) , .QN( u2_uk_n1320 ) );
  DFF_X1 u2_uk_K_r2_reg_10 (.CK( clk ) , .D( u2_uk_K_r1_10 ) , .Q( u2_uk_K_r2_10 ) , .QN( u2_uk_n1327 ) );
  DFF_X1 u2_uk_K_r2_reg_11 (.CK( clk ) , .D( u2_uk_K_r1_11 ) , .Q( u2_uk_K_r2_11 ) , .QN( u2_uk_n1328 ) );
  DFF_X1 u2_uk_K_r2_reg_12 (.CK( clk ) , .D( u2_uk_K_r1_12 ) , .Q( u2_uk_K_r2_12 ) , .QN( u2_uk_n1329 ) );
  DFF_X1 u2_uk_K_r2_reg_13 (.CK( clk ) , .D( u2_uk_K_r1_13 ) , .Q( u2_uk_K_r2_13 ) );
  DFF_X1 u2_uk_K_r2_reg_14 (.CK( clk ) , .D( u2_uk_K_r1_14 ) , .Q( u2_uk_K_r2_14 ) , .QN( u2_uk_n1330 ) );
  DFF_X1 u2_uk_K_r2_reg_15 (.CK( clk ) , .D( u2_uk_K_r1_15 ) , .Q( u2_uk_K_r2_15 ) , .QN( u2_uk_n1331 ) );
  DFF_X1 u2_uk_K_r2_reg_16 (.CK( clk ) , .D( u2_uk_K_r1_16 ) , .Q( u2_uk_K_r2_16 ) );
  DFF_X1 u2_uk_K_r2_reg_17 (.CK( clk ) , .D( u2_uk_K_r1_17 ) , .Q( u2_uk_K_r2_17 ) , .QN( u2_uk_n1333 ) );
  DFF_X1 u2_uk_K_r2_reg_18 (.CK( clk ) , .D( u2_uk_K_r1_18 ) , .Q( u2_uk_K_r2_18 ) );
  DFF_X1 u2_uk_K_r2_reg_19 (.CK( clk ) , .D( u2_uk_K_r1_19 ) , .Q( u2_uk_K_r2_19 ) , .QN( u2_uk_n1335 ) );
  DFF_X1 u2_uk_K_r2_reg_2 (.CK( clk ) , .D( u2_uk_K_r1_2 ) , .Q( u2_uk_K_r2_2 ) , .QN( u2_uk_n1321 ) );
  DFF_X1 u2_uk_K_r2_reg_20 (.CK( clk ) , .D( u2_uk_K_r1_20 ) , .Q( u2_uk_K_r2_20 ) );
  DFF_X1 u2_uk_K_r2_reg_21 (.CK( clk ) , .D( u2_uk_K_r1_21 ) , .Q( u2_uk_K_r2_21 ) );
  DFF_X1 u2_uk_K_r2_reg_22 (.CK( clk ) , .D( u2_uk_K_r1_22 ) , .Q( u2_uk_K_r2_22 ) , .QN( u2_uk_n1336 ) );
  DFF_X1 u2_uk_K_r2_reg_23 (.CK( clk ) , .D( u2_uk_K_r1_23 ) , .Q( u2_uk_K_r2_23 ) , .QN( u2_uk_n1337 ) );
  DFF_X1 u2_uk_K_r2_reg_24 (.CK( clk ) , .D( u2_uk_K_r1_24 ) , .Q( u2_uk_K_r2_24 ) );
  DFF_X1 u2_uk_K_r2_reg_25 (.CK( clk ) , .D( u2_uk_K_r1_25 ) , .Q( u2_uk_K_r2_25 ) );
  DFF_X1 u2_uk_K_r2_reg_26 (.CK( clk ) , .D( u2_uk_K_r1_26 ) , .Q( u2_uk_K_r2_26 ) );
  DFF_X1 u2_uk_K_r2_reg_27 (.CK( clk ) , .D( u2_uk_K_r1_27 ) , .Q( u2_uk_K_r2_27 ) );
  DFF_X1 u2_uk_K_r2_reg_28 (.CK( clk ) , .D( u2_uk_K_r1_28 ) , .Q( u2_uk_K_r2_28 ) );
  DFF_X1 u2_uk_K_r2_reg_29 (.CK( clk ) , .D( u2_uk_K_r1_29 ) , .Q( u2_uk_K_r2_29 ) );
  DFF_X1 u2_uk_K_r2_reg_3 (.CK( clk ) , .D( u2_uk_K_r1_3 ) , .Q( u2_uk_K_r2_3 ) , .QN( u2_uk_n1322 ) );
  DFF_X1 u2_uk_K_r2_reg_30 (.CK( clk ) , .D( u2_uk_K_r1_30 ) , .Q( u2_uk_K_r2_30 ) );
  DFF_X1 u2_uk_K_r2_reg_31 (.CK( clk ) , .D( u2_uk_K_r1_31 ) , .Q( u2_uk_K_r2_31 ) );
  DFF_X1 u2_uk_K_r2_reg_32 (.CK( clk ) , .D( u2_uk_K_r1_32 ) , .Q( u2_uk_K_r2_32 ) , .QN( u2_uk_n1339 ) );
  DFF_X1 u2_uk_K_r2_reg_33 (.CK( clk ) , .D( u2_uk_K_r1_33 ) , .Q( u2_uk_K_r2_33 ) );
  DFF_X1 u2_uk_K_r2_reg_34 (.CK( clk ) , .D( u2_uk_K_r1_34 ) , .Q( u2_uk_K_r2_34 ) , .QN( u2_uk_n1341 ) );
  DFF_X1 u2_uk_K_r2_reg_35 (.CK( clk ) , .D( u2_uk_K_r1_35 ) , .Q( u2_uk_K_r2_35 ) , .QN( u2_uk_n1342 ) );
  DFF_X1 u2_uk_K_r2_reg_36 (.CK( clk ) , .D( u2_uk_K_r1_36 ) , .Q( u2_uk_K_r2_36 ) , .QN( u2_uk_n1344 ) );
  DFF_X1 u2_uk_K_r2_reg_37 (.CK( clk ) , .D( u2_uk_K_r1_37 ) , .Q( u2_uk_K_r2_37 ) , .QN( u2_uk_n1345 ) );
  DFF_X1 u2_uk_K_r2_reg_38 (.CK( clk ) , .D( u2_uk_K_r1_38 ) , .Q( u2_uk_K_r2_38 ) , .QN( u2_uk_n1346 ) );
  DFF_X1 u2_uk_K_r2_reg_39 (.CK( clk ) , .D( u2_uk_K_r1_39 ) , .Q( u2_uk_K_r2_39 ) , .QN( u2_uk_n1347 ) );
  DFF_X1 u2_uk_K_r2_reg_4 (.CK( clk ) , .D( u2_uk_K_r1_4 ) , .Q( u2_uk_K_r2_4 ) );
  DFF_X1 u2_uk_K_r2_reg_40 (.CK( clk ) , .D( u2_uk_K_r1_40 ) , .Q( u2_uk_K_r2_40 ) , .QN( u2_uk_n1348 ) );
  DFF_X1 u2_uk_K_r2_reg_41 (.CK( clk ) , .D( u2_uk_K_r1_41 ) , .Q( u2_uk_K_r2_41 ) );
  DFF_X1 u2_uk_K_r2_reg_42 (.CK( clk ) , .D( u2_uk_K_r1_42 ) , .Q( u2_uk_K_r2_42 ) , .QN( u2_uk_n1350 ) );
  DFF_X1 u2_uk_K_r2_reg_43 (.CK( clk ) , .D( u2_uk_K_r1_43 ) , .Q( u2_uk_K_r2_43 ) , .QN( u2_uk_n1351 ) );
  DFF_X1 u2_uk_K_r2_reg_44 (.CK( clk ) , .D( u2_uk_K_r1_44 ) , .Q( u2_uk_K_r2_44 ) , .QN( u2_uk_n1352 ) );
  DFF_X1 u2_uk_K_r2_reg_45 (.CK( clk ) , .D( u2_uk_K_r1_45 ) , .Q( u2_uk_K_r2_45 ) , .QN( u2_uk_n1353 ) );
  DFF_X1 u2_uk_K_r2_reg_46 (.CK( clk ) , .D( u2_uk_K_r1_46 ) , .Q( u2_uk_K_r2_46 ) );
  DFF_X1 u2_uk_K_r2_reg_47 (.CK( clk ) , .D( u2_uk_K_r1_47 ) , .Q( u2_uk_K_r2_47 ) );
  DFF_X1 u2_uk_K_r2_reg_48 (.CK( clk ) , .D( u2_uk_K_r1_48 ) , .Q( u2_uk_K_r2_48 ) , .QN( u2_uk_n1356 ) );
  DFF_X1 u2_uk_K_r2_reg_49 (.CK( clk ) , .D( u2_uk_K_r1_49 ) , .Q( u2_uk_K_r2_49 ) );
  DFF_X1 u2_uk_K_r2_reg_5 (.CK( clk ) , .D( u2_uk_K_r1_5 ) , .Q( u2_uk_K_r2_5 ) , .QN( u2_uk_n1323 ) );
  DFF_X1 u2_uk_K_r2_reg_50 (.CK( clk ) , .D( u2_uk_K_r1_50 ) , .Q( u2_uk_K_r2_50 ) );
  DFF_X1 u2_uk_K_r2_reg_51 (.CK( clk ) , .D( u2_uk_K_r1_51 ) , .Q( u2_uk_K_r2_51 ) , .QN( u2_uk_n1359 ) );
  DFF_X1 u2_uk_K_r2_reg_52 (.CK( clk ) , .D( u2_uk_K_r1_52 ) , .Q( u2_uk_K_r2_52 ) , .QN( u2_uk_n1360 ) );
  DFF_X1 u2_uk_K_r2_reg_53 (.CK( clk ) , .D( u2_uk_K_r1_53 ) , .Q( u2_uk_K_r2_53 ) );
  DFF_X1 u2_uk_K_r2_reg_54 (.CK( clk ) , .D( u2_uk_K_r1_54 ) , .Q( u2_uk_K_r2_54 ) , .QN( u2_uk_n1361 ) );
  DFF_X1 u2_uk_K_r2_reg_55 (.CK( clk ) , .D( u2_uk_K_r1_55 ) , .Q( u2_uk_K_r2_55 ) , .QN( u2_uk_n1363 ) );
  DFF_X1 u2_uk_K_r2_reg_6 (.CK( clk ) , .D( u2_uk_K_r1_6 ) , .Q( u2_uk_K_r2_6 ) , .QN( u2_uk_n1324 ) );
  DFF_X1 u2_uk_K_r2_reg_7 (.CK( clk ) , .D( u2_uk_K_r1_7 ) , .Q( u2_uk_K_r2_7 ) );
  DFF_X1 u2_uk_K_r2_reg_8 (.CK( clk ) , .D( u2_uk_K_r1_8 ) , .Q( u2_uk_K_r2_8 ) , .QN( u2_uk_n1325 ) );
  DFF_X1 u2_uk_K_r2_reg_9 (.CK( clk ) , .D( u2_uk_K_r1_9 ) , .Q( u2_uk_K_r2_9 ) , .QN( u2_uk_n1326 ) );
  DFF_X1 u2_uk_K_r3_reg_0 (.CK( clk ) , .D( u2_uk_K_r2_0 ) , .Q( u2_uk_K_r3_0 ) , .QN( u2_uk_n1364 ) );
  DFF_X1 u2_uk_K_r3_reg_1 (.CK( clk ) , .D( u2_uk_K_r2_1 ) , .Q( u2_uk_K_r3_1 ) , .QN( u2_uk_n1365 ) );
  DFF_X1 u2_uk_K_r3_reg_10 (.CK( clk ) , .D( u2_uk_K_r2_10 ) , .Q( u2_uk_K_r3_10 ) );
  DFF_X1 u2_uk_K_r3_reg_11 (.CK( clk ) , .D( u2_uk_K_r2_11 ) , .Q( u2_uk_K_r3_11 ) );
  DFF_X1 u2_uk_K_r3_reg_12 (.CK( clk ) , .D( u2_uk_K_r2_12 ) , .Q( u2_uk_K_r3_12 ) , .QN( u2_uk_n1372 ) );
  DFF_X1 u2_uk_K_r3_reg_13 (.CK( clk ) , .D( u2_uk_K_r2_13 ) , .Q( u2_uk_K_r3_13 ) );
  DFF_X1 u2_uk_K_r3_reg_14 (.CK( clk ) , .D( u2_uk_K_r2_14 ) , .Q( u2_uk_K_r3_14 ) );
  DFF_X1 u2_uk_K_r3_reg_15 (.CK( clk ) , .D( u2_uk_K_r2_15 ) , .Q( u2_uk_K_r3_15 ) );
  DFF_X1 u2_uk_K_r3_reg_16 (.CK( clk ) , .D( u2_uk_K_r2_16 ) , .Q( u2_uk_K_r3_16 ) );
  DFF_X1 u2_uk_K_r3_reg_17 (.CK( clk ) , .D( u2_uk_K_r2_17 ) , .Q( u2_uk_K_r3_17 ) , .QN( u2_uk_n1373 ) );
  DFF_X1 u2_uk_K_r3_reg_18 (.CK( clk ) , .D( u2_uk_K_r2_18 ) , .Q( u2_uk_K_r3_18 ) , .QN( u2_uk_n1374 ) );
  DFF_X1 u2_uk_K_r3_reg_19 (.CK( clk ) , .D( u2_uk_K_r2_19 ) , .Q( u2_uk_K_r3_19 ) );
  DFF_X1 u2_uk_K_r3_reg_2 (.CK( clk ) , .D( u2_uk_K_r2_2 ) , .Q( u2_uk_K_r3_2 ) , .QN( u2_uk_n1366 ) );
  DFF_X1 u2_uk_K_r3_reg_20 (.CK( clk ) , .D( u2_uk_K_r2_20 ) , .Q( u2_uk_K_r3_20 ) , .QN( u2_uk_n1375 ) );
  DFF_X1 u2_uk_K_r3_reg_21 (.CK( clk ) , .D( u2_uk_K_r2_21 ) , .Q( u2_uk_K_r3_21 ) , .QN( u2_uk_n1376 ) );
  DFF_X1 u2_uk_K_r3_reg_22 (.CK( clk ) , .D( u2_uk_K_r2_22 ) , .Q( u2_uk_K_r3_22 ) , .QN( u2_uk_n1377 ) );
  DFF_X1 u2_uk_K_r3_reg_23 (.CK( clk ) , .D( u2_uk_K_r2_23 ) , .Q( u2_uk_K_r3_23 ) , .QN( u2_uk_n1378 ) );
  DFF_X1 u2_uk_K_r3_reg_24 (.CK( clk ) , .D( u2_uk_K_r2_24 ) , .Q( u2_uk_K_r3_24 ) );
  DFF_X1 u2_uk_K_r3_reg_25 (.CK( clk ) , .D( u2_uk_K_r2_25 ) , .Q( u2_uk_K_r3_25 ) , .QN( u2_uk_n1379 ) );
  DFF_X1 u2_uk_K_r3_reg_26 (.CK( clk ) , .D( u2_uk_K_r2_26 ) , .Q( u2_uk_K_r3_26 ) , .QN( u2_uk_n1380 ) );
  DFF_X1 u2_uk_K_r3_reg_27 (.CK( clk ) , .D( u2_uk_K_r2_27 ) , .Q( u2_uk_K_r3_27 ) , .QN( u2_uk_n1381 ) );
  DFF_X1 u2_uk_K_r3_reg_28 (.CK( clk ) , .D( u2_uk_K_r2_28 ) , .Q( u2_uk_K_r3_28 ) , .QN( u2_uk_n1382 ) );
  DFF_X1 u2_uk_K_r3_reg_29 (.CK( clk ) , .D( u2_uk_K_r2_29 ) , .Q( u2_uk_K_r3_29 ) );
  DFF_X1 u2_uk_K_r3_reg_3 (.CK( clk ) , .D( u2_uk_K_r2_3 ) , .Q( u2_uk_K_r3_3 ) , .QN( u2_uk_n1367 ) );
  DFF_X1 u2_uk_K_r3_reg_30 (.CK( clk ) , .D( u2_uk_K_r2_30 ) , .Q( u2_uk_K_r3_30 ) , .QN( u2_uk_n1383 ) );
  DFF_X1 u2_uk_K_r3_reg_31 (.CK( clk ) , .D( u2_uk_K_r2_31 ) , .Q( u2_uk_K_r3_31 ) , .QN( u2_uk_n1384 ) );
  DFF_X1 u2_uk_K_r3_reg_32 (.CK( clk ) , .D( u2_uk_K_r2_32 ) , .Q( u2_uk_K_r3_32 ) , .QN( u2_uk_n1385 ) );
  DFF_X1 u2_uk_K_r3_reg_33 (.CK( clk ) , .D( u2_uk_K_r2_33 ) , .Q( u2_uk_K_r3_33 ) , .QN( u2_uk_n1387 ) );
  DFF_X1 u2_uk_K_r3_reg_34 (.CK( clk ) , .D( u2_uk_K_r2_34 ) , .Q( u2_uk_K_r3_34 ) );
  DFF_X1 u2_uk_K_r3_reg_35 (.CK( clk ) , .D( u2_uk_K_r2_35 ) , .Q( u2_uk_K_r3_35 ) );
  DFF_X1 u2_uk_K_r3_reg_36 (.CK( clk ) , .D( u2_uk_K_r2_36 ) , .Q( u2_uk_K_r3_36 ) , .QN( u2_uk_n1388 ) );
  DFF_X1 u2_uk_K_r3_reg_37 (.CK( clk ) , .D( u2_uk_K_r2_37 ) , .Q( u2_uk_K_r3_37 ) , .QN( u2_uk_n1389 ) );
  DFF_X1 u2_uk_K_r3_reg_38 (.CK( clk ) , .D( u2_uk_K_r2_38 ) , .Q( u2_uk_K_r3_38 ) );
  DFF_X1 u2_uk_K_r3_reg_39 (.CK( clk ) , .D( u2_uk_K_r2_39 ) , .Q( u2_uk_K_r3_39 ) , .QN( u2_uk_n1392 ) );
  DFF_X1 u2_uk_K_r3_reg_4 (.CK( clk ) , .D( u2_uk_K_r2_4 ) , .Q( u2_uk_K_r3_4 ) );
  DFF_X1 u2_uk_K_r3_reg_40 (.CK( clk ) , .D( u2_uk_K_r2_40 ) , .Q( u2_uk_K_r3_40 ) , .QN( u2_uk_n1393 ) );
  DFF_X1 u2_uk_K_r3_reg_41 (.CK( clk ) , .D( u2_uk_K_r2_41 ) , .Q( u2_uk_K_r3_41 ) , .QN( u2_uk_n1394 ) );
  DFF_X1 u2_uk_K_r3_reg_42 (.CK( clk ) , .D( u2_uk_K_r2_42 ) , .Q( u2_uk_K_r3_42 ) , .QN( u2_uk_n1395 ) );
  DFF_X1 u2_uk_K_r3_reg_43 (.CK( clk ) , .D( u2_uk_K_r2_43 ) , .Q( u2_uk_K_r3_43 ) );
  DFF_X1 u2_uk_K_r3_reg_44 (.CK( clk ) , .D( u2_uk_K_r2_44 ) , .Q( u2_uk_K_r3_44 ) );
  DFF_X1 u2_uk_K_r3_reg_45 (.CK( clk ) , .D( u2_uk_K_r2_45 ) , .Q( u2_uk_K_r3_45 ) , .QN( u2_uk_n1396 ) );
  DFF_X1 u2_uk_K_r3_reg_46 (.CK( clk ) , .D( u2_uk_K_r2_46 ) , .Q( u2_uk_K_r3_46 ) , .QN( u2_uk_n1397 ) );
  DFF_X1 u2_uk_K_r3_reg_47 (.CK( clk ) , .D( u2_uk_K_r2_47 ) , .Q( u2_uk_K_r3_47 ) );
  DFF_X1 u2_uk_K_r3_reg_48 (.CK( clk ) , .D( u2_uk_K_r2_48 ) , .Q( u2_uk_K_r3_48 ) , .QN( u2_uk_n1399 ) );
  DFF_X1 u2_uk_K_r3_reg_49 (.CK( clk ) , .D( u2_uk_K_r2_49 ) , .Q( u2_uk_K_r3_49 ) , .QN( u2_uk_n1400 ) );
  DFF_X1 u2_uk_K_r3_reg_5 (.CK( clk ) , .D( u2_uk_K_r2_5 ) , .Q( u2_uk_K_r3_5 ) , .QN( u2_uk_n1368 ) );
  DFF_X1 u2_uk_K_r3_reg_50 (.CK( clk ) , .D( u2_uk_K_r2_50 ) , .Q( u2_uk_K_r3_50 ) , .QN( u2_uk_n1401 ) );
  DFF_X1 u2_uk_K_r3_reg_51 (.CK( clk ) , .D( u2_uk_K_r2_51 ) , .Q( u2_uk_K_r3_51 ) , .QN( u2_uk_n1403 ) );
  DFF_X1 u2_uk_K_r3_reg_52 (.CK( clk ) , .D( u2_uk_K_r2_52 ) , .Q( u2_uk_K_r3_52 ) );
  DFF_X1 u2_uk_K_r3_reg_53 (.CK( clk ) , .D( u2_uk_K_r2_53 ) , .Q( u2_uk_K_r3_53 ) , .QN( u2_uk_n1405 ) );
  DFF_X1 u2_uk_K_r3_reg_54 (.CK( clk ) , .D( u2_uk_K_r2_54 ) , .Q( u2_uk_K_r3_54 ) , .QN( u2_uk_n1406 ) );
  DFF_X1 u2_uk_K_r3_reg_55 (.CK( clk ) , .D( u2_uk_K_r2_55 ) , .Q( u2_uk_K_r3_55 ) , .QN( u2_uk_n1407 ) );
  DFF_X1 u2_uk_K_r3_reg_6 (.CK( clk ) , .D( u2_uk_K_r2_6 ) , .Q( u2_uk_K_r3_6 ) , .QN( u2_uk_n1369 ) );
  DFF_X1 u2_uk_K_r3_reg_7 (.CK( clk ) , .D( u2_uk_K_r2_7 ) , .Q( u2_uk_K_r3_7 ) , .QN( u2_uk_n1370 ) );
  DFF_X1 u2_uk_K_r3_reg_8 (.CK( clk ) , .D( u2_uk_K_r2_8 ) , .Q( u2_uk_K_r3_8 ) , .QN( u2_uk_n1371 ) );
  DFF_X1 u2_uk_K_r3_reg_9 (.CK( clk ) , .D( u2_uk_K_r2_9 ) , .Q( u2_uk_K_r3_9 ) );
  DFF_X1 u2_uk_K_r4_reg_0 (.CK( clk ) , .D( u2_uk_K_r3_0 ) , .Q( u2_uk_K_r4_0 ) );
  DFF_X1 u2_uk_K_r4_reg_1 (.CK( clk ) , .D( u2_uk_K_r3_1 ) , .Q( u2_uk_K_r4_1 ) , .QN( u2_uk_n1408 ) );
  DFF_X1 u2_uk_K_r4_reg_10 (.CK( clk ) , .D( u2_uk_K_r3_10 ) , .Q( u2_uk_K_r4_10 ) , .QN( u2_uk_n1414 ) );
  DFF_X1 u2_uk_K_r4_reg_11 (.CK( clk ) , .D( u2_uk_K_r3_11 ) , .Q( u2_uk_K_r4_11 ) );
  DFF_X1 u2_uk_K_r4_reg_12 (.CK( clk ) , .D( u2_uk_K_r3_12 ) , .Q( u2_uk_K_r4_12 ) , .QN( u2_uk_n1416 ) );
  DFF_X1 u2_uk_K_r4_reg_13 (.CK( clk ) , .D( u2_uk_K_r3_13 ) , .Q( u2_uk_K_r4_13 ) , .QN( u2_uk_n1417 ) );
  DFF_X1 u2_uk_K_r4_reg_14 (.CK( clk ) , .D( u2_uk_K_r3_14 ) , .Q( u2_uk_K_r4_14 ) , .QN( u2_uk_n1418 ) );
  DFF_X1 u2_uk_K_r4_reg_15 (.CK( clk ) , .D( u2_uk_K_r3_15 ) , .Q( u2_uk_K_r4_15 ) , .QN( u2_uk_n1419 ) );
  DFF_X1 u2_uk_K_r4_reg_16 (.CK( clk ) , .D( u2_uk_K_r3_16 ) , .Q( u2_uk_K_r4_16 ) , .QN( u2_uk_n1420 ) );
  DFF_X1 u2_uk_K_r4_reg_17 (.CK( clk ) , .D( u2_uk_K_r3_17 ) , .Q( u2_uk_K_r4_17 ) );
  DFF_X1 u2_uk_K_r4_reg_18 (.CK( clk ) , .D( u2_uk_K_r3_18 ) , .Q( u2_uk_K_r4_18 ) );
  DFF_X1 u2_uk_K_r4_reg_19 (.CK( clk ) , .D( u2_uk_K_r3_19 ) , .Q( u2_uk_K_r4_19 ) , .QN( u2_uk_n1422 ) );
  DFF_X1 u2_uk_K_r4_reg_2 (.CK( clk ) , .D( u2_uk_K_r3_2 ) , .Q( u2_uk_K_r4_2 ) );
  DFF_X1 u2_uk_K_r4_reg_20 (.CK( clk ) , .D( u2_uk_K_r3_20 ) , .Q( u2_uk_K_r4_20 ) , .QN( u2_uk_n1423 ) );
  DFF_X1 u2_uk_K_r4_reg_21 (.CK( clk ) , .D( u2_uk_K_r3_21 ) , .Q( u2_uk_K_r4_21 ) , .QN( u2_uk_n1424 ) );
  DFF_X1 u2_uk_K_r4_reg_22 (.CK( clk ) , .D( u2_uk_K_r3_22 ) , .Q( u2_uk_K_r4_22 ) , .QN( u2_uk_n1425 ) );
  DFF_X1 u2_uk_K_r4_reg_23 (.CK( clk ) , .D( u2_uk_K_r3_23 ) , .Q( u2_uk_K_r4_23 ) );
  DFF_X1 u2_uk_K_r4_reg_24 (.CK( clk ) , .D( u2_uk_K_r3_24 ) , .Q( u2_uk_K_r4_24 ) );
  DFF_X1 u2_uk_K_r4_reg_25 (.CK( clk ) , .D( u2_uk_K_r3_25 ) , .Q( u2_uk_K_r4_25 ) , .QN( u2_uk_n1426 ) );
  DFF_X1 u2_uk_K_r4_reg_26 (.CK( clk ) , .D( u2_uk_K_r3_26 ) , .Q( u2_uk_K_r4_26 ) , .QN( u2_uk_n1427 ) );
  DFF_X1 u2_uk_K_r4_reg_27 (.CK( clk ) , .D( u2_uk_K_r3_27 ) , .Q( u2_uk_K_r4_27 ) );
  DFF_X1 u2_uk_K_r4_reg_28 (.CK( clk ) , .D( u2_uk_K_r3_28 ) , .Q( u2_uk_K_r4_28 ) , .QN( u2_uk_n1428 ) );
  DFF_X1 u2_uk_K_r4_reg_29 (.CK( clk ) , .D( u2_uk_K_r3_29 ) , .Q( u2_uk_K_r4_29 ) , .QN( u2_uk_n1429 ) );
  DFF_X1 u2_uk_K_r4_reg_3 (.CK( clk ) , .D( u2_uk_K_r3_3 ) , .Q( u2_uk_K_r4_3 ) );
  DFF_X1 u2_uk_K_r4_reg_30 (.CK( clk ) , .D( u2_uk_K_r3_30 ) , .Q( u2_uk_K_r4_30 ) , .QN( u2_uk_n1430 ) );
  DFF_X1 u2_uk_K_r4_reg_31 (.CK( clk ) , .D( u2_uk_K_r3_31 ) , .Q( u2_uk_K_r4_31 ) );
  DFF_X1 u2_uk_K_r4_reg_32 (.CK( clk ) , .D( u2_uk_K_r3_32 ) , .Q( u2_uk_K_r4_32 ) , .QN( u2_uk_n1431 ) );
  DFF_X1 u2_uk_K_r4_reg_33 (.CK( clk ) , .D( u2_uk_K_r3_33 ) , .Q( u2_uk_K_r4_33 ) );
  DFF_X1 u2_uk_K_r4_reg_34 (.CK( clk ) , .D( u2_uk_K_r3_34 ) , .Q( u2_uk_K_r4_34 ) , .QN( u2_uk_n1432 ) );
  DFF_X1 u2_uk_K_r4_reg_35 (.CK( clk ) , .D( u2_uk_K_r3_35 ) , .Q( u2_uk_K_r4_35 ) );
  DFF_X1 u2_uk_K_r4_reg_36 (.CK( clk ) , .D( u2_uk_K_r3_36 ) , .Q( u2_uk_K_r4_36 ) , .QN( u2_uk_n1433 ) );
  DFF_X1 u2_uk_K_r4_reg_37 (.CK( clk ) , .D( u2_uk_K_r3_37 ) , .Q( u2_uk_K_r4_37 ) , .QN( u2_uk_n1434 ) );
  DFF_X1 u2_uk_K_r4_reg_38 (.CK( clk ) , .D( u2_uk_K_r3_38 ) , .Q( u2_uk_K_r4_38 ) );
  DFF_X1 u2_uk_K_r4_reg_39 (.CK( clk ) , .D( u2_uk_K_r3_39 ) , .Q( u2_uk_K_r4_39 ) , .QN( u2_uk_n1435 ) );
  DFF_X1 u2_uk_K_r4_reg_4 (.CK( clk ) , .D( u2_uk_K_r3_4 ) , .Q( u2_uk_K_r4_4 ) , .QN( u2_uk_n1409 ) );
  DFF_X1 u2_uk_K_r4_reg_40 (.CK( clk ) , .D( u2_uk_K_r3_40 ) , .Q( u2_uk_K_r4_40 ) , .QN( u2_uk_n1436 ) );
  DFF_X1 u2_uk_K_r4_reg_41 (.CK( clk ) , .D( u2_uk_K_r3_41 ) , .Q( u2_uk_K_r4_41 ) );
  DFF_X1 u2_uk_K_r4_reg_42 (.CK( clk ) , .D( u2_uk_K_r3_42 ) , .Q( u2_uk_K_r4_42 ) , .QN( u2_uk_n1438 ) );
  DFF_X1 u2_uk_K_r4_reg_43 (.CK( clk ) , .D( u2_uk_K_r3_43 ) , .Q( u2_uk_K_r4_43 ) , .QN( u2_uk_n1439 ) );
  DFF_X1 u2_uk_K_r4_reg_44 (.CK( clk ) , .D( u2_uk_K_r3_44 ) , .Q( u2_uk_K_r4_44 ) , .QN( u2_uk_n1440 ) );
  DFF_X1 u2_uk_K_r4_reg_45 (.CK( clk ) , .D( u2_uk_K_r3_45 ) , .Q( u2_uk_K_r4_45 ) , .QN( u2_uk_n1441 ) );
  DFF_X1 u2_uk_K_r4_reg_46 (.CK( clk ) , .D( u2_uk_K_r3_46 ) , .Q( u2_uk_K_r4_46 ) , .QN( u2_uk_n1442 ) );
  DFF_X1 u2_uk_K_r4_reg_47 (.CK( clk ) , .D( u2_uk_K_r3_47 ) , .Q( u2_uk_K_r4_47 ) , .QN( u2_uk_n1444 ) );
  DFF_X1 u2_uk_K_r4_reg_48 (.CK( clk ) , .D( u2_uk_K_r3_48 ) , .Q( u2_uk_K_r4_48 ) );
  DFF_X1 u2_uk_K_r4_reg_49 (.CK( clk ) , .D( u2_uk_K_r3_49 ) , .Q( u2_uk_K_r4_49 ) );
  DFF_X1 u2_uk_K_r4_reg_5 (.CK( clk ) , .D( u2_uk_K_r3_5 ) , .Q( u2_uk_K_r4_5 ) );
  DFF_X1 u2_uk_K_r4_reg_50 (.CK( clk ) , .D( u2_uk_K_r3_50 ) , .Q( u2_uk_K_r4_50 ) , .QN( u2_uk_n1445 ) );
  DFF_X1 u2_uk_K_r4_reg_51 (.CK( clk ) , .D( u2_uk_K_r3_51 ) , .Q( u2_uk_K_r4_51 ) , .QN( u2_uk_n1446 ) );
  DFF_X1 u2_uk_K_r4_reg_52 (.CK( clk ) , .D( u2_uk_K_r3_52 ) , .Q( u2_uk_K_r4_52 ) , .QN( u2_uk_n1447 ) );
  DFF_X1 u2_uk_K_r4_reg_53 (.CK( clk ) , .D( u2_uk_K_r3_53 ) , .Q( u2_uk_K_r4_53 ) , .QN( u2_uk_n1448 ) );
  DFF_X1 u2_uk_K_r4_reg_54 (.CK( clk ) , .D( u2_uk_K_r3_54 ) , .Q( u2_uk_K_r4_54 ) );
  DFF_X1 u2_uk_K_r4_reg_55 (.CK( clk ) , .D( u2_uk_K_r3_55 ) , .Q( u2_uk_K_r4_55 ) );
  DFF_X1 u2_uk_K_r4_reg_6 (.CK( clk ) , .D( u2_uk_K_r3_6 ) , .Q( u2_uk_K_r4_6 ) , .QN( u2_uk_n1410 ) );
  DFF_X1 u2_uk_K_r4_reg_7 (.CK( clk ) , .D( u2_uk_K_r3_7 ) , .Q( u2_uk_K_r4_7 ) , .QN( u2_uk_n1411 ) );
  DFF_X1 u2_uk_K_r4_reg_8 (.CK( clk ) , .D( u2_uk_K_r3_8 ) , .Q( u2_uk_K_r4_8 ) , .QN( u2_uk_n1412 ) );
  DFF_X1 u2_uk_K_r4_reg_9 (.CK( clk ) , .D( u2_uk_K_r3_9 ) , .Q( u2_uk_K_r4_9 ) , .QN( u2_uk_n1413 ) );
  DFF_X1 u2_uk_K_r5_reg_0 (.CK( clk ) , .D( u2_uk_K_r4_0 ) , .Q( u2_uk_K_r5_0 ) );
  DFF_X1 u2_uk_K_r5_reg_1 (.CK( clk ) , .D( u2_uk_K_r4_1 ) , .Q( u2_uk_K_r5_1 ) );
  DFF_X1 u2_uk_K_r5_reg_10 (.CK( clk ) , .D( u2_uk_K_r4_10 ) , .Q( u2_uk_K_r5_10 ) );
  DFF_X1 u2_uk_K_r5_reg_11 (.CK( clk ) , .D( u2_uk_K_r4_11 ) , .Q( u2_uk_K_r5_11 ) , .QN( u2_uk_n1457 ) );
  DFF_X1 u2_uk_K_r5_reg_12 (.CK( clk ) , .D( u2_uk_K_r4_12 ) , .Q( u2_uk_K_r5_12 ) , .QN( u2_uk_n1458 ) );
  DFF_X1 u2_uk_K_r5_reg_13 (.CK( clk ) , .D( u2_uk_K_r4_13 ) , .Q( u2_uk_K_r5_13 ) );
  DFF_X1 u2_uk_K_r5_reg_14 (.CK( clk ) , .D( u2_uk_K_r4_14 ) , .Q( u2_uk_K_r5_14 ) , .QN( u2_uk_n1459 ) );
  DFF_X1 u2_uk_K_r5_reg_15 (.CK( clk ) , .D( u2_uk_K_r4_15 ) , .Q( u2_uk_K_r5_15 ) , .QN( u2_uk_n1460 ) );
  DFF_X1 u2_uk_K_r5_reg_16 (.CK( clk ) , .D( u2_uk_K_r4_16 ) , .Q( u2_uk_K_r5_16 ) );
  DFF_X1 u2_uk_K_r5_reg_17 (.CK( clk ) , .D( u2_uk_K_r4_17 ) , .Q( u2_uk_K_r5_17 ) , .QN( u2_uk_n1461 ) );
  DFF_X1 u2_uk_K_r5_reg_18 (.CK( clk ) , .D( u2_uk_K_r4_18 ) , .Q( u2_uk_K_r5_18 ) );
  DFF_X1 u2_uk_K_r5_reg_19 (.CK( clk ) , .D( u2_uk_K_r4_19 ) , .Q( u2_uk_K_r5_19 ) );
  DFF_X1 u2_uk_K_r5_reg_2 (.CK( clk ) , .D( u2_uk_K_r4_2 ) , .Q( u2_uk_K_r5_2 ) , .QN( u2_uk_n1452 ) );
  DFF_X1 u2_uk_K_r5_reg_20 (.CK( clk ) , .D( u2_uk_K_r4_20 ) , .Q( u2_uk_K_r5_20 ) , .QN( u2_uk_n1462 ) );
  DFF_X1 u2_uk_K_r5_reg_21 (.CK( clk ) , .D( u2_uk_K_r4_21 ) , .Q( u2_uk_K_r5_21 ) );
  DFF_X1 u2_uk_K_r5_reg_22 (.CK( clk ) , .D( u2_uk_K_r4_22 ) , .Q( u2_uk_K_r5_22 ) , .QN( u2_uk_n1464 ) );
  DFF_X1 u2_uk_K_r5_reg_23 (.CK( clk ) , .D( u2_uk_K_r4_23 ) , .Q( u2_uk_K_r5_23 ) );
  DFF_X1 u2_uk_K_r5_reg_24 (.CK( clk ) , .D( u2_uk_K_r4_24 ) , .Q( u2_uk_K_r5_24 ) , .QN( u2_uk_n1465 ) );
  DFF_X1 u2_uk_K_r5_reg_25 (.CK( clk ) , .D( u2_uk_K_r4_25 ) , .Q( u2_uk_K_r5_25 ) , .QN( u2_uk_n1466 ) );
  DFF_X1 u2_uk_K_r5_reg_26 (.CK( clk ) , .D( u2_uk_K_r4_26 ) , .Q( u2_uk_K_r5_26 ) );
  DFF_X1 u2_uk_K_r5_reg_27 (.CK( clk ) , .D( u2_uk_K_r4_27 ) , .Q( u2_uk_K_r5_27 ) , .QN( u2_uk_n1468 ) );
  DFF_X1 u2_uk_K_r5_reg_28 (.CK( clk ) , .D( u2_uk_K_r4_28 ) , .Q( u2_uk_K_r5_28 ) , .QN( u2_uk_n1469 ) );
  DFF_X1 u2_uk_K_r5_reg_29 (.CK( clk ) , .D( u2_uk_K_r4_29 ) , .Q( u2_uk_K_r5_29 ) , .QN( u2_uk_n1470 ) );
  DFF_X1 u2_uk_K_r5_reg_3 (.CK( clk ) , .D( u2_uk_K_r4_3 ) , .Q( u2_uk_K_r5_3 ) , .QN( u2_uk_n1453 ) );
  DFF_X1 u2_uk_K_r5_reg_30 (.CK( clk ) , .D( u2_uk_K_r4_30 ) , .Q( u2_uk_K_r5_30 ) , .QN( u2_uk_n1471 ) );
  DFF_X1 u2_uk_K_r5_reg_31 (.CK( clk ) , .D( u2_uk_K_r4_31 ) , .Q( u2_uk_K_r5_31 ) );
  DFF_X1 u2_uk_K_r5_reg_32 (.CK( clk ) , .D( u2_uk_K_r4_32 ) , .Q( u2_uk_K_r5_32 ) );
  DFF_X1 u2_uk_K_r5_reg_33 (.CK( clk ) , .D( u2_uk_K_r4_33 ) , .Q( u2_uk_K_r5_33 ) , .QN( u2_uk_n1474 ) );
  DFF_X1 u2_uk_K_r5_reg_34 (.CK( clk ) , .D( u2_uk_K_r4_34 ) , .Q( u2_uk_K_r5_34 ) , .QN( u2_uk_n1475 ) );
  DFF_X1 u2_uk_K_r5_reg_35 (.CK( clk ) , .D( u2_uk_K_r4_35 ) , .Q( u2_uk_K_r5_35 ) , .QN( u2_uk_n1477 ) );
  DFF_X1 u2_uk_K_r5_reg_36 (.CK( clk ) , .D( u2_uk_K_r4_36 ) , .Q( u2_uk_K_r5_36 ) , .QN( u2_uk_n1478 ) );
  DFF_X1 u2_uk_K_r5_reg_37 (.CK( clk ) , .D( u2_uk_K_r4_37 ) , .Q( u2_uk_K_r5_37 ) );
  DFF_X1 u2_uk_K_r5_reg_38 (.CK( clk ) , .D( u2_uk_K_r4_38 ) , .Q( u2_uk_K_r5_38 ) , .QN( u2_uk_n1480 ) );
  DFF_X1 u2_uk_K_r5_reg_39 (.CK( clk ) , .D( u2_uk_K_r4_39 ) , .Q( u2_uk_K_r5_39 ) );
  DFF_X1 u2_uk_K_r5_reg_4 (.CK( clk ) , .D( u2_uk_K_r4_4 ) , .Q( u2_uk_K_r5_4 ) );
  DFF_X1 u2_uk_K_r5_reg_40 (.CK( clk ) , .D( u2_uk_K_r4_40 ) , .Q( u2_uk_K_r5_40 ) );
  DFF_X1 u2_uk_K_r5_reg_41 (.CK( clk ) , .D( u2_uk_K_r4_41 ) , .Q( u2_uk_K_r5_41 ) );
  DFF_X1 u2_uk_K_r5_reg_42 (.CK( clk ) , .D( u2_uk_K_r4_42 ) , .Q( u2_uk_K_r5_42 ) , .QN( u2_uk_n1484 ) );
  DFF_X1 u2_uk_K_r5_reg_43 (.CK( clk ) , .D( u2_uk_K_r4_43 ) , .Q( u2_uk_K_r5_43 ) );
  DFF_X1 u2_uk_K_r5_reg_44 (.CK( clk ) , .D( u2_uk_K_r4_44 ) , .Q( u2_uk_K_r5_44 ) , .QN( u2_uk_n1486 ) );
  DFF_X1 u2_uk_K_r5_reg_45 (.CK( clk ) , .D( u2_uk_K_r4_45 ) , .Q( u2_uk_K_r5_45 ) );
  DFF_X1 u2_uk_K_r5_reg_46 (.CK( clk ) , .D( u2_uk_K_r4_46 ) , .Q( u2_uk_K_r5_46 ) , .QN( u2_uk_n1487 ) );
  DFF_X1 u2_uk_K_r5_reg_47 (.CK( clk ) , .D( u2_uk_K_r4_47 ) , .Q( u2_uk_K_r5_47 ) , .QN( u2_uk_n1488 ) );
  DFF_X1 u2_uk_K_r5_reg_48 (.CK( clk ) , .D( u2_uk_K_r4_48 ) , .Q( u2_uk_K_r5_48 ) );
  DFF_X1 u2_uk_K_r5_reg_49 (.CK( clk ) , .D( u2_uk_K_r4_49 ) , .Q( u2_uk_K_r5_49 ) , .QN( u2_uk_n1490 ) );
  DFF_X1 u2_uk_K_r5_reg_5 (.CK( clk ) , .D( u2_uk_K_r4_5 ) , .Q( u2_uk_K_r5_5 ) );
  DFF_X1 u2_uk_K_r5_reg_50 (.CK( clk ) , .D( u2_uk_K_r4_50 ) , .Q( u2_uk_K_r5_50 ) , .QN( u2_uk_n1491 ) );
  DFF_X1 u2_uk_K_r5_reg_51 (.CK( clk ) , .D( u2_uk_K_r4_51 ) , .Q( u2_uk_K_r5_51 ) );
  DFF_X1 u2_uk_K_r5_reg_52 (.CK( clk ) , .D( u2_uk_K_r4_52 ) , .Q( u2_uk_K_r5_52 ) , .QN( u2_uk_n1493 ) );
  DFF_X1 u2_uk_K_r5_reg_53 (.CK( clk ) , .D( u2_uk_K_r4_53 ) , .Q( u2_uk_K_r5_53 ) , .QN( u2_uk_n1494 ) );
  DFF_X1 u2_uk_K_r5_reg_54 (.CK( clk ) , .D( u2_uk_K_r4_54 ) , .Q( u2_uk_K_r5_54 ) , .QN( u2_uk_n1496 ) );
  DFF_X1 u2_uk_K_r5_reg_55 (.CK( clk ) , .D( u2_uk_K_r4_55 ) , .Q( u2_uk_K_r5_55 ) , .QN( u2_uk_n1497 ) );
  DFF_X1 u2_uk_K_r5_reg_6 (.CK( clk ) , .D( u2_uk_K_r4_6 ) , .Q( u2_uk_K_r5_6 ) , .QN( u2_uk_n1454 ) );
  DFF_X1 u2_uk_K_r5_reg_7 (.CK( clk ) , .D( u2_uk_K_r4_7 ) , .Q( u2_uk_K_r5_7 ) , .QN( u2_uk_n1455 ) );
  DFF_X1 u2_uk_K_r5_reg_8 (.CK( clk ) , .D( u2_uk_K_r4_8 ) , .Q( u2_uk_K_r5_8 ) );
  DFF_X1 u2_uk_K_r5_reg_9 (.CK( clk ) , .D( u2_uk_K_r4_9 ) , .Q( u2_uk_K_r5_9 ) , .QN( u2_uk_n1456 ) );
  DFF_X1 u2_uk_K_r6_reg_0 (.CK( clk ) , .D( u2_uk_K_r5_0 ) , .Q( u2_uk_K_r6_0 ) );
  DFF_X1 u2_uk_K_r6_reg_1 (.CK( clk ) , .D( u2_uk_K_r5_1 ) , .Q( u2_uk_K_r6_1 ) , .QN( u2_uk_n1498 ) );
  DFF_X1 u2_uk_K_r6_reg_10 (.CK( clk ) , .D( u2_uk_K_r5_10 ) , .Q( u2_uk_K_r6_10 ) );
  DFF_X1 u2_uk_K_r6_reg_11 (.CK( clk ) , .D( u2_uk_K_r5_11 ) , .Q( u2_uk_K_r6_11 ) , .QN( u2_uk_n1506 ) );
  DFF_X1 u2_uk_K_r6_reg_12 (.CK( clk ) , .D( u2_uk_K_r5_12 ) , .Q( u2_uk_K_r6_12 ) , .QN( u2_uk_n1507 ) );
  DFF_X1 u2_uk_K_r6_reg_13 (.CK( clk ) , .D( u2_uk_K_r5_13 ) , .Q( u2_uk_K_r6_13 ) , .QN( u2_uk_n1508 ) );
  DFF_X1 u2_uk_K_r6_reg_14 (.CK( clk ) , .D( u2_uk_K_r5_14 ) , .Q( u2_uk_K_r6_14 ) );
  DFF_X1 u2_uk_K_r6_reg_15 (.CK( clk ) , .D( u2_uk_K_r5_15 ) , .Q( u2_uk_K_r6_15 ) , .QN( u2_uk_n1510 ) );
  DFF_X1 u2_uk_K_r6_reg_16 (.CK( clk ) , .D( u2_uk_K_r5_16 ) , .Q( u2_uk_K_r6_16 ) , .QN( u2_uk_n1511 ) );
  DFF_X1 u2_uk_K_r6_reg_17 (.CK( clk ) , .D( u2_uk_K_r5_17 ) , .Q( u2_uk_K_r6_17 ) , .QN( u2_uk_n1513 ) );
  DFF_X1 u2_uk_K_r6_reg_18 (.CK( clk ) , .D( u2_uk_K_r5_18 ) , .Q( u2_uk_K_r6_18 ) , .QN( u2_uk_n1514 ) );
  DFF_X1 u2_uk_K_r6_reg_19 (.CK( clk ) , .D( u2_uk_K_r5_19 ) , .Q( u2_uk_K_r6_19 ) );
  DFF_X1 u2_uk_K_r6_reg_2 (.CK( clk ) , .D( u2_uk_K_r5_2 ) , .Q( u2_uk_K_r6_2 ) , .QN( u2_uk_n1499 ) );
  DFF_X1 u2_uk_K_r6_reg_20 (.CK( clk ) , .D( u2_uk_K_r5_20 ) , .Q( u2_uk_K_r6_20 ) , .QN( u2_uk_n1515 ) );
  DFF_X1 u2_uk_K_r6_reg_21 (.CK( clk ) , .D( u2_uk_K_r5_21 ) , .Q( u2_uk_K_r6_21 ) );
  DFF_X1 u2_uk_K_r6_reg_22 (.CK( clk ) , .D( u2_uk_K_r5_22 ) , .Q( u2_uk_K_r6_22 ) );
  DFF_X1 u2_uk_K_r6_reg_23 (.CK( clk ) , .D( u2_uk_K_r5_23 ) , .Q( u2_uk_K_r6_23 ) , .QN( u2_uk_n1517 ) );
  DFF_X1 u2_uk_K_r6_reg_24 (.CK( clk ) , .D( u2_uk_K_r5_24 ) , .Q( u2_uk_K_r6_24 ) , .QN( u2_uk_n1518 ) );
  DFF_X1 u2_uk_K_r6_reg_25 (.CK( clk ) , .D( u2_uk_K_r5_25 ) , .Q( u2_uk_K_r6_25 ) , .QN( u2_uk_n1519 ) );
  DFF_X1 u2_uk_K_r6_reg_26 (.CK( clk ) , .D( u2_uk_K_r5_26 ) , .Q( u2_uk_K_r6_26 ) );
  DFF_X1 u2_uk_K_r6_reg_27 (.CK( clk ) , .D( u2_uk_K_r5_27 ) , .Q( u2_uk_K_r6_27 ) );
  DFF_X1 u2_uk_K_r6_reg_28 (.CK( clk ) , .D( u2_uk_K_r5_28 ) , .Q( u2_uk_K_r6_28 ) );
  DFF_X1 u2_uk_K_r6_reg_29 (.CK( clk ) , .D( u2_uk_K_r5_29 ) , .Q( u2_uk_K_r6_29 ) );
  DFF_X1 u2_uk_K_r6_reg_3 (.CK( clk ) , .D( u2_uk_K_r5_3 ) , .Q( u2_uk_K_r6_3 ) );
  DFF_X1 u2_uk_K_r6_reg_30 (.CK( clk ) , .D( u2_uk_K_r5_30 ) , .Q( u2_uk_K_r6_30 ) );
  DFF_X1 u2_uk_K_r6_reg_31 (.CK( clk ) , .D( u2_uk_K_r5_31 ) , .Q( u2_uk_K_r6_31 ) );
  DFF_X1 u2_uk_K_r6_reg_32 (.CK( clk ) , .D( u2_uk_K_r5_32 ) , .Q( u2_uk_K_r6_32 ) , .QN( u2_uk_n1521 ) );
  DFF_X1 u2_uk_K_r6_reg_33 (.CK( clk ) , .D( u2_uk_K_r5_33 ) , .Q( u2_uk_K_r6_33 ) , .QN( u2_uk_n1522 ) );
  DFF_X1 u2_uk_K_r6_reg_34 (.CK( clk ) , .D( u2_uk_K_r5_34 ) , .Q( u2_uk_K_r6_34 ) );
  DFF_X1 u2_uk_K_r6_reg_35 (.CK( clk ) , .D( u2_uk_K_r5_35 ) , .Q( u2_uk_K_r6_35 ) , .QN( u2_uk_n1524 ) );
  DFF_X1 u2_uk_K_r6_reg_36 (.CK( clk ) , .D( u2_uk_K_r5_36 ) , .Q( u2_uk_K_r6_36 ) , .QN( u2_uk_n1525 ) );
  DFF_X1 u2_uk_K_r6_reg_37 (.CK( clk ) , .D( u2_uk_K_r5_37 ) , .Q( u2_uk_K_r6_37 ) );
  DFF_X1 u2_uk_K_r6_reg_38 (.CK( clk ) , .D( u2_uk_K_r5_38 ) , .Q( u2_uk_K_r6_38 ) , .QN( u2_uk_n1526 ) );
  DFF_X1 u2_uk_K_r6_reg_39 (.CK( clk ) , .D( u2_uk_K_r5_39 ) , .Q( u2_uk_K_r6_39 ) , .QN( u2_uk_n1527 ) );
  DFF_X1 u2_uk_K_r6_reg_4 (.CK( clk ) , .D( u2_uk_K_r5_4 ) , .Q( u2_uk_K_r6_4 ) , .QN( u2_uk_n1500 ) );
  DFF_X1 u2_uk_K_r6_reg_40 (.CK( clk ) , .D( u2_uk_K_r5_40 ) , .Q( u2_uk_K_r6_40 ) , .QN( u2_uk_n1528 ) );
  DFF_X1 u2_uk_K_r6_reg_41 (.CK( clk ) , .D( u2_uk_K_r5_41 ) , .Q( u2_uk_K_r6_41 ) , .QN( u2_uk_n1529 ) );
  DFF_X1 u2_uk_K_r6_reg_42 (.CK( clk ) , .D( u2_uk_K_r5_42 ) , .Q( u2_uk_K_r6_42 ) , .QN( u2_uk_n1530 ) );
  DFF_X1 u2_uk_K_r6_reg_43 (.CK( clk ) , .D( u2_uk_K_r5_43 ) , .Q( u2_uk_K_r6_43 ) , .QN( u2_uk_n1531 ) );
  DFF_X1 u2_uk_K_r6_reg_44 (.CK( clk ) , .D( u2_uk_K_r5_44 ) , .Q( u2_uk_K_r6_44 ) , .QN( u2_uk_n1532 ) );
  DFF_X1 u2_uk_K_r6_reg_45 (.CK( clk ) , .D( u2_uk_K_r5_45 ) , .Q( u2_uk_K_r6_45 ) , .QN( u2_uk_n1533 ) );
  DFF_X1 u2_uk_K_r6_reg_46 (.CK( clk ) , .D( u2_uk_K_r5_46 ) , .Q( u2_uk_K_r6_46 ) );
  DFF_X1 u2_uk_K_r6_reg_47 (.CK( clk ) , .D( u2_uk_K_r5_47 ) , .Q( u2_uk_K_r6_47 ) , .QN( u2_uk_n1534 ) );
  DFF_X1 u2_uk_K_r6_reg_48 (.CK( clk ) , .D( u2_uk_K_r5_48 ) , .Q( u2_uk_K_r6_48 ) , .QN( u2_uk_n1535 ) );
  DFF_X1 u2_uk_K_r6_reg_49 (.CK( clk ) , .D( u2_uk_K_r5_49 ) , .Q( u2_uk_K_r6_49 ) , .QN( u2_uk_n1536 ) );
  DFF_X1 u2_uk_K_r6_reg_5 (.CK( clk ) , .D( u2_uk_K_r5_5 ) , .Q( u2_uk_K_r6_5 ) , .QN( u2_uk_n1501 ) );
  DFF_X1 u2_uk_K_r6_reg_50 (.CK( clk ) , .D( u2_uk_K_r5_50 ) , .Q( u2_uk_K_r6_50 ) , .QN( u2_uk_n1537 ) );
  DFF_X1 u2_uk_K_r6_reg_51 (.CK( clk ) , .D( u2_uk_K_r5_51 ) , .Q( u2_uk_K_r6_51 ) );
  DFF_X1 u2_uk_K_r6_reg_52 (.CK( clk ) , .D( u2_uk_K_r5_52 ) , .Q( u2_uk_K_r6_52 ) , .QN( u2_uk_n1538 ) );
  DFF_X1 u2_uk_K_r6_reg_53 (.CK( clk ) , .D( u2_uk_K_r5_53 ) , .Q( u2_uk_K_r6_53 ) );
  DFF_X1 u2_uk_K_r6_reg_54 (.CK( clk ) , .D( u2_uk_K_r5_54 ) , .Q( u2_uk_K_r6_54 ) , .QN( u2_uk_n1540 ) );
  DFF_X1 u2_uk_K_r6_reg_55 (.CK( clk ) , .D( u2_uk_K_r5_55 ) , .Q( u2_uk_K_r6_55 ) );
  DFF_X1 u2_uk_K_r6_reg_6 (.CK( clk ) , .D( u2_uk_K_r5_6 ) , .Q( u2_uk_K_r6_6 ) , .QN( u2_uk_n1502 ) );
  DFF_X1 u2_uk_K_r6_reg_7 (.CK( clk ) , .D( u2_uk_K_r5_7 ) , .Q( u2_uk_K_r6_7 ) );
  DFF_X1 u2_uk_K_r6_reg_8 (.CK( clk ) , .D( u2_uk_K_r5_8 ) , .Q( u2_uk_K_r6_8 ) , .QN( u2_uk_n1503 ) );
  DFF_X1 u2_uk_K_r6_reg_9 (.CK( clk ) , .D( u2_uk_K_r5_9 ) , .Q( u2_uk_K_r6_9 ) , .QN( u2_uk_n1504 ) );
  DFF_X1 u2_uk_K_r7_reg_0 (.CK( clk ) , .D( u2_uk_K_r6_0 ) , .Q( u2_uk_K_r7_0 ) );
  DFF_X1 u2_uk_K_r7_reg_1 (.CK( clk ) , .D( u2_uk_K_r6_1 ) , .Q( u2_uk_K_r7_1 ) , .QN( u2_uk_n1541 ) );
  DFF_X1 u2_uk_K_r7_reg_10 (.CK( clk ) , .D( u2_uk_K_r6_10 ) , .Q( u2_uk_K_r7_10 ) , .QN( u2_uk_n1547 ) );
  DFF_X1 u2_uk_K_r7_reg_11 (.CK( clk ) , .D( u2_uk_K_r6_11 ) , .Q( u2_uk_K_r7_11 ) , .QN( u2_uk_n1548 ) );
  DFF_X1 u2_uk_K_r7_reg_12 (.CK( clk ) , .D( u2_uk_K_r6_12 ) , .Q( u2_uk_K_r7_12 ) , .QN( u2_uk_n1549 ) );
  DFF_X1 u2_uk_K_r7_reg_13 (.CK( clk ) , .D( u2_uk_K_r6_13 ) , .Q( u2_uk_K_r7_13 ) );
  DFF_X1 u2_uk_K_r7_reg_14 (.CK( clk ) , .D( u2_uk_K_r6_14 ) , .Q( u2_uk_K_r7_14 ) , .QN( u2_uk_n1551 ) );
  DFF_X1 u2_uk_K_r7_reg_15 (.CK( clk ) , .D( u2_uk_K_r6_15 ) , .Q( u2_uk_K_r7_15 ) );
  DFF_X1 u2_uk_K_r7_reg_16 (.CK( clk ) , .D( u2_uk_K_r6_16 ) , .Q( u2_uk_K_r7_16 ) );
  DFF_X1 u2_uk_K_r7_reg_17 (.CK( clk ) , .D( u2_uk_K_r6_17 ) , .Q( u2_uk_K_r7_17 ) , .QN( u2_uk_n1554 ) );
  DFF_X1 u2_uk_K_r7_reg_18 (.CK( clk ) , .D( u2_uk_K_r6_18 ) , .Q( u2_uk_K_r7_18 ) , .QN( u2_uk_n1555 ) );
  DFF_X1 u2_uk_K_r7_reg_19 (.CK( clk ) , .D( u2_uk_K_r6_19 ) , .Q( u2_uk_K_r7_19 ) , .QN( u2_uk_n1556 ) );
  DFF_X1 u2_uk_K_r7_reg_2 (.CK( clk ) , .D( u2_uk_K_r6_2 ) , .Q( u2_uk_K_r7_2 ) , .QN( u2_uk_n1542 ) );
  DFF_X1 u2_uk_K_r7_reg_20 (.CK( clk ) , .D( u2_uk_K_r6_20 ) , .Q( u2_uk_K_r7_20 ) );
  DFF_X1 u2_uk_K_r7_reg_21 (.CK( clk ) , .D( u2_uk_K_r6_21 ) , .Q( u2_uk_K_r7_21 ) , .QN( u2_uk_n1558 ) );
  DFF_X1 u2_uk_K_r7_reg_22 (.CK( clk ) , .D( u2_uk_K_r6_22 ) , .Q( u2_uk_K_r7_22 ) );
  DFF_X1 u2_uk_K_r7_reg_23 (.CK( clk ) , .D( u2_uk_K_r6_23 ) , .Q( u2_uk_K_r7_23 ) );
  DFF_X1 u2_uk_K_r7_reg_24 (.CK( clk ) , .D( u2_uk_K_r6_24 ) , .Q( u2_uk_K_r7_24 ) , .QN( u2_uk_n1562 ) );
  DFF_X1 u2_uk_K_r7_reg_25 (.CK( clk ) , .D( u2_uk_K_r6_25 ) , .Q( u2_uk_K_r7_25 ) , .QN( u2_uk_n1563 ) );
  DFF_X1 u2_uk_K_r7_reg_26 (.CK( clk ) , .D( u2_uk_K_r6_26 ) , .Q( u2_uk_K_r7_26 ) );
  DFF_X1 u2_uk_K_r7_reg_27 (.CK( clk ) , .D( u2_uk_K_r6_27 ) , .Q( u2_uk_K_r7_27 ) );
  DFF_X1 u2_uk_K_r7_reg_28 (.CK( clk ) , .D( u2_uk_K_r6_28 ) , .Q( u2_uk_K_r7_28 ) , .QN( u2_uk_n1565 ) );
  DFF_X1 u2_uk_K_r7_reg_29 (.CK( clk ) , .D( u2_uk_K_r6_29 ) , .Q( u2_uk_K_r7_29 ) );
  DFF_X1 u2_uk_K_r7_reg_3 (.CK( clk ) , .D( u2_uk_K_r6_3 ) , .Q( u2_uk_K_r7_3 ) , .QN( u2_uk_n1543 ) );
  DFF_X1 u2_uk_K_r7_reg_30 (.CK( clk ) , .D( u2_uk_K_r6_30 ) , .Q( u2_uk_K_r7_30 ) );
  DFF_X1 u2_uk_K_r7_reg_31 (.CK( clk ) , .D( u2_uk_K_r6_31 ) , .Q( u2_uk_K_r7_31 ) );
  DFF_X1 u2_uk_K_r7_reg_32 (.CK( clk ) , .D( u2_uk_K_r6_32 ) , .Q( u2_uk_K_r7_32 ) );
  DFF_X1 u2_uk_K_r7_reg_33 (.CK( clk ) , .D( u2_uk_K_r6_33 ) , .Q( u2_uk_K_r7_33 ) , .QN( u2_uk_n1568 ) );
  DFF_X1 u2_uk_K_r7_reg_34 (.CK( clk ) , .D( u2_uk_K_r6_34 ) , .Q( u2_uk_K_r7_34 ) );
  DFF_X1 u2_uk_K_r7_reg_35 (.CK( clk ) , .D( u2_uk_K_r6_35 ) , .Q( u2_uk_K_r7_35 ) , .QN( u2_uk_n1569 ) );
  DFF_X1 u2_uk_K_r7_reg_36 (.CK( clk ) , .D( u2_uk_K_r6_36 ) , .Q( u2_uk_K_r7_36 ) , .QN( u2_uk_n1570 ) );
  DFF_X1 u2_uk_K_r7_reg_37 (.CK( clk ) , .D( u2_uk_K_r6_37 ) , .Q( u2_uk_K_r7_37 ) );
  DFF_X1 u2_uk_K_r7_reg_38 (.CK( clk ) , .D( u2_uk_K_r6_38 ) , .Q( u2_uk_K_r7_38 ) , .QN( u2_uk_n1571 ) );
  DFF_X1 u2_uk_K_r7_reg_39 (.CK( clk ) , .D( u2_uk_K_r6_39 ) , .Q( u2_uk_K_r7_39 ) );
  DFF_X1 u2_uk_K_r7_reg_4 (.CK( clk ) , .D( u2_uk_K_r6_4 ) , .Q( u2_uk_K_r7_4 ) , .QN( u2_uk_n1544 ) );
  DFF_X1 u2_uk_K_r7_reg_40 (.CK( clk ) , .D( u2_uk_K_r6_40 ) , .Q( u2_uk_K_r7_40 ) , .QN( u2_uk_n1573 ) );
  DFF_X1 u2_uk_K_r7_reg_41 (.CK( clk ) , .D( u2_uk_K_r6_41 ) , .Q( u2_uk_K_r7_41 ) , .QN( u2_uk_n1574 ) );
  DFF_X1 u2_uk_K_r7_reg_42 (.CK( clk ) , .D( u2_uk_K_r6_42 ) , .Q( u2_uk_K_r7_42 ) , .QN( u2_uk_n1575 ) );
  DFF_X1 u2_uk_K_r7_reg_43 (.CK( clk ) , .D( u2_uk_K_r6_43 ) , .Q( u2_uk_K_r7_43 ) , .QN( u2_uk_n1576 ) );
  DFF_X1 u2_uk_K_r7_reg_44 (.CK( clk ) , .D( u2_uk_K_r6_44 ) , .Q( u2_uk_K_r7_44 ) , .QN( u2_uk_n1577 ) );
  DFF_X1 u2_uk_K_r7_reg_45 (.CK( clk ) , .D( u2_uk_K_r6_45 ) , .Q( u2_uk_K_r7_45 ) , .QN( u2_uk_n1578 ) );
  DFF_X1 u2_uk_K_r7_reg_46 (.CK( clk ) , .D( u2_uk_K_r6_46 ) , .Q( u2_uk_K_r7_46 ) );
  DFF_X1 u2_uk_K_r7_reg_47 (.CK( clk ) , .D( u2_uk_K_r6_47 ) , .Q( u2_uk_K_r7_47 ) , .QN( u2_uk_n1580 ) );
  DFF_X1 u2_uk_K_r7_reg_48 (.CK( clk ) , .D( u2_uk_K_r6_48 ) , .Q( u2_uk_K_r7_48 ) );
  DFF_X1 u2_uk_K_r7_reg_49 (.CK( clk ) , .D( u2_uk_K_r6_49 ) , .Q( u2_uk_K_r7_49 ) , .QN( u2_uk_n1582 ) );
  DFF_X1 u2_uk_K_r7_reg_5 (.CK( clk ) , .D( u2_uk_K_r6_5 ) , .Q( u2_uk_K_r7_5 ) );
  DFF_X1 u2_uk_K_r7_reg_50 (.CK( clk ) , .D( u2_uk_K_r6_50 ) , .Q( u2_uk_K_r7_50 ) , .QN( u2_uk_n1583 ) );
  DFF_X1 u2_uk_K_r7_reg_51 (.CK( clk ) , .D( u2_uk_K_r6_51 ) , .Q( u2_uk_K_r7_51 ) , .QN( u2_uk_n1584 ) );
  DFF_X1 u2_uk_K_r7_reg_52 (.CK( clk ) , .D( u2_uk_K_r6_52 ) , .Q( u2_uk_K_r7_52 ) , .QN( u2_uk_n1585 ) );
  DFF_X1 u2_uk_K_r7_reg_53 (.CK( clk ) , .D( u2_uk_K_r6_53 ) , .Q( u2_uk_K_r7_53 ) );
  DFF_X1 u2_uk_K_r7_reg_54 (.CK( clk ) , .D( u2_uk_K_r6_54 ) , .Q( u2_uk_K_r7_54 ) , .QN( u2_uk_n1586 ) );
  DFF_X1 u2_uk_K_r7_reg_55 (.CK( clk ) , .D( u2_uk_K_r6_55 ) , .Q( u2_uk_K_r7_55 ) );
  DFF_X1 u2_uk_K_r7_reg_6 (.CK( clk ) , .D( u2_uk_K_r6_6 ) , .Q( u2_uk_K_r7_6 ) );
  DFF_X1 u2_uk_K_r7_reg_7 (.CK( clk ) , .D( u2_uk_K_r6_7 ) , .Q( u2_uk_K_r7_7 ) );
  DFF_X1 u2_uk_K_r7_reg_8 (.CK( clk ) , .D( u2_uk_K_r6_8 ) , .Q( u2_uk_K_r7_8 ) );
  DFF_X1 u2_uk_K_r7_reg_9 (.CK( clk ) , .D( u2_uk_K_r6_9 ) , .Q( u2_uk_K_r7_9 ) );
  DFF_X1 u2_uk_K_r8_reg_0 (.CK( clk ) , .D( u2_uk_K_r7_0 ) , .Q( u2_uk_K_r8_0 ) , .QN( u2_uk_n1588 ) );
  DFF_X1 u2_uk_K_r8_reg_1 (.CK( clk ) , .D( u2_uk_K_r7_1 ) , .Q( u2_uk_K_r8_1 ) , .QN( u2_uk_n1589 ) );
  DFF_X1 u2_uk_K_r8_reg_10 (.CK( clk ) , .D( u2_uk_K_r7_10 ) , .Q( u2_uk_K_r8_10 ) );
  DFF_X1 u2_uk_K_r8_reg_11 (.CK( clk ) , .D( u2_uk_K_r7_11 ) , .Q( u2_uk_K_r8_11 ) , .QN( u2_uk_n1595 ) );
  DFF_X1 u2_uk_K_r8_reg_12 (.CK( clk ) , .D( u2_uk_K_r7_12 ) , .Q( u2_uk_K_r8_12 ) , .QN( u2_uk_n1596 ) );
  DFF_X1 u2_uk_K_r8_reg_13 (.CK( clk ) , .D( u2_uk_K_r7_13 ) , .Q( u2_uk_K_r8_13 ) );
  DFF_X1 u2_uk_K_r8_reg_14 (.CK( clk ) , .D( u2_uk_K_r7_14 ) , .Q( u2_uk_K_r8_14 ) , .QN( u2_uk_n1597 ) );
  DFF_X1 u2_uk_K_r8_reg_15 (.CK( clk ) , .D( u2_uk_K_r7_15 ) , .Q( u2_uk_K_r8_15 ) , .QN( u2_uk_n1598 ) );
  DFF_X1 u2_uk_K_r8_reg_16 (.CK( clk ) , .D( u2_uk_K_r7_16 ) , .Q( u2_uk_K_r8_16 ) );
  DFF_X1 u2_uk_K_r8_reg_17 (.CK( clk ) , .D( u2_uk_K_r7_17 ) , .Q( u2_uk_K_r8_17 ) );
  DFF_X1 u2_uk_K_r8_reg_18 (.CK( clk ) , .D( u2_uk_K_r7_18 ) , .Q( u2_uk_K_r8_18 ) , .QN( u2_uk_n1599 ) );
  DFF_X1 u2_uk_K_r8_reg_19 (.CK( clk ) , .D( u2_uk_K_r7_19 ) , .Q( u2_uk_K_r8_19 ) );
  DFF_X1 u2_uk_K_r8_reg_2 (.CK( clk ) , .D( u2_uk_K_r7_2 ) , .Q( u2_uk_K_r8_2 ) );
  DFF_X1 u2_uk_K_r8_reg_20 (.CK( clk ) , .D( u2_uk_K_r7_20 ) , .Q( u2_uk_K_r8_20 ) , .QN( u2_uk_n1600 ) );
  DFF_X1 u2_uk_K_r8_reg_21 (.CK( clk ) , .D( u2_uk_K_r7_21 ) , .Q( u2_uk_K_r8_21 ) );
  DFF_X1 u2_uk_K_r8_reg_22 (.CK( clk ) , .D( u2_uk_K_r7_22 ) , .Q( u2_uk_K_r8_22 ) );
  DFF_X1 u2_uk_K_r8_reg_23 (.CK( clk ) , .D( u2_uk_K_r7_23 ) , .Q( u2_uk_K_r8_23 ) , .QN( u2_uk_n1602 ) );
  DFF_X1 u2_uk_K_r8_reg_24 (.CK( clk ) , .D( u2_uk_K_r7_24 ) , .Q( u2_uk_K_r8_24 ) , .QN( u2_uk_n1603 ) );
  DFF_X1 u2_uk_K_r8_reg_25 (.CK( clk ) , .D( u2_uk_K_r7_25 ) , .Q( u2_uk_K_r8_25 ) , .QN( u2_uk_n1604 ) );
  DFF_X1 u2_uk_K_r8_reg_26 (.CK( clk ) , .D( u2_uk_K_r7_26 ) , .Q( u2_uk_K_r8_26 ) , .QN( u2_uk_n1605 ) );
  DFF_X1 u2_uk_K_r8_reg_27 (.CK( clk ) , .D( u2_uk_K_r7_27 ) , .Q( u2_uk_K_r8_27 ) );
  DFF_X1 u2_uk_K_r8_reg_28 (.CK( clk ) , .D( u2_uk_K_r7_28 ) , .Q( u2_uk_K_r8_28 ) );
  DFF_X1 u2_uk_K_r8_reg_29 (.CK( clk ) , .D( u2_uk_K_r7_29 ) , .Q( u2_uk_K_r8_29 ) , .QN( u2_uk_n1609 ) );
  DFF_X1 u2_uk_K_r8_reg_3 (.CK( clk ) , .D( u2_uk_K_r7_3 ) , .Q( u2_uk_K_r8_3 ) , .QN( u2_uk_n1590 ) );
  DFF_X1 u2_uk_K_r8_reg_30 (.CK( clk ) , .D( u2_uk_K_r7_30 ) , .Q( u2_uk_K_r8_30 ) , .QN( u2_uk_n1610 ) );
  DFF_X1 u2_uk_K_r8_reg_31 (.CK( clk ) , .D( u2_uk_K_r7_31 ) , .Q( u2_uk_K_r8_31 ) , .QN( u2_uk_n1611 ) );
  DFF_X1 u2_uk_K_r8_reg_32 (.CK( clk ) , .D( u2_uk_K_r7_32 ) , .Q( u2_uk_K_r8_32 ) );
  DFF_X1 u2_uk_K_r8_reg_33 (.CK( clk ) , .D( u2_uk_K_r7_33 ) , .Q( u2_uk_K_r8_33 ) , .QN( u2_uk_n1612 ) );
  DFF_X1 u2_uk_K_r8_reg_34 (.CK( clk ) , .D( u2_uk_K_r7_34 ) , .Q( u2_uk_K_r8_34 ) , .QN( u2_uk_n1613 ) );
  DFF_X1 u2_uk_K_r8_reg_35 (.CK( clk ) , .D( u2_uk_K_r7_35 ) , .Q( u2_uk_K_r8_35 ) , .QN( u2_uk_n1614 ) );
  DFF_X1 u2_uk_K_r8_reg_36 (.CK( clk ) , .D( u2_uk_K_r7_36 ) , .Q( u2_uk_K_r8_36 ) , .QN( u2_uk_n1615 ) );
  DFF_X1 u2_uk_K_r8_reg_37 (.CK( clk ) , .D( u2_uk_K_r7_37 ) , .Q( u2_uk_K_r8_37 ) );
  DFF_X1 u2_uk_K_r8_reg_38 (.CK( clk ) , .D( u2_uk_K_r7_38 ) , .Q( u2_uk_K_r8_38 ) , .QN( u2_uk_n1617 ) );
  DFF_X1 u2_uk_K_r8_reg_39 (.CK( clk ) , .D( u2_uk_K_r7_39 ) , .Q( u2_uk_K_r8_39 ) , .QN( u2_uk_n1619 ) );
  DFF_X1 u2_uk_K_r8_reg_4 (.CK( clk ) , .D( u2_uk_K_r7_4 ) , .Q( u2_uk_K_r8_4 ) , .QN( u2_uk_n1591 ) );
  DFF_X1 u2_uk_K_r8_reg_40 (.CK( clk ) , .D( u2_uk_K_r7_40 ) , .Q( u2_uk_K_r8_40 ) );
  DFF_X1 u2_uk_K_r8_reg_41 (.CK( clk ) , .D( u2_uk_K_r7_41 ) , .Q( u2_uk_K_r8_41 ) );
  DFF_X1 u2_uk_K_r8_reg_42 (.CK( clk ) , .D( u2_uk_K_r7_42 ) , .Q( u2_uk_K_r8_42 ) , .QN( u2_uk_n1621 ) );
  DFF_X1 u2_uk_K_r8_reg_43 (.CK( clk ) , .D( u2_uk_K_r7_43 ) , .Q( u2_uk_K_r8_43 ) );
  DFF_X1 u2_uk_K_r8_reg_44 (.CK( clk ) , .D( u2_uk_K_r7_44 ) , .Q( u2_uk_K_r8_44 ) , .QN( u2_uk_n1622 ) );
  DFF_X1 u2_uk_K_r8_reg_45 (.CK( clk ) , .D( u2_uk_K_r7_45 ) , .Q( u2_uk_K_r8_45 ) );
  DFF_X1 u2_uk_K_r8_reg_46 (.CK( clk ) , .D( u2_uk_K_r7_46 ) , .Q( u2_uk_K_r8_46 ) , .QN( u2_uk_n1623 ) );
  DFF_X1 u2_uk_K_r8_reg_47 (.CK( clk ) , .D( u2_uk_K_r7_47 ) , .Q( u2_uk_K_r8_47 ) , .QN( u2_uk_n1624 ) );
  DFF_X1 u2_uk_K_r8_reg_48 (.CK( clk ) , .D( u2_uk_K_r7_48 ) , .Q( u2_uk_K_r8_48 ) );
  DFF_X1 u2_uk_K_r8_reg_49 (.CK( clk ) , .D( u2_uk_K_r7_49 ) , .Q( u2_uk_K_r8_49 ) , .QN( u2_uk_n1625 ) );
  DFF_X1 u2_uk_K_r8_reg_5 (.CK( clk ) , .D( u2_uk_K_r7_5 ) , .Q( u2_uk_K_r8_5 ) );
  DFF_X1 u2_uk_K_r8_reg_50 (.CK( clk ) , .D( u2_uk_K_r7_50 ) , .Q( u2_uk_K_r8_50 ) , .QN( u2_uk_n1626 ) );
  DFF_X1 u2_uk_K_r8_reg_51 (.CK( clk ) , .D( u2_uk_K_r7_51 ) , .Q( u2_uk_K_r8_51 ) );
  DFF_X1 u2_uk_K_r8_reg_52 (.CK( clk ) , .D( u2_uk_K_r7_52 ) , .Q( u2_uk_K_r8_52 ) );
  DFF_X1 u2_uk_K_r8_reg_53 (.CK( clk ) , .D( u2_uk_K_r7_53 ) , .Q( u2_uk_K_r8_53 ) , .QN( u2_uk_n1629 ) );
  DFF_X1 u2_uk_K_r8_reg_54 (.CK( clk ) , .D( u2_uk_K_r7_54 ) , .Q( u2_uk_K_r8_54 ) , .QN( u2_uk_n1630 ) );
  DFF_X1 u2_uk_K_r8_reg_55 (.CK( clk ) , .D( u2_uk_K_r7_55 ) , .Q( u2_uk_K_r8_55 ) , .QN( u2_uk_n1631 ) );
  DFF_X1 u2_uk_K_r8_reg_6 (.CK( clk ) , .D( u2_uk_K_r7_6 ) , .Q( u2_uk_K_r8_6 ) , .QN( u2_uk_n1592 ) );
  DFF_X1 u2_uk_K_r8_reg_7 (.CK( clk ) , .D( u2_uk_K_r7_7 ) , .Q( u2_uk_K_r8_7 ) , .QN( u2_uk_n1593 ) );
  DFF_X1 u2_uk_K_r8_reg_8 (.CK( clk ) , .D( u2_uk_K_r7_8 ) , .Q( u2_uk_K_r8_8 ) );
  DFF_X1 u2_uk_K_r8_reg_9 (.CK( clk ) , .D( u2_uk_K_r7_9 ) , .Q( u2_uk_K_r8_9 ) , .QN( u2_uk_n1594 ) );
  DFF_X1 u2_uk_K_r9_reg_0 (.CK( clk ) , .D( u2_uk_K_r8_0 ) , .Q( u2_uk_K_r9_0 ) );
  DFF_X1 u2_uk_K_r9_reg_1 (.CK( clk ) , .D( u2_uk_K_r8_1 ) , .Q( u2_uk_K_r9_1 ) , .QN( u2_uk_n1632 ) );
  DFF_X1 u2_uk_K_r9_reg_10 (.CK( clk ) , .D( u2_uk_K_r8_10 ) , .Q( u2_uk_K_r9_10 ) );
  DFF_X1 u2_uk_K_r9_reg_11 (.CK( clk ) , .D( u2_uk_K_r8_11 ) , .Q( u2_uk_K_r9_11 ) , .QN( u2_uk_n1637 ) );
  DFF_X1 u2_uk_K_r9_reg_12 (.CK( clk ) , .D( u2_uk_K_r8_12 ) , .Q( u2_uk_K_r9_12 ) );
  DFF_X1 u2_uk_K_r9_reg_13 (.CK( clk ) , .D( u2_uk_K_r8_13 ) , .Q( u2_uk_K_r9_13 ) , .QN( u2_uk_n1639 ) );
  DFF_X1 u2_uk_K_r9_reg_14 (.CK( clk ) , .D( u2_uk_K_r8_14 ) , .Q( u2_uk_K_r9_14 ) , .QN( u2_uk_n1640 ) );
  DFF_X1 u2_uk_K_r9_reg_15 (.CK( clk ) , .D( u2_uk_K_r8_15 ) , .Q( u2_uk_K_r9_15 ) );
  DFF_X1 u2_uk_K_r9_reg_16 (.CK( clk ) , .D( u2_uk_K_r8_16 ) , .Q( u2_uk_K_r9_16 ) , .QN( u2_uk_n1642 ) );
  DFF_X1 u2_uk_K_r9_reg_17 (.CK( clk ) , .D( u2_uk_K_r8_17 ) , .Q( u2_uk_K_r9_17 ) , .QN( u2_uk_n1643 ) );
  DFF_X1 u2_uk_K_r9_reg_18 (.CK( clk ) , .D( u2_uk_K_r8_18 ) , .Q( u2_uk_K_r9_18 ) );
  DFF_X1 u2_uk_K_r9_reg_19 (.CK( clk ) , .D( u2_uk_K_r8_19 ) , .Q( u2_uk_K_r9_19 ) );
  DFF_X1 u2_uk_K_r9_reg_2 (.CK( clk ) , .D( u2_uk_K_r8_2 ) , .Q( u2_uk_K_r9_2 ) );
  DFF_X1 u2_uk_K_r9_reg_20 (.CK( clk ) , .D( u2_uk_K_r8_20 ) , .Q( u2_uk_K_r9_20 ) , .QN( u2_uk_n1646 ) );
  DFF_X1 u2_uk_K_r9_reg_21 (.CK( clk ) , .D( u2_uk_K_r8_21 ) , .Q( u2_uk_K_r9_21 ) , .QN( u2_uk_n1647 ) );
  DFF_X1 u2_uk_K_r9_reg_22 (.CK( clk ) , .D( u2_uk_K_r8_22 ) , .Q( u2_uk_K_r9_22 ) , .QN( u2_uk_n1648 ) );
  DFF_X1 u2_uk_K_r9_reg_23 (.CK( clk ) , .D( u2_uk_K_r8_23 ) , .Q( u2_uk_K_r9_23 ) );
  DFF_X1 u2_uk_K_r9_reg_24 (.CK( clk ) , .D( u2_uk_K_r8_24 ) , .Q( u2_uk_K_r9_24 ) );
  DFF_X1 u2_uk_K_r9_reg_25 (.CK( clk ) , .D( u2_uk_K_r8_25 ) , .Q( u2_uk_K_r9_25 ) );
  DFF_X1 u2_uk_K_r9_reg_26 (.CK( clk ) , .D( u2_uk_K_r8_26 ) , .Q( u2_uk_K_r9_26 ) , .QN( u2_uk_n1652 ) );
  DFF_X1 u2_uk_K_r9_reg_27 (.CK( clk ) , .D( u2_uk_K_r8_27 ) , .Q( u2_uk_K_r9_27 ) );
  DFF_X1 u2_uk_K_r9_reg_28 (.CK( clk ) , .D( u2_uk_K_r8_28 ) , .Q( u2_uk_K_r9_28 ) , .QN( u2_uk_n1653 ) );
  DFF_X1 u2_uk_K_r9_reg_29 (.CK( clk ) , .D( u2_uk_K_r8_29 ) , .Q( u2_uk_K_r9_29 ) , .QN( u2_uk_n1654 ) );
  DFF_X1 u2_uk_K_r9_reg_3 (.CK( clk ) , .D( u2_uk_K_r8_3 ) , .Q( u2_uk_K_r9_3 ) , .QN( u2_uk_n1633 ) );
  DFF_X1 u2_uk_K_r9_reg_30 (.CK( clk ) , .D( u2_uk_K_r8_30 ) , .Q( u2_uk_K_r9_30 ) );
  DFF_X1 u2_uk_K_r9_reg_31 (.CK( clk ) , .D( u2_uk_K_r8_31 ) , .Q( u2_uk_K_r9_31 ) );
  DFF_X1 u2_uk_K_r9_reg_32 (.CK( clk ) , .D( u2_uk_K_r8_32 ) , .Q( u2_uk_K_r9_32 ) , .QN( u2_uk_n1657 ) );
  DFF_X1 u2_uk_K_r9_reg_33 (.CK( clk ) , .D( u2_uk_K_r8_33 ) , .Q( u2_uk_K_r9_33 ) );
  DFF_X1 u2_uk_K_r9_reg_34 (.CK( clk ) , .D( u2_uk_K_r8_34 ) , .Q( u2_uk_K_r9_34 ) , .QN( u2_uk_n1658 ) );
  DFF_X1 u2_uk_K_r9_reg_35 (.CK( clk ) , .D( u2_uk_K_r8_35 ) , .Q( u2_uk_K_r9_35 ) );
  DFF_X1 u2_uk_K_r9_reg_36 (.CK( clk ) , .D( u2_uk_K_r8_36 ) , .Q( u2_uk_K_r9_36 ) , .QN( u2_uk_n1659 ) );
  DFF_X1 u2_uk_K_r9_reg_37 (.CK( clk ) , .D( u2_uk_K_r8_37 ) , .Q( u2_uk_K_r9_37 ) , .QN( u2_uk_n1660 ) );
  DFF_X1 u2_uk_K_r9_reg_38 (.CK( clk ) , .D( u2_uk_K_r8_38 ) , .Q( u2_uk_K_r9_38 ) );
  DFF_X1 u2_uk_K_r9_reg_39 (.CK( clk ) , .D( u2_uk_K_r8_39 ) , .Q( u2_uk_K_r9_39 ) , .QN( u2_uk_n1661 ) );
  DFF_X1 u2_uk_K_r9_reg_4 (.CK( clk ) , .D( u2_uk_K_r8_4 ) , .Q( u2_uk_K_r9_4 ) );
  DFF_X1 u2_uk_K_r9_reg_40 (.CK( clk ) , .D( u2_uk_K_r8_40 ) , .Q( u2_uk_K_r9_40 ) , .QN( u2_uk_n1662 ) );
  DFF_X1 u2_uk_K_r9_reg_41 (.CK( clk ) , .D( u2_uk_K_r8_41 ) , .Q( u2_uk_K_r9_41 ) , .QN( u2_uk_n1663 ) );
  DFF_X1 u2_uk_K_r9_reg_42 (.CK( clk ) , .D( u2_uk_K_r8_42 ) , .Q( u2_uk_K_r9_42 ) , .QN( u2_uk_n1664 ) );
  DFF_X1 u2_uk_K_r9_reg_43 (.CK( clk ) , .D( u2_uk_K_r8_43 ) , .Q( u2_uk_K_r9_43 ) , .QN( u2_uk_n1665 ) );
  DFF_X1 u2_uk_K_r9_reg_44 (.CK( clk ) , .D( u2_uk_K_r8_44 ) , .Q( u2_uk_K_r9_44 ) , .QN( u2_uk_n1666 ) );
  DFF_X1 u2_uk_K_r9_reg_45 (.CK( clk ) , .D( u2_uk_K_r8_45 ) , .Q( u2_uk_K_r9_45 ) );
  DFF_X1 u2_uk_K_r9_reg_46 (.CK( clk ) , .D( u2_uk_K_r8_46 ) , .Q( u2_uk_K_r9_46 ) , .QN( u2_uk_n1668 ) );
  DFF_X1 u2_uk_K_r9_reg_47 (.CK( clk ) , .D( u2_uk_K_r8_47 ) , .Q( u2_uk_K_r9_47 ) , .QN( u2_uk_n1669 ) );
  DFF_X1 u2_uk_K_r9_reg_48 (.CK( clk ) , .D( u2_uk_K_r8_48 ) , .Q( u2_uk_K_r9_48 ) );
  DFF_X1 u2_uk_K_r9_reg_49 (.CK( clk ) , .D( u2_uk_K_r8_49 ) , .Q( u2_uk_K_r9_49 ) );
  DFF_X1 u2_uk_K_r9_reg_5 (.CK( clk ) , .D( u2_uk_K_r8_5 ) , .Q( u2_uk_K_r9_5 ) );
  DFF_X1 u2_uk_K_r9_reg_50 (.CK( clk ) , .D( u2_uk_K_r8_50 ) , .Q( u2_uk_K_r9_50 ) , .QN( u2_uk_n1672 ) );
  DFF_X1 u2_uk_K_r9_reg_51 (.CK( clk ) , .D( u2_uk_K_r8_51 ) , .Q( u2_uk_K_r9_51 ) , .QN( u2_uk_n1673 ) );
  DFF_X1 u2_uk_K_r9_reg_52 (.CK( clk ) , .D( u2_uk_K_r8_52 ) , .Q( u2_uk_K_r9_52 ) , .QN( u2_uk_n1674 ) );
  DFF_X1 u2_uk_K_r9_reg_53 (.CK( clk ) , .D( u2_uk_K_r8_53 ) , .Q( u2_uk_K_r9_53 ) , .QN( u2_uk_n1675 ) );
  DFF_X1 u2_uk_K_r9_reg_54 (.CK( clk ) , .D( u2_uk_K_r8_54 ) , .Q( u2_uk_K_r9_54 ) );
  DFF_X1 u2_uk_K_r9_reg_55 (.CK( clk ) , .D( u2_uk_K_r8_55 ) , .Q( u2_uk_K_r9_55 ) , .QN( u2_uk_n1677 ) );
  DFF_X1 u2_uk_K_r9_reg_6 (.CK( clk ) , .D( u2_uk_K_r8_6 ) , .Q( u2_uk_K_r9_6 ) );
  DFF_X1 u2_uk_K_r9_reg_7 (.CK( clk ) , .D( u2_uk_K_r8_7 ) , .Q( u2_uk_K_r9_7 ) );
  DFF_X1 u2_uk_K_r9_reg_8 (.CK( clk ) , .D( u2_uk_K_r8_8 ) , .Q( u2_uk_K_r9_8 ) , .QN( u2_uk_n1634 ) );
  DFF_X1 u2_uk_K_r9_reg_9 (.CK( clk ) , .D( u2_uk_K_r8_9 ) , .Q( u2_uk_K_r9_9 ) );
  NAND2_X1 u2_uk_U1004 (.A2( decrypt ) , .A1( u2_uk_K_r10_19 ) , .ZN( u2_uk_n520 ) );
  OAI21_X1 u2_uk_U1007 (.B1( decrypt ) , .ZN( u2_K1_37 ) , .B2( u2_uk_n1144 ) , .A( u2_uk_n983 ) );
  OAI22_X1 u2_uk_U101 (.A1( decrypt ) , .ZN( u2_K9_5 ) , .B2( u2_uk_n1580 ) , .A2( u2_uk_n1586 ) , .B1( u2_uk_n191 ) );
  OAI22_X1 u2_uk_U102 (.A1( decrypt ) , .ZN( u2_K7_5 ) , .B2( u2_uk_n1457 ) , .A2( u2_uk_n1474 ) , .B1( u2_uk_n155 ) );
  NAND2_X1 u2_uk_U1020 (.A2( decrypt ) , .A1( u2_uk_K_r10_52 ) , .ZN( u2_uk_n472 ) );
  NAND2_X1 u2_uk_U1022 (.A2( decrypt ) , .A1( u2_uk_K_r4_31 ) , .ZN( u2_uk_n1069 ) );
  OAI21_X1 u2_uk_U1027 (.B1( decrypt ) , .ZN( u2_K7_31 ) , .A( u2_uk_n1087 ) , .B2( u2_uk_n1478 ) );
  OAI22_X1 u2_uk_U103 (.A1( decrypt ) , .ZN( u2_K5_5 ) , .A2( u2_uk_n1368 ) , .B2( u2_uk_n1392 ) , .B1( u2_uk_n146 ) );
  NAND2_X1 u2_uk_U1034 (.A2( decrypt ) , .A1( u2_uk_K_r13_36 ) , .ZN( u2_uk_n941 ) );
  OAI21_X1 u2_uk_U1035 (.B1( decrypt ) , .ZN( u2_K7_38 ) , .A( u2_uk_n1092 ) , .B2( u2_uk_n1469 ) );
  NAND2_X1 u2_uk_U1036 (.A2( decrypt ) , .A1( u2_uk_K_r5_8 ) , .ZN( u2_uk_n1092 ) );
  OAI21_X1 u2_uk_U1039 (.B1( decrypt ) , .ZN( u2_K4_38 ) , .A( u2_uk_n1034 ) , .B2( u2_uk_n1353 ) );
  OAI21_X1 u2_uk_U1041 (.B1( decrypt ) , .ZN( u2_K11_29 ) , .B2( u2_uk_n1634 ) , .A( u2_uk_n366 ) );
  OAI22_X1 u2_uk_U105 (.B1( decrypt ) , .ZN( u2_K1_5 ) , .A2( u2_uk_n1146 ) , .B2( u2_uk_n1150 ) , .A1( u2_uk_n147 ) );
  OAI22_X1 u2_uk_U108 (.A1( decrypt ) , .ZN( u2_K12_41 ) , .B1( u2_uk_n141 ) , .B2( u2_uk_n1705 ) , .A2( u2_uk_n1714 ) );
  AOI22_X1 u2_uk_U1085 (.B1( decrypt ) , .B2( u2_key_r_32 ) , .A2( u2_key_r_39 ) , .A1( u2_uk_n203 ) , .ZN( u2_uk_n967 ) );
  AOI22_X1 u2_uk_U1087 (.B1( decrypt ) , .A2( u2_key_r_5 ) , .B2( u2_key_r_55 ) , .A1( u2_uk_n142 ) , .ZN( u2_uk_n972 ) );
  AOI22_X1 u2_uk_U1097 (.B1( decrypt ) , .B2( u2_uk_K_r9_25 ) , .A2( u2_uk_K_r9_6 ) , .A1( u2_uk_n213 ) , .ZN( u2_uk_n313 ) );
  OAI22_X1 u2_uk_U110 (.B1( decrypt ) , .ZN( u2_K16_47 ) , .B2( u2_uk_n1188 ) , .A2( u2_uk_n1192 ) , .A1( u2_uk_n207 ) );
  AOI22_X1 u2_uk_U1105 (.B1( decrypt ) , .A2( u2_uk_K_r2_4 ) , .B2( u2_uk_K_r2_41 ) , .ZN( u2_uk_n1035 ) , .A1( u2_uk_n230 ) );
  OAI22_X1 u2_uk_U111 (.A1( decrypt ) , .ZN( u2_K13_47 ) , .B2( u2_uk_n1752 ) , .A2( u2_uk_n1762 ) , .B1( u2_uk_n202 ) );
  AOI22_X1 u2_uk_U1111 (.B1( decrypt ) , .B2( u2_uk_K_r10_23 ) , .A2( u2_uk_K_r10_28 ) , .A1( u2_uk_n220 ) , .ZN( u2_uk_n467 ) );
  AOI22_X1 u2_uk_U1115 (.B1( decrypt ) , .B2( u2_uk_K_r3_24 ) , .A2( u2_uk_K_r3_47 ) , .ZN( u2_uk_n1043 ) , .A1( u2_uk_n155 ) );
  OAI22_X1 u2_uk_U112 (.A1( decrypt ) , .ZN( u2_K12_47 ) , .B2( u2_uk_n1679 ) , .A2( u2_uk_n1706 ) , .B1( u2_uk_n222 ) );
  AOI22_X1 u2_uk_U1123 (.B1( decrypt ) , .B2( u2_uk_K_r2_13 ) , .A2( u2_uk_K_r2_33 ) , .ZN( u2_uk_n1024 ) , .A1( u2_uk_n161 ) );
  AOI22_X1 u2_uk_U1127 (.A1( decrypt ) , .B2( u2_uk_K_r3_29 ) , .A2( u2_uk_K_r3_38 ) , .ZN( u2_uk_n1049 ) , .B1( u2_uk_n163 ) );
  AOI22_X1 u2_uk_U1133 (.A1( decrypt ) , .B2( u2_uk_K_r8_17 ) , .A2( u2_uk_K_r8_39 ) , .B1( u2_uk_n191 ) , .ZN( u2_uk_n240 ) );
  AOI22_X1 u2_uk_U1135 (.A1( decrypt ) , .B2( u2_uk_K_r11_34 ) , .A2( u2_uk_K_r11_54 ) , .B1( u2_uk_n238 ) , .ZN( u2_uk_n551 ) );
  AOI22_X1 u2_uk_U1137 (.A1( decrypt ) , .B2( u2_uk_K_r6_10 ) , .A2( u2_uk_K_r6_17 ) , .ZN( u2_uk_n1100 ) , .B1( u2_uk_n188 ) );
  AOI22_X1 u2_uk_U1138 (.A1( decrypt ) , .B2( u2_uk_K_r6_21 ) , .A2( u2_uk_K_r6_28 ) , .ZN( u2_uk_n1113 ) , .B1( u2_uk_n238 ) );
  NAND2_X1 u2_uk_U1141 (.A2( decrypt ) , .A1( u2_uk_K_r14_11 ) , .ZN( u2_uk_n956 ) );
  AOI22_X1 u2_uk_U1142 (.B1( decrypt ) , .A2( u2_uk_K_r13_2 ) , .B2( u2_uk_K_r13_23 ) , .A1( u2_uk_n213 ) , .ZN( u2_uk_n944 ) );
  AOI22_X1 u2_uk_U1144 (.B1( decrypt ) , .B2( u2_uk_K_r10_39 ) , .A2( u2_uk_K_r10_48 ) , .A1( u2_uk_n209 ) , .ZN( u2_uk_n421 ) );
  AOI22_X1 u2_uk_U1148 (.A1( decrypt ) , .B2( u2_uk_K_r11_26 ) , .A2( u2_uk_K_r11_46 ) , .B1( u2_uk_n209 ) , .ZN( u2_uk_n665 ) );
  AOI22_X1 u2_uk_U1152 (.B1( decrypt ) , .B2( u2_uk_K_r7_20 ) , .A2( u2_uk_K_r7_27 ) , .ZN( u2_uk_n1130 ) , .A1( u2_uk_n161 ) );
  AOI22_X1 u2_uk_U1156 (.B1( decrypt ) , .B2( u2_uk_K_r2_26 ) , .A2( u2_uk_K_r2_46 ) , .ZN( u2_uk_n1031 ) , .A1( u2_uk_n187 ) );
  NAND2_X1 u2_uk_U119 (.A2( decrypt ) , .A1( u2_uk_K_r4_23 ) , .ZN( u2_uk_n1070 ) );
  OAI22_X1 u2_uk_U120 (.B1( decrypt ) , .ZN( u2_K5_47 ) , .B2( u2_uk_n1365 ) , .A2( u2_uk_n1389 ) , .A1( u2_uk_n213 ) );
  OAI21_X1 u2_uk_U122 (.B1( decrypt ) , .ZN( u2_K2_47 ) , .A( u2_uk_n1003 ) , .B2( u2_uk_n1241 ) );
  NAND2_X1 u2_uk_U123 (.A2( decrypt ) , .A1( u2_uk_K_r0_52 ) , .ZN( u2_uk_n1003 ) );
  OAI22_X1 u2_uk_U124 (.A1( decrypt ) , .ZN( u2_K1_15 ) , .B2( u2_uk_n1161 ) , .A2( u2_uk_n1167 ) , .B1( u2_uk_n209 ) );
  NAND2_X1 u2_uk_U127 (.A2( decrypt ) , .A1( u2_uk_K_r3_34 ) , .ZN( u2_uk_n1042 ) );
  AOI22_X1 u2_uk_U129 (.B1( decrypt ) , .B2( u2_uk_K_r11_11 ) , .A2( u2_uk_K_r11_48 ) , .A1( u2_uk_n141 ) , .ZN( u2_uk_n586 ) );
  OAI22_X1 u2_uk_U133 (.B1( decrypt ) , .ZN( u2_K3_15 ) , .A2( u2_uk_n1282 ) , .A1( u2_uk_n129 ) , .B2( u2_uk_n1317 ) );
  NAND2_X1 u2_uk_U138 (.A2( decrypt ) , .A1( u2_uk_K_r4_48 ) , .ZN( u2_uk_n1061 ) );
  NAND2_X1 u2_uk_U140 (.A2( decrypt ) , .A1( u2_uk_K_r0_19 ) , .ZN( u2_uk_n994 ) );
  OAI22_X1 u2_uk_U141 (.B1( decrypt ) , .ZN( u2_K1_19 ) , .B2( u2_uk_n1145 ) , .A2( u2_uk_n1185 ) , .A1( u2_uk_n217 ) );
  OAI22_X1 u2_uk_U143 (.A1( decrypt ) , .ZN( u2_K10_15 ) , .A2( u2_uk_n1592 ) , .B2( u2_uk_n1629 ) , .B1( u2_uk_n182 ) );
  NAND2_X1 u2_uk_U155 (.A2( decrypt ) , .A1( u2_uk_K_r1_33 ) , .ZN( u2_uk_n1007 ) );
  AOI22_X1 u2_uk_U165 (.A1( decrypt ) , .B2( u2_uk_K_r10_23 ) , .A2( u2_uk_K_r10_42 ) , .B1( u2_uk_n191 ) , .ZN( u2_uk_n456 ) );
  OAI22_X1 u2_uk_U166 (.A1( decrypt ) , .ZN( u2_K10_30 ) , .B1( u2_uk_n146 ) , .B2( u2_uk_n1598 ) , .A2( u2_uk_n1626 ) );
  OAI22_X1 u2_uk_U167 (.A1( decrypt ) , .ZN( u2_K12_24 ) , .B1( u2_uk_n155 ) , .B2( u2_uk_n1686 ) , .A2( u2_uk_n1715 ) );
  NAND2_X1 u2_uk_U169 (.A2( decrypt ) , .A1( u2_key_r_18 ) , .ZN( u2_uk_n970 ) );
  OAI22_X1 u2_uk_U175 (.A1( decrypt ) , .ZN( u2_K13_14 ) , .B1( u2_uk_n141 ) , .B2( u2_uk_n1726 ) , .A2( u2_uk_n1750 ) );
  AOI22_X1 u2_uk_U178 (.A1( decrypt ) , .B2( u2_uk_K_r9_12 ) , .A2( u2_uk_K_r9_6 ) , .B1( u2_uk_n188 ) , .ZN( u2_uk_n319 ) );
  NAND2_X1 u2_uk_U182 (.A2( decrypt ) , .A1( u2_uk_K_r7_34 ) , .ZN( u2_uk_n1121 ) );
  OAI22_X1 u2_uk_U183 (.A1( decrypt ) , .ZN( u2_K6_14 ) , .A2( u2_uk_n1410 ) , .B2( u2_uk_n1416 ) , .B1( u2_uk_n222 ) );
  OAI22_X1 u2_uk_U186 (.A1( decrypt ) , .ZN( u2_K1_24 ) , .B2( u2_uk_n1150 ) , .A2( u2_uk_n1155 ) , .B1( u2_uk_n238 ) );
  NAND2_X1 u2_uk_U201 (.A2( decrypt ) , .A1( u2_key_r_45 ) , .ZN( u2_uk_n979 ) );
  NAND2_X1 u2_uk_U203 (.A2( decrypt ) , .A1( u2_uk_K_r7_29 ) , .ZN( u2_uk_n1131 ) );
  OAI22_X1 u2_uk_U213 (.A1( decrypt ) , .ZN( u2_K16_31 ) , .A2( u2_uk_n1192 ) , .B2( u2_uk_n1195 ) , .B1( u2_uk_n191 ) );
  OAI22_X1 u2_uk_U214 (.A1( decrypt ) , .ZN( u2_K8_31 ) , .B2( u2_uk_n1499 ) , .A2( u2_uk_n1537 ) , .B1( u2_uk_n208 ) );
  AOI22_X1 u2_uk_U218 (.B1( decrypt ) , .B2( u2_uk_K_r9_22 ) , .A2( u2_uk_K_r9_30 ) , .A1( u2_uk_n203 ) , .ZN( u2_uk_n373 ) );
  AOI22_X1 u2_uk_U221 (.B1( decrypt ) , .B2( u2_uk_K_r9_30 ) , .A2( u2_uk_K_r9_7 ) , .A1( u2_uk_n207 ) , .ZN( u2_uk_n379 ) );
  OAI22_X1 u2_uk_U224 (.B1( decrypt ) , .ZN( u2_K13_31 ) , .A1( u2_uk_n146 ) , .B2( u2_uk_n1742 ) , .A2( u2_uk_n1760 ) );
  OAI21_X1 u2_uk_U229 (.B1( decrypt ) , .ZN( u2_K5_31 ) , .A( u2_uk_n1047 ) , .B2( u2_uk_n1371 ) );
  NAND2_X1 u2_uk_U230 (.A2( decrypt ) , .A1( u2_uk_K_r3_44 ) , .ZN( u2_uk_n1047 ) );
  OAI22_X1 u2_uk_U231 (.B1( decrypt ) , .ZN( u2_K15_31 ) , .B2( u2_uk_n1813 ) , .A2( u2_uk_n1830 ) , .A1( u2_uk_n207 ) );
  NAND2_X1 u2_uk_U233 (.A2( decrypt ) , .A1( u2_key_r_15 ) , .ZN( u2_uk_n984 ) );
  OAI22_X1 u2_uk_U237 (.A1( decrypt ) , .ZN( u2_K15_39 ) , .A2( u2_uk_n1818 ) , .B2( u2_uk_n1836 ) , .B1( u2_uk_n188 ) );
  OAI22_X1 u2_uk_U238 (.A1( decrypt ) , .ZN( u2_K14_39 ) , .B1( u2_uk_n142 ) , .B2( u2_uk_n1802 ) , .A2( u2_uk_n1806 ) );
  OAI21_X1 u2_uk_U243 (.B1( decrypt ) , .ZN( u2_K16_44 ) , .B2( u2_uk_n1216 ) , .A( u2_uk_n964 ) );
  NAND2_X1 u2_uk_U244 (.A2( decrypt ) , .A1( u2_uk_K_r14_43 ) , .ZN( u2_uk_n964 ) );
  OAI22_X1 u2_uk_U245 (.B1( decrypt ) , .ZN( u2_K5_44 ) , .B2( u2_uk_n1389 ) , .A2( u2_uk_n1395 ) , .A1( u2_uk_n207 ) );
  OAI22_X1 u2_uk_U246 (.B1( decrypt ) , .ZN( u2_K5_48 ) , .B2( u2_uk_n1377 ) , .A2( u2_uk_n1384 ) , .A1( u2_uk_n213 ) );
  NAND2_X1 u2_uk_U251 (.A2( decrypt ) , .A1( u2_uk_K_r13_35 ) , .ZN( u2_uk_n945 ) );
  OAI22_X1 u2_uk_U253 (.B1( decrypt ) , .ZN( u2_K13_44 ) , .B2( u2_uk_n1724 ) , .A2( u2_uk_n1739 ) , .A1( u2_uk_n220 ) );
  NAND2_X1 u2_uk_U255 (.A2( decrypt ) , .A1( u2_uk_K_r11_8 ) , .ZN( u2_uk_n677 ) );
  AOI22_X1 u2_uk_U257 (.B1( decrypt ) , .B2( u2_uk_K_r10_37 ) , .A2( u2_uk_K_r10_42 ) , .A1( u2_uk_n230 ) , .ZN( u2_uk_n504 ) );
  OAI22_X1 u2_uk_U260 (.B1( decrypt ) , .ZN( u2_K10_44 ) , .B2( u2_uk_n1597 ) , .A2( u2_uk_n1617 ) , .A1( u2_uk_n188 ) );
  AOI22_X1 u2_uk_U263 (.A1( decrypt ) , .B2( u2_uk_K_r7_16 ) , .A2( u2_uk_K_r7_9 ) , .ZN( u2_uk_n1140 ) , .B1( u2_uk_n231 ) );
  OAI22_X1 u2_uk_U268 (.A1( decrypt ) , .ZN( u2_K7_48 ) , .B2( u2_uk_n1471 ) , .A2( u2_uk_n1491 ) , .B1( u2_uk_n188 ) );
  OAI22_X1 u2_uk_U274 (.A1( decrypt ) , .ZN( u2_K3_48 ) , .B2( u2_uk_n1277 ) , .A2( u2_uk_n1312 ) , .B1( u2_uk_n222 ) );
  OAI22_X1 u2_uk_U275 (.A1( decrypt ) , .ZN( u2_K2_44 ) , .B2( u2_uk_n1251 ) , .A2( u2_uk_n1273 ) , .B1( u2_uk_n208 ) );
  OAI22_X1 u2_uk_U276 (.B1( decrypt ) , .ZN( u2_K16_6 ) , .B2( u2_uk_n1214 ) , .A2( u2_uk_n1219 ) , .A1( u2_uk_n203 ) );
  OAI22_X1 u2_uk_U278 (.B1( decrypt ) , .ZN( u2_K14_6 ) , .A1( u2_uk_n146 ) , .A2( u2_uk_n1773 ) , .B2( u2_uk_n1780 ) );
  OAI22_X1 u2_uk_U279 (.B1( decrypt ) , .ZN( u2_K10_6 ) , .A1( u2_uk_n147 ) , .A2( u2_uk_n1591 ) , .B2( u2_uk_n1619 ) );
  NAND2_X1 u2_uk_U282 (.A2( decrypt ) , .A1( u2_uk_K_r4_18 ) , .ZN( u2_uk_n1073 ) );
  OAI22_X1 u2_uk_U287 (.B1( decrypt ) , .ZN( u2_K12_8 ) , .A1( u2_uk_n129 ) , .B2( u2_uk_n1701 ) , .A2( u2_uk_n1722 ) );
  OAI22_X1 u2_uk_U288 (.B1( decrypt ) , .ZN( u2_K8_8 ) , .B2( u2_uk_n1528 ) , .A2( u2_uk_n1534 ) , .A1( u2_uk_n203 ) );
  AOI22_X1 u2_uk_U290 (.A1( decrypt ) , .B2( u2_uk_K_r5_26 ) , .A2( u2_uk_K_r5_4 ) , .ZN( u2_uk_n1096 ) , .B1( u2_uk_n147 ) );
  OAI22_X1 u2_uk_U291 (.A1( decrypt ) , .ZN( u2_K5_8 ) , .B2( u2_uk_n1385 ) , .A2( u2_uk_n1407 ) , .B1( u2_uk_n222 ) );
  AOI22_X1 u2_uk_U293 (.A1( decrypt ) , .B2( u2_uk_K_r2_41 ) , .A2( u2_uk_K_r2_46 ) , .ZN( u2_uk_n1040 ) , .B1( u2_uk_n188 ) );
  OAI22_X1 u2_uk_U297 (.A1( decrypt ) , .ZN( u2_K7_26 ) , .B2( u2_uk_n1470 ) , .A2( u2_uk_n1490 ) , .B1( u2_uk_n209 ) );
  OAI22_X1 u2_uk_U300 (.B1( decrypt ) , .ZN( u2_K16_8 ) , .A2( u2_uk_n1191 ) , .B2( u2_uk_n1204 ) , .A1( u2_uk_n230 ) );
  AOI22_X1 u2_uk_U302 (.A1( decrypt ) , .B2( u2_uk_K_r7_15 ) , .A2( u2_uk_K_r7_8 ) , .ZN( u2_uk_n1128 ) , .B1( u2_uk_n238 ) );
  AOI22_X1 u2_uk_U304 (.B1( decrypt ) , .B2( u2_uk_K_r2_16 ) , .A2( u2_uk_K_r2_7 ) , .ZN( u2_uk_n1028 ) , .A1( u2_uk_n163 ) );
  AOI22_X1 u2_uk_U306 (.B1( decrypt ) , .B2( u2_uk_K_r13_38 ) , .A2( u2_uk_K_r13_44 ) , .A1( u2_uk_n203 ) , .ZN( u2_uk_n939 ) );
  NAND2_X1 u2_uk_U310 (.A2( decrypt ) , .A1( u2_uk_K_r9_35 ) , .ZN( u2_uk_n363 ) );
  OAI21_X1 u2_uk_U311 (.B1( decrypt ) , .ZN( u2_K13_26 ) , .B2( u2_uk_n1735 ) , .A( u2_uk_n656 ) );
  OAI22_X1 u2_uk_U313 (.B1( decrypt ) , .ZN( u2_K5_26 ) , .A2( u2_uk_n1366 ) , .B2( u2_uk_n1376 ) , .A1( u2_uk_n213 ) );
  OAI22_X1 u2_uk_U315 (.A1( decrypt ) , .ZN( u2_K16_26 ) , .B2( u2_uk_n1211 ) , .A2( u2_uk_n1225 ) , .B1( u2_uk_n223 ) );
  OAI22_X1 u2_uk_U317 (.A1( decrypt ) , .ZN( u2_K12_26 ) , .B1( u2_uk_n146 ) , .A2( u2_uk_n1680 ) , .B2( u2_uk_n1690 ) );
  OAI22_X1 u2_uk_U318 (.B1( decrypt ) , .ZN( u2_K10_26 ) , .B2( u2_uk_n1609 ) , .A2( u2_uk_n1625 ) , .A1( u2_uk_n202 ) );
  OAI22_X1 u2_uk_U319 (.A1( decrypt ) , .ZN( u2_K8_26 ) , .A2( u2_uk_n1503 ) , .B2( u2_uk_n1510 ) , .B1( u2_uk_n220 ) );
  OAI22_X1 u2_uk_U323 (.B1( decrypt ) , .ZN( u2_K13_46 ) , .A1( u2_uk_n145 ) , .B2( u2_uk_n1733 ) , .A2( u2_uk_n1745 ) );
  OAI22_X1 u2_uk_U324 (.B1( decrypt ) , .ZN( u2_K12_46 ) , .B2( u2_uk_n1678 ) , .A2( u2_uk_n1718 ) , .A1( u2_uk_n203 ) );
  OAI22_X1 u2_uk_U328 (.A1( decrypt ) , .ZN( u2_K2_46 ) , .A2( u2_uk_n1236 ) , .B2( u2_uk_n1263 ) , .B1( u2_uk_n163 ) );
  OAI21_X1 u2_uk_U329 (.B1( decrypt ) , .ZN( u2_K1_46 ) , .B2( u2_uk_n1143 ) , .A( u2_uk_n988 ) );
  OAI22_X1 u2_uk_U333 (.A1( decrypt ) , .ZN( u2_K11_4 ) , .B2( u2_uk_n1663 ) , .A2( u2_uk_n1669 ) , .B1( u2_uk_n214 ) );
  AOI22_X1 u2_uk_U335 (.A1( decrypt ) , .B2( u2_uk_K_r9_45 ) , .A2( u2_uk_K_r9_9 ) , .B1( u2_uk_n188 ) , .ZN( u2_uk_n385 ) );
  OAI22_X1 u2_uk_U340 (.B1( decrypt ) , .ZN( u2_K10_4 ) , .B2( u2_uk_n1612 ) , .A2( u2_uk_n1631 ) , .A1( u2_uk_n217 ) );
  OAI22_X1 u2_uk_U341 (.A1( decrypt ) , .ZN( u2_K7_4 ) , .B2( u2_uk_n1474 ) , .A2( u2_uk_n1497 ) , .B1( u2_uk_n214 ) );
  OAI22_X1 u2_uk_U346 (.B1( decrypt ) , .ZN( u2_K1_40 ) , .B2( u2_uk_n1142 ) , .A2( u2_uk_n1183 ) , .A1( u2_uk_n187 ) );
  OAI22_X1 u2_uk_U347 (.A1( decrypt ) , .ZN( u2_K6_40 ) , .A2( u2_uk_n1412 ) , .B2( u2_uk_n1420 ) , .B1( u2_uk_n146 ) );
  AOI22_X1 u2_uk_U349 (.A1( decrypt ) , .B2( u2_uk_K_r5_23 ) , .A2( u2_uk_K_r5_31 ) , .ZN( u2_uk_n1094 ) , .B1( u2_uk_n148 ) );
  NAND2_X1 u2_uk_U353 (.A2( decrypt ) , .A1( u2_uk_K_r12_21 ) , .ZN( u2_uk_n702 ) );
  OAI22_X1 u2_uk_U356 (.A1( decrypt ) , .ZN( u2_K13_40 ) , .B2( u2_uk_n1744 ) , .A2( u2_uk_n1754 ) , .B1( u2_uk_n208 ) );
  OAI22_X1 u2_uk_U361 (.A1( decrypt ) , .ZN( u2_K2_40 ) , .A2( u2_uk_n1235 ) , .B2( u2_uk_n1266 ) , .B1( u2_uk_n163 ) );
  NAND2_X1 u2_uk_U363 (.A2( decrypt ) , .A1( u2_uk_K_r13_31 ) , .ZN( u2_uk_n942 ) );
  OAI22_X1 u2_uk_U366 (.A1( decrypt ) , .ZN( u2_K1_28 ) , .B2( u2_uk_n1143 ) , .A2( u2_uk_n1148 ) , .B1( u2_uk_n214 ) );
  NAND2_X1 u2_uk_U369 (.A2( decrypt ) , .A1( u2_uk_K_r14_8 ) , .ZN( u2_uk_n954 ) );
  OAI22_X1 u2_uk_U370 (.A1( decrypt ) , .ZN( u2_K14_28 ) , .B1( u2_uk_n141 ) , .B2( u2_uk_n1791 ) , .A2( u2_uk_n1797 ) );
  OAI22_X1 u2_uk_U376 (.A1( decrypt ) , .ZN( u2_K15_28 ) , .B2( u2_uk_n1825 ) , .A2( u2_uk_n1853 ) , .B1( u2_uk_n213 ) );
  OAI22_X1 u2_uk_U379 (.A1( decrypt ) , .ZN( u2_K9_28 ) , .B2( u2_uk_n1577 ) , .A2( u2_uk_n1584 ) , .B1( u2_uk_n217 ) );
  OAI22_X1 u2_uk_U381 (.B1( decrypt ) , .ZN( u2_K5_28 ) , .B2( u2_uk_n1366 ) , .A2( u2_uk_n1370 ) , .A1( u2_uk_n213 ) );
  OAI22_X1 u2_uk_U382 (.B1( decrypt ) , .ZN( u2_K15_1 ) , .B2( u2_uk_n1838 ) , .A2( u2_uk_n1857 ) , .A1( u2_uk_n213 ) );
  NAND2_X1 u2_uk_U385 (.A2( decrypt ) , .A1( u2_uk_K_r8_10 ) , .ZN( u2_uk_n251 ) );
  OAI22_X1 u2_uk_U386 (.A1( decrypt ) , .ZN( u2_K6_1 ) , .B2( u2_uk_n1432 ) , .A2( u2_uk_n1448 ) , .B1( u2_uk_n146 ) );
  OAI22_X1 u2_uk_U387 (.B1( decrypt ) , .ZN( u2_K5_1 ) , .B2( u2_uk_n1392 ) , .A2( u2_uk_n1399 ) , .A1( u2_uk_n203 ) );
  OAI22_X1 u2_uk_U394 (.A1( decrypt ) , .ZN( u2_K1_9 ) , .B2( u2_uk_n1179 ) , .A2( u2_uk_n1185 ) , .B1( u2_uk_n145 ) );
  NAND2_X1 u2_uk_U401 (.A2( decrypt ) , .A1( u2_uk_K_r5_32 ) , .ZN( u2_uk_n1077 ) );
  OAI22_X1 u2_uk_U402 (.B1( decrypt ) , .ZN( u2_K6_16 ) , .B2( u2_uk_n1436 ) , .A2( u2_uk_n1442 ) , .A1( u2_uk_n148 ) );
  OAI21_X1 u2_uk_U404 (.B1( decrypt ) , .ZN( u2_K3_16 ) , .A( u2_uk_n1006 ) , .B2( u2_uk_n1318 ) );
  NAND2_X1 u2_uk_U405 (.A2( decrypt ) , .A1( u2_uk_K_r1_6 ) , .ZN( u2_uk_n1006 ) );
  OAI22_X1 u2_uk_U406 (.A1( decrypt ) , .ZN( u2_K1_16 ) , .B2( u2_uk_n1162 ) , .A2( u2_uk_n1168 ) , .B1( u2_uk_n214 ) );
  NAND2_X1 u2_uk_U408 (.A2( decrypt ) , .A1( u2_uk_K_r13_4 ) , .ZN( u2_uk_n947 ) );
  NAND2_X1 u2_uk_U410 (.A2( decrypt ) , .A1( u2_uk_K_r12_18 ) , .ZN( u2_uk_n933 ) );
  OAI22_X1 u2_uk_U413 (.A1( decrypt ) , .ZN( u2_K11_9 ) , .B2( u2_uk_n1633 ) , .A2( u2_uk_n1663 ) , .B1( u2_uk_n188 ) );
  AOI22_X1 u2_uk_U417 (.A1( decrypt ) , .B2( u2_uk_K_r8_28 ) , .A2( u2_uk_K_r8_52 ) , .B1( u2_uk_n147 ) , .ZN( u2_uk_n299 ) );
  AOI22_X1 u2_uk_U423 (.A2( decrypt ) , .B2( u2_uk_K_r7_13 ) , .A1( u2_uk_K_r7_6 ) , .ZN( u2_uk_n1141 ) , .B1( u2_uk_n217 ) );
  AOI22_X1 u2_uk_U425 (.A1( decrypt ) , .B2( u2_uk_K_r4_3 ) , .A2( u2_uk_K_r4_41 ) , .ZN( u2_uk_n1074 ) , .B1( u2_uk_n155 ) );
  OAI22_X1 u2_uk_U427 (.B1( decrypt ) , .ZN( u2_K5_9 ) , .B2( u2_uk_n1397 ) , .A2( u2_uk_n1407 ) , .A1( u2_uk_n213 ) );
  OAI22_X1 u2_uk_U432 (.A1( decrypt ) , .ZN( u2_K2_1 ) , .B2( u2_uk_n1254 ) , .A2( u2_uk_n1275 ) , .B1( u2_uk_n145 ) );
  OAI22_X1 u2_uk_U433 (.B1( decrypt ) , .ZN( u2_K16_9 ) , .B2( u2_uk_n1221 ) , .A2( u2_uk_n1228 ) , .A1( u2_uk_n222 ) );
  OAI22_X1 u2_uk_U435 (.B1( decrypt ) , .ZN( u2_K15_16 ) , .A1( u2_uk_n145 ) , .B2( u2_uk_n1829 ) , .A2( u2_uk_n1844 ) );
  OAI22_X1 u2_uk_U436 (.B1( decrypt ) , .ZN( u2_K5_16 ) , .A2( u2_uk_n1367 ) , .B2( u2_uk_n1380 ) , .A1( u2_uk_n147 ) );
  OAI22_X1 u2_uk_U437 (.A1( decrypt ) , .ZN( u2_K2_16 ) , .B2( u2_uk_n1244 ) , .A2( u2_uk_n1262 ) , .B1( u2_uk_n145 ) );
  OAI22_X1 u2_uk_U443 (.A1( decrypt ) , .ZN( u2_K7_33 ) , .B1( u2_uk_n129 ) , .B2( u2_uk_n1464 ) , .A2( u2_uk_n1484 ) );
  AOI22_X1 u2_uk_U445 (.B1( decrypt ) , .B2( u2_uk_K_r7_1 ) , .A2( u2_uk_K_r7_8 ) , .ZN( u2_uk_n1132 ) , .A1( u2_uk_n207 ) );
  NAND2_X1 u2_uk_U451 (.A2( decrypt ) , .A1( u2_uk_K_r10_14 ) , .ZN( u2_uk_n468 ) );
  OAI22_X1 u2_uk_U458 (.B1( decrypt ) , .ZN( u2_K4_33 ) , .B2( u2_uk_n1319 ) , .A2( u2_uk_n1326 ) , .A1( u2_uk_n182 ) );
  OAI22_X1 u2_uk_U462 (.B1( decrypt ) , .ZN( u2_K13_37 ) , .B2( u2_uk_n1734 ) , .A2( u2_uk_n1746 ) , .A1( u2_uk_n220 ) );
  OAI22_X1 u2_uk_U463 (.B1( decrypt ) , .ZN( u2_K12_37 ) , .B2( u2_uk_n1679 ) , .A2( u2_uk_n1719 ) , .A1( u2_uk_n207 ) );
  NAND2_X1 u2_uk_U465 (.A2( decrypt ) , .A1( u2_uk_K_r9_38 ) , .ZN( u2_uk_n377 ) );
  NAND2_X1 u2_uk_U467 (.A2( decrypt ) , .A1( u2_uk_K_r7_7 ) , .ZN( u2_uk_n1134 ) );
  OAI21_X1 u2_uk_U473 (.B1( decrypt ) , .ZN( u2_K10_36 ) , .B2( u2_uk_n1589 ) , .A( u2_uk_n298 ) );
  NAND2_X1 u2_uk_U476 (.A2( decrypt ) , .A1( u2_uk_K_r12_44 ) , .ZN( u2_uk_n689 ) );
  OAI22_X1 u2_uk_U480 (.A1( decrypt ) , .ZN( u2_K15_29 ) , .A2( u2_uk_n1819 ) , .B2( u2_uk_n1837 ) , .B1( u2_uk_n222 ) );
  AOI22_X1 u2_uk_U482 (.A1( decrypt ) , .B2( u2_uk_K_r14_16 ) , .A2( u2_uk_K_r14_23 ) , .B1( u2_uk_n214 ) , .ZN( u2_uk_n955 ) );
  OAI22_X1 u2_uk_U488 (.B1( decrypt ) , .ZN( u2_K12_29 ) , .B2( u2_uk_n1691 ) , .A2( u2_uk_n1714 ) , .A1( u2_uk_n207 ) );
  OAI22_X1 u2_uk_U490 (.A1( decrypt ) , .ZN( u2_K9_29 ) , .B2( u2_uk_n1565 ) , .A2( u2_uk_n1569 ) , .B1( u2_uk_n163 ) );
  AOI22_X1 u2_uk_U492 (.A1( decrypt ) , .B2( u2_uk_K_r6_28 ) , .A2( u2_uk_K_r6_35 ) , .ZN( u2_uk_n1104 ) , .B1( u2_uk_n188 ) );
  OAI22_X1 u2_uk_U495 (.A1( decrypt ) , .ZN( u2_K15_2 ) , .B2( u2_uk_n1828 ) , .A2( u2_uk_n1857 ) , .B1( u2_uk_n223 ) );
  NAND2_X1 u2_uk_U500 (.A2( decrypt ) , .A1( u2_uk_K_r6_27 ) , .ZN( u2_uk_n1105 ) );
  NAND2_X1 u2_uk_U506 (.A2( decrypt ) , .A1( u2_uk_K_r7_53 ) , .ZN( u2_uk_n1119 ) );
  INV_X1 u2_uk_U51 (.A( decrypt ) , .ZN( u2_uk_n238 ) );
  OAI22_X1 u2_uk_U511 (.A1( decrypt ) , .ZN( u2_K10_17 ) , .B2( u2_uk_n1596 ) , .A2( u2_uk_n1624 ) , .B1( u2_uk_n187 ) );
  OAI22_X1 u2_uk_U522 (.A1( decrypt ) , .ZN( u2_K14_12 ) , .B2( u2_uk_n1801 ) , .A2( u2_uk_n1805 ) , .B1( u2_uk_n223 ) );
  NAND2_X1 u2_uk_U524 (.A2( decrypt ) , .A1( u2_uk_K_r10_11 ) , .ZN( u2_uk_n408 ) );
  OAI22_X1 u2_uk_U538 (.A1( decrypt ) , .ZN( u2_K9_36 ) , .B2( u2_uk_n1569 ) , .A2( u2_uk_n1575 ) , .B1( u2_uk_n230 ) );
  OAI22_X1 u2_uk_U540 (.A1( decrypt ) , .ZN( u2_K14_17 ) , .B1( u2_uk_n141 ) , .B2( u2_uk_n1780 ) , .A2( u2_uk_n1804 ) );
  OAI22_X1 u2_uk_U541 (.A1( decrypt ) , .ZN( u2_K5_17 ) , .B2( u2_uk_n1374 ) , .A2( u2_uk_n1394 ) , .B1( u2_uk_n148 ) );
  AOI22_X1 u2_uk_U543 (.A1( decrypt ) , .B2( u2_uk_K_r10_18 ) , .A2( u2_uk_K_r10_41 ) , .B1( u2_uk_n217 ) , .ZN( u2_uk_n415 ) );
  OAI22_X1 u2_uk_U552 (.A1( decrypt ) , .ZN( u2_K2_36 ) , .B2( u2_uk_n1242 ) , .A2( u2_uk_n1258 ) , .B1( u2_uk_n223 ) );
  OAI22_X1 u2_uk_U555 (.A1( decrypt ) , .ZN( u2_K11_38 ) , .B1( u2_uk_n147 ) , .B2( u2_uk_n1640 ) , .A2( u2_uk_n1648 ) );
  OAI22_X1 u2_uk_U556 (.A1( decrypt ) , .ZN( u2_K9_38 ) , .B2( u2_uk_n1575 ) , .A2( u2_uk_n1582 ) , .B1( u2_uk_n188 ) );
  AOI22_X1 u2_uk_U560 (.A1( decrypt ) , .B2( u2_uk_K_r9_15 ) , .A2( u2_uk_K_r9_7 ) , .B1( u2_uk_n162 ) , .ZN( u2_uk_n376 ) );
  AOI22_X1 u2_uk_U565 (.A1( decrypt ) , .B2( u2_uk_K_r13_23 ) , .A2( u2_uk_K_r13_44 ) , .B1( u2_uk_n163 ) , .ZN( u2_uk_n943 ) );
  AOI22_X1 u2_uk_U57 (.A1( decrypt ) , .B2( u2_uk_K_r6_14 ) , .A2( u2_uk_K_r6_21 ) , .ZN( u2_uk_n1107 ) , .B1( u2_uk_n209 ) );
  OAI22_X1 u2_uk_U570 (.B1( decrypt ) , .ZN( u2_K5_38 ) , .B2( u2_uk_n1364 ) , .A2( u2_uk_n1388 ) , .A1( u2_uk_n213 ) );
  OAI22_X1 u2_uk_U573 (.A1( decrypt ) , .ZN( u2_K14_10 ) , .B2( u2_uk_n1779 ) , .A2( u2_uk_n1784 ) , .B1( u2_uk_n230 ) );
  OAI22_X1 u2_uk_U576 (.A1( decrypt ) , .ZN( u2_K10_10 ) , .B1( u2_uk_n155 ) , .B2( u2_uk_n1595 ) , .A2( u2_uk_n1623 ) );
  OAI22_X1 u2_uk_U577 (.A1( decrypt ) , .ZN( u2_K5_10 ) , .B2( u2_uk_n1373 ) , .A2( u2_uk_n1393 ) , .B1( u2_uk_n162 ) );
  OAI22_X1 u2_uk_U586 (.A1( decrypt ) , .ZN( u2_K12_22 ) , .B1( u2_uk_n141 ) , .B2( u2_uk_n1692 ) , .A2( u2_uk_n1702 ) );
  AOI22_X1 u2_uk_U59 (.A1( decrypt ) , .B2( u2_uk_K_r5_0 ) , .A2( u2_uk_K_r5_35 ) , .ZN( u2_uk_n1089 ) , .B1( u2_uk_n217 ) );
  AOI22_X1 u2_uk_U594 (.B1( decrypt ) , .B2( u2_uk_K_r8_27 ) , .A2( u2_uk_K_r8_5 ) , .A1( u2_uk_n220 ) , .ZN( u2_uk_n257 ) );
  NAND2_X1 u2_uk_U599 (.A2( decrypt ) , .A1( u2_uk_K_r5_5 ) , .ZN( u2_uk_n1081 ) );
  OAI22_X1 u2_uk_U60 (.A1( decrypt ) , .ZN( u2_K15_34 ) , .B1( u2_uk_n141 ) , .B2( u2_uk_n1826 ) , .A2( u2_uk_n1854 ) );
  AOI22_X1 u2_uk_U601 (.A1( decrypt ) , .B2( u2_uk_K_r3_24 ) , .A2( u2_uk_K_r3_33 ) , .ZN( u2_uk_n1044 ) , .B1( u2_uk_n214 ) );
  OAI21_X1 u2_uk_U607 (.B1( decrypt ) , .ZN( u2_K7_35 ) , .A( u2_uk_n1090 ) , .B2( u2_uk_n1452 ) );
  OAI22_X1 u2_uk_U609 (.B1( decrypt ) , .ZN( u2_K15_35 ) , .B2( u2_uk_n1830 ) , .A2( u2_uk_n1845 ) , .A1( u2_uk_n188 ) );
  OAI22_X1 u2_uk_U619 (.B1( decrypt ) , .ZN( u2_K4_35 ) , .B2( u2_uk_n1331 ) , .A2( u2_uk_n1360 ) , .A1( u2_uk_n164 ) );
  OAI22_X1 u2_uk_U620 (.A1( decrypt ) , .ZN( u2_K2_35 ) , .B2( u2_uk_n1245 ) , .A2( u2_uk_n1263 ) , .B1( u2_uk_n164 ) );
  NAND2_X1 u2_uk_U624 (.A2( decrypt ) , .A1( u2_uk_K_r14_39 ) , .ZN( u2_uk_n948 ) );
  OAI22_X1 u2_uk_U628 (.B1( decrypt ) , .ZN( u2_K14_11 ) , .A1( u2_uk_n142 ) , .A2( u2_uk_n1771 ) , .B2( u2_uk_n1778 ) );
  OAI22_X1 u2_uk_U629 (.A1( decrypt ) , .ZN( u2_K11_11 ) , .B1( u2_uk_n145 ) , .B2( u2_uk_n1646 ) , .A2( u2_uk_n1652 ) );
  OAI22_X1 u2_uk_U63 (.A1( decrypt ) , .ZN( u2_K12_34 ) , .B1( u2_uk_n142 ) , .A2( u2_uk_n1685 ) , .B2( u2_uk_n1700 ) );
  AOI22_X1 u2_uk_U631 (.B1( decrypt ) , .B2( u2_uk_K_r11_17 ) , .A2( u2_uk_K_r11_54 ) , .A1( u2_uk_n231 ) , .ZN( u2_uk_n526 ) );
  OAI22_X1 u2_uk_U632 (.B1( decrypt ) , .ZN( u2_K10_11 ) , .B2( u2_uk_n1596 ) , .A2( u2_uk_n1613 ) , .A1( u2_uk_n187 ) );
  NAND2_X1 u2_uk_U634 (.A2( decrypt ) , .A1( u2_uk_K_r6_55 ) , .ZN( u2_uk_n1097 ) );
  OAI22_X1 u2_uk_U637 (.B1( decrypt ) , .ZN( u2_K6_11 ) , .B2( u2_uk_n1423 ) , .A2( u2_uk_n1427 ) , .A1( u2_uk_n163 ) );
  OAI22_X1 u2_uk_U638 (.A1( decrypt ) , .ZN( u2_K5_11 ) , .A2( u2_uk_n1369 ) , .B2( u2_uk_n1393 ) , .B1( u2_uk_n147 ) );
  OAI21_X1 u2_uk_U64 (.B1( decrypt ) , .ZN( u2_K6_34 ) , .A( u2_uk_n1067 ) , .B2( u2_uk_n1441 ) );
  OAI21_X1 u2_uk_U642 (.B1( decrypt ) , .ZN( u2_K4_6 ) , .A( u2_uk_n1039 ) , .B2( u2_uk_n1335 ) );
  OAI22_X1 u2_uk_U649 (.A1( decrypt ) , .ZN( u2_K1_45 ) , .B2( u2_uk_n1171 ) , .A2( u2_uk_n1178 ) , .B1( u2_uk_n230 ) );
  NAND2_X1 u2_uk_U65 (.A2( decrypt ) , .A1( u2_uk_K_r4_49 ) , .ZN( u2_uk_n1067 ) );
  NAND2_X1 u2_uk_U654 (.A2( decrypt ) , .A1( u2_uk_K_r2_29 ) , .ZN( u2_uk_n1036 ) );
  OAI22_X1 u2_uk_U655 (.B1( decrypt ) , .ZN( u2_K3_43 ) , .B2( u2_uk_n1304 ) , .A2( u2_uk_n1308 ) , .A1( u2_uk_n202 ) );
  OAI21_X1 u2_uk_U656 (.B1( decrypt ) , .ZN( u2_K2_43 ) , .A( u2_uk_n1002 ) , .B2( u2_uk_n1246 ) );
  NAND2_X1 u2_uk_U657 (.A2( decrypt ) , .A1( u2_uk_K_r0_2 ) , .ZN( u2_uk_n1002 ) );
  OAI22_X1 u2_uk_U659 (.A1( decrypt ) , .ZN( u2_K4_7 ) , .A2( u2_uk_n1323 ) , .B2( u2_uk_n1327 ) , .B1( u2_uk_n147 ) );
  OAI22_X1 u2_uk_U66 (.A1( decrypt ) , .ZN( u2_K4_34 ) , .B2( u2_uk_n1336 ) , .A2( u2_uk_n1352 ) , .B1( u2_uk_n147 ) );
  OAI22_X1 u2_uk_U660 (.A1( decrypt ) , .ZN( u2_K9_25 ) , .B2( u2_uk_n1578 ) , .A2( u2_uk_n1585 ) , .B1( u2_uk_n238 ) );
  OAI22_X1 u2_uk_U672 (.B1( decrypt ) , .ZN( u2_K10_43 ) , .A2( u2_uk_n1593 ) , .B2( u2_uk_n1621 ) , .A1( u2_uk_n214 ) );
  OAI22_X1 u2_uk_U674 (.B1( decrypt ) , .ZN( u2_K9_45 ) , .B2( u2_uk_n1541 ) , .A2( u2_uk_n1582 ) , .A1( u2_uk_n164 ) );
  OAI22_X1 u2_uk_U675 (.A1( decrypt ) , .ZN( u2_K7_43 ) , .A2( u2_uk_n1455 ) , .B2( u2_uk_n1484 ) , .B1( u2_uk_n164 ) );
  OAI21_X1 u2_uk_U677 (.B1( decrypt ) , .ZN( u2_K14_3 ) , .B2( u2_uk_n1812 ) , .A( u2_uk_n695 ) );
  NAND2_X1 u2_uk_U678 (.A2( decrypt ) , .A1( u2_uk_K_r12_47 ) , .ZN( u2_uk_n695 ) );
  NAND2_X1 u2_uk_U68 (.A2( decrypt ) , .A1( u2_uk_K_r1_36 ) , .ZN( u2_uk_n1011 ) );
  OAI21_X1 u2_uk_U685 (.B1( decrypt ) , .ZN( u2_K11_7 ) , .B2( u2_uk_n1661 ) , .A( u2_uk_n395 ) );
  OAI22_X1 u2_uk_U69 (.B1( decrypt ) , .ZN( u2_K2_34 ) , .B2( u2_uk_n1242 ) , .A2( u2_uk_n1273 ) , .A1( u2_uk_n161 ) );
  OAI21_X1 u2_uk_U690 (.B1( decrypt ) , .ZN( u2_K5_25 ) , .A( u2_uk_n1045 ) , .B2( u2_uk_n1383 ) );
  NAND2_X1 u2_uk_U691 (.A2( decrypt ) , .A1( u2_uk_K_r3_35 ) , .ZN( u2_uk_n1045 ) );
  NAND2_X1 u2_uk_U693 (.A2( decrypt ) , .A1( u2_uk_K_r0_22 ) , .ZN( u2_uk_n996 ) );
  OAI22_X1 u2_uk_U694 (.A1( decrypt ) , .ZN( u2_K12_25 ) , .B1( u2_uk_n148 ) , .B2( u2_uk_n1699 ) , .A2( u2_uk_n1704 ) );
  OAI22_X1 u2_uk_U695 (.A1( decrypt ) , .ZN( u2_K10_25 ) , .B1( u2_uk_n146 ) , .A2( u2_uk_n1593 ) , .B2( u2_uk_n1611 ) );
  AOI22_X1 u2_uk_U698 (.A1( decrypt ) , .B2( u2_uk_K_r11_10 ) , .A2( u2_uk_K_r11_5 ) , .B1( u2_uk_n217 ) , .ZN( u2_uk_n682 ) );
  AOI22_X1 u2_uk_U706 (.A1( decrypt ) , .B2( u2_uk_K_r2_16 ) , .A2( u2_uk_K_r2_49 ) , .ZN( u2_uk_n1027 ) , .B1( u2_uk_n148 ) );
  OAI22_X1 u2_uk_U710 (.B1( decrypt ) , .ZN( u2_K12_2 ) , .A2( u2_uk_n1681 ) , .B2( u2_uk_n1686 ) , .A1( u2_uk_n182 ) );
  OAI22_X1 u2_uk_U717 (.B1( decrypt ) , .ZN( u2_K13_32 ) , .A2( u2_uk_n1728 ) , .B2( u2_uk_n1752 ) , .A1( u2_uk_n220 ) );
  OAI21_X1 u2_uk_U718 (.B1( decrypt ) , .ZN( u2_K10_32 ) , .B2( u2_uk_n1588 ) , .A( u2_uk_n292 ) );
  NAND2_X1 u2_uk_U719 (.A2( decrypt ) , .A1( u2_uk_K_r8_51 ) , .ZN( u2_uk_n292 ) );
  OAI22_X1 u2_uk_U720 (.A1( decrypt ) , .ZN( u2_K6_32 ) , .B2( u2_uk_n1418 ) , .A2( u2_uk_n1434 ) , .B1( u2_uk_n164 ) );
  OAI22_X1 u2_uk_U721 (.A1( decrypt ) , .ZN( u2_K3_32 ) , .B2( u2_uk_n1278 ) , .A2( u2_uk_n1313 ) , .B1( u2_uk_n230 ) );
  OAI22_X1 u2_uk_U722 (.B1( decrypt ) , .ZN( u2_K5_32 ) , .B2( u2_uk_n1378 ) , .A2( u2_uk_n1382 ) , .A1( u2_uk_n238 ) );
  OAI22_X1 u2_uk_U724 (.A1( decrypt ) , .ZN( u2_K9_32 ) , .B1( u2_uk_n148 ) , .B2( u2_uk_n1571 ) , .A2( u2_uk_n1578 ) );
  OAI21_X1 u2_uk_U725 (.B1( decrypt ) , .ZN( u2_K16_42 ) , .B2( u2_uk_n1211 ) , .A( u2_uk_n962 ) );
  NAND2_X1 u2_uk_U726 (.A2( decrypt ) , .A1( u2_uk_K_r14_38 ) , .ZN( u2_uk_n962 ) );
  OAI22_X1 u2_uk_U728 (.A1( decrypt ) , .ZN( u2_K14_42 ) , .B1( u2_uk_n142 ) , .B2( u2_uk_n1768 ) , .A2( u2_uk_n1799 ) );
  OAI22_X1 u2_uk_U729 (.A1( decrypt ) , .ZN( u2_K13_42 ) , .B2( u2_uk_n1733 ) , .A2( u2_uk_n1739 ) , .B1( u2_uk_n203 ) );
  OAI22_X1 u2_uk_U730 (.A1( decrypt ) , .ZN( u2_K11_42 ) , .B1( u2_uk_n147 ) , .B2( u2_uk_n1664 ) , .A2( u2_uk_n1672 ) );
  OAI22_X1 u2_uk_U731 (.A1( decrypt ) , .ZN( u2_K10_42 ) , .B2( u2_uk_n1589 ) , .A2( u2_uk_n1615 ) , .B1( u2_uk_n202 ) );
  NAND2_X1 u2_uk_U733 (.A2( decrypt ) , .A1( u2_uk_K_r6_22 ) , .ZN( u2_uk_n1112 ) );
  OAI22_X1 u2_uk_U734 (.B1( decrypt ) , .ZN( u2_K4_42 ) , .B2( u2_uk_n1330 ) , .A2( u2_uk_n1337 ) , .A1( u2_uk_n231 ) );
  OAI22_X1 u2_uk_U735 (.B1( decrypt ) , .ZN( u2_K3_42 ) , .B2( u2_uk_n1277 ) , .A2( u2_uk_n1304 ) , .A1( u2_uk_n220 ) );
  AOI22_X1 u2_uk_U738 (.A1( decrypt ) , .B2( u2_uk_K_r5_1 ) , .A2( u2_uk_K_r5_36 ) , .ZN( u2_uk_n1093 ) , .B1( u2_uk_n147 ) );
  AOI22_X1 u2_uk_U740 (.B1( decrypt ) , .B2( u2_key_r_31 ) , .A2( u2_key_r_38 ) , .A1( u2_uk_n162 ) , .ZN( u2_uk_n986 ) );
  OAI22_X1 u2_uk_U743 (.A1( decrypt ) , .ZN( u2_K12_27 ) , .B1( u2_uk_n129 ) , .B2( u2_uk_n1687 ) , .A2( u2_uk_n1719 ) );
  OAI22_X1 u2_uk_U749 (.A1( decrypt ) , .ZN( u2_K11_13 ) , .B1( u2_uk_n164 ) , .B2( u2_uk_n1658 ) , .A2( u2_uk_n1662 ) );
  OAI22_X1 u2_uk_U751 (.B1( decrypt ) , .ZN( u2_K6_13 ) , .B2( u2_uk_n1432 ) , .A2( u2_uk_n1436 ) , .A1( u2_uk_n203 ) );
  NAND2_X1 u2_uk_U755 (.A2( decrypt ) , .A1( u2_uk_K_r7_5 ) , .ZN( u2_uk_n1120 ) );
  OAI22_X1 u2_uk_U758 (.A1( decrypt ) , .ZN( u2_K14_21 ) , .B2( u2_uk_n1784 ) , .A2( u2_uk_n1810 ) , .B1( u2_uk_n230 ) );
  OAI21_X1 u2_uk_U759 (.B1( decrypt ) , .ZN( u2_K11_21 ) , .B2( u2_uk_n1637 ) , .A( u2_uk_n346 ) );
  OAI22_X1 u2_uk_U762 (.A1( decrypt ) , .ZN( u2_K5_21 ) , .B2( u2_uk_n1379 ) , .A2( u2_uk_n1399 ) , .B1( u2_uk_n155 ) );
  OAI22_X1 u2_uk_U763 (.B1( decrypt ) , .ZN( u2_K4_21 ) , .B2( u2_uk_n1341 ) , .A2( u2_uk_n1347 ) , .A1( u2_uk_n161 ) );
  OAI22_X1 u2_uk_U765 (.A1( decrypt ) , .ZN( u2_K14_13 ) , .B2( u2_uk_n1782 ) , .A2( u2_uk_n1787 ) , .B1( u2_uk_n223 ) );
  OAI22_X1 u2_uk_U766 (.B1( decrypt ) , .ZN( u2_K15_21 ) , .A1( u2_uk_n148 ) , .A2( u2_uk_n1816 ) , .B2( u2_uk_n1820 ) );
  AOI22_X1 u2_uk_U769 (.A1( decrypt ) , .B2( u2_uk_K_r0_28 ) , .A2( u2_uk_K_r0_7 ) , .B1( u2_uk_n188 ) , .ZN( u2_uk_n997 ) );
  AOI22_X1 u2_uk_U771 (.A1( decrypt ) , .B2( u2_uk_K_r10_25 ) , .A2( u2_uk_K_r10_48 ) , .B1( u2_uk_n214 ) , .ZN( u2_uk_n443 ) );
  OAI22_X1 u2_uk_U774 (.B1( decrypt ) , .ZN( u2_K4_27 ) , .B2( u2_uk_n1320 ) , .A2( u2_uk_n1346 ) , .A1( u2_uk_n182 ) );
  AOI22_X1 u2_uk_U777 (.B1( decrypt ) , .B2( u2_uk_K_r11_34 ) , .A2( u2_uk_K_r11_39 ) , .A1( u2_uk_n203 ) , .ZN( u2_uk_n608 ) );
  OAI22_X1 u2_uk_U78 (.A1( decrypt ) , .ZN( u2_K3_23 ) , .A2( u2_uk_n1281 ) , .B2( u2_uk_n1286 ) , .B1( u2_uk_n141 ) );
  OAI22_X1 u2_uk_U784 (.B1( decrypt ) , .ZN( u2_K6_27 ) , .B2( u2_uk_n1429 ) , .A2( u2_uk_n1434 ) , .A1( u2_uk_n231 ) );
  AOI22_X1 u2_uk_U786 (.A1( decrypt ) , .B2( u2_uk_K_r3_15 ) , .A2( u2_uk_K_r3_51 ) , .ZN( u2_uk_n1046 ) , .B1( u2_uk_n209 ) );
  AOI22_X1 u2_uk_U798 (.B1( decrypt ) , .B2( u2_uk_K_r7_24 ) , .A2( u2_uk_K_r7_6 ) , .ZN( u2_uk_n1125 ) , .A1( u2_uk_n162 ) );
  NAND2_X1 u2_uk_U800 (.A2( decrypt ) , .A1( u2_uk_K_r2_20 ) , .ZN( u2_uk_n1022 ) );
  OAI22_X1 u2_uk_U801 (.B1( decrypt ) , .ZN( u2_K5_18 ) , .A2( u2_uk_n1369 ) , .B2( u2_uk_n1406 ) , .A1( u2_uk_n207 ) );
  OAI21_X1 u2_uk_U803 (.B1( decrypt ) , .ZN( u2_K13_20 ) , .B2( u2_uk_n1732 ) , .A( u2_uk_n605 ) );
  OAI21_X1 u2_uk_U805 (.B1( decrypt ) , .ZN( u2_K8_18 ) , .A( u2_uk_n1102 ) , .B2( u2_uk_n1527 ) );
  OAI22_X1 u2_uk_U807 (.B1( decrypt ) , .ZN( u2_K2_18 ) , .B2( u2_uk_n1239 ) , .A2( u2_uk_n1270 ) , .A1( u2_uk_n223 ) );
  NAND2_X1 u2_uk_U81 (.A2( decrypt ) , .A1( u2_uk_K_r14_42 ) , .ZN( u2_uk_n961 ) );
  OAI22_X1 u2_uk_U811 (.A1( decrypt ) , .ZN( u2_K15_18 ) , .B1( u2_uk_n145 ) , .B2( u2_uk_n1822 ) , .A2( u2_uk_n1852 ) );
  OAI22_X1 u2_uk_U814 (.B1( decrypt ) , .ZN( u2_K3_20 ) , .B2( u2_uk_n1290 ) , .A2( u2_uk_n1296 ) , .A1( u2_uk_n202 ) );
  OAI21_X1 u2_uk_U815 (.B1( decrypt ) , .ZN( u2_K12_20 ) , .B2( u2_uk_n1692 ) , .A( u2_uk_n437 ) );
  NAND2_X1 u2_uk_U816 (.A2( decrypt ) , .A1( u2_uk_K_r10_47 ) , .ZN( u2_uk_n437 ) );
  OAI22_X1 u2_uk_U818 (.B1( decrypt ) , .ZN( u2_K15_20 ) , .A2( u2_uk_n1815 ) , .B2( u2_uk_n1844 ) , .A1( u2_uk_n207 ) );
  AOI22_X1 u2_uk_U827 (.A1( decrypt ) , .B2( u2_uk_K_r5_18 ) , .A2( u2_uk_K_r5_53 ) , .ZN( u2_uk_n1079 ) , .B1( u2_uk_n155 ) );
  OAI22_X1 u2_uk_U829 (.A1( decrypt ) , .ZN( u2_K11_6 ) , .B2( u2_uk_n1669 ) , .A2( u2_uk_n1675 ) , .B1( u2_uk_n209 ) );
  AOI22_X1 u2_uk_U832 (.B1( decrypt ) , .B2( u2_uk_K_r10_18 ) , .A2( u2_uk_K_r10_27 ) , .A1( u2_uk_n163 ) , .ZN( u2_uk_n500 ) );
  OAI21_X1 u2_uk_U833 (.B1( decrypt ) , .ZN( u2_K13_3 ) , .B2( u2_uk_n1751 ) , .A( u2_uk_n672 ) );
  OAI22_X1 u2_uk_U835 (.B1( decrypt ) , .ZN( u2_K5_3 ) , .B2( u2_uk_n1374 ) , .A2( u2_uk_n1381 ) , .A1( u2_uk_n202 ) );
  OAI21_X1 u2_uk_U84 (.B1( decrypt ) , .ZN( u2_K8_41 ) , .A( u2_uk_n1111 ) , .B2( u2_uk_n1517 ) );
  OAI21_X1 u2_uk_U840 (.B1( decrypt ) , .ZN( u2_K5_6 ) , .A( u2_uk_n1056 ) , .B2( u2_uk_n1387 ) );
  OAI22_X1 u2_uk_U842 (.A1( decrypt ) , .ZN( u2_K7_3 ) , .B2( u2_uk_n1465 ) , .A2( u2_uk_n1487 ) , .B1( u2_uk_n187 ) );
  OAI22_X1 u2_uk_U843 (.B1( decrypt ) , .ZN( u2_K1_43 ) , .A2( u2_uk_n1149 ) , .B2( u2_uk_n1152 ) , .A1( u2_uk_n209 ) );
  OAI22_X1 u2_uk_U848 (.B1( decrypt ) , .ZN( u2_K5_41 ) , .B2( u2_uk_n1388 ) , .A2( u2_uk_n1396 ) , .A1( u2_uk_n145 ) );
  NAND2_X1 u2_uk_U85 (.A2( decrypt ) , .A1( u2_uk_K_r6_30 ) , .ZN( u2_uk_n1111 ) );
  OAI22_X1 u2_uk_U850 (.B1( decrypt ) , .ZN( u2_K6_22 ) , .B2( u2_uk_n1417 ) , .A2( u2_uk_n1422 ) , .A1( u2_uk_n155 ) );
  OAI22_X1 u2_uk_U851 (.B1( decrypt ) , .ZN( u2_K15_23 ) , .B2( u2_uk_n1833 ) , .A2( u2_uk_n1851 ) , .A1( u2_uk_n207 ) );
  OAI22_X1 u2_uk_U853 (.B1( decrypt ) , .ZN( u2_K5_23 ) , .B2( u2_uk_n1385 ) , .A2( u2_uk_n1394 ) , .A1( u2_uk_n163 ) );
  OAI22_X1 u2_uk_U854 (.B1( decrypt ) , .ZN( u2_K13_34 ) , .A1( u2_uk_n129 ) , .B2( u2_uk_n1738 ) , .A2( u2_uk_n1754 ) );
  OAI22_X1 u2_uk_U855 (.B1( decrypt ) , .ZN( u2_K5_34 ) , .A2( u2_uk_n1371 ) , .B2( u2_uk_n1384 ) , .A1( u2_uk_n162 ) );
  OAI22_X1 u2_uk_U856 (.B1( decrypt ) , .ZN( u2_K3_47 ) , .B2( u2_uk_n1297 ) , .A2( u2_uk_n1305 ) , .A1( u2_uk_n188 ) );
  OAI22_X1 u2_uk_U857 (.B1( decrypt ) , .ZN( u2_K8_5 ) , .B2( u2_uk_n1534 ) , .A2( u2_uk_n1540 ) , .A1( u2_uk_n231 ) );
  OAI22_X1 u2_uk_U865 (.B1( decrypt ) , .ZN( u2_K13_45 ) , .B2( u2_uk_n1725 ) , .A2( u2_uk_n1763 ) , .A1( u2_uk_n238 ) );
  OAI22_X1 u2_uk_U868 (.B1( decrypt ) , .ZN( u2_K3_30 ) , .B2( u2_uk_n1288 ) , .A1( u2_uk_n129 ) , .A2( u2_uk_n1314 ) );
  AOI22_X1 u2_uk_U87 (.B1( decrypt ) , .B2( u2_uk_K_r0_28 ) , .A2( u2_uk_K_r0_49 ) , .ZN( u2_uk_n1001 ) , .A1( u2_uk_n191 ) );
  OAI22_X1 u2_uk_U872 (.B1( decrypt ) , .ZN( u2_K9_3 ) , .A2( u2_uk_n1543 ) , .B2( u2_uk_n1547 ) , .A1( u2_uk_n238 ) );
  OAI22_X1 u2_uk_U878 (.B1( decrypt ) , .ZN( u2_K6_24 ) , .B2( u2_uk_n1427 ) , .A2( u2_uk_n1431 ) , .A1( u2_uk_n191 ) );
  OAI22_X1 u2_uk_U879 (.B1( decrypt ) , .ZN( u2_K15_13 ) , .A1( u2_uk_n146 ) , .A2( u2_uk_n1814 ) , .B2( u2_uk_n1842 ) );
  OAI22_X1 u2_uk_U882 (.B1( decrypt ) , .ZN( u2_K5_19 ) , .A2( u2_uk_n1368 ) , .B2( u2_uk_n1405 ) , .A1( u2_uk_n203 ) );
  OAI22_X1 u2_uk_U883 (.B1( decrypt ) , .ZN( u2_K5_24 ) , .B2( u2_uk_n1372 ) , .A2( u2_uk_n1397 ) , .A1( u2_uk_n161 ) );
  OAI22_X1 u2_uk_U889 (.B1( decrypt ) , .ZN( u2_K5_13 ) , .B2( u2_uk_n1375 ) , .A2( u2_uk_n1406 ) , .A1( u2_uk_n161 ) );
  OAI22_X1 u2_uk_U890 (.B1( decrypt ) , .ZN( u2_K5_14 ) , .B2( u2_uk_n1373 ) , .A2( u2_uk_n1380 ) , .A1( u2_uk_n213 ) );
  OAI22_X1 u2_uk_U891 (.B1( decrypt ) , .ZN( u2_K4_14 ) , .B2( u2_uk_n1322 ) , .A2( u2_uk_n1348 ) , .A1( u2_uk_n164 ) );
  OAI22_X1 u2_uk_U892 (.B1( decrypt ) , .ZN( u2_K3_13 ) , .B2( u2_uk_n1289 ) , .A2( u2_uk_n1294 ) , .A1( u2_uk_n162 ) );
  OAI22_X1 u2_uk_U902 (.B1( decrypt ) , .ZN( u2_K4_39 ) , .B2( u2_uk_n1321 ) , .A2( u2_uk_n1342 ) , .A1( u2_uk_n164 ) );
  OAI22_X1 u2_uk_U906 (.A1( decrypt ) , .ZN( u2_K14_18 ) , .B1( u2_uk_n141 ) , .B2( u2_uk_n1788 ) , .A2( u2_uk_n1796 ) );
  OAI22_X1 u2_uk_U908 (.A1( decrypt ) , .ZN( u2_K9_23 ) , .B2( u2_uk_n1554 ) , .A2( u2_uk_n1562 ) , .B1( u2_uk_n182 ) );
  OAI22_X1 u2_uk_U911 (.A1( decrypt ) , .ZN( u2_K11_16 ) , .B1( u2_uk_n146 ) , .B2( u2_uk_n1662 ) , .A2( u2_uk_n1668 ) );
  OAI22_X1 u2_uk_U912 (.A1( decrypt ) , .ZN( u2_K11_48 ) , .B2( u2_uk_n1659 ) , .A2( u2_uk_n1666 ) , .B1( u2_uk_n214 ) );
  OAI22_X1 u2_uk_U915 (.A1( decrypt ) , .ZN( u2_K14_8 ) , .B1( u2_uk_n142 ) , .A2( u2_uk_n1771 ) , .B2( u2_uk_n1789 ) );
  OAI22_X1 u2_uk_U918 (.A1( decrypt ) , .ZN( u2_K2_20 ) , .A2( u2_uk_n1233 ) , .B2( u2_uk_n1262 ) , .B1( u2_uk_n142 ) );
  OAI22_X1 u2_uk_U919 (.A1( decrypt ) , .ZN( u2_K14_14 ) , .B1( u2_uk_n145 ) , .B2( u2_uk_n1804 ) , .A2( u2_uk_n1811 ) );
  OAI22_X1 u2_uk_U92 (.A1( decrypt ) , .ZN( u2_K16_5 ) , .A2( u2_uk_n1191 ) , .B2( u2_uk_n1194 ) , .B1( u2_uk_n164 ) );
  OAI22_X1 u2_uk_U921 (.A1( decrypt ) , .ZN( u2_K8_24 ) , .B2( u2_uk_n1500 ) , .A2( u2_uk_n1540 ) , .B1( u2_uk_n191 ) );
  OAI22_X1 u2_uk_U925 (.A1( decrypt ) , .ZN( u2_K10_46 ) , .B2( u2_uk_n1602 ) , .A2( u2_uk_n1611 ) , .B1( u2_uk_n182 ) );
  OAI22_X1 u2_uk_U926 (.A1( decrypt ) , .ZN( u2_K10_34 ) , .B2( u2_uk_n1588 ) , .A2( u2_uk_n1614 ) , .B1( u2_uk_n220 ) );
  OAI22_X1 u2_uk_U93 (.A1( decrypt ) , .ZN( u2_K15_5 ) , .B1( u2_uk_n164 ) , .B2( u2_uk_n1829 ) , .A2( u2_uk_n1832 ) );
  OAI22_X1 u2_uk_U932 (.A1( decrypt ) , .ZN( u2_K2_48 ) , .B2( u2_uk_n1241 ) , .A2( u2_uk_n1256 ) , .B1( u2_uk_n209 ) );
  OAI22_X1 u2_uk_U934 (.A1( decrypt ) , .ZN( u2_K13_8 ) , .B2( u2_uk_n1751 ) , .A2( u2_uk_n1757 ) , .B1( u2_uk_n214 ) );
  OAI22_X1 u2_uk_U935 (.A1( decrypt ) , .ZN( u2_K6_20 ) , .A2( u2_uk_n1409 ) , .B2( u2_uk_n1414 ) , .B1( u2_uk_n164 ) );
  OAI22_X1 u2_uk_U936 (.A1( decrypt ) , .ZN( u2_K11_18 ) , .B2( u2_uk_n1637 ) , .A2( u2_uk_n1643 ) , .B1( u2_uk_n208 ) );
  OAI22_X1 u2_uk_U941 (.A1( decrypt ) , .ZN( u2_K14_16 ) , .B1( u2_uk_n141 ) , .A2( u2_uk_n1774 ) , .B2( u2_uk_n1812 ) );
  OAI22_X1 u2_uk_U942 (.A1( decrypt ) , .ZN( u2_K6_36 ) , .A2( u2_uk_n1411 ) , .B2( u2_uk_n1419 ) , .B1( u2_uk_n182 ) );
  OAI22_X1 u2_uk_U946 (.A1( decrypt ) , .ZN( u2_K7_37 ) , .B2( u2_uk_n1469 ) , .A2( u2_uk_n1493 ) , .B1( u2_uk_n188 ) );
  OAI22_X1 u2_uk_U948 (.A1( decrypt ) , .ZN( u2_K9_40 ) , .B2( u2_uk_n1570 ) , .A2( u2_uk_n1576 ) , .B1( u2_uk_n188 ) );
  OAI22_X1 u2_uk_U951 (.A1( decrypt ) , .ZN( u2_K11_45 ) , .B2( u2_uk_n1647 ) , .A2( u2_uk_n1654 ) , .B1( u2_uk_n214 ) );
  OAI22_X1 u2_uk_U952 (.A1( decrypt ) , .ZN( u2_K8_45 ) , .B2( u2_uk_n1498 ) , .A2( u2_uk_n1536 ) , .B1( u2_uk_n191 ) );
  OAI22_X1 u2_uk_U953 (.A1( decrypt ) , .ZN( u2_K7_45 ) , .B2( u2_uk_n1460 ) , .A2( u2_uk_n1477 ) , .B1( u2_uk_n222 ) );
  OAI22_X1 u2_uk_U956 (.A1( decrypt ) , .ZN( u2_K2_45 ) , .B2( u2_uk_n1252 ) , .A2( u2_uk_n1274 ) , .B1( u2_uk_n129 ) );
  OAI22_X1 u2_uk_U957 (.A1( decrypt ) , .ZN( u2_K6_3 ) , .B2( u2_uk_n1417 ) , .A2( u2_uk_n1431 ) , .B1( u2_uk_n164 ) );
  OAI22_X1 u2_uk_U959 (.A1( decrypt ) , .ZN( u2_K7_7 ) , .B2( u2_uk_n1466 ) , .B1( u2_uk_n148 ) , .A2( u2_uk_n1488 ) );
  OAI22_X1 u2_uk_U960 (.A1( decrypt ) , .ZN( u2_K3_7 ) , .B2( u2_uk_n1293 ) , .A2( u2_uk_n1311 ) , .B1( u2_uk_n230 ) );
  OAI22_X1 u2_uk_U961 (.A1( decrypt ) , .ZN( u2_K9_15 ) , .B2( u2_uk_n1547 ) , .A2( u2_uk_n1554 ) , .B1( u2_uk_n209 ) );
  OAI22_X1 u2_uk_U962 (.A1( decrypt ) , .ZN( u2_K6_15 ) , .B2( u2_uk_n1423 ) , .A2( u2_uk_n1435 ) , .B1( u2_uk_n202 ) );
  OAI22_X1 u2_uk_U963 (.A1( decrypt ) , .ZN( u2_K6_25 ) , .B2( u2_uk_n1424 ) , .A2( u2_uk_n1440 ) , .B1( u2_uk_n182 ) );
  OAI22_X1 u2_uk_U964 (.A1( decrypt ) , .ZN( u2_K14_25 ) , .B1( u2_uk_n142 ) , .B2( u2_uk_n1770 ) , .A2( u2_uk_n1776 ) );
  AOI22_X1 u2_uk_U969 (.B1( decrypt ) , .B2( u2_uk_K_r7_23 ) , .A2( u2_uk_K_r7_30 ) , .ZN( u2_uk_n1136 ) , .A1( u2_uk_n161 ) );
  AOI22_X1 u2_uk_U971 (.B1( decrypt ) , .B2( u2_uk_K_r10_28 ) , .A2( u2_uk_K_r10_9 ) , .A1( u2_uk_n213 ) , .ZN( u2_uk_n503 ) );
  AOI22_X1 u2_uk_U973 (.B1( decrypt ) , .B2( u2_uk_K_r7_15 ) , .A2( u2_uk_K_r7_22 ) , .ZN( u2_uk_n1137 ) , .A1( u2_uk_n161 ) );
  OAI21_X1 u2_uk_U975 (.B1( decrypt ) , .ZN( u2_K4_22 ) , .A( u2_uk_n1025 ) , .B2( u2_uk_n1327 ) );
  NAND2_X1 u2_uk_U976 (.A2( decrypt ) , .A1( u2_uk_K_r2_47 ) , .ZN( u2_uk_n1025 ) );
  NAND2_X1 u2_uk_U978 (.A2( decrypt ) , .A1( u2_uk_K_r5_13 ) , .ZN( u2_uk_n1082 ) );
  NAND2_X1 u2_uk_U980 (.A2( decrypt ) , .A1( u2_uk_K_r4_27 ) , .ZN( u2_uk_n1063 ) );
  OAI21_X1 u2_uk_U981 (.B1( decrypt ) , .ZN( u2_K3_35 ) , .A( u2_uk_n1012 ) , .B2( u2_uk_n1278 ) );
  NAND2_X1 u2_uk_U984 (.A2( decrypt ) , .A1( u2_uk_K_r12_22 ) , .ZN( u2_uk_n931 ) );
  NAND2_X1 u2_uk_U986 (.A2( decrypt ) , .A1( u2_uk_K_r2_53 ) , .ZN( u2_uk_n1038 ) );
  NAND2_X1 u2_uk_U990 (.A2( decrypt ) , .A1( u2_uk_K_r6_19 ) , .ZN( u2_uk_n1116 ) );
  NAND2_X1 u2_uk_U994 (.A2( decrypt ) , .A1( u2_uk_K_r1_10 ) , .ZN( u2_uk_n1018 ) );
endmodule
