module des_des_die_10 ( u0_FP_48, u0_FP_49, u0_FP_50, u0_FP_51, u0_FP_52, u0_FP_53, u0_FP_54, u0_FP_55, u0_FP_56, 
       u0_FP_57, u0_FP_58, u0_FP_59, u0_FP_60, u0_FP_61, u0_K13_30, u0_K13_36, u0_K13_39, u0_K13_40, 
       u0_K13_42, u0_K16_26, u0_K16_38, u0_K1_23, u0_K5_13, u0_K5_14, u0_K5_15, u0_K5_16, u0_K5_18, 
       u0_K5_19, u0_K5_23, u0_K5_24, u0_K5_9, u0_K9_45, u0_L11_11, u0_L11_12, u0_L11_14, u0_L11_19, 
       u0_L11_22, u0_L11_25, u0_L11_29, u0_L11_3, u0_L11_32, u0_L11_4, u0_L11_7, u0_L11_8, u0_L14_11, 
       u0_L14_12, u0_L14_14, u0_L14_19, u0_L14_22, u0_L14_25, u0_L14_29, u0_L14_3, u0_L14_32, u0_L14_4, 
       u0_L14_7, u0_L14_8, u0_L3_1, u0_L3_10, u0_L3_13, u0_L3_16, u0_L3_18, u0_L3_2, u0_L3_20, 
       u0_L3_24, u0_L3_26, u0_L3_28, u0_L3_30, u0_L3_6, u0_L5_11, u0_L5_12, u0_L5_14, u0_L5_19, 
       u0_L5_22, u0_L5_25, u0_L5_29, u0_L5_3, u0_L5_32, u0_L5_4, u0_L5_7, u0_L5_8, u0_L7_1, 
       u0_L7_10, u0_L7_14, u0_L7_15, u0_L7_20, u0_L7_21, u0_L7_25, u0_L7_26, u0_L7_27, u0_L7_3, 
       u0_L7_5, u0_L7_8, u0_R11_16, u0_R11_17, u0_R11_18, u0_R11_19, u0_R11_20, u0_R11_21, u0_R11_22, 
       u0_R11_23, u0_R11_24, u0_R11_25, u0_R11_26, u0_R11_27, u0_R11_28, u0_R11_29, u0_R3_10, u0_R3_11, 
       u0_R3_12, u0_R3_13, u0_R3_14, u0_R3_15, u0_R3_16, u0_R3_17, u0_R3_4, u0_R3_5, u0_R3_6, 
       u0_R3_7, u0_R3_8, u0_R3_9, u0_R5_16, u0_R5_17, u0_R5_18, u0_R5_19, u0_R5_20, u0_R5_21, 
       u0_R5_22, u0_R5_23, u0_R5_24, u0_R5_25, u0_R5_26, u0_R5_27, u0_R5_28, u0_R5_29, u0_R7_1, 
       u0_R7_12, u0_R7_13, u0_R7_14, u0_R7_15, u0_R7_16, u0_R7_17, u0_R7_18, u0_R7_19, u0_R7_20, 
       u0_R7_21, u0_R7_28, u0_R7_29, u0_R7_30, u0_R7_31, u0_R7_32, u0_desIn_r_10, u0_desIn_r_12, u0_desIn_r_14, 
       u0_desIn_r_15, u0_desIn_r_2, u0_desIn_r_23, u0_desIn_r_24, u0_desIn_r_26, u0_desIn_r_29, u0_desIn_r_3, u0_desIn_r_31, u0_desIn_r_36, 
       u0_desIn_r_37, u0_desIn_r_39, u0_desIn_r_4, u0_desIn_r_45, u0_desIn_r_47, u0_desIn_r_48, u0_desIn_r_5, u0_desIn_r_50, u0_desIn_r_53, 
       u0_desIn_r_55, u0_desIn_r_57, u0_desIn_r_6, u0_desIn_r_61, u0_desIn_r_63, u0_desIn_r_7, u0_desIn_r_8, u0_key_r_11, u0_key_r_12, 
       u0_key_r_13, u0_key_r_17, u0_key_r_19, u0_key_r_20, u0_key_r_24, u0_key_r_25, u0_key_r_26, u0_key_r_27, u0_key_r_3, 
       u0_key_r_32, u0_key_r_34, u0_key_r_39, u0_key_r_4, u0_key_r_40, u0_key_r_41, u0_key_r_47, u0_key_r_48, u0_key_r_49, 
       u0_key_r_53, u0_key_r_54, u0_key_r_55, u0_key_r_6, u0_uk_K_r11_21, u0_uk_K_r14_15, u0_uk_K_r14_2, u0_uk_K_r14_45, u0_uk_K_r14_50, 
       u0_uk_K_r14_8, u0_uk_K_r14_9, u0_uk_K_r3_11, u0_uk_K_r3_19, u0_uk_K_r3_24, u0_uk_K_r3_47, u0_uk_K_r4_31, u0_uk_K_r5_0, u0_uk_K_r5_1, 
       u0_uk_K_r5_16, u0_uk_K_r5_21, u0_uk_K_r5_23, u0_uk_K_r5_37, u0_uk_K_r5_43, u0_uk_K_r5_51, u0_uk_K_r5_8, u0_uk_K_r7_0, u0_uk_K_r7_2, 
       u0_uk_K_r7_32, u0_uk_K_r7_39, u0_uk_K_r7_9, u0_uk_n10, u0_uk_n100, u0_uk_n102, u0_uk_n103, u0_uk_n104, u0_uk_n105, 
       u0_uk_n106, u0_uk_n109, u0_uk_n11, u0_uk_n110, u0_uk_n111, u0_uk_n112, u0_uk_n113, u0_uk_n116, u0_uk_n118, 
       u0_uk_n120, u0_uk_n123, u0_uk_n124, u0_uk_n128, u0_uk_n129, u0_uk_n130, u0_uk_n134, u0_uk_n135, u0_uk_n141, 
       u0_uk_n142, u0_uk_n145, u0_uk_n146, u0_uk_n147, u0_uk_n161, u0_uk_n162, u0_uk_n163, u0_uk_n182, u0_uk_n188, 
       u0_uk_n191, u0_uk_n202, u0_uk_n203, u0_uk_n208, u0_uk_n209, u0_uk_n213, u0_uk_n214, u0_uk_n217, u0_uk_n222, 
       u0_uk_n223, u0_uk_n231, u0_uk_n238, u0_uk_n240, u0_uk_n242, u0_uk_n250, u0_uk_n251, u0_uk_n252, u0_uk_n257, 
       u0_uk_n27, u0_uk_n272, u0_uk_n273, u0_uk_n274, u0_uk_n275, u0_uk_n280, u0_uk_n281, u0_uk_n282, u0_uk_n285, 
       u0_uk_n288, u0_uk_n289, u0_uk_n290, u0_uk_n293, u0_uk_n296, u0_uk_n300, u0_uk_n304, u0_uk_n31, u0_uk_n314, 
       u0_uk_n365, u0_uk_n367, u0_uk_n368, u0_uk_n372, u0_uk_n374, u0_uk_n378, u0_uk_n380, u0_uk_n387, u0_uk_n388, 
       u0_uk_n389, u0_uk_n394, u0_uk_n398, u0_uk_n399, u0_uk_n402, u0_uk_n406, u0_uk_n451, u0_uk_n453, u0_uk_n459, 
       u0_uk_n464, u0_uk_n465, u0_uk_n473, u0_uk_n479, u0_uk_n483, u0_uk_n484, u0_uk_n485, u0_uk_n489, u0_uk_n60, 
       u0_uk_n63, u0_uk_n632, u0_uk_n633, u0_uk_n638, u0_uk_n642, u0_uk_n643, u0_uk_n647, u0_uk_n648, u0_uk_n649, 
       u0_uk_n650, u0_uk_n655, u0_uk_n657, u0_uk_n658, u0_uk_n663, u0_uk_n666, u0_uk_n669, u0_uk_n670, u0_uk_n719, 
       u0_uk_n720, u0_uk_n728, u0_uk_n731, u0_uk_n732, u0_uk_n735, u0_uk_n766, u0_uk_n770, u0_uk_n775, u0_uk_n815, 
       u0_uk_n83, u0_uk_n897, u0_uk_n898, u0_uk_n904, u0_uk_n92, u0_uk_n93, u0_uk_n94, u0_uk_n948, u0_uk_n95, 
       u0_uk_n97, u0_uk_n98, u2_K11_11, u2_K11_13, u2_K11_16, u2_K11_18, u2_K11_21, u2_K11_4, u2_K11_6, 
       u2_K11_7, u2_K11_9, u2_K13_20, u2_K13_26, u2_K13_31, u2_K13_32, u2_K13_34, u2_K14_25, u2_K14_28, 
       u2_K3_20, u2_K3_23, u2_K3_30, u2_K3_32, u2_K3_35, u2_K3_42, u2_K3_43, u2_K3_47, u2_K3_48, 
       u2_K4_27, u2_K4_33, u2_K4_34, u2_K4_35, u2_K4_38, u2_K4_39, u2_K4_42, u2_K6_1, u2_K6_11, 
       u2_K6_3, u2_L11_1, u2_L11_10, u2_L11_11, u2_L11_14, u2_L11_19, u2_L11_20, u2_L11_25, u2_L11_26, 
       u2_L11_29, u2_L11_3, u2_L11_4, u2_L11_8, u2_L12_14, u2_L12_25, u2_L12_3, u2_L12_8, u2_L1_1, 
       u2_L1_10, u2_L1_11, u2_L1_12, u2_L1_14, u2_L1_15, u2_L1_19, u2_L1_20, u2_L1_21, u2_L1_22, 
       u2_L1_25, u2_L1_26, u2_L1_27, u2_L1_29, u2_L1_3, u2_L1_32, u2_L1_4, u2_L1_5, u2_L1_7, 
       u2_L1_8, u2_L2_11, u2_L2_12, u2_L2_14, u2_L2_19, u2_L2_22, u2_L2_25, u2_L2_29, u2_L2_3, 
       u2_L2_32, u2_L2_4, u2_L2_7, u2_L2_8, u2_L4_13, u2_L4_15, u2_L4_17, u2_L4_18, u2_L4_2, 
       u2_L4_21, u2_L4_23, u2_L4_27, u2_L4_28, u2_L4_31, u2_L4_5, u2_L4_9, u2_L9_1, u2_L9_10, 
       u2_L9_13, u2_L9_16, u2_L9_17, u2_L9_18, u2_L9_2, u2_L9_20, u2_L9_23, u2_L9_24, u2_L9_26, 
       u2_L9_28, u2_L9_30, u2_L9_31, u2_L9_6, u2_L9_9, u2_R11_12, u2_R11_13, u2_R11_14, u2_R11_15, 
       u2_R11_16, u2_R11_17, u2_R11_18, u2_R11_19, u2_R11_20, u2_R11_21, u2_R11_22, u2_R11_23, u2_R11_24, 
       u2_R11_25, u2_R12_16, u2_R12_17, u2_R12_18, u2_R12_19, u2_R12_20, u2_R12_21, u2_R1_1, u2_R1_12, 
       u2_R1_13, u2_R1_14, u2_R1_15, u2_R1_16, u2_R1_17, u2_R1_18, u2_R1_19, u2_R1_20, u2_R1_21, 
       u2_R1_22, u2_R1_23, u2_R1_24, u2_R1_25, u2_R1_26, u2_R1_27, u2_R1_28, u2_R1_29, u2_R1_30, 
       u2_R1_31, u2_R1_32, u2_R2_16, u2_R2_17, u2_R2_18, u2_R2_19, u2_R2_20, u2_R2_21, u2_R2_22, 
       u2_R2_23, u2_R2_24, u2_R2_25, u2_R2_26, u2_R2_27, u2_R2_28, u2_R2_29, u2_R4_1, u2_R4_2, 
       u2_R4_28, u2_R4_29, u2_R4_3, u2_R4_30, u2_R4_31, u2_R4_32, u2_R4_4, u2_R4_5, u2_R4_6, 
       u2_R4_7, u2_R4_8, u2_R4_9, u2_R9_1, u2_R9_10, u2_R9_11, u2_R9_12, u2_R9_13, u2_R9_14, 
       u2_R9_15, u2_R9_16, u2_R9_17, u2_R9_2, u2_R9_3, u2_R9_32, u2_R9_4, u2_R9_5, u2_R9_6, 
       u2_R9_7, u2_R9_8, u2_R9_9, u2_uk_K_r11_10, u2_uk_K_r11_19, u2_uk_K_r11_21, u2_uk_K_r11_28, u2_uk_K_r11_39, u2_uk_K_r11_4, 
       u2_uk_K_r11_47, u2_uk_K_r12_42, u2_uk_K_r1_15, u2_uk_K_r1_16, u2_uk_K_r1_17, u2_uk_K_r1_21, u2_uk_K_r1_22, u2_uk_K_r1_41, u2_uk_K_r1_42, 
       u2_uk_K_r1_44, u2_uk_K_r2_21, u2_uk_K_r2_24, u2_uk_K_r2_28, u2_uk_K_r2_31, u2_uk_K_r2_36, u2_uk_K_r2_49, u2_uk_K_r3_10, u2_uk_K_r4_17, 
       u2_uk_K_r4_3, u2_uk_K_r4_33, u2_uk_K_r4_41, u2_uk_K_r4_47, u2_uk_K_r4_54, u2_uk_K_r4_55, u2_uk_K_r9_10, u2_uk_K_r9_12, u2_uk_K_r9_13, 
       u2_uk_K_r9_18, u2_uk_K_r9_19, u2_uk_K_r9_25, u2_uk_K_r9_27, u2_uk_K_r9_4, u2_uk_K_r9_48, u2_uk_K_r9_54, u2_uk_K_r9_55, u2_uk_n10, 
       u2_uk_n100, u2_uk_n1007, u2_uk_n1011, u2_uk_n102, u2_uk_n1027, u2_uk_n1028, u2_uk_n1070, u2_uk_n1073, u2_uk_n1074, 
       u2_uk_n109, u2_uk_n11, u2_uk_n110, u2_uk_n117, u2_uk_n118, u2_uk_n1279, u2_uk_n128, u2_uk_n1281, u2_uk_n1283, 
       u2_uk_n1284, u2_uk_n1288, u2_uk_n129, u2_uk_n1291, u2_uk_n1292, u2_uk_n1294, u2_uk_n1297, u2_uk_n1298, u2_uk_n1299, 
       u2_uk_n1300, u2_uk_n1303, u2_uk_n1305, u2_uk_n1308, u2_uk_n1309, u2_uk_n1312, u2_uk_n1313, u2_uk_n1314, u2_uk_n1315, 
       u2_uk_n1316, u2_uk_n1319, u2_uk_n1326, u2_uk_n1331, u2_uk_n1336, u2_uk_n1342, u2_uk_n1345, u2_uk_n1346, u2_uk_n1350, 
       u2_uk_n1351, u2_uk_n1352, u2_uk_n1408, u2_uk_n141, u2_uk_n1410, u2_uk_n1413, u2_uk_n1416, u2_uk_n1419, u2_uk_n142, 
       u2_uk_n1422, u2_uk_n1424, u2_uk_n1426, u2_uk_n1428, u2_uk_n1429, u2_uk_n1433, u2_uk_n1435, u2_uk_n1440, u2_uk_n1441, 
       u2_uk_n1444, u2_uk_n1446, u2_uk_n1447, u2_uk_n1448, u2_uk_n145, u2_uk_n146, u2_uk_n147, u2_uk_n148, u2_uk_n155, 
       u2_uk_n161, u2_uk_n162, u2_uk_n163, u2_uk_n1633, u2_uk_n1639, u2_uk_n164, u2_uk_n1643, u2_uk_n1646, u2_uk_n1652, 
       u2_uk_n1657, u2_uk_n1658, u2_uk_n1661, u2_uk_n1668, u2_uk_n1675, u2_uk_n1677, u2_uk_n17, u2_uk_n1723, u2_uk_n1724, 
       u2_uk_n1726, u2_uk_n1728, u2_uk_n1734, u2_uk_n1735, u2_uk_n1737, u2_uk_n1742, u2_uk_n1745, u2_uk_n1746, u2_uk_n1747, 
       u2_uk_n1753, u2_uk_n1760, u2_uk_n1763, u2_uk_n1767, u2_uk_n1781, u2_uk_n1792, u2_uk_n1807, u2_uk_n1808, u2_uk_n1809, 
       u2_uk_n182, u2_uk_n187, u2_uk_n188, u2_uk_n191, u2_uk_n202, u2_uk_n207, u2_uk_n208, u2_uk_n209, u2_uk_n213, 
       u2_uk_n214, u2_uk_n217, u2_uk_n222, u2_uk_n223, u2_uk_n231, u2_uk_n238, u2_uk_n27, u2_uk_n31, u2_uk_n313, 
       u2_uk_n319, u2_uk_n60, u2_uk_n608, u2_uk_n63, u2_uk_n689, u2_uk_n83, u2_uk_n92, u2_uk_n93, u2_uk_n94, 
       u2_uk_n99, u0_FP_11, u0_FP_12, u0_FP_14, u0_FP_19, u0_FP_22, u0_FP_25, u0_FP_29, u0_FP_3, u0_FP_32, 
        u0_FP_4, u0_FP_7, u0_FP_8, u0_N0, u0_N1, u0_N12, u0_N128, u0_N129, u0_N133, 
        u0_N137, u0_N140, u0_N143, u0_N145, u0_N147, u0_N151, u0_N153, u0_N155, u0_N157, 
        u0_N16, u0_N17, u0_N19, u0_N194, u0_N195, u0_N198, u0_N199, u0_N202, u0_N203, 
        u0_N205, u0_N210, u0_N213, u0_N216, u0_N22, u0_N220, u0_N223, u0_N25, u0_N256, 
        u0_N258, u0_N260, u0_N263, u0_N265, u0_N269, u0_N27, u0_N270, u0_N275, u0_N276, 
        u0_N280, u0_N281, u0_N282, u0_N30, u0_N386, u0_N387, u0_N390, u0_N391, u0_N394, 
        u0_N395, u0_N397, u0_N402, u0_N405, u0_N408, u0_N412, u0_N415, u0_N8, u0_N9, 
        u0_uk_n117, u0_uk_n155, u0_uk_n187, u0_uk_n230, u0_uk_n674, u0_uk_n684, u0_uk_n690, u0_uk_n696, u0_uk_n697, 
        u0_uk_n698, u0_uk_n705, u0_uk_n790, u0_uk_n871, u0_uk_n99, u2_N102, u2_N103, u2_N106, u2_N107, 
        u2_N109, u2_N114, u2_N117, u2_N120, u2_N124, u2_N127, u2_N161, u2_N164, u2_N168, 
        u2_N172, u2_N174, u2_N176, u2_N177, u2_N180, u2_N182, u2_N186, u2_N187, u2_N190, 
        u2_N320, u2_N321, u2_N325, u2_N328, u2_N329, u2_N332, u2_N335, u2_N336, u2_N337, 
        u2_N339, u2_N342, u2_N343, u2_N345, u2_N347, u2_N349, u2_N350, u2_N384, u2_N386, 
        u2_N387, u2_N391, u2_N393, u2_N394, u2_N397, u2_N402, u2_N403, u2_N408, u2_N409, 
        u2_N412, u2_N418, u2_N423, u2_N429, u2_N440, u2_N64, u2_N66, u2_N67, u2_N68, 
        u2_N70, u2_N71, u2_N73, u2_N74, u2_N75, u2_N77, u2_N78, u2_N82, u2_N83, 
        u2_N84, u2_N85, u2_N88, u2_N89, u2_N90, u2_N92, u2_N95, u2_N98, u2_N99, 
        u2_uk_n1039, u2_uk_n1056, u2_uk_n230, u2_uk_n672 );
  input u0_FP_48, u0_FP_49, u0_FP_50, u0_FP_51, u0_FP_52, u0_FP_53, u0_FP_54, u0_FP_55, u0_FP_56, 
        u0_FP_57, u0_FP_58, u0_FP_59, u0_FP_60, u0_FP_61, u0_K13_30, u0_K13_36, u0_K13_39, u0_K13_40, 
        u0_K13_42, u0_K16_26, u0_K16_38, u0_K1_23, u0_K5_13, u0_K5_14, u0_K5_15, u0_K5_16, u0_K5_18, 
        u0_K5_19, u0_K5_23, u0_K5_24, u0_K5_9, u0_K9_45, u0_L11_11, u0_L11_12, u0_L11_14, u0_L11_19, 
        u0_L11_22, u0_L11_25, u0_L11_29, u0_L11_3, u0_L11_32, u0_L11_4, u0_L11_7, u0_L11_8, u0_L14_11, 
        u0_L14_12, u0_L14_14, u0_L14_19, u0_L14_22, u0_L14_25, u0_L14_29, u0_L14_3, u0_L14_32, u0_L14_4, 
        u0_L14_7, u0_L14_8, u0_L3_1, u0_L3_10, u0_L3_13, u0_L3_16, u0_L3_18, u0_L3_2, u0_L3_20, 
        u0_L3_24, u0_L3_26, u0_L3_28, u0_L3_30, u0_L3_6, u0_L5_11, u0_L5_12, u0_L5_14, u0_L5_19, 
        u0_L5_22, u0_L5_25, u0_L5_29, u0_L5_3, u0_L5_32, u0_L5_4, u0_L5_7, u0_L5_8, u0_L7_1, 
        u0_L7_10, u0_L7_14, u0_L7_15, u0_L7_20, u0_L7_21, u0_L7_25, u0_L7_26, u0_L7_27, u0_L7_3, 
        u0_L7_5, u0_L7_8, u0_R11_16, u0_R11_17, u0_R11_18, u0_R11_19, u0_R11_20, u0_R11_21, u0_R11_22, 
        u0_R11_23, u0_R11_24, u0_R11_25, u0_R11_26, u0_R11_27, u0_R11_28, u0_R11_29, u0_R3_10, u0_R3_11, 
        u0_R3_12, u0_R3_13, u0_R3_14, u0_R3_15, u0_R3_16, u0_R3_17, u0_R3_4, u0_R3_5, u0_R3_6, 
        u0_R3_7, u0_R3_8, u0_R3_9, u0_R5_16, u0_R5_17, u0_R5_18, u0_R5_19, u0_R5_20, u0_R5_21, 
        u0_R5_22, u0_R5_23, u0_R5_24, u0_R5_25, u0_R5_26, u0_R5_27, u0_R5_28, u0_R5_29, u0_R7_1, 
        u0_R7_12, u0_R7_13, u0_R7_14, u0_R7_15, u0_R7_16, u0_R7_17, u0_R7_18, u0_R7_19, u0_R7_20, 
        u0_R7_21, u0_R7_28, u0_R7_29, u0_R7_30, u0_R7_31, u0_R7_32, u0_desIn_r_10, u0_desIn_r_12, u0_desIn_r_14, 
        u0_desIn_r_15, u0_desIn_r_2, u0_desIn_r_23, u0_desIn_r_24, u0_desIn_r_26, u0_desIn_r_29, u0_desIn_r_3, u0_desIn_r_31, u0_desIn_r_36, 
        u0_desIn_r_37, u0_desIn_r_39, u0_desIn_r_4, u0_desIn_r_45, u0_desIn_r_47, u0_desIn_r_48, u0_desIn_r_5, u0_desIn_r_50, u0_desIn_r_53, 
        u0_desIn_r_55, u0_desIn_r_57, u0_desIn_r_6, u0_desIn_r_61, u0_desIn_r_63, u0_desIn_r_7, u0_desIn_r_8, u0_key_r_11, u0_key_r_12, 
        u0_key_r_13, u0_key_r_17, u0_key_r_19, u0_key_r_20, u0_key_r_24, u0_key_r_25, u0_key_r_26, u0_key_r_27, u0_key_r_3, 
        u0_key_r_32, u0_key_r_34, u0_key_r_39, u0_key_r_4, u0_key_r_40, u0_key_r_41, u0_key_r_47, u0_key_r_48, u0_key_r_49, 
        u0_key_r_53, u0_key_r_54, u0_key_r_55, u0_key_r_6, u0_uk_K_r11_21, u0_uk_K_r14_15, u0_uk_K_r14_2, u0_uk_K_r14_45, u0_uk_K_r14_50, 
        u0_uk_K_r14_8, u0_uk_K_r14_9, u0_uk_K_r3_11, u0_uk_K_r3_19, u0_uk_K_r3_24, u0_uk_K_r3_47, u0_uk_K_r4_31, u0_uk_K_r5_0, u0_uk_K_r5_1, 
        u0_uk_K_r5_16, u0_uk_K_r5_21, u0_uk_K_r5_23, u0_uk_K_r5_37, u0_uk_K_r5_43, u0_uk_K_r5_51, u0_uk_K_r5_8, u0_uk_K_r7_0, u0_uk_K_r7_2, 
        u0_uk_K_r7_32, u0_uk_K_r7_39, u0_uk_K_r7_9, u0_uk_n10, u0_uk_n100, u0_uk_n102, u0_uk_n103, u0_uk_n104, u0_uk_n105, 
        u0_uk_n106, u0_uk_n109, u0_uk_n11, u0_uk_n110, u0_uk_n111, u0_uk_n112, u0_uk_n113, u0_uk_n116, u0_uk_n118, 
        u0_uk_n120, u0_uk_n123, u0_uk_n124, u0_uk_n128, u0_uk_n129, u0_uk_n130, u0_uk_n134, u0_uk_n135, u0_uk_n141, 
        u0_uk_n142, u0_uk_n145, u0_uk_n146, u0_uk_n147, u0_uk_n161, u0_uk_n162, u0_uk_n163, u0_uk_n182, u0_uk_n188, 
        u0_uk_n191, u0_uk_n202, u0_uk_n203, u0_uk_n208, u0_uk_n209, u0_uk_n213, u0_uk_n214, u0_uk_n217, u0_uk_n222, 
        u0_uk_n223, u0_uk_n231, u0_uk_n238, u0_uk_n240, u0_uk_n242, u0_uk_n250, u0_uk_n251, u0_uk_n252, u0_uk_n257, 
        u0_uk_n27, u0_uk_n272, u0_uk_n273, u0_uk_n274, u0_uk_n275, u0_uk_n280, u0_uk_n281, u0_uk_n282, u0_uk_n285, 
        u0_uk_n288, u0_uk_n289, u0_uk_n290, u0_uk_n293, u0_uk_n296, u0_uk_n300, u0_uk_n304, u0_uk_n31, u0_uk_n314, 
        u0_uk_n365, u0_uk_n367, u0_uk_n368, u0_uk_n372, u0_uk_n374, u0_uk_n378, u0_uk_n380, u0_uk_n387, u0_uk_n388, 
        u0_uk_n389, u0_uk_n394, u0_uk_n398, u0_uk_n399, u0_uk_n402, u0_uk_n406, u0_uk_n451, u0_uk_n453, u0_uk_n459, 
        u0_uk_n464, u0_uk_n465, u0_uk_n473, u0_uk_n479, u0_uk_n483, u0_uk_n484, u0_uk_n485, u0_uk_n489, u0_uk_n60, 
        u0_uk_n63, u0_uk_n632, u0_uk_n633, u0_uk_n638, u0_uk_n642, u0_uk_n643, u0_uk_n647, u0_uk_n648, u0_uk_n649, 
        u0_uk_n650, u0_uk_n655, u0_uk_n657, u0_uk_n658, u0_uk_n663, u0_uk_n666, u0_uk_n669, u0_uk_n670, u0_uk_n719, 
        u0_uk_n720, u0_uk_n728, u0_uk_n731, u0_uk_n732, u0_uk_n735, u0_uk_n766, u0_uk_n770, u0_uk_n775, u0_uk_n815, 
        u0_uk_n83, u0_uk_n897, u0_uk_n898, u0_uk_n904, u0_uk_n92, u0_uk_n93, u0_uk_n94, u0_uk_n948, u0_uk_n95, 
        u0_uk_n97, u0_uk_n98, u2_K11_11, u2_K11_13, u2_K11_16, u2_K11_18, u2_K11_21, u2_K11_4, u2_K11_6, 
        u2_K11_7, u2_K11_9, u2_K13_20, u2_K13_26, u2_K13_31, u2_K13_32, u2_K13_34, u2_K14_25, u2_K14_28, 
        u2_K3_20, u2_K3_23, u2_K3_30, u2_K3_32, u2_K3_35, u2_K3_42, u2_K3_43, u2_K3_47, u2_K3_48, 
        u2_K4_27, u2_K4_33, u2_K4_34, u2_K4_35, u2_K4_38, u2_K4_39, u2_K4_42, u2_K6_1, u2_K6_11, 
        u2_K6_3, u2_L11_1, u2_L11_10, u2_L11_11, u2_L11_14, u2_L11_19, u2_L11_20, u2_L11_25, u2_L11_26, 
        u2_L11_29, u2_L11_3, u2_L11_4, u2_L11_8, u2_L12_14, u2_L12_25, u2_L12_3, u2_L12_8, u2_L1_1, 
        u2_L1_10, u2_L1_11, u2_L1_12, u2_L1_14, u2_L1_15, u2_L1_19, u2_L1_20, u2_L1_21, u2_L1_22, 
        u2_L1_25, u2_L1_26, u2_L1_27, u2_L1_29, u2_L1_3, u2_L1_32, u2_L1_4, u2_L1_5, u2_L1_7, 
        u2_L1_8, u2_L2_11, u2_L2_12, u2_L2_14, u2_L2_19, u2_L2_22, u2_L2_25, u2_L2_29, u2_L2_3, 
        u2_L2_32, u2_L2_4, u2_L2_7, u2_L2_8, u2_L4_13, u2_L4_15, u2_L4_17, u2_L4_18, u2_L4_2, 
        u2_L4_21, u2_L4_23, u2_L4_27, u2_L4_28, u2_L4_31, u2_L4_5, u2_L4_9, u2_L9_1, u2_L9_10, 
        u2_L9_13, u2_L9_16, u2_L9_17, u2_L9_18, u2_L9_2, u2_L9_20, u2_L9_23, u2_L9_24, u2_L9_26, 
        u2_L9_28, u2_L9_30, u2_L9_31, u2_L9_6, u2_L9_9, u2_R11_12, u2_R11_13, u2_R11_14, u2_R11_15, 
        u2_R11_16, u2_R11_17, u2_R11_18, u2_R11_19, u2_R11_20, u2_R11_21, u2_R11_22, u2_R11_23, u2_R11_24, 
        u2_R11_25, u2_R12_16, u2_R12_17, u2_R12_18, u2_R12_19, u2_R12_20, u2_R12_21, u2_R1_1, u2_R1_12, 
        u2_R1_13, u2_R1_14, u2_R1_15, u2_R1_16, u2_R1_17, u2_R1_18, u2_R1_19, u2_R1_20, u2_R1_21, 
        u2_R1_22, u2_R1_23, u2_R1_24, u2_R1_25, u2_R1_26, u2_R1_27, u2_R1_28, u2_R1_29, u2_R1_30, 
        u2_R1_31, u2_R1_32, u2_R2_16, u2_R2_17, u2_R2_18, u2_R2_19, u2_R2_20, u2_R2_21, u2_R2_22, 
        u2_R2_23, u2_R2_24, u2_R2_25, u2_R2_26, u2_R2_27, u2_R2_28, u2_R2_29, u2_R4_1, u2_R4_2, 
        u2_R4_28, u2_R4_29, u2_R4_3, u2_R4_30, u2_R4_31, u2_R4_32, u2_R4_4, u2_R4_5, u2_R4_6, 
        u2_R4_7, u2_R4_8, u2_R4_9, u2_R9_1, u2_R9_10, u2_R9_11, u2_R9_12, u2_R9_13, u2_R9_14, 
        u2_R9_15, u2_R9_16, u2_R9_17, u2_R9_2, u2_R9_3, u2_R9_32, u2_R9_4, u2_R9_5, u2_R9_6, 
        u2_R9_7, u2_R9_8, u2_R9_9, u2_uk_K_r11_10, u2_uk_K_r11_19, u2_uk_K_r11_21, u2_uk_K_r11_28, u2_uk_K_r11_39, u2_uk_K_r11_4, 
        u2_uk_K_r11_47, u2_uk_K_r12_42, u2_uk_K_r1_15, u2_uk_K_r1_16, u2_uk_K_r1_17, u2_uk_K_r1_21, u2_uk_K_r1_22, u2_uk_K_r1_41, u2_uk_K_r1_42, 
        u2_uk_K_r1_44, u2_uk_K_r2_21, u2_uk_K_r2_24, u2_uk_K_r2_28, u2_uk_K_r2_31, u2_uk_K_r2_36, u2_uk_K_r2_49, u2_uk_K_r3_10, u2_uk_K_r4_17, 
        u2_uk_K_r4_3, u2_uk_K_r4_33, u2_uk_K_r4_41, u2_uk_K_r4_47, u2_uk_K_r4_54, u2_uk_K_r4_55, u2_uk_K_r9_10, u2_uk_K_r9_12, u2_uk_K_r9_13, 
        u2_uk_K_r9_18, u2_uk_K_r9_19, u2_uk_K_r9_25, u2_uk_K_r9_27, u2_uk_K_r9_4, u2_uk_K_r9_48, u2_uk_K_r9_54, u2_uk_K_r9_55, u2_uk_n10, 
        u2_uk_n100, u2_uk_n1007, u2_uk_n1011, u2_uk_n102, u2_uk_n1027, u2_uk_n1028, u2_uk_n1070, u2_uk_n1073, u2_uk_n1074, 
        u2_uk_n109, u2_uk_n11, u2_uk_n110, u2_uk_n117, u2_uk_n118, u2_uk_n1279, u2_uk_n128, u2_uk_n1281, u2_uk_n1283, 
        u2_uk_n1284, u2_uk_n1288, u2_uk_n129, u2_uk_n1291, u2_uk_n1292, u2_uk_n1294, u2_uk_n1297, u2_uk_n1298, u2_uk_n1299, 
        u2_uk_n1300, u2_uk_n1303, u2_uk_n1305, u2_uk_n1308, u2_uk_n1309, u2_uk_n1312, u2_uk_n1313, u2_uk_n1314, u2_uk_n1315, 
        u2_uk_n1316, u2_uk_n1319, u2_uk_n1326, u2_uk_n1331, u2_uk_n1336, u2_uk_n1342, u2_uk_n1345, u2_uk_n1346, u2_uk_n1350, 
        u2_uk_n1351, u2_uk_n1352, u2_uk_n1408, u2_uk_n141, u2_uk_n1410, u2_uk_n1413, u2_uk_n1416, u2_uk_n1419, u2_uk_n142, 
        u2_uk_n1422, u2_uk_n1424, u2_uk_n1426, u2_uk_n1428, u2_uk_n1429, u2_uk_n1433, u2_uk_n1435, u2_uk_n1440, u2_uk_n1441, 
        u2_uk_n1444, u2_uk_n1446, u2_uk_n1447, u2_uk_n1448, u2_uk_n145, u2_uk_n146, u2_uk_n147, u2_uk_n148, u2_uk_n155, 
        u2_uk_n161, u2_uk_n162, u2_uk_n163, u2_uk_n1633, u2_uk_n1639, u2_uk_n164, u2_uk_n1643, u2_uk_n1646, u2_uk_n1652, 
        u2_uk_n1657, u2_uk_n1658, u2_uk_n1661, u2_uk_n1668, u2_uk_n1675, u2_uk_n1677, u2_uk_n17, u2_uk_n1723, u2_uk_n1724, 
        u2_uk_n1726, u2_uk_n1728, u2_uk_n1734, u2_uk_n1735, u2_uk_n1737, u2_uk_n1742, u2_uk_n1745, u2_uk_n1746, u2_uk_n1747, 
        u2_uk_n1753, u2_uk_n1760, u2_uk_n1763, u2_uk_n1767, u2_uk_n1781, u2_uk_n1792, u2_uk_n1807, u2_uk_n1808, u2_uk_n1809, 
        u2_uk_n182, u2_uk_n187, u2_uk_n188, u2_uk_n191, u2_uk_n202, u2_uk_n207, u2_uk_n208, u2_uk_n209, u2_uk_n213, 
        u2_uk_n214, u2_uk_n217, u2_uk_n222, u2_uk_n223, u2_uk_n231, u2_uk_n238, u2_uk_n27, u2_uk_n31, u2_uk_n313, 
        u2_uk_n319, u2_uk_n60, u2_uk_n608, u2_uk_n63, u2_uk_n689, u2_uk_n83, u2_uk_n92, u2_uk_n93, u2_uk_n94, 
        u2_uk_n99;
  output u0_FP_11, u0_FP_12, u0_FP_14, u0_FP_19, u0_FP_22, u0_FP_25, u0_FP_29, u0_FP_3, u0_FP_32, 
        u0_FP_4, u0_FP_7, u0_FP_8, u0_N0, u0_N1, u0_N12, u0_N128, u0_N129, u0_N133, 
        u0_N137, u0_N140, u0_N143, u0_N145, u0_N147, u0_N151, u0_N153, u0_N155, u0_N157, 
        u0_N16, u0_N17, u0_N19, u0_N194, u0_N195, u0_N198, u0_N199, u0_N202, u0_N203, 
        u0_N205, u0_N210, u0_N213, u0_N216, u0_N22, u0_N220, u0_N223, u0_N25, u0_N256, 
        u0_N258, u0_N260, u0_N263, u0_N265, u0_N269, u0_N27, u0_N270, u0_N275, u0_N276, 
        u0_N280, u0_N281, u0_N282, u0_N30, u0_N386, u0_N387, u0_N390, u0_N391, u0_N394, 
        u0_N395, u0_N397, u0_N402, u0_N405, u0_N408, u0_N412, u0_N415, u0_N8, u0_N9, 
        u0_uk_n117, u0_uk_n155, u0_uk_n187, u0_uk_n230, u0_uk_n674, u0_uk_n684, u0_uk_n690, u0_uk_n696, u0_uk_n697, 
        u0_uk_n698, u0_uk_n705, u0_uk_n790, u0_uk_n871, u0_uk_n99, u2_N102, u2_N103, u2_N106, u2_N107, 
        u2_N109, u2_N114, u2_N117, u2_N120, u2_N124, u2_N127, u2_N161, u2_N164, u2_N168, 
        u2_N172, u2_N174, u2_N176, u2_N177, u2_N180, u2_N182, u2_N186, u2_N187, u2_N190, 
        u2_N320, u2_N321, u2_N325, u2_N328, u2_N329, u2_N332, u2_N335, u2_N336, u2_N337, 
        u2_N339, u2_N342, u2_N343, u2_N345, u2_N347, u2_N349, u2_N350, u2_N384, u2_N386, 
        u2_N387, u2_N391, u2_N393, u2_N394, u2_N397, u2_N402, u2_N403, u2_N408, u2_N409, 
        u2_N412, u2_N418, u2_N423, u2_N429, u2_N440, u2_N64, u2_N66, u2_N67, u2_N68, 
        u2_N70, u2_N71, u2_N73, u2_N74, u2_N75, u2_N77, u2_N78, u2_N82, u2_N83, 
        u2_N84, u2_N85, u2_N88, u2_N89, u2_N90, u2_N92, u2_N95, u2_N98, u2_N99, 
        u2_uk_n1039, u2_uk_n1056, u2_uk_n230, u2_uk_n672;
  wire u0_K13_25, u0_K13_26, u0_K13_27, u0_K13_28, u0_K13_29, u0_K13_31, u0_K13_32, u0_K13_33, u0_K13_34, 
       u0_K13_35, u0_K13_37, u0_K13_38, u0_K13_41, u0_K16_25, u0_K16_27, u0_K16_28, u0_K16_29, u0_K16_30, 
       u0_K16_31, u0_K16_32, u0_K16_33, u0_K16_34, u0_K16_35, u0_K16_36, u0_K16_37, u0_K16_39, u0_K16_40, 
       u0_K16_41, u0_K16_42, u0_K1_1, u0_K1_10, u0_K1_11, u0_K1_12, u0_K1_19, u0_K1_2, u0_K1_20, 
       u0_K1_21, u0_K1_22, u0_K1_24, u0_K1_3, u0_K1_4, u0_K1_5, u0_K1_6, u0_K1_7, u0_K1_8, 
       u0_K1_9, u0_K5_10, u0_K5_11, u0_K5_12, u0_K5_17, u0_K5_20, u0_K5_21, u0_K5_22, u0_K5_7, 
       u0_K5_8, u0_K7_25, u0_K7_26, u0_K7_27, u0_K7_28, u0_K7_29, u0_K7_30, u0_K7_31, u0_K7_32, 
       u0_K7_33, u0_K7_34, u0_K7_35, u0_K7_36, u0_K7_37, u0_K7_38, u0_K7_39, u0_K7_40, u0_K7_41, 
       u0_K7_42, u0_K9_19, u0_K9_20, u0_K9_21, u0_K9_22, u0_K9_23, u0_K9_24, u0_K9_25, u0_K9_26, 
       u0_K9_27, u0_K9_28, u0_K9_29, u0_K9_30, u0_K9_43, u0_K9_44, u0_K9_46, u0_K9_47, u0_K9_48, 
       u0_out0_1, u0_out0_10, u0_out0_13, u0_out0_17, u0_out0_18, u0_out0_2, u0_out0_20, u0_out0_23, u0_out0_26, 
       u0_out0_28, u0_out0_31, u0_out0_9, u0_out12_11, u0_out12_12, u0_out12_14, u0_out12_19, u0_out12_22, u0_out12_25, 
       u0_out12_29, u0_out12_3, u0_out12_32, u0_out12_4, u0_out12_7, u0_out12_8, u0_out15_11, u0_out15_12, u0_out15_14, 
       u0_out15_19, u0_out15_22, u0_out15_25, u0_out15_29, u0_out15_3, u0_out15_32, u0_out15_4, u0_out15_7, u0_out15_8, 
       u0_out4_1, u0_out4_10, u0_out4_13, u0_out4_16, u0_out4_18, u0_out4_2, u0_out4_20, u0_out4_24, u0_out4_26, 
       u0_out4_28, u0_out4_30, u0_out4_6, u0_out6_11, u0_out6_12, u0_out6_14, u0_out6_19, u0_out6_22, u0_out6_25, 
       u0_out6_29, u0_out6_3, u0_out6_32, u0_out6_4, u0_out6_7, u0_out6_8, u0_out8_1, u0_out8_10, u0_out8_14, 
       u0_out8_15, u0_out8_20, u0_out8_21, u0_out8_25, u0_out8_26, u0_out8_27, u0_out8_3, u0_out8_5, u0_out8_8, 
       u0_u0_X_1, u0_u0_X_10, u0_u0_X_11, u0_u0_X_12, u0_u0_X_19, u0_u0_X_2, u0_u0_X_20, u0_u0_X_21, u0_u0_X_22, 
       u0_u0_X_23, u0_u0_X_24, u0_u0_X_3, u0_u0_X_4, u0_u0_X_5, u0_u0_X_6, u0_u0_X_7, u0_u0_X_8, u0_u0_X_9, 
       u0_u0_u0_n1, u0_u0_u0_n10, u0_u0_u0_n11, u0_u0_u0_n12, u0_u0_u0_n13, u0_u0_u0_n14, u0_u0_u0_n15, u0_u0_u0_n16, u0_u0_u0_n17, 
       u0_u0_u0_n18, u0_u0_u0_n19, u0_u0_u0_n2, u0_u0_u0_n20, u0_u0_u0_n21, u0_u0_u0_n22, u0_u0_u0_n23, u0_u0_u0_n24, u0_u0_u0_n25, 
       u0_u0_u0_n26, u0_u0_u0_n27, u0_u0_u0_n28, u0_u0_u0_n29, u0_u0_u0_n3, u0_u0_u0_n30, u0_u0_u0_n31, u0_u0_u0_n32, u0_u0_u0_n33, 
       u0_u0_u0_n34, u0_u0_u0_n35, u0_u0_u0_n36, u0_u0_u0_n37, u0_u0_u0_n38, u0_u0_u0_n39, u0_u0_u0_n4, u0_u0_u0_n40, u0_u0_u0_n41, 
       u0_u0_u0_n42, u0_u0_u0_n43, u0_u0_u0_n44, u0_u0_u0_n45, u0_u0_u0_n46, u0_u0_u0_n47, u0_u0_u0_n48, u0_u0_u0_n49, u0_u0_u0_n5, 
       u0_u0_u0_n50, u0_u0_u0_n51, u0_u0_u0_n52, u0_u0_u0_n53, u0_u0_u0_n54, u0_u0_u0_n55, u0_u0_u0_n56, u0_u0_u0_n57, u0_u0_u0_n58, 
       u0_u0_u0_n59, u0_u0_u0_n6, u0_u0_u0_n60, u0_u0_u0_n61, u0_u0_u0_n62, u0_u0_u0_n63, u0_u0_u0_n64, u0_u0_u0_n65, u0_u0_u0_n66, 
       u0_u0_u0_n67, u0_u0_u0_n68, u0_u0_u0_n69, u0_u0_u0_n7, u0_u0_u0_n70, u0_u0_u0_n71, u0_u0_u0_n72, u0_u0_u0_n73, u0_u0_u0_n74, 
       u0_u0_u0_n75, u0_u0_u0_n76, u0_u0_u0_n77, u0_u0_u0_n78, u0_u0_u0_n79, u0_u0_u0_n8, u0_u0_u0_n80, u0_u0_u0_n81, u0_u0_u0_n82, 
       u0_u0_u0_n83, u0_u0_u0_n84, u0_u0_u0_n85, u0_u0_u0_n86, u0_u0_u0_n87, u0_u0_u0_n9, u0_u0_u1_n1, u0_u0_u1_n10, u0_u0_u1_n11, 
       u0_u0_u1_n12, u0_u0_u1_n13, u0_u0_u1_n14, u0_u0_u1_n15, u0_u0_u1_n16, u0_u0_u1_n17, u0_u0_u1_n18, u0_u0_u1_n19, u0_u0_u1_n2, 
       u0_u0_u1_n20, u0_u0_u1_n21, u0_u0_u1_n22, u0_u0_u1_n23, u0_u0_u1_n24, u0_u0_u1_n25, u0_u0_u1_n26, u0_u0_u1_n27, u0_u0_u1_n28, 
       u0_u0_u1_n29, u0_u0_u1_n3, u0_u0_u1_n30, u0_u0_u1_n31, u0_u0_u1_n32, u0_u0_u1_n33, u0_u0_u1_n34, u0_u0_u1_n35, u0_u0_u1_n36, 
       u0_u0_u1_n37, u0_u0_u1_n38, u0_u0_u1_n39, u0_u0_u1_n4, u0_u0_u1_n40, u0_u0_u1_n41, u0_u0_u1_n42, u0_u0_u1_n43, u0_u0_u1_n44, 
       u0_u0_u1_n45, u0_u0_u1_n46, u0_u0_u1_n47, u0_u0_u1_n48, u0_u0_u1_n49, u0_u0_u1_n5, u0_u0_u1_n50, u0_u0_u1_n51, u0_u0_u1_n52, 
       u0_u0_u1_n53, u0_u0_u1_n54, u0_u0_u1_n55, u0_u0_u1_n56, u0_u0_u1_n57, u0_u0_u1_n58, u0_u0_u1_n59, u0_u0_u1_n6, u0_u0_u1_n60, 
       u0_u0_u1_n61, u0_u0_u1_n62, u0_u0_u1_n63, u0_u0_u1_n64, u0_u0_u1_n65, u0_u0_u1_n66, u0_u0_u1_n67, u0_u0_u1_n68, u0_u0_u1_n69, 
       u0_u0_u1_n7, u0_u0_u1_n70, u0_u0_u1_n71, u0_u0_u1_n72, u0_u0_u1_n73, u0_u0_u1_n74, u0_u0_u1_n75, u0_u0_u1_n76, u0_u0_u1_n77, 
       u0_u0_u1_n78, u0_u0_u1_n79, u0_u0_u1_n8, u0_u0_u1_n80, u0_u0_u1_n81, u0_u0_u1_n82, u0_u0_u1_n83, u0_u0_u1_n84, u0_u0_u1_n85, 
       u0_u0_u1_n86, u0_u0_u1_n87, u0_u0_u1_n88, u0_u0_u1_n89, u0_u0_u1_n9, u0_u0_u1_n90, u0_u0_u1_n91, u0_u0_u1_n92, u0_u0_u1_n93, 
       u0_u0_u1_n94, u0_u0_u3_n1, u0_u0_u3_n10, u0_u0_u3_n11, u0_u0_u3_n12, u0_u0_u3_n13, u0_u0_u3_n14, u0_u0_u3_n15, u0_u0_u3_n16, 
       u0_u0_u3_n17, u0_u0_u3_n18, u0_u0_u3_n19, u0_u0_u3_n2, u0_u0_u3_n20, u0_u0_u3_n21, u0_u0_u3_n22, u0_u0_u3_n23, u0_u0_u3_n24, 
       u0_u0_u3_n25, u0_u0_u3_n26, u0_u0_u3_n27, u0_u0_u3_n28, u0_u0_u3_n29, u0_u0_u3_n3, u0_u0_u3_n30, u0_u0_u3_n31, u0_u0_u3_n32, 
       u0_u0_u3_n33, u0_u0_u3_n34, u0_u0_u3_n35, u0_u0_u3_n36, u0_u0_u3_n37, u0_u0_u3_n38, u0_u0_u3_n39, u0_u0_u3_n4, u0_u0_u3_n40, 
       u0_u0_u3_n41, u0_u0_u3_n42, u0_u0_u3_n43, u0_u0_u3_n44, u0_u0_u3_n45, u0_u0_u3_n46, u0_u0_u3_n47, u0_u0_u3_n48, u0_u0_u3_n49, 
       u0_u0_u3_n5, u0_u0_u3_n50, u0_u0_u3_n51, u0_u0_u3_n52, u0_u0_u3_n53, u0_u0_u3_n54, u0_u0_u3_n55, u0_u0_u3_n56, u0_u0_u3_n57, 
       u0_u0_u3_n58, u0_u0_u3_n59, u0_u0_u3_n6, u0_u0_u3_n60, u0_u0_u3_n61, u0_u0_u3_n62, u0_u0_u3_n63, u0_u0_u3_n64, u0_u0_u3_n65, 
       u0_u0_u3_n66, u0_u0_u3_n67, u0_u0_u3_n68, u0_u0_u3_n69, u0_u0_u3_n7, u0_u0_u3_n70, u0_u0_u3_n71, u0_u0_u3_n72, u0_u0_u3_n73, 
       u0_u0_u3_n74, u0_u0_u3_n75, u0_u0_u3_n76, u0_u0_u3_n77, u0_u0_u3_n78, u0_u0_u3_n79, u0_u0_u3_n8, u0_u0_u3_n80, u0_u0_u3_n81, 
       u0_u0_u3_n82, u0_u0_u3_n83, u0_u0_u3_n84, u0_u0_u3_n85, u0_u0_u3_n86, u0_u0_u3_n87, u0_u0_u3_n88, u0_u0_u3_n89, u0_u0_u3_n9, 
       u0_u0_u3_n90, u0_u0_u3_n91, u0_u0_u3_n92, u0_u0_u3_n93, u0_u12_X_25, u0_u12_X_26, u0_u12_X_27, u0_u12_X_28, u0_u12_X_29, 
       u0_u12_X_30, u0_u12_X_31, u0_u12_X_32, u0_u12_X_33, u0_u12_X_34, u0_u12_X_35, u0_u12_X_36, u0_u12_X_37, u0_u12_X_38, 
       u0_u12_X_39, u0_u12_X_40, u0_u12_X_41, u0_u12_X_42, u0_u12_u4_n100, u0_u12_u4_n101, u0_u12_u4_n102, u0_u12_u4_n103, u0_u12_u4_n104, 
       u0_u12_u4_n105, u0_u12_u4_n106, u0_u12_u4_n107, u0_u12_u4_n108, u0_u12_u4_n109, u0_u12_u4_n110, u0_u12_u4_n111, u0_u12_u4_n112, u0_u12_u4_n113, 
       u0_u12_u4_n114, u0_u12_u4_n115, u0_u12_u4_n116, u0_u12_u4_n117, u0_u12_u4_n118, u0_u12_u4_n119, u0_u12_u4_n120, u0_u12_u4_n121, u0_u12_u4_n122, 
       u0_u12_u4_n123, u0_u12_u4_n124, u0_u12_u4_n125, u0_u12_u4_n126, u0_u12_u4_n127, u0_u12_u4_n128, u0_u12_u4_n129, u0_u12_u4_n130, u0_u12_u4_n131, 
       u0_u12_u4_n132, u0_u12_u4_n133, u0_u12_u4_n134, u0_u12_u4_n135, u0_u12_u4_n136, u0_u12_u4_n137, u0_u12_u4_n138, u0_u12_u4_n139, u0_u12_u4_n140, 
       u0_u12_u4_n141, u0_u12_u4_n142, u0_u12_u4_n143, u0_u12_u4_n144, u0_u12_u4_n145, u0_u12_u4_n146, u0_u12_u4_n147, u0_u12_u4_n148, u0_u12_u4_n149, 
       u0_u12_u4_n150, u0_u12_u4_n151, u0_u12_u4_n152, u0_u12_u4_n153, u0_u12_u4_n154, u0_u12_u4_n155, u0_u12_u4_n156, u0_u12_u4_n157, u0_u12_u4_n158, 
       u0_u12_u4_n159, u0_u12_u4_n160, u0_u12_u4_n161, u0_u12_u4_n162, u0_u12_u4_n163, u0_u12_u4_n164, u0_u12_u4_n165, u0_u12_u4_n166, u0_u12_u4_n167, 
       u0_u12_u4_n168, u0_u12_u4_n169, u0_u12_u4_n170, u0_u12_u4_n171, u0_u12_u4_n172, u0_u12_u4_n173, u0_u12_u4_n174, u0_u12_u4_n175, u0_u12_u4_n176, 
       u0_u12_u4_n177, u0_u12_u4_n178, u0_u12_u4_n179, u0_u12_u4_n180, u0_u12_u4_n181, u0_u12_u4_n182, u0_u12_u4_n183, u0_u12_u4_n184, u0_u12_u4_n185, 
       u0_u12_u4_n186, u0_u12_u4_n94, u0_u12_u4_n95, u0_u12_u4_n96, u0_u12_u4_n97, u0_u12_u4_n98, u0_u12_u4_n99, u0_u12_u5_n100, u0_u12_u5_n101, 
       u0_u12_u5_n102, u0_u12_u5_n103, u0_u12_u5_n104, u0_u12_u5_n105, u0_u12_u5_n106, u0_u12_u5_n107, u0_u12_u5_n108, u0_u12_u5_n109, u0_u12_u5_n110, 
       u0_u12_u5_n111, u0_u12_u5_n112, u0_u12_u5_n113, u0_u12_u5_n114, u0_u12_u5_n115, u0_u12_u5_n116, u0_u12_u5_n117, u0_u12_u5_n118, u0_u12_u5_n119, 
       u0_u12_u5_n120, u0_u12_u5_n121, u0_u12_u5_n122, u0_u12_u5_n123, u0_u12_u5_n124, u0_u12_u5_n125, u0_u12_u5_n126, u0_u12_u5_n127, u0_u12_u5_n128, 
       u0_u12_u5_n129, u0_u12_u5_n130, u0_u12_u5_n131, u0_u12_u5_n132, u0_u12_u5_n133, u0_u12_u5_n134, u0_u12_u5_n135, u0_u12_u5_n136, u0_u12_u5_n137, 
       u0_u12_u5_n138, u0_u12_u5_n139, u0_u12_u5_n140, u0_u12_u5_n141, u0_u12_u5_n142, u0_u12_u5_n143, u0_u12_u5_n144, u0_u12_u5_n145, u0_u12_u5_n146, 
       u0_u12_u5_n147, u0_u12_u5_n148, u0_u12_u5_n149, u0_u12_u5_n150, u0_u12_u5_n151, u0_u12_u5_n152, u0_u12_u5_n153, u0_u12_u5_n154, u0_u12_u5_n155, 
       u0_u12_u5_n156, u0_u12_u5_n157, u0_u12_u5_n158, u0_u12_u5_n159, u0_u12_u5_n160, u0_u12_u5_n161, u0_u12_u5_n162, u0_u12_u5_n163, u0_u12_u5_n164, 
       u0_u12_u5_n165, u0_u12_u5_n166, u0_u12_u5_n167, u0_u12_u5_n168, u0_u12_u5_n169, u0_u12_u5_n170, u0_u12_u5_n171, u0_u12_u5_n172, u0_u12_u5_n173, 
       u0_u12_u5_n174, u0_u12_u5_n175, u0_u12_u5_n176, u0_u12_u5_n177, u0_u12_u5_n178, u0_u12_u5_n179, u0_u12_u5_n180, u0_u12_u5_n181, u0_u12_u5_n182, 
       u0_u12_u5_n183, u0_u12_u5_n184, u0_u12_u5_n185, u0_u12_u5_n186, u0_u12_u5_n187, u0_u12_u5_n188, u0_u12_u5_n189, u0_u12_u5_n190, u0_u12_u5_n191, 
       u0_u12_u5_n192, u0_u12_u5_n193, u0_u12_u5_n194, u0_u12_u5_n195, u0_u12_u5_n196, u0_u12_u5_n99, u0_u12_u6_n100, u0_u12_u6_n101, u0_u12_u6_n102, 
       u0_u12_u6_n103, u0_u12_u6_n104, u0_u12_u6_n105, u0_u12_u6_n106, u0_u12_u6_n107, u0_u12_u6_n108, u0_u12_u6_n109, u0_u12_u6_n110, u0_u12_u6_n111, 
       u0_u12_u6_n112, u0_u12_u6_n113, u0_u12_u6_n114, u0_u12_u6_n115, u0_u12_u6_n116, u0_u12_u6_n117, u0_u12_u6_n118, u0_u12_u6_n119, u0_u12_u6_n120, 
       u0_u12_u6_n121, u0_u12_u6_n122, u0_u12_u6_n123, u0_u12_u6_n124, u0_u12_u6_n125, u0_u12_u6_n126, u0_u12_u6_n127, u0_u12_u6_n128, u0_u12_u6_n129, 
       u0_u12_u6_n130, u0_u12_u6_n131, u0_u12_u6_n132, u0_u12_u6_n133, u0_u12_u6_n134, u0_u12_u6_n135, u0_u12_u6_n136, u0_u12_u6_n137, u0_u12_u6_n138, 
       u0_u12_u6_n139, u0_u12_u6_n140, u0_u12_u6_n141, u0_u12_u6_n142, u0_u12_u6_n143, u0_u12_u6_n144, u0_u12_u6_n145, u0_u12_u6_n146, u0_u12_u6_n147, 
       u0_u12_u6_n148, u0_u12_u6_n149, u0_u12_u6_n150, u0_u12_u6_n151, u0_u12_u6_n152, u0_u12_u6_n153, u0_u12_u6_n154, u0_u12_u6_n155, u0_u12_u6_n156, 
       u0_u12_u6_n157, u0_u12_u6_n158, u0_u12_u6_n159, u0_u12_u6_n160, u0_u12_u6_n161, u0_u12_u6_n162, u0_u12_u6_n163, u0_u12_u6_n164, u0_u12_u6_n165, 
       u0_u12_u6_n166, u0_u12_u6_n167, u0_u12_u6_n168, u0_u12_u6_n169, u0_u12_u6_n170, u0_u12_u6_n171, u0_u12_u6_n172, u0_u12_u6_n173, u0_u12_u6_n174, 
       u0_u12_u6_n88, u0_u12_u6_n89, u0_u12_u6_n90, u0_u12_u6_n91, u0_u12_u6_n92, u0_u12_u6_n93, u0_u12_u6_n94, u0_u12_u6_n95, u0_u12_u6_n96, 
       u0_u12_u6_n97, u0_u12_u6_n98, u0_u12_u6_n99, u0_u15_X_25, u0_u15_X_26, u0_u15_X_27, u0_u15_X_28, u0_u15_X_29, u0_u15_X_30, 
       u0_u15_X_31, u0_u15_X_32, u0_u15_X_33, u0_u15_X_34, u0_u15_X_35, u0_u15_X_36, u0_u15_X_37, u0_u15_X_38, u0_u15_X_39, 
       u0_u15_X_40, u0_u15_X_41, u0_u15_X_42, u0_u15_u4_n100, u0_u15_u4_n101, u0_u15_u4_n102, u0_u15_u4_n103, u0_u15_u4_n104, u0_u15_u4_n105, 
       u0_u15_u4_n106, u0_u15_u4_n107, u0_u15_u4_n108, u0_u15_u4_n109, u0_u15_u4_n110, u0_u15_u4_n111, u0_u15_u4_n112, u0_u15_u4_n113, u0_u15_u4_n114, 
       u0_u15_u4_n115, u0_u15_u4_n116, u0_u15_u4_n117, u0_u15_u4_n118, u0_u15_u4_n119, u0_u15_u4_n120, u0_u15_u4_n121, u0_u15_u4_n122, u0_u15_u4_n123, 
       u0_u15_u4_n124, u0_u15_u4_n125, u0_u15_u4_n126, u0_u15_u4_n127, u0_u15_u4_n128, u0_u15_u4_n129, u0_u15_u4_n130, u0_u15_u4_n131, u0_u15_u4_n132, 
       u0_u15_u4_n133, u0_u15_u4_n134, u0_u15_u4_n135, u0_u15_u4_n136, u0_u15_u4_n137, u0_u15_u4_n138, u0_u15_u4_n139, u0_u15_u4_n140, u0_u15_u4_n141, 
       u0_u15_u4_n142, u0_u15_u4_n143, u0_u15_u4_n144, u0_u15_u4_n145, u0_u15_u4_n146, u0_u15_u4_n147, u0_u15_u4_n148, u0_u15_u4_n149, u0_u15_u4_n150, 
       u0_u15_u4_n151, u0_u15_u4_n152, u0_u15_u4_n153, u0_u15_u4_n154, u0_u15_u4_n155, u0_u15_u4_n156, u0_u15_u4_n157, u0_u15_u4_n158, u0_u15_u4_n159, 
       u0_u15_u4_n160, u0_u15_u4_n161, u0_u15_u4_n162, u0_u15_u4_n163, u0_u15_u4_n164, u0_u15_u4_n165, u0_u15_u4_n166, u0_u15_u4_n167, u0_u15_u4_n168, 
       u0_u15_u4_n169, u0_u15_u4_n170, u0_u15_u4_n171, u0_u15_u4_n172, u0_u15_u4_n173, u0_u15_u4_n174, u0_u15_u4_n175, u0_u15_u4_n176, u0_u15_u4_n177, 
       u0_u15_u4_n178, u0_u15_u4_n179, u0_u15_u4_n180, u0_u15_u4_n181, u0_u15_u4_n182, u0_u15_u4_n183, u0_u15_u4_n184, u0_u15_u4_n185, u0_u15_u4_n186, 
       u0_u15_u4_n94, u0_u15_u4_n95, u0_u15_u4_n96, u0_u15_u4_n97, u0_u15_u4_n98, u0_u15_u4_n99, u0_u15_u5_n100, u0_u15_u5_n101, u0_u15_u5_n102, 
       u0_u15_u5_n103, u0_u15_u5_n104, u0_u15_u5_n105, u0_u15_u5_n106, u0_u15_u5_n107, u0_u15_u5_n108, u0_u15_u5_n109, u0_u15_u5_n110, u0_u15_u5_n111, 
       u0_u15_u5_n112, u0_u15_u5_n113, u0_u15_u5_n114, u0_u15_u5_n115, u0_u15_u5_n116, u0_u15_u5_n117, u0_u15_u5_n118, u0_u15_u5_n119, u0_u15_u5_n120, 
       u0_u15_u5_n121, u0_u15_u5_n122, u0_u15_u5_n123, u0_u15_u5_n124, u0_u15_u5_n125, u0_u15_u5_n126, u0_u15_u5_n127, u0_u15_u5_n128, u0_u15_u5_n129, 
       u0_u15_u5_n130, u0_u15_u5_n131, u0_u15_u5_n132, u0_u15_u5_n133, u0_u15_u5_n134, u0_u15_u5_n135, u0_u15_u5_n136, u0_u15_u5_n137, u0_u15_u5_n138, 
       u0_u15_u5_n139, u0_u15_u5_n140, u0_u15_u5_n141, u0_u15_u5_n142, u0_u15_u5_n143, u0_u15_u5_n144, u0_u15_u5_n145, u0_u15_u5_n146, u0_u15_u5_n147, 
       u0_u15_u5_n148, u0_u15_u5_n149, u0_u15_u5_n150, u0_u15_u5_n151, u0_u15_u5_n152, u0_u15_u5_n153, u0_u15_u5_n154, u0_u15_u5_n155, u0_u15_u5_n156, 
       u0_u15_u5_n157, u0_u15_u5_n158, u0_u15_u5_n159, u0_u15_u5_n160, u0_u15_u5_n161, u0_u15_u5_n162, u0_u15_u5_n163, u0_u15_u5_n164, u0_u15_u5_n165, 
       u0_u15_u5_n166, u0_u15_u5_n167, u0_u15_u5_n168, u0_u15_u5_n169, u0_u15_u5_n170, u0_u15_u5_n171, u0_u15_u5_n172, u0_u15_u5_n173, u0_u15_u5_n174, 
       u0_u15_u5_n175, u0_u15_u5_n176, u0_u15_u5_n177, u0_u15_u5_n178, u0_u15_u5_n179, u0_u15_u5_n180, u0_u15_u5_n181, u0_u15_u5_n182, u0_u15_u5_n183, 
       u0_u15_u5_n184, u0_u15_u5_n185, u0_u15_u5_n186, u0_u15_u5_n187, u0_u15_u5_n188, u0_u15_u5_n189, u0_u15_u5_n190, u0_u15_u5_n191, u0_u15_u5_n192, 
       u0_u15_u5_n193, u0_u15_u5_n194, u0_u15_u5_n195, u0_u15_u5_n196, u0_u15_u5_n99, u0_u15_u6_n100, u0_u15_u6_n101, u0_u15_u6_n102, u0_u15_u6_n103, 
       u0_u15_u6_n104, u0_u15_u6_n105, u0_u15_u6_n106, u0_u15_u6_n107, u0_u15_u6_n108, u0_u15_u6_n109, u0_u15_u6_n110, u0_u15_u6_n111, u0_u15_u6_n112, 
       u0_u15_u6_n113, u0_u15_u6_n114, u0_u15_u6_n115, u0_u15_u6_n116, u0_u15_u6_n117, u0_u15_u6_n118, u0_u15_u6_n119, u0_u15_u6_n120, u0_u15_u6_n121, 
       u0_u15_u6_n122, u0_u15_u6_n123, u0_u15_u6_n124, u0_u15_u6_n125, u0_u15_u6_n126, u0_u15_u6_n127, u0_u15_u6_n128, u0_u15_u6_n129, u0_u15_u6_n130, 
       u0_u15_u6_n131, u0_u15_u6_n132, u0_u15_u6_n133, u0_u15_u6_n134, u0_u15_u6_n135, u0_u15_u6_n136, u0_u15_u6_n137, u0_u15_u6_n138, u0_u15_u6_n139, 
       u0_u15_u6_n140, u0_u15_u6_n141, u0_u15_u6_n142, u0_u15_u6_n143, u0_u15_u6_n144, u0_u15_u6_n145, u0_u15_u6_n146, u0_u15_u6_n147, u0_u15_u6_n148, 
       u0_u15_u6_n149, u0_u15_u6_n150, u0_u15_u6_n151, u0_u15_u6_n152, u0_u15_u6_n153, u0_u15_u6_n154, u0_u15_u6_n155, u0_u15_u6_n156, u0_u15_u6_n157, 
       u0_u15_u6_n158, u0_u15_u6_n159, u0_u15_u6_n160, u0_u15_u6_n161, u0_u15_u6_n162, u0_u15_u6_n163, u0_u15_u6_n164, u0_u15_u6_n165, u0_u15_u6_n166, 
       u0_u15_u6_n167, u0_u15_u6_n168, u0_u15_u6_n169, u0_u15_u6_n170, u0_u15_u6_n171, u0_u15_u6_n172, u0_u15_u6_n173, u0_u15_u6_n174, u0_u15_u6_n88, 
       u0_u15_u6_n89, u0_u15_u6_n90, u0_u15_u6_n91, u0_u15_u6_n92, u0_u15_u6_n93, u0_u15_u6_n94, u0_u15_u6_n95, u0_u15_u6_n96, u0_u15_u6_n97, 
       u0_u15_u6_n98, u0_u15_u6_n99, u0_u4_X_10, u0_u4_X_11, u0_u4_X_12, u0_u4_X_13, u0_u4_X_14, u0_u4_X_15, u0_u4_X_16, 
       u0_u4_X_17, u0_u4_X_18, u0_u4_X_19, u0_u4_X_20, u0_u4_X_21, u0_u4_X_22, u0_u4_X_23, u0_u4_X_24, u0_u4_X_7, 
       u0_u4_X_8, u0_u4_X_9, u0_u4_u1_n100, u0_u4_u1_n101, u0_u4_u1_n102, u0_u4_u1_n103, u0_u4_u1_n104, u0_u4_u1_n105, u0_u4_u1_n106, 
       u0_u4_u1_n107, u0_u4_u1_n108, u0_u4_u1_n109, u0_u4_u1_n110, u0_u4_u1_n111, u0_u4_u1_n112, u0_u4_u1_n113, u0_u4_u1_n114, u0_u4_u1_n115, 
       u0_u4_u1_n116, u0_u4_u1_n117, u0_u4_u1_n118, u0_u4_u1_n119, u0_u4_u1_n120, u0_u4_u1_n121, u0_u4_u1_n122, u0_u4_u1_n123, u0_u4_u1_n124, 
       u0_u4_u1_n125, u0_u4_u1_n126, u0_u4_u1_n127, u0_u4_u1_n128, u0_u4_u1_n129, u0_u4_u1_n130, u0_u4_u1_n131, u0_u4_u1_n132, u0_u4_u1_n133, 
       u0_u4_u1_n134, u0_u4_u1_n135, u0_u4_u1_n136, u0_u4_u1_n137, u0_u4_u1_n138, u0_u4_u1_n139, u0_u4_u1_n140, u0_u4_u1_n141, u0_u4_u1_n142, 
       u0_u4_u1_n143, u0_u4_u1_n144, u0_u4_u1_n145, u0_u4_u1_n146, u0_u4_u1_n147, u0_u4_u1_n148, u0_u4_u1_n149, u0_u4_u1_n150, u0_u4_u1_n151, 
       u0_u4_u1_n152, u0_u4_u1_n153, u0_u4_u1_n154, u0_u4_u1_n155, u0_u4_u1_n156, u0_u4_u1_n157, u0_u4_u1_n158, u0_u4_u1_n159, u0_u4_u1_n160, 
       u0_u4_u1_n161, u0_u4_u1_n162, u0_u4_u1_n163, u0_u4_u1_n164, u0_u4_u1_n165, u0_u4_u1_n166, u0_u4_u1_n167, u0_u4_u1_n168, u0_u4_u1_n169, 
       u0_u4_u1_n170, u0_u4_u1_n171, u0_u4_u1_n172, u0_u4_u1_n173, u0_u4_u1_n174, u0_u4_u1_n175, u0_u4_u1_n176, u0_u4_u1_n177, u0_u4_u1_n178, 
       u0_u4_u1_n179, u0_u4_u1_n180, u0_u4_u1_n181, u0_u4_u1_n182, u0_u4_u1_n183, u0_u4_u1_n184, u0_u4_u1_n185, u0_u4_u1_n186, u0_u4_u1_n187, 
       u0_u4_u1_n188, u0_u4_u1_n95, u0_u4_u1_n96, u0_u4_u1_n97, u0_u4_u1_n98, u0_u4_u1_n99, u0_u4_u2_n100, u0_u4_u2_n101, u0_u4_u2_n102, 
       u0_u4_u2_n103, u0_u4_u2_n104, u0_u4_u2_n105, u0_u4_u2_n106, u0_u4_u2_n107, u0_u4_u2_n108, u0_u4_u2_n109, u0_u4_u2_n110, u0_u4_u2_n111, 
       u0_u4_u2_n112, u0_u4_u2_n113, u0_u4_u2_n114, u0_u4_u2_n115, u0_u4_u2_n116, u0_u4_u2_n117, u0_u4_u2_n118, u0_u4_u2_n119, u0_u4_u2_n120, 
       u0_u4_u2_n121, u0_u4_u2_n122, u0_u4_u2_n123, u0_u4_u2_n124, u0_u4_u2_n125, u0_u4_u2_n126, u0_u4_u2_n127, u0_u4_u2_n128, u0_u4_u2_n129, 
       u0_u4_u2_n130, u0_u4_u2_n131, u0_u4_u2_n132, u0_u4_u2_n133, u0_u4_u2_n134, u0_u4_u2_n135, u0_u4_u2_n136, u0_u4_u2_n137, u0_u4_u2_n138, 
       u0_u4_u2_n139, u0_u4_u2_n140, u0_u4_u2_n141, u0_u4_u2_n142, u0_u4_u2_n143, u0_u4_u2_n144, u0_u4_u2_n145, u0_u4_u2_n146, u0_u4_u2_n147, 
       u0_u4_u2_n148, u0_u4_u2_n149, u0_u4_u2_n150, u0_u4_u2_n151, u0_u4_u2_n152, u0_u4_u2_n153, u0_u4_u2_n154, u0_u4_u2_n155, u0_u4_u2_n156, 
       u0_u4_u2_n157, u0_u4_u2_n158, u0_u4_u2_n159, u0_u4_u2_n160, u0_u4_u2_n161, u0_u4_u2_n162, u0_u4_u2_n163, u0_u4_u2_n164, u0_u4_u2_n165, 
       u0_u4_u2_n166, u0_u4_u2_n167, u0_u4_u2_n168, u0_u4_u2_n169, u0_u4_u2_n170, u0_u4_u2_n171, u0_u4_u2_n172, u0_u4_u2_n173, u0_u4_u2_n174, 
       u0_u4_u2_n175, u0_u4_u2_n176, u0_u4_u2_n177, u0_u4_u2_n178, u0_u4_u2_n179, u0_u4_u2_n180, u0_u4_u2_n181, u0_u4_u2_n182, u0_u4_u2_n183, 
       u0_u4_u2_n184, u0_u4_u2_n185, u0_u4_u2_n186, u0_u4_u2_n187, u0_u4_u2_n188, u0_u4_u2_n95, u0_u4_u2_n96, u0_u4_u2_n97, u0_u4_u2_n98, 
       u0_u4_u2_n99, u0_u4_u3_n100, u0_u4_u3_n101, u0_u4_u3_n102, u0_u4_u3_n103, u0_u4_u3_n104, u0_u4_u3_n105, u0_u4_u3_n106, u0_u4_u3_n107, 
       u0_u4_u3_n108, u0_u4_u3_n109, u0_u4_u3_n110, u0_u4_u3_n111, u0_u4_u3_n112, u0_u4_u3_n113, u0_u4_u3_n114, u0_u4_u3_n115, u0_u4_u3_n116, 
       u0_u4_u3_n117, u0_u4_u3_n118, u0_u4_u3_n119, u0_u4_u3_n120, u0_u4_u3_n121, u0_u4_u3_n122, u0_u4_u3_n123, u0_u4_u3_n124, u0_u4_u3_n125, 
       u0_u4_u3_n126, u0_u4_u3_n127, u0_u4_u3_n128, u0_u4_u3_n129, u0_u4_u3_n130, u0_u4_u3_n131, u0_u4_u3_n132, u0_u4_u3_n133, u0_u4_u3_n134, 
       u0_u4_u3_n135, u0_u4_u3_n136, u0_u4_u3_n137, u0_u4_u3_n138, u0_u4_u3_n139, u0_u4_u3_n140, u0_u4_u3_n141, u0_u4_u3_n142, u0_u4_u3_n143, 
       u0_u4_u3_n144, u0_u4_u3_n145, u0_u4_u3_n146, u0_u4_u3_n147, u0_u4_u3_n148, u0_u4_u3_n149, u0_u4_u3_n150, u0_u4_u3_n151, u0_u4_u3_n152, 
       u0_u4_u3_n153, u0_u4_u3_n154, u0_u4_u3_n155, u0_u4_u3_n156, u0_u4_u3_n157, u0_u4_u3_n158, u0_u4_u3_n159, u0_u4_u3_n160, u0_u4_u3_n161, 
       u0_u4_u3_n162, u0_u4_u3_n163, u0_u4_u3_n164, u0_u4_u3_n165, u0_u4_u3_n166, u0_u4_u3_n167, u0_u4_u3_n168, u0_u4_u3_n169, u0_u4_u3_n170, 
       u0_u4_u3_n171, u0_u4_u3_n172, u0_u4_u3_n173, u0_u4_u3_n174, u0_u4_u3_n175, u0_u4_u3_n176, u0_u4_u3_n177, u0_u4_u3_n178, u0_u4_u3_n179, 
       u0_u4_u3_n180, u0_u4_u3_n181, u0_u4_u3_n182, u0_u4_u3_n183, u0_u4_u3_n184, u0_u4_u3_n185, u0_u4_u3_n186, u0_u4_u3_n94, u0_u4_u3_n95, 
       u0_u4_u3_n96, u0_u4_u3_n97, u0_u4_u3_n98, u0_u4_u3_n99, u0_u6_X_25, u0_u6_X_26, u0_u6_X_27, u0_u6_X_28, u0_u6_X_29, 
       u0_u6_X_30, u0_u6_X_31, u0_u6_X_32, u0_u6_X_33, u0_u6_X_34, u0_u6_X_35, u0_u6_X_36, u0_u6_X_37, u0_u6_X_38, 
       u0_u6_X_39, u0_u6_X_40, u0_u6_X_41, u0_u6_X_42, u0_u6_u4_n100, u0_u6_u4_n101, u0_u6_u4_n102, u0_u6_u4_n103, u0_u6_u4_n104, 
       u0_u6_u4_n105, u0_u6_u4_n106, u0_u6_u4_n107, u0_u6_u4_n108, u0_u6_u4_n109, u0_u6_u4_n110, u0_u6_u4_n111, u0_u6_u4_n112, u0_u6_u4_n113, 
       u0_u6_u4_n114, u0_u6_u4_n115, u0_u6_u4_n116, u0_u6_u4_n117, u0_u6_u4_n118, u0_u6_u4_n119, u0_u6_u4_n120, u0_u6_u4_n121, u0_u6_u4_n122, 
       u0_u6_u4_n123, u0_u6_u4_n124, u0_u6_u4_n125, u0_u6_u4_n126, u0_u6_u4_n127, u0_u6_u4_n128, u0_u6_u4_n129, u0_u6_u4_n130, u0_u6_u4_n131, 
       u0_u6_u4_n132, u0_u6_u4_n133, u0_u6_u4_n134, u0_u6_u4_n135, u0_u6_u4_n136, u0_u6_u4_n137, u0_u6_u4_n138, u0_u6_u4_n139, u0_u6_u4_n140, 
       u0_u6_u4_n141, u0_u6_u4_n142, u0_u6_u4_n143, u0_u6_u4_n144, u0_u6_u4_n145, u0_u6_u4_n146, u0_u6_u4_n147, u0_u6_u4_n148, u0_u6_u4_n149, 
       u0_u6_u4_n150, u0_u6_u4_n151, u0_u6_u4_n152, u0_u6_u4_n153, u0_u6_u4_n154, u0_u6_u4_n155, u0_u6_u4_n156, u0_u6_u4_n157, u0_u6_u4_n158, 
       u0_u6_u4_n159, u0_u6_u4_n160, u0_u6_u4_n161, u0_u6_u4_n162, u0_u6_u4_n163, u0_u6_u4_n164, u0_u6_u4_n165, u0_u6_u4_n166, u0_u6_u4_n167, 
       u0_u6_u4_n168, u0_u6_u4_n169, u0_u6_u4_n170, u0_u6_u4_n171, u0_u6_u4_n172, u0_u6_u4_n173, u0_u6_u4_n174, u0_u6_u4_n175, u0_u6_u4_n176, 
       u0_u6_u4_n177, u0_u6_u4_n178, u0_u6_u4_n179, u0_u6_u4_n180, u0_u6_u4_n181, u0_u6_u4_n182, u0_u6_u4_n183, u0_u6_u4_n184, u0_u6_u4_n185, 
       u0_u6_u4_n186, u0_u6_u4_n94, u0_u6_u4_n95, u0_u6_u4_n96, u0_u6_u4_n97, u0_u6_u4_n98, u0_u6_u4_n99, u0_u6_u5_n100, u0_u6_u5_n101, 
       u0_u6_u5_n102, u0_u6_u5_n103, u0_u6_u5_n104, u0_u6_u5_n105, u0_u6_u5_n106, u0_u6_u5_n107, u0_u6_u5_n108, u0_u6_u5_n109, u0_u6_u5_n110, 
       u0_u6_u5_n111, u0_u6_u5_n112, u0_u6_u5_n113, u0_u6_u5_n114, u0_u6_u5_n115, u0_u6_u5_n116, u0_u6_u5_n117, u0_u6_u5_n118, u0_u6_u5_n119, 
       u0_u6_u5_n120, u0_u6_u5_n121, u0_u6_u5_n122, u0_u6_u5_n123, u0_u6_u5_n124, u0_u6_u5_n125, u0_u6_u5_n126, u0_u6_u5_n127, u0_u6_u5_n128, 
       u0_u6_u5_n129, u0_u6_u5_n130, u0_u6_u5_n131, u0_u6_u5_n132, u0_u6_u5_n133, u0_u6_u5_n134, u0_u6_u5_n135, u0_u6_u5_n136, u0_u6_u5_n137, 
       u0_u6_u5_n138, u0_u6_u5_n139, u0_u6_u5_n140, u0_u6_u5_n141, u0_u6_u5_n142, u0_u6_u5_n143, u0_u6_u5_n144, u0_u6_u5_n145, u0_u6_u5_n146, 
       u0_u6_u5_n147, u0_u6_u5_n148, u0_u6_u5_n149, u0_u6_u5_n150, u0_u6_u5_n151, u0_u6_u5_n152, u0_u6_u5_n153, u0_u6_u5_n154, u0_u6_u5_n155, 
       u0_u6_u5_n156, u0_u6_u5_n157, u0_u6_u5_n158, u0_u6_u5_n159, u0_u6_u5_n160, u0_u6_u5_n161, u0_u6_u5_n162, u0_u6_u5_n163, u0_u6_u5_n164, 
       u0_u6_u5_n165, u0_u6_u5_n166, u0_u6_u5_n167, u0_u6_u5_n168, u0_u6_u5_n169, u0_u6_u5_n170, u0_u6_u5_n171, u0_u6_u5_n172, u0_u6_u5_n173, 
       u0_u6_u5_n174, u0_u6_u5_n175, u0_u6_u5_n176, u0_u6_u5_n177, u0_u6_u5_n178, u0_u6_u5_n179, u0_u6_u5_n180, u0_u6_u5_n181, u0_u6_u5_n182, 
       u0_u6_u5_n183, u0_u6_u5_n184, u0_u6_u5_n185, u0_u6_u5_n186, u0_u6_u5_n187, u0_u6_u5_n188, u0_u6_u5_n189, u0_u6_u5_n190, u0_u6_u5_n191, 
       u0_u6_u5_n192, u0_u6_u5_n193, u0_u6_u5_n194, u0_u6_u5_n195, u0_u6_u5_n196, u0_u6_u5_n99, u0_u6_u6_n100, u0_u6_u6_n101, u0_u6_u6_n102, 
       u0_u6_u6_n103, u0_u6_u6_n104, u0_u6_u6_n105, u0_u6_u6_n106, u0_u6_u6_n107, u0_u6_u6_n108, u0_u6_u6_n109, u0_u6_u6_n110, u0_u6_u6_n111, 
       u0_u6_u6_n112, u0_u6_u6_n113, u0_u6_u6_n114, u0_u6_u6_n115, u0_u6_u6_n116, u0_u6_u6_n117, u0_u6_u6_n118, u0_u6_u6_n119, u0_u6_u6_n120, 
       u0_u6_u6_n121, u0_u6_u6_n122, u0_u6_u6_n123, u0_u6_u6_n124, u0_u6_u6_n125, u0_u6_u6_n126, u0_u6_u6_n127, u0_u6_u6_n128, u0_u6_u6_n129, 
       u0_u6_u6_n130, u0_u6_u6_n131, u0_u6_u6_n132, u0_u6_u6_n133, u0_u6_u6_n134, u0_u6_u6_n135, u0_u6_u6_n136, u0_u6_u6_n137, u0_u6_u6_n138, 
       u0_u6_u6_n139, u0_u6_u6_n140, u0_u6_u6_n141, u0_u6_u6_n142, u0_u6_u6_n143, u0_u6_u6_n144, u0_u6_u6_n145, u0_u6_u6_n146, u0_u6_u6_n147, 
       u0_u6_u6_n148, u0_u6_u6_n149, u0_u6_u6_n150, u0_u6_u6_n151, u0_u6_u6_n152, u0_u6_u6_n153, u0_u6_u6_n154, u0_u6_u6_n155, u0_u6_u6_n156, 
       u0_u6_u6_n157, u0_u6_u6_n158, u0_u6_u6_n159, u0_u6_u6_n160, u0_u6_u6_n161, u0_u6_u6_n162, u0_u6_u6_n163, u0_u6_u6_n164, u0_u6_u6_n165, 
       u0_u6_u6_n166, u0_u6_u6_n167, u0_u6_u6_n168, u0_u6_u6_n169, u0_u6_u6_n170, u0_u6_u6_n171, u0_u6_u6_n172, u0_u6_u6_n173, u0_u6_u6_n174, 
       u0_u6_u6_n88, u0_u6_u6_n89, u0_u6_u6_n90, u0_u6_u6_n91, u0_u6_u6_n92, u0_u6_u6_n93, u0_u6_u6_n94, u0_u6_u6_n95, u0_u6_u6_n96, 
       u0_u6_u6_n97, u0_u6_u6_n98, u0_u6_u6_n99, u0_u8_X_19, u0_u8_X_20, u0_u8_X_21, u0_u8_X_22, u0_u8_X_23, u0_u8_X_24, 
       u0_u8_X_25, u0_u8_X_26, u0_u8_X_27, u0_u8_X_28, u0_u8_X_29, u0_u8_X_30, u0_u8_X_43, u0_u8_X_44, u0_u8_X_45, 
       u0_u8_X_46, u0_u8_X_47, u0_u8_X_48, u0_u8_u3_n100, u0_u8_u3_n101, u0_u8_u3_n102, u0_u8_u3_n103, u0_u8_u3_n104, u0_u8_u3_n105, 
       u0_u8_u3_n106, u0_u8_u3_n107, u0_u8_u3_n108, u0_u8_u3_n109, u0_u8_u3_n110, u0_u8_u3_n111, u0_u8_u3_n112, u0_u8_u3_n113, u0_u8_u3_n114, 
       u0_u8_u3_n115, u0_u8_u3_n116, u0_u8_u3_n117, u0_u8_u3_n118, u0_u8_u3_n119, u0_u8_u3_n120, u0_u8_u3_n121, u0_u8_u3_n122, u0_u8_u3_n123, 
       u0_u8_u3_n124, u0_u8_u3_n125, u0_u8_u3_n126, u0_u8_u3_n127, u0_u8_u3_n128, u0_u8_u3_n129, u0_u8_u3_n130, u0_u8_u3_n131, u0_u8_u3_n132, 
       u0_u8_u3_n133, u0_u8_u3_n134, u0_u8_u3_n135, u0_u8_u3_n136, u0_u8_u3_n137, u0_u8_u3_n138, u0_u8_u3_n139, u0_u8_u3_n140, u0_u8_u3_n141, 
       u0_u8_u3_n142, u0_u8_u3_n143, u0_u8_u3_n144, u0_u8_u3_n145, u0_u8_u3_n146, u0_u8_u3_n147, u0_u8_u3_n148, u0_u8_u3_n149, u0_u8_u3_n150, 
       u0_u8_u3_n151, u0_u8_u3_n152, u0_u8_u3_n153, u0_u8_u3_n154, u0_u8_u3_n155, u0_u8_u3_n156, u0_u8_u3_n157, u0_u8_u3_n158, u0_u8_u3_n159, 
       u0_u8_u3_n160, u0_u8_u3_n161, u0_u8_u3_n162, u0_u8_u3_n163, u0_u8_u3_n164, u0_u8_u3_n165, u0_u8_u3_n166, u0_u8_u3_n167, u0_u8_u3_n168, 
       u0_u8_u3_n169, u0_u8_u3_n170, u0_u8_u3_n171, u0_u8_u3_n172, u0_u8_u3_n173, u0_u8_u3_n174, u0_u8_u3_n175, u0_u8_u3_n176, u0_u8_u3_n177, 
       u0_u8_u3_n178, u0_u8_u3_n179, u0_u8_u3_n180, u0_u8_u3_n181, u0_u8_u3_n182, u0_u8_u3_n183, u0_u8_u3_n184, u0_u8_u3_n185, u0_u8_u3_n186, 
       u0_u8_u3_n94, u0_u8_u3_n95, u0_u8_u3_n96, u0_u8_u3_n97, u0_u8_u3_n98, u0_u8_u3_n99, u0_u8_u4_n100, u0_u8_u4_n101, u0_u8_u4_n102, 
       u0_u8_u4_n103, u0_u8_u4_n104, u0_u8_u4_n105, u0_u8_u4_n106, u0_u8_u4_n107, u0_u8_u4_n108, u0_u8_u4_n109, u0_u8_u4_n110, u0_u8_u4_n111, 
       u0_u8_u4_n112, u0_u8_u4_n113, u0_u8_u4_n114, u0_u8_u4_n115, u0_u8_u4_n116, u0_u8_u4_n117, u0_u8_u4_n118, u0_u8_u4_n119, u0_u8_u4_n120, 
       u0_u8_u4_n121, u0_u8_u4_n122, u0_u8_u4_n123, u0_u8_u4_n124, u0_u8_u4_n125, u0_u8_u4_n126, u0_u8_u4_n127, u0_u8_u4_n128, u0_u8_u4_n129, 
       u0_u8_u4_n130, u0_u8_u4_n131, u0_u8_u4_n132, u0_u8_u4_n133, u0_u8_u4_n134, u0_u8_u4_n135, u0_u8_u4_n136, u0_u8_u4_n137, u0_u8_u4_n138, 
       u0_u8_u4_n139, u0_u8_u4_n140, u0_u8_u4_n141, u0_u8_u4_n142, u0_u8_u4_n143, u0_u8_u4_n144, u0_u8_u4_n145, u0_u8_u4_n146, u0_u8_u4_n147, 
       u0_u8_u4_n148, u0_u8_u4_n149, u0_u8_u4_n150, u0_u8_u4_n151, u0_u8_u4_n152, u0_u8_u4_n153, u0_u8_u4_n154, u0_u8_u4_n155, u0_u8_u4_n156, 
       u0_u8_u4_n157, u0_u8_u4_n158, u0_u8_u4_n159, u0_u8_u4_n160, u0_u8_u4_n161, u0_u8_u4_n162, u0_u8_u4_n163, u0_u8_u4_n164, u0_u8_u4_n165, 
       u0_u8_u4_n166, u0_u8_u4_n167, u0_u8_u4_n168, u0_u8_u4_n169, u0_u8_u4_n170, u0_u8_u4_n171, u0_u8_u4_n172, u0_u8_u4_n173, u0_u8_u4_n174, 
       u0_u8_u4_n175, u0_u8_u4_n176, u0_u8_u4_n177, u0_u8_u4_n178, u0_u8_u4_n179, u0_u8_u4_n180, u0_u8_u4_n181, u0_u8_u4_n182, u0_u8_u4_n183, 
       u0_u8_u4_n184, u0_u8_u4_n185, u0_u8_u4_n186, u0_u8_u4_n94, u0_u8_u4_n95, u0_u8_u4_n96, u0_u8_u4_n97, u0_u8_u4_n98, u0_u8_u4_n99, 
       u0_u8_u7_n100, u0_u8_u7_n101, u0_u8_u7_n102, u0_u8_u7_n103, u0_u8_u7_n104, u0_u8_u7_n105, u0_u8_u7_n106, u0_u8_u7_n107, u0_u8_u7_n108, 
       u0_u8_u7_n109, u0_u8_u7_n110, u0_u8_u7_n111, u0_u8_u7_n112, u0_u8_u7_n113, u0_u8_u7_n114, u0_u8_u7_n115, u0_u8_u7_n116, u0_u8_u7_n117, 
       u0_u8_u7_n118, u0_u8_u7_n119, u0_u8_u7_n120, u0_u8_u7_n121, u0_u8_u7_n122, u0_u8_u7_n123, u0_u8_u7_n124, u0_u8_u7_n125, u0_u8_u7_n126, 
       u0_u8_u7_n127, u0_u8_u7_n128, u0_u8_u7_n129, u0_u8_u7_n130, u0_u8_u7_n131, u0_u8_u7_n132, u0_u8_u7_n133, u0_u8_u7_n134, u0_u8_u7_n135, 
       u0_u8_u7_n136, u0_u8_u7_n137, u0_u8_u7_n138, u0_u8_u7_n139, u0_u8_u7_n140, u0_u8_u7_n141, u0_u8_u7_n142, u0_u8_u7_n143, u0_u8_u7_n144, 
       u0_u8_u7_n145, u0_u8_u7_n146, u0_u8_u7_n147, u0_u8_u7_n148, u0_u8_u7_n149, u0_u8_u7_n150, u0_u8_u7_n151, u0_u8_u7_n152, u0_u8_u7_n153, 
       u0_u8_u7_n154, u0_u8_u7_n155, u0_u8_u7_n156, u0_u8_u7_n157, u0_u8_u7_n158, u0_u8_u7_n159, u0_u8_u7_n160, u0_u8_u7_n161, u0_u8_u7_n162, 
       u0_u8_u7_n163, u0_u8_u7_n164, u0_u8_u7_n165, u0_u8_u7_n166, u0_u8_u7_n167, u0_u8_u7_n168, u0_u8_u7_n169, u0_u8_u7_n170, u0_u8_u7_n171, 
       u0_u8_u7_n172, u0_u8_u7_n173, u0_u8_u7_n174, u0_u8_u7_n175, u0_u8_u7_n176, u0_u8_u7_n177, u0_u8_u7_n178, u0_u8_u7_n179, u0_u8_u7_n180, 
       u0_u8_u7_n91, u0_u8_u7_n92, u0_u8_u7_n93, u0_u8_u7_n94, u0_u8_u7_n95, u0_u8_u7_n96, u0_u8_u7_n97, u0_u8_u7_n98, u0_u8_u7_n99, 
       u0_uk_n673, u0_uk_n679, u0_uk_n683, u0_uk_n699, u0_uk_n703, u0_uk_n704, u0_uk_n708, u0_uk_n712, u0_uk_n713, 
       u0_uk_n721, u0_uk_n730, u0_uk_n733, u0_uk_n767, u0_uk_n768, u0_uk_n769, u0_uk_n771, u0_uk_n772, u0_uk_n774, 
       u0_uk_n802, u0_uk_n816, u0_uk_n818, u0_uk_n869, u0_uk_n881, u0_uk_n885, u0_uk_n886, u0_uk_n891, u0_uk_n892, 
       u0_uk_n893, u0_uk_n899, u0_uk_n900, u0_uk_n901, u0_uk_n902, u0_uk_n905, u0_uk_n947, u2_K11_1, u2_K11_10, 
       u2_K11_12, u2_K11_14, u2_K11_15, u2_K11_17, u2_K11_19, u2_K11_2, u2_K11_20, u2_K11_22, u2_K11_23, 
       u2_K11_24, u2_K11_3, u2_K11_5, u2_K11_8, u2_K13_19, u2_K13_21, u2_K13_22, u2_K13_23, u2_K13_24, 
       u2_K13_25, u2_K13_27, u2_K13_28, u2_K13_29, u2_K13_30, u2_K13_33, u2_K13_35, u2_K13_36, u2_K14_26, 
       u2_K14_27, u2_K14_29, u2_K14_30, u2_K3_19, u2_K3_21, u2_K3_22, u2_K3_24, u2_K3_25, u2_K3_26, 
       u2_K3_27, u2_K3_28, u2_K3_29, u2_K3_31, u2_K3_33, u2_K3_34, u2_K3_36, u2_K3_37, u2_K3_38, 
       u2_K3_39, u2_K3_40, u2_K3_41, u2_K3_44, u2_K3_45, u2_K3_46, u2_K4_25, u2_K4_26, u2_K4_28, 
       u2_K4_29, u2_K4_30, u2_K4_31, u2_K4_32, u2_K4_36, u2_K4_37, u2_K4_40, u2_K4_41, u2_K6_10, 
       u2_K6_12, u2_K6_2, u2_K6_4, u2_K6_43, u2_K6_44, u2_K6_45, u2_K6_46, u2_K6_47, u2_K6_48, 
       u2_K6_5, u2_K6_6, u2_K6_7, u2_K6_8, u2_K6_9, u2_out10_1, u2_out10_10, u2_out10_13, u2_out10_16, 
       u2_out10_17, u2_out10_18, u2_out10_2, u2_out10_20, u2_out10_23, u2_out10_24, u2_out10_26, u2_out10_28, u2_out10_30, 
       u2_out10_31, u2_out10_6, u2_out10_9, u2_out12_1, u2_out12_10, u2_out12_11, u2_out12_14, u2_out12_19, u2_out12_20, 
       u2_out12_25, u2_out12_26, u2_out12_29, u2_out12_3, u2_out12_4, u2_out12_8, u2_out13_14, u2_out13_25, u2_out13_3, 
       u2_out13_8, u2_out2_1, u2_out2_10, u2_out2_11, u2_out2_12, u2_out2_14, u2_out2_15, u2_out2_19, u2_out2_20, 
       u2_out2_21, u2_out2_22, u2_out2_25, u2_out2_26, u2_out2_27, u2_out2_29, u2_out2_3, u2_out2_32, u2_out2_4, 
       u2_out2_5, u2_out2_7, u2_out2_8, u2_out3_11, u2_out3_12, u2_out3_14, u2_out3_19, u2_out3_22, u2_out3_25, 
       u2_out3_29, u2_out3_3, u2_out3_32, u2_out3_4, u2_out3_7, u2_out3_8, u2_out5_13, u2_out5_15, u2_out5_17, 
       u2_out5_18, u2_out5_2, u2_out5_21, u2_out5_23, u2_out5_27, u2_out5_28, u2_out5_31, u2_out5_5, u2_out5_9, 
       u2_u10_X_1, u2_u10_X_10, u2_u10_X_11, u2_u10_X_12, u2_u10_X_13, u2_u10_X_14, u2_u10_X_15, u2_u10_X_16, u2_u10_X_17, 
       u2_u10_X_18, u2_u10_X_19, u2_u10_X_2, u2_u10_X_20, u2_u10_X_21, u2_u10_X_22, u2_u10_X_23, u2_u10_X_24, u2_u10_X_3, 
       u2_u10_X_4, u2_u10_X_5, u2_u10_X_6, u2_u10_X_7, u2_u10_X_8, u2_u10_X_9, u2_u10_u0_n100, u2_u10_u0_n101, u2_u10_u0_n102, 
       u2_u10_u0_n103, u2_u10_u0_n104, u2_u10_u0_n105, u2_u10_u0_n106, u2_u10_u0_n107, u2_u10_u0_n108, u2_u10_u0_n109, u2_u10_u0_n110, u2_u10_u0_n111, 
       u2_u10_u0_n112, u2_u10_u0_n113, u2_u10_u0_n114, u2_u10_u0_n115, u2_u10_u0_n116, u2_u10_u0_n117, u2_u10_u0_n118, u2_u10_u0_n119, u2_u10_u0_n120, 
       u2_u10_u0_n121, u2_u10_u0_n122, u2_u10_u0_n123, u2_u10_u0_n124, u2_u10_u0_n125, u2_u10_u0_n126, u2_u10_u0_n127, u2_u10_u0_n128, u2_u10_u0_n129, 
       u2_u10_u0_n130, u2_u10_u0_n131, u2_u10_u0_n132, u2_u10_u0_n133, u2_u10_u0_n134, u2_u10_u0_n135, u2_u10_u0_n136, u2_u10_u0_n137, u2_u10_u0_n138, 
       u2_u10_u0_n139, u2_u10_u0_n140, u2_u10_u0_n141, u2_u10_u0_n142, u2_u10_u0_n143, u2_u10_u0_n144, u2_u10_u0_n145, u2_u10_u0_n146, u2_u10_u0_n147, 
       u2_u10_u0_n148, u2_u10_u0_n149, u2_u10_u0_n150, u2_u10_u0_n151, u2_u10_u0_n152, u2_u10_u0_n153, u2_u10_u0_n154, u2_u10_u0_n155, u2_u10_u0_n156, 
       u2_u10_u0_n157, u2_u10_u0_n158, u2_u10_u0_n159, u2_u10_u0_n160, u2_u10_u0_n161, u2_u10_u0_n162, u2_u10_u0_n163, u2_u10_u0_n164, u2_u10_u0_n165, 
       u2_u10_u0_n166, u2_u10_u0_n167, u2_u10_u0_n168, u2_u10_u0_n169, u2_u10_u0_n170, u2_u10_u0_n171, u2_u10_u0_n172, u2_u10_u0_n173, u2_u10_u0_n174, 
       u2_u10_u0_n88, u2_u10_u0_n89, u2_u10_u0_n90, u2_u10_u0_n91, u2_u10_u0_n92, u2_u10_u0_n93, u2_u10_u0_n94, u2_u10_u0_n95, u2_u10_u0_n96, 
       u2_u10_u0_n97, u2_u10_u0_n98, u2_u10_u0_n99, u2_u10_u1_n100, u2_u10_u1_n101, u2_u10_u1_n102, u2_u10_u1_n103, u2_u10_u1_n104, u2_u10_u1_n105, 
       u2_u10_u1_n106, u2_u10_u1_n107, u2_u10_u1_n108, u2_u10_u1_n109, u2_u10_u1_n110, u2_u10_u1_n111, u2_u10_u1_n112, u2_u10_u1_n113, u2_u10_u1_n114, 
       u2_u10_u1_n115, u2_u10_u1_n116, u2_u10_u1_n117, u2_u10_u1_n118, u2_u10_u1_n119, u2_u10_u1_n120, u2_u10_u1_n121, u2_u10_u1_n122, u2_u10_u1_n123, 
       u2_u10_u1_n124, u2_u10_u1_n125, u2_u10_u1_n126, u2_u10_u1_n127, u2_u10_u1_n128, u2_u10_u1_n129, u2_u10_u1_n130, u2_u10_u1_n131, u2_u10_u1_n132, 
       u2_u10_u1_n133, u2_u10_u1_n134, u2_u10_u1_n135, u2_u10_u1_n136, u2_u10_u1_n137, u2_u10_u1_n138, u2_u10_u1_n139, u2_u10_u1_n140, u2_u10_u1_n141, 
       u2_u10_u1_n142, u2_u10_u1_n143, u2_u10_u1_n144, u2_u10_u1_n145, u2_u10_u1_n146, u2_u10_u1_n147, u2_u10_u1_n148, u2_u10_u1_n149, u2_u10_u1_n150, 
       u2_u10_u1_n151, u2_u10_u1_n152, u2_u10_u1_n153, u2_u10_u1_n154, u2_u10_u1_n155, u2_u10_u1_n156, u2_u10_u1_n157, u2_u10_u1_n158, u2_u10_u1_n159, 
       u2_u10_u1_n160, u2_u10_u1_n161, u2_u10_u1_n162, u2_u10_u1_n163, u2_u10_u1_n164, u2_u10_u1_n165, u2_u10_u1_n166, u2_u10_u1_n167, u2_u10_u1_n168, 
       u2_u10_u1_n169, u2_u10_u1_n170, u2_u10_u1_n171, u2_u10_u1_n172, u2_u10_u1_n173, u2_u10_u1_n174, u2_u10_u1_n175, u2_u10_u1_n176, u2_u10_u1_n177, 
       u2_u10_u1_n178, u2_u10_u1_n179, u2_u10_u1_n180, u2_u10_u1_n181, u2_u10_u1_n182, u2_u10_u1_n183, u2_u10_u1_n184, u2_u10_u1_n185, u2_u10_u1_n186, 
       u2_u10_u1_n187, u2_u10_u1_n188, u2_u10_u1_n95, u2_u10_u1_n96, u2_u10_u1_n97, u2_u10_u1_n98, u2_u10_u1_n99, u2_u10_u2_n100, u2_u10_u2_n101, 
       u2_u10_u2_n102, u2_u10_u2_n103, u2_u10_u2_n104, u2_u10_u2_n105, u2_u10_u2_n106, u2_u10_u2_n107, u2_u10_u2_n108, u2_u10_u2_n109, u2_u10_u2_n110, 
       u2_u10_u2_n111, u2_u10_u2_n112, u2_u10_u2_n113, u2_u10_u2_n114, u2_u10_u2_n115, u2_u10_u2_n116, u2_u10_u2_n117, u2_u10_u2_n118, u2_u10_u2_n119, 
       u2_u10_u2_n120, u2_u10_u2_n121, u2_u10_u2_n122, u2_u10_u2_n123, u2_u10_u2_n124, u2_u10_u2_n125, u2_u10_u2_n126, u2_u10_u2_n127, u2_u10_u2_n128, 
       u2_u10_u2_n129, u2_u10_u2_n130, u2_u10_u2_n131, u2_u10_u2_n132, u2_u10_u2_n133, u2_u10_u2_n134, u2_u10_u2_n135, u2_u10_u2_n136, u2_u10_u2_n137, 
       u2_u10_u2_n138, u2_u10_u2_n139, u2_u10_u2_n140, u2_u10_u2_n141, u2_u10_u2_n142, u2_u10_u2_n143, u2_u10_u2_n144, u2_u10_u2_n145, u2_u10_u2_n146, 
       u2_u10_u2_n147, u2_u10_u2_n148, u2_u10_u2_n149, u2_u10_u2_n150, u2_u10_u2_n151, u2_u10_u2_n152, u2_u10_u2_n153, u2_u10_u2_n154, u2_u10_u2_n155, 
       u2_u10_u2_n156, u2_u10_u2_n157, u2_u10_u2_n158, u2_u10_u2_n159, u2_u10_u2_n160, u2_u10_u2_n161, u2_u10_u2_n162, u2_u10_u2_n163, u2_u10_u2_n164, 
       u2_u10_u2_n165, u2_u10_u2_n166, u2_u10_u2_n167, u2_u10_u2_n168, u2_u10_u2_n169, u2_u10_u2_n170, u2_u10_u2_n171, u2_u10_u2_n172, u2_u10_u2_n173, 
       u2_u10_u2_n174, u2_u10_u2_n175, u2_u10_u2_n176, u2_u10_u2_n177, u2_u10_u2_n178, u2_u10_u2_n179, u2_u10_u2_n180, u2_u10_u2_n181, u2_u10_u2_n182, 
       u2_u10_u2_n183, u2_u10_u2_n184, u2_u10_u2_n185, u2_u10_u2_n186, u2_u10_u2_n187, u2_u10_u2_n188, u2_u10_u2_n95, u2_u10_u2_n96, u2_u10_u2_n97, 
       u2_u10_u2_n98, u2_u10_u2_n99, u2_u10_u3_n100, u2_u10_u3_n101, u2_u10_u3_n102, u2_u10_u3_n103, u2_u10_u3_n104, u2_u10_u3_n105, u2_u10_u3_n106, 
       u2_u10_u3_n107, u2_u10_u3_n108, u2_u10_u3_n109, u2_u10_u3_n110, u2_u10_u3_n111, u2_u10_u3_n112, u2_u10_u3_n113, u2_u10_u3_n114, u2_u10_u3_n115, 
       u2_u10_u3_n116, u2_u10_u3_n117, u2_u10_u3_n118, u2_u10_u3_n119, u2_u10_u3_n120, u2_u10_u3_n121, u2_u10_u3_n122, u2_u10_u3_n123, u2_u10_u3_n124, 
       u2_u10_u3_n125, u2_u10_u3_n126, u2_u10_u3_n127, u2_u10_u3_n128, u2_u10_u3_n129, u2_u10_u3_n130, u2_u10_u3_n131, u2_u10_u3_n132, u2_u10_u3_n133, 
       u2_u10_u3_n134, u2_u10_u3_n135, u2_u10_u3_n136, u2_u10_u3_n137, u2_u10_u3_n138, u2_u10_u3_n139, u2_u10_u3_n140, u2_u10_u3_n141, u2_u10_u3_n142, 
       u2_u10_u3_n143, u2_u10_u3_n144, u2_u10_u3_n145, u2_u10_u3_n146, u2_u10_u3_n147, u2_u10_u3_n148, u2_u10_u3_n149, u2_u10_u3_n150, u2_u10_u3_n151, 
       u2_u10_u3_n152, u2_u10_u3_n153, u2_u10_u3_n154, u2_u10_u3_n155, u2_u10_u3_n156, u2_u10_u3_n157, u2_u10_u3_n158, u2_u10_u3_n159, u2_u10_u3_n160, 
       u2_u10_u3_n161, u2_u10_u3_n162, u2_u10_u3_n163, u2_u10_u3_n164, u2_u10_u3_n165, u2_u10_u3_n166, u2_u10_u3_n167, u2_u10_u3_n168, u2_u10_u3_n169, 
       u2_u10_u3_n170, u2_u10_u3_n171, u2_u10_u3_n172, u2_u10_u3_n173, u2_u10_u3_n174, u2_u10_u3_n175, u2_u10_u3_n176, u2_u10_u3_n177, u2_u10_u3_n178, 
       u2_u10_u3_n179, u2_u10_u3_n180, u2_u10_u3_n181, u2_u10_u3_n182, u2_u10_u3_n183, u2_u10_u3_n184, u2_u10_u3_n185, u2_u10_u3_n186, u2_u10_u3_n94, 
       u2_u10_u3_n95, u2_u10_u3_n96, u2_u10_u3_n97, u2_u10_u3_n98, u2_u10_u3_n99, u2_u12_X_19, u2_u12_X_20, u2_u12_X_21, u2_u12_X_22, 
       u2_u12_X_23, u2_u12_X_24, u2_u12_X_25, u2_u12_X_26, u2_u12_X_27, u2_u12_X_28, u2_u12_X_29, u2_u12_X_30, u2_u12_X_31, 
       u2_u12_X_32, u2_u12_X_33, u2_u12_X_34, u2_u12_X_35, u2_u12_X_36, u2_u12_u3_n100, u2_u12_u3_n101, u2_u12_u3_n102, u2_u12_u3_n103, 
       u2_u12_u3_n104, u2_u12_u3_n105, u2_u12_u3_n106, u2_u12_u3_n107, u2_u12_u3_n108, u2_u12_u3_n109, u2_u12_u3_n110, u2_u12_u3_n111, u2_u12_u3_n112, 
       u2_u12_u3_n113, u2_u12_u3_n114, u2_u12_u3_n115, u2_u12_u3_n116, u2_u12_u3_n117, u2_u12_u3_n118, u2_u12_u3_n119, u2_u12_u3_n120, u2_u12_u3_n121, 
       u2_u12_u3_n122, u2_u12_u3_n123, u2_u12_u3_n124, u2_u12_u3_n125, u2_u12_u3_n126, u2_u12_u3_n127, u2_u12_u3_n128, u2_u12_u3_n129, u2_u12_u3_n130, 
       u2_u12_u3_n131, u2_u12_u3_n132, u2_u12_u3_n133, u2_u12_u3_n134, u2_u12_u3_n135, u2_u12_u3_n136, u2_u12_u3_n137, u2_u12_u3_n138, u2_u12_u3_n139, 
       u2_u12_u3_n140, u2_u12_u3_n141, u2_u12_u3_n142, u2_u12_u3_n143, u2_u12_u3_n144, u2_u12_u3_n145, u2_u12_u3_n146, u2_u12_u3_n147, u2_u12_u3_n148, 
       u2_u12_u3_n149, u2_u12_u3_n150, u2_u12_u3_n151, u2_u12_u3_n152, u2_u12_u3_n153, u2_u12_u3_n154, u2_u12_u3_n155, u2_u12_u3_n156, u2_u12_u3_n157, 
       u2_u12_u3_n158, u2_u12_u3_n159, u2_u12_u3_n160, u2_u12_u3_n161, u2_u12_u3_n162, u2_u12_u3_n163, u2_u12_u3_n164, u2_u12_u3_n165, u2_u12_u3_n166, 
       u2_u12_u3_n167, u2_u12_u3_n168, u2_u12_u3_n169, u2_u12_u3_n170, u2_u12_u3_n171, u2_u12_u3_n172, u2_u12_u3_n173, u2_u12_u3_n174, u2_u12_u3_n175, 
       u2_u12_u3_n176, u2_u12_u3_n177, u2_u12_u3_n178, u2_u12_u3_n179, u2_u12_u3_n180, u2_u12_u3_n181, u2_u12_u3_n182, u2_u12_u3_n183, u2_u12_u3_n184, 
       u2_u12_u3_n185, u2_u12_u3_n186, u2_u12_u3_n94, u2_u12_u3_n95, u2_u12_u3_n96, u2_u12_u3_n97, u2_u12_u3_n98, u2_u12_u3_n99, u2_u12_u4_n100, 
       u2_u12_u4_n101, u2_u12_u4_n102, u2_u12_u4_n103, u2_u12_u4_n104, u2_u12_u4_n105, u2_u12_u4_n106, u2_u12_u4_n107, u2_u12_u4_n108, u2_u12_u4_n109, 
       u2_u12_u4_n110, u2_u12_u4_n111, u2_u12_u4_n112, u2_u12_u4_n113, u2_u12_u4_n114, u2_u12_u4_n115, u2_u12_u4_n116, u2_u12_u4_n117, u2_u12_u4_n118, 
       u2_u12_u4_n119, u2_u12_u4_n120, u2_u12_u4_n121, u2_u12_u4_n122, u2_u12_u4_n123, u2_u12_u4_n124, u2_u12_u4_n125, u2_u12_u4_n126, u2_u12_u4_n127, 
       u2_u12_u4_n128, u2_u12_u4_n129, u2_u12_u4_n130, u2_u12_u4_n131, u2_u12_u4_n132, u2_u12_u4_n133, u2_u12_u4_n134, u2_u12_u4_n135, u2_u12_u4_n136, 
       u2_u12_u4_n137, u2_u12_u4_n138, u2_u12_u4_n139, u2_u12_u4_n140, u2_u12_u4_n141, u2_u12_u4_n142, u2_u12_u4_n143, u2_u12_u4_n144, u2_u12_u4_n145, 
       u2_u12_u4_n146, u2_u12_u4_n147, u2_u12_u4_n148, u2_u12_u4_n149, u2_u12_u4_n150, u2_u12_u4_n151, u2_u12_u4_n152, u2_u12_u4_n153, u2_u12_u4_n154, 
       u2_u12_u4_n155, u2_u12_u4_n156, u2_u12_u4_n157, u2_u12_u4_n158, u2_u12_u4_n159, u2_u12_u4_n160, u2_u12_u4_n161, u2_u12_u4_n162, u2_u12_u4_n163, 
       u2_u12_u4_n164, u2_u12_u4_n165, u2_u12_u4_n166, u2_u12_u4_n167, u2_u12_u4_n168, u2_u12_u4_n169, u2_u12_u4_n170, u2_u12_u4_n171, u2_u12_u4_n172, 
       u2_u12_u4_n173, u2_u12_u4_n174, u2_u12_u4_n175, u2_u12_u4_n176, u2_u12_u4_n177, u2_u12_u4_n178, u2_u12_u4_n179, u2_u12_u4_n180, u2_u12_u4_n181, 
       u2_u12_u4_n182, u2_u12_u4_n183, u2_u12_u4_n184, u2_u12_u4_n185, u2_u12_u4_n186, u2_u12_u4_n94, u2_u12_u4_n95, u2_u12_u4_n96, u2_u12_u4_n97, 
       u2_u12_u4_n98, u2_u12_u4_n99, u2_u12_u5_n100, u2_u12_u5_n101, u2_u12_u5_n102, u2_u12_u5_n103, u2_u12_u5_n104, u2_u12_u5_n105, u2_u12_u5_n106, 
       u2_u12_u5_n107, u2_u12_u5_n108, u2_u12_u5_n109, u2_u12_u5_n110, u2_u12_u5_n111, u2_u12_u5_n112, u2_u12_u5_n113, u2_u12_u5_n114, u2_u12_u5_n115, 
       u2_u12_u5_n116, u2_u12_u5_n117, u2_u12_u5_n118, u2_u12_u5_n119, u2_u12_u5_n120, u2_u12_u5_n121, u2_u12_u5_n122, u2_u12_u5_n123, u2_u12_u5_n124, 
       u2_u12_u5_n125, u2_u12_u5_n126, u2_u12_u5_n127, u2_u12_u5_n128, u2_u12_u5_n129, u2_u12_u5_n130, u2_u12_u5_n131, u2_u12_u5_n132, u2_u12_u5_n133, 
       u2_u12_u5_n134, u2_u12_u5_n135, u2_u12_u5_n136, u2_u12_u5_n137, u2_u12_u5_n138, u2_u12_u5_n139, u2_u12_u5_n140, u2_u12_u5_n141, u2_u12_u5_n142, 
       u2_u12_u5_n143, u2_u12_u5_n144, u2_u12_u5_n145, u2_u12_u5_n146, u2_u12_u5_n147, u2_u12_u5_n148, u2_u12_u5_n149, u2_u12_u5_n150, u2_u12_u5_n151, 
       u2_u12_u5_n152, u2_u12_u5_n153, u2_u12_u5_n154, u2_u12_u5_n155, u2_u12_u5_n156, u2_u12_u5_n157, u2_u12_u5_n158, u2_u12_u5_n159, u2_u12_u5_n160, 
       u2_u12_u5_n161, u2_u12_u5_n162, u2_u12_u5_n163, u2_u12_u5_n164, u2_u12_u5_n165, u2_u12_u5_n166, u2_u12_u5_n167, u2_u12_u5_n168, u2_u12_u5_n169, 
       u2_u12_u5_n170, u2_u12_u5_n171, u2_u12_u5_n172, u2_u12_u5_n173, u2_u12_u5_n174, u2_u12_u5_n175, u2_u12_u5_n176, u2_u12_u5_n177, u2_u12_u5_n178, 
       u2_u12_u5_n179, u2_u12_u5_n180, u2_u12_u5_n181, u2_u12_u5_n182, u2_u12_u5_n183, u2_u12_u5_n184, u2_u12_u5_n185, u2_u12_u5_n186, u2_u12_u5_n187, 
       u2_u12_u5_n188, u2_u12_u5_n189, u2_u12_u5_n190, u2_u12_u5_n191, u2_u12_u5_n192, u2_u12_u5_n193, u2_u12_u5_n194, u2_u12_u5_n195, u2_u12_u5_n196, 
       u2_u12_u5_n99, u2_u13_X_25, u2_u13_X_26, u2_u13_X_27, u2_u13_X_28, u2_u13_X_29, u2_u13_X_30, u2_u13_u4_n100, u2_u13_u4_n101, 
       u2_u13_u4_n102, u2_u13_u4_n103, u2_u13_u4_n104, u2_u13_u4_n105, u2_u13_u4_n106, u2_u13_u4_n107, u2_u13_u4_n108, u2_u13_u4_n109, u2_u13_u4_n110, 
       u2_u13_u4_n111, u2_u13_u4_n112, u2_u13_u4_n113, u2_u13_u4_n114, u2_u13_u4_n115, u2_u13_u4_n116, u2_u13_u4_n117, u2_u13_u4_n118, u2_u13_u4_n119, 
       u2_u13_u4_n120, u2_u13_u4_n121, u2_u13_u4_n122, u2_u13_u4_n123, u2_u13_u4_n124, u2_u13_u4_n125, u2_u13_u4_n126, u2_u13_u4_n127, u2_u13_u4_n128, 
       u2_u13_u4_n129, u2_u13_u4_n130, u2_u13_u4_n131, u2_u13_u4_n132, u2_u13_u4_n133, u2_u13_u4_n134, u2_u13_u4_n135, u2_u13_u4_n136, u2_u13_u4_n137, 
       u2_u13_u4_n138, u2_u13_u4_n139, u2_u13_u4_n140, u2_u13_u4_n141, u2_u13_u4_n142, u2_u13_u4_n143, u2_u13_u4_n144, u2_u13_u4_n145, u2_u13_u4_n146, 
       u2_u13_u4_n147, u2_u13_u4_n148, u2_u13_u4_n149, u2_u13_u4_n150, u2_u13_u4_n151, u2_u13_u4_n152, u2_u13_u4_n153, u2_u13_u4_n154, u2_u13_u4_n155, 
       u2_u13_u4_n156, u2_u13_u4_n157, u2_u13_u4_n158, u2_u13_u4_n159, u2_u13_u4_n160, u2_u13_u4_n161, u2_u13_u4_n162, u2_u13_u4_n163, u2_u13_u4_n164, 
       u2_u13_u4_n165, u2_u13_u4_n166, u2_u13_u4_n167, u2_u13_u4_n168, u2_u13_u4_n169, u2_u13_u4_n170, u2_u13_u4_n171, u2_u13_u4_n172, u2_u13_u4_n173, 
       u2_u13_u4_n174, u2_u13_u4_n175, u2_u13_u4_n176, u2_u13_u4_n177, u2_u13_u4_n178, u2_u13_u4_n179, u2_u13_u4_n180, u2_u13_u4_n181, u2_u13_u4_n182, 
       u2_u13_u4_n183, u2_u13_u4_n184, u2_u13_u4_n185, u2_u13_u4_n186, u2_u13_u4_n94, u2_u13_u4_n95, u2_u13_u4_n96, u2_u13_u4_n97, u2_u13_u4_n98, 
       u2_u13_u4_n99, u2_u2_X_19, u2_u2_X_20, u2_u2_X_21, u2_u2_X_22, u2_u2_X_23, u2_u2_X_24, u2_u2_X_25, u2_u2_X_26, 
       u2_u2_X_27, u2_u2_X_28, u2_u2_X_29, u2_u2_X_30, u2_u2_X_31, u2_u2_X_32, u2_u2_X_33, u2_u2_X_34, u2_u2_X_35, 
       u2_u2_X_36, u2_u2_X_37, u2_u2_X_38, u2_u2_X_39, u2_u2_X_40, u2_u2_X_41, u2_u2_X_42, u2_u2_X_43, u2_u2_X_44, 
       u2_u2_X_45, u2_u2_X_46, u2_u2_X_47, u2_u2_X_48, u2_u2_u3_n100, u2_u2_u3_n101, u2_u2_u3_n102, u2_u2_u3_n103, u2_u2_u3_n104, 
       u2_u2_u3_n105, u2_u2_u3_n106, u2_u2_u3_n107, u2_u2_u3_n108, u2_u2_u3_n109, u2_u2_u3_n110, u2_u2_u3_n111, u2_u2_u3_n112, u2_u2_u3_n113, 
       u2_u2_u3_n114, u2_u2_u3_n115, u2_u2_u3_n116, u2_u2_u3_n117, u2_u2_u3_n118, u2_u2_u3_n119, u2_u2_u3_n120, u2_u2_u3_n121, u2_u2_u3_n122, 
       u2_u2_u3_n123, u2_u2_u3_n124, u2_u2_u3_n125, u2_u2_u3_n126, u2_u2_u3_n127, u2_u2_u3_n128, u2_u2_u3_n129, u2_u2_u3_n130, u2_u2_u3_n131, 
       u2_u2_u3_n132, u2_u2_u3_n133, u2_u2_u3_n134, u2_u2_u3_n135, u2_u2_u3_n136, u2_u2_u3_n137, u2_u2_u3_n138, u2_u2_u3_n139, u2_u2_u3_n140, 
       u2_u2_u3_n141, u2_u2_u3_n142, u2_u2_u3_n143, u2_u2_u3_n144, u2_u2_u3_n145, u2_u2_u3_n146, u2_u2_u3_n147, u2_u2_u3_n148, u2_u2_u3_n149, 
       u2_u2_u3_n150, u2_u2_u3_n151, u2_u2_u3_n152, u2_u2_u3_n153, u2_u2_u3_n154, u2_u2_u3_n155, u2_u2_u3_n156, u2_u2_u3_n157, u2_u2_u3_n158, 
       u2_u2_u3_n159, u2_u2_u3_n160, u2_u2_u3_n161, u2_u2_u3_n162, u2_u2_u3_n163, u2_u2_u3_n164, u2_u2_u3_n165, u2_u2_u3_n166, u2_u2_u3_n167, 
       u2_u2_u3_n168, u2_u2_u3_n169, u2_u2_u3_n170, u2_u2_u3_n171, u2_u2_u3_n172, u2_u2_u3_n173, u2_u2_u3_n174, u2_u2_u3_n175, u2_u2_u3_n176, 
       u2_u2_u3_n177, u2_u2_u3_n178, u2_u2_u3_n179, u2_u2_u3_n180, u2_u2_u3_n181, u2_u2_u3_n182, u2_u2_u3_n183, u2_u2_u3_n184, u2_u2_u3_n185, 
       u2_u2_u3_n186, u2_u2_u3_n94, u2_u2_u3_n95, u2_u2_u3_n96, u2_u2_u3_n97, u2_u2_u3_n98, u2_u2_u3_n99, u2_u2_u4_n100, u2_u2_u4_n101, 
       u2_u2_u4_n102, u2_u2_u4_n103, u2_u2_u4_n104, u2_u2_u4_n105, u2_u2_u4_n106, u2_u2_u4_n107, u2_u2_u4_n108, u2_u2_u4_n109, u2_u2_u4_n110, 
       u2_u2_u4_n111, u2_u2_u4_n112, u2_u2_u4_n113, u2_u2_u4_n114, u2_u2_u4_n115, u2_u2_u4_n116, u2_u2_u4_n117, u2_u2_u4_n118, u2_u2_u4_n119, 
       u2_u2_u4_n120, u2_u2_u4_n121, u2_u2_u4_n122, u2_u2_u4_n123, u2_u2_u4_n124, u2_u2_u4_n125, u2_u2_u4_n126, u2_u2_u4_n127, u2_u2_u4_n128, 
       u2_u2_u4_n129, u2_u2_u4_n130, u2_u2_u4_n131, u2_u2_u4_n132, u2_u2_u4_n133, u2_u2_u4_n134, u2_u2_u4_n135, u2_u2_u4_n136, u2_u2_u4_n137, 
       u2_u2_u4_n138, u2_u2_u4_n139, u2_u2_u4_n140, u2_u2_u4_n141, u2_u2_u4_n142, u2_u2_u4_n143, u2_u2_u4_n144, u2_u2_u4_n145, u2_u2_u4_n146, 
       u2_u2_u4_n147, u2_u2_u4_n148, u2_u2_u4_n149, u2_u2_u4_n150, u2_u2_u4_n151, u2_u2_u4_n152, u2_u2_u4_n153, u2_u2_u4_n154, u2_u2_u4_n155, 
       u2_u2_u4_n156, u2_u2_u4_n157, u2_u2_u4_n158, u2_u2_u4_n159, u2_u2_u4_n160, u2_u2_u4_n161, u2_u2_u4_n162, u2_u2_u4_n163, u2_u2_u4_n164, 
       u2_u2_u4_n165, u2_u2_u4_n166, u2_u2_u4_n167, u2_u2_u4_n168, u2_u2_u4_n169, u2_u2_u4_n170, u2_u2_u4_n171, u2_u2_u4_n172, u2_u2_u4_n173, 
       u2_u2_u4_n174, u2_u2_u4_n175, u2_u2_u4_n176, u2_u2_u4_n177, u2_u2_u4_n178, u2_u2_u4_n179, u2_u2_u4_n180, u2_u2_u4_n181, u2_u2_u4_n182, 
       u2_u2_u4_n183, u2_u2_u4_n184, u2_u2_u4_n185, u2_u2_u4_n186, u2_u2_u4_n94, u2_u2_u4_n95, u2_u2_u4_n96, u2_u2_u4_n97, u2_u2_u4_n98, 
       u2_u2_u4_n99, u2_u2_u5_n100, u2_u2_u5_n101, u2_u2_u5_n102, u2_u2_u5_n103, u2_u2_u5_n104, u2_u2_u5_n105, u2_u2_u5_n106, u2_u2_u5_n107, 
       u2_u2_u5_n108, u2_u2_u5_n109, u2_u2_u5_n110, u2_u2_u5_n111, u2_u2_u5_n112, u2_u2_u5_n113, u2_u2_u5_n114, u2_u2_u5_n115, u2_u2_u5_n116, 
       u2_u2_u5_n117, u2_u2_u5_n118, u2_u2_u5_n119, u2_u2_u5_n120, u2_u2_u5_n121, u2_u2_u5_n122, u2_u2_u5_n123, u2_u2_u5_n124, u2_u2_u5_n125, 
       u2_u2_u5_n126, u2_u2_u5_n127, u2_u2_u5_n128, u2_u2_u5_n129, u2_u2_u5_n130, u2_u2_u5_n131, u2_u2_u5_n132, u2_u2_u5_n133, u2_u2_u5_n134, 
       u2_u2_u5_n135, u2_u2_u5_n136, u2_u2_u5_n137, u2_u2_u5_n138, u2_u2_u5_n139, u2_u2_u5_n140, u2_u2_u5_n141, u2_u2_u5_n142, u2_u2_u5_n143, 
       u2_u2_u5_n144, u2_u2_u5_n145, u2_u2_u5_n146, u2_u2_u5_n147, u2_u2_u5_n148, u2_u2_u5_n149, u2_u2_u5_n150, u2_u2_u5_n151, u2_u2_u5_n152, 
       u2_u2_u5_n153, u2_u2_u5_n154, u2_u2_u5_n155, u2_u2_u5_n156, u2_u2_u5_n157, u2_u2_u5_n158, u2_u2_u5_n159, u2_u2_u5_n160, u2_u2_u5_n161, 
       u2_u2_u5_n162, u2_u2_u5_n163, u2_u2_u5_n164, u2_u2_u5_n165, u2_u2_u5_n166, u2_u2_u5_n167, u2_u2_u5_n168, u2_u2_u5_n169, u2_u2_u5_n170, 
       u2_u2_u5_n171, u2_u2_u5_n172, u2_u2_u5_n173, u2_u2_u5_n174, u2_u2_u5_n175, u2_u2_u5_n176, u2_u2_u5_n177, u2_u2_u5_n178, u2_u2_u5_n179, 
       u2_u2_u5_n180, u2_u2_u5_n181, u2_u2_u5_n182, u2_u2_u5_n183, u2_u2_u5_n184, u2_u2_u5_n185, u2_u2_u5_n186, u2_u2_u5_n187, u2_u2_u5_n188, 
       u2_u2_u5_n189, u2_u2_u5_n190, u2_u2_u5_n191, u2_u2_u5_n192, u2_u2_u5_n193, u2_u2_u5_n194, u2_u2_u5_n195, u2_u2_u5_n196, u2_u2_u5_n99, 
       u2_u2_u6_n100, u2_u2_u6_n101, u2_u2_u6_n102, u2_u2_u6_n103, u2_u2_u6_n104, u2_u2_u6_n105, u2_u2_u6_n106, u2_u2_u6_n107, u2_u2_u6_n108, 
       u2_u2_u6_n109, u2_u2_u6_n110, u2_u2_u6_n111, u2_u2_u6_n112, u2_u2_u6_n113, u2_u2_u6_n114, u2_u2_u6_n115, u2_u2_u6_n116, u2_u2_u6_n117, 
       u2_u2_u6_n118, u2_u2_u6_n119, u2_u2_u6_n120, u2_u2_u6_n121, u2_u2_u6_n122, u2_u2_u6_n123, u2_u2_u6_n124, u2_u2_u6_n125, u2_u2_u6_n126, 
       u2_u2_u6_n127, u2_u2_u6_n128, u2_u2_u6_n129, u2_u2_u6_n130, u2_u2_u6_n131, u2_u2_u6_n132, u2_u2_u6_n133, u2_u2_u6_n134, u2_u2_u6_n135, 
       u2_u2_u6_n136, u2_u2_u6_n137, u2_u2_u6_n138, u2_u2_u6_n139, u2_u2_u6_n140, u2_u2_u6_n141, u2_u2_u6_n142, u2_u2_u6_n143, u2_u2_u6_n144, 
       u2_u2_u6_n145, u2_u2_u6_n146, u2_u2_u6_n147, u2_u2_u6_n148, u2_u2_u6_n149, u2_u2_u6_n150, u2_u2_u6_n151, u2_u2_u6_n152, u2_u2_u6_n153, 
       u2_u2_u6_n154, u2_u2_u6_n155, u2_u2_u6_n156, u2_u2_u6_n157, u2_u2_u6_n158, u2_u2_u6_n159, u2_u2_u6_n160, u2_u2_u6_n161, u2_u2_u6_n162, 
       u2_u2_u6_n163, u2_u2_u6_n164, u2_u2_u6_n165, u2_u2_u6_n166, u2_u2_u6_n167, u2_u2_u6_n168, u2_u2_u6_n169, u2_u2_u6_n170, u2_u2_u6_n171, 
       u2_u2_u6_n172, u2_u2_u6_n173, u2_u2_u6_n174, u2_u2_u6_n88, u2_u2_u6_n89, u2_u2_u6_n90, u2_u2_u6_n91, u2_u2_u6_n92, u2_u2_u6_n93, 
       u2_u2_u6_n94, u2_u2_u6_n95, u2_u2_u6_n96, u2_u2_u6_n97, u2_u2_u6_n98, u2_u2_u6_n99, u2_u2_u7_n100, u2_u2_u7_n101, u2_u2_u7_n102, 
       u2_u2_u7_n103, u2_u2_u7_n104, u2_u2_u7_n105, u2_u2_u7_n106, u2_u2_u7_n107, u2_u2_u7_n108, u2_u2_u7_n109, u2_u2_u7_n110, u2_u2_u7_n111, 
       u2_u2_u7_n112, u2_u2_u7_n113, u2_u2_u7_n114, u2_u2_u7_n115, u2_u2_u7_n116, u2_u2_u7_n117, u2_u2_u7_n118, u2_u2_u7_n119, u2_u2_u7_n120, 
       u2_u2_u7_n121, u2_u2_u7_n122, u2_u2_u7_n123, u2_u2_u7_n124, u2_u2_u7_n125, u2_u2_u7_n126, u2_u2_u7_n127, u2_u2_u7_n128, u2_u2_u7_n129, 
       u2_u2_u7_n130, u2_u2_u7_n131, u2_u2_u7_n132, u2_u2_u7_n133, u2_u2_u7_n134, u2_u2_u7_n135, u2_u2_u7_n136, u2_u2_u7_n137, u2_u2_u7_n138, 
       u2_u2_u7_n139, u2_u2_u7_n140, u2_u2_u7_n141, u2_u2_u7_n142, u2_u2_u7_n143, u2_u2_u7_n144, u2_u2_u7_n145, u2_u2_u7_n146, u2_u2_u7_n147, 
       u2_u2_u7_n148, u2_u2_u7_n149, u2_u2_u7_n150, u2_u2_u7_n151, u2_u2_u7_n152, u2_u2_u7_n153, u2_u2_u7_n154, u2_u2_u7_n155, u2_u2_u7_n156, 
       u2_u2_u7_n157, u2_u2_u7_n158, u2_u2_u7_n159, u2_u2_u7_n160, u2_u2_u7_n161, u2_u2_u7_n162, u2_u2_u7_n163, u2_u2_u7_n164, u2_u2_u7_n165, 
       u2_u2_u7_n166, u2_u2_u7_n167, u2_u2_u7_n168, u2_u2_u7_n169, u2_u2_u7_n170, u2_u2_u7_n171, u2_u2_u7_n172, u2_u2_u7_n173, u2_u2_u7_n174, 
       u2_u2_u7_n175, u2_u2_u7_n176, u2_u2_u7_n177, u2_u2_u7_n178, u2_u2_u7_n179, u2_u2_u7_n180, u2_u2_u7_n91, u2_u2_u7_n92, u2_u2_u7_n93, 
       u2_u2_u7_n94, u2_u2_u7_n95, u2_u2_u7_n96, u2_u2_u7_n97, u2_u2_u7_n98, u2_u2_u7_n99, u2_u3_X_25, u2_u3_X_26, u2_u3_X_27, 
       u2_u3_X_28, u2_u3_X_29, u2_u3_X_30, u2_u3_X_31, u2_u3_X_32, u2_u3_X_33, u2_u3_X_34, u2_u3_X_35, u2_u3_X_36, 
       u2_u3_X_37, u2_u3_X_38, u2_u3_X_39, u2_u3_X_40, u2_u3_X_41, u2_u3_X_42, u2_u3_u4_n100, u2_u3_u4_n101, u2_u3_u4_n102, 
       u2_u3_u4_n103, u2_u3_u4_n104, u2_u3_u4_n105, u2_u3_u4_n106, u2_u3_u4_n107, u2_u3_u4_n108, u2_u3_u4_n109, u2_u3_u4_n110, u2_u3_u4_n111, 
       u2_u3_u4_n112, u2_u3_u4_n113, u2_u3_u4_n114, u2_u3_u4_n115, u2_u3_u4_n116, u2_u3_u4_n117, u2_u3_u4_n118, u2_u3_u4_n119, u2_u3_u4_n120, 
       u2_u3_u4_n121, u2_u3_u4_n122, u2_u3_u4_n123, u2_u3_u4_n124, u2_u3_u4_n125, u2_u3_u4_n126, u2_u3_u4_n127, u2_u3_u4_n128, u2_u3_u4_n129, 
       u2_u3_u4_n130, u2_u3_u4_n131, u2_u3_u4_n132, u2_u3_u4_n133, u2_u3_u4_n134, u2_u3_u4_n135, u2_u3_u4_n136, u2_u3_u4_n137, u2_u3_u4_n138, 
       u2_u3_u4_n139, u2_u3_u4_n140, u2_u3_u4_n141, u2_u3_u4_n142, u2_u3_u4_n143, u2_u3_u4_n144, u2_u3_u4_n145, u2_u3_u4_n146, u2_u3_u4_n147, 
       u2_u3_u4_n148, u2_u3_u4_n149, u2_u3_u4_n150, u2_u3_u4_n151, u2_u3_u4_n152, u2_u3_u4_n153, u2_u3_u4_n154, u2_u3_u4_n155, u2_u3_u4_n156, 
       u2_u3_u4_n157, u2_u3_u4_n158, u2_u3_u4_n159, u2_u3_u4_n160, u2_u3_u4_n161, u2_u3_u4_n162, u2_u3_u4_n163, u2_u3_u4_n164, u2_u3_u4_n165, 
       u2_u3_u4_n166, u2_u3_u4_n167, u2_u3_u4_n168, u2_u3_u4_n169, u2_u3_u4_n170, u2_u3_u4_n171, u2_u3_u4_n172, u2_u3_u4_n173, u2_u3_u4_n174, 
       u2_u3_u4_n175, u2_u3_u4_n176, u2_u3_u4_n177, u2_u3_u4_n178, u2_u3_u4_n179, u2_u3_u4_n180, u2_u3_u4_n181, u2_u3_u4_n182, u2_u3_u4_n183, 
       u2_u3_u4_n184, u2_u3_u4_n185, u2_u3_u4_n186, u2_u3_u4_n94, u2_u3_u4_n95, u2_u3_u4_n96, u2_u3_u4_n97, u2_u3_u4_n98, u2_u3_u4_n99, 
       u2_u3_u5_n100, u2_u3_u5_n101, u2_u3_u5_n102, u2_u3_u5_n103, u2_u3_u5_n104, u2_u3_u5_n105, u2_u3_u5_n106, u2_u3_u5_n107, u2_u3_u5_n108, 
       u2_u3_u5_n109, u2_u3_u5_n110, u2_u3_u5_n111, u2_u3_u5_n112, u2_u3_u5_n113, u2_u3_u5_n114, u2_u3_u5_n115, u2_u3_u5_n116, u2_u3_u5_n117, 
       u2_u3_u5_n118, u2_u3_u5_n119, u2_u3_u5_n120, u2_u3_u5_n121, u2_u3_u5_n122, u2_u3_u5_n123, u2_u3_u5_n124, u2_u3_u5_n125, u2_u3_u5_n126, 
       u2_u3_u5_n127, u2_u3_u5_n128, u2_u3_u5_n129, u2_u3_u5_n130, u2_u3_u5_n131, u2_u3_u5_n132, u2_u3_u5_n133, u2_u3_u5_n134, u2_u3_u5_n135, 
       u2_u3_u5_n136, u2_u3_u5_n137, u2_u3_u5_n138, u2_u3_u5_n139, u2_u3_u5_n140, u2_u3_u5_n141, u2_u3_u5_n142, u2_u3_u5_n143, u2_u3_u5_n144, 
       u2_u3_u5_n145, u2_u3_u5_n146, u2_u3_u5_n147, u2_u3_u5_n148, u2_u3_u5_n149, u2_u3_u5_n150, u2_u3_u5_n151, u2_u3_u5_n152, u2_u3_u5_n153, 
       u2_u3_u5_n154, u2_u3_u5_n155, u2_u3_u5_n156, u2_u3_u5_n157, u2_u3_u5_n158, u2_u3_u5_n159, u2_u3_u5_n160, u2_u3_u5_n161, u2_u3_u5_n162, 
       u2_u3_u5_n163, u2_u3_u5_n164, u2_u3_u5_n165, u2_u3_u5_n166, u2_u3_u5_n167, u2_u3_u5_n168, u2_u3_u5_n169, u2_u3_u5_n170, u2_u3_u5_n171, 
       u2_u3_u5_n172, u2_u3_u5_n173, u2_u3_u5_n174, u2_u3_u5_n175, u2_u3_u5_n176, u2_u3_u5_n177, u2_u3_u5_n178, u2_u3_u5_n179, u2_u3_u5_n180, 
       u2_u3_u5_n181, u2_u3_u5_n182, u2_u3_u5_n183, u2_u3_u5_n184, u2_u3_u5_n185, u2_u3_u5_n186, u2_u3_u5_n187, u2_u3_u5_n188, u2_u3_u5_n189, 
       u2_u3_u5_n190, u2_u3_u5_n191, u2_u3_u5_n192, u2_u3_u5_n193, u2_u3_u5_n194, u2_u3_u5_n195, u2_u3_u5_n196, u2_u3_u5_n99, u2_u3_u6_n100, 
       u2_u3_u6_n101, u2_u3_u6_n102, u2_u3_u6_n103, u2_u3_u6_n104, u2_u3_u6_n105, u2_u3_u6_n106, u2_u3_u6_n107, u2_u3_u6_n108, u2_u3_u6_n109, 
       u2_u3_u6_n110, u2_u3_u6_n111, u2_u3_u6_n112, u2_u3_u6_n113, u2_u3_u6_n114, u2_u3_u6_n115, u2_u3_u6_n116, u2_u3_u6_n117, u2_u3_u6_n118, 
       u2_u3_u6_n119, u2_u3_u6_n120, u2_u3_u6_n121, u2_u3_u6_n122, u2_u3_u6_n123, u2_u3_u6_n124, u2_u3_u6_n125, u2_u3_u6_n126, u2_u3_u6_n127, 
       u2_u3_u6_n128, u2_u3_u6_n129, u2_u3_u6_n130, u2_u3_u6_n131, u2_u3_u6_n132, u2_u3_u6_n133, u2_u3_u6_n134, u2_u3_u6_n135, u2_u3_u6_n136, 
       u2_u3_u6_n137, u2_u3_u6_n138, u2_u3_u6_n139, u2_u3_u6_n140, u2_u3_u6_n141, u2_u3_u6_n142, u2_u3_u6_n143, u2_u3_u6_n144, u2_u3_u6_n145, 
       u2_u3_u6_n146, u2_u3_u6_n147, u2_u3_u6_n148, u2_u3_u6_n149, u2_u3_u6_n150, u2_u3_u6_n151, u2_u3_u6_n152, u2_u3_u6_n153, u2_u3_u6_n154, 
       u2_u3_u6_n155, u2_u3_u6_n156, u2_u3_u6_n157, u2_u3_u6_n158, u2_u3_u6_n159, u2_u3_u6_n160, u2_u3_u6_n161, u2_u3_u6_n162, u2_u3_u6_n163, 
       u2_u3_u6_n164, u2_u3_u6_n165, u2_u3_u6_n166, u2_u3_u6_n167, u2_u3_u6_n168, u2_u3_u6_n169, u2_u3_u6_n170, u2_u3_u6_n171, u2_u3_u6_n172, 
       u2_u3_u6_n173, u2_u3_u6_n174, u2_u3_u6_n88, u2_u3_u6_n89, u2_u3_u6_n90, u2_u3_u6_n91, u2_u3_u6_n92, u2_u3_u6_n93, u2_u3_u6_n94, 
       u2_u3_u6_n95, u2_u3_u6_n96, u2_u3_u6_n97, u2_u3_u6_n98, u2_u3_u6_n99, u2_u5_X_1, u2_u5_X_10, u2_u5_X_11, u2_u5_X_12, 
       u2_u5_X_2, u2_u5_X_3, u2_u5_X_4, u2_u5_X_43, u2_u5_X_44, u2_u5_X_45, u2_u5_X_46, u2_u5_X_47, u2_u5_X_48, 
       u2_u5_X_5, u2_u5_X_6, u2_u5_X_7, u2_u5_X_8, u2_u5_X_9, u2_u5_u0_n100, u2_u5_u0_n101, u2_u5_u0_n102, u2_u5_u0_n103, 
       u2_u5_u0_n104, u2_u5_u0_n105, u2_u5_u0_n106, u2_u5_u0_n107, u2_u5_u0_n108, u2_u5_u0_n109, u2_u5_u0_n110, u2_u5_u0_n111, u2_u5_u0_n112, 
       u2_u5_u0_n113, u2_u5_u0_n114, u2_u5_u0_n115, u2_u5_u0_n116, u2_u5_u0_n117, u2_u5_u0_n118, u2_u5_u0_n119, u2_u5_u0_n120, u2_u5_u0_n121, 
       u2_u5_u0_n122, u2_u5_u0_n123, u2_u5_u0_n124, u2_u5_u0_n125, u2_u5_u0_n126, u2_u5_u0_n127, u2_u5_u0_n128, u2_u5_u0_n129, u2_u5_u0_n130, 
       u2_u5_u0_n131, u2_u5_u0_n132, u2_u5_u0_n133, u2_u5_u0_n134, u2_u5_u0_n135, u2_u5_u0_n136, u2_u5_u0_n137, u2_u5_u0_n138, u2_u5_u0_n139, 
       u2_u5_u0_n140, u2_u5_u0_n141, u2_u5_u0_n142, u2_u5_u0_n143, u2_u5_u0_n144, u2_u5_u0_n145, u2_u5_u0_n146, u2_u5_u0_n147, u2_u5_u0_n148, 
       u2_u5_u0_n149, u2_u5_u0_n150, u2_u5_u0_n151, u2_u5_u0_n152, u2_u5_u0_n153, u2_u5_u0_n154, u2_u5_u0_n155, u2_u5_u0_n156, u2_u5_u0_n157, 
       u2_u5_u0_n158, u2_u5_u0_n159, u2_u5_u0_n160, u2_u5_u0_n161, u2_u5_u0_n162, u2_u5_u0_n163, u2_u5_u0_n164, u2_u5_u0_n165, u2_u5_u0_n166, 
       u2_u5_u0_n167, u2_u5_u0_n168, u2_u5_u0_n169, u2_u5_u0_n170, u2_u5_u0_n171, u2_u5_u0_n172, u2_u5_u0_n173, u2_u5_u0_n174, u2_u5_u0_n88, 
       u2_u5_u0_n89, u2_u5_u0_n90, u2_u5_u0_n91, u2_u5_u0_n92, u2_u5_u0_n93, u2_u5_u0_n94, u2_u5_u0_n95, u2_u5_u0_n96, u2_u5_u0_n97, 
       u2_u5_u0_n98, u2_u5_u0_n99, u2_u5_u1_n100, u2_u5_u1_n101, u2_u5_u1_n102, u2_u5_u1_n103, u2_u5_u1_n104, u2_u5_u1_n105, u2_u5_u1_n106, 
       u2_u5_u1_n107, u2_u5_u1_n108, u2_u5_u1_n109, u2_u5_u1_n110, u2_u5_u1_n111, u2_u5_u1_n112, u2_u5_u1_n113, u2_u5_u1_n114, u2_u5_u1_n115, 
       u2_u5_u1_n116, u2_u5_u1_n117, u2_u5_u1_n118, u2_u5_u1_n119, u2_u5_u1_n120, u2_u5_u1_n121, u2_u5_u1_n122, u2_u5_u1_n123, u2_u5_u1_n124, 
       u2_u5_u1_n125, u2_u5_u1_n126, u2_u5_u1_n127, u2_u5_u1_n128, u2_u5_u1_n129, u2_u5_u1_n130, u2_u5_u1_n131, u2_u5_u1_n132, u2_u5_u1_n133, 
       u2_u5_u1_n134, u2_u5_u1_n135, u2_u5_u1_n136, u2_u5_u1_n137, u2_u5_u1_n138, u2_u5_u1_n139, u2_u5_u1_n140, u2_u5_u1_n141, u2_u5_u1_n142, 
       u2_u5_u1_n143, u2_u5_u1_n144, u2_u5_u1_n145, u2_u5_u1_n146, u2_u5_u1_n147, u2_u5_u1_n148, u2_u5_u1_n149, u2_u5_u1_n150, u2_u5_u1_n151, 
       u2_u5_u1_n152, u2_u5_u1_n153, u2_u5_u1_n154, u2_u5_u1_n155, u2_u5_u1_n156, u2_u5_u1_n157, u2_u5_u1_n158, u2_u5_u1_n159, u2_u5_u1_n160, 
       u2_u5_u1_n161, u2_u5_u1_n162, u2_u5_u1_n163, u2_u5_u1_n164, u2_u5_u1_n165, u2_u5_u1_n166, u2_u5_u1_n167, u2_u5_u1_n168, u2_u5_u1_n169, 
       u2_u5_u1_n170, u2_u5_u1_n171, u2_u5_u1_n172, u2_u5_u1_n173, u2_u5_u1_n174, u2_u5_u1_n175, u2_u5_u1_n176, u2_u5_u1_n177, u2_u5_u1_n178, 
       u2_u5_u1_n179, u2_u5_u1_n180, u2_u5_u1_n181, u2_u5_u1_n182, u2_u5_u1_n183, u2_u5_u1_n184, u2_u5_u1_n185, u2_u5_u1_n186, u2_u5_u1_n187, 
       u2_u5_u1_n188, u2_u5_u1_n95, u2_u5_u1_n96, u2_u5_u1_n97, u2_u5_u1_n98, u2_u5_u1_n99, u2_u5_u7_n100, u2_u5_u7_n101, u2_u5_u7_n102, 
       u2_u5_u7_n103, u2_u5_u7_n104, u2_u5_u7_n105, u2_u5_u7_n106, u2_u5_u7_n107, u2_u5_u7_n108, u2_u5_u7_n109, u2_u5_u7_n110, u2_u5_u7_n111, 
       u2_u5_u7_n112, u2_u5_u7_n113, u2_u5_u7_n114, u2_u5_u7_n115, u2_u5_u7_n116, u2_u5_u7_n117, u2_u5_u7_n118, u2_u5_u7_n119, u2_u5_u7_n120, 
       u2_u5_u7_n121, u2_u5_u7_n122, u2_u5_u7_n123, u2_u5_u7_n124, u2_u5_u7_n125, u2_u5_u7_n126, u2_u5_u7_n127, u2_u5_u7_n128, u2_u5_u7_n129, 
       u2_u5_u7_n130, u2_u5_u7_n131, u2_u5_u7_n132, u2_u5_u7_n133, u2_u5_u7_n134, u2_u5_u7_n135, u2_u5_u7_n136, u2_u5_u7_n137, u2_u5_u7_n138, 
       u2_u5_u7_n139, u2_u5_u7_n140, u2_u5_u7_n141, u2_u5_u7_n142, u2_u5_u7_n143, u2_u5_u7_n144, u2_u5_u7_n145, u2_u5_u7_n146, u2_u5_u7_n147, 
       u2_u5_u7_n148, u2_u5_u7_n149, u2_u5_u7_n150, u2_u5_u7_n151, u2_u5_u7_n152, u2_u5_u7_n153, u2_u5_u7_n154, u2_u5_u7_n155, u2_u5_u7_n156, 
       u2_u5_u7_n157, u2_u5_u7_n158, u2_u5_u7_n159, u2_u5_u7_n160, u2_u5_u7_n161, u2_u5_u7_n162, u2_u5_u7_n163, u2_u5_u7_n164, u2_u5_u7_n165, 
       u2_u5_u7_n166, u2_u5_u7_n167, u2_u5_u7_n168, u2_u5_u7_n169, u2_u5_u7_n170, u2_u5_u7_n171, u2_u5_u7_n172, u2_u5_u7_n173, u2_u5_u7_n174, 
       u2_u5_u7_n175, u2_u5_u7_n176, u2_u5_u7_n177, u2_u5_u7_n178, u2_u5_u7_n179, u2_u5_u7_n180, u2_u5_u7_n91, u2_u5_u7_n92, u2_u5_u7_n93, 
       u2_u5_u7_n94, u2_u5_u7_n95, u2_u5_u7_n96, u2_u5_u7_n97, u2_u5_u7_n98, u2_u5_u7_n99, u2_uk_n1008, u2_uk_n1009, u2_uk_n1010, 
       u2_uk_n1014, u2_uk_n1015, u2_uk_n1016, u2_uk_n1017, u2_uk_n1029, u2_uk_n1030, u2_uk_n1032, u2_uk_n1033, u2_uk_n1058, 
       u2_uk_n1066, u2_uk_n1071, u2_uk_n1072, u2_uk_n312, u2_uk_n335, u2_uk_n338, u2_uk_n342, u2_uk_n349, u2_uk_n353, 
       u2_uk_n391, u2_uk_n407, u2_uk_n601, u2_uk_n634, u2_uk_n662, u2_uk_n671,  u2_uk_n688;
  XOR2_X1 u0_U13 (.Z( u0_N9 ) , .B( u0_desIn_r_12 ) , .A( u0_out0_10 ) );
  XOR2_X1 u0_U130 (.B( u0_L11_32 ) , .Z( u0_N415 ) , .A( u0_out12_32 ) );
  XOR2_X1 u0_U133 (.B( u0_L11_29 ) , .Z( u0_N412 ) , .A( u0_out12_29 ) );
  XOR2_X1 u0_U138 (.B( u0_L11_25 ) , .Z( u0_N408 ) , .A( u0_out12_25 ) );
  XOR2_X1 u0_U141 (.B( u0_L11_22 ) , .Z( u0_N405 ) , .A( u0_out12_22 ) );
  XOR2_X1 u0_U144 (.B( u0_L11_19 ) , .Z( u0_N402 ) , .A( u0_out12_19 ) );
  XOR2_X1 u0_U151 (.B( u0_L11_14 ) , .Z( u0_N397 ) , .A( u0_out12_14 ) );
  XOR2_X1 u0_U153 (.B( u0_L11_12 ) , .Z( u0_N395 ) , .A( u0_out12_12 ) );
  XOR2_X1 u0_U154 (.B( u0_L11_11 ) , .Z( u0_N394 ) , .A( u0_out12_11 ) );
  XOR2_X1 u0_U157 (.B( u0_L11_8 ) , .Z( u0_N391 ) , .A( u0_out12_8 ) );
  XOR2_X1 u0_U158 (.B( u0_L11_7 ) , .Z( u0_N390 ) , .A( u0_out12_7 ) );
  XOR2_X1 u0_U162 (.B( u0_L11_4 ) , .Z( u0_N387 ) , .A( u0_out12_4 ) );
  XOR2_X1 u0_U163 (.B( u0_L11_3 ) , .Z( u0_N386 ) , .A( u0_out12_3 ) );
  XOR2_X1 u0_U24 (.Z( u0_N8 ) , .B( u0_desIn_r_4 ) , .A( u0_out0_9 ) );
  XOR2_X1 u0_U258 (.Z( u0_N30 ) , .B( u0_desIn_r_48 ) , .A( u0_out0_31 ) );
  XOR2_X1 u0_U278 (.B( u0_L7_27 ) , .Z( u0_N282 ) , .A( u0_out8_27 ) );
  XOR2_X1 u0_U279 (.B( u0_L7_26 ) , .Z( u0_N281 ) , .A( u0_out8_26 ) );
  XOR2_X1 u0_U280 (.B( u0_L7_25 ) , .Z( u0_N280 ) , .A( u0_out8_25 ) );
  XOR2_X1 u0_U285 (.B( u0_L7_21 ) , .Z( u0_N276 ) , .A( u0_out8_21 ) );
  XOR2_X1 u0_U286 (.B( u0_L7_20 ) , .Z( u0_N275 ) , .A( u0_out8_20 ) );
  XOR2_X1 u0_U291 (.B( u0_L7_15 ) , .Z( u0_N270 ) , .A( u0_out8_15 ) );
  XOR2_X1 u0_U292 (.Z( u0_N27 ) , .B( u0_desIn_r_24 ) , .A( u0_out0_28 ) );
  XOR2_X1 u0_U293 (.B( u0_L7_14 ) , .Z( u0_N269 ) , .A( u0_out8_14 ) );
  XOR2_X1 u0_U297 (.B( u0_L7_10 ) , .Z( u0_N265 ) , .A( u0_out8_10 ) );
  XOR2_X1 u0_U299 (.B( u0_L7_8 ) , .Z( u0_N263 ) , .A( u0_out8_8 ) );
  XOR2_X1 u0_U302 (.B( u0_L7_5 ) , .Z( u0_N260 ) , .A( u0_out8_5 ) );
  XOR2_X1 u0_U305 (.B( u0_L7_3 ) , .Z( u0_N258 ) , .A( u0_out8_3 ) );
  XOR2_X1 u0_U307 (.B( u0_L7_1 ) , .Z( u0_N256 ) , .A( u0_out8_1 ) );
  XOR2_X1 u0_U314 (.Z( u0_N25 ) , .B( u0_desIn_r_8 ) , .A( u0_out0_26 ) );
  XOR2_X1 u0_U343 (.B( u0_L5_32 ) , .Z( u0_N223 ) , .A( u0_out6_32 ) );
  XOR2_X1 u0_U346 (.B( u0_L5_29 ) , .Z( u0_N220 ) , .A( u0_out6_29 ) );
  XOR2_X1 u0_U347 (.Z( u0_N22 ) , .B( u0_desIn_r_50 ) , .A( u0_out0_23 ) );
  XOR2_X1 u0_U351 (.B( u0_L5_25 ) , .Z( u0_N216 ) , .A( u0_out6_25 ) );
  XOR2_X1 u0_U354 (.B( u0_L5_22 ) , .Z( u0_N213 ) , .A( u0_out6_22 ) );
  XOR2_X1 u0_U357 (.B( u0_L5_19 ) , .Z( u0_N210 ) , .A( u0_out6_19 ) );
  XOR2_X1 u0_U363 (.B( u0_L5_14 ) , .Z( u0_N205 ) , .A( u0_out6_14 ) );
  XOR2_X1 u0_U365 (.B( u0_L5_12 ) , .Z( u0_N203 ) , .A( u0_out6_12 ) );
  XOR2_X1 u0_U366 (.B( u0_L5_11 ) , .Z( u0_N202 ) , .A( u0_out6_11 ) );
  XOR2_X1 u0_U371 (.B( u0_L5_8 ) , .Z( u0_N199 ) , .A( u0_out6_8 ) );
  XOR2_X1 u0_U372 (.B( u0_L5_7 ) , .Z( u0_N198 ) , .A( u0_out6_7 ) );
  XOR2_X1 u0_U375 (.B( u0_L5_4 ) , .Z( u0_N195 ) , .A( u0_out6_4 ) );
  XOR2_X1 u0_U376 (.B( u0_L5_3 ) , .Z( u0_N194 ) , .A( u0_out6_3 ) );
  XOR2_X1 u0_U381 (.Z( u0_N19 ) , .B( u0_desIn_r_26 ) , .A( u0_out0_20 ) );
  XOR2_X1 u0_U403 (.Z( u0_N17 ) , .B( u0_desIn_r_10 ) , .A( u0_out0_18 ) );
  XOR2_X1 u0_U414 (.Z( u0_N16 ) , .B( u0_desIn_r_2 ) , .A( u0_out0_17 ) );
  XOR2_X1 u0_U417 (.B( u0_L3_30 ) , .Z( u0_N157 ) , .A( u0_out4_30 ) );
  XOR2_X1 u0_U419 (.B( u0_L3_28 ) , .Z( u0_N155 ) , .A( u0_out4_28 ) );
  XOR2_X1 u0_U421 (.B( u0_L3_26 ) , .Z( u0_N153 ) , .A( u0_out4_26 ) );
  XOR2_X1 u0_U423 (.B( u0_L3_24 ) , .Z( u0_N151 ) , .A( u0_out4_24 ) );
  XOR2_X1 u0_U428 (.B( u0_L3_20 ) , .Z( u0_N147 ) , .A( u0_out4_20 ) );
  XOR2_X1 u0_U430 (.B( u0_L3_18 ) , .Z( u0_N145 ) , .A( u0_out4_18 ) );
  XOR2_X1 u0_U432 (.B( u0_L3_16 ) , .Z( u0_N143 ) , .A( u0_out4_16 ) );
  XOR2_X1 u0_U435 (.B( u0_L3_13 ) , .Z( u0_N140 ) , .A( u0_out4_13 ) );
  XOR2_X1 u0_U439 (.B( u0_L3_10 ) , .Z( u0_N137 ) , .A( u0_out4_10 ) );
  XOR2_X1 u0_U443 (.B( u0_L3_6 ) , .Z( u0_N133 ) , .A( u0_out4_6 ) );
  XOR2_X1 u0_U448 (.B( u0_L3_2 ) , .Z( u0_N129 ) , .A( u0_out4_2 ) );
  XOR2_X1 u0_U449 (.B( u0_L3_1 ) , .Z( u0_N128 ) , .A( u0_out4_1 ) );
  XOR2_X1 u0_U458 (.Z( u0_N12 ) , .B( u0_desIn_r_36 ) , .A( u0_out0_13 ) );
  XOR2_X1 u0_U481 (.Z( u0_N1 ) , .B( u0_desIn_r_14 ) , .A( u0_out0_2 ) );
  XOR2_X1 u0_U482 (.Z( u0_N0 ) , .B( u0_desIn_r_6 ) , .A( u0_out0_1 ) );
  XOR2_X1 u0_U484 (.Z( u0_FP_8 ) , .B( u0_L14_8 ) , .A( u0_out15_8 ) );
  XOR2_X1 u0_U485 (.Z( u0_FP_7 ) , .B( u0_L14_7 ) , .A( u0_out15_7 ) );
  XOR2_X1 u0_U488 (.Z( u0_FP_4 ) , .B( u0_L14_4 ) , .A( u0_out15_4 ) );
  XOR2_X1 u0_U489 (.Z( u0_FP_3 ) , .B( u0_L14_3 ) , .A( u0_out15_3 ) );
  XOR2_X1 u0_U490 (.Z( u0_FP_32 ) , .B( u0_L14_32 ) , .A( u0_out15_32 ) );
  XOR2_X1 u0_U494 (.Z( u0_FP_29 ) , .B( u0_L14_29 ) , .A( u0_out15_29 ) );
  XOR2_X1 u0_U498 (.Z( u0_FP_25 ) , .B( u0_L14_25 ) , .A( u0_out15_25 ) );
  XOR2_X1 u0_U501 (.Z( u0_FP_22 ) , .B( u0_L14_22 ) , .A( u0_out15_22 ) );
  XOR2_X1 u0_U505 (.Z( u0_FP_19 ) , .B( u0_L14_19 ) , .A( u0_out15_19 ) );
  XOR2_X1 u0_U510 (.Z( u0_FP_14 ) , .B( u0_L14_14 ) , .A( u0_out15_14 ) );
  XOR2_X1 u0_U512 (.Z( u0_FP_12 ) , .B( u0_L14_12 ) , .A( u0_out15_12 ) );
  XOR2_X1 u0_U513 (.Z( u0_FP_11 ) , .B( u0_L14_11 ) , .A( u0_out15_11 ) );
  XOR2_X1 u0_u0_U1 (.B( u0_K1_9 ) , .A( u0_desIn_r_47 ) , .Z( u0_u0_X_9 ) );
  XOR2_X1 u0_u0_U16 (.B( u0_K1_3 ) , .A( u0_desIn_r_15 ) , .Z( u0_u0_X_3 ) );
  XOR2_X1 u0_u0_U2 (.B( u0_K1_8 ) , .A( u0_desIn_r_39 ) , .Z( u0_u0_X_8 ) );
  XOR2_X1 u0_u0_U27 (.B( u0_K1_2 ) , .A( u0_desIn_r_7 ) , .Z( u0_u0_X_2 ) );
  XOR2_X1 u0_u0_U3 (.B( u0_K1_7 ) , .A( u0_desIn_r_31 ) , .Z( u0_u0_X_7 ) );
  XOR2_X1 u0_u0_U33 (.B( u0_K1_24 ) , .A( u0_desIn_r_3 ) , .Z( u0_u0_X_24 ) );
  XOR2_X1 u0_u0_U34 (.B( u0_K1_23 ) , .A( u0_desIn_r_61 ) , .Z( u0_u0_X_23 ) );
  XOR2_X1 u0_u0_U35 (.B( u0_K1_22 ) , .A( u0_desIn_r_53 ) , .Z( u0_u0_X_22 ) );
  XOR2_X1 u0_u0_U36 (.B( u0_K1_21 ) , .A( u0_desIn_r_45 ) , .Z( u0_u0_X_21 ) );
  XOR2_X1 u0_u0_U37 (.B( u0_K1_20 ) , .A( u0_desIn_r_37 ) , .Z( u0_u0_X_20 ) );
  XOR2_X1 u0_u0_U38 (.B( u0_K1_1 ) , .A( u0_desIn_r_57 ) , .Z( u0_u0_X_1 ) );
  XOR2_X1 u0_u0_U39 (.B( u0_K1_19 ) , .A( u0_desIn_r_29 ) , .Z( u0_u0_X_19 ) );
  XOR2_X1 u0_u0_U4 (.B( u0_K1_6 ) , .A( u0_desIn_r_39 ) , .Z( u0_u0_X_6 ) );
  XOR2_X1 u0_u0_U46 (.B( u0_K1_12 ) , .A( u0_desIn_r_5 ) , .Z( u0_u0_X_12 ) );
  XOR2_X1 u0_u0_U47 (.B( u0_K1_11 ) , .A( u0_desIn_r_63 ) , .Z( u0_u0_X_11 ) );
  XOR2_X1 u0_u0_U48 (.B( u0_K1_10 ) , .A( u0_desIn_r_55 ) , .Z( u0_u0_X_10 ) );
  XOR2_X1 u0_u0_U5 (.B( u0_K1_5 ) , .A( u0_desIn_r_31 ) , .Z( u0_u0_X_5 ) );
  XOR2_X1 u0_u0_U6 (.B( u0_K1_4 ) , .A( u0_desIn_r_23 ) , .Z( u0_u0_X_4 ) );
  AND3_X1 u0_u0_u0_U10 (.A1( u0_u0_u0_n27 ) , .A3( u0_u0_u0_n45 ) , .ZN( u0_u0_u0_n48 ) , .A2( u0_u0_u0_n63 ) );
  NAND2_X1 u0_u0_u0_U11 (.A2( u0_u0_u0_n26 ) , .A1( u0_u0_u0_n36 ) , .ZN( u0_u0_u0_n62 ) );
  AND2_X1 u0_u0_u0_U12 (.A2( u0_u0_u0_n35 ) , .A1( u0_u0_u0_n45 ) , .ZN( u0_u0_u0_n68 ) );
  AND2_X1 u0_u0_u0_U13 (.ZN( u0_u0_u0_n24 ) , .A1( u0_u0_u0_n45 ) , .A2( u0_u0_u0_n46 ) );
  AND2_X1 u0_u0_u0_U14 (.ZN( u0_u0_u0_n30 ) , .A2( u0_u0_u0_n50 ) , .A1( u0_u0_u0_n67 ) );
  INV_X1 u0_u0_u0_U15 (.ZN( u0_u0_u0_n2 ) , .A( u0_u0_u0_n32 ) );
  NOR2_X1 u0_u0_u0_U16 (.A1( u0_u0_u0_n15 ) , .ZN( u0_u0_u0_n28 ) , .A2( u0_u0_u0_n39 ) );
  AOI21_X1 u0_u0_u0_U17 (.A( u0_u0_u0_n10 ) , .ZN( u0_u0_u0_n43 ) , .B1( u0_u0_u0_n72 ) , .B2( u0_u0_u0_n82 ) );
  INV_X1 u0_u0_u0_U18 (.ZN( u0_u0_u0_n10 ) , .A( u0_u0_u0_n33 ) );
  OAI22_X1 u0_u0_u0_U19 (.B2( u0_u0_u0_n28 ) , .A2( u0_u0_u0_n29 ) , .A1( u0_u0_u0_n37 ) , .ZN( u0_u0_u0_n49 ) , .B1( u0_u0_u0_n50 ) );
  OAI22_X1 u0_u0_u0_U20 (.B2( u0_u0_u0_n28 ) , .A1( u0_u0_u0_n31 ) , .B1( u0_u0_u0_n44 ) , .ZN( u0_u0_u0_n84 ) , .A2( u0_u0_u0_n85 ) );
  AND3_X1 u0_u0_u0_U21 (.A1( u0_u0_u0_n27 ) , .A2( u0_u0_u0_n50 ) , .A3( u0_u0_u0_n54 ) , .ZN( u0_u0_u0_n85 ) );
  NAND2_X1 u0_u0_u0_U22 (.ZN( u0_u0_u0_n50 ) , .A2( u0_u0_u0_n72 ) , .A1( u0_u0_u0_n75 ) );
  INV_X1 u0_u0_u0_U23 (.ZN( u0_u0_u0_n14 ) , .A( u0_u0_u0_n39 ) );
  AOI22_X1 u0_u0_u0_U24 (.A1( u0_u0_u0_n15 ) , .B1( u0_u0_u0_n57 ) , .ZN( u0_u0_u0_n64 ) , .A2( u0_u0_u0_n65 ) , .B2( u0_u0_u0_n66 ) );
  NAND2_X1 u0_u0_u0_U25 (.ZN( u0_u0_u0_n46 ) , .A1( u0_u0_u0_n75 ) , .A2( u0_u0_u0_n80 ) );
  INV_X1 u0_u0_u0_U26 (.ZN( u0_u0_u0_n17 ) , .A( u0_u0_u0_n57 ) );
  AOI21_X1 u0_u0_u0_U27 (.A( u0_u0_u0_n31 ) , .B2( u0_u0_u0_n34 ) , .B1( u0_u0_u0_n68 ) , .ZN( u0_u0_u0_n71 ) );
  AOI21_X1 u0_u0_u0_U28 (.A( u0_u0_u0_n37 ) , .B2( u0_u0_u0_n46 ) , .B1( u0_u0_u0_n48 ) , .ZN( u0_u0_u0_n79 ) );
  AOI21_X1 u0_u0_u0_U29 (.A( u0_u0_u0_n31 ) , .B2( u0_u0_u0_n33 ) , .ZN( u0_u0_u0_n59 ) , .B1( u0_u0_u0_n9 ) );
  INV_X1 u0_u0_u0_U3 (.A( u0_u0_u0_n62 ) , .ZN( u0_u0_u0_n9 ) );
  NOR2_X1 u0_u0_u0_U30 (.ZN( u0_u0_u0_n32 ) , .A1( u0_u0_u0_n55 ) , .A2( u0_u0_u0_n8 ) );
  OAI221_X1 u0_u0_u0_U31 (.C2( u0_u0_u0_n28 ) , .A( u0_u0_u0_n3 ) , .B2( u0_u0_u0_n34 ) , .B1( u0_u0_u0_n37 ) , .ZN( u0_u0_u0_n55 ) , .C1( u0_u0_u0_n63 ) );
  AOI211_X1 u0_u0_u0_U32 (.ZN( u0_u0_u0_n56 ) , .C1( u0_u0_u0_n57 ) , .C2( u0_u0_u0_n58 ) , .A( u0_u0_u0_n59 ) , .B( u0_u0_u0_n60 ) );
  NAND2_X1 u0_u0_u0_U33 (.ZN( u0_u0_u0_n47 ) , .A1( u0_u0_u0_n73 ) , .A2( u0_u0_u0_n80 ) );
  NAND2_X1 u0_u0_u0_U34 (.ZN( u0_u0_u0_n36 ) , .A1( u0_u0_u0_n74 ) , .A2( u0_u0_u0_n75 ) );
  NAND2_X1 u0_u0_u0_U35 (.ZN( u0_u0_u0_n27 ) , .A2( u0_u0_u0_n80 ) , .A1( u0_u0_u0_n82 ) );
  NAND2_X1 u0_u0_u0_U36 (.ZN( u0_u0_u0_n44 ) , .A2( u0_u0_u0_n75 ) , .A1( u0_u0_u0_n83 ) );
  NAND2_X1 u0_u0_u0_U37 (.ZN( u0_u0_u0_n25 ) , .A2( u0_u0_u0_n73 ) , .A1( u0_u0_u0_n74 ) );
  INV_X1 u0_u0_u0_U38 (.ZN( u0_u0_u0_n15 ) , .A( u0_u0_u0_n37 ) );
  NAND2_X1 u0_u0_u0_U39 (.ZN( u0_u0_u0_n26 ) , .A1( u0_u0_u0_n72 ) , .A2( u0_u0_u0_n73 ) );
  AOI21_X1 u0_u0_u0_U4 (.A( u0_u0_u0_n14 ) , .B2( u0_u0_u0_n46 ) , .ZN( u0_u0_u0_n60 ) , .B1( u0_u0_u0_n61 ) );
  NAND2_X1 u0_u0_u0_U40 (.ZN( u0_u0_u0_n61 ) , .A2( u0_u0_u0_n73 ) , .A1( u0_u0_u0_n83 ) );
  INV_X1 u0_u0_u0_U41 (.ZN( u0_u0_u0_n3 ) , .A( u0_u0_u0_n87 ) );
  OAI222_X1 u0_u0_u0_U42 (.C2( u0_u0_u0_n14 ) , .A2( u0_u0_u0_n17 ) , .B1( u0_u0_u0_n31 ) , .B2( u0_u0_u0_n47 ) , .A1( u0_u0_u0_n50 ) , .C1( u0_u0_u0_n67 ) , .ZN( u0_u0_u0_n87 ) );
  NAND2_X1 u0_u0_u0_U43 (.ZN( u0_u0_u0_n54 ) , .A2( u0_u0_u0_n74 ) , .A1( u0_u0_u0_n82 ) );
  NAND2_X1 u0_u0_u0_U44 (.ZN( u0_u0_u0_n63 ) , .A1( u0_u0_u0_n82 ) , .A2( u0_u0_u0_n83 ) );
  OR3_X1 u0_u0_u0_U45 (.ZN( u0_u0_u0_n20 ) , .A1( u0_u0_u0_n21 ) , .A2( u0_u0_u0_n22 ) , .A3( u0_u0_u0_n23 ) );
  AOI21_X1 u0_u0_u0_U46 (.A( u0_u0_u0_n17 ) , .ZN( u0_u0_u0_n23 ) , .B1( u0_u0_u0_n24 ) , .B2( u0_u0_u0_n25 ) );
  AOI21_X1 u0_u0_u0_U47 (.ZN( u0_u0_u0_n21 ) , .B1( u0_u0_u0_n29 ) , .B2( u0_u0_u0_n30 ) , .A( u0_u0_u0_n31 ) );
  AOI21_X1 u0_u0_u0_U48 (.ZN( u0_u0_u0_n22 ) , .B1( u0_u0_u0_n26 ) , .B2( u0_u0_u0_n27 ) , .A( u0_u0_u0_n28 ) );
  INV_X1 u0_u0_u0_U49 (.ZN( u0_u0_u0_n4 ) , .A( u0_u0_u0_n76 ) );
  AOI21_X1 u0_u0_u0_U5 (.A( u0_u0_u0_n17 ) , .B1( u0_u0_u0_n24 ) , .ZN( u0_u0_u0_n41 ) , .B2( u0_u0_u0_n44 ) );
  OAI211_X1 u0_u0_u0_U50 (.C1( u0_u0_u0_n14 ) , .C2( u0_u0_u0_n35 ) , .A( u0_u0_u0_n6 ) , .ZN( u0_u0_u0_n76 ) , .B( u0_u0_u0_n77 ) );
  INV_X1 u0_u0_u0_U51 (.ZN( u0_u0_u0_n6 ) , .A( u0_u0_u0_n84 ) );
  AOI211_X1 u0_u0_u0_U52 (.A( u0_u0_u0_n52 ) , .C1( u0_u0_u0_n57 ) , .ZN( u0_u0_u0_n77 ) , .C2( u0_u0_u0_n78 ) , .B( u0_u0_u0_n79 ) );
  NOR2_X1 u0_u0_u0_U53 (.A2( u0_u0_X_4 ) , .A1( u0_u0_X_5 ) , .ZN( u0_u0_u0_n57 ) );
  NOR2_X1 u0_u0_u0_U54 (.A2( u0_u0_X_2 ) , .A1( u0_u0_u0_n11 ) , .ZN( u0_u0_u0_n72 ) );
  NOR2_X1 u0_u0_u0_U55 (.A2( u0_u0_X_1 ) , .A1( u0_u0_X_2 ) , .ZN( u0_u0_u0_n83 ) );
  NOR2_X1 u0_u0_u0_U56 (.A2( u0_u0_X_1 ) , .A1( u0_u0_u0_n12 ) , .ZN( u0_u0_u0_n74 ) );
  NAND2_X1 u0_u0_u0_U57 (.A2( u0_u0_X_4 ) , .A1( u0_u0_X_5 ) , .ZN( u0_u0_u0_n31 ) );
  NOR2_X1 u0_u0_u0_U58 (.A2( u0_u0_X_5 ) , .A1( u0_u0_u0_n16 ) , .ZN( u0_u0_u0_n39 ) );
  NAND2_X1 u0_u0_u0_U59 (.A1( u0_u0_X_5 ) , .A2( u0_u0_u0_n16 ) , .ZN( u0_u0_u0_n37 ) );
  NOR2_X1 u0_u0_u0_U6 (.A2( u0_u0_u0_n17 ) , .ZN( u0_u0_u0_n52 ) , .A1( u0_u0_u0_n67 ) );
  AND2_X1 u0_u0_u0_U60 (.A2( u0_u0_X_3 ) , .A1( u0_u0_X_6 ) , .ZN( u0_u0_u0_n73 ) );
  AND2_X1 u0_u0_u0_U61 (.A1( u0_u0_X_6 ) , .A2( u0_u0_u0_n13 ) , .ZN( u0_u0_u0_n82 ) );
  INV_X1 u0_u0_u0_U62 (.A( u0_u0_X_4 ) , .ZN( u0_u0_u0_n16 ) );
  INV_X1 u0_u0_u0_U63 (.A( u0_u0_X_2 ) , .ZN( u0_u0_u0_n12 ) );
  INV_X1 u0_u0_u0_U64 (.A( u0_u0_X_3 ) , .ZN( u0_u0_u0_n13 ) );
  AOI211_X1 u0_u0_u0_U65 (.C1( u0_u0_u0_n15 ) , .C2( u0_u0_u0_n62 ) , .ZN( u0_u0_u0_n69 ) , .A( u0_u0_u0_n70 ) , .B( u0_u0_u0_n71 ) );
  INV_X1 u0_u0_u0_U66 (.ZN( u0_u0_u0_n1 ) , .A( u0_u0_u0_n86 ) );
  OR4_X1 u0_u0_u0_U67 (.ZN( u0_out0_17 ) , .A3( u0_u0_u0_n5 ) , .A1( u0_u0_u0_n51 ) , .A2( u0_u0_u0_n52 ) , .A4( u0_u0_u0_n53 ) );
  AOI21_X1 u0_u0_u0_U68 (.A( u0_u0_u0_n14 ) , .B1( u0_u0_u0_n47 ) , .ZN( u0_u0_u0_n51 ) , .B2( u0_u0_u0_n68 ) );
  INV_X1 u0_u0_u0_U69 (.ZN( u0_u0_u0_n5 ) , .A( u0_u0_u0_n64 ) );
  OAI21_X1 u0_u0_u0_U7 (.B2( u0_u0_u0_n17 ) , .B1( u0_u0_u0_n25 ) , .A( u0_u0_u0_n3 ) , .ZN( u0_u0_u0_n86 ) );
  OR4_X1 u0_u0_u0_U70 (.ZN( u0_out0_31 ) , .A1( u0_u0_u0_n18 ) , .A2( u0_u0_u0_n19 ) , .A3( u0_u0_u0_n2 ) , .A4( u0_u0_u0_n20 ) );
  AOI21_X1 u0_u0_u0_U71 (.ZN( u0_u0_u0_n18 ) , .B1( u0_u0_u0_n35 ) , .B2( u0_u0_u0_n36 ) , .A( u0_u0_u0_n37 ) );
  AOI21_X1 u0_u0_u0_U72 (.A( u0_u0_u0_n14 ) , .ZN( u0_u0_u0_n19 ) , .B1( u0_u0_u0_n33 ) , .B2( u0_u0_u0_n34 ) );
  INV_X1 u0_u0_u0_U73 (.A( u0_u0_u0_n49 ) , .ZN( u0_u0_u0_n7 ) );
  AOI211_X1 u0_u0_u0_U74 (.ZN( u0_u0_u0_n38 ) , .C1( u0_u0_u0_n39 ) , .C2( u0_u0_u0_n40 ) , .A( u0_u0_u0_n41 ) , .B( u0_u0_u0_n42 ) );
  NOR2_X1 u0_u0_u0_U75 (.A2( u0_u0_u0_n11 ) , .A1( u0_u0_u0_n12 ) , .ZN( u0_u0_u0_n80 ) );
  OAI221_X1 u0_u0_u0_U76 (.C2( u0_u0_u0_n28 ) , .B1( u0_u0_u0_n31 ) , .A( u0_u0_u0_n32 ) , .B2( u0_u0_u0_n48 ) , .ZN( u0_u0_u0_n53 ) , .C1( u0_u0_u0_n54 ) );
  INV_X1 u0_u0_u0_U77 (.A( u0_u0_X_1 ) , .ZN( u0_u0_u0_n11 ) );
  AOI21_X1 u0_u0_u0_U78 (.A( u0_u0_u0_n31 ) , .ZN( u0_u0_u0_n42 ) , .B1( u0_u0_u0_n43 ) , .B2( u0_u0_u0_n9 ) );
  OAI22_X1 u0_u0_u0_U79 (.B2( u0_u0_u0_n14 ) , .A1( u0_u0_u0_n28 ) , .B1( u0_u0_u0_n29 ) , .A2( u0_u0_u0_n43 ) , .ZN( u0_u0_u0_n70 ) );
  AND2_X1 u0_u0_u0_U8 (.ZN( u0_u0_u0_n29 ) , .A2( u0_u0_u0_n54 ) , .A1( u0_u0_u0_n61 ) );
  NAND2_X1 u0_u0_u0_U80 (.A1( u0_u0_u0_n30 ) , .A2( u0_u0_u0_n43 ) , .ZN( u0_u0_u0_n65 ) );
  INV_X1 u0_u0_u0_U81 (.A( u0_u0_u0_n56 ) , .ZN( u0_u0_u0_n8 ) );
  NAND2_X1 u0_u0_u0_U82 (.ZN( u0_u0_u0_n35 ) , .A2( u0_u0_u0_n72 ) , .A1( u0_u0_u0_n81 ) );
  NAND2_X1 u0_u0_u0_U83 (.ZN( u0_u0_u0_n45 ) , .A1( u0_u0_u0_n74 ) , .A2( u0_u0_u0_n81 ) );
  NAND2_X1 u0_u0_u0_U84 (.ZN( u0_u0_u0_n67 ) , .A2( u0_u0_u0_n81 ) , .A1( u0_u0_u0_n83 ) );
  NAND2_X1 u0_u0_u0_U85 (.ZN( u0_u0_u0_n33 ) , .A2( u0_u0_u0_n80 ) , .A1( u0_u0_u0_n81 ) );
  NOR2_X1 u0_u0_u0_U86 (.A2( u0_u0_X_6 ) , .A1( u0_u0_u0_n13 ) , .ZN( u0_u0_u0_n75 ) );
  NOR2_X1 u0_u0_u0_U87 (.A2( u0_u0_X_3 ) , .A1( u0_u0_X_6 ) , .ZN( u0_u0_u0_n81 ) );
  NAND3_X1 u0_u0_u0_U88 (.ZN( u0_out0_23 ) , .A3( u0_u0_u0_n38 ) , .A2( u0_u0_u0_n4 ) , .A1( u0_u0_u0_n7 ) );
  NAND3_X1 u0_u0_u0_U89 (.A1( u0_u0_u0_n25 ) , .ZN( u0_u0_u0_n40 ) , .A2( u0_u0_u0_n47 ) , .A3( u0_u0_u0_n48 ) );
  AND2_X1 u0_u0_u0_U9 (.A2( u0_u0_u0_n25 ) , .ZN( u0_u0_u0_n34 ) , .A1( u0_u0_u0_n44 ) );
  NAND3_X1 u0_u0_u0_U90 (.A1( u0_u0_u0_n27 ) , .A2( u0_u0_u0_n36 ) , .A3( u0_u0_u0_n43 ) , .ZN( u0_u0_u0_n58 ) );
  NAND3_X1 u0_u0_u0_U91 (.A1( u0_u0_u0_n26 ) , .A3( u0_u0_u0_n35 ) , .A2( u0_u0_u0_n61 ) , .ZN( u0_u0_u0_n66 ) );
  NAND3_X1 u0_u0_u0_U92 (.ZN( u0_out0_9 ) , .A1( u0_u0_u0_n1 ) , .A2( u0_u0_u0_n4 ) , .A3( u0_u0_u0_n69 ) );
  NAND3_X1 u0_u0_u0_U93 (.A3( u0_u0_u0_n29 ) , .A1( u0_u0_u0_n43 ) , .A2( u0_u0_u0_n47 ) , .ZN( u0_u0_u0_n78 ) );
  AOI21_X1 u0_u0_u1_U10 (.A( u0_u0_u1_n15 ) , .ZN( u0_u0_u1_n32 ) , .B1( u0_u0_u1_n33 ) , .B2( u0_u0_u1_n34 ) );
  NAND3_X1 u0_u0_u1_U100 (.A2( u0_u0_u1_n34 ) , .A3( u0_u0_u1_n56 ) , .A1( u0_u0_u1_n69 ) , .ZN( u0_u0_u1_n76 ) );
  NAND2_X1 u0_u0_u1_U11 (.A1( u0_u0_u1_n34 ) , .A2( u0_u0_u1_n39 ) , .ZN( u0_u0_u1_n49 ) );
  NAND2_X1 u0_u0_u1_U12 (.A2( u0_u0_u1_n36 ) , .ZN( u0_u0_u1_n42 ) , .A1( u0_u0_u1_n58 ) );
  AOI22_X1 u0_u0_u1_U13 (.B1( u0_u0_u1_n16 ) , .A1( u0_u0_u1_n18 ) , .ZN( u0_u0_u1_n46 ) , .A2( u0_u0_u1_n52 ) , .B2( u0_u0_u1_n53 ) );
  INV_X1 u0_u0_u1_U14 (.A( u0_u0_u1_n42 ) , .ZN( u0_u0_u1_n8 ) );
  INV_X1 u0_u0_u1_U15 (.ZN( u0_u0_u1_n15 ) , .A( u0_u0_u1_n50 ) );
  OR4_X1 u0_u0_u1_U16 (.A2( u0_u0_u1_n5 ) , .A1( u0_u0_u1_n72 ) , .ZN( u0_u0_u1_n81 ) , .A3( u0_u0_u1_n82 ) , .A4( u0_u0_u1_n83 ) );
  AOI21_X1 u0_u0_u1_U17 (.B2( u0_u0_u1_n33 ) , .B1( u0_u0_u1_n35 ) , .A( u0_u0_u1_n77 ) , .ZN( u0_u0_u1_n83 ) );
  AOI21_X1 u0_u0_u1_U18 (.A( u0_u0_u1_n15 ) , .B2( u0_u0_u1_n40 ) , .B1( u0_u0_u1_n55 ) , .ZN( u0_u0_u1_n82 ) );
  INV_X1 u0_u0_u1_U19 (.ZN( u0_u0_u1_n5 ) , .A( u0_u0_u1_n88 ) );
  INV_X1 u0_u0_u1_U20 (.ZN( u0_u0_u1_n18 ) , .A( u0_u0_u1_n77 ) );
  NAND2_X1 u0_u0_u1_U21 (.A2( u0_u0_u1_n33 ) , .A1( u0_u0_u1_n36 ) , .ZN( u0_u0_u1_n48 ) );
  AND2_X1 u0_u0_u1_U22 (.A2( u0_u0_u1_n28 ) , .ZN( u0_u0_u1_n55 ) , .A1( u0_u0_u1_n66 ) );
  NAND2_X1 u0_u0_u1_U23 (.ZN( u0_u0_u1_n41 ) , .A1( u0_u0_u1_n73 ) , .A2( u0_u0_u1_n74 ) );
  NAND2_X1 u0_u0_u1_U24 (.ZN( u0_u0_u1_n30 ) , .A1( u0_u0_u1_n54 ) , .A2( u0_u0_u1_n56 ) );
  NAND2_X1 u0_u0_u1_U25 (.ZN( u0_u0_u1_n57 ) , .A1( u0_u0_u1_n69 ) , .A2( u0_u0_u1_n74 ) );
  INV_X1 u0_u0_u1_U26 (.ZN( u0_u0_u1_n11 ) , .A( u0_u0_u1_n35 ) );
  INV_X1 u0_u0_u1_U27 (.A( u0_u0_u1_n38 ) , .ZN( u0_u0_u1_n6 ) );
  AND2_X1 u0_u0_u1_U28 (.ZN( u0_u0_u1_n40 ) , .A2( u0_u0_u1_n56 ) , .A1( u0_u0_u1_n60 ) );
  INV_X1 u0_u0_u1_U29 (.A( u0_u0_u1_n58 ) , .ZN( u0_u0_u1_n9 ) );
  INV_X1 u0_u0_u1_U3 (.A( u0_u0_u1_n30 ) , .ZN( u0_u0_u1_n7 ) );
  AOI221_X1 u0_u0_u1_U30 (.A( u0_u0_u1_n1 ) , .C1( u0_u0_u1_n11 ) , .C2( u0_u0_u1_n14 ) , .B2( u0_u0_u1_n17 ) , .ZN( u0_u0_u1_n22 ) , .B1( u0_u0_u1_n49 ) );
  INV_X1 u0_u0_u1_U31 (.ZN( u0_u0_u1_n1 ) , .A( u0_u0_u1_n92 ) );
  AOI211_X1 u0_u0_u1_U32 (.C2( u0_u0_u1_n50 ) , .C1( u0_u0_u1_n57 ) , .A( u0_u0_u1_n71 ) , .ZN( u0_u0_u1_n92 ) , .B( u0_u0_u1_n93 ) );
  AOI21_X1 u0_u0_u1_U33 (.A( u0_u0_u1_n37 ) , .B1( u0_u0_u1_n54 ) , .B2( u0_u0_u1_n68 ) , .ZN( u0_u0_u1_n93 ) );
  OAI221_X1 u0_u0_u1_U34 (.C1( u0_u0_u1_n15 ) , .B1( u0_u0_u1_n2 ) , .B2( u0_u0_u1_n37 ) , .ZN( u0_u0_u1_n51 ) , .C2( u0_u0_u1_n60 ) , .A( u0_u0_u1_n70 ) );
  INV_X1 u0_u0_u1_U35 (.ZN( u0_u0_u1_n2 ) , .A( u0_u0_u1_n41 ) );
  AOI211_X1 u0_u0_u1_U36 (.C1( u0_u0_u1_n30 ) , .C2( u0_u0_u1_n43 ) , .ZN( u0_u0_u1_n70 ) , .A( u0_u0_u1_n71 ) , .B( u0_u0_u1_n72 ) );
  NOR2_X1 u0_u0_u1_U37 (.A2( u0_u0_u1_n13 ) , .A1( u0_u0_u1_n21 ) , .ZN( u0_u0_u1_n91 ) );
  AOI211_X1 u0_u0_u1_U38 (.C1( u0_u0_u1_n18 ) , .ZN( u0_u0_u1_n24 ) , .C2( u0_u0_u1_n25 ) , .A( u0_u0_u1_n26 ) , .B( u0_u0_u1_n27 ) );
  AOI21_X1 u0_u0_u1_U39 (.ZN( u0_u0_u1_n27 ) , .B2( u0_u0_u1_n28 ) , .A( u0_u0_u1_n29 ) , .B1( u0_u0_u1_n7 ) );
  AOI221_X1 u0_u0_u1_U4 (.B1( u0_u0_u1_n14 ) , .ZN( u0_u0_u1_n47 ) , .B2( u0_u0_u1_n48 ) , .C1( u0_u0_u1_n49 ) , .C2( u0_u0_u1_n50 ) , .A( u0_u0_u1_n51 ) );
  OR2_X1 u0_u0_u1_U40 (.ZN( u0_u0_u1_n26 ) , .A1( u0_u0_u1_n31 ) , .A2( u0_u0_u1_n32 ) );
  NAND2_X1 u0_u0_u1_U41 (.A2( u0_u0_u1_n29 ) , .ZN( u0_u0_u1_n43 ) , .A1( u0_u0_u1_n61 ) );
  NAND2_X1 u0_u0_u1_U42 (.A1( u0_u0_u1_n37 ) , .ZN( u0_u0_u1_n50 ) , .A2( u0_u0_u1_n77 ) );
  NAND2_X1 u0_u0_u1_U43 (.ZN( u0_u0_u1_n33 ) , .A1( u0_u0_u1_n84 ) , .A2( u0_u0_u1_n90 ) );
  NOR2_X1 u0_u0_u1_U44 (.A2( u0_u0_u1_n29 ) , .A1( u0_u0_u1_n68 ) , .ZN( u0_u0_u1_n72 ) );
  AOI21_X1 u0_u0_u1_U45 (.B1( u0_u0_u1_n39 ) , .ZN( u0_u0_u1_n59 ) , .B2( u0_u0_u1_n60 ) , .A( u0_u0_u1_n61 ) );
  NAND2_X1 u0_u0_u1_U46 (.A2( u0_u0_u1_n19 ) , .A1( u0_u0_u1_n20 ) , .ZN( u0_u0_u1_n77 ) );
  NAND2_X1 u0_u0_u1_U47 (.ZN( u0_u0_u1_n60 ) , .A1( u0_u0_u1_n91 ) , .A2( u0_u0_u1_n94 ) );
  NAND2_X1 u0_u0_u1_U48 (.ZN( u0_u0_u1_n35 ) , .A1( u0_u0_u1_n87 ) , .A2( u0_u0_u1_n90 ) );
  NAND2_X1 u0_u0_u1_U49 (.ZN( u0_u0_u1_n54 ) , .A2( u0_u0_u1_n89 ) , .A1( u0_u0_u1_n90 ) );
  AOI211_X1 u0_u0_u1_U5 (.C1( u0_u0_u1_n42 ) , .B( u0_u0_u1_n44 ) , .C2( u0_u0_u1_n50 ) , .A( u0_u0_u1_n51 ) , .ZN( u0_u0_u1_n65 ) );
  AOI21_X1 u0_u0_u1_U50 (.ZN( u0_u0_u1_n31 ) , .B1( u0_u0_u1_n35 ) , .B2( u0_u0_u1_n36 ) , .A( u0_u0_u1_n37 ) );
  INV_X1 u0_u0_u1_U51 (.ZN( u0_u0_u1_n14 ) , .A( u0_u0_u1_n29 ) );
  NAND2_X1 u0_u0_u1_U52 (.ZN( u0_u0_u1_n73 ) , .A1( u0_u0_u1_n89 ) , .A2( u0_u0_u1_n94 ) );
  NAND2_X1 u0_u0_u1_U53 (.ZN( u0_u0_u1_n58 ) , .A1( u0_u0_u1_n87 ) , .A2( u0_u0_u1_n94 ) );
  NAND2_X1 u0_u0_u1_U54 (.ZN( u0_u0_u1_n68 ) , .A2( u0_u0_u1_n85 ) , .A1( u0_u0_u1_n91 ) );
  NAND2_X1 u0_u0_u1_U55 (.ZN( u0_u0_u1_n36 ) , .A1( u0_u0_u1_n86 ) , .A2( u0_u0_u1_n91 ) );
  NAND2_X1 u0_u0_u1_U56 (.ZN( u0_u0_u1_n56 ) , .A1( u0_u0_u1_n84 ) , .A2( u0_u0_u1_n85 ) );
  NAND2_X1 u0_u0_u1_U57 (.ZN( u0_u0_u1_n39 ) , .A1( u0_u0_u1_n90 ) , .A2( u0_u0_u1_n91 ) );
  NAND2_X1 u0_u0_u1_U58 (.ZN( u0_u0_u1_n34 ) , .A1( u0_u0_u1_n84 ) , .A2( u0_u0_u1_n94 ) );
  OAI21_X1 u0_u0_u1_U59 (.A( u0_u0_u1_n22 ) , .B2( u0_u0_u1_n29 ) , .B1( u0_u0_u1_n60 ) , .ZN( u0_u0_u1_n80 ) );
  AOI22_X1 u0_u0_u1_U6 (.B1( u0_u0_u1_n16 ) , .A1( u0_u0_u1_n18 ) , .ZN( u0_u0_u1_n64 ) , .A2( u0_u0_u1_n75 ) , .B2( u0_u0_u1_n76 ) );
  NAND2_X1 u0_u0_u1_U60 (.ZN( u0_u0_u1_n69 ) , .A1( u0_u0_u1_n86 ) , .A2( u0_u0_u1_n89 ) );
  NAND2_X1 u0_u0_u1_U61 (.ZN( u0_u0_u1_n74 ) , .A2( u0_u0_u1_n85 ) , .A1( u0_u0_u1_n87 ) );
  NAND2_X1 u0_u0_u1_U62 (.ZN( u0_u0_u1_n38 ) , .A1( u0_u0_u1_n85 ) , .A2( u0_u0_u1_n89 ) );
  NAND2_X1 u0_u0_u1_U63 (.ZN( u0_u0_u1_n28 ) , .A1( u0_u0_u1_n84 ) , .A2( u0_u0_u1_n86 ) );
  INV_X1 u0_u0_u1_U64 (.ZN( u0_u0_u1_n16 ) , .A( u0_u0_u1_n37 ) );
  INV_X1 u0_u0_u1_U65 (.ZN( u0_u0_u1_n17 ) , .A( u0_u0_u1_n61 ) );
  NAND2_X1 u0_u0_u1_U66 (.ZN( u0_u0_u1_n66 ) , .A1( u0_u0_u1_n86 ) , .A2( u0_u0_u1_n87 ) );
  OAI21_X1 u0_u0_u1_U67 (.B1( u0_u0_u1_n29 ) , .A( u0_u0_u1_n4 ) , .ZN( u0_u0_u1_n44 ) , .B2( u0_u0_u1_n66 ) );
  INV_X1 u0_u0_u1_U68 (.ZN( u0_u0_u1_n4 ) , .A( u0_u0_u1_n67 ) );
  AOI21_X1 u0_u0_u1_U69 (.A( u0_u0_u1_n61 ) , .ZN( u0_u0_u1_n67 ) , .B1( u0_u0_u1_n68 ) , .B2( u0_u0_u1_n69 ) );
  NAND2_X1 u0_u0_u1_U7 (.A2( u0_u0_u1_n33 ) , .A1( u0_u0_u1_n55 ) , .ZN( u0_u0_u1_n75 ) );
  NOR2_X1 u0_u0_u1_U70 (.A2( u0_u0_X_7 ) , .A1( u0_u0_X_8 ) , .ZN( u0_u0_u1_n94 ) );
  NOR2_X1 u0_u0_u1_U71 (.A1( u0_u0_X_12 ) , .A2( u0_u0_X_9 ) , .ZN( u0_u0_u1_n89 ) );
  NOR2_X1 u0_u0_u1_U72 (.A2( u0_u0_X_8 ) , .A1( u0_u0_u1_n12 ) , .ZN( u0_u0_u1_n90 ) );
  NOR2_X1 u0_u0_u1_U73 (.A2( u0_u0_X_12 ) , .A1( u0_u0_u1_n13 ) , .ZN( u0_u0_u1_n87 ) );
  NOR2_X1 u0_u0_u1_U74 (.A2( u0_u0_X_9 ) , .A1( u0_u0_u1_n21 ) , .ZN( u0_u0_u1_n84 ) );
  NAND2_X1 u0_u0_u1_U75 (.A1( u0_u0_X_10 ) , .A2( u0_u0_u1_n20 ) , .ZN( u0_u0_u1_n29 ) );
  NAND2_X1 u0_u0_u1_U76 (.A2( u0_u0_X_10 ) , .A1( u0_u0_X_11 ) , .ZN( u0_u0_u1_n37 ) );
  NAND2_X1 u0_u0_u1_U77 (.A1( u0_u0_X_11 ) , .A2( u0_u0_u1_n19 ) , .ZN( u0_u0_u1_n61 ) );
  AND2_X1 u0_u0_u1_U78 (.A2( u0_u0_X_7 ) , .A1( u0_u0_X_8 ) , .ZN( u0_u0_u1_n85 ) );
  AND2_X1 u0_u0_u1_U79 (.A1( u0_u0_X_8 ) , .A2( u0_u0_u1_n12 ) , .ZN( u0_u0_u1_n86 ) );
  NOR2_X1 u0_u0_u1_U8 (.ZN( u0_u0_u1_n71 ) , .A2( u0_u0_u1_n73 ) , .A1( u0_u0_u1_n77 ) );
  INV_X1 u0_u0_u1_U80 (.A( u0_u0_X_10 ) , .ZN( u0_u0_u1_n19 ) );
  INV_X1 u0_u0_u1_U81 (.A( u0_u0_X_9 ) , .ZN( u0_u0_u1_n13 ) );
  INV_X1 u0_u0_u1_U82 (.A( u0_u0_X_11 ) , .ZN( u0_u0_u1_n20 ) );
  INV_X1 u0_u0_u1_U83 (.A( u0_u0_X_12 ) , .ZN( u0_u0_u1_n21 ) );
  INV_X1 u0_u0_u1_U84 (.A( u0_u0_X_7 ) , .ZN( u0_u0_u1_n12 ) );
  NAND4_X1 u0_u0_u1_U85 (.ZN( u0_out0_18 ) , .A1( u0_u0_u1_n22 ) , .A3( u0_u0_u1_n23 ) , .A4( u0_u0_u1_n24 ) , .A2( u0_u0_u1_n3 ) );
  AOI22_X1 u0_u0_u1_U86 (.A1( u0_u0_u1_n17 ) , .ZN( u0_u0_u1_n23 ) , .A2( u0_u0_u1_n41 ) , .B1( u0_u0_u1_n42 ) , .B2( u0_u0_u1_n43 ) );
  INV_X1 u0_u0_u1_U87 (.ZN( u0_u0_u1_n3 ) , .A( u0_u0_u1_n44 ) );
  NAND4_X1 u0_u0_u1_U88 (.ZN( u0_out0_2 ) , .A1( u0_u0_u1_n10 ) , .A2( u0_u0_u1_n45 ) , .A3( u0_u0_u1_n46 ) , .A4( u0_u0_u1_n47 ) );
  OAI21_X1 u0_u0_u1_U89 (.A( u0_u0_u1_n43 ) , .ZN( u0_u0_u1_n45 ) , .B2( u0_u0_u1_n57 ) , .B1( u0_u0_u1_n9 ) );
  OAI21_X1 u0_u0_u1_U9 (.A( u0_u0_u1_n43 ) , .B1( u0_u0_u1_n48 ) , .B2( u0_u0_u1_n6 ) , .ZN( u0_u0_u1_n88 ) );
  INV_X1 u0_u0_u1_U90 (.ZN( u0_u0_u1_n10 ) , .A( u0_u0_u1_n59 ) );
  NAND4_X1 u0_u0_u1_U91 (.ZN( u0_out0_28 ) , .A1( u0_u0_u1_n62 ) , .A2( u0_u0_u1_n63 ) , .A3( u0_u0_u1_n64 ) , .A4( u0_u0_u1_n65 ) );
  OAI21_X1 u0_u0_u1_U92 (.B1( u0_u0_u1_n14 ) , .B2( u0_u0_u1_n50 ) , .A( u0_u0_u1_n6 ) , .ZN( u0_u0_u1_n62 ) );
  OAI21_X1 u0_u0_u1_U93 (.B1( u0_u0_u1_n11 ) , .A( u0_u0_u1_n43 ) , .B2( u0_u0_u1_n49 ) , .ZN( u0_u0_u1_n63 ) );
  OR4_X1 u0_u0_u1_U94 (.ZN( u0_out0_13 ) , .A1( u0_u0_u1_n78 ) , .A2( u0_u0_u1_n79 ) , .A3( u0_u0_u1_n80 ) , .A4( u0_u0_u1_n81 ) );
  AOI21_X1 u0_u0_u1_U95 (.B1( u0_u0_u1_n54 ) , .B2( u0_u0_u1_n58 ) , .A( u0_u0_u1_n61 ) , .ZN( u0_u0_u1_n78 ) );
  AOI21_X1 u0_u0_u1_U96 (.B2( u0_u0_u1_n29 ) , .B1( u0_u0_u1_n37 ) , .A( u0_u0_u1_n73 ) , .ZN( u0_u0_u1_n79 ) );
  NAND3_X1 u0_u0_u1_U97 (.ZN( u0_u0_u1_n25 ) , .A1( u0_u0_u1_n38 ) , .A2( u0_u0_u1_n39 ) , .A3( u0_u0_u1_n40 ) );
  NAND3_X1 u0_u0_u1_U98 (.A1( u0_u0_u1_n38 ) , .ZN( u0_u0_u1_n53 ) , .A2( u0_u0_u1_n54 ) , .A3( u0_u0_u1_n55 ) );
  NAND3_X1 u0_u0_u1_U99 (.A2( u0_u0_u1_n35 ) , .ZN( u0_u0_u1_n52 ) , .A1( u0_u0_u1_n56 ) , .A3( u0_u0_u1_n8 ) );
  OAI22_X1 u0_u0_u3_U10 (.B2( u0_u0_u3_n23 ) , .A1( u0_u0_u3_n37 ) , .A2( u0_u0_u3_n52 ) , .B1( u0_u0_u3_n74 ) , .ZN( u0_u0_u3_n89 ) );
  OAI211_X1 u0_u0_u3_U11 (.C1( u0_u0_u3_n20 ) , .C2( u0_u0_u3_n59 ) , .A( u0_u0_u3_n6 ) , .ZN( u0_u0_u3_n68 ) , .B( u0_u0_u3_n81 ) );
  AOI221_X1 u0_u0_u3_U12 (.B1( u0_u0_u3_n18 ) , .C2( u0_u0_u3_n54 ) , .B2( u0_u0_u3_n55 ) , .A( u0_u0_u3_n56 ) , .ZN( u0_u0_u3_n81 ) , .C1( u0_u0_u3_n82 ) );
  INV_X1 u0_u0_u3_U13 (.ZN( u0_u0_u3_n6 ) , .A( u0_u0_u3_n89 ) );
  NAND2_X1 u0_u0_u3_U14 (.A1( u0_u0_u3_n32 ) , .A2( u0_u0_u3_n57 ) , .ZN( u0_u0_u3_n82 ) );
  AOI22_X1 u0_u0_u3_U15 (.A1( u0_u0_u3_n18 ) , .B2( u0_u0_u3_n54 ) , .ZN( u0_u0_u3_n64 ) , .A2( u0_u0_u3_n71 ) , .B1( u0_u0_u3_n72 ) );
  NAND2_X1 u0_u0_u3_U16 (.A2( u0_u0_u3_n36 ) , .A1( u0_u0_u3_n5 ) , .ZN( u0_u0_u3_n71 ) );
  NOR2_X1 u0_u0_u3_U17 (.A1( u0_u0_u3_n23 ) , .A2( u0_u0_u3_n37 ) , .ZN( u0_u0_u3_n61 ) );
  AOI21_X1 u0_u0_u3_U18 (.A( u0_u0_u3_n20 ) , .B1( u0_u0_u3_n32 ) , .B2( u0_u0_u3_n41 ) , .ZN( u0_u0_u3_n75 ) );
  NAND2_X1 u0_u0_u3_U19 (.A2( u0_u0_u3_n23 ) , .ZN( u0_u0_u3_n45 ) , .A1( u0_u0_u3_n52 ) );
  NAND2_X1 u0_u0_u3_U20 (.A1( u0_u0_u3_n31 ) , .A2( u0_u0_u3_n35 ) , .ZN( u0_u0_u3_n55 ) );
  INV_X1 u0_u0_u3_U21 (.ZN( u0_u0_u3_n22 ) , .A( u0_u0_u3_n54 ) );
  AND2_X1 u0_u0_u3_U22 (.ZN( u0_u0_u3_n36 ) , .A1( u0_u0_u3_n73 ) , .A2( u0_u0_u3_n74 ) );
  INV_X1 u0_u0_u3_U23 (.ZN( u0_u0_u3_n17 ) , .A( u0_u0_u3_n52 ) );
  NAND2_X1 u0_u0_u3_U24 (.ZN( u0_u0_u3_n47 ) , .A2( u0_u0_u3_n79 ) , .A1( u0_u0_u3_n80 ) );
  NAND2_X1 u0_u0_u3_U25 (.A2( u0_u0_u3_n39 ) , .A1( u0_u0_u3_n63 ) , .ZN( u0_u0_u3_n70 ) );
  NAND2_X1 u0_u0_u3_U26 (.A2( u0_u0_u3_n20 ) , .A1( u0_u0_u3_n22 ) , .ZN( u0_u0_u3_n44 ) );
  INV_X1 u0_u0_u3_U27 (.ZN( u0_u0_u3_n10 ) , .A( u0_u0_u3_n57 ) );
  INV_X1 u0_u0_u3_U28 (.ZN( u0_u0_u3_n11 ) , .A( u0_u0_u3_n59 ) );
  INV_X1 u0_u0_u3_U29 (.ZN( u0_u0_u3_n13 ) , .A( u0_u0_u3_n32 ) );
  INV_X1 u0_u0_u3_U3 (.A( u0_u0_u3_n47 ) , .ZN( u0_u0_u3_n5 ) );
  INV_X1 u0_u0_u3_U30 (.ZN( u0_u0_u3_n2 ) , .A( u0_u0_u3_n48 ) );
  NOR2_X1 u0_u0_u3_U31 (.A1( u0_u0_u3_n18 ) , .A2( u0_u0_u3_n46 ) , .ZN( u0_u0_u3_n52 ) );
  OAI222_X1 u0_u0_u3_U32 (.A1( u0_u0_u3_n23 ) , .C1( u0_u0_u3_n33 ) , .B2( u0_u0_u3_n41 ) , .ZN( u0_u0_u3_n49 ) , .B1( u0_u0_u3_n52 ) , .A2( u0_u0_u3_n79 ) , .C2( u0_u0_u3_n80 ) );
  NOR4_X1 u0_u0_u3_U33 (.ZN( u0_u0_u3_n26 ) , .A1( u0_u0_u3_n27 ) , .A2( u0_u0_u3_n28 ) , .A3( u0_u0_u3_n29 ) , .A4( u0_u0_u3_n30 ) );
  AOI21_X1 u0_u0_u3_U34 (.A( u0_u0_u3_n23 ) , .ZN( u0_u0_u3_n29 ) , .B1( u0_u0_u3_n34 ) , .B2( u0_u0_u3_n35 ) );
  AOI21_X1 u0_u0_u3_U35 (.ZN( u0_u0_u3_n30 ) , .B1( u0_u0_u3_n31 ) , .B2( u0_u0_u3_n32 ) , .A( u0_u0_u3_n33 ) );
  AOI21_X1 u0_u0_u3_U36 (.ZN( u0_u0_u3_n28 ) , .B1( u0_u0_u3_n36 ) , .B2( u0_u0_u3_n37 ) , .A( u0_u0_u3_n38 ) );
  OAI211_X1 u0_u0_u3_U37 (.A( u0_u0_u3_n3 ) , .C2( u0_u0_u3_n33 ) , .C1( u0_u0_u3_n37 ) , .ZN( u0_u0_u3_n48 ) , .B( u0_u0_u3_n60 ) );
  INV_X1 u0_u0_u3_U38 (.ZN( u0_u0_u3_n3 ) , .A( u0_u0_u3_n62 ) );
  AOI221_X1 u0_u0_u3_U39 (.B1( u0_u0_u3_n13 ) , .B2( u0_u0_u3_n17 ) , .C1( u0_u0_u3_n18 ) , .C2( u0_u0_u3_n55 ) , .ZN( u0_u0_u3_n60 ) , .A( u0_u0_u3_n61 ) );
  INV_X1 u0_u0_u3_U4 (.ZN( u0_u0_u3_n4 ) , .A( u0_u0_u3_n58 ) );
  OAI22_X1 u0_u0_u3_U40 (.B1( u0_u0_u3_n20 ) , .A2( u0_u0_u3_n22 ) , .B2( u0_u0_u3_n42 ) , .ZN( u0_u0_u3_n62 ) , .A1( u0_u0_u3_n63 ) );
  AOI211_X1 u0_u0_u3_U41 (.C1( u0_u0_u3_n46 ) , .B( u0_u0_u3_n49 ) , .C2( u0_u0_u3_n58 ) , .A( u0_u0_u3_n68 ) , .ZN( u0_u0_u3_n78 ) );
  AOI211_X1 u0_u0_u3_U42 (.ZN( u0_u0_u3_n65 ) , .C2( u0_u0_u3_n66 ) , .A( u0_u0_u3_n67 ) , .B( u0_u0_u3_n68 ) , .C1( u0_u0_u3_n8 ) );
  INV_X1 u0_u0_u3_U43 (.A( u0_u0_u3_n31 ) , .ZN( u0_u0_u3_n8 ) );
  OAI22_X1 u0_u0_u3_U44 (.B2( u0_u0_u3_n33 ) , .A1( u0_u0_u3_n52 ) , .ZN( u0_u0_u3_n67 ) , .B1( u0_u0_u3_n69 ) , .A2( u0_u0_u3_n9 ) );
  AND3_X1 u0_u0_u3_U45 (.A3( u0_u0_u3_n35 ) , .A1( u0_u0_u3_n43 ) , .A2( u0_u0_u3_n63 ) , .ZN( u0_u0_u3_n69 ) );
  INV_X1 u0_u0_u3_U46 (.ZN( u0_u0_u3_n23 ) , .A( u0_u0_u3_n66 ) );
  NAND2_X1 u0_u0_u3_U47 (.A2( u0_u0_u3_n23 ) , .A1( u0_u0_u3_n33 ) , .ZN( u0_u0_u3_n54 ) );
  NOR2_X1 u0_u0_u3_U48 (.A2( u0_u0_u3_n33 ) , .ZN( u0_u0_u3_n56 ) , .A1( u0_u0_u3_n74 ) );
  NAND2_X1 u0_u0_u3_U49 (.ZN( u0_u0_u3_n37 ) , .A1( u0_u0_u3_n84 ) , .A2( u0_u0_u3_n88 ) );
  INV_X1 u0_u0_u3_U5 (.A( u0_u0_u3_n70 ) , .ZN( u0_u0_u3_n9 ) );
  NAND2_X1 u0_u0_u3_U50 (.ZN( u0_u0_u3_n32 ) , .A2( u0_u0_u3_n85 ) , .A1( u0_u0_u3_n90 ) );
  INV_X1 u0_u0_u3_U51 (.ZN( u0_u0_u3_n20 ) , .A( u0_u0_u3_n46 ) );
  AOI21_X1 u0_u0_u3_U52 (.A( u0_u0_u3_n33 ) , .B1( u0_u0_u3_n41 ) , .B2( u0_u0_u3_n73 ) , .ZN( u0_u0_u3_n93 ) );
  AOI21_X1 u0_u0_u3_U53 (.B1( u0_u0_u3_n1 ) , .B2( u0_u0_u3_n45 ) , .ZN( u0_u0_u3_n77 ) , .A( u0_u0_u3_n92 ) );
  INV_X1 u0_u0_u3_U54 (.ZN( u0_u0_u3_n1 ) , .A( u0_u0_u3_n42 ) );
  AOI21_X1 u0_u0_u3_U55 (.B2( u0_u0_u3_n32 ) , .A( u0_u0_u3_n38 ) , .B1( u0_u0_u3_n63 ) , .ZN( u0_u0_u3_n92 ) );
  INV_X1 u0_u0_u3_U56 (.ZN( u0_u0_u3_n18 ) , .A( u0_u0_u3_n38 ) );
  NAND2_X1 u0_u0_u3_U57 (.ZN( u0_u0_u3_n63 ) , .A2( u0_u0_u3_n90 ) , .A1( u0_u0_u3_n91 ) );
  NAND2_X1 u0_u0_u3_U58 (.ZN( u0_u0_u3_n41 ) , .A2( u0_u0_u3_n87 ) , .A1( u0_u0_u3_n91 ) );
  NAND2_X1 u0_u0_u3_U59 (.ZN( u0_u0_u3_n42 ) , .A1( u0_u0_u3_n86 ) , .A2( u0_u0_u3_n88 ) );
  AOI221_X1 u0_u0_u3_U6 (.B2( u0_u0_u3_n10 ) , .B1( u0_u0_u3_n44 ) , .ZN( u0_u0_u3_n53 ) , .C1( u0_u0_u3_n54 ) , .C2( u0_u0_u3_n55 ) , .A( u0_u0_u3_n56 ) );
  NAND2_X1 u0_u0_u3_U60 (.ZN( u0_u0_u3_n31 ) , .A1( u0_u0_u3_n87 ) , .A2( u0_u0_u3_n88 ) );
  NAND2_X1 u0_u0_u3_U61 (.ZN( u0_u0_u3_n39 ) , .A1( u0_u0_u3_n83 ) , .A2( u0_u0_u3_n86 ) );
  NAND2_X1 u0_u0_u3_U62 (.ZN( u0_u0_u3_n59 ) , .A2( u0_u0_u3_n85 ) , .A1( u0_u0_u3_n87 ) );
  NAND2_X1 u0_u0_u3_U63 (.ZN( u0_u0_u3_n35 ) , .A1( u0_u0_u3_n85 ) , .A2( u0_u0_u3_n86 ) );
  NAND2_X1 u0_u0_u3_U64 (.ZN( u0_u0_u3_n73 ) , .A2( u0_u0_u3_n86 ) , .A1( u0_u0_u3_n91 ) );
  NAND2_X1 u0_u0_u3_U65 (.ZN( u0_u0_u3_n80 ) , .A2( u0_u0_u3_n88 ) , .A1( u0_u0_u3_n90 ) );
  NAND2_X1 u0_u0_u3_U66 (.ZN( u0_u0_u3_n74 ) , .A1( u0_u0_u3_n83 ) , .A2( u0_u0_u3_n87 ) );
  NAND2_X1 u0_u0_u3_U67 (.ZN( u0_u0_u3_n34 ) , .A1( u0_u0_u3_n83 ) , .A2( u0_u0_u3_n90 ) );
  NAND2_X1 u0_u0_u3_U68 (.ZN( u0_u0_u3_n57 ) , .A1( u0_u0_u3_n83 ) , .A2( u0_u0_u3_n84 ) );
  NAND2_X1 u0_u0_u3_U69 (.ZN( u0_u0_u3_n43 ) , .A2( u0_u0_u3_n84 ) , .A1( u0_u0_u3_n91 ) );
  OAI22_X1 u0_u0_u3_U7 (.A1( u0_u0_u3_n19 ) , .B1( u0_u0_u3_n22 ) , .ZN( u0_u0_u3_n27 ) , .A2( u0_u0_u3_n39 ) , .B2( u0_u0_u3_n40 ) );
  NAND2_X1 u0_u0_u3_U70 (.ZN( u0_u0_u3_n79 ) , .A2( u0_u0_u3_n84 ) , .A1( u0_u0_u3_n85 ) );
  NOR2_X1 u0_u0_u3_U71 (.A2( u0_u0_X_19 ) , .A1( u0_u0_X_20 ) , .ZN( u0_u0_u3_n88 ) );
  NOR2_X1 u0_u0_u3_U72 (.A2( u0_u0_X_21 ) , .A1( u0_u0_X_24 ) , .ZN( u0_u0_u3_n84 ) );
  NOR2_X1 u0_u0_u3_U73 (.A2( u0_u0_X_24 ) , .A1( u0_u0_u3_n16 ) , .ZN( u0_u0_u3_n90 ) );
  NOR2_X1 u0_u0_u3_U74 (.A2( u0_u0_X_23 ) , .A1( u0_u0_u3_n21 ) , .ZN( u0_u0_u3_n46 ) );
  NOR2_X1 u0_u0_u3_U75 (.A2( u0_u0_X_19 ) , .A1( u0_u0_u3_n15 ) , .ZN( u0_u0_u3_n91 ) );
  NAND2_X1 u0_u0_u3_U76 (.A1( u0_u0_X_22 ) , .A2( u0_u0_X_23 ) , .ZN( u0_u0_u3_n33 ) );
  NAND2_X1 u0_u0_u3_U77 (.A1( u0_u0_X_23 ) , .A2( u0_u0_u3_n21 ) , .ZN( u0_u0_u3_n38 ) );
  NOR2_X1 u0_u0_u3_U78 (.A2( u0_u0_X_22 ) , .A1( u0_u0_X_23 ) , .ZN( u0_u0_u3_n66 ) );
  AND2_X1 u0_u0_u3_U79 (.A1( u0_u0_X_24 ) , .A2( u0_u0_u3_n16 ) , .ZN( u0_u0_u3_n86 ) );
  AND3_X1 u0_u0_u3_U8 (.ZN( u0_u0_u3_n40 ) , .A1( u0_u0_u3_n41 ) , .A2( u0_u0_u3_n42 ) , .A3( u0_u0_u3_n43 ) );
  AND2_X1 u0_u0_u3_U80 (.A1( u0_u0_X_19 ) , .A2( u0_u0_u3_n15 ) , .ZN( u0_u0_u3_n85 ) );
  AND2_X1 u0_u0_u3_U81 (.A1( u0_u0_X_21 ) , .A2( u0_u0_X_24 ) , .ZN( u0_u0_u3_n87 ) );
  AND2_X1 u0_u0_u3_U82 (.A2( u0_u0_X_19 ) , .A1( u0_u0_X_20 ) , .ZN( u0_u0_u3_n83 ) );
  INV_X1 u0_u0_u3_U83 (.A( u0_u0_X_22 ) , .ZN( u0_u0_u3_n21 ) );
  INV_X1 u0_u0_u3_U84 (.A( u0_u0_X_21 ) , .ZN( u0_u0_u3_n16 ) );
  INV_X1 u0_u0_u3_U85 (.A( u0_u0_X_20 ) , .ZN( u0_u0_u3_n15 ) );
  NAND4_X1 u0_u0_u3_U86 (.ZN( u0_out0_26 ) , .A1( u0_u0_u3_n14 ) , .A2( u0_u0_u3_n76 ) , .A3( u0_u0_u3_n77 ) , .A4( u0_u0_u3_n78 ) );
  INV_X1 u0_u0_u3_U87 (.ZN( u0_u0_u3_n14 ) , .A( u0_u0_u3_n93 ) );
  OAI21_X1 u0_u0_u3_U88 (.B1( u0_u0_u3_n11 ) , .A( u0_u0_u3_n54 ) , .B2( u0_u0_u3_n70 ) , .ZN( u0_u0_u3_n76 ) );
  NAND4_X1 u0_u0_u3_U89 (.ZN( u0_out0_1 ) , .A1( u0_u0_u3_n2 ) , .A2( u0_u0_u3_n24 ) , .A3( u0_u0_u3_n25 ) , .A4( u0_u0_u3_n26 ) );
  INV_X1 u0_u0_u3_U9 (.ZN( u0_u0_u3_n19 ) , .A( u0_u0_u3_n44 ) );
  NAND2_X1 u0_u0_u3_U90 (.A1( u0_u0_u3_n11 ) , .A2( u0_u0_u3_n17 ) , .ZN( u0_u0_u3_n24 ) );
  AOI22_X1 u0_u0_u3_U91 (.A1( u0_u0_u3_n10 ) , .ZN( u0_u0_u3_n25 ) , .A2( u0_u0_u3_n45 ) , .B1( u0_u0_u3_n46 ) , .B2( u0_u0_u3_n47 ) );
  NAND4_X1 u0_u0_u3_U92 (.ZN( u0_out0_20 ) , .A1( u0_u0_u3_n12 ) , .A3( u0_u0_u3_n64 ) , .A4( u0_u0_u3_n65 ) , .A2( u0_u0_u3_n7 ) );
  INV_X1 u0_u0_u3_U93 (.A( u0_u0_u3_n61 ) , .ZN( u0_u0_u3_n7 ) );
  INV_X1 u0_u0_u3_U94 (.ZN( u0_u0_u3_n12 ) , .A( u0_u0_u3_n75 ) );
  OR4_X1 u0_u0_u3_U95 (.ZN( u0_out0_10 ) , .A2( u0_u0_u3_n48 ) , .A1( u0_u0_u3_n49 ) , .A3( u0_u0_u3_n50 ) , .A4( u0_u0_u3_n51 ) );
  OAI222_X1 u0_u0_u3_U96 (.A1( u0_u0_u3_n20 ) , .C2( u0_u0_u3_n23 ) , .B2( u0_u0_u3_n33 ) , .A2( u0_u0_u3_n37 ) , .B1( u0_u0_u3_n39 ) , .ZN( u0_u0_u3_n50 ) , .C1( u0_u0_u3_n59 ) );
  OAI221_X1 u0_u0_u3_U97 (.B1( u0_u0_u3_n36 ) , .C1( u0_u0_u3_n38 ) , .C2( u0_u0_u3_n4 ) , .ZN( u0_u0_u3_n51 ) , .B2( u0_u0_u3_n52 ) , .A( u0_u0_u3_n53 ) );
  NAND3_X1 u0_u0_u3_U98 (.A3( u0_u0_u3_n34 ) , .A2( u0_u0_u3_n42 ) , .ZN( u0_u0_u3_n72 ) , .A1( u0_u0_u3_n73 ) );
  NAND3_X1 u0_u0_u3_U99 (.A1( u0_u0_u3_n34 ) , .A2( u0_u0_u3_n43 ) , .A3( u0_u0_u3_n5 ) , .ZN( u0_u0_u3_n58 ) );
  XOR2_X1 u0_u12_U13 (.B( u0_K13_42 ) , .A( u0_R11_29 ) , .Z( u0_u12_X_42 ) );
  XOR2_X1 u0_u12_U14 (.B( u0_K13_41 ) , .A( u0_R11_28 ) , .Z( u0_u12_X_41 ) );
  XOR2_X1 u0_u12_U15 (.B( u0_K13_40 ) , .A( u0_R11_27 ) , .Z( u0_u12_X_40 ) );
  XOR2_X1 u0_u12_U17 (.B( u0_K13_39 ) , .A( u0_R11_26 ) , .Z( u0_u12_X_39 ) );
  XOR2_X1 u0_u12_U18 (.B( u0_K13_38 ) , .A( u0_R11_25 ) , .Z( u0_u12_X_38 ) );
  XOR2_X1 u0_u12_U19 (.B( u0_K13_37 ) , .A( u0_R11_24 ) , .Z( u0_u12_X_37 ) );
  XOR2_X1 u0_u12_U20 (.B( u0_K13_36 ) , .A( u0_R11_25 ) , .Z( u0_u12_X_36 ) );
  XOR2_X1 u0_u12_U21 (.B( u0_K13_35 ) , .A( u0_R11_24 ) , .Z( u0_u12_X_35 ) );
  XOR2_X1 u0_u12_U22 (.B( u0_K13_34 ) , .A( u0_R11_23 ) , .Z( u0_u12_X_34 ) );
  XOR2_X1 u0_u12_U23 (.B( u0_K13_33 ) , .A( u0_R11_22 ) , .Z( u0_u12_X_33 ) );
  XOR2_X1 u0_u12_U24 (.B( u0_K13_32 ) , .A( u0_R11_21 ) , .Z( u0_u12_X_32 ) );
  XOR2_X1 u0_u12_U25 (.B( u0_K13_31 ) , .A( u0_R11_20 ) , .Z( u0_u12_X_31 ) );
  XOR2_X1 u0_u12_U26 (.B( u0_K13_30 ) , .A( u0_R11_21 ) , .Z( u0_u12_X_30 ) );
  XOR2_X1 u0_u12_U28 (.B( u0_K13_29 ) , .A( u0_R11_20 ) , .Z( u0_u12_X_29 ) );
  XOR2_X1 u0_u12_U29 (.B( u0_K13_28 ) , .A( u0_R11_19 ) , .Z( u0_u12_X_28 ) );
  XOR2_X1 u0_u12_U30 (.B( u0_K13_27 ) , .A( u0_R11_18 ) , .Z( u0_u12_X_27 ) );
  XOR2_X1 u0_u12_U31 (.B( u0_K13_26 ) , .A( u0_R11_17 ) , .Z( u0_u12_X_26 ) );
  XOR2_X1 u0_u12_U32 (.B( u0_K13_25 ) , .A( u0_R11_16 ) , .Z( u0_u12_X_25 ) );
  OAI22_X1 u0_u12_u4_U10 (.B2( u0_u12_u4_n135 ) , .ZN( u0_u12_u4_n137 ) , .B1( u0_u12_u4_n153 ) , .A1( u0_u12_u4_n155 ) , .A2( u0_u12_u4_n171 ) );
  AND3_X1 u0_u12_u4_U11 (.A2( u0_u12_u4_n134 ) , .ZN( u0_u12_u4_n135 ) , .A3( u0_u12_u4_n145 ) , .A1( u0_u12_u4_n157 ) );
  NAND2_X1 u0_u12_u4_U12 (.ZN( u0_u12_u4_n132 ) , .A2( u0_u12_u4_n170 ) , .A1( u0_u12_u4_n173 ) );
  AOI21_X1 u0_u12_u4_U13 (.B2( u0_u12_u4_n160 ) , .B1( u0_u12_u4_n161 ) , .ZN( u0_u12_u4_n162 ) , .A( u0_u12_u4_n170 ) );
  AOI21_X1 u0_u12_u4_U14 (.ZN( u0_u12_u4_n107 ) , .B2( u0_u12_u4_n143 ) , .A( u0_u12_u4_n174 ) , .B1( u0_u12_u4_n184 ) );
  AOI21_X1 u0_u12_u4_U15 (.B2( u0_u12_u4_n158 ) , .B1( u0_u12_u4_n159 ) , .ZN( u0_u12_u4_n163 ) , .A( u0_u12_u4_n174 ) );
  AOI21_X1 u0_u12_u4_U16 (.A( u0_u12_u4_n153 ) , .B2( u0_u12_u4_n154 ) , .B1( u0_u12_u4_n155 ) , .ZN( u0_u12_u4_n165 ) );
  AOI21_X1 u0_u12_u4_U17 (.A( u0_u12_u4_n156 ) , .B2( u0_u12_u4_n157 ) , .ZN( u0_u12_u4_n164 ) , .B1( u0_u12_u4_n184 ) );
  INV_X1 u0_u12_u4_U18 (.A( u0_u12_u4_n138 ) , .ZN( u0_u12_u4_n170 ) );
  AND2_X1 u0_u12_u4_U19 (.A2( u0_u12_u4_n120 ) , .ZN( u0_u12_u4_n155 ) , .A1( u0_u12_u4_n160 ) );
  INV_X1 u0_u12_u4_U20 (.A( u0_u12_u4_n156 ) , .ZN( u0_u12_u4_n175 ) );
  NAND2_X1 u0_u12_u4_U21 (.A2( u0_u12_u4_n118 ) , .ZN( u0_u12_u4_n131 ) , .A1( u0_u12_u4_n147 ) );
  NAND2_X1 u0_u12_u4_U22 (.A1( u0_u12_u4_n119 ) , .A2( u0_u12_u4_n120 ) , .ZN( u0_u12_u4_n130 ) );
  NAND2_X1 u0_u12_u4_U23 (.ZN( u0_u12_u4_n117 ) , .A2( u0_u12_u4_n118 ) , .A1( u0_u12_u4_n148 ) );
  NAND2_X1 u0_u12_u4_U24 (.ZN( u0_u12_u4_n129 ) , .A1( u0_u12_u4_n134 ) , .A2( u0_u12_u4_n148 ) );
  AND3_X1 u0_u12_u4_U25 (.A1( u0_u12_u4_n119 ) , .A2( u0_u12_u4_n143 ) , .A3( u0_u12_u4_n154 ) , .ZN( u0_u12_u4_n161 ) );
  AND2_X1 u0_u12_u4_U26 (.A1( u0_u12_u4_n145 ) , .A2( u0_u12_u4_n147 ) , .ZN( u0_u12_u4_n159 ) );
  OR3_X1 u0_u12_u4_U27 (.A3( u0_u12_u4_n114 ) , .A2( u0_u12_u4_n115 ) , .A1( u0_u12_u4_n116 ) , .ZN( u0_u12_u4_n136 ) );
  AOI21_X1 u0_u12_u4_U28 (.A( u0_u12_u4_n113 ) , .ZN( u0_u12_u4_n116 ) , .B2( u0_u12_u4_n173 ) , .B1( u0_u12_u4_n174 ) );
  AOI21_X1 u0_u12_u4_U29 (.ZN( u0_u12_u4_n115 ) , .B2( u0_u12_u4_n145 ) , .B1( u0_u12_u4_n146 ) , .A( u0_u12_u4_n156 ) );
  NOR2_X1 u0_u12_u4_U3 (.ZN( u0_u12_u4_n121 ) , .A1( u0_u12_u4_n181 ) , .A2( u0_u12_u4_n182 ) );
  OAI22_X1 u0_u12_u4_U30 (.ZN( u0_u12_u4_n114 ) , .A2( u0_u12_u4_n121 ) , .B1( u0_u12_u4_n160 ) , .B2( u0_u12_u4_n170 ) , .A1( u0_u12_u4_n171 ) );
  INV_X1 u0_u12_u4_U31 (.A( u0_u12_u4_n158 ) , .ZN( u0_u12_u4_n182 ) );
  INV_X1 u0_u12_u4_U32 (.ZN( u0_u12_u4_n181 ) , .A( u0_u12_u4_n96 ) );
  INV_X1 u0_u12_u4_U33 (.A( u0_u12_u4_n144 ) , .ZN( u0_u12_u4_n179 ) );
  INV_X1 u0_u12_u4_U34 (.A( u0_u12_u4_n157 ) , .ZN( u0_u12_u4_n178 ) );
  NAND2_X1 u0_u12_u4_U35 (.A2( u0_u12_u4_n154 ) , .A1( u0_u12_u4_n96 ) , .ZN( u0_u12_u4_n97 ) );
  INV_X1 u0_u12_u4_U36 (.ZN( u0_u12_u4_n186 ) , .A( u0_u12_u4_n95 ) );
  OAI221_X1 u0_u12_u4_U37 (.C1( u0_u12_u4_n134 ) , .B1( u0_u12_u4_n158 ) , .B2( u0_u12_u4_n171 ) , .C2( u0_u12_u4_n173 ) , .A( u0_u12_u4_n94 ) , .ZN( u0_u12_u4_n95 ) );
  AOI222_X1 u0_u12_u4_U38 (.B2( u0_u12_u4_n132 ) , .A1( u0_u12_u4_n138 ) , .C2( u0_u12_u4_n175 ) , .A2( u0_u12_u4_n179 ) , .C1( u0_u12_u4_n181 ) , .B1( u0_u12_u4_n185 ) , .ZN( u0_u12_u4_n94 ) );
  INV_X1 u0_u12_u4_U39 (.A( u0_u12_u4_n113 ) , .ZN( u0_u12_u4_n185 ) );
  INV_X1 u0_u12_u4_U4 (.A( u0_u12_u4_n117 ) , .ZN( u0_u12_u4_n184 ) );
  INV_X1 u0_u12_u4_U40 (.A( u0_u12_u4_n143 ) , .ZN( u0_u12_u4_n183 ) );
  NOR2_X1 u0_u12_u4_U41 (.ZN( u0_u12_u4_n138 ) , .A1( u0_u12_u4_n168 ) , .A2( u0_u12_u4_n169 ) );
  NOR2_X1 u0_u12_u4_U42 (.A1( u0_u12_u4_n150 ) , .A2( u0_u12_u4_n152 ) , .ZN( u0_u12_u4_n153 ) );
  NOR2_X1 u0_u12_u4_U43 (.A2( u0_u12_u4_n128 ) , .A1( u0_u12_u4_n138 ) , .ZN( u0_u12_u4_n156 ) );
  AOI22_X1 u0_u12_u4_U44 (.B2( u0_u12_u4_n122 ) , .A1( u0_u12_u4_n123 ) , .ZN( u0_u12_u4_n124 ) , .B1( u0_u12_u4_n128 ) , .A2( u0_u12_u4_n172 ) );
  INV_X1 u0_u12_u4_U45 (.A( u0_u12_u4_n153 ) , .ZN( u0_u12_u4_n172 ) );
  NAND2_X1 u0_u12_u4_U46 (.A2( u0_u12_u4_n120 ) , .ZN( u0_u12_u4_n123 ) , .A1( u0_u12_u4_n161 ) );
  AOI22_X1 u0_u12_u4_U47 (.B2( u0_u12_u4_n132 ) , .A2( u0_u12_u4_n133 ) , .ZN( u0_u12_u4_n140 ) , .A1( u0_u12_u4_n150 ) , .B1( u0_u12_u4_n179 ) );
  NAND2_X1 u0_u12_u4_U48 (.ZN( u0_u12_u4_n133 ) , .A2( u0_u12_u4_n146 ) , .A1( u0_u12_u4_n154 ) );
  NAND2_X1 u0_u12_u4_U49 (.A1( u0_u12_u4_n103 ) , .ZN( u0_u12_u4_n154 ) , .A2( u0_u12_u4_n98 ) );
  NOR4_X1 u0_u12_u4_U5 (.A4( u0_u12_u4_n106 ) , .A3( u0_u12_u4_n107 ) , .A2( u0_u12_u4_n108 ) , .A1( u0_u12_u4_n109 ) , .ZN( u0_u12_u4_n110 ) );
  NAND2_X1 u0_u12_u4_U50 (.A1( u0_u12_u4_n101 ) , .ZN( u0_u12_u4_n158 ) , .A2( u0_u12_u4_n99 ) );
  AOI21_X1 u0_u12_u4_U51 (.ZN( u0_u12_u4_n127 ) , .A( u0_u12_u4_n136 ) , .B2( u0_u12_u4_n150 ) , .B1( u0_u12_u4_n180 ) );
  INV_X1 u0_u12_u4_U52 (.A( u0_u12_u4_n160 ) , .ZN( u0_u12_u4_n180 ) );
  NAND2_X1 u0_u12_u4_U53 (.A2( u0_u12_u4_n104 ) , .A1( u0_u12_u4_n105 ) , .ZN( u0_u12_u4_n146 ) );
  NAND2_X1 u0_u12_u4_U54 (.A2( u0_u12_u4_n101 ) , .A1( u0_u12_u4_n102 ) , .ZN( u0_u12_u4_n160 ) );
  NAND2_X1 u0_u12_u4_U55 (.ZN( u0_u12_u4_n134 ) , .A1( u0_u12_u4_n98 ) , .A2( u0_u12_u4_n99 ) );
  NAND2_X1 u0_u12_u4_U56 (.A1( u0_u12_u4_n103 ) , .A2( u0_u12_u4_n104 ) , .ZN( u0_u12_u4_n143 ) );
  NAND2_X1 u0_u12_u4_U57 (.A2( u0_u12_u4_n105 ) , .ZN( u0_u12_u4_n145 ) , .A1( u0_u12_u4_n98 ) );
  NAND2_X1 u0_u12_u4_U58 (.A1( u0_u12_u4_n100 ) , .A2( u0_u12_u4_n105 ) , .ZN( u0_u12_u4_n120 ) );
  NAND2_X1 u0_u12_u4_U59 (.A1( u0_u12_u4_n102 ) , .A2( u0_u12_u4_n104 ) , .ZN( u0_u12_u4_n148 ) );
  AOI21_X1 u0_u12_u4_U6 (.ZN( u0_u12_u4_n106 ) , .B2( u0_u12_u4_n146 ) , .B1( u0_u12_u4_n158 ) , .A( u0_u12_u4_n170 ) );
  NAND2_X1 u0_u12_u4_U60 (.A2( u0_u12_u4_n100 ) , .A1( u0_u12_u4_n103 ) , .ZN( u0_u12_u4_n157 ) );
  INV_X1 u0_u12_u4_U61 (.A( u0_u12_u4_n150 ) , .ZN( u0_u12_u4_n173 ) );
  INV_X1 u0_u12_u4_U62 (.A( u0_u12_u4_n152 ) , .ZN( u0_u12_u4_n171 ) );
  NAND2_X1 u0_u12_u4_U63 (.A1( u0_u12_u4_n100 ) , .ZN( u0_u12_u4_n118 ) , .A2( u0_u12_u4_n99 ) );
  NAND2_X1 u0_u12_u4_U64 (.A2( u0_u12_u4_n100 ) , .A1( u0_u12_u4_n102 ) , .ZN( u0_u12_u4_n144 ) );
  NAND2_X1 u0_u12_u4_U65 (.A2( u0_u12_u4_n101 ) , .A1( u0_u12_u4_n105 ) , .ZN( u0_u12_u4_n96 ) );
  INV_X1 u0_u12_u4_U66 (.A( u0_u12_u4_n128 ) , .ZN( u0_u12_u4_n174 ) );
  NAND2_X1 u0_u12_u4_U67 (.A2( u0_u12_u4_n102 ) , .ZN( u0_u12_u4_n119 ) , .A1( u0_u12_u4_n98 ) );
  NAND2_X1 u0_u12_u4_U68 (.A2( u0_u12_u4_n101 ) , .A1( u0_u12_u4_n103 ) , .ZN( u0_u12_u4_n147 ) );
  NAND2_X1 u0_u12_u4_U69 (.A2( u0_u12_u4_n104 ) , .ZN( u0_u12_u4_n113 ) , .A1( u0_u12_u4_n99 ) );
  AOI21_X1 u0_u12_u4_U7 (.ZN( u0_u12_u4_n108 ) , .B2( u0_u12_u4_n134 ) , .B1( u0_u12_u4_n155 ) , .A( u0_u12_u4_n156 ) );
  NOR2_X1 u0_u12_u4_U70 (.A2( u0_u12_X_28 ) , .ZN( u0_u12_u4_n150 ) , .A1( u0_u12_u4_n168 ) );
  NOR2_X1 u0_u12_u4_U71 (.A2( u0_u12_X_29 ) , .ZN( u0_u12_u4_n152 ) , .A1( u0_u12_u4_n169 ) );
  NOR2_X1 u0_u12_u4_U72 (.A2( u0_u12_X_30 ) , .ZN( u0_u12_u4_n105 ) , .A1( u0_u12_u4_n176 ) );
  NOR2_X1 u0_u12_u4_U73 (.A2( u0_u12_X_26 ) , .ZN( u0_u12_u4_n100 ) , .A1( u0_u12_u4_n177 ) );
  NOR2_X1 u0_u12_u4_U74 (.A2( u0_u12_X_28 ) , .A1( u0_u12_X_29 ) , .ZN( u0_u12_u4_n128 ) );
  NOR2_X1 u0_u12_u4_U75 (.A2( u0_u12_X_27 ) , .A1( u0_u12_X_30 ) , .ZN( u0_u12_u4_n102 ) );
  NOR2_X1 u0_u12_u4_U76 (.A2( u0_u12_X_25 ) , .A1( u0_u12_X_26 ) , .ZN( u0_u12_u4_n98 ) );
  AND2_X1 u0_u12_u4_U77 (.A2( u0_u12_X_25 ) , .A1( u0_u12_X_26 ) , .ZN( u0_u12_u4_n104 ) );
  AND2_X1 u0_u12_u4_U78 (.A1( u0_u12_X_30 ) , .A2( u0_u12_u4_n176 ) , .ZN( u0_u12_u4_n99 ) );
  AND2_X1 u0_u12_u4_U79 (.A1( u0_u12_X_26 ) , .ZN( u0_u12_u4_n101 ) , .A2( u0_u12_u4_n177 ) );
  AOI21_X1 u0_u12_u4_U8 (.ZN( u0_u12_u4_n109 ) , .A( u0_u12_u4_n153 ) , .B1( u0_u12_u4_n159 ) , .B2( u0_u12_u4_n184 ) );
  AND2_X1 u0_u12_u4_U80 (.A1( u0_u12_X_27 ) , .A2( u0_u12_X_30 ) , .ZN( u0_u12_u4_n103 ) );
  INV_X1 u0_u12_u4_U81 (.A( u0_u12_X_28 ) , .ZN( u0_u12_u4_n169 ) );
  INV_X1 u0_u12_u4_U82 (.A( u0_u12_X_29 ) , .ZN( u0_u12_u4_n168 ) );
  INV_X1 u0_u12_u4_U83 (.A( u0_u12_X_25 ) , .ZN( u0_u12_u4_n177 ) );
  INV_X1 u0_u12_u4_U84 (.A( u0_u12_X_27 ) , .ZN( u0_u12_u4_n176 ) );
  NAND4_X1 u0_u12_u4_U85 (.ZN( u0_out12_25 ) , .A4( u0_u12_u4_n139 ) , .A3( u0_u12_u4_n140 ) , .A2( u0_u12_u4_n141 ) , .A1( u0_u12_u4_n142 ) );
  OAI21_X1 u0_u12_u4_U86 (.A( u0_u12_u4_n128 ) , .B2( u0_u12_u4_n129 ) , .B1( u0_u12_u4_n130 ) , .ZN( u0_u12_u4_n142 ) );
  OAI21_X1 u0_u12_u4_U87 (.B2( u0_u12_u4_n131 ) , .ZN( u0_u12_u4_n141 ) , .A( u0_u12_u4_n175 ) , .B1( u0_u12_u4_n183 ) );
  NAND4_X1 u0_u12_u4_U88 (.ZN( u0_out12_14 ) , .A4( u0_u12_u4_n124 ) , .A3( u0_u12_u4_n125 ) , .A2( u0_u12_u4_n126 ) , .A1( u0_u12_u4_n127 ) );
  AOI22_X1 u0_u12_u4_U89 (.B2( u0_u12_u4_n117 ) , .ZN( u0_u12_u4_n126 ) , .A1( u0_u12_u4_n129 ) , .B1( u0_u12_u4_n152 ) , .A2( u0_u12_u4_n175 ) );
  AOI211_X1 u0_u12_u4_U9 (.B( u0_u12_u4_n136 ) , .A( u0_u12_u4_n137 ) , .C2( u0_u12_u4_n138 ) , .ZN( u0_u12_u4_n139 ) , .C1( u0_u12_u4_n182 ) );
  AOI22_X1 u0_u12_u4_U90 (.ZN( u0_u12_u4_n125 ) , .B2( u0_u12_u4_n131 ) , .A2( u0_u12_u4_n132 ) , .B1( u0_u12_u4_n138 ) , .A1( u0_u12_u4_n178 ) );
  NAND4_X1 u0_u12_u4_U91 (.ZN( u0_out12_8 ) , .A4( u0_u12_u4_n110 ) , .A3( u0_u12_u4_n111 ) , .A2( u0_u12_u4_n112 ) , .A1( u0_u12_u4_n186 ) );
  NAND2_X1 u0_u12_u4_U92 (.ZN( u0_u12_u4_n112 ) , .A2( u0_u12_u4_n130 ) , .A1( u0_u12_u4_n150 ) );
  AOI22_X1 u0_u12_u4_U93 (.ZN( u0_u12_u4_n111 ) , .B2( u0_u12_u4_n132 ) , .A1( u0_u12_u4_n152 ) , .B1( u0_u12_u4_n178 ) , .A2( u0_u12_u4_n97 ) );
  AOI22_X1 u0_u12_u4_U94 (.B2( u0_u12_u4_n149 ) , .B1( u0_u12_u4_n150 ) , .A2( u0_u12_u4_n151 ) , .A1( u0_u12_u4_n152 ) , .ZN( u0_u12_u4_n167 ) );
  NOR4_X1 u0_u12_u4_U95 (.A4( u0_u12_u4_n162 ) , .A3( u0_u12_u4_n163 ) , .A2( u0_u12_u4_n164 ) , .A1( u0_u12_u4_n165 ) , .ZN( u0_u12_u4_n166 ) );
  NAND3_X1 u0_u12_u4_U96 (.ZN( u0_out12_3 ) , .A3( u0_u12_u4_n166 ) , .A1( u0_u12_u4_n167 ) , .A2( u0_u12_u4_n186 ) );
  NAND3_X1 u0_u12_u4_U97 (.A3( u0_u12_u4_n146 ) , .A2( u0_u12_u4_n147 ) , .A1( u0_u12_u4_n148 ) , .ZN( u0_u12_u4_n149 ) );
  NAND3_X1 u0_u12_u4_U98 (.A3( u0_u12_u4_n143 ) , .A2( u0_u12_u4_n144 ) , .A1( u0_u12_u4_n145 ) , .ZN( u0_u12_u4_n151 ) );
  NAND3_X1 u0_u12_u4_U99 (.A3( u0_u12_u4_n121 ) , .ZN( u0_u12_u4_n122 ) , .A2( u0_u12_u4_n144 ) , .A1( u0_u12_u4_n154 ) );
  INV_X1 u0_u12_u5_U10 (.A( u0_u12_u5_n121 ) , .ZN( u0_u12_u5_n177 ) );
  NOR3_X1 u0_u12_u5_U100 (.A3( u0_u12_u5_n141 ) , .A1( u0_u12_u5_n142 ) , .ZN( u0_u12_u5_n143 ) , .A2( u0_u12_u5_n191 ) );
  NAND4_X1 u0_u12_u5_U101 (.ZN( u0_out12_4 ) , .A4( u0_u12_u5_n112 ) , .A2( u0_u12_u5_n113 ) , .A1( u0_u12_u5_n114 ) , .A3( u0_u12_u5_n195 ) );
  AOI211_X1 u0_u12_u5_U102 (.A( u0_u12_u5_n110 ) , .C1( u0_u12_u5_n111 ) , .ZN( u0_u12_u5_n112 ) , .B( u0_u12_u5_n118 ) , .C2( u0_u12_u5_n177 ) );
  AOI222_X1 u0_u12_u5_U103 (.ZN( u0_u12_u5_n113 ) , .A1( u0_u12_u5_n131 ) , .C1( u0_u12_u5_n148 ) , .B2( u0_u12_u5_n174 ) , .C2( u0_u12_u5_n178 ) , .A2( u0_u12_u5_n179 ) , .B1( u0_u12_u5_n99 ) );
  NAND3_X1 u0_u12_u5_U104 (.A2( u0_u12_u5_n154 ) , .A3( u0_u12_u5_n158 ) , .A1( u0_u12_u5_n161 ) , .ZN( u0_u12_u5_n99 ) );
  NOR2_X1 u0_u12_u5_U11 (.ZN( u0_u12_u5_n160 ) , .A2( u0_u12_u5_n173 ) , .A1( u0_u12_u5_n177 ) );
  INV_X1 u0_u12_u5_U12 (.A( u0_u12_u5_n150 ) , .ZN( u0_u12_u5_n174 ) );
  AOI21_X1 u0_u12_u5_U13 (.A( u0_u12_u5_n160 ) , .B2( u0_u12_u5_n161 ) , .ZN( u0_u12_u5_n162 ) , .B1( u0_u12_u5_n192 ) );
  INV_X1 u0_u12_u5_U14 (.A( u0_u12_u5_n159 ) , .ZN( u0_u12_u5_n192 ) );
  AOI21_X1 u0_u12_u5_U15 (.A( u0_u12_u5_n156 ) , .B2( u0_u12_u5_n157 ) , .B1( u0_u12_u5_n158 ) , .ZN( u0_u12_u5_n163 ) );
  AOI21_X1 u0_u12_u5_U16 (.B2( u0_u12_u5_n139 ) , .B1( u0_u12_u5_n140 ) , .ZN( u0_u12_u5_n141 ) , .A( u0_u12_u5_n150 ) );
  OAI21_X1 u0_u12_u5_U17 (.A( u0_u12_u5_n133 ) , .B2( u0_u12_u5_n134 ) , .B1( u0_u12_u5_n135 ) , .ZN( u0_u12_u5_n142 ) );
  OAI21_X1 u0_u12_u5_U18 (.ZN( u0_u12_u5_n133 ) , .B2( u0_u12_u5_n147 ) , .A( u0_u12_u5_n173 ) , .B1( u0_u12_u5_n188 ) );
  NAND2_X1 u0_u12_u5_U19 (.A2( u0_u12_u5_n119 ) , .A1( u0_u12_u5_n123 ) , .ZN( u0_u12_u5_n137 ) );
  INV_X1 u0_u12_u5_U20 (.A( u0_u12_u5_n155 ) , .ZN( u0_u12_u5_n194 ) );
  NAND2_X1 u0_u12_u5_U21 (.A1( u0_u12_u5_n121 ) , .ZN( u0_u12_u5_n132 ) , .A2( u0_u12_u5_n172 ) );
  NAND2_X1 u0_u12_u5_U22 (.A2( u0_u12_u5_n122 ) , .ZN( u0_u12_u5_n136 ) , .A1( u0_u12_u5_n154 ) );
  NAND2_X1 u0_u12_u5_U23 (.A2( u0_u12_u5_n119 ) , .A1( u0_u12_u5_n120 ) , .ZN( u0_u12_u5_n159 ) );
  INV_X1 u0_u12_u5_U24 (.A( u0_u12_u5_n156 ) , .ZN( u0_u12_u5_n175 ) );
  INV_X1 u0_u12_u5_U25 (.A( u0_u12_u5_n158 ) , .ZN( u0_u12_u5_n188 ) );
  INV_X1 u0_u12_u5_U26 (.A( u0_u12_u5_n152 ) , .ZN( u0_u12_u5_n179 ) );
  INV_X1 u0_u12_u5_U27 (.A( u0_u12_u5_n140 ) , .ZN( u0_u12_u5_n182 ) );
  INV_X1 u0_u12_u5_U28 (.A( u0_u12_u5_n151 ) , .ZN( u0_u12_u5_n183 ) );
  INV_X1 u0_u12_u5_U29 (.A( u0_u12_u5_n123 ) , .ZN( u0_u12_u5_n185 ) );
  NOR2_X1 u0_u12_u5_U3 (.ZN( u0_u12_u5_n134 ) , .A1( u0_u12_u5_n183 ) , .A2( u0_u12_u5_n190 ) );
  INV_X1 u0_u12_u5_U30 (.A( u0_u12_u5_n161 ) , .ZN( u0_u12_u5_n184 ) );
  INV_X1 u0_u12_u5_U31 (.A( u0_u12_u5_n139 ) , .ZN( u0_u12_u5_n189 ) );
  INV_X1 u0_u12_u5_U32 (.A( u0_u12_u5_n157 ) , .ZN( u0_u12_u5_n190 ) );
  INV_X1 u0_u12_u5_U33 (.A( u0_u12_u5_n120 ) , .ZN( u0_u12_u5_n193 ) );
  NAND2_X1 u0_u12_u5_U34 (.ZN( u0_u12_u5_n111 ) , .A1( u0_u12_u5_n140 ) , .A2( u0_u12_u5_n155 ) );
  NOR2_X1 u0_u12_u5_U35 (.ZN( u0_u12_u5_n100 ) , .A1( u0_u12_u5_n170 ) , .A2( u0_u12_u5_n180 ) );
  INV_X1 u0_u12_u5_U36 (.A( u0_u12_u5_n117 ) , .ZN( u0_u12_u5_n196 ) );
  OAI221_X1 u0_u12_u5_U37 (.A( u0_u12_u5_n116 ) , .ZN( u0_u12_u5_n117 ) , .B2( u0_u12_u5_n119 ) , .C1( u0_u12_u5_n153 ) , .C2( u0_u12_u5_n158 ) , .B1( u0_u12_u5_n172 ) );
  AOI222_X1 u0_u12_u5_U38 (.ZN( u0_u12_u5_n116 ) , .B2( u0_u12_u5_n145 ) , .C1( u0_u12_u5_n148 ) , .A2( u0_u12_u5_n174 ) , .C2( u0_u12_u5_n177 ) , .B1( u0_u12_u5_n187 ) , .A1( u0_u12_u5_n193 ) );
  INV_X1 u0_u12_u5_U39 (.A( u0_u12_u5_n115 ) , .ZN( u0_u12_u5_n187 ) );
  INV_X1 u0_u12_u5_U4 (.A( u0_u12_u5_n138 ) , .ZN( u0_u12_u5_n191 ) );
  AOI22_X1 u0_u12_u5_U40 (.B2( u0_u12_u5_n131 ) , .A2( u0_u12_u5_n146 ) , .ZN( u0_u12_u5_n169 ) , .B1( u0_u12_u5_n174 ) , .A1( u0_u12_u5_n185 ) );
  NOR2_X1 u0_u12_u5_U41 (.A1( u0_u12_u5_n146 ) , .ZN( u0_u12_u5_n150 ) , .A2( u0_u12_u5_n173 ) );
  AOI21_X1 u0_u12_u5_U42 (.A( u0_u12_u5_n118 ) , .B2( u0_u12_u5_n145 ) , .ZN( u0_u12_u5_n168 ) , .B1( u0_u12_u5_n186 ) );
  INV_X1 u0_u12_u5_U43 (.A( u0_u12_u5_n122 ) , .ZN( u0_u12_u5_n186 ) );
  NOR2_X1 u0_u12_u5_U44 (.A1( u0_u12_u5_n146 ) , .ZN( u0_u12_u5_n152 ) , .A2( u0_u12_u5_n176 ) );
  NOR2_X1 u0_u12_u5_U45 (.A1( u0_u12_u5_n115 ) , .ZN( u0_u12_u5_n118 ) , .A2( u0_u12_u5_n153 ) );
  NOR2_X1 u0_u12_u5_U46 (.A2( u0_u12_u5_n145 ) , .ZN( u0_u12_u5_n156 ) , .A1( u0_u12_u5_n174 ) );
  NOR2_X1 u0_u12_u5_U47 (.ZN( u0_u12_u5_n121 ) , .A2( u0_u12_u5_n145 ) , .A1( u0_u12_u5_n176 ) );
  AOI22_X1 u0_u12_u5_U48 (.ZN( u0_u12_u5_n114 ) , .A2( u0_u12_u5_n137 ) , .A1( u0_u12_u5_n145 ) , .B2( u0_u12_u5_n175 ) , .B1( u0_u12_u5_n193 ) );
  OAI211_X1 u0_u12_u5_U49 (.B( u0_u12_u5_n124 ) , .A( u0_u12_u5_n125 ) , .C2( u0_u12_u5_n126 ) , .C1( u0_u12_u5_n127 ) , .ZN( u0_u12_u5_n128 ) );
  OAI21_X1 u0_u12_u5_U5 (.B2( u0_u12_u5_n136 ) , .B1( u0_u12_u5_n137 ) , .ZN( u0_u12_u5_n138 ) , .A( u0_u12_u5_n177 ) );
  NOR3_X1 u0_u12_u5_U50 (.ZN( u0_u12_u5_n127 ) , .A1( u0_u12_u5_n136 ) , .A3( u0_u12_u5_n148 ) , .A2( u0_u12_u5_n182 ) );
  OAI21_X1 u0_u12_u5_U51 (.ZN( u0_u12_u5_n124 ) , .A( u0_u12_u5_n177 ) , .B2( u0_u12_u5_n183 ) , .B1( u0_u12_u5_n189 ) );
  OAI21_X1 u0_u12_u5_U52 (.ZN( u0_u12_u5_n125 ) , .A( u0_u12_u5_n174 ) , .B2( u0_u12_u5_n185 ) , .B1( u0_u12_u5_n190 ) );
  AOI21_X1 u0_u12_u5_U53 (.A( u0_u12_u5_n153 ) , .B2( u0_u12_u5_n154 ) , .B1( u0_u12_u5_n155 ) , .ZN( u0_u12_u5_n164 ) );
  AOI21_X1 u0_u12_u5_U54 (.ZN( u0_u12_u5_n110 ) , .B1( u0_u12_u5_n122 ) , .B2( u0_u12_u5_n139 ) , .A( u0_u12_u5_n153 ) );
  INV_X1 u0_u12_u5_U55 (.A( u0_u12_u5_n153 ) , .ZN( u0_u12_u5_n176 ) );
  INV_X1 u0_u12_u5_U56 (.A( u0_u12_u5_n126 ) , .ZN( u0_u12_u5_n173 ) );
  AND2_X1 u0_u12_u5_U57 (.A2( u0_u12_u5_n104 ) , .A1( u0_u12_u5_n107 ) , .ZN( u0_u12_u5_n147 ) );
  AND2_X1 u0_u12_u5_U58 (.A2( u0_u12_u5_n104 ) , .A1( u0_u12_u5_n108 ) , .ZN( u0_u12_u5_n148 ) );
  NAND2_X1 u0_u12_u5_U59 (.A1( u0_u12_u5_n105 ) , .A2( u0_u12_u5_n106 ) , .ZN( u0_u12_u5_n158 ) );
  INV_X1 u0_u12_u5_U6 (.A( u0_u12_u5_n135 ) , .ZN( u0_u12_u5_n178 ) );
  NAND2_X1 u0_u12_u5_U60 (.A2( u0_u12_u5_n108 ) , .A1( u0_u12_u5_n109 ) , .ZN( u0_u12_u5_n139 ) );
  NAND2_X1 u0_u12_u5_U61 (.A1( u0_u12_u5_n106 ) , .A2( u0_u12_u5_n108 ) , .ZN( u0_u12_u5_n119 ) );
  NAND2_X1 u0_u12_u5_U62 (.A2( u0_u12_u5_n103 ) , .A1( u0_u12_u5_n105 ) , .ZN( u0_u12_u5_n140 ) );
  NAND2_X1 u0_u12_u5_U63 (.A2( u0_u12_u5_n104 ) , .A1( u0_u12_u5_n105 ) , .ZN( u0_u12_u5_n155 ) );
  NAND2_X1 u0_u12_u5_U64 (.A2( u0_u12_u5_n106 ) , .A1( u0_u12_u5_n107 ) , .ZN( u0_u12_u5_n122 ) );
  NAND2_X1 u0_u12_u5_U65 (.A2( u0_u12_u5_n100 ) , .A1( u0_u12_u5_n106 ) , .ZN( u0_u12_u5_n115 ) );
  NAND2_X1 u0_u12_u5_U66 (.A2( u0_u12_u5_n100 ) , .A1( u0_u12_u5_n103 ) , .ZN( u0_u12_u5_n161 ) );
  NAND2_X1 u0_u12_u5_U67 (.A1( u0_u12_u5_n105 ) , .A2( u0_u12_u5_n109 ) , .ZN( u0_u12_u5_n154 ) );
  INV_X1 u0_u12_u5_U68 (.A( u0_u12_u5_n146 ) , .ZN( u0_u12_u5_n172 ) );
  NAND2_X1 u0_u12_u5_U69 (.A1( u0_u12_u5_n103 ) , .A2( u0_u12_u5_n108 ) , .ZN( u0_u12_u5_n123 ) );
  OAI22_X1 u0_u12_u5_U7 (.B2( u0_u12_u5_n149 ) , .B1( u0_u12_u5_n150 ) , .A2( u0_u12_u5_n151 ) , .A1( u0_u12_u5_n152 ) , .ZN( u0_u12_u5_n165 ) );
  NAND2_X1 u0_u12_u5_U70 (.A2( u0_u12_u5_n103 ) , .A1( u0_u12_u5_n107 ) , .ZN( u0_u12_u5_n151 ) );
  NAND2_X1 u0_u12_u5_U71 (.A2( u0_u12_u5_n107 ) , .A1( u0_u12_u5_n109 ) , .ZN( u0_u12_u5_n120 ) );
  NAND2_X1 u0_u12_u5_U72 (.A2( u0_u12_u5_n100 ) , .A1( u0_u12_u5_n109 ) , .ZN( u0_u12_u5_n157 ) );
  AND2_X1 u0_u12_u5_U73 (.A2( u0_u12_u5_n100 ) , .A1( u0_u12_u5_n104 ) , .ZN( u0_u12_u5_n131 ) );
  INV_X1 u0_u12_u5_U74 (.A( u0_u12_u5_n102 ) , .ZN( u0_u12_u5_n195 ) );
  OAI221_X1 u0_u12_u5_U75 (.A( u0_u12_u5_n101 ) , .ZN( u0_u12_u5_n102 ) , .C2( u0_u12_u5_n115 ) , .C1( u0_u12_u5_n126 ) , .B1( u0_u12_u5_n134 ) , .B2( u0_u12_u5_n160 ) );
  OAI21_X1 u0_u12_u5_U76 (.ZN( u0_u12_u5_n101 ) , .B1( u0_u12_u5_n137 ) , .A( u0_u12_u5_n146 ) , .B2( u0_u12_u5_n147 ) );
  NOR2_X1 u0_u12_u5_U77 (.A2( u0_u12_X_34 ) , .A1( u0_u12_X_35 ) , .ZN( u0_u12_u5_n145 ) );
  NOR2_X1 u0_u12_u5_U78 (.A2( u0_u12_X_34 ) , .ZN( u0_u12_u5_n146 ) , .A1( u0_u12_u5_n171 ) );
  NOR2_X1 u0_u12_u5_U79 (.A2( u0_u12_X_31 ) , .A1( u0_u12_X_32 ) , .ZN( u0_u12_u5_n103 ) );
  NOR3_X1 u0_u12_u5_U8 (.A2( u0_u12_u5_n147 ) , .A1( u0_u12_u5_n148 ) , .ZN( u0_u12_u5_n149 ) , .A3( u0_u12_u5_n194 ) );
  NOR2_X1 u0_u12_u5_U80 (.A2( u0_u12_X_36 ) , .ZN( u0_u12_u5_n105 ) , .A1( u0_u12_u5_n180 ) );
  NOR2_X1 u0_u12_u5_U81 (.A2( u0_u12_X_33 ) , .ZN( u0_u12_u5_n108 ) , .A1( u0_u12_u5_n170 ) );
  NOR2_X1 u0_u12_u5_U82 (.A2( u0_u12_X_33 ) , .A1( u0_u12_X_36 ) , .ZN( u0_u12_u5_n107 ) );
  NOR2_X1 u0_u12_u5_U83 (.A2( u0_u12_X_31 ) , .ZN( u0_u12_u5_n104 ) , .A1( u0_u12_u5_n181 ) );
  NAND2_X1 u0_u12_u5_U84 (.A2( u0_u12_X_34 ) , .A1( u0_u12_X_35 ) , .ZN( u0_u12_u5_n153 ) );
  NAND2_X1 u0_u12_u5_U85 (.A1( u0_u12_X_34 ) , .ZN( u0_u12_u5_n126 ) , .A2( u0_u12_u5_n171 ) );
  AND2_X1 u0_u12_u5_U86 (.A1( u0_u12_X_31 ) , .A2( u0_u12_X_32 ) , .ZN( u0_u12_u5_n106 ) );
  AND2_X1 u0_u12_u5_U87 (.A1( u0_u12_X_31 ) , .ZN( u0_u12_u5_n109 ) , .A2( u0_u12_u5_n181 ) );
  INV_X1 u0_u12_u5_U88 (.A( u0_u12_X_33 ) , .ZN( u0_u12_u5_n180 ) );
  INV_X1 u0_u12_u5_U89 (.A( u0_u12_X_35 ) , .ZN( u0_u12_u5_n171 ) );
  NOR2_X1 u0_u12_u5_U9 (.ZN( u0_u12_u5_n135 ) , .A1( u0_u12_u5_n173 ) , .A2( u0_u12_u5_n176 ) );
  INV_X1 u0_u12_u5_U90 (.A( u0_u12_X_36 ) , .ZN( u0_u12_u5_n170 ) );
  INV_X1 u0_u12_u5_U91 (.A( u0_u12_X_32 ) , .ZN( u0_u12_u5_n181 ) );
  NAND4_X1 u0_u12_u5_U92 (.ZN( u0_out12_29 ) , .A4( u0_u12_u5_n129 ) , .A3( u0_u12_u5_n130 ) , .A2( u0_u12_u5_n168 ) , .A1( u0_u12_u5_n196 ) );
  AOI221_X1 u0_u12_u5_U93 (.A( u0_u12_u5_n128 ) , .ZN( u0_u12_u5_n129 ) , .C2( u0_u12_u5_n132 ) , .B2( u0_u12_u5_n159 ) , .B1( u0_u12_u5_n176 ) , .C1( u0_u12_u5_n184 ) );
  AOI222_X1 u0_u12_u5_U94 (.ZN( u0_u12_u5_n130 ) , .A2( u0_u12_u5_n146 ) , .B1( u0_u12_u5_n147 ) , .C2( u0_u12_u5_n175 ) , .B2( u0_u12_u5_n179 ) , .A1( u0_u12_u5_n188 ) , .C1( u0_u12_u5_n194 ) );
  NAND4_X1 u0_u12_u5_U95 (.ZN( u0_out12_19 ) , .A4( u0_u12_u5_n166 ) , .A3( u0_u12_u5_n167 ) , .A2( u0_u12_u5_n168 ) , .A1( u0_u12_u5_n169 ) );
  AOI22_X1 u0_u12_u5_U96 (.B2( u0_u12_u5_n145 ) , .A2( u0_u12_u5_n146 ) , .ZN( u0_u12_u5_n167 ) , .B1( u0_u12_u5_n182 ) , .A1( u0_u12_u5_n189 ) );
  NOR4_X1 u0_u12_u5_U97 (.A4( u0_u12_u5_n162 ) , .A3( u0_u12_u5_n163 ) , .A2( u0_u12_u5_n164 ) , .A1( u0_u12_u5_n165 ) , .ZN( u0_u12_u5_n166 ) );
  NAND4_X1 u0_u12_u5_U98 (.ZN( u0_out12_11 ) , .A4( u0_u12_u5_n143 ) , .A3( u0_u12_u5_n144 ) , .A2( u0_u12_u5_n169 ) , .A1( u0_u12_u5_n196 ) );
  AOI22_X1 u0_u12_u5_U99 (.A2( u0_u12_u5_n132 ) , .ZN( u0_u12_u5_n144 ) , .B2( u0_u12_u5_n145 ) , .B1( u0_u12_u5_n184 ) , .A1( u0_u12_u5_n194 ) );
  AOI22_X1 u0_u12_u6_U10 (.A2( u0_u12_u6_n151 ) , .B2( u0_u12_u6_n161 ) , .A1( u0_u12_u6_n167 ) , .B1( u0_u12_u6_n170 ) , .ZN( u0_u12_u6_n89 ) );
  AOI21_X1 u0_u12_u6_U11 (.B1( u0_u12_u6_n107 ) , .B2( u0_u12_u6_n132 ) , .A( u0_u12_u6_n158 ) , .ZN( u0_u12_u6_n88 ) );
  AOI21_X1 u0_u12_u6_U12 (.B2( u0_u12_u6_n147 ) , .B1( u0_u12_u6_n148 ) , .ZN( u0_u12_u6_n149 ) , .A( u0_u12_u6_n158 ) );
  AOI21_X1 u0_u12_u6_U13 (.ZN( u0_u12_u6_n106 ) , .A( u0_u12_u6_n142 ) , .B2( u0_u12_u6_n159 ) , .B1( u0_u12_u6_n164 ) );
  INV_X1 u0_u12_u6_U14 (.A( u0_u12_u6_n155 ) , .ZN( u0_u12_u6_n161 ) );
  INV_X1 u0_u12_u6_U15 (.A( u0_u12_u6_n128 ) , .ZN( u0_u12_u6_n164 ) );
  NAND2_X1 u0_u12_u6_U16 (.ZN( u0_u12_u6_n110 ) , .A1( u0_u12_u6_n122 ) , .A2( u0_u12_u6_n129 ) );
  NAND2_X1 u0_u12_u6_U17 (.ZN( u0_u12_u6_n124 ) , .A2( u0_u12_u6_n146 ) , .A1( u0_u12_u6_n148 ) );
  INV_X1 u0_u12_u6_U18 (.A( u0_u12_u6_n132 ) , .ZN( u0_u12_u6_n171 ) );
  AND2_X1 u0_u12_u6_U19 (.A1( u0_u12_u6_n100 ) , .ZN( u0_u12_u6_n130 ) , .A2( u0_u12_u6_n147 ) );
  INV_X1 u0_u12_u6_U20 (.A( u0_u12_u6_n127 ) , .ZN( u0_u12_u6_n173 ) );
  INV_X1 u0_u12_u6_U21 (.A( u0_u12_u6_n121 ) , .ZN( u0_u12_u6_n167 ) );
  INV_X1 u0_u12_u6_U22 (.A( u0_u12_u6_n100 ) , .ZN( u0_u12_u6_n169 ) );
  INV_X1 u0_u12_u6_U23 (.A( u0_u12_u6_n123 ) , .ZN( u0_u12_u6_n170 ) );
  INV_X1 u0_u12_u6_U24 (.A( u0_u12_u6_n113 ) , .ZN( u0_u12_u6_n168 ) );
  AND2_X1 u0_u12_u6_U25 (.A1( u0_u12_u6_n107 ) , .A2( u0_u12_u6_n119 ) , .ZN( u0_u12_u6_n133 ) );
  AND2_X1 u0_u12_u6_U26 (.A2( u0_u12_u6_n121 ) , .A1( u0_u12_u6_n122 ) , .ZN( u0_u12_u6_n131 ) );
  AND3_X1 u0_u12_u6_U27 (.ZN( u0_u12_u6_n120 ) , .A2( u0_u12_u6_n127 ) , .A1( u0_u12_u6_n132 ) , .A3( u0_u12_u6_n145 ) );
  INV_X1 u0_u12_u6_U28 (.A( u0_u12_u6_n146 ) , .ZN( u0_u12_u6_n163 ) );
  AOI222_X1 u0_u12_u6_U29 (.ZN( u0_u12_u6_n114 ) , .A1( u0_u12_u6_n118 ) , .A2( u0_u12_u6_n126 ) , .B2( u0_u12_u6_n151 ) , .C2( u0_u12_u6_n159 ) , .C1( u0_u12_u6_n168 ) , .B1( u0_u12_u6_n169 ) );
  INV_X1 u0_u12_u6_U3 (.A( u0_u12_u6_n110 ) , .ZN( u0_u12_u6_n166 ) );
  NOR2_X1 u0_u12_u6_U30 (.A1( u0_u12_u6_n162 ) , .A2( u0_u12_u6_n165 ) , .ZN( u0_u12_u6_n98 ) );
  AOI211_X1 u0_u12_u6_U31 (.B( u0_u12_u6_n134 ) , .A( u0_u12_u6_n135 ) , .C1( u0_u12_u6_n136 ) , .ZN( u0_u12_u6_n137 ) , .C2( u0_u12_u6_n151 ) );
  AOI21_X1 u0_u12_u6_U32 (.B2( u0_u12_u6_n132 ) , .B1( u0_u12_u6_n133 ) , .ZN( u0_u12_u6_n134 ) , .A( u0_u12_u6_n158 ) );
  AOI21_X1 u0_u12_u6_U33 (.B1( u0_u12_u6_n131 ) , .ZN( u0_u12_u6_n135 ) , .A( u0_u12_u6_n144 ) , .B2( u0_u12_u6_n146 ) );
  NAND4_X1 u0_u12_u6_U34 (.A4( u0_u12_u6_n127 ) , .A3( u0_u12_u6_n128 ) , .A2( u0_u12_u6_n129 ) , .A1( u0_u12_u6_n130 ) , .ZN( u0_u12_u6_n136 ) );
  NAND2_X1 u0_u12_u6_U35 (.A1( u0_u12_u6_n144 ) , .ZN( u0_u12_u6_n151 ) , .A2( u0_u12_u6_n158 ) );
  NAND2_X1 u0_u12_u6_U36 (.ZN( u0_u12_u6_n132 ) , .A1( u0_u12_u6_n91 ) , .A2( u0_u12_u6_n97 ) );
  AOI22_X1 u0_u12_u6_U37 (.B2( u0_u12_u6_n110 ) , .B1( u0_u12_u6_n111 ) , .A1( u0_u12_u6_n112 ) , .ZN( u0_u12_u6_n115 ) , .A2( u0_u12_u6_n161 ) );
  NAND4_X1 u0_u12_u6_U38 (.A3( u0_u12_u6_n109 ) , .ZN( u0_u12_u6_n112 ) , .A4( u0_u12_u6_n132 ) , .A2( u0_u12_u6_n147 ) , .A1( u0_u12_u6_n166 ) );
  NOR2_X1 u0_u12_u6_U39 (.ZN( u0_u12_u6_n109 ) , .A1( u0_u12_u6_n170 ) , .A2( u0_u12_u6_n173 ) );
  INV_X1 u0_u12_u6_U4 (.A( u0_u12_u6_n142 ) , .ZN( u0_u12_u6_n174 ) );
  NOR2_X1 u0_u12_u6_U40 (.A2( u0_u12_u6_n126 ) , .ZN( u0_u12_u6_n155 ) , .A1( u0_u12_u6_n160 ) );
  NAND2_X1 u0_u12_u6_U41 (.ZN( u0_u12_u6_n146 ) , .A2( u0_u12_u6_n94 ) , .A1( u0_u12_u6_n99 ) );
  AOI21_X1 u0_u12_u6_U42 (.A( u0_u12_u6_n144 ) , .B2( u0_u12_u6_n145 ) , .B1( u0_u12_u6_n146 ) , .ZN( u0_u12_u6_n150 ) );
  INV_X1 u0_u12_u6_U43 (.A( u0_u12_u6_n111 ) , .ZN( u0_u12_u6_n158 ) );
  NAND2_X1 u0_u12_u6_U44 (.ZN( u0_u12_u6_n127 ) , .A1( u0_u12_u6_n91 ) , .A2( u0_u12_u6_n92 ) );
  NAND2_X1 u0_u12_u6_U45 (.ZN( u0_u12_u6_n129 ) , .A2( u0_u12_u6_n95 ) , .A1( u0_u12_u6_n96 ) );
  INV_X1 u0_u12_u6_U46 (.A( u0_u12_u6_n144 ) , .ZN( u0_u12_u6_n159 ) );
  NAND2_X1 u0_u12_u6_U47 (.ZN( u0_u12_u6_n145 ) , .A2( u0_u12_u6_n97 ) , .A1( u0_u12_u6_n98 ) );
  NAND2_X1 u0_u12_u6_U48 (.ZN( u0_u12_u6_n148 ) , .A2( u0_u12_u6_n92 ) , .A1( u0_u12_u6_n94 ) );
  NAND2_X1 u0_u12_u6_U49 (.ZN( u0_u12_u6_n108 ) , .A2( u0_u12_u6_n139 ) , .A1( u0_u12_u6_n144 ) );
  NAND2_X1 u0_u12_u6_U5 (.A2( u0_u12_u6_n143 ) , .ZN( u0_u12_u6_n152 ) , .A1( u0_u12_u6_n166 ) );
  NAND2_X1 u0_u12_u6_U50 (.ZN( u0_u12_u6_n121 ) , .A2( u0_u12_u6_n95 ) , .A1( u0_u12_u6_n97 ) );
  NAND2_X1 u0_u12_u6_U51 (.ZN( u0_u12_u6_n107 ) , .A2( u0_u12_u6_n92 ) , .A1( u0_u12_u6_n95 ) );
  AND2_X1 u0_u12_u6_U52 (.ZN( u0_u12_u6_n118 ) , .A2( u0_u12_u6_n91 ) , .A1( u0_u12_u6_n99 ) );
  NAND2_X1 u0_u12_u6_U53 (.ZN( u0_u12_u6_n147 ) , .A2( u0_u12_u6_n98 ) , .A1( u0_u12_u6_n99 ) );
  NAND2_X1 u0_u12_u6_U54 (.ZN( u0_u12_u6_n128 ) , .A1( u0_u12_u6_n94 ) , .A2( u0_u12_u6_n96 ) );
  NAND2_X1 u0_u12_u6_U55 (.ZN( u0_u12_u6_n119 ) , .A2( u0_u12_u6_n95 ) , .A1( u0_u12_u6_n99 ) );
  NAND2_X1 u0_u12_u6_U56 (.ZN( u0_u12_u6_n123 ) , .A2( u0_u12_u6_n91 ) , .A1( u0_u12_u6_n96 ) );
  NAND2_X1 u0_u12_u6_U57 (.ZN( u0_u12_u6_n100 ) , .A2( u0_u12_u6_n92 ) , .A1( u0_u12_u6_n98 ) );
  NAND2_X1 u0_u12_u6_U58 (.ZN( u0_u12_u6_n122 ) , .A1( u0_u12_u6_n94 ) , .A2( u0_u12_u6_n97 ) );
  INV_X1 u0_u12_u6_U59 (.A( u0_u12_u6_n139 ) , .ZN( u0_u12_u6_n160 ) );
  AOI22_X1 u0_u12_u6_U6 (.B2( u0_u12_u6_n101 ) , .A1( u0_u12_u6_n102 ) , .ZN( u0_u12_u6_n103 ) , .B1( u0_u12_u6_n160 ) , .A2( u0_u12_u6_n161 ) );
  NAND2_X1 u0_u12_u6_U60 (.ZN( u0_u12_u6_n113 ) , .A1( u0_u12_u6_n96 ) , .A2( u0_u12_u6_n98 ) );
  NOR2_X1 u0_u12_u6_U61 (.A2( u0_u12_X_40 ) , .A1( u0_u12_X_41 ) , .ZN( u0_u12_u6_n126 ) );
  NOR2_X1 u0_u12_u6_U62 (.A2( u0_u12_X_39 ) , .A1( u0_u12_X_42 ) , .ZN( u0_u12_u6_n92 ) );
  NOR2_X1 u0_u12_u6_U63 (.A2( u0_u12_X_39 ) , .A1( u0_u12_u6_n156 ) , .ZN( u0_u12_u6_n97 ) );
  NOR2_X1 u0_u12_u6_U64 (.A2( u0_u12_X_38 ) , .A1( u0_u12_u6_n165 ) , .ZN( u0_u12_u6_n95 ) );
  NOR2_X1 u0_u12_u6_U65 (.A2( u0_u12_X_41 ) , .ZN( u0_u12_u6_n111 ) , .A1( u0_u12_u6_n157 ) );
  NOR2_X1 u0_u12_u6_U66 (.A2( u0_u12_X_37 ) , .A1( u0_u12_u6_n162 ) , .ZN( u0_u12_u6_n94 ) );
  NOR2_X1 u0_u12_u6_U67 (.A2( u0_u12_X_37 ) , .A1( u0_u12_X_38 ) , .ZN( u0_u12_u6_n91 ) );
  NAND2_X1 u0_u12_u6_U68 (.A1( u0_u12_X_41 ) , .ZN( u0_u12_u6_n144 ) , .A2( u0_u12_u6_n157 ) );
  NAND2_X1 u0_u12_u6_U69 (.A2( u0_u12_X_40 ) , .A1( u0_u12_X_41 ) , .ZN( u0_u12_u6_n139 ) );
  NOR2_X1 u0_u12_u6_U7 (.A1( u0_u12_u6_n118 ) , .ZN( u0_u12_u6_n143 ) , .A2( u0_u12_u6_n168 ) );
  AND2_X1 u0_u12_u6_U70 (.A1( u0_u12_X_39 ) , .A2( u0_u12_u6_n156 ) , .ZN( u0_u12_u6_n96 ) );
  AND2_X1 u0_u12_u6_U71 (.A1( u0_u12_X_39 ) , .A2( u0_u12_X_42 ) , .ZN( u0_u12_u6_n99 ) );
  INV_X1 u0_u12_u6_U72 (.A( u0_u12_X_40 ) , .ZN( u0_u12_u6_n157 ) );
  INV_X1 u0_u12_u6_U73 (.A( u0_u12_X_37 ) , .ZN( u0_u12_u6_n165 ) );
  INV_X1 u0_u12_u6_U74 (.A( u0_u12_X_38 ) , .ZN( u0_u12_u6_n162 ) );
  INV_X1 u0_u12_u6_U75 (.A( u0_u12_X_42 ) , .ZN( u0_u12_u6_n156 ) );
  NAND4_X1 u0_u12_u6_U76 (.ZN( u0_out12_32 ) , .A4( u0_u12_u6_n103 ) , .A3( u0_u12_u6_n104 ) , .A2( u0_u12_u6_n105 ) , .A1( u0_u12_u6_n106 ) );
  AOI22_X1 u0_u12_u6_U77 (.ZN( u0_u12_u6_n105 ) , .A2( u0_u12_u6_n108 ) , .A1( u0_u12_u6_n118 ) , .B2( u0_u12_u6_n126 ) , .B1( u0_u12_u6_n171 ) );
  AOI22_X1 u0_u12_u6_U78 (.ZN( u0_u12_u6_n104 ) , .A1( u0_u12_u6_n111 ) , .B1( u0_u12_u6_n124 ) , .B2( u0_u12_u6_n151 ) , .A2( u0_u12_u6_n93 ) );
  NAND4_X1 u0_u12_u6_U79 (.ZN( u0_out12_12 ) , .A4( u0_u12_u6_n114 ) , .A3( u0_u12_u6_n115 ) , .A2( u0_u12_u6_n116 ) , .A1( u0_u12_u6_n117 ) );
  INV_X1 u0_u12_u6_U8 (.ZN( u0_u12_u6_n172 ) , .A( u0_u12_u6_n88 ) );
  OAI22_X1 u0_u12_u6_U80 (.B2( u0_u12_u6_n111 ) , .ZN( u0_u12_u6_n116 ) , .B1( u0_u12_u6_n126 ) , .A2( u0_u12_u6_n164 ) , .A1( u0_u12_u6_n167 ) );
  OAI21_X1 u0_u12_u6_U81 (.A( u0_u12_u6_n108 ) , .ZN( u0_u12_u6_n117 ) , .B2( u0_u12_u6_n141 ) , .B1( u0_u12_u6_n163 ) );
  OAI211_X1 u0_u12_u6_U82 (.ZN( u0_out12_22 ) , .B( u0_u12_u6_n137 ) , .A( u0_u12_u6_n138 ) , .C2( u0_u12_u6_n139 ) , .C1( u0_u12_u6_n140 ) );
  AOI22_X1 u0_u12_u6_U83 (.B1( u0_u12_u6_n124 ) , .A2( u0_u12_u6_n125 ) , .A1( u0_u12_u6_n126 ) , .ZN( u0_u12_u6_n138 ) , .B2( u0_u12_u6_n161 ) );
  AND4_X1 u0_u12_u6_U84 (.A3( u0_u12_u6_n119 ) , .A1( u0_u12_u6_n120 ) , .A4( u0_u12_u6_n129 ) , .ZN( u0_u12_u6_n140 ) , .A2( u0_u12_u6_n143 ) );
  OAI211_X1 u0_u12_u6_U85 (.ZN( u0_out12_7 ) , .B( u0_u12_u6_n153 ) , .C2( u0_u12_u6_n154 ) , .C1( u0_u12_u6_n155 ) , .A( u0_u12_u6_n174 ) );
  NOR3_X1 u0_u12_u6_U86 (.A1( u0_u12_u6_n141 ) , .ZN( u0_u12_u6_n154 ) , .A3( u0_u12_u6_n164 ) , .A2( u0_u12_u6_n171 ) );
  AOI211_X1 u0_u12_u6_U87 (.B( u0_u12_u6_n149 ) , .A( u0_u12_u6_n150 ) , .C2( u0_u12_u6_n151 ) , .C1( u0_u12_u6_n152 ) , .ZN( u0_u12_u6_n153 ) );
  NAND3_X1 u0_u12_u6_U88 (.A2( u0_u12_u6_n123 ) , .ZN( u0_u12_u6_n125 ) , .A1( u0_u12_u6_n130 ) , .A3( u0_u12_u6_n131 ) );
  NAND3_X1 u0_u12_u6_U89 (.A3( u0_u12_u6_n133 ) , .ZN( u0_u12_u6_n141 ) , .A1( u0_u12_u6_n145 ) , .A2( u0_u12_u6_n148 ) );
  OAI21_X1 u0_u12_u6_U9 (.A( u0_u12_u6_n159 ) , .B1( u0_u12_u6_n169 ) , .B2( u0_u12_u6_n173 ) , .ZN( u0_u12_u6_n90 ) );
  NAND3_X1 u0_u12_u6_U90 (.ZN( u0_u12_u6_n101 ) , .A3( u0_u12_u6_n107 ) , .A2( u0_u12_u6_n121 ) , .A1( u0_u12_u6_n127 ) );
  NAND3_X1 u0_u12_u6_U91 (.ZN( u0_u12_u6_n102 ) , .A3( u0_u12_u6_n130 ) , .A2( u0_u12_u6_n145 ) , .A1( u0_u12_u6_n166 ) );
  NAND3_X1 u0_u12_u6_U92 (.A3( u0_u12_u6_n113 ) , .A1( u0_u12_u6_n119 ) , .A2( u0_u12_u6_n123 ) , .ZN( u0_u12_u6_n93 ) );
  NAND3_X1 u0_u12_u6_U93 (.ZN( u0_u12_u6_n142 ) , .A2( u0_u12_u6_n172 ) , .A3( u0_u12_u6_n89 ) , .A1( u0_u12_u6_n90 ) );
  XOR2_X1 u0_u15_U13 (.A( u0_FP_61 ) , .B( u0_K16_42 ) , .Z( u0_u15_X_42 ) );
  XOR2_X1 u0_u15_U14 (.A( u0_FP_60 ) , .B( u0_K16_41 ) , .Z( u0_u15_X_41 ) );
  XOR2_X1 u0_u15_U15 (.A( u0_FP_59 ) , .B( u0_K16_40 ) , .Z( u0_u15_X_40 ) );
  XOR2_X1 u0_u15_U17 (.A( u0_FP_58 ) , .B( u0_K16_39 ) , .Z( u0_u15_X_39 ) );
  XOR2_X1 u0_u15_U18 (.A( u0_FP_57 ) , .B( u0_K16_38 ) , .Z( u0_u15_X_38 ) );
  XOR2_X1 u0_u15_U19 (.A( u0_FP_56 ) , .B( u0_K16_37 ) , .Z( u0_u15_X_37 ) );
  XOR2_X1 u0_u15_U20 (.A( u0_FP_57 ) , .B( u0_K16_36 ) , .Z( u0_u15_X_36 ) );
  XOR2_X1 u0_u15_U21 (.A( u0_FP_56 ) , .B( u0_K16_35 ) , .Z( u0_u15_X_35 ) );
  XOR2_X1 u0_u15_U22 (.A( u0_FP_55 ) , .B( u0_K16_34 ) , .Z( u0_u15_X_34 ) );
  XOR2_X1 u0_u15_U23 (.A( u0_FP_54 ) , .B( u0_K16_33 ) , .Z( u0_u15_X_33 ) );
  XOR2_X1 u0_u15_U24 (.A( u0_FP_53 ) , .B( u0_K16_32 ) , .Z( u0_u15_X_32 ) );
  XOR2_X1 u0_u15_U25 (.A( u0_FP_52 ) , .B( u0_K16_31 ) , .Z( u0_u15_X_31 ) );
  XOR2_X1 u0_u15_U26 (.A( u0_FP_53 ) , .B( u0_K16_30 ) , .Z( u0_u15_X_30 ) );
  XOR2_X1 u0_u15_U28 (.A( u0_FP_52 ) , .B( u0_K16_29 ) , .Z( u0_u15_X_29 ) );
  XOR2_X1 u0_u15_U29 (.A( u0_FP_51 ) , .B( u0_K16_28 ) , .Z( u0_u15_X_28 ) );
  XOR2_X1 u0_u15_U30 (.A( u0_FP_50 ) , .B( u0_K16_27 ) , .Z( u0_u15_X_27 ) );
  XOR2_X1 u0_u15_U31 (.A( u0_FP_49 ) , .B( u0_K16_26 ) , .Z( u0_u15_X_26 ) );
  XOR2_X1 u0_u15_U32 (.A( u0_FP_48 ) , .B( u0_K16_25 ) , .Z( u0_u15_X_25 ) );
  OAI22_X1 u0_u15_u4_U10 (.B2( u0_u15_u4_n135 ) , .ZN( u0_u15_u4_n137 ) , .B1( u0_u15_u4_n153 ) , .A1( u0_u15_u4_n155 ) , .A2( u0_u15_u4_n171 ) );
  AND3_X1 u0_u15_u4_U11 (.A2( u0_u15_u4_n134 ) , .ZN( u0_u15_u4_n135 ) , .A3( u0_u15_u4_n145 ) , .A1( u0_u15_u4_n157 ) );
  OR3_X1 u0_u15_u4_U12 (.A3( u0_u15_u4_n114 ) , .A2( u0_u15_u4_n115 ) , .A1( u0_u15_u4_n116 ) , .ZN( u0_u15_u4_n136 ) );
  AOI21_X1 u0_u15_u4_U13 (.A( u0_u15_u4_n113 ) , .ZN( u0_u15_u4_n116 ) , .B2( u0_u15_u4_n173 ) , .B1( u0_u15_u4_n174 ) );
  AOI21_X1 u0_u15_u4_U14 (.ZN( u0_u15_u4_n115 ) , .B2( u0_u15_u4_n145 ) , .B1( u0_u15_u4_n146 ) , .A( u0_u15_u4_n156 ) );
  OAI22_X1 u0_u15_u4_U15 (.ZN( u0_u15_u4_n114 ) , .A2( u0_u15_u4_n121 ) , .B1( u0_u15_u4_n160 ) , .B2( u0_u15_u4_n170 ) , .A1( u0_u15_u4_n171 ) );
  NAND2_X1 u0_u15_u4_U16 (.ZN( u0_u15_u4_n132 ) , .A2( u0_u15_u4_n170 ) , .A1( u0_u15_u4_n173 ) );
  AOI21_X1 u0_u15_u4_U17 (.B2( u0_u15_u4_n160 ) , .B1( u0_u15_u4_n161 ) , .ZN( u0_u15_u4_n162 ) , .A( u0_u15_u4_n170 ) );
  AOI21_X1 u0_u15_u4_U18 (.ZN( u0_u15_u4_n107 ) , .B2( u0_u15_u4_n143 ) , .A( u0_u15_u4_n174 ) , .B1( u0_u15_u4_n184 ) );
  AOI21_X1 u0_u15_u4_U19 (.B2( u0_u15_u4_n158 ) , .B1( u0_u15_u4_n159 ) , .ZN( u0_u15_u4_n163 ) , .A( u0_u15_u4_n174 ) );
  AOI21_X1 u0_u15_u4_U20 (.A( u0_u15_u4_n153 ) , .B2( u0_u15_u4_n154 ) , .B1( u0_u15_u4_n155 ) , .ZN( u0_u15_u4_n165 ) );
  AOI21_X1 u0_u15_u4_U21 (.A( u0_u15_u4_n156 ) , .B2( u0_u15_u4_n157 ) , .ZN( u0_u15_u4_n164 ) , .B1( u0_u15_u4_n184 ) );
  INV_X1 u0_u15_u4_U22 (.A( u0_u15_u4_n138 ) , .ZN( u0_u15_u4_n170 ) );
  AND2_X1 u0_u15_u4_U23 (.A2( u0_u15_u4_n120 ) , .ZN( u0_u15_u4_n155 ) , .A1( u0_u15_u4_n160 ) );
  INV_X1 u0_u15_u4_U24 (.A( u0_u15_u4_n156 ) , .ZN( u0_u15_u4_n175 ) );
  NAND2_X1 u0_u15_u4_U25 (.A2( u0_u15_u4_n118 ) , .ZN( u0_u15_u4_n131 ) , .A1( u0_u15_u4_n147 ) );
  NAND2_X1 u0_u15_u4_U26 (.A1( u0_u15_u4_n119 ) , .A2( u0_u15_u4_n120 ) , .ZN( u0_u15_u4_n130 ) );
  NAND2_X1 u0_u15_u4_U27 (.ZN( u0_u15_u4_n117 ) , .A2( u0_u15_u4_n118 ) , .A1( u0_u15_u4_n148 ) );
  NAND2_X1 u0_u15_u4_U28 (.ZN( u0_u15_u4_n129 ) , .A1( u0_u15_u4_n134 ) , .A2( u0_u15_u4_n148 ) );
  AND3_X1 u0_u15_u4_U29 (.A1( u0_u15_u4_n119 ) , .A2( u0_u15_u4_n143 ) , .A3( u0_u15_u4_n154 ) , .ZN( u0_u15_u4_n161 ) );
  NOR2_X1 u0_u15_u4_U3 (.ZN( u0_u15_u4_n121 ) , .A1( u0_u15_u4_n181 ) , .A2( u0_u15_u4_n182 ) );
  AND2_X1 u0_u15_u4_U30 (.A1( u0_u15_u4_n145 ) , .A2( u0_u15_u4_n147 ) , .ZN( u0_u15_u4_n159 ) );
  INV_X1 u0_u15_u4_U31 (.A( u0_u15_u4_n158 ) , .ZN( u0_u15_u4_n182 ) );
  INV_X1 u0_u15_u4_U32 (.ZN( u0_u15_u4_n181 ) , .A( u0_u15_u4_n96 ) );
  INV_X1 u0_u15_u4_U33 (.A( u0_u15_u4_n144 ) , .ZN( u0_u15_u4_n179 ) );
  INV_X1 u0_u15_u4_U34 (.A( u0_u15_u4_n157 ) , .ZN( u0_u15_u4_n178 ) );
  NAND2_X1 u0_u15_u4_U35 (.A2( u0_u15_u4_n154 ) , .A1( u0_u15_u4_n96 ) , .ZN( u0_u15_u4_n97 ) );
  INV_X1 u0_u15_u4_U36 (.ZN( u0_u15_u4_n186 ) , .A( u0_u15_u4_n95 ) );
  OAI221_X1 u0_u15_u4_U37 (.C1( u0_u15_u4_n134 ) , .B1( u0_u15_u4_n158 ) , .B2( u0_u15_u4_n171 ) , .C2( u0_u15_u4_n173 ) , .A( u0_u15_u4_n94 ) , .ZN( u0_u15_u4_n95 ) );
  AOI222_X1 u0_u15_u4_U38 (.B2( u0_u15_u4_n132 ) , .A1( u0_u15_u4_n138 ) , .C2( u0_u15_u4_n175 ) , .A2( u0_u15_u4_n179 ) , .C1( u0_u15_u4_n181 ) , .B1( u0_u15_u4_n185 ) , .ZN( u0_u15_u4_n94 ) );
  INV_X1 u0_u15_u4_U39 (.A( u0_u15_u4_n113 ) , .ZN( u0_u15_u4_n185 ) );
  INV_X1 u0_u15_u4_U4 (.A( u0_u15_u4_n117 ) , .ZN( u0_u15_u4_n184 ) );
  INV_X1 u0_u15_u4_U40 (.A( u0_u15_u4_n143 ) , .ZN( u0_u15_u4_n183 ) );
  NOR2_X1 u0_u15_u4_U41 (.ZN( u0_u15_u4_n138 ) , .A1( u0_u15_u4_n168 ) , .A2( u0_u15_u4_n169 ) );
  NOR2_X1 u0_u15_u4_U42 (.A1( u0_u15_u4_n150 ) , .A2( u0_u15_u4_n152 ) , .ZN( u0_u15_u4_n153 ) );
  NOR2_X1 u0_u15_u4_U43 (.A2( u0_u15_u4_n128 ) , .A1( u0_u15_u4_n138 ) , .ZN( u0_u15_u4_n156 ) );
  AOI22_X1 u0_u15_u4_U44 (.B2( u0_u15_u4_n122 ) , .A1( u0_u15_u4_n123 ) , .ZN( u0_u15_u4_n124 ) , .B1( u0_u15_u4_n128 ) , .A2( u0_u15_u4_n172 ) );
  NAND2_X1 u0_u15_u4_U45 (.A2( u0_u15_u4_n120 ) , .ZN( u0_u15_u4_n123 ) , .A1( u0_u15_u4_n161 ) );
  INV_X1 u0_u15_u4_U46 (.A( u0_u15_u4_n153 ) , .ZN( u0_u15_u4_n172 ) );
  AOI22_X1 u0_u15_u4_U47 (.B2( u0_u15_u4_n132 ) , .A2( u0_u15_u4_n133 ) , .ZN( u0_u15_u4_n140 ) , .A1( u0_u15_u4_n150 ) , .B1( u0_u15_u4_n179 ) );
  NAND2_X1 u0_u15_u4_U48 (.ZN( u0_u15_u4_n133 ) , .A2( u0_u15_u4_n146 ) , .A1( u0_u15_u4_n154 ) );
  NAND2_X1 u0_u15_u4_U49 (.A1( u0_u15_u4_n103 ) , .ZN( u0_u15_u4_n154 ) , .A2( u0_u15_u4_n98 ) );
  NOR4_X1 u0_u15_u4_U5 (.A4( u0_u15_u4_n106 ) , .A3( u0_u15_u4_n107 ) , .A2( u0_u15_u4_n108 ) , .A1( u0_u15_u4_n109 ) , .ZN( u0_u15_u4_n110 ) );
  NAND2_X1 u0_u15_u4_U50 (.A1( u0_u15_u4_n101 ) , .ZN( u0_u15_u4_n158 ) , .A2( u0_u15_u4_n99 ) );
  AOI21_X1 u0_u15_u4_U51 (.ZN( u0_u15_u4_n127 ) , .A( u0_u15_u4_n136 ) , .B2( u0_u15_u4_n150 ) , .B1( u0_u15_u4_n180 ) );
  INV_X1 u0_u15_u4_U52 (.A( u0_u15_u4_n160 ) , .ZN( u0_u15_u4_n180 ) );
  NAND2_X1 u0_u15_u4_U53 (.A2( u0_u15_u4_n104 ) , .A1( u0_u15_u4_n105 ) , .ZN( u0_u15_u4_n146 ) );
  NAND2_X1 u0_u15_u4_U54 (.A2( u0_u15_u4_n101 ) , .A1( u0_u15_u4_n102 ) , .ZN( u0_u15_u4_n160 ) );
  NAND2_X1 u0_u15_u4_U55 (.ZN( u0_u15_u4_n134 ) , .A1( u0_u15_u4_n98 ) , .A2( u0_u15_u4_n99 ) );
  NAND2_X1 u0_u15_u4_U56 (.A1( u0_u15_u4_n103 ) , .A2( u0_u15_u4_n104 ) , .ZN( u0_u15_u4_n143 ) );
  NAND2_X1 u0_u15_u4_U57 (.A2( u0_u15_u4_n105 ) , .ZN( u0_u15_u4_n145 ) , .A1( u0_u15_u4_n98 ) );
  NAND2_X1 u0_u15_u4_U58 (.A1( u0_u15_u4_n100 ) , .A2( u0_u15_u4_n105 ) , .ZN( u0_u15_u4_n120 ) );
  NAND2_X1 u0_u15_u4_U59 (.A1( u0_u15_u4_n102 ) , .A2( u0_u15_u4_n104 ) , .ZN( u0_u15_u4_n148 ) );
  AOI21_X1 u0_u15_u4_U6 (.ZN( u0_u15_u4_n106 ) , .B2( u0_u15_u4_n146 ) , .B1( u0_u15_u4_n158 ) , .A( u0_u15_u4_n170 ) );
  NAND2_X1 u0_u15_u4_U60 (.A2( u0_u15_u4_n100 ) , .A1( u0_u15_u4_n103 ) , .ZN( u0_u15_u4_n157 ) );
  INV_X1 u0_u15_u4_U61 (.A( u0_u15_u4_n150 ) , .ZN( u0_u15_u4_n173 ) );
  INV_X1 u0_u15_u4_U62 (.A( u0_u15_u4_n152 ) , .ZN( u0_u15_u4_n171 ) );
  NAND2_X1 u0_u15_u4_U63 (.A1( u0_u15_u4_n100 ) , .ZN( u0_u15_u4_n118 ) , .A2( u0_u15_u4_n99 ) );
  NAND2_X1 u0_u15_u4_U64 (.A2( u0_u15_u4_n100 ) , .A1( u0_u15_u4_n102 ) , .ZN( u0_u15_u4_n144 ) );
  NAND2_X1 u0_u15_u4_U65 (.A2( u0_u15_u4_n101 ) , .A1( u0_u15_u4_n105 ) , .ZN( u0_u15_u4_n96 ) );
  INV_X1 u0_u15_u4_U66 (.A( u0_u15_u4_n128 ) , .ZN( u0_u15_u4_n174 ) );
  NAND2_X1 u0_u15_u4_U67 (.A2( u0_u15_u4_n102 ) , .ZN( u0_u15_u4_n119 ) , .A1( u0_u15_u4_n98 ) );
  NAND2_X1 u0_u15_u4_U68 (.A2( u0_u15_u4_n101 ) , .A1( u0_u15_u4_n103 ) , .ZN( u0_u15_u4_n147 ) );
  NAND2_X1 u0_u15_u4_U69 (.A2( u0_u15_u4_n104 ) , .ZN( u0_u15_u4_n113 ) , .A1( u0_u15_u4_n99 ) );
  AOI21_X1 u0_u15_u4_U7 (.ZN( u0_u15_u4_n108 ) , .B2( u0_u15_u4_n134 ) , .B1( u0_u15_u4_n155 ) , .A( u0_u15_u4_n156 ) );
  NOR2_X1 u0_u15_u4_U70 (.A2( u0_u15_X_28 ) , .ZN( u0_u15_u4_n150 ) , .A1( u0_u15_u4_n168 ) );
  NOR2_X1 u0_u15_u4_U71 (.A2( u0_u15_X_29 ) , .ZN( u0_u15_u4_n152 ) , .A1( u0_u15_u4_n169 ) );
  NOR2_X1 u0_u15_u4_U72 (.A2( u0_u15_X_26 ) , .ZN( u0_u15_u4_n100 ) , .A1( u0_u15_u4_n177 ) );
  NOR2_X1 u0_u15_u4_U73 (.A2( u0_u15_X_30 ) , .ZN( u0_u15_u4_n105 ) , .A1( u0_u15_u4_n176 ) );
  NOR2_X1 u0_u15_u4_U74 (.A2( u0_u15_X_28 ) , .A1( u0_u15_X_29 ) , .ZN( u0_u15_u4_n128 ) );
  NOR2_X1 u0_u15_u4_U75 (.A2( u0_u15_X_25 ) , .A1( u0_u15_X_26 ) , .ZN( u0_u15_u4_n98 ) );
  NOR2_X1 u0_u15_u4_U76 (.A2( u0_u15_X_27 ) , .A1( u0_u15_X_30 ) , .ZN( u0_u15_u4_n102 ) );
  AND2_X1 u0_u15_u4_U77 (.A2( u0_u15_X_25 ) , .A1( u0_u15_X_26 ) , .ZN( u0_u15_u4_n104 ) );
  AND2_X1 u0_u15_u4_U78 (.A1( u0_u15_X_30 ) , .A2( u0_u15_u4_n176 ) , .ZN( u0_u15_u4_n99 ) );
  AND2_X1 u0_u15_u4_U79 (.A1( u0_u15_X_26 ) , .ZN( u0_u15_u4_n101 ) , .A2( u0_u15_u4_n177 ) );
  AOI21_X1 u0_u15_u4_U8 (.ZN( u0_u15_u4_n109 ) , .A( u0_u15_u4_n153 ) , .B1( u0_u15_u4_n159 ) , .B2( u0_u15_u4_n184 ) );
  AND2_X1 u0_u15_u4_U80 (.A1( u0_u15_X_27 ) , .A2( u0_u15_X_30 ) , .ZN( u0_u15_u4_n103 ) );
  INV_X1 u0_u15_u4_U81 (.A( u0_u15_X_28 ) , .ZN( u0_u15_u4_n169 ) );
  INV_X1 u0_u15_u4_U82 (.A( u0_u15_X_29 ) , .ZN( u0_u15_u4_n168 ) );
  INV_X1 u0_u15_u4_U83 (.A( u0_u15_X_25 ) , .ZN( u0_u15_u4_n177 ) );
  INV_X1 u0_u15_u4_U84 (.A( u0_u15_X_27 ) , .ZN( u0_u15_u4_n176 ) );
  NAND4_X1 u0_u15_u4_U85 (.ZN( u0_out15_25 ) , .A4( u0_u15_u4_n139 ) , .A3( u0_u15_u4_n140 ) , .A2( u0_u15_u4_n141 ) , .A1( u0_u15_u4_n142 ) );
  OAI21_X1 u0_u15_u4_U86 (.A( u0_u15_u4_n128 ) , .B2( u0_u15_u4_n129 ) , .B1( u0_u15_u4_n130 ) , .ZN( u0_u15_u4_n142 ) );
  OAI21_X1 u0_u15_u4_U87 (.B2( u0_u15_u4_n131 ) , .ZN( u0_u15_u4_n141 ) , .A( u0_u15_u4_n175 ) , .B1( u0_u15_u4_n183 ) );
  NAND4_X1 u0_u15_u4_U88 (.ZN( u0_out15_14 ) , .A4( u0_u15_u4_n124 ) , .A3( u0_u15_u4_n125 ) , .A2( u0_u15_u4_n126 ) , .A1( u0_u15_u4_n127 ) );
  AOI22_X1 u0_u15_u4_U89 (.B2( u0_u15_u4_n117 ) , .ZN( u0_u15_u4_n126 ) , .A1( u0_u15_u4_n129 ) , .B1( u0_u15_u4_n152 ) , .A2( u0_u15_u4_n175 ) );
  AOI211_X1 u0_u15_u4_U9 (.B( u0_u15_u4_n136 ) , .A( u0_u15_u4_n137 ) , .C2( u0_u15_u4_n138 ) , .ZN( u0_u15_u4_n139 ) , .C1( u0_u15_u4_n182 ) );
  AOI22_X1 u0_u15_u4_U90 (.ZN( u0_u15_u4_n125 ) , .B2( u0_u15_u4_n131 ) , .A2( u0_u15_u4_n132 ) , .B1( u0_u15_u4_n138 ) , .A1( u0_u15_u4_n178 ) );
  AOI22_X1 u0_u15_u4_U91 (.B2( u0_u15_u4_n149 ) , .B1( u0_u15_u4_n150 ) , .A2( u0_u15_u4_n151 ) , .A1( u0_u15_u4_n152 ) , .ZN( u0_u15_u4_n167 ) );
  NOR4_X1 u0_u15_u4_U92 (.A4( u0_u15_u4_n162 ) , .A3( u0_u15_u4_n163 ) , .A2( u0_u15_u4_n164 ) , .A1( u0_u15_u4_n165 ) , .ZN( u0_u15_u4_n166 ) );
  NAND4_X1 u0_u15_u4_U93 (.ZN( u0_out15_8 ) , .A4( u0_u15_u4_n110 ) , .A3( u0_u15_u4_n111 ) , .A2( u0_u15_u4_n112 ) , .A1( u0_u15_u4_n186 ) );
  NAND2_X1 u0_u15_u4_U94 (.ZN( u0_u15_u4_n112 ) , .A2( u0_u15_u4_n130 ) , .A1( u0_u15_u4_n150 ) );
  AOI22_X1 u0_u15_u4_U95 (.ZN( u0_u15_u4_n111 ) , .B2( u0_u15_u4_n132 ) , .A1( u0_u15_u4_n152 ) , .B1( u0_u15_u4_n178 ) , .A2( u0_u15_u4_n97 ) );
  NAND3_X1 u0_u15_u4_U96 (.ZN( u0_out15_3 ) , .A3( u0_u15_u4_n166 ) , .A1( u0_u15_u4_n167 ) , .A2( u0_u15_u4_n186 ) );
  NAND3_X1 u0_u15_u4_U97 (.A3( u0_u15_u4_n146 ) , .A2( u0_u15_u4_n147 ) , .A1( u0_u15_u4_n148 ) , .ZN( u0_u15_u4_n149 ) );
  NAND3_X1 u0_u15_u4_U98 (.A3( u0_u15_u4_n143 ) , .A2( u0_u15_u4_n144 ) , .A1( u0_u15_u4_n145 ) , .ZN( u0_u15_u4_n151 ) );
  NAND3_X1 u0_u15_u4_U99 (.A3( u0_u15_u4_n121 ) , .ZN( u0_u15_u4_n122 ) , .A2( u0_u15_u4_n144 ) , .A1( u0_u15_u4_n154 ) );
  INV_X1 u0_u15_u5_U10 (.A( u0_u15_u5_n121 ) , .ZN( u0_u15_u5_n177 ) );
  AOI222_X1 u0_u15_u5_U100 (.ZN( u0_u15_u5_n113 ) , .A1( u0_u15_u5_n131 ) , .C1( u0_u15_u5_n148 ) , .B2( u0_u15_u5_n174 ) , .C2( u0_u15_u5_n178 ) , .A2( u0_u15_u5_n179 ) , .B1( u0_u15_u5_n99 ) );
  NAND4_X1 u0_u15_u5_U101 (.ZN( u0_out15_29 ) , .A4( u0_u15_u5_n129 ) , .A3( u0_u15_u5_n130 ) , .A2( u0_u15_u5_n168 ) , .A1( u0_u15_u5_n196 ) );
  AOI221_X1 u0_u15_u5_U102 (.A( u0_u15_u5_n128 ) , .ZN( u0_u15_u5_n129 ) , .C2( u0_u15_u5_n132 ) , .B2( u0_u15_u5_n159 ) , .B1( u0_u15_u5_n176 ) , .C1( u0_u15_u5_n184 ) );
  AOI222_X1 u0_u15_u5_U103 (.ZN( u0_u15_u5_n130 ) , .A2( u0_u15_u5_n146 ) , .B1( u0_u15_u5_n147 ) , .C2( u0_u15_u5_n175 ) , .B2( u0_u15_u5_n179 ) , .A1( u0_u15_u5_n188 ) , .C1( u0_u15_u5_n194 ) );
  NAND3_X1 u0_u15_u5_U104 (.A2( u0_u15_u5_n154 ) , .A3( u0_u15_u5_n158 ) , .A1( u0_u15_u5_n161 ) , .ZN( u0_u15_u5_n99 ) );
  NOR2_X1 u0_u15_u5_U11 (.ZN( u0_u15_u5_n160 ) , .A2( u0_u15_u5_n173 ) , .A1( u0_u15_u5_n177 ) );
  INV_X1 u0_u15_u5_U12 (.A( u0_u15_u5_n150 ) , .ZN( u0_u15_u5_n174 ) );
  AOI21_X1 u0_u15_u5_U13 (.A( u0_u15_u5_n160 ) , .B2( u0_u15_u5_n161 ) , .ZN( u0_u15_u5_n162 ) , .B1( u0_u15_u5_n192 ) );
  INV_X1 u0_u15_u5_U14 (.A( u0_u15_u5_n159 ) , .ZN( u0_u15_u5_n192 ) );
  AOI21_X1 u0_u15_u5_U15 (.A( u0_u15_u5_n156 ) , .B2( u0_u15_u5_n157 ) , .B1( u0_u15_u5_n158 ) , .ZN( u0_u15_u5_n163 ) );
  AOI21_X1 u0_u15_u5_U16 (.B2( u0_u15_u5_n139 ) , .B1( u0_u15_u5_n140 ) , .ZN( u0_u15_u5_n141 ) , .A( u0_u15_u5_n150 ) );
  OAI21_X1 u0_u15_u5_U17 (.A( u0_u15_u5_n133 ) , .B2( u0_u15_u5_n134 ) , .B1( u0_u15_u5_n135 ) , .ZN( u0_u15_u5_n142 ) );
  OAI21_X1 u0_u15_u5_U18 (.ZN( u0_u15_u5_n133 ) , .B2( u0_u15_u5_n147 ) , .A( u0_u15_u5_n173 ) , .B1( u0_u15_u5_n188 ) );
  NAND2_X1 u0_u15_u5_U19 (.A2( u0_u15_u5_n119 ) , .A1( u0_u15_u5_n123 ) , .ZN( u0_u15_u5_n137 ) );
  INV_X1 u0_u15_u5_U20 (.A( u0_u15_u5_n155 ) , .ZN( u0_u15_u5_n194 ) );
  NAND2_X1 u0_u15_u5_U21 (.A1( u0_u15_u5_n121 ) , .ZN( u0_u15_u5_n132 ) , .A2( u0_u15_u5_n172 ) );
  NAND2_X1 u0_u15_u5_U22 (.A2( u0_u15_u5_n122 ) , .ZN( u0_u15_u5_n136 ) , .A1( u0_u15_u5_n154 ) );
  NAND2_X1 u0_u15_u5_U23 (.A2( u0_u15_u5_n119 ) , .A1( u0_u15_u5_n120 ) , .ZN( u0_u15_u5_n159 ) );
  INV_X1 u0_u15_u5_U24 (.A( u0_u15_u5_n156 ) , .ZN( u0_u15_u5_n175 ) );
  INV_X1 u0_u15_u5_U25 (.A( u0_u15_u5_n158 ) , .ZN( u0_u15_u5_n188 ) );
  INV_X1 u0_u15_u5_U26 (.A( u0_u15_u5_n152 ) , .ZN( u0_u15_u5_n179 ) );
  INV_X1 u0_u15_u5_U27 (.A( u0_u15_u5_n140 ) , .ZN( u0_u15_u5_n182 ) );
  INV_X1 u0_u15_u5_U28 (.A( u0_u15_u5_n151 ) , .ZN( u0_u15_u5_n183 ) );
  INV_X1 u0_u15_u5_U29 (.A( u0_u15_u5_n123 ) , .ZN( u0_u15_u5_n185 ) );
  NOR2_X1 u0_u15_u5_U3 (.ZN( u0_u15_u5_n134 ) , .A1( u0_u15_u5_n183 ) , .A2( u0_u15_u5_n190 ) );
  INV_X1 u0_u15_u5_U30 (.A( u0_u15_u5_n161 ) , .ZN( u0_u15_u5_n184 ) );
  INV_X1 u0_u15_u5_U31 (.A( u0_u15_u5_n139 ) , .ZN( u0_u15_u5_n189 ) );
  INV_X1 u0_u15_u5_U32 (.A( u0_u15_u5_n157 ) , .ZN( u0_u15_u5_n190 ) );
  INV_X1 u0_u15_u5_U33 (.A( u0_u15_u5_n120 ) , .ZN( u0_u15_u5_n193 ) );
  NAND2_X1 u0_u15_u5_U34 (.ZN( u0_u15_u5_n111 ) , .A1( u0_u15_u5_n140 ) , .A2( u0_u15_u5_n155 ) );
  NOR2_X1 u0_u15_u5_U35 (.ZN( u0_u15_u5_n100 ) , .A1( u0_u15_u5_n170 ) , .A2( u0_u15_u5_n180 ) );
  INV_X1 u0_u15_u5_U36 (.A( u0_u15_u5_n117 ) , .ZN( u0_u15_u5_n196 ) );
  OAI221_X1 u0_u15_u5_U37 (.A( u0_u15_u5_n116 ) , .ZN( u0_u15_u5_n117 ) , .B2( u0_u15_u5_n119 ) , .C1( u0_u15_u5_n153 ) , .C2( u0_u15_u5_n158 ) , .B1( u0_u15_u5_n172 ) );
  AOI222_X1 u0_u15_u5_U38 (.ZN( u0_u15_u5_n116 ) , .B2( u0_u15_u5_n145 ) , .C1( u0_u15_u5_n148 ) , .A2( u0_u15_u5_n174 ) , .C2( u0_u15_u5_n177 ) , .B1( u0_u15_u5_n187 ) , .A1( u0_u15_u5_n193 ) );
  INV_X1 u0_u15_u5_U39 (.A( u0_u15_u5_n115 ) , .ZN( u0_u15_u5_n187 ) );
  INV_X1 u0_u15_u5_U4 (.A( u0_u15_u5_n138 ) , .ZN( u0_u15_u5_n191 ) );
  AOI22_X1 u0_u15_u5_U40 (.B2( u0_u15_u5_n131 ) , .A2( u0_u15_u5_n146 ) , .ZN( u0_u15_u5_n169 ) , .B1( u0_u15_u5_n174 ) , .A1( u0_u15_u5_n185 ) );
  NOR2_X1 u0_u15_u5_U41 (.A1( u0_u15_u5_n146 ) , .ZN( u0_u15_u5_n150 ) , .A2( u0_u15_u5_n173 ) );
  AOI21_X1 u0_u15_u5_U42 (.A( u0_u15_u5_n118 ) , .B2( u0_u15_u5_n145 ) , .ZN( u0_u15_u5_n168 ) , .B1( u0_u15_u5_n186 ) );
  INV_X1 u0_u15_u5_U43 (.A( u0_u15_u5_n122 ) , .ZN( u0_u15_u5_n186 ) );
  NOR2_X1 u0_u15_u5_U44 (.A1( u0_u15_u5_n146 ) , .ZN( u0_u15_u5_n152 ) , .A2( u0_u15_u5_n176 ) );
  NOR2_X1 u0_u15_u5_U45 (.A1( u0_u15_u5_n115 ) , .ZN( u0_u15_u5_n118 ) , .A2( u0_u15_u5_n153 ) );
  NOR2_X1 u0_u15_u5_U46 (.A2( u0_u15_u5_n145 ) , .ZN( u0_u15_u5_n156 ) , .A1( u0_u15_u5_n174 ) );
  NOR2_X1 u0_u15_u5_U47 (.ZN( u0_u15_u5_n121 ) , .A2( u0_u15_u5_n145 ) , .A1( u0_u15_u5_n176 ) );
  AOI22_X1 u0_u15_u5_U48 (.ZN( u0_u15_u5_n114 ) , .A2( u0_u15_u5_n137 ) , .A1( u0_u15_u5_n145 ) , .B2( u0_u15_u5_n175 ) , .B1( u0_u15_u5_n193 ) );
  OAI211_X1 u0_u15_u5_U49 (.B( u0_u15_u5_n124 ) , .A( u0_u15_u5_n125 ) , .C2( u0_u15_u5_n126 ) , .C1( u0_u15_u5_n127 ) , .ZN( u0_u15_u5_n128 ) );
  OAI21_X1 u0_u15_u5_U5 (.B2( u0_u15_u5_n136 ) , .B1( u0_u15_u5_n137 ) , .ZN( u0_u15_u5_n138 ) , .A( u0_u15_u5_n177 ) );
  NOR3_X1 u0_u15_u5_U50 (.ZN( u0_u15_u5_n127 ) , .A1( u0_u15_u5_n136 ) , .A3( u0_u15_u5_n148 ) , .A2( u0_u15_u5_n182 ) );
  OAI21_X1 u0_u15_u5_U51 (.ZN( u0_u15_u5_n124 ) , .A( u0_u15_u5_n177 ) , .B2( u0_u15_u5_n183 ) , .B1( u0_u15_u5_n189 ) );
  OAI21_X1 u0_u15_u5_U52 (.ZN( u0_u15_u5_n125 ) , .A( u0_u15_u5_n174 ) , .B2( u0_u15_u5_n185 ) , .B1( u0_u15_u5_n190 ) );
  AOI21_X1 u0_u15_u5_U53 (.A( u0_u15_u5_n153 ) , .B2( u0_u15_u5_n154 ) , .B1( u0_u15_u5_n155 ) , .ZN( u0_u15_u5_n164 ) );
  AOI21_X1 u0_u15_u5_U54 (.ZN( u0_u15_u5_n110 ) , .B1( u0_u15_u5_n122 ) , .B2( u0_u15_u5_n139 ) , .A( u0_u15_u5_n153 ) );
  INV_X1 u0_u15_u5_U55 (.A( u0_u15_u5_n153 ) , .ZN( u0_u15_u5_n176 ) );
  INV_X1 u0_u15_u5_U56 (.A( u0_u15_u5_n126 ) , .ZN( u0_u15_u5_n173 ) );
  AND2_X1 u0_u15_u5_U57 (.A2( u0_u15_u5_n104 ) , .A1( u0_u15_u5_n107 ) , .ZN( u0_u15_u5_n147 ) );
  AND2_X1 u0_u15_u5_U58 (.A2( u0_u15_u5_n104 ) , .A1( u0_u15_u5_n108 ) , .ZN( u0_u15_u5_n148 ) );
  NAND2_X1 u0_u15_u5_U59 (.A1( u0_u15_u5_n105 ) , .A2( u0_u15_u5_n106 ) , .ZN( u0_u15_u5_n158 ) );
  INV_X1 u0_u15_u5_U6 (.A( u0_u15_u5_n135 ) , .ZN( u0_u15_u5_n178 ) );
  NAND2_X1 u0_u15_u5_U60 (.A2( u0_u15_u5_n108 ) , .A1( u0_u15_u5_n109 ) , .ZN( u0_u15_u5_n139 ) );
  NAND2_X1 u0_u15_u5_U61 (.A1( u0_u15_u5_n106 ) , .A2( u0_u15_u5_n108 ) , .ZN( u0_u15_u5_n119 ) );
  NAND2_X1 u0_u15_u5_U62 (.A2( u0_u15_u5_n103 ) , .A1( u0_u15_u5_n105 ) , .ZN( u0_u15_u5_n140 ) );
  NAND2_X1 u0_u15_u5_U63 (.A2( u0_u15_u5_n104 ) , .A1( u0_u15_u5_n105 ) , .ZN( u0_u15_u5_n155 ) );
  NAND2_X1 u0_u15_u5_U64 (.A2( u0_u15_u5_n106 ) , .A1( u0_u15_u5_n107 ) , .ZN( u0_u15_u5_n122 ) );
  NAND2_X1 u0_u15_u5_U65 (.A2( u0_u15_u5_n100 ) , .A1( u0_u15_u5_n106 ) , .ZN( u0_u15_u5_n115 ) );
  NAND2_X1 u0_u15_u5_U66 (.A2( u0_u15_u5_n100 ) , .A1( u0_u15_u5_n103 ) , .ZN( u0_u15_u5_n161 ) );
  NAND2_X1 u0_u15_u5_U67 (.A1( u0_u15_u5_n105 ) , .A2( u0_u15_u5_n109 ) , .ZN( u0_u15_u5_n154 ) );
  INV_X1 u0_u15_u5_U68 (.A( u0_u15_u5_n146 ) , .ZN( u0_u15_u5_n172 ) );
  NAND2_X1 u0_u15_u5_U69 (.A1( u0_u15_u5_n103 ) , .A2( u0_u15_u5_n108 ) , .ZN( u0_u15_u5_n123 ) );
  OAI22_X1 u0_u15_u5_U7 (.B2( u0_u15_u5_n149 ) , .B1( u0_u15_u5_n150 ) , .A2( u0_u15_u5_n151 ) , .A1( u0_u15_u5_n152 ) , .ZN( u0_u15_u5_n165 ) );
  NAND2_X1 u0_u15_u5_U70 (.A2( u0_u15_u5_n103 ) , .A1( u0_u15_u5_n107 ) , .ZN( u0_u15_u5_n151 ) );
  NAND2_X1 u0_u15_u5_U71 (.A2( u0_u15_u5_n107 ) , .A1( u0_u15_u5_n109 ) , .ZN( u0_u15_u5_n120 ) );
  NAND2_X1 u0_u15_u5_U72 (.A2( u0_u15_u5_n100 ) , .A1( u0_u15_u5_n109 ) , .ZN( u0_u15_u5_n157 ) );
  AND2_X1 u0_u15_u5_U73 (.A2( u0_u15_u5_n100 ) , .A1( u0_u15_u5_n104 ) , .ZN( u0_u15_u5_n131 ) );
  INV_X1 u0_u15_u5_U74 (.A( u0_u15_u5_n102 ) , .ZN( u0_u15_u5_n195 ) );
  OAI221_X1 u0_u15_u5_U75 (.A( u0_u15_u5_n101 ) , .ZN( u0_u15_u5_n102 ) , .C2( u0_u15_u5_n115 ) , .C1( u0_u15_u5_n126 ) , .B1( u0_u15_u5_n134 ) , .B2( u0_u15_u5_n160 ) );
  OAI21_X1 u0_u15_u5_U76 (.ZN( u0_u15_u5_n101 ) , .B1( u0_u15_u5_n137 ) , .A( u0_u15_u5_n146 ) , .B2( u0_u15_u5_n147 ) );
  NOR2_X1 u0_u15_u5_U77 (.A2( u0_u15_X_34 ) , .A1( u0_u15_X_35 ) , .ZN( u0_u15_u5_n145 ) );
  NOR2_X1 u0_u15_u5_U78 (.A2( u0_u15_X_34 ) , .ZN( u0_u15_u5_n146 ) , .A1( u0_u15_u5_n171 ) );
  NOR2_X1 u0_u15_u5_U79 (.A2( u0_u15_X_31 ) , .A1( u0_u15_X_32 ) , .ZN( u0_u15_u5_n103 ) );
  NOR3_X1 u0_u15_u5_U8 (.A2( u0_u15_u5_n147 ) , .A1( u0_u15_u5_n148 ) , .ZN( u0_u15_u5_n149 ) , .A3( u0_u15_u5_n194 ) );
  NOR2_X1 u0_u15_u5_U80 (.A2( u0_u15_X_36 ) , .ZN( u0_u15_u5_n105 ) , .A1( u0_u15_u5_n180 ) );
  NOR2_X1 u0_u15_u5_U81 (.A2( u0_u15_X_33 ) , .ZN( u0_u15_u5_n108 ) , .A1( u0_u15_u5_n170 ) );
  NOR2_X1 u0_u15_u5_U82 (.A2( u0_u15_X_33 ) , .A1( u0_u15_X_36 ) , .ZN( u0_u15_u5_n107 ) );
  NOR2_X1 u0_u15_u5_U83 (.A2( u0_u15_X_31 ) , .ZN( u0_u15_u5_n104 ) , .A1( u0_u15_u5_n181 ) );
  NAND2_X1 u0_u15_u5_U84 (.A2( u0_u15_X_34 ) , .A1( u0_u15_X_35 ) , .ZN( u0_u15_u5_n153 ) );
  NAND2_X1 u0_u15_u5_U85 (.A1( u0_u15_X_34 ) , .ZN( u0_u15_u5_n126 ) , .A2( u0_u15_u5_n171 ) );
  AND2_X1 u0_u15_u5_U86 (.A1( u0_u15_X_31 ) , .A2( u0_u15_X_32 ) , .ZN( u0_u15_u5_n106 ) );
  AND2_X1 u0_u15_u5_U87 (.A1( u0_u15_X_31 ) , .ZN( u0_u15_u5_n109 ) , .A2( u0_u15_u5_n181 ) );
  INV_X1 u0_u15_u5_U88 (.A( u0_u15_X_33 ) , .ZN( u0_u15_u5_n180 ) );
  INV_X1 u0_u15_u5_U89 (.A( u0_u15_X_35 ) , .ZN( u0_u15_u5_n171 ) );
  NOR2_X1 u0_u15_u5_U9 (.ZN( u0_u15_u5_n135 ) , .A1( u0_u15_u5_n173 ) , .A2( u0_u15_u5_n176 ) );
  INV_X1 u0_u15_u5_U90 (.A( u0_u15_X_36 ) , .ZN( u0_u15_u5_n170 ) );
  INV_X1 u0_u15_u5_U91 (.A( u0_u15_X_32 ) , .ZN( u0_u15_u5_n181 ) );
  NAND4_X1 u0_u15_u5_U92 (.ZN( u0_out15_19 ) , .A4( u0_u15_u5_n166 ) , .A3( u0_u15_u5_n167 ) , .A2( u0_u15_u5_n168 ) , .A1( u0_u15_u5_n169 ) );
  AOI22_X1 u0_u15_u5_U93 (.B2( u0_u15_u5_n145 ) , .A2( u0_u15_u5_n146 ) , .ZN( u0_u15_u5_n167 ) , .B1( u0_u15_u5_n182 ) , .A1( u0_u15_u5_n189 ) );
  NOR4_X1 u0_u15_u5_U94 (.A4( u0_u15_u5_n162 ) , .A3( u0_u15_u5_n163 ) , .A2( u0_u15_u5_n164 ) , .A1( u0_u15_u5_n165 ) , .ZN( u0_u15_u5_n166 ) );
  NAND4_X1 u0_u15_u5_U95 (.ZN( u0_out15_11 ) , .A4( u0_u15_u5_n143 ) , .A3( u0_u15_u5_n144 ) , .A2( u0_u15_u5_n169 ) , .A1( u0_u15_u5_n196 ) );
  AOI22_X1 u0_u15_u5_U96 (.A2( u0_u15_u5_n132 ) , .ZN( u0_u15_u5_n144 ) , .B2( u0_u15_u5_n145 ) , .B1( u0_u15_u5_n184 ) , .A1( u0_u15_u5_n194 ) );
  NOR3_X1 u0_u15_u5_U97 (.A3( u0_u15_u5_n141 ) , .A1( u0_u15_u5_n142 ) , .ZN( u0_u15_u5_n143 ) , .A2( u0_u15_u5_n191 ) );
  NAND4_X1 u0_u15_u5_U98 (.ZN( u0_out15_4 ) , .A4( u0_u15_u5_n112 ) , .A2( u0_u15_u5_n113 ) , .A1( u0_u15_u5_n114 ) , .A3( u0_u15_u5_n195 ) );
  AOI211_X1 u0_u15_u5_U99 (.A( u0_u15_u5_n110 ) , .C1( u0_u15_u5_n111 ) , .ZN( u0_u15_u5_n112 ) , .B( u0_u15_u5_n118 ) , .C2( u0_u15_u5_n177 ) );
  INV_X1 u0_u15_u6_U10 (.ZN( u0_u15_u6_n172 ) , .A( u0_u15_u6_n88 ) );
  OAI21_X1 u0_u15_u6_U11 (.A( u0_u15_u6_n159 ) , .B1( u0_u15_u6_n169 ) , .B2( u0_u15_u6_n173 ) , .ZN( u0_u15_u6_n90 ) );
  AOI22_X1 u0_u15_u6_U12 (.A2( u0_u15_u6_n151 ) , .B2( u0_u15_u6_n161 ) , .A1( u0_u15_u6_n167 ) , .B1( u0_u15_u6_n170 ) , .ZN( u0_u15_u6_n89 ) );
  AOI21_X1 u0_u15_u6_U13 (.ZN( u0_u15_u6_n106 ) , .A( u0_u15_u6_n142 ) , .B2( u0_u15_u6_n159 ) , .B1( u0_u15_u6_n164 ) );
  INV_X1 u0_u15_u6_U14 (.A( u0_u15_u6_n155 ) , .ZN( u0_u15_u6_n161 ) );
  INV_X1 u0_u15_u6_U15 (.A( u0_u15_u6_n128 ) , .ZN( u0_u15_u6_n164 ) );
  NAND2_X1 u0_u15_u6_U16 (.ZN( u0_u15_u6_n110 ) , .A1( u0_u15_u6_n122 ) , .A2( u0_u15_u6_n129 ) );
  NAND2_X1 u0_u15_u6_U17 (.ZN( u0_u15_u6_n124 ) , .A2( u0_u15_u6_n146 ) , .A1( u0_u15_u6_n148 ) );
  INV_X1 u0_u15_u6_U18 (.A( u0_u15_u6_n132 ) , .ZN( u0_u15_u6_n171 ) );
  AND2_X1 u0_u15_u6_U19 (.A1( u0_u15_u6_n100 ) , .ZN( u0_u15_u6_n130 ) , .A2( u0_u15_u6_n147 ) );
  INV_X1 u0_u15_u6_U20 (.A( u0_u15_u6_n127 ) , .ZN( u0_u15_u6_n173 ) );
  INV_X1 u0_u15_u6_U21 (.A( u0_u15_u6_n121 ) , .ZN( u0_u15_u6_n167 ) );
  INV_X1 u0_u15_u6_U22 (.A( u0_u15_u6_n100 ) , .ZN( u0_u15_u6_n169 ) );
  INV_X1 u0_u15_u6_U23 (.A( u0_u15_u6_n123 ) , .ZN( u0_u15_u6_n170 ) );
  INV_X1 u0_u15_u6_U24 (.A( u0_u15_u6_n113 ) , .ZN( u0_u15_u6_n168 ) );
  AND2_X1 u0_u15_u6_U25 (.A1( u0_u15_u6_n107 ) , .A2( u0_u15_u6_n119 ) , .ZN( u0_u15_u6_n133 ) );
  AND2_X1 u0_u15_u6_U26 (.A2( u0_u15_u6_n121 ) , .A1( u0_u15_u6_n122 ) , .ZN( u0_u15_u6_n131 ) );
  AND3_X1 u0_u15_u6_U27 (.ZN( u0_u15_u6_n120 ) , .A2( u0_u15_u6_n127 ) , .A1( u0_u15_u6_n132 ) , .A3( u0_u15_u6_n145 ) );
  INV_X1 u0_u15_u6_U28 (.A( u0_u15_u6_n146 ) , .ZN( u0_u15_u6_n163 ) );
  AOI222_X1 u0_u15_u6_U29 (.ZN( u0_u15_u6_n114 ) , .A1( u0_u15_u6_n118 ) , .A2( u0_u15_u6_n126 ) , .B2( u0_u15_u6_n151 ) , .C2( u0_u15_u6_n159 ) , .C1( u0_u15_u6_n168 ) , .B1( u0_u15_u6_n169 ) );
  INV_X1 u0_u15_u6_U3 (.A( u0_u15_u6_n110 ) , .ZN( u0_u15_u6_n166 ) );
  NOR2_X1 u0_u15_u6_U30 (.A1( u0_u15_u6_n162 ) , .A2( u0_u15_u6_n165 ) , .ZN( u0_u15_u6_n98 ) );
  NAND2_X1 u0_u15_u6_U31 (.A1( u0_u15_u6_n144 ) , .ZN( u0_u15_u6_n151 ) , .A2( u0_u15_u6_n158 ) );
  NAND2_X1 u0_u15_u6_U32 (.ZN( u0_u15_u6_n132 ) , .A1( u0_u15_u6_n91 ) , .A2( u0_u15_u6_n97 ) );
  AOI22_X1 u0_u15_u6_U33 (.B2( u0_u15_u6_n110 ) , .B1( u0_u15_u6_n111 ) , .A1( u0_u15_u6_n112 ) , .ZN( u0_u15_u6_n115 ) , .A2( u0_u15_u6_n161 ) );
  NAND4_X1 u0_u15_u6_U34 (.A3( u0_u15_u6_n109 ) , .ZN( u0_u15_u6_n112 ) , .A4( u0_u15_u6_n132 ) , .A2( u0_u15_u6_n147 ) , .A1( u0_u15_u6_n166 ) );
  NOR2_X1 u0_u15_u6_U35 (.ZN( u0_u15_u6_n109 ) , .A1( u0_u15_u6_n170 ) , .A2( u0_u15_u6_n173 ) );
  NOR2_X1 u0_u15_u6_U36 (.A2( u0_u15_u6_n126 ) , .ZN( u0_u15_u6_n155 ) , .A1( u0_u15_u6_n160 ) );
  NAND2_X1 u0_u15_u6_U37 (.ZN( u0_u15_u6_n146 ) , .A2( u0_u15_u6_n94 ) , .A1( u0_u15_u6_n99 ) );
  AOI21_X1 u0_u15_u6_U38 (.A( u0_u15_u6_n144 ) , .B2( u0_u15_u6_n145 ) , .B1( u0_u15_u6_n146 ) , .ZN( u0_u15_u6_n150 ) );
  AOI211_X1 u0_u15_u6_U39 (.B( u0_u15_u6_n134 ) , .A( u0_u15_u6_n135 ) , .C1( u0_u15_u6_n136 ) , .ZN( u0_u15_u6_n137 ) , .C2( u0_u15_u6_n151 ) );
  INV_X1 u0_u15_u6_U4 (.A( u0_u15_u6_n142 ) , .ZN( u0_u15_u6_n174 ) );
  NAND4_X1 u0_u15_u6_U40 (.A4( u0_u15_u6_n127 ) , .A3( u0_u15_u6_n128 ) , .A2( u0_u15_u6_n129 ) , .A1( u0_u15_u6_n130 ) , .ZN( u0_u15_u6_n136 ) );
  AOI21_X1 u0_u15_u6_U41 (.B2( u0_u15_u6_n132 ) , .B1( u0_u15_u6_n133 ) , .ZN( u0_u15_u6_n134 ) , .A( u0_u15_u6_n158 ) );
  AOI21_X1 u0_u15_u6_U42 (.B1( u0_u15_u6_n131 ) , .ZN( u0_u15_u6_n135 ) , .A( u0_u15_u6_n144 ) , .B2( u0_u15_u6_n146 ) );
  INV_X1 u0_u15_u6_U43 (.A( u0_u15_u6_n111 ) , .ZN( u0_u15_u6_n158 ) );
  NAND2_X1 u0_u15_u6_U44 (.ZN( u0_u15_u6_n127 ) , .A1( u0_u15_u6_n91 ) , .A2( u0_u15_u6_n92 ) );
  NAND2_X1 u0_u15_u6_U45 (.ZN( u0_u15_u6_n129 ) , .A2( u0_u15_u6_n95 ) , .A1( u0_u15_u6_n96 ) );
  INV_X1 u0_u15_u6_U46 (.A( u0_u15_u6_n144 ) , .ZN( u0_u15_u6_n159 ) );
  NAND2_X1 u0_u15_u6_U47 (.ZN( u0_u15_u6_n145 ) , .A2( u0_u15_u6_n97 ) , .A1( u0_u15_u6_n98 ) );
  NAND2_X1 u0_u15_u6_U48 (.ZN( u0_u15_u6_n148 ) , .A2( u0_u15_u6_n92 ) , .A1( u0_u15_u6_n94 ) );
  NAND2_X1 u0_u15_u6_U49 (.ZN( u0_u15_u6_n108 ) , .A2( u0_u15_u6_n139 ) , .A1( u0_u15_u6_n144 ) );
  NAND2_X1 u0_u15_u6_U5 (.A2( u0_u15_u6_n143 ) , .ZN( u0_u15_u6_n152 ) , .A1( u0_u15_u6_n166 ) );
  NAND2_X1 u0_u15_u6_U50 (.ZN( u0_u15_u6_n121 ) , .A2( u0_u15_u6_n95 ) , .A1( u0_u15_u6_n97 ) );
  NAND2_X1 u0_u15_u6_U51 (.ZN( u0_u15_u6_n107 ) , .A2( u0_u15_u6_n92 ) , .A1( u0_u15_u6_n95 ) );
  AND2_X1 u0_u15_u6_U52 (.ZN( u0_u15_u6_n118 ) , .A2( u0_u15_u6_n91 ) , .A1( u0_u15_u6_n99 ) );
  NAND2_X1 u0_u15_u6_U53 (.ZN( u0_u15_u6_n147 ) , .A2( u0_u15_u6_n98 ) , .A1( u0_u15_u6_n99 ) );
  NAND2_X1 u0_u15_u6_U54 (.ZN( u0_u15_u6_n128 ) , .A1( u0_u15_u6_n94 ) , .A2( u0_u15_u6_n96 ) );
  NAND2_X1 u0_u15_u6_U55 (.ZN( u0_u15_u6_n119 ) , .A2( u0_u15_u6_n95 ) , .A1( u0_u15_u6_n99 ) );
  NAND2_X1 u0_u15_u6_U56 (.ZN( u0_u15_u6_n123 ) , .A2( u0_u15_u6_n91 ) , .A1( u0_u15_u6_n96 ) );
  NAND2_X1 u0_u15_u6_U57 (.ZN( u0_u15_u6_n100 ) , .A2( u0_u15_u6_n92 ) , .A1( u0_u15_u6_n98 ) );
  NAND2_X1 u0_u15_u6_U58 (.ZN( u0_u15_u6_n122 ) , .A1( u0_u15_u6_n94 ) , .A2( u0_u15_u6_n97 ) );
  INV_X1 u0_u15_u6_U59 (.A( u0_u15_u6_n139 ) , .ZN( u0_u15_u6_n160 ) );
  AOI22_X1 u0_u15_u6_U6 (.B2( u0_u15_u6_n101 ) , .A1( u0_u15_u6_n102 ) , .ZN( u0_u15_u6_n103 ) , .B1( u0_u15_u6_n160 ) , .A2( u0_u15_u6_n161 ) );
  NAND2_X1 u0_u15_u6_U60 (.ZN( u0_u15_u6_n113 ) , .A1( u0_u15_u6_n96 ) , .A2( u0_u15_u6_n98 ) );
  NOR2_X1 u0_u15_u6_U61 (.A2( u0_u15_X_40 ) , .A1( u0_u15_X_41 ) , .ZN( u0_u15_u6_n126 ) );
  NOR2_X1 u0_u15_u6_U62 (.A2( u0_u15_X_39 ) , .A1( u0_u15_X_42 ) , .ZN( u0_u15_u6_n92 ) );
  NOR2_X1 u0_u15_u6_U63 (.A2( u0_u15_X_39 ) , .A1( u0_u15_u6_n156 ) , .ZN( u0_u15_u6_n97 ) );
  NOR2_X1 u0_u15_u6_U64 (.A2( u0_u15_X_38 ) , .A1( u0_u15_u6_n165 ) , .ZN( u0_u15_u6_n95 ) );
  NOR2_X1 u0_u15_u6_U65 (.A2( u0_u15_X_41 ) , .ZN( u0_u15_u6_n111 ) , .A1( u0_u15_u6_n157 ) );
  NOR2_X1 u0_u15_u6_U66 (.A2( u0_u15_X_37 ) , .A1( u0_u15_u6_n162 ) , .ZN( u0_u15_u6_n94 ) );
  NOR2_X1 u0_u15_u6_U67 (.A2( u0_u15_X_37 ) , .A1( u0_u15_X_38 ) , .ZN( u0_u15_u6_n91 ) );
  NAND2_X1 u0_u15_u6_U68 (.A1( u0_u15_X_41 ) , .ZN( u0_u15_u6_n144 ) , .A2( u0_u15_u6_n157 ) );
  NAND2_X1 u0_u15_u6_U69 (.A2( u0_u15_X_40 ) , .A1( u0_u15_X_41 ) , .ZN( u0_u15_u6_n139 ) );
  NOR2_X1 u0_u15_u6_U7 (.A1( u0_u15_u6_n118 ) , .ZN( u0_u15_u6_n143 ) , .A2( u0_u15_u6_n168 ) );
  AND2_X1 u0_u15_u6_U70 (.A1( u0_u15_X_39 ) , .A2( u0_u15_u6_n156 ) , .ZN( u0_u15_u6_n96 ) );
  AND2_X1 u0_u15_u6_U71 (.A1( u0_u15_X_39 ) , .A2( u0_u15_X_42 ) , .ZN( u0_u15_u6_n99 ) );
  INV_X1 u0_u15_u6_U72 (.A( u0_u15_X_40 ) , .ZN( u0_u15_u6_n157 ) );
  INV_X1 u0_u15_u6_U73 (.A( u0_u15_X_37 ) , .ZN( u0_u15_u6_n165 ) );
  INV_X1 u0_u15_u6_U74 (.A( u0_u15_X_38 ) , .ZN( u0_u15_u6_n162 ) );
  INV_X1 u0_u15_u6_U75 (.A( u0_u15_X_42 ) , .ZN( u0_u15_u6_n156 ) );
  NAND4_X1 u0_u15_u6_U76 (.ZN( u0_out15_12 ) , .A4( u0_u15_u6_n114 ) , .A3( u0_u15_u6_n115 ) , .A2( u0_u15_u6_n116 ) , .A1( u0_u15_u6_n117 ) );
  OAI22_X1 u0_u15_u6_U77 (.B2( u0_u15_u6_n111 ) , .ZN( u0_u15_u6_n116 ) , .B1( u0_u15_u6_n126 ) , .A2( u0_u15_u6_n164 ) , .A1( u0_u15_u6_n167 ) );
  OAI21_X1 u0_u15_u6_U78 (.A( u0_u15_u6_n108 ) , .ZN( u0_u15_u6_n117 ) , .B2( u0_u15_u6_n141 ) , .B1( u0_u15_u6_n163 ) );
  NAND4_X1 u0_u15_u6_U79 (.ZN( u0_out15_32 ) , .A4( u0_u15_u6_n103 ) , .A3( u0_u15_u6_n104 ) , .A2( u0_u15_u6_n105 ) , .A1( u0_u15_u6_n106 ) );
  AOI21_X1 u0_u15_u6_U8 (.B1( u0_u15_u6_n107 ) , .B2( u0_u15_u6_n132 ) , .A( u0_u15_u6_n158 ) , .ZN( u0_u15_u6_n88 ) );
  AOI22_X1 u0_u15_u6_U80 (.ZN( u0_u15_u6_n105 ) , .A2( u0_u15_u6_n108 ) , .A1( u0_u15_u6_n118 ) , .B2( u0_u15_u6_n126 ) , .B1( u0_u15_u6_n171 ) );
  AOI22_X1 u0_u15_u6_U81 (.ZN( u0_u15_u6_n104 ) , .A1( u0_u15_u6_n111 ) , .B1( u0_u15_u6_n124 ) , .B2( u0_u15_u6_n151 ) , .A2( u0_u15_u6_n93 ) );
  OAI211_X1 u0_u15_u6_U82 (.ZN( u0_out15_22 ) , .B( u0_u15_u6_n137 ) , .A( u0_u15_u6_n138 ) , .C2( u0_u15_u6_n139 ) , .C1( u0_u15_u6_n140 ) );
  AOI22_X1 u0_u15_u6_U83 (.B1( u0_u15_u6_n124 ) , .A2( u0_u15_u6_n125 ) , .A1( u0_u15_u6_n126 ) , .ZN( u0_u15_u6_n138 ) , .B2( u0_u15_u6_n161 ) );
  AND4_X1 u0_u15_u6_U84 (.A3( u0_u15_u6_n119 ) , .A1( u0_u15_u6_n120 ) , .A4( u0_u15_u6_n129 ) , .ZN( u0_u15_u6_n140 ) , .A2( u0_u15_u6_n143 ) );
  OAI211_X1 u0_u15_u6_U85 (.ZN( u0_out15_7 ) , .B( u0_u15_u6_n153 ) , .C2( u0_u15_u6_n154 ) , .C1( u0_u15_u6_n155 ) , .A( u0_u15_u6_n174 ) );
  NOR3_X1 u0_u15_u6_U86 (.A1( u0_u15_u6_n141 ) , .ZN( u0_u15_u6_n154 ) , .A3( u0_u15_u6_n164 ) , .A2( u0_u15_u6_n171 ) );
  AOI211_X1 u0_u15_u6_U87 (.B( u0_u15_u6_n149 ) , .A( u0_u15_u6_n150 ) , .C2( u0_u15_u6_n151 ) , .C1( u0_u15_u6_n152 ) , .ZN( u0_u15_u6_n153 ) );
  NAND3_X1 u0_u15_u6_U88 (.A2( u0_u15_u6_n123 ) , .ZN( u0_u15_u6_n125 ) , .A1( u0_u15_u6_n130 ) , .A3( u0_u15_u6_n131 ) );
  NAND3_X1 u0_u15_u6_U89 (.A3( u0_u15_u6_n133 ) , .ZN( u0_u15_u6_n141 ) , .A1( u0_u15_u6_n145 ) , .A2( u0_u15_u6_n148 ) );
  AOI21_X1 u0_u15_u6_U9 (.B2( u0_u15_u6_n147 ) , .B1( u0_u15_u6_n148 ) , .ZN( u0_u15_u6_n149 ) , .A( u0_u15_u6_n158 ) );
  NAND3_X1 u0_u15_u6_U90 (.ZN( u0_u15_u6_n101 ) , .A3( u0_u15_u6_n107 ) , .A2( u0_u15_u6_n121 ) , .A1( u0_u15_u6_n127 ) );
  NAND3_X1 u0_u15_u6_U91 (.ZN( u0_u15_u6_n102 ) , .A3( u0_u15_u6_n130 ) , .A2( u0_u15_u6_n145 ) , .A1( u0_u15_u6_n166 ) );
  NAND3_X1 u0_u15_u6_U92 (.A3( u0_u15_u6_n113 ) , .A1( u0_u15_u6_n119 ) , .A2( u0_u15_u6_n123 ) , .ZN( u0_u15_u6_n93 ) );
  NAND3_X1 u0_u15_u6_U93 (.ZN( u0_u15_u6_n142 ) , .A2( u0_u15_u6_n172 ) , .A3( u0_u15_u6_n89 ) , .A1( u0_u15_u6_n90 ) );
  XOR2_X1 u0_u4_U1 (.B( u0_K5_9 ) , .A( u0_R3_6 ) , .Z( u0_u4_X_9 ) );
  XOR2_X1 u0_u4_U2 (.B( u0_K5_8 ) , .A( u0_R3_5 ) , .Z( u0_u4_X_8 ) );
  XOR2_X1 u0_u4_U3 (.B( u0_K5_7 ) , .A( u0_R3_4 ) , .Z( u0_u4_X_7 ) );
  XOR2_X1 u0_u4_U33 (.B( u0_K5_24 ) , .A( u0_R3_17 ) , .Z( u0_u4_X_24 ) );
  XOR2_X1 u0_u4_U34 (.B( u0_K5_23 ) , .A( u0_R3_16 ) , .Z( u0_u4_X_23 ) );
  XOR2_X1 u0_u4_U35 (.B( u0_K5_22 ) , .A( u0_R3_15 ) , .Z( u0_u4_X_22 ) );
  XOR2_X1 u0_u4_U36 (.B( u0_K5_21 ) , .A( u0_R3_14 ) , .Z( u0_u4_X_21 ) );
  XOR2_X1 u0_u4_U37 (.B( u0_K5_20 ) , .A( u0_R3_13 ) , .Z( u0_u4_X_20 ) );
  XOR2_X1 u0_u4_U39 (.B( u0_K5_19 ) , .A( u0_R3_12 ) , .Z( u0_u4_X_19 ) );
  XOR2_X1 u0_u4_U40 (.B( u0_K5_18 ) , .A( u0_R3_13 ) , .Z( u0_u4_X_18 ) );
  XOR2_X1 u0_u4_U41 (.B( u0_K5_17 ) , .A( u0_R3_12 ) , .Z( u0_u4_X_17 ) );
  XOR2_X1 u0_u4_U42 (.B( u0_K5_16 ) , .A( u0_R3_11 ) , .Z( u0_u4_X_16 ) );
  XOR2_X1 u0_u4_U43 (.B( u0_K5_15 ) , .A( u0_R3_10 ) , .Z( u0_u4_X_15 ) );
  XOR2_X1 u0_u4_U44 (.B( u0_K5_14 ) , .A( u0_R3_9 ) , .Z( u0_u4_X_14 ) );
  XOR2_X1 u0_u4_U45 (.B( u0_K5_13 ) , .A( u0_R3_8 ) , .Z( u0_u4_X_13 ) );
  XOR2_X1 u0_u4_U46 (.B( u0_K5_12 ) , .A( u0_R3_9 ) , .Z( u0_u4_X_12 ) );
  XOR2_X1 u0_u4_U47 (.B( u0_K5_11 ) , .A( u0_R3_8 ) , .Z( u0_u4_X_11 ) );
  XOR2_X1 u0_u4_U48 (.B( u0_K5_10 ) , .A( u0_R3_7 ) , .Z( u0_u4_X_10 ) );
  NOR2_X1 u0_u4_u1_U10 (.A1( u0_u4_u1_n112 ) , .A2( u0_u4_u1_n116 ) , .ZN( u0_u4_u1_n118 ) );
  NAND3_X1 u0_u4_u1_U100 (.ZN( u0_u4_u1_n113 ) , .A1( u0_u4_u1_n120 ) , .A3( u0_u4_u1_n133 ) , .A2( u0_u4_u1_n155 ) );
  OAI21_X1 u0_u4_u1_U11 (.ZN( u0_u4_u1_n101 ) , .B1( u0_u4_u1_n141 ) , .A( u0_u4_u1_n146 ) , .B2( u0_u4_u1_n183 ) );
  AOI21_X1 u0_u4_u1_U12 (.B2( u0_u4_u1_n155 ) , .B1( u0_u4_u1_n156 ) , .ZN( u0_u4_u1_n157 ) , .A( u0_u4_u1_n174 ) );
  NAND2_X1 u0_u4_u1_U13 (.ZN( u0_u4_u1_n140 ) , .A2( u0_u4_u1_n150 ) , .A1( u0_u4_u1_n155 ) );
  NAND2_X1 u0_u4_u1_U14 (.A1( u0_u4_u1_n131 ) , .ZN( u0_u4_u1_n147 ) , .A2( u0_u4_u1_n153 ) );
  INV_X1 u0_u4_u1_U15 (.A( u0_u4_u1_n139 ) , .ZN( u0_u4_u1_n174 ) );
  OR4_X1 u0_u4_u1_U16 (.A4( u0_u4_u1_n106 ) , .A3( u0_u4_u1_n107 ) , .ZN( u0_u4_u1_n108 ) , .A1( u0_u4_u1_n117 ) , .A2( u0_u4_u1_n184 ) );
  AOI21_X1 u0_u4_u1_U17 (.ZN( u0_u4_u1_n106 ) , .A( u0_u4_u1_n112 ) , .B1( u0_u4_u1_n154 ) , .B2( u0_u4_u1_n156 ) );
  AOI21_X1 u0_u4_u1_U18 (.ZN( u0_u4_u1_n107 ) , .B1( u0_u4_u1_n134 ) , .B2( u0_u4_u1_n149 ) , .A( u0_u4_u1_n174 ) );
  INV_X1 u0_u4_u1_U19 (.A( u0_u4_u1_n101 ) , .ZN( u0_u4_u1_n184 ) );
  INV_X1 u0_u4_u1_U20 (.A( u0_u4_u1_n112 ) , .ZN( u0_u4_u1_n171 ) );
  NAND2_X1 u0_u4_u1_U21 (.ZN( u0_u4_u1_n141 ) , .A1( u0_u4_u1_n153 ) , .A2( u0_u4_u1_n156 ) );
  AND2_X1 u0_u4_u1_U22 (.A1( u0_u4_u1_n123 ) , .ZN( u0_u4_u1_n134 ) , .A2( u0_u4_u1_n161 ) );
  NAND2_X1 u0_u4_u1_U23 (.A2( u0_u4_u1_n115 ) , .A1( u0_u4_u1_n116 ) , .ZN( u0_u4_u1_n148 ) );
  NAND2_X1 u0_u4_u1_U24 (.A2( u0_u4_u1_n133 ) , .A1( u0_u4_u1_n135 ) , .ZN( u0_u4_u1_n159 ) );
  NAND2_X1 u0_u4_u1_U25 (.A2( u0_u4_u1_n115 ) , .A1( u0_u4_u1_n120 ) , .ZN( u0_u4_u1_n132 ) );
  INV_X1 u0_u4_u1_U26 (.A( u0_u4_u1_n154 ) , .ZN( u0_u4_u1_n178 ) );
  INV_X1 u0_u4_u1_U27 (.A( u0_u4_u1_n151 ) , .ZN( u0_u4_u1_n183 ) );
  AND2_X1 u0_u4_u1_U28 (.A1( u0_u4_u1_n129 ) , .A2( u0_u4_u1_n133 ) , .ZN( u0_u4_u1_n149 ) );
  INV_X1 u0_u4_u1_U29 (.A( u0_u4_u1_n131 ) , .ZN( u0_u4_u1_n180 ) );
  INV_X1 u0_u4_u1_U3 (.A( u0_u4_u1_n159 ) , .ZN( u0_u4_u1_n182 ) );
  OAI221_X1 u0_u4_u1_U30 (.A( u0_u4_u1_n119 ) , .C2( u0_u4_u1_n129 ) , .ZN( u0_u4_u1_n138 ) , .B2( u0_u4_u1_n152 ) , .C1( u0_u4_u1_n174 ) , .B1( u0_u4_u1_n187 ) );
  INV_X1 u0_u4_u1_U31 (.A( u0_u4_u1_n148 ) , .ZN( u0_u4_u1_n187 ) );
  AOI211_X1 u0_u4_u1_U32 (.B( u0_u4_u1_n117 ) , .A( u0_u4_u1_n118 ) , .ZN( u0_u4_u1_n119 ) , .C2( u0_u4_u1_n146 ) , .C1( u0_u4_u1_n159 ) );
  NOR2_X1 u0_u4_u1_U33 (.A1( u0_u4_u1_n168 ) , .A2( u0_u4_u1_n176 ) , .ZN( u0_u4_u1_n98 ) );
  AOI211_X1 u0_u4_u1_U34 (.B( u0_u4_u1_n162 ) , .A( u0_u4_u1_n163 ) , .C2( u0_u4_u1_n164 ) , .ZN( u0_u4_u1_n165 ) , .C1( u0_u4_u1_n171 ) );
  AOI21_X1 u0_u4_u1_U35 (.A( u0_u4_u1_n160 ) , .B2( u0_u4_u1_n161 ) , .ZN( u0_u4_u1_n162 ) , .B1( u0_u4_u1_n182 ) );
  OR2_X1 u0_u4_u1_U36 (.A2( u0_u4_u1_n157 ) , .A1( u0_u4_u1_n158 ) , .ZN( u0_u4_u1_n163 ) );
  NAND2_X1 u0_u4_u1_U37 (.A1( u0_u4_u1_n128 ) , .ZN( u0_u4_u1_n146 ) , .A2( u0_u4_u1_n160 ) );
  NAND2_X1 u0_u4_u1_U38 (.A2( u0_u4_u1_n112 ) , .ZN( u0_u4_u1_n139 ) , .A1( u0_u4_u1_n152 ) );
  NAND2_X1 u0_u4_u1_U39 (.A1( u0_u4_u1_n105 ) , .ZN( u0_u4_u1_n156 ) , .A2( u0_u4_u1_n99 ) );
  AOI221_X1 u0_u4_u1_U4 (.A( u0_u4_u1_n138 ) , .C2( u0_u4_u1_n139 ) , .C1( u0_u4_u1_n140 ) , .B2( u0_u4_u1_n141 ) , .ZN( u0_u4_u1_n142 ) , .B1( u0_u4_u1_n175 ) );
  AOI221_X1 u0_u4_u1_U40 (.B1( u0_u4_u1_n140 ) , .ZN( u0_u4_u1_n167 ) , .B2( u0_u4_u1_n172 ) , .C2( u0_u4_u1_n175 ) , .C1( u0_u4_u1_n178 ) , .A( u0_u4_u1_n188 ) );
  INV_X1 u0_u4_u1_U41 (.ZN( u0_u4_u1_n188 ) , .A( u0_u4_u1_n97 ) );
  AOI211_X1 u0_u4_u1_U42 (.A( u0_u4_u1_n118 ) , .C1( u0_u4_u1_n132 ) , .C2( u0_u4_u1_n139 ) , .B( u0_u4_u1_n96 ) , .ZN( u0_u4_u1_n97 ) );
  AOI21_X1 u0_u4_u1_U43 (.B2( u0_u4_u1_n121 ) , .B1( u0_u4_u1_n135 ) , .A( u0_u4_u1_n152 ) , .ZN( u0_u4_u1_n96 ) );
  NOR2_X1 u0_u4_u1_U44 (.ZN( u0_u4_u1_n117 ) , .A1( u0_u4_u1_n121 ) , .A2( u0_u4_u1_n160 ) );
  OAI21_X1 u0_u4_u1_U45 (.B2( u0_u4_u1_n123 ) , .ZN( u0_u4_u1_n145 ) , .B1( u0_u4_u1_n160 ) , .A( u0_u4_u1_n185 ) );
  INV_X1 u0_u4_u1_U46 (.A( u0_u4_u1_n122 ) , .ZN( u0_u4_u1_n185 ) );
  AOI21_X1 u0_u4_u1_U47 (.B2( u0_u4_u1_n120 ) , .B1( u0_u4_u1_n121 ) , .ZN( u0_u4_u1_n122 ) , .A( u0_u4_u1_n128 ) );
  AOI21_X1 u0_u4_u1_U48 (.A( u0_u4_u1_n128 ) , .B2( u0_u4_u1_n129 ) , .ZN( u0_u4_u1_n130 ) , .B1( u0_u4_u1_n150 ) );
  NAND2_X1 u0_u4_u1_U49 (.ZN( u0_u4_u1_n112 ) , .A1( u0_u4_u1_n169 ) , .A2( u0_u4_u1_n170 ) );
  AOI211_X1 u0_u4_u1_U5 (.ZN( u0_u4_u1_n124 ) , .A( u0_u4_u1_n138 ) , .C2( u0_u4_u1_n139 ) , .B( u0_u4_u1_n145 ) , .C1( u0_u4_u1_n147 ) );
  NAND2_X1 u0_u4_u1_U50 (.ZN( u0_u4_u1_n129 ) , .A2( u0_u4_u1_n95 ) , .A1( u0_u4_u1_n98 ) );
  NAND2_X1 u0_u4_u1_U51 (.A1( u0_u4_u1_n102 ) , .ZN( u0_u4_u1_n154 ) , .A2( u0_u4_u1_n99 ) );
  NAND2_X1 u0_u4_u1_U52 (.A2( u0_u4_u1_n100 ) , .ZN( u0_u4_u1_n135 ) , .A1( u0_u4_u1_n99 ) );
  AOI21_X1 u0_u4_u1_U53 (.A( u0_u4_u1_n152 ) , .B2( u0_u4_u1_n153 ) , .B1( u0_u4_u1_n154 ) , .ZN( u0_u4_u1_n158 ) );
  INV_X1 u0_u4_u1_U54 (.A( u0_u4_u1_n160 ) , .ZN( u0_u4_u1_n175 ) );
  NAND2_X1 u0_u4_u1_U55 (.A1( u0_u4_u1_n100 ) , .ZN( u0_u4_u1_n116 ) , .A2( u0_u4_u1_n95 ) );
  NAND2_X1 u0_u4_u1_U56 (.A1( u0_u4_u1_n102 ) , .ZN( u0_u4_u1_n131 ) , .A2( u0_u4_u1_n95 ) );
  NAND2_X1 u0_u4_u1_U57 (.A2( u0_u4_u1_n104 ) , .ZN( u0_u4_u1_n121 ) , .A1( u0_u4_u1_n98 ) );
  NAND2_X1 u0_u4_u1_U58 (.A1( u0_u4_u1_n103 ) , .ZN( u0_u4_u1_n153 ) , .A2( u0_u4_u1_n98 ) );
  NAND2_X1 u0_u4_u1_U59 (.A2( u0_u4_u1_n104 ) , .A1( u0_u4_u1_n105 ) , .ZN( u0_u4_u1_n133 ) );
  AOI22_X1 u0_u4_u1_U6 (.B2( u0_u4_u1_n113 ) , .A2( u0_u4_u1_n114 ) , .ZN( u0_u4_u1_n125 ) , .A1( u0_u4_u1_n171 ) , .B1( u0_u4_u1_n173 ) );
  NAND2_X1 u0_u4_u1_U60 (.ZN( u0_u4_u1_n150 ) , .A2( u0_u4_u1_n98 ) , .A1( u0_u4_u1_n99 ) );
  NAND2_X1 u0_u4_u1_U61 (.A1( u0_u4_u1_n105 ) , .ZN( u0_u4_u1_n155 ) , .A2( u0_u4_u1_n95 ) );
  OAI21_X1 u0_u4_u1_U62 (.ZN( u0_u4_u1_n109 ) , .B1( u0_u4_u1_n129 ) , .B2( u0_u4_u1_n160 ) , .A( u0_u4_u1_n167 ) );
  NAND2_X1 u0_u4_u1_U63 (.A2( u0_u4_u1_n100 ) , .A1( u0_u4_u1_n103 ) , .ZN( u0_u4_u1_n120 ) );
  NAND2_X1 u0_u4_u1_U64 (.A1( u0_u4_u1_n102 ) , .A2( u0_u4_u1_n104 ) , .ZN( u0_u4_u1_n115 ) );
  NAND2_X1 u0_u4_u1_U65 (.A2( u0_u4_u1_n100 ) , .A1( u0_u4_u1_n104 ) , .ZN( u0_u4_u1_n151 ) );
  NAND2_X1 u0_u4_u1_U66 (.A2( u0_u4_u1_n103 ) , .A1( u0_u4_u1_n105 ) , .ZN( u0_u4_u1_n161 ) );
  INV_X1 u0_u4_u1_U67 (.A( u0_u4_u1_n152 ) , .ZN( u0_u4_u1_n173 ) );
  INV_X1 u0_u4_u1_U68 (.A( u0_u4_u1_n128 ) , .ZN( u0_u4_u1_n172 ) );
  NAND2_X1 u0_u4_u1_U69 (.A2( u0_u4_u1_n102 ) , .A1( u0_u4_u1_n103 ) , .ZN( u0_u4_u1_n123 ) );
  NAND2_X1 u0_u4_u1_U7 (.ZN( u0_u4_u1_n114 ) , .A1( u0_u4_u1_n134 ) , .A2( u0_u4_u1_n156 ) );
  NOR2_X1 u0_u4_u1_U70 (.A2( u0_u4_X_7 ) , .A1( u0_u4_X_8 ) , .ZN( u0_u4_u1_n95 ) );
  NOR2_X1 u0_u4_u1_U71 (.A1( u0_u4_X_12 ) , .A2( u0_u4_X_9 ) , .ZN( u0_u4_u1_n100 ) );
  NOR2_X1 u0_u4_u1_U72 (.A2( u0_u4_X_8 ) , .A1( u0_u4_u1_n177 ) , .ZN( u0_u4_u1_n99 ) );
  NOR2_X1 u0_u4_u1_U73 (.A2( u0_u4_X_12 ) , .ZN( u0_u4_u1_n102 ) , .A1( u0_u4_u1_n176 ) );
  NOR2_X1 u0_u4_u1_U74 (.A2( u0_u4_X_9 ) , .ZN( u0_u4_u1_n105 ) , .A1( u0_u4_u1_n168 ) );
  NAND2_X1 u0_u4_u1_U75 (.A1( u0_u4_X_10 ) , .ZN( u0_u4_u1_n160 ) , .A2( u0_u4_u1_n169 ) );
  NAND2_X1 u0_u4_u1_U76 (.A2( u0_u4_X_10 ) , .A1( u0_u4_X_11 ) , .ZN( u0_u4_u1_n152 ) );
  NAND2_X1 u0_u4_u1_U77 (.A1( u0_u4_X_11 ) , .ZN( u0_u4_u1_n128 ) , .A2( u0_u4_u1_n170 ) );
  AND2_X1 u0_u4_u1_U78 (.A2( u0_u4_X_7 ) , .A1( u0_u4_X_8 ) , .ZN( u0_u4_u1_n104 ) );
  AND2_X1 u0_u4_u1_U79 (.A1( u0_u4_X_8 ) , .ZN( u0_u4_u1_n103 ) , .A2( u0_u4_u1_n177 ) );
  AOI22_X1 u0_u4_u1_U8 (.B2( u0_u4_u1_n136 ) , .A2( u0_u4_u1_n137 ) , .ZN( u0_u4_u1_n143 ) , .A1( u0_u4_u1_n171 ) , .B1( u0_u4_u1_n173 ) );
  INV_X1 u0_u4_u1_U80 (.A( u0_u4_X_10 ) , .ZN( u0_u4_u1_n170 ) );
  INV_X1 u0_u4_u1_U81 (.A( u0_u4_X_9 ) , .ZN( u0_u4_u1_n176 ) );
  INV_X1 u0_u4_u1_U82 (.A( u0_u4_X_11 ) , .ZN( u0_u4_u1_n169 ) );
  INV_X1 u0_u4_u1_U83 (.A( u0_u4_X_12 ) , .ZN( u0_u4_u1_n168 ) );
  INV_X1 u0_u4_u1_U84 (.A( u0_u4_X_7 ) , .ZN( u0_u4_u1_n177 ) );
  NAND4_X1 u0_u4_u1_U85 (.ZN( u0_out4_28 ) , .A4( u0_u4_u1_n124 ) , .A3( u0_u4_u1_n125 ) , .A2( u0_u4_u1_n126 ) , .A1( u0_u4_u1_n127 ) );
  OAI21_X1 u0_u4_u1_U86 (.ZN( u0_u4_u1_n127 ) , .B2( u0_u4_u1_n139 ) , .B1( u0_u4_u1_n175 ) , .A( u0_u4_u1_n183 ) );
  OAI21_X1 u0_u4_u1_U87 (.ZN( u0_u4_u1_n126 ) , .B2( u0_u4_u1_n140 ) , .A( u0_u4_u1_n146 ) , .B1( u0_u4_u1_n178 ) );
  NAND4_X1 u0_u4_u1_U88 (.ZN( u0_out4_18 ) , .A4( u0_u4_u1_n165 ) , .A3( u0_u4_u1_n166 ) , .A1( u0_u4_u1_n167 ) , .A2( u0_u4_u1_n186 ) );
  AOI22_X1 u0_u4_u1_U89 (.B2( u0_u4_u1_n146 ) , .B1( u0_u4_u1_n147 ) , .A2( u0_u4_u1_n148 ) , .ZN( u0_u4_u1_n166 ) , .A1( u0_u4_u1_n172 ) );
  INV_X1 u0_u4_u1_U9 (.A( u0_u4_u1_n147 ) , .ZN( u0_u4_u1_n181 ) );
  INV_X1 u0_u4_u1_U90 (.A( u0_u4_u1_n145 ) , .ZN( u0_u4_u1_n186 ) );
  NAND4_X1 u0_u4_u1_U91 (.ZN( u0_out4_2 ) , .A4( u0_u4_u1_n142 ) , .A3( u0_u4_u1_n143 ) , .A2( u0_u4_u1_n144 ) , .A1( u0_u4_u1_n179 ) );
  OAI21_X1 u0_u4_u1_U92 (.B2( u0_u4_u1_n132 ) , .ZN( u0_u4_u1_n144 ) , .A( u0_u4_u1_n146 ) , .B1( u0_u4_u1_n180 ) );
  INV_X1 u0_u4_u1_U93 (.A( u0_u4_u1_n130 ) , .ZN( u0_u4_u1_n179 ) );
  OR4_X1 u0_u4_u1_U94 (.ZN( u0_out4_13 ) , .A4( u0_u4_u1_n108 ) , .A3( u0_u4_u1_n109 ) , .A2( u0_u4_u1_n110 ) , .A1( u0_u4_u1_n111 ) );
  AOI21_X1 u0_u4_u1_U95 (.ZN( u0_u4_u1_n111 ) , .A( u0_u4_u1_n128 ) , .B2( u0_u4_u1_n131 ) , .B1( u0_u4_u1_n135 ) );
  AOI21_X1 u0_u4_u1_U96 (.ZN( u0_u4_u1_n110 ) , .A( u0_u4_u1_n116 ) , .B1( u0_u4_u1_n152 ) , .B2( u0_u4_u1_n160 ) );
  NAND3_X1 u0_u4_u1_U97 (.A3( u0_u4_u1_n149 ) , .A2( u0_u4_u1_n150 ) , .A1( u0_u4_u1_n151 ) , .ZN( u0_u4_u1_n164 ) );
  NAND3_X1 u0_u4_u1_U98 (.A3( u0_u4_u1_n134 ) , .A2( u0_u4_u1_n135 ) , .ZN( u0_u4_u1_n136 ) , .A1( u0_u4_u1_n151 ) );
  NAND3_X1 u0_u4_u1_U99 (.A1( u0_u4_u1_n133 ) , .ZN( u0_u4_u1_n137 ) , .A2( u0_u4_u1_n154 ) , .A3( u0_u4_u1_n181 ) );
  OAI22_X1 u0_u4_u2_U10 (.ZN( u0_u4_u2_n109 ) , .A2( u0_u4_u2_n113 ) , .B2( u0_u4_u2_n133 ) , .B1( u0_u4_u2_n167 ) , .A1( u0_u4_u2_n168 ) );
  NAND3_X1 u0_u4_u2_U100 (.A2( u0_u4_u2_n100 ) , .A1( u0_u4_u2_n104 ) , .A3( u0_u4_u2_n138 ) , .ZN( u0_u4_u2_n98 ) );
  OAI22_X1 u0_u4_u2_U11 (.B1( u0_u4_u2_n151 ) , .A2( u0_u4_u2_n152 ) , .A1( u0_u4_u2_n153 ) , .ZN( u0_u4_u2_n160 ) , .B2( u0_u4_u2_n168 ) );
  NOR3_X1 u0_u4_u2_U12 (.A1( u0_u4_u2_n150 ) , .ZN( u0_u4_u2_n151 ) , .A3( u0_u4_u2_n175 ) , .A2( u0_u4_u2_n188 ) );
  AOI21_X1 u0_u4_u2_U13 (.ZN( u0_u4_u2_n144 ) , .B2( u0_u4_u2_n155 ) , .A( u0_u4_u2_n172 ) , .B1( u0_u4_u2_n185 ) );
  AOI21_X1 u0_u4_u2_U14 (.B2( u0_u4_u2_n143 ) , .ZN( u0_u4_u2_n145 ) , .B1( u0_u4_u2_n152 ) , .A( u0_u4_u2_n171 ) );
  AOI21_X1 u0_u4_u2_U15 (.B2( u0_u4_u2_n120 ) , .B1( u0_u4_u2_n121 ) , .ZN( u0_u4_u2_n126 ) , .A( u0_u4_u2_n167 ) );
  INV_X1 u0_u4_u2_U16 (.A( u0_u4_u2_n156 ) , .ZN( u0_u4_u2_n171 ) );
  INV_X1 u0_u4_u2_U17 (.A( u0_u4_u2_n120 ) , .ZN( u0_u4_u2_n188 ) );
  NAND2_X1 u0_u4_u2_U18 (.A2( u0_u4_u2_n122 ) , .ZN( u0_u4_u2_n150 ) , .A1( u0_u4_u2_n152 ) );
  INV_X1 u0_u4_u2_U19 (.A( u0_u4_u2_n153 ) , .ZN( u0_u4_u2_n170 ) );
  INV_X1 u0_u4_u2_U20 (.A( u0_u4_u2_n137 ) , .ZN( u0_u4_u2_n173 ) );
  NAND2_X1 u0_u4_u2_U21 (.A1( u0_u4_u2_n132 ) , .A2( u0_u4_u2_n139 ) , .ZN( u0_u4_u2_n157 ) );
  INV_X1 u0_u4_u2_U22 (.A( u0_u4_u2_n113 ) , .ZN( u0_u4_u2_n178 ) );
  INV_X1 u0_u4_u2_U23 (.A( u0_u4_u2_n139 ) , .ZN( u0_u4_u2_n175 ) );
  INV_X1 u0_u4_u2_U24 (.A( u0_u4_u2_n155 ) , .ZN( u0_u4_u2_n181 ) );
  INV_X1 u0_u4_u2_U25 (.A( u0_u4_u2_n119 ) , .ZN( u0_u4_u2_n177 ) );
  INV_X1 u0_u4_u2_U26 (.A( u0_u4_u2_n116 ) , .ZN( u0_u4_u2_n180 ) );
  INV_X1 u0_u4_u2_U27 (.A( u0_u4_u2_n131 ) , .ZN( u0_u4_u2_n179 ) );
  INV_X1 u0_u4_u2_U28 (.A( u0_u4_u2_n154 ) , .ZN( u0_u4_u2_n176 ) );
  NAND2_X1 u0_u4_u2_U29 (.A2( u0_u4_u2_n116 ) , .A1( u0_u4_u2_n117 ) , .ZN( u0_u4_u2_n118 ) );
  NOR2_X1 u0_u4_u2_U3 (.ZN( u0_u4_u2_n121 ) , .A2( u0_u4_u2_n177 ) , .A1( u0_u4_u2_n180 ) );
  INV_X1 u0_u4_u2_U30 (.A( u0_u4_u2_n132 ) , .ZN( u0_u4_u2_n182 ) );
  INV_X1 u0_u4_u2_U31 (.A( u0_u4_u2_n158 ) , .ZN( u0_u4_u2_n183 ) );
  OAI21_X1 u0_u4_u2_U32 (.A( u0_u4_u2_n156 ) , .B1( u0_u4_u2_n157 ) , .ZN( u0_u4_u2_n158 ) , .B2( u0_u4_u2_n179 ) );
  NOR2_X1 u0_u4_u2_U33 (.ZN( u0_u4_u2_n156 ) , .A1( u0_u4_u2_n166 ) , .A2( u0_u4_u2_n169 ) );
  NOR2_X1 u0_u4_u2_U34 (.A2( u0_u4_u2_n114 ) , .ZN( u0_u4_u2_n137 ) , .A1( u0_u4_u2_n140 ) );
  NOR2_X1 u0_u4_u2_U35 (.A2( u0_u4_u2_n138 ) , .ZN( u0_u4_u2_n153 ) , .A1( u0_u4_u2_n156 ) );
  AOI211_X1 u0_u4_u2_U36 (.ZN( u0_u4_u2_n130 ) , .C1( u0_u4_u2_n138 ) , .C2( u0_u4_u2_n179 ) , .B( u0_u4_u2_n96 ) , .A( u0_u4_u2_n97 ) );
  OAI22_X1 u0_u4_u2_U37 (.B1( u0_u4_u2_n133 ) , .A2( u0_u4_u2_n137 ) , .A1( u0_u4_u2_n152 ) , .B2( u0_u4_u2_n168 ) , .ZN( u0_u4_u2_n97 ) );
  OAI221_X1 u0_u4_u2_U38 (.B1( u0_u4_u2_n113 ) , .C1( u0_u4_u2_n132 ) , .A( u0_u4_u2_n149 ) , .B2( u0_u4_u2_n171 ) , .C2( u0_u4_u2_n172 ) , .ZN( u0_u4_u2_n96 ) );
  OAI221_X1 u0_u4_u2_U39 (.A( u0_u4_u2_n115 ) , .C2( u0_u4_u2_n123 ) , .B2( u0_u4_u2_n143 ) , .B1( u0_u4_u2_n153 ) , .ZN( u0_u4_u2_n163 ) , .C1( u0_u4_u2_n168 ) );
  INV_X1 u0_u4_u2_U4 (.A( u0_u4_u2_n134 ) , .ZN( u0_u4_u2_n185 ) );
  OAI21_X1 u0_u4_u2_U40 (.A( u0_u4_u2_n114 ) , .ZN( u0_u4_u2_n115 ) , .B1( u0_u4_u2_n176 ) , .B2( u0_u4_u2_n178 ) );
  OAI221_X1 u0_u4_u2_U41 (.A( u0_u4_u2_n135 ) , .B2( u0_u4_u2_n136 ) , .B1( u0_u4_u2_n137 ) , .ZN( u0_u4_u2_n162 ) , .C2( u0_u4_u2_n167 ) , .C1( u0_u4_u2_n185 ) );
  AND3_X1 u0_u4_u2_U42 (.A3( u0_u4_u2_n131 ) , .A2( u0_u4_u2_n132 ) , .A1( u0_u4_u2_n133 ) , .ZN( u0_u4_u2_n136 ) );
  AOI22_X1 u0_u4_u2_U43 (.ZN( u0_u4_u2_n135 ) , .B1( u0_u4_u2_n140 ) , .A1( u0_u4_u2_n156 ) , .B2( u0_u4_u2_n180 ) , .A2( u0_u4_u2_n188 ) );
  AOI21_X1 u0_u4_u2_U44 (.ZN( u0_u4_u2_n149 ) , .B1( u0_u4_u2_n173 ) , .B2( u0_u4_u2_n188 ) , .A( u0_u4_u2_n95 ) );
  AND3_X1 u0_u4_u2_U45 (.A2( u0_u4_u2_n100 ) , .A1( u0_u4_u2_n104 ) , .A3( u0_u4_u2_n156 ) , .ZN( u0_u4_u2_n95 ) );
  OAI21_X1 u0_u4_u2_U46 (.A( u0_u4_u2_n101 ) , .B2( u0_u4_u2_n121 ) , .B1( u0_u4_u2_n153 ) , .ZN( u0_u4_u2_n164 ) );
  NAND2_X1 u0_u4_u2_U47 (.A2( u0_u4_u2_n100 ) , .A1( u0_u4_u2_n107 ) , .ZN( u0_u4_u2_n155 ) );
  NAND2_X1 u0_u4_u2_U48 (.A2( u0_u4_u2_n105 ) , .A1( u0_u4_u2_n108 ) , .ZN( u0_u4_u2_n143 ) );
  NAND2_X1 u0_u4_u2_U49 (.A1( u0_u4_u2_n104 ) , .A2( u0_u4_u2_n106 ) , .ZN( u0_u4_u2_n152 ) );
  INV_X1 u0_u4_u2_U5 (.A( u0_u4_u2_n150 ) , .ZN( u0_u4_u2_n184 ) );
  NAND2_X1 u0_u4_u2_U50 (.A1( u0_u4_u2_n100 ) , .A2( u0_u4_u2_n105 ) , .ZN( u0_u4_u2_n132 ) );
  INV_X1 u0_u4_u2_U51 (.A( u0_u4_u2_n140 ) , .ZN( u0_u4_u2_n168 ) );
  INV_X1 u0_u4_u2_U52 (.A( u0_u4_u2_n138 ) , .ZN( u0_u4_u2_n167 ) );
  OAI21_X1 u0_u4_u2_U53 (.A( u0_u4_u2_n141 ) , .B2( u0_u4_u2_n142 ) , .ZN( u0_u4_u2_n146 ) , .B1( u0_u4_u2_n153 ) );
  OAI21_X1 u0_u4_u2_U54 (.A( u0_u4_u2_n140 ) , .ZN( u0_u4_u2_n141 ) , .B1( u0_u4_u2_n176 ) , .B2( u0_u4_u2_n177 ) );
  NOR3_X1 u0_u4_u2_U55 (.ZN( u0_u4_u2_n142 ) , .A3( u0_u4_u2_n175 ) , .A2( u0_u4_u2_n178 ) , .A1( u0_u4_u2_n181 ) );
  INV_X1 u0_u4_u2_U56 (.ZN( u0_u4_u2_n187 ) , .A( u0_u4_u2_n99 ) );
  OAI21_X1 u0_u4_u2_U57 (.B1( u0_u4_u2_n137 ) , .B2( u0_u4_u2_n143 ) , .A( u0_u4_u2_n98 ) , .ZN( u0_u4_u2_n99 ) );
  NAND2_X1 u0_u4_u2_U58 (.A1( u0_u4_u2_n102 ) , .A2( u0_u4_u2_n106 ) , .ZN( u0_u4_u2_n113 ) );
  NAND2_X1 u0_u4_u2_U59 (.A1( u0_u4_u2_n106 ) , .A2( u0_u4_u2_n107 ) , .ZN( u0_u4_u2_n131 ) );
  NOR4_X1 u0_u4_u2_U6 (.A4( u0_u4_u2_n124 ) , .A3( u0_u4_u2_n125 ) , .A2( u0_u4_u2_n126 ) , .A1( u0_u4_u2_n127 ) , .ZN( u0_u4_u2_n128 ) );
  NAND2_X1 u0_u4_u2_U60 (.A1( u0_u4_u2_n103 ) , .A2( u0_u4_u2_n107 ) , .ZN( u0_u4_u2_n139 ) );
  NAND2_X1 u0_u4_u2_U61 (.A1( u0_u4_u2_n103 ) , .A2( u0_u4_u2_n105 ) , .ZN( u0_u4_u2_n133 ) );
  NAND2_X1 u0_u4_u2_U62 (.A1( u0_u4_u2_n102 ) , .A2( u0_u4_u2_n103 ) , .ZN( u0_u4_u2_n154 ) );
  NAND2_X1 u0_u4_u2_U63 (.A2( u0_u4_u2_n103 ) , .A1( u0_u4_u2_n104 ) , .ZN( u0_u4_u2_n119 ) );
  NAND2_X1 u0_u4_u2_U64 (.A2( u0_u4_u2_n107 ) , .A1( u0_u4_u2_n108 ) , .ZN( u0_u4_u2_n123 ) );
  NAND2_X1 u0_u4_u2_U65 (.A1( u0_u4_u2_n104 ) , .A2( u0_u4_u2_n108 ) , .ZN( u0_u4_u2_n122 ) );
  INV_X1 u0_u4_u2_U66 (.A( u0_u4_u2_n114 ) , .ZN( u0_u4_u2_n172 ) );
  NAND2_X1 u0_u4_u2_U67 (.A2( u0_u4_u2_n100 ) , .A1( u0_u4_u2_n102 ) , .ZN( u0_u4_u2_n116 ) );
  NAND2_X1 u0_u4_u2_U68 (.A1( u0_u4_u2_n102 ) , .A2( u0_u4_u2_n108 ) , .ZN( u0_u4_u2_n120 ) );
  NAND2_X1 u0_u4_u2_U69 (.A2( u0_u4_u2_n105 ) , .A1( u0_u4_u2_n106 ) , .ZN( u0_u4_u2_n117 ) );
  AOI21_X1 u0_u4_u2_U7 (.B2( u0_u4_u2_n119 ) , .ZN( u0_u4_u2_n127 ) , .A( u0_u4_u2_n137 ) , .B1( u0_u4_u2_n155 ) );
  NOR2_X1 u0_u4_u2_U70 (.A2( u0_u4_X_16 ) , .ZN( u0_u4_u2_n140 ) , .A1( u0_u4_u2_n166 ) );
  NOR2_X1 u0_u4_u2_U71 (.A2( u0_u4_X_13 ) , .A1( u0_u4_X_14 ) , .ZN( u0_u4_u2_n100 ) );
  NOR2_X1 u0_u4_u2_U72 (.A2( u0_u4_X_16 ) , .A1( u0_u4_X_17 ) , .ZN( u0_u4_u2_n138 ) );
  NOR2_X1 u0_u4_u2_U73 (.A2( u0_u4_X_15 ) , .A1( u0_u4_X_18 ) , .ZN( u0_u4_u2_n104 ) );
  NOR2_X1 u0_u4_u2_U74 (.A2( u0_u4_X_14 ) , .ZN( u0_u4_u2_n103 ) , .A1( u0_u4_u2_n174 ) );
  NOR2_X1 u0_u4_u2_U75 (.A2( u0_u4_X_15 ) , .ZN( u0_u4_u2_n102 ) , .A1( u0_u4_u2_n165 ) );
  NOR2_X1 u0_u4_u2_U76 (.A2( u0_u4_X_17 ) , .ZN( u0_u4_u2_n114 ) , .A1( u0_u4_u2_n169 ) );
  AND2_X1 u0_u4_u2_U77 (.A1( u0_u4_X_15 ) , .ZN( u0_u4_u2_n105 ) , .A2( u0_u4_u2_n165 ) );
  AND2_X1 u0_u4_u2_U78 (.A2( u0_u4_X_15 ) , .A1( u0_u4_X_18 ) , .ZN( u0_u4_u2_n107 ) );
  AND2_X1 u0_u4_u2_U79 (.A1( u0_u4_X_14 ) , .ZN( u0_u4_u2_n106 ) , .A2( u0_u4_u2_n174 ) );
  AOI21_X1 u0_u4_u2_U8 (.ZN( u0_u4_u2_n124 ) , .B1( u0_u4_u2_n131 ) , .B2( u0_u4_u2_n143 ) , .A( u0_u4_u2_n172 ) );
  AND2_X1 u0_u4_u2_U80 (.A1( u0_u4_X_13 ) , .A2( u0_u4_X_14 ) , .ZN( u0_u4_u2_n108 ) );
  INV_X1 u0_u4_u2_U81 (.A( u0_u4_X_16 ) , .ZN( u0_u4_u2_n169 ) );
  INV_X1 u0_u4_u2_U82 (.A( u0_u4_X_17 ) , .ZN( u0_u4_u2_n166 ) );
  INV_X1 u0_u4_u2_U83 (.A( u0_u4_X_13 ) , .ZN( u0_u4_u2_n174 ) );
  INV_X1 u0_u4_u2_U84 (.A( u0_u4_X_18 ) , .ZN( u0_u4_u2_n165 ) );
  NAND4_X1 u0_u4_u2_U85 (.ZN( u0_out4_30 ) , .A4( u0_u4_u2_n147 ) , .A3( u0_u4_u2_n148 ) , .A2( u0_u4_u2_n149 ) , .A1( u0_u4_u2_n187 ) );
  NOR3_X1 u0_u4_u2_U86 (.A3( u0_u4_u2_n144 ) , .A2( u0_u4_u2_n145 ) , .A1( u0_u4_u2_n146 ) , .ZN( u0_u4_u2_n147 ) );
  AOI21_X1 u0_u4_u2_U87 (.B2( u0_u4_u2_n138 ) , .ZN( u0_u4_u2_n148 ) , .A( u0_u4_u2_n162 ) , .B1( u0_u4_u2_n182 ) );
  NAND4_X1 u0_u4_u2_U88 (.ZN( u0_out4_24 ) , .A4( u0_u4_u2_n111 ) , .A3( u0_u4_u2_n112 ) , .A1( u0_u4_u2_n130 ) , .A2( u0_u4_u2_n187 ) );
  AOI221_X1 u0_u4_u2_U89 (.A( u0_u4_u2_n109 ) , .B1( u0_u4_u2_n110 ) , .ZN( u0_u4_u2_n111 ) , .C1( u0_u4_u2_n134 ) , .C2( u0_u4_u2_n170 ) , .B2( u0_u4_u2_n173 ) );
  AOI21_X1 u0_u4_u2_U9 (.B2( u0_u4_u2_n123 ) , .ZN( u0_u4_u2_n125 ) , .A( u0_u4_u2_n171 ) , .B1( u0_u4_u2_n184 ) );
  AOI21_X1 u0_u4_u2_U90 (.ZN( u0_u4_u2_n112 ) , .B2( u0_u4_u2_n156 ) , .A( u0_u4_u2_n164 ) , .B1( u0_u4_u2_n181 ) );
  NAND4_X1 u0_u4_u2_U91 (.ZN( u0_out4_16 ) , .A4( u0_u4_u2_n128 ) , .A3( u0_u4_u2_n129 ) , .A1( u0_u4_u2_n130 ) , .A2( u0_u4_u2_n186 ) );
  AOI22_X1 u0_u4_u2_U92 (.A2( u0_u4_u2_n118 ) , .ZN( u0_u4_u2_n129 ) , .A1( u0_u4_u2_n140 ) , .B1( u0_u4_u2_n157 ) , .B2( u0_u4_u2_n170 ) );
  INV_X1 u0_u4_u2_U93 (.A( u0_u4_u2_n163 ) , .ZN( u0_u4_u2_n186 ) );
  OR4_X1 u0_u4_u2_U94 (.ZN( u0_out4_6 ) , .A4( u0_u4_u2_n161 ) , .A3( u0_u4_u2_n162 ) , .A2( u0_u4_u2_n163 ) , .A1( u0_u4_u2_n164 ) );
  OR3_X1 u0_u4_u2_U95 (.A2( u0_u4_u2_n159 ) , .A1( u0_u4_u2_n160 ) , .ZN( u0_u4_u2_n161 ) , .A3( u0_u4_u2_n183 ) );
  AOI21_X1 u0_u4_u2_U96 (.B2( u0_u4_u2_n154 ) , .B1( u0_u4_u2_n155 ) , .ZN( u0_u4_u2_n159 ) , .A( u0_u4_u2_n167 ) );
  NAND3_X1 u0_u4_u2_U97 (.A2( u0_u4_u2_n117 ) , .A1( u0_u4_u2_n122 ) , .A3( u0_u4_u2_n123 ) , .ZN( u0_u4_u2_n134 ) );
  NAND3_X1 u0_u4_u2_U98 (.ZN( u0_u4_u2_n110 ) , .A2( u0_u4_u2_n131 ) , .A3( u0_u4_u2_n139 ) , .A1( u0_u4_u2_n154 ) );
  NAND3_X1 u0_u4_u2_U99 (.A2( u0_u4_u2_n100 ) , .ZN( u0_u4_u2_n101 ) , .A1( u0_u4_u2_n104 ) , .A3( u0_u4_u2_n114 ) );
  OAI22_X1 u0_u4_u3_U10 (.B1( u0_u4_u3_n113 ) , .A2( u0_u4_u3_n135 ) , .A1( u0_u4_u3_n150 ) , .B2( u0_u4_u3_n164 ) , .ZN( u0_u4_u3_n98 ) );
  OAI211_X1 u0_u4_u3_U11 (.B( u0_u4_u3_n106 ) , .ZN( u0_u4_u3_n119 ) , .C2( u0_u4_u3_n128 ) , .C1( u0_u4_u3_n167 ) , .A( u0_u4_u3_n181 ) );
  AOI221_X1 u0_u4_u3_U12 (.C1( u0_u4_u3_n105 ) , .ZN( u0_u4_u3_n106 ) , .A( u0_u4_u3_n131 ) , .B2( u0_u4_u3_n132 ) , .C2( u0_u4_u3_n133 ) , .B1( u0_u4_u3_n169 ) );
  INV_X1 u0_u4_u3_U13 (.ZN( u0_u4_u3_n181 ) , .A( u0_u4_u3_n98 ) );
  NAND2_X1 u0_u4_u3_U14 (.ZN( u0_u4_u3_n105 ) , .A2( u0_u4_u3_n130 ) , .A1( u0_u4_u3_n155 ) );
  AOI22_X1 u0_u4_u3_U15 (.B1( u0_u4_u3_n115 ) , .A2( u0_u4_u3_n116 ) , .ZN( u0_u4_u3_n123 ) , .B2( u0_u4_u3_n133 ) , .A1( u0_u4_u3_n169 ) );
  NAND2_X1 u0_u4_u3_U16 (.ZN( u0_u4_u3_n116 ) , .A2( u0_u4_u3_n151 ) , .A1( u0_u4_u3_n182 ) );
  NOR2_X1 u0_u4_u3_U17 (.ZN( u0_u4_u3_n126 ) , .A2( u0_u4_u3_n150 ) , .A1( u0_u4_u3_n164 ) );
  AOI21_X1 u0_u4_u3_U18 (.ZN( u0_u4_u3_n112 ) , .B2( u0_u4_u3_n146 ) , .B1( u0_u4_u3_n155 ) , .A( u0_u4_u3_n167 ) );
  NAND2_X1 u0_u4_u3_U19 (.A1( u0_u4_u3_n135 ) , .ZN( u0_u4_u3_n142 ) , .A2( u0_u4_u3_n164 ) );
  NAND2_X1 u0_u4_u3_U20 (.ZN( u0_u4_u3_n132 ) , .A2( u0_u4_u3_n152 ) , .A1( u0_u4_u3_n156 ) );
  AND2_X1 u0_u4_u3_U21 (.A2( u0_u4_u3_n113 ) , .A1( u0_u4_u3_n114 ) , .ZN( u0_u4_u3_n151 ) );
  INV_X1 u0_u4_u3_U22 (.A( u0_u4_u3_n133 ) , .ZN( u0_u4_u3_n165 ) );
  INV_X1 u0_u4_u3_U23 (.A( u0_u4_u3_n135 ) , .ZN( u0_u4_u3_n170 ) );
  NAND2_X1 u0_u4_u3_U24 (.A1( u0_u4_u3_n107 ) , .A2( u0_u4_u3_n108 ) , .ZN( u0_u4_u3_n140 ) );
  NAND2_X1 u0_u4_u3_U25 (.ZN( u0_u4_u3_n117 ) , .A1( u0_u4_u3_n124 ) , .A2( u0_u4_u3_n148 ) );
  NAND2_X1 u0_u4_u3_U26 (.ZN( u0_u4_u3_n143 ) , .A1( u0_u4_u3_n165 ) , .A2( u0_u4_u3_n167 ) );
  INV_X1 u0_u4_u3_U27 (.A( u0_u4_u3_n130 ) , .ZN( u0_u4_u3_n177 ) );
  INV_X1 u0_u4_u3_U28 (.A( u0_u4_u3_n128 ) , .ZN( u0_u4_u3_n176 ) );
  INV_X1 u0_u4_u3_U29 (.A( u0_u4_u3_n155 ) , .ZN( u0_u4_u3_n174 ) );
  INV_X1 u0_u4_u3_U3 (.A( u0_u4_u3_n129 ) , .ZN( u0_u4_u3_n183 ) );
  INV_X1 u0_u4_u3_U30 (.A( u0_u4_u3_n139 ) , .ZN( u0_u4_u3_n185 ) );
  NOR2_X1 u0_u4_u3_U31 (.ZN( u0_u4_u3_n135 ) , .A2( u0_u4_u3_n141 ) , .A1( u0_u4_u3_n169 ) );
  OAI222_X1 u0_u4_u3_U32 (.C2( u0_u4_u3_n107 ) , .A2( u0_u4_u3_n108 ) , .B1( u0_u4_u3_n135 ) , .ZN( u0_u4_u3_n138 ) , .B2( u0_u4_u3_n146 ) , .C1( u0_u4_u3_n154 ) , .A1( u0_u4_u3_n164 ) );
  NOR4_X1 u0_u4_u3_U33 (.A4( u0_u4_u3_n157 ) , .A3( u0_u4_u3_n158 ) , .A2( u0_u4_u3_n159 ) , .A1( u0_u4_u3_n160 ) , .ZN( u0_u4_u3_n161 ) );
  AOI21_X1 u0_u4_u3_U34 (.B2( u0_u4_u3_n152 ) , .B1( u0_u4_u3_n153 ) , .ZN( u0_u4_u3_n158 ) , .A( u0_u4_u3_n164 ) );
  AOI21_X1 u0_u4_u3_U35 (.A( u0_u4_u3_n149 ) , .B2( u0_u4_u3_n150 ) , .B1( u0_u4_u3_n151 ) , .ZN( u0_u4_u3_n159 ) );
  AOI21_X1 u0_u4_u3_U36 (.A( u0_u4_u3_n154 ) , .B2( u0_u4_u3_n155 ) , .B1( u0_u4_u3_n156 ) , .ZN( u0_u4_u3_n157 ) );
  AOI211_X1 u0_u4_u3_U37 (.ZN( u0_u4_u3_n109 ) , .A( u0_u4_u3_n119 ) , .C2( u0_u4_u3_n129 ) , .B( u0_u4_u3_n138 ) , .C1( u0_u4_u3_n141 ) );
  AOI211_X1 u0_u4_u3_U38 (.B( u0_u4_u3_n119 ) , .A( u0_u4_u3_n120 ) , .C2( u0_u4_u3_n121 ) , .ZN( u0_u4_u3_n122 ) , .C1( u0_u4_u3_n179 ) );
  INV_X1 u0_u4_u3_U39 (.A( u0_u4_u3_n156 ) , .ZN( u0_u4_u3_n179 ) );
  INV_X1 u0_u4_u3_U4 (.A( u0_u4_u3_n140 ) , .ZN( u0_u4_u3_n182 ) );
  OAI22_X1 u0_u4_u3_U40 (.B1( u0_u4_u3_n118 ) , .ZN( u0_u4_u3_n120 ) , .A1( u0_u4_u3_n135 ) , .B2( u0_u4_u3_n154 ) , .A2( u0_u4_u3_n178 ) );
  AND3_X1 u0_u4_u3_U41 (.ZN( u0_u4_u3_n118 ) , .A2( u0_u4_u3_n124 ) , .A1( u0_u4_u3_n144 ) , .A3( u0_u4_u3_n152 ) );
  INV_X1 u0_u4_u3_U42 (.A( u0_u4_u3_n121 ) , .ZN( u0_u4_u3_n164 ) );
  NAND2_X1 u0_u4_u3_U43 (.ZN( u0_u4_u3_n133 ) , .A1( u0_u4_u3_n154 ) , .A2( u0_u4_u3_n164 ) );
  OAI211_X1 u0_u4_u3_U44 (.B( u0_u4_u3_n127 ) , .ZN( u0_u4_u3_n139 ) , .C1( u0_u4_u3_n150 ) , .C2( u0_u4_u3_n154 ) , .A( u0_u4_u3_n184 ) );
  INV_X1 u0_u4_u3_U45 (.A( u0_u4_u3_n125 ) , .ZN( u0_u4_u3_n184 ) );
  AOI221_X1 u0_u4_u3_U46 (.A( u0_u4_u3_n126 ) , .ZN( u0_u4_u3_n127 ) , .C2( u0_u4_u3_n132 ) , .C1( u0_u4_u3_n169 ) , .B2( u0_u4_u3_n170 ) , .B1( u0_u4_u3_n174 ) );
  OAI22_X1 u0_u4_u3_U47 (.A1( u0_u4_u3_n124 ) , .ZN( u0_u4_u3_n125 ) , .B2( u0_u4_u3_n145 ) , .A2( u0_u4_u3_n165 ) , .B1( u0_u4_u3_n167 ) );
  NOR2_X1 u0_u4_u3_U48 (.A1( u0_u4_u3_n113 ) , .ZN( u0_u4_u3_n131 ) , .A2( u0_u4_u3_n154 ) );
  NAND2_X1 u0_u4_u3_U49 (.A1( u0_u4_u3_n103 ) , .ZN( u0_u4_u3_n150 ) , .A2( u0_u4_u3_n99 ) );
  INV_X1 u0_u4_u3_U5 (.A( u0_u4_u3_n117 ) , .ZN( u0_u4_u3_n178 ) );
  NAND2_X1 u0_u4_u3_U50 (.A2( u0_u4_u3_n102 ) , .ZN( u0_u4_u3_n155 ) , .A1( u0_u4_u3_n97 ) );
  INV_X1 u0_u4_u3_U51 (.A( u0_u4_u3_n141 ) , .ZN( u0_u4_u3_n167 ) );
  AOI21_X1 u0_u4_u3_U52 (.B2( u0_u4_u3_n114 ) , .B1( u0_u4_u3_n146 ) , .A( u0_u4_u3_n154 ) , .ZN( u0_u4_u3_n94 ) );
  AOI21_X1 u0_u4_u3_U53 (.ZN( u0_u4_u3_n110 ) , .B2( u0_u4_u3_n142 ) , .B1( u0_u4_u3_n186 ) , .A( u0_u4_u3_n95 ) );
  INV_X1 u0_u4_u3_U54 (.A( u0_u4_u3_n145 ) , .ZN( u0_u4_u3_n186 ) );
  AOI21_X1 u0_u4_u3_U55 (.B1( u0_u4_u3_n124 ) , .A( u0_u4_u3_n149 ) , .B2( u0_u4_u3_n155 ) , .ZN( u0_u4_u3_n95 ) );
  INV_X1 u0_u4_u3_U56 (.A( u0_u4_u3_n149 ) , .ZN( u0_u4_u3_n169 ) );
  NAND2_X1 u0_u4_u3_U57 (.ZN( u0_u4_u3_n124 ) , .A1( u0_u4_u3_n96 ) , .A2( u0_u4_u3_n97 ) );
  NAND2_X1 u0_u4_u3_U58 (.A2( u0_u4_u3_n100 ) , .ZN( u0_u4_u3_n146 ) , .A1( u0_u4_u3_n96 ) );
  NAND2_X1 u0_u4_u3_U59 (.A1( u0_u4_u3_n101 ) , .ZN( u0_u4_u3_n145 ) , .A2( u0_u4_u3_n99 ) );
  AOI221_X1 u0_u4_u3_U6 (.A( u0_u4_u3_n131 ) , .C2( u0_u4_u3_n132 ) , .C1( u0_u4_u3_n133 ) , .ZN( u0_u4_u3_n134 ) , .B1( u0_u4_u3_n143 ) , .B2( u0_u4_u3_n177 ) );
  NAND2_X1 u0_u4_u3_U60 (.A1( u0_u4_u3_n100 ) , .ZN( u0_u4_u3_n156 ) , .A2( u0_u4_u3_n99 ) );
  NAND2_X1 u0_u4_u3_U61 (.A2( u0_u4_u3_n101 ) , .A1( u0_u4_u3_n104 ) , .ZN( u0_u4_u3_n148 ) );
  NAND2_X1 u0_u4_u3_U62 (.A1( u0_u4_u3_n100 ) , .A2( u0_u4_u3_n102 ) , .ZN( u0_u4_u3_n128 ) );
  NAND2_X1 u0_u4_u3_U63 (.A2( u0_u4_u3_n101 ) , .A1( u0_u4_u3_n102 ) , .ZN( u0_u4_u3_n152 ) );
  NAND2_X1 u0_u4_u3_U64 (.A2( u0_u4_u3_n101 ) , .ZN( u0_u4_u3_n114 ) , .A1( u0_u4_u3_n96 ) );
  NAND2_X1 u0_u4_u3_U65 (.ZN( u0_u4_u3_n107 ) , .A1( u0_u4_u3_n97 ) , .A2( u0_u4_u3_n99 ) );
  NAND2_X1 u0_u4_u3_U66 (.A2( u0_u4_u3_n100 ) , .A1( u0_u4_u3_n104 ) , .ZN( u0_u4_u3_n113 ) );
  NAND2_X1 u0_u4_u3_U67 (.A1( u0_u4_u3_n104 ) , .ZN( u0_u4_u3_n153 ) , .A2( u0_u4_u3_n97 ) );
  NAND2_X1 u0_u4_u3_U68 (.A2( u0_u4_u3_n103 ) , .A1( u0_u4_u3_n104 ) , .ZN( u0_u4_u3_n130 ) );
  NAND2_X1 u0_u4_u3_U69 (.A2( u0_u4_u3_n103 ) , .ZN( u0_u4_u3_n144 ) , .A1( u0_u4_u3_n96 ) );
  OAI22_X1 u0_u4_u3_U7 (.B2( u0_u4_u3_n147 ) , .A2( u0_u4_u3_n148 ) , .ZN( u0_u4_u3_n160 ) , .B1( u0_u4_u3_n165 ) , .A1( u0_u4_u3_n168 ) );
  NAND2_X1 u0_u4_u3_U70 (.A1( u0_u4_u3_n102 ) , .A2( u0_u4_u3_n103 ) , .ZN( u0_u4_u3_n108 ) );
  NOR2_X1 u0_u4_u3_U71 (.A2( u0_u4_X_19 ) , .A1( u0_u4_X_20 ) , .ZN( u0_u4_u3_n99 ) );
  NOR2_X1 u0_u4_u3_U72 (.A2( u0_u4_X_21 ) , .A1( u0_u4_X_24 ) , .ZN( u0_u4_u3_n103 ) );
  NOR2_X1 u0_u4_u3_U73 (.A2( u0_u4_X_24 ) , .A1( u0_u4_u3_n171 ) , .ZN( u0_u4_u3_n97 ) );
  NOR2_X1 u0_u4_u3_U74 (.A2( u0_u4_X_23 ) , .ZN( u0_u4_u3_n141 ) , .A1( u0_u4_u3_n166 ) );
  NOR2_X1 u0_u4_u3_U75 (.A2( u0_u4_X_19 ) , .A1( u0_u4_u3_n172 ) , .ZN( u0_u4_u3_n96 ) );
  NAND2_X1 u0_u4_u3_U76 (.A1( u0_u4_X_22 ) , .A2( u0_u4_X_23 ) , .ZN( u0_u4_u3_n154 ) );
  NAND2_X1 u0_u4_u3_U77 (.A1( u0_u4_X_23 ) , .ZN( u0_u4_u3_n149 ) , .A2( u0_u4_u3_n166 ) );
  NOR2_X1 u0_u4_u3_U78 (.A2( u0_u4_X_22 ) , .A1( u0_u4_X_23 ) , .ZN( u0_u4_u3_n121 ) );
  AND2_X1 u0_u4_u3_U79 (.A1( u0_u4_X_24 ) , .ZN( u0_u4_u3_n101 ) , .A2( u0_u4_u3_n171 ) );
  AND3_X1 u0_u4_u3_U8 (.A3( u0_u4_u3_n144 ) , .A2( u0_u4_u3_n145 ) , .A1( u0_u4_u3_n146 ) , .ZN( u0_u4_u3_n147 ) );
  AND2_X1 u0_u4_u3_U80 (.A1( u0_u4_X_19 ) , .ZN( u0_u4_u3_n102 ) , .A2( u0_u4_u3_n172 ) );
  AND2_X1 u0_u4_u3_U81 (.A1( u0_u4_X_21 ) , .A2( u0_u4_X_24 ) , .ZN( u0_u4_u3_n100 ) );
  AND2_X1 u0_u4_u3_U82 (.A2( u0_u4_X_19 ) , .A1( u0_u4_X_20 ) , .ZN( u0_u4_u3_n104 ) );
  INV_X1 u0_u4_u3_U83 (.A( u0_u4_X_22 ) , .ZN( u0_u4_u3_n166 ) );
  INV_X1 u0_u4_u3_U84 (.A( u0_u4_X_21 ) , .ZN( u0_u4_u3_n171 ) );
  INV_X1 u0_u4_u3_U85 (.A( u0_u4_X_20 ) , .ZN( u0_u4_u3_n172 ) );
  OR4_X1 u0_u4_u3_U86 (.ZN( u0_out4_10 ) , .A4( u0_u4_u3_n136 ) , .A3( u0_u4_u3_n137 ) , .A1( u0_u4_u3_n138 ) , .A2( u0_u4_u3_n139 ) );
  OAI222_X1 u0_u4_u3_U87 (.C1( u0_u4_u3_n128 ) , .ZN( u0_u4_u3_n137 ) , .B1( u0_u4_u3_n148 ) , .A2( u0_u4_u3_n150 ) , .B2( u0_u4_u3_n154 ) , .C2( u0_u4_u3_n164 ) , .A1( u0_u4_u3_n167 ) );
  OAI221_X1 u0_u4_u3_U88 (.A( u0_u4_u3_n134 ) , .B2( u0_u4_u3_n135 ) , .ZN( u0_u4_u3_n136 ) , .C1( u0_u4_u3_n149 ) , .B1( u0_u4_u3_n151 ) , .C2( u0_u4_u3_n183 ) );
  NAND4_X1 u0_u4_u3_U89 (.ZN( u0_out4_26 ) , .A4( u0_u4_u3_n109 ) , .A3( u0_u4_u3_n110 ) , .A2( u0_u4_u3_n111 ) , .A1( u0_u4_u3_n173 ) );
  INV_X1 u0_u4_u3_U9 (.A( u0_u4_u3_n143 ) , .ZN( u0_u4_u3_n168 ) );
  INV_X1 u0_u4_u3_U90 (.ZN( u0_u4_u3_n173 ) , .A( u0_u4_u3_n94 ) );
  OAI21_X1 u0_u4_u3_U91 (.ZN( u0_u4_u3_n111 ) , .B2( u0_u4_u3_n117 ) , .A( u0_u4_u3_n133 ) , .B1( u0_u4_u3_n176 ) );
  NAND4_X1 u0_u4_u3_U92 (.ZN( u0_out4_20 ) , .A4( u0_u4_u3_n122 ) , .A3( u0_u4_u3_n123 ) , .A1( u0_u4_u3_n175 ) , .A2( u0_u4_u3_n180 ) );
  INV_X1 u0_u4_u3_U93 (.A( u0_u4_u3_n126 ) , .ZN( u0_u4_u3_n180 ) );
  INV_X1 u0_u4_u3_U94 (.A( u0_u4_u3_n112 ) , .ZN( u0_u4_u3_n175 ) );
  NAND4_X1 u0_u4_u3_U95 (.ZN( u0_out4_1 ) , .A4( u0_u4_u3_n161 ) , .A3( u0_u4_u3_n162 ) , .A2( u0_u4_u3_n163 ) , .A1( u0_u4_u3_n185 ) );
  NAND2_X1 u0_u4_u3_U96 (.ZN( u0_u4_u3_n163 ) , .A2( u0_u4_u3_n170 ) , .A1( u0_u4_u3_n176 ) );
  AOI22_X1 u0_u4_u3_U97 (.B2( u0_u4_u3_n140 ) , .B1( u0_u4_u3_n141 ) , .A2( u0_u4_u3_n142 ) , .ZN( u0_u4_u3_n162 ) , .A1( u0_u4_u3_n177 ) );
  NAND3_X1 u0_u4_u3_U98 (.A1( u0_u4_u3_n114 ) , .ZN( u0_u4_u3_n115 ) , .A2( u0_u4_u3_n145 ) , .A3( u0_u4_u3_n153 ) );
  NAND3_X1 u0_u4_u3_U99 (.ZN( u0_u4_u3_n129 ) , .A2( u0_u4_u3_n144 ) , .A1( u0_u4_u3_n153 ) , .A3( u0_u4_u3_n182 ) );
  XOR2_X1 u0_u6_U13 (.B( u0_K7_42 ) , .A( u0_R5_29 ) , .Z( u0_u6_X_42 ) );
  XOR2_X1 u0_u6_U14 (.B( u0_K7_41 ) , .A( u0_R5_28 ) , .Z( u0_u6_X_41 ) );
  XOR2_X1 u0_u6_U15 (.B( u0_K7_40 ) , .A( u0_R5_27 ) , .Z( u0_u6_X_40 ) );
  XOR2_X1 u0_u6_U17 (.B( u0_K7_39 ) , .A( u0_R5_26 ) , .Z( u0_u6_X_39 ) );
  XOR2_X1 u0_u6_U18 (.B( u0_K7_38 ) , .A( u0_R5_25 ) , .Z( u0_u6_X_38 ) );
  XOR2_X1 u0_u6_U19 (.B( u0_K7_37 ) , .A( u0_R5_24 ) , .Z( u0_u6_X_37 ) );
  XOR2_X1 u0_u6_U20 (.B( u0_K7_36 ) , .A( u0_R5_25 ) , .Z( u0_u6_X_36 ) );
  XOR2_X1 u0_u6_U21 (.B( u0_K7_35 ) , .A( u0_R5_24 ) , .Z( u0_u6_X_35 ) );
  XOR2_X1 u0_u6_U22 (.B( u0_K7_34 ) , .A( u0_R5_23 ) , .Z( u0_u6_X_34 ) );
  XOR2_X1 u0_u6_U23 (.B( u0_K7_33 ) , .A( u0_R5_22 ) , .Z( u0_u6_X_33 ) );
  XOR2_X1 u0_u6_U24 (.B( u0_K7_32 ) , .A( u0_R5_21 ) , .Z( u0_u6_X_32 ) );
  XOR2_X1 u0_u6_U25 (.B( u0_K7_31 ) , .A( u0_R5_20 ) , .Z( u0_u6_X_31 ) );
  XOR2_X1 u0_u6_U26 (.B( u0_K7_30 ) , .A( u0_R5_21 ) , .Z( u0_u6_X_30 ) );
  XOR2_X1 u0_u6_U28 (.B( u0_K7_29 ) , .A( u0_R5_20 ) , .Z( u0_u6_X_29 ) );
  XOR2_X1 u0_u6_U29 (.B( u0_K7_28 ) , .A( u0_R5_19 ) , .Z( u0_u6_X_28 ) );
  XOR2_X1 u0_u6_U30 (.B( u0_K7_27 ) , .A( u0_R5_18 ) , .Z( u0_u6_X_27 ) );
  XOR2_X1 u0_u6_U31 (.B( u0_K7_26 ) , .A( u0_R5_17 ) , .Z( u0_u6_X_26 ) );
  XOR2_X1 u0_u6_U32 (.B( u0_K7_25 ) , .A( u0_R5_16 ) , .Z( u0_u6_X_25 ) );
  OAI22_X1 u0_u6_u4_U10 (.B2( u0_u6_u4_n135 ) , .ZN( u0_u6_u4_n137 ) , .B1( u0_u6_u4_n153 ) , .A1( u0_u6_u4_n155 ) , .A2( u0_u6_u4_n171 ) );
  AND3_X1 u0_u6_u4_U11 (.A2( u0_u6_u4_n134 ) , .ZN( u0_u6_u4_n135 ) , .A3( u0_u6_u4_n145 ) , .A1( u0_u6_u4_n157 ) );
  NAND2_X1 u0_u6_u4_U12 (.ZN( u0_u6_u4_n132 ) , .A2( u0_u6_u4_n170 ) , .A1( u0_u6_u4_n173 ) );
  AOI21_X1 u0_u6_u4_U13 (.B2( u0_u6_u4_n160 ) , .B1( u0_u6_u4_n161 ) , .ZN( u0_u6_u4_n162 ) , .A( u0_u6_u4_n170 ) );
  AOI21_X1 u0_u6_u4_U14 (.ZN( u0_u6_u4_n107 ) , .B2( u0_u6_u4_n143 ) , .A( u0_u6_u4_n174 ) , .B1( u0_u6_u4_n184 ) );
  AOI21_X1 u0_u6_u4_U15 (.B2( u0_u6_u4_n158 ) , .B1( u0_u6_u4_n159 ) , .ZN( u0_u6_u4_n163 ) , .A( u0_u6_u4_n174 ) );
  AOI21_X1 u0_u6_u4_U16 (.A( u0_u6_u4_n153 ) , .B2( u0_u6_u4_n154 ) , .B1( u0_u6_u4_n155 ) , .ZN( u0_u6_u4_n165 ) );
  AOI21_X1 u0_u6_u4_U17 (.A( u0_u6_u4_n156 ) , .B2( u0_u6_u4_n157 ) , .ZN( u0_u6_u4_n164 ) , .B1( u0_u6_u4_n184 ) );
  INV_X1 u0_u6_u4_U18 (.A( u0_u6_u4_n138 ) , .ZN( u0_u6_u4_n170 ) );
  AND2_X1 u0_u6_u4_U19 (.A2( u0_u6_u4_n120 ) , .ZN( u0_u6_u4_n155 ) , .A1( u0_u6_u4_n160 ) );
  INV_X1 u0_u6_u4_U20 (.A( u0_u6_u4_n156 ) , .ZN( u0_u6_u4_n175 ) );
  NAND2_X1 u0_u6_u4_U21 (.A2( u0_u6_u4_n118 ) , .ZN( u0_u6_u4_n131 ) , .A1( u0_u6_u4_n147 ) );
  NAND2_X1 u0_u6_u4_U22 (.A1( u0_u6_u4_n119 ) , .A2( u0_u6_u4_n120 ) , .ZN( u0_u6_u4_n130 ) );
  NAND2_X1 u0_u6_u4_U23 (.ZN( u0_u6_u4_n117 ) , .A2( u0_u6_u4_n118 ) , .A1( u0_u6_u4_n148 ) );
  NAND2_X1 u0_u6_u4_U24 (.ZN( u0_u6_u4_n129 ) , .A1( u0_u6_u4_n134 ) , .A2( u0_u6_u4_n148 ) );
  AND3_X1 u0_u6_u4_U25 (.A1( u0_u6_u4_n119 ) , .A2( u0_u6_u4_n143 ) , .A3( u0_u6_u4_n154 ) , .ZN( u0_u6_u4_n161 ) );
  AND2_X1 u0_u6_u4_U26 (.A1( u0_u6_u4_n145 ) , .A2( u0_u6_u4_n147 ) , .ZN( u0_u6_u4_n159 ) );
  OR3_X1 u0_u6_u4_U27 (.A3( u0_u6_u4_n114 ) , .A2( u0_u6_u4_n115 ) , .A1( u0_u6_u4_n116 ) , .ZN( u0_u6_u4_n136 ) );
  AOI21_X1 u0_u6_u4_U28 (.A( u0_u6_u4_n113 ) , .ZN( u0_u6_u4_n116 ) , .B2( u0_u6_u4_n173 ) , .B1( u0_u6_u4_n174 ) );
  AOI21_X1 u0_u6_u4_U29 (.ZN( u0_u6_u4_n115 ) , .B2( u0_u6_u4_n145 ) , .B1( u0_u6_u4_n146 ) , .A( u0_u6_u4_n156 ) );
  NOR2_X1 u0_u6_u4_U3 (.ZN( u0_u6_u4_n121 ) , .A1( u0_u6_u4_n181 ) , .A2( u0_u6_u4_n182 ) );
  OAI22_X1 u0_u6_u4_U30 (.ZN( u0_u6_u4_n114 ) , .A2( u0_u6_u4_n121 ) , .B1( u0_u6_u4_n160 ) , .B2( u0_u6_u4_n170 ) , .A1( u0_u6_u4_n171 ) );
  INV_X1 u0_u6_u4_U31 (.A( u0_u6_u4_n158 ) , .ZN( u0_u6_u4_n182 ) );
  INV_X1 u0_u6_u4_U32 (.ZN( u0_u6_u4_n181 ) , .A( u0_u6_u4_n96 ) );
  INV_X1 u0_u6_u4_U33 (.A( u0_u6_u4_n144 ) , .ZN( u0_u6_u4_n179 ) );
  INV_X1 u0_u6_u4_U34 (.A( u0_u6_u4_n157 ) , .ZN( u0_u6_u4_n178 ) );
  NAND2_X1 u0_u6_u4_U35 (.A2( u0_u6_u4_n154 ) , .A1( u0_u6_u4_n96 ) , .ZN( u0_u6_u4_n97 ) );
  INV_X1 u0_u6_u4_U36 (.ZN( u0_u6_u4_n186 ) , .A( u0_u6_u4_n95 ) );
  OAI221_X1 u0_u6_u4_U37 (.C1( u0_u6_u4_n134 ) , .B1( u0_u6_u4_n158 ) , .B2( u0_u6_u4_n171 ) , .C2( u0_u6_u4_n173 ) , .A( u0_u6_u4_n94 ) , .ZN( u0_u6_u4_n95 ) );
  AOI222_X1 u0_u6_u4_U38 (.B2( u0_u6_u4_n132 ) , .A1( u0_u6_u4_n138 ) , .C2( u0_u6_u4_n175 ) , .A2( u0_u6_u4_n179 ) , .C1( u0_u6_u4_n181 ) , .B1( u0_u6_u4_n185 ) , .ZN( u0_u6_u4_n94 ) );
  INV_X1 u0_u6_u4_U39 (.A( u0_u6_u4_n113 ) , .ZN( u0_u6_u4_n185 ) );
  INV_X1 u0_u6_u4_U4 (.A( u0_u6_u4_n117 ) , .ZN( u0_u6_u4_n184 ) );
  INV_X1 u0_u6_u4_U40 (.A( u0_u6_u4_n143 ) , .ZN( u0_u6_u4_n183 ) );
  NOR2_X1 u0_u6_u4_U41 (.ZN( u0_u6_u4_n138 ) , .A1( u0_u6_u4_n168 ) , .A2( u0_u6_u4_n169 ) );
  NOR2_X1 u0_u6_u4_U42 (.A1( u0_u6_u4_n150 ) , .A2( u0_u6_u4_n152 ) , .ZN( u0_u6_u4_n153 ) );
  NOR2_X1 u0_u6_u4_U43 (.A2( u0_u6_u4_n128 ) , .A1( u0_u6_u4_n138 ) , .ZN( u0_u6_u4_n156 ) );
  AOI22_X1 u0_u6_u4_U44 (.B2( u0_u6_u4_n122 ) , .A1( u0_u6_u4_n123 ) , .ZN( u0_u6_u4_n124 ) , .B1( u0_u6_u4_n128 ) , .A2( u0_u6_u4_n172 ) );
  INV_X1 u0_u6_u4_U45 (.A( u0_u6_u4_n153 ) , .ZN( u0_u6_u4_n172 ) );
  NAND2_X1 u0_u6_u4_U46 (.A2( u0_u6_u4_n120 ) , .ZN( u0_u6_u4_n123 ) , .A1( u0_u6_u4_n161 ) );
  AOI22_X1 u0_u6_u4_U47 (.B2( u0_u6_u4_n132 ) , .A2( u0_u6_u4_n133 ) , .ZN( u0_u6_u4_n140 ) , .A1( u0_u6_u4_n150 ) , .B1( u0_u6_u4_n179 ) );
  NAND2_X1 u0_u6_u4_U48 (.ZN( u0_u6_u4_n133 ) , .A2( u0_u6_u4_n146 ) , .A1( u0_u6_u4_n154 ) );
  NAND2_X1 u0_u6_u4_U49 (.A1( u0_u6_u4_n103 ) , .ZN( u0_u6_u4_n154 ) , .A2( u0_u6_u4_n98 ) );
  NOR4_X1 u0_u6_u4_U5 (.A4( u0_u6_u4_n106 ) , .A3( u0_u6_u4_n107 ) , .A2( u0_u6_u4_n108 ) , .A1( u0_u6_u4_n109 ) , .ZN( u0_u6_u4_n110 ) );
  NAND2_X1 u0_u6_u4_U50 (.A1( u0_u6_u4_n101 ) , .ZN( u0_u6_u4_n158 ) , .A2( u0_u6_u4_n99 ) );
  AOI21_X1 u0_u6_u4_U51 (.ZN( u0_u6_u4_n127 ) , .A( u0_u6_u4_n136 ) , .B2( u0_u6_u4_n150 ) , .B1( u0_u6_u4_n180 ) );
  INV_X1 u0_u6_u4_U52 (.A( u0_u6_u4_n160 ) , .ZN( u0_u6_u4_n180 ) );
  NAND2_X1 u0_u6_u4_U53 (.A2( u0_u6_u4_n104 ) , .A1( u0_u6_u4_n105 ) , .ZN( u0_u6_u4_n146 ) );
  NAND2_X1 u0_u6_u4_U54 (.A2( u0_u6_u4_n101 ) , .A1( u0_u6_u4_n102 ) , .ZN( u0_u6_u4_n160 ) );
  NAND2_X1 u0_u6_u4_U55 (.ZN( u0_u6_u4_n134 ) , .A1( u0_u6_u4_n98 ) , .A2( u0_u6_u4_n99 ) );
  NAND2_X1 u0_u6_u4_U56 (.A1( u0_u6_u4_n103 ) , .A2( u0_u6_u4_n104 ) , .ZN( u0_u6_u4_n143 ) );
  NAND2_X1 u0_u6_u4_U57 (.A2( u0_u6_u4_n105 ) , .ZN( u0_u6_u4_n145 ) , .A1( u0_u6_u4_n98 ) );
  NAND2_X1 u0_u6_u4_U58 (.A1( u0_u6_u4_n100 ) , .A2( u0_u6_u4_n105 ) , .ZN( u0_u6_u4_n120 ) );
  NAND2_X1 u0_u6_u4_U59 (.A1( u0_u6_u4_n102 ) , .A2( u0_u6_u4_n104 ) , .ZN( u0_u6_u4_n148 ) );
  AOI21_X1 u0_u6_u4_U6 (.ZN( u0_u6_u4_n106 ) , .B2( u0_u6_u4_n146 ) , .B1( u0_u6_u4_n158 ) , .A( u0_u6_u4_n170 ) );
  NAND2_X1 u0_u6_u4_U60 (.A2( u0_u6_u4_n100 ) , .A1( u0_u6_u4_n103 ) , .ZN( u0_u6_u4_n157 ) );
  INV_X1 u0_u6_u4_U61 (.A( u0_u6_u4_n150 ) , .ZN( u0_u6_u4_n173 ) );
  INV_X1 u0_u6_u4_U62 (.A( u0_u6_u4_n152 ) , .ZN( u0_u6_u4_n171 ) );
  NAND2_X1 u0_u6_u4_U63 (.A1( u0_u6_u4_n100 ) , .ZN( u0_u6_u4_n118 ) , .A2( u0_u6_u4_n99 ) );
  NAND2_X1 u0_u6_u4_U64 (.A2( u0_u6_u4_n100 ) , .A1( u0_u6_u4_n102 ) , .ZN( u0_u6_u4_n144 ) );
  NAND2_X1 u0_u6_u4_U65 (.A2( u0_u6_u4_n101 ) , .A1( u0_u6_u4_n105 ) , .ZN( u0_u6_u4_n96 ) );
  INV_X1 u0_u6_u4_U66 (.A( u0_u6_u4_n128 ) , .ZN( u0_u6_u4_n174 ) );
  NAND2_X1 u0_u6_u4_U67 (.A2( u0_u6_u4_n102 ) , .ZN( u0_u6_u4_n119 ) , .A1( u0_u6_u4_n98 ) );
  NAND2_X1 u0_u6_u4_U68 (.A2( u0_u6_u4_n101 ) , .A1( u0_u6_u4_n103 ) , .ZN( u0_u6_u4_n147 ) );
  NAND2_X1 u0_u6_u4_U69 (.A2( u0_u6_u4_n104 ) , .ZN( u0_u6_u4_n113 ) , .A1( u0_u6_u4_n99 ) );
  AOI21_X1 u0_u6_u4_U7 (.ZN( u0_u6_u4_n108 ) , .B2( u0_u6_u4_n134 ) , .B1( u0_u6_u4_n155 ) , .A( u0_u6_u4_n156 ) );
  NOR2_X1 u0_u6_u4_U70 (.A2( u0_u6_X_28 ) , .ZN( u0_u6_u4_n150 ) , .A1( u0_u6_u4_n168 ) );
  NOR2_X1 u0_u6_u4_U71 (.A2( u0_u6_X_29 ) , .ZN( u0_u6_u4_n152 ) , .A1( u0_u6_u4_n169 ) );
  NOR2_X1 u0_u6_u4_U72 (.A2( u0_u6_X_30 ) , .ZN( u0_u6_u4_n105 ) , .A1( u0_u6_u4_n176 ) );
  NOR2_X1 u0_u6_u4_U73 (.A2( u0_u6_X_26 ) , .ZN( u0_u6_u4_n100 ) , .A1( u0_u6_u4_n177 ) );
  NOR2_X1 u0_u6_u4_U74 (.A2( u0_u6_X_28 ) , .A1( u0_u6_X_29 ) , .ZN( u0_u6_u4_n128 ) );
  NOR2_X1 u0_u6_u4_U75 (.A2( u0_u6_X_27 ) , .A1( u0_u6_X_30 ) , .ZN( u0_u6_u4_n102 ) );
  NOR2_X1 u0_u6_u4_U76 (.A2( u0_u6_X_25 ) , .A1( u0_u6_X_26 ) , .ZN( u0_u6_u4_n98 ) );
  AND2_X1 u0_u6_u4_U77 (.A2( u0_u6_X_25 ) , .A1( u0_u6_X_26 ) , .ZN( u0_u6_u4_n104 ) );
  AND2_X1 u0_u6_u4_U78 (.A1( u0_u6_X_30 ) , .A2( u0_u6_u4_n176 ) , .ZN( u0_u6_u4_n99 ) );
  AND2_X1 u0_u6_u4_U79 (.A1( u0_u6_X_26 ) , .ZN( u0_u6_u4_n101 ) , .A2( u0_u6_u4_n177 ) );
  AOI21_X1 u0_u6_u4_U8 (.ZN( u0_u6_u4_n109 ) , .A( u0_u6_u4_n153 ) , .B1( u0_u6_u4_n159 ) , .B2( u0_u6_u4_n184 ) );
  AND2_X1 u0_u6_u4_U80 (.A1( u0_u6_X_27 ) , .A2( u0_u6_X_30 ) , .ZN( u0_u6_u4_n103 ) );
  INV_X1 u0_u6_u4_U81 (.A( u0_u6_X_28 ) , .ZN( u0_u6_u4_n169 ) );
  INV_X1 u0_u6_u4_U82 (.A( u0_u6_X_29 ) , .ZN( u0_u6_u4_n168 ) );
  INV_X1 u0_u6_u4_U83 (.A( u0_u6_X_25 ) , .ZN( u0_u6_u4_n177 ) );
  INV_X1 u0_u6_u4_U84 (.A( u0_u6_X_27 ) , .ZN( u0_u6_u4_n176 ) );
  NAND4_X1 u0_u6_u4_U85 (.ZN( u0_out6_25 ) , .A4( u0_u6_u4_n139 ) , .A3( u0_u6_u4_n140 ) , .A2( u0_u6_u4_n141 ) , .A1( u0_u6_u4_n142 ) );
  OAI21_X1 u0_u6_u4_U86 (.B2( u0_u6_u4_n131 ) , .ZN( u0_u6_u4_n141 ) , .A( u0_u6_u4_n175 ) , .B1( u0_u6_u4_n183 ) );
  OAI21_X1 u0_u6_u4_U87 (.A( u0_u6_u4_n128 ) , .B2( u0_u6_u4_n129 ) , .B1( u0_u6_u4_n130 ) , .ZN( u0_u6_u4_n142 ) );
  NAND4_X1 u0_u6_u4_U88 (.ZN( u0_out6_14 ) , .A4( u0_u6_u4_n124 ) , .A3( u0_u6_u4_n125 ) , .A2( u0_u6_u4_n126 ) , .A1( u0_u6_u4_n127 ) );
  AOI22_X1 u0_u6_u4_U89 (.B2( u0_u6_u4_n117 ) , .ZN( u0_u6_u4_n126 ) , .A1( u0_u6_u4_n129 ) , .B1( u0_u6_u4_n152 ) , .A2( u0_u6_u4_n175 ) );
  AOI211_X1 u0_u6_u4_U9 (.B( u0_u6_u4_n136 ) , .A( u0_u6_u4_n137 ) , .C2( u0_u6_u4_n138 ) , .ZN( u0_u6_u4_n139 ) , .C1( u0_u6_u4_n182 ) );
  AOI22_X1 u0_u6_u4_U90 (.ZN( u0_u6_u4_n125 ) , .B2( u0_u6_u4_n131 ) , .A2( u0_u6_u4_n132 ) , .B1( u0_u6_u4_n138 ) , .A1( u0_u6_u4_n178 ) );
  NAND4_X1 u0_u6_u4_U91 (.ZN( u0_out6_8 ) , .A4( u0_u6_u4_n110 ) , .A3( u0_u6_u4_n111 ) , .A2( u0_u6_u4_n112 ) , .A1( u0_u6_u4_n186 ) );
  NAND2_X1 u0_u6_u4_U92 (.ZN( u0_u6_u4_n112 ) , .A2( u0_u6_u4_n130 ) , .A1( u0_u6_u4_n150 ) );
  AOI22_X1 u0_u6_u4_U93 (.ZN( u0_u6_u4_n111 ) , .B2( u0_u6_u4_n132 ) , .A1( u0_u6_u4_n152 ) , .B1( u0_u6_u4_n178 ) , .A2( u0_u6_u4_n97 ) );
  AOI22_X1 u0_u6_u4_U94 (.B2( u0_u6_u4_n149 ) , .B1( u0_u6_u4_n150 ) , .A2( u0_u6_u4_n151 ) , .A1( u0_u6_u4_n152 ) , .ZN( u0_u6_u4_n167 ) );
  NOR4_X1 u0_u6_u4_U95 (.A4( u0_u6_u4_n162 ) , .A3( u0_u6_u4_n163 ) , .A2( u0_u6_u4_n164 ) , .A1( u0_u6_u4_n165 ) , .ZN( u0_u6_u4_n166 ) );
  NAND3_X1 u0_u6_u4_U96 (.ZN( u0_out6_3 ) , .A3( u0_u6_u4_n166 ) , .A1( u0_u6_u4_n167 ) , .A2( u0_u6_u4_n186 ) );
  NAND3_X1 u0_u6_u4_U97 (.A3( u0_u6_u4_n146 ) , .A2( u0_u6_u4_n147 ) , .A1( u0_u6_u4_n148 ) , .ZN( u0_u6_u4_n149 ) );
  NAND3_X1 u0_u6_u4_U98 (.A3( u0_u6_u4_n143 ) , .A2( u0_u6_u4_n144 ) , .A1( u0_u6_u4_n145 ) , .ZN( u0_u6_u4_n151 ) );
  NAND3_X1 u0_u6_u4_U99 (.A3( u0_u6_u4_n121 ) , .ZN( u0_u6_u4_n122 ) , .A2( u0_u6_u4_n144 ) , .A1( u0_u6_u4_n154 ) );
  INV_X1 u0_u6_u5_U10 (.A( u0_u6_u5_n121 ) , .ZN( u0_u6_u5_n177 ) );
  NOR3_X1 u0_u6_u5_U100 (.A3( u0_u6_u5_n141 ) , .A1( u0_u6_u5_n142 ) , .ZN( u0_u6_u5_n143 ) , .A2( u0_u6_u5_n191 ) );
  NAND4_X1 u0_u6_u5_U101 (.ZN( u0_out6_4 ) , .A4( u0_u6_u5_n112 ) , .A2( u0_u6_u5_n113 ) , .A1( u0_u6_u5_n114 ) , .A3( u0_u6_u5_n195 ) );
  AOI211_X1 u0_u6_u5_U102 (.A( u0_u6_u5_n110 ) , .C1( u0_u6_u5_n111 ) , .ZN( u0_u6_u5_n112 ) , .B( u0_u6_u5_n118 ) , .C2( u0_u6_u5_n177 ) );
  AOI222_X1 u0_u6_u5_U103 (.ZN( u0_u6_u5_n113 ) , .A1( u0_u6_u5_n131 ) , .C1( u0_u6_u5_n148 ) , .B2( u0_u6_u5_n174 ) , .C2( u0_u6_u5_n178 ) , .A2( u0_u6_u5_n179 ) , .B1( u0_u6_u5_n99 ) );
  NAND3_X1 u0_u6_u5_U104 (.A2( u0_u6_u5_n154 ) , .A3( u0_u6_u5_n158 ) , .A1( u0_u6_u5_n161 ) , .ZN( u0_u6_u5_n99 ) );
  NOR2_X1 u0_u6_u5_U11 (.ZN( u0_u6_u5_n160 ) , .A2( u0_u6_u5_n173 ) , .A1( u0_u6_u5_n177 ) );
  INV_X1 u0_u6_u5_U12 (.A( u0_u6_u5_n150 ) , .ZN( u0_u6_u5_n174 ) );
  AOI21_X1 u0_u6_u5_U13 (.A( u0_u6_u5_n160 ) , .B2( u0_u6_u5_n161 ) , .ZN( u0_u6_u5_n162 ) , .B1( u0_u6_u5_n192 ) );
  INV_X1 u0_u6_u5_U14 (.A( u0_u6_u5_n159 ) , .ZN( u0_u6_u5_n192 ) );
  AOI21_X1 u0_u6_u5_U15 (.A( u0_u6_u5_n156 ) , .B2( u0_u6_u5_n157 ) , .B1( u0_u6_u5_n158 ) , .ZN( u0_u6_u5_n163 ) );
  AOI21_X1 u0_u6_u5_U16 (.B2( u0_u6_u5_n139 ) , .B1( u0_u6_u5_n140 ) , .ZN( u0_u6_u5_n141 ) , .A( u0_u6_u5_n150 ) );
  OAI21_X1 u0_u6_u5_U17 (.A( u0_u6_u5_n133 ) , .B2( u0_u6_u5_n134 ) , .B1( u0_u6_u5_n135 ) , .ZN( u0_u6_u5_n142 ) );
  OAI21_X1 u0_u6_u5_U18 (.ZN( u0_u6_u5_n133 ) , .B2( u0_u6_u5_n147 ) , .A( u0_u6_u5_n173 ) , .B1( u0_u6_u5_n188 ) );
  NAND2_X1 u0_u6_u5_U19 (.A2( u0_u6_u5_n119 ) , .A1( u0_u6_u5_n123 ) , .ZN( u0_u6_u5_n137 ) );
  INV_X1 u0_u6_u5_U20 (.A( u0_u6_u5_n155 ) , .ZN( u0_u6_u5_n194 ) );
  NAND2_X1 u0_u6_u5_U21 (.A1( u0_u6_u5_n121 ) , .ZN( u0_u6_u5_n132 ) , .A2( u0_u6_u5_n172 ) );
  NAND2_X1 u0_u6_u5_U22 (.A2( u0_u6_u5_n122 ) , .ZN( u0_u6_u5_n136 ) , .A1( u0_u6_u5_n154 ) );
  NAND2_X1 u0_u6_u5_U23 (.A2( u0_u6_u5_n119 ) , .A1( u0_u6_u5_n120 ) , .ZN( u0_u6_u5_n159 ) );
  INV_X1 u0_u6_u5_U24 (.A( u0_u6_u5_n156 ) , .ZN( u0_u6_u5_n175 ) );
  INV_X1 u0_u6_u5_U25 (.A( u0_u6_u5_n158 ) , .ZN( u0_u6_u5_n188 ) );
  INV_X1 u0_u6_u5_U26 (.A( u0_u6_u5_n152 ) , .ZN( u0_u6_u5_n179 ) );
  INV_X1 u0_u6_u5_U27 (.A( u0_u6_u5_n140 ) , .ZN( u0_u6_u5_n182 ) );
  INV_X1 u0_u6_u5_U28 (.A( u0_u6_u5_n151 ) , .ZN( u0_u6_u5_n183 ) );
  INV_X1 u0_u6_u5_U29 (.A( u0_u6_u5_n123 ) , .ZN( u0_u6_u5_n185 ) );
  NOR2_X1 u0_u6_u5_U3 (.ZN( u0_u6_u5_n134 ) , .A1( u0_u6_u5_n183 ) , .A2( u0_u6_u5_n190 ) );
  INV_X1 u0_u6_u5_U30 (.A( u0_u6_u5_n161 ) , .ZN( u0_u6_u5_n184 ) );
  INV_X1 u0_u6_u5_U31 (.A( u0_u6_u5_n139 ) , .ZN( u0_u6_u5_n189 ) );
  INV_X1 u0_u6_u5_U32 (.A( u0_u6_u5_n157 ) , .ZN( u0_u6_u5_n190 ) );
  INV_X1 u0_u6_u5_U33 (.A( u0_u6_u5_n120 ) , .ZN( u0_u6_u5_n193 ) );
  NAND2_X1 u0_u6_u5_U34 (.ZN( u0_u6_u5_n111 ) , .A1( u0_u6_u5_n140 ) , .A2( u0_u6_u5_n155 ) );
  INV_X1 u0_u6_u5_U35 (.A( u0_u6_u5_n117 ) , .ZN( u0_u6_u5_n196 ) );
  OAI221_X1 u0_u6_u5_U36 (.A( u0_u6_u5_n116 ) , .ZN( u0_u6_u5_n117 ) , .B2( u0_u6_u5_n119 ) , .C1( u0_u6_u5_n153 ) , .C2( u0_u6_u5_n158 ) , .B1( u0_u6_u5_n172 ) );
  AOI222_X1 u0_u6_u5_U37 (.ZN( u0_u6_u5_n116 ) , .B2( u0_u6_u5_n145 ) , .C1( u0_u6_u5_n148 ) , .A2( u0_u6_u5_n174 ) , .C2( u0_u6_u5_n177 ) , .B1( u0_u6_u5_n187 ) , .A1( u0_u6_u5_n193 ) );
  INV_X1 u0_u6_u5_U38 (.A( u0_u6_u5_n115 ) , .ZN( u0_u6_u5_n187 ) );
  NOR2_X1 u0_u6_u5_U39 (.ZN( u0_u6_u5_n100 ) , .A1( u0_u6_u5_n170 ) , .A2( u0_u6_u5_n180 ) );
  INV_X1 u0_u6_u5_U4 (.A( u0_u6_u5_n138 ) , .ZN( u0_u6_u5_n191 ) );
  AOI22_X1 u0_u6_u5_U40 (.B2( u0_u6_u5_n131 ) , .A2( u0_u6_u5_n146 ) , .ZN( u0_u6_u5_n169 ) , .B1( u0_u6_u5_n174 ) , .A1( u0_u6_u5_n185 ) );
  NOR2_X1 u0_u6_u5_U41 (.A1( u0_u6_u5_n146 ) , .ZN( u0_u6_u5_n150 ) , .A2( u0_u6_u5_n173 ) );
  AOI21_X1 u0_u6_u5_U42 (.A( u0_u6_u5_n118 ) , .B2( u0_u6_u5_n145 ) , .ZN( u0_u6_u5_n168 ) , .B1( u0_u6_u5_n186 ) );
  INV_X1 u0_u6_u5_U43 (.A( u0_u6_u5_n122 ) , .ZN( u0_u6_u5_n186 ) );
  NOR2_X1 u0_u6_u5_U44 (.A1( u0_u6_u5_n146 ) , .ZN( u0_u6_u5_n152 ) , .A2( u0_u6_u5_n176 ) );
  NOR2_X1 u0_u6_u5_U45 (.A1( u0_u6_u5_n115 ) , .ZN( u0_u6_u5_n118 ) , .A2( u0_u6_u5_n153 ) );
  NOR2_X1 u0_u6_u5_U46 (.A2( u0_u6_u5_n145 ) , .ZN( u0_u6_u5_n156 ) , .A1( u0_u6_u5_n174 ) );
  NOR2_X1 u0_u6_u5_U47 (.ZN( u0_u6_u5_n121 ) , .A2( u0_u6_u5_n145 ) , .A1( u0_u6_u5_n176 ) );
  AOI22_X1 u0_u6_u5_U48 (.ZN( u0_u6_u5_n114 ) , .A2( u0_u6_u5_n137 ) , .A1( u0_u6_u5_n145 ) , .B2( u0_u6_u5_n175 ) , .B1( u0_u6_u5_n193 ) );
  OAI211_X1 u0_u6_u5_U49 (.B( u0_u6_u5_n124 ) , .A( u0_u6_u5_n125 ) , .C2( u0_u6_u5_n126 ) , .C1( u0_u6_u5_n127 ) , .ZN( u0_u6_u5_n128 ) );
  OAI21_X1 u0_u6_u5_U5 (.B2( u0_u6_u5_n136 ) , .B1( u0_u6_u5_n137 ) , .ZN( u0_u6_u5_n138 ) , .A( u0_u6_u5_n177 ) );
  NOR3_X1 u0_u6_u5_U50 (.ZN( u0_u6_u5_n127 ) , .A1( u0_u6_u5_n136 ) , .A3( u0_u6_u5_n148 ) , .A2( u0_u6_u5_n182 ) );
  OAI21_X1 u0_u6_u5_U51 (.ZN( u0_u6_u5_n124 ) , .A( u0_u6_u5_n177 ) , .B2( u0_u6_u5_n183 ) , .B1( u0_u6_u5_n189 ) );
  OAI21_X1 u0_u6_u5_U52 (.ZN( u0_u6_u5_n125 ) , .A( u0_u6_u5_n174 ) , .B2( u0_u6_u5_n185 ) , .B1( u0_u6_u5_n190 ) );
  AOI21_X1 u0_u6_u5_U53 (.A( u0_u6_u5_n153 ) , .B2( u0_u6_u5_n154 ) , .B1( u0_u6_u5_n155 ) , .ZN( u0_u6_u5_n164 ) );
  AOI21_X1 u0_u6_u5_U54 (.ZN( u0_u6_u5_n110 ) , .B1( u0_u6_u5_n122 ) , .B2( u0_u6_u5_n139 ) , .A( u0_u6_u5_n153 ) );
  INV_X1 u0_u6_u5_U55 (.A( u0_u6_u5_n153 ) , .ZN( u0_u6_u5_n176 ) );
  INV_X1 u0_u6_u5_U56 (.A( u0_u6_u5_n126 ) , .ZN( u0_u6_u5_n173 ) );
  AND2_X1 u0_u6_u5_U57 (.A2( u0_u6_u5_n104 ) , .A1( u0_u6_u5_n107 ) , .ZN( u0_u6_u5_n147 ) );
  AND2_X1 u0_u6_u5_U58 (.A2( u0_u6_u5_n104 ) , .A1( u0_u6_u5_n108 ) , .ZN( u0_u6_u5_n148 ) );
  NAND2_X1 u0_u6_u5_U59 (.A1( u0_u6_u5_n105 ) , .A2( u0_u6_u5_n106 ) , .ZN( u0_u6_u5_n158 ) );
  INV_X1 u0_u6_u5_U6 (.A( u0_u6_u5_n135 ) , .ZN( u0_u6_u5_n178 ) );
  NAND2_X1 u0_u6_u5_U60 (.A2( u0_u6_u5_n108 ) , .A1( u0_u6_u5_n109 ) , .ZN( u0_u6_u5_n139 ) );
  NAND2_X1 u0_u6_u5_U61 (.A1( u0_u6_u5_n106 ) , .A2( u0_u6_u5_n108 ) , .ZN( u0_u6_u5_n119 ) );
  NAND2_X1 u0_u6_u5_U62 (.A2( u0_u6_u5_n103 ) , .A1( u0_u6_u5_n105 ) , .ZN( u0_u6_u5_n140 ) );
  NAND2_X1 u0_u6_u5_U63 (.A2( u0_u6_u5_n104 ) , .A1( u0_u6_u5_n105 ) , .ZN( u0_u6_u5_n155 ) );
  NAND2_X1 u0_u6_u5_U64 (.A2( u0_u6_u5_n106 ) , .A1( u0_u6_u5_n107 ) , .ZN( u0_u6_u5_n122 ) );
  NAND2_X1 u0_u6_u5_U65 (.A2( u0_u6_u5_n100 ) , .A1( u0_u6_u5_n106 ) , .ZN( u0_u6_u5_n115 ) );
  NAND2_X1 u0_u6_u5_U66 (.A2( u0_u6_u5_n100 ) , .A1( u0_u6_u5_n103 ) , .ZN( u0_u6_u5_n161 ) );
  NAND2_X1 u0_u6_u5_U67 (.A1( u0_u6_u5_n105 ) , .A2( u0_u6_u5_n109 ) , .ZN( u0_u6_u5_n154 ) );
  INV_X1 u0_u6_u5_U68 (.A( u0_u6_u5_n146 ) , .ZN( u0_u6_u5_n172 ) );
  NAND2_X1 u0_u6_u5_U69 (.A1( u0_u6_u5_n103 ) , .A2( u0_u6_u5_n108 ) , .ZN( u0_u6_u5_n123 ) );
  OAI22_X1 u0_u6_u5_U7 (.B2( u0_u6_u5_n149 ) , .B1( u0_u6_u5_n150 ) , .A2( u0_u6_u5_n151 ) , .A1( u0_u6_u5_n152 ) , .ZN( u0_u6_u5_n165 ) );
  NAND2_X1 u0_u6_u5_U70 (.A2( u0_u6_u5_n103 ) , .A1( u0_u6_u5_n107 ) , .ZN( u0_u6_u5_n151 ) );
  NAND2_X1 u0_u6_u5_U71 (.A2( u0_u6_u5_n107 ) , .A1( u0_u6_u5_n109 ) , .ZN( u0_u6_u5_n120 ) );
  NAND2_X1 u0_u6_u5_U72 (.A2( u0_u6_u5_n100 ) , .A1( u0_u6_u5_n109 ) , .ZN( u0_u6_u5_n157 ) );
  AND2_X1 u0_u6_u5_U73 (.A2( u0_u6_u5_n100 ) , .A1( u0_u6_u5_n104 ) , .ZN( u0_u6_u5_n131 ) );
  INV_X1 u0_u6_u5_U74 (.A( u0_u6_u5_n102 ) , .ZN( u0_u6_u5_n195 ) );
  OAI221_X1 u0_u6_u5_U75 (.A( u0_u6_u5_n101 ) , .ZN( u0_u6_u5_n102 ) , .C2( u0_u6_u5_n115 ) , .C1( u0_u6_u5_n126 ) , .B1( u0_u6_u5_n134 ) , .B2( u0_u6_u5_n160 ) );
  OAI21_X1 u0_u6_u5_U76 (.ZN( u0_u6_u5_n101 ) , .B1( u0_u6_u5_n137 ) , .A( u0_u6_u5_n146 ) , .B2( u0_u6_u5_n147 ) );
  NOR2_X1 u0_u6_u5_U77 (.A2( u0_u6_X_34 ) , .A1( u0_u6_X_35 ) , .ZN( u0_u6_u5_n145 ) );
  NOR2_X1 u0_u6_u5_U78 (.A2( u0_u6_X_34 ) , .ZN( u0_u6_u5_n146 ) , .A1( u0_u6_u5_n171 ) );
  NOR2_X1 u0_u6_u5_U79 (.A2( u0_u6_X_31 ) , .A1( u0_u6_X_32 ) , .ZN( u0_u6_u5_n103 ) );
  NOR3_X1 u0_u6_u5_U8 (.A2( u0_u6_u5_n147 ) , .A1( u0_u6_u5_n148 ) , .ZN( u0_u6_u5_n149 ) , .A3( u0_u6_u5_n194 ) );
  NOR2_X1 u0_u6_u5_U80 (.A2( u0_u6_X_36 ) , .ZN( u0_u6_u5_n105 ) , .A1( u0_u6_u5_n180 ) );
  NOR2_X1 u0_u6_u5_U81 (.A2( u0_u6_X_33 ) , .ZN( u0_u6_u5_n108 ) , .A1( u0_u6_u5_n170 ) );
  NOR2_X1 u0_u6_u5_U82 (.A2( u0_u6_X_33 ) , .A1( u0_u6_X_36 ) , .ZN( u0_u6_u5_n107 ) );
  NOR2_X1 u0_u6_u5_U83 (.A2( u0_u6_X_31 ) , .ZN( u0_u6_u5_n104 ) , .A1( u0_u6_u5_n181 ) );
  NAND2_X1 u0_u6_u5_U84 (.A2( u0_u6_X_34 ) , .A1( u0_u6_X_35 ) , .ZN( u0_u6_u5_n153 ) );
  NAND2_X1 u0_u6_u5_U85 (.A1( u0_u6_X_34 ) , .ZN( u0_u6_u5_n126 ) , .A2( u0_u6_u5_n171 ) );
  AND2_X1 u0_u6_u5_U86 (.A1( u0_u6_X_31 ) , .A2( u0_u6_X_32 ) , .ZN( u0_u6_u5_n106 ) );
  AND2_X1 u0_u6_u5_U87 (.A1( u0_u6_X_31 ) , .ZN( u0_u6_u5_n109 ) , .A2( u0_u6_u5_n181 ) );
  INV_X1 u0_u6_u5_U88 (.A( u0_u6_X_33 ) , .ZN( u0_u6_u5_n180 ) );
  INV_X1 u0_u6_u5_U89 (.A( u0_u6_X_35 ) , .ZN( u0_u6_u5_n171 ) );
  NOR2_X1 u0_u6_u5_U9 (.ZN( u0_u6_u5_n135 ) , .A1( u0_u6_u5_n173 ) , .A2( u0_u6_u5_n176 ) );
  INV_X1 u0_u6_u5_U90 (.A( u0_u6_X_36 ) , .ZN( u0_u6_u5_n170 ) );
  INV_X1 u0_u6_u5_U91 (.A( u0_u6_X_32 ) , .ZN( u0_u6_u5_n181 ) );
  NAND4_X1 u0_u6_u5_U92 (.ZN( u0_out6_29 ) , .A4( u0_u6_u5_n129 ) , .A3( u0_u6_u5_n130 ) , .A2( u0_u6_u5_n168 ) , .A1( u0_u6_u5_n196 ) );
  AOI221_X1 u0_u6_u5_U93 (.A( u0_u6_u5_n128 ) , .ZN( u0_u6_u5_n129 ) , .C2( u0_u6_u5_n132 ) , .B2( u0_u6_u5_n159 ) , .B1( u0_u6_u5_n176 ) , .C1( u0_u6_u5_n184 ) );
  AOI222_X1 u0_u6_u5_U94 (.ZN( u0_u6_u5_n130 ) , .A2( u0_u6_u5_n146 ) , .B1( u0_u6_u5_n147 ) , .C2( u0_u6_u5_n175 ) , .B2( u0_u6_u5_n179 ) , .A1( u0_u6_u5_n188 ) , .C1( u0_u6_u5_n194 ) );
  NAND4_X1 u0_u6_u5_U95 (.ZN( u0_out6_19 ) , .A4( u0_u6_u5_n166 ) , .A3( u0_u6_u5_n167 ) , .A2( u0_u6_u5_n168 ) , .A1( u0_u6_u5_n169 ) );
  AOI22_X1 u0_u6_u5_U96 (.B2( u0_u6_u5_n145 ) , .A2( u0_u6_u5_n146 ) , .ZN( u0_u6_u5_n167 ) , .B1( u0_u6_u5_n182 ) , .A1( u0_u6_u5_n189 ) );
  NOR4_X1 u0_u6_u5_U97 (.A4( u0_u6_u5_n162 ) , .A3( u0_u6_u5_n163 ) , .A2( u0_u6_u5_n164 ) , .A1( u0_u6_u5_n165 ) , .ZN( u0_u6_u5_n166 ) );
  NAND4_X1 u0_u6_u5_U98 (.ZN( u0_out6_11 ) , .A4( u0_u6_u5_n143 ) , .A3( u0_u6_u5_n144 ) , .A2( u0_u6_u5_n169 ) , .A1( u0_u6_u5_n196 ) );
  AOI22_X1 u0_u6_u5_U99 (.A2( u0_u6_u5_n132 ) , .ZN( u0_u6_u5_n144 ) , .B2( u0_u6_u5_n145 ) , .B1( u0_u6_u5_n184 ) , .A1( u0_u6_u5_n194 ) );
  AOI21_X1 u0_u6_u6_U10 (.ZN( u0_u6_u6_n106 ) , .A( u0_u6_u6_n142 ) , .B2( u0_u6_u6_n159 ) , .B1( u0_u6_u6_n164 ) );
  INV_X1 u0_u6_u6_U11 (.A( u0_u6_u6_n155 ) , .ZN( u0_u6_u6_n161 ) );
  INV_X1 u0_u6_u6_U12 (.A( u0_u6_u6_n128 ) , .ZN( u0_u6_u6_n164 ) );
  NAND2_X1 u0_u6_u6_U13 (.ZN( u0_u6_u6_n110 ) , .A1( u0_u6_u6_n122 ) , .A2( u0_u6_u6_n129 ) );
  NAND2_X1 u0_u6_u6_U14 (.ZN( u0_u6_u6_n124 ) , .A2( u0_u6_u6_n146 ) , .A1( u0_u6_u6_n148 ) );
  INV_X1 u0_u6_u6_U15 (.A( u0_u6_u6_n132 ) , .ZN( u0_u6_u6_n171 ) );
  AND2_X1 u0_u6_u6_U16 (.A1( u0_u6_u6_n100 ) , .ZN( u0_u6_u6_n130 ) , .A2( u0_u6_u6_n147 ) );
  INV_X1 u0_u6_u6_U17 (.A( u0_u6_u6_n127 ) , .ZN( u0_u6_u6_n173 ) );
  INV_X1 u0_u6_u6_U18 (.A( u0_u6_u6_n121 ) , .ZN( u0_u6_u6_n167 ) );
  INV_X1 u0_u6_u6_U19 (.A( u0_u6_u6_n100 ) , .ZN( u0_u6_u6_n169 ) );
  INV_X1 u0_u6_u6_U20 (.A( u0_u6_u6_n123 ) , .ZN( u0_u6_u6_n170 ) );
  INV_X1 u0_u6_u6_U21 (.A( u0_u6_u6_n113 ) , .ZN( u0_u6_u6_n168 ) );
  AND2_X1 u0_u6_u6_U22 (.A1( u0_u6_u6_n107 ) , .A2( u0_u6_u6_n119 ) , .ZN( u0_u6_u6_n133 ) );
  AND2_X1 u0_u6_u6_U23 (.A2( u0_u6_u6_n121 ) , .A1( u0_u6_u6_n122 ) , .ZN( u0_u6_u6_n131 ) );
  AND3_X1 u0_u6_u6_U24 (.ZN( u0_u6_u6_n120 ) , .A2( u0_u6_u6_n127 ) , .A1( u0_u6_u6_n132 ) , .A3( u0_u6_u6_n145 ) );
  INV_X1 u0_u6_u6_U25 (.A( u0_u6_u6_n146 ) , .ZN( u0_u6_u6_n163 ) );
  AOI222_X1 u0_u6_u6_U26 (.ZN( u0_u6_u6_n114 ) , .A1( u0_u6_u6_n118 ) , .A2( u0_u6_u6_n126 ) , .B2( u0_u6_u6_n151 ) , .C2( u0_u6_u6_n159 ) , .C1( u0_u6_u6_n168 ) , .B1( u0_u6_u6_n169 ) );
  NOR2_X1 u0_u6_u6_U27 (.A1( u0_u6_u6_n162 ) , .A2( u0_u6_u6_n165 ) , .ZN( u0_u6_u6_n98 ) );
  AOI211_X1 u0_u6_u6_U28 (.B( u0_u6_u6_n149 ) , .A( u0_u6_u6_n150 ) , .C2( u0_u6_u6_n151 ) , .C1( u0_u6_u6_n152 ) , .ZN( u0_u6_u6_n153 ) );
  AOI21_X1 u0_u6_u6_U29 (.B2( u0_u6_u6_n147 ) , .B1( u0_u6_u6_n148 ) , .ZN( u0_u6_u6_n149 ) , .A( u0_u6_u6_n158 ) );
  INV_X1 u0_u6_u6_U3 (.A( u0_u6_u6_n110 ) , .ZN( u0_u6_u6_n166 ) );
  AOI21_X1 u0_u6_u6_U30 (.A( u0_u6_u6_n144 ) , .B2( u0_u6_u6_n145 ) , .B1( u0_u6_u6_n146 ) , .ZN( u0_u6_u6_n150 ) );
  NAND2_X1 u0_u6_u6_U31 (.A2( u0_u6_u6_n143 ) , .ZN( u0_u6_u6_n152 ) , .A1( u0_u6_u6_n166 ) );
  NAND2_X1 u0_u6_u6_U32 (.A1( u0_u6_u6_n144 ) , .ZN( u0_u6_u6_n151 ) , .A2( u0_u6_u6_n158 ) );
  NAND2_X1 u0_u6_u6_U33 (.ZN( u0_u6_u6_n132 ) , .A1( u0_u6_u6_n91 ) , .A2( u0_u6_u6_n97 ) );
  AOI22_X1 u0_u6_u6_U34 (.B2( u0_u6_u6_n110 ) , .B1( u0_u6_u6_n111 ) , .A1( u0_u6_u6_n112 ) , .ZN( u0_u6_u6_n115 ) , .A2( u0_u6_u6_n161 ) );
  NAND4_X1 u0_u6_u6_U35 (.A3( u0_u6_u6_n109 ) , .ZN( u0_u6_u6_n112 ) , .A4( u0_u6_u6_n132 ) , .A2( u0_u6_u6_n147 ) , .A1( u0_u6_u6_n166 ) );
  NOR2_X1 u0_u6_u6_U36 (.ZN( u0_u6_u6_n109 ) , .A1( u0_u6_u6_n170 ) , .A2( u0_u6_u6_n173 ) );
  NOR2_X1 u0_u6_u6_U37 (.A2( u0_u6_u6_n126 ) , .ZN( u0_u6_u6_n155 ) , .A1( u0_u6_u6_n160 ) );
  NAND2_X1 u0_u6_u6_U38 (.ZN( u0_u6_u6_n146 ) , .A2( u0_u6_u6_n94 ) , .A1( u0_u6_u6_n99 ) );
  AOI211_X1 u0_u6_u6_U39 (.B( u0_u6_u6_n134 ) , .A( u0_u6_u6_n135 ) , .C1( u0_u6_u6_n136 ) , .ZN( u0_u6_u6_n137 ) , .C2( u0_u6_u6_n151 ) );
  AOI22_X1 u0_u6_u6_U4 (.B2( u0_u6_u6_n101 ) , .A1( u0_u6_u6_n102 ) , .ZN( u0_u6_u6_n103 ) , .B1( u0_u6_u6_n160 ) , .A2( u0_u6_u6_n161 ) );
  NAND4_X1 u0_u6_u6_U40 (.A4( u0_u6_u6_n127 ) , .A3( u0_u6_u6_n128 ) , .A2( u0_u6_u6_n129 ) , .A1( u0_u6_u6_n130 ) , .ZN( u0_u6_u6_n136 ) );
  AOI21_X1 u0_u6_u6_U41 (.B2( u0_u6_u6_n132 ) , .B1( u0_u6_u6_n133 ) , .ZN( u0_u6_u6_n134 ) , .A( u0_u6_u6_n158 ) );
  AOI21_X1 u0_u6_u6_U42 (.B1( u0_u6_u6_n131 ) , .ZN( u0_u6_u6_n135 ) , .A( u0_u6_u6_n144 ) , .B2( u0_u6_u6_n146 ) );
  INV_X1 u0_u6_u6_U43 (.A( u0_u6_u6_n111 ) , .ZN( u0_u6_u6_n158 ) );
  NAND2_X1 u0_u6_u6_U44 (.ZN( u0_u6_u6_n127 ) , .A1( u0_u6_u6_n91 ) , .A2( u0_u6_u6_n92 ) );
  NAND2_X1 u0_u6_u6_U45 (.ZN( u0_u6_u6_n129 ) , .A2( u0_u6_u6_n95 ) , .A1( u0_u6_u6_n96 ) );
  INV_X1 u0_u6_u6_U46 (.A( u0_u6_u6_n144 ) , .ZN( u0_u6_u6_n159 ) );
  NAND2_X1 u0_u6_u6_U47 (.ZN( u0_u6_u6_n145 ) , .A2( u0_u6_u6_n97 ) , .A1( u0_u6_u6_n98 ) );
  NAND2_X1 u0_u6_u6_U48 (.ZN( u0_u6_u6_n148 ) , .A2( u0_u6_u6_n92 ) , .A1( u0_u6_u6_n94 ) );
  NAND2_X1 u0_u6_u6_U49 (.ZN( u0_u6_u6_n108 ) , .A2( u0_u6_u6_n139 ) , .A1( u0_u6_u6_n144 ) );
  NOR2_X1 u0_u6_u6_U5 (.A1( u0_u6_u6_n118 ) , .ZN( u0_u6_u6_n143 ) , .A2( u0_u6_u6_n168 ) );
  NAND2_X1 u0_u6_u6_U50 (.ZN( u0_u6_u6_n121 ) , .A2( u0_u6_u6_n95 ) , .A1( u0_u6_u6_n97 ) );
  NAND2_X1 u0_u6_u6_U51 (.ZN( u0_u6_u6_n107 ) , .A2( u0_u6_u6_n92 ) , .A1( u0_u6_u6_n95 ) );
  AND2_X1 u0_u6_u6_U52 (.ZN( u0_u6_u6_n118 ) , .A2( u0_u6_u6_n91 ) , .A1( u0_u6_u6_n99 ) );
  NAND2_X1 u0_u6_u6_U53 (.ZN( u0_u6_u6_n147 ) , .A2( u0_u6_u6_n98 ) , .A1( u0_u6_u6_n99 ) );
  NAND2_X1 u0_u6_u6_U54 (.ZN( u0_u6_u6_n128 ) , .A1( u0_u6_u6_n94 ) , .A2( u0_u6_u6_n96 ) );
  NAND2_X1 u0_u6_u6_U55 (.ZN( u0_u6_u6_n119 ) , .A2( u0_u6_u6_n95 ) , .A1( u0_u6_u6_n99 ) );
  NAND2_X1 u0_u6_u6_U56 (.ZN( u0_u6_u6_n123 ) , .A2( u0_u6_u6_n91 ) , .A1( u0_u6_u6_n96 ) );
  NAND2_X1 u0_u6_u6_U57 (.ZN( u0_u6_u6_n100 ) , .A2( u0_u6_u6_n92 ) , .A1( u0_u6_u6_n98 ) );
  NAND2_X1 u0_u6_u6_U58 (.ZN( u0_u6_u6_n122 ) , .A1( u0_u6_u6_n94 ) , .A2( u0_u6_u6_n97 ) );
  INV_X1 u0_u6_u6_U59 (.A( u0_u6_u6_n139 ) , .ZN( u0_u6_u6_n160 ) );
  AOI21_X1 u0_u6_u6_U6 (.B1( u0_u6_u6_n107 ) , .B2( u0_u6_u6_n132 ) , .A( u0_u6_u6_n158 ) , .ZN( u0_u6_u6_n88 ) );
  NAND2_X1 u0_u6_u6_U60 (.ZN( u0_u6_u6_n113 ) , .A1( u0_u6_u6_n96 ) , .A2( u0_u6_u6_n98 ) );
  NOR2_X1 u0_u6_u6_U61 (.A2( u0_u6_X_40 ) , .A1( u0_u6_X_41 ) , .ZN( u0_u6_u6_n126 ) );
  NOR2_X1 u0_u6_u6_U62 (.A2( u0_u6_X_39 ) , .A1( u0_u6_X_42 ) , .ZN( u0_u6_u6_n92 ) );
  NOR2_X1 u0_u6_u6_U63 (.A2( u0_u6_X_39 ) , .A1( u0_u6_u6_n156 ) , .ZN( u0_u6_u6_n97 ) );
  NOR2_X1 u0_u6_u6_U64 (.A2( u0_u6_X_38 ) , .A1( u0_u6_u6_n165 ) , .ZN( u0_u6_u6_n95 ) );
  NOR2_X1 u0_u6_u6_U65 (.A2( u0_u6_X_41 ) , .ZN( u0_u6_u6_n111 ) , .A1( u0_u6_u6_n157 ) );
  NOR2_X1 u0_u6_u6_U66 (.A2( u0_u6_X_37 ) , .A1( u0_u6_u6_n162 ) , .ZN( u0_u6_u6_n94 ) );
  NOR2_X1 u0_u6_u6_U67 (.A2( u0_u6_X_37 ) , .A1( u0_u6_X_38 ) , .ZN( u0_u6_u6_n91 ) );
  NAND2_X1 u0_u6_u6_U68 (.A1( u0_u6_X_41 ) , .ZN( u0_u6_u6_n144 ) , .A2( u0_u6_u6_n157 ) );
  NAND2_X1 u0_u6_u6_U69 (.A2( u0_u6_X_40 ) , .A1( u0_u6_X_41 ) , .ZN( u0_u6_u6_n139 ) );
  OAI21_X1 u0_u6_u6_U7 (.A( u0_u6_u6_n159 ) , .B1( u0_u6_u6_n169 ) , .B2( u0_u6_u6_n173 ) , .ZN( u0_u6_u6_n90 ) );
  AND2_X1 u0_u6_u6_U70 (.A1( u0_u6_X_39 ) , .A2( u0_u6_u6_n156 ) , .ZN( u0_u6_u6_n96 ) );
  AND2_X1 u0_u6_u6_U71 (.A1( u0_u6_X_39 ) , .A2( u0_u6_X_42 ) , .ZN( u0_u6_u6_n99 ) );
  INV_X1 u0_u6_u6_U72 (.A( u0_u6_X_40 ) , .ZN( u0_u6_u6_n157 ) );
  INV_X1 u0_u6_u6_U73 (.A( u0_u6_X_37 ) , .ZN( u0_u6_u6_n165 ) );
  INV_X1 u0_u6_u6_U74 (.A( u0_u6_X_38 ) , .ZN( u0_u6_u6_n162 ) );
  INV_X1 u0_u6_u6_U75 (.A( u0_u6_X_42 ) , .ZN( u0_u6_u6_n156 ) );
  NAND4_X1 u0_u6_u6_U76 (.ZN( u0_out6_32 ) , .A4( u0_u6_u6_n103 ) , .A3( u0_u6_u6_n104 ) , .A2( u0_u6_u6_n105 ) , .A1( u0_u6_u6_n106 ) );
  AOI22_X1 u0_u6_u6_U77 (.ZN( u0_u6_u6_n104 ) , .A1( u0_u6_u6_n111 ) , .B1( u0_u6_u6_n124 ) , .B2( u0_u6_u6_n151 ) , .A2( u0_u6_u6_n93 ) );
  AOI22_X1 u0_u6_u6_U78 (.ZN( u0_u6_u6_n105 ) , .A2( u0_u6_u6_n108 ) , .A1( u0_u6_u6_n118 ) , .B2( u0_u6_u6_n126 ) , .B1( u0_u6_u6_n171 ) );
  NAND4_X1 u0_u6_u6_U79 (.ZN( u0_out6_12 ) , .A4( u0_u6_u6_n114 ) , .A3( u0_u6_u6_n115 ) , .A2( u0_u6_u6_n116 ) , .A1( u0_u6_u6_n117 ) );
  INV_X1 u0_u6_u6_U8 (.ZN( u0_u6_u6_n172 ) , .A( u0_u6_u6_n88 ) );
  OAI22_X1 u0_u6_u6_U80 (.B2( u0_u6_u6_n111 ) , .ZN( u0_u6_u6_n116 ) , .B1( u0_u6_u6_n126 ) , .A2( u0_u6_u6_n164 ) , .A1( u0_u6_u6_n167 ) );
  OAI21_X1 u0_u6_u6_U81 (.A( u0_u6_u6_n108 ) , .ZN( u0_u6_u6_n117 ) , .B2( u0_u6_u6_n141 ) , .B1( u0_u6_u6_n163 ) );
  OAI211_X1 u0_u6_u6_U82 (.ZN( u0_out6_22 ) , .B( u0_u6_u6_n137 ) , .A( u0_u6_u6_n138 ) , .C2( u0_u6_u6_n139 ) , .C1( u0_u6_u6_n140 ) );
  AOI22_X1 u0_u6_u6_U83 (.B1( u0_u6_u6_n124 ) , .A2( u0_u6_u6_n125 ) , .A1( u0_u6_u6_n126 ) , .ZN( u0_u6_u6_n138 ) , .B2( u0_u6_u6_n161 ) );
  AND4_X1 u0_u6_u6_U84 (.A3( u0_u6_u6_n119 ) , .A1( u0_u6_u6_n120 ) , .A4( u0_u6_u6_n129 ) , .ZN( u0_u6_u6_n140 ) , .A2( u0_u6_u6_n143 ) );
  OAI211_X1 u0_u6_u6_U85 (.ZN( u0_out6_7 ) , .B( u0_u6_u6_n153 ) , .C2( u0_u6_u6_n154 ) , .C1( u0_u6_u6_n155 ) , .A( u0_u6_u6_n174 ) );
  NOR3_X1 u0_u6_u6_U86 (.A1( u0_u6_u6_n141 ) , .ZN( u0_u6_u6_n154 ) , .A3( u0_u6_u6_n164 ) , .A2( u0_u6_u6_n171 ) );
  INV_X1 u0_u6_u6_U87 (.A( u0_u6_u6_n142 ) , .ZN( u0_u6_u6_n174 ) );
  NAND3_X1 u0_u6_u6_U88 (.A2( u0_u6_u6_n123 ) , .ZN( u0_u6_u6_n125 ) , .A1( u0_u6_u6_n130 ) , .A3( u0_u6_u6_n131 ) );
  NAND3_X1 u0_u6_u6_U89 (.A3( u0_u6_u6_n133 ) , .ZN( u0_u6_u6_n141 ) , .A1( u0_u6_u6_n145 ) , .A2( u0_u6_u6_n148 ) );
  AOI22_X1 u0_u6_u6_U9 (.A2( u0_u6_u6_n151 ) , .B2( u0_u6_u6_n161 ) , .A1( u0_u6_u6_n167 ) , .B1( u0_u6_u6_n170 ) , .ZN( u0_u6_u6_n89 ) );
  NAND3_X1 u0_u6_u6_U90 (.ZN( u0_u6_u6_n101 ) , .A3( u0_u6_u6_n107 ) , .A2( u0_u6_u6_n121 ) , .A1( u0_u6_u6_n127 ) );
  NAND3_X1 u0_u6_u6_U91 (.ZN( u0_u6_u6_n102 ) , .A3( u0_u6_u6_n130 ) , .A2( u0_u6_u6_n145 ) , .A1( u0_u6_u6_n166 ) );
  NAND3_X1 u0_u6_u6_U92 (.A3( u0_u6_u6_n113 ) , .A1( u0_u6_u6_n119 ) , .A2( u0_u6_u6_n123 ) , .ZN( u0_u6_u6_n93 ) );
  NAND3_X1 u0_u6_u6_U93 (.ZN( u0_u6_u6_n142 ) , .A2( u0_u6_u6_n172 ) , .A3( u0_u6_u6_n89 ) , .A1( u0_u6_u6_n90 ) );
  XOR2_X1 u0_u8_U10 (.B( u0_K9_45 ) , .A( u0_R7_30 ) , .Z( u0_u8_X_45 ) );
  XOR2_X1 u0_u8_U11 (.B( u0_K9_44 ) , .A( u0_R7_29 ) , .Z( u0_u8_X_44 ) );
  XOR2_X1 u0_u8_U12 (.B( u0_K9_43 ) , .A( u0_R7_28 ) , .Z( u0_u8_X_43 ) );
  XOR2_X1 u0_u8_U26 (.B( u0_K9_30 ) , .A( u0_R7_21 ) , .Z( u0_u8_X_30 ) );
  XOR2_X1 u0_u8_U28 (.B( u0_K9_29 ) , .A( u0_R7_20 ) , .Z( u0_u8_X_29 ) );
  XOR2_X1 u0_u8_U29 (.B( u0_K9_28 ) , .A( u0_R7_19 ) , .Z( u0_u8_X_28 ) );
  XOR2_X1 u0_u8_U30 (.B( u0_K9_27 ) , .A( u0_R7_18 ) , .Z( u0_u8_X_27 ) );
  XOR2_X1 u0_u8_U31 (.B( u0_K9_26 ) , .A( u0_R7_17 ) , .Z( u0_u8_X_26 ) );
  XOR2_X1 u0_u8_U32 (.B( u0_K9_25 ) , .A( u0_R7_16 ) , .Z( u0_u8_X_25 ) );
  XOR2_X1 u0_u8_U33 (.B( u0_K9_24 ) , .A( u0_R7_17 ) , .Z( u0_u8_X_24 ) );
  XOR2_X1 u0_u8_U34 (.B( u0_K9_23 ) , .A( u0_R7_16 ) , .Z( u0_u8_X_23 ) );
  XOR2_X1 u0_u8_U35 (.B( u0_K9_22 ) , .A( u0_R7_15 ) , .Z( u0_u8_X_22 ) );
  XOR2_X1 u0_u8_U36 (.B( u0_K9_21 ) , .A( u0_R7_14 ) , .Z( u0_u8_X_21 ) );
  XOR2_X1 u0_u8_U37 (.B( u0_K9_20 ) , .A( u0_R7_13 ) , .Z( u0_u8_X_20 ) );
  XOR2_X1 u0_u8_U39 (.B( u0_K9_19 ) , .A( u0_R7_12 ) , .Z( u0_u8_X_19 ) );
  XOR2_X1 u0_u8_U7 (.B( u0_K9_48 ) , .A( u0_R7_1 ) , .Z( u0_u8_X_48 ) );
  XOR2_X1 u0_u8_U8 (.B( u0_K9_47 ) , .A( u0_R7_32 ) , .Z( u0_u8_X_47 ) );
  XOR2_X1 u0_u8_U9 (.B( u0_K9_46 ) , .A( u0_R7_31 ) , .Z( u0_u8_X_46 ) );
  OAI22_X1 u0_u8_u3_U10 (.B1( u0_u8_u3_n113 ) , .A2( u0_u8_u3_n135 ) , .A1( u0_u8_u3_n150 ) , .B2( u0_u8_u3_n164 ) , .ZN( u0_u8_u3_n98 ) );
  OAI211_X1 u0_u8_u3_U11 (.B( u0_u8_u3_n106 ) , .ZN( u0_u8_u3_n119 ) , .C2( u0_u8_u3_n128 ) , .C1( u0_u8_u3_n167 ) , .A( u0_u8_u3_n181 ) );
  AOI221_X1 u0_u8_u3_U12 (.C1( u0_u8_u3_n105 ) , .ZN( u0_u8_u3_n106 ) , .A( u0_u8_u3_n131 ) , .B2( u0_u8_u3_n132 ) , .C2( u0_u8_u3_n133 ) , .B1( u0_u8_u3_n169 ) );
  INV_X1 u0_u8_u3_U13 (.ZN( u0_u8_u3_n181 ) , .A( u0_u8_u3_n98 ) );
  NAND2_X1 u0_u8_u3_U14 (.ZN( u0_u8_u3_n105 ) , .A2( u0_u8_u3_n130 ) , .A1( u0_u8_u3_n155 ) );
  AOI22_X1 u0_u8_u3_U15 (.B1( u0_u8_u3_n115 ) , .A2( u0_u8_u3_n116 ) , .ZN( u0_u8_u3_n123 ) , .B2( u0_u8_u3_n133 ) , .A1( u0_u8_u3_n169 ) );
  NAND2_X1 u0_u8_u3_U16 (.ZN( u0_u8_u3_n116 ) , .A2( u0_u8_u3_n151 ) , .A1( u0_u8_u3_n182 ) );
  NOR2_X1 u0_u8_u3_U17 (.ZN( u0_u8_u3_n126 ) , .A2( u0_u8_u3_n150 ) , .A1( u0_u8_u3_n164 ) );
  AOI21_X1 u0_u8_u3_U18 (.ZN( u0_u8_u3_n112 ) , .B2( u0_u8_u3_n146 ) , .B1( u0_u8_u3_n155 ) , .A( u0_u8_u3_n167 ) );
  NAND2_X1 u0_u8_u3_U19 (.A1( u0_u8_u3_n135 ) , .ZN( u0_u8_u3_n142 ) , .A2( u0_u8_u3_n164 ) );
  NAND2_X1 u0_u8_u3_U20 (.ZN( u0_u8_u3_n132 ) , .A2( u0_u8_u3_n152 ) , .A1( u0_u8_u3_n156 ) );
  AND2_X1 u0_u8_u3_U21 (.A2( u0_u8_u3_n113 ) , .A1( u0_u8_u3_n114 ) , .ZN( u0_u8_u3_n151 ) );
  INV_X1 u0_u8_u3_U22 (.A( u0_u8_u3_n133 ) , .ZN( u0_u8_u3_n165 ) );
  INV_X1 u0_u8_u3_U23 (.A( u0_u8_u3_n135 ) , .ZN( u0_u8_u3_n170 ) );
  NAND2_X1 u0_u8_u3_U24 (.A1( u0_u8_u3_n107 ) , .A2( u0_u8_u3_n108 ) , .ZN( u0_u8_u3_n140 ) );
  NAND2_X1 u0_u8_u3_U25 (.ZN( u0_u8_u3_n117 ) , .A1( u0_u8_u3_n124 ) , .A2( u0_u8_u3_n148 ) );
  NAND2_X1 u0_u8_u3_U26 (.ZN( u0_u8_u3_n143 ) , .A1( u0_u8_u3_n165 ) , .A2( u0_u8_u3_n167 ) );
  INV_X1 u0_u8_u3_U27 (.A( u0_u8_u3_n130 ) , .ZN( u0_u8_u3_n177 ) );
  INV_X1 u0_u8_u3_U28 (.A( u0_u8_u3_n128 ) , .ZN( u0_u8_u3_n176 ) );
  INV_X1 u0_u8_u3_U29 (.A( u0_u8_u3_n155 ) , .ZN( u0_u8_u3_n174 ) );
  INV_X1 u0_u8_u3_U3 (.A( u0_u8_u3_n129 ) , .ZN( u0_u8_u3_n183 ) );
  INV_X1 u0_u8_u3_U30 (.A( u0_u8_u3_n139 ) , .ZN( u0_u8_u3_n185 ) );
  NOR2_X1 u0_u8_u3_U31 (.ZN( u0_u8_u3_n135 ) , .A2( u0_u8_u3_n141 ) , .A1( u0_u8_u3_n169 ) );
  OAI222_X1 u0_u8_u3_U32 (.C2( u0_u8_u3_n107 ) , .A2( u0_u8_u3_n108 ) , .B1( u0_u8_u3_n135 ) , .ZN( u0_u8_u3_n138 ) , .B2( u0_u8_u3_n146 ) , .C1( u0_u8_u3_n154 ) , .A1( u0_u8_u3_n164 ) );
  NOR4_X1 u0_u8_u3_U33 (.A4( u0_u8_u3_n157 ) , .A3( u0_u8_u3_n158 ) , .A2( u0_u8_u3_n159 ) , .A1( u0_u8_u3_n160 ) , .ZN( u0_u8_u3_n161 ) );
  AOI21_X1 u0_u8_u3_U34 (.B2( u0_u8_u3_n152 ) , .B1( u0_u8_u3_n153 ) , .ZN( u0_u8_u3_n158 ) , .A( u0_u8_u3_n164 ) );
  AOI21_X1 u0_u8_u3_U35 (.A( u0_u8_u3_n149 ) , .B2( u0_u8_u3_n150 ) , .B1( u0_u8_u3_n151 ) , .ZN( u0_u8_u3_n159 ) );
  AOI21_X1 u0_u8_u3_U36 (.A( u0_u8_u3_n154 ) , .B2( u0_u8_u3_n155 ) , .B1( u0_u8_u3_n156 ) , .ZN( u0_u8_u3_n157 ) );
  AOI211_X1 u0_u8_u3_U37 (.ZN( u0_u8_u3_n109 ) , .A( u0_u8_u3_n119 ) , .C2( u0_u8_u3_n129 ) , .B( u0_u8_u3_n138 ) , .C1( u0_u8_u3_n141 ) );
  AOI211_X1 u0_u8_u3_U38 (.B( u0_u8_u3_n119 ) , .A( u0_u8_u3_n120 ) , .C2( u0_u8_u3_n121 ) , .ZN( u0_u8_u3_n122 ) , .C1( u0_u8_u3_n179 ) );
  INV_X1 u0_u8_u3_U39 (.A( u0_u8_u3_n156 ) , .ZN( u0_u8_u3_n179 ) );
  INV_X1 u0_u8_u3_U4 (.A( u0_u8_u3_n140 ) , .ZN( u0_u8_u3_n182 ) );
  OAI22_X1 u0_u8_u3_U40 (.B1( u0_u8_u3_n118 ) , .ZN( u0_u8_u3_n120 ) , .A1( u0_u8_u3_n135 ) , .B2( u0_u8_u3_n154 ) , .A2( u0_u8_u3_n178 ) );
  AND3_X1 u0_u8_u3_U41 (.ZN( u0_u8_u3_n118 ) , .A2( u0_u8_u3_n124 ) , .A1( u0_u8_u3_n144 ) , .A3( u0_u8_u3_n152 ) );
  INV_X1 u0_u8_u3_U42 (.A( u0_u8_u3_n121 ) , .ZN( u0_u8_u3_n164 ) );
  NAND2_X1 u0_u8_u3_U43 (.ZN( u0_u8_u3_n133 ) , .A1( u0_u8_u3_n154 ) , .A2( u0_u8_u3_n164 ) );
  OAI211_X1 u0_u8_u3_U44 (.B( u0_u8_u3_n127 ) , .ZN( u0_u8_u3_n139 ) , .C1( u0_u8_u3_n150 ) , .C2( u0_u8_u3_n154 ) , .A( u0_u8_u3_n184 ) );
  INV_X1 u0_u8_u3_U45 (.A( u0_u8_u3_n125 ) , .ZN( u0_u8_u3_n184 ) );
  AOI221_X1 u0_u8_u3_U46 (.A( u0_u8_u3_n126 ) , .ZN( u0_u8_u3_n127 ) , .C2( u0_u8_u3_n132 ) , .C1( u0_u8_u3_n169 ) , .B2( u0_u8_u3_n170 ) , .B1( u0_u8_u3_n174 ) );
  OAI22_X1 u0_u8_u3_U47 (.A1( u0_u8_u3_n124 ) , .ZN( u0_u8_u3_n125 ) , .B2( u0_u8_u3_n145 ) , .A2( u0_u8_u3_n165 ) , .B1( u0_u8_u3_n167 ) );
  NOR2_X1 u0_u8_u3_U48 (.A1( u0_u8_u3_n113 ) , .ZN( u0_u8_u3_n131 ) , .A2( u0_u8_u3_n154 ) );
  NAND2_X1 u0_u8_u3_U49 (.A1( u0_u8_u3_n103 ) , .ZN( u0_u8_u3_n150 ) , .A2( u0_u8_u3_n99 ) );
  INV_X1 u0_u8_u3_U5 (.A( u0_u8_u3_n117 ) , .ZN( u0_u8_u3_n178 ) );
  NAND2_X1 u0_u8_u3_U50 (.A2( u0_u8_u3_n102 ) , .ZN( u0_u8_u3_n155 ) , .A1( u0_u8_u3_n97 ) );
  INV_X1 u0_u8_u3_U51 (.A( u0_u8_u3_n141 ) , .ZN( u0_u8_u3_n167 ) );
  AOI21_X1 u0_u8_u3_U52 (.B2( u0_u8_u3_n114 ) , .B1( u0_u8_u3_n146 ) , .A( u0_u8_u3_n154 ) , .ZN( u0_u8_u3_n94 ) );
  AOI21_X1 u0_u8_u3_U53 (.ZN( u0_u8_u3_n110 ) , .B2( u0_u8_u3_n142 ) , .B1( u0_u8_u3_n186 ) , .A( u0_u8_u3_n95 ) );
  INV_X1 u0_u8_u3_U54 (.A( u0_u8_u3_n145 ) , .ZN( u0_u8_u3_n186 ) );
  AOI21_X1 u0_u8_u3_U55 (.B1( u0_u8_u3_n124 ) , .A( u0_u8_u3_n149 ) , .B2( u0_u8_u3_n155 ) , .ZN( u0_u8_u3_n95 ) );
  INV_X1 u0_u8_u3_U56 (.A( u0_u8_u3_n149 ) , .ZN( u0_u8_u3_n169 ) );
  NAND2_X1 u0_u8_u3_U57 (.ZN( u0_u8_u3_n124 ) , .A1( u0_u8_u3_n96 ) , .A2( u0_u8_u3_n97 ) );
  NAND2_X1 u0_u8_u3_U58 (.A2( u0_u8_u3_n100 ) , .ZN( u0_u8_u3_n146 ) , .A1( u0_u8_u3_n96 ) );
  NAND2_X1 u0_u8_u3_U59 (.A1( u0_u8_u3_n101 ) , .ZN( u0_u8_u3_n145 ) , .A2( u0_u8_u3_n99 ) );
  AOI221_X1 u0_u8_u3_U6 (.A( u0_u8_u3_n131 ) , .C2( u0_u8_u3_n132 ) , .C1( u0_u8_u3_n133 ) , .ZN( u0_u8_u3_n134 ) , .B1( u0_u8_u3_n143 ) , .B2( u0_u8_u3_n177 ) );
  NAND2_X1 u0_u8_u3_U60 (.A1( u0_u8_u3_n100 ) , .ZN( u0_u8_u3_n156 ) , .A2( u0_u8_u3_n99 ) );
  NAND2_X1 u0_u8_u3_U61 (.A2( u0_u8_u3_n101 ) , .A1( u0_u8_u3_n104 ) , .ZN( u0_u8_u3_n148 ) );
  NAND2_X1 u0_u8_u3_U62 (.A1( u0_u8_u3_n100 ) , .A2( u0_u8_u3_n102 ) , .ZN( u0_u8_u3_n128 ) );
  NAND2_X1 u0_u8_u3_U63 (.A2( u0_u8_u3_n101 ) , .A1( u0_u8_u3_n102 ) , .ZN( u0_u8_u3_n152 ) );
  NAND2_X1 u0_u8_u3_U64 (.A2( u0_u8_u3_n101 ) , .ZN( u0_u8_u3_n114 ) , .A1( u0_u8_u3_n96 ) );
  NAND2_X1 u0_u8_u3_U65 (.ZN( u0_u8_u3_n107 ) , .A1( u0_u8_u3_n97 ) , .A2( u0_u8_u3_n99 ) );
  NAND2_X1 u0_u8_u3_U66 (.A2( u0_u8_u3_n100 ) , .A1( u0_u8_u3_n104 ) , .ZN( u0_u8_u3_n113 ) );
  NAND2_X1 u0_u8_u3_U67 (.A1( u0_u8_u3_n104 ) , .ZN( u0_u8_u3_n153 ) , .A2( u0_u8_u3_n97 ) );
  NAND2_X1 u0_u8_u3_U68 (.A2( u0_u8_u3_n103 ) , .A1( u0_u8_u3_n104 ) , .ZN( u0_u8_u3_n130 ) );
  NAND2_X1 u0_u8_u3_U69 (.A2( u0_u8_u3_n103 ) , .ZN( u0_u8_u3_n144 ) , .A1( u0_u8_u3_n96 ) );
  OAI22_X1 u0_u8_u3_U7 (.B2( u0_u8_u3_n147 ) , .A2( u0_u8_u3_n148 ) , .ZN( u0_u8_u3_n160 ) , .B1( u0_u8_u3_n165 ) , .A1( u0_u8_u3_n168 ) );
  NAND2_X1 u0_u8_u3_U70 (.A1( u0_u8_u3_n102 ) , .A2( u0_u8_u3_n103 ) , .ZN( u0_u8_u3_n108 ) );
  NOR2_X1 u0_u8_u3_U71 (.A2( u0_u8_X_19 ) , .A1( u0_u8_X_20 ) , .ZN( u0_u8_u3_n99 ) );
  NOR2_X1 u0_u8_u3_U72 (.A2( u0_u8_X_21 ) , .A1( u0_u8_X_24 ) , .ZN( u0_u8_u3_n103 ) );
  NOR2_X1 u0_u8_u3_U73 (.A2( u0_u8_X_24 ) , .A1( u0_u8_u3_n171 ) , .ZN( u0_u8_u3_n97 ) );
  NOR2_X1 u0_u8_u3_U74 (.A2( u0_u8_X_23 ) , .ZN( u0_u8_u3_n141 ) , .A1( u0_u8_u3_n166 ) );
  NOR2_X1 u0_u8_u3_U75 (.A2( u0_u8_X_19 ) , .A1( u0_u8_u3_n172 ) , .ZN( u0_u8_u3_n96 ) );
  NAND2_X1 u0_u8_u3_U76 (.A1( u0_u8_X_22 ) , .A2( u0_u8_X_23 ) , .ZN( u0_u8_u3_n154 ) );
  NAND2_X1 u0_u8_u3_U77 (.A1( u0_u8_X_23 ) , .ZN( u0_u8_u3_n149 ) , .A2( u0_u8_u3_n166 ) );
  NOR2_X1 u0_u8_u3_U78 (.A2( u0_u8_X_22 ) , .A1( u0_u8_X_23 ) , .ZN( u0_u8_u3_n121 ) );
  AND2_X1 u0_u8_u3_U79 (.A1( u0_u8_X_24 ) , .ZN( u0_u8_u3_n101 ) , .A2( u0_u8_u3_n171 ) );
  AND3_X1 u0_u8_u3_U8 (.A3( u0_u8_u3_n144 ) , .A2( u0_u8_u3_n145 ) , .A1( u0_u8_u3_n146 ) , .ZN( u0_u8_u3_n147 ) );
  AND2_X1 u0_u8_u3_U80 (.A1( u0_u8_X_19 ) , .ZN( u0_u8_u3_n102 ) , .A2( u0_u8_u3_n172 ) );
  AND2_X1 u0_u8_u3_U81 (.A1( u0_u8_X_21 ) , .A2( u0_u8_X_24 ) , .ZN( u0_u8_u3_n100 ) );
  AND2_X1 u0_u8_u3_U82 (.A2( u0_u8_X_19 ) , .A1( u0_u8_X_20 ) , .ZN( u0_u8_u3_n104 ) );
  INV_X1 u0_u8_u3_U83 (.A( u0_u8_X_22 ) , .ZN( u0_u8_u3_n166 ) );
  INV_X1 u0_u8_u3_U84 (.A( u0_u8_X_21 ) , .ZN( u0_u8_u3_n171 ) );
  INV_X1 u0_u8_u3_U85 (.A( u0_u8_X_20 ) , .ZN( u0_u8_u3_n172 ) );
  OR4_X1 u0_u8_u3_U86 (.ZN( u0_out8_10 ) , .A4( u0_u8_u3_n136 ) , .A3( u0_u8_u3_n137 ) , .A1( u0_u8_u3_n138 ) , .A2( u0_u8_u3_n139 ) );
  OAI222_X1 u0_u8_u3_U87 (.C1( u0_u8_u3_n128 ) , .ZN( u0_u8_u3_n137 ) , .B1( u0_u8_u3_n148 ) , .A2( u0_u8_u3_n150 ) , .B2( u0_u8_u3_n154 ) , .C2( u0_u8_u3_n164 ) , .A1( u0_u8_u3_n167 ) );
  OAI221_X1 u0_u8_u3_U88 (.A( u0_u8_u3_n134 ) , .B2( u0_u8_u3_n135 ) , .ZN( u0_u8_u3_n136 ) , .C1( u0_u8_u3_n149 ) , .B1( u0_u8_u3_n151 ) , .C2( u0_u8_u3_n183 ) );
  NAND4_X1 u0_u8_u3_U89 (.ZN( u0_out8_26 ) , .A4( u0_u8_u3_n109 ) , .A3( u0_u8_u3_n110 ) , .A2( u0_u8_u3_n111 ) , .A1( u0_u8_u3_n173 ) );
  INV_X1 u0_u8_u3_U9 (.A( u0_u8_u3_n143 ) , .ZN( u0_u8_u3_n168 ) );
  INV_X1 u0_u8_u3_U90 (.ZN( u0_u8_u3_n173 ) , .A( u0_u8_u3_n94 ) );
  OAI21_X1 u0_u8_u3_U91 (.ZN( u0_u8_u3_n111 ) , .B2( u0_u8_u3_n117 ) , .A( u0_u8_u3_n133 ) , .B1( u0_u8_u3_n176 ) );
  NAND4_X1 u0_u8_u3_U92 (.ZN( u0_out8_20 ) , .A4( u0_u8_u3_n122 ) , .A3( u0_u8_u3_n123 ) , .A1( u0_u8_u3_n175 ) , .A2( u0_u8_u3_n180 ) );
  INV_X1 u0_u8_u3_U93 (.A( u0_u8_u3_n126 ) , .ZN( u0_u8_u3_n180 ) );
  INV_X1 u0_u8_u3_U94 (.A( u0_u8_u3_n112 ) , .ZN( u0_u8_u3_n175 ) );
  NAND4_X1 u0_u8_u3_U95 (.ZN( u0_out8_1 ) , .A4( u0_u8_u3_n161 ) , .A3( u0_u8_u3_n162 ) , .A2( u0_u8_u3_n163 ) , .A1( u0_u8_u3_n185 ) );
  NAND2_X1 u0_u8_u3_U96 (.ZN( u0_u8_u3_n163 ) , .A2( u0_u8_u3_n170 ) , .A1( u0_u8_u3_n176 ) );
  AOI22_X1 u0_u8_u3_U97 (.B2( u0_u8_u3_n140 ) , .B1( u0_u8_u3_n141 ) , .A2( u0_u8_u3_n142 ) , .ZN( u0_u8_u3_n162 ) , .A1( u0_u8_u3_n177 ) );
  NAND3_X1 u0_u8_u3_U98 (.A1( u0_u8_u3_n114 ) , .ZN( u0_u8_u3_n115 ) , .A2( u0_u8_u3_n145 ) , .A3( u0_u8_u3_n153 ) );
  NAND3_X1 u0_u8_u3_U99 (.ZN( u0_u8_u3_n129 ) , .A2( u0_u8_u3_n144 ) , .A1( u0_u8_u3_n153 ) , .A3( u0_u8_u3_n182 ) );
  OAI22_X1 u0_u8_u4_U10 (.B2( u0_u8_u4_n135 ) , .ZN( u0_u8_u4_n137 ) , .B1( u0_u8_u4_n153 ) , .A1( u0_u8_u4_n155 ) , .A2( u0_u8_u4_n171 ) );
  AND3_X1 u0_u8_u4_U11 (.A2( u0_u8_u4_n134 ) , .ZN( u0_u8_u4_n135 ) , .A3( u0_u8_u4_n145 ) , .A1( u0_u8_u4_n157 ) );
  NAND2_X1 u0_u8_u4_U12 (.ZN( u0_u8_u4_n132 ) , .A2( u0_u8_u4_n170 ) , .A1( u0_u8_u4_n173 ) );
  AOI21_X1 u0_u8_u4_U13 (.B2( u0_u8_u4_n160 ) , .B1( u0_u8_u4_n161 ) , .ZN( u0_u8_u4_n162 ) , .A( u0_u8_u4_n170 ) );
  AOI21_X1 u0_u8_u4_U14 (.ZN( u0_u8_u4_n107 ) , .B2( u0_u8_u4_n143 ) , .A( u0_u8_u4_n174 ) , .B1( u0_u8_u4_n184 ) );
  AOI21_X1 u0_u8_u4_U15 (.B2( u0_u8_u4_n158 ) , .B1( u0_u8_u4_n159 ) , .ZN( u0_u8_u4_n163 ) , .A( u0_u8_u4_n174 ) );
  AOI21_X1 u0_u8_u4_U16 (.A( u0_u8_u4_n153 ) , .B2( u0_u8_u4_n154 ) , .B1( u0_u8_u4_n155 ) , .ZN( u0_u8_u4_n165 ) );
  AOI21_X1 u0_u8_u4_U17 (.A( u0_u8_u4_n156 ) , .B2( u0_u8_u4_n157 ) , .ZN( u0_u8_u4_n164 ) , .B1( u0_u8_u4_n184 ) );
  INV_X1 u0_u8_u4_U18 (.A( u0_u8_u4_n138 ) , .ZN( u0_u8_u4_n170 ) );
  AND2_X1 u0_u8_u4_U19 (.A2( u0_u8_u4_n120 ) , .ZN( u0_u8_u4_n155 ) , .A1( u0_u8_u4_n160 ) );
  INV_X1 u0_u8_u4_U20 (.A( u0_u8_u4_n156 ) , .ZN( u0_u8_u4_n175 ) );
  NAND2_X1 u0_u8_u4_U21 (.A2( u0_u8_u4_n118 ) , .ZN( u0_u8_u4_n131 ) , .A1( u0_u8_u4_n147 ) );
  NAND2_X1 u0_u8_u4_U22 (.A1( u0_u8_u4_n119 ) , .A2( u0_u8_u4_n120 ) , .ZN( u0_u8_u4_n130 ) );
  NAND2_X1 u0_u8_u4_U23 (.ZN( u0_u8_u4_n117 ) , .A2( u0_u8_u4_n118 ) , .A1( u0_u8_u4_n148 ) );
  NAND2_X1 u0_u8_u4_U24 (.ZN( u0_u8_u4_n129 ) , .A1( u0_u8_u4_n134 ) , .A2( u0_u8_u4_n148 ) );
  AND3_X1 u0_u8_u4_U25 (.A1( u0_u8_u4_n119 ) , .A2( u0_u8_u4_n143 ) , .A3( u0_u8_u4_n154 ) , .ZN( u0_u8_u4_n161 ) );
  AND2_X1 u0_u8_u4_U26 (.A1( u0_u8_u4_n145 ) , .A2( u0_u8_u4_n147 ) , .ZN( u0_u8_u4_n159 ) );
  OR3_X1 u0_u8_u4_U27 (.A3( u0_u8_u4_n114 ) , .A2( u0_u8_u4_n115 ) , .A1( u0_u8_u4_n116 ) , .ZN( u0_u8_u4_n136 ) );
  AOI21_X1 u0_u8_u4_U28 (.A( u0_u8_u4_n113 ) , .ZN( u0_u8_u4_n116 ) , .B2( u0_u8_u4_n173 ) , .B1( u0_u8_u4_n174 ) );
  AOI21_X1 u0_u8_u4_U29 (.ZN( u0_u8_u4_n115 ) , .B2( u0_u8_u4_n145 ) , .B1( u0_u8_u4_n146 ) , .A( u0_u8_u4_n156 ) );
  NOR2_X1 u0_u8_u4_U3 (.ZN( u0_u8_u4_n121 ) , .A1( u0_u8_u4_n181 ) , .A2( u0_u8_u4_n182 ) );
  OAI22_X1 u0_u8_u4_U30 (.ZN( u0_u8_u4_n114 ) , .A2( u0_u8_u4_n121 ) , .B1( u0_u8_u4_n160 ) , .B2( u0_u8_u4_n170 ) , .A1( u0_u8_u4_n171 ) );
  INV_X1 u0_u8_u4_U31 (.A( u0_u8_u4_n158 ) , .ZN( u0_u8_u4_n182 ) );
  INV_X1 u0_u8_u4_U32 (.ZN( u0_u8_u4_n181 ) , .A( u0_u8_u4_n96 ) );
  INV_X1 u0_u8_u4_U33 (.A( u0_u8_u4_n144 ) , .ZN( u0_u8_u4_n179 ) );
  INV_X1 u0_u8_u4_U34 (.A( u0_u8_u4_n157 ) , .ZN( u0_u8_u4_n178 ) );
  NAND2_X1 u0_u8_u4_U35 (.A2( u0_u8_u4_n154 ) , .A1( u0_u8_u4_n96 ) , .ZN( u0_u8_u4_n97 ) );
  INV_X1 u0_u8_u4_U36 (.ZN( u0_u8_u4_n186 ) , .A( u0_u8_u4_n95 ) );
  OAI221_X1 u0_u8_u4_U37 (.C1( u0_u8_u4_n134 ) , .B1( u0_u8_u4_n158 ) , .B2( u0_u8_u4_n171 ) , .C2( u0_u8_u4_n173 ) , .A( u0_u8_u4_n94 ) , .ZN( u0_u8_u4_n95 ) );
  AOI222_X1 u0_u8_u4_U38 (.B2( u0_u8_u4_n132 ) , .A1( u0_u8_u4_n138 ) , .C2( u0_u8_u4_n175 ) , .A2( u0_u8_u4_n179 ) , .C1( u0_u8_u4_n181 ) , .B1( u0_u8_u4_n185 ) , .ZN( u0_u8_u4_n94 ) );
  INV_X1 u0_u8_u4_U39 (.A( u0_u8_u4_n113 ) , .ZN( u0_u8_u4_n185 ) );
  INV_X1 u0_u8_u4_U4 (.A( u0_u8_u4_n117 ) , .ZN( u0_u8_u4_n184 ) );
  INV_X1 u0_u8_u4_U40 (.A( u0_u8_u4_n143 ) , .ZN( u0_u8_u4_n183 ) );
  NOR2_X1 u0_u8_u4_U41 (.ZN( u0_u8_u4_n138 ) , .A1( u0_u8_u4_n168 ) , .A2( u0_u8_u4_n169 ) );
  NOR2_X1 u0_u8_u4_U42 (.A1( u0_u8_u4_n150 ) , .A2( u0_u8_u4_n152 ) , .ZN( u0_u8_u4_n153 ) );
  NOR2_X1 u0_u8_u4_U43 (.A2( u0_u8_u4_n128 ) , .A1( u0_u8_u4_n138 ) , .ZN( u0_u8_u4_n156 ) );
  AOI22_X1 u0_u8_u4_U44 (.B2( u0_u8_u4_n122 ) , .A1( u0_u8_u4_n123 ) , .ZN( u0_u8_u4_n124 ) , .B1( u0_u8_u4_n128 ) , .A2( u0_u8_u4_n172 ) );
  INV_X1 u0_u8_u4_U45 (.A( u0_u8_u4_n153 ) , .ZN( u0_u8_u4_n172 ) );
  NAND2_X1 u0_u8_u4_U46 (.A2( u0_u8_u4_n120 ) , .ZN( u0_u8_u4_n123 ) , .A1( u0_u8_u4_n161 ) );
  AOI22_X1 u0_u8_u4_U47 (.B2( u0_u8_u4_n132 ) , .A2( u0_u8_u4_n133 ) , .ZN( u0_u8_u4_n140 ) , .A1( u0_u8_u4_n150 ) , .B1( u0_u8_u4_n179 ) );
  NAND2_X1 u0_u8_u4_U48 (.ZN( u0_u8_u4_n133 ) , .A2( u0_u8_u4_n146 ) , .A1( u0_u8_u4_n154 ) );
  NAND2_X1 u0_u8_u4_U49 (.A1( u0_u8_u4_n103 ) , .ZN( u0_u8_u4_n154 ) , .A2( u0_u8_u4_n98 ) );
  NOR4_X1 u0_u8_u4_U5 (.A4( u0_u8_u4_n106 ) , .A3( u0_u8_u4_n107 ) , .A2( u0_u8_u4_n108 ) , .A1( u0_u8_u4_n109 ) , .ZN( u0_u8_u4_n110 ) );
  NAND2_X1 u0_u8_u4_U50 (.A1( u0_u8_u4_n101 ) , .ZN( u0_u8_u4_n158 ) , .A2( u0_u8_u4_n99 ) );
  AOI21_X1 u0_u8_u4_U51 (.ZN( u0_u8_u4_n127 ) , .A( u0_u8_u4_n136 ) , .B2( u0_u8_u4_n150 ) , .B1( u0_u8_u4_n180 ) );
  INV_X1 u0_u8_u4_U52 (.A( u0_u8_u4_n160 ) , .ZN( u0_u8_u4_n180 ) );
  NAND2_X1 u0_u8_u4_U53 (.A2( u0_u8_u4_n104 ) , .A1( u0_u8_u4_n105 ) , .ZN( u0_u8_u4_n146 ) );
  NAND2_X1 u0_u8_u4_U54 (.A2( u0_u8_u4_n101 ) , .A1( u0_u8_u4_n102 ) , .ZN( u0_u8_u4_n160 ) );
  NAND2_X1 u0_u8_u4_U55 (.ZN( u0_u8_u4_n134 ) , .A1( u0_u8_u4_n98 ) , .A2( u0_u8_u4_n99 ) );
  NAND2_X1 u0_u8_u4_U56 (.A1( u0_u8_u4_n103 ) , .A2( u0_u8_u4_n104 ) , .ZN( u0_u8_u4_n143 ) );
  NAND2_X1 u0_u8_u4_U57 (.A2( u0_u8_u4_n105 ) , .ZN( u0_u8_u4_n145 ) , .A1( u0_u8_u4_n98 ) );
  NAND2_X1 u0_u8_u4_U58 (.A1( u0_u8_u4_n100 ) , .A2( u0_u8_u4_n105 ) , .ZN( u0_u8_u4_n120 ) );
  NAND2_X1 u0_u8_u4_U59 (.A1( u0_u8_u4_n102 ) , .A2( u0_u8_u4_n104 ) , .ZN( u0_u8_u4_n148 ) );
  AOI21_X1 u0_u8_u4_U6 (.ZN( u0_u8_u4_n106 ) , .B2( u0_u8_u4_n146 ) , .B1( u0_u8_u4_n158 ) , .A( u0_u8_u4_n170 ) );
  NAND2_X1 u0_u8_u4_U60 (.A2( u0_u8_u4_n100 ) , .A1( u0_u8_u4_n103 ) , .ZN( u0_u8_u4_n157 ) );
  INV_X1 u0_u8_u4_U61 (.A( u0_u8_u4_n150 ) , .ZN( u0_u8_u4_n173 ) );
  INV_X1 u0_u8_u4_U62 (.A( u0_u8_u4_n152 ) , .ZN( u0_u8_u4_n171 ) );
  NAND2_X1 u0_u8_u4_U63 (.A1( u0_u8_u4_n100 ) , .ZN( u0_u8_u4_n118 ) , .A2( u0_u8_u4_n99 ) );
  NAND2_X1 u0_u8_u4_U64 (.A2( u0_u8_u4_n100 ) , .A1( u0_u8_u4_n102 ) , .ZN( u0_u8_u4_n144 ) );
  NAND2_X1 u0_u8_u4_U65 (.A2( u0_u8_u4_n101 ) , .A1( u0_u8_u4_n105 ) , .ZN( u0_u8_u4_n96 ) );
  INV_X1 u0_u8_u4_U66 (.A( u0_u8_u4_n128 ) , .ZN( u0_u8_u4_n174 ) );
  NAND2_X1 u0_u8_u4_U67 (.A2( u0_u8_u4_n102 ) , .ZN( u0_u8_u4_n119 ) , .A1( u0_u8_u4_n98 ) );
  NAND2_X1 u0_u8_u4_U68 (.A2( u0_u8_u4_n101 ) , .A1( u0_u8_u4_n103 ) , .ZN( u0_u8_u4_n147 ) );
  NAND2_X1 u0_u8_u4_U69 (.A2( u0_u8_u4_n104 ) , .ZN( u0_u8_u4_n113 ) , .A1( u0_u8_u4_n99 ) );
  AOI21_X1 u0_u8_u4_U7 (.ZN( u0_u8_u4_n108 ) , .B2( u0_u8_u4_n134 ) , .B1( u0_u8_u4_n155 ) , .A( u0_u8_u4_n156 ) );
  NOR2_X1 u0_u8_u4_U70 (.A2( u0_u8_X_28 ) , .ZN( u0_u8_u4_n150 ) , .A1( u0_u8_u4_n168 ) );
  NOR2_X1 u0_u8_u4_U71 (.A2( u0_u8_X_29 ) , .ZN( u0_u8_u4_n152 ) , .A1( u0_u8_u4_n169 ) );
  NOR2_X1 u0_u8_u4_U72 (.A2( u0_u8_X_30 ) , .ZN( u0_u8_u4_n105 ) , .A1( u0_u8_u4_n176 ) );
  NOR2_X1 u0_u8_u4_U73 (.A2( u0_u8_X_26 ) , .ZN( u0_u8_u4_n100 ) , .A1( u0_u8_u4_n177 ) );
  NOR2_X1 u0_u8_u4_U74 (.A2( u0_u8_X_28 ) , .A1( u0_u8_X_29 ) , .ZN( u0_u8_u4_n128 ) );
  NOR2_X1 u0_u8_u4_U75 (.A2( u0_u8_X_27 ) , .A1( u0_u8_X_30 ) , .ZN( u0_u8_u4_n102 ) );
  NOR2_X1 u0_u8_u4_U76 (.A2( u0_u8_X_25 ) , .A1( u0_u8_X_26 ) , .ZN( u0_u8_u4_n98 ) );
  AND2_X1 u0_u8_u4_U77 (.A2( u0_u8_X_25 ) , .A1( u0_u8_X_26 ) , .ZN( u0_u8_u4_n104 ) );
  AND2_X1 u0_u8_u4_U78 (.A1( u0_u8_X_30 ) , .A2( u0_u8_u4_n176 ) , .ZN( u0_u8_u4_n99 ) );
  AND2_X1 u0_u8_u4_U79 (.A1( u0_u8_X_26 ) , .ZN( u0_u8_u4_n101 ) , .A2( u0_u8_u4_n177 ) );
  AOI21_X1 u0_u8_u4_U8 (.ZN( u0_u8_u4_n109 ) , .A( u0_u8_u4_n153 ) , .B1( u0_u8_u4_n159 ) , .B2( u0_u8_u4_n184 ) );
  AND2_X1 u0_u8_u4_U80 (.A1( u0_u8_X_27 ) , .A2( u0_u8_X_30 ) , .ZN( u0_u8_u4_n103 ) );
  INV_X1 u0_u8_u4_U81 (.A( u0_u8_X_28 ) , .ZN( u0_u8_u4_n169 ) );
  INV_X1 u0_u8_u4_U82 (.A( u0_u8_X_29 ) , .ZN( u0_u8_u4_n168 ) );
  INV_X1 u0_u8_u4_U83 (.A( u0_u8_X_25 ) , .ZN( u0_u8_u4_n177 ) );
  INV_X1 u0_u8_u4_U84 (.A( u0_u8_X_27 ) , .ZN( u0_u8_u4_n176 ) );
  NAND4_X1 u0_u8_u4_U85 (.ZN( u0_out8_25 ) , .A4( u0_u8_u4_n139 ) , .A3( u0_u8_u4_n140 ) , .A2( u0_u8_u4_n141 ) , .A1( u0_u8_u4_n142 ) );
  OAI21_X1 u0_u8_u4_U86 (.B2( u0_u8_u4_n131 ) , .ZN( u0_u8_u4_n141 ) , .A( u0_u8_u4_n175 ) , .B1( u0_u8_u4_n183 ) );
  OAI21_X1 u0_u8_u4_U87 (.A( u0_u8_u4_n128 ) , .B2( u0_u8_u4_n129 ) , .B1( u0_u8_u4_n130 ) , .ZN( u0_u8_u4_n142 ) );
  NAND4_X1 u0_u8_u4_U88 (.ZN( u0_out8_14 ) , .A4( u0_u8_u4_n124 ) , .A3( u0_u8_u4_n125 ) , .A2( u0_u8_u4_n126 ) , .A1( u0_u8_u4_n127 ) );
  AOI22_X1 u0_u8_u4_U89 (.B2( u0_u8_u4_n117 ) , .ZN( u0_u8_u4_n126 ) , .A1( u0_u8_u4_n129 ) , .B1( u0_u8_u4_n152 ) , .A2( u0_u8_u4_n175 ) );
  AOI211_X1 u0_u8_u4_U9 (.B( u0_u8_u4_n136 ) , .A( u0_u8_u4_n137 ) , .C2( u0_u8_u4_n138 ) , .ZN( u0_u8_u4_n139 ) , .C1( u0_u8_u4_n182 ) );
  AOI22_X1 u0_u8_u4_U90 (.ZN( u0_u8_u4_n125 ) , .B2( u0_u8_u4_n131 ) , .A2( u0_u8_u4_n132 ) , .B1( u0_u8_u4_n138 ) , .A1( u0_u8_u4_n178 ) );
  NAND4_X1 u0_u8_u4_U91 (.ZN( u0_out8_8 ) , .A4( u0_u8_u4_n110 ) , .A3( u0_u8_u4_n111 ) , .A2( u0_u8_u4_n112 ) , .A1( u0_u8_u4_n186 ) );
  NAND2_X1 u0_u8_u4_U92 (.ZN( u0_u8_u4_n112 ) , .A2( u0_u8_u4_n130 ) , .A1( u0_u8_u4_n150 ) );
  AOI22_X1 u0_u8_u4_U93 (.ZN( u0_u8_u4_n111 ) , .B2( u0_u8_u4_n132 ) , .A1( u0_u8_u4_n152 ) , .B1( u0_u8_u4_n178 ) , .A2( u0_u8_u4_n97 ) );
  AOI22_X1 u0_u8_u4_U94 (.B2( u0_u8_u4_n149 ) , .B1( u0_u8_u4_n150 ) , .A2( u0_u8_u4_n151 ) , .A1( u0_u8_u4_n152 ) , .ZN( u0_u8_u4_n167 ) );
  NOR4_X1 u0_u8_u4_U95 (.A4( u0_u8_u4_n162 ) , .A3( u0_u8_u4_n163 ) , .A2( u0_u8_u4_n164 ) , .A1( u0_u8_u4_n165 ) , .ZN( u0_u8_u4_n166 ) );
  NAND3_X1 u0_u8_u4_U96 (.ZN( u0_out8_3 ) , .A3( u0_u8_u4_n166 ) , .A1( u0_u8_u4_n167 ) , .A2( u0_u8_u4_n186 ) );
  NAND3_X1 u0_u8_u4_U97 (.A3( u0_u8_u4_n146 ) , .A2( u0_u8_u4_n147 ) , .A1( u0_u8_u4_n148 ) , .ZN( u0_u8_u4_n149 ) );
  NAND3_X1 u0_u8_u4_U98 (.A3( u0_u8_u4_n143 ) , .A2( u0_u8_u4_n144 ) , .A1( u0_u8_u4_n145 ) , .ZN( u0_u8_u4_n151 ) );
  NAND3_X1 u0_u8_u4_U99 (.A3( u0_u8_u4_n121 ) , .ZN( u0_u8_u4_n122 ) , .A2( u0_u8_u4_n144 ) , .A1( u0_u8_u4_n154 ) );
  AND3_X1 u0_u8_u7_U10 (.A3( u0_u8_u7_n110 ) , .A2( u0_u8_u7_n127 ) , .A1( u0_u8_u7_n132 ) , .ZN( u0_u8_u7_n92 ) );
  OAI21_X1 u0_u8_u7_U11 (.A( u0_u8_u7_n161 ) , .B1( u0_u8_u7_n168 ) , .B2( u0_u8_u7_n173 ) , .ZN( u0_u8_u7_n91 ) );
  AOI211_X1 u0_u8_u7_U12 (.A( u0_u8_u7_n117 ) , .ZN( u0_u8_u7_n118 ) , .C2( u0_u8_u7_n126 ) , .C1( u0_u8_u7_n177 ) , .B( u0_u8_u7_n180 ) );
  OAI22_X1 u0_u8_u7_U13 (.B1( u0_u8_u7_n115 ) , .ZN( u0_u8_u7_n117 ) , .A2( u0_u8_u7_n133 ) , .A1( u0_u8_u7_n137 ) , .B2( u0_u8_u7_n162 ) );
  INV_X1 u0_u8_u7_U14 (.A( u0_u8_u7_n116 ) , .ZN( u0_u8_u7_n180 ) );
  NOR3_X1 u0_u8_u7_U15 (.ZN( u0_u8_u7_n115 ) , .A3( u0_u8_u7_n145 ) , .A2( u0_u8_u7_n168 ) , .A1( u0_u8_u7_n169 ) );
  OAI211_X1 u0_u8_u7_U16 (.B( u0_u8_u7_n122 ) , .A( u0_u8_u7_n123 ) , .C2( u0_u8_u7_n124 ) , .ZN( u0_u8_u7_n154 ) , .C1( u0_u8_u7_n162 ) );
  AOI222_X1 u0_u8_u7_U17 (.ZN( u0_u8_u7_n122 ) , .C2( u0_u8_u7_n126 ) , .C1( u0_u8_u7_n145 ) , .B1( u0_u8_u7_n161 ) , .A2( u0_u8_u7_n165 ) , .B2( u0_u8_u7_n170 ) , .A1( u0_u8_u7_n176 ) );
  INV_X1 u0_u8_u7_U18 (.A( u0_u8_u7_n133 ) , .ZN( u0_u8_u7_n176 ) );
  NOR3_X1 u0_u8_u7_U19 (.A2( u0_u8_u7_n134 ) , .A1( u0_u8_u7_n135 ) , .ZN( u0_u8_u7_n136 ) , .A3( u0_u8_u7_n171 ) );
  NOR2_X1 u0_u8_u7_U20 (.A1( u0_u8_u7_n130 ) , .A2( u0_u8_u7_n134 ) , .ZN( u0_u8_u7_n153 ) );
  INV_X1 u0_u8_u7_U21 (.A( u0_u8_u7_n101 ) , .ZN( u0_u8_u7_n165 ) );
  NOR2_X1 u0_u8_u7_U22 (.ZN( u0_u8_u7_n111 ) , .A2( u0_u8_u7_n134 ) , .A1( u0_u8_u7_n169 ) );
  AOI21_X1 u0_u8_u7_U23 (.ZN( u0_u8_u7_n104 ) , .B2( u0_u8_u7_n112 ) , .B1( u0_u8_u7_n127 ) , .A( u0_u8_u7_n164 ) );
  AOI21_X1 u0_u8_u7_U24 (.ZN( u0_u8_u7_n106 ) , .B1( u0_u8_u7_n133 ) , .B2( u0_u8_u7_n146 ) , .A( u0_u8_u7_n162 ) );
  AOI21_X1 u0_u8_u7_U25 (.A( u0_u8_u7_n101 ) , .ZN( u0_u8_u7_n107 ) , .B2( u0_u8_u7_n128 ) , .B1( u0_u8_u7_n175 ) );
  INV_X1 u0_u8_u7_U26 (.A( u0_u8_u7_n138 ) , .ZN( u0_u8_u7_n171 ) );
  INV_X1 u0_u8_u7_U27 (.A( u0_u8_u7_n131 ) , .ZN( u0_u8_u7_n177 ) );
  INV_X1 u0_u8_u7_U28 (.A( u0_u8_u7_n110 ) , .ZN( u0_u8_u7_n174 ) );
  NAND2_X1 u0_u8_u7_U29 (.A1( u0_u8_u7_n129 ) , .A2( u0_u8_u7_n132 ) , .ZN( u0_u8_u7_n149 ) );
  OAI21_X1 u0_u8_u7_U3 (.ZN( u0_u8_u7_n159 ) , .A( u0_u8_u7_n165 ) , .B2( u0_u8_u7_n171 ) , .B1( u0_u8_u7_n174 ) );
  NAND2_X1 u0_u8_u7_U30 (.A1( u0_u8_u7_n113 ) , .A2( u0_u8_u7_n124 ) , .ZN( u0_u8_u7_n130 ) );
  INV_X1 u0_u8_u7_U31 (.A( u0_u8_u7_n112 ) , .ZN( u0_u8_u7_n173 ) );
  INV_X1 u0_u8_u7_U32 (.A( u0_u8_u7_n128 ) , .ZN( u0_u8_u7_n168 ) );
  INV_X1 u0_u8_u7_U33 (.A( u0_u8_u7_n148 ) , .ZN( u0_u8_u7_n169 ) );
  INV_X1 u0_u8_u7_U34 (.A( u0_u8_u7_n127 ) , .ZN( u0_u8_u7_n179 ) );
  NOR2_X1 u0_u8_u7_U35 (.ZN( u0_u8_u7_n101 ) , .A2( u0_u8_u7_n150 ) , .A1( u0_u8_u7_n156 ) );
  AOI211_X1 u0_u8_u7_U36 (.B( u0_u8_u7_n154 ) , .A( u0_u8_u7_n155 ) , .C1( u0_u8_u7_n156 ) , .ZN( u0_u8_u7_n157 ) , .C2( u0_u8_u7_n172 ) );
  INV_X1 u0_u8_u7_U37 (.A( u0_u8_u7_n153 ) , .ZN( u0_u8_u7_n172 ) );
  AOI211_X1 u0_u8_u7_U38 (.B( u0_u8_u7_n139 ) , .A( u0_u8_u7_n140 ) , .C2( u0_u8_u7_n141 ) , .ZN( u0_u8_u7_n142 ) , .C1( u0_u8_u7_n156 ) );
  NAND4_X1 u0_u8_u7_U39 (.A3( u0_u8_u7_n127 ) , .A2( u0_u8_u7_n128 ) , .A1( u0_u8_u7_n129 ) , .ZN( u0_u8_u7_n141 ) , .A4( u0_u8_u7_n147 ) );
  INV_X1 u0_u8_u7_U4 (.A( u0_u8_u7_n111 ) , .ZN( u0_u8_u7_n170 ) );
  AOI21_X1 u0_u8_u7_U40 (.A( u0_u8_u7_n137 ) , .B1( u0_u8_u7_n138 ) , .ZN( u0_u8_u7_n139 ) , .B2( u0_u8_u7_n146 ) );
  OAI22_X1 u0_u8_u7_U41 (.B1( u0_u8_u7_n136 ) , .ZN( u0_u8_u7_n140 ) , .A1( u0_u8_u7_n153 ) , .B2( u0_u8_u7_n162 ) , .A2( u0_u8_u7_n164 ) );
  AOI21_X1 u0_u8_u7_U42 (.ZN( u0_u8_u7_n123 ) , .B1( u0_u8_u7_n165 ) , .B2( u0_u8_u7_n177 ) , .A( u0_u8_u7_n97 ) );
  AOI21_X1 u0_u8_u7_U43 (.B2( u0_u8_u7_n113 ) , .B1( u0_u8_u7_n124 ) , .A( u0_u8_u7_n125 ) , .ZN( u0_u8_u7_n97 ) );
  INV_X1 u0_u8_u7_U44 (.A( u0_u8_u7_n125 ) , .ZN( u0_u8_u7_n161 ) );
  INV_X1 u0_u8_u7_U45 (.A( u0_u8_u7_n152 ) , .ZN( u0_u8_u7_n162 ) );
  AOI22_X1 u0_u8_u7_U46 (.A2( u0_u8_u7_n114 ) , .ZN( u0_u8_u7_n119 ) , .B1( u0_u8_u7_n130 ) , .A1( u0_u8_u7_n156 ) , .B2( u0_u8_u7_n165 ) );
  NAND2_X1 u0_u8_u7_U47 (.A2( u0_u8_u7_n112 ) , .ZN( u0_u8_u7_n114 ) , .A1( u0_u8_u7_n175 ) );
  AND2_X1 u0_u8_u7_U48 (.ZN( u0_u8_u7_n145 ) , .A2( u0_u8_u7_n98 ) , .A1( u0_u8_u7_n99 ) );
  NOR2_X1 u0_u8_u7_U49 (.ZN( u0_u8_u7_n137 ) , .A1( u0_u8_u7_n150 ) , .A2( u0_u8_u7_n161 ) );
  INV_X1 u0_u8_u7_U5 (.A( u0_u8_u7_n149 ) , .ZN( u0_u8_u7_n175 ) );
  AOI21_X1 u0_u8_u7_U50 (.ZN( u0_u8_u7_n105 ) , .B2( u0_u8_u7_n110 ) , .A( u0_u8_u7_n125 ) , .B1( u0_u8_u7_n147 ) );
  NAND2_X1 u0_u8_u7_U51 (.ZN( u0_u8_u7_n146 ) , .A1( u0_u8_u7_n95 ) , .A2( u0_u8_u7_n98 ) );
  NAND2_X1 u0_u8_u7_U52 (.A2( u0_u8_u7_n103 ) , .ZN( u0_u8_u7_n147 ) , .A1( u0_u8_u7_n93 ) );
  NAND2_X1 u0_u8_u7_U53 (.A1( u0_u8_u7_n103 ) , .ZN( u0_u8_u7_n127 ) , .A2( u0_u8_u7_n99 ) );
  OR2_X1 u0_u8_u7_U54 (.ZN( u0_u8_u7_n126 ) , .A2( u0_u8_u7_n152 ) , .A1( u0_u8_u7_n156 ) );
  NAND2_X1 u0_u8_u7_U55 (.A2( u0_u8_u7_n102 ) , .A1( u0_u8_u7_n103 ) , .ZN( u0_u8_u7_n133 ) );
  NAND2_X1 u0_u8_u7_U56 (.ZN( u0_u8_u7_n112 ) , .A2( u0_u8_u7_n96 ) , .A1( u0_u8_u7_n99 ) );
  NAND2_X1 u0_u8_u7_U57 (.A2( u0_u8_u7_n102 ) , .ZN( u0_u8_u7_n128 ) , .A1( u0_u8_u7_n98 ) );
  NAND2_X1 u0_u8_u7_U58 (.A1( u0_u8_u7_n100 ) , .ZN( u0_u8_u7_n113 ) , .A2( u0_u8_u7_n93 ) );
  NAND2_X1 u0_u8_u7_U59 (.A2( u0_u8_u7_n102 ) , .ZN( u0_u8_u7_n124 ) , .A1( u0_u8_u7_n96 ) );
  INV_X1 u0_u8_u7_U6 (.A( u0_u8_u7_n154 ) , .ZN( u0_u8_u7_n178 ) );
  NAND2_X1 u0_u8_u7_U60 (.ZN( u0_u8_u7_n110 ) , .A1( u0_u8_u7_n95 ) , .A2( u0_u8_u7_n96 ) );
  INV_X1 u0_u8_u7_U61 (.A( u0_u8_u7_n150 ) , .ZN( u0_u8_u7_n164 ) );
  AND2_X1 u0_u8_u7_U62 (.ZN( u0_u8_u7_n134 ) , .A1( u0_u8_u7_n93 ) , .A2( u0_u8_u7_n98 ) );
  NAND2_X1 u0_u8_u7_U63 (.A1( u0_u8_u7_n100 ) , .A2( u0_u8_u7_n102 ) , .ZN( u0_u8_u7_n129 ) );
  NAND2_X1 u0_u8_u7_U64 (.A2( u0_u8_u7_n103 ) , .ZN( u0_u8_u7_n131 ) , .A1( u0_u8_u7_n95 ) );
  NAND2_X1 u0_u8_u7_U65 (.A1( u0_u8_u7_n100 ) , .ZN( u0_u8_u7_n138 ) , .A2( u0_u8_u7_n99 ) );
  NAND2_X1 u0_u8_u7_U66 (.ZN( u0_u8_u7_n132 ) , .A1( u0_u8_u7_n93 ) , .A2( u0_u8_u7_n96 ) );
  NAND2_X1 u0_u8_u7_U67 (.A1( u0_u8_u7_n100 ) , .ZN( u0_u8_u7_n148 ) , .A2( u0_u8_u7_n95 ) );
  NOR2_X1 u0_u8_u7_U68 (.A2( u0_u8_X_47 ) , .ZN( u0_u8_u7_n150 ) , .A1( u0_u8_u7_n163 ) );
  NOR2_X1 u0_u8_u7_U69 (.A2( u0_u8_X_43 ) , .A1( u0_u8_X_44 ) , .ZN( u0_u8_u7_n103 ) );
  AOI211_X1 u0_u8_u7_U7 (.ZN( u0_u8_u7_n116 ) , .A( u0_u8_u7_n155 ) , .C1( u0_u8_u7_n161 ) , .C2( u0_u8_u7_n171 ) , .B( u0_u8_u7_n94 ) );
  NOR2_X1 u0_u8_u7_U70 (.A2( u0_u8_X_48 ) , .A1( u0_u8_u7_n166 ) , .ZN( u0_u8_u7_n95 ) );
  NOR2_X1 u0_u8_u7_U71 (.A2( u0_u8_X_45 ) , .A1( u0_u8_X_48 ) , .ZN( u0_u8_u7_n99 ) );
  NOR2_X1 u0_u8_u7_U72 (.A2( u0_u8_X_44 ) , .A1( u0_u8_u7_n167 ) , .ZN( u0_u8_u7_n98 ) );
  NOR2_X1 u0_u8_u7_U73 (.A2( u0_u8_X_46 ) , .A1( u0_u8_X_47 ) , .ZN( u0_u8_u7_n152 ) );
  AND2_X1 u0_u8_u7_U74 (.A1( u0_u8_X_47 ) , .ZN( u0_u8_u7_n156 ) , .A2( u0_u8_u7_n163 ) );
  NAND2_X1 u0_u8_u7_U75 (.A2( u0_u8_X_46 ) , .A1( u0_u8_X_47 ) , .ZN( u0_u8_u7_n125 ) );
  AND2_X1 u0_u8_u7_U76 (.A2( u0_u8_X_45 ) , .A1( u0_u8_X_48 ) , .ZN( u0_u8_u7_n102 ) );
  AND2_X1 u0_u8_u7_U77 (.A2( u0_u8_X_43 ) , .A1( u0_u8_X_44 ) , .ZN( u0_u8_u7_n96 ) );
  AND2_X1 u0_u8_u7_U78 (.A1( u0_u8_X_44 ) , .ZN( u0_u8_u7_n100 ) , .A2( u0_u8_u7_n167 ) );
  AND2_X1 u0_u8_u7_U79 (.A1( u0_u8_X_48 ) , .A2( u0_u8_u7_n166 ) , .ZN( u0_u8_u7_n93 ) );
  OAI222_X1 u0_u8_u7_U8 (.C2( u0_u8_u7_n101 ) , .B2( u0_u8_u7_n111 ) , .A1( u0_u8_u7_n113 ) , .C1( u0_u8_u7_n146 ) , .A2( u0_u8_u7_n162 ) , .B1( u0_u8_u7_n164 ) , .ZN( u0_u8_u7_n94 ) );
  INV_X1 u0_u8_u7_U80 (.A( u0_u8_X_46 ) , .ZN( u0_u8_u7_n163 ) );
  INV_X1 u0_u8_u7_U81 (.A( u0_u8_X_43 ) , .ZN( u0_u8_u7_n167 ) );
  INV_X1 u0_u8_u7_U82 (.A( u0_u8_X_45 ) , .ZN( u0_u8_u7_n166 ) );
  NAND4_X1 u0_u8_u7_U83 (.ZN( u0_out8_27 ) , .A4( u0_u8_u7_n118 ) , .A3( u0_u8_u7_n119 ) , .A2( u0_u8_u7_n120 ) , .A1( u0_u8_u7_n121 ) );
  OAI21_X1 u0_u8_u7_U84 (.ZN( u0_u8_u7_n121 ) , .B2( u0_u8_u7_n145 ) , .A( u0_u8_u7_n150 ) , .B1( u0_u8_u7_n174 ) );
  OAI21_X1 u0_u8_u7_U85 (.ZN( u0_u8_u7_n120 ) , .A( u0_u8_u7_n161 ) , .B2( u0_u8_u7_n170 ) , .B1( u0_u8_u7_n179 ) );
  NAND4_X1 u0_u8_u7_U86 (.ZN( u0_out8_15 ) , .A4( u0_u8_u7_n142 ) , .A3( u0_u8_u7_n143 ) , .A2( u0_u8_u7_n144 ) , .A1( u0_u8_u7_n178 ) );
  OR2_X1 u0_u8_u7_U87 (.A2( u0_u8_u7_n125 ) , .A1( u0_u8_u7_n129 ) , .ZN( u0_u8_u7_n144 ) );
  AOI22_X1 u0_u8_u7_U88 (.A2( u0_u8_u7_n126 ) , .ZN( u0_u8_u7_n143 ) , .B2( u0_u8_u7_n165 ) , .B1( u0_u8_u7_n173 ) , .A1( u0_u8_u7_n174 ) );
  NAND4_X1 u0_u8_u7_U89 (.ZN( u0_out8_5 ) , .A4( u0_u8_u7_n108 ) , .A3( u0_u8_u7_n109 ) , .A1( u0_u8_u7_n116 ) , .A2( u0_u8_u7_n123 ) );
  OAI221_X1 u0_u8_u7_U9 (.C1( u0_u8_u7_n101 ) , .C2( u0_u8_u7_n147 ) , .ZN( u0_u8_u7_n155 ) , .B2( u0_u8_u7_n162 ) , .A( u0_u8_u7_n91 ) , .B1( u0_u8_u7_n92 ) );
  AOI22_X1 u0_u8_u7_U90 (.ZN( u0_u8_u7_n109 ) , .A2( u0_u8_u7_n126 ) , .B2( u0_u8_u7_n145 ) , .B1( u0_u8_u7_n156 ) , .A1( u0_u8_u7_n171 ) );
  NOR4_X1 u0_u8_u7_U91 (.A4( u0_u8_u7_n104 ) , .A3( u0_u8_u7_n105 ) , .A2( u0_u8_u7_n106 ) , .A1( u0_u8_u7_n107 ) , .ZN( u0_u8_u7_n108 ) );
  NAND4_X1 u0_u8_u7_U92 (.ZN( u0_out8_21 ) , .A4( u0_u8_u7_n157 ) , .A3( u0_u8_u7_n158 ) , .A2( u0_u8_u7_n159 ) , .A1( u0_u8_u7_n160 ) );
  OAI21_X1 u0_u8_u7_U93 (.B1( u0_u8_u7_n145 ) , .ZN( u0_u8_u7_n160 ) , .A( u0_u8_u7_n161 ) , .B2( u0_u8_u7_n177 ) );
  AOI22_X1 u0_u8_u7_U94 (.B2( u0_u8_u7_n149 ) , .B1( u0_u8_u7_n150 ) , .A2( u0_u8_u7_n151 ) , .A1( u0_u8_u7_n152 ) , .ZN( u0_u8_u7_n158 ) );
  NAND3_X1 u0_u8_u7_U95 (.A3( u0_u8_u7_n146 ) , .A2( u0_u8_u7_n147 ) , .A1( u0_u8_u7_n148 ) , .ZN( u0_u8_u7_n151 ) );
  NAND3_X1 u0_u8_u7_U96 (.A3( u0_u8_u7_n131 ) , .A2( u0_u8_u7_n132 ) , .A1( u0_u8_u7_n133 ) , .ZN( u0_u8_u7_n135 ) );
  OAI21_X1 u0_uk_U1022 (.ZN( u0_K9_44 ) , .B1( u0_uk_n147 ) , .B2( u0_uk_n273 ) , .A( u0_uk_n721 ) );
  NAND2_X1 u0_uk_U1023 (.A1( u0_uk_K_r7_0 ) , .A2( u0_uk_n217 ) , .ZN( u0_uk_n721 ) );
  OAI21_X1 u0_uk_U1030 (.ZN( u0_K16_41 ) , .B1( u0_uk_n142 ) , .B2( u0_uk_n643 ) , .A( u0_uk_n898 ) );
  NAND2_X1 u0_uk_U1035 (.A1( u0_uk_K_r4_31 ) , .ZN( u0_uk_n790 ) , .A2( u0_uk_n92 ) );
  OAI21_X1 u0_uk_U1036 (.ZN( u0_K16_28 ) , .B1( u0_uk_n60 ) , .B2( u0_uk_n669 ) , .A( u0_uk_n905 ) );
  NAND2_X1 u0_uk_U1037 (.A1( u0_uk_K_r14_8 ) , .A2( u0_uk_n83 ) , .ZN( u0_uk_n905 ) );
  OAI21_X1 u0_uk_U1040 (.ZN( u0_K7_31 ) , .B1( u0_uk_n128 ) , .B2( u0_uk_n380 ) , .A( u0_uk_n772 ) );
  NAND2_X1 u0_uk_U1041 (.A1( u0_uk_K_r5_16 ) , .A2( u0_uk_n102 ) , .ZN( u0_uk_n772 ) );
  OAI21_X1 u0_uk_U1052 (.ZN( u0_K16_42 ) , .B2( u0_uk_n647 ) , .A( u0_uk_n897 ) , .B1( u0_uk_n92 ) );
  OAI21_X1 u0_uk_U1056 (.ZN( u0_K7_38 ) , .B1( u0_uk_n128 ) , .B2( u0_uk_n389 ) , .A( u0_uk_n767 ) );
  NAND2_X1 u0_uk_U1057 (.A1( u0_uk_K_r5_8 ) , .A2( u0_uk_n117 ) , .ZN( u0_uk_n767 ) );
  INV_X1 u0_uk_U1064 (.A( u0_key_r_6 ) , .ZN( u0_uk_n712 ) );
  INV_X1 u0_uk_U1065 (.A( u0_key_r_54 ) , .ZN( u0_uk_n673 ) );
  INV_X1 u0_uk_U1068 (.A( u0_key_r_26 ) , .ZN( u0_uk_n697 ) );
  OAI22_X1 u0_uk_U107 (.ZN( u0_K1_5 ) , .A1( u0_uk_n188 ) , .B2( u0_uk_n708 ) , .A2( u0_uk_n712 ) , .B1( u0_uk_n99 ) );
  INV_X1 u0_uk_U1070 (.A( u0_key_r_34 ) , .ZN( u0_uk_n690 ) );
  INV_X1 u0_uk_U1071 (.A( u0_key_r_27 ) , .ZN( u0_uk_n696 ) );
  INV_X1 u0_uk_U1072 (.A( u0_key_r_24 ) , .ZN( u0_uk_n699 ) );
  INV_X1 u0_uk_U1073 (.A( u0_key_r_20 ) , .ZN( u0_uk_n703 ) );
  INV_X1 u0_uk_U1078 (.A( u0_key_r_13 ) , .ZN( u0_uk_n708 ) );
  INV_X1 u0_uk_U1081 (.A( u0_key_r_19 ) , .ZN( u0_uk_n704 ) );
  INV_X1 u0_uk_U1082 (.A( u0_key_r_4 ) , .ZN( u0_uk_n713 ) );
  INV_X1 u0_uk_U1083 (.A( u0_key_r_17 ) , .ZN( u0_uk_n705 ) );
  INV_X1 u0_uk_U1084 (.A( u0_key_r_53 ) , .ZN( u0_uk_n674 ) );
  OAI21_X1 u0_uk_U1085 (.ZN( u0_K13_28 ) , .B2( u0_uk_n105 ) , .B1( u0_uk_n252 ) , .A( u0_uk_n947 ) );
  NAND2_X1 u0_uk_U1086 (.A1( u0_uk_K_r11_21 ) , .A2( u0_uk_n214 ) , .ZN( u0_uk_n947 ) );
  OAI21_X1 u0_uk_U1093 (.ZN( u0_K16_39 ) , .B1( u0_uk_n250 ) , .B2( u0_uk_n657 ) , .A( u0_uk_n899 ) );
  NAND2_X1 u0_uk_U1094 (.A1( u0_uk_K_r14_15 ) , .A2( u0_uk_n208 ) , .ZN( u0_uk_n899 ) );
  INV_X1 u0_uk_U1099 (.A( u0_key_r_40 ) , .ZN( u0_uk_n684 ) );
  INV_X1 u0_uk_U1100 (.A( u0_key_r_47 ) , .ZN( u0_uk_n679 ) );
  INV_X1 u0_uk_U1103 (.ZN( u0_K1_11 ) , .A( u0_uk_n892 ) );
  AOI22_X1 u0_uk_U1104 (.B2( u0_key_r_32 ) , .A2( u0_key_r_39 ) , .B1( u0_uk_n145 ) , .A1( u0_uk_n240 ) , .ZN( u0_uk_n892 ) );
  INV_X1 u0_uk_U1115 (.ZN( u0_K1_20 ) , .A( u0_uk_n886 ) );
  AOI22_X1 u0_uk_U1116 (.B2( u0_key_r_48 ) , .A2( u0_key_r_55 ) , .B1( u0_uk_n145 ) , .A1( u0_uk_n242 ) , .ZN( u0_uk_n886 ) );
  INV_X1 u0_uk_U1121 (.ZN( u0_K5_20 ) , .A( u0_uk_n816 ) );
  AOI22_X1 u0_uk_U1122 (.B2( u0_uk_K_r3_24 ) , .A2( u0_uk_K_r3_47 ) , .B1( u0_uk_n100 ) , .A1( u0_uk_n257 ) , .ZN( u0_uk_n816 ) );
  INV_X1 u0_uk_U1127 (.ZN( u0_K7_32 ) , .A( u0_uk_n771 ) );
  AOI22_X1 u0_uk_U1128 (.B2( u0_uk_K_r5_0 ) , .A2( u0_uk_K_r5_51 ) , .B1( u0_uk_n146 ) , .A1( u0_uk_n213 ) , .ZN( u0_uk_n771 ) );
  INV_X1 u0_uk_U1139 (.ZN( u0_K7_34 ) , .A( u0_uk_n770 ) );
  OAI22_X1 u0_uk_U1157 (.ZN( u0_K1_1 ) , .A1( u0_uk_n142 ) , .B1( u0_uk_n217 ) , .A2( u0_uk_n679 ) , .B2( u0_uk_n684 ) );
  OAI22_X1 u0_uk_U144 (.ZN( u0_K1_19 ) , .B1( u0_uk_n110 ) , .A1( u0_uk_n187 ) , .A2( u0_uk_n673 ) , .B2( u0_uk_n713 ) );
  INV_X1 u0_uk_U15 (.A( u0_uk_n155 ) , .ZN( u0_uk_n99 ) );
  INV_X1 u0_uk_U153 (.ZN( u0_K9_19 ) , .A( u0_uk_n735 ) );
  INV_X1 u0_uk_U172 (.A( u0_key_r_25 ) , .ZN( u0_uk_n698 ) );
  OAI21_X1 u0_uk_U175 (.ZN( u0_K16_30 ) , .B1( u0_uk_n147 ) , .B2( u0_uk_n632 ) , .A( u0_uk_n902 ) );
  NAND2_X1 u0_uk_U176 (.A1( u0_uk_K_r14_45 ) , .A2( u0_uk_n203 ) , .ZN( u0_uk_n902 ) );
  INV_X1 u0_uk_U18 (.ZN( u0_uk_n117 ) , .A( u0_uk_n182 ) );
  OAI22_X1 u0_uk_U189 (.ZN( u0_K1_24 ) , .A1( u0_uk_n118 ) , .B1( u0_uk_n222 ) , .A2( u0_uk_n703 ) , .B2( u0_uk_n708 ) );
  OAI21_X1 u0_uk_U203 (.ZN( u0_K9_30 ) , .B2( u0_uk_n288 ) , .B1( u0_uk_n60 ) , .A( u0_uk_n728 ) );
  OAI22_X1 u0_uk_U214 (.ZN( u0_K16_31 ) , .B1( u0_uk_n155 ) , .B2( u0_uk_n663 ) , .A2( u0_uk_n666 ) , .A1( u0_uk_n99 ) );
  OAI22_X1 u0_uk_U225 (.ZN( u0_K13_31 ) , .B2( u0_uk_n116 ) , .A1( u0_uk_n209 ) , .B1( u0_uk_n92 ) , .A2( u0_uk_n98 ) );
  INV_X1 u0_uk_U264 (.ZN( u0_K9_48 ) , .A( u0_uk_n719 ) );
  OAI22_X1 u0_uk_U283 (.ZN( u0_K1_8 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n182 ) , .B2( u0_uk_n699 ) , .A2( u0_uk_n712 ) );
  OAI22_X1 u0_uk_U290 (.ZN( u0_K5_8 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n182 ) , .A2( u0_uk_n451 ) , .B2( u0_uk_n473 ) );
  OAI22_X1 u0_uk_U296 (.ZN( u0_K7_26 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n230 ) , .A2( u0_uk_n368 ) , .B2( u0_uk_n388 ) );
  INV_X1 u0_uk_U300 (.ZN( u0_K9_26 ) , .A( u0_uk_n731 ) );
  BUF_X1 u0_uk_U31 (.Z( u0_uk_n155 ) , .A( u0_uk_n223 ) );
  OAI21_X1 u0_uk_U310 (.ZN( u0_K13_26 ) , .B1( u0_uk_n10 ) , .B2( u0_uk_n123 ) , .A( u0_uk_n948 ) );
  OAI21_X1 u0_uk_U323 (.ZN( u0_K9_46 ) , .B1( u0_uk_n11 ) , .B2( u0_uk_n281 ) , .A( u0_uk_n720 ) );
  NAND2_X1 u0_uk_U331 (.A1( u0_key_r_49 ) , .A2( u0_uk_n117 ) , .ZN( u0_uk_n871 ) );
  OAI21_X1 u0_uk_U349 (.ZN( u0_K1_4 ) , .B1( u0_uk_n217 ) , .B2( u0_uk_n674 ) , .A( u0_uk_n869 ) );
  BUF_X1 u0_uk_U35 (.A( u0_uk_n155 ) , .Z( u0_uk_n187 ) );
  NAND2_X1 u0_uk_U350 (.A1( u0_key_r_3 ) , .A2( u0_uk_n251 ) , .ZN( u0_uk_n869 ) );
  OAI22_X1 u0_uk_U351 (.ZN( u0_K16_40 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n155 ) , .A2( u0_uk_n632 ) , .B2( u0_uk_n670 ) );
  OAI22_X1 u0_uk_U364 (.ZN( u0_K7_40 ) , .A1( u0_uk_n223 ) , .B1( u0_uk_n31 ) , .B2( u0_uk_n394 ) , .A2( u0_uk_n406 ) );
  OAI22_X1 u0_uk_U384 (.ZN( u0_K9_28 ) , .B1( u0_uk_n162 ) , .A2( u0_uk_n274 ) , .B2( u0_uk_n281 ) , .A1( u0_uk_n99 ) );
  OAI22_X1 u0_uk_U385 (.ZN( u0_K7_28 ) , .A1( u0_uk_n223 ) , .B1( u0_uk_n31 ) , .A2( u0_uk_n378 ) , .B2( u0_uk_n387 ) );
  OAI22_X1 u0_uk_U391 (.ZN( u0_K1_9 ) , .B1( u0_uk_n231 ) , .A2( u0_uk_n673 ) , .B2( u0_uk_n679 ) , .A1( u0_uk_n94 ) );
  BUF_X1 u0_uk_U40 (.Z( u0_uk_n230 ) , .A( u0_uk_n257 ) );
  OAI22_X1 u0_uk_U443 (.ZN( u0_K16_33 ) , .A1( u0_uk_n187 ) , .B1( u0_uk_n31 ) , .A2( u0_uk_n633 ) , .B2( u0_uk_n638 ) );
  OAI22_X1 u0_uk_U445 (.ZN( u0_K13_33 ) , .A1( u0_uk_n100 ) , .A2( u0_uk_n130 ) , .B2( u0_uk_n135 ) , .B1( u0_uk_n238 ) );
  OAI22_X1 u0_uk_U447 (.ZN( u0_K7_33 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n230 ) , .A2( u0_uk_n374 ) , .B2( u0_uk_n394 ) );
  INV_X1 u0_uk_U452 (.ZN( u0_K16_37 ) , .A( u0_uk_n900 ) );
  AOI22_X1 u0_uk_U453 (.B2( u0_uk_K_r14_2 ) , .A2( u0_uk_K_r14_50 ) , .B1( u0_uk_n141 ) , .A1( u0_uk_n251 ) , .ZN( u0_uk_n900 ) );
  OAI22_X1 u0_uk_U455 (.ZN( u0_K13_37 ) , .A2( u0_uk_n112 ) , .B2( u0_uk_n124 ) , .A1( u0_uk_n209 ) , .B1( u0_uk_n92 ) );
  OAI22_X1 u0_uk_U474 (.ZN( u0_K13_29 ) , .A2( u0_uk_n113 ) , .B2( u0_uk_n116 ) , .A1( u0_uk_n118 ) , .B1( u0_uk_n161 ) );
  OAI22_X1 u0_uk_U484 (.ZN( u0_K9_29 ) , .B1( u0_uk_n161 ) , .A2( u0_uk_n289 ) , .B2( u0_uk_n293 ) , .A1( u0_uk_n99 ) );
  OAI22_X1 u0_uk_U486 (.ZN( u0_K7_29 ) , .A1( u0_uk_n162 ) , .B1( u0_uk_n31 ) , .A2( u0_uk_n368 ) , .B2( u0_uk_n399 ) );
  OAI21_X1 u0_uk_U495 (.ZN( u0_K1_2 ) , .B1( u0_uk_n250 ) , .B2( u0_uk_n713 ) , .A( u0_uk_n881 ) );
  NAND2_X1 u0_uk_U496 (.A1( u0_key_r_11 ) , .A2( u0_uk_n202 ) , .ZN( u0_uk_n881 ) );
  OAI21_X1 u0_uk_U499 (.ZN( u0_K1_12 ) , .B1( u0_uk_n128 ) , .B2( u0_uk_n704 ) , .A( u0_uk_n891 ) );
  NAND2_X1 u0_uk_U500 (.A1( u0_key_r_12 ) , .A2( u0_uk_n10 ) , .ZN( u0_uk_n891 ) );
  OAI21_X1 u0_uk_U524 (.ZN( u0_K5_12 ) , .B1( u0_uk_n202 ) , .B2( u0_uk_n483 ) , .A( u0_uk_n818 ) );
  NAND2_X1 u0_uk_U525 (.A1( u0_uk_K_r3_11 ) , .A2( u0_uk_n208 ) , .ZN( u0_uk_n818 ) );
  OAI22_X1 u0_uk_U539 (.ZN( u0_K5_17 ) , .B1( u0_uk_n203 ) , .A2( u0_uk_n464 ) , .B2( u0_uk_n484 ) , .A1( u0_uk_n99 ) );
  INV_X1 u0_uk_U552 (.ZN( u0_K16_29 ) , .A( u0_uk_n904 ) );
  OAI22_X1 u0_uk_U554 (.ZN( u0_K16_36 ) , .A1( u0_uk_n155 ) , .B1( u0_uk_n63 ) , .A2( u0_uk_n648 ) , .B2( u0_uk_n655 ) );
  INV_X1 u0_uk_U558 (.ZN( u0_K7_36 ) , .A( u0_uk_n768 ) );
  AOI22_X1 u0_uk_U559 (.B2( u0_uk_K_r5_1 ) , .A2( u0_uk_K_r5_21 ) , .B1( u0_uk_n146 ) , .A1( u0_uk_n257 ) , .ZN( u0_uk_n768 ) );
  OAI22_X1 u0_uk_U570 (.ZN( u0_K5_10 ) , .B1( u0_uk_n208 ) , .A2( u0_uk_n465 ) , .B2( u0_uk_n485 ) , .A1( u0_uk_n99 ) );
  INV_X1 u0_uk_U58 (.ZN( u0_K16_34 ) , .A( u0_uk_n901 ) );
  INV_X1 u0_uk_U586 (.ZN( u0_K1_10 ) , .A( u0_uk_n893 ) );
  AOI22_X1 u0_uk_U587 (.B2( u0_key_r_41 ) , .A2( u0_key_r_48 ) , .B1( u0_uk_n142 ) , .A1( u0_uk_n251 ) , .ZN( u0_uk_n893 ) );
  AOI22_X1 u0_uk_U59 (.B2( u0_uk_K_r14_2 ) , .A2( u0_uk_K_r14_9 ) , .A1( u0_uk_n145 ) , .B1( u0_uk_n202 ) , .ZN( u0_uk_n901 ) );
  INV_X1 u0_uk_U596 (.ZN( u0_K9_22 ) , .A( u0_uk_n732 ) );
  INV_X1 u0_uk_U599 (.ZN( u0_K5_22 ) , .A( u0_uk_n815 ) );
  INV_X1 u0_uk_U601 (.ZN( u0_K1_22 ) , .A( u0_uk_n885 ) );
  AOI22_X1 u0_uk_U602 (.B2( u0_key_r_25 ) , .A2( u0_key_r_32 ) , .B1( u0_uk_n145 ) , .A1( u0_uk_n213 ) , .ZN( u0_uk_n885 ) );
  OAI22_X1 u0_uk_U603 (.ZN( u0_K16_35 ) , .B1( u0_uk_n100 ) , .A1( u0_uk_n155 ) , .A2( u0_uk_n643 ) , .B2( u0_uk_n650 ) );
  OAI21_X1 u0_uk_U606 (.ZN( u0_K7_35 ) , .B1( u0_uk_n128 ) , .B2( u0_uk_n406 ) , .A( u0_uk_n769 ) );
  NAND2_X1 u0_uk_U607 (.A1( u0_uk_K_r5_37 ) , .ZN( u0_uk_n769 ) , .A2( u0_uk_n92 ) );
  OAI22_X1 u0_uk_U609 (.ZN( u0_K13_35 ) , .B2( u0_uk_n124 ) , .B1( u0_uk_n214 ) , .A1( u0_uk_n27 ) , .A2( u0_uk_n95 ) );
  OAI22_X1 u0_uk_U640 (.ZN( u0_K5_11 ) , .B1( u0_uk_n208 ) , .B2( u0_uk_n465 ) , .A2( u0_uk_n489 ) , .A1( u0_uk_n99 ) );
  OAI22_X1 u0_uk_U656 (.ZN( u0_K1_7 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n203 ) , .A2( u0_uk_n696 ) , .B2( u0_uk_n703 ) );
  OAI22_X1 u0_uk_U657 (.ZN( u0_K9_25 ) , .B1( u0_uk_n162 ) , .A2( u0_uk_n273 ) , .B2( u0_uk_n280 ) , .A1( u0_uk_n99 ) );
  OAI22_X1 u0_uk_U671 (.ZN( u0_K9_43 ) , .A1( u0_uk_n146 ) , .B1( u0_uk_n155 ) , .A2( u0_uk_n293 ) , .B2( u0_uk_n300 ) );
  OAI22_X1 u0_uk_U689 (.ZN( u0_K13_25 ) , .A1( u0_uk_n118 ) , .B2( u0_uk_n123 ) , .B1( u0_uk_n242 ) , .A2( u0_uk_n98 ) );
  OAI22_X1 u0_uk_U694 (.ZN( u0_K16_25 ) , .B1( u0_uk_n117 ) , .A1( u0_uk_n240 ) , .A2( u0_uk_n642 ) , .B2( u0_uk_n649 ) );
  OAI21_X1 u0_uk_U706 (.ZN( u0_K5_7 ) , .B1( u0_uk_n163 ) , .B2( u0_uk_n453 ) , .A( u0_uk_n802 ) );
  NAND2_X1 u0_uk_U707 (.A1( u0_uk_K_r3_19 ) , .A2( u0_uk_n203 ) , .ZN( u0_uk_n802 ) );
  INV_X1 u0_uk_U708 (.ZN( u0_K7_25 ) , .A( u0_uk_n775 ) );
  OAI22_X1 u0_uk_U717 (.ZN( u0_K16_32 ) , .B1( u0_uk_n118 ) , .A1( u0_uk_n155 ) , .A2( u0_uk_n649 ) , .B2( u0_uk_n657 ) );
  OAI22_X1 u0_uk_U720 (.ZN( u0_K13_32 ) , .B2( u0_uk_n106 ) , .A2( u0_uk_n130 ) , .A1( u0_uk_n191 ) , .B1( u0_uk_n92 ) );
  INV_X1 u0_uk_U736 (.ZN( u0_K7_42 ) , .A( u0_uk_n766 ) );
  OAI22_X1 u0_uk_U750 (.ZN( u0_K16_27 ) , .B1( u0_uk_n109 ) , .A1( u0_uk_n187 ) , .A2( u0_uk_n658 ) , .B2( u0_uk_n663 ) );
  OAI22_X1 u0_uk_U756 (.ZN( u0_K1_21 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n147 ) , .A2( u0_uk_n699 ) , .B2( u0_uk_n705 ) );
  OAI22_X1 u0_uk_U760 (.ZN( u0_K13_27 ) , .A2( u0_uk_n111 ) , .B2( u0_uk_n134 ) , .B1( u0_uk_n238 ) , .A1( u0_uk_n94 ) );
  OAI22_X1 u0_uk_U764 (.ZN( u0_K9_21 ) , .B1( u0_uk_n162 ) , .A2( u0_uk_n285 ) , .B2( u0_uk_n290 ) , .A1( u0_uk_n94 ) );
  OAI22_X1 u0_uk_U765 (.ZN( u0_K5_21 ) , .B1( u0_uk_n163 ) , .A2( u0_uk_n459 ) , .B2( u0_uk_n479 ) , .A1( u0_uk_n99 ) );
  INV_X1 u0_uk_U792 (.ZN( u0_K7_27 ) , .A( u0_uk_n774 ) );
  AOI22_X1 u0_uk_U793 (.B2( u0_uk_K_r5_23 ) , .A2( u0_uk_K_r5_43 ) , .B1( u0_uk_n146 ) , .A1( u0_uk_n223 ) , .ZN( u0_uk_n774 ) );
  INV_X1 u0_uk_U796 (.ZN( u0_K9_27 ) , .A( u0_uk_n730 ) );
  AOI22_X1 u0_uk_U797 (.B2( u0_uk_K_r7_2 ) , .A2( u0_uk_K_r7_9 ) , .A1( u0_uk_n240 ) , .ZN( u0_uk_n730 ) , .B1( u0_uk_n94 ) );
  INV_X1 u0_uk_U831 (.ZN( u0_K9_20 ) , .A( u0_uk_n733 ) );
  AOI22_X1 u0_uk_U832 (.B2( u0_uk_K_r7_32 ) , .A2( u0_uk_K_r7_39 ) , .B1( u0_uk_n10 ) , .A1( u0_uk_n240 ) , .ZN( u0_uk_n733 ) );
  OAI22_X1 u0_uk_U840 (.ZN( u0_K1_6 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n222 ) , .A2( u0_uk_n683 ) , .B2( u0_uk_n690 ) );
  INV_X1 u0_uk_U841 (.A( u0_key_r_41 ) , .ZN( u0_uk_n683 ) );
  OAI22_X1 u0_uk_U876 (.ZN( u0_K13_34 ) , .A2( u0_uk_n104 ) , .B2( u0_uk_n120 ) , .A1( u0_uk_n209 ) , .B1( u0_uk_n92 ) );
  OAI22_X1 u0_uk_U89 (.ZN( u0_K13_41 ) , .A2( u0_uk_n120 ) , .B2( u0_uk_n135 ) , .A1( u0_uk_n209 ) , .B1( u0_uk_n93 ) );
  OAI22_X1 u0_uk_U90 (.ZN( u0_K7_41 ) , .A1( u0_uk_n146 ) , .B1( u0_uk_n250 ) , .B2( u0_uk_n372 ) , .A2( u0_uk_n402 ) );
  OAI22_X1 u0_uk_U904 (.ZN( u0_K9_24 ) , .A1( u0_uk_n257 ) , .B1( u0_uk_n27 ) , .A2( u0_uk_n272 ) , .B2( u0_uk_n314 ) );
  OAI22_X1 u0_uk_U911 (.ZN( u0_K7_30 ) , .A1( u0_uk_n213 ) , .B1( u0_uk_n31 ) , .A2( u0_uk_n367 ) , .B2( u0_uk_n398 ) );
  OAI22_X1 u0_uk_U922 (.ZN( u0_K7_39 ) , .A1( u0_uk_n257 ) , .B1( u0_uk_n31 ) , .A2( u0_uk_n365 ) , .B2( u0_uk_n372 ) );
  OAI22_X1 u0_uk_U930 (.ZN( u0_K9_23 ) , .B1( u0_uk_n162 ) , .A2( u0_uk_n296 ) , .B2( u0_uk_n304 ) , .A1( u0_uk_n99 ) );
  OAI22_X1 u0_uk_U931 (.ZN( u0_K9_47 ) , .A1( u0_uk_n129 ) , .B1( u0_uk_n187 ) , .A2( u0_uk_n275 ) , .B2( u0_uk_n282 ) );
  OAI22_X1 u0_uk_U967 (.ZN( u0_K13_38 ) , .B2( u0_uk_n103 ) , .B1( u0_uk_n147 ) , .A2( u0_uk_n97 ) , .A1( u0_uk_n99 ) );
  OAI22_X1 u0_uk_U969 (.ZN( u0_K7_37 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n230 ) , .A2( u0_uk_n365 ) , .B2( u0_uk_n389 ) );
  OAI22_X1 u0_uk_U993 (.ZN( u0_K1_3 ) , .A1( u0_uk_n142 ) , .B1( u0_uk_n188 ) , .A2( u0_uk_n697 ) , .B2( u0_uk_n704 ) );
  XOR2_X1 u2_U10 (.B( u2_L1_29 ) , .Z( u2_N92 ) , .A( u2_out2_29 ) );
  XOR2_X1 u2_U102 (.B( u2_L12_25 ) , .Z( u2_N440 ) , .A( u2_out13_25 ) );
  XOR2_X1 u2_U115 (.B( u2_L12_14 ) , .Z( u2_N429 ) , .A( u2_out13_14 ) );
  XOR2_X1 u2_U12 (.B( u2_L1_27 ) , .Z( u2_N90 ) , .A( u2_out2_27 ) );
  XOR2_X1 u2_U121 (.B( u2_L12_8 ) , .Z( u2_N423 ) , .A( u2_out13_8 ) );
  XOR2_X1 u2_U127 (.B( u2_L12_3 ) , .Z( u2_N418 ) , .A( u2_out13_3 ) );
  XOR2_X1 u2_U133 (.B( u2_L11_29 ) , .Z( u2_N412 ) , .A( u2_out12_29 ) );
  XOR2_X1 u2_U137 (.B( u2_L11_26 ) , .Z( u2_N409 ) , .A( u2_out12_26 ) );
  XOR2_X1 u2_U138 (.B( u2_L11_25 ) , .Z( u2_N408 ) , .A( u2_out12_25 ) );
  XOR2_X1 u2_U14 (.B( u2_L1_26 ) , .Z( u2_N89 ) , .A( u2_out2_26 ) );
  XOR2_X1 u2_U143 (.B( u2_L11_20 ) , .Z( u2_N403 ) , .A( u2_out12_20 ) );
  XOR2_X1 u2_U144 (.B( u2_L11_19 ) , .Z( u2_N402 ) , .A( u2_out12_19 ) );
  XOR2_X1 u2_U15 (.B( u2_L1_25 ) , .Z( u2_N88 ) , .A( u2_out2_25 ) );
  XOR2_X1 u2_U151 (.B( u2_L11_14 ) , .Z( u2_N397 ) , .A( u2_out12_14 ) );
  XOR2_X1 u2_U154 (.B( u2_L11_11 ) , .Z( u2_N394 ) , .A( u2_out12_11 ) );
  XOR2_X1 u2_U155 (.B( u2_L11_10 ) , .Z( u2_N393 ) , .A( u2_out12_10 ) );
  XOR2_X1 u2_U157 (.B( u2_L11_8 ) , .Z( u2_N391 ) , .A( u2_out12_8 ) );
  XOR2_X1 u2_U162 (.B( u2_L11_4 ) , .Z( u2_N387 ) , .A( u2_out12_4 ) );
  XOR2_X1 u2_U163 (.B( u2_L11_3 ) , .Z( u2_N386 ) , .A( u2_out12_3 ) );
  XOR2_X1 u2_U165 (.B( u2_L11_1 ) , .Z( u2_N384 ) , .A( u2_out12_1 ) );
  XOR2_X1 u2_U18 (.B( u2_L1_22 ) , .Z( u2_N85 ) , .A( u2_out2_22 ) );
  XOR2_X1 u2_U19 (.B( u2_L1_21 ) , .Z( u2_N84 ) , .A( u2_out2_21 ) );
  XOR2_X1 u2_U20 (.B( u2_L1_20 ) , .Z( u2_N83 ) , .A( u2_out2_20 ) );
  XOR2_X1 u2_U202 (.B( u2_L9_31 ) , .Z( u2_N350 ) , .A( u2_out10_31 ) );
  XOR2_X1 u2_U204 (.B( u2_L9_30 ) , .Z( u2_N349 ) , .A( u2_out10_30 ) );
  XOR2_X1 u2_U206 (.B( u2_L9_28 ) , .Z( u2_N347 ) , .A( u2_out10_28 ) );
  XOR2_X1 u2_U208 (.B( u2_L9_26 ) , .Z( u2_N345 ) , .A( u2_out10_26 ) );
  XOR2_X1 u2_U21 (.B( u2_L1_19 ) , .Z( u2_N82 ) , .A( u2_out2_19 ) );
  XOR2_X1 u2_U210 (.B( u2_L9_24 ) , .Z( u2_N343 ) , .A( u2_out10_24 ) );
  XOR2_X1 u2_U211 (.B( u2_L9_23 ) , .Z( u2_N342 ) , .A( u2_out10_23 ) );
  XOR2_X1 u2_U215 (.B( u2_L9_20 ) , .Z( u2_N339 ) , .A( u2_out10_20 ) );
  XOR2_X1 u2_U217 (.B( u2_L9_18 ) , .Z( u2_N337 ) , .A( u2_out10_18 ) );
  XOR2_X1 u2_U218 (.B( u2_L9_17 ) , .Z( u2_N336 ) , .A( u2_out10_17 ) );
  XOR2_X1 u2_U219 (.B( u2_L9_16 ) , .Z( u2_N335 ) , .A( u2_out10_16 ) );
  XOR2_X1 u2_U222 (.B( u2_L9_13 ) , .Z( u2_N332 ) , .A( u2_out10_13 ) );
  XOR2_X1 u2_U226 (.B( u2_L9_10 ) , .Z( u2_N329 ) , .A( u2_out10_10 ) );
  XOR2_X1 u2_U227 (.B( u2_L9_9 ) , .Z( u2_N328 ) , .A( u2_out10_9 ) );
  XOR2_X1 u2_U230 (.B( u2_L9_6 ) , .Z( u2_N325 ) , .A( u2_out10_6 ) );
  XOR2_X1 u2_U234 (.B( u2_L9_2 ) , .Z( u2_N321 ) , .A( u2_out10_2 ) );
  XOR2_X1 u2_U235 (.B( u2_L9_1 ) , .Z( u2_N320 ) , .A( u2_out10_1 ) );
  XOR2_X1 u2_U26 (.B( u2_L1_15 ) , .Z( u2_N78 ) , .A( u2_out2_15 ) );
  XOR2_X1 u2_U27 (.B( u2_L1_14 ) , .Z( u2_N77 ) , .A( u2_out2_14 ) );
  XOR2_X1 u2_U29 (.B( u2_L1_12 ) , .Z( u2_N75 ) , .A( u2_out2_12 ) );
  XOR2_X1 u2_U3 (.B( u2_L2_4 ) , .Z( u2_N99 ) , .A( u2_out3_4 ) );
  XOR2_X1 u2_U30 (.B( u2_L1_11 ) , .Z( u2_N74 ) , .A( u2_out2_11 ) );
  XOR2_X1 u2_U31 (.B( u2_L1_10 ) , .Z( u2_N73 ) , .A( u2_out2_10 ) );
  XOR2_X1 u2_U33 (.B( u2_L1_8 ) , .Z( u2_N71 ) , .A( u2_out2_8 ) );
  XOR2_X1 u2_U34 (.B( u2_L1_7 ) , .Z( u2_N70 ) , .A( u2_out2_7 ) );
  XOR2_X1 u2_U37 (.B( u2_L1_5 ) , .Z( u2_N68 ) , .A( u2_out2_5 ) );
  XOR2_X1 u2_U38 (.B( u2_L1_4 ) , .Z( u2_N67 ) , .A( u2_out2_4 ) );
  XOR2_X1 u2_U380 (.B( u2_L4_31 ) , .Z( u2_N190 ) , .A( u2_out5_31 ) );
  XOR2_X1 u2_U384 (.B( u2_L4_28 ) , .Z( u2_N187 ) , .A( u2_out5_28 ) );
  XOR2_X1 u2_U385 (.B( u2_L4_27 ) , .Z( u2_N186 ) , .A( u2_out5_27 ) );
  XOR2_X1 u2_U389 (.B( u2_L4_23 ) , .Z( u2_N182 ) , .A( u2_out5_23 ) );
  XOR2_X1 u2_U39 (.B( u2_L1_3 ) , .Z( u2_N66 ) , .A( u2_out2_3 ) );
  XOR2_X1 u2_U391 (.B( u2_L4_21 ) , .Z( u2_N180 ) , .A( u2_out5_21 ) );
  XOR2_X1 u2_U395 (.B( u2_L4_18 ) , .Z( u2_N177 ) , .A( u2_out5_18 ) );
  XOR2_X1 u2_U396 (.B( u2_L4_17 ) , .Z( u2_N176 ) , .A( u2_out5_17 ) );
  XOR2_X1 u2_U398 (.B( u2_L4_15 ) , .Z( u2_N174 ) , .A( u2_out5_15 ) );
  XOR2_X1 u2_U4 (.B( u2_L2_3 ) , .Z( u2_N98 ) , .A( u2_out3_3 ) );
  XOR2_X1 u2_U400 (.B( u2_L4_13 ) , .Z( u2_N172 ) , .A( u2_out5_13 ) );
  XOR2_X1 u2_U405 (.B( u2_L4_9 ) , .Z( u2_N168 ) , .A( u2_out5_9 ) );
  XOR2_X1 u2_U409 (.B( u2_L4_5 ) , .Z( u2_N164 ) , .A( u2_out5_5 ) );
  XOR2_X1 u2_U41 (.B( u2_L1_1 ) , .Z( u2_N64 ) , .A( u2_out2_1 ) );
  XOR2_X1 u2_U412 (.B( u2_L4_2 ) , .Z( u2_N161 ) , .A( u2_out5_2 ) );
  XOR2_X1 u2_U450 (.B( u2_L2_32 ) , .Z( u2_N127 ) , .A( u2_out3_32 ) );
  XOR2_X1 u2_U453 (.B( u2_L2_29 ) , .Z( u2_N124 ) , .A( u2_out3_29 ) );
  XOR2_X1 u2_U457 (.B( u2_L2_25 ) , .Z( u2_N120 ) , .A( u2_out3_25 ) );
  XOR2_X1 u2_U461 (.B( u2_L2_22 ) , .Z( u2_N117 ) , .A( u2_out3_22 ) );
  XOR2_X1 u2_U464 (.B( u2_L2_19 ) , .Z( u2_N114 ) , .A( u2_out3_19 ) );
  XOR2_X1 u2_U470 (.B( u2_L2_14 ) , .Z( u2_N109 ) , .A( u2_out3_14 ) );
  XOR2_X1 u2_U472 (.B( u2_L2_12 ) , .Z( u2_N107 ) , .A( u2_out3_12 ) );
  XOR2_X1 u2_U473 (.B( u2_L2_11 ) , .Z( u2_N106 ) , .A( u2_out3_11 ) );
  XOR2_X1 u2_U476 (.B( u2_L2_8 ) , .Z( u2_N103 ) , .A( u2_out3_8 ) );
  XOR2_X1 u2_U477 (.B( u2_L2_7 ) , .Z( u2_N102 ) , .A( u2_out3_7 ) );
  XOR2_X1 u2_U7 (.B( u2_L1_32 ) , .Z( u2_N95 ) , .A( u2_out2_32 ) );
  XOR2_X1 u2_u10_U1 (.B( u2_K11_9 ) , .A( u2_R9_6 ) , .Z( u2_u10_X_9 ) );
  XOR2_X1 u2_u10_U16 (.B( u2_K11_3 ) , .A( u2_R9_2 ) , .Z( u2_u10_X_3 ) );
  XOR2_X1 u2_u10_U2 (.B( u2_K11_8 ) , .A( u2_R9_5 ) , .Z( u2_u10_X_8 ) );
  XOR2_X1 u2_u10_U27 (.B( u2_K11_2 ) , .A( u2_R9_1 ) , .Z( u2_u10_X_2 ) );
  XOR2_X1 u2_u10_U3 (.B( u2_K11_7 ) , .A( u2_R9_4 ) , .Z( u2_u10_X_7 ) );
  XOR2_X1 u2_u10_U33 (.B( u2_K11_24 ) , .A( u2_R9_17 ) , .Z( u2_u10_X_24 ) );
  XOR2_X1 u2_u10_U34 (.B( u2_K11_23 ) , .A( u2_R9_16 ) , .Z( u2_u10_X_23 ) );
  XOR2_X1 u2_u10_U35 (.B( u2_K11_22 ) , .A( u2_R9_15 ) , .Z( u2_u10_X_22 ) );
  XOR2_X1 u2_u10_U36 (.B( u2_K11_21 ) , .A( u2_R9_14 ) , .Z( u2_u10_X_21 ) );
  XOR2_X1 u2_u10_U37 (.B( u2_K11_20 ) , .A( u2_R9_13 ) , .Z( u2_u10_X_20 ) );
  XOR2_X1 u2_u10_U38 (.B( u2_K11_1 ) , .A( u2_R9_32 ) , .Z( u2_u10_X_1 ) );
  XOR2_X1 u2_u10_U39 (.B( u2_K11_19 ) , .A( u2_R9_12 ) , .Z( u2_u10_X_19 ) );
  XOR2_X1 u2_u10_U4 (.B( u2_K11_6 ) , .A( u2_R9_5 ) , .Z( u2_u10_X_6 ) );
  XOR2_X1 u2_u10_U40 (.B( u2_K11_18 ) , .A( u2_R9_13 ) , .Z( u2_u10_X_18 ) );
  XOR2_X1 u2_u10_U41 (.B( u2_K11_17 ) , .A( u2_R9_12 ) , .Z( u2_u10_X_17 ) );
  XOR2_X1 u2_u10_U42 (.B( u2_K11_16 ) , .A( u2_R9_11 ) , .Z( u2_u10_X_16 ) );
  XOR2_X1 u2_u10_U43 (.B( u2_K11_15 ) , .A( u2_R9_10 ) , .Z( u2_u10_X_15 ) );
  XOR2_X1 u2_u10_U44 (.B( u2_K11_14 ) , .A( u2_R9_9 ) , .Z( u2_u10_X_14 ) );
  XOR2_X1 u2_u10_U45 (.B( u2_K11_13 ) , .A( u2_R9_8 ) , .Z( u2_u10_X_13 ) );
  XOR2_X1 u2_u10_U46 (.B( u2_K11_12 ) , .A( u2_R9_9 ) , .Z( u2_u10_X_12 ) );
  XOR2_X1 u2_u10_U47 (.B( u2_K11_11 ) , .A( u2_R9_8 ) , .Z( u2_u10_X_11 ) );
  XOR2_X1 u2_u10_U48 (.B( u2_K11_10 ) , .A( u2_R9_7 ) , .Z( u2_u10_X_10 ) );
  XOR2_X1 u2_u10_U5 (.B( u2_K11_5 ) , .A( u2_R9_4 ) , .Z( u2_u10_X_5 ) );
  XOR2_X1 u2_u10_U6 (.B( u2_K11_4 ) , .A( u2_R9_3 ) , .Z( u2_u10_X_4 ) );
  AND3_X1 u2_u10_u0_U10 (.A2( u2_u10_u0_n112 ) , .ZN( u2_u10_u0_n127 ) , .A3( u2_u10_u0_n130 ) , .A1( u2_u10_u0_n148 ) );
  NAND2_X1 u2_u10_u0_U11 (.ZN( u2_u10_u0_n113 ) , .A1( u2_u10_u0_n139 ) , .A2( u2_u10_u0_n149 ) );
  AND2_X1 u2_u10_u0_U12 (.ZN( u2_u10_u0_n107 ) , .A1( u2_u10_u0_n130 ) , .A2( u2_u10_u0_n140 ) );
  AND2_X1 u2_u10_u0_U13 (.A2( u2_u10_u0_n129 ) , .A1( u2_u10_u0_n130 ) , .ZN( u2_u10_u0_n151 ) );
  AND2_X1 u2_u10_u0_U14 (.A1( u2_u10_u0_n108 ) , .A2( u2_u10_u0_n125 ) , .ZN( u2_u10_u0_n145 ) );
  INV_X1 u2_u10_u0_U15 (.A( u2_u10_u0_n143 ) , .ZN( u2_u10_u0_n173 ) );
  NOR2_X1 u2_u10_u0_U16 (.A2( u2_u10_u0_n136 ) , .ZN( u2_u10_u0_n147 ) , .A1( u2_u10_u0_n160 ) );
  NOR2_X1 u2_u10_u0_U17 (.A1( u2_u10_u0_n163 ) , .A2( u2_u10_u0_n164 ) , .ZN( u2_u10_u0_n95 ) );
  AOI21_X1 u2_u10_u0_U18 (.B1( u2_u10_u0_n103 ) , .ZN( u2_u10_u0_n132 ) , .A( u2_u10_u0_n165 ) , .B2( u2_u10_u0_n93 ) );
  INV_X1 u2_u10_u0_U19 (.A( u2_u10_u0_n142 ) , .ZN( u2_u10_u0_n165 ) );
  OAI221_X1 u2_u10_u0_U20 (.C1( u2_u10_u0_n121 ) , .ZN( u2_u10_u0_n122 ) , .B2( u2_u10_u0_n127 ) , .A( u2_u10_u0_n143 ) , .B1( u2_u10_u0_n144 ) , .C2( u2_u10_u0_n147 ) );
  OAI22_X1 u2_u10_u0_U21 (.B1( u2_u10_u0_n125 ) , .ZN( u2_u10_u0_n126 ) , .A1( u2_u10_u0_n138 ) , .A2( u2_u10_u0_n146 ) , .B2( u2_u10_u0_n147 ) );
  OAI22_X1 u2_u10_u0_U22 (.B1( u2_u10_u0_n131 ) , .A1( u2_u10_u0_n144 ) , .B2( u2_u10_u0_n147 ) , .A2( u2_u10_u0_n90 ) , .ZN( u2_u10_u0_n91 ) );
  AND3_X1 u2_u10_u0_U23 (.A3( u2_u10_u0_n121 ) , .A2( u2_u10_u0_n125 ) , .A1( u2_u10_u0_n148 ) , .ZN( u2_u10_u0_n90 ) );
  NAND2_X1 u2_u10_u0_U24 (.A1( u2_u10_u0_n100 ) , .A2( u2_u10_u0_n103 ) , .ZN( u2_u10_u0_n125 ) );
  INV_X1 u2_u10_u0_U25 (.A( u2_u10_u0_n136 ) , .ZN( u2_u10_u0_n161 ) );
  NOR2_X1 u2_u10_u0_U26 (.A1( u2_u10_u0_n120 ) , .ZN( u2_u10_u0_n143 ) , .A2( u2_u10_u0_n167 ) );
  OAI221_X1 u2_u10_u0_U27 (.C1( u2_u10_u0_n112 ) , .ZN( u2_u10_u0_n120 ) , .B1( u2_u10_u0_n138 ) , .B2( u2_u10_u0_n141 ) , .C2( u2_u10_u0_n147 ) , .A( u2_u10_u0_n172 ) );
  AOI211_X1 u2_u10_u0_U28 (.B( u2_u10_u0_n115 ) , .A( u2_u10_u0_n116 ) , .C2( u2_u10_u0_n117 ) , .C1( u2_u10_u0_n118 ) , .ZN( u2_u10_u0_n119 ) );
  AOI22_X1 u2_u10_u0_U29 (.B2( u2_u10_u0_n109 ) , .A2( u2_u10_u0_n110 ) , .ZN( u2_u10_u0_n111 ) , .B1( u2_u10_u0_n118 ) , .A1( u2_u10_u0_n160 ) );
  INV_X1 u2_u10_u0_U3 (.A( u2_u10_u0_n113 ) , .ZN( u2_u10_u0_n166 ) );
  NAND2_X1 u2_u10_u0_U30 (.A1( u2_u10_u0_n100 ) , .ZN( u2_u10_u0_n129 ) , .A2( u2_u10_u0_n95 ) );
  INV_X1 u2_u10_u0_U31 (.A( u2_u10_u0_n118 ) , .ZN( u2_u10_u0_n158 ) );
  AOI21_X1 u2_u10_u0_U32 (.ZN( u2_u10_u0_n104 ) , .B1( u2_u10_u0_n107 ) , .B2( u2_u10_u0_n141 ) , .A( u2_u10_u0_n144 ) );
  AOI21_X1 u2_u10_u0_U33 (.B1( u2_u10_u0_n127 ) , .B2( u2_u10_u0_n129 ) , .A( u2_u10_u0_n138 ) , .ZN( u2_u10_u0_n96 ) );
  AOI21_X1 u2_u10_u0_U34 (.ZN( u2_u10_u0_n116 ) , .B2( u2_u10_u0_n142 ) , .A( u2_u10_u0_n144 ) , .B1( u2_u10_u0_n166 ) );
  NAND2_X1 u2_u10_u0_U35 (.A2( u2_u10_u0_n100 ) , .A1( u2_u10_u0_n101 ) , .ZN( u2_u10_u0_n139 ) );
  NAND2_X1 u2_u10_u0_U36 (.A2( u2_u10_u0_n100 ) , .ZN( u2_u10_u0_n131 ) , .A1( u2_u10_u0_n92 ) );
  NAND2_X1 u2_u10_u0_U37 (.A1( u2_u10_u0_n101 ) , .A2( u2_u10_u0_n102 ) , .ZN( u2_u10_u0_n150 ) );
  INV_X1 u2_u10_u0_U38 (.A( u2_u10_u0_n138 ) , .ZN( u2_u10_u0_n160 ) );
  NAND2_X1 u2_u10_u0_U39 (.A1( u2_u10_u0_n102 ) , .ZN( u2_u10_u0_n128 ) , .A2( u2_u10_u0_n95 ) );
  AOI21_X1 u2_u10_u0_U4 (.B1( u2_u10_u0_n114 ) , .ZN( u2_u10_u0_n115 ) , .B2( u2_u10_u0_n129 ) , .A( u2_u10_u0_n161 ) );
  NAND2_X1 u2_u10_u0_U40 (.ZN( u2_u10_u0_n148 ) , .A1( u2_u10_u0_n93 ) , .A2( u2_u10_u0_n95 ) );
  NAND2_X1 u2_u10_u0_U41 (.A2( u2_u10_u0_n102 ) , .A1( u2_u10_u0_n103 ) , .ZN( u2_u10_u0_n149 ) );
  NAND2_X1 u2_u10_u0_U42 (.A2( u2_u10_u0_n102 ) , .ZN( u2_u10_u0_n114 ) , .A1( u2_u10_u0_n92 ) );
  NAND2_X1 u2_u10_u0_U43 (.A2( u2_u10_u0_n101 ) , .ZN( u2_u10_u0_n121 ) , .A1( u2_u10_u0_n93 ) );
  INV_X1 u2_u10_u0_U44 (.ZN( u2_u10_u0_n172 ) , .A( u2_u10_u0_n88 ) );
  OAI222_X1 u2_u10_u0_U45 (.C1( u2_u10_u0_n108 ) , .A1( u2_u10_u0_n125 ) , .B2( u2_u10_u0_n128 ) , .B1( u2_u10_u0_n144 ) , .A2( u2_u10_u0_n158 ) , .C2( u2_u10_u0_n161 ) , .ZN( u2_u10_u0_n88 ) );
  NAND2_X1 u2_u10_u0_U46 (.ZN( u2_u10_u0_n112 ) , .A2( u2_u10_u0_n92 ) , .A1( u2_u10_u0_n93 ) );
  OR3_X1 u2_u10_u0_U47 (.A3( u2_u10_u0_n152 ) , .A2( u2_u10_u0_n153 ) , .A1( u2_u10_u0_n154 ) , .ZN( u2_u10_u0_n155 ) );
  AOI21_X1 u2_u10_u0_U48 (.A( u2_u10_u0_n144 ) , .B2( u2_u10_u0_n145 ) , .B1( u2_u10_u0_n146 ) , .ZN( u2_u10_u0_n154 ) );
  AOI21_X1 u2_u10_u0_U49 (.B2( u2_u10_u0_n150 ) , .B1( u2_u10_u0_n151 ) , .ZN( u2_u10_u0_n152 ) , .A( u2_u10_u0_n158 ) );
  AOI21_X1 u2_u10_u0_U5 (.B2( u2_u10_u0_n131 ) , .ZN( u2_u10_u0_n134 ) , .B1( u2_u10_u0_n151 ) , .A( u2_u10_u0_n158 ) );
  AOI21_X1 u2_u10_u0_U50 (.A( u2_u10_u0_n147 ) , .B2( u2_u10_u0_n148 ) , .B1( u2_u10_u0_n149 ) , .ZN( u2_u10_u0_n153 ) );
  INV_X1 u2_u10_u0_U51 (.ZN( u2_u10_u0_n171 ) , .A( u2_u10_u0_n99 ) );
  OAI211_X1 u2_u10_u0_U52 (.C2( u2_u10_u0_n140 ) , .C1( u2_u10_u0_n161 ) , .A( u2_u10_u0_n169 ) , .B( u2_u10_u0_n98 ) , .ZN( u2_u10_u0_n99 ) );
  AOI211_X1 u2_u10_u0_U53 (.C1( u2_u10_u0_n118 ) , .A( u2_u10_u0_n123 ) , .B( u2_u10_u0_n96 ) , .C2( u2_u10_u0_n97 ) , .ZN( u2_u10_u0_n98 ) );
  INV_X1 u2_u10_u0_U54 (.ZN( u2_u10_u0_n169 ) , .A( u2_u10_u0_n91 ) );
  NOR2_X1 u2_u10_u0_U55 (.A2( u2_u10_X_4 ) , .A1( u2_u10_X_5 ) , .ZN( u2_u10_u0_n118 ) );
  NOR2_X1 u2_u10_u0_U56 (.A2( u2_u10_X_2 ) , .ZN( u2_u10_u0_n103 ) , .A1( u2_u10_u0_n164 ) );
  NOR2_X1 u2_u10_u0_U57 (.A2( u2_u10_X_1 ) , .A1( u2_u10_X_2 ) , .ZN( u2_u10_u0_n92 ) );
  NOR2_X1 u2_u10_u0_U58 (.A2( u2_u10_X_1 ) , .ZN( u2_u10_u0_n101 ) , .A1( u2_u10_u0_n163 ) );
  NAND2_X1 u2_u10_u0_U59 (.A2( u2_u10_X_4 ) , .A1( u2_u10_X_5 ) , .ZN( u2_u10_u0_n144 ) );
  NOR2_X1 u2_u10_u0_U6 (.A1( u2_u10_u0_n108 ) , .ZN( u2_u10_u0_n123 ) , .A2( u2_u10_u0_n158 ) );
  NOR2_X1 u2_u10_u0_U60 (.A2( u2_u10_X_5 ) , .ZN( u2_u10_u0_n136 ) , .A1( u2_u10_u0_n159 ) );
  NAND2_X1 u2_u10_u0_U61 (.A1( u2_u10_X_5 ) , .ZN( u2_u10_u0_n138 ) , .A2( u2_u10_u0_n159 ) );
  AND2_X1 u2_u10_u0_U62 (.A2( u2_u10_X_3 ) , .A1( u2_u10_X_6 ) , .ZN( u2_u10_u0_n102 ) );
  AND2_X1 u2_u10_u0_U63 (.A1( u2_u10_X_6 ) , .A2( u2_u10_u0_n162 ) , .ZN( u2_u10_u0_n93 ) );
  INV_X1 u2_u10_u0_U64 (.A( u2_u10_X_4 ) , .ZN( u2_u10_u0_n159 ) );
  INV_X1 u2_u10_u0_U65 (.A( u2_u10_X_1 ) , .ZN( u2_u10_u0_n164 ) );
  INV_X1 u2_u10_u0_U66 (.A( u2_u10_X_2 ) , .ZN( u2_u10_u0_n163 ) );
  INV_X1 u2_u10_u0_U67 (.A( u2_u10_X_3 ) , .ZN( u2_u10_u0_n162 ) );
  INV_X1 u2_u10_u0_U68 (.A( u2_u10_u0_n126 ) , .ZN( u2_u10_u0_n168 ) );
  AOI211_X1 u2_u10_u0_U69 (.B( u2_u10_u0_n133 ) , .A( u2_u10_u0_n134 ) , .C2( u2_u10_u0_n135 ) , .C1( u2_u10_u0_n136 ) , .ZN( u2_u10_u0_n137 ) );
  OAI21_X1 u2_u10_u0_U7 (.B1( u2_u10_u0_n150 ) , .B2( u2_u10_u0_n158 ) , .A( u2_u10_u0_n172 ) , .ZN( u2_u10_u0_n89 ) );
  INV_X1 u2_u10_u0_U70 (.ZN( u2_u10_u0_n174 ) , .A( u2_u10_u0_n89 ) );
  AOI211_X1 u2_u10_u0_U71 (.B( u2_u10_u0_n104 ) , .A( u2_u10_u0_n105 ) , .ZN( u2_u10_u0_n106 ) , .C2( u2_u10_u0_n113 ) , .C1( u2_u10_u0_n160 ) );
  OR4_X1 u2_u10_u0_U72 (.ZN( u2_out10_17 ) , .A4( u2_u10_u0_n122 ) , .A2( u2_u10_u0_n123 ) , .A1( u2_u10_u0_n124 ) , .A3( u2_u10_u0_n170 ) );
  AOI21_X1 u2_u10_u0_U73 (.B2( u2_u10_u0_n107 ) , .ZN( u2_u10_u0_n124 ) , .B1( u2_u10_u0_n128 ) , .A( u2_u10_u0_n161 ) );
  INV_X1 u2_u10_u0_U74 (.A( u2_u10_u0_n111 ) , .ZN( u2_u10_u0_n170 ) );
  OR4_X1 u2_u10_u0_U75 (.ZN( u2_out10_31 ) , .A4( u2_u10_u0_n155 ) , .A2( u2_u10_u0_n156 ) , .A1( u2_u10_u0_n157 ) , .A3( u2_u10_u0_n173 ) );
  AOI21_X1 u2_u10_u0_U76 (.A( u2_u10_u0_n138 ) , .B2( u2_u10_u0_n139 ) , .B1( u2_u10_u0_n140 ) , .ZN( u2_u10_u0_n157 ) );
  AOI21_X1 u2_u10_u0_U77 (.B2( u2_u10_u0_n141 ) , .B1( u2_u10_u0_n142 ) , .ZN( u2_u10_u0_n156 ) , .A( u2_u10_u0_n161 ) );
  AOI21_X1 u2_u10_u0_U78 (.B1( u2_u10_u0_n132 ) , .ZN( u2_u10_u0_n133 ) , .A( u2_u10_u0_n144 ) , .B2( u2_u10_u0_n166 ) );
  OAI22_X1 u2_u10_u0_U79 (.ZN( u2_u10_u0_n105 ) , .A2( u2_u10_u0_n132 ) , .B1( u2_u10_u0_n146 ) , .A1( u2_u10_u0_n147 ) , .B2( u2_u10_u0_n161 ) );
  AND2_X1 u2_u10_u0_U8 (.A1( u2_u10_u0_n114 ) , .A2( u2_u10_u0_n121 ) , .ZN( u2_u10_u0_n146 ) );
  NAND2_X1 u2_u10_u0_U80 (.ZN( u2_u10_u0_n110 ) , .A2( u2_u10_u0_n132 ) , .A1( u2_u10_u0_n145 ) );
  INV_X1 u2_u10_u0_U81 (.A( u2_u10_u0_n119 ) , .ZN( u2_u10_u0_n167 ) );
  NAND2_X1 u2_u10_u0_U82 (.A2( u2_u10_u0_n103 ) , .ZN( u2_u10_u0_n140 ) , .A1( u2_u10_u0_n94 ) );
  NAND2_X1 u2_u10_u0_U83 (.A1( u2_u10_u0_n101 ) , .ZN( u2_u10_u0_n130 ) , .A2( u2_u10_u0_n94 ) );
  NAND2_X1 u2_u10_u0_U84 (.ZN( u2_u10_u0_n108 ) , .A1( u2_u10_u0_n92 ) , .A2( u2_u10_u0_n94 ) );
  NAND2_X1 u2_u10_u0_U85 (.ZN( u2_u10_u0_n142 ) , .A1( u2_u10_u0_n94 ) , .A2( u2_u10_u0_n95 ) );
  NOR2_X1 u2_u10_u0_U86 (.A2( u2_u10_X_6 ) , .ZN( u2_u10_u0_n100 ) , .A1( u2_u10_u0_n162 ) );
  NOR2_X1 u2_u10_u0_U87 (.A2( u2_u10_X_3 ) , .A1( u2_u10_X_6 ) , .ZN( u2_u10_u0_n94 ) );
  NAND3_X1 u2_u10_u0_U88 (.ZN( u2_out10_23 ) , .A3( u2_u10_u0_n137 ) , .A1( u2_u10_u0_n168 ) , .A2( u2_u10_u0_n171 ) );
  NAND3_X1 u2_u10_u0_U89 (.A3( u2_u10_u0_n127 ) , .A2( u2_u10_u0_n128 ) , .ZN( u2_u10_u0_n135 ) , .A1( u2_u10_u0_n150 ) );
  AND2_X1 u2_u10_u0_U9 (.A1( u2_u10_u0_n131 ) , .ZN( u2_u10_u0_n141 ) , .A2( u2_u10_u0_n150 ) );
  NAND3_X1 u2_u10_u0_U90 (.ZN( u2_u10_u0_n117 ) , .A3( u2_u10_u0_n132 ) , .A2( u2_u10_u0_n139 ) , .A1( u2_u10_u0_n148 ) );
  NAND3_X1 u2_u10_u0_U91 (.ZN( u2_u10_u0_n109 ) , .A2( u2_u10_u0_n114 ) , .A3( u2_u10_u0_n140 ) , .A1( u2_u10_u0_n149 ) );
  NAND3_X1 u2_u10_u0_U92 (.ZN( u2_out10_9 ) , .A3( u2_u10_u0_n106 ) , .A2( u2_u10_u0_n171 ) , .A1( u2_u10_u0_n174 ) );
  NAND3_X1 u2_u10_u0_U93 (.A2( u2_u10_u0_n128 ) , .A1( u2_u10_u0_n132 ) , .A3( u2_u10_u0_n146 ) , .ZN( u2_u10_u0_n97 ) );
  AOI21_X1 u2_u10_u1_U10 (.B2( u2_u10_u1_n155 ) , .B1( u2_u10_u1_n156 ) , .ZN( u2_u10_u1_n157 ) , .A( u2_u10_u1_n174 ) );
  NAND3_X1 u2_u10_u1_U100 (.ZN( u2_u10_u1_n113 ) , .A1( u2_u10_u1_n120 ) , .A3( u2_u10_u1_n133 ) , .A2( u2_u10_u1_n155 ) );
  NAND2_X1 u2_u10_u1_U11 (.ZN( u2_u10_u1_n140 ) , .A2( u2_u10_u1_n150 ) , .A1( u2_u10_u1_n155 ) );
  NAND2_X1 u2_u10_u1_U12 (.A1( u2_u10_u1_n131 ) , .ZN( u2_u10_u1_n147 ) , .A2( u2_u10_u1_n153 ) );
  AOI22_X1 u2_u10_u1_U13 (.B2( u2_u10_u1_n136 ) , .A2( u2_u10_u1_n137 ) , .ZN( u2_u10_u1_n143 ) , .A1( u2_u10_u1_n171 ) , .B1( u2_u10_u1_n173 ) );
  INV_X1 u2_u10_u1_U14 (.A( u2_u10_u1_n147 ) , .ZN( u2_u10_u1_n181 ) );
  INV_X1 u2_u10_u1_U15 (.A( u2_u10_u1_n139 ) , .ZN( u2_u10_u1_n174 ) );
  OR4_X1 u2_u10_u1_U16 (.A4( u2_u10_u1_n106 ) , .A3( u2_u10_u1_n107 ) , .ZN( u2_u10_u1_n108 ) , .A1( u2_u10_u1_n117 ) , .A2( u2_u10_u1_n184 ) );
  AOI21_X1 u2_u10_u1_U17 (.ZN( u2_u10_u1_n106 ) , .A( u2_u10_u1_n112 ) , .B1( u2_u10_u1_n154 ) , .B2( u2_u10_u1_n156 ) );
  AOI21_X1 u2_u10_u1_U18 (.ZN( u2_u10_u1_n107 ) , .B1( u2_u10_u1_n134 ) , .B2( u2_u10_u1_n149 ) , .A( u2_u10_u1_n174 ) );
  INV_X1 u2_u10_u1_U19 (.A( u2_u10_u1_n101 ) , .ZN( u2_u10_u1_n184 ) );
  INV_X1 u2_u10_u1_U20 (.A( u2_u10_u1_n112 ) , .ZN( u2_u10_u1_n171 ) );
  NAND2_X1 u2_u10_u1_U21 (.ZN( u2_u10_u1_n141 ) , .A1( u2_u10_u1_n153 ) , .A2( u2_u10_u1_n156 ) );
  AND2_X1 u2_u10_u1_U22 (.A1( u2_u10_u1_n123 ) , .ZN( u2_u10_u1_n134 ) , .A2( u2_u10_u1_n161 ) );
  NAND2_X1 u2_u10_u1_U23 (.A2( u2_u10_u1_n115 ) , .A1( u2_u10_u1_n116 ) , .ZN( u2_u10_u1_n148 ) );
  NAND2_X1 u2_u10_u1_U24 (.A2( u2_u10_u1_n133 ) , .A1( u2_u10_u1_n135 ) , .ZN( u2_u10_u1_n159 ) );
  NAND2_X1 u2_u10_u1_U25 (.A2( u2_u10_u1_n115 ) , .A1( u2_u10_u1_n120 ) , .ZN( u2_u10_u1_n132 ) );
  INV_X1 u2_u10_u1_U26 (.A( u2_u10_u1_n154 ) , .ZN( u2_u10_u1_n178 ) );
  INV_X1 u2_u10_u1_U27 (.A( u2_u10_u1_n151 ) , .ZN( u2_u10_u1_n183 ) );
  AND2_X1 u2_u10_u1_U28 (.A1( u2_u10_u1_n129 ) , .A2( u2_u10_u1_n133 ) , .ZN( u2_u10_u1_n149 ) );
  INV_X1 u2_u10_u1_U29 (.A( u2_u10_u1_n131 ) , .ZN( u2_u10_u1_n180 ) );
  INV_X1 u2_u10_u1_U3 (.A( u2_u10_u1_n159 ) , .ZN( u2_u10_u1_n182 ) );
  OAI221_X1 u2_u10_u1_U30 (.A( u2_u10_u1_n119 ) , .C2( u2_u10_u1_n129 ) , .ZN( u2_u10_u1_n138 ) , .B2( u2_u10_u1_n152 ) , .C1( u2_u10_u1_n174 ) , .B1( u2_u10_u1_n187 ) );
  INV_X1 u2_u10_u1_U31 (.A( u2_u10_u1_n148 ) , .ZN( u2_u10_u1_n187 ) );
  AOI211_X1 u2_u10_u1_U32 (.B( u2_u10_u1_n117 ) , .A( u2_u10_u1_n118 ) , .ZN( u2_u10_u1_n119 ) , .C2( u2_u10_u1_n146 ) , .C1( u2_u10_u1_n159 ) );
  NOR2_X1 u2_u10_u1_U33 (.A1( u2_u10_u1_n168 ) , .A2( u2_u10_u1_n176 ) , .ZN( u2_u10_u1_n98 ) );
  OAI21_X1 u2_u10_u1_U34 (.B2( u2_u10_u1_n123 ) , .ZN( u2_u10_u1_n145 ) , .B1( u2_u10_u1_n160 ) , .A( u2_u10_u1_n185 ) );
  INV_X1 u2_u10_u1_U35 (.A( u2_u10_u1_n122 ) , .ZN( u2_u10_u1_n185 ) );
  AOI21_X1 u2_u10_u1_U36 (.B2( u2_u10_u1_n120 ) , .B1( u2_u10_u1_n121 ) , .ZN( u2_u10_u1_n122 ) , .A( u2_u10_u1_n128 ) );
  NAND2_X1 u2_u10_u1_U37 (.A1( u2_u10_u1_n128 ) , .ZN( u2_u10_u1_n146 ) , .A2( u2_u10_u1_n160 ) );
  NAND2_X1 u2_u10_u1_U38 (.A2( u2_u10_u1_n112 ) , .ZN( u2_u10_u1_n139 ) , .A1( u2_u10_u1_n152 ) );
  NAND2_X1 u2_u10_u1_U39 (.A1( u2_u10_u1_n105 ) , .ZN( u2_u10_u1_n156 ) , .A2( u2_u10_u1_n99 ) );
  AOI221_X1 u2_u10_u1_U4 (.A( u2_u10_u1_n138 ) , .C2( u2_u10_u1_n139 ) , .C1( u2_u10_u1_n140 ) , .B2( u2_u10_u1_n141 ) , .ZN( u2_u10_u1_n142 ) , .B1( u2_u10_u1_n175 ) );
  AOI221_X1 u2_u10_u1_U40 (.B1( u2_u10_u1_n140 ) , .ZN( u2_u10_u1_n167 ) , .B2( u2_u10_u1_n172 ) , .C2( u2_u10_u1_n175 ) , .C1( u2_u10_u1_n178 ) , .A( u2_u10_u1_n188 ) );
  INV_X1 u2_u10_u1_U41 (.ZN( u2_u10_u1_n188 ) , .A( u2_u10_u1_n97 ) );
  AOI211_X1 u2_u10_u1_U42 (.A( u2_u10_u1_n118 ) , .C1( u2_u10_u1_n132 ) , .C2( u2_u10_u1_n139 ) , .B( u2_u10_u1_n96 ) , .ZN( u2_u10_u1_n97 ) );
  AOI21_X1 u2_u10_u1_U43 (.B2( u2_u10_u1_n121 ) , .B1( u2_u10_u1_n135 ) , .A( u2_u10_u1_n152 ) , .ZN( u2_u10_u1_n96 ) );
  NOR2_X1 u2_u10_u1_U44 (.ZN( u2_u10_u1_n117 ) , .A1( u2_u10_u1_n121 ) , .A2( u2_u10_u1_n160 ) );
  AOI21_X1 u2_u10_u1_U45 (.A( u2_u10_u1_n128 ) , .B2( u2_u10_u1_n129 ) , .ZN( u2_u10_u1_n130 ) , .B1( u2_u10_u1_n150 ) );
  NAND2_X1 u2_u10_u1_U46 (.ZN( u2_u10_u1_n112 ) , .A1( u2_u10_u1_n169 ) , .A2( u2_u10_u1_n170 ) );
  NAND2_X1 u2_u10_u1_U47 (.ZN( u2_u10_u1_n129 ) , .A2( u2_u10_u1_n95 ) , .A1( u2_u10_u1_n98 ) );
  NAND2_X1 u2_u10_u1_U48 (.A1( u2_u10_u1_n102 ) , .ZN( u2_u10_u1_n154 ) , .A2( u2_u10_u1_n99 ) );
  NAND2_X1 u2_u10_u1_U49 (.A2( u2_u10_u1_n100 ) , .ZN( u2_u10_u1_n135 ) , .A1( u2_u10_u1_n99 ) );
  AOI211_X1 u2_u10_u1_U5 (.ZN( u2_u10_u1_n124 ) , .A( u2_u10_u1_n138 ) , .C2( u2_u10_u1_n139 ) , .B( u2_u10_u1_n145 ) , .C1( u2_u10_u1_n147 ) );
  AOI21_X1 u2_u10_u1_U50 (.A( u2_u10_u1_n152 ) , .B2( u2_u10_u1_n153 ) , .B1( u2_u10_u1_n154 ) , .ZN( u2_u10_u1_n158 ) );
  INV_X1 u2_u10_u1_U51 (.A( u2_u10_u1_n160 ) , .ZN( u2_u10_u1_n175 ) );
  NAND2_X1 u2_u10_u1_U52 (.A1( u2_u10_u1_n100 ) , .ZN( u2_u10_u1_n116 ) , .A2( u2_u10_u1_n95 ) );
  NAND2_X1 u2_u10_u1_U53 (.A1( u2_u10_u1_n102 ) , .ZN( u2_u10_u1_n131 ) , .A2( u2_u10_u1_n95 ) );
  NAND2_X1 u2_u10_u1_U54 (.A2( u2_u10_u1_n104 ) , .ZN( u2_u10_u1_n121 ) , .A1( u2_u10_u1_n98 ) );
  NAND2_X1 u2_u10_u1_U55 (.A1( u2_u10_u1_n103 ) , .ZN( u2_u10_u1_n153 ) , .A2( u2_u10_u1_n98 ) );
  NAND2_X1 u2_u10_u1_U56 (.A2( u2_u10_u1_n104 ) , .A1( u2_u10_u1_n105 ) , .ZN( u2_u10_u1_n133 ) );
  NAND2_X1 u2_u10_u1_U57 (.ZN( u2_u10_u1_n150 ) , .A2( u2_u10_u1_n98 ) , .A1( u2_u10_u1_n99 ) );
  NAND2_X1 u2_u10_u1_U58 (.A1( u2_u10_u1_n105 ) , .ZN( u2_u10_u1_n155 ) , .A2( u2_u10_u1_n95 ) );
  OAI21_X1 u2_u10_u1_U59 (.ZN( u2_u10_u1_n109 ) , .B1( u2_u10_u1_n129 ) , .B2( u2_u10_u1_n160 ) , .A( u2_u10_u1_n167 ) );
  AOI22_X1 u2_u10_u1_U6 (.B2( u2_u10_u1_n113 ) , .A2( u2_u10_u1_n114 ) , .ZN( u2_u10_u1_n125 ) , .A1( u2_u10_u1_n171 ) , .B1( u2_u10_u1_n173 ) );
  NAND2_X1 u2_u10_u1_U60 (.A2( u2_u10_u1_n100 ) , .A1( u2_u10_u1_n103 ) , .ZN( u2_u10_u1_n120 ) );
  NAND2_X1 u2_u10_u1_U61 (.A1( u2_u10_u1_n102 ) , .A2( u2_u10_u1_n104 ) , .ZN( u2_u10_u1_n115 ) );
  NAND2_X1 u2_u10_u1_U62 (.A2( u2_u10_u1_n100 ) , .A1( u2_u10_u1_n104 ) , .ZN( u2_u10_u1_n151 ) );
  NAND2_X1 u2_u10_u1_U63 (.A2( u2_u10_u1_n103 ) , .A1( u2_u10_u1_n105 ) , .ZN( u2_u10_u1_n161 ) );
  INV_X1 u2_u10_u1_U64 (.A( u2_u10_u1_n152 ) , .ZN( u2_u10_u1_n173 ) );
  INV_X1 u2_u10_u1_U65 (.A( u2_u10_u1_n128 ) , .ZN( u2_u10_u1_n172 ) );
  NAND2_X1 u2_u10_u1_U66 (.A2( u2_u10_u1_n102 ) , .A1( u2_u10_u1_n103 ) , .ZN( u2_u10_u1_n123 ) );
  AOI211_X1 u2_u10_u1_U67 (.B( u2_u10_u1_n162 ) , .A( u2_u10_u1_n163 ) , .C2( u2_u10_u1_n164 ) , .ZN( u2_u10_u1_n165 ) , .C1( u2_u10_u1_n171 ) );
  AOI21_X1 u2_u10_u1_U68 (.A( u2_u10_u1_n160 ) , .B2( u2_u10_u1_n161 ) , .ZN( u2_u10_u1_n162 ) , .B1( u2_u10_u1_n182 ) );
  OR2_X1 u2_u10_u1_U69 (.A2( u2_u10_u1_n157 ) , .A1( u2_u10_u1_n158 ) , .ZN( u2_u10_u1_n163 ) );
  NAND2_X1 u2_u10_u1_U7 (.ZN( u2_u10_u1_n114 ) , .A1( u2_u10_u1_n134 ) , .A2( u2_u10_u1_n156 ) );
  NOR2_X1 u2_u10_u1_U70 (.A2( u2_u10_X_7 ) , .A1( u2_u10_X_8 ) , .ZN( u2_u10_u1_n95 ) );
  NOR2_X1 u2_u10_u1_U71 (.A1( u2_u10_X_12 ) , .A2( u2_u10_X_9 ) , .ZN( u2_u10_u1_n100 ) );
  NOR2_X1 u2_u10_u1_U72 (.A2( u2_u10_X_8 ) , .A1( u2_u10_u1_n177 ) , .ZN( u2_u10_u1_n99 ) );
  NOR2_X1 u2_u10_u1_U73 (.A2( u2_u10_X_12 ) , .ZN( u2_u10_u1_n102 ) , .A1( u2_u10_u1_n176 ) );
  NOR2_X1 u2_u10_u1_U74 (.A2( u2_u10_X_9 ) , .ZN( u2_u10_u1_n105 ) , .A1( u2_u10_u1_n168 ) );
  NAND2_X1 u2_u10_u1_U75 (.A1( u2_u10_X_10 ) , .ZN( u2_u10_u1_n160 ) , .A2( u2_u10_u1_n169 ) );
  NAND2_X1 u2_u10_u1_U76 (.A2( u2_u10_X_10 ) , .A1( u2_u10_X_11 ) , .ZN( u2_u10_u1_n152 ) );
  NAND2_X1 u2_u10_u1_U77 (.A1( u2_u10_X_11 ) , .ZN( u2_u10_u1_n128 ) , .A2( u2_u10_u1_n170 ) );
  AND2_X1 u2_u10_u1_U78 (.A2( u2_u10_X_7 ) , .A1( u2_u10_X_8 ) , .ZN( u2_u10_u1_n104 ) );
  AND2_X1 u2_u10_u1_U79 (.A1( u2_u10_X_8 ) , .ZN( u2_u10_u1_n103 ) , .A2( u2_u10_u1_n177 ) );
  NOR2_X1 u2_u10_u1_U8 (.A1( u2_u10_u1_n112 ) , .A2( u2_u10_u1_n116 ) , .ZN( u2_u10_u1_n118 ) );
  INV_X1 u2_u10_u1_U80 (.A( u2_u10_X_10 ) , .ZN( u2_u10_u1_n170 ) );
  INV_X1 u2_u10_u1_U81 (.A( u2_u10_X_9 ) , .ZN( u2_u10_u1_n176 ) );
  INV_X1 u2_u10_u1_U82 (.A( u2_u10_X_11 ) , .ZN( u2_u10_u1_n169 ) );
  INV_X1 u2_u10_u1_U83 (.A( u2_u10_X_12 ) , .ZN( u2_u10_u1_n168 ) );
  INV_X1 u2_u10_u1_U84 (.A( u2_u10_X_7 ) , .ZN( u2_u10_u1_n177 ) );
  NAND4_X1 u2_u10_u1_U85 (.ZN( u2_out10_28 ) , .A4( u2_u10_u1_n124 ) , .A3( u2_u10_u1_n125 ) , .A2( u2_u10_u1_n126 ) , .A1( u2_u10_u1_n127 ) );
  OAI21_X1 u2_u10_u1_U86 (.ZN( u2_u10_u1_n127 ) , .B2( u2_u10_u1_n139 ) , .B1( u2_u10_u1_n175 ) , .A( u2_u10_u1_n183 ) );
  OAI21_X1 u2_u10_u1_U87 (.ZN( u2_u10_u1_n126 ) , .B2( u2_u10_u1_n140 ) , .A( u2_u10_u1_n146 ) , .B1( u2_u10_u1_n178 ) );
  NAND4_X1 u2_u10_u1_U88 (.ZN( u2_out10_18 ) , .A4( u2_u10_u1_n165 ) , .A3( u2_u10_u1_n166 ) , .A1( u2_u10_u1_n167 ) , .A2( u2_u10_u1_n186 ) );
  AOI22_X1 u2_u10_u1_U89 (.B2( u2_u10_u1_n146 ) , .B1( u2_u10_u1_n147 ) , .A2( u2_u10_u1_n148 ) , .ZN( u2_u10_u1_n166 ) , .A1( u2_u10_u1_n172 ) );
  OAI21_X1 u2_u10_u1_U9 (.ZN( u2_u10_u1_n101 ) , .B1( u2_u10_u1_n141 ) , .A( u2_u10_u1_n146 ) , .B2( u2_u10_u1_n183 ) );
  INV_X1 u2_u10_u1_U90 (.A( u2_u10_u1_n145 ) , .ZN( u2_u10_u1_n186 ) );
  NAND4_X1 u2_u10_u1_U91 (.ZN( u2_out10_2 ) , .A4( u2_u10_u1_n142 ) , .A3( u2_u10_u1_n143 ) , .A2( u2_u10_u1_n144 ) , .A1( u2_u10_u1_n179 ) );
  OAI21_X1 u2_u10_u1_U92 (.B2( u2_u10_u1_n132 ) , .ZN( u2_u10_u1_n144 ) , .A( u2_u10_u1_n146 ) , .B1( u2_u10_u1_n180 ) );
  INV_X1 u2_u10_u1_U93 (.A( u2_u10_u1_n130 ) , .ZN( u2_u10_u1_n179 ) );
  OR4_X1 u2_u10_u1_U94 (.ZN( u2_out10_13 ) , .A4( u2_u10_u1_n108 ) , .A3( u2_u10_u1_n109 ) , .A2( u2_u10_u1_n110 ) , .A1( u2_u10_u1_n111 ) );
  AOI21_X1 u2_u10_u1_U95 (.ZN( u2_u10_u1_n111 ) , .A( u2_u10_u1_n128 ) , .B2( u2_u10_u1_n131 ) , .B1( u2_u10_u1_n135 ) );
  AOI21_X1 u2_u10_u1_U96 (.ZN( u2_u10_u1_n110 ) , .A( u2_u10_u1_n116 ) , .B1( u2_u10_u1_n152 ) , .B2( u2_u10_u1_n160 ) );
  NAND3_X1 u2_u10_u1_U97 (.A3( u2_u10_u1_n149 ) , .A2( u2_u10_u1_n150 ) , .A1( u2_u10_u1_n151 ) , .ZN( u2_u10_u1_n164 ) );
  NAND3_X1 u2_u10_u1_U98 (.A3( u2_u10_u1_n134 ) , .A2( u2_u10_u1_n135 ) , .ZN( u2_u10_u1_n136 ) , .A1( u2_u10_u1_n151 ) );
  NAND3_X1 u2_u10_u1_U99 (.A1( u2_u10_u1_n133 ) , .ZN( u2_u10_u1_n137 ) , .A2( u2_u10_u1_n154 ) , .A3( u2_u10_u1_n181 ) );
  OAI22_X1 u2_u10_u2_U10 (.ZN( u2_u10_u2_n109 ) , .A2( u2_u10_u2_n113 ) , .B2( u2_u10_u2_n133 ) , .B1( u2_u10_u2_n167 ) , .A1( u2_u10_u2_n168 ) );
  NAND3_X1 u2_u10_u2_U100 (.A2( u2_u10_u2_n100 ) , .A1( u2_u10_u2_n104 ) , .A3( u2_u10_u2_n138 ) , .ZN( u2_u10_u2_n98 ) );
  OAI22_X1 u2_u10_u2_U11 (.B1( u2_u10_u2_n151 ) , .A2( u2_u10_u2_n152 ) , .A1( u2_u10_u2_n153 ) , .ZN( u2_u10_u2_n160 ) , .B2( u2_u10_u2_n168 ) );
  NOR3_X1 u2_u10_u2_U12 (.A1( u2_u10_u2_n150 ) , .ZN( u2_u10_u2_n151 ) , .A3( u2_u10_u2_n175 ) , .A2( u2_u10_u2_n188 ) );
  AOI21_X1 u2_u10_u2_U13 (.ZN( u2_u10_u2_n144 ) , .B2( u2_u10_u2_n155 ) , .A( u2_u10_u2_n172 ) , .B1( u2_u10_u2_n185 ) );
  AOI21_X1 u2_u10_u2_U14 (.B2( u2_u10_u2_n143 ) , .ZN( u2_u10_u2_n145 ) , .B1( u2_u10_u2_n152 ) , .A( u2_u10_u2_n171 ) );
  AOI21_X1 u2_u10_u2_U15 (.B2( u2_u10_u2_n120 ) , .B1( u2_u10_u2_n121 ) , .ZN( u2_u10_u2_n126 ) , .A( u2_u10_u2_n167 ) );
  INV_X1 u2_u10_u2_U16 (.A( u2_u10_u2_n156 ) , .ZN( u2_u10_u2_n171 ) );
  INV_X1 u2_u10_u2_U17 (.A( u2_u10_u2_n120 ) , .ZN( u2_u10_u2_n188 ) );
  NAND2_X1 u2_u10_u2_U18 (.A2( u2_u10_u2_n122 ) , .ZN( u2_u10_u2_n150 ) , .A1( u2_u10_u2_n152 ) );
  INV_X1 u2_u10_u2_U19 (.A( u2_u10_u2_n153 ) , .ZN( u2_u10_u2_n170 ) );
  INV_X1 u2_u10_u2_U20 (.A( u2_u10_u2_n137 ) , .ZN( u2_u10_u2_n173 ) );
  NAND2_X1 u2_u10_u2_U21 (.A1( u2_u10_u2_n132 ) , .A2( u2_u10_u2_n139 ) , .ZN( u2_u10_u2_n157 ) );
  INV_X1 u2_u10_u2_U22 (.A( u2_u10_u2_n113 ) , .ZN( u2_u10_u2_n178 ) );
  INV_X1 u2_u10_u2_U23 (.A( u2_u10_u2_n139 ) , .ZN( u2_u10_u2_n175 ) );
  INV_X1 u2_u10_u2_U24 (.A( u2_u10_u2_n155 ) , .ZN( u2_u10_u2_n181 ) );
  INV_X1 u2_u10_u2_U25 (.A( u2_u10_u2_n119 ) , .ZN( u2_u10_u2_n177 ) );
  INV_X1 u2_u10_u2_U26 (.A( u2_u10_u2_n116 ) , .ZN( u2_u10_u2_n180 ) );
  INV_X1 u2_u10_u2_U27 (.A( u2_u10_u2_n131 ) , .ZN( u2_u10_u2_n179 ) );
  INV_X1 u2_u10_u2_U28 (.A( u2_u10_u2_n154 ) , .ZN( u2_u10_u2_n176 ) );
  NAND2_X1 u2_u10_u2_U29 (.A2( u2_u10_u2_n116 ) , .A1( u2_u10_u2_n117 ) , .ZN( u2_u10_u2_n118 ) );
  NOR2_X1 u2_u10_u2_U3 (.ZN( u2_u10_u2_n121 ) , .A2( u2_u10_u2_n177 ) , .A1( u2_u10_u2_n180 ) );
  INV_X1 u2_u10_u2_U30 (.A( u2_u10_u2_n132 ) , .ZN( u2_u10_u2_n182 ) );
  INV_X1 u2_u10_u2_U31 (.A( u2_u10_u2_n158 ) , .ZN( u2_u10_u2_n183 ) );
  OAI21_X1 u2_u10_u2_U32 (.A( u2_u10_u2_n156 ) , .B1( u2_u10_u2_n157 ) , .ZN( u2_u10_u2_n158 ) , .B2( u2_u10_u2_n179 ) );
  NOR2_X1 u2_u10_u2_U33 (.ZN( u2_u10_u2_n156 ) , .A1( u2_u10_u2_n166 ) , .A2( u2_u10_u2_n169 ) );
  NOR2_X1 u2_u10_u2_U34 (.A2( u2_u10_u2_n114 ) , .ZN( u2_u10_u2_n137 ) , .A1( u2_u10_u2_n140 ) );
  NOR2_X1 u2_u10_u2_U35 (.A2( u2_u10_u2_n138 ) , .ZN( u2_u10_u2_n153 ) , .A1( u2_u10_u2_n156 ) );
  AOI211_X1 u2_u10_u2_U36 (.ZN( u2_u10_u2_n130 ) , .C1( u2_u10_u2_n138 ) , .C2( u2_u10_u2_n179 ) , .B( u2_u10_u2_n96 ) , .A( u2_u10_u2_n97 ) );
  OAI22_X1 u2_u10_u2_U37 (.B1( u2_u10_u2_n133 ) , .A2( u2_u10_u2_n137 ) , .A1( u2_u10_u2_n152 ) , .B2( u2_u10_u2_n168 ) , .ZN( u2_u10_u2_n97 ) );
  OAI221_X1 u2_u10_u2_U38 (.B1( u2_u10_u2_n113 ) , .C1( u2_u10_u2_n132 ) , .A( u2_u10_u2_n149 ) , .B2( u2_u10_u2_n171 ) , .C2( u2_u10_u2_n172 ) , .ZN( u2_u10_u2_n96 ) );
  OAI221_X1 u2_u10_u2_U39 (.A( u2_u10_u2_n115 ) , .C2( u2_u10_u2_n123 ) , .B2( u2_u10_u2_n143 ) , .B1( u2_u10_u2_n153 ) , .ZN( u2_u10_u2_n163 ) , .C1( u2_u10_u2_n168 ) );
  INV_X1 u2_u10_u2_U4 (.A( u2_u10_u2_n134 ) , .ZN( u2_u10_u2_n185 ) );
  OAI21_X1 u2_u10_u2_U40 (.A( u2_u10_u2_n114 ) , .ZN( u2_u10_u2_n115 ) , .B1( u2_u10_u2_n176 ) , .B2( u2_u10_u2_n178 ) );
  OAI221_X1 u2_u10_u2_U41 (.A( u2_u10_u2_n135 ) , .B2( u2_u10_u2_n136 ) , .B1( u2_u10_u2_n137 ) , .ZN( u2_u10_u2_n162 ) , .C2( u2_u10_u2_n167 ) , .C1( u2_u10_u2_n185 ) );
  AND3_X1 u2_u10_u2_U42 (.A3( u2_u10_u2_n131 ) , .A2( u2_u10_u2_n132 ) , .A1( u2_u10_u2_n133 ) , .ZN( u2_u10_u2_n136 ) );
  AOI22_X1 u2_u10_u2_U43 (.ZN( u2_u10_u2_n135 ) , .B1( u2_u10_u2_n140 ) , .A1( u2_u10_u2_n156 ) , .B2( u2_u10_u2_n180 ) , .A2( u2_u10_u2_n188 ) );
  AOI21_X1 u2_u10_u2_U44 (.ZN( u2_u10_u2_n149 ) , .B1( u2_u10_u2_n173 ) , .B2( u2_u10_u2_n188 ) , .A( u2_u10_u2_n95 ) );
  AND3_X1 u2_u10_u2_U45 (.A2( u2_u10_u2_n100 ) , .A1( u2_u10_u2_n104 ) , .A3( u2_u10_u2_n156 ) , .ZN( u2_u10_u2_n95 ) );
  OAI21_X1 u2_u10_u2_U46 (.A( u2_u10_u2_n141 ) , .B2( u2_u10_u2_n142 ) , .ZN( u2_u10_u2_n146 ) , .B1( u2_u10_u2_n153 ) );
  OAI21_X1 u2_u10_u2_U47 (.A( u2_u10_u2_n140 ) , .ZN( u2_u10_u2_n141 ) , .B1( u2_u10_u2_n176 ) , .B2( u2_u10_u2_n177 ) );
  NOR3_X1 u2_u10_u2_U48 (.ZN( u2_u10_u2_n142 ) , .A3( u2_u10_u2_n175 ) , .A2( u2_u10_u2_n178 ) , .A1( u2_u10_u2_n181 ) );
  OAI21_X1 u2_u10_u2_U49 (.A( u2_u10_u2_n101 ) , .B2( u2_u10_u2_n121 ) , .B1( u2_u10_u2_n153 ) , .ZN( u2_u10_u2_n164 ) );
  INV_X1 u2_u10_u2_U5 (.A( u2_u10_u2_n150 ) , .ZN( u2_u10_u2_n184 ) );
  NAND2_X1 u2_u10_u2_U50 (.A2( u2_u10_u2_n100 ) , .A1( u2_u10_u2_n107 ) , .ZN( u2_u10_u2_n155 ) );
  NAND2_X1 u2_u10_u2_U51 (.A2( u2_u10_u2_n105 ) , .A1( u2_u10_u2_n108 ) , .ZN( u2_u10_u2_n143 ) );
  NAND2_X1 u2_u10_u2_U52 (.A1( u2_u10_u2_n104 ) , .A2( u2_u10_u2_n106 ) , .ZN( u2_u10_u2_n152 ) );
  NAND2_X1 u2_u10_u2_U53 (.A1( u2_u10_u2_n100 ) , .A2( u2_u10_u2_n105 ) , .ZN( u2_u10_u2_n132 ) );
  INV_X1 u2_u10_u2_U54 (.A( u2_u10_u2_n140 ) , .ZN( u2_u10_u2_n168 ) );
  INV_X1 u2_u10_u2_U55 (.A( u2_u10_u2_n138 ) , .ZN( u2_u10_u2_n167 ) );
  NAND2_X1 u2_u10_u2_U56 (.A1( u2_u10_u2_n102 ) , .A2( u2_u10_u2_n106 ) , .ZN( u2_u10_u2_n113 ) );
  NAND2_X1 u2_u10_u2_U57 (.A1( u2_u10_u2_n106 ) , .A2( u2_u10_u2_n107 ) , .ZN( u2_u10_u2_n131 ) );
  NAND2_X1 u2_u10_u2_U58 (.A1( u2_u10_u2_n103 ) , .A2( u2_u10_u2_n107 ) , .ZN( u2_u10_u2_n139 ) );
  NAND2_X1 u2_u10_u2_U59 (.A1( u2_u10_u2_n103 ) , .A2( u2_u10_u2_n105 ) , .ZN( u2_u10_u2_n133 ) );
  NOR4_X1 u2_u10_u2_U6 (.A4( u2_u10_u2_n124 ) , .A3( u2_u10_u2_n125 ) , .A2( u2_u10_u2_n126 ) , .A1( u2_u10_u2_n127 ) , .ZN( u2_u10_u2_n128 ) );
  NAND2_X1 u2_u10_u2_U60 (.A1( u2_u10_u2_n102 ) , .A2( u2_u10_u2_n103 ) , .ZN( u2_u10_u2_n154 ) );
  NAND2_X1 u2_u10_u2_U61 (.A2( u2_u10_u2_n103 ) , .A1( u2_u10_u2_n104 ) , .ZN( u2_u10_u2_n119 ) );
  NAND2_X1 u2_u10_u2_U62 (.A2( u2_u10_u2_n107 ) , .A1( u2_u10_u2_n108 ) , .ZN( u2_u10_u2_n123 ) );
  NAND2_X1 u2_u10_u2_U63 (.A1( u2_u10_u2_n104 ) , .A2( u2_u10_u2_n108 ) , .ZN( u2_u10_u2_n122 ) );
  INV_X1 u2_u10_u2_U64 (.A( u2_u10_u2_n114 ) , .ZN( u2_u10_u2_n172 ) );
  NAND2_X1 u2_u10_u2_U65 (.A2( u2_u10_u2_n100 ) , .A1( u2_u10_u2_n102 ) , .ZN( u2_u10_u2_n116 ) );
  NAND2_X1 u2_u10_u2_U66 (.A1( u2_u10_u2_n102 ) , .A2( u2_u10_u2_n108 ) , .ZN( u2_u10_u2_n120 ) );
  NAND2_X1 u2_u10_u2_U67 (.A2( u2_u10_u2_n105 ) , .A1( u2_u10_u2_n106 ) , .ZN( u2_u10_u2_n117 ) );
  INV_X1 u2_u10_u2_U68 (.ZN( u2_u10_u2_n187 ) , .A( u2_u10_u2_n99 ) );
  OAI21_X1 u2_u10_u2_U69 (.B1( u2_u10_u2_n137 ) , .B2( u2_u10_u2_n143 ) , .A( u2_u10_u2_n98 ) , .ZN( u2_u10_u2_n99 ) );
  AOI21_X1 u2_u10_u2_U7 (.ZN( u2_u10_u2_n124 ) , .B1( u2_u10_u2_n131 ) , .B2( u2_u10_u2_n143 ) , .A( u2_u10_u2_n172 ) );
  NOR2_X1 u2_u10_u2_U70 (.A2( u2_u10_X_16 ) , .ZN( u2_u10_u2_n140 ) , .A1( u2_u10_u2_n166 ) );
  NOR2_X1 u2_u10_u2_U71 (.A2( u2_u10_X_13 ) , .A1( u2_u10_X_14 ) , .ZN( u2_u10_u2_n100 ) );
  NOR2_X1 u2_u10_u2_U72 (.A2( u2_u10_X_16 ) , .A1( u2_u10_X_17 ) , .ZN( u2_u10_u2_n138 ) );
  NOR2_X1 u2_u10_u2_U73 (.A2( u2_u10_X_15 ) , .A1( u2_u10_X_18 ) , .ZN( u2_u10_u2_n104 ) );
  NOR2_X1 u2_u10_u2_U74 (.A2( u2_u10_X_14 ) , .ZN( u2_u10_u2_n103 ) , .A1( u2_u10_u2_n174 ) );
  NOR2_X1 u2_u10_u2_U75 (.A2( u2_u10_X_15 ) , .ZN( u2_u10_u2_n102 ) , .A1( u2_u10_u2_n165 ) );
  NOR2_X1 u2_u10_u2_U76 (.A2( u2_u10_X_17 ) , .ZN( u2_u10_u2_n114 ) , .A1( u2_u10_u2_n169 ) );
  AND2_X1 u2_u10_u2_U77 (.A1( u2_u10_X_15 ) , .ZN( u2_u10_u2_n105 ) , .A2( u2_u10_u2_n165 ) );
  AND2_X1 u2_u10_u2_U78 (.A2( u2_u10_X_15 ) , .A1( u2_u10_X_18 ) , .ZN( u2_u10_u2_n107 ) );
  AND2_X1 u2_u10_u2_U79 (.A1( u2_u10_X_14 ) , .ZN( u2_u10_u2_n106 ) , .A2( u2_u10_u2_n174 ) );
  AOI21_X1 u2_u10_u2_U8 (.B2( u2_u10_u2_n119 ) , .ZN( u2_u10_u2_n127 ) , .A( u2_u10_u2_n137 ) , .B1( u2_u10_u2_n155 ) );
  AND2_X1 u2_u10_u2_U80 (.A1( u2_u10_X_13 ) , .A2( u2_u10_X_14 ) , .ZN( u2_u10_u2_n108 ) );
  INV_X1 u2_u10_u2_U81 (.A( u2_u10_X_16 ) , .ZN( u2_u10_u2_n169 ) );
  INV_X1 u2_u10_u2_U82 (.A( u2_u10_X_17 ) , .ZN( u2_u10_u2_n166 ) );
  INV_X1 u2_u10_u2_U83 (.A( u2_u10_X_13 ) , .ZN( u2_u10_u2_n174 ) );
  INV_X1 u2_u10_u2_U84 (.A( u2_u10_X_18 ) , .ZN( u2_u10_u2_n165 ) );
  NAND4_X1 u2_u10_u2_U85 (.ZN( u2_out10_24 ) , .A4( u2_u10_u2_n111 ) , .A3( u2_u10_u2_n112 ) , .A1( u2_u10_u2_n130 ) , .A2( u2_u10_u2_n187 ) );
  AOI221_X1 u2_u10_u2_U86 (.A( u2_u10_u2_n109 ) , .B1( u2_u10_u2_n110 ) , .ZN( u2_u10_u2_n111 ) , .C1( u2_u10_u2_n134 ) , .C2( u2_u10_u2_n170 ) , .B2( u2_u10_u2_n173 ) );
  AOI21_X1 u2_u10_u2_U87 (.ZN( u2_u10_u2_n112 ) , .B2( u2_u10_u2_n156 ) , .A( u2_u10_u2_n164 ) , .B1( u2_u10_u2_n181 ) );
  NAND4_X1 u2_u10_u2_U88 (.ZN( u2_out10_16 ) , .A4( u2_u10_u2_n128 ) , .A3( u2_u10_u2_n129 ) , .A1( u2_u10_u2_n130 ) , .A2( u2_u10_u2_n186 ) );
  AOI22_X1 u2_u10_u2_U89 (.A2( u2_u10_u2_n118 ) , .ZN( u2_u10_u2_n129 ) , .A1( u2_u10_u2_n140 ) , .B1( u2_u10_u2_n157 ) , .B2( u2_u10_u2_n170 ) );
  AOI21_X1 u2_u10_u2_U9 (.B2( u2_u10_u2_n123 ) , .ZN( u2_u10_u2_n125 ) , .A( u2_u10_u2_n171 ) , .B1( u2_u10_u2_n184 ) );
  INV_X1 u2_u10_u2_U90 (.A( u2_u10_u2_n163 ) , .ZN( u2_u10_u2_n186 ) );
  NAND4_X1 u2_u10_u2_U91 (.ZN( u2_out10_30 ) , .A4( u2_u10_u2_n147 ) , .A3( u2_u10_u2_n148 ) , .A2( u2_u10_u2_n149 ) , .A1( u2_u10_u2_n187 ) );
  NOR3_X1 u2_u10_u2_U92 (.A3( u2_u10_u2_n144 ) , .A2( u2_u10_u2_n145 ) , .A1( u2_u10_u2_n146 ) , .ZN( u2_u10_u2_n147 ) );
  AOI21_X1 u2_u10_u2_U93 (.B2( u2_u10_u2_n138 ) , .ZN( u2_u10_u2_n148 ) , .A( u2_u10_u2_n162 ) , .B1( u2_u10_u2_n182 ) );
  OR4_X1 u2_u10_u2_U94 (.ZN( u2_out10_6 ) , .A4( u2_u10_u2_n161 ) , .A3( u2_u10_u2_n162 ) , .A2( u2_u10_u2_n163 ) , .A1( u2_u10_u2_n164 ) );
  OR3_X1 u2_u10_u2_U95 (.A2( u2_u10_u2_n159 ) , .A1( u2_u10_u2_n160 ) , .ZN( u2_u10_u2_n161 ) , .A3( u2_u10_u2_n183 ) );
  AOI21_X1 u2_u10_u2_U96 (.B2( u2_u10_u2_n154 ) , .B1( u2_u10_u2_n155 ) , .ZN( u2_u10_u2_n159 ) , .A( u2_u10_u2_n167 ) );
  NAND3_X1 u2_u10_u2_U97 (.A2( u2_u10_u2_n117 ) , .A1( u2_u10_u2_n122 ) , .A3( u2_u10_u2_n123 ) , .ZN( u2_u10_u2_n134 ) );
  NAND3_X1 u2_u10_u2_U98 (.ZN( u2_u10_u2_n110 ) , .A2( u2_u10_u2_n131 ) , .A3( u2_u10_u2_n139 ) , .A1( u2_u10_u2_n154 ) );
  NAND3_X1 u2_u10_u2_U99 (.A2( u2_u10_u2_n100 ) , .ZN( u2_u10_u2_n101 ) , .A1( u2_u10_u2_n104 ) , .A3( u2_u10_u2_n114 ) );
  OAI22_X1 u2_u10_u3_U10 (.B1( u2_u10_u3_n113 ) , .A2( u2_u10_u3_n135 ) , .A1( u2_u10_u3_n150 ) , .B2( u2_u10_u3_n164 ) , .ZN( u2_u10_u3_n98 ) );
  OAI211_X1 u2_u10_u3_U11 (.B( u2_u10_u3_n106 ) , .ZN( u2_u10_u3_n119 ) , .C2( u2_u10_u3_n128 ) , .C1( u2_u10_u3_n167 ) , .A( u2_u10_u3_n181 ) );
  AOI221_X1 u2_u10_u3_U12 (.C1( u2_u10_u3_n105 ) , .ZN( u2_u10_u3_n106 ) , .A( u2_u10_u3_n131 ) , .B2( u2_u10_u3_n132 ) , .C2( u2_u10_u3_n133 ) , .B1( u2_u10_u3_n169 ) );
  INV_X1 u2_u10_u3_U13 (.ZN( u2_u10_u3_n181 ) , .A( u2_u10_u3_n98 ) );
  NAND2_X1 u2_u10_u3_U14 (.ZN( u2_u10_u3_n105 ) , .A2( u2_u10_u3_n130 ) , .A1( u2_u10_u3_n155 ) );
  AOI22_X1 u2_u10_u3_U15 (.B1( u2_u10_u3_n115 ) , .A2( u2_u10_u3_n116 ) , .ZN( u2_u10_u3_n123 ) , .B2( u2_u10_u3_n133 ) , .A1( u2_u10_u3_n169 ) );
  NAND2_X1 u2_u10_u3_U16 (.ZN( u2_u10_u3_n116 ) , .A2( u2_u10_u3_n151 ) , .A1( u2_u10_u3_n182 ) );
  NOR2_X1 u2_u10_u3_U17 (.ZN( u2_u10_u3_n126 ) , .A2( u2_u10_u3_n150 ) , .A1( u2_u10_u3_n164 ) );
  AOI21_X1 u2_u10_u3_U18 (.ZN( u2_u10_u3_n112 ) , .B2( u2_u10_u3_n146 ) , .B1( u2_u10_u3_n155 ) , .A( u2_u10_u3_n167 ) );
  NAND2_X1 u2_u10_u3_U19 (.A1( u2_u10_u3_n135 ) , .ZN( u2_u10_u3_n142 ) , .A2( u2_u10_u3_n164 ) );
  NAND2_X1 u2_u10_u3_U20 (.ZN( u2_u10_u3_n132 ) , .A2( u2_u10_u3_n152 ) , .A1( u2_u10_u3_n156 ) );
  AND2_X1 u2_u10_u3_U21 (.A2( u2_u10_u3_n113 ) , .A1( u2_u10_u3_n114 ) , .ZN( u2_u10_u3_n151 ) );
  INV_X1 u2_u10_u3_U22 (.A( u2_u10_u3_n133 ) , .ZN( u2_u10_u3_n165 ) );
  INV_X1 u2_u10_u3_U23 (.A( u2_u10_u3_n135 ) , .ZN( u2_u10_u3_n170 ) );
  NAND2_X1 u2_u10_u3_U24 (.A1( u2_u10_u3_n107 ) , .A2( u2_u10_u3_n108 ) , .ZN( u2_u10_u3_n140 ) );
  NAND2_X1 u2_u10_u3_U25 (.ZN( u2_u10_u3_n117 ) , .A1( u2_u10_u3_n124 ) , .A2( u2_u10_u3_n148 ) );
  NAND2_X1 u2_u10_u3_U26 (.ZN( u2_u10_u3_n143 ) , .A1( u2_u10_u3_n165 ) , .A2( u2_u10_u3_n167 ) );
  INV_X1 u2_u10_u3_U27 (.A( u2_u10_u3_n130 ) , .ZN( u2_u10_u3_n177 ) );
  INV_X1 u2_u10_u3_U28 (.A( u2_u10_u3_n128 ) , .ZN( u2_u10_u3_n176 ) );
  INV_X1 u2_u10_u3_U29 (.A( u2_u10_u3_n155 ) , .ZN( u2_u10_u3_n174 ) );
  INV_X1 u2_u10_u3_U3 (.A( u2_u10_u3_n129 ) , .ZN( u2_u10_u3_n183 ) );
  INV_X1 u2_u10_u3_U30 (.A( u2_u10_u3_n139 ) , .ZN( u2_u10_u3_n185 ) );
  NOR2_X1 u2_u10_u3_U31 (.ZN( u2_u10_u3_n135 ) , .A2( u2_u10_u3_n141 ) , .A1( u2_u10_u3_n169 ) );
  OAI222_X1 u2_u10_u3_U32 (.C2( u2_u10_u3_n107 ) , .A2( u2_u10_u3_n108 ) , .B1( u2_u10_u3_n135 ) , .ZN( u2_u10_u3_n138 ) , .B2( u2_u10_u3_n146 ) , .C1( u2_u10_u3_n154 ) , .A1( u2_u10_u3_n164 ) );
  NOR4_X1 u2_u10_u3_U33 (.A4( u2_u10_u3_n157 ) , .A3( u2_u10_u3_n158 ) , .A2( u2_u10_u3_n159 ) , .A1( u2_u10_u3_n160 ) , .ZN( u2_u10_u3_n161 ) );
  AOI21_X1 u2_u10_u3_U34 (.B2( u2_u10_u3_n152 ) , .B1( u2_u10_u3_n153 ) , .ZN( u2_u10_u3_n158 ) , .A( u2_u10_u3_n164 ) );
  AOI21_X1 u2_u10_u3_U35 (.A( u2_u10_u3_n154 ) , .B2( u2_u10_u3_n155 ) , .B1( u2_u10_u3_n156 ) , .ZN( u2_u10_u3_n157 ) );
  AOI21_X1 u2_u10_u3_U36 (.A( u2_u10_u3_n149 ) , .B2( u2_u10_u3_n150 ) , .B1( u2_u10_u3_n151 ) , .ZN( u2_u10_u3_n159 ) );
  AOI211_X1 u2_u10_u3_U37 (.ZN( u2_u10_u3_n109 ) , .A( u2_u10_u3_n119 ) , .C2( u2_u10_u3_n129 ) , .B( u2_u10_u3_n138 ) , .C1( u2_u10_u3_n141 ) );
  AOI211_X1 u2_u10_u3_U38 (.B( u2_u10_u3_n119 ) , .A( u2_u10_u3_n120 ) , .C2( u2_u10_u3_n121 ) , .ZN( u2_u10_u3_n122 ) , .C1( u2_u10_u3_n179 ) );
  INV_X1 u2_u10_u3_U39 (.A( u2_u10_u3_n156 ) , .ZN( u2_u10_u3_n179 ) );
  INV_X1 u2_u10_u3_U4 (.A( u2_u10_u3_n140 ) , .ZN( u2_u10_u3_n182 ) );
  OAI22_X1 u2_u10_u3_U40 (.B1( u2_u10_u3_n118 ) , .ZN( u2_u10_u3_n120 ) , .A1( u2_u10_u3_n135 ) , .B2( u2_u10_u3_n154 ) , .A2( u2_u10_u3_n178 ) );
  AND3_X1 u2_u10_u3_U41 (.ZN( u2_u10_u3_n118 ) , .A2( u2_u10_u3_n124 ) , .A1( u2_u10_u3_n144 ) , .A3( u2_u10_u3_n152 ) );
  INV_X1 u2_u10_u3_U42 (.A( u2_u10_u3_n121 ) , .ZN( u2_u10_u3_n164 ) );
  NAND2_X1 u2_u10_u3_U43 (.ZN( u2_u10_u3_n133 ) , .A1( u2_u10_u3_n154 ) , .A2( u2_u10_u3_n164 ) );
  OAI211_X1 u2_u10_u3_U44 (.B( u2_u10_u3_n127 ) , .ZN( u2_u10_u3_n139 ) , .C1( u2_u10_u3_n150 ) , .C2( u2_u10_u3_n154 ) , .A( u2_u10_u3_n184 ) );
  INV_X1 u2_u10_u3_U45 (.A( u2_u10_u3_n125 ) , .ZN( u2_u10_u3_n184 ) );
  AOI221_X1 u2_u10_u3_U46 (.A( u2_u10_u3_n126 ) , .ZN( u2_u10_u3_n127 ) , .C2( u2_u10_u3_n132 ) , .C1( u2_u10_u3_n169 ) , .B2( u2_u10_u3_n170 ) , .B1( u2_u10_u3_n174 ) );
  OAI22_X1 u2_u10_u3_U47 (.A1( u2_u10_u3_n124 ) , .ZN( u2_u10_u3_n125 ) , .B2( u2_u10_u3_n145 ) , .A2( u2_u10_u3_n165 ) , .B1( u2_u10_u3_n167 ) );
  NOR2_X1 u2_u10_u3_U48 (.A1( u2_u10_u3_n113 ) , .ZN( u2_u10_u3_n131 ) , .A2( u2_u10_u3_n154 ) );
  NAND2_X1 u2_u10_u3_U49 (.A1( u2_u10_u3_n103 ) , .ZN( u2_u10_u3_n150 ) , .A2( u2_u10_u3_n99 ) );
  INV_X1 u2_u10_u3_U5 (.A( u2_u10_u3_n117 ) , .ZN( u2_u10_u3_n178 ) );
  NAND2_X1 u2_u10_u3_U50 (.A2( u2_u10_u3_n102 ) , .ZN( u2_u10_u3_n155 ) , .A1( u2_u10_u3_n97 ) );
  INV_X1 u2_u10_u3_U51 (.A( u2_u10_u3_n141 ) , .ZN( u2_u10_u3_n167 ) );
  AOI21_X1 u2_u10_u3_U52 (.B2( u2_u10_u3_n114 ) , .B1( u2_u10_u3_n146 ) , .A( u2_u10_u3_n154 ) , .ZN( u2_u10_u3_n94 ) );
  AOI21_X1 u2_u10_u3_U53 (.ZN( u2_u10_u3_n110 ) , .B2( u2_u10_u3_n142 ) , .B1( u2_u10_u3_n186 ) , .A( u2_u10_u3_n95 ) );
  INV_X1 u2_u10_u3_U54 (.A( u2_u10_u3_n145 ) , .ZN( u2_u10_u3_n186 ) );
  AOI21_X1 u2_u10_u3_U55 (.B1( u2_u10_u3_n124 ) , .A( u2_u10_u3_n149 ) , .B2( u2_u10_u3_n155 ) , .ZN( u2_u10_u3_n95 ) );
  INV_X1 u2_u10_u3_U56 (.A( u2_u10_u3_n149 ) , .ZN( u2_u10_u3_n169 ) );
  NAND2_X1 u2_u10_u3_U57 (.ZN( u2_u10_u3_n124 ) , .A1( u2_u10_u3_n96 ) , .A2( u2_u10_u3_n97 ) );
  NAND2_X1 u2_u10_u3_U58 (.A2( u2_u10_u3_n100 ) , .ZN( u2_u10_u3_n146 ) , .A1( u2_u10_u3_n96 ) );
  NAND2_X1 u2_u10_u3_U59 (.A1( u2_u10_u3_n101 ) , .ZN( u2_u10_u3_n145 ) , .A2( u2_u10_u3_n99 ) );
  AOI221_X1 u2_u10_u3_U6 (.A( u2_u10_u3_n131 ) , .C2( u2_u10_u3_n132 ) , .C1( u2_u10_u3_n133 ) , .ZN( u2_u10_u3_n134 ) , .B1( u2_u10_u3_n143 ) , .B2( u2_u10_u3_n177 ) );
  NAND2_X1 u2_u10_u3_U60 (.A1( u2_u10_u3_n100 ) , .ZN( u2_u10_u3_n156 ) , .A2( u2_u10_u3_n99 ) );
  NAND2_X1 u2_u10_u3_U61 (.A2( u2_u10_u3_n101 ) , .A1( u2_u10_u3_n104 ) , .ZN( u2_u10_u3_n148 ) );
  NAND2_X1 u2_u10_u3_U62 (.A1( u2_u10_u3_n100 ) , .A2( u2_u10_u3_n102 ) , .ZN( u2_u10_u3_n128 ) );
  NAND2_X1 u2_u10_u3_U63 (.A2( u2_u10_u3_n101 ) , .A1( u2_u10_u3_n102 ) , .ZN( u2_u10_u3_n152 ) );
  NAND2_X1 u2_u10_u3_U64 (.A2( u2_u10_u3_n101 ) , .ZN( u2_u10_u3_n114 ) , .A1( u2_u10_u3_n96 ) );
  NAND2_X1 u2_u10_u3_U65 (.ZN( u2_u10_u3_n107 ) , .A1( u2_u10_u3_n97 ) , .A2( u2_u10_u3_n99 ) );
  NAND2_X1 u2_u10_u3_U66 (.A2( u2_u10_u3_n100 ) , .A1( u2_u10_u3_n104 ) , .ZN( u2_u10_u3_n113 ) );
  NAND2_X1 u2_u10_u3_U67 (.A1( u2_u10_u3_n104 ) , .ZN( u2_u10_u3_n153 ) , .A2( u2_u10_u3_n97 ) );
  NAND2_X1 u2_u10_u3_U68 (.A2( u2_u10_u3_n103 ) , .A1( u2_u10_u3_n104 ) , .ZN( u2_u10_u3_n130 ) );
  NAND2_X1 u2_u10_u3_U69 (.A2( u2_u10_u3_n103 ) , .ZN( u2_u10_u3_n144 ) , .A1( u2_u10_u3_n96 ) );
  OAI22_X1 u2_u10_u3_U7 (.B2( u2_u10_u3_n147 ) , .A2( u2_u10_u3_n148 ) , .ZN( u2_u10_u3_n160 ) , .B1( u2_u10_u3_n165 ) , .A1( u2_u10_u3_n168 ) );
  NAND2_X1 u2_u10_u3_U70 (.A1( u2_u10_u3_n102 ) , .A2( u2_u10_u3_n103 ) , .ZN( u2_u10_u3_n108 ) );
  NOR2_X1 u2_u10_u3_U71 (.A2( u2_u10_X_19 ) , .A1( u2_u10_X_20 ) , .ZN( u2_u10_u3_n99 ) );
  NOR2_X1 u2_u10_u3_U72 (.A2( u2_u10_X_21 ) , .A1( u2_u10_X_24 ) , .ZN( u2_u10_u3_n103 ) );
  NOR2_X1 u2_u10_u3_U73 (.A2( u2_u10_X_24 ) , .A1( u2_u10_u3_n171 ) , .ZN( u2_u10_u3_n97 ) );
  NOR2_X1 u2_u10_u3_U74 (.A2( u2_u10_X_23 ) , .ZN( u2_u10_u3_n141 ) , .A1( u2_u10_u3_n166 ) );
  NOR2_X1 u2_u10_u3_U75 (.A2( u2_u10_X_19 ) , .A1( u2_u10_u3_n172 ) , .ZN( u2_u10_u3_n96 ) );
  NAND2_X1 u2_u10_u3_U76 (.A1( u2_u10_X_22 ) , .A2( u2_u10_X_23 ) , .ZN( u2_u10_u3_n154 ) );
  NAND2_X1 u2_u10_u3_U77 (.A1( u2_u10_X_23 ) , .ZN( u2_u10_u3_n149 ) , .A2( u2_u10_u3_n166 ) );
  NOR2_X1 u2_u10_u3_U78 (.A2( u2_u10_X_22 ) , .A1( u2_u10_X_23 ) , .ZN( u2_u10_u3_n121 ) );
  AND2_X1 u2_u10_u3_U79 (.A1( u2_u10_X_24 ) , .ZN( u2_u10_u3_n101 ) , .A2( u2_u10_u3_n171 ) );
  AND3_X1 u2_u10_u3_U8 (.A3( u2_u10_u3_n144 ) , .A2( u2_u10_u3_n145 ) , .A1( u2_u10_u3_n146 ) , .ZN( u2_u10_u3_n147 ) );
  AND2_X1 u2_u10_u3_U80 (.A1( u2_u10_X_19 ) , .ZN( u2_u10_u3_n102 ) , .A2( u2_u10_u3_n172 ) );
  AND2_X1 u2_u10_u3_U81 (.A1( u2_u10_X_21 ) , .A2( u2_u10_X_24 ) , .ZN( u2_u10_u3_n100 ) );
  AND2_X1 u2_u10_u3_U82 (.A2( u2_u10_X_19 ) , .A1( u2_u10_X_20 ) , .ZN( u2_u10_u3_n104 ) );
  INV_X1 u2_u10_u3_U83 (.A( u2_u10_X_22 ) , .ZN( u2_u10_u3_n166 ) );
  INV_X1 u2_u10_u3_U84 (.A( u2_u10_X_21 ) , .ZN( u2_u10_u3_n171 ) );
  INV_X1 u2_u10_u3_U85 (.A( u2_u10_X_20 ) , .ZN( u2_u10_u3_n172 ) );
  OR4_X1 u2_u10_u3_U86 (.ZN( u2_out10_10 ) , .A4( u2_u10_u3_n136 ) , .A3( u2_u10_u3_n137 ) , .A1( u2_u10_u3_n138 ) , .A2( u2_u10_u3_n139 ) );
  OAI222_X1 u2_u10_u3_U87 (.C1( u2_u10_u3_n128 ) , .ZN( u2_u10_u3_n137 ) , .B1( u2_u10_u3_n148 ) , .A2( u2_u10_u3_n150 ) , .B2( u2_u10_u3_n154 ) , .C2( u2_u10_u3_n164 ) , .A1( u2_u10_u3_n167 ) );
  OAI221_X1 u2_u10_u3_U88 (.A( u2_u10_u3_n134 ) , .B2( u2_u10_u3_n135 ) , .ZN( u2_u10_u3_n136 ) , .C1( u2_u10_u3_n149 ) , .B1( u2_u10_u3_n151 ) , .C2( u2_u10_u3_n183 ) );
  NAND4_X1 u2_u10_u3_U89 (.ZN( u2_out10_26 ) , .A4( u2_u10_u3_n109 ) , .A3( u2_u10_u3_n110 ) , .A2( u2_u10_u3_n111 ) , .A1( u2_u10_u3_n173 ) );
  INV_X1 u2_u10_u3_U9 (.A( u2_u10_u3_n143 ) , .ZN( u2_u10_u3_n168 ) );
  INV_X1 u2_u10_u3_U90 (.ZN( u2_u10_u3_n173 ) , .A( u2_u10_u3_n94 ) );
  OAI21_X1 u2_u10_u3_U91 (.ZN( u2_u10_u3_n111 ) , .B2( u2_u10_u3_n117 ) , .A( u2_u10_u3_n133 ) , .B1( u2_u10_u3_n176 ) );
  NAND4_X1 u2_u10_u3_U92 (.ZN( u2_out10_20 ) , .A4( u2_u10_u3_n122 ) , .A3( u2_u10_u3_n123 ) , .A1( u2_u10_u3_n175 ) , .A2( u2_u10_u3_n180 ) );
  INV_X1 u2_u10_u3_U93 (.A( u2_u10_u3_n126 ) , .ZN( u2_u10_u3_n180 ) );
  INV_X1 u2_u10_u3_U94 (.A( u2_u10_u3_n112 ) , .ZN( u2_u10_u3_n175 ) );
  NAND4_X1 u2_u10_u3_U95 (.ZN( u2_out10_1 ) , .A4( u2_u10_u3_n161 ) , .A3( u2_u10_u3_n162 ) , .A2( u2_u10_u3_n163 ) , .A1( u2_u10_u3_n185 ) );
  NAND2_X1 u2_u10_u3_U96 (.ZN( u2_u10_u3_n163 ) , .A2( u2_u10_u3_n170 ) , .A1( u2_u10_u3_n176 ) );
  AOI22_X1 u2_u10_u3_U97 (.B2( u2_u10_u3_n140 ) , .B1( u2_u10_u3_n141 ) , .A2( u2_u10_u3_n142 ) , .ZN( u2_u10_u3_n162 ) , .A1( u2_u10_u3_n177 ) );
  NAND3_X1 u2_u10_u3_U98 (.A1( u2_u10_u3_n114 ) , .ZN( u2_u10_u3_n115 ) , .A2( u2_u10_u3_n145 ) , .A3( u2_u10_u3_n153 ) );
  NAND3_X1 u2_u10_u3_U99 (.ZN( u2_u10_u3_n129 ) , .A2( u2_u10_u3_n144 ) , .A1( u2_u10_u3_n153 ) , .A3( u2_u10_u3_n182 ) );
  XOR2_X1 u2_u12_U20 (.B( u2_K13_36 ) , .A( u2_R11_25 ) , .Z( u2_u12_X_36 ) );
  XOR2_X1 u2_u12_U21 (.B( u2_K13_35 ) , .A( u2_R11_24 ) , .Z( u2_u12_X_35 ) );
  XOR2_X1 u2_u12_U22 (.B( u2_K13_34 ) , .A( u2_R11_23 ) , .Z( u2_u12_X_34 ) );
  XOR2_X1 u2_u12_U23 (.B( u2_K13_33 ) , .A( u2_R11_22 ) , .Z( u2_u12_X_33 ) );
  XOR2_X1 u2_u12_U24 (.B( u2_K13_32 ) , .A( u2_R11_21 ) , .Z( u2_u12_X_32 ) );
  XOR2_X1 u2_u12_U25 (.B( u2_K13_31 ) , .A( u2_R11_20 ) , .Z( u2_u12_X_31 ) );
  XOR2_X1 u2_u12_U26 (.B( u2_K13_30 ) , .A( u2_R11_21 ) , .Z( u2_u12_X_30 ) );
  XOR2_X1 u2_u12_U28 (.B( u2_K13_29 ) , .A( u2_R11_20 ) , .Z( u2_u12_X_29 ) );
  XOR2_X1 u2_u12_U29 (.B( u2_K13_28 ) , .A( u2_R11_19 ) , .Z( u2_u12_X_28 ) );
  XOR2_X1 u2_u12_U30 (.B( u2_K13_27 ) , .A( u2_R11_18 ) , .Z( u2_u12_X_27 ) );
  XOR2_X1 u2_u12_U31 (.B( u2_K13_26 ) , .A( u2_R11_17 ) , .Z( u2_u12_X_26 ) );
  XOR2_X1 u2_u12_U32 (.B( u2_K13_25 ) , .A( u2_R11_16 ) , .Z( u2_u12_X_25 ) );
  XOR2_X1 u2_u12_U33 (.B( u2_K13_24 ) , .A( u2_R11_17 ) , .Z( u2_u12_X_24 ) );
  XOR2_X1 u2_u12_U34 (.B( u2_K13_23 ) , .A( u2_R11_16 ) , .Z( u2_u12_X_23 ) );
  XOR2_X1 u2_u12_U35 (.B( u2_K13_22 ) , .A( u2_R11_15 ) , .Z( u2_u12_X_22 ) );
  XOR2_X1 u2_u12_U36 (.B( u2_K13_21 ) , .A( u2_R11_14 ) , .Z( u2_u12_X_21 ) );
  XOR2_X1 u2_u12_U37 (.B( u2_K13_20 ) , .A( u2_R11_13 ) , .Z( u2_u12_X_20 ) );
  XOR2_X1 u2_u12_U39 (.B( u2_K13_19 ) , .A( u2_R11_12 ) , .Z( u2_u12_X_19 ) );
  OAI22_X1 u2_u12_u3_U10 (.B1( u2_u12_u3_n113 ) , .A2( u2_u12_u3_n135 ) , .A1( u2_u12_u3_n150 ) , .B2( u2_u12_u3_n164 ) , .ZN( u2_u12_u3_n98 ) );
  OAI211_X1 u2_u12_u3_U11 (.B( u2_u12_u3_n106 ) , .ZN( u2_u12_u3_n119 ) , .C2( u2_u12_u3_n128 ) , .C1( u2_u12_u3_n167 ) , .A( u2_u12_u3_n181 ) );
  AOI221_X1 u2_u12_u3_U12 (.C1( u2_u12_u3_n105 ) , .ZN( u2_u12_u3_n106 ) , .A( u2_u12_u3_n131 ) , .B2( u2_u12_u3_n132 ) , .C2( u2_u12_u3_n133 ) , .B1( u2_u12_u3_n169 ) );
  INV_X1 u2_u12_u3_U13 (.ZN( u2_u12_u3_n181 ) , .A( u2_u12_u3_n98 ) );
  NAND2_X1 u2_u12_u3_U14 (.ZN( u2_u12_u3_n105 ) , .A2( u2_u12_u3_n130 ) , .A1( u2_u12_u3_n155 ) );
  AOI22_X1 u2_u12_u3_U15 (.B1( u2_u12_u3_n115 ) , .A2( u2_u12_u3_n116 ) , .ZN( u2_u12_u3_n123 ) , .B2( u2_u12_u3_n133 ) , .A1( u2_u12_u3_n169 ) );
  NAND2_X1 u2_u12_u3_U16 (.ZN( u2_u12_u3_n116 ) , .A2( u2_u12_u3_n151 ) , .A1( u2_u12_u3_n182 ) );
  NOR2_X1 u2_u12_u3_U17 (.ZN( u2_u12_u3_n126 ) , .A2( u2_u12_u3_n150 ) , .A1( u2_u12_u3_n164 ) );
  AOI21_X1 u2_u12_u3_U18 (.ZN( u2_u12_u3_n112 ) , .B2( u2_u12_u3_n146 ) , .B1( u2_u12_u3_n155 ) , .A( u2_u12_u3_n167 ) );
  NAND2_X1 u2_u12_u3_U19 (.A1( u2_u12_u3_n135 ) , .ZN( u2_u12_u3_n142 ) , .A2( u2_u12_u3_n164 ) );
  NAND2_X1 u2_u12_u3_U20 (.ZN( u2_u12_u3_n132 ) , .A2( u2_u12_u3_n152 ) , .A1( u2_u12_u3_n156 ) );
  AND2_X1 u2_u12_u3_U21 (.A2( u2_u12_u3_n113 ) , .A1( u2_u12_u3_n114 ) , .ZN( u2_u12_u3_n151 ) );
  INV_X1 u2_u12_u3_U22 (.A( u2_u12_u3_n133 ) , .ZN( u2_u12_u3_n165 ) );
  INV_X1 u2_u12_u3_U23 (.A( u2_u12_u3_n135 ) , .ZN( u2_u12_u3_n170 ) );
  NAND2_X1 u2_u12_u3_U24 (.A1( u2_u12_u3_n107 ) , .A2( u2_u12_u3_n108 ) , .ZN( u2_u12_u3_n140 ) );
  NAND2_X1 u2_u12_u3_U25 (.ZN( u2_u12_u3_n117 ) , .A1( u2_u12_u3_n124 ) , .A2( u2_u12_u3_n148 ) );
  NAND2_X1 u2_u12_u3_U26 (.ZN( u2_u12_u3_n143 ) , .A1( u2_u12_u3_n165 ) , .A2( u2_u12_u3_n167 ) );
  INV_X1 u2_u12_u3_U27 (.A( u2_u12_u3_n130 ) , .ZN( u2_u12_u3_n177 ) );
  INV_X1 u2_u12_u3_U28 (.A( u2_u12_u3_n128 ) , .ZN( u2_u12_u3_n176 ) );
  INV_X1 u2_u12_u3_U29 (.A( u2_u12_u3_n155 ) , .ZN( u2_u12_u3_n174 ) );
  INV_X1 u2_u12_u3_U3 (.A( u2_u12_u3_n129 ) , .ZN( u2_u12_u3_n183 ) );
  INV_X1 u2_u12_u3_U30 (.A( u2_u12_u3_n139 ) , .ZN( u2_u12_u3_n185 ) );
  NOR2_X1 u2_u12_u3_U31 (.ZN( u2_u12_u3_n135 ) , .A2( u2_u12_u3_n141 ) , .A1( u2_u12_u3_n169 ) );
  OAI222_X1 u2_u12_u3_U32 (.C2( u2_u12_u3_n107 ) , .A2( u2_u12_u3_n108 ) , .B1( u2_u12_u3_n135 ) , .ZN( u2_u12_u3_n138 ) , .B2( u2_u12_u3_n146 ) , .C1( u2_u12_u3_n154 ) , .A1( u2_u12_u3_n164 ) );
  NOR4_X1 u2_u12_u3_U33 (.A4( u2_u12_u3_n157 ) , .A3( u2_u12_u3_n158 ) , .A2( u2_u12_u3_n159 ) , .A1( u2_u12_u3_n160 ) , .ZN( u2_u12_u3_n161 ) );
  AOI21_X1 u2_u12_u3_U34 (.B2( u2_u12_u3_n152 ) , .B1( u2_u12_u3_n153 ) , .ZN( u2_u12_u3_n158 ) , .A( u2_u12_u3_n164 ) );
  AOI21_X1 u2_u12_u3_U35 (.A( u2_u12_u3_n154 ) , .B2( u2_u12_u3_n155 ) , .B1( u2_u12_u3_n156 ) , .ZN( u2_u12_u3_n157 ) );
  AOI21_X1 u2_u12_u3_U36 (.A( u2_u12_u3_n149 ) , .B2( u2_u12_u3_n150 ) , .B1( u2_u12_u3_n151 ) , .ZN( u2_u12_u3_n159 ) );
  AOI211_X1 u2_u12_u3_U37 (.ZN( u2_u12_u3_n109 ) , .A( u2_u12_u3_n119 ) , .C2( u2_u12_u3_n129 ) , .B( u2_u12_u3_n138 ) , .C1( u2_u12_u3_n141 ) );
  AOI211_X1 u2_u12_u3_U38 (.B( u2_u12_u3_n119 ) , .A( u2_u12_u3_n120 ) , .C2( u2_u12_u3_n121 ) , .ZN( u2_u12_u3_n122 ) , .C1( u2_u12_u3_n179 ) );
  INV_X1 u2_u12_u3_U39 (.A( u2_u12_u3_n156 ) , .ZN( u2_u12_u3_n179 ) );
  INV_X1 u2_u12_u3_U4 (.A( u2_u12_u3_n140 ) , .ZN( u2_u12_u3_n182 ) );
  OAI22_X1 u2_u12_u3_U40 (.B1( u2_u12_u3_n118 ) , .ZN( u2_u12_u3_n120 ) , .A1( u2_u12_u3_n135 ) , .B2( u2_u12_u3_n154 ) , .A2( u2_u12_u3_n178 ) );
  AND3_X1 u2_u12_u3_U41 (.ZN( u2_u12_u3_n118 ) , .A2( u2_u12_u3_n124 ) , .A1( u2_u12_u3_n144 ) , .A3( u2_u12_u3_n152 ) );
  INV_X1 u2_u12_u3_U42 (.A( u2_u12_u3_n121 ) , .ZN( u2_u12_u3_n164 ) );
  NAND2_X1 u2_u12_u3_U43 (.ZN( u2_u12_u3_n133 ) , .A1( u2_u12_u3_n154 ) , .A2( u2_u12_u3_n164 ) );
  OAI211_X1 u2_u12_u3_U44 (.B( u2_u12_u3_n127 ) , .ZN( u2_u12_u3_n139 ) , .C1( u2_u12_u3_n150 ) , .C2( u2_u12_u3_n154 ) , .A( u2_u12_u3_n184 ) );
  INV_X1 u2_u12_u3_U45 (.A( u2_u12_u3_n125 ) , .ZN( u2_u12_u3_n184 ) );
  AOI221_X1 u2_u12_u3_U46 (.A( u2_u12_u3_n126 ) , .ZN( u2_u12_u3_n127 ) , .C2( u2_u12_u3_n132 ) , .C1( u2_u12_u3_n169 ) , .B2( u2_u12_u3_n170 ) , .B1( u2_u12_u3_n174 ) );
  OAI22_X1 u2_u12_u3_U47 (.A1( u2_u12_u3_n124 ) , .ZN( u2_u12_u3_n125 ) , .B2( u2_u12_u3_n145 ) , .A2( u2_u12_u3_n165 ) , .B1( u2_u12_u3_n167 ) );
  NOR2_X1 u2_u12_u3_U48 (.A1( u2_u12_u3_n113 ) , .ZN( u2_u12_u3_n131 ) , .A2( u2_u12_u3_n154 ) );
  NAND2_X1 u2_u12_u3_U49 (.A1( u2_u12_u3_n103 ) , .ZN( u2_u12_u3_n150 ) , .A2( u2_u12_u3_n99 ) );
  INV_X1 u2_u12_u3_U5 (.A( u2_u12_u3_n117 ) , .ZN( u2_u12_u3_n178 ) );
  NAND2_X1 u2_u12_u3_U50 (.A2( u2_u12_u3_n102 ) , .ZN( u2_u12_u3_n155 ) , .A1( u2_u12_u3_n97 ) );
  INV_X1 u2_u12_u3_U51 (.A( u2_u12_u3_n141 ) , .ZN( u2_u12_u3_n167 ) );
  AOI21_X1 u2_u12_u3_U52 (.B2( u2_u12_u3_n114 ) , .B1( u2_u12_u3_n146 ) , .A( u2_u12_u3_n154 ) , .ZN( u2_u12_u3_n94 ) );
  AOI21_X1 u2_u12_u3_U53 (.ZN( u2_u12_u3_n110 ) , .B2( u2_u12_u3_n142 ) , .B1( u2_u12_u3_n186 ) , .A( u2_u12_u3_n95 ) );
  INV_X1 u2_u12_u3_U54 (.A( u2_u12_u3_n145 ) , .ZN( u2_u12_u3_n186 ) );
  AOI21_X1 u2_u12_u3_U55 (.B1( u2_u12_u3_n124 ) , .A( u2_u12_u3_n149 ) , .B2( u2_u12_u3_n155 ) , .ZN( u2_u12_u3_n95 ) );
  INV_X1 u2_u12_u3_U56 (.A( u2_u12_u3_n149 ) , .ZN( u2_u12_u3_n169 ) );
  NAND2_X1 u2_u12_u3_U57 (.ZN( u2_u12_u3_n124 ) , .A1( u2_u12_u3_n96 ) , .A2( u2_u12_u3_n97 ) );
  NAND2_X1 u2_u12_u3_U58 (.A2( u2_u12_u3_n100 ) , .ZN( u2_u12_u3_n146 ) , .A1( u2_u12_u3_n96 ) );
  NAND2_X1 u2_u12_u3_U59 (.A1( u2_u12_u3_n101 ) , .ZN( u2_u12_u3_n145 ) , .A2( u2_u12_u3_n99 ) );
  AOI221_X1 u2_u12_u3_U6 (.A( u2_u12_u3_n131 ) , .C2( u2_u12_u3_n132 ) , .C1( u2_u12_u3_n133 ) , .ZN( u2_u12_u3_n134 ) , .B1( u2_u12_u3_n143 ) , .B2( u2_u12_u3_n177 ) );
  NAND2_X1 u2_u12_u3_U60 (.A1( u2_u12_u3_n100 ) , .ZN( u2_u12_u3_n156 ) , .A2( u2_u12_u3_n99 ) );
  NAND2_X1 u2_u12_u3_U61 (.A2( u2_u12_u3_n101 ) , .A1( u2_u12_u3_n104 ) , .ZN( u2_u12_u3_n148 ) );
  NAND2_X1 u2_u12_u3_U62 (.A1( u2_u12_u3_n100 ) , .A2( u2_u12_u3_n102 ) , .ZN( u2_u12_u3_n128 ) );
  NAND2_X1 u2_u12_u3_U63 (.A2( u2_u12_u3_n101 ) , .A1( u2_u12_u3_n102 ) , .ZN( u2_u12_u3_n152 ) );
  NAND2_X1 u2_u12_u3_U64 (.A2( u2_u12_u3_n101 ) , .ZN( u2_u12_u3_n114 ) , .A1( u2_u12_u3_n96 ) );
  NAND2_X1 u2_u12_u3_U65 (.ZN( u2_u12_u3_n107 ) , .A1( u2_u12_u3_n97 ) , .A2( u2_u12_u3_n99 ) );
  NAND2_X1 u2_u12_u3_U66 (.A2( u2_u12_u3_n100 ) , .A1( u2_u12_u3_n104 ) , .ZN( u2_u12_u3_n113 ) );
  NAND2_X1 u2_u12_u3_U67 (.A1( u2_u12_u3_n104 ) , .ZN( u2_u12_u3_n153 ) , .A2( u2_u12_u3_n97 ) );
  NAND2_X1 u2_u12_u3_U68 (.A2( u2_u12_u3_n103 ) , .A1( u2_u12_u3_n104 ) , .ZN( u2_u12_u3_n130 ) );
  NAND2_X1 u2_u12_u3_U69 (.A2( u2_u12_u3_n103 ) , .ZN( u2_u12_u3_n144 ) , .A1( u2_u12_u3_n96 ) );
  OAI22_X1 u2_u12_u3_U7 (.B2( u2_u12_u3_n147 ) , .A2( u2_u12_u3_n148 ) , .ZN( u2_u12_u3_n160 ) , .B1( u2_u12_u3_n165 ) , .A1( u2_u12_u3_n168 ) );
  NAND2_X1 u2_u12_u3_U70 (.A1( u2_u12_u3_n102 ) , .A2( u2_u12_u3_n103 ) , .ZN( u2_u12_u3_n108 ) );
  NOR2_X1 u2_u12_u3_U71 (.A2( u2_u12_X_19 ) , .A1( u2_u12_X_20 ) , .ZN( u2_u12_u3_n99 ) );
  NOR2_X1 u2_u12_u3_U72 (.A2( u2_u12_X_21 ) , .A1( u2_u12_X_24 ) , .ZN( u2_u12_u3_n103 ) );
  NOR2_X1 u2_u12_u3_U73 (.A2( u2_u12_X_24 ) , .A1( u2_u12_u3_n171 ) , .ZN( u2_u12_u3_n97 ) );
  NOR2_X1 u2_u12_u3_U74 (.A2( u2_u12_X_23 ) , .ZN( u2_u12_u3_n141 ) , .A1( u2_u12_u3_n166 ) );
  NOR2_X1 u2_u12_u3_U75 (.A2( u2_u12_X_19 ) , .A1( u2_u12_u3_n172 ) , .ZN( u2_u12_u3_n96 ) );
  NAND2_X1 u2_u12_u3_U76 (.A1( u2_u12_X_22 ) , .A2( u2_u12_X_23 ) , .ZN( u2_u12_u3_n154 ) );
  NAND2_X1 u2_u12_u3_U77 (.A1( u2_u12_X_23 ) , .ZN( u2_u12_u3_n149 ) , .A2( u2_u12_u3_n166 ) );
  NOR2_X1 u2_u12_u3_U78 (.A2( u2_u12_X_22 ) , .A1( u2_u12_X_23 ) , .ZN( u2_u12_u3_n121 ) );
  AND2_X1 u2_u12_u3_U79 (.A1( u2_u12_X_24 ) , .ZN( u2_u12_u3_n101 ) , .A2( u2_u12_u3_n171 ) );
  AND3_X1 u2_u12_u3_U8 (.A3( u2_u12_u3_n144 ) , .A2( u2_u12_u3_n145 ) , .A1( u2_u12_u3_n146 ) , .ZN( u2_u12_u3_n147 ) );
  AND2_X1 u2_u12_u3_U80 (.A1( u2_u12_X_19 ) , .ZN( u2_u12_u3_n102 ) , .A2( u2_u12_u3_n172 ) );
  AND2_X1 u2_u12_u3_U81 (.A1( u2_u12_X_21 ) , .A2( u2_u12_X_24 ) , .ZN( u2_u12_u3_n100 ) );
  AND2_X1 u2_u12_u3_U82 (.A2( u2_u12_X_19 ) , .A1( u2_u12_X_20 ) , .ZN( u2_u12_u3_n104 ) );
  INV_X1 u2_u12_u3_U83 (.A( u2_u12_X_22 ) , .ZN( u2_u12_u3_n166 ) );
  INV_X1 u2_u12_u3_U84 (.A( u2_u12_X_21 ) , .ZN( u2_u12_u3_n171 ) );
  INV_X1 u2_u12_u3_U85 (.A( u2_u12_X_20 ) , .ZN( u2_u12_u3_n172 ) );
  OR4_X1 u2_u12_u3_U86 (.ZN( u2_out12_10 ) , .A4( u2_u12_u3_n136 ) , .A3( u2_u12_u3_n137 ) , .A1( u2_u12_u3_n138 ) , .A2( u2_u12_u3_n139 ) );
  OAI222_X1 u2_u12_u3_U87 (.C1( u2_u12_u3_n128 ) , .ZN( u2_u12_u3_n137 ) , .B1( u2_u12_u3_n148 ) , .A2( u2_u12_u3_n150 ) , .B2( u2_u12_u3_n154 ) , .C2( u2_u12_u3_n164 ) , .A1( u2_u12_u3_n167 ) );
  OAI221_X1 u2_u12_u3_U88 (.A( u2_u12_u3_n134 ) , .B2( u2_u12_u3_n135 ) , .ZN( u2_u12_u3_n136 ) , .C1( u2_u12_u3_n149 ) , .B1( u2_u12_u3_n151 ) , .C2( u2_u12_u3_n183 ) );
  NAND4_X1 u2_u12_u3_U89 (.ZN( u2_out12_26 ) , .A4( u2_u12_u3_n109 ) , .A3( u2_u12_u3_n110 ) , .A2( u2_u12_u3_n111 ) , .A1( u2_u12_u3_n173 ) );
  INV_X1 u2_u12_u3_U9 (.A( u2_u12_u3_n143 ) , .ZN( u2_u12_u3_n168 ) );
  INV_X1 u2_u12_u3_U90 (.ZN( u2_u12_u3_n173 ) , .A( u2_u12_u3_n94 ) );
  OAI21_X1 u2_u12_u3_U91 (.ZN( u2_u12_u3_n111 ) , .B2( u2_u12_u3_n117 ) , .A( u2_u12_u3_n133 ) , .B1( u2_u12_u3_n176 ) );
  NAND4_X1 u2_u12_u3_U92 (.ZN( u2_out12_20 ) , .A4( u2_u12_u3_n122 ) , .A3( u2_u12_u3_n123 ) , .A1( u2_u12_u3_n175 ) , .A2( u2_u12_u3_n180 ) );
  INV_X1 u2_u12_u3_U93 (.A( u2_u12_u3_n126 ) , .ZN( u2_u12_u3_n180 ) );
  INV_X1 u2_u12_u3_U94 (.A( u2_u12_u3_n112 ) , .ZN( u2_u12_u3_n175 ) );
  NAND4_X1 u2_u12_u3_U95 (.ZN( u2_out12_1 ) , .A4( u2_u12_u3_n161 ) , .A3( u2_u12_u3_n162 ) , .A2( u2_u12_u3_n163 ) , .A1( u2_u12_u3_n185 ) );
  NAND2_X1 u2_u12_u3_U96 (.ZN( u2_u12_u3_n163 ) , .A2( u2_u12_u3_n170 ) , .A1( u2_u12_u3_n176 ) );
  AOI22_X1 u2_u12_u3_U97 (.B2( u2_u12_u3_n140 ) , .B1( u2_u12_u3_n141 ) , .A2( u2_u12_u3_n142 ) , .ZN( u2_u12_u3_n162 ) , .A1( u2_u12_u3_n177 ) );
  NAND3_X1 u2_u12_u3_U98 (.A1( u2_u12_u3_n114 ) , .ZN( u2_u12_u3_n115 ) , .A2( u2_u12_u3_n145 ) , .A3( u2_u12_u3_n153 ) );
  NAND3_X1 u2_u12_u3_U99 (.ZN( u2_u12_u3_n129 ) , .A2( u2_u12_u3_n144 ) , .A1( u2_u12_u3_n153 ) , .A3( u2_u12_u3_n182 ) );
  OAI22_X1 u2_u12_u4_U10 (.B2( u2_u12_u4_n135 ) , .ZN( u2_u12_u4_n137 ) , .B1( u2_u12_u4_n153 ) , .A1( u2_u12_u4_n155 ) , .A2( u2_u12_u4_n171 ) );
  AND3_X1 u2_u12_u4_U11 (.A2( u2_u12_u4_n134 ) , .ZN( u2_u12_u4_n135 ) , .A3( u2_u12_u4_n145 ) , .A1( u2_u12_u4_n157 ) );
  NAND2_X1 u2_u12_u4_U12 (.ZN( u2_u12_u4_n132 ) , .A2( u2_u12_u4_n170 ) , .A1( u2_u12_u4_n173 ) );
  AOI21_X1 u2_u12_u4_U13 (.B2( u2_u12_u4_n160 ) , .B1( u2_u12_u4_n161 ) , .ZN( u2_u12_u4_n162 ) , .A( u2_u12_u4_n170 ) );
  AOI21_X1 u2_u12_u4_U14 (.ZN( u2_u12_u4_n107 ) , .B2( u2_u12_u4_n143 ) , .A( u2_u12_u4_n174 ) , .B1( u2_u12_u4_n184 ) );
  AOI21_X1 u2_u12_u4_U15 (.B2( u2_u12_u4_n158 ) , .B1( u2_u12_u4_n159 ) , .ZN( u2_u12_u4_n163 ) , .A( u2_u12_u4_n174 ) );
  AOI21_X1 u2_u12_u4_U16 (.A( u2_u12_u4_n153 ) , .B2( u2_u12_u4_n154 ) , .B1( u2_u12_u4_n155 ) , .ZN( u2_u12_u4_n165 ) );
  AOI21_X1 u2_u12_u4_U17 (.A( u2_u12_u4_n156 ) , .B2( u2_u12_u4_n157 ) , .ZN( u2_u12_u4_n164 ) , .B1( u2_u12_u4_n184 ) );
  INV_X1 u2_u12_u4_U18 (.A( u2_u12_u4_n138 ) , .ZN( u2_u12_u4_n170 ) );
  AND2_X1 u2_u12_u4_U19 (.A2( u2_u12_u4_n120 ) , .ZN( u2_u12_u4_n155 ) , .A1( u2_u12_u4_n160 ) );
  INV_X1 u2_u12_u4_U20 (.A( u2_u12_u4_n156 ) , .ZN( u2_u12_u4_n175 ) );
  NAND2_X1 u2_u12_u4_U21 (.A2( u2_u12_u4_n118 ) , .ZN( u2_u12_u4_n131 ) , .A1( u2_u12_u4_n147 ) );
  NAND2_X1 u2_u12_u4_U22 (.A1( u2_u12_u4_n119 ) , .A2( u2_u12_u4_n120 ) , .ZN( u2_u12_u4_n130 ) );
  NAND2_X1 u2_u12_u4_U23 (.ZN( u2_u12_u4_n117 ) , .A2( u2_u12_u4_n118 ) , .A1( u2_u12_u4_n148 ) );
  NAND2_X1 u2_u12_u4_U24 (.ZN( u2_u12_u4_n129 ) , .A1( u2_u12_u4_n134 ) , .A2( u2_u12_u4_n148 ) );
  AND3_X1 u2_u12_u4_U25 (.A1( u2_u12_u4_n119 ) , .A2( u2_u12_u4_n143 ) , .A3( u2_u12_u4_n154 ) , .ZN( u2_u12_u4_n161 ) );
  AND2_X1 u2_u12_u4_U26 (.A1( u2_u12_u4_n145 ) , .A2( u2_u12_u4_n147 ) , .ZN( u2_u12_u4_n159 ) );
  OR3_X1 u2_u12_u4_U27 (.A3( u2_u12_u4_n114 ) , .A2( u2_u12_u4_n115 ) , .A1( u2_u12_u4_n116 ) , .ZN( u2_u12_u4_n136 ) );
  AOI21_X1 u2_u12_u4_U28 (.A( u2_u12_u4_n113 ) , .ZN( u2_u12_u4_n116 ) , .B2( u2_u12_u4_n173 ) , .B1( u2_u12_u4_n174 ) );
  AOI21_X1 u2_u12_u4_U29 (.ZN( u2_u12_u4_n115 ) , .B2( u2_u12_u4_n145 ) , .B1( u2_u12_u4_n146 ) , .A( u2_u12_u4_n156 ) );
  NOR2_X1 u2_u12_u4_U3 (.ZN( u2_u12_u4_n121 ) , .A1( u2_u12_u4_n181 ) , .A2( u2_u12_u4_n182 ) );
  OAI22_X1 u2_u12_u4_U30 (.ZN( u2_u12_u4_n114 ) , .A2( u2_u12_u4_n121 ) , .B1( u2_u12_u4_n160 ) , .B2( u2_u12_u4_n170 ) , .A1( u2_u12_u4_n171 ) );
  INV_X1 u2_u12_u4_U31 (.A( u2_u12_u4_n158 ) , .ZN( u2_u12_u4_n182 ) );
  INV_X1 u2_u12_u4_U32 (.ZN( u2_u12_u4_n181 ) , .A( u2_u12_u4_n96 ) );
  INV_X1 u2_u12_u4_U33 (.A( u2_u12_u4_n144 ) , .ZN( u2_u12_u4_n179 ) );
  INV_X1 u2_u12_u4_U34 (.A( u2_u12_u4_n157 ) , .ZN( u2_u12_u4_n178 ) );
  NAND2_X1 u2_u12_u4_U35 (.A2( u2_u12_u4_n154 ) , .A1( u2_u12_u4_n96 ) , .ZN( u2_u12_u4_n97 ) );
  INV_X1 u2_u12_u4_U36 (.ZN( u2_u12_u4_n186 ) , .A( u2_u12_u4_n95 ) );
  OAI221_X1 u2_u12_u4_U37 (.C1( u2_u12_u4_n134 ) , .B1( u2_u12_u4_n158 ) , .B2( u2_u12_u4_n171 ) , .C2( u2_u12_u4_n173 ) , .A( u2_u12_u4_n94 ) , .ZN( u2_u12_u4_n95 ) );
  AOI222_X1 u2_u12_u4_U38 (.B2( u2_u12_u4_n132 ) , .A1( u2_u12_u4_n138 ) , .C2( u2_u12_u4_n175 ) , .A2( u2_u12_u4_n179 ) , .C1( u2_u12_u4_n181 ) , .B1( u2_u12_u4_n185 ) , .ZN( u2_u12_u4_n94 ) );
  INV_X1 u2_u12_u4_U39 (.A( u2_u12_u4_n113 ) , .ZN( u2_u12_u4_n185 ) );
  INV_X1 u2_u12_u4_U4 (.A( u2_u12_u4_n117 ) , .ZN( u2_u12_u4_n184 ) );
  INV_X1 u2_u12_u4_U40 (.A( u2_u12_u4_n143 ) , .ZN( u2_u12_u4_n183 ) );
  NOR2_X1 u2_u12_u4_U41 (.ZN( u2_u12_u4_n138 ) , .A1( u2_u12_u4_n168 ) , .A2( u2_u12_u4_n169 ) );
  NOR2_X1 u2_u12_u4_U42 (.A1( u2_u12_u4_n150 ) , .A2( u2_u12_u4_n152 ) , .ZN( u2_u12_u4_n153 ) );
  NOR2_X1 u2_u12_u4_U43 (.A2( u2_u12_u4_n128 ) , .A1( u2_u12_u4_n138 ) , .ZN( u2_u12_u4_n156 ) );
  AOI22_X1 u2_u12_u4_U44 (.B2( u2_u12_u4_n122 ) , .A1( u2_u12_u4_n123 ) , .ZN( u2_u12_u4_n124 ) , .B1( u2_u12_u4_n128 ) , .A2( u2_u12_u4_n172 ) );
  INV_X1 u2_u12_u4_U45 (.A( u2_u12_u4_n153 ) , .ZN( u2_u12_u4_n172 ) );
  NAND2_X1 u2_u12_u4_U46 (.A2( u2_u12_u4_n120 ) , .ZN( u2_u12_u4_n123 ) , .A1( u2_u12_u4_n161 ) );
  AOI22_X1 u2_u12_u4_U47 (.B2( u2_u12_u4_n132 ) , .A2( u2_u12_u4_n133 ) , .ZN( u2_u12_u4_n140 ) , .A1( u2_u12_u4_n150 ) , .B1( u2_u12_u4_n179 ) );
  NAND2_X1 u2_u12_u4_U48 (.ZN( u2_u12_u4_n133 ) , .A2( u2_u12_u4_n146 ) , .A1( u2_u12_u4_n154 ) );
  NAND2_X1 u2_u12_u4_U49 (.A1( u2_u12_u4_n103 ) , .ZN( u2_u12_u4_n154 ) , .A2( u2_u12_u4_n98 ) );
  NOR4_X1 u2_u12_u4_U5 (.A4( u2_u12_u4_n106 ) , .A3( u2_u12_u4_n107 ) , .A2( u2_u12_u4_n108 ) , .A1( u2_u12_u4_n109 ) , .ZN( u2_u12_u4_n110 ) );
  NAND2_X1 u2_u12_u4_U50 (.A1( u2_u12_u4_n101 ) , .ZN( u2_u12_u4_n158 ) , .A2( u2_u12_u4_n99 ) );
  AOI21_X1 u2_u12_u4_U51 (.ZN( u2_u12_u4_n127 ) , .A( u2_u12_u4_n136 ) , .B2( u2_u12_u4_n150 ) , .B1( u2_u12_u4_n180 ) );
  INV_X1 u2_u12_u4_U52 (.A( u2_u12_u4_n160 ) , .ZN( u2_u12_u4_n180 ) );
  NAND2_X1 u2_u12_u4_U53 (.A2( u2_u12_u4_n104 ) , .A1( u2_u12_u4_n105 ) , .ZN( u2_u12_u4_n146 ) );
  NAND2_X1 u2_u12_u4_U54 (.A2( u2_u12_u4_n101 ) , .A1( u2_u12_u4_n102 ) , .ZN( u2_u12_u4_n160 ) );
  NAND2_X1 u2_u12_u4_U55 (.ZN( u2_u12_u4_n134 ) , .A1( u2_u12_u4_n98 ) , .A2( u2_u12_u4_n99 ) );
  NAND2_X1 u2_u12_u4_U56 (.A1( u2_u12_u4_n103 ) , .A2( u2_u12_u4_n104 ) , .ZN( u2_u12_u4_n143 ) );
  NAND2_X1 u2_u12_u4_U57 (.A2( u2_u12_u4_n105 ) , .ZN( u2_u12_u4_n145 ) , .A1( u2_u12_u4_n98 ) );
  NAND2_X1 u2_u12_u4_U58 (.A1( u2_u12_u4_n100 ) , .A2( u2_u12_u4_n105 ) , .ZN( u2_u12_u4_n120 ) );
  NAND2_X1 u2_u12_u4_U59 (.A1( u2_u12_u4_n102 ) , .A2( u2_u12_u4_n104 ) , .ZN( u2_u12_u4_n148 ) );
  AOI21_X1 u2_u12_u4_U6 (.ZN( u2_u12_u4_n106 ) , .B2( u2_u12_u4_n146 ) , .B1( u2_u12_u4_n158 ) , .A( u2_u12_u4_n170 ) );
  NAND2_X1 u2_u12_u4_U60 (.A2( u2_u12_u4_n100 ) , .A1( u2_u12_u4_n103 ) , .ZN( u2_u12_u4_n157 ) );
  INV_X1 u2_u12_u4_U61 (.A( u2_u12_u4_n150 ) , .ZN( u2_u12_u4_n173 ) );
  INV_X1 u2_u12_u4_U62 (.A( u2_u12_u4_n152 ) , .ZN( u2_u12_u4_n171 ) );
  NAND2_X1 u2_u12_u4_U63 (.A1( u2_u12_u4_n100 ) , .ZN( u2_u12_u4_n118 ) , .A2( u2_u12_u4_n99 ) );
  NAND2_X1 u2_u12_u4_U64 (.A2( u2_u12_u4_n100 ) , .A1( u2_u12_u4_n102 ) , .ZN( u2_u12_u4_n144 ) );
  NAND2_X1 u2_u12_u4_U65 (.A2( u2_u12_u4_n101 ) , .A1( u2_u12_u4_n105 ) , .ZN( u2_u12_u4_n96 ) );
  INV_X1 u2_u12_u4_U66 (.A( u2_u12_u4_n128 ) , .ZN( u2_u12_u4_n174 ) );
  NAND2_X1 u2_u12_u4_U67 (.A2( u2_u12_u4_n102 ) , .ZN( u2_u12_u4_n119 ) , .A1( u2_u12_u4_n98 ) );
  NAND2_X1 u2_u12_u4_U68 (.A2( u2_u12_u4_n101 ) , .A1( u2_u12_u4_n103 ) , .ZN( u2_u12_u4_n147 ) );
  NAND2_X1 u2_u12_u4_U69 (.A2( u2_u12_u4_n104 ) , .ZN( u2_u12_u4_n113 ) , .A1( u2_u12_u4_n99 ) );
  AOI21_X1 u2_u12_u4_U7 (.ZN( u2_u12_u4_n108 ) , .B2( u2_u12_u4_n134 ) , .B1( u2_u12_u4_n155 ) , .A( u2_u12_u4_n156 ) );
  NOR2_X1 u2_u12_u4_U70 (.A2( u2_u12_X_28 ) , .ZN( u2_u12_u4_n150 ) , .A1( u2_u12_u4_n168 ) );
  NOR2_X1 u2_u12_u4_U71 (.A2( u2_u12_X_29 ) , .ZN( u2_u12_u4_n152 ) , .A1( u2_u12_u4_n169 ) );
  NOR2_X1 u2_u12_u4_U72 (.A2( u2_u12_X_30 ) , .ZN( u2_u12_u4_n105 ) , .A1( u2_u12_u4_n176 ) );
  NOR2_X1 u2_u12_u4_U73 (.A2( u2_u12_X_26 ) , .ZN( u2_u12_u4_n100 ) , .A1( u2_u12_u4_n177 ) );
  NOR2_X1 u2_u12_u4_U74 (.A2( u2_u12_X_28 ) , .A1( u2_u12_X_29 ) , .ZN( u2_u12_u4_n128 ) );
  NOR2_X1 u2_u12_u4_U75 (.A2( u2_u12_X_27 ) , .A1( u2_u12_X_30 ) , .ZN( u2_u12_u4_n102 ) );
  NOR2_X1 u2_u12_u4_U76 (.A2( u2_u12_X_25 ) , .A1( u2_u12_X_26 ) , .ZN( u2_u12_u4_n98 ) );
  AND2_X1 u2_u12_u4_U77 (.A2( u2_u12_X_25 ) , .A1( u2_u12_X_26 ) , .ZN( u2_u12_u4_n104 ) );
  AND2_X1 u2_u12_u4_U78 (.A1( u2_u12_X_30 ) , .A2( u2_u12_u4_n176 ) , .ZN( u2_u12_u4_n99 ) );
  AND2_X1 u2_u12_u4_U79 (.A1( u2_u12_X_26 ) , .ZN( u2_u12_u4_n101 ) , .A2( u2_u12_u4_n177 ) );
  AOI21_X1 u2_u12_u4_U8 (.ZN( u2_u12_u4_n109 ) , .A( u2_u12_u4_n153 ) , .B1( u2_u12_u4_n159 ) , .B2( u2_u12_u4_n184 ) );
  AND2_X1 u2_u12_u4_U80 (.A1( u2_u12_X_27 ) , .A2( u2_u12_X_30 ) , .ZN( u2_u12_u4_n103 ) );
  INV_X1 u2_u12_u4_U81 (.A( u2_u12_X_28 ) , .ZN( u2_u12_u4_n169 ) );
  INV_X1 u2_u12_u4_U82 (.A( u2_u12_X_29 ) , .ZN( u2_u12_u4_n168 ) );
  INV_X1 u2_u12_u4_U83 (.A( u2_u12_X_25 ) , .ZN( u2_u12_u4_n177 ) );
  INV_X1 u2_u12_u4_U84 (.A( u2_u12_X_27 ) , .ZN( u2_u12_u4_n176 ) );
  NAND4_X1 u2_u12_u4_U85 (.ZN( u2_out12_25 ) , .A4( u2_u12_u4_n139 ) , .A3( u2_u12_u4_n140 ) , .A2( u2_u12_u4_n141 ) , .A1( u2_u12_u4_n142 ) );
  OAI21_X1 u2_u12_u4_U86 (.A( u2_u12_u4_n128 ) , .B2( u2_u12_u4_n129 ) , .B1( u2_u12_u4_n130 ) , .ZN( u2_u12_u4_n142 ) );
  OAI21_X1 u2_u12_u4_U87 (.B2( u2_u12_u4_n131 ) , .ZN( u2_u12_u4_n141 ) , .A( u2_u12_u4_n175 ) , .B1( u2_u12_u4_n183 ) );
  NAND4_X1 u2_u12_u4_U88 (.ZN( u2_out12_14 ) , .A4( u2_u12_u4_n124 ) , .A3( u2_u12_u4_n125 ) , .A2( u2_u12_u4_n126 ) , .A1( u2_u12_u4_n127 ) );
  AOI22_X1 u2_u12_u4_U89 (.B2( u2_u12_u4_n117 ) , .ZN( u2_u12_u4_n126 ) , .A1( u2_u12_u4_n129 ) , .B1( u2_u12_u4_n152 ) , .A2( u2_u12_u4_n175 ) );
  AOI211_X1 u2_u12_u4_U9 (.B( u2_u12_u4_n136 ) , .A( u2_u12_u4_n137 ) , .C2( u2_u12_u4_n138 ) , .ZN( u2_u12_u4_n139 ) , .C1( u2_u12_u4_n182 ) );
  AOI22_X1 u2_u12_u4_U90 (.ZN( u2_u12_u4_n125 ) , .B2( u2_u12_u4_n131 ) , .A2( u2_u12_u4_n132 ) , .B1( u2_u12_u4_n138 ) , .A1( u2_u12_u4_n178 ) );
  NAND4_X1 u2_u12_u4_U91 (.ZN( u2_out12_8 ) , .A4( u2_u12_u4_n110 ) , .A3( u2_u12_u4_n111 ) , .A2( u2_u12_u4_n112 ) , .A1( u2_u12_u4_n186 ) );
  NAND2_X1 u2_u12_u4_U92 (.ZN( u2_u12_u4_n112 ) , .A2( u2_u12_u4_n130 ) , .A1( u2_u12_u4_n150 ) );
  AOI22_X1 u2_u12_u4_U93 (.ZN( u2_u12_u4_n111 ) , .B2( u2_u12_u4_n132 ) , .A1( u2_u12_u4_n152 ) , .B1( u2_u12_u4_n178 ) , .A2( u2_u12_u4_n97 ) );
  AOI22_X1 u2_u12_u4_U94 (.B2( u2_u12_u4_n149 ) , .B1( u2_u12_u4_n150 ) , .A2( u2_u12_u4_n151 ) , .A1( u2_u12_u4_n152 ) , .ZN( u2_u12_u4_n167 ) );
  NOR4_X1 u2_u12_u4_U95 (.A4( u2_u12_u4_n162 ) , .A3( u2_u12_u4_n163 ) , .A2( u2_u12_u4_n164 ) , .A1( u2_u12_u4_n165 ) , .ZN( u2_u12_u4_n166 ) );
  NAND3_X1 u2_u12_u4_U96 (.ZN( u2_out12_3 ) , .A3( u2_u12_u4_n166 ) , .A1( u2_u12_u4_n167 ) , .A2( u2_u12_u4_n186 ) );
  NAND3_X1 u2_u12_u4_U97 (.A3( u2_u12_u4_n146 ) , .A2( u2_u12_u4_n147 ) , .A1( u2_u12_u4_n148 ) , .ZN( u2_u12_u4_n149 ) );
  NAND3_X1 u2_u12_u4_U98 (.A3( u2_u12_u4_n143 ) , .A2( u2_u12_u4_n144 ) , .A1( u2_u12_u4_n145 ) , .ZN( u2_u12_u4_n151 ) );
  NAND3_X1 u2_u12_u4_U99 (.A3( u2_u12_u4_n121 ) , .ZN( u2_u12_u4_n122 ) , .A2( u2_u12_u4_n144 ) , .A1( u2_u12_u4_n154 ) );
  INV_X1 u2_u12_u5_U10 (.A( u2_u12_u5_n121 ) , .ZN( u2_u12_u5_n177 ) );
  NOR3_X1 u2_u12_u5_U100 (.A3( u2_u12_u5_n141 ) , .A1( u2_u12_u5_n142 ) , .ZN( u2_u12_u5_n143 ) , .A2( u2_u12_u5_n191 ) );
  NAND4_X1 u2_u12_u5_U101 (.ZN( u2_out12_4 ) , .A4( u2_u12_u5_n112 ) , .A2( u2_u12_u5_n113 ) , .A1( u2_u12_u5_n114 ) , .A3( u2_u12_u5_n195 ) );
  AOI211_X1 u2_u12_u5_U102 (.A( u2_u12_u5_n110 ) , .C1( u2_u12_u5_n111 ) , .ZN( u2_u12_u5_n112 ) , .B( u2_u12_u5_n118 ) , .C2( u2_u12_u5_n177 ) );
  AOI222_X1 u2_u12_u5_U103 (.ZN( u2_u12_u5_n113 ) , .A1( u2_u12_u5_n131 ) , .C1( u2_u12_u5_n148 ) , .B2( u2_u12_u5_n174 ) , .C2( u2_u12_u5_n178 ) , .A2( u2_u12_u5_n179 ) , .B1( u2_u12_u5_n99 ) );
  NAND3_X1 u2_u12_u5_U104 (.A2( u2_u12_u5_n154 ) , .A3( u2_u12_u5_n158 ) , .A1( u2_u12_u5_n161 ) , .ZN( u2_u12_u5_n99 ) );
  NOR2_X1 u2_u12_u5_U11 (.ZN( u2_u12_u5_n160 ) , .A2( u2_u12_u5_n173 ) , .A1( u2_u12_u5_n177 ) );
  INV_X1 u2_u12_u5_U12 (.A( u2_u12_u5_n150 ) , .ZN( u2_u12_u5_n174 ) );
  AOI21_X1 u2_u12_u5_U13 (.A( u2_u12_u5_n160 ) , .B2( u2_u12_u5_n161 ) , .ZN( u2_u12_u5_n162 ) , .B1( u2_u12_u5_n192 ) );
  INV_X1 u2_u12_u5_U14 (.A( u2_u12_u5_n159 ) , .ZN( u2_u12_u5_n192 ) );
  AOI21_X1 u2_u12_u5_U15 (.A( u2_u12_u5_n156 ) , .B2( u2_u12_u5_n157 ) , .B1( u2_u12_u5_n158 ) , .ZN( u2_u12_u5_n163 ) );
  AOI21_X1 u2_u12_u5_U16 (.B2( u2_u12_u5_n139 ) , .B1( u2_u12_u5_n140 ) , .ZN( u2_u12_u5_n141 ) , .A( u2_u12_u5_n150 ) );
  OAI21_X1 u2_u12_u5_U17 (.A( u2_u12_u5_n133 ) , .B2( u2_u12_u5_n134 ) , .B1( u2_u12_u5_n135 ) , .ZN( u2_u12_u5_n142 ) );
  OAI21_X1 u2_u12_u5_U18 (.ZN( u2_u12_u5_n133 ) , .B2( u2_u12_u5_n147 ) , .A( u2_u12_u5_n173 ) , .B1( u2_u12_u5_n188 ) );
  NAND2_X1 u2_u12_u5_U19 (.A2( u2_u12_u5_n119 ) , .A1( u2_u12_u5_n123 ) , .ZN( u2_u12_u5_n137 ) );
  INV_X1 u2_u12_u5_U20 (.A( u2_u12_u5_n155 ) , .ZN( u2_u12_u5_n194 ) );
  NAND2_X1 u2_u12_u5_U21 (.A1( u2_u12_u5_n121 ) , .ZN( u2_u12_u5_n132 ) , .A2( u2_u12_u5_n172 ) );
  NAND2_X1 u2_u12_u5_U22 (.A2( u2_u12_u5_n122 ) , .ZN( u2_u12_u5_n136 ) , .A1( u2_u12_u5_n154 ) );
  NAND2_X1 u2_u12_u5_U23 (.A2( u2_u12_u5_n119 ) , .A1( u2_u12_u5_n120 ) , .ZN( u2_u12_u5_n159 ) );
  INV_X1 u2_u12_u5_U24 (.A( u2_u12_u5_n156 ) , .ZN( u2_u12_u5_n175 ) );
  INV_X1 u2_u12_u5_U25 (.A( u2_u12_u5_n158 ) , .ZN( u2_u12_u5_n188 ) );
  INV_X1 u2_u12_u5_U26 (.A( u2_u12_u5_n152 ) , .ZN( u2_u12_u5_n179 ) );
  INV_X1 u2_u12_u5_U27 (.A( u2_u12_u5_n140 ) , .ZN( u2_u12_u5_n182 ) );
  INV_X1 u2_u12_u5_U28 (.A( u2_u12_u5_n151 ) , .ZN( u2_u12_u5_n183 ) );
  INV_X1 u2_u12_u5_U29 (.A( u2_u12_u5_n123 ) , .ZN( u2_u12_u5_n185 ) );
  NOR2_X1 u2_u12_u5_U3 (.ZN( u2_u12_u5_n134 ) , .A1( u2_u12_u5_n183 ) , .A2( u2_u12_u5_n190 ) );
  INV_X1 u2_u12_u5_U30 (.A( u2_u12_u5_n161 ) , .ZN( u2_u12_u5_n184 ) );
  INV_X1 u2_u12_u5_U31 (.A( u2_u12_u5_n139 ) , .ZN( u2_u12_u5_n189 ) );
  INV_X1 u2_u12_u5_U32 (.A( u2_u12_u5_n157 ) , .ZN( u2_u12_u5_n190 ) );
  INV_X1 u2_u12_u5_U33 (.A( u2_u12_u5_n120 ) , .ZN( u2_u12_u5_n193 ) );
  NAND2_X1 u2_u12_u5_U34 (.ZN( u2_u12_u5_n111 ) , .A1( u2_u12_u5_n140 ) , .A2( u2_u12_u5_n155 ) );
  NOR2_X1 u2_u12_u5_U35 (.ZN( u2_u12_u5_n100 ) , .A1( u2_u12_u5_n170 ) , .A2( u2_u12_u5_n180 ) );
  INV_X1 u2_u12_u5_U36 (.A( u2_u12_u5_n117 ) , .ZN( u2_u12_u5_n196 ) );
  OAI221_X1 u2_u12_u5_U37 (.A( u2_u12_u5_n116 ) , .ZN( u2_u12_u5_n117 ) , .B2( u2_u12_u5_n119 ) , .C1( u2_u12_u5_n153 ) , .C2( u2_u12_u5_n158 ) , .B1( u2_u12_u5_n172 ) );
  AOI222_X1 u2_u12_u5_U38 (.ZN( u2_u12_u5_n116 ) , .B2( u2_u12_u5_n145 ) , .C1( u2_u12_u5_n148 ) , .A2( u2_u12_u5_n174 ) , .C2( u2_u12_u5_n177 ) , .B1( u2_u12_u5_n187 ) , .A1( u2_u12_u5_n193 ) );
  INV_X1 u2_u12_u5_U39 (.A( u2_u12_u5_n115 ) , .ZN( u2_u12_u5_n187 ) );
  INV_X1 u2_u12_u5_U4 (.A( u2_u12_u5_n138 ) , .ZN( u2_u12_u5_n191 ) );
  AOI22_X1 u2_u12_u5_U40 (.B2( u2_u12_u5_n131 ) , .A2( u2_u12_u5_n146 ) , .ZN( u2_u12_u5_n169 ) , .B1( u2_u12_u5_n174 ) , .A1( u2_u12_u5_n185 ) );
  NOR2_X1 u2_u12_u5_U41 (.A1( u2_u12_u5_n146 ) , .ZN( u2_u12_u5_n150 ) , .A2( u2_u12_u5_n173 ) );
  AOI21_X1 u2_u12_u5_U42 (.A( u2_u12_u5_n118 ) , .B2( u2_u12_u5_n145 ) , .ZN( u2_u12_u5_n168 ) , .B1( u2_u12_u5_n186 ) );
  INV_X1 u2_u12_u5_U43 (.A( u2_u12_u5_n122 ) , .ZN( u2_u12_u5_n186 ) );
  NOR2_X1 u2_u12_u5_U44 (.A1( u2_u12_u5_n146 ) , .ZN( u2_u12_u5_n152 ) , .A2( u2_u12_u5_n176 ) );
  NOR2_X1 u2_u12_u5_U45 (.A1( u2_u12_u5_n115 ) , .ZN( u2_u12_u5_n118 ) , .A2( u2_u12_u5_n153 ) );
  NOR2_X1 u2_u12_u5_U46 (.A2( u2_u12_u5_n145 ) , .ZN( u2_u12_u5_n156 ) , .A1( u2_u12_u5_n174 ) );
  NOR2_X1 u2_u12_u5_U47 (.ZN( u2_u12_u5_n121 ) , .A2( u2_u12_u5_n145 ) , .A1( u2_u12_u5_n176 ) );
  AOI22_X1 u2_u12_u5_U48 (.ZN( u2_u12_u5_n114 ) , .A2( u2_u12_u5_n137 ) , .A1( u2_u12_u5_n145 ) , .B2( u2_u12_u5_n175 ) , .B1( u2_u12_u5_n193 ) );
  OAI211_X1 u2_u12_u5_U49 (.B( u2_u12_u5_n124 ) , .A( u2_u12_u5_n125 ) , .C2( u2_u12_u5_n126 ) , .C1( u2_u12_u5_n127 ) , .ZN( u2_u12_u5_n128 ) );
  OAI21_X1 u2_u12_u5_U5 (.B2( u2_u12_u5_n136 ) , .B1( u2_u12_u5_n137 ) , .ZN( u2_u12_u5_n138 ) , .A( u2_u12_u5_n177 ) );
  NOR3_X1 u2_u12_u5_U50 (.ZN( u2_u12_u5_n127 ) , .A1( u2_u12_u5_n136 ) , .A3( u2_u12_u5_n148 ) , .A2( u2_u12_u5_n182 ) );
  OAI21_X1 u2_u12_u5_U51 (.ZN( u2_u12_u5_n124 ) , .A( u2_u12_u5_n177 ) , .B2( u2_u12_u5_n183 ) , .B1( u2_u12_u5_n189 ) );
  OAI21_X1 u2_u12_u5_U52 (.ZN( u2_u12_u5_n125 ) , .A( u2_u12_u5_n174 ) , .B2( u2_u12_u5_n185 ) , .B1( u2_u12_u5_n190 ) );
  AOI21_X1 u2_u12_u5_U53 (.A( u2_u12_u5_n153 ) , .B2( u2_u12_u5_n154 ) , .B1( u2_u12_u5_n155 ) , .ZN( u2_u12_u5_n164 ) );
  AOI21_X1 u2_u12_u5_U54 (.ZN( u2_u12_u5_n110 ) , .B1( u2_u12_u5_n122 ) , .B2( u2_u12_u5_n139 ) , .A( u2_u12_u5_n153 ) );
  INV_X1 u2_u12_u5_U55 (.A( u2_u12_u5_n153 ) , .ZN( u2_u12_u5_n176 ) );
  INV_X1 u2_u12_u5_U56 (.A( u2_u12_u5_n126 ) , .ZN( u2_u12_u5_n173 ) );
  AND2_X1 u2_u12_u5_U57 (.A2( u2_u12_u5_n104 ) , .A1( u2_u12_u5_n107 ) , .ZN( u2_u12_u5_n147 ) );
  AND2_X1 u2_u12_u5_U58 (.A2( u2_u12_u5_n104 ) , .A1( u2_u12_u5_n108 ) , .ZN( u2_u12_u5_n148 ) );
  NAND2_X1 u2_u12_u5_U59 (.A1( u2_u12_u5_n105 ) , .A2( u2_u12_u5_n106 ) , .ZN( u2_u12_u5_n158 ) );
  INV_X1 u2_u12_u5_U6 (.A( u2_u12_u5_n135 ) , .ZN( u2_u12_u5_n178 ) );
  NAND2_X1 u2_u12_u5_U60 (.A2( u2_u12_u5_n108 ) , .A1( u2_u12_u5_n109 ) , .ZN( u2_u12_u5_n139 ) );
  NAND2_X1 u2_u12_u5_U61 (.A1( u2_u12_u5_n106 ) , .A2( u2_u12_u5_n108 ) , .ZN( u2_u12_u5_n119 ) );
  NAND2_X1 u2_u12_u5_U62 (.A2( u2_u12_u5_n103 ) , .A1( u2_u12_u5_n105 ) , .ZN( u2_u12_u5_n140 ) );
  NAND2_X1 u2_u12_u5_U63 (.A2( u2_u12_u5_n104 ) , .A1( u2_u12_u5_n105 ) , .ZN( u2_u12_u5_n155 ) );
  NAND2_X1 u2_u12_u5_U64 (.A2( u2_u12_u5_n106 ) , .A1( u2_u12_u5_n107 ) , .ZN( u2_u12_u5_n122 ) );
  NAND2_X1 u2_u12_u5_U65 (.A2( u2_u12_u5_n100 ) , .A1( u2_u12_u5_n106 ) , .ZN( u2_u12_u5_n115 ) );
  NAND2_X1 u2_u12_u5_U66 (.A2( u2_u12_u5_n100 ) , .A1( u2_u12_u5_n103 ) , .ZN( u2_u12_u5_n161 ) );
  NAND2_X1 u2_u12_u5_U67 (.A1( u2_u12_u5_n105 ) , .A2( u2_u12_u5_n109 ) , .ZN( u2_u12_u5_n154 ) );
  INV_X1 u2_u12_u5_U68 (.A( u2_u12_u5_n146 ) , .ZN( u2_u12_u5_n172 ) );
  NAND2_X1 u2_u12_u5_U69 (.A1( u2_u12_u5_n103 ) , .A2( u2_u12_u5_n108 ) , .ZN( u2_u12_u5_n123 ) );
  OAI22_X1 u2_u12_u5_U7 (.B2( u2_u12_u5_n149 ) , .B1( u2_u12_u5_n150 ) , .A2( u2_u12_u5_n151 ) , .A1( u2_u12_u5_n152 ) , .ZN( u2_u12_u5_n165 ) );
  NAND2_X1 u2_u12_u5_U70 (.A2( u2_u12_u5_n103 ) , .A1( u2_u12_u5_n107 ) , .ZN( u2_u12_u5_n151 ) );
  NAND2_X1 u2_u12_u5_U71 (.A2( u2_u12_u5_n107 ) , .A1( u2_u12_u5_n109 ) , .ZN( u2_u12_u5_n120 ) );
  NAND2_X1 u2_u12_u5_U72 (.A2( u2_u12_u5_n100 ) , .A1( u2_u12_u5_n109 ) , .ZN( u2_u12_u5_n157 ) );
  AND2_X1 u2_u12_u5_U73 (.A2( u2_u12_u5_n100 ) , .A1( u2_u12_u5_n104 ) , .ZN( u2_u12_u5_n131 ) );
  INV_X1 u2_u12_u5_U74 (.A( u2_u12_u5_n102 ) , .ZN( u2_u12_u5_n195 ) );
  OAI221_X1 u2_u12_u5_U75 (.A( u2_u12_u5_n101 ) , .ZN( u2_u12_u5_n102 ) , .C2( u2_u12_u5_n115 ) , .C1( u2_u12_u5_n126 ) , .B1( u2_u12_u5_n134 ) , .B2( u2_u12_u5_n160 ) );
  OAI21_X1 u2_u12_u5_U76 (.ZN( u2_u12_u5_n101 ) , .B1( u2_u12_u5_n137 ) , .A( u2_u12_u5_n146 ) , .B2( u2_u12_u5_n147 ) );
  NOR2_X1 u2_u12_u5_U77 (.A2( u2_u12_X_34 ) , .A1( u2_u12_X_35 ) , .ZN( u2_u12_u5_n145 ) );
  NOR2_X1 u2_u12_u5_U78 (.A2( u2_u12_X_34 ) , .ZN( u2_u12_u5_n146 ) , .A1( u2_u12_u5_n171 ) );
  NOR2_X1 u2_u12_u5_U79 (.A2( u2_u12_X_31 ) , .A1( u2_u12_X_32 ) , .ZN( u2_u12_u5_n103 ) );
  NOR3_X1 u2_u12_u5_U8 (.A2( u2_u12_u5_n147 ) , .A1( u2_u12_u5_n148 ) , .ZN( u2_u12_u5_n149 ) , .A3( u2_u12_u5_n194 ) );
  NOR2_X1 u2_u12_u5_U80 (.A2( u2_u12_X_36 ) , .ZN( u2_u12_u5_n105 ) , .A1( u2_u12_u5_n180 ) );
  NOR2_X1 u2_u12_u5_U81 (.A2( u2_u12_X_33 ) , .ZN( u2_u12_u5_n108 ) , .A1( u2_u12_u5_n170 ) );
  NOR2_X1 u2_u12_u5_U82 (.A2( u2_u12_X_33 ) , .A1( u2_u12_X_36 ) , .ZN( u2_u12_u5_n107 ) );
  NOR2_X1 u2_u12_u5_U83 (.A2( u2_u12_X_31 ) , .ZN( u2_u12_u5_n104 ) , .A1( u2_u12_u5_n181 ) );
  NAND2_X1 u2_u12_u5_U84 (.A2( u2_u12_X_34 ) , .A1( u2_u12_X_35 ) , .ZN( u2_u12_u5_n153 ) );
  NAND2_X1 u2_u12_u5_U85 (.A1( u2_u12_X_34 ) , .ZN( u2_u12_u5_n126 ) , .A2( u2_u12_u5_n171 ) );
  AND2_X1 u2_u12_u5_U86 (.A1( u2_u12_X_31 ) , .A2( u2_u12_X_32 ) , .ZN( u2_u12_u5_n106 ) );
  AND2_X1 u2_u12_u5_U87 (.A1( u2_u12_X_31 ) , .ZN( u2_u12_u5_n109 ) , .A2( u2_u12_u5_n181 ) );
  INV_X1 u2_u12_u5_U88 (.A( u2_u12_X_33 ) , .ZN( u2_u12_u5_n180 ) );
  INV_X1 u2_u12_u5_U89 (.A( u2_u12_X_35 ) , .ZN( u2_u12_u5_n171 ) );
  NOR2_X1 u2_u12_u5_U9 (.ZN( u2_u12_u5_n135 ) , .A1( u2_u12_u5_n173 ) , .A2( u2_u12_u5_n176 ) );
  INV_X1 u2_u12_u5_U90 (.A( u2_u12_X_36 ) , .ZN( u2_u12_u5_n170 ) );
  INV_X1 u2_u12_u5_U91 (.A( u2_u12_X_32 ) , .ZN( u2_u12_u5_n181 ) );
  NAND4_X1 u2_u12_u5_U92 (.ZN( u2_out12_29 ) , .A4( u2_u12_u5_n129 ) , .A3( u2_u12_u5_n130 ) , .A2( u2_u12_u5_n168 ) , .A1( u2_u12_u5_n196 ) );
  AOI221_X1 u2_u12_u5_U93 (.A( u2_u12_u5_n128 ) , .ZN( u2_u12_u5_n129 ) , .C2( u2_u12_u5_n132 ) , .B2( u2_u12_u5_n159 ) , .B1( u2_u12_u5_n176 ) , .C1( u2_u12_u5_n184 ) );
  AOI222_X1 u2_u12_u5_U94 (.ZN( u2_u12_u5_n130 ) , .A2( u2_u12_u5_n146 ) , .B1( u2_u12_u5_n147 ) , .C2( u2_u12_u5_n175 ) , .B2( u2_u12_u5_n179 ) , .A1( u2_u12_u5_n188 ) , .C1( u2_u12_u5_n194 ) );
  NAND4_X1 u2_u12_u5_U95 (.ZN( u2_out12_19 ) , .A4( u2_u12_u5_n166 ) , .A3( u2_u12_u5_n167 ) , .A2( u2_u12_u5_n168 ) , .A1( u2_u12_u5_n169 ) );
  AOI22_X1 u2_u12_u5_U96 (.B2( u2_u12_u5_n145 ) , .A2( u2_u12_u5_n146 ) , .ZN( u2_u12_u5_n167 ) , .B1( u2_u12_u5_n182 ) , .A1( u2_u12_u5_n189 ) );
  NOR4_X1 u2_u12_u5_U97 (.A4( u2_u12_u5_n162 ) , .A3( u2_u12_u5_n163 ) , .A2( u2_u12_u5_n164 ) , .A1( u2_u12_u5_n165 ) , .ZN( u2_u12_u5_n166 ) );
  NAND4_X1 u2_u12_u5_U98 (.ZN( u2_out12_11 ) , .A4( u2_u12_u5_n143 ) , .A3( u2_u12_u5_n144 ) , .A2( u2_u12_u5_n169 ) , .A1( u2_u12_u5_n196 ) );
  AOI22_X1 u2_u12_u5_U99 (.A2( u2_u12_u5_n132 ) , .ZN( u2_u12_u5_n144 ) , .B2( u2_u12_u5_n145 ) , .B1( u2_u12_u5_n184 ) , .A1( u2_u12_u5_n194 ) );
  XOR2_X1 u2_u13_U26 (.B( u2_K14_30 ) , .A( u2_R12_21 ) , .Z( u2_u13_X_30 ) );
  XOR2_X1 u2_u13_U28 (.B( u2_K14_29 ) , .A( u2_R12_20 ) , .Z( u2_u13_X_29 ) );
  XOR2_X1 u2_u13_U29 (.B( u2_K14_28 ) , .A( u2_R12_19 ) , .Z( u2_u13_X_28 ) );
  XOR2_X1 u2_u13_U30 (.B( u2_K14_27 ) , .A( u2_R12_18 ) , .Z( u2_u13_X_27 ) );
  XOR2_X1 u2_u13_U31 (.B( u2_K14_26 ) , .A( u2_R12_17 ) , .Z( u2_u13_X_26 ) );
  XOR2_X1 u2_u13_U32 (.B( u2_K14_25 ) , .A( u2_R12_16 ) , .Z( u2_u13_X_25 ) );
  AOI21_X1 u2_u13_u4_U10 (.ZN( u2_u13_u4_n106 ) , .B2( u2_u13_u4_n146 ) , .B1( u2_u13_u4_n158 ) , .A( u2_u13_u4_n170 ) );
  AOI21_X1 u2_u13_u4_U11 (.ZN( u2_u13_u4_n108 ) , .B2( u2_u13_u4_n134 ) , .B1( u2_u13_u4_n155 ) , .A( u2_u13_u4_n156 ) );
  AOI21_X1 u2_u13_u4_U12 (.ZN( u2_u13_u4_n109 ) , .A( u2_u13_u4_n153 ) , .B1( u2_u13_u4_n159 ) , .B2( u2_u13_u4_n184 ) );
  AOI211_X1 u2_u13_u4_U13 (.B( u2_u13_u4_n136 ) , .A( u2_u13_u4_n137 ) , .C2( u2_u13_u4_n138 ) , .ZN( u2_u13_u4_n139 ) , .C1( u2_u13_u4_n182 ) );
  OAI22_X1 u2_u13_u4_U14 (.B2( u2_u13_u4_n135 ) , .ZN( u2_u13_u4_n137 ) , .B1( u2_u13_u4_n153 ) , .A1( u2_u13_u4_n155 ) , .A2( u2_u13_u4_n171 ) );
  AND3_X1 u2_u13_u4_U15 (.A2( u2_u13_u4_n134 ) , .ZN( u2_u13_u4_n135 ) , .A3( u2_u13_u4_n145 ) , .A1( u2_u13_u4_n157 ) );
  NAND2_X1 u2_u13_u4_U16 (.ZN( u2_u13_u4_n132 ) , .A2( u2_u13_u4_n170 ) , .A1( u2_u13_u4_n173 ) );
  AOI21_X1 u2_u13_u4_U17 (.B2( u2_u13_u4_n160 ) , .B1( u2_u13_u4_n161 ) , .ZN( u2_u13_u4_n162 ) , .A( u2_u13_u4_n170 ) );
  AOI21_X1 u2_u13_u4_U18 (.ZN( u2_u13_u4_n107 ) , .B2( u2_u13_u4_n143 ) , .A( u2_u13_u4_n174 ) , .B1( u2_u13_u4_n184 ) );
  AOI21_X1 u2_u13_u4_U19 (.B2( u2_u13_u4_n158 ) , .B1( u2_u13_u4_n159 ) , .ZN( u2_u13_u4_n163 ) , .A( u2_u13_u4_n174 ) );
  AOI21_X1 u2_u13_u4_U20 (.A( u2_u13_u4_n153 ) , .B2( u2_u13_u4_n154 ) , .B1( u2_u13_u4_n155 ) , .ZN( u2_u13_u4_n165 ) );
  AOI21_X1 u2_u13_u4_U21 (.A( u2_u13_u4_n156 ) , .B2( u2_u13_u4_n157 ) , .ZN( u2_u13_u4_n164 ) , .B1( u2_u13_u4_n184 ) );
  INV_X1 u2_u13_u4_U22 (.A( u2_u13_u4_n138 ) , .ZN( u2_u13_u4_n170 ) );
  AND2_X1 u2_u13_u4_U23 (.A2( u2_u13_u4_n120 ) , .ZN( u2_u13_u4_n155 ) , .A1( u2_u13_u4_n160 ) );
  INV_X1 u2_u13_u4_U24 (.A( u2_u13_u4_n156 ) , .ZN( u2_u13_u4_n175 ) );
  NAND2_X1 u2_u13_u4_U25 (.A2( u2_u13_u4_n118 ) , .ZN( u2_u13_u4_n131 ) , .A1( u2_u13_u4_n147 ) );
  NAND2_X1 u2_u13_u4_U26 (.A1( u2_u13_u4_n119 ) , .A2( u2_u13_u4_n120 ) , .ZN( u2_u13_u4_n130 ) );
  NAND2_X1 u2_u13_u4_U27 (.ZN( u2_u13_u4_n117 ) , .A2( u2_u13_u4_n118 ) , .A1( u2_u13_u4_n148 ) );
  NAND2_X1 u2_u13_u4_U28 (.ZN( u2_u13_u4_n129 ) , .A1( u2_u13_u4_n134 ) , .A2( u2_u13_u4_n148 ) );
  AND3_X1 u2_u13_u4_U29 (.A1( u2_u13_u4_n119 ) , .A2( u2_u13_u4_n143 ) , .A3( u2_u13_u4_n154 ) , .ZN( u2_u13_u4_n161 ) );
  NOR2_X1 u2_u13_u4_U3 (.ZN( u2_u13_u4_n121 ) , .A1( u2_u13_u4_n181 ) , .A2( u2_u13_u4_n182 ) );
  AND2_X1 u2_u13_u4_U30 (.A1( u2_u13_u4_n145 ) , .A2( u2_u13_u4_n147 ) , .ZN( u2_u13_u4_n159 ) );
  OR3_X1 u2_u13_u4_U31 (.A3( u2_u13_u4_n114 ) , .A2( u2_u13_u4_n115 ) , .A1( u2_u13_u4_n116 ) , .ZN( u2_u13_u4_n136 ) );
  AOI21_X1 u2_u13_u4_U32 (.A( u2_u13_u4_n113 ) , .ZN( u2_u13_u4_n116 ) , .B2( u2_u13_u4_n173 ) , .B1( u2_u13_u4_n174 ) );
  AOI21_X1 u2_u13_u4_U33 (.ZN( u2_u13_u4_n115 ) , .B2( u2_u13_u4_n145 ) , .B1( u2_u13_u4_n146 ) , .A( u2_u13_u4_n156 ) );
  OAI22_X1 u2_u13_u4_U34 (.ZN( u2_u13_u4_n114 ) , .A2( u2_u13_u4_n121 ) , .B1( u2_u13_u4_n160 ) , .B2( u2_u13_u4_n170 ) , .A1( u2_u13_u4_n171 ) );
  INV_X1 u2_u13_u4_U35 (.A( u2_u13_u4_n158 ) , .ZN( u2_u13_u4_n182 ) );
  INV_X1 u2_u13_u4_U36 (.ZN( u2_u13_u4_n181 ) , .A( u2_u13_u4_n96 ) );
  INV_X1 u2_u13_u4_U37 (.A( u2_u13_u4_n144 ) , .ZN( u2_u13_u4_n179 ) );
  INV_X1 u2_u13_u4_U38 (.A( u2_u13_u4_n157 ) , .ZN( u2_u13_u4_n178 ) );
  NAND2_X1 u2_u13_u4_U39 (.A2( u2_u13_u4_n154 ) , .A1( u2_u13_u4_n96 ) , .ZN( u2_u13_u4_n97 ) );
  INV_X1 u2_u13_u4_U4 (.A( u2_u13_u4_n117 ) , .ZN( u2_u13_u4_n184 ) );
  INV_X1 u2_u13_u4_U40 (.A( u2_u13_u4_n143 ) , .ZN( u2_u13_u4_n183 ) );
  NOR2_X1 u2_u13_u4_U41 (.ZN( u2_u13_u4_n138 ) , .A1( u2_u13_u4_n168 ) , .A2( u2_u13_u4_n169 ) );
  NOR2_X1 u2_u13_u4_U42 (.A1( u2_u13_u4_n150 ) , .A2( u2_u13_u4_n152 ) , .ZN( u2_u13_u4_n153 ) );
  NOR2_X1 u2_u13_u4_U43 (.A2( u2_u13_u4_n128 ) , .A1( u2_u13_u4_n138 ) , .ZN( u2_u13_u4_n156 ) );
  AOI22_X1 u2_u13_u4_U44 (.B2( u2_u13_u4_n122 ) , .A1( u2_u13_u4_n123 ) , .ZN( u2_u13_u4_n124 ) , .B1( u2_u13_u4_n128 ) , .A2( u2_u13_u4_n172 ) );
  NAND2_X1 u2_u13_u4_U45 (.A2( u2_u13_u4_n120 ) , .ZN( u2_u13_u4_n123 ) , .A1( u2_u13_u4_n161 ) );
  INV_X1 u2_u13_u4_U46 (.A( u2_u13_u4_n153 ) , .ZN( u2_u13_u4_n172 ) );
  AOI22_X1 u2_u13_u4_U47 (.B2( u2_u13_u4_n132 ) , .A2( u2_u13_u4_n133 ) , .ZN( u2_u13_u4_n140 ) , .A1( u2_u13_u4_n150 ) , .B1( u2_u13_u4_n179 ) );
  NAND2_X1 u2_u13_u4_U48 (.ZN( u2_u13_u4_n133 ) , .A2( u2_u13_u4_n146 ) , .A1( u2_u13_u4_n154 ) );
  NAND2_X1 u2_u13_u4_U49 (.A1( u2_u13_u4_n103 ) , .ZN( u2_u13_u4_n154 ) , .A2( u2_u13_u4_n98 ) );
  INV_X1 u2_u13_u4_U5 (.ZN( u2_u13_u4_n186 ) , .A( u2_u13_u4_n95 ) );
  NAND2_X1 u2_u13_u4_U50 (.A1( u2_u13_u4_n101 ) , .ZN( u2_u13_u4_n158 ) , .A2( u2_u13_u4_n99 ) );
  AOI21_X1 u2_u13_u4_U51 (.ZN( u2_u13_u4_n127 ) , .A( u2_u13_u4_n136 ) , .B2( u2_u13_u4_n150 ) , .B1( u2_u13_u4_n180 ) );
  INV_X1 u2_u13_u4_U52 (.A( u2_u13_u4_n160 ) , .ZN( u2_u13_u4_n180 ) );
  NAND2_X1 u2_u13_u4_U53 (.A2( u2_u13_u4_n104 ) , .A1( u2_u13_u4_n105 ) , .ZN( u2_u13_u4_n146 ) );
  NAND2_X1 u2_u13_u4_U54 (.A2( u2_u13_u4_n101 ) , .A1( u2_u13_u4_n102 ) , .ZN( u2_u13_u4_n160 ) );
  NAND2_X1 u2_u13_u4_U55 (.ZN( u2_u13_u4_n134 ) , .A1( u2_u13_u4_n98 ) , .A2( u2_u13_u4_n99 ) );
  NAND2_X1 u2_u13_u4_U56 (.A1( u2_u13_u4_n103 ) , .A2( u2_u13_u4_n104 ) , .ZN( u2_u13_u4_n143 ) );
  NAND2_X1 u2_u13_u4_U57 (.A2( u2_u13_u4_n105 ) , .ZN( u2_u13_u4_n145 ) , .A1( u2_u13_u4_n98 ) );
  NAND2_X1 u2_u13_u4_U58 (.A1( u2_u13_u4_n100 ) , .A2( u2_u13_u4_n105 ) , .ZN( u2_u13_u4_n120 ) );
  NAND2_X1 u2_u13_u4_U59 (.A1( u2_u13_u4_n102 ) , .A2( u2_u13_u4_n104 ) , .ZN( u2_u13_u4_n148 ) );
  OAI221_X1 u2_u13_u4_U6 (.C1( u2_u13_u4_n134 ) , .B1( u2_u13_u4_n158 ) , .B2( u2_u13_u4_n171 ) , .C2( u2_u13_u4_n173 ) , .A( u2_u13_u4_n94 ) , .ZN( u2_u13_u4_n95 ) );
  NAND2_X1 u2_u13_u4_U60 (.A2( u2_u13_u4_n100 ) , .A1( u2_u13_u4_n103 ) , .ZN( u2_u13_u4_n157 ) );
  INV_X1 u2_u13_u4_U61 (.A( u2_u13_u4_n150 ) , .ZN( u2_u13_u4_n173 ) );
  INV_X1 u2_u13_u4_U62 (.A( u2_u13_u4_n152 ) , .ZN( u2_u13_u4_n171 ) );
  NAND2_X1 u2_u13_u4_U63 (.A1( u2_u13_u4_n100 ) , .ZN( u2_u13_u4_n118 ) , .A2( u2_u13_u4_n99 ) );
  NAND2_X1 u2_u13_u4_U64 (.A2( u2_u13_u4_n100 ) , .A1( u2_u13_u4_n102 ) , .ZN( u2_u13_u4_n144 ) );
  NAND2_X1 u2_u13_u4_U65 (.A2( u2_u13_u4_n101 ) , .A1( u2_u13_u4_n105 ) , .ZN( u2_u13_u4_n96 ) );
  INV_X1 u2_u13_u4_U66 (.A( u2_u13_u4_n128 ) , .ZN( u2_u13_u4_n174 ) );
  NAND2_X1 u2_u13_u4_U67 (.A2( u2_u13_u4_n102 ) , .ZN( u2_u13_u4_n119 ) , .A1( u2_u13_u4_n98 ) );
  NAND2_X1 u2_u13_u4_U68 (.A2( u2_u13_u4_n101 ) , .A1( u2_u13_u4_n103 ) , .ZN( u2_u13_u4_n147 ) );
  NAND2_X1 u2_u13_u4_U69 (.A2( u2_u13_u4_n104 ) , .ZN( u2_u13_u4_n113 ) , .A1( u2_u13_u4_n99 ) );
  AOI222_X1 u2_u13_u4_U7 (.B2( u2_u13_u4_n132 ) , .A1( u2_u13_u4_n138 ) , .C2( u2_u13_u4_n175 ) , .A2( u2_u13_u4_n179 ) , .C1( u2_u13_u4_n181 ) , .B1( u2_u13_u4_n185 ) , .ZN( u2_u13_u4_n94 ) );
  NOR2_X1 u2_u13_u4_U70 (.A2( u2_u13_X_28 ) , .ZN( u2_u13_u4_n150 ) , .A1( u2_u13_u4_n168 ) );
  NOR2_X1 u2_u13_u4_U71 (.A2( u2_u13_X_29 ) , .ZN( u2_u13_u4_n152 ) , .A1( u2_u13_u4_n169 ) );
  NOR2_X1 u2_u13_u4_U72 (.A2( u2_u13_X_30 ) , .ZN( u2_u13_u4_n105 ) , .A1( u2_u13_u4_n176 ) );
  NOR2_X1 u2_u13_u4_U73 (.A2( u2_u13_X_26 ) , .ZN( u2_u13_u4_n100 ) , .A1( u2_u13_u4_n177 ) );
  NOR2_X1 u2_u13_u4_U74 (.A2( u2_u13_X_28 ) , .A1( u2_u13_X_29 ) , .ZN( u2_u13_u4_n128 ) );
  NOR2_X1 u2_u13_u4_U75 (.A2( u2_u13_X_27 ) , .A1( u2_u13_X_30 ) , .ZN( u2_u13_u4_n102 ) );
  NOR2_X1 u2_u13_u4_U76 (.A2( u2_u13_X_25 ) , .A1( u2_u13_X_26 ) , .ZN( u2_u13_u4_n98 ) );
  AND2_X1 u2_u13_u4_U77 (.A2( u2_u13_X_25 ) , .A1( u2_u13_X_26 ) , .ZN( u2_u13_u4_n104 ) );
  AND2_X1 u2_u13_u4_U78 (.A1( u2_u13_X_30 ) , .A2( u2_u13_u4_n176 ) , .ZN( u2_u13_u4_n99 ) );
  AND2_X1 u2_u13_u4_U79 (.A1( u2_u13_X_26 ) , .ZN( u2_u13_u4_n101 ) , .A2( u2_u13_u4_n177 ) );
  INV_X1 u2_u13_u4_U8 (.A( u2_u13_u4_n113 ) , .ZN( u2_u13_u4_n185 ) );
  AND2_X1 u2_u13_u4_U80 (.A1( u2_u13_X_27 ) , .A2( u2_u13_X_30 ) , .ZN( u2_u13_u4_n103 ) );
  INV_X1 u2_u13_u4_U81 (.A( u2_u13_X_28 ) , .ZN( u2_u13_u4_n169 ) );
  INV_X1 u2_u13_u4_U82 (.A( u2_u13_X_29 ) , .ZN( u2_u13_u4_n168 ) );
  INV_X1 u2_u13_u4_U83 (.A( u2_u13_X_25 ) , .ZN( u2_u13_u4_n177 ) );
  INV_X1 u2_u13_u4_U84 (.A( u2_u13_X_27 ) , .ZN( u2_u13_u4_n176 ) );
  NAND4_X1 u2_u13_u4_U85 (.ZN( u2_out13_25 ) , .A4( u2_u13_u4_n139 ) , .A3( u2_u13_u4_n140 ) , .A2( u2_u13_u4_n141 ) , .A1( u2_u13_u4_n142 ) );
  OAI21_X1 u2_u13_u4_U86 (.A( u2_u13_u4_n128 ) , .B2( u2_u13_u4_n129 ) , .B1( u2_u13_u4_n130 ) , .ZN( u2_u13_u4_n142 ) );
  OAI21_X1 u2_u13_u4_U87 (.B2( u2_u13_u4_n131 ) , .ZN( u2_u13_u4_n141 ) , .A( u2_u13_u4_n175 ) , .B1( u2_u13_u4_n183 ) );
  NAND4_X1 u2_u13_u4_U88 (.ZN( u2_out13_14 ) , .A4( u2_u13_u4_n124 ) , .A3( u2_u13_u4_n125 ) , .A2( u2_u13_u4_n126 ) , .A1( u2_u13_u4_n127 ) );
  AOI22_X1 u2_u13_u4_U89 (.B2( u2_u13_u4_n117 ) , .ZN( u2_u13_u4_n126 ) , .A1( u2_u13_u4_n129 ) , .B1( u2_u13_u4_n152 ) , .A2( u2_u13_u4_n175 ) );
  NOR4_X1 u2_u13_u4_U9 (.A4( u2_u13_u4_n106 ) , .A3( u2_u13_u4_n107 ) , .A2( u2_u13_u4_n108 ) , .A1( u2_u13_u4_n109 ) , .ZN( u2_u13_u4_n110 ) );
  AOI22_X1 u2_u13_u4_U90 (.ZN( u2_u13_u4_n125 ) , .B2( u2_u13_u4_n131 ) , .A2( u2_u13_u4_n132 ) , .B1( u2_u13_u4_n138 ) , .A1( u2_u13_u4_n178 ) );
  NAND4_X1 u2_u13_u4_U91 (.ZN( u2_out13_8 ) , .A4( u2_u13_u4_n110 ) , .A3( u2_u13_u4_n111 ) , .A2( u2_u13_u4_n112 ) , .A1( u2_u13_u4_n186 ) );
  NAND2_X1 u2_u13_u4_U92 (.ZN( u2_u13_u4_n112 ) , .A2( u2_u13_u4_n130 ) , .A1( u2_u13_u4_n150 ) );
  AOI22_X1 u2_u13_u4_U93 (.ZN( u2_u13_u4_n111 ) , .B2( u2_u13_u4_n132 ) , .A1( u2_u13_u4_n152 ) , .B1( u2_u13_u4_n178 ) , .A2( u2_u13_u4_n97 ) );
  AOI22_X1 u2_u13_u4_U94 (.B2( u2_u13_u4_n149 ) , .B1( u2_u13_u4_n150 ) , .A2( u2_u13_u4_n151 ) , .A1( u2_u13_u4_n152 ) , .ZN( u2_u13_u4_n167 ) );
  NOR4_X1 u2_u13_u4_U95 (.A4( u2_u13_u4_n162 ) , .A3( u2_u13_u4_n163 ) , .A2( u2_u13_u4_n164 ) , .A1( u2_u13_u4_n165 ) , .ZN( u2_u13_u4_n166 ) );
  NAND3_X1 u2_u13_u4_U96 (.ZN( u2_out13_3 ) , .A3( u2_u13_u4_n166 ) , .A1( u2_u13_u4_n167 ) , .A2( u2_u13_u4_n186 ) );
  NAND3_X1 u2_u13_u4_U97 (.A3( u2_u13_u4_n146 ) , .A2( u2_u13_u4_n147 ) , .A1( u2_u13_u4_n148 ) , .ZN( u2_u13_u4_n149 ) );
  NAND3_X1 u2_u13_u4_U98 (.A3( u2_u13_u4_n143 ) , .A2( u2_u13_u4_n144 ) , .A1( u2_u13_u4_n145 ) , .ZN( u2_u13_u4_n151 ) );
  NAND3_X1 u2_u13_u4_U99 (.A3( u2_u13_u4_n121 ) , .ZN( u2_u13_u4_n122 ) , .A2( u2_u13_u4_n144 ) , .A1( u2_u13_u4_n154 ) );
  XOR2_X1 u2_u2_U10 (.B( u2_K3_45 ) , .A( u2_R1_30 ) , .Z( u2_u2_X_45 ) );
  XOR2_X1 u2_u2_U11 (.B( u2_K3_44 ) , .A( u2_R1_29 ) , .Z( u2_u2_X_44 ) );
  XOR2_X1 u2_u2_U12 (.B( u2_K3_43 ) , .A( u2_R1_28 ) , .Z( u2_u2_X_43 ) );
  XOR2_X1 u2_u2_U13 (.B( u2_K3_42 ) , .A( u2_R1_29 ) , .Z( u2_u2_X_42 ) );
  XOR2_X1 u2_u2_U14 (.B( u2_K3_41 ) , .A( u2_R1_28 ) , .Z( u2_u2_X_41 ) );
  XOR2_X1 u2_u2_U15 (.B( u2_K3_40 ) , .A( u2_R1_27 ) , .Z( u2_u2_X_40 ) );
  XOR2_X1 u2_u2_U17 (.B( u2_K3_39 ) , .A( u2_R1_26 ) , .Z( u2_u2_X_39 ) );
  XOR2_X1 u2_u2_U18 (.B( u2_K3_38 ) , .A( u2_R1_25 ) , .Z( u2_u2_X_38 ) );
  XOR2_X1 u2_u2_U19 (.B( u2_K3_37 ) , .A( u2_R1_24 ) , .Z( u2_u2_X_37 ) );
  XOR2_X1 u2_u2_U20 (.B( u2_K3_36 ) , .A( u2_R1_25 ) , .Z( u2_u2_X_36 ) );
  XOR2_X1 u2_u2_U21 (.B( u2_K3_35 ) , .A( u2_R1_24 ) , .Z( u2_u2_X_35 ) );
  XOR2_X1 u2_u2_U22 (.B( u2_K3_34 ) , .A( u2_R1_23 ) , .Z( u2_u2_X_34 ) );
  XOR2_X1 u2_u2_U23 (.B( u2_K3_33 ) , .A( u2_R1_22 ) , .Z( u2_u2_X_33 ) );
  XOR2_X1 u2_u2_U24 (.B( u2_K3_32 ) , .A( u2_R1_21 ) , .Z( u2_u2_X_32 ) );
  XOR2_X1 u2_u2_U25 (.B( u2_K3_31 ) , .A( u2_R1_20 ) , .Z( u2_u2_X_31 ) );
  XOR2_X1 u2_u2_U26 (.B( u2_K3_30 ) , .A( u2_R1_21 ) , .Z( u2_u2_X_30 ) );
  XOR2_X1 u2_u2_U28 (.B( u2_K3_29 ) , .A( u2_R1_20 ) , .Z( u2_u2_X_29 ) );
  XOR2_X1 u2_u2_U29 (.B( u2_K3_28 ) , .A( u2_R1_19 ) , .Z( u2_u2_X_28 ) );
  XOR2_X1 u2_u2_U30 (.B( u2_K3_27 ) , .A( u2_R1_18 ) , .Z( u2_u2_X_27 ) );
  XOR2_X1 u2_u2_U31 (.B( u2_K3_26 ) , .A( u2_R1_17 ) , .Z( u2_u2_X_26 ) );
  XOR2_X1 u2_u2_U32 (.B( u2_K3_25 ) , .A( u2_R1_16 ) , .Z( u2_u2_X_25 ) );
  XOR2_X1 u2_u2_U33 (.B( u2_K3_24 ) , .A( u2_R1_17 ) , .Z( u2_u2_X_24 ) );
  XOR2_X1 u2_u2_U34 (.B( u2_K3_23 ) , .A( u2_R1_16 ) , .Z( u2_u2_X_23 ) );
  XOR2_X1 u2_u2_U35 (.B( u2_K3_22 ) , .A( u2_R1_15 ) , .Z( u2_u2_X_22 ) );
  XOR2_X1 u2_u2_U36 (.B( u2_K3_21 ) , .A( u2_R1_14 ) , .Z( u2_u2_X_21 ) );
  XOR2_X1 u2_u2_U37 (.B( u2_K3_20 ) , .A( u2_R1_13 ) , .Z( u2_u2_X_20 ) );
  XOR2_X1 u2_u2_U39 (.B( u2_K3_19 ) , .A( u2_R1_12 ) , .Z( u2_u2_X_19 ) );
  XOR2_X1 u2_u2_U7 (.B( u2_K3_48 ) , .A( u2_R1_1 ) , .Z( u2_u2_X_48 ) );
  XOR2_X1 u2_u2_U8 (.B( u2_K3_47 ) , .A( u2_R1_32 ) , .Z( u2_u2_X_47 ) );
  XOR2_X1 u2_u2_U9 (.B( u2_K3_46 ) , .A( u2_R1_31 ) , .Z( u2_u2_X_46 ) );
  OAI22_X1 u2_u2_u3_U10 (.B1( u2_u2_u3_n113 ) , .A2( u2_u2_u3_n135 ) , .A1( u2_u2_u3_n150 ) , .B2( u2_u2_u3_n164 ) , .ZN( u2_u2_u3_n98 ) );
  OAI211_X1 u2_u2_u3_U11 (.B( u2_u2_u3_n106 ) , .ZN( u2_u2_u3_n119 ) , .C2( u2_u2_u3_n128 ) , .C1( u2_u2_u3_n167 ) , .A( u2_u2_u3_n181 ) );
  AOI221_X1 u2_u2_u3_U12 (.C1( u2_u2_u3_n105 ) , .ZN( u2_u2_u3_n106 ) , .A( u2_u2_u3_n131 ) , .B2( u2_u2_u3_n132 ) , .C2( u2_u2_u3_n133 ) , .B1( u2_u2_u3_n169 ) );
  INV_X1 u2_u2_u3_U13 (.ZN( u2_u2_u3_n181 ) , .A( u2_u2_u3_n98 ) );
  NAND2_X1 u2_u2_u3_U14 (.ZN( u2_u2_u3_n105 ) , .A2( u2_u2_u3_n130 ) , .A1( u2_u2_u3_n155 ) );
  AOI22_X1 u2_u2_u3_U15 (.B1( u2_u2_u3_n115 ) , .A2( u2_u2_u3_n116 ) , .ZN( u2_u2_u3_n123 ) , .B2( u2_u2_u3_n133 ) , .A1( u2_u2_u3_n169 ) );
  NAND2_X1 u2_u2_u3_U16 (.ZN( u2_u2_u3_n116 ) , .A2( u2_u2_u3_n151 ) , .A1( u2_u2_u3_n182 ) );
  NOR2_X1 u2_u2_u3_U17 (.ZN( u2_u2_u3_n126 ) , .A2( u2_u2_u3_n150 ) , .A1( u2_u2_u3_n164 ) );
  AOI21_X1 u2_u2_u3_U18 (.ZN( u2_u2_u3_n112 ) , .B2( u2_u2_u3_n146 ) , .B1( u2_u2_u3_n155 ) , .A( u2_u2_u3_n167 ) );
  NAND2_X1 u2_u2_u3_U19 (.A1( u2_u2_u3_n135 ) , .ZN( u2_u2_u3_n142 ) , .A2( u2_u2_u3_n164 ) );
  NAND2_X1 u2_u2_u3_U20 (.ZN( u2_u2_u3_n132 ) , .A2( u2_u2_u3_n152 ) , .A1( u2_u2_u3_n156 ) );
  AND2_X1 u2_u2_u3_U21 (.A2( u2_u2_u3_n113 ) , .A1( u2_u2_u3_n114 ) , .ZN( u2_u2_u3_n151 ) );
  INV_X1 u2_u2_u3_U22 (.A( u2_u2_u3_n133 ) , .ZN( u2_u2_u3_n165 ) );
  INV_X1 u2_u2_u3_U23 (.A( u2_u2_u3_n135 ) , .ZN( u2_u2_u3_n170 ) );
  NAND2_X1 u2_u2_u3_U24 (.A1( u2_u2_u3_n107 ) , .A2( u2_u2_u3_n108 ) , .ZN( u2_u2_u3_n140 ) );
  NAND2_X1 u2_u2_u3_U25 (.ZN( u2_u2_u3_n117 ) , .A1( u2_u2_u3_n124 ) , .A2( u2_u2_u3_n148 ) );
  NAND2_X1 u2_u2_u3_U26 (.ZN( u2_u2_u3_n143 ) , .A1( u2_u2_u3_n165 ) , .A2( u2_u2_u3_n167 ) );
  INV_X1 u2_u2_u3_U27 (.A( u2_u2_u3_n130 ) , .ZN( u2_u2_u3_n177 ) );
  INV_X1 u2_u2_u3_U28 (.A( u2_u2_u3_n128 ) , .ZN( u2_u2_u3_n176 ) );
  INV_X1 u2_u2_u3_U29 (.A( u2_u2_u3_n155 ) , .ZN( u2_u2_u3_n174 ) );
  INV_X1 u2_u2_u3_U3 (.A( u2_u2_u3_n129 ) , .ZN( u2_u2_u3_n183 ) );
  INV_X1 u2_u2_u3_U30 (.A( u2_u2_u3_n139 ) , .ZN( u2_u2_u3_n185 ) );
  NOR2_X1 u2_u2_u3_U31 (.ZN( u2_u2_u3_n135 ) , .A2( u2_u2_u3_n141 ) , .A1( u2_u2_u3_n169 ) );
  OAI222_X1 u2_u2_u3_U32 (.C2( u2_u2_u3_n107 ) , .A2( u2_u2_u3_n108 ) , .B1( u2_u2_u3_n135 ) , .ZN( u2_u2_u3_n138 ) , .B2( u2_u2_u3_n146 ) , .C1( u2_u2_u3_n154 ) , .A1( u2_u2_u3_n164 ) );
  NOR4_X1 u2_u2_u3_U33 (.A4( u2_u2_u3_n157 ) , .A3( u2_u2_u3_n158 ) , .A2( u2_u2_u3_n159 ) , .A1( u2_u2_u3_n160 ) , .ZN( u2_u2_u3_n161 ) );
  AOI21_X1 u2_u2_u3_U34 (.B2( u2_u2_u3_n152 ) , .B1( u2_u2_u3_n153 ) , .ZN( u2_u2_u3_n158 ) , .A( u2_u2_u3_n164 ) );
  AOI21_X1 u2_u2_u3_U35 (.A( u2_u2_u3_n154 ) , .B2( u2_u2_u3_n155 ) , .B1( u2_u2_u3_n156 ) , .ZN( u2_u2_u3_n157 ) );
  AOI21_X1 u2_u2_u3_U36 (.A( u2_u2_u3_n149 ) , .B2( u2_u2_u3_n150 ) , .B1( u2_u2_u3_n151 ) , .ZN( u2_u2_u3_n159 ) );
  AOI211_X1 u2_u2_u3_U37 (.ZN( u2_u2_u3_n109 ) , .A( u2_u2_u3_n119 ) , .C2( u2_u2_u3_n129 ) , .B( u2_u2_u3_n138 ) , .C1( u2_u2_u3_n141 ) );
  AOI211_X1 u2_u2_u3_U38 (.B( u2_u2_u3_n119 ) , .A( u2_u2_u3_n120 ) , .C2( u2_u2_u3_n121 ) , .ZN( u2_u2_u3_n122 ) , .C1( u2_u2_u3_n179 ) );
  INV_X1 u2_u2_u3_U39 (.A( u2_u2_u3_n156 ) , .ZN( u2_u2_u3_n179 ) );
  INV_X1 u2_u2_u3_U4 (.A( u2_u2_u3_n140 ) , .ZN( u2_u2_u3_n182 ) );
  OAI22_X1 u2_u2_u3_U40 (.B1( u2_u2_u3_n118 ) , .ZN( u2_u2_u3_n120 ) , .A1( u2_u2_u3_n135 ) , .B2( u2_u2_u3_n154 ) , .A2( u2_u2_u3_n178 ) );
  AND3_X1 u2_u2_u3_U41 (.ZN( u2_u2_u3_n118 ) , .A2( u2_u2_u3_n124 ) , .A1( u2_u2_u3_n144 ) , .A3( u2_u2_u3_n152 ) );
  INV_X1 u2_u2_u3_U42 (.A( u2_u2_u3_n121 ) , .ZN( u2_u2_u3_n164 ) );
  NAND2_X1 u2_u2_u3_U43 (.ZN( u2_u2_u3_n133 ) , .A1( u2_u2_u3_n154 ) , .A2( u2_u2_u3_n164 ) );
  OAI211_X1 u2_u2_u3_U44 (.B( u2_u2_u3_n127 ) , .ZN( u2_u2_u3_n139 ) , .C1( u2_u2_u3_n150 ) , .C2( u2_u2_u3_n154 ) , .A( u2_u2_u3_n184 ) );
  INV_X1 u2_u2_u3_U45 (.A( u2_u2_u3_n125 ) , .ZN( u2_u2_u3_n184 ) );
  AOI221_X1 u2_u2_u3_U46 (.A( u2_u2_u3_n126 ) , .ZN( u2_u2_u3_n127 ) , .C2( u2_u2_u3_n132 ) , .C1( u2_u2_u3_n169 ) , .B2( u2_u2_u3_n170 ) , .B1( u2_u2_u3_n174 ) );
  OAI22_X1 u2_u2_u3_U47 (.A1( u2_u2_u3_n124 ) , .ZN( u2_u2_u3_n125 ) , .B2( u2_u2_u3_n145 ) , .A2( u2_u2_u3_n165 ) , .B1( u2_u2_u3_n167 ) );
  NOR2_X1 u2_u2_u3_U48 (.A1( u2_u2_u3_n113 ) , .ZN( u2_u2_u3_n131 ) , .A2( u2_u2_u3_n154 ) );
  NAND2_X1 u2_u2_u3_U49 (.A1( u2_u2_u3_n103 ) , .ZN( u2_u2_u3_n150 ) , .A2( u2_u2_u3_n99 ) );
  INV_X1 u2_u2_u3_U5 (.A( u2_u2_u3_n117 ) , .ZN( u2_u2_u3_n178 ) );
  NAND2_X1 u2_u2_u3_U50 (.A2( u2_u2_u3_n102 ) , .ZN( u2_u2_u3_n155 ) , .A1( u2_u2_u3_n97 ) );
  INV_X1 u2_u2_u3_U51 (.A( u2_u2_u3_n141 ) , .ZN( u2_u2_u3_n167 ) );
  AOI21_X1 u2_u2_u3_U52 (.B2( u2_u2_u3_n114 ) , .B1( u2_u2_u3_n146 ) , .A( u2_u2_u3_n154 ) , .ZN( u2_u2_u3_n94 ) );
  AOI21_X1 u2_u2_u3_U53 (.ZN( u2_u2_u3_n110 ) , .B2( u2_u2_u3_n142 ) , .B1( u2_u2_u3_n186 ) , .A( u2_u2_u3_n95 ) );
  INV_X1 u2_u2_u3_U54 (.A( u2_u2_u3_n145 ) , .ZN( u2_u2_u3_n186 ) );
  AOI21_X1 u2_u2_u3_U55 (.B1( u2_u2_u3_n124 ) , .A( u2_u2_u3_n149 ) , .B2( u2_u2_u3_n155 ) , .ZN( u2_u2_u3_n95 ) );
  INV_X1 u2_u2_u3_U56 (.A( u2_u2_u3_n149 ) , .ZN( u2_u2_u3_n169 ) );
  NAND2_X1 u2_u2_u3_U57 (.ZN( u2_u2_u3_n124 ) , .A1( u2_u2_u3_n96 ) , .A2( u2_u2_u3_n97 ) );
  NAND2_X1 u2_u2_u3_U58 (.A2( u2_u2_u3_n100 ) , .ZN( u2_u2_u3_n146 ) , .A1( u2_u2_u3_n96 ) );
  NAND2_X1 u2_u2_u3_U59 (.A1( u2_u2_u3_n101 ) , .ZN( u2_u2_u3_n145 ) , .A2( u2_u2_u3_n99 ) );
  AOI221_X1 u2_u2_u3_U6 (.A( u2_u2_u3_n131 ) , .C2( u2_u2_u3_n132 ) , .C1( u2_u2_u3_n133 ) , .ZN( u2_u2_u3_n134 ) , .B1( u2_u2_u3_n143 ) , .B2( u2_u2_u3_n177 ) );
  NAND2_X1 u2_u2_u3_U60 (.A1( u2_u2_u3_n100 ) , .ZN( u2_u2_u3_n156 ) , .A2( u2_u2_u3_n99 ) );
  NAND2_X1 u2_u2_u3_U61 (.A2( u2_u2_u3_n101 ) , .A1( u2_u2_u3_n104 ) , .ZN( u2_u2_u3_n148 ) );
  NAND2_X1 u2_u2_u3_U62 (.A1( u2_u2_u3_n100 ) , .A2( u2_u2_u3_n102 ) , .ZN( u2_u2_u3_n128 ) );
  NAND2_X1 u2_u2_u3_U63 (.A2( u2_u2_u3_n101 ) , .A1( u2_u2_u3_n102 ) , .ZN( u2_u2_u3_n152 ) );
  NAND2_X1 u2_u2_u3_U64 (.A2( u2_u2_u3_n101 ) , .ZN( u2_u2_u3_n114 ) , .A1( u2_u2_u3_n96 ) );
  NAND2_X1 u2_u2_u3_U65 (.ZN( u2_u2_u3_n107 ) , .A1( u2_u2_u3_n97 ) , .A2( u2_u2_u3_n99 ) );
  NAND2_X1 u2_u2_u3_U66 (.A2( u2_u2_u3_n100 ) , .A1( u2_u2_u3_n104 ) , .ZN( u2_u2_u3_n113 ) );
  NAND2_X1 u2_u2_u3_U67 (.A1( u2_u2_u3_n104 ) , .ZN( u2_u2_u3_n153 ) , .A2( u2_u2_u3_n97 ) );
  NAND2_X1 u2_u2_u3_U68 (.A2( u2_u2_u3_n103 ) , .A1( u2_u2_u3_n104 ) , .ZN( u2_u2_u3_n130 ) );
  NAND2_X1 u2_u2_u3_U69 (.A2( u2_u2_u3_n103 ) , .ZN( u2_u2_u3_n144 ) , .A1( u2_u2_u3_n96 ) );
  OAI22_X1 u2_u2_u3_U7 (.B2( u2_u2_u3_n147 ) , .A2( u2_u2_u3_n148 ) , .ZN( u2_u2_u3_n160 ) , .B1( u2_u2_u3_n165 ) , .A1( u2_u2_u3_n168 ) );
  NAND2_X1 u2_u2_u3_U70 (.A1( u2_u2_u3_n102 ) , .A2( u2_u2_u3_n103 ) , .ZN( u2_u2_u3_n108 ) );
  NOR2_X1 u2_u2_u3_U71 (.A2( u2_u2_X_19 ) , .A1( u2_u2_X_20 ) , .ZN( u2_u2_u3_n99 ) );
  NOR2_X1 u2_u2_u3_U72 (.A2( u2_u2_X_21 ) , .A1( u2_u2_X_24 ) , .ZN( u2_u2_u3_n103 ) );
  NOR2_X1 u2_u2_u3_U73 (.A2( u2_u2_X_24 ) , .A1( u2_u2_u3_n171 ) , .ZN( u2_u2_u3_n97 ) );
  NOR2_X1 u2_u2_u3_U74 (.A2( u2_u2_X_23 ) , .ZN( u2_u2_u3_n141 ) , .A1( u2_u2_u3_n166 ) );
  NOR2_X1 u2_u2_u3_U75 (.A2( u2_u2_X_19 ) , .A1( u2_u2_u3_n172 ) , .ZN( u2_u2_u3_n96 ) );
  NAND2_X1 u2_u2_u3_U76 (.A1( u2_u2_X_22 ) , .A2( u2_u2_X_23 ) , .ZN( u2_u2_u3_n154 ) );
  NAND2_X1 u2_u2_u3_U77 (.A1( u2_u2_X_23 ) , .ZN( u2_u2_u3_n149 ) , .A2( u2_u2_u3_n166 ) );
  NOR2_X1 u2_u2_u3_U78 (.A2( u2_u2_X_22 ) , .A1( u2_u2_X_23 ) , .ZN( u2_u2_u3_n121 ) );
  AND2_X1 u2_u2_u3_U79 (.A1( u2_u2_X_24 ) , .ZN( u2_u2_u3_n101 ) , .A2( u2_u2_u3_n171 ) );
  AND3_X1 u2_u2_u3_U8 (.A3( u2_u2_u3_n144 ) , .A2( u2_u2_u3_n145 ) , .A1( u2_u2_u3_n146 ) , .ZN( u2_u2_u3_n147 ) );
  AND2_X1 u2_u2_u3_U80 (.A1( u2_u2_X_19 ) , .ZN( u2_u2_u3_n102 ) , .A2( u2_u2_u3_n172 ) );
  AND2_X1 u2_u2_u3_U81 (.A1( u2_u2_X_21 ) , .A2( u2_u2_X_24 ) , .ZN( u2_u2_u3_n100 ) );
  AND2_X1 u2_u2_u3_U82 (.A2( u2_u2_X_19 ) , .A1( u2_u2_X_20 ) , .ZN( u2_u2_u3_n104 ) );
  INV_X1 u2_u2_u3_U83 (.A( u2_u2_X_22 ) , .ZN( u2_u2_u3_n166 ) );
  INV_X1 u2_u2_u3_U84 (.A( u2_u2_X_21 ) , .ZN( u2_u2_u3_n171 ) );
  INV_X1 u2_u2_u3_U85 (.A( u2_u2_X_20 ) , .ZN( u2_u2_u3_n172 ) );
  OR4_X1 u2_u2_u3_U86 (.ZN( u2_out2_10 ) , .A4( u2_u2_u3_n136 ) , .A3( u2_u2_u3_n137 ) , .A1( u2_u2_u3_n138 ) , .A2( u2_u2_u3_n139 ) );
  OAI222_X1 u2_u2_u3_U87 (.C1( u2_u2_u3_n128 ) , .ZN( u2_u2_u3_n137 ) , .B1( u2_u2_u3_n148 ) , .A2( u2_u2_u3_n150 ) , .B2( u2_u2_u3_n154 ) , .C2( u2_u2_u3_n164 ) , .A1( u2_u2_u3_n167 ) );
  OAI221_X1 u2_u2_u3_U88 (.A( u2_u2_u3_n134 ) , .B2( u2_u2_u3_n135 ) , .ZN( u2_u2_u3_n136 ) , .C1( u2_u2_u3_n149 ) , .B1( u2_u2_u3_n151 ) , .C2( u2_u2_u3_n183 ) );
  NAND4_X1 u2_u2_u3_U89 (.ZN( u2_out2_26 ) , .A4( u2_u2_u3_n109 ) , .A3( u2_u2_u3_n110 ) , .A2( u2_u2_u3_n111 ) , .A1( u2_u2_u3_n173 ) );
  INV_X1 u2_u2_u3_U9 (.A( u2_u2_u3_n143 ) , .ZN( u2_u2_u3_n168 ) );
  INV_X1 u2_u2_u3_U90 (.ZN( u2_u2_u3_n173 ) , .A( u2_u2_u3_n94 ) );
  OAI21_X1 u2_u2_u3_U91 (.ZN( u2_u2_u3_n111 ) , .B2( u2_u2_u3_n117 ) , .A( u2_u2_u3_n133 ) , .B1( u2_u2_u3_n176 ) );
  NAND4_X1 u2_u2_u3_U92 (.ZN( u2_out2_20 ) , .A4( u2_u2_u3_n122 ) , .A3( u2_u2_u3_n123 ) , .A1( u2_u2_u3_n175 ) , .A2( u2_u2_u3_n180 ) );
  INV_X1 u2_u2_u3_U93 (.A( u2_u2_u3_n112 ) , .ZN( u2_u2_u3_n175 ) );
  INV_X1 u2_u2_u3_U94 (.A( u2_u2_u3_n126 ) , .ZN( u2_u2_u3_n180 ) );
  NAND4_X1 u2_u2_u3_U95 (.ZN( u2_out2_1 ) , .A4( u2_u2_u3_n161 ) , .A3( u2_u2_u3_n162 ) , .A2( u2_u2_u3_n163 ) , .A1( u2_u2_u3_n185 ) );
  NAND2_X1 u2_u2_u3_U96 (.ZN( u2_u2_u3_n163 ) , .A2( u2_u2_u3_n170 ) , .A1( u2_u2_u3_n176 ) );
  AOI22_X1 u2_u2_u3_U97 (.B2( u2_u2_u3_n140 ) , .B1( u2_u2_u3_n141 ) , .A2( u2_u2_u3_n142 ) , .ZN( u2_u2_u3_n162 ) , .A1( u2_u2_u3_n177 ) );
  NAND3_X1 u2_u2_u3_U98 (.A1( u2_u2_u3_n114 ) , .ZN( u2_u2_u3_n115 ) , .A2( u2_u2_u3_n145 ) , .A3( u2_u2_u3_n153 ) );
  NAND3_X1 u2_u2_u3_U99 (.ZN( u2_u2_u3_n129 ) , .A2( u2_u2_u3_n144 ) , .A1( u2_u2_u3_n153 ) , .A3( u2_u2_u3_n182 ) );
  OAI22_X1 u2_u2_u4_U10 (.B2( u2_u2_u4_n135 ) , .ZN( u2_u2_u4_n137 ) , .B1( u2_u2_u4_n153 ) , .A1( u2_u2_u4_n155 ) , .A2( u2_u2_u4_n171 ) );
  AND3_X1 u2_u2_u4_U11 (.A2( u2_u2_u4_n134 ) , .ZN( u2_u2_u4_n135 ) , .A3( u2_u2_u4_n145 ) , .A1( u2_u2_u4_n157 ) );
  NAND2_X1 u2_u2_u4_U12 (.ZN( u2_u2_u4_n132 ) , .A2( u2_u2_u4_n170 ) , .A1( u2_u2_u4_n173 ) );
  AOI21_X1 u2_u2_u4_U13 (.B2( u2_u2_u4_n160 ) , .B1( u2_u2_u4_n161 ) , .ZN( u2_u2_u4_n162 ) , .A( u2_u2_u4_n170 ) );
  AOI21_X1 u2_u2_u4_U14 (.ZN( u2_u2_u4_n107 ) , .B2( u2_u2_u4_n143 ) , .A( u2_u2_u4_n174 ) , .B1( u2_u2_u4_n184 ) );
  AOI21_X1 u2_u2_u4_U15 (.B2( u2_u2_u4_n158 ) , .B1( u2_u2_u4_n159 ) , .ZN( u2_u2_u4_n163 ) , .A( u2_u2_u4_n174 ) );
  AOI21_X1 u2_u2_u4_U16 (.A( u2_u2_u4_n153 ) , .B2( u2_u2_u4_n154 ) , .B1( u2_u2_u4_n155 ) , .ZN( u2_u2_u4_n165 ) );
  AOI21_X1 u2_u2_u4_U17 (.A( u2_u2_u4_n156 ) , .B2( u2_u2_u4_n157 ) , .ZN( u2_u2_u4_n164 ) , .B1( u2_u2_u4_n184 ) );
  INV_X1 u2_u2_u4_U18 (.A( u2_u2_u4_n138 ) , .ZN( u2_u2_u4_n170 ) );
  AND2_X1 u2_u2_u4_U19 (.A2( u2_u2_u4_n120 ) , .ZN( u2_u2_u4_n155 ) , .A1( u2_u2_u4_n160 ) );
  INV_X1 u2_u2_u4_U20 (.A( u2_u2_u4_n156 ) , .ZN( u2_u2_u4_n175 ) );
  NAND2_X1 u2_u2_u4_U21 (.A2( u2_u2_u4_n118 ) , .ZN( u2_u2_u4_n131 ) , .A1( u2_u2_u4_n147 ) );
  NAND2_X1 u2_u2_u4_U22 (.A1( u2_u2_u4_n119 ) , .A2( u2_u2_u4_n120 ) , .ZN( u2_u2_u4_n130 ) );
  NAND2_X1 u2_u2_u4_U23 (.ZN( u2_u2_u4_n117 ) , .A2( u2_u2_u4_n118 ) , .A1( u2_u2_u4_n148 ) );
  NAND2_X1 u2_u2_u4_U24 (.ZN( u2_u2_u4_n129 ) , .A1( u2_u2_u4_n134 ) , .A2( u2_u2_u4_n148 ) );
  AND3_X1 u2_u2_u4_U25 (.A1( u2_u2_u4_n119 ) , .A2( u2_u2_u4_n143 ) , .A3( u2_u2_u4_n154 ) , .ZN( u2_u2_u4_n161 ) );
  AND2_X1 u2_u2_u4_U26 (.A1( u2_u2_u4_n145 ) , .A2( u2_u2_u4_n147 ) , .ZN( u2_u2_u4_n159 ) );
  OR3_X1 u2_u2_u4_U27 (.A3( u2_u2_u4_n114 ) , .A2( u2_u2_u4_n115 ) , .A1( u2_u2_u4_n116 ) , .ZN( u2_u2_u4_n136 ) );
  AOI21_X1 u2_u2_u4_U28 (.A( u2_u2_u4_n113 ) , .ZN( u2_u2_u4_n116 ) , .B2( u2_u2_u4_n173 ) , .B1( u2_u2_u4_n174 ) );
  AOI21_X1 u2_u2_u4_U29 (.ZN( u2_u2_u4_n115 ) , .B2( u2_u2_u4_n145 ) , .B1( u2_u2_u4_n146 ) , .A( u2_u2_u4_n156 ) );
  NOR2_X1 u2_u2_u4_U3 (.ZN( u2_u2_u4_n121 ) , .A1( u2_u2_u4_n181 ) , .A2( u2_u2_u4_n182 ) );
  OAI22_X1 u2_u2_u4_U30 (.ZN( u2_u2_u4_n114 ) , .A2( u2_u2_u4_n121 ) , .B1( u2_u2_u4_n160 ) , .B2( u2_u2_u4_n170 ) , .A1( u2_u2_u4_n171 ) );
  INV_X1 u2_u2_u4_U31 (.A( u2_u2_u4_n158 ) , .ZN( u2_u2_u4_n182 ) );
  INV_X1 u2_u2_u4_U32 (.ZN( u2_u2_u4_n181 ) , .A( u2_u2_u4_n96 ) );
  INV_X1 u2_u2_u4_U33 (.A( u2_u2_u4_n144 ) , .ZN( u2_u2_u4_n179 ) );
  INV_X1 u2_u2_u4_U34 (.A( u2_u2_u4_n157 ) , .ZN( u2_u2_u4_n178 ) );
  NAND2_X1 u2_u2_u4_U35 (.A2( u2_u2_u4_n154 ) , .A1( u2_u2_u4_n96 ) , .ZN( u2_u2_u4_n97 ) );
  INV_X1 u2_u2_u4_U36 (.ZN( u2_u2_u4_n186 ) , .A( u2_u2_u4_n95 ) );
  OAI221_X1 u2_u2_u4_U37 (.C1( u2_u2_u4_n134 ) , .B1( u2_u2_u4_n158 ) , .B2( u2_u2_u4_n171 ) , .C2( u2_u2_u4_n173 ) , .A( u2_u2_u4_n94 ) , .ZN( u2_u2_u4_n95 ) );
  AOI222_X1 u2_u2_u4_U38 (.B2( u2_u2_u4_n132 ) , .A1( u2_u2_u4_n138 ) , .C2( u2_u2_u4_n175 ) , .A2( u2_u2_u4_n179 ) , .C1( u2_u2_u4_n181 ) , .B1( u2_u2_u4_n185 ) , .ZN( u2_u2_u4_n94 ) );
  INV_X1 u2_u2_u4_U39 (.A( u2_u2_u4_n113 ) , .ZN( u2_u2_u4_n185 ) );
  INV_X1 u2_u2_u4_U4 (.A( u2_u2_u4_n117 ) , .ZN( u2_u2_u4_n184 ) );
  INV_X1 u2_u2_u4_U40 (.A( u2_u2_u4_n143 ) , .ZN( u2_u2_u4_n183 ) );
  NOR2_X1 u2_u2_u4_U41 (.ZN( u2_u2_u4_n138 ) , .A1( u2_u2_u4_n168 ) , .A2( u2_u2_u4_n169 ) );
  NOR2_X1 u2_u2_u4_U42 (.A1( u2_u2_u4_n150 ) , .A2( u2_u2_u4_n152 ) , .ZN( u2_u2_u4_n153 ) );
  NOR2_X1 u2_u2_u4_U43 (.A2( u2_u2_u4_n128 ) , .A1( u2_u2_u4_n138 ) , .ZN( u2_u2_u4_n156 ) );
  AOI22_X1 u2_u2_u4_U44 (.B2( u2_u2_u4_n122 ) , .A1( u2_u2_u4_n123 ) , .ZN( u2_u2_u4_n124 ) , .B1( u2_u2_u4_n128 ) , .A2( u2_u2_u4_n172 ) );
  INV_X1 u2_u2_u4_U45 (.A( u2_u2_u4_n153 ) , .ZN( u2_u2_u4_n172 ) );
  NAND2_X1 u2_u2_u4_U46 (.A2( u2_u2_u4_n120 ) , .ZN( u2_u2_u4_n123 ) , .A1( u2_u2_u4_n161 ) );
  AOI22_X1 u2_u2_u4_U47 (.B2( u2_u2_u4_n132 ) , .A2( u2_u2_u4_n133 ) , .ZN( u2_u2_u4_n140 ) , .A1( u2_u2_u4_n150 ) , .B1( u2_u2_u4_n179 ) );
  NAND2_X1 u2_u2_u4_U48 (.ZN( u2_u2_u4_n133 ) , .A2( u2_u2_u4_n146 ) , .A1( u2_u2_u4_n154 ) );
  NAND2_X1 u2_u2_u4_U49 (.A1( u2_u2_u4_n103 ) , .ZN( u2_u2_u4_n154 ) , .A2( u2_u2_u4_n98 ) );
  NOR4_X1 u2_u2_u4_U5 (.A4( u2_u2_u4_n106 ) , .A3( u2_u2_u4_n107 ) , .A2( u2_u2_u4_n108 ) , .A1( u2_u2_u4_n109 ) , .ZN( u2_u2_u4_n110 ) );
  NAND2_X1 u2_u2_u4_U50 (.A1( u2_u2_u4_n101 ) , .ZN( u2_u2_u4_n158 ) , .A2( u2_u2_u4_n99 ) );
  AOI21_X1 u2_u2_u4_U51 (.ZN( u2_u2_u4_n127 ) , .A( u2_u2_u4_n136 ) , .B2( u2_u2_u4_n150 ) , .B1( u2_u2_u4_n180 ) );
  INV_X1 u2_u2_u4_U52 (.A( u2_u2_u4_n160 ) , .ZN( u2_u2_u4_n180 ) );
  NAND2_X1 u2_u2_u4_U53 (.A2( u2_u2_u4_n104 ) , .A1( u2_u2_u4_n105 ) , .ZN( u2_u2_u4_n146 ) );
  NAND2_X1 u2_u2_u4_U54 (.A2( u2_u2_u4_n101 ) , .A1( u2_u2_u4_n102 ) , .ZN( u2_u2_u4_n160 ) );
  NAND2_X1 u2_u2_u4_U55 (.ZN( u2_u2_u4_n134 ) , .A1( u2_u2_u4_n98 ) , .A2( u2_u2_u4_n99 ) );
  NAND2_X1 u2_u2_u4_U56 (.A1( u2_u2_u4_n103 ) , .A2( u2_u2_u4_n104 ) , .ZN( u2_u2_u4_n143 ) );
  NAND2_X1 u2_u2_u4_U57 (.A2( u2_u2_u4_n105 ) , .ZN( u2_u2_u4_n145 ) , .A1( u2_u2_u4_n98 ) );
  NAND2_X1 u2_u2_u4_U58 (.A1( u2_u2_u4_n100 ) , .A2( u2_u2_u4_n105 ) , .ZN( u2_u2_u4_n120 ) );
  NAND2_X1 u2_u2_u4_U59 (.A1( u2_u2_u4_n102 ) , .A2( u2_u2_u4_n104 ) , .ZN( u2_u2_u4_n148 ) );
  AOI21_X1 u2_u2_u4_U6 (.ZN( u2_u2_u4_n106 ) , .B2( u2_u2_u4_n146 ) , .B1( u2_u2_u4_n158 ) , .A( u2_u2_u4_n170 ) );
  NAND2_X1 u2_u2_u4_U60 (.A2( u2_u2_u4_n100 ) , .A1( u2_u2_u4_n103 ) , .ZN( u2_u2_u4_n157 ) );
  INV_X1 u2_u2_u4_U61 (.A( u2_u2_u4_n150 ) , .ZN( u2_u2_u4_n173 ) );
  INV_X1 u2_u2_u4_U62 (.A( u2_u2_u4_n152 ) , .ZN( u2_u2_u4_n171 ) );
  NAND2_X1 u2_u2_u4_U63 (.A1( u2_u2_u4_n100 ) , .ZN( u2_u2_u4_n118 ) , .A2( u2_u2_u4_n99 ) );
  NAND2_X1 u2_u2_u4_U64 (.A2( u2_u2_u4_n100 ) , .A1( u2_u2_u4_n102 ) , .ZN( u2_u2_u4_n144 ) );
  NAND2_X1 u2_u2_u4_U65 (.A2( u2_u2_u4_n101 ) , .A1( u2_u2_u4_n105 ) , .ZN( u2_u2_u4_n96 ) );
  INV_X1 u2_u2_u4_U66 (.A( u2_u2_u4_n128 ) , .ZN( u2_u2_u4_n174 ) );
  NAND2_X1 u2_u2_u4_U67 (.A2( u2_u2_u4_n102 ) , .ZN( u2_u2_u4_n119 ) , .A1( u2_u2_u4_n98 ) );
  NAND2_X1 u2_u2_u4_U68 (.A2( u2_u2_u4_n101 ) , .A1( u2_u2_u4_n103 ) , .ZN( u2_u2_u4_n147 ) );
  NAND2_X1 u2_u2_u4_U69 (.A2( u2_u2_u4_n104 ) , .ZN( u2_u2_u4_n113 ) , .A1( u2_u2_u4_n99 ) );
  AOI21_X1 u2_u2_u4_U7 (.ZN( u2_u2_u4_n108 ) , .B2( u2_u2_u4_n134 ) , .B1( u2_u2_u4_n155 ) , .A( u2_u2_u4_n156 ) );
  NOR2_X1 u2_u2_u4_U70 (.A2( u2_u2_X_28 ) , .ZN( u2_u2_u4_n150 ) , .A1( u2_u2_u4_n168 ) );
  NOR2_X1 u2_u2_u4_U71 (.A2( u2_u2_X_29 ) , .ZN( u2_u2_u4_n152 ) , .A1( u2_u2_u4_n169 ) );
  NOR2_X1 u2_u2_u4_U72 (.A2( u2_u2_X_30 ) , .ZN( u2_u2_u4_n105 ) , .A1( u2_u2_u4_n176 ) );
  NOR2_X1 u2_u2_u4_U73 (.A2( u2_u2_X_26 ) , .ZN( u2_u2_u4_n100 ) , .A1( u2_u2_u4_n177 ) );
  NOR2_X1 u2_u2_u4_U74 (.A2( u2_u2_X_28 ) , .A1( u2_u2_X_29 ) , .ZN( u2_u2_u4_n128 ) );
  NOR2_X1 u2_u2_u4_U75 (.A2( u2_u2_X_27 ) , .A1( u2_u2_X_30 ) , .ZN( u2_u2_u4_n102 ) );
  NOR2_X1 u2_u2_u4_U76 (.A2( u2_u2_X_25 ) , .A1( u2_u2_X_26 ) , .ZN( u2_u2_u4_n98 ) );
  AND2_X1 u2_u2_u4_U77 (.A2( u2_u2_X_25 ) , .A1( u2_u2_X_26 ) , .ZN( u2_u2_u4_n104 ) );
  AND2_X1 u2_u2_u4_U78 (.A1( u2_u2_X_30 ) , .A2( u2_u2_u4_n176 ) , .ZN( u2_u2_u4_n99 ) );
  AND2_X1 u2_u2_u4_U79 (.A1( u2_u2_X_26 ) , .ZN( u2_u2_u4_n101 ) , .A2( u2_u2_u4_n177 ) );
  AOI21_X1 u2_u2_u4_U8 (.ZN( u2_u2_u4_n109 ) , .A( u2_u2_u4_n153 ) , .B1( u2_u2_u4_n159 ) , .B2( u2_u2_u4_n184 ) );
  AND2_X1 u2_u2_u4_U80 (.A1( u2_u2_X_27 ) , .A2( u2_u2_X_30 ) , .ZN( u2_u2_u4_n103 ) );
  INV_X1 u2_u2_u4_U81 (.A( u2_u2_X_28 ) , .ZN( u2_u2_u4_n169 ) );
  INV_X1 u2_u2_u4_U82 (.A( u2_u2_X_29 ) , .ZN( u2_u2_u4_n168 ) );
  INV_X1 u2_u2_u4_U83 (.A( u2_u2_X_25 ) , .ZN( u2_u2_u4_n177 ) );
  INV_X1 u2_u2_u4_U84 (.A( u2_u2_X_27 ) , .ZN( u2_u2_u4_n176 ) );
  NAND4_X1 u2_u2_u4_U85 (.ZN( u2_out2_25 ) , .A4( u2_u2_u4_n139 ) , .A3( u2_u2_u4_n140 ) , .A2( u2_u2_u4_n141 ) , .A1( u2_u2_u4_n142 ) );
  OAI21_X1 u2_u2_u4_U86 (.A( u2_u2_u4_n128 ) , .B2( u2_u2_u4_n129 ) , .B1( u2_u2_u4_n130 ) , .ZN( u2_u2_u4_n142 ) );
  OAI21_X1 u2_u2_u4_U87 (.B2( u2_u2_u4_n131 ) , .ZN( u2_u2_u4_n141 ) , .A( u2_u2_u4_n175 ) , .B1( u2_u2_u4_n183 ) );
  NAND4_X1 u2_u2_u4_U88 (.ZN( u2_out2_14 ) , .A4( u2_u2_u4_n124 ) , .A3( u2_u2_u4_n125 ) , .A2( u2_u2_u4_n126 ) , .A1( u2_u2_u4_n127 ) );
  AOI22_X1 u2_u2_u4_U89 (.B2( u2_u2_u4_n117 ) , .ZN( u2_u2_u4_n126 ) , .A1( u2_u2_u4_n129 ) , .B1( u2_u2_u4_n152 ) , .A2( u2_u2_u4_n175 ) );
  AOI211_X1 u2_u2_u4_U9 (.B( u2_u2_u4_n136 ) , .A( u2_u2_u4_n137 ) , .C2( u2_u2_u4_n138 ) , .ZN( u2_u2_u4_n139 ) , .C1( u2_u2_u4_n182 ) );
  AOI22_X1 u2_u2_u4_U90 (.ZN( u2_u2_u4_n125 ) , .B2( u2_u2_u4_n131 ) , .A2( u2_u2_u4_n132 ) , .B1( u2_u2_u4_n138 ) , .A1( u2_u2_u4_n178 ) );
  NAND4_X1 u2_u2_u4_U91 (.ZN( u2_out2_8 ) , .A4( u2_u2_u4_n110 ) , .A3( u2_u2_u4_n111 ) , .A2( u2_u2_u4_n112 ) , .A1( u2_u2_u4_n186 ) );
  NAND2_X1 u2_u2_u4_U92 (.ZN( u2_u2_u4_n112 ) , .A2( u2_u2_u4_n130 ) , .A1( u2_u2_u4_n150 ) );
  AOI22_X1 u2_u2_u4_U93 (.ZN( u2_u2_u4_n111 ) , .B2( u2_u2_u4_n132 ) , .A1( u2_u2_u4_n152 ) , .B1( u2_u2_u4_n178 ) , .A2( u2_u2_u4_n97 ) );
  AOI22_X1 u2_u2_u4_U94 (.B2( u2_u2_u4_n149 ) , .B1( u2_u2_u4_n150 ) , .A2( u2_u2_u4_n151 ) , .A1( u2_u2_u4_n152 ) , .ZN( u2_u2_u4_n167 ) );
  NOR4_X1 u2_u2_u4_U95 (.A4( u2_u2_u4_n162 ) , .A3( u2_u2_u4_n163 ) , .A2( u2_u2_u4_n164 ) , .A1( u2_u2_u4_n165 ) , .ZN( u2_u2_u4_n166 ) );
  NAND3_X1 u2_u2_u4_U96 (.ZN( u2_out2_3 ) , .A3( u2_u2_u4_n166 ) , .A1( u2_u2_u4_n167 ) , .A2( u2_u2_u4_n186 ) );
  NAND3_X1 u2_u2_u4_U97 (.A3( u2_u2_u4_n146 ) , .A2( u2_u2_u4_n147 ) , .A1( u2_u2_u4_n148 ) , .ZN( u2_u2_u4_n149 ) );
  NAND3_X1 u2_u2_u4_U98 (.A3( u2_u2_u4_n143 ) , .A2( u2_u2_u4_n144 ) , .A1( u2_u2_u4_n145 ) , .ZN( u2_u2_u4_n151 ) );
  NAND3_X1 u2_u2_u4_U99 (.A3( u2_u2_u4_n121 ) , .ZN( u2_u2_u4_n122 ) , .A2( u2_u2_u4_n144 ) , .A1( u2_u2_u4_n154 ) );
  INV_X1 u2_u2_u5_U10 (.A( u2_u2_u5_n121 ) , .ZN( u2_u2_u5_n177 ) );
  NOR3_X1 u2_u2_u5_U100 (.A3( u2_u2_u5_n141 ) , .A1( u2_u2_u5_n142 ) , .ZN( u2_u2_u5_n143 ) , .A2( u2_u2_u5_n191 ) );
  NAND4_X1 u2_u2_u5_U101 (.ZN( u2_out2_4 ) , .A4( u2_u2_u5_n112 ) , .A2( u2_u2_u5_n113 ) , .A1( u2_u2_u5_n114 ) , .A3( u2_u2_u5_n195 ) );
  AOI211_X1 u2_u2_u5_U102 (.A( u2_u2_u5_n110 ) , .C1( u2_u2_u5_n111 ) , .ZN( u2_u2_u5_n112 ) , .B( u2_u2_u5_n118 ) , .C2( u2_u2_u5_n177 ) );
  AOI222_X1 u2_u2_u5_U103 (.ZN( u2_u2_u5_n113 ) , .A1( u2_u2_u5_n131 ) , .C1( u2_u2_u5_n148 ) , .B2( u2_u2_u5_n174 ) , .C2( u2_u2_u5_n178 ) , .A2( u2_u2_u5_n179 ) , .B1( u2_u2_u5_n99 ) );
  NAND3_X1 u2_u2_u5_U104 (.A2( u2_u2_u5_n154 ) , .A3( u2_u2_u5_n158 ) , .A1( u2_u2_u5_n161 ) , .ZN( u2_u2_u5_n99 ) );
  NOR2_X1 u2_u2_u5_U11 (.ZN( u2_u2_u5_n160 ) , .A2( u2_u2_u5_n173 ) , .A1( u2_u2_u5_n177 ) );
  INV_X1 u2_u2_u5_U12 (.A( u2_u2_u5_n150 ) , .ZN( u2_u2_u5_n174 ) );
  AOI21_X1 u2_u2_u5_U13 (.A( u2_u2_u5_n160 ) , .B2( u2_u2_u5_n161 ) , .ZN( u2_u2_u5_n162 ) , .B1( u2_u2_u5_n192 ) );
  INV_X1 u2_u2_u5_U14 (.A( u2_u2_u5_n159 ) , .ZN( u2_u2_u5_n192 ) );
  AOI21_X1 u2_u2_u5_U15 (.A( u2_u2_u5_n156 ) , .B2( u2_u2_u5_n157 ) , .B1( u2_u2_u5_n158 ) , .ZN( u2_u2_u5_n163 ) );
  AOI21_X1 u2_u2_u5_U16 (.B2( u2_u2_u5_n139 ) , .B1( u2_u2_u5_n140 ) , .ZN( u2_u2_u5_n141 ) , .A( u2_u2_u5_n150 ) );
  OAI21_X1 u2_u2_u5_U17 (.A( u2_u2_u5_n133 ) , .B2( u2_u2_u5_n134 ) , .B1( u2_u2_u5_n135 ) , .ZN( u2_u2_u5_n142 ) );
  OAI21_X1 u2_u2_u5_U18 (.ZN( u2_u2_u5_n133 ) , .B2( u2_u2_u5_n147 ) , .A( u2_u2_u5_n173 ) , .B1( u2_u2_u5_n188 ) );
  NAND2_X1 u2_u2_u5_U19 (.A2( u2_u2_u5_n119 ) , .A1( u2_u2_u5_n123 ) , .ZN( u2_u2_u5_n137 ) );
  INV_X1 u2_u2_u5_U20 (.A( u2_u2_u5_n155 ) , .ZN( u2_u2_u5_n194 ) );
  NAND2_X1 u2_u2_u5_U21 (.A1( u2_u2_u5_n121 ) , .ZN( u2_u2_u5_n132 ) , .A2( u2_u2_u5_n172 ) );
  NAND2_X1 u2_u2_u5_U22 (.A2( u2_u2_u5_n122 ) , .ZN( u2_u2_u5_n136 ) , .A1( u2_u2_u5_n154 ) );
  NAND2_X1 u2_u2_u5_U23 (.A2( u2_u2_u5_n119 ) , .A1( u2_u2_u5_n120 ) , .ZN( u2_u2_u5_n159 ) );
  INV_X1 u2_u2_u5_U24 (.A( u2_u2_u5_n156 ) , .ZN( u2_u2_u5_n175 ) );
  INV_X1 u2_u2_u5_U25 (.A( u2_u2_u5_n158 ) , .ZN( u2_u2_u5_n188 ) );
  INV_X1 u2_u2_u5_U26 (.A( u2_u2_u5_n152 ) , .ZN( u2_u2_u5_n179 ) );
  INV_X1 u2_u2_u5_U27 (.A( u2_u2_u5_n140 ) , .ZN( u2_u2_u5_n182 ) );
  INV_X1 u2_u2_u5_U28 (.A( u2_u2_u5_n151 ) , .ZN( u2_u2_u5_n183 ) );
  INV_X1 u2_u2_u5_U29 (.A( u2_u2_u5_n123 ) , .ZN( u2_u2_u5_n185 ) );
  NOR2_X1 u2_u2_u5_U3 (.ZN( u2_u2_u5_n134 ) , .A1( u2_u2_u5_n183 ) , .A2( u2_u2_u5_n190 ) );
  INV_X1 u2_u2_u5_U30 (.A( u2_u2_u5_n161 ) , .ZN( u2_u2_u5_n184 ) );
  INV_X1 u2_u2_u5_U31 (.A( u2_u2_u5_n139 ) , .ZN( u2_u2_u5_n189 ) );
  INV_X1 u2_u2_u5_U32 (.A( u2_u2_u5_n157 ) , .ZN( u2_u2_u5_n190 ) );
  INV_X1 u2_u2_u5_U33 (.A( u2_u2_u5_n120 ) , .ZN( u2_u2_u5_n193 ) );
  NAND2_X1 u2_u2_u5_U34 (.ZN( u2_u2_u5_n111 ) , .A1( u2_u2_u5_n140 ) , .A2( u2_u2_u5_n155 ) );
  INV_X1 u2_u2_u5_U35 (.A( u2_u2_u5_n117 ) , .ZN( u2_u2_u5_n196 ) );
  OAI221_X1 u2_u2_u5_U36 (.A( u2_u2_u5_n116 ) , .ZN( u2_u2_u5_n117 ) , .B2( u2_u2_u5_n119 ) , .C1( u2_u2_u5_n153 ) , .C2( u2_u2_u5_n158 ) , .B1( u2_u2_u5_n172 ) );
  AOI222_X1 u2_u2_u5_U37 (.ZN( u2_u2_u5_n116 ) , .B2( u2_u2_u5_n145 ) , .C1( u2_u2_u5_n148 ) , .A2( u2_u2_u5_n174 ) , .C2( u2_u2_u5_n177 ) , .B1( u2_u2_u5_n187 ) , .A1( u2_u2_u5_n193 ) );
  INV_X1 u2_u2_u5_U38 (.A( u2_u2_u5_n115 ) , .ZN( u2_u2_u5_n187 ) );
  NOR2_X1 u2_u2_u5_U39 (.ZN( u2_u2_u5_n100 ) , .A1( u2_u2_u5_n170 ) , .A2( u2_u2_u5_n180 ) );
  INV_X1 u2_u2_u5_U4 (.A( u2_u2_u5_n138 ) , .ZN( u2_u2_u5_n191 ) );
  AOI22_X1 u2_u2_u5_U40 (.B2( u2_u2_u5_n131 ) , .A2( u2_u2_u5_n146 ) , .ZN( u2_u2_u5_n169 ) , .B1( u2_u2_u5_n174 ) , .A1( u2_u2_u5_n185 ) );
  NOR2_X1 u2_u2_u5_U41 (.A1( u2_u2_u5_n146 ) , .ZN( u2_u2_u5_n150 ) , .A2( u2_u2_u5_n173 ) );
  AOI21_X1 u2_u2_u5_U42 (.A( u2_u2_u5_n118 ) , .B2( u2_u2_u5_n145 ) , .ZN( u2_u2_u5_n168 ) , .B1( u2_u2_u5_n186 ) );
  INV_X1 u2_u2_u5_U43 (.A( u2_u2_u5_n122 ) , .ZN( u2_u2_u5_n186 ) );
  NOR2_X1 u2_u2_u5_U44 (.A1( u2_u2_u5_n146 ) , .ZN( u2_u2_u5_n152 ) , .A2( u2_u2_u5_n176 ) );
  NOR2_X1 u2_u2_u5_U45 (.A1( u2_u2_u5_n115 ) , .ZN( u2_u2_u5_n118 ) , .A2( u2_u2_u5_n153 ) );
  NOR2_X1 u2_u2_u5_U46 (.A2( u2_u2_u5_n145 ) , .ZN( u2_u2_u5_n156 ) , .A1( u2_u2_u5_n174 ) );
  NOR2_X1 u2_u2_u5_U47 (.ZN( u2_u2_u5_n121 ) , .A2( u2_u2_u5_n145 ) , .A1( u2_u2_u5_n176 ) );
  AOI22_X1 u2_u2_u5_U48 (.ZN( u2_u2_u5_n114 ) , .A2( u2_u2_u5_n137 ) , .A1( u2_u2_u5_n145 ) , .B2( u2_u2_u5_n175 ) , .B1( u2_u2_u5_n193 ) );
  AOI21_X1 u2_u2_u5_U49 (.A( u2_u2_u5_n153 ) , .B2( u2_u2_u5_n154 ) , .B1( u2_u2_u5_n155 ) , .ZN( u2_u2_u5_n164 ) );
  OAI21_X1 u2_u2_u5_U5 (.B2( u2_u2_u5_n136 ) , .B1( u2_u2_u5_n137 ) , .ZN( u2_u2_u5_n138 ) , .A( u2_u2_u5_n177 ) );
  AOI21_X1 u2_u2_u5_U50 (.ZN( u2_u2_u5_n110 ) , .B1( u2_u2_u5_n122 ) , .B2( u2_u2_u5_n139 ) , .A( u2_u2_u5_n153 ) );
  INV_X1 u2_u2_u5_U51 (.A( u2_u2_u5_n153 ) , .ZN( u2_u2_u5_n176 ) );
  INV_X1 u2_u2_u5_U52 (.A( u2_u2_u5_n126 ) , .ZN( u2_u2_u5_n173 ) );
  AND2_X1 u2_u2_u5_U53 (.A2( u2_u2_u5_n104 ) , .A1( u2_u2_u5_n107 ) , .ZN( u2_u2_u5_n147 ) );
  AND2_X1 u2_u2_u5_U54 (.A2( u2_u2_u5_n104 ) , .A1( u2_u2_u5_n108 ) , .ZN( u2_u2_u5_n148 ) );
  NAND2_X1 u2_u2_u5_U55 (.A1( u2_u2_u5_n105 ) , .A2( u2_u2_u5_n106 ) , .ZN( u2_u2_u5_n158 ) );
  NAND2_X1 u2_u2_u5_U56 (.A2( u2_u2_u5_n108 ) , .A1( u2_u2_u5_n109 ) , .ZN( u2_u2_u5_n139 ) );
  NAND2_X1 u2_u2_u5_U57 (.A1( u2_u2_u5_n106 ) , .A2( u2_u2_u5_n108 ) , .ZN( u2_u2_u5_n119 ) );
  OAI211_X1 u2_u2_u5_U58 (.B( u2_u2_u5_n124 ) , .A( u2_u2_u5_n125 ) , .C2( u2_u2_u5_n126 ) , .C1( u2_u2_u5_n127 ) , .ZN( u2_u2_u5_n128 ) );
  NOR3_X1 u2_u2_u5_U59 (.ZN( u2_u2_u5_n127 ) , .A1( u2_u2_u5_n136 ) , .A3( u2_u2_u5_n148 ) , .A2( u2_u2_u5_n182 ) );
  INV_X1 u2_u2_u5_U6 (.A( u2_u2_u5_n135 ) , .ZN( u2_u2_u5_n178 ) );
  OAI21_X1 u2_u2_u5_U60 (.ZN( u2_u2_u5_n124 ) , .A( u2_u2_u5_n177 ) , .B2( u2_u2_u5_n183 ) , .B1( u2_u2_u5_n189 ) );
  OAI21_X1 u2_u2_u5_U61 (.ZN( u2_u2_u5_n125 ) , .A( u2_u2_u5_n174 ) , .B2( u2_u2_u5_n185 ) , .B1( u2_u2_u5_n190 ) );
  NAND2_X1 u2_u2_u5_U62 (.A2( u2_u2_u5_n103 ) , .A1( u2_u2_u5_n105 ) , .ZN( u2_u2_u5_n140 ) );
  NAND2_X1 u2_u2_u5_U63 (.A2( u2_u2_u5_n104 ) , .A1( u2_u2_u5_n105 ) , .ZN( u2_u2_u5_n155 ) );
  NAND2_X1 u2_u2_u5_U64 (.A2( u2_u2_u5_n106 ) , .A1( u2_u2_u5_n107 ) , .ZN( u2_u2_u5_n122 ) );
  NAND2_X1 u2_u2_u5_U65 (.A2( u2_u2_u5_n100 ) , .A1( u2_u2_u5_n106 ) , .ZN( u2_u2_u5_n115 ) );
  NAND2_X1 u2_u2_u5_U66 (.A2( u2_u2_u5_n100 ) , .A1( u2_u2_u5_n103 ) , .ZN( u2_u2_u5_n161 ) );
  NAND2_X1 u2_u2_u5_U67 (.A1( u2_u2_u5_n105 ) , .A2( u2_u2_u5_n109 ) , .ZN( u2_u2_u5_n154 ) );
  INV_X1 u2_u2_u5_U68 (.A( u2_u2_u5_n146 ) , .ZN( u2_u2_u5_n172 ) );
  NAND2_X1 u2_u2_u5_U69 (.A1( u2_u2_u5_n103 ) , .A2( u2_u2_u5_n108 ) , .ZN( u2_u2_u5_n123 ) );
  OAI22_X1 u2_u2_u5_U7 (.B2( u2_u2_u5_n149 ) , .B1( u2_u2_u5_n150 ) , .A2( u2_u2_u5_n151 ) , .A1( u2_u2_u5_n152 ) , .ZN( u2_u2_u5_n165 ) );
  NAND2_X1 u2_u2_u5_U70 (.A2( u2_u2_u5_n103 ) , .A1( u2_u2_u5_n107 ) , .ZN( u2_u2_u5_n151 ) );
  NAND2_X1 u2_u2_u5_U71 (.A2( u2_u2_u5_n107 ) , .A1( u2_u2_u5_n109 ) , .ZN( u2_u2_u5_n120 ) );
  NAND2_X1 u2_u2_u5_U72 (.A2( u2_u2_u5_n100 ) , .A1( u2_u2_u5_n109 ) , .ZN( u2_u2_u5_n157 ) );
  AND2_X1 u2_u2_u5_U73 (.A2( u2_u2_u5_n100 ) , .A1( u2_u2_u5_n104 ) , .ZN( u2_u2_u5_n131 ) );
  INV_X1 u2_u2_u5_U74 (.A( u2_u2_u5_n102 ) , .ZN( u2_u2_u5_n195 ) );
  OAI221_X1 u2_u2_u5_U75 (.A( u2_u2_u5_n101 ) , .ZN( u2_u2_u5_n102 ) , .C2( u2_u2_u5_n115 ) , .C1( u2_u2_u5_n126 ) , .B1( u2_u2_u5_n134 ) , .B2( u2_u2_u5_n160 ) );
  OAI21_X1 u2_u2_u5_U76 (.ZN( u2_u2_u5_n101 ) , .B1( u2_u2_u5_n137 ) , .A( u2_u2_u5_n146 ) , .B2( u2_u2_u5_n147 ) );
  NOR2_X1 u2_u2_u5_U77 (.A2( u2_u2_X_34 ) , .A1( u2_u2_X_35 ) , .ZN( u2_u2_u5_n145 ) );
  NOR2_X1 u2_u2_u5_U78 (.A2( u2_u2_X_34 ) , .ZN( u2_u2_u5_n146 ) , .A1( u2_u2_u5_n171 ) );
  NOR2_X1 u2_u2_u5_U79 (.A2( u2_u2_X_31 ) , .A1( u2_u2_X_32 ) , .ZN( u2_u2_u5_n103 ) );
  NOR3_X1 u2_u2_u5_U8 (.A2( u2_u2_u5_n147 ) , .A1( u2_u2_u5_n148 ) , .ZN( u2_u2_u5_n149 ) , .A3( u2_u2_u5_n194 ) );
  NOR2_X1 u2_u2_u5_U80 (.A2( u2_u2_X_36 ) , .ZN( u2_u2_u5_n105 ) , .A1( u2_u2_u5_n180 ) );
  NOR2_X1 u2_u2_u5_U81 (.A2( u2_u2_X_33 ) , .ZN( u2_u2_u5_n108 ) , .A1( u2_u2_u5_n170 ) );
  NOR2_X1 u2_u2_u5_U82 (.A2( u2_u2_X_33 ) , .A1( u2_u2_X_36 ) , .ZN( u2_u2_u5_n107 ) );
  NOR2_X1 u2_u2_u5_U83 (.A2( u2_u2_X_31 ) , .ZN( u2_u2_u5_n104 ) , .A1( u2_u2_u5_n181 ) );
  NAND2_X1 u2_u2_u5_U84 (.A2( u2_u2_X_34 ) , .A1( u2_u2_X_35 ) , .ZN( u2_u2_u5_n153 ) );
  NAND2_X1 u2_u2_u5_U85 (.A1( u2_u2_X_34 ) , .ZN( u2_u2_u5_n126 ) , .A2( u2_u2_u5_n171 ) );
  AND2_X1 u2_u2_u5_U86 (.A1( u2_u2_X_31 ) , .A2( u2_u2_X_32 ) , .ZN( u2_u2_u5_n106 ) );
  AND2_X1 u2_u2_u5_U87 (.A1( u2_u2_X_31 ) , .ZN( u2_u2_u5_n109 ) , .A2( u2_u2_u5_n181 ) );
  INV_X1 u2_u2_u5_U88 (.A( u2_u2_X_33 ) , .ZN( u2_u2_u5_n180 ) );
  INV_X1 u2_u2_u5_U89 (.A( u2_u2_X_35 ) , .ZN( u2_u2_u5_n171 ) );
  NOR2_X1 u2_u2_u5_U9 (.ZN( u2_u2_u5_n135 ) , .A1( u2_u2_u5_n173 ) , .A2( u2_u2_u5_n176 ) );
  INV_X1 u2_u2_u5_U90 (.A( u2_u2_X_36 ) , .ZN( u2_u2_u5_n170 ) );
  INV_X1 u2_u2_u5_U91 (.A( u2_u2_X_32 ) , .ZN( u2_u2_u5_n181 ) );
  NAND4_X1 u2_u2_u5_U92 (.ZN( u2_out2_29 ) , .A4( u2_u2_u5_n129 ) , .A3( u2_u2_u5_n130 ) , .A2( u2_u2_u5_n168 ) , .A1( u2_u2_u5_n196 ) );
  AOI221_X1 u2_u2_u5_U93 (.A( u2_u2_u5_n128 ) , .ZN( u2_u2_u5_n129 ) , .C2( u2_u2_u5_n132 ) , .B2( u2_u2_u5_n159 ) , .B1( u2_u2_u5_n176 ) , .C1( u2_u2_u5_n184 ) );
  AOI222_X1 u2_u2_u5_U94 (.ZN( u2_u2_u5_n130 ) , .A2( u2_u2_u5_n146 ) , .B1( u2_u2_u5_n147 ) , .C2( u2_u2_u5_n175 ) , .B2( u2_u2_u5_n179 ) , .A1( u2_u2_u5_n188 ) , .C1( u2_u2_u5_n194 ) );
  NAND4_X1 u2_u2_u5_U95 (.ZN( u2_out2_19 ) , .A4( u2_u2_u5_n166 ) , .A3( u2_u2_u5_n167 ) , .A2( u2_u2_u5_n168 ) , .A1( u2_u2_u5_n169 ) );
  AOI22_X1 u2_u2_u5_U96 (.B2( u2_u2_u5_n145 ) , .A2( u2_u2_u5_n146 ) , .ZN( u2_u2_u5_n167 ) , .B1( u2_u2_u5_n182 ) , .A1( u2_u2_u5_n189 ) );
  NOR4_X1 u2_u2_u5_U97 (.A4( u2_u2_u5_n162 ) , .A3( u2_u2_u5_n163 ) , .A2( u2_u2_u5_n164 ) , .A1( u2_u2_u5_n165 ) , .ZN( u2_u2_u5_n166 ) );
  NAND4_X1 u2_u2_u5_U98 (.ZN( u2_out2_11 ) , .A4( u2_u2_u5_n143 ) , .A3( u2_u2_u5_n144 ) , .A2( u2_u2_u5_n169 ) , .A1( u2_u2_u5_n196 ) );
  AOI22_X1 u2_u2_u5_U99 (.A2( u2_u2_u5_n132 ) , .ZN( u2_u2_u5_n144 ) , .B2( u2_u2_u5_n145 ) , .B1( u2_u2_u5_n184 ) , .A1( u2_u2_u5_n194 ) );
  OAI21_X1 u2_u2_u6_U10 (.A( u2_u2_u6_n159 ) , .B1( u2_u2_u6_n169 ) , .B2( u2_u2_u6_n173 ) , .ZN( u2_u2_u6_n90 ) );
  INV_X1 u2_u2_u6_U11 (.ZN( u2_u2_u6_n172 ) , .A( u2_u2_u6_n88 ) );
  AOI22_X1 u2_u2_u6_U12 (.A2( u2_u2_u6_n151 ) , .B2( u2_u2_u6_n161 ) , .A1( u2_u2_u6_n167 ) , .B1( u2_u2_u6_n170 ) , .ZN( u2_u2_u6_n89 ) );
  AOI21_X1 u2_u2_u6_U13 (.ZN( u2_u2_u6_n106 ) , .A( u2_u2_u6_n142 ) , .B2( u2_u2_u6_n159 ) , .B1( u2_u2_u6_n164 ) );
  INV_X1 u2_u2_u6_U14 (.A( u2_u2_u6_n155 ) , .ZN( u2_u2_u6_n161 ) );
  INV_X1 u2_u2_u6_U15 (.A( u2_u2_u6_n128 ) , .ZN( u2_u2_u6_n164 ) );
  NAND2_X1 u2_u2_u6_U16 (.ZN( u2_u2_u6_n110 ) , .A1( u2_u2_u6_n122 ) , .A2( u2_u2_u6_n129 ) );
  NAND2_X1 u2_u2_u6_U17 (.ZN( u2_u2_u6_n124 ) , .A2( u2_u2_u6_n146 ) , .A1( u2_u2_u6_n148 ) );
  INV_X1 u2_u2_u6_U18 (.A( u2_u2_u6_n132 ) , .ZN( u2_u2_u6_n171 ) );
  AND2_X1 u2_u2_u6_U19 (.A1( u2_u2_u6_n100 ) , .ZN( u2_u2_u6_n130 ) , .A2( u2_u2_u6_n147 ) );
  INV_X1 u2_u2_u6_U20 (.A( u2_u2_u6_n127 ) , .ZN( u2_u2_u6_n173 ) );
  INV_X1 u2_u2_u6_U21 (.A( u2_u2_u6_n121 ) , .ZN( u2_u2_u6_n167 ) );
  INV_X1 u2_u2_u6_U22 (.A( u2_u2_u6_n100 ) , .ZN( u2_u2_u6_n169 ) );
  INV_X1 u2_u2_u6_U23 (.A( u2_u2_u6_n123 ) , .ZN( u2_u2_u6_n170 ) );
  INV_X1 u2_u2_u6_U24 (.A( u2_u2_u6_n113 ) , .ZN( u2_u2_u6_n168 ) );
  AND2_X1 u2_u2_u6_U25 (.A1( u2_u2_u6_n107 ) , .A2( u2_u2_u6_n119 ) , .ZN( u2_u2_u6_n133 ) );
  AND2_X1 u2_u2_u6_U26 (.A2( u2_u2_u6_n121 ) , .A1( u2_u2_u6_n122 ) , .ZN( u2_u2_u6_n131 ) );
  AND3_X1 u2_u2_u6_U27 (.ZN( u2_u2_u6_n120 ) , .A2( u2_u2_u6_n127 ) , .A1( u2_u2_u6_n132 ) , .A3( u2_u2_u6_n145 ) );
  INV_X1 u2_u2_u6_U28 (.A( u2_u2_u6_n146 ) , .ZN( u2_u2_u6_n163 ) );
  AOI222_X1 u2_u2_u6_U29 (.ZN( u2_u2_u6_n114 ) , .A1( u2_u2_u6_n118 ) , .A2( u2_u2_u6_n126 ) , .B2( u2_u2_u6_n151 ) , .C2( u2_u2_u6_n159 ) , .C1( u2_u2_u6_n168 ) , .B1( u2_u2_u6_n169 ) );
  INV_X1 u2_u2_u6_U3 (.A( u2_u2_u6_n110 ) , .ZN( u2_u2_u6_n166 ) );
  NOR2_X1 u2_u2_u6_U30 (.A1( u2_u2_u6_n162 ) , .A2( u2_u2_u6_n165 ) , .ZN( u2_u2_u6_n98 ) );
  NAND2_X1 u2_u2_u6_U31 (.A1( u2_u2_u6_n144 ) , .ZN( u2_u2_u6_n151 ) , .A2( u2_u2_u6_n158 ) );
  NAND2_X1 u2_u2_u6_U32 (.ZN( u2_u2_u6_n132 ) , .A1( u2_u2_u6_n91 ) , .A2( u2_u2_u6_n97 ) );
  AOI22_X1 u2_u2_u6_U33 (.B2( u2_u2_u6_n110 ) , .B1( u2_u2_u6_n111 ) , .A1( u2_u2_u6_n112 ) , .ZN( u2_u2_u6_n115 ) , .A2( u2_u2_u6_n161 ) );
  NAND4_X1 u2_u2_u6_U34 (.A3( u2_u2_u6_n109 ) , .ZN( u2_u2_u6_n112 ) , .A4( u2_u2_u6_n132 ) , .A2( u2_u2_u6_n147 ) , .A1( u2_u2_u6_n166 ) );
  NOR2_X1 u2_u2_u6_U35 (.ZN( u2_u2_u6_n109 ) , .A1( u2_u2_u6_n170 ) , .A2( u2_u2_u6_n173 ) );
  NOR2_X1 u2_u2_u6_U36 (.A2( u2_u2_u6_n126 ) , .ZN( u2_u2_u6_n155 ) , .A1( u2_u2_u6_n160 ) );
  NAND2_X1 u2_u2_u6_U37 (.ZN( u2_u2_u6_n146 ) , .A2( u2_u2_u6_n94 ) , .A1( u2_u2_u6_n99 ) );
  AOI21_X1 u2_u2_u6_U38 (.A( u2_u2_u6_n144 ) , .B2( u2_u2_u6_n145 ) , .B1( u2_u2_u6_n146 ) , .ZN( u2_u2_u6_n150 ) );
  INV_X1 u2_u2_u6_U39 (.A( u2_u2_u6_n111 ) , .ZN( u2_u2_u6_n158 ) );
  INV_X1 u2_u2_u6_U4 (.A( u2_u2_u6_n142 ) , .ZN( u2_u2_u6_n174 ) );
  NAND2_X1 u2_u2_u6_U40 (.ZN( u2_u2_u6_n127 ) , .A1( u2_u2_u6_n91 ) , .A2( u2_u2_u6_n92 ) );
  NAND2_X1 u2_u2_u6_U41 (.ZN( u2_u2_u6_n129 ) , .A2( u2_u2_u6_n95 ) , .A1( u2_u2_u6_n96 ) );
  INV_X1 u2_u2_u6_U42 (.A( u2_u2_u6_n144 ) , .ZN( u2_u2_u6_n159 ) );
  NAND2_X1 u2_u2_u6_U43 (.ZN( u2_u2_u6_n145 ) , .A2( u2_u2_u6_n97 ) , .A1( u2_u2_u6_n98 ) );
  NAND2_X1 u2_u2_u6_U44 (.ZN( u2_u2_u6_n148 ) , .A2( u2_u2_u6_n92 ) , .A1( u2_u2_u6_n94 ) );
  NAND2_X1 u2_u2_u6_U45 (.ZN( u2_u2_u6_n108 ) , .A2( u2_u2_u6_n139 ) , .A1( u2_u2_u6_n144 ) );
  NAND2_X1 u2_u2_u6_U46 (.ZN( u2_u2_u6_n121 ) , .A2( u2_u2_u6_n95 ) , .A1( u2_u2_u6_n97 ) );
  NAND2_X1 u2_u2_u6_U47 (.ZN( u2_u2_u6_n107 ) , .A2( u2_u2_u6_n92 ) , .A1( u2_u2_u6_n95 ) );
  AND2_X1 u2_u2_u6_U48 (.ZN( u2_u2_u6_n118 ) , .A2( u2_u2_u6_n91 ) , .A1( u2_u2_u6_n99 ) );
  NAND2_X1 u2_u2_u6_U49 (.ZN( u2_u2_u6_n147 ) , .A2( u2_u2_u6_n98 ) , .A1( u2_u2_u6_n99 ) );
  NAND2_X1 u2_u2_u6_U5 (.A2( u2_u2_u6_n143 ) , .ZN( u2_u2_u6_n152 ) , .A1( u2_u2_u6_n166 ) );
  NAND2_X1 u2_u2_u6_U50 (.ZN( u2_u2_u6_n128 ) , .A1( u2_u2_u6_n94 ) , .A2( u2_u2_u6_n96 ) );
  AOI211_X1 u2_u2_u6_U51 (.B( u2_u2_u6_n134 ) , .A( u2_u2_u6_n135 ) , .C1( u2_u2_u6_n136 ) , .ZN( u2_u2_u6_n137 ) , .C2( u2_u2_u6_n151 ) );
  AOI21_X1 u2_u2_u6_U52 (.B2( u2_u2_u6_n132 ) , .B1( u2_u2_u6_n133 ) , .ZN( u2_u2_u6_n134 ) , .A( u2_u2_u6_n158 ) );
  AOI21_X1 u2_u2_u6_U53 (.B1( u2_u2_u6_n131 ) , .ZN( u2_u2_u6_n135 ) , .A( u2_u2_u6_n144 ) , .B2( u2_u2_u6_n146 ) );
  NAND4_X1 u2_u2_u6_U54 (.A4( u2_u2_u6_n127 ) , .A3( u2_u2_u6_n128 ) , .A2( u2_u2_u6_n129 ) , .A1( u2_u2_u6_n130 ) , .ZN( u2_u2_u6_n136 ) );
  NAND2_X1 u2_u2_u6_U55 (.ZN( u2_u2_u6_n119 ) , .A2( u2_u2_u6_n95 ) , .A1( u2_u2_u6_n99 ) );
  NAND2_X1 u2_u2_u6_U56 (.ZN( u2_u2_u6_n123 ) , .A2( u2_u2_u6_n91 ) , .A1( u2_u2_u6_n96 ) );
  NAND2_X1 u2_u2_u6_U57 (.ZN( u2_u2_u6_n100 ) , .A2( u2_u2_u6_n92 ) , .A1( u2_u2_u6_n98 ) );
  NAND2_X1 u2_u2_u6_U58 (.ZN( u2_u2_u6_n122 ) , .A1( u2_u2_u6_n94 ) , .A2( u2_u2_u6_n97 ) );
  INV_X1 u2_u2_u6_U59 (.A( u2_u2_u6_n139 ) , .ZN( u2_u2_u6_n160 ) );
  AOI22_X1 u2_u2_u6_U6 (.B2( u2_u2_u6_n101 ) , .A1( u2_u2_u6_n102 ) , .ZN( u2_u2_u6_n103 ) , .B1( u2_u2_u6_n160 ) , .A2( u2_u2_u6_n161 ) );
  NAND2_X1 u2_u2_u6_U60 (.ZN( u2_u2_u6_n113 ) , .A1( u2_u2_u6_n96 ) , .A2( u2_u2_u6_n98 ) );
  NOR2_X1 u2_u2_u6_U61 (.A2( u2_u2_X_40 ) , .A1( u2_u2_X_41 ) , .ZN( u2_u2_u6_n126 ) );
  NOR2_X1 u2_u2_u6_U62 (.A2( u2_u2_X_39 ) , .A1( u2_u2_X_42 ) , .ZN( u2_u2_u6_n92 ) );
  NOR2_X1 u2_u2_u6_U63 (.A2( u2_u2_X_39 ) , .A1( u2_u2_u6_n156 ) , .ZN( u2_u2_u6_n97 ) );
  NOR2_X1 u2_u2_u6_U64 (.A2( u2_u2_X_38 ) , .A1( u2_u2_u6_n165 ) , .ZN( u2_u2_u6_n95 ) );
  NOR2_X1 u2_u2_u6_U65 (.A2( u2_u2_X_41 ) , .ZN( u2_u2_u6_n111 ) , .A1( u2_u2_u6_n157 ) );
  NOR2_X1 u2_u2_u6_U66 (.A2( u2_u2_X_37 ) , .A1( u2_u2_u6_n162 ) , .ZN( u2_u2_u6_n94 ) );
  NOR2_X1 u2_u2_u6_U67 (.A2( u2_u2_X_37 ) , .A1( u2_u2_X_38 ) , .ZN( u2_u2_u6_n91 ) );
  NAND2_X1 u2_u2_u6_U68 (.A1( u2_u2_X_41 ) , .ZN( u2_u2_u6_n144 ) , .A2( u2_u2_u6_n157 ) );
  NAND2_X1 u2_u2_u6_U69 (.A2( u2_u2_X_40 ) , .A1( u2_u2_X_41 ) , .ZN( u2_u2_u6_n139 ) );
  NOR2_X1 u2_u2_u6_U7 (.A1( u2_u2_u6_n118 ) , .ZN( u2_u2_u6_n143 ) , .A2( u2_u2_u6_n168 ) );
  AND2_X1 u2_u2_u6_U70 (.A1( u2_u2_X_39 ) , .A2( u2_u2_u6_n156 ) , .ZN( u2_u2_u6_n96 ) );
  AND2_X1 u2_u2_u6_U71 (.A1( u2_u2_X_39 ) , .A2( u2_u2_X_42 ) , .ZN( u2_u2_u6_n99 ) );
  INV_X1 u2_u2_u6_U72 (.A( u2_u2_X_40 ) , .ZN( u2_u2_u6_n157 ) );
  INV_X1 u2_u2_u6_U73 (.A( u2_u2_X_37 ) , .ZN( u2_u2_u6_n165 ) );
  INV_X1 u2_u2_u6_U74 (.A( u2_u2_X_38 ) , .ZN( u2_u2_u6_n162 ) );
  INV_X1 u2_u2_u6_U75 (.A( u2_u2_X_42 ) , .ZN( u2_u2_u6_n156 ) );
  NAND4_X1 u2_u2_u6_U76 (.ZN( u2_out2_32 ) , .A4( u2_u2_u6_n103 ) , .A3( u2_u2_u6_n104 ) , .A2( u2_u2_u6_n105 ) , .A1( u2_u2_u6_n106 ) );
  AOI22_X1 u2_u2_u6_U77 (.ZN( u2_u2_u6_n105 ) , .A2( u2_u2_u6_n108 ) , .A1( u2_u2_u6_n118 ) , .B2( u2_u2_u6_n126 ) , .B1( u2_u2_u6_n171 ) );
  AOI22_X1 u2_u2_u6_U78 (.ZN( u2_u2_u6_n104 ) , .A1( u2_u2_u6_n111 ) , .B1( u2_u2_u6_n124 ) , .B2( u2_u2_u6_n151 ) , .A2( u2_u2_u6_n93 ) );
  NAND4_X1 u2_u2_u6_U79 (.ZN( u2_out2_12 ) , .A4( u2_u2_u6_n114 ) , .A3( u2_u2_u6_n115 ) , .A2( u2_u2_u6_n116 ) , .A1( u2_u2_u6_n117 ) );
  AOI21_X1 u2_u2_u6_U8 (.B1( u2_u2_u6_n107 ) , .B2( u2_u2_u6_n132 ) , .A( u2_u2_u6_n158 ) , .ZN( u2_u2_u6_n88 ) );
  OAI22_X1 u2_u2_u6_U80 (.B2( u2_u2_u6_n111 ) , .ZN( u2_u2_u6_n116 ) , .B1( u2_u2_u6_n126 ) , .A2( u2_u2_u6_n164 ) , .A1( u2_u2_u6_n167 ) );
  OAI21_X1 u2_u2_u6_U81 (.A( u2_u2_u6_n108 ) , .ZN( u2_u2_u6_n117 ) , .B2( u2_u2_u6_n141 ) , .B1( u2_u2_u6_n163 ) );
  OAI211_X1 u2_u2_u6_U82 (.ZN( u2_out2_7 ) , .B( u2_u2_u6_n153 ) , .C2( u2_u2_u6_n154 ) , .C1( u2_u2_u6_n155 ) , .A( u2_u2_u6_n174 ) );
  NOR3_X1 u2_u2_u6_U83 (.A1( u2_u2_u6_n141 ) , .ZN( u2_u2_u6_n154 ) , .A3( u2_u2_u6_n164 ) , .A2( u2_u2_u6_n171 ) );
  AOI211_X1 u2_u2_u6_U84 (.B( u2_u2_u6_n149 ) , .A( u2_u2_u6_n150 ) , .C2( u2_u2_u6_n151 ) , .C1( u2_u2_u6_n152 ) , .ZN( u2_u2_u6_n153 ) );
  OAI211_X1 u2_u2_u6_U85 (.ZN( u2_out2_22 ) , .B( u2_u2_u6_n137 ) , .A( u2_u2_u6_n138 ) , .C2( u2_u2_u6_n139 ) , .C1( u2_u2_u6_n140 ) );
  AOI22_X1 u2_u2_u6_U86 (.B1( u2_u2_u6_n124 ) , .A2( u2_u2_u6_n125 ) , .A1( u2_u2_u6_n126 ) , .ZN( u2_u2_u6_n138 ) , .B2( u2_u2_u6_n161 ) );
  AND4_X1 u2_u2_u6_U87 (.A3( u2_u2_u6_n119 ) , .A1( u2_u2_u6_n120 ) , .A4( u2_u2_u6_n129 ) , .ZN( u2_u2_u6_n140 ) , .A2( u2_u2_u6_n143 ) );
  NAND3_X1 u2_u2_u6_U88 (.A2( u2_u2_u6_n123 ) , .ZN( u2_u2_u6_n125 ) , .A1( u2_u2_u6_n130 ) , .A3( u2_u2_u6_n131 ) );
  NAND3_X1 u2_u2_u6_U89 (.A3( u2_u2_u6_n133 ) , .ZN( u2_u2_u6_n141 ) , .A1( u2_u2_u6_n145 ) , .A2( u2_u2_u6_n148 ) );
  AOI21_X1 u2_u2_u6_U9 (.B2( u2_u2_u6_n147 ) , .B1( u2_u2_u6_n148 ) , .ZN( u2_u2_u6_n149 ) , .A( u2_u2_u6_n158 ) );
  NAND3_X1 u2_u2_u6_U90 (.ZN( u2_u2_u6_n101 ) , .A3( u2_u2_u6_n107 ) , .A2( u2_u2_u6_n121 ) , .A1( u2_u2_u6_n127 ) );
  NAND3_X1 u2_u2_u6_U91 (.ZN( u2_u2_u6_n102 ) , .A3( u2_u2_u6_n130 ) , .A2( u2_u2_u6_n145 ) , .A1( u2_u2_u6_n166 ) );
  NAND3_X1 u2_u2_u6_U92 (.A3( u2_u2_u6_n113 ) , .A1( u2_u2_u6_n119 ) , .A2( u2_u2_u6_n123 ) , .ZN( u2_u2_u6_n93 ) );
  NAND3_X1 u2_u2_u6_U93 (.ZN( u2_u2_u6_n142 ) , .A2( u2_u2_u6_n172 ) , .A3( u2_u2_u6_n89 ) , .A1( u2_u2_u6_n90 ) );
  AND3_X1 u2_u2_u7_U10 (.A3( u2_u2_u7_n110 ) , .A2( u2_u2_u7_n127 ) , .A1( u2_u2_u7_n132 ) , .ZN( u2_u2_u7_n92 ) );
  OAI21_X1 u2_u2_u7_U11 (.A( u2_u2_u7_n161 ) , .B1( u2_u2_u7_n168 ) , .B2( u2_u2_u7_n173 ) , .ZN( u2_u2_u7_n91 ) );
  AOI211_X1 u2_u2_u7_U12 (.A( u2_u2_u7_n117 ) , .ZN( u2_u2_u7_n118 ) , .C2( u2_u2_u7_n126 ) , .C1( u2_u2_u7_n177 ) , .B( u2_u2_u7_n180 ) );
  OAI22_X1 u2_u2_u7_U13 (.B1( u2_u2_u7_n115 ) , .ZN( u2_u2_u7_n117 ) , .A2( u2_u2_u7_n133 ) , .A1( u2_u2_u7_n137 ) , .B2( u2_u2_u7_n162 ) );
  INV_X1 u2_u2_u7_U14 (.A( u2_u2_u7_n116 ) , .ZN( u2_u2_u7_n180 ) );
  NOR3_X1 u2_u2_u7_U15 (.ZN( u2_u2_u7_n115 ) , .A3( u2_u2_u7_n145 ) , .A2( u2_u2_u7_n168 ) , .A1( u2_u2_u7_n169 ) );
  OAI211_X1 u2_u2_u7_U16 (.B( u2_u2_u7_n122 ) , .A( u2_u2_u7_n123 ) , .C2( u2_u2_u7_n124 ) , .ZN( u2_u2_u7_n154 ) , .C1( u2_u2_u7_n162 ) );
  AOI222_X1 u2_u2_u7_U17 (.ZN( u2_u2_u7_n122 ) , .C2( u2_u2_u7_n126 ) , .C1( u2_u2_u7_n145 ) , .B1( u2_u2_u7_n161 ) , .A2( u2_u2_u7_n165 ) , .B2( u2_u2_u7_n170 ) , .A1( u2_u2_u7_n176 ) );
  INV_X1 u2_u2_u7_U18 (.A( u2_u2_u7_n133 ) , .ZN( u2_u2_u7_n176 ) );
  NOR3_X1 u2_u2_u7_U19 (.A2( u2_u2_u7_n134 ) , .A1( u2_u2_u7_n135 ) , .ZN( u2_u2_u7_n136 ) , .A3( u2_u2_u7_n171 ) );
  NOR2_X1 u2_u2_u7_U20 (.A1( u2_u2_u7_n130 ) , .A2( u2_u2_u7_n134 ) , .ZN( u2_u2_u7_n153 ) );
  INV_X1 u2_u2_u7_U21 (.A( u2_u2_u7_n101 ) , .ZN( u2_u2_u7_n165 ) );
  NOR2_X1 u2_u2_u7_U22 (.ZN( u2_u2_u7_n111 ) , .A2( u2_u2_u7_n134 ) , .A1( u2_u2_u7_n169 ) );
  AOI21_X1 u2_u2_u7_U23 (.ZN( u2_u2_u7_n104 ) , .B2( u2_u2_u7_n112 ) , .B1( u2_u2_u7_n127 ) , .A( u2_u2_u7_n164 ) );
  AOI21_X1 u2_u2_u7_U24 (.ZN( u2_u2_u7_n106 ) , .B1( u2_u2_u7_n133 ) , .B2( u2_u2_u7_n146 ) , .A( u2_u2_u7_n162 ) );
  AOI21_X1 u2_u2_u7_U25 (.A( u2_u2_u7_n101 ) , .ZN( u2_u2_u7_n107 ) , .B2( u2_u2_u7_n128 ) , .B1( u2_u2_u7_n175 ) );
  INV_X1 u2_u2_u7_U26 (.A( u2_u2_u7_n138 ) , .ZN( u2_u2_u7_n171 ) );
  INV_X1 u2_u2_u7_U27 (.A( u2_u2_u7_n131 ) , .ZN( u2_u2_u7_n177 ) );
  INV_X1 u2_u2_u7_U28 (.A( u2_u2_u7_n110 ) , .ZN( u2_u2_u7_n174 ) );
  NAND2_X1 u2_u2_u7_U29 (.A1( u2_u2_u7_n129 ) , .A2( u2_u2_u7_n132 ) , .ZN( u2_u2_u7_n149 ) );
  OAI21_X1 u2_u2_u7_U3 (.ZN( u2_u2_u7_n159 ) , .A( u2_u2_u7_n165 ) , .B2( u2_u2_u7_n171 ) , .B1( u2_u2_u7_n174 ) );
  NAND2_X1 u2_u2_u7_U30 (.A1( u2_u2_u7_n113 ) , .A2( u2_u2_u7_n124 ) , .ZN( u2_u2_u7_n130 ) );
  INV_X1 u2_u2_u7_U31 (.A( u2_u2_u7_n112 ) , .ZN( u2_u2_u7_n173 ) );
  INV_X1 u2_u2_u7_U32 (.A( u2_u2_u7_n128 ) , .ZN( u2_u2_u7_n168 ) );
  INV_X1 u2_u2_u7_U33 (.A( u2_u2_u7_n148 ) , .ZN( u2_u2_u7_n169 ) );
  INV_X1 u2_u2_u7_U34 (.A( u2_u2_u7_n127 ) , .ZN( u2_u2_u7_n179 ) );
  NOR2_X1 u2_u2_u7_U35 (.ZN( u2_u2_u7_n101 ) , .A2( u2_u2_u7_n150 ) , .A1( u2_u2_u7_n156 ) );
  AOI211_X1 u2_u2_u7_U36 (.B( u2_u2_u7_n154 ) , .A( u2_u2_u7_n155 ) , .C1( u2_u2_u7_n156 ) , .ZN( u2_u2_u7_n157 ) , .C2( u2_u2_u7_n172 ) );
  INV_X1 u2_u2_u7_U37 (.A( u2_u2_u7_n153 ) , .ZN( u2_u2_u7_n172 ) );
  AOI211_X1 u2_u2_u7_U38 (.B( u2_u2_u7_n139 ) , .A( u2_u2_u7_n140 ) , .C2( u2_u2_u7_n141 ) , .ZN( u2_u2_u7_n142 ) , .C1( u2_u2_u7_n156 ) );
  NAND4_X1 u2_u2_u7_U39 (.A3( u2_u2_u7_n127 ) , .A2( u2_u2_u7_n128 ) , .A1( u2_u2_u7_n129 ) , .ZN( u2_u2_u7_n141 ) , .A4( u2_u2_u7_n147 ) );
  INV_X1 u2_u2_u7_U4 (.A( u2_u2_u7_n111 ) , .ZN( u2_u2_u7_n170 ) );
  AOI21_X1 u2_u2_u7_U40 (.A( u2_u2_u7_n137 ) , .B1( u2_u2_u7_n138 ) , .ZN( u2_u2_u7_n139 ) , .B2( u2_u2_u7_n146 ) );
  OAI22_X1 u2_u2_u7_U41 (.B1( u2_u2_u7_n136 ) , .ZN( u2_u2_u7_n140 ) , .A1( u2_u2_u7_n153 ) , .B2( u2_u2_u7_n162 ) , .A2( u2_u2_u7_n164 ) );
  AOI21_X1 u2_u2_u7_U42 (.ZN( u2_u2_u7_n123 ) , .B1( u2_u2_u7_n165 ) , .B2( u2_u2_u7_n177 ) , .A( u2_u2_u7_n97 ) );
  AOI21_X1 u2_u2_u7_U43 (.B2( u2_u2_u7_n113 ) , .B1( u2_u2_u7_n124 ) , .A( u2_u2_u7_n125 ) , .ZN( u2_u2_u7_n97 ) );
  INV_X1 u2_u2_u7_U44 (.A( u2_u2_u7_n125 ) , .ZN( u2_u2_u7_n161 ) );
  INV_X1 u2_u2_u7_U45 (.A( u2_u2_u7_n152 ) , .ZN( u2_u2_u7_n162 ) );
  AOI22_X1 u2_u2_u7_U46 (.A2( u2_u2_u7_n114 ) , .ZN( u2_u2_u7_n119 ) , .B1( u2_u2_u7_n130 ) , .A1( u2_u2_u7_n156 ) , .B2( u2_u2_u7_n165 ) );
  NAND2_X1 u2_u2_u7_U47 (.A2( u2_u2_u7_n112 ) , .ZN( u2_u2_u7_n114 ) , .A1( u2_u2_u7_n175 ) );
  AND2_X1 u2_u2_u7_U48 (.ZN( u2_u2_u7_n145 ) , .A2( u2_u2_u7_n98 ) , .A1( u2_u2_u7_n99 ) );
  NOR2_X1 u2_u2_u7_U49 (.ZN( u2_u2_u7_n137 ) , .A1( u2_u2_u7_n150 ) , .A2( u2_u2_u7_n161 ) );
  INV_X1 u2_u2_u7_U5 (.A( u2_u2_u7_n149 ) , .ZN( u2_u2_u7_n175 ) );
  AOI21_X1 u2_u2_u7_U50 (.ZN( u2_u2_u7_n105 ) , .B2( u2_u2_u7_n110 ) , .A( u2_u2_u7_n125 ) , .B1( u2_u2_u7_n147 ) );
  NAND2_X1 u2_u2_u7_U51 (.ZN( u2_u2_u7_n146 ) , .A1( u2_u2_u7_n95 ) , .A2( u2_u2_u7_n98 ) );
  NAND2_X1 u2_u2_u7_U52 (.A2( u2_u2_u7_n103 ) , .ZN( u2_u2_u7_n147 ) , .A1( u2_u2_u7_n93 ) );
  NAND2_X1 u2_u2_u7_U53 (.A1( u2_u2_u7_n103 ) , .ZN( u2_u2_u7_n127 ) , .A2( u2_u2_u7_n99 ) );
  OR2_X1 u2_u2_u7_U54 (.ZN( u2_u2_u7_n126 ) , .A2( u2_u2_u7_n152 ) , .A1( u2_u2_u7_n156 ) );
  NAND2_X1 u2_u2_u7_U55 (.A2( u2_u2_u7_n102 ) , .A1( u2_u2_u7_n103 ) , .ZN( u2_u2_u7_n133 ) );
  NAND2_X1 u2_u2_u7_U56 (.ZN( u2_u2_u7_n112 ) , .A2( u2_u2_u7_n96 ) , .A1( u2_u2_u7_n99 ) );
  NAND2_X1 u2_u2_u7_U57 (.A2( u2_u2_u7_n102 ) , .ZN( u2_u2_u7_n128 ) , .A1( u2_u2_u7_n98 ) );
  NAND2_X1 u2_u2_u7_U58 (.A1( u2_u2_u7_n100 ) , .ZN( u2_u2_u7_n113 ) , .A2( u2_u2_u7_n93 ) );
  NAND2_X1 u2_u2_u7_U59 (.A2( u2_u2_u7_n102 ) , .ZN( u2_u2_u7_n124 ) , .A1( u2_u2_u7_n96 ) );
  INV_X1 u2_u2_u7_U6 (.A( u2_u2_u7_n154 ) , .ZN( u2_u2_u7_n178 ) );
  NAND2_X1 u2_u2_u7_U60 (.ZN( u2_u2_u7_n110 ) , .A1( u2_u2_u7_n95 ) , .A2( u2_u2_u7_n96 ) );
  INV_X1 u2_u2_u7_U61 (.A( u2_u2_u7_n150 ) , .ZN( u2_u2_u7_n164 ) );
  AND2_X1 u2_u2_u7_U62 (.ZN( u2_u2_u7_n134 ) , .A1( u2_u2_u7_n93 ) , .A2( u2_u2_u7_n98 ) );
  NAND2_X1 u2_u2_u7_U63 (.A1( u2_u2_u7_n100 ) , .A2( u2_u2_u7_n102 ) , .ZN( u2_u2_u7_n129 ) );
  NAND2_X1 u2_u2_u7_U64 (.A2( u2_u2_u7_n103 ) , .ZN( u2_u2_u7_n131 ) , .A1( u2_u2_u7_n95 ) );
  NAND2_X1 u2_u2_u7_U65 (.A1( u2_u2_u7_n100 ) , .ZN( u2_u2_u7_n138 ) , .A2( u2_u2_u7_n99 ) );
  NAND2_X1 u2_u2_u7_U66 (.ZN( u2_u2_u7_n132 ) , .A1( u2_u2_u7_n93 ) , .A2( u2_u2_u7_n96 ) );
  NAND2_X1 u2_u2_u7_U67 (.A1( u2_u2_u7_n100 ) , .ZN( u2_u2_u7_n148 ) , .A2( u2_u2_u7_n95 ) );
  NOR2_X1 u2_u2_u7_U68 (.A2( u2_u2_X_47 ) , .ZN( u2_u2_u7_n150 ) , .A1( u2_u2_u7_n163 ) );
  NOR2_X1 u2_u2_u7_U69 (.A2( u2_u2_X_43 ) , .A1( u2_u2_X_44 ) , .ZN( u2_u2_u7_n103 ) );
  AOI211_X1 u2_u2_u7_U7 (.ZN( u2_u2_u7_n116 ) , .A( u2_u2_u7_n155 ) , .C1( u2_u2_u7_n161 ) , .C2( u2_u2_u7_n171 ) , .B( u2_u2_u7_n94 ) );
  NOR2_X1 u2_u2_u7_U70 (.A2( u2_u2_X_48 ) , .A1( u2_u2_u7_n166 ) , .ZN( u2_u2_u7_n95 ) );
  NOR2_X1 u2_u2_u7_U71 (.A2( u2_u2_X_45 ) , .A1( u2_u2_X_48 ) , .ZN( u2_u2_u7_n99 ) );
  NOR2_X1 u2_u2_u7_U72 (.A2( u2_u2_X_44 ) , .A1( u2_u2_u7_n167 ) , .ZN( u2_u2_u7_n98 ) );
  NOR2_X1 u2_u2_u7_U73 (.A2( u2_u2_X_46 ) , .A1( u2_u2_X_47 ) , .ZN( u2_u2_u7_n152 ) );
  AND2_X1 u2_u2_u7_U74 (.A1( u2_u2_X_47 ) , .ZN( u2_u2_u7_n156 ) , .A2( u2_u2_u7_n163 ) );
  NAND2_X1 u2_u2_u7_U75 (.A2( u2_u2_X_46 ) , .A1( u2_u2_X_47 ) , .ZN( u2_u2_u7_n125 ) );
  AND2_X1 u2_u2_u7_U76 (.A2( u2_u2_X_45 ) , .A1( u2_u2_X_48 ) , .ZN( u2_u2_u7_n102 ) );
  AND2_X1 u2_u2_u7_U77 (.A2( u2_u2_X_43 ) , .A1( u2_u2_X_44 ) , .ZN( u2_u2_u7_n96 ) );
  AND2_X1 u2_u2_u7_U78 (.A1( u2_u2_X_44 ) , .ZN( u2_u2_u7_n100 ) , .A2( u2_u2_u7_n167 ) );
  AND2_X1 u2_u2_u7_U79 (.A1( u2_u2_X_48 ) , .A2( u2_u2_u7_n166 ) , .ZN( u2_u2_u7_n93 ) );
  OAI222_X1 u2_u2_u7_U8 (.C2( u2_u2_u7_n101 ) , .B2( u2_u2_u7_n111 ) , .A1( u2_u2_u7_n113 ) , .C1( u2_u2_u7_n146 ) , .A2( u2_u2_u7_n162 ) , .B1( u2_u2_u7_n164 ) , .ZN( u2_u2_u7_n94 ) );
  INV_X1 u2_u2_u7_U80 (.A( u2_u2_X_46 ) , .ZN( u2_u2_u7_n163 ) );
  INV_X1 u2_u2_u7_U81 (.A( u2_u2_X_43 ) , .ZN( u2_u2_u7_n167 ) );
  INV_X1 u2_u2_u7_U82 (.A( u2_u2_X_45 ) , .ZN( u2_u2_u7_n166 ) );
  NAND4_X1 u2_u2_u7_U83 (.ZN( u2_out2_5 ) , .A4( u2_u2_u7_n108 ) , .A3( u2_u2_u7_n109 ) , .A1( u2_u2_u7_n116 ) , .A2( u2_u2_u7_n123 ) );
  AOI22_X1 u2_u2_u7_U84 (.ZN( u2_u2_u7_n109 ) , .A2( u2_u2_u7_n126 ) , .B2( u2_u2_u7_n145 ) , .B1( u2_u2_u7_n156 ) , .A1( u2_u2_u7_n171 ) );
  NOR4_X1 u2_u2_u7_U85 (.A4( u2_u2_u7_n104 ) , .A3( u2_u2_u7_n105 ) , .A2( u2_u2_u7_n106 ) , .A1( u2_u2_u7_n107 ) , .ZN( u2_u2_u7_n108 ) );
  NAND4_X1 u2_u2_u7_U86 (.ZN( u2_out2_27 ) , .A4( u2_u2_u7_n118 ) , .A3( u2_u2_u7_n119 ) , .A2( u2_u2_u7_n120 ) , .A1( u2_u2_u7_n121 ) );
  OAI21_X1 u2_u2_u7_U87 (.ZN( u2_u2_u7_n121 ) , .B2( u2_u2_u7_n145 ) , .A( u2_u2_u7_n150 ) , .B1( u2_u2_u7_n174 ) );
  OAI21_X1 u2_u2_u7_U88 (.ZN( u2_u2_u7_n120 ) , .A( u2_u2_u7_n161 ) , .B2( u2_u2_u7_n170 ) , .B1( u2_u2_u7_n179 ) );
  NAND4_X1 u2_u2_u7_U89 (.ZN( u2_out2_21 ) , .A4( u2_u2_u7_n157 ) , .A3( u2_u2_u7_n158 ) , .A2( u2_u2_u7_n159 ) , .A1( u2_u2_u7_n160 ) );
  OAI221_X1 u2_u2_u7_U9 (.C1( u2_u2_u7_n101 ) , .C2( u2_u2_u7_n147 ) , .ZN( u2_u2_u7_n155 ) , .B2( u2_u2_u7_n162 ) , .A( u2_u2_u7_n91 ) , .B1( u2_u2_u7_n92 ) );
  OAI21_X1 u2_u2_u7_U90 (.B1( u2_u2_u7_n145 ) , .ZN( u2_u2_u7_n160 ) , .A( u2_u2_u7_n161 ) , .B2( u2_u2_u7_n177 ) );
  AOI22_X1 u2_u2_u7_U91 (.B2( u2_u2_u7_n149 ) , .B1( u2_u2_u7_n150 ) , .A2( u2_u2_u7_n151 ) , .A1( u2_u2_u7_n152 ) , .ZN( u2_u2_u7_n158 ) );
  NAND4_X1 u2_u2_u7_U92 (.ZN( u2_out2_15 ) , .A4( u2_u2_u7_n142 ) , .A3( u2_u2_u7_n143 ) , .A2( u2_u2_u7_n144 ) , .A1( u2_u2_u7_n178 ) );
  OR2_X1 u2_u2_u7_U93 (.A2( u2_u2_u7_n125 ) , .A1( u2_u2_u7_n129 ) , .ZN( u2_u2_u7_n144 ) );
  AOI22_X1 u2_u2_u7_U94 (.A2( u2_u2_u7_n126 ) , .ZN( u2_u2_u7_n143 ) , .B2( u2_u2_u7_n165 ) , .B1( u2_u2_u7_n173 ) , .A1( u2_u2_u7_n174 ) );
  NAND3_X1 u2_u2_u7_U95 (.A3( u2_u2_u7_n146 ) , .A2( u2_u2_u7_n147 ) , .A1( u2_u2_u7_n148 ) , .ZN( u2_u2_u7_n151 ) );
  NAND3_X1 u2_u2_u7_U96 (.A3( u2_u2_u7_n131 ) , .A2( u2_u2_u7_n132 ) , .A1( u2_u2_u7_n133 ) , .ZN( u2_u2_u7_n135 ) );
  XOR2_X1 u2_u3_U13 (.B( u2_K4_42 ) , .A( u2_R2_29 ) , .Z( u2_u3_X_42 ) );
  XOR2_X1 u2_u3_U14 (.B( u2_K4_41 ) , .A( u2_R2_28 ) , .Z( u2_u3_X_41 ) );
  XOR2_X1 u2_u3_U15 (.B( u2_K4_40 ) , .A( u2_R2_27 ) , .Z( u2_u3_X_40 ) );
  XOR2_X1 u2_u3_U17 (.B( u2_K4_39 ) , .A( u2_R2_26 ) , .Z( u2_u3_X_39 ) );
  XOR2_X1 u2_u3_U18 (.B( u2_K4_38 ) , .A( u2_R2_25 ) , .Z( u2_u3_X_38 ) );
  XOR2_X1 u2_u3_U19 (.B( u2_K4_37 ) , .A( u2_R2_24 ) , .Z( u2_u3_X_37 ) );
  XOR2_X1 u2_u3_U20 (.B( u2_K4_36 ) , .A( u2_R2_25 ) , .Z( u2_u3_X_36 ) );
  XOR2_X1 u2_u3_U21 (.B( u2_K4_35 ) , .A( u2_R2_24 ) , .Z( u2_u3_X_35 ) );
  XOR2_X1 u2_u3_U22 (.B( u2_K4_34 ) , .A( u2_R2_23 ) , .Z( u2_u3_X_34 ) );
  XOR2_X1 u2_u3_U23 (.B( u2_K4_33 ) , .A( u2_R2_22 ) , .Z( u2_u3_X_33 ) );
  XOR2_X1 u2_u3_U24 (.B( u2_K4_32 ) , .A( u2_R2_21 ) , .Z( u2_u3_X_32 ) );
  XOR2_X1 u2_u3_U25 (.B( u2_K4_31 ) , .A( u2_R2_20 ) , .Z( u2_u3_X_31 ) );
  XOR2_X1 u2_u3_U26 (.B( u2_K4_30 ) , .A( u2_R2_21 ) , .Z( u2_u3_X_30 ) );
  XOR2_X1 u2_u3_U28 (.B( u2_K4_29 ) , .A( u2_R2_20 ) , .Z( u2_u3_X_29 ) );
  XOR2_X1 u2_u3_U29 (.B( u2_K4_28 ) , .A( u2_R2_19 ) , .Z( u2_u3_X_28 ) );
  XOR2_X1 u2_u3_U30 (.B( u2_K4_27 ) , .A( u2_R2_18 ) , .Z( u2_u3_X_27 ) );
  XOR2_X1 u2_u3_U31 (.B( u2_K4_26 ) , .A( u2_R2_17 ) , .Z( u2_u3_X_26 ) );
  XOR2_X1 u2_u3_U32 (.B( u2_K4_25 ) , .A( u2_R2_16 ) , .Z( u2_u3_X_25 ) );
  OAI22_X1 u2_u3_u4_U10 (.B2( u2_u3_u4_n135 ) , .ZN( u2_u3_u4_n137 ) , .B1( u2_u3_u4_n153 ) , .A1( u2_u3_u4_n155 ) , .A2( u2_u3_u4_n171 ) );
  AND3_X1 u2_u3_u4_U11 (.A2( u2_u3_u4_n134 ) , .ZN( u2_u3_u4_n135 ) , .A3( u2_u3_u4_n145 ) , .A1( u2_u3_u4_n157 ) );
  OR3_X1 u2_u3_u4_U12 (.A3( u2_u3_u4_n114 ) , .A2( u2_u3_u4_n115 ) , .A1( u2_u3_u4_n116 ) , .ZN( u2_u3_u4_n136 ) );
  AOI21_X1 u2_u3_u4_U13 (.A( u2_u3_u4_n113 ) , .ZN( u2_u3_u4_n116 ) , .B2( u2_u3_u4_n173 ) , .B1( u2_u3_u4_n174 ) );
  AOI21_X1 u2_u3_u4_U14 (.ZN( u2_u3_u4_n115 ) , .B2( u2_u3_u4_n145 ) , .B1( u2_u3_u4_n146 ) , .A( u2_u3_u4_n156 ) );
  OAI22_X1 u2_u3_u4_U15 (.ZN( u2_u3_u4_n114 ) , .A2( u2_u3_u4_n121 ) , .B1( u2_u3_u4_n160 ) , .B2( u2_u3_u4_n170 ) , .A1( u2_u3_u4_n171 ) );
  NAND2_X1 u2_u3_u4_U16 (.ZN( u2_u3_u4_n132 ) , .A2( u2_u3_u4_n170 ) , .A1( u2_u3_u4_n173 ) );
  AOI21_X1 u2_u3_u4_U17 (.B2( u2_u3_u4_n160 ) , .B1( u2_u3_u4_n161 ) , .ZN( u2_u3_u4_n162 ) , .A( u2_u3_u4_n170 ) );
  AOI21_X1 u2_u3_u4_U18 (.ZN( u2_u3_u4_n107 ) , .B2( u2_u3_u4_n143 ) , .A( u2_u3_u4_n174 ) , .B1( u2_u3_u4_n184 ) );
  AOI21_X1 u2_u3_u4_U19 (.B2( u2_u3_u4_n158 ) , .B1( u2_u3_u4_n159 ) , .ZN( u2_u3_u4_n163 ) , .A( u2_u3_u4_n174 ) );
  AOI21_X1 u2_u3_u4_U20 (.A( u2_u3_u4_n153 ) , .B2( u2_u3_u4_n154 ) , .B1( u2_u3_u4_n155 ) , .ZN( u2_u3_u4_n165 ) );
  AOI21_X1 u2_u3_u4_U21 (.A( u2_u3_u4_n156 ) , .B2( u2_u3_u4_n157 ) , .ZN( u2_u3_u4_n164 ) , .B1( u2_u3_u4_n184 ) );
  INV_X1 u2_u3_u4_U22 (.A( u2_u3_u4_n138 ) , .ZN( u2_u3_u4_n170 ) );
  AND2_X1 u2_u3_u4_U23 (.A2( u2_u3_u4_n120 ) , .ZN( u2_u3_u4_n155 ) , .A1( u2_u3_u4_n160 ) );
  INV_X1 u2_u3_u4_U24 (.A( u2_u3_u4_n156 ) , .ZN( u2_u3_u4_n175 ) );
  NAND2_X1 u2_u3_u4_U25 (.A2( u2_u3_u4_n118 ) , .ZN( u2_u3_u4_n131 ) , .A1( u2_u3_u4_n147 ) );
  NAND2_X1 u2_u3_u4_U26 (.A1( u2_u3_u4_n119 ) , .A2( u2_u3_u4_n120 ) , .ZN( u2_u3_u4_n130 ) );
  NAND2_X1 u2_u3_u4_U27 (.ZN( u2_u3_u4_n117 ) , .A2( u2_u3_u4_n118 ) , .A1( u2_u3_u4_n148 ) );
  NAND2_X1 u2_u3_u4_U28 (.ZN( u2_u3_u4_n129 ) , .A1( u2_u3_u4_n134 ) , .A2( u2_u3_u4_n148 ) );
  AND3_X1 u2_u3_u4_U29 (.A1( u2_u3_u4_n119 ) , .A2( u2_u3_u4_n143 ) , .A3( u2_u3_u4_n154 ) , .ZN( u2_u3_u4_n161 ) );
  NOR2_X1 u2_u3_u4_U3 (.ZN( u2_u3_u4_n121 ) , .A1( u2_u3_u4_n181 ) , .A2( u2_u3_u4_n182 ) );
  AND2_X1 u2_u3_u4_U30 (.A1( u2_u3_u4_n145 ) , .A2( u2_u3_u4_n147 ) , .ZN( u2_u3_u4_n159 ) );
  INV_X1 u2_u3_u4_U31 (.A( u2_u3_u4_n158 ) , .ZN( u2_u3_u4_n182 ) );
  INV_X1 u2_u3_u4_U32 (.ZN( u2_u3_u4_n181 ) , .A( u2_u3_u4_n96 ) );
  INV_X1 u2_u3_u4_U33 (.A( u2_u3_u4_n144 ) , .ZN( u2_u3_u4_n179 ) );
  INV_X1 u2_u3_u4_U34 (.A( u2_u3_u4_n157 ) , .ZN( u2_u3_u4_n178 ) );
  NAND2_X1 u2_u3_u4_U35 (.A2( u2_u3_u4_n154 ) , .A1( u2_u3_u4_n96 ) , .ZN( u2_u3_u4_n97 ) );
  INV_X1 u2_u3_u4_U36 (.ZN( u2_u3_u4_n186 ) , .A( u2_u3_u4_n95 ) );
  OAI221_X1 u2_u3_u4_U37 (.C1( u2_u3_u4_n134 ) , .B1( u2_u3_u4_n158 ) , .B2( u2_u3_u4_n171 ) , .C2( u2_u3_u4_n173 ) , .A( u2_u3_u4_n94 ) , .ZN( u2_u3_u4_n95 ) );
  AOI222_X1 u2_u3_u4_U38 (.B2( u2_u3_u4_n132 ) , .A1( u2_u3_u4_n138 ) , .C2( u2_u3_u4_n175 ) , .A2( u2_u3_u4_n179 ) , .C1( u2_u3_u4_n181 ) , .B1( u2_u3_u4_n185 ) , .ZN( u2_u3_u4_n94 ) );
  INV_X1 u2_u3_u4_U39 (.A( u2_u3_u4_n113 ) , .ZN( u2_u3_u4_n185 ) );
  INV_X1 u2_u3_u4_U4 (.A( u2_u3_u4_n117 ) , .ZN( u2_u3_u4_n184 ) );
  INV_X1 u2_u3_u4_U40 (.A( u2_u3_u4_n143 ) , .ZN( u2_u3_u4_n183 ) );
  NOR2_X1 u2_u3_u4_U41 (.ZN( u2_u3_u4_n138 ) , .A1( u2_u3_u4_n168 ) , .A2( u2_u3_u4_n169 ) );
  NOR2_X1 u2_u3_u4_U42 (.A1( u2_u3_u4_n150 ) , .A2( u2_u3_u4_n152 ) , .ZN( u2_u3_u4_n153 ) );
  NOR2_X1 u2_u3_u4_U43 (.A2( u2_u3_u4_n128 ) , .A1( u2_u3_u4_n138 ) , .ZN( u2_u3_u4_n156 ) );
  AOI22_X1 u2_u3_u4_U44 (.B2( u2_u3_u4_n122 ) , .A1( u2_u3_u4_n123 ) , .ZN( u2_u3_u4_n124 ) , .B1( u2_u3_u4_n128 ) , .A2( u2_u3_u4_n172 ) );
  INV_X1 u2_u3_u4_U45 (.A( u2_u3_u4_n153 ) , .ZN( u2_u3_u4_n172 ) );
  NAND2_X1 u2_u3_u4_U46 (.A2( u2_u3_u4_n120 ) , .ZN( u2_u3_u4_n123 ) , .A1( u2_u3_u4_n161 ) );
  AOI22_X1 u2_u3_u4_U47 (.B2( u2_u3_u4_n132 ) , .A2( u2_u3_u4_n133 ) , .ZN( u2_u3_u4_n140 ) , .A1( u2_u3_u4_n150 ) , .B1( u2_u3_u4_n179 ) );
  NAND2_X1 u2_u3_u4_U48 (.ZN( u2_u3_u4_n133 ) , .A2( u2_u3_u4_n146 ) , .A1( u2_u3_u4_n154 ) );
  NAND2_X1 u2_u3_u4_U49 (.A1( u2_u3_u4_n103 ) , .ZN( u2_u3_u4_n154 ) , .A2( u2_u3_u4_n98 ) );
  NOR4_X1 u2_u3_u4_U5 (.A4( u2_u3_u4_n106 ) , .A3( u2_u3_u4_n107 ) , .A2( u2_u3_u4_n108 ) , .A1( u2_u3_u4_n109 ) , .ZN( u2_u3_u4_n110 ) );
  NAND2_X1 u2_u3_u4_U50 (.A1( u2_u3_u4_n101 ) , .ZN( u2_u3_u4_n158 ) , .A2( u2_u3_u4_n99 ) );
  AOI21_X1 u2_u3_u4_U51 (.ZN( u2_u3_u4_n127 ) , .A( u2_u3_u4_n136 ) , .B2( u2_u3_u4_n150 ) , .B1( u2_u3_u4_n180 ) );
  INV_X1 u2_u3_u4_U52 (.A( u2_u3_u4_n160 ) , .ZN( u2_u3_u4_n180 ) );
  NAND2_X1 u2_u3_u4_U53 (.A2( u2_u3_u4_n104 ) , .A1( u2_u3_u4_n105 ) , .ZN( u2_u3_u4_n146 ) );
  NAND2_X1 u2_u3_u4_U54 (.A2( u2_u3_u4_n101 ) , .A1( u2_u3_u4_n102 ) , .ZN( u2_u3_u4_n160 ) );
  NAND2_X1 u2_u3_u4_U55 (.ZN( u2_u3_u4_n134 ) , .A1( u2_u3_u4_n98 ) , .A2( u2_u3_u4_n99 ) );
  NAND2_X1 u2_u3_u4_U56 (.A1( u2_u3_u4_n103 ) , .A2( u2_u3_u4_n104 ) , .ZN( u2_u3_u4_n143 ) );
  NAND2_X1 u2_u3_u4_U57 (.A2( u2_u3_u4_n105 ) , .ZN( u2_u3_u4_n145 ) , .A1( u2_u3_u4_n98 ) );
  NAND2_X1 u2_u3_u4_U58 (.A1( u2_u3_u4_n100 ) , .A2( u2_u3_u4_n105 ) , .ZN( u2_u3_u4_n120 ) );
  NAND2_X1 u2_u3_u4_U59 (.A1( u2_u3_u4_n102 ) , .A2( u2_u3_u4_n104 ) , .ZN( u2_u3_u4_n148 ) );
  AOI21_X1 u2_u3_u4_U6 (.ZN( u2_u3_u4_n106 ) , .B2( u2_u3_u4_n146 ) , .B1( u2_u3_u4_n158 ) , .A( u2_u3_u4_n170 ) );
  NAND2_X1 u2_u3_u4_U60 (.A2( u2_u3_u4_n100 ) , .A1( u2_u3_u4_n103 ) , .ZN( u2_u3_u4_n157 ) );
  INV_X1 u2_u3_u4_U61 (.A( u2_u3_u4_n150 ) , .ZN( u2_u3_u4_n173 ) );
  INV_X1 u2_u3_u4_U62 (.A( u2_u3_u4_n152 ) , .ZN( u2_u3_u4_n171 ) );
  NAND2_X1 u2_u3_u4_U63 (.A1( u2_u3_u4_n100 ) , .ZN( u2_u3_u4_n118 ) , .A2( u2_u3_u4_n99 ) );
  NAND2_X1 u2_u3_u4_U64 (.A2( u2_u3_u4_n100 ) , .A1( u2_u3_u4_n102 ) , .ZN( u2_u3_u4_n144 ) );
  NAND2_X1 u2_u3_u4_U65 (.A2( u2_u3_u4_n101 ) , .A1( u2_u3_u4_n105 ) , .ZN( u2_u3_u4_n96 ) );
  INV_X1 u2_u3_u4_U66 (.A( u2_u3_u4_n128 ) , .ZN( u2_u3_u4_n174 ) );
  NAND2_X1 u2_u3_u4_U67 (.A2( u2_u3_u4_n102 ) , .ZN( u2_u3_u4_n119 ) , .A1( u2_u3_u4_n98 ) );
  NAND2_X1 u2_u3_u4_U68 (.A2( u2_u3_u4_n101 ) , .A1( u2_u3_u4_n103 ) , .ZN( u2_u3_u4_n147 ) );
  NAND2_X1 u2_u3_u4_U69 (.A2( u2_u3_u4_n104 ) , .ZN( u2_u3_u4_n113 ) , .A1( u2_u3_u4_n99 ) );
  AOI21_X1 u2_u3_u4_U7 (.ZN( u2_u3_u4_n109 ) , .A( u2_u3_u4_n153 ) , .B1( u2_u3_u4_n159 ) , .B2( u2_u3_u4_n184 ) );
  NOR2_X1 u2_u3_u4_U70 (.A2( u2_u3_X_28 ) , .ZN( u2_u3_u4_n150 ) , .A1( u2_u3_u4_n168 ) );
  NOR2_X1 u2_u3_u4_U71 (.A2( u2_u3_X_29 ) , .ZN( u2_u3_u4_n152 ) , .A1( u2_u3_u4_n169 ) );
  NOR2_X1 u2_u3_u4_U72 (.A2( u2_u3_X_30 ) , .ZN( u2_u3_u4_n105 ) , .A1( u2_u3_u4_n176 ) );
  NOR2_X1 u2_u3_u4_U73 (.A2( u2_u3_X_26 ) , .ZN( u2_u3_u4_n100 ) , .A1( u2_u3_u4_n177 ) );
  NOR2_X1 u2_u3_u4_U74 (.A2( u2_u3_X_28 ) , .A1( u2_u3_X_29 ) , .ZN( u2_u3_u4_n128 ) );
  NOR2_X1 u2_u3_u4_U75 (.A2( u2_u3_X_27 ) , .A1( u2_u3_X_30 ) , .ZN( u2_u3_u4_n102 ) );
  NOR2_X1 u2_u3_u4_U76 (.A2( u2_u3_X_25 ) , .A1( u2_u3_X_26 ) , .ZN( u2_u3_u4_n98 ) );
  AND2_X1 u2_u3_u4_U77 (.A2( u2_u3_X_25 ) , .A1( u2_u3_X_26 ) , .ZN( u2_u3_u4_n104 ) );
  AND2_X1 u2_u3_u4_U78 (.A1( u2_u3_X_30 ) , .A2( u2_u3_u4_n176 ) , .ZN( u2_u3_u4_n99 ) );
  AND2_X1 u2_u3_u4_U79 (.A1( u2_u3_X_26 ) , .ZN( u2_u3_u4_n101 ) , .A2( u2_u3_u4_n177 ) );
  AOI21_X1 u2_u3_u4_U8 (.ZN( u2_u3_u4_n108 ) , .B2( u2_u3_u4_n134 ) , .B1( u2_u3_u4_n155 ) , .A( u2_u3_u4_n156 ) );
  AND2_X1 u2_u3_u4_U80 (.A1( u2_u3_X_27 ) , .A2( u2_u3_X_30 ) , .ZN( u2_u3_u4_n103 ) );
  INV_X1 u2_u3_u4_U81 (.A( u2_u3_X_28 ) , .ZN( u2_u3_u4_n169 ) );
  INV_X1 u2_u3_u4_U82 (.A( u2_u3_X_29 ) , .ZN( u2_u3_u4_n168 ) );
  INV_X1 u2_u3_u4_U83 (.A( u2_u3_X_25 ) , .ZN( u2_u3_u4_n177 ) );
  INV_X1 u2_u3_u4_U84 (.A( u2_u3_X_27 ) , .ZN( u2_u3_u4_n176 ) );
  NAND4_X1 u2_u3_u4_U85 (.ZN( u2_out3_25 ) , .A4( u2_u3_u4_n139 ) , .A3( u2_u3_u4_n140 ) , .A2( u2_u3_u4_n141 ) , .A1( u2_u3_u4_n142 ) );
  OAI21_X1 u2_u3_u4_U86 (.A( u2_u3_u4_n128 ) , .B2( u2_u3_u4_n129 ) , .B1( u2_u3_u4_n130 ) , .ZN( u2_u3_u4_n142 ) );
  OAI21_X1 u2_u3_u4_U87 (.B2( u2_u3_u4_n131 ) , .ZN( u2_u3_u4_n141 ) , .A( u2_u3_u4_n175 ) , .B1( u2_u3_u4_n183 ) );
  NAND4_X1 u2_u3_u4_U88 (.ZN( u2_out3_14 ) , .A4( u2_u3_u4_n124 ) , .A3( u2_u3_u4_n125 ) , .A2( u2_u3_u4_n126 ) , .A1( u2_u3_u4_n127 ) );
  AOI22_X1 u2_u3_u4_U89 (.B2( u2_u3_u4_n117 ) , .ZN( u2_u3_u4_n126 ) , .A1( u2_u3_u4_n129 ) , .B1( u2_u3_u4_n152 ) , .A2( u2_u3_u4_n175 ) );
  AOI211_X1 u2_u3_u4_U9 (.B( u2_u3_u4_n136 ) , .A( u2_u3_u4_n137 ) , .C2( u2_u3_u4_n138 ) , .ZN( u2_u3_u4_n139 ) , .C1( u2_u3_u4_n182 ) );
  AOI22_X1 u2_u3_u4_U90 (.ZN( u2_u3_u4_n125 ) , .B2( u2_u3_u4_n131 ) , .A2( u2_u3_u4_n132 ) , .B1( u2_u3_u4_n138 ) , .A1( u2_u3_u4_n178 ) );
  NAND4_X1 u2_u3_u4_U91 (.ZN( u2_out3_8 ) , .A4( u2_u3_u4_n110 ) , .A3( u2_u3_u4_n111 ) , .A2( u2_u3_u4_n112 ) , .A1( u2_u3_u4_n186 ) );
  NAND2_X1 u2_u3_u4_U92 (.ZN( u2_u3_u4_n112 ) , .A2( u2_u3_u4_n130 ) , .A1( u2_u3_u4_n150 ) );
  AOI22_X1 u2_u3_u4_U93 (.ZN( u2_u3_u4_n111 ) , .B2( u2_u3_u4_n132 ) , .A1( u2_u3_u4_n152 ) , .B1( u2_u3_u4_n178 ) , .A2( u2_u3_u4_n97 ) );
  AOI22_X1 u2_u3_u4_U94 (.B2( u2_u3_u4_n149 ) , .B1( u2_u3_u4_n150 ) , .A2( u2_u3_u4_n151 ) , .A1( u2_u3_u4_n152 ) , .ZN( u2_u3_u4_n167 ) );
  NOR4_X1 u2_u3_u4_U95 (.A4( u2_u3_u4_n162 ) , .A3( u2_u3_u4_n163 ) , .A2( u2_u3_u4_n164 ) , .A1( u2_u3_u4_n165 ) , .ZN( u2_u3_u4_n166 ) );
  NAND3_X1 u2_u3_u4_U96 (.ZN( u2_out3_3 ) , .A3( u2_u3_u4_n166 ) , .A1( u2_u3_u4_n167 ) , .A2( u2_u3_u4_n186 ) );
  NAND3_X1 u2_u3_u4_U97 (.A3( u2_u3_u4_n146 ) , .A2( u2_u3_u4_n147 ) , .A1( u2_u3_u4_n148 ) , .ZN( u2_u3_u4_n149 ) );
  NAND3_X1 u2_u3_u4_U98 (.A3( u2_u3_u4_n143 ) , .A2( u2_u3_u4_n144 ) , .A1( u2_u3_u4_n145 ) , .ZN( u2_u3_u4_n151 ) );
  NAND3_X1 u2_u3_u4_U99 (.A3( u2_u3_u4_n121 ) , .ZN( u2_u3_u4_n122 ) , .A2( u2_u3_u4_n144 ) , .A1( u2_u3_u4_n154 ) );
  INV_X1 u2_u3_u5_U10 (.A( u2_u3_u5_n121 ) , .ZN( u2_u3_u5_n177 ) );
  NOR3_X1 u2_u3_u5_U100 (.A3( u2_u3_u5_n141 ) , .A1( u2_u3_u5_n142 ) , .ZN( u2_u3_u5_n143 ) , .A2( u2_u3_u5_n191 ) );
  NAND4_X1 u2_u3_u5_U101 (.ZN( u2_out3_4 ) , .A4( u2_u3_u5_n112 ) , .A2( u2_u3_u5_n113 ) , .A1( u2_u3_u5_n114 ) , .A3( u2_u3_u5_n195 ) );
  AOI211_X1 u2_u3_u5_U102 (.A( u2_u3_u5_n110 ) , .C1( u2_u3_u5_n111 ) , .ZN( u2_u3_u5_n112 ) , .B( u2_u3_u5_n118 ) , .C2( u2_u3_u5_n177 ) );
  AOI222_X1 u2_u3_u5_U103 (.ZN( u2_u3_u5_n113 ) , .A1( u2_u3_u5_n131 ) , .C1( u2_u3_u5_n148 ) , .B2( u2_u3_u5_n174 ) , .C2( u2_u3_u5_n178 ) , .A2( u2_u3_u5_n179 ) , .B1( u2_u3_u5_n99 ) );
  NAND3_X1 u2_u3_u5_U104 (.A2( u2_u3_u5_n154 ) , .A3( u2_u3_u5_n158 ) , .A1( u2_u3_u5_n161 ) , .ZN( u2_u3_u5_n99 ) );
  NOR2_X1 u2_u3_u5_U11 (.ZN( u2_u3_u5_n160 ) , .A2( u2_u3_u5_n173 ) , .A1( u2_u3_u5_n177 ) );
  INV_X1 u2_u3_u5_U12 (.A( u2_u3_u5_n150 ) , .ZN( u2_u3_u5_n174 ) );
  AOI21_X1 u2_u3_u5_U13 (.A( u2_u3_u5_n160 ) , .B2( u2_u3_u5_n161 ) , .ZN( u2_u3_u5_n162 ) , .B1( u2_u3_u5_n192 ) );
  INV_X1 u2_u3_u5_U14 (.A( u2_u3_u5_n159 ) , .ZN( u2_u3_u5_n192 ) );
  AOI21_X1 u2_u3_u5_U15 (.A( u2_u3_u5_n156 ) , .B2( u2_u3_u5_n157 ) , .B1( u2_u3_u5_n158 ) , .ZN( u2_u3_u5_n163 ) );
  AOI21_X1 u2_u3_u5_U16 (.B2( u2_u3_u5_n139 ) , .B1( u2_u3_u5_n140 ) , .ZN( u2_u3_u5_n141 ) , .A( u2_u3_u5_n150 ) );
  OAI21_X1 u2_u3_u5_U17 (.A( u2_u3_u5_n133 ) , .B2( u2_u3_u5_n134 ) , .B1( u2_u3_u5_n135 ) , .ZN( u2_u3_u5_n142 ) );
  OAI21_X1 u2_u3_u5_U18 (.ZN( u2_u3_u5_n133 ) , .B2( u2_u3_u5_n147 ) , .A( u2_u3_u5_n173 ) , .B1( u2_u3_u5_n188 ) );
  NAND2_X1 u2_u3_u5_U19 (.A2( u2_u3_u5_n119 ) , .A1( u2_u3_u5_n123 ) , .ZN( u2_u3_u5_n137 ) );
  INV_X1 u2_u3_u5_U20 (.A( u2_u3_u5_n155 ) , .ZN( u2_u3_u5_n194 ) );
  NAND2_X1 u2_u3_u5_U21 (.A1( u2_u3_u5_n121 ) , .ZN( u2_u3_u5_n132 ) , .A2( u2_u3_u5_n172 ) );
  NAND2_X1 u2_u3_u5_U22 (.A2( u2_u3_u5_n122 ) , .ZN( u2_u3_u5_n136 ) , .A1( u2_u3_u5_n154 ) );
  NAND2_X1 u2_u3_u5_U23 (.A2( u2_u3_u5_n119 ) , .A1( u2_u3_u5_n120 ) , .ZN( u2_u3_u5_n159 ) );
  INV_X1 u2_u3_u5_U24 (.A( u2_u3_u5_n156 ) , .ZN( u2_u3_u5_n175 ) );
  INV_X1 u2_u3_u5_U25 (.A( u2_u3_u5_n158 ) , .ZN( u2_u3_u5_n188 ) );
  INV_X1 u2_u3_u5_U26 (.A( u2_u3_u5_n152 ) , .ZN( u2_u3_u5_n179 ) );
  INV_X1 u2_u3_u5_U27 (.A( u2_u3_u5_n140 ) , .ZN( u2_u3_u5_n182 ) );
  INV_X1 u2_u3_u5_U28 (.A( u2_u3_u5_n151 ) , .ZN( u2_u3_u5_n183 ) );
  INV_X1 u2_u3_u5_U29 (.A( u2_u3_u5_n123 ) , .ZN( u2_u3_u5_n185 ) );
  NOR2_X1 u2_u3_u5_U3 (.ZN( u2_u3_u5_n134 ) , .A1( u2_u3_u5_n183 ) , .A2( u2_u3_u5_n190 ) );
  INV_X1 u2_u3_u5_U30 (.A( u2_u3_u5_n161 ) , .ZN( u2_u3_u5_n184 ) );
  INV_X1 u2_u3_u5_U31 (.A( u2_u3_u5_n139 ) , .ZN( u2_u3_u5_n189 ) );
  INV_X1 u2_u3_u5_U32 (.A( u2_u3_u5_n157 ) , .ZN( u2_u3_u5_n190 ) );
  INV_X1 u2_u3_u5_U33 (.A( u2_u3_u5_n120 ) , .ZN( u2_u3_u5_n193 ) );
  NAND2_X1 u2_u3_u5_U34 (.ZN( u2_u3_u5_n111 ) , .A1( u2_u3_u5_n140 ) , .A2( u2_u3_u5_n155 ) );
  INV_X1 u2_u3_u5_U35 (.A( u2_u3_u5_n117 ) , .ZN( u2_u3_u5_n196 ) );
  OAI221_X1 u2_u3_u5_U36 (.A( u2_u3_u5_n116 ) , .ZN( u2_u3_u5_n117 ) , .B2( u2_u3_u5_n119 ) , .C1( u2_u3_u5_n153 ) , .C2( u2_u3_u5_n158 ) , .B1( u2_u3_u5_n172 ) );
  AOI222_X1 u2_u3_u5_U37 (.ZN( u2_u3_u5_n116 ) , .B2( u2_u3_u5_n145 ) , .C1( u2_u3_u5_n148 ) , .A2( u2_u3_u5_n174 ) , .C2( u2_u3_u5_n177 ) , .B1( u2_u3_u5_n187 ) , .A1( u2_u3_u5_n193 ) );
  INV_X1 u2_u3_u5_U38 (.A( u2_u3_u5_n115 ) , .ZN( u2_u3_u5_n187 ) );
  NOR2_X1 u2_u3_u5_U39 (.ZN( u2_u3_u5_n100 ) , .A1( u2_u3_u5_n170 ) , .A2( u2_u3_u5_n180 ) );
  INV_X1 u2_u3_u5_U4 (.A( u2_u3_u5_n138 ) , .ZN( u2_u3_u5_n191 ) );
  AOI22_X1 u2_u3_u5_U40 (.B2( u2_u3_u5_n131 ) , .A2( u2_u3_u5_n146 ) , .ZN( u2_u3_u5_n169 ) , .B1( u2_u3_u5_n174 ) , .A1( u2_u3_u5_n185 ) );
  NOR2_X1 u2_u3_u5_U41 (.A1( u2_u3_u5_n146 ) , .ZN( u2_u3_u5_n150 ) , .A2( u2_u3_u5_n173 ) );
  AOI21_X1 u2_u3_u5_U42 (.A( u2_u3_u5_n118 ) , .B2( u2_u3_u5_n145 ) , .ZN( u2_u3_u5_n168 ) , .B1( u2_u3_u5_n186 ) );
  INV_X1 u2_u3_u5_U43 (.A( u2_u3_u5_n122 ) , .ZN( u2_u3_u5_n186 ) );
  NOR2_X1 u2_u3_u5_U44 (.A1( u2_u3_u5_n146 ) , .ZN( u2_u3_u5_n152 ) , .A2( u2_u3_u5_n176 ) );
  NOR2_X1 u2_u3_u5_U45 (.A1( u2_u3_u5_n115 ) , .ZN( u2_u3_u5_n118 ) , .A2( u2_u3_u5_n153 ) );
  NOR2_X1 u2_u3_u5_U46 (.A2( u2_u3_u5_n145 ) , .ZN( u2_u3_u5_n156 ) , .A1( u2_u3_u5_n174 ) );
  NOR2_X1 u2_u3_u5_U47 (.ZN( u2_u3_u5_n121 ) , .A2( u2_u3_u5_n145 ) , .A1( u2_u3_u5_n176 ) );
  AOI22_X1 u2_u3_u5_U48 (.ZN( u2_u3_u5_n114 ) , .A2( u2_u3_u5_n137 ) , .A1( u2_u3_u5_n145 ) , .B2( u2_u3_u5_n175 ) , .B1( u2_u3_u5_n193 ) );
  OAI211_X1 u2_u3_u5_U49 (.B( u2_u3_u5_n124 ) , .A( u2_u3_u5_n125 ) , .C2( u2_u3_u5_n126 ) , .C1( u2_u3_u5_n127 ) , .ZN( u2_u3_u5_n128 ) );
  OAI21_X1 u2_u3_u5_U5 (.B2( u2_u3_u5_n136 ) , .B1( u2_u3_u5_n137 ) , .ZN( u2_u3_u5_n138 ) , .A( u2_u3_u5_n177 ) );
  NOR3_X1 u2_u3_u5_U50 (.ZN( u2_u3_u5_n127 ) , .A1( u2_u3_u5_n136 ) , .A3( u2_u3_u5_n148 ) , .A2( u2_u3_u5_n182 ) );
  OAI21_X1 u2_u3_u5_U51 (.ZN( u2_u3_u5_n124 ) , .A( u2_u3_u5_n177 ) , .B2( u2_u3_u5_n183 ) , .B1( u2_u3_u5_n189 ) );
  OAI21_X1 u2_u3_u5_U52 (.ZN( u2_u3_u5_n125 ) , .A( u2_u3_u5_n174 ) , .B2( u2_u3_u5_n185 ) , .B1( u2_u3_u5_n190 ) );
  AOI21_X1 u2_u3_u5_U53 (.A( u2_u3_u5_n153 ) , .B2( u2_u3_u5_n154 ) , .B1( u2_u3_u5_n155 ) , .ZN( u2_u3_u5_n164 ) );
  AOI21_X1 u2_u3_u5_U54 (.ZN( u2_u3_u5_n110 ) , .B1( u2_u3_u5_n122 ) , .B2( u2_u3_u5_n139 ) , .A( u2_u3_u5_n153 ) );
  INV_X1 u2_u3_u5_U55 (.A( u2_u3_u5_n153 ) , .ZN( u2_u3_u5_n176 ) );
  INV_X1 u2_u3_u5_U56 (.A( u2_u3_u5_n126 ) , .ZN( u2_u3_u5_n173 ) );
  AND2_X1 u2_u3_u5_U57 (.A2( u2_u3_u5_n104 ) , .A1( u2_u3_u5_n107 ) , .ZN( u2_u3_u5_n147 ) );
  AND2_X1 u2_u3_u5_U58 (.A2( u2_u3_u5_n104 ) , .A1( u2_u3_u5_n108 ) , .ZN( u2_u3_u5_n148 ) );
  NAND2_X1 u2_u3_u5_U59 (.A1( u2_u3_u5_n105 ) , .A2( u2_u3_u5_n106 ) , .ZN( u2_u3_u5_n158 ) );
  INV_X1 u2_u3_u5_U6 (.A( u2_u3_u5_n135 ) , .ZN( u2_u3_u5_n178 ) );
  NAND2_X1 u2_u3_u5_U60 (.A2( u2_u3_u5_n108 ) , .A1( u2_u3_u5_n109 ) , .ZN( u2_u3_u5_n139 ) );
  NAND2_X1 u2_u3_u5_U61 (.A1( u2_u3_u5_n106 ) , .A2( u2_u3_u5_n108 ) , .ZN( u2_u3_u5_n119 ) );
  NAND2_X1 u2_u3_u5_U62 (.A2( u2_u3_u5_n103 ) , .A1( u2_u3_u5_n105 ) , .ZN( u2_u3_u5_n140 ) );
  NAND2_X1 u2_u3_u5_U63 (.A2( u2_u3_u5_n104 ) , .A1( u2_u3_u5_n105 ) , .ZN( u2_u3_u5_n155 ) );
  NAND2_X1 u2_u3_u5_U64 (.A2( u2_u3_u5_n106 ) , .A1( u2_u3_u5_n107 ) , .ZN( u2_u3_u5_n122 ) );
  NAND2_X1 u2_u3_u5_U65 (.A2( u2_u3_u5_n100 ) , .A1( u2_u3_u5_n106 ) , .ZN( u2_u3_u5_n115 ) );
  NAND2_X1 u2_u3_u5_U66 (.A2( u2_u3_u5_n100 ) , .A1( u2_u3_u5_n103 ) , .ZN( u2_u3_u5_n161 ) );
  NAND2_X1 u2_u3_u5_U67 (.A1( u2_u3_u5_n105 ) , .A2( u2_u3_u5_n109 ) , .ZN( u2_u3_u5_n154 ) );
  INV_X1 u2_u3_u5_U68 (.A( u2_u3_u5_n146 ) , .ZN( u2_u3_u5_n172 ) );
  NAND2_X1 u2_u3_u5_U69 (.A1( u2_u3_u5_n103 ) , .A2( u2_u3_u5_n108 ) , .ZN( u2_u3_u5_n123 ) );
  OAI22_X1 u2_u3_u5_U7 (.B2( u2_u3_u5_n149 ) , .B1( u2_u3_u5_n150 ) , .A2( u2_u3_u5_n151 ) , .A1( u2_u3_u5_n152 ) , .ZN( u2_u3_u5_n165 ) );
  NAND2_X1 u2_u3_u5_U70 (.A2( u2_u3_u5_n103 ) , .A1( u2_u3_u5_n107 ) , .ZN( u2_u3_u5_n151 ) );
  NAND2_X1 u2_u3_u5_U71 (.A2( u2_u3_u5_n107 ) , .A1( u2_u3_u5_n109 ) , .ZN( u2_u3_u5_n120 ) );
  NAND2_X1 u2_u3_u5_U72 (.A2( u2_u3_u5_n100 ) , .A1( u2_u3_u5_n109 ) , .ZN( u2_u3_u5_n157 ) );
  AND2_X1 u2_u3_u5_U73 (.A2( u2_u3_u5_n100 ) , .A1( u2_u3_u5_n104 ) , .ZN( u2_u3_u5_n131 ) );
  INV_X1 u2_u3_u5_U74 (.A( u2_u3_u5_n102 ) , .ZN( u2_u3_u5_n195 ) );
  OAI221_X1 u2_u3_u5_U75 (.A( u2_u3_u5_n101 ) , .ZN( u2_u3_u5_n102 ) , .C2( u2_u3_u5_n115 ) , .C1( u2_u3_u5_n126 ) , .B1( u2_u3_u5_n134 ) , .B2( u2_u3_u5_n160 ) );
  OAI21_X1 u2_u3_u5_U76 (.ZN( u2_u3_u5_n101 ) , .B1( u2_u3_u5_n137 ) , .A( u2_u3_u5_n146 ) , .B2( u2_u3_u5_n147 ) );
  NOR2_X1 u2_u3_u5_U77 (.A2( u2_u3_X_34 ) , .A1( u2_u3_X_35 ) , .ZN( u2_u3_u5_n145 ) );
  NOR2_X1 u2_u3_u5_U78 (.A2( u2_u3_X_34 ) , .ZN( u2_u3_u5_n146 ) , .A1( u2_u3_u5_n171 ) );
  NOR2_X1 u2_u3_u5_U79 (.A2( u2_u3_X_31 ) , .A1( u2_u3_X_32 ) , .ZN( u2_u3_u5_n103 ) );
  NOR3_X1 u2_u3_u5_U8 (.A2( u2_u3_u5_n147 ) , .A1( u2_u3_u5_n148 ) , .ZN( u2_u3_u5_n149 ) , .A3( u2_u3_u5_n194 ) );
  NOR2_X1 u2_u3_u5_U80 (.A2( u2_u3_X_36 ) , .ZN( u2_u3_u5_n105 ) , .A1( u2_u3_u5_n180 ) );
  NOR2_X1 u2_u3_u5_U81 (.A2( u2_u3_X_33 ) , .ZN( u2_u3_u5_n108 ) , .A1( u2_u3_u5_n170 ) );
  NOR2_X1 u2_u3_u5_U82 (.A2( u2_u3_X_33 ) , .A1( u2_u3_X_36 ) , .ZN( u2_u3_u5_n107 ) );
  NOR2_X1 u2_u3_u5_U83 (.A2( u2_u3_X_31 ) , .ZN( u2_u3_u5_n104 ) , .A1( u2_u3_u5_n181 ) );
  NAND2_X1 u2_u3_u5_U84 (.A2( u2_u3_X_34 ) , .A1( u2_u3_X_35 ) , .ZN( u2_u3_u5_n153 ) );
  NAND2_X1 u2_u3_u5_U85 (.A1( u2_u3_X_34 ) , .ZN( u2_u3_u5_n126 ) , .A2( u2_u3_u5_n171 ) );
  AND2_X1 u2_u3_u5_U86 (.A1( u2_u3_X_31 ) , .A2( u2_u3_X_32 ) , .ZN( u2_u3_u5_n106 ) );
  AND2_X1 u2_u3_u5_U87 (.A1( u2_u3_X_31 ) , .ZN( u2_u3_u5_n109 ) , .A2( u2_u3_u5_n181 ) );
  INV_X1 u2_u3_u5_U88 (.A( u2_u3_X_33 ) , .ZN( u2_u3_u5_n180 ) );
  INV_X1 u2_u3_u5_U89 (.A( u2_u3_X_35 ) , .ZN( u2_u3_u5_n171 ) );
  NOR2_X1 u2_u3_u5_U9 (.ZN( u2_u3_u5_n135 ) , .A1( u2_u3_u5_n173 ) , .A2( u2_u3_u5_n176 ) );
  INV_X1 u2_u3_u5_U90 (.A( u2_u3_X_36 ) , .ZN( u2_u3_u5_n170 ) );
  INV_X1 u2_u3_u5_U91 (.A( u2_u3_X_32 ) , .ZN( u2_u3_u5_n181 ) );
  NAND4_X1 u2_u3_u5_U92 (.ZN( u2_out3_29 ) , .A4( u2_u3_u5_n129 ) , .A3( u2_u3_u5_n130 ) , .A2( u2_u3_u5_n168 ) , .A1( u2_u3_u5_n196 ) );
  AOI221_X1 u2_u3_u5_U93 (.A( u2_u3_u5_n128 ) , .ZN( u2_u3_u5_n129 ) , .C2( u2_u3_u5_n132 ) , .B2( u2_u3_u5_n159 ) , .B1( u2_u3_u5_n176 ) , .C1( u2_u3_u5_n184 ) );
  AOI222_X1 u2_u3_u5_U94 (.ZN( u2_u3_u5_n130 ) , .A2( u2_u3_u5_n146 ) , .B1( u2_u3_u5_n147 ) , .C2( u2_u3_u5_n175 ) , .B2( u2_u3_u5_n179 ) , .A1( u2_u3_u5_n188 ) , .C1( u2_u3_u5_n194 ) );
  NAND4_X1 u2_u3_u5_U95 (.ZN( u2_out3_19 ) , .A4( u2_u3_u5_n166 ) , .A3( u2_u3_u5_n167 ) , .A2( u2_u3_u5_n168 ) , .A1( u2_u3_u5_n169 ) );
  AOI22_X1 u2_u3_u5_U96 (.B2( u2_u3_u5_n145 ) , .A2( u2_u3_u5_n146 ) , .ZN( u2_u3_u5_n167 ) , .B1( u2_u3_u5_n182 ) , .A1( u2_u3_u5_n189 ) );
  NOR4_X1 u2_u3_u5_U97 (.A4( u2_u3_u5_n162 ) , .A3( u2_u3_u5_n163 ) , .A2( u2_u3_u5_n164 ) , .A1( u2_u3_u5_n165 ) , .ZN( u2_u3_u5_n166 ) );
  NAND4_X1 u2_u3_u5_U98 (.ZN( u2_out3_11 ) , .A4( u2_u3_u5_n143 ) , .A3( u2_u3_u5_n144 ) , .A2( u2_u3_u5_n169 ) , .A1( u2_u3_u5_n196 ) );
  AOI22_X1 u2_u3_u5_U99 (.A2( u2_u3_u5_n132 ) , .ZN( u2_u3_u5_n144 ) , .B2( u2_u3_u5_n145 ) , .B1( u2_u3_u5_n184 ) , .A1( u2_u3_u5_n194 ) );
  INV_X1 u2_u3_u6_U10 (.ZN( u2_u3_u6_n172 ) , .A( u2_u3_u6_n88 ) );
  OAI21_X1 u2_u3_u6_U11 (.A( u2_u3_u6_n159 ) , .B1( u2_u3_u6_n169 ) , .B2( u2_u3_u6_n173 ) , .ZN( u2_u3_u6_n90 ) );
  AOI22_X1 u2_u3_u6_U12 (.A2( u2_u3_u6_n151 ) , .B2( u2_u3_u6_n161 ) , .A1( u2_u3_u6_n167 ) , .B1( u2_u3_u6_n170 ) , .ZN( u2_u3_u6_n89 ) );
  AOI21_X1 u2_u3_u6_U13 (.ZN( u2_u3_u6_n106 ) , .A( u2_u3_u6_n142 ) , .B2( u2_u3_u6_n159 ) , .B1( u2_u3_u6_n164 ) );
  INV_X1 u2_u3_u6_U14 (.A( u2_u3_u6_n155 ) , .ZN( u2_u3_u6_n161 ) );
  INV_X1 u2_u3_u6_U15 (.A( u2_u3_u6_n128 ) , .ZN( u2_u3_u6_n164 ) );
  NAND2_X1 u2_u3_u6_U16 (.ZN( u2_u3_u6_n110 ) , .A1( u2_u3_u6_n122 ) , .A2( u2_u3_u6_n129 ) );
  NAND2_X1 u2_u3_u6_U17 (.ZN( u2_u3_u6_n124 ) , .A2( u2_u3_u6_n146 ) , .A1( u2_u3_u6_n148 ) );
  INV_X1 u2_u3_u6_U18 (.A( u2_u3_u6_n132 ) , .ZN( u2_u3_u6_n171 ) );
  AND2_X1 u2_u3_u6_U19 (.A1( u2_u3_u6_n100 ) , .ZN( u2_u3_u6_n130 ) , .A2( u2_u3_u6_n147 ) );
  INV_X1 u2_u3_u6_U20 (.A( u2_u3_u6_n127 ) , .ZN( u2_u3_u6_n173 ) );
  INV_X1 u2_u3_u6_U21 (.A( u2_u3_u6_n121 ) , .ZN( u2_u3_u6_n167 ) );
  INV_X1 u2_u3_u6_U22 (.A( u2_u3_u6_n100 ) , .ZN( u2_u3_u6_n169 ) );
  INV_X1 u2_u3_u6_U23 (.A( u2_u3_u6_n123 ) , .ZN( u2_u3_u6_n170 ) );
  INV_X1 u2_u3_u6_U24 (.A( u2_u3_u6_n113 ) , .ZN( u2_u3_u6_n168 ) );
  AND2_X1 u2_u3_u6_U25 (.A1( u2_u3_u6_n107 ) , .A2( u2_u3_u6_n119 ) , .ZN( u2_u3_u6_n133 ) );
  AND2_X1 u2_u3_u6_U26 (.A2( u2_u3_u6_n121 ) , .A1( u2_u3_u6_n122 ) , .ZN( u2_u3_u6_n131 ) );
  AND3_X1 u2_u3_u6_U27 (.ZN( u2_u3_u6_n120 ) , .A2( u2_u3_u6_n127 ) , .A1( u2_u3_u6_n132 ) , .A3( u2_u3_u6_n145 ) );
  INV_X1 u2_u3_u6_U28 (.A( u2_u3_u6_n146 ) , .ZN( u2_u3_u6_n163 ) );
  AOI222_X1 u2_u3_u6_U29 (.ZN( u2_u3_u6_n114 ) , .A1( u2_u3_u6_n118 ) , .A2( u2_u3_u6_n126 ) , .B2( u2_u3_u6_n151 ) , .C2( u2_u3_u6_n159 ) , .C1( u2_u3_u6_n168 ) , .B1( u2_u3_u6_n169 ) );
  INV_X1 u2_u3_u6_U3 (.A( u2_u3_u6_n110 ) , .ZN( u2_u3_u6_n166 ) );
  NOR2_X1 u2_u3_u6_U30 (.A1( u2_u3_u6_n162 ) , .A2( u2_u3_u6_n165 ) , .ZN( u2_u3_u6_n98 ) );
  NAND2_X1 u2_u3_u6_U31 (.A1( u2_u3_u6_n144 ) , .ZN( u2_u3_u6_n151 ) , .A2( u2_u3_u6_n158 ) );
  NAND2_X1 u2_u3_u6_U32 (.ZN( u2_u3_u6_n132 ) , .A1( u2_u3_u6_n91 ) , .A2( u2_u3_u6_n97 ) );
  AOI22_X1 u2_u3_u6_U33 (.B2( u2_u3_u6_n110 ) , .B1( u2_u3_u6_n111 ) , .A1( u2_u3_u6_n112 ) , .ZN( u2_u3_u6_n115 ) , .A2( u2_u3_u6_n161 ) );
  NAND4_X1 u2_u3_u6_U34 (.A3( u2_u3_u6_n109 ) , .ZN( u2_u3_u6_n112 ) , .A4( u2_u3_u6_n132 ) , .A2( u2_u3_u6_n147 ) , .A1( u2_u3_u6_n166 ) );
  NOR2_X1 u2_u3_u6_U35 (.ZN( u2_u3_u6_n109 ) , .A1( u2_u3_u6_n170 ) , .A2( u2_u3_u6_n173 ) );
  NOR2_X1 u2_u3_u6_U36 (.A2( u2_u3_u6_n126 ) , .ZN( u2_u3_u6_n155 ) , .A1( u2_u3_u6_n160 ) );
  NAND2_X1 u2_u3_u6_U37 (.ZN( u2_u3_u6_n146 ) , .A2( u2_u3_u6_n94 ) , .A1( u2_u3_u6_n99 ) );
  AOI21_X1 u2_u3_u6_U38 (.A( u2_u3_u6_n144 ) , .B2( u2_u3_u6_n145 ) , .B1( u2_u3_u6_n146 ) , .ZN( u2_u3_u6_n150 ) );
  AOI211_X1 u2_u3_u6_U39 (.B( u2_u3_u6_n134 ) , .A( u2_u3_u6_n135 ) , .C1( u2_u3_u6_n136 ) , .ZN( u2_u3_u6_n137 ) , .C2( u2_u3_u6_n151 ) );
  INV_X1 u2_u3_u6_U4 (.A( u2_u3_u6_n142 ) , .ZN( u2_u3_u6_n174 ) );
  AOI21_X1 u2_u3_u6_U40 (.B2( u2_u3_u6_n132 ) , .B1( u2_u3_u6_n133 ) , .ZN( u2_u3_u6_n134 ) , .A( u2_u3_u6_n158 ) );
  NAND4_X1 u2_u3_u6_U41 (.A4( u2_u3_u6_n127 ) , .A3( u2_u3_u6_n128 ) , .A2( u2_u3_u6_n129 ) , .A1( u2_u3_u6_n130 ) , .ZN( u2_u3_u6_n136 ) );
  AOI21_X1 u2_u3_u6_U42 (.B1( u2_u3_u6_n131 ) , .ZN( u2_u3_u6_n135 ) , .A( u2_u3_u6_n144 ) , .B2( u2_u3_u6_n146 ) );
  INV_X1 u2_u3_u6_U43 (.A( u2_u3_u6_n111 ) , .ZN( u2_u3_u6_n158 ) );
  NAND2_X1 u2_u3_u6_U44 (.ZN( u2_u3_u6_n127 ) , .A1( u2_u3_u6_n91 ) , .A2( u2_u3_u6_n92 ) );
  NAND2_X1 u2_u3_u6_U45 (.ZN( u2_u3_u6_n129 ) , .A2( u2_u3_u6_n95 ) , .A1( u2_u3_u6_n96 ) );
  INV_X1 u2_u3_u6_U46 (.A( u2_u3_u6_n144 ) , .ZN( u2_u3_u6_n159 ) );
  NAND2_X1 u2_u3_u6_U47 (.ZN( u2_u3_u6_n145 ) , .A2( u2_u3_u6_n97 ) , .A1( u2_u3_u6_n98 ) );
  NAND2_X1 u2_u3_u6_U48 (.ZN( u2_u3_u6_n148 ) , .A2( u2_u3_u6_n92 ) , .A1( u2_u3_u6_n94 ) );
  NAND2_X1 u2_u3_u6_U49 (.ZN( u2_u3_u6_n108 ) , .A2( u2_u3_u6_n139 ) , .A1( u2_u3_u6_n144 ) );
  NAND2_X1 u2_u3_u6_U5 (.A2( u2_u3_u6_n143 ) , .ZN( u2_u3_u6_n152 ) , .A1( u2_u3_u6_n166 ) );
  NAND2_X1 u2_u3_u6_U50 (.ZN( u2_u3_u6_n121 ) , .A2( u2_u3_u6_n95 ) , .A1( u2_u3_u6_n97 ) );
  NAND2_X1 u2_u3_u6_U51 (.ZN( u2_u3_u6_n107 ) , .A2( u2_u3_u6_n92 ) , .A1( u2_u3_u6_n95 ) );
  AND2_X1 u2_u3_u6_U52 (.ZN( u2_u3_u6_n118 ) , .A2( u2_u3_u6_n91 ) , .A1( u2_u3_u6_n99 ) );
  NAND2_X1 u2_u3_u6_U53 (.ZN( u2_u3_u6_n147 ) , .A2( u2_u3_u6_n98 ) , .A1( u2_u3_u6_n99 ) );
  NAND2_X1 u2_u3_u6_U54 (.ZN( u2_u3_u6_n128 ) , .A1( u2_u3_u6_n94 ) , .A2( u2_u3_u6_n96 ) );
  NAND2_X1 u2_u3_u6_U55 (.ZN( u2_u3_u6_n119 ) , .A2( u2_u3_u6_n95 ) , .A1( u2_u3_u6_n99 ) );
  NAND2_X1 u2_u3_u6_U56 (.ZN( u2_u3_u6_n123 ) , .A2( u2_u3_u6_n91 ) , .A1( u2_u3_u6_n96 ) );
  NAND2_X1 u2_u3_u6_U57 (.ZN( u2_u3_u6_n100 ) , .A2( u2_u3_u6_n92 ) , .A1( u2_u3_u6_n98 ) );
  NAND2_X1 u2_u3_u6_U58 (.ZN( u2_u3_u6_n122 ) , .A1( u2_u3_u6_n94 ) , .A2( u2_u3_u6_n97 ) );
  INV_X1 u2_u3_u6_U59 (.A( u2_u3_u6_n139 ) , .ZN( u2_u3_u6_n160 ) );
  AOI22_X1 u2_u3_u6_U6 (.B2( u2_u3_u6_n101 ) , .A1( u2_u3_u6_n102 ) , .ZN( u2_u3_u6_n103 ) , .B1( u2_u3_u6_n160 ) , .A2( u2_u3_u6_n161 ) );
  NAND2_X1 u2_u3_u6_U60 (.ZN( u2_u3_u6_n113 ) , .A1( u2_u3_u6_n96 ) , .A2( u2_u3_u6_n98 ) );
  NOR2_X1 u2_u3_u6_U61 (.A2( u2_u3_X_40 ) , .A1( u2_u3_X_41 ) , .ZN( u2_u3_u6_n126 ) );
  NOR2_X1 u2_u3_u6_U62 (.A2( u2_u3_X_39 ) , .A1( u2_u3_X_42 ) , .ZN( u2_u3_u6_n92 ) );
  NOR2_X1 u2_u3_u6_U63 (.A2( u2_u3_X_39 ) , .A1( u2_u3_u6_n156 ) , .ZN( u2_u3_u6_n97 ) );
  NOR2_X1 u2_u3_u6_U64 (.A2( u2_u3_X_38 ) , .A1( u2_u3_u6_n165 ) , .ZN( u2_u3_u6_n95 ) );
  NOR2_X1 u2_u3_u6_U65 (.A2( u2_u3_X_41 ) , .ZN( u2_u3_u6_n111 ) , .A1( u2_u3_u6_n157 ) );
  NOR2_X1 u2_u3_u6_U66 (.A2( u2_u3_X_37 ) , .A1( u2_u3_u6_n162 ) , .ZN( u2_u3_u6_n94 ) );
  NOR2_X1 u2_u3_u6_U67 (.A2( u2_u3_X_37 ) , .A1( u2_u3_X_38 ) , .ZN( u2_u3_u6_n91 ) );
  NAND2_X1 u2_u3_u6_U68 (.A1( u2_u3_X_41 ) , .ZN( u2_u3_u6_n144 ) , .A2( u2_u3_u6_n157 ) );
  NAND2_X1 u2_u3_u6_U69 (.A2( u2_u3_X_40 ) , .A1( u2_u3_X_41 ) , .ZN( u2_u3_u6_n139 ) );
  NOR2_X1 u2_u3_u6_U7 (.A1( u2_u3_u6_n118 ) , .ZN( u2_u3_u6_n143 ) , .A2( u2_u3_u6_n168 ) );
  AND2_X1 u2_u3_u6_U70 (.A1( u2_u3_X_39 ) , .A2( u2_u3_u6_n156 ) , .ZN( u2_u3_u6_n96 ) );
  AND2_X1 u2_u3_u6_U71 (.A1( u2_u3_X_39 ) , .A2( u2_u3_X_42 ) , .ZN( u2_u3_u6_n99 ) );
  INV_X1 u2_u3_u6_U72 (.A( u2_u3_X_40 ) , .ZN( u2_u3_u6_n157 ) );
  INV_X1 u2_u3_u6_U73 (.A( u2_u3_X_37 ) , .ZN( u2_u3_u6_n165 ) );
  INV_X1 u2_u3_u6_U74 (.A( u2_u3_X_38 ) , .ZN( u2_u3_u6_n162 ) );
  INV_X1 u2_u3_u6_U75 (.A( u2_u3_X_42 ) , .ZN( u2_u3_u6_n156 ) );
  NAND4_X1 u2_u3_u6_U76 (.ZN( u2_out3_32 ) , .A4( u2_u3_u6_n103 ) , .A3( u2_u3_u6_n104 ) , .A2( u2_u3_u6_n105 ) , .A1( u2_u3_u6_n106 ) );
  AOI22_X1 u2_u3_u6_U77 (.ZN( u2_u3_u6_n105 ) , .A2( u2_u3_u6_n108 ) , .A1( u2_u3_u6_n118 ) , .B2( u2_u3_u6_n126 ) , .B1( u2_u3_u6_n171 ) );
  AOI22_X1 u2_u3_u6_U78 (.ZN( u2_u3_u6_n104 ) , .A1( u2_u3_u6_n111 ) , .B1( u2_u3_u6_n124 ) , .B2( u2_u3_u6_n151 ) , .A2( u2_u3_u6_n93 ) );
  NAND4_X1 u2_u3_u6_U79 (.ZN( u2_out3_12 ) , .A4( u2_u3_u6_n114 ) , .A3( u2_u3_u6_n115 ) , .A2( u2_u3_u6_n116 ) , .A1( u2_u3_u6_n117 ) );
  AOI21_X1 u2_u3_u6_U8 (.B1( u2_u3_u6_n107 ) , .B2( u2_u3_u6_n132 ) , .A( u2_u3_u6_n158 ) , .ZN( u2_u3_u6_n88 ) );
  OAI22_X1 u2_u3_u6_U80 (.B2( u2_u3_u6_n111 ) , .ZN( u2_u3_u6_n116 ) , .B1( u2_u3_u6_n126 ) , .A2( u2_u3_u6_n164 ) , .A1( u2_u3_u6_n167 ) );
  OAI21_X1 u2_u3_u6_U81 (.A( u2_u3_u6_n108 ) , .ZN( u2_u3_u6_n117 ) , .B2( u2_u3_u6_n141 ) , .B1( u2_u3_u6_n163 ) );
  OAI211_X1 u2_u3_u6_U82 (.ZN( u2_out3_22 ) , .B( u2_u3_u6_n137 ) , .A( u2_u3_u6_n138 ) , .C2( u2_u3_u6_n139 ) , .C1( u2_u3_u6_n140 ) );
  AOI22_X1 u2_u3_u6_U83 (.B1( u2_u3_u6_n124 ) , .A2( u2_u3_u6_n125 ) , .A1( u2_u3_u6_n126 ) , .ZN( u2_u3_u6_n138 ) , .B2( u2_u3_u6_n161 ) );
  AND4_X1 u2_u3_u6_U84 (.A3( u2_u3_u6_n119 ) , .A1( u2_u3_u6_n120 ) , .A4( u2_u3_u6_n129 ) , .ZN( u2_u3_u6_n140 ) , .A2( u2_u3_u6_n143 ) );
  OAI211_X1 u2_u3_u6_U85 (.ZN( u2_out3_7 ) , .B( u2_u3_u6_n153 ) , .C2( u2_u3_u6_n154 ) , .C1( u2_u3_u6_n155 ) , .A( u2_u3_u6_n174 ) );
  NOR3_X1 u2_u3_u6_U86 (.A1( u2_u3_u6_n141 ) , .ZN( u2_u3_u6_n154 ) , .A3( u2_u3_u6_n164 ) , .A2( u2_u3_u6_n171 ) );
  AOI211_X1 u2_u3_u6_U87 (.B( u2_u3_u6_n149 ) , .A( u2_u3_u6_n150 ) , .C2( u2_u3_u6_n151 ) , .C1( u2_u3_u6_n152 ) , .ZN( u2_u3_u6_n153 ) );
  NAND3_X1 u2_u3_u6_U88 (.A2( u2_u3_u6_n123 ) , .ZN( u2_u3_u6_n125 ) , .A1( u2_u3_u6_n130 ) , .A3( u2_u3_u6_n131 ) );
  NAND3_X1 u2_u3_u6_U89 (.A3( u2_u3_u6_n133 ) , .ZN( u2_u3_u6_n141 ) , .A1( u2_u3_u6_n145 ) , .A2( u2_u3_u6_n148 ) );
  AOI21_X1 u2_u3_u6_U9 (.B2( u2_u3_u6_n147 ) , .B1( u2_u3_u6_n148 ) , .ZN( u2_u3_u6_n149 ) , .A( u2_u3_u6_n158 ) );
  NAND3_X1 u2_u3_u6_U90 (.ZN( u2_u3_u6_n101 ) , .A3( u2_u3_u6_n107 ) , .A2( u2_u3_u6_n121 ) , .A1( u2_u3_u6_n127 ) );
  NAND3_X1 u2_u3_u6_U91 (.ZN( u2_u3_u6_n102 ) , .A3( u2_u3_u6_n130 ) , .A2( u2_u3_u6_n145 ) , .A1( u2_u3_u6_n166 ) );
  NAND3_X1 u2_u3_u6_U92 (.A3( u2_u3_u6_n113 ) , .A1( u2_u3_u6_n119 ) , .A2( u2_u3_u6_n123 ) , .ZN( u2_u3_u6_n93 ) );
  NAND3_X1 u2_u3_u6_U93 (.ZN( u2_u3_u6_n142 ) , .A2( u2_u3_u6_n172 ) , .A3( u2_u3_u6_n89 ) , .A1( u2_u3_u6_n90 ) );
  XOR2_X1 u2_u5_U1 (.B( u2_K6_9 ) , .A( u2_R4_6 ) , .Z( u2_u5_X_9 ) );
  XOR2_X1 u2_u5_U10 (.B( u2_K6_45 ) , .A( u2_R4_30 ) , .Z( u2_u5_X_45 ) );
  XOR2_X1 u2_u5_U11 (.B( u2_K6_44 ) , .A( u2_R4_29 ) , .Z( u2_u5_X_44 ) );
  XOR2_X1 u2_u5_U12 (.B( u2_K6_43 ) , .A( u2_R4_28 ) , .Z( u2_u5_X_43 ) );
  XOR2_X1 u2_u5_U16 (.B( u2_K6_3 ) , .A( u2_R4_2 ) , .Z( u2_u5_X_3 ) );
  XOR2_X1 u2_u5_U2 (.B( u2_K6_8 ) , .A( u2_R4_5 ) , .Z( u2_u5_X_8 ) );
  XOR2_X1 u2_u5_U27 (.B( u2_K6_2 ) , .A( u2_R4_1 ) , .Z( u2_u5_X_2 ) );
  XOR2_X1 u2_u5_U3 (.B( u2_K6_7 ) , .A( u2_R4_4 ) , .Z( u2_u5_X_7 ) );
  XOR2_X1 u2_u5_U38 (.B( u2_K6_1 ) , .A( u2_R4_32 ) , .Z( u2_u5_X_1 ) );
  XOR2_X1 u2_u5_U4 (.B( u2_K6_6 ) , .A( u2_R4_5 ) , .Z( u2_u5_X_6 ) );
  XOR2_X1 u2_u5_U46 (.B( u2_K6_12 ) , .A( u2_R4_9 ) , .Z( u2_u5_X_12 ) );
  XOR2_X1 u2_u5_U47 (.B( u2_K6_11 ) , .A( u2_R4_8 ) , .Z( u2_u5_X_11 ) );
  XOR2_X1 u2_u5_U48 (.B( u2_K6_10 ) , .A( u2_R4_7 ) , .Z( u2_u5_X_10 ) );
  XOR2_X1 u2_u5_U5 (.B( u2_K6_5 ) , .A( u2_R4_4 ) , .Z( u2_u5_X_5 ) );
  XOR2_X1 u2_u5_U6 (.B( u2_K6_4 ) , .A( u2_R4_3 ) , .Z( u2_u5_X_4 ) );
  XOR2_X1 u2_u5_U7 (.B( u2_K6_48 ) , .A( u2_R4_1 ) , .Z( u2_u5_X_48 ) );
  XOR2_X1 u2_u5_U8 (.B( u2_K6_47 ) , .A( u2_R4_32 ) , .Z( u2_u5_X_47 ) );
  XOR2_X1 u2_u5_U9 (.B( u2_K6_46 ) , .A( u2_R4_31 ) , .Z( u2_u5_X_46 ) );
  AND3_X1 u2_u5_u0_U10 (.A2( u2_u5_u0_n112 ) , .ZN( u2_u5_u0_n127 ) , .A3( u2_u5_u0_n130 ) , .A1( u2_u5_u0_n148 ) );
  NAND2_X1 u2_u5_u0_U11 (.ZN( u2_u5_u0_n113 ) , .A1( u2_u5_u0_n139 ) , .A2( u2_u5_u0_n149 ) );
  AND2_X1 u2_u5_u0_U12 (.ZN( u2_u5_u0_n107 ) , .A1( u2_u5_u0_n130 ) , .A2( u2_u5_u0_n140 ) );
  AND2_X1 u2_u5_u0_U13 (.A2( u2_u5_u0_n129 ) , .A1( u2_u5_u0_n130 ) , .ZN( u2_u5_u0_n151 ) );
  AND2_X1 u2_u5_u0_U14 (.A1( u2_u5_u0_n108 ) , .A2( u2_u5_u0_n125 ) , .ZN( u2_u5_u0_n145 ) );
  INV_X1 u2_u5_u0_U15 (.A( u2_u5_u0_n143 ) , .ZN( u2_u5_u0_n173 ) );
  NOR2_X1 u2_u5_u0_U16 (.A2( u2_u5_u0_n136 ) , .ZN( u2_u5_u0_n147 ) , .A1( u2_u5_u0_n160 ) );
  AOI21_X1 u2_u5_u0_U17 (.B1( u2_u5_u0_n103 ) , .ZN( u2_u5_u0_n132 ) , .A( u2_u5_u0_n165 ) , .B2( u2_u5_u0_n93 ) );
  INV_X1 u2_u5_u0_U18 (.A( u2_u5_u0_n142 ) , .ZN( u2_u5_u0_n165 ) );
  OAI22_X1 u2_u5_u0_U19 (.B1( u2_u5_u0_n125 ) , .ZN( u2_u5_u0_n126 ) , .A1( u2_u5_u0_n138 ) , .A2( u2_u5_u0_n146 ) , .B2( u2_u5_u0_n147 ) );
  OAI22_X1 u2_u5_u0_U20 (.B1( u2_u5_u0_n131 ) , .A1( u2_u5_u0_n144 ) , .B2( u2_u5_u0_n147 ) , .A2( u2_u5_u0_n90 ) , .ZN( u2_u5_u0_n91 ) );
  AND3_X1 u2_u5_u0_U21 (.A3( u2_u5_u0_n121 ) , .A2( u2_u5_u0_n125 ) , .A1( u2_u5_u0_n148 ) , .ZN( u2_u5_u0_n90 ) );
  INV_X1 u2_u5_u0_U22 (.A( u2_u5_u0_n136 ) , .ZN( u2_u5_u0_n161 ) );
  AOI22_X1 u2_u5_u0_U23 (.B2( u2_u5_u0_n109 ) , .A2( u2_u5_u0_n110 ) , .ZN( u2_u5_u0_n111 ) , .B1( u2_u5_u0_n118 ) , .A1( u2_u5_u0_n160 ) );
  INV_X1 u2_u5_u0_U24 (.A( u2_u5_u0_n118 ) , .ZN( u2_u5_u0_n158 ) );
  AOI21_X1 u2_u5_u0_U25 (.ZN( u2_u5_u0_n104 ) , .B1( u2_u5_u0_n107 ) , .B2( u2_u5_u0_n141 ) , .A( u2_u5_u0_n144 ) );
  AOI21_X1 u2_u5_u0_U26 (.B1( u2_u5_u0_n127 ) , .B2( u2_u5_u0_n129 ) , .A( u2_u5_u0_n138 ) , .ZN( u2_u5_u0_n96 ) );
  AOI21_X1 u2_u5_u0_U27 (.ZN( u2_u5_u0_n116 ) , .B2( u2_u5_u0_n142 ) , .A( u2_u5_u0_n144 ) , .B1( u2_u5_u0_n166 ) );
  NOR2_X1 u2_u5_u0_U28 (.A1( u2_u5_u0_n120 ) , .ZN( u2_u5_u0_n143 ) , .A2( u2_u5_u0_n167 ) );
  OAI221_X1 u2_u5_u0_U29 (.C1( u2_u5_u0_n112 ) , .ZN( u2_u5_u0_n120 ) , .B1( u2_u5_u0_n138 ) , .B2( u2_u5_u0_n141 ) , .C2( u2_u5_u0_n147 ) , .A( u2_u5_u0_n172 ) );
  INV_X1 u2_u5_u0_U3 (.A( u2_u5_u0_n113 ) , .ZN( u2_u5_u0_n166 ) );
  AOI211_X1 u2_u5_u0_U30 (.B( u2_u5_u0_n115 ) , .A( u2_u5_u0_n116 ) , .C2( u2_u5_u0_n117 ) , .C1( u2_u5_u0_n118 ) , .ZN( u2_u5_u0_n119 ) );
  NAND2_X1 u2_u5_u0_U31 (.A1( u2_u5_u0_n100 ) , .A2( u2_u5_u0_n103 ) , .ZN( u2_u5_u0_n125 ) );
  NAND2_X1 u2_u5_u0_U32 (.A2( u2_u5_u0_n103 ) , .ZN( u2_u5_u0_n140 ) , .A1( u2_u5_u0_n94 ) );
  NAND2_X1 u2_u5_u0_U33 (.A1( u2_u5_u0_n101 ) , .A2( u2_u5_u0_n102 ) , .ZN( u2_u5_u0_n150 ) );
  INV_X1 u2_u5_u0_U34 (.A( u2_u5_u0_n138 ) , .ZN( u2_u5_u0_n160 ) );
  NAND2_X1 u2_u5_u0_U35 (.A2( u2_u5_u0_n102 ) , .A1( u2_u5_u0_n103 ) , .ZN( u2_u5_u0_n149 ) );
  NAND2_X1 u2_u5_u0_U36 (.A2( u2_u5_u0_n100 ) , .A1( u2_u5_u0_n101 ) , .ZN( u2_u5_u0_n139 ) );
  NAND2_X1 u2_u5_u0_U37 (.A2( u2_u5_u0_n100 ) , .ZN( u2_u5_u0_n131 ) , .A1( u2_u5_u0_n92 ) );
  NAND2_X1 u2_u5_u0_U38 (.ZN( u2_u5_u0_n108 ) , .A1( u2_u5_u0_n92 ) , .A2( u2_u5_u0_n94 ) );
  NAND2_X1 u2_u5_u0_U39 (.A2( u2_u5_u0_n102 ) , .ZN( u2_u5_u0_n114 ) , .A1( u2_u5_u0_n92 ) );
  AOI21_X1 u2_u5_u0_U4 (.B1( u2_u5_u0_n114 ) , .ZN( u2_u5_u0_n115 ) , .B2( u2_u5_u0_n129 ) , .A( u2_u5_u0_n161 ) );
  NAND2_X1 u2_u5_u0_U40 (.A1( u2_u5_u0_n101 ) , .ZN( u2_u5_u0_n130 ) , .A2( u2_u5_u0_n94 ) );
  NAND2_X1 u2_u5_u0_U41 (.A2( u2_u5_u0_n101 ) , .ZN( u2_u5_u0_n121 ) , .A1( u2_u5_u0_n93 ) );
  INV_X1 u2_u5_u0_U42 (.ZN( u2_u5_u0_n172 ) , .A( u2_u5_u0_n88 ) );
  OAI222_X1 u2_u5_u0_U43 (.C1( u2_u5_u0_n108 ) , .A1( u2_u5_u0_n125 ) , .B2( u2_u5_u0_n128 ) , .B1( u2_u5_u0_n144 ) , .A2( u2_u5_u0_n158 ) , .C2( u2_u5_u0_n161 ) , .ZN( u2_u5_u0_n88 ) );
  NAND2_X1 u2_u5_u0_U44 (.ZN( u2_u5_u0_n112 ) , .A2( u2_u5_u0_n92 ) , .A1( u2_u5_u0_n93 ) );
  OR3_X1 u2_u5_u0_U45 (.A3( u2_u5_u0_n152 ) , .A2( u2_u5_u0_n153 ) , .A1( u2_u5_u0_n154 ) , .ZN( u2_u5_u0_n155 ) );
  AOI21_X1 u2_u5_u0_U46 (.A( u2_u5_u0_n144 ) , .B2( u2_u5_u0_n145 ) , .B1( u2_u5_u0_n146 ) , .ZN( u2_u5_u0_n154 ) );
  AOI21_X1 u2_u5_u0_U47 (.B2( u2_u5_u0_n150 ) , .B1( u2_u5_u0_n151 ) , .ZN( u2_u5_u0_n152 ) , .A( u2_u5_u0_n158 ) );
  AOI21_X1 u2_u5_u0_U48 (.A( u2_u5_u0_n147 ) , .B2( u2_u5_u0_n148 ) , .B1( u2_u5_u0_n149 ) , .ZN( u2_u5_u0_n153 ) );
  INV_X1 u2_u5_u0_U49 (.ZN( u2_u5_u0_n171 ) , .A( u2_u5_u0_n99 ) );
  AOI21_X1 u2_u5_u0_U5 (.B2( u2_u5_u0_n131 ) , .ZN( u2_u5_u0_n134 ) , .B1( u2_u5_u0_n151 ) , .A( u2_u5_u0_n158 ) );
  OAI211_X1 u2_u5_u0_U50 (.C2( u2_u5_u0_n140 ) , .C1( u2_u5_u0_n161 ) , .A( u2_u5_u0_n169 ) , .B( u2_u5_u0_n98 ) , .ZN( u2_u5_u0_n99 ) );
  AOI211_X1 u2_u5_u0_U51 (.C1( u2_u5_u0_n118 ) , .A( u2_u5_u0_n123 ) , .B( u2_u5_u0_n96 ) , .C2( u2_u5_u0_n97 ) , .ZN( u2_u5_u0_n98 ) );
  INV_X1 u2_u5_u0_U52 (.ZN( u2_u5_u0_n169 ) , .A( u2_u5_u0_n91 ) );
  NOR2_X1 u2_u5_u0_U53 (.A2( u2_u5_X_2 ) , .ZN( u2_u5_u0_n103 ) , .A1( u2_u5_u0_n164 ) );
  NOR2_X1 u2_u5_u0_U54 (.A2( u2_u5_X_4 ) , .A1( u2_u5_X_5 ) , .ZN( u2_u5_u0_n118 ) );
  NOR2_X1 u2_u5_u0_U55 (.A2( u2_u5_X_1 ) , .A1( u2_u5_X_2 ) , .ZN( u2_u5_u0_n92 ) );
  NOR2_X1 u2_u5_u0_U56 (.A2( u2_u5_X_1 ) , .ZN( u2_u5_u0_n101 ) , .A1( u2_u5_u0_n163 ) );
  NOR2_X1 u2_u5_u0_U57 (.A2( u2_u5_X_3 ) , .A1( u2_u5_X_6 ) , .ZN( u2_u5_u0_n94 ) );
  NOR2_X1 u2_u5_u0_U58 (.A2( u2_u5_X_6 ) , .ZN( u2_u5_u0_n100 ) , .A1( u2_u5_u0_n162 ) );
  NAND2_X1 u2_u5_u0_U59 (.A2( u2_u5_X_4 ) , .A1( u2_u5_X_5 ) , .ZN( u2_u5_u0_n144 ) );
  NOR2_X1 u2_u5_u0_U6 (.A1( u2_u5_u0_n108 ) , .ZN( u2_u5_u0_n123 ) , .A2( u2_u5_u0_n158 ) );
  NOR2_X1 u2_u5_u0_U60 (.A2( u2_u5_X_5 ) , .ZN( u2_u5_u0_n136 ) , .A1( u2_u5_u0_n159 ) );
  NAND2_X1 u2_u5_u0_U61 (.A1( u2_u5_X_5 ) , .ZN( u2_u5_u0_n138 ) , .A2( u2_u5_u0_n159 ) );
  AND2_X1 u2_u5_u0_U62 (.A2( u2_u5_X_3 ) , .A1( u2_u5_X_6 ) , .ZN( u2_u5_u0_n102 ) );
  AND2_X1 u2_u5_u0_U63 (.A1( u2_u5_X_6 ) , .A2( u2_u5_u0_n162 ) , .ZN( u2_u5_u0_n93 ) );
  INV_X1 u2_u5_u0_U64 (.A( u2_u5_X_4 ) , .ZN( u2_u5_u0_n159 ) );
  INV_X1 u2_u5_u0_U65 (.A( u2_u5_X_1 ) , .ZN( u2_u5_u0_n164 ) );
  INV_X1 u2_u5_u0_U66 (.A( u2_u5_X_2 ) , .ZN( u2_u5_u0_n163 ) );
  INV_X1 u2_u5_u0_U67 (.A( u2_u5_X_3 ) , .ZN( u2_u5_u0_n162 ) );
  INV_X1 u2_u5_u0_U68 (.A( u2_u5_u0_n126 ) , .ZN( u2_u5_u0_n168 ) );
  AOI211_X1 u2_u5_u0_U69 (.B( u2_u5_u0_n133 ) , .A( u2_u5_u0_n134 ) , .C2( u2_u5_u0_n135 ) , .C1( u2_u5_u0_n136 ) , .ZN( u2_u5_u0_n137 ) );
  OAI21_X1 u2_u5_u0_U7 (.B1( u2_u5_u0_n150 ) , .B2( u2_u5_u0_n158 ) , .A( u2_u5_u0_n172 ) , .ZN( u2_u5_u0_n89 ) );
  OR4_X1 u2_u5_u0_U70 (.ZN( u2_out5_17 ) , .A4( u2_u5_u0_n122 ) , .A2( u2_u5_u0_n123 ) , .A1( u2_u5_u0_n124 ) , .A3( u2_u5_u0_n170 ) );
  AOI21_X1 u2_u5_u0_U71 (.B2( u2_u5_u0_n107 ) , .ZN( u2_u5_u0_n124 ) , .B1( u2_u5_u0_n128 ) , .A( u2_u5_u0_n161 ) );
  INV_X1 u2_u5_u0_U72 (.A( u2_u5_u0_n111 ) , .ZN( u2_u5_u0_n170 ) );
  OR4_X1 u2_u5_u0_U73 (.ZN( u2_out5_31 ) , .A4( u2_u5_u0_n155 ) , .A2( u2_u5_u0_n156 ) , .A1( u2_u5_u0_n157 ) , .A3( u2_u5_u0_n173 ) );
  AOI21_X1 u2_u5_u0_U74 (.A( u2_u5_u0_n138 ) , .B2( u2_u5_u0_n139 ) , .B1( u2_u5_u0_n140 ) , .ZN( u2_u5_u0_n157 ) );
  AOI21_X1 u2_u5_u0_U75 (.B2( u2_u5_u0_n141 ) , .B1( u2_u5_u0_n142 ) , .ZN( u2_u5_u0_n156 ) , .A( u2_u5_u0_n161 ) );
  INV_X1 u2_u5_u0_U76 (.ZN( u2_u5_u0_n174 ) , .A( u2_u5_u0_n89 ) );
  AOI211_X1 u2_u5_u0_U77 (.B( u2_u5_u0_n104 ) , .A( u2_u5_u0_n105 ) , .ZN( u2_u5_u0_n106 ) , .C2( u2_u5_u0_n113 ) , .C1( u2_u5_u0_n160 ) );
  NOR2_X1 u2_u5_u0_U78 (.A1( u2_u5_u0_n163 ) , .A2( u2_u5_u0_n164 ) , .ZN( u2_u5_u0_n95 ) );
  OAI221_X1 u2_u5_u0_U79 (.C1( u2_u5_u0_n121 ) , .ZN( u2_u5_u0_n122 ) , .B2( u2_u5_u0_n127 ) , .A( u2_u5_u0_n143 ) , .B1( u2_u5_u0_n144 ) , .C2( u2_u5_u0_n147 ) );
  AND2_X1 u2_u5_u0_U8 (.A1( u2_u5_u0_n114 ) , .A2( u2_u5_u0_n121 ) , .ZN( u2_u5_u0_n146 ) );
  AOI21_X1 u2_u5_u0_U80 (.B1( u2_u5_u0_n132 ) , .ZN( u2_u5_u0_n133 ) , .A( u2_u5_u0_n144 ) , .B2( u2_u5_u0_n166 ) );
  OAI22_X1 u2_u5_u0_U81 (.ZN( u2_u5_u0_n105 ) , .A2( u2_u5_u0_n132 ) , .B1( u2_u5_u0_n146 ) , .A1( u2_u5_u0_n147 ) , .B2( u2_u5_u0_n161 ) );
  NAND2_X1 u2_u5_u0_U82 (.ZN( u2_u5_u0_n110 ) , .A2( u2_u5_u0_n132 ) , .A1( u2_u5_u0_n145 ) );
  INV_X1 u2_u5_u0_U83 (.A( u2_u5_u0_n119 ) , .ZN( u2_u5_u0_n167 ) );
  NAND2_X1 u2_u5_u0_U84 (.ZN( u2_u5_u0_n148 ) , .A1( u2_u5_u0_n93 ) , .A2( u2_u5_u0_n95 ) );
  NAND2_X1 u2_u5_u0_U85 (.A1( u2_u5_u0_n100 ) , .ZN( u2_u5_u0_n129 ) , .A2( u2_u5_u0_n95 ) );
  NAND2_X1 u2_u5_u0_U86 (.A1( u2_u5_u0_n102 ) , .ZN( u2_u5_u0_n128 ) , .A2( u2_u5_u0_n95 ) );
  NAND2_X1 u2_u5_u0_U87 (.ZN( u2_u5_u0_n142 ) , .A1( u2_u5_u0_n94 ) , .A2( u2_u5_u0_n95 ) );
  NAND3_X1 u2_u5_u0_U88 (.ZN( u2_out5_23 ) , .A3( u2_u5_u0_n137 ) , .A1( u2_u5_u0_n168 ) , .A2( u2_u5_u0_n171 ) );
  NAND3_X1 u2_u5_u0_U89 (.A3( u2_u5_u0_n127 ) , .A2( u2_u5_u0_n128 ) , .ZN( u2_u5_u0_n135 ) , .A1( u2_u5_u0_n150 ) );
  AND2_X1 u2_u5_u0_U9 (.A1( u2_u5_u0_n131 ) , .ZN( u2_u5_u0_n141 ) , .A2( u2_u5_u0_n150 ) );
  NAND3_X1 u2_u5_u0_U90 (.ZN( u2_u5_u0_n117 ) , .A3( u2_u5_u0_n132 ) , .A2( u2_u5_u0_n139 ) , .A1( u2_u5_u0_n148 ) );
  NAND3_X1 u2_u5_u0_U91 (.ZN( u2_u5_u0_n109 ) , .A2( u2_u5_u0_n114 ) , .A3( u2_u5_u0_n140 ) , .A1( u2_u5_u0_n149 ) );
  NAND3_X1 u2_u5_u0_U92 (.ZN( u2_out5_9 ) , .A3( u2_u5_u0_n106 ) , .A2( u2_u5_u0_n171 ) , .A1( u2_u5_u0_n174 ) );
  NAND3_X1 u2_u5_u0_U93 (.A2( u2_u5_u0_n128 ) , .A1( u2_u5_u0_n132 ) , .A3( u2_u5_u0_n146 ) , .ZN( u2_u5_u0_n97 ) );
  NOR2_X1 u2_u5_u1_U10 (.A1( u2_u5_u1_n112 ) , .A2( u2_u5_u1_n116 ) , .ZN( u2_u5_u1_n118 ) );
  NAND3_X1 u2_u5_u1_U100 (.ZN( u2_u5_u1_n113 ) , .A1( u2_u5_u1_n120 ) , .A3( u2_u5_u1_n133 ) , .A2( u2_u5_u1_n155 ) );
  OAI21_X1 u2_u5_u1_U11 (.ZN( u2_u5_u1_n101 ) , .B1( u2_u5_u1_n141 ) , .A( u2_u5_u1_n146 ) , .B2( u2_u5_u1_n183 ) );
  AOI21_X1 u2_u5_u1_U12 (.B2( u2_u5_u1_n155 ) , .B1( u2_u5_u1_n156 ) , .ZN( u2_u5_u1_n157 ) , .A( u2_u5_u1_n174 ) );
  NAND2_X1 u2_u5_u1_U13 (.ZN( u2_u5_u1_n140 ) , .A2( u2_u5_u1_n150 ) , .A1( u2_u5_u1_n155 ) );
  NAND2_X1 u2_u5_u1_U14 (.A1( u2_u5_u1_n131 ) , .ZN( u2_u5_u1_n147 ) , .A2( u2_u5_u1_n153 ) );
  INV_X1 u2_u5_u1_U15 (.A( u2_u5_u1_n139 ) , .ZN( u2_u5_u1_n174 ) );
  OR4_X1 u2_u5_u1_U16 (.A4( u2_u5_u1_n106 ) , .A3( u2_u5_u1_n107 ) , .ZN( u2_u5_u1_n108 ) , .A1( u2_u5_u1_n117 ) , .A2( u2_u5_u1_n184 ) );
  AOI21_X1 u2_u5_u1_U17 (.ZN( u2_u5_u1_n106 ) , .A( u2_u5_u1_n112 ) , .B1( u2_u5_u1_n154 ) , .B2( u2_u5_u1_n156 ) );
  INV_X1 u2_u5_u1_U18 (.A( u2_u5_u1_n101 ) , .ZN( u2_u5_u1_n184 ) );
  AOI21_X1 u2_u5_u1_U19 (.ZN( u2_u5_u1_n107 ) , .B1( u2_u5_u1_n134 ) , .B2( u2_u5_u1_n149 ) , .A( u2_u5_u1_n174 ) );
  INV_X1 u2_u5_u1_U20 (.A( u2_u5_u1_n112 ) , .ZN( u2_u5_u1_n171 ) );
  NAND2_X1 u2_u5_u1_U21 (.ZN( u2_u5_u1_n141 ) , .A1( u2_u5_u1_n153 ) , .A2( u2_u5_u1_n156 ) );
  AND2_X1 u2_u5_u1_U22 (.A1( u2_u5_u1_n123 ) , .ZN( u2_u5_u1_n134 ) , .A2( u2_u5_u1_n161 ) );
  NAND2_X1 u2_u5_u1_U23 (.A2( u2_u5_u1_n115 ) , .A1( u2_u5_u1_n116 ) , .ZN( u2_u5_u1_n148 ) );
  NAND2_X1 u2_u5_u1_U24 (.A2( u2_u5_u1_n133 ) , .A1( u2_u5_u1_n135 ) , .ZN( u2_u5_u1_n159 ) );
  NAND2_X1 u2_u5_u1_U25 (.A2( u2_u5_u1_n115 ) , .A1( u2_u5_u1_n120 ) , .ZN( u2_u5_u1_n132 ) );
  INV_X1 u2_u5_u1_U26 (.A( u2_u5_u1_n154 ) , .ZN( u2_u5_u1_n178 ) );
  INV_X1 u2_u5_u1_U27 (.A( u2_u5_u1_n151 ) , .ZN( u2_u5_u1_n183 ) );
  AND2_X1 u2_u5_u1_U28 (.A1( u2_u5_u1_n129 ) , .A2( u2_u5_u1_n133 ) , .ZN( u2_u5_u1_n149 ) );
  INV_X1 u2_u5_u1_U29 (.A( u2_u5_u1_n131 ) , .ZN( u2_u5_u1_n180 ) );
  INV_X1 u2_u5_u1_U3 (.A( u2_u5_u1_n159 ) , .ZN( u2_u5_u1_n182 ) );
  OAI221_X1 u2_u5_u1_U30 (.A( u2_u5_u1_n119 ) , .C2( u2_u5_u1_n129 ) , .ZN( u2_u5_u1_n138 ) , .B2( u2_u5_u1_n152 ) , .C1( u2_u5_u1_n174 ) , .B1( u2_u5_u1_n187 ) );
  INV_X1 u2_u5_u1_U31 (.A( u2_u5_u1_n148 ) , .ZN( u2_u5_u1_n187 ) );
  AOI211_X1 u2_u5_u1_U32 (.B( u2_u5_u1_n117 ) , .A( u2_u5_u1_n118 ) , .ZN( u2_u5_u1_n119 ) , .C2( u2_u5_u1_n146 ) , .C1( u2_u5_u1_n159 ) );
  NOR2_X1 u2_u5_u1_U33 (.A1( u2_u5_u1_n168 ) , .A2( u2_u5_u1_n176 ) , .ZN( u2_u5_u1_n98 ) );
  OAI21_X1 u2_u5_u1_U34 (.B2( u2_u5_u1_n123 ) , .ZN( u2_u5_u1_n145 ) , .B1( u2_u5_u1_n160 ) , .A( u2_u5_u1_n185 ) );
  INV_X1 u2_u5_u1_U35 (.A( u2_u5_u1_n122 ) , .ZN( u2_u5_u1_n185 ) );
  AOI21_X1 u2_u5_u1_U36 (.B2( u2_u5_u1_n120 ) , .B1( u2_u5_u1_n121 ) , .ZN( u2_u5_u1_n122 ) , .A( u2_u5_u1_n128 ) );
  NAND2_X1 u2_u5_u1_U37 (.A1( u2_u5_u1_n128 ) , .ZN( u2_u5_u1_n146 ) , .A2( u2_u5_u1_n160 ) );
  NAND2_X1 u2_u5_u1_U38 (.A2( u2_u5_u1_n112 ) , .ZN( u2_u5_u1_n139 ) , .A1( u2_u5_u1_n152 ) );
  NAND2_X1 u2_u5_u1_U39 (.A1( u2_u5_u1_n105 ) , .ZN( u2_u5_u1_n156 ) , .A2( u2_u5_u1_n99 ) );
  AOI221_X1 u2_u5_u1_U4 (.A( u2_u5_u1_n138 ) , .C2( u2_u5_u1_n139 ) , .C1( u2_u5_u1_n140 ) , .B2( u2_u5_u1_n141 ) , .ZN( u2_u5_u1_n142 ) , .B1( u2_u5_u1_n175 ) );
  AOI221_X1 u2_u5_u1_U40 (.B1( u2_u5_u1_n140 ) , .ZN( u2_u5_u1_n167 ) , .B2( u2_u5_u1_n172 ) , .C2( u2_u5_u1_n175 ) , .C1( u2_u5_u1_n178 ) , .A( u2_u5_u1_n188 ) );
  INV_X1 u2_u5_u1_U41 (.ZN( u2_u5_u1_n188 ) , .A( u2_u5_u1_n97 ) );
  AOI211_X1 u2_u5_u1_U42 (.A( u2_u5_u1_n118 ) , .C1( u2_u5_u1_n132 ) , .C2( u2_u5_u1_n139 ) , .B( u2_u5_u1_n96 ) , .ZN( u2_u5_u1_n97 ) );
  AOI21_X1 u2_u5_u1_U43 (.B2( u2_u5_u1_n121 ) , .B1( u2_u5_u1_n135 ) , .A( u2_u5_u1_n152 ) , .ZN( u2_u5_u1_n96 ) );
  NOR2_X1 u2_u5_u1_U44 (.ZN( u2_u5_u1_n117 ) , .A1( u2_u5_u1_n121 ) , .A2( u2_u5_u1_n160 ) );
  AOI21_X1 u2_u5_u1_U45 (.A( u2_u5_u1_n128 ) , .B2( u2_u5_u1_n129 ) , .ZN( u2_u5_u1_n130 ) , .B1( u2_u5_u1_n150 ) );
  NAND2_X1 u2_u5_u1_U46 (.ZN( u2_u5_u1_n112 ) , .A1( u2_u5_u1_n169 ) , .A2( u2_u5_u1_n170 ) );
  NAND2_X1 u2_u5_u1_U47 (.ZN( u2_u5_u1_n129 ) , .A2( u2_u5_u1_n95 ) , .A1( u2_u5_u1_n98 ) );
  NAND2_X1 u2_u5_u1_U48 (.A1( u2_u5_u1_n102 ) , .ZN( u2_u5_u1_n154 ) , .A2( u2_u5_u1_n99 ) );
  NAND2_X1 u2_u5_u1_U49 (.A2( u2_u5_u1_n100 ) , .ZN( u2_u5_u1_n135 ) , .A1( u2_u5_u1_n99 ) );
  AOI211_X1 u2_u5_u1_U5 (.ZN( u2_u5_u1_n124 ) , .A( u2_u5_u1_n138 ) , .C2( u2_u5_u1_n139 ) , .B( u2_u5_u1_n145 ) , .C1( u2_u5_u1_n147 ) );
  AOI21_X1 u2_u5_u1_U50 (.A( u2_u5_u1_n152 ) , .B2( u2_u5_u1_n153 ) , .B1( u2_u5_u1_n154 ) , .ZN( u2_u5_u1_n158 ) );
  INV_X1 u2_u5_u1_U51 (.A( u2_u5_u1_n160 ) , .ZN( u2_u5_u1_n175 ) );
  NAND2_X1 u2_u5_u1_U52 (.A1( u2_u5_u1_n100 ) , .ZN( u2_u5_u1_n116 ) , .A2( u2_u5_u1_n95 ) );
  NAND2_X1 u2_u5_u1_U53 (.A1( u2_u5_u1_n102 ) , .ZN( u2_u5_u1_n131 ) , .A2( u2_u5_u1_n95 ) );
  NAND2_X1 u2_u5_u1_U54 (.A2( u2_u5_u1_n104 ) , .ZN( u2_u5_u1_n121 ) , .A1( u2_u5_u1_n98 ) );
  NAND2_X1 u2_u5_u1_U55 (.A1( u2_u5_u1_n103 ) , .ZN( u2_u5_u1_n153 ) , .A2( u2_u5_u1_n98 ) );
  NAND2_X1 u2_u5_u1_U56 (.A2( u2_u5_u1_n104 ) , .A1( u2_u5_u1_n105 ) , .ZN( u2_u5_u1_n133 ) );
  NAND2_X1 u2_u5_u1_U57 (.ZN( u2_u5_u1_n150 ) , .A2( u2_u5_u1_n98 ) , .A1( u2_u5_u1_n99 ) );
  NAND2_X1 u2_u5_u1_U58 (.A1( u2_u5_u1_n105 ) , .ZN( u2_u5_u1_n155 ) , .A2( u2_u5_u1_n95 ) );
  OAI21_X1 u2_u5_u1_U59 (.ZN( u2_u5_u1_n109 ) , .B1( u2_u5_u1_n129 ) , .B2( u2_u5_u1_n160 ) , .A( u2_u5_u1_n167 ) );
  AOI22_X1 u2_u5_u1_U6 (.B2( u2_u5_u1_n136 ) , .A2( u2_u5_u1_n137 ) , .ZN( u2_u5_u1_n143 ) , .A1( u2_u5_u1_n171 ) , .B1( u2_u5_u1_n173 ) );
  NAND2_X1 u2_u5_u1_U60 (.A2( u2_u5_u1_n100 ) , .A1( u2_u5_u1_n103 ) , .ZN( u2_u5_u1_n120 ) );
  NAND2_X1 u2_u5_u1_U61 (.A1( u2_u5_u1_n102 ) , .A2( u2_u5_u1_n104 ) , .ZN( u2_u5_u1_n115 ) );
  NAND2_X1 u2_u5_u1_U62 (.A2( u2_u5_u1_n100 ) , .A1( u2_u5_u1_n104 ) , .ZN( u2_u5_u1_n151 ) );
  NAND2_X1 u2_u5_u1_U63 (.A2( u2_u5_u1_n103 ) , .A1( u2_u5_u1_n105 ) , .ZN( u2_u5_u1_n161 ) );
  INV_X1 u2_u5_u1_U64 (.A( u2_u5_u1_n152 ) , .ZN( u2_u5_u1_n173 ) );
  INV_X1 u2_u5_u1_U65 (.A( u2_u5_u1_n128 ) , .ZN( u2_u5_u1_n172 ) );
  NAND2_X1 u2_u5_u1_U66 (.A2( u2_u5_u1_n102 ) , .A1( u2_u5_u1_n103 ) , .ZN( u2_u5_u1_n123 ) );
  AOI211_X1 u2_u5_u1_U67 (.B( u2_u5_u1_n162 ) , .A( u2_u5_u1_n163 ) , .C2( u2_u5_u1_n164 ) , .ZN( u2_u5_u1_n165 ) , .C1( u2_u5_u1_n171 ) );
  AOI21_X1 u2_u5_u1_U68 (.A( u2_u5_u1_n160 ) , .B2( u2_u5_u1_n161 ) , .ZN( u2_u5_u1_n162 ) , .B1( u2_u5_u1_n182 ) );
  OR2_X1 u2_u5_u1_U69 (.A2( u2_u5_u1_n157 ) , .A1( u2_u5_u1_n158 ) , .ZN( u2_u5_u1_n163 ) );
  INV_X1 u2_u5_u1_U7 (.A( u2_u5_u1_n147 ) , .ZN( u2_u5_u1_n181 ) );
  NOR2_X1 u2_u5_u1_U70 (.A2( u2_u5_X_7 ) , .A1( u2_u5_X_8 ) , .ZN( u2_u5_u1_n95 ) );
  NOR2_X1 u2_u5_u1_U71 (.A1( u2_u5_X_12 ) , .A2( u2_u5_X_9 ) , .ZN( u2_u5_u1_n100 ) );
  NOR2_X1 u2_u5_u1_U72 (.A2( u2_u5_X_8 ) , .A1( u2_u5_u1_n177 ) , .ZN( u2_u5_u1_n99 ) );
  NOR2_X1 u2_u5_u1_U73 (.A2( u2_u5_X_12 ) , .ZN( u2_u5_u1_n102 ) , .A1( u2_u5_u1_n176 ) );
  NOR2_X1 u2_u5_u1_U74 (.A2( u2_u5_X_9 ) , .ZN( u2_u5_u1_n105 ) , .A1( u2_u5_u1_n168 ) );
  NAND2_X1 u2_u5_u1_U75 (.A1( u2_u5_X_10 ) , .ZN( u2_u5_u1_n160 ) , .A2( u2_u5_u1_n169 ) );
  NAND2_X1 u2_u5_u1_U76 (.A2( u2_u5_X_10 ) , .A1( u2_u5_X_11 ) , .ZN( u2_u5_u1_n152 ) );
  NAND2_X1 u2_u5_u1_U77 (.A1( u2_u5_X_11 ) , .ZN( u2_u5_u1_n128 ) , .A2( u2_u5_u1_n170 ) );
  AND2_X1 u2_u5_u1_U78 (.A2( u2_u5_X_7 ) , .A1( u2_u5_X_8 ) , .ZN( u2_u5_u1_n104 ) );
  AND2_X1 u2_u5_u1_U79 (.A1( u2_u5_X_8 ) , .ZN( u2_u5_u1_n103 ) , .A2( u2_u5_u1_n177 ) );
  AOI22_X1 u2_u5_u1_U8 (.B2( u2_u5_u1_n113 ) , .A2( u2_u5_u1_n114 ) , .ZN( u2_u5_u1_n125 ) , .A1( u2_u5_u1_n171 ) , .B1( u2_u5_u1_n173 ) );
  INV_X1 u2_u5_u1_U80 (.A( u2_u5_X_10 ) , .ZN( u2_u5_u1_n170 ) );
  INV_X1 u2_u5_u1_U81 (.A( u2_u5_X_9 ) , .ZN( u2_u5_u1_n176 ) );
  INV_X1 u2_u5_u1_U82 (.A( u2_u5_X_11 ) , .ZN( u2_u5_u1_n169 ) );
  INV_X1 u2_u5_u1_U83 (.A( u2_u5_X_12 ) , .ZN( u2_u5_u1_n168 ) );
  INV_X1 u2_u5_u1_U84 (.A( u2_u5_X_7 ) , .ZN( u2_u5_u1_n177 ) );
  NAND4_X1 u2_u5_u1_U85 (.ZN( u2_out5_28 ) , .A4( u2_u5_u1_n124 ) , .A3( u2_u5_u1_n125 ) , .A2( u2_u5_u1_n126 ) , .A1( u2_u5_u1_n127 ) );
  OAI21_X1 u2_u5_u1_U86 (.ZN( u2_u5_u1_n127 ) , .B2( u2_u5_u1_n139 ) , .B1( u2_u5_u1_n175 ) , .A( u2_u5_u1_n183 ) );
  OAI21_X1 u2_u5_u1_U87 (.ZN( u2_u5_u1_n126 ) , .B2( u2_u5_u1_n140 ) , .A( u2_u5_u1_n146 ) , .B1( u2_u5_u1_n178 ) );
  NAND4_X1 u2_u5_u1_U88 (.ZN( u2_out5_18 ) , .A4( u2_u5_u1_n165 ) , .A3( u2_u5_u1_n166 ) , .A1( u2_u5_u1_n167 ) , .A2( u2_u5_u1_n186 ) );
  AOI22_X1 u2_u5_u1_U89 (.B2( u2_u5_u1_n146 ) , .B1( u2_u5_u1_n147 ) , .A2( u2_u5_u1_n148 ) , .ZN( u2_u5_u1_n166 ) , .A1( u2_u5_u1_n172 ) );
  NAND2_X1 u2_u5_u1_U9 (.ZN( u2_u5_u1_n114 ) , .A1( u2_u5_u1_n134 ) , .A2( u2_u5_u1_n156 ) );
  INV_X1 u2_u5_u1_U90 (.A( u2_u5_u1_n145 ) , .ZN( u2_u5_u1_n186 ) );
  NAND4_X1 u2_u5_u1_U91 (.ZN( u2_out5_2 ) , .A4( u2_u5_u1_n142 ) , .A3( u2_u5_u1_n143 ) , .A2( u2_u5_u1_n144 ) , .A1( u2_u5_u1_n179 ) );
  OAI21_X1 u2_u5_u1_U92 (.B2( u2_u5_u1_n132 ) , .ZN( u2_u5_u1_n144 ) , .A( u2_u5_u1_n146 ) , .B1( u2_u5_u1_n180 ) );
  INV_X1 u2_u5_u1_U93 (.A( u2_u5_u1_n130 ) , .ZN( u2_u5_u1_n179 ) );
  OR4_X1 u2_u5_u1_U94 (.ZN( u2_out5_13 ) , .A4( u2_u5_u1_n108 ) , .A3( u2_u5_u1_n109 ) , .A2( u2_u5_u1_n110 ) , .A1( u2_u5_u1_n111 ) );
  AOI21_X1 u2_u5_u1_U95 (.ZN( u2_u5_u1_n110 ) , .A( u2_u5_u1_n116 ) , .B1( u2_u5_u1_n152 ) , .B2( u2_u5_u1_n160 ) );
  AOI21_X1 u2_u5_u1_U96 (.ZN( u2_u5_u1_n111 ) , .A( u2_u5_u1_n128 ) , .B2( u2_u5_u1_n131 ) , .B1( u2_u5_u1_n135 ) );
  NAND3_X1 u2_u5_u1_U97 (.A3( u2_u5_u1_n149 ) , .A2( u2_u5_u1_n150 ) , .A1( u2_u5_u1_n151 ) , .ZN( u2_u5_u1_n164 ) );
  NAND3_X1 u2_u5_u1_U98 (.A3( u2_u5_u1_n134 ) , .A2( u2_u5_u1_n135 ) , .ZN( u2_u5_u1_n136 ) , .A1( u2_u5_u1_n151 ) );
  NAND3_X1 u2_u5_u1_U99 (.A1( u2_u5_u1_n133 ) , .ZN( u2_u5_u1_n137 ) , .A2( u2_u5_u1_n154 ) , .A3( u2_u5_u1_n181 ) );
  AND3_X1 u2_u5_u7_U10 (.A3( u2_u5_u7_n110 ) , .A2( u2_u5_u7_n127 ) , .A1( u2_u5_u7_n132 ) , .ZN( u2_u5_u7_n92 ) );
  OAI21_X1 u2_u5_u7_U11 (.A( u2_u5_u7_n161 ) , .B1( u2_u5_u7_n168 ) , .B2( u2_u5_u7_n173 ) , .ZN( u2_u5_u7_n91 ) );
  AOI211_X1 u2_u5_u7_U12 (.A( u2_u5_u7_n117 ) , .ZN( u2_u5_u7_n118 ) , .C2( u2_u5_u7_n126 ) , .C1( u2_u5_u7_n177 ) , .B( u2_u5_u7_n180 ) );
  OAI22_X1 u2_u5_u7_U13 (.B1( u2_u5_u7_n115 ) , .ZN( u2_u5_u7_n117 ) , .A2( u2_u5_u7_n133 ) , .A1( u2_u5_u7_n137 ) , .B2( u2_u5_u7_n162 ) );
  INV_X1 u2_u5_u7_U14 (.A( u2_u5_u7_n116 ) , .ZN( u2_u5_u7_n180 ) );
  NOR3_X1 u2_u5_u7_U15 (.ZN( u2_u5_u7_n115 ) , .A3( u2_u5_u7_n145 ) , .A2( u2_u5_u7_n168 ) , .A1( u2_u5_u7_n169 ) );
  OAI211_X1 u2_u5_u7_U16 (.B( u2_u5_u7_n122 ) , .A( u2_u5_u7_n123 ) , .C2( u2_u5_u7_n124 ) , .ZN( u2_u5_u7_n154 ) , .C1( u2_u5_u7_n162 ) );
  AOI222_X1 u2_u5_u7_U17 (.ZN( u2_u5_u7_n122 ) , .C2( u2_u5_u7_n126 ) , .C1( u2_u5_u7_n145 ) , .B1( u2_u5_u7_n161 ) , .A2( u2_u5_u7_n165 ) , .B2( u2_u5_u7_n170 ) , .A1( u2_u5_u7_n176 ) );
  INV_X1 u2_u5_u7_U18 (.A( u2_u5_u7_n133 ) , .ZN( u2_u5_u7_n176 ) );
  NOR3_X1 u2_u5_u7_U19 (.A2( u2_u5_u7_n134 ) , .A1( u2_u5_u7_n135 ) , .ZN( u2_u5_u7_n136 ) , .A3( u2_u5_u7_n171 ) );
  NOR2_X1 u2_u5_u7_U20 (.A1( u2_u5_u7_n130 ) , .A2( u2_u5_u7_n134 ) , .ZN( u2_u5_u7_n153 ) );
  INV_X1 u2_u5_u7_U21 (.A( u2_u5_u7_n101 ) , .ZN( u2_u5_u7_n165 ) );
  NOR2_X1 u2_u5_u7_U22 (.ZN( u2_u5_u7_n111 ) , .A2( u2_u5_u7_n134 ) , .A1( u2_u5_u7_n169 ) );
  AOI21_X1 u2_u5_u7_U23 (.ZN( u2_u5_u7_n104 ) , .B2( u2_u5_u7_n112 ) , .B1( u2_u5_u7_n127 ) , .A( u2_u5_u7_n164 ) );
  AOI21_X1 u2_u5_u7_U24 (.ZN( u2_u5_u7_n106 ) , .B1( u2_u5_u7_n133 ) , .B2( u2_u5_u7_n146 ) , .A( u2_u5_u7_n162 ) );
  AOI21_X1 u2_u5_u7_U25 (.A( u2_u5_u7_n101 ) , .ZN( u2_u5_u7_n107 ) , .B2( u2_u5_u7_n128 ) , .B1( u2_u5_u7_n175 ) );
  INV_X1 u2_u5_u7_U26 (.A( u2_u5_u7_n138 ) , .ZN( u2_u5_u7_n171 ) );
  INV_X1 u2_u5_u7_U27 (.A( u2_u5_u7_n131 ) , .ZN( u2_u5_u7_n177 ) );
  INV_X1 u2_u5_u7_U28 (.A( u2_u5_u7_n110 ) , .ZN( u2_u5_u7_n174 ) );
  NAND2_X1 u2_u5_u7_U29 (.A1( u2_u5_u7_n129 ) , .A2( u2_u5_u7_n132 ) , .ZN( u2_u5_u7_n149 ) );
  OAI21_X1 u2_u5_u7_U3 (.ZN( u2_u5_u7_n159 ) , .A( u2_u5_u7_n165 ) , .B2( u2_u5_u7_n171 ) , .B1( u2_u5_u7_n174 ) );
  NAND2_X1 u2_u5_u7_U30 (.A1( u2_u5_u7_n113 ) , .A2( u2_u5_u7_n124 ) , .ZN( u2_u5_u7_n130 ) );
  INV_X1 u2_u5_u7_U31 (.A( u2_u5_u7_n112 ) , .ZN( u2_u5_u7_n173 ) );
  INV_X1 u2_u5_u7_U32 (.A( u2_u5_u7_n128 ) , .ZN( u2_u5_u7_n168 ) );
  INV_X1 u2_u5_u7_U33 (.A( u2_u5_u7_n148 ) , .ZN( u2_u5_u7_n169 ) );
  INV_X1 u2_u5_u7_U34 (.A( u2_u5_u7_n127 ) , .ZN( u2_u5_u7_n179 ) );
  NOR2_X1 u2_u5_u7_U35 (.ZN( u2_u5_u7_n101 ) , .A2( u2_u5_u7_n150 ) , .A1( u2_u5_u7_n156 ) );
  AOI211_X1 u2_u5_u7_U36 (.B( u2_u5_u7_n154 ) , .A( u2_u5_u7_n155 ) , .C1( u2_u5_u7_n156 ) , .ZN( u2_u5_u7_n157 ) , .C2( u2_u5_u7_n172 ) );
  INV_X1 u2_u5_u7_U37 (.A( u2_u5_u7_n153 ) , .ZN( u2_u5_u7_n172 ) );
  AOI211_X1 u2_u5_u7_U38 (.B( u2_u5_u7_n139 ) , .A( u2_u5_u7_n140 ) , .C2( u2_u5_u7_n141 ) , .ZN( u2_u5_u7_n142 ) , .C1( u2_u5_u7_n156 ) );
  NAND4_X1 u2_u5_u7_U39 (.A3( u2_u5_u7_n127 ) , .A2( u2_u5_u7_n128 ) , .A1( u2_u5_u7_n129 ) , .ZN( u2_u5_u7_n141 ) , .A4( u2_u5_u7_n147 ) );
  INV_X1 u2_u5_u7_U4 (.A( u2_u5_u7_n111 ) , .ZN( u2_u5_u7_n170 ) );
  AOI21_X1 u2_u5_u7_U40 (.A( u2_u5_u7_n137 ) , .B1( u2_u5_u7_n138 ) , .ZN( u2_u5_u7_n139 ) , .B2( u2_u5_u7_n146 ) );
  OAI22_X1 u2_u5_u7_U41 (.B1( u2_u5_u7_n136 ) , .ZN( u2_u5_u7_n140 ) , .A1( u2_u5_u7_n153 ) , .B2( u2_u5_u7_n162 ) , .A2( u2_u5_u7_n164 ) );
  AOI21_X1 u2_u5_u7_U42 (.ZN( u2_u5_u7_n123 ) , .B1( u2_u5_u7_n165 ) , .B2( u2_u5_u7_n177 ) , .A( u2_u5_u7_n97 ) );
  AOI21_X1 u2_u5_u7_U43 (.B2( u2_u5_u7_n113 ) , .B1( u2_u5_u7_n124 ) , .A( u2_u5_u7_n125 ) , .ZN( u2_u5_u7_n97 ) );
  INV_X1 u2_u5_u7_U44 (.A( u2_u5_u7_n125 ) , .ZN( u2_u5_u7_n161 ) );
  INV_X1 u2_u5_u7_U45 (.A( u2_u5_u7_n152 ) , .ZN( u2_u5_u7_n162 ) );
  AOI22_X1 u2_u5_u7_U46 (.A2( u2_u5_u7_n114 ) , .ZN( u2_u5_u7_n119 ) , .B1( u2_u5_u7_n130 ) , .A1( u2_u5_u7_n156 ) , .B2( u2_u5_u7_n165 ) );
  NAND2_X1 u2_u5_u7_U47 (.A2( u2_u5_u7_n112 ) , .ZN( u2_u5_u7_n114 ) , .A1( u2_u5_u7_n175 ) );
  AND2_X1 u2_u5_u7_U48 (.ZN( u2_u5_u7_n145 ) , .A2( u2_u5_u7_n98 ) , .A1( u2_u5_u7_n99 ) );
  NOR2_X1 u2_u5_u7_U49 (.ZN( u2_u5_u7_n137 ) , .A1( u2_u5_u7_n150 ) , .A2( u2_u5_u7_n161 ) );
  INV_X1 u2_u5_u7_U5 (.A( u2_u5_u7_n149 ) , .ZN( u2_u5_u7_n175 ) );
  AOI21_X1 u2_u5_u7_U50 (.ZN( u2_u5_u7_n105 ) , .B2( u2_u5_u7_n110 ) , .A( u2_u5_u7_n125 ) , .B1( u2_u5_u7_n147 ) );
  NAND2_X1 u2_u5_u7_U51 (.ZN( u2_u5_u7_n146 ) , .A1( u2_u5_u7_n95 ) , .A2( u2_u5_u7_n98 ) );
  NAND2_X1 u2_u5_u7_U52 (.A2( u2_u5_u7_n103 ) , .ZN( u2_u5_u7_n147 ) , .A1( u2_u5_u7_n93 ) );
  NAND2_X1 u2_u5_u7_U53 (.A1( u2_u5_u7_n103 ) , .ZN( u2_u5_u7_n127 ) , .A2( u2_u5_u7_n99 ) );
  OR2_X1 u2_u5_u7_U54 (.ZN( u2_u5_u7_n126 ) , .A2( u2_u5_u7_n152 ) , .A1( u2_u5_u7_n156 ) );
  NAND2_X1 u2_u5_u7_U55 (.A2( u2_u5_u7_n102 ) , .A1( u2_u5_u7_n103 ) , .ZN( u2_u5_u7_n133 ) );
  NAND2_X1 u2_u5_u7_U56 (.ZN( u2_u5_u7_n112 ) , .A2( u2_u5_u7_n96 ) , .A1( u2_u5_u7_n99 ) );
  NAND2_X1 u2_u5_u7_U57 (.A2( u2_u5_u7_n102 ) , .ZN( u2_u5_u7_n128 ) , .A1( u2_u5_u7_n98 ) );
  NAND2_X1 u2_u5_u7_U58 (.A1( u2_u5_u7_n100 ) , .ZN( u2_u5_u7_n113 ) , .A2( u2_u5_u7_n93 ) );
  NAND2_X1 u2_u5_u7_U59 (.A2( u2_u5_u7_n102 ) , .ZN( u2_u5_u7_n124 ) , .A1( u2_u5_u7_n96 ) );
  INV_X1 u2_u5_u7_U6 (.A( u2_u5_u7_n154 ) , .ZN( u2_u5_u7_n178 ) );
  NAND2_X1 u2_u5_u7_U60 (.ZN( u2_u5_u7_n110 ) , .A1( u2_u5_u7_n95 ) , .A2( u2_u5_u7_n96 ) );
  INV_X1 u2_u5_u7_U61 (.A( u2_u5_u7_n150 ) , .ZN( u2_u5_u7_n164 ) );
  AND2_X1 u2_u5_u7_U62 (.ZN( u2_u5_u7_n134 ) , .A1( u2_u5_u7_n93 ) , .A2( u2_u5_u7_n98 ) );
  NAND2_X1 u2_u5_u7_U63 (.A1( u2_u5_u7_n100 ) , .A2( u2_u5_u7_n102 ) , .ZN( u2_u5_u7_n129 ) );
  NAND2_X1 u2_u5_u7_U64 (.A2( u2_u5_u7_n103 ) , .ZN( u2_u5_u7_n131 ) , .A1( u2_u5_u7_n95 ) );
  NAND2_X1 u2_u5_u7_U65 (.A1( u2_u5_u7_n100 ) , .ZN( u2_u5_u7_n138 ) , .A2( u2_u5_u7_n99 ) );
  NAND2_X1 u2_u5_u7_U66 (.ZN( u2_u5_u7_n132 ) , .A1( u2_u5_u7_n93 ) , .A2( u2_u5_u7_n96 ) );
  NAND2_X1 u2_u5_u7_U67 (.A1( u2_u5_u7_n100 ) , .ZN( u2_u5_u7_n148 ) , .A2( u2_u5_u7_n95 ) );
  NOR2_X1 u2_u5_u7_U68 (.A2( u2_u5_X_47 ) , .ZN( u2_u5_u7_n150 ) , .A1( u2_u5_u7_n163 ) );
  NOR2_X1 u2_u5_u7_U69 (.A2( u2_u5_X_43 ) , .A1( u2_u5_X_44 ) , .ZN( u2_u5_u7_n103 ) );
  AOI211_X1 u2_u5_u7_U7 (.ZN( u2_u5_u7_n116 ) , .A( u2_u5_u7_n155 ) , .C1( u2_u5_u7_n161 ) , .C2( u2_u5_u7_n171 ) , .B( u2_u5_u7_n94 ) );
  NOR2_X1 u2_u5_u7_U70 (.A2( u2_u5_X_48 ) , .A1( u2_u5_u7_n166 ) , .ZN( u2_u5_u7_n95 ) );
  NOR2_X1 u2_u5_u7_U71 (.A2( u2_u5_X_45 ) , .A1( u2_u5_X_48 ) , .ZN( u2_u5_u7_n99 ) );
  NOR2_X1 u2_u5_u7_U72 (.A2( u2_u5_X_44 ) , .A1( u2_u5_u7_n167 ) , .ZN( u2_u5_u7_n98 ) );
  NOR2_X1 u2_u5_u7_U73 (.A2( u2_u5_X_46 ) , .A1( u2_u5_X_47 ) , .ZN( u2_u5_u7_n152 ) );
  AND2_X1 u2_u5_u7_U74 (.A1( u2_u5_X_47 ) , .ZN( u2_u5_u7_n156 ) , .A2( u2_u5_u7_n163 ) );
  NAND2_X1 u2_u5_u7_U75 (.A2( u2_u5_X_46 ) , .A1( u2_u5_X_47 ) , .ZN( u2_u5_u7_n125 ) );
  AND2_X1 u2_u5_u7_U76 (.A2( u2_u5_X_45 ) , .A1( u2_u5_X_48 ) , .ZN( u2_u5_u7_n102 ) );
  AND2_X1 u2_u5_u7_U77 (.A2( u2_u5_X_43 ) , .A1( u2_u5_X_44 ) , .ZN( u2_u5_u7_n96 ) );
  AND2_X1 u2_u5_u7_U78 (.A1( u2_u5_X_44 ) , .ZN( u2_u5_u7_n100 ) , .A2( u2_u5_u7_n167 ) );
  AND2_X1 u2_u5_u7_U79 (.A1( u2_u5_X_48 ) , .A2( u2_u5_u7_n166 ) , .ZN( u2_u5_u7_n93 ) );
  OAI222_X1 u2_u5_u7_U8 (.C2( u2_u5_u7_n101 ) , .B2( u2_u5_u7_n111 ) , .A1( u2_u5_u7_n113 ) , .C1( u2_u5_u7_n146 ) , .A2( u2_u5_u7_n162 ) , .B1( u2_u5_u7_n164 ) , .ZN( u2_u5_u7_n94 ) );
  INV_X1 u2_u5_u7_U80 (.A( u2_u5_X_46 ) , .ZN( u2_u5_u7_n163 ) );
  INV_X1 u2_u5_u7_U81 (.A( u2_u5_X_43 ) , .ZN( u2_u5_u7_n167 ) );
  INV_X1 u2_u5_u7_U82 (.A( u2_u5_X_45 ) , .ZN( u2_u5_u7_n166 ) );
  NAND4_X1 u2_u5_u7_U83 (.ZN( u2_out5_27 ) , .A4( u2_u5_u7_n118 ) , .A3( u2_u5_u7_n119 ) , .A2( u2_u5_u7_n120 ) , .A1( u2_u5_u7_n121 ) );
  OAI21_X1 u2_u5_u7_U84 (.ZN( u2_u5_u7_n121 ) , .B2( u2_u5_u7_n145 ) , .A( u2_u5_u7_n150 ) , .B1( u2_u5_u7_n174 ) );
  OAI21_X1 u2_u5_u7_U85 (.ZN( u2_u5_u7_n120 ) , .A( u2_u5_u7_n161 ) , .B2( u2_u5_u7_n170 ) , .B1( u2_u5_u7_n179 ) );
  NAND4_X1 u2_u5_u7_U86 (.ZN( u2_out5_21 ) , .A4( u2_u5_u7_n157 ) , .A3( u2_u5_u7_n158 ) , .A2( u2_u5_u7_n159 ) , .A1( u2_u5_u7_n160 ) );
  OAI21_X1 u2_u5_u7_U87 (.B1( u2_u5_u7_n145 ) , .ZN( u2_u5_u7_n160 ) , .A( u2_u5_u7_n161 ) , .B2( u2_u5_u7_n177 ) );
  AOI22_X1 u2_u5_u7_U88 (.B2( u2_u5_u7_n149 ) , .B1( u2_u5_u7_n150 ) , .A2( u2_u5_u7_n151 ) , .A1( u2_u5_u7_n152 ) , .ZN( u2_u5_u7_n158 ) );
  NAND4_X1 u2_u5_u7_U89 (.ZN( u2_out5_15 ) , .A4( u2_u5_u7_n142 ) , .A3( u2_u5_u7_n143 ) , .A2( u2_u5_u7_n144 ) , .A1( u2_u5_u7_n178 ) );
  OAI221_X1 u2_u5_u7_U9 (.C1( u2_u5_u7_n101 ) , .C2( u2_u5_u7_n147 ) , .ZN( u2_u5_u7_n155 ) , .B2( u2_u5_u7_n162 ) , .A( u2_u5_u7_n91 ) , .B1( u2_u5_u7_n92 ) );
  OR2_X1 u2_u5_u7_U90 (.A2( u2_u5_u7_n125 ) , .A1( u2_u5_u7_n129 ) , .ZN( u2_u5_u7_n144 ) );
  AOI22_X1 u2_u5_u7_U91 (.A2( u2_u5_u7_n126 ) , .ZN( u2_u5_u7_n143 ) , .B2( u2_u5_u7_n165 ) , .B1( u2_u5_u7_n173 ) , .A1( u2_u5_u7_n174 ) );
  NAND4_X1 u2_u5_u7_U92 (.ZN( u2_out5_5 ) , .A4( u2_u5_u7_n108 ) , .A3( u2_u5_u7_n109 ) , .A1( u2_u5_u7_n116 ) , .A2( u2_u5_u7_n123 ) );
  AOI22_X1 u2_u5_u7_U93 (.ZN( u2_u5_u7_n109 ) , .A2( u2_u5_u7_n126 ) , .B2( u2_u5_u7_n145 ) , .B1( u2_u5_u7_n156 ) , .A1( u2_u5_u7_n171 ) );
  NOR4_X1 u2_u5_u7_U94 (.A4( u2_u5_u7_n104 ) , .A3( u2_u5_u7_n105 ) , .A2( u2_u5_u7_n106 ) , .A1( u2_u5_u7_n107 ) , .ZN( u2_u5_u7_n108 ) );
  NAND3_X1 u2_u5_u7_U95 (.A3( u2_u5_u7_n146 ) , .A2( u2_u5_u7_n147 ) , .A1( u2_u5_u7_n148 ) , .ZN( u2_u5_u7_n151 ) );
  NAND3_X1 u2_u5_u7_U96 (.A3( u2_u5_u7_n131 ) , .A2( u2_u5_u7_n132 ) , .A1( u2_u5_u7_n133 ) , .ZN( u2_u5_u7_n135 ) );
  AOI22_X1 u2_uk_U100 (.B2( u2_uk_K_r9_19 ) , .A2( u2_uk_K_r9_25 ) , .B1( u2_uk_n118 ) , .A1( u2_uk_n142 ) , .ZN( u2_uk_n391 ) );
  OAI21_X1 u2_uk_U1025 (.ZN( u2_K4_28 ) , .A( u2_uk_n1029 ) , .B2( u2_uk_n1351 ) , .B1( u2_uk_n17 ) );
  NAND2_X1 u2_uk_U1026 (.A1( u2_uk_K_r2_21 ) , .ZN( u2_uk_n1029 ) , .A2( u2_uk_n99 ) );
  OAI21_X1 u2_uk_U1066 (.ZN( u2_K13_28 ) , .B2( u2_uk_n1753 ) , .B1( u2_uk_n208 ) , .A( u2_uk_n662 ) );
  NAND2_X1 u2_uk_U1067 (.A1( u2_uk_K_r11_21 ) , .A2( u2_uk_n238 ) , .ZN( u2_uk_n662 ) );
  OAI21_X1 u2_uk_U1072 (.ZN( u2_K3_40 ) , .A( u2_uk_n1014 ) , .B2( u2_uk_n1300 ) , .B1( u2_uk_n230 ) );
  NAND2_X1 u2_uk_U1073 (.A1( u2_uk_K_r1_21 ) , .ZN( u2_uk_n1014 ) , .A2( u2_uk_n148 ) );
  OAI22_X1 u2_uk_U109 (.ZN( u2_K3_41 ) , .A2( u2_uk_n1283 ) , .B2( u2_uk_n1288 ) , .B1( u2_uk_n141 ) , .A1( u2_uk_n83 ) );
  INV_X1 u2_uk_U1094 (.ZN( u2_K11_8 ) , .A( u2_uk_n407 ) );
  AOI22_X1 u2_uk_U1095 (.B2( u2_uk_K_r9_12 ) , .A2( u2_uk_K_r9_18 ) , .B1( u2_uk_n118 ) , .A1( u2_uk_n230 ) , .ZN( u2_uk_n407 ) );
  INV_X1 u2_uk_U1096 (.ZN( u2_K11_12 ) , .A( u2_uk_n313 ) );
  INV_X1 u2_uk_U1128 (.ZN( u2_K6_4 ) , .A( u2_uk_n1071 ) );
  AOI22_X1 u2_uk_U1129 (.B2( u2_uk_K_r4_41 ) , .A2( u2_uk_K_r4_47 ) , .ZN( u2_uk_n1071 ) , .B1( u2_uk_n148 ) , .A1( u2_uk_n60 ) );
  AOI22_X1 u2_uk_U1154 (.B2( u2_uk_K_r4_17 ) , .A2( u2_uk_K_r4_55 ) , .ZN( u2_uk_n1066 ) , .B1( u2_uk_n148 ) , .A1( u2_uk_n63 ) );
  INV_X1 u2_uk_U1155 (.ZN( u2_K6_2 ) , .A( u2_uk_n1066 ) );
  OAI21_X1 u2_uk_U118 (.ZN( u2_K6_47 ) , .A( u2_uk_n1070 ) , .B2( u2_uk_n1419 ) , .B1( u2_uk_n60 ) );
  INV_X1 u2_uk_U134 (.ZN( u2_K13_19 ) , .A( u2_uk_n601 ) );
  AOI22_X1 u2_uk_U135 (.B2( u2_uk_K_r11_19 ) , .A2( u2_uk_K_r11_39 ) , .B1( u2_uk_n191 ) , .ZN( u2_uk_n601 ) , .A1( u2_uk_n83 ) );
  OAI22_X1 u2_uk_U136 (.ZN( u2_K11_15 ) , .A1( u2_uk_n163 ) , .B2( u2_uk_n1646 ) , .A2( u2_uk_n1661 ) , .B1( u2_uk_n63 ) );
  INV_X1 u2_uk_U149 (.ZN( u2_K11_19 ) , .A( u2_uk_n338 ) );
  AOI22_X1 u2_uk_U150 (.B2( u2_uk_K_r9_10 ) , .A2( u2_uk_K_r9_48 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n163 ) , .ZN( u2_uk_n338 ) );
  OAI21_X1 u2_uk_U154 (.ZN( u2_K3_19 ) , .A( u2_uk_n1007 ) , .B2( u2_uk_n1294 ) , .B1( u2_uk_n83 ) );
  OAI22_X1 u2_uk_U163 (.ZN( u2_K14_30 ) , .B1( u2_uk_n142 ) , .B2( u2_uk_n1781 ) , .A2( u2_uk_n1808 ) , .A1( u2_uk_n94 ) );
  INV_X1 u2_uk_U177 (.ZN( u2_K11_14 ) , .A( u2_uk_n319 ) );
  OAI21_X1 u2_uk_U190 (.ZN( u2_K13_30 ) , .B1( u2_uk_n110 ) , .B2( u2_uk_n1746 ) , .A( u2_uk_n671 ) );
  NAND2_X1 u2_uk_U191 (.A1( u2_uk_K_r11_28 ) , .A2( u2_uk_n17 ) , .ZN( u2_uk_n671 ) );
  INV_X1 u2_uk_U197 (.ZN( u2_K3_24 ) , .A( u2_uk_n1008 ) );
  AOI22_X1 u2_uk_U198 (.B2( u2_uk_K_r1_17 ) , .A2( u2_uk_K_r1_41 ) , .ZN( u2_uk_n1008 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n202 ) );
  OAI21_X1 u2_uk_U204 (.ZN( u2_K4_30 ) , .A( u2_uk_n1032 ) , .B2( u2_uk_n1345 ) , .B1( u2_uk_n187 ) );
  NAND2_X1 u2_uk_U205 (.A1( u2_uk_K_r2_28 ) , .ZN( u2_uk_n1032 ) , .A2( u2_uk_n148 ) );
  INV_X1 u2_uk_U209 (.ZN( u2_K4_31 ) , .A( u2_uk_n1033 ) );
  AOI22_X1 u2_uk_U210 (.B2( u2_uk_K_r2_31 ) , .A2( u2_uk_K_r2_49 ) , .B1( u2_uk_n10 ) , .ZN( u2_uk_n1033 ) , .A1( u2_uk_n188 ) );
  OAI22_X1 u2_uk_U228 (.ZN( u2_K3_31 ) , .B1( u2_uk_n110 ) , .B2( u2_uk_n1303 ) , .A2( u2_uk_n1309 ) , .A1( u2_uk_n213 ) );
  OAI22_X1 u2_uk_U269 (.ZN( u2_K6_44 ) , .B2( u2_uk_n1428 ) , .A2( u2_uk_n1446 ) , .B1( u2_uk_n182 ) , .A1( u2_uk_n93 ) );
  OAI22_X1 u2_uk_U270 (.ZN( u2_K6_48 ) , .B2( u2_uk_n1433 ) , .A2( u2_uk_n1440 ) , .A1( u2_uk_n222 ) , .B1( u2_uk_n60 ) );
  OAI21_X1 u2_uk_U272 (.ZN( u2_K3_44 ) , .A( u2_uk_n1015 ) , .B1( u2_uk_n109 ) , .B2( u2_uk_n1284 ) );
  NAND2_X1 u2_uk_U273 (.A1( u2_uk_K_r1_15 ) , .ZN( u2_uk_n1015 ) , .A2( u2_uk_n60 ) );
  OAI22_X1 u2_uk_U280 (.ZN( u2_K6_6 ) , .B2( u2_uk_n1444 ) , .A2( u2_uk_n1448 ) , .A1( u2_uk_n162 ) , .B1( u2_uk_n60 ) );
  OAI21_X1 u2_uk_U281 (.ZN( u2_K6_8 ) , .A( u2_uk_n1073 ) , .B2( u2_uk_n1416 ) , .B1( u2_uk_n31 ) );
  INV_X1 u2_uk_U303 (.ZN( u2_K4_26 ) , .A( u2_uk_n1028 ) );
  OAI22_X1 u2_uk_U316 (.ZN( u2_K14_26 ) , .B2( u2_uk_n1792 ) , .A2( u2_uk_n1809 ) , .A1( u2_uk_n191 ) , .B1( u2_uk_n63 ) );
  OAI22_X1 u2_uk_U320 (.ZN( u2_K3_26 ) , .B2( u2_uk_n1299 ) , .A2( u2_uk_n1315 ) , .B1( u2_uk_n141 ) , .A1( u2_uk_n92 ) );
  OAI21_X1 u2_uk_U326 (.ZN( u2_K3_46 ) , .A( u2_uk_n1017 ) , .B2( u2_uk_n1297 ) , .B1( u2_uk_n202 ) );
  NAND2_X1 u2_uk_U327 (.A1( u2_uk_K_r1_22 ) , .ZN( u2_uk_n1017 ) , .A2( u2_uk_n148 ) );
  OAI22_X1 u2_uk_U360 (.ZN( u2_K4_40 ) , .B2( u2_uk_n1342 ) , .A2( u2_uk_n1352 ) , .A1( u2_uk_n146 ) , .B1( u2_uk_n31 ) );
  OAI22_X1 u2_uk_U373 (.ZN( u2_K3_28 ) , .B2( u2_uk_n1298 ) , .A2( u2_uk_n1303 ) , .A1( u2_uk_n162 ) , .B1( u2_uk_n99 ) );
  INV_X1 u2_uk_U424 (.ZN( u2_K6_9 ) , .A( u2_uk_n1074 ) );
  OAI22_X1 u2_uk_U431 (.ZN( u2_K11_1 ) , .A1( u2_uk_n163 ) , .B2( u2_uk_n1658 ) , .A2( u2_uk_n1675 ) , .B1( u2_uk_n63 ) );
  OAI22_X1 u2_uk_U438 (.ZN( u2_K4_37 ) , .A1( u2_uk_n118 ) , .B2( u2_uk_n1331 ) , .A2( u2_uk_n1345 ) , .B1( u2_uk_n238 ) );
  OAI22_X1 u2_uk_U454 (.ZN( u2_K13_33 ) , .B2( u2_uk_n1723 ) , .A2( u2_uk_n1728 ) , .B1( u2_uk_n223 ) , .A1( u2_uk_n92 ) );
  OAI22_X1 u2_uk_U459 (.ZN( u2_K3_33 ) , .A1( u2_uk_n128 ) , .B2( u2_uk_n1292 ) , .A2( u2_uk_n1309 ) , .B1( u2_uk_n145 ) );
  OAI22_X1 u2_uk_U471 (.ZN( u2_K3_37 ) , .B2( u2_uk_n1292 ) , .A2( u2_uk_n1298 ) , .A1( u2_uk_n202 ) , .B1( u2_uk_n92 ) );
  OAI21_X1 u2_uk_U475 (.ZN( u2_K14_29 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1807 ) , .A( u2_uk_n689 ) );
  OAI22_X1 u2_uk_U477 (.ZN( u2_K13_29 ) , .B2( u2_uk_n1742 ) , .A2( u2_uk_n1745 ) , .B1( u2_uk_n222 ) , .A1( u2_uk_n99 ) );
  INV_X1 u2_uk_U483 (.ZN( u2_K4_29 ) , .A( u2_uk_n1030 ) );
  AOI22_X1 u2_uk_U484 (.B2( u2_uk_K_r2_31 ) , .A2( u2_uk_K_r2_36 ) , .ZN( u2_uk_n1030 ) , .B1( u2_uk_n191 ) , .A1( u2_uk_n83 ) );
  OAI21_X1 u2_uk_U485 (.ZN( u2_K3_29 ) , .A( u2_uk_n1010 ) , .B2( u2_uk_n1313 ) , .B1( u2_uk_n187 ) );
  NAND2_X1 u2_uk_U486 (.A1( u2_uk_K_r1_44 ) , .ZN( u2_uk_n1010 ) , .A2( u2_uk_n223 ) );
  BUF_X1 u2_uk_U50 (.Z( u2_uk_n230 ) , .A( u2_uk_n238 ) );
  OAI22_X1 u2_uk_U520 (.ZN( u2_K11_2 ) , .B1( u2_uk_n147 ) , .B2( u2_uk_n1643 ) , .A2( u2_uk_n1677 ) , .A1( u2_uk_n93 ) );
  INV_X1 u2_uk_U544 (.ZN( u2_K11_17 ) , .A( u2_uk_n335 ) );
  AOI22_X1 u2_uk_U545 (.B2( u2_uk_K_r9_4 ) , .A2( u2_uk_K_r9_55 ) , .A1( u2_uk_n109 ) , .B1( u2_uk_n231 ) , .ZN( u2_uk_n335 ) );
  OAI22_X1 u2_uk_U550 (.ZN( u2_K13_36 ) , .B2( u2_uk_n1747 ) , .A2( u2_uk_n1753 ) , .B1( u2_uk_n202 ) , .A1( u2_uk_n99 ) );
  OAI22_X1 u2_uk_U551 (.ZN( u2_K3_36 ) , .B2( u2_uk_n1279 ) , .A1( u2_uk_n128 ) , .A2( u2_uk_n1314 ) , .B1( u2_uk_n145 ) );
  OAI21_X1 u2_uk_U574 (.ZN( u2_K11_10 ) , .B2( u2_uk_n1633 ) , .A( u2_uk_n312 ) , .B1( u2_uk_n83 ) );
  NAND2_X1 u2_uk_U575 (.A1( u2_uk_K_r9_54 ) , .A2( u2_uk_n31 ) , .ZN( u2_uk_n312 ) );
  INV_X1 u2_uk_U582 (.ZN( u2_K6_10 ) , .A( u2_uk_n1058 ) );
  AOI22_X1 u2_uk_U583 (.B2( u2_uk_K_r4_3 ) , .A2( u2_uk_K_r4_54 ) , .ZN( u2_uk_n1058 ) , .B1( u2_uk_n118 ) , .A1( u2_uk_n148 ) );
  OAI22_X1 u2_uk_U587 (.ZN( u2_K3_22 ) , .B2( u2_uk_n1281 ) , .A2( u2_uk_n1316 ) , .B1( u2_uk_n141 ) , .A1( u2_uk_n94 ) );
  INV_X1 u2_uk_U589 (.ZN( u2_K13_22 ) , .A( u2_uk_n634 ) );
  AOI22_X1 u2_uk_U590 (.B2( u2_uk_K_r11_10 ) , .A2( u2_uk_K_r11_47 ) , .A1( u2_uk_n207 ) , .ZN( u2_uk_n634 ) , .B1( u2_uk_n94 ) );
  INV_X1 u2_uk_U591 (.ZN( u2_K11_22 ) , .A( u2_uk_n349 ) );
  AOI22_X1 u2_uk_U592 (.B2( u2_uk_K_r9_13 ) , .A2( u2_uk_K_r9_19 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n207 ) , .ZN( u2_uk_n349 ) );
  OAI22_X1 u2_uk_U610 (.ZN( u2_K13_35 ) , .B2( u2_uk_n1734 ) , .A2( u2_uk_n1763 ) , .B1( u2_uk_n214 ) , .A1( u2_uk_n99 ) );
  NAND2_X1 u2_uk_U643 (.A1( u2_uk_K_r2_24 ) , .ZN( u2_uk_n1039 ) , .A2( u2_uk_n60 ) );
  OAI21_X1 u2_uk_U67 (.ZN( u2_K3_34 ) , .A( u2_uk_n1011 ) , .B1( u2_uk_n110 ) , .B2( u2_uk_n1299 ) );
  OAI21_X1 u2_uk_U680 (.ZN( u2_K6_7 ) , .A( u2_uk_n1072 ) , .B2( u2_uk_n1435 ) , .B1( u2_uk_n238 ) );
  NAND2_X1 u2_uk_U681 (.A1( u2_uk_K_r4_33 ) , .ZN( u2_uk_n1072 ) , .A2( u2_uk_n217 ) );
  OAI22_X1 u2_uk_U689 (.ZN( u2_K13_25 ) , .A1( u2_uk_n110 ) , .B2( u2_uk_n1735 ) , .A2( u2_uk_n1760 ) , .B1( u2_uk_n223 ) );
  INV_X1 u2_uk_U705 (.ZN( u2_K4_25 ) , .A( u2_uk_n1027 ) );
  OAI21_X1 u2_uk_U71 (.ZN( u2_K11_23 ) , .B1( u2_uk_n164 ) , .B2( u2_uk_n1668 ) , .A( u2_uk_n353 ) );
  OAI22_X1 u2_uk_U713 (.ZN( u2_K4_32 ) , .A1( u2_uk_n109 ) , .A2( u2_uk_n1326 ) , .B2( u2_uk_n1350 ) , .B1( u2_uk_n209 ) );
  NAND2_X1 u2_uk_U72 (.A1( u2_uk_K_r9_27 ) , .A2( u2_uk_n155 ) , .ZN( u2_uk_n353 ) );
  OAI21_X1 u2_uk_U741 (.ZN( u2_K14_27 ) , .B1( u2_uk_n100 ) , .B2( u2_uk_n1809 ) , .A( u2_uk_n688 ) );
  NAND2_X1 u2_uk_U742 (.A1( u2_uk_K_r12_42 ) , .A2( u2_uk_n31 ) , .ZN( u2_uk_n688 ) );
  OAI22_X1 u2_uk_U757 (.ZN( u2_K13_27 ) , .A1( u2_uk_n128 ) , .B2( u2_uk_n1724 ) , .A2( u2_uk_n1747 ) , .B1( u2_uk_n222 ) );
  OAI21_X1 u2_uk_U772 (.ZN( u2_K3_27 ) , .A( u2_uk_n1009 ) , .B2( u2_uk_n1315 ) , .B1( u2_uk_n208 ) );
  NAND2_X1 u2_uk_U773 (.A1( u2_uk_K_r1_42 ) , .ZN( u2_uk_n1009 ) , .A2( u2_uk_n188 ) );
  INV_X1 u2_uk_U776 (.ZN( u2_K13_21 ) , .A( u2_uk_n608 ) );
  INV_X1 u2_uk_U824 (.ZN( u2_K11_20 ) , .A( u2_uk_n342 ) );
  AOI22_X1 u2_uk_U825 (.B2( u2_uk_K_r9_10 ) , .A2( u2_uk_K_r9_4 ) , .A1( u2_uk_n110 ) , .B1( u2_uk_n162 ) , .ZN( u2_uk_n342 ) );
  NAND2_X1 u2_uk_U834 (.A1( u2_uk_K_r11_4 ) , .A2( u2_uk_n128 ) , .ZN( u2_uk_n672 ) );
  OAI22_X1 u2_uk_U837 (.ZN( u2_K11_3 ) , .B2( u2_uk_n1639 ) , .A2( u2_uk_n1657 ) , .A1( u2_uk_n207 ) , .B1( u2_uk_n63 ) );
  NAND2_X1 u2_uk_U841 (.A1( u2_uk_K_r3_10 ) , .ZN( u2_uk_n1056 ) , .A2( u2_uk_n60 ) );
  OAI22_X1 u2_uk_U858 (.ZN( u2_K6_5 ) , .B2( u2_uk_n1422 ) , .A2( u2_uk_n1426 ) , .A1( u2_uk_n230 ) , .B1( u2_uk_n60 ) );
  OAI22_X1 u2_uk_U867 (.ZN( u2_K6_45 ) , .A1( u2_uk_n129 ) , .B2( u2_uk_n1424 ) , .A2( u2_uk_n1429 ) , .B1( u2_uk_n60 ) );
  OAI22_X1 u2_uk_U874 (.ZN( u2_K6_12 ) , .A2( u2_uk_n1410 ) , .B2( u2_uk_n1426 ) , .A1( u2_uk_n207 ) , .B1( u2_uk_n93 ) );
  OAI22_X1 u2_uk_U877 (.ZN( u2_K13_24 ) , .B2( u2_uk_n1726 ) , .A2( u2_uk_n1767 ) , .A1( u2_uk_n202 ) , .B1( u2_uk_n92 ) );
  OAI22_X1 u2_uk_U880 (.ZN( u2_K3_21 ) , .B1( u2_uk_n109 ) , .B2( u2_uk_n1291 ) , .A2( u2_uk_n1316 ) , .A1( u2_uk_n161 ) );
  OAI22_X1 u2_uk_U893 (.ZN( u2_K4_36 ) , .B1( u2_uk_n109 ) , .B2( u2_uk_n1346 ) , .A2( u2_uk_n1351 ) , .A1( u2_uk_n161 ) );
  OAI22_X1 u2_uk_U896 (.ZN( u2_K3_25 ) , .B1( u2_uk_n117 ) , .B2( u2_uk_n1279 ) , .A2( u2_uk_n1283 ) , .A1( u2_uk_n207 ) );
  OAI22_X1 u2_uk_U903 (.ZN( u2_K3_38 ) , .B1( u2_uk_n128 ) , .A2( u2_uk_n1284 ) , .A1( u2_uk_n129 ) , .B2( u2_uk_n1300 ) );
  OAI22_X1 u2_uk_U904 (.ZN( u2_K3_39 ) , .B1( u2_uk_n118 ) , .B2( u2_uk_n1308 ) , .A2( u2_uk_n1312 ) , .A1( u2_uk_n202 ) );
  OAI22_X1 u2_uk_U907 (.ZN( u2_K13_23 ) , .A1( u2_uk_n110 ) , .B2( u2_uk_n1737 ) , .A2( u2_uk_n1767 ) , .B1( u2_uk_n223 ) );
  OAI22_X1 u2_uk_U91 (.ZN( u2_K4_41 ) , .B2( u2_uk_n1319 ) , .A2( u2_uk_n1336 ) , .B1( u2_uk_n162 ) , .A1( u2_uk_n83 ) );
  OAI22_X1 u2_uk_U920 (.ZN( u2_K11_24 ) , .B1( u2_uk_n147 ) , .B2( u2_uk_n1652 ) , .A2( u2_uk_n1657 ) , .A1( u2_uk_n93 ) );
  OAI22_X1 u2_uk_U928 (.ZN( u2_K6_46 ) , .A2( u2_uk_n1413 ) , .B2( u2_uk_n1441 ) , .B1( u2_uk_n208 ) , .A1( u2_uk_n93 ) );
  OAI22_X1 u2_uk_U954 (.ZN( u2_K6_43 ) , .B2( u2_uk_n1408 ) , .A2( u2_uk_n1447 ) , .B1( u2_uk_n182 ) , .A1( u2_uk_n93 ) );
  INV_X1 u2_uk_U99 (.ZN( u2_K11_5 ) , .A( u2_uk_n391 ) );
  OAI21_X1 u2_uk_U997 (.ZN( u2_K3_45 ) , .A( u2_uk_n1016 ) , .B1( u2_uk_n102 ) , .B2( u2_uk_n1305 ) );
  NAND2_X1 u2_uk_U998 (.A1( u2_uk_K_r1_16 ) , .ZN( u2_uk_n1016 ) , .A2( u2_uk_n27 ) );
endmodule

