module aes_aes ( clk, key, ld, rst, text_in, done, text_out );
  input clk;
  input [127:0] key;
  input ld;
  input rst;
  input [127:0] text_in;
  output done;
  output [127:0] text_out;

  wire sa00_0, sa00_1, sa00_2, sa00_3, sa00_4, sa00_5, sa00_6, sa00_7, 
       sa00_sr_0, sa00_sr_1, sa00_sr_2, sa00_sr_3, sa00_sr_4, sa00_sr_5, sa00_sr_6, sa00_sr_7, sa01_0, 
       sa01_1, sa01_2, sa01_3, sa01_4, sa01_5, sa01_6, sa01_7, sa01_sr_0, sa01_sr_1, 
       sa01_sr_2, sa01_sr_3, sa01_sr_4, sa01_sr_5, sa01_sr_6, sa01_sr_7, sa02_0, sa02_1, sa02_2, 
       sa02_3, sa02_4, sa02_5, sa02_6, sa02_7, sa02_sr_0, sa02_sr_1, sa02_sr_2, sa02_sr_3, 
       sa02_sr_4, sa02_sr_5, sa02_sr_6, sa02_sr_7, sa03_0, sa03_1, sa03_2, sa03_3, sa03_4, 
       sa03_5, sa03_6, sa03_7, sa03_sr_0, sa03_sr_1, sa03_sr_2, sa03_sr_3, sa03_sr_4, sa03_sr_5, 
       sa03_sr_6, sa03_sr_7, sa10_0, sa10_1, sa10_2, sa10_3, sa10_4, sa10_5, sa10_6, 
       sa10_7, sa10_sr_0, sa10_sr_1, sa10_sr_2, sa10_sr_3, sa10_sr_4, sa10_sr_5, sa10_sr_6, sa10_sr_7, 
       sa11_0, sa11_1, sa11_2, sa11_3, sa11_4, sa11_5, sa11_6, sa11_7, sa11_sr_0, 
       sa11_sr_1, sa11_sr_2, sa11_sr_3, sa11_sr_4, sa11_sr_5, sa11_sr_6, sa11_sr_7, sa12_0, sa12_1, 
       sa12_2, sa12_3, sa12_4, sa12_5, sa12_6, sa12_7, sa12_sr_0, sa12_sr_1, sa12_sr_2, 
       sa12_sr_3, sa12_sr_4, sa12_sr_5, sa12_sr_6, sa12_sr_7, sa13_0, sa13_1, sa13_2, sa13_3, 
       sa13_4, sa13_5, sa13_6, sa13_7, sa13_sr_0, sa13_sr_1, sa13_sr_2, sa13_sr_3, sa13_sr_4, 
       sa13_sr_5, sa13_sr_6, sa13_sr_7, sa20_0, sa20_1, sa20_2, sa20_3, sa20_4, sa20_5, 
       sa20_6, sa20_7, sa21_0, sa21_1, sa21_2, sa21_3, sa21_4, sa21_5, sa21_6, 
       sa21_7, sa21_sr_0, sa21_sr_1, sa21_sr_2, sa21_sr_3, sa21_sr_4, sa21_sr_5, sa21_sr_6, sa21_sr_7, 
       sa22_sr_0, sa22_sr_1, sa22_sr_2, sa22_sr_3, sa22_sr_4, sa22_sr_5, sa22_sr_6, sa22_sr_7, sa23_0, 
       sa23_1, sa23_2, sa23_3, sa23_4, sa23_5, sa23_6, sa23_7, sa23_sr_0, sa23_sr_1, 
       sa23_sr_2, sa23_sr_3, sa23_sr_4, sa23_sr_5, sa23_sr_6, sa23_sr_7, sa30_0, sa30_1, sa30_2, 
       sa30_3, sa30_4, sa30_5, sa30_6, sa30_7, sa30_sr_0, sa30_sr_1, sa30_sr_2, sa30_sr_3, 
       sa30_sr_4, sa30_sr_5, sa30_sr_6, sa30_sr_7, sa31_0, sa31_1, sa31_2, sa31_3, sa31_4, 
       sa31_5, sa31_6, sa31_7, sa31_sr_0, sa31_sr_1, sa31_sr_2, sa31_sr_3, sa31_sr_4, sa31_sr_5, 
       sa31_sr_6, sa31_sr_7, sa32_0, sa32_1, sa32_2, sa32_3, sa32_4, sa32_5, sa32_6, 
       sa32_7, sa32_sr_0, sa32_sr_1, sa32_sr_2, sa32_sr_3, sa32_sr_4, sa32_sr_5, sa32_sr_6, sa32_sr_7, 
       sa33_0, sa33_1, sa33_2, sa33_3, sa33_4, sa33_5, sa33_6, sa33_7, sa33_sr_0, 
       sa33_sr_1, sa33_sr_2, sa33_sr_3, sa33_sr_4, sa33_sr_5, sa33_sr_6, sa33_sr_7, u0_n268, u0_n270, 
       u0_n272, u0_n274, u0_subword_0, u0_subword_1, u0_subword_10, u0_subword_11, u0_subword_12, u0_subword_13, u0_subword_14, 
       u0_subword_15, u0_subword_16, u0_subword_17, u0_subword_18, u0_subword_19, u0_subword_2, u0_subword_20, u0_subword_21, u0_subword_22, 
       u0_subword_23, u0_subword_3, u0_subword_4, u0_subword_5, u0_subword_6, u0_subword_7, u0_subword_8, u0_subword_9, w3_0, 
       w3_1, w3_10, w3_11, w3_2, w3_24, w3_25, w3_26, w3_27, w3_28, 
       w3_29, w3_3, w3_30, w3_31, w3_4, w3_5, w3_6, w3_7, w3_8, 
       w3_9 ;

  aes_aes_die_0 u0 ( clk, key, ld, rst, text_in, done, text_out, sa00_sr_0, sa00_sr_1, sa00_sr_2, sa00_sr_3, sa00_sr_4, sa00_sr_5, sa00_sr_6, sa00_sr_7, 
      sa01_sr_0, sa01_sr_1, sa01_sr_2, sa01_sr_3, sa01_sr_4, sa01_sr_5, sa01_sr_6, sa01_sr_7, sa02_sr_0, 
      sa02_sr_1, sa02_sr_2, sa02_sr_3, sa02_sr_4, sa02_sr_5, sa02_sr_6, sa02_sr_7, sa03_sr_0, sa03_sr_1, 
      sa03_sr_2, sa03_sr_3, sa03_sr_4, sa03_sr_5, sa03_sr_6, sa03_sr_7, sa10_sr_0, sa10_sr_1, sa10_sr_2, 
      sa10_sr_3, sa10_sr_4, sa10_sr_5, sa10_sr_6, sa10_sr_7, sa11_sr_0, sa11_sr_1, sa11_sr_2, sa11_sr_3, 
      sa11_sr_4, sa11_sr_5, sa11_sr_6, sa11_sr_7, sa12_sr_0, sa12_sr_1, sa12_sr_2, sa12_sr_3, sa12_sr_4, 
      sa12_sr_5, sa12_sr_6, sa12_sr_7, sa13_sr_0, sa13_sr_1, sa13_sr_2, sa13_sr_3, sa13_sr_4, sa13_sr_5, 
      sa13_sr_6, sa13_sr_7, sa21_sr_0, sa21_sr_1, sa21_sr_2, sa21_sr_3, sa21_sr_4, sa21_sr_5, sa21_sr_6, 
      sa21_sr_7, sa22_sr_0, sa22_sr_1, sa22_sr_2, sa22_sr_3, sa22_sr_4, sa22_sr_5, sa22_sr_6, sa22_sr_7, 
      sa23_sr_0, sa23_sr_1, sa23_sr_2, sa23_sr_3, sa23_sr_4, sa23_sr_5, sa23_sr_6, sa23_sr_7, sa30_sr_0, 
      sa30_sr_1, sa30_sr_2, sa30_sr_3, sa30_sr_4, sa30_sr_5, sa30_sr_6, sa30_sr_7, sa31_sr_0, sa31_sr_1, 
      sa31_sr_2, sa31_sr_3, sa31_sr_4, sa31_sr_5, sa31_sr_6, sa31_sr_7, sa32_sr_0, sa32_sr_1, sa32_sr_2, 
      sa32_sr_3, sa32_sr_4, sa32_sr_5, sa32_sr_6, sa32_sr_7, sa33_sr_0, sa33_sr_1, sa33_sr_2, sa33_sr_3, 
      sa33_sr_4, sa33_sr_5, sa33_sr_6, sa33_sr_7, u0_subword_0, u0_subword_1, u0_subword_10, u0_subword_11, u0_subword_12, 
      u0_subword_13, u0_subword_14, u0_subword_15, u0_subword_16, u0_subword_17, u0_subword_18, u0_subword_19, u0_subword_2, u0_subword_20, 
      u0_subword_21, u0_subword_22, u0_subword_23, u0_subword_3, u0_subword_4, u0_subword_5, u0_subword_6, u0_subword_7, u0_subword_8, 
      u0_subword_9, sa00_0, sa00_1, sa00_2, sa00_3, sa00_4, sa00_5, sa00_6, sa00_7, 
      sa01_0, sa01_1, sa01_2, sa01_3, sa01_4, sa01_5, sa01_6, sa01_7, sa02_0, 
      sa02_1, sa02_2, sa02_3, sa02_4, sa02_5, sa02_6, sa02_7, sa03_0, sa03_1, 
      sa03_2, sa03_3, sa03_4, sa03_5, sa03_6, sa03_7, sa10_0, sa10_1, sa10_2, 
      sa10_3, sa10_4, sa10_5, sa10_6, sa10_7, sa11_0, sa11_1, sa11_2, sa11_3, 
      sa11_4, sa11_5, sa11_6, sa11_7, sa12_0, sa12_1, sa12_2, sa12_3, sa12_4, 
      sa12_5, sa12_6, sa12_7, sa13_0, sa13_1, sa13_2, sa13_3, sa13_4, sa13_5, 
      sa13_6, sa13_7, sa20_0, sa20_1, sa20_2, sa20_3, sa20_4, sa20_5, sa20_6, 
      sa20_7, sa21_0, sa21_1, sa21_2, sa21_3, sa21_4, sa21_5, sa21_6, sa21_7, 
      sa23_0, sa23_1, sa23_2, sa23_3, sa23_4, sa23_5, sa23_6, sa23_7, sa30_0, 
      sa30_1, sa30_2, sa30_3, sa30_4, sa30_5, sa30_6, sa30_7, sa31_0, sa31_1, 
      sa31_2, sa31_3, sa31_4, sa31_5, sa31_6, sa31_7, sa32_0, sa32_1, sa32_2, 
      sa32_3, sa32_4, sa32_5, sa32_6, sa32_7, sa33_0, sa33_1, sa33_2, sa33_3, 
      sa33_4, sa33_5, sa33_6, sa33_7, u0_n268, u0_n270, u0_n272, u0_n274, w3_0, 
      w3_1, w3_10, w3_11, w3_2, w3_24, w3_25, w3_26, w3_27, w3_28, 
      w3_29, w3_3, w3_30, w3_31, w3_4, w3_5, w3_6, w3_7, w3_8, 
      w3_9 );
  aes_aes_die_1 u1 ( sa00_0, sa00_1, sa00_2, sa00_3, sa00_4, sa00_5, sa00_6, sa00_7, sa03_0, 
      sa03_1, sa03_2, sa03_3, sa03_4, sa03_5, sa03_6, sa03_7, sa12_0, sa12_1, 
      sa12_2, sa12_3, sa12_4, sa12_5, sa12_6, sa12_7, sa31_0, sa31_1, sa31_2, 
      sa31_3, sa31_4, sa31_5, sa31_6, sa31_7, w3_0, w3_1, w3_2, w3_24, 
      w3_25, w3_26, w3_27, w3_28, w3_29, w3_3, w3_30, w3_31, w3_4, 
      w3_5, w3_6, w3_7, sa00_sr_0, sa00_sr_1, sa00_sr_2, sa00_sr_3, sa00_sr_4, sa00_sr_5, 
      sa00_sr_6, sa00_sr_7, sa03_sr_0, sa03_sr_1, sa03_sr_2, sa03_sr_3, sa03_sr_4, sa03_sr_5, sa03_sr_6, 
      sa03_sr_7, sa11_sr_0, sa11_sr_1, sa11_sr_2, sa11_sr_3, sa11_sr_4, sa11_sr_5, sa11_sr_6, sa11_sr_7, 
      sa32_sr_0, sa32_sr_1, sa32_sr_2, sa32_sr_3, sa32_sr_4, sa32_sr_5, sa32_sr_6, sa32_sr_7, u0_subword_0, 
      u0_subword_1, u0_subword_10, u0_subword_11, u0_subword_12, u0_subword_13, u0_subword_14, u0_subword_15, u0_subword_2, u0_subword_3, 
      u0_subword_4, u0_subword_5, u0_subword_6, u0_subword_7, u0_subword_8, u0_subword_9 );
  aes_aes_die_2 u2 ( sa01_0, sa01_1, sa01_2, sa01_3, sa01_4, sa01_5, sa01_6, sa01_7, sa10_0, 
      sa10_1, sa10_2, sa10_3, sa10_4, sa10_5, sa10_6, sa10_7, sa11_0, sa11_1, 
      sa11_2, sa11_3, sa11_4, sa11_5, sa11_6, sa11_7, sa13_0, sa13_1, sa13_2, 
      sa13_3, sa13_4, sa13_5, sa13_6, sa13_7, sa20_0, sa20_1, sa20_2, sa20_3, 
      sa20_4, sa20_5, sa20_6, sa20_7, sa33_0, sa33_1, sa33_2, sa33_3, sa33_4, 
      sa33_5, sa33_6, sa33_7, sa01_sr_0, sa01_sr_1, sa01_sr_2, sa01_sr_3, sa01_sr_4, sa01_sr_5, 
      sa01_sr_6, sa01_sr_7, sa10_sr_0, sa10_sr_1, sa10_sr_2, sa10_sr_3, sa10_sr_4, sa10_sr_5, sa10_sr_6, 
      sa10_sr_7, sa12_sr_0, sa12_sr_1, sa12_sr_2, sa12_sr_3, sa12_sr_4, sa12_sr_5, sa12_sr_6, sa12_sr_7, 
      sa13_sr_0, sa13_sr_1, sa13_sr_2, sa13_sr_3, sa13_sr_4, sa13_sr_5, sa13_sr_6, sa13_sr_7, sa22_sr_0, 
      sa22_sr_1, sa22_sr_2, sa22_sr_3, sa22_sr_4, sa22_sr_5, sa22_sr_6, sa22_sr_7, sa30_sr_0, sa30_sr_1, 
      sa30_sr_2, sa30_sr_3, sa30_sr_4, sa30_sr_5, sa30_sr_6, sa30_sr_7 );
  aes_aes_die_3 u3 ( sa02_0, sa02_1, sa02_2, sa02_3, sa02_4, sa02_5, sa02_6, sa02_7, sa21_0, 
      sa21_1, sa21_2, sa21_3, sa21_4, sa21_5, sa21_6, sa21_7, sa23_0, sa23_1, 
      sa23_2, sa23_3, sa23_4, sa23_5, sa23_6, sa23_7, sa30_0, sa30_1, sa30_2, 
      sa30_3, sa30_4, sa30_5, sa30_6, sa30_7, sa32_0, sa32_1, sa32_2, sa32_3, 
      sa32_4, sa32_5, sa32_6, sa32_7, u0_n268, u0_n270, u0_n272, u0_n274, w3_10, 
      w3_11, w3_8, w3_9, sa02_sr_0, sa02_sr_1, sa02_sr_2, sa02_sr_3, sa02_sr_4, sa02_sr_5, 
      sa02_sr_6, sa02_sr_7, sa21_sr_0, sa21_sr_1, sa21_sr_2, sa21_sr_3, sa21_sr_4, sa21_sr_5, sa21_sr_6, 
      sa21_sr_7, sa23_sr_0, sa23_sr_1, sa23_sr_2, sa23_sr_3, sa23_sr_4, sa23_sr_5, sa23_sr_6, sa23_sr_7, 
      sa31_sr_0, sa31_sr_1, sa31_sr_2, sa31_sr_3, sa31_sr_4, sa31_sr_5, sa31_sr_6, sa31_sr_7, sa33_sr_0, 
      sa33_sr_1, sa33_sr_2, sa33_sr_3, sa33_sr_4, sa33_sr_5, sa33_sr_6, sa33_sr_7, u0_subword_16, u0_subword_17, 
      u0_subword_18, u0_subword_19, u0_subword_20, u0_subword_21, u0_subword_22, u0_subword_23 );
endmodule
module aes_aes_die_0 ( clk, key, ld, rst, text_in, done, text_out, sa00_sr_0, sa00_sr_1, 
       sa00_sr_2, sa00_sr_3, sa00_sr_4, sa00_sr_5, sa00_sr_6, sa00_sr_7, sa01_sr_0, sa01_sr_1, sa01_sr_2, 
       sa01_sr_3, sa01_sr_4, sa01_sr_5, sa01_sr_6, sa01_sr_7, sa02_sr_0, sa02_sr_1, sa02_sr_2, sa02_sr_3, 
       sa02_sr_4, sa02_sr_5, sa02_sr_6, sa02_sr_7, sa03_sr_0, sa03_sr_1, sa03_sr_2, sa03_sr_3, sa03_sr_4, 
       sa03_sr_5, sa03_sr_6, sa03_sr_7, sa10_sr_0, sa10_sr_1, sa10_sr_2, sa10_sr_3, sa10_sr_4, sa10_sr_5, 
       sa10_sr_6, sa10_sr_7, sa11_sr_0, sa11_sr_1, sa11_sr_2, sa11_sr_3, sa11_sr_4, sa11_sr_5, sa11_sr_6, 
       sa11_sr_7, sa12_sr_0, sa12_sr_1, sa12_sr_2, sa12_sr_3, sa12_sr_4, sa12_sr_5, sa12_sr_6, sa12_sr_7, 
       sa13_sr_0, sa13_sr_1, sa13_sr_2, sa13_sr_3, sa13_sr_4, sa13_sr_5, sa13_sr_6, sa13_sr_7, sa21_sr_0, 
       sa21_sr_1, sa21_sr_2, sa21_sr_3, sa21_sr_4, sa21_sr_5, sa21_sr_6, sa21_sr_7, sa22_sr_0, sa22_sr_1, 
       sa22_sr_2, sa22_sr_3, sa22_sr_4, sa22_sr_5, sa22_sr_6, sa22_sr_7, sa23_sr_0, sa23_sr_1, sa23_sr_2, 
       sa23_sr_3, sa23_sr_4, sa23_sr_5, sa23_sr_6, sa23_sr_7, sa30_sr_0, sa30_sr_1, sa30_sr_2, sa30_sr_3, 
       sa30_sr_4, sa30_sr_5, sa30_sr_6, sa30_sr_7, sa31_sr_0, sa31_sr_1, sa31_sr_2, sa31_sr_3, sa31_sr_4, 
       sa31_sr_5, sa31_sr_6, sa31_sr_7, sa32_sr_0, sa32_sr_1, sa32_sr_2, sa32_sr_3, sa32_sr_4, sa32_sr_5, 
       sa32_sr_6, sa32_sr_7, sa33_sr_0, sa33_sr_1, sa33_sr_2, sa33_sr_3, sa33_sr_4, sa33_sr_5, sa33_sr_6, 
       sa33_sr_7, u0_subword_0, u0_subword_1, u0_subword_10, u0_subword_11, u0_subword_12, u0_subword_13, u0_subword_14, u0_subword_15, 
       u0_subword_16, u0_subword_17, u0_subword_18, u0_subword_19, u0_subword_2, u0_subword_20, u0_subword_21, u0_subword_22, u0_subword_23, 
       u0_subword_3, u0_subword_4, u0_subword_5, u0_subword_6, u0_subword_7, u0_subword_8, u0_subword_9, sa00_0, sa00_1, sa00_2, sa00_3, sa00_4, sa00_5, sa00_6, sa00_7, sa01_0, 
        sa01_1, sa01_2, sa01_3, sa01_4, sa01_5, sa01_6, sa01_7, sa02_0, sa02_1, 
        sa02_2, sa02_3, sa02_4, sa02_5, sa02_6, sa02_7, sa03_0, sa03_1, sa03_2, 
        sa03_3, sa03_4, sa03_5, sa03_6, sa03_7, sa10_0, sa10_1, sa10_2, sa10_3, 
        sa10_4, sa10_5, sa10_6, sa10_7, sa11_0, sa11_1, sa11_2, sa11_3, sa11_4, 
        sa11_5, sa11_6, sa11_7, sa12_0, sa12_1, sa12_2, sa12_3, sa12_4, sa12_5, 
        sa12_6, sa12_7, sa13_0, sa13_1, sa13_2, sa13_3, sa13_4, sa13_5, sa13_6, 
        sa13_7, sa20_0, sa20_1, sa20_2, sa20_3, sa20_4, sa20_5, sa20_6, sa20_7, 
        sa21_0, sa21_1, sa21_2, sa21_3, sa21_4, sa21_5, sa21_6, sa21_7, sa23_0, 
        sa23_1, sa23_2, sa23_3, sa23_4, sa23_5, sa23_6, sa23_7, sa30_0, sa30_1, 
        sa30_2, sa30_3, sa30_4, sa30_5, sa30_6, sa30_7, sa31_0, sa31_1, sa31_2, 
        sa31_3, sa31_4, sa31_5, sa31_6, sa31_7, sa32_0, sa32_1, sa32_2, sa32_3, 
        sa32_4, sa32_5, sa32_6, sa32_7, sa33_0, sa33_1, sa33_2, sa33_3, sa33_4, 
        sa33_5, sa33_6, sa33_7, u0_n268, u0_n270, u0_n272, u0_n274, w3_0, w3_1, 
        w3_10, w3_11, w3_2, w3_24, w3_25, w3_26, w3_27, w3_28, w3_29, 
        w3_3, w3_30, w3_31, w3_4, w3_5, w3_6, w3_7, w3_8, w3_9 );
  input clk;
  input [127:0] key;
  input ld;
  input rst;
  input [127:0] text_in;
  output done;
  output [127:0] text_out;
  input sa00_sr_0, sa00_sr_1, sa00_sr_2, sa00_sr_3, sa00_sr_4, sa00_sr_5, sa00_sr_6, sa00_sr_7, sa01_sr_0, 
        sa01_sr_1, sa01_sr_2, sa01_sr_3, sa01_sr_4, sa01_sr_5, sa01_sr_6, sa01_sr_7, sa02_sr_0, sa02_sr_1, 
        sa02_sr_2, sa02_sr_3, sa02_sr_4, sa02_sr_5, sa02_sr_6, sa02_sr_7, sa03_sr_0, sa03_sr_1, sa03_sr_2, 
        sa03_sr_3, sa03_sr_4, sa03_sr_5, sa03_sr_6, sa03_sr_7, sa10_sr_0, sa10_sr_1, sa10_sr_2, sa10_sr_3, 
        sa10_sr_4, sa10_sr_5, sa10_sr_6, sa10_sr_7, sa11_sr_0, sa11_sr_1, sa11_sr_2, sa11_sr_3, sa11_sr_4, 
        sa11_sr_5, sa11_sr_6, sa11_sr_7, sa12_sr_0, sa12_sr_1, sa12_sr_2, sa12_sr_3, sa12_sr_4, sa12_sr_5, 
        sa12_sr_6, sa12_sr_7, sa13_sr_0, sa13_sr_1, sa13_sr_2, sa13_sr_3, sa13_sr_4, sa13_sr_5, sa13_sr_6, 
        sa13_sr_7, sa21_sr_0, sa21_sr_1, sa21_sr_2, sa21_sr_3, sa21_sr_4, sa21_sr_5, sa21_sr_6, sa21_sr_7, 
        sa22_sr_0, sa22_sr_1, sa22_sr_2, sa22_sr_3, sa22_sr_4, sa22_sr_5, sa22_sr_6, sa22_sr_7, sa23_sr_0, 
        sa23_sr_1, sa23_sr_2, sa23_sr_3, sa23_sr_4, sa23_sr_5, sa23_sr_6, sa23_sr_7, sa30_sr_0, sa30_sr_1, 
        sa30_sr_2, sa30_sr_3, sa30_sr_4, sa30_sr_5, sa30_sr_6, sa30_sr_7, sa31_sr_0, sa31_sr_1, sa31_sr_2, 
        sa31_sr_3, sa31_sr_4, sa31_sr_5, sa31_sr_6, sa31_sr_7, sa32_sr_0, sa32_sr_1, sa32_sr_2, sa32_sr_3, 
        sa32_sr_4, sa32_sr_5, sa32_sr_6, sa32_sr_7, sa33_sr_0, sa33_sr_1, sa33_sr_2, sa33_sr_3, sa33_sr_4, 
        sa33_sr_5, sa33_sr_6, sa33_sr_7, u0_subword_0, u0_subword_1, u0_subword_10, u0_subword_11, u0_subword_12, u0_subword_13, 
        u0_subword_14, u0_subword_15, u0_subword_16, u0_subword_17, u0_subword_18, u0_subword_19, u0_subword_2, u0_subword_20, u0_subword_21, 
        u0_subword_22, u0_subword_23, u0_subword_3, u0_subword_4, u0_subword_5, u0_subword_6, u0_subword_7, u0_subword_8, u0_subword_9;
  output sa00_0, sa00_1, sa00_2, sa00_3, sa00_4, sa00_5, sa00_6, sa00_7, sa01_0, 
        sa01_1, sa01_2, sa01_3, sa01_4, sa01_5, sa01_6, sa01_7, sa02_0, sa02_1, 
        sa02_2, sa02_3, sa02_4, sa02_5, sa02_6, sa02_7, sa03_0, sa03_1, sa03_2, 
        sa03_3, sa03_4, sa03_5, sa03_6, sa03_7, sa10_0, sa10_1, sa10_2, sa10_3, 
        sa10_4, sa10_5, sa10_6, sa10_7, sa11_0, sa11_1, sa11_2, sa11_3, sa11_4, 
        sa11_5, sa11_6, sa11_7, sa12_0, sa12_1, sa12_2, sa12_3, sa12_4, sa12_5, 
        sa12_6, sa12_7, sa13_0, sa13_1, sa13_2, sa13_3, sa13_4, sa13_5, sa13_6, 
        sa13_7, sa20_0, sa20_1, sa20_2, sa20_3, sa20_4, sa20_5, sa20_6, sa20_7, 
        sa21_0, sa21_1, sa21_2, sa21_3, sa21_4, sa21_5, sa21_6, sa21_7, sa23_0, 
        sa23_1, sa23_2, sa23_3, sa23_4, sa23_5, sa23_6, sa23_7, sa30_0, sa30_1, 
        sa30_2, sa30_3, sa30_4, sa30_5, sa30_6, sa30_7, sa31_0, sa31_1, sa31_2, 
        sa31_3, sa31_4, sa31_5, sa31_6, sa31_7, sa32_0, sa32_1, sa32_2, sa32_3, 
        sa32_4, sa32_5, sa32_6, sa32_7, sa33_0, sa33_1, sa33_2, sa33_3, sa33_4, 
        sa33_5, sa33_6, sa33_7, u0_n268, u0_n270, u0_n272, u0_n274, w3_0, w3_1, 
        w3_10, w3_11, w3_2, w3_24, w3_25, w3_26, w3_27, w3_28, w3_29, 
        w3_3, w3_30, w3_31, w3_4, w3_5, w3_6, w3_7, w3_8, w3_9;
  wire N100, N101, N102, N103, N104, N105, N114, N115, N116, 
       N117, N118, N119, N120, N121, N130, N131, N132, N133, 
       N134, N135, N136, N137, N146, N147, N148, N149, N150, 
       N151, N152, N153, N162, N163, N164, N165, N166, N167, 
       N168, N169, N178, N179, N180, N181, N182, N183, N184, 
       N185, N194, N195, N196, N197, N198, N199, N200, N201, 
       N210, N211, N212, N213, N214, N215, N216, N217, N226, 
       N227, N228, N229, N23, N230, N231, N232, N233, N242, 
       N243, N244, N245, N246, N247, N248, N249, N258, N259, 
       N260, N261, N262, N263, N264, N265, N274, N275, N276, 
       N277, N278, N279, N280, N281, N34, N35, N36, N37, 
       N378, N379, N38, N380, N381, N382, N383, N384, N385, 
       N386, N387, N388, N389, N39, N390, N391, N392, N393, 
       N394, N395, N396, N397, N398, N399, N40, N400, N401, 
       N402, N403, N404, N405, N406, N407, N408, N409, N41, 
       N410, N411, N412, N413, N414, N415, N416, N417, N418, 
       N419, N420, N421, N422, N423, N424, N425, N426, N427, 
       N428, N429, N430, N431, N432, N433, N434, N435, N436, 
       N437, N438, N439, N440, N441, N442, N443, N444, N445, 
       N446, N447, N448, N449, N450, N451, N452, N453, N454, 
       N455, N456, N457, N458, N459, N460, N461, N462, N463, 
       N464, N465, N466, N467, N468, N469, N470, N471, N472, 
       N473, N474, N475, N476, N477, N478, N479, N480, N481, 
       N482, N483, N484, N485, N486, N487, N488, N489, N490, 
       N491, N492, N493, N494, N495, N496, N497, N498, N499, 
       N50, N500, N501, N502, N503, N504, N505, N51, N52, 
       N53, N54, N55, N56, N57, N66, N67, N68, N69, 
       N70, N71, N72, N73, N82, N83, N84, N85, N86, 
       N87, N88, N89, N98, N99, n1, n10, n100, n1000, 
       n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, 
       n101, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, 
       n1018, n1019, n102, n1020, n1021, n1022, n1023, n1024, n1025, 
       n1026, n1027, n1028, n1029, n103, n1030, n1031, n1032, n1033, 
       n1034, n1035, n1036, n1037, n1038, n1039, n104, n1040, n1041, 
       n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n105, 
       n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, 
       n1059, n106, n1060, n1061, n1062, n1063, n1064, n1065, n1066, 
       n1067, n1068, n1069, n107, n1070, n1071, n1072, n1073, n1074, 
       n1075, n1076, n1077, n1078, n1079, n108, n1080, n1081, n1082, 
       n1083, n1084, n1085, n1086, n1087, n1088, n1089, n109, n1090, 
       n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, 
       n11, n110, n1100, n1101, n1102, n1103, n1104, n1105, n1106, 
       n1107, n1108, n1109, n111, n1110, n1111, n1112, n1113, n1114, 
       n1115, n1116, n1117, n1118, n1119, n112, n1120, n1121, n1122, 
       n1123, n1124, n1125, n1126, n1127, n1128, n1129, n113, n1130, 
       n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, 
       n114, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, 
       n1148, n1149, n115, n1150, n1151, n1152, n1153, n1154, n1155, 
       n1156, n1157, n1158, n1159, n116, n1160, n1161, n1162, n1163, 
       n1164, n1165, n1166, n1167, n1168, n1169, n117, n1170, n1171, 
       n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n118, 
       n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, 
       n1189, n119, n1190, n1191, n1192, n1193, n1194, n1195, n1196, 
       n1197, n1198, n1199, n12, n120, n1200, n1201, n1202, n1203, 
       n1204, n1205, n1206, n1207, n1208, n1209, n121, n1210, n1211, 
       n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n122, 
       n1220, n1221, n1222, n123, n124, n125, n126, n127, n128, 
       n129, n13, n130, n131, n132, n133, n134, n135, n136, 
       n137, n138, n139, n14, n140, n141, n142, n143, n144, 
       n145, n146, n147, n148, n149, n15, n150, n151, n152, 
       n153, n154, n155, n156, n157, n158, n159, n16, n160, 
       n161, n162, n163, n164, n165, n166, n167, n168, n169, 
       n17, n170, n171, n172, n173, n174, n175, n176, n177, 
       n178, n179, n18, n180, n181, n182, n183, n184, n185, 
       n186, n187, n188, n189, n19, n190, n191, n192, n193, 
       n194, n195, n196, n197, n198, n199, n2, n20, n200, 
       n201, n202, n203, n204, n205, n206, n207, n208, n209, 
       n21, n210, n211, n212, n213, n214, n215, n216, n217, 
       n218, n219, n22, n220, n221, n222, n223, n224, n225, 
       n226, n227, n228, n229, n23, n230, n231, n232, n233, 
       n234, n235, n236, n237, n238, n239, n24, n240, n241, 
       n242, n243, n244, n245, n246, n247, n248, n249, n25, 
       n250, n251, n252, n253, n254, n255, n256, n258, n259, 
       n26, n260, n261, n262, n263, n264, n265, n266, n267, 
       n268, n269, n27, n270, n271, n272, n275, n276, n277, 
       n278, n279, n28, n280, n281, n283, n284, n285, n286, 
       n288, n289, n29, n290, n291, n292, n294, n295, n296, 
       n297, n298, n3, n30, n300, n301, n302, n303, n304, 
       n305, n306, n307, n308, n309, n31, n310, n311, n312, 
       n314, n315, n316, n317, n318, n319, n32, n321, n322, 
       n323, n324, n325, n327, n328, n329, n33, n330, n331, 
       n332, n334, n335, n336, n337, n338, n339, n34, n341, 
       n342, n343, n345, n347, n348, n349, n35, n350, n351, 
       n352, n353, n354, n355, n356, n357, n358, n359, n36, 
       n360, n361, n362, n363, n365, n366, n367, n368, n369, 
       n37, n370, n372, n373, n374, n375, n376, n378, n379, 
       n38, n380, n381, n382, n384, n385, n386, n387, n388, 
       n39, n390, n391, n392, n394, n395, n396, n398, n399, 
       n4, n40, n400, n401, n402, n403, n404, n405, n407, 
       n408, n409, n41, n410, n412, n413, n414, n416, n417, 
       n418, n419, n42, n421, n422, n423, n424, n425, n426, 
       n427, n428, n429, n43, n431, n432, n433, n434, n436, 
       n437, n438, n439, n44, n440, n441, n442, n443, n444, 
       n445, n446, n448, n449, n45, n450, n451, n452, n453, 
       n454, n455, n456, n457, n459, n46, n460, n461, n462, 
       n464, n465, n466, n468, n469, n47, n470, n471, n472, 
       n473, n475, n476, n477, n478, n479, n48, n481, n482, 
       n483, n484, n485, n486, n487, n488, n489, n49, n490, 
       n491, n492, n493, n495, n496, n497, n498, n499, n5, 
       n50, n500, n502, n503, n504, n505, n506, n508, n509, 
       n51, n510, n511, n512, n513, n515, n516, n517, n518, 
       n519, n52, n520, n521, n522, n523, n524, n526, n528, 
       n529, n53, n530, n531, n532, n533, n534, n535, n536, 
       n537, n538, n539, n54, n540, n541, n542, n543, n544, 
       n546, n547, n548, n55, n550, n551, n552, n554, n555, 
       n556, n557, n558, n56, n560, n561, n562, n564, n565, 
       n566, n568, n569, n57, n570, n571, n572, n573, n574, 
       n575, n576, n577, n578, n579, n58, n581, n582, n583, 
       n584, n586, n587, n588, n59, n590, n591, n592, n593, 
       n595, n596, n597, n598, n599, n6, n60, n600, n601, 
       n602, n603, n605, n606, n607, n608, n609, n61, n610, 
       n611, n612, n613, n614, n615, n616, n617, n618, n619, 
       n62, n620, n622, n623, n624, n625, n626, n628, n629, 
       n63, n630, n632, n633, n634, n635, n636, n638, n639, 
       n64, n640, n642, n643, n644, n645, n646, n647, n649, 
       n65, n650, n651, n652, n653, n655, n656, n657, n658, 
       n659, n66, n660, n661, n662, n663, n664, n665, n666, 
       n667, n669, n67, n670, n671, n672, n673, n674, n676, 
       n677, n678, n679, n68, n680, n682, n683, n684, n685, 
       n686, n687, n689, n69, n690, n691, n692, n693, n694, 
       n696, n697, n698, n7, n70, n700, n702, n703, n704, 
       n705, n706, n707, n708, n709, n71, n710, n711, n712, 
       n713, n714, n715, n716, n718, n719, n72, n720, n721, 
       n722, n724, n725, n726, n728, n729, n73, n730, n731, 
       n732, n734, n735, n736, n738, n739, n74, n740, n742, 
       n743, n744, n745, n746, n747, n748, n749, n75, n750, 
       n751, n752, n753, n755, n756, n757, n758, n76, n760, 
       n761, n762, n764, n765, n766, n767, n769, n77, n770, 
       n771, n772, n773, n774, n775, n776, n777, n778, n779, 
       n78, n780, n781, n782, n783, n784, n785, n786, n787, 
       n788, n789, n79, n790, n791, n792, n793, n794, n796, 
       n797, n798, n799, n8, n80, n800, n801, n802, n803, 
       n804, n806, n807, n808, n809, n81, n810, n812, n813, 
       n814, n816, n817, n818, n819, n82, n820, n821, n823, 
       n824, n825, n826, n827, n828, n829, n83, n830, n831, 
       n832, n833, n834, n835, n836, n837, n838, n839, n84, 
       n840, n841, n843, n844, n845, n846, n847, n848, n85, 
       n850, n851, n852, n853, n854, n856, n857, n858, n859, 
       n86, n861, n862, n863, n864, n865, n866, n867, n868, 
       n869, n87, n870, n872, n874, n875, n876, n877, n878, 
       n879, n88, n880, n881, n882, n883, n884, n885, n886, 
       n887, n888, n889, n89, n890, n892, n893, n894, n896, 
       n898, n899, n9, n90, n900, n901, n902, n903, n904, 
       n905, n907, n908, n909, n91, n911, n912, n913, n915, 
       n916, n917, n918, n919, n92, n920, n921, n922, n923, 
       n924, n925, n926, n927, n929, n93, n930, n931, n932, 
       n933, n935, n936, n937, n939, n94, n940, n941, n942, 
       n944, n945, n946, n947, n948, n949, n95, n950, n951, 
       n952, n954, n955, n956, n957, n958, n959, n96, n960, 
       n961, n962, n964, n965, n966, n967, n969, n97, n970, 
       n971, n972, n973, n974, n975, n976, n977, n978, n979, 
       n98, n980, n981, n982, n983, n984, n985, n986, n987, 
       n988, n989, n99, n990, n991, n992, n993, n994, n995, 
       n996, n997, n998, n999, sa20_sr_0, sa20_sr_1, sa20_sr_2, sa20_sr_3, sa20_sr_4, 
       sa20_sr_5, sa20_sr_6, sa20_sr_7, sa22_0, sa22_1, sa22_2, sa22_3, sa22_4, sa22_5, 
       sa22_6, sa22_7, u0_N108, u0_N109, u0_N110, u0_N111, u0_N112, u0_N113, u0_N114, 
       u0_N115, u0_N116, u0_N117, u0_N118, u0_N119, u0_N120, u0_N121, u0_N122, u0_N123, 
       u0_N124, u0_N125, u0_N126, u0_N127, u0_N128, u0_N129, u0_N130, u0_N131, u0_N132, 
       u0_N133, u0_N134, u0_N135, u0_N136, u0_N137, u0_N138, u0_N139, u0_N174, u0_N175, 
       u0_N176, u0_N177, u0_N178, u0_N179, u0_N180, u0_N181, u0_N182, u0_N183, u0_N184, 
       u0_N185, u0_N186, u0_N187, u0_N188, u0_N189, u0_N190, u0_N191, u0_N192, u0_N193, 
       u0_N194, u0_N195, u0_N196, u0_N197, u0_N198, u0_N199, u0_N200, u0_N201, u0_N202, 
       u0_N203, u0_N204, u0_N205, u0_N240, u0_N241, u0_N242, u0_N243, u0_N244, u0_N245, 
       u0_N246, u0_N247, u0_N248, u0_N249, u0_N250, u0_N251, u0_N252, u0_N253, u0_N254, 
       u0_N255, u0_N256, u0_N257, u0_N258, u0_N259, u0_N260, u0_N261, u0_N262, u0_N263, 
       u0_N264, u0_N265, u0_N266, u0_N267, u0_N268, u0_N269, u0_N270, u0_N271, u0_N42, 
       u0_N43, u0_N44, u0_N45, u0_N46, u0_N47, u0_N48, u0_N49, u0_N50, u0_N51, 
       u0_N52, u0_N53, u0_N54, u0_N55, u0_N56, u0_N57, u0_N58, u0_N59, u0_N60, 
       u0_N61, u0_N62, u0_N63, u0_N64, u0_N65, u0_N66, u0_N67, u0_N68, u0_N69, 
       u0_N70, u0_N71, u0_N72, u0_N73, u0_n1, u0_n10, u0_n100, u0_n101, u0_n102, 
       u0_n103, u0_n104, u0_n105, u0_n106, u0_n107, u0_n108, u0_n109, u0_n11, u0_n110, 
       u0_n111, u0_n112, u0_n113, u0_n114, u0_n115, u0_n116, u0_n117, u0_n118, u0_n119, 
       u0_n12, u0_n120, u0_n121, u0_n122, u0_n123, u0_n124, u0_n125, u0_n126, u0_n127, 
       u0_n128, u0_n129, u0_n13, u0_n130, u0_n131, u0_n132, u0_n133, u0_n134, u0_n135, 
       u0_n136, u0_n137, u0_n138, u0_n139, u0_n14, u0_n140, u0_n141, u0_n142, u0_n143, 
       u0_n144, u0_n145, u0_n146, u0_n147, u0_n148, u0_n149, u0_n15, u0_n150, u0_n151, 
       u0_n152, u0_n153, u0_n154, u0_n155, u0_n156, u0_n157, u0_n158, u0_n159, u0_n16, 
       u0_n160, u0_n161, u0_n162, u0_n163, u0_n164, u0_n165, u0_n166, u0_n167, u0_n168, 
       u0_n169, u0_n17, u0_n170, u0_n171, u0_n172, u0_n173, u0_n174, u0_n175, u0_n176, 
       u0_n177, u0_n178, u0_n179, u0_n18, u0_n180, u0_n181, u0_n182, u0_n183, u0_n184, 
       u0_n185, u0_n186, u0_n187, u0_n188, u0_n189, u0_n19, u0_n190, u0_n191, u0_n192, 
       u0_n193, u0_n194, u0_n195, u0_n196, u0_n197, u0_n198, u0_n199, u0_n2, u0_n20, 
       u0_n200, u0_n201, u0_n202, u0_n203, u0_n204, u0_n205, u0_n206, u0_n207, u0_n208, 
       u0_n209, u0_n21, u0_n210, u0_n211, u0_n212, u0_n213, u0_n214, u0_n215, u0_n216, 
       u0_n217, u0_n218, u0_n219, u0_n22, u0_n220, u0_n221, u0_n222, u0_n223, u0_n224, 
       u0_n225, u0_n226, u0_n227, u0_n228, u0_n229, u0_n23, u0_n230, u0_n231, u0_n232, 
       u0_n233, u0_n234, u0_n235, u0_n236, u0_n237, u0_n238, u0_n239, u0_n24, u0_n240, 
       u0_n241, u0_n242, u0_n243, u0_n244, u0_n245, u0_n246, u0_n247, u0_n248, u0_n249, 
       u0_n25, u0_n250, u0_n251, u0_n253, u0_n254, u0_n255, u0_n257, u0_n258, u0_n259, 
       u0_n26, u0_n261, u0_n262, u0_n263, u0_n264, u0_n265, u0_n267, u0_n269, u0_n27, 
       u0_n271, u0_n273, u0_n275, u0_n277, u0_n279, u0_n28, u0_n281, u0_n283, u0_n285, 
       u0_n287, u0_n29, u0_n3, u0_n30, u0_n31, u0_n32, u0_n33, u0_n34, u0_n35, 
       u0_n36, u0_n37, u0_n38, u0_n39, u0_n4, u0_n40, u0_n41, u0_n42, u0_n43, 
       u0_n44, u0_n45, u0_n46, u0_n47, u0_n48, u0_n49, u0_n5, u0_n50, u0_n51, 
       u0_n52, u0_n53, u0_n54, u0_n55, u0_n56, u0_n57, u0_n58, u0_n59, u0_n6, 
       u0_n60, u0_n61, u0_n62, u0_n63, u0_n64, u0_n65, u0_n66, u0_n67, u0_n68, 
       u0_n69, u0_n7, u0_n70, u0_n71, u0_n72, u0_n73, u0_n74, u0_n75, u0_n76, 
       u0_n77, u0_n78, u0_n79, u0_n8, u0_n80, u0_n81, u0_n82, u0_n83, u0_n84, 
       u0_n85, u0_n86, u0_n87, u0_n88, u0_n89, u0_n9, u0_n90, u0_n91, u0_n92, 
       u0_n93, u0_n94, u0_n95, u0_n96, u0_n97, u0_n98, u0_n99, u0_r0_N70, u0_r0_N71, 
       u0_r0_N72, u0_r0_N73, u0_r0_N74, u0_r0_N75, u0_r0_N76, u0_r0_N77, u0_r0_N78, u0_r0_N79, u0_r0_N80, 
       u0_r0_N81, u0_r0_n1, u0_r0_n10, u0_r0_n11, u0_r0_n12, u0_r0_n13, u0_r0_n14, u0_r0_n15, u0_r0_n16, 
       u0_r0_n17, u0_r0_n18, u0_r0_n19, u0_r0_n2, u0_r0_n20, u0_r0_n21, u0_r0_n22, u0_r0_n23, u0_r0_n24, 
       u0_r0_n25, u0_r0_n3, u0_r0_n4, u0_r0_n5, u0_r0_n6, u0_r0_n7, u0_r0_n8, u0_r0_n9, u0_r0_rcnt_0, 
       u0_r0_rcnt_1, u0_r0_rcnt_2, u0_rcon_24, u0_rcon_25, u0_rcon_26, u0_rcon_27, u0_rcon_28, u0_rcon_29, u0_rcon_30, 
       u0_rcon_31, u0_subword_24, u0_subword_25, u0_subword_26, u0_subword_27, u0_subword_28, u0_subword_29, u0_subword_30, u0_subword_31, 
       u0_u0_n1, u0_u0_n171, u0_u0_n22, u0_u0_n438, u0_u0_n439, u0_u0_n440, u0_u0_n441, u0_u0_n442, u0_u0_n443, 
       u0_u0_n444, u0_u0_n445, u0_u0_n446, u0_u0_n447, u0_u0_n448, u0_u0_n449, u0_u0_n450, u0_u0_n451, u0_u0_n452, 
       u0_u0_n453, u0_u0_n454, u0_u0_n455, u0_u0_n456, u0_u0_n457, u0_u0_n458, u0_u0_n459, u0_u0_n460, u0_u0_n461, 
       u0_u0_n462, u0_u0_n463, u0_u0_n464, u0_u0_n465, u0_u0_n466, u0_u0_n467, u0_u0_n468, u0_u0_n469, u0_u0_n470, 
       u0_u0_n471, u0_u0_n472, u0_u0_n473, u0_u0_n474, u0_u0_n475, u0_u0_n476, u0_u0_n477, u0_u0_n478, u0_u0_n479, 
       u0_u0_n480, u0_u0_n481, u0_u0_n482, u0_u0_n483, u0_u0_n484, u0_u0_n485, u0_u0_n486, u0_u0_n487, u0_u0_n488, 
       u0_u0_n489, u0_u0_n490, u0_u0_n491, u0_u0_n492, u0_u0_n493, u0_u0_n494, u0_u0_n495, u0_u0_n496, u0_u0_n497, 
       u0_u0_n498, u0_u0_n499, u0_u0_n500, u0_u0_n501, u0_u0_n502, u0_u0_n503, u0_u0_n504, u0_u0_n505, u0_u0_n506, 
       u0_u0_n507, u0_u0_n508, u0_u0_n509, u0_u0_n510, u0_u0_n511, u0_u0_n512, u0_u0_n513, u0_u0_n514, u0_u0_n515, 
       u0_u0_n516, u0_u0_n517, u0_u0_n518, u0_u0_n519, u0_u0_n520, u0_u0_n521, u0_u0_n522, u0_u0_n523, u0_u0_n524, 
       u0_u0_n525, u0_u0_n526, u0_u0_n527, u0_u0_n528, u0_u0_n529, u0_u0_n530, u0_u0_n531, u0_u0_n532, u0_u0_n533, 
       u0_u0_n534, u0_u0_n535, u0_u0_n536, u0_u0_n537, u0_u0_n538, u0_u0_n539, u0_u0_n540, u0_u0_n541, u0_u0_n542, 
       u0_u0_n543, u0_u0_n544, u0_u0_n545, u0_u0_n546, u0_u0_n547, u0_u0_n548, u0_u0_n549, u0_u0_n550, u0_u0_n551, 
       u0_u0_n552, u0_u0_n553, u0_u0_n554, u0_u0_n555, u0_u0_n556, u0_u0_n557, u0_u0_n558, u0_u0_n559, u0_u0_n560, 
       u0_u0_n561, u0_u0_n562, u0_u0_n563, u0_u0_n564, u0_u0_n565, u0_u0_n566, u0_u0_n567, u0_u0_n568, u0_u0_n569, 
       u0_u0_n570, u0_u0_n571, u0_u0_n572, u0_u0_n573, u0_u0_n574, u0_u0_n575, u0_u0_n576, u0_u0_n577, u0_u0_n578, 
       u0_u0_n579, u0_u0_n580, u0_u0_n581, u0_u0_n582, u0_u0_n583, u0_u0_n584, u0_u0_n585, u0_u0_n586, u0_u0_n587, 
       u0_u0_n588, u0_u0_n589, u0_u0_n590, u0_u0_n591, u0_u0_n592, u0_u0_n593, u0_u0_n594, u0_u0_n595, u0_u0_n596, 
       u0_u0_n597, u0_u0_n598, u0_u0_n599, u0_u0_n600, u0_u0_n601, u0_u0_n602, u0_u0_n603, u0_u0_n604, u0_u0_n605, 
       u0_u0_n606, u0_u0_n607, u0_u0_n608, u0_u0_n609, u0_u0_n610, u0_u0_n611, u0_u0_n612, u0_u0_n613, u0_u0_n614, 
       u0_u0_n615, u0_u0_n616, u0_u0_n617, u0_u0_n618, u0_u0_n619, u0_u0_n620, u0_u0_n621, u0_u0_n622, u0_u0_n623, 
       u0_u0_n624, u0_u0_n625, u0_u0_n626, u0_u0_n627, u0_u0_n628, u0_u0_n629, u0_u0_n630, u0_u0_n631, u0_u0_n632, 
       u0_u0_n633, u0_u0_n634, u0_u0_n635, u0_u0_n636, u0_u0_n637, u0_u0_n638, u0_u0_n639, u0_u0_n640, u0_u0_n641, 
       u0_u0_n642, u0_u0_n643, u0_u0_n644, u0_u0_n645, u0_u0_n646, u0_u0_n647, u0_u0_n648, u0_u0_n649, u0_u0_n650, 
       u0_u0_n651, u0_u0_n652, u0_u0_n653, u0_u0_n654, u0_u0_n655, u0_u0_n656, u0_u0_n657, u0_u0_n658, u0_u0_n659, 
       u0_u0_n660, u0_u0_n661, u0_u0_n662, u0_u0_n663, u0_u0_n664, u0_u0_n665, u0_u0_n666, u0_u0_n667, u0_u0_n668, 
       u0_u0_n669, u0_u0_n670, u0_u0_n671, u0_u0_n672, u0_u0_n673, u0_u0_n674, u0_u0_n675, u0_u0_n676, u0_u0_n677, 
       u0_u0_n678, u0_u0_n679, u0_u0_n680, u0_u0_n681, u0_u0_n682, u0_u0_n683, u0_u0_n684, u0_u0_n685, u0_u0_n686, 
       u0_u0_n687, u0_u0_n688, u0_u0_n689, u0_u0_n690, u0_u0_n691, u0_u0_n692, u0_u0_n693, u0_u0_n694, u0_u0_n695, 
       u0_u0_n696, u0_u0_n697, u0_u0_n698, u0_u0_n699, u0_u0_n700, u0_u0_n701, u0_u0_n702, u0_u0_n703, u0_u0_n704, 
       u0_u0_n705, u0_u0_n706, u0_u0_n707, u0_u0_n708, u0_u0_n709, u0_u0_n710, u0_u0_n711, u0_u0_n712, u0_u0_n713, 
       u0_u0_n714, u0_u0_n715, u0_u0_n716, u0_u0_n717, u0_u0_n718, u0_u0_n719, u0_u0_n720, u0_u0_n721, u0_u0_n722, 
       u0_u0_n723, u0_u0_n724, u0_u0_n725, u0_u0_n726, u0_u0_n727, u0_u0_n728, u0_u0_n729, u0_u0_n730, u0_u0_n731, 
       u0_u0_n732, u0_u0_n733, u0_u0_n734, u0_u0_n735, u0_u0_n736, u0_u0_n737, u0_u0_n738, u0_u0_n739, u0_u0_n740, 
       u0_u0_n741, u0_u0_n742, u0_u0_n743, u0_u0_n744, u0_u0_n745, u0_u0_n746, u0_u0_n747, u0_u0_n748, u0_u0_n749, 
       u0_u0_n750, u0_u0_n751, u0_u0_n752, u0_u0_n753, u0_u0_n754, u0_u0_n755, u0_u0_n756, u0_u0_n757, u0_u0_n758, 
       u0_u0_n759, u0_u0_n760, u0_u0_n761, u0_u0_n762, u0_u0_n763, u0_u0_n764, u0_u0_n765, u0_u0_n766, u0_u0_n767, 
       u0_u0_n768, u0_u0_n769, u0_u0_n770, u0_u0_n771, u0_u0_n772, u0_u0_n773, u0_u0_n774, u0_u0_n775, u0_u0_n776, 
       u0_u0_n777, u0_u0_n778, u0_u0_n779, u0_u0_n780, u0_u0_n781, u0_u0_n782, u0_u0_n783, u0_u0_n784, u0_u0_n785, 
       u0_u0_n786, u0_u0_n787, u0_u0_n788, u0_u0_n789, u0_u0_n790, u0_u0_n791, u0_u0_n792, u0_u0_n793, u0_u0_n794, 
       u0_u0_n795, u0_u0_n796, u0_u0_n797, u0_u0_n798, u0_u0_n799, u0_u0_n800, u0_u0_n801, u0_u0_n802, u0_u0_n803, 
       u0_u0_n804, u0_u0_n805, u0_u0_n806, u0_u0_n807, u0_u0_n808, u0_u0_n809, u0_u0_n810, u0_u0_n811, u0_u0_n812, 
       u0_u0_n813, u0_u0_n814, u0_u0_n815, u0_u0_n816, u0_u0_n817, u0_u0_n818, u0_u0_n819, u0_u0_n820, u0_u0_n821, 
       u0_u0_n822, u0_u0_n823, u0_u0_n824, u0_u0_n825, u0_u0_n826, u0_u0_n827, u0_u0_n828, u0_u0_n829, u0_u0_n830, 
       u0_u0_n831, u0_u0_n832, u0_u0_n833, u0_u0_n834, u0_u0_n835, u0_u0_n836, u0_u0_n837, u0_u0_n838, u0_u0_n839, 
       u0_u0_n840, u0_u0_n841, u0_u0_n842, u0_u0_n843, u0_u0_n844, u0_u0_n845, u0_u0_n846, u0_u0_n847, u0_u0_n848, 
       u0_u0_n849, u0_u0_n850, u0_u0_n851, u0_u0_n852, u0_u0_n853, u0_u0_n854, u0_u0_n855, u0_u0_n856, u0_u0_n857, 
       u0_u0_n858, u0_u0_n859, u0_u0_n860, u0_u0_n861, u0_u0_n862, u0_u0_n863, u0_u0_n864, u0_u0_n865, u0_u0_n866, 
       u0_u0_n867, u0_u0_n868, u0_u0_n869, u0_u0_n870, u0_u0_n871, u0_u0_n872, u0_u0_n873, u0_u0_n874, u0_u0_n875, 
       u0_u0_n876, u0_u0_n877, u0_u0_n878, u0_u0_n879, us22_n438, us22_n439, us22_n440, us22_n441, us22_n442, 
       us22_n443, us22_n444, us22_n445, us22_n446, us22_n447, us22_n448, us22_n449, us22_n450, us22_n451, 
       us22_n452, us22_n453, us22_n454, us22_n455, us22_n456, us22_n457, us22_n458, us22_n459, us22_n460, 
       us22_n461, us22_n462, us22_n463, us22_n464, us22_n465, us22_n466, us22_n467, us22_n468, us22_n469, 
       us22_n470, us22_n471, us22_n472, us22_n473, us22_n474, us22_n475, us22_n476, us22_n477, us22_n478, 
       us22_n479, us22_n480, us22_n481, us22_n482, us22_n483, us22_n484, us22_n485, us22_n486, us22_n487, 
       us22_n488, us22_n489, us22_n490, us22_n491, us22_n492, us22_n493, us22_n494, us22_n495, us22_n496, 
       us22_n497, us22_n498, us22_n499, us22_n500, us22_n501, us22_n502, us22_n503, us22_n504, us22_n505, 
       us22_n506, us22_n507, us22_n508, us22_n509, us22_n510, us22_n511, us22_n512, us22_n513, us22_n514, 
       us22_n515, us22_n516, us22_n517, us22_n518, us22_n519, us22_n520, us22_n521, us22_n522, us22_n523, 
       us22_n524, us22_n525, us22_n526, us22_n527, us22_n528, us22_n529, us22_n530, us22_n531, us22_n532, 
       us22_n533, us22_n534, us22_n535, us22_n536, us22_n537, us22_n538, us22_n539, us22_n540, us22_n541, 
       us22_n542, us22_n543, us22_n544, us22_n545, us22_n546, us22_n547, us22_n548, us22_n549, us22_n550, 
       us22_n551, us22_n552, us22_n553, us22_n554, us22_n555, us22_n556, us22_n557, us22_n558, us22_n559, 
       us22_n560, us22_n561, us22_n562, us22_n563, us22_n564, us22_n565, us22_n566, us22_n567, us22_n568, 
       us22_n569, us22_n570, us22_n571, us22_n572, us22_n573, us22_n574, us22_n575, us22_n576, us22_n577, 
       us22_n578, us22_n579, us22_n580, us22_n581, us22_n582, us22_n583, us22_n584, us22_n585, us22_n586, 
       us22_n587, us22_n588, us22_n589, us22_n590, us22_n591, us22_n592, us22_n593, us22_n594, us22_n595, 
       us22_n596, us22_n597, us22_n598, us22_n599, us22_n600, us22_n601, us22_n602, us22_n603, us22_n604, 
       us22_n605, us22_n606, us22_n607, us22_n608, us22_n609, us22_n610, us22_n611, us22_n612, us22_n613, 
       us22_n614, us22_n615, us22_n616, us22_n617, us22_n618, us22_n619, us22_n620, us22_n621, us22_n622, 
       us22_n623, us22_n624, us22_n625, us22_n626, us22_n627, us22_n628, us22_n629, us22_n630, us22_n631, 
       us22_n632, us22_n633, us22_n634, us22_n635, us22_n636, us22_n637, us22_n638, us22_n639, us22_n640, 
       us22_n641, us22_n642, us22_n643, us22_n644, us22_n645, us22_n646, us22_n647, us22_n648, us22_n649, 
       us22_n650, us22_n651, us22_n652, us22_n653, us22_n654, us22_n655, us22_n656, us22_n657, us22_n658, 
       us22_n659, us22_n660, us22_n661, us22_n662, us22_n663, us22_n664, us22_n665, us22_n666, us22_n667, 
       us22_n668, us22_n669, us22_n670, us22_n671, us22_n672, us22_n673, us22_n674, us22_n675, us22_n676, 
       us22_n677, us22_n678, us22_n679, us22_n680, us22_n681, us22_n682, us22_n683, us22_n684, us22_n685, 
       us22_n686, us22_n687, us22_n688, us22_n689, us22_n690, us22_n691, us22_n692, us22_n693, us22_n694, 
       us22_n695, us22_n696, us22_n697, us22_n698, us22_n699, us22_n700, us22_n701, us22_n702, us22_n703, 
       us22_n704, us22_n705, us22_n706, us22_n707, us22_n708, us22_n709, us22_n710, us22_n711, us22_n712, 
       us22_n713, us22_n714, us22_n715, us22_n716, us22_n717, us22_n718, us22_n719, us22_n720, us22_n721, 
       us22_n722, us22_n723, us22_n724, us22_n725, us22_n726, us22_n727, us22_n728, us22_n729, us22_n730, 
       us22_n731, us22_n732, us22_n733, us22_n734, us22_n735, us22_n736, us22_n737, us22_n738, us22_n739, 
       us22_n740, us22_n741, us22_n742, us22_n743, us22_n744, us22_n745, us22_n746, us22_n747, us22_n748, 
       us22_n749, us22_n750, us22_n751, us22_n752, us22_n753, us22_n754, us22_n755, us22_n756, us22_n757, 
       us22_n758, us22_n759, us22_n760, us22_n761, us22_n762, us22_n763, us22_n764, us22_n765, us22_n766, 
       us22_n767, us22_n768, us22_n769, us22_n770, us22_n771, us22_n772, us22_n773, us22_n774, us22_n775, 
       us22_n776, us22_n777, us22_n778, us22_n779, us22_n780, us22_n781, us22_n782, us22_n783, us22_n784, 
       us22_n785, us22_n786, us22_n787, us22_n788, us22_n789, us22_n790, us22_n791, us22_n792, us22_n793, 
       us22_n794, us22_n795, us22_n796, us22_n797, us22_n798, us22_n799, us22_n800, us22_n801, us22_n802, 
       us22_n803, us22_n804, us22_n805, us22_n806, us22_n807, us22_n808, us22_n809, us22_n810, us22_n811, 
       us22_n812, us22_n813, us22_n814, us22_n815, us22_n816, us22_n817, us22_n818, us22_n819, us22_n820, 
       us22_n821, us22_n822, us22_n823, us22_n824, us22_n825, us22_n826, us22_n827, us22_n828, us22_n829, 
       us22_n830, us22_n831, us22_n832, us22_n833, us22_n834, us22_n835, us22_n836, us22_n837, us22_n838, 
       us22_n839, us22_n840, us22_n841, us22_n842, us22_n843, us22_n844, us22_n845, us22_n846, us22_n847, 
       us22_n848, us22_n849, us22_n850, us22_n851, us22_n852, us22_n853, us22_n854, us22_n855, us22_n856, 
       us22_n857, us22_n858, us22_n859, us22_n860, us22_n861, us22_n862, us22_n863, us22_n864, us22_n865, 
       us22_n866, us22_n867, us22_n868, us22_n869, us22_n870, us22_n871, us22_n872, us22_n873, us22_n874, 
       w0_0, w0_1, w0_10, w0_11, w0_12, w0_13, w0_14, w0_15, w0_16, 
       w0_17, w0_18, w0_19, w0_2, w0_20, w0_21, w0_22, w0_23, w0_24, 
       w0_25, w0_26, w0_27, w0_28, w0_29, w0_3, w0_30, w0_31, w0_4, 
       w0_5, w0_6, w0_7, w0_8, w0_9, w1_0, w1_1, w1_10, w1_11, 
       w1_12, w1_13, w1_14, w1_15, w1_16, w1_17, w1_18, w1_19, w1_2, 
       w1_20, w1_21, w1_22, w1_23, w1_24, w1_25, w1_26, w1_27, w1_28, 
       w1_29, w1_3, w1_30, w1_31, w1_4, w1_5, w1_6, w1_7, w1_8, 
       w1_9, w2_0, w2_1, w2_10, w2_11, w2_12, w2_13, w2_14, w2_15, 
       w2_16, w2_17, w2_18, w2_19, w2_2, w2_20, w2_21, w2_22, w2_23, 
       w2_24, w2_25, w2_26, w2_27, w2_28, w2_29, w2_3, w2_30, w2_31, 
       w2_4, w2_5, w2_6, w2_7, w2_8, w2_9, w3_12, w3_13, w3_14, 
       w3_15, w3_16, w3_17, w3_18, w3_19, w3_20, w3_21, w3_22,  w3_23;
  NAND2_X1 U10 (.A2( ld ) , .ZN( n8 ) , .A1( text_in[3] ) );
  NAND2_X1 U100 (.A2( ld ) , .ZN( n98 ) , .A1( text_in[48] ) );
  XOR2_X1 U1001 (.Z( n728 ) , .B( n729 ) , .A( sa11_sr_0 ) );
  XOR2_X1 U1002 (.Z( n729 ) , .B( sa21_sr_0 ) , .A( w1_17 ) );
  XNOR2_X1 U1004 (.B( n683 ) , .ZN( n730 ) , .A( sa01_sr_1 ) );
  XOR2_X1 U1005 (.A( n163 ) , .Z( n725 ) , .B( w1_17 ) );
  OAI22_X1 U1007 (.ZN( N194 ) , .A1( n1214 ) , .B2( n1221 ) , .A2( n731 ) , .B1( n732 ) );
  XOR2_X1 U1009 (.A( n690 ) , .B( n713 ) , .Z( n734 ) );
  OAI21_X1 U101 (.B1( ld ) , .A( n100 ) , .ZN( n1027 ) , .B2( n99 ) );
  XOR2_X1 U1010 (.Z( n713 ) , .A( sa11_sr_7 ) , .B( sa21_sr_7 ) );
  XOR2_X1 U1012 (.A( n161 ) , .Z( n731 ) , .B( w1_16 ) );
  OAI22_X1 U1014 (.ZN( N185 ) , .A1( n1214 ) , .B2( n1220 ) , .A2( n735 ) , .B1( n736 ) );
  XOR2_X1 U1016 (.A( n650 ) , .B( n665 ) , .Z( n738 ) );
  XOR2_X1 U1017 (.Z( n650 ) , .A( sa21_sr_6 ) , .B( sa31_sr_6 ) );
  XOR2_X1 U1019 (.A( n159 ) , .Z( n735 ) , .B( w1_15 ) );
  NAND2_X1 U102 (.A2( ld ) , .ZN( n100 ) , .A1( text_in[49] ) );
  OAI22_X1 U1021 (.ZN( N184 ) , .A1( n1214 ) , .B2( n1220 ) , .A2( n739 ) , .B1( n740 ) );
  XOR2_X1 U1023 (.A( n644 ) , .B( n656 ) , .Z( n742 ) );
  XOR2_X1 U1024 (.Z( n656 ) , .A( sa21_sr_5 ) , .B( sa31_sr_5 ) );
  XOR2_X1 U1026 (.A( n157 ) , .Z( n739 ) , .B( w1_14 ) );
  OAI22_X1 U1028 (.ZN( N183 ) , .A1( n1109 ) , .B2( n1221 ) , .A2( n743 ) , .B1( n744 ) );
  XOR2_X1 U1029 (.Z( n744 ) , .A( n745 ) , .B( n746 ) );
  OAI21_X1 U103 (.B1( ld ) , .B2( n101 ) , .A( n102 ) , .ZN( n1028 ) );
  XOR2_X1 U1030 (.A( n651 ) , .B( n663 ) , .Z( n746 ) );
  XOR2_X1 U1031 (.Z( n663 ) , .A( sa21_sr_4 ) , .B( sa31_sr_4 ) );
  XNOR2_X1 U1032 (.ZN( n745 ) , .B( sa31_sr_5 ) , .A( w1_13 ) );
  XOR2_X1 U1033 (.A( n155 ) , .Z( n743 ) , .B( w1_13 ) );
  OAI22_X1 U1035 (.ZN( N182 ) , .A1( n1213 ) , .B2( n1221 ) , .A2( n747 ) , .B1( n748 ) );
  XOR2_X1 U1036 (.Z( n748 ) , .A( n749 ) , .B( n750 ) );
  XOR2_X1 U1037 (.A( n657 ) , .B( n670 ) , .Z( n750 ) );
  XOR2_X1 U1038 (.Z( n670 ) , .A( sa21_sr_3 ) , .B( sa31_sr_3 ) );
  XOR2_X1 U1039 (.B( n643 ) , .Z( n749 ) , .A( n751 ) );
  NAND2_X1 U104 (.A2( ld ) , .ZN( n102 ) , .A1( text_in[50] ) );
  XNOR2_X1 U1040 (.ZN( n751 ) , .B( sa31_sr_4 ) , .A( w1_12 ) );
  XOR2_X1 U1041 (.A( n153 ) , .Z( n747 ) , .B( w1_12 ) );
  OAI22_X1 U1043 (.ZN( N181 ) , .A1( n1214 ) , .B2( n1220 ) , .A2( n752 ) , .B1( n753 ) );
  XOR2_X1 U1045 (.A( n662 ) , .B( n677 ) , .Z( n755 ) );
  XOR2_X1 U1046 (.Z( n677 ) , .A( sa21_sr_2 ) , .B( sa31_sr_2 ) );
  XNOR2_X1 U1048 (.ZN( n756 ) , .B( sa31_sr_3 ) , .A( w1_11 ) );
  XOR2_X1 U1049 (.A( n151 ) , .Z( n752 ) , .B( w1_11 ) );
  OAI21_X1 U105 (.B1( ld ) , .ZN( n1029 ) , .B2( n103 ) , .A( n104 ) );
  OAI22_X1 U1051 (.ZN( N180 ) , .A1( n1109 ) , .B2( n1217 ) , .A2( n757 ) , .B1( n758 ) );
  XOR2_X1 U1053 (.A( n671 ) , .B( n683 ) , .Z( n760 ) );
  XOR2_X1 U1054 (.Z( n683 ) , .A( sa21_sr_1 ) , .B( sa31_sr_1 ) );
  XOR2_X1 U1056 (.A( n149 ) , .Z( n757 ) , .B( w1_10 ) );
  OAI22_X1 U1058 (.ZN( N179 ) , .A1( n1214 ) , .B2( n1220 ) , .A2( n761 ) , .B1( n762 ) );
  NAND2_X1 U106 (.A2( ld ) , .ZN( n104 ) , .A1( text_in[51] ) );
  XOR2_X1 U1060 (.A( n678 ) , .B( n690 ) , .Z( n764 ) );
  XOR2_X1 U1061 (.Z( n690 ) , .A( sa21_sr_0 ) , .B( sa31_sr_0 ) );
  XNOR2_X1 U1063 (.ZN( n765 ) , .B( sa31_sr_1 ) , .A( w1_9 ) );
  XOR2_X1 U1064 (.A( n147 ) , .Z( n761 ) , .B( w1_9 ) );
  OAI22_X1 U1066 (.ZN( N178 ) , .A1( n1214 ) , .B2( n1218 ) , .A2( n766 ) , .B1( n767 ) );
  XOR2_X1 U1068 (.A( n643 ) , .B( n684 ) , .Z( n769 ) );
  XOR2_X1 U1069 (.Z( n643 ) , .A( sa21_sr_7 ) , .B( sa31_sr_7 ) );
  OAI21_X1 U107 (.B1( ld ) , .ZN( n1030 ) , .B2( n105 ) , .A( n106 ) );
  XOR2_X1 U1071 (.A( n145 ) , .Z( n766 ) , .B( w1_8 ) );
  OAI22_X1 U1073 (.ZN( N169 ) , .A1( n1109 ) , .B2( n1217 ) , .A2( n770 ) , .B1( n771 ) );
  XOR2_X1 U1074 (.Z( n771 ) , .A( n772 ) , .B( n773 ) );
  XOR2_X1 U1075 (.B( n665 ) , .Z( n773 ) , .A( sa01_sr_6 ) );
  XOR2_X1 U1076 (.Z( n665 ) , .A( sa01_sr_7 ) , .B( sa11_sr_7 ) );
  XNOR2_X1 U1077 (.ZN( n772 ) , .B( n774 ) , .A( sa21_sr_7 ) );
  XOR2_X1 U1078 (.Z( n774 ) , .B( sa31_sr_6 ) , .A( w1_7 ) );
  XOR2_X1 U1079 (.A( n143 ) , .Z( n770 ) , .B( w1_7 ) );
  NAND2_X1 U108 (.A2( ld ) , .ZN( n106 ) , .A1( text_in[52] ) );
  OAI22_X1 U1081 (.ZN( N168 ) , .A1( n1213 ) , .B2( n1218 ) , .A2( n775 ) , .B1( n776 ) );
  XOR2_X1 U1082 (.Z( n776 ) , .A( n777 ) , .B( n778 ) );
  XOR2_X1 U1083 (.Z( n778 ) , .B( n779 ) , .A( sa21_sr_6 ) );
  XOR2_X1 U1084 (.Z( n779 ) , .B( sa31_sr_5 ) , .A( w1_6 ) );
  XNOR2_X1 U1085 (.B( n644 ) , .ZN( n777 ) , .A( sa01_sr_5 ) );
  XOR2_X1 U1086 (.Z( n644 ) , .A( sa01_sr_6 ) , .B( sa11_sr_6 ) );
  XOR2_X1 U1087 (.A( n141 ) , .Z( n775 ) , .B( w1_6 ) );
  OAI22_X1 U1089 (.ZN( N167 ) , .A1( n1212 ) , .B2( n1217 ) , .A2( n780 ) , .B1( n781 ) );
  OAI21_X1 U109 (.B1( ld ) , .ZN( n1031 ) , .B2( n107 ) , .A( n108 ) );
  XOR2_X1 U1090 (.Z( n781 ) , .A( n782 ) , .B( n783 ) );
  XOR2_X1 U1091 (.Z( n783 ) , .B( n784 ) , .A( sa21_sr_5 ) );
  XOR2_X1 U1092 (.Z( n784 ) , .B( sa31_sr_4 ) , .A( w1_5 ) );
  XNOR2_X1 U1093 (.B( n651 ) , .ZN( n782 ) , .A( sa01_sr_4 ) );
  XOR2_X1 U1094 (.Z( n651 ) , .A( sa01_sr_5 ) , .B( sa11_sr_5 ) );
  XOR2_X1 U1095 (.A( n139 ) , .Z( n780 ) , .B( w1_5 ) );
  OAI22_X1 U1097 (.ZN( N166 ) , .A1( n1213 ) , .B2( n1220 ) , .A2( n785 ) , .B1( n786 ) );
  XOR2_X1 U1098 (.Z( n786 ) , .A( n787 ) , .B( n788 ) );
  XOR2_X1 U1099 (.Z( n788 ) , .B( n789 ) , .A( sa21_sr_4 ) );
  OAI21_X1 U11 (.B1( ld ) , .A( n10 ) , .B2( n9 ) , .ZN( n982 ) );
  NAND2_X1 U110 (.A2( ld ) , .ZN( n108 ) , .A1( text_in[53] ) );
  XOR2_X1 U1100 (.Z( n789 ) , .B( sa31_sr_3 ) , .A( w1_4 ) );
  XOR2_X1 U1101 (.Z( n787 ) , .A( n790 ) , .B( n791 ) );
  XNOR2_X1 U1102 (.B( n657 ) , .ZN( n790 ) , .A( sa01_sr_3 ) );
  XOR2_X1 U1103 (.Z( n657 ) , .A( sa01_sr_4 ) , .B( sa11_sr_4 ) );
  XOR2_X1 U1104 (.A( n137 ) , .Z( n785 ) , .B( w1_4 ) );
  OAI22_X1 U1106 (.ZN( N165 ) , .A1( n1216 ) , .B2( n1217 ) , .A2( n792 ) , .B1( n793 ) );
  XOR2_X1 U1109 (.Z( n796 ) , .B( sa31_sr_2 ) , .A( w1_3 ) );
  OAI21_X1 U111 (.B1( ld ) , .ZN( n1032 ) , .B2( n109 ) , .A( n110 ) );
  XOR2_X1 U1110 (.B( n791 ) , .Z( n794 ) , .A( n797 ) );
  XNOR2_X1 U1111 (.B( n662 ) , .ZN( n797 ) , .A( sa01_sr_2 ) );
  XOR2_X1 U1112 (.Z( n662 ) , .A( sa01_sr_3 ) , .B( sa11_sr_3 ) );
  XOR2_X1 U1113 (.A( n135 ) , .Z( n792 ) , .B( w1_3 ) );
  OAI22_X1 U1115 (.ZN( N164 ) , .A1( n1213 ) , .B2( n1218 ) , .A2( n798 ) , .B1( n799 ) );
  XOR2_X1 U1116 (.Z( n799 ) , .A( n800 ) , .B( n801 ) );
  XOR2_X1 U1117 (.Z( n801 ) , .B( n802 ) , .A( sa21_sr_2 ) );
  XOR2_X1 U1118 (.Z( n802 ) , .B( sa31_sr_1 ) , .A( w1_2 ) );
  XNOR2_X1 U1119 (.B( n671 ) , .ZN( n800 ) , .A( sa01_sr_1 ) );
  NAND2_X1 U112 (.A2( ld ) , .ZN( n110 ) , .A1( text_in[54] ) );
  XOR2_X1 U1120 (.Z( n671 ) , .A( sa01_sr_2 ) , .B( sa11_sr_2 ) );
  XOR2_X1 U1121 (.A( n133 ) , .Z( n798 ) , .B( w1_2 ) );
  OAI22_X1 U1123 (.ZN( N163 ) , .A1( n1215 ) , .B2( n1220 ) , .A2( n803 ) , .B1( n804 ) );
  XOR2_X1 U1125 (.Z( n806 ) , .B( n807 ) , .A( sa21_sr_1 ) );
  XOR2_X1 U1126 (.Z( n807 ) , .B( sa31_sr_0 ) , .A( w1_1 ) );
  XNOR2_X1 U1128 (.B( n678 ) , .ZN( n808 ) , .A( sa01_sr_0 ) );
  XOR2_X1 U1129 (.Z( n678 ) , .A( sa01_sr_1 ) , .B( sa11_sr_1 ) );
  OAI21_X1 U113 (.B1( ld ) , .ZN( n1033 ) , .B2( n111 ) , .A( n112 ) );
  XOR2_X1 U1130 (.A( n131 ) , .Z( n803 ) , .B( w1_1 ) );
  OAI22_X1 U1132 (.ZN( N162 ) , .A1( n1215 ) , .B2( n1217 ) , .A2( n809 ) , .B1( n810 ) );
  XOR2_X1 U1134 (.A( n684 ) , .B( n791 ) , .Z( n812 ) );
  XOR2_X1 U1135 (.Z( n791 ) , .A( sa01_sr_7 ) , .B( sa31_sr_7 ) );
  XOR2_X1 U1136 (.Z( n684 ) , .A( sa01_sr_0 ) , .B( sa11_sr_0 ) );
  XOR2_X1 U1138 (.A( n129 ) , .Z( n809 ) , .B( w1_0 ) );
  NAND2_X1 U114 (.A2( ld ) , .ZN( n112 ) , .A1( text_in[55] ) );
  OAI22_X1 U1140 (.ZN( N153 ) , .A1( n1215 ) , .B2( n1218 ) , .A2( n813 ) , .B1( n814 ) );
  XOR2_X1 U1142 (.Z( n816 ) , .A( n817 ) , .B( n818 ) );
  INV_X1 U1144 (.ZN( n819 ) , .A( sa12_sr_7 ) );
  XOR2_X1 U1145 (.A( n127 ) , .Z( n813 ) , .B( w2_31 ) );
  OAI22_X1 U1147 (.ZN( N152 ) , .A1( n1215 ) , .B2( n1217 ) , .A2( n820 ) , .B1( n821 ) );
  XOR2_X1 U1149 (.Z( n823 ) , .A( n824 ) , .B( n825 ) );
  OAI21_X1 U115 (.B1( ld ) , .ZN( n1034 ) , .B2( n113 ) , .A( n114 ) );
  XOR2_X1 U1151 (.A( n125 ) , .Z( n820 ) , .B( w2_30 ) );
  OAI22_X1 U1153 (.ZN( N151 ) , .A1( n1215 ) , .B2( n1218 ) , .A2( n826 ) , .B1( n827 ) );
  XOR2_X1 U1154 (.Z( n827 ) , .A( n828 ) , .B( n829 ) );
  XOR2_X1 U1155 (.Z( n829 ) , .A( n830 ) , .B( n831 ) );
  XNOR2_X1 U1156 (.ZN( n828 ) , .B( sa12_sr_5 ) , .A( w2_29 ) );
  XOR2_X1 U1157 (.A( n123 ) , .Z( n826 ) , .B( w2_29 ) );
  OAI22_X1 U1159 (.ZN( N150 ) , .A1( n1215 ) , .B2( n1221 ) , .A2( n832 ) , .B1( n833 ) );
  NAND2_X1 U116 (.A2( ld ) , .ZN( n114 ) , .A1( text_in[56] ) );
  XOR2_X1 U1160 (.Z( n833 ) , .A( n834 ) , .B( n835 ) );
  XOR2_X1 U1161 (.Z( n835 ) , .A( n836 ) , .B( n837 ) );
  XOR2_X1 U1162 (.Z( n834 ) , .A( n838 ) , .B( n839 ) );
  XNOR2_X1 U1163 (.ZN( n838 ) , .B( sa12_sr_4 ) , .A( w2_28 ) );
  XOR2_X1 U1164 (.A( n121 ) , .Z( n832 ) , .B( w2_28 ) );
  OAI22_X1 U1166 (.ZN( N149 ) , .A1( n1215 ) , .B2( n1221 ) , .A2( n840 ) , .B1( n841 ) );
  XOR2_X1 U1168 (.Z( n843 ) , .B( n844 ) , .A( n845 ) );
  OAI21_X1 U117 (.B1( ld ) , .ZN( n1035 ) , .B2( n115 ) , .A( n116 ) );
  XNOR2_X1 U1170 (.ZN( n846 ) , .B( sa12_sr_3 ) , .A( w2_27 ) );
  XOR2_X1 U1171 (.A( n119 ) , .Z( n840 ) , .B( w2_27 ) );
  OAI22_X1 U1173 (.ZN( N148 ) , .A1( n1215 ) , .B2( n1219 ) , .A2( n847 ) , .B1( n848 ) );
  XOR2_X1 U1175 (.A( n277 ) , .Z( n850 ) , .B( n851 ) );
  XOR2_X1 U1177 (.A( n117 ) , .Z( n847 ) , .B( w2_26 ) );
  OAI22_X1 U1179 (.ZN( N147 ) , .A1( n1215 ) , .B2( n1221 ) , .A2( n852 ) , .B1( n853 ) );
  NAND2_X1 U118 (.A2( ld ) , .ZN( n116 ) , .A1( text_in[57] ) );
  XOR2_X1 U1182 (.B( n284 ) , .Z( n854 ) , .A( n857 ) );
  XNOR2_X1 U1183 (.ZN( n857 ) , .B( sa12_sr_1 ) , .A( w2_25 ) );
  XOR2_X1 U1184 (.A( n115 ) , .Z( n852 ) , .B( w2_25 ) );
  OAI22_X1 U1186 (.ZN( N146 ) , .A1( n1215 ) , .B2( n1217 ) , .A2( n858 ) , .B1( n859 ) );
  XOR2_X1 U1188 (.A( n836 ) , .Z( n861 ) , .B( n862 ) );
  OAI21_X1 U119 (.B1( ld ) , .ZN( n1036 ) , .B2( n117 ) , .A( n118 ) );
  XOR2_X1 U1190 (.A( n113 ) , .Z( n858 ) , .B( w2_24 ) );
  OAI22_X1 U1192 (.ZN( N137 ) , .A1( n1215 ) , .B2( n1218 ) , .A2( n863 ) , .B1( n864 ) );
  XOR2_X1 U1193 (.Z( n864 ) , .A( n865 ) , .B( n866 ) );
  XOR2_X1 U1194 (.B( n817 ) , .Z( n866 ) , .A( sa02_sr_7 ) );
  XNOR2_X1 U1195 (.ZN( n865 ) , .B( n867 ) , .A( sa12_sr_6 ) );
  XOR2_X1 U1196 (.Z( n867 ) , .B( sa22_sr_6 ) , .A( w2_23 ) );
  XOR2_X1 U1197 (.A( n111 ) , .Z( n863 ) , .B( w2_23 ) );
  OAI22_X1 U1199 (.ZN( N136 ) , .A1( n1215 ) , .B2( n1219 ) , .A2( n868 ) , .B1( n869 ) );
  NAND2_X1 U12 (.A2( ld ) , .ZN( n10 ) , .A1( text_in[4] ) );
  NAND2_X1 U120 (.A2( ld ) , .ZN( n118 ) , .A1( text_in[58] ) );
  XOR2_X1 U1202 (.Z( n872 ) , .B( sa22_sr_5 ) , .A( w2_22 ) );
  XOR2_X1 U1205 (.A( n109 ) , .Z( n868 ) , .B( w2_22 ) );
  OAI22_X1 U1207 (.ZN( N135 ) , .A1( n1213 ) , .B2( n1219 ) , .A2( n874 ) , .B1( n875 ) );
  XOR2_X1 U1208 (.Z( n875 ) , .A( n876 ) , .B( n877 ) );
  XOR2_X1 U1209 (.Z( n877 ) , .B( n878 ) , .A( sa12_sr_4 ) );
  OAI21_X1 U121 (.B1( ld ) , .ZN( n1037 ) , .B2( n119 ) , .A( n120 ) );
  XOR2_X1 U1210 (.Z( n878 ) , .B( sa22_sr_4 ) , .A( w2_21 ) );
  XNOR2_X1 U1211 (.B( n831 ) , .ZN( n876 ) , .A( sa02_sr_5 ) );
  XOR2_X1 U1212 (.A( n107 ) , .Z( n874 ) , .B( w2_21 ) );
  OAI22_X1 U1214 (.ZN( N134 ) , .A1( n1212 ) , .B2( n1219 ) , .A2( n879 ) , .B1( n880 ) );
  XOR2_X1 U1215 (.Z( n880 ) , .A( n881 ) , .B( n882 ) );
  XOR2_X1 U1216 (.Z( n882 ) , .B( n883 ) , .A( sa12_sr_3 ) );
  XOR2_X1 U1217 (.Z( n883 ) , .B( sa22_sr_3 ) , .A( w2_20 ) );
  XOR2_X1 U1218 (.Z( n881 ) , .A( n884 ) , .B( n885 ) );
  XNOR2_X1 U1219 (.B( n839 ) , .ZN( n884 ) , .A( sa02_sr_4 ) );
  NAND2_X1 U122 (.A2( ld ) , .ZN( n120 ) , .A1( text_in[59] ) );
  XOR2_X1 U1220 (.A( n105 ) , .Z( n879 ) , .B( w2_20 ) );
  OAI22_X1 U1222 (.ZN( N133 ) , .A1( n1213 ) , .B2( n1219 ) , .A2( n886 ) , .B1( n887 ) );
  XOR2_X1 U1223 (.Z( n887 ) , .A( n888 ) , .B( n889 ) );
  XOR2_X1 U1224 (.Z( n889 ) , .B( n890 ) , .A( sa12_sr_2 ) );
  XOR2_X1 U1225 (.Z( n890 ) , .B( sa22_sr_2 ) , .A( w2_19 ) );
  XOR2_X1 U1228 (.A( n103 ) , .Z( n886 ) , .B( w2_19 ) );
  OAI21_X1 U123 (.B1( ld ) , .ZN( n1038 ) , .B2( n121 ) , .A( n122 ) );
  OAI22_X1 U1230 (.ZN( N132 ) , .A1( n1212 ) , .B2( n1219 ) , .A2( n892 ) , .B1( n893 ) );
  XOR2_X1 U1233 (.Z( n896 ) , .B( sa22_sr_1 ) , .A( w2_18 ) );
  XOR2_X1 U1236 (.A( n101 ) , .Z( n892 ) , .B( w2_18 ) );
  OAI22_X1 U1238 (.ZN( N131 ) , .A1( n1212 ) , .B2( n1219 ) , .A2( n898 ) , .B1( n899 ) );
  XOR2_X1 U1239 (.Z( n899 ) , .A( n900 ) , .B( n901 ) );
  NAND2_X1 U124 (.A2( ld ) , .ZN( n122 ) , .A1( text_in[60] ) );
  XOR2_X1 U1240 (.Z( n901 ) , .B( n902 ) , .A( sa12_sr_0 ) );
  XOR2_X1 U1241 (.Z( n902 ) , .B( sa22_sr_0 ) , .A( w2_17 ) );
  XOR2_X1 U1242 (.B( n885 ) , .Z( n900 ) , .A( n903 ) );
  XNOR2_X1 U1243 (.B( n856 ) , .ZN( n903 ) , .A( sa02_sr_1 ) );
  XOR2_X1 U1244 (.Z( n898 ) , .A( n99 ) , .B( w2_17 ) );
  OAI22_X1 U1246 (.ZN( N130 ) , .A1( n1213 ) , .B2( n1219 ) , .A2( n904 ) , .B1( n905 ) );
  XOR2_X1 U1248 (.A( n862 ) , .B( n885 ) , .Z( n907 ) );
  XOR2_X1 U1249 (.Z( n885 ) , .A( sa12_sr_7 ) , .B( sa22_sr_7 ) );
  OAI21_X1 U125 (.B1( ld ) , .ZN( n1039 ) , .B2( n123 ) , .A( n124 ) );
  XOR2_X1 U1251 (.Z( n904 ) , .A( n97 ) , .B( w2_16 ) );
  OAI22_X1 U1253 (.ZN( N121 ) , .A1( n1109 ) , .B2( n1219 ) , .A2( n908 ) , .B1( n909 ) );
  XOR2_X1 U1255 (.A( n824 ) , .B( n836 ) , .Z( n911 ) );
  XOR2_X1 U1256 (.Z( n824 ) , .A( sa22_sr_6 ) , .B( sa32_sr_6 ) );
  XOR2_X1 U1258 (.Z( n908 ) , .A( n95 ) , .B( w2_15 ) );
  NAND2_X1 U126 (.A2( ld ) , .ZN( n124 ) , .A1( text_in[61] ) );
  OAI22_X1 U1260 (.ZN( N120 ) , .A1( n1109 ) , .B2( n1220 ) , .A2( n912 ) , .B1( n913 ) );
  XOR2_X1 U1262 (.A( n818 ) , .B( n831 ) , .Z( n915 ) );
  XOR2_X1 U1263 (.Z( n831 ) , .A( sa22_sr_5 ) , .B( sa32_sr_5 ) );
  XOR2_X1 U1265 (.Z( n912 ) , .A( n93 ) , .B( w2_14 ) );
  OAI22_X1 U1267 (.ZN( N119 ) , .A1( n1109 ) , .B2( n1218 ) , .A2( n916 ) , .B1( n917 ) );
  XOR2_X1 U1268 (.Z( n917 ) , .A( n918 ) , .B( n919 ) );
  XOR2_X1 U1269 (.A( n825 ) , .B( n839 ) , .Z( n919 ) );
  OAI21_X1 U127 (.B1( ld ) , .ZN( n1040 ) , .B2( n125 ) , .A( n126 ) );
  XOR2_X1 U1270 (.Z( n839 ) , .A( sa22_sr_4 ) , .B( sa32_sr_4 ) );
  XNOR2_X1 U1271 (.ZN( n918 ) , .B( sa32_sr_5 ) , .A( w2_13 ) );
  XOR2_X1 U1272 (.A( n91 ) , .Z( n916 ) , .B( w2_13 ) );
  OAI22_X1 U1274 (.ZN( N118 ) , .A1( n1109 ) , .B2( n1220 ) , .A2( n920 ) , .B1( n921 ) );
  XOR2_X1 U1275 (.Z( n921 ) , .A( n922 ) , .B( n923 ) );
  XOR2_X1 U1276 (.A( n830 ) , .B( n844 ) , .Z( n923 ) );
  XOR2_X1 U1277 (.Z( n844 ) , .A( sa22_sr_3 ) , .B( sa32_sr_3 ) );
  INV_X1 U1278 (.ZN( n830 ) , .A( n924 ) );
  XOR2_X1 U1279 (.B( n817 ) , .Z( n922 ) , .A( n925 ) );
  NAND2_X1 U128 (.A2( ld ) , .ZN( n126 ) , .A1( text_in[62] ) );
  XNOR2_X1 U1280 (.ZN( n925 ) , .B( sa32_sr_4 ) , .A( w2_12 ) );
  XOR2_X1 U1281 (.A( n89 ) , .Z( n920 ) , .B( w2_12 ) );
  OAI22_X1 U1283 (.ZN( N117 ) , .A1( n1212 ) , .B2( n1220 ) , .A2( n926 ) , .B1( n927 ) );
  XOR2_X1 U1285 (.A( n837 ) , .B( n851 ) , .Z( n929 ) );
  INV_X1 U1287 (.ZN( n837 ) , .A( n930 ) );
  XNOR2_X1 U1289 (.ZN( n931 ) , .B( sa32_sr_3 ) , .A( w2_11 ) );
  OAI21_X1 U129 (.B1( ld ) , .ZN( n1041 ) , .B2( n127 ) , .A( n128 ) );
  XOR2_X1 U1290 (.A( n87 ) , .Z( n926 ) , .B( w2_11 ) );
  OAI22_X1 U1292 (.ZN( N116 ) , .A1( n1213 ) , .B2( n1217 ) , .A2( n932 ) , .B1( n933 ) );
  XOR2_X1 U1294 (.A( n845 ) , .B( n856 ) , .Z( n935 ) );
  XOR2_X1 U1295 (.Z( n856 ) , .A( sa22_sr_1 ) , .B( sa32_sr_1 ) );
  XOR2_X1 U1297 (.A( n85 ) , .Z( n932 ) , .B( w2_10 ) );
  OAI22_X1 U1299 (.ZN( N115 ) , .B2( n1114 ) , .A1( n1216 ) , .A2( n936 ) , .B1( n937 ) );
  OAI21_X1 U13 (.B1( ld ) , .B2( n11 ) , .A( n12 ) , .ZN( n983 ) );
  NAND2_X1 U130 (.A2( ld ) , .ZN( n128 ) , .A1( text_in[63] ) );
  XOR2_X1 U1301 (.A( n817 ) , .B( n862 ) , .Z( n939 ) );
  XOR2_X1 U1302 (.Z( n862 ) , .A( sa22_sr_0 ) , .B( sa32_sr_0 ) );
  XOR2_X1 U1304 (.Z( n277 ) , .A( sa02_sr_1 ) , .B( sa12_sr_1 ) );
  XNOR2_X1 U1305 (.ZN( n940 ) , .B( sa32_sr_1 ) , .A( w2_9 ) );
  XOR2_X1 U1306 (.A( n83 ) , .Z( n936 ) , .B( w2_9 ) );
  OAI22_X1 U1308 (.ZN( N114 ) , .B2( n1114 ) , .A1( n1216 ) , .A2( n941 ) , .B1( n942 ) );
  OAI21_X1 U131 (.B1( ld ) , .ZN( n1042 ) , .B2( n129 ) , .A( n130 ) );
  XOR2_X1 U1310 (.A( n284 ) , .B( n817 ) , .Z( n944 ) );
  XOR2_X1 U1311 (.Z( n817 ) , .A( sa22_sr_7 ) , .B( sa32_sr_7 ) );
  XOR2_X1 U1312 (.Z( n284 ) , .A( sa02_sr_0 ) , .B( sa12_sr_0 ) );
  XOR2_X1 U1314 (.A( n81 ) , .Z( n941 ) , .B( w2_8 ) );
  OAI22_X1 U1316 (.ZN( N105 ) , .B2( n1114 ) , .A1( n1216 ) , .A2( n945 ) , .B1( n946 ) );
  XOR2_X1 U1317 (.Z( n946 ) , .A( n947 ) , .B( n948 ) );
  XOR2_X1 U1318 (.B( n836 ) , .Z( n948 ) , .A( sa02_sr_6 ) );
  XOR2_X1 U1319 (.Z( n836 ) , .A( sa02_sr_7 ) , .B( sa12_sr_7 ) );
  NAND2_X1 U132 (.A2( ld ) , .ZN( n130 ) , .A1( text_in[64] ) );
  XNOR2_X1 U1320 (.ZN( n947 ) , .B( n949 ) , .A( sa22_sr_7 ) );
  XOR2_X1 U1321 (.Z( n949 ) , .B( sa32_sr_6 ) , .A( w2_7 ) );
  XOR2_X1 U1322 (.A( n79 ) , .Z( n945 ) , .B( w2_7 ) );
  OAI22_X1 U1324 (.ZN( N104 ) , .B2( n1114 ) , .A1( n1216 ) , .A2( n950 ) , .B1( n951 ) );
  XOR2_X1 U1327 (.Z( n954 ) , .B( sa32_sr_5 ) , .A( w2_6 ) );
  XNOR2_X1 U1328 (.B( n818 ) , .ZN( n952 ) , .A( sa02_sr_5 ) );
  XOR2_X1 U1329 (.Z( n818 ) , .A( sa02_sr_6 ) , .B( sa12_sr_6 ) );
  OAI21_X1 U133 (.B1( ld ) , .ZN( n1043 ) , .B2( n131 ) , .A( n132 ) );
  XOR2_X1 U1330 (.A( n77 ) , .Z( n950 ) , .B( w2_6 ) );
  OAI22_X1 U1332 (.ZN( N103 ) , .B2( n1114 ) , .A1( n1216 ) , .A2( n955 ) , .B1( n956 ) );
  XOR2_X1 U1333 (.Z( n956 ) , .A( n957 ) , .B( n958 ) );
  XOR2_X1 U1334 (.Z( n958 ) , .B( n959 ) , .A( sa22_sr_5 ) );
  XOR2_X1 U1335 (.Z( n959 ) , .B( sa32_sr_4 ) , .A( w2_5 ) );
  XNOR2_X1 U1336 (.B( n825 ) , .ZN( n957 ) , .A( sa02_sr_4 ) );
  XOR2_X1 U1337 (.Z( n825 ) , .A( sa02_sr_5 ) , .B( sa12_sr_5 ) );
  XOR2_X1 U1338 (.A( n75 ) , .Z( n955 ) , .B( w2_5 ) );
  NAND2_X1 U134 (.A2( ld ) , .ZN( n132 ) , .A1( text_in[65] ) );
  OAI22_X1 U1340 (.ZN( N102 ) , .B2( n1114 ) , .A1( n1216 ) , .A2( n960 ) , .B1( n961 ) );
  XOR2_X1 U1343 (.Z( n964 ) , .B( sa32_sr_3 ) , .A( w2_4 ) );
  XOR2_X1 U1344 (.A( n924 ) , .Z( n962 ) , .B( n965 ) );
  XOR2_X1 U1345 (.B( n279 ) , .Z( n965 ) , .A( sa02_sr_3 ) );
  XNOR2_X1 U1346 (.ZN( n924 ) , .A( sa02_sr_4 ) , .B( sa12_sr_4 ) );
  XOR2_X1 U1347 (.A( n73 ) , .Z( n960 ) , .B( w2_4 ) );
  OAI22_X1 U1349 (.ZN( N101 ) , .B2( n1114 ) , .A1( n1216 ) , .A2( n966 ) , .B1( n967 ) );
  OAI21_X1 U135 (.B1( ld ) , .ZN( n1044 ) , .B2( n133 ) , .A( n134 ) );
  XOR2_X1 U1351 (.Z( n969 ) , .B( n970 ) , .A( sa22_sr_3 ) );
  XOR2_X1 U1352 (.Z( n970 ) , .B( sa32_sr_2 ) , .A( w2_3 ) );
  XOR2_X1 U1354 (.B( n279 ) , .Z( n971 ) , .A( sa02_sr_2 ) );
  XOR2_X1 U1355 (.Z( n279 ) , .A( sa02_sr_7 ) , .B( sa32_sr_7 ) );
  XNOR2_X1 U1356 (.ZN( n930 ) , .A( sa02_sr_3 ) , .B( sa12_sr_3 ) );
  XOR2_X1 U1357 (.A( n71 ) , .Z( n966 ) , .B( w2_3 ) );
  OAI22_X1 U1359 (.ZN( N100 ) , .B2( n1114 ) , .A1( n1216 ) , .A2( n972 ) , .B1( n973 ) );
  NAND2_X1 U136 (.A2( ld ) , .ZN( n134 ) , .A1( text_in[66] ) );
  XOR2_X1 U1361 (.Z( n973 ) , .A( n974 ) , .B( n975 ) );
  XOR2_X1 U1362 (.Z( n975 ) , .B( n976 ) , .A( sa22_sr_2 ) );
  XOR2_X1 U1363 (.Z( n976 ) , .B( sa32_sr_1 ) , .A( w2_2 ) );
  XNOR2_X1 U1364 (.B( n845 ) , .ZN( n974 ) , .A( sa02_sr_1 ) );
  XOR2_X1 U1365 (.Z( n845 ) , .B( sa02_sr_2 ) , .A( sa12_sr_2 ) );
  XOR2_X1 U1366 (.A( n69 ) , .Z( n972 ) , .B( w2_2 ) );
  CLKBUF_X1 U1368 (.Z( n1219 ) , .A( n1220 ) );
  CLKBUF_X1 U1369 (.A( n1109 ) , .Z( n1212 ) );
  OAI21_X1 U137 (.B1( ld ) , .ZN( n1045 ) , .B2( n135 ) , .A( n136 ) );
  XOR2_X1 U1370 (.A( n1115 ) , .Z( n382 ) , .B( n384 ) );
  XOR2_X1 U1371 (.Z( n1115 ) , .B( n386 ) , .A( w3_16 ) );
  XNOR2_X1 U1372 (.B( n1116 ) , .ZN( n338 ) , .A( sa13_sr_6 ) );
  XOR2_X1 U1373 (.Z( n1116 ) , .B( sa23_sr_6 ) , .A( w3_23 ) );
  XOR2_X1 U1374 (.Z( N495 ) , .B( sa32_sr_2 ) , .A( w2_2 ) );
  XNOR2_X1 U1375 (.A( n1117 ) , .B( n885 ) , .ZN( n888 ) );
  XOR2_X1 U1376 (.Z( n1117 ) , .B( n844 ) , .A( sa02_sr_3 ) );
  XNOR2_X1 U1377 (.A( n1118 ) , .B( n539 ) , .ZN( n542 ) );
  XOR2_X1 U1378 (.Z( n1118 ) , .B( n496 ) , .A( sa00_sr_3 ) );
  XNOR2_X1 U1379 (.B( n476 ) , .ZN( n524 ) , .A( sa00_sr_6 ) );
  NAND2_X1 U138 (.A2( ld ) , .ZN( n136 ) , .A1( text_in[67] ) );
  XNOR2_X1 U1380 (.B( n824 ) , .ZN( n870 ) , .A( sa02_sr_6 ) );
  XNOR2_X1 U1381 (.B( n650 ) , .ZN( n698 ) , .A( sa01_sr_6 ) );
  XNOR2_X1 U1382 (.B( n295 ) , .ZN( n343 ) , .A( sa03_sr_6 ) );
  XNOR2_X1 U1383 (.B( n851 ) , .ZN( n894 ) , .A( sa02_sr_2 ) );
  INV_X1 U1384 (.A( n1114 ) , .ZN( n1214 ) );
  BUF_X1 U1385 (.Z( n1217 ) , .A( n1221 ) );
  BUF_X1 U1386 (.Z( n1218 ) , .A( n1221 ) );
  XNOR2_X1 U1387 (.A( n1119 ) , .ZN( n405 ) , .B( n407 ) );
  XNOR2_X1 U1388 (.ZN( n1119 ) , .B( n289 ) , .A( n408 ) );
  XNOR2_X1 U1389 (.A( n1120 ) , .ZN( n312 ) , .B( n314 ) );
  OAI21_X1 U139 (.B1( ld ) , .ZN( n1046 ) , .B2( n137 ) , .A( n138 ) );
  XNOR2_X1 U1390 (.ZN( n1120 ) , .B( n307 ) , .A( n317 ) );
  XNOR2_X1 U1391 (.A( n1121 ) , .ZN( n392 ) , .B( n394 ) );
  XOR2_X1 U1392 (.Z( n1121 ) , .B( sa33_sr_6 ) , .A( w3_14 ) );
  XNOR2_X1 U1393 (.B( n1122 ) , .ZN( n428 ) , .A( n429 ) );
  XNOR2_X1 U1394 (.ZN( n1122 ) , .B( n431 ) , .A( sa23_sr_6 ) );
  XNOR2_X1 U1395 (.A( n1123 ) , .ZN( n388 ) , .B( n390 ) );
  XOR2_X1 U1396 (.Z( n1123 ) , .B( sa33_sr_7 ) , .A( w3_15 ) );
  XNOR2_X1 U1397 (.A( n1124 ) , .ZN( n396 ) , .B( n398 ) );
  XOR2_X1 U1398 (.Z( n1124 ) , .B( sa33_sr_5 ) , .A( w3_13 ) );
  INV_X1 U1399 (.A( n1213 ) , .ZN( n1221 ) );
  NAND2_X1 U14 (.A2( ld ) , .ZN( n12 ) , .A1( text_in[5] ) );
  NAND2_X1 U140 (.A2( ld ) , .ZN( n138 ) , .A1( text_in[68] ) );
  INV_X1 U1400 (.A( n1212 ) , .ZN( n1220 ) );
  XNOR2_X1 U1401 (.A( n1125 ) , .ZN( n753 ) , .B( n755 ) );
  XNOR2_X1 U1402 (.ZN( n1125 ) , .B( n643 ) , .A( n756 ) );
  XNOR2_X1 U1403 (.A( n1126 ) , .ZN( n493 ) , .B( n495 ) );
  XNOR2_X1 U1404 (.ZN( n1126 ) , .B( n488 ) , .A( n498 ) );
  XNOR2_X1 U1405 (.A( n1127 ) , .ZN( n841 ) , .B( n843 ) );
  XNOR2_X1 U1406 (.ZN( n1127 ) , .B( n836 ) , .A( n846 ) );
  XNOR2_X1 U1407 (.A( n1128 ) , .ZN( n933 ) , .B( n935 ) );
  XOR2_X1 U1408 (.Z( n1128 ) , .B( sa32_sr_2 ) , .A( w2_10 ) );
  XNOR2_X1 U1409 (.A( n1129 ) , .ZN( n667 ) , .B( n669 ) );
  OAI21_X1 U141 (.B1( ld ) , .ZN( n1047 ) , .B2( n139 ) , .A( n140 ) );
  XNOR2_X1 U1410 (.ZN( n1129 ) , .B( n665 ) , .A( n672 ) );
  XNOR2_X1 U1411 (.A( n1130 ) , .ZN( n848 ) , .B( n850 ) );
  XOR2_X1 U1412 (.Z( n1130 ) , .B( sa12_sr_2 ) , .A( w2_26 ) );
  XNOR2_X1 U1413 (.B( n1131 ) , .ZN( n602 ) , .A( n603 ) );
  XNOR2_X1 U1414 (.ZN( n1131 ) , .B( n605 ) , .A( sa20_sr_6 ) );
  XNOR2_X1 U1415 (.A( n1132 ) , .ZN( n479 ) , .B( n481 ) );
  XOR2_X1 U1416 (.Z( n1132 ) , .B( sa10_sr_5 ) , .A( w0_29 ) );
  XNOR2_X1 U1417 (.A( n1133 ) , .ZN( n272 ) , .B( n275 ) );
  XOR2_X1 U1418 (.Z( n1133 ) , .A( n277 ) , .B( n278 ) );
  XNOR2_X1 U1419 (.B( n1134 ) , .ZN( n433 ) , .A( n434 ) );
  NAND2_X1 U142 (.A2( ld ) , .ZN( n140 ) , .A1( text_in[69] ) );
  XNOR2_X1 U1420 (.ZN( n1134 ) , .B( n436 ) , .A( sa23_sr_5 ) );
  XNOR2_X1 U1421 (.A( n1135 ) , .ZN( n579 ) , .B( n581 ) );
  XNOR2_X1 U1422 (.ZN( n1135 ) , .B( n469 ) , .A( n582 ) );
  XNOR2_X1 U1423 (.A( n1136 ) , .ZN( n814 ) , .B( n816 ) );
  XNOR2_X1 U1424 (.ZN( n1136 ) , .B( n819 ) , .A( w2_31 ) );
  XNOR2_X1 U1425 (.A( n1137 ) , .ZN( n325 ) , .B( n327 ) );
  XNOR2_X1 U1426 (.ZN( n1137 ) , .B( n307 ) , .A( n330 ) );
  XNOR2_X1 U1427 (.A( n1138 ) , .ZN( n927 ) , .B( n929 ) );
  XNOR2_X1 U1428 (.ZN( n1138 ) , .B( n817 ) , .A( n931 ) );
  XNOR2_X1 U1429 (.B( n1139 ) , .ZN( n893 ) , .A( n894 ) );
  OAI21_X1 U143 (.B1( ld ) , .ZN( n1048 ) , .B2( n141 ) , .A( n142 ) );
  XNOR2_X1 U1430 (.ZN( n1139 ) , .B( n896 ) , .A( sa12_sr_1 ) );
  XNOR2_X1 U1431 (.B( n1140 ) , .ZN( n445 ) , .A( n446 ) );
  XNOR2_X1 U1432 (.ZN( n1140 ) , .B( n448 ) , .A( sa23_sr_3 ) );
  XNOR2_X1 U1433 (.B( n1141 ) , .ZN( n362 ) , .A( n363 ) );
  XNOR2_X1 U1434 (.ZN( n1141 ) , .B( n365 ) , .A( sa13_sr_2 ) );
  XNOR2_X1 U1435 (.B( n1142 ) , .ZN( n369 ) , .A( n370 ) );
  XNOR2_X1 U1436 (.ZN( n1142 ) , .B( n372 ) , .A( sa13_sr_1 ) );
  XNOR2_X1 U1437 (.B( n1143 ) , .ZN( n715 ) , .A( n716 ) );
  XNOR2_X1 U1438 (.ZN( n1143 ) , .B( n718 ) , .A( sa11_sr_2 ) );
  XNOR2_X1 U1439 (.A( n1144 ) , .ZN( n500 ) , .B( n502 ) );
  NAND2_X1 U144 (.A2( ld ) , .ZN( n142 ) , .A1( text_in[70] ) );
  XOR2_X1 U1440 (.Z( n1144 ) , .B( sa10_sr_2 ) , .A( w0_26 ) );
  XNOR2_X1 U1441 (.A( n1145 ) , .ZN( n967 ) , .B( n969 ) );
  XNOR2_X1 U1442 (.ZN( n1145 ) , .A( n930 ) , .B( n971 ) );
  XNOR2_X1 U1443 (.A( n1146 ) , .ZN( n640 ) , .B( n642 ) );
  XNOR2_X1 U1444 (.ZN( n1146 ) , .B( n645 ) , .A( w1_31 ) );
  XNOR2_X1 U1445 (.A( n1147 ) , .ZN( n687 ) , .B( n689 ) );
  XOR2_X1 U1446 (.Z( n1147 ) , .B( sa11_sr_0 ) , .A( w1_24 ) );
  XNOR2_X1 U1447 (.A( n1148 ) , .ZN( n281 ) , .B( n283 ) );
  XOR2_X1 U1448 (.Z( n1148 ) , .B( sa22_sr_0 ) , .A( w2_0 ) );
  XNOR2_X1 U1449 (.B( n1149 ) , .ZN( n619 ) , .A( n620 ) );
  OAI21_X1 U145 (.B1( ld ) , .ZN( n1049 ) , .B2( n143 ) , .A( n144 ) );
  XNOR2_X1 U1450 (.ZN( n1149 ) , .B( n622 ) , .A( sa20_sr_3 ) );
  XNOR2_X1 U1451 (.A( n1150 ) , .ZN( n937 ) , .B( n939 ) );
  XNOR2_X1 U1452 (.ZN( n1150 ) , .B( n277 ) , .A( n940 ) );
  XNOR2_X1 U1453 (.A( n1151 ) , .ZN( n859 ) , .B( n861 ) );
  XOR2_X1 U1454 (.Z( n1151 ) , .B( sa12_sr_0 ) , .A( w2_24 ) );
  XNOR2_X1 U1455 (.A( n1152 ) , .ZN( n736 ) , .B( n738 ) );
  XOR2_X1 U1456 (.Z( n1152 ) , .B( sa31_sr_7 ) , .A( w1_15 ) );
  XNOR2_X1 U1457 (.A( n1153 ) , .ZN( n562 ) , .B( n564 ) );
  XOR2_X1 U1458 (.Z( n1153 ) , .B( sa30_sr_7 ) , .A( w0_15 ) );
  XNOR2_X1 U1459 (.A( n1154 ) , .ZN( n909 ) , .B( n911 ) );
  NAND2_X1 U146 (.A2( ld ) , .ZN( n144 ) , .A1( text_in[71] ) );
  XOR2_X1 U1460 (.Z( n1154 ) , .B( sa32_sr_7 ) , .A( w2_15 ) );
  XNOR2_X1 U1461 (.A( n1155 ) , .ZN( n473 ) , .B( n475 ) );
  XOR2_X1 U1462 (.Z( n1155 ) , .B( sa10_sr_6 ) , .A( w0_30 ) );
  XNOR2_X1 U1463 (.A( n1156 ) , .ZN( n821 ) , .B( n823 ) );
  XOR2_X1 U1464 (.Z( n1156 ) , .B( sa12_sr_6 ) , .A( w2_30 ) );
  XNOR2_X1 U1465 (.A( n1157 ) , .ZN( n647 ) , .B( n649 ) );
  XOR2_X1 U1466 (.Z( n1157 ) , .B( sa11_sr_6 ) , .A( w1_30 ) );
  XNOR2_X1 U1467 (.A( n1158 ) , .ZN( n588 ) , .B( n590 ) );
  XNOR2_X1 U1468 (.ZN( n1158 ) , .B( n469 ) , .A( n591 ) );
  XNOR2_X1 U1469 (.A( n1159 ) , .ZN( n762 ) , .B( n764 ) );
  OAI21_X1 U147 (.B1( ld ) , .ZN( n1050 ) , .B2( n145 ) , .A( n146 ) );
  XNOR2_X1 U1470 (.ZN( n1159 ) , .B( n643 ) , .A( n765 ) );
  XNOR2_X1 U1471 (.B( n1160 ) , .ZN( n523 ) , .A( n524 ) );
  XNOR2_X1 U1472 (.ZN( n1160 ) , .B( n526 ) , .A( sa10_sr_5 ) );
  XNOR2_X1 U1473 (.B( n1161 ) , .ZN( n869 ) , .A( n870 ) );
  XNOR2_X1 U1474 (.ZN( n1161 ) , .B( n872 ) , .A( sa12_sr_5 ) );
  XNOR2_X1 U1475 (.B( n1162 ) , .ZN( n697 ) , .A( n698 ) );
  XNOR2_X1 U1476 (.ZN( n1162 ) , .B( n700 ) , .A( sa11_sr_5 ) );
  XNOR2_X1 U1477 (.A( n1163 ) , .ZN( n740 ) , .B( n742 ) );
  XOR2_X1 U1478 (.Z( n1163 ) , .B( sa31_sr_6 ) , .A( w1_14 ) );
  XNOR2_X1 U1479 (.A( n1164 ) , .ZN( n913 ) , .B( n915 ) );
  NAND2_X1 U148 (.A2( ld ) , .ZN( n146 ) , .A1( text_in[72] ) );
  XOR2_X1 U1480 (.Z( n1164 ) , .B( sa32_sr_6 ) , .A( w2_14 ) );
  XNOR2_X1 U1481 (.A( n1165 ) , .ZN( n414 ) , .B( n416 ) );
  XNOR2_X1 U1482 (.ZN( n1165 ) , .B( n289 ) , .A( n417 ) );
  XNOR2_X1 U1483 (.A( n1166 ) , .ZN( n506 ) , .B( n508 ) );
  XNOR2_X1 U1484 (.ZN( n1166 ) , .B( n488 ) , .A( n511 ) );
  XNOR2_X1 U1485 (.B( n1167 ) , .ZN( n793 ) , .A( n794 ) );
  XNOR2_X1 U1486 (.ZN( n1167 ) , .B( n796 ) , .A( sa21_sr_3 ) );
  XNOR2_X1 U1487 (.A( n1168 ) , .ZN( n942 ) , .B( n944 ) );
  XOR2_X1 U1488 (.Z( n1168 ) , .B( sa32_sr_0 ) , .A( w2_8 ) );
  XNOR2_X1 U1489 (.A( n1169 ) , .ZN( n566 ) , .B( n568 ) );
  OAI21_X1 U149 (.B1( ld ) , .ZN( n1051 ) , .B2( n147 ) , .A( n148 ) );
  XOR2_X1 U1490 (.Z( n1169 ) , .B( sa30_sr_6 ) , .A( w0_14 ) );
  XNOR2_X1 U1491 (.A( n1170 ) , .ZN( n767 ) , .B( n769 ) );
  XOR2_X1 U1492 (.Z( n1170 ) , .B( sa31_sr_0 ) , .A( w1_8 ) );
  XNOR2_X1 U1493 (.A( n1171 ) , .ZN( n732 ) , .B( n734 ) );
  XOR2_X1 U1494 (.Z( n1171 ) , .B( sa01_sr_0 ) , .A( w1_16 ) );
  XNOR2_X1 U1495 (.B( n1172 ) , .ZN( n853 ) , .A( n854 ) );
  XNOR2_X1 U1496 (.ZN( n1172 ) , .A( n836 ) , .B( n856 ) );
  XNOR2_X1 U1497 (.A( n1173 ) , .ZN( n905 ) , .B( n907 ) );
  XOR2_X1 U1498 (.Z( n1173 ) , .B( sa02_sr_0 ) , .A( w2_16 ) );
  XNOR2_X1 U1499 (.A( n1174 ) , .ZN( n653 ) , .B( n655 ) );
  OAI21_X1 U15 (.B1( ld ) , .B2( n13 ) , .A( n14 ) , .ZN( n984 ) );
  NAND2_X1 U150 (.A2( ld ) , .ZN( n148 ) , .A1( text_in[73] ) );
  XOR2_X1 U1500 (.Z( n1174 ) , .B( sa11_sr_5 ) , .A( w1_29 ) );
  XNOR2_X1 U1501 (.B( n1175 ) , .ZN( n456 ) , .A( n457 ) );
  XNOR2_X1 U1502 (.ZN( n1175 ) , .B( n459 ) , .A( sa23_sr_1 ) );
  XNOR2_X1 U1503 (.B( n1176 ) , .ZN( n721 ) , .A( n722 ) );
  XNOR2_X1 U1504 (.ZN( n1176 ) , .B( n724 ) , .A( sa11_sr_1 ) );
  XNOR2_X1 U1505 (.A( n1177 ) , .ZN( n680 ) , .B( n682 ) );
  XNOR2_X1 U1506 (.ZN( n1177 ) , .B( n665 ) , .A( n685 ) );
  XNOR2_X1 U1507 (.B( n1178 ) , .ZN( n625 ) , .A( n626 ) );
  XNOR2_X1 U1508 (.ZN( n1178 ) , .B( n628 ) , .A( sa20_sr_2 ) );
  XNOR2_X1 U1509 (.B( n1179 ) , .ZN( n547 ) , .A( n548 ) );
  OAI21_X1 U151 (.B1( ld ) , .ZN( n1052 ) , .B2( n149 ) , .A( n150 ) );
  XNOR2_X1 U1510 (.ZN( n1179 ) , .B( n550 ) , .A( sa10_sr_1 ) );
  XNOR2_X1 U1511 (.B( n1180 ) , .ZN( n375 ) , .A( n376 ) );
  XNOR2_X1 U1512 (.ZN( n1180 ) , .B( n378 ) , .A( sa13_sr_0 ) );
  XNOR2_X1 U1513 (.B( n1181 ) , .ZN( n961 ) , .A( n962 ) );
  XNOR2_X1 U1514 (.ZN( n1181 ) , .B( n964 ) , .A( sa22_sr_4 ) );
  XNOR2_X1 U1515 (.B( n1182 ) , .ZN( n342 ) , .A( n343 ) );
  XNOR2_X1 U1516 (.ZN( n1182 ) , .B( n345 ) , .A( sa13_sr_5 ) );
  XNOR2_X1 U1517 (.A( n1183 ) , .ZN( n552 ) , .B( n554 ) );
  XNOR2_X1 U1518 (.ZN( n1183 ) , .B( n539 ) , .A( n556 ) );
  XNOR2_X1 U1519 (.A( n1184 ) , .ZN( n810 ) , .B( n812 ) );
  NAND2_X1 U152 (.A2( ld ) , .ZN( n150 ) , .A1( text_in[74] ) );
  XOR2_X1 U1520 (.Z( n1184 ) , .B( sa21_sr_0 ) , .A( w1_0 ) );
  XNOR2_X1 U1521 (.A( n1185 ) , .ZN( n726 ) , .B( n728 ) );
  XNOR2_X1 U1522 (.ZN( n1185 ) , .B( n713 ) , .A( n730 ) );
  XNOR2_X1 U1523 (.B( n1186 ) , .ZN( n951 ) , .A( n952 ) );
  XNOR2_X1 U1524 (.ZN( n1186 ) , .B( n954 ) , .A( sa22_sr_6 ) );
  XNOR2_X1 U1525 (.A( n1187 ) , .ZN( n804 ) , .B( n806 ) );
  XNOR2_X1 U1526 (.ZN( n1187 ) , .B( n791 ) , .A( n808 ) );
  XNOR2_X1 U1527 (.A( n1188 ) , .ZN( n630 ) , .B( n632 ) );
  XNOR2_X1 U1528 (.ZN( n1188 ) , .B( n617 ) , .A( n634 ) );
  XOR2_X1 U1529 (.B( n1189 ) , .Z( n693 ) , .A( sa11_sr_6 ) );
  OAI21_X1 U153 (.B1( ld ) , .ZN( n1053 ) , .B2( n151 ) , .A( n152 ) );
  XNOR2_X1 U1530 (.ZN( n1189 ) , .B( sa21_sr_6 ) , .A( w1_23 ) );
  XNOR2_X1 U1531 (.A( n1190 ) , .ZN( n419 ) , .B( n421 ) );
  XOR2_X1 U1532 (.Z( n1190 ) , .B( sa33_sr_0 ) , .A( w3_8 ) );
  XNOR2_X1 U1533 (.A( n1191 ) , .ZN( n466 ) , .B( n468 ) );
  XNOR2_X1 U1534 (.ZN( n1191 ) , .B( n471 ) , .A( w0_31 ) );
  XNOR2_X1 U1535 (.A( n1192 ) , .ZN( n513 ) , .B( n515 ) );
  XOR2_X1 U1536 (.Z( n1192 ) , .B( sa10_sr_0 ) , .A( w0_24 ) );
  XNOR2_X1 U1537 (.A( n1193 ) , .ZN( n332 ) , .B( n334 ) );
  XOR2_X1 U1538 (.Z( n1193 ) , .B( sa13_sr_0 ) , .A( w3_24 ) );
  XNOR2_X1 U1539 (.A( n1194 ) , .ZN( n593 ) , .B( n595 ) );
  NAND2_X1 U154 (.A2( ld ) , .ZN( n152 ) , .A1( text_in[75] ) );
  XOR2_X1 U1540 (.Z( n1194 ) , .B( sa30_sr_0 ) , .A( w0_8 ) );
  XNOR2_X1 U1541 (.A( n1195 ) , .ZN( n286 ) , .B( n288 ) );
  XOR2_X1 U1542 (.Z( n1195 ) , .B( sa13_sr_7 ) , .A( w3_31 ) );
  XNOR2_X1 U1543 (.A( n1196 ) , .ZN( n584 ) , .B( n586 ) );
  XOR2_X1 U1544 (.Z( n1196 ) , .B( sa30_sr_2 ) , .A( w0_10 ) );
  XNOR2_X1 U1545 (.A( n1197 ) , .ZN( n674 ) , .B( n676 ) );
  XOR2_X1 U1546 (.Z( n1197 ) , .B( sa11_sr_2 ) , .A( w1_26 ) );
  XNOR2_X1 U1547 (.A( n1198 ) , .ZN( n758 ) , .B( n760 ) );
  XOR2_X1 U1548 (.Z( n1198 ) , .B( sa31_sr_2 ) , .A( w1_10 ) );
  XNOR2_X1 U1549 (.A( n1199 ) , .ZN( n298 ) , .B( n300 ) );
  OAI21_X1 U155 (.B1( ld ) , .ZN( n1054 ) , .B2( n153 ) , .A( n154 ) );
  XOR2_X1 U1550 (.Z( n1199 ) , .B( sa13_sr_5 ) , .A( w3_29 ) );
  XNOR2_X1 U1551 (.A( n1200 ) , .ZN( n319 ) , .B( n321 ) );
  XOR2_X1 U1552 (.Z( n1200 ) , .B( sa13_sr_2 ) , .A( w3_26 ) );
  XNOR2_X1 U1553 (.A( n1201 ) , .ZN( n410 ) , .B( n412 ) );
  XOR2_X1 U1554 (.Z( n1201 ) , .B( sa33_sr_2 ) , .A( w3_10 ) );
  XNOR2_X1 U1555 (.A( n1202 ) , .ZN( n462 ) , .B( n464 ) );
  XOR2_X1 U1556 (.Z( n1202 ) , .B( sa23_sr_0 ) , .A( w3_0 ) );
  XNOR2_X1 U1557 (.A( n1203 ) , .ZN( n558 ) , .B( n560 ) );
  XOR2_X1 U1558 (.Z( n1203 ) , .B( sa00_sr_0 ) , .A( w0_16 ) );
  XNOR2_X1 U1559 (.A( n1204 ) , .ZN( n636 ) , .B( n638 ) );
  NAND2_X1 U156 (.A2( ld ) , .ZN( n154 ) , .A1( text_in[76] ) );
  XOR2_X1 U1560 (.Z( n1204 ) , .B( sa20_sr_0 ) , .A( w0_0 ) );
  XNOR2_X1 U1561 (.A( n1205 ) , .ZN( n292 ) , .B( n294 ) );
  XOR2_X1 U1562 (.Z( n1205 ) , .B( sa13_sr_6 ) , .A( w3_30 ) );
  XNOR2_X1 U1563 (.ZN( N415 ) , .B( n1206 ) , .A( w0_18 ) );
  XNOR2_X1 U1564 (.ZN( N463 ) , .B( n1208 ) , .A( w2_10 ) );
  BUF_X1 U1565 (.A( n1109 ) , .Z( n1213 ) );
  XNOR2_X1 U1566 (.ZN( N423 ) , .B( n1207 ) , .A( w1_18 ) );
  INV_X1 U1567 (.ZN( n1206 ) , .A( sa10_sr_2 ) );
  INV_X1 U1568 (.ZN( n1207 ) , .A( sa11_sr_2 ) );
  NAND2_X1 U1569 (.A2( n1209 ) , .ZN( n1210 ) , .A1( sa22_sr_2 ) );
  OAI21_X1 U157 (.B1( ld ) , .ZN( n1055 ) , .B2( n155 ) , .A( n156 ) );
  NAND2_X1 U1570 (.A1( n1208 ) , .ZN( n1211 ) , .A2( sa32_sr_2 ) );
  NAND2_X1 U1571 (.A1( n1210 ) , .A2( n1211 ) , .ZN( n851 ) );
  INV_X1 U1572 (.ZN( n1208 ) , .A( sa22_sr_2 ) );
  INV_X1 U1573 (.ZN( n1209 ) , .A( sa32_sr_2 ) );
  INV_X1 U1574 (.ZN( n1215 ) , .A( n1221 ) );
  INV_X1 U1575 (.ZN( n1216 ) , .A( n1221 ) );
  INV_X1 U1576 (.A( ld ) , .ZN( n1222 ) );
  NAND2_X1 U158 (.A2( ld ) , .ZN( n156 ) , .A1( text_in[77] ) );
  OAI21_X1 U159 (.B1( ld ) , .ZN( n1056 ) , .B2( n157 ) , .A( n158 ) );
  NAND2_X1 U16 (.A2( ld ) , .ZN( n14 ) , .A1( text_in[6] ) );
  NAND2_X1 U160 (.A2( ld ) , .ZN( n158 ) , .A1( text_in[78] ) );
  OAI21_X1 U161 (.B1( ld ) , .ZN( n1057 ) , .B2( n159 ) , .A( n160 ) );
  NAND2_X1 U162 (.A2( ld ) , .ZN( n160 ) , .A1( text_in[79] ) );
  OAI21_X1 U163 (.B1( ld ) , .ZN( n1058 ) , .B2( n161 ) , .A( n162 ) );
  NAND2_X1 U164 (.A2( ld ) , .ZN( n162 ) , .A1( text_in[80] ) );
  OAI21_X1 U165 (.B1( ld ) , .ZN( n1059 ) , .B2( n163 ) , .A( n164 ) );
  NAND2_X1 U166 (.A2( ld ) , .ZN( n164 ) , .A1( text_in[81] ) );
  OAI21_X1 U167 (.B1( ld ) , .ZN( n1060 ) , .B2( n165 ) , .A( n166 ) );
  NAND2_X1 U168 (.A2( ld ) , .ZN( n166 ) , .A1( text_in[82] ) );
  OAI21_X1 U169 (.B1( ld ) , .ZN( n1061 ) , .B2( n167 ) , .A( n168 ) );
  OAI21_X1 U17 (.B1( ld ) , .B2( n15 ) , .A( n16 ) , .ZN( n985 ) );
  NAND2_X1 U170 (.A2( ld ) , .ZN( n168 ) , .A1( text_in[83] ) );
  OAI21_X1 U171 (.B1( ld ) , .ZN( n1062 ) , .B2( n169 ) , .A( n170 ) );
  NAND2_X1 U172 (.A2( ld ) , .ZN( n170 ) , .A1( text_in[84] ) );
  OAI21_X1 U173 (.B1( ld ) , .ZN( n1063 ) , .B2( n171 ) , .A( n172 ) );
  NAND2_X1 U174 (.A2( ld ) , .ZN( n172 ) , .A1( text_in[85] ) );
  OAI21_X1 U175 (.B1( ld ) , .ZN( n1064 ) , .B2( n173 ) , .A( n174 ) );
  NAND2_X1 U176 (.A2( ld ) , .ZN( n174 ) , .A1( text_in[86] ) );
  OAI21_X1 U177 (.B1( ld ) , .ZN( n1065 ) , .B2( n175 ) , .A( n176 ) );
  NAND2_X1 U178 (.A2( ld ) , .ZN( n176 ) , .A1( text_in[87] ) );
  OAI21_X1 U179 (.B1( ld ) , .ZN( n1066 ) , .B2( n177 ) , .A( n178 ) );
  NAND2_X1 U18 (.A2( ld ) , .ZN( n16 ) , .A1( text_in[7] ) );
  NAND2_X1 U180 (.A2( ld ) , .ZN( n178 ) , .A1( text_in[88] ) );
  OAI21_X1 U181 (.B1( ld ) , .ZN( n1067 ) , .B2( n179 ) , .A( n180 ) );
  NAND2_X1 U182 (.A2( ld ) , .ZN( n180 ) , .A1( text_in[89] ) );
  OAI21_X1 U183 (.B1( ld ) , .ZN( n1068 ) , .B2( n181 ) , .A( n182 ) );
  NAND2_X1 U184 (.A2( ld ) , .ZN( n182 ) , .A1( text_in[90] ) );
  OAI21_X1 U185 (.B1( ld ) , .ZN( n1069 ) , .B2( n183 ) , .A( n184 ) );
  NAND2_X1 U186 (.A2( ld ) , .ZN( n184 ) , .A1( text_in[91] ) );
  OAI21_X1 U187 (.B1( ld ) , .ZN( n1070 ) , .B2( n185 ) , .A( n186 ) );
  NAND2_X1 U188 (.A2( ld ) , .ZN( n186 ) , .A1( text_in[92] ) );
  OAI21_X1 U189 (.B1( ld ) , .ZN( n1071 ) , .B2( n187 ) , .A( n188 ) );
  OAI21_X1 U19 (.B1( ld ) , .B2( n17 ) , .A( n18 ) , .ZN( n986 ) );
  NAND2_X1 U190 (.A2( ld ) , .ZN( n188 ) , .A1( text_in[93] ) );
  OAI21_X1 U191 (.B1( ld ) , .ZN( n1072 ) , .B2( n189 ) , .A( n190 ) );
  NAND2_X1 U192 (.A2( ld ) , .ZN( n190 ) , .A1( text_in[94] ) );
  OAI21_X1 U193 (.B1( ld ) , .ZN( n1073 ) , .B2( n191 ) , .A( n192 ) );
  NAND2_X1 U194 (.A2( ld ) , .ZN( n192 ) , .A1( text_in[95] ) );
  OAI21_X1 U195 (.B1( ld ) , .ZN( n1074 ) , .B2( n193 ) , .A( n194 ) );
  NAND2_X1 U196 (.A2( ld ) , .ZN( n194 ) , .A1( text_in[96] ) );
  OAI21_X1 U197 (.B1( ld ) , .ZN( n1075 ) , .B2( n195 ) , .A( n196 ) );
  NAND2_X1 U198 (.A2( ld ) , .ZN( n196 ) , .A1( text_in[97] ) );
  OAI21_X1 U199 (.B1( ld ) , .ZN( n1076 ) , .B2( n197 ) , .A( n198 ) );
  NAND2_X1 U20 (.A2( ld ) , .ZN( n18 ) , .A1( text_in[8] ) );
  NAND2_X1 U200 (.A2( ld ) , .ZN( n198 ) , .A1( text_in[98] ) );
  OAI21_X1 U201 (.B1( ld ) , .ZN( n1077 ) , .B2( n199 ) , .A( n200 ) );
  NAND2_X1 U202 (.A2( ld ) , .ZN( n200 ) , .A1( text_in[99] ) );
  OAI21_X1 U203 (.B1( ld ) , .ZN( n1078 ) , .B2( n201 ) , .A( n202 ) );
  NAND2_X1 U204 (.A2( ld ) , .ZN( n202 ) , .A1( text_in[100] ) );
  OAI21_X1 U205 (.B1( ld ) , .ZN( n1079 ) , .B2( n203 ) , .A( n204 ) );
  NAND2_X1 U206 (.A2( ld ) , .ZN( n204 ) , .A1( text_in[101] ) );
  OAI21_X1 U207 (.B1( ld ) , .ZN( n1080 ) , .B2( n205 ) , .A( n206 ) );
  NAND2_X1 U208 (.A2( ld ) , .ZN( n206 ) , .A1( text_in[102] ) );
  OAI21_X1 U209 (.B1( ld ) , .ZN( n1081 ) , .B2( n207 ) , .A( n208 ) );
  OAI21_X1 U21 (.B1( ld ) , .B2( n19 ) , .A( n20 ) , .ZN( n987 ) );
  NAND2_X1 U210 (.A2( ld ) , .ZN( n208 ) , .A1( text_in[103] ) );
  OAI21_X1 U211 (.B1( ld ) , .ZN( n1082 ) , .B2( n209 ) , .A( n210 ) );
  NAND2_X1 U212 (.A2( ld ) , .ZN( n210 ) , .A1( text_in[104] ) );
  OAI21_X1 U213 (.B1( ld ) , .ZN( n1083 ) , .B2( n211 ) , .A( n212 ) );
  NAND2_X1 U214 (.A2( ld ) , .ZN( n212 ) , .A1( text_in[105] ) );
  OAI21_X1 U215 (.B1( ld ) , .ZN( n1084 ) , .B2( n213 ) , .A( n214 ) );
  NAND2_X1 U216 (.A2( ld ) , .ZN( n214 ) , .A1( text_in[106] ) );
  OAI21_X1 U217 (.B1( ld ) , .ZN( n1085 ) , .B2( n215 ) , .A( n216 ) );
  NAND2_X1 U218 (.A2( ld ) , .ZN( n216 ) , .A1( text_in[107] ) );
  OAI21_X1 U219 (.B1( ld ) , .ZN( n1086 ) , .B2( n217 ) , .A( n218 ) );
  NAND2_X1 U22 (.A2( ld ) , .ZN( n20 ) , .A1( text_in[9] ) );
  NAND2_X1 U220 (.A2( ld ) , .ZN( n218 ) , .A1( text_in[108] ) );
  OAI21_X1 U221 (.B1( ld ) , .ZN( n1087 ) , .B2( n219 ) , .A( n220 ) );
  NAND2_X1 U222 (.A2( ld ) , .ZN( n220 ) , .A1( text_in[109] ) );
  OAI21_X1 U223 (.B1( ld ) , .ZN( n1088 ) , .B2( n221 ) , .A( n222 ) );
  NAND2_X1 U224 (.A2( ld ) , .ZN( n222 ) , .A1( text_in[110] ) );
  OAI21_X1 U225 (.B1( ld ) , .ZN( n1089 ) , .B2( n223 ) , .A( n224 ) );
  NAND2_X1 U226 (.A2( ld ) , .ZN( n224 ) , .A1( text_in[111] ) );
  OAI21_X1 U227 (.B1( ld ) , .ZN( n1090 ) , .B2( n225 ) , .A( n226 ) );
  NAND2_X1 U228 (.A2( ld ) , .ZN( n226 ) , .A1( text_in[112] ) );
  OAI21_X1 U229 (.B1( ld ) , .ZN( n1091 ) , .B2( n227 ) , .A( n228 ) );
  OAI21_X1 U23 (.B1( ld ) , .B2( n21 ) , .A( n22 ) , .ZN( n988 ) );
  NAND2_X1 U230 (.A2( ld ) , .ZN( n228 ) , .A1( text_in[113] ) );
  OAI21_X1 U231 (.B1( ld ) , .ZN( n1092 ) , .B2( n229 ) , .A( n230 ) );
  NAND2_X1 U232 (.A2( ld ) , .ZN( n230 ) , .A1( text_in[114] ) );
  OAI21_X1 U233 (.B1( ld ) , .ZN( n1093 ) , .B2( n231 ) , .A( n232 ) );
  NAND2_X1 U234 (.A2( ld ) , .ZN( n232 ) , .A1( text_in[115] ) );
  OAI21_X1 U235 (.B1( ld ) , .ZN( n1094 ) , .B2( n233 ) , .A( n234 ) );
  NAND2_X1 U236 (.A2( ld ) , .ZN( n234 ) , .A1( text_in[116] ) );
  OAI21_X1 U237 (.B1( ld ) , .ZN( n1095 ) , .B2( n235 ) , .A( n236 ) );
  NAND2_X1 U238 (.A2( ld ) , .ZN( n236 ) , .A1( text_in[117] ) );
  OAI21_X1 U239 (.B1( ld ) , .ZN( n1096 ) , .B2( n237 ) , .A( n238 ) );
  NAND2_X1 U24 (.A2( ld ) , .ZN( n22 ) , .A1( text_in[10] ) );
  NAND2_X1 U240 (.A2( ld ) , .ZN( n238 ) , .A1( text_in[118] ) );
  OAI21_X1 U241 (.B1( ld ) , .ZN( n1097 ) , .B2( n239 ) , .A( n240 ) );
  NAND2_X1 U242 (.A2( ld ) , .ZN( n240 ) , .A1( text_in[119] ) );
  OAI21_X1 U243 (.B1( ld ) , .ZN( n1098 ) , .B2( n241 ) , .A( n242 ) );
  NAND2_X1 U244 (.A2( ld ) , .ZN( n242 ) , .A1( text_in[120] ) );
  OAI21_X1 U245 (.B1( ld ) , .ZN( n1099 ) , .B2( n243 ) , .A( n244 ) );
  NAND2_X1 U246 (.A2( ld ) , .ZN( n244 ) , .A1( text_in[121] ) );
  OAI21_X1 U247 (.B1( ld ) , .ZN( n1100 ) , .B2( n245 ) , .A( n246 ) );
  NAND2_X1 U248 (.A2( ld ) , .ZN( n246 ) , .A1( text_in[122] ) );
  OAI21_X1 U249 (.B1( ld ) , .ZN( n1101 ) , .B2( n247 ) , .A( n248 ) );
  OAI21_X1 U25 (.B1( ld ) , .B2( n23 ) , .A( n24 ) , .ZN( n989 ) );
  NAND2_X1 U250 (.A2( ld ) , .ZN( n248 ) , .A1( text_in[123] ) );
  OAI21_X1 U251 (.B1( ld ) , .ZN( n1102 ) , .B2( n249 ) , .A( n250 ) );
  NAND2_X1 U252 (.A2( ld ) , .ZN( n250 ) , .A1( text_in[124] ) );
  OAI21_X1 U253 (.B1( ld ) , .ZN( n1103 ) , .B2( n251 ) , .A( n252 ) );
  NAND2_X1 U254 (.A2( ld ) , .ZN( n252 ) , .A1( text_in[125] ) );
  OAI21_X1 U255 (.B1( ld ) , .ZN( n1104 ) , .B2( n253 ) , .A( n254 ) );
  NAND2_X1 U256 (.A2( ld ) , .ZN( n254 ) , .A1( text_in[126] ) );
  OAI21_X1 U257 (.B1( ld ) , .ZN( n1105 ) , .B2( n255 ) , .A( n256 ) );
  NAND2_X1 U258 (.A2( ld ) , .ZN( n256 ) , .A1( text_in[127] ) );
  AOI21_X1 U259 (.ZN( n1110 ) , .B1( n1222 ) , .B2( n258 ) , .A( n259 ) );
  NAND2_X1 U26 (.A2( ld ) , .ZN( n24 ) , .A1( text_in[11] ) );
  OAI21_X1 U260 (.ZN( n258 ) , .B1( n260 ) , .B2( n261 ) , .A( n262 ) );
  NOR3_X1 U261 (.A2( ld ) , .ZN( n1111 ) , .A1( n259 ) , .A3( n263 ) );
  AOI22_X1 U262 (.ZN( n263 ) , .A1( n264 ) , .A2( n265 ) , .B1( n266 ) , .B2( n267 ) );
  NOR2_X1 U263 (.A1( n1106 ) , .ZN( n264 ) , .A2( n267 ) );
  INV_X1 U265 (.ZN( n1112 ) , .A( n268 ) );
  OAI21_X1 U266 (.B1( ld ) , .ZN( n268 ) , .B2( n269 ) , .A( rst ) );
  AOI21_X1 U267 (.A( n1106 ) , .B1( n1107 ) , .B2( n265 ) , .ZN( n269 ) );
  INV_X1 U268 (.ZN( n265 ) , .A( n266 ) );
  NAND2_X1 U269 (.A1( n1108 ) , .A2( n262 ) , .ZN( n266 ) );
  OAI21_X1 U27 (.B1( ld ) , .B2( n25 ) , .A( n26 ) , .ZN( n990 ) );
  XNOR2_X1 U270 (.B( n261 ) , .ZN( n262 ) , .A( n977 ) );
  AOI21_X1 U272 (.ZN( n1113 ) , .B1( n1222 ) , .A( n259 ) , .B2( n270 ) );
  INV_X1 U273 (.ZN( n259 ) , .A( rst ) );
  OAI21_X1 U274 (.A( n1108 ) , .B2( n260 ) , .ZN( n270 ) , .B1( n977 ) );
  OAI22_X1 U276 (.ZN( N99 ) , .A1( n1216 ) , .B2( n1220 ) , .A2( n271 ) , .B1( n272 ) );
  XOR2_X1 U278 (.Z( n275 ) , .B( n276 ) , .A( sa22_sr_1 ) );
  XOR2_X1 U279 (.Z( n276 ) , .B( sa32_sr_0 ) , .A( w2_1 ) );
  NAND2_X1 U28 (.A2( ld ) , .ZN( n26 ) , .A1( text_in[12] ) );
  XOR2_X1 U281 (.Z( n278 ) , .B( n279 ) , .A( sa02_sr_0 ) );
  XOR2_X1 U282 (.Z( n271 ) , .A( n67 ) , .B( w2_1 ) );
  OAI22_X1 U284 (.ZN( N98 ) , .A1( n1215 ) , .B2( n1220 ) , .A2( n280 ) , .B1( n281 ) );
  XOR2_X1 U286 (.A( n279 ) , .Z( n283 ) , .B( n284 ) );
  XOR2_X1 U288 (.Z( n280 ) , .A( n65 ) , .B( w2_0 ) );
  OAI21_X1 U29 (.B1( ld ) , .B2( n27 ) , .A( n28 ) , .ZN( n991 ) );
  OAI22_X1 U290 (.ZN( N89 ) , .A1( n1216 ) , .B2( n1217 ) , .A2( n285 ) , .B1( n286 ) );
  XOR2_X1 U292 (.Z( n288 ) , .A( n289 ) , .B( n290 ) );
  XOR2_X1 U294 (.Z( n285 ) , .A( n63 ) , .B( w3_31 ) );
  OAI22_X1 U296 (.ZN( N88 ) , .B2( n1114 ) , .A1( n1212 ) , .A2( n291 ) , .B1( n292 ) );
  XOR2_X1 U298 (.Z( n294 ) , .A( n295 ) , .B( n296 ) );
  OAI21_X1 U3 (.B1( ld ) , .B2( n1 ) , .A( n2 ) , .ZN( n978 ) );
  NAND2_X1 U30 (.A2( ld ) , .ZN( n28 ) , .A1( text_in[13] ) );
  XOR2_X1 U300 (.Z( n291 ) , .A( n61 ) , .B( w3_30 ) );
  OAI22_X1 U302 (.ZN( N87 ) , .A1( n1212 ) , .B2( n1221 ) , .A2( n297 ) , .B1( n298 ) );
  XOR2_X1 U304 (.Z( n300 ) , .A( n301 ) , .B( n302 ) );
  XOR2_X1 U306 (.Z( n297 ) , .A( n59 ) , .B( w3_29 ) );
  OAI22_X1 U308 (.ZN( N86 ) , .B2( n1114 ) , .A1( n1212 ) , .A2( n303 ) , .B1( n304 ) );
  XOR2_X1 U309 (.Z( n304 ) , .A( n305 ) , .B( n306 ) );
  OAI21_X1 U31 (.B1( ld ) , .B2( n29 ) , .A( n30 ) , .ZN( n992 ) );
  XOR2_X1 U310 (.Z( n306 ) , .A( n307 ) , .B( n308 ) );
  XOR2_X1 U311 (.Z( n305 ) , .A( n309 ) , .B( n310 ) );
  XNOR2_X1 U312 (.ZN( n309 ) , .B( sa13_sr_4 ) , .A( w3_28 ) );
  XOR2_X1 U313 (.Z( n303 ) , .A( n57 ) , .B( w3_28 ) );
  OAI22_X1 U315 (.ZN( N85 ) , .B2( n1114 ) , .A1( n1213 ) , .A2( n311 ) , .B1( n312 ) );
  XOR2_X1 U317 (.Z( n314 ) , .A( n315 ) , .B( n316 ) );
  XNOR2_X1 U319 (.ZN( n317 ) , .B( sa13_sr_3 ) , .A( w3_27 ) );
  NAND2_X1 U32 (.A2( ld ) , .ZN( n30 ) , .A1( text_in[14] ) );
  XOR2_X1 U320 (.Z( n311 ) , .A( n55 ) , .B( w3_27 ) );
  OAI22_X1 U322 (.ZN( N84 ) , .B2( n1114 ) , .A1( n1212 ) , .A2( n318 ) , .B1( n319 ) );
  XOR2_X1 U324 (.Z( n321 ) , .A( n322 ) , .B( n323 ) );
  XOR2_X1 U326 (.Z( n318 ) , .A( n53 ) , .B( w3_26 ) );
  OAI22_X1 U328 (.ZN( N83 ) , .B2( n1114 ) , .A1( n1213 ) , .A2( n324 ) , .B1( n325 ) );
  OAI21_X1 U33 (.B1( ld ) , .B2( n31 ) , .A( n32 ) , .ZN( n993 ) );
  XOR2_X1 U330 (.Z( n327 ) , .A( n328 ) , .B( n329 ) );
  XNOR2_X1 U332 (.ZN( n330 ) , .B( sa13_sr_1 ) , .A( w3_25 ) );
  XOR2_X1 U333 (.Z( n324 ) , .A( n51 ) , .B( w3_25 ) );
  OAI22_X1 U335 (.ZN( N82 ) , .B2( n1114 ) , .A1( n1212 ) , .A2( n331 ) , .B1( n332 ) );
  XOR2_X1 U337 (.A( n307 ) , .Z( n334 ) , .B( n335 ) );
  XOR2_X1 U339 (.Z( n331 ) , .A( n49 ) , .B( w3_24 ) );
  NAND2_X1 U34 (.A2( ld ) , .ZN( n32 ) , .A1( text_in[15] ) );
  OAI22_X1 U341 (.ZN( N73 ) , .A1( n1213 ) , .B2( n1219 ) , .A2( n336 ) , .B1( n337 ) );
  XOR2_X1 U342 (.Z( n337 ) , .A( n338 ) , .B( n339 ) );
  XOR2_X1 U343 (.B( n289 ) , .Z( n339 ) , .A( sa03_sr_7 ) );
  XOR2_X1 U346 (.Z( n336 ) , .A( n47 ) , .B( w3_23 ) );
  OAI22_X1 U348 (.ZN( N72 ) , .A1( n1212 ) , .B2( n1217 ) , .A2( n341 ) , .B1( n342 ) );
  OAI21_X1 U35 (.B1( ld ) , .B2( n33 ) , .A( n34 ) , .ZN( n994 ) );
  XOR2_X1 U351 (.Z( n345 ) , .B( sa23_sr_5 ) , .A( w3_22 ) );
  XOR2_X1 U354 (.Z( n341 ) , .A( n45 ) , .B( w3_22 ) );
  OAI22_X1 U356 (.ZN( N71 ) , .A1( n1214 ) , .B2( n1221 ) , .A2( n347 ) , .B1( n348 ) );
  XOR2_X1 U357 (.Z( n348 ) , .A( n349 ) , .B( n350 ) );
  XOR2_X1 U358 (.Z( n350 ) , .B( n351 ) , .A( sa13_sr_4 ) );
  XOR2_X1 U359 (.Z( n351 ) , .B( sa23_sr_4 ) , .A( w3_21 ) );
  NAND2_X1 U36 (.A2( ld ) , .ZN( n34 ) , .A1( text_in[16] ) );
  XOR2_X1 U360 (.B( n301 ) , .Z( n349 ) , .A( n352 ) );
  XOR2_X1 U361 (.Z( n347 ) , .A( n43 ) , .B( w3_21 ) );
  OAI22_X1 U363 (.ZN( N70 ) , .B2( n1114 ) , .A1( n1213 ) , .A2( n353 ) , .B1( n354 ) );
  XOR2_X1 U364 (.Z( n354 ) , .A( n355 ) , .B( n356 ) );
  XOR2_X1 U365 (.Z( n356 ) , .B( n357 ) , .A( sa13_sr_3 ) );
  XOR2_X1 U366 (.Z( n357 ) , .B( sa23_sr_3 ) , .A( w3_20 ) );
  XOR2_X1 U367 (.Z( n355 ) , .A( n358 ) , .B( n359 ) );
  XOR2_X1 U368 (.B( n310 ) , .Z( n358 ) , .A( n360 ) );
  XOR2_X1 U369 (.Z( n353 ) , .A( n41 ) , .B( w3_20 ) );
  OAI21_X1 U37 (.B1( ld ) , .B2( n35 ) , .A( n36 ) , .ZN( n995 ) );
  OAI22_X1 U371 (.ZN( N69 ) , .B2( n1114 ) , .A1( n1212 ) , .A2( n361 ) , .B1( n362 ) );
  XOR2_X1 U374 (.Z( n365 ) , .B( sa23_sr_2 ) , .A( w3_19 ) );
  XOR2_X1 U375 (.B( n359 ) , .Z( n363 ) , .A( n366 ) );
  XOR2_X1 U376 (.B( n315 ) , .Z( n366 ) , .A( n367 ) );
  XOR2_X1 U377 (.Z( n361 ) , .A( n39 ) , .B( w3_19 ) );
  OAI22_X1 U379 (.ZN( N68 ) , .A1( n1214 ) , .B2( n1221 ) , .A2( n368 ) , .B1( n369 ) );
  NAND2_X1 U38 (.A2( ld ) , .ZN( n36 ) , .A1( text_in[17] ) );
  XOR2_X1 U382 (.Z( n372 ) , .B( sa23_sr_1 ) , .A( w3_18 ) );
  XOR2_X1 U383 (.B( n322 ) , .Z( n370 ) , .A( n373 ) );
  XOR2_X1 U384 (.Z( n368 ) , .A( n37 ) , .B( w3_18 ) );
  OAI22_X1 U386 (.ZN( N67 ) , .B2( n1114 ) , .A1( n1213 ) , .A2( n374 ) , .B1( n375 ) );
  XOR2_X1 U389 (.Z( n378 ) , .B( sa23_sr_0 ) , .A( w3_17 ) );
  OAI21_X1 U39 (.B1( ld ) , .B2( n37 ) , .A( n38 ) , .ZN( n996 ) );
  XOR2_X1 U390 (.B( n359 ) , .Z( n376 ) , .A( n379 ) );
  XOR2_X1 U391 (.B( n328 ) , .Z( n379 ) , .A( n380 ) );
  XOR2_X1 U392 (.A( n35 ) , .Z( n374 ) , .B( w3_17 ) );
  OAI22_X1 U394 (.ZN( N66 ) , .A1( n1214 ) , .B2( n1220 ) , .A2( n381 ) , .B1( n382 ) );
  XOR2_X1 U396 (.A( n335 ) , .B( n359 ) , .Z( n384 ) );
  XNOR2_X1 U397 (.ZN( n359 ) , .B( n385 ) , .A( sa13_sr_7 ) );
  XOR2_X1 U399 (.A( n33 ) , .Z( n381 ) , .B( w3_16 ) );
  NAND2_X1 U4 (.A2( ld ) , .ZN( n2 ) , .A1( text_in[0] ) );
  NAND2_X1 U40 (.A2( ld ) , .ZN( n38 ) , .A1( text_in[18] ) );
  OAI22_X1 U401 (.ZN( N57 ) , .A1( n1212 ) , .B2( n1221 ) , .A2( n387 ) , .B1( n388 ) );
  XOR2_X1 U403 (.A( n295 ) , .B( n307 ) , .Z( n390 ) );
  XOR2_X1 U404 (.Z( n295 ) , .A( sa23_sr_6 ) , .B( sa33_sr_6 ) );
  XOR2_X1 U406 (.A( n31 ) , .Z( n387 ) , .B( w3_15 ) );
  OAI22_X1 U408 (.ZN( N56 ) , .B2( n1114 ) , .A1( n1213 ) , .A2( n391 ) , .B1( n392 ) );
  OAI21_X1 U41 (.B1( ld ) , .B2( n39 ) , .A( n40 ) , .ZN( n997 ) );
  XOR2_X1 U410 (.A( n290 ) , .B( n301 ) , .Z( n394 ) );
  XOR2_X1 U411 (.Z( n301 ) , .A( sa23_sr_5 ) , .B( sa33_sr_5 ) );
  XOR2_X1 U413 (.A( n29 ) , .Z( n391 ) , .B( w3_14 ) );
  OAI22_X1 U415 (.ZN( N55 ) , .A1( n1216 ) , .B2( n1221 ) , .A2( n395 ) , .B1( n396 ) );
  XOR2_X1 U417 (.A( n296 ) , .B( n310 ) , .Z( n398 ) );
  XOR2_X1 U418 (.Z( n310 ) , .A( sa23_sr_4 ) , .B( sa33_sr_4 ) );
  NAND2_X1 U42 (.A2( ld ) , .ZN( n40 ) , .A1( text_in[19] ) );
  XOR2_X1 U420 (.A( n27 ) , .Z( n395 ) , .B( w3_13 ) );
  OAI22_X1 U422 (.ZN( N54 ) , .A1( n1216 ) , .B2( n1220 ) , .A2( n399 ) , .B1( n400 ) );
  XOR2_X1 U423 (.Z( n400 ) , .A( n401 ) , .B( n402 ) );
  XOR2_X1 U424 (.A( n302 ) , .B( n315 ) , .Z( n402 ) );
  XOR2_X1 U425 (.Z( n315 ) , .A( sa23_sr_3 ) , .B( sa33_sr_3 ) );
  XOR2_X1 U426 (.B( n289 ) , .Z( n401 ) , .A( n403 ) );
  XNOR2_X1 U427 (.ZN( n403 ) , .B( sa33_sr_4 ) , .A( w3_12 ) );
  XOR2_X1 U428 (.A( n25 ) , .Z( n399 ) , .B( w3_12 ) );
  OAI21_X1 U43 (.B1( ld ) , .B2( n41 ) , .A( n42 ) , .ZN( n998 ) );
  OAI22_X1 U430 (.ZN( N53 ) , .A1( n1216 ) , .B2( n1220 ) , .A2( n404 ) , .B1( n405 ) );
  XOR2_X1 U432 (.A( n308 ) , .B( n322 ) , .Z( n407 ) );
  XOR2_X1 U433 (.Z( n322 ) , .A( sa23_sr_2 ) , .B( sa33_sr_2 ) );
  XNOR2_X1 U435 (.ZN( n408 ) , .B( sa33_sr_3 ) , .A( w3_11 ) );
  XOR2_X1 U436 (.A( n23 ) , .Z( n404 ) , .B( w3_11 ) );
  OAI22_X1 U438 (.ZN( N52 ) , .B2( n1114 ) , .A1( n1214 ) , .A2( n409 ) , .B1( n410 ) );
  NAND2_X1 U44 (.A2( ld ) , .ZN( n42 ) , .A1( text_in[20] ) );
  XOR2_X1 U440 (.A( n316 ) , .B( n328 ) , .Z( n412 ) );
  XOR2_X1 U441 (.Z( n328 ) , .A( sa23_sr_1 ) , .B( sa33_sr_1 ) );
  XOR2_X1 U443 (.A( n21 ) , .Z( n409 ) , .B( w3_10 ) );
  OAI22_X1 U445 (.ZN( N51 ) , .A1( n1214 ) , .B2( n1217 ) , .A2( n413 ) , .B1( n414 ) );
  XOR2_X1 U447 (.A( n323 ) , .B( n335 ) , .Z( n416 ) );
  XOR2_X1 U448 (.Z( n335 ) , .A( sa23_sr_0 ) , .B( sa33_sr_0 ) );
  OAI21_X1 U45 (.B1( ld ) , .B2( n43 ) , .A( n44 ) , .ZN( n999 ) );
  XNOR2_X1 U450 (.ZN( n417 ) , .B( sa33_sr_1 ) , .A( w3_9 ) );
  XOR2_X1 U451 (.A( n19 ) , .Z( n413 ) , .B( w3_9 ) );
  XOR2_X1 U453 (.Z( N505 ) , .B( sa33_sr_0 ) , .A( w3_0 ) );
  XOR2_X1 U454 (.Z( N504 ) , .B( sa33_sr_1 ) , .A( w3_1 ) );
  XOR2_X1 U455 (.Z( N503 ) , .B( sa33_sr_2 ) , .A( w3_2 ) );
  XOR2_X1 U456 (.Z( N502 ) , .B( sa33_sr_3 ) , .A( w3_3 ) );
  XOR2_X1 U457 (.Z( N501 ) , .B( sa33_sr_4 ) , .A( w3_4 ) );
  XOR2_X1 U458 (.Z( N500 ) , .B( sa33_sr_5 ) , .A( w3_5 ) );
  OAI22_X1 U459 (.ZN( N50 ) , .A1( n1214 ) , .B2( n1218 ) , .A2( n418 ) , .B1( n419 ) );
  NAND2_X1 U46 (.A2( ld ) , .ZN( n44 ) , .A1( text_in[21] ) );
  XOR2_X1 U461 (.A( n289 ) , .B( n329 ) , .Z( n421 ) );
  XOR2_X1 U462 (.Z( n289 ) , .A( sa23_sr_7 ) , .B( sa33_sr_7 ) );
  XOR2_X1 U464 (.A( n17 ) , .Z( n418 ) , .B( w3_8 ) );
  XOR2_X1 U466 (.Z( N499 ) , .B( sa33_sr_6 ) , .A( w3_6 ) );
  XOR2_X1 U467 (.Z( N498 ) , .B( sa33_sr_7 ) , .A( w3_7 ) );
  XOR2_X1 U468 (.Z( N497 ) , .B( sa32_sr_0 ) , .A( w2_0 ) );
  XOR2_X1 U469 (.Z( N496 ) , .B( sa32_sr_1 ) , .A( w2_1 ) );
  OAI21_X1 U47 (.B1( ld ) , .ZN( n1000 ) , .B2( n45 ) , .A( n46 ) );
  XOR2_X1 U471 (.Z( N494 ) , .B( sa32_sr_3 ) , .A( w2_3 ) );
  XOR2_X1 U472 (.Z( N493 ) , .B( sa32_sr_4 ) , .A( w2_4 ) );
  XOR2_X1 U473 (.Z( N492 ) , .B( sa32_sr_5 ) , .A( w2_5 ) );
  XOR2_X1 U474 (.Z( N491 ) , .B( sa32_sr_6 ) , .A( w2_6 ) );
  XOR2_X1 U475 (.Z( N490 ) , .B( sa32_sr_7 ) , .A( w2_7 ) );
  XOR2_X1 U476 (.Z( N489 ) , .B( sa31_sr_0 ) , .A( w1_0 ) );
  XOR2_X1 U477 (.Z( N488 ) , .B( sa31_sr_1 ) , .A( w1_1 ) );
  XOR2_X1 U478 (.Z( N487 ) , .B( sa31_sr_2 ) , .A( w1_2 ) );
  XOR2_X1 U479 (.Z( N486 ) , .B( sa31_sr_3 ) , .A( w1_3 ) );
  NAND2_X1 U48 (.A2( ld ) , .ZN( n46 ) , .A1( text_in[22] ) );
  XOR2_X1 U480 (.Z( N485 ) , .B( sa31_sr_4 ) , .A( w1_4 ) );
  XOR2_X1 U481 (.Z( N484 ) , .B( sa31_sr_5 ) , .A( w1_5 ) );
  XOR2_X1 U482 (.Z( N483 ) , .B( sa31_sr_6 ) , .A( w1_6 ) );
  XOR2_X1 U483 (.Z( N482 ) , .B( sa31_sr_7 ) , .A( w1_7 ) );
  XOR2_X1 U484 (.Z( N481 ) , .B( sa30_sr_0 ) , .A( w0_0 ) );
  XOR2_X1 U485 (.Z( N480 ) , .B( sa30_sr_1 ) , .A( w0_1 ) );
  XOR2_X1 U486 (.Z( N479 ) , .B( sa30_sr_2 ) , .A( w0_2 ) );
  XOR2_X1 U487 (.Z( N478 ) , .B( sa30_sr_3 ) , .A( w0_3 ) );
  XOR2_X1 U488 (.Z( N477 ) , .B( sa30_sr_4 ) , .A( w0_4 ) );
  XOR2_X1 U489 (.Z( N476 ) , .B( sa30_sr_5 ) , .A( w0_5 ) );
  OAI21_X1 U49 (.B1( ld ) , .ZN( n1001 ) , .B2( n47 ) , .A( n48 ) );
  XOR2_X1 U490 (.Z( N475 ) , .B( sa30_sr_6 ) , .A( w0_6 ) );
  XOR2_X1 U491 (.Z( N474 ) , .B( sa30_sr_7 ) , .A( w0_7 ) );
  XOR2_X1 U492 (.Z( N473 ) , .B( sa23_sr_0 ) , .A( w3_8 ) );
  XOR2_X1 U493 (.Z( N472 ) , .B( sa23_sr_1 ) , .A( w3_9 ) );
  XOR2_X1 U494 (.Z( N471 ) , .B( sa23_sr_2 ) , .A( w3_10 ) );
  XOR2_X1 U495 (.Z( N470 ) , .B( sa23_sr_3 ) , .A( w3_11 ) );
  XOR2_X1 U496 (.Z( N469 ) , .B( sa23_sr_4 ) , .A( w3_12 ) );
  XOR2_X1 U497 (.Z( N468 ) , .B( sa23_sr_5 ) , .A( w3_13 ) );
  XOR2_X1 U498 (.Z( N467 ) , .B( sa23_sr_6 ) , .A( w3_14 ) );
  XOR2_X1 U499 (.Z( N466 ) , .B( sa23_sr_7 ) , .A( w3_15 ) );
  OAI21_X1 U5 (.B1( ld ) , .B2( n3 ) , .A( n4 ) , .ZN( n979 ) );
  NAND2_X1 U50 (.A2( ld ) , .ZN( n48 ) , .A1( text_in[23] ) );
  XOR2_X1 U500 (.Z( N465 ) , .B( sa22_sr_0 ) , .A( w2_8 ) );
  XOR2_X1 U501 (.Z( N464 ) , .B( sa22_sr_1 ) , .A( w2_9 ) );
  XOR2_X1 U503 (.Z( N462 ) , .B( sa22_sr_3 ) , .A( w2_11 ) );
  XOR2_X1 U504 (.Z( N461 ) , .B( sa22_sr_4 ) , .A( w2_12 ) );
  XOR2_X1 U505 (.Z( N460 ) , .B( sa22_sr_5 ) , .A( w2_13 ) );
  XOR2_X1 U506 (.Z( N459 ) , .B( sa22_sr_6 ) , .A( w2_14 ) );
  XOR2_X1 U507 (.Z( N458 ) , .B( sa22_sr_7 ) , .A( w2_15 ) );
  XOR2_X1 U508 (.Z( N457 ) , .B( sa21_sr_0 ) , .A( w1_8 ) );
  XOR2_X1 U509 (.Z( N456 ) , .B( sa21_sr_1 ) , .A( w1_9 ) );
  OAI21_X1 U51 (.B1( ld ) , .ZN( n1002 ) , .B2( n49 ) , .A( n50 ) );
  XOR2_X1 U510 (.Z( N455 ) , .B( sa21_sr_2 ) , .A( w1_10 ) );
  XOR2_X1 U511 (.Z( N454 ) , .B( sa21_sr_3 ) , .A( w1_11 ) );
  XOR2_X1 U512 (.Z( N453 ) , .B( sa21_sr_4 ) , .A( w1_12 ) );
  XOR2_X1 U513 (.Z( N452 ) , .B( sa21_sr_5 ) , .A( w1_13 ) );
  XOR2_X1 U514 (.Z( N451 ) , .B( sa21_sr_6 ) , .A( w1_14 ) );
  XOR2_X1 U515 (.Z( N450 ) , .B( sa21_sr_7 ) , .A( w1_15 ) );
  XOR2_X1 U516 (.Z( N449 ) , .B( sa20_sr_0 ) , .A( w0_8 ) );
  XOR2_X1 U517 (.Z( N448 ) , .B( sa20_sr_1 ) , .A( w0_9 ) );
  XOR2_X1 U518 (.Z( N447 ) , .B( sa20_sr_2 ) , .A( w0_10 ) );
  XOR2_X1 U519 (.Z( N446 ) , .B( sa20_sr_3 ) , .A( w0_11 ) );
  NAND2_X1 U52 (.A2( ld ) , .ZN( n50 ) , .A1( text_in[24] ) );
  XOR2_X1 U520 (.Z( N445 ) , .B( sa20_sr_4 ) , .A( w0_12 ) );
  XOR2_X1 U521 (.Z( N444 ) , .B( sa20_sr_5 ) , .A( w0_13 ) );
  XOR2_X1 U522 (.Z( N443 ) , .B( sa20_sr_6 ) , .A( w0_14 ) );
  XOR2_X1 U523 (.Z( N442 ) , .B( sa20_sr_7 ) , .A( w0_15 ) );
  XOR2_X1 U524 (.Z( N441 ) , .B( sa13_sr_0 ) , .A( w3_16 ) );
  XOR2_X1 U525 (.Z( N440 ) , .B( sa13_sr_1 ) , .A( w3_17 ) );
  XOR2_X1 U526 (.Z( N439 ) , .B( sa13_sr_2 ) , .A( w3_18 ) );
  XOR2_X1 U527 (.Z( N438 ) , .B( sa13_sr_3 ) , .A( w3_19 ) );
  XOR2_X1 U528 (.Z( N437 ) , .B( sa13_sr_4 ) , .A( w3_20 ) );
  XOR2_X1 U529 (.Z( N436 ) , .B( sa13_sr_5 ) , .A( w3_21 ) );
  OAI21_X1 U53 (.B1( ld ) , .ZN( n1003 ) , .B2( n51 ) , .A( n52 ) );
  XOR2_X1 U530 (.Z( N435 ) , .B( sa13_sr_6 ) , .A( w3_22 ) );
  XOR2_X1 U531 (.Z( N434 ) , .B( sa13_sr_7 ) , .A( w3_23 ) );
  XOR2_X1 U532 (.Z( N433 ) , .B( sa12_sr_0 ) , .A( w2_16 ) );
  XOR2_X1 U533 (.Z( N432 ) , .B( sa12_sr_1 ) , .A( w2_17 ) );
  XOR2_X1 U534 (.Z( N431 ) , .B( sa12_sr_2 ) , .A( w2_18 ) );
  XOR2_X1 U535 (.Z( N430 ) , .B( sa12_sr_3 ) , .A( w2_19 ) );
  XOR2_X1 U536 (.Z( N429 ) , .B( sa12_sr_4 ) , .A( w2_20 ) );
  XOR2_X1 U537 (.Z( N428 ) , .B( sa12_sr_5 ) , .A( w2_21 ) );
  XOR2_X1 U538 (.Z( N427 ) , .B( sa12_sr_6 ) , .A( w2_22 ) );
  XOR2_X1 U539 (.Z( N426 ) , .B( sa12_sr_7 ) , .A( w2_23 ) );
  NAND2_X1 U54 (.A2( ld ) , .ZN( n52 ) , .A1( text_in[25] ) );
  XOR2_X1 U540 (.Z( N425 ) , .B( sa11_sr_0 ) , .A( w1_16 ) );
  XOR2_X1 U541 (.Z( N424 ) , .B( sa11_sr_1 ) , .A( w1_17 ) );
  XOR2_X1 U543 (.Z( N422 ) , .B( sa11_sr_3 ) , .A( w1_19 ) );
  XOR2_X1 U544 (.Z( N421 ) , .B( sa11_sr_4 ) , .A( w1_20 ) );
  XOR2_X1 U545 (.Z( N420 ) , .B( sa11_sr_5 ) , .A( w1_21 ) );
  XOR2_X1 U546 (.Z( N419 ) , .B( sa11_sr_6 ) , .A( w1_22 ) );
  XOR2_X1 U547 (.Z( N418 ) , .B( sa11_sr_7 ) , .A( w1_23 ) );
  XOR2_X1 U548 (.Z( N417 ) , .B( sa10_sr_0 ) , .A( w0_16 ) );
  XOR2_X1 U549 (.Z( N416 ) , .B( sa10_sr_1 ) , .A( w0_17 ) );
  OAI21_X1 U55 (.B1( ld ) , .ZN( n1004 ) , .B2( n53 ) , .A( n54 ) );
  XOR2_X1 U551 (.Z( N414 ) , .B( sa10_sr_3 ) , .A( w0_19 ) );
  XOR2_X1 U552 (.Z( N413 ) , .B( sa10_sr_4 ) , .A( w0_20 ) );
  XOR2_X1 U553 (.Z( N412 ) , .B( sa10_sr_5 ) , .A( w0_21 ) );
  XOR2_X1 U554 (.Z( N411 ) , .B( sa10_sr_6 ) , .A( w0_22 ) );
  XOR2_X1 U555 (.Z( N410 ) , .B( sa10_sr_7 ) , .A( w0_23 ) );
  OAI22_X1 U556 (.ZN( N41 ) , .B2( n1114 ) , .A1( n1214 ) , .A2( n422 ) , .B1( n423 ) );
  XOR2_X1 U557 (.Z( n423 ) , .A( n424 ) , .B( n425 ) );
  XOR2_X1 U558 (.B( n307 ) , .Z( n425 ) , .A( sa03_sr_6 ) );
  XOR2_X1 U559 (.Z( n307 ) , .A( sa03_sr_7 ) , .B( sa13_sr_7 ) );
  NAND2_X1 U56 (.A2( ld ) , .ZN( n54 ) , .A1( text_in[26] ) );
  XOR2_X1 U560 (.A( n385 ) , .Z( n424 ) , .B( n426 ) );
  XOR2_X1 U561 (.Z( n426 ) , .B( sa33_sr_6 ) , .A( w3_7 ) );
  INV_X1 U562 (.ZN( n385 ) , .A( sa23_sr_7 ) );
  XOR2_X1 U563 (.A( n15 ) , .Z( n422 ) , .B( w3_7 ) );
  XOR2_X1 U565 (.Z( N409 ) , .B( sa03_sr_0 ) , .A( w3_24 ) );
  XOR2_X1 U566 (.Z( N408 ) , .B( sa03_sr_1 ) , .A( w3_25 ) );
  XOR2_X1 U567 (.Z( N407 ) , .B( sa03_sr_2 ) , .A( w3_26 ) );
  XOR2_X1 U568 (.Z( N406 ) , .B( sa03_sr_3 ) , .A( w3_27 ) );
  XOR2_X1 U569 (.Z( N405 ) , .B( sa03_sr_4 ) , .A( w3_28 ) );
  OAI21_X1 U57 (.B1( ld ) , .ZN( n1005 ) , .B2( n55 ) , .A( n56 ) );
  XOR2_X1 U570 (.Z( N404 ) , .B( sa03_sr_5 ) , .A( w3_29 ) );
  XOR2_X1 U571 (.Z( N403 ) , .B( sa03_sr_6 ) , .A( w3_30 ) );
  XOR2_X1 U572 (.Z( N402 ) , .B( sa03_sr_7 ) , .A( w3_31 ) );
  XOR2_X1 U573 (.Z( N401 ) , .B( sa02_sr_0 ) , .A( w2_24 ) );
  XOR2_X1 U574 (.Z( N400 ) , .B( sa02_sr_1 ) , .A( w2_25 ) );
  OAI22_X1 U575 (.ZN( N40 ) , .A1( n1214 ) , .B2( n1221 ) , .A2( n427 ) , .B1( n428 ) );
  XOR2_X1 U578 (.Z( n431 ) , .B( sa33_sr_5 ) , .A( w3_6 ) );
  XOR2_X1 U579 (.B( n290 ) , .A( n352 ) , .Z( n429 ) );
  NAND2_X1 U58 (.A2( ld ) , .ZN( n56 ) , .A1( text_in[27] ) );
  XOR2_X1 U580 (.Z( n290 ) , .A( sa03_sr_6 ) , .B( sa13_sr_6 ) );
  INV_X1 U581 (.ZN( n352 ) , .A( sa03_sr_5 ) );
  XOR2_X1 U582 (.A( n13 ) , .Z( n427 ) , .B( w3_6 ) );
  XOR2_X1 U584 (.Z( N399 ) , .B( sa02_sr_2 ) , .A( w2_26 ) );
  XOR2_X1 U585 (.Z( N398 ) , .B( sa02_sr_3 ) , .A( w2_27 ) );
  XOR2_X1 U586 (.Z( N397 ) , .B( sa02_sr_4 ) , .A( w2_28 ) );
  XOR2_X1 U587 (.Z( N396 ) , .B( sa02_sr_5 ) , .A( w2_29 ) );
  XOR2_X1 U588 (.Z( N395 ) , .B( sa02_sr_6 ) , .A( w2_30 ) );
  XOR2_X1 U589 (.Z( N394 ) , .B( sa02_sr_7 ) , .A( w2_31 ) );
  OAI21_X1 U59 (.B1( ld ) , .ZN( n1006 ) , .B2( n57 ) , .A( n58 ) );
  XOR2_X1 U590 (.Z( N393 ) , .B( sa01_sr_0 ) , .A( w1_24 ) );
  XOR2_X1 U591 (.Z( N392 ) , .B( sa01_sr_1 ) , .A( w1_25 ) );
  XOR2_X1 U592 (.Z( N391 ) , .B( sa01_sr_2 ) , .A( w1_26 ) );
  XOR2_X1 U593 (.Z( N390 ) , .B( sa01_sr_3 ) , .A( w1_27 ) );
  OAI22_X1 U594 (.ZN( N39 ) , .A1( n1214 ) , .B2( n1218 ) , .A2( n432 ) , .B1( n433 ) );
  XOR2_X1 U597 (.Z( n436 ) , .B( sa33_sr_4 ) , .A( w3_5 ) );
  XOR2_X1 U598 (.B( n296 ) , .A( n360 ) , .Z( n434 ) );
  XOR2_X1 U599 (.Z( n296 ) , .A( sa03_sr_5 ) , .B( sa13_sr_5 ) );
  NAND2_X1 U6 (.A2( ld ) , .ZN( n4 ) , .A1( text_in[1] ) );
  NAND2_X1 U60 (.A2( ld ) , .ZN( n58 ) , .A1( text_in[28] ) );
  INV_X1 U600 (.ZN( n360 ) , .A( sa03_sr_4 ) );
  XOR2_X1 U601 (.A( n11 ) , .Z( n432 ) , .B( w3_5 ) );
  XOR2_X1 U603 (.Z( N389 ) , .B( sa01_sr_4 ) , .A( w1_28 ) );
  XOR2_X1 U604 (.Z( N388 ) , .B( sa01_sr_5 ) , .A( w1_29 ) );
  XOR2_X1 U605 (.Z( N387 ) , .B( sa01_sr_6 ) , .A( w1_30 ) );
  XOR2_X1 U606 (.Z( N386 ) , .B( sa01_sr_7 ) , .A( w1_31 ) );
  XOR2_X1 U607 (.Z( N385 ) , .B( sa00_sr_0 ) , .A( w0_24 ) );
  XOR2_X1 U608 (.Z( N384 ) , .B( sa00_sr_1 ) , .A( w0_25 ) );
  XOR2_X1 U609 (.Z( N383 ) , .B( sa00_sr_2 ) , .A( w0_26 ) );
  OAI21_X1 U61 (.B1( ld ) , .ZN( n1007 ) , .B2( n59 ) , .A( n60 ) );
  XOR2_X1 U610 (.Z( N382 ) , .B( sa00_sr_3 ) , .A( w0_27 ) );
  XOR2_X1 U611 (.Z( N381 ) , .B( sa00_sr_4 ) , .A( w0_28 ) );
  XOR2_X1 U612 (.Z( N380 ) , .B( sa00_sr_5 ) , .A( w0_29 ) );
  OAI22_X1 U613 (.ZN( N38 ) , .A1( n1214 ) , .B2( n1221 ) , .A2( n437 ) , .B1( n438 ) );
  XOR2_X1 U614 (.Z( n438 ) , .A( n439 ) , .B( n440 ) );
  XOR2_X1 U615 (.Z( n440 ) , .B( n441 ) , .A( sa23_sr_4 ) );
  XOR2_X1 U616 (.Z( n441 ) , .B( sa33_sr_3 ) , .A( w3_4 ) );
  XOR2_X1 U617 (.Z( n439 ) , .A( n442 ) , .B( n443 ) );
  XOR2_X1 U618 (.B( n302 ) , .A( n367 ) , .Z( n442 ) );
  XOR2_X1 U619 (.Z( n302 ) , .A( sa03_sr_4 ) , .B( sa13_sr_4 ) );
  NAND2_X1 U62 (.A2( ld ) , .ZN( n60 ) , .A1( text_in[29] ) );
  INV_X1 U620 (.ZN( n367 ) , .A( sa03_sr_3 ) );
  XOR2_X1 U621 (.Z( n437 ) , .A( n9 ) , .B( w3_4 ) );
  XOR2_X1 U623 (.Z( N379 ) , .B( sa00_sr_6 ) , .A( w0_30 ) );
  XOR2_X1 U624 (.Z( N378 ) , .B( sa00_sr_7 ) , .A( w0_31 ) );
  OAI22_X1 U625 (.ZN( N37 ) , .B2( n1114 ) , .A1( n1214 ) , .A2( n444 ) , .B1( n445 ) );
  XOR2_X1 U628 (.Z( n448 ) , .B( sa33_sr_2 ) , .A( w3_3 ) );
  XOR2_X1 U629 (.B( n443 ) , .Z( n446 ) , .A( n449 ) );
  OAI21_X1 U63 (.B1( ld ) , .ZN( n1008 ) , .B2( n61 ) , .A( n62 ) );
  XOR2_X1 U630 (.B( n308 ) , .A( n373 ) , .Z( n449 ) );
  XOR2_X1 U631 (.Z( n308 ) , .A( sa03_sr_3 ) , .B( sa13_sr_3 ) );
  INV_X1 U632 (.ZN( n373 ) , .A( sa03_sr_2 ) );
  XOR2_X1 U633 (.Z( n444 ) , .A( n7 ) , .B( w3_3 ) );
  OAI22_X1 U635 (.ZN( N36 ) , .A1( n1214 ) , .B2( n1220 ) , .A2( n450 ) , .B1( n451 ) );
  XOR2_X1 U636 (.Z( n451 ) , .A( n452 ) , .B( n453 ) );
  XOR2_X1 U637 (.Z( n453 ) , .B( n454 ) , .A( sa23_sr_2 ) );
  XOR2_X1 U638 (.Z( n454 ) , .B( sa33_sr_1 ) , .A( w3_2 ) );
  XOR2_X1 U639 (.B( n316 ) , .A( n380 ) , .Z( n452 ) );
  NAND2_X1 U64 (.A2( ld ) , .ZN( n62 ) , .A1( text_in[30] ) );
  XOR2_X1 U640 (.Z( n316 ) , .A( sa03_sr_2 ) , .B( sa13_sr_2 ) );
  INV_X1 U641 (.ZN( n380 ) , .A( sa03_sr_1 ) );
  XOR2_X1 U642 (.Z( n450 ) , .A( n5 ) , .B( w3_2 ) );
  OAI22_X1 U644 (.ZN( N35 ) , .A1( n1214 ) , .B2( n1217 ) , .A2( n455 ) , .B1( n456 ) );
  XOR2_X1 U647 (.Z( n459 ) , .B( sa33_sr_0 ) , .A( w3_1 ) );
  XOR2_X1 U648 (.B( n443 ) , .Z( n457 ) , .A( n460 ) );
  XOR2_X1 U649 (.B( n323 ) , .A( n386 ) , .Z( n460 ) );
  OAI21_X1 U65 (.B1( ld ) , .ZN( n1009 ) , .B2( n63 ) , .A( n64 ) );
  XOR2_X1 U650 (.Z( n323 ) , .A( sa03_sr_1 ) , .B( sa13_sr_1 ) );
  INV_X1 U651 (.ZN( n386 ) , .A( sa03_sr_0 ) );
  XOR2_X1 U652 (.A( n3 ) , .Z( n455 ) , .B( w3_1 ) );
  OAI22_X1 U654 (.ZN( N34 ) , .A1( n1214 ) , .B2( n1218 ) , .A2( n461 ) , .B1( n462 ) );
  XOR2_X1 U656 (.A( n329 ) , .B( n443 ) , .Z( n464 ) );
  XOR2_X1 U657 (.Z( n443 ) , .A( sa03_sr_7 ) , .B( sa33_sr_7 ) );
  XOR2_X1 U658 (.Z( n329 ) , .A( sa03_sr_0 ) , .B( sa13_sr_0 ) );
  NAND2_X1 U66 (.A2( ld ) , .ZN( n64 ) , .A1( text_in[31] ) );
  XOR2_X1 U660 (.A( n1 ) , .Z( n461 ) , .B( w3_0 ) );
  OAI22_X1 U662 (.ZN( N281 ) , .A1( n1214 ) , .B2( n1221 ) , .A2( n465 ) , .B1( n466 ) );
  XOR2_X1 U664 (.Z( n468 ) , .A( n469 ) , .B( n470 ) );
  INV_X1 U666 (.ZN( n471 ) , .A( sa10_sr_7 ) );
  XOR2_X1 U667 (.A( n255 ) , .Z( n465 ) , .B( w0_31 ) );
  OAI22_X1 U669 (.ZN( N280 ) , .B2( n1114 ) , .A1( n1214 ) , .A2( n472 ) , .B1( n473 ) );
  OAI21_X1 U67 (.B1( ld ) , .ZN( n1010 ) , .B2( n65 ) , .A( n66 ) );
  XOR2_X1 U671 (.Z( n475 ) , .A( n476 ) , .B( n477 ) );
  XOR2_X1 U673 (.A( n253 ) , .Z( n472 ) , .B( w0_30 ) );
  OAI22_X1 U675 (.ZN( N279 ) , .A1( n1212 ) , .B2( n1218 ) , .A2( n478 ) , .B1( n479 ) );
  XOR2_X1 U677 (.Z( n481 ) , .A( n482 ) , .B( n483 ) );
  XOR2_X1 U679 (.A( n251 ) , .Z( n478 ) , .B( w0_29 ) );
  NAND2_X1 U68 (.A2( ld ) , .ZN( n66 ) , .A1( text_in[32] ) );
  OAI22_X1 U681 (.ZN( N278 ) , .B2( n1114 ) , .A1( n1213 ) , .A2( n484 ) , .B1( n485 ) );
  XOR2_X1 U682 (.Z( n485 ) , .A( n486 ) , .B( n487 ) );
  XOR2_X1 U683 (.Z( n487 ) , .A( n488 ) , .B( n489 ) );
  XOR2_X1 U684 (.Z( n486 ) , .A( n490 ) , .B( n491 ) );
  XNOR2_X1 U685 (.ZN( n490 ) , .B( sa10_sr_4 ) , .A( w0_28 ) );
  XOR2_X1 U686 (.A( n249 ) , .Z( n484 ) , .B( w0_28 ) );
  OAI22_X1 U688 (.ZN( N277 ) , .A1( n1212 ) , .B2( n1219 ) , .A2( n492 ) , .B1( n493 ) );
  OAI21_X1 U69 (.B1( ld ) , .ZN( n1011 ) , .B2( n67 ) , .A( n68 ) );
  XOR2_X1 U690 (.Z( n495 ) , .A( n496 ) , .B( n497 ) );
  XNOR2_X1 U692 (.ZN( n498 ) , .B( sa10_sr_3 ) , .A( w0_27 ) );
  XOR2_X1 U693 (.A( n247 ) , .Z( n492 ) , .B( w0_27 ) );
  OAI22_X1 U695 (.ZN( N276 ) , .A1( n1212 ) , .B2( n1220 ) , .A2( n499 ) , .B1( n500 ) );
  XOR2_X1 U697 (.Z( n502 ) , .A( n503 ) , .B( n504 ) );
  XOR2_X1 U699 (.A( n245 ) , .Z( n499 ) , .B( w0_26 ) );
  OAI21_X1 U7 (.B1( ld ) , .B2( n5 ) , .A( n6 ) , .ZN( n980 ) );
  NAND2_X1 U70 (.A2( ld ) , .ZN( n68 ) , .A1( text_in[33] ) );
  OAI22_X1 U701 (.ZN( N275 ) , .A1( n1213 ) , .B2( n1220 ) , .A2( n505 ) , .B1( n506 ) );
  XOR2_X1 U703 (.Z( n508 ) , .A( n509 ) , .B( n510 ) );
  XNOR2_X1 U705 (.ZN( n511 ) , .B( sa10_sr_1 ) , .A( w0_25 ) );
  XOR2_X1 U706 (.A( n243 ) , .Z( n505 ) , .B( w0_25 ) );
  OAI22_X1 U708 (.ZN( N274 ) , .A1( n1216 ) , .B2( n1221 ) , .A2( n512 ) , .B1( n513 ) );
  OAI21_X1 U71 (.B1( ld ) , .ZN( n1012 ) , .B2( n69 ) , .A( n70 ) );
  XOR2_X1 U710 (.A( n488 ) , .Z( n515 ) , .B( n516 ) );
  XOR2_X1 U712 (.A( n241 ) , .Z( n512 ) , .B( w0_24 ) );
  OAI22_X1 U714 (.ZN( N265 ) , .B2( n1114 ) , .A1( n1215 ) , .A2( n517 ) , .B1( n518 ) );
  XOR2_X1 U715 (.Z( n518 ) , .A( n519 ) , .B( n520 ) );
  XOR2_X1 U716 (.B( n469 ) , .Z( n520 ) , .A( sa00_sr_7 ) );
  XNOR2_X1 U717 (.ZN( n519 ) , .B( n521 ) , .A( sa10_sr_6 ) );
  XOR2_X1 U718 (.Z( n521 ) , .B( sa20_sr_6 ) , .A( w0_23 ) );
  XOR2_X1 U719 (.A( n239 ) , .Z( n517 ) , .B( w0_23 ) );
  NAND2_X1 U72 (.A2( ld ) , .ZN( n70 ) , .A1( text_in[34] ) );
  OAI22_X1 U721 (.ZN( N264 ) , .A1( n1213 ) , .B2( n1220 ) , .A2( n522 ) , .B1( n523 ) );
  XOR2_X1 U724 (.Z( n526 ) , .B( sa20_sr_5 ) , .A( w0_22 ) );
  XOR2_X1 U727 (.A( n237 ) , .Z( n522 ) , .B( w0_22 ) );
  OAI22_X1 U729 (.ZN( N263 ) , .A1( n1213 ) , .B2( n1221 ) , .A2( n528 ) , .B1( n529 ) );
  OAI21_X1 U73 (.B1( ld ) , .ZN( n1013 ) , .B2( n71 ) , .A( n72 ) );
  XOR2_X1 U730 (.Z( n529 ) , .A( n530 ) , .B( n531 ) );
  XOR2_X1 U731 (.Z( n531 ) , .B( n532 ) , .A( sa10_sr_4 ) );
  XOR2_X1 U732 (.Z( n532 ) , .B( sa20_sr_4 ) , .A( w0_21 ) );
  XNOR2_X1 U733 (.B( n482 ) , .ZN( n530 ) , .A( sa00_sr_5 ) );
  XOR2_X1 U734 (.A( n235 ) , .Z( n528 ) , .B( w0_21 ) );
  OAI22_X1 U736 (.ZN( N262 ) , .A1( n1213 ) , .B2( n1218 ) , .A2( n533 ) , .B1( n534 ) );
  XOR2_X1 U737 (.Z( n534 ) , .A( n535 ) , .B( n536 ) );
  XOR2_X1 U738 (.Z( n536 ) , .B( n537 ) , .A( sa10_sr_3 ) );
  XOR2_X1 U739 (.Z( n537 ) , .B( sa20_sr_3 ) , .A( w0_20 ) );
  NAND2_X1 U74 (.A2( ld ) , .ZN( n72 ) , .A1( text_in[35] ) );
  XOR2_X1 U740 (.Z( n535 ) , .A( n538 ) , .B( n539 ) );
  XNOR2_X1 U741 (.B( n491 ) , .ZN( n538 ) , .A( sa00_sr_4 ) );
  XOR2_X1 U742 (.A( n233 ) , .Z( n533 ) , .B( w0_20 ) );
  OAI22_X1 U744 (.ZN( N261 ) , .A1( n1213 ) , .B2( n1220 ) , .A2( n540 ) , .B1( n541 ) );
  XOR2_X1 U745 (.Z( n541 ) , .A( n542 ) , .B( n543 ) );
  XOR2_X1 U746 (.Z( n543 ) , .B( n544 ) , .A( sa10_sr_2 ) );
  XOR2_X1 U747 (.Z( n544 ) , .B( sa20_sr_2 ) , .A( w0_19 ) );
  OAI21_X1 U75 (.B1( ld ) , .ZN( n1014 ) , .B2( n73 ) , .A( n74 ) );
  XOR2_X1 U750 (.A( n231 ) , .Z( n540 ) , .B( w0_19 ) );
  OAI22_X1 U752 (.ZN( N260 ) , .A1( n1213 ) , .B2( n1218 ) , .A2( n546 ) , .B1( n547 ) );
  XOR2_X1 U755 (.Z( n550 ) , .B( sa20_sr_1 ) , .A( w0_18 ) );
  XNOR2_X1 U756 (.B( n503 ) , .ZN( n548 ) , .A( sa00_sr_2 ) );
  XOR2_X1 U757 (.A( n229 ) , .Z( n546 ) , .B( w0_18 ) );
  OAI22_X1 U759 (.ZN( N259 ) , .A1( n1109 ) , .B2( n1218 ) , .A2( n551 ) , .B1( n552 ) );
  NAND2_X1 U76 (.A2( ld ) , .ZN( n74 ) , .A1( text_in[36] ) );
  XOR2_X1 U761 (.Z( n554 ) , .B( n555 ) , .A( sa10_sr_0 ) );
  XOR2_X1 U762 (.Z( n555 ) , .B( sa20_sr_0 ) , .A( w0_17 ) );
  XNOR2_X1 U764 (.B( n509 ) , .ZN( n556 ) , .A( sa00_sr_1 ) );
  XOR2_X1 U765 (.A( n227 ) , .Z( n551 ) , .B( w0_17 ) );
  OAI22_X1 U767 (.ZN( N258 ) , .A1( n1109 ) , .B2( n1220 ) , .A2( n557 ) , .B1( n558 ) );
  XOR2_X1 U769 (.A( n516 ) , .B( n539 ) , .Z( n560 ) );
  OAI21_X1 U77 (.B1( ld ) , .ZN( n1015 ) , .B2( n75 ) , .A( n76 ) );
  XOR2_X1 U770 (.Z( n539 ) , .A( sa10_sr_7 ) , .B( sa20_sr_7 ) );
  XOR2_X1 U772 (.A( n225 ) , .Z( n557 ) , .B( w0_16 ) );
  OAI22_X1 U774 (.ZN( N249 ) , .A1( n1109 ) , .B2( n1217 ) , .A2( n561 ) , .B1( n562 ) );
  XOR2_X1 U776 (.A( n476 ) , .B( n488 ) , .Z( n564 ) );
  XOR2_X1 U777 (.Z( n476 ) , .A( sa20_sr_6 ) , .B( sa30_sr_6 ) );
  XOR2_X1 U779 (.A( n223 ) , .Z( n561 ) , .B( w0_15 ) );
  NAND2_X1 U78 (.A2( ld ) , .ZN( n76 ) , .A1( text_in[37] ) );
  OAI22_X1 U781 (.ZN( N248 ) , .A1( n1109 ) , .B2( n1220 ) , .A2( n565 ) , .B1( n566 ) );
  XOR2_X1 U783 (.A( n470 ) , .B( n482 ) , .Z( n568 ) );
  XOR2_X1 U784 (.Z( n482 ) , .A( sa20_sr_5 ) , .B( sa30_sr_5 ) );
  XOR2_X1 U786 (.A( n221 ) , .Z( n565 ) , .B( w0_14 ) );
  OAI22_X1 U788 (.ZN( N247 ) , .A1( n1212 ) , .B2( n1221 ) , .A2( n569 ) , .B1( n570 ) );
  XOR2_X1 U789 (.Z( n570 ) , .A( n571 ) , .B( n572 ) );
  OAI21_X1 U79 (.B1( ld ) , .ZN( n1016 ) , .B2( n77 ) , .A( n78 ) );
  XOR2_X1 U790 (.A( n477 ) , .B( n491 ) , .Z( n572 ) );
  XOR2_X1 U791 (.Z( n491 ) , .A( sa20_sr_4 ) , .B( sa30_sr_4 ) );
  XNOR2_X1 U792 (.ZN( n571 ) , .B( sa30_sr_5 ) , .A( w0_13 ) );
  XOR2_X1 U793 (.A( n219 ) , .Z( n569 ) , .B( w0_13 ) );
  OAI22_X1 U795 (.ZN( N246 ) , .A1( n1213 ) , .B2( n1217 ) , .A2( n573 ) , .B1( n574 ) );
  XOR2_X1 U796 (.Z( n574 ) , .A( n575 ) , .B( n576 ) );
  XOR2_X1 U797 (.A( n483 ) , .B( n496 ) , .Z( n576 ) );
  XOR2_X1 U798 (.Z( n496 ) , .A( sa20_sr_3 ) , .B( sa30_sr_3 ) );
  XOR2_X1 U799 (.B( n469 ) , .Z( n575 ) , .A( n577 ) );
  NAND2_X1 U8 (.A2( ld ) , .ZN( n6 ) , .A1( text_in[2] ) );
  NAND2_X1 U80 (.A2( ld ) , .ZN( n78 ) , .A1( text_in[38] ) );
  XNOR2_X1 U800 (.ZN( n577 ) , .B( sa30_sr_4 ) , .A( w0_12 ) );
  XOR2_X1 U801 (.A( n217 ) , .Z( n573 ) , .B( w0_12 ) );
  OAI22_X1 U803 (.ZN( N245 ) , .B2( n1114 ) , .A1( n1216 ) , .A2( n578 ) , .B1( n579 ) );
  XOR2_X1 U805 (.A( n489 ) , .B( n503 ) , .Z( n581 ) );
  XOR2_X1 U806 (.Z( n503 ) , .A( sa20_sr_2 ) , .B( sa30_sr_2 ) );
  XNOR2_X1 U808 (.ZN( n582 ) , .B( sa30_sr_3 ) , .A( w0_11 ) );
  XOR2_X1 U809 (.A( n215 ) , .Z( n578 ) , .B( w0_11 ) );
  OAI21_X1 U81 (.B1( ld ) , .ZN( n1017 ) , .B2( n79 ) , .A( n80 ) );
  OAI22_X1 U811 (.ZN( N244 ) , .A1( n1212 ) , .B2( n1220 ) , .A2( n583 ) , .B1( n584 ) );
  XOR2_X1 U813 (.A( n497 ) , .B( n509 ) , .Z( n586 ) );
  XOR2_X1 U814 (.Z( n509 ) , .A( sa20_sr_1 ) , .B( sa30_sr_1 ) );
  XOR2_X1 U816 (.A( n213 ) , .Z( n583 ) , .B( w0_10 ) );
  OAI22_X1 U818 (.ZN( N243 ) , .A1( n1212 ) , .B2( n1220 ) , .A2( n587 ) , .B1( n588 ) );
  NAND2_X1 U82 (.A2( ld ) , .ZN( n80 ) , .A1( text_in[39] ) );
  XOR2_X1 U820 (.A( n504 ) , .B( n516 ) , .Z( n590 ) );
  XOR2_X1 U821 (.Z( n516 ) , .A( sa20_sr_0 ) , .B( sa30_sr_0 ) );
  XNOR2_X1 U823 (.ZN( n591 ) , .B( sa30_sr_1 ) , .A( w0_9 ) );
  XOR2_X1 U824 (.A( n211 ) , .Z( n587 ) , .B( w0_9 ) );
  OAI22_X1 U826 (.ZN( N242 ) , .A1( n1215 ) , .B2( n1220 ) , .A2( n592 ) , .B1( n593 ) );
  XOR2_X1 U828 (.A( n469 ) , .B( n510 ) , .Z( n595 ) );
  XOR2_X1 U829 (.Z( n469 ) , .A( sa20_sr_7 ) , .B( sa30_sr_7 ) );
  OAI21_X1 U83 (.B1( ld ) , .ZN( n1018 ) , .B2( n81 ) , .A( n82 ) );
  XOR2_X1 U831 (.A( n209 ) , .Z( n592 ) , .B( w0_8 ) );
  OAI22_X1 U833 (.ZN( N233 ) , .A1( n1213 ) , .B2( n1221 ) , .A2( n596 ) , .B1( n597 ) );
  XOR2_X1 U834 (.Z( n597 ) , .A( n598 ) , .B( n599 ) );
  XOR2_X1 U835 (.B( n488 ) , .Z( n599 ) , .A( sa00_sr_6 ) );
  XOR2_X1 U836 (.Z( n488 ) , .A( sa00_sr_7 ) , .B( sa10_sr_7 ) );
  XNOR2_X1 U837 (.ZN( n598 ) , .B( n600 ) , .A( sa20_sr_7 ) );
  XOR2_X1 U838 (.Z( n600 ) , .B( sa30_sr_6 ) , .A( w0_7 ) );
  XOR2_X1 U839 (.A( n207 ) , .Z( n596 ) , .B( w0_7 ) );
  NAND2_X1 U84 (.A2( ld ) , .ZN( n82 ) , .A1( text_in[40] ) );
  OAI22_X1 U841 (.ZN( N232 ) , .A1( n1109 ) , .B2( n1217 ) , .A2( n601 ) , .B1( n602 ) );
  XOR2_X1 U844 (.Z( n605 ) , .B( sa30_sr_5 ) , .A( w0_6 ) );
  XNOR2_X1 U845 (.B( n470 ) , .ZN( n603 ) , .A( sa00_sr_5 ) );
  XOR2_X1 U846 (.Z( n470 ) , .A( sa00_sr_6 ) , .B( sa10_sr_6 ) );
  XOR2_X1 U847 (.A( n205 ) , .Z( n601 ) , .B( w0_6 ) );
  OAI22_X1 U849 (.ZN( N231 ) , .A1( n1109 ) , .B2( n1217 ) , .A2( n606 ) , .B1( n607 ) );
  OAI21_X1 U85 (.B1( ld ) , .ZN( n1019 ) , .B2( n83 ) , .A( n84 ) );
  XOR2_X1 U850 (.Z( n607 ) , .A( n608 ) , .B( n609 ) );
  XOR2_X1 U851 (.Z( n609 ) , .B( n610 ) , .A( sa20_sr_5 ) );
  XOR2_X1 U852 (.Z( n610 ) , .B( sa30_sr_4 ) , .A( w0_5 ) );
  XNOR2_X1 U853 (.B( n477 ) , .ZN( n608 ) , .A( sa00_sr_4 ) );
  XOR2_X1 U854 (.Z( n477 ) , .A( sa00_sr_5 ) , .B( sa10_sr_5 ) );
  XOR2_X1 U855 (.A( n203 ) , .Z( n606 ) , .B( w0_5 ) );
  OAI22_X1 U857 (.ZN( N230 ) , .A1( n1109 ) , .B2( n1217 ) , .A2( n611 ) , .B1( n612 ) );
  XOR2_X1 U858 (.Z( n612 ) , .A( n613 ) , .B( n614 ) );
  XOR2_X1 U859 (.Z( n614 ) , .B( n615 ) , .A( sa20_sr_4 ) );
  NAND2_X1 U86 (.A2( ld ) , .ZN( n84 ) , .A1( text_in[41] ) );
  XOR2_X1 U860 (.Z( n615 ) , .B( sa30_sr_3 ) , .A( w0_4 ) );
  XOR2_X1 U861 (.Z( n613 ) , .A( n616 ) , .B( n617 ) );
  XNOR2_X1 U862 (.B( n483 ) , .ZN( n616 ) , .A( sa00_sr_3 ) );
  XOR2_X1 U863 (.Z( n483 ) , .A( sa00_sr_4 ) , .B( sa10_sr_4 ) );
  XOR2_X1 U864 (.A( n201 ) , .Z( n611 ) , .B( w0_4 ) );
  NOR4_X1 U866 (.ZN( N23 ) , .A3( ld ) , .A2( n1108 ) , .A4( n260 ) , .A1( n977 ) );
  NAND2_X1 U867 (.A1( n1106 ) , .A2( n1107 ) , .ZN( n260 ) );
  OAI22_X1 U868 (.ZN( N229 ) , .A1( n1109 ) , .B2( n1217 ) , .A2( n618 ) , .B1( n619 ) );
  OAI21_X1 U87 (.B1( ld ) , .ZN( n1020 ) , .B2( n85 ) , .A( n86 ) );
  XOR2_X1 U871 (.Z( n622 ) , .B( sa30_sr_2 ) , .A( w0_3 ) );
  XOR2_X1 U872 (.B( n617 ) , .Z( n620 ) , .A( n623 ) );
  XNOR2_X1 U873 (.B( n489 ) , .ZN( n623 ) , .A( sa00_sr_2 ) );
  XOR2_X1 U874 (.Z( n489 ) , .A( sa00_sr_3 ) , .B( sa10_sr_3 ) );
  XOR2_X1 U875 (.A( n199 ) , .Z( n618 ) , .B( w0_3 ) );
  OAI22_X1 U877 (.ZN( N228 ) , .A1( n1109 ) , .B2( n1217 ) , .A2( n624 ) , .B1( n625 ) );
  NAND2_X1 U88 (.A2( ld ) , .ZN( n86 ) , .A1( text_in[42] ) );
  XOR2_X1 U880 (.Z( n628 ) , .B( sa30_sr_1 ) , .A( w0_2 ) );
  XNOR2_X1 U881 (.B( n497 ) , .ZN( n626 ) , .A( sa00_sr_1 ) );
  XOR2_X1 U882 (.Z( n497 ) , .A( sa00_sr_2 ) , .B( sa10_sr_2 ) );
  XOR2_X1 U883 (.A( n197 ) , .Z( n624 ) , .B( w0_2 ) );
  OAI22_X1 U885 (.ZN( N227 ) , .A1( n1109 ) , .B2( n1217 ) , .A2( n629 ) , .B1( n630 ) );
  XOR2_X1 U887 (.Z( n632 ) , .B( n633 ) , .A( sa20_sr_1 ) );
  XOR2_X1 U888 (.Z( n633 ) , .B( sa30_sr_0 ) , .A( w0_1 ) );
  OAI21_X1 U89 (.B1( ld ) , .ZN( n1021 ) , .B2( n87 ) , .A( n88 ) );
  XNOR2_X1 U890 (.B( n504 ) , .ZN( n634 ) , .A( sa00_sr_0 ) );
  XOR2_X1 U891 (.Z( n504 ) , .A( sa00_sr_1 ) , .B( sa10_sr_1 ) );
  XOR2_X1 U892 (.A( n195 ) , .Z( n629 ) , .B( w0_1 ) );
  OAI22_X1 U894 (.ZN( N226 ) , .A1( n1109 ) , .B2( n1217 ) , .A2( n635 ) , .B1( n636 ) );
  XOR2_X1 U896 (.A( n510 ) , .B( n617 ) , .Z( n638 ) );
  XOR2_X1 U897 (.Z( n617 ) , .A( sa00_sr_7 ) , .B( sa30_sr_7 ) );
  XOR2_X1 U898 (.Z( n510 ) , .A( sa00_sr_0 ) , .B( sa10_sr_0 ) );
  OAI21_X1 U9 (.B1( ld ) , .B2( n7 ) , .A( n8 ) , .ZN( n981 ) );
  NAND2_X1 U90 (.A2( ld ) , .ZN( n88 ) , .A1( text_in[43] ) );
  XOR2_X1 U900 (.A( n193 ) , .Z( n635 ) , .B( w0_0 ) );
  OAI22_X1 U902 (.ZN( N217 ) , .A1( n1109 ) , .B2( n1218 ) , .A2( n639 ) , .B1( n640 ) );
  XOR2_X1 U904 (.Z( n642 ) , .A( n643 ) , .B( n644 ) );
  INV_X1 U906 (.ZN( n645 ) , .A( sa11_sr_7 ) );
  XOR2_X1 U907 (.A( n191 ) , .Z( n639 ) , .B( w1_31 ) );
  OAI22_X1 U909 (.ZN( N216 ) , .A1( n1109 ) , .B2( n1218 ) , .A2( n646 ) , .B1( n647 ) );
  OAI21_X1 U91 (.B1( ld ) , .ZN( n1022 ) , .B2( n89 ) , .A( n90 ) );
  XOR2_X1 U911 (.Z( n649 ) , .A( n650 ) , .B( n651 ) );
  XOR2_X1 U913 (.A( n189 ) , .Z( n646 ) , .B( w1_30 ) );
  OAI22_X1 U915 (.ZN( N215 ) , .A1( n1109 ) , .B2( n1218 ) , .A2( n652 ) , .B1( n653 ) );
  XOR2_X1 U917 (.Z( n655 ) , .A( n656 ) , .B( n657 ) );
  XOR2_X1 U919 (.A( n187 ) , .Z( n652 ) , .B( w1_29 ) );
  NAND2_X1 U92 (.A2( ld ) , .ZN( n90 ) , .A1( text_in[44] ) );
  OAI22_X1 U921 (.ZN( N214 ) , .A1( n1109 ) , .B2( n1218 ) , .A2( n658 ) , .B1( n659 ) );
  XOR2_X1 U922 (.Z( n659 ) , .A( n660 ) , .B( n661 ) );
  XOR2_X1 U923 (.Z( n661 ) , .A( n662 ) , .B( n663 ) );
  XOR2_X1 U924 (.Z( n660 ) , .A( n664 ) , .B( n665 ) );
  XNOR2_X1 U925 (.ZN( n664 ) , .B( sa11_sr_4 ) , .A( w1_28 ) );
  XOR2_X1 U926 (.A( n185 ) , .Z( n658 ) , .B( w1_28 ) );
  OAI22_X1 U928 (.ZN( N213 ) , .A1( n1213 ) , .B2( n1218 ) , .A2( n666 ) , .B1( n667 ) );
  OAI21_X1 U93 (.B1( ld ) , .ZN( n1023 ) , .B2( n91 ) , .A( n92 ) );
  XOR2_X1 U930 (.Z( n669 ) , .A( n670 ) , .B( n671 ) );
  XNOR2_X1 U932 (.ZN( n672 ) , .B( sa11_sr_3 ) , .A( w1_27 ) );
  XOR2_X1 U933 (.A( n183 ) , .Z( n666 ) , .B( w1_27 ) );
  OAI22_X1 U935 (.ZN( N212 ) , .A1( n1214 ) , .B2( n1218 ) , .A2( n673 ) , .B1( n674 ) );
  XOR2_X1 U937 (.Z( n676 ) , .A( n677 ) , .B( n678 ) );
  XOR2_X1 U939 (.A( n181 ) , .Z( n673 ) , .B( w1_26 ) );
  NAND2_X1 U94 (.A2( ld ) , .ZN( n92 ) , .A1( text_in[45] ) );
  OAI22_X1 U941 (.ZN( N211 ) , .A1( n1214 ) , .B2( n1218 ) , .A2( n679 ) , .B1( n680 ) );
  XOR2_X1 U943 (.Z( n682 ) , .A( n683 ) , .B( n684 ) );
  XNOR2_X1 U945 (.ZN( n685 ) , .B( sa11_sr_1 ) , .A( w1_25 ) );
  XOR2_X1 U946 (.A( n179 ) , .Z( n679 ) , .B( w1_25 ) );
  OAI22_X1 U948 (.ZN( N210 ) , .A1( n1109 ) , .B2( n1219 ) , .A2( n686 ) , .B1( n687 ) );
  OAI21_X1 U95 (.B1( ld ) , .ZN( n1024 ) , .B2( n93 ) , .A( n94 ) );
  XOR2_X1 U950 (.A( n665 ) , .Z( n689 ) , .B( n690 ) );
  XOR2_X1 U952 (.A( n177 ) , .Z( n686 ) , .B( w1_24 ) );
  OAI22_X1 U954 (.ZN( N201 ) , .A1( n1214 ) , .B2( n1217 ) , .A2( n691 ) , .B1( n692 ) );
  XOR2_X1 U955 (.Z( n692 ) , .A( n693 ) , .B( n694 ) );
  XOR2_X1 U956 (.B( n643 ) , .Z( n694 ) , .A( sa01_sr_7 ) );
  XOR2_X1 U959 (.A( n175 ) , .Z( n691 ) , .B( w1_23 ) );
  NAND2_X1 U96 (.A2( ld ) , .ZN( n94 ) , .A1( text_in[46] ) );
  OAI22_X1 U961 (.ZN( N200 ) , .A1( n1212 ) , .B2( n1219 ) , .A2( n696 ) , .B1( n697 ) );
  XOR2_X1 U964 (.Z( n700 ) , .B( sa21_sr_5 ) , .A( w1_22 ) );
  XOR2_X1 U967 (.A( n173 ) , .Z( n696 ) , .B( w1_22 ) );
  OAI22_X1 U969 (.ZN( N199 ) , .A1( n1215 ) , .B2( n1218 ) , .A2( n702 ) , .B1( n703 ) );
  OAI21_X1 U97 (.B1( ld ) , .ZN( n1025 ) , .B2( n95 ) , .A( n96 ) );
  XOR2_X1 U970 (.Z( n703 ) , .A( n704 ) , .B( n705 ) );
  XOR2_X1 U971 (.Z( n705 ) , .B( n706 ) , .A( sa11_sr_4 ) );
  XOR2_X1 U972 (.Z( n706 ) , .B( sa21_sr_4 ) , .A( w1_21 ) );
  XNOR2_X1 U973 (.B( n656 ) , .ZN( n704 ) , .A( sa01_sr_5 ) );
  XOR2_X1 U974 (.A( n171 ) , .Z( n702 ) , .B( w1_21 ) );
  OAI22_X1 U976 (.ZN( N198 ) , .A1( n1216 ) , .B2( n1217 ) , .A2( n707 ) , .B1( n708 ) );
  XOR2_X1 U977 (.Z( n708 ) , .A( n709 ) , .B( n710 ) );
  XOR2_X1 U978 (.Z( n710 ) , .B( n711 ) , .A( sa11_sr_3 ) );
  XOR2_X1 U979 (.Z( n711 ) , .B( sa21_sr_3 ) , .A( w1_20 ) );
  NAND2_X1 U98 (.A2( ld ) , .ZN( n96 ) , .A1( text_in[47] ) );
  XOR2_X1 U980 (.Z( n709 ) , .A( n712 ) , .B( n713 ) );
  XNOR2_X1 U981 (.B( n663 ) , .ZN( n712 ) , .A( sa01_sr_4 ) );
  XOR2_X1 U982 (.A( n169 ) , .Z( n707 ) , .B( w1_20 ) );
  OAI22_X1 U984 (.ZN( N197 ) , .A1( n1109 ) , .B2( n1220 ) , .A2( n714 ) , .B1( n715 ) );
  XOR2_X1 U987 (.Z( n718 ) , .B( sa21_sr_2 ) , .A( w1_19 ) );
  XOR2_X1 U988 (.B( n713 ) , .Z( n716 ) , .A( n719 ) );
  XNOR2_X1 U989 (.B( n670 ) , .ZN( n719 ) , .A( sa01_sr_3 ) );
  OAI21_X1 U99 (.B1( ld ) , .ZN( n1026 ) , .B2( n97 ) , .A( n98 ) );
  XOR2_X1 U990 (.A( n167 ) , .Z( n714 ) , .B( w1_19 ) );
  OAI22_X1 U992 (.ZN( N196 ) , .A1( n1212 ) , .B2( n1218 ) , .A2( n720 ) , .B1( n721 ) );
  XOR2_X1 U995 (.Z( n724 ) , .B( sa21_sr_1 ) , .A( w1_18 ) );
  XNOR2_X1 U996 (.B( n677 ) , .ZN( n722 ) , .A( sa01_sr_2 ) );
  XOR2_X1 U997 (.A( n165 ) , .Z( n720 ) , .B( w1_18 ) );
  OAI22_X1 U999 (.ZN( N195 ) , .A1( n1215 ) , .B2( n1221 ) , .A2( n725 ) , .B1( n726 ) );
  DFF_X1 dcnt_reg_0 (.CK( clk ) , .QN( n1108 ) , .D( n1113 ) , .Q( n261 ) );
  DFF_X1 dcnt_reg_1 (.CK( clk ) , .D( n1110 ) , .Q( n977 ) );
  DFF_X1 dcnt_reg_2 (.CK( clk ) , .QN( n1107 ) , .D( n1111 ) , .Q( n267 ) );
  DFF_X1 dcnt_reg_3 (.CK( clk ) , .QN( n1106 ) , .D( n1112 ) );
  DFF_X1 done_reg (.D( N23 ) , .CK( clk ) , .Q( done ) );
  DFF_X1 ld_r_reg (.CK( clk ) , .D( ld ) , .QN( n1109 ) , .Q( n1114 ) );
  DFF_X1 sa00_reg_0 (.D( N274 ) , .CK( clk ) , .Q( sa00_0 ) );
  DFF_X1 sa00_reg_1 (.D( N275 ) , .CK( clk ) , .Q( sa00_1 ) );
  DFF_X1 sa00_reg_2 (.D( N276 ) , .CK( clk ) , .Q( sa00_2 ) );
  DFF_X1 sa00_reg_3 (.D( N277 ) , .CK( clk ) , .Q( sa00_3 ) );
  DFF_X1 sa00_reg_4 (.D( N278 ) , .CK( clk ) , .Q( sa00_4 ) );
  DFF_X1 sa00_reg_5 (.D( N279 ) , .CK( clk ) , .Q( sa00_5 ) );
  DFF_X1 sa00_reg_6 (.D( N280 ) , .CK( clk ) , .Q( sa00_6 ) );
  DFF_X1 sa00_reg_7 (.D( N281 ) , .CK( clk ) , .Q( sa00_7 ) );
  DFF_X1 sa01_reg_0 (.D( N210 ) , .CK( clk ) , .Q( sa01_0 ) );
  DFF_X1 sa01_reg_1 (.D( N211 ) , .CK( clk ) , .Q( sa01_1 ) );
  DFF_X1 sa01_reg_2 (.D( N212 ) , .CK( clk ) , .Q( sa01_2 ) );
  DFF_X1 sa01_reg_3 (.D( N213 ) , .CK( clk ) , .Q( sa01_3 ) );
  DFF_X1 sa01_reg_4 (.D( N214 ) , .CK( clk ) , .Q( sa01_4 ) );
  DFF_X1 sa01_reg_5 (.D( N215 ) , .CK( clk ) , .Q( sa01_5 ) );
  DFF_X1 sa01_reg_6 (.D( N216 ) , .CK( clk ) , .Q( sa01_6 ) );
  DFF_X1 sa01_reg_7 (.D( N217 ) , .CK( clk ) , .Q( sa01_7 ) );
  DFF_X1 sa02_reg_0 (.D( N146 ) , .CK( clk ) , .Q( sa02_0 ) );
  DFF_X1 sa02_reg_1 (.D( N147 ) , .CK( clk ) , .Q( sa02_1 ) );
  DFF_X1 sa02_reg_2 (.D( N148 ) , .CK( clk ) , .Q( sa02_2 ) );
  DFF_X1 sa02_reg_3 (.D( N149 ) , .CK( clk ) , .Q( sa02_3 ) );
  DFF_X1 sa02_reg_4 (.D( N150 ) , .CK( clk ) , .Q( sa02_4 ) );
  DFF_X1 sa02_reg_5 (.D( N151 ) , .CK( clk ) , .Q( sa02_5 ) );
  DFF_X1 sa02_reg_6 (.D( N152 ) , .CK( clk ) , .Q( sa02_6 ) );
  DFF_X1 sa02_reg_7 (.D( N153 ) , .CK( clk ) , .Q( sa02_7 ) );
  DFF_X1 sa03_reg_0 (.D( N82 ) , .CK( clk ) , .Q( sa03_0 ) );
  DFF_X1 sa03_reg_1 (.D( N83 ) , .CK( clk ) , .Q( sa03_1 ) );
  DFF_X1 sa03_reg_2 (.D( N84 ) , .CK( clk ) , .Q( sa03_2 ) );
  DFF_X1 sa03_reg_3 (.D( N85 ) , .CK( clk ) , .Q( sa03_3 ) );
  DFF_X1 sa03_reg_4 (.D( N86 ) , .CK( clk ) , .Q( sa03_4 ) );
  DFF_X1 sa03_reg_5 (.D( N87 ) , .CK( clk ) , .Q( sa03_5 ) );
  DFF_X1 sa03_reg_6 (.D( N88 ) , .CK( clk ) , .Q( sa03_6 ) );
  DFF_X1 sa03_reg_7 (.D( N89 ) , .CK( clk ) , .Q( sa03_7 ) );
  DFF_X1 sa10_reg_0 (.D( N258 ) , .CK( clk ) , .Q( sa10_0 ) );
  DFF_X1 sa10_reg_1 (.D( N259 ) , .CK( clk ) , .Q( sa10_1 ) );
  DFF_X1 sa10_reg_2 (.D( N260 ) , .CK( clk ) , .Q( sa10_2 ) );
  DFF_X1 sa10_reg_3 (.D( N261 ) , .CK( clk ) , .Q( sa10_3 ) );
  DFF_X1 sa10_reg_4 (.D( N262 ) , .CK( clk ) , .Q( sa10_4 ) );
  DFF_X1 sa10_reg_5 (.D( N263 ) , .CK( clk ) , .Q( sa10_5 ) );
  DFF_X1 sa10_reg_6 (.D( N264 ) , .CK( clk ) , .Q( sa10_6 ) );
  DFF_X1 sa10_reg_7 (.D( N265 ) , .CK( clk ) , .Q( sa10_7 ) );
  DFF_X1 sa11_reg_0 (.D( N194 ) , .CK( clk ) , .Q( sa11_0 ) );
  DFF_X1 sa11_reg_1 (.D( N195 ) , .CK( clk ) , .Q( sa11_1 ) );
  DFF_X1 sa11_reg_2 (.D( N196 ) , .CK( clk ) , .Q( sa11_2 ) );
  DFF_X1 sa11_reg_3 (.D( N197 ) , .CK( clk ) , .Q( sa11_3 ) );
  DFF_X1 sa11_reg_4 (.D( N198 ) , .CK( clk ) , .Q( sa11_4 ) );
  DFF_X1 sa11_reg_5 (.D( N199 ) , .CK( clk ) , .Q( sa11_5 ) );
  DFF_X1 sa11_reg_6 (.D( N200 ) , .CK( clk ) , .Q( sa11_6 ) );
  DFF_X1 sa11_reg_7 (.D( N201 ) , .CK( clk ) , .Q( sa11_7 ) );
  DFF_X1 sa12_reg_0 (.D( N130 ) , .CK( clk ) , .Q( sa12_0 ) );
  DFF_X1 sa12_reg_1 (.D( N131 ) , .CK( clk ) , .Q( sa12_1 ) );
  DFF_X1 sa12_reg_2 (.D( N132 ) , .CK( clk ) , .Q( sa12_2 ) );
  DFF_X1 sa12_reg_3 (.D( N133 ) , .CK( clk ) , .Q( sa12_3 ) );
  DFF_X1 sa12_reg_4 (.D( N134 ) , .CK( clk ) , .Q( sa12_4 ) );
  DFF_X1 sa12_reg_5 (.D( N135 ) , .CK( clk ) , .Q( sa12_5 ) );
  DFF_X1 sa12_reg_6 (.D( N136 ) , .CK( clk ) , .Q( sa12_6 ) );
  DFF_X1 sa12_reg_7 (.D( N137 ) , .CK( clk ) , .Q( sa12_7 ) );
  DFF_X1 sa13_reg_0 (.D( N66 ) , .CK( clk ) , .Q( sa13_0 ) );
  DFF_X1 sa13_reg_1 (.D( N67 ) , .CK( clk ) , .Q( sa13_1 ) );
  DFF_X1 sa13_reg_2 (.D( N68 ) , .CK( clk ) , .Q( sa13_2 ) );
  DFF_X1 sa13_reg_3 (.D( N69 ) , .CK( clk ) , .Q( sa13_3 ) );
  DFF_X1 sa13_reg_4 (.D( N70 ) , .CK( clk ) , .Q( sa13_4 ) );
  DFF_X1 sa13_reg_5 (.D( N71 ) , .CK( clk ) , .Q( sa13_5 ) );
  DFF_X1 sa13_reg_6 (.D( N72 ) , .CK( clk ) , .Q( sa13_6 ) );
  DFF_X1 sa13_reg_7 (.D( N73 ) , .CK( clk ) , .Q( sa13_7 ) );
  DFF_X1 sa20_reg_0 (.D( N242 ) , .CK( clk ) , .Q( sa20_0 ) );
  DFF_X1 sa20_reg_1 (.D( N243 ) , .CK( clk ) , .Q( sa20_1 ) );
  DFF_X1 sa20_reg_2 (.D( N244 ) , .CK( clk ) , .Q( sa20_2 ) );
  DFF_X1 sa20_reg_3 (.D( N245 ) , .CK( clk ) , .Q( sa20_3 ) );
  DFF_X1 sa20_reg_4 (.D( N246 ) , .CK( clk ) , .Q( sa20_4 ) );
  DFF_X1 sa20_reg_5 (.D( N247 ) , .CK( clk ) , .Q( sa20_5 ) );
  DFF_X1 sa20_reg_6 (.D( N248 ) , .CK( clk ) , .Q( sa20_6 ) );
  DFF_X1 sa20_reg_7 (.D( N249 ) , .CK( clk ) , .Q( sa20_7 ) );
  DFF_X1 sa21_reg_0 (.D( N178 ) , .CK( clk ) , .Q( sa21_0 ) );
  DFF_X1 sa21_reg_1 (.D( N179 ) , .CK( clk ) , .Q( sa21_1 ) );
  DFF_X1 sa21_reg_2 (.D( N180 ) , .CK( clk ) , .Q( sa21_2 ) );
  DFF_X1 sa21_reg_3 (.D( N181 ) , .CK( clk ) , .Q( sa21_3 ) );
  DFF_X1 sa21_reg_4 (.D( N182 ) , .CK( clk ) , .Q( sa21_4 ) );
  DFF_X1 sa21_reg_5 (.D( N183 ) , .CK( clk ) , .Q( sa21_5 ) );
  DFF_X1 sa21_reg_6 (.D( N184 ) , .CK( clk ) , .Q( sa21_6 ) );
  DFF_X1 sa21_reg_7 (.D( N185 ) , .CK( clk ) , .Q( sa21_7 ) );
  DFF_X1 sa22_reg_0 (.D( N114 ) , .CK( clk ) , .Q( sa22_0 ) );
  DFF_X1 sa22_reg_1 (.D( N115 ) , .CK( clk ) , .Q( sa22_1 ) );
  DFF_X1 sa22_reg_2 (.D( N116 ) , .CK( clk ) , .Q( sa22_2 ) );
  DFF_X1 sa22_reg_3 (.D( N117 ) , .CK( clk ) , .Q( sa22_3 ) );
  DFF_X1 sa22_reg_4 (.D( N118 ) , .CK( clk ) , .Q( sa22_4 ) );
  DFF_X1 sa22_reg_5 (.D( N119 ) , .CK( clk ) , .Q( sa22_5 ) );
  DFF_X1 sa22_reg_6 (.D( N120 ) , .CK( clk ) , .Q( sa22_6 ) );
  DFF_X1 sa22_reg_7 (.D( N121 ) , .CK( clk ) , .Q( sa22_7 ) );
  DFF_X1 sa23_reg_0 (.D( N50 ) , .CK( clk ) , .Q( sa23_0 ) );
  DFF_X1 sa23_reg_1 (.D( N51 ) , .CK( clk ) , .Q( sa23_1 ) );
  DFF_X1 sa23_reg_2 (.D( N52 ) , .CK( clk ) , .Q( sa23_2 ) );
  DFF_X1 sa23_reg_3 (.D( N53 ) , .CK( clk ) , .Q( sa23_3 ) );
  DFF_X1 sa23_reg_4 (.D( N54 ) , .CK( clk ) , .Q( sa23_4 ) );
  DFF_X1 sa23_reg_5 (.D( N55 ) , .CK( clk ) , .Q( sa23_5 ) );
  DFF_X1 sa23_reg_6 (.D( N56 ) , .CK( clk ) , .Q( sa23_6 ) );
  DFF_X1 sa23_reg_7 (.D( N57 ) , .CK( clk ) , .Q( sa23_7 ) );
  DFF_X1 sa30_reg_0 (.D( N226 ) , .CK( clk ) , .Q( sa30_0 ) );
  DFF_X1 sa30_reg_1 (.D( N227 ) , .CK( clk ) , .Q( sa30_1 ) );
  DFF_X1 sa30_reg_2 (.D( N228 ) , .CK( clk ) , .Q( sa30_2 ) );
  DFF_X1 sa30_reg_3 (.D( N229 ) , .CK( clk ) , .Q( sa30_3 ) );
  DFF_X1 sa30_reg_4 (.D( N230 ) , .CK( clk ) , .Q( sa30_4 ) );
  DFF_X1 sa30_reg_5 (.D( N231 ) , .CK( clk ) , .Q( sa30_5 ) );
  DFF_X1 sa30_reg_6 (.D( N232 ) , .CK( clk ) , .Q( sa30_6 ) );
  DFF_X1 sa30_reg_7 (.D( N233 ) , .CK( clk ) , .Q( sa30_7 ) );
  DFF_X1 sa31_reg_0 (.D( N162 ) , .CK( clk ) , .Q( sa31_0 ) );
  DFF_X1 sa31_reg_1 (.D( N163 ) , .CK( clk ) , .Q( sa31_1 ) );
  DFF_X1 sa31_reg_2 (.D( N164 ) , .CK( clk ) , .Q( sa31_2 ) );
  DFF_X1 sa31_reg_3 (.D( N165 ) , .CK( clk ) , .Q( sa31_3 ) );
  DFF_X1 sa31_reg_4 (.D( N166 ) , .CK( clk ) , .Q( sa31_4 ) );
  DFF_X1 sa31_reg_5 (.D( N167 ) , .CK( clk ) , .Q( sa31_5 ) );
  DFF_X1 sa31_reg_6 (.D( N168 ) , .CK( clk ) , .Q( sa31_6 ) );
  DFF_X1 sa31_reg_7 (.D( N169 ) , .CK( clk ) , .Q( sa31_7 ) );
  DFF_X1 sa32_reg_0 (.D( N98 ) , .CK( clk ) , .Q( sa32_0 ) );
  DFF_X1 sa32_reg_1 (.D( N99 ) , .CK( clk ) , .Q( sa32_1 ) );
  DFF_X1 sa32_reg_2 (.D( N100 ) , .CK( clk ) , .Q( sa32_2 ) );
  DFF_X1 sa32_reg_3 (.D( N101 ) , .CK( clk ) , .Q( sa32_3 ) );
  DFF_X1 sa32_reg_4 (.D( N102 ) , .CK( clk ) , .Q( sa32_4 ) );
  DFF_X1 sa32_reg_5 (.D( N103 ) , .CK( clk ) , .Q( sa32_5 ) );
  DFF_X1 sa32_reg_6 (.D( N104 ) , .CK( clk ) , .Q( sa32_6 ) );
  DFF_X1 sa32_reg_7 (.D( N105 ) , .CK( clk ) , .Q( sa32_7 ) );
  DFF_X1 sa33_reg_0 (.D( N34 ) , .CK( clk ) , .Q( sa33_0 ) );
  DFF_X1 sa33_reg_1 (.D( N35 ) , .CK( clk ) , .Q( sa33_1 ) );
  DFF_X1 sa33_reg_2 (.D( N36 ) , .CK( clk ) , .Q( sa33_2 ) );
  DFF_X1 sa33_reg_3 (.D( N37 ) , .CK( clk ) , .Q( sa33_3 ) );
  DFF_X1 sa33_reg_4 (.D( N38 ) , .CK( clk ) , .Q( sa33_4 ) );
  DFF_X1 sa33_reg_5 (.D( N39 ) , .CK( clk ) , .Q( sa33_5 ) );
  DFF_X1 sa33_reg_6 (.D( N40 ) , .CK( clk ) , .Q( sa33_6 ) );
  DFF_X1 sa33_reg_7 (.D( N41 ) , .CK( clk ) , .Q( sa33_7 ) );
  DFF_X1 text_in_r_reg_0 (.CK( clk ) , .QN( n1 ) , .D( n978 ) );
  DFF_X1 text_in_r_reg_1 (.CK( clk ) , .QN( n3 ) , .D( n979 ) );
  DFF_X1 text_in_r_reg_10 (.CK( clk ) , .QN( n21 ) , .D( n988 ) );
  DFF_X1 text_in_r_reg_100 (.CK( clk ) , .D( n1078 ) , .QN( n201 ) );
  DFF_X1 text_in_r_reg_101 (.CK( clk ) , .D( n1079 ) , .QN( n203 ) );
  DFF_X1 text_in_r_reg_102 (.CK( clk ) , .D( n1080 ) , .QN( n205 ) );
  DFF_X1 text_in_r_reg_103 (.CK( clk ) , .D( n1081 ) , .QN( n207 ) );
  DFF_X1 text_in_r_reg_104 (.CK( clk ) , .D( n1082 ) , .QN( n209 ) );
  DFF_X1 text_in_r_reg_105 (.CK( clk ) , .D( n1083 ) , .QN( n211 ) );
  DFF_X1 text_in_r_reg_106 (.CK( clk ) , .D( n1084 ) , .QN( n213 ) );
  DFF_X1 text_in_r_reg_107 (.CK( clk ) , .D( n1085 ) , .QN( n215 ) );
  DFF_X1 text_in_r_reg_108 (.CK( clk ) , .D( n1086 ) , .QN( n217 ) );
  DFF_X1 text_in_r_reg_109 (.CK( clk ) , .D( n1087 ) , .QN( n219 ) );
  DFF_X1 text_in_r_reg_11 (.CK( clk ) , .QN( n23 ) , .D( n989 ) );
  DFF_X1 text_in_r_reg_110 (.CK( clk ) , .D( n1088 ) , .QN( n221 ) );
  DFF_X1 text_in_r_reg_111 (.CK( clk ) , .D( n1089 ) , .QN( n223 ) );
  DFF_X1 text_in_r_reg_112 (.CK( clk ) , .D( n1090 ) , .QN( n225 ) );
  DFF_X1 text_in_r_reg_113 (.CK( clk ) , .D( n1091 ) , .QN( n227 ) );
  DFF_X1 text_in_r_reg_114 (.CK( clk ) , .D( n1092 ) , .QN( n229 ) );
  DFF_X1 text_in_r_reg_115 (.CK( clk ) , .D( n1093 ) , .QN( n231 ) );
  DFF_X1 text_in_r_reg_116 (.CK( clk ) , .D( n1094 ) , .QN( n233 ) );
  DFF_X1 text_in_r_reg_117 (.CK( clk ) , .D( n1095 ) , .QN( n235 ) );
  DFF_X1 text_in_r_reg_118 (.CK( clk ) , .D( n1096 ) , .QN( n237 ) );
  DFF_X1 text_in_r_reg_119 (.CK( clk ) , .D( n1097 ) , .QN( n239 ) );
  DFF_X1 text_in_r_reg_12 (.CK( clk ) , .QN( n25 ) , .D( n990 ) );
  DFF_X1 text_in_r_reg_120 (.CK( clk ) , .D( n1098 ) , .QN( n241 ) );
  DFF_X1 text_in_r_reg_121 (.CK( clk ) , .D( n1099 ) , .QN( n243 ) );
  DFF_X1 text_in_r_reg_122 (.CK( clk ) , .D( n1100 ) , .QN( n245 ) );
  DFF_X1 text_in_r_reg_123 (.CK( clk ) , .D( n1101 ) , .QN( n247 ) );
  DFF_X1 text_in_r_reg_124 (.CK( clk ) , .D( n1102 ) , .QN( n249 ) );
  DFF_X1 text_in_r_reg_125 (.CK( clk ) , .D( n1103 ) , .QN( n251 ) );
  DFF_X1 text_in_r_reg_126 (.CK( clk ) , .D( n1104 ) , .QN( n253 ) );
  DFF_X1 text_in_r_reg_127 (.CK( clk ) , .D( n1105 ) , .QN( n255 ) );
  DFF_X1 text_in_r_reg_13 (.CK( clk ) , .QN( n27 ) , .D( n991 ) );
  DFF_X1 text_in_r_reg_14 (.CK( clk ) , .QN( n29 ) , .D( n992 ) );
  DFF_X1 text_in_r_reg_15 (.CK( clk ) , .QN( n31 ) , .D( n993 ) );
  DFF_X1 text_in_r_reg_16 (.CK( clk ) , .QN( n33 ) , .D( n994 ) );
  DFF_X1 text_in_r_reg_17 (.CK( clk ) , .QN( n35 ) , .D( n995 ) );
  DFF_X1 text_in_r_reg_18 (.CK( clk ) , .QN( n37 ) , .D( n996 ) );
  DFF_X1 text_in_r_reg_19 (.CK( clk ) , .QN( n39 ) , .D( n997 ) );
  DFF_X1 text_in_r_reg_2 (.CK( clk ) , .QN( n5 ) , .D( n980 ) );
  DFF_X1 text_in_r_reg_20 (.CK( clk ) , .QN( n41 ) , .D( n998 ) );
  DFF_X1 text_in_r_reg_21 (.CK( clk ) , .QN( n43 ) , .D( n999 ) );
  DFF_X1 text_in_r_reg_22 (.CK( clk ) , .D( n1000 ) , .QN( n45 ) );
  DFF_X1 text_in_r_reg_23 (.CK( clk ) , .D( n1001 ) , .QN( n47 ) );
  DFF_X1 text_in_r_reg_24 (.CK( clk ) , .D( n1002 ) , .QN( n49 ) );
  DFF_X1 text_in_r_reg_25 (.CK( clk ) , .D( n1003 ) , .QN( n51 ) );
  DFF_X1 text_in_r_reg_26 (.CK( clk ) , .D( n1004 ) , .QN( n53 ) );
  DFF_X1 text_in_r_reg_27 (.CK( clk ) , .D( n1005 ) , .QN( n55 ) );
  DFF_X1 text_in_r_reg_28 (.CK( clk ) , .D( n1006 ) , .QN( n57 ) );
  DFF_X1 text_in_r_reg_29 (.CK( clk ) , .D( n1007 ) , .QN( n59 ) );
  DFF_X1 text_in_r_reg_3 (.CK( clk ) , .QN( n7 ) , .D( n981 ) );
  DFF_X1 text_in_r_reg_30 (.CK( clk ) , .D( n1008 ) , .QN( n61 ) );
  DFF_X1 text_in_r_reg_31 (.CK( clk ) , .D( n1009 ) , .QN( n63 ) );
  DFF_X1 text_in_r_reg_32 (.CK( clk ) , .D( n1010 ) , .QN( n65 ) );
  DFF_X1 text_in_r_reg_33 (.CK( clk ) , .D( n1011 ) , .QN( n67 ) );
  DFF_X1 text_in_r_reg_34 (.CK( clk ) , .D( n1012 ) , .QN( n69 ) );
  DFF_X1 text_in_r_reg_35 (.CK( clk ) , .D( n1013 ) , .QN( n71 ) );
  DFF_X1 text_in_r_reg_36 (.CK( clk ) , .D( n1014 ) , .QN( n73 ) );
  DFF_X1 text_in_r_reg_37 (.CK( clk ) , .D( n1015 ) , .QN( n75 ) );
  DFF_X1 text_in_r_reg_38 (.CK( clk ) , .D( n1016 ) , .QN( n77 ) );
  DFF_X1 text_in_r_reg_39 (.CK( clk ) , .D( n1017 ) , .QN( n79 ) );
  DFF_X1 text_in_r_reg_4 (.CK( clk ) , .QN( n9 ) , .D( n982 ) );
  DFF_X1 text_in_r_reg_40 (.CK( clk ) , .D( n1018 ) , .QN( n81 ) );
  DFF_X1 text_in_r_reg_41 (.CK( clk ) , .D( n1019 ) , .QN( n83 ) );
  DFF_X1 text_in_r_reg_42 (.CK( clk ) , .D( n1020 ) , .QN( n85 ) );
  DFF_X1 text_in_r_reg_43 (.CK( clk ) , .D( n1021 ) , .QN( n87 ) );
  DFF_X1 text_in_r_reg_44 (.CK( clk ) , .D( n1022 ) , .QN( n89 ) );
  DFF_X1 text_in_r_reg_45 (.CK( clk ) , .D( n1023 ) , .QN( n91 ) );
  DFF_X1 text_in_r_reg_46 (.CK( clk ) , .D( n1024 ) , .QN( n93 ) );
  DFF_X1 text_in_r_reg_47 (.CK( clk ) , .D( n1025 ) , .QN( n95 ) );
  DFF_X1 text_in_r_reg_48 (.CK( clk ) , .D( n1026 ) , .QN( n97 ) );
  DFF_X1 text_in_r_reg_49 (.CK( clk ) , .D( n1027 ) , .QN( n99 ) );
  DFF_X1 text_in_r_reg_5 (.CK( clk ) , .QN( n11 ) , .D( n983 ) );
  DFF_X1 text_in_r_reg_50 (.CK( clk ) , .QN( n101 ) , .D( n1028 ) );
  DFF_X1 text_in_r_reg_51 (.CK( clk ) , .D( n1029 ) , .QN( n103 ) );
  DFF_X1 text_in_r_reg_52 (.CK( clk ) , .D( n1030 ) , .QN( n105 ) );
  DFF_X1 text_in_r_reg_53 (.CK( clk ) , .D( n1031 ) , .QN( n107 ) );
  DFF_X1 text_in_r_reg_54 (.CK( clk ) , .D( n1032 ) , .QN( n109 ) );
  DFF_X1 text_in_r_reg_55 (.CK( clk ) , .D( n1033 ) , .QN( n111 ) );
  DFF_X1 text_in_r_reg_56 (.CK( clk ) , .D( n1034 ) , .QN( n113 ) );
  DFF_X1 text_in_r_reg_57 (.CK( clk ) , .D( n1035 ) , .QN( n115 ) );
  DFF_X1 text_in_r_reg_58 (.CK( clk ) , .D( n1036 ) , .QN( n117 ) );
  DFF_X1 text_in_r_reg_59 (.CK( clk ) , .D( n1037 ) , .QN( n119 ) );
  DFF_X1 text_in_r_reg_6 (.CK( clk ) , .QN( n13 ) , .D( n984 ) );
  DFF_X1 text_in_r_reg_60 (.CK( clk ) , .D( n1038 ) , .QN( n121 ) );
  DFF_X1 text_in_r_reg_61 (.CK( clk ) , .D( n1039 ) , .QN( n123 ) );
  DFF_X1 text_in_r_reg_62 (.CK( clk ) , .D( n1040 ) , .QN( n125 ) );
  DFF_X1 text_in_r_reg_63 (.CK( clk ) , .D( n1041 ) , .QN( n127 ) );
  DFF_X1 text_in_r_reg_64 (.CK( clk ) , .D( n1042 ) , .QN( n129 ) );
  DFF_X1 text_in_r_reg_65 (.CK( clk ) , .D( n1043 ) , .QN( n131 ) );
  DFF_X1 text_in_r_reg_66 (.CK( clk ) , .D( n1044 ) , .QN( n133 ) );
  DFF_X1 text_in_r_reg_67 (.CK( clk ) , .D( n1045 ) , .QN( n135 ) );
  DFF_X1 text_in_r_reg_68 (.CK( clk ) , .D( n1046 ) , .QN( n137 ) );
  DFF_X1 text_in_r_reg_69 (.CK( clk ) , .D( n1047 ) , .QN( n139 ) );
  DFF_X1 text_in_r_reg_7 (.CK( clk ) , .QN( n15 ) , .D( n985 ) );
  DFF_X1 text_in_r_reg_70 (.CK( clk ) , .D( n1048 ) , .QN( n141 ) );
  DFF_X1 text_in_r_reg_71 (.CK( clk ) , .D( n1049 ) , .QN( n143 ) );
  DFF_X1 text_in_r_reg_72 (.CK( clk ) , .D( n1050 ) , .QN( n145 ) );
  DFF_X1 text_in_r_reg_73 (.CK( clk ) , .D( n1051 ) , .QN( n147 ) );
  DFF_X1 text_in_r_reg_74 (.CK( clk ) , .D( n1052 ) , .QN( n149 ) );
  DFF_X1 text_in_r_reg_75 (.CK( clk ) , .D( n1053 ) , .QN( n151 ) );
  DFF_X1 text_in_r_reg_76 (.CK( clk ) , .D( n1054 ) , .QN( n153 ) );
  DFF_X1 text_in_r_reg_77 (.CK( clk ) , .D( n1055 ) , .QN( n155 ) );
  DFF_X1 text_in_r_reg_78 (.CK( clk ) , .D( n1056 ) , .QN( n157 ) );
  DFF_X1 text_in_r_reg_79 (.CK( clk ) , .D( n1057 ) , .QN( n159 ) );
  DFF_X1 text_in_r_reg_8 (.CK( clk ) , .QN( n17 ) , .D( n986 ) );
  DFF_X1 text_in_r_reg_80 (.CK( clk ) , .D( n1058 ) , .QN( n161 ) );
  DFF_X1 text_in_r_reg_81 (.CK( clk ) , .D( n1059 ) , .QN( n163 ) );
  DFF_X1 text_in_r_reg_82 (.CK( clk ) , .D( n1060 ) , .QN( n165 ) );
  DFF_X1 text_in_r_reg_83 (.CK( clk ) , .D( n1061 ) , .QN( n167 ) );
  DFF_X1 text_in_r_reg_84 (.CK( clk ) , .D( n1062 ) , .QN( n169 ) );
  DFF_X1 text_in_r_reg_85 (.CK( clk ) , .D( n1063 ) , .QN( n171 ) );
  DFF_X1 text_in_r_reg_86 (.CK( clk ) , .D( n1064 ) , .QN( n173 ) );
  DFF_X1 text_in_r_reg_87 (.CK( clk ) , .D( n1065 ) , .QN( n175 ) );
  DFF_X1 text_in_r_reg_88 (.CK( clk ) , .D( n1066 ) , .QN( n177 ) );
  DFF_X1 text_in_r_reg_89 (.CK( clk ) , .D( n1067 ) , .QN( n179 ) );
  DFF_X1 text_in_r_reg_9 (.CK( clk ) , .QN( n19 ) , .D( n987 ) );
  DFF_X1 text_in_r_reg_90 (.CK( clk ) , .D( n1068 ) , .QN( n181 ) );
  DFF_X1 text_in_r_reg_91 (.CK( clk ) , .D( n1069 ) , .QN( n183 ) );
  DFF_X1 text_in_r_reg_92 (.CK( clk ) , .D( n1070 ) , .QN( n185 ) );
  DFF_X1 text_in_r_reg_93 (.CK( clk ) , .D( n1071 ) , .QN( n187 ) );
  DFF_X1 text_in_r_reg_94 (.CK( clk ) , .D( n1072 ) , .QN( n189 ) );
  DFF_X1 text_in_r_reg_95 (.CK( clk ) , .D( n1073 ) , .QN( n191 ) );
  DFF_X1 text_in_r_reg_96 (.CK( clk ) , .D( n1074 ) , .QN( n193 ) );
  DFF_X1 text_in_r_reg_97 (.CK( clk ) , .D( n1075 ) , .QN( n195 ) );
  DFF_X1 text_in_r_reg_98 (.CK( clk ) , .D( n1076 ) , .QN( n197 ) );
  DFF_X1 text_in_r_reg_99 (.CK( clk ) , .D( n1077 ) , .QN( n199 ) );
  DFF_X1 text_out_reg_0 (.D( N505 ) , .CK( clk ) , .Q( text_out[0] ) );
  DFF_X1 text_out_reg_1 (.D( N504 ) , .CK( clk ) , .Q( text_out[1] ) );
  DFF_X1 text_out_reg_10 (.D( N471 ) , .CK( clk ) , .Q( text_out[10] ) );
  DFF_X1 text_out_reg_100 (.D( N477 ) , .CK( clk ) , .Q( text_out[100] ) );
  DFF_X1 text_out_reg_101 (.D( N476 ) , .CK( clk ) , .Q( text_out[101] ) );
  DFF_X1 text_out_reg_102 (.D( N475 ) , .CK( clk ) , .Q( text_out[102] ) );
  DFF_X1 text_out_reg_103 (.D( N474 ) , .CK( clk ) , .Q( text_out[103] ) );
  DFF_X1 text_out_reg_104 (.D( N449 ) , .CK( clk ) , .Q( text_out[104] ) );
  DFF_X1 text_out_reg_105 (.D( N448 ) , .CK( clk ) , .Q( text_out[105] ) );
  DFF_X1 text_out_reg_106 (.D( N447 ) , .CK( clk ) , .Q( text_out[106] ) );
  DFF_X1 text_out_reg_107 (.D( N446 ) , .CK( clk ) , .Q( text_out[107] ) );
  DFF_X1 text_out_reg_108 (.D( N445 ) , .CK( clk ) , .Q( text_out[108] ) );
  DFF_X1 text_out_reg_109 (.D( N444 ) , .CK( clk ) , .Q( text_out[109] ) );
  DFF_X1 text_out_reg_11 (.D( N470 ) , .CK( clk ) , .Q( text_out[11] ) );
  DFF_X1 text_out_reg_110 (.D( N443 ) , .CK( clk ) , .Q( text_out[110] ) );
  DFF_X1 text_out_reg_111 (.D( N442 ) , .CK( clk ) , .Q( text_out[111] ) );
  DFF_X1 text_out_reg_112 (.D( N417 ) , .CK( clk ) , .Q( text_out[112] ) );
  DFF_X1 text_out_reg_113 (.D( N416 ) , .CK( clk ) , .Q( text_out[113] ) );
  DFF_X1 text_out_reg_114 (.D( N415 ) , .CK( clk ) , .Q( text_out[114] ) );
  DFF_X1 text_out_reg_115 (.D( N414 ) , .CK( clk ) , .Q( text_out[115] ) );
  DFF_X1 text_out_reg_116 (.D( N413 ) , .CK( clk ) , .Q( text_out[116] ) );
  DFF_X1 text_out_reg_117 (.D( N412 ) , .CK( clk ) , .Q( text_out[117] ) );
  DFF_X1 text_out_reg_118 (.D( N411 ) , .CK( clk ) , .Q( text_out[118] ) );
  DFF_X1 text_out_reg_119 (.D( N410 ) , .CK( clk ) , .Q( text_out[119] ) );
  DFF_X1 text_out_reg_12 (.D( N469 ) , .CK( clk ) , .Q( text_out[12] ) );
  DFF_X1 text_out_reg_120 (.D( N385 ) , .CK( clk ) , .Q( text_out[120] ) );
  DFF_X1 text_out_reg_121 (.D( N384 ) , .CK( clk ) , .Q( text_out[121] ) );
  DFF_X1 text_out_reg_122 (.D( N383 ) , .CK( clk ) , .Q( text_out[122] ) );
  DFF_X1 text_out_reg_123 (.D( N382 ) , .CK( clk ) , .Q( text_out[123] ) );
  DFF_X1 text_out_reg_124 (.D( N381 ) , .CK( clk ) , .Q( text_out[124] ) );
  DFF_X1 text_out_reg_125 (.D( N380 ) , .CK( clk ) , .Q( text_out[125] ) );
  DFF_X1 text_out_reg_126 (.D( N379 ) , .CK( clk ) , .Q( text_out[126] ) );
  DFF_X1 text_out_reg_127 (.D( N378 ) , .CK( clk ) , .Q( text_out[127] ) );
  DFF_X1 text_out_reg_13 (.D( N468 ) , .CK( clk ) , .Q( text_out[13] ) );
  DFF_X1 text_out_reg_14 (.D( N467 ) , .CK( clk ) , .Q( text_out[14] ) );
  DFF_X1 text_out_reg_15 (.D( N466 ) , .CK( clk ) , .Q( text_out[15] ) );
  DFF_X1 text_out_reg_16 (.D( N441 ) , .CK( clk ) , .Q( text_out[16] ) );
  DFF_X1 text_out_reg_17 (.D( N440 ) , .CK( clk ) , .Q( text_out[17] ) );
  DFF_X1 text_out_reg_18 (.D( N439 ) , .CK( clk ) , .Q( text_out[18] ) );
  DFF_X1 text_out_reg_19 (.D( N438 ) , .CK( clk ) , .Q( text_out[19] ) );
  DFF_X1 text_out_reg_2 (.D( N503 ) , .CK( clk ) , .Q( text_out[2] ) );
  DFF_X1 text_out_reg_20 (.D( N437 ) , .CK( clk ) , .Q( text_out[20] ) );
  DFF_X1 text_out_reg_21 (.D( N436 ) , .CK( clk ) , .Q( text_out[21] ) );
  DFF_X1 text_out_reg_22 (.D( N435 ) , .CK( clk ) , .Q( text_out[22] ) );
  DFF_X1 text_out_reg_23 (.D( N434 ) , .CK( clk ) , .Q( text_out[23] ) );
  DFF_X1 text_out_reg_24 (.D( N409 ) , .CK( clk ) , .Q( text_out[24] ) );
  DFF_X1 text_out_reg_25 (.D( N408 ) , .CK( clk ) , .Q( text_out[25] ) );
  DFF_X1 text_out_reg_26 (.D( N407 ) , .CK( clk ) , .Q( text_out[26] ) );
  DFF_X1 text_out_reg_27 (.D( N406 ) , .CK( clk ) , .Q( text_out[27] ) );
  DFF_X1 text_out_reg_28 (.D( N405 ) , .CK( clk ) , .Q( text_out[28] ) );
  DFF_X1 text_out_reg_29 (.D( N404 ) , .CK( clk ) , .Q( text_out[29] ) );
  DFF_X1 text_out_reg_3 (.D( N502 ) , .CK( clk ) , .Q( text_out[3] ) );
  DFF_X1 text_out_reg_30 (.D( N403 ) , .CK( clk ) , .Q( text_out[30] ) );
  DFF_X1 text_out_reg_31 (.D( N402 ) , .CK( clk ) , .Q( text_out[31] ) );
  DFF_X1 text_out_reg_32 (.D( N497 ) , .CK( clk ) , .Q( text_out[32] ) );
  DFF_X1 text_out_reg_33 (.D( N496 ) , .CK( clk ) , .Q( text_out[33] ) );
  DFF_X1 text_out_reg_34 (.D( N495 ) , .CK( clk ) , .Q( text_out[34] ) );
  DFF_X1 text_out_reg_35 (.D( N494 ) , .CK( clk ) , .Q( text_out[35] ) );
  DFF_X1 text_out_reg_36 (.D( N493 ) , .CK( clk ) , .Q( text_out[36] ) );
  DFF_X1 text_out_reg_37 (.D( N492 ) , .CK( clk ) , .Q( text_out[37] ) );
  DFF_X1 text_out_reg_38 (.D( N491 ) , .CK( clk ) , .Q( text_out[38] ) );
  DFF_X1 text_out_reg_39 (.D( N490 ) , .CK( clk ) , .Q( text_out[39] ) );
  DFF_X1 text_out_reg_4 (.D( N501 ) , .CK( clk ) , .Q( text_out[4] ) );
  DFF_X1 text_out_reg_40 (.D( N465 ) , .CK( clk ) , .Q( text_out[40] ) );
  DFF_X1 text_out_reg_41 (.D( N464 ) , .CK( clk ) , .Q( text_out[41] ) );
  DFF_X1 text_out_reg_42 (.D( N463 ) , .CK( clk ) , .Q( text_out[42] ) );
  DFF_X1 text_out_reg_43 (.D( N462 ) , .CK( clk ) , .Q( text_out[43] ) );
  DFF_X1 text_out_reg_44 (.D( N461 ) , .CK( clk ) , .Q( text_out[44] ) );
  DFF_X1 text_out_reg_45 (.D( N460 ) , .CK( clk ) , .Q( text_out[45] ) );
  DFF_X1 text_out_reg_46 (.D( N459 ) , .CK( clk ) , .Q( text_out[46] ) );
  DFF_X1 text_out_reg_47 (.D( N458 ) , .CK( clk ) , .Q( text_out[47] ) );
  DFF_X1 text_out_reg_48 (.D( N433 ) , .CK( clk ) , .Q( text_out[48] ) );
  DFF_X1 text_out_reg_49 (.D( N432 ) , .CK( clk ) , .Q( text_out[49] ) );
  DFF_X1 text_out_reg_5 (.D( N500 ) , .CK( clk ) , .Q( text_out[5] ) );
  DFF_X1 text_out_reg_50 (.D( N431 ) , .CK( clk ) , .Q( text_out[50] ) );
  DFF_X1 text_out_reg_51 (.D( N430 ) , .CK( clk ) , .Q( text_out[51] ) );
  DFF_X1 text_out_reg_52 (.D( N429 ) , .CK( clk ) , .Q( text_out[52] ) );
  DFF_X1 text_out_reg_53 (.D( N428 ) , .CK( clk ) , .Q( text_out[53] ) );
  DFF_X1 text_out_reg_54 (.D( N427 ) , .CK( clk ) , .Q( text_out[54] ) );
  DFF_X1 text_out_reg_55 (.D( N426 ) , .CK( clk ) , .Q( text_out[55] ) );
  DFF_X1 text_out_reg_56 (.D( N401 ) , .CK( clk ) , .Q( text_out[56] ) );
  DFF_X1 text_out_reg_57 (.D( N400 ) , .CK( clk ) , .Q( text_out[57] ) );
  DFF_X1 text_out_reg_58 (.D( N399 ) , .CK( clk ) , .Q( text_out[58] ) );
  DFF_X1 text_out_reg_59 (.D( N398 ) , .CK( clk ) , .Q( text_out[59] ) );
  DFF_X1 text_out_reg_6 (.D( N499 ) , .CK( clk ) , .Q( text_out[6] ) );
  DFF_X1 text_out_reg_60 (.D( N397 ) , .CK( clk ) , .Q( text_out[60] ) );
  DFF_X1 text_out_reg_61 (.D( N396 ) , .CK( clk ) , .Q( text_out[61] ) );
  DFF_X1 text_out_reg_62 (.D( N395 ) , .CK( clk ) , .Q( text_out[62] ) );
  DFF_X1 text_out_reg_63 (.D( N394 ) , .CK( clk ) , .Q( text_out[63] ) );
  DFF_X1 text_out_reg_64 (.D( N489 ) , .CK( clk ) , .Q( text_out[64] ) );
  DFF_X1 text_out_reg_65 (.D( N488 ) , .CK( clk ) , .Q( text_out[65] ) );
  DFF_X1 text_out_reg_66 (.D( N487 ) , .CK( clk ) , .Q( text_out[66] ) );
  DFF_X1 text_out_reg_67 (.D( N486 ) , .CK( clk ) , .Q( text_out[67] ) );
  DFF_X1 text_out_reg_68 (.D( N485 ) , .CK( clk ) , .Q( text_out[68] ) );
  DFF_X1 text_out_reg_69 (.D( N484 ) , .CK( clk ) , .Q( text_out[69] ) );
  DFF_X1 text_out_reg_7 (.D( N498 ) , .CK( clk ) , .Q( text_out[7] ) );
  DFF_X1 text_out_reg_70 (.D( N483 ) , .CK( clk ) , .Q( text_out[70] ) );
  DFF_X1 text_out_reg_71 (.D( N482 ) , .CK( clk ) , .Q( text_out[71] ) );
  DFF_X1 text_out_reg_72 (.D( N457 ) , .CK( clk ) , .Q( text_out[72] ) );
  DFF_X1 text_out_reg_73 (.D( N456 ) , .CK( clk ) , .Q( text_out[73] ) );
  DFF_X1 text_out_reg_74 (.D( N455 ) , .CK( clk ) , .Q( text_out[74] ) );
  DFF_X1 text_out_reg_75 (.D( N454 ) , .CK( clk ) , .Q( text_out[75] ) );
  DFF_X1 text_out_reg_76 (.D( N453 ) , .CK( clk ) , .Q( text_out[76] ) );
  DFF_X1 text_out_reg_77 (.D( N452 ) , .CK( clk ) , .Q( text_out[77] ) );
  DFF_X1 text_out_reg_78 (.D( N451 ) , .CK( clk ) , .Q( text_out[78] ) );
  DFF_X1 text_out_reg_79 (.D( N450 ) , .CK( clk ) , .Q( text_out[79] ) );
  DFF_X1 text_out_reg_8 (.D( N473 ) , .CK( clk ) , .Q( text_out[8] ) );
  DFF_X1 text_out_reg_80 (.D( N425 ) , .CK( clk ) , .Q( text_out[80] ) );
  DFF_X1 text_out_reg_81 (.D( N424 ) , .CK( clk ) , .Q( text_out[81] ) );
  DFF_X1 text_out_reg_82 (.D( N423 ) , .CK( clk ) , .Q( text_out[82] ) );
  DFF_X1 text_out_reg_83 (.D( N422 ) , .CK( clk ) , .Q( text_out[83] ) );
  DFF_X1 text_out_reg_84 (.D( N421 ) , .CK( clk ) , .Q( text_out[84] ) );
  DFF_X1 text_out_reg_85 (.D( N420 ) , .CK( clk ) , .Q( text_out[85] ) );
  DFF_X1 text_out_reg_86 (.D( N419 ) , .CK( clk ) , .Q( text_out[86] ) );
  DFF_X1 text_out_reg_87 (.D( N418 ) , .CK( clk ) , .Q( text_out[87] ) );
  DFF_X1 text_out_reg_88 (.D( N393 ) , .CK( clk ) , .Q( text_out[88] ) );
  DFF_X1 text_out_reg_89 (.D( N392 ) , .CK( clk ) , .Q( text_out[89] ) );
  DFF_X1 text_out_reg_9 (.D( N472 ) , .CK( clk ) , .Q( text_out[9] ) );
  DFF_X1 text_out_reg_90 (.D( N391 ) , .CK( clk ) , .Q( text_out[90] ) );
  DFF_X1 text_out_reg_91 (.D( N390 ) , .CK( clk ) , .Q( text_out[91] ) );
  DFF_X1 text_out_reg_92 (.D( N389 ) , .CK( clk ) , .Q( text_out[92] ) );
  DFF_X1 text_out_reg_93 (.D( N388 ) , .CK( clk ) , .Q( text_out[93] ) );
  DFF_X1 text_out_reg_94 (.D( N387 ) , .CK( clk ) , .Q( text_out[94] ) );
  DFF_X1 text_out_reg_95 (.D( N386 ) , .CK( clk ) , .Q( text_out[95] ) );
  DFF_X1 text_out_reg_96 (.D( N481 ) , .CK( clk ) , .Q( text_out[96] ) );
  DFF_X1 text_out_reg_97 (.D( N480 ) , .CK( clk ) , .Q( text_out[97] ) );
  DFF_X1 text_out_reg_98 (.D( N479 ) , .CK( clk ) , .Q( text_out[98] ) );
  DFF_X1 text_out_reg_99 (.D( N478 ) , .CK( clk ) , .Q( text_out[99] ) );
  XNOR2_X1 u0_U10 (.ZN( u0_n57 ) , .B( u0_subword_3 ) , .A( w0_3 ) );
  NAND2_X1 u0_U100 (.A1( key[62] ) , .A2( ld ) , .ZN( u0_n163 ) );
  NAND2_X1 u0_U101 (.A1( key[15] ) , .A2( ld ) , .ZN( u0_n114 ) );
  NAND2_X1 u0_U102 (.A1( key[74] ) , .A2( ld ) , .ZN( u0_n267 ) );
  NAND2_X1 u0_U103 (.A1( key[10] ) , .A2( ld ) , .ZN( u0_n129 ) );
  NAND2_X1 u0_U104 (.A1( key[72] ) , .A2( ld ) , .ZN( u0_n271 ) );
  NAND2_X1 u0_U105 (.A2( key[127] ) , .A1( ld ) , .ZN( u0_n2 ) );
  NAND2_X1 u0_U106 (.A1( key[6] ) , .A2( ld ) , .ZN( u0_n141 ) );
  NAND2_X1 u0_U107 (.A1( key[2] ) , .A2( ld ) , .ZN( u0_n153 ) );
  NAND2_X1 u0_U108 (.A1( key[73] ) , .A2( ld ) , .ZN( u0_n269 ) );
  NAND2_X1 u0_U109 (.A1( key[30] ) , .A2( ld ) , .ZN( u0_n69 ) );
  XNOR2_X1 u0_U11 (.ZN( u0_n41 ) , .B( u0_subword_11 ) , .A( w0_11 ) );
  NAND2_X1 u0_U110 (.A1( key[29] ) , .A2( ld ) , .ZN( u0_n72 ) );
  NAND2_X1 u0_U111 (.A1( key[17] ) , .A2( ld ) , .ZN( u0_n108 ) );
  NAND2_X1 u0_U112 (.A1( key[18] ) , .A2( ld ) , .ZN( u0_n105 ) );
  NAND2_X1 u0_U113 (.A1( key[16] ) , .A2( ld ) , .ZN( u0_n111 ) );
  NAND2_X1 u0_U114 (.A1( key[9] ) , .A2( ld ) , .ZN( u0_n132 ) );
  NAND2_X1 u0_U115 (.A1( key[19] ) , .A2( ld ) , .ZN( u0_n102 ) );
  NAND2_X1 u0_U116 (.A1( key[8] ) , .A2( ld ) , .ZN( u0_n135 ) );
  NAND2_X1 u0_U117 (.A1( key[3] ) , .A2( ld ) , .ZN( u0_n150 ) );
  NAND2_X1 u0_U118 (.A1( key[0] ) , .A2( ld ) , .ZN( u0_n159 ) );
  NAND2_X1 u0_U119 (.A1( key[5] ) , .A2( ld ) , .ZN( u0_n144 ) );
  XNOR2_X1 u0_U12 (.ZN( u0_n33 ) , .B( u0_subword_15 ) , .A( w0_15 ) );
  NAND2_X1 u0_U120 (.A1( key[1] ) , .A2( ld ) , .ZN( u0_n156 ) );
  OAI21_X1 u0_U121 (.B1( ld ) , .ZN( u0_N181 ) , .B2( u0_n139 ) , .A( u0_n209 ) );
  NAND2_X1 u0_U122 (.A1( key[39] ) , .A2( ld ) , .ZN( u0_n209 ) );
  OAI21_X1 u0_U123 (.B1( ld ) , .ZN( u0_N135 ) , .B2( u0_n170 ) , .A( u0_n233 ) );
  NAND2_X1 u0_U124 (.A1( key[91] ) , .A2( ld ) , .ZN( u0_n233 ) );
  OAI21_X1 u0_U125 (.B1( ld ) , .ZN( u0_N57 ) , .B2( u0_n33 ) , .A( u0_n34 ) );
  NAND2_X1 u0_U126 (.A1( key[111] ) , .A2( ld ) , .ZN( u0_n34 ) );
  OAI21_X1 u0_U127 (.B1( ld ) , .ZN( u0_N46 ) , .B2( u0_n55 ) , .A( u0_n56 ) );
  NAND2_X1 u0_U128 (.A1( key[100] ) , .A2( ld ) , .ZN( u0_n56 ) );
  OAI21_X1 u0_U129 (.B1( ld ) , .ZN( u0_N45 ) , .B2( u0_n57 ) , .A( u0_n58 ) );
  XNOR2_X1 u0_U13 (.ZN( u0_n17 ) , .B( u0_subword_23 ) , .A( w0_23 ) );
  NAND2_X1 u0_U130 (.A1( key[99] ) , .A2( ld ) , .ZN( u0_n58 ) );
  OAI21_X1 u0_U131 (.B1( ld ) , .ZN( u0_N43 ) , .B2( u0_n61 ) , .A( u0_n62 ) );
  NAND2_X1 u0_U132 (.A1( key[97] ) , .A2( ld ) , .ZN( u0_n62 ) );
  OAI21_X1 u0_U133 (.B1( ld ) , .ZN( u0_N54 ) , .B2( u0_n39 ) , .A( u0_n40 ) );
  NAND2_X1 u0_U134 (.A1( key[108] ) , .A2( ld ) , .ZN( u0_n40 ) );
  OAI21_X1 u0_U135 (.B1( ld ) , .ZN( u0_N51 ) , .B2( u0_n45 ) , .A( u0_n46 ) );
  NAND2_X1 u0_U136 (.A1( key[105] ) , .A2( ld ) , .ZN( u0_n46 ) );
  OAI21_X1 u0_U137 (.B1( ld ) , .ZN( u0_N65 ) , .B2( u0_n17 ) , .A( u0_n18 ) );
  NAND2_X1 u0_U138 (.A1( key[119] ) , .A2( ld ) , .ZN( u0_n18 ) );
  OAI21_X1 u0_U139 (.B1( ld ) , .ZN( u0_N71 ) , .B2( u0_n5 ) , .A( u0_n6 ) );
  XNOR2_X1 u0_U14 (.ZN( u0_n45 ) , .B( u0_subword_9 ) , .A( w0_9 ) );
  NAND2_X1 u0_U140 (.A1( key[125] ) , .A2( ld ) , .ZN( u0_n6 ) );
  OAI21_X1 u0_U141 (.B1( ld ) , .ZN( u0_N70 ) , .B2( u0_n7 ) , .A( u0_n8 ) );
  NAND2_X1 u0_U142 (.A1( key[124] ) , .A2( ld ) , .ZN( u0_n8 ) );
  OAI21_X1 u0_U143 (.B1( ld ) , .ZN( u0_N69 ) , .A( u0_n10 ) , .B2( u0_n9 ) );
  NAND2_X1 u0_U144 (.A1( key[123] ) , .A2( ld ) , .ZN( u0_n10 ) );
  OAI21_X1 u0_U145 (.B1( ld ) , .ZN( u0_N123 ) , .B2( u0_n194 ) , .A( u0_n257 ) );
  NAND2_X1 u0_U146 (.A1( key[79] ) , .A2( ld ) , .ZN( u0_n257 ) );
  OAI21_X1 u0_U147 (.B1( ld ) , .ZN( u0_N131 ) , .B2( u0_n178 ) , .A( u0_n241 ) );
  NAND2_X1 u0_U148 (.A1( key[87] ) , .A2( ld ) , .ZN( u0_n241 ) );
  OAI21_X1 u0_U149 (.B1( ld ) , .ZN( u0_N121 ) , .B2( u0_n198 ) , .A( u0_n261 ) );
  XNOR2_X1 u0_U15 (.ZN( u0_n23 ) , .B( u0_subword_20 ) , .A( w0_20 ) );
  NAND2_X1 u0_U150 (.A1( key[77] ) , .A2( ld ) , .ZN( u0_n261 ) );
  OAI21_X1 u0_U151 (.B1( ld ) , .ZN( u0_N47 ) , .B2( u0_n53 ) , .A( u0_n54 ) );
  NAND2_X1 u0_U152 (.A1( key[101] ) , .A2( ld ) , .ZN( u0_n54 ) );
  OAI21_X1 u0_U153 (.B1( ld ) , .ZN( u0_N63 ) , .B2( u0_n21 ) , .A( u0_n22 ) );
  NAND2_X1 u0_U154 (.A1( key[117] ) , .A2( ld ) , .ZN( u0_n22 ) );
  OAI21_X1 u0_U155 (.B1( ld ) , .ZN( u0_N129 ) , .B2( u0_n182 ) , .A( u0_n245 ) );
  NAND2_X1 u0_U156 (.A1( key[85] ) , .A2( ld ) , .ZN( u0_n245 ) );
  OAI21_X1 u0_U157 (.B1( ld ) , .ZN( u0_N62 ) , .B2( u0_n23 ) , .A( u0_n24 ) );
  NAND2_X1 u0_U158 (.A1( key[116] ) , .A2( ld ) , .ZN( u0_n24 ) );
  OAI21_X1 u0_U159 (.B1( ld ) , .ZN( u0_N55 ) , .B2( u0_n37 ) , .A( u0_n38 ) );
  XNOR2_X1 u0_U16 (.ZN( u0_n37 ) , .B( u0_subword_13 ) , .A( w0_13 ) );
  NAND2_X1 u0_U160 (.A1( key[109] ) , .A2( ld ) , .ZN( u0_n38 ) );
  OAI21_X1 u0_U161 (.B1( ld ) , .ZN( u0_N120 ) , .B2( u0_n200 ) , .A( u0_n263 ) );
  NAND2_X1 u0_U162 (.A1( key[76] ) , .A2( ld ) , .ZN( u0_n263 ) );
  OAI21_X1 u0_U163 (.B1( ld ) , .ZN( u0_N53 ) , .B2( u0_n41 ) , .A( u0_n42 ) );
  NAND2_X1 u0_U164 (.A1( key[107] ) , .A2( ld ) , .ZN( u0_n42 ) );
  OAI21_X1 u0_U165 (.B1( ld ) , .ZN( u0_N268 ) , .B2( u0_n74 ) , .A( u0_n75 ) );
  NAND2_X1 u0_U166 (.A1( key[28] ) , .A2( ld ) , .ZN( u0_n75 ) );
  OAI21_X1 u0_U167 (.B1( ld ) , .ZN( u0_N271 ) , .B2( u0_n65 ) , .A( u0_n66 ) );
  NAND2_X1 u0_U168 (.A1( key[31] ) , .A2( ld ) , .ZN( u0_n66 ) );
  OAI21_X1 u0_U169 (.B1( ld ) , .ZN( u0_N260 ) , .B2( u0_n98 ) , .A( u0_n99 ) );
  XNOR2_X1 u0_U17 (.ZN( u0_n53 ) , .B( u0_subword_5 ) , .A( w0_5 ) );
  NAND2_X1 u0_U170 (.A1( key[20] ) , .A2( ld ) , .ZN( u0_n99 ) );
  OAI21_X1 u0_U171 (.B1( ld ) , .ZN( u0_N251 ) , .B2( u0_n125 ) , .A( u0_n126 ) );
  NAND2_X1 u0_U172 (.A1( key[11] ) , .A2( ld ) , .ZN( u0_n126 ) );
  OAI21_X1 u0_U173 (.B1( ld ) , .ZN( u0_N244 ) , .B2( u0_n146 ) , .A( u0_n147 ) );
  NAND2_X1 u0_U174 (.A1( key[4] ) , .A2( ld ) , .ZN( u0_n147 ) );
  OAI21_X1 u0_U175 (.B1( ld ) , .ZN( u0_N115 ) , .B2( u0_n210 ) , .A( u0_n273 ) );
  NAND2_X1 u0_U176 (.A1( key[71] ) , .A2( ld ) , .ZN( u0_n273 ) );
  OAI21_X1 u0_U177 (.B1( ld ) , .ZN( u0_N113 ) , .B2( u0_n214 ) , .A( u0_n277 ) );
  NAND2_X1 u0_U178 (.A1( key[69] ) , .A2( ld ) , .ZN( u0_n277 ) );
  OAI21_X1 u0_U179 (.B1( ld ) , .ZN( u0_N111 ) , .B2( u0_n218 ) , .A( u0_n281 ) );
  XNOR2_X1 u0_U18 (.ZN( u0_n21 ) , .B( u0_subword_21 ) , .A( w0_21 ) );
  NAND2_X1 u0_U180 (.A1( key[67] ) , .A2( ld ) , .ZN( u0_n281 ) );
  XNOR2_X1 u0_U181 (.ZN( u0_n226 ) , .B( u0_subword_31 ) , .A( w0_31 ) );
  OAI21_X1 u0_U182 (.B1( ld ) , .ZN( u0_N42 ) , .B2( u0_n63 ) , .A( u0_n64 ) );
  XNOR2_X1 u0_U183 (.ZN( u0_n61 ) , .B( u0_subword_1 ) , .A( w0_1 ) );
  OAI21_X1 u0_U184 (.B1( ld ) , .ZN( u0_N50 ) , .B2( u0_n47 ) , .A( u0_n48 ) );
  XNOR2_X1 u0_U185 (.ZN( u0_n55 ) , .B( u0_subword_4 ) , .A( w0_4 ) );
  OAI21_X1 u0_U186 (.B1( ld ) , .ZN( u0_N44 ) , .B2( u0_n59 ) , .A( u0_n60 ) );
  OAI21_X1 u0_U187 (.B1( ld ) , .ZN( u0_N59 ) , .B2( u0_n29 ) , .A( u0_n30 ) );
  OAI21_X1 u0_U188 (.B1( ld ) , .ZN( u0_N247 ) , .B2( u0_n137 ) , .A( u0_n138 ) );
  OAI21_X1 u0_U189 (.B1( ld ) , .ZN( u0_N67 ) , .B2( u0_n13 ) , .A( u0_n14 ) );
  NAND2_X1 u0_U19 (.A1( key[22] ) , .A2( ld ) , .ZN( u0_n93 ) );
  OAI21_X1 u0_U190 (.B1( ld ) , .ZN( u0_N252 ) , .B2( u0_n122 ) , .A( u0_n123 ) );
  OAI21_X1 u0_U191 (.B1( ld ) , .ZN( u0_N186 ) , .B2( u0_n124 ) , .A( u0_n199 ) );
  OAI21_X1 u0_U192 (.B1( ld ) , .ZN( u0_N269 ) , .B2( u0_n71 ) , .A( u0_n72 ) );
  OAI21_X1 u0_U193 (.B1( ld ) , .ZN( u0_N73 ) , .B2( u0_n1 ) , .A( u0_n2 ) );
  XNOR2_X1 u0_U194 (.ZN( u0_n15 ) , .A( u0_n240 ) , .B( u0_n246 ) );
  XNOR2_X1 u0_U195 (.B( u0_n248 ) , .ZN( u0_n86 ) , .A( u0_n88 ) );
  OAI21_X1 u0_U196 (.B1( ld ) , .ZN( u0_N254 ) , .B2( u0_n116 ) , .A( u0_n117 ) );
  OAI21_X1 u0_U197 (.B1( ld ) , .ZN( u0_N109 ) , .B2( u0_n222 ) , .A( u0_n285 ) );
  OAI21_X1 u0_U198 (.B1( ld ) , .ZN( u0_N119 ) , .B2( u0_n202 ) , .A( u0_n265 ) );
  OAI21_X1 u0_U199 (.B1( ld ) , .ZN( u0_N185 ) , .B2( u0_n127 ) , .A( u0_n201 ) );
  XNOR2_X1 u0_U20 (.ZN( u0_n25 ) , .B( u0_subword_19 ) , .A( w0_19 ) );
  OAI21_X1 u0_U200 (.B1( ld ) , .ZN( u0_N136 ) , .B2( u0_n168 ) , .A( u0_n231 ) );
  OAI21_X1 u0_U201 (.B1( ld ) , .ZN( u0_N202 ) , .A( u0_n167 ) , .B2( u0_n76 ) );
  XNOR2_X1 u0_U202 (.ZN( u0_n31 ) , .B( u0_subword_16 ) , .A( w0_16 ) );
  INV_X1 u0_U203 (.A( u0_n250 ) , .ZN( w3_13 ) );
  OAI21_X1 u0_U204 (.B1( ld ) , .ZN( u0_N128 ) , .B2( u0_n184 ) , .A( u0_n247 ) );
  OAI21_X1 u0_U205 (.B1( ld ) , .ZN( u0_N194 ) , .B2( u0_n100 ) , .A( u0_n183 ) );
  INV_X1 u0_U206 (.A( u0_n254 ) , .ZN( w3_14 ) );
  OAI21_X1 u0_U207 (.B1( ld ) , .ZN( u0_N245 ) , .B2( u0_n143 ) , .A( u0_n144 ) );
  OAI21_X1 u0_U208 (.B1( ld ) , .ZN( u0_N179 ) , .B2( u0_n145 ) , .A( u0_n213 ) );
  OAI21_X1 u0_U209 (.B1( ld ) , .ZN( u0_N249 ) , .B2( u0_n131 ) , .A( u0_n132 ) );
  XNOR2_X1 u0_U21 (.ZN( u0_n49 ) , .B( u0_subword_7 ) , .A( w0_7 ) );
  INV_X1 u0_U210 (.A( u0_n258 ) , .ZN( w3_12 ) );
  XNOR2_X1 u0_U211 (.ZN( u0_n43 ) , .B( u0_subword_10 ) , .A( w0_10 ) );
  XNOR2_X1 u0_U212 (.ZN( u0_n59 ) , .A( u0_subword_2 ) , .B( w0_2 ) );
  OAI21_X1 u0_U213 (.B1( ld ) , .ZN( u0_N49 ) , .B2( u0_n49 ) , .A( u0_n50 ) );
  OAI21_X1 u0_U214 (.B1( ld ) , .ZN( u0_N125 ) , .B2( u0_n190 ) , .A( u0_n253 ) );
  XNOR2_X1 u0_U215 (.ZN( u0_n164 ) , .B( u0_n262 ) , .A( u0_n3 ) );
  OAI21_X1 u0_U216 (.B1( ld ) , .ZN( u0_N262 ) , .B2( u0_n92 ) , .A( u0_n93 ) );
  XNOR2_X1 u0_U217 (.ZN( u0_n27 ) , .B( u0_subword_18 ) , .A( w0_18 ) );
  OAI21_X1 u0_U218 (.B1( ld ) , .ZN( u0_N139 ) , .B2( u0_n162 ) , .A( u0_n225 ) );
  OAI21_X1 u0_U219 (.B1( ld ) , .ZN( u0_N205 ) , .A( u0_n161 ) , .B2( u0_n67 ) );
  XNOR2_X1 u0_U22 (.ZN( u0_n29 ) , .B( u0_subword_17 ) , .A( w0_17 ) );
  OAI21_X1 u0_U220 (.B1( ld ) , .ZN( u0_N112 ) , .B2( u0_n216 ) , .A( u0_n279 ) );
  OAI21_X1 u0_U221 (.B1( ld ) , .ZN( u0_N178 ) , .B2( u0_n148 ) , .A( u0_n215 ) );
  OAI21_X1 u0_U222 (.B1( ld ) , .ZN( u0_N246 ) , .B2( u0_n140 ) , .A( u0_n141 ) );
  OAI21_X1 u0_U223 (.B1( ld ) , .ZN( u0_N243 ) , .B2( u0_n149 ) , .A( u0_n150 ) );
  OAI21_X1 u0_U224 (.B1( ld ) , .ZN( u0_N177 ) , .B2( u0_n151 ) , .A( u0_n217 ) );
  OAI21_X1 u0_U225 (.B1( ld ) , .ZN( u0_N133 ) , .B2( u0_n174 ) , .A( u0_n237 ) );
  OAI21_X1 u0_U226 (.B1( ld ) , .ZN( u0_N259 ) , .B2( u0_n101 ) , .A( u0_n102 ) );
  OAI21_X1 u0_U227 (.B1( ld ) , .ZN( u0_N61 ) , .B2( u0_n25 ) , .A( u0_n26 ) );
  OAI21_X1 u0_U228 (.B1( ld ) , .ZN( u0_N255 ) , .B2( u0_n113 ) , .A( u0_n114 ) );
  OAI21_X1 u0_U229 (.B1( ld ) , .ZN( u0_N189 ) , .B2( u0_n115 ) , .A( u0_n193 ) );
  XNOR2_X1 u0_U23 (.ZN( u0_n39 ) , .B( u0_subword_12 ) , .A( w0_12 ) );
  INV_X1 u0_U230 (.A( u0_n264 ) , .ZN( w3_15 ) );
  OAI21_X1 u0_U231 (.B1( ld ) , .ZN( u0_N263 ) , .B2( u0_n89 ) , .A( u0_n90 ) );
  OAI21_X1 u0_U232 (.B1( ld ) , .ZN( u0_N197 ) , .A( u0_n177 ) , .B2( u0_n91 ) );
  OAI21_X1 u0_U233 (.B1( ld ) , .ZN( u0_N117 ) , .B2( u0_n206 ) , .A( u0_n269 ) );
  OAI21_X1 u0_U234 (.B1( ld ) , .ZN( u0_N183 ) , .B2( u0_n133 ) , .A( u0_n205 ) );
  XNOR2_X1 u0_U235 (.ZN( u0_n47 ) , .B( u0_subword_8 ) , .A( w0_8 ) );
  OAI21_X1 u0_U236 (.B1( ld ) , .ZN( u0_N127 ) , .B2( u0_n186 ) , .A( u0_n249 ) );
  OAI21_X1 u0_U237 (.B1( ld ) , .ZN( u0_N193 ) , .B2( u0_n103 ) , .A( u0_n185 ) );
  OAI21_X1 u0_U238 (.B1( ld ) , .ZN( u0_N241 ) , .B2( u0_n155 ) , .A( u0_n156 ) );
  OAI21_X1 u0_U239 (.B1( ld ) , .ZN( u0_N175 ) , .B2( u0_n157 ) , .A( u0_n221 ) );
  NAND2_X1 u0_U24 (.A1( key[47] ) , .A2( ld ) , .ZN( u0_n193 ) );
  XNOR2_X1 u0_U240 (.ZN( u0_n35 ) , .B( u0_subword_14 ) , .A( w0_14 ) );
  OAI21_X1 u0_U241 (.B1( ld ) , .ZN( u0_N257 ) , .B2( u0_n107 ) , .A( u0_n108 ) );
  OAI21_X1 u0_U242 (.B1( ld ) , .ZN( u0_N191 ) , .B2( u0_n109 ) , .A( u0_n189 ) );
  OAI21_X1 u0_U243 (.B1( ld ) , .ZN( u0_N48 ) , .B2( u0_n51 ) , .A( u0_n52 ) );
  OAI21_X1 u0_U244 (.B1( ld ) , .ZN( u0_N116 ) , .B2( u0_n208 ) , .A( u0_n271 ) );
  OAI21_X1 u0_U245 (.B1( ld ) , .ZN( u0_N264 ) , .B2( u0_n86 ) , .A( u0_n87 ) );
  OAI21_X1 u0_U246 (.B1( ld ) , .ZN( u0_N66 ) , .B2( u0_n15 ) , .A( u0_n16 ) );
  OAI21_X1 u0_U247 (.B1( ld ) , .ZN( u0_N64 ) , .B2( u0_n19 ) , .A( u0_n20 ) );
  XNOR2_X1 u0_U248 (.ZN( u0_n63 ) , .B( u0_subword_0 ) , .A( w0_0 ) );
  OAI21_X1 u0_U249 (.B1( ld ) , .ZN( u0_N265 ) , .B2( u0_n83 ) , .A( u0_n84 ) );
  NAND2_X1 u0_U25 (.A1( key[55] ) , .A2( ld ) , .ZN( u0_n177 ) );
  OAI21_X1 u0_U250 (.B1( ld ) , .ZN( u0_N199 ) , .A( u0_n173 ) , .B2( u0_n85 ) );
  OAI21_X1 u0_U251 (.B1( ld ) , .ZN( u0_N108 ) , .B2( u0_n224 ) , .A( u0_n287 ) );
  OAI21_X1 u0_U252 (.B1( ld ) , .ZN( u0_N256 ) , .B2( u0_n110 ) , .A( u0_n111 ) );
  OAI21_X1 u0_U253 (.B1( ld ) , .ZN( u0_N58 ) , .B2( u0_n31 ) , .A( u0_n32 ) );
  XNOR2_X1 u0_U254 (.ZN( u0_n240 ) , .B( u0_subword_24 ) , .A( w0_24 ) );
  OAI21_X1 u0_U255 (.B1( ld ) , .ZN( u0_N267 ) , .B2( u0_n77 ) , .A( u0_n78 ) );
  OAI21_X1 u0_U256 (.B1( ld ) , .ZN( u0_N201 ) , .A( u0_n169 ) , .B2( u0_n79 ) );
  OAI21_X1 u0_U257 (.B1( ld ) , .ZN( u0_N72 ) , .B2( u0_n3 ) , .A( u0_n4 ) );
  OAI21_X1 u0_U258 (.B1( ld ) , .ZN( u0_N138 ) , .B2( u0_n164 ) , .A( u0_n227 ) );
  XNOR2_X1 u0_U259 (.ZN( u0_n51 ) , .B( u0_subword_6 ) , .A( w0_6 ) );
  NAND2_X1 u0_U26 (.A1( key[37] ) , .A2( ld ) , .ZN( u0_n213 ) );
  XNOR2_X1 u0_U260 (.ZN( u0_n230 ) , .B( u0_subword_29 ) , .A( w0_29 ) );
  OAI21_X1 u0_U261 (.B1( ld ) , .ZN( u0_N56 ) , .B2( u0_n35 ) , .A( u0_n36 ) );
  XNOR2_X1 u0_U262 (.ZN( u0_n19 ) , .B( u0_subword_22 ) , .A( w0_22 ) );
  OAI21_X1 u0_U263 (.B1( ld ) , .ZN( u0_N261 ) , .B2( u0_n95 ) , .A( u0_n96 ) );
  OAI21_X1 u0_U264 (.B1( ld ) , .ZN( u0_N195 ) , .A( u0_n181 ) , .B2( u0_n97 ) );
  OAI21_X1 u0_U265 (.B1( ld ) , .ZN( u0_N137 ) , .B2( u0_n166 ) , .A( u0_n229 ) );
  OAI21_X1 u0_U266 (.B1( ld ) , .ZN( u0_N203 ) , .A( u0_n165 ) , .B2( u0_n73 ) );
  OAI21_X1 u0_U267 (.B1( ld ) , .ZN( u0_N266 ) , .B2( u0_n80 ) , .A( u0_n81 ) );
  OAI21_X1 u0_U268 (.B1( ld ) , .ZN( u0_N114 ) , .B2( u0_n212 ) , .A( u0_n275 ) );
  OAI21_X1 u0_U269 (.B1( ld ) , .ZN( u0_N180 ) , .B2( u0_n142 ) , .A( u0_n211 ) );
  NAND2_X1 u0_U27 (.A1( key[35] ) , .A2( ld ) , .ZN( u0_n217 ) );
  OAI21_X1 u0_U270 (.B1( ld ) , .ZN( u0_N130 ) , .B2( u0_n180 ) , .A( u0_n243 ) );
  OAI21_X1 u0_U271 (.B1( ld ) , .ZN( u0_N196 ) , .A( u0_n179 ) , .B2( u0_n94 ) );
  OAI21_X1 u0_U272 (.B1( ld ) , .ZN( u0_N242 ) , .B2( u0_n152 ) , .A( u0_n153 ) );
  OAI21_X1 u0_U273 (.B1( ld ) , .ZN( u0_N122 ) , .B2( u0_n196 ) , .A( u0_n259 ) );
  OAI21_X1 u0_U274 (.B1( ld ) , .ZN( u0_N188 ) , .B2( u0_n118 ) , .A( u0_n195 ) );
  OAI21_X1 u0_U275 (.B1( ld ) , .ZN( u0_N253 ) , .B2( u0_n119 ) , .A( u0_n120 ) );
  OAI21_X1 u0_U276 (.B1( ld ) , .ZN( u0_N187 ) , .B2( u0_n121 ) , .A( u0_n197 ) );
  OAI21_X1 u0_U277 (.B1( ld ) , .ZN( u0_N270 ) , .B2( u0_n68 ) , .A( u0_n69 ) );
  OAI21_X1 u0_U278 (.B1( ld ) , .ZN( u0_N204 ) , .A( u0_n163 ) , .B2( u0_n70 ) );
  OAI21_X1 u0_U279 (.B1( ld ) , .ZN( u0_N124 ) , .B2( u0_n192 ) , .A( u0_n255 ) );
  NAND2_X1 u0_U28 (.A1( key[93] ) , .A2( ld ) , .ZN( u0_n229 ) );
  OAI21_X1 u0_U280 (.B1( ld ) , .ZN( u0_N190 ) , .B2( u0_n112 ) , .A( u0_n191 ) );
  OAI21_X1 u0_U281 (.B1( ld ) , .ZN( u0_N248 ) , .B2( u0_n134 ) , .A( u0_n135 ) );
  OAI21_X1 u0_U282 (.B1( ld ) , .ZN( u0_N182 ) , .B2( u0_n136 ) , .A( u0_n207 ) );
  OAI21_X1 u0_U283 (.B1( ld ) , .ZN( u0_N132 ) , .B2( u0_n176 ) , .A( u0_n239 ) );
  OAI21_X1 u0_U284 (.B1( ld ) , .ZN( u0_N198 ) , .A( u0_n175 ) , .B2( u0_n88 ) );
  OAI21_X1 u0_U285 (.B1( ld ) , .ZN( u0_N240 ) , .B2( u0_n158 ) , .A( u0_n159 ) );
  OAI21_X1 u0_U286 (.B1( ld ) , .ZN( u0_N174 ) , .B2( u0_n160 ) , .A( u0_n223 ) );
  XNOR2_X1 u0_U287 (.ZN( u0_n236 ) , .A( u0_subword_26 ) , .B( w0_26 ) );
  OAI21_X1 u0_U288 (.B1( ld ) , .ZN( u0_N52 ) , .B2( u0_n43 ) , .A( u0_n44 ) );
  OAI21_X1 u0_U289 (.B1( ld ) , .ZN( u0_N118 ) , .B2( u0_n204 ) , .A( u0_n267 ) );
  NAND2_X1 u0_U29 (.A1( key[92] ) , .A2( ld ) , .ZN( u0_n231 ) );
  OAI21_X1 u0_U290 (.B1( ld ) , .ZN( u0_N60 ) , .B2( u0_n27 ) , .A( u0_n28 ) );
  XOR2_X1 u0_U291 (.Z( u0_n65 ) , .A( u0_n67 ) , .B( w3_31 ) );
  XOR2_X1 u0_U292 (.Z( u0_n68 ) , .A( u0_n70 ) , .B( w3_30 ) );
  XOR2_X1 u0_U293 (.Z( u0_n71 ) , .A( u0_n73 ) , .B( w3_29 ) );
  XOR2_X1 u0_U294 (.Z( u0_n74 ) , .A( u0_n76 ) , .B( w3_28 ) );
  XOR2_X1 u0_U295 (.Z( u0_n77 ) , .A( u0_n79 ) , .B( w3_27 ) );
  XOR2_X1 u0_U296 (.Z( u0_n80 ) , .A( u0_n82 ) , .B( w3_26 ) );
  XOR2_X1 u0_U297 (.Z( u0_n83 ) , .A( u0_n85 ) , .B( w3_25 ) );
  OAI21_X1 u0_U298 (.B1( ld ) , .ZN( u0_N126 ) , .B2( u0_n188 ) , .A( u0_n251 ) );
  XOR2_X1 u0_U299 (.Z( u0_n89 ) , .A( u0_n91 ) , .B( w3_23 ) );
  XNOR2_X1 u0_U3 (.A( u0_n11 ) , .ZN( u0_n172 ) , .B( u0_n242 ) );
  NAND2_X1 u0_U30 (.A1( key[59] ) , .A2( ld ) , .ZN( u0_n169 ) );
  XOR2_X1 u0_U300 (.Z( u0_n92 ) , .A( u0_n94 ) , .B( w3_22 ) );
  XOR2_X1 u0_U301 (.Z( u0_n95 ) , .A( u0_n97 ) , .B( w3_21 ) );
  XOR2_X1 u0_U302 (.A( u0_n100 ) , .Z( u0_n98 ) , .B( w3_20 ) );
  XOR2_X1 u0_U303 (.Z( u0_n101 ) , .A( u0_n103 ) , .B( w3_19 ) );
  XOR2_X1 u0_U304 (.Z( u0_n104 ) , .A( u0_n106 ) , .B( w3_18 ) );
  XOR2_X1 u0_U305 (.Z( u0_n107 ) , .A( u0_n109 ) , .B( w3_17 ) );
  XOR2_X1 u0_U306 (.Z( u0_n110 ) , .A( u0_n112 ) , .B( w3_16 ) );
  XOR2_X1 u0_U307 (.Z( u0_n113 ) , .A( u0_n115 ) , .B( w3_15 ) );
  XOR2_X1 u0_U308 (.Z( u0_n116 ) , .A( u0_n118 ) , .B( w3_14 ) );
  XOR2_X1 u0_U309 (.Z( u0_n119 ) , .A( u0_n121 ) , .B( w3_13 ) );
  NAND2_X1 u0_U31 (.A1( key[53] ) , .A2( ld ) , .ZN( u0_n181 ) );
  XOR2_X1 u0_U310 (.Z( u0_n122 ) , .A( u0_n124 ) , .B( w3_12 ) );
  XOR2_X1 u0_U311 (.Z( u0_n125 ) , .A( u0_n127 ) , .B( w3_11 ) );
  XOR2_X1 u0_U312 (.Z( u0_n128 ) , .A( u0_n130 ) , .B( w3_10 ) );
  XOR2_X1 u0_U313 (.Z( u0_n131 ) , .A( u0_n133 ) , .B( w3_9 ) );
  XOR2_X1 u0_U314 (.Z( u0_n134 ) , .A( u0_n136 ) , .B( w3_8 ) );
  XOR2_X1 u0_U315 (.Z( u0_n137 ) , .A( u0_n139 ) , .B( w3_7 ) );
  XOR2_X1 u0_U316 (.Z( u0_n140 ) , .A( u0_n142 ) , .B( w3_6 ) );
  XOR2_X1 u0_U317 (.Z( u0_n143 ) , .A( u0_n145 ) , .B( w3_5 ) );
  XOR2_X1 u0_U318 (.Z( u0_n146 ) , .A( u0_n148 ) , .B( w3_4 ) );
  XOR2_X1 u0_U319 (.Z( u0_n149 ) , .A( u0_n151 ) , .B( w3_3 ) );
  NAND2_X1 u0_U32 (.A1( key[45] ) , .A2( ld ) , .ZN( u0_n197 ) );
  XOR2_X1 u0_U320 (.Z( u0_n152 ) , .A( u0_n154 ) , .B( w3_2 ) );
  XOR2_X1 u0_U321 (.Z( u0_n155 ) , .A( u0_n157 ) , .B( w3_1 ) );
  XOR2_X1 u0_U322 (.Z( u0_n158 ) , .A( u0_n160 ) , .B( w3_0 ) );
  XOR2_X1 u0_U323 (.A( u0_n162 ) , .Z( u0_n67 ) , .B( w2_31 ) );
  XOR2_X1 u0_U324 (.A( u0_n164 ) , .Z( u0_n70 ) , .B( w2_30 ) );
  XOR2_X1 u0_U325 (.A( u0_n166 ) , .Z( u0_n73 ) , .B( w2_29 ) );
  XOR2_X1 u0_U326 (.A( u0_n168 ) , .Z( u0_n76 ) , .B( w2_28 ) );
  XOR2_X1 u0_U327 (.A( u0_n170 ) , .Z( u0_n79 ) , .B( w2_27 ) );
  OAI21_X1 u0_U328 (.B1( ld ) , .ZN( u0_N68 ) , .B2( u0_n11 ) , .A( u0_n12 ) );
  XOR2_X1 u0_U329 (.A( u0_n174 ) , .Z( u0_n85 ) , .B( w2_25 ) );
  NAND2_X1 u0_U33 (.A1( key[44] ) , .A2( ld ) , .ZN( u0_n199 ) );
  XOR2_X1 u0_U330 (.A( u0_n176 ) , .Z( u0_n88 ) , .B( w2_24 ) );
  XOR2_X1 u0_U331 (.A( u0_n178 ) , .Z( u0_n91 ) , .B( w2_23 ) );
  XOR2_X1 u0_U332 (.A( u0_n180 ) , .Z( u0_n94 ) , .B( w2_22 ) );
  XOR2_X1 u0_U333 (.A( u0_n182 ) , .Z( u0_n97 ) , .B( w2_21 ) );
  XOR2_X1 u0_U334 (.Z( u0_n100 ) , .A( u0_n184 ) , .B( w2_20 ) );
  XOR2_X1 u0_U335 (.Z( u0_n103 ) , .A( u0_n186 ) , .B( w2_19 ) );
  XOR2_X1 u0_U336 (.Z( u0_n106 ) , .A( u0_n188 ) , .B( w2_18 ) );
  XOR2_X1 u0_U337 (.Z( u0_n109 ) , .A( u0_n190 ) , .B( w2_17 ) );
  XOR2_X1 u0_U338 (.Z( u0_n112 ) , .A( u0_n192 ) , .B( w2_16 ) );
  XOR2_X1 u0_U339 (.Z( u0_n115 ) , .A( u0_n194 ) , .B( w2_15 ) );
  NAND2_X1 u0_U34 (.A1( key[65] ) , .A2( ld ) , .ZN( u0_n285 ) );
  XOR2_X1 u0_U340 (.Z( u0_n118 ) , .A( u0_n196 ) , .B( w2_14 ) );
  XOR2_X1 u0_U341 (.Z( u0_n121 ) , .A( u0_n198 ) , .B( w2_13 ) );
  XOR2_X1 u0_U342 (.Z( u0_n124 ) , .A( u0_n200 ) , .B( w2_12 ) );
  XOR2_X1 u0_U343 (.Z( u0_n127 ) , .A( u0_n202 ) , .B( w2_11 ) );
  XOR2_X1 u0_U344 (.Z( u0_n130 ) , .A( u0_n204 ) , .B( w2_10 ) );
  XOR2_X1 u0_U345 (.Z( u0_n133 ) , .A( u0_n206 ) , .B( w2_9 ) );
  XOR2_X1 u0_U346 (.Z( u0_n136 ) , .A( u0_n208 ) , .B( w2_8 ) );
  XOR2_X1 u0_U347 (.Z( u0_n139 ) , .A( u0_n210 ) , .B( w2_7 ) );
  XOR2_X1 u0_U348 (.Z( u0_n142 ) , .A( u0_n212 ) , .B( w2_6 ) );
  XOR2_X1 u0_U349 (.Z( u0_n145 ) , .A( u0_n214 ) , .B( w2_5 ) );
  NAND2_X1 u0_U35 (.A1( key[68] ) , .A2( ld ) , .ZN( u0_n279 ) );
  XOR2_X1 u0_U350 (.Z( u0_n148 ) , .A( u0_n216 ) , .B( w2_4 ) );
  XOR2_X1 u0_U351 (.Z( u0_n151 ) , .A( u0_n218 ) , .B( w2_3 ) );
  XOR2_X1 u0_U352 (.Z( u0_n154 ) , .A( u0_n220 ) , .B( w2_2 ) );
  XOR2_X1 u0_U353 (.Z( u0_n157 ) , .A( u0_n222 ) , .B( w2_1 ) );
  XOR2_X1 u0_U354 (.Z( u0_n160 ) , .A( u0_n224 ) , .B( w2_0 ) );
  XOR2_X1 u0_U355 (.A( u0_n1 ) , .Z( u0_n162 ) , .B( w1_31 ) );
  XOR2_X1 u0_U356 (.Z( u0_n1 ) , .A( u0_n226 ) , .B( u0_rcon_31 ) );
  OAI21_X1 u0_U357 (.B1( ld ) , .ZN( u0_N258 ) , .B2( u0_n104 ) , .A( u0_n105 ) );
  XOR2_X1 u0_U358 (.A( u0_n228 ) , .Z( u0_n3 ) , .B( u0_rcon_30 ) );
  XOR2_X1 u0_U359 (.Z( u0_n166 ) , .A( u0_n5 ) , .B( w1_29 ) );
  NAND2_X1 u0_U36 (.A1( key[103] ) , .A2( ld ) , .ZN( u0_n50 ) );
  XOR2_X1 u0_U360 (.A( u0_n230 ) , .Z( u0_n5 ) , .B( u0_rcon_29 ) );
  XOR2_X1 u0_U361 (.Z( u0_n168 ) , .A( u0_n7 ) , .B( w1_28 ) );
  XOR2_X1 u0_U362 (.A( u0_n232 ) , .Z( u0_n7 ) , .B( u0_rcon_28 ) );
  XOR2_X1 u0_U363 (.Z( u0_n170 ) , .A( u0_n9 ) , .B( w1_27 ) );
  XOR2_X1 u0_U364 (.A( u0_n234 ) , .Z( u0_n9 ) , .B( u0_rcon_27 ) );
  OAI21_X1 u0_U365 (.B1( ld ) , .ZN( u0_N192 ) , .B2( u0_n106 ) , .A( u0_n187 ) );
  XOR2_X1 u0_U366 (.Z( u0_n11 ) , .A( u0_n236 ) , .B( u0_rcon_26 ) );
  XOR2_X1 u0_U367 (.A( u0_n13 ) , .Z( u0_n174 ) , .B( w1_25 ) );
  XOR2_X1 u0_U368 (.Z( u0_n13 ) , .A( u0_n238 ) , .B( u0_rcon_25 ) );
  XOR2_X1 u0_U369 (.A( u0_n15 ) , .Z( u0_n176 ) , .B( w1_24 ) );
  NAND2_X1 u0_U37 (.A1( key[102] ) , .A2( ld ) , .ZN( u0_n52 ) );
  OAI21_X1 u0_U370 (.B1( ld ) , .ZN( u0_N110 ) , .B2( u0_n220 ) , .A( u0_n283 ) );
  XOR2_X1 u0_U371 (.A( u0_n17 ) , .Z( u0_n178 ) , .B( w1_23 ) );
  OAI21_X1 u0_U372 (.B1( ld ) , .ZN( u0_N176 ) , .B2( u0_n154 ) , .A( u0_n219 ) );
  XOR2_X1 u0_U373 (.Z( u0_n180 ) , .A( u0_n19 ) , .B( w1_22 ) );
  OAI21_X1 u0_U374 (.B1( ld ) , .ZN( u0_N250 ) , .B2( u0_n128 ) , .A( u0_n129 ) );
  XOR2_X1 u0_U375 (.Z( u0_n182 ) , .A( u0_n21 ) , .B( w1_21 ) );
  OAI21_X1 u0_U376 (.B1( ld ) , .ZN( u0_N184 ) , .B2( u0_n130 ) , .A( u0_n203 ) );
  XOR2_X1 u0_U377 (.Z( u0_n184 ) , .A( u0_n23 ) , .B( w1_20 ) );
  OAI21_X1 u0_U378 (.B1( ld ) , .ZN( u0_N134 ) , .B2( u0_n172 ) , .A( u0_n235 ) );
  XOR2_X1 u0_U379 (.Z( u0_n186 ) , .A( u0_n25 ) , .B( w1_19 ) );
  NAND2_X1 u0_U38 (.A1( key[96] ) , .A2( ld ) , .ZN( u0_n64 ) );
  OAI21_X1 u0_U380 (.B1( ld ) , .ZN( u0_N200 ) , .A( u0_n171 ) , .B2( u0_n82 ) );
  XOR2_X1 u0_U381 (.Z( u0_n188 ) , .A( u0_n27 ) , .B( w1_18 ) );
  XOR2_X1 u0_U383 (.Z( u0_n190 ) , .A( u0_n29 ) , .B( w1_17 ) );
  XOR2_X1 u0_U385 (.Z( u0_n192 ) , .A( u0_n31 ) , .B( w1_16 ) );
  XOR2_X1 u0_U387 (.Z( u0_n194 ) , .A( u0_n33 ) , .B( w1_15 ) );
  XOR2_X1 u0_U389 (.Z( u0_n196 ) , .A( u0_n35 ) , .B( w1_14 ) );
  NAND2_X1 u0_U39 (.A1( key[115] ) , .A2( ld ) , .ZN( u0_n26 ) );
  XOR2_X1 u0_U391 (.Z( u0_n198 ) , .A( u0_n37 ) , .B( w1_13 ) );
  XOR2_X1 u0_U393 (.Z( u0_n200 ) , .A( u0_n39 ) , .B( w1_12 ) );
  XOR2_X1 u0_U395 (.Z( u0_n202 ) , .A( u0_n41 ) , .B( w1_11 ) );
  XOR2_X1 u0_U397 (.Z( u0_n204 ) , .A( u0_n43 ) , .B( w1_10 ) );
  XOR2_X1 u0_U399 (.Z( u0_n206 ) , .A( u0_n45 ) , .B( w1_9 ) );
  XNOR2_X1 u0_U4 (.A( u0_n172 ) , .B( u0_n244 ) , .ZN( u0_n82 ) );
  NAND2_X1 u0_U40 (.A1( key[114] ) , .A2( ld ) , .ZN( u0_n28 ) );
  XOR2_X1 u0_U401 (.Z( u0_n208 ) , .A( u0_n47 ) , .B( w1_8 ) );
  XOR2_X1 u0_U403 (.Z( u0_n210 ) , .A( u0_n49 ) , .B( w1_7 ) );
  XOR2_X1 u0_U405 (.Z( u0_n212 ) , .A( u0_n51 ) , .B( w1_6 ) );
  XOR2_X1 u0_U407 (.Z( u0_n214 ) , .A( u0_n53 ) , .B( w1_5 ) );
  XOR2_X1 u0_U409 (.Z( u0_n216 ) , .A( u0_n55 ) , .B( w1_4 ) );
  NAND2_X1 u0_U41 (.A1( key[112] ) , .A2( ld ) , .ZN( u0_n32 ) );
  XOR2_X1 u0_U411 (.Z( u0_n218 ) , .A( u0_n57 ) , .B( w1_3 ) );
  XOR2_X1 u0_U413 (.Z( u0_n220 ) , .A( u0_n59 ) , .B( w1_2 ) );
  XOR2_X1 u0_U415 (.Z( u0_n222 ) , .A( u0_n61 ) , .B( w1_1 ) );
  XOR2_X1 u0_U417 (.Z( u0_n224 ) , .A( u0_n63 ) , .B( w1_0 ) );
  NAND2_X1 u0_U42 (.A1( key[106] ) , .A2( ld ) , .ZN( u0_n44 ) );
  NAND2_X1 u0_U43 (.A1( key[64] ) , .A2( ld ) , .ZN( u0_n287 ) );
  NAND2_X1 u0_U44 (.A1( key[126] ) , .A2( ld ) , .ZN( u0_n4 ) );
  NAND2_X1 u0_U45 (.A1( key[23] ) , .A2( ld ) , .ZN( u0_n90 ) );
  NAND2_X1 u0_U46 (.A1( key[21] ) , .A2( ld ) , .ZN( u0_n96 ) );
  NAND2_X1 u0_U47 (.A1( key[24] ) , .A2( ld ) , .ZN( u0_n87 ) );
  NAND2_X1 u0_U48 (.A1( key[25] ) , .A2( ld ) , .ZN( u0_n84 ) );
  NAND2_X1 u0_U49 (.A1( key[122] ) , .A2( ld ) , .ZN( u0_n12 ) );
  XNOR2_X1 u0_U5 (.ZN( u0_n232 ) , .B( u0_subword_28 ) , .A( w0_28 ) );
  NAND2_X1 u0_U50 (.A1( key[118] ) , .A2( ld ) , .ZN( u0_n20 ) );
  NAND2_X1 u0_U51 (.A1( key[89] ) , .A2( ld ) , .ZN( u0_n237 ) );
  NAND2_X1 u0_U52 (.A1( key[120] ) , .A2( ld ) , .ZN( u0_n16 ) );
  NAND2_X1 u0_U53 (.A1( key[88] ) , .A2( ld ) , .ZN( u0_n239 ) );
  NAND2_X1 u0_U54 (.A1( key[86] ) , .A2( ld ) , .ZN( u0_n243 ) );
  NAND2_X1 u0_U55 (.A1( key[82] ) , .A2( ld ) , .ZN( u0_n251 ) );
  NAND2_X1 u0_U56 (.A1( key[80] ) , .A2( ld ) , .ZN( u0_n255 ) );
  NAND2_X1 u0_U57 (.A1( key[78] ) , .A2( ld ) , .ZN( u0_n259 ) );
  NAND2_X1 u0_U58 (.A1( key[26] ) , .A2( ld ) , .ZN( u0_n81 ) );
  NAND2_X1 u0_U59 (.A1( key[27] ) , .A2( ld ) , .ZN( u0_n78 ) );
  XNOR2_X1 u0_U6 (.ZN( u0_n234 ) , .B( u0_subword_27 ) , .A( w0_27 ) );
  NAND2_X1 u0_U60 (.A1( key[98] ) , .A2( ld ) , .ZN( u0_n60 ) );
  NAND2_X1 u0_U61 (.A1( key[121] ) , .A2( ld ) , .ZN( u0_n14 ) );
  NAND2_X1 u0_U62 (.A1( key[84] ) , .A2( ld ) , .ZN( u0_n247 ) );
  NAND2_X1 u0_U63 (.A1( key[83] ) , .A2( ld ) , .ZN( u0_n249 ) );
  NAND2_X1 u0_U64 (.A1( key[113] ) , .A2( ld ) , .ZN( u0_n30 ) );
  NAND2_X1 u0_U65 (.A1( key[81] ) , .A2( ld ) , .ZN( u0_n253 ) );
  NAND2_X1 u0_U66 (.A1( key[110] ) , .A2( ld ) , .ZN( u0_n36 ) );
  NAND2_X1 u0_U67 (.A1( key[75] ) , .A2( ld ) , .ZN( u0_n265 ) );
  NAND2_X1 u0_U68 (.A1( key[104] ) , .A2( ld ) , .ZN( u0_n48 ) );
  NAND2_X1 u0_U69 (.A1( key[95] ) , .A2( ld ) , .ZN( u0_n225 ) );
  XNOR2_X1 u0_U7 (.ZN( u0_n228 ) , .B( u0_subword_30 ) , .A( w0_30 ) );
  NAND2_X1 u0_U70 (.A1( key[63] ) , .A2( ld ) , .ZN( u0_n161 ) );
  NAND2_X1 u0_U71 (.A1( key[38] ) , .A2( ld ) , .ZN( u0_n211 ) );
  NAND2_X1 u0_U72 (.A1( key[36] ) , .A2( ld ) , .ZN( u0_n215 ) );
  NAND2_X1 u0_U73 (.A1( key[34] ) , .A2( ld ) , .ZN( u0_n219 ) );
  NAND2_X1 u0_U74 (.A1( key[33] ) , .A2( ld ) , .ZN( u0_n221 ) );
  NAND2_X1 u0_U75 (.A1( key[32] ) , .A2( ld ) , .ZN( u0_n223 ) );
  NAND2_X1 u0_U76 (.A1( key[94] ) , .A2( ld ) , .ZN( u0_n227 ) );
  NAND2_X1 u0_U77 (.A1( key[61] ) , .A2( ld ) , .ZN( u0_n165 ) );
  NAND2_X1 u0_U78 (.A1( key[60] ) , .A2( ld ) , .ZN( u0_n167 ) );
  NAND2_X1 u0_U79 (.A1( key[90] ) , .A2( ld ) , .ZN( u0_n235 ) );
  XNOR2_X1 u0_U8 (.ZN( u0_n238 ) , .B( u0_subword_25 ) , .A( w0_25 ) );
  NAND2_X1 u0_U80 (.A1( key[58] ) , .A2( ld ) , .ZN( u0_n171 ) );
  NAND2_X1 u0_U81 (.A1( key[57] ) , .A2( ld ) , .ZN( u0_n173 ) );
  NAND2_X1 u0_U82 (.A1( key[56] ) , .A2( ld ) , .ZN( u0_n175 ) );
  NAND2_X1 u0_U83 (.A1( key[54] ) , .A2( ld ) , .ZN( u0_n179 ) );
  NAND2_X1 u0_U84 (.A1( key[52] ) , .A2( ld ) , .ZN( u0_n183 ) );
  NAND2_X1 u0_U85 (.A1( key[51] ) , .A2( ld ) , .ZN( u0_n185 ) );
  NAND2_X1 u0_U86 (.A1( key[50] ) , .A2( ld ) , .ZN( u0_n187 ) );
  NAND2_X1 u0_U87 (.A1( key[49] ) , .A2( ld ) , .ZN( u0_n189 ) );
  NAND2_X1 u0_U88 (.A1( key[48] ) , .A2( ld ) , .ZN( u0_n191 ) );
  NAND2_X1 u0_U89 (.A1( key[46] ) , .A2( ld ) , .ZN( u0_n195 ) );
  INV_X1 u0_U9 (.ZN( u0_n246 ) , .A( u0_rcon_24 ) );
  NAND2_X1 u0_U90 (.A1( key[43] ) , .A2( ld ) , .ZN( u0_n201 ) );
  NAND2_X1 u0_U91 (.A1( key[42] ) , .A2( ld ) , .ZN( u0_n203 ) );
  NAND2_X1 u0_U92 (.A1( key[41] ) , .A2( ld ) , .ZN( u0_n205 ) );
  NAND2_X1 u0_U93 (.A1( key[40] ) , .A2( ld ) , .ZN( u0_n207 ) );
  NAND2_X1 u0_U94 (.A1( key[13] ) , .A2( ld ) , .ZN( u0_n120 ) );
  NAND2_X1 u0_U95 (.A1( key[14] ) , .A2( ld ) , .ZN( u0_n117 ) );
  NAND2_X1 u0_U96 (.A1( key[12] ) , .A2( ld ) , .ZN( u0_n123 ) );
  NAND2_X1 u0_U97 (.A1( key[7] ) , .A2( ld ) , .ZN( u0_n138 ) );
  NAND2_X1 u0_U98 (.A1( key[70] ) , .A2( ld ) , .ZN( u0_n275 ) );
  NAND2_X1 u0_U99 (.A1( key[66] ) , .A2( ld ) , .ZN( u0_n283 ) );
  OAI21_X1 u0_r0_U27 (.ZN( u0_r0_N70 ) , .B1( u0_r0_n4 ) , .B2( u0_r0_n5 ) , .A( u0_r0_n9 ) );
  NAND4_X1 u0_r0_U28 (.A3( u0_r0_N78 ) , .A2( u0_r0_n12 ) , .ZN( u0_r0_n14 ) , .A1( u0_r0_n18 ) , .A4( u0_r0_n2 ) );
  NAND2_X1 u0_r0_U29 (.A1( u0_r0_N80 ) , .ZN( u0_r0_n11 ) , .A2( u0_r0_n17 ) );
  NOR2_X1 u0_r0_U30 (.A2( ld ) , .ZN( u0_r0_N79 ) , .A1( u0_r0_n12 ) );
  NOR2_X1 u0_r0_U31 (.A2( ld ) , .ZN( u0_r0_N80 ) , .A1( u0_r0_n18 ) );
  NAND2_X1 u0_r0_U32 (.ZN( u0_r0_N71 ) , .A1( u0_r0_n10 ) , .A2( u0_r0_n23 ) );
  INV_X1 u0_r0_U33 (.A( u0_r0_n17 ) , .ZN( u0_r0_n2 ) );
  INV_X1 u0_r0_U34 (.A( u0_r0_n24 ) , .ZN( u0_r0_n5 ) );
  INV_X1 u0_r0_U35 (.A( u0_r0_n25 ) , .ZN( u0_r0_n4 ) );
  XNOR2_X1 u0_r0_U36 (.ZN( u0_r0_n12 ) , .B( u0_r0_rcnt_0 ) , .A( u0_r0_rcnt_1 ) );
  OAI21_X1 u0_r0_U37 (.B1( u0_r0_n12 ) , .A( u0_r0_n21 ) , .ZN( u0_r0_n25 ) , .B2( u0_r0_n6 ) );
  NAND4_X1 u0_r0_U38 (.ZN( u0_r0_n10 ) , .A1( u0_r0_n24 ) , .A2( u0_r0_n25 ) , .A4( u0_r0_n3 ) , .A3( u0_r0_n9 ) );
  OAI22_X1 u0_r0_U39 (.ZN( u0_r0_N73 ) , .B1( u0_r0_n16 ) , .A2( u0_r0_n19 ) , .B2( u0_r0_n20 ) , .A1( u0_r0_rcnt_0 ) );
  NAND2_X1 u0_r0_U40 (.A1( u0_r0_n12 ) , .ZN( u0_r0_n20 ) , .A2( u0_r0_rcnt_0 ) );
  NOR3_X1 u0_r0_U41 (.ZN( u0_r0_N76 ) , .A1( u0_r0_n11 ) , .A2( u0_r0_n12 ) , .A3( u0_r0_n8 ) );
  NOR3_X1 u0_r0_U42 (.ZN( u0_r0_N77 ) , .A1( u0_r0_n11 ) , .A3( u0_r0_n12 ) , .A2( u0_r0_rcnt_0 ) );
  NAND2_X1 u0_r0_U43 (.ZN( u0_r0_n21 ) , .A1( u0_r0_rcnt_0 ) , .A2( u0_r0_rcnt_1 ) );
  NOR2_X1 u0_r0_U44 (.A2( ld ) , .ZN( u0_r0_N78 ) , .A1( u0_r0_rcnt_0 ) );
  OAI21_X1 u0_r0_U45 (.ZN( u0_r0_N72 ) , .A( u0_r0_n14 ) , .B2( u0_r0_n19 ) , .B1( u0_r0_n8 ) );
  OAI21_X1 u0_r0_U46 (.ZN( u0_r0_N75 ) , .B1( u0_r0_n11 ) , .B2( u0_r0_n13 ) , .A( u0_r0_n14 ) );
  NAND2_X1 u0_r0_U47 (.A1( u0_r0_n12 ) , .ZN( u0_r0_n13 ) , .A2( u0_r0_n8 ) );
  NOR2_X1 u0_r0_U48 (.A2( u0_r0_n21 ) , .ZN( u0_r0_n22 ) , .A1( u0_r0_n6 ) );
  OAI21_X1 u0_r0_U49 (.B1( u0_r0_N70 ) , .ZN( u0_r0_N81 ) , .A( u0_r0_n10 ) , .B2( u0_r0_n3 ) );
  NAND2_X1 u0_r0_U50 (.ZN( u0_r0_N74 ) , .A2( u0_r0_n1 ) , .A1( u0_r0_n14 ) );
  INV_X1 u0_r0_U51 (.ZN( u0_r0_n1 ) , .A( u0_r0_n15 ) );
  AOI211_X1 u0_r0_U52 (.C2( u0_r0_n11 ) , .ZN( u0_r0_n15 ) , .C1( u0_r0_n16 ) , .B( u0_r0_n7 ) , .A( u0_r0_n8 ) );
  INV_X1 u0_r0_U53 (.A( u0_r0_n12 ) , .ZN( u0_r0_n7 ) );
  INV_X1 u0_r0_U54 (.A( ld ) , .ZN( u0_r0_n9 ) );
  NAND3_X1 u0_r0_U55 (.ZN( u0_r0_n16 ) , .A3( u0_r0_n18 ) , .A1( u0_r0_n2 ) , .A2( u0_r0_n9 ) );
  NAND3_X1 u0_r0_U56 (.A3( u0_r0_N79 ) , .A1( u0_r0_n17 ) , .A2( u0_r0_n18 ) , .ZN( u0_r0_n19 ) );
  XOR2_X1 u0_r0_U57 (.Z( u0_r0_n18 ) , .A( u0_r0_n21 ) , .B( u0_r0_rcnt_2 ) );
  XOR2_X1 u0_r0_U58 (.Z( u0_r0_n17 ) , .B( u0_r0_n22 ) , .A( u0_r0_n3 ) );
  NAND3_X1 u0_r0_U59 (.ZN( u0_r0_n23 ) , .A3( u0_r0_n4 ) , .A1( u0_r0_n5 ) , .A2( u0_r0_n9 ) );
  XOR2_X1 u0_r0_U60 (.B( u0_r0_n12 ) , .Z( u0_r0_n24 ) , .A( u0_r0_n6 ) );
  DFF_X1 u0_r0_out_reg_24 (.CK( clk ) , .D( u0_r0_N70 ) , .Q( u0_rcon_24 ) );
  DFF_X1 u0_r0_out_reg_25 (.CK( clk ) , .D( u0_r0_N71 ) , .Q( u0_rcon_25 ) );
  DFF_X1 u0_r0_out_reg_26 (.CK( clk ) , .D( u0_r0_N72 ) , .Q( u0_rcon_26 ) );
  DFF_X1 u0_r0_out_reg_27 (.CK( clk ) , .D( u0_r0_N73 ) , .Q( u0_rcon_27 ) );
  DFF_X1 u0_r0_out_reg_28 (.CK( clk ) , .D( u0_r0_N74 ) , .Q( u0_rcon_28 ) );
  DFF_X1 u0_r0_out_reg_29 (.CK( clk ) , .D( u0_r0_N75 ) , .Q( u0_rcon_29 ) );
  DFF_X1 u0_r0_out_reg_30 (.CK( clk ) , .D( u0_r0_N76 ) , .Q( u0_rcon_30 ) );
  DFF_X1 u0_r0_out_reg_31 (.CK( clk ) , .D( u0_r0_N77 ) , .Q( u0_rcon_31 ) );
  DFF_X1 u0_r0_rcnt_reg_0 (.CK( clk ) , .D( u0_r0_N78 ) , .QN( u0_r0_n8 ) , .Q( u0_r0_rcnt_0 ) );
  DFF_X1 u0_r0_rcnt_reg_1 (.CK( clk ) , .D( u0_r0_N79 ) , .Q( u0_r0_rcnt_1 ) );
  DFF_X1 u0_r0_rcnt_reg_2 (.CK( clk ) , .D( u0_r0_N80 ) , .QN( u0_r0_n6 ) , .Q( u0_r0_rcnt_2 ) );
  DFF_X1 u0_r0_rcnt_reg_3 (.CK( clk ) , .D( u0_r0_N81 ) , .QN( u0_r0_n3 ) );
  INV_X1 u0_u0_U10 (.A( u0_u0_n1 ) , .ZN( u0_u0_n440 ) );
  AOI22_X1 u0_u0_U100 (.A2( u0_u0_n787 ) , .ZN( u0_u0_n788 ) , .B2( u0_u0_n836 ) , .A1( u0_u0_n839 ) , .B1( u0_u0_n867 ) );
  INV_X1 u0_u0_U101 (.A( u0_u0_n767 ) , .ZN( u0_u0_n835 ) );
  NOR2_X1 u0_u0_U102 (.ZN( u0_u0_n653 ) , .A1( u0_u0_n859 ) , .A2( u0_u0_n872 ) );
  INV_X1 u0_u0_U103 (.A( u0_u0_n759 ) , .ZN( u0_u0_n873 ) );
  OAI21_X1 u0_u0_U104 (.A( u0_u0_n439 ) , .B1( u0_u0_n758 ) , .ZN( u0_u0_n759 ) , .B2( u0_u0_n872 ) );
  NOR4_X1 u0_u0_U105 (.A4( u0_u0_n671 ) , .A3( u0_u0_n672 ) , .A2( u0_u0_n673 ) , .A1( u0_u0_n674 ) , .ZN( u0_u0_n682 ) );
  NOR4_X1 u0_u0_U106 (.A4( u0_u0_n667 ) , .A3( u0_u0_n668 ) , .A2( u0_u0_n669 ) , .A1( u0_u0_n670 ) , .ZN( u0_u0_n683 ) );
  NOR2_X1 u0_u0_U107 (.ZN( u0_u0_n738 ) , .A2( u0_u0_n837 ) , .A1( u0_u0_n850 ) );
  OR4_X1 u0_u0_U108 (.ZN( u0_u0_n472 ) , .A4( u0_u0_n524 ) , .A3( u0_u0_n535 ) , .A2( u0_u0_n584 ) , .A1( u0_u0_n717 ) );
  OR4_X1 u0_u0_U109 (.A4( u0_u0_n524 ) , .A2( u0_u0_n525 ) , .A1( u0_u0_n526 ) , .ZN( u0_u0_n528 ) , .A3( u0_u0_n826 ) );
  NAND2_X2 u0_u0_U11 (.A1( u0_u0_n455 ) , .A2( u0_u0_n466 ) , .ZN( u0_u0_n797 ) );
  OR4_X1 u0_u0_U110 (.A4( u0_u0_n688 ) , .A3( u0_u0_n689 ) , .A2( u0_u0_n690 ) , .A1( u0_u0_n691 ) , .ZN( u0_u0_n696 ) );
  OR4_X1 u0_u0_U111 (.A4( u0_u0_n572 ) , .A3( u0_u0_n573 ) , .A2( u0_u0_n574 ) , .ZN( u0_u0_n578 ) , .A1( u0_u0_n671 ) );
  OR4_X1 u0_u0_U112 (.ZN( u0_u0_n498 ) , .A4( u0_u0_n540 ) , .A2( u0_u0_n553 ) , .A1( u0_u0_n565 ) , .A3( u0_u0_n638 ) );
  INV_X1 u0_u0_U113 (.A( u0_u0_n442 ) , .ZN( u0_u0_n843 ) );
  OR3_X1 u0_u0_U114 (.A3( u0_u0_n512 ) , .A2( u0_u0_n513 ) , .A1( u0_u0_n514 ) , .ZN( u0_u0_n517 ) );
  INV_X1 u0_u0_U115 (.A( u0_u0_n469 ) , .ZN( u0_u0_n868 ) );
  OAI21_X1 u0_u0_U116 (.ZN( u0_u0_n469 ) , .B1( u0_u0_n814 ) , .A( u0_u0_n839 ) , .B2( u0_u0_n856 ) );
  AOI221_X1 u0_u0_U117 (.A( u0_u0_n718 ) , .B2( u0_u0_n719 ) , .ZN( u0_u0_n725 ) , .C1( u0_u0_n837 ) , .B1( u0_u0_n844 ) , .C2( u0_u0_n867 ) );
  OR2_X1 u0_u0_U118 (.A2( u0_u0_n716 ) , .A1( u0_u0_n717 ) , .ZN( u0_u0_n718 ) );
  NOR4_X1 u0_u0_U119 (.A4( u0_u0_n504 ) , .A3( u0_u0_n505 ) , .A2( u0_u0_n506 ) , .ZN( u0_u0_n507 ) , .A1( u0_u0_n533 ) );
  NAND2_X1 u0_u0_U12 (.A1( u0_u0_n457 ) , .A2( u0_u0_n477 ) , .ZN( u0_u0_n821 ) );
  NOR4_X1 u0_u0_U120 (.A4( u0_u0_n823 ) , .A3( u0_u0_n824 ) , .A2( u0_u0_n825 ) , .A1( u0_u0_n826 ) , .ZN( u0_u0_n827 ) );
  INV_X1 u0_u0_U121 (.A( u0_u0_n754 ) , .ZN( u0_u0_n867 ) );
  AOI221_X1 u0_u0_U122 (.C1( u0_u0_n444 ) , .A( u0_u0_n769 ) , .ZN( u0_u0_n779 ) , .C2( u0_u0_n815 ) , .B2( u0_u0_n840 ) , .B1( u0_u0_n870 ) );
  INV_X1 u0_u0_U123 (.A( u0_u0_n766 ) , .ZN( u0_u0_n840 ) );
  INV_X1 u0_u0_U124 (.A( u0_u0_n735 ) , .ZN( u0_u0_n844 ) );
  INV_X1 u0_u0_U125 (.A( u0_u0_n795 ) , .ZN( u0_u0_n837 ) );
  AOI211_X1 u0_u0_U126 (.B( u0_u0_n595 ) , .A( u0_u0_n596 ) , .ZN( u0_u0_n602 ) , .C2( u0_u0_n816 ) , .C1( u0_u0_n838 ) );
  AOI211_X1 u0_u0_U127 (.A( u0_u0_n502 ) , .ZN( u0_u0_n509 ) , .B( u0_u0_n807 ) , .C2( u0_u0_n844 ) , .C1( u0_u0_n856 ) );
  OAI221_X1 u0_u0_U128 (.A( u0_u0_n732 ) , .C2( u0_u0_n733 ) , .B2( u0_u0_n734 ) , .B1( u0_u0_n735 ) , .ZN( u0_u0_n742 ) , .C1( u0_u0_n822 ) );
  AOI22_X1 u0_u0_U129 (.ZN( u0_u0_n732 ) , .B1( u0_u0_n837 ) , .A2( u0_u0_n843 ) , .A1( u0_u0_n867 ) , .B2( u0_u0_n870 ) );
  NAND2_X1 u0_u0_U13 (.A2( u0_u0_n459 ) , .A1( u0_u0_n461 ) , .ZN( u0_u0_n811 ) );
  NOR4_X1 u0_u0_U130 (.A4( u0_u0_n645 ) , .A3( u0_u0_n646 ) , .A2( u0_u0_n647 ) , .A1( u0_u0_n648 ) , .ZN( u0_u0_n649 ) );
  AOI21_X1 u0_u0_U131 (.ZN( u0_u0_n645 ) , .B2( u0_u0_n754 ) , .A( u0_u0_n793 ) , .B1( u0_u0_n817 ) );
  NOR4_X1 u0_u0_U132 (.A4( u0_u0_n798 ) , .A3( u0_u0_n799 ) , .A2( u0_u0_n800 ) , .A1( u0_u0_n801 ) , .ZN( u0_u0_n802 ) );
  OAI21_X1 u0_u0_U133 (.A( u0_u0_n792 ) , .B2( u0_u0_n793 ) , .B1( u0_u0_n794 ) , .ZN( u0_u0_n800 ) );
  OAI221_X1 u0_u0_U134 (.A( u0_u0_n788 ) , .C2( u0_u0_n789 ) , .B2( u0_u0_n790 ) , .B1( u0_u0_n791 ) , .ZN( u0_u0_n801 ) , .C1( u0_u0_n818 ) );
  NOR3_X1 u0_u0_U135 (.ZN( u0_u0_n496 ) , .A1( u0_u0_n787 ) , .A2( u0_u0_n855 ) , .A3( u0_u0_n867 ) );
  AOI211_X1 u0_u0_U136 (.B( u0_u0_n750 ) , .A( u0_u0_n751 ) , .ZN( u0_u0_n764 ) , .C1( u0_u0_n837 ) , .C2( u0_u0_n858 ) );
  AOI211_X1 u0_u0_U137 (.B( u0_u0_n700 ) , .A( u0_u0_n701 ) , .ZN( u0_u0_n711 ) , .C2( u0_u0_n836 ) , .C1( u0_u0_n856 ) );
  AOI211_X1 u0_u0_U138 (.C2( u0_u0_n444 ) , .B( u0_u0_n730 ) , .A( u0_u0_n731 ) , .ZN( u0_u0_n744 ) , .C1( u0_u0_n848 ) );
  INV_X1 u0_u0_U139 (.A( u0_u0_n793 ) , .ZN( u0_u0_n850 ) );
  NOR3_X1 u0_u0_U14 (.A3( u0_u0_n171 ) , .A1( u0_u0_n622 ) , .A2( u0_u0_n623 ) , .ZN( u0_u0_n624 ) );
  NOR2_X1 u0_u0_U140 (.ZN( u0_u0_n672 ) , .A1( u0_u0_n733 ) , .A2( u0_u0_n808 ) );
  NOR2_X1 u0_u0_U141 (.ZN( u0_u0_n576 ) , .A1( u0_u0_n733 ) , .A2( u0_u0_n811 ) );
  NOR2_X1 u0_u0_U142 (.ZN( u0_u0_n538 ) , .A2( u0_u0_n754 ) , .A1( u0_u0_n755 ) );
  NOR2_X1 u0_u0_U143 (.ZN( u0_u0_n512 ) , .A2( u0_u0_n733 ) , .A1( u0_u0_n767 ) );
  BUF_X2 u0_u0_U144 (.Z( u0_u0_n441 ) , .A( u0_u0_n796 ) );
  CLKBUF_X3 u0_u0_U145 (.Z( u0_u0_n442 ) , .A( u0_u0_n703 ) );
  NOR2_X1 u0_u0_U146 (.ZN( u0_u0_n667 ) , .A1( u0_u0_n734 ) , .A2( u0_u0_n795 ) );
  NOR2_X1 u0_u0_U147 (.ZN( u0_u0_n515 ) , .A1( u0_u0_n734 ) , .A2( u0_u0_n784 ) );
  NOR2_X1 u0_u0_U148 (.ZN( u0_u0_n673 ) , .A1( u0_u0_n755 ) , .A2( u0_u0_n820 ) );
  INV_X1 u0_u0_U149 (.A( u0_u0_n819 ) , .ZN( u0_u0_n838 ) );
  NOR3_X1 u0_u0_U15 (.A3( u0_u0_n438 ) , .A1( u0_u0_n781 ) , .ZN( u0_u0_n804 ) , .A2( u0_u0_n806 ) );
  NOR2_X1 u0_u0_U150 (.A2( u0_u0_n442 ) , .ZN( u0_u0_n668 ) , .A1( u0_u0_n734 ) );
  NOR2_X1 u0_u0_U151 (.ZN( u0_u0_n669 ) , .A1( u0_u0_n734 ) , .A2( u0_u0_n790 ) );
  NOR2_X1 u0_u0_U152 (.ZN( u0_u0_n513 ) , .A1( u0_u0_n817 ) , .A2( u0_u0_n822 ) );
  NOR2_X1 u0_u0_U153 (.ZN( u0_u0_n661 ) , .A1( u0_u0_n795 ) , .A2( u0_u0_n820 ) );
  NOR2_X1 u0_u0_U154 (.ZN( u0_u0_n551 ) , .A1( u0_u0_n754 ) , .A2( u0_u0_n819 ) );
  NOR2_X1 u0_u0_U155 (.ZN( u0_u0_n636 ) , .A1( u0_u0_n752 ) , .A2( u0_u0_n820 ) );
  NOR2_X1 u0_u0_U156 (.A1( u0_u0_n754 ) , .ZN( u0_u0_n772 ) , .A2( u0_u0_n808 ) );
  NOR2_X1 u0_u0_U157 (.A1( u0_u0_n442 ) , .ZN( u0_u0_n775 ) , .A2( u0_u0_n820 ) );
  INV_X1 u0_u0_U158 (.A( u0_u0_n752 ) , .ZN( u0_u0_n839 ) );
  INV_X1 u0_u0_U159 (.A( u0_u0_n755 ) , .ZN( u0_u0_n847 ) );
  OR4_X1 u0_u0_U16 (.A4( u0_u0_n586 ) , .A3( u0_u0_n587 ) , .A2( u0_u0_n588 ) , .A1( u0_u0_n589 ) , .ZN( u0_u0_n590 ) );
  NOR2_X1 u0_u0_U160 (.ZN( u0_u0_n621 ) , .A1( u0_u0_n790 ) , .A2( u0_u0_n820 ) );
  NOR2_X1 u0_u0_U161 (.ZN( u0_u0_n635 ) , .A2( u0_u0_n733 ) , .A1( u0_u0_n790 ) );
  NOR2_X1 u0_u0_U162 (.ZN( u0_u0_n716 ) , .A1( u0_u0_n767 ) , .A2( u0_u0_n768 ) );
  NOR2_X1 u0_u0_U163 (.A2( u0_u0_n442 ) , .ZN( u0_u0_n600 ) , .A1( u0_u0_n733 ) );
  NOR2_X1 u0_u0_U164 (.ZN( u0_u0_n620 ) , .A1( u0_u0_n767 ) , .A2( u0_u0_n817 ) );
  AOI21_X1 u0_u0_U165 (.B1( u0_u0_n631 ) , .ZN( u0_u0_n633 ) , .A( u0_u0_n768 ) , .B2( u0_u0_n819 ) );
  AOI21_X1 u0_u0_U166 (.ZN( u0_u0_n597 ) , .B2( u0_u0_n768 ) , .A( u0_u0_n790 ) , .B1( u0_u0_n817 ) );
  AOI21_X1 u0_u0_U167 (.ZN( u0_u0_n521 ) , .A( u0_u0_n734 ) , .B1( u0_u0_n755 ) , .B2( u0_u0_n808 ) );
  AOI21_X1 u0_u0_U168 (.ZN( u0_u0_n545 ) , .B2( u0_u0_n817 ) , .A( u0_u0_n819 ) , .B1( u0_u0_n820 ) );
  INV_X1 u0_u0_U169 (.A( u0_u0_n808 ) , .ZN( u0_u0_n848 ) );
  NOR2_X1 u0_u0_U17 (.A2( u0_u0_n22 ) , .A1( u0_u0_n590 ) , .ZN( u0_u0_n591 ) );
  AOI21_X1 u0_u0_U170 (.ZN( u0_u0_n546 ) , .A( u0_u0_n768 ) , .B2( u0_u0_n784 ) , .B1( u0_u0_n822 ) );
  NOR2_X1 u0_u0_U171 (.ZN( u0_u0_n574 ) , .A1( u0_u0_n734 ) , .A2( u0_u0_n767 ) );
  AOI21_X1 u0_u0_U172 (.B1( u0_u0_n692 ) , .ZN( u0_u0_n693 ) , .A( u0_u0_n733 ) , .B2( u0_u0_n766 ) );
  NOR2_X1 u0_u0_U173 (.A2( u0_u0_n442 ) , .ZN( u0_u0_n572 ) , .A1( u0_u0_n768 ) );
  INV_X1 u0_u0_U174 (.A( u0_u0_n733 ) , .ZN( u0_u0_n857 ) );
  INV_X1 u0_u0_U175 (.A( u0_u0_n734 ) , .ZN( u0_u0_n872 ) );
  AOI21_X1 u0_u0_U176 (.B2( u0_u0_n442 ) , .ZN( u0_u0_n577 ) , .B1( u0_u0_n811 ) , .A( u0_u0_n817 ) );
  NOR2_X1 u0_u0_U177 (.ZN( u0_u0_n527 ) , .A1( u0_u0_n795 ) , .A2( u0_u0_n817 ) );
  AOI21_X1 u0_u0_U178 (.ZN( u0_u0_n695 ) , .B2( u0_u0_n754 ) , .B1( u0_u0_n768 ) , .A( u0_u0_n811 ) );
  AOI21_X1 u0_u0_U179 (.B2( u0_u0_n442 ) , .ZN( u0_u0_n484 ) , .A( u0_u0_n754 ) , .B1( u0_u0_n784 ) );
  NOR3_X1 u0_u0_U18 (.A3( u0_u0_n805 ) , .A2( u0_u0_n806 ) , .A1( u0_u0_n807 ) , .ZN( u0_u0_n830 ) );
  INV_X1 u0_u0_U180 (.A( u0_u0_n817 ) , .ZN( u0_u0_n859 ) );
  INV_X1 u0_u0_U181 (.A( u0_u0_n811 ) , .ZN( u0_u0_n846 ) );
  INV_X1 u0_u0_U182 (.A( u0_u0_n768 ) , .ZN( u0_u0_n870 ) );
  OAI21_X1 u0_u0_U183 (.A( u0_u0_n704 ) , .ZN( u0_u0_n708 ) , .B2( u0_u0_n755 ) , .B1( u0_u0_n809 ) );
  OAI21_X1 u0_u0_U184 (.ZN( u0_u0_n704 ) , .B2( u0_u0_n838 ) , .B1( u0_u0_n843 ) , .A( u0_u0_n864 ) );
  NOR2_X1 u0_u0_U185 (.ZN( u0_u0_n476 ) , .A2( u0_u0_n784 ) , .A1( u0_u0_n820 ) );
  NAND2_X1 u0_u0_U186 (.A2( u0_u0_n767 ) , .A1( u0_u0_n811 ) , .ZN( u0_u0_n815 ) );
  BUF_X1 u0_u0_U187 (.Z( u0_u0_n443 ) , .A( u0_u0_n818 ) );
  INV_X1 u0_u0_U188 (.A( u0_u0_n790 ) , .ZN( u0_u0_n851 ) );
  INV_X1 u0_u0_U189 (.A( u0_u0_n822 ) , .ZN( u0_u0_n849 ) );
  NOR3_X1 u0_u0_U19 (.ZN( u0_u0_n604 ) , .A1( u0_u0_n614 ) , .A3( u0_u0_n728 ) , .A2( u0_u0_n747 ) );
  OAI22_X1 u0_u0_U190 (.B2( u0_u0_n755 ) , .B1( u0_u0_n756 ) , .A1( u0_u0_n757 ) , .ZN( u0_u0_n761 ) , .A2( u0_u0_n811 ) );
  NOR3_X1 u0_u0_U191 (.ZN( u0_u0_n757 ) , .A2( u0_u0_n858 ) , .A1( u0_u0_n867 ) , .A3( u0_u0_n869 ) );
  NOR2_X1 u0_u0_U192 (.ZN( u0_u0_n756 ) , .A2( u0_u0_n857 ) , .A1( u0_u0_n864 ) );
  AND2_X1 u0_u0_U193 (.ZN( u0_u0_n753 ) , .A1( u0_u0_n789 ) , .A2( u0_u0_n791 ) );
  AND2_X1 u0_u0_U194 (.ZN( u0_u0_n737 ) , .A1( u0_u0_n784 ) , .A2( u0_u0_n790 ) );
  AOI221_X1 u0_u0_U195 (.A( u0_u0_n503 ) , .ZN( u0_u0_n508 ) , .B2( u0_u0_n848 ) , .C1( u0_u0_n851 ) , .C2( u0_u0_n864 ) , .B1( u0_u0_n866 ) );
  AOI221_X1 u0_u0_U196 (.A( u0_u0_n687 ) , .ZN( u0_u0_n698 ) , .B2( u0_u0_n845 ) , .C1( u0_u0_n847 ) , .C2( u0_u0_n866 ) , .B1( u0_u0_n869 ) );
  INV_X1 u0_u0_U197 (.A( u0_u0_n686 ) , .ZN( u0_u0_n845 ) );
  OAI221_X1 u0_u0_U198 (.A( u0_u0_n702 ) , .ZN( u0_u0_n709 ) , .C2( u0_u0_n789 ) , .C1( u0_u0_n790 ) , .B1( u0_u0_n791 ) , .B2( u0_u0_n811 ) );
  AOI22_X1 u0_u0_U199 (.ZN( u0_u0_n702 ) , .A1( u0_u0_n835 ) , .B2( u0_u0_n848 ) , .A2( u0_u0_n869 ) , .B1( u0_u0_n872 ) );
  NOR3_X1 u0_u0_U20 (.A1( u0_u0_n1 ) , .ZN( u0_u0_n510 ) , .A2( u0_u0_n685 ) , .A3( u0_u0_n782 ) );
  OAI222_X1 u0_u0_U200 (.A2( u0_u0_n675 ) , .ZN( u0_u0_n680 ) , .B1( u0_u0_n752 ) , .B2( u0_u0_n789 ) , .C2( u0_u0_n793 ) , .C1( u0_u0_n820 ) , .A1( u0_u0_n822 ) );
  NAND2_X1 u0_u0_U201 (.A2( u0_u0_n454 ) , .A1( u0_u0_n466 ) , .ZN( u0_u0_n733 ) );
  NAND2_X1 u0_u0_U202 (.A2( u0_u0_n454 ) , .A1( u0_u0_n458 ) , .ZN( u0_u0_n734 ) );
  NAND2_X1 u0_u0_U203 (.A2( u0_u0_n455 ) , .A1( u0_u0_n458 ) , .ZN( u0_u0_n768 ) );
  NAND2_X1 u0_u0_U204 (.A2( u0_u0_n454 ) , .A1( u0_u0_n470 ) , .ZN( u0_u0_n820 ) );
  NAND2_X1 u0_u0_U205 (.A2( u0_u0_n466 ) , .A1( u0_u0_n471 ) , .ZN( u0_u0_n785 ) );
  NAND2_X1 u0_u0_U206 (.A1( u0_u0_n453 ) , .A2( u0_u0_n471 ) , .ZN( u0_u0_n754 ) );
  NOR2_X1 u0_u0_U207 (.ZN( u0_u0_n471 ) , .A2( u0_u0_n852 ) , .A1( u0_u0_n853 ) );
  NAND2_X1 u0_u0_U208 (.A2( u0_u0_n467 ) , .A1( u0_u0_n468 ) , .ZN( u0_u0_n752 ) );
  NAND2_X1 u0_u0_U209 (.A1( u0_u0_n468 ) , .A2( u0_u0_n478 ) , .ZN( u0_u0_n793 ) );
  NOR3_X1 u0_u0_U21 (.A2( u0_u0_n613 ) , .A1( u0_u0_n614 ) , .ZN( u0_u0_n652 ) , .A3( u0_u0_n727 ) );
  NOR4_X1 u0_u0_U210 (.A4( u0_u0_n739 ) , .A3( u0_u0_n740 ) , .A2( u0_u0_n741 ) , .A1( u0_u0_n742 ) , .ZN( u0_u0_n743 ) );
  NOR4_X1 u0_u0_U211 (.A4( u0_u0_n706 ) , .A3( u0_u0_n707 ) , .A2( u0_u0_n708 ) , .A1( u0_u0_n709 ) , .ZN( u0_u0_n710 ) );
  NOR4_X1 u0_u0_U212 (.A3( u0_u0_n760 ) , .A2( u0_u0_n761 ) , .A1( u0_u0_n762 ) , .ZN( u0_u0_n763 ) , .A4( u0_u0_n873 ) );
  NOR2_X1 u0_u0_U213 (.ZN( u0_u0_n477 ) , .A1( u0_u0_n831 ) , .A2( w3_17 ) );
  AOI221_X1 u0_u0_U214 (.A( u0_u0_n786 ) , .ZN( u0_u0_n803 ) , .C2( u0_u0_n842 ) , .B2( u0_u0_n843 ) , .B1( u0_u0_n869 ) , .C1( u0_u0_n870 ) );
  NAND4_X1 u0_u0_U215 (.ZN( u0_subword_25 ) , .A4( u0_u0_n601 ) , .A3( u0_u0_n602 ) , .A2( u0_u0_n603 ) , .A1( u0_u0_n604 ) );
  NOR4_X1 u0_u0_U216 (.A4( u0_u0_n597 ) , .A3( u0_u0_n598 ) , .A2( u0_u0_n599 ) , .A1( u0_u0_n600 ) , .ZN( u0_u0_n601 ) );
  NAND4_X1 u0_u0_U217 (.ZN( u0_subword_24 ) , .A4( u0_u0_n507 ) , .A3( u0_u0_n508 ) , .A2( u0_u0_n509 ) , .A1( u0_u0_n510 ) );
  AOI222_X1 u0_u0_U218 (.B2( u0_u0_n644 ) , .ZN( u0_u0_n650 ) , .B1( u0_u0_n846 ) , .A1( u0_u0_n847 ) , .C2( u0_u0_n851 ) , .C1( u0_u0_n867 ) , .A2( u0_u0_n869 ) );
  AND2_X1 u0_u0_U219 (.ZN( u0_u0_n453 ) , .A2( w3_22 ) , .A1( w3_23 ) );
  NOR3_X1 u0_u0_U22 (.A3( u0_u0_n746 ) , .A2( u0_u0_n747 ) , .A1( u0_u0_n748 ) , .ZN( u0_u0_n765 ) );
  NAND4_X1 u0_u0_U220 (.ZN( u0_subword_31 ) , .A4( u0_u0_n827 ) , .A3( u0_u0_n828 ) , .A2( u0_u0_n829 ) , .A1( u0_u0_n830 ) );
  AOI222_X1 u0_u0_U221 (.C2( u0_u0_n814 ) , .B2( u0_u0_n815 ) , .A2( u0_u0_n816 ) , .ZN( u0_u0_n828 ) , .C1( u0_u0_n837 ) , .A1( u0_u0_n844 ) , .B1( u0_u0_n858 ) );
  INV_X1 u0_u0_U222 (.ZN( u0_u0_n853 ) , .A( w3_21 ) );
  NAND4_X1 u0_u0_U223 (.A4( u0_u0_n697 ) , .A3( u0_u0_n698 ) , .A1( u0_u0_n699 ) , .ZN( u0_u0_n781 ) , .A2( u0_u0_n876 ) );
  NAND2_X2 u0_u0_U224 (.A2( u0_u0_n470 ) , .A1( u0_u0_n471 ) , .ZN( u0_u0_n817 ) );
  NAND2_X1 u0_u0_U225 (.A2( u0_u0_n447 ) , .A1( u0_u0_n458 ) , .ZN( u0_u0_n796 ) );
  AOI222_X1 u0_u0_U226 (.ZN( u0_u0_n780 ) , .A1( u0_u0_n835 ) , .C1( u0_u0_n839 ) , .B2( u0_u0_n846 ) , .A2( u0_u0_n855 ) , .B1( u0_u0_n865 ) , .C2( u0_u0_n877 ) );
  OAI21_X1 u0_u0_U227 (.ZN( u0_u0_n736 ) , .A( u0_u0_n838 ) , .B2( u0_u0_n857 ) , .B1( u0_u0_n877 ) );
  AOI222_X1 u0_u0_U228 (.ZN( u0_u0_n569 ) , .B1( u0_u0_n835 ) , .C1( u0_u0_n846 ) , .A2( u0_u0_n848 ) , .A1( u0_u0_n859 ) , .B2( u0_u0_n867 ) , .C2( u0_u0_n877 ) );
  OAI21_X1 u0_u0_U229 (.ZN( u0_u0_n792 ) , .A( u0_u0_n844 ) , .B1( u0_u0_n867 ) , .B2( u0_u0_n877 ) );
  NOR3_X1 u0_u0_U23 (.A3( u0_u0_n727 ) , .A1( u0_u0_n728 ) , .ZN( u0_u0_n745 ) , .A2( u0_u0_n746 ) );
  NAND4_X1 u0_u0_U230 (.A4( u0_u0_n479 ) , .A3( u0_u0_n480 ) , .A2( u0_u0_n481 ) , .A1( u0_u0_n482 ) , .ZN( u0_u0_n684 ) );
  NOR4_X1 u0_u0_U231 (.ZN( u0_u0_n479 ) , .A2( u0_u0_n527 ) , .A4( u0_u0_n600 ) , .A1( u0_u0_n615 ) , .A3( u0_u0_n635 ) );
  NAND2_X1 u0_u0_U232 (.A2( u0_u0_n467 ) , .A1( u0_u0_n477 ) , .ZN( u0_u0_n703 ) );
  NAND2_X1 u0_u0_U233 (.A2( u0_u0_n460 ) , .A1( u0_u0_n461 ) , .ZN( u0_u0_n735 ) );
  NAND2_X1 u0_u0_U234 (.A1( u0_u0_n460 ) , .A2( u0_u0_n467 ) , .ZN( u0_u0_n818 ) );
  NOR2_X1 u0_u0_U235 (.ZN( u0_u0_n461 ) , .A1( u0_u0_n833 ) , .A2( w3_19 ) );
  NAND2_X2 u0_u0_U236 (.A1( u0_u0_n457 ) , .A2( u0_u0_n460 ) , .ZN( u0_u0_n819 ) );
  AOI211_X1 u0_u0_U237 (.B( u0_u0_n812 ) , .A( u0_u0_n813 ) , .ZN( u0_u0_n829 ) , .C1( u0_u0_n847 ) , .C2( u0_u0_n855 ) );
  NOR2_X1 u0_u0_U238 (.A1( u0_u0_n684 ) , .ZN( u0_u0_n699 ) , .A2( u0_u0_n812 ) );
  OAI222_X1 u0_u0_U239 (.B1( u0_u0_n442 ) , .ZN( u0_u0_n623 ) , .C1( u0_u0_n729 ) , .C2( u0_u0_n752 ) , .B2( u0_u0_n791 ) , .A2( u0_u0_n797 ) , .A1( u0_u0_n821 ) );
  NOR2_X1 u0_u0_U24 (.ZN( u0_u0_n581 ) , .A1( u0_u0_n628 ) , .A2( u0_u0_n750 ) );
  AOI21_X1 u0_u0_U240 (.A( u0_u0_n676 ) , .B1( u0_u0_n677 ) , .ZN( u0_u0_n678 ) , .B2( u0_u0_n860 ) );
  AOI21_X1 u0_u0_U241 (.B1( u0_u0_n445 ) , .ZN( u0_u0_n516 ) , .B2( u0_u0_n675 ) , .A( u0_u0_n735 ) );
  INV_X1 u0_u0_U242 (.A( u0_u0_n675 ) , .ZN( u0_u0_n869 ) );
  NOR2_X1 u0_u0_U243 (.ZN( u0_u0_n658 ) , .A1( u0_u0_n675 ) , .A2( u0_u0_n819 ) );
  NOR2_X1 u0_u0_U244 (.ZN( u0_u0_n533 ) , .A1( u0_u0_n675 ) , .A2( u0_u0_n784 ) );
  AOI21_X1 u0_u0_U245 (.ZN( u0_u0_n483 ) , .A( u0_u0_n675 ) , .B1( u0_u0_n755 ) , .B2( u0_u0_n811 ) );
  NOR2_X1 u0_u0_U246 (.ZN( u0_u0_n608 ) , .A1( u0_u0_n675 ) , .A2( u0_u0_n808 ) );
  NOR2_X1 u0_u0_U247 (.ZN( u0_u0_n634 ) , .A2( u0_u0_n675 ) , .A1( u0_u0_n790 ) );
  NOR2_X1 u0_u0_U248 (.ZN( u0_u0_n587 ) , .A1( u0_u0_n675 ) , .A2( u0_u0_n793 ) );
  NAND2_X2 u0_u0_U249 (.A1( u0_u0_n458 ) , .A2( u0_u0_n471 ) , .ZN( u0_u0_n675 ) );
  NOR2_X1 u0_u0_U25 (.ZN( u0_u0_n501 ) , .A1( u0_u0_n684 ) , .A2( u0_u0_n700 ) );
  NAND4_X1 u0_u0_U250 (.A4( u0_u0_n541 ) , .A3( u0_u0_n542 ) , .A2( u0_u0_n543 ) , .A1( u0_u0_n544 ) , .ZN( u0_u0_n628 ) );
  OAI222_X1 u0_u0_U251 (.A2( u0_u0_n445 ) , .B2( u0_u0_n713 ) , .ZN( u0_u0_n714 ) , .C2( u0_u0_n729 ) , .B1( u0_u0_n752 ) , .A1( u0_u0_n811 ) , .C1( u0_u0_n819 ) );
  NOR2_X1 u0_u0_U252 (.ZN( u0_u0_n524 ) , .A1( u0_u0_n713 ) , .A2( u0_u0_n793 ) );
  NOR2_X1 u0_u0_U253 (.ZN( u0_u0_n526 ) , .A2( u0_u0_n713 ) , .A1( u0_u0_n819 ) );
  NOR2_X1 u0_u0_U254 (.A2( u0_u0_n713 ) , .A1( u0_u0_n767 ) , .ZN( u0_u0_n799 ) );
  NOR2_X1 u0_u0_U255 (.A2( u0_u0_n713 ) , .A1( u0_u0_n755 ) , .ZN( u0_u0_n776 ) );
  NOR2_X1 u0_u0_U256 (.ZN( u0_u0_n523 ) , .A1( u0_u0_n713 ) , .A2( u0_u0_n808 ) );
  NOR2_X1 u0_u0_U257 (.ZN( u0_u0_n688 ) , .A2( u0_u0_n713 ) , .A1( u0_u0_n822 ) );
  OAI22_X1 u0_u0_U258 (.ZN( u0_u0_n489 ) , .A1( u0_u0_n713 ) , .B2( u0_u0_n790 ) , .A2( u0_u0_n811 ) , .B1( u0_u0_n817 ) );
  NOR2_X1 u0_u0_U259 (.ZN( u0_u0_n549 ) , .A2( u0_u0_n713 ) , .A1( u0_u0_n790 ) );
  NOR2_X1 u0_u0_U26 (.ZN( u0_u0_n712 ) , .A2( u0_u0_n781 ) , .A1( u0_u0_n805 ) );
  NOR2_X1 u0_u0_U260 (.ZN( u0_u0_n585 ) , .A2( u0_u0_n713 ) , .A1( u0_u0_n735 ) );
  NOR2_X1 u0_u0_U261 (.ZN( u0_u0_n535 ) , .A1( u0_u0_n713 ) , .A2( u0_u0_n784 ) );
  NOR2_X1 u0_u0_U262 (.ZN( u0_u0_n674 ) , .A2( u0_u0_n713 ) , .A1( u0_u0_n795 ) );
  AOI222_X1 u0_u0_U263 (.ZN( u0_u0_n531 ) , .A1( u0_u0_n839 ) , .B2( u0_u0_n842 ) , .C1( u0_u0_n849 ) , .C2( u0_u0_n855 ) , .A2( u0_u0_n857 ) , .B1( u0_u0_n870 ) );
  AOI222_X1 u0_u0_U264 (.ZN( u0_u0_n612 ) , .A1( u0_u0_n835 ) , .C2( u0_u0_n842 ) , .B1( u0_u0_n847 ) , .A2( u0_u0_n860 ) , .B2( u0_u0_n865 ) , .C1( u0_u0_n872 ) );
  NOR3_X1 u0_u0_U265 (.ZN( u0_u0_n446 ) , .A2( u0_u0_n841 ) , .A3( u0_u0_n842 ) , .A1( u0_u0_n851 ) );
  NAND2_X1 u0_u0_U266 (.ZN( u0_u0_n619 ) , .A2( u0_u0_n842 ) , .A1( u0_u0_n877 ) );
  OAI22_X1 u0_u0_U267 (.A1( u0_u0_n445 ) , .B2( u0_u0_n784 ) , .B1( u0_u0_n785 ) , .ZN( u0_u0_n786 ) , .A2( u0_u0_n819 ) );
  NAND4_X1 u0_u0_U268 (.A4( u0_u0_n499 ) , .A3( u0_u0_n500 ) , .A1( u0_u0_n501 ) , .ZN( u0_u0_n807 ) , .A2( u0_u0_n871 ) );
  AOI21_X1 u0_u0_U269 (.ZN( u0_u0_n575 ) , .B1( u0_u0_n755 ) , .B2( u0_u0_n767 ) , .A( u0_u0_n785 ) );
  AOI222_X1 u0_u0_U27 (.ZN( u0_u0_n666 ) , .A2( u0_u0_n844 ) , .B1( u0_u0_n846 ) , .C2( u0_u0_n850 ) , .A1( u0_u0_n864 ) , .C1( u0_u0_n867 ) , .B2( u0_u0_n874 ) );
  NAND2_X1 u0_u0_U270 (.ZN( u0_u0_n719 ) , .A1( u0_u0_n733 ) , .A2( u0_u0_n785 ) );
  OAI22_X1 u0_u0_U271 (.B1( u0_u0_n496 ) , .ZN( u0_u0_n497 ) , .A1( u0_u0_n692 ) , .A2( u0_u0_n768 ) , .B2( u0_u0_n822 ) );
  NOR2_X1 u0_u0_U272 (.ZN( u0_u0_n662 ) , .A1( u0_u0_n752 ) , .A2( u0_u0_n785 ) );
  NOR2_X1 u0_u0_U273 (.A2( u0_u0_n442 ) , .A1( u0_u0_n785 ) , .ZN( u0_u0_n825 ) );
  NOR2_X1 u0_u0_U274 (.ZN( u0_u0_n514 ) , .A2( u0_u0_n785 ) , .A1( u0_u0_n790 ) );
  NOR2_X1 u0_u0_U275 (.ZN( u0_u0_n607 ) , .A2( u0_u0_n785 ) , .A1( u0_u0_n808 ) );
  NOR2_X1 u0_u0_U276 (.ZN( u0_u0_n617 ) , .A2( u0_u0_n785 ) , .A1( u0_u0_n811 ) );
  NOR2_X1 u0_u0_U277 (.ZN( u0_u0_n552 ) , .A2( u0_u0_n785 ) , .A1( u0_u0_n819 ) );
  INV_X1 u0_u0_U278 (.A( u0_u0_n785 ) , .ZN( u0_u0_n855 ) );
  AOI21_X1 u0_u0_U279 (.ZN( u0_u0_n646 ) , .B2( u0_u0_n752 ) , .A( u0_u0_n797 ) , .B1( u0_u0_n808 ) );
  INV_X1 u0_u0_U28 (.A( u0_u0_n653 ) , .ZN( u0_u0_n874 ) );
  AOI21_X1 u0_u0_U280 (.A( u0_u0_n738 ) , .ZN( u0_u0_n739 ) , .B2( u0_u0_n785 ) , .B1( u0_u0_n797 ) );
  NAND4_X1 u0_u0_U281 (.A4( u0_u0_n554 ) , .A3( u0_u0_n555 ) , .A2( u0_u0_n556 ) , .A1( u0_u0_n557 ) , .ZN( u0_u0_n750 ) );
  AOI21_X1 u0_u0_U282 (.ZN( u0_u0_n520 ) , .A( u0_u0_n784 ) , .B2( u0_u0_n797 ) , .B1( u0_u0_n817 ) );
  AOI21_X1 u0_u0_U283 (.B2( u0_u0_n768 ) , .ZN( u0_u0_n769 ) , .A( u0_u0_n793 ) , .B1( u0_u0_n797 ) );
  AOI21_X1 u0_u0_U284 (.ZN( u0_u0_n456 ) , .B2( u0_u0_n797 ) , .A( u0_u0_n808 ) , .B1( u0_u0_n820 ) );
  INV_X1 u0_u0_U285 (.A( u0_u0_n797 ) , .ZN( u0_u0_n856 ) );
  NOR2_X1 u0_u0_U286 (.A2( u0_u0_n442 ) , .ZN( u0_u0_n721 ) , .A1( u0_u0_n797 ) );
  NOR2_X1 u0_u0_U287 (.ZN( u0_u0_n563 ) , .A1( u0_u0_n797 ) , .A2( u0_u0_n819 ) );
  NOR2_X1 u0_u0_U288 (.ZN( u0_u0_n589 ) , .A1( u0_u0_n797 ) , .A2( u0_u0_n822 ) );
  NOR2_X1 u0_u0_U289 (.ZN( u0_u0_n550 ) , .A2( u0_u0_n790 ) , .A1( u0_u0_n797 ) );
  NOR4_X1 u0_u0_U29 (.ZN( u0_u0_n491 ) , .A2( u0_u0_n539 ) , .A1( u0_u0_n564 ) , .A3( u0_u0_n637 ) , .A4( u0_u0_n723 ) );
  INV_X1 u0_u0_U290 (.ZN( u0_u0_n444 ) , .A( u0_u0_n820 ) );
  INV_X1 u0_u0_U291 (.A( u0_u0_n444 ) , .ZN( u0_u0_n445 ) );
  NOR4_X1 u0_u0_U292 (.A2( u0_u0_n497 ) , .A1( u0_u0_n498 ) , .ZN( u0_u0_n499 ) , .A3( u0_u0_n586 ) , .A4( u0_u0_n618 ) );
  INV_X1 u0_u0_U293 (.ZN( u0_u0_n832 ) , .A( w3_17 ) );
  AOI21_X1 u0_u0_U294 (.B1( u0_u0_n445 ) , .ZN( u0_u0_n595 ) , .B2( u0_u0_n705 ) , .A( u0_u0_n822 ) );
  AOI21_X1 u0_u0_U295 (.B1( u0_u0_n705 ) , .ZN( u0_u0_n706 ) , .A( u0_u0_n737 ) , .B2( u0_u0_n768 ) );
  INV_X1 u0_u0_U296 (.A( u0_u0_n705 ) , .ZN( u0_u0_n858 ) );
  AOI21_X1 u0_u0_U297 (.ZN( u0_u0_n448 ) , .A( u0_u0_n705 ) , .B1( u0_u0_n738 ) , .B2( u0_u0_n755 ) );
  NOR2_X1 u0_u0_U298 (.ZN( u0_u0_n583 ) , .A2( u0_u0_n705 ) , .A1( u0_u0_n819 ) );
  NOR2_X1 u0_u0_U299 (.ZN( u0_u0_n689 ) , .A2( u0_u0_n705 ) , .A1( u0_u0_n808 ) );
  OR4_X1 u0_u0_U3 (.ZN( u0_u0_n1 ) , .A4( u0_u0_n451 ) , .A3( u0_u0_n452 ) , .A2( u0_u0_n522 ) , .A1( u0_u0_n547 ) );
  NOR4_X1 u0_u0_U30 (.ZN( u0_u0_n485 ) , .A1( u0_u0_n526 ) , .A4( u0_u0_n563 ) , .A3( u0_u0_n588 ) , .A2( u0_u0_n636 ) );
  NOR2_X1 u0_u0_U300 (.A2( u0_u0_n442 ) , .ZN( u0_u0_n547 ) , .A1( u0_u0_n705 ) );
  NAND2_X1 u0_u0_U301 (.A1( u0_u0_n705 ) , .A2( u0_u0_n734 ) , .ZN( u0_u0_n787 ) );
  NAND2_X2 u0_u0_U302 (.A1( u0_u0_n447 ) , .A2( u0_u0_n466 ) , .ZN( u0_u0_n705 ) );
  NOR4_X1 u0_u0_U303 (.A3( u0_u0_n679 ) , .A1( u0_u0_n680 ) , .ZN( u0_u0_n681 ) , .A4( u0_u0_n720 ) , .A2( u0_u0_n863 ) );
  INV_X1 u0_u0_U304 (.A( u0_u0_n678 ) , .ZN( u0_u0_n863 ) );
  NOR2_X1 u0_u0_U305 (.ZN( u0_u0_n459 ) , .A1( u0_u0_n831 ) , .A2( u0_u0_n832 ) );
  AOI21_X1 u0_u0_U306 (.ZN( u0_u0_n504 ) , .A( u0_u0_n729 ) , .B2( u0_u0_n767 ) , .B1( u0_u0_n819 ) );
  OAI22_X1 u0_u0_U307 (.ZN( u0_u0_n495 ) , .A1( u0_u0_n729 ) , .B2( u0_u0_n733 ) , .B1( u0_u0_n735 ) , .A2( u0_u0_n784 ) );
  NOR2_X1 u0_u0_U308 (.ZN( u0_u0_n717 ) , .A2( u0_u0_n729 ) , .A1( u0_u0_n795 ) );
  NOR2_X1 u0_u0_U309 (.ZN( u0_u0_n534 ) , .A2( u0_u0_n729 ) , .A1( u0_u0_n808 ) );
  NOR4_X1 u0_u0_U31 (.ZN( u0_u0_n462 ) , .A2( u0_u0_n523 ) , .A1( u0_u0_n549 ) , .A3( u0_u0_n585 ) , .A4( u0_u0_n621 ) );
  NOR2_X1 u0_u0_U310 (.ZN( u0_u0_n532 ) , .A1( u0_u0_n729 ) , .A2( u0_u0_n755 ) );
  NOR2_X1 u0_u0_U311 (.ZN( u0_u0_n615 ) , .A2( u0_u0_n729 ) , .A1( u0_u0_n822 ) );
  NOR2_X1 u0_u0_U312 (.A2( u0_u0_n442 ) , .ZN( u0_u0_n638 ) , .A1( u0_u0_n729 ) );
  NOR2_X1 u0_u0_U313 (.ZN( u0_u0_n540 ) , .A1( u0_u0_n729 ) , .A2( u0_u0_n793 ) );
  NOR2_X1 u0_u0_U314 (.ZN( u0_u0_n539 ) , .A2( u0_u0_n729 ) , .A1( u0_u0_n735 ) );
  INV_X1 u0_u0_U315 (.A( u0_u0_n729 ) , .ZN( u0_u0_n860 ) );
  NAND2_X2 u0_u0_U316 (.A1( u0_u0_n447 ) , .A2( u0_u0_n470 ) , .ZN( u0_u0_n713 ) );
  NAND2_X2 u0_u0_U317 (.A1( u0_u0_n455 ) , .A2( u0_u0_n470 ) , .ZN( u0_u0_n729 ) );
  AOI211_X1 u0_u0_U318 (.C1( u0_u0_n439 ) , .C2( u0_u0_n444 ) , .A( u0_u0_n594 ) , .ZN( u0_u0_n603 ) , .B( u0_u0_n627 ) );
  NOR3_X1 u0_u0_U319 (.A2( u0_u0_n627 ) , .A3( u0_u0_n628 ) , .ZN( u0_u0_n642 ) , .A1( u0_u0_n730 ) );
  OR3_X1 u0_u0_U32 (.ZN( u0_u0_n452 ) , .A1( u0_u0_n534 ) , .A3( u0_u0_n583 ) , .A2( u0_u0_n879 ) );
  AOI21_X1 u0_u0_U320 (.B2( u0_u0_n443 ) , .ZN( u0_u0_n599 ) , .B1( u0_u0_n755 ) , .A( u0_u0_n797 ) );
  AOI21_X1 u0_u0_U321 (.A( u0_u0_n817 ) , .B2( u0_u0_n818 ) , .B1( u0_u0_n819 ) , .ZN( u0_u0_n824 ) );
  AOI21_X1 u0_u0_U322 (.A( u0_u0_n443 ) , .ZN( u0_u0_n655 ) , .B1( u0_u0_n734 ) , .B2( u0_u0_n768 ) );
  NOR2_X1 u0_u0_U323 (.A2( u0_u0_n818 ) , .A1( u0_u0_n820 ) , .ZN( u0_u0_n826 ) );
  NOR2_X1 u0_u0_U324 (.A2( u0_u0_n443 ) , .A1( u0_u0_n675 ) , .ZN( u0_u0_n771 ) );
  NOR2_X1 u0_u0_U325 (.ZN( u0_u0_n584 ) , .A1( u0_u0_n713 ) , .A2( u0_u0_n818 ) );
  NOR2_X1 u0_u0_U326 (.ZN( u0_u0_n671 ) , .A1( u0_u0_n785 ) , .A2( u0_u0_n818 ) );
  NAND2_X2 u0_u0_U327 (.A2( u0_u0_n460 ) , .A1( u0_u0_n478 ) , .ZN( u0_u0_n784 ) );
  NOR2_X1 u0_u0_U328 (.A1( u0_u0_n705 ) , .ZN( u0_u0_n773 ) , .A2( u0_u0_n818 ) );
  NOR2_X1 u0_u0_U329 (.A2( u0_u0_n443 ) , .ZN( u0_u0_n660 ) , .A1( u0_u0_n733 ) );
  INV_X1 u0_u0_U33 (.A( u0_u0_n619 ) , .ZN( u0_u0_n879 ) );
  NOR2_X1 u0_u0_U330 (.A2( u0_u0_n443 ) , .ZN( u0_u0_n637 ) , .A1( u0_u0_n729 ) );
  INV_X1 u0_u0_U331 (.A( u0_u0_n818 ) , .ZN( u0_u0_n841 ) );
  NAND2_X2 u0_u0_U332 (.A1( u0_u0_n457 ) , .A2( u0_u0_n459 ) , .ZN( u0_u0_n767 ) );
  NOR2_X1 u0_u0_U333 (.ZN( u0_u0_n478 ) , .A1( w3_18 ) , .A2( w3_19 ) );
  AOI21_X1 u0_u0_U334 (.A( u0_u0_n441 ) , .ZN( u0_u0_n647 ) , .B1( u0_u0_n686 ) , .B2( u0_u0_n822 ) );
  NAND2_X2 u0_u0_U335 (.A1( u0_u0_n453 ) , .A2( u0_u0_n455 ) , .ZN( u0_u0_n810 ) );
  AOI21_X1 u0_u0_U336 (.B2( u0_u0_n441 ) , .A( u0_u0_n795 ) , .B1( u0_u0_n797 ) , .ZN( u0_u0_n798 ) );
  OAI22_X1 u0_u0_U337 (.B1( u0_u0_n441 ) , .ZN( u0_u0_n701 ) , .A2( u0_u0_n735 ) , .A1( u0_u0_n785 ) , .B2( u0_u0_n822 ) );
  AOI21_X1 u0_u0_U338 (.B2( u0_u0_n441 ) , .ZN( u0_u0_n503 ) , .A( u0_u0_n784 ) , .B1( u0_u0_n809 ) );
  AOI21_X1 u0_u0_U339 (.B1( u0_u0_n441 ) , .ZN( u0_u0_n632 ) , .B2( u0_u0_n675 ) , .A( u0_u0_n795 ) );
  NOR4_X1 u0_u0_U34 (.A1( u0_u0_n537 ) , .ZN( u0_u0_n542 ) , .A2( u0_u0_n660 ) , .A4( u0_u0_n674 ) , .A3( u0_u0_n770 ) );
  NAND2_X2 u0_u0_U340 (.A1( u0_u0_n461 ) , .A2( u0_u0_n468 ) , .ZN( u0_u0_n755 ) );
  AOI21_X1 u0_u0_U341 (.B2( u0_u0_n441 ) , .ZN( u0_u0_n570 ) , .B1( u0_u0_n729 ) , .A( u0_u0_n784 ) );
  NAND2_X2 u0_u0_U342 (.A1( u0_u0_n457 ) , .A2( u0_u0_n468 ) , .ZN( u0_u0_n795 ) );
  AOI21_X1 u0_u0_U343 (.B2( u0_u0_n441 ) , .ZN( u0_u0_n449 ) , .B1( u0_u0_n794 ) , .A( u0_u0_n819 ) );
  NOR2_X1 u0_u0_U344 (.A2( u0_u0_n441 ) , .ZN( u0_u0_n670 ) , .A1( u0_u0_n790 ) );
  NOR2_X1 u0_u0_U345 (.A2( u0_u0_n441 ) , .ZN( u0_u0_n561 ) , .A1( u0_u0_n755 ) );
  NOR2_X1 u0_u0_U346 (.A2( u0_u0_n441 ) , .ZN( u0_u0_n565 ) , .A1( u0_u0_n808 ) );
  NOR2_X1 u0_u0_U347 (.A1( u0_u0_n441 ) , .A2( u0_u0_n443 ) , .ZN( u0_u0_n690 ) );
  NOR2_X1 u0_u0_U348 (.A1( u0_u0_n441 ) , .ZN( u0_u0_n648 ) , .A2( u0_u0_n793 ) );
  NAND2_X2 u0_u0_U349 (.A1( u0_u0_n453 ) , .A2( u0_u0_n454 ) , .ZN( u0_u0_n791 ) );
  NOR4_X1 u0_u0_U35 (.A4( u0_u0_n547 ) , .A3( u0_u0_n548 ) , .A2( u0_u0_n549 ) , .ZN( u0_u0_n556 ) , .A1( u0_u0_n694 ) );
  NOR2_X1 u0_u0_U350 (.A2( u0_u0_n441 ) , .ZN( u0_u0_n548 ) , .A1( u0_u0_n767 ) );
  INV_X1 u0_u0_U351 (.A( u0_u0_n796 ) , .ZN( u0_u0_n877 ) );
  NOR2_X1 u0_u0_U352 (.ZN( u0_u0_n586 ) , .A2( u0_u0_n703 ) , .A1( u0_u0_n796 ) );
  NOR2_X1 u0_u0_U353 (.ZN( u0_u0_n467 ) , .A1( u0_u0_n834 ) , .A2( w3_18 ) );
  AOI221_X1 u0_u0_U354 (.A( u0_u0_n582 ) , .ZN( u0_u0_n593 ) , .B2( u0_u0_n836 ) , .C2( u0_u0_n848 ) , .B1( u0_u0_n859 ) , .C1( u0_u0_n865 ) );
  NOR2_X1 u0_u0_U355 (.ZN( u0_u0_n457 ) , .A1( u0_u0_n833 ) , .A2( u0_u0_n834 ) );
  INV_X1 u0_u0_U356 (.ZN( u0_u0_n834 ) , .A( w3_19 ) );
  NAND2_X2 u0_u0_U357 (.A1( u0_u0_n459 ) , .A2( u0_u0_n478 ) , .ZN( u0_u0_n790 ) );
  INV_X1 u0_u0_U358 (.ZN( u0_u0_n833 ) , .A( w3_18 ) );
  AOI222_X1 u0_u0_U359 (.ZN( u0_u0_n611 ) , .B2( u0_u0_n677 ) , .B1( u0_u0_n758 ) , .C2( u0_u0_n836 ) , .A1( u0_u0_n838 ) , .A2( u0_u0_n866 ) , .C1( u0_u0_n867 ) );
  NOR4_X1 u0_u0_U36 (.A4( u0_u0_n583 ) , .A3( u0_u0_n584 ) , .A2( u0_u0_n585 ) , .ZN( u0_u0_n592 ) , .A1( u0_u0_n689 ) );
  AOI222_X1 u0_u0_U360 (.ZN( u0_u0_n519 ) , .C1( u0_u0_n837 ) , .B2( u0_u0_n842 ) , .A2( u0_u0_n848 ) , .C2( u0_u0_n866 ) , .B1( u0_u0_n867 ) , .A1( u0_u0_n870 ) );
  AOI221_X1 u0_u0_U361 (.A( u0_u0_n489 ) , .ZN( u0_u0_n494 ) , .B1( u0_u0_n836 ) , .C2( u0_u0_n849 ) , .C1( u0_u0_n857 ) , .B2( u0_u0_n866 ) );
  NOR2_X1 u0_u0_U362 (.ZN( u0_u0_n794 ) , .A2( u0_u0_n866 ) , .A1( u0_u0_n872 ) );
  INV_X1 u0_u0_U363 (.A( u0_u0_n791 ) , .ZN( u0_u0_n866 ) );
  OAI22_X1 u0_u0_U364 (.ZN( u0_u0_n643 ) , .A1( u0_u0_n705 ) , .B2( u0_u0_n733 ) , .A2( u0_u0_n767 ) , .B1( u0_u0_n821 ) );
  OAI22_X1 u0_u0_U365 (.A1( u0_u0_n729 ) , .ZN( u0_u0_n731 ) , .B2( u0_u0_n755 ) , .B1( u0_u0_n817 ) , .A2( u0_u0_n821 ) );
  AOI21_X1 u0_u0_U366 (.ZN( u0_u0_n505 ) , .B1( u0_u0_n686 ) , .A( u0_u0_n817 ) , .B2( u0_u0_n821 ) );
  AOI21_X1 u0_u0_U367 (.A( u0_u0_n445 ) , .B2( u0_u0_n821 ) , .B1( u0_u0_n822 ) , .ZN( u0_u0_n823 ) );
  OAI22_X1 u0_u0_U368 (.A1( u0_u0_n445 ) , .ZN( u0_u0_n630 ) , .B1( u0_u0_n675 ) , .B2( u0_u0_n752 ) , .A2( u0_u0_n821 ) );
  NOR2_X1 u0_u0_U369 (.A2( u0_u0_n441 ) , .ZN( u0_u0_n605 ) , .A1( u0_u0_n821 ) );
  NOR3_X1 u0_u0_U37 (.ZN( u0_u0_n555 ) , .A2( u0_u0_n657 ) , .A1( u0_u0_n673 ) , .A3( u0_u0_n776 ) );
  NOR2_X1 u0_u0_U370 (.ZN( u0_u0_n537 ) , .A2( u0_u0_n785 ) , .A1( u0_u0_n821 ) );
  NOR2_X1 u0_u0_U371 (.ZN( u0_u0_n525 ) , .A2( u0_u0_n705 ) , .A1( u0_u0_n821 ) );
  NAND2_X2 u0_u0_U372 (.A1( u0_u0_n461 ) , .A2( u0_u0_n477 ) , .ZN( u0_u0_n808 ) );
  NOR2_X1 u0_u0_U373 (.A1( u0_u0_n675 ) , .ZN( u0_u0_n694 ) , .A2( u0_u0_n821 ) );
  NOR2_X1 u0_u0_U374 (.ZN( u0_u0_n564 ) , .A1( u0_u0_n713 ) , .A2( u0_u0_n821 ) );
  NAND2_X2 u0_u0_U375 (.A1( u0_u0_n459 ) , .A2( u0_u0_n467 ) , .ZN( u0_u0_n749 ) );
  NOR2_X1 u0_u0_U376 (.ZN( u0_u0_n691 ) , .A1( u0_u0_n734 ) , .A2( u0_u0_n821 ) );
  INV_X1 u0_u0_U377 (.A( u0_u0_n821 ) , .ZN( u0_u0_n836 ) );
  NAND2_X1 u0_u0_U378 (.ZN( u0_u0_n677 ) , .A1( u0_u0_n811 ) , .A2( u0_u0_n821 ) );
  NOR2_X1 u0_u0_U379 (.ZN( u0_u0_n460 ) , .A1( u0_u0_n832 ) , .A2( w3_16 ) );
  AOI211_X1 u0_u0_U38 (.B( u0_u0_n545 ) , .A( u0_u0_n546 ) , .ZN( u0_u0_n557 ) , .C2( u0_u0_n844 ) , .C1( u0_u0_n856 ) );
  NOR2_X1 u0_u0_U380 (.ZN( u0_u0_n468 ) , .A2( w3_16 ) , .A1( w3_17 ) );
  INV_X1 u0_u0_U381 (.ZN( u0_u0_n831 ) , .A( w3_16 ) );
  AOI211_X1 u0_u0_U382 (.A( u0_u0_n643 ) , .ZN( u0_u0_n651 ) , .B( u0_u0_n748 ) , .C2( u0_u0_n844 ) , .C1( u0_u0_n859 ) );
  NAND4_X1 u0_u0_U383 (.A4( u0_u0_n639 ) , .A3( u0_u0_n640 ) , .A2( u0_u0_n641 ) , .A1( u0_u0_n642 ) , .ZN( u0_u0_n748 ) );
  AOI21_X1 u0_u0_U384 (.ZN( u0_u0_n582 ) , .B2( u0_u0_n729 ) , .B1( u0_u0_n753 ) , .A( u0_u0_n790 ) );
  NAND2_X2 u0_u0_U385 (.A2( u0_u0_n447 ) , .A1( u0_u0_n453 ) , .ZN( u0_u0_n789 ) );
  NOR2_X1 u0_u0_U386 (.ZN( u0_u0_n466 ) , .A1( u0_u0_n854 ) , .A2( w3_23 ) );
  INV_X1 u0_u0_U387 (.ZN( u0_u0_n862 ) , .A( w3_23 ) );
  NOR2_X1 u0_u0_U388 (.ZN( u0_u0_n447 ) , .A2( w3_20 ) , .A1( w3_21 ) );
  NOR2_X1 u0_u0_U389 (.ZN( u0_u0_n454 ) , .A1( u0_u0_n852 ) , .A2( w3_21 ) );
  NOR4_X1 u0_u0_U39 (.A4( u0_u0_n550 ) , .A3( u0_u0_n551 ) , .A2( u0_u0_n552 ) , .A1( u0_u0_n553 ) , .ZN( u0_u0_n554 ) );
  OAI21_X1 u0_u0_U390 (.A( u0_u0_n736 ) , .B1( u0_u0_n737 ) , .ZN( u0_u0_n741 ) , .B2( u0_u0_n810 ) );
  OAI222_X1 u0_u0_U391 (.B2( u0_u0_n752 ) , .B1( u0_u0_n753 ) , .A2( u0_u0_n754 ) , .ZN( u0_u0_n762 ) , .C2( u0_u0_n810 ) , .C1( u0_u0_n819 ) , .A1( u0_u0_n822 ) );
  OAI22_X1 u0_u0_U392 (.B2( u0_u0_n808 ) , .B1( u0_u0_n809 ) , .A2( u0_u0_n810 ) , .A1( u0_u0_n811 ) , .ZN( u0_u0_n813 ) );
  OAI222_X1 u0_u0_U393 (.ZN( u0_u0_n511 ) , .C2( u0_u0_n631 ) , .B2( u0_u0_n653 ) , .B1( u0_u0_n752 ) , .A2( u0_u0_n753 ) , .C1( u0_u0_n810 ) , .A1( u0_u0_n811 ) );
  AOI21_X1 u0_u0_U394 (.ZN( u0_u0_n656 ) , .A( u0_u0_n784 ) , .B1( u0_u0_n797 ) , .B2( u0_u0_n810 ) );
  INV_X1 u0_u0_U395 (.A( u0_u0_n810 ) , .ZN( u0_u0_n864 ) );
  NOR2_X1 u0_u0_U396 (.ZN( u0_u0_n740 ) , .A2( u0_u0_n808 ) , .A1( u0_u0_n810 ) );
  NOR2_X1 u0_u0_U397 (.ZN( u0_u0_n490 ) , .A1( u0_u0_n793 ) , .A2( u0_u0_n810 ) );
  NOR2_X1 u0_u0_U398 (.ZN( u0_u0_n573 ) , .A1( u0_u0_n752 ) , .A2( u0_u0_n810 ) );
  AOI21_X1 u0_u0_U399 (.A( u0_u0_n442 ) , .ZN( u0_u0_n558 ) , .B1( u0_u0_n675 ) , .B2( u0_u0_n810 ) );
  OR4_X1 u0_u0_U4 (.A4( u0_u0_n448 ) , .A2( u0_u0_n449 ) , .A1( u0_u0_n450 ) , .ZN( u0_u0_n451 ) , .A3( u0_u0_n559 ) );
  AOI221_X1 u0_u0_U40 (.A( u0_u0_n495 ) , .ZN( u0_u0_n500 ) , .B2( u0_u0_n841 ) , .C2( u0_u0_n846 ) , .C1( u0_u0_n856 ) , .B1( u0_u0_n864 ) );
  NAND2_X1 u0_u0_U400 (.ZN( u0_u0_n758 ) , .A1( u0_u0_n768 ) , .A2( u0_u0_n810 ) );
  NOR2_X1 u0_u0_U401 (.ZN( u0_u0_n720 ) , .A1( u0_u0_n810 ) , .A2( u0_u0_n822 ) );
  NOR2_X1 u0_u0_U402 (.ZN( u0_u0_n562 ) , .A1( u0_u0_n767 ) , .A2( u0_u0_n810 ) );
  NOR2_X1 u0_u0_U403 (.ZN( u0_u0_n676 ) , .A1( u0_u0_n795 ) , .A2( u0_u0_n810 ) );
  NAND4_X1 u0_u0_U404 (.ZN( u0_subword_27 ) , .A2( u0_u0_n440 ) , .A4( u0_u0_n710 ) , .A3( u0_u0_n711 ) , .A1( u0_u0_n712 ) );
  OAI22_X1 u0_u0_U405 (.B2( u0_u0_n749 ) , .ZN( u0_u0_n751 ) , .A2( u0_u0_n767 ) , .B1( u0_u0_n785 ) , .A1( u0_u0_n797 ) );
  OAI22_X1 u0_u0_U406 (.B1( u0_u0_n441 ) , .ZN( u0_u0_n502 ) , .A2( u0_u0_n749 ) , .A1( u0_u0_n785 ) , .B2( u0_u0_n811 ) );
  NOR2_X1 u0_u0_U407 (.ZN( u0_u0_n522 ) , .A1( u0_u0_n713 ) , .A2( u0_u0_n749 ) );
  OAI22_X1 u0_u0_U408 (.ZN( u0_u0_n715 ) , .A2( u0_u0_n733 ) , .B2( u0_u0_n734 ) , .A1( u0_u0_n749 ) , .B1( u0_u0_n818 ) );
  NOR2_X1 u0_u0_U409 (.A2( u0_u0_n749 ) , .ZN( u0_u0_n774 ) , .A1( u0_u0_n817 ) );
  INV_X1 u0_u0_U41 (.A( u0_u0_n783 ) , .ZN( u0_u0_n871 ) );
  OAI22_X1 u0_u0_U410 (.B1( u0_u0_n446 ) , .ZN( u0_u0_n450 ) , .A2( u0_u0_n733 ) , .A1( u0_u0_n749 ) , .B2( u0_u0_n754 ) );
  NOR2_X1 u0_u0_U411 (.ZN( u0_u0_n553 ) , .A1( u0_u0_n705 ) , .A2( u0_u0_n749 ) );
  NOR2_X1 u0_u0_U412 (.ZN( u0_u0_n536 ) , .A2( u0_u0_n749 ) , .A1( u0_u0_n797 ) );
  NOR2_X1 u0_u0_U413 (.A2( u0_u0_n749 ) , .ZN( u0_u0_n760 ) , .A1( u0_u0_n810 ) );
  NOR2_X1 u0_u0_U414 (.A1( u0_u0_n675 ) , .ZN( u0_u0_n679 ) , .A2( u0_u0_n749 ) );
  NOR2_X1 u0_u0_U415 (.ZN( u0_u0_n723 ) , .A2( u0_u0_n729 ) , .A1( u0_u0_n749 ) );
  NOR2_X1 u0_u0_U416 (.ZN( u0_u0_n588 ) , .A1( u0_u0_n749 ) , .A2( u0_u0_n820 ) );
  INV_X1 u0_u0_U417 (.A( u0_u0_n749 ) , .ZN( u0_u0_n842 ) );
  NAND4_X1 u0_u0_U418 (.ZN( u0_subword_26 ) , .A4( u0_u0_n649 ) , .A3( u0_u0_n650 ) , .A1( u0_u0_n651 ) , .A2( u0_u0_n652 ) );
  OAI22_X1 u0_u0_U419 (.ZN( u0_u0_n594 ) , .A2( u0_u0_n752 ) , .B2( u0_u0_n767 ) , .A1( u0_u0_n768 ) , .B1( u0_u0_n789 ) );
  NOR2_X1 u0_u0_U42 (.ZN( u0_u0_n686 ) , .A2( u0_u0_n839 ) , .A1( u0_u0_n844 ) );
  NAND2_X1 u0_u0_U420 (.A1( u0_u0_n734 ) , .A2( u0_u0_n789 ) , .ZN( u0_u0_n816 ) );
  AOI21_X1 u0_u0_U421 (.ZN( u0_u0_n598 ) , .B1( u0_u0_n733 ) , .B2( u0_u0_n789 ) , .A( u0_u0_n795 ) );
  AOI21_X1 u0_u0_U422 (.ZN( u0_u0_n654 ) , .A( u0_u0_n767 ) , .B2( u0_u0_n789 ) , .B1( u0_u0_n797 ) );
  AOI21_X1 u0_u0_U423 (.ZN( u0_u0_n629 ) , .B1( u0_u0_n705 ) , .A( u0_u0_n784 ) , .B2( u0_u0_n789 ) );
  OAI22_X1 u0_u0_U424 (.ZN( u0_u0_n687 ) , .A1( u0_u0_n705 ) , .A2( u0_u0_n735 ) , .B2( u0_u0_n789 ) , .B1( u0_u0_n822 ) );
  NOR2_X1 u0_u0_U425 (.ZN( u0_u0_n657 ) , .A1( u0_u0_n789 ) , .A2( u0_u0_n793 ) );
  OAI21_X1 u0_u0_U426 (.A( u0_u0_n619 ) , .ZN( u0_u0_n622 ) , .B1( u0_u0_n631 ) , .B2( u0_u0_n789 ) );
  NOR2_X1 u0_u0_U427 (.ZN( u0_u0_n559 ) , .A2( u0_u0_n749 ) , .A1( u0_u0_n789 ) );
  NOR2_X1 u0_u0_U428 (.ZN( u0_u0_n616 ) , .A1( u0_u0_n789 ) , .A2( u0_u0_n821 ) );
  NOR2_X1 u0_u0_U429 (.A2( u0_u0_n442 ) , .ZN( u0_u0_n606 ) , .A1( u0_u0_n789 ) );
  NAND4_X1 u0_u0_U43 (.A4( u0_u0_n609 ) , .A3( u0_u0_n610 ) , .A2( u0_u0_n611 ) , .A1( u0_u0_n612 ) , .ZN( u0_u0_n727 ) );
  INV_X1 u0_u0_U430 (.A( u0_u0_n789 ) , .ZN( u0_u0_n865 ) );
  NOR2_X1 u0_u0_U431 (.ZN( u0_u0_n470 ) , .A2( w3_22 ) , .A1( w3_23 ) );
  NOR2_X1 u0_u0_U432 (.ZN( u0_u0_n458 ) , .A1( u0_u0_n862 ) , .A2( w3_22 ) );
  INV_X1 u0_u0_U433 (.ZN( u0_u0_n854 ) , .A( w3_22 ) );
  AOI21_X1 u0_u0_U434 (.A( u0_u0_n442 ) , .ZN( u0_u0_n506 ) , .B1( u0_u0_n713 ) , .B2( u0_u0_n791 ) );
  OAI22_X1 u0_u0_U435 (.ZN( u0_u0_n596 ) , .B1( u0_u0_n735 ) , .B2( u0_u0_n754 ) , .A2( u0_u0_n791 ) , .A1( u0_u0_n808 ) );
  NOR2_X1 u0_u0_U436 (.ZN( u0_u0_n659 ) , .A1( u0_u0_n767 ) , .A2( u0_u0_n791 ) );
  NAND3_X1 u0_u0_U437 (.ZN( u0_subword_30 ) , .A3( u0_u0_n802 ) , .A2( u0_u0_n803 ) , .A1( u0_u0_n804 ) );
  NAND3_X1 u0_u0_U438 (.ZN( u0_subword_29 ) , .A3( u0_u0_n763 ) , .A2( u0_u0_n764 ) , .A1( u0_u0_n765 ) );
  NAND3_X1 u0_u0_U439 (.ZN( u0_subword_28 ) , .A3( u0_u0_n743 ) , .A2( u0_u0_n744 ) , .A1( u0_u0_n745 ) );
  NOR4_X1 u0_u0_U44 (.A3( u0_u0_n606 ) , .A2( u0_u0_n607 ) , .A1( u0_u0_n608 ) , .ZN( u0_u0_n609 ) , .A4( u0_u0_n661 ) );
  NAND3_X1 u0_u0_U440 (.A3( u0_u0_n681 ) , .A2( u0_u0_n682 ) , .A1( u0_u0_n683 ) , .ZN( u0_u0_n812 ) );
  NAND3_X1 u0_u0_U441 (.ZN( u0_u0_n644 ) , .A3( u0_u0_n713 ) , .A2( u0_u0_n729 ) , .A1( u0_u0_n797 ) );
  NAND3_X1 u0_u0_U442 (.A3( u0_u0_n624 ) , .A2( u0_u0_n625 ) , .A1( u0_u0_n626 ) , .ZN( u0_u0_n730 ) );
  NAND3_X1 u0_u0_U443 (.A1( u0_u0_n591 ) , .A2( u0_u0_n592 ) , .A3( u0_u0_n593 ) , .ZN( u0_u0_n627 ) );
  NAND3_X1 u0_u0_U444 (.ZN( u0_u0_n571 ) , .A3( u0_u0_n686 ) , .A2( u0_u0_n755 ) , .A1( u0_u0_n790 ) );
  NAND3_X1 u0_u0_U445 (.A3( u0_u0_n529 ) , .A2( u0_u0_n530 ) , .A1( u0_u0_n531 ) , .ZN( u0_u0_n747 ) );
  NAND3_X1 u0_u0_U446 (.A3( u0_u0_n518 ) , .A1( u0_u0_n519 ) , .ZN( u0_u0_n614 ) , .A2( u0_u0_n875 ) );
  NAND3_X1 u0_u0_U447 (.A3( u0_u0_n473 ) , .A2( u0_u0_n474 ) , .A1( u0_u0_n475 ) , .ZN( u0_u0_n782 ) );
  NAND2_X1 u0_u0_U448 (.A2( u0_u0_n754 ) , .A1( u0_u0_n791 ) , .ZN( u0_u0_n814 ) );
  NOR2_X1 u0_u0_U449 (.A2( u0_u0_n443 ) , .ZN( u0_u0_n560 ) , .A1( u0_u0_n791 ) );
  NOR3_X1 u0_u0_U45 (.A1( u0_u0_n605 ) , .ZN( u0_u0_n610 ) , .A3( u0_u0_n669 ) , .A2( u0_u0_n775 ) );
  NOR2_X1 u0_u0_U450 (.ZN( u0_u0_n618 ) , .A1( u0_u0_n784 ) , .A2( u0_u0_n791 ) );
  NOR2_X1 u0_u0_U451 (.ZN( u0_u0_n722 ) , .A2( u0_u0_n749 ) , .A1( u0_u0_n791 ) );
  NOR2_X1 u0_u0_U452 (.ZN( u0_u0_n707 ) , .A2( u0_u0_n791 ) , .A1( u0_u0_n822 ) );
  NOR2_X1 u0_u0_U453 (.A1( u0_u0_n735 ) , .ZN( u0_u0_n770 ) , .A2( u0_u0_n791 ) );
  NOR2_X1 u0_u0_U454 (.ZN( u0_u0_n455 ) , .A1( u0_u0_n853 ) , .A2( w3_20 ) );
  INV_X1 u0_u0_U455 (.ZN( u0_u0_n852 ) , .A( w3_20 ) );
  NAND4_X1 u0_u0_U46 (.A4( u0_u0_n566 ) , .A3( u0_u0_n567 ) , .A2( u0_u0_n568 ) , .A1( u0_u0_n569 ) , .ZN( u0_u0_n613 ) );
  NOR4_X1 u0_u0_U47 (.ZN( u0_u0_n567 ) , .A1( u0_u0_n659 ) , .A3( u0_u0_n667 ) , .A4( u0_u0_n691 ) , .A2( u0_u0_n773 ) );
  NOR4_X1 u0_u0_U48 (.A4( u0_u0_n558 ) , .A3( u0_u0_n559 ) , .A2( u0_u0_n560 ) , .A1( u0_u0_n561 ) , .ZN( u0_u0_n568 ) );
  NOR4_X1 u0_u0_U49 (.A4( u0_u0_n562 ) , .A3( u0_u0_n563 ) , .A2( u0_u0_n564 ) , .A1( u0_u0_n565 ) , .ZN( u0_u0_n566 ) );
  OR3_X1 u0_u0_U5 (.ZN( u0_u0_n22 ) , .A3( u0_u0_n658 ) , .A1( u0_u0_n668 ) , .A2( u0_u0_n772 ) );
  NOR4_X1 u0_u0_U50 (.A4( u0_u0_n693 ) , .A3( u0_u0_n694 ) , .A2( u0_u0_n695 ) , .A1( u0_u0_n696 ) , .ZN( u0_u0_n697 ) );
  INV_X1 u0_u0_U51 (.A( u0_u0_n685 ) , .ZN( u0_u0_n876 ) );
  NOR4_X1 u0_u0_U52 (.A4( u0_u0_n532 ) , .A2( u0_u0_n533 ) , .A1( u0_u0_n534 ) , .ZN( u0_u0_n544 ) , .A3( u0_u0_n707 ) );
  NOR4_X1 u0_u0_U53 (.A4( u0_u0_n535 ) , .A3( u0_u0_n536 ) , .ZN( u0_u0_n543 ) , .A2( u0_u0_n690 ) , .A1( u0_u0_n799 ) );
  NOR4_X1 u0_u0_U54 (.A4( u0_u0_n538 ) , .A3( u0_u0_n539 ) , .A2( u0_u0_n540 ) , .ZN( u0_u0_n541 ) , .A1( u0_u0_n825 ) );
  NOR4_X1 u0_u0_U55 (.A4( u0_u0_n520 ) , .A3( u0_u0_n521 ) , .A2( u0_u0_n522 ) , .A1( u0_u0_n523 ) , .ZN( u0_u0_n530 ) );
  NOR4_X1 u0_u0_U56 (.A3( u0_u0_n527 ) , .A1( u0_u0_n528 ) , .ZN( u0_u0_n529 ) , .A2( u0_u0_n679 ) , .A4( u0_u0_n774 ) );
  NOR4_X1 u0_u0_U57 (.A4( u0_u0_n476 ) , .ZN( u0_u0_n482 ) , .A3( u0_u0_n562 ) , .A1( u0_u0_n740 ) , .A2( u0_u0_n760 ) );
  NOR4_X1 u0_u0_U58 (.ZN( u0_u0_n481 ) , .A1( u0_u0_n537 ) , .A3( u0_u0_n574 ) , .A4( u0_u0_n606 ) , .A2( u0_u0_n648 ) );
  NOR4_X1 u0_u0_U59 (.ZN( u0_u0_n480 ) , .A1( u0_u0_n512 ) , .A3( u0_u0_n550 ) , .A2( u0_u0_n589 ) , .A4( u0_u0_n721 ) );
  OR2_X1 u0_u0_U6 (.ZN( u0_u0_n171 ) , .A2( u0_u0_n620 ) , .A1( u0_u0_n621 ) );
  NOR4_X1 u0_u0_U60 (.A4( u0_u0_n635 ) , .A3( u0_u0_n636 ) , .A2( u0_u0_n637 ) , .A1( u0_u0_n638 ) , .ZN( u0_u0_n639 ) );
  NOR4_X1 u0_u0_U61 (.A4( u0_u0_n632 ) , .A3( u0_u0_n633 ) , .A2( u0_u0_n634 ) , .ZN( u0_u0_n640 ) , .A1( u0_u0_n670 ) );
  AOI211_X1 u0_u0_U62 (.B( u0_u0_n629 ) , .A( u0_u0_n630 ) , .ZN( u0_u0_n641 ) , .C2( u0_u0_n841 ) , .C1( u0_u0_n867 ) );
  NAND4_X1 u0_u0_U63 (.A4( u0_u0_n777 ) , .A3( u0_u0_n778 ) , .A2( u0_u0_n779 ) , .A1( u0_u0_n780 ) , .ZN( u0_u0_n806 ) );
  NOR3_X1 u0_u0_U64 (.A3( u0_u0_n770 ) , .A2( u0_u0_n771 ) , .A1( u0_u0_n772 ) , .ZN( u0_u0_n778 ) );
  NOR4_X1 u0_u0_U65 (.A4( u0_u0_n773 ) , .A3( u0_u0_n774 ) , .A2( u0_u0_n775 ) , .A1( u0_u0_n776 ) , .ZN( u0_u0_n777 ) );
  NAND4_X1 u0_u0_U66 (.A4( u0_u0_n663 ) , .A3( u0_u0_n664 ) , .A2( u0_u0_n665 ) , .A1( u0_u0_n666 ) , .ZN( u0_u0_n805 ) );
  NOR3_X1 u0_u0_U67 (.A3( u0_u0_n654 ) , .A2( u0_u0_n655 ) , .A1( u0_u0_n656 ) , .ZN( u0_u0_n665 ) );
  NOR3_X1 u0_u0_U68 (.A3( u0_u0_n657 ) , .A2( u0_u0_n658 ) , .A1( u0_u0_n659 ) , .ZN( u0_u0_n664 ) );
  NOR3_X1 u0_u0_U69 (.A3( u0_u0_n660 ) , .A2( u0_u0_n661 ) , .A1( u0_u0_n662 ) , .ZN( u0_u0_n663 ) );
  OR2_X1 u0_u0_U7 (.ZN( u0_u0_n438 ) , .A1( u0_u0_n782 ) , .A2( u0_u0_n783 ) );
  NOR4_X1 u0_u0_U70 (.A4( u0_u0_n515 ) , .A2( u0_u0_n516 ) , .A1( u0_u0_n517 ) , .ZN( u0_u0_n518 ) , .A3( u0_u0_n676 ) );
  INV_X1 u0_u0_U71 (.A( u0_u0_n511 ) , .ZN( u0_u0_n875 ) );
  NOR2_X1 u0_u0_U72 (.ZN( u0_u0_n809 ) , .A1( u0_u0_n859 ) , .A2( u0_u0_n865 ) );
  NAND4_X1 u0_u0_U73 (.A4( u0_u0_n491 ) , .A3( u0_u0_n492 ) , .A2( u0_u0_n493 ) , .A1( u0_u0_n494 ) , .ZN( u0_u0_n783 ) );
  NOR4_X1 u0_u0_U74 (.A4( u0_u0_n490 ) , .ZN( u0_u0_n493 ) , .A1( u0_u0_n572 ) , .A2( u0_u0_n587 ) , .A3( u0_u0_n608 ) );
  NOR4_X1 u0_u0_U75 (.ZN( u0_u0_n492 ) , .A1( u0_u0_n513 ) , .A2( u0_u0_n525 ) , .A4( u0_u0_n552 ) , .A3( u0_u0_n617 ) );
  NAND4_X1 u0_u0_U76 (.A4( u0_u0_n462 ) , .A3( u0_u0_n463 ) , .A2( u0_u0_n464 ) , .A1( u0_u0_n465 ) , .ZN( u0_u0_n685 ) );
  NOR3_X1 u0_u0_U77 (.ZN( u0_u0_n463 ) , .A3( u0_u0_n536 ) , .A1( u0_u0_n561 ) , .A2( u0_u0_n576 ) );
  AOI221_X1 u0_u0_U78 (.A( u0_u0_n456 ) , .ZN( u0_u0_n465 ) , .C2( u0_u0_n758 ) , .B1( u0_u0_n837 ) , .C1( u0_u0_n847 ) , .B2( u0_u0_n865 ) );
  NOR4_X1 u0_u0_U79 (.ZN( u0_u0_n464 ) , .A2( u0_u0_n515 ) , .A1( u0_u0_n605 ) , .A4( u0_u0_n634 ) , .A3( u0_u0_n716 ) );
  NAND2_X2 u0_u0_U8 (.A2( u0_u0_n477 ) , .A1( u0_u0_n478 ) , .ZN( u0_u0_n822 ) );
  NOR2_X1 u0_u0_U80 (.ZN( u0_u0_n766 ) , .A1( u0_u0_n838 ) , .A2( u0_u0_n839 ) );
  NOR2_X1 u0_u0_U81 (.ZN( u0_u0_n631 ) , .A2( u0_u0_n841 ) , .A1( u0_u0_n844 ) );
  NAND4_X1 u0_u0_U82 (.A4( u0_u0_n485 ) , .A3( u0_u0_n486 ) , .A2( u0_u0_n487 ) , .A1( u0_u0_n488 ) , .ZN( u0_u0_n700 ) );
  NOR3_X1 u0_u0_U83 (.ZN( u0_u0_n486 ) , .A2( u0_u0_n514 ) , .A3( u0_u0_n607 ) , .A1( u0_u0_n616 ) );
  NOR4_X1 u0_u0_U84 (.ZN( u0_u0_n487 ) , .A3( u0_u0_n538 ) , .A4( u0_u0_n551 ) , .A2( u0_u0_n573 ) , .A1( u0_u0_n722 ) );
  AOI211_X1 u0_u0_U85 (.B( u0_u0_n483 ) , .A( u0_u0_n484 ) , .ZN( u0_u0_n488 ) , .C2( u0_u0_n838 ) , .C1( u0_u0_n865 ) );
  AOI222_X1 u0_u0_U86 (.A2( u0_u0_n444 ) , .ZN( u0_u0_n475 ) , .B1( u0_u0_n837 ) , .A1( u0_u0_n844 ) , .C1( u0_u0_n847 ) , .C2( u0_u0_n856 ) , .B2( u0_u0_n869 ) );
  NOR4_X1 u0_u0_U87 (.A1( u0_u0_n472 ) , .ZN( u0_u0_n473 ) , .A4( u0_u0_n548 ) , .A2( u0_u0_n560 ) , .A3( u0_u0_n620 ) );
  AOI221_X1 u0_u0_U88 (.ZN( u0_u0_n474 ) , .C2( u0_u0_n719 ) , .B2( u0_u0_n836 ) , .C1( u0_u0_n850 ) , .B1( u0_u0_n864 ) , .A( u0_u0_n868 ) );
  NAND4_X1 u0_u0_U89 (.A4( u0_u0_n724 ) , .A3( u0_u0_n725 ) , .A2( u0_u0_n726 ) , .ZN( u0_u0_n746 ) , .A1( u0_u0_n861 ) );
  CLKBUF_X1 u0_u0_U9 (.Z( u0_u0_n439 ) , .A( u0_u0_n850 ) );
  INV_X1 u0_u0_U90 (.A( u0_u0_n714 ) , .ZN( u0_u0_n861 ) );
  NOR4_X1 u0_u0_U91 (.A4( u0_u0_n720 ) , .A3( u0_u0_n721 ) , .A2( u0_u0_n722 ) , .A1( u0_u0_n723 ) , .ZN( u0_u0_n724 ) );
  AOI221_X1 u0_u0_U92 (.B2( u0_u0_n439 ) , .A( u0_u0_n715 ) , .ZN( u0_u0_n726 ) , .C2( u0_u0_n849 ) , .C1( u0_u0_n865 ) , .B1( u0_u0_n866 ) );
  NAND4_X1 u0_u0_U93 (.A4( u0_u0_n579 ) , .A3( u0_u0_n580 ) , .A1( u0_u0_n581 ) , .ZN( u0_u0_n728 ) , .A2( u0_u0_n878 ) );
  AOI221_X1 u0_u0_U94 (.A( u0_u0_n570 ) , .C2( u0_u0_n571 ) , .ZN( u0_u0_n580 ) , .B2( u0_u0_n850 ) , .B1( u0_u0_n857 ) , .C1( u0_u0_n858 ) );
  NOR4_X1 u0_u0_U95 (.A4( u0_u0_n575 ) , .A3( u0_u0_n576 ) , .A2( u0_u0_n577 ) , .A1( u0_u0_n578 ) , .ZN( u0_u0_n579 ) );
  INV_X1 u0_u0_U96 (.A( u0_u0_n613 ) , .ZN( u0_u0_n878 ) );
  NOR4_X1 u0_u0_U97 (.A4( u0_u0_n615 ) , .A3( u0_u0_n616 ) , .A2( u0_u0_n617 ) , .A1( u0_u0_n618 ) , .ZN( u0_u0_n625 ) );
  NOR4_X1 u0_u0_U98 (.ZN( u0_u0_n626 ) , .A1( u0_u0_n662 ) , .A3( u0_u0_n672 ) , .A4( u0_u0_n688 ) , .A2( u0_u0_n771 ) );
  NOR2_X1 u0_u0_U99 (.ZN( u0_u0_n692 ) , .A1( u0_u0_n836 ) , .A2( u0_u0_n837 ) );
  DFF_X1 u0_w_reg_0_0 (.CK( clk ) , .D( u0_N42 ) , .Q( w0_0 ) );
  DFF_X1 u0_w_reg_0_1 (.CK( clk ) , .D( u0_N43 ) , .Q( w0_1 ) );
  DFF_X1 u0_w_reg_0_10 (.CK( clk ) , .D( u0_N52 ) , .Q( w0_10 ) );
  DFF_X1 u0_w_reg_0_11 (.CK( clk ) , .D( u0_N53 ) , .Q( w0_11 ) );
  DFF_X1 u0_w_reg_0_12 (.CK( clk ) , .D( u0_N54 ) , .Q( w0_12 ) );
  DFF_X1 u0_w_reg_0_13 (.CK( clk ) , .D( u0_N55 ) , .Q( w0_13 ) );
  DFF_X1 u0_w_reg_0_14 (.CK( clk ) , .D( u0_N56 ) , .Q( w0_14 ) );
  DFF_X1 u0_w_reg_0_15 (.CK( clk ) , .D( u0_N57 ) , .Q( w0_15 ) );
  DFF_X1 u0_w_reg_0_16 (.CK( clk ) , .D( u0_N58 ) , .Q( w0_16 ) );
  DFF_X1 u0_w_reg_0_17 (.CK( clk ) , .D( u0_N59 ) , .Q( w0_17 ) );
  DFF_X1 u0_w_reg_0_18 (.CK( clk ) , .D( u0_N60 ) , .Q( w0_18 ) );
  DFF_X1 u0_w_reg_0_19 (.CK( clk ) , .D( u0_N61 ) , .Q( w0_19 ) );
  DFF_X1 u0_w_reg_0_2 (.CK( clk ) , .D( u0_N44 ) , .Q( w0_2 ) );
  DFF_X1 u0_w_reg_0_20 (.CK( clk ) , .D( u0_N62 ) , .Q( w0_20 ) );
  DFF_X1 u0_w_reg_0_21 (.CK( clk ) , .D( u0_N63 ) , .Q( w0_21 ) );
  DFF_X1 u0_w_reg_0_22 (.CK( clk ) , .D( u0_N64 ) , .Q( w0_22 ) );
  DFF_X1 u0_w_reg_0_23 (.CK( clk ) , .D( u0_N65 ) , .Q( w0_23 ) );
  DFF_X1 u0_w_reg_0_24 (.CK( clk ) , .D( u0_N66 ) , .Q( w0_24 ) );
  DFF_X1 u0_w_reg_0_25 (.CK( clk ) , .D( u0_N67 ) , .Q( w0_25 ) );
  DFF_X1 u0_w_reg_0_26 (.CK( clk ) , .D( u0_N68 ) , .Q( w0_26 ) );
  DFF_X1 u0_w_reg_0_27 (.CK( clk ) , .D( u0_N69 ) , .Q( w0_27 ) );
  DFF_X1 u0_w_reg_0_28 (.CK( clk ) , .D( u0_N70 ) , .Q( w0_28 ) );
  DFF_X1 u0_w_reg_0_29 (.CK( clk ) , .D( u0_N71 ) , .Q( w0_29 ) );
  DFF_X1 u0_w_reg_0_3 (.CK( clk ) , .D( u0_N45 ) , .Q( w0_3 ) );
  DFF_X1 u0_w_reg_0_30 (.CK( clk ) , .D( u0_N72 ) , .Q( w0_30 ) );
  DFF_X1 u0_w_reg_0_31 (.CK( clk ) , .D( u0_N73 ) , .Q( w0_31 ) );
  DFF_X1 u0_w_reg_0_4 (.CK( clk ) , .D( u0_N46 ) , .Q( w0_4 ) );
  DFF_X1 u0_w_reg_0_5 (.CK( clk ) , .D( u0_N47 ) , .Q( w0_5 ) );
  DFF_X1 u0_w_reg_0_6 (.CK( clk ) , .D( u0_N48 ) , .Q( w0_6 ) );
  DFF_X1 u0_w_reg_0_7 (.CK( clk ) , .D( u0_N49 ) , .Q( w0_7 ) );
  DFF_X1 u0_w_reg_0_8 (.CK( clk ) , .D( u0_N50 ) , .Q( w0_8 ) );
  DFF_X1 u0_w_reg_0_9 (.CK( clk ) , .D( u0_N51 ) , .Q( w0_9 ) );
  DFF_X1 u0_w_reg_1_0 (.CK( clk ) , .D( u0_N108 ) , .Q( w1_0 ) );
  DFF_X1 u0_w_reg_1_1 (.CK( clk ) , .D( u0_N109 ) , .Q( w1_1 ) );
  DFF_X1 u0_w_reg_1_10 (.CK( clk ) , .D( u0_N118 ) , .Q( w1_10 ) );
  DFF_X1 u0_w_reg_1_11 (.CK( clk ) , .D( u0_N119 ) , .Q( w1_11 ) );
  DFF_X1 u0_w_reg_1_12 (.CK( clk ) , .D( u0_N120 ) , .Q( w1_12 ) );
  DFF_X1 u0_w_reg_1_13 (.CK( clk ) , .D( u0_N121 ) , .Q( w1_13 ) );
  DFF_X1 u0_w_reg_1_14 (.CK( clk ) , .D( u0_N122 ) , .Q( w1_14 ) );
  DFF_X1 u0_w_reg_1_15 (.CK( clk ) , .D( u0_N123 ) , .Q( w1_15 ) );
  DFF_X1 u0_w_reg_1_16 (.CK( clk ) , .D( u0_N124 ) , .Q( w1_16 ) );
  DFF_X1 u0_w_reg_1_17 (.CK( clk ) , .D( u0_N125 ) , .Q( w1_17 ) );
  DFF_X1 u0_w_reg_1_18 (.CK( clk ) , .D( u0_N126 ) , .Q( w1_18 ) );
  DFF_X1 u0_w_reg_1_19 (.CK( clk ) , .D( u0_N127 ) , .Q( w1_19 ) );
  DFF_X1 u0_w_reg_1_2 (.CK( clk ) , .D( u0_N110 ) , .Q( w1_2 ) );
  DFF_X1 u0_w_reg_1_20 (.CK( clk ) , .D( u0_N128 ) , .Q( w1_20 ) );
  DFF_X1 u0_w_reg_1_21 (.CK( clk ) , .D( u0_N129 ) , .Q( w1_21 ) );
  DFF_X1 u0_w_reg_1_22 (.CK( clk ) , .D( u0_N130 ) , .Q( w1_22 ) );
  DFF_X1 u0_w_reg_1_23 (.CK( clk ) , .D( u0_N131 ) , .Q( w1_23 ) );
  DFF_X1 u0_w_reg_1_24 (.CK( clk ) , .D( u0_N132 ) , .Q( w1_24 ) );
  DFF_X1 u0_w_reg_1_25 (.CK( clk ) , .D( u0_N133 ) , .Q( w1_25 ) );
  DFF_X1 u0_w_reg_1_26 (.CK( clk ) , .D( u0_N134 ) , .QN( u0_n242 ) , .Q( w1_26 ) );
  DFF_X1 u0_w_reg_1_27 (.CK( clk ) , .D( u0_N135 ) , .Q( w1_27 ) );
  DFF_X1 u0_w_reg_1_28 (.CK( clk ) , .D( u0_N136 ) , .Q( w1_28 ) );
  DFF_X1 u0_w_reg_1_29 (.CK( clk ) , .D( u0_N137 ) , .Q( w1_29 ) );
  DFF_X1 u0_w_reg_1_3 (.CK( clk ) , .D( u0_N111 ) , .Q( w1_3 ) );
  DFF_X1 u0_w_reg_1_30 (.CK( clk ) , .D( u0_N138 ) , .QN( u0_n262 ) , .Q( w1_30 ) );
  DFF_X1 u0_w_reg_1_31 (.CK( clk ) , .D( u0_N139 ) , .Q( w1_31 ) );
  DFF_X1 u0_w_reg_1_4 (.CK( clk ) , .D( u0_N112 ) , .Q( w1_4 ) );
  DFF_X1 u0_w_reg_1_5 (.CK( clk ) , .D( u0_N113 ) , .Q( w1_5 ) );
  DFF_X1 u0_w_reg_1_6 (.CK( clk ) , .D( u0_N114 ) , .Q( w1_6 ) );
  DFF_X1 u0_w_reg_1_7 (.CK( clk ) , .D( u0_N115 ) , .Q( w1_7 ) );
  DFF_X1 u0_w_reg_1_8 (.CK( clk ) , .D( u0_N116 ) , .Q( w1_8 ) );
  DFF_X1 u0_w_reg_1_9 (.CK( clk ) , .D( u0_N117 ) , .Q( w1_9 ) );
  DFF_X1 u0_w_reg_2_0 (.CK( clk ) , .D( u0_N174 ) , .Q( w2_0 ) );
  DFF_X1 u0_w_reg_2_1 (.CK( clk ) , .D( u0_N175 ) , .Q( w2_1 ) );
  DFF_X1 u0_w_reg_2_10 (.CK( clk ) , .D( u0_N184 ) , .Q( w2_10 ) );
  DFF_X1 u0_w_reg_2_11 (.CK( clk ) , .D( u0_N185 ) , .Q( w2_11 ) );
  DFF_X1 u0_w_reg_2_12 (.CK( clk ) , .D( u0_N186 ) , .Q( w2_12 ) );
  DFF_X1 u0_w_reg_2_13 (.CK( clk ) , .D( u0_N187 ) , .Q( w2_13 ) );
  DFF_X1 u0_w_reg_2_14 (.CK( clk ) , .D( u0_N188 ) , .Q( w2_14 ) );
  DFF_X1 u0_w_reg_2_15 (.CK( clk ) , .D( u0_N189 ) , .Q( w2_15 ) );
  DFF_X1 u0_w_reg_2_16 (.CK( clk ) , .D( u0_N190 ) , .Q( w2_16 ) );
  DFF_X1 u0_w_reg_2_17 (.CK( clk ) , .D( u0_N191 ) , .Q( w2_17 ) );
  DFF_X1 u0_w_reg_2_18 (.CK( clk ) , .D( u0_N192 ) , .Q( w2_18 ) );
  DFF_X1 u0_w_reg_2_19 (.CK( clk ) , .D( u0_N193 ) , .Q( w2_19 ) );
  DFF_X1 u0_w_reg_2_2 (.CK( clk ) , .D( u0_N176 ) , .Q( w2_2 ) );
  DFF_X1 u0_w_reg_2_20 (.CK( clk ) , .D( u0_N194 ) , .Q( w2_20 ) );
  DFF_X1 u0_w_reg_2_21 (.CK( clk ) , .D( u0_N195 ) , .Q( w2_21 ) );
  DFF_X1 u0_w_reg_2_22 (.CK( clk ) , .D( u0_N196 ) , .Q( w2_22 ) );
  DFF_X1 u0_w_reg_2_23 (.CK( clk ) , .D( u0_N197 ) , .Q( w2_23 ) );
  DFF_X1 u0_w_reg_2_24 (.CK( clk ) , .D( u0_N198 ) , .Q( w2_24 ) );
  DFF_X1 u0_w_reg_2_25 (.CK( clk ) , .D( u0_N199 ) , .Q( w2_25 ) );
  DFF_X1 u0_w_reg_2_26 (.CK( clk ) , .D( u0_N200 ) , .QN( u0_n244 ) , .Q( w2_26 ) );
  DFF_X1 u0_w_reg_2_27 (.CK( clk ) , .D( u0_N201 ) , .Q( w2_27 ) );
  DFF_X1 u0_w_reg_2_28 (.CK( clk ) , .D( u0_N202 ) , .Q( w2_28 ) );
  DFF_X1 u0_w_reg_2_29 (.CK( clk ) , .D( u0_N203 ) , .Q( w2_29 ) );
  DFF_X1 u0_w_reg_2_3 (.CK( clk ) , .D( u0_N177 ) , .Q( w2_3 ) );
  DFF_X1 u0_w_reg_2_30 (.CK( clk ) , .D( u0_N204 ) , .Q( w2_30 ) );
  DFF_X1 u0_w_reg_2_31 (.CK( clk ) , .D( u0_N205 ) , .Q( w2_31 ) );
  DFF_X1 u0_w_reg_2_4 (.CK( clk ) , .D( u0_N178 ) , .Q( w2_4 ) );
  DFF_X1 u0_w_reg_2_5 (.CK( clk ) , .D( u0_N179 ) , .Q( w2_5 ) );
  DFF_X1 u0_w_reg_2_6 (.CK( clk ) , .D( u0_N180 ) , .Q( w2_6 ) );
  DFF_X1 u0_w_reg_2_7 (.CK( clk ) , .D( u0_N181 ) , .Q( w2_7 ) );
  DFF_X1 u0_w_reg_2_8 (.CK( clk ) , .D( u0_N182 ) , .Q( w2_8 ) );
  DFF_X1 u0_w_reg_2_9 (.CK( clk ) , .D( u0_N183 ) , .Q( w2_9 ) );
  DFF_X1 u0_w_reg_3_0 (.CK( clk ) , .D( u0_N240 ) , .Q( w3_0 ) );
  DFF_X1 u0_w_reg_3_1 (.CK( clk ) , .D( u0_N241 ) , .Q( w3_1 ) );
  DFF_X1 u0_w_reg_3_10 (.CK( clk ) , .D( u0_N250 ) , .Q( w3_10 ) );
  DFF_X1 u0_w_reg_3_11 (.CK( clk ) , .D( u0_N251 ) , .Q( w3_11 ) );
  DFF_X1 u0_w_reg_3_12 (.CK( clk ) , .D( u0_N252 ) , .QN( u0_n258 ) , .Q( u0_n274 ) );
  DFF_X1 u0_w_reg_3_13 (.CK( clk ) , .D( u0_N253 ) , .QN( u0_n250 ) , .Q( u0_n272 ) );
  DFF_X1 u0_w_reg_3_14 (.CK( clk ) , .D( u0_N254 ) , .QN( u0_n254 ) , .Q( u0_n270 ) );
  DFF_X1 u0_w_reg_3_15 (.CK( clk ) , .D( u0_N255 ) , .QN( u0_n264 ) , .Q( u0_n268 ) );
  DFF_X1 u0_w_reg_3_16 (.CK( clk ) , .D( u0_N256 ) , .Q( w3_16 ) );
  DFF_X1 u0_w_reg_3_17 (.CK( clk ) , .D( u0_N257 ) , .Q( w3_17 ) );
  DFF_X1 u0_w_reg_3_18 (.CK( clk ) , .D( u0_N258 ) , .Q( w3_18 ) );
  DFF_X1 u0_w_reg_3_19 (.CK( clk ) , .D( u0_N259 ) , .Q( w3_19 ) );
  DFF_X1 u0_w_reg_3_2 (.CK( clk ) , .D( u0_N242 ) , .Q( w3_2 ) );
  DFF_X1 u0_w_reg_3_20 (.CK( clk ) , .D( u0_N260 ) , .Q( w3_20 ) );
  DFF_X1 u0_w_reg_3_21 (.CK( clk ) , .D( u0_N261 ) , .Q( w3_21 ) );
  DFF_X1 u0_w_reg_3_22 (.CK( clk ) , .D( u0_N262 ) , .Q( w3_22 ) );
  DFF_X1 u0_w_reg_3_23 (.CK( clk ) , .D( u0_N263 ) , .Q( w3_23 ) );
  DFF_X1 u0_w_reg_3_24 (.CK( clk ) , .D( u0_N264 ) , .QN( u0_n248 ) , .Q( w3_24 ) );
  DFF_X1 u0_w_reg_3_25 (.CK( clk ) , .D( u0_N265 ) , .Q( w3_25 ) );
  DFF_X1 u0_w_reg_3_26 (.CK( clk ) , .D( u0_N266 ) , .Q( w3_26 ) );
  DFF_X1 u0_w_reg_3_27 (.CK( clk ) , .D( u0_N267 ) , .Q( w3_27 ) );
  DFF_X1 u0_w_reg_3_28 (.CK( clk ) , .D( u0_N268 ) , .Q( w3_28 ) );
  DFF_X1 u0_w_reg_3_29 (.CK( clk ) , .D( u0_N269 ) , .Q( w3_29 ) );
  DFF_X1 u0_w_reg_3_3 (.CK( clk ) , .D( u0_N243 ) , .Q( w3_3 ) );
  DFF_X1 u0_w_reg_3_30 (.CK( clk ) , .D( u0_N270 ) , .Q( w3_30 ) );
  DFF_X1 u0_w_reg_3_31 (.CK( clk ) , .D( u0_N271 ) , .Q( w3_31 ) );
  DFF_X1 u0_w_reg_3_4 (.CK( clk ) , .D( u0_N244 ) , .Q( w3_4 ) );
  DFF_X1 u0_w_reg_3_5 (.CK( clk ) , .D( u0_N245 ) , .Q( w3_5 ) );
  DFF_X1 u0_w_reg_3_6 (.CK( clk ) , .D( u0_N246 ) , .Q( w3_6 ) );
  DFF_X1 u0_w_reg_3_7 (.CK( clk ) , .D( u0_N247 ) , .Q( w3_7 ) );
  DFF_X1 u0_w_reg_3_8 (.CK( clk ) , .D( u0_N248 ) , .Q( w3_8 ) );
  DFF_X1 u0_w_reg_3_9 (.CK( clk ) , .D( u0_N249 ) , .Q( w3_9 ) );
  NOR2_X1 us22_U10 (.ZN( us22_n573 ) , .A1( us22_n620 ) , .A2( us22_n743 ) );
  NOR4_X1 us22_U100 (.A4( us22_n527 ) , .A3( us22_n528 ) , .ZN( us22_n535 ) , .A2( us22_n682 ) , .A1( us22_n792 ) );
  NAND4_X1 us22_U101 (.A4( us22_n477 ) , .A3( us22_n478 ) , .A2( us22_n479 ) , .A1( us22_n480 ) , .ZN( us22_n692 ) );
  NOR3_X1 us22_U102 (.ZN( us22_n478 ) , .A2( us22_n506 ) , .A3( us22_n599 ) , .A1( us22_n608 ) );
  AOI211_X1 us22_U103 (.B( us22_n475 ) , .A( us22_n476 ) , .ZN( us22_n480 ) , .C2( us22_n831 ) , .C1( us22_n859 ) );
  NOR4_X1 us22_U104 (.ZN( us22_n479 ) , .A3( us22_n530 ) , .A4( us22_n543 ) , .A2( us22_n565 ) , .A1( us22_n715 ) );
  NAND4_X1 us22_U105 (.A4( us22_n546 ) , .A3( us22_n547 ) , .A2( us22_n548 ) , .A1( us22_n549 ) , .ZN( us22_n743 ) );
  NOR3_X1 us22_U106 (.ZN( us22_n547 ) , .A2( us22_n649 ) , .A1( us22_n665 ) , .A3( us22_n769 ) );
  AOI211_X1 us22_U107 (.B( us22_n537 ) , .A( us22_n538 ) , .ZN( us22_n549 ) , .C2( us22_n837 ) , .C1( us22_n849 ) );
  NOR4_X1 us22_U108 (.A4( us22_n542 ) , .A3( us22_n543 ) , .A2( us22_n544 ) , .A1( us22_n545 ) , .ZN( us22_n546 ) );
  NOR2_X1 us22_U109 (.ZN( us22_n684 ) , .A1( us22_n829 ) , .A2( us22_n830 ) );
  NOR2_X1 us22_U11 (.A1( us22_n676 ) , .ZN( us22_n691 ) , .A2( us22_n805 ) );
  NOR4_X1 us22_U110 (.ZN( us22_n618 ) , .A1( us22_n654 ) , .A3( us22_n664 ) , .A4( us22_n680 ) , .A2( us22_n764 ) );
  NOR4_X1 us22_U111 (.A4( us22_n607 ) , .A3( us22_n608 ) , .A2( us22_n609 ) , .A1( us22_n610 ) , .ZN( us22_n617 ) );
  NOR4_X1 us22_U112 (.A4( us22_n612 ) , .A3( us22_n613 ) , .A2( us22_n614 ) , .A1( us22_n615 ) , .ZN( us22_n616 ) );
  NAND4_X1 us22_U113 (.A4( us22_n483 ) , .A3( us22_n484 ) , .A2( us22_n485 ) , .A1( us22_n486 ) , .ZN( us22_n776 ) );
  NOR4_X1 us22_U114 (.A4( us22_n482 ) , .ZN( us22_n485 ) , .A1( us22_n564 ) , .A2( us22_n579 ) , .A3( us22_n600 ) );
  NOR4_X1 us22_U115 (.ZN( us22_n484 ) , .A1( us22_n505 ) , .A2( us22_n517 ) , .A4( us22_n544 ) , .A3( us22_n609 ) );
  NOR4_X1 us22_U116 (.ZN( us22_n483 ) , .A2( us22_n531 ) , .A1( us22_n556 ) , .A3( us22_n629 ) , .A4( us22_n716 ) );
  NAND4_X1 us22_U117 (.A4( us22_n689 ) , .A3( us22_n690 ) , .A1( us22_n691 ) , .ZN( us22_n774 ) , .A2( us22_n870 ) );
  AOI221_X1 us22_U118 (.A( us22_n679 ) , .ZN( us22_n690 ) , .B2( us22_n838 ) , .C1( us22_n840 ) , .C2( us22_n860 ) , .B1( us22_n863 ) );
  INV_X1 us22_U119 (.A( us22_n677 ) , .ZN( us22_n870 ) );
  INV_X1 us22_U12 (.A( us22_n678 ) , .ZN( us22_n838 ) );
  NOR4_X1 us22_U120 (.A4( us22_n685 ) , .A3( us22_n686 ) , .A2( us22_n687 ) , .A1( us22_n688 ) , .ZN( us22_n689 ) );
  NAND4_X1 us22_U121 (.A4( us22_n717 ) , .A3( us22_n718 ) , .A2( us22_n719 ) , .ZN( us22_n739 ) , .A1( us22_n855 ) );
  INV_X1 us22_U122 (.A( us22_n707 ) , .ZN( us22_n855 ) );
  AOI221_X1 us22_U123 (.A( us22_n708 ) , .ZN( us22_n719 ) , .C2( us22_n842 ) , .B2( us22_n843 ) , .C1( us22_n859 ) , .B1( us22_n860 ) );
  NOR4_X1 us22_U124 (.A4( us22_n713 ) , .A3( us22_n714 ) , .A2( us22_n715 ) , .A1( us22_n716 ) , .ZN( us22_n717 ) );
  NAND4_X1 us22_U125 (.A4( us22_n471 ) , .A3( us22_n472 ) , .A2( us22_n473 ) , .A1( us22_n474 ) , .ZN( us22_n676 ) );
  NOR4_X1 us22_U126 (.A4( us22_n468 ) , .ZN( us22_n474 ) , .A3( us22_n554 ) , .A1( us22_n733 ) , .A2( us22_n753 ) );
  NOR4_X1 us22_U127 (.ZN( us22_n473 ) , .A1( us22_n529 ) , .A3( us22_n566 ) , .A4( us22_n598 ) , .A2( us22_n640 ) );
  NOR4_X1 us22_U128 (.ZN( us22_n472 ) , .A1( us22_n504 ) , .A3( us22_n542 ) , .A2( us22_n581 ) , .A4( us22_n714 ) );
  NOR2_X1 us22_U129 (.ZN( us22_n731 ) , .A2( us22_n830 ) , .A1( us22_n843 ) );
  NOR4_X1 us22_U13 (.A4( us22_n443 ) , .A3( us22_n444 ) , .A2( us22_n514 ) , .A1( us22_n539 ) , .ZN( us22_n704 ) );
  NOR2_X1 us22_U130 (.ZN( us22_n787 ) , .A2( us22_n860 ) , .A1( us22_n866 ) );
  NOR2_X1 us22_U131 (.ZN( us22_n645 ) , .A1( us22_n852 ) , .A2( us22_n866 ) );
  NAND4_X1 us22_U132 (.A4( us22_n571 ) , .A3( us22_n572 ) , .A1( us22_n573 ) , .ZN( us22_n721 ) , .A2( us22_n872 ) );
  NOR4_X1 us22_U133 (.A4( us22_n567 ) , .A3( us22_n568 ) , .A2( us22_n569 ) , .A1( us22_n570 ) , .ZN( us22_n571 ) );
  AOI221_X1 us22_U134 (.A( us22_n562 ) , .C2( us22_n563 ) , .ZN( us22_n572 ) , .B2( us22_n843 ) , .B1( us22_n850 ) , .C1( us22_n851 ) );
  INV_X1 us22_U135 (.A( us22_n605 ) , .ZN( us22_n872 ) );
  NAND4_X1 us22_U136 (.A4( us22_n491 ) , .A3( us22_n492 ) , .A1( us22_n493 ) , .ZN( us22_n800 ) , .A2( us22_n865 ) );
  AOI221_X1 us22_U137 (.A( us22_n487 ) , .ZN( us22_n492 ) , .B2( us22_n834 ) , .C2( us22_n839 ) , .C1( us22_n849 ) , .B1( us22_n858 ) );
  INV_X1 us22_U138 (.A( us22_n776 ) , .ZN( us22_n865 ) );
  NOR2_X1 us22_U139 (.ZN( us22_n493 ) , .A1( us22_n676 ) , .A2( us22_n692 ) );
  OR3_X1 us22_U14 (.ZN( us22_n444 ) , .A1( us22_n526 ) , .A3( us22_n575 ) , .A2( us22_n873 ) );
  INV_X1 us22_U140 (.A( us22_n760 ) , .ZN( us22_n828 ) );
  INV_X1 us22_U141 (.A( us22_n461 ) , .ZN( us22_n862 ) );
  OAI21_X1 us22_U142 (.ZN( us22_n461 ) , .B1( us22_n807 ) , .A( us22_n832 ) , .B2( us22_n849 ) );
  OR4_X1 us22_U143 (.A4( us22_n578 ) , .A3( us22_n579 ) , .A2( us22_n580 ) , .A1( us22_n581 ) , .ZN( us22_n582 ) );
  OR4_X1 us22_U144 (.A4( us22_n680 ) , .A3( us22_n681 ) , .A2( us22_n682 ) , .A1( us22_n683 ) , .ZN( us22_n688 ) );
  OR4_X1 us22_U145 (.A4( us22_n564 ) , .A3( us22_n565 ) , .A2( us22_n566 ) , .ZN( us22_n570 ) , .A1( us22_n663 ) );
  OR4_X1 us22_U146 (.A4( us22_n516 ) , .A2( us22_n517 ) , .A1( us22_n518 ) , .ZN( us22_n520 ) , .A3( us22_n819 ) );
  OR4_X1 us22_U147 (.ZN( us22_n464 ) , .A4( us22_n516 ) , .A3( us22_n527 ) , .A2( us22_n576 ) , .A1( us22_n710 ) );
  NAND2_X1 us22_U148 (.ZN( us22_n611 ) , .A2( us22_n835 ) , .A1( us22_n871 ) );
  OR3_X1 us22_U149 (.A3( us22_n504 ) , .A2( us22_n505 ) , .A1( us22_n506 ) , .ZN( us22_n509 ) );
  OR4_X1 us22_U15 (.A4( us22_n440 ) , .A2( us22_n441 ) , .A1( us22_n442 ) , .ZN( us22_n443 ) , .A3( us22_n551 ) );
  AOI221_X1 us22_U150 (.A( us22_n711 ) , .B2( us22_n712 ) , .ZN( us22_n718 ) , .C1( us22_n830 ) , .B1( us22_n837 ) , .C2( us22_n861 ) );
  OR2_X1 us22_U151 (.A2( us22_n709 ) , .A1( us22_n710 ) , .ZN( us22_n711 ) );
  INV_X1 us22_U152 (.A( us22_n752 ) , .ZN( us22_n867 ) );
  OAI21_X1 us22_U153 (.B1( us22_n751 ) , .ZN( us22_n752 ) , .A( us22_n843 ) , .B2( us22_n866 ) );
  INV_X1 us22_U154 (.A( us22_n670 ) , .ZN( us22_n857 ) );
  AOI21_X1 us22_U155 (.A( us22_n668 ) , .B1( us22_n669 ) , .ZN( us22_n670 ) , .B2( us22_n854 ) );
  NAND2_X1 us22_U156 (.A1( us22_n445 ) , .A2( us22_n463 ) , .ZN( us22_n747 ) );
  OAI222_X1 us22_U157 (.B2( us22_n745 ) , .B1( us22_n746 ) , .A2( us22_n747 ) , .ZN( us22_n755 ) , .C2( us22_n803 ) , .C1( us22_n812 ) , .A1( us22_n815 ) );
  OAI222_X1 us22_U158 (.B2( us22_n706 ) , .ZN( us22_n707 ) , .C2( us22_n722 ) , .B1( us22_n745 ) , .A1( us22_n804 ) , .C1( us22_n812 ) , .A2( us22_n813 ) );
  OAI222_X1 us22_U159 (.ZN( us22_n615 ) , .B1( us22_n695 ) , .C1( us22_n722 ) , .C2( us22_n745 ) , .B2( us22_n784 ) , .A2( us22_n790 ) , .A1( us22_n814 ) );
  INV_X1 us22_U16 (.A( us22_n611 ) , .ZN( us22_n873 ) );
  OAI222_X1 us22_U160 (.ZN( us22_n503 ) , .C2( us22_n623 ) , .B2( us22_n645 ) , .B1( us22_n745 ) , .A2( us22_n746 ) , .C1( us22_n803 ) , .A1( us22_n804 ) );
  NOR4_X1 us22_U161 (.A2( us22_n489 ) , .A1( us22_n490 ) , .ZN( us22_n491 ) , .A3( us22_n578 ) , .A4( us22_n610 ) );
  OR4_X1 us22_U162 (.ZN( us22_n490 ) , .A4( us22_n532 ) , .A2( us22_n545 ) , .A1( us22_n557 ) , .A3( us22_n630 ) );
  OAI22_X1 us22_U163 (.B1( us22_n488 ) , .ZN( us22_n489 ) , .A1( us22_n684 ) , .A2( us22_n761 ) , .B2( us22_n815 ) );
  NOR3_X1 us22_U164 (.ZN( us22_n488 ) , .A1( us22_n780 ) , .A2( us22_n848 ) , .A3( us22_n861 ) );
  AOI22_X1 us22_U165 (.ZN( us22_n694 ) , .A1( us22_n828 ) , .B2( us22_n841 ) , .A2( us22_n863 ) , .B1( us22_n866 ) );
  AOI22_X1 us22_U166 (.A2( us22_n780 ) , .ZN( us22_n781 ) , .B2( us22_n829 ) , .A1( us22_n832 ) , .B1( us22_n861 ) );
  INV_X1 us22_U167 (.A( us22_n728 ) , .ZN( us22_n837 ) );
  AOI221_X1 us22_U168 (.A( us22_n481 ) , .ZN( us22_n486 ) , .B1( us22_n829 ) , .C2( us22_n842 ) , .C1( us22_n850 ) , .B2( us22_n860 ) );
  OAI22_X1 us22_U169 (.ZN( us22_n481 ) , .A1( us22_n706 ) , .B2( us22_n783 ) , .A2( us22_n804 ) , .B1( us22_n810 ) );
  INV_X1 us22_U17 (.A( us22_n747 ) , .ZN( us22_n861 ) );
  INV_X1 us22_U170 (.A( us22_n788 ) , .ZN( us22_n830 ) );
  NAND2_X1 us22_U171 (.A1( us22_n449 ) , .A2( us22_n451 ) , .ZN( us22_n760 ) );
  OAI22_X1 us22_U172 (.ZN( us22_n635 ) , .A1( us22_n697 ) , .B2( us22_n726 ) , .A2( us22_n760 ) , .B1( us22_n814 ) );
  OAI221_X1 us22_U173 (.A( us22_n725 ) , .C2( us22_n726 ) , .B2( us22_n727 ) , .B1( us22_n728 ) , .ZN( us22_n735 ) , .C1( us22_n815 ) );
  AOI22_X1 us22_U174 (.ZN( us22_n725 ) , .B1( us22_n830 ) , .A2( us22_n836 ) , .A1( us22_n861 ) , .B2( us22_n864 ) );
  OAI22_X1 us22_U175 (.ZN( us22_n708 ) , .A2( us22_n726 ) , .B2( us22_n727 ) , .A1( us22_n742 ) , .B1( us22_n811 ) );
  INV_X1 us22_U176 (.A( us22_n814 ) , .ZN( us22_n829 ) );
  OAI22_X1 us22_U177 (.ZN( us22_n487 ) , .A1( us22_n722 ) , .B2( us22_n726 ) , .B1( us22_n728 ) , .A2( us22_n777 ) );
  OAI22_X1 us22_U178 (.ZN( us22_n622 ) , .B1( us22_n667 ) , .B2( us22_n745 ) , .A1( us22_n813 ) , .A2( us22_n814 ) );
  INV_X1 us22_U179 (.A( us22_n742 ) , .ZN( us22_n835 ) );
  AOI222_X1 us22_U18 (.ZN( us22_n603 ) , .B2( us22_n669 ) , .B1( us22_n751 ) , .C2( us22_n829 ) , .A1( us22_n831 ) , .A2( us22_n860 ) , .C1( us22_n861 ) );
  OAI22_X1 us22_U180 (.A1( us22_n722 ) , .ZN( us22_n724 ) , .B2( us22_n748 ) , .B1( us22_n810 ) , .A2( us22_n814 ) );
  OAI22_X1 us22_U181 (.B2( us22_n777 ) , .B1( us22_n778 ) , .ZN( us22_n779 ) , .A2( us22_n812 ) , .A1( us22_n813 ) );
  INV_X1 us22_U182 (.A( us22_n786 ) , .ZN( us22_n843 ) );
  INV_X1 us22_U183 (.A( us22_n812 ) , .ZN( us22_n831 ) );
  OAI22_X1 us22_U184 (.B2( us22_n742 ) , .ZN( us22_n744 ) , .A2( us22_n760 ) , .B1( us22_n778 ) , .A1( us22_n790 ) );
  OAI22_X1 us22_U185 (.B2( us22_n801 ) , .B1( us22_n802 ) , .A2( us22_n803 ) , .A1( us22_n804 ) , .ZN( us22_n806 ) );
  INV_X1 us22_U186 (.A( us22_n667 ) , .ZN( us22_n863 ) );
  OAI22_X1 us22_U187 (.ZN( us22_n494 ) , .A2( us22_n742 ) , .A1( us22_n778 ) , .B1( us22_n789 ) , .B2( us22_n804 ) );
  INV_X1 us22_U188 (.A( us22_n748 ) , .ZN( us22_n840 ) );
  OAI22_X1 us22_U189 (.ZN( us22_n588 ) , .B1( us22_n728 ) , .B2( us22_n747 ) , .A2( us22_n784 ) , .A1( us22_n801 ) );
  AOI222_X1 us22_U19 (.ZN( us22_n561 ) , .B1( us22_n828 ) , .C1( us22_n839 ) , .A2( us22_n841 ) , .A1( us22_n852 ) , .B2( us22_n861 ) , .C2( us22_n871 ) );
  OAI22_X1 us22_U190 (.ZN( us22_n693 ) , .A2( us22_n728 ) , .A1( us22_n778 ) , .B1( us22_n789 ) , .B2( us22_n815 ) );
  INV_X1 us22_U191 (.A( us22_n801 ) , .ZN( us22_n841 ) );
  NOR2_X1 us22_U192 (.A1( us22_n695 ) , .ZN( us22_n768 ) , .A2( us22_n813 ) );
  NOR2_X1 us22_U193 (.ZN( us22_n664 ) , .A1( us22_n726 ) , .A2( us22_n801 ) );
  NOR2_X1 us22_U194 (.ZN( us22_n592 ) , .A2( us22_n695 ) , .A1( us22_n726 ) );
  NOR2_X1 us22_U195 (.ZN( us22_n568 ) , .A1( us22_n726 ) , .A2( us22_n804 ) );
  NOR2_X1 us22_U196 (.ZN( us22_n716 ) , .A2( us22_n722 ) , .A1( us22_n742 ) );
  NOR2_X1 us22_U197 (.ZN( us22_n544 ) , .A2( us22_n778 ) , .A1( us22_n812 ) );
  NOR2_X1 us22_U198 (.ZN( us22_n575 ) , .A2( us22_n697 ) , .A1( us22_n812 ) );
  NOR2_X1 us22_U199 (.ZN( us22_n652 ) , .A1( us22_n726 ) , .A2( us22_n811 ) );
  AOI222_X1 us22_U20 (.ZN( us22_n658 ) , .A2( us22_n837 ) , .B1( us22_n839 ) , .C2( us22_n843 ) , .A1( us22_n858 ) , .C1( us22_n861 ) , .B2( us22_n868 ) );
  NOR2_X1 us22_U200 (.ZN( us22_n610 ) , .A1( us22_n777 ) , .A2( us22_n784 ) );
  NOR2_X1 us22_U201 (.ZN( us22_n530 ) , .A2( us22_n747 ) , .A1( us22_n748 ) );
  NOR2_X1 us22_U202 (.ZN( us22_n627 ) , .A2( us22_n726 ) , .A1( us22_n783 ) );
  NOR2_X1 us22_U203 (.ZN( us22_n613 ) , .A1( us22_n783 ) , .A2( us22_n813 ) );
  NOR2_X1 us22_U204 (.ZN( us22_n599 ) , .A2( us22_n778 ) , .A1( us22_n801 ) );
  NOR2_X1 us22_U205 (.ZN( us22_n609 ) , .A2( us22_n778 ) , .A1( us22_n804 ) );
  INV_X1 us22_U206 (.A( us22_n745 ) , .ZN( us22_n832 ) );
  NOR2_X1 us22_U207 (.A2( us22_n742 ) , .ZN( us22_n767 ) , .A1( us22_n810 ) );
  NOR2_X1 us22_U208 (.ZN( us22_n526 ) , .A2( us22_n722 ) , .A1( us22_n801 ) );
  NOR2_X1 us22_U209 (.ZN( us22_n529 ) , .A2( us22_n778 ) , .A1( us22_n814 ) );
  INV_X1 us22_U21 (.A( us22_n645 ) , .ZN( us22_n868 ) );
  NOR2_X1 us22_U210 (.ZN( us22_n626 ) , .A2( us22_n667 ) , .A1( us22_n783 ) );
  NOR2_X1 us22_U211 (.ZN( us22_n597 ) , .A2( us22_n789 ) , .A1( us22_n814 ) );
  INV_X1 us22_U212 (.A( us22_n790 ) , .ZN( us22_n849 ) );
  INV_X1 us22_U213 (.A( us22_n726 ) , .ZN( us22_n850 ) );
  NOR2_X1 us22_U214 (.ZN( us22_n650 ) , .A1( us22_n667 ) , .A2( us22_n812 ) );
  NOR2_X1 us22_U215 (.A1( us22_n667 ) , .ZN( us22_n671 ) , .A2( us22_n742 ) );
  INV_X1 us22_U216 (.A( us22_n803 ) , .ZN( us22_n858 ) );
  NOR2_X1 us22_U217 (.ZN( us22_n600 ) , .A1( us22_n667 ) , .A2( us22_n801 ) );
  NOR2_X1 us22_U218 (.A1( us22_n667 ) , .ZN( us22_n686 ) , .A2( us22_n814 ) );
  NOR2_X1 us22_U219 (.A2( us22_n706 ) , .A1( us22_n748 ) , .ZN( us22_n769 ) );
  NOR4_X1 us22_U22 (.ZN( us22_n471 ) , .A2( us22_n519 ) , .A4( us22_n592 ) , .A1( us22_n607 ) , .A3( us22_n627 ) );
  NOR2_X1 us22_U220 (.A1( us22_n667 ) , .ZN( us22_n764 ) , .A2( us22_n811 ) );
  NOR2_X1 us22_U221 (.A1( us22_n697 ) , .ZN( us22_n766 ) , .A2( us22_n811 ) );
  NOR2_X1 us22_U222 (.ZN( us22_n539 ) , .A2( us22_n695 ) , .A1( us22_n697 ) );
  NOR2_X1 us22_U223 (.ZN( us22_n525 ) , .A1( us22_n667 ) , .A2( us22_n777 ) );
  NOR2_X1 us22_U224 (.ZN( us22_n665 ) , .A1( us22_n748 ) , .A2( us22_n813 ) );
  NOR2_X1 us22_U225 (.ZN( us22_n553 ) , .A1( us22_n748 ) , .A2( us22_n789 ) );
  NOR2_X1 us22_U226 (.ZN( us22_n506 ) , .A2( us22_n778 ) , .A1( us22_n783 ) );
  NOR2_X1 us22_U227 (.ZN( us22_n541 ) , .A2( us22_n706 ) , .A1( us22_n783 ) );
  NOR2_X1 us22_U228 (.ZN( us22_n662 ) , .A1( us22_n783 ) , .A2( us22_n789 ) );
  NOR2_X1 us22_U229 (.A2( us22_n695 ) , .ZN( us22_n714 ) , .A1( us22_n790 ) );
  NOR4_X1 us22_U23 (.ZN( us22_n477 ) , .A1( us22_n518 ) , .A4( us22_n555 ) , .A3( us22_n580 ) , .A2( us22_n628 ) );
  NOR2_X1 us22_U230 (.ZN( us22_n505 ) , .A1( us22_n810 ) , .A2( us22_n815 ) );
  INV_X1 us22_U231 (.A( us22_n804 ) , .ZN( us22_n839 ) );
  NOR2_X1 us22_U232 (.ZN( us22_n659 ) , .A1( us22_n727 ) , .A2( us22_n788 ) );
  NOR2_X1 us22_U233 (.ZN( us22_n660 ) , .A2( us22_n695 ) , .A1( us22_n727 ) );
  NOR2_X1 us22_U234 (.ZN( us22_n555 ) , .A1( us22_n790 ) , .A2( us22_n812 ) );
  NOR2_X1 us22_U235 (.ZN( us22_n543 ) , .A1( us22_n747 ) , .A2( us22_n812 ) );
  NOR2_X1 us22_U236 (.ZN( us22_n507 ) , .A1( us22_n727 ) , .A2( us22_n777 ) );
  NOR2_X1 us22_U237 (.A2( us22_n695 ) , .A1( us22_n778 ) , .ZN( us22_n818 ) );
  OAI22_X1 us22_U238 (.B2( us22_n748 ) , .B1( us22_n749 ) , .A1( us22_n750 ) , .ZN( us22_n754 ) , .A2( us22_n804 ) );
  NOR2_X1 us22_U239 (.ZN( us22_n749 ) , .A2( us22_n850 ) , .A1( us22_n858 ) );
  NOR4_X1 us22_U24 (.ZN( us22_n454 ) , .A2( us22_n515 ) , .A1( us22_n541 ) , .A3( us22_n577 ) , .A4( us22_n613 ) );
  NOR3_X1 us22_U240 (.ZN( us22_n750 ) , .A2( us22_n851 ) , .A1( us22_n861 ) , .A3( us22_n863 ) );
  NOR2_X1 us22_U241 (.ZN( us22_n528 ) , .A2( us22_n742 ) , .A1( us22_n790 ) );
  NOR2_X1 us22_U242 (.A1( us22_n747 ) , .ZN( us22_n765 ) , .A2( us22_n801 ) );
  NOR2_X1 us22_U243 (.A2( us22_n742 ) , .ZN( us22_n753 ) , .A1( us22_n803 ) );
  NOR2_X1 us22_U244 (.ZN( us22_n542 ) , .A2( us22_n783 ) , .A1( us22_n790 ) );
  NOR2_X1 us22_U245 (.ZN( us22_n661 ) , .A1( us22_n727 ) , .A2( us22_n783 ) );
  NOR2_X1 us22_U246 (.ZN( us22_n629 ) , .A1( us22_n722 ) , .A2( us22_n811 ) );
  NOR2_X1 us22_U247 (.ZN( us22_n733 ) , .A2( us22_n801 ) , .A1( us22_n803 ) );
  NOR2_X1 us22_U248 (.ZN( us22_n612 ) , .A1( us22_n760 ) , .A2( us22_n810 ) );
  OAI22_X1 us22_U249 (.B1( us22_n438 ) , .ZN( us22_n442 ) , .A2( us22_n726 ) , .A1( us22_n742 ) , .B2( us22_n747 ) );
  NOR4_X1 us22_U25 (.A4( us22_n530 ) , .A3( us22_n531 ) , .A2( us22_n532 ) , .ZN( us22_n533 ) , .A1( us22_n818 ) );
  NOR3_X1 us22_U250 (.ZN( us22_n438 ) , .A2( us22_n834 ) , .A3( us22_n835 ) , .A1( us22_n844 ) );
  NOR2_X1 us22_U251 (.ZN( us22_n504 ) , .A2( us22_n726 ) , .A1( us22_n760 ) );
  NOR2_X1 us22_U252 (.ZN( us22_n514 ) , .A1( us22_n706 ) , .A2( us22_n742 ) );
  NOR2_X1 us22_U253 (.ZN( us22_n715 ) , .A2( us22_n742 ) , .A1( us22_n784 ) );
  NOR2_X1 us22_U254 (.ZN( us22_n552 ) , .A1( us22_n784 ) , .A2( us22_n811 ) );
  NOR2_X1 us22_U255 (.ZN( us22_n515 ) , .A1( us22_n706 ) , .A2( us22_n801 ) );
  NOR2_X1 us22_U256 (.ZN( us22_n556 ) , .A1( us22_n706 ) , .A2( us22_n814 ) );
  NOR2_X1 us22_U257 (.ZN( us22_n519 ) , .A1( us22_n788 ) , .A2( us22_n810 ) );
  NOR2_X1 us22_U258 (.ZN( us22_n628 ) , .A1( us22_n745 ) , .A2( us22_n813 ) );
  NOR2_X1 us22_U259 (.ZN( us22_n713 ) , .A1( us22_n803 ) , .A2( us22_n815 ) );
  NOR4_X1 us22_U26 (.A4( us22_n539 ) , .A3( us22_n540 ) , .A2( us22_n541 ) , .ZN( us22_n548 ) , .A1( us22_n686 ) );
  AOI21_X1 us22_U260 (.ZN( us22_n569 ) , .B2( us22_n695 ) , .B1( us22_n804 ) , .A( us22_n810 ) );
  INV_X1 us22_U261 (.A( us22_n761 ) , .ZN( us22_n864 ) );
  NOR2_X1 us22_U262 (.ZN( us22_n653 ) , .A1( us22_n788 ) , .A2( us22_n813 ) );
  NOR2_X1 us22_U263 (.ZN( us22_n666 ) , .A2( us22_n706 ) , .A1( us22_n788 ) );
  NOR2_X1 us22_U264 (.ZN( us22_n654 ) , .A1( us22_n745 ) , .A2( us22_n778 ) );
  NOR2_X1 us22_U265 (.ZN( us22_n554 ) , .A1( us22_n760 ) , .A2( us22_n803 ) );
  NOR2_X1 us22_U266 (.ZN( us22_n540 ) , .A1( us22_n760 ) , .A2( us22_n789 ) );
  NOR2_X1 us22_U267 (.ZN( us22_n699 ) , .A2( us22_n784 ) , .A1( us22_n815 ) );
  NOR2_X1 us22_U268 (.ZN( us22_n607 ) , .A2( us22_n722 ) , .A1( us22_n815 ) );
  NOR2_X1 us22_U269 (.A1( us22_n728 ) , .ZN( us22_n763 ) , .A2( us22_n784 ) );
  NOR2_X1 us22_U27 (.ZN( us22_n678 ) , .A2( us22_n832 ) , .A1( us22_n837 ) );
  AOI21_X1 us22_U270 (.A( us22_n813 ) , .B2( us22_n814 ) , .B1( us22_n815 ) , .ZN( us22_n816 ) );
  INV_X1 us22_U271 (.A( us22_n727 ) , .ZN( us22_n866 ) );
  NOR2_X1 us22_U272 (.ZN( us22_n577 ) , .A2( us22_n706 ) , .A1( us22_n728 ) );
  NOR2_X1 us22_U273 (.ZN( us22_n531 ) , .A2( us22_n722 ) , .A1( us22_n728 ) );
  AOI21_X1 us22_U274 (.B1( us22_n623 ) , .ZN( us22_n625 ) , .A( us22_n761 ) , .B2( us22_n812 ) );
  AOI21_X1 us22_U275 (.A( us22_n810 ) , .B2( us22_n811 ) , .B1( us22_n812 ) , .ZN( us22_n817 ) );
  AOI21_X1 us22_U276 (.ZN( us22_n513 ) , .A( us22_n727 ) , .B1( us22_n748 ) , .B2( us22_n801 ) );
  AOI21_X1 us22_U277 (.ZN( us22_n497 ) , .B1( us22_n678 ) , .A( us22_n810 ) , .B2( us22_n814 ) );
  AOI21_X1 us22_U278 (.ZN( us22_n476 ) , .B2( us22_n695 ) , .A( us22_n747 ) , .B1( us22_n777 ) );
  NOR2_X1 us22_U279 (.ZN( us22_n580 ) , .A1( us22_n742 ) , .A2( us22_n813 ) );
  NOR4_X1 us22_U28 (.A4( us22_n512 ) , .A3( us22_n513 ) , .A2( us22_n514 ) , .A1( us22_n515 ) , .ZN( us22_n522 ) );
  NOR2_X1 us22_U280 (.ZN( us22_n640 ) , .A2( us22_n786 ) , .A1( us22_n789 ) );
  AOI21_X1 us22_U281 (.ZN( us22_n591 ) , .B1( us22_n748 ) , .A( us22_n790 ) , .B2( us22_n811 ) );
  NOR2_X1 us22_U282 (.A2( us22_n706 ) , .A1( us22_n760 ) , .ZN( us22_n792 ) );
  AOI21_X1 us22_U283 (.ZN( us22_n624 ) , .B2( us22_n667 ) , .A( us22_n788 ) , .B1( us22_n789 ) );
  NOR2_X1 us22_U284 (.ZN( us22_n668 ) , .A1( us22_n788 ) , .A2( us22_n803 ) );
  NOR2_X1 us22_U285 (.ZN( us22_n518 ) , .A2( us22_n706 ) , .A1( us22_n812 ) );
  AOI21_X1 us22_U286 (.ZN( us22_n475 ) , .A( us22_n667 ) , .B1( us22_n748 ) , .B2( us22_n804 ) );
  NOR2_X1 us22_U287 (.ZN( us22_n557 ) , .A2( us22_n789 ) , .A1( us22_n801 ) );
  NOR2_X1 us22_U288 (.ZN( us22_n517 ) , .A2( us22_n697 ) , .A1( us22_n814 ) );
  NOR2_X1 us22_U289 (.ZN( us22_n681 ) , .A2( us22_n697 ) , .A1( us22_n801 ) );
  AOI222_X1 us22_U29 (.ZN( us22_n523 ) , .A1( us22_n832 ) , .B2( us22_n835 ) , .C1( us22_n842 ) , .C2( us22_n848 ) , .A2( us22_n850 ) , .B1( us22_n864 ) );
  NOR2_X1 us22_U290 (.ZN( us22_n651 ) , .A1( us22_n760 ) , .A2( us22_n784 ) );
  INV_X1 us22_U291 (.A( us22_n811 ) , .ZN( us22_n834 ) );
  AOI21_X1 us22_U292 (.ZN( us22_n508 ) , .B2( us22_n667 ) , .A( us22_n728 ) , .B1( us22_n813 ) );
  AOI21_X1 us22_U293 (.ZN( us22_n537 ) , .B2( us22_n810 ) , .A( us22_n812 ) , .B1( us22_n813 ) );
  AOI21_X1 us22_U294 (.ZN( us22_n538 ) , .A( us22_n761 ) , .B2( us22_n777 ) , .B1( us22_n815 ) );
  NOR2_X1 us22_U295 (.ZN( us22_n579 ) , .A1( us22_n667 ) , .A2( us22_n786 ) );
  AOI21_X1 us22_U296 (.ZN( us22_n587 ) , .B2( us22_n697 ) , .B1( us22_n813 ) , .A( us22_n815 ) );
  AOI21_X1 us22_U297 (.B1( us22_n697 ) , .ZN( us22_n698 ) , .A( us22_n730 ) , .B2( us22_n761 ) );
  AOI21_X1 us22_U298 (.ZN( us22_n589 ) , .B2( us22_n761 ) , .A( us22_n783 ) , .B1( us22_n810 ) );
  AOI21_X1 us22_U299 (.ZN( us22_n496 ) , .A( us22_n722 ) , .B2( us22_n760 ) , .B1( us22_n812 ) );
  NAND2_X2 us22_U3 (.A1( us22_n445 ) , .A2( us22_n446 ) , .ZN( us22_n784 ) );
  NOR4_X1 us22_U30 (.A3( us22_n519 ) , .A1( us22_n520 ) , .ZN( us22_n521 ) , .A2( us22_n671 ) , .A4( us22_n767 ) );
  AOI21_X1 us22_U300 (.ZN( us22_n550 ) , .B1( us22_n667 ) , .A( us22_n695 ) , .B2( us22_n803 ) );
  NOR2_X1 us22_U301 (.ZN( us22_n545 ) , .A1( us22_n697 ) , .A2( us22_n742 ) );
  INV_X1 us22_U302 (.A( us22_n789 ) , .ZN( us22_n871 ) );
  INV_X1 us22_U303 (.A( us22_n810 ) , .ZN( us22_n852 ) );
  AOI21_X1 us22_U304 (.ZN( us22_n638 ) , .B2( us22_n745 ) , .A( us22_n790 ) , .B1( us22_n801 ) );
  AOI21_X1 us22_U305 (.ZN( us22_n647 ) , .B1( us22_n727 ) , .B2( us22_n761 ) , .A( us22_n811 ) );
  NOR2_X1 us22_U306 (.ZN( us22_n683 ) , .A1( us22_n727 ) , .A2( us22_n814 ) );
  AOI21_X1 us22_U307 (.B1( us22_n684 ) , .ZN( us22_n685 ) , .A( us22_n726 ) , .B2( us22_n759 ) );
  AOI21_X1 us22_U308 (.ZN( us22_n567 ) , .B1( us22_n748 ) , .B2( us22_n760 ) , .A( us22_n778 ) );
  AOI21_X1 us22_U309 (.ZN( us22_n498 ) , .A( us22_n695 ) , .B1( us22_n706 ) , .B2( us22_n784 ) );
  AOI221_X1 us22_U31 (.A( us22_n779 ) , .ZN( us22_n796 ) , .C2( us22_n835 ) , .B2( us22_n836 ) , .B1( us22_n863 ) , .C1( us22_n864 ) );
  NOR2_X1 us22_U310 (.ZN( us22_n566 ) , .A1( us22_n727 ) , .A2( us22_n760 ) );
  AOI21_X1 us22_U311 (.ZN( us22_n637 ) , .B2( us22_n747 ) , .A( us22_n786 ) , .B1( us22_n810 ) );
  NOR2_X1 us22_U312 (.ZN( us22_n564 ) , .A2( us22_n695 ) , .A1( us22_n761 ) );
  NOR2_X1 us22_U313 (.ZN( us22_n578 ) , .A2( us22_n695 ) , .A1( us22_n789 ) );
  AOI21_X1 us22_U314 (.ZN( us22_n512 ) , .A( us22_n777 ) , .B2( us22_n790 ) , .B1( us22_n810 ) );
  INV_X1 us22_U315 (.A( us22_n697 ) , .ZN( us22_n851 ) );
  NOR2_X1 us22_U316 (.ZN( us22_n663 ) , .A1( us22_n778 ) , .A2( us22_n811 ) );
  AOI21_X1 us22_U317 (.ZN( us22_n448 ) , .B2( us22_n790 ) , .A( us22_n801 ) , .B1( us22_n813 ) );
  NOR2_X1 us22_U318 (.ZN( us22_n630 ) , .A2( us22_n695 ) , .A1( us22_n722 ) );
  AOI21_X1 us22_U319 (.ZN( us22_n562 ) , .B1( us22_n722 ) , .A( us22_n777 ) , .B2( us22_n789 ) );
  NOR4_X1 us22_U32 (.A4( us22_n791 ) , .A3( us22_n792 ) , .A2( us22_n793 ) , .A1( us22_n794 ) , .ZN( us22_n795 ) );
  AOI21_X1 us22_U320 (.ZN( us22_n495 ) , .A( us22_n777 ) , .B2( us22_n789 ) , .B1( us22_n802 ) );
  AOI21_X1 us22_U321 (.ZN( us22_n687 ) , .B2( us22_n747 ) , .B1( us22_n761 ) , .A( us22_n804 ) );
  NOR2_X1 us22_U322 (.ZN( us22_n527 ) , .A1( us22_n706 ) , .A2( us22_n777 ) );
  NOR2_X1 us22_U323 (.ZN( us22_n576 ) , .A1( us22_n706 ) , .A2( us22_n811 ) );
  AOI21_X1 us22_U324 (.ZN( us22_n648 ) , .A( us22_n777 ) , .B1( us22_n790 ) , .B2( us22_n803 ) );
  NOR2_X1 us22_U325 (.ZN( us22_n682 ) , .A1( us22_n789 ) , .A2( us22_n811 ) );
  NOR2_X1 us22_U326 (.A2( us22_n811 ) , .A1( us22_n813 ) , .ZN( us22_n819 ) );
  AOI21_X1 us22_U327 (.A( us22_n788 ) , .B2( us22_n789 ) , .B1( us22_n790 ) , .ZN( us22_n791 ) );
  AOI21_X1 us22_U328 (.A( us22_n731 ) , .ZN( us22_n732 ) , .B2( us22_n778 ) , .B1( us22_n790 ) );
  NOR2_X1 us22_U329 (.ZN( us22_n565 ) , .A1( us22_n745 ) , .A2( us22_n803 ) );
  NOR4_X1 us22_U33 (.A4( us22_n774 ) , .A3( us22_n775 ) , .A1( us22_n776 ) , .ZN( us22_n797 ) , .A2( us22_n799 ) );
  NOR2_X1 us22_U330 (.ZN( us22_n581 ) , .A1( us22_n790 ) , .A2( us22_n815 ) );
  NOR2_X1 us22_U331 (.ZN( us22_n532 ) , .A1( us22_n722 ) , .A2( us22_n786 ) );
  AOI21_X1 us22_U332 (.ZN( us22_n639 ) , .B1( us22_n678 ) , .A( us22_n789 ) , .B2( us22_n815 ) );
  NOR2_X1 us22_U333 (.ZN( us22_n709 ) , .A1( us22_n760 ) , .A2( us22_n761 ) );
  NOR2_X1 us22_U334 (.ZN( us22_n680 ) , .A2( us22_n706 ) , .A1( us22_n815 ) );
  INV_X1 us22_U335 (.A( us22_n695 ) , .ZN( us22_n836 ) );
  INV_X1 us22_U336 (.A( us22_n813 ) , .ZN( us22_n853 ) );
  AOI21_X1 us22_U337 (.ZN( us22_n440 ) , .A( us22_n697 ) , .B1( us22_n731 ) , .B2( us22_n748 ) );
  OAI21_X1 us22_U338 (.A( us22_n696 ) , .ZN( us22_n700 ) , .B2( us22_n748 ) , .B1( us22_n802 ) );
  OAI21_X1 us22_U339 (.ZN( us22_n696 ) , .B2( us22_n831 ) , .B1( us22_n836 ) , .A( us22_n858 ) );
  NOR4_X1 us22_U34 (.A3( us22_n753 ) , .A2( us22_n754 ) , .A1( us22_n755 ) , .ZN( us22_n756 ) , .A4( us22_n867 ) );
  NAND2_X1 us22_U340 (.ZN( us22_n751 ) , .A1( us22_n761 ) , .A2( us22_n803 ) );
  INV_X1 us22_U341 (.A( us22_n778 ) , .ZN( us22_n848 ) );
  INV_X1 us22_U342 (.A( us22_n783 ) , .ZN( us22_n844 ) );
  NAND2_X1 us22_U343 (.ZN( us22_n669 ) , .A1( us22_n804 ) , .A2( us22_n814 ) );
  NAND2_X1 us22_U344 (.ZN( us22_n712 ) , .A1( us22_n726 ) , .A2( us22_n778 ) );
  NAND2_X1 us22_U345 (.A2( us22_n760 ) , .A1( us22_n804 ) , .ZN( us22_n808 ) );
  NAND2_X2 us22_U346 (.A2( us22_n439 ) , .A1( us22_n445 ) , .ZN( us22_n782 ) );
  AOI21_X1 us22_U347 (.ZN( us22_n441 ) , .B1( us22_n787 ) , .B2( us22_n789 ) , .A( us22_n812 ) );
  NOR2_X1 us22_U348 (.ZN( us22_n468 ) , .A2( us22_n777 ) , .A1( us22_n813 ) );
  OAI21_X1 us22_U349 (.A( us22_n785 ) , .B2( us22_n786 ) , .B1( us22_n787 ) , .ZN( us22_n793 ) );
  AOI211_X1 us22_U35 (.B( us22_n743 ) , .A( us22_n744 ) , .ZN( us22_n757 ) , .C1( us22_n830 ) , .C2( us22_n851 ) );
  OAI21_X1 us22_U350 (.ZN( us22_n785 ) , .A( us22_n837 ) , .B1( us22_n861 ) , .B2( us22_n871 ) );
  NOR2_X1 us22_U351 (.ZN( us22_n524 ) , .A1( us22_n722 ) , .A2( us22_n748 ) );
  NOR2_X1 us22_U352 (.ZN( us22_n710 ) , .A2( us22_n722 ) , .A1( us22_n788 ) );
  NOR2_X1 us22_U353 (.ZN( us22_n482 ) , .A1( us22_n786 ) , .A2( us22_n803 ) );
  NAND2_X1 us22_U354 (.A1( us22_n697 ) , .A2( us22_n727 ) , .ZN( us22_n780 ) );
  NOR2_X1 us22_U355 (.ZN( us22_n516 ) , .A1( us22_n706 ) , .A2( us22_n786 ) );
  NAND2_X1 us22_U356 (.A2( us22_n747 ) , .A1( us22_n784 ) , .ZN( us22_n807 ) );
  OAI21_X1 us22_U357 (.A( us22_n729 ) , .B1( us22_n730 ) , .ZN( us22_n734 ) , .B2( us22_n803 ) );
  OAI21_X1 us22_U358 (.ZN( us22_n729 ) , .A( us22_n831 ) , .B2( us22_n850 ) , .B1( us22_n871 ) );
  INV_X1 us22_U359 (.A( us22_n815 ) , .ZN( us22_n842 ) );
  NOR3_X1 us22_U36 (.A3( us22_n739 ) , .A2( us22_n740 ) , .A1( us22_n741 ) , .ZN( us22_n758 ) );
  INV_X1 us22_U360 (.A( us22_n722 ) , .ZN( us22_n854 ) );
  AND2_X1 us22_U361 (.ZN( us22_n730 ) , .A1( us22_n777 ) , .A2( us22_n783 ) );
  AOI221_X1 us22_U362 (.A( us22_n762 ) , .ZN( us22_n772 ) , .C2( us22_n808 ) , .B2( us22_n833 ) , .C1( us22_n853 ) , .B1( us22_n864 ) );
  AOI21_X1 us22_U363 (.B2( us22_n761 ) , .ZN( us22_n762 ) , .A( us22_n786 ) , .B1( us22_n790 ) );
  INV_X1 us22_U364 (.A( us22_n759 ) , .ZN( us22_n833 ) );
  NAND2_X1 us22_U365 (.A1( us22_n453 ) , .A2( us22_n469 ) , .ZN( us22_n801 ) );
  NAND2_X1 us22_U366 (.A1( us22_n449 ) , .A2( us22_n452 ) , .ZN( us22_n812 ) );
  NAND2_X1 us22_U367 (.A1( us22_n449 ) , .A2( us22_n469 ) , .ZN( us22_n814 ) );
  NAND2_X1 us22_U368 (.A1( us22_n452 ) , .A2( us22_n459 ) , .ZN( us22_n811 ) );
  NAND2_X1 us22_U369 (.A1( us22_n451 ) , .A2( us22_n459 ) , .ZN( us22_n742 ) );
  NOR4_X1 us22_U37 (.A4( us22_n732 ) , .A3( us22_n733 ) , .A2( us22_n734 ) , .A1( us22_n735 ) , .ZN( us22_n736 ) );
  NAND2_X1 us22_U370 (.A1( us22_n450 ) , .A2( us22_n463 ) , .ZN( us22_n667 ) );
  NAND2_X1 us22_U371 (.A2( us22_n446 ) , .A1( us22_n458 ) , .ZN( us22_n726 ) );
  NAND2_X1 us22_U372 (.A1( us22_n453 ) , .A2( us22_n460 ) , .ZN( us22_n748 ) );
  NAND2_X1 us22_U373 (.A2( us22_n451 ) , .A1( us22_n453 ) , .ZN( us22_n804 ) );
  NAND2_X1 us22_U374 (.A2( us22_n452 ) , .A1( us22_n470 ) , .ZN( us22_n777 ) );
  NAND2_X1 us22_U375 (.A1( us22_n451 ) , .A2( us22_n470 ) , .ZN( us22_n783 ) );
  NAND2_X1 us22_U376 (.A2( us22_n462 ) , .A1( us22_n463 ) , .ZN( us22_n810 ) );
  NAND2_X1 us22_U377 (.A1( us22_n439 ) , .A2( us22_n458 ) , .ZN( us22_n697 ) );
  NAND2_X1 us22_U378 (.A2( us22_n447 ) , .A1( us22_n450 ) , .ZN( us22_n761 ) );
  NAND2_X1 us22_U379 (.A2( us22_n446 ) , .A1( us22_n450 ) , .ZN( us22_n727 ) );
  AOI211_X1 us22_U38 (.B( us22_n723 ) , .A( us22_n724 ) , .ZN( us22_n737 ) , .C1( us22_n841 ) , .C2( us22_n853 ) );
  NAND2_X2 us22_U380 (.A2( us22_n459 ) , .A1( us22_n469 ) , .ZN( us22_n695 ) );
  NOR2_X1 us22_U381 (.ZN( us22_n445 ) , .A2( us22_n847 ) , .A1( us22_n856 ) );
  NAND2_X1 us22_U382 (.A2( us22_n459 ) , .A1( us22_n460 ) , .ZN( us22_n745 ) );
  NAND2_X1 us22_U383 (.A1( us22_n460 ) , .A2( us22_n470 ) , .ZN( us22_n786 ) );
  NOR2_X1 us22_U384 (.ZN( us22_n463 ) , .A2( us22_n845 ) , .A1( us22_n846 ) );
  NOR2_X1 us22_U385 (.ZN( us22_n451 ) , .A1( us22_n824 ) , .A2( us22_n825 ) );
  NOR2_X1 us22_U386 (.ZN( us22_n449 ) , .A1( us22_n826 ) , .A2( us22_n827 ) );
  NAND2_X1 us22_U387 (.A2( us22_n452 ) , .A1( us22_n453 ) , .ZN( us22_n728 ) );
  NAND2_X1 us22_U388 (.A1( us22_n449 ) , .A2( us22_n460 ) , .ZN( us22_n788 ) );
  NAND2_X2 us22_U389 (.A2( us22_n446 ) , .A1( us22_n462 ) , .ZN( us22_n813 ) );
  NOR3_X1 us22_U39 (.A3( us22_n720 ) , .A1( us22_n721 ) , .ZN( us22_n738 ) , .A2( us22_n739 ) );
  NAND2_X2 us22_U390 (.A2( us22_n439 ) , .A1( us22_n450 ) , .ZN( us22_n789 ) );
  NAND2_X2 us22_U391 (.A1( us22_n447 ) , .A2( us22_n462 ) , .ZN( us22_n722 ) );
  NAND2_X2 us22_U392 (.A1( us22_n447 ) , .A2( us22_n458 ) , .ZN( us22_n790 ) );
  NAND2_X2 us22_U393 (.A1( us22_n439 ) , .A2( us22_n462 ) , .ZN( us22_n706 ) );
  NAND2_X2 us22_U394 (.A2( us22_n469 ) , .A1( us22_n470 ) , .ZN( us22_n815 ) );
  NAND2_X2 us22_U395 (.A2( us22_n458 ) , .A1( us22_n463 ) , .ZN( us22_n778 ) );
  NAND2_X1 us22_U396 (.A1( us22_n445 ) , .A2( us22_n447 ) , .ZN( us22_n803 ) );
  NOR2_X1 us22_U397 (.A2( sa22_6 ) , .A1( sa22_7 ) , .ZN( us22_n462 ) );
  NOR2_X1 us22_U398 (.A2( sa22_4 ) , .ZN( us22_n447 ) , .A1( us22_n846 ) );
  NOR2_X1 us22_U399 (.A2( sa22_5 ) , .ZN( us22_n446 ) , .A1( us22_n845 ) );
  INV_X1 us22_U4 (.A( us22_n784 ) , .ZN( us22_n860 ) );
  NAND4_X1 us22_U40 (.ZN( sa20_sr_3 ) , .A4( us22_n702 ) , .A3( us22_n703 ) , .A2( us22_n704 ) , .A1( us22_n705 ) );
  NOR2_X1 us22_U400 (.A2( sa22_7 ) , .ZN( us22_n458 ) , .A1( us22_n847 ) );
  NOR2_X1 us22_U401 (.A2( sa22_4 ) , .A1( sa22_5 ) , .ZN( us22_n439 ) );
  NOR2_X1 us22_U402 (.A2( sa22_1 ) , .ZN( us22_n469 ) , .A1( us22_n824 ) );
  NOR2_X1 us22_U403 (.A2( sa22_2 ) , .A1( sa22_3 ) , .ZN( us22_n470 ) );
  NOR2_X1 us22_U404 (.A2( sa22_6 ) , .ZN( us22_n450 ) , .A1( us22_n856 ) );
  NOR2_X1 us22_U405 (.A2( sa22_2 ) , .ZN( us22_n459 ) , .A1( us22_n827 ) );
  NOR2_X1 us22_U406 (.A2( sa22_0 ) , .ZN( us22_n452 ) , .A1( us22_n825 ) );
  NOR2_X1 us22_U407 (.A2( sa22_0 ) , .A1( sa22_1 ) , .ZN( us22_n460 ) );
  NOR2_X1 us22_U408 (.A2( sa22_3 ) , .ZN( us22_n453 ) , .A1( us22_n826 ) );
  INV_X1 us22_U409 (.A( sa22_6 ) , .ZN( us22_n847 ) );
  NOR4_X1 us22_U41 (.A4( us22_n698 ) , .A3( us22_n699 ) , .A2( us22_n700 ) , .A1( us22_n701 ) , .ZN( us22_n702 ) );
  INV_X1 us22_U410 (.A( sa22_3 ) , .ZN( us22_n827 ) );
  INV_X1 us22_U411 (.A( sa22_1 ) , .ZN( us22_n825 ) );
  INV_X1 us22_U412 (.A( sa22_2 ) , .ZN( us22_n826 ) );
  INV_X1 us22_U413 (.A( sa22_0 ) , .ZN( us22_n824 ) );
  INV_X1 us22_U414 (.A( sa22_7 ) , .ZN( us22_n856 ) );
  INV_X1 us22_U415 (.A( sa22_5 ) , .ZN( us22_n846 ) );
  OAI221_X1 us22_U416 (.A( us22_n781 ) , .C2( us22_n782 ) , .B2( us22_n783 ) , .B1( us22_n784 ) , .ZN( us22_n794 ) , .C1( us22_n811 ) );
  NAND2_X1 us22_U417 (.A1( us22_n727 ) , .A2( us22_n782 ) , .ZN( us22_n809 ) );
  OAI22_X1 us22_U418 (.ZN( us22_n586 ) , .A2( us22_n745 ) , .B2( us22_n760 ) , .A1( us22_n761 ) , .B1( us22_n782 ) );
  OAI221_X1 us22_U419 (.A( us22_n694 ) , .ZN( us22_n701 ) , .C2( us22_n782 ) , .C1( us22_n783 ) , .B1( us22_n784 ) , .B2( us22_n804 ) );
  AOI211_X1 us22_U42 (.B( us22_n692 ) , .A( us22_n693 ) , .ZN( us22_n703 ) , .C2( us22_n829 ) , .C1( us22_n849 ) );
  AOI21_X1 us22_U420 (.ZN( us22_n590 ) , .B1( us22_n726 ) , .B2( us22_n782 ) , .A( us22_n788 ) );
  AOI21_X1 us22_U421 (.ZN( us22_n621 ) , .B1( us22_n697 ) , .A( us22_n777 ) , .B2( us22_n782 ) );
  AOI21_X1 us22_U422 (.ZN( us22_n646 ) , .A( us22_n760 ) , .B2( us22_n782 ) , .B1( us22_n790 ) );
  OAI22_X1 us22_U423 (.ZN( us22_n679 ) , .A1( us22_n697 ) , .A2( us22_n728 ) , .B2( us22_n782 ) , .B1( us22_n815 ) );
  OAI21_X1 us22_U424 (.A( us22_n611 ) , .ZN( us22_n614 ) , .B1( us22_n623 ) , .B2( us22_n782 ) );
  NOR2_X1 us22_U425 (.ZN( us22_n608 ) , .A1( us22_n782 ) , .A2( us22_n814 ) );
  OAI222_X1 us22_U426 (.A2( us22_n667 ) , .ZN( us22_n672 ) , .B1( us22_n745 ) , .B2( us22_n782 ) , .C2( us22_n786 ) , .C1( us22_n813 ) , .A1( us22_n815 ) );
  NOR2_X1 us22_U427 (.ZN( us22_n649 ) , .A1( us22_n782 ) , .A2( us22_n786 ) );
  NOR2_X1 us22_U428 (.ZN( us22_n598 ) , .A2( us22_n695 ) , .A1( us22_n782 ) );
  NOR2_X1 us22_U429 (.ZN( us22_n551 ) , .A2( us22_n742 ) , .A1( us22_n782 ) );
  NOR2_X1 us22_U43 (.ZN( us22_n705 ) , .A2( us22_n774 ) , .A1( us22_n798 ) );
  INV_X1 us22_U430 (.A( us22_n782 ) , .ZN( us22_n859 ) );
  NAND4_X1 us22_U431 (.ZN( sa20_sr_2 ) , .A4( us22_n641 ) , .A3( us22_n642 ) , .A1( us22_n643 ) , .A2( us22_n644 ) );
  AOI221_X1 us22_U432 (.A( us22_n574 ) , .ZN( us22_n585 ) , .B2( us22_n829 ) , .C2( us22_n841 ) , .B1( us22_n852 ) , .C1( us22_n859 ) );
  AOI21_X1 us22_U433 (.ZN( us22_n574 ) , .B2( us22_n722 ) , .B1( us22_n746 ) , .A( us22_n783 ) );
  AOI211_X1 us22_U434 (.A( us22_n635 ) , .ZN( us22_n643 ) , .B( us22_n741 ) , .C2( us22_n837 ) , .C1( us22_n852 ) );
  NAND4_X1 us22_U435 (.A4( us22_n631 ) , .A3( us22_n632 ) , .A2( us22_n633 ) , .A1( us22_n634 ) , .ZN( us22_n741 ) );
  INV_X1 us22_U436 (.A( sa22_4 ) , .ZN( us22_n845 ) );
  NAND3_X1 us22_U437 (.ZN( sa20_sr_6 ) , .A3( us22_n795 ) , .A2( us22_n796 ) , .A1( us22_n797 ) );
  NAND3_X1 us22_U438 (.ZN( sa20_sr_5 ) , .A3( us22_n756 ) , .A2( us22_n757 ) , .A1( us22_n758 ) );
  NAND3_X1 us22_U439 (.ZN( sa20_sr_4 ) , .A3( us22_n736 ) , .A2( us22_n737 ) , .A1( us22_n738 ) );
  AOI222_X1 us22_U44 (.B2( us22_n636 ) , .ZN( us22_n642 ) , .B1( us22_n839 ) , .A1( us22_n840 ) , .C2( us22_n844 ) , .C1( us22_n861 ) , .A2( us22_n863 ) );
  NAND3_X1 us22_U440 (.A3( us22_n673 ) , .A2( us22_n674 ) , .A1( us22_n675 ) , .ZN( us22_n805 ) );
  NAND3_X1 us22_U441 (.ZN( us22_n636 ) , .A3( us22_n706 ) , .A2( us22_n722 ) , .A1( us22_n790 ) );
  NAND3_X1 us22_U442 (.A3( us22_n616 ) , .A2( us22_n617 ) , .A1( us22_n618 ) , .ZN( us22_n723 ) );
  NAND3_X1 us22_U443 (.A3( us22_n583 ) , .A2( us22_n584 ) , .A1( us22_n585 ) , .ZN( us22_n619 ) );
  NAND3_X1 us22_U444 (.ZN( us22_n563 ) , .A3( us22_n678 ) , .A2( us22_n748 ) , .A1( us22_n783 ) );
  NAND3_X1 us22_U445 (.A3( us22_n521 ) , .A2( us22_n522 ) , .A1( us22_n523 ) , .ZN( us22_n740 ) );
  NAND3_X1 us22_U446 (.A3( us22_n510 ) , .A1( us22_n511 ) , .ZN( us22_n606 ) , .A2( us22_n869 ) );
  NAND3_X1 us22_U447 (.A3( us22_n465 ) , .A2( us22_n466 ) , .A1( us22_n467 ) , .ZN( us22_n775 ) );
  NOR4_X1 us22_U45 (.A4( us22_n637 ) , .A3( us22_n638 ) , .A2( us22_n639 ) , .A1( us22_n640 ) , .ZN( us22_n641 ) );
  NOR3_X1 us22_U46 (.A2( us22_n605 ) , .A1( us22_n606 ) , .ZN( us22_n644 ) , .A3( us22_n720 ) );
  NOR2_X1 us22_U47 (.ZN( us22_n802 ) , .A1( us22_n852 ) , .A2( us22_n859 ) );
  NAND4_X1 us22_U48 (.ZN( sa20_sr_7 ) , .A4( us22_n820 ) , .A3( us22_n821 ) , .A2( us22_n822 ) , .A1( us22_n823 ) );
  NOR4_X1 us22_U49 (.A4( us22_n816 ) , .A3( us22_n817 ) , .A2( us22_n818 ) , .A1( us22_n819 ) , .ZN( us22_n820 ) );
  NOR3_X1 us22_U5 (.ZN( us22_n596 ) , .A1( us22_n606 ) , .A3( us22_n721 ) , .A2( us22_n740 ) );
  AOI222_X1 us22_U50 (.C2( us22_n807 ) , .B2( us22_n808 ) , .A2( us22_n809 ) , .ZN( us22_n821 ) , .C1( us22_n830 ) , .A1( us22_n837 ) , .B1( us22_n851 ) );
  AOI211_X1 us22_U51 (.B( us22_n805 ) , .A( us22_n806 ) , .ZN( us22_n822 ) , .C1( us22_n840 ) , .C2( us22_n848 ) );
  NAND4_X1 us22_U52 (.ZN( sa20_sr_0 ) , .A4( us22_n499 ) , .A3( us22_n500 ) , .A2( us22_n501 ) , .A1( us22_n502 ) );
  AOI221_X1 us22_U53 (.A( us22_n495 ) , .ZN( us22_n500 ) , .B2( us22_n841 ) , .C1( us22_n844 ) , .C2( us22_n858 ) , .B1( us22_n860 ) );
  NOR4_X1 us22_U54 (.A4( us22_n496 ) , .A3( us22_n497 ) , .A2( us22_n498 ) , .ZN( us22_n499 ) , .A1( us22_n525 ) );
  AOI211_X1 us22_U55 (.A( us22_n494 ) , .ZN( us22_n501 ) , .B( us22_n800 ) , .C2( us22_n837 ) , .C1( us22_n849 ) );
  NOR2_X1 us22_U56 (.ZN( us22_n746 ) , .A1( us22_n859 ) , .A2( us22_n860 ) );
  NAND4_X1 us22_U57 (.ZN( sa20_sr_1 ) , .A4( us22_n593 ) , .A3( us22_n594 ) , .A2( us22_n595 ) , .A1( us22_n596 ) );
  NOR4_X1 us22_U58 (.A4( us22_n589 ) , .A3( us22_n590 ) , .A2( us22_n591 ) , .A1( us22_n592 ) , .ZN( us22_n593 ) );
  AOI211_X1 us22_U59 (.B( us22_n587 ) , .A( us22_n588 ) , .ZN( us22_n594 ) , .C2( us22_n809 ) , .C1( us22_n831 ) );
  NOR3_X1 us22_U6 (.A3( us22_n798 ) , .A2( us22_n799 ) , .A1( us22_n800 ) , .ZN( us22_n823 ) );
  AOI211_X1 us22_U60 (.A( us22_n586 ) , .ZN( us22_n595 ) , .B( us22_n619 ) , .C1( us22_n843 ) , .C2( us22_n853 ) );
  NOR2_X1 us22_U61 (.ZN( us22_n623 ) , .A2( us22_n834 ) , .A1( us22_n837 ) );
  AOI222_X1 us22_U62 (.ZN( us22_n467 ) , .B1( us22_n830 ) , .A1( us22_n837 ) , .C1( us22_n840 ) , .C2( us22_n849 ) , .A2( us22_n853 ) , .B2( us22_n863 ) );
  NOR4_X1 us22_U63 (.A1( us22_n464 ) , .ZN( us22_n465 ) , .A4( us22_n540 ) , .A2( us22_n552 ) , .A3( us22_n612 ) );
  AOI221_X1 us22_U64 (.ZN( us22_n466 ) , .C2( us22_n712 ) , .B2( us22_n829 ) , .C1( us22_n843 ) , .B1( us22_n858 ) , .A( us22_n862 ) );
  NAND4_X1 us22_U65 (.A4( us22_n601 ) , .A3( us22_n602 ) , .A2( us22_n603 ) , .A1( us22_n604 ) , .ZN( us22_n720 ) );
  NOR3_X1 us22_U66 (.A1( us22_n597 ) , .ZN( us22_n602 ) , .A3( us22_n661 ) , .A2( us22_n768 ) );
  NOR4_X1 us22_U67 (.A3( us22_n598 ) , .A2( us22_n599 ) , .A1( us22_n600 ) , .ZN( us22_n601 ) , .A4( us22_n653 ) );
  AOI222_X1 us22_U68 (.ZN( us22_n604 ) , .A1( us22_n828 ) , .C2( us22_n835 ) , .B1( us22_n840 ) , .A2( us22_n854 ) , .B2( us22_n859 ) , .C1( us22_n866 ) );
  NOR4_X1 us22_U69 (.A4( us22_n575 ) , .A3( us22_n576 ) , .A2( us22_n577 ) , .ZN( us22_n584 ) , .A1( us22_n681 ) );
  NOR3_X1 us22_U7 (.ZN( us22_n502 ) , .A2( us22_n677 ) , .A3( us22_n775 ) , .A1( us22_n874 ) );
  NOR4_X1 us22_U70 (.A1( us22_n582 ) , .ZN( us22_n583 ) , .A3( us22_n650 ) , .A2( us22_n660 ) , .A4( us22_n765 ) );
  AOI211_X1 us22_U71 (.B( us22_n621 ) , .A( us22_n622 ) , .ZN( us22_n633 ) , .C2( us22_n834 ) , .C1( us22_n861 ) );
  NOR4_X1 us22_U72 (.A4( us22_n627 ) , .A3( us22_n628 ) , .A2( us22_n629 ) , .A1( us22_n630 ) , .ZN( us22_n631 ) );
  NOR4_X1 us22_U73 (.A4( us22_n624 ) , .A3( us22_n625 ) , .A2( us22_n626 ) , .ZN( us22_n632 ) , .A1( us22_n662 ) );
  NAND4_X1 us22_U74 (.A4( us22_n655 ) , .A3( us22_n656 ) , .A2( us22_n657 ) , .A1( us22_n658 ) , .ZN( us22_n798 ) );
  NOR3_X1 us22_U75 (.A3( us22_n646 ) , .A2( us22_n647 ) , .A1( us22_n648 ) , .ZN( us22_n657 ) );
  NOR3_X1 us22_U76 (.A3( us22_n649 ) , .A2( us22_n650 ) , .A1( us22_n651 ) , .ZN( us22_n656 ) );
  NOR3_X1 us22_U77 (.A3( us22_n652 ) , .A2( us22_n653 ) , .A1( us22_n654 ) , .ZN( us22_n655 ) );
  NAND4_X1 us22_U78 (.A4( us22_n558 ) , .A3( us22_n559 ) , .A2( us22_n560 ) , .A1( us22_n561 ) , .ZN( us22_n605 ) );
  NOR4_X1 us22_U79 (.A4( us22_n554 ) , .A3( us22_n555 ) , .A2( us22_n556 ) , .A1( us22_n557 ) , .ZN( us22_n558 ) );
  INV_X1 us22_U8 (.A( us22_n704 ) , .ZN( us22_n874 ) );
  NOR4_X1 us22_U80 (.ZN( us22_n559 ) , .A1( us22_n651 ) , .A3( us22_n659 ) , .A4( us22_n683 ) , .A2( us22_n766 ) );
  NOR4_X1 us22_U81 (.A4( us22_n550 ) , .A3( us22_n551 ) , .A2( us22_n552 ) , .A1( us22_n553 ) , .ZN( us22_n560 ) );
  NAND4_X1 us22_U82 (.A4( us22_n770 ) , .A3( us22_n771 ) , .A2( us22_n772 ) , .A1( us22_n773 ) , .ZN( us22_n799 ) );
  NOR3_X1 us22_U83 (.A3( us22_n763 ) , .A2( us22_n764 ) , .A1( us22_n765 ) , .ZN( us22_n771 ) );
  NOR4_X1 us22_U84 (.A4( us22_n766 ) , .A3( us22_n767 ) , .A2( us22_n768 ) , .A1( us22_n769 ) , .ZN( us22_n770 ) );
  AOI222_X1 us22_U85 (.ZN( us22_n773 ) , .A1( us22_n828 ) , .C1( us22_n832 ) , .B2( us22_n839 ) , .A2( us22_n848 ) , .B1( us22_n859 ) , .C2( us22_n871 ) );
  NOR4_X1 us22_U86 (.A4( us22_n663 ) , .A3( us22_n664 ) , .A2( us22_n665 ) , .A1( us22_n666 ) , .ZN( us22_n674 ) );
  NOR4_X1 us22_U87 (.A4( us22_n659 ) , .A3( us22_n660 ) , .A2( us22_n661 ) , .A1( us22_n662 ) , .ZN( us22_n675 ) );
  NOR4_X1 us22_U88 (.A3( us22_n671 ) , .A1( us22_n672 ) , .ZN( us22_n673 ) , .A4( us22_n713 ) , .A2( us22_n857 ) );
  NOR2_X1 us22_U89 (.ZN( us22_n759 ) , .A1( us22_n831 ) , .A2( us22_n832 ) );
  NOR3_X1 us22_U9 (.A3( us22_n619 ) , .A2( us22_n620 ) , .ZN( us22_n634 ) , .A1( us22_n723 ) );
  AOI222_X1 us22_U90 (.ZN( us22_n511 ) , .C1( us22_n830 ) , .B2( us22_n835 ) , .A2( us22_n841 ) , .C2( us22_n860 ) , .B1( us22_n861 ) , .A1( us22_n864 ) );
  NOR4_X1 us22_U91 (.A4( us22_n507 ) , .A2( us22_n508 ) , .A1( us22_n509 ) , .ZN( us22_n510 ) , .A3( us22_n668 ) );
  INV_X1 us22_U92 (.A( us22_n503 ) , .ZN( us22_n869 ) );
  NAND4_X1 us22_U93 (.A4( us22_n454 ) , .A3( us22_n455 ) , .A2( us22_n456 ) , .A1( us22_n457 ) , .ZN( us22_n677 ) );
  NOR3_X1 us22_U94 (.ZN( us22_n455 ) , .A3( us22_n528 ) , .A1( us22_n553 ) , .A2( us22_n568 ) );
  AOI221_X1 us22_U95 (.A( us22_n448 ) , .ZN( us22_n457 ) , .C2( us22_n751 ) , .B1( us22_n830 ) , .C1( us22_n840 ) , .B2( us22_n859 ) );
  NOR4_X1 us22_U96 (.ZN( us22_n456 ) , .A2( us22_n507 ) , .A1( us22_n597 ) , .A4( us22_n626 ) , .A3( us22_n709 ) );
  NAND4_X1 us22_U97 (.A4( us22_n533 ) , .A3( us22_n534 ) , .A2( us22_n535 ) , .A1( us22_n536 ) , .ZN( us22_n620 ) );
  NOR4_X1 us22_U98 (.A4( us22_n524 ) , .A2( us22_n525 ) , .A1( us22_n526 ) , .ZN( us22_n536 ) , .A3( us22_n699 ) );
  NOR4_X1 us22_U99 (.A1( us22_n529 ) , .ZN( us22_n534 ) , .A2( us22_n652 ) , .A4( us22_n666 ) , .A3( us22_n763 ) );
endmodule
module aes_aes_die_1 ( sa00_0, sa00_1, sa00_2, sa00_3, sa00_4, sa00_5, sa00_6, sa00_7, sa03_0, 
       sa03_1, sa03_2, sa03_3, sa03_4, sa03_5, sa03_6, sa03_7, sa12_0, sa12_1, 
       sa12_2, sa12_3, sa12_4, sa12_5, sa12_6, sa12_7, sa31_0, sa31_1, sa31_2, 
       sa31_3, sa31_4, sa31_5, sa31_6, sa31_7, w3_0, w3_1, w3_2, w3_24, 
       w3_25, w3_26, w3_27, w3_28, w3_29, w3_3, w3_30, w3_31, w3_4, 
       w3_5, w3_6, w3_7, sa00_sr_0, sa00_sr_1, sa00_sr_2, sa00_sr_3, sa00_sr_4, sa00_sr_5, sa00_sr_6, sa00_sr_7, sa03_sr_0, 
        sa03_sr_1, sa03_sr_2, sa03_sr_3, sa03_sr_4, sa03_sr_5, sa03_sr_6, sa03_sr_7, sa11_sr_0, sa11_sr_1, 
        sa11_sr_2, sa11_sr_3, sa11_sr_4, sa11_sr_5, sa11_sr_6, sa11_sr_7, sa32_sr_0, sa32_sr_1, sa32_sr_2, 
        sa32_sr_3, sa32_sr_4, sa32_sr_5, sa32_sr_6, sa32_sr_7, u0_subword_0, u0_subword_1, u0_subword_10, u0_subword_11, 
        u0_subword_12, u0_subword_13, u0_subword_14, u0_subword_15, u0_subword_2, u0_subword_3, u0_subword_4, u0_subword_5, u0_subword_6, 
        u0_subword_7, u0_subword_8, u0_subword_9 );
  input sa00_0, sa00_1, sa00_2, sa00_3, sa00_4, sa00_5, sa00_6, sa00_7, sa03_0, 
        sa03_1, sa03_2, sa03_3, sa03_4, sa03_5, sa03_6, sa03_7, sa12_0, sa12_1, 
        sa12_2, sa12_3, sa12_4, sa12_5, sa12_6, sa12_7, sa31_0, sa31_1, sa31_2, 
        sa31_3, sa31_4, sa31_5, sa31_6, sa31_7, w3_0, w3_1, w3_2, w3_24, 
        w3_25, w3_26, w3_27, w3_28, w3_29, w3_3, w3_30, w3_31, w3_4, 
        w3_5, w3_6, w3_7;
  output sa00_sr_0, sa00_sr_1, sa00_sr_2, sa00_sr_3, sa00_sr_4, sa00_sr_5, sa00_sr_6, sa00_sr_7, sa03_sr_0, 
        sa03_sr_1, sa03_sr_2, sa03_sr_3, sa03_sr_4, sa03_sr_5, sa03_sr_6, sa03_sr_7, sa11_sr_0, sa11_sr_1, 
        sa11_sr_2, sa11_sr_3, sa11_sr_4, sa11_sr_5, sa11_sr_6, sa11_sr_7, sa32_sr_0, sa32_sr_1, sa32_sr_2, 
        sa32_sr_3, sa32_sr_4, sa32_sr_5, sa32_sr_6, sa32_sr_7, u0_subword_0, u0_subword_1, u0_subword_10, u0_subword_11, 
        u0_subword_12, u0_subword_13, u0_subword_14, u0_subword_15, u0_subword_2, u0_subword_3, u0_subword_4, u0_subword_5, u0_subword_6, 
        u0_subword_7, u0_subword_8, u0_subword_9;
  wire u0_u2_n438, u0_u2_n439, u0_u2_n440, u0_u2_n441, u0_u2_n442, u0_u2_n443, u0_u2_n444, u0_u2_n445, u0_u2_n446, 
       u0_u2_n447, u0_u2_n448, u0_u2_n449, u0_u2_n450, u0_u2_n451, u0_u2_n452, u0_u2_n453, u0_u2_n454, u0_u2_n455, 
       u0_u2_n456, u0_u2_n457, u0_u2_n458, u0_u2_n459, u0_u2_n460, u0_u2_n461, u0_u2_n462, u0_u2_n463, u0_u2_n464, 
       u0_u2_n465, u0_u2_n466, u0_u2_n467, u0_u2_n468, u0_u2_n469, u0_u2_n470, u0_u2_n471, u0_u2_n472, u0_u2_n473, 
       u0_u2_n474, u0_u2_n475, u0_u2_n476, u0_u2_n477, u0_u2_n478, u0_u2_n479, u0_u2_n480, u0_u2_n481, u0_u2_n482, 
       u0_u2_n483, u0_u2_n484, u0_u2_n485, u0_u2_n486, u0_u2_n487, u0_u2_n488, u0_u2_n489, u0_u2_n490, u0_u2_n491, 
       u0_u2_n492, u0_u2_n493, u0_u2_n494, u0_u2_n495, u0_u2_n496, u0_u2_n497, u0_u2_n498, u0_u2_n499, u0_u2_n500, 
       u0_u2_n501, u0_u2_n502, u0_u2_n503, u0_u2_n504, u0_u2_n505, u0_u2_n506, u0_u2_n507, u0_u2_n508, u0_u2_n509, 
       u0_u2_n510, u0_u2_n511, u0_u2_n512, u0_u2_n513, u0_u2_n514, u0_u2_n515, u0_u2_n516, u0_u2_n517, u0_u2_n518, 
       u0_u2_n519, u0_u2_n520, u0_u2_n521, u0_u2_n522, u0_u2_n523, u0_u2_n524, u0_u2_n525, u0_u2_n526, u0_u2_n527, 
       u0_u2_n528, u0_u2_n529, u0_u2_n530, u0_u2_n531, u0_u2_n532, u0_u2_n533, u0_u2_n534, u0_u2_n535, u0_u2_n536, 
       u0_u2_n537, u0_u2_n538, u0_u2_n539, u0_u2_n540, u0_u2_n541, u0_u2_n542, u0_u2_n543, u0_u2_n544, u0_u2_n545, 
       u0_u2_n546, u0_u2_n547, u0_u2_n548, u0_u2_n549, u0_u2_n550, u0_u2_n551, u0_u2_n552, u0_u2_n553, u0_u2_n554, 
       u0_u2_n555, u0_u2_n556, u0_u2_n557, u0_u2_n558, u0_u2_n559, u0_u2_n560, u0_u2_n561, u0_u2_n562, u0_u2_n563, 
       u0_u2_n564, u0_u2_n565, u0_u2_n566, u0_u2_n567, u0_u2_n568, u0_u2_n569, u0_u2_n570, u0_u2_n571, u0_u2_n572, 
       u0_u2_n573, u0_u2_n574, u0_u2_n575, u0_u2_n576, u0_u2_n577, u0_u2_n578, u0_u2_n579, u0_u2_n580, u0_u2_n581, 
       u0_u2_n582, u0_u2_n583, u0_u2_n584, u0_u2_n585, u0_u2_n586, u0_u2_n587, u0_u2_n588, u0_u2_n589, u0_u2_n590, 
       u0_u2_n591, u0_u2_n592, u0_u2_n593, u0_u2_n594, u0_u2_n595, u0_u2_n596, u0_u2_n597, u0_u2_n598, u0_u2_n599, 
       u0_u2_n600, u0_u2_n601, u0_u2_n602, u0_u2_n603, u0_u2_n604, u0_u2_n605, u0_u2_n606, u0_u2_n607, u0_u2_n608, 
       u0_u2_n609, u0_u2_n610, u0_u2_n611, u0_u2_n612, u0_u2_n613, u0_u2_n614, u0_u2_n615, u0_u2_n616, u0_u2_n617, 
       u0_u2_n618, u0_u2_n619, u0_u2_n620, u0_u2_n621, u0_u2_n622, u0_u2_n623, u0_u2_n624, u0_u2_n625, u0_u2_n626, 
       u0_u2_n627, u0_u2_n628, u0_u2_n629, u0_u2_n630, u0_u2_n631, u0_u2_n632, u0_u2_n633, u0_u2_n634, u0_u2_n635, 
       u0_u2_n636, u0_u2_n637, u0_u2_n638, u0_u2_n639, u0_u2_n640, u0_u2_n641, u0_u2_n642, u0_u2_n643, u0_u2_n644, 
       u0_u2_n645, u0_u2_n646, u0_u2_n647, u0_u2_n648, u0_u2_n649, u0_u2_n650, u0_u2_n651, u0_u2_n652, u0_u2_n653, 
       u0_u2_n654, u0_u2_n655, u0_u2_n656, u0_u2_n657, u0_u2_n658, u0_u2_n659, u0_u2_n660, u0_u2_n661, u0_u2_n662, 
       u0_u2_n663, u0_u2_n664, u0_u2_n665, u0_u2_n666, u0_u2_n667, u0_u2_n668, u0_u2_n669, u0_u2_n670, u0_u2_n671, 
       u0_u2_n672, u0_u2_n673, u0_u2_n674, u0_u2_n675, u0_u2_n676, u0_u2_n677, u0_u2_n678, u0_u2_n679, u0_u2_n680, 
       u0_u2_n681, u0_u2_n682, u0_u2_n683, u0_u2_n684, u0_u2_n685, u0_u2_n686, u0_u2_n687, u0_u2_n688, u0_u2_n689, 
       u0_u2_n690, u0_u2_n691, u0_u2_n692, u0_u2_n693, u0_u2_n694, u0_u2_n695, u0_u2_n696, u0_u2_n697, u0_u2_n698, 
       u0_u2_n699, u0_u2_n700, u0_u2_n701, u0_u2_n702, u0_u2_n703, u0_u2_n704, u0_u2_n705, u0_u2_n706, u0_u2_n707, 
       u0_u2_n708, u0_u2_n709, u0_u2_n710, u0_u2_n711, u0_u2_n712, u0_u2_n713, u0_u2_n714, u0_u2_n715, u0_u2_n716, 
       u0_u2_n717, u0_u2_n718, u0_u2_n719, u0_u2_n720, u0_u2_n721, u0_u2_n722, u0_u2_n723, u0_u2_n724, u0_u2_n725, 
       u0_u2_n726, u0_u2_n727, u0_u2_n728, u0_u2_n729, u0_u2_n730, u0_u2_n731, u0_u2_n732, u0_u2_n733, u0_u2_n734, 
       u0_u2_n735, u0_u2_n736, u0_u2_n737, u0_u2_n738, u0_u2_n739, u0_u2_n740, u0_u2_n741, u0_u2_n742, u0_u2_n743, 
       u0_u2_n744, u0_u2_n745, u0_u2_n746, u0_u2_n747, u0_u2_n748, u0_u2_n749, u0_u2_n750, u0_u2_n751, u0_u2_n752, 
       u0_u2_n753, u0_u2_n754, u0_u2_n755, u0_u2_n756, u0_u2_n757, u0_u2_n758, u0_u2_n759, u0_u2_n760, u0_u2_n761, 
       u0_u2_n762, u0_u2_n763, u0_u2_n764, u0_u2_n765, u0_u2_n766, u0_u2_n767, u0_u2_n768, u0_u2_n769, u0_u2_n770, 
       u0_u2_n771, u0_u2_n772, u0_u2_n773, u0_u2_n774, u0_u2_n775, u0_u2_n776, u0_u2_n777, u0_u2_n778, u0_u2_n779, 
       u0_u2_n780, u0_u2_n781, u0_u2_n782, u0_u2_n783, u0_u2_n784, u0_u2_n785, u0_u2_n786, u0_u2_n787, u0_u2_n788, 
       u0_u2_n789, u0_u2_n790, u0_u2_n791, u0_u2_n792, u0_u2_n793, u0_u2_n794, u0_u2_n795, u0_u2_n796, u0_u2_n797, 
       u0_u2_n798, u0_u2_n799, u0_u2_n800, u0_u2_n801, u0_u2_n802, u0_u2_n803, u0_u2_n804, u0_u2_n805, u0_u2_n806, 
       u0_u2_n807, u0_u2_n808, u0_u2_n809, u0_u2_n810, u0_u2_n811, u0_u2_n812, u0_u2_n813, u0_u2_n814, u0_u2_n815, 
       u0_u2_n816, u0_u2_n817, u0_u2_n818, u0_u2_n819, u0_u2_n820, u0_u2_n821, u0_u2_n822, u0_u2_n823, u0_u2_n824, 
       u0_u2_n825, u0_u2_n826, u0_u2_n827, u0_u2_n828, u0_u2_n829, u0_u2_n830, u0_u2_n831, u0_u2_n832, u0_u2_n833, 
       u0_u2_n834, u0_u2_n835, u0_u2_n836, u0_u2_n837, u0_u2_n838, u0_u2_n839, u0_u2_n840, u0_u2_n841, u0_u2_n842, 
       u0_u2_n843, u0_u2_n844, u0_u2_n845, u0_u2_n846, u0_u2_n847, u0_u2_n848, u0_u2_n849, u0_u2_n850, u0_u2_n851, 
       u0_u2_n852, u0_u2_n853, u0_u2_n854, u0_u2_n855, u0_u2_n856, u0_u2_n857, u0_u2_n858, u0_u2_n859, u0_u2_n860, 
       u0_u2_n861, u0_u2_n862, u0_u2_n863, u0_u2_n864, u0_u2_n865, u0_u2_n866, u0_u2_n867, u0_u2_n868, u0_u2_n869, 
       u0_u2_n870, u0_u2_n871, u0_u2_n872, u0_u2_n873, u0_u2_n874, u0_u2_n875, u0_u2_n876, u0_u2_n877, u0_u2_n878, 
       u0_u2_n879, u0_u2_n880, u0_u2_n881, u0_u2_n882, u0_u2_n883, u0_u3_n41, u0_u3_n438, u0_u3_n439, u0_u3_n440, 
       u0_u3_n441, u0_u3_n442, u0_u3_n443, u0_u3_n444, u0_u3_n445, u0_u3_n446, u0_u3_n447, u0_u3_n448, u0_u3_n449, 
       u0_u3_n450, u0_u3_n451, u0_u3_n452, u0_u3_n453, u0_u3_n454, u0_u3_n455, u0_u3_n456, u0_u3_n457, u0_u3_n458, 
       u0_u3_n459, u0_u3_n460, u0_u3_n461, u0_u3_n462, u0_u3_n463, u0_u3_n464, u0_u3_n465, u0_u3_n466, u0_u3_n467, 
       u0_u3_n468, u0_u3_n469, u0_u3_n470, u0_u3_n471, u0_u3_n472, u0_u3_n473, u0_u3_n474, u0_u3_n475, u0_u3_n476, 
       u0_u3_n477, u0_u3_n478, u0_u3_n479, u0_u3_n480, u0_u3_n481, u0_u3_n482, u0_u3_n483, u0_u3_n484, u0_u3_n485, 
       u0_u3_n486, u0_u3_n487, u0_u3_n488, u0_u3_n489, u0_u3_n490, u0_u3_n491, u0_u3_n492, u0_u3_n493, u0_u3_n494, 
       u0_u3_n495, u0_u3_n496, u0_u3_n497, u0_u3_n498, u0_u3_n499, u0_u3_n500, u0_u3_n501, u0_u3_n502, u0_u3_n503, 
       u0_u3_n504, u0_u3_n505, u0_u3_n506, u0_u3_n507, u0_u3_n508, u0_u3_n509, u0_u3_n510, u0_u3_n511, u0_u3_n512, 
       u0_u3_n513, u0_u3_n514, u0_u3_n515, u0_u3_n516, u0_u3_n517, u0_u3_n518, u0_u3_n519, u0_u3_n520, u0_u3_n521, 
       u0_u3_n522, u0_u3_n523, u0_u3_n524, u0_u3_n525, u0_u3_n526, u0_u3_n527, u0_u3_n528, u0_u3_n529, u0_u3_n530, 
       u0_u3_n531, u0_u3_n532, u0_u3_n533, u0_u3_n534, u0_u3_n535, u0_u3_n536, u0_u3_n537, u0_u3_n538, u0_u3_n539, 
       u0_u3_n540, u0_u3_n541, u0_u3_n542, u0_u3_n543, u0_u3_n544, u0_u3_n545, u0_u3_n546, u0_u3_n547, u0_u3_n548, 
       u0_u3_n549, u0_u3_n550, u0_u3_n551, u0_u3_n552, u0_u3_n553, u0_u3_n554, u0_u3_n555, u0_u3_n556, u0_u3_n557, 
       u0_u3_n558, u0_u3_n559, u0_u3_n560, u0_u3_n561, u0_u3_n562, u0_u3_n563, u0_u3_n564, u0_u3_n565, u0_u3_n566, 
       u0_u3_n567, u0_u3_n568, u0_u3_n569, u0_u3_n570, u0_u3_n571, u0_u3_n572, u0_u3_n573, u0_u3_n574, u0_u3_n575, 
       u0_u3_n576, u0_u3_n577, u0_u3_n578, u0_u3_n579, u0_u3_n580, u0_u3_n581, u0_u3_n582, u0_u3_n583, u0_u3_n584, 
       u0_u3_n585, u0_u3_n586, u0_u3_n587, u0_u3_n588, u0_u3_n589, u0_u3_n590, u0_u3_n591, u0_u3_n592, u0_u3_n593, 
       u0_u3_n594, u0_u3_n595, u0_u3_n596, u0_u3_n597, u0_u3_n598, u0_u3_n599, u0_u3_n600, u0_u3_n601, u0_u3_n602, 
       u0_u3_n603, u0_u3_n604, u0_u3_n605, u0_u3_n606, u0_u3_n607, u0_u3_n608, u0_u3_n609, u0_u3_n610, u0_u3_n611, 
       u0_u3_n612, u0_u3_n613, u0_u3_n614, u0_u3_n615, u0_u3_n616, u0_u3_n617, u0_u3_n618, u0_u3_n619, u0_u3_n620, 
       u0_u3_n621, u0_u3_n622, u0_u3_n623, u0_u3_n624, u0_u3_n625, u0_u3_n626, u0_u3_n627, u0_u3_n628, u0_u3_n629, 
       u0_u3_n630, u0_u3_n631, u0_u3_n632, u0_u3_n633, u0_u3_n634, u0_u3_n635, u0_u3_n636, u0_u3_n637, u0_u3_n638, 
       u0_u3_n639, u0_u3_n640, u0_u3_n641, u0_u3_n642, u0_u3_n643, u0_u3_n644, u0_u3_n645, u0_u3_n646, u0_u3_n647, 
       u0_u3_n648, u0_u3_n649, u0_u3_n650, u0_u3_n651, u0_u3_n652, u0_u3_n653, u0_u3_n654, u0_u3_n655, u0_u3_n656, 
       u0_u3_n657, u0_u3_n658, u0_u3_n659, u0_u3_n660, u0_u3_n661, u0_u3_n662, u0_u3_n663, u0_u3_n664, u0_u3_n665, 
       u0_u3_n666, u0_u3_n667, u0_u3_n668, u0_u3_n669, u0_u3_n670, u0_u3_n671, u0_u3_n672, u0_u3_n673, u0_u3_n674, 
       u0_u3_n675, u0_u3_n676, u0_u3_n677, u0_u3_n678, u0_u3_n679, u0_u3_n680, u0_u3_n681, u0_u3_n682, u0_u3_n683, 
       u0_u3_n684, u0_u3_n685, u0_u3_n686, u0_u3_n687, u0_u3_n688, u0_u3_n689, u0_u3_n690, u0_u3_n691, u0_u3_n692, 
       u0_u3_n693, u0_u3_n694, u0_u3_n695, u0_u3_n696, u0_u3_n697, u0_u3_n698, u0_u3_n699, u0_u3_n700, u0_u3_n701, 
       u0_u3_n702, u0_u3_n703, u0_u3_n704, u0_u3_n705, u0_u3_n706, u0_u3_n707, u0_u3_n708, u0_u3_n709, u0_u3_n710, 
       u0_u3_n711, u0_u3_n712, u0_u3_n713, u0_u3_n714, u0_u3_n715, u0_u3_n716, u0_u3_n717, u0_u3_n718, u0_u3_n719, 
       u0_u3_n720, u0_u3_n721, u0_u3_n722, u0_u3_n723, u0_u3_n724, u0_u3_n725, u0_u3_n726, u0_u3_n727, u0_u3_n728, 
       u0_u3_n729, u0_u3_n730, u0_u3_n731, u0_u3_n732, u0_u3_n733, u0_u3_n734, u0_u3_n735, u0_u3_n736, u0_u3_n737, 
       u0_u3_n738, u0_u3_n739, u0_u3_n740, u0_u3_n741, u0_u3_n742, u0_u3_n743, u0_u3_n744, u0_u3_n745, u0_u3_n746, 
       u0_u3_n747, u0_u3_n748, u0_u3_n749, u0_u3_n750, u0_u3_n751, u0_u3_n752, u0_u3_n753, u0_u3_n754, u0_u3_n755, 
       u0_u3_n756, u0_u3_n757, u0_u3_n758, u0_u3_n759, u0_u3_n760, u0_u3_n761, u0_u3_n762, u0_u3_n763, u0_u3_n764, 
       u0_u3_n765, u0_u3_n766, u0_u3_n767, u0_u3_n768, u0_u3_n769, u0_u3_n770, u0_u3_n771, u0_u3_n772, u0_u3_n773, 
       u0_u3_n774, u0_u3_n775, u0_u3_n776, u0_u3_n777, u0_u3_n778, u0_u3_n779, u0_u3_n780, u0_u3_n781, u0_u3_n782, 
       u0_u3_n783, u0_u3_n784, u0_u3_n785, u0_u3_n786, u0_u3_n787, u0_u3_n788, u0_u3_n789, u0_u3_n790, u0_u3_n791, 
       u0_u3_n792, u0_u3_n793, u0_u3_n794, u0_u3_n795, u0_u3_n796, u0_u3_n797, u0_u3_n798, u0_u3_n799, u0_u3_n800, 
       u0_u3_n801, u0_u3_n802, u0_u3_n803, u0_u3_n804, u0_u3_n805, u0_u3_n806, u0_u3_n807, u0_u3_n808, u0_u3_n809, 
       u0_u3_n810, u0_u3_n811, u0_u3_n812, u0_u3_n813, u0_u3_n814, u0_u3_n815, u0_u3_n816, u0_u3_n817, u0_u3_n818, 
       u0_u3_n819, u0_u3_n820, u0_u3_n821, u0_u3_n822, u0_u3_n823, u0_u3_n824, u0_u3_n825, u0_u3_n826, u0_u3_n827, 
       u0_u3_n828, u0_u3_n829, u0_u3_n830, u0_u3_n831, u0_u3_n832, u0_u3_n833, u0_u3_n834, u0_u3_n835, u0_u3_n836, 
       u0_u3_n837, u0_u3_n838, u0_u3_n839, u0_u3_n840, u0_u3_n841, u0_u3_n842, u0_u3_n843, u0_u3_n844, u0_u3_n845, 
       u0_u3_n846, u0_u3_n847, u0_u3_n848, u0_u3_n849, u0_u3_n850, u0_u3_n851, u0_u3_n852, u0_u3_n853, u0_u3_n854, 
       u0_u3_n855, u0_u3_n856, u0_u3_n857, u0_u3_n858, u0_u3_n859, u0_u3_n860, u0_u3_n861, u0_u3_n862, u0_u3_n863, 
       u0_u3_n864, u0_u3_n865, u0_u3_n866, u0_u3_n867, u0_u3_n868, u0_u3_n869, u0_u3_n870, u0_u3_n871, u0_u3_n872, 
       u0_u3_n873, u0_u3_n874, u0_u3_n875, u0_u3_n876, u0_u3_n877, u0_u3_n878, us00_n1, us00_n10, us00_n100, 
       us00_n101, us00_n102, us00_n103, us00_n104, us00_n105, us00_n106, us00_n107, us00_n108, us00_n109, 
       us00_n11, us00_n110, us00_n111, us00_n112, us00_n113, us00_n114, us00_n115, us00_n116, us00_n117, 
       us00_n118, us00_n119, us00_n12, us00_n120, us00_n121, us00_n122, us00_n123, us00_n124, us00_n125, 
       us00_n126, us00_n127, us00_n128, us00_n129, us00_n13, us00_n130, us00_n131, us00_n132, us00_n133, 
       us00_n134, us00_n135, us00_n136, us00_n137, us00_n138, us00_n139, us00_n14, us00_n140, us00_n141, 
       us00_n142, us00_n143, us00_n144, us00_n145, us00_n146, us00_n147, us00_n148, us00_n149, us00_n15, 
       us00_n150, us00_n151, us00_n152, us00_n153, us00_n154, us00_n155, us00_n156, us00_n157, us00_n158, 
       us00_n159, us00_n16, us00_n160, us00_n161, us00_n162, us00_n163, us00_n164, us00_n165, us00_n166, 
       us00_n167, us00_n168, us00_n169, us00_n17, us00_n170, us00_n171, us00_n172, us00_n173, us00_n174, 
       us00_n175, us00_n176, us00_n177, us00_n178, us00_n179, us00_n18, us00_n180, us00_n181, us00_n182, 
       us00_n183, us00_n184, us00_n185, us00_n186, us00_n187, us00_n188, us00_n189, us00_n19, us00_n190, 
       us00_n191, us00_n192, us00_n193, us00_n194, us00_n195, us00_n196, us00_n197, us00_n198, us00_n199, 
       us00_n2, us00_n20, us00_n200, us00_n201, us00_n202, us00_n203, us00_n204, us00_n205, us00_n206, 
       us00_n207, us00_n208, us00_n209, us00_n21, us00_n210, us00_n211, us00_n212, us00_n213, us00_n214, 
       us00_n215, us00_n216, us00_n217, us00_n218, us00_n219, us00_n22, us00_n220, us00_n221, us00_n222, 
       us00_n223, us00_n224, us00_n225, us00_n226, us00_n227, us00_n228, us00_n229, us00_n23, us00_n230, 
       us00_n231, us00_n232, us00_n233, us00_n234, us00_n235, us00_n236, us00_n237, us00_n238, us00_n239, 
       us00_n24, us00_n240, us00_n241, us00_n242, us00_n243, us00_n244, us00_n245, us00_n246, us00_n247, 
       us00_n248, us00_n249, us00_n25, us00_n250, us00_n251, us00_n252, us00_n253, us00_n254, us00_n255, 
       us00_n256, us00_n257, us00_n258, us00_n259, us00_n26, us00_n260, us00_n261, us00_n262, us00_n263, 
       us00_n264, us00_n265, us00_n266, us00_n267, us00_n268, us00_n269, us00_n27, us00_n270, us00_n271, 
       us00_n272, us00_n273, us00_n274, us00_n275, us00_n276, us00_n277, us00_n278, us00_n279, us00_n28, 
       us00_n280, us00_n281, us00_n282, us00_n283, us00_n284, us00_n285, us00_n286, us00_n287, us00_n288, 
       us00_n289, us00_n29, us00_n290, us00_n291, us00_n292, us00_n293, us00_n294, us00_n295, us00_n296, 
       us00_n297, us00_n298, us00_n299, us00_n3, us00_n30, us00_n300, us00_n301, us00_n302, us00_n303, 
       us00_n304, us00_n305, us00_n306, us00_n307, us00_n308, us00_n309, us00_n31, us00_n310, us00_n311, 
       us00_n312, us00_n313, us00_n314, us00_n315, us00_n316, us00_n317, us00_n318, us00_n319, us00_n32, 
       us00_n320, us00_n321, us00_n322, us00_n323, us00_n324, us00_n325, us00_n326, us00_n327, us00_n328, 
       us00_n329, us00_n33, us00_n330, us00_n331, us00_n332, us00_n333, us00_n334, us00_n335, us00_n336, 
       us00_n337, us00_n338, us00_n339, us00_n34, us00_n340, us00_n341, us00_n342, us00_n343, us00_n344, 
       us00_n345, us00_n346, us00_n347, us00_n348, us00_n349, us00_n35, us00_n350, us00_n351, us00_n352, 
       us00_n353, us00_n354, us00_n355, us00_n356, us00_n357, us00_n358, us00_n359, us00_n36, us00_n360, 
       us00_n361, us00_n362, us00_n363, us00_n364, us00_n365, us00_n366, us00_n367, us00_n368, us00_n369, 
       us00_n37, us00_n370, us00_n371, us00_n372, us00_n373, us00_n374, us00_n375, us00_n376, us00_n377, 
       us00_n378, us00_n379, us00_n38, us00_n380, us00_n381, us00_n382, us00_n383, us00_n384, us00_n385, 
       us00_n386, us00_n387, us00_n388, us00_n389, us00_n39, us00_n390, us00_n391, us00_n392, us00_n393, 
       us00_n394, us00_n395, us00_n396, us00_n397, us00_n398, us00_n399, us00_n4, us00_n40, us00_n400, 
       us00_n401, us00_n402, us00_n403, us00_n404, us00_n405, us00_n406, us00_n407, us00_n408, us00_n409, 
       us00_n41, us00_n410, us00_n411, us00_n412, us00_n413, us00_n414, us00_n415, us00_n416, us00_n417, 
       us00_n418, us00_n419, us00_n42, us00_n420, us00_n421, us00_n422, us00_n423, us00_n424, us00_n425, 
       us00_n426, us00_n427, us00_n428, us00_n429, us00_n43, us00_n430, us00_n431, us00_n432, us00_n433, 
       us00_n434, us00_n435, us00_n436, us00_n437, us00_n44, us00_n45, us00_n46, us00_n47, us00_n48, 
       us00_n49, us00_n5, us00_n50, us00_n51, us00_n52, us00_n53, us00_n54, us00_n55, us00_n56, 
       us00_n57, us00_n58, us00_n59, us00_n6, us00_n60, us00_n61, us00_n62, us00_n63, us00_n64, 
       us00_n65, us00_n66, us00_n67, us00_n68, us00_n69, us00_n7, us00_n70, us00_n71, us00_n72, 
       us00_n73, us00_n74, us00_n75, us00_n76, us00_n77, us00_n78, us00_n79, us00_n8, us00_n80, 
       us00_n81, us00_n82, us00_n83, us00_n84, us00_n85, us00_n86, us00_n87, us00_n88, us00_n89, 
       us00_n9, us00_n90, us00_n91, us00_n92, us00_n93, us00_n94, us00_n95, us00_n96, us00_n97, 
       us00_n98, us00_n99, us03_n438, us03_n439, us03_n440, us03_n441, us03_n442, us03_n443, us03_n444, 
       us03_n445, us03_n446, us03_n447, us03_n448, us03_n449, us03_n450, us03_n451, us03_n452, us03_n453, 
       us03_n454, us03_n455, us03_n456, us03_n457, us03_n458, us03_n459, us03_n460, us03_n461, us03_n462, 
       us03_n463, us03_n464, us03_n465, us03_n466, us03_n467, us03_n468, us03_n469, us03_n470, us03_n471, 
       us03_n472, us03_n473, us03_n474, us03_n475, us03_n476, us03_n477, us03_n478, us03_n479, us03_n480, 
       us03_n481, us03_n482, us03_n483, us03_n484, us03_n485, us03_n486, us03_n487, us03_n488, us03_n489, 
       us03_n490, us03_n491, us03_n492, us03_n493, us03_n494, us03_n495, us03_n496, us03_n497, us03_n498, 
       us03_n499, us03_n500, us03_n501, us03_n502, us03_n503, us03_n504, us03_n505, us03_n506, us03_n507, 
       us03_n508, us03_n509, us03_n510, us03_n511, us03_n512, us03_n513, us03_n514, us03_n515, us03_n516, 
       us03_n517, us03_n518, us03_n519, us03_n520, us03_n521, us03_n522, us03_n523, us03_n524, us03_n525, 
       us03_n526, us03_n527, us03_n528, us03_n529, us03_n530, us03_n531, us03_n532, us03_n533, us03_n534, 
       us03_n535, us03_n536, us03_n537, us03_n538, us03_n539, us03_n540, us03_n541, us03_n542, us03_n543, 
       us03_n544, us03_n545, us03_n546, us03_n547, us03_n548, us03_n549, us03_n550, us03_n551, us03_n552, 
       us03_n553, us03_n554, us03_n555, us03_n556, us03_n557, us03_n558, us03_n559, us03_n560, us03_n561, 
       us03_n562, us03_n563, us03_n564, us03_n565, us03_n566, us03_n567, us03_n568, us03_n569, us03_n570, 
       us03_n571, us03_n572, us03_n573, us03_n574, us03_n575, us03_n576, us03_n577, us03_n578, us03_n579, 
       us03_n580, us03_n581, us03_n582, us03_n583, us03_n584, us03_n585, us03_n586, us03_n587, us03_n588, 
       us03_n589, us03_n590, us03_n591, us03_n592, us03_n593, us03_n594, us03_n595, us03_n596, us03_n597, 
       us03_n598, us03_n599, us03_n600, us03_n601, us03_n602, us03_n603, us03_n604, us03_n605, us03_n606, 
       us03_n607, us03_n608, us03_n609, us03_n610, us03_n611, us03_n612, us03_n613, us03_n614, us03_n615, 
       us03_n616, us03_n617, us03_n618, us03_n619, us03_n620, us03_n621, us03_n622, us03_n623, us03_n624, 
       us03_n625, us03_n626, us03_n627, us03_n628, us03_n629, us03_n630, us03_n631, us03_n632, us03_n633, 
       us03_n634, us03_n635, us03_n636, us03_n637, us03_n638, us03_n639, us03_n640, us03_n641, us03_n642, 
       us03_n643, us03_n644, us03_n645, us03_n646, us03_n647, us03_n648, us03_n649, us03_n650, us03_n651, 
       us03_n652, us03_n653, us03_n654, us03_n655, us03_n656, us03_n657, us03_n658, us03_n659, us03_n660, 
       us03_n661, us03_n662, us03_n663, us03_n664, us03_n665, us03_n666, us03_n667, us03_n668, us03_n669, 
       us03_n670, us03_n671, us03_n672, us03_n673, us03_n674, us03_n675, us03_n676, us03_n677, us03_n678, 
       us03_n679, us03_n680, us03_n681, us03_n682, us03_n683, us03_n684, us03_n685, us03_n686, us03_n687, 
       us03_n688, us03_n689, us03_n690, us03_n691, us03_n692, us03_n693, us03_n694, us03_n695, us03_n696, 
       us03_n697, us03_n698, us03_n699, us03_n700, us03_n701, us03_n702, us03_n703, us03_n704, us03_n705, 
       us03_n706, us03_n707, us03_n708, us03_n709, us03_n710, us03_n711, us03_n712, us03_n713, us03_n714, 
       us03_n715, us03_n716, us03_n717, us03_n718, us03_n719, us03_n720, us03_n721, us03_n722, us03_n723, 
       us03_n724, us03_n725, us03_n726, us03_n727, us03_n728, us03_n729, us03_n730, us03_n731, us03_n732, 
       us03_n733, us03_n734, us03_n735, us03_n736, us03_n737, us03_n738, us03_n739, us03_n740, us03_n741, 
       us03_n742, us03_n743, us03_n744, us03_n745, us03_n746, us03_n747, us03_n748, us03_n749, us03_n750, 
       us03_n751, us03_n752, us03_n753, us03_n754, us03_n755, us03_n756, us03_n757, us03_n758, us03_n759, 
       us03_n760, us03_n761, us03_n762, us03_n763, us03_n764, us03_n765, us03_n766, us03_n767, us03_n768, 
       us03_n769, us03_n770, us03_n771, us03_n772, us03_n773, us03_n774, us03_n775, us03_n776, us03_n777, 
       us03_n778, us03_n779, us03_n780, us03_n781, us03_n782, us03_n783, us03_n784, us03_n785, us03_n786, 
       us03_n787, us03_n788, us03_n789, us03_n790, us03_n791, us03_n792, us03_n793, us03_n794, us03_n795, 
       us03_n796, us03_n797, us03_n798, us03_n799, us03_n800, us03_n801, us03_n802, us03_n803, us03_n804, 
       us03_n805, us03_n806, us03_n807, us03_n808, us03_n809, us03_n810, us03_n811, us03_n812, us03_n813, 
       us03_n814, us03_n815, us03_n816, us03_n817, us03_n818, us03_n819, us03_n820, us03_n821, us03_n822, 
       us03_n823, us03_n824, us03_n825, us03_n826, us03_n827, us03_n828, us03_n829, us03_n830, us03_n831, 
       us03_n832, us03_n833, us03_n834, us03_n835, us03_n836, us03_n837, us03_n838, us03_n839, us03_n840, 
       us03_n841, us03_n842, us03_n843, us03_n844, us03_n845, us03_n846, us03_n847, us03_n848, us03_n849, 
       us03_n850, us03_n851, us03_n852, us03_n853, us03_n854, us03_n855, us03_n856, us03_n857, us03_n858, 
       us03_n859, us03_n860, us03_n861, us03_n862, us03_n863, us03_n864, us03_n865, us03_n866, us03_n867, 
       us03_n868, us03_n869, us03_n870, us03_n871, us03_n872, us03_n873, us03_n874, us12_n438, us12_n439, 
       us12_n440, us12_n441, us12_n442, us12_n443, us12_n444, us12_n445, us12_n446, us12_n447, us12_n448, 
       us12_n449, us12_n450, us12_n451, us12_n452, us12_n453, us12_n454, us12_n455, us12_n456, us12_n457, 
       us12_n458, us12_n459, us12_n460, us12_n461, us12_n462, us12_n463, us12_n464, us12_n465, us12_n466, 
       us12_n467, us12_n468, us12_n469, us12_n470, us12_n471, us12_n472, us12_n473, us12_n474, us12_n475, 
       us12_n476, us12_n477, us12_n478, us12_n479, us12_n480, us12_n481, us12_n482, us12_n483, us12_n484, 
       us12_n485, us12_n486, us12_n487, us12_n488, us12_n489, us12_n490, us12_n491, us12_n492, us12_n493, 
       us12_n494, us12_n495, us12_n496, us12_n497, us12_n498, us12_n499, us12_n500, us12_n501, us12_n502, 
       us12_n503, us12_n504, us12_n505, us12_n506, us12_n507, us12_n508, us12_n509, us12_n510, us12_n511, 
       us12_n512, us12_n513, us12_n514, us12_n515, us12_n516, us12_n517, us12_n518, us12_n519, us12_n520, 
       us12_n521, us12_n522, us12_n523, us12_n524, us12_n525, us12_n526, us12_n527, us12_n528, us12_n529, 
       us12_n530, us12_n531, us12_n532, us12_n533, us12_n534, us12_n535, us12_n536, us12_n537, us12_n538, 
       us12_n539, us12_n540, us12_n541, us12_n542, us12_n543, us12_n544, us12_n545, us12_n546, us12_n547, 
       us12_n548, us12_n549, us12_n550, us12_n551, us12_n552, us12_n553, us12_n554, us12_n555, us12_n556, 
       us12_n557, us12_n558, us12_n559, us12_n560, us12_n561, us12_n562, us12_n563, us12_n564, us12_n565, 
       us12_n566, us12_n567, us12_n568, us12_n569, us12_n570, us12_n571, us12_n572, us12_n573, us12_n574, 
       us12_n575, us12_n576, us12_n577, us12_n578, us12_n579, us12_n580, us12_n581, us12_n582, us12_n583, 
       us12_n584, us12_n585, us12_n586, us12_n587, us12_n588, us12_n589, us12_n590, us12_n591, us12_n592, 
       us12_n593, us12_n594, us12_n595, us12_n596, us12_n597, us12_n598, us12_n599, us12_n600, us12_n601, 
       us12_n602, us12_n603, us12_n604, us12_n605, us12_n606, us12_n607, us12_n608, us12_n609, us12_n610, 
       us12_n611, us12_n612, us12_n613, us12_n614, us12_n615, us12_n616, us12_n617, us12_n618, us12_n619, 
       us12_n620, us12_n621, us12_n622, us12_n623, us12_n624, us12_n625, us12_n626, us12_n627, us12_n628, 
       us12_n629, us12_n630, us12_n631, us12_n632, us12_n633, us12_n634, us12_n635, us12_n636, us12_n637, 
       us12_n638, us12_n639, us12_n640, us12_n641, us12_n642, us12_n643, us12_n644, us12_n645, us12_n646, 
       us12_n647, us12_n648, us12_n649, us12_n650, us12_n651, us12_n652, us12_n653, us12_n654, us12_n655, 
       us12_n656, us12_n657, us12_n658, us12_n659, us12_n660, us12_n661, us12_n662, us12_n663, us12_n664, 
       us12_n665, us12_n666, us12_n667, us12_n668, us12_n669, us12_n670, us12_n671, us12_n672, us12_n673, 
       us12_n674, us12_n675, us12_n676, us12_n677, us12_n678, us12_n679, us12_n680, us12_n681, us12_n682, 
       us12_n683, us12_n684, us12_n685, us12_n686, us12_n687, us12_n688, us12_n689, us12_n690, us12_n691, 
       us12_n692, us12_n693, us12_n694, us12_n695, us12_n696, us12_n697, us12_n698, us12_n699, us12_n700, 
       us12_n701, us12_n702, us12_n703, us12_n704, us12_n705, us12_n706, us12_n707, us12_n708, us12_n709, 
       us12_n710, us12_n711, us12_n712, us12_n713, us12_n714, us12_n715, us12_n716, us12_n717, us12_n718, 
       us12_n719, us12_n720, us12_n721, us12_n722, us12_n723, us12_n724, us12_n725, us12_n726, us12_n727, 
       us12_n728, us12_n729, us12_n730, us12_n731, us12_n732, us12_n733, us12_n734, us12_n735, us12_n736, 
       us12_n737, us12_n738, us12_n739, us12_n740, us12_n741, us12_n742, us12_n743, us12_n744, us12_n745, 
       us12_n746, us12_n747, us12_n748, us12_n749, us12_n750, us12_n751, us12_n752, us12_n753, us12_n754, 
       us12_n755, us12_n756, us12_n757, us12_n758, us12_n759, us12_n760, us12_n761, us12_n762, us12_n763, 
       us12_n764, us12_n765, us12_n766, us12_n767, us12_n768, us12_n769, us12_n770, us12_n771, us12_n772, 
       us12_n773, us12_n774, us12_n775, us12_n776, us12_n777, us12_n778, us12_n779, us12_n780, us12_n781, 
       us12_n782, us12_n783, us12_n784, us12_n785, us12_n786, us12_n787, us12_n788, us12_n789, us12_n790, 
       us12_n791, us12_n792, us12_n793, us12_n794, us12_n795, us12_n796, us12_n797, us12_n798, us12_n799, 
       us12_n800, us12_n801, us12_n802, us12_n803, us12_n804, us12_n805, us12_n806, us12_n807, us12_n808, 
       us12_n809, us12_n810, us12_n811, us12_n812, us12_n813, us12_n814, us12_n815, us12_n816, us12_n817, 
       us12_n818, us12_n819, us12_n820, us12_n821, us12_n822, us12_n823, us12_n824, us12_n825, us12_n826, 
       us12_n827, us12_n828, us12_n829, us12_n830, us12_n831, us12_n832, us12_n833, us12_n834, us12_n835, 
       us12_n836, us12_n837, us12_n838, us12_n839, us12_n840, us12_n841, us12_n842, us12_n843, us12_n844, 
       us12_n845, us12_n846, us12_n847, us12_n848, us12_n849, us12_n850, us12_n851, us12_n852, us12_n853, 
       us12_n854, us12_n855, us12_n856, us12_n857, us12_n858, us12_n859, us12_n860, us12_n861, us12_n862, 
       us12_n863, us12_n864, us12_n865, us12_n866, us12_n867, us12_n868, us12_n869, us12_n870, us12_n871, 
       us12_n872, us12_n873, us12_n874, us12_n875, us12_n876, us31_n438, us31_n439, us31_n440, us31_n441, 
       us31_n442, us31_n443, us31_n444, us31_n445, us31_n446, us31_n447, us31_n448, us31_n449, us31_n450, 
       us31_n451, us31_n452, us31_n453, us31_n454, us31_n455, us31_n456, us31_n457, us31_n458, us31_n459, 
       us31_n460, us31_n461, us31_n462, us31_n463, us31_n464, us31_n465, us31_n466, us31_n467, us31_n468, 
       us31_n469, us31_n470, us31_n471, us31_n472, us31_n473, us31_n474, us31_n475, us31_n476, us31_n477, 
       us31_n478, us31_n479, us31_n480, us31_n481, us31_n482, us31_n483, us31_n484, us31_n485, us31_n486, 
       us31_n487, us31_n488, us31_n489, us31_n490, us31_n491, us31_n492, us31_n493, us31_n494, us31_n495, 
       us31_n496, us31_n497, us31_n498, us31_n499, us31_n500, us31_n501, us31_n502, us31_n503, us31_n504, 
       us31_n505, us31_n506, us31_n507, us31_n508, us31_n509, us31_n510, us31_n511, us31_n512, us31_n513, 
       us31_n514, us31_n515, us31_n516, us31_n517, us31_n518, us31_n519, us31_n520, us31_n521, us31_n522, 
       us31_n523, us31_n524, us31_n525, us31_n526, us31_n527, us31_n528, us31_n529, us31_n530, us31_n531, 
       us31_n532, us31_n533, us31_n534, us31_n535, us31_n536, us31_n537, us31_n538, us31_n539, us31_n540, 
       us31_n541, us31_n542, us31_n543, us31_n544, us31_n545, us31_n546, us31_n547, us31_n548, us31_n549, 
       us31_n550, us31_n551, us31_n552, us31_n553, us31_n554, us31_n555, us31_n556, us31_n557, us31_n558, 
       us31_n559, us31_n560, us31_n561, us31_n562, us31_n563, us31_n564, us31_n565, us31_n566, us31_n567, 
       us31_n568, us31_n569, us31_n570, us31_n571, us31_n572, us31_n573, us31_n574, us31_n575, us31_n576, 
       us31_n577, us31_n578, us31_n579, us31_n580, us31_n581, us31_n582, us31_n583, us31_n584, us31_n585, 
       us31_n586, us31_n587, us31_n588, us31_n589, us31_n590, us31_n591, us31_n592, us31_n593, us31_n594, 
       us31_n595, us31_n596, us31_n597, us31_n598, us31_n599, us31_n600, us31_n601, us31_n602, us31_n603, 
       us31_n604, us31_n605, us31_n606, us31_n607, us31_n608, us31_n609, us31_n610, us31_n611, us31_n612, 
       us31_n613, us31_n614, us31_n615, us31_n616, us31_n617, us31_n618, us31_n619, us31_n620, us31_n621, 
       us31_n622, us31_n623, us31_n624, us31_n625, us31_n626, us31_n627, us31_n628, us31_n629, us31_n630, 
       us31_n631, us31_n632, us31_n633, us31_n634, us31_n635, us31_n636, us31_n637, us31_n638, us31_n639, 
       us31_n640, us31_n641, us31_n642, us31_n643, us31_n644, us31_n645, us31_n646, us31_n647, us31_n648, 
       us31_n649, us31_n650, us31_n651, us31_n652, us31_n653, us31_n654, us31_n655, us31_n656, us31_n657, 
       us31_n658, us31_n659, us31_n660, us31_n661, us31_n662, us31_n663, us31_n664, us31_n665, us31_n666, 
       us31_n667, us31_n668, us31_n669, us31_n670, us31_n671, us31_n672, us31_n673, us31_n674, us31_n675, 
       us31_n676, us31_n677, us31_n678, us31_n679, us31_n680, us31_n681, us31_n682, us31_n683, us31_n684, 
       us31_n685, us31_n686, us31_n687, us31_n688, us31_n689, us31_n690, us31_n691, us31_n692, us31_n693, 
       us31_n694, us31_n695, us31_n696, us31_n697, us31_n698, us31_n699, us31_n700, us31_n701, us31_n702, 
       us31_n703, us31_n704, us31_n705, us31_n706, us31_n707, us31_n708, us31_n709, us31_n710, us31_n711, 
       us31_n712, us31_n713, us31_n714, us31_n715, us31_n716, us31_n717, us31_n718, us31_n719, us31_n720, 
       us31_n721, us31_n722, us31_n723, us31_n724, us31_n725, us31_n726, us31_n727, us31_n728, us31_n729, 
       us31_n730, us31_n731, us31_n732, us31_n733, us31_n734, us31_n735, us31_n736, us31_n737, us31_n738, 
       us31_n739, us31_n740, us31_n741, us31_n742, us31_n743, us31_n744, us31_n745, us31_n746, us31_n747, 
       us31_n748, us31_n749, us31_n750, us31_n751, us31_n752, us31_n753, us31_n754, us31_n755, us31_n756, 
       us31_n757, us31_n758, us31_n759, us31_n760, us31_n761, us31_n762, us31_n763, us31_n764, us31_n765, 
       us31_n766, us31_n767, us31_n768, us31_n769, us31_n770, us31_n771, us31_n772, us31_n773, us31_n774, 
       us31_n775, us31_n776, us31_n777, us31_n778, us31_n779, us31_n780, us31_n781, us31_n782, us31_n783, 
       us31_n784, us31_n785, us31_n786, us31_n787, us31_n788, us31_n789, us31_n790, us31_n791, us31_n792, 
       us31_n793, us31_n794, us31_n795, us31_n796, us31_n797, us31_n798, us31_n799, us31_n800, us31_n801, 
       us31_n802, us31_n803, us31_n804, us31_n805, us31_n806, us31_n807, us31_n808, us31_n809, us31_n810, 
       us31_n811, us31_n812, us31_n813, us31_n814, us31_n815, us31_n816, us31_n817, us31_n818, us31_n819, 
       us31_n820, us31_n821, us31_n822, us31_n823, us31_n824, us31_n825, us31_n826, us31_n827, us31_n828, 
       us31_n829, us31_n830, us31_n831, us31_n832, us31_n833, us31_n834, us31_n835, us31_n836, us31_n837, 
       us31_n838, us31_n839, us31_n840, us31_n841, us31_n842, us31_n843, us31_n844, us31_n845, us31_n846, 
       us31_n847, us31_n848, us31_n849, us31_n850, us31_n851, us31_n852, us31_n853, us31_n854, us31_n855, 
       us31_n856, us31_n857, us31_n858, us31_n859, us31_n860, us31_n861, us31_n862, us31_n863, us31_n864, 
       us31_n865, us31_n866, us31_n867, us31_n868, us31_n869, us31_n870, us31_n871, us31_n872, us31_n873, 
       us31_n874, us31_n875,  us31_n876;
  NOR2_X1 u0_u2_U10 (.ZN( u0_u2_n714 ) , .A2( u0_u2_n783 ) , .A1( u0_u2_n807 ) );
  OR4_X1 u0_u2_U100 (.ZN( u0_u2_n473 ) , .A4( u0_u2_n525 ) , .A3( u0_u2_n536 ) , .A2( u0_u2_n585 ) , .A1( u0_u2_n719 ) );
  NOR4_X1 u0_u2_U101 (.A4( u0_u2_n584 ) , .A3( u0_u2_n585 ) , .A2( u0_u2_n586 ) , .ZN( u0_u2_n593 ) , .A1( u0_u2_n690 ) );
  NOR4_X1 u0_u2_U102 (.A1( u0_u2_n591 ) , .ZN( u0_u2_n592 ) , .A3( u0_u2_n659 ) , .A2( u0_u2_n669 ) , .A4( u0_u2_n774 ) );
  OR4_X1 u0_u2_U103 (.ZN( u0_u2_n499 ) , .A4( u0_u2_n541 ) , .A2( u0_u2_n554 ) , .A1( u0_u2_n566 ) , .A3( u0_u2_n639 ) );
  OR3_X1 u0_u2_U104 (.A3( u0_u2_n513 ) , .A2( u0_u2_n514 ) , .A1( u0_u2_n515 ) , .ZN( u0_u2_n518 ) );
  AOI21_X1 u0_u2_U105 (.A( u0_u2_n677 ) , .B1( u0_u2_n678 ) , .ZN( u0_u2_n679 ) , .B2( u0_u2_n863 ) );
  INV_X1 u0_u2_U106 (.A( u0_u2_n761 ) , .ZN( u0_u2_n876 ) );
  OAI21_X1 u0_u2_U107 (.B1( u0_u2_n760 ) , .ZN( u0_u2_n761 ) , .A( u0_u2_n852 ) , .B2( u0_u2_n875 ) );
  AOI221_X1 u0_u2_U108 (.A( u0_u2_n720 ) , .B2( u0_u2_n721 ) , .ZN( u0_u2_n727 ) , .C1( u0_u2_n839 ) , .B1( u0_u2_n846 ) , .C2( u0_u2_n870 ) );
  OR2_X1 u0_u2_U109 (.A2( u0_u2_n718 ) , .A1( u0_u2_n719 ) , .ZN( u0_u2_n720 ) );
  INV_X1 u0_u2_U11 (.A( u0_u2_n785 ) , .ZN( u0_u2_n874 ) );
  INV_X1 u0_u2_U110 (.A( u0_u2_n470 ) , .ZN( u0_u2_n871 ) );
  OAI21_X1 u0_u2_U111 (.ZN( u0_u2_n470 ) , .B1( u0_u2_n816 ) , .A( u0_u2_n841 ) , .B2( u0_u2_n858 ) );
  NAND2_X1 u0_u2_U112 (.ZN( u0_u2_n439 ) , .A2( u0_u2_n850 ) , .A1( u0_u2_n868 ) );
  NAND2_X1 u0_u2_U113 (.ZN( u0_u2_n440 ) , .A2( u0_u2_n838 ) , .A1( u0_u2_n861 ) );
  AOI221_X1 u0_u2_U114 (.A( u0_u2_n771 ) , .ZN( u0_u2_n781 ) , .C2( u0_u2_n817 ) , .B2( u0_u2_n842 ) , .C1( u0_u2_n862 ) , .B1( u0_u2_n873 ) );
  INV_X1 u0_u2_U115 (.A( u0_u2_n768 ) , .ZN( u0_u2_n842 ) );
  NAND2_X1 u0_u2_U116 (.A1( u0_u2_n454 ) , .A2( u0_u2_n472 ) , .ZN( u0_u2_n756 ) );
  AOI211_X1 u0_u2_U117 (.B( u0_u2_n814 ) , .A( u0_u2_n815 ) , .ZN( u0_u2_n831 ) , .C1( u0_u2_n849 ) , .C2( u0_u2_n857 ) );
  AOI211_X1 u0_u2_U118 (.A( u0_u2_n595 ) , .ZN( u0_u2_n604 ) , .B( u0_u2_n628 ) , .C1( u0_u2_n852 ) , .C2( u0_u2_n862 ) );
  INV_X1 u0_u2_U119 (.A( u0_u2_n737 ) , .ZN( u0_u2_n846 ) );
  INV_X1 u0_u2_U12 (.A( u0_u2_n686 ) , .ZN( u0_u2_n879 ) );
  NAND2_X1 u0_u2_U120 (.A1( u0_u2_n458 ) , .A2( u0_u2_n460 ) , .ZN( u0_u2_n769 ) );
  NOR3_X1 u0_u2_U121 (.ZN( u0_u2_n497 ) , .A1( u0_u2_n789 ) , .A2( u0_u2_n857 ) , .A3( u0_u2_n870 ) );
  OAI22_X1 u0_u2_U122 (.B2( u0_u2_n757 ) , .B1( u0_u2_n758 ) , .A1( u0_u2_n759 ) , .ZN( u0_u2_n763 ) , .A2( u0_u2_n813 ) );
  NOR2_X1 u0_u2_U123 (.ZN( u0_u2_n758 ) , .A2( u0_u2_n859 ) , .A1( u0_u2_n867 ) );
  NOR3_X1 u0_u2_U124 (.ZN( u0_u2_n759 ) , .A2( u0_u2_n860 ) , .A1( u0_u2_n870 ) , .A3( u0_u2_n872 ) );
  NOR2_X1 u0_u2_U125 (.ZN( u0_u2_n539 ) , .A2( u0_u2_n756 ) , .A1( u0_u2_n757 ) );
  NOR2_X1 u0_u2_U126 (.ZN( u0_u2_n577 ) , .A1( u0_u2_n735 ) , .A2( u0_u2_n813 ) );
  OAI21_X1 u0_u2_U127 (.ZN( u0_u2_n794 ) , .A( u0_u2_n846 ) , .B1( u0_u2_n870 ) , .B2( u0_u2_n880 ) );
  NOR2_X1 u0_u2_U128 (.A2( u0_u2_n715 ) , .A1( u0_u2_n757 ) , .ZN( u0_u2_n778 ) );
  NOR2_X1 u0_u2_U129 (.ZN( u0_u2_n516 ) , .A1( u0_u2_n736 ) , .A2( u0_u2_n786 ) );
  INV_X1 u0_u2_U13 (.A( u0_u2_n687 ) , .ZN( u0_u2_n847 ) );
  NOR2_X1 u0_u2_U130 (.ZN( u0_u2_n553 ) , .A2( u0_u2_n787 ) , .A1( u0_u2_n821 ) );
  NOR2_X1 u0_u2_U131 (.ZN( u0_u2_n618 ) , .A2( u0_u2_n787 ) , .A1( u0_u2_n813 ) );
  NOR2_X1 u0_u2_U132 (.ZN( u0_u2_n514 ) , .A1( u0_u2_n819 ) , .A2( u0_u2_n824 ) );
  NOR2_X1 u0_u2_U133 (.A2( u0_u2_n715 ) , .A1( u0_u2_n769 ) , .ZN( u0_u2_n801 ) );
  NOR2_X1 u0_u2_U134 (.ZN( u0_u2_n663 ) , .A1( u0_u2_n754 ) , .A2( u0_u2_n787 ) );
  NOR2_X1 u0_u2_U135 (.ZN( u0_u2_n513 ) , .A2( u0_u2_n735 ) , .A1( u0_u2_n769 ) );
  INV_X1 u0_u2_U136 (.A( u0_u2_n754 ) , .ZN( u0_u2_n841 ) );
  NOR2_X1 u0_u2_U137 (.ZN( u0_u2_n689 ) , .A2( u0_u2_n715 ) , .A1( u0_u2_n824 ) );
  INV_X1 u0_u2_U138 (.A( u0_u2_n735 ) , .ZN( u0_u2_n859 ) );
  AOI21_X1 u0_u2_U139 (.B1( u0_u2_n706 ) , .ZN( u0_u2_n707 ) , .A( u0_u2_n739 ) , .B2( u0_u2_n770 ) );
  AOI222_X1 u0_u2_U14 (.ZN( u0_u2_n570 ) , .B1( u0_u2_n837 ) , .C1( u0_u2_n848 ) , .A2( u0_u2_n850 ) , .A1( u0_u2_n861 ) , .B2( u0_u2_n870 ) , .C2( u0_u2_n880 ) );
  INV_X1 u0_u2_U140 (.A( u0_u2_n757 ) , .ZN( u0_u2_n849 ) );
  AOI21_X1 u0_u2_U141 (.ZN( u0_u2_n547 ) , .A( u0_u2_n770 ) , .B2( u0_u2_n786 ) , .B1( u0_u2_n824 ) );
  AOI21_X1 u0_u2_U142 (.ZN( u0_u2_n576 ) , .B1( u0_u2_n757 ) , .B2( u0_u2_n769 ) , .A( u0_u2_n787 ) );
  AOI21_X1 u0_u2_U143 (.B1( u0_u2_n693 ) , .ZN( u0_u2_n694 ) , .A( u0_u2_n735 ) , .B2( u0_u2_n768 ) );
  NOR2_X1 u0_u2_U144 (.ZN( u0_u2_n575 ) , .A1( u0_u2_n736 ) , .A2( u0_u2_n769 ) );
  NOR2_X1 u0_u2_U145 (.ZN( u0_u2_n536 ) , .A1( u0_u2_n715 ) , .A2( u0_u2_n786 ) );
  AOI21_X1 u0_u2_U146 (.ZN( u0_u2_n696 ) , .B2( u0_u2_n756 ) , .B1( u0_u2_n770 ) , .A( u0_u2_n813 ) );
  NOR2_X1 u0_u2_U147 (.ZN( u0_u2_n718 ) , .A1( u0_u2_n769 ) , .A2( u0_u2_n770 ) );
  INV_X1 u0_u2_U148 (.A( u0_u2_n787 ) , .ZN( u0_u2_n857 ) );
  NOR2_X1 u0_u2_U149 (.ZN( u0_u2_n621 ) , .A1( u0_u2_n769 ) , .A2( u0_u2_n819 ) );
  AOI222_X1 u0_u2_U15 (.ZN( u0_u2_n667 ) , .A2( u0_u2_n846 ) , .B1( u0_u2_n848 ) , .C2( u0_u2_n852 ) , .A1( u0_u2_n867 ) , .C1( u0_u2_n870 ) , .B2( u0_u2_n877 ) );
  AOI21_X1 u0_u2_U150 (.B1( u0_u2_n444 ) , .ZN( u0_u2_n634 ) , .A( u0_u2_n770 ) , .B2( u0_u2_n821 ) );
  INV_X1 u0_u2_U151 (.A( u0_u2_n736 ) , .ZN( u0_u2_n875 ) );
  NOR2_X1 u0_u2_U152 (.ZN( u0_u2_n527 ) , .A2( u0_u2_n715 ) , .A1( u0_u2_n821 ) );
  NOR2_X1 u0_u2_U153 (.ZN( u0_u2_n584 ) , .A2( u0_u2_n706 ) , .A1( u0_u2_n821 ) );
  INV_X1 u0_u2_U154 (.A( u0_u2_n706 ) , .ZN( u0_u2_n860 ) );
  OAI21_X1 u0_u2_U155 (.A( u0_u2_n705 ) , .ZN( u0_u2_n709 ) , .B2( u0_u2_n757 ) , .B1( u0_u2_n811 ) );
  OAI21_X1 u0_u2_U156 (.ZN( u0_u2_n705 ) , .B2( u0_u2_n840 ) , .B1( u0_u2_n845 ) , .A( u0_u2_n867 ) );
  INV_X1 u0_u2_U157 (.A( u0_u2_n770 ) , .ZN( u0_u2_n873 ) );
  NAND2_X1 u0_u2_U158 (.A1( u0_u2_n706 ) , .A2( u0_u2_n736 ) , .ZN( u0_u2_n789 ) );
  BUF_X1 u0_u2_U159 (.Z( u0_u2_n443 ) , .A( u0_u2_n822 ) );
  INV_X1 u0_u2_U16 (.A( u0_u2_n654 ) , .ZN( u0_u2_n877 ) );
  INV_X1 u0_u2_U160 (.A( u0_u2_n824 ) , .ZN( u0_u2_n851 ) );
  NAND2_X1 u0_u2_U161 (.ZN( u0_u2_n721 ) , .A1( u0_u2_n735 ) , .A2( u0_u2_n787 ) );
  BUF_X1 u0_u2_U162 (.Z( u0_u2_n442 ) , .A( u0_u2_n676 ) );
  BUF_X1 u0_u2_U163 (.Z( u0_u2_n441 ) , .A( u0_u2_n704 ) );
  OR4_X1 u0_u2_U164 (.A3( u0_u2_n587 ) , .A4( u0_u2_n588 ) , .A2( u0_u2_n589 ) , .A1( u0_u2_n590 ) , .ZN( u0_u2_n591 ) );
  OAI222_X1 u0_u2_U165 (.A2( u0_u2_n443 ) , .B2( u0_u2_n715 ) , .ZN( u0_u2_n716 ) , .C2( u0_u2_n731 ) , .B1( u0_u2_n754 ) , .A1( u0_u2_n813 ) , .C1( u0_u2_n821 ) );
  AOI221_X1 u0_u2_U166 (.A( u0_u2_n457 ) , .ZN( u0_u2_n466 ) , .C2( u0_u2_n760 ) , .B1( u0_u2_n839 ) , .C1( u0_u2_n849 ) , .B2( u0_u2_n868 ) );
  OAI221_X1 u0_u2_U167 (.A( u0_u2_n790 ) , .C2( u0_u2_n791 ) , .B2( u0_u2_n792 ) , .B1( u0_u2_n793 ) , .ZN( u0_u2_n803 ) , .C1( u0_u2_n820 ) );
  OAI221_X1 u0_u2_U168 (.A( u0_u2_n703 ) , .ZN( u0_u2_n710 ) , .C2( u0_u2_n791 ) , .C1( u0_u2_n792 ) , .B1( u0_u2_n793 ) , .B2( u0_u2_n813 ) );
  AOI22_X1 u0_u2_U169 (.ZN( u0_u2_n703 ) , .A1( u0_u2_n837 ) , .B2( u0_u2_n850 ) , .A2( u0_u2_n872 ) , .B1( u0_u2_n875 ) );
  NOR4_X1 u0_u2_U17 (.A4( u0_u2_n551 ) , .A3( u0_u2_n552 ) , .A2( u0_u2_n553 ) , .A1( u0_u2_n554 ) , .ZN( u0_u2_n555 ) );
  OAI221_X1 u0_u2_U170 (.A( u0_u2_n734 ) , .C2( u0_u2_n735 ) , .B2( u0_u2_n736 ) , .B1( u0_u2_n737 ) , .ZN( u0_u2_n744 ) , .C1( u0_u2_n824 ) );
  NAND2_X1 u0_u2_U171 (.A2( u0_u2_n467 ) , .A1( u0_u2_n472 ) , .ZN( u0_u2_n787 ) );
  NAND2_X1 u0_u2_U172 (.A2( u0_u2_n478 ) , .A1( u0_u2_n479 ) , .ZN( u0_u2_n824 ) );
  NAND2_X1 u0_u2_U173 (.A1( u0_u2_n456 ) , .A2( u0_u2_n467 ) , .ZN( u0_u2_n799 ) );
  NAND2_X1 u0_u2_U174 (.A2( u0_u2_n455 ) , .A1( u0_u2_n467 ) , .ZN( u0_u2_n735 ) );
  NAND2_X1 u0_u2_U175 (.A2( u0_u2_n456 ) , .A1( u0_u2_n459 ) , .ZN( u0_u2_n770 ) );
  NAND2_X1 u0_u2_U176 (.A2( u0_u2_n461 ) , .A1( u0_u2_n479 ) , .ZN( u0_u2_n786 ) );
  NAND2_X1 u0_u2_U177 (.A1( u0_u2_n448 ) , .A2( u0_u2_n467 ) , .ZN( u0_u2_n706 ) );
  NAND2_X1 u0_u2_U178 (.A1( u0_u2_n460 ) , .A2( u0_u2_n479 ) , .ZN( u0_u2_n792 ) );
  NAND2_X1 u0_u2_U179 (.A2( u0_u2_n455 ) , .A1( u0_u2_n459 ) , .ZN( u0_u2_n736 ) );
  NOR4_X1 u0_u2_U18 (.A4( u0_u2_n539 ) , .A3( u0_u2_n540 ) , .A2( u0_u2_n541 ) , .ZN( u0_u2_n542 ) , .A1( u0_u2_n827 ) );
  NAND2_X1 u0_u2_U180 (.A2( u0_u2_n471 ) , .A1( u0_u2_n472 ) , .ZN( u0_u2_n819 ) );
  NAND2_X1 u0_u2_U181 (.A1( u0_u2_n462 ) , .A2( u0_u2_n478 ) , .ZN( u0_u2_n810 ) );
  NAND2_X1 u0_u2_U182 (.A1( u0_u2_n458 ) , .A2( u0_u2_n478 ) , .ZN( u0_u2_n823 ) );
  NAND2_X1 u0_u2_U183 (.A2( u0_u2_n448 ) , .A1( u0_u2_n454 ) , .ZN( u0_u2_n791 ) );
  NAND2_X1 u0_u2_U184 (.A1( u0_u2_n461 ) , .A2( u0_u2_n468 ) , .ZN( u0_u2_n820 ) );
  NOR2_X1 u0_u2_U185 (.ZN( u0_u2_n460 ) , .A1( u0_u2_n833 ) , .A2( u0_u2_n834 ) );
  NAND2_X1 u0_u2_U186 (.A2( u0_u2_n468 ) , .A1( u0_u2_n469 ) , .ZN( u0_u2_n754 ) );
  NAND2_X1 u0_u2_U187 (.A1( u0_u2_n454 ) , .A2( u0_u2_n455 ) , .ZN( u0_u2_n793 ) );
  NAND2_X1 u0_u2_U188 (.A1( u0_u2_n448 ) , .A2( u0_u2_n471 ) , .ZN( u0_u2_n715 ) );
  NAND2_X1 u0_u2_U189 (.A1( u0_u2_n469 ) , .A2( u0_u2_n479 ) , .ZN( u0_u2_n795 ) );
  NOR4_X1 u0_u2_U19 (.A4( u0_u2_n452 ) , .A3( u0_u2_n453 ) , .A2( u0_u2_n523 ) , .A1( u0_u2_n548 ) , .ZN( u0_u2_n713 ) );
  NAND2_X1 u0_u2_U190 (.A2( u0_u2_n448 ) , .A1( u0_u2_n459 ) , .ZN( u0_u2_n798 ) );
  NAND2_X1 u0_u2_U191 (.A1( u0_u2_n458 ) , .A2( u0_u2_n469 ) , .ZN( u0_u2_n797 ) );
  NAND2_X1 u0_u2_U192 (.A2( u0_u2_n461 ) , .A1( u0_u2_n462 ) , .ZN( u0_u2_n737 ) );
  AOI222_X1 u0_u2_U193 (.B2( u0_u2_n645 ) , .ZN( u0_u2_n651 ) , .B1( u0_u2_n848 ) , .A1( u0_u2_n849 ) , .C2( u0_u2_n853 ) , .C1( u0_u2_n870 ) , .A2( u0_u2_n872 ) );
  NOR4_X1 u0_u2_U194 (.A4( u0_u2_n646 ) , .A3( u0_u2_n647 ) , .A2( u0_u2_n648 ) , .A1( u0_u2_n649 ) , .ZN( u0_u2_n650 ) );
  NAND4_X1 u0_u2_U195 (.ZN( u0_subword_8 ) , .A4( u0_u2_n508 ) , .A3( u0_u2_n509 ) , .A2( u0_u2_n510 ) , .A1( u0_u2_n511 ) );
  NOR4_X1 u0_u2_U196 (.A4( u0_u2_n505 ) , .A3( u0_u2_n506 ) , .A2( u0_u2_n507 ) , .ZN( u0_u2_n508 ) , .A1( u0_u2_n534 ) );
  AOI221_X1 u0_u2_U197 (.A( u0_u2_n504 ) , .ZN( u0_u2_n509 ) , .B2( u0_u2_n850 ) , .C1( u0_u2_n853 ) , .C2( u0_u2_n867 ) , .B1( u0_u2_n869 ) );
  AOI221_X1 u0_u2_U198 (.A( u0_u2_n788 ) , .ZN( u0_u2_n805 ) , .C2( u0_u2_n844 ) , .B2( u0_u2_n845 ) , .B1( u0_u2_n872 ) , .C1( u0_u2_n873 ) );
  NOR4_X1 u0_u2_U199 (.A4( u0_u2_n800 ) , .A3( u0_u2_n801 ) , .A2( u0_u2_n802 ) , .A1( u0_u2_n803 ) , .ZN( u0_u2_n804 ) );
  OR4_X1 u0_u2_U20 (.A4( u0_u2_n449 ) , .A2( u0_u2_n450 ) , .A1( u0_u2_n451 ) , .ZN( u0_u2_n452 ) , .A3( u0_u2_n560 ) );
  NOR4_X1 u0_u2_U200 (.A4( u0_u2_n707 ) , .A3( u0_u2_n708 ) , .A2( u0_u2_n709 ) , .A1( u0_u2_n710 ) , .ZN( u0_u2_n711 ) );
  AOI211_X1 u0_u2_U201 (.B( u0_u2_n701 ) , .A( u0_u2_n702 ) , .ZN( u0_u2_n712 ) , .C2( u0_u2_n838 ) , .C1( u0_u2_n858 ) );
  NAND4_X1 u0_u2_U202 (.ZN( u0_subword_15 ) , .A4( u0_u2_n829 ) , .A3( u0_u2_n830 ) , .A2( u0_u2_n831 ) , .A1( u0_u2_n832 ) );
  NOR4_X1 u0_u2_U203 (.A4( u0_u2_n825 ) , .A3( u0_u2_n826 ) , .A2( u0_u2_n827 ) , .A1( u0_u2_n828 ) , .ZN( u0_u2_n829 ) );
  NAND4_X1 u0_u2_U204 (.ZN( u0_subword_9 ) , .A4( u0_u2_n602 ) , .A3( u0_u2_n603 ) , .A2( u0_u2_n604 ) , .A1( u0_u2_n605 ) );
  NOR4_X1 u0_u2_U205 (.A4( u0_u2_n598 ) , .A3( u0_u2_n599 ) , .A2( u0_u2_n600 ) , .A1( u0_u2_n601 ) , .ZN( u0_u2_n602 ) );
  AOI211_X1 u0_u2_U206 (.B( u0_u2_n596 ) , .A( u0_u2_n597 ) , .ZN( u0_u2_n603 ) , .C2( u0_u2_n818 ) , .C1( u0_u2_n840 ) );
  NOR4_X1 u0_u2_U207 (.A3( u0_u2_n762 ) , .A2( u0_u2_n763 ) , .A1( u0_u2_n764 ) , .ZN( u0_u2_n765 ) , .A4( u0_u2_n876 ) );
  AOI211_X1 u0_u2_U208 (.B( u0_u2_n752 ) , .A( u0_u2_n753 ) , .ZN( u0_u2_n766 ) , .C1( u0_u2_n839 ) , .C2( u0_u2_n860 ) );
  NOR4_X1 u0_u2_U209 (.A4( u0_u2_n741 ) , .A3( u0_u2_n742 ) , .A2( u0_u2_n743 ) , .A1( u0_u2_n744 ) , .ZN( u0_u2_n745 ) );
  INV_X1 u0_u2_U21 (.A( u0_u2_n620 ) , .ZN( u0_u2_n882 ) );
  AOI211_X1 u0_u2_U210 (.B( u0_u2_n732 ) , .A( u0_u2_n733 ) , .ZN( u0_u2_n746 ) , .C1( u0_u2_n850 ) , .C2( u0_u2_n862 ) );
  AOI221_X1 u0_u2_U211 (.ZN( u0_u2_n475 ) , .C2( u0_u2_n721 ) , .B2( u0_u2_n838 ) , .C1( u0_u2_n852 ) , .B1( u0_u2_n867 ) , .A( u0_u2_n871 ) );
  AOI22_X1 u0_u2_U212 (.A2( u0_u2_n789 ) , .ZN( u0_u2_n790 ) , .B2( u0_u2_n838 ) , .A1( u0_u2_n841 ) , .B1( u0_u2_n870 ) );
  NAND2_X1 u0_u2_U213 (.A1( u0_u2_n460 ) , .A2( u0_u2_n468 ) , .ZN( u0_u2_n751 ) );
  NAND2_X1 u0_u2_U214 (.A1( u0_u2_n454 ) , .A2( u0_u2_n456 ) , .ZN( u0_u2_n812 ) );
  NAND2_X1 u0_u2_U215 (.A2( u0_u2_n460 ) , .A1( u0_u2_n462 ) , .ZN( u0_u2_n813 ) );
  NAND2_X1 u0_u2_U216 (.A1( u0_u2_n456 ) , .A2( u0_u2_n471 ) , .ZN( u0_u2_n731 ) );
  AOI21_X1 u0_u2_U217 (.ZN( u0_u2_n522 ) , .A( u0_u2_n736 ) , .B1( u0_u2_n757 ) , .B2( u0_u2_n810 ) );
  NOR2_X1 u0_u2_U218 (.ZN( u0_u2_n690 ) , .A2( u0_u2_n706 ) , .A1( u0_u2_n810 ) );
  NOR2_X1 u0_u2_U219 (.A1( u0_u2_n756 ) , .ZN( u0_u2_n774 ) , .A2( u0_u2_n810 ) );
  NOR4_X1 u0_u2_U22 (.ZN( u0_u2_n493 ) , .A1( u0_u2_n514 ) , .A2( u0_u2_n526 ) , .A4( u0_u2_n553 ) , .A3( u0_u2_n618 ) );
  NOR2_X1 u0_u2_U220 (.ZN( u0_u2_n524 ) , .A1( u0_u2_n715 ) , .A2( u0_u2_n810 ) );
  NOR2_X1 u0_u2_U221 (.ZN( u0_u2_n673 ) , .A1( u0_u2_n735 ) , .A2( u0_u2_n810 ) );
  NOR2_X1 u0_u2_U222 (.ZN( u0_u2_n608 ) , .A2( u0_u2_n787 ) , .A1( u0_u2_n810 ) );
  NAND2_X1 u0_u2_U223 (.A2( u0_u2_n468 ) , .A1( u0_u2_n478 ) , .ZN( u0_u2_n704 ) );
  NAND2_X1 u0_u2_U224 (.A1( u0_u2_n459 ) , .A2( u0_u2_n472 ) , .ZN( u0_u2_n676 ) );
  NAND2_X1 u0_u2_U225 (.A2( u0_u2_n455 ) , .A1( u0_u2_n471 ) , .ZN( u0_u2_n822 ) );
  NOR2_X1 u0_u2_U226 (.ZN( u0_u2_n458 ) , .A1( u0_u2_n835 ) , .A2( u0_u2_n836 ) );
  OR3_X1 u0_u2_U227 (.ZN( u0_u2_n453 ) , .A1( u0_u2_n535 ) , .A3( u0_u2_n584 ) , .A2( u0_u2_n882 ) );
  NAND2_X1 u0_u2_U228 (.A1( u0_u2_n458 ) , .A2( u0_u2_n461 ) , .ZN( u0_u2_n821 ) );
  AOI211_X1 u0_u2_U229 (.A( u0_u2_n503 ) , .ZN( u0_u2_n510 ) , .B( u0_u2_n809 ) , .C2( u0_u2_n846 ) , .C1( u0_u2_n858 ) );
  NOR4_X1 u0_u2_U23 (.ZN( u0_u2_n482 ) , .A1( u0_u2_n538 ) , .A3( u0_u2_n575 ) , .A4( u0_u2_n607 ) , .A2( u0_u2_n649 ) );
  NAND4_X1 u0_u2_U230 (.A4( u0_u2_n500 ) , .A3( u0_u2_n501 ) , .A1( u0_u2_n502 ) , .ZN( u0_u2_n809 ) , .A2( u0_u2_n874 ) );
  NOR4_X1 u0_u2_U231 (.A3( u0_u2_n445 ) , .A2( u0_u2_n498 ) , .A1( u0_u2_n499 ) , .ZN( u0_u2_n500 ) , .A4( u0_u2_n619 ) );
  OAI22_X1 u0_u2_U232 (.B1( u0_u2_n497 ) , .ZN( u0_u2_n498 ) , .A1( u0_u2_n693 ) , .A2( u0_u2_n770 ) , .B2( u0_u2_n824 ) );
  NOR2_X1 u0_u2_U233 (.ZN( u0_u2_n444 ) , .A2( u0_u2_n843 ) , .A1( u0_u2_n846 ) );
  NOR2_X1 u0_u2_U234 (.ZN( u0_u2_n632 ) , .A2( u0_u2_n843 ) , .A1( u0_u2_n846 ) );
  NOR2_X1 u0_u2_U235 (.ZN( u0_u2_n445 ) , .A2( u0_u2_n704 ) , .A1( u0_u2_n798 ) );
  OAI222_X1 u0_u2_U236 (.A2( u0_u2_n442 ) , .C1( u0_u2_n443 ) , .ZN( u0_u2_n681 ) , .B1( u0_u2_n754 ) , .B2( u0_u2_n791 ) , .C2( u0_u2_n795 ) , .A1( u0_u2_n824 ) );
  NOR4_X1 u0_u2_U237 (.A4( u0_u2_n491 ) , .ZN( u0_u2_n494 ) , .A1( u0_u2_n573 ) , .A2( u0_u2_n588 ) , .A3( u0_u2_n609 ) );
  AOI222_X1 u0_u2_U238 (.ZN( u0_u2_n613 ) , .A1( u0_u2_n837 ) , .C2( u0_u2_n844 ) , .B1( u0_u2_n849 ) , .A2( u0_u2_n863 ) , .B2( u0_u2_n868 ) , .C1( u0_u2_n875 ) );
  AOI222_X1 u0_u2_U239 (.ZN( u0_u2_n532 ) , .A1( u0_u2_n841 ) , .B2( u0_u2_n844 ) , .C1( u0_u2_n851 ) , .C2( u0_u2_n857 ) , .A2( u0_u2_n859 ) , .B1( u0_u2_n873 ) );
  INV_X1 u0_u2_U24 (.A( u0_u2_n756 ) , .ZN( u0_u2_n870 ) );
  NAND2_X1 u0_u2_U240 (.ZN( u0_u2_n620 ) , .A2( u0_u2_n844 ) , .A1( u0_u2_n880 ) );
  NAND4_X1 u0_u2_U241 (.A4( u0_u2_n486 ) , .A3( u0_u2_n487 ) , .A2( u0_u2_n488 ) , .A1( u0_u2_n489 ) , .ZN( u0_u2_n701 ) );
  NOR2_X1 u0_u2_U242 (.ZN( u0_u2_n586 ) , .A2( u0_u2_n715 ) , .A1( u0_u2_n737 ) );
  OAI21_X1 u0_u2_U243 (.A( u0_u2_n794 ) , .B2( u0_u2_n795 ) , .B1( u0_u2_n796 ) , .ZN( u0_u2_n802 ) );
  AOI21_X1 u0_u2_U244 (.ZN( u0_u2_n646 ) , .B2( u0_u2_n756 ) , .A( u0_u2_n795 ) , .B1( u0_u2_n819 ) );
  AOI21_X1 u0_u2_U245 (.ZN( u0_u2_n449 ) , .A( u0_u2_n706 ) , .B1( u0_u2_n740 ) , .B2( u0_u2_n757 ) );
  NOR2_X1 u0_u2_U246 (.ZN( u0_u2_n525 ) , .A1( u0_u2_n715 ) , .A2( u0_u2_n795 ) );
  INV_X1 u0_u2_U247 (.A( u0_u2_n795 ) , .ZN( u0_u2_n852 ) );
  NOR2_X1 u0_u2_U248 (.ZN( u0_u2_n456 ) , .A1( u0_u2_n855 ) , .A2( w3_4 ) );
  NOR2_X1 u0_u2_U249 (.ZN( u0_u2_n472 ) , .A2( u0_u2_n854 ) , .A1( u0_u2_n855 ) );
  NOR4_X1 u0_u2_U25 (.ZN( u0_u2_n486 ) , .A1( u0_u2_n527 ) , .A4( u0_u2_n564 ) , .A3( u0_u2_n589 ) , .A2( u0_u2_n637 ) );
  OAI222_X1 u0_u2_U250 (.B1( u0_u2_n441 ) , .ZN( u0_u2_n624 ) , .C1( u0_u2_n731 ) , .C2( u0_u2_n754 ) , .B2( u0_u2_n793 ) , .A2( u0_u2_n799 ) , .A1( u0_u2_n823 ) );
  NOR2_X1 u0_u2_U251 (.ZN( u0_u2_n467 ) , .A1( u0_u2_n856 ) , .A2( w3_7 ) );
  AOI21_X1 u0_u2_U252 (.ZN( u0_u2_n647 ) , .B2( u0_u2_n754 ) , .A( u0_u2_n799 ) , .B1( u0_u2_n810 ) );
  AOI21_X1 u0_u2_U253 (.A( u0_u2_n740 ) , .ZN( u0_u2_n741 ) , .B2( u0_u2_n787 ) , .B1( u0_u2_n799 ) );
  AOI21_X1 u0_u2_U254 (.ZN( u0_u2_n521 ) , .A( u0_u2_n786 ) , .B2( u0_u2_n799 ) , .B1( u0_u2_n819 ) );
  AOI21_X1 u0_u2_U255 (.B2( u0_u2_n770 ) , .ZN( u0_u2_n771 ) , .A( u0_u2_n795 ) , .B1( u0_u2_n799 ) );
  INV_X1 u0_u2_U256 (.A( u0_u2_n799 ) , .ZN( u0_u2_n858 ) );
  NOR2_X1 u0_u2_U257 (.ZN( u0_u2_n564 ) , .A1( u0_u2_n799 ) , .A2( u0_u2_n821 ) );
  NOR2_X1 u0_u2_U258 (.ZN( u0_u2_n590 ) , .A1( u0_u2_n799 ) , .A2( u0_u2_n824 ) );
  AOI221_X1 u0_u2_U259 (.A( u0_u2_n496 ) , .ZN( u0_u2_n501 ) , .B2( u0_u2_n843 ) , .C2( u0_u2_n848 ) , .C1( u0_u2_n858 ) , .B1( u0_u2_n867 ) );
  NOR3_X1 u0_u2_U26 (.ZN( u0_u2_n487 ) , .A2( u0_u2_n515 ) , .A3( u0_u2_n608 ) , .A1( u0_u2_n617 ) );
  NOR3_X1 u0_u2_U260 (.ZN( u0_u2_n447 ) , .A2( u0_u2_n843 ) , .A3( u0_u2_n844 ) , .A1( u0_u2_n853 ) );
  NOR4_X1 u0_u2_U261 (.A3( u0_u2_n680 ) , .A1( u0_u2_n681 ) , .ZN( u0_u2_n682 ) , .A4( u0_u2_n722 ) , .A2( u0_u2_n866 ) );
  INV_X1 u0_u2_U262 (.A( u0_u2_n679 ) , .ZN( u0_u2_n866 ) );
  NOR2_X1 u0_u2_U263 (.ZN( u0_u2_n478 ) , .A1( u0_u2_n833 ) , .A2( w3_1 ) );
  INV_X1 u0_u2_U264 (.ZN( u0_u2_n834 ) , .A( w3_1 ) );
  CLKBUF_X1 u0_u2_U265 (.Z( u0_u2_n446 ) , .A( u0_u2_n798 ) );
  NOR2_X1 u0_u2_U266 (.A2( u0_u2_n438 ) , .A1( u0_u2_n583 ) , .ZN( u0_u2_n594 ) );
  OAI22_X1 u0_u2_U267 (.B2( u0_u2_n786 ) , .B1( u0_u2_n787 ) , .ZN( u0_u2_n788 ) , .A2( u0_u2_n821 ) , .A1( u0_u2_n822 ) );
  AOI21_X1 u0_u2_U268 (.B1( u0_u2_n443 ) , .ZN( u0_u2_n596 ) , .B2( u0_u2_n706 ) , .A( u0_u2_n824 ) );
  INV_X1 u0_u2_U269 (.A( u0_u2_n822 ) , .ZN( u0_u2_n862 ) );
  AOI211_X1 u0_u2_U27 (.B( u0_u2_n484 ) , .A( u0_u2_n485 ) , .ZN( u0_u2_n489 ) , .C2( u0_u2_n840 ) , .C1( u0_u2_n868 ) );
  NOR2_X1 u0_u2_U270 (.ZN( u0_u2_n674 ) , .A1( u0_u2_n757 ) , .A2( u0_u2_n822 ) );
  NOR2_X1 u0_u2_U271 (.A1( u0_u2_n443 ) , .ZN( u0_u2_n477 ) , .A2( u0_u2_n786 ) );
  AOI21_X1 u0_u2_U272 (.B1( u0_u2_n443 ) , .ZN( u0_u2_n546 ) , .B2( u0_u2_n819 ) , .A( u0_u2_n821 ) );
  AOI21_X1 u0_u2_U273 (.B1( u0_u2_n443 ) , .ZN( u0_u2_n457 ) , .B2( u0_u2_n799 ) , .A( u0_u2_n810 ) );
  NOR2_X1 u0_u2_U274 (.A2( u0_u2_n443 ) , .ZN( u0_u2_n637 ) , .A1( u0_u2_n754 ) );
  INV_X1 u0_u2_U275 (.ZN( u0_u2_n865 ) , .A( w3_7 ) );
  AOI222_X1 u0_u2_U276 (.C2( u0_u2_n816 ) , .B2( u0_u2_n817 ) , .A2( u0_u2_n818 ) , .ZN( u0_u2_n830 ) , .C1( u0_u2_n839 ) , .A1( u0_u2_n846 ) , .B1( u0_u2_n860 ) );
  AOI22_X1 u0_u2_U277 (.ZN( u0_u2_n734 ) , .B1( u0_u2_n839 ) , .A2( u0_u2_n845 ) , .A1( u0_u2_n870 ) , .B2( u0_u2_n873 ) );
  AOI222_X1 u0_u2_U278 (.ZN( u0_u2_n476 ) , .B1( u0_u2_n839 ) , .A1( u0_u2_n846 ) , .C1( u0_u2_n849 ) , .C2( u0_u2_n858 ) , .A2( u0_u2_n862 ) , .B2( u0_u2_n872 ) );
  NOR2_X1 u0_u2_U279 (.A2( u0_u2_n443 ) , .ZN( u0_u2_n662 ) , .A1( u0_u2_n797 ) );
  NOR4_X1 u0_u2_U28 (.ZN( u0_u2_n488 ) , .A3( u0_u2_n539 ) , .A4( u0_u2_n552 ) , .A2( u0_u2_n574 ) , .A1( u0_u2_n724 ) );
  NOR2_X1 u0_u2_U280 (.ZN( u0_u2_n693 ) , .A1( u0_u2_n838 ) , .A2( u0_u2_n839 ) );
  NOR2_X1 u0_u2_U281 (.ZN( u0_u2_n528 ) , .A1( u0_u2_n797 ) , .A2( u0_u2_n819 ) );
  NOR2_X1 u0_u2_U282 (.ZN( u0_u2_n740 ) , .A2( u0_u2_n839 ) , .A1( u0_u2_n852 ) );
  NOR2_X1 u0_u2_U283 (.ZN( u0_u2_n668 ) , .A1( u0_u2_n736 ) , .A2( u0_u2_n797 ) );
  NOR2_X1 u0_u2_U284 (.ZN( u0_u2_n675 ) , .A2( u0_u2_n715 ) , .A1( u0_u2_n797 ) );
  INV_X1 u0_u2_U285 (.A( u0_u2_n797 ) , .ZN( u0_u2_n839 ) );
  NOR2_X1 u0_u2_U286 (.ZN( u0_u2_n468 ) , .A1( u0_u2_n836 ) , .A2( w3_2 ) );
  INV_X1 u0_u2_U287 (.ZN( u0_u2_n835 ) , .A( w3_2 ) );
  AOI21_X1 u0_u2_U288 (.ZN( u0_u2_n600 ) , .B1( u0_u2_n757 ) , .A( u0_u2_n799 ) , .B2( u0_u2_n820 ) );
  AOI21_X1 u0_u2_U289 (.A( u0_u2_n819 ) , .B2( u0_u2_n820 ) , .B1( u0_u2_n821 ) , .ZN( u0_u2_n826 ) );
  NOR2_X1 u0_u2_U29 (.ZN( u0_u2_n687 ) , .A2( u0_u2_n841 ) , .A1( u0_u2_n846 ) );
  AOI21_X1 u0_u2_U290 (.ZN( u0_u2_n656 ) , .B1( u0_u2_n736 ) , .B2( u0_u2_n770 ) , .A( u0_u2_n820 ) );
  NOR2_X1 u0_u2_U291 (.A2( u0_u2_n820 ) , .A1( u0_u2_n822 ) , .ZN( u0_u2_n828 ) );
  NOR2_X1 u0_u2_U292 (.ZN( u0_u2_n585 ) , .A1( u0_u2_n715 ) , .A2( u0_u2_n820 ) );
  NOR2_X1 u0_u2_U293 (.ZN( u0_u2_n672 ) , .A1( u0_u2_n787 ) , .A2( u0_u2_n820 ) );
  NOR2_X1 u0_u2_U294 (.A1( u0_u2_n706 ) , .ZN( u0_u2_n775 ) , .A2( u0_u2_n820 ) );
  NOR2_X1 u0_u2_U295 (.ZN( u0_u2_n661 ) , .A1( u0_u2_n735 ) , .A2( u0_u2_n820 ) );
  INV_X1 u0_u2_U296 (.A( u0_u2_n820 ) , .ZN( u0_u2_n843 ) );
  AOI21_X1 u0_u2_U297 (.ZN( u0_u2_n598 ) , .B2( u0_u2_n770 ) , .A( u0_u2_n792 ) , .B1( u0_u2_n819 ) );
  AND2_X1 u0_u2_U298 (.ZN( u0_u2_n739 ) , .A1( u0_u2_n786 ) , .A2( u0_u2_n792 ) );
  NOR2_X1 u0_u2_U299 (.ZN( u0_u2_n670 ) , .A1( u0_u2_n736 ) , .A2( u0_u2_n792 ) );
  NAND2_X1 u0_u2_U3 (.ZN( u0_u2_n438 ) , .A1( u0_u2_n439 ) , .A2( u0_u2_n440 ) );
  NAND4_X1 u0_u2_U30 (.A4( u0_u2_n610 ) , .A3( u0_u2_n611 ) , .A2( u0_u2_n612 ) , .A1( u0_u2_n613 ) , .ZN( u0_u2_n729 ) );
  NOR2_X1 u0_u2_U300 (.ZN( u0_u2_n515 ) , .A2( u0_u2_n787 ) , .A1( u0_u2_n792 ) );
  NOR2_X1 u0_u2_U301 (.A2( u0_u2_n443 ) , .ZN( u0_u2_n622 ) , .A1( u0_u2_n792 ) );
  INV_X1 u0_u2_U302 (.A( u0_u2_n792 ) , .ZN( u0_u2_n853 ) );
  OAI22_X1 u0_u2_U303 (.ZN( u0_u2_n490 ) , .A1( u0_u2_n715 ) , .B2( u0_u2_n792 ) , .A2( u0_u2_n813 ) , .B1( u0_u2_n819 ) );
  NOR2_X1 u0_u2_U304 (.ZN( u0_u2_n636 ) , .A2( u0_u2_n735 ) , .A1( u0_u2_n792 ) );
  NOR2_X1 u0_u2_U305 (.ZN( u0_u2_n550 ) , .A2( u0_u2_n715 ) , .A1( u0_u2_n792 ) );
  NOR2_X1 u0_u2_U306 (.ZN( u0_u2_n551 ) , .A2( u0_u2_n792 ) , .A1( u0_u2_n799 ) );
  NAND4_X1 u0_u2_U307 (.A4( u0_u2_n698 ) , .A3( u0_u2_n699 ) , .A1( u0_u2_n700 ) , .ZN( u0_u2_n783 ) , .A2( u0_u2_n879 ) );
  NOR4_X1 u0_u2_U308 (.A4( u0_u2_n783 ) , .A3( u0_u2_n784 ) , .A1( u0_u2_n785 ) , .ZN( u0_u2_n806 ) , .A2( u0_u2_n808 ) );
  AOI211_X1 u0_u2_U309 (.A( u0_u2_n644 ) , .ZN( u0_u2_n652 ) , .B( u0_u2_n750 ) , .C2( u0_u2_n846 ) , .C1( u0_u2_n861 ) );
  NOR3_X1 u0_u2_U31 (.A1( u0_u2_n606 ) , .ZN( u0_u2_n611 ) , .A3( u0_u2_n670 ) , .A2( u0_u2_n777 ) );
  NOR3_X1 u0_u2_U310 (.A3( u0_u2_n748 ) , .A2( u0_u2_n749 ) , .A1( u0_u2_n750 ) , .ZN( u0_u2_n767 ) );
  NAND4_X1 u0_u2_U311 (.A4( u0_u2_n640 ) , .A3( u0_u2_n641 ) , .A2( u0_u2_n642 ) , .A1( u0_u2_n643 ) , .ZN( u0_u2_n750 ) );
  NOR3_X1 u0_u2_U312 (.A3( u0_u2_n628 ) , .A2( u0_u2_n629 ) , .ZN( u0_u2_n643 ) , .A1( u0_u2_n732 ) );
  NOR4_X1 u0_u2_U313 (.A4( u0_u2_n621 ) , .A3( u0_u2_n622 ) , .A2( u0_u2_n623 ) , .A1( u0_u2_n624 ) , .ZN( u0_u2_n625 ) );
  NOR2_X1 u0_u2_U314 (.ZN( u0_u2_n459 ) , .A1( u0_u2_n865 ) , .A2( w3_6 ) );
  NOR2_X1 u0_u2_U315 (.ZN( u0_u2_n454 ) , .A2( u0_u2_n856 ) , .A1( u0_u2_n865 ) );
  NOR2_X1 u0_u2_U316 (.ZN( u0_u2_n471 ) , .A2( w3_6 ) , .A1( w3_7 ) );
  INV_X1 u0_u2_U317 (.ZN( u0_u2_n856 ) , .A( w3_6 ) );
  AOI21_X1 u0_u2_U318 (.ZN( u0_u2_n505 ) , .A( u0_u2_n731 ) , .B2( u0_u2_n769 ) , .B1( u0_u2_n821 ) );
  OAI22_X1 u0_u2_U319 (.ZN( u0_u2_n496 ) , .A1( u0_u2_n731 ) , .B2( u0_u2_n735 ) , .B1( u0_u2_n737 ) , .A2( u0_u2_n786 ) );
  NOR4_X1 u0_u2_U32 (.A3( u0_u2_n607 ) , .A2( u0_u2_n608 ) , .A1( u0_u2_n609 ) , .ZN( u0_u2_n610 ) , .A4( u0_u2_n662 ) );
  NOR2_X1 u0_u2_U320 (.ZN( u0_u2_n719 ) , .A2( u0_u2_n731 ) , .A1( u0_u2_n797 ) );
  NOR2_X1 u0_u2_U321 (.ZN( u0_u2_n535 ) , .A2( u0_u2_n731 ) , .A1( u0_u2_n810 ) );
  NOR2_X1 u0_u2_U322 (.ZN( u0_u2_n616 ) , .A2( u0_u2_n731 ) , .A1( u0_u2_n824 ) );
  NOR2_X1 u0_u2_U323 (.ZN( u0_u2_n533 ) , .A1( u0_u2_n731 ) , .A2( u0_u2_n757 ) );
  NOR2_X1 u0_u2_U324 (.ZN( u0_u2_n541 ) , .A1( u0_u2_n731 ) , .A2( u0_u2_n795 ) );
  NOR2_X1 u0_u2_U325 (.ZN( u0_u2_n638 ) , .A1( u0_u2_n731 ) , .A2( u0_u2_n820 ) );
  NOR2_X1 u0_u2_U326 (.ZN( u0_u2_n540 ) , .A2( u0_u2_n731 ) , .A1( u0_u2_n737 ) );
  INV_X1 u0_u2_U327 (.A( u0_u2_n731 ) , .ZN( u0_u2_n863 ) );
  NOR2_X1 u0_u2_U328 (.ZN( u0_u2_n455 ) , .A1( u0_u2_n854 ) , .A2( w3_5 ) );
  NOR2_X1 u0_u2_U329 (.ZN( u0_u2_n448 ) , .A2( w3_4 ) , .A1( w3_5 ) );
  NOR4_X1 u0_u2_U33 (.A4( u0_u2_n694 ) , .A3( u0_u2_n695 ) , .A2( u0_u2_n696 ) , .A1( u0_u2_n697 ) , .ZN( u0_u2_n698 ) );
  INV_X1 u0_u2_U330 (.ZN( u0_u2_n855 ) , .A( w3_5 ) );
  AOI21_X1 u0_u2_U331 (.A( u0_u2_n446 ) , .ZN( u0_u2_n648 ) , .B1( u0_u2_n687 ) , .B2( u0_u2_n824 ) );
  AOI21_X1 u0_u2_U332 (.B2( u0_u2_n446 ) , .A( u0_u2_n797 ) , .B1( u0_u2_n799 ) , .ZN( u0_u2_n800 ) );
  OAI22_X1 u0_u2_U333 (.B1( u0_u2_n446 ) , .ZN( u0_u2_n702 ) , .A2( u0_u2_n737 ) , .A1( u0_u2_n787 ) , .B2( u0_u2_n824 ) );
  AOI21_X1 u0_u2_U334 (.B2( u0_u2_n446 ) , .ZN( u0_u2_n504 ) , .A( u0_u2_n786 ) , .B1( u0_u2_n811 ) );
  AOI21_X1 u0_u2_U335 (.B2( u0_u2_n446 ) , .ZN( u0_u2_n571 ) , .B1( u0_u2_n731 ) , .A( u0_u2_n786 ) );
  AOI21_X1 u0_u2_U336 (.ZN( u0_u2_n450 ) , .B1( u0_u2_n796 ) , .B2( u0_u2_n798 ) , .A( u0_u2_n821 ) );
  NOR2_X1 u0_u2_U337 (.ZN( u0_u2_n671 ) , .A1( u0_u2_n792 ) , .A2( u0_u2_n798 ) );
  NOR2_X1 u0_u2_U338 (.ZN( u0_u2_n562 ) , .A1( u0_u2_n757 ) , .A2( u0_u2_n798 ) );
  NOR2_X1 u0_u2_U339 (.ZN( u0_u2_n566 ) , .A2( u0_u2_n798 ) , .A1( u0_u2_n810 ) );
  AOI221_X1 u0_u2_U34 (.A( u0_u2_n688 ) , .ZN( u0_u2_n699 ) , .B2( u0_u2_n847 ) , .C1( u0_u2_n849 ) , .C2( u0_u2_n869 ) , .B1( u0_u2_n872 ) );
  NAND2_X2 u0_u2_U340 (.A1( u0_u2_n462 ) , .A2( u0_u2_n469 ) , .ZN( u0_u2_n757 ) );
  NOR2_X1 u0_u2_U341 (.ZN( u0_u2_n649 ) , .A2( u0_u2_n795 ) , .A1( u0_u2_n798 ) );
  NOR2_X1 u0_u2_U342 (.ZN( u0_u2_n691 ) , .A1( u0_u2_n798 ) , .A2( u0_u2_n820 ) );
  NOR2_X1 u0_u2_U343 (.ZN( u0_u2_n549 ) , .A1( u0_u2_n769 ) , .A2( u0_u2_n798 ) );
  INV_X1 u0_u2_U344 (.A( u0_u2_n798 ) , .ZN( u0_u2_n880 ) );
  AOI21_X1 u0_u2_U345 (.B2( u0_u2_n442 ) , .ZN( u0_u2_n517 ) , .A( u0_u2_n737 ) , .B1( u0_u2_n822 ) );
  AOI21_X1 u0_u2_U346 (.B1( u0_u2_n446 ) , .ZN( u0_u2_n633 ) , .B2( u0_u2_n676 ) , .A( u0_u2_n797 ) );
  INV_X1 u0_u2_U347 (.A( u0_u2_n676 ) , .ZN( u0_u2_n872 ) );
  NOR2_X1 u0_u2_U348 (.A1( u0_u2_n442 ) , .ZN( u0_u2_n773 ) , .A2( u0_u2_n820 ) );
  NOR2_X1 u0_u2_U349 (.A1( u0_u2_n442 ) , .ZN( u0_u2_n659 ) , .A2( u0_u2_n821 ) );
  NOR2_X1 u0_u2_U35 (.A1( u0_u2_n685 ) , .ZN( u0_u2_n700 ) , .A2( u0_u2_n814 ) );
  AOI21_X1 u0_u2_U350 (.A( u0_u2_n442 ) , .ZN( u0_u2_n484 ) , .B1( u0_u2_n757 ) , .B2( u0_u2_n813 ) );
  NOR2_X1 u0_u2_U351 (.A1( u0_u2_n442 ) , .ZN( u0_u2_n534 ) , .A2( u0_u2_n786 ) );
  NOR2_X1 u0_u2_U352 (.A1( u0_u2_n442 ) , .ZN( u0_u2_n609 ) , .A2( u0_u2_n810 ) );
  NOR2_X1 u0_u2_U353 (.A2( u0_u2_n442 ) , .ZN( u0_u2_n635 ) , .A1( u0_u2_n792 ) );
  NOR2_X1 u0_u2_U354 (.ZN( u0_u2_n588 ) , .A1( u0_u2_n676 ) , .A2( u0_u2_n795 ) );
  OAI22_X1 u0_u2_U355 (.ZN( u0_u2_n644 ) , .A1( u0_u2_n706 ) , .B2( u0_u2_n735 ) , .A2( u0_u2_n769 ) , .B1( u0_u2_n823 ) );
  AOI21_X1 u0_u2_U356 (.ZN( u0_u2_n506 ) , .B1( u0_u2_n687 ) , .A( u0_u2_n819 ) , .B2( u0_u2_n823 ) );
  OAI22_X1 u0_u2_U357 (.A1( u0_u2_n731 ) , .ZN( u0_u2_n733 ) , .B2( u0_u2_n757 ) , .B1( u0_u2_n819 ) , .A2( u0_u2_n823 ) );
  AOI21_X1 u0_u2_U358 (.A( u0_u2_n443 ) , .B2( u0_u2_n823 ) , .B1( u0_u2_n824 ) , .ZN( u0_u2_n825 ) );
  OAI22_X1 u0_u2_U359 (.B1( u0_u2_n442 ) , .A1( u0_u2_n443 ) , .ZN( u0_u2_n631 ) , .B2( u0_u2_n754 ) , .A2( u0_u2_n823 ) );
  NOR2_X1 u0_u2_U36 (.ZN( u0_u2_n552 ) , .A1( u0_u2_n756 ) , .A2( u0_u2_n821 ) );
  NOR2_X1 u0_u2_U360 (.ZN( u0_u2_n606 ) , .A2( u0_u2_n798 ) , .A1( u0_u2_n823 ) );
  NOR2_X1 u0_u2_U361 (.ZN( u0_u2_n538 ) , .A2( u0_u2_n787 ) , .A1( u0_u2_n823 ) );
  NOR2_X1 u0_u2_U362 (.ZN( u0_u2_n526 ) , .A2( u0_u2_n706 ) , .A1( u0_u2_n823 ) );
  NOR2_X1 u0_u2_U363 (.A1( u0_u2_n442 ) , .ZN( u0_u2_n695 ) , .A2( u0_u2_n823 ) );
  NOR2_X1 u0_u2_U364 (.ZN( u0_u2_n565 ) , .A1( u0_u2_n715 ) , .A2( u0_u2_n823 ) );
  NOR2_X1 u0_u2_U365 (.ZN( u0_u2_n692 ) , .A1( u0_u2_n736 ) , .A2( u0_u2_n823 ) );
  NAND2_X1 u0_u2_U366 (.ZN( u0_u2_n678 ) , .A1( u0_u2_n813 ) , .A2( u0_u2_n823 ) );
  NOR2_X1 u0_u2_U367 (.ZN( u0_u2_n469 ) , .A2( w3_0 ) , .A1( w3_1 ) );
  NOR2_X1 u0_u2_U368 (.ZN( u0_u2_n461 ) , .A1( u0_u2_n834 ) , .A2( w3_0 ) );
  INV_X1 u0_u2_U369 (.ZN( u0_u2_n833 ) , .A( w3_0 ) );
  NOR2_X1 u0_u2_U37 (.ZN( u0_u2_n502 ) , .A1( u0_u2_n685 ) , .A2( u0_u2_n701 ) );
  INV_X1 u0_u2_U370 (.A( u0_u2_n819 ) , .ZN( u0_u2_n861 ) );
  INV_X1 u0_u2_U371 (.A( u0_u2_n823 ) , .ZN( u0_u2_n838 ) );
  INV_X1 u0_u2_U372 (.A( u0_u2_n810 ) , .ZN( u0_u2_n850 ) );
  INV_X1 u0_u2_U373 (.ZN( u0_u2_n854 ) , .A( w3_4 ) );
  INV_X1 u0_u2_U374 (.A( u0_u2_n441 ) , .ZN( u0_u2_n845 ) );
  NOR2_X1 u0_u2_U375 (.A1( u0_u2_n704 ) , .ZN( u0_u2_n777 ) , .A2( u0_u2_n822 ) );
  AOI21_X1 u0_u2_U376 (.B2( u0_u2_n441 ) , .ZN( u0_u2_n578 ) , .B1( u0_u2_n813 ) , .A( u0_u2_n819 ) );
  NOR2_X1 u0_u2_U377 (.ZN( u0_u2_n639 ) , .A2( u0_u2_n704 ) , .A1( u0_u2_n731 ) );
  NOR2_X1 u0_u2_U378 (.A2( u0_u2_n441 ) , .A1( u0_u2_n787 ) , .ZN( u0_u2_n827 ) );
  AOI21_X1 u0_u2_U379 (.B2( u0_u2_n441 ) , .ZN( u0_u2_n485 ) , .A( u0_u2_n756 ) , .B1( u0_u2_n786 ) );
  INV_X1 u0_u2_U38 (.A( u0_u2_n821 ) , .ZN( u0_u2_n840 ) );
  NOR2_X1 u0_u2_U380 (.A2( u0_u2_n441 ) , .ZN( u0_u2_n573 ) , .A1( u0_u2_n770 ) );
  NOR2_X1 u0_u2_U381 (.ZN( u0_u2_n669 ) , .A2( u0_u2_n704 ) , .A1( u0_u2_n736 ) );
  NOR2_X1 u0_u2_U382 (.A2( u0_u2_n441 ) , .ZN( u0_u2_n723 ) , .A1( u0_u2_n799 ) );
  NOR2_X1 u0_u2_U383 (.A2( u0_u2_n441 ) , .ZN( u0_u2_n601 ) , .A1( u0_u2_n735 ) );
  NOR2_X1 u0_u2_U384 (.A2( u0_u2_n441 ) , .ZN( u0_u2_n548 ) , .A1( u0_u2_n706 ) );
  NOR2_X1 u0_u2_U385 (.ZN( u0_u2_n587 ) , .A2( u0_u2_n704 ) , .A1( u0_u2_n798 ) );
  NOR2_X1 u0_u2_U386 (.ZN( u0_u2_n479 ) , .A2( w3_2 ) , .A1( w3_3 ) );
  NOR2_X1 u0_u2_U387 (.ZN( u0_u2_n462 ) , .A1( u0_u2_n835 ) , .A2( w3_3 ) );
  INV_X1 u0_u2_U388 (.ZN( u0_u2_n836 ) , .A( w3_3 ) );
  AOI21_X1 u0_u2_U389 (.ZN( u0_u2_n583 ) , .B2( u0_u2_n731 ) , .B1( u0_u2_n755 ) , .A( u0_u2_n792 ) );
  NAND4_X1 u0_u2_U39 (.A4( u0_u2_n664 ) , .A3( u0_u2_n665 ) , .A2( u0_u2_n666 ) , .A1( u0_u2_n667 ) , .ZN( u0_u2_n807 ) );
  OAI222_X1 u0_u2_U390 (.B2( u0_u2_n754 ) , .B1( u0_u2_n755 ) , .A2( u0_u2_n756 ) , .ZN( u0_u2_n764 ) , .C2( u0_u2_n812 ) , .C1( u0_u2_n821 ) , .A1( u0_u2_n824 ) );
  OAI21_X1 u0_u2_U391 (.A( u0_u2_n738 ) , .B1( u0_u2_n739 ) , .ZN( u0_u2_n743 ) , .B2( u0_u2_n812 ) );
  OAI22_X1 u0_u2_U392 (.B2( u0_u2_n810 ) , .B1( u0_u2_n811 ) , .A2( u0_u2_n812 ) , .A1( u0_u2_n813 ) , .ZN( u0_u2_n815 ) );
  OAI222_X1 u0_u2_U393 (.C2( u0_u2_n444 ) , .ZN( u0_u2_n512 ) , .B2( u0_u2_n654 ) , .B1( u0_u2_n754 ) , .A2( u0_u2_n755 ) , .C1( u0_u2_n812 ) , .A1( u0_u2_n813 ) );
  AOI21_X1 u0_u2_U394 (.ZN( u0_u2_n657 ) , .A( u0_u2_n786 ) , .B1( u0_u2_n799 ) , .B2( u0_u2_n812 ) );
  INV_X1 u0_u2_U395 (.A( u0_u2_n812 ) , .ZN( u0_u2_n867 ) );
  NOR2_X1 u0_u2_U396 (.ZN( u0_u2_n742 ) , .A2( u0_u2_n810 ) , .A1( u0_u2_n812 ) );
  NOR2_X1 u0_u2_U397 (.ZN( u0_u2_n491 ) , .A1( u0_u2_n795 ) , .A2( u0_u2_n812 ) );
  NOR2_X1 u0_u2_U398 (.ZN( u0_u2_n574 ) , .A1( u0_u2_n754 ) , .A2( u0_u2_n812 ) );
  AOI21_X1 u0_u2_U399 (.A( u0_u2_n441 ) , .B1( u0_u2_n442 ) , .ZN( u0_u2_n559 ) , .B2( u0_u2_n812 ) );
  NOR3_X1 u0_u2_U4 (.A3( u0_u2_n807 ) , .A2( u0_u2_n808 ) , .A1( u0_u2_n809 ) , .ZN( u0_u2_n832 ) );
  NOR3_X1 u0_u2_U40 (.A3( u0_u2_n661 ) , .A2( u0_u2_n662 ) , .A1( u0_u2_n663 ) , .ZN( u0_u2_n664 ) );
  NAND2_X1 u0_u2_U400 (.ZN( u0_u2_n760 ) , .A1( u0_u2_n770 ) , .A2( u0_u2_n812 ) );
  NOR2_X1 u0_u2_U401 (.ZN( u0_u2_n722 ) , .A1( u0_u2_n812 ) , .A2( u0_u2_n824 ) );
  NOR2_X1 u0_u2_U402 (.ZN( u0_u2_n563 ) , .A1( u0_u2_n769 ) , .A2( u0_u2_n812 ) );
  NOR2_X1 u0_u2_U403 (.ZN( u0_u2_n677 ) , .A1( u0_u2_n797 ) , .A2( u0_u2_n812 ) );
  NAND4_X1 u0_u2_U404 (.ZN( u0_subword_11 ) , .A4( u0_u2_n711 ) , .A3( u0_u2_n712 ) , .A2( u0_u2_n713 ) , .A1( u0_u2_n714 ) );
  INV_X1 u0_u2_U405 (.A( u0_u2_n713 ) , .ZN( u0_u2_n883 ) );
  OAI22_X1 u0_u2_U406 (.B2( u0_u2_n751 ) , .ZN( u0_u2_n753 ) , .A2( u0_u2_n769 ) , .B1( u0_u2_n787 ) , .A1( u0_u2_n799 ) );
  OAI22_X1 u0_u2_U407 (.B1( u0_u2_n446 ) , .ZN( u0_u2_n503 ) , .A2( u0_u2_n751 ) , .A1( u0_u2_n787 ) , .B2( u0_u2_n813 ) );
  NOR2_X1 u0_u2_U408 (.ZN( u0_u2_n523 ) , .A1( u0_u2_n715 ) , .A2( u0_u2_n751 ) );
  OAI22_X1 u0_u2_U409 (.ZN( u0_u2_n717 ) , .A2( u0_u2_n735 ) , .B2( u0_u2_n736 ) , .A1( u0_u2_n751 ) , .B1( u0_u2_n820 ) );
  NOR3_X1 u0_u2_U41 (.A3( u0_u2_n655 ) , .A2( u0_u2_n656 ) , .A1( u0_u2_n657 ) , .ZN( u0_u2_n666 ) );
  NOR2_X1 u0_u2_U410 (.A2( u0_u2_n751 ) , .ZN( u0_u2_n776 ) , .A1( u0_u2_n819 ) );
  OAI22_X1 u0_u2_U411 (.B1( u0_u2_n447 ) , .ZN( u0_u2_n451 ) , .A2( u0_u2_n735 ) , .A1( u0_u2_n751 ) , .B2( u0_u2_n756 ) );
  NOR2_X1 u0_u2_U412 (.ZN( u0_u2_n554 ) , .A1( u0_u2_n706 ) , .A2( u0_u2_n751 ) );
  NOR2_X1 u0_u2_U413 (.ZN( u0_u2_n537 ) , .A2( u0_u2_n751 ) , .A1( u0_u2_n799 ) );
  NOR2_X1 u0_u2_U414 (.A2( u0_u2_n751 ) , .ZN( u0_u2_n762 ) , .A1( u0_u2_n812 ) );
  NOR2_X1 u0_u2_U415 (.A1( u0_u2_n442 ) , .ZN( u0_u2_n680 ) , .A2( u0_u2_n751 ) );
  NOR2_X1 u0_u2_U416 (.ZN( u0_u2_n725 ) , .A2( u0_u2_n731 ) , .A1( u0_u2_n751 ) );
  NOR2_X1 u0_u2_U417 (.ZN( u0_u2_n589 ) , .A1( u0_u2_n751 ) , .A2( u0_u2_n822 ) );
  INV_X1 u0_u2_U418 (.A( u0_u2_n751 ) , .ZN( u0_u2_n844 ) );
  NAND4_X1 u0_u2_U419 (.ZN( u0_subword_10 ) , .A4( u0_u2_n650 ) , .A3( u0_u2_n651 ) , .A2( u0_u2_n652 ) , .A1( u0_u2_n653 ) );
  NOR3_X1 u0_u2_U42 (.A3( u0_u2_n658 ) , .A2( u0_u2_n659 ) , .A1( u0_u2_n660 ) , .ZN( u0_u2_n665 ) );
  OAI22_X1 u0_u2_U420 (.ZN( u0_u2_n595 ) , .A2( u0_u2_n754 ) , .B2( u0_u2_n769 ) , .A1( u0_u2_n770 ) , .B1( u0_u2_n791 ) );
  NAND2_X1 u0_u2_U421 (.A1( u0_u2_n736 ) , .A2( u0_u2_n791 ) , .ZN( u0_u2_n818 ) );
  AOI21_X1 u0_u2_U422 (.ZN( u0_u2_n599 ) , .B1( u0_u2_n735 ) , .B2( u0_u2_n791 ) , .A( u0_u2_n797 ) );
  AOI21_X1 u0_u2_U423 (.ZN( u0_u2_n655 ) , .A( u0_u2_n769 ) , .B2( u0_u2_n791 ) , .B1( u0_u2_n799 ) );
  AOI21_X1 u0_u2_U424 (.ZN( u0_u2_n630 ) , .B1( u0_u2_n706 ) , .A( u0_u2_n786 ) , .B2( u0_u2_n791 ) );
  OAI22_X1 u0_u2_U425 (.ZN( u0_u2_n688 ) , .A1( u0_u2_n706 ) , .A2( u0_u2_n737 ) , .B2( u0_u2_n791 ) , .B1( u0_u2_n824 ) );
  OAI21_X1 u0_u2_U426 (.A( u0_u2_n620 ) , .ZN( u0_u2_n623 ) , .B1( u0_u2_n632 ) , .B2( u0_u2_n791 ) );
  NOR2_X1 u0_u2_U427 (.ZN( u0_u2_n658 ) , .A1( u0_u2_n791 ) , .A2( u0_u2_n795 ) );
  NOR2_X1 u0_u2_U428 (.ZN( u0_u2_n617 ) , .A1( u0_u2_n791 ) , .A2( u0_u2_n823 ) );
  NOR2_X1 u0_u2_U429 (.ZN( u0_u2_n560 ) , .A2( u0_u2_n751 ) , .A1( u0_u2_n791 ) );
  NAND4_X1 u0_u2_U43 (.A4( u0_u2_n567 ) , .A3( u0_u2_n568 ) , .A2( u0_u2_n569 ) , .A1( u0_u2_n570 ) , .ZN( u0_u2_n614 ) );
  NOR2_X1 u0_u2_U430 (.A2( u0_u2_n441 ) , .ZN( u0_u2_n607 ) , .A1( u0_u2_n791 ) );
  INV_X1 u0_u2_U431 (.A( u0_u2_n791 ) , .ZN( u0_u2_n868 ) );
  AOI21_X1 u0_u2_U432 (.ZN( u0_u2_n507 ) , .A( u0_u2_n704 ) , .B1( u0_u2_n715 ) , .B2( u0_u2_n793 ) );
  OAI22_X1 u0_u2_U433 (.ZN( u0_u2_n597 ) , .B1( u0_u2_n737 ) , .B2( u0_u2_n756 ) , .A2( u0_u2_n793 ) , .A1( u0_u2_n810 ) );
  AOI222_X1 u0_u2_U434 (.ZN( u0_u2_n520 ) , .C1( u0_u2_n839 ) , .B2( u0_u2_n844 ) , .A2( u0_u2_n850 ) , .C2( u0_u2_n869 ) , .B1( u0_u2_n870 ) , .A1( u0_u2_n873 ) );
  AOI222_X1 u0_u2_U435 (.ZN( u0_u2_n612 ) , .B2( u0_u2_n678 ) , .B1( u0_u2_n760 ) , .C2( u0_u2_n838 ) , .A1( u0_u2_n840 ) , .A2( u0_u2_n869 ) , .C1( u0_u2_n870 ) );
  AOI221_X1 u0_u2_U436 (.A( u0_u2_n490 ) , .ZN( u0_u2_n495 ) , .B1( u0_u2_n838 ) , .C2( u0_u2_n851 ) , .C1( u0_u2_n859 ) , .B2( u0_u2_n869 ) );
  NAND3_X1 u0_u2_U437 (.ZN( u0_subword_14 ) , .A3( u0_u2_n804 ) , .A2( u0_u2_n805 ) , .A1( u0_u2_n806 ) );
  NAND3_X1 u0_u2_U438 (.ZN( u0_subword_13 ) , .A3( u0_u2_n765 ) , .A2( u0_u2_n766 ) , .A1( u0_u2_n767 ) );
  NAND3_X1 u0_u2_U439 (.ZN( u0_subword_12 ) , .A3( u0_u2_n745 ) , .A2( u0_u2_n746 ) , .A1( u0_u2_n747 ) );
  NOR4_X1 u0_u2_U44 (.ZN( u0_u2_n568 ) , .A1( u0_u2_n660 ) , .A3( u0_u2_n668 ) , .A4( u0_u2_n692 ) , .A2( u0_u2_n775 ) );
  NAND3_X1 u0_u2_U440 (.A3( u0_u2_n682 ) , .A2( u0_u2_n683 ) , .A1( u0_u2_n684 ) , .ZN( u0_u2_n814 ) );
  NAND3_X1 u0_u2_U441 (.ZN( u0_u2_n645 ) , .A3( u0_u2_n715 ) , .A2( u0_u2_n731 ) , .A1( u0_u2_n799 ) );
  NAND3_X1 u0_u2_U442 (.A3( u0_u2_n625 ) , .A2( u0_u2_n626 ) , .A1( u0_u2_n627 ) , .ZN( u0_u2_n732 ) );
  NAND3_X1 u0_u2_U443 (.A3( u0_u2_n592 ) , .A2( u0_u2_n593 ) , .A1( u0_u2_n594 ) , .ZN( u0_u2_n628 ) );
  NAND3_X1 u0_u2_U444 (.ZN( u0_u2_n572 ) , .A3( u0_u2_n687 ) , .A2( u0_u2_n757 ) , .A1( u0_u2_n792 ) );
  NAND3_X1 u0_u2_U445 (.A3( u0_u2_n530 ) , .A2( u0_u2_n531 ) , .A1( u0_u2_n532 ) , .ZN( u0_u2_n749 ) );
  NAND3_X1 u0_u2_U446 (.A3( u0_u2_n519 ) , .A1( u0_u2_n520 ) , .ZN( u0_u2_n615 ) , .A2( u0_u2_n878 ) );
  NAND3_X1 u0_u2_U447 (.A3( u0_u2_n474 ) , .A2( u0_u2_n475 ) , .A1( u0_u2_n476 ) , .ZN( u0_u2_n784 ) );
  NOR2_X1 u0_u2_U448 (.ZN( u0_u2_n660 ) , .A1( u0_u2_n769 ) , .A2( u0_u2_n793 ) );
  NAND2_X1 u0_u2_U449 (.A2( u0_u2_n756 ) , .A1( u0_u2_n793 ) , .ZN( u0_u2_n816 ) );
  NOR4_X1 u0_u2_U45 (.A4( u0_u2_n559 ) , .A3( u0_u2_n560 ) , .A2( u0_u2_n561 ) , .A1( u0_u2_n562 ) , .ZN( u0_u2_n569 ) );
  NOR2_X1 u0_u2_U450 (.ZN( u0_u2_n561 ) , .A1( u0_u2_n793 ) , .A2( u0_u2_n820 ) );
  NOR2_X1 u0_u2_U451 (.ZN( u0_u2_n619 ) , .A1( u0_u2_n786 ) , .A2( u0_u2_n793 ) );
  NOR2_X1 u0_u2_U452 (.ZN( u0_u2_n724 ) , .A2( u0_u2_n751 ) , .A1( u0_u2_n793 ) );
  NOR2_X1 u0_u2_U453 (.ZN( u0_u2_n796 ) , .A2( u0_u2_n869 ) , .A1( u0_u2_n875 ) );
  NOR2_X1 u0_u2_U454 (.ZN( u0_u2_n708 ) , .A2( u0_u2_n793 ) , .A1( u0_u2_n824 ) );
  NOR2_X1 u0_u2_U455 (.A1( u0_u2_n737 ) , .ZN( u0_u2_n772 ) , .A2( u0_u2_n793 ) );
  INV_X1 u0_u2_U456 (.A( u0_u2_n793 ) , .ZN( u0_u2_n869 ) );
  NOR4_X1 u0_u2_U46 (.A4( u0_u2_n563 ) , .A3( u0_u2_n564 ) , .A2( u0_u2_n565 ) , .A1( u0_u2_n566 ) , .ZN( u0_u2_n567 ) );
  NOR4_X1 u0_u2_U47 (.A4( u0_u2_n516 ) , .A2( u0_u2_n517 ) , .A1( u0_u2_n518 ) , .ZN( u0_u2_n519 ) , .A3( u0_u2_n677 ) );
  INV_X1 u0_u2_U48 (.A( u0_u2_n512 ) , .ZN( u0_u2_n878 ) );
  NOR4_X1 u0_u2_U49 (.A4( u0_u2_n668 ) , .A3( u0_u2_n669 ) , .A2( u0_u2_n670 ) , .A1( u0_u2_n671 ) , .ZN( u0_u2_n684 ) );
  NOR3_X1 u0_u2_U5 (.ZN( u0_u2_n605 ) , .A1( u0_u2_n615 ) , .A3( u0_u2_n730 ) , .A2( u0_u2_n749 ) );
  NOR4_X1 u0_u2_U50 (.A4( u0_u2_n672 ) , .A3( u0_u2_n673 ) , .A2( u0_u2_n674 ) , .A1( u0_u2_n675 ) , .ZN( u0_u2_n683 ) );
  NOR2_X1 u0_u2_U51 (.ZN( u0_u2_n811 ) , .A1( u0_u2_n861 ) , .A2( u0_u2_n868 ) );
  NOR4_X1 u0_u2_U52 (.A1( u0_u2_n473 ) , .ZN( u0_u2_n474 ) , .A4( u0_u2_n549 ) , .A2( u0_u2_n561 ) , .A3( u0_u2_n621 ) );
  NAND4_X1 u0_u2_U53 (.A4( u0_u2_n492 ) , .A3( u0_u2_n493 ) , .A2( u0_u2_n494 ) , .A1( u0_u2_n495 ) , .ZN( u0_u2_n785 ) );
  NOR4_X1 u0_u2_U54 (.ZN( u0_u2_n492 ) , .A2( u0_u2_n540 ) , .A1( u0_u2_n565 ) , .A3( u0_u2_n638 ) , .A4( u0_u2_n725 ) );
  NOR4_X1 u0_u2_U55 (.A4( u0_u2_n521 ) , .A3( u0_u2_n522 ) , .A2( u0_u2_n523 ) , .A1( u0_u2_n524 ) , .ZN( u0_u2_n531 ) );
  NOR4_X1 u0_u2_U56 (.A3( u0_u2_n528 ) , .A1( u0_u2_n529 ) , .ZN( u0_u2_n530 ) , .A2( u0_u2_n680 ) , .A4( u0_u2_n776 ) );
  NOR2_X1 u0_u2_U57 (.ZN( u0_u2_n768 ) , .A1( u0_u2_n840 ) , .A2( u0_u2_n841 ) );
  NAND4_X1 u0_u2_U58 (.A4( u0_u2_n779 ) , .A3( u0_u2_n780 ) , .A2( u0_u2_n781 ) , .A1( u0_u2_n782 ) , .ZN( u0_u2_n808 ) );
  NOR3_X1 u0_u2_U59 (.A3( u0_u2_n772 ) , .A2( u0_u2_n773 ) , .A1( u0_u2_n774 ) , .ZN( u0_u2_n780 ) );
  NOR3_X1 u0_u2_U6 (.ZN( u0_u2_n511 ) , .A2( u0_u2_n686 ) , .A3( u0_u2_n784 ) , .A1( u0_u2_n883 ) );
  NOR4_X1 u0_u2_U60 (.A4( u0_u2_n775 ) , .A3( u0_u2_n776 ) , .A2( u0_u2_n777 ) , .A1( u0_u2_n778 ) , .ZN( u0_u2_n779 ) );
  AOI222_X1 u0_u2_U61 (.ZN( u0_u2_n782 ) , .A1( u0_u2_n837 ) , .C1( u0_u2_n841 ) , .B2( u0_u2_n848 ) , .A2( u0_u2_n857 ) , .B1( u0_u2_n868 ) , .C2( u0_u2_n880 ) );
  NAND4_X1 u0_u2_U62 (.A4( u0_u2_n480 ) , .A3( u0_u2_n481 ) , .A2( u0_u2_n482 ) , .A1( u0_u2_n483 ) , .ZN( u0_u2_n685 ) );
  NOR4_X1 u0_u2_U63 (.A4( u0_u2_n477 ) , .ZN( u0_u2_n483 ) , .A3( u0_u2_n563 ) , .A1( u0_u2_n742 ) , .A2( u0_u2_n762 ) );
  NOR4_X1 u0_u2_U64 (.ZN( u0_u2_n480 ) , .A2( u0_u2_n528 ) , .A4( u0_u2_n601 ) , .A1( u0_u2_n616 ) , .A3( u0_u2_n636 ) );
  NOR4_X1 u0_u2_U65 (.ZN( u0_u2_n481 ) , .A1( u0_u2_n513 ) , .A3( u0_u2_n551 ) , .A2( u0_u2_n590 ) , .A4( u0_u2_n723 ) );
  NAND4_X1 u0_u2_U66 (.A4( u0_u2_n463 ) , .A3( u0_u2_n464 ) , .A2( u0_u2_n465 ) , .A1( u0_u2_n466 ) , .ZN( u0_u2_n686 ) );
  NOR3_X1 u0_u2_U67 (.ZN( u0_u2_n464 ) , .A3( u0_u2_n537 ) , .A1( u0_u2_n562 ) , .A2( u0_u2_n577 ) );
  NOR4_X1 u0_u2_U68 (.ZN( u0_u2_n463 ) , .A2( u0_u2_n524 ) , .A1( u0_u2_n550 ) , .A3( u0_u2_n586 ) , .A4( u0_u2_n622 ) );
  NOR4_X1 u0_u2_U69 (.ZN( u0_u2_n465 ) , .A2( u0_u2_n516 ) , .A1( u0_u2_n606 ) , .A4( u0_u2_n635 ) , .A3( u0_u2_n718 ) );
  NOR3_X1 u0_u2_U7 (.A2( u0_u2_n614 ) , .A1( u0_u2_n615 ) , .ZN( u0_u2_n653 ) , .A3( u0_u2_n729 ) );
  NAND4_X1 u0_u2_U70 (.A4( u0_u2_n580 ) , .A3( u0_u2_n581 ) , .A1( u0_u2_n582 ) , .ZN( u0_u2_n730 ) , .A2( u0_u2_n881 ) );
  NOR4_X1 u0_u2_U71 (.A4( u0_u2_n576 ) , .A3( u0_u2_n577 ) , .A2( u0_u2_n578 ) , .A1( u0_u2_n579 ) , .ZN( u0_u2_n580 ) );
  AOI221_X1 u0_u2_U72 (.A( u0_u2_n571 ) , .C2( u0_u2_n572 ) , .ZN( u0_u2_n581 ) , .B2( u0_u2_n852 ) , .B1( u0_u2_n859 ) , .C1( u0_u2_n860 ) );
  INV_X1 u0_u2_U73 (.A( u0_u2_n614 ) , .ZN( u0_u2_n881 ) );
  NOR4_X1 u0_u2_U74 (.A4( u0_u2_n636 ) , .A3( u0_u2_n637 ) , .A2( u0_u2_n638 ) , .A1( u0_u2_n639 ) , .ZN( u0_u2_n640 ) );
  AOI211_X1 u0_u2_U75 (.B( u0_u2_n630 ) , .A( u0_u2_n631 ) , .ZN( u0_u2_n642 ) , .C2( u0_u2_n843 ) , .C1( u0_u2_n870 ) );
  NOR4_X1 u0_u2_U76 (.A4( u0_u2_n633 ) , .A3( u0_u2_n634 ) , .A2( u0_u2_n635 ) , .ZN( u0_u2_n641 ) , .A1( u0_u2_n671 ) );
  NAND4_X1 u0_u2_U77 (.A4( u0_u2_n542 ) , .A3( u0_u2_n543 ) , .A2( u0_u2_n544 ) , .A1( u0_u2_n545 ) , .ZN( u0_u2_n629 ) );
  NOR4_X1 u0_u2_U78 (.A4( u0_u2_n533 ) , .A2( u0_u2_n534 ) , .A1( u0_u2_n535 ) , .ZN( u0_u2_n545 ) , .A3( u0_u2_n708 ) );
  NOR4_X1 u0_u2_U79 (.A1( u0_u2_n538 ) , .ZN( u0_u2_n543 ) , .A2( u0_u2_n661 ) , .A4( u0_u2_n675 ) , .A3( u0_u2_n772 ) );
  NOR3_X1 u0_u2_U8 (.A3( u0_u2_n729 ) , .A1( u0_u2_n730 ) , .ZN( u0_u2_n747 ) , .A2( u0_u2_n748 ) );
  NOR4_X1 u0_u2_U80 (.A4( u0_u2_n536 ) , .A3( u0_u2_n537 ) , .ZN( u0_u2_n544 ) , .A2( u0_u2_n691 ) , .A1( u0_u2_n801 ) );
  NOR2_X1 u0_u2_U81 (.ZN( u0_u2_n755 ) , .A1( u0_u2_n868 ) , .A2( u0_u2_n869 ) );
  NAND4_X1 u0_u2_U82 (.A4( u0_u2_n555 ) , .A3( u0_u2_n556 ) , .A2( u0_u2_n557 ) , .A1( u0_u2_n558 ) , .ZN( u0_u2_n752 ) );
  NOR3_X1 u0_u2_U83 (.ZN( u0_u2_n556 ) , .A2( u0_u2_n658 ) , .A1( u0_u2_n674 ) , .A3( u0_u2_n778 ) );
  AOI211_X1 u0_u2_U84 (.B( u0_u2_n546 ) , .A( u0_u2_n547 ) , .ZN( u0_u2_n558 ) , .C2( u0_u2_n846 ) , .C1( u0_u2_n858 ) );
  NOR4_X1 u0_u2_U85 (.A4( u0_u2_n548 ) , .A3( u0_u2_n549 ) , .A2( u0_u2_n550 ) , .ZN( u0_u2_n557 ) , .A1( u0_u2_n695 ) );
  NOR4_X1 u0_u2_U86 (.A4( u0_u2_n616 ) , .A3( u0_u2_n617 ) , .A2( u0_u2_n618 ) , .A1( u0_u2_n619 ) , .ZN( u0_u2_n626 ) );
  NOR4_X1 u0_u2_U87 (.ZN( u0_u2_n627 ) , .A1( u0_u2_n663 ) , .A3( u0_u2_n673 ) , .A4( u0_u2_n689 ) , .A2( u0_u2_n773 ) );
  NOR2_X1 u0_u2_U88 (.ZN( u0_u2_n654 ) , .A1( u0_u2_n861 ) , .A2( u0_u2_n875 ) );
  INV_X1 u0_u2_U89 (.A( u0_u2_n813 ) , .ZN( u0_u2_n848 ) );
  NOR2_X1 u0_u2_U9 (.ZN( u0_u2_n582 ) , .A1( u0_u2_n629 ) , .A2( u0_u2_n752 ) );
  NAND4_X1 u0_u2_U90 (.A4( u0_u2_n726 ) , .A3( u0_u2_n727 ) , .A2( u0_u2_n728 ) , .ZN( u0_u2_n748 ) , .A1( u0_u2_n864 ) );
  NOR4_X1 u0_u2_U91 (.A4( u0_u2_n722 ) , .A3( u0_u2_n723 ) , .A2( u0_u2_n724 ) , .A1( u0_u2_n725 ) , .ZN( u0_u2_n726 ) );
  AOI221_X1 u0_u2_U92 (.A( u0_u2_n717 ) , .ZN( u0_u2_n728 ) , .C2( u0_u2_n851 ) , .B2( u0_u2_n852 ) , .C1( u0_u2_n868 ) , .B1( u0_u2_n869 ) );
  INV_X1 u0_u2_U93 (.A( u0_u2_n716 ) , .ZN( u0_u2_n864 ) );
  INV_X1 u0_u2_U94 (.A( u0_u2_n769 ) , .ZN( u0_u2_n837 ) );
  NAND2_X1 u0_u2_U95 (.A2( u0_u2_n769 ) , .A1( u0_u2_n813 ) , .ZN( u0_u2_n817 ) );
  OAI21_X1 u0_u2_U96 (.ZN( u0_u2_n738 ) , .A( u0_u2_n840 ) , .B2( u0_u2_n859 ) , .B1( u0_u2_n880 ) );
  OR4_X1 u0_u2_U97 (.A4( u0_u2_n525 ) , .A2( u0_u2_n526 ) , .A1( u0_u2_n527 ) , .ZN( u0_u2_n529 ) , .A3( u0_u2_n828 ) );
  OR4_X1 u0_u2_U98 (.A4( u0_u2_n573 ) , .A3( u0_u2_n574 ) , .A2( u0_u2_n575 ) , .ZN( u0_u2_n579 ) , .A1( u0_u2_n672 ) );
  OR4_X1 u0_u2_U99 (.A4( u0_u2_n689 ) , .A3( u0_u2_n690 ) , .A2( u0_u2_n691 ) , .A1( u0_u2_n692 ) , .ZN( u0_u2_n697 ) );
  NOR2_X1 u0_u3_U10 (.ZN( u0_u3_n578 ) , .A1( u0_u3_n625 ) , .A2( u0_u3_n748 ) );
  NOR2_X1 u0_u3_U100 (.ZN( u0_u3_n669 ) , .A1( u0_u3_n731 ) , .A2( u0_u3_n806 ) );
  NOR2_X1 u0_u3_U101 (.ZN( u0_u3_n535 ) , .A2( u0_u3_n752 ) , .A1( u0_u3_n753 ) );
  NOR2_X1 u0_u3_U102 (.A2( u0_u3_n711 ) , .A1( u0_u3_n765 ) , .ZN( u0_u3_n797 ) );
  OAI22_X1 u0_u3_U103 (.B1( u0_u3_n493 ) , .ZN( u0_u3_n494 ) , .A1( u0_u3_n689 ) , .A2( u0_u3_n766 ) , .B2( u0_u3_n820 ) );
  NOR3_X1 u0_u3_U104 (.ZN( u0_u3_n493 ) , .A1( u0_u3_n785 ) , .A2( u0_u3_n852 ) , .A3( u0_u3_n865 ) );
  NOR2_X1 u0_u3_U105 (.ZN( u0_u3_n509 ) , .A2( u0_u3_n731 ) , .A1( u0_u3_n765 ) );
  NOR2_X1 u0_u3_U106 (.ZN( u0_u3_n520 ) , .A1( u0_u3_n711 ) , .A2( u0_u3_n806 ) );
  OAI21_X1 u0_u3_U107 (.ZN( u0_u3_n734 ) , .A( u0_u3_n836 ) , .B2( u0_u3_n854 ) , .B1( u0_u3_n875 ) );
  NOR2_X1 u0_u3_U108 (.ZN( u0_u3_n604 ) , .A2( u0_u3_n783 ) , .A1( u0_u3_n806 ) );
  NOR2_X1 u0_u3_U109 (.A2( u0_u3_n711 ) , .A1( u0_u3_n753 ) , .ZN( u0_u3_n774 ) );
  NOR2_X1 u0_u3_U11 (.A1( u0_u3_n681 ) , .ZN( u0_u3_n696 ) , .A2( u0_u3_n810 ) );
  NOR2_X1 u0_u3_U110 (.A2( u0_u3_n438 ) , .ZN( u0_u3_n670 ) , .A1( u0_u3_n753 ) );
  BUF_X2 u0_u3_U111 (.Z( u0_u3_n439 ) , .A( u0_u3_n794 ) );
  OAI21_X1 u0_u3_U112 (.ZN( u0_u3_n790 ) , .A( u0_u3_n841 ) , .B1( u0_u3_n865 ) , .B2( u0_u3_n875 ) );
  BUF_X2 u0_u3_U113 (.Z( u0_u3_n41 ) , .A( u0_u3_n700 ) );
  NOR2_X1 u0_u3_U114 (.ZN( u0_u3_n632 ) , .A2( u0_u3_n731 ) , .A1( u0_u3_n788 ) );
  NOR2_X1 u0_u3_U115 (.ZN( u0_u3_n512 ) , .A1( u0_u3_n732 ) , .A2( u0_u3_n782 ) );
  NOR2_X1 u0_u3_U116 (.ZN( u0_u3_n510 ) , .A1( u0_u3_n815 ) , .A2( u0_u3_n820 ) );
  NOR2_X1 u0_u3_U117 (.ZN( u0_u3_n666 ) , .A1( u0_u3_n732 ) , .A2( u0_u3_n788 ) );
  NOR2_X1 u0_u3_U118 (.ZN( u0_u3_n546 ) , .A2( u0_u3_n711 ) , .A1( u0_u3_n788 ) );
  NOR2_X1 u0_u3_U119 (.ZN( u0_u3_n511 ) , .A2( u0_u3_n783 ) , .A1( u0_u3_n788 ) );
  INV_X1 u0_u3_U12 (.A( u0_u3_n683 ) , .ZN( u0_u3_n842 ) );
  NOR2_X1 u0_u3_U120 (.ZN( u0_u3_n547 ) , .A2( u0_u3_n788 ) , .A1( u0_u3_n795 ) );
  NOR2_X1 u0_u3_U121 (.ZN( u0_u3_n685 ) , .A2( u0_u3_n711 ) , .A1( u0_u3_n820 ) );
  AOI21_X1 u0_u3_U122 (.ZN( u0_u3_n572 ) , .B1( u0_u3_n753 ) , .B2( u0_u3_n765 ) , .A( u0_u3_n783 ) );
  NOR2_X1 u0_u3_U123 (.ZN( u0_u3_n714 ) , .A1( u0_u3_n765 ) , .A2( u0_u3_n766 ) );
  NOR2_X1 u0_u3_U124 (.ZN( u0_u3_n532 ) , .A1( u0_u3_n711 ) , .A2( u0_u3_n782 ) );
  AOI21_X1 u0_u3_U125 (.ZN( u0_u3_n518 ) , .A( u0_u3_n732 ) , .B1( u0_u3_n753 ) , .B2( u0_u3_n806 ) );
  NOR2_X1 u0_u3_U126 (.ZN( u0_u3_n617 ) , .A1( u0_u3_n765 ) , .A2( u0_u3_n815 ) );
  INV_X1 u0_u3_U127 (.A( u0_u3_n753 ) , .ZN( u0_u3_n844 ) );
  AOI21_X1 u0_u3_U128 (.ZN( u0_u3_n594 ) , .B2( u0_u3_n766 ) , .A( u0_u3_n788 ) , .B1( u0_u3_n815 ) );
  AOI21_X1 u0_u3_U129 (.ZN( u0_u3_n517 ) , .A( u0_u3_n782 ) , .B2( u0_u3_n795 ) , .B1( u0_u3_n815 ) );
  INV_X1 u0_u3_U13 (.A( u0_u3_n650 ) , .ZN( u0_u3_n872 ) );
  AOI21_X1 u0_u3_U130 (.B1( u0_u3_n689 ) , .ZN( u0_u3_n690 ) , .A( u0_u3_n731 ) , .B2( u0_u3_n764 ) );
  INV_X1 u0_u3_U131 (.A( u0_u3_n731 ) , .ZN( u0_u3_n854 ) );
  NOR2_X1 u0_u3_U132 (.ZN( u0_u3_n571 ) , .A1( u0_u3_n732 ) , .A2( u0_u3_n765 ) );
  INV_X1 u0_u3_U133 (.A( u0_u3_n795 ) , .ZN( u0_u3_n853 ) );
  NOR2_X1 u0_u3_U134 (.A1( u0_u3_n752 ) , .ZN( u0_u3_n770 ) , .A2( u0_u3_n806 ) );
  NOR2_X1 u0_u3_U135 (.A2( u0_u3_n438 ) , .ZN( u0_u3_n618 ) , .A1( u0_u3_n788 ) );
  AOI211_X1 u0_u3_U136 (.C2( u0_u3_n440 ) , .B( u0_u3_n626 ) , .A( u0_u3_n627 ) , .ZN( u0_u3_n638 ) , .C1( u0_u3_n865 ) );
  NOR4_X1 u0_u3_U137 (.A4( u0_u3_n632 ) , .A3( u0_u3_n633 ) , .A2( u0_u3_n634 ) , .A1( u0_u3_n635 ) , .ZN( u0_u3_n636 ) );
  NOR4_X1 u0_u3_U138 (.A4( u0_u3_n629 ) , .A3( u0_u3_n630 ) , .A2( u0_u3_n631 ) , .ZN( u0_u3_n637 ) , .A1( u0_u3_n667 ) );
  INV_X1 u0_u3_U139 (.A( u0_u3_n783 ) , .ZN( u0_u3_n852 ) );
  NOR4_X1 u0_u3_U14 (.A4( u0_u3_n547 ) , .A3( u0_u3_n548 ) , .A2( u0_u3_n549 ) , .A1( u0_u3_n550 ) , .ZN( u0_u3_n551 ) );
  OAI21_X1 u0_u3_U140 (.A( u0_u3_n701 ) , .ZN( u0_u3_n705 ) , .B2( u0_u3_n753 ) , .B1( u0_u3_n807 ) );
  OAI21_X1 u0_u3_U141 (.ZN( u0_u3_n701 ) , .B2( u0_u3_n836 ) , .B1( u0_u3_n840 ) , .A( u0_u3_n862 ) );
  INV_X1 u0_u3_U142 (.A( u0_u3_n732 ) , .ZN( u0_u3_n870 ) );
  NOR2_X1 u0_u3_U143 (.A2( u0_u3_n440 ) , .ZN( u0_u3_n628 ) , .A1( u0_u3_n841 ) );
  INV_X1 u0_u3_U144 (.A( u0_u3_n766 ) , .ZN( u0_u3_n868 ) );
  NOR2_X1 u0_u3_U145 (.ZN( u0_u3_n473 ) , .A2( u0_u3_n782 ) , .A1( u0_u3_n818 ) );
  INV_X1 u0_u3_U146 (.A( u0_u3_n440 ) , .ZN( u0_u3_n816 ) );
  INV_X1 u0_u3_U147 (.A( u0_u3_n820 ) , .ZN( u0_u3_n846 ) );
  NAND2_X1 u0_u3_U148 (.ZN( u0_u3_n717 ) , .A1( u0_u3_n731 ) , .A2( u0_u3_n783 ) );
  INV_X1 u0_u3_U149 (.A( u0_u3_n788 ) , .ZN( u0_u3_n848 ) );
  NOR4_X1 u0_u3_U15 (.A4( u0_u3_n448 ) , .A3( u0_u3_n449 ) , .A2( u0_u3_n519 ) , .A1( u0_u3_n544 ) , .ZN( u0_u3_n709 ) );
  AOI221_X1 u0_u3_U150 (.A( u0_u3_n767 ) , .ZN( u0_u3_n777 ) , .C2( u0_u3_n813 ) , .B2( u0_u3_n838 ) , .C1( u0_u3_n857 ) , .B1( u0_u3_n868 ) );
  INV_X1 u0_u3_U151 (.A( u0_u3_n764 ) , .ZN( u0_u3_n838 ) );
  AND2_X1 u0_u3_U152 (.ZN( u0_u3_n735 ) , .A1( u0_u3_n782 ) , .A2( u0_u3_n788 ) );
  AOI221_X1 u0_u3_U153 (.A( u0_u3_n453 ) , .ZN( u0_u3_n462 ) , .C2( u0_u3_n756 ) , .B1( u0_u3_n835 ) , .C1( u0_u3_n844 ) , .B2( u0_u3_n863 ) );
  AOI21_X1 u0_u3_U154 (.ZN( u0_u3_n453 ) , .B2( u0_u3_n795 ) , .A( u0_u3_n806 ) , .B1( u0_u3_n818 ) );
  AOI211_X1 u0_u3_U155 (.A( u0_u3_n591 ) , .ZN( u0_u3_n600 ) , .B( u0_u3_n624 ) , .C1( u0_u3_n847 ) , .C2( u0_u3_n857 ) );
  OAI221_X1 u0_u3_U156 (.A( u0_u3_n730 ) , .C2( u0_u3_n731 ) , .B2( u0_u3_n732 ) , .B1( u0_u3_n733 ) , .ZN( u0_u3_n740 ) , .C1( u0_u3_n820 ) );
  NAND2_X1 u0_u3_U157 (.A1( u0_u3_n444 ) , .A2( u0_u3_n467 ) , .ZN( u0_u3_n711 ) );
  NAND2_X1 u0_u3_U158 (.A2( u0_u3_n474 ) , .A1( u0_u3_n475 ) , .ZN( u0_u3_n820 ) );
  NAND2_X1 u0_u3_U159 (.A2( u0_u3_n463 ) , .A1( u0_u3_n468 ) , .ZN( u0_u3_n783 ) );
  OR3_X1 u0_u3_U16 (.ZN( u0_u3_n449 ) , .A1( u0_u3_n531 ) , .A3( u0_u3_n580 ) , .A2( u0_u3_n877 ) );
  NAND2_X1 u0_u3_U160 (.A1( u0_u3_n458 ) , .A2( u0_u3_n474 ) , .ZN( u0_u3_n806 ) );
  NAND2_X1 u0_u3_U161 (.A2( u0_u3_n451 ) , .A1( u0_u3_n463 ) , .ZN( u0_u3_n731 ) );
  NAND2_X1 u0_u3_U162 (.A1( u0_u3_n452 ) , .A2( u0_u3_n467 ) , .ZN( u0_u3_n727 ) );
  NAND2_X1 u0_u3_U163 (.A2( u0_u3_n457 ) , .A1( u0_u3_n475 ) , .ZN( u0_u3_n782 ) );
  NOR2_X1 u0_u3_U164 (.ZN( u0_u3_n456 ) , .A1( u0_u3_n829 ) , .A2( u0_u3_n830 ) );
  NAND2_X1 u0_u3_U165 (.A2( u0_u3_n467 ) , .A1( u0_u3_n468 ) , .ZN( u0_u3_n815 ) );
  NAND2_X1 u0_u3_U166 (.A2( u0_u3_n451 ) , .A1( u0_u3_n455 ) , .ZN( u0_u3_n732 ) );
  NAND2_X1 u0_u3_U167 (.A2( u0_u3_n452 ) , .A1( u0_u3_n455 ) , .ZN( u0_u3_n766 ) );
  NAND2_X1 u0_u3_U168 (.A1( u0_u3_n454 ) , .A2( u0_u3_n474 ) , .ZN( u0_u3_n819 ) );
  NAND2_X1 u0_u3_U169 (.A1( u0_u3_n456 ) , .A2( u0_u3_n464 ) , .ZN( u0_u3_n747 ) );
  OR4_X1 u0_u3_U17 (.A4( u0_u3_n445 ) , .A2( u0_u3_n446 ) , .A1( u0_u3_n447 ) , .ZN( u0_u3_n448 ) , .A3( u0_u3_n556 ) );
  NAND2_X1 u0_u3_U170 (.A2( u0_u3_n444 ) , .A1( u0_u3_n450 ) , .ZN( u0_u3_n787 ) );
  NAND2_X1 u0_u3_U171 (.A1( u0_u3_n454 ) , .A2( u0_u3_n457 ) , .ZN( u0_u3_n817 ) );
  NAND2_X1 u0_u3_U172 (.A1( u0_u3_n450 ) , .A2( u0_u3_n452 ) , .ZN( u0_u3_n808 ) );
  NAND2_X1 u0_u3_U173 (.A2( u0_u3_n456 ) , .A1( u0_u3_n458 ) , .ZN( u0_u3_n809 ) );
  NAND2_X1 u0_u3_U174 (.A1( u0_u3_n450 ) , .A2( u0_u3_n451 ) , .ZN( u0_u3_n789 ) );
  NAND2_X1 u0_u3_U175 (.A2( u0_u3_n464 ) , .A1( u0_u3_n465 ) , .ZN( u0_u3_n750 ) );
  NAND2_X1 u0_u3_U176 (.A1( u0_u3_n465 ) , .A2( u0_u3_n475 ) , .ZN( u0_u3_n791 ) );
  NAND2_X1 u0_u3_U177 (.A2( u0_u3_n457 ) , .A1( u0_u3_n458 ) , .ZN( u0_u3_n733 ) );
  NAND2_X1 u0_u3_U178 (.A1( u0_u3_n454 ) , .A2( u0_u3_n465 ) , .ZN( u0_u3_n793 ) );
  AND2_X1 u0_u3_U179 (.ZN( u0_u3_n440 ) , .A1( u0_u3_n457 ) , .A2( u0_u3_n464 ) );
  INV_X1 u0_u3_U18 (.A( u0_u3_n616 ) , .ZN( u0_u3_n877 ) );
  NOR2_X1 u0_u3_U180 (.ZN( u0_u3_n452 ) , .A1( u0_u3_n850 ) , .A2( w3_28 ) );
  NAND4_X1 u0_u3_U181 (.ZN( u0_subword_1 ) , .A4( u0_u3_n598 ) , .A3( u0_u3_n599 ) , .A2( u0_u3_n600 ) , .A1( u0_u3_n601 ) );
  AOI211_X1 u0_u3_U182 (.B( u0_u3_n592 ) , .A( u0_u3_n593 ) , .ZN( u0_u3_n599 ) , .C2( u0_u3_n814 ) , .C1( u0_u3_n836 ) );
  NOR4_X1 u0_u3_U183 (.A4( u0_u3_n594 ) , .A3( u0_u3_n595 ) , .A2( u0_u3_n596 ) , .A1( u0_u3_n597 ) , .ZN( u0_u3_n598 ) );
  NOR4_X1 u0_u3_U184 (.A4( u0_u3_n737 ) , .A3( u0_u3_n738 ) , .A2( u0_u3_n739 ) , .A1( u0_u3_n740 ) , .ZN( u0_u3_n741 ) );
  AOI211_X1 u0_u3_U185 (.B( u0_u3_n728 ) , .A( u0_u3_n729 ) , .ZN( u0_u3_n742 ) , .C1( u0_u3_n845 ) , .C2( u0_u3_n857 ) );
  AOI222_X1 u0_u3_U186 (.B2( u0_u3_n641 ) , .ZN( u0_u3_n647 ) , .B1( u0_u3_n843 ) , .A1( u0_u3_n844 ) , .C2( u0_u3_n848 ) , .C1( u0_u3_n865 ) , .A2( u0_u3_n867 ) );
  NOR4_X1 u0_u3_U187 (.A4( u0_u3_n642 ) , .A3( u0_u3_n643 ) , .A2( u0_u3_n644 ) , .A1( u0_u3_n645 ) , .ZN( u0_u3_n646 ) );
  AOI221_X1 u0_u3_U188 (.A( u0_u3_n784 ) , .ZN( u0_u3_n801 ) , .C2( u0_u3_n839 ) , .B2( u0_u3_n840 ) , .B1( u0_u3_n867 ) , .C1( u0_u3_n868 ) );
  NOR4_X1 u0_u3_U189 (.A4( u0_u3_n796 ) , .A3( u0_u3_n797 ) , .A2( u0_u3_n798 ) , .A1( u0_u3_n799 ) , .ZN( u0_u3_n800 ) );
  NOR4_X1 u0_u3_U19 (.ZN( u0_u3_n478 ) , .A1( u0_u3_n534 ) , .A3( u0_u3_n571 ) , .A4( u0_u3_n603 ) , .A2( u0_u3_n645 ) );
  NAND4_X1 u0_u3_U190 (.ZN( u0_subword_0 ) , .A4( u0_u3_n504 ) , .A3( u0_u3_n505 ) , .A2( u0_u3_n506 ) , .A1( u0_u3_n507 ) );
  NOR4_X1 u0_u3_U191 (.A4( u0_u3_n501 ) , .A3( u0_u3_n502 ) , .A2( u0_u3_n503 ) , .ZN( u0_u3_n504 ) , .A1( u0_u3_n530 ) );
  AOI221_X1 u0_u3_U192 (.A( u0_u3_n500 ) , .ZN( u0_u3_n505 ) , .B2( u0_u3_n845 ) , .C1( u0_u3_n848 ) , .C2( u0_u3_n862 ) , .B1( u0_u3_n864 ) );
  NOR4_X1 u0_u3_U193 (.A4( u0_u3_n703 ) , .A3( u0_u3_n704 ) , .A2( u0_u3_n705 ) , .A1( u0_u3_n706 ) , .ZN( u0_u3_n707 ) );
  NOR4_X1 u0_u3_U194 (.A3( u0_u3_n758 ) , .A2( u0_u3_n759 ) , .A1( u0_u3_n760 ) , .ZN( u0_u3_n761 ) , .A4( u0_u3_n871 ) );
  AOI211_X1 u0_u3_U195 (.B( u0_u3_n748 ) , .A( u0_u3_n749 ) , .ZN( u0_u3_n762 ) , .C1( u0_u3_n835 ) , .C2( u0_u3_n855 ) );
  NAND4_X1 u0_u3_U196 (.ZN( u0_subword_7 ) , .A4( u0_u3_n825 ) , .A3( u0_u3_n826 ) , .A2( u0_u3_n827 ) , .A1( u0_u3_n828 ) );
  NOR4_X1 u0_u3_U197 (.A4( u0_u3_n821 ) , .A3( u0_u3_n822 ) , .A2( u0_u3_n823 ) , .A1( u0_u3_n824 ) , .ZN( u0_u3_n825 ) );
  NAND2_X1 u0_u3_U198 (.A2( u0_u3_n464 ) , .A1( u0_u3_n474 ) , .ZN( u0_u3_n700 ) );
  NAND2_X1 u0_u3_U199 (.A2( u0_u3_n451 ) , .A1( u0_u3_n467 ) , .ZN( u0_u3_n818 ) );
  INV_X1 u0_u3_U20 (.A( u0_u3_n752 ) , .ZN( u0_u3_n865 ) );
  OAI21_X1 u0_u3_U200 (.B1( u0_u3_n756 ) , .ZN( u0_u3_n757 ) , .A( u0_u3_n847 ) , .B2( u0_u3_n870 ) );
  AOI221_X1 u0_u3_U201 (.A( u0_u3_n567 ) , .C2( u0_u3_n568 ) , .ZN( u0_u3_n577 ) , .B2( u0_u3_n847 ) , .B1( u0_u3_n854 ) , .C1( u0_u3_n855 ) );
  AOI222_X1 u0_u3_U202 (.ZN( u0_u3_n663 ) , .A2( u0_u3_n841 ) , .B1( u0_u3_n843 ) , .C2( u0_u3_n847 ) , .A1( u0_u3_n862 ) , .C1( u0_u3_n865 ) , .B2( u0_u3_n872 ) );
  AOI221_X1 u0_u3_U203 (.A( u0_u3_n713 ) , .ZN( u0_u3_n724 ) , .C2( u0_u3_n846 ) , .B2( u0_u3_n847 ) , .C1( u0_u3_n863 ) , .B1( u0_u3_n864 ) );
  NAND4_X1 u0_u3_U204 (.A4( u0_u3_n538 ) , .A3( u0_u3_n539 ) , .A2( u0_u3_n540 ) , .A1( u0_u3_n541 ) , .ZN( u0_u3_n625 ) );
  NOR4_X1 u0_u3_U205 (.A1( u0_u3_n534 ) , .ZN( u0_u3_n539 ) , .A2( u0_u3_n657 ) , .A4( u0_u3_n671 ) , .A3( u0_u3_n768 ) );
  NAND4_X1 u0_u3_U206 (.A4( u0_u3_n496 ) , .A3( u0_u3_n497 ) , .A1( u0_u3_n498 ) , .ZN( u0_u3_n805 ) , .A2( u0_u3_n869 ) );
  NOR4_X1 u0_u3_U207 (.A2( u0_u3_n494 ) , .A1( u0_u3_n495 ) , .ZN( u0_u3_n496 ) , .A3( u0_u3_n583 ) , .A4( u0_u3_n615 ) );
  NAND2_X1 u0_u3_U208 (.A1( u0_u3_n444 ) , .A2( u0_u3_n463 ) , .ZN( u0_u3_n702 ) );
  NAND2_X1 u0_u3_U209 (.A1( u0_u3_n455 ) , .A2( u0_u3_n468 ) , .ZN( u0_u3_n672 ) );
  AOI222_X1 u0_u3_U21 (.ZN( u0_u3_n566 ) , .B1( u0_u3_n833 ) , .C1( u0_u3_n843 ) , .A2( u0_u3_n845 ) , .A1( u0_u3_n856 ) , .B2( u0_u3_n865 ) , .C2( u0_u3_n875 ) );
  NAND4_X1 u0_u3_U210 (.A4( u0_u3_n563 ) , .A3( u0_u3_n564 ) , .A2( u0_u3_n565 ) , .A1( u0_u3_n566 ) , .ZN( u0_u3_n610 ) );
  NOR4_X1 u0_u3_U211 (.ZN( u0_u3_n564 ) , .A1( u0_u3_n656 ) , .A3( u0_u3_n664 ) , .A4( u0_u3_n688 ) , .A2( u0_u3_n771 ) );
  NOR2_X1 u0_u3_U212 (.ZN( u0_u3_n454 ) , .A1( u0_u3_n831 ) , .A2( u0_u3_n832 ) );
  INV_X1 u0_u3_U213 (.ZN( u0_u3_n831 ) , .A( w3_26 ) );
  NOR2_X1 u0_u3_U214 (.ZN( u0_u3_n710 ) , .A2( u0_u3_n779 ) , .A1( u0_u3_n803 ) );
  OAI21_X1 u0_u3_U215 (.A( u0_u3_n734 ) , .B1( u0_u3_n735 ) , .ZN( u0_u3_n739 ) , .B2( u0_u3_n808 ) );
  AOI21_X1 u0_u3_U216 (.ZN( u0_u3_n653 ) , .A( u0_u3_n782 ) , .B1( u0_u3_n795 ) , .B2( u0_u3_n808 ) );
  INV_X1 u0_u3_U217 (.A( u0_u3_n808 ) , .ZN( u0_u3_n862 ) );
  NOR2_X1 u0_u3_U218 (.ZN( u0_u3_n738 ) , .A2( u0_u3_n806 ) , .A1( u0_u3_n808 ) );
  NAND2_X1 u0_u3_U219 (.ZN( u0_u3_n756 ) , .A1( u0_u3_n766 ) , .A2( u0_u3_n808 ) );
  NOR4_X1 u0_u3_U22 (.ZN( u0_u3_n482 ) , .A1( u0_u3_n523 ) , .A4( u0_u3_n560 ) , .A3( u0_u3_n585 ) , .A2( u0_u3_n633 ) );
  NOR2_X1 u0_u3_U220 (.ZN( u0_u3_n559 ) , .A1( u0_u3_n765 ) , .A2( u0_u3_n808 ) );
  OAI221_X1 u0_u3_U221 (.A( u0_u3_n699 ) , .ZN( u0_u3_n706 ) , .C2( u0_u3_n787 ) , .C1( u0_u3_n788 ) , .B1( u0_u3_n789 ) , .B2( u0_u3_n809 ) );
  OAI222_X1 u0_u3_U222 (.B1( u0_u3_n41 ) , .ZN( u0_u3_n620 ) , .C1( u0_u3_n727 ) , .C2( u0_u3_n750 ) , .B2( u0_u3_n789 ) , .A2( u0_u3_n795 ) , .A1( u0_u3_n819 ) );
  NAND2_X1 u0_u3_U223 (.A2( u0_u3_n444 ) , .A1( u0_u3_n455 ) , .ZN( u0_u3_n794 ) );
  OAI222_X1 u0_u3_U224 (.B2( u0_u3_n711 ) , .ZN( u0_u3_n712 ) , .C2( u0_u3_n727 ) , .B1( u0_u3_n750 ) , .A1( u0_u3_n809 ) , .C1( u0_u3_n817 ) , .A2( u0_u3_n818 ) );
  INV_X1 u0_u3_U225 (.A( u0_u3_n675 ) , .ZN( u0_u3_n861 ) );
  NOR2_X1 u0_u3_U226 (.ZN( u0_u3_n531 ) , .A2( u0_u3_n727 ) , .A1( u0_u3_n806 ) );
  NOR2_X1 u0_u3_U227 (.ZN( u0_u3_n529 ) , .A1( u0_u3_n727 ) , .A2( u0_u3_n753 ) );
  INV_X1 u0_u3_U228 (.A( u0_u3_n727 ) , .ZN( u0_u3_n858 ) );
  NOR2_X1 u0_u3_U229 (.ZN( u0_u3_n450 ) , .A2( u0_u3_n851 ) , .A1( u0_u3_n860 ) );
  NOR4_X1 u0_u3_U23 (.A4( u0_u3_n559 ) , .A3( u0_u3_n560 ) , .A2( u0_u3_n561 ) , .A1( u0_u3_n562 ) , .ZN( u0_u3_n563 ) );
  AOI222_X1 u0_u3_U230 (.ZN( u0_u3_n528 ) , .A1( u0_u3_n837 ) , .B2( u0_u3_n839 ) , .C1( u0_u3_n846 ) , .C2( u0_u3_n852 ) , .A2( u0_u3_n854 ) , .B1( u0_u3_n868 ) );
  NOR3_X1 u0_u3_U231 (.A2( u0_u3_n440 ) , .ZN( u0_u3_n443 ) , .A3( u0_u3_n839 ) , .A1( u0_u3_n848 ) );
  NAND2_X1 u0_u3_U232 (.ZN( u0_u3_n616 ) , .A2( u0_u3_n839 ) , .A1( u0_u3_n875 ) );
  NOR2_X1 u0_u3_U233 (.ZN( u0_u3_n498 ) , .A1( u0_u3_n681 ) , .A2( u0_u3_n697 ) );
  AOI211_X1 u0_u3_U234 (.B( u0_u3_n697 ) , .A( u0_u3_n698 ) , .ZN( u0_u3_n708 ) , .C2( u0_u3_n834 ) , .C1( u0_u3_n853 ) );
  NOR2_X1 u0_u3_U235 (.ZN( u0_u3_n586 ) , .A1( u0_u3_n795 ) , .A2( u0_u3_n820 ) );
  AOI21_X1 u0_u3_U236 (.ZN( u0_u3_n543 ) , .A( u0_u3_n766 ) , .B2( u0_u3_n782 ) , .B1( u0_u3_n820 ) );
  NOR2_X1 u0_u3_U237 (.ZN( u0_u3_n612 ) , .A2( u0_u3_n727 ) , .A1( u0_u3_n820 ) );
  NOR2_X1 u0_u3_U238 (.ZN( u0_u3_n718 ) , .A1( u0_u3_n808 ) , .A2( u0_u3_n820 ) );
  OAI21_X1 u0_u3_U239 (.A( u0_u3_n790 ) , .B2( u0_u3_n791 ) , .B1( u0_u3_n792 ) , .ZN( u0_u3_n798 ) );
  NOR4_X1 u0_u3_U24 (.A4( u0_u3_n555 ) , .A3( u0_u3_n556 ) , .A2( u0_u3_n557 ) , .A1( u0_u3_n558 ) , .ZN( u0_u3_n565 ) );
  AOI21_X1 u0_u3_U240 (.ZN( u0_u3_n642 ) , .B2( u0_u3_n752 ) , .A( u0_u3_n791 ) , .B1( u0_u3_n815 ) );
  AOI21_X1 u0_u3_U241 (.A( u0_u3_n736 ) , .ZN( u0_u3_n737 ) , .B2( u0_u3_n783 ) , .B1( u0_u3_n795 ) );
  AOI21_X1 u0_u3_U242 (.B2( u0_u3_n766 ) , .ZN( u0_u3_n767 ) , .A( u0_u3_n791 ) , .B1( u0_u3_n795 ) );
  NOR2_X1 u0_u3_U243 (.ZN( u0_u3_n521 ) , .A1( u0_u3_n711 ) , .A2( u0_u3_n791 ) );
  NOR2_X1 u0_u3_U244 (.ZN( u0_u3_n487 ) , .A1( u0_u3_n791 ) , .A2( u0_u3_n808 ) );
  NOR2_X1 u0_u3_U245 (.ZN( u0_u3_n537 ) , .A1( u0_u3_n727 ) , .A2( u0_u3_n791 ) );
  INV_X1 u0_u3_U246 (.A( u0_u3_n791 ) , .ZN( u0_u3_n847 ) );
  OAI22_X1 u0_u3_U247 (.B2( u0_u3_n782 ) , .B1( u0_u3_n783 ) , .ZN( u0_u3_n784 ) , .A2( u0_u3_n817 ) , .A1( u0_u3_n818 ) );
  AOI21_X1 u0_u3_U248 (.ZN( u0_u3_n501 ) , .A( u0_u3_n727 ) , .B2( u0_u3_n765 ) , .B1( u0_u3_n817 ) );
  NAND4_X1 u0_u3_U249 (.A4( u0_u3_n482 ) , .A3( u0_u3_n483 ) , .A2( u0_u3_n484 ) , .A1( u0_u3_n485 ) , .ZN( u0_u3_n697 ) );
  NOR4_X1 u0_u3_U25 (.A4( u0_u3_n771 ) , .A3( u0_u3_n772 ) , .A2( u0_u3_n773 ) , .A1( u0_u3_n774 ) , .ZN( u0_u3_n775 ) );
  AOI21_X1 u0_u3_U250 (.ZN( u0_u3_n542 ) , .B2( u0_u3_n815 ) , .A( u0_u3_n817 ) , .B1( u0_u3_n818 ) );
  NOR2_X1 u0_u3_U251 (.ZN( u0_u3_n523 ) , .A2( u0_u3_n711 ) , .A1( u0_u3_n817 ) );
  NOR2_X1 u0_u3_U252 (.ZN( u0_u3_n549 ) , .A2( u0_u3_n783 ) , .A1( u0_u3_n817 ) );
  INV_X1 u0_u3_U253 (.A( u0_u3_n817 ) , .ZN( u0_u3_n836 ) );
  NOR2_X1 u0_u3_U254 (.ZN( u0_u3_n548 ) , .A1( u0_u3_n752 ) , .A2( u0_u3_n817 ) );
  NOR2_X1 u0_u3_U255 (.ZN( u0_u3_n560 ) , .A1( u0_u3_n795 ) , .A2( u0_u3_n817 ) );
  AOI21_X1 u0_u3_U256 (.A( u0_u3_n673 ) , .B1( u0_u3_n674 ) , .ZN( u0_u3_n675 ) , .B2( u0_u3_n858 ) );
  AOI22_X1 u0_u3_U257 (.A2( u0_u3_n785 ) , .ZN( u0_u3_n786 ) , .B2( u0_u3_n834 ) , .A1( u0_u3_n837 ) , .B1( u0_u3_n865 ) );
  AOI21_X1 u0_u3_U258 (.ZN( u0_u3_n643 ) , .B2( u0_u3_n750 ) , .A( u0_u3_n795 ) , .B1( u0_u3_n806 ) );
  NAND4_X1 u0_u3_U259 (.A4( u0_u3_n775 ) , .A3( u0_u3_n776 ) , .A2( u0_u3_n777 ) , .A1( u0_u3_n778 ) , .ZN( u0_u3_n804 ) );
  NOR3_X1 u0_u3_U26 (.A3( u0_u3_n768 ) , .A2( u0_u3_n769 ) , .A1( u0_u3_n770 ) , .ZN( u0_u3_n776 ) );
  OAI21_X1 u0_u3_U260 (.ZN( u0_u3_n466 ) , .B1( u0_u3_n812 ) , .A( u0_u3_n837 ) , .B2( u0_u3_n853 ) );
  NOR2_X1 u0_u3_U261 (.ZN( u0_u3_n659 ) , .A1( u0_u3_n750 ) , .A2( u0_u3_n783 ) );
  NOR2_X1 u0_u3_U262 (.ZN( u0_u3_n683 ) , .A2( u0_u3_n837 ) , .A1( u0_u3_n841 ) );
  NOR2_X1 u0_u3_U263 (.ZN( u0_u3_n764 ) , .A1( u0_u3_n836 ) , .A2( u0_u3_n837 ) );
  NOR2_X1 u0_u3_U264 (.ZN( u0_u3_n570 ) , .A1( u0_u3_n750 ) , .A2( u0_u3_n808 ) );
  NOR2_X1 u0_u3_U265 (.A2( u0_u3_n438 ) , .ZN( u0_u3_n633 ) , .A1( u0_u3_n750 ) );
  INV_X1 u0_u3_U266 (.A( u0_u3_n750 ) , .ZN( u0_u3_n837 ) );
  NOR4_X1 u0_u3_U267 (.ZN( u0_u3_n488 ) , .A2( u0_u3_n536 ) , .A1( u0_u3_n561 ) , .A3( u0_u3_n634 ) , .A4( u0_u3_n721 ) );
  NAND4_X1 u0_u3_U268 (.A4( u0_u3_n488 ) , .A3( u0_u3_n489 ) , .A2( u0_u3_n490 ) , .A1( u0_u3_n491 ) , .ZN( u0_u3_n781 ) );
  AOI21_X1 u0_u3_U269 (.B1( u0_u3_n438 ) , .ZN( u0_u3_n592 ) , .B2( u0_u3_n702 ) , .A( u0_u3_n820 ) );
  NAND4_X1 u0_u3_U27 (.A4( u0_u3_n606 ) , .A3( u0_u3_n607 ) , .A2( u0_u3_n608 ) , .A1( u0_u3_n609 ) , .ZN( u0_u3_n725 ) );
  AOI21_X1 u0_u3_U270 (.B1( u0_u3_n702 ) , .ZN( u0_u3_n703 ) , .A( u0_u3_n735 ) , .B2( u0_u3_n766 ) );
  INV_X1 u0_u3_U271 (.A( u0_u3_n702 ) , .ZN( u0_u3_n855 ) );
  AOI21_X1 u0_u3_U272 (.ZN( u0_u3_n445 ) , .A( u0_u3_n702 ) , .B1( u0_u3_n736 ) , .B2( u0_u3_n753 ) );
  NOR2_X1 u0_u3_U273 (.ZN( u0_u3_n686 ) , .A2( u0_u3_n702 ) , .A1( u0_u3_n806 ) );
  NOR2_X1 u0_u3_U274 (.ZN( u0_u3_n580 ) , .A2( u0_u3_n702 ) , .A1( u0_u3_n817 ) );
  NAND2_X1 u0_u3_U275 (.A1( u0_u3_n702 ) , .A2( u0_u3_n732 ) , .ZN( u0_u3_n785 ) );
  NOR3_X1 u0_u3_U276 (.A3( u0_u3_n744 ) , .A2( u0_u3_n745 ) , .A1( u0_u3_n746 ) , .ZN( u0_u3_n763 ) );
  OAI22_X1 u0_u3_U277 (.ZN( u0_u3_n492 ) , .A1( u0_u3_n727 ) , .B2( u0_u3_n731 ) , .B1( u0_u3_n733 ) , .A2( u0_u3_n782 ) );
  NOR2_X1 u0_u3_U278 (.ZN( u0_u3_n582 ) , .A2( u0_u3_n711 ) , .A1( u0_u3_n733 ) );
  NOR2_X1 u0_u3_U279 (.ZN( u0_u3_n536 ) , .A2( u0_u3_n727 ) , .A1( u0_u3_n733 ) );
  NOR3_X1 u0_u3_U28 (.A1( u0_u3_n602 ) , .ZN( u0_u3_n607 ) , .A3( u0_u3_n666 ) , .A2( u0_u3_n773 ) );
  AOI222_X1 u0_u3_U280 (.ZN( u0_u3_n608 ) , .B2( u0_u3_n674 ) , .B1( u0_u3_n756 ) , .C2( u0_u3_n834 ) , .A1( u0_u3_n836 ) , .A2( u0_u3_n864 ) , .C1( u0_u3_n865 ) );
  AOI221_X1 u0_u3_U281 (.A( u0_u3_n486 ) , .ZN( u0_u3_n491 ) , .B1( u0_u3_n834 ) , .C2( u0_u3_n846 ) , .C1( u0_u3_n854 ) , .B2( u0_u3_n864 ) );
  NOR2_X1 u0_u3_U282 (.ZN( u0_u3_n792 ) , .A2( u0_u3_n864 ) , .A1( u0_u3_n870 ) );
  NOR2_X1 u0_u3_U283 (.ZN( u0_u3_n464 ) , .A1( u0_u3_n832 ) , .A2( w3_26 ) );
  NOR2_X1 u0_u3_U284 (.ZN( u0_u3_n474 ) , .A1( u0_u3_n829 ) , .A2( w3_25 ) );
  AOI21_X1 u0_u3_U285 (.A( u0_u3_n439 ) , .ZN( u0_u3_n644 ) , .B1( u0_u3_n683 ) , .B2( u0_u3_n820 ) );
  AOI21_X1 u0_u3_U286 (.B2( u0_u3_n439 ) , .ZN( u0_u3_n500 ) , .A( u0_u3_n782 ) , .B1( u0_u3_n807 ) );
  OAI22_X1 u0_u3_U287 (.B1( u0_u3_n439 ) , .ZN( u0_u3_n698 ) , .A2( u0_u3_n733 ) , .A1( u0_u3_n783 ) , .B2( u0_u3_n820 ) );
  AOI21_X1 u0_u3_U288 (.B2( u0_u3_n439 ) , .ZN( u0_u3_n567 ) , .B1( u0_u3_n727 ) , .A( u0_u3_n782 ) );
  AOI21_X1 u0_u3_U289 (.B2( u0_u3_n439 ) , .ZN( u0_u3_n446 ) , .B1( u0_u3_n792 ) , .A( u0_u3_n817 ) );
  NOR4_X1 u0_u3_U29 (.A3( u0_u3_n603 ) , .A2( u0_u3_n604 ) , .A1( u0_u3_n605 ) , .ZN( u0_u3_n606 ) , .A4( u0_u3_n658 ) );
  NOR2_X1 u0_u3_U290 (.A2( u0_u3_n439 ) , .ZN( u0_u3_n667 ) , .A1( u0_u3_n788 ) );
  NOR2_X1 u0_u3_U291 (.A2( u0_u3_n439 ) , .ZN( u0_u3_n558 ) , .A1( u0_u3_n753 ) );
  NOR2_X1 u0_u3_U292 (.A2( u0_u3_n439 ) , .ZN( u0_u3_n562 ) , .A1( u0_u3_n806 ) );
  NOR2_X1 u0_u3_U293 (.A1( u0_u3_n439 ) , .ZN( u0_u3_n645 ) , .A2( u0_u3_n791 ) );
  NOR2_X1 u0_u3_U294 (.A2( u0_u3_n439 ) , .ZN( u0_u3_n545 ) , .A1( u0_u3_n765 ) );
  INV_X1 u0_u3_U295 (.A( u0_u3_n794 ) , .ZN( u0_u3_n875 ) );
  NOR2_X1 u0_u3_U296 (.ZN( u0_u3_n463 ) , .A1( u0_u3_n851 ) , .A2( w3_31 ) );
  AOI21_X1 u0_u3_U297 (.B2( u0_u3_n439 ) , .A( u0_u3_n793 ) , .B1( u0_u3_n795 ) , .ZN( u0_u3_n796 ) );
  AOI222_X1 u0_u3_U298 (.C2( u0_u3_n812 ) , .B2( u0_u3_n813 ) , .A2( u0_u3_n814 ) , .ZN( u0_u3_n826 ) , .C1( u0_u3_n835 ) , .A1( u0_u3_n841 ) , .B1( u0_u3_n855 ) );
  AOI22_X1 u0_u3_U299 (.ZN( u0_u3_n730 ) , .B1( u0_u3_n835 ) , .A2( u0_u3_n840 ) , .A1( u0_u3_n865 ) , .B2( u0_u3_n868 ) );
  BUF_X1 u0_u3_U3 (.Z( u0_u3_n438 ) , .A( u0_u3_n818 ) );
  NOR4_X1 u0_u3_U30 (.A4( u0_u3_n487 ) , .ZN( u0_u3_n490 ) , .A1( u0_u3_n569 ) , .A2( u0_u3_n584 ) , .A3( u0_u3_n605 ) );
  AOI222_X1 u0_u3_U300 (.ZN( u0_u3_n516 ) , .C1( u0_u3_n835 ) , .B2( u0_u3_n839 ) , .A2( u0_u3_n845 ) , .C2( u0_u3_n864 ) , .B1( u0_u3_n865 ) , .A1( u0_u3_n868 ) );
  AOI222_X1 u0_u3_U301 (.ZN( u0_u3_n472 ) , .B1( u0_u3_n835 ) , .A1( u0_u3_n841 ) , .C1( u0_u3_n844 ) , .C2( u0_u3_n853 ) , .A2( u0_u3_n857 ) , .B2( u0_u3_n867 ) );
  NOR2_X1 u0_u3_U302 (.A2( u0_u3_n438 ) , .ZN( u0_u3_n658 ) , .A1( u0_u3_n793 ) );
  NOR2_X1 u0_u3_U303 (.ZN( u0_u3_n715 ) , .A2( u0_u3_n727 ) , .A1( u0_u3_n793 ) );
  NOR2_X1 u0_u3_U304 (.ZN( u0_u3_n689 ) , .A1( u0_u3_n834 ) , .A2( u0_u3_n835 ) );
  NOR2_X1 u0_u3_U305 (.ZN( u0_u3_n524 ) , .A1( u0_u3_n793 ) , .A2( u0_u3_n815 ) );
  NOR2_X1 u0_u3_U306 (.ZN( u0_u3_n664 ) , .A1( u0_u3_n732 ) , .A2( u0_u3_n793 ) );
  NOR2_X1 u0_u3_U307 (.ZN( u0_u3_n736 ) , .A2( u0_u3_n835 ) , .A1( u0_u3_n847 ) );
  NOR2_X1 u0_u3_U308 (.ZN( u0_u3_n671 ) , .A2( u0_u3_n711 ) , .A1( u0_u3_n793 ) );
  NOR2_X1 u0_u3_U309 (.ZN( u0_u3_n673 ) , .A1( u0_u3_n793 ) , .A2( u0_u3_n808 ) );
  NOR4_X1 u0_u3_U31 (.ZN( u0_u3_n489 ) , .A1( u0_u3_n510 ) , .A2( u0_u3_n522 ) , .A4( u0_u3_n549 ) , .A3( u0_u3_n614 ) );
  INV_X1 u0_u3_U310 (.A( u0_u3_n793 ) , .ZN( u0_u3_n835 ) );
  AOI21_X1 u0_u3_U311 (.B1( u0_u3_n438 ) , .ZN( u0_u3_n513 ) , .B2( u0_u3_n672 ) , .A( u0_u3_n733 ) );
  AOI21_X1 u0_u3_U312 (.B1( u0_u3_n439 ) , .ZN( u0_u3_n629 ) , .B2( u0_u3_n672 ) , .A( u0_u3_n793 ) );
  INV_X1 u0_u3_U313 (.A( u0_u3_n672 ) , .ZN( u0_u3_n867 ) );
  NOR2_X1 u0_u3_U314 (.ZN( u0_u3_n655 ) , .A1( u0_u3_n672 ) , .A2( u0_u3_n817 ) );
  NOR2_X1 u0_u3_U315 (.ZN( u0_u3_n631 ) , .A2( u0_u3_n672 ) , .A1( u0_u3_n788 ) );
  NOR2_X1 u0_u3_U316 (.ZN( u0_u3_n605 ) , .A1( u0_u3_n672 ) , .A2( u0_u3_n806 ) );
  NOR2_X1 u0_u3_U317 (.ZN( u0_u3_n530 ) , .A1( u0_u3_n672 ) , .A2( u0_u3_n782 ) );
  NOR2_X1 u0_u3_U318 (.ZN( u0_u3_n584 ) , .A1( u0_u3_n672 ) , .A2( u0_u3_n791 ) );
  NOR2_X1 u0_u3_U319 (.ZN( u0_u3_n444 ) , .A2( w3_28 ) , .A1( w3_29 ) );
  NOR4_X1 u0_u3_U32 (.A4( u0_u3_n529 ) , .A2( u0_u3_n530 ) , .A1( u0_u3_n531 ) , .ZN( u0_u3_n541 ) , .A3( u0_u3_n704 ) );
  NOR2_X1 u0_u3_U320 (.ZN( u0_u3_n468 ) , .A2( u0_u3_n849 ) , .A1( u0_u3_n850 ) );
  OAI222_X1 u0_u3_U321 (.B2( u0_u3_n750 ) , .B1( u0_u3_n751 ) , .A2( u0_u3_n752 ) , .ZN( u0_u3_n760 ) , .C2( u0_u3_n808 ) , .C1( u0_u3_n817 ) , .A1( u0_u3_n820 ) );
  INV_X1 u0_u3_U322 (.A( u0_u3_n789 ) , .ZN( u0_u3_n864 ) );
  NOR4_X1 u0_u3_U323 (.A4( u0_u3_n617 ) , .A3( u0_u3_n618 ) , .A1( u0_u3_n619 ) , .A2( u0_u3_n620 ) , .ZN( u0_u3_n621 ) );
  INV_X1 u0_u3_U324 (.ZN( u0_u3_n830 ) , .A( w3_25 ) );
  OAI22_X1 u0_u3_U325 (.B2( u0_u3_n753 ) , .B1( u0_u3_n754 ) , .A1( u0_u3_n755 ) , .ZN( u0_u3_n759 ) , .A2( u0_u3_n809 ) );
  OAI22_X1 u0_u3_U326 (.B2( u0_u3_n806 ) , .B1( u0_u3_n807 ) , .A2( u0_u3_n808 ) , .A1( u0_u3_n809 ) , .ZN( u0_u3_n811 ) );
  AOI21_X1 u0_u3_U327 (.ZN( u0_u3_n692 ) , .B2( u0_u3_n752 ) , .B1( u0_u3_n766 ) , .A( u0_u3_n809 ) );
  NAND2_X1 u0_u3_U328 (.A2( u0_u3_n765 ) , .A1( u0_u3_n809 ) , .ZN( u0_u3_n813 ) );
  NOR2_X1 u0_u3_U329 (.ZN( u0_u3_n573 ) , .A1( u0_u3_n731 ) , .A2( u0_u3_n809 ) );
  NOR4_X1 u0_u3_U33 (.A4( u0_u3_n535 ) , .A3( u0_u3_n536 ) , .A2( u0_u3_n537 ) , .ZN( u0_u3_n538 ) , .A1( u0_u3_n823 ) );
  NOR2_X1 u0_u3_U330 (.ZN( u0_u3_n614 ) , .A2( u0_u3_n783 ) , .A1( u0_u3_n809 ) );
  OAI22_X1 u0_u3_U331 (.ZN( u0_u3_n486 ) , .A1( u0_u3_n711 ) , .B2( u0_u3_n788 ) , .A2( u0_u3_n809 ) , .B1( u0_u3_n815 ) );
  AOI21_X1 u0_u3_U332 (.ZN( u0_u3_n480 ) , .A( u0_u3_n672 ) , .B1( u0_u3_n753 ) , .B2( u0_u3_n809 ) );
  INV_X1 u0_u3_U333 (.A( u0_u3_n809 ) , .ZN( u0_u3_n843 ) );
  OAI221_X1 u0_u3_U334 (.A( u0_u3_n786 ) , .C2( u0_u3_n787 ) , .B2( u0_u3_n788 ) , .B1( u0_u3_n789 ) , .ZN( u0_u3_n799 ) , .C1( u0_u3_n816 ) );
  NAND2_X1 u0_u3_U335 (.A1( u0_u3_n732 ) , .A2( u0_u3_n787 ) , .ZN( u0_u3_n814 ) );
  OAI22_X1 u0_u3_U336 (.ZN( u0_u3_n591 ) , .A2( u0_u3_n750 ) , .B2( u0_u3_n765 ) , .A1( u0_u3_n766 ) , .B1( u0_u3_n787 ) );
  AOI21_X1 u0_u3_U337 (.ZN( u0_u3_n595 ) , .B1( u0_u3_n731 ) , .B2( u0_u3_n787 ) , .A( u0_u3_n793 ) );
  NOR2_X1 u0_u3_U338 (.ZN( u0_u3_n807 ) , .A1( u0_u3_n856 ) , .A2( u0_u3_n863 ) );
  AOI21_X1 u0_u3_U339 (.ZN( u0_u3_n626 ) , .B1( u0_u3_n702 ) , .A( u0_u3_n782 ) , .B2( u0_u3_n787 ) );
  NOR4_X1 u0_u3_U34 (.A4( u0_u3_n532 ) , .A3( u0_u3_n533 ) , .ZN( u0_u3_n540 ) , .A2( u0_u3_n687 ) , .A1( u0_u3_n797 ) );
  NAND2_X2 u0_u3_U340 (.A1( u0_u3_n458 ) , .A2( u0_u3_n465 ) , .ZN( u0_u3_n753 ) );
  AOI222_X1 u0_u3_U341 (.ZN( u0_u3_n778 ) , .A1( u0_u3_n833 ) , .C1( u0_u3_n837 ) , .B2( u0_u3_n843 ) , .A2( u0_u3_n852 ) , .B1( u0_u3_n863 ) , .C2( u0_u3_n875 ) );
  AOI222_X1 u0_u3_U342 (.ZN( u0_u3_n609 ) , .A1( u0_u3_n833 ) , .C2( u0_u3_n839 ) , .B1( u0_u3_n844 ) , .A2( u0_u3_n858 ) , .B2( u0_u3_n863 ) , .C1( u0_u3_n870 ) );
  AOI21_X1 u0_u3_U343 (.ZN( u0_u3_n651 ) , .A( u0_u3_n765 ) , .B2( u0_u3_n787 ) , .B1( u0_u3_n795 ) );
  OAI22_X1 u0_u3_U344 (.ZN( u0_u3_n684 ) , .A1( u0_u3_n702 ) , .A2( u0_u3_n733 ) , .B2( u0_u3_n787 ) , .B1( u0_u3_n820 ) );
  NOR2_X1 u0_u3_U345 (.ZN( u0_u3_n654 ) , .A1( u0_u3_n787 ) , .A2( u0_u3_n791 ) );
  NOR2_X1 u0_u3_U346 (.ZN( u0_u3_n751 ) , .A1( u0_u3_n863 ) , .A2( u0_u3_n864 ) );
  NOR2_X1 u0_u3_U347 (.ZN( u0_u3_n455 ) , .A1( u0_u3_n860 ) , .A2( w3_30 ) );
  NOR2_X1 u0_u3_U348 (.ZN( u0_u3_n467 ) , .A2( w3_30 ) , .A1( w3_31 ) );
  AND2_X1 u0_u3_U349 (.ZN( u0_u3_n441 ) , .A2( u0_u3_n834 ) , .A1( u0_u3_n856 ) );
  NOR3_X1 u0_u3_U35 (.A3( u0_u3_n803 ) , .A2( u0_u3_n804 ) , .A1( u0_u3_n805 ) , .ZN( u0_u3_n828 ) );
  AND2_X1 u0_u3_U350 (.ZN( u0_u3_n442 ) , .A2( u0_u3_n845 ) , .A1( u0_u3_n863 ) );
  NOR3_X1 u0_u3_U351 (.A3( u0_u3_n441 ) , .A2( u0_u3_n442 ) , .A1( u0_u3_n579 ) , .ZN( u0_u3_n590 ) );
  INV_X1 u0_u3_U352 (.A( u0_u3_n815 ) , .ZN( u0_u3_n856 ) );
  INV_X1 u0_u3_U353 (.A( u0_u3_n787 ) , .ZN( u0_u3_n863 ) );
  INV_X1 u0_u3_U354 (.A( u0_u3_n806 ) , .ZN( u0_u3_n845 ) );
  INV_X1 u0_u3_U355 (.A( u0_u3_n41 ) , .ZN( u0_u3_n840 ) );
  NOR2_X1 u0_u3_U356 (.A1( u0_u3_n41 ) , .ZN( u0_u3_n773 ) , .A2( u0_u3_n818 ) );
  AOI21_X1 u0_u3_U357 (.B2( u0_u3_n41 ) , .ZN( u0_u3_n574 ) , .B1( u0_u3_n809 ) , .A( u0_u3_n815 ) );
  NOR2_X1 u0_u3_U358 (.A2( u0_u3_n41 ) , .ZN( u0_u3_n665 ) , .A1( u0_u3_n732 ) );
  NOR2_X1 u0_u3_U359 (.A2( u0_u3_n41 ) , .ZN( u0_u3_n635 ) , .A1( u0_u3_n727 ) );
  NAND4_X1 u0_u3_U36 (.A4( u0_u3_n660 ) , .A3( u0_u3_n661 ) , .A2( u0_u3_n662 ) , .A1( u0_u3_n663 ) , .ZN( u0_u3_n803 ) );
  NOR2_X1 u0_u3_U360 (.A2( u0_u3_n41 ) , .A1( u0_u3_n783 ) , .ZN( u0_u3_n823 ) );
  AOI21_X1 u0_u3_U361 (.B2( u0_u3_n41 ) , .ZN( u0_u3_n481 ) , .A( u0_u3_n752 ) , .B1( u0_u3_n782 ) );
  NOR2_X1 u0_u3_U362 (.A2( u0_u3_n41 ) , .ZN( u0_u3_n569 ) , .A1( u0_u3_n766 ) );
  NOR2_X1 u0_u3_U363 (.A2( u0_u3_n41 ) , .ZN( u0_u3_n719 ) , .A1( u0_u3_n795 ) );
  NOR2_X1 u0_u3_U364 (.A2( u0_u3_n41 ) , .ZN( u0_u3_n597 ) , .A1( u0_u3_n731 ) );
  AOI21_X1 u0_u3_U365 (.A( u0_u3_n41 ) , .ZN( u0_u3_n555 ) , .B1( u0_u3_n672 ) , .B2( u0_u3_n808 ) );
  NOR2_X1 u0_u3_U366 (.A2( u0_u3_n41 ) , .ZN( u0_u3_n544 ) , .A1( u0_u3_n702 ) );
  NOR2_X1 u0_u3_U367 (.ZN( u0_u3_n583 ) , .A2( u0_u3_n700 ) , .A1( u0_u3_n794 ) );
  NOR4_X1 u0_u3_U368 (.A4( u0_u3_n779 ) , .A3( u0_u3_n780 ) , .A1( u0_u3_n781 ) , .ZN( u0_u3_n802 ) , .A2( u0_u3_n804 ) );
  NAND4_X1 u0_u3_U369 (.A4( u0_u3_n694 ) , .A3( u0_u3_n695 ) , .A1( u0_u3_n696 ) , .ZN( u0_u3_n779 ) , .A2( u0_u3_n874 ) );
  NOR3_X1 u0_u3_U37 (.A3( u0_u3_n654 ) , .A2( u0_u3_n655 ) , .A1( u0_u3_n656 ) , .ZN( u0_u3_n661 ) );
  AOI21_X1 u0_u3_U370 (.ZN( u0_u3_n596 ) , .B1( u0_u3_n753 ) , .A( u0_u3_n795 ) , .B2( u0_u3_n816 ) );
  AOI21_X1 u0_u3_U371 (.A( u0_u3_n815 ) , .B2( u0_u3_n816 ) , .B1( u0_u3_n817 ) , .ZN( u0_u3_n822 ) );
  OAI222_X1 u0_u3_U372 (.ZN( u0_u3_n508 ) , .C2( u0_u3_n628 ) , .B2( u0_u3_n650 ) , .B1( u0_u3_n750 ) , .A2( u0_u3_n751 ) , .C1( u0_u3_n808 ) , .A1( u0_u3_n809 ) );
  AOI21_X1 u0_u3_U373 (.B1( u0_u3_n628 ) , .ZN( u0_u3_n630 ) , .A( u0_u3_n766 ) , .B2( u0_u3_n817 ) );
  AOI21_X1 u0_u3_U374 (.ZN( u0_u3_n652 ) , .B1( u0_u3_n732 ) , .B2( u0_u3_n766 ) , .A( u0_u3_n816 ) );
  OAI21_X1 u0_u3_U375 (.A( u0_u3_n616 ) , .ZN( u0_u3_n619 ) , .B1( u0_u3_n628 ) , .B2( u0_u3_n787 ) );
  NOR2_X1 u0_u3_U376 (.A1( u0_u3_n672 ) , .ZN( u0_u3_n769 ) , .A2( u0_u3_n816 ) );
  NOR2_X1 u0_u3_U377 (.A2( u0_u3_n816 ) , .A1( u0_u3_n818 ) , .ZN( u0_u3_n824 ) );
  NOR2_X1 u0_u3_U378 (.ZN( u0_u3_n581 ) , .A1( u0_u3_n711 ) , .A2( u0_u3_n816 ) );
  NOR2_X1 u0_u3_U379 (.A1( u0_u3_n439 ) , .ZN( u0_u3_n687 ) , .A2( u0_u3_n816 ) );
  NOR3_X1 u0_u3_U38 (.A3( u0_u3_n651 ) , .A2( u0_u3_n652 ) , .A1( u0_u3_n653 ) , .ZN( u0_u3_n662 ) );
  NOR2_X1 u0_u3_U380 (.ZN( u0_u3_n657 ) , .A1( u0_u3_n731 ) , .A2( u0_u3_n816 ) );
  NOR2_X1 u0_u3_U381 (.A1( u0_u3_n702 ) , .ZN( u0_u3_n771 ) , .A2( u0_u3_n816 ) );
  NOR2_X1 u0_u3_U382 (.ZN( u0_u3_n668 ) , .A1( u0_u3_n783 ) , .A2( u0_u3_n816 ) );
  NOR2_X1 u0_u3_U383 (.ZN( u0_u3_n634 ) , .A1( u0_u3_n727 ) , .A2( u0_u3_n816 ) );
  NOR2_X1 u0_u3_U384 (.ZN( u0_u3_n475 ) , .A2( w3_26 ) , .A1( w3_27 ) );
  NOR2_X1 u0_u3_U385 (.ZN( u0_u3_n458 ) , .A1( u0_u3_n831 ) , .A2( w3_27 ) );
  INV_X1 u0_u3_U386 (.ZN( u0_u3_n832 ) , .A( w3_27 ) );
  NOR3_X1 u0_u3_U387 (.A3( u0_u3_n624 ) , .A2( u0_u3_n625 ) , .ZN( u0_u3_n639 ) , .A1( u0_u3_n728 ) );
  NOR4_X1 u0_u3_U388 (.A1( u0_u3_n587 ) , .ZN( u0_u3_n588 ) , .A3( u0_u3_n655 ) , .A2( u0_u3_n665 ) , .A4( u0_u3_n770 ) );
  OAI22_X1 u0_u3_U389 (.ZN( u0_u3_n640 ) , .A1( u0_u3_n702 ) , .B2( u0_u3_n731 ) , .A2( u0_u3_n765 ) , .B1( u0_u3_n819 ) );
  NOR3_X1 u0_u3_U39 (.A3( u0_u3_n657 ) , .A2( u0_u3_n658 ) , .A1( u0_u3_n659 ) , .ZN( u0_u3_n660 ) );
  AOI21_X1 u0_u3_U390 (.ZN( u0_u3_n502 ) , .B1( u0_u3_n683 ) , .A( u0_u3_n815 ) , .B2( u0_u3_n819 ) );
  OAI22_X1 u0_u3_U391 (.A1( u0_u3_n727 ) , .ZN( u0_u3_n729 ) , .B2( u0_u3_n753 ) , .B1( u0_u3_n815 ) , .A2( u0_u3_n819 ) );
  AOI21_X1 u0_u3_U392 (.A( u0_u3_n438 ) , .B2( u0_u3_n819 ) , .B1( u0_u3_n820 ) , .ZN( u0_u3_n821 ) );
  OAI22_X1 u0_u3_U393 (.A1( u0_u3_n438 ) , .ZN( u0_u3_n627 ) , .B1( u0_u3_n672 ) , .B2( u0_u3_n750 ) , .A2( u0_u3_n819 ) );
  NOR2_X1 u0_u3_U394 (.ZN( u0_u3_n522 ) , .A2( u0_u3_n702 ) , .A1( u0_u3_n819 ) );
  NOR2_X1 u0_u3_U395 (.A1( u0_u3_n672 ) , .ZN( u0_u3_n691 ) , .A2( u0_u3_n819 ) );
  NOR2_X1 u0_u3_U396 (.A2( u0_u3_n439 ) , .ZN( u0_u3_n602 ) , .A1( u0_u3_n819 ) );
  NOR2_X1 u0_u3_U397 (.ZN( u0_u3_n534 ) , .A2( u0_u3_n783 ) , .A1( u0_u3_n819 ) );
  NOR2_X1 u0_u3_U398 (.ZN( u0_u3_n561 ) , .A1( u0_u3_n711 ) , .A2( u0_u3_n819 ) );
  NOR2_X1 u0_u3_U399 (.ZN( u0_u3_n688 ) , .A1( u0_u3_n732 ) , .A2( u0_u3_n819 ) );
  NAND2_X1 u0_u3_U4 (.A1( u0_u3_n452 ) , .A2( u0_u3_n463 ) , .ZN( u0_u3_n795 ) );
  NOR4_X1 u0_u3_U40 (.A4( u0_u3_n664 ) , .A3( u0_u3_n665 ) , .A2( u0_u3_n666 ) , .A1( u0_u3_n667 ) , .ZN( u0_u3_n680 ) );
  INV_X1 u0_u3_U400 (.A( u0_u3_n819 ) , .ZN( u0_u3_n834 ) );
  NAND2_X1 u0_u3_U401 (.ZN( u0_u3_n674 ) , .A1( u0_u3_n809 ) , .A2( u0_u3_n819 ) );
  NOR2_X1 u0_u3_U402 (.ZN( u0_u3_n465 ) , .A2( w3_24 ) , .A1( w3_25 ) );
  NOR2_X1 u0_u3_U403 (.ZN( u0_u3_n457 ) , .A1( u0_u3_n830 ) , .A2( w3_24 ) );
  INV_X1 u0_u3_U404 (.ZN( u0_u3_n829 ) , .A( w3_24 ) );
  INV_X1 u0_u3_U405 (.ZN( u0_u3_n850 ) , .A( w3_29 ) );
  NOR2_X1 u0_u3_U406 (.ZN( u0_u3_n451 ) , .A1( u0_u3_n849 ) , .A2( w3_29 ) );
  NAND4_X1 u0_u3_U407 (.ZN( u0_subword_3 ) , .A4( u0_u3_n707 ) , .A3( u0_u3_n708 ) , .A2( u0_u3_n709 ) , .A1( u0_u3_n710 ) );
  INV_X1 u0_u3_U408 (.A( u0_u3_n709 ) , .ZN( u0_u3_n878 ) );
  OAI22_X1 u0_u3_U409 (.B2( u0_u3_n747 ) , .ZN( u0_u3_n749 ) , .A2( u0_u3_n765 ) , .B1( u0_u3_n783 ) , .A1( u0_u3_n795 ) );
  NOR4_X1 u0_u3_U41 (.A4( u0_u3_n668 ) , .A3( u0_u3_n669 ) , .A2( u0_u3_n670 ) , .A1( u0_u3_n671 ) , .ZN( u0_u3_n679 ) );
  OAI22_X1 u0_u3_U410 (.B1( u0_u3_n439 ) , .ZN( u0_u3_n499 ) , .A2( u0_u3_n747 ) , .A1( u0_u3_n783 ) , .B2( u0_u3_n809 ) );
  NOR2_X1 u0_u3_U411 (.ZN( u0_u3_n519 ) , .A1( u0_u3_n711 ) , .A2( u0_u3_n747 ) );
  OAI22_X1 u0_u3_U412 (.ZN( u0_u3_n713 ) , .A2( u0_u3_n731 ) , .B2( u0_u3_n732 ) , .A1( u0_u3_n747 ) , .B1( u0_u3_n816 ) );
  NOR2_X1 u0_u3_U413 (.A2( u0_u3_n747 ) , .ZN( u0_u3_n772 ) , .A1( u0_u3_n815 ) );
  OAI22_X1 u0_u3_U414 (.B1( u0_u3_n443 ) , .ZN( u0_u3_n447 ) , .A2( u0_u3_n731 ) , .A1( u0_u3_n747 ) , .B2( u0_u3_n752 ) );
  NOR2_X1 u0_u3_U415 (.ZN( u0_u3_n550 ) , .A1( u0_u3_n702 ) , .A2( u0_u3_n747 ) );
  NOR2_X1 u0_u3_U416 (.ZN( u0_u3_n556 ) , .A2( u0_u3_n747 ) , .A1( u0_u3_n787 ) );
  NOR2_X1 u0_u3_U417 (.A2( u0_u3_n747 ) , .ZN( u0_u3_n758 ) , .A1( u0_u3_n808 ) );
  NOR2_X1 u0_u3_U418 (.A1( u0_u3_n672 ) , .ZN( u0_u3_n676 ) , .A2( u0_u3_n747 ) );
  NOR2_X1 u0_u3_U419 (.ZN( u0_u3_n533 ) , .A2( u0_u3_n747 ) , .A1( u0_u3_n795 ) );
  NOR4_X1 u0_u3_U42 (.A3( u0_u3_n676 ) , .A1( u0_u3_n677 ) , .ZN( u0_u3_n678 ) , .A4( u0_u3_n718 ) , .A2( u0_u3_n861 ) );
  NOR2_X1 u0_u3_U420 (.ZN( u0_u3_n721 ) , .A2( u0_u3_n727 ) , .A1( u0_u3_n747 ) );
  NOR2_X1 u0_u3_U421 (.ZN( u0_u3_n585 ) , .A1( u0_u3_n747 ) , .A2( u0_u3_n818 ) );
  INV_X1 u0_u3_U422 (.A( u0_u3_n747 ) , .ZN( u0_u3_n839 ) );
  AOI21_X1 u0_u3_U423 (.ZN( u0_u3_n579 ) , .B2( u0_u3_n727 ) , .B1( u0_u3_n751 ) , .A( u0_u3_n788 ) );
  NAND4_X1 u0_u3_U424 (.A4( u0_u3_n636 ) , .A3( u0_u3_n637 ) , .A2( u0_u3_n638 ) , .A1( u0_u3_n639 ) , .ZN( u0_u3_n746 ) );
  INV_X1 u0_u3_U425 (.ZN( u0_u3_n851 ) , .A( w3_30 ) );
  INV_X1 u0_u3_U426 (.ZN( u0_u3_n860 ) , .A( w3_31 ) );
  NAND4_X1 u0_u3_U427 (.ZN( u0_subword_2 ) , .A4( u0_u3_n646 ) , .A3( u0_u3_n647 ) , .A2( u0_u3_n648 ) , .A1( u0_u3_n649 ) );
  AOI211_X1 u0_u3_U428 (.A( u0_u3_n640 ) , .ZN( u0_u3_n648 ) , .B( u0_u3_n746 ) , .C2( u0_u3_n841 ) , .C1( u0_u3_n856 ) );
  NOR2_X1 u0_u3_U429 (.A2( u0_u3_n41 ) , .ZN( u0_u3_n603 ) , .A1( u0_u3_n787 ) );
  NOR4_X1 u0_u3_U43 (.A1( u0_u3_n469 ) , .ZN( u0_u3_n470 ) , .A4( u0_u3_n545 ) , .A2( u0_u3_n557 ) , .A3( u0_u3_n617 ) );
  OAI222_X1 u0_u3_U430 (.A2( u0_u3_n672 ) , .ZN( u0_u3_n677 ) , .B1( u0_u3_n750 ) , .B2( u0_u3_n787 ) , .C2( u0_u3_n791 ) , .C1( u0_u3_n818 ) , .A1( u0_u3_n820 ) );
  NOR2_X1 u0_u3_U431 (.ZN( u0_u3_n613 ) , .A1( u0_u3_n787 ) , .A2( u0_u3_n819 ) );
  AOI21_X1 u0_u3_U432 (.A( u0_u3_n41 ) , .ZN( u0_u3_n503 ) , .B1( u0_u3_n711 ) , .B2( u0_u3_n789 ) );
  OAI22_X1 u0_u3_U433 (.ZN( u0_u3_n593 ) , .B1( u0_u3_n733 ) , .B2( u0_u3_n752 ) , .A2( u0_u3_n789 ) , .A1( u0_u3_n806 ) );
  NOR2_X1 u0_u3_U434 (.ZN( u0_u3_n656 ) , .A1( u0_u3_n765 ) , .A2( u0_u3_n789 ) );
  NAND2_X1 u0_u3_U435 (.A2( u0_u3_n752 ) , .A1( u0_u3_n789 ) , .ZN( u0_u3_n812 ) );
  NOR2_X1 u0_u3_U436 (.ZN( u0_u3_n557 ) , .A1( u0_u3_n789 ) , .A2( u0_u3_n816 ) );
  NAND3_X1 u0_u3_U437 (.ZN( u0_subword_6 ) , .A3( u0_u3_n800 ) , .A2( u0_u3_n801 ) , .A1( u0_u3_n802 ) );
  NAND3_X1 u0_u3_U438 (.ZN( u0_subword_5 ) , .A3( u0_u3_n761 ) , .A2( u0_u3_n762 ) , .A1( u0_u3_n763 ) );
  NAND3_X1 u0_u3_U439 (.ZN( u0_subword_4 ) , .A3( u0_u3_n741 ) , .A2( u0_u3_n742 ) , .A1( u0_u3_n743 ) );
  AOI221_X1 u0_u3_U44 (.ZN( u0_u3_n471 ) , .C2( u0_u3_n717 ) , .B2( u0_u3_n834 ) , .C1( u0_u3_n847 ) , .B1( u0_u3_n862 ) , .A( u0_u3_n866 ) );
  NAND3_X1 u0_u3_U440 (.A3( u0_u3_n678 ) , .A2( u0_u3_n679 ) , .A1( u0_u3_n680 ) , .ZN( u0_u3_n810 ) );
  NAND3_X1 u0_u3_U441 (.ZN( u0_u3_n641 ) , .A3( u0_u3_n711 ) , .A2( u0_u3_n727 ) , .A1( u0_u3_n795 ) );
  NAND3_X1 u0_u3_U442 (.A3( u0_u3_n621 ) , .A2( u0_u3_n622 ) , .A1( u0_u3_n623 ) , .ZN( u0_u3_n728 ) );
  NAND3_X1 u0_u3_U443 (.A3( u0_u3_n588 ) , .A2( u0_u3_n589 ) , .A1( u0_u3_n590 ) , .ZN( u0_u3_n624 ) );
  NAND3_X1 u0_u3_U444 (.ZN( u0_u3_n568 ) , .A3( u0_u3_n683 ) , .A2( u0_u3_n753 ) , .A1( u0_u3_n788 ) );
  NAND3_X1 u0_u3_U445 (.A3( u0_u3_n526 ) , .A2( u0_u3_n527 ) , .A1( u0_u3_n528 ) , .ZN( u0_u3_n745 ) );
  NAND3_X1 u0_u3_U446 (.A3( u0_u3_n515 ) , .A1( u0_u3_n516 ) , .ZN( u0_u3_n611 ) , .A2( u0_u3_n873 ) );
  NAND3_X1 u0_u3_U447 (.A3( u0_u3_n470 ) , .A2( u0_u3_n471 ) , .A1( u0_u3_n472 ) , .ZN( u0_u3_n780 ) );
  NOR2_X1 u0_u3_U448 (.ZN( u0_u3_n615 ) , .A1( u0_u3_n782 ) , .A2( u0_u3_n789 ) );
  NOR2_X1 u0_u3_U449 (.ZN( u0_u3_n720 ) , .A2( u0_u3_n747 ) , .A1( u0_u3_n789 ) );
  NOR4_X1 u0_u3_U45 (.A4( u0_u3_n517 ) , .A3( u0_u3_n518 ) , .A2( u0_u3_n519 ) , .A1( u0_u3_n520 ) , .ZN( u0_u3_n527 ) );
  NOR2_X1 u0_u3_U450 (.ZN( u0_u3_n704 ) , .A2( u0_u3_n789 ) , .A1( u0_u3_n820 ) );
  NOR2_X1 u0_u3_U451 (.A1( u0_u3_n733 ) , .ZN( u0_u3_n768 ) , .A2( u0_u3_n789 ) );
  INV_X1 u0_u3_U452 (.ZN( u0_u3_n849 ) , .A( w3_28 ) );
  NOR4_X1 u0_u3_U46 (.A3( u0_u3_n524 ) , .A1( u0_u3_n525 ) , .ZN( u0_u3_n526 ) , .A2( u0_u3_n676 ) , .A4( u0_u3_n772 ) );
  NAND4_X1 u0_u3_U47 (.A4( u0_u3_n576 ) , .A3( u0_u3_n577 ) , .A1( u0_u3_n578 ) , .ZN( u0_u3_n726 ) , .A2( u0_u3_n876 ) );
  NOR4_X1 u0_u3_U48 (.A4( u0_u3_n572 ) , .A3( u0_u3_n573 ) , .A2( u0_u3_n574 ) , .A1( u0_u3_n575 ) , .ZN( u0_u3_n576 ) );
  INV_X1 u0_u3_U49 (.A( u0_u3_n610 ) , .ZN( u0_u3_n876 ) );
  NAND2_X1 u0_u3_U5 (.A1( u0_u3_n456 ) , .A2( u0_u3_n475 ) , .ZN( u0_u3_n788 ) );
  NAND4_X1 u0_u3_U50 (.A4( u0_u3_n459 ) , .A3( u0_u3_n460 ) , .A2( u0_u3_n461 ) , .A1( u0_u3_n462 ) , .ZN( u0_u3_n682 ) );
  NOR3_X1 u0_u3_U51 (.ZN( u0_u3_n460 ) , .A3( u0_u3_n533 ) , .A1( u0_u3_n558 ) , .A2( u0_u3_n573 ) );
  NOR4_X1 u0_u3_U52 (.ZN( u0_u3_n459 ) , .A2( u0_u3_n520 ) , .A1( u0_u3_n546 ) , .A3( u0_u3_n582 ) , .A4( u0_u3_n618 ) );
  NOR4_X1 u0_u3_U53 (.ZN( u0_u3_n461 ) , .A2( u0_u3_n512 ) , .A1( u0_u3_n602 ) , .A4( u0_u3_n631 ) , .A3( u0_u3_n714 ) );
  NAND4_X1 u0_u3_U54 (.A4( u0_u3_n722 ) , .A3( u0_u3_n723 ) , .A2( u0_u3_n724 ) , .ZN( u0_u3_n744 ) , .A1( u0_u3_n859 ) );
  INV_X1 u0_u3_U55 (.A( u0_u3_n712 ) , .ZN( u0_u3_n859 ) );
  NOR4_X1 u0_u3_U56 (.A4( u0_u3_n718 ) , .A3( u0_u3_n719 ) , .A2( u0_u3_n720 ) , .A1( u0_u3_n721 ) , .ZN( u0_u3_n722 ) );
  NOR3_X1 u0_u3_U57 (.ZN( u0_u3_n483 ) , .A2( u0_u3_n511 ) , .A3( u0_u3_n604 ) , .A1( u0_u3_n613 ) );
  NOR4_X1 u0_u3_U58 (.ZN( u0_u3_n484 ) , .A3( u0_u3_n535 ) , .A4( u0_u3_n548 ) , .A2( u0_u3_n570 ) , .A1( u0_u3_n720 ) );
  AOI211_X1 u0_u3_U59 (.B( u0_u3_n480 ) , .A( u0_u3_n481 ) , .ZN( u0_u3_n485 ) , .C2( u0_u3_n836 ) , .C1( u0_u3_n863 ) );
  NOR3_X1 u0_u3_U6 (.ZN( u0_u3_n601 ) , .A1( u0_u3_n611 ) , .A3( u0_u3_n726 ) , .A2( u0_u3_n745 ) );
  INV_X1 u0_u3_U60 (.A( u0_u3_n682 ) , .ZN( u0_u3_n874 ) );
  NOR4_X1 u0_u3_U61 (.A4( u0_u3_n690 ) , .A3( u0_u3_n691 ) , .A2( u0_u3_n692 ) , .A1( u0_u3_n693 ) , .ZN( u0_u3_n694 ) );
  AOI221_X1 u0_u3_U62 (.A( u0_u3_n684 ) , .ZN( u0_u3_n695 ) , .B2( u0_u3_n842 ) , .C1( u0_u3_n844 ) , .C2( u0_u3_n864 ) , .B1( u0_u3_n867 ) );
  NAND4_X1 u0_u3_U63 (.A4( u0_u3_n476 ) , .A3( u0_u3_n477 ) , .A2( u0_u3_n478 ) , .A1( u0_u3_n479 ) , .ZN( u0_u3_n681 ) );
  NOR4_X1 u0_u3_U64 (.A4( u0_u3_n473 ) , .ZN( u0_u3_n479 ) , .A3( u0_u3_n559 ) , .A1( u0_u3_n738 ) , .A2( u0_u3_n758 ) );
  NOR4_X1 u0_u3_U65 (.ZN( u0_u3_n477 ) , .A1( u0_u3_n509 ) , .A3( u0_u3_n547 ) , .A2( u0_u3_n586 ) , .A4( u0_u3_n719 ) );
  NOR4_X1 u0_u3_U66 (.ZN( u0_u3_n476 ) , .A2( u0_u3_n524 ) , .A4( u0_u3_n597 ) , .A1( u0_u3_n612 ) , .A3( u0_u3_n632 ) );
  NAND4_X1 u0_u3_U67 (.A4( u0_u3_n551 ) , .A3( u0_u3_n552 ) , .A2( u0_u3_n553 ) , .A1( u0_u3_n554 ) , .ZN( u0_u3_n748 ) );
  AOI211_X1 u0_u3_U68 (.B( u0_u3_n542 ) , .A( u0_u3_n543 ) , .ZN( u0_u3_n554 ) , .C2( u0_u3_n841 ) , .C1( u0_u3_n853 ) );
  NOR3_X1 u0_u3_U69 (.ZN( u0_u3_n552 ) , .A2( u0_u3_n654 ) , .A1( u0_u3_n670 ) , .A3( u0_u3_n774 ) );
  NOR3_X1 u0_u3_U7 (.ZN( u0_u3_n507 ) , .A2( u0_u3_n682 ) , .A3( u0_u3_n780 ) , .A1( u0_u3_n878 ) );
  NOR4_X1 u0_u3_U70 (.A4( u0_u3_n544 ) , .A3( u0_u3_n545 ) , .A2( u0_u3_n546 ) , .ZN( u0_u3_n553 ) , .A1( u0_u3_n691 ) );
  NOR4_X1 u0_u3_U71 (.A4( u0_u3_n612 ) , .A3( u0_u3_n613 ) , .A2( u0_u3_n614 ) , .A1( u0_u3_n615 ) , .ZN( u0_u3_n622 ) );
  NOR4_X1 u0_u3_U72 (.ZN( u0_u3_n623 ) , .A1( u0_u3_n659 ) , .A3( u0_u3_n669 ) , .A4( u0_u3_n685 ) , .A2( u0_u3_n769 ) );
  INV_X1 u0_u3_U73 (.A( u0_u3_n765 ) , .ZN( u0_u3_n833 ) );
  NOR2_X1 u0_u3_U74 (.ZN( u0_u3_n650 ) , .A1( u0_u3_n856 ) , .A2( u0_u3_n870 ) );
  NOR4_X1 u0_u3_U75 (.A4( u0_u3_n580 ) , .A3( u0_u3_n581 ) , .A2( u0_u3_n582 ) , .ZN( u0_u3_n589 ) , .A1( u0_u3_n686 ) );
  INV_X1 u0_u3_U76 (.A( u0_u3_n818 ) , .ZN( u0_u3_n857 ) );
  OR4_X1 u0_u3_U77 (.A4( u0_u3_n685 ) , .A3( u0_u3_n686 ) , .A2( u0_u3_n687 ) , .A1( u0_u3_n688 ) , .ZN( u0_u3_n693 ) );
  OR4_X1 u0_u3_U78 (.ZN( u0_u3_n469 ) , .A4( u0_u3_n521 ) , .A3( u0_u3_n532 ) , .A2( u0_u3_n581 ) , .A1( u0_u3_n715 ) );
  OR4_X1 u0_u3_U79 (.A4( u0_u3_n569 ) , .A3( u0_u3_n570 ) , .A2( u0_u3_n571 ) , .ZN( u0_u3_n575 ) , .A1( u0_u3_n668 ) );
  NOR3_X1 u0_u3_U8 (.A2( u0_u3_n610 ) , .A1( u0_u3_n611 ) , .ZN( u0_u3_n649 ) , .A3( u0_u3_n725 ) );
  OR4_X1 u0_u3_U80 (.A4( u0_u3_n521 ) , .A2( u0_u3_n522 ) , .A1( u0_u3_n523 ) , .ZN( u0_u3_n525 ) , .A3( u0_u3_n824 ) );
  OR4_X1 u0_u3_U81 (.A4( u0_u3_n583 ) , .A3( u0_u3_n584 ) , .A2( u0_u3_n585 ) , .A1( u0_u3_n586 ) , .ZN( u0_u3_n587 ) );
  OR4_X1 u0_u3_U82 (.ZN( u0_u3_n495 ) , .A4( u0_u3_n537 ) , .A2( u0_u3_n550 ) , .A1( u0_u3_n562 ) , .A3( u0_u3_n635 ) );
  NOR4_X1 u0_u3_U83 (.A4( u0_u3_n512 ) , .A2( u0_u3_n513 ) , .A1( u0_u3_n514 ) , .ZN( u0_u3_n515 ) , .A3( u0_u3_n673 ) );
  INV_X1 u0_u3_U84 (.A( u0_u3_n508 ) , .ZN( u0_u3_n873 ) );
  OR3_X1 u0_u3_U85 (.A3( u0_u3_n509 ) , .A2( u0_u3_n510 ) , .A1( u0_u3_n511 ) , .ZN( u0_u3_n514 ) );
  INV_X1 u0_u3_U86 (.A( u0_u3_n757 ) , .ZN( u0_u3_n871 ) );
  AOI221_X1 u0_u3_U87 (.A( u0_u3_n716 ) , .B2( u0_u3_n717 ) , .ZN( u0_u3_n723 ) , .C1( u0_u3_n835 ) , .B1( u0_u3_n841 ) , .C2( u0_u3_n865 ) );
  OR2_X1 u0_u3_U88 (.A2( u0_u3_n714 ) , .A1( u0_u3_n715 ) , .ZN( u0_u3_n716 ) );
  INV_X1 u0_u3_U89 (.A( u0_u3_n466 ) , .ZN( u0_u3_n866 ) );
  NOR3_X1 u0_u3_U9 (.A3( u0_u3_n725 ) , .A1( u0_u3_n726 ) , .ZN( u0_u3_n743 ) , .A2( u0_u3_n744 ) );
  NAND2_X1 u0_u3_U90 (.A1( u0_u3_n454 ) , .A2( u0_u3_n456 ) , .ZN( u0_u3_n765 ) );
  AOI22_X1 u0_u3_U91 (.ZN( u0_u3_n699 ) , .A1( u0_u3_n833 ) , .B2( u0_u3_n845 ) , .A2( u0_u3_n867 ) , .B1( u0_u3_n870 ) );
  NOR3_X1 u0_u3_U92 (.ZN( u0_u3_n755 ) , .A2( u0_u3_n855 ) , .A1( u0_u3_n865 ) , .A3( u0_u3_n867 ) );
  NOR2_X1 u0_u3_U93 (.ZN( u0_u3_n754 ) , .A2( u0_u3_n854 ) , .A1( u0_u3_n862 ) );
  AOI211_X1 u0_u3_U94 (.A( u0_u3_n499 ) , .ZN( u0_u3_n506 ) , .B( u0_u3_n805 ) , .C2( u0_u3_n841 ) , .C1( u0_u3_n853 ) );
  AOI211_X1 u0_u3_U95 (.B( u0_u3_n810 ) , .A( u0_u3_n811 ) , .ZN( u0_u3_n827 ) , .C1( u0_u3_n844 ) , .C2( u0_u3_n852 ) );
  NAND2_X1 u0_u3_U96 (.A1( u0_u3_n450 ) , .A2( u0_u3_n468 ) , .ZN( u0_u3_n752 ) );
  INV_X1 u0_u3_U97 (.A( u0_u3_n733 ) , .ZN( u0_u3_n841 ) );
  AOI221_X1 u0_u3_U98 (.B2( u0_u3_n440 ) , .A( u0_u3_n492 ) , .ZN( u0_u3_n497 ) , .C2( u0_u3_n843 ) , .C1( u0_u3_n853 ) , .B1( u0_u3_n862 ) );
  INV_X1 u0_u3_U99 (.A( u0_u3_n781 ) , .ZN( u0_u3_n869 ) );
  NOR2_X1 us00_U10 (.A2( us00_n132 ) , .A1( us00_n255 ) , .ZN( us00_n302 ) );
  NOR4_X1 us00_U100 (.A2( us00_n193 ) , .ZN( us00_n340 ) , .A3( us00_n347 ) , .A4( us00_n348 ) , .A1( us00_n83 ) );
  NAND4_X1 us00_U101 (.ZN( us00_n183 ) , .A1( us00_n395 ) , .A2( us00_n396 ) , .A3( us00_n397 ) , .A4( us00_n398 ) );
  NOR3_X1 us00_U102 (.A1( us00_n267 ) , .A3( us00_n276 ) , .A2( us00_n369 ) , .ZN( us00_n397 ) );
  AOI211_X1 us00_U103 (.C1( us00_n16 ) , .ZN( us00_n395 ) , .A( us00_n399 ) , .B( us00_n400 ) , .C2( us00_n44 ) );
  NOR4_X1 us00_U104 (.A1( us00_n160 ) , .A2( us00_n310 ) , .A4( us00_n332 ) , .A3( us00_n345 ) , .ZN( us00_n396 ) );
  NAND4_X1 us00_U105 (.ZN( us00_n132 ) , .A1( us00_n326 ) , .A2( us00_n327 ) , .A3( us00_n328 ) , .A4( us00_n329 ) );
  NOR3_X1 us00_U106 (.A3( us00_n106 ) , .A1( us00_n210 ) , .A2( us00_n226 ) , .ZN( us00_n328 ) );
  AOI211_X1 us00_U107 (.C1( us00_n26 ) , .ZN( us00_n326 ) , .A( us00_n337 ) , .B( us00_n338 ) , .C2( us00_n38 ) );
  NOR4_X1 us00_U108 (.ZN( us00_n329 ) , .A1( us00_n330 ) , .A2( us00_n331 ) , .A3( us00_n332 ) , .A4( us00_n333 ) );
  NOR2_X1 us00_U109 (.ZN( us00_n191 ) , .A2( us00_n45 ) , .A1( us00_n46 ) );
  NOR2_X1 us00_U11 (.ZN( us00_n184 ) , .A1( us00_n199 ) , .A2( us00_n70 ) );
  NOR4_X1 us00_U110 (.A2( us00_n111 ) , .A4( us00_n195 ) , .A3( us00_n211 ) , .A1( us00_n221 ) , .ZN( us00_n257 ) );
  NOR4_X1 us00_U111 (.ZN( us00_n258 ) , .A1( us00_n265 ) , .A2( us00_n266 ) , .A3( us00_n267 ) , .A4( us00_n268 ) );
  NOR4_X1 us00_U112 (.ZN( us00_n259 ) , .A1( us00_n260 ) , .A2( us00_n261 ) , .A3( us00_n262 ) , .A4( us00_n263 ) );
  NAND4_X1 us00_U113 (.A1( us00_n389 ) , .A2( us00_n390 ) , .A3( us00_n391 ) , .A4( us00_n392 ) , .ZN( us00_n99 ) );
  NOR4_X1 us00_U114 (.A3( us00_n275 ) , .A2( us00_n296 ) , .A1( us00_n311 ) , .ZN( us00_n390 ) , .A4( us00_n393 ) );
  NOR4_X1 us00_U115 (.A3( us00_n266 ) , .A4( us00_n331 ) , .A2( us00_n358 ) , .A1( us00_n370 ) , .ZN( us00_n391 ) );
  NOR4_X1 us00_U116 (.A4( us00_n159 ) , .A3( us00_n246 ) , .A1( us00_n319 ) , .A2( us00_n344 ) , .ZN( us00_n392 ) );
  NAND4_X1 us00_U117 (.ZN( us00_n101 ) , .A1( us00_n184 ) , .A3( us00_n185 ) , .A4( us00_n186 ) , .A2( us00_n5 ) );
  AOI221_X1 us00_U118 (.B1( us00_n12 ) , .C2( us00_n15 ) , .ZN( us00_n185 ) , .A( us00_n196 ) , .C1( us00_n35 ) , .B2( us00_n37 ) );
  INV_X1 us00_U119 (.A( us00_n198 ) , .ZN( us00_n5 ) );
  INV_X1 us00_U12 (.A( us00_n197 ) , .ZN( us00_n37 ) );
  NOR4_X1 us00_U120 (.ZN( us00_n186 ) , .A1( us00_n187 ) , .A2( us00_n188 ) , .A3( us00_n189 ) , .A4( us00_n190 ) );
  NAND4_X1 us00_U121 (.ZN( us00_n136 ) , .A2( us00_n156 ) , .A3( us00_n157 ) , .A4( us00_n158 ) , .A1( us00_n20 ) );
  INV_X1 us00_U122 (.A( us00_n168 ) , .ZN( us00_n20 ) );
  AOI221_X1 us00_U123 (.B1( us00_n15 ) , .ZN( us00_n156 ) , .C1( us00_n16 ) , .A( us00_n167 ) , .B2( us00_n32 ) , .C2( us00_n33 ) );
  NOR4_X1 us00_U124 (.ZN( us00_n158 ) , .A1( us00_n159 ) , .A2( us00_n160 ) , .A3( us00_n161 ) , .A4( us00_n162 ) );
  NAND4_X1 us00_U125 (.ZN( us00_n199 ) , .A1( us00_n401 ) , .A2( us00_n402 ) , .A3( us00_n403 ) , .A4( us00_n404 ) );
  NOR4_X1 us00_U126 (.A2( us00_n122 ) , .A1( us00_n142 ) , .A3( us00_n321 ) , .ZN( us00_n401 ) , .A4( us00_n407 ) );
  NOR4_X1 us00_U127 (.A2( us00_n235 ) , .A4( us00_n277 ) , .A3( us00_n309 ) , .A1( us00_n346 ) , .ZN( us00_n402 ) );
  NOR4_X1 us00_U128 (.A4( us00_n161 ) , .A2( us00_n294 ) , .A3( us00_n333 ) , .A1( us00_n371 ) , .ZN( us00_n403 ) );
  NOR2_X1 us00_U129 (.ZN( us00_n144 ) , .A1( us00_n32 ) , .A2( us00_n45 ) );
  NOR4_X1 us00_U13 (.ZN( us00_n171 ) , .A1( us00_n336 ) , .A2( us00_n361 ) , .A3( us00_n431 ) , .A4( us00_n432 ) );
  NOR2_X1 us00_U130 (.A2( us00_n15 ) , .ZN( us00_n88 ) , .A1( us00_n9 ) );
  NOR2_X1 us00_U131 (.A1( us00_n23 ) , .ZN( us00_n230 ) , .A2( us00_n9 ) );
  NAND4_X1 us00_U132 (.ZN( us00_n154 ) , .A2( us00_n3 ) , .A1( us00_n302 ) , .A3( us00_n303 ) , .A4( us00_n304 ) );
  NOR4_X1 us00_U133 (.ZN( us00_n304 ) , .A1( us00_n305 ) , .A2( us00_n306 ) , .A3( us00_n307 ) , .A4( us00_n308 ) );
  AOI221_X1 us00_U134 (.C1( us00_n24 ) , .B1( us00_n25 ) , .ZN( us00_n303 ) , .C2( us00_n312 ) , .A( us00_n313 ) , .B2( us00_n32 ) );
  INV_X1 us00_U135 (.A( us00_n270 ) , .ZN( us00_n3 ) );
  NAND4_X1 us00_U136 (.A2( us00_n10 ) , .A1( us00_n382 ) , .A3( us00_n383 ) , .A4( us00_n384 ) , .ZN( us00_n75 ) );
  AOI221_X1 us00_U137 (.B1( us00_n17 ) , .C1( us00_n26 ) , .C2( us00_n36 ) , .ZN( us00_n383 ) , .A( us00_n388 ) , .B2( us00_n41 ) );
  INV_X1 us00_U138 (.ZN( us00_n10 ) , .A( us00_n99 ) );
  NOR2_X1 us00_U139 (.A2( us00_n183 ) , .A1( us00_n199 ) , .ZN( us00_n382 ) );
  OR3_X1 us00_U14 (.A2( us00_n2 ) , .A3( us00_n300 ) , .A1( us00_n349 ) , .ZN( us00_n431 ) );
  INV_X1 us00_U140 (.A( us00_n115 ) , .ZN( us00_n47 ) );
  INV_X1 us00_U141 (.ZN( us00_n13 ) , .A( us00_n414 ) );
  OAI21_X1 us00_U142 (.B2( us00_n26 ) , .ZN( us00_n414 ) , .A( us00_n43 ) , .B1( us00_n68 ) );
  OR4_X1 us00_U143 (.A1( us00_n212 ) , .ZN( us00_n305 ) , .A2( us00_n309 ) , .A3( us00_n310 ) , .A4( us00_n311 ) );
  OR4_X1 us00_U144 (.ZN( us00_n355 ) , .A1( us00_n357 ) , .A2( us00_n358 ) , .A4( us00_n359 ) , .A3( us00_n56 ) );
  OR4_X1 us00_U145 (.A1( us00_n165 ) , .A2( us00_n299 ) , .A3( us00_n348 ) , .A4( us00_n359 ) , .ZN( us00_n411 ) );
  OR4_X1 us00_U146 (.ZN( us00_n187 ) , .A1( us00_n192 ) , .A2( us00_n193 ) , .A3( us00_n194 ) , .A4( us00_n195 ) );
  OR4_X1 us00_U147 (.ZN( us00_n293 ) , .A1( us00_n294 ) , .A2( us00_n295 ) , .A3( us00_n296 ) , .A4( us00_n297 ) );
  NAND2_X1 us00_U148 (.ZN( us00_n264 ) , .A1( us00_n4 ) , .A2( us00_n40 ) );
  OR3_X1 us00_U149 (.ZN( us00_n366 ) , .A1( us00_n369 ) , .A2( us00_n370 ) , .A3( us00_n371 ) );
  OR4_X1 us00_U15 (.A3( us00_n324 ) , .ZN( us00_n432 ) , .A1( us00_n433 ) , .A2( us00_n434 ) , .A4( us00_n435 ) );
  AOI221_X1 us00_U150 (.C2( us00_n14 ) , .ZN( us00_n157 ) , .B2( us00_n163 ) , .A( us00_n164 ) , .B1( us00_n38 ) , .C1( us00_n45 ) );
  OR2_X1 us00_U151 (.ZN( us00_n164 ) , .A1( us00_n165 ) , .A2( us00_n166 ) );
  INV_X1 us00_U152 (.A( us00_n123 ) , .ZN( us00_n8 ) );
  OAI21_X1 us00_U153 (.ZN( us00_n123 ) , .B1( us00_n124 ) , .A( us00_n32 ) , .B2( us00_n9 ) );
  INV_X1 us00_U154 (.ZN( us00_n18 ) , .A( us00_n205 ) );
  AOI21_X1 us00_U155 (.ZN( us00_n205 ) , .B1( us00_n206 ) , .A( us00_n207 ) , .B2( us00_n21 ) );
  NAND2_X1 us00_U156 (.ZN( us00_n128 ) , .A2( us00_n412 ) , .A1( us00_n430 ) );
  OAI222_X1 us00_U157 (.ZN( us00_n120 ) , .A2( us00_n128 ) , .B1( us00_n129 ) , .B2( us00_n130 ) , .A1( us00_n60 ) , .C1( us00_n63 ) , .C2( us00_n72 ) );
  OAI222_X1 us00_U158 (.A2( us00_n129 ) , .B1( us00_n130 ) , .B2( us00_n230 ) , .C2( us00_n252 ) , .ZN( us00_n372 ) , .A1( us00_n71 ) , .C1( us00_n72 ) );
  OAI222_X1 us00_U159 (.B1( us00_n130 ) , .C2( us00_n153 ) , .ZN( us00_n168 ) , .B2( us00_n169 ) , .A2( us00_n62 ) , .C1( us00_n63 ) , .A1( us00_n71 ) );
  INV_X1 us00_U16 (.ZN( us00_n2 ) , .A( us00_n264 ) );
  OAI222_X1 us00_U160 (.C2( us00_n130 ) , .C1( us00_n153 ) , .B1( us00_n180 ) , .ZN( us00_n260 ) , .A1( us00_n61 ) , .A2( us00_n85 ) , .B2( us00_n91 ) );
  NOR4_X1 us00_U161 (.A4( us00_n265 ) , .A3( us00_n297 ) , .ZN( us00_n384 ) , .A1( us00_n385 ) , .A2( us00_n386 ) );
  OR4_X1 us00_U162 (.A3( us00_n245 ) , .A1( us00_n318 ) , .A2( us00_n330 ) , .A4( us00_n343 ) , .ZN( us00_n385 ) );
  OAI22_X1 us00_U163 (.A2( us00_n114 ) , .A1( us00_n191 ) , .ZN( us00_n386 ) , .B1( us00_n387 ) , .B2( us00_n60 ) );
  NOR3_X1 us00_U164 (.A3( us00_n14 ) , .A2( us00_n27 ) , .ZN( us00_n387 ) , .A1( us00_n95 ) );
  AOI22_X1 us00_U165 (.A2( us00_n12 ) , .ZN( us00_n181 ) , .B2( us00_n34 ) , .A1( us00_n47 ) , .B1( us00_n9 ) );
  INV_X1 us00_U166 (.A( us00_n147 ) , .ZN( us00_n38 ) );
  AOI221_X1 us00_U167 (.B2( us00_n15 ) , .C1( us00_n25 ) , .C2( us00_n33 ) , .ZN( us00_n389 ) , .A( us00_n394 ) , .B1( us00_n46 ) );
  OAI22_X1 us00_U168 (.A1( us00_n169 ) , .ZN( us00_n394 ) , .B1( us00_n65 ) , .A2( us00_n71 ) , .B2( us00_n92 ) );
  INV_X1 us00_U169 (.ZN( us00_n45 ) , .A( us00_n87 ) );
  INV_X1 us00_U17 (.A( us00_n128 ) , .ZN( us00_n14 ) );
  NAND2_X1 us00_U170 (.ZN( us00_n115 ) , .A2( us00_n424 ) , .A1( us00_n426 ) );
  OAI22_X1 us00_U171 (.A2( us00_n115 ) , .B2( us00_n149 ) , .A1( us00_n178 ) , .ZN( us00_n240 ) , .B1( us00_n61 ) );
  OAI221_X1 us00_U172 (.ZN( us00_n140 ) , .B1( us00_n147 ) , .B2( us00_n148 ) , .C2( us00_n149 ) , .A( us00_n150 ) , .C1( us00_n60 ) );
  AOI22_X1 us00_U173 (.B2( us00_n11 ) , .A1( us00_n14 ) , .ZN( us00_n150 ) , .A2( us00_n39 ) , .B1( us00_n45 ) );
  INV_X1 us00_U174 (.ZN( us00_n15 ) , .A( us00_n91 ) );
  OAI22_X1 us00_U175 (.A1( us00_n133 ) , .B2( us00_n148 ) , .A2( us00_n149 ) , .ZN( us00_n167 ) , .B1( us00_n64 ) );
  INV_X1 us00_U176 (.ZN( us00_n46 ) , .A( us00_n61 ) );
  OAI22_X1 us00_U177 (.B1( us00_n147 ) , .B2( us00_n149 ) , .A1( us00_n153 ) , .ZN( us00_n388 ) , .A2( us00_n98 ) );
  OAI22_X1 us00_U178 (.B2( us00_n130 ) , .B1( us00_n208 ) , .ZN( us00_n253 ) , .A2( us00_n61 ) , .A1( us00_n62 ) );
  INV_X1 us00_U179 (.A( us00_n133 ) , .ZN( us00_n40 ) );
  AOI222_X1 us00_U18 (.B1( us00_n124 ) , .C1( us00_n14 ) , .A2( us00_n15 ) , .B2( us00_n206 ) , .ZN( us00_n272 ) , .A1( us00_n44 ) , .C2( us00_n46 ) );
  OAI22_X1 us00_U180 (.B2( us00_n127 ) , .ZN( us00_n151 ) , .A1( us00_n153 ) , .A2( us00_n61 ) , .B1( us00_n65 ) );
  OAI22_X1 us00_U181 (.A1( us00_n62 ) , .A2( us00_n63 ) , .ZN( us00_n96 ) , .B1( us00_n97 ) , .B2( us00_n98 ) );
  INV_X1 us00_U182 (.ZN( us00_n32 ) , .A( us00_n89 ) );
  INV_X1 us00_U183 (.ZN( us00_n17 ) , .A( us00_n72 ) );
  INV_X1 us00_U184 (.ZN( us00_n44 ) , .A( us00_n63 ) );
  OAI22_X1 us00_U185 (.A2( us00_n115 ) , .ZN( us00_n131 ) , .B2( us00_n133 ) , .A1( us00_n85 ) , .B1( us00_n97 ) );
  OAI22_X1 us00_U186 (.ZN( us00_n69 ) , .A1( us00_n71 ) , .A2( us00_n72 ) , .B1( us00_n73 ) , .B2( us00_n74 ) );
  INV_X1 us00_U187 (.ZN( us00_n12 ) , .A( us00_n208 ) );
  OAI22_X1 us00_U188 (.A2( us00_n133 ) , .ZN( us00_n381 ) , .B2( us00_n71 ) , .B1( us00_n86 ) , .A1( us00_n97 ) );
  INV_X1 us00_U189 (.A( us00_n127 ) , .ZN( us00_n35 ) );
  AOI222_X1 us00_U19 (.B2( us00_n14 ) , .A1( us00_n23 ) , .ZN( us00_n314 ) , .A2( us00_n34 ) , .C1( us00_n36 ) , .C2( us00_n4 ) , .B1( us00_n47 ) );
  OAI22_X1 us00_U190 (.B2( us00_n128 ) , .B1( us00_n147 ) , .ZN( us00_n287 ) , .A1( us00_n74 ) , .A2( us00_n91 ) );
  OAI22_X1 us00_U191 (.A2( us00_n147 ) , .ZN( us00_n182 ) , .B2( us00_n60 ) , .B1( us00_n86 ) , .A1( us00_n97 ) );
  INV_X1 us00_U192 (.ZN( us00_n34 ) , .A( us00_n74 ) );
  NOR2_X1 us00_U193 (.ZN( us00_n162 ) , .A2( us00_n60 ) , .A1( us00_n72 ) );
  NOR2_X1 us00_U194 (.ZN( us00_n107 ) , .A1( us00_n180 ) , .A2( us00_n62 ) );
  NOR2_X1 us00_U195 (.A1( us00_n149 ) , .ZN( us00_n211 ) , .A2( us00_n74 ) );
  NOR2_X1 us00_U196 (.A1( us00_n149 ) , .A2( us00_n180 ) , .ZN( us00_n283 ) );
  NOR2_X1 us00_U197 (.A1( us00_n149 ) , .ZN( us00_n307 ) , .A2( us00_n71 ) );
  NOR2_X1 us00_U198 (.ZN( us00_n122 ) , .A2( us00_n133 ) , .A1( us00_n72 ) );
  NOR2_X1 us00_U199 (.A1( us00_n133 ) , .A2( us00_n153 ) , .ZN( us00_n159 ) );
  AOI222_X1 us00_U20 (.C1( us00_n14 ) , .A1( us00_n17 ) , .ZN( us00_n217 ) , .C2( us00_n32 ) , .B1( us00_n36 ) , .A2( us00_n38 ) , .B2( us00_n7 ) );
  NOR2_X1 us00_U200 (.ZN( us00_n142 ) , .A1( us00_n72 ) , .A2( us00_n74 ) );
  NOR2_X1 us00_U201 (.ZN( us00_n331 ) , .A1( us00_n63 ) , .A2( us00_n97 ) );
  NOR2_X1 us00_U202 (.A2( us00_n178 ) , .ZN( us00_n300 ) , .A1( us00_n63 ) );
  NOR2_X1 us00_U203 (.A1( us00_n149 ) , .ZN( us00_n223 ) , .A2( us00_n64 ) );
  NOR2_X1 us00_U204 (.ZN( us00_n265 ) , .A2( us00_n91 ) , .A1( us00_n98 ) );
  NOR2_X1 us00_U205 (.A1( us00_n127 ) , .A2( us00_n128 ) , .ZN( us00_n345 ) );
  NOR2_X1 us00_U206 (.ZN( us00_n262 ) , .A2( us00_n62 ) , .A1( us00_n92 ) );
  NOR2_X1 us00_U207 (.A2( us00_n149 ) , .ZN( us00_n248 ) , .A1( us00_n92 ) );
  NOR2_X1 us00_U208 (.ZN( us00_n276 ) , .A1( us00_n74 ) , .A2( us00_n97 ) );
  NOR2_X1 us00_U209 (.ZN( us00_n266 ) , .A1( us00_n71 ) , .A2( us00_n97 ) );
  INV_X1 us00_U21 (.A( us00_n230 ) , .ZN( us00_n7 ) );
  INV_X1 us00_U210 (.A( us00_n130 ) , .ZN( us00_n43 ) );
  NOR2_X1 us00_U211 (.ZN( us00_n108 ) , .A2( us00_n133 ) , .A1( us00_n65 ) );
  NOR2_X1 us00_U212 (.A2( us00_n153 ) , .ZN( us00_n349 ) , .A1( us00_n74 ) );
  NOR2_X1 us00_U213 (.ZN( us00_n346 ) , .A1( us00_n61 ) , .A2( us00_n97 ) );
  NOR2_X1 us00_U214 (.A2( us00_n208 ) , .ZN( us00_n249 ) , .A1( us00_n92 ) );
  NOR2_X1 us00_U215 (.ZN( us00_n278 ) , .A1( us00_n61 ) , .A2( us00_n86 ) );
  INV_X1 us00_U216 (.A( us00_n149 ) , .ZN( us00_n25 ) );
  NOR2_X1 us00_U217 (.A1( us00_n208 ) , .ZN( us00_n225 ) , .A2( us00_n63 ) );
  NOR2_X1 us00_U218 (.A2( us00_n133 ) , .ZN( us00_n204 ) , .A1( us00_n208 ) );
  NOR2_X1 us00_U219 (.A1( us00_n208 ) , .ZN( us00_n275 ) , .A2( us00_n74 ) );
  NOR4_X1 us00_U22 (.A3( us00_n248 ) , .A1( us00_n268 ) , .A4( us00_n283 ) , .A2( us00_n356 ) , .ZN( us00_n404 ) );
  NOR2_X1 us00_U220 (.ZN( us00_n189 ) , .A1( us00_n208 ) , .A2( us00_n61 ) );
  INV_X1 us00_U221 (.ZN( us00_n26 ) , .A( us00_n85 ) );
  NOR2_X1 us00_U222 (.ZN( us00_n106 ) , .A1( us00_n127 ) , .A2( us00_n169 ) );
  NOR2_X1 us00_U223 (.ZN( us00_n111 ) , .A1( us00_n208 ) , .A2( us00_n64 ) );
  NOR2_X1 us00_U224 (.ZN( us00_n109 ) , .A1( us00_n178 ) , .A2( us00_n64 ) );
  NOR2_X1 us00_U225 (.A1( us00_n178 ) , .A2( us00_n180 ) , .ZN( us00_n336 ) );
  NOR2_X1 us00_U226 (.A1( us00_n208 ) , .ZN( us00_n350 ) , .A2( us00_n98 ) );
  NOR2_X1 us00_U227 (.A1( us00_n127 ) , .ZN( us00_n210 ) , .A2( us00_n62 ) );
  NOR2_X1 us00_U228 (.A1( us00_n127 ) , .ZN( us00_n322 ) , .A2( us00_n86 ) );
  NOR2_X1 us00_U229 (.ZN( us00_n369 ) , .A1( us00_n92 ) , .A2( us00_n97 ) );
  NOR4_X1 us00_U23 (.A2( us00_n247 ) , .A3( us00_n295 ) , .A4( us00_n320 ) , .A1( us00_n357 ) , .ZN( us00_n398 ) );
  NOR2_X1 us00_U230 (.A2( us00_n169 ) , .ZN( us00_n334 ) , .A1( us00_n92 ) );
  NOR2_X1 us00_U231 (.ZN( us00_n213 ) , .A2( us00_n86 ) , .A1( us00_n92 ) );
  NOR2_X1 us00_U232 (.ZN( us00_n161 ) , .A2( us00_n180 ) , .A1( us00_n85 ) );
  NOR2_X1 us00_U233 (.ZN( us00_n370 ) , .A2( us00_n60 ) , .A1( us00_n65 ) );
  NOR2_X1 us00_U234 (.A1( us00_n115 ) , .ZN( us00_n321 ) , .A2( us00_n72 ) );
  INV_X1 us00_U235 (.ZN( us00_n36 ) , .A( us00_n71 ) );
  NOR2_X1 us00_U236 (.A1( us00_n148 ) , .ZN( us00_n216 ) , .A2( us00_n87 ) );
  NOR2_X1 us00_U237 (.A1( us00_n148 ) , .A2( us00_n180 ) , .ZN( us00_n215 ) );
  NOR2_X1 us00_U238 (.ZN( us00_n320 ) , .A2( us00_n63 ) , .A1( us00_n85 ) );
  NOR2_X1 us00_U239 (.A1( us00_n128 ) , .ZN( us00_n332 ) , .A2( us00_n63 ) );
  NOR4_X1 us00_U24 (.ZN( us00_n342 ) , .A2( us00_n343 ) , .A3( us00_n344 ) , .A4( us00_n345 ) , .A1( us00_n57 ) );
  NOR2_X1 us00_U240 (.A1( us00_n148 ) , .ZN( us00_n368 ) , .A2( us00_n98 ) );
  NOR2_X1 us00_U241 (.A2( us00_n180 ) , .ZN( us00_n57 ) , .A1( us00_n97 ) );
  OAI22_X1 us00_U242 (.ZN( us00_n121 ) , .A1( us00_n125 ) , .B1( us00_n126 ) , .B2( us00_n127 ) , .A2( us00_n71 ) );
  NOR2_X1 us00_U243 (.ZN( us00_n126 ) , .A1( us00_n17 ) , .A2( us00_n25 ) );
  NOR3_X1 us00_U244 (.A3( us00_n12 ) , .ZN( us00_n125 ) , .A1( us00_n14 ) , .A2( us00_n24 ) );
  NOR2_X1 us00_U245 (.A2( us00_n133 ) , .ZN( us00_n347 ) , .A1( us00_n85 ) );
  NOR2_X1 us00_U246 (.ZN( us00_n110 ) , .A1( us00_n128 ) , .A2( us00_n74 ) );
  NOR2_X1 us00_U247 (.ZN( us00_n333 ) , .A1( us00_n85 ) , .A2( us00_n92 ) );
  NOR2_X1 us00_U248 (.A1( us00_n148 ) , .ZN( us00_n214 ) , .A2( us00_n92 ) );
  NOR2_X1 us00_U249 (.A1( us00_n153 ) , .ZN( us00_n246 ) , .A2( us00_n64 ) );
  NOR4_X1 us00_U25 (.A4( us00_n262 ) , .A3( us00_n298 ) , .A1( us00_n334 ) , .A2( us00_n360 ) , .ZN( us00_n421 ) );
  NOR2_X1 us00_U250 (.A1( us00_n115 ) , .ZN( us00_n263 ) , .A2( us00_n65 ) );
  OAI22_X1 us00_U251 (.B2( us00_n128 ) , .A1( us00_n133 ) , .A2( us00_n149 ) , .ZN( us00_n433 ) , .B1( us00_n437 ) );
  NOR3_X1 us00_U252 (.A1( us00_n31 ) , .A3( us00_n40 ) , .A2( us00_n41 ) , .ZN( us00_n437 ) );
  NOR2_X1 us00_U253 (.A1( us00_n115 ) , .A2( us00_n149 ) , .ZN( us00_n371 ) );
  NOR2_X1 us00_U254 (.A2( us00_n133 ) , .A1( us00_n169 ) , .ZN( us00_n361 ) );
  NOR2_X1 us00_U255 (.A2( us00_n133 ) , .ZN( us00_n160 ) , .A1( us00_n91 ) );
  NOR2_X1 us00_U256 (.ZN( us00_n323 ) , .A2( us00_n64 ) , .A1( us00_n91 ) );
  NOR2_X1 us00_U257 (.A1( us00_n169 ) , .ZN( us00_n360 ) , .A2( us00_n74 ) );
  NOR2_X1 us00_U258 (.A1( us00_n169 ) , .ZN( us00_n319 ) , .A2( us00_n61 ) );
  NOR2_X1 us00_U259 (.ZN( us00_n207 ) , .A2( us00_n72 ) , .A1( us00_n87 ) );
  NOR4_X1 us00_U26 (.A1( us00_n189 ) , .ZN( us00_n327 ) , .A2( us00_n334 ) , .A3( us00_n335 ) , .A4( us00_n336 ) );
  NOR2_X1 us00_U260 (.ZN( us00_n356 ) , .A2( us00_n65 ) , .A1( us00_n87 ) );
  NOR2_X1 us00_U261 (.A1( us00_n130 ) , .ZN( us00_n247 ) , .A2( us00_n62 ) );
  AOI21_X1 us00_U262 (.B2( us00_n180 ) , .ZN( us00_n306 ) , .A( us00_n65 ) , .B1( us00_n71 ) );
  NOR2_X1 us00_U263 (.ZN( us00_n222 ) , .A2( us00_n62 ) , .A1( us00_n87 ) );
  INV_X1 us00_U264 (.ZN( us00_n11 ) , .A( us00_n114 ) );
  AOI21_X1 us00_U265 (.A( us00_n180 ) , .B1( us00_n208 ) , .ZN( us00_n325 ) , .B2( us00_n72 ) );
  NOR2_X1 us00_U266 (.A2( us00_n169 ) , .ZN( us00_n209 ) , .A1( us00_n87 ) );
  NOR2_X1 us00_U267 (.A1( us00_n130 ) , .ZN( us00_n221 ) , .A2( us00_n97 ) );
  NOR2_X1 us00_U268 (.A1( us00_n115 ) , .ZN( us00_n335 ) , .A2( us00_n86 ) );
  NOR2_X1 us00_U269 (.ZN( us00_n176 ) , .A1( us00_n60 ) , .A2( us00_n91 ) );
  NOR2_X1 us00_U27 (.ZN( us00_n197 ) , .A1( us00_n38 ) , .A2( us00_n43 ) );
  NOR2_X1 us00_U270 (.A2( us00_n153 ) , .ZN( us00_n268 ) , .A1( us00_n60 ) );
  NOR2_X1 us00_U271 (.ZN( us00_n112 ) , .A1( us00_n147 ) , .A2( us00_n91 ) );
  AOI21_X1 us00_U272 (.ZN( us00_n59 ) , .B1( us00_n60 ) , .B2( us00_n61 ) , .A( us00_n62 ) );
  INV_X1 us00_U273 (.A( us00_n148 ) , .ZN( us00_n9 ) );
  NOR2_X1 us00_U274 (.A1( us00_n147 ) , .A2( us00_n169 ) , .ZN( us00_n298 ) );
  NOR2_X1 us00_U275 (.A1( us00_n147 ) , .A2( us00_n153 ) , .ZN( us00_n344 ) );
  AOI21_X1 us00_U276 (.A( us00_n114 ) , .ZN( us00_n250 ) , .B1( us00_n252 ) , .B2( us00_n63 ) );
  AOI21_X1 us00_U277 (.ZN( us00_n58 ) , .B1( us00_n63 ) , .B2( us00_n64 ) , .A( us00_n65 ) );
  AOI21_X1 us00_U278 (.B1( us00_n127 ) , .A( us00_n148 ) , .ZN( us00_n362 ) , .B2( us00_n74 ) );
  AOI21_X1 us00_U279 (.B1( us00_n197 ) , .ZN( us00_n378 ) , .B2( us00_n61 ) , .A( us00_n65 ) );
  AOI222_X1 us00_U28 (.B2( us00_n12 ) , .A2( us00_n22 ) , .C2( us00_n26 ) , .C1( us00_n35 ) , .A1( us00_n38 ) , .ZN( us00_n408 ) , .B1( us00_n45 ) );
  AOI21_X1 us00_U280 (.ZN( us00_n227 ) , .B2( us00_n72 ) , .B1( us00_n85 ) , .A( us00_n98 ) );
  AOI21_X1 us00_U281 (.A( us00_n128 ) , .B2( us00_n180 ) , .ZN( us00_n399 ) , .B1( us00_n98 ) );
  NOR2_X1 us00_U282 (.A1( us00_n133 ) , .ZN( us00_n295 ) , .A2( us00_n62 ) );
  NOR2_X1 us00_U283 (.ZN( us00_n235 ) , .A1( us00_n86 ) , .A2( us00_n89 ) );
  AOI21_X1 us00_U284 (.B1( us00_n127 ) , .ZN( us00_n284 ) , .B2( us00_n64 ) , .A( us00_n85 ) );
  NOR2_X1 us00_U285 (.A1( us00_n115 ) , .A2( us00_n169 ) , .ZN( us00_n83 ) );
  AOI21_X1 us00_U286 (.B2( us00_n208 ) , .ZN( us00_n251 ) , .B1( us00_n86 ) , .A( us00_n87 ) );
  NOR2_X1 us00_U287 (.A2( us00_n169 ) , .ZN( us00_n357 ) , .A1( us00_n63 ) );
  AOI21_X1 us00_U288 (.B1( us00_n127 ) , .A( us00_n208 ) , .ZN( us00_n400 ) , .B2( us00_n71 ) );
  NOR2_X1 us00_U289 (.ZN( us00_n318 ) , .A1( us00_n74 ) , .A2( us00_n86 ) );
  NOR4_X1 us00_U29 (.A3( us00_n263 ) , .A2( us00_n323 ) , .A4( us00_n335 ) , .ZN( us00_n410 ) , .A1( us00_n411 ) );
  NOR2_X1 us00_U290 (.A2( us00_n178 ) , .ZN( us00_n358 ) , .A1( us00_n61 ) );
  NOR2_X1 us00_U291 (.A2( us00_n178 ) , .ZN( us00_n194 ) , .A1( us00_n74 ) );
  NOR2_X1 us00_U292 (.A1( us00_n115 ) , .ZN( us00_n224 ) , .A2( us00_n91 ) );
  INV_X1 us00_U293 (.ZN( us00_n41 ) , .A( us00_n64 ) );
  AOI21_X1 us00_U294 (.A( us00_n147 ) , .B2( us00_n208 ) , .ZN( us00_n367 ) , .B1( us00_n62 ) );
  AOI21_X1 us00_U295 (.ZN( us00_n338 ) , .B1( us00_n62 ) , .A( us00_n63 ) , .B2( us00_n65 ) );
  AOI21_X1 us00_U296 (.A( us00_n114 ) , .ZN( us00_n337 ) , .B1( us00_n60 ) , .B2( us00_n98 ) );
  NOR2_X1 us00_U297 (.A1( us00_n208 ) , .ZN( us00_n296 ) , .A2( us00_n89 ) );
  AOI21_X1 us00_U298 (.B2( us00_n178 ) , .ZN( us00_n288 ) , .A( us00_n60 ) , .B1( us00_n62 ) );
  AOI21_X1 us00_U299 (.B2( us00_n114 ) , .A( us00_n145 ) , .ZN( us00_n177 ) , .B1( us00_n178 ) );
  NAND2_X1 us00_U3 (.ZN( us00_n169 ) , .A2( us00_n413 ) , .A1( us00_n436 ) );
  AOI221_X1 us00_U30 (.A( us00_n13 ) , .C2( us00_n163 ) , .B1( us00_n17 ) , .C1( us00_n32 ) , .ZN( us00_n409 ) , .B2( us00_n46 ) );
  AOI21_X1 us00_U300 (.B2( us00_n114 ) , .ZN( us00_n286 ) , .B1( us00_n65 ) , .A( us00_n92 ) );
  AOI21_X1 us00_U301 (.B2( us00_n115 ) , .A( us00_n153 ) , .ZN( us00_n379 ) , .B1( us00_n63 ) );
  NOR2_X1 us00_U302 (.A2( us00_n133 ) , .A1( us00_n178 ) , .ZN( us00_n330 ) );
  INV_X1 us00_U303 (.ZN( us00_n4 ) , .A( us00_n86 ) );
  INV_X1 us00_U304 (.ZN( us00_n23 ) , .A( us00_n65 ) );
  AOI21_X1 us00_U305 (.B2( us00_n130 ) , .ZN( us00_n237 ) , .B1( us00_n74 ) , .A( us00_n85 ) );
  AOI21_X1 us00_U306 (.B2( us00_n114 ) , .B1( us00_n148 ) , .ZN( us00_n228 ) , .A( us00_n64 ) );
  NOR2_X1 us00_U307 (.A1( us00_n148 ) , .ZN( us00_n192 ) , .A2( us00_n61 ) );
  AOI21_X1 us00_U308 (.B2( us00_n116 ) , .A( us00_n149 ) , .ZN( us00_n190 ) , .B1( us00_n191 ) );
  AOI21_X1 us00_U309 (.B2( us00_n115 ) , .B1( us00_n127 ) , .ZN( us00_n308 ) , .A( us00_n97 ) );
  NOR4_X1 us00_U31 (.ZN( us00_n353 ) , .A1( us00_n360 ) , .A2( us00_n361 ) , .A3( us00_n362 ) , .A4( us00_n363 ) );
  AOI21_X1 us00_U310 (.B1( us00_n169 ) , .A( us00_n180 ) , .ZN( us00_n377 ) , .B2( us00_n91 ) );
  NOR2_X1 us00_U311 (.A2( us00_n115 ) , .A1( us00_n148 ) , .ZN( us00_n309 ) );
  NOR2_X1 us00_U312 (.A2( us00_n180 ) , .ZN( us00_n297 ) , .A1( us00_n86 ) );
  NOR2_X1 us00_U313 (.A1( us00_n114 ) , .A2( us00_n180 ) , .ZN( us00_n311 ) );
  AOI21_X1 us00_U314 (.ZN( us00_n363 ) , .B1( us00_n65 ) , .B2( us00_n85 ) , .A( us00_n98 ) );
  AOI21_X1 us00_U315 (.B2( us00_n128 ) , .ZN( us00_n238 ) , .B1( us00_n65 ) , .A( us00_n89 ) );
  INV_X1 us00_U316 (.A( us00_n178 ) , .ZN( us00_n24 ) );
  NOR2_X1 us00_U317 (.ZN( us00_n212 ) , .A2( us00_n64 ) , .A1( us00_n97 ) );
  AOI21_X1 us00_U318 (.ZN( us00_n427 ) , .B1( us00_n62 ) , .A( us00_n74 ) , .B2( us00_n85 ) );
  NOR2_X1 us00_U319 (.A1( us00_n153 ) , .A2( us00_n180 ) , .ZN( us00_n245 ) );
  AOI222_X1 us00_U32 (.B1( us00_n11 ) , .A2( us00_n25 ) , .C2( us00_n27 ) , .C1( us00_n33 ) , .ZN( us00_n352 ) , .B2( us00_n40 ) , .A1( us00_n43 ) );
  AOI21_X1 us00_U320 (.B1( us00_n153 ) , .ZN( us00_n313 ) , .B2( us00_n86 ) , .A( us00_n98 ) );
  AOI21_X1 us00_U321 (.ZN( us00_n380 ) , .B1( us00_n73 ) , .B2( us00_n86 ) , .A( us00_n98 ) );
  NAND2_X1 us00_U322 (.A1( us00_n114 ) , .ZN( us00_n124 ) , .A2( us00_n72 ) );
  NOR2_X1 us00_U323 (.A1( us00_n169 ) , .ZN( us00_n348 ) , .A2( us00_n98 ) );
  NOR2_X1 us00_U324 (.A1( us00_n169 ) , .ZN( us00_n299 ) , .A2( us00_n64 ) );
  AOI21_X1 us00_U325 (.B1( us00_n114 ) , .B2( us00_n128 ) , .ZN( us00_n188 ) , .A( us00_n71 ) );
  NOR2_X1 us00_U326 (.A1( us00_n130 ) , .ZN( us00_n310 ) , .A2( us00_n72 ) );
  NOR2_X1 us00_U327 (.ZN( us00_n193 ) , .A2( us00_n64 ) , .A1( us00_n86 ) );
  NOR2_X1 us00_U328 (.ZN( us00_n56 ) , .A1( us00_n62 ) , .A2( us00_n64 ) );
  AOI21_X1 us00_U329 (.ZN( us00_n84 ) , .B1( us00_n85 ) , .B2( us00_n86 ) , .A( us00_n87 ) );
  NOR4_X1 us00_U33 (.A4( us00_n108 ) , .A2( us00_n204 ) , .ZN( us00_n354 ) , .A1( us00_n355 ) , .A3( us00_n356 ) );
  AOI21_X1 us00_U330 (.ZN( us00_n143 ) , .A( us00_n144 ) , .B1( us00_n85 ) , .B2( us00_n97 ) );
  AOI21_X1 us00_U331 (.B1( us00_n197 ) , .ZN( us00_n236 ) , .B2( us00_n60 ) , .A( us00_n86 ) );
  NOR2_X1 us00_U332 (.A2( us00_n114 ) , .A1( us00_n115 ) , .ZN( us00_n166 ) );
  NOR2_X1 us00_U333 (.ZN( us00_n294 ) , .A2( us00_n60 ) , .A1( us00_n85 ) );
  NOR2_X1 us00_U334 (.A1( us00_n153 ) , .ZN( us00_n343 ) , .A2( us00_n89 ) );
  NOR2_X1 us00_U335 (.A2( us00_n169 ) , .ZN( us00_n195 ) , .A1( us00_n60 ) );
  INV_X1 us00_U336 (.A( us00_n180 ) , .ZN( us00_n39 ) );
  INV_X1 us00_U337 (.ZN( us00_n22 ) , .A( us00_n62 ) );
  AOI21_X1 us00_U338 (.B2( us00_n127 ) , .B1( us00_n144 ) , .A( us00_n178 ) , .ZN( us00_n435 ) );
  OAI21_X1 us00_U339 (.B2( us00_n127 ) , .ZN( us00_n175 ) , .A( us00_n179 ) , .B1( us00_n73 ) );
  NOR4_X1 us00_U34 (.ZN( us00_n139 ) , .A1( us00_n140 ) , .A2( us00_n141 ) , .A3( us00_n142 ) , .A4( us00_n143 ) );
  OAI21_X1 us00_U340 (.A( us00_n17 ) , .ZN( us00_n179 ) , .B1( us00_n39 ) , .B2( us00_n44 ) );
  INV_X1 us00_U341 (.ZN( us00_n27 ) , .A( us00_n97 ) );
  INV_X1 us00_U342 (.ZN( us00_n31 ) , .A( us00_n92 ) );
  AOI22_X1 us00_U343 (.B1( us00_n14 ) , .A1( us00_n43 ) , .B2( us00_n46 ) , .ZN( us00_n94 ) , .A2( us00_n95 ) );
  NAND2_X1 us00_U344 (.ZN( us00_n206 ) , .A2( us00_n61 ) , .A1( us00_n71 ) );
  NAND2_X1 us00_U345 (.A1( us00_n149 ) , .ZN( us00_n163 ) , .A2( us00_n97 ) );
  NAND2_X1 us00_U346 (.A2( us00_n115 ) , .ZN( us00_n67 ) , .A1( us00_n71 ) );
  AOI21_X1 us00_U347 (.ZN( us00_n434 ) , .A( us00_n63 ) , .B2( us00_n86 ) , .B1( us00_n88 ) );
  NOR2_X1 us00_U348 (.ZN( us00_n393 ) , .A2( us00_n72 ) , .A1( us00_n89 ) );
  NOR2_X1 us00_U349 (.ZN( us00_n407 ) , .A1( us00_n62 ) , .A2( us00_n98 ) );
  AOI211_X1 us00_U35 (.ZN( us00_n138 ) , .A( us00_n151 ) , .B( us00_n152 ) , .C2( us00_n22 ) , .C1( us00_n34 ) );
  OAI21_X1 us00_U350 (.ZN( us00_n82 ) , .B1( us00_n88 ) , .B2( us00_n89 ) , .A( us00_n90 ) );
  OAI21_X1 us00_U351 (.B1( us00_n14 ) , .A( us00_n38 ) , .B2( us00_n4 ) , .ZN( us00_n90 ) );
  NOR2_X1 us00_U352 (.A2( us00_n153 ) , .ZN( us00_n165 ) , .A1( us00_n87 ) );
  NOR2_X1 us00_U353 (.A2( us00_n127 ) , .A1( us00_n153 ) , .ZN( us00_n351 ) );
  NAND2_X1 us00_U354 (.A2( us00_n148 ) , .A1( us00_n178 ) , .ZN( us00_n95 ) );
  NOR2_X1 us00_U355 (.A1( us00_n169 ) , .ZN( us00_n359 ) , .A2( us00_n89 ) );
  OAI21_X1 us00_U356 (.ZN( us00_n141 ) , .B1( us00_n145 ) , .A( us00_n146 ) , .B2( us00_n72 ) );
  OAI21_X1 us00_U357 (.ZN( us00_n146 ) , .B2( us00_n25 ) , .B1( us00_n4 ) , .A( us00_n44 ) );
  NAND2_X1 us00_U358 (.A2( us00_n128 ) , .ZN( us00_n68 ) , .A1( us00_n91 ) );
  INV_X1 us00_U359 (.ZN( us00_n33 ) , .A( us00_n60 ) );
  NOR3_X1 us00_U36 (.A2( us00_n136 ) , .ZN( us00_n137 ) , .A1( us00_n154 ) , .A3( us00_n155 ) );
  INV_X1 us00_U360 (.A( us00_n153 ) , .ZN( us00_n21 ) );
  AND2_X1 us00_U361 (.ZN( us00_n145 ) , .A2( us00_n92 ) , .A1( us00_n98 ) );
  AOI221_X1 us00_U362 (.ZN( us00_n103 ) , .B1( us00_n11 ) , .A( us00_n113 ) , .C1( us00_n22 ) , .B2( us00_n42 ) , .C2( us00_n67 ) );
  AOI21_X1 us00_U363 (.ZN( us00_n113 ) , .B2( us00_n114 ) , .B1( us00_n85 ) , .A( us00_n89 ) );
  INV_X1 us00_U364 (.A( us00_n116 ) , .ZN( us00_n42 ) );
  NAND2_X1 us00_U365 (.A2( us00_n428 ) , .A1( us00_n430 ) , .ZN( us00_n72 ) );
  NAND2_X1 us00_U366 (.A2( us00_n406 ) , .A1( us00_n422 ) , .ZN( us00_n74 ) );
  NAND2_X1 us00_U367 (.A2( us00_n423 ) , .A1( us00_n426 ) , .ZN( us00_n63 ) );
  NAND2_X1 us00_U368 (.A2( us00_n406 ) , .A1( us00_n426 ) , .ZN( us00_n61 ) );
  NAND2_X1 us00_U369 (.A2( us00_n416 ) , .A1( us00_n423 ) , .ZN( us00_n64 ) );
  NOR4_X1 us00_U37 (.ZN( us00_n119 ) , .A1( us00_n120 ) , .A2( us00_n121 ) , .A3( us00_n122 ) , .A4( us00_n8 ) );
  NAND2_X1 us00_U370 (.ZN( us00_n133 ) , .A2( us00_n416 ) , .A1( us00_n424 ) );
  NAND2_X1 us00_U371 (.ZN( us00_n208 ) , .A2( us00_n412 ) , .A1( us00_n425 ) );
  NAND2_X1 us00_U372 (.ZN( us00_n149 ) , .A1( us00_n417 ) , .A2( us00_n429 ) );
  NAND2_X1 us00_U373 (.ZN( us00_n127 ) , .A2( us00_n415 ) , .A1( us00_n422 ) );
  NAND2_X1 us00_U374 (.A1( us00_n422 ) , .A2( us00_n424 ) , .ZN( us00_n71 ) );
  NAND2_X1 us00_U375 (.A1( us00_n405 ) , .A2( us00_n423 ) , .ZN( us00_n98 ) );
  NAND2_X1 us00_U376 (.A2( us00_n405 ) , .A1( us00_n424 ) , .ZN( us00_n92 ) );
  NAND2_X1 us00_U377 (.A1( us00_n412 ) , .A2( us00_n413 ) , .ZN( us00_n65 ) );
  NAND2_X1 us00_U378 (.ZN( us00_n178 ) , .A2( us00_n417 ) , .A1( us00_n436 ) );
  NAND2_X1 us00_U379 (.ZN( us00_n114 ) , .A1( us00_n425 ) , .A2( us00_n428 ) );
  AOI211_X1 us00_U38 (.ZN( us00_n118 ) , .A( us00_n131 ) , .B( us00_n132 ) , .C2( us00_n24 ) , .C1( us00_n45 ) );
  NAND2_X2 us00_U380 (.ZN( us00_n180 ) , .A1( us00_n406 ) , .A2( us00_n416 ) );
  NAND2_X1 us00_U381 (.ZN( us00_n148 ) , .A1( us00_n425 ) , .A2( us00_n429 ) );
  NAND2_X1 us00_U382 (.ZN( us00_n130 ) , .A1( us00_n415 ) , .A2( us00_n416 ) );
  NAND2_X1 us00_U383 (.A2( us00_n405 ) , .A1( us00_n415 ) , .ZN( us00_n89 ) );
  NOR2_X1 us00_U384 (.A1( us00_n29 ) , .A2( us00_n30 ) , .ZN( us00_n412 ) );
  NOR2_X1 us00_U385 (.ZN( us00_n424 ) , .A2( us00_n50 ) , .A1( us00_n51 ) );
  NOR2_X1 us00_U386 (.ZN( us00_n426 ) , .A2( us00_n48 ) , .A1( us00_n49 ) );
  NOR2_X1 us00_U387 (.A1( us00_n19 ) , .A2( us00_n28 ) , .ZN( us00_n430 ) );
  NAND2_X1 us00_U388 (.ZN( us00_n147 ) , .A1( us00_n422 ) , .A2( us00_n423 ) );
  NAND2_X1 us00_U389 (.A2( us00_n415 ) , .A1( us00_n426 ) , .ZN( us00_n87 ) );
  NOR3_X1 us00_U39 (.ZN( us00_n117 ) , .A1( us00_n134 ) , .A2( us00_n135 ) , .A3( us00_n136 ) );
  NAND2_X2 us00_U390 (.A1( us00_n413 ) , .A2( us00_n429 ) , .ZN( us00_n62 ) );
  NAND2_X2 us00_U391 (.A1( us00_n425 ) , .A2( us00_n436 ) , .ZN( us00_n86 ) );
  NAND2_X2 us00_U392 (.ZN( us00_n153 ) , .A2( us00_n413 ) , .A1( us00_n428 ) );
  NAND2_X1 us00_U393 (.A1( us00_n430 ) , .A2( us00_n436 ) , .ZN( us00_n93 ) );
  NAND2_X2 us00_U394 (.A2( us00_n417 ) , .A1( us00_n428 ) , .ZN( us00_n85 ) );
  NAND2_X2 us00_U395 (.A1( us00_n412 ) , .A2( us00_n417 ) , .ZN( us00_n97 ) );
  NAND2_X1 us00_U396 (.A2( us00_n429 ) , .A1( us00_n430 ) , .ZN( us00_n91 ) );
  NOR2_X1 us00_U397 (.A2( sa00_6 ) , .A1( sa00_7 ) , .ZN( us00_n413 ) );
  NOR2_X1 us00_U398 (.A2( sa00_5 ) , .A1( us00_n30 ) , .ZN( us00_n429 ) );
  NOR2_X1 us00_U399 (.A2( sa00_7 ) , .A1( us00_n28 ) , .ZN( us00_n417 ) );
  NAND2_X1 us00_U4 (.A1( us00_n405 ) , .A2( us00_n406 ) , .ZN( us00_n60 ) );
  AOI221_X1 us00_U40 (.C1( us00_n11 ) , .B1( us00_n12 ) , .B2( us00_n39 ) , .C2( us00_n40 ) , .ZN( us00_n79 ) , .A( us00_n96 ) );
  NOR2_X1 us00_U400 (.A2( sa00_4 ) , .A1( us00_n29 ) , .ZN( us00_n428 ) );
  NOR2_X1 us00_U401 (.A2( sa00_4 ) , .A1( sa00_5 ) , .ZN( us00_n436 ) );
  NOR2_X1 us00_U402 (.A2( sa00_1 ) , .ZN( us00_n406 ) , .A1( us00_n51 ) );
  NOR2_X1 us00_U403 (.A2( sa00_2 ) , .A1( sa00_3 ) , .ZN( us00_n405 ) );
  NOR2_X1 us00_U404 (.A2( sa00_6 ) , .A1( us00_n19 ) , .ZN( us00_n425 ) );
  NOR2_X1 us00_U405 (.A2( sa00_2 ) , .ZN( us00_n416 ) , .A1( us00_n48 ) );
  NOR2_X1 us00_U406 (.A2( sa00_0 ) , .ZN( us00_n423 ) , .A1( us00_n50 ) );
  NOR2_X1 us00_U407 (.A2( sa00_0 ) , .A1( sa00_1 ) , .ZN( us00_n415 ) );
  NOR2_X1 us00_U408 (.A2( sa00_3 ) , .ZN( us00_n422 ) , .A1( us00_n49 ) );
  INV_X1 us00_U409 (.A( sa00_6 ) , .ZN( us00_n28 ) );
  NOR4_X1 us00_U41 (.ZN( us00_n80 ) , .A1( us00_n81 ) , .A2( us00_n82 ) , .A3( us00_n83 ) , .A4( us00_n84 ) );
  INV_X1 us00_U410 (.A( sa00_1 ) , .ZN( us00_n50 ) );
  INV_X1 us00_U411 (.A( sa00_3 ) , .ZN( us00_n48 ) );
  INV_X1 us00_U412 (.A( sa00_2 ) , .ZN( us00_n49 ) );
  INV_X1 us00_U413 (.A( sa00_0 ) , .ZN( us00_n51 ) );
  INV_X1 us00_U414 (.A( sa00_5 ) , .ZN( us00_n29 ) );
  INV_X1 us00_U415 (.A( sa00_7 ) , .ZN( us00_n19 ) );
  OAI221_X1 us00_U416 (.C1( us00_n64 ) , .ZN( us00_n81 ) , .B1( us00_n91 ) , .B2( us00_n92 ) , .C2( us00_n93 ) , .A( us00_n94 ) );
  NAND2_X1 us00_U417 (.A1( us00_n148 ) , .ZN( us00_n66 ) , .A2( us00_n93 ) );
  OAI22_X1 us00_U418 (.A1( us00_n114 ) , .B2( us00_n115 ) , .A2( us00_n130 ) , .ZN( us00_n289 ) , .B1( us00_n93 ) );
  OAI221_X1 us00_U419 (.ZN( us00_n174 ) , .A( us00_n181 ) , .B2( us00_n71 ) , .B1( us00_n91 ) , .C1( us00_n92 ) , .C2( us00_n93 ) );
  NOR4_X1 us00_U42 (.A3( us00_n100 ) , .A4( us00_n101 ) , .A2( us00_n76 ) , .ZN( us00_n78 ) , .A1( us00_n99 ) );
  AOI21_X1 us00_U420 (.B1( us00_n149 ) , .ZN( us00_n285 ) , .A( us00_n87 ) , .B2( us00_n93 ) );
  AOI21_X1 us00_U421 (.B1( us00_n178 ) , .ZN( us00_n254 ) , .B2( us00_n93 ) , .A( us00_n98 ) );
  AOI21_X1 us00_U422 (.A( us00_n115 ) , .ZN( us00_n229 ) , .B1( us00_n85 ) , .B2( us00_n93 ) );
  OAI22_X1 us00_U423 (.A2( us00_n147 ) , .A1( us00_n178 ) , .ZN( us00_n196 ) , .B1( us00_n60 ) , .B2( us00_n93 ) );
  OAI21_X1 us00_U424 (.B1( us00_n252 ) , .ZN( us00_n261 ) , .A( us00_n264 ) , .B2( us00_n93 ) );
  NOR2_X1 us00_U425 (.ZN( us00_n267 ) , .A2( us00_n61 ) , .A1( us00_n93 ) );
  OAI222_X1 us00_U426 (.B1( us00_n130 ) , .ZN( us00_n203 ) , .A2( us00_n208 ) , .A1( us00_n60 ) , .C1( us00_n62 ) , .C2( us00_n89 ) , .B2( us00_n93 ) );
  NOR2_X1 us00_U427 (.ZN( us00_n226 ) , .A2( us00_n89 ) , .A1( us00_n93 ) );
  NOR2_X1 us00_U428 (.A2( us00_n180 ) , .ZN( us00_n277 ) , .A1( us00_n93 ) );
  NOR2_X1 us00_U429 (.A2( us00_n133 ) , .ZN( us00_n324 ) , .A1( us00_n93 ) );
  NOR2_X1 us00_U43 (.A2( us00_n16 ) , .A1( us00_n23 ) , .ZN( us00_n73 ) );
  INV_X1 us00_U430 (.ZN( us00_n16 ) , .A( us00_n93 ) );
  NAND4_X1 us00_U431 (.ZN( sa00_sr_2 ) , .A2( us00_n231 ) , .A1( us00_n232 ) , .A3( us00_n233 ) , .A4( us00_n234 ) );
  AOI221_X1 us00_U432 (.C1( us00_n16 ) , .B1( us00_n23 ) , .ZN( us00_n290 ) , .A( us00_n301 ) , .C2( us00_n34 ) , .B2( us00_n46 ) );
  AOI21_X1 us00_U433 (.B1( us00_n129 ) , .B2( us00_n153 ) , .ZN( us00_n301 ) , .A( us00_n92 ) );
  AOI211_X1 us00_U434 (.B( us00_n134 ) , .C1( us00_n23 ) , .ZN( us00_n232 ) , .A( us00_n240 ) , .C2( us00_n38 ) );
  NAND4_X1 us00_U435 (.ZN( us00_n134 ) , .A1( us00_n241 ) , .A2( us00_n242 ) , .A3( us00_n243 ) , .A4( us00_n244 ) );
  INV_X1 us00_U436 (.A( sa00_4 ) , .ZN( us00_n30 ) );
  NAND3_X1 us00_U437 (.ZN( sa00_sr_6 ) , .A1( us00_n78 ) , .A2( us00_n79 ) , .A3( us00_n80 ) );
  NAND3_X1 us00_U438 (.ZN( sa00_sr_5 ) , .A1( us00_n117 ) , .A2( us00_n118 ) , .A3( us00_n119 ) );
  NAND3_X1 us00_U439 (.ZN( sa00_sr_4 ) , .A1( us00_n137 ) , .A2( us00_n138 ) , .A3( us00_n139 ) );
  NAND4_X1 us00_U44 (.ZN( sa00_sr_3 ) , .A1( us00_n170 ) , .A2( us00_n171 ) , .A3( us00_n172 ) , .A4( us00_n173 ) );
  NAND3_X1 us00_U440 (.A1( us00_n200 ) , .A2( us00_n201 ) , .A3( us00_n202 ) , .ZN( us00_n70 ) );
  NAND3_X1 us00_U441 (.A2( us00_n153 ) , .A3( us00_n169 ) , .ZN( us00_n239 ) , .A1( us00_n85 ) );
  NAND3_X1 us00_U442 (.ZN( us00_n152 ) , .A1( us00_n257 ) , .A2( us00_n258 ) , .A3( us00_n259 ) );
  NAND3_X1 us00_U443 (.ZN( us00_n256 ) , .A1( us00_n290 ) , .A2( us00_n291 ) , .A3( us00_n292 ) );
  NAND3_X1 us00_U444 (.A2( us00_n127 ) , .A3( us00_n197 ) , .ZN( us00_n312 ) , .A1( us00_n92 ) );
  NAND3_X1 us00_U445 (.ZN( us00_n135 ) , .A1( us00_n352 ) , .A2( us00_n353 ) , .A3( us00_n354 ) );
  NAND3_X1 us00_U446 (.ZN( us00_n269 ) , .A1( us00_n364 ) , .A3( us00_n365 ) , .A2( us00_n6 ) );
  NAND3_X1 us00_U447 (.ZN( us00_n100 ) , .A1( us00_n408 ) , .A2( us00_n409 ) , .A3( us00_n410 ) );
  NOR4_X1 us00_U45 (.ZN( us00_n173 ) , .A1( us00_n174 ) , .A2( us00_n175 ) , .A3( us00_n176 ) , .A4( us00_n177 ) );
  AOI211_X1 us00_U46 (.ZN( us00_n172 ) , .A( us00_n182 ) , .B( us00_n183 ) , .C1( us00_n26 ) , .C2( us00_n46 ) );
  NOR2_X1 us00_U47 (.A2( us00_n101 ) , .ZN( us00_n170 ) , .A1( us00_n77 ) );
  NAND4_X1 us00_U48 (.ZN( sa00_sr_7 ) , .A1( us00_n52 ) , .A2( us00_n53 ) , .A3( us00_n54 ) , .A4( us00_n55 ) );
  NOR4_X1 us00_U49 (.ZN( us00_n55 ) , .A1( us00_n56 ) , .A2( us00_n57 ) , .A3( us00_n58 ) , .A4( us00_n59 ) );
  NOR3_X1 us00_U5 (.A2( us00_n135 ) , .A3( us00_n154 ) , .A1( us00_n269 ) , .ZN( us00_n279 ) );
  AOI222_X1 us00_U50 (.B1( us00_n24 ) , .A1( us00_n38 ) , .C1( us00_n45 ) , .ZN( us00_n54 ) , .A2( us00_n66 ) , .B2( us00_n67 ) , .C2( us00_n68 ) );
  AOI211_X1 us00_U51 (.C2( us00_n27 ) , .C1( us00_n35 ) , .ZN( us00_n53 ) , .A( us00_n69 ) , .B( us00_n70 ) );
  NOR2_X1 us00_U52 (.ZN( us00_n129 ) , .A2( us00_n15 ) , .A1( us00_n16 ) );
  NAND4_X1 us00_U53 (.ZN( sa00_sr_0 ) , .A1( us00_n373 ) , .A2( us00_n374 ) , .A3( us00_n375 ) , .A4( us00_n376 ) );
  AOI221_X1 us00_U54 (.B1( us00_n15 ) , .C2( us00_n17 ) , .C1( us00_n31 ) , .B2( us00_n34 ) , .ZN( us00_n375 ) , .A( us00_n380 ) );
  NOR4_X1 us00_U55 (.A1( us00_n350 ) , .ZN( us00_n376 ) , .A2( us00_n377 ) , .A3( us00_n378 ) , .A4( us00_n379 ) );
  AOI211_X1 us00_U56 (.C1( us00_n26 ) , .ZN( us00_n374 ) , .C2( us00_n38 ) , .A( us00_n381 ) , .B( us00_n75 ) );
  NAND4_X1 us00_U57 (.ZN( sa00_sr_1 ) , .A1( us00_n279 ) , .A2( us00_n280 ) , .A3( us00_n281 ) , .A4( us00_n282 ) );
  NOR4_X1 us00_U58 (.ZN( us00_n282 ) , .A1( us00_n283 ) , .A2( us00_n284 ) , .A3( us00_n285 ) , .A4( us00_n286 ) );
  AOI211_X1 us00_U59 (.ZN( us00_n281 ) , .A( us00_n287 ) , .B( us00_n288 ) , .C1( us00_n44 ) , .C2( us00_n66 ) );
  NOR3_X1 us00_U6 (.ZN( us00_n52 ) , .A1( us00_n75 ) , .A2( us00_n76 ) , .A3( us00_n77 ) );
  AOI211_X1 us00_U60 (.C2( us00_n22 ) , .B( us00_n256 ) , .ZN( us00_n280 ) , .A( us00_n289 ) , .C1( us00_n32 ) );
  NOR2_X1 us00_U61 (.ZN( us00_n252 ) , .A1( us00_n38 ) , .A2( us00_n41 ) );
  NAND4_X1 us00_U62 (.ZN( us00_n155 ) , .A1( us00_n271 ) , .A2( us00_n272 ) , .A3( us00_n273 ) , .A4( us00_n274 ) );
  NOR3_X1 us00_U63 (.A2( us00_n107 ) , .A3( us00_n214 ) , .ZN( us00_n273 ) , .A1( us00_n278 ) );
  NOR4_X1 us00_U64 (.A4( us00_n222 ) , .ZN( us00_n274 ) , .A1( us00_n275 ) , .A2( us00_n276 ) , .A3( us00_n277 ) );
  AOI222_X1 us00_U65 (.B2( us00_n16 ) , .A2( us00_n21 ) , .ZN( us00_n271 ) , .B1( us00_n35 ) , .C2( us00_n40 ) , .A1( us00_n47 ) , .C1( us00_n9 ) );
  NOR4_X1 us00_U66 (.A1( us00_n194 ) , .ZN( us00_n291 ) , .A2( us00_n298 ) , .A3( us00_n299 ) , .A4( us00_n300 ) );
  NOR4_X1 us00_U67 (.A4( us00_n110 ) , .A2( us00_n215 ) , .A3( us00_n225 ) , .ZN( us00_n292 ) , .A1( us00_n293 ) );
  AOI211_X1 us00_U68 (.C1( us00_n14 ) , .ZN( us00_n242 ) , .A( us00_n253 ) , .B( us00_n254 ) , .C2( us00_n41 ) );
  NOR4_X1 us00_U69 (.ZN( us00_n244 ) , .A1( us00_n245 ) , .A2( us00_n246 ) , .A3( us00_n247 ) , .A4( us00_n248 ) );
  NOR3_X1 us00_U7 (.A1( us00_n1 ) , .A3( us00_n100 ) , .A2( us00_n198 ) , .ZN( us00_n373 ) );
  NOR4_X1 us00_U70 (.A1( us00_n213 ) , .ZN( us00_n243 ) , .A2( us00_n249 ) , .A3( us00_n250 ) , .A4( us00_n251 ) );
  NAND4_X1 us00_U71 (.A1( us00_n217 ) , .A2( us00_n218 ) , .A3( us00_n219 ) , .A4( us00_n220 ) , .ZN( us00_n77 ) );
  NOR3_X1 us00_U72 (.ZN( us00_n218 ) , .A1( us00_n227 ) , .A2( us00_n228 ) , .A3( us00_n229 ) );
  NOR3_X1 us00_U73 (.ZN( us00_n219 ) , .A1( us00_n224 ) , .A2( us00_n225 ) , .A3( us00_n226 ) );
  NOR3_X1 us00_U74 (.ZN( us00_n220 ) , .A1( us00_n221 ) , .A2( us00_n222 ) , .A3( us00_n223 ) );
  NAND4_X1 us00_U75 (.ZN( us00_n270 ) , .A1( us00_n314 ) , .A2( us00_n315 ) , .A3( us00_n316 ) , .A4( us00_n317 ) );
  NOR4_X1 us00_U76 (.A2( us00_n109 ) , .A4( us00_n192 ) , .A3( us00_n216 ) , .A1( us00_n224 ) , .ZN( us00_n316 ) );
  NOR4_X1 us00_U77 (.ZN( us00_n315 ) , .A1( us00_n322 ) , .A2( us00_n323 ) , .A3( us00_n324 ) , .A4( us00_n325 ) );
  NOR4_X1 us00_U78 (.ZN( us00_n317 ) , .A1( us00_n318 ) , .A2( us00_n319 ) , .A3( us00_n320 ) , .A4( us00_n321 ) );
  NAND4_X1 us00_U79 (.A1( us00_n102 ) , .A2( us00_n103 ) , .A3( us00_n104 ) , .A4( us00_n105 ) , .ZN( us00_n76 ) );
  INV_X1 us00_U8 (.ZN( us00_n1 ) , .A( us00_n171 ) );
  NOR3_X1 us00_U80 (.ZN( us00_n104 ) , .A1( us00_n110 ) , .A2( us00_n111 ) , .A3( us00_n112 ) );
  NOR4_X1 us00_U81 (.ZN( us00_n105 ) , .A1( us00_n106 ) , .A2( us00_n107 ) , .A3( us00_n108 ) , .A4( us00_n109 ) );
  AOI222_X1 us00_U82 (.ZN( us00_n102 ) , .B1( us00_n16 ) , .A2( us00_n27 ) , .B2( us00_n36 ) , .C2( us00_n4 ) , .C1( us00_n43 ) , .A1( us00_n47 ) );
  NOR4_X1 us00_U83 (.ZN( us00_n201 ) , .A1( us00_n209 ) , .A2( us00_n210 ) , .A3( us00_n211 ) , .A4( us00_n212 ) );
  NOR4_X1 us00_U84 (.ZN( us00_n200 ) , .A1( us00_n213 ) , .A2( us00_n214 ) , .A3( us00_n215 ) , .A4( us00_n216 ) );
  NOR4_X1 us00_U85 (.A4( us00_n162 ) , .A2( us00_n18 ) , .ZN( us00_n202 ) , .A1( us00_n203 ) , .A3( us00_n204 ) );
  NOR2_X1 us00_U86 (.ZN( us00_n116 ) , .A2( us00_n43 ) , .A1( us00_n44 ) );
  AOI222_X1 us00_U87 (.A2( us00_n12 ) , .C1( us00_n14 ) , .ZN( us00_n233 ) , .B2( us00_n239 ) , .C2( us00_n31 ) , .A1( us00_n35 ) , .B1( us00_n36 ) );
  NOR4_X1 us00_U88 (.ZN( us00_n234 ) , .A1( us00_n235 ) , .A2( us00_n236 ) , .A3( us00_n237 ) , .A4( us00_n238 ) );
  NOR3_X1 us00_U89 (.A3( us00_n155 ) , .ZN( us00_n231 ) , .A1( us00_n269 ) , .A2( us00_n270 ) );
  NOR3_X1 us00_U9 (.A1( us00_n152 ) , .ZN( us00_n241 ) , .A2( us00_n255 ) , .A3( us00_n256 ) );
  AOI222_X1 us00_U90 (.A1( us00_n11 ) , .B1( us00_n14 ) , .C2( us00_n15 ) , .A2( us00_n34 ) , .ZN( us00_n364 ) , .B2( us00_n40 ) , .C1( us00_n45 ) );
  NOR4_X1 us00_U91 (.A3( us00_n207 ) , .ZN( us00_n365 ) , .A1( us00_n366 ) , .A2( us00_n367 ) , .A4( us00_n368 ) );
  INV_X1 us00_U92 (.A( us00_n372 ) , .ZN( us00_n6 ) );
  NAND4_X1 us00_U93 (.ZN( us00_n198 ) , .A1( us00_n418 ) , .A2( us00_n419 ) , .A3( us00_n420 ) , .A4( us00_n421 ) );
  NOR3_X1 us00_U94 (.A2( us00_n307 ) , .A1( us00_n322 ) , .A3( us00_n347 ) , .ZN( us00_n420 ) );
  AOI221_X1 us00_U95 (.C2( us00_n124 ) , .B2( us00_n16 ) , .C1( us00_n35 ) , .ZN( us00_n418 ) , .A( us00_n427 ) , .B1( us00_n45 ) );
  NOR4_X1 us00_U96 (.A3( us00_n166 ) , .A4( us00_n249 ) , .A1( us00_n278 ) , .A2( us00_n368 ) , .ZN( us00_n419 ) );
  NAND4_X1 us00_U97 (.ZN( us00_n255 ) , .A1( us00_n339 ) , .A2( us00_n340 ) , .A3( us00_n341 ) , .A4( us00_n342 ) );
  NOR4_X1 us00_U98 (.A3( us00_n176 ) , .ZN( us00_n339 ) , .A1( us00_n349 ) , .A2( us00_n350 ) , .A4( us00_n351 ) );
  NOR4_X1 us00_U99 (.A3( us00_n112 ) , .A4( us00_n209 ) , .A2( us00_n223 ) , .ZN( us00_n341 ) , .A1( us00_n346 ) );
  INV_X1 us03_U10 (.A( us03_n678 ) , .ZN( us03_n838 ) );
  NOR4_X1 us03_U100 (.A4( us03_n607 ) , .A3( us03_n608 ) , .A2( us03_n609 ) , .A1( us03_n610 ) , .ZN( us03_n617 ) );
  NOR4_X1 us03_U101 (.A4( us03_n612 ) , .A3( us03_n613 ) , .A2( us03_n614 ) , .A1( us03_n615 ) , .ZN( us03_n616 ) );
  NOR2_X1 us03_U102 (.ZN( us03_n684 ) , .A1( us03_n829 ) , .A2( us03_n830 ) );
  NAND4_X1 us03_U103 (.A4( us03_n471 ) , .A3( us03_n472 ) , .A2( us03_n473 ) , .A1( us03_n474 ) , .ZN( us03_n676 ) );
  NOR4_X1 us03_U104 (.A4( us03_n468 ) , .ZN( us03_n474 ) , .A3( us03_n554 ) , .A1( us03_n733 ) , .A2( us03_n753 ) );
  NOR4_X1 us03_U105 (.ZN( us03_n473 ) , .A1( us03_n529 ) , .A3( us03_n566 ) , .A4( us03_n598 ) , .A2( us03_n640 ) );
  NOR4_X1 us03_U106 (.ZN( us03_n472 ) , .A1( us03_n504 ) , .A3( us03_n542 ) , .A2( us03_n581 ) , .A4( us03_n714 ) );
  NAND4_X1 us03_U107 (.ZN( sa03_sr_1 ) , .A4( us03_n593 ) , .A3( us03_n594 ) , .A2( us03_n595 ) , .A1( us03_n596 ) );
  AOI211_X1 us03_U108 (.B( us03_n587 ) , .A( us03_n588 ) , .ZN( us03_n594 ) , .C2( us03_n809 ) , .C1( us03_n831 ) );
  NOR4_X1 us03_U109 (.A4( us03_n589 ) , .A3( us03_n590 ) , .A2( us03_n591 ) , .A1( us03_n592 ) , .ZN( us03_n593 ) );
  NOR4_X1 us03_U11 (.A4( us03_n443 ) , .A3( us03_n444 ) , .A2( us03_n514 ) , .A1( us03_n539 ) , .ZN( us03_n704 ) );
  AOI211_X1 us03_U110 (.A( us03_n586 ) , .ZN( us03_n595 ) , .B( us03_n619 ) , .C1( us03_n843 ) , .C2( us03_n853 ) );
  NAND4_X1 us03_U111 (.ZN( sa03_sr_0 ) , .A4( us03_n499 ) , .A3( us03_n500 ) , .A2( us03_n501 ) , .A1( us03_n502 ) );
  NOR4_X1 us03_U112 (.A4( us03_n496 ) , .A3( us03_n497 ) , .A2( us03_n498 ) , .ZN( us03_n499 ) , .A1( us03_n525 ) );
  AOI221_X1 us03_U113 (.A( us03_n495 ) , .ZN( us03_n500 ) , .B2( us03_n841 ) , .C1( us03_n844 ) , .C2( us03_n858 ) , .B1( us03_n860 ) );
  AOI211_X1 us03_U114 (.A( us03_n494 ) , .ZN( us03_n501 ) , .B( us03_n800 ) , .C2( us03_n837 ) , .C1( us03_n849 ) );
  NAND4_X1 us03_U115 (.A4( us03_n689 ) , .A3( us03_n690 ) , .A1( us03_n691 ) , .ZN( us03_n774 ) , .A2( us03_n870 ) );
  INV_X1 us03_U116 (.A( us03_n677 ) , .ZN( us03_n870 ) );
  AOI221_X1 us03_U117 (.A( us03_n679 ) , .ZN( us03_n690 ) , .B2( us03_n838 ) , .C1( us03_n840 ) , .C2( us03_n860 ) , .B1( us03_n863 ) );
  NOR4_X1 us03_U118 (.A4( us03_n685 ) , .A3( us03_n686 ) , .A2( us03_n687 ) , .A1( us03_n688 ) , .ZN( us03_n689 ) );
  NOR2_X1 us03_U119 (.ZN( us03_n731 ) , .A2( us03_n830 ) , .A1( us03_n843 ) );
  OR3_X1 us03_U12 (.ZN( us03_n444 ) , .A1( us03_n526 ) , .A3( us03_n575 ) , .A2( us03_n873 ) );
  NAND4_X1 us03_U120 (.A4( us03_n717 ) , .A3( us03_n718 ) , .A2( us03_n719 ) , .ZN( us03_n739 ) , .A1( us03_n855 ) );
  INV_X1 us03_U121 (.A( us03_n707 ) , .ZN( us03_n855 ) );
  NOR4_X1 us03_U122 (.A4( us03_n713 ) , .A3( us03_n714 ) , .A2( us03_n715 ) , .A1( us03_n716 ) , .ZN( us03_n717 ) );
  AOI221_X1 us03_U123 (.A( us03_n708 ) , .ZN( us03_n719 ) , .C2( us03_n842 ) , .B2( us03_n843 ) , .C1( us03_n859 ) , .B1( us03_n860 ) );
  NOR2_X1 us03_U124 (.ZN( us03_n645 ) , .A1( us03_n852 ) , .A2( us03_n866 ) );
  NAND4_X1 us03_U125 (.A4( us03_n571 ) , .A3( us03_n572 ) , .A1( us03_n573 ) , .ZN( us03_n721 ) , .A2( us03_n872 ) );
  NOR4_X1 us03_U126 (.A4( us03_n567 ) , .A3( us03_n568 ) , .A2( us03_n569 ) , .A1( us03_n570 ) , .ZN( us03_n571 ) );
  AOI221_X1 us03_U127 (.A( us03_n562 ) , .C2( us03_n563 ) , .ZN( us03_n572 ) , .B2( us03_n843 ) , .B1( us03_n850 ) , .C1( us03_n851 ) );
  INV_X1 us03_U128 (.A( us03_n605 ) , .ZN( us03_n872 ) );
  NAND4_X1 us03_U129 (.A4( us03_n491 ) , .A3( us03_n492 ) , .A1( us03_n493 ) , .ZN( us03_n800 ) , .A2( us03_n865 ) );
  OR4_X1 us03_U13 (.A4( us03_n440 ) , .A2( us03_n441 ) , .A1( us03_n442 ) , .ZN( us03_n443 ) , .A3( us03_n551 ) );
  AOI221_X1 us03_U130 (.A( us03_n487 ) , .ZN( us03_n492 ) , .B2( us03_n834 ) , .C2( us03_n839 ) , .C1( us03_n849 ) , .B1( us03_n858 ) );
  INV_X1 us03_U131 (.A( us03_n776 ) , .ZN( us03_n865 ) );
  NOR2_X1 us03_U132 (.ZN( us03_n493 ) , .A1( us03_n676 ) , .A2( us03_n692 ) );
  INV_X1 us03_U133 (.A( us03_n760 ) , .ZN( us03_n828 ) );
  INV_X1 us03_U134 (.A( us03_n461 ) , .ZN( us03_n862 ) );
  OAI21_X1 us03_U135 (.ZN( us03_n461 ) , .B1( us03_n807 ) , .A( us03_n832 ) , .B2( us03_n849 ) );
  OR4_X1 us03_U136 (.A4( us03_n578 ) , .A3( us03_n579 ) , .A2( us03_n580 ) , .A1( us03_n581 ) , .ZN( us03_n582 ) );
  OR4_X1 us03_U137 (.A4( us03_n564 ) , .A3( us03_n565 ) , .A2( us03_n566 ) , .ZN( us03_n570 ) , .A1( us03_n663 ) );
  OR4_X1 us03_U138 (.A4( us03_n516 ) , .A2( us03_n517 ) , .A1( us03_n518 ) , .ZN( us03_n520 ) , .A3( us03_n819 ) );
  OR4_X1 us03_U139 (.A4( us03_n680 ) , .A3( us03_n681 ) , .A2( us03_n682 ) , .A1( us03_n683 ) , .ZN( us03_n688 ) );
  INV_X1 us03_U14 (.A( us03_n611 ) , .ZN( us03_n873 ) );
  OR4_X1 us03_U140 (.ZN( us03_n464 ) , .A4( us03_n516 ) , .A3( us03_n527 ) , .A2( us03_n576 ) , .A1( us03_n710 ) );
  NAND2_X1 us03_U141 (.ZN( us03_n611 ) , .A2( us03_n835 ) , .A1( us03_n871 ) );
  OR3_X1 us03_U142 (.A3( us03_n504 ) , .A2( us03_n505 ) , .A1( us03_n506 ) , .ZN( us03_n509 ) );
  AOI221_X1 us03_U143 (.A( us03_n711 ) , .B2( us03_n712 ) , .ZN( us03_n718 ) , .C1( us03_n830 ) , .B1( us03_n837 ) , .C2( us03_n861 ) );
  OR2_X1 us03_U144 (.A2( us03_n709 ) , .A1( us03_n710 ) , .ZN( us03_n711 ) );
  INV_X1 us03_U145 (.A( us03_n752 ) , .ZN( us03_n867 ) );
  OAI21_X1 us03_U146 (.B1( us03_n751 ) , .ZN( us03_n752 ) , .A( us03_n843 ) , .B2( us03_n866 ) );
  INV_X1 us03_U147 (.A( us03_n670 ) , .ZN( us03_n857 ) );
  AOI21_X1 us03_U148 (.A( us03_n668 ) , .B1( us03_n669 ) , .ZN( us03_n670 ) , .B2( us03_n854 ) );
  AOI222_X1 us03_U149 (.ZN( us03_n658 ) , .A2( us03_n837 ) , .B1( us03_n839 ) , .C2( us03_n843 ) , .A1( us03_n858 ) , .C1( us03_n861 ) , .B2( us03_n868 ) );
  INV_X1 us03_U15 (.A( us03_n747 ) , .ZN( us03_n861 ) );
  INV_X1 us03_U150 (.A( us03_n645 ) , .ZN( us03_n868 ) );
  OAI22_X1 us03_U151 (.ZN( us03_n481 ) , .A1( us03_n706 ) , .B2( us03_n783 ) , .A2( us03_n804 ) , .B1( us03_n810 ) );
  NAND2_X1 us03_U152 (.A1( us03_n445 ) , .A2( us03_n463 ) , .ZN( us03_n747 ) );
  OAI222_X1 us03_U153 (.B2( us03_n745 ) , .B1( us03_n746 ) , .A2( us03_n747 ) , .ZN( us03_n755 ) , .C2( us03_n803 ) , .C1( us03_n812 ) , .A1( us03_n815 ) );
  OAI222_X1 us03_U154 (.B2( us03_n706 ) , .ZN( us03_n707 ) , .C2( us03_n722 ) , .B1( us03_n745 ) , .A1( us03_n804 ) , .C1( us03_n812 ) , .A2( us03_n813 ) );
  OAI222_X1 us03_U155 (.ZN( us03_n615 ) , .B1( us03_n695 ) , .C1( us03_n722 ) , .C2( us03_n745 ) , .B2( us03_n784 ) , .A2( us03_n790 ) , .A1( us03_n814 ) );
  OAI222_X1 us03_U156 (.ZN( us03_n503 ) , .C2( us03_n623 ) , .B2( us03_n645 ) , .B1( us03_n745 ) , .A2( us03_n746 ) , .C1( us03_n803 ) , .A1( us03_n804 ) );
  AOI22_X1 us03_U157 (.ZN( us03_n694 ) , .A1( us03_n828 ) , .B2( us03_n841 ) , .A2( us03_n863 ) , .B1( us03_n866 ) );
  INV_X1 us03_U158 (.A( us03_n728 ) , .ZN( us03_n837 ) );
  AOI221_X1 us03_U159 (.A( us03_n762 ) , .ZN( us03_n772 ) , .C2( us03_n808 ) , .B2( us03_n833 ) , .C1( us03_n853 ) , .B1( us03_n864 ) );
  AOI222_X1 us03_U16 (.ZN( us03_n561 ) , .B1( us03_n828 ) , .C1( us03_n839 ) , .A2( us03_n841 ) , .A1( us03_n852 ) , .B2( us03_n861 ) , .C2( us03_n871 ) );
  AOI21_X1 us03_U160 (.B2( us03_n761 ) , .ZN( us03_n762 ) , .A( us03_n786 ) , .B1( us03_n790 ) );
  INV_X1 us03_U161 (.A( us03_n759 ) , .ZN( us03_n833 ) );
  NAND2_X1 us03_U162 (.A1( us03_n449 ) , .A2( us03_n451 ) , .ZN( us03_n760 ) );
  INV_X1 us03_U163 (.A( us03_n788 ) , .ZN( us03_n830 ) );
  OAI22_X1 us03_U164 (.ZN( us03_n635 ) , .A1( us03_n697 ) , .B2( us03_n726 ) , .A2( us03_n760 ) , .B1( us03_n814 ) );
  OAI221_X1 us03_U165 (.A( us03_n725 ) , .C2( us03_n726 ) , .B2( us03_n727 ) , .B1( us03_n728 ) , .ZN( us03_n735 ) , .C1( us03_n815 ) );
  AOI22_X1 us03_U166 (.ZN( us03_n725 ) , .B1( us03_n830 ) , .A2( us03_n836 ) , .A1( us03_n861 ) , .B2( us03_n864 ) );
  OAI22_X1 us03_U167 (.ZN( us03_n487 ) , .A1( us03_n722 ) , .B2( us03_n726 ) , .B1( us03_n728 ) , .A2( us03_n777 ) );
  OAI22_X1 us03_U168 (.ZN( us03_n622 ) , .B1( us03_n667 ) , .B2( us03_n745 ) , .A1( us03_n813 ) , .A2( us03_n814 ) );
  OAI22_X1 us03_U169 (.A1( us03_n722 ) , .ZN( us03_n724 ) , .B2( us03_n748 ) , .B1( us03_n810 ) , .A2( us03_n814 ) );
  NOR4_X1 us03_U17 (.ZN( us03_n471 ) , .A2( us03_n519 ) , .A4( us03_n592 ) , .A1( us03_n607 ) , .A3( us03_n627 ) );
  OAI22_X1 us03_U170 (.B2( us03_n777 ) , .B1( us03_n778 ) , .ZN( us03_n779 ) , .A2( us03_n812 ) , .A1( us03_n813 ) );
  OAI22_X1 us03_U171 (.B2( us03_n742 ) , .ZN( us03_n744 ) , .A2( us03_n760 ) , .B1( us03_n778 ) , .A1( us03_n790 ) );
  OAI22_X1 us03_U172 (.B2( us03_n801 ) , .B1( us03_n802 ) , .A2( us03_n803 ) , .A1( us03_n804 ) , .ZN( us03_n806 ) );
  OAI22_X1 us03_U173 (.ZN( us03_n494 ) , .A2( us03_n742 ) , .A1( us03_n778 ) , .B1( us03_n789 ) , .B2( us03_n804 ) );
  INV_X1 us03_U174 (.A( us03_n742 ) , .ZN( us03_n835 ) );
  INV_X1 us03_U175 (.A( us03_n814 ) , .ZN( us03_n829 ) );
  INV_X1 us03_U176 (.A( us03_n786 ) , .ZN( us03_n843 ) );
  INV_X1 us03_U177 (.A( us03_n812 ) , .ZN( us03_n831 ) );
  OAI22_X1 us03_U178 (.ZN( us03_n588 ) , .B1( us03_n728 ) , .B2( us03_n747 ) , .A2( us03_n784 ) , .A1( us03_n801 ) );
  OAI22_X1 us03_U179 (.ZN( us03_n693 ) , .A2( us03_n728 ) , .A1( us03_n778 ) , .B1( us03_n789 ) , .B2( us03_n815 ) );
  NOR4_X1 us03_U18 (.ZN( us03_n477 ) , .A1( us03_n518 ) , .A4( us03_n555 ) , .A3( us03_n580 ) , .A2( us03_n628 ) );
  OAI22_X1 us03_U180 (.ZN( us03_n708 ) , .A2( us03_n726 ) , .B2( us03_n727 ) , .A1( us03_n742 ) , .B1( us03_n811 ) );
  INV_X1 us03_U181 (.A( us03_n667 ) , .ZN( us03_n863 ) );
  NOR2_X1 us03_U182 (.A1( us03_n695 ) , .ZN( us03_n768 ) , .A2( us03_n813 ) );
  NOR2_X1 us03_U183 (.ZN( us03_n664 ) , .A1( us03_n726 ) , .A2( us03_n801 ) );
  NOR2_X1 us03_U184 (.ZN( us03_n592 ) , .A2( us03_n695 ) , .A1( us03_n726 ) );
  NOR2_X1 us03_U185 (.ZN( us03_n568 ) , .A1( us03_n726 ) , .A2( us03_n804 ) );
  NOR2_X1 us03_U186 (.ZN( us03_n716 ) , .A2( us03_n722 ) , .A1( us03_n742 ) );
  NOR2_X1 us03_U187 (.ZN( us03_n544 ) , .A2( us03_n778 ) , .A1( us03_n812 ) );
  NOR2_X1 us03_U188 (.ZN( us03_n575 ) , .A2( us03_n697 ) , .A1( us03_n812 ) );
  NOR2_X1 us03_U189 (.ZN( us03_n652 ) , .A1( us03_n726 ) , .A2( us03_n811 ) );
  NOR4_X1 us03_U19 (.A4( us03_n530 ) , .A3( us03_n531 ) , .A2( us03_n532 ) , .ZN( us03_n533 ) , .A1( us03_n818 ) );
  NOR2_X1 us03_U190 (.ZN( us03_n610 ) , .A1( us03_n777 ) , .A2( us03_n784 ) );
  INV_X1 us03_U191 (.A( us03_n748 ) , .ZN( us03_n840 ) );
  NOR2_X1 us03_U192 (.ZN( us03_n530 ) , .A2( us03_n747 ) , .A1( us03_n748 ) );
  NOR2_X1 us03_U193 (.ZN( us03_n627 ) , .A2( us03_n726 ) , .A1( us03_n783 ) );
  NOR2_X1 us03_U194 (.ZN( us03_n613 ) , .A1( us03_n783 ) , .A2( us03_n813 ) );
  NOR2_X1 us03_U195 (.ZN( us03_n599 ) , .A2( us03_n778 ) , .A1( us03_n801 ) );
  NOR2_X1 us03_U196 (.ZN( us03_n609 ) , .A2( us03_n778 ) , .A1( us03_n804 ) );
  INV_X1 us03_U197 (.A( us03_n745 ) , .ZN( us03_n832 ) );
  NOR2_X1 us03_U198 (.A2( us03_n742 ) , .ZN( us03_n767 ) , .A1( us03_n810 ) );
  NOR2_X1 us03_U199 (.ZN( us03_n526 ) , .A2( us03_n722 ) , .A1( us03_n801 ) );
  NOR4_X1 us03_U20 (.ZN( us03_n454 ) , .A2( us03_n515 ) , .A1( us03_n541 ) , .A3( us03_n577 ) , .A4( us03_n613 ) );
  NOR2_X1 us03_U200 (.ZN( us03_n529 ) , .A2( us03_n778 ) , .A1( us03_n814 ) );
  NOR2_X1 us03_U201 (.ZN( us03_n626 ) , .A2( us03_n667 ) , .A1( us03_n783 ) );
  NOR2_X1 us03_U202 (.ZN( us03_n597 ) , .A2( us03_n789 ) , .A1( us03_n814 ) );
  INV_X1 us03_U203 (.A( us03_n790 ) , .ZN( us03_n849 ) );
  NOR2_X1 us03_U204 (.ZN( us03_n650 ) , .A1( us03_n667 ) , .A2( us03_n812 ) );
  NOR2_X1 us03_U205 (.A1( us03_n667 ) , .ZN( us03_n671 ) , .A2( us03_n742 ) );
  NOR2_X1 us03_U206 (.ZN( us03_n600 ) , .A1( us03_n667 ) , .A2( us03_n801 ) );
  NOR2_X1 us03_U207 (.A1( us03_n667 ) , .ZN( us03_n686 ) , .A2( us03_n814 ) );
  NOR2_X1 us03_U208 (.A2( us03_n706 ) , .A1( us03_n748 ) , .ZN( us03_n769 ) );
  NOR2_X1 us03_U209 (.A1( us03_n667 ) , .ZN( us03_n764 ) , .A2( us03_n811 ) );
  NOR4_X1 us03_U21 (.A4( us03_n539 ) , .A3( us03_n540 ) , .A2( us03_n541 ) , .ZN( us03_n548 ) , .A1( us03_n686 ) );
  NOR2_X1 us03_U210 (.A1( us03_n697 ) , .ZN( us03_n766 ) , .A2( us03_n811 ) );
  NOR2_X1 us03_U211 (.ZN( us03_n539 ) , .A2( us03_n695 ) , .A1( us03_n697 ) );
  NOR2_X1 us03_U212 (.ZN( us03_n525 ) , .A1( us03_n667 ) , .A2( us03_n777 ) );
  NOR2_X1 us03_U213 (.ZN( us03_n665 ) , .A1( us03_n748 ) , .A2( us03_n813 ) );
  NOR2_X1 us03_U214 (.ZN( us03_n553 ) , .A1( us03_n748 ) , .A2( us03_n789 ) );
  NOR2_X1 us03_U215 (.ZN( us03_n506 ) , .A2( us03_n778 ) , .A1( us03_n783 ) );
  NOR2_X1 us03_U216 (.ZN( us03_n541 ) , .A2( us03_n706 ) , .A1( us03_n783 ) );
  NOR2_X1 us03_U217 (.ZN( us03_n662 ) , .A1( us03_n783 ) , .A2( us03_n789 ) );
  NOR2_X1 us03_U218 (.A2( us03_n695 ) , .ZN( us03_n714 ) , .A1( us03_n790 ) );
  OAI22_X1 us03_U219 (.B1( us03_n438 ) , .ZN( us03_n442 ) , .A2( us03_n726 ) , .A1( us03_n742 ) , .B2( us03_n747 ) );
  NOR2_X1 us03_U22 (.ZN( us03_n678 ) , .A2( us03_n832 ) , .A1( us03_n837 ) );
  NOR3_X1 us03_U220 (.ZN( us03_n438 ) , .A2( us03_n834 ) , .A3( us03_n835 ) , .A1( us03_n844 ) );
  NOR2_X1 us03_U221 (.ZN( us03_n505 ) , .A1( us03_n810 ) , .A2( us03_n815 ) );
  INV_X1 us03_U222 (.A( us03_n804 ) , .ZN( us03_n839 ) );
  NOR2_X1 us03_U223 (.ZN( us03_n659 ) , .A1( us03_n727 ) , .A2( us03_n788 ) );
  NOR2_X1 us03_U224 (.ZN( us03_n660 ) , .A2( us03_n695 ) , .A1( us03_n727 ) );
  NOR2_X1 us03_U225 (.ZN( us03_n555 ) , .A1( us03_n790 ) , .A2( us03_n812 ) );
  NOR2_X1 us03_U226 (.ZN( us03_n543 ) , .A1( us03_n747 ) , .A2( us03_n812 ) );
  NOR2_X1 us03_U227 (.ZN( us03_n507 ) , .A1( us03_n727 ) , .A2( us03_n777 ) );
  INV_X1 us03_U228 (.A( us03_n801 ) , .ZN( us03_n841 ) );
  NOR2_X1 us03_U229 (.A2( us03_n695 ) , .A1( us03_n778 ) , .ZN( us03_n818 ) );
  NOR4_X1 us03_U23 (.A4( us03_n512 ) , .A3( us03_n513 ) , .A2( us03_n514 ) , .A1( us03_n515 ) , .ZN( us03_n522 ) );
  NOR2_X1 us03_U230 (.ZN( us03_n528 ) , .A2( us03_n742 ) , .A1( us03_n790 ) );
  OAI22_X1 us03_U231 (.B2( us03_n748 ) , .B1( us03_n749 ) , .A1( us03_n750 ) , .ZN( us03_n754 ) , .A2( us03_n804 ) );
  NOR2_X1 us03_U232 (.ZN( us03_n749 ) , .A2( us03_n850 ) , .A1( us03_n858 ) );
  NOR3_X1 us03_U233 (.ZN( us03_n750 ) , .A2( us03_n851 ) , .A1( us03_n861 ) , .A3( us03_n863 ) );
  NOR2_X1 us03_U234 (.A1( us03_n747 ) , .ZN( us03_n765 ) , .A2( us03_n801 ) );
  NOR2_X1 us03_U235 (.A2( us03_n742 ) , .ZN( us03_n753 ) , .A1( us03_n803 ) );
  NOR2_X1 us03_U236 (.ZN( us03_n542 ) , .A2( us03_n783 ) , .A1( us03_n790 ) );
  NOR2_X1 us03_U237 (.ZN( us03_n661 ) , .A1( us03_n727 ) , .A2( us03_n783 ) );
  INV_X1 us03_U238 (.A( us03_n726 ) , .ZN( us03_n850 ) );
  NOR2_X1 us03_U239 (.ZN( us03_n629 ) , .A1( us03_n722 ) , .A2( us03_n811 ) );
  AOI222_X1 us03_U24 (.ZN( us03_n523 ) , .A1( us03_n832 ) , .B2( us03_n835 ) , .C1( us03_n842 ) , .C2( us03_n848 ) , .A2( us03_n850 ) , .B1( us03_n864 ) );
  NOR2_X1 us03_U240 (.ZN( us03_n733 ) , .A2( us03_n801 ) , .A1( us03_n803 ) );
  NOR2_X1 us03_U241 (.ZN( us03_n612 ) , .A1( us03_n760 ) , .A2( us03_n810 ) );
  NOR4_X1 us03_U242 (.A2( us03_n489 ) , .A1( us03_n490 ) , .ZN( us03_n491 ) , .A3( us03_n578 ) , .A4( us03_n610 ) );
  OR4_X1 us03_U243 (.ZN( us03_n490 ) , .A4( us03_n532 ) , .A2( us03_n545 ) , .A1( us03_n557 ) , .A3( us03_n630 ) );
  OAI22_X1 us03_U244 (.B1( us03_n488 ) , .ZN( us03_n489 ) , .A1( us03_n684 ) , .A2( us03_n761 ) , .B2( us03_n815 ) );
  NOR3_X1 us03_U245 (.ZN( us03_n488 ) , .A1( us03_n780 ) , .A2( us03_n848 ) , .A3( us03_n861 ) );
  NOR2_X1 us03_U246 (.ZN( us03_n504 ) , .A2( us03_n726 ) , .A1( us03_n760 ) );
  NOR2_X1 us03_U247 (.ZN( us03_n514 ) , .A1( us03_n706 ) , .A2( us03_n742 ) );
  NOR2_X1 us03_U248 (.ZN( us03_n715 ) , .A2( us03_n742 ) , .A1( us03_n784 ) );
  NOR2_X1 us03_U249 (.ZN( us03_n552 ) , .A1( us03_n784 ) , .A2( us03_n811 ) );
  NOR4_X1 us03_U25 (.A3( us03_n519 ) , .A1( us03_n520 ) , .ZN( us03_n521 ) , .A2( us03_n671 ) , .A4( us03_n767 ) );
  NOR2_X1 us03_U250 (.ZN( us03_n515 ) , .A1( us03_n706 ) , .A2( us03_n801 ) );
  NOR2_X1 us03_U251 (.ZN( us03_n556 ) , .A1( us03_n706 ) , .A2( us03_n814 ) );
  NOR2_X1 us03_U252 (.ZN( us03_n519 ) , .A1( us03_n788 ) , .A2( us03_n810 ) );
  INV_X1 us03_U253 (.A( us03_n803 ) , .ZN( us03_n858 ) );
  NOR2_X1 us03_U254 (.ZN( us03_n628 ) , .A1( us03_n745 ) , .A2( us03_n813 ) );
  NOR2_X1 us03_U255 (.ZN( us03_n713 ) , .A1( us03_n803 ) , .A2( us03_n815 ) );
  AOI21_X1 us03_U256 (.ZN( us03_n569 ) , .B2( us03_n695 ) , .B1( us03_n804 ) , .A( us03_n810 ) );
  NOR2_X1 us03_U257 (.ZN( us03_n653 ) , .A1( us03_n788 ) , .A2( us03_n813 ) );
  NOR2_X1 us03_U258 (.ZN( us03_n666 ) , .A2( us03_n706 ) , .A1( us03_n788 ) );
  NOR2_X1 us03_U259 (.ZN( us03_n654 ) , .A1( us03_n745 ) , .A2( us03_n778 ) );
  AOI222_X1 us03_U26 (.B2( us03_n636 ) , .ZN( us03_n642 ) , .B1( us03_n839 ) , .A1( us03_n840 ) , .C2( us03_n844 ) , .C1( us03_n861 ) , .A2( us03_n863 ) );
  NOR2_X1 us03_U260 (.ZN( us03_n554 ) , .A1( us03_n760 ) , .A2( us03_n803 ) );
  NOR2_X1 us03_U261 (.ZN( us03_n540 ) , .A1( us03_n760 ) , .A2( us03_n789 ) );
  NOR2_X1 us03_U262 (.ZN( us03_n699 ) , .A2( us03_n784 ) , .A1( us03_n815 ) );
  NOR2_X1 us03_U263 (.ZN( us03_n607 ) , .A2( us03_n722 ) , .A1( us03_n815 ) );
  NOR2_X1 us03_U264 (.A1( us03_n728 ) , .ZN( us03_n763 ) , .A2( us03_n784 ) );
  AOI21_X1 us03_U265 (.A( us03_n813 ) , .B2( us03_n814 ) , .B1( us03_n815 ) , .ZN( us03_n816 ) );
  NOR2_X1 us03_U266 (.ZN( us03_n577 ) , .A2( us03_n706 ) , .A1( us03_n728 ) );
  NOR2_X1 us03_U267 (.ZN( us03_n531 ) , .A2( us03_n722 ) , .A1( us03_n728 ) );
  AOI21_X1 us03_U268 (.B1( us03_n623 ) , .ZN( us03_n625 ) , .A( us03_n761 ) , .B2( us03_n812 ) );
  AOI21_X1 us03_U269 (.A( us03_n810 ) , .B2( us03_n811 ) , .B1( us03_n812 ) , .ZN( us03_n817 ) );
  NOR4_X1 us03_U27 (.A4( us03_n637 ) , .A3( us03_n638 ) , .A2( us03_n639 ) , .A1( us03_n640 ) , .ZN( us03_n641 ) );
  AOI21_X1 us03_U270 (.ZN( us03_n513 ) , .A( us03_n727 ) , .B1( us03_n748 ) , .B2( us03_n801 ) );
  AOI21_X1 us03_U271 (.ZN( us03_n497 ) , .B1( us03_n678 ) , .A( us03_n810 ) , .B2( us03_n814 ) );
  AOI21_X1 us03_U272 (.ZN( us03_n476 ) , .B2( us03_n695 ) , .A( us03_n747 ) , .B1( us03_n777 ) );
  NOR2_X1 us03_U273 (.ZN( us03_n580 ) , .A1( us03_n742 ) , .A2( us03_n813 ) );
  NOR2_X1 us03_U274 (.ZN( us03_n640 ) , .A2( us03_n786 ) , .A1( us03_n789 ) );
  AOI21_X1 us03_U275 (.ZN( us03_n591 ) , .B1( us03_n748 ) , .A( us03_n790 ) , .B2( us03_n811 ) );
  NOR2_X1 us03_U276 (.A2( us03_n706 ) , .A1( us03_n760 ) , .ZN( us03_n792 ) );
  AOI21_X1 us03_U277 (.ZN( us03_n624 ) , .B2( us03_n667 ) , .A( us03_n788 ) , .B1( us03_n789 ) );
  NOR2_X1 us03_U278 (.ZN( us03_n668 ) , .A1( us03_n788 ) , .A2( us03_n803 ) );
  NOR2_X1 us03_U279 (.ZN( us03_n518 ) , .A2( us03_n706 ) , .A1( us03_n812 ) );
  NOR3_X1 us03_U28 (.A2( us03_n605 ) , .A1( us03_n606 ) , .ZN( us03_n644 ) , .A3( us03_n720 ) );
  AOI21_X1 us03_U280 (.ZN( us03_n475 ) , .A( us03_n667 ) , .B1( us03_n748 ) , .B2( us03_n804 ) );
  NOR2_X1 us03_U281 (.ZN( us03_n557 ) , .A2( us03_n789 ) , .A1( us03_n801 ) );
  NOR2_X1 us03_U282 (.ZN( us03_n517 ) , .A2( us03_n697 ) , .A1( us03_n814 ) );
  NOR2_X1 us03_U283 (.ZN( us03_n681 ) , .A2( us03_n697 ) , .A1( us03_n801 ) );
  NOR2_X1 us03_U284 (.ZN( us03_n651 ) , .A1( us03_n760 ) , .A2( us03_n784 ) );
  INV_X1 us03_U285 (.A( us03_n811 ) , .ZN( us03_n834 ) );
  AOI21_X1 us03_U286 (.ZN( us03_n508 ) , .B2( us03_n667 ) , .A( us03_n728 ) , .B1( us03_n813 ) );
  AOI21_X1 us03_U287 (.ZN( us03_n537 ) , .B2( us03_n810 ) , .A( us03_n812 ) , .B1( us03_n813 ) );
  INV_X1 us03_U288 (.A( us03_n761 ) , .ZN( us03_n864 ) );
  AOI21_X1 us03_U289 (.ZN( us03_n538 ) , .A( us03_n761 ) , .B2( us03_n777 ) , .B1( us03_n815 ) );
  AOI221_X1 us03_U29 (.A( us03_n779 ) , .ZN( us03_n796 ) , .C2( us03_n835 ) , .B2( us03_n836 ) , .B1( us03_n863 ) , .C1( us03_n864 ) );
  NOR2_X1 us03_U290 (.ZN( us03_n579 ) , .A1( us03_n667 ) , .A2( us03_n786 ) );
  AOI21_X1 us03_U291 (.ZN( us03_n587 ) , .B2( us03_n697 ) , .B1( us03_n813 ) , .A( us03_n815 ) );
  AOI21_X1 us03_U292 (.B1( us03_n697 ) , .ZN( us03_n698 ) , .A( us03_n730 ) , .B2( us03_n761 ) );
  AOI21_X1 us03_U293 (.ZN( us03_n589 ) , .B2( us03_n761 ) , .A( us03_n783 ) , .B1( us03_n810 ) );
  AOI21_X1 us03_U294 (.ZN( us03_n496 ) , .A( us03_n722 ) , .B2( us03_n760 ) , .B1( us03_n812 ) );
  AOI21_X1 us03_U295 (.ZN( us03_n550 ) , .B1( us03_n667 ) , .A( us03_n695 ) , .B2( us03_n803 ) );
  NOR2_X1 us03_U296 (.ZN( us03_n545 ) , .A1( us03_n697 ) , .A2( us03_n742 ) );
  INV_X1 us03_U297 (.A( us03_n727 ) , .ZN( us03_n866 ) );
  INV_X1 us03_U298 (.A( us03_n789 ) , .ZN( us03_n871 ) );
  INV_X1 us03_U299 (.A( us03_n810 ) , .ZN( us03_n852 ) );
  NOR3_X1 us03_U3 (.ZN( us03_n596 ) , .A1( us03_n606 ) , .A3( us03_n721 ) , .A2( us03_n740 ) );
  NOR4_X1 us03_U30 (.A4( us03_n791 ) , .A3( us03_n792 ) , .A2( us03_n793 ) , .A1( us03_n794 ) , .ZN( us03_n795 ) );
  AOI21_X1 us03_U300 (.ZN( us03_n638 ) , .B2( us03_n745 ) , .A( us03_n790 ) , .B1( us03_n801 ) );
  AOI21_X1 us03_U301 (.ZN( us03_n647 ) , .B1( us03_n727 ) , .B2( us03_n761 ) , .A( us03_n811 ) );
  INV_X1 us03_U302 (.A( us03_n784 ) , .ZN( us03_n860 ) );
  NOR2_X1 us03_U303 (.ZN( us03_n683 ) , .A1( us03_n727 ) , .A2( us03_n814 ) );
  AOI21_X1 us03_U304 (.B1( us03_n684 ) , .ZN( us03_n685 ) , .A( us03_n726 ) , .B2( us03_n759 ) );
  AOI21_X1 us03_U305 (.ZN( us03_n567 ) , .B1( us03_n748 ) , .B2( us03_n760 ) , .A( us03_n778 ) );
  AOI21_X1 us03_U306 (.ZN( us03_n498 ) , .A( us03_n695 ) , .B1( us03_n706 ) , .B2( us03_n784 ) );
  NOR2_X1 us03_U307 (.ZN( us03_n566 ) , .A1( us03_n727 ) , .A2( us03_n760 ) );
  AOI21_X1 us03_U308 (.ZN( us03_n637 ) , .B2( us03_n747 ) , .A( us03_n786 ) , .B1( us03_n810 ) );
  NOR2_X1 us03_U309 (.ZN( us03_n564 ) , .A2( us03_n695 ) , .A1( us03_n761 ) );
  NOR4_X1 us03_U31 (.A4( us03_n774 ) , .A3( us03_n775 ) , .A1( us03_n776 ) , .ZN( us03_n797 ) , .A2( us03_n799 ) );
  NOR2_X1 us03_U310 (.ZN( us03_n578 ) , .A2( us03_n695 ) , .A1( us03_n789 ) );
  AOI21_X1 us03_U311 (.ZN( us03_n512 ) , .A( us03_n777 ) , .B2( us03_n790 ) , .B1( us03_n810 ) );
  INV_X1 us03_U312 (.A( us03_n697 ) , .ZN( us03_n851 ) );
  NOR2_X1 us03_U313 (.ZN( us03_n663 ) , .A1( us03_n778 ) , .A2( us03_n811 ) );
  AOI21_X1 us03_U314 (.ZN( us03_n448 ) , .B2( us03_n790 ) , .A( us03_n801 ) , .B1( us03_n813 ) );
  NOR2_X1 us03_U315 (.ZN( us03_n630 ) , .A2( us03_n695 ) , .A1( us03_n722 ) );
  AOI21_X1 us03_U316 (.ZN( us03_n562 ) , .B1( us03_n722 ) , .A( us03_n777 ) , .B2( us03_n789 ) );
  AOI21_X1 us03_U317 (.ZN( us03_n687 ) , .B2( us03_n747 ) , .B1( us03_n761 ) , .A( us03_n804 ) );
  NOR2_X1 us03_U318 (.ZN( us03_n527 ) , .A1( us03_n706 ) , .A2( us03_n777 ) );
  NOR2_X1 us03_U319 (.ZN( us03_n576 ) , .A1( us03_n706 ) , .A2( us03_n811 ) );
  NOR2_X1 us03_U32 (.ZN( us03_n802 ) , .A1( us03_n852 ) , .A2( us03_n859 ) );
  AOI21_X1 us03_U320 (.ZN( us03_n648 ) , .A( us03_n777 ) , .B1( us03_n790 ) , .B2( us03_n803 ) );
  NOR2_X1 us03_U321 (.ZN( us03_n682 ) , .A1( us03_n789 ) , .A2( us03_n811 ) );
  NOR2_X1 us03_U322 (.A2( us03_n811 ) , .A1( us03_n813 ) , .ZN( us03_n819 ) );
  AOI21_X1 us03_U323 (.A( us03_n788 ) , .B2( us03_n789 ) , .B1( us03_n790 ) , .ZN( us03_n791 ) );
  AOI21_X1 us03_U324 (.A( us03_n731 ) , .ZN( us03_n732 ) , .B2( us03_n778 ) , .B1( us03_n790 ) );
  NOR2_X1 us03_U325 (.ZN( us03_n565 ) , .A1( us03_n745 ) , .A2( us03_n803 ) );
  NOR2_X1 us03_U326 (.ZN( us03_n581 ) , .A1( us03_n790 ) , .A2( us03_n815 ) );
  NOR2_X1 us03_U327 (.ZN( us03_n532 ) , .A1( us03_n722 ) , .A2( us03_n786 ) );
  AOI21_X1 us03_U328 (.ZN( us03_n639 ) , .B1( us03_n678 ) , .A( us03_n789 ) , .B2( us03_n815 ) );
  NOR2_X1 us03_U329 (.ZN( us03_n709 ) , .A1( us03_n760 ) , .A2( us03_n761 ) );
  NAND4_X1 us03_U33 (.ZN( sa03_sr_7 ) , .A4( us03_n820 ) , .A3( us03_n821 ) , .A2( us03_n822 ) , .A1( us03_n823 ) );
  NOR2_X1 us03_U330 (.ZN( us03_n680 ) , .A2( us03_n706 ) , .A1( us03_n815 ) );
  INV_X1 us03_U331 (.A( us03_n695 ) , .ZN( us03_n836 ) );
  INV_X1 us03_U332 (.A( us03_n813 ) , .ZN( us03_n853 ) );
  AOI21_X1 us03_U333 (.ZN( us03_n440 ) , .A( us03_n697 ) , .B1( us03_n731 ) , .B2( us03_n748 ) );
  OAI21_X1 us03_U334 (.A( us03_n696 ) , .ZN( us03_n700 ) , .B2( us03_n748 ) , .B1( us03_n802 ) );
  OAI21_X1 us03_U335 (.ZN( us03_n696 ) , .B2( us03_n831 ) , .B1( us03_n836 ) , .A( us03_n858 ) );
  INV_X1 us03_U336 (.A( us03_n778 ) , .ZN( us03_n848 ) );
  AOI22_X1 us03_U337 (.A2( us03_n780 ) , .ZN( us03_n781 ) , .B2( us03_n829 ) , .A1( us03_n832 ) , .B1( us03_n861 ) );
  NAND2_X1 us03_U338 (.ZN( us03_n712 ) , .A1( us03_n726 ) , .A2( us03_n778 ) );
  NAND2_X1 us03_U339 (.ZN( us03_n751 ) , .A1( us03_n761 ) , .A2( us03_n803 ) );
  NOR4_X1 us03_U34 (.A4( us03_n816 ) , .A3( us03_n817 ) , .A2( us03_n818 ) , .A1( us03_n819 ) , .ZN( us03_n820 ) );
  NAND2_X1 us03_U340 (.A2( us03_n760 ) , .A1( us03_n804 ) , .ZN( us03_n808 ) );
  AOI21_X1 us03_U341 (.ZN( us03_n441 ) , .B1( us03_n787 ) , .B2( us03_n789 ) , .A( us03_n812 ) );
  NAND2_X2 us03_U342 (.A1( us03_n449 ) , .A2( us03_n460 ) , .ZN( us03_n788 ) );
  OAI21_X1 us03_U343 (.A( us03_n785 ) , .B2( us03_n786 ) , .B1( us03_n787 ) , .ZN( us03_n793 ) );
  OAI21_X1 us03_U344 (.ZN( us03_n785 ) , .A( us03_n837 ) , .B1( us03_n861 ) , .B2( us03_n871 ) );
  AOI21_X1 us03_U345 (.ZN( us03_n495 ) , .A( us03_n777 ) , .B2( us03_n789 ) , .B1( us03_n802 ) );
  NAND2_X2 us03_U346 (.A2( us03_n439 ) , .A1( us03_n445 ) , .ZN( us03_n782 ) );
  INV_X1 us03_U347 (.A( us03_n783 ) , .ZN( us03_n844 ) );
  NOR2_X1 us03_U348 (.ZN( us03_n468 ) , .A2( us03_n777 ) , .A1( us03_n813 ) );
  OAI21_X1 us03_U349 (.A( us03_n729 ) , .B1( us03_n730 ) , .ZN( us03_n734 ) , .B2( us03_n803 ) );
  AOI222_X1 us03_U35 (.C2( us03_n807 ) , .B2( us03_n808 ) , .A2( us03_n809 ) , .ZN( us03_n821 ) , .C1( us03_n830 ) , .A1( us03_n837 ) , .B1( us03_n851 ) );
  OAI21_X1 us03_U350 (.ZN( us03_n729 ) , .A( us03_n831 ) , .B2( us03_n850 ) , .B1( us03_n871 ) );
  NOR2_X1 us03_U351 (.ZN( us03_n524 ) , .A1( us03_n722 ) , .A2( us03_n748 ) );
  NOR2_X1 us03_U352 (.ZN( us03_n710 ) , .A2( us03_n722 ) , .A1( us03_n788 ) );
  NOR2_X1 us03_U353 (.ZN( us03_n482 ) , .A1( us03_n786 ) , .A2( us03_n803 ) );
  NAND2_X1 us03_U354 (.A1( us03_n697 ) , .A2( us03_n727 ) , .ZN( us03_n780 ) );
  NOR2_X1 us03_U355 (.ZN( us03_n516 ) , .A1( us03_n706 ) , .A2( us03_n786 ) );
  NAND2_X1 us03_U356 (.ZN( us03_n669 ) , .A1( us03_n804 ) , .A2( us03_n814 ) );
  NAND2_X1 us03_U357 (.A2( us03_n747 ) , .A1( us03_n784 ) , .ZN( us03_n807 ) );
  INV_X1 us03_U358 (.A( us03_n722 ) , .ZN( us03_n854 ) );
  INV_X1 us03_U359 (.A( us03_n815 ) , .ZN( us03_n842 ) );
  AOI211_X1 us03_U36 (.B( us03_n805 ) , .A( us03_n806 ) , .ZN( us03_n822 ) , .C1( us03_n840 ) , .C2( us03_n848 ) );
  AND2_X1 us03_U360 (.ZN( us03_n730 ) , .A1( us03_n777 ) , .A2( us03_n783 ) );
  NAND2_X1 us03_U361 (.A1( us03_n453 ) , .A2( us03_n469 ) , .ZN( us03_n801 ) );
  NAND2_X1 us03_U362 (.A1( us03_n449 ) , .A2( us03_n452 ) , .ZN( us03_n812 ) );
  NAND2_X1 us03_U363 (.A1( us03_n449 ) , .A2( us03_n469 ) , .ZN( us03_n814 ) );
  NAND2_X1 us03_U364 (.A1( us03_n452 ) , .A2( us03_n459 ) , .ZN( us03_n811 ) );
  NAND2_X1 us03_U365 (.A1( us03_n451 ) , .A2( us03_n459 ) , .ZN( us03_n742 ) );
  NAND2_X1 us03_U366 (.A1( us03_n450 ) , .A2( us03_n463 ) , .ZN( us03_n667 ) );
  NAND2_X1 us03_U367 (.A2( us03_n446 ) , .A1( us03_n458 ) , .ZN( us03_n726 ) );
  NAND2_X1 us03_U368 (.A1( us03_n453 ) , .A2( us03_n460 ) , .ZN( us03_n748 ) );
  NAND2_X1 us03_U369 (.A2( us03_n451 ) , .A1( us03_n453 ) , .ZN( us03_n804 ) );
  NOR2_X1 us03_U37 (.ZN( us03_n746 ) , .A1( us03_n859 ) , .A2( us03_n860 ) );
  NAND2_X1 us03_U370 (.A2( us03_n452 ) , .A1( us03_n470 ) , .ZN( us03_n777 ) );
  NAND2_X1 us03_U371 (.A1( us03_n451 ) , .A2( us03_n470 ) , .ZN( us03_n783 ) );
  NAND2_X1 us03_U372 (.A2( us03_n462 ) , .A1( us03_n463 ) , .ZN( us03_n810 ) );
  NAND2_X1 us03_U373 (.A1( us03_n439 ) , .A2( us03_n458 ) , .ZN( us03_n697 ) );
  NAND2_X1 us03_U374 (.A2( us03_n447 ) , .A1( us03_n450 ) , .ZN( us03_n761 ) );
  NAND2_X1 us03_U375 (.A2( us03_n446 ) , .A1( us03_n450 ) , .ZN( us03_n727 ) );
  NOR2_X1 us03_U376 (.ZN( us03_n445 ) , .A2( us03_n847 ) , .A1( us03_n856 ) );
  NAND2_X1 us03_U377 (.A2( us03_n459 ) , .A1( us03_n460 ) , .ZN( us03_n745 ) );
  NAND2_X1 us03_U378 (.A1( us03_n460 ) , .A2( us03_n470 ) , .ZN( us03_n786 ) );
  NOR2_X1 us03_U379 (.ZN( us03_n463 ) , .A2( us03_n845 ) , .A1( us03_n846 ) );
  NOR2_X1 us03_U38 (.ZN( us03_n623 ) , .A2( us03_n834 ) , .A1( us03_n837 ) );
  NAND2_X2 us03_U380 (.A2( us03_n459 ) , .A1( us03_n469 ) , .ZN( us03_n695 ) );
  NOR2_X1 us03_U381 (.ZN( us03_n451 ) , .A1( us03_n824 ) , .A2( us03_n825 ) );
  NOR2_X1 us03_U382 (.ZN( us03_n449 ) , .A1( us03_n826 ) , .A2( us03_n827 ) );
  NAND2_X1 us03_U383 (.A2( us03_n452 ) , .A1( us03_n453 ) , .ZN( us03_n728 ) );
  NAND2_X2 us03_U384 (.A2( us03_n446 ) , .A1( us03_n462 ) , .ZN( us03_n813 ) );
  NAND2_X2 us03_U385 (.A2( us03_n439 ) , .A1( us03_n450 ) , .ZN( us03_n789 ) );
  NAND2_X2 us03_U386 (.A1( us03_n447 ) , .A2( us03_n462 ) , .ZN( us03_n722 ) );
  NAND2_X2 us03_U387 (.A1( us03_n447 ) , .A2( us03_n458 ) , .ZN( us03_n790 ) );
  NAND2_X2 us03_U388 (.A1( us03_n439 ) , .A2( us03_n462 ) , .ZN( us03_n706 ) );
  NAND2_X2 us03_U389 (.A2( us03_n469 ) , .A1( us03_n470 ) , .ZN( us03_n815 ) );
  NAND4_X1 us03_U39 (.A4( us03_n601 ) , .A3( us03_n602 ) , .A2( us03_n603 ) , .A1( us03_n604 ) , .ZN( us03_n720 ) );
  NAND2_X2 us03_U390 (.A2( us03_n458 ) , .A1( us03_n463 ) , .ZN( us03_n778 ) );
  NAND2_X1 us03_U391 (.A1( us03_n445 ) , .A2( us03_n447 ) , .ZN( us03_n803 ) );
  NAND2_X2 us03_U392 (.A1( us03_n445 ) , .A2( us03_n446 ) , .ZN( us03_n784 ) );
  NOR2_X1 us03_U393 (.A2( sa03_6 ) , .A1( sa03_7 ) , .ZN( us03_n462 ) );
  NOR2_X1 us03_U394 (.A2( sa03_4 ) , .ZN( us03_n447 ) , .A1( us03_n846 ) );
  NOR2_X1 us03_U395 (.A2( sa03_5 ) , .ZN( us03_n446 ) , .A1( us03_n845 ) );
  NOR2_X1 us03_U396 (.A2( sa03_7 ) , .ZN( us03_n458 ) , .A1( us03_n847 ) );
  NOR2_X1 us03_U397 (.A2( sa03_4 ) , .A1( sa03_5 ) , .ZN( us03_n439 ) );
  NOR2_X1 us03_U398 (.A2( sa03_1 ) , .ZN( us03_n469 ) , .A1( us03_n824 ) );
  NOR2_X1 us03_U399 (.A2( sa03_2 ) , .A1( sa03_3 ) , .ZN( us03_n470 ) );
  NOR3_X1 us03_U4 (.A3( us03_n798 ) , .A2( us03_n799 ) , .A1( us03_n800 ) , .ZN( us03_n823 ) );
  NOR3_X1 us03_U40 (.A1( us03_n597 ) , .ZN( us03_n602 ) , .A3( us03_n661 ) , .A2( us03_n768 ) );
  NOR2_X1 us03_U400 (.A2( sa03_6 ) , .ZN( us03_n450 ) , .A1( us03_n856 ) );
  NOR2_X1 us03_U401 (.A2( sa03_2 ) , .ZN( us03_n459 ) , .A1( us03_n827 ) );
  NOR2_X1 us03_U402 (.A2( sa03_0 ) , .ZN( us03_n452 ) , .A1( us03_n825 ) );
  NOR2_X1 us03_U403 (.A2( sa03_0 ) , .A1( sa03_1 ) , .ZN( us03_n460 ) );
  NOR2_X1 us03_U404 (.A2( sa03_3 ) , .ZN( us03_n453 ) , .A1( us03_n826 ) );
  INV_X1 us03_U405 (.A( sa03_6 ) , .ZN( us03_n847 ) );
  INV_X1 us03_U406 (.A( sa03_3 ) , .ZN( us03_n827 ) );
  INV_X1 us03_U407 (.A( sa03_1 ) , .ZN( us03_n825 ) );
  INV_X1 us03_U408 (.A( sa03_0 ) , .ZN( us03_n824 ) );
  INV_X1 us03_U409 (.A( sa03_2 ) , .ZN( us03_n826 ) );
  NOR4_X1 us03_U41 (.A3( us03_n598 ) , .A2( us03_n599 ) , .A1( us03_n600 ) , .ZN( us03_n601 ) , .A4( us03_n653 ) );
  INV_X1 us03_U410 (.A( sa03_7 ) , .ZN( us03_n856 ) );
  INV_X1 us03_U411 (.A( sa03_5 ) , .ZN( us03_n846 ) );
  AOI222_X1 us03_U412 (.ZN( us03_n603 ) , .B2( us03_n669 ) , .B1( us03_n751 ) , .C2( us03_n829 ) , .A1( us03_n831 ) , .A2( us03_n860 ) , .C1( us03_n861 ) );
  AOI222_X1 us03_U413 (.ZN( us03_n511 ) , .C1( us03_n830 ) , .B2( us03_n835 ) , .A2( us03_n841 ) , .C2( us03_n860 ) , .B1( us03_n861 ) , .A1( us03_n864 ) );
  AOI221_X1 us03_U414 (.A( us03_n481 ) , .ZN( us03_n486 ) , .B1( us03_n829 ) , .C2( us03_n842 ) , .C1( us03_n850 ) , .B2( us03_n860 ) );
  NOR2_X1 us03_U415 (.ZN( us03_n787 ) , .A2( us03_n860 ) , .A1( us03_n866 ) );
  NAND4_X1 us03_U416 (.ZN( sa03_sr_2 ) , .A4( us03_n641 ) , .A3( us03_n642 ) , .A2( us03_n643 ) , .A1( us03_n644 ) );
  OAI221_X1 us03_U417 (.A( us03_n781 ) , .C2( us03_n782 ) , .B2( us03_n783 ) , .B1( us03_n784 ) , .ZN( us03_n794 ) , .C1( us03_n811 ) );
  NAND2_X1 us03_U418 (.A1( us03_n727 ) , .A2( us03_n782 ) , .ZN( us03_n809 ) );
  OAI22_X1 us03_U419 (.ZN( us03_n586 ) , .A2( us03_n745 ) , .B2( us03_n760 ) , .A1( us03_n761 ) , .B1( us03_n782 ) );
  AOI222_X1 us03_U42 (.ZN( us03_n604 ) , .A1( us03_n828 ) , .C2( us03_n835 ) , .B1( us03_n840 ) , .A2( us03_n854 ) , .B2( us03_n859 ) , .C1( us03_n866 ) );
  OAI221_X1 us03_U420 (.A( us03_n694 ) , .ZN( us03_n701 ) , .C2( us03_n782 ) , .C1( us03_n783 ) , .B1( us03_n784 ) , .B2( us03_n804 ) );
  AOI21_X1 us03_U421 (.ZN( us03_n590 ) , .B1( us03_n726 ) , .B2( us03_n782 ) , .A( us03_n788 ) );
  AOI21_X1 us03_U422 (.ZN( us03_n621 ) , .B1( us03_n697 ) , .A( us03_n777 ) , .B2( us03_n782 ) );
  AOI21_X1 us03_U423 (.ZN( us03_n646 ) , .A( us03_n760 ) , .B2( us03_n782 ) , .B1( us03_n790 ) );
  OAI22_X1 us03_U424 (.ZN( us03_n679 ) , .A1( us03_n697 ) , .A2( us03_n728 ) , .B2( us03_n782 ) , .B1( us03_n815 ) );
  OAI21_X1 us03_U425 (.A( us03_n611 ) , .ZN( us03_n614 ) , .B1( us03_n623 ) , .B2( us03_n782 ) );
  NOR2_X1 us03_U426 (.ZN( us03_n608 ) , .A1( us03_n782 ) , .A2( us03_n814 ) );
  OAI222_X1 us03_U427 (.A2( us03_n667 ) , .ZN( us03_n672 ) , .B1( us03_n745 ) , .B2( us03_n782 ) , .C2( us03_n786 ) , .C1( us03_n813 ) , .A1( us03_n815 ) );
  NOR2_X1 us03_U428 (.ZN( us03_n649 ) , .A1( us03_n782 ) , .A2( us03_n786 ) );
  NOR2_X1 us03_U429 (.ZN( us03_n598 ) , .A2( us03_n695 ) , .A1( us03_n782 ) );
  NAND4_X1 us03_U43 (.ZN( sa03_sr_3 ) , .A4( us03_n702 ) , .A3( us03_n703 ) , .A2( us03_n704 ) , .A1( us03_n705 ) );
  NOR2_X1 us03_U430 (.ZN( us03_n551 ) , .A2( us03_n742 ) , .A1( us03_n782 ) );
  INV_X1 us03_U431 (.A( us03_n782 ) , .ZN( us03_n859 ) );
  AOI221_X1 us03_U432 (.A( us03_n574 ) , .ZN( us03_n585 ) , .B2( us03_n829 ) , .C2( us03_n841 ) , .B1( us03_n852 ) , .C1( us03_n859 ) );
  AOI21_X1 us03_U433 (.ZN( us03_n574 ) , .B2( us03_n722 ) , .B1( us03_n746 ) , .A( us03_n783 ) );
  AOI211_X1 us03_U434 (.A( us03_n635 ) , .ZN( us03_n643 ) , .B( us03_n741 ) , .C2( us03_n837 ) , .C1( us03_n852 ) );
  NAND4_X1 us03_U435 (.A4( us03_n631 ) , .A3( us03_n632 ) , .A2( us03_n633 ) , .A1( us03_n634 ) , .ZN( us03_n741 ) );
  INV_X1 us03_U436 (.A( sa03_4 ) , .ZN( us03_n845 ) );
  NAND3_X1 us03_U437 (.ZN( sa03_sr_6 ) , .A3( us03_n795 ) , .A2( us03_n796 ) , .A1( us03_n797 ) );
  NAND3_X1 us03_U438 (.ZN( sa03_sr_5 ) , .A3( us03_n756 ) , .A2( us03_n757 ) , .A1( us03_n758 ) );
  NAND3_X1 us03_U439 (.ZN( sa03_sr_4 ) , .A3( us03_n736 ) , .A2( us03_n737 ) , .A1( us03_n738 ) );
  NOR4_X1 us03_U44 (.A4( us03_n698 ) , .A3( us03_n699 ) , .A2( us03_n700 ) , .A1( us03_n701 ) , .ZN( us03_n702 ) );
  NAND3_X1 us03_U440 (.A3( us03_n673 ) , .A2( us03_n674 ) , .A1( us03_n675 ) , .ZN( us03_n805 ) );
  NAND3_X1 us03_U441 (.ZN( us03_n636 ) , .A3( us03_n706 ) , .A2( us03_n722 ) , .A1( us03_n790 ) );
  NAND3_X1 us03_U442 (.A3( us03_n616 ) , .A2( us03_n617 ) , .A1( us03_n618 ) , .ZN( us03_n723 ) );
  NAND3_X1 us03_U443 (.A3( us03_n583 ) , .A2( us03_n584 ) , .A1( us03_n585 ) , .ZN( us03_n619 ) );
  NAND3_X1 us03_U444 (.ZN( us03_n563 ) , .A3( us03_n678 ) , .A2( us03_n748 ) , .A1( us03_n783 ) );
  NAND3_X1 us03_U445 (.A3( us03_n521 ) , .A2( us03_n522 ) , .A1( us03_n523 ) , .ZN( us03_n740 ) );
  NAND3_X1 us03_U446 (.A3( us03_n510 ) , .A1( us03_n511 ) , .ZN( us03_n606 ) , .A2( us03_n869 ) );
  NAND3_X1 us03_U447 (.A3( us03_n465 ) , .A2( us03_n466 ) , .A1( us03_n467 ) , .ZN( us03_n775 ) );
  AOI211_X1 us03_U45 (.B( us03_n692 ) , .A( us03_n693 ) , .ZN( us03_n703 ) , .C2( us03_n829 ) , .C1( us03_n849 ) );
  NOR2_X1 us03_U46 (.ZN( us03_n705 ) , .A2( us03_n774 ) , .A1( us03_n798 ) );
  AOI222_X1 us03_U47 (.ZN( us03_n467 ) , .B1( us03_n830 ) , .A1( us03_n837 ) , .C1( us03_n840 ) , .C2( us03_n849 ) , .A2( us03_n853 ) , .B2( us03_n863 ) );
  NOR4_X1 us03_U48 (.A1( us03_n464 ) , .ZN( us03_n465 ) , .A4( us03_n540 ) , .A2( us03_n552 ) , .A3( us03_n612 ) );
  AOI221_X1 us03_U49 (.ZN( us03_n466 ) , .C2( us03_n712 ) , .B2( us03_n829 ) , .C1( us03_n843 ) , .B1( us03_n858 ) , .A( us03_n862 ) );
  NOR3_X1 us03_U5 (.ZN( us03_n502 ) , .A2( us03_n677 ) , .A3( us03_n775 ) , .A1( us03_n874 ) );
  NOR4_X1 us03_U50 (.A4( us03_n575 ) , .A3( us03_n576 ) , .A2( us03_n577 ) , .ZN( us03_n584 ) , .A1( us03_n681 ) );
  NOR4_X1 us03_U51 (.A1( us03_n582 ) , .ZN( us03_n583 ) , .A3( us03_n650 ) , .A2( us03_n660 ) , .A4( us03_n765 ) );
  NAND4_X1 us03_U52 (.A4( us03_n483 ) , .A3( us03_n484 ) , .A2( us03_n485 ) , .A1( us03_n486 ) , .ZN( us03_n776 ) );
  NOR4_X1 us03_U53 (.A4( us03_n482 ) , .ZN( us03_n485 ) , .A1( us03_n564 ) , .A2( us03_n579 ) , .A3( us03_n600 ) );
  NOR4_X1 us03_U54 (.ZN( us03_n484 ) , .A1( us03_n505 ) , .A2( us03_n517 ) , .A4( us03_n544 ) , .A3( us03_n609 ) );
  NOR4_X1 us03_U55 (.ZN( us03_n483 ) , .A2( us03_n531 ) , .A1( us03_n556 ) , .A3( us03_n629 ) , .A4( us03_n716 ) );
  AOI211_X1 us03_U56 (.B( us03_n621 ) , .A( us03_n622 ) , .ZN( us03_n633 ) , .C2( us03_n834 ) , .C1( us03_n861 ) );
  NOR4_X1 us03_U57 (.A4( us03_n627 ) , .A3( us03_n628 ) , .A2( us03_n629 ) , .A1( us03_n630 ) , .ZN( us03_n631 ) );
  NOR4_X1 us03_U58 (.A4( us03_n624 ) , .A3( us03_n625 ) , .A2( us03_n626 ) , .ZN( us03_n632 ) , .A1( us03_n662 ) );
  NAND4_X1 us03_U59 (.A4( us03_n655 ) , .A3( us03_n656 ) , .A2( us03_n657 ) , .A1( us03_n658 ) , .ZN( us03_n798 ) );
  INV_X1 us03_U6 (.A( us03_n704 ) , .ZN( us03_n874 ) );
  NOR3_X1 us03_U60 (.A3( us03_n646 ) , .A2( us03_n647 ) , .A1( us03_n648 ) , .ZN( us03_n657 ) );
  NOR3_X1 us03_U61 (.A3( us03_n649 ) , .A2( us03_n650 ) , .A1( us03_n651 ) , .ZN( us03_n656 ) );
  NOR3_X1 us03_U62 (.A3( us03_n652 ) , .A2( us03_n653 ) , .A1( us03_n654 ) , .ZN( us03_n655 ) );
  NAND4_X1 us03_U63 (.A4( us03_n558 ) , .A3( us03_n559 ) , .A2( us03_n560 ) , .A1( us03_n561 ) , .ZN( us03_n605 ) );
  NOR4_X1 us03_U64 (.A4( us03_n554 ) , .A3( us03_n555 ) , .A2( us03_n556 ) , .A1( us03_n557 ) , .ZN( us03_n558 ) );
  NOR4_X1 us03_U65 (.ZN( us03_n559 ) , .A1( us03_n651 ) , .A3( us03_n659 ) , .A4( us03_n683 ) , .A2( us03_n766 ) );
  NOR4_X1 us03_U66 (.A4( us03_n550 ) , .A3( us03_n551 ) , .A2( us03_n552 ) , .A1( us03_n553 ) , .ZN( us03_n560 ) );
  NAND4_X1 us03_U67 (.A4( us03_n770 ) , .A3( us03_n771 ) , .A2( us03_n772 ) , .A1( us03_n773 ) , .ZN( us03_n799 ) );
  NOR3_X1 us03_U68 (.A3( us03_n763 ) , .A2( us03_n764 ) , .A1( us03_n765 ) , .ZN( us03_n771 ) );
  NOR4_X1 us03_U69 (.A4( us03_n766 ) , .A3( us03_n767 ) , .A2( us03_n768 ) , .A1( us03_n769 ) , .ZN( us03_n770 ) );
  NOR3_X1 us03_U7 (.A3( us03_n619 ) , .A2( us03_n620 ) , .ZN( us03_n634 ) , .A1( us03_n723 ) );
  AOI222_X1 us03_U70 (.ZN( us03_n773 ) , .A1( us03_n828 ) , .C1( us03_n832 ) , .B2( us03_n839 ) , .A2( us03_n848 ) , .B1( us03_n859 ) , .C2( us03_n871 ) );
  NOR4_X1 us03_U71 (.A4( us03_n507 ) , .A2( us03_n508 ) , .A1( us03_n509 ) , .ZN( us03_n510 ) , .A3( us03_n668 ) );
  INV_X1 us03_U72 (.A( us03_n503 ) , .ZN( us03_n869 ) );
  NOR4_X1 us03_U73 (.A4( us03_n663 ) , .A3( us03_n664 ) , .A2( us03_n665 ) , .A1( us03_n666 ) , .ZN( us03_n674 ) );
  NOR4_X1 us03_U74 (.A4( us03_n659 ) , .A3( us03_n660 ) , .A2( us03_n661 ) , .A1( us03_n662 ) , .ZN( us03_n675 ) );
  NOR4_X1 us03_U75 (.A3( us03_n671 ) , .A1( us03_n672 ) , .ZN( us03_n673 ) , .A4( us03_n713 ) , .A2( us03_n857 ) );
  NOR2_X1 us03_U76 (.ZN( us03_n759 ) , .A1( us03_n831 ) , .A2( us03_n832 ) );
  NOR4_X1 us03_U77 (.A4( us03_n732 ) , .A3( us03_n733 ) , .A2( us03_n734 ) , .A1( us03_n735 ) , .ZN( us03_n736 ) );
  AOI211_X1 us03_U78 (.B( us03_n723 ) , .A( us03_n724 ) , .ZN( us03_n737 ) , .C1( us03_n841 ) , .C2( us03_n853 ) );
  NOR3_X1 us03_U79 (.A3( us03_n720 ) , .A1( us03_n721 ) , .ZN( us03_n738 ) , .A2( us03_n739 ) );
  NOR2_X1 us03_U8 (.ZN( us03_n573 ) , .A1( us03_n620 ) , .A2( us03_n743 ) );
  NOR4_X1 us03_U80 (.A3( us03_n753 ) , .A2( us03_n754 ) , .A1( us03_n755 ) , .ZN( us03_n756 ) , .A4( us03_n867 ) );
  AOI211_X1 us03_U81 (.B( us03_n743 ) , .A( us03_n744 ) , .ZN( us03_n757 ) , .C1( us03_n830 ) , .C2( us03_n851 ) );
  NOR3_X1 us03_U82 (.A3( us03_n739 ) , .A2( us03_n740 ) , .A1( us03_n741 ) , .ZN( us03_n758 ) );
  NAND4_X1 us03_U83 (.A4( us03_n454 ) , .A3( us03_n455 ) , .A2( us03_n456 ) , .A1( us03_n457 ) , .ZN( us03_n677 ) );
  NOR3_X1 us03_U84 (.ZN( us03_n455 ) , .A3( us03_n528 ) , .A1( us03_n553 ) , .A2( us03_n568 ) );
  AOI221_X1 us03_U85 (.A( us03_n448 ) , .ZN( us03_n457 ) , .C2( us03_n751 ) , .B1( us03_n830 ) , .C1( us03_n840 ) , .B2( us03_n859 ) );
  NOR4_X1 us03_U86 (.ZN( us03_n456 ) , .A2( us03_n507 ) , .A1( us03_n597 ) , .A4( us03_n626 ) , .A3( us03_n709 ) );
  NAND4_X1 us03_U87 (.A4( us03_n533 ) , .A3( us03_n534 ) , .A2( us03_n535 ) , .A1( us03_n536 ) , .ZN( us03_n620 ) );
  NOR4_X1 us03_U88 (.A4( us03_n524 ) , .A2( us03_n525 ) , .A1( us03_n526 ) , .ZN( us03_n536 ) , .A3( us03_n699 ) );
  NOR4_X1 us03_U89 (.A1( us03_n529 ) , .ZN( us03_n534 ) , .A2( us03_n652 ) , .A4( us03_n666 ) , .A3( us03_n763 ) );
  NOR2_X1 us03_U9 (.A1( us03_n676 ) , .ZN( us03_n691 ) , .A2( us03_n805 ) );
  NOR4_X1 us03_U90 (.A4( us03_n527 ) , .A3( us03_n528 ) , .ZN( us03_n535 ) , .A2( us03_n682 ) , .A1( us03_n792 ) );
  NAND4_X1 us03_U91 (.A4( us03_n477 ) , .A3( us03_n478 ) , .A2( us03_n479 ) , .A1( us03_n480 ) , .ZN( us03_n692 ) );
  NOR3_X1 us03_U92 (.ZN( us03_n478 ) , .A2( us03_n506 ) , .A3( us03_n599 ) , .A1( us03_n608 ) );
  AOI211_X1 us03_U93 (.B( us03_n475 ) , .A( us03_n476 ) , .ZN( us03_n480 ) , .C2( us03_n831 ) , .C1( us03_n859 ) );
  NOR4_X1 us03_U94 (.ZN( us03_n479 ) , .A3( us03_n530 ) , .A4( us03_n543 ) , .A2( us03_n565 ) , .A1( us03_n715 ) );
  NAND4_X1 us03_U95 (.A4( us03_n546 ) , .A3( us03_n547 ) , .A2( us03_n548 ) , .A1( us03_n549 ) , .ZN( us03_n743 ) );
  NOR3_X1 us03_U96 (.ZN( us03_n547 ) , .A2( us03_n649 ) , .A1( us03_n665 ) , .A3( us03_n769 ) );
  AOI211_X1 us03_U97 (.B( us03_n537 ) , .A( us03_n538 ) , .ZN( us03_n549 ) , .C2( us03_n837 ) , .C1( us03_n849 ) );
  NOR4_X1 us03_U98 (.A4( us03_n542 ) , .A3( us03_n543 ) , .A2( us03_n544 ) , .A1( us03_n545 ) , .ZN( us03_n546 ) );
  NOR4_X1 us03_U99 (.ZN( us03_n618 ) , .A1( us03_n654 ) , .A3( us03_n664 ) , .A4( us03_n680 ) , .A2( us03_n764 ) );
  NOR3_X1 us12_U10 (.ZN( us12_n504 ) , .A2( us12_n679 ) , .A3( us12_n777 ) , .A1( us12_n876 ) );
  NOR4_X1 us12_U100 (.A4( us12_n529 ) , .A3( us12_n530 ) , .ZN( us12_n537 ) , .A2( us12_n684 ) , .A1( us12_n794 ) );
  NAND4_X1 us12_U101 (.A4( us12_n479 ) , .A3( us12_n480 ) , .A2( us12_n481 ) , .A1( us12_n482 ) , .ZN( us12_n694 ) );
  NOR3_X1 us12_U102 (.ZN( us12_n480 ) , .A2( us12_n508 ) , .A3( us12_n601 ) , .A1( us12_n610 ) );
  AOI211_X1 us12_U103 (.B( us12_n477 ) , .A( us12_n478 ) , .ZN( us12_n482 ) , .C2( us12_n833 ) , .C1( us12_n861 ) );
  NOR4_X1 us12_U104 (.ZN( us12_n481 ) , .A3( us12_n532 ) , .A4( us12_n545 ) , .A2( us12_n567 ) , .A1( us12_n717 ) );
  NAND4_X1 us12_U105 (.A4( us12_n548 ) , .A3( us12_n549 ) , .A2( us12_n550 ) , .A1( us12_n551 ) , .ZN( us12_n745 ) );
  NOR3_X1 us12_U106 (.ZN( us12_n549 ) , .A2( us12_n651 ) , .A1( us12_n667 ) , .A3( us12_n771 ) );
  AOI211_X1 us12_U107 (.B( us12_n539 ) , .A( us12_n540 ) , .ZN( us12_n551 ) , .C2( us12_n839 ) , .C1( us12_n851 ) );
  NOR4_X1 us12_U108 (.A4( us12_n541 ) , .A3( us12_n542 ) , .A2( us12_n543 ) , .ZN( us12_n550 ) , .A1( us12_n688 ) );
  NOR4_X1 us12_U109 (.ZN( us12_n620 ) , .A1( us12_n656 ) , .A3( us12_n666 ) , .A4( us12_n682 ) , .A2( us12_n766 ) );
  INV_X1 us12_U11 (.A( us12_n706 ) , .ZN( us12_n876 ) );
  NOR4_X1 us12_U110 (.A4( us12_n609 ) , .A3( us12_n610 ) , .A2( us12_n611 ) , .A1( us12_n612 ) , .ZN( us12_n619 ) );
  NOR4_X1 us12_U111 (.A4( us12_n614 ) , .A3( us12_n615 ) , .A2( us12_n616 ) , .A1( us12_n617 ) , .ZN( us12_n618 ) );
  NOR2_X1 us12_U112 (.ZN( us12_n686 ) , .A1( us12_n831 ) , .A2( us12_n832 ) );
  NAND4_X1 us12_U113 (.A4( us12_n485 ) , .A3( us12_n486 ) , .A2( us12_n487 ) , .A1( us12_n488 ) , .ZN( us12_n778 ) );
  NOR4_X1 us12_U114 (.A4( us12_n484 ) , .ZN( us12_n487 ) , .A1( us12_n566 ) , .A2( us12_n581 ) , .A3( us12_n602 ) );
  NOR4_X1 us12_U115 (.ZN( us12_n486 ) , .A1( us12_n507 ) , .A2( us12_n519 ) , .A4( us12_n546 ) , .A3( us12_n611 ) );
  NOR4_X1 us12_U116 (.ZN( us12_n485 ) , .A2( us12_n533 ) , .A1( us12_n558 ) , .A3( us12_n631 ) , .A4( us12_n718 ) );
  NAND4_X1 us12_U117 (.A4( us12_n691 ) , .A3( us12_n692 ) , .A1( us12_n693 ) , .ZN( us12_n776 ) , .A2( us12_n872 ) );
  AOI221_X1 us12_U118 (.A( us12_n681 ) , .ZN( us12_n692 ) , .B2( us12_n840 ) , .C1( us12_n842 ) , .C2( us12_n862 ) , .B1( us12_n865 ) );
  INV_X1 us12_U119 (.A( us12_n679 ) , .ZN( us12_n872 ) );
  NOR3_X1 us12_U12 (.A3( us12_n621 ) , .A2( us12_n622 ) , .ZN( us12_n636 ) , .A1( us12_n725 ) );
  NOR4_X1 us12_U120 (.A4( us12_n687 ) , .A3( us12_n688 ) , .A2( us12_n689 ) , .A1( us12_n690 ) , .ZN( us12_n691 ) );
  NAND4_X1 us12_U121 (.A4( us12_n719 ) , .A3( us12_n720 ) , .A2( us12_n721 ) , .ZN( us12_n741 ) , .A1( us12_n857 ) );
  INV_X1 us12_U122 (.A( us12_n709 ) , .ZN( us12_n857 ) );
  AOI221_X1 us12_U123 (.A( us12_n710 ) , .ZN( us12_n721 ) , .C2( us12_n844 ) , .B2( us12_n845 ) , .C1( us12_n861 ) , .B1( us12_n862 ) );
  NOR4_X1 us12_U124 (.A4( us12_n715 ) , .A3( us12_n716 ) , .A2( us12_n717 ) , .A1( us12_n718 ) , .ZN( us12_n719 ) );
  NAND4_X1 us12_U125 (.A4( us12_n473 ) , .A3( us12_n474 ) , .A2( us12_n475 ) , .A1( us12_n476 ) , .ZN( us12_n678 ) );
  NOR4_X1 us12_U126 (.ZN( us12_n475 ) , .A1( us12_n531 ) , .A3( us12_n568 ) , .A4( us12_n600 ) , .A2( us12_n642 ) );
  NOR4_X1 us12_U127 (.A4( us12_n470 ) , .ZN( us12_n476 ) , .A3( us12_n556 ) , .A1( us12_n735 ) , .A2( us12_n755 ) );
  NOR4_X1 us12_U128 (.ZN( us12_n474 ) , .A1( us12_n506 ) , .A3( us12_n544 ) , .A2( us12_n583 ) , .A4( us12_n716 ) );
  NOR2_X1 us12_U129 (.ZN( us12_n733 ) , .A2( us12_n832 ) , .A1( us12_n845 ) );
  NOR2_X1 us12_U13 (.ZN( us12_n495 ) , .A1( us12_n678 ) , .A2( us12_n694 ) );
  NOR2_X1 us12_U130 (.ZN( us12_n789 ) , .A2( us12_n862 ) , .A1( us12_n868 ) );
  NAND4_X1 us12_U131 (.A4( us12_n573 ) , .A3( us12_n574 ) , .A1( us12_n575 ) , .ZN( us12_n723 ) , .A2( us12_n874 ) );
  NOR4_X1 us12_U132 (.A4( us12_n569 ) , .A3( us12_n570 ) , .A2( us12_n571 ) , .A1( us12_n572 ) , .ZN( us12_n573 ) );
  AOI221_X1 us12_U133 (.A( us12_n564 ) , .C2( us12_n565 ) , .ZN( us12_n574 ) , .B2( us12_n845 ) , .B1( us12_n852 ) , .C1( us12_n853 ) );
  NOR2_X1 us12_U134 (.ZN( us12_n575 ) , .A1( us12_n622 ) , .A2( us12_n745 ) );
  NAND4_X1 us12_U135 (.A4( us12_n633 ) , .A3( us12_n634 ) , .A2( us12_n635 ) , .A1( us12_n636 ) , .ZN( us12_n743 ) );
  AOI211_X1 us12_U136 (.B( us12_n623 ) , .A( us12_n624 ) , .ZN( us12_n635 ) , .C2( us12_n836 ) , .C1( us12_n863 ) );
  NOR4_X1 us12_U137 (.A4( us12_n629 ) , .A3( us12_n630 ) , .A2( us12_n631 ) , .A1( us12_n632 ) , .ZN( us12_n633 ) );
  NOR4_X1 us12_U138 (.A4( us12_n626 ) , .A3( us12_n627 ) , .A2( us12_n628 ) , .ZN( us12_n634 ) , .A1( us12_n664 ) );
  NAND4_X1 us12_U139 (.A4( us12_n493 ) , .A3( us12_n494 ) , .A1( us12_n495 ) , .ZN( us12_n802 ) , .A2( us12_n867 ) );
  NOR2_X1 us12_U14 (.A1( us12_n678 ) , .ZN( us12_n693 ) , .A2( us12_n807 ) );
  AOI221_X1 us12_U140 (.A( us12_n489 ) , .ZN( us12_n494 ) , .B2( us12_n836 ) , .C2( us12_n841 ) , .C1( us12_n851 ) , .B1( us12_n860 ) );
  INV_X1 us12_U141 (.A( us12_n778 ) , .ZN( us12_n867 ) );
  NOR4_X1 us12_U142 (.A2( us12_n491 ) , .A1( us12_n492 ) , .ZN( us12_n493 ) , .A3( us12_n580 ) , .A4( us12_n612 ) );
  NOR4_X1 us12_U143 (.A3( us12_n755 ) , .A2( us12_n756 ) , .A1( us12_n757 ) , .ZN( us12_n758 ) , .A4( us12_n869 ) );
  AOI211_X1 us12_U144 (.B( us12_n745 ) , .A( us12_n746 ) , .ZN( us12_n759 ) , .C1( us12_n832 ) , .C2( us12_n853 ) );
  NOR3_X1 us12_U145 (.A3( us12_n741 ) , .A2( us12_n742 ) , .A1( us12_n743 ) , .ZN( us12_n760 ) );
  NOR2_X1 us12_U146 (.ZN( us12_n647 ) , .A1( us12_n854 ) , .A2( us12_n868 ) );
  INV_X1 us12_U147 (.A( us12_n762 ) , .ZN( us12_n830 ) );
  INV_X1 us12_U148 (.A( us12_n754 ) , .ZN( us12_n869 ) );
  OAI21_X1 us12_U149 (.B1( us12_n753 ) , .ZN( us12_n754 ) , .A( us12_n845 ) , .B2( us12_n868 ) );
  INV_X1 us12_U15 (.A( us12_n607 ) , .ZN( us12_n874 ) );
  OR4_X1 us12_U150 (.ZN( us12_n466 ) , .A4( us12_n518 ) , .A3( us12_n529 ) , .A2( us12_n578 ) , .A1( us12_n712 ) );
  OR4_X1 us12_U151 (.A4( us12_n566 ) , .A3( us12_n567 ) , .A2( us12_n568 ) , .ZN( us12_n572 ) , .A1( us12_n665 ) );
  OR4_X1 us12_U152 (.ZN( us12_n492 ) , .A4( us12_n534 ) , .A2( us12_n547 ) , .A1( us12_n559 ) , .A3( us12_n632 ) );
  OR4_X1 us12_U153 (.A4( us12_n518 ) , .A2( us12_n519 ) , .A1( us12_n520 ) , .ZN( us12_n522 ) , .A3( us12_n821 ) );
  OR4_X1 us12_U154 (.A4( us12_n682 ) , .A3( us12_n683 ) , .A2( us12_n684 ) , .A1( us12_n685 ) , .ZN( us12_n690 ) );
  OR4_X1 us12_U155 (.A4( us12_n580 ) , .A3( us12_n581 ) , .A2( us12_n582 ) , .A1( us12_n583 ) , .ZN( us12_n584 ) );
  NAND2_X1 us12_U156 (.ZN( us12_n613 ) , .A2( us12_n837 ) , .A1( us12_n873 ) );
  OR3_X1 us12_U157 (.A3( us12_n506 ) , .A2( us12_n507 ) , .A1( us12_n508 ) , .ZN( us12_n511 ) );
  INV_X1 us12_U158 (.A( us12_n463 ) , .ZN( us12_n864 ) );
  OAI21_X1 us12_U159 (.ZN( us12_n463 ) , .B1( us12_n809 ) , .A( us12_n834 ) , .B2( us12_n851 ) );
  INV_X1 us12_U16 (.A( us12_n680 ) , .ZN( us12_n840 ) );
  INV_X1 us12_U160 (.A( us12_n672 ) , .ZN( us12_n859 ) );
  AOI21_X1 us12_U161 (.A( us12_n670 ) , .B1( us12_n671 ) , .ZN( us12_n672 ) , .B2( us12_n856 ) );
  OAI222_X1 us12_U162 (.B2( us12_n708 ) , .ZN( us12_n709 ) , .C2( us12_n724 ) , .B1( us12_n747 ) , .A1( us12_n806 ) , .C1( us12_n814 ) , .A2( us12_n815 ) );
  AOI22_X1 us12_U163 (.ZN( us12_n696 ) , .A1( us12_n830 ) , .B2( us12_n843 ) , .A2( us12_n865 ) , .B1( us12_n868 ) );
  INV_X1 us12_U164 (.A( us12_n730 ) , .ZN( us12_n839 ) );
  NAND2_X1 us12_U165 (.A1( us12_n447 ) , .A2( us12_n465 ) , .ZN( us12_n749 ) );
  AOI221_X1 us12_U166 (.A( us12_n483 ) , .ZN( us12_n488 ) , .B1( us12_n831 ) , .C2( us12_n844 ) , .C1( us12_n852 ) , .B2( us12_n862 ) );
  OAI22_X1 us12_U167 (.ZN( us12_n483 ) , .A1( us12_n708 ) , .B2( us12_n785 ) , .A2( us12_n806 ) , .B1( us12_n812 ) );
  INV_X1 us12_U168 (.A( us12_n790 ) , .ZN( us12_n832 ) );
  NAND2_X1 us12_U169 (.A1( us12_n451 ) , .A2( us12_n453 ) , .ZN( us12_n762 ) );
  NOR4_X1 us12_U17 (.A4( us12_n445 ) , .A3( us12_n446 ) , .A2( us12_n516 ) , .A1( us12_n541 ) , .ZN( us12_n706 ) );
  AOI211_X1 us12_U170 (.A( us12_n637 ) , .ZN( us12_n645 ) , .B( us12_n743 ) , .C2( us12_n839 ) , .C1( us12_n854 ) );
  OAI22_X1 us12_U171 (.ZN( us12_n637 ) , .A1( us12_n699 ) , .B2( us12_n728 ) , .A2( us12_n762 ) , .B1( us12_n816 ) );
  INV_X1 us12_U172 (.A( us12_n786 ) , .ZN( us12_n862 ) );
  OAI22_X1 us12_U173 (.B2( us12_n779 ) , .B1( us12_n780 ) , .ZN( us12_n781 ) , .A2( us12_n814 ) , .A1( us12_n815 ) );
  OAI22_X1 us12_U174 (.ZN( us12_n489 ) , .A1( us12_n724 ) , .B2( us12_n728 ) , .B1( us12_n730 ) , .A2( us12_n779 ) );
  INV_X1 us12_U175 (.A( us12_n788 ) , .ZN( us12_n845 ) );
  INV_X1 us12_U176 (.A( us12_n816 ) , .ZN( us12_n831 ) );
  OAI22_X1 us12_U177 (.A1( us12_n724 ) , .ZN( us12_n726 ) , .B2( us12_n750 ) , .B1( us12_n812 ) , .A2( us12_n816 ) );
  OAI22_X1 us12_U178 (.B2( us12_n803 ) , .B1( us12_n804 ) , .A2( us12_n805 ) , .A1( us12_n806 ) , .ZN( us12_n808 ) );
  OAI22_X1 us12_U179 (.ZN( us12_n496 ) , .A2( us12_n744 ) , .A1( us12_n780 ) , .B1( us12_n791 ) , .B2( us12_n806 ) );
  OR3_X1 us12_U18 (.ZN( us12_n446 ) , .A1( us12_n528 ) , .A3( us12_n577 ) , .A2( us12_n875 ) );
  INV_X1 us12_U180 (.A( us12_n814 ) , .ZN( us12_n833 ) );
  INV_X1 us12_U181 (.A( us12_n805 ) , .ZN( us12_n860 ) );
  OAI22_X1 us12_U182 (.ZN( us12_n710 ) , .A2( us12_n728 ) , .B2( us12_n729 ) , .A1( us12_n744 ) , .B1( us12_n813 ) );
  INV_X1 us12_U183 (.A( us12_n750 ) , .ZN( us12_n842 ) );
  OAI22_X1 us12_U184 (.B1( us12_n490 ) , .ZN( us12_n491 ) , .A1( us12_n686 ) , .A2( us12_n763 ) , .B2( us12_n817 ) );
  NOR3_X1 us12_U185 (.ZN( us12_n490 ) , .A1( us12_n782 ) , .A2( us12_n850 ) , .A3( us12_n863 ) );
  OAI22_X1 us12_U186 (.ZN( us12_n695 ) , .A2( us12_n730 ) , .A1( us12_n780 ) , .B1( us12_n791 ) , .B2( us12_n817 ) );
  OAI22_X1 us12_U187 (.B2( us12_n744 ) , .ZN( us12_n746 ) , .A2( us12_n762 ) , .B1( us12_n780 ) , .A1( us12_n792 ) );
  NOR2_X1 us12_U188 (.ZN( us12_n532 ) , .A2( us12_n749 ) , .A1( us12_n750 ) );
  INV_X1 us12_U189 (.A( us12_n744 ) , .ZN( us12_n837 ) );
  OR4_X1 us12_U19 (.A4( us12_n442 ) , .A2( us12_n443 ) , .A1( us12_n444 ) , .ZN( us12_n445 ) , .A3( us12_n553 ) );
  NOR2_X1 us12_U190 (.ZN( us12_n666 ) , .A1( us12_n728 ) , .A2( us12_n803 ) );
  NOR2_X1 us12_U191 (.ZN( us12_n615 ) , .A1( us12_n785 ) , .A2( us12_n815 ) );
  NOR2_X1 us12_U192 (.ZN( us12_n629 ) , .A2( us12_n728 ) , .A1( us12_n785 ) );
  NOR2_X1 us12_U193 (.ZN( us12_n715 ) , .A1( us12_n805 ) , .A2( us12_n817 ) );
  NOR2_X1 us12_U194 (.ZN( us12_n570 ) , .A1( us12_n728 ) , .A2( us12_n806 ) );
  NOR2_X1 us12_U195 (.A2( us12_n708 ) , .A1( us12_n750 ) , .ZN( us12_n771 ) );
  NOR2_X1 us12_U196 (.ZN( us12_n611 ) , .A2( us12_n780 ) , .A1( us12_n806 ) );
  NOR2_X1 us12_U197 (.ZN( us12_n601 ) , .A2( us12_n780 ) , .A1( us12_n803 ) );
  NOR2_X1 us12_U198 (.ZN( us12_n667 ) , .A1( us12_n750 ) , .A2( us12_n815 ) );
  NOR2_X1 us12_U199 (.ZN( us12_n555 ) , .A1( us12_n750 ) , .A2( us12_n791 ) );
  INV_X1 us12_U20 (.A( us12_n613 ) , .ZN( us12_n875 ) );
  NOR2_X1 us12_U200 (.ZN( us12_n654 ) , .A1( us12_n728 ) , .A2( us12_n813 ) );
  NOR2_X1 us12_U201 (.ZN( us12_n528 ) , .A2( us12_n724 ) , .A1( us12_n803 ) );
  NOR2_X1 us12_U202 (.ZN( us12_n546 ) , .A2( us12_n780 ) , .A1( us12_n814 ) );
  NOR2_X1 us12_U203 (.ZN( us12_n577 ) , .A2( us12_n699 ) , .A1( us12_n814 ) );
  NOR2_X1 us12_U204 (.ZN( us12_n508 ) , .A2( us12_n780 ) , .A1( us12_n785 ) );
  NOR2_X1 us12_U205 (.ZN( us12_n543 ) , .A2( us12_n708 ) , .A1( us12_n785 ) );
  NOR2_X1 us12_U206 (.ZN( us12_n664 ) , .A1( us12_n785 ) , .A2( us12_n791 ) );
  NOR2_X1 us12_U207 (.A2( us12_n744 ) , .ZN( us12_n755 ) , .A1( us12_n805 ) );
  NOR2_X1 us12_U208 (.ZN( us12_n735 ) , .A2( us12_n803 ) , .A1( us12_n805 ) );
  INV_X1 us12_U209 (.A( us12_n792 ) , .ZN( us12_n851 ) );
  INV_X1 us12_U21 (.A( us12_n749 ) , .ZN( us12_n863 ) );
  INV_X1 us12_U210 (.A( us12_n728 ) , .ZN( us12_n852 ) );
  NOR2_X1 us12_U211 (.A2( us12_n744 ) , .ZN( us12_n769 ) , .A1( us12_n812 ) );
  INV_X1 us12_U212 (.A( us12_n747 ) , .ZN( us12_n834 ) );
  NOR2_X1 us12_U213 (.A1( us12_n699 ) , .ZN( us12_n768 ) , .A2( us12_n813 ) );
  INV_X1 us12_U214 (.A( us12_n806 ) , .ZN( us12_n841 ) );
  NOR2_X1 us12_U215 (.ZN( us12_n531 ) , .A2( us12_n780 ) , .A1( us12_n816 ) );
  NOR2_X1 us12_U216 (.ZN( us12_n509 ) , .A1( us12_n729 ) , .A2( us12_n779 ) );
  NOR2_X1 us12_U217 (.ZN( us12_n599 ) , .A2( us12_n791 ) , .A1( us12_n816 ) );
  NOR2_X1 us12_U218 (.ZN( us12_n661 ) , .A1( us12_n729 ) , .A2( us12_n790 ) );
  NOR2_X1 us12_U219 (.ZN( us12_n507 ) , .A1( us12_n812 ) , .A2( us12_n817 ) );
  AOI222_X1 us12_U22 (.ZN( us12_n605 ) , .B2( us12_n671 ) , .B1( us12_n753 ) , .C2( us12_n831 ) , .A1( us12_n833 ) , .A2( us12_n862 ) , .C1( us12_n863 ) );
  NOR2_X1 us12_U220 (.ZN( us12_n544 ) , .A2( us12_n785 ) , .A1( us12_n792 ) );
  NOR2_X1 us12_U221 (.A1( us12_n749 ) , .ZN( us12_n767 ) , .A2( us12_n803 ) );
  NOR2_X1 us12_U222 (.ZN( us12_n545 ) , .A1( us12_n749 ) , .A2( us12_n814 ) );
  NOR2_X1 us12_U223 (.ZN( us12_n557 ) , .A1( us12_n792 ) , .A2( us12_n814 ) );
  NOR2_X1 us12_U224 (.ZN( us12_n556 ) , .A1( us12_n762 ) , .A2( us12_n805 ) );
  NOR2_X1 us12_U225 (.ZN( us12_n609 ) , .A2( us12_n724 ) , .A1( us12_n817 ) );
  NOR2_X1 us12_U226 (.ZN( us12_n663 ) , .A1( us12_n729 ) , .A2( us12_n785 ) );
  NOR2_X1 us12_U227 (.ZN( us12_n517 ) , .A1( us12_n708 ) , .A2( us12_n803 ) );
  NOR2_X1 us12_U228 (.ZN( us12_n506 ) , .A2( us12_n728 ) , .A1( us12_n762 ) );
  OAI22_X1 us12_U229 (.B1( us12_n440 ) , .ZN( us12_n444 ) , .A2( us12_n728 ) , .A1( us12_n744 ) , .B2( us12_n749 ) );
  AOI222_X1 us12_U23 (.ZN( us12_n563 ) , .B1( us12_n830 ) , .C1( us12_n841 ) , .A2( us12_n843 ) , .A1( us12_n854 ) , .B2( us12_n863 ) , .C2( us12_n873 ) );
  NOR3_X1 us12_U230 (.ZN( us12_n440 ) , .A2( us12_n836 ) , .A3( us12_n837 ) , .A1( us12_n846 ) );
  NOR2_X1 us12_U231 (.ZN( us12_n614 ) , .A1( us12_n762 ) , .A2( us12_n812 ) );
  NOR2_X1 us12_U232 (.ZN( us12_n533 ) , .A2( us12_n724 ) , .A1( us12_n730 ) );
  NOR2_X1 us12_U233 (.ZN( us12_n579 ) , .A2( us12_n708 ) , .A1( us12_n730 ) );
  NOR2_X1 us12_U234 (.ZN( us12_n521 ) , .A1( us12_n790 ) , .A2( us12_n812 ) );
  NOR2_X1 us12_U235 (.ZN( us12_n558 ) , .A1( us12_n708 ) , .A2( us12_n816 ) );
  NOR2_X1 us12_U236 (.ZN( us12_n655 ) , .A1( us12_n790 ) , .A2( us12_n815 ) );
  NOR2_X1 us12_U237 (.ZN( us12_n670 ) , .A1( us12_n790 ) , .A2( us12_n805 ) );
  NOR2_X1 us12_U238 (.ZN( us12_n668 ) , .A2( us12_n708 ) , .A1( us12_n790 ) );
  NOR2_X1 us12_U239 (.ZN( us12_n530 ) , .A2( us12_n744 ) , .A1( us12_n792 ) );
  AOI222_X1 us12_U24 (.ZN( us12_n660 ) , .A2( us12_n839 ) , .B1( us12_n841 ) , .C2( us12_n845 ) , .A1( us12_n860 ) , .C1( us12_n863 ) , .B2( us12_n870 ) );
  NOR2_X1 us12_U240 (.ZN( us12_n631 ) , .A1( us12_n724 ) , .A2( us12_n813 ) );
  NOR2_X1 us12_U241 (.ZN( us12_n630 ) , .A1( us12_n747 ) , .A2( us12_n815 ) );
  NOR2_X1 us12_U242 (.ZN( us12_n542 ) , .A1( us12_n762 ) , .A2( us12_n791 ) );
  INV_X1 us12_U243 (.A( us12_n763 ) , .ZN( us12_n866 ) );
  AOI21_X1 us12_U244 (.ZN( us12_n515 ) , .A( us12_n729 ) , .B1( us12_n750 ) , .B2( us12_n803 ) );
  NOR2_X1 us12_U245 (.ZN( us12_n718 ) , .A2( us12_n724 ) , .A1( us12_n744 ) );
  NOR2_X1 us12_U246 (.ZN( us12_n516 ) , .A1( us12_n708 ) , .A2( us12_n744 ) );
  INV_X1 us12_U247 (.A( us12_n729 ) , .ZN( us12_n868 ) );
  NOR2_X1 us12_U248 (.ZN( us12_n656 ) , .A1( us12_n747 ) , .A2( us12_n780 ) );
  AOI21_X1 us12_U249 (.ZN( us12_n540 ) , .A( us12_n763 ) , .B2( us12_n779 ) , .B1( us12_n817 ) );
  INV_X1 us12_U25 (.A( us12_n647 ) , .ZN( us12_n870 ) );
  NOR2_X1 us12_U250 (.ZN( us12_n559 ) , .A2( us12_n791 ) , .A1( us12_n803 ) );
  NOR2_X1 us12_U251 (.A2( us12_n708 ) , .A1( us12_n762 ) , .ZN( us12_n794 ) );
  NOR2_X1 us12_U252 (.ZN( us12_n642 ) , .A2( us12_n788 ) , .A1( us12_n791 ) );
  NOR2_X1 us12_U253 (.ZN( us12_n683 ) , .A2( us12_n699 ) , .A1( us12_n803 ) );
  AOI21_X1 us12_U254 (.B1( us12_n625 ) , .ZN( us12_n627 ) , .A( us12_n763 ) , .B2( us12_n814 ) );
  AOI21_X1 us12_U255 (.A( us12_n815 ) , .B2( us12_n816 ) , .B1( us12_n817 ) , .ZN( us12_n818 ) );
  AOI21_X1 us12_U256 (.ZN( us12_n650 ) , .A( us12_n779 ) , .B1( us12_n792 ) , .B2( us12_n805 ) );
  AOI21_X1 us12_U257 (.ZN( us12_n499 ) , .B1( us12_n680 ) , .A( us12_n812 ) , .B2( us12_n816 ) );
  NOR2_X1 us12_U258 (.ZN( us12_n520 ) , .A2( us12_n708 ) , .A1( us12_n814 ) );
  AOI21_X1 us12_U259 (.ZN( us12_n569 ) , .B1( us12_n750 ) , .B2( us12_n762 ) , .A( us12_n780 ) );
  NOR4_X1 us12_U26 (.ZN( us12_n473 ) , .A2( us12_n521 ) , .A4( us12_n594 ) , .A1( us12_n609 ) , .A3( us12_n629 ) );
  OAI221_X1 us12_U260 (.A( us12_n727 ) , .C2( us12_n728 ) , .B2( us12_n729 ) , .B1( us12_n730 ) , .ZN( us12_n737 ) , .C1( us12_n817 ) );
  AOI22_X1 us12_U261 (.ZN( us12_n727 ) , .B1( us12_n832 ) , .A2( us12_n838 ) , .A1( us12_n863 ) , .B2( us12_n866 ) );
  AOI21_X1 us12_U262 (.ZN( us12_n589 ) , .B2( us12_n699 ) , .B1( us12_n815 ) , .A( us12_n817 ) );
  NOR2_X1 us12_U263 (.ZN( us12_n519 ) , .A2( us12_n699 ) , .A1( us12_n816 ) );
  AOI21_X1 us12_U264 (.ZN( us12_n539 ) , .B2( us12_n812 ) , .A( us12_n814 ) , .B1( us12_n815 ) );
  AOI21_X1 us12_U265 (.ZN( us12_n640 ) , .B2( us12_n747 ) , .A( us12_n792 ) , .B1( us12_n803 ) );
  AOI21_X1 us12_U266 (.ZN( us12_n514 ) , .A( us12_n779 ) , .B2( us12_n792 ) , .B1( us12_n812 ) );
  AOI21_X1 us12_U267 (.B1( us12_n699 ) , .ZN( us12_n700 ) , .A( us12_n732 ) , .B2( us12_n763 ) );
  AOI21_X1 us12_U268 (.ZN( us12_n591 ) , .B2( us12_n763 ) , .A( us12_n785 ) , .B1( us12_n812 ) );
  AOI21_X1 us12_U269 (.ZN( us12_n593 ) , .B1( us12_n750 ) , .A( us12_n792 ) , .B2( us12_n813 ) );
  NOR4_X1 us12_U27 (.A4( us12_n544 ) , .A3( us12_n545 ) , .A2( us12_n546 ) , .A1( us12_n547 ) , .ZN( us12_n548 ) );
  NOR2_X1 us12_U270 (.ZN( us12_n547 ) , .A1( us12_n699 ) , .A2( us12_n744 ) );
  INV_X1 us12_U271 (.A( us12_n791 ) , .ZN( us12_n873 ) );
  AOI21_X1 us12_U272 (.ZN( us12_n564 ) , .B1( us12_n724 ) , .A( us12_n779 ) , .B2( us12_n791 ) );
  AOI21_X1 us12_U273 (.ZN( us12_n497 ) , .A( us12_n779 ) , .B2( us12_n791 ) , .B1( us12_n804 ) );
  AOI21_X1 us12_U274 (.ZN( us12_n498 ) , .A( us12_n724 ) , .B2( us12_n762 ) , .B1( us12_n814 ) );
  AOI21_X1 us12_U275 (.ZN( us12_n649 ) , .B1( us12_n729 ) , .B2( us12_n763 ) , .A( us12_n813 ) );
  NOR2_X1 us12_U276 (.ZN( us12_n529 ) , .A1( us12_n708 ) , .A2( us12_n779 ) );
  NOR2_X1 us12_U277 (.ZN( us12_n685 ) , .A1( us12_n729 ) , .A2( us12_n816 ) );
  AOI21_X1 us12_U278 (.B1( us12_n686 ) , .ZN( us12_n687 ) , .A( us12_n728 ) , .B2( us12_n761 ) );
  AOI21_X1 us12_U279 (.A( us12_n812 ) , .B2( us12_n813 ) , .B1( us12_n814 ) , .ZN( us12_n819 ) );
  NOR4_X1 us12_U28 (.A4( us12_n532 ) , .A3( us12_n533 ) , .A2( us12_n534 ) , .ZN( us12_n535 ) , .A1( us12_n820 ) );
  AOI21_X1 us12_U280 (.ZN( us12_n450 ) , .B2( us12_n792 ) , .A( us12_n803 ) , .B1( us12_n815 ) );
  NOR2_X1 us12_U281 (.ZN( us12_n568 ) , .A1( us12_n729 ) , .A2( us12_n762 ) );
  NOR2_X1 us12_U282 (.ZN( us12_n682 ) , .A2( us12_n708 ) , .A1( us12_n817 ) );
  AOI21_X1 us12_U283 (.ZN( us12_n641 ) , .B1( us12_n680 ) , .A( us12_n791 ) , .B2( us12_n817 ) );
  INV_X1 us12_U284 (.A( us12_n699 ) , .ZN( us12_n853 ) );
  AOI21_X1 us12_U285 (.ZN( us12_n689 ) , .B2( us12_n749 ) , .B1( us12_n763 ) , .A( us12_n806 ) );
  AOI21_X1 us12_U286 (.ZN( us12_n639 ) , .B2( us12_n749 ) , .A( us12_n788 ) , .B1( us12_n812 ) );
  AOI21_X1 us12_U287 (.A( us12_n790 ) , .B2( us12_n791 ) , .B1( us12_n792 ) , .ZN( us12_n793 ) );
  AOI21_X1 us12_U288 (.A( us12_n733 ) , .ZN( us12_n734 ) , .B2( us12_n780 ) , .B1( us12_n792 ) );
  NOR2_X1 us12_U289 (.ZN( us12_n567 ) , .A1( us12_n747 ) , .A2( us12_n805 ) );
  NOR4_X1 us12_U29 (.ZN( us12_n479 ) , .A1( us12_n520 ) , .A4( us12_n557 ) , .A3( us12_n582 ) , .A2( us12_n630 ) );
  NAND2_X1 us12_U290 (.ZN( us12_n753 ) , .A1( us12_n763 ) , .A2( us12_n805 ) );
  NOR2_X1 us12_U291 (.A2( us12_n813 ) , .A1( us12_n815 ) , .ZN( us12_n821 ) );
  NOR2_X1 us12_U292 (.ZN( us12_n578 ) , .A1( us12_n708 ) , .A2( us12_n813 ) );
  NOR2_X1 us12_U293 (.ZN( us12_n665 ) , .A1( us12_n780 ) , .A2( us12_n813 ) );
  NOR2_X1 us12_U294 (.ZN( us12_n711 ) , .A1( us12_n762 ) , .A2( us12_n763 ) );
  NOR2_X1 us12_U295 (.ZN( us12_n583 ) , .A1( us12_n792 ) , .A2( us12_n817 ) );
  AOI21_X1 us12_U296 (.ZN( us12_n442 ) , .A( us12_n699 ) , .B1( us12_n733 ) , .B2( us12_n750 ) );
  NOR2_X1 us12_U297 (.ZN( us12_n534 ) , .A1( us12_n724 ) , .A2( us12_n788 ) );
  NOR2_X1 us12_U298 (.ZN( us12_n582 ) , .A1( us12_n744 ) , .A2( us12_n815 ) );
  NOR2_X1 us12_U299 (.ZN( us12_n684 ) , .A1( us12_n791 ) , .A2( us12_n813 ) );
  NAND2_X1 us12_U3 (.A1( us12_n449 ) , .A2( us12_n460 ) , .ZN( us12_n792 ) );
  NOR4_X1 us12_U30 (.ZN( us12_n456 ) , .A2( us12_n517 ) , .A1( us12_n543 ) , .A3( us12_n579 ) , .A4( us12_n615 ) );
  OAI21_X1 us12_U300 (.A( us12_n698 ) , .ZN( us12_n702 ) , .B2( us12_n750 ) , .B1( us12_n804 ) );
  OAI21_X1 us12_U301 (.ZN( us12_n698 ) , .B2( us12_n833 ) , .B1( us12_n838 ) , .A( us12_n860 ) );
  INV_X1 us12_U302 (.A( us12_n815 ) , .ZN( us12_n855 ) );
  INV_X1 us12_U303 (.A( us12_n785 ) , .ZN( us12_n846 ) );
  OAI21_X1 us12_U304 (.A( us12_n731 ) , .B1( us12_n732 ) , .ZN( us12_n736 ) , .B2( us12_n805 ) );
  OAI21_X1 us12_U305 (.ZN( us12_n731 ) , .A( us12_n833 ) , .B2( us12_n852 ) , .B1( us12_n873 ) );
  INV_X1 us12_U306 (.A( us12_n780 ) , .ZN( us12_n850 ) );
  INV_X1 us12_U307 (.A( us12_n813 ) , .ZN( us12_n836 ) );
  OAI221_X1 us12_U308 (.A( us12_n783 ) , .C2( us12_n784 ) , .B2( us12_n785 ) , .B1( us12_n786 ) , .ZN( us12_n796 ) , .C1( us12_n813 ) );
  AOI22_X1 us12_U309 (.A2( us12_n782 ) , .ZN( us12_n783 ) , .B2( us12_n831 ) , .A1( us12_n834 ) , .B1( us12_n863 ) );
  AOI221_X1 us12_U31 (.A( us12_n713 ) , .B2( us12_n714 ) , .ZN( us12_n720 ) , .C1( us12_n832 ) , .B1( us12_n839 ) , .C2( us12_n863 ) );
  OAI21_X1 us12_U310 (.A( us12_n787 ) , .B2( us12_n788 ) , .B1( us12_n789 ) , .ZN( us12_n795 ) );
  OAI21_X1 us12_U311 (.ZN( us12_n787 ) , .A( us12_n839 ) , .B1( us12_n863 ) , .B2( us12_n873 ) );
  NAND2_X1 us12_U312 (.A2( us12_n762 ) , .A1( us12_n806 ) , .ZN( us12_n810 ) );
  NOR2_X1 us12_U313 (.ZN( us12_n470 ) , .A2( us12_n779 ) , .A1( us12_n815 ) );
  NOR2_X1 us12_U314 (.ZN( us12_n484 ) , .A1( us12_n788 ) , .A2( us12_n805 ) );
  NAND2_X1 us12_U315 (.ZN( us12_n714 ) , .A1( us12_n728 ) , .A2( us12_n780 ) );
  NAND2_X1 us12_U316 (.ZN( us12_n671 ) , .A1( us12_n806 ) , .A2( us12_n816 ) );
  NOR2_X1 us12_U317 (.ZN( us12_n526 ) , .A1( us12_n724 ) , .A2( us12_n750 ) );
  AOI21_X1 us12_U318 (.ZN( us12_n443 ) , .B1( us12_n789 ) , .B2( us12_n791 ) , .A( us12_n814 ) );
  INV_X1 us12_U319 (.A( us12_n817 ) , .ZN( us12_n844 ) );
  OR2_X1 us12_U32 (.A2( us12_n711 ) , .A1( us12_n712 ) , .ZN( us12_n713 ) );
  NOR2_X1 us12_U320 (.ZN( us12_n712 ) , .A2( us12_n724 ) , .A1( us12_n790 ) );
  NAND2_X1 us12_U321 (.A1( us12_n699 ) , .A2( us12_n729 ) , .ZN( us12_n782 ) );
  NOR2_X1 us12_U322 (.ZN( us12_n518 ) , .A1( us12_n708 ) , .A2( us12_n788 ) );
  OAI22_X1 us12_U323 (.B2( us12_n750 ) , .B1( us12_n751 ) , .A1( us12_n752 ) , .ZN( us12_n756 ) , .A2( us12_n806 ) );
  NOR3_X1 us12_U324 (.ZN( us12_n752 ) , .A2( us12_n853 ) , .A1( us12_n863 ) , .A3( us12_n865 ) );
  NOR2_X1 us12_U325 (.ZN( us12_n751 ) , .A2( us12_n852 ) , .A1( us12_n860 ) );
  INV_X1 us12_U326 (.A( us12_n724 ) , .ZN( us12_n856 ) );
  NAND2_X2 us12_U327 (.A2( us12_n454 ) , .A1( us12_n472 ) , .ZN( us12_n779 ) );
  AND2_X1 us12_U328 (.ZN( us12_n732 ) , .A1( us12_n779 ) , .A2( us12_n785 ) );
  AOI221_X1 us12_U329 (.A( us12_n764 ) , .ZN( us12_n774 ) , .C2( us12_n810 ) , .B2( us12_n835 ) , .C1( us12_n855 ) , .B1( us12_n866 ) );
  NOR2_X1 us12_U33 (.ZN( us12_n680 ) , .A2( us12_n834 ) , .A1( us12_n839 ) );
  AOI21_X1 us12_U330 (.B2( us12_n763 ) , .ZN( us12_n764 ) , .A( us12_n788 ) , .B1( us12_n792 ) );
  INV_X1 us12_U331 (.A( us12_n761 ) , .ZN( us12_n835 ) );
  NAND2_X1 us12_U332 (.A2( us12_n448 ) , .A1( us12_n460 ) , .ZN( us12_n728 ) );
  NAND2_X1 us12_U333 (.A1( us12_n451 ) , .A2( us12_n454 ) , .ZN( us12_n814 ) );
  NAND2_X1 us12_U334 (.A1( us12_n447 ) , .A2( us12_n449 ) , .ZN( us12_n805 ) );
  NAND2_X1 us12_U335 (.A1( us12_n451 ) , .A2( us12_n471 ) , .ZN( us12_n816 ) );
  NAND2_X1 us12_U336 (.A2( us12_n453 ) , .A1( us12_n455 ) , .ZN( us12_n806 ) );
  NAND2_X1 us12_U337 (.A2( us12_n464 ) , .A1( us12_n465 ) , .ZN( us12_n812 ) );
  NAND2_X1 us12_U338 (.A1( us12_n441 ) , .A2( us12_n460 ) , .ZN( us12_n699 ) );
  NAND2_X1 us12_U339 (.A2( us12_n449 ) , .A1( us12_n452 ) , .ZN( us12_n763 ) );
  AOI222_X1 us12_U34 (.ZN( us12_n469 ) , .B1( us12_n832 ) , .A1( us12_n839 ) , .C1( us12_n842 ) , .C2( us12_n851 ) , .A2( us12_n855 ) , .B2( us12_n865 ) );
  NAND2_X2 us12_U340 (.A1( us12_n455 ) , .A2( us12_n462 ) , .ZN( us12_n750 ) );
  NAND2_X1 us12_U341 (.A2( us12_n448 ) , .A1( us12_n452 ) , .ZN( us12_n729 ) );
  NOR2_X1 us12_U342 (.ZN( us12_n453 ) , .A1( us12_n826 ) , .A2( us12_n827 ) );
  NOR2_X1 us12_U343 (.ZN( us12_n465 ) , .A2( us12_n847 ) , .A1( us12_n848 ) );
  NOR2_X1 us12_U344 (.ZN( us12_n451 ) , .A1( us12_n828 ) , .A2( us12_n829 ) );
  NAND2_X1 us12_U345 (.A1( us12_n462 ) , .A2( us12_n472 ) , .ZN( us12_n788 ) );
  NAND2_X1 us12_U346 (.A2( us12_n461 ) , .A1( us12_n471 ) , .ZN( us12_n697 ) );
  NAND2_X1 us12_U347 (.A2( us12_n461 ) , .A1( us12_n462 ) , .ZN( us12_n747 ) );
  NAND2_X1 us12_U348 (.A1( us12_n451 ) , .A2( us12_n462 ) , .ZN( us12_n790 ) );
  NAND2_X1 us12_U349 (.A1( us12_n452 ) , .A2( us12_n465 ) , .ZN( us12_n669 ) );
  NOR4_X1 us12_U35 (.A1( us12_n466 ) , .ZN( us12_n467 ) , .A4( us12_n542 ) , .A2( us12_n554 ) , .A3( us12_n614 ) );
  NAND2_X1 us12_U350 (.A2( us12_n441 ) , .A1( us12_n447 ) , .ZN( us12_n784 ) );
  NAND2_X2 us12_U351 (.A1( us12_n441 ) , .A2( us12_n464 ) , .ZN( us12_n708 ) );
  NAND2_X1 us12_U352 (.A2( us12_n471 ) , .A1( us12_n472 ) , .ZN( us12_n817 ) );
  NAND2_X1 us12_U353 (.A2( us12_n454 ) , .A1( us12_n455 ) , .ZN( us12_n730 ) );
  NOR2_X1 us12_U354 (.ZN( us12_n447 ) , .A2( us12_n849 ) , .A1( us12_n858 ) );
  NAND2_X1 us12_U355 (.A1( us12_n447 ) , .A2( us12_n448 ) , .ZN( us12_n786 ) );
  NAND2_X1 us12_U356 (.A1( us12_n454 ) , .A2( us12_n461 ) , .ZN( us12_n813 ) );
  NAND2_X2 us12_U357 (.A1( us12_n453 ) , .A2( us12_n472 ) , .ZN( us12_n785 ) );
  NAND2_X1 us12_U358 (.A1( us12_n453 ) , .A2( us12_n461 ) , .ZN( us12_n744 ) );
  NOR2_X1 us12_U359 (.A2( sa12_6 ) , .A1( sa12_7 ) , .ZN( us12_n464 ) );
  AOI221_X1 us12_U36 (.ZN( us12_n468 ) , .C2( us12_n714 ) , .B2( us12_n831 ) , .C1( us12_n845 ) , .B1( us12_n860 ) , .A( us12_n864 ) );
  NOR2_X1 us12_U360 (.A2( sa12_2 ) , .ZN( us12_n461 ) , .A1( us12_n829 ) );
  NOR2_X1 us12_U361 (.A2( sa12_7 ) , .ZN( us12_n460 ) , .A1( us12_n849 ) );
  NOR2_X1 us12_U362 (.A2( sa12_4 ) , .ZN( us12_n449 ) , .A1( us12_n848 ) );
  NOR2_X1 us12_U363 (.A2( sa12_4 ) , .A1( sa12_5 ) , .ZN( us12_n441 ) );
  NOR2_X1 us12_U364 (.A2( sa12_5 ) , .ZN( us12_n448 ) , .A1( us12_n847 ) );
  NOR2_X1 us12_U365 (.A2( sa12_0 ) , .ZN( us12_n454 ) , .A1( us12_n827 ) );
  NOR2_X1 us12_U366 (.A2( sa12_1 ) , .ZN( us12_n471 ) , .A1( us12_n826 ) );
  NOR2_X1 us12_U367 (.A2( sa12_6 ) , .ZN( us12_n452 ) , .A1( us12_n858 ) );
  NOR2_X1 us12_U368 (.A2( sa12_0 ) , .A1( sa12_1 ) , .ZN( us12_n462 ) );
  INV_X1 us12_U369 (.A( sa12_6 ) , .ZN( us12_n849 ) );
  NOR4_X1 us12_U37 (.A4( us12_n577 ) , .A3( us12_n578 ) , .A2( us12_n579 ) , .ZN( us12_n586 ) , .A1( us12_n683 ) );
  INV_X1 us12_U370 (.A( sa12_4 ) , .ZN( us12_n847 ) );
  INV_X1 us12_U371 (.A( sa12_1 ) , .ZN( us12_n827 ) );
  NAND2_X2 us12_U372 (.A1( us12_n455 ) , .A2( us12_n471 ) , .ZN( us12_n803 ) );
  INV_X1 us12_U373 (.A( sa12_0 ) , .ZN( us12_n826 ) );
  INV_X1 us12_U374 (.A( sa12_7 ) , .ZN( us12_n858 ) );
  INV_X1 us12_U375 (.A( sa12_5 ) , .ZN( us12_n848 ) );
  INV_X1 us12_U376 (.A( sa12_2 ) , .ZN( us12_n828 ) );
  AOI21_X1 us12_U377 (.ZN( us12_n510 ) , .B2( us12_n669 ) , .A( us12_n730 ) , .B1( us12_n815 ) );
  OAI22_X1 us12_U378 (.ZN( us12_n624 ) , .B1( us12_n669 ) , .B2( us12_n747 ) , .A1( us12_n815 ) , .A2( us12_n816 ) );
  AOI21_X1 us12_U379 (.ZN( us12_n626 ) , .B2( us12_n669 ) , .A( us12_n790 ) , .B1( us12_n791 ) );
  NOR4_X1 us12_U38 (.A1( us12_n584 ) , .ZN( us12_n585 ) , .A3( us12_n652 ) , .A2( us12_n662 ) , .A4( us12_n767 ) );
  INV_X1 us12_U380 (.A( us12_n669 ) , .ZN( us12_n865 ) );
  NOR2_X1 us12_U381 (.A1( us12_n669 ) , .ZN( us12_n766 ) , .A2( us12_n813 ) );
  AOI21_X1 us12_U382 (.ZN( us12_n477 ) , .A( us12_n669 ) , .B1( us12_n750 ) , .B2( us12_n806 ) );
  NOR2_X1 us12_U383 (.A1( us12_n669 ) , .ZN( us12_n673 ) , .A2( us12_n744 ) );
  NOR2_X1 us12_U384 (.ZN( us12_n602 ) , .A1( us12_n669 ) , .A2( us12_n803 ) );
  NOR2_X1 us12_U385 (.A1( us12_n669 ) , .ZN( us12_n688 ) , .A2( us12_n816 ) );
  NOR2_X1 us12_U386 (.ZN( us12_n527 ) , .A1( us12_n669 ) , .A2( us12_n779 ) );
  NOR2_X1 us12_U387 (.ZN( us12_n652 ) , .A1( us12_n669 ) , .A2( us12_n814 ) );
  NOR2_X1 us12_U388 (.ZN( us12_n628 ) , .A2( us12_n669 ) , .A1( us12_n785 ) );
  NOR2_X1 us12_U389 (.ZN( us12_n581 ) , .A1( us12_n669 ) , .A2( us12_n788 ) );
  NOR4_X1 us12_U39 (.A4( us12_n661 ) , .A3( us12_n662 ) , .A2( us12_n663 ) , .A1( us12_n664 ) , .ZN( us12_n677 ) );
  OAI22_X1 us12_U390 (.ZN( us12_n590 ) , .B1( us12_n730 ) , .B2( us12_n749 ) , .A2( us12_n786 ) , .A1( us12_n803 ) );
  NAND2_X1 us12_U391 (.A2( us12_n749 ) , .A1( us12_n786 ) , .ZN( us12_n809 ) );
  NOR2_X1 us12_U392 (.ZN( us12_n612 ) , .A1( us12_n779 ) , .A2( us12_n786 ) );
  NOR2_X1 us12_U393 (.ZN( us12_n717 ) , .A2( us12_n744 ) , .A1( us12_n786 ) );
  NOR2_X1 us12_U394 (.ZN( us12_n653 ) , .A1( us12_n762 ) , .A2( us12_n786 ) );
  NOR2_X1 us12_U395 (.ZN( us12_n554 ) , .A1( us12_n786 ) , .A2( us12_n813 ) );
  NOR2_X1 us12_U396 (.ZN( us12_n701 ) , .A2( us12_n786 ) , .A1( us12_n817 ) );
  OAI222_X1 us12_U397 (.ZN( us12_n617 ) , .B1( us12_n697 ) , .C1( us12_n724 ) , .C2( us12_n747 ) , .B2( us12_n786 ) , .A2( us12_n792 ) , .A1( us12_n816 ) );
  NOR2_X1 us12_U398 (.A1( us12_n730 ) , .ZN( us12_n765 ) , .A2( us12_n786 ) );
  NAND2_X1 us12_U399 (.A1( us12_n729 ) , .A2( us12_n784 ) , .ZN( us12_n811 ) );
  NAND2_X1 us12_U4 (.A1( us12_n449 ) , .A2( us12_n464 ) , .ZN( us12_n724 ) );
  NOR4_X1 us12_U40 (.A4( us12_n665 ) , .A3( us12_n666 ) , .A2( us12_n667 ) , .A1( us12_n668 ) , .ZN( us12_n676 ) );
  OAI22_X1 us12_U400 (.ZN( us12_n588 ) , .A2( us12_n747 ) , .B2( us12_n762 ) , .A1( us12_n763 ) , .B1( us12_n784 ) );
  OAI221_X1 us12_U401 (.A( us12_n696 ) , .ZN( us12_n703 ) , .C2( us12_n784 ) , .C1( us12_n785 ) , .B1( us12_n786 ) , .B2( us12_n806 ) );
  AOI21_X1 us12_U402 (.ZN( us12_n592 ) , .B1( us12_n728 ) , .B2( us12_n784 ) , .A( us12_n790 ) );
  AOI21_X1 us12_U403 (.ZN( us12_n648 ) , .A( us12_n762 ) , .B2( us12_n784 ) , .B1( us12_n792 ) );
  AOI21_X1 us12_U404 (.ZN( us12_n623 ) , .B1( us12_n699 ) , .A( us12_n779 ) , .B2( us12_n784 ) );
  OAI22_X1 us12_U405 (.ZN( us12_n681 ) , .A1( us12_n699 ) , .A2( us12_n730 ) , .B2( us12_n784 ) , .B1( us12_n817 ) );
  OAI21_X1 us12_U406 (.A( us12_n613 ) , .ZN( us12_n616 ) , .B1( us12_n625 ) , .B2( us12_n784 ) );
  NOR2_X1 us12_U407 (.ZN( us12_n610 ) , .A1( us12_n784 ) , .A2( us12_n816 ) );
  NOR2_X1 us12_U408 (.ZN( us12_n651 ) , .A1( us12_n784 ) , .A2( us12_n788 ) );
  OAI222_X1 us12_U409 (.A2( us12_n669 ) , .ZN( us12_n674 ) , .B1( us12_n747 ) , .B2( us12_n784 ) , .C2( us12_n788 ) , .C1( us12_n815 ) , .A1( us12_n817 ) );
  NOR4_X1 us12_U41 (.A3( us12_n673 ) , .A1( us12_n674 ) , .ZN( us12_n675 ) , .A4( us12_n715 ) , .A2( us12_n859 ) );
  NOR2_X1 us12_U410 (.ZN( us12_n553 ) , .A2( us12_n744 ) , .A1( us12_n784 ) );
  INV_X1 us12_U411 (.A( us12_n784 ) , .ZN( us12_n861 ) );
  AOI21_X1 us12_U412 (.ZN( us12_n500 ) , .A( us12_n697 ) , .B1( us12_n708 ) , .B2( us12_n786 ) );
  INV_X1 us12_U413 (.A( us12_n697 ) , .ZN( us12_n838 ) );
  NOR2_X1 us12_U414 (.A1( us12_n697 ) , .ZN( us12_n770 ) , .A2( us12_n815 ) );
  AOI21_X1 us12_U415 (.ZN( us12_n571 ) , .B2( us12_n697 ) , .B1( us12_n806 ) , .A( us12_n812 ) );
  NOR2_X1 us12_U416 (.ZN( us12_n632 ) , .A2( us12_n697 ) , .A1( us12_n724 ) );
  AOI21_X1 us12_U417 (.ZN( us12_n478 ) , .B2( us12_n697 ) , .A( us12_n749 ) , .B1( us12_n779 ) );
  NOR2_X1 us12_U418 (.A2( us12_n697 ) , .A1( us12_n780 ) , .ZN( us12_n820 ) );
  NOR2_X1 us12_U419 (.ZN( us12_n662 ) , .A2( us12_n697 ) , .A1( us12_n729 ) );
  AOI221_X1 us12_U42 (.A( us12_n781 ) , .ZN( us12_n798 ) , .C2( us12_n837 ) , .B2( us12_n838 ) , .B1( us12_n865 ) , .C1( us12_n866 ) );
  NOR2_X1 us12_U420 (.ZN( us12_n566 ) , .A2( us12_n697 ) , .A1( us12_n763 ) );
  NOR2_X1 us12_U421 (.ZN( us12_n600 ) , .A2( us12_n697 ) , .A1( us12_n784 ) );
  NOR2_X1 us12_U422 (.A2( us12_n697 ) , .ZN( us12_n716 ) , .A1( us12_n792 ) );
  NOR2_X1 us12_U423 (.ZN( us12_n594 ) , .A2( us12_n697 ) , .A1( us12_n728 ) );
  AOI21_X1 us12_U424 (.ZN( us12_n552 ) , .B1( us12_n669 ) , .A( us12_n697 ) , .B2( us12_n805 ) );
  NOR2_X1 us12_U425 (.ZN( us12_n541 ) , .A2( us12_n697 ) , .A1( us12_n699 ) );
  NOR2_X1 us12_U426 (.ZN( us12_n580 ) , .A2( us12_n697 ) , .A1( us12_n791 ) );
  NOR2_X1 us12_U427 (.A2( sa12_2 ) , .A1( sa12_3 ) , .ZN( us12_n472 ) );
  NOR2_X1 us12_U428 (.A2( sa12_3 ) , .ZN( us12_n455 ) , .A1( us12_n828 ) );
  INV_X1 us12_U429 (.A( sa12_3 ) , .ZN( us12_n829 ) );
  NOR4_X1 us12_U43 (.A4( us12_n793 ) , .A3( us12_n794 ) , .A2( us12_n795 ) , .A1( us12_n796 ) , .ZN( us12_n797 ) );
  OAI222_X1 us12_U430 (.ZN( us12_n505 ) , .C2( us12_n625 ) , .B2( us12_n647 ) , .B1( us12_n747 ) , .A2( us12_n748 ) , .C1( us12_n805 ) , .A1( us12_n806 ) );
  OAI222_X1 us12_U431 (.B2( us12_n747 ) , .B1( us12_n748 ) , .A2( us12_n749 ) , .ZN( us12_n757 ) , .C2( us12_n805 ) , .C1( us12_n814 ) , .A1( us12_n817 ) );
  NOR2_X1 us12_U432 (.ZN( us12_n748 ) , .A1( us12_n861 ) , .A2( us12_n862 ) );
  AND2_X1 us12_U433 (.ZN( us12_n438 ) , .A2( us12_n831 ) , .A1( us12_n854 ) );
  AND2_X1 us12_U434 (.ZN( us12_n439 ) , .A2( us12_n843 ) , .A1( us12_n861 ) );
  NOR3_X1 us12_U435 (.A1( us12_n438 ) , .A2( us12_n439 ) , .A3( us12_n576 ) , .ZN( us12_n587 ) );
  INV_X1 us12_U436 (.A( us12_n812 ) , .ZN( us12_n854 ) );
  NAND3_X1 us12_U437 (.ZN( sa11_sr_6 ) , .A3( us12_n797 ) , .A2( us12_n798 ) , .A1( us12_n799 ) );
  NAND3_X1 us12_U438 (.ZN( sa11_sr_5 ) , .A3( us12_n758 ) , .A2( us12_n759 ) , .A1( us12_n760 ) );
  NAND3_X1 us12_U439 (.ZN( sa11_sr_4 ) , .A3( us12_n738 ) , .A2( us12_n739 ) , .A1( us12_n740 ) );
  NOR4_X1 us12_U44 (.A4( us12_n776 ) , .A3( us12_n777 ) , .A1( us12_n778 ) , .ZN( us12_n799 ) , .A2( us12_n801 ) );
  NAND3_X1 us12_U440 (.A3( us12_n675 ) , .A2( us12_n676 ) , .A1( us12_n677 ) , .ZN( us12_n807 ) );
  NAND3_X1 us12_U441 (.ZN( us12_n638 ) , .A3( us12_n708 ) , .A2( us12_n724 ) , .A1( us12_n792 ) );
  NAND3_X1 us12_U442 (.A3( us12_n618 ) , .A2( us12_n619 ) , .A1( us12_n620 ) , .ZN( us12_n725 ) );
  NAND3_X1 us12_U443 (.A3( us12_n585 ) , .A2( us12_n586 ) , .A1( us12_n587 ) , .ZN( us12_n621 ) );
  NAND3_X1 us12_U444 (.ZN( us12_n565 ) , .A3( us12_n680 ) , .A2( us12_n750 ) , .A1( us12_n785 ) );
  NAND3_X1 us12_U445 (.A3( us12_n523 ) , .A2( us12_n524 ) , .A1( us12_n525 ) , .ZN( us12_n742 ) );
  NAND3_X1 us12_U446 (.A3( us12_n512 ) , .A1( us12_n513 ) , .ZN( us12_n608 ) , .A2( us12_n871 ) );
  NAND3_X1 us12_U447 (.A3( us12_n467 ) , .A2( us12_n468 ) , .A1( us12_n469 ) , .ZN( us12_n777 ) );
  INV_X1 us12_U448 (.A( us12_n803 ) , .ZN( us12_n843 ) );
  AOI21_X1 us12_U449 (.ZN( us12_n576 ) , .B2( us12_n724 ) , .B1( us12_n748 ) , .A( us12_n785 ) );
  NOR4_X1 us12_U45 (.A4( us12_n734 ) , .A3( us12_n735 ) , .A2( us12_n736 ) , .A1( us12_n737 ) , .ZN( us12_n738 ) );
  AOI211_X1 us12_U46 (.B( us12_n725 ) , .A( us12_n726 ) , .ZN( us12_n739 ) , .C1( us12_n843 ) , .C2( us12_n855 ) );
  NOR3_X1 us12_U47 (.A3( us12_n722 ) , .A1( us12_n723 ) , .ZN( us12_n740 ) , .A2( us12_n741 ) );
  NAND4_X1 us12_U48 (.ZN( sa11_sr_3 ) , .A4( us12_n704 ) , .A3( us12_n705 ) , .A2( us12_n706 ) , .A1( us12_n707 ) );
  NOR4_X1 us12_U49 (.A4( us12_n700 ) , .A3( us12_n701 ) , .A2( us12_n702 ) , .A1( us12_n703 ) , .ZN( us12_n704 ) );
  NAND2_X1 us12_U5 (.A2( us12_n448 ) , .A1( us12_n464 ) , .ZN( us12_n815 ) );
  AOI211_X1 us12_U50 (.B( us12_n694 ) , .A( us12_n695 ) , .ZN( us12_n705 ) , .C2( us12_n831 ) , .C1( us12_n851 ) );
  NOR2_X1 us12_U51 (.ZN( us12_n707 ) , .A2( us12_n776 ) , .A1( us12_n800 ) );
  NOR2_X1 us12_U52 (.ZN( us12_n804 ) , .A1( us12_n854 ) , .A2( us12_n861 ) );
  NAND4_X1 us12_U53 (.ZN( sa11_sr_0 ) , .A4( us12_n501 ) , .A3( us12_n502 ) , .A2( us12_n503 ) , .A1( us12_n504 ) );
  AOI221_X1 us12_U54 (.A( us12_n497 ) , .ZN( us12_n502 ) , .B2( us12_n843 ) , .C1( us12_n846 ) , .C2( us12_n860 ) , .B1( us12_n862 ) );
  NOR4_X1 us12_U55 (.A4( us12_n498 ) , .A3( us12_n499 ) , .A2( us12_n500 ) , .ZN( us12_n501 ) , .A1( us12_n527 ) );
  AOI211_X1 us12_U56 (.A( us12_n496 ) , .ZN( us12_n503 ) , .B( us12_n802 ) , .C2( us12_n839 ) , .C1( us12_n851 ) );
  NAND4_X1 us12_U57 (.ZN( sa11_sr_1 ) , .A4( us12_n595 ) , .A3( us12_n596 ) , .A2( us12_n597 ) , .A1( us12_n598 ) );
  AOI211_X1 us12_U58 (.B( us12_n589 ) , .A( us12_n590 ) , .ZN( us12_n596 ) , .C2( us12_n811 ) , .C1( us12_n833 ) );
  NOR4_X1 us12_U59 (.A4( us12_n591 ) , .A3( us12_n592 ) , .A2( us12_n593 ) , .A1( us12_n594 ) , .ZN( us12_n595 ) );
  NAND2_X1 us12_U6 (.A2( us12_n441 ) , .A1( us12_n452 ) , .ZN( us12_n791 ) );
  AOI211_X1 us12_U60 (.A( us12_n588 ) , .ZN( us12_n597 ) , .B( us12_n621 ) , .C1( us12_n845 ) , .C2( us12_n855 ) );
  NAND4_X1 us12_U61 (.ZN( sa11_sr_7 ) , .A4( us12_n822 ) , .A3( us12_n823 ) , .A2( us12_n824 ) , .A1( us12_n825 ) );
  NOR4_X1 us12_U62 (.A4( us12_n818 ) , .A3( us12_n819 ) , .A2( us12_n820 ) , .A1( us12_n821 ) , .ZN( us12_n822 ) );
  AOI222_X1 us12_U63 (.C2( us12_n809 ) , .B2( us12_n810 ) , .A2( us12_n811 ) , .ZN( us12_n823 ) , .C1( us12_n832 ) , .A1( us12_n839 ) , .B1( us12_n853 ) );
  AOI211_X1 us12_U64 (.B( us12_n807 ) , .A( us12_n808 ) , .ZN( us12_n824 ) , .C1( us12_n842 ) , .C2( us12_n850 ) );
  NAND4_X1 us12_U65 (.ZN( sa11_sr_2 ) , .A4( us12_n643 ) , .A3( us12_n644 ) , .A2( us12_n645 ) , .A1( us12_n646 ) );
  AOI222_X1 us12_U66 (.B2( us12_n638 ) , .ZN( us12_n644 ) , .B1( us12_n841 ) , .A1( us12_n842 ) , .C2( us12_n846 ) , .C1( us12_n863 ) , .A2( us12_n865 ) );
  NOR4_X1 us12_U67 (.A4( us12_n639 ) , .A3( us12_n640 ) , .A2( us12_n641 ) , .A1( us12_n642 ) , .ZN( us12_n643 ) );
  NOR3_X1 us12_U68 (.A2( us12_n607 ) , .A1( us12_n608 ) , .ZN( us12_n646 ) , .A3( us12_n722 ) );
  NAND4_X1 us12_U69 (.A4( us12_n603 ) , .A3( us12_n604 ) , .A2( us12_n605 ) , .A1( us12_n606 ) , .ZN( us12_n722 ) );
  NAND2_X1 us12_U7 (.A2( us12_n460 ) , .A1( us12_n465 ) , .ZN( us12_n780 ) );
  NOR3_X1 us12_U70 (.A1( us12_n599 ) , .ZN( us12_n604 ) , .A3( us12_n663 ) , .A2( us12_n770 ) );
  NOR4_X1 us12_U71 (.A3( us12_n600 ) , .A2( us12_n601 ) , .A1( us12_n602 ) , .ZN( us12_n603 ) , .A4( us12_n655 ) );
  AOI222_X1 us12_U72 (.ZN( us12_n606 ) , .A1( us12_n830 ) , .C2( us12_n837 ) , .B1( us12_n842 ) , .A2( us12_n856 ) , .B2( us12_n861 ) , .C1( us12_n868 ) );
  NOR4_X1 us12_U73 (.A4( us12_n514 ) , .A3( us12_n515 ) , .A2( us12_n516 ) , .A1( us12_n517 ) , .ZN( us12_n524 ) );
  AOI222_X1 us12_U74 (.ZN( us12_n525 ) , .A1( us12_n834 ) , .B2( us12_n837 ) , .C1( us12_n844 ) , .C2( us12_n850 ) , .A2( us12_n852 ) , .B1( us12_n866 ) );
  NOR4_X1 us12_U75 (.A3( us12_n521 ) , .A1( us12_n522 ) , .ZN( us12_n523 ) , .A2( us12_n673 ) , .A4( us12_n769 ) );
  NAND4_X1 us12_U76 (.A4( us12_n657 ) , .A3( us12_n658 ) , .A2( us12_n659 ) , .A1( us12_n660 ) , .ZN( us12_n800 ) );
  NOR3_X1 us12_U77 (.A3( us12_n648 ) , .A2( us12_n649 ) , .A1( us12_n650 ) , .ZN( us12_n659 ) );
  NOR3_X1 us12_U78 (.A3( us12_n651 ) , .A2( us12_n652 ) , .A1( us12_n653 ) , .ZN( us12_n658 ) );
  NOR3_X1 us12_U79 (.A3( us12_n654 ) , .A2( us12_n655 ) , .A1( us12_n656 ) , .ZN( us12_n657 ) );
  NOR3_X1 us12_U8 (.ZN( us12_n598 ) , .A1( us12_n608 ) , .A3( us12_n723 ) , .A2( us12_n742 ) );
  NAND4_X1 us12_U80 (.A4( us12_n560 ) , .A3( us12_n561 ) , .A2( us12_n562 ) , .A1( us12_n563 ) , .ZN( us12_n607 ) );
  NOR4_X1 us12_U81 (.A4( us12_n552 ) , .A3( us12_n553 ) , .A2( us12_n554 ) , .A1( us12_n555 ) , .ZN( us12_n562 ) );
  NOR4_X1 us12_U82 (.ZN( us12_n561 ) , .A1( us12_n653 ) , .A3( us12_n661 ) , .A4( us12_n685 ) , .A2( us12_n768 ) );
  NOR4_X1 us12_U83 (.A4( us12_n556 ) , .A3( us12_n557 ) , .A2( us12_n558 ) , .A1( us12_n559 ) , .ZN( us12_n560 ) );
  NAND4_X1 us12_U84 (.A4( us12_n772 ) , .A3( us12_n773 ) , .A2( us12_n774 ) , .A1( us12_n775 ) , .ZN( us12_n801 ) );
  NOR3_X1 us12_U85 (.A3( us12_n765 ) , .A2( us12_n766 ) , .A1( us12_n767 ) , .ZN( us12_n773 ) );
  NOR4_X1 us12_U86 (.A4( us12_n768 ) , .A3( us12_n769 ) , .A2( us12_n770 ) , .A1( us12_n771 ) , .ZN( us12_n772 ) );
  AOI222_X1 us12_U87 (.ZN( us12_n775 ) , .A1( us12_n830 ) , .C1( us12_n834 ) , .B2( us12_n841 ) , .A2( us12_n850 ) , .B1( us12_n861 ) , .C2( us12_n873 ) );
  NOR2_X1 us12_U88 (.ZN( us12_n625 ) , .A2( us12_n836 ) , .A1( us12_n839 ) );
  NOR2_X1 us12_U89 (.ZN( us12_n761 ) , .A1( us12_n833 ) , .A2( us12_n834 ) );
  NOR3_X1 us12_U9 (.A3( us12_n800 ) , .A2( us12_n801 ) , .A1( us12_n802 ) , .ZN( us12_n825 ) );
  AOI222_X1 us12_U90 (.ZN( us12_n513 ) , .C1( us12_n832 ) , .B2( us12_n837 ) , .A2( us12_n843 ) , .C2( us12_n862 ) , .B1( us12_n863 ) , .A1( us12_n866 ) );
  NOR4_X1 us12_U91 (.A4( us12_n509 ) , .A2( us12_n510 ) , .A1( us12_n511 ) , .ZN( us12_n512 ) , .A3( us12_n670 ) );
  INV_X1 us12_U92 (.A( us12_n505 ) , .ZN( us12_n871 ) );
  NAND4_X1 us12_U93 (.A4( us12_n456 ) , .A3( us12_n457 ) , .A2( us12_n458 ) , .A1( us12_n459 ) , .ZN( us12_n679 ) );
  NOR3_X1 us12_U94 (.ZN( us12_n457 ) , .A3( us12_n530 ) , .A1( us12_n555 ) , .A2( us12_n570 ) );
  AOI221_X1 us12_U95 (.A( us12_n450 ) , .ZN( us12_n459 ) , .C2( us12_n753 ) , .B1( us12_n832 ) , .C1( us12_n842 ) , .B2( us12_n861 ) );
  NOR4_X1 us12_U96 (.ZN( us12_n458 ) , .A2( us12_n509 ) , .A1( us12_n599 ) , .A4( us12_n628 ) , .A3( us12_n711 ) );
  NAND4_X1 us12_U97 (.A4( us12_n535 ) , .A3( us12_n536 ) , .A2( us12_n537 ) , .A1( us12_n538 ) , .ZN( us12_n622 ) );
  NOR4_X1 us12_U98 (.A4( us12_n526 ) , .A2( us12_n527 ) , .A1( us12_n528 ) , .ZN( us12_n538 ) , .A3( us12_n701 ) );
  NOR4_X1 us12_U99 (.A1( us12_n531 ) , .ZN( us12_n536 ) , .A2( us12_n654 ) , .A4( us12_n668 ) , .A3( us12_n765 ) );
  NOR3_X1 us31_U10 (.A3( us31_n621 ) , .A2( us31_n622 ) , .ZN( us31_n636 ) , .A1( us31_n725 ) );
  NOR4_X1 us31_U100 (.ZN( us31_n458 ) , .A2( us31_n509 ) , .A1( us31_n599 ) , .A4( us31_n628 ) , .A3( us31_n711 ) );
  NAND4_X1 us31_U101 (.A4( us31_n535 ) , .A3( us31_n536 ) , .A2( us31_n537 ) , .A1( us31_n538 ) , .ZN( us31_n622 ) );
  NOR4_X1 us31_U102 (.A4( us31_n526 ) , .A2( us31_n527 ) , .A1( us31_n528 ) , .ZN( us31_n538 ) , .A3( us31_n701 ) );
  NOR4_X1 us31_U103 (.A1( us31_n531 ) , .ZN( us31_n536 ) , .A2( us31_n654 ) , .A4( us31_n668 ) , .A3( us31_n765 ) );
  NOR4_X1 us31_U104 (.A4( us31_n529 ) , .A3( us31_n530 ) , .ZN( us31_n537 ) , .A2( us31_n684 ) , .A1( us31_n794 ) );
  NOR2_X1 us31_U105 (.ZN( us31_n647 ) , .A1( us31_n854 ) , .A2( us31_n868 ) );
  NAND4_X1 us31_U106 (.A4( us31_n548 ) , .A3( us31_n549 ) , .A2( us31_n550 ) , .A1( us31_n551 ) , .ZN( us31_n745 ) );
  NOR3_X1 us31_U107 (.ZN( us31_n549 ) , .A2( us31_n651 ) , .A1( us31_n667 ) , .A3( us31_n771 ) );
  AOI211_X1 us31_U108 (.B( us31_n539 ) , .A( us31_n540 ) , .ZN( us31_n551 ) , .C2( us31_n839 ) , .C1( us31_n851 ) );
  NOR4_X1 us31_U109 (.A4( us31_n541 ) , .A3( us31_n542 ) , .A2( us31_n543 ) , .ZN( us31_n550 ) , .A1( us31_n688 ) );
  NOR2_X1 us31_U11 (.A1( us31_n678 ) , .ZN( us31_n693 ) , .A2( us31_n807 ) );
  NAND4_X1 us31_U110 (.A4( us31_n479 ) , .A3( us31_n480 ) , .A2( us31_n481 ) , .A1( us31_n482 ) , .ZN( us31_n694 ) );
  NOR3_X1 us31_U111 (.ZN( us31_n480 ) , .A2( us31_n508 ) , .A3( us31_n601 ) , .A1( us31_n610 ) );
  AOI211_X1 us31_U112 (.B( us31_n477 ) , .A( us31_n478 ) , .ZN( us31_n482 ) , .C2( us31_n833 ) , .C1( us31_n861 ) );
  NOR4_X1 us31_U113 (.ZN( us31_n481 ) , .A3( us31_n532 ) , .A4( us31_n545 ) , .A2( us31_n567 ) , .A1( us31_n717 ) );
  NOR2_X1 us31_U114 (.ZN( us31_n686 ) , .A1( us31_n831 ) , .A2( us31_n832 ) );
  NAND4_X1 us31_U115 (.A4( us31_n485 ) , .A3( us31_n486 ) , .A2( us31_n487 ) , .A1( us31_n488 ) , .ZN( us31_n778 ) );
  NOR4_X1 us31_U116 (.A4( us31_n484 ) , .ZN( us31_n487 ) , .A1( us31_n566 ) , .A2( us31_n581 ) , .A3( us31_n602 ) );
  NOR4_X1 us31_U117 (.ZN( us31_n486 ) , .A1( us31_n507 ) , .A2( us31_n519 ) , .A4( us31_n546 ) , .A3( us31_n611 ) );
  NOR4_X1 us31_U118 (.ZN( us31_n485 ) , .A2( us31_n533 ) , .A1( us31_n558 ) , .A3( us31_n631 ) , .A4( us31_n718 ) );
  NAND4_X1 us31_U119 (.A4( us31_n691 ) , .A3( us31_n692 ) , .A1( us31_n693 ) , .ZN( us31_n776 ) , .A2( us31_n872 ) );
  NOR2_X1 us31_U12 (.ZN( us31_n495 ) , .A1( us31_n678 ) , .A2( us31_n694 ) );
  AOI221_X1 us31_U120 (.A( us31_n681 ) , .ZN( us31_n692 ) , .B2( us31_n840 ) , .C1( us31_n842 ) , .C2( us31_n862 ) , .B1( us31_n865 ) );
  INV_X1 us31_U121 (.A( us31_n679 ) , .ZN( us31_n872 ) );
  NOR4_X1 us31_U122 (.A4( us31_n687 ) , .A3( us31_n688 ) , .A2( us31_n689 ) , .A1( us31_n690 ) , .ZN( us31_n691 ) );
  NAND4_X1 us31_U123 (.A4( us31_n719 ) , .A3( us31_n720 ) , .A2( us31_n721 ) , .ZN( us31_n741 ) , .A1( us31_n857 ) );
  INV_X1 us31_U124 (.A( us31_n709 ) , .ZN( us31_n857 ) );
  AOI221_X1 us31_U125 (.A( us31_n710 ) , .ZN( us31_n721 ) , .C2( us31_n844 ) , .B2( us31_n845 ) , .C1( us31_n861 ) , .B1( us31_n862 ) );
  NOR4_X1 us31_U126 (.A4( us31_n715 ) , .A3( us31_n716 ) , .A2( us31_n717 ) , .A1( us31_n718 ) , .ZN( us31_n719 ) );
  NAND4_X1 us31_U127 (.A4( us31_n473 ) , .A3( us31_n474 ) , .A2( us31_n475 ) , .A1( us31_n476 ) , .ZN( us31_n678 ) );
  NOR4_X1 us31_U128 (.ZN( us31_n475 ) , .A1( us31_n531 ) , .A3( us31_n568 ) , .A4( us31_n600 ) , .A2( us31_n642 ) );
  NOR4_X1 us31_U129 (.ZN( us31_n473 ) , .A2( us31_n521 ) , .A4( us31_n594 ) , .A1( us31_n609 ) , .A3( us31_n629 ) );
  NOR3_X1 us31_U13 (.ZN( us31_n504 ) , .A2( us31_n679 ) , .A3( us31_n777 ) , .A1( us31_n876 ) );
  NOR4_X1 us31_U130 (.A4( us31_n470 ) , .ZN( us31_n476 ) , .A3( us31_n556 ) , .A1( us31_n735 ) , .A2( us31_n755 ) );
  NOR2_X1 us31_U131 (.ZN( us31_n733 ) , .A2( us31_n832 ) , .A1( us31_n845 ) );
  NOR2_X1 us31_U132 (.ZN( us31_n789 ) , .A2( us31_n862 ) , .A1( us31_n868 ) );
  NAND4_X1 us31_U133 (.A4( us31_n573 ) , .A3( us31_n574 ) , .A1( us31_n575 ) , .ZN( us31_n723 ) , .A2( us31_n874 ) );
  NOR4_X1 us31_U134 (.A4( us31_n569 ) , .A3( us31_n570 ) , .A2( us31_n571 ) , .A1( us31_n572 ) , .ZN( us31_n573 ) );
  AOI221_X1 us31_U135 (.A( us31_n564 ) , .C2( us31_n565 ) , .ZN( us31_n574 ) , .B2( us31_n845 ) , .B1( us31_n852 ) , .C1( us31_n853 ) );
  NOR2_X1 us31_U136 (.ZN( us31_n575 ) , .A1( us31_n622 ) , .A2( us31_n745 ) );
  NAND4_X1 us31_U137 (.A4( us31_n633 ) , .A3( us31_n634 ) , .A2( us31_n635 ) , .A1( us31_n636 ) , .ZN( us31_n743 ) );
  AOI211_X1 us31_U138 (.B( us31_n623 ) , .A( us31_n624 ) , .ZN( us31_n635 ) , .C2( us31_n836 ) , .C1( us31_n863 ) );
  NOR4_X1 us31_U139 (.A4( us31_n629 ) , .A3( us31_n630 ) , .A2( us31_n631 ) , .A1( us31_n632 ) , .ZN( us31_n633 ) );
  INV_X1 us31_U14 (.A( us31_n706 ) , .ZN( us31_n876 ) );
  NOR4_X1 us31_U140 (.A4( us31_n626 ) , .A3( us31_n627 ) , .A2( us31_n628 ) , .ZN( us31_n634 ) , .A1( us31_n664 ) );
  NAND4_X1 us31_U141 (.A4( us31_n493 ) , .A3( us31_n494 ) , .A1( us31_n495 ) , .ZN( us31_n802 ) , .A2( us31_n867 ) );
  AOI221_X1 us31_U142 (.A( us31_n489 ) , .ZN( us31_n494 ) , .B2( us31_n836 ) , .C2( us31_n841 ) , .C1( us31_n851 ) , .B1( us31_n860 ) );
  INV_X1 us31_U143 (.A( us31_n778 ) , .ZN( us31_n867 ) );
  NOR4_X1 us31_U144 (.A2( us31_n491 ) , .A1( us31_n492 ) , .ZN( us31_n493 ) , .A3( us31_n580 ) , .A4( us31_n612 ) );
  NOR4_X1 us31_U145 (.A4( us31_n734 ) , .A3( us31_n735 ) , .A2( us31_n736 ) , .A1( us31_n737 ) , .ZN( us31_n738 ) );
  AOI211_X1 us31_U146 (.B( us31_n725 ) , .A( us31_n726 ) , .ZN( us31_n739 ) , .C1( us31_n843 ) , .C2( us31_n855 ) );
  NOR3_X1 us31_U147 (.A3( us31_n722 ) , .A1( us31_n723 ) , .ZN( us31_n740 ) , .A2( us31_n741 ) );
  INV_X1 us31_U148 (.A( us31_n762 ) , .ZN( us31_n830 ) );
  INV_X1 us31_U149 (.A( us31_n697 ) , .ZN( us31_n838 ) );
  INV_X1 us31_U15 (.A( us31_n607 ) , .ZN( us31_n874 ) );
  OR4_X1 us31_U150 (.A4( us31_n566 ) , .A3( us31_n567 ) , .A2( us31_n568 ) , .ZN( us31_n572 ) , .A1( us31_n665 ) );
  OR4_X1 us31_U151 (.A4( us31_n682 ) , .A3( us31_n683 ) , .A2( us31_n684 ) , .A1( us31_n685 ) , .ZN( us31_n690 ) );
  OR4_X1 us31_U152 (.ZN( us31_n466 ) , .A4( us31_n518 ) , .A3( us31_n529 ) , .A2( us31_n578 ) , .A1( us31_n712 ) );
  OR4_X1 us31_U153 (.A4( us31_n518 ) , .A2( us31_n519 ) , .A1( us31_n520 ) , .ZN( us31_n522 ) , .A3( us31_n821 ) );
  OR4_X1 us31_U154 (.ZN( us31_n492 ) , .A4( us31_n534 ) , .A2( us31_n547 ) , .A1( us31_n559 ) , .A3( us31_n632 ) );
  OR4_X1 us31_U155 (.A4( us31_n580 ) , .A3( us31_n581 ) , .A2( us31_n582 ) , .A1( us31_n583 ) , .ZN( us31_n584 ) );
  NAND2_X1 us31_U156 (.ZN( us31_n613 ) , .A2( us31_n837 ) , .A1( us31_n873 ) );
  OR3_X1 us31_U157 (.A3( us31_n506 ) , .A2( us31_n507 ) , .A1( us31_n508 ) , .ZN( us31_n511 ) );
  INV_X1 us31_U158 (.A( us31_n463 ) , .ZN( us31_n864 ) );
  OAI21_X1 us31_U159 (.ZN( us31_n463 ) , .B1( us31_n809 ) , .A( us31_n834 ) , .B2( us31_n851 ) );
  INV_X1 us31_U16 (.A( us31_n680 ) , .ZN( us31_n840 ) );
  INV_X1 us31_U160 (.A( us31_n754 ) , .ZN( us31_n869 ) );
  OAI21_X1 us31_U161 (.B1( us31_n753 ) , .ZN( us31_n754 ) , .A( us31_n845 ) , .B2( us31_n868 ) );
  INV_X1 us31_U162 (.A( us31_n672 ) , .ZN( us31_n859 ) );
  AOI21_X1 us31_U163 (.A( us31_n670 ) , .B1( us31_n671 ) , .ZN( us31_n672 ) , .B2( us31_n856 ) );
  OAI222_X1 us31_U164 (.B2( us31_n747 ) , .B1( us31_n748 ) , .A2( us31_n749 ) , .ZN( us31_n757 ) , .C2( us31_n805 ) , .C1( us31_n814 ) , .A1( us31_n817 ) );
  OAI222_X1 us31_U165 (.ZN( us31_n505 ) , .C2( us31_n625 ) , .B2( us31_n647 ) , .B1( us31_n747 ) , .A2( us31_n748 ) , .C1( us31_n805 ) , .A1( us31_n806 ) );
  OAI222_X1 us31_U166 (.B2( us31_n708 ) , .ZN( us31_n709 ) , .C2( us31_n724 ) , .B1( us31_n747 ) , .A1( us31_n806 ) , .C1( us31_n814 ) , .A2( us31_n815 ) );
  NAND2_X1 us31_U167 (.A1( us31_n447 ) , .A2( us31_n465 ) , .ZN( us31_n749 ) );
  AOI22_X1 us31_U168 (.ZN( us31_n696 ) , .A1( us31_n830 ) , .B2( us31_n843 ) , .A2( us31_n865 ) , .B1( us31_n868 ) );
  AOI22_X1 us31_U169 (.A2( us31_n782 ) , .ZN( us31_n783 ) , .B2( us31_n831 ) , .A1( us31_n834 ) , .B1( us31_n863 ) );
  NOR4_X1 us31_U17 (.A4( us31_n445 ) , .A3( us31_n446 ) , .A2( us31_n516 ) , .A1( us31_n541 ) , .ZN( us31_n706 ) );
  INV_X1 us31_U170 (.A( us31_n730 ) , .ZN( us31_n839 ) );
  AOI221_X1 us31_U171 (.A( us31_n764 ) , .ZN( us31_n774 ) , .C2( us31_n810 ) , .B2( us31_n835 ) , .C1( us31_n855 ) , .B1( us31_n866 ) );
  AOI21_X1 us31_U172 (.B2( us31_n763 ) , .ZN( us31_n764 ) , .A( us31_n788 ) , .B1( us31_n792 ) );
  INV_X1 us31_U173 (.A( us31_n761 ) , .ZN( us31_n835 ) );
  AOI221_X1 us31_U174 (.A( us31_n483 ) , .ZN( us31_n488 ) , .B1( us31_n831 ) , .C2( us31_n844 ) , .C1( us31_n852 ) , .B2( us31_n862 ) );
  OAI22_X1 us31_U175 (.ZN( us31_n483 ) , .A1( us31_n708 ) , .B2( us31_n785 ) , .A2( us31_n806 ) , .B1( us31_n812 ) );
  INV_X1 us31_U176 (.A( us31_n790 ) , .ZN( us31_n832 ) );
  NAND2_X1 us31_U177 (.A1( us31_n451 ) , .A2( us31_n453 ) , .ZN( us31_n762 ) );
  AOI211_X1 us31_U178 (.A( us31_n637 ) , .ZN( us31_n645 ) , .B( us31_n743 ) , .C2( us31_n839 ) , .C1( us31_n854 ) );
  OAI22_X1 us31_U179 (.ZN( us31_n637 ) , .A1( us31_n699 ) , .B2( us31_n728 ) , .A2( us31_n762 ) , .B1( us31_n816 ) );
  OR3_X1 us31_U18 (.ZN( us31_n446 ) , .A1( us31_n528 ) , .A3( us31_n577 ) , .A2( us31_n875 ) );
  INV_X1 us31_U180 (.A( us31_n786 ) , .ZN( us31_n862 ) );
  OAI221_X1 us31_U181 (.A( us31_n727 ) , .C2( us31_n728 ) , .B2( us31_n729 ) , .B1( us31_n730 ) , .ZN( us31_n737 ) , .C1( us31_n817 ) );
  AOI22_X1 us31_U182 (.ZN( us31_n727 ) , .B1( us31_n832 ) , .A2( us31_n838 ) , .A1( us31_n863 ) , .B2( us31_n866 ) );
  OAI22_X1 us31_U183 (.ZN( us31_n710 ) , .A2( us31_n728 ) , .B2( us31_n729 ) , .A1( us31_n744 ) , .B1( us31_n813 ) );
  INV_X1 us31_U184 (.A( us31_n816 ) , .ZN( us31_n831 ) );
  OAI22_X1 us31_U185 (.ZN( us31_n624 ) , .B1( us31_n669 ) , .B2( us31_n747 ) , .A1( us31_n815 ) , .A2( us31_n816 ) );
  INV_X1 us31_U186 (.A( us31_n744 ) , .ZN( us31_n837 ) );
  INV_X1 us31_U187 (.A( us31_n788 ) , .ZN( us31_n845 ) );
  OAI22_X1 us31_U188 (.B2( us31_n779 ) , .B1( us31_n780 ) , .ZN( us31_n781 ) , .A2( us31_n814 ) , .A1( us31_n815 ) );
  OAI22_X1 us31_U189 (.A1( us31_n724 ) , .ZN( us31_n726 ) , .B2( us31_n750 ) , .B1( us31_n812 ) , .A2( us31_n816 ) );
  OR4_X1 us31_U19 (.A4( us31_n442 ) , .A2( us31_n443 ) , .A1( us31_n444 ) , .ZN( us31_n445 ) , .A3( us31_n553 ) );
  INV_X1 us31_U190 (.A( us31_n805 ) , .ZN( us31_n860 ) );
  INV_X1 us31_U191 (.A( us31_n814 ) , .ZN( us31_n833 ) );
  INV_X1 us31_U192 (.A( us31_n669 ) , .ZN( us31_n865 ) );
  OAI22_X1 us31_U193 (.B2( us31_n744 ) , .ZN( us31_n746 ) , .A2( us31_n762 ) , .B1( us31_n780 ) , .A1( us31_n792 ) );
  OAI22_X1 us31_U194 (.ZN( us31_n496 ) , .A2( us31_n744 ) , .A1( us31_n780 ) , .B1( us31_n791 ) , .B2( us31_n806 ) );
  OAI22_X1 us31_U195 (.B2( us31_n803 ) , .B1( us31_n804 ) , .A2( us31_n805 ) , .A1( us31_n806 ) , .ZN( us31_n808 ) );
  OAI22_X1 us31_U196 (.ZN( us31_n489 ) , .A1( us31_n724 ) , .B2( us31_n728 ) , .B1( us31_n730 ) , .A2( us31_n779 ) );
  OAI22_X1 us31_U197 (.ZN( us31_n695 ) , .A2( us31_n730 ) , .A1( us31_n780 ) , .B1( us31_n791 ) , .B2( us31_n817 ) );
  OAI22_X1 us31_U198 (.B1( us31_n490 ) , .ZN( us31_n491 ) , .A1( us31_n686 ) , .A2( us31_n763 ) , .B2( us31_n817 ) );
  NOR3_X1 us31_U199 (.ZN( us31_n490 ) , .A1( us31_n782 ) , .A2( us31_n850 ) , .A3( us31_n863 ) );
  INV_X1 us31_U20 (.A( us31_n613 ) , .ZN( us31_n875 ) );
  INV_X1 us31_U200 (.A( us31_n750 ) , .ZN( us31_n842 ) );
  NOR2_X1 us31_U201 (.ZN( us31_n715 ) , .A1( us31_n805 ) , .A2( us31_n817 ) );
  NOR2_X1 us31_U202 (.A2( us31_n744 ) , .ZN( us31_n755 ) , .A1( us31_n805 ) );
  NOR2_X1 us31_U203 (.ZN( us31_n735 ) , .A2( us31_n803 ) , .A1( us31_n805 ) );
  NOR2_X1 us31_U204 (.ZN( us31_n546 ) , .A2( us31_n780 ) , .A1( us31_n814 ) );
  NOR2_X1 us31_U205 (.ZN( us31_n577 ) , .A2( us31_n699 ) , .A1( us31_n814 ) );
  NOR2_X1 us31_U206 (.ZN( us31_n718 ) , .A2( us31_n724 ) , .A1( us31_n744 ) );
  NOR2_X1 us31_U207 (.ZN( us31_n532 ) , .A2( us31_n749 ) , .A1( us31_n750 ) );
  NOR2_X1 us31_U208 (.ZN( us31_n615 ) , .A1( us31_n785 ) , .A2( us31_n815 ) );
  NOR2_X1 us31_U209 (.ZN( us31_n629 ) , .A2( us31_n728 ) , .A1( us31_n785 ) );
  INV_X1 us31_U21 (.A( us31_n749 ) , .ZN( us31_n863 ) );
  NOR2_X1 us31_U210 (.ZN( us31_n611 ) , .A2( us31_n780 ) , .A1( us31_n806 ) );
  NOR2_X1 us31_U211 (.ZN( us31_n652 ) , .A1( us31_n669 ) , .A2( us31_n814 ) );
  NOR2_X1 us31_U212 (.A1( us31_n669 ) , .ZN( us31_n673 ) , .A2( us31_n744 ) );
  NOR2_X1 us31_U213 (.ZN( us31_n602 ) , .A1( us31_n669 ) , .A2( us31_n803 ) );
  NOR2_X1 us31_U214 (.A1( us31_n669 ) , .ZN( us31_n688 ) , .A2( us31_n816 ) );
  NOR2_X1 us31_U215 (.ZN( us31_n628 ) , .A2( us31_n669 ) , .A1( us31_n785 ) );
  INV_X1 us31_U216 (.A( us31_n747 ) , .ZN( us31_n834 ) );
  NOR2_X1 us31_U217 (.A1( us31_n669 ) , .ZN( us31_n766 ) , .A2( us31_n813 ) );
  NOR2_X1 us31_U218 (.A2( us31_n744 ) , .ZN( us31_n769 ) , .A1( us31_n812 ) );
  NOR2_X1 us31_U219 (.ZN( us31_n527 ) , .A1( us31_n669 ) , .A2( us31_n779 ) );
  AOI222_X1 us31_U22 (.ZN( us31_n605 ) , .B2( us31_n671 ) , .B1( us31_n753 ) , .C2( us31_n831 ) , .A1( us31_n833 ) , .A2( us31_n862 ) , .C1( us31_n863 ) );
  NOR2_X1 us31_U220 (.ZN( us31_n531 ) , .A2( us31_n780 ) , .A1( us31_n816 ) );
  INV_X1 us31_U221 (.A( us31_n792 ) , .ZN( us31_n851 ) );
  NOR2_X1 us31_U222 (.A2( us31_n708 ) , .A1( us31_n750 ) , .ZN( us31_n771 ) );
  NOR2_X1 us31_U223 (.ZN( us31_n599 ) , .A2( us31_n791 ) , .A1( us31_n816 ) );
  NOR2_X1 us31_U224 (.ZN( us31_n601 ) , .A2( us31_n780 ) , .A1( us31_n803 ) );
  NOR2_X1 us31_U225 (.A1( us31_n699 ) , .ZN( us31_n768 ) , .A2( us31_n813 ) );
  NOR2_X1 us31_U226 (.ZN( us31_n541 ) , .A2( us31_n697 ) , .A1( us31_n699 ) );
  NOR2_X1 us31_U227 (.ZN( us31_n667 ) , .A1( us31_n750 ) , .A2( us31_n815 ) );
  NOR2_X1 us31_U228 (.ZN( us31_n555 ) , .A1( us31_n750 ) , .A2( us31_n791 ) );
  NOR2_X1 us31_U229 (.ZN( us31_n508 ) , .A2( us31_n780 ) , .A1( us31_n785 ) );
  AOI222_X1 us31_U23 (.ZN( us31_n563 ) , .B1( us31_n830 ) , .C1( us31_n841 ) , .A2( us31_n843 ) , .A1( us31_n854 ) , .B2( us31_n863 ) , .C2( us31_n873 ) );
  NOR2_X1 us31_U230 (.ZN( us31_n543 ) , .A2( us31_n708 ) , .A1( us31_n785 ) );
  NOR2_X1 us31_U231 (.ZN( us31_n528 ) , .A2( us31_n724 ) , .A1( us31_n803 ) );
  NOR2_X1 us31_U232 (.ZN( us31_n664 ) , .A1( us31_n785 ) , .A2( us31_n791 ) );
  NOR2_X1 us31_U233 (.ZN( us31_n556 ) , .A1( us31_n762 ) , .A2( us31_n805 ) );
  INV_X1 us31_U234 (.A( us31_n806 ) , .ZN( us31_n841 ) );
  OAI22_X1 us31_U235 (.B1( us31_n440 ) , .ZN( us31_n444 ) , .A2( us31_n728 ) , .A1( us31_n744 ) , .B2( us31_n749 ) );
  NOR3_X1 us31_U236 (.ZN( us31_n440 ) , .A2( us31_n836 ) , .A3( us31_n837 ) , .A1( us31_n846 ) );
  NOR2_X1 us31_U237 (.ZN( us31_n507 ) , .A1( us31_n812 ) , .A2( us31_n817 ) );
  NOR2_X1 us31_U238 (.ZN( us31_n557 ) , .A1( us31_n792 ) , .A2( us31_n814 ) );
  NOR2_X1 us31_U239 (.ZN( us31_n545 ) , .A1( us31_n749 ) , .A2( us31_n814 ) );
  AOI222_X1 us31_U24 (.ZN( us31_n660 ) , .A2( us31_n839 ) , .B1( us31_n841 ) , .C2( us31_n845 ) , .A1( us31_n860 ) , .C1( us31_n863 ) , .B2( us31_n870 ) );
  OAI22_X1 us31_U240 (.B2( us31_n750 ) , .B1( us31_n751 ) , .A1( us31_n752 ) , .ZN( us31_n756 ) , .A2( us31_n806 ) );
  NOR2_X1 us31_U241 (.ZN( us31_n751 ) , .A2( us31_n852 ) , .A1( us31_n860 ) );
  NOR3_X1 us31_U242 (.ZN( us31_n752 ) , .A2( us31_n853 ) , .A1( us31_n863 ) , .A3( us31_n865 ) );
  NOR2_X1 us31_U243 (.ZN( us31_n544 ) , .A2( us31_n785 ) , .A1( us31_n792 ) );
  NOR2_X1 us31_U244 (.ZN( us31_n530 ) , .A2( us31_n744 ) , .A1( us31_n792 ) );
  NOR2_X1 us31_U245 (.ZN( us31_n509 ) , .A1( us31_n729 ) , .A2( us31_n779 ) );
  NOR2_X1 us31_U246 (.ZN( us31_n570 ) , .A1( us31_n728 ) , .A2( us31_n806 ) );
  NOR2_X1 us31_U247 (.ZN( us31_n666 ) , .A1( us31_n728 ) , .A2( us31_n803 ) );
  NOR2_X1 us31_U248 (.ZN( us31_n631 ) , .A1( us31_n724 ) , .A2( us31_n813 ) );
  NOR2_X1 us31_U249 (.ZN( us31_n614 ) , .A1( us31_n762 ) , .A2( us31_n812 ) );
  INV_X1 us31_U25 (.A( us31_n647 ) , .ZN( us31_n870 ) );
  NOR2_X1 us31_U250 (.A1( us31_n749 ) , .ZN( us31_n767 ) , .A2( us31_n803 ) );
  NOR2_X1 us31_U251 (.ZN( us31_n654 ) , .A1( us31_n728 ) , .A2( us31_n813 ) );
  NOR2_X1 us31_U252 (.ZN( us31_n516 ) , .A1( us31_n708 ) , .A2( us31_n744 ) );
  NOR2_X1 us31_U253 (.ZN( us31_n670 ) , .A1( us31_n790 ) , .A2( us31_n805 ) );
  NOR2_X1 us31_U254 (.ZN( us31_n558 ) , .A1( us31_n708 ) , .A2( us31_n816 ) );
  INV_X1 us31_U255 (.A( us31_n763 ) , .ZN( us31_n866 ) );
  NOR2_X1 us31_U256 (.ZN( us31_n663 ) , .A1( us31_n729 ) , .A2( us31_n785 ) );
  NOR2_X1 us31_U257 (.A2( us31_n697 ) , .ZN( us31_n716 ) , .A1( us31_n792 ) );
  NOR2_X1 us31_U258 (.ZN( us31_n517 ) , .A1( us31_n708 ) , .A2( us31_n803 ) );
  NOR2_X1 us31_U259 (.ZN( us31_n521 ) , .A1( us31_n790 ) , .A2( us31_n812 ) );
  NOR4_X1 us31_U26 (.A4( us31_n544 ) , .A3( us31_n545 ) , .A2( us31_n546 ) , .A1( us31_n547 ) , .ZN( us31_n548 ) );
  NOR2_X1 us31_U260 (.ZN( us31_n630 ) , .A1( us31_n747 ) , .A2( us31_n815 ) );
  NOR2_X1 us31_U261 (.ZN( us31_n655 ) , .A1( us31_n790 ) , .A2( us31_n815 ) );
  AOI21_X1 us31_U262 (.ZN( us31_n552 ) , .B1( us31_n669 ) , .A( us31_n697 ) , .B2( us31_n805 ) );
  NOR2_X1 us31_U263 (.ZN( us31_n668 ) , .A2( us31_n708 ) , .A1( us31_n790 ) );
  NOR2_X1 us31_U264 (.ZN( us31_n594 ) , .A2( us31_n697 ) , .A1( us31_n728 ) );
  NOR2_X1 us31_U265 (.ZN( us31_n542 ) , .A1( us31_n762 ) , .A2( us31_n791 ) );
  NOR2_X1 us31_U266 (.ZN( us31_n656 ) , .A1( us31_n747 ) , .A2( us31_n780 ) );
  NOR2_X1 us31_U267 (.ZN( us31_n609 ) , .A2( us31_n724 ) , .A1( us31_n817 ) );
  AOI21_X1 us31_U268 (.B1( us31_n625 ) , .ZN( us31_n627 ) , .A( us31_n763 ) , .B2( us31_n814 ) );
  NOR2_X1 us31_U269 (.ZN( us31_n661 ) , .A1( us31_n729 ) , .A2( us31_n790 ) );
  NOR4_X1 us31_U27 (.ZN( us31_n479 ) , .A1( us31_n520 ) , .A4( us31_n557 ) , .A3( us31_n582 ) , .A2( us31_n630 ) );
  NOR2_X1 us31_U270 (.ZN( us31_n642 ) , .A2( us31_n788 ) , .A1( us31_n791 ) );
  AOI21_X1 us31_U271 (.ZN( us31_n650 ) , .A( us31_n779 ) , .B1( us31_n792 ) , .B2( us31_n805 ) );
  AOI21_X1 us31_U272 (.ZN( us31_n626 ) , .B2( us31_n669 ) , .A( us31_n790 ) , .B1( us31_n791 ) );
  AOI21_X1 us31_U273 (.A( us31_n815 ) , .B2( us31_n816 ) , .B1( us31_n817 ) , .ZN( us31_n818 ) );
  NOR2_X1 us31_U274 (.ZN( us31_n579 ) , .A2( us31_n708 ) , .A1( us31_n730 ) );
  NOR2_X1 us31_U275 (.ZN( us31_n533 ) , .A2( us31_n724 ) , .A1( us31_n730 ) );
  AOI21_X1 us31_U276 (.A( us31_n812 ) , .B2( us31_n813 ) , .B1( us31_n814 ) , .ZN( us31_n819 ) );
  NOR2_X1 us31_U277 (.A2( us31_n708 ) , .A1( us31_n762 ) , .ZN( us31_n794 ) );
  NOR2_X1 us31_U278 (.A2( us31_n697 ) , .A1( us31_n780 ) , .ZN( us31_n820 ) );
  AOI21_X1 us31_U279 (.ZN( us31_n499 ) , .B1( us31_n680 ) , .A( us31_n812 ) , .B2( us31_n816 ) );
  NOR4_X1 us31_U28 (.ZN( us31_n456 ) , .A2( us31_n517 ) , .A1( us31_n543 ) , .A3( us31_n579 ) , .A4( us31_n615 ) );
  NOR2_X1 us31_U280 (.ZN( us31_n520 ) , .A2( us31_n708 ) , .A1( us31_n814 ) );
  AOI21_X1 us31_U281 (.ZN( us31_n477 ) , .A( us31_n669 ) , .B1( us31_n750 ) , .B2( us31_n806 ) );
  NOR2_X1 us31_U282 (.ZN( us31_n582 ) , .A1( us31_n744 ) , .A2( us31_n815 ) );
  NOR2_X1 us31_U283 (.ZN( us31_n662 ) , .A2( us31_n697 ) , .A1( us31_n729 ) );
  AOI21_X1 us31_U284 (.ZN( us31_n593 ) , .B1( us31_n750 ) , .A( us31_n792 ) , .B2( us31_n813 ) );
  AOI21_X1 us31_U285 (.ZN( us31_n515 ) , .A( us31_n729 ) , .B1( us31_n750 ) , .B2( us31_n803 ) );
  AOI21_X1 us31_U286 (.ZN( us31_n510 ) , .B2( us31_n669 ) , .A( us31_n730 ) , .B1( us31_n815 ) );
  NOR2_X1 us31_U287 (.ZN( us31_n506 ) , .A2( us31_n728 ) , .A1( us31_n762 ) );
  NOR2_X1 us31_U288 (.A1( us31_n697 ) , .ZN( us31_n770 ) , .A2( us31_n815 ) );
  NOR2_X1 us31_U289 (.ZN( us31_n519 ) , .A2( us31_n699 ) , .A1( us31_n816 ) );
  NOR4_X1 us31_U29 (.A4( us31_n532 ) , .A3( us31_n533 ) , .A2( us31_n534 ) , .ZN( us31_n535 ) , .A1( us31_n820 ) );
  NOR2_X1 us31_U290 (.ZN( us31_n581 ) , .A1( us31_n669 ) , .A2( us31_n788 ) );
  NOR2_X1 us31_U291 (.ZN( us31_n559 ) , .A2( us31_n791 ) , .A1( us31_n803 ) );
  AOI21_X1 us31_U292 (.B1( us31_n699 ) , .ZN( us31_n700 ) , .A( us31_n732 ) , .B2( us31_n763 ) );
  AOI21_X1 us31_U293 (.ZN( us31_n591 ) , .B2( us31_n763 ) , .A( us31_n785 ) , .B1( us31_n812 ) );
  INV_X1 us31_U294 (.A( us31_n813 ) , .ZN( us31_n836 ) );
  NOR2_X1 us31_U295 (.ZN( us31_n683 ) , .A2( us31_n699 ) , .A1( us31_n803 ) );
  AOI21_X1 us31_U296 (.ZN( us31_n589 ) , .B2( us31_n699 ) , .B1( us31_n815 ) , .A( us31_n817 ) );
  AOI21_X1 us31_U297 (.ZN( us31_n539 ) , .B2( us31_n812 ) , .A( us31_n814 ) , .B1( us31_n815 ) );
  INV_X1 us31_U298 (.A( us31_n728 ) , .ZN( us31_n852 ) );
  AOI21_X1 us31_U299 (.ZN( us31_n540 ) , .A( us31_n763 ) , .B2( us31_n779 ) , .B1( us31_n817 ) );
  NAND2_X1 us31_U3 (.A1( us31_n449 ) , .A2( us31_n460 ) , .ZN( us31_n792 ) );
  NOR4_X1 us31_U30 (.ZN( us31_n474 ) , .A1( us31_n506 ) , .A3( us31_n544 ) , .A2( us31_n583 ) , .A4( us31_n716 ) );
  INV_X1 us31_U300 (.A( us31_n791 ) , .ZN( us31_n873 ) );
  AOI21_X1 us31_U301 (.ZN( us31_n498 ) , .A( us31_n724 ) , .B2( us31_n762 ) , .B1( us31_n814 ) );
  AOI21_X1 us31_U302 (.ZN( us31_n649 ) , .B1( us31_n729 ) , .B2( us31_n763 ) , .A( us31_n813 ) );
  NOR2_X1 us31_U303 (.ZN( us31_n547 ) , .A1( us31_n699 ) , .A2( us31_n744 ) );
  NOR2_X1 us31_U304 (.ZN( us31_n566 ) , .A2( us31_n697 ) , .A1( us31_n763 ) );
  AOI21_X1 us31_U305 (.ZN( us31_n569 ) , .B1( us31_n750 ) , .B2( us31_n762 ) , .A( us31_n780 ) );
  AOI21_X1 us31_U306 (.ZN( us31_n571 ) , .B2( us31_n697 ) , .B1( us31_n806 ) , .A( us31_n812 ) );
  AOI21_X1 us31_U307 (.ZN( us31_n640 ) , .B2( us31_n747 ) , .A( us31_n792 ) , .B1( us31_n803 ) );
  INV_X1 us31_U308 (.A( us31_n699 ) , .ZN( us31_n853 ) );
  AOI21_X1 us31_U309 (.ZN( us31_n514 ) , .A( us31_n779 ) , .B2( us31_n792 ) , .B1( us31_n812 ) );
  AOI221_X1 us31_U31 (.A( us31_n713 ) , .B2( us31_n714 ) , .ZN( us31_n720 ) , .C1( us31_n832 ) , .B1( us31_n839 ) , .C2( us31_n863 ) );
  AOI21_X1 us31_U310 (.ZN( us31_n639 ) , .B2( us31_n749 ) , .A( us31_n788 ) , .B1( us31_n812 ) );
  NAND2_X1 us31_U311 (.ZN( us31_n753 ) , .A1( us31_n763 ) , .A2( us31_n805 ) );
  NOR2_X1 us31_U312 (.ZN( us31_n665 ) , .A1( us31_n780 ) , .A2( us31_n813 ) );
  INV_X1 us31_U313 (.A( us31_n729 ) , .ZN( us31_n868 ) );
  NOR2_X1 us31_U314 (.ZN( us31_n685 ) , .A1( us31_n729 ) , .A2( us31_n816 ) );
  AOI21_X1 us31_U315 (.ZN( us31_n564 ) , .B1( us31_n724 ) , .A( us31_n779 ) , .B2( us31_n791 ) );
  AOI21_X1 us31_U316 (.ZN( us31_n497 ) , .A( us31_n779 ) , .B2( us31_n791 ) , .B1( us31_n804 ) );
  AOI21_X1 us31_U317 (.ZN( us31_n689 ) , .B2( us31_n749 ) , .B1( us31_n763 ) , .A( us31_n806 ) );
  AOI21_X1 us31_U318 (.ZN( us31_n450 ) , .B2( us31_n792 ) , .A( us31_n803 ) , .B1( us31_n815 ) );
  NOR2_X1 us31_U319 (.ZN( us31_n567 ) , .A1( us31_n747 ) , .A2( us31_n805 ) );
  OR2_X1 us31_U32 (.A2( us31_n711 ) , .A1( us31_n712 ) , .ZN( us31_n713 ) );
  NOR2_X1 us31_U320 (.ZN( us31_n529 ) , .A1( us31_n708 ) , .A2( us31_n779 ) );
  NOR2_X1 us31_U321 (.ZN( us31_n578 ) , .A1( us31_n708 ) , .A2( us31_n813 ) );
  AOI21_X1 us31_U322 (.ZN( us31_n478 ) , .B2( us31_n697 ) , .A( us31_n749 ) , .B1( us31_n779 ) );
  AOI21_X1 us31_U323 (.A( us31_n790 ) , .B2( us31_n791 ) , .B1( us31_n792 ) , .ZN( us31_n793 ) );
  NOR2_X1 us31_U324 (.ZN( us31_n684 ) , .A1( us31_n791 ) , .A2( us31_n813 ) );
  AOI21_X1 us31_U325 (.A( us31_n733 ) , .ZN( us31_n734 ) , .B2( us31_n780 ) , .B1( us31_n792 ) );
  NOR2_X1 us31_U326 (.A2( us31_n813 ) , .A1( us31_n815 ) , .ZN( us31_n821 ) );
  NOR2_X1 us31_U327 (.ZN( us31_n711 ) , .A1( us31_n762 ) , .A2( us31_n763 ) );
  AOI21_X1 us31_U328 (.ZN( us31_n641 ) , .B1( us31_n680 ) , .A( us31_n791 ) , .B2( us31_n817 ) );
  NOR2_X1 us31_U329 (.ZN( us31_n580 ) , .A2( us31_n697 ) , .A1( us31_n791 ) );
  NOR2_X1 us31_U33 (.ZN( us31_n680 ) , .A2( us31_n834 ) , .A1( us31_n839 ) );
  NOR2_X1 us31_U330 (.ZN( us31_n583 ) , .A1( us31_n792 ) , .A2( us31_n817 ) );
  NOR2_X1 us31_U331 (.ZN( us31_n534 ) , .A1( us31_n724 ) , .A2( us31_n788 ) );
  NOR2_X1 us31_U332 (.ZN( us31_n632 ) , .A2( us31_n697 ) , .A1( us31_n724 ) );
  NOR2_X1 us31_U333 (.ZN( us31_n682 ) , .A2( us31_n708 ) , .A1( us31_n817 ) );
  AOI21_X1 us31_U334 (.B1( us31_n686 ) , .ZN( us31_n687 ) , .A( us31_n728 ) , .B2( us31_n761 ) );
  INV_X1 us31_U335 (.A( us31_n815 ) , .ZN( us31_n855 ) );
  AOI21_X1 us31_U336 (.ZN( us31_n442 ) , .A( us31_n699 ) , .B1( us31_n733 ) , .B2( us31_n750 ) );
  NOR2_X1 us31_U337 (.ZN( us31_n568 ) , .A1( us31_n729 ) , .A2( us31_n762 ) );
  INV_X1 us31_U338 (.A( us31_n780 ) , .ZN( us31_n850 ) );
  INV_X1 us31_U339 (.A( us31_n785 ) , .ZN( us31_n846 ) );
  AOI222_X1 us31_U34 (.ZN( us31_n469 ) , .B1( us31_n832 ) , .A1( us31_n839 ) , .C1( us31_n842 ) , .C2( us31_n851 ) , .A2( us31_n855 ) , .B2( us31_n865 ) );
  NAND2_X1 us31_U340 (.A2( us31_n762 ) , .A1( us31_n806 ) , .ZN( us31_n810 ) );
  AOI21_X1 us31_U341 (.ZN( us31_n443 ) , .B1( us31_n789 ) , .B2( us31_n791 ) , .A( us31_n814 ) );
  NAND2_X1 us31_U342 (.ZN( us31_n671 ) , .A1( us31_n806 ) , .A2( us31_n816 ) );
  NOR2_X1 us31_U343 (.ZN( us31_n484 ) , .A1( us31_n788 ) , .A2( us31_n805 ) );
  NOR2_X1 us31_U344 (.ZN( us31_n470 ) , .A2( us31_n779 ) , .A1( us31_n815 ) );
  NOR2_X1 us31_U345 (.ZN( us31_n712 ) , .A2( us31_n724 ) , .A1( us31_n790 ) );
  OAI21_X1 us31_U346 (.A( us31_n787 ) , .B2( us31_n788 ) , .B1( us31_n789 ) , .ZN( us31_n795 ) );
  OAI21_X1 us31_U347 (.ZN( us31_n787 ) , .A( us31_n839 ) , .B1( us31_n863 ) , .B2( us31_n873 ) );
  NOR2_X1 us31_U348 (.ZN( us31_n526 ) , .A1( us31_n724 ) , .A2( us31_n750 ) );
  NAND2_X1 us31_U349 (.A1( us31_n699 ) , .A2( us31_n729 ) , .ZN( us31_n782 ) );
  NOR4_X1 us31_U35 (.A1( us31_n466 ) , .ZN( us31_n467 ) , .A4( us31_n542 ) , .A2( us31_n554 ) , .A3( us31_n614 ) );
  NOR2_X1 us31_U350 (.ZN( us31_n518 ) , .A1( us31_n708 ) , .A2( us31_n788 ) );
  OAI21_X1 us31_U351 (.A( us31_n698 ) , .ZN( us31_n702 ) , .B2( us31_n750 ) , .B1( us31_n804 ) );
  OAI21_X1 us31_U352 (.ZN( us31_n698 ) , .B2( us31_n833 ) , .B1( us31_n838 ) , .A( us31_n860 ) );
  INV_X1 us31_U353 (.A( us31_n817 ) , .ZN( us31_n844 ) );
  OAI21_X1 us31_U354 (.A( us31_n731 ) , .B1( us31_n732 ) , .ZN( us31_n736 ) , .B2( us31_n805 ) );
  OAI21_X1 us31_U355 (.ZN( us31_n731 ) , .A( us31_n833 ) , .B2( us31_n852 ) , .B1( us31_n873 ) );
  NAND2_X1 us31_U356 (.ZN( us31_n714 ) , .A1( us31_n728 ) , .A2( us31_n780 ) );
  INV_X1 us31_U357 (.A( us31_n724 ) , .ZN( us31_n856 ) );
  AND2_X1 us31_U358 (.ZN( us31_n732 ) , .A1( us31_n779 ) , .A2( us31_n785 ) );
  NAND2_X1 us31_U359 (.A1( us31_n447 ) , .A2( us31_n449 ) , .ZN( us31_n805 ) );
  AOI221_X1 us31_U36 (.ZN( us31_n468 ) , .C2( us31_n714 ) , .B2( us31_n831 ) , .C1( us31_n845 ) , .B1( us31_n860 ) , .A( us31_n864 ) );
  NAND2_X1 us31_U360 (.A1( us31_n451 ) , .A2( us31_n454 ) , .ZN( us31_n814 ) );
  NAND2_X1 us31_U361 (.A1( us31_n452 ) , .A2( us31_n465 ) , .ZN( us31_n669 ) );
  NAND2_X1 us31_U362 (.A1( us31_n455 ) , .A2( us31_n462 ) , .ZN( us31_n750 ) );
  NAND2_X1 us31_U363 (.A2( us31_n453 ) , .A1( us31_n455 ) , .ZN( us31_n806 ) );
  NAND2_X1 us31_U364 (.A1( us31_n451 ) , .A2( us31_n471 ) , .ZN( us31_n816 ) );
  NAND2_X1 us31_U365 (.A1( us31_n454 ) , .A2( us31_n461 ) , .ZN( us31_n813 ) );
  NAND2_X1 us31_U366 (.A1( us31_n455 ) , .A2( us31_n471 ) , .ZN( us31_n803 ) );
  NAND2_X1 us31_U367 (.A1( us31_n453 ) , .A2( us31_n461 ) , .ZN( us31_n744 ) );
  NAND2_X1 us31_U368 (.A1( us31_n453 ) , .A2( us31_n472 ) , .ZN( us31_n785 ) );
  NAND2_X1 us31_U369 (.A2( us31_n454 ) , .A1( us31_n472 ) , .ZN( us31_n779 ) );
  NOR4_X1 us31_U37 (.A4( us31_n577 ) , .A3( us31_n578 ) , .A2( us31_n579 ) , .ZN( us31_n586 ) , .A1( us31_n683 ) );
  NAND2_X1 us31_U370 (.A2( us31_n464 ) , .A1( us31_n465 ) , .ZN( us31_n812 ) );
  NAND2_X1 us31_U371 (.A1( us31_n441 ) , .A2( us31_n460 ) , .ZN( us31_n699 ) );
  NAND2_X1 us31_U372 (.A2( us31_n449 ) , .A1( us31_n452 ) , .ZN( us31_n763 ) );
  NAND2_X1 us31_U373 (.A2( us31_n461 ) , .A1( us31_n462 ) , .ZN( us31_n747 ) );
  NAND2_X1 us31_U374 (.A1( us31_n462 ) , .A2( us31_n472 ) , .ZN( us31_n788 ) );
  NOR2_X1 us31_U375 (.ZN( us31_n465 ) , .A2( us31_n847 ) , .A1( us31_n848 ) );
  NOR2_X1 us31_U376 (.ZN( us31_n453 ) , .A1( us31_n826 ) , .A2( us31_n827 ) );
  NOR2_X1 us31_U377 (.ZN( us31_n451 ) , .A1( us31_n828 ) , .A2( us31_n829 ) );
  NAND2_X1 us31_U378 (.A1( us31_n451 ) , .A2( us31_n462 ) , .ZN( us31_n790 ) );
  NAND2_X1 us31_U379 (.A2( us31_n441 ) , .A1( us31_n447 ) , .ZN( us31_n784 ) );
  NOR4_X1 us31_U38 (.A1( us31_n584 ) , .ZN( us31_n585 ) , .A3( us31_n652 ) , .A2( us31_n662 ) , .A4( us31_n767 ) );
  NAND2_X1 us31_U380 (.A2( us31_n454 ) , .A1( us31_n455 ) , .ZN( us31_n730 ) );
  NAND2_X2 us31_U381 (.A1( us31_n449 ) , .A2( us31_n464 ) , .ZN( us31_n724 ) );
  NAND2_X2 us31_U382 (.A2( us31_n460 ) , .A1( us31_n465 ) , .ZN( us31_n780 ) );
  NOR2_X1 us31_U383 (.ZN( us31_n447 ) , .A2( us31_n849 ) , .A1( us31_n858 ) );
  NAND2_X1 us31_U384 (.A1( us31_n447 ) , .A2( us31_n448 ) , .ZN( us31_n786 ) );
  NAND2_X1 us31_U385 (.A2( us31_n448 ) , .A1( us31_n460 ) , .ZN( us31_n728 ) );
  NAND2_X1 us31_U386 (.A2( us31_n448 ) , .A1( us31_n452 ) , .ZN( us31_n729 ) );
  NOR2_X1 us31_U387 (.A2( sa31_5 ) , .ZN( us31_n448 ) , .A1( us31_n847 ) );
  NOR2_X1 us31_U388 (.A2( sa31_7 ) , .ZN( us31_n460 ) , .A1( us31_n849 ) );
  NOR2_X1 us31_U389 (.A2( sa31_6 ) , .A1( sa31_7 ) , .ZN( us31_n464 ) );
  NOR4_X1 us31_U39 (.ZN( us31_n620 ) , .A1( us31_n656 ) , .A3( us31_n666 ) , .A4( us31_n682 ) , .A2( us31_n766 ) );
  NOR2_X1 us31_U390 (.A2( sa31_4 ) , .ZN( us31_n449 ) , .A1( us31_n848 ) );
  NOR2_X1 us31_U391 (.A2( sa31_4 ) , .A1( sa31_5 ) , .ZN( us31_n441 ) );
  NOR2_X1 us31_U392 (.A2( sa31_6 ) , .ZN( us31_n452 ) , .A1( us31_n858 ) );
  NOR2_X1 us31_U393 (.A2( sa31_2 ) , .A1( sa31_3 ) , .ZN( us31_n472 ) );
  NOR2_X1 us31_U394 (.A2( sa31_1 ) , .ZN( us31_n471 ) , .A1( us31_n826 ) );
  NOR2_X1 us31_U395 (.A2( sa31_0 ) , .ZN( us31_n454 ) , .A1( us31_n827 ) );
  NOR2_X1 us31_U396 (.A2( sa31_0 ) , .A1( sa31_1 ) , .ZN( us31_n462 ) );
  NOR2_X1 us31_U397 (.A2( sa31_3 ) , .ZN( us31_n455 ) , .A1( us31_n828 ) );
  NOR2_X1 us31_U398 (.A2( sa31_2 ) , .ZN( us31_n461 ) , .A1( us31_n829 ) );
  INV_X1 us31_U399 (.A( sa31_4 ) , .ZN( us31_n847 ) );
  NAND2_X1 us31_U4 (.A2( us31_n448 ) , .A1( us31_n464 ) , .ZN( us31_n815 ) );
  NOR4_X1 us31_U40 (.A4( us31_n609 ) , .A3( us31_n610 ) , .A2( us31_n611 ) , .A1( us31_n612 ) , .ZN( us31_n619 ) );
  INV_X1 us31_U400 (.A( sa31_6 ) , .ZN( us31_n849 ) );
  INV_X1 us31_U401 (.A( sa31_3 ) , .ZN( us31_n829 ) );
  INV_X1 us31_U402 (.A( sa31_1 ) , .ZN( us31_n827 ) );
  INV_X1 us31_U403 (.A( sa31_0 ) , .ZN( us31_n826 ) );
  INV_X1 us31_U404 (.A( sa31_2 ) , .ZN( us31_n828 ) );
  INV_X1 us31_U405 (.A( sa31_5 ) , .ZN( us31_n848 ) );
  INV_X1 us31_U406 (.A( sa31_7 ) , .ZN( us31_n858 ) );
  NAND2_X1 us31_U407 (.A2( us31_n461 ) , .A1( us31_n471 ) , .ZN( us31_n697 ) );
  OAI22_X1 us31_U408 (.ZN( us31_n588 ) , .A2( us31_n747 ) , .B2( us31_n762 ) , .A1( us31_n763 ) , .B1( us31_n784 ) );
  AOI21_X1 us31_U409 (.ZN( us31_n592 ) , .B1( us31_n728 ) , .B2( us31_n784 ) , .A( us31_n790 ) );
  NOR4_X1 us31_U41 (.A4( us31_n614 ) , .A3( us31_n615 ) , .A2( us31_n616 ) , .A1( us31_n617 ) , .ZN( us31_n618 ) );
  NAND2_X1 us31_U410 (.A1( us31_n729 ) , .A2( us31_n784 ) , .ZN( us31_n811 ) );
  AOI21_X1 us31_U411 (.ZN( us31_n623 ) , .B1( us31_n699 ) , .A( us31_n779 ) , .B2( us31_n784 ) );
  OAI22_X1 us31_U412 (.ZN( us31_n681 ) , .A1( us31_n699 ) , .A2( us31_n730 ) , .B2( us31_n784 ) , .B1( us31_n817 ) );
  AOI21_X1 us31_U413 (.ZN( us31_n648 ) , .A( us31_n762 ) , .B2( us31_n784 ) , .B1( us31_n792 ) );
  OAI21_X1 us31_U414 (.A( us31_n613 ) , .ZN( us31_n616 ) , .B1( us31_n625 ) , .B2( us31_n784 ) );
  OAI222_X1 us31_U415 (.A2( us31_n669 ) , .ZN( us31_n674 ) , .B1( us31_n747 ) , .B2( us31_n784 ) , .C2( us31_n788 ) , .C1( us31_n815 ) , .A1( us31_n817 ) );
  NOR2_X1 us31_U416 (.ZN( us31_n610 ) , .A1( us31_n784 ) , .A2( us31_n816 ) );
  NOR2_X1 us31_U417 (.ZN( us31_n651 ) , .A1( us31_n784 ) , .A2( us31_n788 ) );
  NOR2_X1 us31_U418 (.ZN( us31_n553 ) , .A2( us31_n744 ) , .A1( us31_n784 ) );
  NOR2_X1 us31_U419 (.ZN( us31_n600 ) , .A2( us31_n697 ) , .A1( us31_n784 ) );
  NOR4_X1 us31_U42 (.A4( us31_n514 ) , .A3( us31_n515 ) , .A2( us31_n516 ) , .A1( us31_n517 ) , .ZN( us31_n524 ) );
  INV_X1 us31_U420 (.A( us31_n784 ) , .ZN( us31_n861 ) );
  AND2_X1 us31_U421 (.ZN( us31_n438 ) , .A2( us31_n831 ) , .A1( us31_n854 ) );
  AND2_X1 us31_U422 (.ZN( us31_n439 ) , .A2( us31_n843 ) , .A1( us31_n861 ) );
  NOR3_X1 us31_U423 (.A1( us31_n438 ) , .A2( us31_n439 ) , .A3( us31_n576 ) , .ZN( us31_n587 ) );
  INV_X1 us31_U424 (.A( us31_n812 ) , .ZN( us31_n854 ) );
  INV_X1 us31_U425 (.A( us31_n803 ) , .ZN( us31_n843 ) );
  AOI21_X1 us31_U426 (.ZN( us31_n576 ) , .B2( us31_n724 ) , .B1( us31_n748 ) , .A( us31_n785 ) );
  OAI221_X1 us31_U427 (.A( us31_n783 ) , .C2( us31_n784 ) , .B2( us31_n785 ) , .B1( us31_n786 ) , .ZN( us31_n796 ) , .C1( us31_n813 ) );
  AOI21_X1 us31_U428 (.ZN( us31_n500 ) , .A( us31_n697 ) , .B1( us31_n708 ) , .B2( us31_n786 ) );
  OAI221_X1 us31_U429 (.A( us31_n696 ) , .ZN( us31_n703 ) , .C2( us31_n784 ) , .C1( us31_n785 ) , .B1( us31_n786 ) , .B2( us31_n806 ) );
  AOI222_X1 us31_U43 (.ZN( us31_n525 ) , .A1( us31_n834 ) , .B2( us31_n837 ) , .C1( us31_n844 ) , .C2( us31_n850 ) , .A2( us31_n852 ) , .B1( us31_n866 ) );
  OAI22_X1 us31_U430 (.ZN( us31_n590 ) , .B1( us31_n730 ) , .B2( us31_n749 ) , .A2( us31_n786 ) , .A1( us31_n803 ) );
  NAND2_X1 us31_U431 (.A2( us31_n749 ) , .A1( us31_n786 ) , .ZN( us31_n809 ) );
  NOR2_X1 us31_U432 (.ZN( us31_n612 ) , .A1( us31_n779 ) , .A2( us31_n786 ) );
  OAI222_X1 us31_U433 (.ZN( us31_n617 ) , .B1( us31_n697 ) , .C1( us31_n724 ) , .C2( us31_n747 ) , .B2( us31_n786 ) , .A2( us31_n792 ) , .A1( us31_n816 ) );
  NOR2_X1 us31_U434 (.ZN( us31_n653 ) , .A1( us31_n762 ) , .A2( us31_n786 ) );
  NOR2_X1 us31_U435 (.ZN( us31_n554 ) , .A1( us31_n786 ) , .A2( us31_n813 ) );
  NOR2_X1 us31_U436 (.ZN( us31_n717 ) , .A2( us31_n744 ) , .A1( us31_n786 ) );
  NAND3_X1 us31_U437 (.ZN( sa32_sr_6 ) , .A3( us31_n797 ) , .A2( us31_n798 ) , .A1( us31_n799 ) );
  NAND3_X1 us31_U438 (.ZN( sa32_sr_5 ) , .A3( us31_n758 ) , .A2( us31_n759 ) , .A1( us31_n760 ) );
  NAND3_X1 us31_U439 (.ZN( sa32_sr_4 ) , .A3( us31_n738 ) , .A2( us31_n739 ) , .A1( us31_n740 ) );
  NOR4_X1 us31_U44 (.A3( us31_n521 ) , .A1( us31_n522 ) , .ZN( us31_n523 ) , .A2( us31_n673 ) , .A4( us31_n769 ) );
  NAND3_X1 us31_U440 (.A3( us31_n675 ) , .A2( us31_n676 ) , .A1( us31_n677 ) , .ZN( us31_n807 ) );
  NAND3_X1 us31_U441 (.ZN( us31_n638 ) , .A3( us31_n708 ) , .A2( us31_n724 ) , .A1( us31_n792 ) );
  NAND3_X1 us31_U442 (.A3( us31_n618 ) , .A2( us31_n619 ) , .A1( us31_n620 ) , .ZN( us31_n725 ) );
  NAND3_X1 us31_U443 (.A3( us31_n585 ) , .A2( us31_n586 ) , .A1( us31_n587 ) , .ZN( us31_n621 ) );
  NAND3_X1 us31_U444 (.ZN( us31_n565 ) , .A3( us31_n680 ) , .A2( us31_n750 ) , .A1( us31_n785 ) );
  NAND3_X1 us31_U445 (.A3( us31_n523 ) , .A2( us31_n524 ) , .A1( us31_n525 ) , .ZN( us31_n742 ) );
  NAND3_X1 us31_U446 (.A3( us31_n512 ) , .A1( us31_n513 ) , .ZN( us31_n608 ) , .A2( us31_n871 ) );
  NAND3_X1 us31_U447 (.A3( us31_n467 ) , .A2( us31_n468 ) , .A1( us31_n469 ) , .ZN( us31_n777 ) );
  NOR2_X1 us31_U448 (.ZN( us31_n701 ) , .A2( us31_n786 ) , .A1( us31_n817 ) );
  NOR2_X1 us31_U449 (.A1( us31_n730 ) , .ZN( us31_n765 ) , .A2( us31_n786 ) );
  AOI221_X1 us31_U45 (.A( us31_n781 ) , .ZN( us31_n798 ) , .C2( us31_n837 ) , .B2( us31_n838 ) , .B1( us31_n865 ) , .C1( us31_n866 ) );
  NOR4_X1 us31_U46 (.A4( us31_n793 ) , .A3( us31_n794 ) , .A2( us31_n795 ) , .A1( us31_n796 ) , .ZN( us31_n797 ) );
  NOR4_X1 us31_U47 (.A4( us31_n776 ) , .A3( us31_n777 ) , .A1( us31_n778 ) , .ZN( us31_n799 ) , .A2( us31_n801 ) );
  NOR4_X1 us31_U48 (.A3( us31_n755 ) , .A2( us31_n756 ) , .A1( us31_n757 ) , .ZN( us31_n758 ) , .A4( us31_n869 ) );
  AOI211_X1 us31_U49 (.B( us31_n745 ) , .A( us31_n746 ) , .ZN( us31_n759 ) , .C1( us31_n832 ) , .C2( us31_n853 ) );
  NAND2_X1 us31_U5 (.A1( us31_n441 ) , .A2( us31_n464 ) , .ZN( us31_n708 ) );
  NOR3_X1 us31_U50 (.A3( us31_n741 ) , .A2( us31_n742 ) , .A1( us31_n743 ) , .ZN( us31_n760 ) );
  NAND4_X1 us31_U51 (.ZN( sa32_sr_3 ) , .A4( us31_n704 ) , .A3( us31_n705 ) , .A2( us31_n706 ) , .A1( us31_n707 ) );
  NOR4_X1 us31_U52 (.A4( us31_n700 ) , .A3( us31_n701 ) , .A2( us31_n702 ) , .A1( us31_n703 ) , .ZN( us31_n704 ) );
  AOI211_X1 us31_U53 (.B( us31_n694 ) , .A( us31_n695 ) , .ZN( us31_n705 ) , .C2( us31_n831 ) , .C1( us31_n851 ) );
  NOR2_X1 us31_U54 (.ZN( us31_n707 ) , .A2( us31_n776 ) , .A1( us31_n800 ) );
  NOR2_X1 us31_U55 (.ZN( us31_n804 ) , .A1( us31_n854 ) , .A2( us31_n861 ) );
  NAND4_X1 us31_U56 (.ZN( sa32_sr_7 ) , .A4( us31_n822 ) , .A3( us31_n823 ) , .A2( us31_n824 ) , .A1( us31_n825 ) );
  NOR4_X1 us31_U57 (.A4( us31_n818 ) , .A3( us31_n819 ) , .A2( us31_n820 ) , .A1( us31_n821 ) , .ZN( us31_n822 ) );
  AOI222_X1 us31_U58 (.C2( us31_n809 ) , .B2( us31_n810 ) , .A2( us31_n811 ) , .ZN( us31_n823 ) , .C1( us31_n832 ) , .A1( us31_n839 ) , .B1( us31_n853 ) );
  AOI211_X1 us31_U59 (.B( us31_n807 ) , .A( us31_n808 ) , .ZN( us31_n824 ) , .C1( us31_n842 ) , .C2( us31_n850 ) );
  NAND2_X1 us31_U6 (.A2( us31_n441 ) , .A1( us31_n452 ) , .ZN( us31_n791 ) );
  NAND4_X1 us31_U60 (.ZN( sa32_sr_0 ) , .A4( us31_n501 ) , .A3( us31_n502 ) , .A2( us31_n503 ) , .A1( us31_n504 ) );
  AOI221_X1 us31_U61 (.A( us31_n497 ) , .ZN( us31_n502 ) , .B2( us31_n843 ) , .C1( us31_n846 ) , .C2( us31_n860 ) , .B1( us31_n862 ) );
  NOR4_X1 us31_U62 (.A4( us31_n498 ) , .A3( us31_n499 ) , .A2( us31_n500 ) , .ZN( us31_n501 ) , .A1( us31_n527 ) );
  AOI211_X1 us31_U63 (.A( us31_n496 ) , .ZN( us31_n503 ) , .B( us31_n802 ) , .C2( us31_n839 ) , .C1( us31_n851 ) );
  NAND4_X1 us31_U64 (.ZN( sa32_sr_1 ) , .A4( us31_n595 ) , .A3( us31_n596 ) , .A2( us31_n597 ) , .A1( us31_n598 ) );
  NOR4_X1 us31_U65 (.A4( us31_n591 ) , .A3( us31_n592 ) , .A2( us31_n593 ) , .A1( us31_n594 ) , .ZN( us31_n595 ) );
  AOI211_X1 us31_U66 (.B( us31_n589 ) , .A( us31_n590 ) , .ZN( us31_n596 ) , .C2( us31_n811 ) , .C1( us31_n833 ) );
  AOI211_X1 us31_U67 (.A( us31_n588 ) , .ZN( us31_n597 ) , .B( us31_n621 ) , .C1( us31_n845 ) , .C2( us31_n855 ) );
  NAND4_X1 us31_U68 (.ZN( sa32_sr_2 ) , .A4( us31_n643 ) , .A3( us31_n644 ) , .A2( us31_n645 ) , .A1( us31_n646 ) );
  AOI222_X1 us31_U69 (.B2( us31_n638 ) , .ZN( us31_n644 ) , .B1( us31_n841 ) , .A1( us31_n842 ) , .C2( us31_n846 ) , .C1( us31_n863 ) , .A2( us31_n865 ) );
  NAND2_X1 us31_U7 (.A2( us31_n471 ) , .A1( us31_n472 ) , .ZN( us31_n817 ) );
  NOR4_X1 us31_U70 (.A4( us31_n639 ) , .A3( us31_n640 ) , .A2( us31_n641 ) , .A1( us31_n642 ) , .ZN( us31_n643 ) );
  NOR3_X1 us31_U71 (.A2( us31_n607 ) , .A1( us31_n608 ) , .ZN( us31_n646 ) , .A3( us31_n722 ) );
  NOR2_X1 us31_U72 (.ZN( us31_n748 ) , .A1( us31_n861 ) , .A2( us31_n862 ) );
  NOR2_X1 us31_U73 (.ZN( us31_n625 ) , .A2( us31_n836 ) , .A1( us31_n839 ) );
  NAND4_X1 us31_U74 (.A4( us31_n603 ) , .A3( us31_n604 ) , .A2( us31_n605 ) , .A1( us31_n606 ) , .ZN( us31_n722 ) );
  NOR3_X1 us31_U75 (.A1( us31_n599 ) , .ZN( us31_n604 ) , .A3( us31_n663 ) , .A2( us31_n770 ) );
  NOR4_X1 us31_U76 (.A3( us31_n600 ) , .A2( us31_n601 ) , .A1( us31_n602 ) , .ZN( us31_n603 ) , .A4( us31_n655 ) );
  AOI222_X1 us31_U77 (.ZN( us31_n606 ) , .A1( us31_n830 ) , .C2( us31_n837 ) , .B1( us31_n842 ) , .A2( us31_n856 ) , .B2( us31_n861 ) , .C1( us31_n868 ) );
  NAND4_X1 us31_U78 (.A4( us31_n657 ) , .A3( us31_n658 ) , .A2( us31_n659 ) , .A1( us31_n660 ) , .ZN( us31_n800 ) );
  NOR3_X1 us31_U79 (.A3( us31_n648 ) , .A2( us31_n649 ) , .A1( us31_n650 ) , .ZN( us31_n659 ) );
  NOR3_X1 us31_U8 (.ZN( us31_n598 ) , .A1( us31_n608 ) , .A3( us31_n723 ) , .A2( us31_n742 ) );
  NOR3_X1 us31_U80 (.A3( us31_n651 ) , .A2( us31_n652 ) , .A1( us31_n653 ) , .ZN( us31_n658 ) );
  NOR3_X1 us31_U81 (.A3( us31_n654 ) , .A2( us31_n655 ) , .A1( us31_n656 ) , .ZN( us31_n657 ) );
  NAND4_X1 us31_U82 (.A4( us31_n560 ) , .A3( us31_n561 ) , .A2( us31_n562 ) , .A1( us31_n563 ) , .ZN( us31_n607 ) );
  NOR4_X1 us31_U83 (.ZN( us31_n561 ) , .A1( us31_n653 ) , .A3( us31_n661 ) , .A4( us31_n685 ) , .A2( us31_n768 ) );
  NOR4_X1 us31_U84 (.A4( us31_n552 ) , .A3( us31_n553 ) , .A2( us31_n554 ) , .A1( us31_n555 ) , .ZN( us31_n562 ) );
  NOR4_X1 us31_U85 (.A4( us31_n556 ) , .A3( us31_n557 ) , .A2( us31_n558 ) , .A1( us31_n559 ) , .ZN( us31_n560 ) );
  NAND4_X1 us31_U86 (.A4( us31_n772 ) , .A3( us31_n773 ) , .A2( us31_n774 ) , .A1( us31_n775 ) , .ZN( us31_n801 ) );
  NOR3_X1 us31_U87 (.A3( us31_n765 ) , .A2( us31_n766 ) , .A1( us31_n767 ) , .ZN( us31_n773 ) );
  NOR4_X1 us31_U88 (.A4( us31_n768 ) , .A3( us31_n769 ) , .A2( us31_n770 ) , .A1( us31_n771 ) , .ZN( us31_n772 ) );
  AOI222_X1 us31_U89 (.ZN( us31_n775 ) , .A1( us31_n830 ) , .C1( us31_n834 ) , .B2( us31_n841 ) , .A2( us31_n850 ) , .B1( us31_n861 ) , .C2( us31_n873 ) );
  NOR3_X1 us31_U9 (.A3( us31_n800 ) , .A2( us31_n801 ) , .A1( us31_n802 ) , .ZN( us31_n825 ) );
  NOR4_X1 us31_U90 (.A4( us31_n661 ) , .A3( us31_n662 ) , .A2( us31_n663 ) , .A1( us31_n664 ) , .ZN( us31_n677 ) );
  NOR4_X1 us31_U91 (.A4( us31_n665 ) , .A3( us31_n666 ) , .A2( us31_n667 ) , .A1( us31_n668 ) , .ZN( us31_n676 ) );
  NOR4_X1 us31_U92 (.A3( us31_n673 ) , .A1( us31_n674 ) , .ZN( us31_n675 ) , .A4( us31_n715 ) , .A2( us31_n859 ) );
  NOR2_X1 us31_U93 (.ZN( us31_n761 ) , .A1( us31_n833 ) , .A2( us31_n834 ) );
  AOI222_X1 us31_U94 (.ZN( us31_n513 ) , .C1( us31_n832 ) , .B2( us31_n837 ) , .A2( us31_n843 ) , .C2( us31_n862 ) , .B1( us31_n863 ) , .A1( us31_n866 ) );
  NOR4_X1 us31_U95 (.A4( us31_n509 ) , .A2( us31_n510 ) , .A1( us31_n511 ) , .ZN( us31_n512 ) , .A3( us31_n670 ) );
  INV_X1 us31_U96 (.A( us31_n505 ) , .ZN( us31_n871 ) );
  NAND4_X1 us31_U97 (.A4( us31_n456 ) , .A3( us31_n457 ) , .A2( us31_n458 ) , .A1( us31_n459 ) , .ZN( us31_n679 ) );
  NOR3_X1 us31_U98 (.ZN( us31_n457 ) , .A3( us31_n530 ) , .A1( us31_n555 ) , .A2( us31_n570 ) );
  AOI221_X1 us31_U99 (.A( us31_n450 ) , .ZN( us31_n459 ) , .C2( us31_n753 ) , .B1( us31_n832 ) , .C1( us31_n842 ) , .B2( us31_n861 ) );
endmodule

module aes_aes_die_2 ( sa01_0, sa01_1, sa01_2, sa01_3, sa01_4, sa01_5, sa01_6, sa01_7, sa10_0, 
       sa10_1, sa10_2, sa10_3, sa10_4, sa10_5, sa10_6, sa10_7, sa11_0, sa11_1, 
       sa11_2, sa11_3, sa11_4, sa11_5, sa11_6, sa11_7, sa13_0, sa13_1, sa13_2, 
       sa13_3, sa13_4, sa13_5, sa13_6, sa13_7, sa20_0, sa20_1, sa20_2, sa20_3, 
       sa20_4, sa20_5, sa20_6, sa20_7, sa33_0, sa33_1, sa33_2, sa33_3, sa33_4, 
       sa33_5, sa33_6, sa33_7, sa01_sr_0, sa01_sr_1, sa01_sr_2, sa01_sr_3, sa01_sr_4, sa01_sr_5, sa01_sr_6, sa01_sr_7, sa10_sr_0, 
        sa10_sr_1, sa10_sr_2, sa10_sr_3, sa10_sr_4, sa10_sr_5, sa10_sr_6, sa10_sr_7, sa12_sr_0, sa12_sr_1, 
        sa12_sr_2, sa12_sr_3, sa12_sr_4, sa12_sr_5, sa12_sr_6, sa12_sr_7, sa13_sr_0, sa13_sr_1, sa13_sr_2, 
        sa13_sr_3, sa13_sr_4, sa13_sr_5, sa13_sr_6, sa13_sr_7, sa22_sr_0, sa22_sr_1, sa22_sr_2, sa22_sr_3, 
        sa22_sr_4, sa22_sr_5, sa22_sr_6, sa22_sr_7, sa30_sr_0, sa30_sr_1, sa30_sr_2, sa30_sr_3, sa30_sr_4, 
        sa30_sr_5, sa30_sr_6, sa30_sr_7 );
  input sa01_0, sa01_1, sa01_2, sa01_3, sa01_4, sa01_5, sa01_6, sa01_7, sa10_0, 
        sa10_1, sa10_2, sa10_3, sa10_4, sa10_5, sa10_6, sa10_7, sa11_0, sa11_1, 
        sa11_2, sa11_3, sa11_4, sa11_5, sa11_6, sa11_7, sa13_0, sa13_1, sa13_2, 
        sa13_3, sa13_4, sa13_5, sa13_6, sa13_7, sa20_0, sa20_1, sa20_2, sa20_3, 
        sa20_4, sa20_5, sa20_6, sa20_7, sa33_0, sa33_1, sa33_2, sa33_3, sa33_4, 
        sa33_5, sa33_6, sa33_7;
  output sa01_sr_0, sa01_sr_1, sa01_sr_2, sa01_sr_3, sa01_sr_4, sa01_sr_5, sa01_sr_6, sa01_sr_7, sa10_sr_0, 
        sa10_sr_1, sa10_sr_2, sa10_sr_3, sa10_sr_4, sa10_sr_5, sa10_sr_6, sa10_sr_7, sa12_sr_0, sa12_sr_1, 
        sa12_sr_2, sa12_sr_3, sa12_sr_4, sa12_sr_5, sa12_sr_6, sa12_sr_7, sa13_sr_0, sa13_sr_1, sa13_sr_2, 
        sa13_sr_3, sa13_sr_4, sa13_sr_5, sa13_sr_6, sa13_sr_7, sa22_sr_0, sa22_sr_1, sa22_sr_2, sa22_sr_3, 
        sa22_sr_4, sa22_sr_5, sa22_sr_6, sa22_sr_7, sa30_sr_0, sa30_sr_1, sa30_sr_2, sa30_sr_3, sa30_sr_4, 
        sa30_sr_5, sa30_sr_6, sa30_sr_7;
  wire us01_n438, us01_n439, us01_n440, us01_n441, us01_n442, us01_n443, us01_n444, us01_n445, us01_n446, 
       us01_n447, us01_n448, us01_n449, us01_n450, us01_n451, us01_n452, us01_n453, us01_n454, us01_n455, 
       us01_n456, us01_n457, us01_n458, us01_n459, us01_n460, us01_n461, us01_n462, us01_n463, us01_n464, 
       us01_n465, us01_n466, us01_n467, us01_n468, us01_n469, us01_n470, us01_n471, us01_n472, us01_n473, 
       us01_n474, us01_n475, us01_n476, us01_n477, us01_n478, us01_n479, us01_n480, us01_n481, us01_n482, 
       us01_n483, us01_n484, us01_n485, us01_n486, us01_n487, us01_n488, us01_n489, us01_n490, us01_n491, 
       us01_n492, us01_n493, us01_n494, us01_n495, us01_n496, us01_n497, us01_n498, us01_n499, us01_n500, 
       us01_n501, us01_n502, us01_n503, us01_n504, us01_n505, us01_n506, us01_n507, us01_n508, us01_n509, 
       us01_n510, us01_n511, us01_n512, us01_n513, us01_n514, us01_n515, us01_n516, us01_n517, us01_n518, 
       us01_n519, us01_n520, us01_n521, us01_n522, us01_n523, us01_n524, us01_n525, us01_n526, us01_n527, 
       us01_n528, us01_n529, us01_n530, us01_n531, us01_n532, us01_n533, us01_n534, us01_n535, us01_n536, 
       us01_n537, us01_n538, us01_n539, us01_n540, us01_n541, us01_n542, us01_n543, us01_n544, us01_n545, 
       us01_n546, us01_n547, us01_n548, us01_n549, us01_n550, us01_n551, us01_n552, us01_n553, us01_n554, 
       us01_n555, us01_n556, us01_n557, us01_n558, us01_n559, us01_n560, us01_n561, us01_n562, us01_n563, 
       us01_n564, us01_n565, us01_n566, us01_n567, us01_n568, us01_n569, us01_n570, us01_n571, us01_n572, 
       us01_n573, us01_n574, us01_n575, us01_n576, us01_n577, us01_n578, us01_n579, us01_n580, us01_n581, 
       us01_n582, us01_n583, us01_n584, us01_n585, us01_n586, us01_n587, us01_n588, us01_n589, us01_n590, 
       us01_n591, us01_n592, us01_n593, us01_n594, us01_n595, us01_n596, us01_n597, us01_n598, us01_n599, 
       us01_n600, us01_n601, us01_n602, us01_n603, us01_n604, us01_n605, us01_n606, us01_n607, us01_n608, 
       us01_n609, us01_n610, us01_n611, us01_n612, us01_n613, us01_n614, us01_n615, us01_n616, us01_n617, 
       us01_n618, us01_n619, us01_n620, us01_n621, us01_n622, us01_n623, us01_n624, us01_n625, us01_n626, 
       us01_n627, us01_n628, us01_n629, us01_n630, us01_n631, us01_n632, us01_n633, us01_n634, us01_n635, 
       us01_n636, us01_n637, us01_n638, us01_n639, us01_n640, us01_n641, us01_n642, us01_n643, us01_n644, 
       us01_n645, us01_n646, us01_n647, us01_n648, us01_n649, us01_n650, us01_n651, us01_n652, us01_n653, 
       us01_n654, us01_n655, us01_n656, us01_n657, us01_n658, us01_n659, us01_n660, us01_n661, us01_n662, 
       us01_n663, us01_n664, us01_n665, us01_n666, us01_n667, us01_n668, us01_n669, us01_n670, us01_n671, 
       us01_n672, us01_n673, us01_n674, us01_n675, us01_n676, us01_n677, us01_n678, us01_n679, us01_n680, 
       us01_n681, us01_n682, us01_n683, us01_n684, us01_n685, us01_n686, us01_n687, us01_n688, us01_n689, 
       us01_n690, us01_n691, us01_n692, us01_n693, us01_n694, us01_n695, us01_n696, us01_n697, us01_n698, 
       us01_n699, us01_n700, us01_n701, us01_n702, us01_n703, us01_n704, us01_n705, us01_n706, us01_n707, 
       us01_n708, us01_n709, us01_n710, us01_n711, us01_n712, us01_n713, us01_n714, us01_n715, us01_n716, 
       us01_n717, us01_n718, us01_n719, us01_n720, us01_n721, us01_n722, us01_n723, us01_n724, us01_n725, 
       us01_n726, us01_n727, us01_n728, us01_n729, us01_n730, us01_n731, us01_n732, us01_n733, us01_n734, 
       us01_n735, us01_n736, us01_n737, us01_n738, us01_n739, us01_n740, us01_n741, us01_n742, us01_n743, 
       us01_n744, us01_n745, us01_n746, us01_n747, us01_n748, us01_n749, us01_n750, us01_n751, us01_n752, 
       us01_n753, us01_n754, us01_n755, us01_n756, us01_n757, us01_n758, us01_n759, us01_n760, us01_n761, 
       us01_n762, us01_n763, us01_n764, us01_n765, us01_n766, us01_n767, us01_n768, us01_n769, us01_n770, 
       us01_n771, us01_n772, us01_n773, us01_n774, us01_n775, us01_n776, us01_n777, us01_n778, us01_n779, 
       us01_n780, us01_n781, us01_n782, us01_n783, us01_n784, us01_n785, us01_n786, us01_n787, us01_n788, 
       us01_n789, us01_n790, us01_n791, us01_n792, us01_n793, us01_n794, us01_n795, us01_n796, us01_n797, 
       us01_n798, us01_n799, us01_n800, us01_n801, us01_n802, us01_n803, us01_n804, us01_n805, us01_n806, 
       us01_n807, us01_n808, us01_n809, us01_n810, us01_n811, us01_n812, us01_n813, us01_n814, us01_n815, 
       us01_n816, us01_n817, us01_n818, us01_n819, us01_n820, us01_n821, us01_n822, us01_n823, us01_n824, 
       us01_n825, us01_n826, us01_n827, us01_n828, us01_n829, us01_n830, us01_n831, us01_n832, us01_n833, 
       us01_n834, us01_n835, us01_n836, us01_n837, us01_n838, us01_n839, us01_n840, us01_n841, us01_n842, 
       us01_n843, us01_n844, us01_n845, us01_n846, us01_n847, us01_n848, us01_n849, us01_n850, us01_n851, 
       us01_n852, us01_n853, us01_n854, us01_n855, us01_n856, us01_n857, us01_n858, us01_n859, us01_n860, 
       us01_n861, us01_n862, us01_n863, us01_n864, us01_n865, us01_n866, us01_n867, us01_n868, us01_n869, 
       us01_n870, us01_n871, us01_n872, us01_n873, us01_n874, us10_n438, us10_n439, us10_n440, us10_n441, 
       us10_n442, us10_n443, us10_n444, us10_n445, us10_n446, us10_n447, us10_n448, us10_n449, us10_n450, 
       us10_n451, us10_n452, us10_n453, us10_n454, us10_n455, us10_n456, us10_n457, us10_n458, us10_n459, 
       us10_n460, us10_n461, us10_n462, us10_n463, us10_n464, us10_n465, us10_n466, us10_n467, us10_n468, 
       us10_n469, us10_n470, us10_n471, us10_n472, us10_n473, us10_n474, us10_n475, us10_n476, us10_n477, 
       us10_n478, us10_n479, us10_n480, us10_n481, us10_n482, us10_n483, us10_n484, us10_n485, us10_n486, 
       us10_n487, us10_n488, us10_n489, us10_n490, us10_n491, us10_n492, us10_n493, us10_n494, us10_n495, 
       us10_n496, us10_n497, us10_n498, us10_n499, us10_n500, us10_n501, us10_n502, us10_n503, us10_n504, 
       us10_n505, us10_n506, us10_n507, us10_n508, us10_n509, us10_n510, us10_n511, us10_n512, us10_n513, 
       us10_n514, us10_n515, us10_n516, us10_n517, us10_n518, us10_n519, us10_n520, us10_n521, us10_n522, 
       us10_n523, us10_n524, us10_n525, us10_n526, us10_n527, us10_n528, us10_n529, us10_n530, us10_n531, 
       us10_n532, us10_n533, us10_n534, us10_n535, us10_n536, us10_n537, us10_n538, us10_n539, us10_n540, 
       us10_n541, us10_n542, us10_n543, us10_n544, us10_n545, us10_n546, us10_n547, us10_n548, us10_n549, 
       us10_n550, us10_n551, us10_n552, us10_n553, us10_n554, us10_n555, us10_n556, us10_n557, us10_n558, 
       us10_n559, us10_n560, us10_n561, us10_n562, us10_n563, us10_n564, us10_n565, us10_n566, us10_n567, 
       us10_n568, us10_n569, us10_n570, us10_n571, us10_n572, us10_n573, us10_n574, us10_n575, us10_n576, 
       us10_n577, us10_n578, us10_n579, us10_n580, us10_n581, us10_n582, us10_n583, us10_n584, us10_n585, 
       us10_n586, us10_n587, us10_n588, us10_n589, us10_n590, us10_n591, us10_n592, us10_n593, us10_n594, 
       us10_n595, us10_n596, us10_n597, us10_n598, us10_n599, us10_n600, us10_n601, us10_n602, us10_n603, 
       us10_n604, us10_n605, us10_n606, us10_n607, us10_n608, us10_n609, us10_n610, us10_n611, us10_n612, 
       us10_n613, us10_n614, us10_n615, us10_n616, us10_n617, us10_n618, us10_n619, us10_n620, us10_n621, 
       us10_n622, us10_n623, us10_n624, us10_n625, us10_n626, us10_n627, us10_n628, us10_n629, us10_n630, 
       us10_n631, us10_n632, us10_n633, us10_n634, us10_n635, us10_n636, us10_n637, us10_n638, us10_n639, 
       us10_n640, us10_n641, us10_n642, us10_n643, us10_n644, us10_n645, us10_n646, us10_n647, us10_n648, 
       us10_n649, us10_n650, us10_n651, us10_n652, us10_n653, us10_n654, us10_n655, us10_n656, us10_n657, 
       us10_n658, us10_n659, us10_n660, us10_n661, us10_n662, us10_n663, us10_n664, us10_n665, us10_n666, 
       us10_n667, us10_n668, us10_n669, us10_n670, us10_n671, us10_n672, us10_n673, us10_n674, us10_n675, 
       us10_n676, us10_n677, us10_n678, us10_n679, us10_n680, us10_n681, us10_n682, us10_n683, us10_n684, 
       us10_n685, us10_n686, us10_n687, us10_n688, us10_n689, us10_n690, us10_n691, us10_n692, us10_n693, 
       us10_n694, us10_n695, us10_n696, us10_n697, us10_n698, us10_n699, us10_n700, us10_n701, us10_n702, 
       us10_n703, us10_n704, us10_n705, us10_n706, us10_n707, us10_n708, us10_n709, us10_n710, us10_n711, 
       us10_n712, us10_n713, us10_n714, us10_n715, us10_n716, us10_n717, us10_n718, us10_n719, us10_n720, 
       us10_n721, us10_n722, us10_n723, us10_n724, us10_n725, us10_n726, us10_n727, us10_n728, us10_n729, 
       us10_n730, us10_n731, us10_n732, us10_n733, us10_n734, us10_n735, us10_n736, us10_n737, us10_n738, 
       us10_n739, us10_n740, us10_n741, us10_n742, us10_n743, us10_n744, us10_n745, us10_n746, us10_n747, 
       us10_n748, us10_n749, us10_n750, us10_n751, us10_n752, us10_n753, us10_n754, us10_n755, us10_n756, 
       us10_n757, us10_n758, us10_n759, us10_n760, us10_n761, us10_n762, us10_n763, us10_n764, us10_n765, 
       us10_n766, us10_n767, us10_n768, us10_n769, us10_n770, us10_n771, us10_n772, us10_n773, us10_n774, 
       us10_n775, us10_n776, us10_n777, us10_n778, us10_n779, us10_n780, us10_n781, us10_n782, us10_n783, 
       us10_n784, us10_n785, us10_n786, us10_n787, us10_n788, us10_n789, us10_n790, us10_n791, us10_n792, 
       us10_n793, us10_n794, us10_n795, us10_n796, us10_n797, us10_n798, us10_n799, us10_n800, us10_n801, 
       us10_n802, us10_n803, us10_n804, us10_n805, us10_n806, us10_n807, us10_n808, us10_n809, us10_n810, 
       us10_n811, us10_n812, us10_n813, us10_n814, us10_n815, us10_n816, us10_n817, us10_n818, us10_n819, 
       us10_n820, us10_n821, us10_n822, us10_n823, us10_n824, us10_n825, us10_n826, us10_n827, us10_n828, 
       us10_n829, us10_n830, us10_n831, us10_n832, us10_n833, us10_n834, us10_n835, us10_n836, us10_n837, 
       us10_n838, us10_n839, us10_n840, us10_n841, us10_n842, us10_n843, us10_n844, us10_n845, us10_n846, 
       us10_n847, us10_n848, us10_n849, us10_n850, us10_n851, us10_n852, us10_n853, us10_n854, us10_n855, 
       us10_n856, us10_n857, us10_n858, us10_n859, us10_n860, us10_n861, us10_n862, us10_n863, us10_n864, 
       us10_n865, us10_n866, us10_n867, us10_n868, us10_n869, us10_n870, us10_n871, us10_n872, us10_n873, 
       us10_n874, us10_n875, us10_n876, us11_n438, us11_n439, us11_n440, us11_n441, us11_n442, us11_n443, 
       us11_n444, us11_n445, us11_n446, us11_n447, us11_n448, us11_n449, us11_n450, us11_n451, us11_n452, 
       us11_n453, us11_n454, us11_n455, us11_n456, us11_n457, us11_n458, us11_n459, us11_n460, us11_n461, 
       us11_n462, us11_n463, us11_n464, us11_n465, us11_n466, us11_n467, us11_n468, us11_n469, us11_n470, 
       us11_n471, us11_n472, us11_n473, us11_n474, us11_n475, us11_n476, us11_n477, us11_n478, us11_n479, 
       us11_n480, us11_n481, us11_n482, us11_n483, us11_n484, us11_n485, us11_n486, us11_n487, us11_n488, 
       us11_n489, us11_n490, us11_n491, us11_n492, us11_n493, us11_n494, us11_n495, us11_n496, us11_n497, 
       us11_n498, us11_n499, us11_n500, us11_n501, us11_n502, us11_n503, us11_n504, us11_n505, us11_n506, 
       us11_n507, us11_n508, us11_n509, us11_n510, us11_n511, us11_n512, us11_n513, us11_n514, us11_n515, 
       us11_n516, us11_n517, us11_n518, us11_n519, us11_n520, us11_n521, us11_n522, us11_n523, us11_n524, 
       us11_n525, us11_n526, us11_n527, us11_n528, us11_n529, us11_n530, us11_n531, us11_n532, us11_n533, 
       us11_n534, us11_n535, us11_n536, us11_n537, us11_n538, us11_n539, us11_n540, us11_n541, us11_n542, 
       us11_n543, us11_n544, us11_n545, us11_n546, us11_n547, us11_n548, us11_n549, us11_n550, us11_n551, 
       us11_n552, us11_n553, us11_n554, us11_n555, us11_n556, us11_n557, us11_n558, us11_n559, us11_n560, 
       us11_n561, us11_n562, us11_n563, us11_n564, us11_n565, us11_n566, us11_n567, us11_n568, us11_n569, 
       us11_n570, us11_n571, us11_n572, us11_n573, us11_n574, us11_n575, us11_n576, us11_n577, us11_n578, 
       us11_n579, us11_n580, us11_n581, us11_n582, us11_n583, us11_n584, us11_n585, us11_n586, us11_n587, 
       us11_n588, us11_n589, us11_n590, us11_n591, us11_n592, us11_n593, us11_n594, us11_n595, us11_n596, 
       us11_n597, us11_n598, us11_n599, us11_n600, us11_n601, us11_n602, us11_n603, us11_n604, us11_n605, 
       us11_n606, us11_n607, us11_n608, us11_n609, us11_n610, us11_n611, us11_n612, us11_n613, us11_n614, 
       us11_n615, us11_n616, us11_n617, us11_n618, us11_n619, us11_n620, us11_n621, us11_n622, us11_n623, 
       us11_n624, us11_n625, us11_n626, us11_n627, us11_n628, us11_n629, us11_n630, us11_n631, us11_n632, 
       us11_n633, us11_n634, us11_n635, us11_n636, us11_n637, us11_n638, us11_n639, us11_n640, us11_n641, 
       us11_n642, us11_n643, us11_n644, us11_n645, us11_n646, us11_n647, us11_n648, us11_n649, us11_n650, 
       us11_n651, us11_n652, us11_n653, us11_n654, us11_n655, us11_n656, us11_n657, us11_n658, us11_n659, 
       us11_n660, us11_n661, us11_n662, us11_n663, us11_n664, us11_n665, us11_n666, us11_n667, us11_n668, 
       us11_n669, us11_n670, us11_n671, us11_n672, us11_n673, us11_n674, us11_n675, us11_n676, us11_n677, 
       us11_n678, us11_n679, us11_n680, us11_n681, us11_n682, us11_n683, us11_n684, us11_n685, us11_n686, 
       us11_n687, us11_n688, us11_n689, us11_n690, us11_n691, us11_n692, us11_n693, us11_n694, us11_n695, 
       us11_n696, us11_n697, us11_n698, us11_n699, us11_n700, us11_n701, us11_n702, us11_n703, us11_n704, 
       us11_n705, us11_n706, us11_n707, us11_n708, us11_n709, us11_n710, us11_n711, us11_n712, us11_n713, 
       us11_n714, us11_n715, us11_n716, us11_n717, us11_n718, us11_n719, us11_n720, us11_n721, us11_n722, 
       us11_n723, us11_n724, us11_n725, us11_n726, us11_n727, us11_n728, us11_n729, us11_n730, us11_n731, 
       us11_n732, us11_n733, us11_n734, us11_n735, us11_n736, us11_n737, us11_n738, us11_n739, us11_n740, 
       us11_n741, us11_n742, us11_n743, us11_n744, us11_n745, us11_n746, us11_n747, us11_n748, us11_n749, 
       us11_n750, us11_n751, us11_n752, us11_n753, us11_n754, us11_n755, us11_n756, us11_n757, us11_n758, 
       us11_n759, us11_n760, us11_n761, us11_n762, us11_n763, us11_n764, us11_n765, us11_n766, us11_n767, 
       us11_n768, us11_n769, us11_n770, us11_n771, us11_n772, us11_n773, us11_n774, us11_n775, us11_n776, 
       us11_n777, us11_n778, us11_n779, us11_n780, us11_n781, us11_n782, us11_n783, us11_n784, us11_n785, 
       us11_n786, us11_n787, us11_n788, us11_n789, us11_n790, us11_n791, us11_n792, us11_n793, us11_n794, 
       us11_n795, us11_n796, us11_n797, us11_n798, us11_n799, us11_n800, us11_n801, us11_n802, us11_n803, 
       us11_n804, us11_n805, us11_n806, us11_n807, us11_n808, us11_n809, us11_n810, us11_n811, us11_n812, 
       us11_n813, us11_n814, us11_n815, us11_n816, us11_n817, us11_n818, us11_n819, us11_n820, us11_n821, 
       us11_n822, us11_n823, us11_n824, us11_n825, us11_n826, us11_n827, us11_n828, us11_n829, us11_n830, 
       us11_n831, us11_n832, us11_n833, us11_n834, us11_n835, us11_n836, us11_n837, us11_n838, us11_n839, 
       us11_n840, us11_n841, us11_n842, us11_n843, us11_n844, us11_n845, us11_n846, us11_n847, us11_n848, 
       us11_n849, us11_n850, us11_n851, us11_n852, us11_n853, us11_n854, us11_n855, us11_n856, us11_n857, 
       us11_n858, us11_n859, us11_n860, us11_n861, us11_n862, us11_n863, us11_n864, us11_n865, us11_n866, 
       us11_n867, us11_n868, us11_n869, us11_n870, us11_n871, us11_n872, us11_n873, us11_n874, us11_n875, 
       us11_n876, us13_n438, us13_n439, us13_n440, us13_n441, us13_n442, us13_n443, us13_n444, us13_n445, 
       us13_n446, us13_n447, us13_n448, us13_n449, us13_n450, us13_n451, us13_n452, us13_n453, us13_n454, 
       us13_n455, us13_n456, us13_n457, us13_n458, us13_n459, us13_n460, us13_n461, us13_n462, us13_n463, 
       us13_n464, us13_n465, us13_n466, us13_n467, us13_n468, us13_n469, us13_n470, us13_n471, us13_n472, 
       us13_n473, us13_n474, us13_n475, us13_n476, us13_n477, us13_n478, us13_n479, us13_n480, us13_n481, 
       us13_n482, us13_n483, us13_n484, us13_n485, us13_n486, us13_n487, us13_n488, us13_n489, us13_n490, 
       us13_n491, us13_n492, us13_n493, us13_n494, us13_n495, us13_n496, us13_n497, us13_n498, us13_n499, 
       us13_n500, us13_n501, us13_n502, us13_n503, us13_n504, us13_n505, us13_n506, us13_n507, us13_n508, 
       us13_n509, us13_n510, us13_n511, us13_n512, us13_n513, us13_n514, us13_n515, us13_n516, us13_n517, 
       us13_n518, us13_n519, us13_n520, us13_n521, us13_n522, us13_n523, us13_n524, us13_n525, us13_n526, 
       us13_n527, us13_n528, us13_n529, us13_n530, us13_n531, us13_n532, us13_n533, us13_n534, us13_n535, 
       us13_n536, us13_n537, us13_n538, us13_n539, us13_n540, us13_n541, us13_n542, us13_n543, us13_n544, 
       us13_n545, us13_n546, us13_n547, us13_n548, us13_n549, us13_n550, us13_n551, us13_n552, us13_n553, 
       us13_n554, us13_n555, us13_n556, us13_n557, us13_n558, us13_n559, us13_n560, us13_n561, us13_n562, 
       us13_n563, us13_n564, us13_n565, us13_n566, us13_n567, us13_n568, us13_n569, us13_n570, us13_n571, 
       us13_n572, us13_n573, us13_n574, us13_n575, us13_n576, us13_n577, us13_n578, us13_n579, us13_n580, 
       us13_n581, us13_n582, us13_n583, us13_n584, us13_n585, us13_n586, us13_n587, us13_n588, us13_n589, 
       us13_n590, us13_n591, us13_n592, us13_n593, us13_n594, us13_n595, us13_n596, us13_n597, us13_n598, 
       us13_n599, us13_n600, us13_n601, us13_n602, us13_n603, us13_n604, us13_n605, us13_n606, us13_n607, 
       us13_n608, us13_n609, us13_n610, us13_n611, us13_n612, us13_n613, us13_n614, us13_n615, us13_n616, 
       us13_n617, us13_n618, us13_n619, us13_n620, us13_n621, us13_n622, us13_n623, us13_n624, us13_n625, 
       us13_n626, us13_n627, us13_n628, us13_n629, us13_n630, us13_n631, us13_n632, us13_n633, us13_n634, 
       us13_n635, us13_n636, us13_n637, us13_n638, us13_n639, us13_n640, us13_n641, us13_n642, us13_n643, 
       us13_n644, us13_n645, us13_n646, us13_n647, us13_n648, us13_n649, us13_n650, us13_n651, us13_n652, 
       us13_n653, us13_n654, us13_n655, us13_n656, us13_n657, us13_n658, us13_n659, us13_n660, us13_n661, 
       us13_n662, us13_n663, us13_n664, us13_n665, us13_n666, us13_n667, us13_n668, us13_n669, us13_n670, 
       us13_n671, us13_n672, us13_n673, us13_n674, us13_n675, us13_n676, us13_n677, us13_n678, us13_n679, 
       us13_n680, us13_n681, us13_n682, us13_n683, us13_n684, us13_n685, us13_n686, us13_n687, us13_n688, 
       us13_n689, us13_n690, us13_n691, us13_n692, us13_n693, us13_n694, us13_n695, us13_n696, us13_n697, 
       us13_n698, us13_n699, us13_n700, us13_n701, us13_n702, us13_n703, us13_n704, us13_n705, us13_n706, 
       us13_n707, us13_n708, us13_n709, us13_n710, us13_n711, us13_n712, us13_n713, us13_n714, us13_n715, 
       us13_n716, us13_n717, us13_n718, us13_n719, us13_n720, us13_n721, us13_n722, us13_n723, us13_n724, 
       us13_n725, us13_n726, us13_n727, us13_n728, us13_n729, us13_n730, us13_n731, us13_n732, us13_n733, 
       us13_n734, us13_n735, us13_n736, us13_n737, us13_n738, us13_n739, us13_n740, us13_n741, us13_n742, 
       us13_n743, us13_n744, us13_n745, us13_n746, us13_n747, us13_n748, us13_n749, us13_n750, us13_n751, 
       us13_n752, us13_n753, us13_n754, us13_n755, us13_n756, us13_n757, us13_n758, us13_n759, us13_n760, 
       us13_n761, us13_n762, us13_n763, us13_n764, us13_n765, us13_n766, us13_n767, us13_n768, us13_n769, 
       us13_n770, us13_n771, us13_n772, us13_n773, us13_n774, us13_n775, us13_n776, us13_n777, us13_n778, 
       us13_n779, us13_n780, us13_n781, us13_n782, us13_n783, us13_n784, us13_n785, us13_n786, us13_n787, 
       us13_n788, us13_n789, us13_n790, us13_n791, us13_n792, us13_n793, us13_n794, us13_n795, us13_n796, 
       us13_n797, us13_n798, us13_n799, us13_n800, us13_n801, us13_n802, us13_n803, us13_n804, us13_n805, 
       us13_n806, us13_n807, us13_n808, us13_n809, us13_n810, us13_n811, us13_n812, us13_n813, us13_n814, 
       us13_n815, us13_n816, us13_n817, us13_n818, us13_n819, us13_n820, us13_n821, us13_n822, us13_n823, 
       us13_n824, us13_n825, us13_n826, us13_n827, us13_n828, us13_n829, us13_n830, us13_n831, us13_n832, 
       us13_n833, us13_n834, us13_n835, us13_n836, us13_n837, us13_n838, us13_n839, us13_n840, us13_n841, 
       us13_n842, us13_n843, us13_n844, us13_n845, us13_n846, us13_n847, us13_n848, us13_n849, us13_n850, 
       us13_n851, us13_n852, us13_n853, us13_n854, us13_n855, us13_n856, us13_n857, us13_n858, us13_n859, 
       us13_n860, us13_n861, us13_n862, us13_n863, us13_n864, us13_n865, us13_n866, us13_n867, us13_n868, 
       us13_n869, us13_n870, us13_n871, us13_n872, us13_n873, us13_n874, us13_n875, us13_n876, us20_n438, 
       us20_n439, us20_n440, us20_n441, us20_n442, us20_n443, us20_n444, us20_n445, us20_n446, us20_n447, 
       us20_n448, us20_n449, us20_n450, us20_n451, us20_n452, us20_n453, us20_n454, us20_n455, us20_n456, 
       us20_n457, us20_n458, us20_n459, us20_n460, us20_n461, us20_n462, us20_n463, us20_n464, us20_n465, 
       us20_n466, us20_n467, us20_n468, us20_n469, us20_n470, us20_n471, us20_n472, us20_n473, us20_n474, 
       us20_n475, us20_n476, us20_n477, us20_n478, us20_n479, us20_n480, us20_n481, us20_n482, us20_n483, 
       us20_n484, us20_n485, us20_n486, us20_n487, us20_n488, us20_n489, us20_n490, us20_n491, us20_n492, 
       us20_n493, us20_n494, us20_n495, us20_n496, us20_n497, us20_n498, us20_n499, us20_n500, us20_n501, 
       us20_n502, us20_n503, us20_n504, us20_n505, us20_n506, us20_n507, us20_n508, us20_n509, us20_n510, 
       us20_n511, us20_n512, us20_n513, us20_n514, us20_n515, us20_n516, us20_n517, us20_n518, us20_n519, 
       us20_n520, us20_n521, us20_n522, us20_n523, us20_n524, us20_n525, us20_n526, us20_n527, us20_n528, 
       us20_n529, us20_n530, us20_n531, us20_n532, us20_n533, us20_n534, us20_n535, us20_n536, us20_n537, 
       us20_n538, us20_n539, us20_n540, us20_n541, us20_n542, us20_n543, us20_n544, us20_n545, us20_n546, 
       us20_n547, us20_n548, us20_n549, us20_n550, us20_n551, us20_n552, us20_n553, us20_n554, us20_n555, 
       us20_n556, us20_n557, us20_n558, us20_n559, us20_n560, us20_n561, us20_n562, us20_n563, us20_n564, 
       us20_n565, us20_n566, us20_n567, us20_n568, us20_n569, us20_n570, us20_n571, us20_n572, us20_n573, 
       us20_n574, us20_n575, us20_n576, us20_n577, us20_n578, us20_n579, us20_n580, us20_n581, us20_n582, 
       us20_n583, us20_n584, us20_n585, us20_n586, us20_n587, us20_n588, us20_n589, us20_n590, us20_n591, 
       us20_n592, us20_n593, us20_n594, us20_n595, us20_n596, us20_n597, us20_n598, us20_n599, us20_n600, 
       us20_n601, us20_n602, us20_n603, us20_n604, us20_n605, us20_n606, us20_n607, us20_n608, us20_n609, 
       us20_n610, us20_n611, us20_n612, us20_n613, us20_n614, us20_n615, us20_n616, us20_n617, us20_n618, 
       us20_n619, us20_n620, us20_n621, us20_n622, us20_n623, us20_n624, us20_n625, us20_n626, us20_n627, 
       us20_n628, us20_n629, us20_n630, us20_n631, us20_n632, us20_n633, us20_n634, us20_n635, us20_n636, 
       us20_n637, us20_n638, us20_n639, us20_n640, us20_n641, us20_n642, us20_n643, us20_n644, us20_n645, 
       us20_n646, us20_n647, us20_n648, us20_n649, us20_n650, us20_n651, us20_n652, us20_n653, us20_n654, 
       us20_n655, us20_n656, us20_n657, us20_n658, us20_n659, us20_n660, us20_n661, us20_n662, us20_n663, 
       us20_n664, us20_n665, us20_n666, us20_n667, us20_n668, us20_n669, us20_n670, us20_n671, us20_n672, 
       us20_n673, us20_n674, us20_n675, us20_n676, us20_n677, us20_n678, us20_n679, us20_n680, us20_n681, 
       us20_n682, us20_n683, us20_n684, us20_n685, us20_n686, us20_n687, us20_n688, us20_n689, us20_n690, 
       us20_n691, us20_n692, us20_n693, us20_n694, us20_n695, us20_n696, us20_n697, us20_n698, us20_n699, 
       us20_n700, us20_n701, us20_n702, us20_n703, us20_n704, us20_n705, us20_n706, us20_n707, us20_n708, 
       us20_n709, us20_n710, us20_n711, us20_n712, us20_n713, us20_n714, us20_n715, us20_n716, us20_n717, 
       us20_n718, us20_n719, us20_n720, us20_n721, us20_n722, us20_n723, us20_n724, us20_n725, us20_n726, 
       us20_n727, us20_n728, us20_n729, us20_n730, us20_n731, us20_n732, us20_n733, us20_n734, us20_n735, 
       us20_n736, us20_n737, us20_n738, us20_n739, us20_n740, us20_n741, us20_n742, us20_n743, us20_n744, 
       us20_n745, us20_n746, us20_n747, us20_n748, us20_n749, us20_n750, us20_n751, us20_n752, us20_n753, 
       us20_n754, us20_n755, us20_n756, us20_n757, us20_n758, us20_n759, us20_n760, us20_n761, us20_n762, 
       us20_n763, us20_n764, us20_n765, us20_n766, us20_n767, us20_n768, us20_n769, us20_n770, us20_n771, 
       us20_n772, us20_n773, us20_n774, us20_n775, us20_n776, us20_n777, us20_n778, us20_n779, us20_n780, 
       us20_n781, us20_n782, us20_n783, us20_n784, us20_n785, us20_n786, us20_n787, us20_n788, us20_n789, 
       us20_n790, us20_n791, us20_n792, us20_n793, us20_n794, us20_n795, us20_n796, us20_n797, us20_n798, 
       us20_n799, us20_n800, us20_n801, us20_n802, us20_n803, us20_n804, us20_n805, us20_n806, us20_n807, 
       us20_n808, us20_n809, us20_n810, us20_n811, us20_n812, us20_n813, us20_n814, us20_n815, us20_n816, 
       us20_n817, us20_n818, us20_n819, us20_n820, us20_n821, us20_n822, us20_n823, us20_n824, us20_n825, 
       us20_n826, us20_n827, us20_n828, us20_n829, us20_n830, us20_n831, us20_n832, us20_n833, us20_n834, 
       us20_n835, us20_n836, us20_n837, us20_n838, us20_n839, us20_n840, us20_n841, us20_n842, us20_n843, 
       us20_n844, us20_n845, us20_n846, us20_n847, us20_n848, us20_n849, us20_n850, us20_n851, us20_n852, 
       us20_n853, us20_n854, us20_n855, us20_n856, us20_n857, us20_n858, us20_n859, us20_n860, us20_n861, 
       us20_n862, us20_n863, us20_n864, us20_n865, us20_n866, us20_n867, us20_n868, us20_n869, us20_n870, 
       us20_n871, us20_n872, us20_n873, us20_n874, us20_n875, us20_n876, us33_n438, us33_n439, us33_n440, 
       us33_n441, us33_n442, us33_n443, us33_n444, us33_n445, us33_n446, us33_n447, us33_n448, us33_n449, 
       us33_n450, us33_n451, us33_n452, us33_n453, us33_n454, us33_n455, us33_n456, us33_n457, us33_n458, 
       us33_n459, us33_n460, us33_n461, us33_n462, us33_n463, us33_n464, us33_n465, us33_n466, us33_n467, 
       us33_n468, us33_n469, us33_n470, us33_n471, us33_n472, us33_n473, us33_n474, us33_n475, us33_n476, 
       us33_n477, us33_n478, us33_n479, us33_n480, us33_n481, us33_n482, us33_n483, us33_n484, us33_n485, 
       us33_n486, us33_n487, us33_n488, us33_n489, us33_n490, us33_n491, us33_n492, us33_n493, us33_n494, 
       us33_n495, us33_n496, us33_n497, us33_n498, us33_n499, us33_n500, us33_n501, us33_n502, us33_n503, 
       us33_n504, us33_n505, us33_n506, us33_n507, us33_n508, us33_n509, us33_n510, us33_n511, us33_n512, 
       us33_n513, us33_n514, us33_n515, us33_n516, us33_n517, us33_n518, us33_n519, us33_n520, us33_n521, 
       us33_n522, us33_n523, us33_n524, us33_n525, us33_n526, us33_n527, us33_n528, us33_n529, us33_n530, 
       us33_n531, us33_n532, us33_n533, us33_n534, us33_n535, us33_n536, us33_n537, us33_n538, us33_n539, 
       us33_n540, us33_n541, us33_n542, us33_n543, us33_n544, us33_n545, us33_n546, us33_n547, us33_n548, 
       us33_n549, us33_n550, us33_n551, us33_n552, us33_n553, us33_n554, us33_n555, us33_n556, us33_n557, 
       us33_n558, us33_n559, us33_n560, us33_n561, us33_n562, us33_n563, us33_n564, us33_n565, us33_n566, 
       us33_n567, us33_n568, us33_n569, us33_n570, us33_n571, us33_n572, us33_n573, us33_n574, us33_n575, 
       us33_n576, us33_n577, us33_n578, us33_n579, us33_n580, us33_n581, us33_n582, us33_n583, us33_n584, 
       us33_n585, us33_n586, us33_n587, us33_n588, us33_n589, us33_n590, us33_n591, us33_n592, us33_n593, 
       us33_n594, us33_n595, us33_n596, us33_n597, us33_n598, us33_n599, us33_n600, us33_n601, us33_n602, 
       us33_n603, us33_n604, us33_n605, us33_n606, us33_n607, us33_n608, us33_n609, us33_n610, us33_n611, 
       us33_n612, us33_n613, us33_n614, us33_n615, us33_n616, us33_n617, us33_n618, us33_n619, us33_n620, 
       us33_n621, us33_n622, us33_n623, us33_n624, us33_n625, us33_n626, us33_n627, us33_n628, us33_n629, 
       us33_n630, us33_n631, us33_n632, us33_n633, us33_n634, us33_n635, us33_n636, us33_n637, us33_n638, 
       us33_n639, us33_n640, us33_n641, us33_n642, us33_n643, us33_n644, us33_n645, us33_n646, us33_n647, 
       us33_n648, us33_n649, us33_n650, us33_n651, us33_n652, us33_n653, us33_n654, us33_n655, us33_n656, 
       us33_n657, us33_n658, us33_n659, us33_n660, us33_n661, us33_n662, us33_n663, us33_n664, us33_n665, 
       us33_n666, us33_n667, us33_n668, us33_n669, us33_n670, us33_n671, us33_n672, us33_n673, us33_n674, 
       us33_n675, us33_n676, us33_n677, us33_n678, us33_n679, us33_n680, us33_n681, us33_n682, us33_n683, 
       us33_n684, us33_n685, us33_n686, us33_n687, us33_n688, us33_n689, us33_n690, us33_n691, us33_n692, 
       us33_n693, us33_n694, us33_n695, us33_n696, us33_n697, us33_n698, us33_n699, us33_n700, us33_n701, 
       us33_n702, us33_n703, us33_n704, us33_n705, us33_n706, us33_n707, us33_n708, us33_n709, us33_n710, 
       us33_n711, us33_n712, us33_n713, us33_n714, us33_n715, us33_n716, us33_n717, us33_n718, us33_n719, 
       us33_n720, us33_n721, us33_n722, us33_n723, us33_n724, us33_n725, us33_n726, us33_n727, us33_n728, 
       us33_n729, us33_n730, us33_n731, us33_n732, us33_n733, us33_n734, us33_n735, us33_n736, us33_n737, 
       us33_n738, us33_n739, us33_n740, us33_n741, us33_n742, us33_n743, us33_n744, us33_n745, us33_n746, 
       us33_n747, us33_n748, us33_n749, us33_n750, us33_n751, us33_n752, us33_n753, us33_n754, us33_n755, 
       us33_n756, us33_n757, us33_n758, us33_n759, us33_n760, us33_n761, us33_n762, us33_n763, us33_n764, 
       us33_n765, us33_n766, us33_n767, us33_n768, us33_n769, us33_n770, us33_n771, us33_n772, us33_n773, 
       us33_n774, us33_n775, us33_n776, us33_n777, us33_n778, us33_n779, us33_n780, us33_n781, us33_n782, 
       us33_n783, us33_n784, us33_n785, us33_n786, us33_n787, us33_n788, us33_n789, us33_n790, us33_n791, 
       us33_n792, us33_n793, us33_n794, us33_n795, us33_n796, us33_n797, us33_n798, us33_n799, us33_n800, 
       us33_n801, us33_n802, us33_n803, us33_n804, us33_n805, us33_n806, us33_n807, us33_n808, us33_n809, 
       us33_n810, us33_n811, us33_n812, us33_n813, us33_n814, us33_n815, us33_n816, us33_n817, us33_n818, 
       us33_n819, us33_n820, us33_n821, us33_n822, us33_n823, us33_n824, us33_n825, us33_n826, us33_n827, 
       us33_n828, us33_n829, us33_n830, us33_n831, us33_n832, us33_n833, us33_n834, us33_n835, us33_n836, 
       us33_n837, us33_n838, us33_n839, us33_n840, us33_n841, us33_n842, us33_n843, us33_n844, us33_n845, 
       us33_n846, us33_n847, us33_n848, us33_n849, us33_n850, us33_n851, us33_n852, us33_n853, us33_n854, 
       us33_n855, us33_n856, us33_n857, us33_n858, us33_n859, us33_n860, us33_n861, us33_n862, us33_n863, 
       us33_n864, us33_n865, us33_n866, us33_n867, us33_n868, us33_n869, us33_n870, us33_n871, us33_n872, 
       us33_n873, us33_n874, us33_n875,  us33_n876;
  NOR2_X1 us01_U10 (.ZN( us01_n573 ) , .A1( us01_n620 ) , .A2( us01_n743 ) );
  AOI211_X1 us01_U100 (.B( us01_n537 ) , .A( us01_n538 ) , .ZN( us01_n549 ) , .C2( us01_n837 ) , .C1( us01_n849 ) );
  NOR4_X1 us01_U101 (.A4( us01_n542 ) , .A3( us01_n543 ) , .A2( us01_n544 ) , .A1( us01_n545 ) , .ZN( us01_n546 ) );
  NOR4_X1 us01_U102 (.A4( us01_n607 ) , .A3( us01_n608 ) , .A2( us01_n609 ) , .A1( us01_n610 ) , .ZN( us01_n617 ) );
  NOR4_X1 us01_U103 (.ZN( us01_n618 ) , .A1( us01_n654 ) , .A3( us01_n664 ) , .A4( us01_n680 ) , .A2( us01_n764 ) );
  NOR4_X1 us01_U104 (.A4( us01_n612 ) , .A3( us01_n613 ) , .A2( us01_n614 ) , .A1( us01_n615 ) , .ZN( us01_n616 ) );
  NOR2_X1 us01_U105 (.ZN( us01_n684 ) , .A1( us01_n829 ) , .A2( us01_n830 ) );
  NAND4_X1 us01_U106 (.A4( us01_n471 ) , .A3( us01_n472 ) , .A2( us01_n473 ) , .A1( us01_n474 ) , .ZN( us01_n676 ) );
  NOR4_X1 us01_U107 (.A4( us01_n468 ) , .ZN( us01_n474 ) , .A3( us01_n554 ) , .A1( us01_n733 ) , .A2( us01_n753 ) );
  NOR4_X1 us01_U108 (.ZN( us01_n473 ) , .A1( us01_n529 ) , .A3( us01_n566 ) , .A4( us01_n598 ) , .A2( us01_n640 ) );
  NOR4_X1 us01_U109 (.ZN( us01_n472 ) , .A1( us01_n504 ) , .A3( us01_n542 ) , .A2( us01_n581 ) , .A4( us01_n714 ) );
  NOR2_X1 us01_U11 (.ZN( us01_n493 ) , .A1( us01_n676 ) , .A2( us01_n692 ) );
  NAND4_X1 us01_U110 (.A4( us01_n689 ) , .A3( us01_n690 ) , .A1( us01_n691 ) , .ZN( us01_n774 ) , .A2( us01_n870 ) );
  INV_X1 us01_U111 (.A( us01_n677 ) , .ZN( us01_n870 ) );
  AOI221_X1 us01_U112 (.A( us01_n679 ) , .ZN( us01_n690 ) , .B2( us01_n838 ) , .C1( us01_n840 ) , .C2( us01_n860 ) , .B1( us01_n863 ) );
  NOR4_X1 us01_U113 (.A4( us01_n685 ) , .A3( us01_n686 ) , .A2( us01_n687 ) , .A1( us01_n688 ) , .ZN( us01_n689 ) );
  NOR2_X1 us01_U114 (.ZN( us01_n731 ) , .A2( us01_n830 ) , .A1( us01_n843 ) );
  NAND4_X1 us01_U115 (.A4( us01_n717 ) , .A3( us01_n718 ) , .A2( us01_n719 ) , .ZN( us01_n739 ) , .A1( us01_n855 ) );
  AOI221_X1 us01_U116 (.A( us01_n708 ) , .ZN( us01_n719 ) , .C2( us01_n842 ) , .B2( us01_n843 ) , .C1( us01_n859 ) , .B1( us01_n860 ) );
  INV_X1 us01_U117 (.A( us01_n707 ) , .ZN( us01_n855 ) );
  NOR4_X1 us01_U118 (.A4( us01_n713 ) , .A3( us01_n714 ) , .A2( us01_n715 ) , .A1( us01_n716 ) , .ZN( us01_n717 ) );
  NOR2_X1 us01_U119 (.ZN( us01_n645 ) , .A1( us01_n852 ) , .A2( us01_n866 ) );
  NOR2_X1 us01_U12 (.A1( us01_n676 ) , .ZN( us01_n691 ) , .A2( us01_n805 ) );
  NAND4_X1 us01_U120 (.A4( us01_n571 ) , .A3( us01_n572 ) , .A1( us01_n573 ) , .ZN( us01_n721 ) , .A2( us01_n872 ) );
  AOI221_X1 us01_U121 (.A( us01_n562 ) , .C2( us01_n563 ) , .ZN( us01_n572 ) , .B2( us01_n843 ) , .B1( us01_n850 ) , .C1( us01_n851 ) );
  NOR4_X1 us01_U122 (.A4( us01_n567 ) , .A3( us01_n568 ) , .A2( us01_n569 ) , .A1( us01_n570 ) , .ZN( us01_n571 ) );
  INV_X1 us01_U123 (.A( us01_n605 ) , .ZN( us01_n872 ) );
  NAND4_X1 us01_U124 (.A4( us01_n491 ) , .A3( us01_n492 ) , .A1( us01_n493 ) , .ZN( us01_n800 ) , .A2( us01_n865 ) );
  AOI221_X1 us01_U125 (.A( us01_n487 ) , .ZN( us01_n492 ) , .B2( us01_n834 ) , .C2( us01_n839 ) , .C1( us01_n849 ) , .B1( us01_n858 ) );
  INV_X1 us01_U126 (.A( us01_n776 ) , .ZN( us01_n865 ) );
  NOR4_X1 us01_U127 (.A2( us01_n489 ) , .A1( us01_n490 ) , .ZN( us01_n491 ) , .A3( us01_n578 ) , .A4( us01_n610 ) );
  NOR4_X1 us01_U128 (.A3( us01_n753 ) , .A2( us01_n754 ) , .A1( us01_n755 ) , .ZN( us01_n756 ) , .A4( us01_n867 ) );
  AOI211_X1 us01_U129 (.B( us01_n743 ) , .A( us01_n744 ) , .ZN( us01_n757 ) , .C1( us01_n830 ) , .C2( us01_n851 ) );
  NOR3_X1 us01_U13 (.ZN( us01_n502 ) , .A2( us01_n677 ) , .A3( us01_n775 ) , .A1( us01_n874 ) );
  NOR3_X1 us01_U130 (.A3( us01_n739 ) , .A2( us01_n740 ) , .A1( us01_n741 ) , .ZN( us01_n758 ) );
  NOR4_X1 us01_U131 (.A4( us01_n732 ) , .A3( us01_n733 ) , .A2( us01_n734 ) , .A1( us01_n735 ) , .ZN( us01_n736 ) );
  AOI211_X1 us01_U132 (.B( us01_n723 ) , .A( us01_n724 ) , .ZN( us01_n737 ) , .C1( us01_n841 ) , .C2( us01_n853 ) );
  NOR3_X1 us01_U133 (.A3( us01_n720 ) , .A1( us01_n721 ) , .ZN( us01_n738 ) , .A2( us01_n739 ) );
  INV_X1 us01_U134 (.A( us01_n760 ) , .ZN( us01_n828 ) );
  NAND4_X1 us01_U135 (.ZN( sa01_sr_3 ) , .A4( us01_n702 ) , .A3( us01_n703 ) , .A2( us01_n704 ) , .A1( us01_n705 ) );
  NOR4_X1 us01_U136 (.A4( us01_n698 ) , .A3( us01_n699 ) , .A2( us01_n700 ) , .A1( us01_n701 ) , .ZN( us01_n702 ) );
  AOI211_X1 us01_U137 (.B( us01_n692 ) , .A( us01_n693 ) , .ZN( us01_n703 ) , .C2( us01_n829 ) , .C1( us01_n849 ) );
  NOR2_X1 us01_U138 (.ZN( us01_n705 ) , .A2( us01_n774 ) , .A1( us01_n798 ) );
  OR4_X1 us01_U139 (.A4( us01_n680 ) , .A3( us01_n681 ) , .A2( us01_n682 ) , .A1( us01_n683 ) , .ZN( us01_n688 ) );
  INV_X1 us01_U14 (.A( us01_n704 ) , .ZN( us01_n874 ) );
  OR4_X1 us01_U140 (.ZN( us01_n464 ) , .A4( us01_n516 ) , .A3( us01_n527 ) , .A2( us01_n576 ) , .A1( us01_n710 ) );
  OR4_X1 us01_U141 (.A4( us01_n564 ) , .A3( us01_n565 ) , .A2( us01_n566 ) , .ZN( us01_n570 ) , .A1( us01_n663 ) );
  OR4_X1 us01_U142 (.A4( us01_n516 ) , .A2( us01_n517 ) , .A1( us01_n518 ) , .ZN( us01_n520 ) , .A3( us01_n819 ) );
  OR4_X1 us01_U143 (.ZN( us01_n490 ) , .A4( us01_n532 ) , .A2( us01_n545 ) , .A1( us01_n557 ) , .A3( us01_n630 ) );
  OR4_X1 us01_U144 (.A4( us01_n578 ) , .A3( us01_n579 ) , .A2( us01_n580 ) , .A1( us01_n581 ) , .ZN( us01_n582 ) );
  INV_X1 us01_U145 (.A( us01_n695 ) , .ZN( us01_n836 ) );
  NAND2_X1 us01_U146 (.ZN( us01_n611 ) , .A2( us01_n835 ) , .A1( us01_n871 ) );
  OR3_X1 us01_U147 (.A3( us01_n504 ) , .A2( us01_n505 ) , .A1( us01_n506 ) , .ZN( us01_n509 ) );
  AOI221_X1 us01_U148 (.A( us01_n711 ) , .B2( us01_n712 ) , .ZN( us01_n718 ) , .C1( us01_n830 ) , .B1( us01_n837 ) , .C2( us01_n861 ) );
  OR2_X1 us01_U149 (.A2( us01_n709 ) , .A1( us01_n710 ) , .ZN( us01_n711 ) );
  INV_X1 us01_U15 (.A( us01_n678 ) , .ZN( us01_n838 ) );
  INV_X1 us01_U150 (.A( us01_n461 ) , .ZN( us01_n862 ) );
  OAI21_X1 us01_U151 (.ZN( us01_n461 ) , .B1( us01_n807 ) , .A( us01_n832 ) , .B2( us01_n849 ) );
  INV_X1 us01_U152 (.A( us01_n752 ) , .ZN( us01_n867 ) );
  OAI21_X1 us01_U153 (.B1( us01_n751 ) , .ZN( us01_n752 ) , .A( us01_n843 ) , .B2( us01_n866 ) );
  INV_X1 us01_U154 (.A( us01_n670 ) , .ZN( us01_n857 ) );
  AOI21_X1 us01_U155 (.A( us01_n668 ) , .B1( us01_n669 ) , .ZN( us01_n670 ) , .B2( us01_n854 ) );
  AOI222_X1 us01_U156 (.ZN( us01_n658 ) , .A2( us01_n837 ) , .B1( us01_n839 ) , .C2( us01_n843 ) , .A1( us01_n858 ) , .C1( us01_n861 ) , .B2( us01_n868 ) );
  INV_X1 us01_U157 (.A( us01_n645 ) , .ZN( us01_n868 ) );
  OAI22_X1 us01_U158 (.ZN( us01_n481 ) , .A1( us01_n706 ) , .B2( us01_n783 ) , .A2( us01_n804 ) , .B1( us01_n810 ) );
  OAI22_X1 us01_U159 (.ZN( us01_n635 ) , .A1( us01_n697 ) , .B2( us01_n726 ) , .A2( us01_n760 ) , .B1( us01_n814 ) );
  NOR4_X1 us01_U16 (.A4( us01_n443 ) , .A3( us01_n444 ) , .A2( us01_n514 ) , .A1( us01_n539 ) , .ZN( us01_n704 ) );
  OAI222_X1 us01_U160 (.ZN( us01_n503 ) , .C2( us01_n623 ) , .B2( us01_n645 ) , .B1( us01_n745 ) , .A2( us01_n746 ) , .C1( us01_n803 ) , .A1( us01_n804 ) );
  OAI222_X1 us01_U161 (.B2( us01_n745 ) , .B1( us01_n746 ) , .A2( us01_n747 ) , .ZN( us01_n755 ) , .C2( us01_n803 ) , .C1( us01_n812 ) , .A1( us01_n815 ) );
  OAI222_X1 us01_U162 (.B2( us01_n706 ) , .ZN( us01_n707 ) , .C2( us01_n722 ) , .B1( us01_n745 ) , .A1( us01_n804 ) , .C1( us01_n812 ) , .A2( us01_n813 ) );
  AOI22_X1 us01_U163 (.ZN( us01_n694 ) , .A1( us01_n828 ) , .B2( us01_n841 ) , .A2( us01_n863 ) , .B1( us01_n866 ) );
  AOI22_X1 us01_U164 (.A2( us01_n780 ) , .ZN( us01_n781 ) , .B2( us01_n829 ) , .A1( us01_n832 ) , .B1( us01_n861 ) );
  INV_X1 us01_U165 (.A( us01_n728 ) , .ZN( us01_n837 ) );
  AOI221_X1 us01_U166 (.A( us01_n762 ) , .ZN( us01_n772 ) , .C2( us01_n808 ) , .B2( us01_n833 ) , .C1( us01_n853 ) , .B1( us01_n864 ) );
  AOI21_X1 us01_U167 (.B2( us01_n761 ) , .ZN( us01_n762 ) , .A( us01_n786 ) , .B1( us01_n790 ) );
  INV_X1 us01_U168 (.A( us01_n759 ) , .ZN( us01_n833 ) );
  INV_X1 us01_U169 (.A( us01_n788 ) , .ZN( us01_n830 ) );
  OR3_X1 us01_U17 (.ZN( us01_n444 ) , .A1( us01_n526 ) , .A3( us01_n575 ) , .A2( us01_n873 ) );
  OAI221_X1 us01_U170 (.A( us01_n725 ) , .C2( us01_n726 ) , .B2( us01_n727 ) , .B1( us01_n728 ) , .ZN( us01_n735 ) , .C1( us01_n815 ) );
  AOI22_X1 us01_U171 (.ZN( us01_n725 ) , .B1( us01_n830 ) , .A2( us01_n836 ) , .A1( us01_n861 ) , .B2( us01_n864 ) );
  NAND2_X1 us01_U172 (.A1( us01_n449 ) , .A2( us01_n451 ) , .ZN( us01_n760 ) );
  OAI22_X1 us01_U173 (.ZN( us01_n622 ) , .B1( us01_n667 ) , .B2( us01_n745 ) , .A1( us01_n813 ) , .A2( us01_n814 ) );
  OAI22_X1 us01_U174 (.A1( us01_n722 ) , .ZN( us01_n724 ) , .B2( us01_n748 ) , .B1( us01_n810 ) , .A2( us01_n814 ) );
  OAI22_X1 us01_U175 (.ZN( us01_n487 ) , .A1( us01_n722 ) , .B2( us01_n726 ) , .B1( us01_n728 ) , .A2( us01_n777 ) );
  OAI22_X1 us01_U176 (.B2( us01_n777 ) , .B1( us01_n778 ) , .ZN( us01_n779 ) , .A2( us01_n812 ) , .A1( us01_n813 ) );
  OAI22_X1 us01_U177 (.B2( us01_n748 ) , .B1( us01_n749 ) , .A1( us01_n750 ) , .ZN( us01_n754 ) , .A2( us01_n804 ) );
  NOR3_X1 us01_U178 (.ZN( us01_n750 ) , .A2( us01_n851 ) , .A1( us01_n861 ) , .A3( us01_n863 ) );
  NOR2_X1 us01_U179 (.ZN( us01_n749 ) , .A2( us01_n850 ) , .A1( us01_n858 ) );
  OR4_X1 us01_U18 (.A4( us01_n440 ) , .A2( us01_n441 ) , .A1( us01_n442 ) , .ZN( us01_n443 ) , .A3( us01_n551 ) );
  INV_X1 us01_U180 (.A( us01_n803 ) , .ZN( us01_n858 ) );
  OAI22_X1 us01_U181 (.B2( us01_n742 ) , .ZN( us01_n744 ) , .A2( us01_n760 ) , .B1( us01_n778 ) , .A1( us01_n790 ) );
  OAI22_X1 us01_U182 (.ZN( us01_n494 ) , .A2( us01_n742 ) , .A1( us01_n778 ) , .B1( us01_n789 ) , .B2( us01_n804 ) );
  OAI22_X1 us01_U183 (.B2( us01_n801 ) , .B1( us01_n802 ) , .A2( us01_n803 ) , .A1( us01_n804 ) , .ZN( us01_n806 ) );
  OAI22_X1 us01_U184 (.ZN( us01_n693 ) , .A2( us01_n728 ) , .A1( us01_n778 ) , .B1( us01_n789 ) , .B2( us01_n815 ) );
  NOR2_X1 us01_U185 (.ZN( us01_n713 ) , .A1( us01_n803 ) , .A2( us01_n815 ) );
  NOR2_X1 us01_U186 (.A1( us01_n697 ) , .ZN( us01_n766 ) , .A2( us01_n811 ) );
  INV_X1 us01_U187 (.A( us01_n786 ) , .ZN( us01_n843 ) );
  NOR2_X1 us01_U188 (.ZN( us01_n539 ) , .A2( us01_n695 ) , .A1( us01_n697 ) );
  INV_X1 us01_U189 (.A( us01_n742 ) , .ZN( us01_n835 ) );
  INV_X1 us01_U19 (.A( us01_n611 ) , .ZN( us01_n873 ) );
  INV_X1 us01_U190 (.A( us01_n814 ) , .ZN( us01_n829 ) );
  INV_X1 us01_U191 (.A( us01_n812 ) , .ZN( us01_n831 ) );
  OAI22_X1 us01_U192 (.B1( us01_n488 ) , .ZN( us01_n489 ) , .A1( us01_n684 ) , .A2( us01_n761 ) , .B2( us01_n815 ) );
  NOR3_X1 us01_U193 (.ZN( us01_n488 ) , .A1( us01_n780 ) , .A2( us01_n848 ) , .A3( us01_n861 ) );
  NOR2_X1 us01_U194 (.A2( us01_n742 ) , .ZN( us01_n753 ) , .A1( us01_n803 ) );
  NOR2_X1 us01_U195 (.ZN( us01_n733 ) , .A2( us01_n801 ) , .A1( us01_n803 ) );
  INV_X1 us01_U196 (.A( us01_n790 ) , .ZN( us01_n849 ) );
  NOR2_X1 us01_U197 (.A2( us01_n742 ) , .ZN( us01_n767 ) , .A1( us01_n810 ) );
  NOR2_X1 us01_U198 (.ZN( us01_n664 ) , .A1( us01_n726 ) , .A2( us01_n801 ) );
  OAI22_X1 us01_U199 (.ZN( us01_n708 ) , .A2( us01_n726 ) , .B2( us01_n727 ) , .A1( us01_n742 ) , .B1( us01_n811 ) );
  AOI222_X1 us01_U20 (.ZN( us01_n561 ) , .B1( us01_n828 ) , .C1( us01_n839 ) , .A2( us01_n841 ) , .A1( us01_n852 ) , .B2( us01_n861 ) , .C2( us01_n871 ) );
  NOR2_X1 us01_U200 (.ZN( us01_n650 ) , .A1( us01_n667 ) , .A2( us01_n812 ) );
  NOR2_X1 us01_U201 (.ZN( us01_n592 ) , .A2( us01_n695 ) , .A1( us01_n726 ) );
  NOR2_X1 us01_U202 (.A1( us01_n667 ) , .ZN( us01_n671 ) , .A2( us01_n742 ) );
  NOR2_X1 us01_U203 (.ZN( us01_n600 ) , .A1( us01_n667 ) , .A2( us01_n801 ) );
  NOR2_X1 us01_U204 (.A1( us01_n667 ) , .ZN( us01_n686 ) , .A2( us01_n814 ) );
  NOR2_X1 us01_U205 (.ZN( us01_n568 ) , .A1( us01_n726 ) , .A2( us01_n804 ) );
  NOR2_X1 us01_U206 (.A1( us01_n667 ) , .ZN( us01_n764 ) , .A2( us01_n811 ) );
  NOR2_X1 us01_U207 (.ZN( us01_n525 ) , .A1( us01_n667 ) , .A2( us01_n777 ) );
  NOR2_X1 us01_U208 (.ZN( us01_n652 ) , .A1( us01_n726 ) , .A2( us01_n811 ) );
  NOR2_X1 us01_U209 (.ZN( us01_n505 ) , .A1( us01_n810 ) , .A2( us01_n815 ) );
  NOR4_X1 us01_U21 (.ZN( us01_n471 ) , .A2( us01_n519 ) , .A4( us01_n592 ) , .A1( us01_n607 ) , .A3( us01_n627 ) );
  NOR2_X1 us01_U210 (.ZN( us01_n659 ) , .A1( us01_n727 ) , .A2( us01_n788 ) );
  NOR2_X1 us01_U211 (.ZN( us01_n544 ) , .A2( us01_n778 ) , .A1( us01_n812 ) );
  NOR2_X1 us01_U212 (.ZN( us01_n575 ) , .A2( us01_n697 ) , .A1( us01_n812 ) );
  NOR2_X1 us01_U213 (.ZN( us01_n507 ) , .A1( us01_n727 ) , .A2( us01_n777 ) );
  NOR2_X1 us01_U214 (.ZN( us01_n716 ) , .A2( us01_n722 ) , .A1( us01_n742 ) );
  INV_X1 us01_U215 (.A( us01_n748 ) , .ZN( us01_n840 ) );
  NOR2_X1 us01_U216 (.ZN( us01_n530 ) , .A2( us01_n747 ) , .A1( us01_n748 ) );
  NOR2_X1 us01_U217 (.ZN( us01_n660 ) , .A2( us01_n695 ) , .A1( us01_n727 ) );
  NOR2_X1 us01_U218 (.ZN( us01_n613 ) , .A1( us01_n783 ) , .A2( us01_n813 ) );
  NOR2_X1 us01_U219 (.ZN( us01_n627 ) , .A2( us01_n726 ) , .A1( us01_n783 ) );
  NOR4_X1 us01_U22 (.ZN( us01_n477 ) , .A1( us01_n518 ) , .A4( us01_n555 ) , .A3( us01_n580 ) , .A2( us01_n628 ) );
  NOR2_X1 us01_U220 (.ZN( us01_n609 ) , .A2( us01_n778 ) , .A1( us01_n804 ) );
  NOR2_X1 us01_U221 (.ZN( us01_n661 ) , .A1( us01_n727 ) , .A2( us01_n783 ) );
  NOR2_X1 us01_U222 (.ZN( us01_n626 ) , .A2( us01_n667 ) , .A1( us01_n783 ) );
  NOR2_X1 us01_U223 (.ZN( us01_n599 ) , .A2( us01_n778 ) , .A1( us01_n801 ) );
  INV_X1 us01_U224 (.A( us01_n745 ) , .ZN( us01_n832 ) );
  NOR2_X1 us01_U225 (.ZN( us01_n554 ) , .A1( us01_n760 ) , .A2( us01_n803 ) );
  NOR2_X1 us01_U226 (.ZN( us01_n529 ) , .A2( us01_n778 ) , .A1( us01_n814 ) );
  NOR2_X1 us01_U227 (.ZN( us01_n526 ) , .A2( us01_n722 ) , .A1( us01_n801 ) );
  NOR2_X1 us01_U228 (.A2( us01_n706 ) , .A1( us01_n748 ) , .ZN( us01_n769 ) );
  NOR2_X1 us01_U229 (.ZN( us01_n597 ) , .A2( us01_n789 ) , .A1( us01_n814 ) );
  NOR4_X1 us01_U23 (.ZN( us01_n454 ) , .A2( us01_n515 ) , .A1( us01_n541 ) , .A3( us01_n577 ) , .A4( us01_n613 ) );
  NOR2_X1 us01_U230 (.ZN( us01_n555 ) , .A1( us01_n790 ) , .A2( us01_n812 ) );
  NOR2_X1 us01_U231 (.ZN( us01_n542 ) , .A2( us01_n783 ) , .A1( us01_n790 ) );
  NOR2_X1 us01_U232 (.A2( us01_n695 ) , .ZN( us01_n714 ) , .A1( us01_n790 ) );
  NOR2_X1 us01_U233 (.ZN( us01_n665 ) , .A1( us01_n748 ) , .A2( us01_n813 ) );
  NOR2_X1 us01_U234 (.ZN( us01_n543 ) , .A1( us01_n747 ) , .A2( us01_n812 ) );
  NOR2_X1 us01_U235 (.ZN( us01_n553 ) , .A1( us01_n748 ) , .A2( us01_n789 ) );
  NOR2_X1 us01_U236 (.ZN( us01_n506 ) , .A2( us01_n778 ) , .A1( us01_n783 ) );
  NOR2_X1 us01_U237 (.ZN( us01_n541 ) , .A2( us01_n706 ) , .A1( us01_n783 ) );
  NOR2_X1 us01_U238 (.ZN( us01_n514 ) , .A1( us01_n706 ) , .A2( us01_n742 ) );
  NOR2_X1 us01_U239 (.ZN( us01_n662 ) , .A1( us01_n783 ) , .A2( us01_n789 ) );
  NOR4_X1 us01_U24 (.A4( us01_n530 ) , .A3( us01_n531 ) , .A2( us01_n532 ) , .ZN( us01_n533 ) , .A1( us01_n818 ) );
  NOR2_X1 us01_U240 (.ZN( us01_n556 ) , .A1( us01_n706 ) , .A2( us01_n814 ) );
  NOR2_X1 us01_U241 (.ZN( us01_n515 ) , .A1( us01_n706 ) , .A2( us01_n801 ) );
  NOR2_X1 us01_U242 (.ZN( us01_n612 ) , .A1( us01_n760 ) , .A2( us01_n810 ) );
  NOR2_X1 us01_U243 (.ZN( us01_n629 ) , .A1( us01_n722 ) , .A2( us01_n811 ) );
  NOR2_X1 us01_U244 (.A1( us01_n747 ) , .ZN( us01_n765 ) , .A2( us01_n801 ) );
  NOR2_X1 us01_U245 (.ZN( us01_n528 ) , .A2( us01_n742 ) , .A1( us01_n790 ) );
  INV_X1 us01_U246 (.A( us01_n804 ) , .ZN( us01_n839 ) );
  OAI22_X1 us01_U247 (.B1( us01_n438 ) , .ZN( us01_n442 ) , .A2( us01_n726 ) , .A1( us01_n742 ) , .B2( us01_n747 ) );
  NOR3_X1 us01_U248 (.ZN( us01_n438 ) , .A2( us01_n834 ) , .A3( us01_n835 ) , .A1( us01_n844 ) );
  INV_X1 us01_U249 (.A( us01_n726 ) , .ZN( us01_n850 ) );
  NOR4_X1 us01_U25 (.A4( us01_n539 ) , .A3( us01_n540 ) , .A2( us01_n541 ) , .ZN( us01_n548 ) , .A1( us01_n686 ) );
  NOR2_X1 us01_U250 (.ZN( us01_n519 ) , .A1( us01_n788 ) , .A2( us01_n810 ) );
  NOR2_X1 us01_U251 (.ZN( us01_n668 ) , .A1( us01_n788 ) , .A2( us01_n803 ) );
  AOI21_X1 us01_U252 (.ZN( us01_n550 ) , .B1( us01_n667 ) , .A( us01_n695 ) , .B2( us01_n803 ) );
  AOI21_X1 us01_U253 (.ZN( us01_n587 ) , .B2( us01_n697 ) , .B1( us01_n813 ) , .A( us01_n815 ) );
  NOR2_X1 us01_U254 (.ZN( us01_n504 ) , .A2( us01_n726 ) , .A1( us01_n760 ) );
  NOR2_X1 us01_U255 (.ZN( us01_n653 ) , .A1( us01_n788 ) , .A2( us01_n813 ) );
  INV_X1 us01_U256 (.A( us01_n801 ) , .ZN( us01_n841 ) );
  NOR2_X1 us01_U257 (.ZN( us01_n628 ) , .A1( us01_n745 ) , .A2( us01_n813 ) );
  NOR2_X1 us01_U258 (.ZN( us01_n545 ) , .A1( us01_n697 ) , .A2( us01_n742 ) );
  INV_X1 us01_U259 (.A( us01_n697 ) , .ZN( us01_n851 ) );
  NOR2_X1 us01_U26 (.ZN( us01_n678 ) , .A2( us01_n832 ) , .A1( us01_n837 ) );
  NOR2_X1 us01_U260 (.ZN( us01_n640 ) , .A2( us01_n786 ) , .A1( us01_n789 ) );
  AOI21_X1 us01_U261 (.ZN( us01_n648 ) , .A( us01_n777 ) , .B1( us01_n790 ) , .B2( us01_n803 ) );
  NOR2_X1 us01_U262 (.ZN( us01_n666 ) , .A2( us01_n706 ) , .A1( us01_n788 ) );
  NOR2_X1 us01_U263 (.A2( us01_n695 ) , .A1( us01_n778 ) , .ZN( us01_n818 ) );
  NOR2_X1 us01_U264 (.A1( us01_n695 ) , .ZN( us01_n768 ) , .A2( us01_n813 ) );
  AOI21_X1 us01_U265 (.ZN( us01_n624 ) , .B2( us01_n667 ) , .A( us01_n788 ) , .B1( us01_n789 ) );
  NOR2_X1 us01_U266 (.ZN( us01_n577 ) , .A2( us01_n706 ) , .A1( us01_n728 ) );
  INV_X1 us01_U267 (.A( us01_n761 ) , .ZN( us01_n864 ) );
  NOR2_X1 us01_U268 (.A2( us01_n706 ) , .A1( us01_n760 ) , .ZN( us01_n792 ) );
  NOR2_X1 us01_U269 (.ZN( us01_n607 ) , .A2( us01_n722 ) , .A1( us01_n815 ) );
  AOI222_X1 us01_U27 (.ZN( us01_n467 ) , .B1( us01_n830 ) , .A1( us01_n837 ) , .C1( us01_n840 ) , .C2( us01_n849 ) , .A2( us01_n853 ) , .B2( us01_n863 ) );
  NOR2_X1 us01_U270 (.ZN( us01_n531 ) , .A2( us01_n722 ) , .A1( us01_n728 ) );
  AOI21_X1 us01_U271 (.ZN( us01_n508 ) , .B2( us01_n667 ) , .A( us01_n728 ) , .B1( us01_n813 ) );
  AOI21_X1 us01_U272 (.ZN( us01_n537 ) , .B2( us01_n810 ) , .A( us01_n812 ) , .B1( us01_n813 ) );
  INV_X1 us01_U273 (.A( us01_n727 ) , .ZN( us01_n866 ) );
  NOR2_X1 us01_U274 (.ZN( us01_n540 ) , .A1( us01_n760 ) , .A2( us01_n789 ) );
  INV_X1 us01_U275 (.A( us01_n810 ) , .ZN( us01_n852 ) );
  AOI21_X1 us01_U276 (.B1( us01_n697 ) , .ZN( us01_n698 ) , .A( us01_n730 ) , .B2( us01_n761 ) );
  NOR2_X1 us01_U277 (.ZN( us01_n579 ) , .A1( us01_n667 ) , .A2( us01_n786 ) );
  AOI21_X1 us01_U278 (.ZN( us01_n589 ) , .B2( us01_n761 ) , .A( us01_n783 ) , .B1( us01_n810 ) );
  NOR2_X1 us01_U279 (.ZN( us01_n654 ) , .A1( us01_n745 ) , .A2( us01_n778 ) );
  NOR4_X1 us01_U28 (.A1( us01_n464 ) , .ZN( us01_n465 ) , .A4( us01_n540 ) , .A2( us01_n552 ) , .A3( us01_n612 ) );
  INV_X1 us01_U280 (.A( us01_n789 ) , .ZN( us01_n871 ) );
  AOI21_X1 us01_U281 (.B1( us01_n623 ) , .ZN( us01_n625 ) , .A( us01_n761 ) , .B2( us01_n812 ) );
  NOR2_X1 us01_U282 (.ZN( us01_n683 ) , .A1( us01_n727 ) , .A2( us01_n814 ) );
  AOI21_X1 us01_U283 (.A( us01_n813 ) , .B2( us01_n814 ) , .B1( us01_n815 ) , .ZN( us01_n816 ) );
  AOI21_X1 us01_U284 (.ZN( us01_n647 ) , .B1( us01_n727 ) , .B2( us01_n761 ) , .A( us01_n811 ) );
  AOI21_X1 us01_U285 (.A( us01_n810 ) , .B2( us01_n811 ) , .B1( us01_n812 ) , .ZN( us01_n817 ) );
  AOI21_X1 us01_U286 (.ZN( us01_n513 ) , .A( us01_n727 ) , .B1( us01_n748 ) , .B2( us01_n801 ) );
  AOI21_X1 us01_U287 (.ZN( us01_n497 ) , .B1( us01_n678 ) , .A( us01_n810 ) , .B2( us01_n814 ) );
  NOR2_X1 us01_U288 (.ZN( us01_n518 ) , .A2( us01_n706 ) , .A1( us01_n812 ) );
  AOI21_X1 us01_U289 (.ZN( us01_n475 ) , .A( us01_n667 ) , .B1( us01_n748 ) , .B2( us01_n804 ) );
  AOI221_X1 us01_U29 (.ZN( us01_n466 ) , .C2( us01_n712 ) , .B2( us01_n829 ) , .C1( us01_n843 ) , .B1( us01_n858 ) , .A( us01_n862 ) );
  NOR2_X1 us01_U290 (.ZN( us01_n566 ) , .A1( us01_n727 ) , .A2( us01_n760 ) );
  NOR2_X1 us01_U291 (.ZN( us01_n580 ) , .A1( us01_n742 ) , .A2( us01_n813 ) );
  AOI21_X1 us01_U292 (.ZN( us01_n591 ) , .B1( us01_n748 ) , .A( us01_n790 ) , .B2( us01_n811 ) );
  NOR2_X1 us01_U293 (.ZN( us01_n564 ) , .A2( us01_n695 ) , .A1( us01_n761 ) );
  AOI21_X1 us01_U294 (.ZN( us01_n512 ) , .A( us01_n777 ) , .B2( us01_n790 ) , .B1( us01_n810 ) );
  NAND2_X2 us01_U295 (.A2( us01_n462 ) , .A1( us01_n463 ) , .ZN( us01_n810 ) );
  AOI21_X1 us01_U296 (.ZN( us01_n637 ) , .B2( us01_n747 ) , .A( us01_n786 ) , .B1( us01_n810 ) );
  NOR2_X1 us01_U297 (.ZN( us01_n557 ) , .A2( us01_n789 ) , .A1( us01_n801 ) );
  NOR2_X1 us01_U298 (.A2( us01_n811 ) , .A1( us01_n813 ) , .ZN( us01_n819 ) );
  NOR2_X1 us01_U299 (.ZN( us01_n527 ) , .A1( us01_n706 ) , .A2( us01_n777 ) );
  NAND2_X2 us01_U3 (.A1( us01_n447 ) , .A2( us01_n462 ) , .ZN( us01_n722 ) );
  NOR4_X1 us01_U30 (.A4( us01_n512 ) , .A3( us01_n513 ) , .A2( us01_n514 ) , .A1( us01_n515 ) , .ZN( us01_n522 ) );
  NOR2_X1 us01_U300 (.ZN( us01_n517 ) , .A2( us01_n697 ) , .A1( us01_n814 ) );
  NOR2_X1 us01_U301 (.ZN( us01_n681 ) , .A2( us01_n697 ) , .A1( us01_n801 ) );
  NOR2_X1 us01_U302 (.ZN( us01_n576 ) , .A1( us01_n706 ) , .A2( us01_n811 ) );
  INV_X1 us01_U303 (.A( us01_n813 ) , .ZN( us01_n853 ) );
  INV_X1 us01_U304 (.A( us01_n811 ) , .ZN( us01_n834 ) );
  AOI21_X1 us01_U305 (.ZN( us01_n448 ) , .B2( us01_n790 ) , .A( us01_n801 ) , .B1( us01_n813 ) );
  AOI21_X1 us01_U306 (.ZN( us01_n538 ) , .A( us01_n761 ) , .B2( us01_n777 ) , .B1( us01_n815 ) );
  AOI21_X1 us01_U307 (.ZN( us01_n496 ) , .A( us01_n722 ) , .B2( us01_n760 ) , .B1( us01_n812 ) );
  AOI21_X1 us01_U308 (.ZN( us01_n687 ) , .B2( us01_n747 ) , .B1( us01_n761 ) , .A( us01_n804 ) );
  AOI21_X1 us01_U309 (.B1( us01_n684 ) , .ZN( us01_n685 ) , .A( us01_n726 ) , .B2( us01_n759 ) );
  AOI222_X1 us01_U31 (.ZN( us01_n523 ) , .A1( us01_n832 ) , .B2( us01_n835 ) , .C1( us01_n842 ) , .C2( us01_n848 ) , .A2( us01_n850 ) , .B1( us01_n864 ) );
  NOR2_X1 us01_U310 (.ZN( us01_n581 ) , .A1( us01_n790 ) , .A2( us01_n815 ) );
  NOR2_X1 us01_U311 (.ZN( us01_n532 ) , .A1( us01_n722 ) , .A2( us01_n786 ) );
  NOR2_X1 us01_U312 (.ZN( us01_n630 ) , .A2( us01_n695 ) , .A1( us01_n722 ) );
  AOI21_X1 us01_U313 (.A( us01_n788 ) , .B2( us01_n789 ) , .B1( us01_n790 ) , .ZN( us01_n791 ) );
  AOI21_X1 us01_U314 (.A( us01_n731 ) , .ZN( us01_n732 ) , .B2( us01_n778 ) , .B1( us01_n790 ) );
  NOR2_X1 us01_U315 (.ZN( us01_n565 ) , .A1( us01_n745 ) , .A2( us01_n803 ) );
  AOI21_X1 us01_U316 (.ZN( us01_n567 ) , .B1( us01_n748 ) , .B2( us01_n760 ) , .A( us01_n778 ) );
  AOI21_X1 us01_U317 (.ZN( us01_n638 ) , .B2( us01_n745 ) , .A( us01_n790 ) , .B1( us01_n801 ) );
  AOI21_X1 us01_U318 (.ZN( us01_n562 ) , .B1( us01_n722 ) , .A( us01_n777 ) , .B2( us01_n789 ) );
  AOI21_X1 us01_U319 (.ZN( us01_n569 ) , .B2( us01_n695 ) , .B1( us01_n804 ) , .A( us01_n810 ) );
  NOR4_X1 us01_U32 (.A3( us01_n519 ) , .A1( us01_n520 ) , .ZN( us01_n521 ) , .A2( us01_n671 ) , .A4( us01_n767 ) );
  NOR2_X1 us01_U320 (.ZN( us01_n663 ) , .A1( us01_n778 ) , .A2( us01_n811 ) );
  NOR2_X1 us01_U321 (.ZN( us01_n578 ) , .A2( us01_n695 ) , .A1( us01_n789 ) );
  NOR2_X1 us01_U322 (.ZN( us01_n682 ) , .A1( us01_n789 ) , .A2( us01_n811 ) );
  NAND2_X2 us01_U323 (.A1( us01_n450 ) , .A2( us01_n463 ) , .ZN( us01_n667 ) );
  NAND2_X1 us01_U324 (.ZN( us01_n751 ) , .A1( us01_n761 ) , .A2( us01_n803 ) );
  NOR2_X1 us01_U325 (.ZN( us01_n709 ) , .A1( us01_n760 ) , .A2( us01_n761 ) );
  AOI21_X1 us01_U326 (.ZN( us01_n476 ) , .B2( us01_n695 ) , .A( us01_n747 ) , .B1( us01_n777 ) );
  NOR2_X1 us01_U327 (.ZN( us01_n680 ) , .A2( us01_n706 ) , .A1( us01_n815 ) );
  INV_X1 us01_U328 (.A( us01_n778 ) , .ZN( us01_n848 ) );
  OAI21_X1 us01_U329 (.A( us01_n729 ) , .B1( us01_n730 ) , .ZN( us01_n734 ) , .B2( us01_n803 ) );
  AOI221_X1 us01_U33 (.A( us01_n779 ) , .ZN( us01_n796 ) , .C2( us01_n835 ) , .B2( us01_n836 ) , .B1( us01_n863 ) , .C1( us01_n864 ) );
  OAI21_X1 us01_U330 (.ZN( us01_n729 ) , .A( us01_n831 ) , .B2( us01_n850 ) , .B1( us01_n871 ) );
  AOI21_X1 us01_U331 (.ZN( us01_n639 ) , .B1( us01_n678 ) , .A( us01_n789 ) , .B2( us01_n815 ) );
  AOI21_X1 us01_U332 (.ZN( us01_n440 ) , .A( us01_n697 ) , .B1( us01_n731 ) , .B2( us01_n748 ) );
  NAND2_X1 us01_U333 (.A1( us01_n697 ) , .A2( us01_n727 ) , .ZN( us01_n780 ) );
  NOR2_X1 us01_U334 (.ZN( us01_n468 ) , .A2( us01_n777 ) , .A1( us01_n813 ) );
  NOR2_X1 us01_U335 (.ZN( us01_n516 ) , .A1( us01_n706 ) , .A2( us01_n786 ) );
  NAND2_X2 us01_U336 (.A2( us01_n447 ) , .A1( us01_n450 ) , .ZN( us01_n761 ) );
  OAI21_X1 us01_U337 (.A( us01_n696 ) , .ZN( us01_n700 ) , .B2( us01_n748 ) , .B1( us01_n802 ) );
  OAI21_X1 us01_U338 (.ZN( us01_n696 ) , .B2( us01_n831 ) , .B1( us01_n836 ) , .A( us01_n858 ) );
  NOR2_X1 us01_U339 (.ZN( us01_n524 ) , .A1( us01_n722 ) , .A2( us01_n748 ) );
  NOR4_X1 us01_U34 (.A4( us01_n791 ) , .A3( us01_n792 ) , .A2( us01_n793 ) , .A1( us01_n794 ) , .ZN( us01_n795 ) );
  AOI21_X1 us01_U340 (.ZN( us01_n441 ) , .B1( us01_n787 ) , .B2( us01_n789 ) , .A( us01_n812 ) );
  AOI21_X1 us01_U341 (.ZN( us01_n495 ) , .A( us01_n777 ) , .B2( us01_n789 ) , .B1( us01_n802 ) );
  NAND2_X1 us01_U342 (.ZN( us01_n712 ) , .A1( us01_n726 ) , .A2( us01_n778 ) );
  NOR2_X1 us01_U343 (.ZN( us01_n482 ) , .A1( us01_n786 ) , .A2( us01_n803 ) );
  NAND2_X1 us01_U344 (.A2( us01_n760 ) , .A1( us01_n804 ) , .ZN( us01_n808 ) );
  OAI21_X1 us01_U345 (.A( us01_n785 ) , .B2( us01_n786 ) , .B1( us01_n787 ) , .ZN( us01_n793 ) );
  OAI21_X1 us01_U346 (.ZN( us01_n785 ) , .A( us01_n837 ) , .B1( us01_n861 ) , .B2( us01_n871 ) );
  INV_X1 us01_U347 (.A( us01_n783 ) , .ZN( us01_n844 ) );
  NOR2_X1 us01_U348 (.ZN( us01_n710 ) , .A2( us01_n722 ) , .A1( us01_n788 ) );
  NAND2_X1 us01_U349 (.ZN( us01_n669 ) , .A1( us01_n804 ) , .A2( us01_n814 ) );
  NOR4_X1 us01_U35 (.A4( us01_n774 ) , .A3( us01_n775 ) , .A1( us01_n776 ) , .ZN( us01_n797 ) , .A2( us01_n799 ) );
  NAND2_X2 us01_U350 (.A2( us01_n446 ) , .A1( us01_n450 ) , .ZN( us01_n727 ) );
  INV_X1 us01_U351 (.A( us01_n722 ) , .ZN( us01_n854 ) );
  NAND2_X2 us01_U352 (.A1( us01_n445 ) , .A2( us01_n463 ) , .ZN( us01_n747 ) );
  INV_X1 us01_U353 (.A( us01_n815 ) , .ZN( us01_n842 ) );
  AND2_X1 us01_U354 (.ZN( us01_n730 ) , .A1( us01_n777 ) , .A2( us01_n783 ) );
  NAND2_X1 us01_U355 (.A1( us01_n445 ) , .A2( us01_n447 ) , .ZN( us01_n803 ) );
  NAND2_X1 us01_U356 (.A1( us01_n449 ) , .A2( us01_n452 ) , .ZN( us01_n812 ) );
  NAND2_X1 us01_U357 (.A1( us01_n453 ) , .A2( us01_n469 ) , .ZN( us01_n801 ) );
  NAND2_X1 us01_U358 (.A1( us01_n453 ) , .A2( us01_n460 ) , .ZN( us01_n748 ) );
  NAND2_X2 us01_U359 (.A2( us01_n446 ) , .A1( us01_n458 ) , .ZN( us01_n726 ) );
  NOR2_X1 us01_U36 (.ZN( us01_n802 ) , .A1( us01_n852 ) , .A2( us01_n859 ) );
  NAND2_X1 us01_U360 (.A2( us01_n451 ) , .A1( us01_n453 ) , .ZN( us01_n804 ) );
  NAND2_X1 us01_U361 (.A1( us01_n449 ) , .A2( us01_n469 ) , .ZN( us01_n814 ) );
  NAND2_X1 us01_U362 (.A1( us01_n452 ) , .A2( us01_n459 ) , .ZN( us01_n811 ) );
  NAND2_X1 us01_U363 (.A1( us01_n451 ) , .A2( us01_n459 ) , .ZN( us01_n742 ) );
  NAND2_X1 us01_U364 (.A1( us01_n451 ) , .A2( us01_n470 ) , .ZN( us01_n783 ) );
  NAND2_X1 us01_U365 (.A2( us01_n452 ) , .A1( us01_n470 ) , .ZN( us01_n777 ) );
  NAND2_X1 us01_U366 (.A2( us01_n459 ) , .A1( us01_n460 ) , .ZN( us01_n745 ) );
  NAND2_X2 us01_U367 (.A2( us01_n446 ) , .A1( us01_n462 ) , .ZN( us01_n813 ) );
  NAND2_X1 us01_U368 (.A1( us01_n460 ) , .A2( us01_n470 ) , .ZN( us01_n786 ) );
  NOR2_X1 us01_U369 (.ZN( us01_n451 ) , .A1( us01_n824 ) , .A2( us01_n825 ) );
  NAND4_X1 us01_U37 (.ZN( sa01_sr_2 ) , .A4( us01_n641 ) , .A3( us01_n642 ) , .A2( us01_n643 ) , .A1( us01_n644 ) );
  NOR2_X1 us01_U370 (.ZN( us01_n449 ) , .A1( us01_n826 ) , .A2( us01_n827 ) );
  NAND2_X1 us01_U371 (.A1( us01_n449 ) , .A2( us01_n460 ) , .ZN( us01_n788 ) );
  NAND2_X2 us01_U372 (.A1( us01_n447 ) , .A2( us01_n458 ) , .ZN( us01_n790 ) );
  NAND2_X2 us01_U373 (.A2( us01_n439 ) , .A1( us01_n450 ) , .ZN( us01_n789 ) );
  NAND2_X1 us01_U374 (.A2( us01_n452 ) , .A1( us01_n453 ) , .ZN( us01_n728 ) );
  NAND2_X2 us01_U375 (.A2( us01_n469 ) , .A1( us01_n470 ) , .ZN( us01_n815 ) );
  NAND2_X1 us01_U376 (.A1( us01_n445 ) , .A2( us01_n446 ) , .ZN( us01_n784 ) );
  NAND2_X2 us01_U377 (.A2( us01_n439 ) , .A1( us01_n445 ) , .ZN( us01_n782 ) );
  NOR2_X1 us01_U378 (.A2( sa01_7 ) , .ZN( us01_n458 ) , .A1( us01_n847 ) );
  NOR2_X1 us01_U379 (.A2( sa01_2 ) , .A1( sa01_3 ) , .ZN( us01_n470 ) );
  AOI222_X1 us01_U38 (.B2( us01_n636 ) , .ZN( us01_n642 ) , .B1( us01_n839 ) , .A1( us01_n840 ) , .C2( us01_n844 ) , .C1( us01_n861 ) , .A2( us01_n863 ) );
  NOR2_X1 us01_U380 (.A2( sa01_1 ) , .ZN( us01_n469 ) , .A1( us01_n824 ) );
  NOR2_X1 us01_U381 (.A2( sa01_0 ) , .ZN( us01_n452 ) , .A1( us01_n825 ) );
  NOR2_X1 us01_U382 (.A2( sa01_0 ) , .A1( sa01_1 ) , .ZN( us01_n460 ) );
  NAND2_X2 us01_U383 (.A1( us01_n439 ) , .A2( us01_n458 ) , .ZN( us01_n697 ) );
  NOR2_X1 us01_U384 (.A2( sa01_3 ) , .ZN( us01_n453 ) , .A1( us01_n826 ) );
  NOR2_X1 us01_U385 (.A2( sa01_2 ) , .ZN( us01_n459 ) , .A1( us01_n827 ) );
  INV_X1 us01_U386 (.A( sa01_3 ) , .ZN( us01_n827 ) );
  INV_X1 us01_U387 (.A( sa01_1 ) , .ZN( us01_n825 ) );
  INV_X1 us01_U388 (.A( sa01_0 ) , .ZN( us01_n824 ) );
  INV_X1 us01_U389 (.A( sa01_2 ) , .ZN( us01_n826 ) );
  NOR4_X1 us01_U39 (.A4( us01_n637 ) , .A3( us01_n638 ) , .A2( us01_n639 ) , .A1( us01_n640 ) , .ZN( us01_n641 ) );
  INV_X1 us01_U390 (.A( sa01_5 ) , .ZN( us01_n846 ) );
  NAND2_X1 us01_U391 (.A1( us01_n727 ) , .A2( us01_n782 ) , .ZN( us01_n809 ) );
  OAI22_X1 us01_U392 (.ZN( us01_n586 ) , .A2( us01_n745 ) , .B2( us01_n760 ) , .A1( us01_n761 ) , .B1( us01_n782 ) );
  AOI21_X1 us01_U393 (.ZN( us01_n590 ) , .B1( us01_n726 ) , .B2( us01_n782 ) , .A( us01_n788 ) );
  AOI21_X1 us01_U394 (.ZN( us01_n646 ) , .A( us01_n760 ) , .B2( us01_n782 ) , .B1( us01_n790 ) );
  AOI21_X1 us01_U395 (.ZN( us01_n621 ) , .B1( us01_n697 ) , .A( us01_n777 ) , .B2( us01_n782 ) );
  OAI22_X1 us01_U396 (.ZN( us01_n679 ) , .A1( us01_n697 ) , .A2( us01_n728 ) , .B2( us01_n782 ) , .B1( us01_n815 ) );
  OAI21_X1 us01_U397 (.A( us01_n611 ) , .ZN( us01_n614 ) , .B1( us01_n623 ) , .B2( us01_n782 ) );
  NOR2_X1 us01_U398 (.ZN( us01_n608 ) , .A1( us01_n782 ) , .A2( us01_n814 ) );
  INV_X2 us01_U399 (.A( us01_n747 ) , .ZN( us01_n861 ) );
  NAND2_X2 us01_U4 (.A1( us01_n439 ) , .A2( us01_n462 ) , .ZN( us01_n706 ) );
  NOR3_X1 us01_U40 (.A2( us01_n605 ) , .A1( us01_n606 ) , .ZN( us01_n644 ) , .A3( us01_n720 ) );
  OAI222_X1 us01_U400 (.A2( us01_n667 ) , .ZN( us01_n672 ) , .B1( us01_n745 ) , .B2( us01_n782 ) , .C2( us01_n786 ) , .C1( us01_n813 ) , .A1( us01_n815 ) );
  NOR2_X1 us01_U401 (.ZN( us01_n649 ) , .A1( us01_n782 ) , .A2( us01_n786 ) );
  NOR2_X1 us01_U402 (.ZN( us01_n598 ) , .A2( us01_n695 ) , .A1( us01_n782 ) );
  NOR2_X1 us01_U403 (.ZN( us01_n551 ) , .A2( us01_n742 ) , .A1( us01_n782 ) );
  INV_X1 us01_U404 (.A( us01_n782 ) , .ZN( us01_n859 ) );
  NAND2_X1 us01_U405 (.A2( us01_n459 ) , .A1( us01_n469 ) , .ZN( us01_n695 ) );
  INV_X1 us01_U406 (.A( sa01_7 ) , .ZN( us01_n856 ) );
  OAI221_X1 us01_U407 (.A( us01_n781 ) , .C2( us01_n782 ) , .B2( us01_n783 ) , .B1( us01_n784 ) , .ZN( us01_n794 ) , .C1( us01_n811 ) );
  AOI21_X1 us01_U408 (.ZN( us01_n498 ) , .A( us01_n695 ) , .B1( us01_n706 ) , .B2( us01_n784 ) );
  OAI221_X1 us01_U409 (.A( us01_n694 ) , .ZN( us01_n701 ) , .C2( us01_n782 ) , .C1( us01_n783 ) , .B1( us01_n784 ) , .B2( us01_n804 ) );
  NAND4_X1 us01_U41 (.ZN( sa01_sr_7 ) , .A4( us01_n820 ) , .A3( us01_n821 ) , .A2( us01_n822 ) , .A1( us01_n823 ) );
  OAI22_X1 us01_U410 (.ZN( us01_n588 ) , .B1( us01_n728 ) , .B2( us01_n747 ) , .A2( us01_n784 ) , .A1( us01_n801 ) );
  AOI222_X1 us01_U411 (.ZN( us01_n511 ) , .C1( us01_n830 ) , .B2( us01_n835 ) , .A2( us01_n841 ) , .C2( us01_n860 ) , .B1( us01_n861 ) , .A1( us01_n864 ) );
  AOI222_X1 us01_U412 (.ZN( us01_n603 ) , .B2( us01_n669 ) , .B1( us01_n751 ) , .C2( us01_n829 ) , .A1( us01_n831 ) , .A2( us01_n860 ) , .C1( us01_n861 ) );
  AOI221_X1 us01_U413 (.A( us01_n481 ) , .ZN( us01_n486 ) , .B1( us01_n829 ) , .C2( us01_n842 ) , .C1( us01_n850 ) , .B2( us01_n860 ) );
  NAND2_X1 us01_U414 (.A2( us01_n747 ) , .A1( us01_n784 ) , .ZN( us01_n807 ) );
  NOR2_X1 us01_U415 (.ZN( us01_n610 ) , .A1( us01_n777 ) , .A2( us01_n784 ) );
  NOR2_X1 us01_U416 (.ZN( us01_n715 ) , .A2( us01_n742 ) , .A1( us01_n784 ) );
  OAI222_X1 us01_U417 (.ZN( us01_n615 ) , .B1( us01_n695 ) , .C1( us01_n722 ) , .C2( us01_n745 ) , .B2( us01_n784 ) , .A2( us01_n790 ) , .A1( us01_n814 ) );
  NOR2_X1 us01_U418 (.ZN( us01_n651 ) , .A1( us01_n760 ) , .A2( us01_n784 ) );
  NOR2_X1 us01_U419 (.ZN( us01_n552 ) , .A1( us01_n784 ) , .A2( us01_n811 ) );
  AOI222_X1 us01_U42 (.C2( us01_n807 ) , .B2( us01_n808 ) , .A2( us01_n809 ) , .ZN( us01_n821 ) , .C1( us01_n830 ) , .A1( us01_n837 ) , .B1( us01_n851 ) );
  NOR2_X1 us01_U420 (.ZN( us01_n787 ) , .A2( us01_n860 ) , .A1( us01_n866 ) );
  NOR2_X1 us01_U421 (.ZN( us01_n699 ) , .A2( us01_n784 ) , .A1( us01_n815 ) );
  NOR2_X1 us01_U422 (.A1( us01_n728 ) , .ZN( us01_n763 ) , .A2( us01_n784 ) );
  INV_X1 us01_U423 (.A( us01_n784 ) , .ZN( us01_n860 ) );
  NOR2_X1 us01_U424 (.A2( sa01_4 ) , .ZN( us01_n447 ) , .A1( us01_n846 ) );
  NOR2_X1 us01_U425 (.ZN( us01_n463 ) , .A2( us01_n845 ) , .A1( us01_n846 ) );
  NOR2_X1 us01_U426 (.A2( sa01_5 ) , .ZN( us01_n446 ) , .A1( us01_n845 ) );
  NOR2_X1 us01_U427 (.A2( sa01_4 ) , .A1( sa01_5 ) , .ZN( us01_n439 ) );
  INV_X1 us01_U428 (.A( sa01_6 ) , .ZN( us01_n847 ) );
  NOR2_X1 us01_U429 (.ZN( us01_n445 ) , .A2( us01_n847 ) , .A1( us01_n856 ) );
  NOR4_X1 us01_U43 (.A4( us01_n816 ) , .A3( us01_n817 ) , .A2( us01_n818 ) , .A1( us01_n819 ) , .ZN( us01_n820 ) );
  NOR2_X1 us01_U430 (.A2( sa01_6 ) , .ZN( us01_n450 ) , .A1( us01_n856 ) );
  NOR2_X1 us01_U431 (.A2( sa01_6 ) , .A1( sa01_7 ) , .ZN( us01_n462 ) );
  AOI221_X1 us01_U432 (.A( us01_n574 ) , .ZN( us01_n585 ) , .B2( us01_n829 ) , .C2( us01_n841 ) , .B1( us01_n852 ) , .C1( us01_n859 ) );
  AOI21_X1 us01_U433 (.ZN( us01_n574 ) , .B2( us01_n722 ) , .B1( us01_n746 ) , .A( us01_n783 ) );
  INV_X1 us01_U434 (.A( sa01_4 ) , .ZN( us01_n845 ) );
  AOI211_X1 us01_U435 (.A( us01_n635 ) , .ZN( us01_n643 ) , .B( us01_n741 ) , .C2( us01_n837 ) , .C1( us01_n852 ) );
  NAND4_X1 us01_U436 (.A4( us01_n631 ) , .A3( us01_n632 ) , .A2( us01_n633 ) , .A1( us01_n634 ) , .ZN( us01_n741 ) );
  NAND3_X1 us01_U437 (.ZN( sa01_sr_6 ) , .A3( us01_n795 ) , .A2( us01_n796 ) , .A1( us01_n797 ) );
  NAND3_X1 us01_U438 (.ZN( sa01_sr_5 ) , .A3( us01_n756 ) , .A2( us01_n757 ) , .A1( us01_n758 ) );
  NAND3_X1 us01_U439 (.ZN( sa01_sr_4 ) , .A3( us01_n736 ) , .A2( us01_n737 ) , .A1( us01_n738 ) );
  AOI211_X1 us01_U44 (.B( us01_n805 ) , .A( us01_n806 ) , .ZN( us01_n822 ) , .C1( us01_n840 ) , .C2( us01_n848 ) );
  NAND3_X1 us01_U440 (.A3( us01_n673 ) , .A2( us01_n674 ) , .A1( us01_n675 ) , .ZN( us01_n805 ) );
  NAND3_X1 us01_U441 (.ZN( us01_n636 ) , .A3( us01_n706 ) , .A2( us01_n722 ) , .A1( us01_n790 ) );
  NAND3_X1 us01_U442 (.A3( us01_n616 ) , .A2( us01_n617 ) , .A1( us01_n618 ) , .ZN( us01_n723 ) );
  NAND3_X1 us01_U443 (.A3( us01_n583 ) , .A2( us01_n584 ) , .A1( us01_n585 ) , .ZN( us01_n619 ) );
  NAND3_X1 us01_U444 (.ZN( us01_n563 ) , .A3( us01_n678 ) , .A2( us01_n748 ) , .A1( us01_n783 ) );
  NAND3_X1 us01_U445 (.A3( us01_n521 ) , .A2( us01_n522 ) , .A1( us01_n523 ) , .ZN( us01_n740 ) );
  NAND3_X1 us01_U446 (.A3( us01_n510 ) , .A1( us01_n511 ) , .ZN( us01_n606 ) , .A2( us01_n869 ) );
  NAND3_X1 us01_U447 (.A3( us01_n465 ) , .A2( us01_n466 ) , .A1( us01_n467 ) , .ZN( us01_n775 ) );
  NAND4_X1 us01_U45 (.ZN( sa01_sr_0 ) , .A4( us01_n499 ) , .A3( us01_n500 ) , .A2( us01_n501 ) , .A1( us01_n502 ) );
  NOR4_X1 us01_U46 (.A4( us01_n496 ) , .A3( us01_n497 ) , .A2( us01_n498 ) , .ZN( us01_n499 ) , .A1( us01_n525 ) );
  AOI221_X1 us01_U47 (.A( us01_n495 ) , .ZN( us01_n500 ) , .B2( us01_n841 ) , .C1( us01_n844 ) , .C2( us01_n858 ) , .B1( us01_n860 ) );
  AOI211_X1 us01_U48 (.A( us01_n494 ) , .ZN( us01_n501 ) , .B( us01_n800 ) , .C2( us01_n837 ) , .C1( us01_n849 ) );
  NOR2_X1 us01_U49 (.ZN( us01_n746 ) , .A1( us01_n859 ) , .A2( us01_n860 ) );
  NAND2_X2 us01_U5 (.A2( us01_n458 ) , .A1( us01_n463 ) , .ZN( us01_n778 ) );
  NAND4_X1 us01_U50 (.ZN( sa01_sr_1 ) , .A4( us01_n593 ) , .A3( us01_n594 ) , .A2( us01_n595 ) , .A1( us01_n596 ) );
  AOI211_X1 us01_U51 (.B( us01_n587 ) , .A( us01_n588 ) , .ZN( us01_n594 ) , .C2( us01_n809 ) , .C1( us01_n831 ) );
  NOR4_X1 us01_U52 (.A4( us01_n589 ) , .A3( us01_n590 ) , .A2( us01_n591 ) , .A1( us01_n592 ) , .ZN( us01_n593 ) );
  AOI211_X1 us01_U53 (.A( us01_n586 ) , .ZN( us01_n595 ) , .B( us01_n619 ) , .C1( us01_n843 ) , .C2( us01_n853 ) );
  NOR2_X1 us01_U54 (.ZN( us01_n623 ) , .A2( us01_n834 ) , .A1( us01_n837 ) );
  NAND4_X1 us01_U55 (.A4( us01_n601 ) , .A3( us01_n602 ) , .A2( us01_n603 ) , .A1( us01_n604 ) , .ZN( us01_n720 ) );
  NOR3_X1 us01_U56 (.A1( us01_n597 ) , .ZN( us01_n602 ) , .A3( us01_n661 ) , .A2( us01_n768 ) );
  NOR4_X1 us01_U57 (.A3( us01_n598 ) , .A2( us01_n599 ) , .A1( us01_n600 ) , .ZN( us01_n601 ) , .A4( us01_n653 ) );
  AOI222_X1 us01_U58 (.ZN( us01_n604 ) , .A1( us01_n828 ) , .C2( us01_n835 ) , .B1( us01_n840 ) , .A2( us01_n854 ) , .B2( us01_n859 ) , .C1( us01_n866 ) );
  NOR4_X1 us01_U59 (.A4( us01_n575 ) , .A3( us01_n576 ) , .A2( us01_n577 ) , .ZN( us01_n584 ) , .A1( us01_n681 ) );
  INV_X1 us01_U6 (.A( us01_n667 ) , .ZN( us01_n863 ) );
  NOR4_X1 us01_U60 (.A1( us01_n582 ) , .ZN( us01_n583 ) , .A3( us01_n650 ) , .A2( us01_n660 ) , .A4( us01_n765 ) );
  NAND4_X1 us01_U61 (.A4( us01_n483 ) , .A3( us01_n484 ) , .A2( us01_n485 ) , .A1( us01_n486 ) , .ZN( us01_n776 ) );
  NOR4_X1 us01_U62 (.A4( us01_n482 ) , .ZN( us01_n485 ) , .A1( us01_n564 ) , .A2( us01_n579 ) , .A3( us01_n600 ) );
  NOR4_X1 us01_U63 (.ZN( us01_n483 ) , .A2( us01_n531 ) , .A1( us01_n556 ) , .A3( us01_n629 ) , .A4( us01_n716 ) );
  NOR4_X1 us01_U64 (.ZN( us01_n484 ) , .A1( us01_n505 ) , .A2( us01_n517 ) , .A4( us01_n544 ) , .A3( us01_n609 ) );
  NOR4_X1 us01_U65 (.A4( us01_n627 ) , .A3( us01_n628 ) , .A2( us01_n629 ) , .A1( us01_n630 ) , .ZN( us01_n631 ) );
  AOI211_X1 us01_U66 (.B( us01_n621 ) , .A( us01_n622 ) , .ZN( us01_n633 ) , .C2( us01_n834 ) , .C1( us01_n861 ) );
  NOR4_X1 us01_U67 (.A4( us01_n624 ) , .A3( us01_n625 ) , .A2( us01_n626 ) , .ZN( us01_n632 ) , .A1( us01_n662 ) );
  NAND4_X1 us01_U68 (.A4( us01_n655 ) , .A3( us01_n656 ) , .A2( us01_n657 ) , .A1( us01_n658 ) , .ZN( us01_n798 ) );
  NOR3_X1 us01_U69 (.A3( us01_n649 ) , .A2( us01_n650 ) , .A1( us01_n651 ) , .ZN( us01_n656 ) );
  NOR3_X1 us01_U7 (.ZN( us01_n596 ) , .A1( us01_n606 ) , .A3( us01_n721 ) , .A2( us01_n740 ) );
  NOR3_X1 us01_U70 (.A3( us01_n652 ) , .A2( us01_n653 ) , .A1( us01_n654 ) , .ZN( us01_n655 ) );
  NOR3_X1 us01_U71 (.A3( us01_n646 ) , .A2( us01_n647 ) , .A1( us01_n648 ) , .ZN( us01_n657 ) );
  NAND4_X1 us01_U72 (.A4( us01_n558 ) , .A3( us01_n559 ) , .A2( us01_n560 ) , .A1( us01_n561 ) , .ZN( us01_n605 ) );
  NOR4_X1 us01_U73 (.ZN( us01_n559 ) , .A1( us01_n651 ) , .A3( us01_n659 ) , .A4( us01_n683 ) , .A2( us01_n766 ) );
  NOR4_X1 us01_U74 (.A4( us01_n550 ) , .A3( us01_n551 ) , .A2( us01_n552 ) , .A1( us01_n553 ) , .ZN( us01_n560 ) );
  NOR4_X1 us01_U75 (.A4( us01_n554 ) , .A3( us01_n555 ) , .A2( us01_n556 ) , .A1( us01_n557 ) , .ZN( us01_n558 ) );
  NAND4_X1 us01_U76 (.A4( us01_n770 ) , .A3( us01_n771 ) , .A2( us01_n772 ) , .A1( us01_n773 ) , .ZN( us01_n799 ) );
  NOR3_X1 us01_U77 (.A3( us01_n763 ) , .A2( us01_n764 ) , .A1( us01_n765 ) , .ZN( us01_n771 ) );
  NOR4_X1 us01_U78 (.A4( us01_n766 ) , .A3( us01_n767 ) , .A2( us01_n768 ) , .A1( us01_n769 ) , .ZN( us01_n770 ) );
  AOI222_X1 us01_U79 (.ZN( us01_n773 ) , .A1( us01_n828 ) , .C1( us01_n832 ) , .B2( us01_n839 ) , .A2( us01_n848 ) , .B1( us01_n859 ) , .C2( us01_n871 ) );
  NOR3_X1 us01_U8 (.A3( us01_n798 ) , .A2( us01_n799 ) , .A1( us01_n800 ) , .ZN( us01_n823 ) );
  NOR4_X1 us01_U80 (.A4( us01_n507 ) , .A2( us01_n508 ) , .A1( us01_n509 ) , .ZN( us01_n510 ) , .A3( us01_n668 ) );
  INV_X1 us01_U81 (.A( us01_n503 ) , .ZN( us01_n869 ) );
  NOR4_X1 us01_U82 (.A4( us01_n663 ) , .A3( us01_n664 ) , .A2( us01_n665 ) , .A1( us01_n666 ) , .ZN( us01_n674 ) );
  NOR4_X1 us01_U83 (.A4( us01_n659 ) , .A3( us01_n660 ) , .A2( us01_n661 ) , .A1( us01_n662 ) , .ZN( us01_n675 ) );
  NOR4_X1 us01_U84 (.A3( us01_n671 ) , .A1( us01_n672 ) , .ZN( us01_n673 ) , .A4( us01_n713 ) , .A2( us01_n857 ) );
  NOR2_X1 us01_U85 (.ZN( us01_n759 ) , .A1( us01_n831 ) , .A2( us01_n832 ) );
  NAND4_X1 us01_U86 (.A4( us01_n454 ) , .A3( us01_n455 ) , .A2( us01_n456 ) , .A1( us01_n457 ) , .ZN( us01_n677 ) );
  NOR3_X1 us01_U87 (.ZN( us01_n455 ) , .A3( us01_n528 ) , .A1( us01_n553 ) , .A2( us01_n568 ) );
  AOI221_X1 us01_U88 (.A( us01_n448 ) , .ZN( us01_n457 ) , .C2( us01_n751 ) , .B1( us01_n830 ) , .C1( us01_n840 ) , .B2( us01_n859 ) );
  NOR4_X1 us01_U89 (.ZN( us01_n456 ) , .A2( us01_n507 ) , .A1( us01_n597 ) , .A4( us01_n626 ) , .A3( us01_n709 ) );
  NOR3_X1 us01_U9 (.A3( us01_n619 ) , .A2( us01_n620 ) , .ZN( us01_n634 ) , .A1( us01_n723 ) );
  NAND4_X1 us01_U90 (.A4( us01_n533 ) , .A3( us01_n534 ) , .A2( us01_n535 ) , .A1( us01_n536 ) , .ZN( us01_n620 ) );
  NOR4_X1 us01_U91 (.A4( us01_n524 ) , .A2( us01_n525 ) , .A1( us01_n526 ) , .ZN( us01_n536 ) , .A3( us01_n699 ) );
  NOR4_X1 us01_U92 (.A1( us01_n529 ) , .ZN( us01_n534 ) , .A2( us01_n652 ) , .A4( us01_n666 ) , .A3( us01_n763 ) );
  NOR4_X1 us01_U93 (.A4( us01_n527 ) , .A3( us01_n528 ) , .ZN( us01_n535 ) , .A2( us01_n682 ) , .A1( us01_n792 ) );
  NAND4_X1 us01_U94 (.A4( us01_n477 ) , .A3( us01_n478 ) , .A2( us01_n479 ) , .A1( us01_n480 ) , .ZN( us01_n692 ) );
  NOR3_X1 us01_U95 (.ZN( us01_n478 ) , .A2( us01_n506 ) , .A3( us01_n599 ) , .A1( us01_n608 ) );
  AOI211_X1 us01_U96 (.B( us01_n475 ) , .A( us01_n476 ) , .ZN( us01_n480 ) , .C2( us01_n831 ) , .C1( us01_n859 ) );
  NOR4_X1 us01_U97 (.ZN( us01_n479 ) , .A3( us01_n530 ) , .A4( us01_n543 ) , .A2( us01_n565 ) , .A1( us01_n715 ) );
  NAND4_X1 us01_U98 (.A4( us01_n546 ) , .A3( us01_n547 ) , .A2( us01_n548 ) , .A1( us01_n549 ) , .ZN( us01_n743 ) );
  NOR3_X1 us01_U99 (.ZN( us01_n547 ) , .A2( us01_n649 ) , .A1( us01_n665 ) , .A3( us01_n769 ) );
  NOR2_X1 us10_U10 (.A1( us10_n678 ) , .ZN( us10_n693 ) , .A2( us10_n807 ) );
  NOR3_X1 us10_U100 (.ZN( us10_n549 ) , .A2( us10_n651 ) , .A1( us10_n667 ) , .A3( us10_n771 ) );
  AOI211_X1 us10_U101 (.B( us10_n539 ) , .A( us10_n540 ) , .ZN( us10_n551 ) , .C2( us10_n839 ) , .C1( us10_n851 ) );
  NOR4_X1 us10_U102 (.A4( us10_n544 ) , .A3( us10_n545 ) , .A2( us10_n546 ) , .A1( us10_n547 ) , .ZN( us10_n548 ) );
  NOR4_X1 us10_U103 (.ZN( us10_n620 ) , .A1( us10_n656 ) , .A3( us10_n666 ) , .A4( us10_n682 ) , .A2( us10_n766 ) );
  NOR4_X1 us10_U104 (.A4( us10_n609 ) , .A3( us10_n610 ) , .A2( us10_n611 ) , .A1( us10_n612 ) , .ZN( us10_n619 ) );
  NOR4_X1 us10_U105 (.A4( us10_n614 ) , .A3( us10_n615 ) , .A2( us10_n616 ) , .A1( us10_n617 ) , .ZN( us10_n618 ) );
  NAND4_X1 us10_U106 (.A4( us10_n485 ) , .A3( us10_n486 ) , .A2( us10_n487 ) , .A1( us10_n488 ) , .ZN( us10_n778 ) );
  NOR4_X1 us10_U107 (.A4( us10_n484 ) , .ZN( us10_n487 ) , .A1( us10_n566 ) , .A2( us10_n581 ) , .A3( us10_n602 ) );
  NOR4_X1 us10_U108 (.ZN( us10_n486 ) , .A1( us10_n507 ) , .A2( us10_n519 ) , .A4( us10_n546 ) , .A3( us10_n611 ) );
  NOR4_X1 us10_U109 (.ZN( us10_n485 ) , .A2( us10_n533 ) , .A1( us10_n558 ) , .A3( us10_n631 ) , .A4( us10_n718 ) );
  INV_X1 us10_U11 (.A( us10_n680 ) , .ZN( us10_n840 ) );
  NAND4_X1 us10_U110 (.A4( us10_n691 ) , .A3( us10_n692 ) , .A1( us10_n693 ) , .ZN( us10_n776 ) , .A2( us10_n872 ) );
  AOI221_X1 us10_U111 (.A( us10_n681 ) , .ZN( us10_n692 ) , .B2( us10_n840 ) , .C1( us10_n842 ) , .C2( us10_n862 ) , .B1( us10_n865 ) );
  INV_X1 us10_U112 (.A( us10_n679 ) , .ZN( us10_n872 ) );
  NOR4_X1 us10_U113 (.A4( us10_n687 ) , .A3( us10_n688 ) , .A2( us10_n689 ) , .A1( us10_n690 ) , .ZN( us10_n691 ) );
  NAND4_X1 us10_U114 (.A4( us10_n473 ) , .A3( us10_n474 ) , .A2( us10_n475 ) , .A1( us10_n476 ) , .ZN( us10_n678 ) );
  NOR4_X1 us10_U115 (.A4( us10_n470 ) , .ZN( us10_n476 ) , .A3( us10_n556 ) , .A1( us10_n735 ) , .A2( us10_n755 ) );
  NOR4_X1 us10_U116 (.ZN( us10_n475 ) , .A1( us10_n531 ) , .A3( us10_n568 ) , .A4( us10_n600 ) , .A2( us10_n642 ) );
  NOR4_X1 us10_U117 (.ZN( us10_n474 ) , .A1( us10_n506 ) , .A3( us10_n544 ) , .A2( us10_n583 ) , .A4( us10_n716 ) );
  NAND4_X1 us10_U118 (.A4( us10_n719 ) , .A3( us10_n720 ) , .A2( us10_n721 ) , .ZN( us10_n741 ) , .A1( us10_n857 ) );
  INV_X1 us10_U119 (.A( us10_n709 ) , .ZN( us10_n857 ) );
  NOR4_X1 us10_U12 (.A4( us10_n445 ) , .A3( us10_n446 ) , .A2( us10_n516 ) , .A1( us10_n541 ) , .ZN( us10_n706 ) );
  NOR4_X1 us10_U120 (.A4( us10_n715 ) , .A3( us10_n716 ) , .A2( us10_n717 ) , .A1( us10_n718 ) , .ZN( us10_n719 ) );
  AOI221_X1 us10_U121 (.A( us10_n710 ) , .ZN( us10_n721 ) , .C2( us10_n844 ) , .B2( us10_n845 ) , .C1( us10_n861 ) , .B1( us10_n862 ) );
  NOR2_X1 us10_U122 (.ZN( us10_n789 ) , .A2( us10_n862 ) , .A1( us10_n868 ) );
  NOR2_X1 us10_U123 (.ZN( us10_n733 ) , .A2( us10_n832 ) , .A1( us10_n845 ) );
  NAND4_X1 us10_U124 (.A4( us10_n573 ) , .A3( us10_n574 ) , .A1( us10_n575 ) , .ZN( us10_n723 ) , .A2( us10_n874 ) );
  NOR4_X1 us10_U125 (.A4( us10_n569 ) , .A3( us10_n570 ) , .A2( us10_n571 ) , .A1( us10_n572 ) , .ZN( us10_n573 ) );
  AOI221_X1 us10_U126 (.A( us10_n564 ) , .C2( us10_n565 ) , .ZN( us10_n574 ) , .B2( us10_n845 ) , .B1( us10_n852 ) , .C1( us10_n853 ) );
  INV_X1 us10_U127 (.A( us10_n607 ) , .ZN( us10_n874 ) );
  NAND4_X1 us10_U128 (.A4( us10_n633 ) , .A3( us10_n634 ) , .A2( us10_n635 ) , .A1( us10_n636 ) , .ZN( us10_n743 ) );
  AOI211_X1 us10_U129 (.B( us10_n623 ) , .A( us10_n624 ) , .ZN( us10_n635 ) , .C2( us10_n836 ) , .C1( us10_n863 ) );
  OR3_X1 us10_U13 (.ZN( us10_n446 ) , .A1( us10_n528 ) , .A3( us10_n577 ) , .A2( us10_n875 ) );
  NOR4_X1 us10_U130 (.A4( us10_n629 ) , .A3( us10_n630 ) , .A2( us10_n631 ) , .A1( us10_n632 ) , .ZN( us10_n633 ) );
  NOR4_X1 us10_U131 (.A4( us10_n626 ) , .A3( us10_n627 ) , .A2( us10_n628 ) , .ZN( us10_n634 ) , .A1( us10_n664 ) );
  NAND4_X1 us10_U132 (.A4( us10_n493 ) , .A3( us10_n494 ) , .A1( us10_n495 ) , .ZN( us10_n802 ) , .A2( us10_n867 ) );
  AOI221_X1 us10_U133 (.A( us10_n489 ) , .ZN( us10_n494 ) , .B2( us10_n836 ) , .C2( us10_n841 ) , .C1( us10_n851 ) , .B1( us10_n860 ) );
  INV_X1 us10_U134 (.A( us10_n778 ) , .ZN( us10_n867 ) );
  NOR2_X1 us10_U135 (.ZN( us10_n495 ) , .A1( us10_n678 ) , .A2( us10_n694 ) );
  NOR2_X1 us10_U136 (.ZN( us10_n748 ) , .A1( us10_n861 ) , .A2( us10_n862 ) );
  NOR2_X1 us10_U137 (.ZN( us10_n647 ) , .A1( us10_n854 ) , .A2( us10_n868 ) );
  INV_X1 us10_U138 (.A( us10_n762 ) , .ZN( us10_n830 ) );
  OR4_X1 us10_U139 (.ZN( us10_n466 ) , .A4( us10_n518 ) , .A3( us10_n529 ) , .A2( us10_n578 ) , .A1( us10_n712 ) );
  OR4_X1 us10_U14 (.A4( us10_n442 ) , .A2( us10_n443 ) , .A1( us10_n444 ) , .ZN( us10_n445 ) , .A3( us10_n553 ) );
  OR4_X1 us10_U140 (.A4( us10_n566 ) , .A3( us10_n567 ) , .A2( us10_n568 ) , .ZN( us10_n572 ) , .A1( us10_n665 ) );
  OR4_X1 us10_U141 (.A4( us10_n518 ) , .A2( us10_n519 ) , .A1( us10_n520 ) , .ZN( us10_n522 ) , .A3( us10_n821 ) );
  OR4_X1 us10_U142 (.A4( us10_n682 ) , .A3( us10_n683 ) , .A2( us10_n684 ) , .A1( us10_n685 ) , .ZN( us10_n690 ) );
  OR4_X1 us10_U143 (.A4( us10_n580 ) , .A3( us10_n581 ) , .A2( us10_n582 ) , .A1( us10_n583 ) , .ZN( us10_n584 ) );
  NAND2_X1 us10_U144 (.ZN( us10_n613 ) , .A2( us10_n837 ) , .A1( us10_n873 ) );
  OR3_X1 us10_U145 (.A3( us10_n506 ) , .A2( us10_n507 ) , .A1( us10_n508 ) , .ZN( us10_n511 ) );
  INV_X1 us10_U146 (.A( us10_n672 ) , .ZN( us10_n859 ) );
  AOI21_X1 us10_U147 (.A( us10_n670 ) , .B1( us10_n671 ) , .ZN( us10_n672 ) , .B2( us10_n856 ) );
  INV_X1 us10_U148 (.A( us10_n754 ) , .ZN( us10_n869 ) );
  OAI21_X1 us10_U149 (.B1( us10_n753 ) , .ZN( us10_n754 ) , .A( us10_n845 ) , .B2( us10_n868 ) );
  INV_X1 us10_U15 (.A( us10_n613 ) , .ZN( us10_n875 ) );
  INV_X1 us10_U150 (.A( us10_n463 ) , .ZN( us10_n864 ) );
  OAI21_X1 us10_U151 (.ZN( us10_n463 ) , .B1( us10_n809 ) , .A( us10_n834 ) , .B2( us10_n851 ) );
  AOI222_X1 us10_U152 (.ZN( us10_n660 ) , .A2( us10_n839 ) , .B1( us10_n841 ) , .C2( us10_n845 ) , .A1( us10_n860 ) , .C1( us10_n863 ) , .B2( us10_n870 ) );
  INV_X1 us10_U153 (.A( us10_n647 ) , .ZN( us10_n870 ) );
  NAND2_X1 us10_U154 (.A1( us10_n447 ) , .A2( us10_n465 ) , .ZN( us10_n749 ) );
  OAI222_X1 us10_U155 (.B2( us10_n708 ) , .ZN( us10_n709 ) , .C2( us10_n724 ) , .B1( us10_n747 ) , .A1( us10_n806 ) , .C1( us10_n814 ) , .A2( us10_n815 ) );
  OAI222_X1 us10_U156 (.A2( us10_n669 ) , .ZN( us10_n674 ) , .B1( us10_n747 ) , .B2( us10_n784 ) , .C2( us10_n788 ) , .C1( us10_n815 ) , .A1( us10_n817 ) );
  OAI222_X1 us10_U157 (.ZN( us10_n617 ) , .B1( us10_n697 ) , .C1( us10_n724 ) , .C2( us10_n747 ) , .B2( us10_n786 ) , .A2( us10_n792 ) , .A1( us10_n816 ) );
  NOR4_X1 us10_U158 (.A2( us10_n491 ) , .A1( us10_n492 ) , .ZN( us10_n493 ) , .A3( us10_n580 ) , .A4( us10_n612 ) );
  OR4_X1 us10_U159 (.ZN( us10_n492 ) , .A4( us10_n534 ) , .A2( us10_n547 ) , .A1( us10_n559 ) , .A3( us10_n632 ) );
  INV_X1 us10_U16 (.A( us10_n749 ) , .ZN( us10_n863 ) );
  OAI22_X1 us10_U160 (.B1( us10_n490 ) , .ZN( us10_n491 ) , .A1( us10_n686 ) , .A2( us10_n763 ) , .B2( us10_n817 ) );
  NOR3_X1 us10_U161 (.ZN( us10_n490 ) , .A1( us10_n782 ) , .A2( us10_n850 ) , .A3( us10_n863 ) );
  INV_X1 us10_U162 (.A( us10_n730 ) , .ZN( us10_n839 ) );
  AOI221_X1 us10_U163 (.A( us10_n450 ) , .ZN( us10_n459 ) , .C2( us10_n753 ) , .B1( us10_n832 ) , .C1( us10_n842 ) , .B2( us10_n861 ) );
  AOI21_X1 us10_U164 (.ZN( us10_n450 ) , .B2( us10_n792 ) , .A( us10_n803 ) , .B1( us10_n815 ) );
  AOI221_X1 us10_U165 (.A( us10_n483 ) , .ZN( us10_n488 ) , .B1( us10_n831 ) , .C2( us10_n844 ) , .C1( us10_n852 ) , .B2( us10_n862 ) );
  OAI22_X1 us10_U166 (.ZN( us10_n483 ) , .A1( us10_n708 ) , .B2( us10_n785 ) , .A2( us10_n806 ) , .B1( us10_n812 ) );
  INV_X1 us10_U167 (.A( us10_n790 ) , .ZN( us10_n832 ) );
  NAND2_X1 us10_U168 (.A1( us10_n451 ) , .A2( us10_n453 ) , .ZN( us10_n762 ) );
  INV_X1 us10_U169 (.A( us10_n786 ) , .ZN( us10_n862 ) );
  AOI222_X1 us10_U17 (.ZN( us10_n605 ) , .B2( us10_n671 ) , .B1( us10_n753 ) , .C2( us10_n831 ) , .A1( us10_n833 ) , .A2( us10_n862 ) , .C1( us10_n863 ) );
  OAI221_X1 us10_U170 (.A( us10_n783 ) , .C2( us10_n784 ) , .B2( us10_n785 ) , .B1( us10_n786 ) , .ZN( us10_n796 ) , .C1( us10_n813 ) );
  AOI22_X1 us10_U171 (.A2( us10_n782 ) , .ZN( us10_n783 ) , .B2( us10_n831 ) , .A1( us10_n834 ) , .B1( us10_n863 ) );
  OAI221_X1 us10_U172 (.A( us10_n696 ) , .ZN( us10_n703 ) , .C2( us10_n784 ) , .C1( us10_n785 ) , .B1( us10_n786 ) , .B2( us10_n806 ) );
  AOI22_X1 us10_U173 (.ZN( us10_n696 ) , .A1( us10_n830 ) , .B2( us10_n843 ) , .A2( us10_n865 ) , .B1( us10_n868 ) );
  OAI221_X1 us10_U174 (.A( us10_n727 ) , .C2( us10_n728 ) , .B2( us10_n729 ) , .B1( us10_n730 ) , .ZN( us10_n737 ) , .C1( us10_n817 ) );
  AOI22_X1 us10_U175 (.ZN( us10_n727 ) , .B1( us10_n832 ) , .A2( us10_n838 ) , .A1( us10_n863 ) , .B2( us10_n866 ) );
  INV_X1 us10_U176 (.A( us10_n784 ) , .ZN( us10_n861 ) );
  OAI22_X1 us10_U177 (.ZN( us10_n710 ) , .A2( us10_n728 ) , .B2( us10_n729 ) , .A1( us10_n744 ) , .B1( us10_n813 ) );
  INV_X1 us10_U178 (.A( us10_n816 ) , .ZN( us10_n831 ) );
  INV_X1 us10_U179 (.A( us10_n788 ) , .ZN( us10_n845 ) );
  AOI222_X1 us10_U18 (.ZN( us10_n563 ) , .B1( us10_n830 ) , .C1( us10_n841 ) , .A2( us10_n843 ) , .A1( us10_n854 ) , .B2( us10_n863 ) , .C2( us10_n873 ) );
  OAI22_X1 us10_U180 (.ZN( us10_n588 ) , .A2( us10_n747 ) , .B2( us10_n762 ) , .A1( us10_n763 ) , .B1( us10_n784 ) );
  OAI22_X1 us10_U181 (.ZN( us10_n489 ) , .A1( us10_n724 ) , .B2( us10_n728 ) , .B1( us10_n730 ) , .A2( us10_n779 ) );
  OAI22_X1 us10_U182 (.ZN( us10_n624 ) , .B1( us10_n669 ) , .B2( us10_n747 ) , .A1( us10_n815 ) , .A2( us10_n816 ) );
  INV_X1 us10_U183 (.A( us10_n744 ) , .ZN( us10_n837 ) );
  OAI22_X1 us10_U184 (.ZN( us10_n681 ) , .A1( us10_n699 ) , .A2( us10_n730 ) , .B2( us10_n784 ) , .B1( us10_n817 ) );
  OAI22_X1 us10_U185 (.B2( us10_n779 ) , .B1( us10_n780 ) , .ZN( us10_n781 ) , .A2( us10_n814 ) , .A1( us10_n815 ) );
  OAI22_X1 us10_U186 (.A1( us10_n724 ) , .ZN( us10_n726 ) , .B2( us10_n750 ) , .B1( us10_n812 ) , .A2( us10_n816 ) );
  INV_X1 us10_U187 (.A( us10_n814 ) , .ZN( us10_n833 ) );
  OAI22_X1 us10_U188 (.B2( us10_n744 ) , .ZN( us10_n746 ) , .A2( us10_n762 ) , .B1( us10_n780 ) , .A1( us10_n792 ) );
  INV_X1 us10_U189 (.A( us10_n669 ) , .ZN( us10_n865 ) );
  NOR4_X1 us10_U19 (.ZN( us10_n473 ) , .A2( us10_n521 ) , .A4( us10_n594 ) , .A1( us10_n609 ) , .A3( us10_n629 ) );
  OAI22_X1 us10_U190 (.ZN( us10_n496 ) , .A2( us10_n744 ) , .A1( us10_n780 ) , .B1( us10_n791 ) , .B2( us10_n806 ) );
  INV_X1 us10_U191 (.A( us10_n750 ) , .ZN( us10_n842 ) );
  AOI211_X1 us10_U192 (.A( us10_n637 ) , .ZN( us10_n645 ) , .B( us10_n743 ) , .C2( us10_n839 ) , .C1( us10_n854 ) );
  OAI22_X1 us10_U193 (.ZN( us10_n637 ) , .A1( us10_n699 ) , .B2( us10_n728 ) , .A2( us10_n762 ) , .B1( us10_n816 ) );
  OAI22_X1 us10_U194 (.ZN( us10_n590 ) , .B1( us10_n730 ) , .B2( us10_n749 ) , .A2( us10_n786 ) , .A1( us10_n803 ) );
  OAI22_X1 us10_U195 (.ZN( us10_n695 ) , .A2( us10_n730 ) , .A1( us10_n780 ) , .B1( us10_n791 ) , .B2( us10_n817 ) );
  INV_X1 us10_U196 (.A( us10_n747 ) , .ZN( us10_n834 ) );
  NOR2_X1 us10_U197 (.A1( us10_n697 ) , .ZN( us10_n770 ) , .A2( us10_n815 ) );
  NOR2_X1 us10_U198 (.ZN( us10_n666 ) , .A1( us10_n728 ) , .A2( us10_n803 ) );
  NOR2_X1 us10_U199 (.ZN( us10_n594 ) , .A2( us10_n697 ) , .A1( us10_n728 ) );
  NOR4_X1 us10_U20 (.ZN( us10_n479 ) , .A1( us10_n520 ) , .A4( us10_n557 ) , .A3( us10_n582 ) , .A2( us10_n630 ) );
  NOR2_X1 us10_U200 (.ZN( us10_n600 ) , .A2( us10_n697 ) , .A1( us10_n784 ) );
  NOR2_X1 us10_U201 (.ZN( us10_n570 ) , .A1( us10_n728 ) , .A2( us10_n806 ) );
  NOR2_X1 us10_U202 (.ZN( us10_n532 ) , .A2( us10_n749 ) , .A1( us10_n750 ) );
  NOR2_X1 us10_U203 (.ZN( us10_n615 ) , .A1( us10_n785 ) , .A2( us10_n815 ) );
  NOR2_X1 us10_U204 (.ZN( us10_n629 ) , .A2( us10_n728 ) , .A1( us10_n785 ) );
  NOR2_X1 us10_U205 (.ZN( us10_n654 ) , .A1( us10_n728 ) , .A2( us10_n813 ) );
  NOR2_X1 us10_U206 (.ZN( us10_n546 ) , .A2( us10_n780 ) , .A1( us10_n814 ) );
  NOR2_X1 us10_U207 (.ZN( us10_n718 ) , .A2( us10_n724 ) , .A1( us10_n744 ) );
  NOR2_X1 us10_U208 (.ZN( us10_n577 ) , .A2( us10_n699 ) , .A1( us10_n814 ) );
  NOR2_X1 us10_U209 (.ZN( us10_n612 ) , .A1( us10_n779 ) , .A2( us10_n786 ) );
  NOR4_X1 us10_U21 (.A4( us10_n532 ) , .A3( us10_n533 ) , .A2( us10_n534 ) , .ZN( us10_n535 ) , .A1( us10_n820 ) );
  NOR2_X1 us10_U210 (.ZN( us10_n628 ) , .A2( us10_n669 ) , .A1( us10_n785 ) );
  NOR2_X1 us10_U211 (.ZN( us10_n610 ) , .A1( us10_n784 ) , .A2( us10_n816 ) );
  NOR2_X1 us10_U212 (.ZN( us10_n651 ) , .A1( us10_n784 ) , .A2( us10_n788 ) );
  NOR2_X1 us10_U213 (.ZN( us10_n531 ) , .A2( us10_n780 ) , .A1( us10_n816 ) );
  NOR2_X1 us10_U214 (.ZN( us10_n599 ) , .A2( us10_n791 ) , .A1( us10_n816 ) );
  INV_X1 us10_U215 (.A( us10_n728 ) , .ZN( us10_n852 ) );
  NOR2_X1 us10_U216 (.A2( us10_n708 ) , .A1( us10_n750 ) , .ZN( us10_n771 ) );
  NOR2_X1 us10_U217 (.A1( us10_n699 ) , .ZN( us10_n768 ) , .A2( us10_n813 ) );
  NOR2_X1 us10_U218 (.ZN( us10_n667 ) , .A1( us10_n750 ) , .A2( us10_n815 ) );
  NOR2_X1 us10_U219 (.ZN( us10_n541 ) , .A2( us10_n697 ) , .A1( us10_n699 ) );
  NOR4_X1 us10_U22 (.A4( us10_n541 ) , .A3( us10_n542 ) , .A2( us10_n543 ) , .ZN( us10_n550 ) , .A1( us10_n688 ) );
  NOR2_X1 us10_U220 (.ZN( us10_n508 ) , .A2( us10_n780 ) , .A1( us10_n785 ) );
  NOR2_X1 us10_U221 (.ZN( us10_n543 ) , .A2( us10_n708 ) , .A1( us10_n785 ) );
  NOR2_X1 us10_U222 (.ZN( us10_n555 ) , .A1( us10_n750 ) , .A2( us10_n791 ) );
  NOR2_X1 us10_U223 (.ZN( us10_n611 ) , .A2( us10_n780 ) , .A1( us10_n806 ) );
  NOR2_X1 us10_U224 (.ZN( us10_n664 ) , .A1( us10_n785 ) , .A2( us10_n791 ) );
  NOR2_X1 us10_U225 (.ZN( us10_n652 ) , .A1( us10_n669 ) , .A2( us10_n814 ) );
  NOR2_X1 us10_U226 (.A1( us10_n669 ) , .ZN( us10_n673 ) , .A2( us10_n744 ) );
  NOR2_X1 us10_U227 (.ZN( us10_n602 ) , .A1( us10_n669 ) , .A2( us10_n803 ) );
  NOR2_X1 us10_U228 (.A1( us10_n669 ) , .ZN( us10_n688 ) , .A2( us10_n816 ) );
  NOR2_X1 us10_U229 (.A2( us10_n744 ) , .ZN( us10_n769 ) , .A1( us10_n812 ) );
  AOI221_X1 us10_U23 (.A( us10_n713 ) , .B2( us10_n714 ) , .ZN( us10_n720 ) , .C1( us10_n832 ) , .B1( us10_n839 ) , .C2( us10_n863 ) );
  INV_X1 us10_U230 (.A( us10_n792 ) , .ZN( us10_n851 ) );
  NOR2_X1 us10_U231 (.A1( us10_n669 ) , .ZN( us10_n766 ) , .A2( us10_n813 ) );
  NOR2_X1 us10_U232 (.ZN( us10_n527 ) , .A1( us10_n669 ) , .A2( us10_n779 ) );
  NOR2_X1 us10_U233 (.A2( us10_n697 ) , .ZN( us10_n716 ) , .A1( us10_n792 ) );
  OAI22_X1 us10_U234 (.B1( us10_n440 ) , .ZN( us10_n444 ) , .A2( us10_n728 ) , .A1( us10_n744 ) , .B2( us10_n749 ) );
  NOR3_X1 us10_U235 (.ZN( us10_n440 ) , .A2( us10_n836 ) , .A3( us10_n837 ) , .A1( us10_n846 ) );
  NOR2_X1 us10_U236 (.ZN( us10_n601 ) , .A2( us10_n780 ) , .A1( us10_n803 ) );
  NOR2_X1 us10_U237 (.ZN( us10_n661 ) , .A1( us10_n729 ) , .A2( us10_n790 ) );
  NOR2_X1 us10_U238 (.ZN( us10_n631 ) , .A1( us10_n724 ) , .A2( us10_n813 ) );
  NOR2_X1 us10_U239 (.ZN( us10_n528 ) , .A2( us10_n724 ) , .A1( us10_n803 ) );
  OR2_X1 us10_U24 (.A2( us10_n711 ) , .A1( us10_n712 ) , .ZN( us10_n713 ) );
  NOR2_X1 us10_U240 (.ZN( us10_n509 ) , .A1( us10_n729 ) , .A2( us10_n779 ) );
  NOR2_X1 us10_U241 (.ZN( us10_n507 ) , .A1( us10_n812 ) , .A2( us10_n817 ) );
  NOR2_X1 us10_U242 (.ZN( us10_n662 ) , .A2( us10_n697 ) , .A1( us10_n729 ) );
  NOR2_X1 us10_U243 (.ZN( us10_n630 ) , .A1( us10_n747 ) , .A2( us10_n815 ) );
  NOR2_X1 us10_U244 (.ZN( us10_n554 ) , .A1( us10_n786 ) , .A2( us10_n813 ) );
  NOR2_X1 us10_U245 (.ZN( us10_n545 ) , .A1( us10_n749 ) , .A2( us10_n814 ) );
  NOR2_X1 us10_U246 (.ZN( us10_n557 ) , .A1( us10_n792 ) , .A2( us10_n814 ) );
  NOR2_X1 us10_U247 (.ZN( us10_n717 ) , .A2( us10_n744 ) , .A1( us10_n786 ) );
  NOR2_X1 us10_U248 (.ZN( us10_n544 ) , .A2( us10_n785 ) , .A1( us10_n792 ) );
  INV_X1 us10_U249 (.A( us10_n806 ) , .ZN( us10_n841 ) );
  NOR2_X1 us10_U25 (.ZN( us10_n680 ) , .A2( us10_n834 ) , .A1( us10_n839 ) );
  OAI21_X1 us10_U250 (.ZN( us10_n731 ) , .A( us10_n833 ) , .B2( us10_n852 ) , .B1( us10_n873 ) );
  NOR2_X1 us10_U251 (.A2( us10_n697 ) , .A1( us10_n780 ) , .ZN( us10_n820 ) );
  NOR2_X1 us10_U252 (.ZN( us10_n663 ) , .A1( us10_n729 ) , .A2( us10_n785 ) );
  OAI22_X1 us10_U253 (.B2( us10_n750 ) , .B1( us10_n751 ) , .A1( us10_n752 ) , .ZN( us10_n756 ) , .A2( us10_n806 ) );
  NOR2_X1 us10_U254 (.ZN( us10_n751 ) , .A2( us10_n852 ) , .A1( us10_n860 ) );
  NOR3_X1 us10_U255 (.ZN( us10_n752 ) , .A2( us10_n853 ) , .A1( us10_n863 ) , .A3( us10_n865 ) );
  NOR2_X1 us10_U256 (.ZN( us10_n656 ) , .A1( us10_n747 ) , .A2( us10_n780 ) );
  NOR2_X1 us10_U257 (.ZN( us10_n530 ) , .A2( us10_n744 ) , .A1( us10_n792 ) );
  NOR2_X1 us10_U258 (.ZN( us10_n506 ) , .A2( us10_n728 ) , .A1( us10_n762 ) );
  NOR2_X1 us10_U259 (.ZN( us10_n558 ) , .A1( us10_n708 ) , .A2( us10_n816 ) );
  NOR4_X1 us10_U26 (.A4( us10_n514 ) , .A3( us10_n515 ) , .A2( us10_n516 ) , .A1( us10_n517 ) , .ZN( us10_n524 ) );
  NOR2_X1 us10_U260 (.ZN( us10_n516 ) , .A1( us10_n708 ) , .A2( us10_n744 ) );
  NOR2_X1 us10_U261 (.ZN( us10_n614 ) , .A1( us10_n762 ) , .A2( us10_n812 ) );
  AOI21_X1 us10_U262 (.A( us10_n812 ) , .B2( us10_n813 ) , .B1( us10_n814 ) , .ZN( us10_n819 ) );
  NOR2_X1 us10_U263 (.A1( us10_n749 ) , .ZN( us10_n767 ) , .A2( us10_n803 ) );
  AOI21_X1 us10_U264 (.ZN( us10_n593 ) , .B1( us10_n750 ) , .A( us10_n792 ) , .B2( us10_n813 ) );
  NOR2_X1 us10_U265 (.A1( us10_n730 ) , .ZN( us10_n765 ) , .A2( us10_n786 ) );
  NOR2_X1 us10_U266 (.ZN( us10_n655 ) , .A1( us10_n790 ) , .A2( us10_n815 ) );
  NOR2_X1 us10_U267 (.ZN( us10_n701 ) , .A2( us10_n786 ) , .A1( us10_n817 ) );
  NOR2_X1 us10_U268 (.ZN( us10_n579 ) , .A2( us10_n708 ) , .A1( us10_n730 ) );
  NOR2_X1 us10_U269 (.ZN( us10_n533 ) , .A2( us10_n724 ) , .A1( us10_n730 ) );
  AOI222_X1 us10_U27 (.ZN( us10_n525 ) , .A1( us10_n834 ) , .B2( us10_n837 ) , .C1( us10_n844 ) , .C2( us10_n850 ) , .A2( us10_n852 ) , .B1( us10_n866 ) );
  NOR2_X1 us10_U270 (.ZN( us10_n668 ) , .A2( us10_n708 ) , .A1( us10_n790 ) );
  INV_X1 us10_U271 (.A( us10_n813 ) , .ZN( us10_n836 ) );
  NOR2_X1 us10_U272 (.ZN( us10_n521 ) , .A1( us10_n790 ) , .A2( us10_n812 ) );
  AOI21_X1 us10_U273 (.ZN( us10_n571 ) , .B2( us10_n697 ) , .B1( us10_n806 ) , .A( us10_n812 ) );
  INV_X1 us10_U274 (.A( us10_n763 ) , .ZN( us10_n866 ) );
  NOR2_X1 us10_U275 (.ZN( us10_n517 ) , .A1( us10_n708 ) , .A2( us10_n803 ) );
  AOI21_X1 us10_U276 (.A( us10_n815 ) , .B2( us10_n816 ) , .B1( us10_n817 ) , .ZN( us10_n818 ) );
  INV_X1 us10_U277 (.A( us10_n729 ) , .ZN( us10_n868 ) );
  NOR2_X1 us10_U278 (.ZN( us10_n542 ) , .A1( us10_n762 ) , .A2( us10_n791 ) );
  AOI21_X1 us10_U279 (.ZN( us10_n499 ) , .B1( us10_n680 ) , .A( us10_n812 ) , .B2( us10_n816 ) );
  NOR4_X1 us10_U28 (.A3( us10_n521 ) , .A1( us10_n522 ) , .ZN( us10_n523 ) , .A2( us10_n673 ) , .A4( us10_n769 ) );
  NOR2_X1 us10_U280 (.ZN( us10_n609 ) , .A2( us10_n724 ) , .A1( us10_n817 ) );
  NOR2_X1 us10_U281 (.ZN( us10_n642 ) , .A2( us10_n788 ) , .A1( us10_n791 ) );
  AOI21_X1 us10_U282 (.ZN( us10_n592 ) , .B1( us10_n728 ) , .B2( us10_n784 ) , .A( us10_n790 ) );
  NOR2_X1 us10_U283 (.ZN( us10_n653 ) , .A1( us10_n762 ) , .A2( us10_n786 ) );
  AOI21_X1 us10_U284 (.B1( us10_n625 ) , .ZN( us10_n627 ) , .A( us10_n763 ) , .B2( us10_n814 ) );
  AOI21_X1 us10_U285 (.ZN( us10_n478 ) , .B2( us10_n697 ) , .A( us10_n749 ) , .B1( us10_n779 ) );
  AOI21_X1 us10_U286 (.ZN( us10_n648 ) , .A( us10_n762 ) , .B2( us10_n784 ) , .B1( us10_n792 ) );
  AOI21_X1 us10_U287 (.ZN( us10_n623 ) , .B1( us10_n699 ) , .A( us10_n779 ) , .B2( us10_n784 ) );
  NOR2_X1 us10_U288 (.ZN( us10_n582 ) , .A1( us10_n744 ) , .A2( us10_n815 ) );
  NOR2_X1 us10_U289 (.A2( us10_n708 ) , .A1( us10_n762 ) , .ZN( us10_n794 ) );
  AOI221_X1 us10_U29 (.A( us10_n781 ) , .ZN( us10_n798 ) , .C2( us10_n837 ) , .B2( us10_n838 ) , .B1( us10_n865 ) , .C1( us10_n866 ) );
  NOR2_X1 us10_U290 (.ZN( us10_n553 ) , .A2( us10_n744 ) , .A1( us10_n784 ) );
  NOR2_X1 us10_U291 (.ZN( us10_n519 ) , .A2( us10_n699 ) , .A1( us10_n816 ) );
  AOI21_X1 us10_U292 (.ZN( us10_n626 ) , .B2( us10_n669 ) , .A( us10_n790 ) , .B1( us10_n791 ) );
  NOR2_X1 us10_U293 (.ZN( us10_n520 ) , .A2( us10_n708 ) , .A1( us10_n814 ) );
  AOI21_X1 us10_U294 (.ZN( us10_n477 ) , .A( us10_n669 ) , .B1( us10_n750 ) , .B2( us10_n806 ) );
  AOI21_X1 us10_U295 (.ZN( us10_n589 ) , .B2( us10_n699 ) , .B1( us10_n815 ) , .A( us10_n817 ) );
  AOI21_X1 us10_U296 (.ZN( us10_n510 ) , .B2( us10_n669 ) , .A( us10_n730 ) , .B1( us10_n815 ) );
  AOI21_X1 us10_U297 (.ZN( us10_n540 ) , .A( us10_n763 ) , .B2( us10_n779 ) , .B1( us10_n817 ) );
  AOI21_X1 us10_U298 (.ZN( us10_n515 ) , .A( us10_n729 ) , .B1( us10_n750 ) , .B2( us10_n803 ) );
  NOR2_X1 us10_U299 (.ZN( us10_n547 ) , .A1( us10_n699 ) , .A2( us10_n744 ) );
  NAND4_X1 us10_U3 (.ZN( sa13_sr_0 ) , .A4( us10_n501 ) , .A3( us10_n502 ) , .A2( us10_n503 ) , .A1( us10_n504 ) );
  NOR4_X1 us10_U30 (.A4( us10_n793 ) , .A3( us10_n794 ) , .A2( us10_n795 ) , .A1( us10_n796 ) , .ZN( us10_n797 ) );
  NOR2_X1 us10_U300 (.ZN( us10_n581 ) , .A1( us10_n669 ) , .A2( us10_n788 ) );
  AOI21_X1 us10_U301 (.ZN( us10_n539 ) , .B2( us10_n812 ) , .A( us10_n814 ) , .B1( us10_n815 ) );
  NOR2_X1 us10_U302 (.ZN( us10_n559 ) , .A2( us10_n791 ) , .A1( us10_n803 ) );
  AOI21_X1 us10_U303 (.ZN( us10_n498 ) , .A( us10_n724 ) , .B2( us10_n762 ) , .B1( us10_n814 ) );
  NAND2_X2 us10_U304 (.A2( us10_n461 ) , .A1( us10_n462 ) , .ZN( us10_n747 ) );
  AOI21_X1 us10_U305 (.B1( us10_n699 ) , .ZN( us10_n700 ) , .A( us10_n732 ) , .B2( us10_n763 ) );
  AOI21_X1 us10_U306 (.ZN( us10_n591 ) , .B2( us10_n763 ) , .A( us10_n785 ) , .B1( us10_n812 ) );
  AOI21_X1 us10_U307 (.ZN( us10_n640 ) , .B2( us10_n747 ) , .A( us10_n792 ) , .B1( us10_n803 ) );
  AOI21_X1 us10_U308 (.ZN( us10_n569 ) , .B1( us10_n750 ) , .B2( us10_n762 ) , .A( us10_n780 ) );
  NOR2_X1 us10_U309 (.ZN( us10_n683 ) , .A2( us10_n699 ) , .A1( us10_n803 ) );
  NOR4_X1 us10_U31 (.A4( us10_n776 ) , .A3( us10_n777 ) , .A1( us10_n778 ) , .ZN( us10_n799 ) , .A2( us10_n801 ) );
  NOR2_X1 us10_U310 (.ZN( us10_n665 ) , .A1( us10_n780 ) , .A2( us10_n813 ) );
  AOI21_X1 us10_U311 (.ZN( us10_n500 ) , .A( us10_n697 ) , .B1( us10_n708 ) , .B2( us10_n786 ) );
  NOR2_X1 us10_U312 (.ZN( us10_n685 ) , .A1( us10_n729 ) , .A2( us10_n816 ) );
  INV_X1 us10_U313 (.A( us10_n791 ) , .ZN( us10_n873 ) );
  AOI21_X1 us10_U314 (.ZN( us10_n649 ) , .B1( us10_n729 ) , .B2( us10_n763 ) , .A( us10_n813 ) );
  AOI21_X1 us10_U315 (.B1( us10_n686 ) , .ZN( us10_n687 ) , .A( us10_n728 ) , .B2( us10_n761 ) );
  INV_X1 us10_U316 (.A( us10_n699 ) , .ZN( us10_n853 ) );
  NOR2_X1 us10_U317 (.ZN( us10_n568 ) , .A1( us10_n729 ) , .A2( us10_n762 ) );
  NOR2_X1 us10_U318 (.ZN( us10_n578 ) , .A1( us10_n708 ) , .A2( us10_n813 ) );
  AOI21_X1 us10_U319 (.ZN( us10_n514 ) , .A( us10_n779 ) , .B2( us10_n792 ) , .B1( us10_n812 ) );
  NOR4_X1 us10_U32 (.A4( us10_n734 ) , .A3( us10_n735 ) , .A2( us10_n736 ) , .A1( us10_n737 ) , .ZN( us10_n738 ) );
  NOR2_X1 us10_U320 (.ZN( us10_n684 ) , .A1( us10_n791 ) , .A2( us10_n813 ) );
  NOR2_X1 us10_U321 (.ZN( us10_n580 ) , .A2( us10_n697 ) , .A1( us10_n791 ) );
  NOR2_X1 us10_U322 (.A2( us10_n813 ) , .A1( us10_n815 ) , .ZN( us10_n821 ) );
  NOR2_X1 us10_U323 (.ZN( us10_n566 ) , .A2( us10_n697 ) , .A1( us10_n763 ) );
  AOI21_X1 us10_U324 (.ZN( us10_n497 ) , .A( us10_n779 ) , .B2( us10_n791 ) , .B1( us10_n804 ) );
  AOI21_X1 us10_U325 (.ZN( us10_n564 ) , .B1( us10_n724 ) , .A( us10_n779 ) , .B2( us10_n791 ) );
  NOR2_X1 us10_U326 (.ZN( us10_n632 ) , .A2( us10_n697 ) , .A1( us10_n724 ) );
  NAND2_X2 us10_U327 (.A2( us10_n454 ) , .A1( us10_n472 ) , .ZN( us10_n779 ) );
  NOR2_X1 us10_U328 (.ZN( us10_n529 ) , .A1( us10_n708 ) , .A2( us10_n779 ) );
  AOI21_X1 us10_U329 (.ZN( us10_n639 ) , .B2( us10_n749 ) , .A( us10_n788 ) , .B1( us10_n812 ) );
  AOI211_X1 us10_U33 (.B( us10_n725 ) , .A( us10_n726 ) , .ZN( us10_n739 ) , .C1( us10_n843 ) , .C2( us10_n855 ) );
  AOI21_X1 us10_U330 (.ZN( us10_n689 ) , .B2( us10_n749 ) , .B1( us10_n763 ) , .A( us10_n806 ) );
  AOI21_X1 us10_U331 (.A( us10_n790 ) , .B2( us10_n791 ) , .B1( us10_n792 ) , .ZN( us10_n793 ) );
  AOI21_X1 us10_U332 (.A( us10_n733 ) , .ZN( us10_n734 ) , .B2( us10_n780 ) , .B1( us10_n792 ) );
  AOI21_X1 us10_U333 (.ZN( us10_n641 ) , .B1( us10_n680 ) , .A( us10_n791 ) , .B2( us10_n817 ) );
  NOR2_X1 us10_U334 (.ZN( us10_n583 ) , .A1( us10_n792 ) , .A2( us10_n817 ) );
  NOR2_X1 us10_U335 (.ZN( us10_n711 ) , .A1( us10_n762 ) , .A2( us10_n763 ) );
  NOR2_X1 us10_U336 (.ZN( us10_n534 ) , .A1( us10_n724 ) , .A2( us10_n788 ) );
  NOR2_X1 us10_U337 (.ZN( us10_n682 ) , .A2( us10_n708 ) , .A1( us10_n817 ) );
  INV_X1 us10_U338 (.A( us10_n697 ) , .ZN( us10_n838 ) );
  AOI21_X1 us10_U339 (.ZN( us10_n442 ) , .A( us10_n699 ) , .B1( us10_n733 ) , .B2( us10_n750 ) );
  NOR3_X1 us10_U34 (.A3( us10_n722 ) , .A1( us10_n723 ) , .ZN( us10_n740 ) , .A2( us10_n741 ) );
  NAND2_X2 us10_U340 (.A1( us10_n455 ) , .A2( us10_n462 ) , .ZN( us10_n750 ) );
  INV_X1 us10_U341 (.A( us10_n815 ) , .ZN( us10_n855 ) );
  OAI21_X1 us10_U342 (.A( us10_n613 ) , .ZN( us10_n616 ) , .B1( us10_n625 ) , .B2( us10_n784 ) );
  NAND2_X2 us10_U343 (.A1( us10_n462 ) , .A2( us10_n472 ) , .ZN( us10_n788 ) );
  OAI21_X1 us10_U344 (.A( us10_n698 ) , .ZN( us10_n702 ) , .B2( us10_n750 ) , .B1( us10_n804 ) );
  OAI21_X1 us10_U345 (.ZN( us10_n698 ) , .B2( us10_n833 ) , .B1( us10_n838 ) , .A( us10_n860 ) );
  INV_X1 us10_U346 (.A( us10_n785 ) , .ZN( us10_n846 ) );
  INV_X1 us10_U347 (.A( us10_n780 ) , .ZN( us10_n850 ) );
  OAI21_X1 us10_U348 (.A( us10_n787 ) , .B2( us10_n788 ) , .B1( us10_n789 ) , .ZN( us10_n795 ) );
  OAI21_X1 us10_U349 (.ZN( us10_n787 ) , .A( us10_n839 ) , .B1( us10_n863 ) , .B2( us10_n873 ) );
  NOR4_X1 us10_U35 (.A3( us10_n755 ) , .A2( us10_n756 ) , .A1( us10_n757 ) , .ZN( us10_n758 ) , .A4( us10_n869 ) );
  NAND2_X1 us10_U350 (.A1( us10_n729 ) , .A2( us10_n784 ) , .ZN( us10_n811 ) );
  NAND2_X1 us10_U351 (.ZN( us10_n671 ) , .A1( us10_n806 ) , .A2( us10_n816 ) );
  NAND2_X1 us10_U352 (.ZN( us10_n714 ) , .A1( us10_n728 ) , .A2( us10_n780 ) );
  AOI21_X1 us10_U353 (.ZN( us10_n443 ) , .B1( us10_n789 ) , .B2( us10_n791 ) , .A( us10_n814 ) );
  NOR2_X1 us10_U354 (.ZN( us10_n712 ) , .A2( us10_n724 ) , .A1( us10_n790 ) );
  NAND2_X1 us10_U355 (.A2( us10_n762 ) , .A1( us10_n806 ) , .ZN( us10_n810 ) );
  NAND2_X2 us10_U356 (.A1( us10_n454 ) , .A2( us10_n461 ) , .ZN( us10_n813 ) );
  NOR2_X1 us10_U357 (.ZN( us10_n470 ) , .A2( us10_n779 ) , .A1( us10_n815 ) );
  NAND2_X1 us10_U358 (.A1( us10_n699 ) , .A2( us10_n729 ) , .ZN( us10_n782 ) );
  NOR2_X1 us10_U359 (.ZN( us10_n526 ) , .A1( us10_n724 ) , .A2( us10_n750 ) );
  AOI211_X1 us10_U36 (.B( us10_n745 ) , .A( us10_n746 ) , .ZN( us10_n759 ) , .C1( us10_n832 ) , .C2( us10_n853 ) );
  NOR2_X1 us10_U360 (.ZN( us10_n518 ) , .A1( us10_n708 ) , .A2( us10_n788 ) );
  NAND2_X1 us10_U361 (.A2( us10_n749 ) , .A1( us10_n786 ) , .ZN( us10_n809 ) );
  INV_X1 us10_U362 (.A( us10_n817 ) , .ZN( us10_n844 ) );
  NAND2_X2 us10_U363 (.A1( us10_n451 ) , .A2( us10_n454 ) , .ZN( us10_n814 ) );
  INV_X1 us10_U364 (.A( us10_n724 ) , .ZN( us10_n856 ) );
  AND2_X1 us10_U365 (.ZN( us10_n732 ) , .A1( us10_n779 ) , .A2( us10_n785 ) );
  AOI221_X1 us10_U366 (.A( us10_n764 ) , .ZN( us10_n774 ) , .C2( us10_n810 ) , .B2( us10_n835 ) , .C1( us10_n855 ) , .B1( us10_n866 ) );
  AOI21_X1 us10_U367 (.B2( us10_n763 ) , .ZN( us10_n764 ) , .A( us10_n788 ) , .B1( us10_n792 ) );
  INV_X1 us10_U368 (.A( us10_n761 ) , .ZN( us10_n835 ) );
  NAND2_X1 us10_U369 (.A1( us10_n451 ) , .A2( us10_n471 ) , .ZN( us10_n816 ) );
  NOR3_X1 us10_U37 (.A3( us10_n741 ) , .A2( us10_n742 ) , .A1( us10_n743 ) , .ZN( us10_n760 ) );
  NAND2_X1 us10_U370 (.A2( us10_n441 ) , .A1( us10_n447 ) , .ZN( us10_n784 ) );
  NAND2_X1 us10_U371 (.A2( us10_n448 ) , .A1( us10_n460 ) , .ZN( us10_n728 ) );
  NAND2_X1 us10_U372 (.A1( us10_n453 ) , .A2( us10_n472 ) , .ZN( us10_n785 ) );
  NAND2_X1 us10_U373 (.A1( us10_n453 ) , .A2( us10_n461 ) , .ZN( us10_n744 ) );
  NAND2_X1 us10_U374 (.A1( us10_n452 ) , .A2( us10_n465 ) , .ZN( us10_n669 ) );
  NAND2_X1 us10_U375 (.A2( us10_n453 ) , .A1( us10_n455 ) , .ZN( us10_n806 ) );
  NAND2_X1 us10_U376 (.A1( us10_n441 ) , .A2( us10_n460 ) , .ZN( us10_n699 ) );
  NAND2_X1 us10_U377 (.A1( us10_n455 ) , .A2( us10_n471 ) , .ZN( us10_n803 ) );
  NAND2_X1 us10_U378 (.A2( us10_n464 ) , .A1( us10_n465 ) , .ZN( us10_n812 ) );
  NAND2_X1 us10_U379 (.A1( us10_n447 ) , .A2( us10_n448 ) , .ZN( us10_n786 ) );
  NAND4_X1 us10_U38 (.ZN( sa13_sr_3 ) , .A4( us10_n704 ) , .A3( us10_n705 ) , .A2( us10_n706 ) , .A1( us10_n707 ) );
  NAND2_X2 us10_U380 (.A2( us10_n461 ) , .A1( us10_n471 ) , .ZN( us10_n697 ) );
  NAND2_X1 us10_U381 (.A2( us10_n448 ) , .A1( us10_n452 ) , .ZN( us10_n729 ) );
  NAND2_X1 us10_U382 (.A2( us10_n449 ) , .A1( us10_n452 ) , .ZN( us10_n763 ) );
  NAND2_X1 us10_U383 (.A2( us10_n454 ) , .A1( us10_n455 ) , .ZN( us10_n730 ) );
  NOR2_X1 us10_U384 (.ZN( us10_n465 ) , .A2( us10_n847 ) , .A1( us10_n848 ) );
  NOR2_X1 us10_U385 (.ZN( us10_n453 ) , .A1( us10_n826 ) , .A2( us10_n827 ) );
  NOR2_X1 us10_U386 (.ZN( us10_n451 ) , .A1( us10_n828 ) , .A2( us10_n829 ) );
  NAND2_X1 us10_U387 (.A1( us10_n451 ) , .A2( us10_n462 ) , .ZN( us10_n790 ) );
  NAND2_X2 us10_U388 (.A2( us10_n448 ) , .A1( us10_n464 ) , .ZN( us10_n815 ) );
  NAND2_X2 us10_U389 (.A2( us10_n441 ) , .A1( us10_n452 ) , .ZN( us10_n791 ) );
  NOR4_X1 us10_U39 (.A4( us10_n700 ) , .A3( us10_n701 ) , .A2( us10_n702 ) , .A1( us10_n703 ) , .ZN( us10_n704 ) );
  NAND2_X2 us10_U390 (.A1( us10_n449 ) , .A2( us10_n464 ) , .ZN( us10_n724 ) );
  NAND2_X1 us10_U391 (.A1( us10_n447 ) , .A2( us10_n449 ) , .ZN( us10_n805 ) );
  NAND2_X2 us10_U392 (.A1( us10_n449 ) , .A2( us10_n460 ) , .ZN( us10_n792 ) );
  NAND2_X2 us10_U393 (.A1( us10_n441 ) , .A2( us10_n464 ) , .ZN( us10_n708 ) );
  NAND2_X2 us10_U394 (.A2( us10_n471 ) , .A1( us10_n472 ) , .ZN( us10_n817 ) );
  NAND2_X2 us10_U395 (.A2( us10_n460 ) , .A1( us10_n465 ) , .ZN( us10_n780 ) );
  NOR2_X1 us10_U396 (.ZN( us10_n447 ) , .A2( us10_n849 ) , .A1( us10_n858 ) );
  NOR2_X1 us10_U397 (.A2( sa10_6 ) , .A1( sa10_7 ) , .ZN( us10_n464 ) );
  NOR2_X1 us10_U398 (.A2( sa10_7 ) , .ZN( us10_n460 ) , .A1( us10_n849 ) );
  NOR2_X1 us10_U399 (.A2( sa10_4 ) , .ZN( us10_n449 ) , .A1( us10_n848 ) );
  NOR3_X1 us10_U4 (.ZN( us10_n598 ) , .A1( us10_n608 ) , .A3( us10_n723 ) , .A2( us10_n742 ) );
  AOI211_X1 us10_U40 (.B( us10_n694 ) , .A( us10_n695 ) , .ZN( us10_n705 ) , .C2( us10_n831 ) , .C1( us10_n851 ) );
  NOR2_X1 us10_U400 (.A2( sa10_4 ) , .A1( sa10_5 ) , .ZN( us10_n441 ) );
  NOR2_X1 us10_U401 (.A2( sa10_5 ) , .ZN( us10_n448 ) , .A1( us10_n847 ) );
  NOR2_X1 us10_U402 (.A2( sa10_1 ) , .ZN( us10_n471 ) , .A1( us10_n826 ) );
  NOR2_X1 us10_U403 (.A2( sa10_2 ) , .A1( sa10_3 ) , .ZN( us10_n472 ) );
  NOR2_X1 us10_U404 (.A2( sa10_6 ) , .ZN( us10_n452 ) , .A1( us10_n858 ) );
  NOR2_X1 us10_U405 (.A2( sa10_2 ) , .ZN( us10_n461 ) , .A1( us10_n829 ) );
  NOR2_X1 us10_U406 (.A2( sa10_3 ) , .ZN( us10_n455 ) , .A1( us10_n828 ) );
  INV_X1 us10_U407 (.A( sa10_6 ) , .ZN( us10_n849 ) );
  INV_X1 us10_U408 (.A( sa10_4 ) , .ZN( us10_n847 ) );
  INV_X1 us10_U409 (.A( sa10_3 ) , .ZN( us10_n829 ) );
  NOR2_X1 us10_U41 (.ZN( us10_n707 ) , .A2( us10_n776 ) , .A1( us10_n800 ) );
  INV_X1 us10_U410 (.A( sa10_2 ) , .ZN( us10_n828 ) );
  INV_X1 us10_U411 (.A( sa10_7 ) , .ZN( us10_n858 ) );
  INV_X1 us10_U412 (.A( sa10_5 ) , .ZN( us10_n848 ) );
  INV_X1 us10_U413 (.A( sa10_1 ) , .ZN( us10_n827 ) );
  INV_X1 us10_U414 (.A( sa10_0 ) , .ZN( us10_n826 ) );
  NOR2_X1 us10_U415 (.A2( sa10_0 ) , .A1( sa10_1 ) , .ZN( us10_n462 ) );
  NOR2_X1 us10_U416 (.A2( sa10_0 ) , .ZN( us10_n454 ) , .A1( us10_n827 ) );
  OAI222_X1 us10_U417 (.B2( us10_n747 ) , .B1( us10_n748 ) , .A2( us10_n749 ) , .ZN( us10_n757 ) , .C2( us10_n805 ) , .C1( us10_n814 ) , .A1( us10_n817 ) );
  OAI22_X1 us10_U418 (.B2( us10_n803 ) , .B1( us10_n804 ) , .A2( us10_n805 ) , .A1( us10_n806 ) , .ZN( us10_n808 ) );
  OAI21_X1 us10_U419 (.A( us10_n731 ) , .B1( us10_n732 ) , .ZN( us10_n736 ) , .B2( us10_n805 ) );
  NAND4_X1 us10_U42 (.ZN( sa13_sr_7 ) , .A4( us10_n822 ) , .A3( us10_n823 ) , .A2( us10_n824 ) , .A1( us10_n825 ) );
  OAI222_X1 us10_U420 (.ZN( us10_n505 ) , .C2( us10_n625 ) , .B2( us10_n647 ) , .B1( us10_n747 ) , .A2( us10_n748 ) , .C1( us10_n805 ) , .A1( us10_n806 ) );
  AOI21_X1 us10_U421 (.ZN( us10_n650 ) , .A( us10_n779 ) , .B1( us10_n792 ) , .B2( us10_n805 ) );
  INV_X1 us10_U422 (.A( us10_n805 ) , .ZN( us10_n860 ) );
  NOR2_X1 us10_U423 (.ZN( us10_n735 ) , .A2( us10_n803 ) , .A1( us10_n805 ) );
  NOR2_X1 us10_U424 (.ZN( us10_n484 ) , .A1( us10_n788 ) , .A2( us10_n805 ) );
  NOR2_X1 us10_U425 (.A2( us10_n744 ) , .ZN( us10_n755 ) , .A1( us10_n805 ) );
  NAND2_X1 us10_U426 (.ZN( us10_n753 ) , .A1( us10_n763 ) , .A2( us10_n805 ) );
  NOR2_X1 us10_U427 (.ZN( us10_n715 ) , .A1( us10_n805 ) , .A2( us10_n817 ) );
  NOR2_X1 us10_U428 (.ZN( us10_n567 ) , .A1( us10_n747 ) , .A2( us10_n805 ) );
  AOI21_X1 us10_U429 (.ZN( us10_n552 ) , .B1( us10_n669 ) , .A( us10_n697 ) , .B2( us10_n805 ) );
  NOR4_X1 us10_U43 (.A4( us10_n818 ) , .A3( us10_n819 ) , .A2( us10_n820 ) , .A1( us10_n821 ) , .ZN( us10_n822 ) );
  NOR2_X1 us10_U430 (.ZN( us10_n556 ) , .A1( us10_n762 ) , .A2( us10_n805 ) );
  NOR2_X1 us10_U431 (.ZN( us10_n670 ) , .A1( us10_n790 ) , .A2( us10_n805 ) );
  AND2_X1 us10_U432 (.ZN( us10_n438 ) , .A2( us10_n831 ) , .A1( us10_n854 ) );
  AND2_X1 us10_U433 (.ZN( us10_n439 ) , .A2( us10_n843 ) , .A1( us10_n861 ) );
  NOR3_X1 us10_U434 (.A1( us10_n438 ) , .A2( us10_n439 ) , .A3( us10_n576 ) , .ZN( us10_n587 ) );
  NAND4_X1 us10_U435 (.ZN( sa13_sr_2 ) , .A4( us10_n643 ) , .A3( us10_n644 ) , .A2( us10_n645 ) , .A1( us10_n646 ) );
  INV_X1 us10_U436 (.A( us10_n812 ) , .ZN( us10_n854 ) );
  NAND3_X1 us10_U437 (.ZN( sa13_sr_6 ) , .A3( us10_n797 ) , .A2( us10_n798 ) , .A1( us10_n799 ) );
  NAND3_X1 us10_U438 (.ZN( sa13_sr_5 ) , .A3( us10_n758 ) , .A2( us10_n759 ) , .A1( us10_n760 ) );
  NAND3_X1 us10_U439 (.ZN( sa13_sr_4 ) , .A3( us10_n738 ) , .A2( us10_n739 ) , .A1( us10_n740 ) );
  AOI222_X1 us10_U44 (.C2( us10_n809 ) , .B2( us10_n810 ) , .A2( us10_n811 ) , .ZN( us10_n823 ) , .C1( us10_n832 ) , .A1( us10_n839 ) , .B1( us10_n853 ) );
  NAND3_X1 us10_U440 (.A3( us10_n675 ) , .A2( us10_n676 ) , .A1( us10_n677 ) , .ZN( us10_n807 ) );
  NAND3_X1 us10_U441 (.ZN( us10_n638 ) , .A3( us10_n708 ) , .A2( us10_n724 ) , .A1( us10_n792 ) );
  NAND3_X1 us10_U442 (.A3( us10_n618 ) , .A2( us10_n619 ) , .A1( us10_n620 ) , .ZN( us10_n725 ) );
  NAND3_X1 us10_U443 (.A3( us10_n585 ) , .A2( us10_n586 ) , .A1( us10_n587 ) , .ZN( us10_n621 ) );
  NAND3_X1 us10_U444 (.ZN( us10_n565 ) , .A3( us10_n680 ) , .A2( us10_n750 ) , .A1( us10_n785 ) );
  NAND3_X1 us10_U445 (.A3( us10_n523 ) , .A2( us10_n524 ) , .A1( us10_n525 ) , .ZN( us10_n742 ) );
  NAND3_X1 us10_U446 (.A3( us10_n512 ) , .A1( us10_n513 ) , .ZN( us10_n608 ) , .A2( us10_n871 ) );
  NAND3_X1 us10_U447 (.A3( us10_n467 ) , .A2( us10_n468 ) , .A1( us10_n469 ) , .ZN( us10_n777 ) );
  INV_X1 us10_U448 (.A( us10_n803 ) , .ZN( us10_n843 ) );
  AOI21_X1 us10_U449 (.ZN( us10_n576 ) , .B2( us10_n724 ) , .B1( us10_n748 ) , .A( us10_n785 ) );
  AOI211_X1 us10_U45 (.B( us10_n807 ) , .A( us10_n808 ) , .ZN( us10_n824 ) , .C1( us10_n842 ) , .C2( us10_n850 ) );
  NOR4_X1 us10_U46 (.A4( us10_n498 ) , .A3( us10_n499 ) , .A2( us10_n500 ) , .ZN( us10_n501 ) , .A1( us10_n527 ) );
  AOI221_X1 us10_U47 (.A( us10_n497 ) , .ZN( us10_n502 ) , .B2( us10_n843 ) , .C1( us10_n846 ) , .C2( us10_n860 ) , .B1( us10_n862 ) );
  AOI211_X1 us10_U48 (.A( us10_n496 ) , .ZN( us10_n503 ) , .B( us10_n802 ) , .C2( us10_n839 ) , .C1( us10_n851 ) );
  NAND4_X1 us10_U49 (.ZN( sa13_sr_1 ) , .A4( us10_n595 ) , .A3( us10_n596 ) , .A2( us10_n597 ) , .A1( us10_n598 ) );
  NOR3_X1 us10_U5 (.A3( us10_n800 ) , .A2( us10_n801 ) , .A1( us10_n802 ) , .ZN( us10_n825 ) );
  NOR4_X1 us10_U50 (.A4( us10_n591 ) , .A3( us10_n592 ) , .A2( us10_n593 ) , .A1( us10_n594 ) , .ZN( us10_n595 ) );
  AOI211_X1 us10_U51 (.B( us10_n589 ) , .A( us10_n590 ) , .ZN( us10_n596 ) , .C2( us10_n811 ) , .C1( us10_n833 ) );
  AOI211_X1 us10_U52 (.A( us10_n588 ) , .ZN( us10_n597 ) , .B( us10_n621 ) , .C1( us10_n845 ) , .C2( us10_n855 ) );
  NOR2_X1 us10_U53 (.ZN( us10_n804 ) , .A1( us10_n854 ) , .A2( us10_n861 ) );
  NOR2_X1 us10_U54 (.ZN( us10_n625 ) , .A2( us10_n836 ) , .A1( us10_n839 ) );
  AOI222_X1 us10_U55 (.ZN( us10_n469 ) , .B1( us10_n832 ) , .A1( us10_n839 ) , .C1( us10_n842 ) , .C2( us10_n851 ) , .A2( us10_n855 ) , .B2( us10_n865 ) );
  NOR4_X1 us10_U56 (.A1( us10_n466 ) , .ZN( us10_n467 ) , .A4( us10_n542 ) , .A2( us10_n554 ) , .A3( us10_n614 ) );
  AOI221_X1 us10_U57 (.ZN( us10_n468 ) , .C2( us10_n714 ) , .B2( us10_n831 ) , .C1( us10_n845 ) , .B1( us10_n860 ) , .A( us10_n864 ) );
  NAND4_X1 us10_U58 (.A4( us10_n603 ) , .A3( us10_n604 ) , .A2( us10_n605 ) , .A1( us10_n606 ) , .ZN( us10_n722 ) );
  NOR3_X1 us10_U59 (.A1( us10_n599 ) , .ZN( us10_n604 ) , .A3( us10_n663 ) , .A2( us10_n770 ) );
  NOR3_X1 us10_U6 (.ZN( us10_n504 ) , .A2( us10_n679 ) , .A3( us10_n777 ) , .A1( us10_n876 ) );
  NOR4_X1 us10_U60 (.A3( us10_n600 ) , .A2( us10_n601 ) , .A1( us10_n602 ) , .ZN( us10_n603 ) , .A4( us10_n655 ) );
  AOI222_X1 us10_U61 (.ZN( us10_n606 ) , .A1( us10_n830 ) , .C2( us10_n837 ) , .B1( us10_n842 ) , .A2( us10_n856 ) , .B2( us10_n861 ) , .C1( us10_n868 ) );
  AOI222_X1 us10_U62 (.B2( us10_n638 ) , .ZN( us10_n644 ) , .B1( us10_n841 ) , .A1( us10_n842 ) , .C2( us10_n846 ) , .C1( us10_n863 ) , .A2( us10_n865 ) );
  NOR4_X1 us10_U63 (.A4( us10_n639 ) , .A3( us10_n640 ) , .A2( us10_n641 ) , .A1( us10_n642 ) , .ZN( us10_n643 ) );
  NOR3_X1 us10_U64 (.A2( us10_n607 ) , .A1( us10_n608 ) , .ZN( us10_n646 ) , .A3( us10_n722 ) );
  NAND4_X1 us10_U65 (.A4( us10_n657 ) , .A3( us10_n658 ) , .A2( us10_n659 ) , .A1( us10_n660 ) , .ZN( us10_n800 ) );
  NOR3_X1 us10_U66 (.A3( us10_n648 ) , .A2( us10_n649 ) , .A1( us10_n650 ) , .ZN( us10_n659 ) );
  NOR3_X1 us10_U67 (.A3( us10_n651 ) , .A2( us10_n652 ) , .A1( us10_n653 ) , .ZN( us10_n658 ) );
  NOR3_X1 us10_U68 (.A3( us10_n654 ) , .A2( us10_n655 ) , .A1( us10_n656 ) , .ZN( us10_n657 ) );
  NAND4_X1 us10_U69 (.A4( us10_n560 ) , .A3( us10_n561 ) , .A2( us10_n562 ) , .A1( us10_n563 ) , .ZN( us10_n607 ) );
  INV_X1 us10_U7 (.A( us10_n706 ) , .ZN( us10_n876 ) );
  NOR4_X1 us10_U70 (.A4( us10_n552 ) , .A3( us10_n553 ) , .A2( us10_n554 ) , .A1( us10_n555 ) , .ZN( us10_n562 ) );
  NOR4_X1 us10_U71 (.A4( us10_n556 ) , .A3( us10_n557 ) , .A2( us10_n558 ) , .A1( us10_n559 ) , .ZN( us10_n560 ) );
  NOR4_X1 us10_U72 (.ZN( us10_n561 ) , .A1( us10_n653 ) , .A3( us10_n661 ) , .A4( us10_n685 ) , .A2( us10_n768 ) );
  NAND4_X1 us10_U73 (.A4( us10_n772 ) , .A3( us10_n773 ) , .A2( us10_n774 ) , .A1( us10_n775 ) , .ZN( us10_n801 ) );
  NOR3_X1 us10_U74 (.A3( us10_n765 ) , .A2( us10_n766 ) , .A1( us10_n767 ) , .ZN( us10_n773 ) );
  NOR4_X1 us10_U75 (.A4( us10_n768 ) , .A3( us10_n769 ) , .A2( us10_n770 ) , .A1( us10_n771 ) , .ZN( us10_n772 ) );
  AOI222_X1 us10_U76 (.ZN( us10_n775 ) , .A1( us10_n830 ) , .C1( us10_n834 ) , .B2( us10_n841 ) , .A2( us10_n850 ) , .B1( us10_n861 ) , .C2( us10_n873 ) );
  NOR4_X1 us10_U77 (.A4( us10_n665 ) , .A3( us10_n666 ) , .A2( us10_n667 ) , .A1( us10_n668 ) , .ZN( us10_n676 ) );
  NOR4_X1 us10_U78 (.A4( us10_n661 ) , .A3( us10_n662 ) , .A2( us10_n663 ) , .A1( us10_n664 ) , .ZN( us10_n677 ) );
  NOR4_X1 us10_U79 (.A3( us10_n673 ) , .A1( us10_n674 ) , .ZN( us10_n675 ) , .A4( us10_n715 ) , .A2( us10_n859 ) );
  NOR3_X1 us10_U8 (.A3( us10_n621 ) , .A2( us10_n622 ) , .ZN( us10_n636 ) , .A1( us10_n725 ) );
  NOR2_X1 us10_U80 (.ZN( us10_n761 ) , .A1( us10_n833 ) , .A2( us10_n834 ) );
  NOR4_X1 us10_U81 (.A4( us10_n577 ) , .A3( us10_n578 ) , .A2( us10_n579 ) , .ZN( us10_n586 ) , .A1( us10_n683 ) );
  NOR4_X1 us10_U82 (.A1( us10_n584 ) , .ZN( us10_n585 ) , .A3( us10_n652 ) , .A2( us10_n662 ) , .A4( us10_n767 ) );
  AOI222_X1 us10_U83 (.ZN( us10_n513 ) , .C1( us10_n832 ) , .B2( us10_n837 ) , .A2( us10_n843 ) , .C2( us10_n862 ) , .B1( us10_n863 ) , .A1( us10_n866 ) );
  NOR4_X1 us10_U84 (.A4( us10_n509 ) , .A2( us10_n510 ) , .A1( us10_n511 ) , .ZN( us10_n512 ) , .A3( us10_n670 ) );
  INV_X1 us10_U85 (.A( us10_n505 ) , .ZN( us10_n871 ) );
  NAND4_X1 us10_U86 (.A4( us10_n456 ) , .A3( us10_n457 ) , .A2( us10_n458 ) , .A1( us10_n459 ) , .ZN( us10_n679 ) );
  NOR3_X1 us10_U87 (.ZN( us10_n457 ) , .A3( us10_n530 ) , .A1( us10_n555 ) , .A2( us10_n570 ) );
  NOR4_X1 us10_U88 (.ZN( us10_n458 ) , .A2( us10_n509 ) , .A1( us10_n599 ) , .A4( us10_n628 ) , .A3( us10_n711 ) );
  NOR4_X1 us10_U89 (.ZN( us10_n456 ) , .A2( us10_n517 ) , .A1( us10_n543 ) , .A3( us10_n579 ) , .A4( us10_n615 ) );
  NOR2_X1 us10_U9 (.ZN( us10_n575 ) , .A1( us10_n622 ) , .A2( us10_n745 ) );
  NAND4_X1 us10_U90 (.A4( us10_n535 ) , .A3( us10_n536 ) , .A2( us10_n537 ) , .A1( us10_n538 ) , .ZN( us10_n622 ) );
  NOR4_X1 us10_U91 (.A4( us10_n526 ) , .A2( us10_n527 ) , .A1( us10_n528 ) , .ZN( us10_n538 ) , .A3( us10_n701 ) );
  NOR4_X1 us10_U92 (.A1( us10_n531 ) , .ZN( us10_n536 ) , .A2( us10_n654 ) , .A4( us10_n668 ) , .A3( us10_n765 ) );
  NOR4_X1 us10_U93 (.A4( us10_n529 ) , .A3( us10_n530 ) , .ZN( us10_n537 ) , .A2( us10_n684 ) , .A1( us10_n794 ) );
  NOR2_X1 us10_U94 (.ZN( us10_n686 ) , .A1( us10_n831 ) , .A2( us10_n832 ) );
  NAND4_X1 us10_U95 (.A4( us10_n479 ) , .A3( us10_n480 ) , .A2( us10_n481 ) , .A1( us10_n482 ) , .ZN( us10_n694 ) );
  NOR3_X1 us10_U96 (.ZN( us10_n480 ) , .A2( us10_n508 ) , .A3( us10_n601 ) , .A1( us10_n610 ) );
  AOI211_X1 us10_U97 (.B( us10_n477 ) , .A( us10_n478 ) , .ZN( us10_n482 ) , .C2( us10_n833 ) , .C1( us10_n861 ) );
  NOR4_X1 us10_U98 (.ZN( us10_n481 ) , .A3( us10_n532 ) , .A4( us10_n545 ) , .A2( us10_n567 ) , .A1( us10_n717 ) );
  NAND4_X1 us10_U99 (.A4( us10_n548 ) , .A3( us10_n549 ) , .A2( us10_n550 ) , .A1( us10_n551 ) , .ZN( us10_n745 ) );
  NOR3_X1 us11_U10 (.ZN( us11_n504 ) , .A2( us11_n679 ) , .A3( us11_n777 ) , .A1( us11_n876 ) );
  NOR4_X1 us11_U100 (.A4( us11_n529 ) , .A3( us11_n530 ) , .ZN( us11_n537 ) , .A2( us11_n684 ) , .A1( us11_n794 ) );
  NAND4_X1 us11_U101 (.A4( us11_n479 ) , .A3( us11_n480 ) , .A2( us11_n481 ) , .A1( us11_n482 ) , .ZN( us11_n694 ) );
  NOR3_X1 us11_U102 (.ZN( us11_n480 ) , .A2( us11_n508 ) , .A3( us11_n601 ) , .A1( us11_n610 ) );
  AOI211_X1 us11_U103 (.B( us11_n477 ) , .A( us11_n478 ) , .ZN( us11_n482 ) , .C2( us11_n833 ) , .C1( us11_n861 ) );
  NOR4_X1 us11_U104 (.ZN( us11_n481 ) , .A3( us11_n532 ) , .A4( us11_n545 ) , .A2( us11_n567 ) , .A1( us11_n717 ) );
  NAND4_X1 us11_U105 (.A4( us11_n548 ) , .A3( us11_n549 ) , .A2( us11_n550 ) , .A1( us11_n551 ) , .ZN( us11_n745 ) );
  NOR3_X1 us11_U106 (.ZN( us11_n549 ) , .A2( us11_n651 ) , .A1( us11_n667 ) , .A3( us11_n771 ) );
  AOI211_X1 us11_U107 (.B( us11_n539 ) , .A( us11_n540 ) , .ZN( us11_n551 ) , .C2( us11_n839 ) , .C1( us11_n851 ) );
  NOR4_X1 us11_U108 (.A4( us11_n544 ) , .A3( us11_n545 ) , .A2( us11_n546 ) , .A1( us11_n547 ) , .ZN( us11_n548 ) );
  NOR4_X1 us11_U109 (.ZN( us11_n620 ) , .A1( us11_n656 ) , .A3( us11_n666 ) , .A4( us11_n682 ) , .A2( us11_n766 ) );
  INV_X1 us11_U11 (.A( us11_n706 ) , .ZN( us11_n876 ) );
  NOR4_X1 us11_U110 (.A4( us11_n609 ) , .A3( us11_n610 ) , .A2( us11_n611 ) , .A1( us11_n612 ) , .ZN( us11_n619 ) );
  NOR4_X1 us11_U111 (.A4( us11_n614 ) , .A3( us11_n615 ) , .A2( us11_n616 ) , .A1( us11_n617 ) , .ZN( us11_n618 ) );
  NOR2_X1 us11_U112 (.ZN( us11_n686 ) , .A1( us11_n831 ) , .A2( us11_n832 ) );
  NAND4_X1 us11_U113 (.A4( us11_n473 ) , .A3( us11_n474 ) , .A2( us11_n475 ) , .A1( us11_n476 ) , .ZN( us11_n678 ) );
  NOR4_X1 us11_U114 (.A4( us11_n470 ) , .ZN( us11_n476 ) , .A3( us11_n556 ) , .A1( us11_n735 ) , .A2( us11_n755 ) );
  NOR4_X1 us11_U115 (.ZN( us11_n475 ) , .A1( us11_n531 ) , .A3( us11_n568 ) , .A4( us11_n600 ) , .A2( us11_n642 ) );
  NOR4_X1 us11_U116 (.ZN( us11_n474 ) , .A1( us11_n506 ) , .A3( us11_n544 ) , .A2( us11_n583 ) , .A4( us11_n716 ) );
  NAND4_X1 us11_U117 (.A4( us11_n691 ) , .A3( us11_n692 ) , .A1( us11_n693 ) , .ZN( us11_n776 ) , .A2( us11_n872 ) );
  INV_X1 us11_U118 (.A( us11_n679 ) , .ZN( us11_n872 ) );
  NOR4_X1 us11_U119 (.A4( us11_n687 ) , .A3( us11_n688 ) , .A2( us11_n689 ) , .A1( us11_n690 ) , .ZN( us11_n691 ) );
  NOR3_X1 us11_U12 (.A3( us11_n621 ) , .A2( us11_n622 ) , .ZN( us11_n636 ) , .A1( us11_n725 ) );
  AOI221_X1 us11_U120 (.A( us11_n681 ) , .ZN( us11_n692 ) , .B2( us11_n840 ) , .C1( us11_n842 ) , .C2( us11_n862 ) , .B1( us11_n865 ) );
  NOR2_X1 us11_U121 (.ZN( us11_n733 ) , .A2( us11_n832 ) , .A1( us11_n845 ) );
  NAND4_X1 us11_U122 (.A4( us11_n719 ) , .A3( us11_n720 ) , .A2( us11_n721 ) , .ZN( us11_n741 ) , .A1( us11_n857 ) );
  AOI221_X1 us11_U123 (.A( us11_n710 ) , .ZN( us11_n721 ) , .C2( us11_n844 ) , .B2( us11_n845 ) , .C1( us11_n861 ) , .B1( us11_n862 ) );
  INV_X1 us11_U124 (.A( us11_n709 ) , .ZN( us11_n857 ) );
  NOR4_X1 us11_U125 (.A4( us11_n715 ) , .A3( us11_n716 ) , .A2( us11_n717 ) , .A1( us11_n718 ) , .ZN( us11_n719 ) );
  NAND4_X1 us11_U126 (.A4( us11_n573 ) , .A3( us11_n574 ) , .A1( us11_n575 ) , .ZN( us11_n723 ) , .A2( us11_n874 ) );
  NOR4_X1 us11_U127 (.A4( us11_n569 ) , .A3( us11_n570 ) , .A2( us11_n571 ) , .A1( us11_n572 ) , .ZN( us11_n573 ) );
  INV_X1 us11_U128 (.A( us11_n607 ) , .ZN( us11_n874 ) );
  NOR2_X1 us11_U129 (.ZN( us11_n575 ) , .A1( us11_n622 ) , .A2( us11_n745 ) );
  NOR2_X1 us11_U13 (.ZN( us11_n495 ) , .A1( us11_n678 ) , .A2( us11_n694 ) );
  NAND4_X1 us11_U130 (.A4( us11_n493 ) , .A3( us11_n494 ) , .A1( us11_n495 ) , .ZN( us11_n802 ) , .A2( us11_n867 ) );
  AOI221_X1 us11_U131 (.A( us11_n489 ) , .ZN( us11_n494 ) , .B2( us11_n836 ) , .C2( us11_n841 ) , .C1( us11_n851 ) , .B1( us11_n860 ) );
  INV_X1 us11_U132 (.A( us11_n778 ) , .ZN( us11_n867 ) );
  NOR4_X1 us11_U133 (.A2( us11_n491 ) , .A1( us11_n492 ) , .ZN( us11_n493 ) , .A3( us11_n580 ) , .A4( us11_n612 ) );
  NOR2_X1 us11_U134 (.ZN( us11_n647 ) , .A1( us11_n854 ) , .A2( us11_n868 ) );
  INV_X1 us11_U135 (.A( us11_n762 ) , .ZN( us11_n830 ) );
  NAND4_X1 us11_U136 (.A4( us11_n633 ) , .A3( us11_n634 ) , .A2( us11_n635 ) , .A1( us11_n636 ) , .ZN( us11_n743 ) );
  AOI211_X1 us11_U137 (.B( us11_n623 ) , .A( us11_n624 ) , .ZN( us11_n635 ) , .C2( us11_n836 ) , .C1( us11_n863 ) );
  NOR4_X1 us11_U138 (.A4( us11_n629 ) , .A3( us11_n630 ) , .A2( us11_n631 ) , .A1( us11_n632 ) , .ZN( us11_n633 ) );
  NOR4_X1 us11_U139 (.A4( us11_n626 ) , .A3( us11_n627 ) , .A2( us11_n628 ) , .ZN( us11_n634 ) , .A1( us11_n664 ) );
  NOR2_X1 us11_U14 (.A1( us11_n678 ) , .ZN( us11_n693 ) , .A2( us11_n807 ) );
  OR4_X1 us11_U140 (.A4( us11_n566 ) , .A3( us11_n567 ) , .A2( us11_n568 ) , .ZN( us11_n572 ) , .A1( us11_n665 ) );
  OR4_X1 us11_U141 (.A4( us11_n518 ) , .A2( us11_n519 ) , .A1( us11_n520 ) , .ZN( us11_n522 ) , .A3( us11_n821 ) );
  OR4_X1 us11_U142 (.ZN( us11_n492 ) , .A4( us11_n534 ) , .A2( us11_n547 ) , .A1( us11_n559 ) , .A3( us11_n632 ) );
  OR4_X1 us11_U143 (.A4( us11_n682 ) , .A3( us11_n683 ) , .A2( us11_n684 ) , .A1( us11_n685 ) , .ZN( us11_n690 ) );
  OR4_X1 us11_U144 (.ZN( us11_n466 ) , .A4( us11_n518 ) , .A3( us11_n529 ) , .A2( us11_n578 ) , .A1( us11_n712 ) );
  INV_X1 us11_U145 (.A( us11_n697 ) , .ZN( us11_n838 ) );
  OR4_X1 us11_U146 (.A4( us11_n580 ) , .A3( us11_n581 ) , .A2( us11_n582 ) , .A1( us11_n583 ) , .ZN( us11_n584 ) );
  NAND2_X1 us11_U147 (.ZN( us11_n613 ) , .A2( us11_n837 ) , .A1( us11_n873 ) );
  OR3_X1 us11_U148 (.A3( us11_n506 ) , .A2( us11_n507 ) , .A1( us11_n508 ) , .ZN( us11_n511 ) );
  INV_X1 us11_U149 (.A( us11_n463 ) , .ZN( us11_n864 ) );
  INV_X1 us11_U15 (.A( us11_n680 ) , .ZN( us11_n840 ) );
  OAI21_X1 us11_U150 (.ZN( us11_n463 ) , .B1( us11_n809 ) , .A( us11_n834 ) , .B2( us11_n851 ) );
  INV_X1 us11_U151 (.A( us11_n754 ) , .ZN( us11_n869 ) );
  OAI21_X1 us11_U152 (.B1( us11_n753 ) , .ZN( us11_n754 ) , .A( us11_n845 ) , .B2( us11_n868 ) );
  INV_X1 us11_U153 (.A( us11_n672 ) , .ZN( us11_n859 ) );
  AOI21_X1 us11_U154 (.A( us11_n670 ) , .B1( us11_n671 ) , .ZN( us11_n672 ) , .B2( us11_n856 ) );
  AOI222_X1 us11_U155 (.ZN( us11_n660 ) , .A2( us11_n839 ) , .B1( us11_n841 ) , .C2( us11_n845 ) , .A1( us11_n860 ) , .C1( us11_n863 ) , .B2( us11_n870 ) );
  INV_X1 us11_U156 (.A( us11_n647 ) , .ZN( us11_n870 ) );
  NAND2_X1 us11_U157 (.A1( us11_n447 ) , .A2( us11_n465 ) , .ZN( us11_n749 ) );
  OAI222_X1 us11_U158 (.ZN( us11_n617 ) , .B1( us11_n697 ) , .C1( us11_n724 ) , .C2( us11_n747 ) , .B2( us11_n786 ) , .A2( us11_n792 ) , .A1( us11_n816 ) );
  OAI222_X1 us11_U159 (.B2( us11_n708 ) , .ZN( us11_n709 ) , .C2( us11_n724 ) , .B1( us11_n747 ) , .A1( us11_n806 ) , .C1( us11_n814 ) , .A2( us11_n815 ) );
  NOR4_X1 us11_U16 (.A4( us11_n445 ) , .A3( us11_n446 ) , .A2( us11_n516 ) , .A1( us11_n541 ) , .ZN( us11_n706 ) );
  AOI22_X1 us11_U160 (.ZN( us11_n696 ) , .A1( us11_n830 ) , .B2( us11_n843 ) , .A2( us11_n865 ) , .B1( us11_n868 ) );
  AOI22_X1 us11_U161 (.A2( us11_n782 ) , .ZN( us11_n783 ) , .B2( us11_n831 ) , .A1( us11_n834 ) , .B1( us11_n863 ) );
  INV_X1 us11_U162 (.A( us11_n730 ) , .ZN( us11_n839 ) );
  AOI221_X1 us11_U163 (.A( us11_n564 ) , .C2( us11_n565 ) , .ZN( us11_n574 ) , .B2( us11_n845 ) , .B1( us11_n852 ) , .C1( us11_n853 ) );
  AOI21_X1 us11_U164 (.ZN( us11_n564 ) , .B1( us11_n724 ) , .A( us11_n779 ) , .B2( us11_n791 ) );
  NAND2_X1 us11_U165 (.A1( us11_n451 ) , .A2( us11_n453 ) , .ZN( us11_n762 ) );
  INV_X1 us11_U166 (.A( us11_n790 ) , .ZN( us11_n832 ) );
  OAI22_X1 us11_U167 (.ZN( us11_n637 ) , .A1( us11_n699 ) , .B2( us11_n728 ) , .A2( us11_n762 ) , .B1( us11_n816 ) );
  OAI221_X1 us11_U168 (.A( us11_n727 ) , .C2( us11_n728 ) , .B2( us11_n729 ) , .B1( us11_n730 ) , .ZN( us11_n737 ) , .C1( us11_n817 ) );
  AOI22_X1 us11_U169 (.ZN( us11_n727 ) , .B1( us11_n832 ) , .A2( us11_n838 ) , .A1( us11_n863 ) , .B2( us11_n866 ) );
  OR3_X1 us11_U17 (.ZN( us11_n446 ) , .A1( us11_n528 ) , .A3( us11_n577 ) , .A2( us11_n875 ) );
  INV_X1 us11_U170 (.A( us11_n747 ) , .ZN( us11_n834 ) );
  OAI22_X1 us11_U171 (.ZN( us11_n624 ) , .B1( us11_n669 ) , .B2( us11_n747 ) , .A1( us11_n815 ) , .A2( us11_n816 ) );
  OAI22_X1 us11_U172 (.ZN( us11_n489 ) , .A1( us11_n724 ) , .B2( us11_n728 ) , .B1( us11_n730 ) , .A2( us11_n779 ) );
  OAI22_X1 us11_U173 (.B2( us11_n779 ) , .B1( us11_n780 ) , .ZN( us11_n781 ) , .A2( us11_n814 ) , .A1( us11_n815 ) );
  OAI22_X1 us11_U174 (.A1( us11_n724 ) , .ZN( us11_n726 ) , .B2( us11_n750 ) , .B1( us11_n812 ) , .A2( us11_n816 ) );
  NOR2_X1 us11_U175 (.ZN( us11_n630 ) , .A1( us11_n747 ) , .A2( us11_n815 ) );
  OAI22_X1 us11_U176 (.B2( us11_n750 ) , .B1( us11_n751 ) , .A1( us11_n752 ) , .ZN( us11_n756 ) , .A2( us11_n806 ) );
  NOR3_X1 us11_U177 (.ZN( us11_n752 ) , .A2( us11_n853 ) , .A1( us11_n863 ) , .A3( us11_n865 ) );
  NOR2_X1 us11_U178 (.ZN( us11_n751 ) , .A2( us11_n852 ) , .A1( us11_n860 ) );
  OAI22_X1 us11_U179 (.B2( us11_n803 ) , .B1( us11_n804 ) , .A2( us11_n805 ) , .A1( us11_n806 ) , .ZN( us11_n808 ) );
  OR4_X1 us11_U18 (.A4( us11_n442 ) , .A2( us11_n443 ) , .A1( us11_n444 ) , .ZN( us11_n445 ) , .A3( us11_n553 ) );
  NOR2_X1 us11_U180 (.ZN( us11_n656 ) , .A1( us11_n747 ) , .A2( us11_n780 ) );
  OAI22_X1 us11_U181 (.B2( us11_n744 ) , .ZN( us11_n746 ) , .A2( us11_n762 ) , .B1( us11_n780 ) , .A1( us11_n792 ) );
  OAI22_X1 us11_U182 (.ZN( us11_n496 ) , .A2( us11_n744 ) , .A1( us11_n780 ) , .B1( us11_n791 ) , .B2( us11_n806 ) );
  OAI22_X1 us11_U183 (.ZN( us11_n695 ) , .A2( us11_n730 ) , .A1( us11_n780 ) , .B1( us11_n791 ) , .B2( us11_n817 ) );
  INV_X1 us11_U184 (.A( us11_n744 ) , .ZN( us11_n837 ) );
  INV_X1 us11_U185 (.A( us11_n805 ) , .ZN( us11_n860 ) );
  INV_X1 us11_U186 (.A( us11_n816 ) , .ZN( us11_n831 ) );
  INV_X1 us11_U187 (.A( us11_n788 ) , .ZN( us11_n845 ) );
  OAI22_X1 us11_U188 (.ZN( us11_n590 ) , .B1( us11_n730 ) , .B2( us11_n749 ) , .A2( us11_n786 ) , .A1( us11_n803 ) );
  OAI22_X1 us11_U189 (.B1( us11_n490 ) , .ZN( us11_n491 ) , .A1( us11_n686 ) , .A2( us11_n763 ) , .B2( us11_n817 ) );
  INV_X1 us11_U19 (.A( us11_n613 ) , .ZN( us11_n875 ) );
  NOR3_X1 us11_U190 (.ZN( us11_n490 ) , .A1( us11_n782 ) , .A2( us11_n850 ) , .A3( us11_n863 ) );
  OAI22_X1 us11_U191 (.ZN( us11_n710 ) , .A2( us11_n728 ) , .B2( us11_n729 ) , .A1( us11_n744 ) , .B1( us11_n813 ) );
  INV_X1 us11_U192 (.A( us11_n792 ) , .ZN( us11_n851 ) );
  NOR2_X1 us11_U193 (.ZN( us11_n715 ) , .A1( us11_n805 ) , .A2( us11_n817 ) );
  NOR2_X1 us11_U194 (.A1( us11_n699 ) , .ZN( us11_n768 ) , .A2( us11_n813 ) );
  NOR2_X1 us11_U195 (.ZN( us11_n541 ) , .A2( us11_n697 ) , .A1( us11_n699 ) );
  INV_X1 us11_U196 (.A( us11_n814 ) , .ZN( us11_n833 ) );
  NOR2_X1 us11_U197 (.A1( us11_n669 ) , .ZN( us11_n673 ) , .A2( us11_n744 ) );
  NOR2_X1 us11_U198 (.ZN( us11_n602 ) , .A1( us11_n669 ) , .A2( us11_n803 ) );
  NOR2_X1 us11_U199 (.A1( us11_n669 ) , .ZN( us11_n688 ) , .A2( us11_n816 ) );
  INV_X1 us11_U20 (.A( us11_n749 ) , .ZN( us11_n863 ) );
  NOR2_X1 us11_U200 (.A2( us11_n744 ) , .ZN( us11_n755 ) , .A1( us11_n805 ) );
  NOR2_X1 us11_U201 (.ZN( us11_n735 ) , .A2( us11_n803 ) , .A1( us11_n805 ) );
  NOR2_X1 us11_U202 (.A1( us11_n669 ) , .ZN( us11_n766 ) , .A2( us11_n813 ) );
  NOR2_X1 us11_U203 (.ZN( us11_n527 ) , .A1( us11_n669 ) , .A2( us11_n779 ) );
  NOR2_X1 us11_U204 (.ZN( us11_n666 ) , .A1( us11_n728 ) , .A2( us11_n803 ) );
  NOR2_X1 us11_U205 (.ZN( us11_n594 ) , .A2( us11_n697 ) , .A1( us11_n728 ) );
  NOR2_X1 us11_U206 (.ZN( us11_n718 ) , .A2( us11_n724 ) , .A1( us11_n744 ) );
  NOR2_X1 us11_U207 (.ZN( us11_n570 ) , .A1( us11_n728 ) , .A2( us11_n806 ) );
  NOR2_X1 us11_U208 (.ZN( us11_n661 ) , .A1( us11_n729 ) , .A2( us11_n790 ) );
  OAI22_X1 us11_U209 (.ZN( us11_n483 ) , .A1( us11_n708 ) , .B2( us11_n785 ) , .A2( us11_n806 ) , .B1( us11_n812 ) );
  AOI222_X1 us11_U21 (.ZN( us11_n563 ) , .B1( us11_n830 ) , .C1( us11_n841 ) , .A2( us11_n843 ) , .A1( us11_n854 ) , .B2( us11_n863 ) , .C2( us11_n873 ) );
  NOR2_X1 us11_U210 (.ZN( us11_n601 ) , .A2( us11_n780 ) , .A1( us11_n803 ) );
  NOR2_X1 us11_U211 (.ZN( us11_n531 ) , .A2( us11_n780 ) , .A1( us11_n816 ) );
  NOR2_X1 us11_U212 (.ZN( us11_n654 ) , .A1( us11_n728 ) , .A2( us11_n813 ) );
  NOR2_X1 us11_U213 (.ZN( us11_n509 ) , .A1( us11_n729 ) , .A2( us11_n779 ) );
  NOR2_X1 us11_U214 (.ZN( us11_n599 ) , .A2( us11_n791 ) , .A1( us11_n816 ) );
  NOR2_X1 us11_U215 (.ZN( us11_n612 ) , .A1( us11_n779 ) , .A2( us11_n786 ) );
  NOR2_X1 us11_U216 (.ZN( us11_n546 ) , .A2( us11_n780 ) , .A1( us11_n814 ) );
  INV_X1 us11_U217 (.A( us11_n750 ) , .ZN( us11_n842 ) );
  NOR2_X1 us11_U218 (.ZN( us11_n532 ) , .A2( us11_n749 ) , .A1( us11_n750 ) );
  NOR2_X1 us11_U219 (.ZN( us11_n528 ) , .A2( us11_n724 ) , .A1( us11_n803 ) );
  NOR4_X1 us11_U22 (.ZN( us11_n479 ) , .A1( us11_n520 ) , .A4( us11_n557 ) , .A3( us11_n582 ) , .A2( us11_n630 ) );
  NOR2_X1 us11_U220 (.ZN( us11_n577 ) , .A2( us11_n699 ) , .A1( us11_n814 ) );
  AOI21_X1 us11_U221 (.ZN( us11_n640 ) , .B2( us11_n747 ) , .A( us11_n792 ) , .B1( us11_n803 ) );
  NOR2_X1 us11_U222 (.ZN( us11_n615 ) , .A1( us11_n785 ) , .A2( us11_n815 ) );
  NOR2_X1 us11_U223 (.ZN( us11_n629 ) , .A2( us11_n728 ) , .A1( us11_n785 ) );
  NOR2_X1 us11_U224 (.ZN( us11_n663 ) , .A1( us11_n729 ) , .A2( us11_n785 ) );
  NOR2_X1 us11_U225 (.ZN( us11_n628 ) , .A2( us11_n669 ) , .A1( us11_n785 ) );
  NOR2_X1 us11_U226 (.ZN( us11_n611 ) , .A2( us11_n780 ) , .A1( us11_n806 ) );
  NOR2_X1 us11_U227 (.A2( us11_n744 ) , .ZN( us11_n769 ) , .A1( us11_n812 ) );
  NOR2_X1 us11_U228 (.ZN( us11_n567 ) , .A1( us11_n747 ) , .A2( us11_n805 ) );
  NOR2_X1 us11_U229 (.A2( us11_n708 ) , .A1( us11_n750 ) , .ZN( us11_n771 ) );
  NOR4_X1 us11_U23 (.ZN( us11_n473 ) , .A2( us11_n521 ) , .A4( us11_n594 ) , .A1( us11_n609 ) , .A3( us11_n629 ) );
  NOR2_X1 us11_U230 (.ZN( us11_n557 ) , .A1( us11_n792 ) , .A2( us11_n814 ) );
  NOR2_X1 us11_U231 (.A2( us11_n697 ) , .ZN( us11_n716 ) , .A1( us11_n792 ) );
  NOR2_X1 us11_U232 (.ZN( us11_n544 ) , .A2( us11_n785 ) , .A1( us11_n792 ) );
  NOR2_X1 us11_U233 (.ZN( us11_n667 ) , .A1( us11_n750 ) , .A2( us11_n815 ) );
  NOR2_X1 us11_U234 (.ZN( us11_n555 ) , .A1( us11_n750 ) , .A2( us11_n791 ) );
  NOR2_X1 us11_U235 (.ZN( us11_n508 ) , .A2( us11_n780 ) , .A1( us11_n785 ) );
  NOR2_X1 us11_U236 (.ZN( us11_n543 ) , .A2( us11_n708 ) , .A1( us11_n785 ) );
  NOR2_X1 us11_U237 (.ZN( us11_n664 ) , .A1( us11_n785 ) , .A2( us11_n791 ) );
  OAI22_X1 us11_U238 (.B1( us11_n440 ) , .ZN( us11_n444 ) , .A2( us11_n728 ) , .A1( us11_n744 ) , .B2( us11_n749 ) );
  NOR3_X1 us11_U239 (.ZN( us11_n440 ) , .A2( us11_n836 ) , .A3( us11_n837 ) , .A1( us11_n846 ) );
  NOR4_X1 us11_U24 (.ZN( us11_n485 ) , .A2( us11_n533 ) , .A1( us11_n558 ) , .A3( us11_n631 ) , .A4( us11_n718 ) );
  NOR2_X1 us11_U240 (.ZN( us11_n631 ) , .A1( us11_n724 ) , .A2( us11_n813 ) );
  NOR2_X1 us11_U241 (.ZN( us11_n556 ) , .A1( us11_n762 ) , .A2( us11_n805 ) );
  NOR2_X1 us11_U242 (.ZN( us11_n530 ) , .A2( us11_n744 ) , .A1( us11_n792 ) );
  NOR2_X1 us11_U243 (.ZN( us11_n507 ) , .A1( us11_n812 ) , .A2( us11_n817 ) );
  NOR2_X1 us11_U244 (.ZN( us11_n516 ) , .A1( us11_n708 ) , .A2( us11_n744 ) );
  NOR2_X1 us11_U245 (.ZN( us11_n558 ) , .A1( us11_n708 ) , .A2( us11_n816 ) );
  NOR2_X1 us11_U246 (.ZN( us11_n517 ) , .A1( us11_n708 ) , .A2( us11_n803 ) );
  INV_X1 us11_U247 (.A( us11_n806 ) , .ZN( us11_n841 ) );
  NOR2_X1 us11_U248 (.ZN( us11_n545 ) , .A1( us11_n749 ) , .A2( us11_n814 ) );
  INV_X1 us11_U249 (.A( us11_n728 ) , .ZN( us11_n852 ) );
  NOR4_X1 us11_U25 (.A4( us11_n532 ) , .A3( us11_n533 ) , .A2( us11_n534 ) , .ZN( us11_n535 ) , .A1( us11_n820 ) );
  NOR2_X1 us11_U250 (.ZN( us11_n554 ) , .A1( us11_n786 ) , .A2( us11_n813 ) );
  NOR2_X1 us11_U251 (.ZN( us11_n670 ) , .A1( us11_n790 ) , .A2( us11_n805 ) );
  NOR2_X1 us11_U252 (.ZN( us11_n717 ) , .A2( us11_n744 ) , .A1( us11_n786 ) );
  NOR2_X1 us11_U253 (.ZN( us11_n506 ) , .A2( us11_n728 ) , .A1( us11_n762 ) );
  NOR2_X1 us11_U254 (.ZN( us11_n642 ) , .A2( us11_n788 ) , .A1( us11_n791 ) );
  NOR2_X1 us11_U255 (.ZN( us11_n614 ) , .A1( us11_n762 ) , .A2( us11_n812 ) );
  AOI21_X1 us11_U256 (.ZN( us11_n626 ) , .B2( us11_n669 ) , .A( us11_n790 ) , .B1( us11_n791 ) );
  AOI21_X1 us11_U257 (.ZN( us11_n552 ) , .B1( us11_n669 ) , .A( us11_n697 ) , .B2( us11_n805 ) );
  AOI21_X1 us11_U258 (.ZN( us11_n589 ) , .B2( us11_n699 ) , .B1( us11_n815 ) , .A( us11_n817 ) );
  INV_X1 us11_U259 (.A( us11_n763 ) , .ZN( us11_n866 ) );
  NOR4_X1 us11_U26 (.ZN( us11_n456 ) , .A2( us11_n517 ) , .A1( us11_n543 ) , .A3( us11_n579 ) , .A4( us11_n615 ) );
  NOR2_X1 us11_U260 (.ZN( us11_n609 ) , .A2( us11_n724 ) , .A1( us11_n817 ) );
  NOR2_X1 us11_U261 (.ZN( us11_n668 ) , .A2( us11_n708 ) , .A1( us11_n790 ) );
  NOR2_X1 us11_U262 (.ZN( us11_n533 ) , .A2( us11_n724 ) , .A1( us11_n730 ) );
  NOR2_X1 us11_U263 (.ZN( us11_n521 ) , .A1( us11_n790 ) , .A2( us11_n812 ) );
  AOI21_X1 us11_U264 (.A( us11_n815 ) , .B2( us11_n816 ) , .B1( us11_n817 ) , .ZN( us11_n818 ) );
  NOR2_X1 us11_U265 (.ZN( us11_n547 ) , .A1( us11_n699 ) , .A2( us11_n744 ) );
  AOI21_X1 us11_U266 (.ZN( us11_n510 ) , .B2( us11_n669 ) , .A( us11_n730 ) , .B1( us11_n815 ) );
  NOR2_X1 us11_U267 (.ZN( us11_n655 ) , .A1( us11_n790 ) , .A2( us11_n815 ) );
  NOR2_X1 us11_U268 (.ZN( us11_n579 ) , .A2( us11_n708 ) , .A1( us11_n730 ) );
  INV_X1 us11_U269 (.A( us11_n729 ) , .ZN( us11_n868 ) );
  NOR4_X1 us11_U27 (.A4( us11_n577 ) , .A3( us11_n578 ) , .A2( us11_n579 ) , .ZN( us11_n586 ) , .A1( us11_n683 ) );
  NOR2_X1 us11_U270 (.ZN( us11_n542 ) , .A1( us11_n762 ) , .A2( us11_n791 ) );
  NOR2_X1 us11_U271 (.ZN( us11_n701 ) , .A2( us11_n786 ) , .A1( us11_n817 ) );
  NOR2_X1 us11_U272 (.A2( us11_n708 ) , .A1( us11_n762 ) , .ZN( us11_n794 ) );
  AOI21_X1 us11_U273 (.ZN( us11_n499 ) , .B1( us11_n680 ) , .A( us11_n812 ) , .B2( us11_n816 ) );
  AOI21_X1 us11_U274 (.ZN( us11_n650 ) , .A( us11_n779 ) , .B1( us11_n792 ) , .B2( us11_n805 ) );
  INV_X1 us11_U275 (.A( us11_n699 ) , .ZN( us11_n853 ) );
  NOR2_X1 us11_U276 (.ZN( us11_n652 ) , .A1( us11_n669 ) , .A2( us11_n814 ) );
  NOR2_X1 us11_U277 (.ZN( us11_n581 ) , .A1( us11_n669 ) , .A2( us11_n788 ) );
  AOI21_X1 us11_U278 (.ZN( us11_n515 ) , .A( us11_n729 ) , .B1( us11_n750 ) , .B2( us11_n803 ) );
  AOI21_X1 us11_U279 (.B1( us11_n699 ) , .ZN( us11_n700 ) , .A( us11_n732 ) , .B2( us11_n763 ) );
  AOI222_X1 us11_U28 (.B2( us11_n638 ) , .ZN( us11_n644 ) , .B1( us11_n841 ) , .A1( us11_n842 ) , .C2( us11_n846 ) , .C1( us11_n863 ) , .A2( us11_n865 ) );
  AOI21_X1 us11_U280 (.ZN( us11_n591 ) , .B2( us11_n763 ) , .A( us11_n785 ) , .B1( us11_n812 ) );
  AOI21_X1 us11_U281 (.A( us11_n812 ) , .B2( us11_n813 ) , .B1( us11_n814 ) , .ZN( us11_n819 ) );
  NOR2_X1 us11_U282 (.A1( us11_n730 ) , .ZN( us11_n765 ) , .A2( us11_n786 ) );
  INV_X1 us11_U283 (.A( us11_n791 ) , .ZN( us11_n873 ) );
  AOI21_X1 us11_U284 (.ZN( us11_n593 ) , .B1( us11_n750 ) , .A( us11_n792 ) , .B2( us11_n813 ) );
  NOR2_X1 us11_U285 (.ZN( us11_n582 ) , .A1( us11_n744 ) , .A2( us11_n815 ) );
  NOR2_X1 us11_U286 (.ZN( us11_n519 ) , .A2( us11_n699 ) , .A1( us11_n816 ) );
  NOR2_X1 us11_U287 (.ZN( us11_n685 ) , .A1( us11_n729 ) , .A2( us11_n816 ) );
  NOR2_X1 us11_U288 (.ZN( us11_n559 ) , .A2( us11_n791 ) , .A1( us11_n803 ) );
  AOI21_X1 us11_U289 (.ZN( us11_n649 ) , .B1( us11_n729 ) , .B2( us11_n763 ) , .A( us11_n813 ) );
  NOR4_X1 us11_U29 (.A4( us11_n639 ) , .A3( us11_n640 ) , .A2( us11_n641 ) , .A1( us11_n642 ) , .ZN( us11_n643 ) );
  AOI21_X1 us11_U290 (.B1( us11_n625 ) , .ZN( us11_n627 ) , .A( us11_n763 ) , .B2( us11_n814 ) );
  NOR2_X1 us11_U291 (.ZN( us11_n683 ) , .A2( us11_n699 ) , .A1( us11_n803 ) );
  NOR2_X1 us11_U292 (.A2( us11_n697 ) , .A1( us11_n780 ) , .ZN( us11_n820 ) );
  NOR2_X1 us11_U293 (.ZN( us11_n653 ) , .A1( us11_n762 ) , .A2( us11_n786 ) );
  NOR2_X1 us11_U294 (.ZN( us11_n568 ) , .A1( us11_n729 ) , .A2( us11_n762 ) );
  NOR2_X1 us11_U295 (.ZN( us11_n662 ) , .A2( us11_n697 ) , .A1( us11_n729 ) );
  INV_X1 us11_U296 (.A( us11_n813 ) , .ZN( us11_n836 ) );
  NOR2_X1 us11_U297 (.ZN( us11_n566 ) , .A2( us11_n697 ) , .A1( us11_n763 ) );
  NOR2_X1 us11_U298 (.ZN( us11_n520 ) , .A2( us11_n708 ) , .A1( us11_n814 ) );
  AOI21_X1 us11_U299 (.ZN( us11_n477 ) , .A( us11_n669 ) , .B1( us11_n750 ) , .B2( us11_n806 ) );
  NAND2_X2 us11_U3 (.A2( us11_n460 ) , .A1( us11_n465 ) , .ZN( us11_n780 ) );
  NOR3_X1 us11_U30 (.A2( us11_n607 ) , .A1( us11_n608 ) , .ZN( us11_n646 ) , .A3( us11_n722 ) );
  NOR2_X1 us11_U300 (.A1( us11_n697 ) , .ZN( us11_n770 ) , .A2( us11_n815 ) );
  AOI21_X1 us11_U301 (.ZN( us11_n514 ) , .A( us11_n779 ) , .B2( us11_n792 ) , .B1( us11_n812 ) );
  INV_X1 us11_U302 (.A( us11_n786 ) , .ZN( us11_n862 ) );
  AOI21_X1 us11_U303 (.ZN( us11_n540 ) , .A( us11_n763 ) , .B2( us11_n779 ) , .B1( us11_n817 ) );
  AOI21_X1 us11_U304 (.ZN( us11_n450 ) , .B2( us11_n792 ) , .A( us11_n803 ) , .B1( us11_n815 ) );
  AOI21_X1 us11_U305 (.ZN( us11_n539 ) , .B2( us11_n812 ) , .A( us11_n814 ) , .B1( us11_n815 ) );
  NOR2_X1 us11_U306 (.ZN( us11_n529 ) , .A1( us11_n708 ) , .A2( us11_n779 ) );
  NOR2_X1 us11_U307 (.ZN( us11_n578 ) , .A1( us11_n708 ) , .A2( us11_n813 ) );
  NOR2_X1 us11_U308 (.ZN( us11_n583 ) , .A1( us11_n792 ) , .A2( us11_n817 ) );
  NOR2_X1 us11_U309 (.ZN( us11_n534 ) , .A1( us11_n724 ) , .A2( us11_n788 ) );
  NOR4_X1 us11_U31 (.A4( us11_n541 ) , .A3( us11_n542 ) , .A2( us11_n543 ) , .ZN( us11_n550 ) , .A1( us11_n688 ) );
  NOR2_X1 us11_U310 (.ZN( us11_n632 ) , .A2( us11_n697 ) , .A1( us11_n724 ) );
  AOI21_X1 us11_U311 (.ZN( us11_n498 ) , .A( us11_n724 ) , .B2( us11_n762 ) , .B1( us11_n814 ) );
  AOI21_X1 us11_U312 (.A( us11_n790 ) , .B2( us11_n791 ) , .B1( us11_n792 ) , .ZN( us11_n793 ) );
  AOI21_X1 us11_U313 (.ZN( us11_n689 ) , .B2( us11_n749 ) , .B1( us11_n763 ) , .A( us11_n806 ) );
  AOI21_X1 us11_U314 (.B1( us11_n686 ) , .ZN( us11_n687 ) , .A( us11_n728 ) , .B2( us11_n761 ) );
  AOI21_X1 us11_U315 (.ZN( us11_n569 ) , .B1( us11_n750 ) , .B2( us11_n762 ) , .A( us11_n780 ) );
  AOI21_X1 us11_U316 (.ZN( us11_n500 ) , .A( us11_n697 ) , .B1( us11_n708 ) , .B2( us11_n786 ) );
  NOR2_X1 us11_U317 (.ZN( us11_n665 ) , .A1( us11_n780 ) , .A2( us11_n813 ) );
  NOR2_X1 us11_U318 (.ZN( us11_n580 ) , .A2( us11_n697 ) , .A1( us11_n791 ) );
  AOI21_X1 us11_U319 (.ZN( us11_n571 ) , .B2( us11_n697 ) , .B1( us11_n806 ) , .A( us11_n812 ) );
  AOI221_X1 us11_U32 (.A( us11_n713 ) , .B2( us11_n714 ) , .ZN( us11_n720 ) , .C1( us11_n832 ) , .B1( us11_n839 ) , .C2( us11_n863 ) );
  NOR2_X1 us11_U320 (.ZN( us11_n684 ) , .A1( us11_n791 ) , .A2( us11_n813 ) );
  AOI21_X1 us11_U321 (.ZN( us11_n639 ) , .B2( us11_n749 ) , .A( us11_n788 ) , .B1( us11_n812 ) );
  AOI21_X1 us11_U322 (.A( us11_n733 ) , .ZN( us11_n734 ) , .B2( us11_n780 ) , .B1( us11_n792 ) );
  NAND2_X2 us11_U323 (.A1( us11_n452 ) , .A2( us11_n465 ) , .ZN( us11_n669 ) );
  NOR2_X1 us11_U324 (.ZN( us11_n711 ) , .A1( us11_n762 ) , .A2( us11_n763 ) );
  AOI21_X1 us11_U325 (.ZN( us11_n478 ) , .B2( us11_n697 ) , .A( us11_n749 ) , .B1( us11_n779 ) );
  NOR2_X1 us11_U326 (.A2( us11_n813 ) , .A1( us11_n815 ) , .ZN( us11_n821 ) );
  NOR2_X1 us11_U327 (.A1( us11_n749 ) , .ZN( us11_n767 ) , .A2( us11_n803 ) );
  NOR2_X1 us11_U328 (.ZN( us11_n682 ) , .A2( us11_n708 ) , .A1( us11_n817 ) );
  NAND2_X2 us11_U329 (.A1( us11_n451 ) , .A2( us11_n471 ) , .ZN( us11_n816 ) );
  OR2_X1 us11_U33 (.A2( us11_n711 ) , .A1( us11_n712 ) , .ZN( us11_n713 ) );
  AOI21_X1 us11_U330 (.ZN( us11_n641 ) , .B1( us11_n680 ) , .A( us11_n791 ) , .B2( us11_n817 ) );
  NAND2_X1 us11_U331 (.ZN( us11_n753 ) , .A1( us11_n763 ) , .A2( us11_n805 ) );
  OAI21_X1 us11_U332 (.A( us11_n731 ) , .B1( us11_n732 ) , .ZN( us11_n736 ) , .B2( us11_n805 ) );
  OAI21_X1 us11_U333 (.ZN( us11_n731 ) , .A( us11_n833 ) , .B2( us11_n852 ) , .B1( us11_n873 ) );
  INV_X1 us11_U334 (.A( us11_n815 ) , .ZN( us11_n855 ) );
  NAND2_X2 us11_U335 (.A1( us11_n447 ) , .A2( us11_n449 ) , .ZN( us11_n805 ) );
  NAND2_X2 us11_U336 (.A2( us11_n449 ) , .A1( us11_n452 ) , .ZN( us11_n763 ) );
  AOI21_X1 us11_U337 (.ZN( us11_n442 ) , .A( us11_n699 ) , .B1( us11_n733 ) , .B2( us11_n750 ) );
  OAI21_X1 us11_U338 (.A( us11_n698 ) , .ZN( us11_n702 ) , .B2( us11_n750 ) , .B1( us11_n804 ) );
  OAI21_X1 us11_U339 (.ZN( us11_n698 ) , .B2( us11_n833 ) , .B1( us11_n838 ) , .A( us11_n860 ) );
  NOR2_X1 us11_U34 (.ZN( us11_n680 ) , .A2( us11_n834 ) , .A1( us11_n839 ) );
  NAND2_X1 us11_U340 (.A1( us11_n699 ) , .A2( us11_n729 ) , .ZN( us11_n782 ) );
  NOR2_X1 us11_U341 (.ZN( us11_n526 ) , .A1( us11_n724 ) , .A2( us11_n750 ) );
  INV_X1 us11_U342 (.A( us11_n780 ) , .ZN( us11_n850 ) );
  NOR2_X1 us11_U343 (.ZN( us11_n518 ) , .A1( us11_n708 ) , .A2( us11_n788 ) );
  AOI21_X1 us11_U344 (.ZN( us11_n443 ) , .B1( us11_n789 ) , .B2( us11_n791 ) , .A( us11_n814 ) );
  AOI21_X1 us11_U345 (.ZN( us11_n497 ) , .A( us11_n779 ) , .B2( us11_n791 ) , .B1( us11_n804 ) );
  NAND2_X2 us11_U346 (.A2( us11_n441 ) , .A1( us11_n447 ) , .ZN( us11_n784 ) );
  NAND2_X1 us11_U347 (.ZN( us11_n714 ) , .A1( us11_n728 ) , .A2( us11_n780 ) );
  NOR2_X1 us11_U348 (.ZN( us11_n484 ) , .A1( us11_n788 ) , .A2( us11_n805 ) );
  OAI21_X1 us11_U349 (.A( us11_n787 ) , .B2( us11_n788 ) , .B1( us11_n789 ) , .ZN( us11_n795 ) );
  AOI222_X1 us11_U35 (.ZN( us11_n469 ) , .B1( us11_n832 ) , .A1( us11_n839 ) , .C1( us11_n842 ) , .C2( us11_n851 ) , .A2( us11_n855 ) , .B2( us11_n865 ) );
  NAND2_X2 us11_U350 (.A2( us11_n448 ) , .A1( us11_n452 ) , .ZN( us11_n729 ) );
  OAI21_X1 us11_U351 (.ZN( us11_n787 ) , .A( us11_n839 ) , .B1( us11_n863 ) , .B2( us11_n873 ) );
  NAND2_X1 us11_U352 (.A2( us11_n762 ) , .A1( us11_n806 ) , .ZN( us11_n810 ) );
  INV_X1 us11_U353 (.A( us11_n785 ) , .ZN( us11_n846 ) );
  NOR2_X1 us11_U354 (.ZN( us11_n470 ) , .A2( us11_n779 ) , .A1( us11_n815 ) );
  NOR2_X1 us11_U355 (.ZN( us11_n712 ) , .A2( us11_n724 ) , .A1( us11_n790 ) );
  NAND2_X1 us11_U356 (.ZN( us11_n671 ) , .A1( us11_n806 ) , .A2( us11_n816 ) );
  NAND2_X1 us11_U357 (.A2( us11_n749 ) , .A1( us11_n786 ) , .ZN( us11_n809 ) );
  INV_X1 us11_U358 (.A( us11_n724 ) , .ZN( us11_n856 ) );
  INV_X1 us11_U359 (.A( us11_n817 ) , .ZN( us11_n844 ) );
  NOR4_X1 us11_U36 (.A1( us11_n466 ) , .ZN( us11_n467 ) , .A4( us11_n542 ) , .A2( us11_n554 ) , .A3( us11_n614 ) );
  AND2_X1 us11_U360 (.ZN( us11_n732 ) , .A1( us11_n779 ) , .A2( us11_n785 ) );
  AOI221_X1 us11_U361 (.A( us11_n764 ) , .ZN( us11_n774 ) , .C2( us11_n810 ) , .B2( us11_n835 ) , .C1( us11_n855 ) , .B1( us11_n866 ) );
  AOI21_X1 us11_U362 (.B2( us11_n763 ) , .ZN( us11_n764 ) , .A( us11_n788 ) , .B1( us11_n792 ) );
  INV_X1 us11_U363 (.A( us11_n761 ) , .ZN( us11_n835 ) );
  NAND2_X1 us11_U364 (.A2( us11_n448 ) , .A1( us11_n460 ) , .ZN( us11_n728 ) );
  NAND2_X1 us11_U365 (.A1( us11_n451 ) , .A2( us11_n454 ) , .ZN( us11_n814 ) );
  NAND2_X1 us11_U366 (.A1( us11_n455 ) , .A2( us11_n462 ) , .ZN( us11_n750 ) );
  NAND2_X1 us11_U367 (.A2( us11_n454 ) , .A1( us11_n472 ) , .ZN( us11_n779 ) );
  NAND2_X1 us11_U368 (.A2( us11_n453 ) , .A1( us11_n455 ) , .ZN( us11_n806 ) );
  NAND2_X1 us11_U369 (.A1( us11_n453 ) , .A2( us11_n472 ) , .ZN( us11_n785 ) );
  AOI221_X1 us11_U37 (.ZN( us11_n468 ) , .C2( us11_n714 ) , .B2( us11_n831 ) , .C1( us11_n845 ) , .B1( us11_n860 ) , .A( us11_n864 ) );
  NAND2_X1 us11_U370 (.A2( us11_n464 ) , .A1( us11_n465 ) , .ZN( us11_n812 ) );
  NAND2_X1 us11_U371 (.A1( us11_n447 ) , .A2( us11_n448 ) , .ZN( us11_n786 ) );
  NAND2_X2 us11_U372 (.A1( us11_n455 ) , .A2( us11_n471 ) , .ZN( us11_n803 ) );
  NAND2_X1 us11_U373 (.A1( us11_n462 ) , .A2( us11_n472 ) , .ZN( us11_n788 ) );
  NOR2_X1 us11_U374 (.ZN( us11_n465 ) , .A2( us11_n847 ) , .A1( us11_n848 ) );
  NAND2_X2 us11_U375 (.A1( us11_n453 ) , .A2( us11_n461 ) , .ZN( us11_n744 ) );
  NOR2_X1 us11_U376 (.ZN( us11_n453 ) , .A1( us11_n826 ) , .A2( us11_n827 ) );
  NOR2_X1 us11_U377 (.ZN( us11_n451 ) , .A1( us11_n828 ) , .A2( us11_n829 ) );
  NAND2_X1 us11_U378 (.A2( us11_n454 ) , .A1( us11_n455 ) , .ZN( us11_n730 ) );
  NAND2_X1 us11_U379 (.A1( us11_n451 ) , .A2( us11_n462 ) , .ZN( us11_n790 ) );
  NOR4_X1 us11_U38 (.A4( us11_n514 ) , .A3( us11_n515 ) , .A2( us11_n516 ) , .A1( us11_n517 ) , .ZN( us11_n524 ) );
  NAND2_X2 us11_U380 (.A1( us11_n449 ) , .A2( us11_n460 ) , .ZN( us11_n792 ) );
  NAND2_X2 us11_U381 (.A2( us11_n448 ) , .A1( us11_n464 ) , .ZN( us11_n815 ) );
  NAND2_X2 us11_U382 (.A2( us11_n471 ) , .A1( us11_n472 ) , .ZN( us11_n817 ) );
  NAND2_X2 us11_U383 (.A1( us11_n441 ) , .A2( us11_n460 ) , .ZN( us11_n699 ) );
  NOR2_X1 us11_U384 (.ZN( us11_n447 ) , .A2( us11_n849 ) , .A1( us11_n858 ) );
  NOR2_X1 us11_U385 (.A2( sa11_6 ) , .A1( sa11_7 ) , .ZN( us11_n464 ) );
  NOR2_X1 us11_U386 (.A2( sa11_7 ) , .ZN( us11_n460 ) , .A1( us11_n849 ) );
  NOR2_X1 us11_U387 (.A2( sa11_5 ) , .ZN( us11_n448 ) , .A1( us11_n847 ) );
  NOR2_X1 us11_U388 (.A2( sa11_2 ) , .A1( sa11_3 ) , .ZN( us11_n472 ) );
  NOR2_X1 us11_U389 (.A2( sa11_0 ) , .ZN( us11_n454 ) , .A1( us11_n827 ) );
  AOI222_X1 us11_U39 (.ZN( us11_n525 ) , .A1( us11_n834 ) , .B2( us11_n837 ) , .C1( us11_n844 ) , .C2( us11_n850 ) , .A2( us11_n852 ) , .B1( us11_n866 ) );
  NOR2_X1 us11_U390 (.A2( sa11_3 ) , .ZN( us11_n455 ) , .A1( us11_n828 ) );
  NOR2_X1 us11_U391 (.A2( sa11_0 ) , .A1( sa11_1 ) , .ZN( us11_n462 ) );
  INV_X1 us11_U392 (.A( sa11_6 ) , .ZN( us11_n849 ) );
  INV_X1 us11_U393 (.A( sa11_1 ) , .ZN( us11_n827 ) );
  INV_X1 us11_U394 (.A( sa11_2 ) , .ZN( us11_n828 ) );
  INV_X1 us11_U395 (.A( sa11_5 ) , .ZN( us11_n848 ) );
  NAND2_X1 us11_U396 (.A2( us11_n461 ) , .A1( us11_n471 ) , .ZN( us11_n697 ) );
  NOR2_X1 us11_U397 (.A2( sa11_6 ) , .ZN( us11_n452 ) , .A1( us11_n858 ) );
  INV_X1 us11_U398 (.A( sa11_7 ) , .ZN( us11_n858 ) );
  NAND2_X1 us11_U399 (.A2( us11_n461 ) , .A1( us11_n462 ) , .ZN( us11_n747 ) );
  NAND2_X2 us11_U4 (.A1( us11_n441 ) , .A2( us11_n464 ) , .ZN( us11_n708 ) );
  NOR4_X1 us11_U40 (.A3( us11_n521 ) , .A1( us11_n522 ) , .ZN( us11_n523 ) , .A2( us11_n673 ) , .A4( us11_n769 ) );
  NAND2_X2 us11_U400 (.A1( us11_n454 ) , .A2( us11_n461 ) , .ZN( us11_n813 ) );
  NOR2_X1 us11_U401 (.A2( sa11_1 ) , .ZN( us11_n471 ) , .A1( us11_n826 ) );
  INV_X1 us11_U402 (.A( sa11_0 ) , .ZN( us11_n826 ) );
  OAI221_X1 us11_U403 (.A( us11_n783 ) , .C2( us11_n784 ) , .B2( us11_n785 ) , .B1( us11_n786 ) , .ZN( us11_n796 ) , .C1( us11_n813 ) );
  NAND2_X1 us11_U404 (.A1( us11_n729 ) , .A2( us11_n784 ) , .ZN( us11_n811 ) );
  OAI22_X1 us11_U405 (.ZN( us11_n588 ) , .A2( us11_n747 ) , .B2( us11_n762 ) , .A1( us11_n763 ) , .B1( us11_n784 ) );
  OAI221_X1 us11_U406 (.A( us11_n696 ) , .ZN( us11_n703 ) , .C2( us11_n784 ) , .C1( us11_n785 ) , .B1( us11_n786 ) , .B2( us11_n806 ) );
  AOI21_X1 us11_U407 (.ZN( us11_n592 ) , .B1( us11_n728 ) , .B2( us11_n784 ) , .A( us11_n790 ) );
  AOI21_X1 us11_U408 (.ZN( us11_n648 ) , .A( us11_n762 ) , .B2( us11_n784 ) , .B1( us11_n792 ) );
  AOI21_X1 us11_U409 (.ZN( us11_n623 ) , .B1( us11_n699 ) , .A( us11_n779 ) , .B2( us11_n784 ) );
  AOI221_X1 us11_U41 (.A( us11_n781 ) , .ZN( us11_n798 ) , .C2( us11_n837 ) , .B2( us11_n838 ) , .B1( us11_n865 ) , .C1( us11_n866 ) );
  OAI22_X1 us11_U410 (.ZN( us11_n681 ) , .A1( us11_n699 ) , .A2( us11_n730 ) , .B2( us11_n784 ) , .B1( us11_n817 ) );
  OAI21_X1 us11_U411 (.A( us11_n613 ) , .ZN( us11_n616 ) , .B1( us11_n625 ) , .B2( us11_n784 ) );
  NOR2_X1 us11_U412 (.ZN( us11_n610 ) , .A1( us11_n784 ) , .A2( us11_n816 ) );
  NOR2_X1 us11_U413 (.ZN( us11_n651 ) , .A1( us11_n784 ) , .A2( us11_n788 ) );
  OAI222_X1 us11_U414 (.A2( us11_n669 ) , .ZN( us11_n674 ) , .B1( us11_n747 ) , .B2( us11_n784 ) , .C2( us11_n788 ) , .C1( us11_n815 ) , .A1( us11_n817 ) );
  NOR2_X1 us11_U415 (.ZN( us11_n600 ) , .A2( us11_n697 ) , .A1( us11_n784 ) );
  NOR2_X1 us11_U416 (.ZN( us11_n553 ) , .A2( us11_n744 ) , .A1( us11_n784 ) );
  INV_X1 us11_U417 (.A( us11_n784 ) , .ZN( us11_n861 ) );
  NAND4_X1 us11_U418 (.ZN( sa10_sr_2 ) , .A4( us11_n643 ) , .A3( us11_n644 ) , .A2( us11_n645 ) , .A1( us11_n646 ) );
  AOI211_X1 us11_U419 (.A( us11_n637 ) , .ZN( us11_n645 ) , .B( us11_n743 ) , .C2( us11_n839 ) , .C1( us11_n854 ) );
  NOR4_X1 us11_U42 (.A4( us11_n793 ) , .A3( us11_n794 ) , .A2( us11_n795 ) , .A1( us11_n796 ) , .ZN( us11_n797 ) );
  NOR4_X1 us11_U420 (.A1( us11_n584 ) , .ZN( us11_n585 ) , .A3( us11_n652 ) , .A2( us11_n662 ) , .A4( us11_n767 ) );
  NOR2_X1 us11_U421 (.A2( sa11_2 ) , .ZN( us11_n461 ) , .A1( us11_n829 ) );
  INV_X1 us11_U422 (.A( sa11_3 ) , .ZN( us11_n829 ) );
  OAI222_X1 us11_U423 (.B2( us11_n747 ) , .B1( us11_n748 ) , .A2( us11_n749 ) , .ZN( us11_n757 ) , .C2( us11_n805 ) , .C1( us11_n814 ) , .A1( us11_n817 ) );
  OAI222_X1 us11_U424 (.ZN( us11_n505 ) , .C2( us11_n625 ) , .B2( us11_n647 ) , .B1( us11_n747 ) , .A2( us11_n748 ) , .C1( us11_n805 ) , .A1( us11_n806 ) );
  AOI222_X1 us11_U425 (.ZN( us11_n605 ) , .B2( us11_n671 ) , .B1( us11_n753 ) , .C2( us11_n831 ) , .A1( us11_n833 ) , .A2( us11_n862 ) , .C1( us11_n863 ) );
  AOI222_X1 us11_U426 (.ZN( us11_n513 ) , .C1( us11_n832 ) , .B2( us11_n837 ) , .A2( us11_n843 ) , .C2( us11_n862 ) , .B1( us11_n863 ) , .A1( us11_n866 ) );
  AOI221_X1 us11_U427 (.A( us11_n483 ) , .ZN( us11_n488 ) , .B1( us11_n831 ) , .C2( us11_n844 ) , .C1( us11_n852 ) , .B2( us11_n862 ) );
  NOR2_X1 us11_U428 (.ZN( us11_n789 ) , .A2( us11_n862 ) , .A1( us11_n868 ) );
  NOR2_X1 us11_U429 (.ZN( us11_n748 ) , .A1( us11_n861 ) , .A2( us11_n862 ) );
  NOR4_X1 us11_U43 (.A4( us11_n776 ) , .A3( us11_n777 ) , .A1( us11_n778 ) , .ZN( us11_n799 ) , .A2( us11_n801 ) );
  NOR2_X1 us11_U430 (.A2( sa11_4 ) , .ZN( us11_n449 ) , .A1( us11_n848 ) );
  NOR2_X1 us11_U431 (.A2( sa11_4 ) , .A1( sa11_5 ) , .ZN( us11_n441 ) );
  INV_X1 us11_U432 (.A( sa11_4 ) , .ZN( us11_n847 ) );
  AND2_X1 us11_U433 (.ZN( us11_n438 ) , .A2( us11_n831 ) , .A1( us11_n854 ) );
  AND2_X1 us11_U434 (.ZN( us11_n439 ) , .A2( us11_n843 ) , .A1( us11_n861 ) );
  NOR3_X1 us11_U435 (.A1( us11_n438 ) , .A2( us11_n439 ) , .A3( us11_n576 ) , .ZN( us11_n587 ) );
  INV_X1 us11_U436 (.A( us11_n812 ) , .ZN( us11_n854 ) );
  NAND3_X1 us11_U437 (.ZN( sa10_sr_6 ) , .A3( us11_n797 ) , .A2( us11_n798 ) , .A1( us11_n799 ) );
  NAND3_X1 us11_U438 (.ZN( sa10_sr_5 ) , .A3( us11_n758 ) , .A2( us11_n759 ) , .A1( us11_n760 ) );
  NAND3_X1 us11_U439 (.ZN( sa10_sr_4 ) , .A3( us11_n738 ) , .A2( us11_n739 ) , .A1( us11_n740 ) );
  NOR4_X1 us11_U44 (.A4( us11_n734 ) , .A3( us11_n735 ) , .A2( us11_n736 ) , .A1( us11_n737 ) , .ZN( us11_n738 ) );
  NAND3_X1 us11_U440 (.A3( us11_n675 ) , .A2( us11_n676 ) , .A1( us11_n677 ) , .ZN( us11_n807 ) );
  NAND3_X1 us11_U441 (.ZN( us11_n638 ) , .A3( us11_n708 ) , .A2( us11_n724 ) , .A1( us11_n792 ) );
  NAND3_X1 us11_U442 (.A3( us11_n618 ) , .A2( us11_n619 ) , .A1( us11_n620 ) , .ZN( us11_n725 ) );
  NAND3_X1 us11_U443 (.A3( us11_n585 ) , .A2( us11_n586 ) , .A1( us11_n587 ) , .ZN( us11_n621 ) );
  NAND3_X1 us11_U444 (.ZN( us11_n565 ) , .A3( us11_n680 ) , .A2( us11_n750 ) , .A1( us11_n785 ) );
  NAND3_X1 us11_U445 (.A3( us11_n523 ) , .A2( us11_n524 ) , .A1( us11_n525 ) , .ZN( us11_n742 ) );
  NAND3_X1 us11_U446 (.A3( us11_n512 ) , .A1( us11_n513 ) , .ZN( us11_n608 ) , .A2( us11_n871 ) );
  NAND3_X1 us11_U447 (.A3( us11_n467 ) , .A2( us11_n468 ) , .A1( us11_n469 ) , .ZN( us11_n777 ) );
  INV_X1 us11_U448 (.A( us11_n803 ) , .ZN( us11_n843 ) );
  AOI21_X1 us11_U449 (.ZN( us11_n576 ) , .B2( us11_n724 ) , .B1( us11_n748 ) , .A( us11_n785 ) );
  AOI211_X1 us11_U45 (.B( us11_n725 ) , .A( us11_n726 ) , .ZN( us11_n739 ) , .C1( us11_n843 ) , .C2( us11_n855 ) );
  NOR3_X1 us11_U46 (.A3( us11_n722 ) , .A1( us11_n723 ) , .ZN( us11_n740 ) , .A2( us11_n741 ) );
  NOR4_X1 us11_U47 (.A3( us11_n755 ) , .A2( us11_n756 ) , .A1( us11_n757 ) , .ZN( us11_n758 ) , .A4( us11_n869 ) );
  AOI211_X1 us11_U48 (.B( us11_n745 ) , .A( us11_n746 ) , .ZN( us11_n759 ) , .C1( us11_n832 ) , .C2( us11_n853 ) );
  NOR3_X1 us11_U49 (.A3( us11_n741 ) , .A2( us11_n742 ) , .A1( us11_n743 ) , .ZN( us11_n760 ) );
  NAND2_X2 us11_U5 (.A2( us11_n441 ) , .A1( us11_n452 ) , .ZN( us11_n791 ) );
  NAND4_X1 us11_U50 (.ZN( sa10_sr_3 ) , .A4( us11_n704 ) , .A3( us11_n705 ) , .A2( us11_n706 ) , .A1( us11_n707 ) );
  NOR4_X1 us11_U51 (.A4( us11_n700 ) , .A3( us11_n701 ) , .A2( us11_n702 ) , .A1( us11_n703 ) , .ZN( us11_n704 ) );
  AOI211_X1 us11_U52 (.B( us11_n694 ) , .A( us11_n695 ) , .ZN( us11_n705 ) , .C2( us11_n831 ) , .C1( us11_n851 ) );
  NOR2_X1 us11_U53 (.ZN( us11_n707 ) , .A2( us11_n776 ) , .A1( us11_n800 ) );
  NOR2_X1 us11_U54 (.ZN( us11_n804 ) , .A1( us11_n854 ) , .A2( us11_n861 ) );
  NAND4_X1 us11_U55 (.ZN( sa10_sr_1 ) , .A4( us11_n595 ) , .A3( us11_n596 ) , .A2( us11_n597 ) , .A1( us11_n598 ) );
  AOI211_X1 us11_U56 (.B( us11_n589 ) , .A( us11_n590 ) , .ZN( us11_n596 ) , .C2( us11_n811 ) , .C1( us11_n833 ) );
  NOR4_X1 us11_U57 (.A4( us11_n591 ) , .A3( us11_n592 ) , .A2( us11_n593 ) , .A1( us11_n594 ) , .ZN( us11_n595 ) );
  AOI211_X1 us11_U58 (.A( us11_n588 ) , .ZN( us11_n597 ) , .B( us11_n621 ) , .C1( us11_n845 ) , .C2( us11_n855 ) );
  NAND4_X1 us11_U59 (.ZN( sa10_sr_0 ) , .A4( us11_n501 ) , .A3( us11_n502 ) , .A2( us11_n503 ) , .A1( us11_n504 ) );
  INV_X1 us11_U6 (.A( us11_n669 ) , .ZN( us11_n865 ) );
  AOI221_X1 us11_U60 (.A( us11_n497 ) , .ZN( us11_n502 ) , .B2( us11_n843 ) , .C1( us11_n846 ) , .C2( us11_n860 ) , .B1( us11_n862 ) );
  NOR4_X1 us11_U61 (.A4( us11_n498 ) , .A3( us11_n499 ) , .A2( us11_n500 ) , .ZN( us11_n501 ) , .A1( us11_n527 ) );
  AOI211_X1 us11_U62 (.A( us11_n496 ) , .ZN( us11_n503 ) , .B( us11_n802 ) , .C2( us11_n839 ) , .C1( us11_n851 ) );
  NAND4_X1 us11_U63 (.ZN( sa10_sr_7 ) , .A4( us11_n822 ) , .A3( us11_n823 ) , .A2( us11_n824 ) , .A1( us11_n825 ) );
  AOI222_X1 us11_U64 (.C2( us11_n809 ) , .B2( us11_n810 ) , .A2( us11_n811 ) , .ZN( us11_n823 ) , .C1( us11_n832 ) , .A1( us11_n839 ) , .B1( us11_n853 ) );
  NOR4_X1 us11_U65 (.A4( us11_n818 ) , .A3( us11_n819 ) , .A2( us11_n820 ) , .A1( us11_n821 ) , .ZN( us11_n822 ) );
  AOI211_X1 us11_U66 (.B( us11_n807 ) , .A( us11_n808 ) , .ZN( us11_n824 ) , .C1( us11_n842 ) , .C2( us11_n850 ) );
  NAND4_X1 us11_U67 (.A4( us11_n603 ) , .A3( us11_n604 ) , .A2( us11_n605 ) , .A1( us11_n606 ) , .ZN( us11_n722 ) );
  NOR3_X1 us11_U68 (.A1( us11_n599 ) , .ZN( us11_n604 ) , .A3( us11_n663 ) , .A2( us11_n770 ) );
  NOR4_X1 us11_U69 (.A3( us11_n600 ) , .A2( us11_n601 ) , .A1( us11_n602 ) , .ZN( us11_n603 ) , .A4( us11_n655 ) );
  NAND2_X1 us11_U7 (.A1( us11_n449 ) , .A2( us11_n464 ) , .ZN( us11_n724 ) );
  AOI222_X1 us11_U70 (.ZN( us11_n606 ) , .A1( us11_n830 ) , .C2( us11_n837 ) , .B1( us11_n842 ) , .A2( us11_n856 ) , .B2( us11_n861 ) , .C1( us11_n868 ) );
  NAND4_X1 us11_U71 (.A4( us11_n485 ) , .A3( us11_n486 ) , .A2( us11_n487 ) , .A1( us11_n488 ) , .ZN( us11_n778 ) );
  NOR4_X1 us11_U72 (.A4( us11_n484 ) , .ZN( us11_n487 ) , .A1( us11_n566 ) , .A2( us11_n581 ) , .A3( us11_n602 ) );
  NOR4_X1 us11_U73 (.ZN( us11_n486 ) , .A1( us11_n507 ) , .A2( us11_n519 ) , .A4( us11_n546 ) , .A3( us11_n611 ) );
  NAND4_X1 us11_U74 (.A4( us11_n657 ) , .A3( us11_n658 ) , .A2( us11_n659 ) , .A1( us11_n660 ) , .ZN( us11_n800 ) );
  NOR3_X1 us11_U75 (.A3( us11_n654 ) , .A2( us11_n655 ) , .A1( us11_n656 ) , .ZN( us11_n657 ) );
  NOR3_X1 us11_U76 (.A3( us11_n651 ) , .A2( us11_n652 ) , .A1( us11_n653 ) , .ZN( us11_n658 ) );
  NOR3_X1 us11_U77 (.A3( us11_n648 ) , .A2( us11_n649 ) , .A1( us11_n650 ) , .ZN( us11_n659 ) );
  NAND4_X1 us11_U78 (.A4( us11_n560 ) , .A3( us11_n561 ) , .A2( us11_n562 ) , .A1( us11_n563 ) , .ZN( us11_n607 ) );
  NOR4_X1 us11_U79 (.ZN( us11_n561 ) , .A1( us11_n653 ) , .A3( us11_n661 ) , .A4( us11_n685 ) , .A2( us11_n768 ) );
  NOR3_X1 us11_U8 (.ZN( us11_n598 ) , .A1( us11_n608 ) , .A3( us11_n723 ) , .A2( us11_n742 ) );
  NOR4_X1 us11_U80 (.A4( us11_n552 ) , .A3( us11_n553 ) , .A2( us11_n554 ) , .A1( us11_n555 ) , .ZN( us11_n562 ) );
  NOR4_X1 us11_U81 (.A4( us11_n556 ) , .A3( us11_n557 ) , .A2( us11_n558 ) , .A1( us11_n559 ) , .ZN( us11_n560 ) );
  NAND4_X1 us11_U82 (.A4( us11_n772 ) , .A3( us11_n773 ) , .A2( us11_n774 ) , .A1( us11_n775 ) , .ZN( us11_n801 ) );
  NOR3_X1 us11_U83 (.A3( us11_n765 ) , .A2( us11_n766 ) , .A1( us11_n767 ) , .ZN( us11_n773 ) );
  NOR4_X1 us11_U84 (.A4( us11_n768 ) , .A3( us11_n769 ) , .A2( us11_n770 ) , .A1( us11_n771 ) , .ZN( us11_n772 ) );
  AOI222_X1 us11_U85 (.ZN( us11_n775 ) , .A1( us11_n830 ) , .C1( us11_n834 ) , .B2( us11_n841 ) , .A2( us11_n850 ) , .B1( us11_n861 ) , .C2( us11_n873 ) );
  NOR4_X1 us11_U86 (.A4( us11_n509 ) , .A2( us11_n510 ) , .A1( us11_n511 ) , .ZN( us11_n512 ) , .A3( us11_n670 ) );
  INV_X1 us11_U87 (.A( us11_n505 ) , .ZN( us11_n871 ) );
  NOR4_X1 us11_U88 (.A4( us11_n665 ) , .A3( us11_n666 ) , .A2( us11_n667 ) , .A1( us11_n668 ) , .ZN( us11_n676 ) );
  NOR4_X1 us11_U89 (.A4( us11_n661 ) , .A3( us11_n662 ) , .A2( us11_n663 ) , .A1( us11_n664 ) , .ZN( us11_n677 ) );
  NOR3_X1 us11_U9 (.A3( us11_n800 ) , .A2( us11_n801 ) , .A1( us11_n802 ) , .ZN( us11_n825 ) );
  NOR4_X1 us11_U90 (.A3( us11_n673 ) , .A1( us11_n674 ) , .ZN( us11_n675 ) , .A4( us11_n715 ) , .A2( us11_n859 ) );
  NOR2_X1 us11_U91 (.ZN( us11_n625 ) , .A2( us11_n836 ) , .A1( us11_n839 ) );
  NOR2_X1 us11_U92 (.ZN( us11_n761 ) , .A1( us11_n833 ) , .A2( us11_n834 ) );
  NAND4_X1 us11_U93 (.A4( us11_n456 ) , .A3( us11_n457 ) , .A2( us11_n458 ) , .A1( us11_n459 ) , .ZN( us11_n679 ) );
  AOI221_X1 us11_U94 (.A( us11_n450 ) , .ZN( us11_n459 ) , .C2( us11_n753 ) , .B1( us11_n832 ) , .C1( us11_n842 ) , .B2( us11_n861 ) );
  NOR3_X1 us11_U95 (.ZN( us11_n457 ) , .A3( us11_n530 ) , .A1( us11_n555 ) , .A2( us11_n570 ) );
  NOR4_X1 us11_U96 (.ZN( us11_n458 ) , .A2( us11_n509 ) , .A1( us11_n599 ) , .A4( us11_n628 ) , .A3( us11_n711 ) );
  NAND4_X1 us11_U97 (.A4( us11_n535 ) , .A3( us11_n536 ) , .A2( us11_n537 ) , .A1( us11_n538 ) , .ZN( us11_n622 ) );
  NOR4_X1 us11_U98 (.A1( us11_n531 ) , .ZN( us11_n536 ) , .A2( us11_n654 ) , .A4( us11_n668 ) , .A3( us11_n765 ) );
  NOR4_X1 us11_U99 (.A4( us11_n526 ) , .A2( us11_n527 ) , .A1( us11_n528 ) , .ZN( us11_n538 ) , .A3( us11_n701 ) );
  NOR3_X1 us13_U10 (.A3( us13_n621 ) , .A2( us13_n622 ) , .ZN( us13_n636 ) , .A1( us13_n725 ) );
  NOR4_X1 us13_U100 (.ZN( us13_n458 ) , .A2( us13_n509 ) , .A1( us13_n599 ) , .A4( us13_n628 ) , .A3( us13_n711 ) );
  NAND4_X1 us13_U101 (.A4( us13_n535 ) , .A3( us13_n536 ) , .A2( us13_n537 ) , .A1( us13_n538 ) , .ZN( us13_n622 ) );
  NOR4_X1 us13_U102 (.A4( us13_n526 ) , .A2( us13_n527 ) , .A1( us13_n528 ) , .ZN( us13_n538 ) , .A3( us13_n701 ) );
  NOR4_X1 us13_U103 (.A4( us13_n529 ) , .A3( us13_n530 ) , .ZN( us13_n537 ) , .A2( us13_n684 ) , .A1( us13_n794 ) );
  NOR4_X1 us13_U104 (.A4( us13_n532 ) , .A3( us13_n533 ) , .A2( us13_n534 ) , .ZN( us13_n535 ) , .A1( us13_n820 ) );
  NAND4_X1 us13_U105 (.A4( us13_n548 ) , .A3( us13_n549 ) , .A2( us13_n550 ) , .A1( us13_n551 ) , .ZN( us13_n745 ) );
  NOR3_X1 us13_U106 (.ZN( us13_n549 ) , .A2( us13_n651 ) , .A1( us13_n667 ) , .A3( us13_n771 ) );
  AOI211_X1 us13_U107 (.B( us13_n539 ) , .A( us13_n540 ) , .ZN( us13_n551 ) , .C2( us13_n839 ) , .C1( us13_n851 ) );
  NOR4_X1 us13_U108 (.A4( us13_n541 ) , .A3( us13_n542 ) , .A2( us13_n543 ) , .ZN( us13_n550 ) , .A1( us13_n688 ) );
  NAND4_X1 us13_U109 (.A4( us13_n479 ) , .A3( us13_n480 ) , .A2( us13_n481 ) , .A1( us13_n482 ) , .ZN( us13_n694 ) );
  NOR2_X1 us13_U11 (.A1( us13_n678 ) , .ZN( us13_n693 ) , .A2( us13_n807 ) );
  NOR3_X1 us13_U110 (.ZN( us13_n480 ) , .A2( us13_n508 ) , .A3( us13_n601 ) , .A1( us13_n610 ) );
  AOI211_X1 us13_U111 (.B( us13_n477 ) , .A( us13_n478 ) , .ZN( us13_n482 ) , .C2( us13_n833 ) , .C1( us13_n861 ) );
  NOR4_X1 us13_U112 (.ZN( us13_n481 ) , .A3( us13_n532 ) , .A4( us13_n545 ) , .A2( us13_n567 ) , .A1( us13_n717 ) );
  NOR2_X1 us13_U113 (.ZN( us13_n647 ) , .A1( us13_n854 ) , .A2( us13_n868 ) );
  NOR4_X1 us13_U114 (.ZN( us13_n620 ) , .A1( us13_n656 ) , .A3( us13_n666 ) , .A4( us13_n682 ) , .A2( us13_n766 ) );
  NOR4_X1 us13_U115 (.A4( us13_n609 ) , .A3( us13_n610 ) , .A2( us13_n611 ) , .A1( us13_n612 ) , .ZN( us13_n619 ) );
  NOR4_X1 us13_U116 (.A4( us13_n614 ) , .A3( us13_n615 ) , .A2( us13_n616 ) , .A1( us13_n617 ) , .ZN( us13_n618 ) );
  NOR2_X1 us13_U117 (.ZN( us13_n686 ) , .A1( us13_n831 ) , .A2( us13_n832 ) );
  NAND4_X1 us13_U118 (.A4( us13_n473 ) , .A3( us13_n474 ) , .A2( us13_n475 ) , .A1( us13_n476 ) , .ZN( us13_n678 ) );
  NOR4_X1 us13_U119 (.ZN( us13_n475 ) , .A1( us13_n531 ) , .A3( us13_n568 ) , .A4( us13_n600 ) , .A2( us13_n642 ) );
  INV_X1 us13_U12 (.A( us13_n607 ) , .ZN( us13_n874 ) );
  NOR4_X1 us13_U120 (.A4( us13_n470 ) , .ZN( us13_n476 ) , .A3( us13_n556 ) , .A1( us13_n735 ) , .A2( us13_n755 ) );
  NOR4_X1 us13_U121 (.ZN( us13_n474 ) , .A1( us13_n506 ) , .A3( us13_n544 ) , .A2( us13_n583 ) , .A4( us13_n716 ) );
  NOR2_X1 us13_U122 (.ZN( us13_n733 ) , .A2( us13_n832 ) , .A1( us13_n845 ) );
  NAND4_X1 us13_U123 (.A4( us13_n719 ) , .A3( us13_n720 ) , .A2( us13_n721 ) , .ZN( us13_n741 ) , .A1( us13_n857 ) );
  INV_X1 us13_U124 (.A( us13_n709 ) , .ZN( us13_n857 ) );
  NOR4_X1 us13_U125 (.A4( us13_n715 ) , .A3( us13_n716 ) , .A2( us13_n717 ) , .A1( us13_n718 ) , .ZN( us13_n719 ) );
  AOI221_X1 us13_U126 (.A( us13_n710 ) , .ZN( us13_n721 ) , .C2( us13_n844 ) , .B2( us13_n845 ) , .C1( us13_n861 ) , .B1( us13_n862 ) );
  NAND4_X1 us13_U127 (.A4( us13_n573 ) , .A3( us13_n574 ) , .A1( us13_n575 ) , .ZN( us13_n723 ) , .A2( us13_n874 ) );
  NOR4_X1 us13_U128 (.A4( us13_n569 ) , .A3( us13_n570 ) , .A2( us13_n571 ) , .A1( us13_n572 ) , .ZN( us13_n573 ) );
  AOI221_X1 us13_U129 (.A( us13_n564 ) , .C2( us13_n565 ) , .ZN( us13_n574 ) , .B2( us13_n845 ) , .B1( us13_n852 ) , .C1( us13_n853 ) );
  INV_X1 us13_U13 (.A( us13_n680 ) , .ZN( us13_n840 ) );
  NOR2_X1 us13_U130 (.ZN( us13_n575 ) , .A1( us13_n622 ) , .A2( us13_n745 ) );
  NAND4_X1 us13_U131 (.A4( us13_n633 ) , .A3( us13_n634 ) , .A2( us13_n635 ) , .A1( us13_n636 ) , .ZN( us13_n743 ) );
  AOI211_X1 us13_U132 (.B( us13_n623 ) , .A( us13_n624 ) , .ZN( us13_n635 ) , .C2( us13_n836 ) , .C1( us13_n863 ) );
  NOR4_X1 us13_U133 (.A4( us13_n629 ) , .A3( us13_n630 ) , .A2( us13_n631 ) , .A1( us13_n632 ) , .ZN( us13_n633 ) );
  NOR4_X1 us13_U134 (.A4( us13_n626 ) , .A3( us13_n627 ) , .A2( us13_n628 ) , .ZN( us13_n634 ) , .A1( us13_n664 ) );
  NAND4_X1 us13_U135 (.A4( us13_n493 ) , .A3( us13_n494 ) , .A1( us13_n495 ) , .ZN( us13_n802 ) , .A2( us13_n867 ) );
  AOI221_X1 us13_U136 (.A( us13_n489 ) , .ZN( us13_n494 ) , .B2( us13_n836 ) , .C2( us13_n841 ) , .C1( us13_n851 ) , .B1( us13_n860 ) );
  INV_X1 us13_U137 (.A( us13_n778 ) , .ZN( us13_n867 ) );
  NOR2_X1 us13_U138 (.ZN( us13_n495 ) , .A1( us13_n678 ) , .A2( us13_n694 ) );
  INV_X1 us13_U139 (.A( us13_n762 ) , .ZN( us13_n830 ) );
  NOR4_X1 us13_U14 (.A4( us13_n445 ) , .A3( us13_n446 ) , .A2( us13_n516 ) , .A1( us13_n541 ) , .ZN( us13_n706 ) );
  OR4_X1 us13_U140 (.A4( us13_n566 ) , .A3( us13_n567 ) , .A2( us13_n568 ) , .ZN( us13_n572 ) , .A1( us13_n665 ) );
  OR4_X1 us13_U141 (.A4( us13_n518 ) , .A2( us13_n519 ) , .A1( us13_n520 ) , .ZN( us13_n522 ) , .A3( us13_n821 ) );
  OR4_X1 us13_U142 (.ZN( us13_n466 ) , .A4( us13_n518 ) , .A3( us13_n529 ) , .A2( us13_n578 ) , .A1( us13_n712 ) );
  OR4_X1 us13_U143 (.A4( us13_n682 ) , .A3( us13_n683 ) , .A2( us13_n684 ) , .A1( us13_n685 ) , .ZN( us13_n690 ) );
  OR4_X1 us13_U144 (.A4( us13_n580 ) , .A3( us13_n581 ) , .A2( us13_n582 ) , .A1( us13_n583 ) , .ZN( us13_n584 ) );
  NAND2_X1 us13_U145 (.ZN( us13_n613 ) , .A2( us13_n837 ) , .A1( us13_n873 ) );
  OR3_X1 us13_U146 (.A3( us13_n506 ) , .A2( us13_n507 ) , .A1( us13_n508 ) , .ZN( us13_n511 ) );
  AOI221_X1 us13_U147 (.A( us13_n713 ) , .B2( us13_n714 ) , .ZN( us13_n720 ) , .C1( us13_n832 ) , .B1( us13_n839 ) , .C2( us13_n863 ) );
  OR2_X1 us13_U148 (.A2( us13_n711 ) , .A1( us13_n712 ) , .ZN( us13_n713 ) );
  INV_X1 us13_U149 (.A( us13_n463 ) , .ZN( us13_n864 ) );
  OR3_X1 us13_U15 (.ZN( us13_n446 ) , .A1( us13_n528 ) , .A3( us13_n577 ) , .A2( us13_n875 ) );
  OAI21_X1 us13_U150 (.ZN( us13_n463 ) , .B1( us13_n809 ) , .A( us13_n834 ) , .B2( us13_n851 ) );
  INV_X1 us13_U151 (.A( us13_n754 ) , .ZN( us13_n869 ) );
  OAI21_X1 us13_U152 (.B1( us13_n753 ) , .ZN( us13_n754 ) , .A( us13_n845 ) , .B2( us13_n868 ) );
  INV_X1 us13_U153 (.A( us13_n672 ) , .ZN( us13_n859 ) );
  AOI21_X1 us13_U154 (.A( us13_n670 ) , .B1( us13_n671 ) , .ZN( us13_n672 ) , .B2( us13_n856 ) );
  NAND2_X1 us13_U155 (.A1( us13_n447 ) , .A2( us13_n465 ) , .ZN( us13_n749 ) );
  OAI222_X1 us13_U156 (.B2( us13_n747 ) , .B1( us13_n748 ) , .A2( us13_n749 ) , .ZN( us13_n757 ) , .C2( us13_n805 ) , .C1( us13_n814 ) , .A1( us13_n817 ) );
  OAI222_X1 us13_U157 (.B2( us13_n708 ) , .ZN( us13_n709 ) , .C2( us13_n724 ) , .B1( us13_n747 ) , .A1( us13_n806 ) , .C1( us13_n814 ) , .A2( us13_n815 ) );
  OAI222_X1 us13_U158 (.ZN( us13_n505 ) , .C2( us13_n625 ) , .B2( us13_n647 ) , .B1( us13_n747 ) , .A2( us13_n748 ) , .C1( us13_n805 ) , .A1( us13_n806 ) );
  NOR4_X1 us13_U159 (.A2( us13_n491 ) , .A1( us13_n492 ) , .ZN( us13_n493 ) , .A3( us13_n580 ) , .A4( us13_n612 ) );
  OR4_X1 us13_U16 (.A4( us13_n442 ) , .A2( us13_n443 ) , .A1( us13_n444 ) , .ZN( us13_n445 ) , .A3( us13_n553 ) );
  OR4_X1 us13_U160 (.ZN( us13_n492 ) , .A4( us13_n534 ) , .A2( us13_n547 ) , .A1( us13_n559 ) , .A3( us13_n632 ) );
  OAI22_X1 us13_U161 (.B1( us13_n490 ) , .ZN( us13_n491 ) , .A1( us13_n686 ) , .A2( us13_n763 ) , .B2( us13_n817 ) );
  NOR3_X1 us13_U162 (.ZN( us13_n490 ) , .A1( us13_n782 ) , .A2( us13_n850 ) , .A3( us13_n863 ) );
  INV_X1 us13_U163 (.A( us13_n730 ) , .ZN( us13_n839 ) );
  INV_X1 us13_U164 (.A( us13_n790 ) , .ZN( us13_n832 ) );
  NAND2_X1 us13_U165 (.A1( us13_n451 ) , .A2( us13_n453 ) , .ZN( us13_n762 ) );
  AOI211_X1 us13_U166 (.A( us13_n637 ) , .ZN( us13_n645 ) , .B( us13_n743 ) , .C2( us13_n839 ) , .C1( us13_n854 ) );
  OAI22_X1 us13_U167 (.ZN( us13_n637 ) , .A1( us13_n699 ) , .B2( us13_n728 ) , .A2( us13_n762 ) , .B1( us13_n816 ) );
  OAI221_X1 us13_U168 (.A( us13_n727 ) , .C2( us13_n728 ) , .B2( us13_n729 ) , .B1( us13_n730 ) , .ZN( us13_n737 ) , .C1( us13_n817 ) );
  AOI22_X1 us13_U169 (.ZN( us13_n727 ) , .B1( us13_n832 ) , .A2( us13_n838 ) , .A1( us13_n863 ) , .B2( us13_n866 ) );
  INV_X1 us13_U17 (.A( us13_n613 ) , .ZN( us13_n875 ) );
  INV_X1 us13_U170 (.A( us13_n744 ) , .ZN( us13_n837 ) );
  OAI22_X1 us13_U171 (.ZN( us13_n489 ) , .A1( us13_n724 ) , .B2( us13_n728 ) , .B1( us13_n730 ) , .A2( us13_n779 ) );
  OAI22_X1 us13_U172 (.ZN( us13_n624 ) , .B1( us13_n669 ) , .B2( us13_n747 ) , .A1( us13_n815 ) , .A2( us13_n816 ) );
  OAI22_X1 us13_U173 (.B2( us13_n779 ) , .B1( us13_n780 ) , .ZN( us13_n781 ) , .A2( us13_n814 ) , .A1( us13_n815 ) );
  OAI22_X1 us13_U174 (.A1( us13_n724 ) , .ZN( us13_n726 ) , .B2( us13_n750 ) , .B1( us13_n812 ) , .A2( us13_n816 ) );
  INV_X1 us13_U175 (.A( us13_n805 ) , .ZN( us13_n860 ) );
  OAI22_X1 us13_U176 (.B2( us13_n744 ) , .ZN( us13_n746 ) , .A2( us13_n762 ) , .B1( us13_n780 ) , .A1( us13_n792 ) );
  OAI22_X1 us13_U177 (.B2( us13_n803 ) , .B1( us13_n804 ) , .A2( us13_n805 ) , .A1( us13_n806 ) , .ZN( us13_n808 ) );
  OAI22_X1 us13_U178 (.ZN( us13_n496 ) , .A2( us13_n744 ) , .A1( us13_n780 ) , .B1( us13_n791 ) , .B2( us13_n806 ) );
  OAI22_X1 us13_U179 (.ZN( us13_n710 ) , .A2( us13_n728 ) , .B2( us13_n729 ) , .A1( us13_n744 ) , .B1( us13_n813 ) );
  INV_X1 us13_U18 (.A( us13_n749 ) , .ZN( us13_n863 ) );
  INV_X1 us13_U180 (.A( us13_n788 ) , .ZN( us13_n845 ) );
  INV_X1 us13_U181 (.A( us13_n814 ) , .ZN( us13_n833 ) );
  OAI22_X1 us13_U182 (.ZN( us13_n590 ) , .B1( us13_n730 ) , .B2( us13_n749 ) , .A2( us13_n786 ) , .A1( us13_n803 ) );
  OAI22_X1 us13_U183 (.ZN( us13_n695 ) , .A2( us13_n730 ) , .A1( us13_n780 ) , .B1( us13_n791 ) , .B2( us13_n817 ) );
  INV_X1 us13_U184 (.A( us13_n816 ) , .ZN( us13_n831 ) );
  INV_X1 us13_U185 (.A( us13_n669 ) , .ZN( us13_n865 ) );
  NOR2_X1 us13_U186 (.ZN( us13_n715 ) , .A1( us13_n805 ) , .A2( us13_n817 ) );
  NOR2_X1 us13_U187 (.ZN( us13_n718 ) , .A2( us13_n724 ) , .A1( us13_n744 ) );
  NOR2_X1 us13_U188 (.ZN( us13_n666 ) , .A1( us13_n728 ) , .A2( us13_n803 ) );
  NOR2_X1 us13_U189 (.ZN( us13_n546 ) , .A2( us13_n780 ) , .A1( us13_n814 ) );
  AOI222_X1 us13_U19 (.ZN( us13_n563 ) , .B1( us13_n830 ) , .C1( us13_n841 ) , .A2( us13_n843 ) , .A1( us13_n854 ) , .B2( us13_n863 ) , .C2( us13_n873 ) );
  NOR2_X1 us13_U190 (.ZN( us13_n577 ) , .A2( us13_n699 ) , .A1( us13_n814 ) );
  NOR2_X1 us13_U191 (.ZN( us13_n570 ) , .A1( us13_n728 ) , .A2( us13_n806 ) );
  NOR2_X1 us13_U192 (.A2( us13_n744 ) , .ZN( us13_n755 ) , .A1( us13_n805 ) );
  INV_X1 us13_U193 (.A( us13_n750 ) , .ZN( us13_n842 ) );
  NOR2_X1 us13_U194 (.ZN( us13_n735 ) , .A2( us13_n803 ) , .A1( us13_n805 ) );
  NOR2_X1 us13_U195 (.ZN( us13_n532 ) , .A2( us13_n749 ) , .A1( us13_n750 ) );
  NOR2_X1 us13_U196 (.ZN( us13_n654 ) , .A1( us13_n728 ) , .A2( us13_n813 ) );
  OAI22_X1 us13_U197 (.ZN( us13_n483 ) , .A1( us13_n708 ) , .B2( us13_n785 ) , .A2( us13_n806 ) , .B1( us13_n812 ) );
  NOR2_X1 us13_U198 (.ZN( us13_n629 ) , .A2( us13_n728 ) , .A1( us13_n785 ) );
  NOR2_X1 us13_U199 (.ZN( us13_n615 ) , .A1( us13_n785 ) , .A2( us13_n815 ) );
  AOI222_X1 us13_U20 (.ZN( us13_n660 ) , .A2( us13_n839 ) , .B1( us13_n841 ) , .C2( us13_n845 ) , .A1( us13_n860 ) , .C1( us13_n863 ) , .B2( us13_n870 ) );
  NOR2_X1 us13_U200 (.ZN( us13_n612 ) , .A1( us13_n779 ) , .A2( us13_n786 ) );
  NOR2_X1 us13_U201 (.ZN( us13_n628 ) , .A2( us13_n669 ) , .A1( us13_n785 ) );
  NOR2_X1 us13_U202 (.ZN( us13_n611 ) , .A2( us13_n780 ) , .A1( us13_n806 ) );
  NOR2_X1 us13_U203 (.ZN( us13_n601 ) , .A2( us13_n780 ) , .A1( us13_n803 ) );
  INV_X1 us13_U204 (.A( us13_n747 ) , .ZN( us13_n834 ) );
  NOR2_X1 us13_U205 (.ZN( us13_n528 ) , .A2( us13_n724 ) , .A1( us13_n803 ) );
  NOR2_X1 us13_U206 (.ZN( us13_n531 ) , .A2( us13_n780 ) , .A1( us13_n816 ) );
  NOR2_X1 us13_U207 (.A2( us13_n708 ) , .A1( us13_n750 ) , .ZN( us13_n771 ) );
  NOR2_X1 us13_U208 (.ZN( us13_n599 ) , .A2( us13_n791 ) , .A1( us13_n816 ) );
  NOR2_X1 us13_U209 (.ZN( us13_n652 ) , .A1( us13_n669 ) , .A2( us13_n814 ) );
  INV_X1 us13_U21 (.A( us13_n647 ) , .ZN( us13_n870 ) );
  INV_X1 us13_U210 (.A( us13_n792 ) , .ZN( us13_n851 ) );
  NOR2_X1 us13_U211 (.A1( us13_n669 ) , .ZN( us13_n673 ) , .A2( us13_n744 ) );
  NOR2_X1 us13_U212 (.ZN( us13_n602 ) , .A1( us13_n669 ) , .A2( us13_n803 ) );
  NOR2_X1 us13_U213 (.A1( us13_n669 ) , .ZN( us13_n688 ) , .A2( us13_n816 ) );
  NOR2_X1 us13_U214 (.ZN( us13_n667 ) , .A1( us13_n750 ) , .A2( us13_n815 ) );
  NOR2_X1 us13_U215 (.A2( us13_n744 ) , .ZN( us13_n769 ) , .A1( us13_n812 ) );
  NOR2_X1 us13_U216 (.ZN( us13_n555 ) , .A1( us13_n750 ) , .A2( us13_n791 ) );
  NOR2_X1 us13_U217 (.ZN( us13_n508 ) , .A2( us13_n780 ) , .A1( us13_n785 ) );
  NOR2_X1 us13_U218 (.ZN( us13_n543 ) , .A2( us13_n708 ) , .A1( us13_n785 ) );
  NOR2_X1 us13_U219 (.ZN( us13_n664 ) , .A1( us13_n785 ) , .A2( us13_n791 ) );
  NOR4_X1 us13_U22 (.ZN( us13_n473 ) , .A2( us13_n521 ) , .A4( us13_n594 ) , .A1( us13_n609 ) , .A3( us13_n629 ) );
  NOR2_X1 us13_U220 (.A1( us13_n669 ) , .ZN( us13_n766 ) , .A2( us13_n813 ) );
  NOR2_X1 us13_U221 (.A1( us13_n699 ) , .ZN( us13_n768 ) , .A2( us13_n813 ) );
  NOR2_X1 us13_U222 (.ZN( us13_n527 ) , .A1( us13_n669 ) , .A2( us13_n779 ) );
  NOR2_X1 us13_U223 (.ZN( us13_n557 ) , .A1( us13_n792 ) , .A2( us13_n814 ) );
  NOR2_X1 us13_U224 (.ZN( us13_n545 ) , .A1( us13_n749 ) , .A2( us13_n814 ) );
  NOR2_X1 us13_U225 (.ZN( us13_n556 ) , .A1( us13_n762 ) , .A2( us13_n805 ) );
  NOR2_X1 us13_U226 (.ZN( us13_n661 ) , .A1( us13_n729 ) , .A2( us13_n790 ) );
  NOR2_X1 us13_U227 (.ZN( us13_n507 ) , .A1( us13_n812 ) , .A2( us13_n817 ) );
  INV_X1 us13_U228 (.A( us13_n806 ) , .ZN( us13_n841 ) );
  NOR2_X1 us13_U229 (.ZN( us13_n554 ) , .A1( us13_n786 ) , .A2( us13_n813 ) );
  NOR4_X1 us13_U23 (.A4( us13_n544 ) , .A3( us13_n545 ) , .A2( us13_n546 ) , .A1( us13_n547 ) , .ZN( us13_n548 ) );
  NOR2_X1 us13_U230 (.ZN( us13_n509 ) , .A1( us13_n729 ) , .A2( us13_n779 ) );
  NOR2_X1 us13_U231 (.ZN( us13_n530 ) , .A2( us13_n744 ) , .A1( us13_n792 ) );
  OAI22_X1 us13_U232 (.B2( us13_n750 ) , .B1( us13_n751 ) , .A1( us13_n752 ) , .ZN( us13_n756 ) , .A2( us13_n806 ) );
  NOR2_X1 us13_U233 (.ZN( us13_n751 ) , .A2( us13_n852 ) , .A1( us13_n860 ) );
  NOR3_X1 us13_U234 (.ZN( us13_n752 ) , .A2( us13_n853 ) , .A1( us13_n863 ) , .A3( us13_n865 ) );
  NOR2_X1 us13_U235 (.ZN( us13_n544 ) , .A2( us13_n785 ) , .A1( us13_n792 ) );
  NOR2_X1 us13_U236 (.A1( us13_n749 ) , .ZN( us13_n767 ) , .A2( us13_n803 ) );
  NOR2_X1 us13_U237 (.ZN( us13_n516 ) , .A1( us13_n708 ) , .A2( us13_n744 ) );
  NOR2_X1 us13_U238 (.ZN( us13_n663 ) , .A1( us13_n729 ) , .A2( us13_n785 ) );
  OAI22_X1 us13_U239 (.B1( us13_n440 ) , .ZN( us13_n444 ) , .A2( us13_n728 ) , .A1( us13_n744 ) , .B2( us13_n749 ) );
  NOR4_X1 us13_U24 (.ZN( us13_n479 ) , .A1( us13_n520 ) , .A4( us13_n557 ) , .A3( us13_n582 ) , .A2( us13_n630 ) );
  NOR3_X1 us13_U240 (.ZN( us13_n440 ) , .A2( us13_n836 ) , .A3( us13_n837 ) , .A1( us13_n846 ) );
  NOR2_X1 us13_U241 (.ZN( us13_n717 ) , .A2( us13_n744 ) , .A1( us13_n786 ) );
  INV_X1 us13_U242 (.A( us13_n728 ) , .ZN( us13_n852 ) );
  NOR2_X1 us13_U243 (.ZN( us13_n506 ) , .A2( us13_n728 ) , .A1( us13_n762 ) );
  NOR2_X1 us13_U244 (.ZN( us13_n614 ) , .A1( us13_n762 ) , .A2( us13_n812 ) );
  NOR2_X1 us13_U245 (.ZN( us13_n517 ) , .A1( us13_n708 ) , .A2( us13_n803 ) );
  NOR2_X1 us13_U246 (.ZN( us13_n558 ) , .A1( us13_n708 ) , .A2( us13_n816 ) );
  AOI21_X1 us13_U247 (.A( us13_n812 ) , .B2( us13_n813 ) , .B1( us13_n814 ) , .ZN( us13_n819 ) );
  NOR2_X1 us13_U248 (.ZN( us13_n670 ) , .A1( us13_n790 ) , .A2( us13_n805 ) );
  NOR2_X1 us13_U249 (.ZN( us13_n630 ) , .A1( us13_n747 ) , .A2( us13_n815 ) );
  NOR4_X1 us13_U25 (.ZN( us13_n456 ) , .A2( us13_n517 ) , .A1( us13_n543 ) , .A3( us13_n579 ) , .A4( us13_n615 ) );
  NOR2_X1 us13_U250 (.ZN( us13_n655 ) , .A1( us13_n790 ) , .A2( us13_n815 ) );
  NOR2_X1 us13_U251 (.ZN( us13_n521 ) , .A1( us13_n790 ) , .A2( us13_n812 ) );
  NOR2_X1 us13_U252 (.ZN( us13_n668 ) , .A2( us13_n708 ) , .A1( us13_n790 ) );
  NOR2_X1 us13_U253 (.ZN( us13_n542 ) , .A1( us13_n762 ) , .A2( us13_n791 ) );
  NOR2_X1 us13_U254 (.ZN( us13_n701 ) , .A2( us13_n786 ) , .A1( us13_n817 ) );
  NOR2_X1 us13_U255 (.ZN( us13_n631 ) , .A1( us13_n724 ) , .A2( us13_n813 ) );
  NOR2_X1 us13_U256 (.ZN( us13_n656 ) , .A1( us13_n747 ) , .A2( us13_n780 ) );
  INV_X1 us13_U257 (.A( us13_n763 ) , .ZN( us13_n866 ) );
  NOR2_X1 us13_U258 (.ZN( us13_n609 ) , .A2( us13_n724 ) , .A1( us13_n817 ) );
  NOR2_X1 us13_U259 (.A1( us13_n730 ) , .ZN( us13_n765 ) , .A2( us13_n786 ) );
  NOR4_X1 us13_U26 (.ZN( us13_n485 ) , .A2( us13_n533 ) , .A1( us13_n558 ) , .A3( us13_n631 ) , .A4( us13_n718 ) );
  NOR2_X1 us13_U260 (.ZN( us13_n533 ) , .A2( us13_n724 ) , .A1( us13_n730 ) );
  NOR2_X1 us13_U261 (.ZN( us13_n579 ) , .A2( us13_n708 ) , .A1( us13_n730 ) );
  AOI21_X1 us13_U262 (.B1( us13_n625 ) , .ZN( us13_n627 ) , .A( us13_n763 ) , .B2( us13_n814 ) );
  AOI21_X1 us13_U263 (.A( us13_n815 ) , .B2( us13_n816 ) , .B1( us13_n817 ) , .ZN( us13_n818 ) );
  NOR2_X1 us13_U264 (.ZN( us13_n582 ) , .A1( us13_n744 ) , .A2( us13_n815 ) );
  NOR2_X1 us13_U265 (.A2( us13_n708 ) , .A1( us13_n762 ) , .ZN( us13_n794 ) );
  AOI21_X1 us13_U266 (.ZN( us13_n515 ) , .A( us13_n729 ) , .B1( us13_n750 ) , .B2( us13_n803 ) );
  NOR2_X1 us13_U267 (.ZN( us13_n642 ) , .A2( us13_n788 ) , .A1( us13_n791 ) );
  AOI21_X1 us13_U268 (.ZN( us13_n499 ) , .B1( us13_n680 ) , .A( us13_n812 ) , .B2( us13_n816 ) );
  AOI21_X1 us13_U269 (.ZN( us13_n650 ) , .A( us13_n779 ) , .B1( us13_n792 ) , .B2( us13_n805 ) );
  NOR4_X1 us13_U27 (.A1( us13_n531 ) , .ZN( us13_n536 ) , .A2( us13_n654 ) , .A4( us13_n668 ) , .A3( us13_n765 ) );
  NOR2_X1 us13_U270 (.ZN( us13_n520 ) , .A2( us13_n708 ) , .A1( us13_n814 ) );
  AOI21_X1 us13_U271 (.ZN( us13_n626 ) , .B2( us13_n669 ) , .A( us13_n790 ) , .B1( us13_n791 ) );
  NOR2_X1 us13_U272 (.ZN( us13_n653 ) , .A1( us13_n762 ) , .A2( us13_n786 ) );
  AOI21_X1 us13_U273 (.ZN( us13_n477 ) , .A( us13_n669 ) , .B1( us13_n750 ) , .B2( us13_n806 ) );
  NOR2_X1 us13_U274 (.ZN( us13_n559 ) , .A2( us13_n791 ) , .A1( us13_n803 ) );
  NOR2_X1 us13_U275 (.ZN( us13_n519 ) , .A2( us13_n699 ) , .A1( us13_n816 ) );
  NOR2_X1 us13_U276 (.ZN( us13_n683 ) , .A2( us13_n699 ) , .A1( us13_n803 ) );
  AOI21_X1 us13_U277 (.ZN( us13_n510 ) , .B2( us13_n669 ) , .A( us13_n730 ) , .B1( us13_n815 ) );
  AOI21_X1 us13_U278 (.ZN( us13_n540 ) , .A( us13_n763 ) , .B2( us13_n779 ) , .B1( us13_n817 ) );
  NOR2_X1 us13_U279 (.ZN( us13_n581 ) , .A1( us13_n669 ) , .A2( us13_n788 ) );
  NOR2_X1 us13_U28 (.ZN( us13_n680 ) , .A2( us13_n834 ) , .A1( us13_n839 ) );
  AOI21_X1 us13_U280 (.ZN( us13_n589 ) , .B2( us13_n699 ) , .B1( us13_n815 ) , .A( us13_n817 ) );
  AOI21_X1 us13_U281 (.ZN( us13_n498 ) , .A( us13_n724 ) , .B2( us13_n762 ) , .B1( us13_n814 ) );
  AOI21_X1 us13_U282 (.ZN( us13_n539 ) , .B2( us13_n812 ) , .A( us13_n814 ) , .B1( us13_n815 ) );
  AOI21_X1 us13_U283 (.B1( us13_n699 ) , .ZN( us13_n700 ) , .A( us13_n732 ) , .B2( us13_n763 ) );
  AOI21_X1 us13_U284 (.ZN( us13_n591 ) , .B2( us13_n763 ) , .A( us13_n785 ) , .B1( us13_n812 ) );
  INV_X1 us13_U285 (.A( us13_n791 ) , .ZN( us13_n873 ) );
  NOR2_X1 us13_U286 (.ZN( us13_n547 ) , .A1( us13_n699 ) , .A2( us13_n744 ) );
  NOR2_X1 us13_U287 (.ZN( us13_n665 ) , .A1( us13_n780 ) , .A2( us13_n813 ) );
  INV_X1 us13_U288 (.A( us13_n729 ) , .ZN( us13_n868 ) );
  AOI21_X1 us13_U289 (.ZN( us13_n640 ) , .B2( us13_n747 ) , .A( us13_n792 ) , .B1( us13_n803 ) );
  AOI221_X1 us13_U29 (.A( us13_n781 ) , .ZN( us13_n798 ) , .C2( us13_n837 ) , .B2( us13_n838 ) , .B1( us13_n865 ) , .C1( us13_n866 ) );
  AOI21_X1 us13_U290 (.ZN( us13_n569 ) , .B1( us13_n750 ) , .B2( us13_n762 ) , .A( us13_n780 ) );
  AOI21_X1 us13_U291 (.ZN( us13_n649 ) , .B1( us13_n729 ) , .B2( us13_n763 ) , .A( us13_n813 ) );
  NOR2_X1 us13_U292 (.ZN( us13_n685 ) , .A1( us13_n729 ) , .A2( us13_n816 ) );
  AOI21_X1 us13_U293 (.B1( us13_n686 ) , .ZN( us13_n687 ) , .A( us13_n728 ) , .B2( us13_n761 ) );
  NOR2_X1 us13_U294 (.ZN( us13_n568 ) , .A1( us13_n729 ) , .A2( us13_n762 ) );
  NOR2_X1 us13_U295 (.ZN( us13_n684 ) , .A1( us13_n791 ) , .A2( us13_n813 ) );
  AOI21_X1 us13_U296 (.ZN( us13_n514 ) , .A( us13_n779 ) , .B2( us13_n792 ) , .B1( us13_n812 ) );
  AOI21_X1 us13_U297 (.ZN( us13_n593 ) , .B1( us13_n750 ) , .A( us13_n792 ) , .B2( us13_n813 ) );
  AOI21_X1 us13_U298 (.ZN( us13_n450 ) , .B2( us13_n792 ) , .A( us13_n803 ) , .B1( us13_n815 ) );
  AOI21_X1 us13_U299 (.ZN( us13_n639 ) , .B2( us13_n749 ) , .A( us13_n788 ) , .B1( us13_n812 ) );
  NAND4_X1 us13_U3 (.ZN( sa12_sr_2 ) , .A4( us13_n643 ) , .A3( us13_n644 ) , .A2( us13_n645 ) , .A1( us13_n646 ) );
  NOR4_X1 us13_U30 (.A4( us13_n793 ) , .A3( us13_n794 ) , .A2( us13_n795 ) , .A1( us13_n796 ) , .ZN( us13_n797 ) );
  INV_X1 us13_U300 (.A( us13_n699 ) , .ZN( us13_n853 ) );
  AOI21_X1 us13_U301 (.ZN( us13_n564 ) , .B1( us13_n724 ) , .A( us13_n779 ) , .B2( us13_n791 ) );
  AOI21_X1 us13_U302 (.ZN( us13_n497 ) , .A( us13_n779 ) , .B2( us13_n791 ) , .B1( us13_n804 ) );
  NOR2_X1 us13_U303 (.ZN( us13_n529 ) , .A1( us13_n708 ) , .A2( us13_n779 ) );
  AOI21_X1 us13_U304 (.ZN( us13_n689 ) , .B2( us13_n749 ) , .B1( us13_n763 ) , .A( us13_n806 ) );
  NOR2_X1 us13_U305 (.ZN( us13_n567 ) , .A1( us13_n747 ) , .A2( us13_n805 ) );
  AOI21_X1 us13_U306 (.A( us13_n790 ) , .B2( us13_n791 ) , .B1( us13_n792 ) , .ZN( us13_n793 ) );
  AOI21_X1 us13_U307 (.A( us13_n733 ) , .ZN( us13_n734 ) , .B2( us13_n780 ) , .B1( us13_n792 ) );
  NOR2_X1 us13_U308 (.A2( us13_n813 ) , .A1( us13_n815 ) , .ZN( us13_n821 ) );
  AOI21_X1 us13_U309 (.ZN( us13_n641 ) , .B1( us13_n680 ) , .A( us13_n791 ) , .B2( us13_n817 ) );
  NOR4_X1 us13_U31 (.A4( us13_n776 ) , .A3( us13_n777 ) , .A1( us13_n778 ) , .ZN( us13_n799 ) , .A2( us13_n801 ) );
  NOR2_X1 us13_U310 (.ZN( us13_n578 ) , .A1( us13_n708 ) , .A2( us13_n813 ) );
  NOR2_X1 us13_U311 (.ZN( us13_n682 ) , .A2( us13_n708 ) , .A1( us13_n817 ) );
  NOR2_X1 us13_U312 (.ZN( us13_n711 ) , .A1( us13_n762 ) , .A2( us13_n763 ) );
  NOR2_X1 us13_U313 (.ZN( us13_n583 ) , .A1( us13_n792 ) , .A2( us13_n817 ) );
  NOR2_X1 us13_U314 (.ZN( us13_n534 ) , .A1( us13_n724 ) , .A2( us13_n788 ) );
  NAND2_X1 us13_U315 (.ZN( us13_n753 ) , .A1( us13_n763 ) , .A2( us13_n805 ) );
  INV_X1 us13_U316 (.A( us13_n815 ) , .ZN( us13_n855 ) );
  AOI21_X1 us13_U317 (.ZN( us13_n442 ) , .A( us13_n699 ) , .B1( us13_n733 ) , .B2( us13_n750 ) );
  OAI21_X1 us13_U318 (.A( us13_n731 ) , .B1( us13_n732 ) , .ZN( us13_n736 ) , .B2( us13_n805 ) );
  OAI21_X1 us13_U319 (.ZN( us13_n731 ) , .A( us13_n833 ) , .B2( us13_n852 ) , .B1( us13_n873 ) );
  NOR4_X1 us13_U32 (.A3( us13_n755 ) , .A2( us13_n756 ) , .A1( us13_n757 ) , .ZN( us13_n758 ) , .A4( us13_n869 ) );
  INV_X1 us13_U320 (.A( us13_n780 ) , .ZN( us13_n850 ) );
  INV_X1 us13_U321 (.A( us13_n785 ) , .ZN( us13_n846 ) );
  AOI22_X1 us13_U322 (.ZN( us13_n696 ) , .A1( us13_n830 ) , .B2( us13_n843 ) , .A2( us13_n865 ) , .B1( us13_n868 ) );
  AOI22_X1 us13_U323 (.A2( us13_n782 ) , .ZN( us13_n783 ) , .B2( us13_n831 ) , .A1( us13_n834 ) , .B1( us13_n863 ) );
  AOI21_X1 us13_U324 (.ZN( us13_n443 ) , .B1( us13_n789 ) , .B2( us13_n791 ) , .A( us13_n814 ) );
  NAND2_X1 us13_U325 (.ZN( us13_n714 ) , .A1( us13_n728 ) , .A2( us13_n780 ) );
  OAI21_X1 us13_U326 (.A( us13_n787 ) , .B2( us13_n788 ) , .B1( us13_n789 ) , .ZN( us13_n795 ) );
  OAI21_X1 us13_U327 (.ZN( us13_n787 ) , .A( us13_n839 ) , .B1( us13_n863 ) , .B2( us13_n873 ) );
  NAND2_X1 us13_U328 (.A2( us13_n762 ) , .A1( us13_n806 ) , .ZN( us13_n810 ) );
  NOR2_X1 us13_U329 (.ZN( us13_n484 ) , .A1( us13_n788 ) , .A2( us13_n805 ) );
  AOI211_X1 us13_U33 (.B( us13_n745 ) , .A( us13_n746 ) , .ZN( us13_n759 ) , .C1( us13_n832 ) , .C2( us13_n853 ) );
  NOR2_X1 us13_U330 (.ZN( us13_n470 ) , .A2( us13_n779 ) , .A1( us13_n815 ) );
  NOR2_X1 us13_U331 (.ZN( us13_n712 ) , .A2( us13_n724 ) , .A1( us13_n790 ) );
  NOR2_X1 us13_U332 (.ZN( us13_n526 ) , .A1( us13_n724 ) , .A2( us13_n750 ) );
  NAND2_X1 us13_U333 (.A1( us13_n699 ) , .A2( us13_n729 ) , .ZN( us13_n782 ) );
  NOR2_X1 us13_U334 (.ZN( us13_n518 ) , .A1( us13_n708 ) , .A2( us13_n788 ) );
  INV_X1 us13_U335 (.A( us13_n813 ) , .ZN( us13_n836 ) );
  NAND2_X1 us13_U336 (.ZN( us13_n671 ) , .A1( us13_n806 ) , .A2( us13_n816 ) );
  OAI21_X1 us13_U337 (.A( us13_n698 ) , .ZN( us13_n702 ) , .B2( us13_n750 ) , .B1( us13_n804 ) );
  OAI21_X1 us13_U338 (.ZN( us13_n698 ) , .B2( us13_n833 ) , .B1( us13_n838 ) , .A( us13_n860 ) );
  NAND2_X1 us13_U339 (.A2( us13_n749 ) , .A1( us13_n786 ) , .ZN( us13_n809 ) );
  NOR3_X1 us13_U34 (.A3( us13_n741 ) , .A2( us13_n742 ) , .A1( us13_n743 ) , .ZN( us13_n760 ) );
  INV_X1 us13_U340 (.A( us13_n724 ) , .ZN( us13_n856 ) );
  INV_X1 us13_U341 (.A( us13_n817 ) , .ZN( us13_n844 ) );
  NAND2_X2 us13_U342 (.A1( us13_n451 ) , .A2( us13_n462 ) , .ZN( us13_n790 ) );
  AND2_X1 us13_U343 (.ZN( us13_n732 ) , .A1( us13_n779 ) , .A2( us13_n785 ) );
  OAI222_X1 us13_U344 (.ZN( us13_n617 ) , .B1( us13_n697 ) , .C1( us13_n724 ) , .C2( us13_n747 ) , .B2( us13_n786 ) , .A2( us13_n792 ) , .A1( us13_n816 ) );
  AOI221_X1 us13_U345 (.A( us13_n764 ) , .ZN( us13_n774 ) , .C2( us13_n810 ) , .B2( us13_n835 ) , .C1( us13_n855 ) , .B1( us13_n866 ) );
  AOI21_X1 us13_U346 (.B2( us13_n763 ) , .ZN( us13_n764 ) , .A( us13_n788 ) , .B1( us13_n792 ) );
  INV_X1 us13_U347 (.A( us13_n761 ) , .ZN( us13_n835 ) );
  NAND2_X1 us13_U348 (.A1( us13_n451 ) , .A2( us13_n454 ) , .ZN( us13_n814 ) );
  NAND2_X1 us13_U349 (.A1( us13_n447 ) , .A2( us13_n449 ) , .ZN( us13_n805 ) );
  NOR4_X1 us13_U35 (.A4( us13_n734 ) , .A3( us13_n735 ) , .A2( us13_n736 ) , .A1( us13_n737 ) , .ZN( us13_n738 ) );
  NAND2_X1 us13_U350 (.A1( us13_n453 ) , .A2( us13_n461 ) , .ZN( us13_n744 ) );
  NAND2_X1 us13_U351 (.A1( us13_n455 ) , .A2( us13_n471 ) , .ZN( us13_n803 ) );
  NAND2_X1 us13_U352 (.A1( us13_n455 ) , .A2( us13_n462 ) , .ZN( us13_n750 ) );
  NAND2_X1 us13_U353 (.A1( us13_n451 ) , .A2( us13_n471 ) , .ZN( us13_n816 ) );
  NAND2_X1 us13_U354 (.A1( us13_n452 ) , .A2( us13_n465 ) , .ZN( us13_n669 ) );
  NAND2_X1 us13_U355 (.A2( us13_n448 ) , .A1( us13_n460 ) , .ZN( us13_n728 ) );
  NAND2_X1 us13_U356 (.A2( us13_n453 ) , .A1( us13_n455 ) , .ZN( us13_n806 ) );
  NAND2_X1 us13_U357 (.A1( us13_n453 ) , .A2( us13_n472 ) , .ZN( us13_n785 ) );
  NAND2_X1 us13_U358 (.A2( us13_n454 ) , .A1( us13_n472 ) , .ZN( us13_n779 ) );
  NAND2_X1 us13_U359 (.A2( us13_n464 ) , .A1( us13_n465 ) , .ZN( us13_n812 ) );
  AOI211_X1 us13_U36 (.B( us13_n725 ) , .A( us13_n726 ) , .ZN( us13_n739 ) , .C1( us13_n843 ) , .C2( us13_n855 ) );
  NAND2_X1 us13_U360 (.A1( us13_n441 ) , .A2( us13_n460 ) , .ZN( us13_n699 ) );
  NAND2_X1 us13_U361 (.A2( us13_n449 ) , .A1( us13_n452 ) , .ZN( us13_n763 ) );
  NAND2_X1 us13_U362 (.A2( us13_n448 ) , .A1( us13_n452 ) , .ZN( us13_n729 ) );
  NAND2_X1 us13_U363 (.A1( us13_n447 ) , .A2( us13_n448 ) , .ZN( us13_n786 ) );
  NAND2_X1 us13_U364 (.A2( us13_n461 ) , .A1( us13_n462 ) , .ZN( us13_n747 ) );
  NAND2_X1 us13_U365 (.A1( us13_n462 ) , .A2( us13_n472 ) , .ZN( us13_n788 ) );
  NOR2_X1 us13_U366 (.ZN( us13_n465 ) , .A2( us13_n847 ) , .A1( us13_n848 ) );
  NOR2_X1 us13_U367 (.ZN( us13_n453 ) , .A1( us13_n826 ) , .A2( us13_n827 ) );
  NOR2_X1 us13_U368 (.ZN( us13_n451 ) , .A1( us13_n828 ) , .A2( us13_n829 ) );
  NAND2_X1 us13_U369 (.A2( us13_n461 ) , .A1( us13_n471 ) , .ZN( us13_n697 ) );
  NOR3_X1 us13_U37 (.A3( us13_n722 ) , .A1( us13_n723 ) , .ZN( us13_n740 ) , .A2( us13_n741 ) );
  NAND2_X1 us13_U370 (.A2( us13_n454 ) , .A1( us13_n455 ) , .ZN( us13_n730 ) );
  NAND2_X1 us13_U371 (.A2( us13_n441 ) , .A1( us13_n447 ) , .ZN( us13_n784 ) );
  NAND2_X2 us13_U372 (.A2( us13_n448 ) , .A1( us13_n464 ) , .ZN( us13_n815 ) );
  NAND2_X2 us13_U373 (.A2( us13_n441 ) , .A1( us13_n452 ) , .ZN( us13_n791 ) );
  NAND2_X2 us13_U374 (.A1( us13_n449 ) , .A2( us13_n460 ) , .ZN( us13_n792 ) );
  NAND2_X2 us13_U375 (.A1( us13_n441 ) , .A2( us13_n464 ) , .ZN( us13_n708 ) );
  NAND2_X2 us13_U376 (.A2( us13_n460 ) , .A1( us13_n465 ) , .ZN( us13_n780 ) );
  NOR2_X1 us13_U377 (.ZN( us13_n447 ) , .A2( us13_n849 ) , .A1( us13_n858 ) );
  NOR2_X1 us13_U378 (.A2( sa13_6 ) , .A1( sa13_7 ) , .ZN( us13_n464 ) );
  NOR2_X1 us13_U379 (.A2( sa13_7 ) , .ZN( us13_n460 ) , .A1( us13_n849 ) );
  NAND4_X1 us13_U38 (.ZN( sa12_sr_3 ) , .A4( us13_n704 ) , .A3( us13_n705 ) , .A2( us13_n706 ) , .A1( us13_n707 ) );
  NOR2_X1 us13_U380 (.A2( sa13_4 ) , .ZN( us13_n449 ) , .A1( us13_n848 ) );
  NOR2_X1 us13_U381 (.A2( sa13_4 ) , .A1( sa13_5 ) , .ZN( us13_n441 ) );
  NOR2_X1 us13_U382 (.A2( sa13_5 ) , .ZN( us13_n448 ) , .A1( us13_n847 ) );
  NOR2_X1 us13_U383 (.A2( sa13_1 ) , .ZN( us13_n471 ) , .A1( us13_n826 ) );
  NOR2_X1 us13_U384 (.A2( sa13_2 ) , .A1( sa13_3 ) , .ZN( us13_n472 ) );
  NOR2_X1 us13_U385 (.A2( sa13_6 ) , .ZN( us13_n452 ) , .A1( us13_n858 ) );
  NOR2_X1 us13_U386 (.A2( sa13_0 ) , .A1( sa13_1 ) , .ZN( us13_n462 ) );
  NOR2_X1 us13_U387 (.A2( sa13_3 ) , .ZN( us13_n455 ) , .A1( us13_n828 ) );
  NOR2_X1 us13_U388 (.A2( sa13_2 ) , .ZN( us13_n461 ) , .A1( us13_n829 ) );
  NOR2_X1 us13_U389 (.A2( sa13_0 ) , .ZN( us13_n454 ) , .A1( us13_n827 ) );
  NOR4_X1 us13_U39 (.A4( us13_n700 ) , .A3( us13_n701 ) , .A2( us13_n702 ) , .A1( us13_n703 ) , .ZN( us13_n704 ) );
  INV_X1 us13_U390 (.A( sa13_4 ) , .ZN( us13_n847 ) );
  INV_X1 us13_U391 (.A( sa13_6 ) , .ZN( us13_n849 ) );
  INV_X1 us13_U392 (.A( sa13_1 ) , .ZN( us13_n827 ) );
  INV_X1 us13_U393 (.A( sa13_3 ) , .ZN( us13_n829 ) );
  INV_X1 us13_U394 (.A( sa13_0 ) , .ZN( us13_n826 ) );
  INV_X1 us13_U395 (.A( sa13_2 ) , .ZN( us13_n828 ) );
  INV_X1 us13_U396 (.A( sa13_7 ) , .ZN( us13_n858 ) );
  INV_X1 us13_U397 (.A( sa13_5 ) , .ZN( us13_n848 ) );
  AOI21_X1 us13_U398 (.ZN( us13_n500 ) , .A( us13_n697 ) , .B1( us13_n708 ) , .B2( us13_n786 ) );
  INV_X1 us13_U399 (.A( us13_n697 ) , .ZN( us13_n838 ) );
  NAND2_X1 us13_U4 (.A1( us13_n449 ) , .A2( us13_n464 ) , .ZN( us13_n724 ) );
  AOI211_X1 us13_U40 (.B( us13_n694 ) , .A( us13_n695 ) , .ZN( us13_n705 ) , .C2( us13_n831 ) , .C1( us13_n851 ) );
  AOI21_X1 us13_U400 (.ZN( us13_n571 ) , .B2( us13_n697 ) , .B1( us13_n806 ) , .A( us13_n812 ) );
  NOR2_X1 us13_U401 (.A1( us13_n697 ) , .ZN( us13_n770 ) , .A2( us13_n815 ) );
  NOR2_X1 us13_U402 (.ZN( us13_n566 ) , .A2( us13_n697 ) , .A1( us13_n763 ) );
  AOI21_X1 us13_U403 (.ZN( us13_n552 ) , .B1( us13_n669 ) , .A( us13_n697 ) , .B2( us13_n805 ) );
  NOR2_X1 us13_U404 (.ZN( us13_n632 ) , .A2( us13_n697 ) , .A1( us13_n724 ) );
  NOR2_X1 us13_U405 (.ZN( us13_n541 ) , .A2( us13_n697 ) , .A1( us13_n699 ) );
  AOI21_X1 us13_U406 (.ZN( us13_n478 ) , .B2( us13_n697 ) , .A( us13_n749 ) , .B1( us13_n779 ) );
  NOR2_X1 us13_U407 (.A2( us13_n697 ) , .A1( us13_n780 ) , .ZN( us13_n820 ) );
  NOR2_X1 us13_U408 (.ZN( us13_n662 ) , .A2( us13_n697 ) , .A1( us13_n729 ) );
  NOR2_X1 us13_U409 (.A2( us13_n697 ) , .ZN( us13_n716 ) , .A1( us13_n792 ) );
  NOR2_X1 us13_U41 (.ZN( us13_n707 ) , .A2( us13_n776 ) , .A1( us13_n800 ) );
  NOR2_X1 us13_U410 (.ZN( us13_n594 ) , .A2( us13_n697 ) , .A1( us13_n728 ) );
  NOR2_X1 us13_U411 (.ZN( us13_n580 ) , .A2( us13_n697 ) , .A1( us13_n791 ) );
  OAI221_X1 us13_U412 (.A( us13_n783 ) , .C2( us13_n784 ) , .B2( us13_n785 ) , .B1( us13_n786 ) , .ZN( us13_n796 ) , .C1( us13_n813 ) );
  OAI22_X1 us13_U413 (.ZN( us13_n588 ) , .A2( us13_n747 ) , .B2( us13_n762 ) , .A1( us13_n763 ) , .B1( us13_n784 ) );
  AOI21_X1 us13_U414 (.ZN( us13_n592 ) , .B1( us13_n728 ) , .B2( us13_n784 ) , .A( us13_n790 ) );
  OAI221_X1 us13_U415 (.A( us13_n696 ) , .ZN( us13_n703 ) , .C2( us13_n784 ) , .C1( us13_n785 ) , .B1( us13_n786 ) , .B2( us13_n806 ) );
  NAND2_X1 us13_U416 (.A1( us13_n729 ) , .A2( us13_n784 ) , .ZN( us13_n811 ) );
  AOI21_X1 us13_U417 (.ZN( us13_n623 ) , .B1( us13_n699 ) , .A( us13_n779 ) , .B2( us13_n784 ) );
  AOI21_X1 us13_U418 (.ZN( us13_n648 ) , .A( us13_n762 ) , .B2( us13_n784 ) , .B1( us13_n792 ) );
  OAI22_X1 us13_U419 (.ZN( us13_n681 ) , .A1( us13_n699 ) , .A2( us13_n730 ) , .B2( us13_n784 ) , .B1( us13_n817 ) );
  NOR2_X1 us13_U42 (.ZN( us13_n804 ) , .A1( us13_n854 ) , .A2( us13_n861 ) );
  NOR2_X1 us13_U420 (.ZN( us13_n651 ) , .A1( us13_n784 ) , .A2( us13_n788 ) );
  NOR2_X1 us13_U421 (.ZN( us13_n553 ) , .A2( us13_n744 ) , .A1( us13_n784 ) );
  OAI21_X1 us13_U422 (.A( us13_n613 ) , .ZN( us13_n616 ) , .B1( us13_n625 ) , .B2( us13_n784 ) );
  NOR2_X1 us13_U423 (.ZN( us13_n610 ) , .A1( us13_n784 ) , .A2( us13_n816 ) );
  OAI222_X1 us13_U424 (.A2( us13_n669 ) , .ZN( us13_n674 ) , .B1( us13_n747 ) , .B2( us13_n784 ) , .C2( us13_n788 ) , .C1( us13_n815 ) , .A1( us13_n817 ) );
  NOR2_X1 us13_U425 (.ZN( us13_n600 ) , .A2( us13_n697 ) , .A1( us13_n784 ) );
  INV_X1 us13_U426 (.A( us13_n784 ) , .ZN( us13_n861 ) );
  NAND2_X1 us13_U427 (.A1( us13_n454 ) , .A2( us13_n461 ) , .ZN( us13_n813 ) );
  NOR2_X1 us13_U428 (.ZN( us13_n789 ) , .A2( us13_n862 ) , .A1( us13_n868 ) );
  AOI221_X1 us13_U429 (.A( us13_n483 ) , .ZN( us13_n488 ) , .B1( us13_n831 ) , .C2( us13_n844 ) , .C1( us13_n852 ) , .B2( us13_n862 ) );
  AOI222_X1 us13_U43 (.B2( us13_n638 ) , .ZN( us13_n644 ) , .B1( us13_n841 ) , .A1( us13_n842 ) , .C2( us13_n846 ) , .C1( us13_n863 ) , .A2( us13_n865 ) );
  AOI221_X1 us13_U430 (.A( us13_n681 ) , .ZN( us13_n692 ) , .B2( us13_n840 ) , .C1( us13_n842 ) , .C2( us13_n862 ) , .B1( us13_n865 ) );
  AOI222_X1 us13_U431 (.ZN( us13_n605 ) , .B2( us13_n671 ) , .B1( us13_n753 ) , .C2( us13_n831 ) , .A1( us13_n833 ) , .A2( us13_n862 ) , .C1( us13_n863 ) );
  INV_X1 us13_U432 (.A( us13_n786 ) , .ZN( us13_n862 ) );
  AND2_X1 us13_U433 (.ZN( us13_n438 ) , .A2( us13_n831 ) , .A1( us13_n854 ) );
  AND2_X1 us13_U434 (.ZN( us13_n439 ) , .A2( us13_n843 ) , .A1( us13_n861 ) );
  NOR3_X1 us13_U435 (.A1( us13_n438 ) , .A2( us13_n439 ) , .A3( us13_n576 ) , .ZN( us13_n587 ) );
  INV_X1 us13_U436 (.A( us13_n812 ) , .ZN( us13_n854 ) );
  NAND3_X1 us13_U437 (.ZN( sa12_sr_6 ) , .A3( us13_n797 ) , .A2( us13_n798 ) , .A1( us13_n799 ) );
  NAND3_X1 us13_U438 (.ZN( sa12_sr_5 ) , .A3( us13_n758 ) , .A2( us13_n759 ) , .A1( us13_n760 ) );
  NAND3_X1 us13_U439 (.ZN( sa12_sr_4 ) , .A3( us13_n738 ) , .A2( us13_n739 ) , .A1( us13_n740 ) );
  NOR4_X1 us13_U44 (.A4( us13_n639 ) , .A3( us13_n640 ) , .A2( us13_n641 ) , .A1( us13_n642 ) , .ZN( us13_n643 ) );
  NAND3_X1 us13_U440 (.A3( us13_n675 ) , .A2( us13_n676 ) , .A1( us13_n677 ) , .ZN( us13_n807 ) );
  NAND3_X1 us13_U441 (.ZN( us13_n638 ) , .A3( us13_n708 ) , .A2( us13_n724 ) , .A1( us13_n792 ) );
  NAND3_X1 us13_U442 (.A3( us13_n618 ) , .A2( us13_n619 ) , .A1( us13_n620 ) , .ZN( us13_n725 ) );
  NAND3_X1 us13_U443 (.A3( us13_n585 ) , .A2( us13_n586 ) , .A1( us13_n587 ) , .ZN( us13_n621 ) );
  NAND3_X1 us13_U444 (.ZN( us13_n565 ) , .A3( us13_n680 ) , .A2( us13_n750 ) , .A1( us13_n785 ) );
  NAND3_X1 us13_U445 (.A3( us13_n523 ) , .A2( us13_n524 ) , .A1( us13_n525 ) , .ZN( us13_n742 ) );
  NAND3_X1 us13_U446 (.A3( us13_n512 ) , .A1( us13_n513 ) , .ZN( us13_n608 ) , .A2( us13_n871 ) );
  NAND3_X1 us13_U447 (.A3( us13_n467 ) , .A2( us13_n468 ) , .A1( us13_n469 ) , .ZN( us13_n777 ) );
  INV_X1 us13_U448 (.A( us13_n803 ) , .ZN( us13_n843 ) );
  AOI21_X1 us13_U449 (.ZN( us13_n576 ) , .B2( us13_n724 ) , .B1( us13_n748 ) , .A( us13_n785 ) );
  NOR3_X1 us13_U45 (.A2( us13_n607 ) , .A1( us13_n608 ) , .ZN( us13_n646 ) , .A3( us13_n722 ) );
  NAND4_X1 us13_U46 (.ZN( sa12_sr_0 ) , .A4( us13_n501 ) , .A3( us13_n502 ) , .A2( us13_n503 ) , .A1( us13_n504 ) );
  AOI221_X1 us13_U47 (.A( us13_n497 ) , .ZN( us13_n502 ) , .B2( us13_n843 ) , .C1( us13_n846 ) , .C2( us13_n860 ) , .B1( us13_n862 ) );
  NOR4_X1 us13_U48 (.A4( us13_n498 ) , .A3( us13_n499 ) , .A2( us13_n500 ) , .ZN( us13_n501 ) , .A1( us13_n527 ) );
  AOI211_X1 us13_U49 (.A( us13_n496 ) , .ZN( us13_n503 ) , .B( us13_n802 ) , .C2( us13_n839 ) , .C1( us13_n851 ) );
  NAND2_X1 us13_U5 (.A2( us13_n471 ) , .A1( us13_n472 ) , .ZN( us13_n817 ) );
  NAND4_X1 us13_U50 (.ZN( sa12_sr_1 ) , .A4( us13_n595 ) , .A3( us13_n596 ) , .A2( us13_n597 ) , .A1( us13_n598 ) );
  AOI211_X1 us13_U51 (.B( us13_n589 ) , .A( us13_n590 ) , .ZN( us13_n596 ) , .C2( us13_n811 ) , .C1( us13_n833 ) );
  NOR4_X1 us13_U52 (.A4( us13_n591 ) , .A3( us13_n592 ) , .A2( us13_n593 ) , .A1( us13_n594 ) , .ZN( us13_n595 ) );
  AOI211_X1 us13_U53 (.A( us13_n588 ) , .ZN( us13_n597 ) , .B( us13_n621 ) , .C1( us13_n845 ) , .C2( us13_n855 ) );
  NOR2_X1 us13_U54 (.ZN( us13_n748 ) , .A1( us13_n861 ) , .A2( us13_n862 ) );
  NAND4_X1 us13_U55 (.ZN( sa12_sr_7 ) , .A4( us13_n822 ) , .A3( us13_n823 ) , .A2( us13_n824 ) , .A1( us13_n825 ) );
  AOI222_X1 us13_U56 (.C2( us13_n809 ) , .B2( us13_n810 ) , .A2( us13_n811 ) , .ZN( us13_n823 ) , .C1( us13_n832 ) , .A1( us13_n839 ) , .B1( us13_n853 ) );
  NOR4_X1 us13_U57 (.A4( us13_n818 ) , .A3( us13_n819 ) , .A2( us13_n820 ) , .A1( us13_n821 ) , .ZN( us13_n822 ) );
  AOI211_X1 us13_U58 (.B( us13_n807 ) , .A( us13_n808 ) , .ZN( us13_n824 ) , .C1( us13_n842 ) , .C2( us13_n850 ) );
  NOR2_X1 us13_U59 (.ZN( us13_n625 ) , .A2( us13_n836 ) , .A1( us13_n839 ) );
  NOR3_X1 us13_U6 (.ZN( us13_n598 ) , .A1( us13_n608 ) , .A3( us13_n723 ) , .A2( us13_n742 ) );
  NAND4_X1 us13_U60 (.A4( us13_n603 ) , .A3( us13_n604 ) , .A2( us13_n605 ) , .A1( us13_n606 ) , .ZN( us13_n722 ) );
  NOR3_X1 us13_U61 (.A1( us13_n599 ) , .ZN( us13_n604 ) , .A3( us13_n663 ) , .A2( us13_n770 ) );
  NOR4_X1 us13_U62 (.A3( us13_n600 ) , .A2( us13_n601 ) , .A1( us13_n602 ) , .ZN( us13_n603 ) , .A4( us13_n655 ) );
  AOI222_X1 us13_U63 (.ZN( us13_n606 ) , .A1( us13_n830 ) , .C2( us13_n837 ) , .B1( us13_n842 ) , .A2( us13_n856 ) , .B2( us13_n861 ) , .C1( us13_n868 ) );
  AOI222_X1 us13_U64 (.ZN( us13_n469 ) , .B1( us13_n832 ) , .A1( us13_n839 ) , .C1( us13_n842 ) , .C2( us13_n851 ) , .A2( us13_n855 ) , .B2( us13_n865 ) );
  NOR4_X1 us13_U65 (.A1( us13_n466 ) , .ZN( us13_n467 ) , .A4( us13_n542 ) , .A2( us13_n554 ) , .A3( us13_n614 ) );
  AOI221_X1 us13_U66 (.ZN( us13_n468 ) , .C2( us13_n714 ) , .B2( us13_n831 ) , .C1( us13_n845 ) , .B1( us13_n860 ) , .A( us13_n864 ) );
  NAND4_X1 us13_U67 (.A4( us13_n485 ) , .A3( us13_n486 ) , .A2( us13_n487 ) , .A1( us13_n488 ) , .ZN( us13_n778 ) );
  NOR4_X1 us13_U68 (.A4( us13_n484 ) , .ZN( us13_n487 ) , .A1( us13_n566 ) , .A2( us13_n581 ) , .A3( us13_n602 ) );
  NOR4_X1 us13_U69 (.ZN( us13_n486 ) , .A1( us13_n507 ) , .A2( us13_n519 ) , .A4( us13_n546 ) , .A3( us13_n611 ) );
  NOR3_X1 us13_U7 (.A3( us13_n800 ) , .A2( us13_n801 ) , .A1( us13_n802 ) , .ZN( us13_n825 ) );
  NOR4_X1 us13_U70 (.A4( us13_n514 ) , .A3( us13_n515 ) , .A2( us13_n516 ) , .A1( us13_n517 ) , .ZN( us13_n524 ) );
  AOI222_X1 us13_U71 (.ZN( us13_n525 ) , .A1( us13_n834 ) , .B2( us13_n837 ) , .C1( us13_n844 ) , .C2( us13_n850 ) , .A2( us13_n852 ) , .B1( us13_n866 ) );
  NOR4_X1 us13_U72 (.A3( us13_n521 ) , .A1( us13_n522 ) , .ZN( us13_n523 ) , .A2( us13_n673 ) , .A4( us13_n769 ) );
  NAND4_X1 us13_U73 (.A4( us13_n657 ) , .A3( us13_n658 ) , .A2( us13_n659 ) , .A1( us13_n660 ) , .ZN( us13_n800 ) );
  NOR3_X1 us13_U74 (.A3( us13_n651 ) , .A2( us13_n652 ) , .A1( us13_n653 ) , .ZN( us13_n658 ) );
  NOR3_X1 us13_U75 (.A3( us13_n648 ) , .A2( us13_n649 ) , .A1( us13_n650 ) , .ZN( us13_n659 ) );
  NOR3_X1 us13_U76 (.A3( us13_n654 ) , .A2( us13_n655 ) , .A1( us13_n656 ) , .ZN( us13_n657 ) );
  NAND4_X1 us13_U77 (.A4( us13_n560 ) , .A3( us13_n561 ) , .A2( us13_n562 ) , .A1( us13_n563 ) , .ZN( us13_n607 ) );
  NOR4_X1 us13_U78 (.A4( us13_n552 ) , .A3( us13_n553 ) , .A2( us13_n554 ) , .A1( us13_n555 ) , .ZN( us13_n562 ) );
  NOR4_X1 us13_U79 (.ZN( us13_n561 ) , .A1( us13_n653 ) , .A3( us13_n661 ) , .A4( us13_n685 ) , .A2( us13_n768 ) );
  NOR3_X1 us13_U8 (.ZN( us13_n504 ) , .A2( us13_n679 ) , .A3( us13_n777 ) , .A1( us13_n876 ) );
  NOR4_X1 us13_U80 (.A4( us13_n556 ) , .A3( us13_n557 ) , .A2( us13_n558 ) , .A1( us13_n559 ) , .ZN( us13_n560 ) );
  NAND4_X1 us13_U81 (.A4( us13_n772 ) , .A3( us13_n773 ) , .A2( us13_n774 ) , .A1( us13_n775 ) , .ZN( us13_n801 ) );
  NOR3_X1 us13_U82 (.A3( us13_n765 ) , .A2( us13_n766 ) , .A1( us13_n767 ) , .ZN( us13_n773 ) );
  AOI222_X1 us13_U83 (.ZN( us13_n775 ) , .A1( us13_n830 ) , .C1( us13_n834 ) , .B2( us13_n841 ) , .A2( us13_n850 ) , .B1( us13_n861 ) , .C2( us13_n873 ) );
  NOR4_X1 us13_U84 (.A4( us13_n768 ) , .A3( us13_n769 ) , .A2( us13_n770 ) , .A1( us13_n771 ) , .ZN( us13_n772 ) );
  NAND4_X1 us13_U85 (.A4( us13_n691 ) , .A3( us13_n692 ) , .A1( us13_n693 ) , .ZN( us13_n776 ) , .A2( us13_n872 ) );
  INV_X1 us13_U86 (.A( us13_n679 ) , .ZN( us13_n872 ) );
  NOR4_X1 us13_U87 (.A4( us13_n687 ) , .A3( us13_n688 ) , .A2( us13_n689 ) , .A1( us13_n690 ) , .ZN( us13_n691 ) );
  NOR4_X1 us13_U88 (.A4( us13_n661 ) , .A3( us13_n662 ) , .A2( us13_n663 ) , .A1( us13_n664 ) , .ZN( us13_n677 ) );
  NOR4_X1 us13_U89 (.A4( us13_n665 ) , .A3( us13_n666 ) , .A2( us13_n667 ) , .A1( us13_n668 ) , .ZN( us13_n676 ) );
  INV_X1 us13_U9 (.A( us13_n706 ) , .ZN( us13_n876 ) );
  NOR4_X1 us13_U90 (.A3( us13_n673 ) , .A1( us13_n674 ) , .ZN( us13_n675 ) , .A4( us13_n715 ) , .A2( us13_n859 ) );
  NOR2_X1 us13_U91 (.ZN( us13_n761 ) , .A1( us13_n833 ) , .A2( us13_n834 ) );
  NOR4_X1 us13_U92 (.A4( us13_n577 ) , .A3( us13_n578 ) , .A2( us13_n579 ) , .ZN( us13_n586 ) , .A1( us13_n683 ) );
  NOR4_X1 us13_U93 (.A1( us13_n584 ) , .ZN( us13_n585 ) , .A3( us13_n652 ) , .A2( us13_n662 ) , .A4( us13_n767 ) );
  AOI222_X1 us13_U94 (.ZN( us13_n513 ) , .C1( us13_n832 ) , .B2( us13_n837 ) , .A2( us13_n843 ) , .C2( us13_n862 ) , .B1( us13_n863 ) , .A1( us13_n866 ) );
  NOR4_X1 us13_U95 (.A4( us13_n509 ) , .A2( us13_n510 ) , .A1( us13_n511 ) , .ZN( us13_n512 ) , .A3( us13_n670 ) );
  INV_X1 us13_U96 (.A( us13_n505 ) , .ZN( us13_n871 ) );
  NAND4_X1 us13_U97 (.A4( us13_n456 ) , .A3( us13_n457 ) , .A2( us13_n458 ) , .A1( us13_n459 ) , .ZN( us13_n679 ) );
  NOR3_X1 us13_U98 (.ZN( us13_n457 ) , .A3( us13_n530 ) , .A1( us13_n555 ) , .A2( us13_n570 ) );
  AOI221_X1 us13_U99 (.A( us13_n450 ) , .ZN( us13_n459 ) , .C2( us13_n753 ) , .B1( us13_n832 ) , .C1( us13_n842 ) , .B2( us13_n861 ) );
  INV_X1 us20_U10 (.A( us20_n706 ) , .ZN( us20_n876 ) );
  NOR4_X1 us20_U100 (.A1( us20_n531 ) , .ZN( us20_n536 ) , .A2( us20_n654 ) , .A4( us20_n668 ) , .A3( us20_n765 ) );
  NOR4_X1 us20_U101 (.A4( us20_n529 ) , .A3( us20_n530 ) , .ZN( us20_n537 ) , .A2( us20_n684 ) , .A1( us20_n794 ) );
  NAND4_X1 us20_U102 (.A4( us20_n548 ) , .A3( us20_n549 ) , .A2( us20_n550 ) , .A1( us20_n551 ) , .ZN( us20_n745 ) );
  NOR3_X1 us20_U103 (.ZN( us20_n549 ) , .A2( us20_n651 ) , .A1( us20_n667 ) , .A3( us20_n771 ) );
  AOI211_X1 us20_U104 (.B( us20_n539 ) , .A( us20_n540 ) , .ZN( us20_n551 ) , .C2( us20_n839 ) , .C1( us20_n851 ) );
  NOR4_X1 us20_U105 (.A4( us20_n541 ) , .A3( us20_n542 ) , .A2( us20_n543 ) , .ZN( us20_n550 ) , .A1( us20_n688 ) );
  NAND4_X1 us20_U106 (.A4( us20_n479 ) , .A3( us20_n480 ) , .A2( us20_n481 ) , .A1( us20_n482 ) , .ZN( us20_n694 ) );
  NOR3_X1 us20_U107 (.ZN( us20_n480 ) , .A2( us20_n508 ) , .A3( us20_n601 ) , .A1( us20_n610 ) );
  AOI211_X1 us20_U108 (.B( us20_n477 ) , .A( us20_n478 ) , .ZN( us20_n482 ) , .C2( us20_n833 ) , .C1( us20_n861 ) );
  NOR4_X1 us20_U109 (.ZN( us20_n481 ) , .A3( us20_n532 ) , .A4( us20_n545 ) , .A2( us20_n567 ) , .A1( us20_n717 ) );
  INV_X1 us20_U11 (.A( us20_n607 ) , .ZN( us20_n874 ) );
  NOR2_X1 us20_U110 (.ZN( us20_n647 ) , .A1( us20_n854 ) , .A2( us20_n868 ) );
  NAND4_X1 us20_U111 (.A4( us20_n473 ) , .A3( us20_n474 ) , .A2( us20_n475 ) , .A1( us20_n476 ) , .ZN( us20_n678 ) );
  NOR4_X1 us20_U112 (.ZN( us20_n475 ) , .A1( us20_n531 ) , .A3( us20_n568 ) , .A4( us20_n600 ) , .A2( us20_n642 ) );
  NOR4_X1 us20_U113 (.A4( us20_n470 ) , .ZN( us20_n476 ) , .A3( us20_n556 ) , .A1( us20_n735 ) , .A2( us20_n755 ) );
  NOR4_X1 us20_U114 (.ZN( us20_n474 ) , .A1( us20_n506 ) , .A3( us20_n544 ) , .A2( us20_n583 ) , .A4( us20_n716 ) );
  NAND4_X1 us20_U115 (.A4( us20_n691 ) , .A3( us20_n692 ) , .A1( us20_n693 ) , .ZN( us20_n776 ) , .A2( us20_n872 ) );
  INV_X1 us20_U116 (.A( us20_n679 ) , .ZN( us20_n872 ) );
  AOI221_X1 us20_U117 (.A( us20_n681 ) , .ZN( us20_n692 ) , .B2( us20_n840 ) , .C1( us20_n842 ) , .C2( us20_n862 ) , .B1( us20_n865 ) );
  NOR4_X1 us20_U118 (.A4( us20_n687 ) , .A3( us20_n688 ) , .A2( us20_n689 ) , .A1( us20_n690 ) , .ZN( us20_n691 ) );
  NOR2_X1 us20_U119 (.ZN( us20_n733 ) , .A2( us20_n832 ) , .A1( us20_n845 ) );
  INV_X1 us20_U12 (.A( us20_n680 ) , .ZN( us20_n840 ) );
  NAND4_X1 us20_U120 (.A4( us20_n719 ) , .A3( us20_n720 ) , .A2( us20_n721 ) , .ZN( us20_n741 ) , .A1( us20_n857 ) );
  INV_X1 us20_U121 (.A( us20_n709 ) , .ZN( us20_n857 ) );
  NOR4_X1 us20_U122 (.A4( us20_n715 ) , .A3( us20_n716 ) , .A2( us20_n717 ) , .A1( us20_n718 ) , .ZN( us20_n719 ) );
  AOI221_X1 us20_U123 (.A( us20_n710 ) , .ZN( us20_n721 ) , .C2( us20_n844 ) , .B2( us20_n845 ) , .C1( us20_n861 ) , .B1( us20_n862 ) );
  NAND4_X1 us20_U124 (.A4( us20_n573 ) , .A3( us20_n574 ) , .A1( us20_n575 ) , .ZN( us20_n723 ) , .A2( us20_n874 ) );
  NOR4_X1 us20_U125 (.A4( us20_n569 ) , .A3( us20_n570 ) , .A2( us20_n571 ) , .A1( us20_n572 ) , .ZN( us20_n573 ) );
  AOI221_X1 us20_U126 (.A( us20_n564 ) , .C2( us20_n565 ) , .ZN( us20_n574 ) , .B2( us20_n845 ) , .B1( us20_n852 ) , .C1( us20_n853 ) );
  NOR2_X1 us20_U127 (.ZN( us20_n575 ) , .A1( us20_n622 ) , .A2( us20_n745 ) );
  NAND4_X1 us20_U128 (.A4( us20_n633 ) , .A3( us20_n634 ) , .A2( us20_n635 ) , .A1( us20_n636 ) , .ZN( us20_n743 ) );
  AOI211_X1 us20_U129 (.B( us20_n623 ) , .A( us20_n624 ) , .ZN( us20_n635 ) , .C2( us20_n836 ) , .C1( us20_n863 ) );
  NOR4_X1 us20_U13 (.A4( us20_n445 ) , .A3( us20_n446 ) , .A2( us20_n516 ) , .A1( us20_n541 ) , .ZN( us20_n706 ) );
  NOR4_X1 us20_U130 (.A4( us20_n629 ) , .A3( us20_n630 ) , .A2( us20_n631 ) , .A1( us20_n632 ) , .ZN( us20_n633 ) );
  NOR4_X1 us20_U131 (.A4( us20_n626 ) , .A3( us20_n627 ) , .A2( us20_n628 ) , .ZN( us20_n634 ) , .A1( us20_n664 ) );
  NAND4_X1 us20_U132 (.A4( us20_n493 ) , .A3( us20_n494 ) , .A1( us20_n495 ) , .ZN( us20_n802 ) , .A2( us20_n867 ) );
  AOI221_X1 us20_U133 (.A( us20_n489 ) , .ZN( us20_n494 ) , .B2( us20_n836 ) , .C2( us20_n841 ) , .C1( us20_n851 ) , .B1( us20_n860 ) );
  INV_X1 us20_U134 (.A( us20_n778 ) , .ZN( us20_n867 ) );
  NOR4_X1 us20_U135 (.A2( us20_n491 ) , .A1( us20_n492 ) , .ZN( us20_n493 ) , .A3( us20_n580 ) , .A4( us20_n612 ) );
  INV_X1 us20_U136 (.A( us20_n762 ) , .ZN( us20_n830 ) );
  OR4_X1 us20_U137 (.A4( us20_n580 ) , .A3( us20_n581 ) , .A2( us20_n582 ) , .A1( us20_n583 ) , .ZN( us20_n584 ) );
  OR4_X1 us20_U138 (.A4( us20_n566 ) , .A3( us20_n567 ) , .A2( us20_n568 ) , .ZN( us20_n572 ) , .A1( us20_n665 ) );
  OR4_X1 us20_U139 (.A4( us20_n682 ) , .A3( us20_n683 ) , .A2( us20_n684 ) , .A1( us20_n685 ) , .ZN( us20_n690 ) );
  OR3_X1 us20_U14 (.ZN( us20_n446 ) , .A1( us20_n528 ) , .A3( us20_n577 ) , .A2( us20_n875 ) );
  OR4_X1 us20_U140 (.ZN( us20_n466 ) , .A4( us20_n518 ) , .A3( us20_n529 ) , .A2( us20_n578 ) , .A1( us20_n712 ) );
  OR4_X1 us20_U141 (.A4( us20_n518 ) , .A2( us20_n519 ) , .A1( us20_n520 ) , .ZN( us20_n522 ) , .A3( us20_n821 ) );
  OR4_X1 us20_U142 (.ZN( us20_n492 ) , .A4( us20_n534 ) , .A2( us20_n547 ) , .A1( us20_n559 ) , .A3( us20_n632 ) );
  NAND2_X1 us20_U143 (.ZN( us20_n613 ) , .A2( us20_n837 ) , .A1( us20_n873 ) );
  OR3_X1 us20_U144 (.A3( us20_n506 ) , .A2( us20_n507 ) , .A1( us20_n508 ) , .ZN( us20_n511 ) );
  AOI221_X1 us20_U145 (.A( us20_n713 ) , .B2( us20_n714 ) , .ZN( us20_n720 ) , .C1( us20_n832 ) , .B1( us20_n839 ) , .C2( us20_n863 ) );
  OR2_X1 us20_U146 (.A2( us20_n711 ) , .A1( us20_n712 ) , .ZN( us20_n713 ) );
  INV_X1 us20_U147 (.A( us20_n463 ) , .ZN( us20_n864 ) );
  OAI21_X1 us20_U148 (.ZN( us20_n463 ) , .B1( us20_n809 ) , .A( us20_n834 ) , .B2( us20_n851 ) );
  INV_X1 us20_U149 (.A( us20_n754 ) , .ZN( us20_n869 ) );
  OR4_X1 us20_U15 (.A4( us20_n442 ) , .A2( us20_n443 ) , .A1( us20_n444 ) , .ZN( us20_n445 ) , .A3( us20_n553 ) );
  OAI21_X1 us20_U150 (.B1( us20_n753 ) , .ZN( us20_n754 ) , .A( us20_n845 ) , .B2( us20_n868 ) );
  AOI222_X1 us20_U151 (.ZN( us20_n660 ) , .A2( us20_n839 ) , .B1( us20_n841 ) , .C2( us20_n845 ) , .A1( us20_n860 ) , .C1( us20_n863 ) , .B2( us20_n870 ) );
  INV_X1 us20_U152 (.A( us20_n647 ) , .ZN( us20_n870 ) );
  INV_X1 us20_U153 (.A( us20_n672 ) , .ZN( us20_n859 ) );
  AOI21_X1 us20_U154 (.A( us20_n670 ) , .B1( us20_n671 ) , .ZN( us20_n672 ) , .B2( us20_n856 ) );
  OAI22_X1 us20_U155 (.ZN( us20_n483 ) , .A1( us20_n708 ) , .B2( us20_n785 ) , .A2( us20_n806 ) , .B1( us20_n812 ) );
  OAI222_X1 us20_U156 (.B2( us20_n747 ) , .B1( us20_n748 ) , .A2( us20_n749 ) , .ZN( us20_n757 ) , .C2( us20_n805 ) , .C1( us20_n814 ) , .A1( us20_n817 ) );
  OAI222_X1 us20_U157 (.B2( us20_n708 ) , .ZN( us20_n709 ) , .C2( us20_n724 ) , .B1( us20_n747 ) , .A1( us20_n806 ) , .C1( us20_n814 ) , .A2( us20_n815 ) );
  OAI222_X1 us20_U158 (.ZN( us20_n505 ) , .C2( us20_n625 ) , .B2( us20_n647 ) , .B1( us20_n747 ) , .A2( us20_n748 ) , .C1( us20_n805 ) , .A1( us20_n806 ) );
  NAND2_X1 us20_U159 (.A1( us20_n447 ) , .A2( us20_n465 ) , .ZN( us20_n749 ) );
  INV_X1 us20_U16 (.A( us20_n613 ) , .ZN( us20_n875 ) );
  AOI22_X1 us20_U160 (.ZN( us20_n696 ) , .A1( us20_n830 ) , .B2( us20_n843 ) , .A2( us20_n865 ) , .B1( us20_n868 ) );
  AOI22_X1 us20_U161 (.A2( us20_n782 ) , .ZN( us20_n783 ) , .B2( us20_n831 ) , .A1( us20_n834 ) , .B1( us20_n863 ) );
  INV_X1 us20_U162 (.A( us20_n730 ) , .ZN( us20_n839 ) );
  INV_X1 us20_U163 (.A( us20_n790 ) , .ZN( us20_n832 ) );
  NAND2_X1 us20_U164 (.A1( us20_n451 ) , .A2( us20_n453 ) , .ZN( us20_n762 ) );
  AOI211_X1 us20_U165 (.A( us20_n637 ) , .ZN( us20_n645 ) , .B( us20_n743 ) , .C2( us20_n839 ) , .C1( us20_n854 ) );
  OAI22_X1 us20_U166 (.ZN( us20_n637 ) , .A1( us20_n699 ) , .B2( us20_n728 ) , .A2( us20_n762 ) , .B1( us20_n816 ) );
  OAI221_X1 us20_U167 (.A( us20_n727 ) , .C2( us20_n728 ) , .B2( us20_n729 ) , .B1( us20_n730 ) , .ZN( us20_n737 ) , .C1( us20_n817 ) );
  AOI22_X1 us20_U168 (.ZN( us20_n727 ) , .B1( us20_n832 ) , .A2( us20_n838 ) , .A1( us20_n863 ) , .B2( us20_n866 ) );
  OAI22_X1 us20_U169 (.ZN( us20_n489 ) , .A1( us20_n724 ) , .B2( us20_n728 ) , .B1( us20_n730 ) , .A2( us20_n779 ) );
  INV_X1 us20_U17 (.A( us20_n749 ) , .ZN( us20_n863 ) );
  OAI22_X1 us20_U170 (.ZN( us20_n624 ) , .B1( us20_n669 ) , .B2( us20_n747 ) , .A1( us20_n815 ) , .A2( us20_n816 ) );
  OAI22_X1 us20_U171 (.B2( us20_n779 ) , .B1( us20_n780 ) , .ZN( us20_n781 ) , .A2( us20_n814 ) , .A1( us20_n815 ) );
  OAI22_X1 us20_U172 (.A1( us20_n724 ) , .ZN( us20_n726 ) , .B2( us20_n750 ) , .B1( us20_n812 ) , .A2( us20_n816 ) );
  OAI22_X1 us20_U173 (.B2( us20_n744 ) , .ZN( us20_n746 ) , .A2( us20_n762 ) , .B1( us20_n780 ) , .A1( us20_n792 ) );
  OAI22_X1 us20_U174 (.ZN( us20_n496 ) , .A2( us20_n744 ) , .A1( us20_n780 ) , .B1( us20_n791 ) , .B2( us20_n806 ) );
  OAI22_X1 us20_U175 (.B2( us20_n803 ) , .B1( us20_n804 ) , .A2( us20_n805 ) , .A1( us20_n806 ) , .ZN( us20_n808 ) );
  INV_X1 us20_U176 (.A( us20_n788 ) , .ZN( us20_n845 ) );
  INV_X1 us20_U177 (.A( us20_n744 ) , .ZN( us20_n837 ) );
  INV_X1 us20_U178 (.A( us20_n814 ) , .ZN( us20_n833 ) );
  OAI22_X1 us20_U179 (.B1( us20_n490 ) , .ZN( us20_n491 ) , .A1( us20_n686 ) , .A2( us20_n763 ) , .B2( us20_n817 ) );
  AOI222_X1 us20_U18 (.ZN( us20_n563 ) , .B1( us20_n830 ) , .C1( us20_n841 ) , .A2( us20_n843 ) , .A1( us20_n854 ) , .B2( us20_n863 ) , .C2( us20_n873 ) );
  NOR3_X1 us20_U180 (.ZN( us20_n490 ) , .A1( us20_n782 ) , .A2( us20_n850 ) , .A3( us20_n863 ) );
  OAI22_X1 us20_U181 (.ZN( us20_n695 ) , .A2( us20_n730 ) , .A1( us20_n780 ) , .B1( us20_n791 ) , .B2( us20_n817 ) );
  INV_X1 us20_U182 (.A( us20_n805 ) , .ZN( us20_n860 ) );
  INV_X1 us20_U183 (.A( us20_n669 ) , .ZN( us20_n865 ) );
  NOR2_X1 us20_U184 (.ZN( us20_n715 ) , .A1( us20_n805 ) , .A2( us20_n817 ) );
  NOR2_X1 us20_U185 (.ZN( us20_n666 ) , .A1( us20_n728 ) , .A2( us20_n803 ) );
  NOR2_X1 us20_U186 (.ZN( us20_n546 ) , .A2( us20_n780 ) , .A1( us20_n814 ) );
  NOR2_X1 us20_U187 (.ZN( us20_n577 ) , .A2( us20_n699 ) , .A1( us20_n814 ) );
  NOR2_X1 us20_U188 (.ZN( us20_n570 ) , .A1( us20_n728 ) , .A2( us20_n806 ) );
  NOR2_X1 us20_U189 (.A2( us20_n744 ) , .ZN( us20_n755 ) , .A1( us20_n805 ) );
  NOR4_X1 us20_U19 (.ZN( us20_n473 ) , .A2( us20_n521 ) , .A4( us20_n594 ) , .A1( us20_n609 ) , .A3( us20_n629 ) );
  NOR2_X1 us20_U190 (.ZN( us20_n718 ) , .A2( us20_n724 ) , .A1( us20_n744 ) );
  NOR2_X1 us20_U191 (.ZN( us20_n735 ) , .A2( us20_n803 ) , .A1( us20_n805 ) );
  INV_X1 us20_U192 (.A( us20_n750 ) , .ZN( us20_n842 ) );
  NOR2_X1 us20_U193 (.ZN( us20_n532 ) , .A2( us20_n749 ) , .A1( us20_n750 ) );
  NOR2_X1 us20_U194 (.ZN( us20_n654 ) , .A1( us20_n728 ) , .A2( us20_n813 ) );
  NOR2_X1 us20_U195 (.ZN( us20_n615 ) , .A1( us20_n785 ) , .A2( us20_n815 ) );
  NOR2_X1 us20_U196 (.ZN( us20_n629 ) , .A2( us20_n728 ) , .A1( us20_n785 ) );
  NOR2_X1 us20_U197 (.ZN( us20_n628 ) , .A2( us20_n669 ) , .A1( us20_n785 ) );
  NOR2_X1 us20_U198 (.ZN( us20_n611 ) , .A2( us20_n780 ) , .A1( us20_n806 ) );
  INV_X1 us20_U199 (.A( us20_n747 ) , .ZN( us20_n834 ) );
  NOR4_X1 us20_U20 (.A4( us20_n544 ) , .A3( us20_n545 ) , .A2( us20_n546 ) , .A1( us20_n547 ) , .ZN( us20_n548 ) );
  NOR2_X1 us20_U200 (.ZN( us20_n601 ) , .A2( us20_n780 ) , .A1( us20_n803 ) );
  NOR2_X1 us20_U201 (.A2( us20_n708 ) , .A1( us20_n750 ) , .ZN( us20_n771 ) );
  NOR2_X1 us20_U202 (.ZN( us20_n652 ) , .A1( us20_n669 ) , .A2( us20_n814 ) );
  INV_X1 us20_U203 (.A( us20_n792 ) , .ZN( us20_n851 ) );
  NOR2_X1 us20_U204 (.A1( us20_n669 ) , .ZN( us20_n673 ) , .A2( us20_n744 ) );
  NOR2_X1 us20_U205 (.ZN( us20_n602 ) , .A1( us20_n669 ) , .A2( us20_n803 ) );
  NOR2_X1 us20_U206 (.A1( us20_n669 ) , .ZN( us20_n688 ) , .A2( us20_n816 ) );
  NOR2_X1 us20_U207 (.ZN( us20_n667 ) , .A1( us20_n750 ) , .A2( us20_n815 ) );
  NOR2_X1 us20_U208 (.A2( us20_n744 ) , .ZN( us20_n769 ) , .A1( us20_n812 ) );
  NOR2_X1 us20_U209 (.ZN( us20_n555 ) , .A1( us20_n750 ) , .A2( us20_n791 ) );
  NOR4_X1 us20_U21 (.ZN( us20_n479 ) , .A1( us20_n520 ) , .A4( us20_n557 ) , .A3( us20_n582 ) , .A2( us20_n630 ) );
  NOR2_X1 us20_U210 (.ZN( us20_n528 ) , .A2( us20_n724 ) , .A1( us20_n803 ) );
  NOR2_X1 us20_U211 (.ZN( us20_n508 ) , .A2( us20_n780 ) , .A1( us20_n785 ) );
  NOR2_X1 us20_U212 (.ZN( us20_n543 ) , .A2( us20_n708 ) , .A1( us20_n785 ) );
  NOR2_X1 us20_U213 (.ZN( us20_n531 ) , .A2( us20_n780 ) , .A1( us20_n816 ) );
  NOR2_X1 us20_U214 (.ZN( us20_n664 ) , .A1( us20_n785 ) , .A2( us20_n791 ) );
  NOR2_X1 us20_U215 (.ZN( us20_n599 ) , .A2( us20_n791 ) , .A1( us20_n816 ) );
  NOR2_X1 us20_U216 (.A1( us20_n669 ) , .ZN( us20_n766 ) , .A2( us20_n813 ) );
  NOR2_X1 us20_U217 (.A1( us20_n699 ) , .ZN( us20_n768 ) , .A2( us20_n813 ) );
  NOR2_X1 us20_U218 (.ZN( us20_n527 ) , .A1( us20_n669 ) , .A2( us20_n779 ) );
  OAI22_X1 us20_U219 (.B1( us20_n440 ) , .ZN( us20_n444 ) , .A2( us20_n728 ) , .A1( us20_n744 ) , .B2( us20_n749 ) );
  NOR4_X1 us20_U22 (.A4( us20_n532 ) , .A3( us20_n533 ) , .A2( us20_n534 ) , .ZN( us20_n535 ) , .A1( us20_n820 ) );
  NOR3_X1 us20_U220 (.ZN( us20_n440 ) , .A2( us20_n836 ) , .A3( us20_n837 ) , .A1( us20_n846 ) );
  OAI22_X1 us20_U221 (.ZN( us20_n710 ) , .A2( us20_n728 ) , .B2( us20_n729 ) , .A1( us20_n744 ) , .B1( us20_n813 ) );
  NOR2_X1 us20_U222 (.ZN( us20_n557 ) , .A1( us20_n792 ) , .A2( us20_n814 ) );
  NOR2_X1 us20_U223 (.ZN( us20_n545 ) , .A1( us20_n749 ) , .A2( us20_n814 ) );
  NOR2_X1 us20_U224 (.ZN( us20_n556 ) , .A1( us20_n762 ) , .A2( us20_n805 ) );
  NOR2_X1 us20_U225 (.ZN( us20_n661 ) , .A1( us20_n729 ) , .A2( us20_n790 ) );
  NOR2_X1 us20_U226 (.ZN( us20_n507 ) , .A1( us20_n812 ) , .A2( us20_n817 ) );
  INV_X1 us20_U227 (.A( us20_n806 ) , .ZN( us20_n841 ) );
  NOR2_X1 us20_U228 (.ZN( us20_n509 ) , .A1( us20_n729 ) , .A2( us20_n779 ) );
  NOR2_X1 us20_U229 (.ZN( us20_n544 ) , .A2( us20_n785 ) , .A1( us20_n792 ) );
  NOR4_X1 us20_U23 (.ZN( us20_n456 ) , .A2( us20_n517 ) , .A1( us20_n543 ) , .A3( us20_n579 ) , .A4( us20_n615 ) );
  OAI22_X1 us20_U230 (.B2( us20_n750 ) , .B1( us20_n751 ) , .A1( us20_n752 ) , .ZN( us20_n756 ) , .A2( us20_n806 ) );
  NOR2_X1 us20_U231 (.ZN( us20_n751 ) , .A2( us20_n852 ) , .A1( us20_n860 ) );
  NOR3_X1 us20_U232 (.ZN( us20_n752 ) , .A2( us20_n853 ) , .A1( us20_n863 ) , .A3( us20_n865 ) );
  NOR2_X1 us20_U233 (.ZN( us20_n530 ) , .A2( us20_n744 ) , .A1( us20_n792 ) );
  NOR2_X1 us20_U234 (.ZN( us20_n663 ) , .A1( us20_n729 ) , .A2( us20_n785 ) );
  INV_X1 us20_U235 (.A( us20_n728 ) , .ZN( us20_n852 ) );
  NOR2_X1 us20_U236 (.A1( us20_n749 ) , .ZN( us20_n767 ) , .A2( us20_n803 ) );
  NOR2_X1 us20_U237 (.ZN( us20_n506 ) , .A2( us20_n728 ) , .A1( us20_n762 ) );
  NOR2_X1 us20_U238 (.ZN( us20_n516 ) , .A1( us20_n708 ) , .A2( us20_n744 ) );
  NOR2_X1 us20_U239 (.ZN( us20_n614 ) , .A1( us20_n762 ) , .A2( us20_n812 ) );
  NOR2_X1 us20_U24 (.ZN( us20_n680 ) , .A2( us20_n834 ) , .A1( us20_n839 ) );
  NOR2_X1 us20_U240 (.ZN( us20_n670 ) , .A1( us20_n790 ) , .A2( us20_n805 ) );
  NOR2_X1 us20_U241 (.ZN( us20_n517 ) , .A1( us20_n708 ) , .A2( us20_n803 ) );
  NOR2_X1 us20_U242 (.ZN( us20_n558 ) , .A1( us20_n708 ) , .A2( us20_n816 ) );
  NOR2_X1 us20_U243 (.ZN( us20_n630 ) , .A1( us20_n747 ) , .A2( us20_n815 ) );
  NOR2_X1 us20_U244 (.ZN( us20_n655 ) , .A1( us20_n790 ) , .A2( us20_n815 ) );
  NOR2_X1 us20_U245 (.ZN( us20_n521 ) , .A1( us20_n790 ) , .A2( us20_n812 ) );
  NOR2_X1 us20_U246 (.ZN( us20_n668 ) , .A2( us20_n708 ) , .A1( us20_n790 ) );
  NOR2_X1 us20_U247 (.ZN( us20_n631 ) , .A1( us20_n724 ) , .A2( us20_n813 ) );
  NOR2_X1 us20_U248 (.ZN( us20_n656 ) , .A1( us20_n747 ) , .A2( us20_n780 ) );
  NOR2_X1 us20_U249 (.ZN( us20_n542 ) , .A1( us20_n762 ) , .A2( us20_n791 ) );
  NOR4_X1 us20_U25 (.ZN( us20_n620 ) , .A1( us20_n656 ) , .A3( us20_n666 ) , .A4( us20_n682 ) , .A2( us20_n766 ) );
  NOR2_X1 us20_U250 (.ZN( us20_n609 ) , .A2( us20_n724 ) , .A1( us20_n817 ) );
  AOI21_X1 us20_U251 (.B1( us20_n625 ) , .ZN( us20_n627 ) , .A( us20_n763 ) , .B2( us20_n814 ) );
  NOR2_X1 us20_U252 (.ZN( us20_n579 ) , .A2( us20_n708 ) , .A1( us20_n730 ) );
  NOR2_X1 us20_U253 (.ZN( us20_n533 ) , .A2( us20_n724 ) , .A1( us20_n730 ) );
  NOR2_X1 us20_U254 (.ZN( us20_n642 ) , .A2( us20_n788 ) , .A1( us20_n791 ) );
  NOR2_X1 us20_U255 (.A2( us20_n708 ) , .A1( us20_n762 ) , .ZN( us20_n794 ) );
  AOI21_X1 us20_U256 (.ZN( us20_n650 ) , .A( us20_n779 ) , .B1( us20_n792 ) , .B2( us20_n805 ) );
  AOI21_X1 us20_U257 (.A( us20_n815 ) , .B2( us20_n816 ) , .B1( us20_n817 ) , .ZN( us20_n818 ) );
  NOR2_X1 us20_U258 (.ZN( us20_n520 ) , .A2( us20_n708 ) , .A1( us20_n814 ) );
  NOR2_X1 us20_U259 (.ZN( us20_n582 ) , .A1( us20_n744 ) , .A2( us20_n815 ) );
  NOR4_X1 us20_U26 (.A4( us20_n609 ) , .A3( us20_n610 ) , .A2( us20_n611 ) , .A1( us20_n612 ) , .ZN( us20_n619 ) );
  AOI21_X1 us20_U260 (.ZN( us20_n515 ) , .A( us20_n729 ) , .B1( us20_n750 ) , .B2( us20_n803 ) );
  AOI21_X1 us20_U261 (.ZN( us20_n626 ) , .B2( us20_n669 ) , .A( us20_n790 ) , .B1( us20_n791 ) );
  AOI21_X1 us20_U262 (.ZN( us20_n499 ) , .B1( us20_n680 ) , .A( us20_n812 ) , .B2( us20_n816 ) );
  AOI21_X1 us20_U263 (.ZN( us20_n477 ) , .A( us20_n669 ) , .B1( us20_n750 ) , .B2( us20_n806 ) );
  NOR2_X1 us20_U264 (.ZN( us20_n559 ) , .A2( us20_n791 ) , .A1( us20_n803 ) );
  AOI21_X1 us20_U265 (.ZN( us20_n510 ) , .B2( us20_n669 ) , .A( us20_n730 ) , .B1( us20_n815 ) );
  NOR2_X1 us20_U266 (.ZN( us20_n519 ) , .A2( us20_n699 ) , .A1( us20_n816 ) );
  NOR2_X1 us20_U267 (.ZN( us20_n683 ) , .A2( us20_n699 ) , .A1( us20_n803 ) );
  NOR2_X1 us20_U268 (.ZN( us20_n581 ) , .A1( us20_n669 ) , .A2( us20_n788 ) );
  AOI21_X1 us20_U269 (.ZN( us20_n589 ) , .B2( us20_n699 ) , .B1( us20_n815 ) , .A( us20_n817 ) );
  NOR4_X1 us20_U27 (.A4( us20_n614 ) , .A3( us20_n615 ) , .A2( us20_n616 ) , .A1( us20_n617 ) , .ZN( us20_n618 ) );
  INV_X1 us20_U270 (.A( us20_n763 ) , .ZN( us20_n866 ) );
  AOI21_X1 us20_U271 (.ZN( us20_n498 ) , .A( us20_n724 ) , .B2( us20_n762 ) , .B1( us20_n814 ) );
  AOI21_X1 us20_U272 (.ZN( us20_n539 ) , .B2( us20_n812 ) , .A( us20_n814 ) , .B1( us20_n815 ) );
  AOI21_X1 us20_U273 (.ZN( us20_n540 ) , .A( us20_n763 ) , .B2( us20_n779 ) , .B1( us20_n817 ) );
  AOI21_X1 us20_U274 (.B1( us20_n699 ) , .ZN( us20_n700 ) , .A( us20_n732 ) , .B2( us20_n763 ) );
  AOI21_X1 us20_U275 (.ZN( us20_n591 ) , .B2( us20_n763 ) , .A( us20_n785 ) , .B1( us20_n812 ) );
  AOI21_X1 us20_U276 (.A( us20_n812 ) , .B2( us20_n813 ) , .B1( us20_n814 ) , .ZN( us20_n819 ) );
  INV_X1 us20_U277 (.A( us20_n791 ) , .ZN( us20_n873 ) );
  NOR2_X1 us20_U278 (.ZN( us20_n547 ) , .A1( us20_n699 ) , .A2( us20_n744 ) );
  INV_X1 us20_U279 (.A( us20_n729 ) , .ZN( us20_n868 ) );
  NOR4_X1 us20_U28 (.A4( us20_n514 ) , .A3( us20_n515 ) , .A2( us20_n516 ) , .A1( us20_n517 ) , .ZN( us20_n524 ) );
  AOI21_X1 us20_U280 (.ZN( us20_n569 ) , .B1( us20_n750 ) , .B2( us20_n762 ) , .A( us20_n780 ) );
  AOI21_X1 us20_U281 (.ZN( us20_n649 ) , .B1( us20_n729 ) , .B2( us20_n763 ) , .A( us20_n813 ) );
  NOR2_X1 us20_U282 (.ZN( us20_n685 ) , .A1( us20_n729 ) , .A2( us20_n816 ) );
  AOI21_X1 us20_U283 (.B1( us20_n686 ) , .ZN( us20_n687 ) , .A( us20_n728 ) , .B2( us20_n761 ) );
  AOI21_X1 us20_U284 (.ZN( us20_n640 ) , .B2( us20_n747 ) , .A( us20_n792 ) , .B1( us20_n803 ) );
  NOR2_X1 us20_U285 (.ZN( us20_n568 ) , .A1( us20_n729 ) , .A2( us20_n762 ) );
  AOI21_X1 us20_U286 (.ZN( us20_n593 ) , .B1( us20_n750 ) , .A( us20_n792 ) , .B2( us20_n813 ) );
  AOI21_X1 us20_U287 (.ZN( us20_n514 ) , .A( us20_n779 ) , .B2( us20_n792 ) , .B1( us20_n812 ) );
  INV_X1 us20_U288 (.A( us20_n699 ) , .ZN( us20_n853 ) );
  AOI21_X1 us20_U289 (.ZN( us20_n450 ) , .B2( us20_n792 ) , .A( us20_n803 ) , .B1( us20_n815 ) );
  AOI222_X1 us20_U29 (.ZN( us20_n525 ) , .A1( us20_n834 ) , .B2( us20_n837 ) , .C1( us20_n844 ) , .C2( us20_n850 ) , .A2( us20_n852 ) , .B1( us20_n866 ) );
  AOI21_X1 us20_U290 (.ZN( us20_n639 ) , .B2( us20_n749 ) , .A( us20_n788 ) , .B1( us20_n812 ) );
  AOI21_X1 us20_U291 (.ZN( us20_n564 ) , .B1( us20_n724 ) , .A( us20_n779 ) , .B2( us20_n791 ) );
  AOI21_X1 us20_U292 (.ZN( us20_n689 ) , .B2( us20_n749 ) , .B1( us20_n763 ) , .A( us20_n806 ) );
  NOR2_X1 us20_U293 (.ZN( us20_n529 ) , .A1( us20_n708 ) , .A2( us20_n779 ) );
  NOR2_X1 us20_U294 (.ZN( us20_n567 ) , .A1( us20_n747 ) , .A2( us20_n805 ) );
  AOI21_X1 us20_U295 (.A( us20_n790 ) , .B2( us20_n791 ) , .B1( us20_n792 ) , .ZN( us20_n793 ) );
  AOI21_X1 us20_U296 (.A( us20_n733 ) , .ZN( us20_n734 ) , .B2( us20_n780 ) , .B1( us20_n792 ) );
  NOR2_X1 us20_U297 (.A2( us20_n813 ) , .A1( us20_n815 ) , .ZN( us20_n821 ) );
  AOI21_X1 us20_U298 (.ZN( us20_n641 ) , .B1( us20_n680 ) , .A( us20_n791 ) , .B2( us20_n817 ) );
  NOR2_X1 us20_U299 (.ZN( us20_n578 ) , .A1( us20_n708 ) , .A2( us20_n813 ) );
  NAND4_X1 us20_U3 (.ZN( sa22_sr_2 ) , .A4( us20_n643 ) , .A3( us20_n644 ) , .A2( us20_n645 ) , .A1( us20_n646 ) );
  NOR4_X1 us20_U30 (.A3( us20_n521 ) , .A1( us20_n522 ) , .ZN( us20_n523 ) , .A2( us20_n673 ) , .A4( us20_n769 ) );
  NOR2_X1 us20_U300 (.ZN( us20_n665 ) , .A1( us20_n780 ) , .A2( us20_n813 ) );
  NOR2_X1 us20_U301 (.ZN( us20_n711 ) , .A1( us20_n762 ) , .A2( us20_n763 ) );
  NOR2_X1 us20_U302 (.ZN( us20_n583 ) , .A1( us20_n792 ) , .A2( us20_n817 ) );
  NOR2_X1 us20_U303 (.ZN( us20_n682 ) , .A2( us20_n708 ) , .A1( us20_n817 ) );
  NOR2_X1 us20_U304 (.ZN( us20_n534 ) , .A1( us20_n724 ) , .A2( us20_n788 ) );
  NOR2_X1 us20_U305 (.ZN( us20_n684 ) , .A1( us20_n791 ) , .A2( us20_n813 ) );
  NAND2_X1 us20_U306 (.ZN( us20_n753 ) , .A1( us20_n763 ) , .A2( us20_n805 ) );
  INV_X1 us20_U307 (.A( us20_n815 ) , .ZN( us20_n855 ) );
  AOI21_X1 us20_U308 (.ZN( us20_n442 ) , .A( us20_n699 ) , .B1( us20_n733 ) , .B2( us20_n750 ) );
  OAI21_X1 us20_U309 (.A( us20_n731 ) , .B1( us20_n732 ) , .ZN( us20_n736 ) , .B2( us20_n805 ) );
  AOI221_X1 us20_U31 (.A( us20_n781 ) , .ZN( us20_n798 ) , .C2( us20_n837 ) , .B2( us20_n838 ) , .B1( us20_n865 ) , .C1( us20_n866 ) );
  OAI21_X1 us20_U310 (.ZN( us20_n731 ) , .A( us20_n833 ) , .B2( us20_n852 ) , .B1( us20_n873 ) );
  INV_X1 us20_U311 (.A( us20_n780 ) , .ZN( us20_n850 ) );
  AOI21_X1 us20_U312 (.ZN( us20_n443 ) , .B1( us20_n789 ) , .B2( us20_n791 ) , .A( us20_n814 ) );
  NAND2_X1 us20_U313 (.ZN( us20_n714 ) , .A1( us20_n728 ) , .A2( us20_n780 ) );
  NAND2_X1 us20_U314 (.A2( us20_n762 ) , .A1( us20_n806 ) , .ZN( us20_n810 ) );
  INV_X1 us20_U315 (.A( us20_n785 ) , .ZN( us20_n846 ) );
  NOR2_X1 us20_U316 (.ZN( us20_n484 ) , .A1( us20_n788 ) , .A2( us20_n805 ) );
  AOI21_X1 us20_U317 (.ZN( us20_n497 ) , .A( us20_n779 ) , .B2( us20_n791 ) , .B1( us20_n804 ) );
  NOR2_X1 us20_U318 (.ZN( us20_n470 ) , .A2( us20_n779 ) , .A1( us20_n815 ) );
  NOR2_X1 us20_U319 (.ZN( us20_n712 ) , .A2( us20_n724 ) , .A1( us20_n790 ) );
  NOR4_X1 us20_U32 (.A4( us20_n793 ) , .A3( us20_n794 ) , .A2( us20_n795 ) , .A1( us20_n796 ) , .ZN( us20_n797 ) );
  NOR2_X1 us20_U320 (.ZN( us20_n526 ) , .A1( us20_n724 ) , .A2( us20_n750 ) );
  OAI21_X1 us20_U321 (.A( us20_n787 ) , .B2( us20_n788 ) , .B1( us20_n789 ) , .ZN( us20_n795 ) );
  OAI21_X1 us20_U322 (.ZN( us20_n787 ) , .A( us20_n839 ) , .B1( us20_n863 ) , .B2( us20_n873 ) );
  NAND2_X1 us20_U323 (.A1( us20_n699 ) , .A2( us20_n729 ) , .ZN( us20_n782 ) );
  NOR2_X1 us20_U324 (.ZN( us20_n518 ) , .A1( us20_n708 ) , .A2( us20_n788 ) );
  INV_X1 us20_U325 (.A( us20_n813 ) , .ZN( us20_n836 ) );
  NAND2_X1 us20_U326 (.ZN( us20_n671 ) , .A1( us20_n806 ) , .A2( us20_n816 ) );
  OAI21_X1 us20_U327 (.A( us20_n698 ) , .ZN( us20_n702 ) , .B2( us20_n750 ) , .B1( us20_n804 ) );
  OAI21_X1 us20_U328 (.ZN( us20_n698 ) , .B2( us20_n833 ) , .B1( us20_n838 ) , .A( us20_n860 ) );
  INV_X1 us20_U329 (.A( us20_n724 ) , .ZN( us20_n856 ) );
  NOR4_X1 us20_U33 (.A4( us20_n776 ) , .A3( us20_n777 ) , .A1( us20_n778 ) , .ZN( us20_n799 ) , .A2( us20_n801 ) );
  INV_X1 us20_U330 (.A( us20_n817 ) , .ZN( us20_n844 ) );
  AND2_X1 us20_U331 (.ZN( us20_n732 ) , .A1( us20_n779 ) , .A2( us20_n785 ) );
  OAI222_X1 us20_U332 (.ZN( us20_n617 ) , .B1( us20_n697 ) , .C1( us20_n724 ) , .C2( us20_n747 ) , .B2( us20_n786 ) , .A2( us20_n792 ) , .A1( us20_n816 ) );
  AOI221_X1 us20_U333 (.A( us20_n764 ) , .ZN( us20_n774 ) , .C2( us20_n810 ) , .B2( us20_n835 ) , .C1( us20_n855 ) , .B1( us20_n866 ) );
  AOI21_X1 us20_U334 (.B2( us20_n763 ) , .ZN( us20_n764 ) , .A( us20_n788 ) , .B1( us20_n792 ) );
  INV_X1 us20_U335 (.A( us20_n761 ) , .ZN( us20_n835 ) );
  NAND2_X1 us20_U336 (.A1( us20_n451 ) , .A2( us20_n454 ) , .ZN( us20_n814 ) );
  NAND2_X1 us20_U337 (.A1( us20_n447 ) , .A2( us20_n449 ) , .ZN( us20_n805 ) );
  NAND2_X1 us20_U338 (.A1( us20_n455 ) , .A2( us20_n462 ) , .ZN( us20_n750 ) );
  NAND2_X1 us20_U339 (.A1( us20_n455 ) , .A2( us20_n471 ) , .ZN( us20_n803 ) );
  NOR4_X1 us20_U34 (.A4( us20_n734 ) , .A3( us20_n735 ) , .A2( us20_n736 ) , .A1( us20_n737 ) , .ZN( us20_n738 ) );
  NAND2_X1 us20_U340 (.A1( us20_n453 ) , .A2( us20_n461 ) , .ZN( us20_n744 ) );
  NAND2_X1 us20_U341 (.A1( us20_n452 ) , .A2( us20_n465 ) , .ZN( us20_n669 ) );
  NAND2_X1 us20_U342 (.A2( us20_n448 ) , .A1( us20_n460 ) , .ZN( us20_n728 ) );
  NAND2_X1 us20_U343 (.A2( us20_n453 ) , .A1( us20_n455 ) , .ZN( us20_n806 ) );
  NAND2_X1 us20_U344 (.A1( us20_n451 ) , .A2( us20_n471 ) , .ZN( us20_n816 ) );
  NAND2_X1 us20_U345 (.A1( us20_n453 ) , .A2( us20_n472 ) , .ZN( us20_n785 ) );
  NAND2_X1 us20_U346 (.A2( us20_n454 ) , .A1( us20_n472 ) , .ZN( us20_n779 ) );
  NAND2_X1 us20_U347 (.A2( us20_n464 ) , .A1( us20_n465 ) , .ZN( us20_n812 ) );
  NAND2_X1 us20_U348 (.A1( us20_n441 ) , .A2( us20_n460 ) , .ZN( us20_n699 ) );
  NAND2_X1 us20_U349 (.A2( us20_n449 ) , .A1( us20_n452 ) , .ZN( us20_n763 ) );
  AOI211_X1 us20_U35 (.B( us20_n725 ) , .A( us20_n726 ) , .ZN( us20_n739 ) , .C1( us20_n843 ) , .C2( us20_n855 ) );
  NAND2_X1 us20_U350 (.A2( us20_n448 ) , .A1( us20_n452 ) , .ZN( us20_n729 ) );
  NAND2_X1 us20_U351 (.A2( us20_n461 ) , .A1( us20_n462 ) , .ZN( us20_n747 ) );
  NAND2_X1 us20_U352 (.A1( us20_n462 ) , .A2( us20_n472 ) , .ZN( us20_n788 ) );
  NOR2_X1 us20_U353 (.ZN( us20_n465 ) , .A2( us20_n847 ) , .A1( us20_n848 ) );
  NOR2_X1 us20_U354 (.ZN( us20_n453 ) , .A1( us20_n826 ) , .A2( us20_n827 ) );
  NOR2_X1 us20_U355 (.ZN( us20_n451 ) , .A1( us20_n828 ) , .A2( us20_n829 ) );
  NAND2_X1 us20_U356 (.A2( us20_n461 ) , .A1( us20_n471 ) , .ZN( us20_n697 ) );
  NAND2_X1 us20_U357 (.A1( us20_n451 ) , .A2( us20_n462 ) , .ZN( us20_n790 ) );
  NAND2_X1 us20_U358 (.A2( us20_n441 ) , .A1( us20_n447 ) , .ZN( us20_n784 ) );
  NAND2_X2 us20_U359 (.A2( us20_n448 ) , .A1( us20_n464 ) , .ZN( us20_n815 ) );
  NOR3_X1 us20_U36 (.A3( us20_n722 ) , .A1( us20_n723 ) , .ZN( us20_n740 ) , .A2( us20_n741 ) );
  NAND2_X1 us20_U360 (.A2( us20_n454 ) , .A1( us20_n455 ) , .ZN( us20_n730 ) );
  NAND2_X2 us20_U361 (.A2( us20_n441 ) , .A1( us20_n452 ) , .ZN( us20_n791 ) );
  NAND2_X2 us20_U362 (.A1( us20_n449 ) , .A2( us20_n464 ) , .ZN( us20_n724 ) );
  NAND2_X2 us20_U363 (.A1( us20_n449 ) , .A2( us20_n460 ) , .ZN( us20_n792 ) );
  NAND2_X2 us20_U364 (.A1( us20_n441 ) , .A2( us20_n464 ) , .ZN( us20_n708 ) );
  NAND2_X2 us20_U365 (.A2( us20_n471 ) , .A1( us20_n472 ) , .ZN( us20_n817 ) );
  NAND2_X2 us20_U366 (.A2( us20_n460 ) , .A1( us20_n465 ) , .ZN( us20_n780 ) );
  NOR2_X1 us20_U367 (.ZN( us20_n447 ) , .A2( us20_n849 ) , .A1( us20_n858 ) );
  NAND2_X1 us20_U368 (.A1( us20_n447 ) , .A2( us20_n448 ) , .ZN( us20_n786 ) );
  NOR2_X1 us20_U369 (.A2( sa20_6 ) , .A1( sa20_7 ) , .ZN( us20_n464 ) );
  NOR4_X1 us20_U37 (.A3( us20_n755 ) , .A2( us20_n756 ) , .A1( us20_n757 ) , .ZN( us20_n758 ) , .A4( us20_n869 ) );
  NOR2_X1 us20_U370 (.A2( sa20_7 ) , .ZN( us20_n460 ) , .A1( us20_n849 ) );
  NOR2_X1 us20_U371 (.A2( sa20_4 ) , .ZN( us20_n449 ) , .A1( us20_n848 ) );
  NOR2_X1 us20_U372 (.A2( sa20_4 ) , .A1( sa20_5 ) , .ZN( us20_n441 ) );
  NOR2_X1 us20_U373 (.A2( sa20_5 ) , .ZN( us20_n448 ) , .A1( us20_n847 ) );
  NOR2_X1 us20_U374 (.A2( sa20_1 ) , .ZN( us20_n471 ) , .A1( us20_n826 ) );
  NOR2_X1 us20_U375 (.A2( sa20_2 ) , .A1( sa20_3 ) , .ZN( us20_n472 ) );
  NOR2_X1 us20_U376 (.A2( sa20_6 ) , .ZN( us20_n452 ) , .A1( us20_n858 ) );
  NOR2_X1 us20_U377 (.A2( sa20_0 ) , .A1( sa20_1 ) , .ZN( us20_n462 ) );
  NOR2_X1 us20_U378 (.A2( sa20_3 ) , .ZN( us20_n455 ) , .A1( us20_n828 ) );
  NOR2_X1 us20_U379 (.A2( sa20_2 ) , .ZN( us20_n461 ) , .A1( us20_n829 ) );
  AOI211_X1 us20_U38 (.B( us20_n745 ) , .A( us20_n746 ) , .ZN( us20_n759 ) , .C1( us20_n832 ) , .C2( us20_n853 ) );
  NOR2_X1 us20_U380 (.A2( sa20_0 ) , .ZN( us20_n454 ) , .A1( us20_n827 ) );
  INV_X1 us20_U381 (.A( sa20_4 ) , .ZN( us20_n847 ) );
  INV_X1 us20_U382 (.A( sa20_6 ) , .ZN( us20_n849 ) );
  INV_X1 us20_U383 (.A( sa20_3 ) , .ZN( us20_n829 ) );
  INV_X1 us20_U384 (.A( sa20_1 ) , .ZN( us20_n827 ) );
  INV_X1 us20_U385 (.A( sa20_2 ) , .ZN( us20_n828 ) );
  INV_X1 us20_U386 (.A( sa20_0 ) , .ZN( us20_n826 ) );
  INV_X1 us20_U387 (.A( sa20_5 ) , .ZN( us20_n848 ) );
  INV_X1 us20_U388 (.A( sa20_7 ) , .ZN( us20_n858 ) );
  NAND2_X1 us20_U389 (.A1( us20_n729 ) , .A2( us20_n784 ) , .ZN( us20_n811 ) );
  NOR3_X1 us20_U39 (.A3( us20_n741 ) , .A2( us20_n742 ) , .A1( us20_n743 ) , .ZN( us20_n760 ) );
  OAI22_X1 us20_U390 (.ZN( us20_n588 ) , .A2( us20_n747 ) , .B2( us20_n762 ) , .A1( us20_n763 ) , .B1( us20_n784 ) );
  AOI21_X1 us20_U391 (.ZN( us20_n592 ) , .B1( us20_n728 ) , .B2( us20_n784 ) , .A( us20_n790 ) );
  AOI21_X1 us20_U392 (.ZN( us20_n648 ) , .A( us20_n762 ) , .B2( us20_n784 ) , .B1( us20_n792 ) );
  AOI21_X1 us20_U393 (.ZN( us20_n623 ) , .B1( us20_n699 ) , .A( us20_n779 ) , .B2( us20_n784 ) );
  OAI22_X1 us20_U394 (.ZN( us20_n681 ) , .A1( us20_n699 ) , .A2( us20_n730 ) , .B2( us20_n784 ) , .B1( us20_n817 ) );
  OAI21_X1 us20_U395 (.A( us20_n613 ) , .ZN( us20_n616 ) , .B1( us20_n625 ) , .B2( us20_n784 ) );
  NOR2_X1 us20_U396 (.ZN( us20_n610 ) , .A1( us20_n784 ) , .A2( us20_n816 ) );
  OAI222_X1 us20_U397 (.A2( us20_n669 ) , .ZN( us20_n674 ) , .B1( us20_n747 ) , .B2( us20_n784 ) , .C2( us20_n788 ) , .C1( us20_n815 ) , .A1( us20_n817 ) );
  NOR2_X1 us20_U398 (.ZN( us20_n651 ) , .A1( us20_n784 ) , .A2( us20_n788 ) );
  NOR2_X1 us20_U399 (.ZN( us20_n553 ) , .A2( us20_n744 ) , .A1( us20_n784 ) );
  NOR3_X1 us20_U4 (.ZN( us20_n598 ) , .A1( us20_n608 ) , .A3( us20_n723 ) , .A2( us20_n742 ) );
  NOR2_X1 us20_U40 (.ZN( us20_n804 ) , .A1( us20_n854 ) , .A2( us20_n861 ) );
  INV_X1 us20_U400 (.A( us20_n784 ) , .ZN( us20_n861 ) );
  INV_X1 us20_U401 (.A( us20_n697 ) , .ZN( us20_n838 ) );
  NOR2_X1 us20_U402 (.A1( us20_n697 ) , .ZN( us20_n770 ) , .A2( us20_n815 ) );
  AOI21_X1 us20_U403 (.ZN( us20_n571 ) , .B2( us20_n697 ) , .B1( us20_n806 ) , .A( us20_n812 ) );
  NOR2_X1 us20_U404 (.ZN( us20_n632 ) , .A2( us20_n697 ) , .A1( us20_n724 ) );
  AOI21_X1 us20_U405 (.ZN( us20_n478 ) , .B2( us20_n697 ) , .A( us20_n749 ) , .B1( us20_n779 ) );
  NOR2_X1 us20_U406 (.ZN( us20_n662 ) , .A2( us20_n697 ) , .A1( us20_n729 ) );
  NOR2_X1 us20_U407 (.A2( us20_n697 ) , .A1( us20_n780 ) , .ZN( us20_n820 ) );
  NOR2_X1 us20_U408 (.ZN( us20_n600 ) , .A2( us20_n697 ) , .A1( us20_n784 ) );
  NOR2_X1 us20_U409 (.A2( us20_n697 ) , .ZN( us20_n716 ) , .A1( us20_n792 ) );
  NAND4_X1 us20_U41 (.ZN( sa22_sr_3 ) , .A4( us20_n704 ) , .A3( us20_n705 ) , .A2( us20_n706 ) , .A1( us20_n707 ) );
  NOR2_X1 us20_U410 (.ZN( us20_n566 ) , .A2( us20_n697 ) , .A1( us20_n763 ) );
  NOR2_X1 us20_U411 (.ZN( us20_n594 ) , .A2( us20_n697 ) , .A1( us20_n728 ) );
  AOI21_X1 us20_U412 (.ZN( us20_n552 ) , .B1( us20_n669 ) , .A( us20_n697 ) , .B2( us20_n805 ) );
  NOR2_X1 us20_U413 (.ZN( us20_n541 ) , .A2( us20_n697 ) , .A1( us20_n699 ) );
  NOR2_X1 us20_U414 (.ZN( us20_n580 ) , .A2( us20_n697 ) , .A1( us20_n791 ) );
  NAND2_X1 us20_U415 (.A1( us20_n454 ) , .A2( us20_n461 ) , .ZN( us20_n813 ) );
  AND2_X1 us20_U416 (.ZN( us20_n438 ) , .A2( us20_n831 ) , .A1( us20_n854 ) );
  AND2_X1 us20_U417 (.ZN( us20_n439 ) , .A2( us20_n843 ) , .A1( us20_n861 ) );
  NOR3_X1 us20_U418 (.A1( us20_n438 ) , .A2( us20_n439 ) , .A3( us20_n576 ) , .ZN( us20_n587 ) );
  INV_X1 us20_U419 (.A( us20_n812 ) , .ZN( us20_n854 ) );
  NOR4_X1 us20_U42 (.A4( us20_n700 ) , .A3( us20_n701 ) , .A2( us20_n702 ) , .A1( us20_n703 ) , .ZN( us20_n704 ) );
  INV_X1 us20_U420 (.A( us20_n816 ) , .ZN( us20_n831 ) );
  INV_X1 us20_U421 (.A( us20_n803 ) , .ZN( us20_n843 ) );
  AOI21_X1 us20_U422 (.ZN( us20_n576 ) , .B2( us20_n724 ) , .B1( us20_n748 ) , .A( us20_n785 ) );
  OAI221_X1 us20_U423 (.A( us20_n783 ) , .C2( us20_n784 ) , .B2( us20_n785 ) , .B1( us20_n786 ) , .ZN( us20_n796 ) , .C1( us20_n813 ) );
  AOI21_X1 us20_U424 (.ZN( us20_n500 ) , .A( us20_n697 ) , .B1( us20_n708 ) , .B2( us20_n786 ) );
  OAI221_X1 us20_U425 (.A( us20_n696 ) , .ZN( us20_n703 ) , .C2( us20_n784 ) , .C1( us20_n785 ) , .B1( us20_n786 ) , .B2( us20_n806 ) );
  OAI22_X1 us20_U426 (.ZN( us20_n590 ) , .B1( us20_n730 ) , .B2( us20_n749 ) , .A2( us20_n786 ) , .A1( us20_n803 ) );
  AOI222_X1 us20_U427 (.ZN( us20_n605 ) , .B2( us20_n671 ) , .B1( us20_n753 ) , .C2( us20_n831 ) , .A1( us20_n833 ) , .A2( us20_n862 ) , .C1( us20_n863 ) );
  AOI222_X1 us20_U428 (.ZN( us20_n513 ) , .C1( us20_n832 ) , .B2( us20_n837 ) , .A2( us20_n843 ) , .C2( us20_n862 ) , .B1( us20_n863 ) , .A1( us20_n866 ) );
  AOI221_X1 us20_U429 (.A( us20_n483 ) , .ZN( us20_n488 ) , .B1( us20_n831 ) , .C2( us20_n844 ) , .C1( us20_n852 ) , .B2( us20_n862 ) );
  AOI211_X1 us20_U43 (.B( us20_n694 ) , .A( us20_n695 ) , .ZN( us20_n705 ) , .C2( us20_n831 ) , .C1( us20_n851 ) );
  NAND2_X1 us20_U430 (.A2( us20_n749 ) , .A1( us20_n786 ) , .ZN( us20_n809 ) );
  NOR2_X1 us20_U431 (.ZN( us20_n612 ) , .A1( us20_n779 ) , .A2( us20_n786 ) );
  NOR2_X1 us20_U432 (.ZN( us20_n717 ) , .A2( us20_n744 ) , .A1( us20_n786 ) );
  NOR2_X1 us20_U433 (.ZN( us20_n653 ) , .A1( us20_n762 ) , .A2( us20_n786 ) );
  NOR2_X1 us20_U434 (.ZN( us20_n554 ) , .A1( us20_n786 ) , .A2( us20_n813 ) );
  NOR2_X1 us20_U435 (.ZN( us20_n789 ) , .A2( us20_n862 ) , .A1( us20_n868 ) );
  NOR2_X1 us20_U436 (.ZN( us20_n701 ) , .A2( us20_n786 ) , .A1( us20_n817 ) );
  NAND3_X1 us20_U437 (.ZN( sa22_sr_6 ) , .A3( us20_n797 ) , .A2( us20_n798 ) , .A1( us20_n799 ) );
  NAND3_X1 us20_U438 (.ZN( sa22_sr_5 ) , .A3( us20_n758 ) , .A2( us20_n759 ) , .A1( us20_n760 ) );
  NAND3_X1 us20_U439 (.ZN( sa22_sr_4 ) , .A3( us20_n738 ) , .A2( us20_n739 ) , .A1( us20_n740 ) );
  NOR2_X1 us20_U44 (.ZN( us20_n707 ) , .A2( us20_n776 ) , .A1( us20_n800 ) );
  NAND3_X1 us20_U440 (.A3( us20_n675 ) , .A2( us20_n676 ) , .A1( us20_n677 ) , .ZN( us20_n807 ) );
  NAND3_X1 us20_U441 (.ZN( us20_n638 ) , .A3( us20_n708 ) , .A2( us20_n724 ) , .A1( us20_n792 ) );
  NAND3_X1 us20_U442 (.A3( us20_n618 ) , .A2( us20_n619 ) , .A1( us20_n620 ) , .ZN( us20_n725 ) );
  NAND3_X1 us20_U443 (.A3( us20_n585 ) , .A2( us20_n586 ) , .A1( us20_n587 ) , .ZN( us20_n621 ) );
  NAND3_X1 us20_U444 (.ZN( us20_n565 ) , .A3( us20_n680 ) , .A2( us20_n750 ) , .A1( us20_n785 ) );
  NAND3_X1 us20_U445 (.A3( us20_n523 ) , .A2( us20_n524 ) , .A1( us20_n525 ) , .ZN( us20_n742 ) );
  NAND3_X1 us20_U446 (.A3( us20_n512 ) , .A1( us20_n513 ) , .ZN( us20_n608 ) , .A2( us20_n871 ) );
  NAND3_X1 us20_U447 (.A3( us20_n467 ) , .A2( us20_n468 ) , .A1( us20_n469 ) , .ZN( us20_n777 ) );
  NOR2_X1 us20_U448 (.A1( us20_n730 ) , .ZN( us20_n765 ) , .A2( us20_n786 ) );
  INV_X1 us20_U449 (.A( us20_n786 ) , .ZN( us20_n862 ) );
  NAND4_X1 us20_U45 (.ZN( sa22_sr_7 ) , .A4( us20_n822 ) , .A3( us20_n823 ) , .A2( us20_n824 ) , .A1( us20_n825 ) );
  NOR4_X1 us20_U46 (.A4( us20_n818 ) , .A3( us20_n819 ) , .A2( us20_n820 ) , .A1( us20_n821 ) , .ZN( us20_n822 ) );
  AOI222_X1 us20_U47 (.C2( us20_n809 ) , .B2( us20_n810 ) , .A2( us20_n811 ) , .ZN( us20_n823 ) , .C1( us20_n832 ) , .A1( us20_n839 ) , .B1( us20_n853 ) );
  AOI211_X1 us20_U48 (.B( us20_n807 ) , .A( us20_n808 ) , .ZN( us20_n824 ) , .C1( us20_n842 ) , .C2( us20_n850 ) );
  NAND4_X1 us20_U49 (.ZN( sa22_sr_0 ) , .A4( us20_n501 ) , .A3( us20_n502 ) , .A2( us20_n503 ) , .A1( us20_n504 ) );
  NOR3_X1 us20_U5 (.A3( us20_n800 ) , .A2( us20_n801 ) , .A1( us20_n802 ) , .ZN( us20_n825 ) );
  NOR4_X1 us20_U50 (.A4( us20_n498 ) , .A3( us20_n499 ) , .A2( us20_n500 ) , .ZN( us20_n501 ) , .A1( us20_n527 ) );
  AOI221_X1 us20_U51 (.A( us20_n497 ) , .ZN( us20_n502 ) , .B2( us20_n843 ) , .C1( us20_n846 ) , .C2( us20_n860 ) , .B1( us20_n862 ) );
  AOI211_X1 us20_U52 (.A( us20_n496 ) , .ZN( us20_n503 ) , .B( us20_n802 ) , .C2( us20_n839 ) , .C1( us20_n851 ) );
  NAND4_X1 us20_U53 (.ZN( sa22_sr_1 ) , .A4( us20_n595 ) , .A3( us20_n596 ) , .A2( us20_n597 ) , .A1( us20_n598 ) );
  NOR4_X1 us20_U54 (.A4( us20_n591 ) , .A3( us20_n592 ) , .A2( us20_n593 ) , .A1( us20_n594 ) , .ZN( us20_n595 ) );
  AOI211_X1 us20_U55 (.B( us20_n589 ) , .A( us20_n590 ) , .ZN( us20_n596 ) , .C2( us20_n811 ) , .C1( us20_n833 ) );
  AOI211_X1 us20_U56 (.A( us20_n588 ) , .ZN( us20_n597 ) , .B( us20_n621 ) , .C1( us20_n845 ) , .C2( us20_n855 ) );
  NOR2_X1 us20_U57 (.ZN( us20_n748 ) , .A1( us20_n861 ) , .A2( us20_n862 ) );
  NOR2_X1 us20_U58 (.ZN( us20_n625 ) , .A2( us20_n836 ) , .A1( us20_n839 ) );
  AOI222_X1 us20_U59 (.B2( us20_n638 ) , .ZN( us20_n644 ) , .B1( us20_n841 ) , .A1( us20_n842 ) , .C2( us20_n846 ) , .C1( us20_n863 ) , .A2( us20_n865 ) );
  NOR3_X1 us20_U6 (.A3( us20_n621 ) , .A2( us20_n622 ) , .ZN( us20_n636 ) , .A1( us20_n725 ) );
  NOR4_X1 us20_U60 (.A4( us20_n639 ) , .A3( us20_n640 ) , .A2( us20_n641 ) , .A1( us20_n642 ) , .ZN( us20_n643 ) );
  NOR3_X1 us20_U61 (.A2( us20_n607 ) , .A1( us20_n608 ) , .ZN( us20_n646 ) , .A3( us20_n722 ) );
  NAND4_X1 us20_U62 (.A4( us20_n603 ) , .A3( us20_n604 ) , .A2( us20_n605 ) , .A1( us20_n606 ) , .ZN( us20_n722 ) );
  NOR3_X1 us20_U63 (.A1( us20_n599 ) , .ZN( us20_n604 ) , .A3( us20_n663 ) , .A2( us20_n770 ) );
  NOR4_X1 us20_U64 (.A3( us20_n600 ) , .A2( us20_n601 ) , .A1( us20_n602 ) , .ZN( us20_n603 ) , .A4( us20_n655 ) );
  AOI222_X1 us20_U65 (.ZN( us20_n606 ) , .A1( us20_n830 ) , .C2( us20_n837 ) , .B1( us20_n842 ) , .A2( us20_n856 ) , .B2( us20_n861 ) , .C1( us20_n868 ) );
  AOI222_X1 us20_U66 (.ZN( us20_n469 ) , .B1( us20_n832 ) , .A1( us20_n839 ) , .C1( us20_n842 ) , .C2( us20_n851 ) , .A2( us20_n855 ) , .B2( us20_n865 ) );
  NOR4_X1 us20_U67 (.A1( us20_n466 ) , .ZN( us20_n467 ) , .A4( us20_n542 ) , .A2( us20_n554 ) , .A3( us20_n614 ) );
  AOI221_X1 us20_U68 (.ZN( us20_n468 ) , .C2( us20_n714 ) , .B2( us20_n831 ) , .C1( us20_n845 ) , .B1( us20_n860 ) , .A( us20_n864 ) );
  NAND4_X1 us20_U69 (.A4( us20_n485 ) , .A3( us20_n486 ) , .A2( us20_n487 ) , .A1( us20_n488 ) , .ZN( us20_n778 ) );
  NOR2_X1 us20_U7 (.ZN( us20_n495 ) , .A1( us20_n678 ) , .A2( us20_n694 ) );
  NOR4_X1 us20_U70 (.A4( us20_n484 ) , .ZN( us20_n487 ) , .A1( us20_n566 ) , .A2( us20_n581 ) , .A3( us20_n602 ) );
  NOR4_X1 us20_U71 (.ZN( us20_n486 ) , .A1( us20_n507 ) , .A2( us20_n519 ) , .A4( us20_n546 ) , .A3( us20_n611 ) );
  NOR4_X1 us20_U72 (.ZN( us20_n485 ) , .A2( us20_n533 ) , .A1( us20_n558 ) , .A3( us20_n631 ) , .A4( us20_n718 ) );
  NAND4_X1 us20_U73 (.A4( us20_n657 ) , .A3( us20_n658 ) , .A2( us20_n659 ) , .A1( us20_n660 ) , .ZN( us20_n800 ) );
  NOR3_X1 us20_U74 (.A3( us20_n648 ) , .A2( us20_n649 ) , .A1( us20_n650 ) , .ZN( us20_n659 ) );
  NOR3_X1 us20_U75 (.A3( us20_n651 ) , .A2( us20_n652 ) , .A1( us20_n653 ) , .ZN( us20_n658 ) );
  NOR3_X1 us20_U76 (.A3( us20_n654 ) , .A2( us20_n655 ) , .A1( us20_n656 ) , .ZN( us20_n657 ) );
  NAND4_X1 us20_U77 (.A4( us20_n560 ) , .A3( us20_n561 ) , .A2( us20_n562 ) , .A1( us20_n563 ) , .ZN( us20_n607 ) );
  NOR4_X1 us20_U78 (.A4( us20_n552 ) , .A3( us20_n553 ) , .A2( us20_n554 ) , .A1( us20_n555 ) , .ZN( us20_n562 ) );
  NOR4_X1 us20_U79 (.ZN( us20_n561 ) , .A1( us20_n653 ) , .A3( us20_n661 ) , .A4( us20_n685 ) , .A2( us20_n768 ) );
  NOR2_X1 us20_U8 (.A1( us20_n678 ) , .ZN( us20_n693 ) , .A2( us20_n807 ) );
  NOR4_X1 us20_U80 (.A4( us20_n556 ) , .A3( us20_n557 ) , .A2( us20_n558 ) , .A1( us20_n559 ) , .ZN( us20_n560 ) );
  NAND4_X1 us20_U81 (.A4( us20_n772 ) , .A3( us20_n773 ) , .A2( us20_n774 ) , .A1( us20_n775 ) , .ZN( us20_n801 ) );
  NOR3_X1 us20_U82 (.A3( us20_n765 ) , .A2( us20_n766 ) , .A1( us20_n767 ) , .ZN( us20_n773 ) );
  NOR4_X1 us20_U83 (.A4( us20_n768 ) , .A3( us20_n769 ) , .A2( us20_n770 ) , .A1( us20_n771 ) , .ZN( us20_n772 ) );
  AOI222_X1 us20_U84 (.ZN( us20_n775 ) , .A1( us20_n830 ) , .C1( us20_n834 ) , .B2( us20_n841 ) , .A2( us20_n850 ) , .B1( us20_n861 ) , .C2( us20_n873 ) );
  NOR4_X1 us20_U85 (.A4( us20_n509 ) , .A2( us20_n510 ) , .A1( us20_n511 ) , .ZN( us20_n512 ) , .A3( us20_n670 ) );
  INV_X1 us20_U86 (.A( us20_n505 ) , .ZN( us20_n871 ) );
  NOR4_X1 us20_U87 (.A4( us20_n661 ) , .A3( us20_n662 ) , .A2( us20_n663 ) , .A1( us20_n664 ) , .ZN( us20_n677 ) );
  NOR4_X1 us20_U88 (.A4( us20_n665 ) , .A3( us20_n666 ) , .A2( us20_n667 ) , .A1( us20_n668 ) , .ZN( us20_n676 ) );
  NOR4_X1 us20_U89 (.A3( us20_n673 ) , .A1( us20_n674 ) , .ZN( us20_n675 ) , .A4( us20_n715 ) , .A2( us20_n859 ) );
  NOR3_X1 us20_U9 (.ZN( us20_n504 ) , .A2( us20_n679 ) , .A3( us20_n777 ) , .A1( us20_n876 ) );
  NOR2_X1 us20_U90 (.ZN( us20_n761 ) , .A1( us20_n833 ) , .A2( us20_n834 ) );
  NOR2_X1 us20_U91 (.ZN( us20_n686 ) , .A1( us20_n831 ) , .A2( us20_n832 ) );
  NOR4_X1 us20_U92 (.A4( us20_n577 ) , .A3( us20_n578 ) , .A2( us20_n579 ) , .ZN( us20_n586 ) , .A1( us20_n683 ) );
  NOR4_X1 us20_U93 (.A1( us20_n584 ) , .ZN( us20_n585 ) , .A3( us20_n652 ) , .A2( us20_n662 ) , .A4( us20_n767 ) );
  NAND4_X1 us20_U94 (.A4( us20_n456 ) , .A3( us20_n457 ) , .A2( us20_n458 ) , .A1( us20_n459 ) , .ZN( us20_n679 ) );
  NOR3_X1 us20_U95 (.ZN( us20_n457 ) , .A3( us20_n530 ) , .A1( us20_n555 ) , .A2( us20_n570 ) );
  AOI221_X1 us20_U96 (.A( us20_n450 ) , .ZN( us20_n459 ) , .C2( us20_n753 ) , .B1( us20_n832 ) , .C1( us20_n842 ) , .B2( us20_n861 ) );
  NOR4_X1 us20_U97 (.ZN( us20_n458 ) , .A2( us20_n509 ) , .A1( us20_n599 ) , .A4( us20_n628 ) , .A3( us20_n711 ) );
  NAND4_X1 us20_U98 (.A4( us20_n535 ) , .A3( us20_n536 ) , .A2( us20_n537 ) , .A1( us20_n538 ) , .ZN( us20_n622 ) );
  NOR4_X1 us20_U99 (.A4( us20_n526 ) , .A2( us20_n527 ) , .A1( us20_n528 ) , .ZN( us20_n538 ) , .A3( us20_n701 ) );
  NOR2_X1 us33_U10 (.ZN( us33_n495 ) , .A1( us33_n678 ) , .A2( us33_n694 ) );
  NAND4_X1 us33_U100 (.A4( us33_n479 ) , .A3( us33_n480 ) , .A2( us33_n481 ) , .A1( us33_n482 ) , .ZN( us33_n694 ) );
  NOR3_X1 us33_U101 (.ZN( us33_n480 ) , .A2( us33_n508 ) , .A3( us33_n601 ) , .A1( us33_n610 ) );
  AOI211_X1 us33_U102 (.B( us33_n477 ) , .A( us33_n478 ) , .ZN( us33_n482 ) , .C2( us33_n833 ) , .C1( us33_n861 ) );
  NOR4_X1 us33_U103 (.ZN( us33_n481 ) , .A3( us33_n532 ) , .A4( us33_n545 ) , .A2( us33_n567 ) , .A1( us33_n717 ) );
  NAND4_X1 us33_U104 (.A4( us33_n548 ) , .A3( us33_n549 ) , .A2( us33_n550 ) , .A1( us33_n551 ) , .ZN( us33_n745 ) );
  NOR3_X1 us33_U105 (.ZN( us33_n549 ) , .A2( us33_n651 ) , .A1( us33_n667 ) , .A3( us33_n771 ) );
  AOI211_X1 us33_U106 (.B( us33_n539 ) , .A( us33_n540 ) , .ZN( us33_n551 ) , .C2( us33_n839 ) , .C1( us33_n851 ) );
  NOR4_X1 us33_U107 (.A4( us33_n544 ) , .A3( us33_n545 ) , .A2( us33_n546 ) , .A1( us33_n547 ) , .ZN( us33_n548 ) );
  NOR4_X1 us33_U108 (.ZN( us33_n620 ) , .A1( us33_n656 ) , .A3( us33_n666 ) , .A4( us33_n682 ) , .A2( us33_n766 ) );
  NOR4_X1 us33_U109 (.A4( us33_n609 ) , .A3( us33_n610 ) , .A2( us33_n611 ) , .A1( us33_n612 ) , .ZN( us33_n619 ) );
  NOR2_X1 us33_U11 (.A1( us33_n678 ) , .ZN( us33_n693 ) , .A2( us33_n807 ) );
  NOR4_X1 us33_U110 (.A4( us33_n614 ) , .A3( us33_n615 ) , .A2( us33_n616 ) , .A1( us33_n617 ) , .ZN( us33_n618 ) );
  NOR2_X1 us33_U111 (.ZN( us33_n686 ) , .A1( us33_n831 ) , .A2( us33_n832 ) );
  NAND4_X1 us33_U112 (.A4( us33_n485 ) , .A3( us33_n486 ) , .A2( us33_n487 ) , .A1( us33_n488 ) , .ZN( us33_n778 ) );
  NOR4_X1 us33_U113 (.A4( us33_n484 ) , .ZN( us33_n487 ) , .A1( us33_n566 ) , .A2( us33_n581 ) , .A3( us33_n602 ) );
  NOR4_X1 us33_U114 (.ZN( us33_n486 ) , .A1( us33_n507 ) , .A2( us33_n519 ) , .A4( us33_n546 ) , .A3( us33_n611 ) );
  NOR4_X1 us33_U115 (.ZN( us33_n485 ) , .A2( us33_n533 ) , .A1( us33_n558 ) , .A3( us33_n631 ) , .A4( us33_n718 ) );
  NAND4_X1 us33_U116 (.A4( us33_n691 ) , .A3( us33_n692 ) , .A1( us33_n693 ) , .ZN( us33_n776 ) , .A2( us33_n872 ) );
  AOI221_X1 us33_U117 (.A( us33_n681 ) , .ZN( us33_n692 ) , .B2( us33_n840 ) , .C1( us33_n842 ) , .C2( us33_n862 ) , .B1( us33_n865 ) );
  INV_X1 us33_U118 (.A( us33_n679 ) , .ZN( us33_n872 ) );
  NOR4_X1 us33_U119 (.A4( us33_n687 ) , .A3( us33_n688 ) , .A2( us33_n689 ) , .A1( us33_n690 ) , .ZN( us33_n691 ) );
  NOR3_X1 us33_U12 (.ZN( us33_n504 ) , .A2( us33_n679 ) , .A3( us33_n777 ) , .A1( us33_n876 ) );
  NAND4_X1 us33_U120 (.A4( us33_n719 ) , .A3( us33_n720 ) , .A2( us33_n721 ) , .ZN( us33_n741 ) , .A1( us33_n857 ) );
  INV_X1 us33_U121 (.A( us33_n709 ) , .ZN( us33_n857 ) );
  AOI221_X1 us33_U122 (.A( us33_n710 ) , .ZN( us33_n721 ) , .C2( us33_n844 ) , .B2( us33_n845 ) , .C1( us33_n861 ) , .B1( us33_n862 ) );
  NOR4_X1 us33_U123 (.A4( us33_n715 ) , .A3( us33_n716 ) , .A2( us33_n717 ) , .A1( us33_n718 ) , .ZN( us33_n719 ) );
  NAND4_X1 us33_U124 (.A4( us33_n473 ) , .A3( us33_n474 ) , .A2( us33_n475 ) , .A1( us33_n476 ) , .ZN( us33_n678 ) );
  NOR4_X1 us33_U125 (.ZN( us33_n475 ) , .A1( us33_n531 ) , .A3( us33_n568 ) , .A4( us33_n600 ) , .A2( us33_n642 ) );
  NOR4_X1 us33_U126 (.A4( us33_n470 ) , .ZN( us33_n476 ) , .A3( us33_n556 ) , .A1( us33_n735 ) , .A2( us33_n755 ) );
  NOR4_X1 us33_U127 (.ZN( us33_n474 ) , .A1( us33_n506 ) , .A3( us33_n544 ) , .A2( us33_n583 ) , .A4( us33_n716 ) );
  NOR2_X1 us33_U128 (.ZN( us33_n733 ) , .A2( us33_n832 ) , .A1( us33_n845 ) );
  NOR2_X1 us33_U129 (.ZN( us33_n789 ) , .A2( us33_n862 ) , .A1( us33_n868 ) );
  INV_X1 us33_U13 (.A( us33_n706 ) , .ZN( us33_n876 ) );
  NAND4_X1 us33_U130 (.A4( us33_n573 ) , .A3( us33_n574 ) , .A1( us33_n575 ) , .ZN( us33_n723 ) , .A2( us33_n874 ) );
  AOI221_X1 us33_U131 (.A( us33_n564 ) , .C2( us33_n565 ) , .ZN( us33_n574 ) , .B2( us33_n845 ) , .B1( us33_n852 ) , .C1( us33_n853 ) );
  NOR4_X1 us33_U132 (.A4( us33_n569 ) , .A3( us33_n570 ) , .A2( us33_n571 ) , .A1( us33_n572 ) , .ZN( us33_n573 ) );
  INV_X1 us33_U133 (.A( us33_n607 ) , .ZN( us33_n874 ) );
  NAND4_X1 us33_U134 (.A4( us33_n633 ) , .A3( us33_n634 ) , .A2( us33_n635 ) , .A1( us33_n636 ) , .ZN( us33_n743 ) );
  AOI211_X1 us33_U135 (.B( us33_n623 ) , .A( us33_n624 ) , .ZN( us33_n635 ) , .C2( us33_n836 ) , .C1( us33_n863 ) );
  NOR4_X1 us33_U136 (.A4( us33_n629 ) , .A3( us33_n630 ) , .A2( us33_n631 ) , .A1( us33_n632 ) , .ZN( us33_n633 ) );
  NOR4_X1 us33_U137 (.A4( us33_n626 ) , .A3( us33_n627 ) , .A2( us33_n628 ) , .ZN( us33_n634 ) , .A1( us33_n664 ) );
  NAND4_X1 us33_U138 (.A4( us33_n493 ) , .A3( us33_n494 ) , .A1( us33_n495 ) , .ZN( us33_n802 ) , .A2( us33_n867 ) );
  AOI221_X1 us33_U139 (.A( us33_n489 ) , .ZN( us33_n494 ) , .B2( us33_n836 ) , .C2( us33_n841 ) , .C1( us33_n851 ) , .B1( us33_n860 ) );
  INV_X1 us33_U14 (.A( us33_n680 ) , .ZN( us33_n840 ) );
  INV_X1 us33_U140 (.A( us33_n778 ) , .ZN( us33_n867 ) );
  NOR4_X1 us33_U141 (.A2( us33_n491 ) , .A1( us33_n492 ) , .ZN( us33_n493 ) , .A3( us33_n580 ) , .A4( us33_n612 ) );
  NOR4_X1 us33_U142 (.A4( us33_n734 ) , .A3( us33_n735 ) , .A2( us33_n736 ) , .A1( us33_n737 ) , .ZN( us33_n738 ) );
  AOI211_X1 us33_U143 (.B( us33_n725 ) , .A( us33_n726 ) , .ZN( us33_n739 ) , .C1( us33_n843 ) , .C2( us33_n855 ) );
  NOR3_X1 us33_U144 (.A3( us33_n722 ) , .A1( us33_n723 ) , .ZN( us33_n740 ) , .A2( us33_n741 ) );
  INV_X1 us33_U145 (.A( us33_n762 ) , .ZN( us33_n830 ) );
  OR4_X1 us33_U146 (.A4( us33_n566 ) , .A3( us33_n567 ) , .A2( us33_n568 ) , .ZN( us33_n572 ) , .A1( us33_n665 ) );
  OR4_X1 us33_U147 (.A4( us33_n682 ) , .A3( us33_n683 ) , .A2( us33_n684 ) , .A1( us33_n685 ) , .ZN( us33_n690 ) );
  OR4_X1 us33_U148 (.ZN( us33_n466 ) , .A4( us33_n518 ) , .A3( us33_n529 ) , .A2( us33_n578 ) , .A1( us33_n712 ) );
  OR4_X1 us33_U149 (.A4( us33_n518 ) , .A2( us33_n519 ) , .A1( us33_n520 ) , .ZN( us33_n522 ) , .A3( us33_n821 ) );
  NOR4_X1 us33_U15 (.A4( us33_n445 ) , .A3( us33_n446 ) , .A2( us33_n516 ) , .A1( us33_n541 ) , .ZN( us33_n706 ) );
  OR4_X1 us33_U150 (.ZN( us33_n492 ) , .A4( us33_n534 ) , .A2( us33_n547 ) , .A1( us33_n559 ) , .A3( us33_n632 ) );
  OR4_X1 us33_U151 (.A4( us33_n580 ) , .A3( us33_n581 ) , .A2( us33_n582 ) , .A1( us33_n583 ) , .ZN( us33_n584 ) );
  INV_X1 us33_U152 (.A( us33_n697 ) , .ZN( us33_n838 ) );
  NAND2_X1 us33_U153 (.ZN( us33_n613 ) , .A2( us33_n837 ) , .A1( us33_n873 ) );
  OR3_X1 us33_U154 (.A3( us33_n506 ) , .A2( us33_n507 ) , .A1( us33_n508 ) , .ZN( us33_n511 ) );
  INV_X1 us33_U155 (.A( us33_n754 ) , .ZN( us33_n869 ) );
  OAI21_X1 us33_U156 (.B1( us33_n753 ) , .ZN( us33_n754 ) , .A( us33_n845 ) , .B2( us33_n868 ) );
  INV_X1 us33_U157 (.A( us33_n463 ) , .ZN( us33_n864 ) );
  OAI21_X1 us33_U158 (.ZN( us33_n463 ) , .B1( us33_n809 ) , .A( us33_n834 ) , .B2( us33_n851 ) );
  INV_X1 us33_U159 (.A( us33_n672 ) , .ZN( us33_n859 ) );
  OR3_X1 us33_U16 (.ZN( us33_n446 ) , .A1( us33_n528 ) , .A3( us33_n577 ) , .A2( us33_n875 ) );
  AOI21_X1 us33_U160 (.A( us33_n670 ) , .B1( us33_n671 ) , .ZN( us33_n672 ) , .B2( us33_n856 ) );
  OAI222_X1 us33_U161 (.B2( us33_n747 ) , .B1( us33_n748 ) , .A2( us33_n749 ) , .ZN( us33_n757 ) , .C2( us33_n805 ) , .C1( us33_n814 ) , .A1( us33_n817 ) );
  OAI222_X1 us33_U162 (.ZN( us33_n505 ) , .C2( us33_n625 ) , .B2( us33_n647 ) , .B1( us33_n747 ) , .A2( us33_n748 ) , .C1( us33_n805 ) , .A1( us33_n806 ) );
  OAI222_X1 us33_U163 (.B2( us33_n708 ) , .ZN( us33_n709 ) , .C2( us33_n724 ) , .B1( us33_n747 ) , .A1( us33_n806 ) , .C1( us33_n814 ) , .A2( us33_n815 ) );
  NAND2_X1 us33_U164 (.A1( us33_n447 ) , .A2( us33_n465 ) , .ZN( us33_n749 ) );
  AOI22_X1 us33_U165 (.ZN( us33_n696 ) , .A1( us33_n830 ) , .B2( us33_n843 ) , .A2( us33_n865 ) , .B1( us33_n868 ) );
  AOI22_X1 us33_U166 (.A2( us33_n782 ) , .ZN( us33_n783 ) , .B2( us33_n831 ) , .A1( us33_n834 ) , .B1( us33_n863 ) );
  INV_X1 us33_U167 (.A( us33_n730 ) , .ZN( us33_n839 ) );
  AOI221_X1 us33_U168 (.A( us33_n764 ) , .ZN( us33_n774 ) , .C2( us33_n810 ) , .B2( us33_n835 ) , .C1( us33_n855 ) , .B1( us33_n866 ) );
  AOI21_X1 us33_U169 (.B2( us33_n763 ) , .ZN( us33_n764 ) , .A( us33_n788 ) , .B1( us33_n792 ) );
  OR4_X1 us33_U17 (.A4( us33_n442 ) , .A2( us33_n443 ) , .A1( us33_n444 ) , .ZN( us33_n445 ) , .A3( us33_n553 ) );
  INV_X1 us33_U170 (.A( us33_n761 ) , .ZN( us33_n835 ) );
  AOI221_X1 us33_U171 (.A( us33_n483 ) , .ZN( us33_n488 ) , .B1( us33_n831 ) , .C2( us33_n844 ) , .C1( us33_n852 ) , .B2( us33_n862 ) );
  OAI22_X1 us33_U172 (.ZN( us33_n483 ) , .A1( us33_n708 ) , .B2( us33_n785 ) , .A2( us33_n806 ) , .B1( us33_n812 ) );
  INV_X1 us33_U173 (.A( us33_n790 ) , .ZN( us33_n832 ) );
  NAND2_X1 us33_U174 (.A1( us33_n451 ) , .A2( us33_n453 ) , .ZN( us33_n762 ) );
  OAI221_X1 us33_U175 (.A( us33_n727 ) , .C2( us33_n728 ) , .B2( us33_n729 ) , .B1( us33_n730 ) , .ZN( us33_n737 ) , .C1( us33_n817 ) );
  AOI22_X1 us33_U176 (.ZN( us33_n727 ) , .B1( us33_n832 ) , .A2( us33_n838 ) , .A1( us33_n863 ) , .B2( us33_n866 ) );
  INV_X1 us33_U177 (.A( us33_n786 ) , .ZN( us33_n862 ) );
  OAI22_X1 us33_U178 (.ZN( us33_n710 ) , .A2( us33_n728 ) , .B2( us33_n729 ) , .A1( us33_n744 ) , .B1( us33_n813 ) );
  INV_X1 us33_U179 (.A( us33_n816 ) , .ZN( us33_n831 ) );
  INV_X1 us33_U18 (.A( us33_n613 ) , .ZN( us33_n875 ) );
  OAI22_X1 us33_U180 (.ZN( us33_n489 ) , .A1( us33_n724 ) , .B2( us33_n728 ) , .B1( us33_n730 ) , .A2( us33_n779 ) );
  OAI22_X1 us33_U181 (.ZN( us33_n624 ) , .B1( us33_n669 ) , .B2( us33_n747 ) , .A1( us33_n815 ) , .A2( us33_n816 ) );
  INV_X1 us33_U182 (.A( us33_n744 ) , .ZN( us33_n837 ) );
  INV_X1 us33_U183 (.A( us33_n788 ) , .ZN( us33_n845 ) );
  OAI22_X1 us33_U184 (.B2( us33_n779 ) , .B1( us33_n780 ) , .ZN( us33_n781 ) , .A2( us33_n814 ) , .A1( us33_n815 ) );
  OAI22_X1 us33_U185 (.A1( us33_n724 ) , .ZN( us33_n726 ) , .B2( us33_n750 ) , .B1( us33_n812 ) , .A2( us33_n816 ) );
  INV_X1 us33_U186 (.A( us33_n805 ) , .ZN( us33_n860 ) );
  INV_X1 us33_U187 (.A( us33_n814 ) , .ZN( us33_n833 ) );
  INV_X1 us33_U188 (.A( us33_n669 ) , .ZN( us33_n865 ) );
  OAI22_X1 us33_U189 (.B2( us33_n744 ) , .ZN( us33_n746 ) , .A2( us33_n762 ) , .B1( us33_n780 ) , .A1( us33_n792 ) );
  INV_X1 us33_U19 (.A( us33_n749 ) , .ZN( us33_n863 ) );
  OAI22_X1 us33_U190 (.ZN( us33_n496 ) , .A2( us33_n744 ) , .A1( us33_n780 ) , .B1( us33_n791 ) , .B2( us33_n806 ) );
  OAI22_X1 us33_U191 (.B2( us33_n803 ) , .B1( us33_n804 ) , .A2( us33_n805 ) , .A1( us33_n806 ) , .ZN( us33_n808 ) );
  AOI211_X1 us33_U192 (.A( us33_n637 ) , .ZN( us33_n645 ) , .B( us33_n743 ) , .C2( us33_n839 ) , .C1( us33_n854 ) );
  OAI22_X1 us33_U193 (.ZN( us33_n637 ) , .A1( us33_n699 ) , .B2( us33_n728 ) , .A2( us33_n762 ) , .B1( us33_n816 ) );
  OAI22_X1 us33_U194 (.B1( us33_n490 ) , .ZN( us33_n491 ) , .A1( us33_n686 ) , .A2( us33_n763 ) , .B2( us33_n817 ) );
  NOR3_X1 us33_U195 (.ZN( us33_n490 ) , .A1( us33_n782 ) , .A2( us33_n850 ) , .A3( us33_n863 ) );
  INV_X1 us33_U196 (.A( us33_n750 ) , .ZN( us33_n842 ) );
  OAI22_X1 us33_U197 (.ZN( us33_n695 ) , .A2( us33_n730 ) , .A1( us33_n780 ) , .B1( us33_n791 ) , .B2( us33_n817 ) );
  NOR2_X1 us33_U198 (.ZN( us33_n715 ) , .A1( us33_n805 ) , .A2( us33_n817 ) );
  NOR2_X1 us33_U199 (.ZN( us33_n666 ) , .A1( us33_n728 ) , .A2( us33_n803 ) );
  AOI222_X1 us33_U20 (.ZN( us33_n605 ) , .B2( us33_n671 ) , .B1( us33_n753 ) , .C2( us33_n831 ) , .A1( us33_n833 ) , .A2( us33_n862 ) , .C1( us33_n863 ) );
  NOR2_X1 us33_U200 (.ZN( us33_n594 ) , .A2( us33_n697 ) , .A1( us33_n728 ) );
  NOR2_X1 us33_U201 (.ZN( us33_n570 ) , .A1( us33_n728 ) , .A2( us33_n806 ) );
  NOR2_X1 us33_U202 (.A2( us33_n744 ) , .ZN( us33_n755 ) , .A1( us33_n805 ) );
  NOR2_X1 us33_U203 (.ZN( us33_n735 ) , .A2( us33_n803 ) , .A1( us33_n805 ) );
  NOR2_X1 us33_U204 (.ZN( us33_n546 ) , .A2( us33_n780 ) , .A1( us33_n814 ) );
  NOR2_X1 us33_U205 (.ZN( us33_n577 ) , .A2( us33_n699 ) , .A1( us33_n814 ) );
  NOR2_X1 us33_U206 (.ZN( us33_n654 ) , .A1( us33_n728 ) , .A2( us33_n813 ) );
  NOR2_X1 us33_U207 (.ZN( us33_n718 ) , .A2( us33_n724 ) , .A1( us33_n744 ) );
  NOR2_X1 us33_U208 (.ZN( us33_n532 ) , .A2( us33_n749 ) , .A1( us33_n750 ) );
  NOR2_X1 us33_U209 (.ZN( us33_n615 ) , .A1( us33_n785 ) , .A2( us33_n815 ) );
  AOI222_X1 us33_U21 (.ZN( us33_n563 ) , .B1( us33_n830 ) , .C1( us33_n841 ) , .A2( us33_n843 ) , .A1( us33_n854 ) , .B2( us33_n863 ) , .C2( us33_n873 ) );
  NOR2_X1 us33_U210 (.ZN( us33_n629 ) , .A2( us33_n728 ) , .A1( us33_n785 ) );
  NOR2_X1 us33_U211 (.ZN( us33_n611 ) , .A2( us33_n780 ) , .A1( us33_n806 ) );
  NOR2_X1 us33_U212 (.ZN( us33_n628 ) , .A2( us33_n669 ) , .A1( us33_n785 ) );
  INV_X1 us33_U213 (.A( us33_n747 ) , .ZN( us33_n834 ) );
  INV_X1 us33_U214 (.A( us33_n728 ) , .ZN( us33_n852 ) );
  NOR2_X1 us33_U215 (.ZN( us33_n652 ) , .A1( us33_n669 ) , .A2( us33_n814 ) );
  NOR2_X1 us33_U216 (.A1( us33_n669 ) , .ZN( us33_n673 ) , .A2( us33_n744 ) );
  NOR2_X1 us33_U217 (.ZN( us33_n602 ) , .A1( us33_n669 ) , .A2( us33_n803 ) );
  NOR2_X1 us33_U218 (.A1( us33_n669 ) , .ZN( us33_n688 ) , .A2( us33_n816 ) );
  NOR2_X1 us33_U219 (.A2( us33_n744 ) , .ZN( us33_n769 ) , .A1( us33_n812 ) );
  AOI222_X1 us33_U22 (.ZN( us33_n660 ) , .A2( us33_n839 ) , .B1( us33_n841 ) , .C2( us33_n845 ) , .A1( us33_n860 ) , .C1( us33_n863 ) , .B2( us33_n870 ) );
  NOR2_X1 us33_U220 (.ZN( us33_n531 ) , .A2( us33_n780 ) , .A1( us33_n816 ) );
  INV_X1 us33_U221 (.A( us33_n792 ) , .ZN( us33_n851 ) );
  NOR2_X1 us33_U222 (.A2( us33_n708 ) , .A1( us33_n750 ) , .ZN( us33_n771 ) );
  NOR2_X1 us33_U223 (.ZN( us33_n599 ) , .A2( us33_n791 ) , .A1( us33_n816 ) );
  NOR2_X1 us33_U224 (.A1( us33_n669 ) , .ZN( us33_n766 ) , .A2( us33_n813 ) );
  NOR2_X1 us33_U225 (.ZN( us33_n601 ) , .A2( us33_n780 ) , .A1( us33_n803 ) );
  NOR2_X1 us33_U226 (.A1( us33_n699 ) , .ZN( us33_n768 ) , .A2( us33_n813 ) );
  NOR2_X1 us33_U227 (.ZN( us33_n541 ) , .A2( us33_n697 ) , .A1( us33_n699 ) );
  NOR2_X1 us33_U228 (.ZN( us33_n527 ) , .A1( us33_n669 ) , .A2( us33_n779 ) );
  NOR2_X1 us33_U229 (.ZN( us33_n667 ) , .A1( us33_n750 ) , .A2( us33_n815 ) );
  INV_X1 us33_U23 (.A( us33_n647 ) , .ZN( us33_n870 ) );
  NOR2_X1 us33_U230 (.ZN( us33_n555 ) , .A1( us33_n750 ) , .A2( us33_n791 ) );
  NOR2_X1 us33_U231 (.ZN( us33_n508 ) , .A2( us33_n780 ) , .A1( us33_n785 ) );
  NOR2_X1 us33_U232 (.ZN( us33_n543 ) , .A2( us33_n708 ) , .A1( us33_n785 ) );
  NOR2_X1 us33_U233 (.ZN( us33_n528 ) , .A2( us33_n724 ) , .A1( us33_n803 ) );
  NOR2_X1 us33_U234 (.ZN( us33_n664 ) , .A1( us33_n785 ) , .A2( us33_n791 ) );
  NOR2_X1 us33_U235 (.ZN( us33_n556 ) , .A1( us33_n762 ) , .A2( us33_n805 ) );
  INV_X1 us33_U236 (.A( us33_n806 ) , .ZN( us33_n841 ) );
  NOR2_X1 us33_U237 (.ZN( us33_n661 ) , .A1( us33_n729 ) , .A2( us33_n790 ) );
  OAI22_X1 us33_U238 (.B1( us33_n440 ) , .ZN( us33_n444 ) , .A2( us33_n728 ) , .A1( us33_n744 ) , .B2( us33_n749 ) );
  NOR3_X1 us33_U239 (.ZN( us33_n440 ) , .A2( us33_n836 ) , .A3( us33_n837 ) , .A1( us33_n846 ) );
  NOR4_X1 us33_U24 (.ZN( us33_n473 ) , .A2( us33_n521 ) , .A4( us33_n594 ) , .A1( us33_n609 ) , .A3( us33_n629 ) );
  NOR2_X1 us33_U240 (.ZN( us33_n507 ) , .A1( us33_n812 ) , .A2( us33_n817 ) );
  NOR2_X1 us33_U241 (.ZN( us33_n557 ) , .A1( us33_n792 ) , .A2( us33_n814 ) );
  NOR2_X1 us33_U242 (.ZN( us33_n545 ) , .A1( us33_n749 ) , .A2( us33_n814 ) );
  NOR2_X1 us33_U243 (.ZN( us33_n509 ) , .A1( us33_n729 ) , .A2( us33_n779 ) );
  NOR2_X1 us33_U244 (.ZN( us33_n662 ) , .A2( us33_n697 ) , .A1( us33_n729 ) );
  OAI22_X1 us33_U245 (.B2( us33_n750 ) , .B1( us33_n751 ) , .A1( us33_n752 ) , .ZN( us33_n756 ) , .A2( us33_n806 ) );
  NOR2_X1 us33_U246 (.ZN( us33_n751 ) , .A2( us33_n852 ) , .A1( us33_n860 ) );
  NOR3_X1 us33_U247 (.ZN( us33_n752 ) , .A2( us33_n853 ) , .A1( us33_n863 ) , .A3( us33_n865 ) );
  NOR2_X1 us33_U248 (.ZN( us33_n544 ) , .A2( us33_n785 ) , .A1( us33_n792 ) );
  NOR2_X1 us33_U249 (.ZN( us33_n663 ) , .A1( us33_n729 ) , .A2( us33_n785 ) );
  NOR4_X1 us33_U25 (.ZN( us33_n479 ) , .A1( us33_n520 ) , .A4( us33_n557 ) , .A3( us33_n582 ) , .A2( us33_n630 ) );
  NOR2_X1 us33_U250 (.ZN( us33_n530 ) , .A2( us33_n744 ) , .A1( us33_n792 ) );
  NOR2_X1 us33_U251 (.ZN( us33_n506 ) , .A2( us33_n728 ) , .A1( us33_n762 ) );
  NOR2_X1 us33_U252 (.ZN( us33_n631 ) , .A1( us33_n724 ) , .A2( us33_n813 ) );
  NOR2_X1 us33_U253 (.ZN( us33_n614 ) , .A1( us33_n762 ) , .A2( us33_n812 ) );
  NOR2_X1 us33_U254 (.A1( us33_n749 ) , .ZN( us33_n767 ) , .A2( us33_n803 ) );
  NOR2_X1 us33_U255 (.ZN( us33_n516 ) , .A1( us33_n708 ) , .A2( us33_n744 ) );
  NOR2_X1 us33_U256 (.ZN( us33_n670 ) , .A1( us33_n790 ) , .A2( us33_n805 ) );
  NOR2_X1 us33_U257 (.ZN( us33_n558 ) , .A1( us33_n708 ) , .A2( us33_n816 ) );
  NOR2_X1 us33_U258 (.A2( us33_n697 ) , .ZN( us33_n716 ) , .A1( us33_n792 ) );
  NOR2_X1 us33_U259 (.ZN( us33_n517 ) , .A1( us33_n708 ) , .A2( us33_n803 ) );
  NOR4_X1 us33_U26 (.A4( us33_n532 ) , .A3( us33_n533 ) , .A2( us33_n534 ) , .ZN( us33_n535 ) , .A1( us33_n820 ) );
  NOR2_X1 us33_U260 (.ZN( us33_n521 ) , .A1( us33_n790 ) , .A2( us33_n812 ) );
  NOR2_X1 us33_U261 (.ZN( us33_n630 ) , .A1( us33_n747 ) , .A2( us33_n815 ) );
  NOR2_X1 us33_U262 (.ZN( us33_n655 ) , .A1( us33_n790 ) , .A2( us33_n815 ) );
  INV_X1 us33_U263 (.A( us33_n763 ) , .ZN( us33_n866 ) );
  AOI21_X1 us33_U264 (.ZN( us33_n552 ) , .B1( us33_n669 ) , .A( us33_n697 ) , .B2( us33_n805 ) );
  NOR2_X1 us33_U265 (.ZN( us33_n668 ) , .A2( us33_n708 ) , .A1( us33_n790 ) );
  NOR2_X1 us33_U266 (.ZN( us33_n542 ) , .A1( us33_n762 ) , .A2( us33_n791 ) );
  NOR2_X1 us33_U267 (.ZN( us33_n656 ) , .A1( us33_n747 ) , .A2( us33_n780 ) );
  NOR2_X1 us33_U268 (.ZN( us33_n609 ) , .A2( us33_n724 ) , .A1( us33_n817 ) );
  INV_X1 us33_U269 (.A( us33_n729 ) , .ZN( us33_n868 ) );
  NOR4_X1 us33_U27 (.ZN( us33_n456 ) , .A2( us33_n517 ) , .A1( us33_n543 ) , .A3( us33_n579 ) , .A4( us33_n615 ) );
  AOI21_X1 us33_U270 (.B1( us33_n625 ) , .ZN( us33_n627 ) , .A( us33_n763 ) , .B2( us33_n814 ) );
  AOI21_X1 us33_U271 (.ZN( us33_n650 ) , .A( us33_n779 ) , .B1( us33_n792 ) , .B2( us33_n805 ) );
  AOI21_X1 us33_U272 (.A( us33_n815 ) , .B2( us33_n816 ) , .B1( us33_n817 ) , .ZN( us33_n818 ) );
  NOR2_X1 us33_U273 (.ZN( us33_n579 ) , .A2( us33_n708 ) , .A1( us33_n730 ) );
  NOR2_X1 us33_U274 (.ZN( us33_n533 ) , .A2( us33_n724 ) , .A1( us33_n730 ) );
  NOR2_X1 us33_U275 (.ZN( us33_n642 ) , .A2( us33_n788 ) , .A1( us33_n791 ) );
  AOI21_X1 us33_U276 (.A( us33_n812 ) , .B2( us33_n813 ) , .B1( us33_n814 ) , .ZN( us33_n819 ) );
  NOR2_X1 us33_U277 (.A2( us33_n708 ) , .A1( us33_n762 ) , .ZN( us33_n794 ) );
  NOR2_X1 us33_U278 (.A2( us33_n697 ) , .A1( us33_n780 ) , .ZN( us33_n820 ) );
  AOI21_X1 us33_U279 (.ZN( us33_n626 ) , .B2( us33_n669 ) , .A( us33_n790 ) , .B1( us33_n791 ) );
  NOR4_X1 us33_U28 (.A4( us33_n541 ) , .A3( us33_n542 ) , .A2( us33_n543 ) , .ZN( us33_n550 ) , .A1( us33_n688 ) );
  AOI21_X1 us33_U280 (.ZN( us33_n499 ) , .B1( us33_n680 ) , .A( us33_n812 ) , .B2( us33_n816 ) );
  NOR2_X1 us33_U281 (.ZN( us33_n520 ) , .A2( us33_n708 ) , .A1( us33_n814 ) );
  AOI21_X1 us33_U282 (.ZN( us33_n477 ) , .A( us33_n669 ) , .B1( us33_n750 ) , .B2( us33_n806 ) );
  NOR2_X1 us33_U283 (.ZN( us33_n582 ) , .A1( us33_n744 ) , .A2( us33_n815 ) );
  AOI21_X1 us33_U284 (.ZN( us33_n593 ) , .B1( us33_n750 ) , .A( us33_n792 ) , .B2( us33_n813 ) );
  AOI21_X1 us33_U285 (.ZN( us33_n515 ) , .A( us33_n729 ) , .B1( us33_n750 ) , .B2( us33_n803 ) );
  NOR2_X1 us33_U286 (.A1( us33_n697 ) , .ZN( us33_n770 ) , .A2( us33_n815 ) );
  AOI21_X1 us33_U287 (.ZN( us33_n510 ) , .B2( us33_n669 ) , .A( us33_n730 ) , .B1( us33_n815 ) );
  NOR2_X1 us33_U288 (.ZN( us33_n519 ) , .A2( us33_n699 ) , .A1( us33_n816 ) );
  NOR2_X1 us33_U289 (.ZN( us33_n559 ) , .A2( us33_n791 ) , .A1( us33_n803 ) );
  AOI221_X1 us33_U29 (.A( us33_n713 ) , .B2( us33_n714 ) , .ZN( us33_n720 ) , .C1( us33_n832 ) , .B1( us33_n839 ) , .C2( us33_n863 ) );
  NOR2_X1 us33_U290 (.ZN( us33_n581 ) , .A1( us33_n669 ) , .A2( us33_n788 ) );
  INV_X1 us33_U291 (.A( us33_n813 ) , .ZN( us33_n836 ) );
  NOR2_X1 us33_U292 (.ZN( us33_n683 ) , .A2( us33_n699 ) , .A1( us33_n803 ) );
  AOI21_X1 us33_U293 (.ZN( us33_n589 ) , .B2( us33_n699 ) , .B1( us33_n815 ) , .A( us33_n817 ) );
  AOI21_X1 us33_U294 (.ZN( us33_n539 ) , .B2( us33_n812 ) , .A( us33_n814 ) , .B1( us33_n815 ) );
  AOI21_X1 us33_U295 (.ZN( us33_n540 ) , .A( us33_n763 ) , .B2( us33_n779 ) , .B1( us33_n817 ) );
  AOI21_X1 us33_U296 (.B1( us33_n699 ) , .ZN( us33_n700 ) , .A( us33_n732 ) , .B2( us33_n763 ) );
  AOI21_X1 us33_U297 (.ZN( us33_n591 ) , .B2( us33_n763 ) , .A( us33_n785 ) , .B1( us33_n812 ) );
  AOI21_X1 us33_U298 (.ZN( us33_n498 ) , .A( us33_n724 ) , .B2( us33_n762 ) , .B1( us33_n814 ) );
  NOR2_X1 us33_U299 (.ZN( us33_n547 ) , .A1( us33_n699 ) , .A2( us33_n744 ) );
  NAND2_X1 us33_U3 (.A1( us33_n441 ) , .A2( us33_n464 ) , .ZN( us33_n708 ) );
  OR2_X1 us33_U30 (.A2( us33_n711 ) , .A1( us33_n712 ) , .ZN( us33_n713 ) );
  INV_X1 us33_U300 (.A( us33_n791 ) , .ZN( us33_n873 ) );
  AOI21_X1 us33_U301 (.ZN( us33_n649 ) , .B1( us33_n729 ) , .B2( us33_n763 ) , .A( us33_n813 ) );
  NOR2_X1 us33_U302 (.ZN( us33_n685 ) , .A1( us33_n729 ) , .A2( us33_n816 ) );
  AOI21_X1 us33_U303 (.B1( us33_n686 ) , .ZN( us33_n687 ) , .A( us33_n728 ) , .B2( us33_n761 ) );
  AOI21_X1 us33_U304 (.ZN( us33_n569 ) , .B1( us33_n750 ) , .B2( us33_n762 ) , .A( us33_n780 ) );
  AOI21_X1 us33_U305 (.ZN( us33_n571 ) , .B2( us33_n697 ) , .B1( us33_n806 ) , .A( us33_n812 ) );
  NOR2_X1 us33_U306 (.ZN( us33_n568 ) , .A1( us33_n729 ) , .A2( us33_n762 ) );
  NOR2_X1 us33_U307 (.ZN( us33_n566 ) , .A2( us33_n697 ) , .A1( us33_n763 ) );
  AOI21_X1 us33_U308 (.ZN( us33_n640 ) , .B2( us33_n747 ) , .A( us33_n792 ) , .B1( us33_n803 ) );
  INV_X1 us33_U309 (.A( us33_n699 ) , .ZN( us33_n853 ) );
  NOR2_X1 us33_U31 (.ZN( us33_n680 ) , .A2( us33_n834 ) , .A1( us33_n839 ) );
  AOI21_X1 us33_U310 (.ZN( us33_n514 ) , .A( us33_n779 ) , .B2( us33_n792 ) , .B1( us33_n812 ) );
  AOI21_X1 us33_U311 (.ZN( us33_n639 ) , .B2( us33_n749 ) , .A( us33_n788 ) , .B1( us33_n812 ) );
  NAND2_X1 us33_U312 (.ZN( us33_n753 ) , .A1( us33_n763 ) , .A2( us33_n805 ) );
  NOR2_X1 us33_U313 (.ZN( us33_n665 ) , .A1( us33_n780 ) , .A2( us33_n813 ) );
  AOI21_X1 us33_U314 (.ZN( us33_n564 ) , .B1( us33_n724 ) , .A( us33_n779 ) , .B2( us33_n791 ) );
  AOI21_X1 us33_U315 (.ZN( us33_n497 ) , .A( us33_n779 ) , .B2( us33_n791 ) , .B1( us33_n804 ) );
  AOI21_X1 us33_U316 (.ZN( us33_n689 ) , .B2( us33_n749 ) , .B1( us33_n763 ) , .A( us33_n806 ) );
  AOI21_X1 us33_U317 (.ZN( us33_n450 ) , .B2( us33_n792 ) , .A( us33_n803 ) , .B1( us33_n815 ) );
  NOR2_X1 us33_U318 (.ZN( us33_n567 ) , .A1( us33_n747 ) , .A2( us33_n805 ) );
  NOR2_X1 us33_U319 (.ZN( us33_n529 ) , .A1( us33_n708 ) , .A2( us33_n779 ) );
  AOI222_X1 us33_U32 (.ZN( us33_n469 ) , .B1( us33_n832 ) , .A1( us33_n839 ) , .C1( us33_n842 ) , .C2( us33_n851 ) , .A2( us33_n855 ) , .B2( us33_n865 ) );
  NOR2_X1 us33_U320 (.ZN( us33_n578 ) , .A1( us33_n708 ) , .A2( us33_n813 ) );
  AOI21_X1 us33_U321 (.ZN( us33_n478 ) , .B2( us33_n697 ) , .A( us33_n749 ) , .B1( us33_n779 ) );
  AOI21_X1 us33_U322 (.A( us33_n790 ) , .B2( us33_n791 ) , .B1( us33_n792 ) , .ZN( us33_n793 ) );
  NOR2_X1 us33_U323 (.ZN( us33_n684 ) , .A1( us33_n791 ) , .A2( us33_n813 ) );
  AOI21_X1 us33_U324 (.A( us33_n733 ) , .ZN( us33_n734 ) , .B2( us33_n780 ) , .B1( us33_n792 ) );
  NOR2_X1 us33_U325 (.A2( us33_n813 ) , .A1( us33_n815 ) , .ZN( us33_n821 ) );
  AOI21_X1 us33_U326 (.ZN( us33_n641 ) , .B1( us33_n680 ) , .A( us33_n791 ) , .B2( us33_n817 ) );
  NOR2_X1 us33_U327 (.ZN( us33_n711 ) , .A1( us33_n762 ) , .A2( us33_n763 ) );
  NOR2_X1 us33_U328 (.ZN( us33_n583 ) , .A1( us33_n792 ) , .A2( us33_n817 ) );
  NOR2_X1 us33_U329 (.ZN( us33_n534 ) , .A1( us33_n724 ) , .A2( us33_n788 ) );
  NOR4_X1 us33_U33 (.A1( us33_n466 ) , .ZN( us33_n467 ) , .A4( us33_n542 ) , .A2( us33_n554 ) , .A3( us33_n614 ) );
  NOR2_X1 us33_U330 (.ZN( us33_n632 ) , .A2( us33_n697 ) , .A1( us33_n724 ) );
  NOR2_X1 us33_U331 (.ZN( us33_n682 ) , .A2( us33_n708 ) , .A1( us33_n817 ) );
  NOR2_X1 us33_U332 (.ZN( us33_n580 ) , .A2( us33_n697 ) , .A1( us33_n791 ) );
  INV_X1 us33_U333 (.A( us33_n815 ) , .ZN( us33_n855 ) );
  AOI21_X1 us33_U334 (.ZN( us33_n442 ) , .A( us33_n699 ) , .B1( us33_n733 ) , .B2( us33_n750 ) );
  INV_X1 us33_U335 (.A( us33_n780 ) , .ZN( us33_n850 ) );
  INV_X1 us33_U336 (.A( us33_n785 ) , .ZN( us33_n846 ) );
  NAND2_X1 us33_U337 (.ZN( us33_n714 ) , .A1( us33_n728 ) , .A2( us33_n780 ) );
  NAND2_X1 us33_U338 (.A2( us33_n762 ) , .A1( us33_n806 ) , .ZN( us33_n810 ) );
  AOI21_X1 us33_U339 (.ZN( us33_n443 ) , .B1( us33_n789 ) , .B2( us33_n791 ) , .A( us33_n814 ) );
  AOI221_X1 us33_U34 (.ZN( us33_n468 ) , .C2( us33_n714 ) , .B2( us33_n831 ) , .C1( us33_n845 ) , .B1( us33_n860 ) , .A( us33_n864 ) );
  NAND2_X1 us33_U340 (.ZN( us33_n671 ) , .A1( us33_n806 ) , .A2( us33_n816 ) );
  NOR2_X1 us33_U341 (.ZN( us33_n484 ) , .A1( us33_n788 ) , .A2( us33_n805 ) );
  NOR2_X1 us33_U342 (.ZN( us33_n470 ) , .A2( us33_n779 ) , .A1( us33_n815 ) );
  NOR2_X1 us33_U343 (.ZN( us33_n712 ) , .A2( us33_n724 ) , .A1( us33_n790 ) );
  OAI21_X1 us33_U344 (.A( us33_n787 ) , .B2( us33_n788 ) , .B1( us33_n789 ) , .ZN( us33_n795 ) );
  OAI21_X1 us33_U345 (.ZN( us33_n787 ) , .A( us33_n839 ) , .B1( us33_n863 ) , .B2( us33_n873 ) );
  NOR2_X1 us33_U346 (.ZN( us33_n526 ) , .A1( us33_n724 ) , .A2( us33_n750 ) );
  NAND2_X1 us33_U347 (.A1( us33_n699 ) , .A2( us33_n729 ) , .ZN( us33_n782 ) );
  NOR2_X1 us33_U348 (.ZN( us33_n518 ) , .A1( us33_n708 ) , .A2( us33_n788 ) );
  OAI21_X1 us33_U349 (.A( us33_n698 ) , .ZN( us33_n702 ) , .B2( us33_n750 ) , .B1( us33_n804 ) );
  NOR4_X1 us33_U35 (.A4( us33_n514 ) , .A3( us33_n515 ) , .A2( us33_n516 ) , .A1( us33_n517 ) , .ZN( us33_n524 ) );
  OAI21_X1 us33_U350 (.ZN( us33_n698 ) , .B2( us33_n833 ) , .B1( us33_n838 ) , .A( us33_n860 ) );
  OAI21_X1 us33_U351 (.A( us33_n731 ) , .B1( us33_n732 ) , .ZN( us33_n736 ) , .B2( us33_n805 ) );
  OAI21_X1 us33_U352 (.ZN( us33_n731 ) , .A( us33_n833 ) , .B2( us33_n852 ) , .B1( us33_n873 ) );
  INV_X1 us33_U353 (.A( us33_n817 ) , .ZN( us33_n844 ) );
  INV_X1 us33_U354 (.A( us33_n724 ) , .ZN( us33_n856 ) );
  AND2_X1 us33_U355 (.ZN( us33_n732 ) , .A1( us33_n779 ) , .A2( us33_n785 ) );
  NAND2_X1 us33_U356 (.A1( us33_n447 ) , .A2( us33_n449 ) , .ZN( us33_n805 ) );
  NAND2_X1 us33_U357 (.A1( us33_n451 ) , .A2( us33_n454 ) , .ZN( us33_n814 ) );
  NAND2_X1 us33_U358 (.A1( us33_n452 ) , .A2( us33_n465 ) , .ZN( us33_n669 ) );
  NAND2_X1 us33_U359 (.A2( us33_n448 ) , .A1( us33_n460 ) , .ZN( us33_n728 ) );
  AOI222_X1 us33_U36 (.ZN( us33_n525 ) , .A1( us33_n834 ) , .B2( us33_n837 ) , .C1( us33_n844 ) , .C2( us33_n850 ) , .A2( us33_n852 ) , .B1( us33_n866 ) );
  NAND2_X1 us33_U360 (.A1( us33_n455 ) , .A2( us33_n462 ) , .ZN( us33_n750 ) );
  NAND2_X1 us33_U361 (.A2( us33_n453 ) , .A1( us33_n455 ) , .ZN( us33_n806 ) );
  NAND2_X1 us33_U362 (.A1( us33_n451 ) , .A2( us33_n471 ) , .ZN( us33_n816 ) );
  NAND2_X1 us33_U363 (.A1( us33_n454 ) , .A2( us33_n461 ) , .ZN( us33_n813 ) );
  NAND2_X1 us33_U364 (.A1( us33_n455 ) , .A2( us33_n471 ) , .ZN( us33_n803 ) );
  NAND2_X1 us33_U365 (.A1( us33_n453 ) , .A2( us33_n461 ) , .ZN( us33_n744 ) );
  NAND2_X1 us33_U366 (.A1( us33_n453 ) , .A2( us33_n472 ) , .ZN( us33_n785 ) );
  NAND2_X1 us33_U367 (.A2( us33_n454 ) , .A1( us33_n472 ) , .ZN( us33_n779 ) );
  NAND2_X1 us33_U368 (.A2( us33_n464 ) , .A1( us33_n465 ) , .ZN( us33_n812 ) );
  NAND2_X1 us33_U369 (.A1( us33_n441 ) , .A2( us33_n460 ) , .ZN( us33_n699 ) );
  NOR4_X1 us33_U37 (.A3( us33_n521 ) , .A1( us33_n522 ) , .ZN( us33_n523 ) , .A2( us33_n673 ) , .A4( us33_n769 ) );
  NAND2_X1 us33_U370 (.A2( us33_n449 ) , .A1( us33_n452 ) , .ZN( us33_n763 ) );
  NAND2_X1 us33_U371 (.A2( us33_n448 ) , .A1( us33_n452 ) , .ZN( us33_n729 ) );
  NAND2_X1 us33_U372 (.A2( us33_n461 ) , .A1( us33_n462 ) , .ZN( us33_n747 ) );
  NAND2_X1 us33_U373 (.A1( us33_n462 ) , .A2( us33_n472 ) , .ZN( us33_n788 ) );
  NOR2_X1 us33_U374 (.ZN( us33_n465 ) , .A2( us33_n847 ) , .A1( us33_n848 ) );
  NOR2_X1 us33_U375 (.ZN( us33_n453 ) , .A1( us33_n826 ) , .A2( us33_n827 ) );
  NOR2_X1 us33_U376 (.ZN( us33_n451 ) , .A1( us33_n828 ) , .A2( us33_n829 ) );
  NAND2_X1 us33_U377 (.A1( us33_n451 ) , .A2( us33_n462 ) , .ZN( us33_n790 ) );
  NAND2_X2 us33_U378 (.A2( us33_n448 ) , .A1( us33_n464 ) , .ZN( us33_n815 ) );
  NAND2_X1 us33_U379 (.A2( us33_n441 ) , .A1( us33_n447 ) , .ZN( us33_n784 ) );
  AOI221_X1 us33_U38 (.A( us33_n781 ) , .ZN( us33_n798 ) , .C2( us33_n837 ) , .B2( us33_n838 ) , .B1( us33_n865 ) , .C1( us33_n866 ) );
  NAND2_X1 us33_U380 (.A2( us33_n454 ) , .A1( us33_n455 ) , .ZN( us33_n730 ) );
  NAND2_X2 us33_U381 (.A1( us33_n449 ) , .A2( us33_n464 ) , .ZN( us33_n724 ) );
  NAND2_X2 us33_U382 (.A1( us33_n449 ) , .A2( us33_n460 ) , .ZN( us33_n792 ) );
  NAND2_X2 us33_U383 (.A2( us33_n460 ) , .A1( us33_n465 ) , .ZN( us33_n780 ) );
  NOR2_X1 us33_U384 (.ZN( us33_n447 ) , .A2( us33_n849 ) , .A1( us33_n858 ) );
  NAND2_X1 us33_U385 (.A1( us33_n447 ) , .A2( us33_n448 ) , .ZN( us33_n786 ) );
  NOR2_X1 us33_U386 (.A2( sa33_6 ) , .A1( sa33_7 ) , .ZN( us33_n464 ) );
  NOR2_X1 us33_U387 (.A2( sa33_7 ) , .ZN( us33_n460 ) , .A1( us33_n849 ) );
  NOR2_X1 us33_U388 (.A2( sa33_4 ) , .ZN( us33_n449 ) , .A1( us33_n848 ) );
  NOR2_X1 us33_U389 (.A2( sa33_4 ) , .A1( sa33_5 ) , .ZN( us33_n441 ) );
  NOR4_X1 us33_U39 (.A4( us33_n793 ) , .A3( us33_n794 ) , .A2( us33_n795 ) , .A1( us33_n796 ) , .ZN( us33_n797 ) );
  NOR2_X1 us33_U390 (.A2( sa33_5 ) , .ZN( us33_n448 ) , .A1( us33_n847 ) );
  NOR2_X1 us33_U391 (.A2( sa33_2 ) , .A1( sa33_3 ) , .ZN( us33_n472 ) );
  NOR2_X1 us33_U392 (.A2( sa33_6 ) , .ZN( us33_n452 ) , .A1( us33_n858 ) );
  NOR2_X1 us33_U393 (.A2( sa33_1 ) , .ZN( us33_n471 ) , .A1( us33_n826 ) );
  NOR2_X1 us33_U394 (.A2( sa33_0 ) , .ZN( us33_n454 ) , .A1( us33_n827 ) );
  NOR2_X1 us33_U395 (.A2( sa33_0 ) , .A1( sa33_1 ) , .ZN( us33_n462 ) );
  NOR2_X1 us33_U396 (.A2( sa33_3 ) , .ZN( us33_n455 ) , .A1( us33_n828 ) );
  NOR2_X1 us33_U397 (.A2( sa33_2 ) , .ZN( us33_n461 ) , .A1( us33_n829 ) );
  INV_X1 us33_U398 (.A( sa33_6 ) , .ZN( us33_n849 ) );
  INV_X1 us33_U399 (.A( sa33_4 ) , .ZN( us33_n847 ) );
  NAND2_X1 us33_U4 (.A2( us33_n441 ) , .A1( us33_n452 ) , .ZN( us33_n791 ) );
  NOR4_X1 us33_U40 (.A4( us33_n776 ) , .A3( us33_n777 ) , .A1( us33_n778 ) , .ZN( us33_n799 ) , .A2( us33_n801 ) );
  INV_X1 us33_U400 (.A( sa33_3 ) , .ZN( us33_n829 ) );
  INV_X1 us33_U401 (.A( sa33_1 ) , .ZN( us33_n827 ) );
  INV_X1 us33_U402 (.A( sa33_0 ) , .ZN( us33_n826 ) );
  INV_X1 us33_U403 (.A( sa33_2 ) , .ZN( us33_n828 ) );
  INV_X1 us33_U404 (.A( sa33_7 ) , .ZN( us33_n858 ) );
  INV_X1 us33_U405 (.A( sa33_5 ) , .ZN( us33_n848 ) );
  NAND2_X1 us33_U406 (.A2( us33_n461 ) , .A1( us33_n471 ) , .ZN( us33_n697 ) );
  OAI221_X1 us33_U407 (.A( us33_n783 ) , .C2( us33_n784 ) , .B2( us33_n785 ) , .B1( us33_n786 ) , .ZN( us33_n796 ) , .C1( us33_n813 ) );
  NAND2_X1 us33_U408 (.A1( us33_n729 ) , .A2( us33_n784 ) , .ZN( us33_n811 ) );
  OAI22_X1 us33_U409 (.ZN( us33_n588 ) , .A2( us33_n747 ) , .B2( us33_n762 ) , .A1( us33_n763 ) , .B1( us33_n784 ) );
  NOR4_X1 us33_U41 (.A3( us33_n755 ) , .A2( us33_n756 ) , .A1( us33_n757 ) , .ZN( us33_n758 ) , .A4( us33_n869 ) );
  AOI21_X1 us33_U410 (.ZN( us33_n592 ) , .B1( us33_n728 ) , .B2( us33_n784 ) , .A( us33_n790 ) );
  AOI21_X1 us33_U411 (.ZN( us33_n623 ) , .B1( us33_n699 ) , .A( us33_n779 ) , .B2( us33_n784 ) );
  AOI21_X1 us33_U412 (.ZN( us33_n648 ) , .A( us33_n762 ) , .B2( us33_n784 ) , .B1( us33_n792 ) );
  OAI22_X1 us33_U413 (.ZN( us33_n681 ) , .A1( us33_n699 ) , .A2( us33_n730 ) , .B2( us33_n784 ) , .B1( us33_n817 ) );
  OAI21_X1 us33_U414 (.A( us33_n613 ) , .ZN( us33_n616 ) , .B1( us33_n625 ) , .B2( us33_n784 ) );
  NOR2_X1 us33_U415 (.ZN( us33_n610 ) , .A1( us33_n784 ) , .A2( us33_n816 ) );
  OAI222_X1 us33_U416 (.A2( us33_n669 ) , .ZN( us33_n674 ) , .B1( us33_n747 ) , .B2( us33_n784 ) , .C2( us33_n788 ) , .C1( us33_n815 ) , .A1( us33_n817 ) );
  NOR2_X1 us33_U417 (.ZN( us33_n651 ) , .A1( us33_n784 ) , .A2( us33_n788 ) );
  NOR2_X1 us33_U418 (.ZN( us33_n600 ) , .A2( us33_n697 ) , .A1( us33_n784 ) );
  NOR2_X1 us33_U419 (.ZN( us33_n553 ) , .A2( us33_n744 ) , .A1( us33_n784 ) );
  AOI211_X1 us33_U42 (.B( us33_n745 ) , .A( us33_n746 ) , .ZN( us33_n759 ) , .C1( us33_n832 ) , .C2( us33_n853 ) );
  INV_X1 us33_U420 (.A( us33_n784 ) , .ZN( us33_n861 ) );
  AOI21_X1 us33_U421 (.ZN( us33_n500 ) , .A( us33_n697 ) , .B1( us33_n708 ) , .B2( us33_n786 ) );
  OAI221_X1 us33_U422 (.A( us33_n696 ) , .ZN( us33_n703 ) , .C2( us33_n784 ) , .C1( us33_n785 ) , .B1( us33_n786 ) , .B2( us33_n806 ) );
  OAI22_X1 us33_U423 (.ZN( us33_n590 ) , .B1( us33_n730 ) , .B2( us33_n749 ) , .A2( us33_n786 ) , .A1( us33_n803 ) );
  NOR2_X1 us33_U424 (.ZN( us33_n612 ) , .A1( us33_n779 ) , .A2( us33_n786 ) );
  NAND2_X1 us33_U425 (.A2( us33_n749 ) , .A1( us33_n786 ) , .ZN( us33_n809 ) );
  OAI222_X1 us33_U426 (.ZN( us33_n617 ) , .B1( us33_n697 ) , .C1( us33_n724 ) , .C2( us33_n747 ) , .B2( us33_n786 ) , .A2( us33_n792 ) , .A1( us33_n816 ) );
  NOR2_X1 us33_U427 (.ZN( us33_n717 ) , .A2( us33_n744 ) , .A1( us33_n786 ) );
  NOR2_X1 us33_U428 (.ZN( us33_n653 ) , .A1( us33_n762 ) , .A2( us33_n786 ) );
  NOR2_X1 us33_U429 (.ZN( us33_n554 ) , .A1( us33_n786 ) , .A2( us33_n813 ) );
  NOR3_X1 us33_U43 (.A3( us33_n741 ) , .A2( us33_n742 ) , .A1( us33_n743 ) , .ZN( us33_n760 ) );
  NOR2_X1 us33_U430 (.ZN( us33_n701 ) , .A2( us33_n786 ) , .A1( us33_n817 ) );
  NOR2_X1 us33_U431 (.A1( us33_n730 ) , .ZN( us33_n765 ) , .A2( us33_n786 ) );
  AND2_X1 us33_U432 (.ZN( us33_n438 ) , .A2( us33_n831 ) , .A1( us33_n854 ) );
  AND2_X1 us33_U433 (.ZN( us33_n439 ) , .A2( us33_n843 ) , .A1( us33_n861 ) );
  NOR3_X1 us33_U434 (.A1( us33_n438 ) , .A2( us33_n439 ) , .A3( us33_n576 ) , .ZN( us33_n587 ) );
  NAND4_X1 us33_U435 (.ZN( sa30_sr_2 ) , .A4( us33_n643 ) , .A3( us33_n644 ) , .A2( us33_n645 ) , .A1( us33_n646 ) );
  INV_X1 us33_U436 (.A( us33_n812 ) , .ZN( us33_n854 ) );
  NAND3_X1 us33_U437 (.ZN( sa30_sr_6 ) , .A3( us33_n797 ) , .A2( us33_n798 ) , .A1( us33_n799 ) );
  NAND3_X1 us33_U438 (.ZN( sa30_sr_5 ) , .A3( us33_n758 ) , .A2( us33_n759 ) , .A1( us33_n760 ) );
  NAND3_X1 us33_U439 (.ZN( sa30_sr_4 ) , .A3( us33_n738 ) , .A2( us33_n739 ) , .A1( us33_n740 ) );
  NAND4_X1 us33_U44 (.ZN( sa30_sr_3 ) , .A4( us33_n704 ) , .A3( us33_n705 ) , .A2( us33_n706 ) , .A1( us33_n707 ) );
  NAND3_X1 us33_U440 (.A3( us33_n675 ) , .A2( us33_n676 ) , .A1( us33_n677 ) , .ZN( us33_n807 ) );
  NAND3_X1 us33_U441 (.ZN( us33_n638 ) , .A3( us33_n708 ) , .A2( us33_n724 ) , .A1( us33_n792 ) );
  NAND3_X1 us33_U442 (.A3( us33_n618 ) , .A2( us33_n619 ) , .A1( us33_n620 ) , .ZN( us33_n725 ) );
  NAND3_X1 us33_U443 (.A3( us33_n585 ) , .A2( us33_n586 ) , .A1( us33_n587 ) , .ZN( us33_n621 ) );
  NAND3_X1 us33_U444 (.ZN( us33_n565 ) , .A3( us33_n680 ) , .A2( us33_n750 ) , .A1( us33_n785 ) );
  NAND3_X1 us33_U445 (.A3( us33_n523 ) , .A2( us33_n524 ) , .A1( us33_n525 ) , .ZN( us33_n742 ) );
  NAND3_X1 us33_U446 (.A3( us33_n512 ) , .A1( us33_n513 ) , .ZN( us33_n608 ) , .A2( us33_n871 ) );
  NAND3_X1 us33_U447 (.A3( us33_n467 ) , .A2( us33_n468 ) , .A1( us33_n469 ) , .ZN( us33_n777 ) );
  INV_X1 us33_U448 (.A( us33_n803 ) , .ZN( us33_n843 ) );
  AOI21_X1 us33_U449 (.ZN( us33_n576 ) , .B2( us33_n724 ) , .B1( us33_n748 ) , .A( us33_n785 ) );
  NOR4_X1 us33_U45 (.A4( us33_n700 ) , .A3( us33_n701 ) , .A2( us33_n702 ) , .A1( us33_n703 ) , .ZN( us33_n704 ) );
  AOI211_X1 us33_U46 (.B( us33_n694 ) , .A( us33_n695 ) , .ZN( us33_n705 ) , .C2( us33_n831 ) , .C1( us33_n851 ) );
  NOR2_X1 us33_U47 (.ZN( us33_n707 ) , .A2( us33_n776 ) , .A1( us33_n800 ) );
  AOI222_X1 us33_U48 (.B2( us33_n638 ) , .ZN( us33_n644 ) , .B1( us33_n841 ) , .A1( us33_n842 ) , .C2( us33_n846 ) , .C1( us33_n863 ) , .A2( us33_n865 ) );
  NOR4_X1 us33_U49 (.A4( us33_n639 ) , .A3( us33_n640 ) , .A2( us33_n641 ) , .A1( us33_n642 ) , .ZN( us33_n643 ) );
  NAND2_X1 us33_U5 (.A2( us33_n471 ) , .A1( us33_n472 ) , .ZN( us33_n817 ) );
  NOR3_X1 us33_U50 (.A2( us33_n607 ) , .A1( us33_n608 ) , .ZN( us33_n646 ) , .A3( us33_n722 ) );
  NOR2_X1 us33_U51 (.ZN( us33_n804 ) , .A1( us33_n854 ) , .A2( us33_n861 ) );
  NAND4_X1 us33_U52 (.ZN( sa30_sr_7 ) , .A4( us33_n822 ) , .A3( us33_n823 ) , .A2( us33_n824 ) , .A1( us33_n825 ) );
  NOR4_X1 us33_U53 (.A4( us33_n818 ) , .A3( us33_n819 ) , .A2( us33_n820 ) , .A1( us33_n821 ) , .ZN( us33_n822 ) );
  AOI222_X1 us33_U54 (.C2( us33_n809 ) , .B2( us33_n810 ) , .A2( us33_n811 ) , .ZN( us33_n823 ) , .C1( us33_n832 ) , .A1( us33_n839 ) , .B1( us33_n853 ) );
  AOI211_X1 us33_U55 (.B( us33_n807 ) , .A( us33_n808 ) , .ZN( us33_n824 ) , .C1( us33_n842 ) , .C2( us33_n850 ) );
  NAND4_X1 us33_U56 (.ZN( sa30_sr_0 ) , .A4( us33_n501 ) , .A3( us33_n502 ) , .A2( us33_n503 ) , .A1( us33_n504 ) );
  AOI221_X1 us33_U57 (.A( us33_n497 ) , .ZN( us33_n502 ) , .B2( us33_n843 ) , .C1( us33_n846 ) , .C2( us33_n860 ) , .B1( us33_n862 ) );
  NOR4_X1 us33_U58 (.A4( us33_n498 ) , .A3( us33_n499 ) , .A2( us33_n500 ) , .ZN( us33_n501 ) , .A1( us33_n527 ) );
  AOI211_X1 us33_U59 (.A( us33_n496 ) , .ZN( us33_n503 ) , .B( us33_n802 ) , .C2( us33_n839 ) , .C1( us33_n851 ) );
  NOR3_X1 us33_U6 (.ZN( us33_n598 ) , .A1( us33_n608 ) , .A3( us33_n723 ) , .A2( us33_n742 ) );
  NAND4_X1 us33_U60 (.ZN( sa30_sr_1 ) , .A4( us33_n595 ) , .A3( us33_n596 ) , .A2( us33_n597 ) , .A1( us33_n598 ) );
  NOR4_X1 us33_U61 (.A4( us33_n591 ) , .A3( us33_n592 ) , .A2( us33_n593 ) , .A1( us33_n594 ) , .ZN( us33_n595 ) );
  AOI211_X1 us33_U62 (.B( us33_n589 ) , .A( us33_n590 ) , .ZN( us33_n596 ) , .C2( us33_n811 ) , .C1( us33_n833 ) );
  AOI211_X1 us33_U63 (.A( us33_n588 ) , .ZN( us33_n597 ) , .B( us33_n621 ) , .C1( us33_n845 ) , .C2( us33_n855 ) );
  NOR2_X1 us33_U64 (.ZN( us33_n748 ) , .A1( us33_n861 ) , .A2( us33_n862 ) );
  NOR2_X1 us33_U65 (.ZN( us33_n625 ) , .A2( us33_n836 ) , .A1( us33_n839 ) );
  NAND4_X1 us33_U66 (.A4( us33_n603 ) , .A3( us33_n604 ) , .A2( us33_n605 ) , .A1( us33_n606 ) , .ZN( us33_n722 ) );
  NOR3_X1 us33_U67 (.A1( us33_n599 ) , .ZN( us33_n604 ) , .A3( us33_n663 ) , .A2( us33_n770 ) );
  NOR4_X1 us33_U68 (.A3( us33_n600 ) , .A2( us33_n601 ) , .A1( us33_n602 ) , .ZN( us33_n603 ) , .A4( us33_n655 ) );
  AOI222_X1 us33_U69 (.ZN( us33_n606 ) , .A1( us33_n830 ) , .C2( us33_n837 ) , .B1( us33_n842 ) , .A2( us33_n856 ) , .B2( us33_n861 ) , .C1( us33_n868 ) );
  NOR3_X1 us33_U7 (.A3( us33_n800 ) , .A2( us33_n801 ) , .A1( us33_n802 ) , .ZN( us33_n825 ) );
  NAND4_X1 us33_U70 (.A4( us33_n657 ) , .A3( us33_n658 ) , .A2( us33_n659 ) , .A1( us33_n660 ) , .ZN( us33_n800 ) );
  NOR3_X1 us33_U71 (.A3( us33_n648 ) , .A2( us33_n649 ) , .A1( us33_n650 ) , .ZN( us33_n659 ) );
  NOR3_X1 us33_U72 (.A3( us33_n651 ) , .A2( us33_n652 ) , .A1( us33_n653 ) , .ZN( us33_n658 ) );
  NOR3_X1 us33_U73 (.A3( us33_n654 ) , .A2( us33_n655 ) , .A1( us33_n656 ) , .ZN( us33_n657 ) );
  NAND4_X1 us33_U74 (.A4( us33_n560 ) , .A3( us33_n561 ) , .A2( us33_n562 ) , .A1( us33_n563 ) , .ZN( us33_n607 ) );
  NOR4_X1 us33_U75 (.ZN( us33_n561 ) , .A1( us33_n653 ) , .A3( us33_n661 ) , .A4( us33_n685 ) , .A2( us33_n768 ) );
  NOR4_X1 us33_U76 (.A4( us33_n552 ) , .A3( us33_n553 ) , .A2( us33_n554 ) , .A1( us33_n555 ) , .ZN( us33_n562 ) );
  NOR4_X1 us33_U77 (.A4( us33_n556 ) , .A3( us33_n557 ) , .A2( us33_n558 ) , .A1( us33_n559 ) , .ZN( us33_n560 ) );
  NAND4_X1 us33_U78 (.A4( us33_n772 ) , .A3( us33_n773 ) , .A2( us33_n774 ) , .A1( us33_n775 ) , .ZN( us33_n801 ) );
  NOR3_X1 us33_U79 (.A3( us33_n765 ) , .A2( us33_n766 ) , .A1( us33_n767 ) , .ZN( us33_n773 ) );
  NOR3_X1 us33_U8 (.A3( us33_n621 ) , .A2( us33_n622 ) , .ZN( us33_n636 ) , .A1( us33_n725 ) );
  NOR4_X1 us33_U80 (.A4( us33_n768 ) , .A3( us33_n769 ) , .A2( us33_n770 ) , .A1( us33_n771 ) , .ZN( us33_n772 ) );
  AOI222_X1 us33_U81 (.ZN( us33_n775 ) , .A1( us33_n830 ) , .C1( us33_n834 ) , .B2( us33_n841 ) , .A2( us33_n850 ) , .B1( us33_n861 ) , .C2( us33_n873 ) );
  NOR4_X1 us33_U82 (.A4( us33_n665 ) , .A3( us33_n666 ) , .A2( us33_n667 ) , .A1( us33_n668 ) , .ZN( us33_n676 ) );
  NOR4_X1 us33_U83 (.A4( us33_n661 ) , .A3( us33_n662 ) , .A2( us33_n663 ) , .A1( us33_n664 ) , .ZN( us33_n677 ) );
  NOR4_X1 us33_U84 (.A3( us33_n673 ) , .A1( us33_n674 ) , .ZN( us33_n675 ) , .A4( us33_n715 ) , .A2( us33_n859 ) );
  NOR2_X1 us33_U85 (.ZN( us33_n761 ) , .A1( us33_n833 ) , .A2( us33_n834 ) );
  NOR4_X1 us33_U86 (.A4( us33_n577 ) , .A3( us33_n578 ) , .A2( us33_n579 ) , .ZN( us33_n586 ) , .A1( us33_n683 ) );
  NOR4_X1 us33_U87 (.A1( us33_n584 ) , .ZN( us33_n585 ) , .A3( us33_n652 ) , .A2( us33_n662 ) , .A4( us33_n767 ) );
  AOI222_X1 us33_U88 (.ZN( us33_n513 ) , .C1( us33_n832 ) , .B2( us33_n837 ) , .A2( us33_n843 ) , .C2( us33_n862 ) , .B1( us33_n863 ) , .A1( us33_n866 ) );
  NOR4_X1 us33_U89 (.A4( us33_n509 ) , .A2( us33_n510 ) , .A1( us33_n511 ) , .ZN( us33_n512 ) , .A3( us33_n670 ) );
  NOR2_X1 us33_U9 (.ZN( us33_n575 ) , .A1( us33_n622 ) , .A2( us33_n745 ) );
  INV_X1 us33_U90 (.A( us33_n505 ) , .ZN( us33_n871 ) );
  NAND4_X1 us33_U91 (.A4( us33_n456 ) , .A3( us33_n457 ) , .A2( us33_n458 ) , .A1( us33_n459 ) , .ZN( us33_n679 ) );
  NOR3_X1 us33_U92 (.ZN( us33_n457 ) , .A3( us33_n530 ) , .A1( us33_n555 ) , .A2( us33_n570 ) );
  AOI221_X1 us33_U93 (.A( us33_n450 ) , .ZN( us33_n459 ) , .C2( us33_n753 ) , .B1( us33_n832 ) , .C1( us33_n842 ) , .B2( us33_n861 ) );
  NOR4_X1 us33_U94 (.ZN( us33_n458 ) , .A2( us33_n509 ) , .A1( us33_n599 ) , .A4( us33_n628 ) , .A3( us33_n711 ) );
  NAND4_X1 us33_U95 (.A4( us33_n535 ) , .A3( us33_n536 ) , .A2( us33_n537 ) , .A1( us33_n538 ) , .ZN( us33_n622 ) );
  NOR4_X1 us33_U96 (.A4( us33_n526 ) , .A2( us33_n527 ) , .A1( us33_n528 ) , .ZN( us33_n538 ) , .A3( us33_n701 ) );
  NOR4_X1 us33_U97 (.A1( us33_n531 ) , .ZN( us33_n536 ) , .A2( us33_n654 ) , .A4( us33_n668 ) , .A3( us33_n765 ) );
  NOR4_X1 us33_U98 (.A4( us33_n529 ) , .A3( us33_n530 ) , .ZN( us33_n537 ) , .A2( us33_n684 ) , .A1( us33_n794 ) );
  NOR2_X1 us33_U99 (.ZN( us33_n647 ) , .A1( us33_n854 ) , .A2( us33_n868 ) );
endmodule

module aes_aes_die_3 ( sa02_0, sa02_1, sa02_2, sa02_3, sa02_4, sa02_5, sa02_6, sa02_7, sa21_0, 
       sa21_1, sa21_2, sa21_3, sa21_4, sa21_5, sa21_6, sa21_7, sa23_0, sa23_1, 
       sa23_2, sa23_3, sa23_4, sa23_5, sa23_6, sa23_7, sa30_0, sa30_1, sa30_2, 
       sa30_3, sa30_4, sa30_5, sa30_6, sa30_7, sa32_0, sa32_1, sa32_2, sa32_3, 
       sa32_4, sa32_5, sa32_6, sa32_7, u0_n268, u0_n270, u0_n272, u0_n274, w3_10, 
       w3_11, w3_8, w3_9, sa02_sr_0, sa02_sr_1, sa02_sr_2, sa02_sr_3, sa02_sr_4, sa02_sr_5, sa02_sr_6, sa02_sr_7, sa21_sr_0, 
        sa21_sr_1, sa21_sr_2, sa21_sr_3, sa21_sr_4, sa21_sr_5, sa21_sr_6, sa21_sr_7, sa23_sr_0, sa23_sr_1, 
        sa23_sr_2, sa23_sr_3, sa23_sr_4, sa23_sr_5, sa23_sr_6, sa23_sr_7, sa31_sr_0, sa31_sr_1, sa31_sr_2, 
        sa31_sr_3, sa31_sr_4, sa31_sr_5, sa31_sr_6, sa31_sr_7, sa33_sr_0, sa33_sr_1, sa33_sr_2, sa33_sr_3, 
        sa33_sr_4, sa33_sr_5, sa33_sr_6, sa33_sr_7, u0_subword_16, u0_subword_17, u0_subword_18, u0_subword_19, u0_subword_20, 
        u0_subword_21, u0_subword_22, u0_subword_23 );
  input sa02_0, sa02_1, sa02_2, sa02_3, sa02_4, sa02_5, sa02_6, sa02_7, sa21_0, 
        sa21_1, sa21_2, sa21_3, sa21_4, sa21_5, sa21_6, sa21_7, sa23_0, sa23_1, 
        sa23_2, sa23_3, sa23_4, sa23_5, sa23_6, sa23_7, sa30_0, sa30_1, sa30_2, 
        sa30_3, sa30_4, sa30_5, sa30_6, sa30_7, sa32_0, sa32_1, sa32_2, sa32_3, 
        sa32_4, sa32_5, sa32_6, sa32_7, u0_n268, u0_n270, u0_n272, u0_n274, w3_10, 
        w3_11, w3_8, w3_9;
  output sa02_sr_0, sa02_sr_1, sa02_sr_2, sa02_sr_3, sa02_sr_4, sa02_sr_5, sa02_sr_6, sa02_sr_7, sa21_sr_0, 
        sa21_sr_1, sa21_sr_2, sa21_sr_3, sa21_sr_4, sa21_sr_5, sa21_sr_6, sa21_sr_7, sa23_sr_0, sa23_sr_1, 
        sa23_sr_2, sa23_sr_3, sa23_sr_4, sa23_sr_5, sa23_sr_6, sa23_sr_7, sa31_sr_0, sa31_sr_1, sa31_sr_2, 
        sa31_sr_3, sa31_sr_4, sa31_sr_5, sa31_sr_6, sa31_sr_7, sa33_sr_0, sa33_sr_1, sa33_sr_2, sa33_sr_3, 
        sa33_sr_4, sa33_sr_5, sa33_sr_6, sa33_sr_7, u0_subword_16, u0_subword_17, u0_subword_18, u0_subword_19, u0_subword_20, 
        u0_subword_21, u0_subword_22, u0_subword_23;
  wire u0_u1_n41, u0_u1_n438, u0_u1_n439, u0_u1_n440, u0_u1_n441, u0_u1_n442, u0_u1_n443, u0_u1_n444, u0_u1_n445, 
       u0_u1_n446, u0_u1_n447, u0_u1_n448, u0_u1_n449, u0_u1_n450, u0_u1_n451, u0_u1_n452, u0_u1_n453, u0_u1_n454, 
       u0_u1_n455, u0_u1_n456, u0_u1_n457, u0_u1_n458, u0_u1_n459, u0_u1_n460, u0_u1_n461, u0_u1_n462, u0_u1_n463, 
       u0_u1_n464, u0_u1_n465, u0_u1_n466, u0_u1_n467, u0_u1_n468, u0_u1_n469, u0_u1_n470, u0_u1_n471, u0_u1_n472, 
       u0_u1_n473, u0_u1_n474, u0_u1_n475, u0_u1_n476, u0_u1_n477, u0_u1_n478, u0_u1_n479, u0_u1_n480, u0_u1_n481, 
       u0_u1_n482, u0_u1_n483, u0_u1_n484, u0_u1_n485, u0_u1_n486, u0_u1_n487, u0_u1_n488, u0_u1_n489, u0_u1_n490, 
       u0_u1_n491, u0_u1_n492, u0_u1_n493, u0_u1_n494, u0_u1_n495, u0_u1_n496, u0_u1_n497, u0_u1_n498, u0_u1_n499, 
       u0_u1_n500, u0_u1_n501, u0_u1_n502, u0_u1_n503, u0_u1_n504, u0_u1_n505, u0_u1_n506, u0_u1_n507, u0_u1_n508, 
       u0_u1_n509, u0_u1_n510, u0_u1_n511, u0_u1_n512, u0_u1_n513, u0_u1_n514, u0_u1_n515, u0_u1_n516, u0_u1_n517, 
       u0_u1_n518, u0_u1_n519, u0_u1_n520, u0_u1_n521, u0_u1_n522, u0_u1_n523, u0_u1_n524, u0_u1_n525, u0_u1_n526, 
       u0_u1_n527, u0_u1_n528, u0_u1_n529, u0_u1_n530, u0_u1_n531, u0_u1_n532, u0_u1_n533, u0_u1_n534, u0_u1_n535, 
       u0_u1_n536, u0_u1_n537, u0_u1_n538, u0_u1_n539, u0_u1_n540, u0_u1_n541, u0_u1_n542, u0_u1_n543, u0_u1_n544, 
       u0_u1_n545, u0_u1_n546, u0_u1_n547, u0_u1_n548, u0_u1_n549, u0_u1_n550, u0_u1_n551, u0_u1_n552, u0_u1_n553, 
       u0_u1_n554, u0_u1_n555, u0_u1_n556, u0_u1_n557, u0_u1_n558, u0_u1_n559, u0_u1_n560, u0_u1_n561, u0_u1_n562, 
       u0_u1_n563, u0_u1_n564, u0_u1_n565, u0_u1_n566, u0_u1_n567, u0_u1_n568, u0_u1_n569, u0_u1_n570, u0_u1_n571, 
       u0_u1_n572, u0_u1_n573, u0_u1_n574, u0_u1_n575, u0_u1_n576, u0_u1_n577, u0_u1_n578, u0_u1_n579, u0_u1_n580, 
       u0_u1_n581, u0_u1_n582, u0_u1_n583, u0_u1_n584, u0_u1_n585, u0_u1_n586, u0_u1_n587, u0_u1_n588, u0_u1_n589, 
       u0_u1_n590, u0_u1_n591, u0_u1_n592, u0_u1_n593, u0_u1_n594, u0_u1_n595, u0_u1_n596, u0_u1_n597, u0_u1_n598, 
       u0_u1_n599, u0_u1_n600, u0_u1_n601, u0_u1_n602, u0_u1_n603, u0_u1_n604, u0_u1_n605, u0_u1_n606, u0_u1_n607, 
       u0_u1_n608, u0_u1_n609, u0_u1_n610, u0_u1_n611, u0_u1_n612, u0_u1_n613, u0_u1_n614, u0_u1_n615, u0_u1_n616, 
       u0_u1_n617, u0_u1_n618, u0_u1_n619, u0_u1_n620, u0_u1_n621, u0_u1_n622, u0_u1_n623, u0_u1_n624, u0_u1_n625, 
       u0_u1_n626, u0_u1_n627, u0_u1_n628, u0_u1_n629, u0_u1_n630, u0_u1_n631, u0_u1_n632, u0_u1_n633, u0_u1_n634, 
       u0_u1_n635, u0_u1_n636, u0_u1_n637, u0_u1_n638, u0_u1_n639, u0_u1_n640, u0_u1_n641, u0_u1_n642, u0_u1_n643, 
       u0_u1_n644, u0_u1_n645, u0_u1_n646, u0_u1_n647, u0_u1_n648, u0_u1_n649, u0_u1_n650, u0_u1_n651, u0_u1_n652, 
       u0_u1_n653, u0_u1_n654, u0_u1_n655, u0_u1_n656, u0_u1_n657, u0_u1_n658, u0_u1_n659, u0_u1_n660, u0_u1_n661, 
       u0_u1_n662, u0_u1_n663, u0_u1_n664, u0_u1_n665, u0_u1_n666, u0_u1_n667, u0_u1_n668, u0_u1_n669, u0_u1_n670, 
       u0_u1_n671, u0_u1_n672, u0_u1_n673, u0_u1_n674, u0_u1_n675, u0_u1_n676, u0_u1_n677, u0_u1_n678, u0_u1_n679, 
       u0_u1_n680, u0_u1_n681, u0_u1_n682, u0_u1_n683, u0_u1_n684, u0_u1_n685, u0_u1_n686, u0_u1_n687, u0_u1_n688, 
       u0_u1_n689, u0_u1_n690, u0_u1_n691, u0_u1_n692, u0_u1_n693, u0_u1_n694, u0_u1_n695, u0_u1_n696, u0_u1_n697, 
       u0_u1_n698, u0_u1_n699, u0_u1_n700, u0_u1_n701, u0_u1_n702, u0_u1_n703, u0_u1_n704, u0_u1_n705, u0_u1_n706, 
       u0_u1_n707, u0_u1_n708, u0_u1_n709, u0_u1_n710, u0_u1_n711, u0_u1_n712, u0_u1_n713, u0_u1_n714, u0_u1_n715, 
       u0_u1_n716, u0_u1_n717, u0_u1_n718, u0_u1_n719, u0_u1_n720, u0_u1_n721, u0_u1_n722, u0_u1_n723, u0_u1_n724, 
       u0_u1_n725, u0_u1_n726, u0_u1_n727, u0_u1_n728, u0_u1_n729, u0_u1_n730, u0_u1_n731, u0_u1_n732, u0_u1_n733, 
       u0_u1_n734, u0_u1_n735, u0_u1_n736, u0_u1_n737, u0_u1_n738, u0_u1_n739, u0_u1_n740, u0_u1_n741, u0_u1_n742, 
       u0_u1_n743, u0_u1_n744, u0_u1_n745, u0_u1_n746, u0_u1_n747, u0_u1_n748, u0_u1_n749, u0_u1_n750, u0_u1_n751, 
       u0_u1_n752, u0_u1_n753, u0_u1_n754, u0_u1_n755, u0_u1_n756, u0_u1_n757, u0_u1_n758, u0_u1_n759, u0_u1_n760, 
       u0_u1_n761, u0_u1_n762, u0_u1_n763, u0_u1_n764, u0_u1_n765, u0_u1_n766, u0_u1_n767, u0_u1_n768, u0_u1_n769, 
       u0_u1_n770, u0_u1_n771, u0_u1_n772, u0_u1_n773, u0_u1_n774, u0_u1_n775, u0_u1_n776, u0_u1_n777, u0_u1_n778, 
       u0_u1_n779, u0_u1_n780, u0_u1_n781, u0_u1_n782, u0_u1_n783, u0_u1_n784, u0_u1_n785, u0_u1_n786, u0_u1_n787, 
       u0_u1_n788, u0_u1_n789, u0_u1_n790, u0_u1_n791, u0_u1_n792, u0_u1_n793, u0_u1_n794, u0_u1_n795, u0_u1_n796, 
       u0_u1_n797, u0_u1_n798, u0_u1_n799, u0_u1_n800, u0_u1_n801, u0_u1_n802, u0_u1_n803, u0_u1_n804, u0_u1_n805, 
       u0_u1_n806, u0_u1_n807, u0_u1_n808, u0_u1_n809, u0_u1_n810, u0_u1_n811, u0_u1_n812, u0_u1_n813, u0_u1_n814, 
       u0_u1_n815, u0_u1_n816, u0_u1_n817, u0_u1_n818, u0_u1_n819, u0_u1_n820, u0_u1_n821, u0_u1_n822, u0_u1_n823, 
       u0_u1_n824, u0_u1_n825, u0_u1_n826, u0_u1_n827, u0_u1_n828, u0_u1_n829, u0_u1_n830, u0_u1_n831, u0_u1_n832, 
       u0_u1_n833, u0_u1_n834, u0_u1_n835, u0_u1_n836, u0_u1_n837, u0_u1_n838, u0_u1_n839, u0_u1_n840, u0_u1_n841, 
       u0_u1_n842, u0_u1_n843, u0_u1_n844, u0_u1_n845, u0_u1_n846, u0_u1_n847, u0_u1_n848, u0_u1_n849, u0_u1_n850, 
       u0_u1_n851, u0_u1_n852, u0_u1_n853, u0_u1_n854, u0_u1_n855, u0_u1_n856, u0_u1_n857, u0_u1_n858, u0_u1_n859, 
       u0_u1_n860, u0_u1_n861, u0_u1_n862, u0_u1_n863, u0_u1_n864, u0_u1_n865, u0_u1_n866, u0_u1_n867, u0_u1_n868, 
       u0_u1_n869, u0_u1_n870, u0_u1_n871, u0_u1_n872, u0_u1_n873, u0_u1_n874, u0_u1_n875, u0_u1_n876, u0_u1_n877, 
       us02_n438, us02_n439, us02_n440, us02_n441, us02_n442, us02_n443, us02_n444, us02_n445, us02_n446, 
       us02_n447, us02_n448, us02_n449, us02_n450, us02_n451, us02_n452, us02_n453, us02_n454, us02_n455, 
       us02_n456, us02_n457, us02_n458, us02_n459, us02_n460, us02_n461, us02_n462, us02_n463, us02_n464, 
       us02_n465, us02_n466, us02_n467, us02_n468, us02_n469, us02_n470, us02_n471, us02_n472, us02_n473, 
       us02_n474, us02_n475, us02_n476, us02_n477, us02_n478, us02_n479, us02_n480, us02_n481, us02_n482, 
       us02_n483, us02_n484, us02_n485, us02_n486, us02_n487, us02_n488, us02_n489, us02_n490, us02_n491, 
       us02_n492, us02_n493, us02_n494, us02_n495, us02_n496, us02_n497, us02_n498, us02_n499, us02_n500, 
       us02_n501, us02_n502, us02_n503, us02_n504, us02_n505, us02_n506, us02_n507, us02_n508, us02_n509, 
       us02_n510, us02_n511, us02_n512, us02_n513, us02_n514, us02_n515, us02_n516, us02_n517, us02_n518, 
       us02_n519, us02_n520, us02_n521, us02_n522, us02_n523, us02_n524, us02_n525, us02_n526, us02_n527, 
       us02_n528, us02_n529, us02_n530, us02_n531, us02_n532, us02_n533, us02_n534, us02_n535, us02_n536, 
       us02_n537, us02_n538, us02_n539, us02_n540, us02_n541, us02_n542, us02_n543, us02_n544, us02_n545, 
       us02_n546, us02_n547, us02_n548, us02_n549, us02_n550, us02_n551, us02_n552, us02_n553, us02_n554, 
       us02_n555, us02_n556, us02_n557, us02_n558, us02_n559, us02_n560, us02_n561, us02_n562, us02_n563, 
       us02_n564, us02_n565, us02_n566, us02_n567, us02_n568, us02_n569, us02_n570, us02_n571, us02_n572, 
       us02_n573, us02_n574, us02_n575, us02_n576, us02_n577, us02_n578, us02_n579, us02_n580, us02_n581, 
       us02_n582, us02_n583, us02_n584, us02_n585, us02_n586, us02_n587, us02_n588, us02_n589, us02_n590, 
       us02_n591, us02_n592, us02_n593, us02_n594, us02_n595, us02_n596, us02_n597, us02_n598, us02_n599, 
       us02_n600, us02_n601, us02_n602, us02_n603, us02_n604, us02_n605, us02_n606, us02_n607, us02_n608, 
       us02_n609, us02_n610, us02_n611, us02_n612, us02_n613, us02_n614, us02_n615, us02_n616, us02_n617, 
       us02_n618, us02_n619, us02_n620, us02_n621, us02_n622, us02_n623, us02_n624, us02_n625, us02_n626, 
       us02_n627, us02_n628, us02_n629, us02_n630, us02_n631, us02_n632, us02_n633, us02_n634, us02_n635, 
       us02_n636, us02_n637, us02_n638, us02_n639, us02_n640, us02_n641, us02_n642, us02_n643, us02_n644, 
       us02_n645, us02_n646, us02_n647, us02_n648, us02_n649, us02_n650, us02_n651, us02_n652, us02_n653, 
       us02_n654, us02_n655, us02_n656, us02_n657, us02_n658, us02_n659, us02_n660, us02_n661, us02_n662, 
       us02_n663, us02_n664, us02_n665, us02_n666, us02_n667, us02_n668, us02_n669, us02_n670, us02_n671, 
       us02_n672, us02_n673, us02_n674, us02_n675, us02_n676, us02_n677, us02_n678, us02_n679, us02_n680, 
       us02_n681, us02_n682, us02_n683, us02_n684, us02_n685, us02_n686, us02_n687, us02_n688, us02_n689, 
       us02_n690, us02_n691, us02_n692, us02_n693, us02_n694, us02_n695, us02_n696, us02_n697, us02_n698, 
       us02_n699, us02_n700, us02_n701, us02_n702, us02_n703, us02_n704, us02_n705, us02_n706, us02_n707, 
       us02_n708, us02_n709, us02_n710, us02_n711, us02_n712, us02_n713, us02_n714, us02_n715, us02_n716, 
       us02_n717, us02_n718, us02_n719, us02_n720, us02_n721, us02_n722, us02_n723, us02_n724, us02_n725, 
       us02_n726, us02_n727, us02_n728, us02_n729, us02_n730, us02_n731, us02_n732, us02_n733, us02_n734, 
       us02_n735, us02_n736, us02_n737, us02_n738, us02_n739, us02_n740, us02_n741, us02_n742, us02_n743, 
       us02_n744, us02_n745, us02_n746, us02_n747, us02_n748, us02_n749, us02_n750, us02_n751, us02_n752, 
       us02_n753, us02_n754, us02_n755, us02_n756, us02_n757, us02_n758, us02_n759, us02_n760, us02_n761, 
       us02_n762, us02_n763, us02_n764, us02_n765, us02_n766, us02_n767, us02_n768, us02_n769, us02_n770, 
       us02_n771, us02_n772, us02_n773, us02_n774, us02_n775, us02_n776, us02_n777, us02_n778, us02_n779, 
       us02_n780, us02_n781, us02_n782, us02_n783, us02_n784, us02_n785, us02_n786, us02_n787, us02_n788, 
       us02_n789, us02_n790, us02_n791, us02_n792, us02_n793, us02_n794, us02_n795, us02_n796, us02_n797, 
       us02_n798, us02_n799, us02_n800, us02_n801, us02_n802, us02_n803, us02_n804, us02_n805, us02_n806, 
       us02_n807, us02_n808, us02_n809, us02_n810, us02_n811, us02_n812, us02_n813, us02_n814, us02_n815, 
       us02_n816, us02_n817, us02_n818, us02_n819, us02_n820, us02_n821, us02_n822, us02_n823, us02_n824, 
       us02_n825, us02_n826, us02_n827, us02_n828, us02_n829, us02_n830, us02_n831, us02_n832, us02_n833, 
       us02_n834, us02_n835, us02_n836, us02_n837, us02_n838, us02_n839, us02_n840, us02_n841, us02_n842, 
       us02_n843, us02_n844, us02_n845, us02_n846, us02_n847, us02_n848, us02_n849, us02_n850, us02_n851, 
       us02_n852, us02_n853, us02_n854, us02_n855, us02_n856, us02_n857, us02_n858, us02_n859, us02_n860, 
       us02_n861, us02_n862, us02_n863, us02_n864, us02_n865, us02_n866, us02_n867, us02_n868, us02_n869, 
       us02_n870, us02_n871, us02_n872, us02_n873, us02_n874, us02_n875, us21_n438, us21_n439, us21_n440, 
       us21_n441, us21_n442, us21_n443, us21_n444, us21_n445, us21_n446, us21_n447, us21_n448, us21_n449, 
       us21_n450, us21_n451, us21_n452, us21_n453, us21_n454, us21_n455, us21_n456, us21_n457, us21_n458, 
       us21_n459, us21_n460, us21_n461, us21_n462, us21_n463, us21_n464, us21_n465, us21_n466, us21_n467, 
       us21_n468, us21_n469, us21_n470, us21_n471, us21_n472, us21_n473, us21_n474, us21_n475, us21_n476, 
       us21_n477, us21_n478, us21_n479, us21_n480, us21_n481, us21_n482, us21_n483, us21_n484, us21_n485, 
       us21_n486, us21_n487, us21_n488, us21_n489, us21_n490, us21_n491, us21_n492, us21_n493, us21_n494, 
       us21_n495, us21_n496, us21_n497, us21_n498, us21_n499, us21_n500, us21_n501, us21_n502, us21_n503, 
       us21_n504, us21_n505, us21_n506, us21_n507, us21_n508, us21_n509, us21_n510, us21_n511, us21_n512, 
       us21_n513, us21_n514, us21_n515, us21_n516, us21_n517, us21_n518, us21_n519, us21_n520, us21_n521, 
       us21_n522, us21_n523, us21_n524, us21_n525, us21_n526, us21_n527, us21_n528, us21_n529, us21_n530, 
       us21_n531, us21_n532, us21_n533, us21_n534, us21_n535, us21_n536, us21_n537, us21_n538, us21_n539, 
       us21_n540, us21_n541, us21_n542, us21_n543, us21_n544, us21_n545, us21_n546, us21_n547, us21_n548, 
       us21_n549, us21_n550, us21_n551, us21_n552, us21_n553, us21_n554, us21_n555, us21_n556, us21_n557, 
       us21_n558, us21_n559, us21_n560, us21_n561, us21_n562, us21_n563, us21_n564, us21_n565, us21_n566, 
       us21_n567, us21_n568, us21_n569, us21_n570, us21_n571, us21_n572, us21_n573, us21_n574, us21_n575, 
       us21_n576, us21_n577, us21_n578, us21_n579, us21_n580, us21_n581, us21_n582, us21_n583, us21_n584, 
       us21_n585, us21_n586, us21_n587, us21_n588, us21_n589, us21_n590, us21_n591, us21_n592, us21_n593, 
       us21_n594, us21_n595, us21_n596, us21_n597, us21_n598, us21_n599, us21_n600, us21_n601, us21_n602, 
       us21_n603, us21_n604, us21_n605, us21_n606, us21_n607, us21_n608, us21_n609, us21_n610, us21_n611, 
       us21_n612, us21_n613, us21_n614, us21_n615, us21_n616, us21_n617, us21_n618, us21_n619, us21_n620, 
       us21_n621, us21_n622, us21_n623, us21_n624, us21_n625, us21_n626, us21_n627, us21_n628, us21_n629, 
       us21_n630, us21_n631, us21_n632, us21_n633, us21_n634, us21_n635, us21_n636, us21_n637, us21_n638, 
       us21_n639, us21_n640, us21_n641, us21_n642, us21_n643, us21_n644, us21_n645, us21_n646, us21_n647, 
       us21_n648, us21_n649, us21_n650, us21_n651, us21_n652, us21_n653, us21_n654, us21_n655, us21_n656, 
       us21_n657, us21_n658, us21_n659, us21_n660, us21_n661, us21_n662, us21_n663, us21_n664, us21_n665, 
       us21_n666, us21_n667, us21_n668, us21_n669, us21_n670, us21_n671, us21_n672, us21_n673, us21_n674, 
       us21_n675, us21_n676, us21_n677, us21_n678, us21_n679, us21_n680, us21_n681, us21_n682, us21_n683, 
       us21_n684, us21_n685, us21_n686, us21_n687, us21_n688, us21_n689, us21_n690, us21_n691, us21_n692, 
       us21_n693, us21_n694, us21_n695, us21_n696, us21_n697, us21_n698, us21_n699, us21_n700, us21_n701, 
       us21_n702, us21_n703, us21_n704, us21_n705, us21_n706, us21_n707, us21_n708, us21_n709, us21_n710, 
       us21_n711, us21_n712, us21_n713, us21_n714, us21_n715, us21_n716, us21_n717, us21_n718, us21_n719, 
       us21_n720, us21_n721, us21_n722, us21_n723, us21_n724, us21_n725, us21_n726, us21_n727, us21_n728, 
       us21_n729, us21_n730, us21_n731, us21_n732, us21_n733, us21_n734, us21_n735, us21_n736, us21_n737, 
       us21_n738, us21_n739, us21_n740, us21_n741, us21_n742, us21_n743, us21_n744, us21_n745, us21_n746, 
       us21_n747, us21_n748, us21_n749, us21_n750, us21_n751, us21_n752, us21_n753, us21_n754, us21_n755, 
       us21_n756, us21_n757, us21_n758, us21_n759, us21_n760, us21_n761, us21_n762, us21_n763, us21_n764, 
       us21_n765, us21_n766, us21_n767, us21_n768, us21_n769, us21_n770, us21_n771, us21_n772, us21_n773, 
       us21_n774, us21_n775, us21_n776, us21_n777, us21_n778, us21_n779, us21_n780, us21_n781, us21_n782, 
       us21_n783, us21_n784, us21_n785, us21_n786, us21_n787, us21_n788, us21_n789, us21_n790, us21_n791, 
       us21_n792, us21_n793, us21_n794, us21_n795, us21_n796, us21_n797, us21_n798, us21_n799, us21_n800, 
       us21_n801, us21_n802, us21_n803, us21_n804, us21_n805, us21_n806, us21_n807, us21_n808, us21_n809, 
       us21_n810, us21_n811, us21_n812, us21_n813, us21_n814, us21_n815, us21_n816, us21_n817, us21_n818, 
       us21_n819, us21_n820, us21_n821, us21_n822, us21_n823, us21_n824, us21_n825, us21_n826, us21_n827, 
       us21_n828, us21_n829, us21_n830, us21_n831, us21_n832, us21_n833, us21_n834, us21_n835, us21_n836, 
       us21_n837, us21_n838, us21_n839, us21_n840, us21_n841, us21_n842, us21_n843, us21_n844, us21_n845, 
       us21_n846, us21_n847, us21_n848, us21_n849, us21_n850, us21_n851, us21_n852, us21_n853, us21_n854, 
       us21_n855, us21_n856, us21_n857, us21_n858, us21_n859, us21_n860, us21_n861, us21_n862, us21_n863, 
       us21_n864, us21_n865, us21_n866, us21_n867, us21_n868, us21_n869, us21_n870, us21_n871, us21_n872, 
       us21_n873, us21_n874, us23_n438, us23_n439, us23_n440, us23_n441, us23_n442, us23_n443, us23_n444, 
       us23_n445, us23_n446, us23_n447, us23_n448, us23_n449, us23_n450, us23_n451, us23_n452, us23_n453, 
       us23_n454, us23_n455, us23_n456, us23_n457, us23_n458, us23_n459, us23_n460, us23_n461, us23_n462, 
       us23_n463, us23_n464, us23_n465, us23_n466, us23_n467, us23_n468, us23_n469, us23_n470, us23_n471, 
       us23_n472, us23_n473, us23_n474, us23_n475, us23_n476, us23_n477, us23_n478, us23_n479, us23_n480, 
       us23_n481, us23_n482, us23_n483, us23_n484, us23_n485, us23_n486, us23_n487, us23_n488, us23_n489, 
       us23_n490, us23_n491, us23_n492, us23_n493, us23_n494, us23_n495, us23_n496, us23_n497, us23_n498, 
       us23_n499, us23_n500, us23_n501, us23_n502, us23_n503, us23_n504, us23_n505, us23_n506, us23_n507, 
       us23_n508, us23_n509, us23_n510, us23_n511, us23_n512, us23_n513, us23_n514, us23_n515, us23_n516, 
       us23_n517, us23_n518, us23_n519, us23_n520, us23_n521, us23_n522, us23_n523, us23_n524, us23_n525, 
       us23_n526, us23_n527, us23_n528, us23_n529, us23_n530, us23_n531, us23_n532, us23_n533, us23_n534, 
       us23_n535, us23_n536, us23_n537, us23_n538, us23_n539, us23_n540, us23_n541, us23_n542, us23_n543, 
       us23_n544, us23_n545, us23_n546, us23_n547, us23_n548, us23_n549, us23_n550, us23_n551, us23_n552, 
       us23_n553, us23_n554, us23_n555, us23_n556, us23_n557, us23_n558, us23_n559, us23_n560, us23_n561, 
       us23_n562, us23_n563, us23_n564, us23_n565, us23_n566, us23_n567, us23_n568, us23_n569, us23_n570, 
       us23_n571, us23_n572, us23_n573, us23_n574, us23_n575, us23_n576, us23_n577, us23_n578, us23_n579, 
       us23_n580, us23_n581, us23_n582, us23_n583, us23_n584, us23_n585, us23_n586, us23_n587, us23_n588, 
       us23_n589, us23_n590, us23_n591, us23_n592, us23_n593, us23_n594, us23_n595, us23_n596, us23_n597, 
       us23_n598, us23_n599, us23_n600, us23_n601, us23_n602, us23_n603, us23_n604, us23_n605, us23_n606, 
       us23_n607, us23_n608, us23_n609, us23_n610, us23_n611, us23_n612, us23_n613, us23_n614, us23_n615, 
       us23_n616, us23_n617, us23_n618, us23_n619, us23_n620, us23_n621, us23_n622, us23_n623, us23_n624, 
       us23_n625, us23_n626, us23_n627, us23_n628, us23_n629, us23_n630, us23_n631, us23_n632, us23_n633, 
       us23_n634, us23_n635, us23_n636, us23_n637, us23_n638, us23_n639, us23_n640, us23_n641, us23_n642, 
       us23_n643, us23_n644, us23_n645, us23_n646, us23_n647, us23_n648, us23_n649, us23_n650, us23_n651, 
       us23_n652, us23_n653, us23_n654, us23_n655, us23_n656, us23_n657, us23_n658, us23_n659, us23_n660, 
       us23_n661, us23_n662, us23_n663, us23_n664, us23_n665, us23_n666, us23_n667, us23_n668, us23_n669, 
       us23_n670, us23_n671, us23_n672, us23_n673, us23_n674, us23_n675, us23_n676, us23_n677, us23_n678, 
       us23_n679, us23_n680, us23_n681, us23_n682, us23_n683, us23_n684, us23_n685, us23_n686, us23_n687, 
       us23_n688, us23_n689, us23_n690, us23_n691, us23_n692, us23_n693, us23_n694, us23_n695, us23_n696, 
       us23_n697, us23_n698, us23_n699, us23_n700, us23_n701, us23_n702, us23_n703, us23_n704, us23_n705, 
       us23_n706, us23_n707, us23_n708, us23_n709, us23_n710, us23_n711, us23_n712, us23_n713, us23_n714, 
       us23_n715, us23_n716, us23_n717, us23_n718, us23_n719, us23_n720, us23_n721, us23_n722, us23_n723, 
       us23_n724, us23_n725, us23_n726, us23_n727, us23_n728, us23_n729, us23_n730, us23_n731, us23_n732, 
       us23_n733, us23_n734, us23_n735, us23_n736, us23_n737, us23_n738, us23_n739, us23_n740, us23_n741, 
       us23_n742, us23_n743, us23_n744, us23_n745, us23_n746, us23_n747, us23_n748, us23_n749, us23_n750, 
       us23_n751, us23_n752, us23_n753, us23_n754, us23_n755, us23_n756, us23_n757, us23_n758, us23_n759, 
       us23_n760, us23_n761, us23_n762, us23_n763, us23_n764, us23_n765, us23_n766, us23_n767, us23_n768, 
       us23_n769, us23_n770, us23_n771, us23_n772, us23_n773, us23_n774, us23_n775, us23_n776, us23_n777, 
       us23_n778, us23_n779, us23_n780, us23_n781, us23_n782, us23_n783, us23_n784, us23_n785, us23_n786, 
       us23_n787, us23_n788, us23_n789, us23_n790, us23_n791, us23_n792, us23_n793, us23_n794, us23_n795, 
       us23_n796, us23_n797, us23_n798, us23_n799, us23_n800, us23_n801, us23_n802, us23_n803, us23_n804, 
       us23_n805, us23_n806, us23_n807, us23_n808, us23_n809, us23_n810, us23_n811, us23_n812, us23_n813, 
       us23_n814, us23_n815, us23_n816, us23_n817, us23_n818, us23_n819, us23_n820, us23_n821, us23_n822, 
       us23_n823, us23_n824, us23_n825, us23_n826, us23_n827, us23_n828, us23_n829, us23_n830, us23_n831, 
       us23_n832, us23_n833, us23_n834, us23_n835, us23_n836, us23_n837, us23_n838, us23_n839, us23_n840, 
       us23_n841, us23_n842, us23_n843, us23_n844, us23_n845, us23_n846, us23_n847, us23_n848, us23_n849, 
       us23_n850, us23_n851, us23_n852, us23_n853, us23_n854, us23_n855, us23_n856, us23_n857, us23_n858, 
       us23_n859, us23_n860, us23_n861, us23_n862, us23_n863, us23_n864, us23_n865, us23_n866, us23_n867, 
       us23_n868, us23_n869, us23_n870, us23_n871, us23_n872, us23_n873, us23_n874, us23_n875, us30_n438, 
       us30_n439, us30_n440, us30_n441, us30_n442, us30_n443, us30_n444, us30_n445, us30_n446, us30_n447, 
       us30_n448, us30_n449, us30_n450, us30_n451, us30_n452, us30_n453, us30_n454, us30_n455, us30_n456, 
       us30_n457, us30_n458, us30_n459, us30_n460, us30_n461, us30_n462, us30_n463, us30_n464, us30_n465, 
       us30_n466, us30_n467, us30_n468, us30_n469, us30_n470, us30_n471, us30_n472, us30_n473, us30_n474, 
       us30_n475, us30_n476, us30_n477, us30_n478, us30_n479, us30_n480, us30_n481, us30_n482, us30_n483, 
       us30_n484, us30_n485, us30_n486, us30_n487, us30_n488, us30_n489, us30_n490, us30_n491, us30_n492, 
       us30_n493, us30_n494, us30_n495, us30_n496, us30_n497, us30_n498, us30_n499, us30_n500, us30_n501, 
       us30_n502, us30_n503, us30_n504, us30_n505, us30_n506, us30_n507, us30_n508, us30_n509, us30_n510, 
       us30_n511, us30_n512, us30_n513, us30_n514, us30_n515, us30_n516, us30_n517, us30_n518, us30_n519, 
       us30_n520, us30_n521, us30_n522, us30_n523, us30_n524, us30_n525, us30_n526, us30_n527, us30_n528, 
       us30_n529, us30_n530, us30_n531, us30_n532, us30_n533, us30_n534, us30_n535, us30_n536, us30_n537, 
       us30_n538, us30_n539, us30_n540, us30_n541, us30_n542, us30_n543, us30_n544, us30_n545, us30_n546, 
       us30_n547, us30_n548, us30_n549, us30_n550, us30_n551, us30_n552, us30_n553, us30_n554, us30_n555, 
       us30_n556, us30_n557, us30_n558, us30_n559, us30_n560, us30_n561, us30_n562, us30_n563, us30_n564, 
       us30_n565, us30_n566, us30_n567, us30_n568, us30_n569, us30_n570, us30_n571, us30_n572, us30_n573, 
       us30_n574, us30_n575, us30_n576, us30_n577, us30_n578, us30_n579, us30_n580, us30_n581, us30_n582, 
       us30_n583, us30_n584, us30_n585, us30_n586, us30_n587, us30_n588, us30_n589, us30_n590, us30_n591, 
       us30_n592, us30_n593, us30_n594, us30_n595, us30_n596, us30_n597, us30_n598, us30_n599, us30_n600, 
       us30_n601, us30_n602, us30_n603, us30_n604, us30_n605, us30_n606, us30_n607, us30_n608, us30_n609, 
       us30_n610, us30_n611, us30_n612, us30_n613, us30_n614, us30_n615, us30_n616, us30_n617, us30_n618, 
       us30_n619, us30_n620, us30_n621, us30_n622, us30_n623, us30_n624, us30_n625, us30_n626, us30_n627, 
       us30_n628, us30_n629, us30_n630, us30_n631, us30_n632, us30_n633, us30_n634, us30_n635, us30_n636, 
       us30_n637, us30_n638, us30_n639, us30_n640, us30_n641, us30_n642, us30_n643, us30_n644, us30_n645, 
       us30_n646, us30_n647, us30_n648, us30_n649, us30_n650, us30_n651, us30_n652, us30_n653, us30_n654, 
       us30_n655, us30_n656, us30_n657, us30_n658, us30_n659, us30_n660, us30_n661, us30_n662, us30_n663, 
       us30_n664, us30_n665, us30_n666, us30_n667, us30_n668, us30_n669, us30_n670, us30_n671, us30_n672, 
       us30_n673, us30_n674, us30_n675, us30_n676, us30_n677, us30_n678, us30_n679, us30_n680, us30_n681, 
       us30_n682, us30_n683, us30_n684, us30_n685, us30_n686, us30_n687, us30_n688, us30_n689, us30_n690, 
       us30_n691, us30_n692, us30_n693, us30_n694, us30_n695, us30_n696, us30_n697, us30_n698, us30_n699, 
       us30_n700, us30_n701, us30_n702, us30_n703, us30_n704, us30_n705, us30_n706, us30_n707, us30_n708, 
       us30_n709, us30_n710, us30_n711, us30_n712, us30_n713, us30_n714, us30_n715, us30_n716, us30_n717, 
       us30_n718, us30_n719, us30_n720, us30_n721, us30_n722, us30_n723, us30_n724, us30_n725, us30_n726, 
       us30_n727, us30_n728, us30_n729, us30_n730, us30_n731, us30_n732, us30_n733, us30_n734, us30_n735, 
       us30_n736, us30_n737, us30_n738, us30_n739, us30_n740, us30_n741, us30_n742, us30_n743, us30_n744, 
       us30_n745, us30_n746, us30_n747, us30_n748, us30_n749, us30_n750, us30_n751, us30_n752, us30_n753, 
       us30_n754, us30_n755, us30_n756, us30_n757, us30_n758, us30_n759, us30_n760, us30_n761, us30_n762, 
       us30_n763, us30_n764, us30_n765, us30_n766, us30_n767, us30_n768, us30_n769, us30_n770, us30_n771, 
       us30_n772, us30_n773, us30_n774, us30_n775, us30_n776, us30_n777, us30_n778, us30_n779, us30_n780, 
       us30_n781, us30_n782, us30_n783, us30_n784, us30_n785, us30_n786, us30_n787, us30_n788, us30_n789, 
       us30_n790, us30_n791, us30_n792, us30_n793, us30_n794, us30_n795, us30_n796, us30_n797, us30_n798, 
       us30_n799, us30_n800, us30_n801, us30_n802, us30_n803, us30_n804, us30_n805, us30_n806, us30_n807, 
       us30_n808, us30_n809, us30_n810, us30_n811, us30_n812, us30_n813, us30_n814, us30_n815, us30_n816, 
       us30_n817, us30_n818, us30_n819, us30_n820, us30_n821, us30_n822, us30_n823, us30_n824, us30_n825, 
       us30_n826, us30_n827, us30_n828, us30_n829, us30_n830, us30_n831, us30_n832, us30_n833, us30_n834, 
       us30_n835, us30_n836, us30_n837, us30_n838, us30_n839, us30_n840, us30_n841, us30_n842, us30_n843, 
       us30_n844, us30_n845, us30_n846, us30_n847, us30_n848, us30_n849, us30_n850, us30_n851, us30_n852, 
       us30_n853, us30_n854, us30_n855, us30_n856, us30_n857, us30_n858, us30_n859, us30_n860, us30_n861, 
       us30_n862, us30_n863, us30_n864, us30_n865, us30_n866, us30_n867, us30_n868, us30_n869, us30_n870, 
       us30_n871, us30_n872, us30_n873, us30_n874, us30_n875, us30_n876, us32_n438, us32_n439, us32_n440, 
       us32_n441, us32_n442, us32_n443, us32_n444, us32_n445, us32_n446, us32_n447, us32_n448, us32_n449, 
       us32_n450, us32_n451, us32_n452, us32_n453, us32_n454, us32_n455, us32_n456, us32_n457, us32_n458, 
       us32_n459, us32_n460, us32_n461, us32_n462, us32_n463, us32_n464, us32_n465, us32_n466, us32_n467, 
       us32_n468, us32_n469, us32_n470, us32_n471, us32_n472, us32_n473, us32_n474, us32_n475, us32_n476, 
       us32_n477, us32_n478, us32_n479, us32_n480, us32_n481, us32_n482, us32_n483, us32_n484, us32_n485, 
       us32_n486, us32_n487, us32_n488, us32_n489, us32_n490, us32_n491, us32_n492, us32_n493, us32_n494, 
       us32_n495, us32_n496, us32_n497, us32_n498, us32_n499, us32_n500, us32_n501, us32_n502, us32_n503, 
       us32_n504, us32_n505, us32_n506, us32_n507, us32_n508, us32_n509, us32_n510, us32_n511, us32_n512, 
       us32_n513, us32_n514, us32_n515, us32_n516, us32_n517, us32_n518, us32_n519, us32_n520, us32_n521, 
       us32_n522, us32_n523, us32_n524, us32_n525, us32_n526, us32_n527, us32_n528, us32_n529, us32_n530, 
       us32_n531, us32_n532, us32_n533, us32_n534, us32_n535, us32_n536, us32_n537, us32_n538, us32_n539, 
       us32_n540, us32_n541, us32_n542, us32_n543, us32_n544, us32_n545, us32_n546, us32_n547, us32_n548, 
       us32_n549, us32_n550, us32_n551, us32_n552, us32_n553, us32_n554, us32_n555, us32_n556, us32_n557, 
       us32_n558, us32_n559, us32_n560, us32_n561, us32_n562, us32_n563, us32_n564, us32_n565, us32_n566, 
       us32_n567, us32_n568, us32_n569, us32_n570, us32_n571, us32_n572, us32_n573, us32_n574, us32_n575, 
       us32_n576, us32_n577, us32_n578, us32_n579, us32_n580, us32_n581, us32_n582, us32_n583, us32_n584, 
       us32_n585, us32_n586, us32_n587, us32_n588, us32_n589, us32_n590, us32_n591, us32_n592, us32_n593, 
       us32_n594, us32_n595, us32_n596, us32_n597, us32_n598, us32_n599, us32_n600, us32_n601, us32_n602, 
       us32_n603, us32_n604, us32_n605, us32_n606, us32_n607, us32_n608, us32_n609, us32_n610, us32_n611, 
       us32_n612, us32_n613, us32_n614, us32_n615, us32_n616, us32_n617, us32_n618, us32_n619, us32_n620, 
       us32_n621, us32_n622, us32_n623, us32_n624, us32_n625, us32_n626, us32_n627, us32_n628, us32_n629, 
       us32_n630, us32_n631, us32_n632, us32_n633, us32_n634, us32_n635, us32_n636, us32_n637, us32_n638, 
       us32_n639, us32_n640, us32_n641, us32_n642, us32_n643, us32_n644, us32_n645, us32_n646, us32_n647, 
       us32_n648, us32_n649, us32_n650, us32_n651, us32_n652, us32_n653, us32_n654, us32_n655, us32_n656, 
       us32_n657, us32_n658, us32_n659, us32_n660, us32_n661, us32_n662, us32_n663, us32_n664, us32_n665, 
       us32_n666, us32_n667, us32_n668, us32_n669, us32_n670, us32_n671, us32_n672, us32_n673, us32_n674, 
       us32_n675, us32_n676, us32_n677, us32_n678, us32_n679, us32_n680, us32_n681, us32_n682, us32_n683, 
       us32_n684, us32_n685, us32_n686, us32_n687, us32_n688, us32_n689, us32_n690, us32_n691, us32_n692, 
       us32_n693, us32_n694, us32_n695, us32_n696, us32_n697, us32_n698, us32_n699, us32_n700, us32_n701, 
       us32_n702, us32_n703, us32_n704, us32_n705, us32_n706, us32_n707, us32_n708, us32_n709, us32_n710, 
       us32_n711, us32_n712, us32_n713, us32_n714, us32_n715, us32_n716, us32_n717, us32_n718, us32_n719, 
       us32_n720, us32_n721, us32_n722, us32_n723, us32_n724, us32_n725, us32_n726, us32_n727, us32_n728, 
       us32_n729, us32_n730, us32_n731, us32_n732, us32_n733, us32_n734, us32_n735, us32_n736, us32_n737, 
       us32_n738, us32_n739, us32_n740, us32_n741, us32_n742, us32_n743, us32_n744, us32_n745, us32_n746, 
       us32_n747, us32_n748, us32_n749, us32_n750, us32_n751, us32_n752, us32_n753, us32_n754, us32_n755, 
       us32_n756, us32_n757, us32_n758, us32_n759, us32_n760, us32_n761, us32_n762, us32_n763, us32_n764, 
       us32_n765, us32_n766, us32_n767, us32_n768, us32_n769, us32_n770, us32_n771, us32_n772, us32_n773, 
       us32_n774, us32_n775, us32_n776, us32_n777, us32_n778, us32_n779, us32_n780, us32_n781, us32_n782, 
       us32_n783, us32_n784, us32_n785, us32_n786, us32_n787, us32_n788, us32_n789, us32_n790, us32_n791, 
       us32_n792, us32_n793, us32_n794, us32_n795, us32_n796, us32_n797, us32_n798, us32_n799, us32_n800, 
       us32_n801, us32_n802, us32_n803, us32_n804, us32_n805, us32_n806, us32_n807, us32_n808, us32_n809, 
       us32_n810, us32_n811, us32_n812, us32_n813, us32_n814, us32_n815, us32_n816, us32_n817, us32_n818, 
       us32_n819, us32_n820, us32_n821, us32_n822, us32_n823, us32_n824, us32_n825, us32_n826, us32_n827, 
       us32_n828, us32_n829, us32_n830, us32_n831, us32_n832, us32_n833, us32_n834, us32_n835, us32_n836, 
       us32_n837, us32_n838, us32_n839, us32_n840, us32_n841, us32_n842, us32_n843, us32_n844, us32_n845, 
       us32_n846, us32_n847, us32_n848, us32_n849, us32_n850, us32_n851, us32_n852, us32_n853, us32_n854, 
       us32_n855, us32_n856, us32_n857, us32_n858, us32_n859, us32_n860, us32_n861, us32_n862, us32_n863, 
       us32_n864, us32_n865, us32_n866, us32_n867, us32_n868, us32_n869, us32_n870, us32_n871, us32_n872, 
       us32_n873, us32_n874, us32_n875,  us32_n876;
  NOR2_X1 u0_u1_U10 (.ZN( u0_u1_n709 ) , .A2( u0_u1_n778 ) , .A1( u0_u1_n802 ) );
  INV_X1 u0_u1_U100 (.A( u0_u1_n819 ) , .ZN( u0_u1_n845 ) );
  INV_X1 u0_u1_U101 (.A( u0_u1_n674 ) , .ZN( u0_u1_n860 ) );
  AOI21_X1 u0_u1_U102 (.A( u0_u1_n672 ) , .B1( u0_u1_n673 ) , .ZN( u0_u1_n674 ) , .B2( u0_u1_n857 ) );
  INV_X1 u0_u1_U103 (.A( u0_u1_n756 ) , .ZN( u0_u1_n870 ) );
  OAI21_X1 u0_u1_U104 (.B1( u0_u1_n755 ) , .ZN( u0_u1_n756 ) , .A( u0_u1_n846 ) , .B2( u0_u1_n869 ) );
  AOI221_X1 u0_u1_U105 (.A( u0_u1_n715 ) , .B2( u0_u1_n716 ) , .ZN( u0_u1_n722 ) , .C1( u0_u1_n834 ) , .B1( u0_u1_n840 ) , .C2( u0_u1_n864 ) );
  OR2_X1 u0_u1_U106 (.A2( u0_u1_n713 ) , .A1( u0_u1_n714 ) , .ZN( u0_u1_n715 ) );
  NAND2_X1 u0_u1_U107 (.A1( u0_u1_n449 ) , .A2( u0_u1_n451 ) , .ZN( u0_u1_n807 ) );
  NOR3_X1 u0_u1_U108 (.ZN( u0_u1_n754 ) , .A2( u0_u1_n854 ) , .A1( u0_u1_n864 ) , .A3( u0_u1_n866 ) );
  NOR2_X1 u0_u1_U109 (.ZN( u0_u1_n753 ) , .A2( u0_u1_n853 ) , .A1( u0_u1_n861 ) );
  NOR2_X1 u0_u1_U11 (.A1( u0_u1_n680 ) , .ZN( u0_u1_n695 ) , .A2( u0_u1_n809 ) );
  INV_X1 u0_u1_U110 (.A( u0_u1_n440 ) , .ZN( u0_u1_n815 ) );
  NAND2_X1 u0_u1_U111 (.A1( u0_u1_n449 ) , .A2( u0_u1_n467 ) , .ZN( u0_u1_n751 ) );
  AOI211_X1 u0_u1_U112 (.B( u0_u1_n809 ) , .A( u0_u1_n810 ) , .ZN( u0_u1_n826 ) , .C1( u0_u1_n843 ) , .C2( u0_u1_n851 ) );
  NOR2_X1 u0_u1_U113 (.ZN( u0_u1_n509 ) , .A1( u0_u1_n814 ) , .A2( u0_u1_n819 ) );
  OAI22_X1 u0_u1_U114 (.B1( u0_u1_n492 ) , .ZN( u0_u1_n493 ) , .A1( u0_u1_n688 ) , .A2( u0_u1_n765 ) , .B2( u0_u1_n819 ) );
  NOR3_X1 u0_u1_U115 (.ZN( u0_u1_n492 ) , .A1( u0_u1_n784 ) , .A2( u0_u1_n851 ) , .A3( u0_u1_n864 ) );
  NOR2_X1 u0_u1_U116 (.ZN( u0_u1_n579 ) , .A2( u0_u1_n701 ) , .A1( u0_u1_n816 ) );
  NOR2_X1 u0_u1_U117 (.ZN( u0_u1_n548 ) , .A2( u0_u1_n782 ) , .A1( u0_u1_n816 ) );
  NOR2_X1 u0_u1_U118 (.ZN( u0_u1_n508 ) , .A2( u0_u1_n730 ) , .A1( u0_u1_n764 ) );
  INV_X1 u0_u1_U119 (.A( u0_u1_n814 ) , .ZN( u0_u1_n855 ) );
  INV_X1 u0_u1_U12 (.A( u0_u1_n609 ) , .ZN( u0_u1_n875 ) );
  NOR2_X1 u0_u1_U120 (.ZN( u0_u1_n534 ) , .A2( u0_u1_n751 ) , .A1( u0_u1_n752 ) );
  NOR2_X1 u0_u1_U121 (.ZN( u0_u1_n603 ) , .A2( u0_u1_n782 ) , .A1( u0_u1_n805 ) );
  NOR2_X1 u0_u1_U122 (.ZN( u0_u1_n530 ) , .A2( u0_u1_n726 ) , .A1( u0_u1_n805 ) );
  INV_X1 u0_u1_U123 (.A( u0_u1_n816 ) , .ZN( u0_u1_n835 ) );
  AOI21_X1 u0_u1_U124 (.B1( u0_u1_n701 ) , .ZN( u0_u1_n702 ) , .A( u0_u1_n734 ) , .B2( u0_u1_n765 ) );
  NOR2_X1 u0_u1_U125 (.ZN( u0_u1_n557 ) , .A1( u0_u1_n752 ) , .A2( u0_u1_n793 ) );
  NOR2_X1 u0_u1_U126 (.ZN( u0_u1_n668 ) , .A1( u0_u1_n730 ) , .A2( u0_u1_n805 ) );
  NOR2_X1 u0_u1_U127 (.ZN( u0_u1_n547 ) , .A1( u0_u1_n751 ) , .A2( u0_u1_n816 ) );
  NOR2_X1 u0_u1_U128 (.ZN( u0_u1_n511 ) , .A1( u0_u1_n731 ) , .A2( u0_u1_n781 ) );
  NOR2_X1 u0_u1_U129 (.A1( u0_u1_n751 ) , .ZN( u0_u1_n769 ) , .A2( u0_u1_n805 ) );
  INV_X1 u0_u1_U13 (.A( u0_u1_n649 ) , .ZN( u0_u1_n871 ) );
  NOR2_X1 u0_u1_U130 (.ZN( u0_u1_n654 ) , .A1( u0_u1_n671 ) , .A2( u0_u1_n816 ) );
  NOR2_X1 u0_u1_U131 (.ZN( u0_u1_n604 ) , .A1( u0_u1_n671 ) , .A2( u0_u1_n805 ) );
  NOR2_X1 u0_u1_U132 (.ZN( u0_u1_n658 ) , .A1( u0_u1_n749 ) , .A2( u0_u1_n782 ) );
  NOR2_X1 u0_u1_U133 (.ZN( u0_u1_n529 ) , .A1( u0_u1_n671 ) , .A2( u0_u1_n781 ) );
  INV_X1 u0_u1_U134 (.A( u0_u1_n701 ) , .ZN( u0_u1_n854 ) );
  NOR2_X1 u0_u1_U135 (.ZN( u0_u1_n611 ) , .A2( u0_u1_n726 ) , .A1( u0_u1_n819 ) );
  AOI21_X1 u0_u1_U136 (.ZN( u0_u1_n571 ) , .B1( u0_u1_n752 ) , .B2( u0_u1_n764 ) , .A( u0_u1_n782 ) );
  AOI21_X1 u0_u1_U137 (.ZN( u0_u1_n500 ) , .A( u0_u1_n726 ) , .B2( u0_u1_n764 ) , .B1( u0_u1_n816 ) );
  NOR2_X1 u0_u1_U138 (.ZN( u0_u1_n685 ) , .A2( u0_u1_n701 ) , .A1( u0_u1_n805 ) );
  NOR2_X1 u0_u1_U139 (.ZN( u0_u1_n713 ) , .A1( u0_u1_n764 ) , .A2( u0_u1_n765 ) );
  NOR4_X1 u0_u1_U14 (.ZN( u0_u1_n458 ) , .A2( u0_u1_n519 ) , .A1( u0_u1_n545 ) , .A3( u0_u1_n581 ) , .A4( u0_u1_n617 ) );
  INV_X1 u0_u1_U140 (.A( u0_u1_n805 ) , .ZN( u0_u1_n844 ) );
  AOI21_X1 u0_u1_U141 (.ZN( u0_u1_n517 ) , .A( u0_u1_n731 ) , .B1( u0_u1_n752 ) , .B2( u0_u1_n805 ) );
  AOI21_X1 u0_u1_U142 (.B1( u0_u1_n627 ) , .ZN( u0_u1_n629 ) , .A( u0_u1_n765 ) , .B2( u0_u1_n816 ) );
  INV_X1 u0_u1_U143 (.A( u0_u1_n792 ) , .ZN( u0_u1_n834 ) );
  NOR2_X1 u0_u1_U144 (.ZN( u0_u1_n616 ) , .A1( u0_u1_n764 ) , .A2( u0_u1_n814 ) );
  NOR2_X1 u0_u1_U145 (.ZN( u0_u1_n561 ) , .A2( u0_u1_n793 ) , .A1( u0_u1_n805 ) );
  NAND2_X1 u0_u1_U146 (.A1( u0_u1_n701 ) , .A2( u0_u1_n731 ) , .ZN( u0_u1_n784 ) );
  INV_X1 u0_u1_U147 (.A( u0_u1_n749 ) , .ZN( u0_u1_n836 ) );
  INV_X1 u0_u1_U148 (.A( u0_u1_n752 ) , .ZN( u0_u1_n843 ) );
  NOR2_X1 u0_u1_U149 (.ZN( u0_u1_n570 ) , .A1( u0_u1_n731 ) , .A2( u0_u1_n764 ) );
  NOR4_X1 u0_u1_U15 (.ZN( u0_u1_n487 ) , .A2( u0_u1_n535 ) , .A1( u0_u1_n560 ) , .A3( u0_u1_n633 ) , .A4( u0_u1_n720 ) );
  INV_X1 u0_u1_U150 (.A( u0_u1_n730 ) , .ZN( u0_u1_n853 ) );
  AOI21_X1 u0_u1_U151 (.ZN( u0_u1_n566 ) , .B1( u0_u1_n726 ) , .A( u0_u1_n781 ) , .B2( u0_u1_n793 ) );
  AOI21_X1 u0_u1_U152 (.B1( u0_u1_n688 ) , .ZN( u0_u1_n689 ) , .A( u0_u1_n730 ) , .B2( u0_u1_n763 ) );
  INV_X1 u0_u1_U153 (.A( u0_u1_n731 ) , .ZN( u0_u1_n869 ) );
  AOI211_X1 u0_u1_U154 (.C2( u0_u1_n440 ) , .B( u0_u1_n625 ) , .A( u0_u1_n626 ) , .ZN( u0_u1_n637 ) , .C1( u0_u1_n864 ) );
  NOR4_X1 u0_u1_U155 (.A4( u0_u1_n631 ) , .A3( u0_u1_n632 ) , .A2( u0_u1_n633 ) , .A1( u0_u1_n634 ) , .ZN( u0_u1_n635 ) );
  NOR4_X1 u0_u1_U156 (.A4( u0_u1_n628 ) , .A3( u0_u1_n629 ) , .A2( u0_u1_n630 ) , .ZN( u0_u1_n636 ) , .A1( u0_u1_n666 ) );
  AOI21_X1 u0_u1_U157 (.ZN( u0_u1_n542 ) , .A( u0_u1_n765 ) , .B2( u0_u1_n781 ) , .B1( u0_u1_n819 ) );
  OAI21_X1 u0_u1_U158 (.A( u0_u1_n700 ) , .ZN( u0_u1_n704 ) , .B2( u0_u1_n752 ) , .B1( u0_u1_n806 ) );
  OAI21_X1 u0_u1_U159 (.ZN( u0_u1_n700 ) , .B2( u0_u1_n835 ) , .B1( u0_u1_n839 ) , .A( u0_u1_n861 ) );
  NOR4_X1 u0_u1_U16 (.A4( u0_u1_n447 ) , .A3( u0_u1_n448 ) , .A2( u0_u1_n518 ) , .A1( u0_u1_n543 ) , .ZN( u0_u1_n708 ) );
  INV_X1 u0_u1_U160 (.A( u0_u1_n765 ) , .ZN( u0_u1_n867 ) );
  NOR2_X1 u0_u1_U161 (.ZN( u0_u1_n528 ) , .A1( u0_u1_n726 ) , .A2( u0_u1_n752 ) );
  AOI21_X1 u0_u1_U162 (.ZN( u0_u1_n445 ) , .B1( u0_u1_n791 ) , .B2( u0_u1_n793 ) , .A( u0_u1_n816 ) );
  NAND4_X1 u0_u1_U163 (.A4( u0_u1_n495 ) , .A3( u0_u1_n496 ) , .A1( u0_u1_n497 ) , .ZN( u0_u1_n804 ) , .A2( u0_u1_n868 ) );
  AOI221_X1 u0_u1_U164 (.B2( u0_u1_n440 ) , .A( u0_u1_n491 ) , .ZN( u0_u1_n496 ) , .C2( u0_u1_n842 ) , .C1( u0_u1_n852 ) , .B1( u0_u1_n861 ) );
  NOR4_X1 u0_u1_U165 (.A3( u0_u1_n439 ) , .A2( u0_u1_n493 ) , .A1( u0_u1_n494 ) , .ZN( u0_u1_n495 ) , .A4( u0_u1_n614 ) );
  INV_X1 u0_u1_U166 (.A( u0_u1_n780 ) , .ZN( u0_u1_n868 ) );
  AOI21_X1 u0_u1_U167 (.ZN( u0_u1_n499 ) , .A( u0_u1_n781 ) , .B2( u0_u1_n793 ) , .B1( u0_u1_n806 ) );
  INV_X1 u0_u1_U168 (.A( u0_u1_n782 ) , .ZN( u0_u1_n851 ) );
  NAND2_X1 u0_u1_U169 (.ZN( u0_u1_n716 ) , .A1( u0_u1_n730 ) , .A2( u0_u1_n782 ) );
  OR3_X1 u0_u1_U17 (.ZN( u0_u1_n448 ) , .A1( u0_u1_n530 ) , .A3( u0_u1_n579 ) , .A2( u0_u1_n876 ) );
  BUF_X2 u0_u1_U170 (.Z( u0_u1_n41 ) , .A( u0_u1_n699 ) );
  OR4_X1 u0_u1_U171 (.A4( u0_u1_n582 ) , .A3( u0_u1_n583 ) , .A2( u0_u1_n584 ) , .A1( u0_u1_n585 ) , .ZN( u0_u1_n586 ) );
  INV_X1 u0_u1_U172 (.A( u0_u1_n726 ) , .ZN( u0_u1_n857 ) );
  OAI222_X1 u0_u1_U173 (.B2( u0_u1_n710 ) , .ZN( u0_u1_n711 ) , .C2( u0_u1_n726 ) , .B1( u0_u1_n749 ) , .A1( u0_u1_n808 ) , .C1( u0_u1_n816 ) , .A2( u0_u1_n817 ) );
  AOI221_X1 u0_u1_U174 (.A( u0_u1_n766 ) , .ZN( u0_u1_n776 ) , .C2( u0_u1_n812 ) , .B2( u0_u1_n837 ) , .C1( u0_u1_n856 ) , .B1( u0_u1_n867 ) );
  INV_X1 u0_u1_U175 (.A( u0_u1_n763 ) , .ZN( u0_u1_n837 ) );
  OAI221_X1 u0_u1_U176 (.A( u0_u1_n729 ) , .C2( u0_u1_n730 ) , .B2( u0_u1_n731 ) , .B1( u0_u1_n732 ) , .ZN( u0_u1_n739 ) , .C1( u0_u1_n819 ) );
  OAI221_X1 u0_u1_U177 (.C2( u0_u1_n441 ) , .A( u0_u1_n785 ) , .B2( u0_u1_n787 ) , .B1( u0_u1_n788 ) , .ZN( u0_u1_n798 ) , .C1( u0_u1_n815 ) );
  AOI22_X1 u0_u1_U178 (.A2( u0_u1_n784 ) , .ZN( u0_u1_n785 ) , .B2( u0_u1_n833 ) , .A1( u0_u1_n836 ) , .B1( u0_u1_n864 ) );
  OAI221_X1 u0_u1_U179 (.C2( u0_u1_n441 ) , .A( u0_u1_n698 ) , .ZN( u0_u1_n705 ) , .C1( u0_u1_n787 ) , .B1( u0_u1_n788 ) , .B2( u0_u1_n808 ) );
  OR4_X1 u0_u1_U18 (.A4( u0_u1_n444 ) , .A2( u0_u1_n445 ) , .A1( u0_u1_n446 ) , .ZN( u0_u1_n447 ) , .A3( u0_u1_n555 ) );
  AOI22_X1 u0_u1_U180 (.ZN( u0_u1_n698 ) , .A1( u0_u1_n832 ) , .B2( u0_u1_n844 ) , .A2( u0_u1_n866 ) , .B1( u0_u1_n869 ) );
  OAI222_X1 u0_u1_U181 (.B1( u0_u1_n41 ) , .ZN( u0_u1_n619 ) , .C1( u0_u1_n726 ) , .C2( u0_u1_n749 ) , .B2( u0_u1_n788 ) , .A2( u0_u1_n794 ) , .A1( u0_u1_n818 ) );
  NAND2_X1 u0_u1_U182 (.A2( u0_u1_n450 ) , .A1( u0_u1_n466 ) , .ZN( u0_u1_n817 ) );
  NAND2_X1 u0_u1_U183 (.A2( u0_u1_n456 ) , .A1( u0_u1_n474 ) , .ZN( u0_u1_n781 ) );
  NAND2_X1 u0_u1_U184 (.A2( u0_u1_n450 ) , .A1( u0_u1_n454 ) , .ZN( u0_u1_n731 ) );
  NAND2_X1 u0_u1_U185 (.A1( u0_u1_n455 ) , .A2( u0_u1_n474 ) , .ZN( u0_u1_n787 ) );
  NAND2_X1 u0_u1_U186 (.A1( u0_u1_n455 ) , .A2( u0_u1_n463 ) , .ZN( u0_u1_n746 ) );
  NAND2_X1 u0_u1_U187 (.A1( u0_u1_n453 ) , .A2( u0_u1_n473 ) , .ZN( u0_u1_n818 ) );
  NAND2_X1 u0_u1_U188 (.A2( u0_u1_n455 ) , .A1( u0_u1_n457 ) , .ZN( u0_u1_n808 ) );
  NOR2_X1 u0_u1_U189 (.ZN( u0_u1_n467 ) , .A2( u0_u1_n848 ) , .A1( u0_u1_n849 ) );
  INV_X1 u0_u1_U19 (.A( u0_u1_n615 ) , .ZN( u0_u1_n876 ) );
  NAND2_X1 u0_u1_U190 (.A1( u0_u1_n449 ) , .A2( u0_u1_n450 ) , .ZN( u0_u1_n788 ) );
  NAND2_X1 u0_u1_U191 (.A2( u0_u1_n463 ) , .A1( u0_u1_n464 ) , .ZN( u0_u1_n749 ) );
  NAND2_X1 u0_u1_U192 (.A1( u0_u1_n464 ) , .A2( u0_u1_n474 ) , .ZN( u0_u1_n790 ) );
  NAND2_X1 u0_u1_U193 (.A1( u0_u1_n453 ) , .A2( u0_u1_n464 ) , .ZN( u0_u1_n792 ) );
  AND2_X1 u0_u1_U194 (.ZN( u0_u1_n440 ) , .A1( u0_u1_n456 ) , .A2( u0_u1_n463 ) );
  NOR2_X1 u0_u1_U195 (.A2( u0_n268 ) , .ZN( u0_u1_n462 ) , .A1( u0_u1_n850 ) );
  AOI222_X1 u0_u1_U196 (.B2( u0_u1_n640 ) , .ZN( u0_u1_n646 ) , .B1( u0_u1_n842 ) , .A1( u0_u1_n843 ) , .C2( u0_u1_n847 ) , .C1( u0_u1_n864 ) , .A2( u0_u1_n866 ) );
  NOR4_X1 u0_u1_U197 (.A4( u0_u1_n641 ) , .A3( u0_u1_n642 ) , .A2( u0_u1_n643 ) , .A1( u0_u1_n644 ) , .ZN( u0_u1_n645 ) );
  NOR4_X1 u0_u1_U198 (.A4( u0_u1_n500 ) , .A3( u0_u1_n501 ) , .A2( u0_u1_n502 ) , .ZN( u0_u1_n503 ) , .A1( u0_u1_n529 ) );
  AOI221_X1 u0_u1_U199 (.A( u0_u1_n499 ) , .ZN( u0_u1_n504 ) , .B2( u0_u1_n844 ) , .C1( u0_u1_n847 ) , .C2( u0_u1_n861 ) , .B1( u0_u1_n863 ) );
  NOR4_X1 u0_u1_U20 (.ZN( u0_u1_n622 ) , .A1( u0_u1_n658 ) , .A3( u0_u1_n668 ) , .A4( u0_u1_n684 ) , .A2( u0_u1_n768 ) );
  AOI221_X1 u0_u1_U200 (.A( u0_u1_n783 ) , .ZN( u0_u1_n800 ) , .C2( u0_u1_n838 ) , .B2( u0_u1_n839 ) , .B1( u0_u1_n866 ) , .C1( u0_u1_n867 ) );
  NOR4_X1 u0_u1_U201 (.A4( u0_u1_n795 ) , .A3( u0_u1_n796 ) , .A2( u0_u1_n797 ) , .A1( u0_u1_n798 ) , .ZN( u0_u1_n799 ) );
  NAND4_X1 u0_u1_U202 (.ZN( u0_subword_23 ) , .A4( u0_u1_n824 ) , .A3( u0_u1_n825 ) , .A2( u0_u1_n826 ) , .A1( u0_u1_n827 ) );
  NOR4_X1 u0_u1_U203 (.A4( u0_u1_n820 ) , .A3( u0_u1_n821 ) , .A2( u0_u1_n822 ) , .A1( u0_u1_n823 ) , .ZN( u0_u1_n824 ) );
  NOR4_X1 u0_u1_U204 (.A4( u0_u1_n736 ) , .A3( u0_u1_n737 ) , .A2( u0_u1_n738 ) , .A1( u0_u1_n739 ) , .ZN( u0_u1_n740 ) );
  NOR4_X1 u0_u1_U205 (.A3( u0_u1_n757 ) , .A2( u0_u1_n758 ) , .A1( u0_u1_n759 ) , .ZN( u0_u1_n760 ) , .A4( u0_u1_n870 ) );
  AOI211_X1 u0_u1_U206 (.B( u0_u1_n747 ) , .A( u0_u1_n748 ) , .ZN( u0_u1_n761 ) , .C1( u0_u1_n834 ) , .C2( u0_u1_n854 ) );
  NOR4_X1 u0_u1_U207 (.A4( u0_u1_n702 ) , .A3( u0_u1_n703 ) , .A2( u0_u1_n704 ) , .A1( u0_u1_n705 ) , .ZN( u0_u1_n706 ) );
  AOI211_X1 u0_u1_U208 (.B( u0_u1_n696 ) , .A( u0_u1_n697 ) , .ZN( u0_u1_n707 ) , .C2( u0_u1_n833 ) , .C1( u0_u1_n852 ) );
  NAND4_X1 u0_u1_U209 (.ZN( u0_subword_17 ) , .A4( u0_u1_n597 ) , .A3( u0_u1_n598 ) , .A2( u0_u1_n599 ) , .A1( u0_u1_n600 ) );
  NOR4_X1 u0_u1_U21 (.A4( u0_u1_n611 ) , .A3( u0_u1_n612 ) , .A2( u0_u1_n613 ) , .A1( u0_u1_n614 ) , .ZN( u0_u1_n621 ) );
  NOR4_X1 u0_u1_U210 (.A4( u0_u1_n593 ) , .A3( u0_u1_n594 ) , .A2( u0_u1_n595 ) , .A1( u0_u1_n596 ) , .ZN( u0_u1_n597 ) );
  AOI211_X1 u0_u1_U211 (.B( u0_u1_n591 ) , .A( u0_u1_n592 ) , .ZN( u0_u1_n598 ) , .C2( u0_u1_n813 ) , .C1( u0_u1_n835 ) );
  NAND2_X1 u0_u1_U212 (.A2( u0_u1_n443 ) , .A1( u0_u1_n454 ) , .ZN( u0_u1_n793 ) );
  AOI21_X1 u0_u1_U213 (.ZN( u0_u1_n642 ) , .B2( u0_u1_n749 ) , .A( u0_u1_n794 ) , .B1( u0_u1_n805 ) );
  AOI21_X1 u0_u1_U214 (.ZN( u0_u1_n516 ) , .A( u0_u1_n781 ) , .B2( u0_u1_n794 ) , .B1( u0_u1_n814 ) );
  INV_X1 u0_u1_U215 (.A( u0_u1_n794 ) , .ZN( u0_u1_n852 ) );
  NOR2_X1 u0_u1_U216 (.ZN( u0_u1_n559 ) , .A1( u0_u1_n794 ) , .A2( u0_u1_n816 ) );
  NOR2_X1 u0_u1_U217 (.ZN( u0_u1_n585 ) , .A1( u0_u1_n794 ) , .A2( u0_u1_n819 ) );
  NAND2_X2 u0_u1_U218 (.A1( u0_u1_n453 ) , .A2( u0_u1_n455 ) , .ZN( u0_u1_n764 ) );
  NAND2_X2 u0_u1_U219 (.A1( u0_u1_n453 ) , .A2( u0_u1_n456 ) , .ZN( u0_u1_n816 ) );
  NOR4_X1 u0_u1_U22 (.ZN( u0_u1_n563 ) , .A1( u0_u1_n655 ) , .A3( u0_u1_n663 ) , .A4( u0_u1_n687 ) , .A2( u0_u1_n770 ) );
  NOR2_X1 u0_u1_U220 (.ZN( u0_u1_n453 ) , .A1( u0_u1_n830 ) , .A2( u0_u1_n831 ) );
  NAND2_X1 u0_u1_U221 (.A1( u0_u1_n454 ) , .A2( u0_u1_n467 ) , .ZN( u0_u1_n671 ) );
  NAND2_X1 u0_u1_U222 (.A1( u0_u1_n443 ) , .A2( u0_u1_n462 ) , .ZN( u0_u1_n701 ) );
  NOR2_X1 u0_u1_U223 (.ZN( u0_u1_n455 ) , .A1( u0_u1_n828 ) , .A2( u0_u1_n829 ) );
  AOI211_X1 u0_u1_U224 (.B( u0_u1_n727 ) , .A( u0_u1_n728 ) , .ZN( u0_u1_n741 ) , .C1( u0_u1_n844 ) , .C2( u0_u1_n856 ) );
  NOR2_X1 u0_u1_U225 (.A2( u0_u1_n710 ) , .A1( u0_u1_n764 ) , .ZN( u0_u1_n796 ) );
  NOR2_X1 u0_u1_U226 (.ZN( u0_u1_n519 ) , .A1( u0_u1_n710 ) , .A2( u0_u1_n805 ) );
  NOR2_X1 u0_u1_U227 (.ZN( u0_u1_n684 ) , .A2( u0_u1_n710 ) , .A1( u0_u1_n819 ) );
  NOR2_X1 u0_u1_U228 (.A2( u0_u1_n710 ) , .A1( u0_u1_n752 ) , .ZN( u0_u1_n773 ) );
  NOR2_X1 u0_u1_U229 (.ZN( u0_u1_n522 ) , .A2( u0_u1_n710 ) , .A1( u0_u1_n816 ) );
  NOR4_X1 u0_u1_U23 (.ZN( u0_u1_n477 ) , .A1( u0_u1_n533 ) , .A3( u0_u1_n570 ) , .A4( u0_u1_n602 ) , .A2( u0_u1_n644 ) );
  NOR2_X1 u0_u1_U230 (.ZN( u0_u1_n531 ) , .A1( u0_u1_n710 ) , .A2( u0_u1_n781 ) );
  INV_X1 u0_u1_U231 (.A( u0_u1_n682 ) , .ZN( u0_u1_n841 ) );
  AOI21_X1 u0_u1_U232 (.ZN( u0_u1_n643 ) , .B1( u0_u1_n682 ) , .A( u0_u1_n793 ) , .B2( u0_u1_n819 ) );
  OAI22_X1 u0_u1_U233 (.B2( u0_u1_n781 ) , .B1( u0_u1_n782 ) , .ZN( u0_u1_n783 ) , .A2( u0_u1_n816 ) , .A1( u0_u1_n817 ) );
  AOI21_X1 u0_u1_U234 (.ZN( u0_u1_n591 ) , .B2( u0_u1_n701 ) , .B1( u0_u1_n817 ) , .A( u0_u1_n819 ) );
  INV_X1 u0_u1_U235 (.A( u0_u1_n817 ) , .ZN( u0_u1_n856 ) );
  NOR2_X1 u0_u1_U236 (.ZN( u0_u1_n669 ) , .A1( u0_u1_n752 ) , .A2( u0_u1_n817 ) );
  AOI21_X1 u0_u1_U237 (.ZN( u0_u1_n541 ) , .B2( u0_u1_n814 ) , .A( u0_u1_n816 ) , .B1( u0_u1_n817 ) );
  AOI21_X1 u0_u1_U238 (.ZN( u0_u1_n452 ) , .B2( u0_u1_n794 ) , .A( u0_u1_n805 ) , .B1( u0_u1_n817 ) );
  NOR2_X1 u0_u1_U239 (.ZN( u0_u1_n472 ) , .A2( u0_u1_n781 ) , .A1( u0_u1_n817 ) );
  NOR4_X1 u0_u1_U24 (.ZN( u0_u1_n483 ) , .A3( u0_u1_n534 ) , .A4( u0_u1_n547 ) , .A2( u0_u1_n569 ) , .A1( u0_u1_n719 ) );
  OAI222_X1 u0_u1_U240 (.A2( u0_u1_n671 ) , .ZN( u0_u1_n676 ) , .B1( u0_u1_n749 ) , .B2( u0_u1_n786 ) , .C2( u0_u1_n790 ) , .C1( u0_u1_n817 ) , .A1( u0_u1_n819 ) );
  NOR2_X1 u0_u1_U241 (.ZN( u0_u1_n632 ) , .A1( u0_u1_n749 ) , .A2( u0_u1_n817 ) );
  NAND2_X1 u0_u1_U242 (.A1( u0_u1_n443 ) , .A2( u0_u1_n466 ) , .ZN( u0_u1_n710 ) );
  NAND2_X1 u0_u1_U243 (.A2( u0_u1_n463 ) , .A1( u0_u1_n473 ) , .ZN( u0_u1_n699 ) );
  INV_X1 u0_u1_U244 (.ZN( u0_u1_n438 ) , .A( u0_u1_n788 ) );
  INV_X1 u0_u1_U245 (.ZN( u0_u1_n828 ) , .A( w3_8 ) );
  NOR2_X1 u0_u1_U246 (.ZN( u0_u1_n456 ) , .A1( u0_u1_n829 ) , .A2( w3_8 ) );
  NOR2_X1 u0_u1_U247 (.A2( u0_n270 ) , .ZN( u0_u1_n454 ) , .A1( u0_u1_n859 ) );
  OAI21_X1 u0_u1_U248 (.A( u0_u1_n789 ) , .B2( u0_u1_n790 ) , .B1( u0_u1_n791 ) , .ZN( u0_u1_n797 ) );
  AOI21_X1 u0_u1_U249 (.ZN( u0_u1_n641 ) , .B2( u0_u1_n751 ) , .A( u0_u1_n790 ) , .B1( u0_u1_n814 ) );
  INV_X1 u0_u1_U25 (.A( u0_u1_n751 ) , .ZN( u0_u1_n864 ) );
  AOI21_X1 u0_u1_U250 (.A( u0_u1_n735 ) , .ZN( u0_u1_n736 ) , .B2( u0_u1_n782 ) , .B1( u0_u1_n794 ) );
  AOI21_X1 u0_u1_U251 (.B2( u0_u1_n765 ) , .ZN( u0_u1_n766 ) , .A( u0_u1_n790 ) , .B1( u0_u1_n794 ) );
  AOI21_X1 u0_u1_U252 (.ZN( u0_u1_n444 ) , .A( u0_u1_n701 ) , .B1( u0_u1_n735 ) , .B2( u0_u1_n752 ) );
  NOR2_X1 u0_u1_U253 (.ZN( u0_u1_n520 ) , .A1( u0_u1_n710 ) , .A2( u0_u1_n790 ) );
  NOR2_X1 u0_u1_U254 (.ZN( u0_u1_n536 ) , .A1( u0_u1_n726 ) , .A2( u0_u1_n790 ) );
  NOR2_X1 u0_u1_U255 (.ZN( u0_u1_n644 ) , .A2( u0_u1_n790 ) , .A1( u0_u1_n793 ) );
  NOR2_X1 u0_u1_U256 (.ZN( u0_u1_n583 ) , .A1( u0_u1_n671 ) , .A2( u0_u1_n790 ) );
  INV_X1 u0_u1_U257 (.A( u0_u1_n790 ) , .ZN( u0_u1_n846 ) );
  AOI222_X1 u0_u1_U258 (.ZN( u0_u1_n527 ) , .A1( u0_u1_n836 ) , .B2( u0_u1_n838 ) , .C1( u0_u1_n845 ) , .C2( u0_u1_n851 ) , .A2( u0_u1_n853 ) , .B1( u0_u1_n867 ) );
  NOR3_X1 u0_u1_U259 (.A2( u0_u1_n440 ) , .ZN( u0_u1_n442 ) , .A3( u0_u1_n838 ) , .A1( u0_u1_n847 ) );
  NOR4_X1 u0_u1_U26 (.A1( u0_u1_n533 ) , .ZN( u0_u1_n538 ) , .A2( u0_u1_n656 ) , .A4( u0_u1_n670 ) , .A3( u0_u1_n767 ) );
  NAND2_X1 u0_u1_U260 (.ZN( u0_u1_n615 ) , .A2( u0_u1_n838 ) , .A1( u0_u1_n874 ) );
  AND2_X1 u0_u1_U261 (.ZN( u0_u1_n627 ) , .A1( u0_u1_n732 ) , .A2( u0_u1_n815 ) );
  NAND2_X1 u0_u1_U262 (.A2( u0_u1_n456 ) , .A1( u0_u1_n457 ) , .ZN( u0_u1_n732 ) );
  NOR2_X1 u0_u1_U263 (.A2( u0_u1_n41 ) , .ZN( u0_u1_n439 ) , .A1( u0_u1_n793 ) );
  AOI21_X1 u0_u1_U264 (.ZN( u0_u1_n593 ) , .B2( u0_u1_n765 ) , .A( u0_u1_n787 ) , .B1( u0_u1_n814 ) );
  AND2_X1 u0_u1_U265 (.ZN( u0_u1_n734 ) , .A1( u0_u1_n781 ) , .A2( u0_u1_n787 ) );
  NAND4_X1 u0_u1_U266 (.A4( u0_u1_n550 ) , .A3( u0_u1_n551 ) , .A2( u0_u1_n552 ) , .A1( u0_u1_n553 ) , .ZN( u0_u1_n747 ) );
  NOR2_X1 u0_u1_U267 (.ZN( u0_u1_n666 ) , .A1( u0_u1_n787 ) , .A2( u0_u1_n793 ) );
  NOR2_X1 u0_u1_U268 (.ZN( u0_u1_n665 ) , .A1( u0_u1_n731 ) , .A2( u0_u1_n787 ) );
  NOR2_X1 u0_u1_U269 (.ZN( u0_u1_n510 ) , .A2( u0_u1_n782 ) , .A1( u0_u1_n787 ) );
  NOR4_X1 u0_u1_U27 (.A4( u0_u1_n543 ) , .A3( u0_u1_n544 ) , .A2( u0_u1_n545 ) , .ZN( u0_u1_n552 ) , .A1( u0_u1_n690 ) );
  NOR2_X1 u0_u1_U270 (.ZN( u0_u1_n630 ) , .A2( u0_u1_n671 ) , .A1( u0_u1_n787 ) );
  NOR2_X1 u0_u1_U271 (.ZN( u0_u1_n617 ) , .A1( u0_u1_n787 ) , .A2( u0_u1_n817 ) );
  INV_X1 u0_u1_U272 (.A( u0_u1_n787 ) , .ZN( u0_u1_n847 ) );
  NOR2_X1 u0_u1_U273 (.ZN( u0_u1_n545 ) , .A2( u0_u1_n710 ) , .A1( u0_u1_n787 ) );
  NOR2_X1 u0_u1_U274 (.ZN( u0_u1_n546 ) , .A2( u0_u1_n787 ) , .A1( u0_u1_n794 ) );
  NAND2_X1 u0_u1_U275 (.A2( u0_u1_n473 ) , .A1( u0_u1_n474 ) , .ZN( u0_u1_n819 ) );
  AOI222_X1 u0_u1_U276 (.C2( u0_u1_n811 ) , .B2( u0_u1_n812 ) , .A2( u0_u1_n813 ) , .ZN( u0_u1_n825 ) , .C1( u0_u1_n834 ) , .A1( u0_u1_n840 ) , .B1( u0_u1_n854 ) );
  AOI22_X1 u0_u1_U277 (.ZN( u0_u1_n729 ) , .B1( u0_u1_n834 ) , .A2( u0_u1_n839 ) , .A1( u0_u1_n864 ) , .B2( u0_u1_n867 ) );
  AOI222_X1 u0_u1_U278 (.ZN( u0_u1_n471 ) , .B1( u0_u1_n834 ) , .A1( u0_u1_n840 ) , .C1( u0_u1_n843 ) , .C2( u0_u1_n852 ) , .A2( u0_u1_n856 ) , .B2( u0_u1_n866 ) );
  NOR2_X1 u0_u1_U279 (.ZN( u0_u1_n688 ) , .A1( u0_u1_n833 ) , .A2( u0_u1_n834 ) );
  NOR2_X1 u0_u1_U28 (.ZN( u0_u1_n544 ) , .A1( u0_u1_n764 ) , .A2( u0_u1_n793 ) );
  NOR2_X1 u0_u1_U280 (.ZN( u0_u1_n735 ) , .A2( u0_u1_n834 ) , .A1( u0_u1_n846 ) );
  NAND4_X1 u0_u1_U281 (.A4( u0_u1_n537 ) , .A3( u0_u1_n538 ) , .A2( u0_u1_n539 ) , .A1( u0_u1_n540 ) , .ZN( u0_u1_n624 ) );
  NAND2_X2 u0_u1_U282 (.A1( u0_u1_n451 ) , .A2( u0_u1_n462 ) , .ZN( u0_u1_n794 ) );
  NAND2_X1 u0_u1_U283 (.A2( u0_u1_n466 ) , .A1( u0_u1_n467 ) , .ZN( u0_u1_n814 ) );
  NOR2_X1 u0_u1_U284 (.ZN( u0_u1_n631 ) , .A2( u0_u1_n730 ) , .A1( u0_u1_n787 ) );
  NAND2_X2 u0_u1_U285 (.A2( u0_u1_n450 ) , .A1( u0_u1_n462 ) , .ZN( u0_u1_n730 ) );
  NOR2_X1 u0_u1_U286 (.A2( u0_n274 ) , .ZN( u0_u1_n451 ) , .A1( u0_u1_n849 ) );
  NOR2_X1 u0_u1_U287 (.A1( u0_n272 ) , .A2( u0_n274 ) , .ZN( u0_u1_n443 ) );
  OAI22_X1 u0_u1_U288 (.ZN( u0_u1_n697 ) , .A2( u0_u1_n732 ) , .A1( u0_u1_n782 ) , .B1( u0_u1_n793 ) , .B2( u0_u1_n819 ) );
  AOI21_X1 u0_u1_U289 (.ZN( u0_u1_n512 ) , .B2( u0_u1_n671 ) , .A( u0_u1_n732 ) , .B1( u0_u1_n817 ) );
  NAND4_X1 u0_u1_U29 (.A4( u0_u1_n605 ) , .A3( u0_u1_n606 ) , .A2( u0_u1_n607 ) , .A1( u0_u1_n608 ) , .ZN( u0_u1_n724 ) );
  OAI22_X1 u0_u1_U290 (.ZN( u0_u1_n491 ) , .A1( u0_u1_n726 ) , .B2( u0_u1_n730 ) , .B1( u0_u1_n732 ) , .A2( u0_u1_n781 ) );
  NOR2_X1 u0_u1_U291 (.ZN( u0_u1_n581 ) , .A2( u0_u1_n710 ) , .A1( u0_u1_n732 ) );
  NOR2_X1 u0_u1_U292 (.ZN( u0_u1_n535 ) , .A2( u0_u1_n726 ) , .A1( u0_u1_n732 ) );
  INV_X1 u0_u1_U293 (.A( u0_u1_n732 ) , .ZN( u0_u1_n840 ) );
  AOI211_X1 u0_u1_U294 (.A( u0_u1_n498 ) , .ZN( u0_u1_n505 ) , .B( u0_u1_n804 ) , .C2( u0_u1_n840 ) , .C1( u0_u1_n852 ) );
  OAI21_X1 u0_u1_U295 (.ZN( u0_u1_n789 ) , .A( u0_u1_n840 ) , .B1( u0_u1_n864 ) , .B2( u0_u1_n874 ) );
  AOI222_X1 u0_u1_U296 (.ZN( u0_u1_n662 ) , .A2( u0_u1_n840 ) , .B1( u0_u1_n842 ) , .C2( u0_u1_n846 ) , .A1( u0_u1_n861 ) , .C1( u0_u1_n864 ) , .B2( u0_u1_n871 ) );
  AOI211_X1 u0_u1_U297 (.B( u0_u1_n541 ) , .A( u0_u1_n542 ) , .ZN( u0_u1_n553 ) , .C2( u0_u1_n840 ) , .C1( u0_u1_n852 ) );
  NOR2_X1 u0_u1_U298 (.ZN( u0_u1_n682 ) , .A2( u0_u1_n836 ) , .A1( u0_u1_n840 ) );
  NAND4_X1 u0_u1_U299 (.ZN( u0_subword_16 ) , .A4( u0_u1_n503 ) , .A3( u0_u1_n504 ) , .A2( u0_u1_n505 ) , .A1( u0_u1_n506 ) );
  NAND2_X1 u0_u1_U3 (.A1( u0_u1_n451 ) , .A2( u0_u1_n466 ) , .ZN( u0_u1_n726 ) );
  NOR4_X1 u0_u1_U30 (.A3( u0_u1_n602 ) , .A2( u0_u1_n603 ) , .A1( u0_u1_n604 ) , .ZN( u0_u1_n605 ) , .A4( u0_u1_n657 ) );
  AOI21_X1 u0_u1_U300 (.A( u0_u1_n792 ) , .B2( u0_u1_n793 ) , .B1( u0_u1_n794 ) , .ZN( u0_u1_n795 ) );
  AOI21_X1 u0_u1_U301 (.ZN( u0_u1_n628 ) , .B2( u0_u1_n671 ) , .A( u0_u1_n792 ) , .B1( u0_u1_n793 ) );
  NOR2_X1 u0_u1_U302 (.ZN( u0_u1_n657 ) , .A1( u0_u1_n792 ) , .A2( u0_u1_n817 ) );
  NOR2_X1 u0_u1_U303 (.ZN( u0_u1_n714 ) , .A2( u0_u1_n726 ) , .A1( u0_u1_n792 ) );
  NOR2_X1 u0_u1_U304 (.ZN( u0_u1_n523 ) , .A1( u0_u1_n792 ) , .A2( u0_u1_n814 ) );
  NOR2_X1 u0_u1_U305 (.ZN( u0_u1_n663 ) , .A1( u0_u1_n731 ) , .A2( u0_u1_n792 ) );
  NOR2_X1 u0_u1_U306 (.ZN( u0_u1_n670 ) , .A2( u0_u1_n710 ) , .A1( u0_u1_n792 ) );
  NOR3_X1 u0_u1_U307 (.A3( u0_u1_n743 ) , .A2( u0_u1_n744 ) , .A1( u0_u1_n745 ) , .ZN( u0_u1_n762 ) );
  NAND2_X2 u0_u1_U308 (.A2( u0_u1_n451 ) , .A1( u0_u1_n454 ) , .ZN( u0_u1_n765 ) );
  OAI22_X1 u0_u1_U309 (.ZN( u0_u1_n639 ) , .A1( u0_u1_n701 ) , .B2( u0_u1_n730 ) , .A2( u0_u1_n764 ) , .B1( u0_u1_n818 ) );
  NOR3_X1 u0_u1_U31 (.A1( u0_u1_n601 ) , .ZN( u0_u1_n606 ) , .A3( u0_u1_n665 ) , .A2( u0_u1_n772 ) );
  AOI21_X1 u0_u1_U310 (.ZN( u0_u1_n501 ) , .B1( u0_u1_n682 ) , .A( u0_u1_n814 ) , .B2( u0_u1_n818 ) );
  OAI22_X1 u0_u1_U311 (.A1( u0_u1_n726 ) , .ZN( u0_u1_n728 ) , .B2( u0_u1_n752 ) , .B1( u0_u1_n814 ) , .A2( u0_u1_n818 ) );
  AOI21_X1 u0_u1_U312 (.A( u0_u1_n817 ) , .B2( u0_u1_n818 ) , .B1( u0_u1_n819 ) , .ZN( u0_u1_n820 ) );
  OAI22_X1 u0_u1_U313 (.ZN( u0_u1_n626 ) , .B1( u0_u1_n671 ) , .B2( u0_u1_n749 ) , .A1( u0_u1_n817 ) , .A2( u0_u1_n818 ) );
  NOR2_X1 u0_u1_U314 (.ZN( u0_u1_n601 ) , .A2( u0_u1_n793 ) , .A1( u0_u1_n818 ) );
  NOR2_X1 u0_u1_U315 (.ZN( u0_u1_n533 ) , .A2( u0_u1_n782 ) , .A1( u0_u1_n818 ) );
  NOR2_X1 u0_u1_U316 (.A1( u0_u1_n671 ) , .ZN( u0_u1_n690 ) , .A2( u0_u1_n818 ) );
  NOR2_X1 u0_u1_U317 (.ZN( u0_u1_n521 ) , .A2( u0_u1_n701 ) , .A1( u0_u1_n818 ) );
  NOR2_X1 u0_u1_U318 (.ZN( u0_u1_n560 ) , .A1( u0_u1_n710 ) , .A2( u0_u1_n818 ) );
  NOR2_X1 u0_u1_U319 (.ZN( u0_u1_n687 ) , .A1( u0_u1_n731 ) , .A2( u0_u1_n818 ) );
  NOR3_X1 u0_u1_U32 (.ZN( u0_u1_n551 ) , .A2( u0_u1_n653 ) , .A1( u0_u1_n669 ) , .A3( u0_u1_n773 ) );
  INV_X1 u0_u1_U320 (.A( u0_u1_n818 ) , .ZN( u0_u1_n833 ) );
  BUF_X2 u0_u1_U321 (.Z( u0_u1_n441 ) , .A( u0_u1_n786 ) );
  NAND2_X1 u0_u1_U322 (.A2( u0_u1_n443 ) , .A1( u0_u1_n449 ) , .ZN( u0_u1_n786 ) );
  AOI222_X1 u0_u1_U323 (.ZN( u0_u1_n777 ) , .A1( u0_u1_n832 ) , .C1( u0_u1_n836 ) , .B2( u0_u1_n842 ) , .A2( u0_u1_n851 ) , .B1( u0_u1_n862 ) , .C2( u0_u1_n874 ) );
  INV_X1 u0_u1_U324 (.A( u0_n268 ) , .ZN( u0_u1_n859 ) );
  INV_X1 u0_u1_U325 (.A( u0_n274 ) , .ZN( u0_u1_n848 ) );
  INV_X1 u0_u1_U326 (.A( u0_u1_n786 ) , .ZN( u0_u1_n862 ) );
  OAI22_X1 u0_u1_U327 (.B2( u0_u1_n752 ) , .B1( u0_u1_n753 ) , .A1( u0_u1_n754 ) , .ZN( u0_u1_n758 ) , .A2( u0_u1_n808 ) );
  OAI222_X1 u0_u1_U328 (.ZN( u0_u1_n507 ) , .C2( u0_u1_n627 ) , .B2( u0_u1_n649 ) , .B1( u0_u1_n749 ) , .A2( u0_u1_n750 ) , .C1( u0_u1_n807 ) , .A1( u0_u1_n808 ) );
  AOI21_X1 u0_u1_U329 (.ZN( u0_u1_n691 ) , .B2( u0_u1_n751 ) , .B1( u0_u1_n765 ) , .A( u0_u1_n808 ) );
  NOR4_X1 u0_u1_U33 (.A4( u0_u1_n546 ) , .A3( u0_u1_n547 ) , .A2( u0_u1_n548 ) , .A1( u0_u1_n549 ) , .ZN( u0_u1_n550 ) );
  NAND2_X1 u0_u1_U330 (.A2( u0_u1_n764 ) , .A1( u0_u1_n808 ) , .ZN( u0_u1_n812 ) );
  NOR2_X1 u0_u1_U331 (.ZN( u0_u1_n572 ) , .A1( u0_u1_n730 ) , .A2( u0_u1_n808 ) );
  AOI21_X1 u0_u1_U332 (.ZN( u0_u1_n479 ) , .A( u0_u1_n671 ) , .B1( u0_u1_n752 ) , .B2( u0_u1_n808 ) );
  OAI22_X1 u0_u1_U333 (.ZN( u0_u1_n485 ) , .A1( u0_u1_n710 ) , .B2( u0_u1_n787 ) , .A2( u0_u1_n808 ) , .B1( u0_u1_n814 ) );
  NOR2_X1 u0_u1_U334 (.ZN( u0_u1_n613 ) , .A2( u0_u1_n782 ) , .A1( u0_u1_n808 ) );
  INV_X1 u0_u1_U335 (.A( u0_u1_n808 ) , .ZN( u0_u1_n842 ) );
  NAND2_X1 u0_u1_U336 (.ZN( u0_u1_n673 ) , .A1( u0_u1_n808 ) , .A2( u0_u1_n818 ) );
  NOR2_X1 u0_u1_U337 (.ZN( u0_u1_n464 ) , .A2( w3_8 ) , .A1( w3_9 ) );
  NOR2_X1 u0_u1_U338 (.ZN( u0_u1_n473 ) , .A1( u0_u1_n828 ) , .A2( w3_9 ) );
  INV_X1 u0_u1_U339 (.ZN( u0_u1_n829 ) , .A( w3_9 ) );
  NOR2_X1 u0_u1_U34 (.ZN( u0_u1_n806 ) , .A1( u0_u1_n855 ) , .A2( u0_u1_n862 ) );
  NAND2_X2 u0_u1_U340 (.A1( u0_u1_n457 ) , .A2( u0_u1_n464 ) , .ZN( u0_u1_n752 ) );
  NOR2_X1 u0_u1_U341 (.ZN( u0_u1_n463 ) , .A1( u0_u1_n831 ) , .A2( w3_10 ) );
  INV_X1 u0_u1_U342 (.ZN( u0_u1_n830 ) , .A( w3_10 ) );
  AOI211_X1 u0_u1_U343 (.A( u0_u1_n590 ) , .ZN( u0_u1_n599 ) , .B( u0_u1_n623 ) , .C1( u0_u1_n846 ) , .C2( u0_u1_n856 ) );
  NOR3_X1 u0_u1_U344 (.A3( u0_u1_n623 ) , .A2( u0_u1_n624 ) , .ZN( u0_u1_n638 ) , .A1( u0_u1_n727 ) );
  AOI211_X1 u0_u1_U345 (.B( u0_u1_n479 ) , .A( u0_u1_n480 ) , .ZN( u0_u1_n484 ) , .C2( u0_u1_n835 ) , .C1( u0_u1_n862 ) );
  AOI222_X1 u0_u1_U346 (.ZN( u0_u1_n608 ) , .A1( u0_u1_n832 ) , .C2( u0_u1_n838 ) , .B1( u0_u1_n843 ) , .A2( u0_u1_n857 ) , .B2( u0_u1_n862 ) , .C1( u0_u1_n869 ) );
  AOI21_X1 u0_u1_U347 (.ZN( u0_u1_n595 ) , .B1( u0_u1_n752 ) , .A( u0_u1_n794 ) , .B2( u0_u1_n815 ) );
  AOI21_X1 u0_u1_U348 (.A( u0_u1_n814 ) , .B2( u0_u1_n815 ) , .B1( u0_u1_n816 ) , .ZN( u0_u1_n821 ) );
  AOI21_X1 u0_u1_U349 (.ZN( u0_u1_n651 ) , .B1( u0_u1_n731 ) , .B2( u0_u1_n765 ) , .A( u0_u1_n815 ) );
  NAND4_X1 u0_u1_U35 (.A4( u0_u1_n659 ) , .A3( u0_u1_n660 ) , .A2( u0_u1_n661 ) , .A1( u0_u1_n662 ) , .ZN( u0_u1_n802 ) );
  NOR4_X1 u0_u1_U350 (.A4( u0_u1_n616 ) , .A3( u0_u1_n617 ) , .A2( u0_u1_n618 ) , .A1( u0_u1_n619 ) , .ZN( u0_u1_n620 ) );
  NOR2_X1 u0_u1_U351 (.A1( u0_u1_n671 ) , .ZN( u0_u1_n768 ) , .A2( u0_u1_n815 ) );
  NOR2_X1 u0_u1_U352 (.A2( u0_u1_n815 ) , .A1( u0_u1_n817 ) , .ZN( u0_u1_n823 ) );
  NOR2_X1 u0_u1_U353 (.ZN( u0_u1_n580 ) , .A1( u0_u1_n710 ) , .A2( u0_u1_n815 ) );
  NOR2_X1 u0_u1_U354 (.ZN( u0_u1_n667 ) , .A1( u0_u1_n782 ) , .A2( u0_u1_n815 ) );
  NOR2_X1 u0_u1_U355 (.ZN( u0_u1_n686 ) , .A1( u0_u1_n793 ) , .A2( u0_u1_n815 ) );
  NOR2_X1 u0_u1_U356 (.A1( u0_u1_n701 ) , .ZN( u0_u1_n770 ) , .A2( u0_u1_n815 ) );
  NOR2_X1 u0_u1_U357 (.ZN( u0_u1_n656 ) , .A1( u0_u1_n730 ) , .A2( u0_u1_n815 ) );
  NOR2_X1 u0_u1_U358 (.ZN( u0_u1_n633 ) , .A1( u0_u1_n726 ) , .A2( u0_u1_n815 ) );
  NOR2_X1 u0_u1_U359 (.ZN( u0_u1_n457 ) , .A1( u0_u1_n830 ) , .A2( w3_11 ) );
  NOR3_X1 u0_u1_U36 (.A3( u0_u1_n650 ) , .A2( u0_u1_n651 ) , .A1( u0_u1_n652 ) , .ZN( u0_u1_n661 ) );
  NOR2_X1 u0_u1_U360 (.ZN( u0_u1_n474 ) , .A2( w3_10 ) , .A1( w3_11 ) );
  INV_X1 u0_u1_U361 (.ZN( u0_u1_n831 ) , .A( w3_11 ) );
  INV_X1 u0_u1_U362 (.A( u0_n270 ) , .ZN( u0_u1_n850 ) );
  NOR2_X1 u0_u1_U363 (.A1( u0_n268 ) , .A2( u0_n270 ) , .ZN( u0_u1_n466 ) );
  NOR2_X1 u0_u1_U364 (.ZN( u0_u1_n449 ) , .A2( u0_u1_n850 ) , .A1( u0_u1_n859 ) );
  INV_X1 u0_u1_U365 (.A( u0_n272 ) , .ZN( u0_u1_n849 ) );
  NOR2_X1 u0_u1_U366 (.A2( u0_n272 ) , .ZN( u0_u1_n450 ) , .A1( u0_u1_n848 ) );
  NOR2_X1 u0_u1_U367 (.A2( u0_u1_n438 ) , .ZN( u0_u1_n750 ) , .A1( u0_u1_n862 ) );
  NOR4_X1 u0_u1_U368 (.A4( u0_u1_n778 ) , .A3( u0_u1_n779 ) , .A1( u0_u1_n780 ) , .ZN( u0_u1_n801 ) , .A2( u0_u1_n803 ) );
  NAND4_X1 u0_u1_U369 (.A4( u0_u1_n693 ) , .A3( u0_u1_n694 ) , .A1( u0_u1_n695 ) , .ZN( u0_u1_n778 ) , .A2( u0_u1_n873 ) );
  NOR3_X1 u0_u1_U37 (.A3( u0_u1_n653 ) , .A2( u0_u1_n654 ) , .A1( u0_u1_n655 ) , .ZN( u0_u1_n660 ) );
  INV_X1 u0_u1_U370 (.A( u0_u1_n41 ) , .ZN( u0_u1_n839 ) );
  NOR2_X1 u0_u1_U371 (.A1( u0_u1_n41 ) , .ZN( u0_u1_n772 ) , .A2( u0_u1_n817 ) );
  NAND2_X2 u0_u1_U372 (.A1( u0_u1_n457 ) , .A2( u0_u1_n473 ) , .ZN( u0_u1_n805 ) );
  AOI21_X1 u0_u1_U373 (.B2( u0_u1_n41 ) , .ZN( u0_u1_n573 ) , .B1( u0_u1_n808 ) , .A( u0_u1_n814 ) );
  NOR2_X1 u0_u1_U374 (.A2( u0_u1_n41 ) , .A1( u0_u1_n782 ) , .ZN( u0_u1_n822 ) );
  NOR2_X1 u0_u1_U375 (.A2( u0_u1_n41 ) , .ZN( u0_u1_n634 ) , .A1( u0_u1_n726 ) );
  NOR2_X1 u0_u1_U376 (.A2( u0_u1_n41 ) , .ZN( u0_u1_n568 ) , .A1( u0_u1_n765 ) );
  NOR2_X1 u0_u1_U377 (.A2( u0_u1_n41 ) , .ZN( u0_u1_n664 ) , .A1( u0_u1_n731 ) );
  AOI21_X1 u0_u1_U378 (.B2( u0_u1_n41 ) , .ZN( u0_u1_n480 ) , .A( u0_u1_n751 ) , .B1( u0_u1_n781 ) );
  NOR2_X1 u0_u1_U379 (.A2( u0_u1_n41 ) , .ZN( u0_u1_n718 ) , .A1( u0_u1_n794 ) );
  NOR3_X1 u0_u1_U38 (.A3( u0_u1_n656 ) , .A2( u0_u1_n657 ) , .A1( u0_u1_n658 ) , .ZN( u0_u1_n659 ) );
  NOR2_X1 u0_u1_U380 (.A2( u0_u1_n41 ) , .ZN( u0_u1_n596 ) , .A1( u0_u1_n730 ) );
  NOR2_X1 u0_u1_U381 (.A2( u0_u1_n41 ) , .ZN( u0_u1_n543 ) , .A1( u0_u1_n701 ) );
  NOR2_X1 u0_u1_U382 (.ZN( u0_u1_n582 ) , .A2( u0_u1_n699 ) , .A1( u0_u1_n793 ) );
  NAND4_X1 u0_u1_U383 (.ZN( u0_subword_18 ) , .A4( u0_u1_n645 ) , .A3( u0_u1_n646 ) , .A2( u0_u1_n647 ) , .A1( u0_u1_n648 ) );
  OAI21_X1 u0_u1_U384 (.A( u0_u1_n733 ) , .B1( u0_u1_n734 ) , .ZN( u0_u1_n738 ) , .B2( u0_u1_n807 ) );
  OAI222_X1 u0_u1_U385 (.B2( u0_u1_n749 ) , .B1( u0_u1_n750 ) , .A2( u0_u1_n751 ) , .ZN( u0_u1_n759 ) , .C2( u0_u1_n807 ) , .C1( u0_u1_n816 ) , .A1( u0_u1_n819 ) );
  OAI22_X1 u0_u1_U386 (.B2( u0_u1_n805 ) , .B1( u0_u1_n806 ) , .A2( u0_u1_n807 ) , .A1( u0_u1_n808 ) , .ZN( u0_u1_n810 ) );
  AOI21_X1 u0_u1_U387 (.ZN( u0_u1_n652 ) , .A( u0_u1_n781 ) , .B1( u0_u1_n794 ) , .B2( u0_u1_n807 ) );
  INV_X1 u0_u1_U388 (.A( u0_u1_n807 ) , .ZN( u0_u1_n861 ) );
  NOR2_X1 u0_u1_U389 (.ZN( u0_u1_n737 ) , .A2( u0_u1_n805 ) , .A1( u0_u1_n807 ) );
  OAI21_X1 u0_u1_U39 (.ZN( u0_u1_n733 ) , .A( u0_u1_n835 ) , .B2( u0_u1_n853 ) , .B1( u0_u1_n874 ) );
  NOR2_X1 u0_u1_U390 (.ZN( u0_u1_n486 ) , .A1( u0_u1_n790 ) , .A2( u0_u1_n807 ) );
  NOR2_X1 u0_u1_U391 (.ZN( u0_u1_n569 ) , .A1( u0_u1_n749 ) , .A2( u0_u1_n807 ) );
  AOI21_X1 u0_u1_U392 (.A( u0_u1_n41 ) , .ZN( u0_u1_n554 ) , .B1( u0_u1_n671 ) , .B2( u0_u1_n807 ) );
  NAND2_X1 u0_u1_U393 (.ZN( u0_u1_n755 ) , .A1( u0_u1_n765 ) , .A2( u0_u1_n807 ) );
  NOR2_X1 u0_u1_U394 (.ZN( u0_u1_n717 ) , .A1( u0_u1_n807 ) , .A2( u0_u1_n819 ) );
  NOR2_X1 u0_u1_U395 (.ZN( u0_u1_n558 ) , .A1( u0_u1_n764 ) , .A2( u0_u1_n807 ) );
  NOR2_X1 u0_u1_U396 (.ZN( u0_u1_n672 ) , .A1( u0_u1_n792 ) , .A2( u0_u1_n807 ) );
  NAND4_X1 u0_u1_U397 (.ZN( u0_subword_19 ) , .A4( u0_u1_n706 ) , .A3( u0_u1_n707 ) , .A2( u0_u1_n708 ) , .A1( u0_u1_n709 ) );
  INV_X1 u0_u1_U398 (.A( u0_u1_n708 ) , .ZN( u0_u1_n877 ) );
  OAI22_X1 u0_u1_U399 (.B2( u0_u1_n746 ) , .ZN( u0_u1_n748 ) , .A2( u0_u1_n764 ) , .B1( u0_u1_n782 ) , .A1( u0_u1_n794 ) );
  NAND2_X1 u0_u1_U4 (.A2( u0_u1_n462 ) , .A1( u0_u1_n467 ) , .ZN( u0_u1_n782 ) );
  INV_X1 u0_u1_U40 (.A( u0_u1_n681 ) , .ZN( u0_u1_n873 ) );
  OAI22_X1 u0_u1_U400 (.ZN( u0_u1_n498 ) , .A2( u0_u1_n746 ) , .A1( u0_u1_n782 ) , .B1( u0_u1_n793 ) , .B2( u0_u1_n808 ) );
  NOR2_X1 u0_u1_U401 (.ZN( u0_u1_n518 ) , .A1( u0_u1_n710 ) , .A2( u0_u1_n746 ) );
  OAI22_X1 u0_u1_U402 (.ZN( u0_u1_n712 ) , .A2( u0_u1_n730 ) , .B2( u0_u1_n731 ) , .A1( u0_u1_n746 ) , .B1( u0_u1_n815 ) );
  NOR2_X1 u0_u1_U403 (.A2( u0_u1_n746 ) , .ZN( u0_u1_n771 ) , .A1( u0_u1_n814 ) );
  OAI22_X1 u0_u1_U404 (.B1( u0_u1_n442 ) , .ZN( u0_u1_n446 ) , .A2( u0_u1_n730 ) , .A1( u0_u1_n746 ) , .B2( u0_u1_n751 ) );
  NOR2_X1 u0_u1_U405 (.ZN( u0_u1_n549 ) , .A1( u0_u1_n701 ) , .A2( u0_u1_n746 ) );
  NOR2_X1 u0_u1_U406 (.ZN( u0_u1_n532 ) , .A2( u0_u1_n746 ) , .A1( u0_u1_n794 ) );
  NOR2_X1 u0_u1_U407 (.A2( u0_u1_n746 ) , .ZN( u0_u1_n757 ) , .A1( u0_u1_n807 ) );
  NOR2_X1 u0_u1_U408 (.A1( u0_u1_n671 ) , .ZN( u0_u1_n675 ) , .A2( u0_u1_n746 ) );
  NOR2_X1 u0_u1_U409 (.ZN( u0_u1_n720 ) , .A2( u0_u1_n726 ) , .A1( u0_u1_n746 ) );
  NOR4_X1 u0_u1_U41 (.A4( u0_u1_n689 ) , .A3( u0_u1_n690 ) , .A2( u0_u1_n691 ) , .A1( u0_u1_n692 ) , .ZN( u0_u1_n693 ) );
  NOR2_X1 u0_u1_U410 (.ZN( u0_u1_n584 ) , .A1( u0_u1_n746 ) , .A2( u0_u1_n817 ) );
  INV_X1 u0_u1_U411 (.A( u0_u1_n746 ) , .ZN( u0_u1_n838 ) );
  AOI221_X1 u0_u1_U412 (.A( u0_u1_n578 ) , .ZN( u0_u1_n589 ) , .B2( u0_u1_n833 ) , .C2( u0_u1_n844 ) , .B1( u0_u1_n855 ) , .C1( u0_u1_n862 ) );
  AOI21_X1 u0_u1_U413 (.ZN( u0_u1_n578 ) , .B2( u0_u1_n726 ) , .B1( u0_u1_n750 ) , .A( u0_u1_n787 ) );
  AOI211_X1 u0_u1_U414 (.A( u0_u1_n639 ) , .ZN( u0_u1_n647 ) , .B( u0_u1_n745 ) , .C2( u0_u1_n840 ) , .C1( u0_u1_n855 ) );
  NAND4_X1 u0_u1_U415 (.A4( u0_u1_n635 ) , .A3( u0_u1_n636 ) , .A2( u0_u1_n637 ) , .A1( u0_u1_n638 ) , .ZN( u0_u1_n745 ) );
  OAI22_X1 u0_u1_U416 (.B1( u0_u1_n441 ) , .ZN( u0_u1_n590 ) , .A2( u0_u1_n749 ) , .B2( u0_u1_n764 ) , .A1( u0_u1_n765 ) );
  NAND2_X1 u0_u1_U417 (.A2( u0_u1_n441 ) , .A1( u0_u1_n731 ) , .ZN( u0_u1_n813 ) );
  AOI21_X1 u0_u1_U418 (.B2( u0_u1_n441 ) , .ZN( u0_u1_n594 ) , .B1( u0_u1_n730 ) , .A( u0_u1_n792 ) );
  AOI21_X1 u0_u1_U419 (.B2( u0_u1_n441 ) , .ZN( u0_u1_n650 ) , .A( u0_u1_n764 ) , .B1( u0_u1_n794 ) );
  AOI221_X1 u0_u1_U42 (.A( u0_u1_n683 ) , .ZN( u0_u1_n694 ) , .B2( u0_u1_n841 ) , .C1( u0_u1_n843 ) , .C2( u0_u1_n863 ) , .B1( u0_u1_n866 ) );
  AOI21_X1 u0_u1_U420 (.B2( u0_u1_n441 ) , .ZN( u0_u1_n625 ) , .B1( u0_u1_n701 ) , .A( u0_u1_n781 ) );
  OAI22_X1 u0_u1_U421 (.B2( u0_u1_n441 ) , .ZN( u0_u1_n683 ) , .A1( u0_u1_n701 ) , .A2( u0_u1_n732 ) , .B1( u0_u1_n819 ) );
  NOR2_X1 u0_u1_U422 (.ZN( u0_u1_n653 ) , .A1( u0_u1_n786 ) , .A2( u0_u1_n790 ) );
  OAI21_X1 u0_u1_U423 (.B2( u0_u1_n441 ) , .A( u0_u1_n615 ) , .ZN( u0_u1_n618 ) , .B1( u0_u1_n627 ) );
  NOR2_X1 u0_u1_U424 (.A1( u0_u1_n441 ) , .ZN( u0_u1_n612 ) , .A2( u0_u1_n818 ) );
  NOR2_X1 u0_u1_U425 (.ZN( u0_u1_n555 ) , .A2( u0_u1_n746 ) , .A1( u0_u1_n786 ) );
  NOR2_X1 u0_u1_U426 (.A2( u0_u1_n41 ) , .ZN( u0_u1_n602 ) , .A1( u0_u1_n786 ) );
  AOI21_X1 u0_u1_U427 (.A( u0_u1_n41 ) , .ZN( u0_u1_n502 ) , .B1( u0_u1_n710 ) , .B2( u0_u1_n788 ) );
  OAI22_X1 u0_u1_U428 (.ZN( u0_u1_n592 ) , .B1( u0_u1_n732 ) , .B2( u0_u1_n751 ) , .A2( u0_u1_n788 ) , .A1( u0_u1_n805 ) );
  AOI222_X1 u0_u1_U429 (.ZN( u0_u1_n515 ) , .C1( u0_u1_n834 ) , .B2( u0_u1_n838 ) , .A2( u0_u1_n844 ) , .C2( u0_u1_n863 ) , .B1( u0_u1_n864 ) , .A1( u0_u1_n867 ) );
  NOR4_X1 u0_u1_U43 (.A4( u0_u1_n528 ) , .A2( u0_u1_n529 ) , .A1( u0_u1_n530 ) , .ZN( u0_u1_n540 ) , .A3( u0_u1_n703 ) );
  AOI222_X1 u0_u1_U430 (.ZN( u0_u1_n607 ) , .B2( u0_u1_n673 ) , .B1( u0_u1_n755 ) , .C2( u0_u1_n833 ) , .A1( u0_u1_n835 ) , .A2( u0_u1_n863 ) , .C1( u0_u1_n864 ) );
  AOI221_X1 u0_u1_U431 (.A( u0_u1_n485 ) , .ZN( u0_u1_n490 ) , .B1( u0_u1_n833 ) , .C2( u0_u1_n845 ) , .C1( u0_u1_n853 ) , .B2( u0_u1_n863 ) );
  NOR2_X1 u0_u1_U432 (.ZN( u0_u1_n655 ) , .A1( u0_u1_n764 ) , .A2( u0_u1_n788 ) );
  NAND2_X1 u0_u1_U433 (.A2( u0_u1_n751 ) , .A1( u0_u1_n788 ) , .ZN( u0_u1_n811 ) );
  NOR2_X1 u0_u1_U434 (.ZN( u0_u1_n556 ) , .A1( u0_u1_n788 ) , .A2( u0_u1_n815 ) );
  NOR2_X1 u0_u1_U435 (.ZN( u0_u1_n614 ) , .A1( u0_u1_n781 ) , .A2( u0_u1_n788 ) );
  NOR2_X1 u0_u1_U436 (.ZN( u0_u1_n719 ) , .A2( u0_u1_n746 ) , .A1( u0_u1_n788 ) );
  NAND3_X1 u0_u1_U437 (.ZN( u0_subword_22 ) , .A3( u0_u1_n799 ) , .A2( u0_u1_n800 ) , .A1( u0_u1_n801 ) );
  NAND3_X1 u0_u1_U438 (.ZN( u0_subword_21 ) , .A3( u0_u1_n760 ) , .A2( u0_u1_n761 ) , .A1( u0_u1_n762 ) );
  NAND3_X1 u0_u1_U439 (.ZN( u0_subword_20 ) , .A3( u0_u1_n740 ) , .A2( u0_u1_n741 ) , .A1( u0_u1_n742 ) );
  NOR4_X1 u0_u1_U44 (.A4( u0_u1_n534 ) , .A3( u0_u1_n535 ) , .A2( u0_u1_n536 ) , .ZN( u0_u1_n537 ) , .A1( u0_u1_n822 ) );
  NAND3_X1 u0_u1_U440 (.A3( u0_u1_n677 ) , .A2( u0_u1_n678 ) , .A1( u0_u1_n679 ) , .ZN( u0_u1_n809 ) );
  NAND3_X1 u0_u1_U441 (.ZN( u0_u1_n640 ) , .A3( u0_u1_n710 ) , .A2( u0_u1_n726 ) , .A1( u0_u1_n794 ) );
  NAND3_X1 u0_u1_U442 (.A3( u0_u1_n620 ) , .A2( u0_u1_n621 ) , .A1( u0_u1_n622 ) , .ZN( u0_u1_n727 ) );
  NAND3_X1 u0_u1_U443 (.A3( u0_u1_n587 ) , .A2( u0_u1_n588 ) , .A1( u0_u1_n589 ) , .ZN( u0_u1_n623 ) );
  NAND3_X1 u0_u1_U444 (.ZN( u0_u1_n567 ) , .A3( u0_u1_n682 ) , .A2( u0_u1_n752 ) , .A1( u0_u1_n787 ) );
  NAND3_X1 u0_u1_U445 (.A3( u0_u1_n525 ) , .A2( u0_u1_n526 ) , .A1( u0_u1_n527 ) , .ZN( u0_u1_n744 ) );
  NAND3_X1 u0_u1_U446 (.A3( u0_u1_n514 ) , .A1( u0_u1_n515 ) , .ZN( u0_u1_n610 ) , .A2( u0_u1_n872 ) );
  NAND3_X1 u0_u1_U447 (.A3( u0_u1_n469 ) , .A2( u0_u1_n470 ) , .A1( u0_u1_n471 ) , .ZN( u0_u1_n779 ) );
  NOR2_X1 u0_u1_U448 (.ZN( u0_u1_n791 ) , .A2( u0_u1_n863 ) , .A1( u0_u1_n869 ) );
  NOR2_X1 u0_u1_U449 (.ZN( u0_u1_n703 ) , .A2( u0_u1_n788 ) , .A1( u0_u1_n819 ) );
  NOR4_X1 u0_u1_U45 (.A4( u0_u1_n531 ) , .A3( u0_u1_n532 ) , .ZN( u0_u1_n539 ) , .A2( u0_u1_n686 ) , .A1( u0_u1_n796 ) );
  NOR2_X1 u0_u1_U450 (.A1( u0_u1_n732 ) , .ZN( u0_u1_n767 ) , .A2( u0_u1_n788 ) );
  INV_X1 u0_u1_U451 (.A( u0_u1_n788 ) , .ZN( u0_u1_n863 ) );
  NOR3_X1 u0_u1_U46 (.A3( u0_u1_n802 ) , .A2( u0_u1_n803 ) , .A1( u0_u1_n804 ) , .ZN( u0_u1_n827 ) );
  NAND4_X1 u0_u1_U47 (.A4( u0_u1_n481 ) , .A3( u0_u1_n482 ) , .A2( u0_u1_n483 ) , .A1( u0_u1_n484 ) , .ZN( u0_u1_n696 ) );
  NOR3_X1 u0_u1_U48 (.ZN( u0_u1_n482 ) , .A2( u0_u1_n510 ) , .A3( u0_u1_n603 ) , .A1( u0_u1_n612 ) );
  NOR4_X1 u0_u1_U49 (.ZN( u0_u1_n481 ) , .A1( u0_u1_n522 ) , .A4( u0_u1_n559 ) , .A3( u0_u1_n584 ) , .A2( u0_u1_n632 ) );
  NOR3_X1 u0_u1_U5 (.ZN( u0_u1_n600 ) , .A1( u0_u1_n610 ) , .A3( u0_u1_n725 ) , .A2( u0_u1_n744 ) );
  NAND4_X1 u0_u1_U50 (.A4( u0_u1_n774 ) , .A3( u0_u1_n775 ) , .A2( u0_u1_n776 ) , .A1( u0_u1_n777 ) , .ZN( u0_u1_n803 ) );
  NOR3_X1 u0_u1_U51 (.A3( u0_u1_n767 ) , .A2( u0_u1_n768 ) , .A1( u0_u1_n769 ) , .ZN( u0_u1_n775 ) );
  NOR4_X1 u0_u1_U52 (.A4( u0_u1_n770 ) , .A3( u0_u1_n771 ) , .A2( u0_u1_n772 ) , .A1( u0_u1_n773 ) , .ZN( u0_u1_n774 ) );
  NAND4_X1 u0_u1_U53 (.A4( u0_u1_n562 ) , .A3( u0_u1_n563 ) , .A2( u0_u1_n564 ) , .A1( u0_u1_n565 ) , .ZN( u0_u1_n609 ) );
  NOR4_X1 u0_u1_U54 (.A4( u0_u1_n554 ) , .A3( u0_u1_n555 ) , .A2( u0_u1_n556 ) , .A1( u0_u1_n557 ) , .ZN( u0_u1_n564 ) );
  AOI222_X1 u0_u1_U55 (.ZN( u0_u1_n565 ) , .B1( u0_u1_n832 ) , .C1( u0_u1_n842 ) , .A2( u0_u1_n844 ) , .A1( u0_u1_n855 ) , .B2( u0_u1_n864 ) , .C2( u0_u1_n874 ) );
  NOR4_X1 u0_u1_U56 (.A4( u0_u1_n558 ) , .A3( u0_u1_n559 ) , .A2( u0_u1_n560 ) , .A1( u0_u1_n561 ) , .ZN( u0_u1_n562 ) );
  INV_X1 u0_u1_U57 (.A( u0_u1_n507 ) , .ZN( u0_u1_n872 ) );
  NOR4_X1 u0_u1_U58 (.A4( u0_u1_n511 ) , .A2( u0_u1_n512 ) , .A1( u0_u1_n513 ) , .ZN( u0_u1_n514 ) , .A3( u0_u1_n672 ) );
  NOR4_X1 u0_u1_U59 (.A4( u0_u1_n663 ) , .A3( u0_u1_n664 ) , .A2( u0_u1_n665 ) , .A1( u0_u1_n666 ) , .ZN( u0_u1_n679 ) );
  NOR3_X1 u0_u1_U6 (.A2( u0_u1_n609 ) , .A1( u0_u1_n610 ) , .ZN( u0_u1_n648 ) , .A3( u0_u1_n724 ) );
  NOR4_X1 u0_u1_U60 (.A4( u0_u1_n667 ) , .A3( u0_u1_n668 ) , .A2( u0_u1_n669 ) , .A1( u0_u1_n670 ) , .ZN( u0_u1_n678 ) );
  NOR4_X1 u0_u1_U61 (.A3( u0_u1_n675 ) , .A1( u0_u1_n676 ) , .ZN( u0_u1_n677 ) , .A4( u0_u1_n717 ) , .A2( u0_u1_n860 ) );
  AOI221_X1 u0_u1_U62 (.ZN( u0_u1_n470 ) , .C2( u0_u1_n716 ) , .B2( u0_u1_n833 ) , .C1( u0_u1_n846 ) , .B1( u0_u1_n861 ) , .A( u0_u1_n865 ) );
  NOR4_X1 u0_u1_U63 (.A1( u0_u1_n468 ) , .ZN( u0_u1_n469 ) , .A4( u0_u1_n544 ) , .A2( u0_u1_n556 ) , .A3( u0_u1_n616 ) );
  NAND4_X1 u0_u1_U64 (.A4( u0_u1_n487 ) , .A3( u0_u1_n488 ) , .A2( u0_u1_n489 ) , .A1( u0_u1_n490 ) , .ZN( u0_u1_n780 ) );
  NOR4_X1 u0_u1_U65 (.A4( u0_u1_n486 ) , .ZN( u0_u1_n489 ) , .A1( u0_u1_n568 ) , .A2( u0_u1_n583 ) , .A3( u0_u1_n604 ) );
  NOR4_X1 u0_u1_U66 (.ZN( u0_u1_n488 ) , .A1( u0_u1_n509 ) , .A2( u0_u1_n521 ) , .A4( u0_u1_n548 ) , .A3( u0_u1_n613 ) );
  NOR2_X1 u0_u1_U67 (.ZN( u0_u1_n763 ) , .A1( u0_u1_n835 ) , .A2( u0_u1_n836 ) );
  NOR4_X1 u0_u1_U68 (.A4( u0_u1_n516 ) , .A3( u0_u1_n517 ) , .A2( u0_u1_n518 ) , .A1( u0_u1_n519 ) , .ZN( u0_u1_n526 ) );
  NOR4_X1 u0_u1_U69 (.A3( u0_u1_n523 ) , .A1( u0_u1_n524 ) , .ZN( u0_u1_n525 ) , .A2( u0_u1_n675 ) , .A4( u0_u1_n771 ) );
  NOR3_X1 u0_u1_U7 (.A3( u0_u1_n724 ) , .A1( u0_u1_n725 ) , .ZN( u0_u1_n742 ) , .A2( u0_u1_n743 ) );
  NAND4_X1 u0_u1_U70 (.A4( u0_u1_n475 ) , .A3( u0_u1_n476 ) , .A2( u0_u1_n477 ) , .A1( u0_u1_n478 ) , .ZN( u0_u1_n680 ) );
  NOR4_X1 u0_u1_U71 (.ZN( u0_u1_n476 ) , .A1( u0_u1_n508 ) , .A3( u0_u1_n546 ) , .A2( u0_u1_n585 ) , .A4( u0_u1_n718 ) );
  NOR4_X1 u0_u1_U72 (.ZN( u0_u1_n475 ) , .A2( u0_u1_n523 ) , .A4( u0_u1_n596 ) , .A1( u0_u1_n611 ) , .A3( u0_u1_n631 ) );
  NOR4_X1 u0_u1_U73 (.A4( u0_u1_n472 ) , .ZN( u0_u1_n478 ) , .A3( u0_u1_n558 ) , .A1( u0_u1_n737 ) , .A2( u0_u1_n757 ) );
  NAND4_X1 u0_u1_U74 (.A4( u0_u1_n458 ) , .A3( u0_u1_n459 ) , .A2( u0_u1_n460 ) , .A1( u0_u1_n461 ) , .ZN( u0_u1_n681 ) );
  NOR3_X1 u0_u1_U75 (.ZN( u0_u1_n459 ) , .A3( u0_u1_n532 ) , .A1( u0_u1_n557 ) , .A2( u0_u1_n572 ) );
  AOI221_X1 u0_u1_U76 (.A( u0_u1_n452 ) , .ZN( u0_u1_n461 ) , .C2( u0_u1_n755 ) , .B1( u0_u1_n834 ) , .C1( u0_u1_n843 ) , .B2( u0_u1_n862 ) );
  NOR4_X1 u0_u1_U77 (.ZN( u0_u1_n460 ) , .A2( u0_u1_n511 ) , .A1( u0_u1_n601 ) , .A4( u0_u1_n630 ) , .A3( u0_u1_n713 ) );
  INV_X1 u0_u1_U78 (.A( u0_u1_n671 ) , .ZN( u0_u1_n866 ) );
  NAND4_X1 u0_u1_U79 (.A4( u0_u1_n575 ) , .A3( u0_u1_n576 ) , .A1( u0_u1_n577 ) , .ZN( u0_u1_n725 ) , .A2( u0_u1_n875 ) );
  NOR3_X1 u0_u1_U8 (.ZN( u0_u1_n506 ) , .A2( u0_u1_n681 ) , .A3( u0_u1_n779 ) , .A1( u0_u1_n877 ) );
  NOR4_X1 u0_u1_U80 (.A4( u0_u1_n571 ) , .A3( u0_u1_n572 ) , .A2( u0_u1_n573 ) , .A1( u0_u1_n574 ) , .ZN( u0_u1_n575 ) );
  AOI221_X1 u0_u1_U81 (.A( u0_u1_n566 ) , .C2( u0_u1_n567 ) , .ZN( u0_u1_n576 ) , .B2( u0_u1_n846 ) , .B1( u0_u1_n853 ) , .C1( u0_u1_n854 ) );
  NOR2_X1 u0_u1_U82 (.ZN( u0_u1_n577 ) , .A1( u0_u1_n624 ) , .A2( u0_u1_n747 ) );
  INV_X1 u0_u1_U83 (.A( u0_u1_n764 ) , .ZN( u0_u1_n832 ) );
  NOR2_X1 u0_u1_U84 (.ZN( u0_u1_n649 ) , .A1( u0_u1_n855 ) , .A2( u0_u1_n869 ) );
  NOR4_X1 u0_u1_U85 (.A4( u0_u1_n579 ) , .A3( u0_u1_n580 ) , .A2( u0_u1_n581 ) , .ZN( u0_u1_n588 ) , .A1( u0_u1_n685 ) );
  NOR4_X1 u0_u1_U86 (.A1( u0_u1_n586 ) , .ZN( u0_u1_n587 ) , .A3( u0_u1_n654 ) , .A2( u0_u1_n664 ) , .A4( u0_u1_n769 ) );
  NAND4_X1 u0_u1_U87 (.A4( u0_u1_n721 ) , .A3( u0_u1_n722 ) , .A2( u0_u1_n723 ) , .ZN( u0_u1_n743 ) , .A1( u0_u1_n858 ) );
  NOR4_X1 u0_u1_U88 (.A4( u0_u1_n717 ) , .A3( u0_u1_n718 ) , .A2( u0_u1_n719 ) , .A1( u0_u1_n720 ) , .ZN( u0_u1_n721 ) );
  INV_X1 u0_u1_U89 (.A( u0_u1_n711 ) , .ZN( u0_u1_n858 ) );
  NOR2_X1 u0_u1_U9 (.ZN( u0_u1_n497 ) , .A1( u0_u1_n680 ) , .A2( u0_u1_n696 ) );
  AOI221_X1 u0_u1_U90 (.A( u0_u1_n712 ) , .ZN( u0_u1_n723 ) , .C2( u0_u1_n845 ) , .B2( u0_u1_n846 ) , .C1( u0_u1_n862 ) , .B1( u0_u1_n863 ) );
  INV_X1 u0_u1_U91 (.A( u0_u1_n465 ) , .ZN( u0_u1_n865 ) );
  OAI21_X1 u0_u1_U92 (.ZN( u0_u1_n465 ) , .B1( u0_u1_n811 ) , .A( u0_u1_n836 ) , .B2( u0_u1_n852 ) );
  INV_X1 u0_u1_U93 (.A( u0_u1_n793 ) , .ZN( u0_u1_n874 ) );
  OR4_X1 u0_u1_U94 (.A4( u0_u1_n568 ) , .A3( u0_u1_n569 ) , .A2( u0_u1_n570 ) , .ZN( u0_u1_n574 ) , .A1( u0_u1_n667 ) );
  OR4_X1 u0_u1_U95 (.A4( u0_u1_n520 ) , .A2( u0_u1_n521 ) , .A1( u0_u1_n522 ) , .ZN( u0_u1_n524 ) , .A3( u0_u1_n823 ) );
  OR4_X1 u0_u1_U96 (.ZN( u0_u1_n494 ) , .A4( u0_u1_n536 ) , .A2( u0_u1_n549 ) , .A1( u0_u1_n561 ) , .A3( u0_u1_n634 ) );
  OR4_X1 u0_u1_U97 (.ZN( u0_u1_n468 ) , .A4( u0_u1_n520 ) , .A3( u0_u1_n531 ) , .A2( u0_u1_n580 ) , .A1( u0_u1_n714 ) );
  OR4_X1 u0_u1_U98 (.A4( u0_u1_n684 ) , .A3( u0_u1_n685 ) , .A2( u0_u1_n686 ) , .A1( u0_u1_n687 ) , .ZN( u0_u1_n692 ) );
  OR3_X1 u0_u1_U99 (.A3( u0_u1_n508 ) , .A2( u0_u1_n509 ) , .A1( u0_u1_n510 ) , .ZN( u0_u1_n513 ) );
  NOR2_X1 us02_U10 (.ZN( us02_n574 ) , .A1( us02_n621 ) , .A2( us02_n744 ) );
  NOR2_X1 us02_U100 (.ZN( us02_n685 ) , .A1( us02_n830 ) , .A2( us02_n831 ) );
  NOR4_X1 us02_U101 (.ZN( us02_n619 ) , .A1( us02_n655 ) , .A3( us02_n665 ) , .A4( us02_n681 ) , .A2( us02_n765 ) );
  NOR4_X1 us02_U102 (.A4( us02_n608 ) , .A3( us02_n609 ) , .A2( us02_n610 ) , .A1( us02_n611 ) , .ZN( us02_n618 ) );
  NOR4_X1 us02_U103 (.A4( us02_n613 ) , .A3( us02_n614 ) , .A2( us02_n615 ) , .A1( us02_n616 ) , .ZN( us02_n617 ) );
  NAND4_X1 us02_U104 (.A4( us02_n484 ) , .A3( us02_n485 ) , .A2( us02_n486 ) , .A1( us02_n487 ) , .ZN( us02_n777 ) );
  NOR4_X1 us02_U105 (.A4( us02_n483 ) , .ZN( us02_n486 ) , .A1( us02_n565 ) , .A2( us02_n580 ) , .A3( us02_n601 ) );
  NOR4_X1 us02_U106 (.ZN( us02_n485 ) , .A1( us02_n506 ) , .A2( us02_n518 ) , .A4( us02_n545 ) , .A3( us02_n610 ) );
  NOR4_X1 us02_U107 (.ZN( us02_n484 ) , .A2( us02_n532 ) , .A1( us02_n557 ) , .A3( us02_n630 ) , .A4( us02_n717 ) );
  NAND4_X1 us02_U108 (.A4( us02_n690 ) , .A3( us02_n691 ) , .A1( us02_n692 ) , .ZN( us02_n775 ) , .A2( us02_n871 ) );
  AOI221_X1 us02_U109 (.A( us02_n680 ) , .ZN( us02_n691 ) , .B2( us02_n839 ) , .C1( us02_n841 ) , .C2( us02_n861 ) , .B1( us02_n864 ) );
  NOR2_X1 us02_U11 (.A1( us02_n677 ) , .ZN( us02_n692 ) , .A2( us02_n806 ) );
  INV_X1 us02_U110 (.A( us02_n678 ) , .ZN( us02_n871 ) );
  NOR4_X1 us02_U111 (.A4( us02_n686 ) , .A3( us02_n687 ) , .A2( us02_n688 ) , .A1( us02_n689 ) , .ZN( us02_n690 ) );
  NAND4_X1 us02_U112 (.A4( us02_n559 ) , .A3( us02_n560 ) , .A2( us02_n561 ) , .A1( us02_n562 ) , .ZN( us02_n606 ) );
  NOR4_X1 us02_U113 (.ZN( us02_n560 ) , .A1( us02_n652 ) , .A3( us02_n660 ) , .A4( us02_n684 ) , .A2( us02_n767 ) );
  NOR4_X1 us02_U114 (.A4( us02_n551 ) , .A3( us02_n552 ) , .A2( us02_n553 ) , .A1( us02_n554 ) , .ZN( us02_n561 ) );
  NOR4_X1 us02_U115 (.A4( us02_n555 ) , .A3( us02_n556 ) , .A2( us02_n557 ) , .A1( us02_n558 ) , .ZN( us02_n559 ) );
  NAND4_X1 us02_U116 (.A4( us02_n718 ) , .A3( us02_n719 ) , .A2( us02_n720 ) , .ZN( us02_n740 ) , .A1( us02_n856 ) );
  INV_X1 us02_U117 (.A( us02_n708 ) , .ZN( us02_n856 ) );
  AOI221_X1 us02_U118 (.A( us02_n709 ) , .ZN( us02_n720 ) , .C2( us02_n843 ) , .B2( us02_n844 ) , .C1( us02_n860 ) , .B1( us02_n861 ) );
  NOR4_X1 us02_U119 (.A4( us02_n714 ) , .A3( us02_n715 ) , .A2( us02_n716 ) , .A1( us02_n717 ) , .ZN( us02_n718 ) );
  INV_X1 us02_U12 (.A( us02_n679 ) , .ZN( us02_n839 ) );
  NAND4_X1 us02_U120 (.A4( us02_n472 ) , .A3( us02_n473 ) , .A2( us02_n474 ) , .A1( us02_n475 ) , .ZN( us02_n677 ) );
  NOR4_X1 us02_U121 (.A4( us02_n469 ) , .ZN( us02_n475 ) , .A3( us02_n555 ) , .A1( us02_n734 ) , .A2( us02_n754 ) );
  NOR4_X1 us02_U122 (.ZN( us02_n474 ) , .A1( us02_n530 ) , .A3( us02_n567 ) , .A4( us02_n599 ) , .A2( us02_n641 ) );
  NOR4_X1 us02_U123 (.ZN( us02_n473 ) , .A1( us02_n505 ) , .A3( us02_n543 ) , .A2( us02_n582 ) , .A4( us02_n715 ) );
  NOR2_X1 us02_U124 (.ZN( us02_n732 ) , .A2( us02_n831 ) , .A1( us02_n844 ) );
  NOR2_X1 us02_U125 (.ZN( us02_n788 ) , .A2( us02_n861 ) , .A1( us02_n867 ) );
  NOR2_X1 us02_U126 (.ZN( us02_n646 ) , .A1( us02_n853 ) , .A2( us02_n867 ) );
  NAND4_X1 us02_U127 (.A4( us02_n572 ) , .A3( us02_n573 ) , .A1( us02_n574 ) , .ZN( us02_n722 ) , .A2( us02_n873 ) );
  NOR4_X1 us02_U128 (.A4( us02_n568 ) , .A3( us02_n569 ) , .A2( us02_n570 ) , .A1( us02_n571 ) , .ZN( us02_n572 ) );
  AOI221_X1 us02_U129 (.A( us02_n563 ) , .C2( us02_n564 ) , .ZN( us02_n573 ) , .B2( us02_n844 ) , .B1( us02_n851 ) , .C1( us02_n852 ) );
  NOR4_X1 us02_U13 (.A4( us02_n444 ) , .A3( us02_n445 ) , .A2( us02_n515 ) , .A1( us02_n540 ) , .ZN( us02_n705 ) );
  INV_X1 us02_U130 (.A( us02_n606 ) , .ZN( us02_n873 ) );
  NAND4_X1 us02_U131 (.A4( us02_n492 ) , .A3( us02_n493 ) , .A1( us02_n494 ) , .ZN( us02_n801 ) , .A2( us02_n866 ) );
  AOI221_X1 us02_U132 (.A( us02_n488 ) , .ZN( us02_n493 ) , .B2( us02_n835 ) , .C2( us02_n840 ) , .C1( us02_n850 ) , .B1( us02_n859 ) );
  INV_X1 us02_U133 (.A( us02_n777 ) , .ZN( us02_n866 ) );
  NOR2_X1 us02_U134 (.ZN( us02_n494 ) , .A1( us02_n677 ) , .A2( us02_n693 ) );
  AOI222_X1 us02_U135 (.ZN( us02_n512 ) , .C1( us02_n831 ) , .B2( us02_n836 ) , .A2( us02_n842 ) , .C2( us02_n861 ) , .B1( us02_n862 ) , .A1( us02_n865 ) );
  NOR4_X1 us02_U136 (.A4( us02_n508 ) , .A2( us02_n509 ) , .A1( us02_n510 ) , .ZN( us02_n511 ) , .A3( us02_n669 ) );
  INV_X1 us02_U137 (.A( us02_n504 ) , .ZN( us02_n870 ) );
  INV_X1 us02_U138 (.A( us02_n761 ) , .ZN( us02_n829 ) );
  INV_X1 us02_U139 (.A( us02_n462 ) , .ZN( us02_n863 ) );
  OR3_X1 us02_U14 (.ZN( us02_n445 ) , .A1( us02_n527 ) , .A3( us02_n576 ) , .A2( us02_n874 ) );
  OAI21_X1 us02_U140 (.ZN( us02_n462 ) , .B1( us02_n808 ) , .A( us02_n833 ) , .B2( us02_n850 ) );
  OR4_X1 us02_U141 (.A4( us02_n565 ) , .A3( us02_n566 ) , .A2( us02_n567 ) , .ZN( us02_n571 ) , .A1( us02_n664 ) );
  OR4_X1 us02_U142 (.A4( us02_n517 ) , .A2( us02_n518 ) , .A1( us02_n519 ) , .ZN( us02_n521 ) , .A3( us02_n820 ) );
  OR4_X1 us02_U143 (.ZN( us02_n465 ) , .A4( us02_n517 ) , .A3( us02_n528 ) , .A2( us02_n577 ) , .A1( us02_n711 ) );
  OR4_X1 us02_U144 (.A4( us02_n681 ) , .A3( us02_n682 ) , .A2( us02_n683 ) , .A1( us02_n684 ) , .ZN( us02_n689 ) );
  OR4_X1 us02_U145 (.A4( us02_n579 ) , .A3( us02_n580 ) , .A2( us02_n581 ) , .A1( us02_n582 ) , .ZN( us02_n583 ) );
  NAND2_X1 us02_U146 (.ZN( us02_n612 ) , .A2( us02_n836 ) , .A1( us02_n872 ) );
  OR3_X1 us02_U147 (.A3( us02_n505 ) , .A2( us02_n506 ) , .A1( us02_n507 ) , .ZN( us02_n510 ) );
  AOI221_X1 us02_U148 (.A( us02_n712 ) , .B2( us02_n713 ) , .ZN( us02_n719 ) , .C1( us02_n831 ) , .B1( us02_n838 ) , .C2( us02_n862 ) );
  OR2_X1 us02_U149 (.A2( us02_n710 ) , .A1( us02_n711 ) , .ZN( us02_n712 ) );
  OR4_X1 us02_U15 (.A4( us02_n441 ) , .A2( us02_n442 ) , .A1( us02_n443 ) , .ZN( us02_n444 ) , .A3( us02_n552 ) );
  INV_X1 us02_U150 (.A( us02_n753 ) , .ZN( us02_n868 ) );
  OAI21_X1 us02_U151 (.B1( us02_n752 ) , .ZN( us02_n753 ) , .A( us02_n844 ) , .B2( us02_n867 ) );
  INV_X1 us02_U152 (.A( us02_n671 ) , .ZN( us02_n858 ) );
  AOI21_X1 us02_U153 (.A( us02_n669 ) , .B1( us02_n670 ) , .ZN( us02_n671 ) , .B2( us02_n855 ) );
  NAND2_X1 us02_U154 (.A1( us02_n446 ) , .A2( us02_n464 ) , .ZN( us02_n748 ) );
  OAI222_X1 us02_U155 (.B2( us02_n746 ) , .B1( us02_n747 ) , .A2( us02_n748 ) , .ZN( us02_n756 ) , .C2( us02_n804 ) , .C1( us02_n813 ) , .A1( us02_n816 ) );
  OAI222_X1 us02_U156 (.ZN( us02_n504 ) , .C2( us02_n624 ) , .B2( us02_n646 ) , .B1( us02_n746 ) , .A2( us02_n747 ) , .C1( us02_n804 ) , .A1( us02_n805 ) );
  OAI222_X1 us02_U157 (.B2( us02_n707 ) , .ZN( us02_n708 ) , .C2( us02_n723 ) , .B1( us02_n746 ) , .A1( us02_n805 ) , .C1( us02_n813 ) , .A2( us02_n814 ) );
  OAI222_X1 us02_U158 (.ZN( us02_n616 ) , .B1( us02_n696 ) , .C1( us02_n723 ) , .C2( us02_n746 ) , .B2( us02_n785 ) , .A2( us02_n791 ) , .A1( us02_n815 ) );
  NOR4_X1 us02_U159 (.A2( us02_n490 ) , .A1( us02_n491 ) , .ZN( us02_n492 ) , .A3( us02_n579 ) , .A4( us02_n611 ) );
  INV_X1 us02_U16 (.A( us02_n612 ) , .ZN( us02_n874 ) );
  OR4_X1 us02_U160 (.ZN( us02_n491 ) , .A4( us02_n533 ) , .A2( us02_n546 ) , .A1( us02_n558 ) , .A3( us02_n631 ) );
  OAI22_X1 us02_U161 (.B1( us02_n489 ) , .ZN( us02_n490 ) , .A1( us02_n685 ) , .A2( us02_n762 ) , .B2( us02_n816 ) );
  NOR3_X1 us02_U162 (.ZN( us02_n489 ) , .A1( us02_n781 ) , .A2( us02_n849 ) , .A3( us02_n862 ) );
  AOI22_X1 us02_U163 (.ZN( us02_n695 ) , .A1( us02_n829 ) , .B2( us02_n842 ) , .A2( us02_n864 ) , .B1( us02_n867 ) );
  INV_X1 us02_U164 (.A( us02_n729 ) , .ZN( us02_n838 ) );
  AOI221_X1 us02_U165 (.A( us02_n763 ) , .ZN( us02_n773 ) , .C2( us02_n809 ) , .B2( us02_n834 ) , .C1( us02_n854 ) , .B1( us02_n865 ) );
  AOI21_X1 us02_U166 (.B2( us02_n762 ) , .ZN( us02_n763 ) , .A( us02_n787 ) , .B1( us02_n791 ) );
  INV_X1 us02_U167 (.A( us02_n760 ) , .ZN( us02_n834 ) );
  AOI221_X1 us02_U168 (.A( us02_n482 ) , .ZN( us02_n487 ) , .B1( us02_n830 ) , .C2( us02_n843 ) , .C1( us02_n851 ) , .B2( us02_n861 ) );
  OAI22_X1 us02_U169 (.ZN( us02_n482 ) , .A1( us02_n707 ) , .B2( us02_n784 ) , .A2( us02_n805 ) , .B1( us02_n811 ) );
  INV_X1 us02_U17 (.A( us02_n748 ) , .ZN( us02_n862 ) );
  INV_X1 us02_U170 (.A( us02_n789 ) , .ZN( us02_n831 ) );
  NAND2_X1 us02_U171 (.A1( us02_n450 ) , .A2( us02_n452 ) , .ZN( us02_n761 ) );
  OAI221_X1 us02_U172 (.A( us02_n726 ) , .C2( us02_n727 ) , .B2( us02_n728 ) , .B1( us02_n729 ) , .ZN( us02_n736 ) , .C1( us02_n816 ) );
  AOI22_X1 us02_U173 (.ZN( us02_n726 ) , .B1( us02_n831 ) , .A2( us02_n837 ) , .A1( us02_n862 ) , .B2( us02_n865 ) );
  INV_X1 us02_U174 (.A( us02_n785 ) , .ZN( us02_n861 ) );
  OAI22_X1 us02_U175 (.ZN( us02_n709 ) , .A2( us02_n727 ) , .B2( us02_n728 ) , .A1( us02_n743 ) , .B1( us02_n812 ) );
  INV_X1 us02_U176 (.A( us02_n815 ) , .ZN( us02_n830 ) );
  OAI22_X1 us02_U177 (.ZN( us02_n488 ) , .A1( us02_n723 ) , .B2( us02_n727 ) , .B1( us02_n729 ) , .A2( us02_n778 ) );
  OAI22_X1 us02_U178 (.ZN( us02_n623 ) , .B1( us02_n668 ) , .B2( us02_n746 ) , .A1( us02_n814 ) , .A2( us02_n815 ) );
  INV_X1 us02_U179 (.A( us02_n743 ) , .ZN( us02_n836 ) );
  AOI222_X1 us02_U18 (.ZN( us02_n604 ) , .B2( us02_n670 ) , .B1( us02_n752 ) , .C2( us02_n830 ) , .A1( us02_n832 ) , .A2( us02_n861 ) , .C1( us02_n862 ) );
  OAI22_X1 us02_U180 (.A1( us02_n723 ) , .ZN( us02_n725 ) , .B2( us02_n749 ) , .B1( us02_n811 ) , .A2( us02_n815 ) );
  OAI22_X1 us02_U181 (.B2( us02_n778 ) , .B1( us02_n779 ) , .ZN( us02_n780 ) , .A2( us02_n813 ) , .A1( us02_n814 ) );
  INV_X1 us02_U182 (.A( us02_n787 ) , .ZN( us02_n844 ) );
  INV_X1 us02_U183 (.A( us02_n804 ) , .ZN( us02_n859 ) );
  INV_X1 us02_U184 (.A( us02_n813 ) , .ZN( us02_n832 ) );
  OAI22_X1 us02_U185 (.B2( us02_n743 ) , .ZN( us02_n745 ) , .A2( us02_n761 ) , .B1( us02_n779 ) , .A1( us02_n791 ) );
  OAI22_X1 us02_U186 (.B2( us02_n802 ) , .B1( us02_n803 ) , .A2( us02_n804 ) , .A1( us02_n805 ) , .ZN( us02_n807 ) );
  OAI22_X1 us02_U187 (.ZN( us02_n495 ) , .A2( us02_n743 ) , .A1( us02_n779 ) , .B1( us02_n790 ) , .B2( us02_n805 ) );
  OAI22_X1 us02_U188 (.ZN( us02_n589 ) , .B1( us02_n729 ) , .B2( us02_n748 ) , .A2( us02_n785 ) , .A1( us02_n802 ) );
  OAI22_X1 us02_U189 (.ZN( us02_n694 ) , .A2( us02_n729 ) , .A1( us02_n779 ) , .B1( us02_n790 ) , .B2( us02_n816 ) );
  AOI222_X1 us02_U19 (.ZN( us02_n562 ) , .B1( us02_n829 ) , .C1( us02_n840 ) , .A2( us02_n842 ) , .A1( us02_n853 ) , .B2( us02_n862 ) , .C2( us02_n872 ) );
  INV_X1 us02_U190 (.A( us02_n802 ) , .ZN( us02_n842 ) );
  INV_X1 us02_U191 (.A( us02_n668 ) , .ZN( us02_n864 ) );
  OAI22_X1 us02_U192 (.ZN( us02_n636 ) , .A1( us02_n698 ) , .B2( us02_n727 ) , .A2( us02_n761 ) , .B1( us02_n815 ) );
  NOR2_X1 us02_U193 (.ZN( us02_n714 ) , .A1( us02_n804 ) , .A2( us02_n816 ) );
  NOR2_X1 us02_U194 (.A1( us02_n696 ) , .ZN( us02_n769 ) , .A2( us02_n814 ) );
  NOR2_X1 us02_U195 (.ZN( us02_n665 ) , .A1( us02_n727 ) , .A2( us02_n802 ) );
  NOR2_X1 us02_U196 (.ZN( us02_n593 ) , .A2( us02_n696 ) , .A1( us02_n727 ) );
  NOR2_X1 us02_U197 (.ZN( us02_n569 ) , .A1( us02_n727 ) , .A2( us02_n805 ) );
  NOR2_X1 us02_U198 (.A2( us02_n743 ) , .ZN( us02_n754 ) , .A1( us02_n804 ) );
  NOR2_X1 us02_U199 (.ZN( us02_n717 ) , .A2( us02_n723 ) , .A1( us02_n743 ) );
  AOI222_X1 us02_U20 (.ZN( us02_n659 ) , .A2( us02_n838 ) , .B1( us02_n840 ) , .C2( us02_n844 ) , .A1( us02_n859 ) , .C1( us02_n862 ) , .B2( us02_n869 ) );
  NOR2_X1 us02_U200 (.ZN( us02_n734 ) , .A2( us02_n802 ) , .A1( us02_n804 ) );
  NOR2_X1 us02_U201 (.ZN( us02_n545 ) , .A2( us02_n779 ) , .A1( us02_n813 ) );
  NOR2_X1 us02_U202 (.ZN( us02_n576 ) , .A2( us02_n698 ) , .A1( us02_n813 ) );
  NOR2_X1 us02_U203 (.ZN( us02_n653 ) , .A1( us02_n727 ) , .A2( us02_n812 ) );
  NOR2_X1 us02_U204 (.ZN( us02_n611 ) , .A1( us02_n778 ) , .A2( us02_n785 ) );
  INV_X1 us02_U205 (.A( us02_n749 ) , .ZN( us02_n841 ) );
  NOR2_X1 us02_U206 (.ZN( us02_n531 ) , .A2( us02_n748 ) , .A1( us02_n749 ) );
  NOR2_X1 us02_U207 (.ZN( us02_n628 ) , .A2( us02_n727 ) , .A1( us02_n784 ) );
  NOR2_X1 us02_U208 (.ZN( us02_n614 ) , .A1( us02_n784 ) , .A2( us02_n814 ) );
  NOR2_X1 us02_U209 (.ZN( us02_n600 ) , .A2( us02_n779 ) , .A1( us02_n802 ) );
  INV_X1 us02_U21 (.A( us02_n646 ) , .ZN( us02_n869 ) );
  NOR2_X1 us02_U210 (.ZN( us02_n610 ) , .A2( us02_n779 ) , .A1( us02_n805 ) );
  INV_X1 us02_U211 (.A( us02_n746 ) , .ZN( us02_n833 ) );
  NOR2_X1 us02_U212 (.A2( us02_n743 ) , .ZN( us02_n768 ) , .A1( us02_n811 ) );
  NOR2_X1 us02_U213 (.ZN( us02_n527 ) , .A2( us02_n723 ) , .A1( us02_n802 ) );
  NOR2_X1 us02_U214 (.ZN( us02_n530 ) , .A2( us02_n779 ) , .A1( us02_n815 ) );
  NOR2_X1 us02_U215 (.ZN( us02_n627 ) , .A2( us02_n668 ) , .A1( us02_n784 ) );
  NOR2_X1 us02_U216 (.ZN( us02_n598 ) , .A2( us02_n790 ) , .A1( us02_n815 ) );
  INV_X1 us02_U217 (.A( us02_n727 ) , .ZN( us02_n851 ) );
  NOR2_X1 us02_U218 (.ZN( us02_n651 ) , .A1( us02_n668 ) , .A2( us02_n813 ) );
  NOR2_X1 us02_U219 (.A1( us02_n668 ) , .ZN( us02_n672 ) , .A2( us02_n743 ) );
  NOR4_X1 us02_U22 (.ZN( us02_n472 ) , .A2( us02_n520 ) , .A4( us02_n593 ) , .A1( us02_n608 ) , .A3( us02_n628 ) );
  NOR2_X1 us02_U220 (.ZN( us02_n601 ) , .A1( us02_n668 ) , .A2( us02_n802 ) );
  NOR2_X1 us02_U221 (.A1( us02_n668 ) , .ZN( us02_n687 ) , .A2( us02_n815 ) );
  INV_X1 us02_U222 (.A( us02_n791 ) , .ZN( us02_n850 ) );
  NOR2_X1 us02_U223 (.A2( us02_n707 ) , .A1( us02_n749 ) , .ZN( us02_n770 ) );
  NOR2_X1 us02_U224 (.A1( us02_n668 ) , .ZN( us02_n765 ) , .A2( us02_n812 ) );
  NOR2_X1 us02_U225 (.A1( us02_n698 ) , .ZN( us02_n767 ) , .A2( us02_n812 ) );
  NOR2_X1 us02_U226 (.ZN( us02_n540 ) , .A2( us02_n696 ) , .A1( us02_n698 ) );
  NOR2_X1 us02_U227 (.ZN( us02_n526 ) , .A1( us02_n668 ) , .A2( us02_n778 ) );
  NOR2_X1 us02_U228 (.ZN( us02_n666 ) , .A1( us02_n749 ) , .A2( us02_n814 ) );
  NOR2_X1 us02_U229 (.ZN( us02_n554 ) , .A1( us02_n749 ) , .A2( us02_n790 ) );
  NOR4_X1 us02_U23 (.ZN( us02_n478 ) , .A1( us02_n519 ) , .A4( us02_n556 ) , .A3( us02_n581 ) , .A2( us02_n629 ) );
  NOR2_X1 us02_U230 (.ZN( us02_n507 ) , .A2( us02_n779 ) , .A1( us02_n784 ) );
  NOR2_X1 us02_U231 (.ZN( us02_n542 ) , .A2( us02_n707 ) , .A1( us02_n784 ) );
  NOR2_X1 us02_U232 (.ZN( us02_n663 ) , .A1( us02_n784 ) , .A2( us02_n790 ) );
  NOR2_X1 us02_U233 (.A2( us02_n696 ) , .ZN( us02_n715 ) , .A1( us02_n791 ) );
  NOR2_X1 us02_U234 (.ZN( us02_n506 ) , .A1( us02_n811 ) , .A2( us02_n816 ) );
  NOR2_X1 us02_U235 (.ZN( us02_n555 ) , .A1( us02_n761 ) , .A2( us02_n804 ) );
  NOR2_X1 us02_U236 (.ZN( us02_n660 ) , .A1( us02_n728 ) , .A2( us02_n789 ) );
  NOR2_X1 us02_U237 (.ZN( us02_n661 ) , .A2( us02_n696 ) , .A1( us02_n728 ) );
  NOR2_X1 us02_U238 (.ZN( us02_n556 ) , .A1( us02_n791 ) , .A2( us02_n813 ) );
  NOR2_X1 us02_U239 (.ZN( us02_n544 ) , .A1( us02_n748 ) , .A2( us02_n813 ) );
  NOR4_X1 us02_U24 (.A4( us02_n531 ) , .A3( us02_n532 ) , .A2( us02_n533 ) , .ZN( us02_n534 ) , .A1( us02_n819 ) );
  NOR2_X1 us02_U240 (.ZN( us02_n508 ) , .A1( us02_n728 ) , .A2( us02_n778 ) );
  NOR2_X1 us02_U241 (.A2( us02_n696 ) , .A1( us02_n779 ) , .ZN( us02_n819 ) );
  OAI22_X1 us02_U242 (.B2( us02_n749 ) , .B1( us02_n750 ) , .A1( us02_n751 ) , .ZN( us02_n755 ) , .A2( us02_n805 ) );
  NOR2_X1 us02_U243 (.ZN( us02_n750 ) , .A2( us02_n851 ) , .A1( us02_n859 ) );
  NOR3_X1 us02_U244 (.ZN( us02_n751 ) , .A2( us02_n852 ) , .A1( us02_n862 ) , .A3( us02_n864 ) );
  NOR2_X1 us02_U245 (.ZN( us02_n529 ) , .A2( us02_n743 ) , .A1( us02_n791 ) );
  NOR2_X1 us02_U246 (.A1( us02_n748 ) , .ZN( us02_n766 ) , .A2( us02_n802 ) );
  NOR2_X1 us02_U247 (.ZN( us02_n543 ) , .A2( us02_n784 ) , .A1( us02_n791 ) );
  NOR2_X1 us02_U248 (.ZN( us02_n662 ) , .A1( us02_n728 ) , .A2( us02_n784 ) );
  NOR2_X1 us02_U249 (.ZN( us02_n630 ) , .A1( us02_n723 ) , .A2( us02_n812 ) );
  NOR4_X1 us02_U25 (.ZN( us02_n455 ) , .A2( us02_n516 ) , .A1( us02_n542 ) , .A3( us02_n578 ) , .A4( us02_n614 ) );
  NOR2_X1 us02_U250 (.ZN( us02_n613 ) , .A1( us02_n761 ) , .A2( us02_n811 ) );
  OAI22_X1 us02_U251 (.B1( us02_n439 ) , .ZN( us02_n443 ) , .A2( us02_n727 ) , .A1( us02_n743 ) , .B2( us02_n748 ) );
  NOR3_X1 us02_U252 (.ZN( us02_n439 ) , .A2( us02_n835 ) , .A3( us02_n836 ) , .A1( us02_n845 ) );
  NOR2_X1 us02_U253 (.ZN( us02_n505 ) , .A2( us02_n727 ) , .A1( us02_n761 ) );
  NOR2_X1 us02_U254 (.ZN( us02_n515 ) , .A1( us02_n707 ) , .A2( us02_n743 ) );
  NOR2_X1 us02_U255 (.ZN( us02_n716 ) , .A2( us02_n743 ) , .A1( us02_n785 ) );
  NOR2_X1 us02_U256 (.ZN( us02_n553 ) , .A1( us02_n785 ) , .A2( us02_n812 ) );
  NOR2_X1 us02_U257 (.ZN( us02_n516 ) , .A1( us02_n707 ) , .A2( us02_n802 ) );
  NOR2_X1 us02_U258 (.ZN( us02_n557 ) , .A1( us02_n707 ) , .A2( us02_n815 ) );
  NOR2_X1 us02_U259 (.ZN( us02_n669 ) , .A1( us02_n789 ) , .A2( us02_n804 ) );
  NOR4_X1 us02_U26 (.A4( us02_n540 ) , .A3( us02_n541 ) , .A2( us02_n542 ) , .ZN( us02_n549 ) , .A1( us02_n687 ) );
  NOR2_X1 us02_U260 (.ZN( us02_n520 ) , .A1( us02_n789 ) , .A2( us02_n811 ) );
  NOR2_X1 us02_U261 (.ZN( us02_n629 ) , .A1( us02_n746 ) , .A2( us02_n814 ) );
  INV_X1 us02_U262 (.A( us02_n805 ) , .ZN( us02_n840 ) );
  AOI21_X1 us02_U263 (.ZN( us02_n570 ) , .B2( us02_n696 ) , .B1( us02_n805 ) , .A( us02_n811 ) );
  NOR2_X1 us02_U264 (.ZN( us02_n654 ) , .A1( us02_n789 ) , .A2( us02_n814 ) );
  INV_X1 us02_U265 (.A( us02_n762 ) , .ZN( us02_n865 ) );
  AOI21_X1 us02_U266 (.ZN( us02_n551 ) , .B1( us02_n668 ) , .A( us02_n696 ) , .B2( us02_n804 ) );
  NOR2_X1 us02_U267 (.ZN( us02_n667 ) , .A2( us02_n707 ) , .A1( us02_n789 ) );
  NOR2_X1 us02_U268 (.ZN( us02_n655 ) , .A1( us02_n746 ) , .A2( us02_n779 ) );
  NOR2_X1 us02_U269 (.ZN( us02_n541 ) , .A1( us02_n761 ) , .A2( us02_n790 ) );
  NOR2_X1 us02_U27 (.ZN( us02_n679 ) , .A2( us02_n833 ) , .A1( us02_n838 ) );
  NOR2_X1 us02_U270 (.ZN( us02_n700 ) , .A2( us02_n785 ) , .A1( us02_n816 ) );
  NOR2_X1 us02_U271 (.ZN( us02_n608 ) , .A2( us02_n723 ) , .A1( us02_n816 ) );
  NOR2_X1 us02_U272 (.A1( us02_n729 ) , .ZN( us02_n764 ) , .A2( us02_n785 ) );
  AOI21_X1 us02_U273 (.A( us02_n814 ) , .B2( us02_n815 ) , .B1( us02_n816 ) , .ZN( us02_n817 ) );
  INV_X1 us02_U274 (.A( us02_n728 ) , .ZN( us02_n867 ) );
  NOR2_X1 us02_U275 (.ZN( us02_n578 ) , .A2( us02_n707 ) , .A1( us02_n729 ) );
  NOR2_X1 us02_U276 (.ZN( us02_n532 ) , .A2( us02_n723 ) , .A1( us02_n729 ) );
  AOI21_X1 us02_U277 (.B1( us02_n624 ) , .ZN( us02_n626 ) , .A( us02_n762 ) , .B2( us02_n813 ) );
  AOI21_X1 us02_U278 (.A( us02_n811 ) , .B2( us02_n812 ) , .B1( us02_n813 ) , .ZN( us02_n818 ) );
  AOI21_X1 us02_U279 (.ZN( us02_n514 ) , .A( us02_n728 ) , .B1( us02_n749 ) , .B2( us02_n802 ) );
  AOI222_X1 us02_U28 (.ZN( us02_n468 ) , .B1( us02_n831 ) , .A1( us02_n838 ) , .C1( us02_n841 ) , .C2( us02_n850 ) , .A2( us02_n854 ) , .B2( us02_n864 ) );
  AOI21_X1 us02_U280 (.ZN( us02_n498 ) , .B1( us02_n679 ) , .A( us02_n811 ) , .B2( us02_n815 ) );
  AOI21_X1 us02_U281 (.ZN( us02_n649 ) , .A( us02_n778 ) , .B1( us02_n791 ) , .B2( us02_n804 ) );
  AOI21_X1 us02_U282 (.ZN( us02_n477 ) , .B2( us02_n696 ) , .A( us02_n748 ) , .B1( us02_n778 ) );
  NOR2_X1 us02_U283 (.ZN( us02_n581 ) , .A1( us02_n743 ) , .A2( us02_n814 ) );
  AOI21_X1 us02_U284 (.ZN( us02_n592 ) , .B1( us02_n749 ) , .A( us02_n791 ) , .B2( us02_n812 ) );
  NOR2_X1 us02_U285 (.A2( us02_n707 ) , .A1( us02_n761 ) , .ZN( us02_n793 ) );
  AOI21_X1 us02_U286 (.ZN( us02_n625 ) , .B2( us02_n668 ) , .A( us02_n789 ) , .B1( us02_n790 ) );
  NOR2_X1 us02_U287 (.ZN( us02_n519 ) , .A2( us02_n707 ) , .A1( us02_n813 ) );
  AOI21_X1 us02_U288 (.ZN( us02_n476 ) , .A( us02_n668 ) , .B1( us02_n749 ) , .B2( us02_n805 ) );
  NOR2_X1 us02_U289 (.ZN( us02_n558 ) , .A2( us02_n790 ) , .A1( us02_n802 ) );
  NOR4_X1 us02_U29 (.A1( us02_n465 ) , .ZN( us02_n466 ) , .A4( us02_n541 ) , .A2( us02_n553 ) , .A3( us02_n613 ) );
  NOR2_X1 us02_U290 (.ZN( us02_n518 ) , .A2( us02_n698 ) , .A1( us02_n815 ) );
  NOR2_X1 us02_U291 (.ZN( us02_n682 ) , .A2( us02_n698 ) , .A1( us02_n802 ) );
  NOR2_X1 us02_U292 (.ZN( us02_n652 ) , .A1( us02_n761 ) , .A2( us02_n785 ) );
  INV_X1 us02_U293 (.A( us02_n812 ) , .ZN( us02_n835 ) );
  AOI21_X1 us02_U294 (.ZN( us02_n509 ) , .B2( us02_n668 ) , .A( us02_n729 ) , .B1( us02_n814 ) );
  AOI21_X1 us02_U295 (.ZN( us02_n538 ) , .B2( us02_n811 ) , .A( us02_n813 ) , .B1( us02_n814 ) );
  AOI21_X1 us02_U296 (.ZN( us02_n539 ) , .A( us02_n762 ) , .B2( us02_n778 ) , .B1( us02_n816 ) );
  NOR2_X1 us02_U297 (.ZN( us02_n580 ) , .A1( us02_n668 ) , .A2( us02_n787 ) );
  AOI21_X1 us02_U298 (.ZN( us02_n588 ) , .B2( us02_n698 ) , .B1( us02_n814 ) , .A( us02_n816 ) );
  AOI21_X1 us02_U299 (.B1( us02_n698 ) , .ZN( us02_n699 ) , .A( us02_n731 ) , .B2( us02_n762 ) );
  NAND2_X1 us02_U3 (.A1( us02_n440 ) , .A2( us02_n463 ) , .ZN( us02_n707 ) );
  AOI221_X1 us02_U30 (.ZN( us02_n467 ) , .C2( us02_n713 ) , .B2( us02_n830 ) , .C1( us02_n844 ) , .B1( us02_n859 ) , .A( us02_n863 ) );
  AOI21_X1 us02_U300 (.ZN( us02_n590 ) , .B2( us02_n762 ) , .A( us02_n784 ) , .B1( us02_n811 ) );
  AOI21_X1 us02_U301 (.ZN( us02_n497 ) , .A( us02_n723 ) , .B2( us02_n761 ) , .B1( us02_n813 ) );
  NOR2_X1 us02_U302 (.ZN( us02_n546 ) , .A1( us02_n698 ) , .A2( us02_n743 ) );
  INV_X1 us02_U303 (.A( us02_n790 ) , .ZN( us02_n872 ) );
  INV_X1 us02_U304 (.A( us02_n811 ) , .ZN( us02_n853 ) );
  AOI21_X1 us02_U305 (.ZN( us02_n648 ) , .B1( us02_n728 ) , .B2( us02_n762 ) , .A( us02_n812 ) );
  NOR2_X1 us02_U306 (.ZN( us02_n684 ) , .A1( us02_n728 ) , .A2( us02_n815 ) );
  AOI21_X1 us02_U307 (.B1( us02_n685 ) , .ZN( us02_n686 ) , .A( us02_n727 ) , .B2( us02_n760 ) );
  AOI21_X1 us02_U308 (.ZN( us02_n568 ) , .B1( us02_n749 ) , .B2( us02_n761 ) , .A( us02_n779 ) );
  AOI21_X1 us02_U309 (.ZN( us02_n499 ) , .A( us02_n696 ) , .B1( us02_n707 ) , .B2( us02_n785 ) );
  NOR4_X1 us02_U31 (.A4( us02_n513 ) , .A3( us02_n514 ) , .A2( us02_n515 ) , .A1( us02_n516 ) , .ZN( us02_n523 ) );
  NOR2_X1 us02_U310 (.ZN( us02_n567 ) , .A1( us02_n728 ) , .A2( us02_n761 ) );
  NOR2_X1 us02_U311 (.ZN( us02_n579 ) , .A2( us02_n696 ) , .A1( us02_n790 ) );
  NOR2_X1 us02_U312 (.ZN( us02_n565 ) , .A2( us02_n696 ) , .A1( us02_n762 ) );
  AOI21_X1 us02_U313 (.ZN( us02_n513 ) , .A( us02_n778 ) , .B2( us02_n791 ) , .B1( us02_n811 ) );
  INV_X1 us02_U314 (.A( us02_n698 ) , .ZN( us02_n852 ) );
  NOR2_X1 us02_U315 (.ZN( us02_n664 ) , .A1( us02_n779 ) , .A2( us02_n812 ) );
  AOI21_X1 us02_U316 (.ZN( us02_n449 ) , .B2( us02_n791 ) , .A( us02_n802 ) , .B1( us02_n814 ) );
  NOR2_X1 us02_U317 (.ZN( us02_n631 ) , .A2( us02_n696 ) , .A1( us02_n723 ) );
  AOI21_X1 us02_U318 (.ZN( us02_n563 ) , .B1( us02_n723 ) , .A( us02_n778 ) , .B2( us02_n790 ) );
  AOI21_X1 us02_U319 (.ZN( us02_n496 ) , .A( us02_n778 ) , .B2( us02_n790 ) , .B1( us02_n803 ) );
  AOI222_X1 us02_U32 (.ZN( us02_n524 ) , .A1( us02_n833 ) , .B2( us02_n836 ) , .C1( us02_n843 ) , .C2( us02_n849 ) , .A2( us02_n851 ) , .B1( us02_n865 ) );
  NAND2_X1 us02_U320 (.ZN( us02_n752 ) , .A1( us02_n762 ) , .A2( us02_n804 ) );
  NOR2_X1 us02_U321 (.ZN( us02_n528 ) , .A1( us02_n707 ) , .A2( us02_n778 ) );
  NOR2_X1 us02_U322 (.ZN( us02_n577 ) , .A1( us02_n707 ) , .A2( us02_n812 ) );
  AOI21_X1 us02_U323 (.ZN( us02_n688 ) , .B2( us02_n748 ) , .B1( us02_n762 ) , .A( us02_n805 ) );
  NOR2_X1 us02_U324 (.ZN( us02_n566 ) , .A1( us02_n746 ) , .A2( us02_n804 ) );
  NOR2_X1 us02_U325 (.ZN( us02_n683 ) , .A1( us02_n790 ) , .A2( us02_n812 ) );
  NOR2_X1 us02_U326 (.A2( us02_n812 ) , .A1( us02_n814 ) , .ZN( us02_n820 ) );
  AOI21_X1 us02_U327 (.A( us02_n789 ) , .B2( us02_n790 ) , .B1( us02_n791 ) , .ZN( us02_n792 ) );
  AOI21_X1 us02_U328 (.A( us02_n732 ) , .ZN( us02_n733 ) , .B2( us02_n779 ) , .B1( us02_n791 ) );
  NOR2_X1 us02_U329 (.ZN( us02_n710 ) , .A1( us02_n761 ) , .A2( us02_n762 ) );
  NOR4_X1 us02_U33 (.A3( us02_n520 ) , .A1( us02_n521 ) , .ZN( us02_n522 ) , .A2( us02_n672 ) , .A4( us02_n768 ) );
  NOR2_X1 us02_U330 (.ZN( us02_n582 ) , .A1( us02_n791 ) , .A2( us02_n816 ) );
  NOR2_X1 us02_U331 (.ZN( us02_n533 ) , .A1( us02_n723 ) , .A2( us02_n787 ) );
  NOR2_X1 us02_U332 (.ZN( us02_n681 ) , .A2( us02_n707 ) , .A1( us02_n816 ) );
  INV_X1 us02_U333 (.A( us02_n696 ) , .ZN( us02_n837 ) );
  NOR2_X1 us02_U334 (.ZN( us02_n641 ) , .A2( us02_n787 ) , .A1( us02_n790 ) );
  INV_X1 us02_U335 (.A( us02_n814 ) , .ZN( us02_n854 ) );
  AOI21_X1 us02_U336 (.ZN( us02_n441 ) , .A( us02_n698 ) , .B1( us02_n732 ) , .B2( us02_n749 ) );
  INV_X1 us02_U337 (.A( us02_n779 ) , .ZN( us02_n849 ) );
  AOI22_X1 us02_U338 (.A2( us02_n781 ) , .ZN( us02_n782 ) , .B2( us02_n830 ) , .A1( us02_n833 ) , .B1( us02_n862 ) );
  NAND2_X1 us02_U339 (.ZN( us02_n670 ) , .A1( us02_n805 ) , .A2( us02_n815 ) );
  NOR4_X1 us02_U34 (.A3( us02_n754 ) , .A2( us02_n755 ) , .A1( us02_n756 ) , .ZN( us02_n757 ) , .A4( us02_n868 ) );
  NAND2_X1 us02_U340 (.ZN( us02_n713 ) , .A1( us02_n727 ) , .A2( us02_n779 ) );
  NAND2_X1 us02_U341 (.A2( us02_n761 ) , .A1( us02_n805 ) , .ZN( us02_n809 ) );
  AOI21_X1 us02_U342 (.ZN( us02_n442 ) , .B1( us02_n788 ) , .B2( us02_n790 ) , .A( us02_n813 ) );
  NOR2_X1 us02_U343 (.ZN( us02_n483 ) , .A1( us02_n787 ) , .A2( us02_n804 ) );
  NOR2_X1 us02_U344 (.ZN( us02_n469 ) , .A2( us02_n778 ) , .A1( us02_n814 ) );
  INV_X1 us02_U345 (.A( us02_n784 ) , .ZN( us02_n845 ) );
  OAI21_X1 us02_U346 (.A( us02_n786 ) , .B2( us02_n787 ) , .B1( us02_n788 ) , .ZN( us02_n794 ) );
  OAI21_X1 us02_U347 (.ZN( us02_n786 ) , .A( us02_n838 ) , .B1( us02_n862 ) , .B2( us02_n872 ) );
  NOR2_X1 us02_U348 (.ZN( us02_n711 ) , .A2( us02_n723 ) , .A1( us02_n789 ) );
  NOR2_X1 us02_U349 (.ZN( us02_n525 ) , .A1( us02_n723 ) , .A2( us02_n749 ) );
  AOI211_X1 us02_U35 (.B( us02_n744 ) , .A( us02_n745 ) , .ZN( us02_n758 ) , .C1( us02_n831 ) , .C2( us02_n852 ) );
  NAND2_X1 us02_U350 (.A1( us02_n698 ) , .A2( us02_n728 ) , .ZN( us02_n781 ) );
  AOI21_X1 us02_U351 (.ZN( us02_n638 ) , .B2( us02_n748 ) , .A( us02_n787 ) , .B1( us02_n811 ) );
  AOI21_X1 us02_U352 (.ZN( us02_n639 ) , .B2( us02_n746 ) , .A( us02_n791 ) , .B1( us02_n802 ) );
  AOI21_X1 us02_U353 (.ZN( us02_n640 ) , .B1( us02_n679 ) , .A( us02_n790 ) , .B2( us02_n816 ) );
  NOR2_X1 us02_U354 (.ZN( us02_n517 ) , .A1( us02_n707 ) , .A2( us02_n787 ) );
  OAI21_X1 us02_U355 (.A( us02_n697 ) , .ZN( us02_n701 ) , .B2( us02_n749 ) , .B1( us02_n803 ) );
  OAI21_X1 us02_U356 (.ZN( us02_n697 ) , .B2( us02_n832 ) , .B1( us02_n837 ) , .A( us02_n859 ) );
  OAI21_X1 us02_U357 (.A( us02_n730 ) , .B1( us02_n731 ) , .ZN( us02_n735 ) , .B2( us02_n804 ) );
  OAI21_X1 us02_U358 (.ZN( us02_n730 ) , .A( us02_n832 ) , .B2( us02_n851 ) , .B1( us02_n872 ) );
  NAND2_X1 us02_U359 (.A2( us02_n748 ) , .A1( us02_n785 ) , .ZN( us02_n808 ) );
  NOR3_X1 us02_U36 (.A3( us02_n740 ) , .A2( us02_n741 ) , .A1( us02_n742 ) , .ZN( us02_n759 ) );
  INV_X1 us02_U360 (.A( us02_n816 ) , .ZN( us02_n843 ) );
  INV_X1 us02_U361 (.A( us02_n723 ) , .ZN( us02_n855 ) );
  AND2_X1 us02_U362 (.ZN( us02_n731 ) , .A1( us02_n778 ) , .A2( us02_n784 ) );
  NAND2_X1 us02_U363 (.A1( us02_n446 ) , .A2( us02_n448 ) , .ZN( us02_n804 ) );
  NAND2_X1 us02_U364 (.A1( us02_n454 ) , .A2( us02_n470 ) , .ZN( us02_n802 ) );
  NAND2_X1 us02_U365 (.A1( us02_n450 ) , .A2( us02_n453 ) , .ZN( us02_n813 ) );
  NAND2_X1 us02_U366 (.A1( us02_n450 ) , .A2( us02_n470 ) , .ZN( us02_n815 ) );
  NAND2_X1 us02_U367 (.A1( us02_n453 ) , .A2( us02_n460 ) , .ZN( us02_n812 ) );
  NAND2_X1 us02_U368 (.A1( us02_n452 ) , .A2( us02_n460 ) , .ZN( us02_n743 ) );
  NAND2_X1 us02_U369 (.A1( us02_n451 ) , .A2( us02_n464 ) , .ZN( us02_n668 ) );
  NOR4_X1 us02_U37 (.A4( us02_n733 ) , .A3( us02_n734 ) , .A2( us02_n735 ) , .A1( us02_n736 ) , .ZN( us02_n737 ) );
  NAND2_X1 us02_U370 (.A2( us02_n447 ) , .A1( us02_n459 ) , .ZN( us02_n727 ) );
  NAND2_X1 us02_U371 (.A1( us02_n454 ) , .A2( us02_n461 ) , .ZN( us02_n749 ) );
  NAND2_X1 us02_U372 (.A2( us02_n452 ) , .A1( us02_n454 ) , .ZN( us02_n805 ) );
  NAND2_X1 us02_U373 (.A2( us02_n453 ) , .A1( us02_n471 ) , .ZN( us02_n778 ) );
  NAND2_X1 us02_U374 (.A1( us02_n452 ) , .A2( us02_n471 ) , .ZN( us02_n784 ) );
  NAND2_X1 us02_U375 (.A2( us02_n463 ) , .A1( us02_n464 ) , .ZN( us02_n811 ) );
  NAND2_X1 us02_U376 (.A1( us02_n440 ) , .A2( us02_n459 ) , .ZN( us02_n698 ) );
  NAND2_X1 us02_U377 (.A2( us02_n448 ) , .A1( us02_n451 ) , .ZN( us02_n762 ) );
  NAND2_X1 us02_U378 (.A2( us02_n447 ) , .A1( us02_n451 ) , .ZN( us02_n728 ) );
  NAND2_X1 us02_U379 (.A2( us02_n460 ) , .A1( us02_n461 ) , .ZN( us02_n746 ) );
  AOI211_X1 us02_U38 (.B( us02_n724 ) , .A( us02_n725 ) , .ZN( us02_n738 ) , .C1( us02_n842 ) , .C2( us02_n854 ) );
  NAND2_X2 us02_U380 (.A2( us02_n460 ) , .A1( us02_n470 ) , .ZN( us02_n696 ) );
  NAND2_X1 us02_U381 (.A1( us02_n461 ) , .A2( us02_n471 ) , .ZN( us02_n787 ) );
  NOR2_X1 us02_U382 (.ZN( us02_n464 ) , .A2( us02_n846 ) , .A1( us02_n847 ) );
  NOR2_X1 us02_U383 (.ZN( us02_n452 ) , .A1( us02_n825 ) , .A2( us02_n826 ) );
  NOR2_X1 us02_U384 (.ZN( us02_n450 ) , .A1( us02_n827 ) , .A2( us02_n828 ) );
  NOR2_X1 us02_U385 (.ZN( us02_n446 ) , .A2( us02_n848 ) , .A1( us02_n857 ) );
  NAND2_X1 us02_U386 (.A2( us02_n453 ) , .A1( us02_n454 ) , .ZN( us02_n729 ) );
  NAND2_X1 us02_U387 (.A1( us02_n450 ) , .A2( us02_n461 ) , .ZN( us02_n789 ) );
  NAND2_X2 us02_U388 (.A2( us02_n447 ) , .A1( us02_n463 ) , .ZN( us02_n814 ) );
  NAND2_X2 us02_U389 (.A2( us02_n440 ) , .A1( us02_n451 ) , .ZN( us02_n790 ) );
  NOR3_X1 us02_U39 (.A3( us02_n721 ) , .A1( us02_n722 ) , .ZN( us02_n739 ) , .A2( us02_n740 ) );
  NAND2_X2 us02_U390 (.A1( us02_n448 ) , .A2( us02_n463 ) , .ZN( us02_n723 ) );
  NAND2_X1 us02_U391 (.A2( us02_n440 ) , .A1( us02_n446 ) , .ZN( us02_n783 ) );
  NAND2_X2 us02_U392 (.A1( us02_n448 ) , .A2( us02_n459 ) , .ZN( us02_n791 ) );
  NAND2_X2 us02_U393 (.A2( us02_n459 ) , .A1( us02_n464 ) , .ZN( us02_n779 ) );
  NAND2_X1 us02_U394 (.A1( us02_n446 ) , .A2( us02_n447 ) , .ZN( us02_n785 ) );
  NOR2_X1 us02_U395 (.A2( sa02_6 ) , .A1( sa02_7 ) , .ZN( us02_n463 ) );
  NOR2_X1 us02_U396 (.A2( sa02_5 ) , .ZN( us02_n447 ) , .A1( us02_n846 ) );
  NOR2_X1 us02_U397 (.A2( sa02_7 ) , .ZN( us02_n459 ) , .A1( us02_n848 ) );
  NOR2_X1 us02_U398 (.A2( sa02_4 ) , .ZN( us02_n448 ) , .A1( us02_n847 ) );
  NOR2_X1 us02_U399 (.A2( sa02_4 ) , .A1( sa02_5 ) , .ZN( us02_n440 ) );
  NAND2_X1 us02_U4 (.A2( us02_n470 ) , .A1( us02_n471 ) , .ZN( us02_n816 ) );
  AOI221_X1 us02_U40 (.A( us02_n780 ) , .ZN( us02_n797 ) , .C2( us02_n836 ) , .B2( us02_n837 ) , .B1( us02_n864 ) , .C1( us02_n865 ) );
  NOR2_X1 us02_U400 (.A2( sa02_1 ) , .ZN( us02_n470 ) , .A1( us02_n825 ) );
  NOR2_X1 us02_U401 (.A2( sa02_2 ) , .A1( sa02_3 ) , .ZN( us02_n471 ) );
  NOR2_X1 us02_U402 (.A2( sa02_6 ) , .ZN( us02_n451 ) , .A1( us02_n857 ) );
  NOR2_X1 us02_U403 (.A2( sa02_2 ) , .ZN( us02_n460 ) , .A1( us02_n828 ) );
  NOR2_X1 us02_U404 (.A2( sa02_0 ) , .ZN( us02_n453 ) , .A1( us02_n826 ) );
  NOR2_X1 us02_U405 (.A2( sa02_0 ) , .A1( sa02_1 ) , .ZN( us02_n461 ) );
  NOR2_X1 us02_U406 (.A2( sa02_3 ) , .ZN( us02_n454 ) , .A1( us02_n827 ) );
  INV_X1 us02_U407 (.A( sa02_6 ) , .ZN( us02_n848 ) );
  INV_X1 us02_U408 (.A( sa02_1 ) , .ZN( us02_n826 ) );
  INV_X1 us02_U409 (.A( sa02_3 ) , .ZN( us02_n828 ) );
  NOR4_X1 us02_U41 (.A4( us02_n792 ) , .A3( us02_n793 ) , .A2( us02_n794 ) , .A1( us02_n795 ) , .ZN( us02_n796 ) );
  INV_X1 us02_U410 (.A( sa02_2 ) , .ZN( us02_n827 ) );
  INV_X1 us02_U411 (.A( sa02_0 ) , .ZN( us02_n825 ) );
  INV_X1 us02_U412 (.A( sa02_5 ) , .ZN( us02_n847 ) );
  INV_X1 us02_U413 (.A( sa02_7 ) , .ZN( us02_n857 ) );
  OAI221_X1 us02_U414 (.A( us02_n782 ) , .C2( us02_n783 ) , .B2( us02_n784 ) , .B1( us02_n785 ) , .ZN( us02_n795 ) , .C1( us02_n812 ) );
  OAI22_X1 us02_U415 (.ZN( us02_n587 ) , .A2( us02_n746 ) , .B2( us02_n761 ) , .A1( us02_n762 ) , .B1( us02_n783 ) );
  AOI21_X1 us02_U416 (.ZN( us02_n591 ) , .B1( us02_n727 ) , .B2( us02_n783 ) , .A( us02_n789 ) );
  OAI221_X1 us02_U417 (.A( us02_n695 ) , .ZN( us02_n702 ) , .C2( us02_n783 ) , .C1( us02_n784 ) , .B1( us02_n785 ) , .B2( us02_n805 ) );
  NAND2_X1 us02_U418 (.A1( us02_n728 ) , .A2( us02_n783 ) , .ZN( us02_n810 ) );
  AOI21_X1 us02_U419 (.ZN( us02_n622 ) , .B1( us02_n698 ) , .A( us02_n778 ) , .B2( us02_n783 ) );
  NOR4_X1 us02_U42 (.A4( us02_n775 ) , .A3( us02_n776 ) , .A1( us02_n777 ) , .ZN( us02_n798 ) , .A2( us02_n800 ) );
  OAI22_X1 us02_U420 (.ZN( us02_n680 ) , .A1( us02_n698 ) , .A2( us02_n729 ) , .B2( us02_n783 ) , .B1( us02_n816 ) );
  AOI21_X1 us02_U421 (.ZN( us02_n647 ) , .A( us02_n761 ) , .B2( us02_n783 ) , .B1( us02_n791 ) );
  OAI21_X1 us02_U422 (.A( us02_n612 ) , .ZN( us02_n615 ) , .B1( us02_n624 ) , .B2( us02_n783 ) );
  NOR2_X1 us02_U423 (.ZN( us02_n650 ) , .A1( us02_n783 ) , .A2( us02_n787 ) );
  NOR2_X1 us02_U424 (.ZN( us02_n552 ) , .A2( us02_n743 ) , .A1( us02_n783 ) );
  NOR2_X1 us02_U425 (.ZN( us02_n609 ) , .A1( us02_n783 ) , .A2( us02_n815 ) );
  OAI222_X1 us02_U426 (.A2( us02_n668 ) , .ZN( us02_n673 ) , .B1( us02_n746 ) , .B2( us02_n783 ) , .C2( us02_n787 ) , .C1( us02_n814 ) , .A1( us02_n816 ) );
  NOR2_X1 us02_U427 (.ZN( us02_n599 ) , .A2( us02_n696 ) , .A1( us02_n783 ) );
  INV_X1 us02_U428 (.A( us02_n783 ) , .ZN( us02_n860 ) );
  AOI221_X1 us02_U429 (.A( us02_n575 ) , .ZN( us02_n586 ) , .B2( us02_n830 ) , .C2( us02_n842 ) , .B1( us02_n853 ) , .C1( us02_n860 ) );
  NOR2_X1 us02_U43 (.ZN( us02_n803 ) , .A1( us02_n853 ) , .A2( us02_n860 ) );
  AOI21_X1 us02_U430 (.ZN( us02_n575 ) , .B2( us02_n723 ) , .B1( us02_n747 ) , .A( us02_n784 ) );
  INV_X1 us02_U431 (.A( sa02_4 ) , .ZN( us02_n846 ) );
  NAND2_X1 us02_U432 (.ZN( sa02_sr_2 ) , .A2( us02_n438 ) , .A1( us02_n644 ) );
  NOR3_X1 us02_U433 (.A2( us02_n606 ) , .A1( us02_n607 ) , .ZN( us02_n645 ) , .A3( us02_n721 ) );
  AOI222_X1 us02_U434 (.B2( us02_n637 ) , .ZN( us02_n643 ) , .B1( us02_n840 ) , .A1( us02_n841 ) , .C2( us02_n845 ) , .C1( us02_n862 ) , .A2( us02_n864 ) );
  NOR4_X1 us02_U435 (.A4( us02_n638 ) , .A3( us02_n639 ) , .A2( us02_n640 ) , .A1( us02_n641 ) , .ZN( us02_n642 ) );
  AOI211_X1 us02_U436 (.A( us02_n636 ) , .ZN( us02_n644 ) , .B( us02_n742 ) , .C2( us02_n838 ) , .C1( us02_n853 ) );
  NAND3_X1 us02_U437 (.ZN( sa02_sr_6 ) , .A3( us02_n796 ) , .A2( us02_n797 ) , .A1( us02_n798 ) );
  NAND3_X1 us02_U438 (.ZN( sa02_sr_5 ) , .A3( us02_n757 ) , .A2( us02_n758 ) , .A1( us02_n759 ) );
  NAND3_X1 us02_U439 (.ZN( sa02_sr_4 ) , .A3( us02_n737 ) , .A2( us02_n738 ) , .A1( us02_n739 ) );
  NAND4_X1 us02_U44 (.ZN( sa02_sr_3 ) , .A4( us02_n703 ) , .A3( us02_n704 ) , .A2( us02_n705 ) , .A1( us02_n706 ) );
  NAND3_X1 us02_U440 (.A3( us02_n674 ) , .A2( us02_n675 ) , .A1( us02_n676 ) , .ZN( us02_n806 ) );
  NAND3_X1 us02_U441 (.ZN( us02_n637 ) , .A3( us02_n707 ) , .A2( us02_n723 ) , .A1( us02_n791 ) );
  NAND3_X1 us02_U442 (.A3( us02_n617 ) , .A2( us02_n618 ) , .A1( us02_n619 ) , .ZN( us02_n724 ) );
  NAND3_X1 us02_U443 (.A3( us02_n584 ) , .A2( us02_n585 ) , .A1( us02_n586 ) , .ZN( us02_n620 ) );
  NAND3_X1 us02_U444 (.ZN( us02_n564 ) , .A3( us02_n679 ) , .A2( us02_n749 ) , .A1( us02_n784 ) );
  NAND3_X1 us02_U445 (.A3( us02_n522 ) , .A2( us02_n523 ) , .A1( us02_n524 ) , .ZN( us02_n741 ) );
  NAND3_X1 us02_U446 (.A3( us02_n511 ) , .A1( us02_n512 ) , .ZN( us02_n607 ) , .A2( us02_n870 ) );
  NAND3_X1 us02_U447 (.A3( us02_n466 ) , .A2( us02_n467 ) , .A1( us02_n468 ) , .ZN( us02_n776 ) );
  NAND4_X1 us02_U448 (.A4( us02_n632 ) , .A3( us02_n633 ) , .A2( us02_n634 ) , .A1( us02_n635 ) , .ZN( us02_n742 ) );
  NOR4_X1 us02_U45 (.A4( us02_n699 ) , .A3( us02_n700 ) , .A2( us02_n701 ) , .A1( us02_n702 ) , .ZN( us02_n703 ) );
  AOI211_X1 us02_U46 (.B( us02_n693 ) , .A( us02_n694 ) , .ZN( us02_n704 ) , .C2( us02_n830 ) , .C1( us02_n850 ) );
  NOR2_X1 us02_U47 (.ZN( us02_n706 ) , .A2( us02_n775 ) , .A1( us02_n799 ) );
  NAND4_X1 us02_U48 (.ZN( sa02_sr_7 ) , .A4( us02_n821 ) , .A3( us02_n822 ) , .A2( us02_n823 ) , .A1( us02_n824 ) );
  NOR4_X1 us02_U49 (.A4( us02_n817 ) , .A3( us02_n818 ) , .A2( us02_n819 ) , .A1( us02_n820 ) , .ZN( us02_n821 ) );
  NOR3_X1 us02_U5 (.ZN( us02_n597 ) , .A1( us02_n607 ) , .A3( us02_n722 ) , .A2( us02_n741 ) );
  AOI222_X1 us02_U50 (.C2( us02_n808 ) , .B2( us02_n809 ) , .A2( us02_n810 ) , .ZN( us02_n822 ) , .C1( us02_n831 ) , .A1( us02_n838 ) , .B1( us02_n852 ) );
  AOI211_X1 us02_U51 (.B( us02_n806 ) , .A( us02_n807 ) , .ZN( us02_n823 ) , .C1( us02_n841 ) , .C2( us02_n849 ) );
  NOR2_X1 us02_U52 (.ZN( us02_n747 ) , .A1( us02_n860 ) , .A2( us02_n861 ) );
  NAND4_X1 us02_U53 (.ZN( sa02_sr_0 ) , .A4( us02_n500 ) , .A3( us02_n501 ) , .A2( us02_n502 ) , .A1( us02_n503 ) );
  AOI221_X1 us02_U54 (.A( us02_n496 ) , .ZN( us02_n501 ) , .B2( us02_n842 ) , .C1( us02_n845 ) , .C2( us02_n859 ) , .B1( us02_n861 ) );
  NOR4_X1 us02_U55 (.A4( us02_n497 ) , .A3( us02_n498 ) , .A2( us02_n499 ) , .ZN( us02_n500 ) , .A1( us02_n526 ) );
  AOI211_X1 us02_U56 (.A( us02_n495 ) , .ZN( us02_n502 ) , .B( us02_n801 ) , .C2( us02_n838 ) , .C1( us02_n850 ) );
  NAND4_X1 us02_U57 (.ZN( sa02_sr_1 ) , .A4( us02_n594 ) , .A3( us02_n595 ) , .A2( us02_n596 ) , .A1( us02_n597 ) );
  NOR4_X1 us02_U58 (.A4( us02_n590 ) , .A3( us02_n591 ) , .A2( us02_n592 ) , .A1( us02_n593 ) , .ZN( us02_n594 ) );
  AOI211_X1 us02_U59 (.B( us02_n588 ) , .A( us02_n589 ) , .ZN( us02_n595 ) , .C2( us02_n810 ) , .C1( us02_n832 ) );
  NOR3_X1 us02_U6 (.A3( us02_n799 ) , .A2( us02_n800 ) , .A1( us02_n801 ) , .ZN( us02_n824 ) );
  AOI211_X1 us02_U60 (.A( us02_n587 ) , .ZN( us02_n596 ) , .B( us02_n620 ) , .C1( us02_n844 ) , .C2( us02_n854 ) );
  NOR2_X1 us02_U61 (.ZN( us02_n624 ) , .A2( us02_n835 ) , .A1( us02_n838 ) );
  AND3_X1 us02_U62 (.ZN( us02_n438 ) , .A2( us02_n642 ) , .A3( us02_n643 ) , .A1( us02_n645 ) );
  NOR4_X1 us02_U63 (.A4( us02_n576 ) , .A3( us02_n577 ) , .A2( us02_n578 ) , .ZN( us02_n585 ) , .A1( us02_n682 ) );
  NOR4_X1 us02_U64 (.A1( us02_n583 ) , .ZN( us02_n584 ) , .A3( us02_n651 ) , .A2( us02_n661 ) , .A4( us02_n766 ) );
  AOI211_X1 us02_U65 (.B( us02_n622 ) , .A( us02_n623 ) , .ZN( us02_n634 ) , .C2( us02_n835 ) , .C1( us02_n862 ) );
  NOR4_X1 us02_U66 (.A4( us02_n628 ) , .A3( us02_n629 ) , .A2( us02_n630 ) , .A1( us02_n631 ) , .ZN( us02_n632 ) );
  NOR4_X1 us02_U67 (.A4( us02_n625 ) , .A3( us02_n626 ) , .A2( us02_n627 ) , .ZN( us02_n633 ) , .A1( us02_n663 ) );
  NAND4_X1 us02_U68 (.A4( us02_n656 ) , .A3( us02_n657 ) , .A2( us02_n658 ) , .A1( us02_n659 ) , .ZN( us02_n799 ) );
  NOR3_X1 us02_U69 (.A3( us02_n647 ) , .A2( us02_n648 ) , .A1( us02_n649 ) , .ZN( us02_n658 ) );
  NOR3_X1 us02_U7 (.ZN( us02_n503 ) , .A2( us02_n678 ) , .A3( us02_n776 ) , .A1( us02_n875 ) );
  NOR3_X1 us02_U70 (.A3( us02_n650 ) , .A2( us02_n651 ) , .A1( us02_n652 ) , .ZN( us02_n657 ) );
  NOR3_X1 us02_U71 (.A3( us02_n653 ) , .A2( us02_n654 ) , .A1( us02_n655 ) , .ZN( us02_n656 ) );
  NAND4_X1 us02_U72 (.A4( us02_n771 ) , .A3( us02_n772 ) , .A2( us02_n773 ) , .A1( us02_n774 ) , .ZN( us02_n800 ) );
  NOR3_X1 us02_U73 (.A3( us02_n764 ) , .A2( us02_n765 ) , .A1( us02_n766 ) , .ZN( us02_n772 ) );
  NOR4_X1 us02_U74 (.A4( us02_n767 ) , .A3( us02_n768 ) , .A2( us02_n769 ) , .A1( us02_n770 ) , .ZN( us02_n771 ) );
  AOI222_X1 us02_U75 (.ZN( us02_n774 ) , .A1( us02_n829 ) , .C1( us02_n833 ) , .B2( us02_n840 ) , .A2( us02_n849 ) , .B1( us02_n860 ) , .C2( us02_n872 ) );
  NOR4_X1 us02_U76 (.A4( us02_n664 ) , .A3( us02_n665 ) , .A2( us02_n666 ) , .A1( us02_n667 ) , .ZN( us02_n675 ) );
  NOR4_X1 us02_U77 (.A4( us02_n660 ) , .A3( us02_n661 ) , .A2( us02_n662 ) , .A1( us02_n663 ) , .ZN( us02_n676 ) );
  NOR4_X1 us02_U78 (.A3( us02_n672 ) , .A1( us02_n673 ) , .ZN( us02_n674 ) , .A4( us02_n714 ) , .A2( us02_n858 ) );
  NOR2_X1 us02_U79 (.ZN( us02_n760 ) , .A1( us02_n832 ) , .A2( us02_n833 ) );
  INV_X1 us02_U8 (.A( us02_n705 ) , .ZN( us02_n875 ) );
  NAND4_X1 us02_U80 (.A4( us02_n455 ) , .A3( us02_n456 ) , .A2( us02_n457 ) , .A1( us02_n458 ) , .ZN( us02_n678 ) );
  NOR3_X1 us02_U81 (.ZN( us02_n456 ) , .A3( us02_n529 ) , .A1( us02_n554 ) , .A2( us02_n569 ) );
  AOI221_X1 us02_U82 (.A( us02_n449 ) , .ZN( us02_n458 ) , .C2( us02_n752 ) , .B1( us02_n831 ) , .C1( us02_n841 ) , .B2( us02_n860 ) );
  NOR4_X1 us02_U83 (.ZN( us02_n457 ) , .A2( us02_n508 ) , .A1( us02_n598 ) , .A4( us02_n627 ) , .A3( us02_n710 ) );
  NAND4_X1 us02_U84 (.A4( us02_n602 ) , .A3( us02_n603 ) , .A2( us02_n604 ) , .A1( us02_n605 ) , .ZN( us02_n721 ) );
  NOR3_X1 us02_U85 (.A1( us02_n598 ) , .ZN( us02_n603 ) , .A3( us02_n662 ) , .A2( us02_n769 ) );
  NOR4_X1 us02_U86 (.A3( us02_n599 ) , .A2( us02_n600 ) , .A1( us02_n601 ) , .ZN( us02_n602 ) , .A4( us02_n654 ) );
  AOI222_X1 us02_U87 (.ZN( us02_n605 ) , .A1( us02_n829 ) , .C2( us02_n836 ) , .B1( us02_n841 ) , .A2( us02_n855 ) , .B2( us02_n860 ) , .C1( us02_n867 ) );
  NAND4_X1 us02_U88 (.A4( us02_n534 ) , .A3( us02_n535 ) , .A2( us02_n536 ) , .A1( us02_n537 ) , .ZN( us02_n621 ) );
  NOR4_X1 us02_U89 (.A4( us02_n525 ) , .A2( us02_n526 ) , .A1( us02_n527 ) , .ZN( us02_n537 ) , .A3( us02_n700 ) );
  NOR3_X1 us02_U9 (.A3( us02_n620 ) , .A2( us02_n621 ) , .ZN( us02_n635 ) , .A1( us02_n724 ) );
  NOR4_X1 us02_U90 (.A1( us02_n530 ) , .ZN( us02_n535 ) , .A2( us02_n653 ) , .A4( us02_n667 ) , .A3( us02_n764 ) );
  NOR4_X1 us02_U91 (.A4( us02_n528 ) , .A3( us02_n529 ) , .ZN( us02_n536 ) , .A2( us02_n683 ) , .A1( us02_n793 ) );
  NAND4_X1 us02_U92 (.A4( us02_n547 ) , .A3( us02_n548 ) , .A2( us02_n549 ) , .A1( us02_n550 ) , .ZN( us02_n744 ) );
  NOR3_X1 us02_U93 (.ZN( us02_n548 ) , .A2( us02_n650 ) , .A1( us02_n666 ) , .A3( us02_n770 ) );
  AOI211_X1 us02_U94 (.B( us02_n538 ) , .A( us02_n539 ) , .ZN( us02_n550 ) , .C2( us02_n838 ) , .C1( us02_n850 ) );
  NOR4_X1 us02_U95 (.A4( us02_n543 ) , .A3( us02_n544 ) , .A2( us02_n545 ) , .A1( us02_n546 ) , .ZN( us02_n547 ) );
  NAND4_X1 us02_U96 (.A4( us02_n478 ) , .A3( us02_n479 ) , .A2( us02_n480 ) , .A1( us02_n481 ) , .ZN( us02_n693 ) );
  NOR3_X1 us02_U97 (.ZN( us02_n479 ) , .A2( us02_n507 ) , .A3( us02_n600 ) , .A1( us02_n609 ) );
  AOI211_X1 us02_U98 (.B( us02_n476 ) , .A( us02_n477 ) , .ZN( us02_n481 ) , .C2( us02_n832 ) , .C1( us02_n860 ) );
  NOR4_X1 us02_U99 (.ZN( us02_n480 ) , .A3( us02_n531 ) , .A4( us02_n544 ) , .A2( us02_n566 ) , .A1( us02_n716 ) );
  NOR3_X1 us21_U10 (.A3( us21_n619 ) , .A2( us21_n620 ) , .ZN( us21_n634 ) , .A1( us21_n723 ) );
  NOR4_X1 us21_U100 (.A4( us21_n524 ) , .A2( us21_n525 ) , .A1( us21_n526 ) , .ZN( us21_n536 ) , .A3( us21_n699 ) );
  NOR4_X1 us21_U101 (.A1( us21_n529 ) , .ZN( us21_n534 ) , .A2( us21_n652 ) , .A4( us21_n666 ) , .A3( us21_n763 ) );
  NOR4_X1 us21_U102 (.A4( us21_n527 ) , .A3( us21_n528 ) , .ZN( us21_n535 ) , .A2( us21_n682 ) , .A1( us21_n792 ) );
  NAND4_X1 us21_U103 (.A4( us21_n546 ) , .A3( us21_n547 ) , .A2( us21_n548 ) , .A1( us21_n549 ) , .ZN( us21_n743 ) );
  NOR3_X1 us21_U104 (.ZN( us21_n547 ) , .A2( us21_n649 ) , .A1( us21_n665 ) , .A3( us21_n769 ) );
  AOI211_X1 us21_U105 (.B( us21_n537 ) , .A( us21_n538 ) , .ZN( us21_n549 ) , .C2( us21_n837 ) , .C1( us21_n849 ) );
  NOR4_X1 us21_U106 (.A4( us21_n539 ) , .A3( us21_n540 ) , .A2( us21_n541 ) , .ZN( us21_n548 ) , .A1( us21_n686 ) );
  NAND4_X1 us21_U107 (.A4( us21_n477 ) , .A3( us21_n478 ) , .A2( us21_n479 ) , .A1( us21_n480 ) , .ZN( us21_n692 ) );
  NOR3_X1 us21_U108 (.ZN( us21_n478 ) , .A2( us21_n506 ) , .A3( us21_n599 ) , .A1( us21_n608 ) );
  AOI211_X1 us21_U109 (.B( us21_n475 ) , .A( us21_n476 ) , .ZN( us21_n480 ) , .C2( us21_n831 ) , .C1( us21_n859 ) );
  NOR2_X1 us21_U11 (.ZN( us21_n493 ) , .A1( us21_n676 ) , .A2( us21_n692 ) );
  NOR4_X1 us21_U110 (.ZN( us21_n479 ) , .A3( us21_n530 ) , .A4( us21_n543 ) , .A2( us21_n565 ) , .A1( us21_n715 ) );
  NOR4_X1 us21_U111 (.A4( us21_n607 ) , .A3( us21_n608 ) , .A2( us21_n609 ) , .A1( us21_n610 ) , .ZN( us21_n617 ) );
  NOR4_X1 us21_U112 (.ZN( us21_n618 ) , .A1( us21_n654 ) , .A3( us21_n664 ) , .A4( us21_n680 ) , .A2( us21_n764 ) );
  NOR4_X1 us21_U113 (.A4( us21_n612 ) , .A3( us21_n613 ) , .A2( us21_n614 ) , .A1( us21_n615 ) , .ZN( us21_n616 ) );
  NOR2_X1 us21_U114 (.ZN( us21_n684 ) , .A1( us21_n829 ) , .A2( us21_n830 ) );
  NAND4_X1 us21_U115 (.A4( us21_n471 ) , .A3( us21_n472 ) , .A2( us21_n473 ) , .A1( us21_n474 ) , .ZN( us21_n676 ) );
  NOR4_X1 us21_U116 (.A4( us21_n468 ) , .ZN( us21_n474 ) , .A3( us21_n554 ) , .A1( us21_n733 ) , .A2( us21_n753 ) );
  NOR4_X1 us21_U117 (.ZN( us21_n473 ) , .A1( us21_n529 ) , .A3( us21_n566 ) , .A4( us21_n598 ) , .A2( us21_n640 ) );
  NOR4_X1 us21_U118 (.ZN( us21_n472 ) , .A1( us21_n504 ) , .A3( us21_n542 ) , .A2( us21_n581 ) , .A4( us21_n714 ) );
  NAND4_X1 us21_U119 (.A4( us21_n689 ) , .A3( us21_n690 ) , .A1( us21_n691 ) , .ZN( us21_n774 ) , .A2( us21_n870 ) );
  NOR2_X1 us21_U12 (.A1( us21_n676 ) , .ZN( us21_n691 ) , .A2( us21_n805 ) );
  INV_X1 us21_U120 (.A( us21_n677 ) , .ZN( us21_n870 ) );
  AOI221_X1 us21_U121 (.A( us21_n679 ) , .ZN( us21_n690 ) , .B2( us21_n838 ) , .C1( us21_n840 ) , .C2( us21_n860 ) , .B1( us21_n863 ) );
  NOR4_X1 us21_U122 (.A4( us21_n685 ) , .A3( us21_n686 ) , .A2( us21_n687 ) , .A1( us21_n688 ) , .ZN( us21_n689 ) );
  NOR2_X1 us21_U123 (.ZN( us21_n731 ) , .A2( us21_n830 ) , .A1( us21_n843 ) );
  NAND4_X1 us21_U124 (.A4( us21_n717 ) , .A3( us21_n718 ) , .A2( us21_n719 ) , .ZN( us21_n739 ) , .A1( us21_n855 ) );
  INV_X1 us21_U125 (.A( us21_n707 ) , .ZN( us21_n855 ) );
  NOR4_X1 us21_U126 (.A4( us21_n713 ) , .A3( us21_n714 ) , .A2( us21_n715 ) , .A1( us21_n716 ) , .ZN( us21_n717 ) );
  AOI221_X1 us21_U127 (.A( us21_n708 ) , .ZN( us21_n719 ) , .C2( us21_n842 ) , .B2( us21_n843 ) , .C1( us21_n859 ) , .B1( us21_n860 ) );
  NAND4_X1 us21_U128 (.A4( us21_n571 ) , .A3( us21_n572 ) , .A1( us21_n573 ) , .ZN( us21_n721 ) , .A2( us21_n872 ) );
  NOR4_X1 us21_U129 (.A4( us21_n567 ) , .A3( us21_n568 ) , .A2( us21_n569 ) , .A1( us21_n570 ) , .ZN( us21_n571 ) );
  INV_X1 us21_U13 (.A( us21_n605 ) , .ZN( us21_n872 ) );
  AOI221_X1 us21_U130 (.A( us21_n562 ) , .C2( us21_n563 ) , .ZN( us21_n572 ) , .B2( us21_n843 ) , .B1( us21_n850 ) , .C1( us21_n851 ) );
  NOR2_X1 us21_U131 (.ZN( us21_n573 ) , .A1( us21_n620 ) , .A2( us21_n743 ) );
  NAND4_X1 us21_U132 (.A4( us21_n491 ) , .A3( us21_n492 ) , .A1( us21_n493 ) , .ZN( us21_n800 ) , .A2( us21_n865 ) );
  AOI221_X1 us21_U133 (.A( us21_n487 ) , .ZN( us21_n492 ) , .B2( us21_n834 ) , .C2( us21_n839 ) , .C1( us21_n849 ) , .B1( us21_n858 ) );
  INV_X1 us21_U134 (.A( us21_n776 ) , .ZN( us21_n865 ) );
  NOR4_X1 us21_U135 (.A2( us21_n489 ) , .A1( us21_n490 ) , .ZN( us21_n491 ) , .A3( us21_n578 ) , .A4( us21_n610 ) );
  INV_X1 us21_U136 (.A( us21_n760 ) , .ZN( us21_n828 ) );
  NOR2_X1 us21_U137 (.ZN( us21_n645 ) , .A1( us21_n852 ) , .A2( us21_n866 ) );
  INV_X1 us21_U138 (.A( us21_n461 ) , .ZN( us21_n862 ) );
  OAI21_X1 us21_U139 (.ZN( us21_n461 ) , .B1( us21_n807 ) , .A( us21_n832 ) , .B2( us21_n849 ) );
  INV_X1 us21_U14 (.A( us21_n678 ) , .ZN( us21_n838 ) );
  OR4_X1 us21_U140 (.ZN( us21_n490 ) , .A4( us21_n532 ) , .A2( us21_n545 ) , .A1( us21_n557 ) , .A3( us21_n630 ) );
  OR4_X1 us21_U141 (.A4( us21_n564 ) , .A3( us21_n565 ) , .A2( us21_n566 ) , .ZN( us21_n570 ) , .A1( us21_n663 ) );
  OR4_X1 us21_U142 (.A4( us21_n680 ) , .A3( us21_n681 ) , .A2( us21_n682 ) , .A1( us21_n683 ) , .ZN( us21_n688 ) );
  OR4_X1 us21_U143 (.ZN( us21_n464 ) , .A4( us21_n516 ) , .A3( us21_n527 ) , .A2( us21_n576 ) , .A1( us21_n710 ) );
  OR4_X1 us21_U144 (.A4( us21_n516 ) , .A2( us21_n517 ) , .A1( us21_n518 ) , .ZN( us21_n520 ) , .A3( us21_n819 ) );
  OR4_X1 us21_U145 (.A4( us21_n578 ) , .A3( us21_n579 ) , .A2( us21_n580 ) , .A1( us21_n581 ) , .ZN( us21_n582 ) );
  NAND2_X1 us21_U146 (.ZN( us21_n611 ) , .A2( us21_n835 ) , .A1( us21_n871 ) );
  OR3_X1 us21_U147 (.A3( us21_n504 ) , .A2( us21_n505 ) , .A1( us21_n506 ) , .ZN( us21_n509 ) );
  AOI221_X1 us21_U148 (.A( us21_n711 ) , .B2( us21_n712 ) , .ZN( us21_n718 ) , .C1( us21_n830 ) , .B1( us21_n837 ) , .C2( us21_n861 ) );
  OR2_X1 us21_U149 (.A2( us21_n709 ) , .A1( us21_n710 ) , .ZN( us21_n711 ) );
  NOR4_X1 us21_U15 (.A4( us21_n443 ) , .A3( us21_n444 ) , .A2( us21_n514 ) , .A1( us21_n539 ) , .ZN( us21_n704 ) );
  INV_X1 us21_U150 (.A( us21_n752 ) , .ZN( us21_n867 ) );
  OAI21_X1 us21_U151 (.B1( us21_n751 ) , .ZN( us21_n752 ) , .A( us21_n843 ) , .B2( us21_n866 ) );
  INV_X1 us21_U152 (.A( us21_n670 ) , .ZN( us21_n857 ) );
  AOI21_X1 us21_U153 (.A( us21_n668 ) , .B1( us21_n669 ) , .ZN( us21_n670 ) , .B2( us21_n854 ) );
  AOI222_X1 us21_U154 (.ZN( us21_n658 ) , .A2( us21_n837 ) , .B1( us21_n839 ) , .C2( us21_n843 ) , .A1( us21_n858 ) , .C1( us21_n861 ) , .B2( us21_n868 ) );
  INV_X1 us21_U155 (.A( us21_n645 ) , .ZN( us21_n868 ) );
  OAI22_X1 us21_U156 (.ZN( us21_n481 ) , .A1( us21_n706 ) , .B2( us21_n783 ) , .A2( us21_n804 ) , .B1( us21_n810 ) );
  OAI22_X1 us21_U157 (.ZN( us21_n635 ) , .A1( us21_n697 ) , .B2( us21_n726 ) , .A2( us21_n760 ) , .B1( us21_n814 ) );
  OAI222_X1 us21_U158 (.B2( us21_n706 ) , .ZN( us21_n707 ) , .C2( us21_n722 ) , .B1( us21_n745 ) , .A1( us21_n804 ) , .C1( us21_n812 ) , .A2( us21_n813 ) );
  NAND2_X1 us21_U159 (.A1( us21_n445 ) , .A2( us21_n463 ) , .ZN( us21_n747 ) );
  OR3_X1 us21_U16 (.ZN( us21_n444 ) , .A1( us21_n526 ) , .A3( us21_n575 ) , .A2( us21_n873 ) );
  AOI22_X1 us21_U160 (.ZN( us21_n694 ) , .A1( us21_n828 ) , .B2( us21_n841 ) , .A2( us21_n863 ) , .B1( us21_n866 ) );
  INV_X1 us21_U161 (.A( us21_n728 ) , .ZN( us21_n837 ) );
  NAND2_X1 us21_U162 (.A1( us21_n449 ) , .A2( us21_n451 ) , .ZN( us21_n760 ) );
  INV_X1 us21_U163 (.A( us21_n788 ) , .ZN( us21_n830 ) );
  OAI221_X1 us21_U164 (.A( us21_n725 ) , .C2( us21_n726 ) , .B2( us21_n727 ) , .B1( us21_n728 ) , .ZN( us21_n735 ) , .C1( us21_n815 ) );
  AOI22_X1 us21_U165 (.ZN( us21_n725 ) , .B1( us21_n830 ) , .A2( us21_n836 ) , .A1( us21_n861 ) , .B2( us21_n864 ) );
  AND2_X1 us21_U166 (.ZN( us21_n746 ) , .A1( us21_n782 ) , .A2( us21_n784 ) );
  OAI22_X1 us21_U167 (.ZN( us21_n487 ) , .A1( us21_n722 ) , .B2( us21_n726 ) , .B1( us21_n728 ) , .A2( us21_n777 ) );
  OAI22_X1 us21_U168 (.ZN( us21_n622 ) , .B1( us21_n667 ) , .B2( us21_n745 ) , .A1( us21_n813 ) , .A2( us21_n814 ) );
  OAI22_X1 us21_U169 (.B2( us21_n777 ) , .B1( us21_n778 ) , .ZN( us21_n779 ) , .A2( us21_n812 ) , .A1( us21_n813 ) );
  OR4_X1 us21_U17 (.A4( us21_n440 ) , .A2( us21_n441 ) , .A1( us21_n442 ) , .ZN( us21_n443 ) , .A3( us21_n551 ) );
  OAI22_X1 us21_U170 (.A1( us21_n722 ) , .ZN( us21_n724 ) , .B2( us21_n748 ) , .B1( us21_n810 ) , .A2( us21_n814 ) );
  OAI22_X1 us21_U171 (.B2( us21_n742 ) , .ZN( us21_n744 ) , .A2( us21_n760 ) , .B1( us21_n778 ) , .A1( us21_n790 ) );
  OAI22_X1 us21_U172 (.B2( us21_n801 ) , .B1( us21_n802 ) , .A2( us21_n803 ) , .A1( us21_n804 ) , .ZN( us21_n806 ) );
  OAI22_X1 us21_U173 (.ZN( us21_n494 ) , .A2( us21_n742 ) , .A1( us21_n778 ) , .B1( us21_n789 ) , .B2( us21_n804 ) );
  INV_X1 us21_U174 (.A( us21_n742 ) , .ZN( us21_n835 ) );
  INV_X1 us21_U175 (.A( us21_n786 ) , .ZN( us21_n843 ) );
  INV_X1 us21_U176 (.A( us21_n814 ) , .ZN( us21_n829 ) );
  OAI22_X1 us21_U177 (.B1( us21_n488 ) , .ZN( us21_n489 ) , .A1( us21_n684 ) , .A2( us21_n761 ) , .B2( us21_n815 ) );
  NOR3_X1 us21_U178 (.ZN( us21_n488 ) , .A1( us21_n780 ) , .A2( us21_n848 ) , .A3( us21_n861 ) );
  OAI22_X1 us21_U179 (.ZN( us21_n588 ) , .B1( us21_n728 ) , .B2( us21_n747 ) , .A2( us21_n784 ) , .A1( us21_n801 ) );
  INV_X1 us21_U18 (.A( us21_n611 ) , .ZN( us21_n873 ) );
  OAI22_X1 us21_U180 (.ZN( us21_n693 ) , .A2( us21_n728 ) , .A1( us21_n778 ) , .B1( us21_n789 ) , .B2( us21_n815 ) );
  OAI22_X1 us21_U181 (.ZN( us21_n708 ) , .A2( us21_n726 ) , .B2( us21_n727 ) , .A1( us21_n742 ) , .B1( us21_n811 ) );
  INV_X1 us21_U182 (.A( us21_n812 ) , .ZN( us21_n831 ) );
  INV_X1 us21_U183 (.A( us21_n667 ) , .ZN( us21_n863 ) );
  NOR2_X1 us21_U184 (.ZN( us21_n716 ) , .A2( us21_n722 ) , .A1( us21_n742 ) );
  NOR2_X1 us21_U185 (.ZN( us21_n664 ) , .A1( us21_n726 ) , .A2( us21_n801 ) );
  NOR2_X1 us21_U186 (.ZN( us21_n568 ) , .A1( us21_n726 ) , .A2( us21_n804 ) );
  NOR2_X1 us21_U187 (.ZN( us21_n544 ) , .A2( us21_n778 ) , .A1( us21_n812 ) );
  INV_X1 us21_U188 (.A( us21_n748 ) , .ZN( us21_n840 ) );
  NOR2_X1 us21_U189 (.ZN( us21_n530 ) , .A2( us21_n747 ) , .A1( us21_n748 ) );
  INV_X1 us21_U19 (.A( us21_n747 ) , .ZN( us21_n861 ) );
  NOR2_X1 us21_U190 (.ZN( us21_n575 ) , .A2( us21_n697 ) , .A1( us21_n812 ) );
  NOR2_X1 us21_U191 (.ZN( us21_n652 ) , .A1( us21_n726 ) , .A2( us21_n811 ) );
  NOR2_X1 us21_U192 (.ZN( us21_n613 ) , .A1( us21_n783 ) , .A2( us21_n813 ) );
  NOR2_X1 us21_U193 (.ZN( us21_n627 ) , .A2( us21_n726 ) , .A1( us21_n783 ) );
  NOR2_X1 us21_U194 (.ZN( us21_n599 ) , .A2( us21_n778 ) , .A1( us21_n801 ) );
  NOR2_X1 us21_U195 (.ZN( us21_n610 ) , .A1( us21_n777 ) , .A2( us21_n784 ) );
  NOR2_X1 us21_U196 (.ZN( us21_n526 ) , .A2( us21_n722 ) , .A1( us21_n801 ) );
  NOR2_X1 us21_U197 (.ZN( us21_n626 ) , .A2( us21_n667 ) , .A1( us21_n783 ) );
  INV_X1 us21_U198 (.A( us21_n790 ) , .ZN( us21_n849 ) );
  NOR2_X1 us21_U199 (.A2( us21_n742 ) , .ZN( us21_n767 ) , .A1( us21_n810 ) );
  AOI222_X1 us21_U20 (.ZN( us21_n561 ) , .B1( us21_n828 ) , .C1( us21_n839 ) , .A2( us21_n841 ) , .A1( us21_n852 ) , .B2( us21_n861 ) , .C2( us21_n871 ) );
  NOR2_X1 us21_U200 (.ZN( us21_n529 ) , .A2( us21_n778 ) , .A1( us21_n814 ) );
  NOR2_X1 us21_U201 (.A2( us21_n706 ) , .A1( us21_n748 ) , .ZN( us21_n769 ) );
  NOR2_X1 us21_U202 (.ZN( us21_n597 ) , .A2( us21_n789 ) , .A1( us21_n814 ) );
  NOR2_X1 us21_U203 (.ZN( us21_n609 ) , .A2( us21_n778 ) , .A1( us21_n804 ) );
  NOR2_X1 us21_U204 (.ZN( us21_n650 ) , .A1( us21_n667 ) , .A2( us21_n812 ) );
  INV_X1 us21_U205 (.A( us21_n745 ) , .ZN( us21_n832 ) );
  NOR2_X1 us21_U206 (.A1( us21_n667 ) , .ZN( us21_n671 ) , .A2( us21_n742 ) );
  NOR2_X1 us21_U207 (.ZN( us21_n600 ) , .A1( us21_n667 ) , .A2( us21_n801 ) );
  NOR2_X1 us21_U208 (.A1( us21_n667 ) , .ZN( us21_n686 ) , .A2( us21_n814 ) );
  NOR2_X1 us21_U209 (.ZN( us21_n665 ) , .A1( us21_n748 ) , .A2( us21_n813 ) );
  NOR4_X1 us21_U21 (.ZN( us21_n471 ) , .A2( us21_n519 ) , .A4( us21_n592 ) , .A1( us21_n607 ) , .A3( us21_n627 ) );
  NOR2_X1 us21_U210 (.ZN( us21_n553 ) , .A1( us21_n748 ) , .A2( us21_n789 ) );
  NOR2_X1 us21_U211 (.ZN( us21_n506 ) , .A2( us21_n778 ) , .A1( us21_n783 ) );
  NOR2_X1 us21_U212 (.ZN( us21_n541 ) , .A2( us21_n706 ) , .A1( us21_n783 ) );
  NOR2_X1 us21_U213 (.ZN( us21_n662 ) , .A1( us21_n783 ) , .A2( us21_n789 ) );
  NOR2_X1 us21_U214 (.A1( us21_n667 ) , .ZN( us21_n764 ) , .A2( us21_n811 ) );
  NOR2_X1 us21_U215 (.A1( us21_n697 ) , .ZN( us21_n766 ) , .A2( us21_n811 ) );
  OAI22_X1 us21_U216 (.B1( us21_n438 ) , .ZN( us21_n442 ) , .A2( us21_n726 ) , .A1( us21_n742 ) , .B2( us21_n747 ) );
  NOR3_X1 us21_U217 (.ZN( us21_n438 ) , .A2( us21_n834 ) , .A3( us21_n835 ) , .A1( us21_n844 ) );
  NOR2_X1 us21_U218 (.ZN( us21_n525 ) , .A1( us21_n667 ) , .A2( us21_n777 ) );
  NOR2_X1 us21_U219 (.ZN( us21_n505 ) , .A1( us21_n810 ) , .A2( us21_n815 ) );
  NOR4_X1 us21_U22 (.A4( us21_n542 ) , .A3( us21_n543 ) , .A2( us21_n544 ) , .A1( us21_n545 ) , .ZN( us21_n546 ) );
  NOR2_X1 us21_U220 (.ZN( us21_n659 ) , .A1( us21_n727 ) , .A2( us21_n788 ) );
  INV_X1 us21_U221 (.A( us21_n801 ) , .ZN( us21_n841 ) );
  NOR2_X1 us21_U222 (.ZN( us21_n555 ) , .A1( us21_n790 ) , .A2( us21_n812 ) );
  NOR2_X1 us21_U223 (.ZN( us21_n543 ) , .A1( us21_n747 ) , .A2( us21_n812 ) );
  NOR2_X1 us21_U224 (.ZN( us21_n507 ) , .A1( us21_n727 ) , .A2( us21_n777 ) );
  NOR2_X1 us21_U225 (.ZN( us21_n528 ) , .A2( us21_n742 ) , .A1( us21_n790 ) );
  NOR2_X1 us21_U226 (.A1( us21_n747 ) , .ZN( us21_n765 ) , .A2( us21_n801 ) );
  NOR2_X1 us21_U227 (.A2( us21_n742 ) , .ZN( us21_n753 ) , .A1( us21_n803 ) );
  OAI22_X1 us21_U228 (.B2( us21_n748 ) , .B1( us21_n749 ) , .A1( us21_n750 ) , .ZN( us21_n754 ) , .A2( us21_n804 ) );
  NOR2_X1 us21_U229 (.ZN( us21_n749 ) , .A2( us21_n850 ) , .A1( us21_n858 ) );
  NOR4_X1 us21_U23 (.ZN( us21_n477 ) , .A1( us21_n518 ) , .A4( us21_n555 ) , .A3( us21_n580 ) , .A2( us21_n628 ) );
  NOR3_X1 us21_U230 (.ZN( us21_n750 ) , .A2( us21_n851 ) , .A1( us21_n861 ) , .A3( us21_n863 ) );
  NOR2_X1 us21_U231 (.ZN( us21_n542 ) , .A2( us21_n783 ) , .A1( us21_n790 ) );
  INV_X1 us21_U232 (.A( us21_n804 ) , .ZN( us21_n839 ) );
  NOR2_X1 us21_U233 (.ZN( us21_n629 ) , .A1( us21_n722 ) , .A2( us21_n811 ) );
  NOR2_X1 us21_U234 (.ZN( us21_n733 ) , .A2( us21_n801 ) , .A1( us21_n803 ) );
  NOR2_X1 us21_U235 (.ZN( us21_n514 ) , .A1( us21_n706 ) , .A2( us21_n742 ) );
  NOR2_X1 us21_U236 (.ZN( us21_n661 ) , .A1( us21_n727 ) , .A2( us21_n783 ) );
  NOR2_X1 us21_U237 (.ZN( us21_n715 ) , .A2( us21_n742 ) , .A1( us21_n784 ) );
  NOR2_X1 us21_U238 (.ZN( us21_n612 ) , .A1( us21_n760 ) , .A2( us21_n810 ) );
  INV_X1 us21_U239 (.A( us21_n726 ) , .ZN( us21_n850 ) );
  NOR4_X1 us21_U24 (.ZN( us21_n454 ) , .A2( us21_n515 ) , .A1( us21_n541 ) , .A3( us21_n577 ) , .A4( us21_n613 ) );
  NOR2_X1 us21_U240 (.ZN( us21_n552 ) , .A1( us21_n784 ) , .A2( us21_n811 ) );
  NOR2_X1 us21_U241 (.ZN( us21_n515 ) , .A1( us21_n706 ) , .A2( us21_n801 ) );
  NOR2_X1 us21_U242 (.ZN( us21_n504 ) , .A2( us21_n726 ) , .A1( us21_n760 ) );
  NOR2_X1 us21_U243 (.ZN( us21_n556 ) , .A1( us21_n706 ) , .A2( us21_n814 ) );
  NOR2_X1 us21_U244 (.ZN( us21_n519 ) , .A1( us21_n788 ) , .A2( us21_n810 ) );
  INV_X1 us21_U245 (.A( us21_n803 ) , .ZN( us21_n858 ) );
  NOR2_X1 us21_U246 (.ZN( us21_n713 ) , .A1( us21_n803 ) , .A2( us21_n815 ) );
  NOR2_X1 us21_U247 (.ZN( us21_n653 ) , .A1( us21_n788 ) , .A2( us21_n813 ) );
  NOR2_X1 us21_U248 (.ZN( us21_n666 ) , .A2( us21_n706 ) , .A1( us21_n788 ) );
  NOR2_X1 us21_U249 (.ZN( us21_n628 ) , .A1( us21_n745 ) , .A2( us21_n813 ) );
  NOR4_X1 us21_U25 (.A4( us21_n530 ) , .A3( us21_n531 ) , .A2( us21_n532 ) , .ZN( us21_n533 ) , .A1( us21_n818 ) );
  NOR2_X1 us21_U250 (.ZN( us21_n554 ) , .A1( us21_n760 ) , .A2( us21_n803 ) );
  NOR2_X1 us21_U251 (.ZN( us21_n540 ) , .A1( us21_n760 ) , .A2( us21_n789 ) );
  NOR2_X1 us21_U252 (.ZN( us21_n699 ) , .A2( us21_n784 ) , .A1( us21_n815 ) );
  NOR2_X1 us21_U253 (.A1( us21_n728 ) , .ZN( us21_n763 ) , .A2( us21_n784 ) );
  NOR2_X1 us21_U254 (.ZN( us21_n607 ) , .A2( us21_n722 ) , .A1( us21_n815 ) );
  NOR2_X1 us21_U255 (.ZN( us21_n577 ) , .A2( us21_n706 ) , .A1( us21_n728 ) );
  NOR2_X1 us21_U256 (.ZN( us21_n531 ) , .A2( us21_n722 ) , .A1( us21_n728 ) );
  AOI21_X1 us21_U257 (.A( us21_n810 ) , .B2( us21_n811 ) , .B1( us21_n812 ) , .ZN( us21_n817 ) );
  AOI21_X1 us21_U258 (.ZN( us21_n513 ) , .A( us21_n727 ) , .B1( us21_n748 ) , .B2( us21_n801 ) );
  NOR2_X1 us21_U259 (.ZN( us21_n654 ) , .A1( us21_n745 ) , .A2( us21_n778 ) );
  NOR2_X1 us21_U26 (.ZN( us21_n678 ) , .A2( us21_n832 ) , .A1( us21_n837 ) );
  AOI21_X1 us21_U260 (.A( us21_n813 ) , .B2( us21_n814 ) , .B1( us21_n815 ) , .ZN( us21_n816 ) );
  NOR2_X1 us21_U261 (.ZN( us21_n580 ) , .A1( us21_n742 ) , .A2( us21_n813 ) );
  AOI21_X1 us21_U262 (.ZN( us21_n591 ) , .B1( us21_n748 ) , .A( us21_n790 ) , .B2( us21_n811 ) );
  AOI21_X1 us21_U263 (.B1( us21_n623 ) , .ZN( us21_n625 ) , .A( us21_n761 ) , .B2( us21_n812 ) );
  NOR2_X1 us21_U264 (.A2( us21_n706 ) , .A1( us21_n760 ) , .ZN( us21_n792 ) );
  NOR2_X1 us21_U265 (.ZN( us21_n640 ) , .A2( us21_n786 ) , .A1( us21_n789 ) );
  AOI21_X1 us21_U266 (.ZN( us21_n497 ) , .B1( us21_n678 ) , .A( us21_n810 ) , .B2( us21_n814 ) );
  NOR2_X1 us21_U267 (.ZN( us21_n668 ) , .A1( us21_n788 ) , .A2( us21_n803 ) );
  NOR2_X1 us21_U268 (.ZN( us21_n557 ) , .A2( us21_n789 ) , .A1( us21_n801 ) );
  AOI21_X1 us21_U269 (.ZN( us21_n624 ) , .B2( us21_n667 ) , .A( us21_n788 ) , .B1( us21_n789 ) );
  NOR4_X1 us21_U27 (.A4( us21_n575 ) , .A3( us21_n576 ) , .A2( us21_n577 ) , .ZN( us21_n584 ) , .A1( us21_n681 ) );
  NOR2_X1 us21_U270 (.ZN( us21_n681 ) , .A2( us21_n697 ) , .A1( us21_n801 ) );
  NOR2_X1 us21_U271 (.ZN( us21_n651 ) , .A1( us21_n760 ) , .A2( us21_n784 ) );
  NOR2_X1 us21_U272 (.ZN( us21_n518 ) , .A2( us21_n706 ) , .A1( us21_n812 ) );
  INV_X1 us21_U273 (.A( us21_n811 ) , .ZN( us21_n834 ) );
  NOR2_X1 us21_U274 (.ZN( us21_n517 ) , .A2( us21_n697 ) , .A1( us21_n814 ) );
  AOI21_X1 us21_U275 (.ZN( us21_n475 ) , .A( us21_n667 ) , .B1( us21_n748 ) , .B2( us21_n804 ) );
  AOI21_X1 us21_U276 (.ZN( us21_n508 ) , .B2( us21_n667 ) , .A( us21_n728 ) , .B1( us21_n813 ) );
  AOI21_X1 us21_U277 (.ZN( us21_n537 ) , .B2( us21_n810 ) , .A( us21_n812 ) , .B1( us21_n813 ) );
  INV_X1 us21_U278 (.A( us21_n761 ) , .ZN( us21_n864 ) );
  AOI21_X1 us21_U279 (.ZN( us21_n538 ) , .A( us21_n761 ) , .B2( us21_n777 ) , .B1( us21_n815 ) );
  NOR4_X1 us21_U28 (.A1( us21_n582 ) , .ZN( us21_n583 ) , .A3( us21_n650 ) , .A2( us21_n660 ) , .A4( us21_n765 ) );
  NOR2_X1 us21_U280 (.ZN( us21_n579 ) , .A1( us21_n667 ) , .A2( us21_n786 ) );
  AOI21_X1 us21_U281 (.ZN( us21_n587 ) , .B2( us21_n697 ) , .B1( us21_n813 ) , .A( us21_n815 ) );
  AOI21_X1 us21_U282 (.ZN( us21_n589 ) , .B2( us21_n761 ) , .A( us21_n783 ) , .B1( us21_n810 ) );
  AOI21_X1 us21_U283 (.B1( us21_n697 ) , .ZN( us21_n698 ) , .A( us21_n730 ) , .B2( us21_n761 ) );
  AOI21_X1 us21_U284 (.ZN( us21_n638 ) , .B2( us21_n745 ) , .A( us21_n790 ) , .B1( us21_n801 ) );
  AOI21_X1 us21_U285 (.ZN( us21_n496 ) , .A( us21_n722 ) , .B2( us21_n760 ) , .B1( us21_n812 ) );
  INV_X1 us21_U286 (.A( us21_n789 ) , .ZN( us21_n871 ) );
  NOR2_X1 us21_U287 (.ZN( us21_n545 ) , .A1( us21_n697 ) , .A2( us21_n742 ) );
  INV_X1 us21_U288 (.A( us21_n727 ) , .ZN( us21_n866 ) );
  AOI21_X1 us21_U289 (.ZN( us21_n647 ) , .B1( us21_n727 ) , .B2( us21_n761 ) , .A( us21_n811 ) );
  AOI221_X1 us21_U29 (.A( us21_n779 ) , .ZN( us21_n796 ) , .C2( us21_n835 ) , .B2( us21_n836 ) , .B1( us21_n863 ) , .C1( us21_n864 ) );
  AOI21_X1 us21_U290 (.ZN( us21_n567 ) , .B1( us21_n748 ) , .B2( us21_n760 ) , .A( us21_n778 ) );
  INV_X1 us21_U291 (.A( us21_n810 ) , .ZN( us21_n852 ) );
  NOR2_X1 us21_U292 (.ZN( us21_n683 ) , .A1( us21_n727 ) , .A2( us21_n814 ) );
  AOI21_X1 us21_U293 (.B1( us21_n684 ) , .ZN( us21_n685 ) , .A( us21_n726 ) , .B2( us21_n759 ) );
  NOR2_X1 us21_U294 (.ZN( us21_n566 ) , .A1( us21_n727 ) , .A2( us21_n760 ) );
  NOR2_X1 us21_U295 (.ZN( us21_n663 ) , .A1( us21_n778 ) , .A2( us21_n811 ) );
  AOI21_X1 us21_U296 (.ZN( us21_n448 ) , .B2( us21_n790 ) , .A( us21_n801 ) , .B1( us21_n813 ) );
  AOI21_X1 us21_U297 (.ZN( us21_n512 ) , .A( us21_n777 ) , .B2( us21_n790 ) , .B1( us21_n810 ) );
  AOI21_X1 us21_U298 (.ZN( us21_n637 ) , .B2( us21_n747 ) , .A( us21_n786 ) , .B1( us21_n810 ) );
  INV_X1 us21_U299 (.A( us21_n697 ) , .ZN( us21_n851 ) );
  NAND2_X2 us21_U3 (.A2( us21_n458 ) , .A1( us21_n463 ) , .ZN( us21_n778 ) );
  NOR4_X1 us21_U30 (.A4( us21_n791 ) , .A3( us21_n792 ) , .A2( us21_n793 ) , .A1( us21_n794 ) , .ZN( us21_n795 ) );
  AOI21_X1 us21_U300 (.ZN( us21_n562 ) , .B1( us21_n722 ) , .A( us21_n777 ) , .B2( us21_n789 ) );
  NOR2_X1 us21_U301 (.ZN( us21_n576 ) , .A1( us21_n706 ) , .A2( us21_n811 ) );
  NOR2_X1 us21_U302 (.ZN( us21_n527 ) , .A1( us21_n706 ) , .A2( us21_n777 ) );
  AOI21_X1 us21_U303 (.ZN( us21_n687 ) , .B2( us21_n747 ) , .B1( us21_n761 ) , .A( us21_n804 ) );
  NOR2_X1 us21_U304 (.ZN( us21_n682 ) , .A1( us21_n789 ) , .A2( us21_n811 ) );
  AOI21_X1 us21_U305 (.ZN( us21_n648 ) , .A( us21_n777 ) , .B1( us21_n790 ) , .B2( us21_n803 ) );
  NOR2_X1 us21_U306 (.A2( us21_n811 ) , .A1( us21_n813 ) , .ZN( us21_n819 ) );
  AOI21_X1 us21_U307 (.A( us21_n788 ) , .B2( us21_n789 ) , .B1( us21_n790 ) , .ZN( us21_n791 ) );
  AOI21_X1 us21_U308 (.A( us21_n731 ) , .ZN( us21_n732 ) , .B2( us21_n778 ) , .B1( us21_n790 ) );
  NOR2_X1 us21_U309 (.ZN( us21_n581 ) , .A1( us21_n790 ) , .A2( us21_n815 ) );
  NOR4_X1 us21_U31 (.A4( us21_n774 ) , .A3( us21_n775 ) , .A1( us21_n776 ) , .ZN( us21_n797 ) , .A2( us21_n799 ) );
  NOR2_X1 us21_U310 (.ZN( us21_n532 ) , .A1( us21_n722 ) , .A2( us21_n786 ) );
  AOI21_X1 us21_U311 (.ZN( us21_n639 ) , .B1( us21_n678 ) , .A( us21_n789 ) , .B2( us21_n815 ) );
  NOR2_X1 us21_U312 (.ZN( us21_n709 ) , .A1( us21_n760 ) , .A2( us21_n761 ) );
  NOR2_X1 us21_U313 (.ZN( us21_n565 ) , .A1( us21_n745 ) , .A2( us21_n803 ) );
  NOR2_X1 us21_U314 (.ZN( us21_n680 ) , .A2( us21_n706 ) , .A1( us21_n815 ) );
  INV_X1 us21_U315 (.A( us21_n813 ) , .ZN( us21_n853 ) );
  AOI21_X1 us21_U316 (.ZN( us21_n440 ) , .A( us21_n697 ) , .B1( us21_n731 ) , .B2( us21_n748 ) );
  INV_X1 us21_U317 (.A( us21_n778 ) , .ZN( us21_n848 ) );
  AOI22_X1 us21_U318 (.A2( us21_n780 ) , .ZN( us21_n781 ) , .B2( us21_n829 ) , .A1( us21_n832 ) , .B1( us21_n861 ) );
  NAND2_X1 us21_U319 (.ZN( us21_n712 ) , .A1( us21_n726 ) , .A2( us21_n778 ) );
  NOR4_X1 us21_U32 (.A3( us21_n753 ) , .A2( us21_n754 ) , .A1( us21_n755 ) , .ZN( us21_n756 ) , .A4( us21_n867 ) );
  NAND2_X1 us21_U320 (.ZN( us21_n751 ) , .A1( us21_n761 ) , .A2( us21_n803 ) );
  AOI21_X1 us21_U321 (.ZN( us21_n441 ) , .B1( us21_n787 ) , .B2( us21_n789 ) , .A( us21_n812 ) );
  INV_X1 us21_U322 (.A( us21_n783 ) , .ZN( us21_n844 ) );
  AOI21_X1 us21_U323 (.ZN( us21_n495 ) , .A( us21_n777 ) , .B2( us21_n789 ) , .B1( us21_n802 ) );
  NAND2_X1 us21_U324 (.A2( us21_n760 ) , .A1( us21_n804 ) , .ZN( us21_n808 ) );
  NOR2_X1 us21_U325 (.ZN( us21_n468 ) , .A2( us21_n777 ) , .A1( us21_n813 ) );
  NOR2_X1 us21_U326 (.ZN( us21_n710 ) , .A2( us21_n722 ) , .A1( us21_n788 ) );
  NOR2_X1 us21_U327 (.ZN( us21_n482 ) , .A1( us21_n786 ) , .A2( us21_n803 ) );
  NOR2_X1 us21_U328 (.ZN( us21_n524 ) , .A1( us21_n722 ) , .A2( us21_n748 ) );
  OAI21_X1 us21_U329 (.A( us21_n729 ) , .B1( us21_n730 ) , .ZN( us21_n734 ) , .B2( us21_n803 ) );
  AOI211_X1 us21_U33 (.B( us21_n743 ) , .A( us21_n744 ) , .ZN( us21_n757 ) , .C1( us21_n830 ) , .C2( us21_n851 ) );
  OAI21_X1 us21_U330 (.ZN( us21_n729 ) , .A( us21_n831 ) , .B2( us21_n850 ) , .B1( us21_n871 ) );
  OAI21_X1 us21_U331 (.A( us21_n785 ) , .B2( us21_n786 ) , .B1( us21_n787 ) , .ZN( us21_n793 ) );
  OAI21_X1 us21_U332 (.ZN( us21_n785 ) , .A( us21_n837 ) , .B1( us21_n861 ) , .B2( us21_n871 ) );
  NAND2_X1 us21_U333 (.A1( us21_n697 ) , .A2( us21_n727 ) , .ZN( us21_n780 ) );
  NOR2_X1 us21_U334 (.ZN( us21_n516 ) , .A1( us21_n706 ) , .A2( us21_n786 ) );
  NAND2_X1 us21_U335 (.ZN( us21_n669 ) , .A1( us21_n804 ) , .A2( us21_n814 ) );
  OAI21_X1 us21_U336 (.A( us21_n696 ) , .ZN( us21_n700 ) , .B2( us21_n748 ) , .B1( us21_n802 ) );
  OAI21_X1 us21_U337 (.ZN( us21_n696 ) , .B2( us21_n831 ) , .B1( us21_n836 ) , .A( us21_n858 ) );
  NAND2_X1 us21_U338 (.A2( us21_n747 ) , .A1( us21_n784 ) , .ZN( us21_n807 ) );
  INV_X1 us21_U339 (.A( us21_n722 ) , .ZN( us21_n854 ) );
  NOR3_X1 us21_U34 (.A3( us21_n739 ) , .A2( us21_n740 ) , .A1( us21_n741 ) , .ZN( us21_n758 ) );
  INV_X1 us21_U340 (.A( us21_n815 ) , .ZN( us21_n842 ) );
  AND2_X1 us21_U341 (.ZN( us21_n730 ) , .A1( us21_n777 ) , .A2( us21_n783 ) );
  OAI222_X1 us21_U342 (.ZN( us21_n615 ) , .B1( us21_n695 ) , .C1( us21_n722 ) , .C2( us21_n745 ) , .B2( us21_n784 ) , .A2( us21_n790 ) , .A1( us21_n814 ) );
  AOI221_X1 us21_U343 (.A( us21_n762 ) , .ZN( us21_n772 ) , .C2( us21_n808 ) , .B2( us21_n833 ) , .C1( us21_n853 ) , .B1( us21_n864 ) );
  AOI21_X1 us21_U344 (.B2( us21_n761 ) , .ZN( us21_n762 ) , .A( us21_n786 ) , .B1( us21_n790 ) );
  INV_X1 us21_U345 (.A( us21_n759 ) , .ZN( us21_n833 ) );
  NAND2_X2 us21_U346 (.A2( us21_n439 ) , .A1( us21_n445 ) , .ZN( us21_n782 ) );
  NAND2_X1 us21_U347 (.A1( us21_n453 ) , .A2( us21_n469 ) , .ZN( us21_n801 ) );
  NAND2_X1 us21_U348 (.A1( us21_n452 ) , .A2( us21_n459 ) , .ZN( us21_n811 ) );
  NAND2_X1 us21_U349 (.A1( us21_n451 ) , .A2( us21_n459 ) , .ZN( us21_n742 ) );
  NOR4_X1 us21_U35 (.A4( us21_n732 ) , .A3( us21_n733 ) , .A2( us21_n734 ) , .A1( us21_n735 ) , .ZN( us21_n736 ) );
  NAND2_X1 us21_U350 (.A1( us21_n449 ) , .A2( us21_n452 ) , .ZN( us21_n812 ) );
  NAND2_X1 us21_U351 (.A1( us21_n453 ) , .A2( us21_n460 ) , .ZN( us21_n748 ) );
  NAND2_X1 us21_U352 (.A1( us21_n449 ) , .A2( us21_n469 ) , .ZN( us21_n814 ) );
  NAND2_X1 us21_U353 (.A1( us21_n450 ) , .A2( us21_n463 ) , .ZN( us21_n667 ) );
  NAND2_X1 us21_U354 (.A2( us21_n446 ) , .A1( us21_n458 ) , .ZN( us21_n726 ) );
  NAND2_X1 us21_U355 (.A1( us21_n451 ) , .A2( us21_n470 ) , .ZN( us21_n783 ) );
  NAND2_X1 us21_U356 (.A2( us21_n452 ) , .A1( us21_n470 ) , .ZN( us21_n777 ) );
  NAND2_X1 us21_U357 (.A2( us21_n451 ) , .A1( us21_n453 ) , .ZN( us21_n804 ) );
  NAND2_X1 us21_U358 (.A2( us21_n462 ) , .A1( us21_n463 ) , .ZN( us21_n810 ) );
  NAND2_X1 us21_U359 (.A1( us21_n439 ) , .A2( us21_n458 ) , .ZN( us21_n697 ) );
  AOI211_X1 us21_U36 (.B( us21_n723 ) , .A( us21_n724 ) , .ZN( us21_n737 ) , .C1( us21_n841 ) , .C2( us21_n853 ) );
  NAND2_X1 us21_U360 (.A2( us21_n447 ) , .A1( us21_n450 ) , .ZN( us21_n761 ) );
  NAND2_X1 us21_U361 (.A2( us21_n446 ) , .A1( us21_n450 ) , .ZN( us21_n727 ) );
  NOR2_X1 us21_U362 (.ZN( us21_n445 ) , .A2( us21_n847 ) , .A1( us21_n856 ) );
  NAND2_X1 us21_U363 (.A1( us21_n460 ) , .A2( us21_n470 ) , .ZN( us21_n786 ) );
  NOR2_X1 us21_U364 (.ZN( us21_n463 ) , .A2( us21_n845 ) , .A1( us21_n846 ) );
  NOR2_X1 us21_U365 (.ZN( us21_n451 ) , .A1( us21_n824 ) , .A2( us21_n825 ) );
  NAND2_X1 us21_U366 (.A2( us21_n459 ) , .A1( us21_n460 ) , .ZN( us21_n745 ) );
  NOR2_X1 us21_U367 (.ZN( us21_n449 ) , .A1( us21_n826 ) , .A2( us21_n827 ) );
  NAND2_X1 us21_U368 (.A2( us21_n459 ) , .A1( us21_n469 ) , .ZN( us21_n695 ) );
  NAND2_X1 us21_U369 (.A2( us21_n452 ) , .A1( us21_n453 ) , .ZN( us21_n728 ) );
  NOR3_X1 us21_U37 (.A3( us21_n720 ) , .A1( us21_n721 ) , .ZN( us21_n738 ) , .A2( us21_n739 ) );
  NAND2_X1 us21_U370 (.A1( us21_n449 ) , .A2( us21_n460 ) , .ZN( us21_n788 ) );
  NAND2_X2 us21_U371 (.A2( us21_n446 ) , .A1( us21_n462 ) , .ZN( us21_n813 ) );
  NAND2_X2 us21_U372 (.A2( us21_n439 ) , .A1( us21_n450 ) , .ZN( us21_n789 ) );
  NAND2_X2 us21_U373 (.A1( us21_n447 ) , .A2( us21_n458 ) , .ZN( us21_n790 ) );
  NAND2_X2 us21_U374 (.A1( us21_n439 ) , .A2( us21_n462 ) , .ZN( us21_n706 ) );
  NAND2_X2 us21_U375 (.A2( us21_n469 ) , .A1( us21_n470 ) , .ZN( us21_n815 ) );
  NAND2_X2 us21_U376 (.A1( us21_n445 ) , .A2( us21_n446 ) , .ZN( us21_n784 ) );
  NOR2_X1 us21_U377 (.A2( sa21_6 ) , .A1( sa21_7 ) , .ZN( us21_n462 ) );
  NOR2_X1 us21_U378 (.A2( sa21_4 ) , .ZN( us21_n447 ) , .A1( us21_n846 ) );
  NOR2_X1 us21_U379 (.A2( sa21_5 ) , .ZN( us21_n446 ) , .A1( us21_n845 ) );
  NAND4_X1 us21_U38 (.ZN( sa23_sr_3 ) , .A4( us21_n702 ) , .A3( us21_n703 ) , .A2( us21_n704 ) , .A1( us21_n705 ) );
  NOR2_X1 us21_U380 (.A2( sa21_7 ) , .ZN( us21_n458 ) , .A1( us21_n847 ) );
  NOR2_X1 us21_U381 (.A2( sa21_4 ) , .A1( sa21_5 ) , .ZN( us21_n439 ) );
  NOR2_X1 us21_U382 (.A2( sa21_1 ) , .ZN( us21_n469 ) , .A1( us21_n824 ) );
  NOR2_X1 us21_U383 (.A2( sa21_2 ) , .A1( sa21_3 ) , .ZN( us21_n470 ) );
  NOR2_X1 us21_U384 (.A2( sa21_6 ) , .ZN( us21_n450 ) , .A1( us21_n856 ) );
  NOR2_X1 us21_U385 (.A2( sa21_2 ) , .ZN( us21_n459 ) , .A1( us21_n827 ) );
  NOR2_X1 us21_U386 (.A2( sa21_0 ) , .ZN( us21_n452 ) , .A1( us21_n825 ) );
  NOR2_X1 us21_U387 (.A2( sa21_0 ) , .A1( sa21_1 ) , .ZN( us21_n460 ) );
  NOR2_X1 us21_U388 (.A2( sa21_3 ) , .ZN( us21_n453 ) , .A1( us21_n826 ) );
  INV_X1 us21_U389 (.A( sa21_6 ) , .ZN( us21_n847 ) );
  NOR4_X1 us21_U39 (.A4( us21_n698 ) , .A3( us21_n699 ) , .A2( us21_n700 ) , .A1( us21_n701 ) , .ZN( us21_n702 ) );
  INV_X1 us21_U390 (.A( sa21_3 ) , .ZN( us21_n827 ) );
  INV_X1 us21_U391 (.A( sa21_1 ) , .ZN( us21_n825 ) );
  INV_X1 us21_U392 (.A( sa21_0 ) , .ZN( us21_n824 ) );
  INV_X1 us21_U393 (.A( sa21_2 ) , .ZN( us21_n826 ) );
  INV_X1 us21_U394 (.A( sa21_5 ) , .ZN( us21_n846 ) );
  INV_X1 us21_U395 (.A( sa21_7 ) , .ZN( us21_n856 ) );
  INV_X1 us21_U396 (.A( us21_n784 ) , .ZN( us21_n860 ) );
  AOI21_X1 us21_U397 (.ZN( us21_n498 ) , .A( us21_n695 ) , .B1( us21_n706 ) , .B2( us21_n784 ) );
  INV_X1 us21_U398 (.A( us21_n695 ) , .ZN( us21_n836 ) );
  NOR2_X1 us21_U399 (.A1( us21_n695 ) , .ZN( us21_n768 ) , .A2( us21_n813 ) );
  NAND2_X1 us21_U4 (.A1( us21_n447 ) , .A2( us21_n462 ) , .ZN( us21_n722 ) );
  AOI211_X1 us21_U40 (.B( us21_n692 ) , .A( us21_n693 ) , .ZN( us21_n703 ) , .C2( us21_n829 ) , .C1( us21_n849 ) );
  AOI21_X1 us21_U400 (.ZN( us21_n569 ) , .B2( us21_n695 ) , .B1( us21_n804 ) , .A( us21_n810 ) );
  NOR2_X1 us21_U401 (.ZN( us21_n630 ) , .A2( us21_n695 ) , .A1( us21_n722 ) );
  AOI21_X1 us21_U402 (.ZN( us21_n476 ) , .B2( us21_n695 ) , .A( us21_n747 ) , .B1( us21_n777 ) );
  NOR2_X1 us21_U403 (.ZN( us21_n660 ) , .A2( us21_n695 ) , .A1( us21_n727 ) );
  NOR2_X1 us21_U404 (.A2( us21_n695 ) , .A1( us21_n778 ) , .ZN( us21_n818 ) );
  NOR2_X1 us21_U405 (.A2( us21_n695 ) , .ZN( us21_n714 ) , .A1( us21_n790 ) );
  NOR2_X1 us21_U406 (.ZN( us21_n564 ) , .A2( us21_n695 ) , .A1( us21_n761 ) );
  NOR2_X1 us21_U407 (.ZN( us21_n592 ) , .A2( us21_n695 ) , .A1( us21_n726 ) );
  AOI21_X1 us21_U408 (.ZN( us21_n550 ) , .B1( us21_n667 ) , .A( us21_n695 ) , .B2( us21_n803 ) );
  NOR2_X1 us21_U409 (.ZN( us21_n539 ) , .A2( us21_n695 ) , .A1( us21_n697 ) );
  NOR2_X1 us21_U41 (.ZN( us21_n705 ) , .A2( us21_n774 ) , .A1( us21_n798 ) );
  NOR2_X1 us21_U410 (.ZN( us21_n578 ) , .A2( us21_n695 ) , .A1( us21_n789 ) );
  OAI222_X1 us21_U411 (.B2( us21_n745 ) , .B1( us21_n746 ) , .A2( us21_n747 ) , .ZN( us21_n755 ) , .C2( us21_n803 ) , .C1( us21_n812 ) , .A1( us21_n815 ) );
  OAI222_X1 us21_U412 (.ZN( us21_n503 ) , .C2( us21_n623 ) , .B2( us21_n645 ) , .B1( us21_n745 ) , .A2( us21_n746 ) , .C1( us21_n803 ) , .A1( us21_n804 ) );
  AOI222_X1 us21_U413 (.ZN( us21_n511 ) , .C1( us21_n830 ) , .B2( us21_n835 ) , .A2( us21_n841 ) , .C2( us21_n860 ) , .B1( us21_n861 ) , .A1( us21_n864 ) );
  AOI222_X1 us21_U414 (.ZN( us21_n603 ) , .B2( us21_n669 ) , .B1( us21_n751 ) , .C2( us21_n829 ) , .A1( us21_n831 ) , .A2( us21_n860 ) , .C1( us21_n861 ) );
  AOI221_X1 us21_U415 (.A( us21_n481 ) , .ZN( us21_n486 ) , .B1( us21_n829 ) , .C2( us21_n842 ) , .C1( us21_n850 ) , .B2( us21_n860 ) );
  NOR2_X1 us21_U416 (.ZN( us21_n787 ) , .A2( us21_n860 ) , .A1( us21_n866 ) );
  OAI221_X1 us21_U417 (.A( us21_n781 ) , .C2( us21_n782 ) , .B2( us21_n783 ) , .B1( us21_n784 ) , .ZN( us21_n794 ) , .C1( us21_n811 ) );
  NAND2_X1 us21_U418 (.A1( us21_n727 ) , .A2( us21_n782 ) , .ZN( us21_n809 ) );
  OAI22_X1 us21_U419 (.ZN( us21_n586 ) , .A2( us21_n745 ) , .B2( us21_n760 ) , .A1( us21_n761 ) , .B1( us21_n782 ) );
  NOR2_X1 us21_U42 (.ZN( us21_n802 ) , .A1( us21_n852 ) , .A2( us21_n859 ) );
  OAI221_X1 us21_U420 (.A( us21_n694 ) , .ZN( us21_n701 ) , .C2( us21_n782 ) , .C1( us21_n783 ) , .B1( us21_n784 ) , .B2( us21_n804 ) );
  AOI21_X1 us21_U421 (.ZN( us21_n590 ) , .B1( us21_n726 ) , .B2( us21_n782 ) , .A( us21_n788 ) );
  AOI21_X1 us21_U422 (.ZN( us21_n646 ) , .A( us21_n760 ) , .B2( us21_n782 ) , .B1( us21_n790 ) );
  AOI21_X1 us21_U423 (.ZN( us21_n621 ) , .B1( us21_n697 ) , .A( us21_n777 ) , .B2( us21_n782 ) );
  OAI22_X1 us21_U424 (.ZN( us21_n679 ) , .A1( us21_n697 ) , .A2( us21_n728 ) , .B2( us21_n782 ) , .B1( us21_n815 ) );
  OAI21_X1 us21_U425 (.A( us21_n611 ) , .ZN( us21_n614 ) , .B1( us21_n623 ) , .B2( us21_n782 ) );
  NOR2_X1 us21_U426 (.ZN( us21_n608 ) , .A1( us21_n782 ) , .A2( us21_n814 ) );
  OAI222_X1 us21_U427 (.A2( us21_n667 ) , .ZN( us21_n672 ) , .B1( us21_n745 ) , .B2( us21_n782 ) , .C2( us21_n786 ) , .C1( us21_n813 ) , .A1( us21_n815 ) );
  NOR2_X1 us21_U428 (.ZN( us21_n649 ) , .A1( us21_n782 ) , .A2( us21_n786 ) );
  NOR2_X1 us21_U429 (.ZN( us21_n598 ) , .A2( us21_n695 ) , .A1( us21_n782 ) );
  NAND4_X1 us21_U43 (.ZN( sa23_sr_2 ) , .A4( us21_n641 ) , .A3( us21_n642 ) , .A2( us21_n643 ) , .A1( us21_n644 ) );
  NOR2_X1 us21_U430 (.ZN( us21_n551 ) , .A2( us21_n742 ) , .A1( us21_n782 ) );
  INV_X1 us21_U431 (.A( us21_n782 ) , .ZN( us21_n859 ) );
  AOI221_X1 us21_U432 (.A( us21_n574 ) , .ZN( us21_n585 ) , .B2( us21_n829 ) , .C2( us21_n841 ) , .B1( us21_n852 ) , .C1( us21_n859 ) );
  AOI21_X1 us21_U433 (.ZN( us21_n574 ) , .B2( us21_n722 ) , .B1( us21_n746 ) , .A( us21_n783 ) );
  INV_X1 us21_U434 (.A( sa21_4 ) , .ZN( us21_n845 ) );
  AOI211_X1 us21_U435 (.A( us21_n635 ) , .ZN( us21_n643 ) , .B( us21_n741 ) , .C2( us21_n837 ) , .C1( us21_n852 ) );
  NAND4_X1 us21_U436 (.A4( us21_n631 ) , .A3( us21_n632 ) , .A2( us21_n633 ) , .A1( us21_n634 ) , .ZN( us21_n741 ) );
  NAND3_X1 us21_U437 (.ZN( sa23_sr_6 ) , .A3( us21_n795 ) , .A2( us21_n796 ) , .A1( us21_n797 ) );
  NAND3_X1 us21_U438 (.ZN( sa23_sr_5 ) , .A3( us21_n756 ) , .A2( us21_n757 ) , .A1( us21_n758 ) );
  NAND3_X1 us21_U439 (.ZN( sa23_sr_4 ) , .A3( us21_n736 ) , .A2( us21_n737 ) , .A1( us21_n738 ) );
  AOI222_X1 us21_U44 (.B2( us21_n636 ) , .ZN( us21_n642 ) , .B1( us21_n839 ) , .A1( us21_n840 ) , .C2( us21_n844 ) , .C1( us21_n861 ) , .A2( us21_n863 ) );
  NAND3_X1 us21_U440 (.A3( us21_n673 ) , .A2( us21_n674 ) , .A1( us21_n675 ) , .ZN( us21_n805 ) );
  NAND3_X1 us21_U441 (.ZN( us21_n636 ) , .A3( us21_n706 ) , .A2( us21_n722 ) , .A1( us21_n790 ) );
  NAND3_X1 us21_U442 (.A3( us21_n616 ) , .A2( us21_n617 ) , .A1( us21_n618 ) , .ZN( us21_n723 ) );
  NAND3_X1 us21_U443 (.A3( us21_n583 ) , .A2( us21_n584 ) , .A1( us21_n585 ) , .ZN( us21_n619 ) );
  NAND3_X1 us21_U444 (.ZN( us21_n563 ) , .A3( us21_n678 ) , .A2( us21_n748 ) , .A1( us21_n783 ) );
  NAND3_X1 us21_U445 (.A3( us21_n521 ) , .A2( us21_n522 ) , .A1( us21_n523 ) , .ZN( us21_n740 ) );
  NAND3_X1 us21_U446 (.A3( us21_n510 ) , .A1( us21_n511 ) , .ZN( us21_n606 ) , .A2( us21_n869 ) );
  NAND3_X1 us21_U447 (.A3( us21_n465 ) , .A2( us21_n466 ) , .A1( us21_n467 ) , .ZN( us21_n775 ) );
  NOR4_X1 us21_U45 (.A4( us21_n637 ) , .A3( us21_n638 ) , .A2( us21_n639 ) , .A1( us21_n640 ) , .ZN( us21_n641 ) );
  NOR3_X1 us21_U46 (.A2( us21_n605 ) , .A1( us21_n606 ) , .ZN( us21_n644 ) , .A3( us21_n720 ) );
  NAND4_X1 us21_U47 (.ZN( sa23_sr_0 ) , .A4( us21_n499 ) , .A3( us21_n500 ) , .A2( us21_n501 ) , .A1( us21_n502 ) );
  NOR4_X1 us21_U48 (.A4( us21_n496 ) , .A3( us21_n497 ) , .A2( us21_n498 ) , .ZN( us21_n499 ) , .A1( us21_n525 ) );
  AOI221_X1 us21_U49 (.A( us21_n495 ) , .ZN( us21_n500 ) , .B2( us21_n841 ) , .C1( us21_n844 ) , .C2( us21_n858 ) , .B1( us21_n860 ) );
  NAND2_X1 us21_U5 (.A1( us21_n445 ) , .A2( us21_n447 ) , .ZN( us21_n803 ) );
  AOI211_X1 us21_U50 (.A( us21_n494 ) , .ZN( us21_n501 ) , .B( us21_n800 ) , .C2( us21_n837 ) , .C1( us21_n849 ) );
  NAND4_X1 us21_U51 (.ZN( sa23_sr_1 ) , .A4( us21_n593 ) , .A3( us21_n594 ) , .A2( us21_n595 ) , .A1( us21_n596 ) );
  AOI211_X1 us21_U52 (.B( us21_n587 ) , .A( us21_n588 ) , .ZN( us21_n594 ) , .C2( us21_n809 ) , .C1( us21_n831 ) );
  NOR4_X1 us21_U53 (.A4( us21_n589 ) , .A3( us21_n590 ) , .A2( us21_n591 ) , .A1( us21_n592 ) , .ZN( us21_n593 ) );
  AOI211_X1 us21_U54 (.A( us21_n586 ) , .ZN( us21_n595 ) , .B( us21_n619 ) , .C1( us21_n843 ) , .C2( us21_n853 ) );
  NAND4_X1 us21_U55 (.A4( us21_n601 ) , .A3( us21_n602 ) , .A2( us21_n603 ) , .A1( us21_n604 ) , .ZN( us21_n720 ) );
  NOR3_X1 us21_U56 (.A1( us21_n597 ) , .ZN( us21_n602 ) , .A3( us21_n661 ) , .A2( us21_n768 ) );
  NOR4_X1 us21_U57 (.A3( us21_n598 ) , .A2( us21_n599 ) , .A1( us21_n600 ) , .ZN( us21_n601 ) , .A4( us21_n653 ) );
  AOI222_X1 us21_U58 (.ZN( us21_n604 ) , .A1( us21_n828 ) , .C2( us21_n835 ) , .B1( us21_n840 ) , .A2( us21_n854 ) , .B2( us21_n859 ) , .C1( us21_n866 ) );
  AOI222_X1 us21_U59 (.ZN( us21_n467 ) , .B1( us21_n830 ) , .A1( us21_n837 ) , .C1( us21_n840 ) , .C2( us21_n849 ) , .A2( us21_n853 ) , .B2( us21_n863 ) );
  NOR3_X1 us21_U6 (.ZN( us21_n596 ) , .A1( us21_n606 ) , .A3( us21_n721 ) , .A2( us21_n740 ) );
  NOR4_X1 us21_U60 (.A1( us21_n464 ) , .ZN( us21_n465 ) , .A4( us21_n540 ) , .A2( us21_n552 ) , .A3( us21_n612 ) );
  AOI221_X1 us21_U61 (.ZN( us21_n466 ) , .C2( us21_n712 ) , .B2( us21_n829 ) , .C1( us21_n843 ) , .B1( us21_n858 ) , .A( us21_n862 ) );
  NAND4_X1 us21_U62 (.A4( us21_n483 ) , .A3( us21_n484 ) , .A2( us21_n485 ) , .A1( us21_n486 ) , .ZN( us21_n776 ) );
  NOR4_X1 us21_U63 (.ZN( us21_n484 ) , .A1( us21_n505 ) , .A2( us21_n517 ) , .A4( us21_n544 ) , .A3( us21_n609 ) );
  NOR4_X1 us21_U64 (.A4( us21_n482 ) , .ZN( us21_n485 ) , .A1( us21_n564 ) , .A2( us21_n579 ) , .A3( us21_n600 ) );
  NOR4_X1 us21_U65 (.ZN( us21_n483 ) , .A2( us21_n531 ) , .A1( us21_n556 ) , .A3( us21_n629 ) , .A4( us21_n716 ) );
  AOI211_X1 us21_U66 (.B( us21_n621 ) , .A( us21_n622 ) , .ZN( us21_n633 ) , .C2( us21_n834 ) , .C1( us21_n861 ) );
  NOR4_X1 us21_U67 (.A4( us21_n627 ) , .A3( us21_n628 ) , .A2( us21_n629 ) , .A1( us21_n630 ) , .ZN( us21_n631 ) );
  NOR4_X1 us21_U68 (.A4( us21_n624 ) , .A3( us21_n625 ) , .A2( us21_n626 ) , .ZN( us21_n632 ) , .A1( us21_n662 ) );
  NOR4_X1 us21_U69 (.A4( us21_n512 ) , .A3( us21_n513 ) , .A2( us21_n514 ) , .A1( us21_n515 ) , .ZN( us21_n522 ) );
  NOR3_X1 us21_U7 (.A3( us21_n798 ) , .A2( us21_n799 ) , .A1( us21_n800 ) , .ZN( us21_n823 ) );
  AOI222_X1 us21_U70 (.ZN( us21_n523 ) , .A1( us21_n832 ) , .B2( us21_n835 ) , .C1( us21_n842 ) , .C2( us21_n848 ) , .A2( us21_n850 ) , .B1( us21_n864 ) );
  NOR4_X1 us21_U71 (.A3( us21_n519 ) , .A1( us21_n520 ) , .ZN( us21_n521 ) , .A2( us21_n671 ) , .A4( us21_n767 ) );
  NAND4_X1 us21_U72 (.A4( us21_n655 ) , .A3( us21_n656 ) , .A2( us21_n657 ) , .A1( us21_n658 ) , .ZN( us21_n798 ) );
  NOR3_X1 us21_U73 (.A3( us21_n646 ) , .A2( us21_n647 ) , .A1( us21_n648 ) , .ZN( us21_n657 ) );
  NOR3_X1 us21_U74 (.A3( us21_n649 ) , .A2( us21_n650 ) , .A1( us21_n651 ) , .ZN( us21_n656 ) );
  NOR3_X1 us21_U75 (.A3( us21_n652 ) , .A2( us21_n653 ) , .A1( us21_n654 ) , .ZN( us21_n655 ) );
  NAND4_X1 us21_U76 (.A4( us21_n558 ) , .A3( us21_n559 ) , .A2( us21_n560 ) , .A1( us21_n561 ) , .ZN( us21_n605 ) );
  NOR4_X1 us21_U77 (.A4( us21_n550 ) , .A3( us21_n551 ) , .A2( us21_n552 ) , .A1( us21_n553 ) , .ZN( us21_n560 ) );
  NOR4_X1 us21_U78 (.A4( us21_n554 ) , .A3( us21_n555 ) , .A2( us21_n556 ) , .A1( us21_n557 ) , .ZN( us21_n558 ) );
  NOR4_X1 us21_U79 (.ZN( us21_n559 ) , .A1( us21_n651 ) , .A3( us21_n659 ) , .A4( us21_n683 ) , .A2( us21_n766 ) );
  NOR3_X1 us21_U8 (.ZN( us21_n502 ) , .A2( us21_n677 ) , .A3( us21_n775 ) , .A1( us21_n874 ) );
  NAND4_X1 us21_U80 (.A4( us21_n770 ) , .A3( us21_n771 ) , .A2( us21_n772 ) , .A1( us21_n773 ) , .ZN( us21_n799 ) );
  NOR3_X1 us21_U81 (.A3( us21_n763 ) , .A2( us21_n764 ) , .A1( us21_n765 ) , .ZN( us21_n771 ) );
  NOR4_X1 us21_U82 (.A4( us21_n766 ) , .A3( us21_n767 ) , .A2( us21_n768 ) , .A1( us21_n769 ) , .ZN( us21_n770 ) );
  AOI222_X1 us21_U83 (.ZN( us21_n773 ) , .A1( us21_n828 ) , .C1( us21_n832 ) , .B2( us21_n839 ) , .A2( us21_n848 ) , .B1( us21_n859 ) , .C2( us21_n871 ) );
  NOR4_X1 us21_U84 (.A4( us21_n507 ) , .A2( us21_n508 ) , .A1( us21_n509 ) , .ZN( us21_n510 ) , .A3( us21_n668 ) );
  INV_X1 us21_U85 (.A( us21_n503 ) , .ZN( us21_n869 ) );
  NOR4_X1 us21_U86 (.A4( us21_n659 ) , .A3( us21_n660 ) , .A2( us21_n661 ) , .A1( us21_n662 ) , .ZN( us21_n675 ) );
  NOR4_X1 us21_U87 (.A4( us21_n663 ) , .A3( us21_n664 ) , .A2( us21_n665 ) , .A1( us21_n666 ) , .ZN( us21_n674 ) );
  NOR4_X1 us21_U88 (.A3( us21_n671 ) , .A1( us21_n672 ) , .ZN( us21_n673 ) , .A4( us21_n713 ) , .A2( us21_n857 ) );
  NOR2_X1 us21_U89 (.ZN( us21_n623 ) , .A2( us21_n834 ) , .A1( us21_n837 ) );
  INV_X1 us21_U9 (.A( us21_n704 ) , .ZN( us21_n874 ) );
  NOR2_X1 us21_U90 (.ZN( us21_n759 ) , .A1( us21_n831 ) , .A2( us21_n832 ) );
  NAND4_X1 us21_U91 (.A4( us21_n454 ) , .A3( us21_n455 ) , .A2( us21_n456 ) , .A1( us21_n457 ) , .ZN( us21_n677 ) );
  NOR3_X1 us21_U92 (.ZN( us21_n455 ) , .A3( us21_n528 ) , .A1( us21_n553 ) , .A2( us21_n568 ) );
  AOI221_X1 us21_U93 (.A( us21_n448 ) , .ZN( us21_n457 ) , .C2( us21_n751 ) , .B1( us21_n830 ) , .C1( us21_n840 ) , .B2( us21_n859 ) );
  NOR4_X1 us21_U94 (.ZN( us21_n456 ) , .A2( us21_n507 ) , .A1( us21_n597 ) , .A4( us21_n626 ) , .A3( us21_n709 ) );
  NAND4_X1 us21_U95 (.ZN( sa23_sr_7 ) , .A4( us21_n820 ) , .A3( us21_n821 ) , .A2( us21_n822 ) , .A1( us21_n823 ) );
  NOR4_X1 us21_U96 (.A4( us21_n816 ) , .A3( us21_n817 ) , .A2( us21_n818 ) , .A1( us21_n819 ) , .ZN( us21_n820 ) );
  AOI222_X1 us21_U97 (.C2( us21_n807 ) , .B2( us21_n808 ) , .A2( us21_n809 ) , .ZN( us21_n821 ) , .C1( us21_n830 ) , .A1( us21_n837 ) , .B1( us21_n851 ) );
  AOI211_X1 us21_U98 (.B( us21_n805 ) , .A( us21_n806 ) , .ZN( us21_n822 ) , .C1( us21_n840 ) , .C2( us21_n848 ) );
  NAND4_X1 us21_U99 (.A4( us21_n533 ) , .A3( us21_n534 ) , .A2( us21_n535 ) , .A1( us21_n536 ) , .ZN( us21_n620 ) );
  INV_X1 us23_U10 (.A( us23_n679 ) , .ZN( us23_n839 ) );
  NOR4_X1 us23_U100 (.A4( us23_n483 ) , .ZN( us23_n486 ) , .A1( us23_n565 ) , .A2( us23_n580 ) , .A3( us23_n601 ) );
  NOR4_X1 us23_U101 (.ZN( us23_n485 ) , .A1( us23_n506 ) , .A2( us23_n518 ) , .A4( us23_n545 ) , .A3( us23_n610 ) );
  NOR4_X1 us23_U102 (.ZN( us23_n484 ) , .A2( us23_n532 ) , .A1( us23_n557 ) , .A3( us23_n630 ) , .A4( us23_n717 ) );
  NAND4_X1 us23_U103 (.A4( us23_n690 ) , .A3( us23_n691 ) , .A1( us23_n692 ) , .ZN( us23_n775 ) , .A2( us23_n871 ) );
  AOI221_X1 us23_U104 (.A( us23_n680 ) , .ZN( us23_n691 ) , .B2( us23_n839 ) , .C1( us23_n841 ) , .C2( us23_n861 ) , .B1( us23_n864 ) );
  INV_X1 us23_U105 (.A( us23_n678 ) , .ZN( us23_n871 ) );
  NOR4_X1 us23_U106 (.A4( us23_n686 ) , .A3( us23_n687 ) , .A2( us23_n688 ) , .A1( us23_n689 ) , .ZN( us23_n690 ) );
  NAND4_X1 us23_U107 (.A4( us23_n559 ) , .A3( us23_n560 ) , .A2( us23_n561 ) , .A1( us23_n562 ) , .ZN( us23_n606 ) );
  NOR4_X1 us23_U108 (.ZN( us23_n560 ) , .A1( us23_n652 ) , .A3( us23_n660 ) , .A4( us23_n684 ) , .A2( us23_n767 ) );
  NOR4_X1 us23_U109 (.A4( us23_n551 ) , .A3( us23_n552 ) , .A2( us23_n553 ) , .A1( us23_n554 ) , .ZN( us23_n561 ) );
  NOR4_X1 us23_U11 (.A4( us23_n444 ) , .A3( us23_n445 ) , .A2( us23_n515 ) , .A1( us23_n540 ) , .ZN( us23_n705 ) );
  NOR4_X1 us23_U110 (.A4( us23_n555 ) , .A3( us23_n556 ) , .A2( us23_n557 ) , .A1( us23_n558 ) , .ZN( us23_n559 ) );
  NAND4_X1 us23_U111 (.A4( us23_n718 ) , .A3( us23_n719 ) , .A2( us23_n720 ) , .ZN( us23_n740 ) , .A1( us23_n856 ) );
  INV_X1 us23_U112 (.A( us23_n708 ) , .ZN( us23_n856 ) );
  AOI221_X1 us23_U113 (.A( us23_n709 ) , .ZN( us23_n720 ) , .C2( us23_n843 ) , .B2( us23_n844 ) , .C1( us23_n860 ) , .B1( us23_n861 ) );
  NOR4_X1 us23_U114 (.A4( us23_n714 ) , .A3( us23_n715 ) , .A2( us23_n716 ) , .A1( us23_n717 ) , .ZN( us23_n718 ) );
  NAND4_X1 us23_U115 (.A4( us23_n472 ) , .A3( us23_n473 ) , .A2( us23_n474 ) , .A1( us23_n475 ) , .ZN( us23_n677 ) );
  NOR4_X1 us23_U116 (.A4( us23_n469 ) , .ZN( us23_n475 ) , .A3( us23_n555 ) , .A1( us23_n734 ) , .A2( us23_n754 ) );
  NOR4_X1 us23_U117 (.ZN( us23_n474 ) , .A1( us23_n530 ) , .A3( us23_n567 ) , .A4( us23_n599 ) , .A2( us23_n641 ) );
  NOR4_X1 us23_U118 (.ZN( us23_n473 ) , .A1( us23_n505 ) , .A3( us23_n543 ) , .A2( us23_n582 ) , .A4( us23_n715 ) );
  NOR2_X1 us23_U119 (.ZN( us23_n732 ) , .A2( us23_n831 ) , .A1( us23_n844 ) );
  OR3_X1 us23_U12 (.ZN( us23_n445 ) , .A1( us23_n527 ) , .A3( us23_n576 ) , .A2( us23_n874 ) );
  NOR2_X1 us23_U120 (.ZN( us23_n788 ) , .A2( us23_n861 ) , .A1( us23_n867 ) );
  NAND4_X1 us23_U121 (.A4( us23_n572 ) , .A3( us23_n573 ) , .A1( us23_n574 ) , .ZN( us23_n722 ) , .A2( us23_n873 ) );
  NOR4_X1 us23_U122 (.A4( us23_n568 ) , .A3( us23_n569 ) , .A2( us23_n570 ) , .A1( us23_n571 ) , .ZN( us23_n572 ) );
  AOI221_X1 us23_U123 (.A( us23_n563 ) , .C2( us23_n564 ) , .ZN( us23_n573 ) , .B2( us23_n844 ) , .B1( us23_n851 ) , .C1( us23_n852 ) );
  INV_X1 us23_U124 (.A( us23_n606 ) , .ZN( us23_n873 ) );
  NAND4_X1 us23_U125 (.A4( us23_n492 ) , .A3( us23_n493 ) , .A1( us23_n494 ) , .ZN( us23_n801 ) , .A2( us23_n866 ) );
  AOI221_X1 us23_U126 (.A( us23_n488 ) , .ZN( us23_n493 ) , .B2( us23_n835 ) , .C2( us23_n840 ) , .C1( us23_n850 ) , .B1( us23_n859 ) );
  INV_X1 us23_U127 (.A( us23_n777 ) , .ZN( us23_n866 ) );
  NOR2_X1 us23_U128 (.ZN( us23_n494 ) , .A1( us23_n677 ) , .A2( us23_n693 ) );
  NOR2_X1 us23_U129 (.ZN( us23_n747 ) , .A1( us23_n860 ) , .A2( us23_n861 ) );
  OR4_X1 us23_U13 (.A4( us23_n441 ) , .A2( us23_n442 ) , .A1( us23_n443 ) , .ZN( us23_n444 ) , .A3( us23_n552 ) );
  AOI222_X1 us23_U130 (.ZN( us23_n512 ) , .C1( us23_n831 ) , .B2( us23_n836 ) , .A2( us23_n842 ) , .C2( us23_n861 ) , .B1( us23_n862 ) , .A1( us23_n865 ) );
  NOR4_X1 us23_U131 (.A4( us23_n508 ) , .A2( us23_n509 ) , .A1( us23_n510 ) , .ZN( us23_n511 ) , .A3( us23_n669 ) );
  INV_X1 us23_U132 (.A( us23_n504 ) , .ZN( us23_n870 ) );
  INV_X1 us23_U133 (.A( us23_n761 ) , .ZN( us23_n829 ) );
  NOR2_X1 us23_U134 (.ZN( us23_n646 ) , .A1( us23_n853 ) , .A2( us23_n867 ) );
  OR4_X1 us23_U135 (.A4( us23_n579 ) , .A3( us23_n580 ) , .A2( us23_n581 ) , .A1( us23_n582 ) , .ZN( us23_n583 ) );
  OR4_X1 us23_U136 (.A4( us23_n681 ) , .A3( us23_n682 ) , .A2( us23_n683 ) , .A1( us23_n684 ) , .ZN( us23_n689 ) );
  OR4_X1 us23_U137 (.A4( us23_n565 ) , .A3( us23_n566 ) , .A2( us23_n567 ) , .ZN( us23_n571 ) , .A1( us23_n664 ) );
  OR4_X1 us23_U138 (.A4( us23_n517 ) , .A2( us23_n518 ) , .A1( us23_n519 ) , .ZN( us23_n521 ) , .A3( us23_n820 ) );
  OR4_X1 us23_U139 (.ZN( us23_n465 ) , .A4( us23_n517 ) , .A3( us23_n528 ) , .A2( us23_n577 ) , .A1( us23_n711 ) );
  INV_X1 us23_U14 (.A( us23_n612 ) , .ZN( us23_n874 ) );
  NAND2_X1 us23_U140 (.ZN( us23_n612 ) , .A2( us23_n836 ) , .A1( us23_n872 ) );
  OR3_X1 us23_U141 (.A3( us23_n505 ) , .A2( us23_n506 ) , .A1( us23_n507 ) , .ZN( us23_n510 ) );
  AOI221_X1 us23_U142 (.A( us23_n712 ) , .B2( us23_n713 ) , .ZN( us23_n719 ) , .C1( us23_n831 ) , .B1( us23_n838 ) , .C2( us23_n862 ) );
  OR2_X1 us23_U143 (.A2( us23_n710 ) , .A1( us23_n711 ) , .ZN( us23_n712 ) );
  INV_X1 us23_U144 (.A( us23_n462 ) , .ZN( us23_n863 ) );
  OAI21_X1 us23_U145 (.ZN( us23_n462 ) , .B1( us23_n808 ) , .A( us23_n833 ) , .B2( us23_n850 ) );
  INV_X1 us23_U146 (.A( us23_n753 ) , .ZN( us23_n868 ) );
  OAI21_X1 us23_U147 (.B1( us23_n752 ) , .ZN( us23_n753 ) , .A( us23_n844 ) , .B2( us23_n867 ) );
  INV_X1 us23_U148 (.A( us23_n671 ) , .ZN( us23_n858 ) );
  AOI21_X1 us23_U149 (.A( us23_n669 ) , .B1( us23_n670 ) , .ZN( us23_n671 ) , .B2( us23_n855 ) );
  INV_X1 us23_U15 (.A( us23_n748 ) , .ZN( us23_n862 ) );
  AOI222_X1 us23_U150 (.ZN( us23_n659 ) , .A2( us23_n838 ) , .B1( us23_n840 ) , .C2( us23_n844 ) , .A1( us23_n859 ) , .C1( us23_n862 ) , .B2( us23_n869 ) );
  INV_X1 us23_U151 (.A( us23_n646 ) , .ZN( us23_n869 ) );
  OAI222_X1 us23_U152 (.B2( us23_n707 ) , .ZN( us23_n708 ) , .C2( us23_n723 ) , .B1( us23_n746 ) , .A1( us23_n805 ) , .C1( us23_n813 ) , .A2( us23_n814 ) );
  OAI222_X1 us23_U153 (.A2( us23_n668 ) , .ZN( us23_n673 ) , .B1( us23_n746 ) , .B2( us23_n783 ) , .C2( us23_n787 ) , .C1( us23_n814 ) , .A1( us23_n816 ) );
  NAND2_X1 us23_U154 (.A1( us23_n446 ) , .A2( us23_n464 ) , .ZN( us23_n748 ) );
  NOR4_X1 us23_U155 (.A2( us23_n490 ) , .A1( us23_n491 ) , .ZN( us23_n492 ) , .A3( us23_n579 ) , .A4( us23_n611 ) );
  OR4_X1 us23_U156 (.ZN( us23_n491 ) , .A4( us23_n533 ) , .A2( us23_n546 ) , .A1( us23_n558 ) , .A3( us23_n631 ) );
  OAI22_X1 us23_U157 (.B1( us23_n489 ) , .ZN( us23_n490 ) , .A1( us23_n685 ) , .A2( us23_n762 ) , .B2( us23_n816 ) );
  NOR3_X1 us23_U158 (.ZN( us23_n489 ) , .A1( us23_n781 ) , .A2( us23_n849 ) , .A3( us23_n862 ) );
  AOI22_X1 us23_U159 (.ZN( us23_n695 ) , .A1( us23_n829 ) , .B2( us23_n842 ) , .A2( us23_n864 ) , .B1( us23_n867 ) );
  AOI222_X1 us23_U16 (.ZN( us23_n604 ) , .B2( us23_n670 ) , .B1( us23_n752 ) , .C2( us23_n830 ) , .A1( us23_n832 ) , .A2( us23_n861 ) , .C1( us23_n862 ) );
  AOI21_X1 us23_U160 (.ZN( us23_n638 ) , .B2( us23_n748 ) , .A( us23_n787 ) , .B1( us23_n811 ) );
  AOI21_X1 us23_U161 (.ZN( us23_n639 ) , .B2( us23_n746 ) , .A( us23_n791 ) , .B1( us23_n802 ) );
  AOI21_X1 us23_U162 (.ZN( us23_n640 ) , .B1( us23_n679 ) , .A( us23_n790 ) , .B2( us23_n816 ) );
  INV_X1 us23_U163 (.A( us23_n729 ) , .ZN( us23_n838 ) );
  AOI221_X1 us23_U164 (.A( us23_n763 ) , .ZN( us23_n773 ) , .C2( us23_n809 ) , .B2( us23_n834 ) , .C1( us23_n854 ) , .B1( us23_n865 ) );
  AOI21_X1 us23_U165 (.B2( us23_n762 ) , .ZN( us23_n763 ) , .A( us23_n787 ) , .B1( us23_n791 ) );
  INV_X1 us23_U166 (.A( us23_n760 ) , .ZN( us23_n834 ) );
  AOI221_X1 us23_U167 (.A( us23_n449 ) , .ZN( us23_n458 ) , .C2( us23_n752 ) , .B1( us23_n831 ) , .C1( us23_n841 ) , .B2( us23_n860 ) );
  AOI21_X1 us23_U168 (.ZN( us23_n449 ) , .B2( us23_n791 ) , .A( us23_n802 ) , .B1( us23_n814 ) );
  AOI221_X1 us23_U169 (.A( us23_n482 ) , .ZN( us23_n487 ) , .B1( us23_n830 ) , .C2( us23_n843 ) , .C1( us23_n851 ) , .B2( us23_n861 ) );
  AOI222_X1 us23_U17 (.ZN( us23_n562 ) , .B1( us23_n829 ) , .C1( us23_n840 ) , .A2( us23_n842 ) , .A1( us23_n853 ) , .B2( us23_n862 ) , .C2( us23_n872 ) );
  OAI22_X1 us23_U170 (.ZN( us23_n482 ) , .A1( us23_n707 ) , .B2( us23_n784 ) , .A2( us23_n805 ) , .B1( us23_n811 ) );
  INV_X1 us23_U171 (.A( us23_n789 ) , .ZN( us23_n831 ) );
  NAND2_X1 us23_U172 (.A1( us23_n450 ) , .A2( us23_n452 ) , .ZN( us23_n761 ) );
  INV_X1 us23_U173 (.A( us23_n783 ) , .ZN( us23_n860 ) );
  INV_X1 us23_U174 (.A( us23_n785 ) , .ZN( us23_n861 ) );
  INV_X1 us23_U175 (.A( us23_n815 ) , .ZN( us23_n830 ) );
  OAI22_X1 us23_U176 (.ZN( us23_n709 ) , .A2( us23_n727 ) , .B2( us23_n728 ) , .A1( us23_n743 ) , .B1( us23_n812 ) );
  OAI22_X1 us23_U177 (.ZN( us23_n623 ) , .B1( us23_n668 ) , .B2( us23_n746 ) , .A1( us23_n814 ) , .A2( us23_n815 ) );
  OAI22_X1 us23_U178 (.ZN( us23_n587 ) , .A2( us23_n746 ) , .B2( us23_n761 ) , .A1( us23_n762 ) , .B1( us23_n783 ) );
  INV_X1 us23_U179 (.A( us23_n743 ) , .ZN( us23_n836 ) );
  NOR4_X1 us23_U18 (.ZN( us23_n472 ) , .A2( us23_n520 ) , .A4( us23_n593 ) , .A1( us23_n608 ) , .A3( us23_n628 ) );
  INV_X1 us23_U180 (.A( us23_n787 ) , .ZN( us23_n844 ) );
  OAI22_X1 us23_U181 (.A1( us23_n723 ) , .ZN( us23_n725 ) , .B2( us23_n749 ) , .B1( us23_n811 ) , .A2( us23_n815 ) );
  OAI22_X1 us23_U182 (.B2( us23_n778 ) , .B1( us23_n779 ) , .ZN( us23_n780 ) , .A2( us23_n813 ) , .A1( us23_n814 ) );
  OAI22_X1 us23_U183 (.ZN( us23_n680 ) , .A1( us23_n698 ) , .A2( us23_n729 ) , .B2( us23_n783 ) , .B1( us23_n816 ) );
  OAI22_X1 us23_U184 (.B2( us23_n749 ) , .B1( us23_n750 ) , .A1( us23_n751 ) , .ZN( us23_n755 ) , .A2( us23_n805 ) );
  NOR2_X1 us23_U185 (.ZN( us23_n750 ) , .A2( us23_n851 ) , .A1( us23_n859 ) );
  NOR3_X1 us23_U186 (.ZN( us23_n751 ) , .A2( us23_n852 ) , .A1( us23_n862 ) , .A3( us23_n864 ) );
  OAI22_X1 us23_U187 (.B2( us23_n743 ) , .ZN( us23_n745 ) , .A2( us23_n761 ) , .B1( us23_n779 ) , .A1( us23_n791 ) );
  INV_X1 us23_U188 (.A( us23_n802 ) , .ZN( us23_n842 ) );
  INV_X1 us23_U189 (.A( us23_n813 ) , .ZN( us23_n832 ) );
  NOR4_X1 us23_U19 (.A4( us23_n531 ) , .A3( us23_n532 ) , .A2( us23_n533 ) , .ZN( us23_n534 ) , .A1( us23_n819 ) );
  INV_X1 us23_U190 (.A( us23_n804 ) , .ZN( us23_n859 ) );
  OAI22_X1 us23_U191 (.B2( us23_n802 ) , .B1( us23_n803 ) , .A2( us23_n804 ) , .A1( us23_n805 ) , .ZN( us23_n807 ) );
  OAI22_X1 us23_U192 (.ZN( us23_n495 ) , .A2( us23_n743 ) , .A1( us23_n779 ) , .B1( us23_n790 ) , .B2( us23_n805 ) );
  OAI22_X1 us23_U193 (.ZN( us23_n488 ) , .A1( us23_n723 ) , .B2( us23_n727 ) , .B1( us23_n729 ) , .A2( us23_n778 ) );
  INV_X1 us23_U194 (.A( us23_n668 ) , .ZN( us23_n864 ) );
  OAI22_X1 us23_U195 (.ZN( us23_n694 ) , .A2( us23_n729 ) , .A1( us23_n779 ) , .B1( us23_n790 ) , .B2( us23_n816 ) );
  OAI22_X1 us23_U196 (.ZN( us23_n636 ) , .A1( us23_n698 ) , .B2( us23_n727 ) , .A2( us23_n761 ) , .B1( us23_n815 ) );
  NOR2_X1 us23_U197 (.A1( us23_n696 ) , .ZN( us23_n769 ) , .A2( us23_n814 ) );
  NOR2_X1 us23_U198 (.ZN( us23_n714 ) , .A1( us23_n804 ) , .A2( us23_n816 ) );
  NOR2_X1 us23_U199 (.ZN( us23_n717 ) , .A2( us23_n723 ) , .A1( us23_n743 ) );
  NOR4_X1 us23_U20 (.ZN( us23_n478 ) , .A1( us23_n519 ) , .A4( us23_n556 ) , .A3( us23_n581 ) , .A2( us23_n629 ) );
  NOR2_X1 us23_U200 (.ZN( us23_n545 ) , .A2( us23_n779 ) , .A1( us23_n813 ) );
  INV_X1 us23_U201 (.A( us23_n749 ) , .ZN( us23_n841 ) );
  NOR2_X1 us23_U202 (.ZN( us23_n651 ) , .A1( us23_n668 ) , .A2( us23_n813 ) );
  NOR2_X1 us23_U203 (.ZN( us23_n531 ) , .A2( us23_n748 ) , .A1( us23_n749 ) );
  NOR2_X1 us23_U204 (.ZN( us23_n576 ) , .A2( us23_n698 ) , .A1( us23_n813 ) );
  NOR2_X1 us23_U205 (.ZN( us23_n599 ) , .A2( us23_n696 ) , .A1( us23_n783 ) );
  NOR2_X1 us23_U206 (.A1( us23_n668 ) , .ZN( us23_n672 ) , .A2( us23_n743 ) );
  NOR2_X1 us23_U207 (.ZN( us23_n601 ) , .A1( us23_n668 ) , .A2( us23_n802 ) );
  NOR2_X1 us23_U208 (.A1( us23_n668 ) , .ZN( us23_n687 ) , .A2( us23_n815 ) );
  NOR2_X1 us23_U209 (.ZN( us23_n628 ) , .A2( us23_n727 ) , .A1( us23_n784 ) );
  NOR4_X1 us23_U21 (.A4( us23_n540 ) , .A3( us23_n541 ) , .A2( us23_n542 ) , .ZN( us23_n549 ) , .A1( us23_n687 ) );
  NOR2_X1 us23_U210 (.ZN( us23_n614 ) , .A1( us23_n784 ) , .A2( us23_n814 ) );
  NOR2_X1 us23_U211 (.A2( us23_n743 ) , .ZN( us23_n754 ) , .A1( us23_n804 ) );
  NOR2_X1 us23_U212 (.A1( us23_n668 ) , .ZN( us23_n765 ) , .A2( us23_n812 ) );
  NOR2_X1 us23_U213 (.ZN( us23_n734 ) , .A2( us23_n802 ) , .A1( us23_n804 ) );
  NOR2_X1 us23_U214 (.A1( us23_n698 ) , .ZN( us23_n767 ) , .A2( us23_n812 ) );
  NOR2_X1 us23_U215 (.A2( us23_n743 ) , .ZN( us23_n768 ) , .A1( us23_n811 ) );
  NOR2_X1 us23_U216 (.ZN( us23_n530 ) , .A2( us23_n779 ) , .A1( us23_n815 ) );
  NOR2_X1 us23_U217 (.ZN( us23_n526 ) , .A1( us23_n668 ) , .A2( us23_n778 ) );
  NOR2_X1 us23_U218 (.ZN( us23_n540 ) , .A2( us23_n696 ) , .A1( us23_n698 ) );
  NOR2_X1 us23_U219 (.ZN( us23_n598 ) , .A2( us23_n790 ) , .A1( us23_n815 ) );
  NOR2_X1 us23_U22 (.ZN( us23_n679 ) , .A2( us23_n833 ) , .A1( us23_n838 ) );
  NOR2_X1 us23_U220 (.ZN( us23_n627 ) , .A2( us23_n668 ) , .A1( us23_n784 ) );
  NOR2_X1 us23_U221 (.ZN( us23_n600 ) , .A2( us23_n779 ) , .A1( us23_n802 ) );
  INV_X1 us23_U222 (.A( us23_n746 ) , .ZN( us23_n833 ) );
  NOR2_X1 us23_U223 (.ZN( us23_n610 ) , .A2( us23_n779 ) , .A1( us23_n805 ) );
  NOR2_X1 us23_U224 (.ZN( us23_n527 ) , .A2( us23_n723 ) , .A1( us23_n802 ) );
  NOR2_X1 us23_U225 (.ZN( us23_n609 ) , .A1( us23_n783 ) , .A2( us23_n815 ) );
  INV_X1 us23_U226 (.A( us23_n791 ) , .ZN( us23_n850 ) );
  NOR2_X1 us23_U227 (.ZN( us23_n650 ) , .A1( us23_n783 ) , .A2( us23_n787 ) );
  NOR2_X1 us23_U228 (.A2( us23_n707 ) , .A1( us23_n749 ) , .ZN( us23_n770 ) );
  NOR2_X1 us23_U229 (.ZN( us23_n666 ) , .A1( us23_n749 ) , .A2( us23_n814 ) );
  AOI222_X1 us23_U23 (.ZN( us23_n468 ) , .B1( us23_n831 ) , .A1( us23_n838 ) , .C1( us23_n841 ) , .C2( us23_n850 ) , .A2( us23_n854 ) , .B2( us23_n864 ) );
  NOR2_X1 us23_U230 (.ZN( us23_n554 ) , .A1( us23_n749 ) , .A2( us23_n790 ) );
  NOR2_X1 us23_U231 (.ZN( us23_n507 ) , .A2( us23_n779 ) , .A1( us23_n784 ) );
  NOR2_X1 us23_U232 (.ZN( us23_n542 ) , .A2( us23_n707 ) , .A1( us23_n784 ) );
  NOR2_X1 us23_U233 (.ZN( us23_n663 ) , .A1( us23_n784 ) , .A2( us23_n790 ) );
  OAI22_X1 us23_U234 (.B1( us23_n439 ) , .ZN( us23_n443 ) , .A2( us23_n727 ) , .A1( us23_n743 ) , .B2( us23_n748 ) );
  NOR3_X1 us23_U235 (.ZN( us23_n439 ) , .A2( us23_n835 ) , .A3( us23_n836 ) , .A1( us23_n845 ) );
  NOR2_X1 us23_U236 (.A2( us23_n696 ) , .ZN( us23_n715 ) , .A1( us23_n791 ) );
  NOR2_X1 us23_U237 (.ZN( us23_n506 ) , .A1( us23_n811 ) , .A2( us23_n816 ) );
  NOR2_X1 us23_U238 (.ZN( us23_n593 ) , .A2( us23_n696 ) , .A1( us23_n727 ) );
  NOR2_X1 us23_U239 (.ZN( us23_n661 ) , .A2( us23_n696 ) , .A1( us23_n728 ) );
  NOR4_X1 us23_U24 (.A1( us23_n465 ) , .ZN( us23_n466 ) , .A4( us23_n541 ) , .A2( us23_n553 ) , .A3( us23_n613 ) );
  NOR2_X1 us23_U240 (.ZN( us23_n556 ) , .A1( us23_n791 ) , .A2( us23_n813 ) );
  NOR2_X1 us23_U241 (.ZN( us23_n544 ) , .A1( us23_n748 ) , .A2( us23_n813 ) );
  NOR2_X1 us23_U242 (.ZN( us23_n555 ) , .A1( us23_n761 ) , .A2( us23_n804 ) );
  NOR2_X1 us23_U243 (.ZN( us23_n529 ) , .A2( us23_n743 ) , .A1( us23_n791 ) );
  NOR2_X1 us23_U244 (.A2( us23_n696 ) , .A1( us23_n779 ) , .ZN( us23_n819 ) );
  NOR2_X1 us23_U245 (.ZN( us23_n508 ) , .A1( us23_n728 ) , .A2( us23_n778 ) );
  NOR2_X1 us23_U246 (.ZN( us23_n665 ) , .A1( us23_n727 ) , .A2( us23_n802 ) );
  NOR2_X1 us23_U247 (.ZN( us23_n543 ) , .A2( us23_n784 ) , .A1( us23_n791 ) );
  NOR2_X1 us23_U248 (.A1( us23_n748 ) , .ZN( us23_n766 ) , .A2( us23_n802 ) );
  NOR2_X1 us23_U249 (.ZN( us23_n613 ) , .A1( us23_n761 ) , .A2( us23_n811 ) );
  AOI221_X1 us23_U25 (.ZN( us23_n467 ) , .C2( us23_n713 ) , .B2( us23_n830 ) , .C1( us23_n844 ) , .B1( us23_n859 ) , .A( us23_n863 ) );
  NOR2_X1 us23_U250 (.ZN( us23_n515 ) , .A1( us23_n707 ) , .A2( us23_n743 ) );
  NOR2_X1 us23_U251 (.ZN( us23_n630 ) , .A1( us23_n723 ) , .A2( us23_n812 ) );
  NOR2_X1 us23_U252 (.ZN( us23_n569 ) , .A1( us23_n727 ) , .A2( us23_n805 ) );
  NOR2_X1 us23_U253 (.ZN( us23_n557 ) , .A1( us23_n707 ) , .A2( us23_n815 ) );
  INV_X1 us23_U254 (.A( us23_n762 ) , .ZN( us23_n865 ) );
  NOR2_X1 us23_U255 (.ZN( us23_n653 ) , .A1( us23_n727 ) , .A2( us23_n812 ) );
  NOR2_X1 us23_U256 (.ZN( us23_n516 ) , .A1( us23_n707 ) , .A2( us23_n802 ) );
  NOR2_X1 us23_U257 (.ZN( us23_n520 ) , .A1( us23_n789 ) , .A2( us23_n811 ) );
  NOR2_X1 us23_U258 (.ZN( us23_n662 ) , .A1( us23_n728 ) , .A2( us23_n784 ) );
  NOR2_X1 us23_U259 (.ZN( us23_n654 ) , .A1( us23_n789 ) , .A2( us23_n814 ) );
  NOR4_X1 us23_U26 (.A4( us23_n664 ) , .A3( us23_n665 ) , .A2( us23_n666 ) , .A1( us23_n667 ) , .ZN( us23_n675 ) );
  NOR2_X1 us23_U260 (.ZN( us23_n629 ) , .A1( us23_n746 ) , .A2( us23_n814 ) );
  NOR2_X1 us23_U261 (.ZN( us23_n667 ) , .A2( us23_n707 ) , .A1( us23_n789 ) );
  NOR2_X1 us23_U262 (.ZN( us23_n669 ) , .A1( us23_n789 ) , .A2( us23_n804 ) );
  AOI21_X1 us23_U263 (.ZN( us23_n570 ) , .B2( us23_n696 ) , .B1( us23_n805 ) , .A( us23_n811 ) );
  NOR2_X1 us23_U264 (.ZN( us23_n541 ) , .A1( us23_n761 ) , .A2( us23_n790 ) );
  NOR2_X1 us23_U265 (.ZN( us23_n655 ) , .A1( us23_n746 ) , .A2( us23_n779 ) );
  INV_X1 us23_U266 (.A( us23_n805 ) , .ZN( us23_n840 ) );
  NOR2_X1 us23_U267 (.ZN( us23_n608 ) , .A2( us23_n723 ) , .A1( us23_n816 ) );
  AOI21_X1 us23_U268 (.A( us23_n814 ) , .B2( us23_n815 ) , .B1( us23_n816 ) , .ZN( us23_n817 ) );
  AOI21_X1 us23_U269 (.ZN( us23_n625 ) , .B2( us23_n668 ) , .A( us23_n789 ) , .B1( us23_n790 ) );
  NOR4_X1 us23_U27 (.A4( us23_n660 ) , .A3( us23_n661 ) , .A2( us23_n662 ) , .A1( us23_n663 ) , .ZN( us23_n676 ) );
  NOR2_X1 us23_U270 (.ZN( us23_n660 ) , .A1( us23_n728 ) , .A2( us23_n789 ) );
  INV_X1 us23_U271 (.A( us23_n811 ) , .ZN( us23_n853 ) );
  NOR2_X1 us23_U272 (.ZN( us23_n578 ) , .A2( us23_n707 ) , .A1( us23_n729 ) );
  NOR2_X1 us23_U273 (.ZN( us23_n532 ) , .A2( us23_n723 ) , .A1( us23_n729 ) );
  AOI21_X1 us23_U274 (.ZN( us23_n498 ) , .B1( us23_n679 ) , .A( us23_n811 ) , .B2( us23_n815 ) );
  AOI21_X1 us23_U275 (.ZN( us23_n551 ) , .B1( us23_n668 ) , .A( us23_n696 ) , .B2( us23_n804 ) );
  NOR2_X1 us23_U276 (.ZN( us23_n581 ) , .A1( us23_n743 ) , .A2( us23_n814 ) );
  NOR2_X1 us23_U277 (.A2( us23_n707 ) , .A1( us23_n761 ) , .ZN( us23_n793 ) );
  AOI21_X1 us23_U278 (.B1( us23_n624 ) , .ZN( us23_n626 ) , .A( us23_n762 ) , .B2( us23_n813 ) );
  AOI21_X1 us23_U279 (.ZN( us23_n514 ) , .A( us23_n728 ) , .B1( us23_n749 ) , .B2( us23_n802 ) );
  NOR4_X1 us23_U28 (.A3( us23_n672 ) , .A1( us23_n673 ) , .ZN( us23_n674 ) , .A4( us23_n714 ) , .A2( us23_n858 ) );
  AOI21_X1 us23_U280 (.A( us23_n811 ) , .B2( us23_n812 ) , .B1( us23_n813 ) , .ZN( us23_n818 ) );
  AOI21_X1 us23_U281 (.ZN( us23_n477 ) , .B2( us23_n696 ) , .A( us23_n748 ) , .B1( us23_n778 ) );
  AOI21_X1 us23_U282 (.ZN( us23_n509 ) , .B2( us23_n668 ) , .A( us23_n729 ) , .B1( us23_n814 ) );
  NOR2_X1 us23_U283 (.ZN( us23_n505 ) , .A2( us23_n727 ) , .A1( us23_n761 ) );
  AOI21_X1 us23_U284 (.ZN( us23_n591 ) , .B1( us23_n727 ) , .B2( us23_n783 ) , .A( us23_n789 ) );
  NOR2_X1 us23_U285 (.ZN( us23_n518 ) , .A2( us23_n698 ) , .A1( us23_n815 ) );
  AOI21_X1 us23_U286 (.ZN( us23_n592 ) , .B1( us23_n749 ) , .A( us23_n791 ) , .B2( us23_n812 ) );
  AOI21_X1 us23_U287 (.ZN( us23_n649 ) , .A( us23_n778 ) , .B1( us23_n791 ) , .B2( us23_n804 ) );
  NOR2_X1 us23_U288 (.ZN( us23_n580 ) , .A1( us23_n668 ) , .A2( us23_n787 ) );
  NOR2_X1 us23_U289 (.ZN( us23_n519 ) , .A2( us23_n707 ) , .A1( us23_n813 ) );
  NOR4_X1 us23_U29 (.A4( us23_n513 ) , .A3( us23_n514 ) , .A2( us23_n515 ) , .A1( us23_n516 ) , .ZN( us23_n523 ) );
  AOI21_X1 us23_U290 (.ZN( us23_n476 ) , .A( us23_n668 ) , .B1( us23_n749 ) , .B2( us23_n805 ) );
  NOR2_X1 us23_U291 (.ZN( us23_n558 ) , .A2( us23_n790 ) , .A1( us23_n802 ) );
  AOI21_X1 us23_U292 (.ZN( us23_n647 ) , .A( us23_n761 ) , .B2( us23_n783 ) , .B1( us23_n791 ) );
  AOI21_X1 us23_U293 (.ZN( us23_n622 ) , .B1( us23_n698 ) , .A( us23_n778 ) , .B2( us23_n783 ) );
  AOI21_X1 us23_U294 (.ZN( us23_n588 ) , .B2( us23_n698 ) , .B1( us23_n814 ) , .A( us23_n816 ) );
  NOR2_X1 us23_U295 (.ZN( us23_n552 ) , .A2( us23_n743 ) , .A1( us23_n783 ) );
  NOR2_X1 us23_U296 (.ZN( us23_n682 ) , .A2( us23_n698 ) , .A1( us23_n802 ) );
  AOI21_X1 us23_U297 (.B1( us23_n698 ) , .ZN( us23_n699 ) , .A( us23_n731 ) , .B2( us23_n762 ) );
  AOI21_X1 us23_U298 (.ZN( us23_n590 ) , .B2( us23_n762 ) , .A( us23_n784 ) , .B1( us23_n811 ) );
  AOI21_X1 us23_U299 (.ZN( us23_n538 ) , .B2( us23_n811 ) , .A( us23_n813 ) , .B1( us23_n814 ) );
  NOR3_X1 us23_U3 (.ZN( us23_n597 ) , .A1( us23_n607 ) , .A3( us23_n722 ) , .A2( us23_n741 ) );
  AOI222_X1 us23_U30 (.ZN( us23_n524 ) , .A1( us23_n833 ) , .B2( us23_n836 ) , .C1( us23_n843 ) , .C2( us23_n849 ) , .A2( us23_n851 ) , .B1( us23_n865 ) );
  AOI21_X1 us23_U300 (.ZN( us23_n539 ) , .A( us23_n762 ) , .B2( us23_n778 ) , .B1( us23_n816 ) );
  NOR2_X1 us23_U301 (.ZN( us23_n546 ) , .A1( us23_n698 ) , .A2( us23_n743 ) );
  INV_X1 us23_U302 (.A( us23_n812 ) , .ZN( us23_n835 ) );
  INV_X1 us23_U303 (.A( us23_n727 ) , .ZN( us23_n851 ) );
  AOI21_X1 us23_U304 (.ZN( us23_n648 ) , .B1( us23_n728 ) , .B2( us23_n762 ) , .A( us23_n812 ) );
  INV_X1 us23_U305 (.A( us23_n790 ) , .ZN( us23_n872 ) );
  OAI221_X1 us23_U306 (.A( us23_n726 ) , .C2( us23_n727 ) , .B2( us23_n728 ) , .B1( us23_n729 ) , .ZN( us23_n736 ) , .C1( us23_n816 ) );
  AOI22_X1 us23_U307 (.ZN( us23_n726 ) , .B1( us23_n831 ) , .A2( us23_n837 ) , .A1( us23_n862 ) , .B2( us23_n865 ) );
  AOI21_X1 us23_U308 (.ZN( us23_n497 ) , .A( us23_n723 ) , .B2( us23_n761 ) , .B1( us23_n813 ) );
  NOR2_X1 us23_U309 (.ZN( us23_n565 ) , .A2( us23_n696 ) , .A1( us23_n762 ) );
  NOR4_X1 us23_U31 (.A3( us23_n520 ) , .A1( us23_n521 ) , .ZN( us23_n522 ) , .A2( us23_n672 ) , .A4( us23_n768 ) );
  INV_X1 us23_U310 (.A( us23_n698 ) , .ZN( us23_n852 ) );
  AOI21_X1 us23_U311 (.ZN( us23_n568 ) , .B1( us23_n749 ) , .B2( us23_n761 ) , .A( us23_n779 ) );
  AOI21_X1 us23_U312 (.ZN( us23_n513 ) , .A( us23_n778 ) , .B2( us23_n791 ) , .B1( us23_n811 ) );
  NOR2_X1 us23_U313 (.ZN( us23_n579 ) , .A2( us23_n696 ) , .A1( us23_n790 ) );
  NOR2_X1 us23_U314 (.ZN( us23_n684 ) , .A1( us23_n728 ) , .A2( us23_n815 ) );
  AOI21_X1 us23_U315 (.ZN( us23_n563 ) , .B1( us23_n723 ) , .A( us23_n778 ) , .B2( us23_n790 ) );
  AOI21_X1 us23_U316 (.ZN( us23_n496 ) , .A( us23_n778 ) , .B2( us23_n790 ) , .B1( us23_n803 ) );
  INV_X1 us23_U317 (.A( us23_n728 ) , .ZN( us23_n867 ) );
  NOR2_X1 us23_U318 (.ZN( us23_n664 ) , .A1( us23_n779 ) , .A2( us23_n812 ) );
  NOR2_X1 us23_U319 (.ZN( us23_n631 ) , .A2( us23_n696 ) , .A1( us23_n723 ) );
  AOI221_X1 us23_U32 (.A( us23_n780 ) , .ZN( us23_n797 ) , .C2( us23_n836 ) , .B2( us23_n837 ) , .B1( us23_n864 ) , .C1( us23_n865 ) );
  NOR2_X1 us23_U320 (.ZN( us23_n528 ) , .A1( us23_n707 ) , .A2( us23_n778 ) );
  NOR2_X1 us23_U321 (.ZN( us23_n577 ) , .A1( us23_n707 ) , .A2( us23_n812 ) );
  AOI21_X1 us23_U322 (.A( us23_n789 ) , .B2( us23_n790 ) , .B1( us23_n791 ) , .ZN( us23_n792 ) );
  AOI21_X1 us23_U323 (.ZN( us23_n688 ) , .B2( us23_n748 ) , .B1( us23_n762 ) , .A( us23_n805 ) );
  NOR2_X1 us23_U324 (.ZN( us23_n683 ) , .A1( us23_n790 ) , .A2( us23_n812 ) );
  NOR2_X1 us23_U325 (.ZN( us23_n566 ) , .A1( us23_n746 ) , .A2( us23_n804 ) );
  NAND2_X1 us23_U326 (.ZN( us23_n752 ) , .A1( us23_n762 ) , .A2( us23_n804 ) );
  AOI21_X1 us23_U327 (.A( us23_n732 ) , .ZN( us23_n733 ) , .B2( us23_n779 ) , .B1( us23_n791 ) );
  NOR2_X1 us23_U328 (.A2( us23_n812 ) , .A1( us23_n814 ) , .ZN( us23_n820 ) );
  NOR2_X1 us23_U329 (.ZN( us23_n710 ) , .A1( us23_n761 ) , .A2( us23_n762 ) );
  NOR4_X1 us23_U33 (.A4( us23_n792 ) , .A3( us23_n793 ) , .A2( us23_n794 ) , .A1( us23_n795 ) , .ZN( us23_n796 ) );
  NOR2_X1 us23_U330 (.ZN( us23_n641 ) , .A2( us23_n787 ) , .A1( us23_n790 ) );
  NOR2_X1 us23_U331 (.ZN( us23_n582 ) , .A1( us23_n791 ) , .A2( us23_n816 ) );
  NOR2_X1 us23_U332 (.ZN( us23_n681 ) , .A2( us23_n707 ) , .A1( us23_n816 ) );
  NOR2_X1 us23_U333 (.ZN( us23_n533 ) , .A1( us23_n723 ) , .A2( us23_n787 ) );
  AOI21_X1 us23_U334 (.B1( us23_n685 ) , .ZN( us23_n686 ) , .A( us23_n727 ) , .B2( us23_n760 ) );
  INV_X1 us23_U335 (.A( us23_n696 ) , .ZN( us23_n837 ) );
  INV_X1 us23_U336 (.A( us23_n814 ) , .ZN( us23_n854 ) );
  NOR2_X1 us23_U337 (.ZN( us23_n567 ) , .A1( us23_n728 ) , .A2( us23_n761 ) );
  AOI21_X1 us23_U338 (.ZN( us23_n441 ) , .A( us23_n698 ) , .B1( us23_n732 ) , .B2( us23_n749 ) );
  OAI21_X1 us23_U339 (.A( us23_n730 ) , .B1( us23_n731 ) , .ZN( us23_n735 ) , .B2( us23_n804 ) );
  NOR4_X1 us23_U34 (.A4( us23_n775 ) , .A3( us23_n776 ) , .A1( us23_n777 ) , .ZN( us23_n798 ) , .A2( us23_n800 ) );
  OAI21_X1 us23_U340 (.ZN( us23_n730 ) , .A( us23_n832 ) , .B2( us23_n851 ) , .B1( us23_n872 ) );
  OAI21_X1 us23_U341 (.A( us23_n697 ) , .ZN( us23_n701 ) , .B2( us23_n749 ) , .B1( us23_n803 ) );
  OAI21_X1 us23_U342 (.ZN( us23_n697 ) , .B2( us23_n832 ) , .B1( us23_n837 ) , .A( us23_n859 ) );
  OAI21_X1 us23_U343 (.A( us23_n612 ) , .ZN( us23_n615 ) , .B1( us23_n624 ) , .B2( us23_n783 ) );
  INV_X1 us23_U344 (.A( us23_n779 ) , .ZN( us23_n849 ) );
  AOI22_X1 us23_U345 (.A2( us23_n781 ) , .ZN( us23_n782 ) , .B2( us23_n830 ) , .A1( us23_n833 ) , .B1( us23_n862 ) );
  NAND2_X1 us23_U346 (.ZN( us23_n670 ) , .A1( us23_n805 ) , .A2( us23_n815 ) );
  OAI21_X1 us23_U347 (.A( us23_n786 ) , .B2( us23_n787 ) , .B1( us23_n788 ) , .ZN( us23_n794 ) );
  OAI21_X1 us23_U348 (.ZN( us23_n786 ) , .A( us23_n838 ) , .B1( us23_n862 ) , .B2( us23_n872 ) );
  NAND2_X1 us23_U349 (.A1( us23_n728 ) , .A2( us23_n783 ) , .ZN( us23_n810 ) );
  NOR4_X1 us23_U35 (.A4( us23_n733 ) , .A3( us23_n734 ) , .A2( us23_n735 ) , .A1( us23_n736 ) , .ZN( us23_n737 ) );
  NOR2_X1 us23_U350 (.ZN( us23_n483 ) , .A1( us23_n787 ) , .A2( us23_n804 ) );
  AOI21_X1 us23_U351 (.ZN( us23_n442 ) , .B1( us23_n788 ) , .B2( us23_n790 ) , .A( us23_n813 ) );
  NAND2_X1 us23_U352 (.A2( us23_n761 ) , .A1( us23_n805 ) , .ZN( us23_n809 ) );
  NOR2_X1 us23_U353 (.ZN( us23_n469 ) , .A2( us23_n778 ) , .A1( us23_n814 ) );
  NAND2_X1 us23_U354 (.A1( us23_n698 ) , .A2( us23_n728 ) , .ZN( us23_n781 ) );
  NOR2_X1 us23_U355 (.ZN( us23_n711 ) , .A2( us23_n723 ) , .A1( us23_n789 ) );
  INV_X1 us23_U356 (.A( us23_n784 ) , .ZN( us23_n845 ) );
  NOR2_X1 us23_U357 (.ZN( us23_n525 ) , .A1( us23_n723 ) , .A2( us23_n749 ) );
  NOR2_X1 us23_U358 (.ZN( us23_n517 ) , .A1( us23_n707 ) , .A2( us23_n787 ) );
  INV_X1 us23_U359 (.A( us23_n816 ) , .ZN( us23_n843 ) );
  AOI211_X1 us23_U36 (.B( us23_n724 ) , .A( us23_n725 ) , .ZN( us23_n738 ) , .C1( us23_n842 ) , .C2( us23_n854 ) );
  NAND2_X1 us23_U360 (.ZN( us23_n713 ) , .A1( us23_n727 ) , .A2( us23_n779 ) );
  INV_X1 us23_U361 (.A( us23_n723 ) , .ZN( us23_n855 ) );
  AND2_X1 us23_U362 (.ZN( us23_n731 ) , .A1( us23_n778 ) , .A2( us23_n784 ) );
  NAND2_X1 us23_U363 (.A2( us23_n460 ) , .A1( us23_n470 ) , .ZN( us23_n696 ) );
  NAND2_X1 us23_U364 (.A1( us23_n451 ) , .A2( us23_n464 ) , .ZN( us23_n668 ) );
  NAND2_X1 us23_U365 (.A1( us23_n450 ) , .A2( us23_n470 ) , .ZN( us23_n815 ) );
  NAND2_X1 us23_U366 (.A1( us23_n452 ) , .A2( us23_n460 ) , .ZN( us23_n743 ) );
  NAND2_X1 us23_U367 (.A1( us23_n454 ) , .A2( us23_n470 ) , .ZN( us23_n802 ) );
  NAND2_X1 us23_U368 (.A1( us23_n450 ) , .A2( us23_n453 ) , .ZN( us23_n813 ) );
  NAND2_X1 us23_U369 (.A1( us23_n454 ) , .A2( us23_n461 ) , .ZN( us23_n749 ) );
  NOR3_X1 us23_U37 (.A3( us23_n721 ) , .A1( us23_n722 ) , .ZN( us23_n739 ) , .A2( us23_n740 ) );
  NAND2_X1 us23_U370 (.A1( us23_n446 ) , .A2( us23_n448 ) , .ZN( us23_n804 ) );
  NAND2_X1 us23_U371 (.A1( us23_n453 ) , .A2( us23_n460 ) , .ZN( us23_n812 ) );
  NAND2_X1 us23_U372 (.A2( us23_n440 ) , .A1( us23_n446 ) , .ZN( us23_n783 ) );
  NAND2_X1 us23_U373 (.A2( us23_n453 ) , .A1( us23_n471 ) , .ZN( us23_n778 ) );
  NAND2_X1 us23_U374 (.A2( us23_n452 ) , .A1( us23_n454 ) , .ZN( us23_n805 ) );
  NAND2_X1 us23_U375 (.A1( us23_n452 ) , .A2( us23_n471 ) , .ZN( us23_n784 ) );
  NAND2_X1 us23_U376 (.A1( us23_n440 ) , .A2( us23_n459 ) , .ZN( us23_n698 ) );
  NAND2_X1 us23_U377 (.A2( us23_n463 ) , .A1( us23_n464 ) , .ZN( us23_n811 ) );
  NAND2_X1 us23_U378 (.A2( us23_n448 ) , .A1( us23_n451 ) , .ZN( us23_n762 ) );
  NAND2_X1 us23_U379 (.A1( us23_n461 ) , .A2( us23_n471 ) , .ZN( us23_n787 ) );
  NOR4_X1 us23_U38 (.A3( us23_n754 ) , .A2( us23_n755 ) , .A1( us23_n756 ) , .ZN( us23_n757 ) , .A4( us23_n868 ) );
  NAND2_X1 us23_U380 (.A2( us23_n460 ) , .A1( us23_n461 ) , .ZN( us23_n746 ) );
  NOR2_X1 us23_U381 (.ZN( us23_n464 ) , .A2( us23_n846 ) , .A1( us23_n847 ) );
  NOR2_X1 us23_U382 (.ZN( us23_n452 ) , .A1( us23_n825 ) , .A2( us23_n826 ) );
  NAND2_X1 us23_U383 (.A1( us23_n450 ) , .A2( us23_n461 ) , .ZN( us23_n789 ) );
  NOR2_X1 us23_U384 (.ZN( us23_n450 ) , .A1( us23_n827 ) , .A2( us23_n828 ) );
  NAND2_X2 us23_U385 (.A2( us23_n447 ) , .A1( us23_n463 ) , .ZN( us23_n814 ) );
  NAND2_X1 us23_U386 (.A2( us23_n453 ) , .A1( us23_n454 ) , .ZN( us23_n729 ) );
  NAND2_X2 us23_U387 (.A2( us23_n440 ) , .A1( us23_n451 ) , .ZN( us23_n790 ) );
  NAND2_X2 us23_U388 (.A1( us23_n448 ) , .A2( us23_n459 ) , .ZN( us23_n791 ) );
  NAND2_X2 us23_U389 (.A1( us23_n448 ) , .A2( us23_n463 ) , .ZN( us23_n723 ) );
  AOI211_X1 us23_U39 (.B( us23_n744 ) , .A( us23_n745 ) , .ZN( us23_n758 ) , .C1( us23_n831 ) , .C2( us23_n852 ) );
  NAND2_X2 us23_U390 (.A1( us23_n440 ) , .A2( us23_n463 ) , .ZN( us23_n707 ) );
  NAND2_X2 us23_U391 (.A2( us23_n470 ) , .A1( us23_n471 ) , .ZN( us23_n816 ) );
  NAND2_X2 us23_U392 (.A2( us23_n459 ) , .A1( us23_n464 ) , .ZN( us23_n779 ) );
  NOR2_X1 us23_U393 (.ZN( us23_n446 ) , .A2( us23_n848 ) , .A1( us23_n857 ) );
  NAND2_X1 us23_U394 (.A1( us23_n446 ) , .A2( us23_n447 ) , .ZN( us23_n785 ) );
  NAND2_X1 us23_U395 (.A2( us23_n447 ) , .A1( us23_n459 ) , .ZN( us23_n727 ) );
  NAND2_X1 us23_U396 (.A2( us23_n447 ) , .A1( us23_n451 ) , .ZN( us23_n728 ) );
  NOR2_X1 us23_U397 (.A2( sa23_5 ) , .ZN( us23_n447 ) , .A1( us23_n846 ) );
  NOR2_X1 us23_U398 (.A2( sa23_7 ) , .ZN( us23_n459 ) , .A1( us23_n848 ) );
  NOR2_X1 us23_U399 (.A2( sa23_6 ) , .A1( sa23_7 ) , .ZN( us23_n463 ) );
  NOR3_X1 us23_U4 (.A3( us23_n799 ) , .A2( us23_n800 ) , .A1( us23_n801 ) , .ZN( us23_n824 ) );
  NOR3_X1 us23_U40 (.A3( us23_n740 ) , .A2( us23_n741 ) , .A1( us23_n742 ) , .ZN( us23_n759 ) );
  NOR2_X1 us23_U400 (.A2( sa23_4 ) , .ZN( us23_n448 ) , .A1( us23_n847 ) );
  NOR2_X1 us23_U401 (.A2( sa23_4 ) , .A1( sa23_5 ) , .ZN( us23_n440 ) );
  NOR2_X1 us23_U402 (.A2( sa23_6 ) , .ZN( us23_n451 ) , .A1( us23_n857 ) );
  NOR2_X1 us23_U403 (.A2( sa23_1 ) , .ZN( us23_n470 ) , .A1( us23_n825 ) );
  NOR2_X1 us23_U404 (.A2( sa23_2 ) , .A1( sa23_3 ) , .ZN( us23_n471 ) );
  NOR2_X1 us23_U405 (.A2( sa23_2 ) , .ZN( us23_n460 ) , .A1( us23_n828 ) );
  NOR2_X1 us23_U406 (.A2( sa23_0 ) , .ZN( us23_n453 ) , .A1( us23_n826 ) );
  NOR2_X1 us23_U407 (.A2( sa23_0 ) , .A1( sa23_1 ) , .ZN( us23_n461 ) );
  NOR2_X1 us23_U408 (.A2( sa23_3 ) , .ZN( us23_n454 ) , .A1( us23_n827 ) );
  INV_X1 us23_U409 (.A( sa23_6 ) , .ZN( us23_n848 ) );
  NAND4_X1 us23_U41 (.ZN( sa21_sr_3 ) , .A4( us23_n703 ) , .A3( us23_n704 ) , .A2( us23_n705 ) , .A1( us23_n706 ) );
  INV_X1 us23_U410 (.A( sa23_4 ) , .ZN( us23_n846 ) );
  INV_X1 us23_U411 (.A( sa23_1 ) , .ZN( us23_n826 ) );
  INV_X1 us23_U412 (.A( sa23_3 ) , .ZN( us23_n828 ) );
  INV_X1 us23_U413 (.A( sa23_2 ) , .ZN( us23_n827 ) );
  INV_X1 us23_U414 (.A( sa23_0 ) , .ZN( us23_n825 ) );
  INV_X1 us23_U415 (.A( sa23_7 ) , .ZN( us23_n857 ) );
  INV_X1 us23_U416 (.A( sa23_5 ) , .ZN( us23_n847 ) );
  OAI221_X1 us23_U417 (.A( us23_n782 ) , .C2( us23_n783 ) , .B2( us23_n784 ) , .B1( us23_n785 ) , .ZN( us23_n795 ) , .C1( us23_n812 ) );
  OAI222_X1 us23_U418 (.B2( us23_n746 ) , .B1( us23_n747 ) , .A2( us23_n748 ) , .ZN( us23_n756 ) , .C2( us23_n804 ) , .C1( us23_n813 ) , .A1( us23_n816 ) );
  AOI21_X1 us23_U419 (.ZN( us23_n499 ) , .A( us23_n696 ) , .B1( us23_n707 ) , .B2( us23_n785 ) );
  NOR4_X1 us23_U42 (.A4( us23_n699 ) , .A3( us23_n700 ) , .A2( us23_n701 ) , .A1( us23_n702 ) , .ZN( us23_n703 ) );
  OAI221_X1 us23_U420 (.A( us23_n695 ) , .ZN( us23_n702 ) , .C2( us23_n783 ) , .C1( us23_n784 ) , .B1( us23_n785 ) , .B2( us23_n805 ) );
  OAI22_X1 us23_U421 (.ZN( us23_n589 ) , .B1( us23_n729 ) , .B2( us23_n748 ) , .A2( us23_n785 ) , .A1( us23_n802 ) );
  OAI222_X1 us23_U422 (.ZN( us23_n504 ) , .C2( us23_n624 ) , .B2( us23_n646 ) , .B1( us23_n746 ) , .A2( us23_n747 ) , .C1( us23_n804 ) , .A1( us23_n805 ) );
  NOR2_X1 us23_U423 (.ZN( us23_n611 ) , .A1( us23_n778 ) , .A2( us23_n785 ) );
  OAI222_X1 us23_U424 (.ZN( us23_n616 ) , .B1( us23_n696 ) , .C1( us23_n723 ) , .C2( us23_n746 ) , .B2( us23_n785 ) , .A2( us23_n791 ) , .A1( us23_n815 ) );
  NAND2_X1 us23_U425 (.A2( us23_n748 ) , .A1( us23_n785 ) , .ZN( us23_n808 ) );
  AOI21_X1 us23_U426 (.ZN( us23_n575 ) , .B2( us23_n723 ) , .B1( us23_n747 ) , .A( us23_n784 ) );
  NOR2_X1 us23_U427 (.ZN( us23_n716 ) , .A2( us23_n743 ) , .A1( us23_n785 ) );
  NOR2_X1 us23_U428 (.ZN( us23_n652 ) , .A1( us23_n761 ) , .A2( us23_n785 ) );
  NOR2_X1 us23_U429 (.ZN( us23_n553 ) , .A1( us23_n785 ) , .A2( us23_n812 ) );
  AOI211_X1 us23_U43 (.B( us23_n693 ) , .A( us23_n694 ) , .ZN( us23_n704 ) , .C2( us23_n830 ) , .C1( us23_n850 ) );
  NOR2_X1 us23_U430 (.ZN( us23_n700 ) , .A2( us23_n785 ) , .A1( us23_n816 ) );
  NOR2_X1 us23_U431 (.A1( us23_n729 ) , .ZN( us23_n764 ) , .A2( us23_n785 ) );
  NAND2_X1 us23_U432 (.ZN( sa21_sr_2 ) , .A1( us23_n438 ) , .A2( us23_n644 ) );
  NOR3_X1 us23_U433 (.A2( us23_n606 ) , .A1( us23_n607 ) , .ZN( us23_n645 ) , .A3( us23_n721 ) );
  AOI222_X1 us23_U434 (.B2( us23_n637 ) , .ZN( us23_n643 ) , .B1( us23_n840 ) , .A1( us23_n841 ) , .C2( us23_n845 ) , .C1( us23_n862 ) , .A2( us23_n864 ) );
  NOR4_X1 us23_U435 (.A4( us23_n638 ) , .A3( us23_n639 ) , .A2( us23_n640 ) , .A1( us23_n641 ) , .ZN( us23_n642 ) );
  AOI211_X1 us23_U436 (.A( us23_n636 ) , .ZN( us23_n644 ) , .B( us23_n742 ) , .C2( us23_n838 ) , .C1( us23_n853 ) );
  NAND3_X1 us23_U437 (.ZN( sa21_sr_6 ) , .A3( us23_n796 ) , .A2( us23_n797 ) , .A1( us23_n798 ) );
  NAND3_X1 us23_U438 (.ZN( sa21_sr_5 ) , .A3( us23_n757 ) , .A2( us23_n758 ) , .A1( us23_n759 ) );
  NAND3_X1 us23_U439 (.ZN( sa21_sr_4 ) , .A3( us23_n737 ) , .A2( us23_n738 ) , .A1( us23_n739 ) );
  NOR2_X1 us23_U44 (.ZN( us23_n706 ) , .A2( us23_n775 ) , .A1( us23_n799 ) );
  NAND3_X1 us23_U440 (.A3( us23_n674 ) , .A2( us23_n675 ) , .A1( us23_n676 ) , .ZN( us23_n806 ) );
  NAND3_X1 us23_U441 (.ZN( us23_n637 ) , .A3( us23_n707 ) , .A2( us23_n723 ) , .A1( us23_n791 ) );
  NAND3_X1 us23_U442 (.A3( us23_n617 ) , .A2( us23_n618 ) , .A1( us23_n619 ) , .ZN( us23_n724 ) );
  NAND3_X1 us23_U443 (.A3( us23_n584 ) , .A2( us23_n585 ) , .A1( us23_n586 ) , .ZN( us23_n620 ) );
  NAND3_X1 us23_U444 (.ZN( us23_n564 ) , .A3( us23_n679 ) , .A2( us23_n749 ) , .A1( us23_n784 ) );
  NAND3_X1 us23_U445 (.A3( us23_n522 ) , .A2( us23_n523 ) , .A1( us23_n524 ) , .ZN( us23_n741 ) );
  NAND3_X1 us23_U446 (.A3( us23_n511 ) , .A1( us23_n512 ) , .ZN( us23_n607 ) , .A2( us23_n870 ) );
  NAND3_X1 us23_U447 (.A3( us23_n466 ) , .A2( us23_n467 ) , .A1( us23_n468 ) , .ZN( us23_n776 ) );
  NAND4_X1 us23_U448 (.A4( us23_n632 ) , .A3( us23_n633 ) , .A2( us23_n634 ) , .A1( us23_n635 ) , .ZN( us23_n742 ) );
  NOR2_X1 us23_U45 (.ZN( us23_n803 ) , .A1( us23_n853 ) , .A2( us23_n860 ) );
  NAND4_X1 us23_U46 (.ZN( sa21_sr_7 ) , .A4( us23_n821 ) , .A3( us23_n822 ) , .A2( us23_n823 ) , .A1( us23_n824 ) );
  AOI222_X1 us23_U47 (.C2( us23_n808 ) , .B2( us23_n809 ) , .A2( us23_n810 ) , .ZN( us23_n822 ) , .C1( us23_n831 ) , .A1( us23_n838 ) , .B1( us23_n852 ) );
  NOR4_X1 us23_U48 (.A4( us23_n817 ) , .A3( us23_n818 ) , .A2( us23_n819 ) , .A1( us23_n820 ) , .ZN( us23_n821 ) );
  AOI211_X1 us23_U49 (.B( us23_n806 ) , .A( us23_n807 ) , .ZN( us23_n823 ) , .C1( us23_n841 ) , .C2( us23_n849 ) );
  NOR3_X1 us23_U5 (.ZN( us23_n503 ) , .A2( us23_n678 ) , .A3( us23_n776 ) , .A1( us23_n875 ) );
  NAND4_X1 us23_U50 (.ZN( sa21_sr_0 ) , .A4( us23_n500 ) , .A3( us23_n501 ) , .A2( us23_n502 ) , .A1( us23_n503 ) );
  NOR4_X1 us23_U51 (.A4( us23_n497 ) , .A3( us23_n498 ) , .A2( us23_n499 ) , .ZN( us23_n500 ) , .A1( us23_n526 ) );
  AOI221_X1 us23_U52 (.A( us23_n496 ) , .ZN( us23_n501 ) , .B2( us23_n842 ) , .C1( us23_n845 ) , .C2( us23_n859 ) , .B1( us23_n861 ) );
  AOI211_X1 us23_U53 (.A( us23_n495 ) , .ZN( us23_n502 ) , .B( us23_n801 ) , .C2( us23_n838 ) , .C1( us23_n850 ) );
  AND3_X1 us23_U54 (.ZN( us23_n438 ) , .A2( us23_n642 ) , .A3( us23_n643 ) , .A1( us23_n645 ) );
  NAND4_X1 us23_U55 (.ZN( sa21_sr_1 ) , .A4( us23_n594 ) , .A3( us23_n595 ) , .A2( us23_n596 ) , .A1( us23_n597 ) );
  NOR4_X1 us23_U56 (.A4( us23_n590 ) , .A3( us23_n591 ) , .A2( us23_n592 ) , .A1( us23_n593 ) , .ZN( us23_n594 ) );
  AOI211_X1 us23_U57 (.B( us23_n588 ) , .A( us23_n589 ) , .ZN( us23_n595 ) , .C2( us23_n810 ) , .C1( us23_n832 ) );
  AOI211_X1 us23_U58 (.A( us23_n587 ) , .ZN( us23_n596 ) , .B( us23_n620 ) , .C1( us23_n844 ) , .C2( us23_n854 ) );
  NOR2_X1 us23_U59 (.ZN( us23_n624 ) , .A2( us23_n835 ) , .A1( us23_n838 ) );
  INV_X1 us23_U6 (.A( us23_n705 ) , .ZN( us23_n875 ) );
  NOR4_X1 us23_U60 (.A4( us23_n628 ) , .A3( us23_n629 ) , .A2( us23_n630 ) , .A1( us23_n631 ) , .ZN( us23_n632 ) );
  AOI211_X1 us23_U61 (.B( us23_n622 ) , .A( us23_n623 ) , .ZN( us23_n634 ) , .C2( us23_n835 ) , .C1( us23_n862 ) );
  NOR4_X1 us23_U62 (.A4( us23_n625 ) , .A3( us23_n626 ) , .A2( us23_n627 ) , .ZN( us23_n633 ) , .A1( us23_n663 ) );
  NAND4_X1 us23_U63 (.A4( us23_n656 ) , .A3( us23_n657 ) , .A2( us23_n658 ) , .A1( us23_n659 ) , .ZN( us23_n799 ) );
  NOR3_X1 us23_U64 (.A3( us23_n650 ) , .A2( us23_n651 ) , .A1( us23_n652 ) , .ZN( us23_n657 ) );
  NOR3_X1 us23_U65 (.A3( us23_n647 ) , .A2( us23_n648 ) , .A1( us23_n649 ) , .ZN( us23_n658 ) );
  NOR3_X1 us23_U66 (.A3( us23_n653 ) , .A2( us23_n654 ) , .A1( us23_n655 ) , .ZN( us23_n656 ) );
  NAND4_X1 us23_U67 (.A4( us23_n771 ) , .A3( us23_n772 ) , .A2( us23_n773 ) , .A1( us23_n774 ) , .ZN( us23_n800 ) );
  NOR3_X1 us23_U68 (.A3( us23_n764 ) , .A2( us23_n765 ) , .A1( us23_n766 ) , .ZN( us23_n772 ) );
  NOR4_X1 us23_U69 (.A4( us23_n767 ) , .A3( us23_n768 ) , .A2( us23_n769 ) , .A1( us23_n770 ) , .ZN( us23_n771 ) );
  NOR3_X1 us23_U7 (.A3( us23_n620 ) , .A2( us23_n621 ) , .ZN( us23_n635 ) , .A1( us23_n724 ) );
  AOI222_X1 us23_U70 (.ZN( us23_n774 ) , .A1( us23_n829 ) , .C1( us23_n833 ) , .B2( us23_n840 ) , .A2( us23_n849 ) , .B1( us23_n860 ) , .C2( us23_n872 ) );
  NOR4_X1 us23_U71 (.A4( us23_n576 ) , .A3( us23_n577 ) , .A2( us23_n578 ) , .ZN( us23_n585 ) , .A1( us23_n682 ) );
  NOR4_X1 us23_U72 (.A1( us23_n583 ) , .ZN( us23_n584 ) , .A3( us23_n651 ) , .A2( us23_n661 ) , .A4( us23_n766 ) );
  AOI221_X1 us23_U73 (.A( us23_n575 ) , .ZN( us23_n586 ) , .B2( us23_n830 ) , .C2( us23_n842 ) , .B1( us23_n853 ) , .C1( us23_n860 ) );
  NOR2_X1 us23_U74 (.ZN( us23_n760 ) , .A1( us23_n832 ) , .A2( us23_n833 ) );
  NAND4_X1 us23_U75 (.A4( us23_n455 ) , .A3( us23_n456 ) , .A2( us23_n457 ) , .A1( us23_n458 ) , .ZN( us23_n678 ) );
  NOR3_X1 us23_U76 (.ZN( us23_n456 ) , .A3( us23_n529 ) , .A1( us23_n554 ) , .A2( us23_n569 ) );
  NOR4_X1 us23_U77 (.ZN( us23_n457 ) , .A2( us23_n508 ) , .A1( us23_n598 ) , .A4( us23_n627 ) , .A3( us23_n710 ) );
  NOR4_X1 us23_U78 (.ZN( us23_n455 ) , .A2( us23_n516 ) , .A1( us23_n542 ) , .A3( us23_n578 ) , .A4( us23_n614 ) );
  NAND4_X1 us23_U79 (.A4( us23_n602 ) , .A3( us23_n603 ) , .A2( us23_n604 ) , .A1( us23_n605 ) , .ZN( us23_n721 ) );
  NOR2_X1 us23_U8 (.ZN( us23_n574 ) , .A1( us23_n621 ) , .A2( us23_n744 ) );
  NOR3_X1 us23_U80 (.A1( us23_n598 ) , .ZN( us23_n603 ) , .A3( us23_n662 ) , .A2( us23_n769 ) );
  NOR4_X1 us23_U81 (.A3( us23_n599 ) , .A2( us23_n600 ) , .A1( us23_n601 ) , .ZN( us23_n602 ) , .A4( us23_n654 ) );
  AOI222_X1 us23_U82 (.ZN( us23_n605 ) , .A1( us23_n829 ) , .C2( us23_n836 ) , .B1( us23_n841 ) , .A2( us23_n855 ) , .B2( us23_n860 ) , .C1( us23_n867 ) );
  NAND4_X1 us23_U83 (.A4( us23_n534 ) , .A3( us23_n535 ) , .A2( us23_n536 ) , .A1( us23_n537 ) , .ZN( us23_n621 ) );
  NOR4_X1 us23_U84 (.A4( us23_n525 ) , .A2( us23_n526 ) , .A1( us23_n527 ) , .ZN( us23_n537 ) , .A3( us23_n700 ) );
  NOR4_X1 us23_U85 (.A1( us23_n530 ) , .ZN( us23_n535 ) , .A2( us23_n653 ) , .A4( us23_n667 ) , .A3( us23_n764 ) );
  NOR4_X1 us23_U86 (.A4( us23_n528 ) , .A3( us23_n529 ) , .ZN( us23_n536 ) , .A2( us23_n683 ) , .A1( us23_n793 ) );
  NOR2_X1 us23_U87 (.ZN( us23_n685 ) , .A1( us23_n830 ) , .A2( us23_n831 ) );
  NAND4_X1 us23_U88 (.A4( us23_n547 ) , .A3( us23_n548 ) , .A2( us23_n549 ) , .A1( us23_n550 ) , .ZN( us23_n744 ) );
  NOR3_X1 us23_U89 (.ZN( us23_n548 ) , .A2( us23_n650 ) , .A1( us23_n666 ) , .A3( us23_n770 ) );
  NOR2_X1 us23_U9 (.A1( us23_n677 ) , .ZN( us23_n692 ) , .A2( us23_n806 ) );
  AOI211_X1 us23_U90 (.B( us23_n538 ) , .A( us23_n539 ) , .ZN( us23_n550 ) , .C2( us23_n838 ) , .C1( us23_n850 ) );
  NOR4_X1 us23_U91 (.A4( us23_n543 ) , .A3( us23_n544 ) , .A2( us23_n545 ) , .A1( us23_n546 ) , .ZN( us23_n547 ) );
  NAND4_X1 us23_U92 (.A4( us23_n478 ) , .A3( us23_n479 ) , .A2( us23_n480 ) , .A1( us23_n481 ) , .ZN( us23_n693 ) );
  NOR3_X1 us23_U93 (.ZN( us23_n479 ) , .A2( us23_n507 ) , .A3( us23_n600 ) , .A1( us23_n609 ) );
  AOI211_X1 us23_U94 (.B( us23_n476 ) , .A( us23_n477 ) , .ZN( us23_n481 ) , .C2( us23_n832 ) , .C1( us23_n860 ) );
  NOR4_X1 us23_U95 (.ZN( us23_n480 ) , .A3( us23_n531 ) , .A4( us23_n544 ) , .A2( us23_n566 ) , .A1( us23_n716 ) );
  NOR4_X1 us23_U96 (.ZN( us23_n619 ) , .A1( us23_n655 ) , .A3( us23_n665 ) , .A4( us23_n681 ) , .A2( us23_n765 ) );
  NOR4_X1 us23_U97 (.A4( us23_n608 ) , .A3( us23_n609 ) , .A2( us23_n610 ) , .A1( us23_n611 ) , .ZN( us23_n618 ) );
  NOR4_X1 us23_U98 (.A4( us23_n613 ) , .A3( us23_n614 ) , .A2( us23_n615 ) , .A1( us23_n616 ) , .ZN( us23_n617 ) );
  NAND4_X1 us23_U99 (.A4( us23_n484 ) , .A3( us23_n485 ) , .A2( us23_n486 ) , .A1( us23_n487 ) , .ZN( us23_n777 ) );
  NOR2_X1 us30_U10 (.ZN( us30_n575 ) , .A1( us30_n622 ) , .A2( us30_n745 ) );
  NOR2_X1 us30_U100 (.ZN( us30_n647 ) , .A1( us30_n854 ) , .A2( us30_n868 ) );
  NAND4_X1 us30_U101 (.A4( us30_n479 ) , .A3( us30_n480 ) , .A2( us30_n481 ) , .A1( us30_n482 ) , .ZN( us30_n694 ) );
  NOR3_X1 us30_U102 (.ZN( us30_n480 ) , .A2( us30_n508 ) , .A3( us30_n601 ) , .A1( us30_n610 ) );
  AOI211_X1 us30_U103 (.B( us30_n477 ) , .A( us30_n478 ) , .ZN( us30_n482 ) , .C2( us30_n833 ) , .C1( us30_n861 ) );
  NOR4_X1 us30_U104 (.ZN( us30_n481 ) , .A3( us30_n532 ) , .A4( us30_n545 ) , .A2( us30_n567 ) , .A1( us30_n717 ) );
  NAND4_X1 us30_U105 (.A4( us30_n548 ) , .A3( us30_n549 ) , .A2( us30_n550 ) , .A1( us30_n551 ) , .ZN( us30_n745 ) );
  NOR3_X1 us30_U106 (.ZN( us30_n549 ) , .A2( us30_n651 ) , .A1( us30_n667 ) , .A3( us30_n771 ) );
  AOI211_X1 us30_U107 (.B( us30_n539 ) , .A( us30_n540 ) , .ZN( us30_n551 ) , .C2( us30_n839 ) , .C1( us30_n851 ) );
  NOR4_X1 us30_U108 (.A4( us30_n544 ) , .A3( us30_n545 ) , .A2( us30_n546 ) , .A1( us30_n547 ) , .ZN( us30_n548 ) );
  NOR4_X1 us30_U109 (.ZN( us30_n620 ) , .A1( us30_n656 ) , .A3( us30_n666 ) , .A4( us30_n682 ) , .A2( us30_n766 ) );
  NOR2_X1 us30_U11 (.ZN( us30_n495 ) , .A1( us30_n678 ) , .A2( us30_n694 ) );
  NOR4_X1 us30_U110 (.A4( us30_n609 ) , .A3( us30_n610 ) , .A2( us30_n611 ) , .A1( us30_n612 ) , .ZN( us30_n619 ) );
  NOR4_X1 us30_U111 (.A4( us30_n614 ) , .A3( us30_n615 ) , .A2( us30_n616 ) , .A1( us30_n617 ) , .ZN( us30_n618 ) );
  NOR2_X1 us30_U112 (.ZN( us30_n686 ) , .A1( us30_n831 ) , .A2( us30_n832 ) );
  NAND4_X1 us30_U113 (.A4( us30_n485 ) , .A3( us30_n486 ) , .A2( us30_n487 ) , .A1( us30_n488 ) , .ZN( us30_n778 ) );
  NOR4_X1 us30_U114 (.A4( us30_n484 ) , .ZN( us30_n487 ) , .A1( us30_n566 ) , .A2( us30_n581 ) , .A3( us30_n602 ) );
  NOR4_X1 us30_U115 (.ZN( us30_n486 ) , .A1( us30_n507 ) , .A2( us30_n519 ) , .A4( us30_n546 ) , .A3( us30_n611 ) );
  NOR4_X1 us30_U116 (.ZN( us30_n485 ) , .A2( us30_n533 ) , .A1( us30_n558 ) , .A3( us30_n631 ) , .A4( us30_n718 ) );
  NAND4_X1 us30_U117 (.A4( us30_n691 ) , .A3( us30_n692 ) , .A1( us30_n693 ) , .ZN( us30_n776 ) , .A2( us30_n872 ) );
  AOI221_X1 us30_U118 (.A( us30_n681 ) , .ZN( us30_n692 ) , .B2( us30_n840 ) , .C1( us30_n842 ) , .C2( us30_n862 ) , .B1( us30_n865 ) );
  INV_X1 us30_U119 (.A( us30_n679 ) , .ZN( us30_n872 ) );
  NOR2_X1 us30_U12 (.A1( us30_n678 ) , .ZN( us30_n693 ) , .A2( us30_n807 ) );
  NOR4_X1 us30_U120 (.A4( us30_n687 ) , .A3( us30_n688 ) , .A2( us30_n689 ) , .A1( us30_n690 ) , .ZN( us30_n691 ) );
  NAND4_X1 us30_U121 (.A4( us30_n719 ) , .A3( us30_n720 ) , .A2( us30_n721 ) , .ZN( us30_n741 ) , .A1( us30_n857 ) );
  INV_X1 us30_U122 (.A( us30_n709 ) , .ZN( us30_n857 ) );
  AOI221_X1 us30_U123 (.A( us30_n710 ) , .ZN( us30_n721 ) , .C2( us30_n844 ) , .B2( us30_n845 ) , .C1( us30_n861 ) , .B1( us30_n862 ) );
  NOR4_X1 us30_U124 (.A4( us30_n715 ) , .A3( us30_n716 ) , .A2( us30_n717 ) , .A1( us30_n718 ) , .ZN( us30_n719 ) );
  NAND4_X1 us30_U125 (.A4( us30_n473 ) , .A3( us30_n474 ) , .A2( us30_n475 ) , .A1( us30_n476 ) , .ZN( us30_n678 ) );
  NOR4_X1 us30_U126 (.ZN( us30_n475 ) , .A1( us30_n531 ) , .A3( us30_n568 ) , .A4( us30_n600 ) , .A2( us30_n642 ) );
  NOR4_X1 us30_U127 (.A4( us30_n470 ) , .ZN( us30_n476 ) , .A3( us30_n556 ) , .A1( us30_n735 ) , .A2( us30_n755 ) );
  NOR4_X1 us30_U128 (.ZN( us30_n474 ) , .A1( us30_n506 ) , .A3( us30_n544 ) , .A2( us30_n583 ) , .A4( us30_n716 ) );
  NOR2_X1 us30_U129 (.ZN( us30_n733 ) , .A2( us30_n832 ) , .A1( us30_n845 ) );
  NOR3_X1 us30_U13 (.ZN( us30_n504 ) , .A2( us30_n679 ) , .A3( us30_n777 ) , .A1( us30_n876 ) );
  NOR2_X1 us30_U130 (.ZN( us30_n789 ) , .A2( us30_n862 ) , .A1( us30_n868 ) );
  NAND4_X1 us30_U131 (.A4( us30_n573 ) , .A3( us30_n574 ) , .A1( us30_n575 ) , .ZN( us30_n723 ) , .A2( us30_n874 ) );
  AOI221_X1 us30_U132 (.A( us30_n564 ) , .C2( us30_n565 ) , .ZN( us30_n574 ) , .B2( us30_n845 ) , .B1( us30_n852 ) , .C1( us30_n853 ) );
  NOR4_X1 us30_U133 (.A4( us30_n569 ) , .A3( us30_n570 ) , .A2( us30_n571 ) , .A1( us30_n572 ) , .ZN( us30_n573 ) );
  INV_X1 us30_U134 (.A( us30_n607 ) , .ZN( us30_n874 ) );
  NAND4_X1 us30_U135 (.A4( us30_n633 ) , .A3( us30_n634 ) , .A2( us30_n635 ) , .A1( us30_n636 ) , .ZN( us30_n743 ) );
  AOI211_X1 us30_U136 (.B( us30_n623 ) , .A( us30_n624 ) , .ZN( us30_n635 ) , .C2( us30_n836 ) , .C1( us30_n863 ) );
  NOR4_X1 us30_U137 (.A4( us30_n629 ) , .A3( us30_n630 ) , .A2( us30_n631 ) , .A1( us30_n632 ) , .ZN( us30_n633 ) );
  NOR4_X1 us30_U138 (.A4( us30_n626 ) , .A3( us30_n627 ) , .A2( us30_n628 ) , .ZN( us30_n634 ) , .A1( us30_n664 ) );
  NAND4_X1 us30_U139 (.A4( us30_n493 ) , .A3( us30_n494 ) , .A1( us30_n495 ) , .ZN( us30_n802 ) , .A2( us30_n867 ) );
  INV_X1 us30_U14 (.A( us30_n706 ) , .ZN( us30_n876 ) );
  AOI221_X1 us30_U140 (.A( us30_n489 ) , .ZN( us30_n494 ) , .B2( us30_n836 ) , .C2( us30_n841 ) , .C1( us30_n851 ) , .B1( us30_n860 ) );
  INV_X1 us30_U141 (.A( us30_n778 ) , .ZN( us30_n867 ) );
  NOR4_X1 us30_U142 (.A2( us30_n491 ) , .A1( us30_n492 ) , .ZN( us30_n493 ) , .A3( us30_n580 ) , .A4( us30_n612 ) );
  NOR4_X1 us30_U143 (.A4( us30_n734 ) , .A3( us30_n735 ) , .A2( us30_n736 ) , .A1( us30_n737 ) , .ZN( us30_n738 ) );
  AOI211_X1 us30_U144 (.B( us30_n725 ) , .A( us30_n726 ) , .ZN( us30_n739 ) , .C1( us30_n843 ) , .C2( us30_n855 ) );
  NOR3_X1 us30_U145 (.A3( us30_n722 ) , .A1( us30_n723 ) , .ZN( us30_n740 ) , .A2( us30_n741 ) );
  INV_X1 us30_U146 (.A( us30_n762 ) , .ZN( us30_n830 ) );
  OR4_X1 us30_U147 (.A4( us30_n566 ) , .A3( us30_n567 ) , .A2( us30_n568 ) , .ZN( us30_n572 ) , .A1( us30_n665 ) );
  OR4_X1 us30_U148 (.A4( us30_n682 ) , .A3( us30_n683 ) , .A2( us30_n684 ) , .A1( us30_n685 ) , .ZN( us30_n690 ) );
  OR4_X1 us30_U149 (.ZN( us30_n466 ) , .A4( us30_n518 ) , .A3( us30_n529 ) , .A2( us30_n578 ) , .A1( us30_n712 ) );
  INV_X1 us30_U15 (.A( us30_n680 ) , .ZN( us30_n840 ) );
  OR4_X1 us30_U150 (.A4( us30_n518 ) , .A2( us30_n519 ) , .A1( us30_n520 ) , .ZN( us30_n522 ) , .A3( us30_n821 ) );
  OR4_X1 us30_U151 (.ZN( us30_n492 ) , .A4( us30_n534 ) , .A2( us30_n547 ) , .A1( us30_n559 ) , .A3( us30_n632 ) );
  OR4_X1 us30_U152 (.A4( us30_n580 ) , .A3( us30_n581 ) , .A2( us30_n582 ) , .A1( us30_n583 ) , .ZN( us30_n584 ) );
  INV_X1 us30_U153 (.A( us30_n697 ) , .ZN( us30_n838 ) );
  NAND2_X1 us30_U154 (.ZN( us30_n613 ) , .A2( us30_n837 ) , .A1( us30_n873 ) );
  OR3_X1 us30_U155 (.A3( us30_n506 ) , .A2( us30_n507 ) , .A1( us30_n508 ) , .ZN( us30_n511 ) );
  INV_X1 us30_U156 (.A( us30_n754 ) , .ZN( us30_n869 ) );
  OAI21_X1 us30_U157 (.B1( us30_n753 ) , .ZN( us30_n754 ) , .A( us30_n845 ) , .B2( us30_n868 ) );
  INV_X1 us30_U158 (.A( us30_n463 ) , .ZN( us30_n864 ) );
  OAI21_X1 us30_U159 (.ZN( us30_n463 ) , .B1( us30_n809 ) , .A( us30_n834 ) , .B2( us30_n851 ) );
  NOR4_X1 us30_U16 (.A4( us30_n445 ) , .A3( us30_n446 ) , .A2( us30_n516 ) , .A1( us30_n541 ) , .ZN( us30_n706 ) );
  INV_X1 us30_U160 (.A( us30_n672 ) , .ZN( us30_n859 ) );
  AOI21_X1 us30_U161 (.A( us30_n670 ) , .B1( us30_n671 ) , .ZN( us30_n672 ) , .B2( us30_n856 ) );
  OAI222_X1 us30_U162 (.B2( us30_n747 ) , .B1( us30_n748 ) , .A2( us30_n749 ) , .ZN( us30_n757 ) , .C2( us30_n805 ) , .C1( us30_n814 ) , .A1( us30_n817 ) );
  OAI222_X1 us30_U163 (.ZN( us30_n505 ) , .C2( us30_n625 ) , .B2( us30_n647 ) , .B1( us30_n747 ) , .A2( us30_n748 ) , .C1( us30_n805 ) , .A1( us30_n806 ) );
  OAI222_X1 us30_U164 (.B2( us30_n708 ) , .ZN( us30_n709 ) , .C2( us30_n724 ) , .B1( us30_n747 ) , .A1( us30_n806 ) , .C1( us30_n814 ) , .A2( us30_n815 ) );
  NAND2_X1 us30_U165 (.A1( us30_n447 ) , .A2( us30_n465 ) , .ZN( us30_n749 ) );
  AOI22_X1 us30_U166 (.ZN( us30_n696 ) , .A1( us30_n830 ) , .B2( us30_n843 ) , .A2( us30_n865 ) , .B1( us30_n868 ) );
  AOI22_X1 us30_U167 (.A2( us30_n782 ) , .ZN( us30_n783 ) , .B2( us30_n831 ) , .A1( us30_n834 ) , .B1( us30_n863 ) );
  INV_X1 us30_U168 (.A( us30_n730 ) , .ZN( us30_n839 ) );
  AOI221_X1 us30_U169 (.A( us30_n764 ) , .ZN( us30_n774 ) , .C2( us30_n810 ) , .B2( us30_n835 ) , .C1( us30_n855 ) , .B1( us30_n866 ) );
  OR3_X1 us30_U17 (.ZN( us30_n446 ) , .A1( us30_n528 ) , .A3( us30_n577 ) , .A2( us30_n875 ) );
  AOI21_X1 us30_U170 (.B2( us30_n763 ) , .ZN( us30_n764 ) , .A( us30_n788 ) , .B1( us30_n792 ) );
  INV_X1 us30_U171 (.A( us30_n761 ) , .ZN( us30_n835 ) );
  AOI221_X1 us30_U172 (.A( us30_n483 ) , .ZN( us30_n488 ) , .B1( us30_n831 ) , .C2( us30_n844 ) , .C1( us30_n852 ) , .B2( us30_n862 ) );
  OAI22_X1 us30_U173 (.ZN( us30_n483 ) , .A1( us30_n708 ) , .B2( us30_n785 ) , .A2( us30_n806 ) , .B1( us30_n812 ) );
  INV_X1 us30_U174 (.A( us30_n790 ) , .ZN( us30_n832 ) );
  NAND2_X1 us30_U175 (.A1( us30_n451 ) , .A2( us30_n453 ) , .ZN( us30_n762 ) );
  OAI221_X1 us30_U176 (.A( us30_n727 ) , .C2( us30_n728 ) , .B2( us30_n729 ) , .B1( us30_n730 ) , .ZN( us30_n737 ) , .C1( us30_n817 ) );
  AOI22_X1 us30_U177 (.ZN( us30_n727 ) , .B1( us30_n832 ) , .A2( us30_n838 ) , .A1( us30_n863 ) , .B2( us30_n866 ) );
  INV_X1 us30_U178 (.A( us30_n786 ) , .ZN( us30_n862 ) );
  OAI22_X1 us30_U179 (.ZN( us30_n710 ) , .A2( us30_n728 ) , .B2( us30_n729 ) , .A1( us30_n744 ) , .B1( us30_n813 ) );
  OR4_X1 us30_U18 (.A4( us30_n442 ) , .A2( us30_n443 ) , .A1( us30_n444 ) , .ZN( us30_n445 ) , .A3( us30_n553 ) );
  INV_X1 us30_U180 (.A( us30_n816 ) , .ZN( us30_n831 ) );
  OAI22_X1 us30_U181 (.ZN( us30_n489 ) , .A1( us30_n724 ) , .B2( us30_n728 ) , .B1( us30_n730 ) , .A2( us30_n779 ) );
  OAI22_X1 us30_U182 (.ZN( us30_n624 ) , .B1( us30_n669 ) , .B2( us30_n747 ) , .A1( us30_n815 ) , .A2( us30_n816 ) );
  INV_X1 us30_U183 (.A( us30_n744 ) , .ZN( us30_n837 ) );
  INV_X1 us30_U184 (.A( us30_n788 ) , .ZN( us30_n845 ) );
  OAI22_X1 us30_U185 (.B2( us30_n779 ) , .B1( us30_n780 ) , .ZN( us30_n781 ) , .A2( us30_n814 ) , .A1( us30_n815 ) );
  OAI22_X1 us30_U186 (.A1( us30_n724 ) , .ZN( us30_n726 ) , .B2( us30_n750 ) , .B1( us30_n812 ) , .A2( us30_n816 ) );
  INV_X1 us30_U187 (.A( us30_n805 ) , .ZN( us30_n860 ) );
  INV_X1 us30_U188 (.A( us30_n814 ) , .ZN( us30_n833 ) );
  INV_X1 us30_U189 (.A( us30_n669 ) , .ZN( us30_n865 ) );
  INV_X1 us30_U19 (.A( us30_n613 ) , .ZN( us30_n875 ) );
  OAI22_X1 us30_U190 (.B2( us30_n744 ) , .ZN( us30_n746 ) , .A2( us30_n762 ) , .B1( us30_n780 ) , .A1( us30_n792 ) );
  OAI22_X1 us30_U191 (.ZN( us30_n496 ) , .A2( us30_n744 ) , .A1( us30_n780 ) , .B1( us30_n791 ) , .B2( us30_n806 ) );
  OAI22_X1 us30_U192 (.B2( us30_n803 ) , .B1( us30_n804 ) , .A2( us30_n805 ) , .A1( us30_n806 ) , .ZN( us30_n808 ) );
  AOI211_X1 us30_U193 (.A( us30_n637 ) , .ZN( us30_n645 ) , .B( us30_n743 ) , .C2( us30_n839 ) , .C1( us30_n854 ) );
  OAI22_X1 us30_U194 (.ZN( us30_n637 ) , .A1( us30_n699 ) , .B2( us30_n728 ) , .A2( us30_n762 ) , .B1( us30_n816 ) );
  OAI22_X1 us30_U195 (.B1( us30_n490 ) , .ZN( us30_n491 ) , .A1( us30_n686 ) , .A2( us30_n763 ) , .B2( us30_n817 ) );
  NOR3_X1 us30_U196 (.ZN( us30_n490 ) , .A1( us30_n782 ) , .A2( us30_n850 ) , .A3( us30_n863 ) );
  INV_X1 us30_U197 (.A( us30_n750 ) , .ZN( us30_n842 ) );
  OAI22_X1 us30_U198 (.ZN( us30_n695 ) , .A2( us30_n730 ) , .A1( us30_n780 ) , .B1( us30_n791 ) , .B2( us30_n817 ) );
  NOR2_X1 us30_U199 (.ZN( us30_n715 ) , .A1( us30_n805 ) , .A2( us30_n817 ) );
  INV_X1 us30_U20 (.A( us30_n749 ) , .ZN( us30_n863 ) );
  NOR2_X1 us30_U200 (.ZN( us30_n666 ) , .A1( us30_n728 ) , .A2( us30_n803 ) );
  NOR2_X1 us30_U201 (.ZN( us30_n594 ) , .A2( us30_n697 ) , .A1( us30_n728 ) );
  NOR2_X1 us30_U202 (.ZN( us30_n570 ) , .A1( us30_n728 ) , .A2( us30_n806 ) );
  NOR2_X1 us30_U203 (.A2( us30_n744 ) , .ZN( us30_n755 ) , .A1( us30_n805 ) );
  NOR2_X1 us30_U204 (.ZN( us30_n735 ) , .A2( us30_n803 ) , .A1( us30_n805 ) );
  NOR2_X1 us30_U205 (.ZN( us30_n546 ) , .A2( us30_n780 ) , .A1( us30_n814 ) );
  NOR2_X1 us30_U206 (.ZN( us30_n577 ) , .A2( us30_n699 ) , .A1( us30_n814 ) );
  NOR2_X1 us30_U207 (.ZN( us30_n654 ) , .A1( us30_n728 ) , .A2( us30_n813 ) );
  NOR2_X1 us30_U208 (.ZN( us30_n718 ) , .A2( us30_n724 ) , .A1( us30_n744 ) );
  NOR2_X1 us30_U209 (.ZN( us30_n532 ) , .A2( us30_n749 ) , .A1( us30_n750 ) );
  AOI222_X1 us30_U21 (.ZN( us30_n605 ) , .B2( us30_n671 ) , .B1( us30_n753 ) , .C2( us30_n831 ) , .A1( us30_n833 ) , .A2( us30_n862 ) , .C1( us30_n863 ) );
  NOR2_X1 us30_U210 (.ZN( us30_n615 ) , .A1( us30_n785 ) , .A2( us30_n815 ) );
  NOR2_X1 us30_U211 (.ZN( us30_n629 ) , .A2( us30_n728 ) , .A1( us30_n785 ) );
  NOR2_X1 us30_U212 (.ZN( us30_n611 ) , .A2( us30_n780 ) , .A1( us30_n806 ) );
  NOR2_X1 us30_U213 (.ZN( us30_n628 ) , .A2( us30_n669 ) , .A1( us30_n785 ) );
  INV_X1 us30_U214 (.A( us30_n747 ) , .ZN( us30_n834 ) );
  INV_X1 us30_U215 (.A( us30_n728 ) , .ZN( us30_n852 ) );
  NOR2_X1 us30_U216 (.ZN( us30_n652 ) , .A1( us30_n669 ) , .A2( us30_n814 ) );
  NOR2_X1 us30_U217 (.A1( us30_n669 ) , .ZN( us30_n673 ) , .A2( us30_n744 ) );
  NOR2_X1 us30_U218 (.ZN( us30_n602 ) , .A1( us30_n669 ) , .A2( us30_n803 ) );
  NOR2_X1 us30_U219 (.A1( us30_n669 ) , .ZN( us30_n688 ) , .A2( us30_n816 ) );
  AOI222_X1 us30_U22 (.ZN( us30_n563 ) , .B1( us30_n830 ) , .C1( us30_n841 ) , .A2( us30_n843 ) , .A1( us30_n854 ) , .B2( us30_n863 ) , .C2( us30_n873 ) );
  NOR2_X1 us30_U220 (.A2( us30_n744 ) , .ZN( us30_n769 ) , .A1( us30_n812 ) );
  NOR2_X1 us30_U221 (.ZN( us30_n531 ) , .A2( us30_n780 ) , .A1( us30_n816 ) );
  INV_X1 us30_U222 (.A( us30_n792 ) , .ZN( us30_n851 ) );
  NOR2_X1 us30_U223 (.A2( us30_n708 ) , .A1( us30_n750 ) , .ZN( us30_n771 ) );
  NOR2_X1 us30_U224 (.ZN( us30_n599 ) , .A2( us30_n791 ) , .A1( us30_n816 ) );
  NOR2_X1 us30_U225 (.A1( us30_n669 ) , .ZN( us30_n766 ) , .A2( us30_n813 ) );
  NOR2_X1 us30_U226 (.ZN( us30_n601 ) , .A2( us30_n780 ) , .A1( us30_n803 ) );
  NOR2_X1 us30_U227 (.A1( us30_n699 ) , .ZN( us30_n768 ) , .A2( us30_n813 ) );
  NOR2_X1 us30_U228 (.ZN( us30_n541 ) , .A2( us30_n697 ) , .A1( us30_n699 ) );
  NOR2_X1 us30_U229 (.ZN( us30_n527 ) , .A1( us30_n669 ) , .A2( us30_n779 ) );
  AOI222_X1 us30_U23 (.ZN( us30_n660 ) , .A2( us30_n839 ) , .B1( us30_n841 ) , .C2( us30_n845 ) , .A1( us30_n860 ) , .C1( us30_n863 ) , .B2( us30_n870 ) );
  NOR2_X1 us30_U230 (.ZN( us30_n667 ) , .A1( us30_n750 ) , .A2( us30_n815 ) );
  NOR2_X1 us30_U231 (.ZN( us30_n555 ) , .A1( us30_n750 ) , .A2( us30_n791 ) );
  NOR2_X1 us30_U232 (.ZN( us30_n508 ) , .A2( us30_n780 ) , .A1( us30_n785 ) );
  NOR2_X1 us30_U233 (.ZN( us30_n543 ) , .A2( us30_n708 ) , .A1( us30_n785 ) );
  NOR2_X1 us30_U234 (.ZN( us30_n528 ) , .A2( us30_n724 ) , .A1( us30_n803 ) );
  NOR2_X1 us30_U235 (.ZN( us30_n664 ) , .A1( us30_n785 ) , .A2( us30_n791 ) );
  NOR2_X1 us30_U236 (.ZN( us30_n556 ) , .A1( us30_n762 ) , .A2( us30_n805 ) );
  INV_X1 us30_U237 (.A( us30_n806 ) , .ZN( us30_n841 ) );
  NOR2_X1 us30_U238 (.ZN( us30_n661 ) , .A1( us30_n729 ) , .A2( us30_n790 ) );
  OAI22_X1 us30_U239 (.B1( us30_n440 ) , .ZN( us30_n444 ) , .A2( us30_n728 ) , .A1( us30_n744 ) , .B2( us30_n749 ) );
  INV_X1 us30_U24 (.A( us30_n647 ) , .ZN( us30_n870 ) );
  NOR3_X1 us30_U240 (.ZN( us30_n440 ) , .A2( us30_n836 ) , .A3( us30_n837 ) , .A1( us30_n846 ) );
  NOR2_X1 us30_U241 (.ZN( us30_n507 ) , .A1( us30_n812 ) , .A2( us30_n817 ) );
  NOR2_X1 us30_U242 (.ZN( us30_n557 ) , .A1( us30_n792 ) , .A2( us30_n814 ) );
  NOR2_X1 us30_U243 (.ZN( us30_n545 ) , .A1( us30_n749 ) , .A2( us30_n814 ) );
  NOR2_X1 us30_U244 (.ZN( us30_n509 ) , .A1( us30_n729 ) , .A2( us30_n779 ) );
  NOR2_X1 us30_U245 (.ZN( us30_n662 ) , .A2( us30_n697 ) , .A1( us30_n729 ) );
  OAI22_X1 us30_U246 (.B2( us30_n750 ) , .B1( us30_n751 ) , .A1( us30_n752 ) , .ZN( us30_n756 ) , .A2( us30_n806 ) );
  NOR2_X1 us30_U247 (.ZN( us30_n751 ) , .A2( us30_n852 ) , .A1( us30_n860 ) );
  NOR3_X1 us30_U248 (.ZN( us30_n752 ) , .A2( us30_n853 ) , .A1( us30_n863 ) , .A3( us30_n865 ) );
  NOR2_X1 us30_U249 (.ZN( us30_n544 ) , .A2( us30_n785 ) , .A1( us30_n792 ) );
  NOR4_X1 us30_U25 (.ZN( us30_n473 ) , .A2( us30_n521 ) , .A4( us30_n594 ) , .A1( us30_n609 ) , .A3( us30_n629 ) );
  NOR2_X1 us30_U250 (.ZN( us30_n663 ) , .A1( us30_n729 ) , .A2( us30_n785 ) );
  NOR2_X1 us30_U251 (.ZN( us30_n530 ) , .A2( us30_n744 ) , .A1( us30_n792 ) );
  NOR2_X1 us30_U252 (.ZN( us30_n506 ) , .A2( us30_n728 ) , .A1( us30_n762 ) );
  NOR2_X1 us30_U253 (.ZN( us30_n631 ) , .A1( us30_n724 ) , .A2( us30_n813 ) );
  NOR2_X1 us30_U254 (.ZN( us30_n614 ) , .A1( us30_n762 ) , .A2( us30_n812 ) );
  NOR2_X1 us30_U255 (.A1( us30_n749 ) , .ZN( us30_n767 ) , .A2( us30_n803 ) );
  NOR2_X1 us30_U256 (.ZN( us30_n516 ) , .A1( us30_n708 ) , .A2( us30_n744 ) );
  NOR2_X1 us30_U257 (.ZN( us30_n670 ) , .A1( us30_n790 ) , .A2( us30_n805 ) );
  NOR2_X1 us30_U258 (.ZN( us30_n558 ) , .A1( us30_n708 ) , .A2( us30_n816 ) );
  NOR2_X1 us30_U259 (.A2( us30_n697 ) , .ZN( us30_n716 ) , .A1( us30_n792 ) );
  NOR4_X1 us30_U26 (.ZN( us30_n479 ) , .A1( us30_n520 ) , .A4( us30_n557 ) , .A3( us30_n582 ) , .A2( us30_n630 ) );
  NOR2_X1 us30_U260 (.ZN( us30_n517 ) , .A1( us30_n708 ) , .A2( us30_n803 ) );
  NOR2_X1 us30_U261 (.ZN( us30_n521 ) , .A1( us30_n790 ) , .A2( us30_n812 ) );
  NOR2_X1 us30_U262 (.ZN( us30_n630 ) , .A1( us30_n747 ) , .A2( us30_n815 ) );
  NOR2_X1 us30_U263 (.ZN( us30_n655 ) , .A1( us30_n790 ) , .A2( us30_n815 ) );
  INV_X1 us30_U264 (.A( us30_n763 ) , .ZN( us30_n866 ) );
  AOI21_X1 us30_U265 (.ZN( us30_n552 ) , .B1( us30_n669 ) , .A( us30_n697 ) , .B2( us30_n805 ) );
  NOR2_X1 us30_U266 (.ZN( us30_n668 ) , .A2( us30_n708 ) , .A1( us30_n790 ) );
  NOR2_X1 us30_U267 (.ZN( us30_n542 ) , .A1( us30_n762 ) , .A2( us30_n791 ) );
  NOR2_X1 us30_U268 (.ZN( us30_n656 ) , .A1( us30_n747 ) , .A2( us30_n780 ) );
  NOR2_X1 us30_U269 (.ZN( us30_n609 ) , .A2( us30_n724 ) , .A1( us30_n817 ) );
  NOR4_X1 us30_U27 (.A4( us30_n532 ) , .A3( us30_n533 ) , .A2( us30_n534 ) , .ZN( us30_n535 ) , .A1( us30_n820 ) );
  INV_X1 us30_U270 (.A( us30_n729 ) , .ZN( us30_n868 ) );
  AOI21_X1 us30_U271 (.B1( us30_n625 ) , .ZN( us30_n627 ) , .A( us30_n763 ) , .B2( us30_n814 ) );
  AOI21_X1 us30_U272 (.ZN( us30_n650 ) , .A( us30_n779 ) , .B1( us30_n792 ) , .B2( us30_n805 ) );
  AOI21_X1 us30_U273 (.A( us30_n815 ) , .B2( us30_n816 ) , .B1( us30_n817 ) , .ZN( us30_n818 ) );
  NOR2_X1 us30_U274 (.ZN( us30_n579 ) , .A2( us30_n708 ) , .A1( us30_n730 ) );
  NOR2_X1 us30_U275 (.ZN( us30_n533 ) , .A2( us30_n724 ) , .A1( us30_n730 ) );
  NOR2_X1 us30_U276 (.ZN( us30_n642 ) , .A2( us30_n788 ) , .A1( us30_n791 ) );
  AOI21_X1 us30_U277 (.A( us30_n812 ) , .B2( us30_n813 ) , .B1( us30_n814 ) , .ZN( us30_n819 ) );
  NOR2_X1 us30_U278 (.A2( us30_n708 ) , .A1( us30_n762 ) , .ZN( us30_n794 ) );
  NOR2_X1 us30_U279 (.A2( us30_n697 ) , .A1( us30_n780 ) , .ZN( us30_n820 ) );
  NOR4_X1 us30_U28 (.ZN( us30_n456 ) , .A2( us30_n517 ) , .A1( us30_n543 ) , .A3( us30_n579 ) , .A4( us30_n615 ) );
  AOI21_X1 us30_U280 (.ZN( us30_n626 ) , .B2( us30_n669 ) , .A( us30_n790 ) , .B1( us30_n791 ) );
  AOI21_X1 us30_U281 (.ZN( us30_n499 ) , .B1( us30_n680 ) , .A( us30_n812 ) , .B2( us30_n816 ) );
  NOR2_X1 us30_U282 (.ZN( us30_n520 ) , .A2( us30_n708 ) , .A1( us30_n814 ) );
  AOI21_X1 us30_U283 (.ZN( us30_n477 ) , .A( us30_n669 ) , .B1( us30_n750 ) , .B2( us30_n806 ) );
  NOR2_X1 us30_U284 (.ZN( us30_n582 ) , .A1( us30_n744 ) , .A2( us30_n815 ) );
  AOI21_X1 us30_U285 (.ZN( us30_n593 ) , .B1( us30_n750 ) , .A( us30_n792 ) , .B2( us30_n813 ) );
  AOI21_X1 us30_U286 (.ZN( us30_n515 ) , .A( us30_n729 ) , .B1( us30_n750 ) , .B2( us30_n803 ) );
  NOR2_X1 us30_U287 (.A1( us30_n697 ) , .ZN( us30_n770 ) , .A2( us30_n815 ) );
  AOI21_X1 us30_U288 (.ZN( us30_n510 ) , .B2( us30_n669 ) , .A( us30_n730 ) , .B1( us30_n815 ) );
  NOR2_X1 us30_U289 (.ZN( us30_n519 ) , .A2( us30_n699 ) , .A1( us30_n816 ) );
  NOR4_X1 us30_U29 (.A4( us30_n541 ) , .A3( us30_n542 ) , .A2( us30_n543 ) , .ZN( us30_n550 ) , .A1( us30_n688 ) );
  NOR2_X1 us30_U290 (.ZN( us30_n559 ) , .A2( us30_n791 ) , .A1( us30_n803 ) );
  NOR2_X1 us30_U291 (.ZN( us30_n581 ) , .A1( us30_n669 ) , .A2( us30_n788 ) );
  INV_X1 us30_U292 (.A( us30_n813 ) , .ZN( us30_n836 ) );
  NOR2_X1 us30_U293 (.ZN( us30_n683 ) , .A2( us30_n699 ) , .A1( us30_n803 ) );
  AOI21_X1 us30_U294 (.ZN( us30_n589 ) , .B2( us30_n699 ) , .B1( us30_n815 ) , .A( us30_n817 ) );
  AOI21_X1 us30_U295 (.ZN( us30_n539 ) , .B2( us30_n812 ) , .A( us30_n814 ) , .B1( us30_n815 ) );
  AOI21_X1 us30_U296 (.ZN( us30_n540 ) , .A( us30_n763 ) , .B2( us30_n779 ) , .B1( us30_n817 ) );
  AOI21_X1 us30_U297 (.B1( us30_n699 ) , .ZN( us30_n700 ) , .A( us30_n732 ) , .B2( us30_n763 ) );
  AOI21_X1 us30_U298 (.ZN( us30_n591 ) , .B2( us30_n763 ) , .A( us30_n785 ) , .B1( us30_n812 ) );
  AOI21_X1 us30_U299 (.ZN( us30_n498 ) , .A( us30_n724 ) , .B2( us30_n762 ) , .B1( us30_n814 ) );
  NAND2_X1 us30_U3 (.A2( us30_n448 ) , .A1( us30_n464 ) , .ZN( us30_n815 ) );
  AOI221_X1 us30_U30 (.A( us30_n713 ) , .B2( us30_n714 ) , .ZN( us30_n720 ) , .C1( us30_n832 ) , .B1( us30_n839 ) , .C2( us30_n863 ) );
  NOR2_X1 us30_U300 (.ZN( us30_n547 ) , .A1( us30_n699 ) , .A2( us30_n744 ) );
  INV_X1 us30_U301 (.A( us30_n791 ) , .ZN( us30_n873 ) );
  AOI21_X1 us30_U302 (.ZN( us30_n649 ) , .B1( us30_n729 ) , .B2( us30_n763 ) , .A( us30_n813 ) );
  NOR2_X1 us30_U303 (.ZN( us30_n685 ) , .A1( us30_n729 ) , .A2( us30_n816 ) );
  AOI21_X1 us30_U304 (.B1( us30_n686 ) , .ZN( us30_n687 ) , .A( us30_n728 ) , .B2( us30_n761 ) );
  AOI21_X1 us30_U305 (.ZN( us30_n569 ) , .B1( us30_n750 ) , .B2( us30_n762 ) , .A( us30_n780 ) );
  AOI21_X1 us30_U306 (.ZN( us30_n571 ) , .B2( us30_n697 ) , .B1( us30_n806 ) , .A( us30_n812 ) );
  NOR2_X1 us30_U307 (.ZN( us30_n568 ) , .A1( us30_n729 ) , .A2( us30_n762 ) );
  NOR2_X1 us30_U308 (.ZN( us30_n566 ) , .A2( us30_n697 ) , .A1( us30_n763 ) );
  AOI21_X1 us30_U309 (.ZN( us30_n640 ) , .B2( us30_n747 ) , .A( us30_n792 ) , .B1( us30_n803 ) );
  OR2_X1 us30_U31 (.A2( us30_n711 ) , .A1( us30_n712 ) , .ZN( us30_n713 ) );
  INV_X1 us30_U310 (.A( us30_n699 ) , .ZN( us30_n853 ) );
  AOI21_X1 us30_U311 (.ZN( us30_n514 ) , .A( us30_n779 ) , .B2( us30_n792 ) , .B1( us30_n812 ) );
  AOI21_X1 us30_U312 (.ZN( us30_n639 ) , .B2( us30_n749 ) , .A( us30_n788 ) , .B1( us30_n812 ) );
  NAND2_X1 us30_U313 (.ZN( us30_n753 ) , .A1( us30_n763 ) , .A2( us30_n805 ) );
  NOR2_X1 us30_U314 (.ZN( us30_n665 ) , .A1( us30_n780 ) , .A2( us30_n813 ) );
  AOI21_X1 us30_U315 (.ZN( us30_n564 ) , .B1( us30_n724 ) , .A( us30_n779 ) , .B2( us30_n791 ) );
  AOI21_X1 us30_U316 (.ZN( us30_n497 ) , .A( us30_n779 ) , .B2( us30_n791 ) , .B1( us30_n804 ) );
  AOI21_X1 us30_U317 (.ZN( us30_n689 ) , .B2( us30_n749 ) , .B1( us30_n763 ) , .A( us30_n806 ) );
  AOI21_X1 us30_U318 (.ZN( us30_n450 ) , .B2( us30_n792 ) , .A( us30_n803 ) , .B1( us30_n815 ) );
  NOR2_X1 us30_U319 (.ZN( us30_n567 ) , .A1( us30_n747 ) , .A2( us30_n805 ) );
  NOR2_X1 us30_U32 (.ZN( us30_n680 ) , .A2( us30_n834 ) , .A1( us30_n839 ) );
  NOR2_X1 us30_U320 (.ZN( us30_n529 ) , .A1( us30_n708 ) , .A2( us30_n779 ) );
  NOR2_X1 us30_U321 (.ZN( us30_n578 ) , .A1( us30_n708 ) , .A2( us30_n813 ) );
  AOI21_X1 us30_U322 (.ZN( us30_n478 ) , .B2( us30_n697 ) , .A( us30_n749 ) , .B1( us30_n779 ) );
  AOI21_X1 us30_U323 (.A( us30_n790 ) , .B2( us30_n791 ) , .B1( us30_n792 ) , .ZN( us30_n793 ) );
  NOR2_X1 us30_U324 (.ZN( us30_n684 ) , .A1( us30_n791 ) , .A2( us30_n813 ) );
  AOI21_X1 us30_U325 (.A( us30_n733 ) , .ZN( us30_n734 ) , .B2( us30_n780 ) , .B1( us30_n792 ) );
  NOR2_X1 us30_U326 (.A2( us30_n813 ) , .A1( us30_n815 ) , .ZN( us30_n821 ) );
  AOI21_X1 us30_U327 (.ZN( us30_n641 ) , .B1( us30_n680 ) , .A( us30_n791 ) , .B2( us30_n817 ) );
  NOR2_X1 us30_U328 (.ZN( us30_n711 ) , .A1( us30_n762 ) , .A2( us30_n763 ) );
  NOR2_X1 us30_U329 (.ZN( us30_n583 ) , .A1( us30_n792 ) , .A2( us30_n817 ) );
  AOI222_X1 us30_U33 (.ZN( us30_n469 ) , .B1( us30_n832 ) , .A1( us30_n839 ) , .C1( us30_n842 ) , .C2( us30_n851 ) , .A2( us30_n855 ) , .B2( us30_n865 ) );
  NOR2_X1 us30_U330 (.ZN( us30_n534 ) , .A1( us30_n724 ) , .A2( us30_n788 ) );
  NOR2_X1 us30_U331 (.ZN( us30_n632 ) , .A2( us30_n697 ) , .A1( us30_n724 ) );
  NOR2_X1 us30_U332 (.ZN( us30_n682 ) , .A2( us30_n708 ) , .A1( us30_n817 ) );
  NOR2_X1 us30_U333 (.ZN( us30_n580 ) , .A2( us30_n697 ) , .A1( us30_n791 ) );
  INV_X1 us30_U334 (.A( us30_n815 ) , .ZN( us30_n855 ) );
  AOI21_X1 us30_U335 (.ZN( us30_n442 ) , .A( us30_n699 ) , .B1( us30_n733 ) , .B2( us30_n750 ) );
  INV_X1 us30_U336 (.A( us30_n780 ) , .ZN( us30_n850 ) );
  INV_X1 us30_U337 (.A( us30_n785 ) , .ZN( us30_n846 ) );
  NAND2_X1 us30_U338 (.ZN( us30_n714 ) , .A1( us30_n728 ) , .A2( us30_n780 ) );
  NAND2_X1 us30_U339 (.A2( us30_n762 ) , .A1( us30_n806 ) , .ZN( us30_n810 ) );
  NOR4_X1 us30_U34 (.A1( us30_n466 ) , .ZN( us30_n467 ) , .A4( us30_n542 ) , .A2( us30_n554 ) , .A3( us30_n614 ) );
  AOI21_X1 us30_U340 (.ZN( us30_n443 ) , .B1( us30_n789 ) , .B2( us30_n791 ) , .A( us30_n814 ) );
  NAND2_X1 us30_U341 (.ZN( us30_n671 ) , .A1( us30_n806 ) , .A2( us30_n816 ) );
  NOR2_X1 us30_U342 (.ZN( us30_n484 ) , .A1( us30_n788 ) , .A2( us30_n805 ) );
  NOR2_X1 us30_U343 (.ZN( us30_n470 ) , .A2( us30_n779 ) , .A1( us30_n815 ) );
  NOR2_X1 us30_U344 (.ZN( us30_n712 ) , .A2( us30_n724 ) , .A1( us30_n790 ) );
  OAI21_X1 us30_U345 (.A( us30_n787 ) , .B2( us30_n788 ) , .B1( us30_n789 ) , .ZN( us30_n795 ) );
  OAI21_X1 us30_U346 (.ZN( us30_n787 ) , .A( us30_n839 ) , .B1( us30_n863 ) , .B2( us30_n873 ) );
  NOR2_X1 us30_U347 (.ZN( us30_n526 ) , .A1( us30_n724 ) , .A2( us30_n750 ) );
  NAND2_X1 us30_U348 (.A1( us30_n699 ) , .A2( us30_n729 ) , .ZN( us30_n782 ) );
  NOR2_X1 us30_U349 (.ZN( us30_n518 ) , .A1( us30_n708 ) , .A2( us30_n788 ) );
  AOI221_X1 us30_U35 (.ZN( us30_n468 ) , .C2( us30_n714 ) , .B2( us30_n831 ) , .C1( us30_n845 ) , .B1( us30_n860 ) , .A( us30_n864 ) );
  OAI21_X1 us30_U350 (.A( us30_n698 ) , .ZN( us30_n702 ) , .B2( us30_n750 ) , .B1( us30_n804 ) );
  OAI21_X1 us30_U351 (.ZN( us30_n698 ) , .B2( us30_n833 ) , .B1( us30_n838 ) , .A( us30_n860 ) );
  OAI21_X1 us30_U352 (.A( us30_n731 ) , .B1( us30_n732 ) , .ZN( us30_n736 ) , .B2( us30_n805 ) );
  OAI21_X1 us30_U353 (.ZN( us30_n731 ) , .A( us30_n833 ) , .B2( us30_n852 ) , .B1( us30_n873 ) );
  INV_X1 us30_U354 (.A( us30_n817 ) , .ZN( us30_n844 ) );
  INV_X1 us30_U355 (.A( us30_n724 ) , .ZN( us30_n856 ) );
  AND2_X1 us30_U356 (.ZN( us30_n732 ) , .A1( us30_n779 ) , .A2( us30_n785 ) );
  NAND2_X1 us30_U357 (.A1( us30_n447 ) , .A2( us30_n449 ) , .ZN( us30_n805 ) );
  NAND2_X1 us30_U358 (.A1( us30_n451 ) , .A2( us30_n454 ) , .ZN( us30_n814 ) );
  NAND2_X1 us30_U359 (.A1( us30_n452 ) , .A2( us30_n465 ) , .ZN( us30_n669 ) );
  NOR4_X1 us30_U36 (.A4( us30_n514 ) , .A3( us30_n515 ) , .A2( us30_n516 ) , .A1( us30_n517 ) , .ZN( us30_n524 ) );
  NAND2_X1 us30_U360 (.A2( us30_n448 ) , .A1( us30_n460 ) , .ZN( us30_n728 ) );
  NAND2_X1 us30_U361 (.A1( us30_n455 ) , .A2( us30_n462 ) , .ZN( us30_n750 ) );
  NAND2_X1 us30_U362 (.A2( us30_n453 ) , .A1( us30_n455 ) , .ZN( us30_n806 ) );
  NAND2_X1 us30_U363 (.A1( us30_n451 ) , .A2( us30_n471 ) , .ZN( us30_n816 ) );
  NAND2_X1 us30_U364 (.A1( us30_n454 ) , .A2( us30_n461 ) , .ZN( us30_n813 ) );
  NAND2_X1 us30_U365 (.A1( us30_n455 ) , .A2( us30_n471 ) , .ZN( us30_n803 ) );
  NAND2_X1 us30_U366 (.A1( us30_n453 ) , .A2( us30_n461 ) , .ZN( us30_n744 ) );
  NAND2_X1 us30_U367 (.A1( us30_n453 ) , .A2( us30_n472 ) , .ZN( us30_n785 ) );
  NAND2_X1 us30_U368 (.A2( us30_n454 ) , .A1( us30_n472 ) , .ZN( us30_n779 ) );
  NAND2_X1 us30_U369 (.A2( us30_n464 ) , .A1( us30_n465 ) , .ZN( us30_n812 ) );
  AOI222_X1 us30_U37 (.ZN( us30_n525 ) , .A1( us30_n834 ) , .B2( us30_n837 ) , .C1( us30_n844 ) , .C2( us30_n850 ) , .A2( us30_n852 ) , .B1( us30_n866 ) );
  NAND2_X1 us30_U370 (.A1( us30_n441 ) , .A2( us30_n460 ) , .ZN( us30_n699 ) );
  NAND2_X1 us30_U371 (.A2( us30_n449 ) , .A1( us30_n452 ) , .ZN( us30_n763 ) );
  NAND2_X1 us30_U372 (.A2( us30_n448 ) , .A1( us30_n452 ) , .ZN( us30_n729 ) );
  NAND2_X1 us30_U373 (.A2( us30_n461 ) , .A1( us30_n462 ) , .ZN( us30_n747 ) );
  NAND2_X1 us30_U374 (.A1( us30_n462 ) , .A2( us30_n472 ) , .ZN( us30_n788 ) );
  NOR2_X1 us30_U375 (.ZN( us30_n465 ) , .A2( us30_n847 ) , .A1( us30_n848 ) );
  NOR2_X1 us30_U376 (.ZN( us30_n453 ) , .A1( us30_n826 ) , .A2( us30_n827 ) );
  NOR2_X1 us30_U377 (.ZN( us30_n451 ) , .A1( us30_n828 ) , .A2( us30_n829 ) );
  NAND2_X1 us30_U378 (.A1( us30_n451 ) , .A2( us30_n462 ) , .ZN( us30_n790 ) );
  NAND2_X1 us30_U379 (.A2( us30_n441 ) , .A1( us30_n447 ) , .ZN( us30_n784 ) );
  NOR4_X1 us30_U38 (.A3( us30_n521 ) , .A1( us30_n522 ) , .ZN( us30_n523 ) , .A2( us30_n673 ) , .A4( us30_n769 ) );
  NAND2_X1 us30_U380 (.A2( us30_n454 ) , .A1( us30_n455 ) , .ZN( us30_n730 ) );
  NAND2_X2 us30_U381 (.A1( us30_n449 ) , .A2( us30_n464 ) , .ZN( us30_n724 ) );
  NAND2_X2 us30_U382 (.A1( us30_n449 ) , .A2( us30_n460 ) , .ZN( us30_n792 ) );
  NAND2_X2 us30_U383 (.A2( us30_n460 ) , .A1( us30_n465 ) , .ZN( us30_n780 ) );
  NOR2_X1 us30_U384 (.ZN( us30_n447 ) , .A2( us30_n849 ) , .A1( us30_n858 ) );
  NAND2_X1 us30_U385 (.A1( us30_n447 ) , .A2( us30_n448 ) , .ZN( us30_n786 ) );
  NOR2_X1 us30_U386 (.A2( sa30_6 ) , .A1( sa30_7 ) , .ZN( us30_n464 ) );
  NOR2_X1 us30_U387 (.A2( sa30_7 ) , .ZN( us30_n460 ) , .A1( us30_n849 ) );
  NOR2_X1 us30_U388 (.A2( sa30_4 ) , .ZN( us30_n449 ) , .A1( us30_n848 ) );
  NOR2_X1 us30_U389 (.A2( sa30_4 ) , .A1( sa30_5 ) , .ZN( us30_n441 ) );
  AOI221_X1 us30_U39 (.A( us30_n781 ) , .ZN( us30_n798 ) , .C2( us30_n837 ) , .B2( us30_n838 ) , .B1( us30_n865 ) , .C1( us30_n866 ) );
  NOR2_X1 us30_U390 (.A2( sa30_5 ) , .ZN( us30_n448 ) , .A1( us30_n847 ) );
  NOR2_X1 us30_U391 (.A2( sa30_2 ) , .A1( sa30_3 ) , .ZN( us30_n472 ) );
  NOR2_X1 us30_U392 (.A2( sa30_6 ) , .ZN( us30_n452 ) , .A1( us30_n858 ) );
  NOR2_X1 us30_U393 (.A2( sa30_1 ) , .ZN( us30_n471 ) , .A1( us30_n826 ) );
  NOR2_X1 us30_U394 (.A2( sa30_0 ) , .ZN( us30_n454 ) , .A1( us30_n827 ) );
  NOR2_X1 us30_U395 (.A2( sa30_0 ) , .A1( sa30_1 ) , .ZN( us30_n462 ) );
  NOR2_X1 us30_U396 (.A2( sa30_3 ) , .ZN( us30_n455 ) , .A1( us30_n828 ) );
  NOR2_X1 us30_U397 (.A2( sa30_2 ) , .ZN( us30_n461 ) , .A1( us30_n829 ) );
  INV_X1 us30_U398 (.A( sa30_6 ) , .ZN( us30_n849 ) );
  INV_X1 us30_U399 (.A( sa30_4 ) , .ZN( us30_n847 ) );
  NAND2_X1 us30_U4 (.A1( us30_n441 ) , .A2( us30_n464 ) , .ZN( us30_n708 ) );
  NOR4_X1 us30_U40 (.A4( us30_n793 ) , .A3( us30_n794 ) , .A2( us30_n795 ) , .A1( us30_n796 ) , .ZN( us30_n797 ) );
  INV_X1 us30_U400 (.A( sa30_3 ) , .ZN( us30_n829 ) );
  INV_X1 us30_U401 (.A( sa30_1 ) , .ZN( us30_n827 ) );
  INV_X1 us30_U402 (.A( sa30_0 ) , .ZN( us30_n826 ) );
  INV_X1 us30_U403 (.A( sa30_2 ) , .ZN( us30_n828 ) );
  INV_X1 us30_U404 (.A( sa30_7 ) , .ZN( us30_n858 ) );
  INV_X1 us30_U405 (.A( sa30_5 ) , .ZN( us30_n848 ) );
  NAND2_X1 us30_U406 (.A2( us30_n461 ) , .A1( us30_n471 ) , .ZN( us30_n697 ) );
  OAI221_X1 us30_U407 (.A( us30_n783 ) , .C2( us30_n784 ) , .B2( us30_n785 ) , .B1( us30_n786 ) , .ZN( us30_n796 ) , .C1( us30_n813 ) );
  NAND2_X1 us30_U408 (.A1( us30_n729 ) , .A2( us30_n784 ) , .ZN( us30_n811 ) );
  OAI22_X1 us30_U409 (.ZN( us30_n588 ) , .A2( us30_n747 ) , .B2( us30_n762 ) , .A1( us30_n763 ) , .B1( us30_n784 ) );
  NOR4_X1 us30_U41 (.A4( us30_n776 ) , .A3( us30_n777 ) , .A1( us30_n778 ) , .ZN( us30_n799 ) , .A2( us30_n801 ) );
  AOI21_X1 us30_U410 (.ZN( us30_n592 ) , .B1( us30_n728 ) , .B2( us30_n784 ) , .A( us30_n790 ) );
  AOI21_X1 us30_U411 (.ZN( us30_n623 ) , .B1( us30_n699 ) , .A( us30_n779 ) , .B2( us30_n784 ) );
  AOI21_X1 us30_U412 (.ZN( us30_n648 ) , .A( us30_n762 ) , .B2( us30_n784 ) , .B1( us30_n792 ) );
  OAI22_X1 us30_U413 (.ZN( us30_n681 ) , .A1( us30_n699 ) , .A2( us30_n730 ) , .B2( us30_n784 ) , .B1( us30_n817 ) );
  OAI21_X1 us30_U414 (.A( us30_n613 ) , .ZN( us30_n616 ) , .B1( us30_n625 ) , .B2( us30_n784 ) );
  NOR2_X1 us30_U415 (.ZN( us30_n610 ) , .A1( us30_n784 ) , .A2( us30_n816 ) );
  OAI222_X1 us30_U416 (.A2( us30_n669 ) , .ZN( us30_n674 ) , .B1( us30_n747 ) , .B2( us30_n784 ) , .C2( us30_n788 ) , .C1( us30_n815 ) , .A1( us30_n817 ) );
  NOR2_X1 us30_U417 (.ZN( us30_n651 ) , .A1( us30_n784 ) , .A2( us30_n788 ) );
  NOR2_X1 us30_U418 (.ZN( us30_n600 ) , .A2( us30_n697 ) , .A1( us30_n784 ) );
  NOR2_X1 us30_U419 (.ZN( us30_n553 ) , .A2( us30_n744 ) , .A1( us30_n784 ) );
  NOR4_X1 us30_U42 (.A3( us30_n755 ) , .A2( us30_n756 ) , .A1( us30_n757 ) , .ZN( us30_n758 ) , .A4( us30_n869 ) );
  INV_X1 us30_U420 (.A( us30_n784 ) , .ZN( us30_n861 ) );
  AOI21_X1 us30_U421 (.ZN( us30_n500 ) , .A( us30_n697 ) , .B1( us30_n708 ) , .B2( us30_n786 ) );
  OAI221_X1 us30_U422 (.A( us30_n696 ) , .ZN( us30_n703 ) , .C2( us30_n784 ) , .C1( us30_n785 ) , .B1( us30_n786 ) , .B2( us30_n806 ) );
  OAI22_X1 us30_U423 (.ZN( us30_n590 ) , .B1( us30_n730 ) , .B2( us30_n749 ) , .A2( us30_n786 ) , .A1( us30_n803 ) );
  NOR2_X1 us30_U424 (.ZN( us30_n612 ) , .A1( us30_n779 ) , .A2( us30_n786 ) );
  NAND2_X1 us30_U425 (.A2( us30_n749 ) , .A1( us30_n786 ) , .ZN( us30_n809 ) );
  OAI222_X1 us30_U426 (.ZN( us30_n617 ) , .B1( us30_n697 ) , .C1( us30_n724 ) , .C2( us30_n747 ) , .B2( us30_n786 ) , .A2( us30_n792 ) , .A1( us30_n816 ) );
  NOR2_X1 us30_U427 (.ZN( us30_n717 ) , .A2( us30_n744 ) , .A1( us30_n786 ) );
  NOR2_X1 us30_U428 (.ZN( us30_n653 ) , .A1( us30_n762 ) , .A2( us30_n786 ) );
  NOR2_X1 us30_U429 (.ZN( us30_n554 ) , .A1( us30_n786 ) , .A2( us30_n813 ) );
  AOI211_X1 us30_U43 (.B( us30_n745 ) , .A( us30_n746 ) , .ZN( us30_n759 ) , .C1( us30_n832 ) , .C2( us30_n853 ) );
  NOR2_X1 us30_U430 (.ZN( us30_n701 ) , .A2( us30_n786 ) , .A1( us30_n817 ) );
  NOR2_X1 us30_U431 (.A1( us30_n730 ) , .ZN( us30_n765 ) , .A2( us30_n786 ) );
  AND2_X1 us30_U432 (.ZN( us30_n438 ) , .A2( us30_n831 ) , .A1( us30_n854 ) );
  AND2_X1 us30_U433 (.ZN( us30_n439 ) , .A2( us30_n843 ) , .A1( us30_n861 ) );
  NOR3_X1 us30_U434 (.A1( us30_n438 ) , .A2( us30_n439 ) , .A3( us30_n576 ) , .ZN( us30_n587 ) );
  NAND4_X1 us30_U435 (.ZN( sa31_sr_2 ) , .A4( us30_n643 ) , .A3( us30_n644 ) , .A2( us30_n645 ) , .A1( us30_n646 ) );
  INV_X1 us30_U436 (.A( us30_n812 ) , .ZN( us30_n854 ) );
  NAND3_X1 us30_U437 (.ZN( sa31_sr_6 ) , .A3( us30_n797 ) , .A2( us30_n798 ) , .A1( us30_n799 ) );
  NAND3_X1 us30_U438 (.ZN( sa31_sr_5 ) , .A3( us30_n758 ) , .A2( us30_n759 ) , .A1( us30_n760 ) );
  NAND3_X1 us30_U439 (.ZN( sa31_sr_4 ) , .A3( us30_n738 ) , .A2( us30_n739 ) , .A1( us30_n740 ) );
  NOR3_X1 us30_U44 (.A3( us30_n741 ) , .A2( us30_n742 ) , .A1( us30_n743 ) , .ZN( us30_n760 ) );
  NAND3_X1 us30_U440 (.A3( us30_n675 ) , .A2( us30_n676 ) , .A1( us30_n677 ) , .ZN( us30_n807 ) );
  NAND3_X1 us30_U441 (.ZN( us30_n638 ) , .A3( us30_n708 ) , .A2( us30_n724 ) , .A1( us30_n792 ) );
  NAND3_X1 us30_U442 (.A3( us30_n618 ) , .A2( us30_n619 ) , .A1( us30_n620 ) , .ZN( us30_n725 ) );
  NAND3_X1 us30_U443 (.A3( us30_n585 ) , .A2( us30_n586 ) , .A1( us30_n587 ) , .ZN( us30_n621 ) );
  NAND3_X1 us30_U444 (.ZN( us30_n565 ) , .A3( us30_n680 ) , .A2( us30_n750 ) , .A1( us30_n785 ) );
  NAND3_X1 us30_U445 (.A3( us30_n523 ) , .A2( us30_n524 ) , .A1( us30_n525 ) , .ZN( us30_n742 ) );
  NAND3_X1 us30_U446 (.A3( us30_n512 ) , .A1( us30_n513 ) , .ZN( us30_n608 ) , .A2( us30_n871 ) );
  NAND3_X1 us30_U447 (.A3( us30_n467 ) , .A2( us30_n468 ) , .A1( us30_n469 ) , .ZN( us30_n777 ) );
  INV_X1 us30_U448 (.A( us30_n803 ) , .ZN( us30_n843 ) );
  AOI21_X1 us30_U449 (.ZN( us30_n576 ) , .B2( us30_n724 ) , .B1( us30_n748 ) , .A( us30_n785 ) );
  NAND4_X1 us30_U45 (.ZN( sa31_sr_3 ) , .A4( us30_n704 ) , .A3( us30_n705 ) , .A2( us30_n706 ) , .A1( us30_n707 ) );
  NOR4_X1 us30_U46 (.A4( us30_n700 ) , .A3( us30_n701 ) , .A2( us30_n702 ) , .A1( us30_n703 ) , .ZN( us30_n704 ) );
  AOI211_X1 us30_U47 (.B( us30_n694 ) , .A( us30_n695 ) , .ZN( us30_n705 ) , .C2( us30_n831 ) , .C1( us30_n851 ) );
  NOR2_X1 us30_U48 (.ZN( us30_n707 ) , .A2( us30_n776 ) , .A1( us30_n800 ) );
  AOI222_X1 us30_U49 (.B2( us30_n638 ) , .ZN( us30_n644 ) , .B1( us30_n841 ) , .A1( us30_n842 ) , .C2( us30_n846 ) , .C1( us30_n863 ) , .A2( us30_n865 ) );
  NAND2_X1 us30_U5 (.A2( us30_n441 ) , .A1( us30_n452 ) , .ZN( us30_n791 ) );
  NOR4_X1 us30_U50 (.A4( us30_n639 ) , .A3( us30_n640 ) , .A2( us30_n641 ) , .A1( us30_n642 ) , .ZN( us30_n643 ) );
  NOR3_X1 us30_U51 (.A2( us30_n607 ) , .A1( us30_n608 ) , .ZN( us30_n646 ) , .A3( us30_n722 ) );
  NOR2_X1 us30_U52 (.ZN( us30_n804 ) , .A1( us30_n854 ) , .A2( us30_n861 ) );
  NAND4_X1 us30_U53 (.ZN( sa31_sr_7 ) , .A4( us30_n822 ) , .A3( us30_n823 ) , .A2( us30_n824 ) , .A1( us30_n825 ) );
  NOR4_X1 us30_U54 (.A4( us30_n818 ) , .A3( us30_n819 ) , .A2( us30_n820 ) , .A1( us30_n821 ) , .ZN( us30_n822 ) );
  AOI222_X1 us30_U55 (.C2( us30_n809 ) , .B2( us30_n810 ) , .A2( us30_n811 ) , .ZN( us30_n823 ) , .C1( us30_n832 ) , .A1( us30_n839 ) , .B1( us30_n853 ) );
  AOI211_X1 us30_U56 (.B( us30_n807 ) , .A( us30_n808 ) , .ZN( us30_n824 ) , .C1( us30_n842 ) , .C2( us30_n850 ) );
  NAND4_X1 us30_U57 (.ZN( sa31_sr_0 ) , .A4( us30_n501 ) , .A3( us30_n502 ) , .A2( us30_n503 ) , .A1( us30_n504 ) );
  AOI221_X1 us30_U58 (.A( us30_n497 ) , .ZN( us30_n502 ) , .B2( us30_n843 ) , .C1( us30_n846 ) , .C2( us30_n860 ) , .B1( us30_n862 ) );
  NOR4_X1 us30_U59 (.A4( us30_n498 ) , .A3( us30_n499 ) , .A2( us30_n500 ) , .ZN( us30_n501 ) , .A1( us30_n527 ) );
  NAND2_X1 us30_U6 (.A2( us30_n471 ) , .A1( us30_n472 ) , .ZN( us30_n817 ) );
  AOI211_X1 us30_U60 (.A( us30_n496 ) , .ZN( us30_n503 ) , .B( us30_n802 ) , .C2( us30_n839 ) , .C1( us30_n851 ) );
  NAND4_X1 us30_U61 (.ZN( sa31_sr_1 ) , .A4( us30_n595 ) , .A3( us30_n596 ) , .A2( us30_n597 ) , .A1( us30_n598 ) );
  NOR4_X1 us30_U62 (.A4( us30_n591 ) , .A3( us30_n592 ) , .A2( us30_n593 ) , .A1( us30_n594 ) , .ZN( us30_n595 ) );
  AOI211_X1 us30_U63 (.B( us30_n589 ) , .A( us30_n590 ) , .ZN( us30_n596 ) , .C2( us30_n811 ) , .C1( us30_n833 ) );
  AOI211_X1 us30_U64 (.A( us30_n588 ) , .ZN( us30_n597 ) , .B( us30_n621 ) , .C1( us30_n845 ) , .C2( us30_n855 ) );
  NOR2_X1 us30_U65 (.ZN( us30_n748 ) , .A1( us30_n861 ) , .A2( us30_n862 ) );
  NOR2_X1 us30_U66 (.ZN( us30_n625 ) , .A2( us30_n836 ) , .A1( us30_n839 ) );
  NAND4_X1 us30_U67 (.A4( us30_n603 ) , .A3( us30_n604 ) , .A2( us30_n605 ) , .A1( us30_n606 ) , .ZN( us30_n722 ) );
  NOR3_X1 us30_U68 (.A1( us30_n599 ) , .ZN( us30_n604 ) , .A3( us30_n663 ) , .A2( us30_n770 ) );
  NOR4_X1 us30_U69 (.A3( us30_n600 ) , .A2( us30_n601 ) , .A1( us30_n602 ) , .ZN( us30_n603 ) , .A4( us30_n655 ) );
  NOR3_X1 us30_U7 (.ZN( us30_n598 ) , .A1( us30_n608 ) , .A3( us30_n723 ) , .A2( us30_n742 ) );
  AOI222_X1 us30_U70 (.ZN( us30_n606 ) , .A1( us30_n830 ) , .C2( us30_n837 ) , .B1( us30_n842 ) , .A2( us30_n856 ) , .B2( us30_n861 ) , .C1( us30_n868 ) );
  NAND4_X1 us30_U71 (.A4( us30_n657 ) , .A3( us30_n658 ) , .A2( us30_n659 ) , .A1( us30_n660 ) , .ZN( us30_n800 ) );
  NOR3_X1 us30_U72 (.A3( us30_n648 ) , .A2( us30_n649 ) , .A1( us30_n650 ) , .ZN( us30_n659 ) );
  NOR3_X1 us30_U73 (.A3( us30_n651 ) , .A2( us30_n652 ) , .A1( us30_n653 ) , .ZN( us30_n658 ) );
  NOR3_X1 us30_U74 (.A3( us30_n654 ) , .A2( us30_n655 ) , .A1( us30_n656 ) , .ZN( us30_n657 ) );
  NAND4_X1 us30_U75 (.A4( us30_n560 ) , .A3( us30_n561 ) , .A2( us30_n562 ) , .A1( us30_n563 ) , .ZN( us30_n607 ) );
  NOR4_X1 us30_U76 (.ZN( us30_n561 ) , .A1( us30_n653 ) , .A3( us30_n661 ) , .A4( us30_n685 ) , .A2( us30_n768 ) );
  NOR4_X1 us30_U77 (.A4( us30_n552 ) , .A3( us30_n553 ) , .A2( us30_n554 ) , .A1( us30_n555 ) , .ZN( us30_n562 ) );
  NOR4_X1 us30_U78 (.A4( us30_n556 ) , .A3( us30_n557 ) , .A2( us30_n558 ) , .A1( us30_n559 ) , .ZN( us30_n560 ) );
  NAND4_X1 us30_U79 (.A4( us30_n772 ) , .A3( us30_n773 ) , .A2( us30_n774 ) , .A1( us30_n775 ) , .ZN( us30_n801 ) );
  NOR3_X1 us30_U8 (.A3( us30_n800 ) , .A2( us30_n801 ) , .A1( us30_n802 ) , .ZN( us30_n825 ) );
  NOR3_X1 us30_U80 (.A3( us30_n765 ) , .A2( us30_n766 ) , .A1( us30_n767 ) , .ZN( us30_n773 ) );
  NOR4_X1 us30_U81 (.A4( us30_n768 ) , .A3( us30_n769 ) , .A2( us30_n770 ) , .A1( us30_n771 ) , .ZN( us30_n772 ) );
  AOI222_X1 us30_U82 (.ZN( us30_n775 ) , .A1( us30_n830 ) , .C1( us30_n834 ) , .B2( us30_n841 ) , .A2( us30_n850 ) , .B1( us30_n861 ) , .C2( us30_n873 ) );
  NOR4_X1 us30_U83 (.A4( us30_n665 ) , .A3( us30_n666 ) , .A2( us30_n667 ) , .A1( us30_n668 ) , .ZN( us30_n676 ) );
  NOR4_X1 us30_U84 (.A4( us30_n661 ) , .A3( us30_n662 ) , .A2( us30_n663 ) , .A1( us30_n664 ) , .ZN( us30_n677 ) );
  NOR4_X1 us30_U85 (.A3( us30_n673 ) , .A1( us30_n674 ) , .ZN( us30_n675 ) , .A4( us30_n715 ) , .A2( us30_n859 ) );
  NOR2_X1 us30_U86 (.ZN( us30_n761 ) , .A1( us30_n833 ) , .A2( us30_n834 ) );
  NOR4_X1 us30_U87 (.A4( us30_n577 ) , .A3( us30_n578 ) , .A2( us30_n579 ) , .ZN( us30_n586 ) , .A1( us30_n683 ) );
  NOR4_X1 us30_U88 (.A1( us30_n584 ) , .ZN( us30_n585 ) , .A3( us30_n652 ) , .A2( us30_n662 ) , .A4( us30_n767 ) );
  AOI222_X1 us30_U89 (.ZN( us30_n513 ) , .C1( us30_n832 ) , .B2( us30_n837 ) , .A2( us30_n843 ) , .C2( us30_n862 ) , .B1( us30_n863 ) , .A1( us30_n866 ) );
  NOR3_X1 us30_U9 (.A3( us30_n621 ) , .A2( us30_n622 ) , .ZN( us30_n636 ) , .A1( us30_n725 ) );
  NOR4_X1 us30_U90 (.A4( us30_n509 ) , .A2( us30_n510 ) , .A1( us30_n511 ) , .ZN( us30_n512 ) , .A3( us30_n670 ) );
  INV_X1 us30_U91 (.A( us30_n505 ) , .ZN( us30_n871 ) );
  NAND4_X1 us30_U92 (.A4( us30_n456 ) , .A3( us30_n457 ) , .A2( us30_n458 ) , .A1( us30_n459 ) , .ZN( us30_n679 ) );
  NOR3_X1 us30_U93 (.ZN( us30_n457 ) , .A3( us30_n530 ) , .A1( us30_n555 ) , .A2( us30_n570 ) );
  AOI221_X1 us30_U94 (.A( us30_n450 ) , .ZN( us30_n459 ) , .C2( us30_n753 ) , .B1( us30_n832 ) , .C1( us30_n842 ) , .B2( us30_n861 ) );
  NOR4_X1 us30_U95 (.ZN( us30_n458 ) , .A2( us30_n509 ) , .A1( us30_n599 ) , .A4( us30_n628 ) , .A3( us30_n711 ) );
  NAND4_X1 us30_U96 (.A4( us30_n535 ) , .A3( us30_n536 ) , .A2( us30_n537 ) , .A1( us30_n538 ) , .ZN( us30_n622 ) );
  NOR4_X1 us30_U97 (.A4( us30_n526 ) , .A2( us30_n527 ) , .A1( us30_n528 ) , .ZN( us30_n538 ) , .A3( us30_n701 ) );
  NOR4_X1 us30_U98 (.A1( us30_n531 ) , .ZN( us30_n536 ) , .A2( us30_n654 ) , .A4( us30_n668 ) , .A3( us30_n765 ) );
  NOR4_X1 us30_U99 (.A4( us30_n529 ) , .A3( us30_n530 ) , .ZN( us30_n537 ) , .A2( us30_n684 ) , .A1( us30_n794 ) );
  NOR2_X1 us32_U10 (.A1( us32_n678 ) , .ZN( us32_n693 ) , .A2( us32_n807 ) );
  AOI211_X1 us32_U100 (.B( us32_n477 ) , .A( us32_n478 ) , .ZN( us32_n482 ) , .C2( us32_n833 ) , .C1( us32_n861 ) );
  NOR4_X1 us32_U101 (.ZN( us32_n481 ) , .A3( us32_n532 ) , .A4( us32_n545 ) , .A2( us32_n567 ) , .A1( us32_n717 ) );
  NAND4_X1 us32_U102 (.A4( us32_n548 ) , .A3( us32_n549 ) , .A2( us32_n550 ) , .A1( us32_n551 ) , .ZN( us32_n745 ) );
  NOR3_X1 us32_U103 (.ZN( us32_n549 ) , .A2( us32_n651 ) , .A1( us32_n667 ) , .A3( us32_n771 ) );
  AOI211_X1 us32_U104 (.B( us32_n539 ) , .A( us32_n540 ) , .ZN( us32_n551 ) , .C2( us32_n839 ) , .C1( us32_n851 ) );
  NOR4_X1 us32_U105 (.A4( us32_n541 ) , .A3( us32_n542 ) , .A2( us32_n543 ) , .ZN( us32_n550 ) , .A1( us32_n688 ) );
  NOR4_X1 us32_U106 (.ZN( us32_n620 ) , .A1( us32_n656 ) , .A3( us32_n666 ) , .A4( us32_n682 ) , .A2( us32_n766 ) );
  NOR4_X1 us32_U107 (.A4( us32_n609 ) , .A3( us32_n610 ) , .A2( us32_n611 ) , .A1( us32_n612 ) , .ZN( us32_n619 ) );
  NOR4_X1 us32_U108 (.A4( us32_n614 ) , .A3( us32_n615 ) , .A2( us32_n616 ) , .A1( us32_n617 ) , .ZN( us32_n618 ) );
  NOR2_X1 us32_U109 (.ZN( us32_n686 ) , .A1( us32_n831 ) , .A2( us32_n832 ) );
  NOR3_X1 us32_U11 (.ZN( us32_n504 ) , .A2( us32_n679 ) , .A3( us32_n777 ) , .A1( us32_n876 ) );
  NAND4_X1 us32_U110 (.A4( us32_n485 ) , .A3( us32_n486 ) , .A2( us32_n487 ) , .A1( us32_n488 ) , .ZN( us32_n778 ) );
  NOR4_X1 us32_U111 (.A4( us32_n484 ) , .ZN( us32_n487 ) , .A1( us32_n566 ) , .A2( us32_n581 ) , .A3( us32_n602 ) );
  NOR4_X1 us32_U112 (.ZN( us32_n486 ) , .A1( us32_n507 ) , .A2( us32_n519 ) , .A4( us32_n546 ) , .A3( us32_n611 ) );
  NOR4_X1 us32_U113 (.ZN( us32_n485 ) , .A2( us32_n533 ) , .A1( us32_n558 ) , .A3( us32_n631 ) , .A4( us32_n718 ) );
  NAND4_X1 us32_U114 (.A4( us32_n691 ) , .A3( us32_n692 ) , .A1( us32_n693 ) , .ZN( us32_n776 ) , .A2( us32_n872 ) );
  AOI221_X1 us32_U115 (.A( us32_n681 ) , .ZN( us32_n692 ) , .B2( us32_n840 ) , .C1( us32_n842 ) , .C2( us32_n862 ) , .B1( us32_n865 ) );
  INV_X1 us32_U116 (.A( us32_n679 ) , .ZN( us32_n872 ) );
  NOR4_X1 us32_U117 (.A4( us32_n687 ) , .A3( us32_n688 ) , .A2( us32_n689 ) , .A1( us32_n690 ) , .ZN( us32_n691 ) );
  NAND4_X1 us32_U118 (.A4( us32_n473 ) , .A3( us32_n474 ) , .A2( us32_n475 ) , .A1( us32_n476 ) , .ZN( us32_n678 ) );
  NOR4_X1 us32_U119 (.ZN( us32_n475 ) , .A1( us32_n531 ) , .A3( us32_n568 ) , .A4( us32_n600 ) , .A2( us32_n642 ) );
  INV_X1 us32_U12 (.A( us32_n706 ) , .ZN( us32_n876 ) );
  NOR4_X1 us32_U120 (.A4( us32_n470 ) , .ZN( us32_n476 ) , .A3( us32_n556 ) , .A1( us32_n735 ) , .A2( us32_n755 ) );
  NOR4_X1 us32_U121 (.ZN( us32_n473 ) , .A2( us32_n521 ) , .A4( us32_n594 ) , .A1( us32_n609 ) , .A3( us32_n629 ) );
  NAND4_X1 us32_U122 (.A4( us32_n719 ) , .A3( us32_n720 ) , .A2( us32_n721 ) , .ZN( us32_n741 ) , .A1( us32_n857 ) );
  INV_X1 us32_U123 (.A( us32_n709 ) , .ZN( us32_n857 ) );
  AOI221_X1 us32_U124 (.A( us32_n710 ) , .ZN( us32_n721 ) , .C2( us32_n844 ) , .B2( us32_n845 ) , .C1( us32_n861 ) , .B1( us32_n862 ) );
  NOR4_X1 us32_U125 (.A4( us32_n715 ) , .A3( us32_n716 ) , .A2( us32_n717 ) , .A1( us32_n718 ) , .ZN( us32_n719 ) );
  NOR2_X1 us32_U126 (.ZN( us32_n733 ) , .A2( us32_n832 ) , .A1( us32_n845 ) );
  NOR2_X1 us32_U127 (.ZN( us32_n789 ) , .A2( us32_n862 ) , .A1( us32_n868 ) );
  NAND4_X1 us32_U128 (.A4( us32_n573 ) , .A3( us32_n574 ) , .A1( us32_n575 ) , .ZN( us32_n723 ) , .A2( us32_n874 ) );
  AOI221_X1 us32_U129 (.A( us32_n564 ) , .C2( us32_n565 ) , .ZN( us32_n574 ) , .B2( us32_n845 ) , .B1( us32_n852 ) , .C1( us32_n853 ) );
  INV_X1 us32_U13 (.A( us32_n607 ) , .ZN( us32_n874 ) );
  NOR4_X1 us32_U130 (.A4( us32_n569 ) , .A3( us32_n570 ) , .A2( us32_n571 ) , .A1( us32_n572 ) , .ZN( us32_n573 ) );
  NOR2_X1 us32_U131 (.ZN( us32_n575 ) , .A1( us32_n622 ) , .A2( us32_n745 ) );
  NOR2_X1 us32_U132 (.ZN( us32_n748 ) , .A1( us32_n861 ) , .A2( us32_n862 ) );
  NAND4_X1 us32_U133 (.A4( us32_n633 ) , .A3( us32_n634 ) , .A2( us32_n635 ) , .A1( us32_n636 ) , .ZN( us32_n743 ) );
  AOI211_X1 us32_U134 (.B( us32_n623 ) , .A( us32_n624 ) , .ZN( us32_n635 ) , .C2( us32_n836 ) , .C1( us32_n863 ) );
  NOR4_X1 us32_U135 (.A4( us32_n629 ) , .A3( us32_n630 ) , .A2( us32_n631 ) , .A1( us32_n632 ) , .ZN( us32_n633 ) );
  NOR4_X1 us32_U136 (.A4( us32_n626 ) , .A3( us32_n627 ) , .A2( us32_n628 ) , .ZN( us32_n634 ) , .A1( us32_n664 ) );
  NAND4_X1 us32_U137 (.A4( us32_n493 ) , .A3( us32_n494 ) , .A1( us32_n495 ) , .ZN( us32_n802 ) , .A2( us32_n867 ) );
  AOI221_X1 us32_U138 (.A( us32_n489 ) , .ZN( us32_n494 ) , .B2( us32_n836 ) , .C2( us32_n841 ) , .C1( us32_n851 ) , .B1( us32_n860 ) );
  INV_X1 us32_U139 (.A( us32_n778 ) , .ZN( us32_n867 ) );
  INV_X1 us32_U14 (.A( us32_n680 ) , .ZN( us32_n840 ) );
  NOR4_X1 us32_U140 (.A2( us32_n491 ) , .A1( us32_n492 ) , .ZN( us32_n493 ) , .A3( us32_n580 ) , .A4( us32_n612 ) );
  NOR4_X1 us32_U141 (.A4( us32_n734 ) , .A3( us32_n735 ) , .A2( us32_n736 ) , .A1( us32_n737 ) , .ZN( us32_n738 ) );
  AOI211_X1 us32_U142 (.B( us32_n725 ) , .A( us32_n726 ) , .ZN( us32_n739 ) , .C1( us32_n843 ) , .C2( us32_n855 ) );
  NOR3_X1 us32_U143 (.A3( us32_n722 ) , .A1( us32_n723 ) , .ZN( us32_n740 ) , .A2( us32_n741 ) );
  NOR2_X1 us32_U144 (.ZN( us32_n647 ) , .A1( us32_n854 ) , .A2( us32_n868 ) );
  INV_X1 us32_U145 (.A( us32_n762 ) , .ZN( us32_n830 ) );
  INV_X1 us32_U146 (.A( us32_n754 ) , .ZN( us32_n869 ) );
  OAI21_X1 us32_U147 (.B1( us32_n753 ) , .ZN( us32_n754 ) , .A( us32_n845 ) , .B2( us32_n868 ) );
  INV_X1 us32_U148 (.A( us32_n697 ) , .ZN( us32_n838 ) );
  OR4_X1 us32_U149 (.ZN( us32_n492 ) , .A4( us32_n534 ) , .A2( us32_n547 ) , .A1( us32_n559 ) , .A3( us32_n632 ) );
  NOR4_X1 us32_U15 (.A4( us32_n445 ) , .A3( us32_n446 ) , .A2( us32_n516 ) , .A1( us32_n541 ) , .ZN( us32_n706 ) );
  OR4_X1 us32_U150 (.A4( us32_n566 ) , .A3( us32_n567 ) , .A2( us32_n568 ) , .ZN( us32_n572 ) , .A1( us32_n665 ) );
  OR4_X1 us32_U151 (.A4( us32_n682 ) , .A3( us32_n683 ) , .A2( us32_n684 ) , .A1( us32_n685 ) , .ZN( us32_n690 ) );
  OR4_X1 us32_U152 (.ZN( us32_n466 ) , .A4( us32_n518 ) , .A3( us32_n529 ) , .A2( us32_n578 ) , .A1( us32_n712 ) );
  OR4_X1 us32_U153 (.A4( us32_n518 ) , .A2( us32_n519 ) , .A1( us32_n520 ) , .ZN( us32_n522 ) , .A3( us32_n821 ) );
  OR4_X1 us32_U154 (.A4( us32_n580 ) , .A3( us32_n581 ) , .A2( us32_n582 ) , .A1( us32_n583 ) , .ZN( us32_n584 ) );
  NAND2_X1 us32_U155 (.ZN( us32_n613 ) , .A2( us32_n837 ) , .A1( us32_n873 ) );
  OR3_X1 us32_U156 (.A3( us32_n506 ) , .A2( us32_n507 ) , .A1( us32_n508 ) , .ZN( us32_n511 ) );
  INV_X1 us32_U157 (.A( us32_n672 ) , .ZN( us32_n859 ) );
  AOI21_X1 us32_U158 (.A( us32_n670 ) , .B1( us32_n671 ) , .ZN( us32_n672 ) , .B2( us32_n856 ) );
  INV_X1 us32_U159 (.A( us32_n463 ) , .ZN( us32_n864 ) );
  OR3_X1 us32_U16 (.ZN( us32_n446 ) , .A1( us32_n528 ) , .A3( us32_n577 ) , .A2( us32_n875 ) );
  OAI21_X1 us32_U160 (.ZN( us32_n463 ) , .B1( us32_n809 ) , .A( us32_n834 ) , .B2( us32_n851 ) );
  OAI222_X1 us32_U161 (.B2( us32_n708 ) , .ZN( us32_n709 ) , .C2( us32_n724 ) , .B1( us32_n747 ) , .A1( us32_n806 ) , .C1( us32_n814 ) , .A2( us32_n815 ) );
  NAND2_X1 us32_U162 (.A1( us32_n447 ) , .A2( us32_n465 ) , .ZN( us32_n749 ) );
  AOI22_X1 us32_U163 (.A2( us32_n782 ) , .ZN( us32_n783 ) , .B2( us32_n831 ) , .A1( us32_n834 ) , .B1( us32_n863 ) );
  AOI22_X1 us32_U164 (.ZN( us32_n696 ) , .A1( us32_n830 ) , .B2( us32_n843 ) , .A2( us32_n865 ) , .B1( us32_n868 ) );
  INV_X1 us32_U165 (.A( us32_n730 ) , .ZN( us32_n839 ) );
  AOI221_X1 us32_U166 (.A( us32_n483 ) , .ZN( us32_n488 ) , .B1( us32_n831 ) , .C2( us32_n844 ) , .C1( us32_n852 ) , .B2( us32_n862 ) );
  OAI22_X1 us32_U167 (.ZN( us32_n483 ) , .A1( us32_n708 ) , .B2( us32_n785 ) , .A2( us32_n806 ) , .B1( us32_n812 ) );
  INV_X1 us32_U168 (.A( us32_n790 ) , .ZN( us32_n832 ) );
  OAI221_X1 us32_U169 (.A( us32_n727 ) , .C2( us32_n728 ) , .B2( us32_n729 ) , .B1( us32_n730 ) , .ZN( us32_n737 ) , .C1( us32_n817 ) );
  OR4_X1 us32_U17 (.A4( us32_n442 ) , .A2( us32_n443 ) , .A1( us32_n444 ) , .ZN( us32_n445 ) , .A3( us32_n553 ) );
  AOI22_X1 us32_U170 (.ZN( us32_n727 ) , .B1( us32_n832 ) , .A2( us32_n838 ) , .A1( us32_n863 ) , .B2( us32_n866 ) );
  NAND2_X1 us32_U171 (.A1( us32_n451 ) , .A2( us32_n453 ) , .ZN( us32_n762 ) );
  INV_X1 us32_U172 (.A( us32_n786 ) , .ZN( us32_n862 ) );
  OAI22_X1 us32_U173 (.ZN( us32_n710 ) , .A2( us32_n728 ) , .B2( us32_n729 ) , .A1( us32_n744 ) , .B1( us32_n813 ) );
  INV_X1 us32_U174 (.A( us32_n816 ) , .ZN( us32_n831 ) );
  OAI22_X1 us32_U175 (.ZN( us32_n489 ) , .A1( us32_n724 ) , .B2( us32_n728 ) , .B1( us32_n730 ) , .A2( us32_n779 ) );
  OAI22_X1 us32_U176 (.ZN( us32_n624 ) , .B1( us32_n669 ) , .B2( us32_n747 ) , .A1( us32_n815 ) , .A2( us32_n816 ) );
  INV_X1 us32_U177 (.A( us32_n788 ) , .ZN( us32_n845 ) );
  OAI22_X1 us32_U178 (.A1( us32_n724 ) , .ZN( us32_n726 ) , .B2( us32_n750 ) , .B1( us32_n812 ) , .A2( us32_n816 ) );
  INV_X1 us32_U179 (.A( us32_n744 ) , .ZN( us32_n837 ) );
  INV_X1 us32_U18 (.A( us32_n613 ) , .ZN( us32_n875 ) );
  OAI22_X1 us32_U180 (.B2( us32_n779 ) , .B1( us32_n780 ) , .ZN( us32_n781 ) , .A2( us32_n814 ) , .A1( us32_n815 ) );
  INV_X1 us32_U181 (.A( us32_n814 ) , .ZN( us32_n833 ) );
  INV_X1 us32_U182 (.A( us32_n669 ) , .ZN( us32_n865 ) );
  OAI22_X1 us32_U183 (.B2( us32_n744 ) , .ZN( us32_n746 ) , .A2( us32_n762 ) , .B1( us32_n780 ) , .A1( us32_n792 ) );
  OAI22_X1 us32_U184 (.ZN( us32_n496 ) , .A2( us32_n744 ) , .A1( us32_n780 ) , .B1( us32_n791 ) , .B2( us32_n806 ) );
  AOI211_X1 us32_U185 (.A( us32_n637 ) , .ZN( us32_n645 ) , .B( us32_n743 ) , .C2( us32_n839 ) , .C1( us32_n854 ) );
  OAI22_X1 us32_U186 (.ZN( us32_n637 ) , .A1( us32_n699 ) , .B2( us32_n728 ) , .A2( us32_n762 ) , .B1( us32_n816 ) );
  INV_X1 us32_U187 (.A( us32_n750 ) , .ZN( us32_n842 ) );
  OAI22_X1 us32_U188 (.B1( us32_n490 ) , .ZN( us32_n491 ) , .A1( us32_n686 ) , .A2( us32_n763 ) , .B2( us32_n817 ) );
  NOR3_X1 us32_U189 (.ZN( us32_n490 ) , .A1( us32_n782 ) , .A2( us32_n850 ) , .A3( us32_n863 ) );
  INV_X1 us32_U19 (.A( us32_n749 ) , .ZN( us32_n863 ) );
  OAI22_X1 us32_U190 (.ZN( us32_n695 ) , .A2( us32_n730 ) , .A1( us32_n780 ) , .B1( us32_n791 ) , .B2( us32_n817 ) );
  NOR2_X1 us32_U191 (.ZN( us32_n666 ) , .A1( us32_n728 ) , .A2( us32_n803 ) );
  NOR2_X1 us32_U192 (.ZN( us32_n594 ) , .A2( us32_n697 ) , .A1( us32_n728 ) );
  NOR2_X1 us32_U193 (.ZN( us32_n570 ) , .A1( us32_n728 ) , .A2( us32_n806 ) );
  NOR2_X1 us32_U194 (.ZN( us32_n654 ) , .A1( us32_n728 ) , .A2( us32_n813 ) );
  NOR2_X1 us32_U195 (.ZN( us32_n546 ) , .A2( us32_n780 ) , .A1( us32_n814 ) );
  NOR2_X1 us32_U196 (.ZN( us32_n532 ) , .A2( us32_n749 ) , .A1( us32_n750 ) );
  NOR2_X1 us32_U197 (.ZN( us32_n577 ) , .A2( us32_n699 ) , .A1( us32_n814 ) );
  NOR2_X1 us32_U198 (.ZN( us32_n615 ) , .A1( us32_n785 ) , .A2( us32_n815 ) );
  NOR2_X1 us32_U199 (.ZN( us32_n629 ) , .A2( us32_n728 ) , .A1( us32_n785 ) );
  AOI222_X1 us32_U20 (.ZN( us32_n605 ) , .B2( us32_n671 ) , .B1( us32_n753 ) , .C2( us32_n831 ) , .A1( us32_n833 ) , .A2( us32_n862 ) , .C1( us32_n863 ) );
  NOR2_X1 us32_U200 (.ZN( us32_n718 ) , .A2( us32_n724 ) , .A1( us32_n744 ) );
  NOR2_X1 us32_U201 (.ZN( us32_n628 ) , .A2( us32_n669 ) , .A1( us32_n785 ) );
  INV_X1 us32_U202 (.A( us32_n728 ) , .ZN( us32_n852 ) );
  NOR2_X1 us32_U203 (.A2( us32_n744 ) , .ZN( us32_n769 ) , .A1( us32_n812 ) );
  NOR2_X1 us32_U204 (.ZN( us32_n531 ) , .A2( us32_n780 ) , .A1( us32_n816 ) );
  NOR2_X1 us32_U205 (.A2( us32_n708 ) , .A1( us32_n750 ) , .ZN( us32_n771 ) );
  NOR2_X1 us32_U206 (.ZN( us32_n599 ) , .A2( us32_n791 ) , .A1( us32_n816 ) );
  NOR2_X1 us32_U207 (.ZN( us32_n611 ) , .A2( us32_n780 ) , .A1( us32_n806 ) );
  NOR2_X1 us32_U208 (.ZN( us32_n652 ) , .A1( us32_n669 ) , .A2( us32_n814 ) );
  INV_X1 us32_U209 (.A( us32_n792 ) , .ZN( us32_n851 ) );
  AOI222_X1 us32_U21 (.ZN( us32_n563 ) , .B1( us32_n830 ) , .C1( us32_n841 ) , .A2( us32_n843 ) , .A1( us32_n854 ) , .B2( us32_n863 ) , .C2( us32_n873 ) );
  NOR2_X1 us32_U210 (.A1( us32_n699 ) , .ZN( us32_n768 ) , .A2( us32_n813 ) );
  NOR2_X1 us32_U211 (.A1( us32_n669 ) , .ZN( us32_n673 ) , .A2( us32_n744 ) );
  NOR2_X1 us32_U212 (.ZN( us32_n541 ) , .A2( us32_n697 ) , .A1( us32_n699 ) );
  NOR2_X1 us32_U213 (.ZN( us32_n602 ) , .A1( us32_n669 ) , .A2( us32_n803 ) );
  NOR2_X1 us32_U214 (.A1( us32_n669 ) , .ZN( us32_n688 ) , .A2( us32_n816 ) );
  NOR2_X1 us32_U215 (.ZN( us32_n667 ) , .A1( us32_n750 ) , .A2( us32_n815 ) );
  NOR2_X1 us32_U216 (.ZN( us32_n555 ) , .A1( us32_n750 ) , .A2( us32_n791 ) );
  NOR2_X1 us32_U217 (.ZN( us32_n508 ) , .A2( us32_n780 ) , .A1( us32_n785 ) );
  NOR2_X1 us32_U218 (.ZN( us32_n543 ) , .A2( us32_n708 ) , .A1( us32_n785 ) );
  INV_X1 us32_U219 (.A( us32_n747 ) , .ZN( us32_n834 ) );
  AOI222_X1 us32_U22 (.ZN( us32_n660 ) , .A2( us32_n839 ) , .B1( us32_n841 ) , .C2( us32_n845 ) , .A1( us32_n860 ) , .C1( us32_n863 ) , .B2( us32_n870 ) );
  NOR2_X1 us32_U220 (.ZN( us32_n664 ) , .A1( us32_n785 ) , .A2( us32_n791 ) );
  NOR2_X1 us32_U221 (.A1( us32_n669 ) , .ZN( us32_n766 ) , .A2( us32_n813 ) );
  NOR2_X1 us32_U222 (.ZN( us32_n527 ) , .A1( us32_n669 ) , .A2( us32_n779 ) );
  NOR2_X1 us32_U223 (.ZN( us32_n661 ) , .A1( us32_n729 ) , .A2( us32_n790 ) );
  NOR2_X1 us32_U224 (.ZN( us32_n601 ) , .A2( us32_n780 ) , .A1( us32_n803 ) );
  NOR2_X1 us32_U225 (.ZN( us32_n507 ) , .A1( us32_n812 ) , .A2( us32_n817 ) );
  NOR2_X1 us32_U226 (.ZN( us32_n528 ) , .A2( us32_n724 ) , .A1( us32_n803 ) );
  NOR2_X1 us32_U227 (.ZN( us32_n509 ) , .A1( us32_n729 ) , .A2( us32_n779 ) );
  NOR2_X1 us32_U228 (.ZN( us32_n557 ) , .A1( us32_n792 ) , .A2( us32_n814 ) );
  NOR2_X1 us32_U229 (.ZN( us32_n545 ) , .A1( us32_n749 ) , .A2( us32_n814 ) );
  INV_X1 us32_U23 (.A( us32_n647 ) , .ZN( us32_n870 ) );
  OAI22_X1 us32_U230 (.B1( us32_n440 ) , .ZN( us32_n444 ) , .A2( us32_n728 ) , .A1( us32_n744 ) , .B2( us32_n749 ) );
  NOR3_X1 us32_U231 (.ZN( us32_n440 ) , .A2( us32_n836 ) , .A3( us32_n837 ) , .A1( us32_n846 ) );
  NOR2_X1 us32_U232 (.ZN( us32_n662 ) , .A2( us32_n697 ) , .A1( us32_n729 ) );
  OAI22_X1 us32_U233 (.B2( us32_n750 ) , .B1( us32_n751 ) , .A1( us32_n752 ) , .ZN( us32_n756 ) , .A2( us32_n806 ) );
  NOR2_X1 us32_U234 (.ZN( us32_n751 ) , .A2( us32_n852 ) , .A1( us32_n860 ) );
  NOR3_X1 us32_U235 (.ZN( us32_n752 ) , .A2( us32_n853 ) , .A1( us32_n863 ) , .A3( us32_n865 ) );
  NOR2_X1 us32_U236 (.ZN( us32_n544 ) , .A2( us32_n785 ) , .A1( us32_n792 ) );
  NOR2_X1 us32_U237 (.ZN( us32_n663 ) , .A1( us32_n729 ) , .A2( us32_n785 ) );
  INV_X1 us32_U238 (.A( us32_n806 ) , .ZN( us32_n841 ) );
  NOR2_X1 us32_U239 (.ZN( us32_n506 ) , .A2( us32_n728 ) , .A1( us32_n762 ) );
  NOR4_X1 us32_U24 (.A4( us32_n544 ) , .A3( us32_n545 ) , .A2( us32_n546 ) , .A1( us32_n547 ) , .ZN( us32_n548 ) );
  NOR2_X1 us32_U240 (.ZN( us32_n631 ) , .A1( us32_n724 ) , .A2( us32_n813 ) );
  NOR2_X1 us32_U241 (.ZN( us32_n614 ) , .A1( us32_n762 ) , .A2( us32_n812 ) );
  NOR2_X1 us32_U242 (.ZN( us32_n530 ) , .A2( us32_n744 ) , .A1( us32_n792 ) );
  NOR2_X1 us32_U243 (.ZN( us32_n558 ) , .A1( us32_n708 ) , .A2( us32_n816 ) );
  NOR2_X1 us32_U244 (.ZN( us32_n516 ) , .A1( us32_n708 ) , .A2( us32_n744 ) );
  NOR2_X1 us32_U245 (.A2( us32_n697 ) , .ZN( us32_n716 ) , .A1( us32_n792 ) );
  NOR2_X1 us32_U246 (.A1( us32_n749 ) , .ZN( us32_n767 ) , .A2( us32_n803 ) );
  NOR2_X1 us32_U247 (.ZN( us32_n521 ) , .A1( us32_n790 ) , .A2( us32_n812 ) );
  NOR2_X1 us32_U248 (.ZN( us32_n655 ) , .A1( us32_n790 ) , .A2( us32_n815 ) );
  NOR2_X1 us32_U249 (.ZN( us32_n668 ) , .A2( us32_n708 ) , .A1( us32_n790 ) );
  NOR4_X1 us32_U25 (.ZN( us32_n479 ) , .A1( us32_n520 ) , .A4( us32_n557 ) , .A3( us32_n582 ) , .A2( us32_n630 ) );
  NOR2_X1 us32_U250 (.ZN( us32_n517 ) , .A1( us32_n708 ) , .A2( us32_n803 ) );
  INV_X1 us32_U251 (.A( us32_n763 ) , .ZN( us32_n866 ) );
  NOR2_X1 us32_U252 (.ZN( us32_n542 ) , .A1( us32_n762 ) , .A2( us32_n791 ) );
  NOR2_X1 us32_U253 (.ZN( us32_n630 ) , .A1( us32_n747 ) , .A2( us32_n815 ) );
  INV_X1 us32_U254 (.A( us32_n729 ) , .ZN( us32_n868 ) );
  NOR2_X1 us32_U255 (.ZN( us32_n609 ) , .A2( us32_n724 ) , .A1( us32_n817 ) );
  AOI21_X1 us32_U256 (.A( us32_n815 ) , .B2( us32_n816 ) , .B1( us32_n817 ) , .ZN( us32_n818 ) );
  NOR2_X1 us32_U257 (.ZN( us32_n579 ) , .A2( us32_n708 ) , .A1( us32_n730 ) );
  NOR2_X1 us32_U258 (.ZN( us32_n533 ) , .A2( us32_n724 ) , .A1( us32_n730 ) );
  NOR2_X1 us32_U259 (.ZN( us32_n642 ) , .A2( us32_n788 ) , .A1( us32_n791 ) );
  NOR4_X1 us32_U26 (.ZN( us32_n456 ) , .A2( us32_n517 ) , .A1( us32_n543 ) , .A3( us32_n579 ) , .A4( us32_n615 ) );
  AOI21_X1 us32_U260 (.B1( us32_n625 ) , .ZN( us32_n627 ) , .A( us32_n763 ) , .B2( us32_n814 ) );
  NOR2_X1 us32_U261 (.ZN( us32_n656 ) , .A1( us32_n747 ) , .A2( us32_n780 ) );
  AOI21_X1 us32_U262 (.A( us32_n812 ) , .B2( us32_n813 ) , .B1( us32_n814 ) , .ZN( us32_n819 ) );
  NOR2_X1 us32_U263 (.A2( us32_n697 ) , .A1( us32_n780 ) , .ZN( us32_n820 ) );
  AOI21_X1 us32_U264 (.ZN( us32_n499 ) , .B1( us32_n680 ) , .A( us32_n812 ) , .B2( us32_n816 ) );
  NOR2_X1 us32_U265 (.A2( us32_n708 ) , .A1( us32_n762 ) , .ZN( us32_n794 ) );
  AOI21_X1 us32_U266 (.ZN( us32_n593 ) , .B1( us32_n750 ) , .A( us32_n792 ) , .B2( us32_n813 ) );
  AOI21_X1 us32_U267 (.ZN( us32_n626 ) , .B2( us32_n669 ) , .A( us32_n790 ) , .B1( us32_n791 ) );
  NOR2_X1 us32_U268 (.ZN( us32_n520 ) , .A2( us32_n708 ) , .A1( us32_n814 ) );
  NOR2_X1 us32_U269 (.A1( us32_n697 ) , .ZN( us32_n770 ) , .A2( us32_n815 ) );
  NOR4_X1 us32_U27 (.A4( us32_n532 ) , .A3( us32_n533 ) , .A2( us32_n534 ) , .ZN( us32_n535 ) , .A1( us32_n820 ) );
  NOR2_X1 us32_U270 (.ZN( us32_n582 ) , .A1( us32_n744 ) , .A2( us32_n815 ) );
  NOR2_X1 us32_U271 (.ZN( us32_n519 ) , .A2( us32_n699 ) , .A1( us32_n816 ) );
  AOI21_X1 us32_U272 (.ZN( us32_n477 ) , .A( us32_n669 ) , .B1( us32_n750 ) , .B2( us32_n806 ) );
  AOI21_X1 us32_U273 (.ZN( us32_n510 ) , .B2( us32_n669 ) , .A( us32_n730 ) , .B1( us32_n815 ) );
  INV_X1 us32_U274 (.A( us32_n813 ) , .ZN( us32_n836 ) );
  AOI21_X1 us32_U275 (.ZN( us32_n589 ) , .B2( us32_n699 ) , .B1( us32_n815 ) , .A( us32_n817 ) );
  AOI21_X1 us32_U276 (.ZN( us32_n515 ) , .A( us32_n729 ) , .B1( us32_n750 ) , .B2( us32_n803 ) );
  AOI21_X1 us32_U277 (.ZN( us32_n539 ) , .B2( us32_n812 ) , .A( us32_n814 ) , .B1( us32_n815 ) );
  NOR2_X1 us32_U278 (.ZN( us32_n581 ) , .A1( us32_n669 ) , .A2( us32_n788 ) );
  NOR2_X1 us32_U279 (.ZN( us32_n547 ) , .A1( us32_n699 ) , .A2( us32_n744 ) );
  NOR4_X1 us32_U28 (.ZN( us32_n474 ) , .A1( us32_n506 ) , .A3( us32_n544 ) , .A2( us32_n583 ) , .A4( us32_n716 ) );
  AOI21_X1 us32_U280 (.ZN( us32_n540 ) , .A( us32_n763 ) , .B2( us32_n779 ) , .B1( us32_n817 ) );
  AOI21_X1 us32_U281 (.B1( us32_n699 ) , .ZN( us32_n700 ) , .A( us32_n732 ) , .B2( us32_n763 ) );
  AOI21_X1 us32_U282 (.ZN( us32_n591 ) , .B2( us32_n763 ) , .A( us32_n785 ) , .B1( us32_n812 ) );
  INV_X1 us32_U283 (.A( us32_n791 ) , .ZN( us32_n873 ) );
  NOR2_X1 us32_U284 (.ZN( us32_n559 ) , .A2( us32_n791 ) , .A1( us32_n803 ) );
  AOI21_X1 us32_U285 (.ZN( us32_n498 ) , .A( us32_n724 ) , .B2( us32_n762 ) , .B1( us32_n814 ) );
  NOR2_X1 us32_U286 (.ZN( us32_n683 ) , .A2( us32_n699 ) , .A1( us32_n803 ) );
  NOR2_X1 us32_U287 (.ZN( us32_n685 ) , .A1( us32_n729 ) , .A2( us32_n816 ) );
  AOI21_X1 us32_U288 (.B1( us32_n686 ) , .ZN( us32_n687 ) , .A( us32_n728 ) , .B2( us32_n761 ) );
  AOI21_X1 us32_U289 (.ZN( us32_n569 ) , .B1( us32_n750 ) , .B2( us32_n762 ) , .A( us32_n780 ) );
  AOI221_X1 us32_U29 (.A( us32_n713 ) , .B2( us32_n714 ) , .ZN( us32_n720 ) , .C1( us32_n832 ) , .B1( us32_n839 ) , .C2( us32_n863 ) );
  AOI21_X1 us32_U290 (.ZN( us32_n649 ) , .B1( us32_n729 ) , .B2( us32_n763 ) , .A( us32_n813 ) );
  NOR2_X1 us32_U291 (.ZN( us32_n568 ) , .A1( us32_n729 ) , .A2( us32_n762 ) );
  INV_X1 us32_U292 (.A( us32_n699 ) , .ZN( us32_n853 ) );
  NOR2_X1 us32_U293 (.ZN( us32_n566 ) , .A2( us32_n697 ) , .A1( us32_n763 ) );
  AOI21_X1 us32_U294 (.ZN( us32_n514 ) , .A( us32_n779 ) , .B2( us32_n792 ) , .B1( us32_n812 ) );
  AOI21_X1 us32_U295 (.ZN( us32_n639 ) , .B2( us32_n749 ) , .A( us32_n788 ) , .B1( us32_n812 ) );
  NOR2_X1 us32_U296 (.ZN( us32_n665 ) , .A1( us32_n780 ) , .A2( us32_n813 ) );
  AOI21_X1 us32_U297 (.ZN( us32_n571 ) , .B2( us32_n697 ) , .B1( us32_n806 ) , .A( us32_n812 ) );
  AOI21_X1 us32_U298 (.ZN( us32_n564 ) , .B1( us32_n724 ) , .A( us32_n779 ) , .B2( us32_n791 ) );
  AOI21_X1 us32_U299 (.ZN( us32_n497 ) , .A( us32_n779 ) , .B2( us32_n791 ) , .B1( us32_n804 ) );
  NAND2_X1 us32_U3 (.A1( us32_n449 ) , .A2( us32_n464 ) , .ZN( us32_n724 ) );
  OR2_X1 us32_U30 (.A2( us32_n711 ) , .A1( us32_n712 ) , .ZN( us32_n713 ) );
  AOI21_X1 us32_U300 (.ZN( us32_n640 ) , .B2( us32_n747 ) , .A( us32_n792 ) , .B1( us32_n803 ) );
  NOR2_X1 us32_U301 (.ZN( us32_n578 ) , .A1( us32_n708 ) , .A2( us32_n813 ) );
  NOR2_X1 us32_U302 (.ZN( us32_n529 ) , .A1( us32_n708 ) , .A2( us32_n779 ) );
  AOI21_X1 us32_U303 (.ZN( us32_n689 ) , .B2( us32_n749 ) , .B1( us32_n763 ) , .A( us32_n806 ) );
  AOI21_X1 us32_U304 (.A( us32_n790 ) , .B2( us32_n791 ) , .B1( us32_n792 ) , .ZN( us32_n793 ) );
  AOI21_X1 us32_U305 (.ZN( us32_n478 ) , .B2( us32_n697 ) , .A( us32_n749 ) , .B1( us32_n779 ) );
  NOR2_X1 us32_U306 (.ZN( us32_n684 ) , .A1( us32_n791 ) , .A2( us32_n813 ) );
  AOI21_X1 us32_U307 (.ZN( us32_n450 ) , .B2( us32_n792 ) , .A( us32_n803 ) , .B1( us32_n815 ) );
  AOI21_X1 us32_U308 (.A( us32_n733 ) , .ZN( us32_n734 ) , .B2( us32_n780 ) , .B1( us32_n792 ) );
  NOR2_X1 us32_U309 (.A2( us32_n813 ) , .A1( us32_n815 ) , .ZN( us32_n821 ) );
  NOR2_X1 us32_U31 (.ZN( us32_n680 ) , .A2( us32_n834 ) , .A1( us32_n839 ) );
  AOI21_X1 us32_U310 (.ZN( us32_n641 ) , .B1( us32_n680 ) , .A( us32_n791 ) , .B2( us32_n817 ) );
  NOR2_X1 us32_U311 (.ZN( us32_n583 ) , .A1( us32_n792 ) , .A2( us32_n817 ) );
  NOR2_X1 us32_U312 (.ZN( us32_n711 ) , .A1( us32_n762 ) , .A2( us32_n763 ) );
  NOR2_X1 us32_U313 (.ZN( us32_n534 ) , .A1( us32_n724 ) , .A2( us32_n788 ) );
  NOR2_X1 us32_U314 (.ZN( us32_n632 ) , .A2( us32_n697 ) , .A1( us32_n724 ) );
  NOR2_X1 us32_U315 (.ZN( us32_n580 ) , .A2( us32_n697 ) , .A1( us32_n791 ) );
  NOR2_X1 us32_U316 (.ZN( us32_n682 ) , .A2( us32_n708 ) , .A1( us32_n817 ) );
  INV_X1 us32_U317 (.A( us32_n815 ) , .ZN( us32_n855 ) );
  AOI21_X1 us32_U318 (.ZN( us32_n442 ) , .A( us32_n699 ) , .B1( us32_n733 ) , .B2( us32_n750 ) );
  INV_X1 us32_U319 (.A( us32_n780 ) , .ZN( us32_n850 ) );
  NOR4_X1 us32_U32 (.A4( us32_n514 ) , .A3( us32_n515 ) , .A2( us32_n516 ) , .A1( us32_n517 ) , .ZN( us32_n524 ) );
  INV_X1 us32_U320 (.A( us32_n785 ) , .ZN( us32_n846 ) );
  NAND2_X1 us32_U321 (.ZN( us32_n714 ) , .A1( us32_n728 ) , .A2( us32_n780 ) );
  NAND2_X1 us32_U322 (.ZN( us32_n671 ) , .A1( us32_n806 ) , .A2( us32_n816 ) );
  AOI21_X1 us32_U323 (.ZN( us32_n443 ) , .B1( us32_n789 ) , .B2( us32_n791 ) , .A( us32_n814 ) );
  NOR2_X1 us32_U324 (.ZN( us32_n470 ) , .A2( us32_n779 ) , .A1( us32_n815 ) );
  NAND2_X1 us32_U325 (.A2( us32_n762 ) , .A1( us32_n806 ) , .ZN( us32_n810 ) );
  NOR2_X1 us32_U326 (.ZN( us32_n526 ) , .A1( us32_n724 ) , .A2( us32_n750 ) );
  OAI21_X1 us32_U327 (.A( us32_n787 ) , .B2( us32_n788 ) , .B1( us32_n789 ) , .ZN( us32_n795 ) );
  OAI21_X1 us32_U328 (.ZN( us32_n787 ) , .A( us32_n839 ) , .B1( us32_n863 ) , .B2( us32_n873 ) );
  NAND2_X1 us32_U329 (.A1( us32_n699 ) , .A2( us32_n729 ) , .ZN( us32_n782 ) );
  AOI222_X1 us32_U33 (.ZN( us32_n525 ) , .A1( us32_n834 ) , .B2( us32_n837 ) , .C1( us32_n844 ) , .C2( us32_n850 ) , .A2( us32_n852 ) , .B1( us32_n866 ) );
  NOR2_X1 us32_U330 (.ZN( us32_n712 ) , .A2( us32_n724 ) , .A1( us32_n790 ) );
  NOR2_X1 us32_U331 (.ZN( us32_n518 ) , .A1( us32_n708 ) , .A2( us32_n788 ) );
  OAI21_X1 us32_U332 (.A( us32_n698 ) , .ZN( us32_n702 ) , .B2( us32_n750 ) , .B1( us32_n804 ) );
  OAI21_X1 us32_U333 (.ZN( us32_n698 ) , .B2( us32_n833 ) , .B1( us32_n838 ) , .A( us32_n860 ) );
  INV_X1 us32_U334 (.A( us32_n817 ) , .ZN( us32_n844 ) );
  INV_X1 us32_U335 (.A( us32_n724 ) , .ZN( us32_n856 ) );
  OAI21_X1 us32_U336 (.ZN( us32_n731 ) , .A( us32_n833 ) , .B2( us32_n852 ) , .B1( us32_n873 ) );
  AND2_X1 us32_U337 (.ZN( us32_n732 ) , .A1( us32_n779 ) , .A2( us32_n785 ) );
  AOI221_X1 us32_U338 (.A( us32_n764 ) , .ZN( us32_n774 ) , .C2( us32_n810 ) , .B2( us32_n835 ) , .C1( us32_n855 ) , .B1( us32_n866 ) );
  AOI21_X1 us32_U339 (.B2( us32_n763 ) , .ZN( us32_n764 ) , .A( us32_n788 ) , .B1( us32_n792 ) );
  NOR4_X1 us32_U34 (.A3( us32_n521 ) , .A1( us32_n522 ) , .ZN( us32_n523 ) , .A2( us32_n673 ) , .A4( us32_n769 ) );
  INV_X1 us32_U340 (.A( us32_n761 ) , .ZN( us32_n835 ) );
  NAND2_X1 us32_U341 (.A2( us32_n448 ) , .A1( us32_n460 ) , .ZN( us32_n728 ) );
  NAND2_X1 us32_U342 (.A1( us32_n451 ) , .A2( us32_n454 ) , .ZN( us32_n814 ) );
  NAND2_X1 us32_U343 (.A1( us32_n455 ) , .A2( us32_n462 ) , .ZN( us32_n750 ) );
  NAND2_X1 us32_U344 (.A1( us32_n451 ) , .A2( us32_n471 ) , .ZN( us32_n816 ) );
  NAND2_X1 us32_U345 (.A1( us32_n454 ) , .A2( us32_n461 ) , .ZN( us32_n813 ) );
  NAND2_X1 us32_U346 (.A1( us32_n452 ) , .A2( us32_n465 ) , .ZN( us32_n669 ) );
  NAND2_X1 us32_U347 (.A1( us32_n453 ) , .A2( us32_n472 ) , .ZN( us32_n785 ) );
  NAND2_X1 us32_U348 (.A1( us32_n453 ) , .A2( us32_n461 ) , .ZN( us32_n744 ) );
  NAND2_X1 us32_U349 (.A2( us32_n453 ) , .A1( us32_n455 ) , .ZN( us32_n806 ) );
  AOI221_X1 us32_U35 (.A( us32_n781 ) , .ZN( us32_n798 ) , .C2( us32_n837 ) , .B2( us32_n838 ) , .B1( us32_n865 ) , .C1( us32_n866 ) );
  NAND2_X1 us32_U350 (.A1( us32_n455 ) , .A2( us32_n471 ) , .ZN( us32_n803 ) );
  NAND2_X1 us32_U351 (.A2( us32_n454 ) , .A1( us32_n472 ) , .ZN( us32_n779 ) );
  NAND2_X1 us32_U352 (.A2( us32_n464 ) , .A1( us32_n465 ) , .ZN( us32_n812 ) );
  NAND2_X1 us32_U353 (.A1( us32_n441 ) , .A2( us32_n460 ) , .ZN( us32_n699 ) );
  NAND2_X1 us32_U354 (.A2( us32_n448 ) , .A1( us32_n452 ) , .ZN( us32_n729 ) );
  NAND2_X1 us32_U355 (.A2( us32_n449 ) , .A1( us32_n452 ) , .ZN( us32_n763 ) );
  NOR2_X1 us32_U356 (.ZN( us32_n465 ) , .A2( us32_n847 ) , .A1( us32_n848 ) );
  NOR2_X1 us32_U357 (.ZN( us32_n453 ) , .A1( us32_n826 ) , .A2( us32_n827 ) );
  NAND2_X1 us32_U358 (.A1( us32_n462 ) , .A2( us32_n472 ) , .ZN( us32_n788 ) );
  NOR2_X1 us32_U359 (.ZN( us32_n451 ) , .A1( us32_n828 ) , .A2( us32_n829 ) );
  NOR4_X1 us32_U36 (.A4( us32_n793 ) , .A3( us32_n794 ) , .A2( us32_n795 ) , .A1( us32_n796 ) , .ZN( us32_n797 ) );
  NAND2_X1 us32_U360 (.A2( us32_n461 ) , .A1( us32_n462 ) , .ZN( us32_n747 ) );
  NAND2_X1 us32_U361 (.A1( us32_n451 ) , .A2( us32_n462 ) , .ZN( us32_n790 ) );
  NAND2_X2 us32_U362 (.A2( us32_n448 ) , .A1( us32_n464 ) , .ZN( us32_n815 ) );
  NAND2_X1 us32_U363 (.A2( us32_n441 ) , .A1( us32_n447 ) , .ZN( us32_n784 ) );
  NAND2_X1 us32_U364 (.A1( us32_n447 ) , .A2( us32_n449 ) , .ZN( us32_n805 ) );
  NAND2_X1 us32_U365 (.A2( us32_n454 ) , .A1( us32_n455 ) , .ZN( us32_n730 ) );
  NAND2_X2 us32_U366 (.A1( us32_n449 ) , .A2( us32_n460 ) , .ZN( us32_n792 ) );
  NAND2_X2 us32_U367 (.A2( us32_n460 ) , .A1( us32_n465 ) , .ZN( us32_n780 ) );
  NOR2_X1 us32_U368 (.ZN( us32_n447 ) , .A2( us32_n849 ) , .A1( us32_n858 ) );
  NAND2_X1 us32_U369 (.A1( us32_n447 ) , .A2( us32_n448 ) , .ZN( us32_n786 ) );
  NOR4_X1 us32_U37 (.A4( us32_n776 ) , .A3( us32_n777 ) , .A1( us32_n778 ) , .ZN( us32_n799 ) , .A2( us32_n801 ) );
  NAND2_X1 us32_U370 (.A2( us32_n471 ) , .A1( us32_n472 ) , .ZN( us32_n817 ) );
  NOR2_X1 us32_U371 (.A2( sa32_6 ) , .A1( sa32_7 ) , .ZN( us32_n464 ) );
  NOR2_X1 us32_U372 (.A2( sa32_7 ) , .ZN( us32_n460 ) , .A1( us32_n849 ) );
  NOR2_X1 us32_U373 (.A2( sa32_4 ) , .ZN( us32_n449 ) , .A1( us32_n848 ) );
  NOR2_X1 us32_U374 (.A2( sa32_4 ) , .A1( sa32_5 ) , .ZN( us32_n441 ) );
  NOR2_X1 us32_U375 (.A2( sa32_5 ) , .ZN( us32_n448 ) , .A1( us32_n847 ) );
  NOR2_X1 us32_U376 (.A2( sa32_2 ) , .A1( sa32_3 ) , .ZN( us32_n472 ) );
  NOR2_X1 us32_U377 (.A2( sa32_6 ) , .ZN( us32_n452 ) , .A1( us32_n858 ) );
  NOR2_X1 us32_U378 (.A2( sa32_1 ) , .ZN( us32_n471 ) , .A1( us32_n826 ) );
  NOR2_X1 us32_U379 (.A2( sa32_0 ) , .ZN( us32_n454 ) , .A1( us32_n827 ) );
  NOR4_X1 us32_U38 (.A3( us32_n755 ) , .A2( us32_n756 ) , .A1( us32_n757 ) , .ZN( us32_n758 ) , .A4( us32_n869 ) );
  NOR2_X1 us32_U380 (.A2( sa32_0 ) , .A1( sa32_1 ) , .ZN( us32_n462 ) );
  NOR2_X1 us32_U381 (.A2( sa32_3 ) , .ZN( us32_n455 ) , .A1( us32_n828 ) );
  NOR2_X1 us32_U382 (.A2( sa32_2 ) , .ZN( us32_n461 ) , .A1( us32_n829 ) );
  INV_X1 us32_U383 (.A( sa32_4 ) , .ZN( us32_n847 ) );
  INV_X1 us32_U384 (.A( sa32_6 ) , .ZN( us32_n849 ) );
  INV_X1 us32_U385 (.A( sa32_3 ) , .ZN( us32_n829 ) );
  INV_X1 us32_U386 (.A( sa32_1 ) , .ZN( us32_n827 ) );
  INV_X1 us32_U387 (.A( sa32_0 ) , .ZN( us32_n826 ) );
  INV_X1 us32_U388 (.A( sa32_2 ) , .ZN( us32_n828 ) );
  INV_X1 us32_U389 (.A( sa32_5 ) , .ZN( us32_n848 ) );
  AOI211_X1 us32_U39 (.B( us32_n745 ) , .A( us32_n746 ) , .ZN( us32_n759 ) , .C1( us32_n832 ) , .C2( us32_n853 ) );
  INV_X1 us32_U390 (.A( sa32_7 ) , .ZN( us32_n858 ) );
  NAND2_X1 us32_U391 (.A2( us32_n461 ) , .A1( us32_n471 ) , .ZN( us32_n697 ) );
  OAI222_X1 us32_U392 (.B2( us32_n747 ) , .B1( us32_n748 ) , .A2( us32_n749 ) , .ZN( us32_n757 ) , .C2( us32_n805 ) , .C1( us32_n814 ) , .A1( us32_n817 ) );
  OAI22_X1 us32_U393 (.B2( us32_n803 ) , .B1( us32_n804 ) , .A2( us32_n805 ) , .A1( us32_n806 ) , .ZN( us32_n808 ) );
  OAI21_X1 us32_U394 (.A( us32_n731 ) , .B1( us32_n732 ) , .ZN( us32_n736 ) , .B2( us32_n805 ) );
  OAI222_X1 us32_U395 (.ZN( us32_n505 ) , .C2( us32_n625 ) , .B2( us32_n647 ) , .B1( us32_n747 ) , .A2( us32_n748 ) , .C1( us32_n805 ) , .A1( us32_n806 ) );
  AOI21_X1 us32_U396 (.ZN( us32_n650 ) , .A( us32_n779 ) , .B1( us32_n792 ) , .B2( us32_n805 ) );
  INV_X1 us32_U397 (.A( us32_n805 ) , .ZN( us32_n860 ) );
  NOR2_X1 us32_U398 (.ZN( us32_n735 ) , .A2( us32_n803 ) , .A1( us32_n805 ) );
  NOR2_X1 us32_U399 (.ZN( us32_n484 ) , .A1( us32_n788 ) , .A2( us32_n805 ) );
  NAND2_X1 us32_U4 (.A1( us32_n441 ) , .A2( us32_n464 ) , .ZN( us32_n708 ) );
  NOR3_X1 us32_U40 (.A3( us32_n741 ) , .A2( us32_n742 ) , .A1( us32_n743 ) , .ZN( us32_n760 ) );
  NOR2_X1 us32_U400 (.A2( us32_n744 ) , .ZN( us32_n755 ) , .A1( us32_n805 ) );
  NAND2_X1 us32_U401 (.ZN( us32_n753 ) , .A1( us32_n763 ) , .A2( us32_n805 ) );
  NOR2_X1 us32_U402 (.ZN( us32_n715 ) , .A1( us32_n805 ) , .A2( us32_n817 ) );
  NOR2_X1 us32_U403 (.ZN( us32_n567 ) , .A1( us32_n747 ) , .A2( us32_n805 ) );
  AOI21_X1 us32_U404 (.ZN( us32_n552 ) , .B1( us32_n669 ) , .A( us32_n697 ) , .B2( us32_n805 ) );
  NOR2_X1 us32_U405 (.ZN( us32_n556 ) , .A1( us32_n762 ) , .A2( us32_n805 ) );
  NOR2_X1 us32_U406 (.ZN( us32_n670 ) , .A1( us32_n790 ) , .A2( us32_n805 ) );
  OAI221_X1 us32_U407 (.A( us32_n783 ) , .C2( us32_n784 ) , .B2( us32_n785 ) , .B1( us32_n786 ) , .ZN( us32_n796 ) , .C1( us32_n813 ) );
  NAND2_X1 us32_U408 (.A1( us32_n729 ) , .A2( us32_n784 ) , .ZN( us32_n811 ) );
  OAI22_X1 us32_U409 (.ZN( us32_n588 ) , .A2( us32_n747 ) , .B2( us32_n762 ) , .A1( us32_n763 ) , .B1( us32_n784 ) );
  NAND4_X1 us32_U41 (.ZN( sa33_sr_3 ) , .A4( us32_n704 ) , .A3( us32_n705 ) , .A2( us32_n706 ) , .A1( us32_n707 ) );
  AOI21_X1 us32_U410 (.ZN( us32_n592 ) , .B1( us32_n728 ) , .B2( us32_n784 ) , .A( us32_n790 ) );
  AOI21_X1 us32_U411 (.ZN( us32_n623 ) , .B1( us32_n699 ) , .A( us32_n779 ) , .B2( us32_n784 ) );
  AOI21_X1 us32_U412 (.ZN( us32_n648 ) , .A( us32_n762 ) , .B2( us32_n784 ) , .B1( us32_n792 ) );
  OAI22_X1 us32_U413 (.ZN( us32_n681 ) , .A1( us32_n699 ) , .A2( us32_n730 ) , .B2( us32_n784 ) , .B1( us32_n817 ) );
  OAI21_X1 us32_U414 (.A( us32_n613 ) , .ZN( us32_n616 ) , .B1( us32_n625 ) , .B2( us32_n784 ) );
  NOR2_X1 us32_U415 (.ZN( us32_n610 ) , .A1( us32_n784 ) , .A2( us32_n816 ) );
  OAI222_X1 us32_U416 (.A2( us32_n669 ) , .ZN( us32_n674 ) , .B1( us32_n747 ) , .B2( us32_n784 ) , .C2( us32_n788 ) , .C1( us32_n815 ) , .A1( us32_n817 ) );
  NOR2_X1 us32_U417 (.ZN( us32_n651 ) , .A1( us32_n784 ) , .A2( us32_n788 ) );
  NOR2_X1 us32_U418 (.ZN( us32_n600 ) , .A2( us32_n697 ) , .A1( us32_n784 ) );
  NOR2_X1 us32_U419 (.ZN( us32_n553 ) , .A2( us32_n744 ) , .A1( us32_n784 ) );
  NOR4_X1 us32_U42 (.A4( us32_n700 ) , .A3( us32_n701 ) , .A2( us32_n702 ) , .A1( us32_n703 ) , .ZN( us32_n704 ) );
  INV_X1 us32_U420 (.A( us32_n784 ) , .ZN( us32_n861 ) );
  AOI21_X1 us32_U421 (.ZN( us32_n500 ) , .A( us32_n697 ) , .B1( us32_n708 ) , .B2( us32_n786 ) );
  OAI221_X1 us32_U422 (.A( us32_n696 ) , .ZN( us32_n703 ) , .C2( us32_n784 ) , .C1( us32_n785 ) , .B1( us32_n786 ) , .B2( us32_n806 ) );
  OAI22_X1 us32_U423 (.ZN( us32_n590 ) , .B1( us32_n730 ) , .B2( us32_n749 ) , .A2( us32_n786 ) , .A1( us32_n803 ) );
  NOR2_X1 us32_U424 (.ZN( us32_n612 ) , .A1( us32_n779 ) , .A2( us32_n786 ) );
  NAND2_X1 us32_U425 (.A2( us32_n749 ) , .A1( us32_n786 ) , .ZN( us32_n809 ) );
  OAI222_X1 us32_U426 (.ZN( us32_n617 ) , .B1( us32_n697 ) , .C1( us32_n724 ) , .C2( us32_n747 ) , .B2( us32_n786 ) , .A2( us32_n792 ) , .A1( us32_n816 ) );
  NOR2_X1 us32_U427 (.ZN( us32_n717 ) , .A2( us32_n744 ) , .A1( us32_n786 ) );
  NOR2_X1 us32_U428 (.ZN( us32_n653 ) , .A1( us32_n762 ) , .A2( us32_n786 ) );
  NOR2_X1 us32_U429 (.ZN( us32_n554 ) , .A1( us32_n786 ) , .A2( us32_n813 ) );
  AOI211_X1 us32_U43 (.B( us32_n694 ) , .A( us32_n695 ) , .ZN( us32_n705 ) , .C2( us32_n831 ) , .C1( us32_n851 ) );
  NOR2_X1 us32_U430 (.ZN( us32_n701 ) , .A2( us32_n786 ) , .A1( us32_n817 ) );
  NOR2_X1 us32_U431 (.A1( us32_n730 ) , .ZN( us32_n765 ) , .A2( us32_n786 ) );
  AND2_X1 us32_U432 (.ZN( us32_n438 ) , .A2( us32_n831 ) , .A1( us32_n854 ) );
  AND2_X1 us32_U433 (.ZN( us32_n439 ) , .A2( us32_n843 ) , .A1( us32_n861 ) );
  NOR3_X1 us32_U434 (.A1( us32_n438 ) , .A2( us32_n439 ) , .A3( us32_n576 ) , .ZN( us32_n587 ) );
  NAND4_X1 us32_U435 (.ZN( sa33_sr_2 ) , .A4( us32_n643 ) , .A3( us32_n644 ) , .A2( us32_n645 ) , .A1( us32_n646 ) );
  INV_X1 us32_U436 (.A( us32_n812 ) , .ZN( us32_n854 ) );
  NAND3_X1 us32_U437 (.ZN( sa33_sr_6 ) , .A3( us32_n797 ) , .A2( us32_n798 ) , .A1( us32_n799 ) );
  NAND3_X1 us32_U438 (.ZN( sa33_sr_5 ) , .A3( us32_n758 ) , .A2( us32_n759 ) , .A1( us32_n760 ) );
  NAND3_X1 us32_U439 (.ZN( sa33_sr_4 ) , .A3( us32_n738 ) , .A2( us32_n739 ) , .A1( us32_n740 ) );
  NOR2_X1 us32_U44 (.ZN( us32_n707 ) , .A2( us32_n776 ) , .A1( us32_n800 ) );
  NAND3_X1 us32_U440 (.A3( us32_n675 ) , .A2( us32_n676 ) , .A1( us32_n677 ) , .ZN( us32_n807 ) );
  NAND3_X1 us32_U441 (.ZN( us32_n638 ) , .A3( us32_n708 ) , .A2( us32_n724 ) , .A1( us32_n792 ) );
  NAND3_X1 us32_U442 (.A3( us32_n618 ) , .A2( us32_n619 ) , .A1( us32_n620 ) , .ZN( us32_n725 ) );
  NAND3_X1 us32_U443 (.A3( us32_n585 ) , .A2( us32_n586 ) , .A1( us32_n587 ) , .ZN( us32_n621 ) );
  NAND3_X1 us32_U444 (.ZN( us32_n565 ) , .A3( us32_n680 ) , .A2( us32_n750 ) , .A1( us32_n785 ) );
  NAND3_X1 us32_U445 (.A3( us32_n523 ) , .A2( us32_n524 ) , .A1( us32_n525 ) , .ZN( us32_n742 ) );
  NAND3_X1 us32_U446 (.A3( us32_n512 ) , .A1( us32_n513 ) , .ZN( us32_n608 ) , .A2( us32_n871 ) );
  NAND3_X1 us32_U447 (.A3( us32_n467 ) , .A2( us32_n468 ) , .A1( us32_n469 ) , .ZN( us32_n777 ) );
  INV_X1 us32_U448 (.A( us32_n803 ) , .ZN( us32_n843 ) );
  AOI21_X1 us32_U449 (.ZN( us32_n576 ) , .B2( us32_n724 ) , .B1( us32_n748 ) , .A( us32_n785 ) );
  AOI222_X1 us32_U45 (.B2( us32_n638 ) , .ZN( us32_n644 ) , .B1( us32_n841 ) , .A1( us32_n842 ) , .C2( us32_n846 ) , .C1( us32_n863 ) , .A2( us32_n865 ) );
  NOR4_X1 us32_U46 (.A4( us32_n639 ) , .A3( us32_n640 ) , .A2( us32_n641 ) , .A1( us32_n642 ) , .ZN( us32_n643 ) );
  NOR3_X1 us32_U47 (.A2( us32_n607 ) , .A1( us32_n608 ) , .ZN( us32_n646 ) , .A3( us32_n722 ) );
  NAND4_X1 us32_U48 (.ZN( sa33_sr_7 ) , .A4( us32_n822 ) , .A3( us32_n823 ) , .A2( us32_n824 ) , .A1( us32_n825 ) );
  NOR4_X1 us32_U49 (.A4( us32_n818 ) , .A3( us32_n819 ) , .A2( us32_n820 ) , .A1( us32_n821 ) , .ZN( us32_n822 ) );
  NAND2_X1 us32_U5 (.A2( us32_n441 ) , .A1( us32_n452 ) , .ZN( us32_n791 ) );
  AOI222_X1 us32_U50 (.C2( us32_n809 ) , .B2( us32_n810 ) , .A2( us32_n811 ) , .ZN( us32_n823 ) , .C1( us32_n832 ) , .A1( us32_n839 ) , .B1( us32_n853 ) );
  AOI211_X1 us32_U51 (.B( us32_n807 ) , .A( us32_n808 ) , .ZN( us32_n824 ) , .C1( us32_n842 ) , .C2( us32_n850 ) );
  NAND4_X1 us32_U52 (.ZN( sa33_sr_0 ) , .A4( us32_n501 ) , .A3( us32_n502 ) , .A2( us32_n503 ) , .A1( us32_n504 ) );
  AOI221_X1 us32_U53 (.A( us32_n497 ) , .ZN( us32_n502 ) , .B2( us32_n843 ) , .C1( us32_n846 ) , .C2( us32_n860 ) , .B1( us32_n862 ) );
  NOR4_X1 us32_U54 (.A4( us32_n498 ) , .A3( us32_n499 ) , .A2( us32_n500 ) , .ZN( us32_n501 ) , .A1( us32_n527 ) );
  AOI211_X1 us32_U55 (.A( us32_n496 ) , .ZN( us32_n503 ) , .B( us32_n802 ) , .C2( us32_n839 ) , .C1( us32_n851 ) );
  NAND4_X1 us32_U56 (.ZN( sa33_sr_1 ) , .A4( us32_n595 ) , .A3( us32_n596 ) , .A2( us32_n597 ) , .A1( us32_n598 ) );
  NOR4_X1 us32_U57 (.A4( us32_n591 ) , .A3( us32_n592 ) , .A2( us32_n593 ) , .A1( us32_n594 ) , .ZN( us32_n595 ) );
  AOI211_X1 us32_U58 (.B( us32_n589 ) , .A( us32_n590 ) , .ZN( us32_n596 ) , .C2( us32_n811 ) , .C1( us32_n833 ) );
  AOI211_X1 us32_U59 (.A( us32_n588 ) , .ZN( us32_n597 ) , .B( us32_n621 ) , .C1( us32_n845 ) , .C2( us32_n855 ) );
  NOR3_X1 us32_U6 (.ZN( us32_n598 ) , .A1( us32_n608 ) , .A3( us32_n723 ) , .A2( us32_n742 ) );
  NOR2_X1 us32_U60 (.ZN( us32_n804 ) , .A1( us32_n854 ) , .A2( us32_n861 ) );
  AOI222_X1 us32_U61 (.ZN( us32_n469 ) , .B1( us32_n832 ) , .A1( us32_n839 ) , .C1( us32_n842 ) , .C2( us32_n851 ) , .A2( us32_n855 ) , .B2( us32_n865 ) );
  NOR4_X1 us32_U62 (.A1( us32_n466 ) , .ZN( us32_n467 ) , .A4( us32_n542 ) , .A2( us32_n554 ) , .A3( us32_n614 ) );
  AOI221_X1 us32_U63 (.ZN( us32_n468 ) , .C2( us32_n714 ) , .B2( us32_n831 ) , .C1( us32_n845 ) , .B1( us32_n860 ) , .A( us32_n864 ) );
  NAND4_X1 us32_U64 (.A4( us32_n603 ) , .A3( us32_n604 ) , .A2( us32_n605 ) , .A1( us32_n606 ) , .ZN( us32_n722 ) );
  NOR3_X1 us32_U65 (.A1( us32_n599 ) , .ZN( us32_n604 ) , .A3( us32_n663 ) , .A2( us32_n770 ) );
  NOR4_X1 us32_U66 (.A3( us32_n600 ) , .A2( us32_n601 ) , .A1( us32_n602 ) , .ZN( us32_n603 ) , .A4( us32_n655 ) );
  AOI222_X1 us32_U67 (.ZN( us32_n606 ) , .A1( us32_n830 ) , .C2( us32_n837 ) , .B1( us32_n842 ) , .A2( us32_n856 ) , .B2( us32_n861 ) , .C1( us32_n868 ) );
  NAND4_X1 us32_U68 (.A4( us32_n657 ) , .A3( us32_n658 ) , .A2( us32_n659 ) , .A1( us32_n660 ) , .ZN( us32_n800 ) );
  NOR3_X1 us32_U69 (.A3( us32_n648 ) , .A2( us32_n649 ) , .A1( us32_n650 ) , .ZN( us32_n659 ) );
  NOR3_X1 us32_U7 (.A3( us32_n800 ) , .A2( us32_n801 ) , .A1( us32_n802 ) , .ZN( us32_n825 ) );
  NOR3_X1 us32_U70 (.A3( us32_n651 ) , .A2( us32_n652 ) , .A1( us32_n653 ) , .ZN( us32_n658 ) );
  NOR3_X1 us32_U71 (.A3( us32_n654 ) , .A2( us32_n655 ) , .A1( us32_n656 ) , .ZN( us32_n657 ) );
  NAND4_X1 us32_U72 (.A4( us32_n560 ) , .A3( us32_n561 ) , .A2( us32_n562 ) , .A1( us32_n563 ) , .ZN( us32_n607 ) );
  NOR4_X1 us32_U73 (.A4( us32_n556 ) , .A3( us32_n557 ) , .A2( us32_n558 ) , .A1( us32_n559 ) , .ZN( us32_n560 ) );
  NOR4_X1 us32_U74 (.ZN( us32_n561 ) , .A1( us32_n653 ) , .A3( us32_n661 ) , .A4( us32_n685 ) , .A2( us32_n768 ) );
  NOR4_X1 us32_U75 (.A4( us32_n552 ) , .A3( us32_n553 ) , .A2( us32_n554 ) , .A1( us32_n555 ) , .ZN( us32_n562 ) );
  NAND4_X1 us32_U76 (.A4( us32_n772 ) , .A3( us32_n773 ) , .A2( us32_n774 ) , .A1( us32_n775 ) , .ZN( us32_n801 ) );
  NOR3_X1 us32_U77 (.A3( us32_n765 ) , .A2( us32_n766 ) , .A1( us32_n767 ) , .ZN( us32_n773 ) );
  NOR4_X1 us32_U78 (.A4( us32_n768 ) , .A3( us32_n769 ) , .A2( us32_n770 ) , .A1( us32_n771 ) , .ZN( us32_n772 ) );
  AOI222_X1 us32_U79 (.ZN( us32_n775 ) , .A1( us32_n830 ) , .C1( us32_n834 ) , .B2( us32_n841 ) , .A2( us32_n850 ) , .B1( us32_n861 ) , .C2( us32_n873 ) );
  NOR3_X1 us32_U8 (.A3( us32_n621 ) , .A2( us32_n622 ) , .ZN( us32_n636 ) , .A1( us32_n725 ) );
  NOR4_X1 us32_U80 (.A4( us32_n665 ) , .A3( us32_n666 ) , .A2( us32_n667 ) , .A1( us32_n668 ) , .ZN( us32_n676 ) );
  NOR4_X1 us32_U81 (.A4( us32_n661 ) , .A3( us32_n662 ) , .A2( us32_n663 ) , .A1( us32_n664 ) , .ZN( us32_n677 ) );
  NOR4_X1 us32_U82 (.A3( us32_n673 ) , .A1( us32_n674 ) , .ZN( us32_n675 ) , .A4( us32_n715 ) , .A2( us32_n859 ) );
  NOR2_X1 us32_U83 (.ZN( us32_n625 ) , .A2( us32_n836 ) , .A1( us32_n839 ) );
  NOR2_X1 us32_U84 (.ZN( us32_n761 ) , .A1( us32_n833 ) , .A2( us32_n834 ) );
  NOR4_X1 us32_U85 (.A4( us32_n577 ) , .A3( us32_n578 ) , .A2( us32_n579 ) , .ZN( us32_n586 ) , .A1( us32_n683 ) );
  NOR4_X1 us32_U86 (.A1( us32_n584 ) , .ZN( us32_n585 ) , .A3( us32_n652 ) , .A2( us32_n662 ) , .A4( us32_n767 ) );
  AOI222_X1 us32_U87 (.ZN( us32_n513 ) , .C1( us32_n832 ) , .B2( us32_n837 ) , .A2( us32_n843 ) , .C2( us32_n862 ) , .B1( us32_n863 ) , .A1( us32_n866 ) );
  NOR4_X1 us32_U88 (.A4( us32_n509 ) , .A2( us32_n510 ) , .A1( us32_n511 ) , .ZN( us32_n512 ) , .A3( us32_n670 ) );
  INV_X1 us32_U89 (.A( us32_n505 ) , .ZN( us32_n871 ) );
  NOR2_X1 us32_U9 (.ZN( us32_n495 ) , .A1( us32_n678 ) , .A2( us32_n694 ) );
  NAND4_X1 us32_U90 (.A4( us32_n456 ) , .A3( us32_n457 ) , .A2( us32_n458 ) , .A1( us32_n459 ) , .ZN( us32_n679 ) );
  NOR3_X1 us32_U91 (.ZN( us32_n457 ) , .A3( us32_n530 ) , .A1( us32_n555 ) , .A2( us32_n570 ) );
  AOI221_X1 us32_U92 (.A( us32_n450 ) , .ZN( us32_n459 ) , .C2( us32_n753 ) , .B1( us32_n832 ) , .C1( us32_n842 ) , .B2( us32_n861 ) );
  NOR4_X1 us32_U93 (.ZN( us32_n458 ) , .A2( us32_n509 ) , .A1( us32_n599 ) , .A4( us32_n628 ) , .A3( us32_n711 ) );
  NAND4_X1 us32_U94 (.A4( us32_n535 ) , .A3( us32_n536 ) , .A2( us32_n537 ) , .A1( us32_n538 ) , .ZN( us32_n622 ) );
  NOR4_X1 us32_U95 (.A4( us32_n526 ) , .A2( us32_n527 ) , .A1( us32_n528 ) , .ZN( us32_n538 ) , .A3( us32_n701 ) );
  NOR4_X1 us32_U96 (.A1( us32_n531 ) , .ZN( us32_n536 ) , .A2( us32_n654 ) , .A4( us32_n668 ) , .A3( us32_n765 ) );
  NOR4_X1 us32_U97 (.A4( us32_n529 ) , .A3( us32_n530 ) , .ZN( us32_n537 ) , .A2( us32_n684 ) , .A1( us32_n794 ) );
  NAND4_X1 us32_U98 (.A4( us32_n479 ) , .A3( us32_n480 ) , .A2( us32_n481 ) , .A1( us32_n482 ) , .ZN( us32_n694 ) );
  NOR3_X1 us32_U99 (.ZN( us32_n480 ) , .A2( us32_n508 ) , .A3( us32_n601 ) , .A1( us32_n610 ) );
endmodule

