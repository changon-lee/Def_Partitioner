module des_des_die_5 ( u0_FP_33, u0_FP_34, u0_FP_36, u0_FP_37, u0_FP_38, u0_FP_39, u0_FP_40, u0_FP_41, u0_FP_42, 
       u0_FP_43, u0_FP_45, u0_FP_48, u0_FP_49, u0_FP_64, u0_K13_8, u0_K14_42, u0_K16_11, u0_K16_18, 
       u0_K16_24, u0_K16_8, u0_K1_31, u0_K1_47, u0_K2_5, u0_K2_6, u0_K2_8, u0_K6_11, u0_K6_13, 
       u0_K6_20, u0_K6_23, u0_K8_19, u0_K8_23, u0_R0_4, u0_R0_5, u0_R11_28, u0_R11_3, u0_R11_32, 
       u0_R11_4, u0_R11_5, u0_R11_6, u0_R11_7, u0_R11_8, u0_R11_9, u0_R12_1, u0_R12_20, u0_R12_21, 
       u0_R12_22, u0_R12_23, u0_R12_24, u0_R12_25, u0_R12_26, u0_R12_28, u0_R12_29, u0_R12_30, u0_R12_32, 
       u0_R2_1, u0_R2_10, u0_R2_11, u0_R2_12, u0_R2_13, u0_R2_3, u0_R2_32, u0_R2_4, u0_R2_6, 
       u0_R2_7, u0_R2_8, u0_R2_9, u0_R4_13, u0_R4_14, u0_R4_16, u0_R4_8, u0_R6_1, u0_R6_12, 
       u0_R6_13, u0_R6_14, u0_R6_16, u0_R6_17, u0_R6_18, u0_R6_20, u0_R6_21, u0_R6_23, u0_R6_24, 
       u0_R6_28, u0_R6_29, u0_R6_32, u0_R9_10, u0_R9_11, u0_R9_12, u0_R9_13, u0_R9_15, u0_R9_16, 
       u0_R9_17, u0_R9_8, u0_R9_9, u0_desIn_r_1, u0_desIn_r_11, u0_desIn_r_25, u0_desIn_r_27, u0_desIn_r_3, u0_desIn_r_33, 
       u0_desIn_r_51, u0_desIn_r_57, u0_desIn_r_59, u0_desIn_r_7, u0_key_r_14, u0_key_r_16, u0_key_r_2, u0_key_r_21, u0_key_r_23, 
       u0_key_r_28, u0_key_r_30, u0_key_r_31, u0_key_r_35, u0_key_r_36, u0_key_r_37, u0_key_r_38, u0_key_r_42, u0_key_r_43, 
       u0_key_r_50, u0_key_r_51, u0_key_r_9, u0_u0_X_25, u0_u0_X_28, u0_u0_X_30, u0_u0_X_32, u0_u0_X_33, u0_u0_X_39, 
       u0_u0_X_40, u0_u0_X_45, u0_u0_X_46, u0_u10_X_21, u0_u12_X_2, u0_u12_X_3, u0_u12_X_44, u0_u12_X_45, u0_u12_X_46, 
       u0_u12_X_48, u0_u13_X_40, u0_u13_X_46, u0_u15_X_17, u0_u15_X_19, u0_u15_X_21, u0_u15_X_22, u0_u15_X_4, u0_u1_X_1, 
       u0_u1_X_10, u0_u1_X_11, u0_u1_X_12, u0_u1_X_2, u0_u1_X_3, u0_u1_X_4, u0_u1_X_9, u0_u3_X_3, u0_u3_X_6, 
       u0_u3_X_8, u0_u5_X_10, u0_u5_X_12, u0_u5_X_14, u0_u5_X_15, u0_u5_X_16, u0_u5_X_17, u0_u5_X_19, u0_u5_X_22, 
       u0_u5_X_24, u0_u5_X_26, u0_u5_X_27, u0_u5_X_28, u0_u5_X_29, u0_u5_X_30, u0_u5_X_7, u0_u5_X_8, u0_u5_X_9, 
       u0_u7_X_22, u0_u7_X_28, u0_u7_X_33, u0_u7_X_36, u0_u7_X_45, u0_u7_X_46, u0_uk_K_r11_17, u0_uk_K_r11_25, u0_uk_K_r11_29, 
       u0_uk_K_r11_34, u0_uk_K_r11_48, u0_uk_K_r11_53, u0_uk_K_r11_54, u0_uk_K_r12_15, u0_uk_K_r12_16, u0_uk_K_r14_11, u0_uk_K_r14_12, u0_uk_K_r14_18, 
       u0_uk_K_r14_46, u0_uk_K_r2_13, u0_uk_K_r2_18, u0_uk_K_r2_20, u0_uk_K_r2_25, u0_uk_K_r2_27, u0_uk_K_r2_53, u0_uk_K_r6_0, u0_uk_K_r6_14, 
       u0_uk_K_r6_21, u0_uk_K_r6_29, u0_uk_K_r9_13, u0_uk_K_r9_19, u0_uk_K_r9_27, u0_uk_n10, u0_uk_n100, u0_uk_n1000, u0_uk_n1001, 
       u0_uk_n1002, u0_uk_n102, u0_uk_n106, u0_uk_n109, u0_uk_n11, u0_uk_n115, u0_uk_n117, u0_uk_n118, u0_uk_n121, 
       u0_uk_n126, u0_uk_n127, u0_uk_n128, u0_uk_n129, u0_uk_n131, u0_uk_n141, u0_uk_n142, u0_uk_n145, u0_uk_n146, 
       u0_uk_n161, u0_uk_n163, u0_uk_n182, u0_uk_n187, u0_uk_n188, u0_uk_n190, u0_uk_n196, u0_uk_n197, u0_uk_n200, 
       u0_uk_n201, u0_uk_n202, u0_uk_n203, u0_uk_n206, u0_uk_n208, u0_uk_n212, u0_uk_n213, u0_uk_n214, u0_uk_n215, 
       u0_uk_n217, u0_uk_n220, u0_uk_n221, u0_uk_n223, u0_uk_n240, u0_uk_n242, u0_uk_n251, u0_uk_n257, u0_uk_n27, 
       u0_uk_n318, u0_uk_n320, u0_uk_n321, u0_uk_n325, u0_uk_n327, u0_uk_n330, u0_uk_n331, u0_uk_n332, u0_uk_n333, 
       u0_uk_n336, u0_uk_n337, u0_uk_n341, u0_uk_n347, u0_uk_n348, u0_uk_n354, u0_uk_n355, u0_uk_n358, u0_uk_n359, 
       u0_uk_n418, u0_uk_n434, u0_uk_n497, u0_uk_n50, u0_uk_n502, u0_uk_n51, u0_uk_n510, u0_uk_n517, u0_uk_n519, 
       u0_uk_n52, u0_uk_n525, u0_uk_n529, u0_uk_n530, u0_uk_n531, u0_uk_n534, u0_uk_n535, u0_uk_n536, u0_uk_n55, 
       u0_uk_n56, u0_uk_n58, u0_uk_n59, u0_uk_n61, u0_uk_n629, u0_uk_n630, u0_uk_n631, u0_uk_n636, u0_uk_n637, 
       u0_uk_n639, u0_uk_n640, u0_uk_n644, u0_uk_n645, u0_uk_n65, u0_uk_n651, u0_uk_n652, u0_uk_n653, u0_uk_n659, 
       u0_uk_n660, u0_uk_n664, u0_uk_n667, u0_uk_n668, u0_uk_n67, u0_uk_n68, u0_uk_n73, u0_uk_n746, u0_uk_n755, 
       u0_uk_n77, u0_uk_n797, u0_uk_n799, u0_uk_n81, u0_uk_n82, u0_uk_n828, u0_uk_n83, u0_uk_n839, u0_uk_n855, 
       u0_uk_n88, u0_uk_n89, u0_uk_n90, u0_uk_n92, u0_uk_n93, u0_uk_n933, u0_uk_n934, u0_uk_n939, u0_uk_n94, 
       u0_uk_n940, u0_uk_n96, u0_uk_n960, u0_uk_n99, u0_uk_n999, u1_FP_34, u1_FP_35, u1_FP_37, u1_FP_38, 
       u1_FP_39, u1_K10_15, u1_K10_16, u1_K10_17, u1_K10_18, u1_K10_19, u1_K10_20, u1_K10_21, u1_K10_45, 
       u1_K10_46, u1_K11_10, u1_K11_11, u1_K11_13, u1_K11_15, u1_K11_16, u1_K11_9, u1_K12_10, u1_K12_11, 
       u1_K12_12, u1_K12_13, u1_K12_14, u1_K12_16, u1_K12_5, u1_K12_7, u1_K12_9, u1_K13_1, u1_K13_24, 
       u1_K13_26, u1_K13_27, u1_K13_28, u1_K13_3, u1_K13_4, u1_K13_45, u1_K13_46, u1_K13_47, u1_K15_14, 
       u1_K15_15, u1_K15_16, u1_K15_17, u1_K15_18, u1_K15_19, u1_K15_20, u1_K15_21, u1_K15_22, u1_K16_10, 
       u1_K16_3, u1_K16_4, u1_K16_6, u1_K16_8, u1_K16_9, u1_K1_21, u1_K1_3, u1_K1_4, u1_K2_33, 
       u1_K2_34, u1_K3_10, u1_K3_3, u1_K3_4, u1_K3_5, u1_K3_7, u1_K3_9, u1_K4_45, u1_K4_46, 
       u1_K5_10, u1_K5_9, u1_K6_1, u1_K6_22, u1_K6_3, u1_K6_33, u1_K6_34, u1_K6_35, u1_K6_36, 
       u1_K6_37, u1_K6_38, u1_K6_39, u1_K6_40, u1_K6_41, u1_K6_42, u1_K6_43, u1_K6_44, u1_K6_45, 
       u1_K6_46, u1_K6_47, u1_K6_48, u1_K6_6, u1_K6_8, u1_K8_45, u1_K8_46, u1_R0_22, u1_R0_23, 
       u1_R10_10, u1_R10_11, u1_R10_2, u1_R10_3, u1_R10_4, u1_R10_6, u1_R10_7, u1_R10_8, u1_R10_9, 
       u1_R11_14, u1_R11_15, u1_R11_17, u1_R11_18, u1_R11_19, u1_R11_2, u1_R11_3, u1_R11_30, u1_R11_31, 
       u1_R11_32, u1_R11_5, u1_R13_10, u1_R13_11, u1_R13_12, u1_R13_13, u1_R13_14, u1_R13_15, u1_R13_9, 
       u1_R1_2, u1_R1_3, u1_R1_4, u1_R1_6, u1_R1_7, u1_R2_30, u1_R2_31, u1_R3_6, u1_R3_7, 
       u1_R4_1, u1_R4_14, u1_R4_15, u1_R4_2, u1_R4_22, u1_R4_23, u1_R4_24, u1_R4_25, u1_R4_26, 
       u1_R4_27, u1_R4_28, u1_R4_29, u1_R4_3, u1_R4_30, u1_R4_31, u1_R4_32, u1_R4_5, u1_R4_6, 
       u1_R4_7, u1_R6_30, u1_R6_31, u1_R7_6, u1_R7_7, u1_R7_8, u1_R8_10, u1_R8_11, u1_R8_12, 
       u1_R8_13, u1_R8_14, u1_R8_15, u1_R8_30, u1_R8_31, u1_R9_10, u1_R9_11, u1_R9_5, u1_R9_6, 
       u1_R9_7, u1_R9_8, u1_R9_9, u1_desIn_r_15, u1_desIn_r_23, u1_desIn_r_45, u1_desIn_r_53, u1_u0_X_1, u1_u0_X_19, 
       u1_u0_X_2, u1_u0_X_20, u1_u0_X_23, u1_u0_X_24, u1_u0_X_5, u1_u0_X_6, u1_u10_X_17, u1_u10_X_18, u1_u10_X_7, 
       u1_u11_X_1, u1_u11_X_17, u1_u11_X_18, u1_u11_X_2, u1_u11_X_6, u1_u11_X_8, u1_u12_X_19, u1_u12_X_2, u1_u12_X_20, 
       u1_u12_X_23, u1_u12_X_25, u1_u12_X_29, u1_u12_X_30, u1_u12_X_43, u1_u12_X_44, u1_u12_X_48, u1_u12_X_5, u1_u14_X_13, 
       u1_u14_X_23, u1_u14_X_24, u1_u15_X_1, u1_u15_X_11, u1_u15_X_12, u1_u15_X_2, u1_u15_X_5, u1_u15_X_7, u1_u1_X_31, 
       u1_u1_X_32, u1_u1_X_35, u1_u1_X_36, u1_u2_X_1, u1_u2_X_11, u1_u2_X_12, u1_u2_X_2, u1_u2_X_6, u1_u2_X_8, 
       u1_u3_X_43, u1_u3_X_44, u1_u3_X_47, u1_u3_X_48, u1_u4_X_11, u1_u4_X_12, u1_u4_X_7, u1_u4_X_8, u1_u5_X_11, 
       u1_u5_X_12, u1_u5_X_19, u1_u5_X_20, u1_u5_X_23, u1_u5_X_24, u1_u5_X_31, u1_u5_X_32, u1_u5_X_5, u1_u5_X_7, 
       u1_u7_X_43, u1_u7_X_44, u1_u7_X_47, u1_u7_X_48, u1_u8_X_12, u1_u8_X_7, u1_u8_X_8, u1_u9_X_13, u1_u9_X_14, 
       u1_u9_X_23, u1_u9_X_24, u1_u9_X_43, u1_u9_X_44, u1_u9_X_47, u1_u9_X_48, u1_uk_n1004, u1_uk_n1088, u1_uk_n1092, 
       u1_uk_n1096, u1_uk_n1101, u1_uk_n1104, u1_uk_n1147, u1_uk_n1148, u1_uk_n1171, u1_uk_n312, u1_uk_n379, u1_uk_n382, 
       u1_uk_n501, u1_uk_n504, u1_uk_n601, u1_uk_n656, u1_uk_n689, u1_uk_n692, u1_uk_n949, u2_K10_36, u2_K15_29, 
       u2_K15_31, u2_K15_35, u2_K1_30, u2_K1_37, u2_K1_43, u2_R13_17, u2_R13_18, u2_R13_20, u2_R13_22, 
       u2_R13_24, u2_R13_25, u2_R8_20, u2_R8_22, u2_R8_24, u2_R8_25, u2_desIn_r_1, u2_desIn_r_11, u2_desIn_r_25, 
       u2_desIn_r_27, u2_desIn_r_3, u2_desIn_r_33, u2_desIn_r_35, u2_desIn_r_43, u2_desIn_r_57, u2_desIn_r_59, u2_desIn_r_61, u2_desIn_r_7, 
       u2_desIn_r_9, u2_key_r_0, u2_key_r_14, u2_key_r_16, u2_key_r_21, u2_key_r_22, u2_key_r_23, u2_key_r_28, u2_key_r_29, 
       u2_key_r_30, u2_key_r_31, u2_key_r_35, u2_key_r_36, u2_key_r_37, u2_key_r_42, u2_key_r_43, u2_key_r_44, u2_key_r_51, 
       u2_key_r_7, u2_u0_X_28, u2_u0_X_34, u2_u0_X_40, u2_u0_X_45, u2_u0_X_46, u2_u14_X_25, u2_u14_X_28, u2_u14_X_30, 
       u2_u14_X_32, u2_u14_X_34, u2_u9_X_32, u2_u9_X_34, u2_uk_K_r8_16, u2_uk_K_r8_2, u2_uk_K_r8_22, u2_uk_K_r8_37, u2_uk_K_r8_42, 
       u2_uk_n10, u2_uk_n100, u2_uk_n102, u2_uk_n109, u2_uk_n117, u2_uk_n118, u2_uk_n128, u2_uk_n142, u2_uk_n155, 
       u2_uk_n1615, u2_uk_n162, u2_uk_n163, u2_uk_n164, u2_uk_n1817, u2_uk_n182, u2_uk_n1826, u2_uk_n1835, u2_uk_n1840, 
       u2_uk_n203, u2_uk_n207, u2_uk_n208, u2_uk_n217, u2_uk_n222, u2_uk_n238, u2_uk_n31, u2_uk_n60, u2_uk_n63, 
       u2_uk_n92, u2_uk_n939, u2_uk_n94, u2_uk_n942, u2_uk_n984, u2_uk_n986, u2_uk_n99, u0_out0_11, u0_out0_12, u0_out0_14, u0_out0_15, u0_out0_19, u0_out0_21, u0_out0_22, u0_out0_25, u0_out0_27, 
        u0_out0_29, u0_out0_3, u0_out0_32, u0_out0_4, u0_out0_5, u0_out0_7, u0_out0_8, u0_out10_1, u0_out10_10, 
        u0_out10_16, u0_out10_20, u0_out10_24, u0_out10_26, u0_out10_30, u0_out10_6, u0_out12_13, u0_out12_15, u0_out12_17, 
        u0_out12_18, u0_out12_2, u0_out12_21, u0_out12_23, u0_out12_27, u0_out12_28, u0_out12_31, u0_out12_5, u0_out12_9, 
        u0_out13_11, u0_out13_12, u0_out13_15, u0_out13_19, u0_out13_21, u0_out13_22, u0_out13_27, u0_out13_29, u0_out13_32, 
        u0_out13_4, u0_out13_5, u0_out13_7, u0_out15_1, u0_out15_10, u0_out15_13, u0_out15_16, u0_out15_17, u0_out15_18, 
        u0_out15_2, u0_out15_20, u0_out15_23, u0_out15_24, u0_out15_26, u0_out15_28, u0_out15_30, u0_out15_31, u0_out15_6, 
        u0_out15_9, u0_out1_13, u0_out1_17, u0_out1_18, u0_out1_2, u0_out1_23, u0_out1_28, u0_out1_31, u0_out1_9, 
        u0_out3_13, u0_out3_16, u0_out3_17, u0_out3_18, u0_out3_2, u0_out3_23, u0_out3_24, u0_out3_28, u0_out3_30, 
        u0_out3_31, u0_out3_6, u0_out3_9, u0_out5_1, u0_out5_10, u0_out5_13, u0_out5_14, u0_out5_16, u0_out5_18, 
        u0_out5_2, u0_out5_20, u0_out5_24, u0_out5_25, u0_out5_26, u0_out5_28, u0_out5_3, u0_out5_30, u0_out5_6, 
        u0_out5_8, u0_out7_1, u0_out7_10, u0_out7_11, u0_out7_14, u0_out7_15, u0_out7_19, u0_out7_20, u0_out7_21, 
        u0_out7_25, u0_out7_26, u0_out7_27, u0_out7_29, u0_out7_3, u0_out7_4, u0_out7_5, u0_out7_8, u0_uk_n110, 
        u0_uk_n147, u0_uk_n155, u0_uk_n164, u0_uk_n17, u0_uk_n207, u0_uk_n222, u0_uk_n230, u0_uk_n231, u0_uk_n238, 
        u0_uk_n250, u0_uk_n252, u0_uk_n31, u0_uk_n60, u0_uk_n687, u0_uk_n707, u1_out0_1, u1_out0_10, u1_out0_17, 
        u1_out0_20, u1_out0_23, u1_out0_26, u1_out0_31, u1_out0_9, u1_out10_13, u1_out10_16, u1_out10_18, u1_out10_2, 
        u1_out10_24, u1_out10_28, u1_out10_30, u1_out10_6, u1_out11_13, u1_out11_16, u1_out11_17, u1_out11_18, u1_out11_2, 
        u1_out11_23, u1_out11_24, u1_out11_28, u1_out11_30, u1_out11_31, u1_out11_6, u1_out11_9, u1_out12_1, u1_out12_10, 
        u1_out12_14, u1_out12_15, u1_out12_17, u1_out12_20, u1_out12_21, u1_out12_23, u1_out12_25, u1_out12_26, u1_out12_27, 
        u1_out12_3, u1_out12_31, u1_out12_5, u1_out12_8, u1_out12_9, u1_out14_1, u1_out14_10, u1_out14_16, u1_out14_20, 
        u1_out14_24, u1_out14_26, u1_out14_30, u1_out14_6, u1_out15_13, u1_out15_17, u1_out15_18, u1_out15_2, u1_out15_23, 
        u1_out15_28, u1_out15_31, u1_out15_9, u1_out1_11, u1_out1_19, u1_out1_29, u1_out1_4, u1_out2_13, u1_out2_17, 
        u1_out2_18, u1_out2_2, u1_out2_23, u1_out2_28, u1_out2_31, u1_out2_9, u1_out3_15, u1_out3_21, u1_out3_27, 
        u1_out3_5, u1_out4_13, u1_out4_18, u1_out4_2, u1_out4_28, u1_out5_1, u1_out5_10, u1_out5_11, u1_out5_12, 
        u1_out5_13, u1_out5_15, u1_out5_17, u1_out5_18, u1_out5_19, u1_out5_2, u1_out5_20, u1_out5_21, u1_out5_22, 
        u1_out5_23, u1_out5_26, u1_out5_27, u1_out5_28, u1_out5_29, u1_out5_31, u1_out5_32, u1_out5_4, u1_out5_5, 
        u1_out5_7, u1_out5_9, u1_out7_15, u1_out7_21, u1_out7_27, u1_out7_5, u1_out8_13, u1_out8_18, u1_out8_2, 
        u1_out8_28, u1_out9_1, u1_out9_10, u1_out9_15, u1_out9_16, u1_out9_20, u1_out9_21, u1_out9_24, u1_out9_26, 
        u1_out9_27, u1_out9_30, u1_out9_5, u1_out9_6, u2_out0_11, u2_out0_12, u2_out0_14, u2_out0_15, u2_out0_19, 
        u2_out0_21, u2_out0_22, u2_out0_25, u2_out0_27, u2_out0_29, u2_out0_3, u2_out0_32, u2_out0_4, u2_out0_5, 
        u2_out0_7, u2_out0_8, u2_out14_11, u2_out14_14, u2_out14_19, u2_out14_25, u2_out14_29, u2_out14_3, u2_out14_4, 
        u2_out14_8, u2_out9_11, u2_out9_19, u2_out9_29, u2_out9_4, u2_uk_n1142, u2_uk_n1152, u2_uk_n1171, u2_uk_n1178 );
  input u0_FP_33, u0_FP_34, u0_FP_36, u0_FP_37, u0_FP_38, u0_FP_39, u0_FP_40, u0_FP_41, u0_FP_42, 
        u0_FP_43, u0_FP_45, u0_FP_48, u0_FP_49, u0_FP_64, u0_K13_8, u0_K14_42, u0_K16_11, u0_K16_18, 
        u0_K16_24, u0_K16_8, u0_K1_31, u0_K1_47, u0_K2_5, u0_K2_6, u0_K2_8, u0_K6_11, u0_K6_13, 
        u0_K6_20, u0_K6_23, u0_K8_19, u0_K8_23, u0_R0_4, u0_R0_5, u0_R11_28, u0_R11_3, u0_R11_32, 
        u0_R11_4, u0_R11_5, u0_R11_6, u0_R11_7, u0_R11_8, u0_R11_9, u0_R12_1, u0_R12_20, u0_R12_21, 
        u0_R12_22, u0_R12_23, u0_R12_24, u0_R12_25, u0_R12_26, u0_R12_28, u0_R12_29, u0_R12_30, u0_R12_32, 
        u0_R2_1, u0_R2_10, u0_R2_11, u0_R2_12, u0_R2_13, u0_R2_3, u0_R2_32, u0_R2_4, u0_R2_6, 
        u0_R2_7, u0_R2_8, u0_R2_9, u0_R4_13, u0_R4_14, u0_R4_16, u0_R4_8, u0_R6_1, u0_R6_12, 
        u0_R6_13, u0_R6_14, u0_R6_16, u0_R6_17, u0_R6_18, u0_R6_20, u0_R6_21, u0_R6_23, u0_R6_24, 
        u0_R6_28, u0_R6_29, u0_R6_32, u0_R9_10, u0_R9_11, u0_R9_12, u0_R9_13, u0_R9_15, u0_R9_16, 
        u0_R9_17, u0_R9_8, u0_R9_9, u0_desIn_r_1, u0_desIn_r_11, u0_desIn_r_25, u0_desIn_r_27, u0_desIn_r_3, u0_desIn_r_33, 
        u0_desIn_r_51, u0_desIn_r_57, u0_desIn_r_59, u0_desIn_r_7, u0_key_r_14, u0_key_r_16, u0_key_r_2, u0_key_r_21, u0_key_r_23, 
        u0_key_r_28, u0_key_r_30, u0_key_r_31, u0_key_r_35, u0_key_r_36, u0_key_r_37, u0_key_r_38, u0_key_r_42, u0_key_r_43, 
        u0_key_r_50, u0_key_r_51, u0_key_r_9, u0_u0_X_25, u0_u0_X_28, u0_u0_X_30, u0_u0_X_32, u0_u0_X_33, u0_u0_X_39, 
        u0_u0_X_40, u0_u0_X_45, u0_u0_X_46, u0_u10_X_21, u0_u12_X_2, u0_u12_X_3, u0_u12_X_44, u0_u12_X_45, u0_u12_X_46, 
        u0_u12_X_48, u0_u13_X_40, u0_u13_X_46, u0_u15_X_17, u0_u15_X_19, u0_u15_X_21, u0_u15_X_22, u0_u15_X_4, u0_u1_X_1, 
        u0_u1_X_10, u0_u1_X_11, u0_u1_X_12, u0_u1_X_2, u0_u1_X_3, u0_u1_X_4, u0_u1_X_9, u0_u3_X_3, u0_u3_X_6, 
        u0_u3_X_8, u0_u5_X_10, u0_u5_X_12, u0_u5_X_14, u0_u5_X_15, u0_u5_X_16, u0_u5_X_17, u0_u5_X_19, u0_u5_X_22, 
        u0_u5_X_24, u0_u5_X_26, u0_u5_X_27, u0_u5_X_28, u0_u5_X_29, u0_u5_X_30, u0_u5_X_7, u0_u5_X_8, u0_u5_X_9, 
        u0_u7_X_22, u0_u7_X_28, u0_u7_X_33, u0_u7_X_36, u0_u7_X_45, u0_u7_X_46, u0_uk_K_r11_17, u0_uk_K_r11_25, u0_uk_K_r11_29, 
        u0_uk_K_r11_34, u0_uk_K_r11_48, u0_uk_K_r11_53, u0_uk_K_r11_54, u0_uk_K_r12_15, u0_uk_K_r12_16, u0_uk_K_r14_11, u0_uk_K_r14_12, u0_uk_K_r14_18, 
        u0_uk_K_r14_46, u0_uk_K_r2_13, u0_uk_K_r2_18, u0_uk_K_r2_20, u0_uk_K_r2_25, u0_uk_K_r2_27, u0_uk_K_r2_53, u0_uk_K_r6_0, u0_uk_K_r6_14, 
        u0_uk_K_r6_21, u0_uk_K_r6_29, u0_uk_K_r9_13, u0_uk_K_r9_19, u0_uk_K_r9_27, u0_uk_n10, u0_uk_n100, u0_uk_n1000, u0_uk_n1001, 
        u0_uk_n1002, u0_uk_n102, u0_uk_n106, u0_uk_n109, u0_uk_n11, u0_uk_n115, u0_uk_n117, u0_uk_n118, u0_uk_n121, 
        u0_uk_n126, u0_uk_n127, u0_uk_n128, u0_uk_n129, u0_uk_n131, u0_uk_n141, u0_uk_n142, u0_uk_n145, u0_uk_n146, 
        u0_uk_n161, u0_uk_n163, u0_uk_n182, u0_uk_n187, u0_uk_n188, u0_uk_n190, u0_uk_n196, u0_uk_n197, u0_uk_n200, 
        u0_uk_n201, u0_uk_n202, u0_uk_n203, u0_uk_n206, u0_uk_n208, u0_uk_n212, u0_uk_n213, u0_uk_n214, u0_uk_n215, 
        u0_uk_n217, u0_uk_n220, u0_uk_n221, u0_uk_n223, u0_uk_n240, u0_uk_n242, u0_uk_n251, u0_uk_n257, u0_uk_n27, 
        u0_uk_n318, u0_uk_n320, u0_uk_n321, u0_uk_n325, u0_uk_n327, u0_uk_n330, u0_uk_n331, u0_uk_n332, u0_uk_n333, 
        u0_uk_n336, u0_uk_n337, u0_uk_n341, u0_uk_n347, u0_uk_n348, u0_uk_n354, u0_uk_n355, u0_uk_n358, u0_uk_n359, 
        u0_uk_n418, u0_uk_n434, u0_uk_n497, u0_uk_n50, u0_uk_n502, u0_uk_n51, u0_uk_n510, u0_uk_n517, u0_uk_n519, 
        u0_uk_n52, u0_uk_n525, u0_uk_n529, u0_uk_n530, u0_uk_n531, u0_uk_n534, u0_uk_n535, u0_uk_n536, u0_uk_n55, 
        u0_uk_n56, u0_uk_n58, u0_uk_n59, u0_uk_n61, u0_uk_n629, u0_uk_n630, u0_uk_n631, u0_uk_n636, u0_uk_n637, 
        u0_uk_n639, u0_uk_n640, u0_uk_n644, u0_uk_n645, u0_uk_n65, u0_uk_n651, u0_uk_n652, u0_uk_n653, u0_uk_n659, 
        u0_uk_n660, u0_uk_n664, u0_uk_n667, u0_uk_n668, u0_uk_n67, u0_uk_n68, u0_uk_n73, u0_uk_n746, u0_uk_n755, 
        u0_uk_n77, u0_uk_n797, u0_uk_n799, u0_uk_n81, u0_uk_n82, u0_uk_n828, u0_uk_n83, u0_uk_n839, u0_uk_n855, 
        u0_uk_n88, u0_uk_n89, u0_uk_n90, u0_uk_n92, u0_uk_n93, u0_uk_n933, u0_uk_n934, u0_uk_n939, u0_uk_n94, 
        u0_uk_n940, u0_uk_n96, u0_uk_n960, u0_uk_n99, u0_uk_n999, u1_FP_34, u1_FP_35, u1_FP_37, u1_FP_38, 
        u1_FP_39, u1_K10_15, u1_K10_16, u1_K10_17, u1_K10_18, u1_K10_19, u1_K10_20, u1_K10_21, u1_K10_45, 
        u1_K10_46, u1_K11_10, u1_K11_11, u1_K11_13, u1_K11_15, u1_K11_16, u1_K11_9, u1_K12_10, u1_K12_11, 
        u1_K12_12, u1_K12_13, u1_K12_14, u1_K12_16, u1_K12_5, u1_K12_7, u1_K12_9, u1_K13_1, u1_K13_24, 
        u1_K13_26, u1_K13_27, u1_K13_28, u1_K13_3, u1_K13_4, u1_K13_45, u1_K13_46, u1_K13_47, u1_K15_14, 
        u1_K15_15, u1_K15_16, u1_K15_17, u1_K15_18, u1_K15_19, u1_K15_20, u1_K15_21, u1_K15_22, u1_K16_10, 
        u1_K16_3, u1_K16_4, u1_K16_6, u1_K16_8, u1_K16_9, u1_K1_21, u1_K1_3, u1_K1_4, u1_K2_33, 
        u1_K2_34, u1_K3_10, u1_K3_3, u1_K3_4, u1_K3_5, u1_K3_7, u1_K3_9, u1_K4_45, u1_K4_46, 
        u1_K5_10, u1_K5_9, u1_K6_1, u1_K6_22, u1_K6_3, u1_K6_33, u1_K6_34, u1_K6_35, u1_K6_36, 
        u1_K6_37, u1_K6_38, u1_K6_39, u1_K6_40, u1_K6_41, u1_K6_42, u1_K6_43, u1_K6_44, u1_K6_45, 
        u1_K6_46, u1_K6_47, u1_K6_48, u1_K6_6, u1_K6_8, u1_K8_45, u1_K8_46, u1_R0_22, u1_R0_23, 
        u1_R10_10, u1_R10_11, u1_R10_2, u1_R10_3, u1_R10_4, u1_R10_6, u1_R10_7, u1_R10_8, u1_R10_9, 
        u1_R11_14, u1_R11_15, u1_R11_17, u1_R11_18, u1_R11_19, u1_R11_2, u1_R11_3, u1_R11_30, u1_R11_31, 
        u1_R11_32, u1_R11_5, u1_R13_10, u1_R13_11, u1_R13_12, u1_R13_13, u1_R13_14, u1_R13_15, u1_R13_9, 
        u1_R1_2, u1_R1_3, u1_R1_4, u1_R1_6, u1_R1_7, u1_R2_30, u1_R2_31, u1_R3_6, u1_R3_7, 
        u1_R4_1, u1_R4_14, u1_R4_15, u1_R4_2, u1_R4_22, u1_R4_23, u1_R4_24, u1_R4_25, u1_R4_26, 
        u1_R4_27, u1_R4_28, u1_R4_29, u1_R4_3, u1_R4_30, u1_R4_31, u1_R4_32, u1_R4_5, u1_R4_6, 
        u1_R4_7, u1_R6_30, u1_R6_31, u1_R7_6, u1_R7_7, u1_R7_8, u1_R8_10, u1_R8_11, u1_R8_12, 
        u1_R8_13, u1_R8_14, u1_R8_15, u1_R8_30, u1_R8_31, u1_R9_10, u1_R9_11, u1_R9_5, u1_R9_6, 
        u1_R9_7, u1_R9_8, u1_R9_9, u1_desIn_r_15, u1_desIn_r_23, u1_desIn_r_45, u1_desIn_r_53, u1_u0_X_1, u1_u0_X_19, 
        u1_u0_X_2, u1_u0_X_20, u1_u0_X_23, u1_u0_X_24, u1_u0_X_5, u1_u0_X_6, u1_u10_X_17, u1_u10_X_18, u1_u10_X_7, 
        u1_u11_X_1, u1_u11_X_17, u1_u11_X_18, u1_u11_X_2, u1_u11_X_6, u1_u11_X_8, u1_u12_X_19, u1_u12_X_2, u1_u12_X_20, 
        u1_u12_X_23, u1_u12_X_25, u1_u12_X_29, u1_u12_X_30, u1_u12_X_43, u1_u12_X_44, u1_u12_X_48, u1_u12_X_5, u1_u14_X_13, 
        u1_u14_X_23, u1_u14_X_24, u1_u15_X_1, u1_u15_X_11, u1_u15_X_12, u1_u15_X_2, u1_u15_X_5, u1_u15_X_7, u1_u1_X_31, 
        u1_u1_X_32, u1_u1_X_35, u1_u1_X_36, u1_u2_X_1, u1_u2_X_11, u1_u2_X_12, u1_u2_X_2, u1_u2_X_6, u1_u2_X_8, 
        u1_u3_X_43, u1_u3_X_44, u1_u3_X_47, u1_u3_X_48, u1_u4_X_11, u1_u4_X_12, u1_u4_X_7, u1_u4_X_8, u1_u5_X_11, 
        u1_u5_X_12, u1_u5_X_19, u1_u5_X_20, u1_u5_X_23, u1_u5_X_24, u1_u5_X_31, u1_u5_X_32, u1_u5_X_5, u1_u5_X_7, 
        u1_u7_X_43, u1_u7_X_44, u1_u7_X_47, u1_u7_X_48, u1_u8_X_12, u1_u8_X_7, u1_u8_X_8, u1_u9_X_13, u1_u9_X_14, 
        u1_u9_X_23, u1_u9_X_24, u1_u9_X_43, u1_u9_X_44, u1_u9_X_47, u1_u9_X_48, u1_uk_n1004, u1_uk_n1088, u1_uk_n1092, 
        u1_uk_n1096, u1_uk_n1101, u1_uk_n1104, u1_uk_n1147, u1_uk_n1148, u1_uk_n1171, u1_uk_n312, u1_uk_n379, u1_uk_n382, 
        u1_uk_n501, u1_uk_n504, u1_uk_n601, u1_uk_n656, u1_uk_n689, u1_uk_n692, u1_uk_n949, u2_K10_36, u2_K15_29, 
        u2_K15_31, u2_K15_35, u2_K1_30, u2_K1_37, u2_K1_43, u2_R13_17, u2_R13_18, u2_R13_20, u2_R13_22, 
        u2_R13_24, u2_R13_25, u2_R8_20, u2_R8_22, u2_R8_24, u2_R8_25, u2_desIn_r_1, u2_desIn_r_11, u2_desIn_r_25, 
        u2_desIn_r_27, u2_desIn_r_3, u2_desIn_r_33, u2_desIn_r_35, u2_desIn_r_43, u2_desIn_r_57, u2_desIn_r_59, u2_desIn_r_61, u2_desIn_r_7, 
        u2_desIn_r_9, u2_key_r_0, u2_key_r_14, u2_key_r_16, u2_key_r_21, u2_key_r_22, u2_key_r_23, u2_key_r_28, u2_key_r_29, 
        u2_key_r_30, u2_key_r_31, u2_key_r_35, u2_key_r_36, u2_key_r_37, u2_key_r_42, u2_key_r_43, u2_key_r_44, u2_key_r_51, 
        u2_key_r_7, u2_u0_X_28, u2_u0_X_34, u2_u0_X_40, u2_u0_X_45, u2_u0_X_46, u2_u14_X_25, u2_u14_X_28, u2_u14_X_30, 
        u2_u14_X_32, u2_u14_X_34, u2_u9_X_32, u2_u9_X_34, u2_uk_K_r8_16, u2_uk_K_r8_2, u2_uk_K_r8_22, u2_uk_K_r8_37, u2_uk_K_r8_42, 
        u2_uk_n10, u2_uk_n100, u2_uk_n102, u2_uk_n109, u2_uk_n117, u2_uk_n118, u2_uk_n128, u2_uk_n142, u2_uk_n155, 
        u2_uk_n1615, u2_uk_n162, u2_uk_n163, u2_uk_n164, u2_uk_n1817, u2_uk_n182, u2_uk_n1826, u2_uk_n1835, u2_uk_n1840, 
        u2_uk_n203, u2_uk_n207, u2_uk_n208, u2_uk_n217, u2_uk_n222, u2_uk_n238, u2_uk_n31, u2_uk_n60, u2_uk_n63, 
        u2_uk_n92, u2_uk_n939, u2_uk_n94, u2_uk_n942, u2_uk_n984, u2_uk_n986, u2_uk_n99;
  output u0_out0_11, u0_out0_12, u0_out0_14, u0_out0_15, u0_out0_19, u0_out0_21, u0_out0_22, u0_out0_25, u0_out0_27, 
        u0_out0_29, u0_out0_3, u0_out0_32, u0_out0_4, u0_out0_5, u0_out0_7, u0_out0_8, u0_out10_1, u0_out10_10, 
        u0_out10_16, u0_out10_20, u0_out10_24, u0_out10_26, u0_out10_30, u0_out10_6, u0_out12_13, u0_out12_15, u0_out12_17, 
        u0_out12_18, u0_out12_2, u0_out12_21, u0_out12_23, u0_out12_27, u0_out12_28, u0_out12_31, u0_out12_5, u0_out12_9, 
        u0_out13_11, u0_out13_12, u0_out13_15, u0_out13_19, u0_out13_21, u0_out13_22, u0_out13_27, u0_out13_29, u0_out13_32, 
        u0_out13_4, u0_out13_5, u0_out13_7, u0_out15_1, u0_out15_10, u0_out15_13, u0_out15_16, u0_out15_17, u0_out15_18, 
        u0_out15_2, u0_out15_20, u0_out15_23, u0_out15_24, u0_out15_26, u0_out15_28, u0_out15_30, u0_out15_31, u0_out15_6, 
        u0_out15_9, u0_out1_13, u0_out1_17, u0_out1_18, u0_out1_2, u0_out1_23, u0_out1_28, u0_out1_31, u0_out1_9, 
        u0_out3_13, u0_out3_16, u0_out3_17, u0_out3_18, u0_out3_2, u0_out3_23, u0_out3_24, u0_out3_28, u0_out3_30, 
        u0_out3_31, u0_out3_6, u0_out3_9, u0_out5_1, u0_out5_10, u0_out5_13, u0_out5_14, u0_out5_16, u0_out5_18, 
        u0_out5_2, u0_out5_20, u0_out5_24, u0_out5_25, u0_out5_26, u0_out5_28, u0_out5_3, u0_out5_30, u0_out5_6, 
        u0_out5_8, u0_out7_1, u0_out7_10, u0_out7_11, u0_out7_14, u0_out7_15, u0_out7_19, u0_out7_20, u0_out7_21, 
        u0_out7_25, u0_out7_26, u0_out7_27, u0_out7_29, u0_out7_3, u0_out7_4, u0_out7_5, u0_out7_8, u0_uk_n110, 
        u0_uk_n147, u0_uk_n155, u0_uk_n164, u0_uk_n17, u0_uk_n207, u0_uk_n222, u0_uk_n230, u0_uk_n231, u0_uk_n238, 
        u0_uk_n250, u0_uk_n252, u0_uk_n31, u0_uk_n60, u0_uk_n687, u0_uk_n707, u1_out0_1, u1_out0_10, u1_out0_17, 
        u1_out0_20, u1_out0_23, u1_out0_26, u1_out0_31, u1_out0_9, u1_out10_13, u1_out10_16, u1_out10_18, u1_out10_2, 
        u1_out10_24, u1_out10_28, u1_out10_30, u1_out10_6, u1_out11_13, u1_out11_16, u1_out11_17, u1_out11_18, u1_out11_2, 
        u1_out11_23, u1_out11_24, u1_out11_28, u1_out11_30, u1_out11_31, u1_out11_6, u1_out11_9, u1_out12_1, u1_out12_10, 
        u1_out12_14, u1_out12_15, u1_out12_17, u1_out12_20, u1_out12_21, u1_out12_23, u1_out12_25, u1_out12_26, u1_out12_27, 
        u1_out12_3, u1_out12_31, u1_out12_5, u1_out12_8, u1_out12_9, u1_out14_1, u1_out14_10, u1_out14_16, u1_out14_20, 
        u1_out14_24, u1_out14_26, u1_out14_30, u1_out14_6, u1_out15_13, u1_out15_17, u1_out15_18, u1_out15_2, u1_out15_23, 
        u1_out15_28, u1_out15_31, u1_out15_9, u1_out1_11, u1_out1_19, u1_out1_29, u1_out1_4, u1_out2_13, u1_out2_17, 
        u1_out2_18, u1_out2_2, u1_out2_23, u1_out2_28, u1_out2_31, u1_out2_9, u1_out3_15, u1_out3_21, u1_out3_27, 
        u1_out3_5, u1_out4_13, u1_out4_18, u1_out4_2, u1_out4_28, u1_out5_1, u1_out5_10, u1_out5_11, u1_out5_12, 
        u1_out5_13, u1_out5_15, u1_out5_17, u1_out5_18, u1_out5_19, u1_out5_2, u1_out5_20, u1_out5_21, u1_out5_22, 
        u1_out5_23, u1_out5_26, u1_out5_27, u1_out5_28, u1_out5_29, u1_out5_31, u1_out5_32, u1_out5_4, u1_out5_5, 
        u1_out5_7, u1_out5_9, u1_out7_15, u1_out7_21, u1_out7_27, u1_out7_5, u1_out8_13, u1_out8_18, u1_out8_2, 
        u1_out8_28, u1_out9_1, u1_out9_10, u1_out9_15, u1_out9_16, u1_out9_20, u1_out9_21, u1_out9_24, u1_out9_26, 
        u1_out9_27, u1_out9_30, u1_out9_5, u1_out9_6, u2_out0_11, u2_out0_12, u2_out0_14, u2_out0_15, u2_out0_19, 
        u2_out0_21, u2_out0_22, u2_out0_25, u2_out0_27, u2_out0_29, u2_out0_3, u2_out0_32, u2_out0_4, u2_out0_5, 
        u2_out0_7, u2_out0_8, u2_out14_11, u2_out14_14, u2_out14_19, u2_out14_25, u2_out14_29, u2_out14_3, u2_out14_4, 
        u2_out14_8, u2_out9_11, u2_out9_19, u2_out9_29, u2_out9_4, u2_uk_n1142, u2_uk_n1152, u2_uk_n1171, u2_uk_n1178;
  wire u0_K11_13, u0_K11_14, u0_K11_15, u0_K11_16, u0_K11_17, u0_K11_18, u0_K11_19, u0_K11_20, u0_K11_22, 
       u0_K11_23, u0_K11_24, u0_K13_1, u0_K13_10, u0_K13_11, u0_K13_12, u0_K13_4, u0_K13_43, u0_K13_47, 
       u0_K13_5, u0_K13_6, u0_K13_7, u0_K13_9, u0_K14_31, u0_K14_32, u0_K14_33, u0_K14_34, u0_K14_35, 
       u0_K14_36, u0_K14_37, u0_K14_38, u0_K14_39, u0_K14_41, u0_K14_43, u0_K14_44, u0_K14_45, u0_K14_47, 
       u0_K14_48, u0_K16_1, u0_K16_10, u0_K16_12, u0_K16_13, u0_K16_14, u0_K16_15, u0_K16_16, u0_K16_2, 
       u0_K16_20, u0_K16_23, u0_K16_3, u0_K16_5, u0_K16_6, u0_K16_7, u0_K16_9, u0_K1_26, u0_K1_27, 
       u0_K1_29, u0_K1_34, u0_K1_35, u0_K1_36, u0_K1_37, u0_K1_38, u0_K1_41, u0_K1_42, u0_K1_43, 
       u0_K1_44, u0_K1_48, u0_K2_7, u0_K4_1, u0_K4_10, u0_K4_11, u0_K4_12, u0_K4_13, u0_K4_14, 
       u0_K4_15, u0_K4_16, u0_K4_17, u0_K4_18, u0_K4_2, u0_K4_4, u0_K4_5, u0_K4_7, u0_K4_9, 
       u0_K6_18, u0_K6_21, u0_K6_25, u0_K8_20, u0_K8_21, u0_K8_24, u0_K8_25, u0_K8_26, u0_K8_27, 
       u0_K8_29, u0_K8_30, u0_K8_31, u0_K8_32, u0_K8_34, u0_K8_35, u0_K8_43, u0_K8_44, u0_K8_47, 
       u0_K8_48, u0_u0_X_26, u0_u0_X_27, u0_u0_X_29, u0_u0_X_31, u0_u0_X_34, u0_u0_X_35, u0_u0_X_36, u0_u0_X_37, 
       u0_u0_X_38, u0_u0_X_41, u0_u0_X_42, u0_u0_X_43, u0_u0_X_44, u0_u0_X_47, u0_u0_X_48, u0_u0_u4_n1, u0_u0_u4_n10, 
       u0_u0_u4_n11, u0_u0_u4_n12, u0_u0_u4_n13, u0_u0_u4_n14, u0_u0_u4_n15, u0_u0_u4_n16, u0_u0_u4_n17, u0_u0_u4_n18, u0_u0_u4_n19, 
       u0_u0_u4_n2, u0_u0_u4_n20, u0_u0_u4_n21, u0_u0_u4_n22, u0_u0_u4_n23, u0_u0_u4_n24, u0_u0_u4_n25, u0_u0_u4_n26, u0_u0_u4_n27, 
       u0_u0_u4_n28, u0_u0_u4_n29, u0_u0_u4_n3, u0_u0_u4_n30, u0_u0_u4_n31, u0_u0_u4_n32, u0_u0_u4_n33, u0_u0_u4_n34, u0_u0_u4_n35, 
       u0_u0_u4_n36, u0_u0_u4_n37, u0_u0_u4_n38, u0_u0_u4_n39, u0_u0_u4_n4, u0_u0_u4_n40, u0_u0_u4_n41, u0_u0_u4_n42, u0_u0_u4_n43, 
       u0_u0_u4_n44, u0_u0_u4_n45, u0_u0_u4_n46, u0_u0_u4_n47, u0_u0_u4_n48, u0_u0_u4_n49, u0_u0_u4_n5, u0_u0_u4_n50, u0_u0_u4_n51, 
       u0_u0_u4_n52, u0_u0_u4_n53, u0_u0_u4_n54, u0_u0_u4_n55, u0_u0_u4_n56, u0_u0_u4_n57, u0_u0_u4_n58, u0_u0_u4_n59, u0_u0_u4_n6, 
       u0_u0_u4_n60, u0_u0_u4_n61, u0_u0_u4_n62, u0_u0_u4_n63, u0_u0_u4_n64, u0_u0_u4_n65, u0_u0_u4_n66, u0_u0_u4_n67, u0_u0_u4_n68, 
       u0_u0_u4_n69, u0_u0_u4_n7, u0_u0_u4_n70, u0_u0_u4_n71, u0_u0_u4_n72, u0_u0_u4_n73, u0_u0_u4_n74, u0_u0_u4_n75, u0_u0_u4_n76, 
       u0_u0_u4_n77, u0_u0_u4_n78, u0_u0_u4_n79, u0_u0_u4_n8, u0_u0_u4_n80, u0_u0_u4_n81, u0_u0_u4_n82, u0_u0_u4_n83, u0_u0_u4_n84, 
       u0_u0_u4_n85, u0_u0_u4_n86, u0_u0_u4_n87, u0_u0_u4_n88, u0_u0_u4_n89, u0_u0_u4_n9, u0_u0_u4_n90, u0_u0_u4_n91, u0_u0_u4_n92, 
       u0_u0_u4_n93, u0_u0_u5_n1, u0_u0_u5_n10, u0_u0_u5_n11, u0_u0_u5_n12, u0_u0_u5_n13, u0_u0_u5_n14, u0_u0_u5_n15, u0_u0_u5_n16, 
       u0_u0_u5_n17, u0_u0_u5_n18, u0_u0_u5_n19, u0_u0_u5_n2, u0_u0_u5_n20, u0_u0_u5_n21, u0_u0_u5_n22, u0_u0_u5_n23, u0_u0_u5_n24, 
       u0_u0_u5_n25, u0_u0_u5_n26, u0_u0_u5_n27, u0_u0_u5_n28, u0_u0_u5_n29, u0_u0_u5_n3, u0_u0_u5_n30, u0_u0_u5_n31, u0_u0_u5_n32, 
       u0_u0_u5_n33, u0_u0_u5_n34, u0_u0_u5_n35, u0_u0_u5_n36, u0_u0_u5_n37, u0_u0_u5_n38, u0_u0_u5_n39, u0_u0_u5_n4, u0_u0_u5_n40, 
       u0_u0_u5_n41, u0_u0_u5_n42, u0_u0_u5_n43, u0_u0_u5_n44, u0_u0_u5_n45, u0_u0_u5_n46, u0_u0_u5_n47, u0_u0_u5_n48, u0_u0_u5_n49, 
       u0_u0_u5_n5, u0_u0_u5_n50, u0_u0_u5_n51, u0_u0_u5_n52, u0_u0_u5_n53, u0_u0_u5_n54, u0_u0_u5_n55, u0_u0_u5_n56, u0_u0_u5_n57, 
       u0_u0_u5_n58, u0_u0_u5_n59, u0_u0_u5_n6, u0_u0_u5_n60, u0_u0_u5_n61, u0_u0_u5_n62, u0_u0_u5_n63, u0_u0_u5_n64, u0_u0_u5_n65, 
       u0_u0_u5_n66, u0_u0_u5_n67, u0_u0_u5_n68, u0_u0_u5_n69, u0_u0_u5_n7, u0_u0_u5_n70, u0_u0_u5_n71, u0_u0_u5_n72, u0_u0_u5_n73, 
       u0_u0_u5_n74, u0_u0_u5_n75, u0_u0_u5_n76, u0_u0_u5_n77, u0_u0_u5_n78, u0_u0_u5_n79, u0_u0_u5_n8, u0_u0_u5_n80, u0_u0_u5_n81, 
       u0_u0_u5_n82, u0_u0_u5_n83, u0_u0_u5_n84, u0_u0_u5_n85, u0_u0_u5_n86, u0_u0_u5_n87, u0_u0_u5_n88, u0_u0_u5_n89, u0_u0_u5_n9, 
       u0_u0_u5_n90, u0_u0_u5_n91, u0_u0_u5_n92, u0_u0_u5_n93, u0_u0_u5_n94, u0_u0_u5_n95, u0_u0_u5_n96, u0_u0_u5_n97, u0_u0_u5_n98, 
       u0_u0_u6_n1, u0_u0_u6_n10, u0_u0_u6_n11, u0_u0_u6_n12, u0_u0_u6_n13, u0_u0_u6_n14, u0_u0_u6_n15, u0_u0_u6_n16, u0_u0_u6_n17, 
       u0_u0_u6_n18, u0_u0_u6_n19, u0_u0_u6_n2, u0_u0_u6_n20, u0_u0_u6_n21, u0_u0_u6_n22, u0_u0_u6_n23, u0_u0_u6_n24, u0_u0_u6_n25, 
       u0_u0_u6_n26, u0_u0_u6_n27, u0_u0_u6_n28, u0_u0_u6_n29, u0_u0_u6_n3, u0_u0_u6_n30, u0_u0_u6_n31, u0_u0_u6_n32, u0_u0_u6_n33, 
       u0_u0_u6_n34, u0_u0_u6_n35, u0_u0_u6_n36, u0_u0_u6_n37, u0_u0_u6_n38, u0_u0_u6_n39, u0_u0_u6_n4, u0_u0_u6_n40, u0_u0_u6_n41, 
       u0_u0_u6_n42, u0_u0_u6_n43, u0_u0_u6_n44, u0_u0_u6_n45, u0_u0_u6_n46, u0_u0_u6_n47, u0_u0_u6_n48, u0_u0_u6_n49, u0_u0_u6_n5, 
       u0_u0_u6_n50, u0_u0_u6_n51, u0_u0_u6_n52, u0_u0_u6_n53, u0_u0_u6_n54, u0_u0_u6_n55, u0_u0_u6_n56, u0_u0_u6_n57, u0_u0_u6_n58, 
       u0_u0_u6_n59, u0_u0_u6_n6, u0_u0_u6_n60, u0_u0_u6_n61, u0_u0_u6_n62, u0_u0_u6_n63, u0_u0_u6_n64, u0_u0_u6_n65, u0_u0_u6_n66, 
       u0_u0_u6_n67, u0_u0_u6_n68, u0_u0_u6_n69, u0_u0_u6_n7, u0_u0_u6_n70, u0_u0_u6_n71, u0_u0_u6_n72, u0_u0_u6_n73, u0_u0_u6_n74, 
       u0_u0_u6_n75, u0_u0_u6_n76, u0_u0_u6_n77, u0_u0_u6_n78, u0_u0_u6_n79, u0_u0_u6_n8, u0_u0_u6_n80, u0_u0_u6_n81, u0_u0_u6_n82, 
       u0_u0_u6_n83, u0_u0_u6_n84, u0_u0_u6_n85, u0_u0_u6_n86, u0_u0_u6_n87, u0_u0_u6_n9, u0_u0_u7_n1, u0_u0_u7_n10, u0_u0_u7_n11, 
       u0_u0_u7_n12, u0_u0_u7_n13, u0_u0_u7_n14, u0_u0_u7_n15, u0_u0_u7_n16, u0_u0_u7_n17, u0_u0_u7_n18, u0_u0_u7_n19, u0_u0_u7_n2, 
       u0_u0_u7_n20, u0_u0_u7_n21, u0_u0_u7_n22, u0_u0_u7_n23, u0_u0_u7_n24, u0_u0_u7_n25, u0_u0_u7_n26, u0_u0_u7_n27, u0_u0_u7_n28, 
       u0_u0_u7_n29, u0_u0_u7_n3, u0_u0_u7_n30, u0_u0_u7_n31, u0_u0_u7_n32, u0_u0_u7_n33, u0_u0_u7_n34, u0_u0_u7_n35, u0_u0_u7_n36, 
       u0_u0_u7_n37, u0_u0_u7_n38, u0_u0_u7_n39, u0_u0_u7_n4, u0_u0_u7_n40, u0_u0_u7_n41, u0_u0_u7_n42, u0_u0_u7_n43, u0_u0_u7_n44, 
       u0_u0_u7_n45, u0_u0_u7_n46, u0_u0_u7_n47, u0_u0_u7_n48, u0_u0_u7_n49, u0_u0_u7_n5, u0_u0_u7_n50, u0_u0_u7_n51, u0_u0_u7_n52, 
       u0_u0_u7_n53, u0_u0_u7_n54, u0_u0_u7_n55, u0_u0_u7_n56, u0_u0_u7_n57, u0_u0_u7_n58, u0_u0_u7_n59, u0_u0_u7_n6, u0_u0_u7_n60, 
       u0_u0_u7_n61, u0_u0_u7_n62, u0_u0_u7_n63, u0_u0_u7_n64, u0_u0_u7_n65, u0_u0_u7_n66, u0_u0_u7_n67, u0_u0_u7_n68, u0_u0_u7_n69, 
       u0_u0_u7_n7, u0_u0_u7_n70, u0_u0_u7_n71, u0_u0_u7_n72, u0_u0_u7_n73, u0_u0_u7_n74, u0_u0_u7_n75, u0_u0_u7_n76, u0_u0_u7_n77, 
       u0_u0_u7_n78, u0_u0_u7_n79, u0_u0_u7_n8, u0_u0_u7_n80, u0_u0_u7_n81, u0_u0_u7_n82, u0_u0_u7_n83, u0_u0_u7_n84, u0_u0_u7_n85, 
       u0_u0_u7_n86, u0_u0_u7_n87, u0_u0_u7_n88, u0_u0_u7_n89, u0_u0_u7_n9, u0_u0_u7_n90, u0_u10_X_13, u0_u10_X_14, u0_u10_X_15, 
       u0_u10_X_16, u0_u10_X_17, u0_u10_X_18, u0_u10_X_19, u0_u10_X_20, u0_u10_X_22, u0_u10_X_23, u0_u10_X_24, u0_u10_u2_n100, 
       u0_u10_u2_n101, u0_u10_u2_n102, u0_u10_u2_n103, u0_u10_u2_n104, u0_u10_u2_n105, u0_u10_u2_n106, u0_u10_u2_n107, u0_u10_u2_n108, u0_u10_u2_n109, 
       u0_u10_u2_n110, u0_u10_u2_n111, u0_u10_u2_n112, u0_u10_u2_n113, u0_u10_u2_n114, u0_u10_u2_n115, u0_u10_u2_n116, u0_u10_u2_n117, u0_u10_u2_n118, 
       u0_u10_u2_n119, u0_u10_u2_n120, u0_u10_u2_n121, u0_u10_u2_n122, u0_u10_u2_n123, u0_u10_u2_n124, u0_u10_u2_n125, u0_u10_u2_n126, u0_u10_u2_n127, 
       u0_u10_u2_n128, u0_u10_u2_n129, u0_u10_u2_n130, u0_u10_u2_n131, u0_u10_u2_n132, u0_u10_u2_n133, u0_u10_u2_n134, u0_u10_u2_n135, u0_u10_u2_n136, 
       u0_u10_u2_n137, u0_u10_u2_n138, u0_u10_u2_n139, u0_u10_u2_n140, u0_u10_u2_n141, u0_u10_u2_n142, u0_u10_u2_n143, u0_u10_u2_n144, u0_u10_u2_n145, 
       u0_u10_u2_n146, u0_u10_u2_n147, u0_u10_u2_n148, u0_u10_u2_n149, u0_u10_u2_n150, u0_u10_u2_n151, u0_u10_u2_n152, u0_u10_u2_n153, u0_u10_u2_n154, 
       u0_u10_u2_n155, u0_u10_u2_n156, u0_u10_u2_n157, u0_u10_u2_n158, u0_u10_u2_n159, u0_u10_u2_n160, u0_u10_u2_n161, u0_u10_u2_n162, u0_u10_u2_n163, 
       u0_u10_u2_n164, u0_u10_u2_n165, u0_u10_u2_n166, u0_u10_u2_n167, u0_u10_u2_n168, u0_u10_u2_n169, u0_u10_u2_n170, u0_u10_u2_n171, u0_u10_u2_n172, 
       u0_u10_u2_n173, u0_u10_u2_n174, u0_u10_u2_n175, u0_u10_u2_n176, u0_u10_u2_n177, u0_u10_u2_n178, u0_u10_u2_n179, u0_u10_u2_n180, u0_u10_u2_n181, 
       u0_u10_u2_n182, u0_u10_u2_n183, u0_u10_u2_n184, u0_u10_u2_n185, u0_u10_u2_n186, u0_u10_u2_n187, u0_u10_u2_n188, u0_u10_u2_n95, u0_u10_u2_n96, 
       u0_u10_u2_n97, u0_u10_u2_n98, u0_u10_u2_n99, u0_u10_u3_n100, u0_u10_u3_n101, u0_u10_u3_n102, u0_u10_u3_n103, u0_u10_u3_n104, u0_u10_u3_n105, 
       u0_u10_u3_n106, u0_u10_u3_n107, u0_u10_u3_n108, u0_u10_u3_n109, u0_u10_u3_n110, u0_u10_u3_n111, u0_u10_u3_n112, u0_u10_u3_n113, u0_u10_u3_n114, 
       u0_u10_u3_n115, u0_u10_u3_n116, u0_u10_u3_n117, u0_u10_u3_n118, u0_u10_u3_n119, u0_u10_u3_n120, u0_u10_u3_n121, u0_u10_u3_n122, u0_u10_u3_n123, 
       u0_u10_u3_n124, u0_u10_u3_n125, u0_u10_u3_n126, u0_u10_u3_n127, u0_u10_u3_n128, u0_u10_u3_n129, u0_u10_u3_n130, u0_u10_u3_n131, u0_u10_u3_n132, 
       u0_u10_u3_n133, u0_u10_u3_n134, u0_u10_u3_n135, u0_u10_u3_n136, u0_u10_u3_n137, u0_u10_u3_n138, u0_u10_u3_n139, u0_u10_u3_n140, u0_u10_u3_n141, 
       u0_u10_u3_n142, u0_u10_u3_n143, u0_u10_u3_n144, u0_u10_u3_n145, u0_u10_u3_n146, u0_u10_u3_n147, u0_u10_u3_n148, u0_u10_u3_n149, u0_u10_u3_n150, 
       u0_u10_u3_n151, u0_u10_u3_n152, u0_u10_u3_n153, u0_u10_u3_n154, u0_u10_u3_n155, u0_u10_u3_n156, u0_u10_u3_n157, u0_u10_u3_n158, u0_u10_u3_n159, 
       u0_u10_u3_n160, u0_u10_u3_n161, u0_u10_u3_n162, u0_u10_u3_n163, u0_u10_u3_n164, u0_u10_u3_n165, u0_u10_u3_n166, u0_u10_u3_n167, u0_u10_u3_n168, 
       u0_u10_u3_n169, u0_u10_u3_n170, u0_u10_u3_n171, u0_u10_u3_n172, u0_u10_u3_n173, u0_u10_u3_n174, u0_u10_u3_n175, u0_u10_u3_n176, u0_u10_u3_n177, 
       u0_u10_u3_n178, u0_u10_u3_n179, u0_u10_u3_n180, u0_u10_u3_n181, u0_u10_u3_n182, u0_u10_u3_n183, u0_u10_u3_n184, u0_u10_u3_n185, u0_u10_u3_n186, 
       u0_u10_u3_n94, u0_u10_u3_n95, u0_u10_u3_n96, u0_u10_u3_n97, u0_u10_u3_n98, u0_u10_u3_n99, u0_u12_X_1, u0_u12_X_10, u0_u12_X_11, 
       u0_u12_X_12, u0_u12_X_4, u0_u12_X_43, u0_u12_X_47, u0_u12_X_5, u0_u12_X_6, u0_u12_X_7, u0_u12_X_8, u0_u12_X_9, 
       u0_u12_u0_n100, u0_u12_u0_n101, u0_u12_u0_n102, u0_u12_u0_n103, u0_u12_u0_n104, u0_u12_u0_n105, u0_u12_u0_n106, u0_u12_u0_n107, u0_u12_u0_n108, 
       u0_u12_u0_n109, u0_u12_u0_n110, u0_u12_u0_n111, u0_u12_u0_n112, u0_u12_u0_n113, u0_u12_u0_n114, u0_u12_u0_n115, u0_u12_u0_n116, u0_u12_u0_n117, 
       u0_u12_u0_n118, u0_u12_u0_n119, u0_u12_u0_n120, u0_u12_u0_n121, u0_u12_u0_n122, u0_u12_u0_n123, u0_u12_u0_n124, u0_u12_u0_n125, u0_u12_u0_n126, 
       u0_u12_u0_n127, u0_u12_u0_n128, u0_u12_u0_n129, u0_u12_u0_n130, u0_u12_u0_n131, u0_u12_u0_n132, u0_u12_u0_n133, u0_u12_u0_n134, u0_u12_u0_n135, 
       u0_u12_u0_n136, u0_u12_u0_n137, u0_u12_u0_n138, u0_u12_u0_n139, u0_u12_u0_n140, u0_u12_u0_n141, u0_u12_u0_n142, u0_u12_u0_n143, u0_u12_u0_n144, 
       u0_u12_u0_n145, u0_u12_u0_n146, u0_u12_u0_n147, u0_u12_u0_n148, u0_u12_u0_n149, u0_u12_u0_n150, u0_u12_u0_n151, u0_u12_u0_n152, u0_u12_u0_n153, 
       u0_u12_u0_n154, u0_u12_u0_n155, u0_u12_u0_n156, u0_u12_u0_n157, u0_u12_u0_n158, u0_u12_u0_n159, u0_u12_u0_n160, u0_u12_u0_n161, u0_u12_u0_n162, 
       u0_u12_u0_n163, u0_u12_u0_n164, u0_u12_u0_n165, u0_u12_u0_n166, u0_u12_u0_n167, u0_u12_u0_n168, u0_u12_u0_n169, u0_u12_u0_n170, u0_u12_u0_n171, 
       u0_u12_u0_n172, u0_u12_u0_n173, u0_u12_u0_n174, u0_u12_u0_n88, u0_u12_u0_n89, u0_u12_u0_n90, u0_u12_u0_n91, u0_u12_u0_n92, u0_u12_u0_n93, 
       u0_u12_u0_n94, u0_u12_u0_n95, u0_u12_u0_n96, u0_u12_u0_n97, u0_u12_u0_n98, u0_u12_u0_n99, u0_u12_u1_n100, u0_u12_u1_n101, u0_u12_u1_n102, 
       u0_u12_u1_n103, u0_u12_u1_n104, u0_u12_u1_n105, u0_u12_u1_n106, u0_u12_u1_n107, u0_u12_u1_n108, u0_u12_u1_n109, u0_u12_u1_n110, u0_u12_u1_n111, 
       u0_u12_u1_n112, u0_u12_u1_n113, u0_u12_u1_n114, u0_u12_u1_n115, u0_u12_u1_n116, u0_u12_u1_n117, u0_u12_u1_n118, u0_u12_u1_n119, u0_u12_u1_n120, 
       u0_u12_u1_n121, u0_u12_u1_n122, u0_u12_u1_n123, u0_u12_u1_n124, u0_u12_u1_n125, u0_u12_u1_n126, u0_u12_u1_n127, u0_u12_u1_n128, u0_u12_u1_n129, 
       u0_u12_u1_n130, u0_u12_u1_n131, u0_u12_u1_n132, u0_u12_u1_n133, u0_u12_u1_n134, u0_u12_u1_n135, u0_u12_u1_n136, u0_u12_u1_n137, u0_u12_u1_n138, 
       u0_u12_u1_n139, u0_u12_u1_n140, u0_u12_u1_n141, u0_u12_u1_n142, u0_u12_u1_n143, u0_u12_u1_n144, u0_u12_u1_n145, u0_u12_u1_n146, u0_u12_u1_n147, 
       u0_u12_u1_n148, u0_u12_u1_n149, u0_u12_u1_n150, u0_u12_u1_n151, u0_u12_u1_n152, u0_u12_u1_n153, u0_u12_u1_n154, u0_u12_u1_n155, u0_u12_u1_n156, 
       u0_u12_u1_n157, u0_u12_u1_n158, u0_u12_u1_n159, u0_u12_u1_n160, u0_u12_u1_n161, u0_u12_u1_n162, u0_u12_u1_n163, u0_u12_u1_n164, u0_u12_u1_n165, 
       u0_u12_u1_n166, u0_u12_u1_n167, u0_u12_u1_n168, u0_u12_u1_n169, u0_u12_u1_n170, u0_u12_u1_n171, u0_u12_u1_n172, u0_u12_u1_n173, u0_u12_u1_n174, 
       u0_u12_u1_n175, u0_u12_u1_n176, u0_u12_u1_n177, u0_u12_u1_n178, u0_u12_u1_n179, u0_u12_u1_n180, u0_u12_u1_n181, u0_u12_u1_n182, u0_u12_u1_n183, 
       u0_u12_u1_n184, u0_u12_u1_n185, u0_u12_u1_n186, u0_u12_u1_n187, u0_u12_u1_n188, u0_u12_u1_n95, u0_u12_u1_n96, u0_u12_u1_n97, u0_u12_u1_n98, 
       u0_u12_u1_n99, u0_u12_u7_n100, u0_u12_u7_n101, u0_u12_u7_n102, u0_u12_u7_n103, u0_u12_u7_n104, u0_u12_u7_n105, u0_u12_u7_n106, u0_u12_u7_n107, 
       u0_u12_u7_n108, u0_u12_u7_n109, u0_u12_u7_n110, u0_u12_u7_n111, u0_u12_u7_n112, u0_u12_u7_n113, u0_u12_u7_n114, u0_u12_u7_n115, u0_u12_u7_n116, 
       u0_u12_u7_n117, u0_u12_u7_n118, u0_u12_u7_n119, u0_u12_u7_n120, u0_u12_u7_n121, u0_u12_u7_n122, u0_u12_u7_n123, u0_u12_u7_n124, u0_u12_u7_n125, 
       u0_u12_u7_n126, u0_u12_u7_n127, u0_u12_u7_n128, u0_u12_u7_n129, u0_u12_u7_n130, u0_u12_u7_n131, u0_u12_u7_n132, u0_u12_u7_n133, u0_u12_u7_n134, 
       u0_u12_u7_n135, u0_u12_u7_n136, u0_u12_u7_n137, u0_u12_u7_n138, u0_u12_u7_n139, u0_u12_u7_n140, u0_u12_u7_n141, u0_u12_u7_n142, u0_u12_u7_n143, 
       u0_u12_u7_n144, u0_u12_u7_n145, u0_u12_u7_n146, u0_u12_u7_n147, u0_u12_u7_n148, u0_u12_u7_n149, u0_u12_u7_n150, u0_u12_u7_n151, u0_u12_u7_n152, 
       u0_u12_u7_n153, u0_u12_u7_n154, u0_u12_u7_n155, u0_u12_u7_n156, u0_u12_u7_n157, u0_u12_u7_n158, u0_u12_u7_n159, u0_u12_u7_n160, u0_u12_u7_n161, 
       u0_u12_u7_n162, u0_u12_u7_n163, u0_u12_u7_n164, u0_u12_u7_n165, u0_u12_u7_n166, u0_u12_u7_n167, u0_u12_u7_n168, u0_u12_u7_n169, u0_u12_u7_n170, 
       u0_u12_u7_n171, u0_u12_u7_n172, u0_u12_u7_n173, u0_u12_u7_n174, u0_u12_u7_n175, u0_u12_u7_n176, u0_u12_u7_n177, u0_u12_u7_n178, u0_u12_u7_n179, 
       u0_u12_u7_n180, u0_u12_u7_n91, u0_u12_u7_n92, u0_u12_u7_n93, u0_u12_u7_n94, u0_u12_u7_n95, u0_u12_u7_n96, u0_u12_u7_n97, u0_u12_u7_n98, 
       u0_u12_u7_n99, u0_u13_X_31, u0_u13_X_32, u0_u13_X_33, u0_u13_X_34, u0_u13_X_35, u0_u13_X_36, u0_u13_X_37, u0_u13_X_38, 
       u0_u13_X_39, u0_u13_X_41, u0_u13_X_42, u0_u13_X_43, u0_u13_X_44, u0_u13_X_45, u0_u13_X_47, u0_u13_X_48, u0_u13_u5_n100, 
       u0_u13_u5_n101, u0_u13_u5_n102, u0_u13_u5_n103, u0_u13_u5_n104, u0_u13_u5_n105, u0_u13_u5_n106, u0_u13_u5_n107, u0_u13_u5_n108, u0_u13_u5_n109, 
       u0_u13_u5_n110, u0_u13_u5_n111, u0_u13_u5_n112, u0_u13_u5_n113, u0_u13_u5_n114, u0_u13_u5_n115, u0_u13_u5_n116, u0_u13_u5_n117, u0_u13_u5_n118, 
       u0_u13_u5_n119, u0_u13_u5_n120, u0_u13_u5_n121, u0_u13_u5_n122, u0_u13_u5_n123, u0_u13_u5_n124, u0_u13_u5_n125, u0_u13_u5_n126, u0_u13_u5_n127, 
       u0_u13_u5_n128, u0_u13_u5_n129, u0_u13_u5_n130, u0_u13_u5_n131, u0_u13_u5_n132, u0_u13_u5_n133, u0_u13_u5_n134, u0_u13_u5_n135, u0_u13_u5_n136, 
       u0_u13_u5_n137, u0_u13_u5_n138, u0_u13_u5_n139, u0_u13_u5_n140, u0_u13_u5_n141, u0_u13_u5_n142, u0_u13_u5_n143, u0_u13_u5_n144, u0_u13_u5_n145, 
       u0_u13_u5_n146, u0_u13_u5_n147, u0_u13_u5_n148, u0_u13_u5_n149, u0_u13_u5_n150, u0_u13_u5_n151, u0_u13_u5_n152, u0_u13_u5_n153, u0_u13_u5_n154, 
       u0_u13_u5_n155, u0_u13_u5_n156, u0_u13_u5_n157, u0_u13_u5_n158, u0_u13_u5_n159, u0_u13_u5_n160, u0_u13_u5_n161, u0_u13_u5_n162, u0_u13_u5_n163, 
       u0_u13_u5_n164, u0_u13_u5_n165, u0_u13_u5_n166, u0_u13_u5_n167, u0_u13_u5_n168, u0_u13_u5_n169, u0_u13_u5_n170, u0_u13_u5_n171, u0_u13_u5_n172, 
       u0_u13_u5_n173, u0_u13_u5_n174, u0_u13_u5_n175, u0_u13_u5_n176, u0_u13_u5_n177, u0_u13_u5_n178, u0_u13_u5_n179, u0_u13_u5_n180, u0_u13_u5_n181, 
       u0_u13_u5_n182, u0_u13_u5_n183, u0_u13_u5_n184, u0_u13_u5_n185, u0_u13_u5_n186, u0_u13_u5_n187, u0_u13_u5_n188, u0_u13_u5_n189, u0_u13_u5_n190, 
       u0_u13_u5_n191, u0_u13_u5_n192, u0_u13_u5_n193, u0_u13_u5_n194, u0_u13_u5_n195, u0_u13_u5_n196, u0_u13_u5_n99, u0_u13_u6_n100, u0_u13_u6_n101, 
       u0_u13_u6_n102, u0_u13_u6_n103, u0_u13_u6_n104, u0_u13_u6_n105, u0_u13_u6_n106, u0_u13_u6_n107, u0_u13_u6_n108, u0_u13_u6_n109, u0_u13_u6_n110, 
       u0_u13_u6_n111, u0_u13_u6_n112, u0_u13_u6_n113, u0_u13_u6_n114, u0_u13_u6_n115, u0_u13_u6_n116, u0_u13_u6_n117, u0_u13_u6_n118, u0_u13_u6_n119, 
       u0_u13_u6_n120, u0_u13_u6_n121, u0_u13_u6_n122, u0_u13_u6_n123, u0_u13_u6_n124, u0_u13_u6_n125, u0_u13_u6_n126, u0_u13_u6_n127, u0_u13_u6_n128, 
       u0_u13_u6_n129, u0_u13_u6_n130, u0_u13_u6_n131, u0_u13_u6_n132, u0_u13_u6_n133, u0_u13_u6_n134, u0_u13_u6_n135, u0_u13_u6_n136, u0_u13_u6_n137, 
       u0_u13_u6_n138, u0_u13_u6_n139, u0_u13_u6_n140, u0_u13_u6_n141, u0_u13_u6_n142, u0_u13_u6_n143, u0_u13_u6_n144, u0_u13_u6_n145, u0_u13_u6_n146, 
       u0_u13_u6_n147, u0_u13_u6_n148, u0_u13_u6_n149, u0_u13_u6_n150, u0_u13_u6_n151, u0_u13_u6_n152, u0_u13_u6_n153, u0_u13_u6_n154, u0_u13_u6_n155, 
       u0_u13_u6_n156, u0_u13_u6_n157, u0_u13_u6_n158, u0_u13_u6_n159, u0_u13_u6_n160, u0_u13_u6_n161, u0_u13_u6_n162, u0_u13_u6_n163, u0_u13_u6_n164, 
       u0_u13_u6_n165, u0_u13_u6_n166, u0_u13_u6_n167, u0_u13_u6_n168, u0_u13_u6_n169, u0_u13_u6_n170, u0_u13_u6_n171, u0_u13_u6_n172, u0_u13_u6_n173, 
       u0_u13_u6_n174, u0_u13_u6_n88, u0_u13_u6_n89, u0_u13_u6_n90, u0_u13_u6_n91, u0_u13_u6_n92, u0_u13_u6_n93, u0_u13_u6_n94, u0_u13_u6_n95, 
       u0_u13_u6_n96, u0_u13_u6_n97, u0_u13_u6_n98, u0_u13_u6_n99, u0_u13_u7_n100, u0_u13_u7_n101, u0_u13_u7_n102, u0_u13_u7_n103, u0_u13_u7_n104, 
       u0_u13_u7_n105, u0_u13_u7_n106, u0_u13_u7_n107, u0_u13_u7_n108, u0_u13_u7_n109, u0_u13_u7_n110, u0_u13_u7_n111, u0_u13_u7_n112, u0_u13_u7_n113, 
       u0_u13_u7_n114, u0_u13_u7_n115, u0_u13_u7_n116, u0_u13_u7_n117, u0_u13_u7_n118, u0_u13_u7_n119, u0_u13_u7_n120, u0_u13_u7_n121, u0_u13_u7_n122, 
       u0_u13_u7_n123, u0_u13_u7_n124, u0_u13_u7_n125, u0_u13_u7_n126, u0_u13_u7_n127, u0_u13_u7_n128, u0_u13_u7_n129, u0_u13_u7_n130, u0_u13_u7_n131, 
       u0_u13_u7_n132, u0_u13_u7_n133, u0_u13_u7_n134, u0_u13_u7_n135, u0_u13_u7_n136, u0_u13_u7_n137, u0_u13_u7_n138, u0_u13_u7_n139, u0_u13_u7_n140, 
       u0_u13_u7_n141, u0_u13_u7_n142, u0_u13_u7_n143, u0_u13_u7_n144, u0_u13_u7_n145, u0_u13_u7_n146, u0_u13_u7_n147, u0_u13_u7_n148, u0_u13_u7_n149, 
       u0_u13_u7_n150, u0_u13_u7_n151, u0_u13_u7_n152, u0_u13_u7_n153, u0_u13_u7_n154, u0_u13_u7_n155, u0_u13_u7_n156, u0_u13_u7_n157, u0_u13_u7_n158, 
       u0_u13_u7_n159, u0_u13_u7_n160, u0_u13_u7_n161, u0_u13_u7_n162, u0_u13_u7_n163, u0_u13_u7_n164, u0_u13_u7_n165, u0_u13_u7_n166, u0_u13_u7_n167, 
       u0_u13_u7_n168, u0_u13_u7_n169, u0_u13_u7_n170, u0_u13_u7_n171, u0_u13_u7_n172, u0_u13_u7_n173, u0_u13_u7_n174, u0_u13_u7_n175, u0_u13_u7_n176, 
       u0_u13_u7_n177, u0_u13_u7_n178, u0_u13_u7_n179, u0_u13_u7_n180, u0_u13_u7_n91, u0_u13_u7_n92, u0_u13_u7_n93, u0_u13_u7_n94, u0_u13_u7_n95, 
       u0_u13_u7_n96, u0_u13_u7_n97, u0_u13_u7_n98, u0_u13_u7_n99, u0_u15_X_1, u0_u15_X_10, u0_u15_X_11, u0_u15_X_12, u0_u15_X_13, 
       u0_u15_X_14, u0_u15_X_15, u0_u15_X_16, u0_u15_X_18, u0_u15_X_2, u0_u15_X_20, u0_u15_X_23, u0_u15_X_24, u0_u15_X_3, 
       u0_u15_X_5, u0_u15_X_6, u0_u15_X_7, u0_u15_X_8, u0_u15_X_9, u0_u15_u0_n100, u0_u15_u0_n101, u0_u15_u0_n102, u0_u15_u0_n103, 
       u0_u15_u0_n104, u0_u15_u0_n105, u0_u15_u0_n106, u0_u15_u0_n107, u0_u15_u0_n108, u0_u15_u0_n109, u0_u15_u0_n110, u0_u15_u0_n111, u0_u15_u0_n112, 
       u0_u15_u0_n113, u0_u15_u0_n114, u0_u15_u0_n115, u0_u15_u0_n116, u0_u15_u0_n117, u0_u15_u0_n118, u0_u15_u0_n119, u0_u15_u0_n120, u0_u15_u0_n121, 
       u0_u15_u0_n122, u0_u15_u0_n123, u0_u15_u0_n124, u0_u15_u0_n125, u0_u15_u0_n126, u0_u15_u0_n127, u0_u15_u0_n128, u0_u15_u0_n129, u0_u15_u0_n130, 
       u0_u15_u0_n131, u0_u15_u0_n132, u0_u15_u0_n133, u0_u15_u0_n134, u0_u15_u0_n135, u0_u15_u0_n136, u0_u15_u0_n137, u0_u15_u0_n138, u0_u15_u0_n139, 
       u0_u15_u0_n140, u0_u15_u0_n141, u0_u15_u0_n142, u0_u15_u0_n143, u0_u15_u0_n144, u0_u15_u0_n145, u0_u15_u0_n146, u0_u15_u0_n147, u0_u15_u0_n148, 
       u0_u15_u0_n149, u0_u15_u0_n150, u0_u15_u0_n151, u0_u15_u0_n152, u0_u15_u0_n153, u0_u15_u0_n154, u0_u15_u0_n155, u0_u15_u0_n156, u0_u15_u0_n157, 
       u0_u15_u0_n158, u0_u15_u0_n159, u0_u15_u0_n160, u0_u15_u0_n161, u0_u15_u0_n162, u0_u15_u0_n163, u0_u15_u0_n164, u0_u15_u0_n165, u0_u15_u0_n166, 
       u0_u15_u0_n167, u0_u15_u0_n168, u0_u15_u0_n169, u0_u15_u0_n170, u0_u15_u0_n171, u0_u15_u0_n172, u0_u15_u0_n173, u0_u15_u0_n174, u0_u15_u0_n88, 
       u0_u15_u0_n89, u0_u15_u0_n90, u0_u15_u0_n91, u0_u15_u0_n92, u0_u15_u0_n93, u0_u15_u0_n94, u0_u15_u0_n95, u0_u15_u0_n96, u0_u15_u0_n97, 
       u0_u15_u0_n98, u0_u15_u0_n99, u0_u15_u1_n100, u0_u15_u1_n101, u0_u15_u1_n102, u0_u15_u1_n103, u0_u15_u1_n104, u0_u15_u1_n105, u0_u15_u1_n106, 
       u0_u15_u1_n107, u0_u15_u1_n108, u0_u15_u1_n109, u0_u15_u1_n110, u0_u15_u1_n111, u0_u15_u1_n112, u0_u15_u1_n113, u0_u15_u1_n114, u0_u15_u1_n115, 
       u0_u15_u1_n116, u0_u15_u1_n117, u0_u15_u1_n118, u0_u15_u1_n119, u0_u15_u1_n120, u0_u15_u1_n121, u0_u15_u1_n122, u0_u15_u1_n123, u0_u15_u1_n124, 
       u0_u15_u1_n125, u0_u15_u1_n126, u0_u15_u1_n127, u0_u15_u1_n128, u0_u15_u1_n129, u0_u15_u1_n130, u0_u15_u1_n131, u0_u15_u1_n132, u0_u15_u1_n133, 
       u0_u15_u1_n134, u0_u15_u1_n135, u0_u15_u1_n136, u0_u15_u1_n137, u0_u15_u1_n138, u0_u15_u1_n139, u0_u15_u1_n140, u0_u15_u1_n141, u0_u15_u1_n142, 
       u0_u15_u1_n143, u0_u15_u1_n144, u0_u15_u1_n145, u0_u15_u1_n146, u0_u15_u1_n147, u0_u15_u1_n148, u0_u15_u1_n149, u0_u15_u1_n150, u0_u15_u1_n151, 
       u0_u15_u1_n152, u0_u15_u1_n153, u0_u15_u1_n154, u0_u15_u1_n155, u0_u15_u1_n156, u0_u15_u1_n157, u0_u15_u1_n158, u0_u15_u1_n159, u0_u15_u1_n160, 
       u0_u15_u1_n161, u0_u15_u1_n162, u0_u15_u1_n163, u0_u15_u1_n164, u0_u15_u1_n165, u0_u15_u1_n166, u0_u15_u1_n167, u0_u15_u1_n168, u0_u15_u1_n169, 
       u0_u15_u1_n170, u0_u15_u1_n171, u0_u15_u1_n172, u0_u15_u1_n173, u0_u15_u1_n174, u0_u15_u1_n175, u0_u15_u1_n176, u0_u15_u1_n177, u0_u15_u1_n178, 
       u0_u15_u1_n179, u0_u15_u1_n180, u0_u15_u1_n181, u0_u15_u1_n182, u0_u15_u1_n183, u0_u15_u1_n184, u0_u15_u1_n185, u0_u15_u1_n186, u0_u15_u1_n187, 
       u0_u15_u1_n188, u0_u15_u1_n95, u0_u15_u1_n96, u0_u15_u1_n97, u0_u15_u1_n98, u0_u15_u1_n99, u0_u15_u2_n100, u0_u15_u2_n101, u0_u15_u2_n102, 
       u0_u15_u2_n103, u0_u15_u2_n104, u0_u15_u2_n105, u0_u15_u2_n106, u0_u15_u2_n107, u0_u15_u2_n108, u0_u15_u2_n109, u0_u15_u2_n110, u0_u15_u2_n111, 
       u0_u15_u2_n112, u0_u15_u2_n113, u0_u15_u2_n114, u0_u15_u2_n115, u0_u15_u2_n116, u0_u15_u2_n117, u0_u15_u2_n118, u0_u15_u2_n119, u0_u15_u2_n120, 
       u0_u15_u2_n121, u0_u15_u2_n122, u0_u15_u2_n123, u0_u15_u2_n124, u0_u15_u2_n125, u0_u15_u2_n126, u0_u15_u2_n127, u0_u15_u2_n128, u0_u15_u2_n129, 
       u0_u15_u2_n130, u0_u15_u2_n131, u0_u15_u2_n132, u0_u15_u2_n133, u0_u15_u2_n134, u0_u15_u2_n135, u0_u15_u2_n136, u0_u15_u2_n137, u0_u15_u2_n138, 
       u0_u15_u2_n139, u0_u15_u2_n140, u0_u15_u2_n141, u0_u15_u2_n142, u0_u15_u2_n143, u0_u15_u2_n144, u0_u15_u2_n145, u0_u15_u2_n146, u0_u15_u2_n147, 
       u0_u15_u2_n148, u0_u15_u2_n149, u0_u15_u2_n150, u0_u15_u2_n151, u0_u15_u2_n152, u0_u15_u2_n153, u0_u15_u2_n154, u0_u15_u2_n155, u0_u15_u2_n156, 
       u0_u15_u2_n157, u0_u15_u2_n158, u0_u15_u2_n159, u0_u15_u2_n160, u0_u15_u2_n161, u0_u15_u2_n162, u0_u15_u2_n163, u0_u15_u2_n164, u0_u15_u2_n165, 
       u0_u15_u2_n166, u0_u15_u2_n167, u0_u15_u2_n168, u0_u15_u2_n169, u0_u15_u2_n170, u0_u15_u2_n171, u0_u15_u2_n172, u0_u15_u2_n173, u0_u15_u2_n174, 
       u0_u15_u2_n175, u0_u15_u2_n176, u0_u15_u2_n177, u0_u15_u2_n178, u0_u15_u2_n179, u0_u15_u2_n180, u0_u15_u2_n181, u0_u15_u2_n182, u0_u15_u2_n183, 
       u0_u15_u2_n184, u0_u15_u2_n185, u0_u15_u2_n186, u0_u15_u2_n187, u0_u15_u2_n188, u0_u15_u2_n95, u0_u15_u2_n96, u0_u15_u2_n97, u0_u15_u2_n98, 
       u0_u15_u2_n99, u0_u15_u3_n100, u0_u15_u3_n101, u0_u15_u3_n102, u0_u15_u3_n103, u0_u15_u3_n104, u0_u15_u3_n105, u0_u15_u3_n106, u0_u15_u3_n107, 
       u0_u15_u3_n108, u0_u15_u3_n109, u0_u15_u3_n110, u0_u15_u3_n111, u0_u15_u3_n112, u0_u15_u3_n113, u0_u15_u3_n114, u0_u15_u3_n115, u0_u15_u3_n116, 
       u0_u15_u3_n117, u0_u15_u3_n118, u0_u15_u3_n119, u0_u15_u3_n120, u0_u15_u3_n121, u0_u15_u3_n122, u0_u15_u3_n123, u0_u15_u3_n124, u0_u15_u3_n125, 
       u0_u15_u3_n126, u0_u15_u3_n127, u0_u15_u3_n128, u0_u15_u3_n129, u0_u15_u3_n130, u0_u15_u3_n131, u0_u15_u3_n132, u0_u15_u3_n133, u0_u15_u3_n134, 
       u0_u15_u3_n135, u0_u15_u3_n136, u0_u15_u3_n137, u0_u15_u3_n138, u0_u15_u3_n139, u0_u15_u3_n140, u0_u15_u3_n141, u0_u15_u3_n142, u0_u15_u3_n143, 
       u0_u15_u3_n144, u0_u15_u3_n145, u0_u15_u3_n146, u0_u15_u3_n147, u0_u15_u3_n148, u0_u15_u3_n149, u0_u15_u3_n150, u0_u15_u3_n151, u0_u15_u3_n152, 
       u0_u15_u3_n153, u0_u15_u3_n154, u0_u15_u3_n155, u0_u15_u3_n156, u0_u15_u3_n157, u0_u15_u3_n158, u0_u15_u3_n159, u0_u15_u3_n160, u0_u15_u3_n161, 
       u0_u15_u3_n162, u0_u15_u3_n163, u0_u15_u3_n164, u0_u15_u3_n165, u0_u15_u3_n166, u0_u15_u3_n167, u0_u15_u3_n168, u0_u15_u3_n169, u0_u15_u3_n170, 
       u0_u15_u3_n171, u0_u15_u3_n172, u0_u15_u3_n173, u0_u15_u3_n174, u0_u15_u3_n175, u0_u15_u3_n176, u0_u15_u3_n177, u0_u15_u3_n178, u0_u15_u3_n179, 
       u0_u15_u3_n180, u0_u15_u3_n181, u0_u15_u3_n182, u0_u15_u3_n183, u0_u15_u3_n184, u0_u15_u3_n185, u0_u15_u3_n186, u0_u15_u3_n94, u0_u15_u3_n95, 
       u0_u15_u3_n96, u0_u15_u3_n97, u0_u15_u3_n98, u0_u15_u3_n99, u0_u1_X_5, u0_u1_X_6, u0_u1_X_7, u0_u1_X_8, u0_u1_u0_n100, 
       u0_u1_u0_n101, u0_u1_u0_n102, u0_u1_u0_n103, u0_u1_u0_n104, u0_u1_u0_n105, u0_u1_u0_n106, u0_u1_u0_n107, u0_u1_u0_n108, u0_u1_u0_n109, 
       u0_u1_u0_n110, u0_u1_u0_n111, u0_u1_u0_n112, u0_u1_u0_n113, u0_u1_u0_n114, u0_u1_u0_n115, u0_u1_u0_n116, u0_u1_u0_n117, u0_u1_u0_n118, 
       u0_u1_u0_n119, u0_u1_u0_n120, u0_u1_u0_n121, u0_u1_u0_n122, u0_u1_u0_n123, u0_u1_u0_n124, u0_u1_u0_n125, u0_u1_u0_n126, u0_u1_u0_n127, 
       u0_u1_u0_n128, u0_u1_u0_n129, u0_u1_u0_n130, u0_u1_u0_n131, u0_u1_u0_n132, u0_u1_u0_n133, u0_u1_u0_n134, u0_u1_u0_n135, u0_u1_u0_n136, 
       u0_u1_u0_n137, u0_u1_u0_n138, u0_u1_u0_n139, u0_u1_u0_n140, u0_u1_u0_n141, u0_u1_u0_n142, u0_u1_u0_n143, u0_u1_u0_n144, u0_u1_u0_n145, 
       u0_u1_u0_n146, u0_u1_u0_n147, u0_u1_u0_n148, u0_u1_u0_n149, u0_u1_u0_n150, u0_u1_u0_n151, u0_u1_u0_n152, u0_u1_u0_n153, u0_u1_u0_n154, 
       u0_u1_u0_n155, u0_u1_u0_n156, u0_u1_u0_n157, u0_u1_u0_n158, u0_u1_u0_n159, u0_u1_u0_n160, u0_u1_u0_n161, u0_u1_u0_n162, u0_u1_u0_n163, 
       u0_u1_u0_n164, u0_u1_u0_n165, u0_u1_u0_n166, u0_u1_u0_n167, u0_u1_u0_n168, u0_u1_u0_n169, u0_u1_u0_n170, u0_u1_u0_n171, u0_u1_u0_n172, 
       u0_u1_u0_n173, u0_u1_u0_n174, u0_u1_u0_n88, u0_u1_u0_n89, u0_u1_u0_n90, u0_u1_u0_n91, u0_u1_u0_n92, u0_u1_u0_n93, u0_u1_u0_n94, 
       u0_u1_u0_n95, u0_u1_u0_n96, u0_u1_u0_n97, u0_u1_u0_n98, u0_u1_u0_n99, u0_u1_u1_n100, u0_u1_u1_n101, u0_u1_u1_n102, u0_u1_u1_n103, 
       u0_u1_u1_n104, u0_u1_u1_n105, u0_u1_u1_n106, u0_u1_u1_n107, u0_u1_u1_n108, u0_u1_u1_n109, u0_u1_u1_n110, u0_u1_u1_n111, u0_u1_u1_n112, 
       u0_u1_u1_n113, u0_u1_u1_n114, u0_u1_u1_n115, u0_u1_u1_n116, u0_u1_u1_n117, u0_u1_u1_n118, u0_u1_u1_n119, u0_u1_u1_n120, u0_u1_u1_n121, 
       u0_u1_u1_n122, u0_u1_u1_n123, u0_u1_u1_n124, u0_u1_u1_n125, u0_u1_u1_n126, u0_u1_u1_n127, u0_u1_u1_n128, u0_u1_u1_n129, u0_u1_u1_n130, 
       u0_u1_u1_n131, u0_u1_u1_n132, u0_u1_u1_n133, u0_u1_u1_n134, u0_u1_u1_n135, u0_u1_u1_n136, u0_u1_u1_n137, u0_u1_u1_n138, u0_u1_u1_n139, 
       u0_u1_u1_n140, u0_u1_u1_n141, u0_u1_u1_n142, u0_u1_u1_n143, u0_u1_u1_n144, u0_u1_u1_n145, u0_u1_u1_n146, u0_u1_u1_n147, u0_u1_u1_n148, 
       u0_u1_u1_n149, u0_u1_u1_n150, u0_u1_u1_n151, u0_u1_u1_n152, u0_u1_u1_n153, u0_u1_u1_n154, u0_u1_u1_n155, u0_u1_u1_n156, u0_u1_u1_n157, 
       u0_u1_u1_n158, u0_u1_u1_n159, u0_u1_u1_n160, u0_u1_u1_n161, u0_u1_u1_n162, u0_u1_u1_n163, u0_u1_u1_n164, u0_u1_u1_n165, u0_u1_u1_n166, 
       u0_u1_u1_n167, u0_u1_u1_n168, u0_u1_u1_n169, u0_u1_u1_n170, u0_u1_u1_n171, u0_u1_u1_n172, u0_u1_u1_n173, u0_u1_u1_n174, u0_u1_u1_n175, 
       u0_u1_u1_n176, u0_u1_u1_n177, u0_u1_u1_n178, u0_u1_u1_n179, u0_u1_u1_n180, u0_u1_u1_n181, u0_u1_u1_n182, u0_u1_u1_n183, u0_u1_u1_n184, 
       u0_u1_u1_n185, u0_u1_u1_n186, u0_u1_u1_n187, u0_u1_u1_n188, u0_u1_u1_n95, u0_u1_u1_n96, u0_u1_u1_n97, u0_u1_u1_n98, u0_u1_u1_n99, 
       u0_u3_X_1, u0_u3_X_10, u0_u3_X_11, u0_u3_X_12, u0_u3_X_13, u0_u3_X_14, u0_u3_X_15, u0_u3_X_16, u0_u3_X_17, 
       u0_u3_X_18, u0_u3_X_2, u0_u3_X_4, u0_u3_X_5, u0_u3_X_7, u0_u3_X_9, u0_u3_u0_n100, u0_u3_u0_n101, u0_u3_u0_n102, 
       u0_u3_u0_n103, u0_u3_u0_n104, u0_u3_u0_n105, u0_u3_u0_n106, u0_u3_u0_n107, u0_u3_u0_n108, u0_u3_u0_n109, u0_u3_u0_n110, u0_u3_u0_n111, 
       u0_u3_u0_n112, u0_u3_u0_n113, u0_u3_u0_n114, u0_u3_u0_n115, u0_u3_u0_n116, u0_u3_u0_n117, u0_u3_u0_n118, u0_u3_u0_n119, u0_u3_u0_n120, 
       u0_u3_u0_n121, u0_u3_u0_n122, u0_u3_u0_n123, u0_u3_u0_n124, u0_u3_u0_n125, u0_u3_u0_n126, u0_u3_u0_n127, u0_u3_u0_n128, u0_u3_u0_n129, 
       u0_u3_u0_n130, u0_u3_u0_n131, u0_u3_u0_n132, u0_u3_u0_n133, u0_u3_u0_n134, u0_u3_u0_n135, u0_u3_u0_n136, u0_u3_u0_n137, u0_u3_u0_n138, 
       u0_u3_u0_n139, u0_u3_u0_n140, u0_u3_u0_n141, u0_u3_u0_n142, u0_u3_u0_n143, u0_u3_u0_n144, u0_u3_u0_n145, u0_u3_u0_n146, u0_u3_u0_n147, 
       u0_u3_u0_n148, u0_u3_u0_n149, u0_u3_u0_n150, u0_u3_u0_n151, u0_u3_u0_n152, u0_u3_u0_n153, u0_u3_u0_n154, u0_u3_u0_n155, u0_u3_u0_n156, 
       u0_u3_u0_n157, u0_u3_u0_n158, u0_u3_u0_n159, u0_u3_u0_n160, u0_u3_u0_n161, u0_u3_u0_n162, u0_u3_u0_n163, u0_u3_u0_n164, u0_u3_u0_n165, 
       u0_u3_u0_n166, u0_u3_u0_n167, u0_u3_u0_n168, u0_u3_u0_n169, u0_u3_u0_n170, u0_u3_u0_n171, u0_u3_u0_n172, u0_u3_u0_n173, u0_u3_u0_n174, 
       u0_u3_u0_n175, u0_u3_u0_n176, u0_u3_u0_n88, u0_u3_u0_n89, u0_u3_u0_n90, u0_u3_u0_n91, u0_u3_u0_n92, u0_u3_u0_n93, u0_u3_u0_n94, 
       u0_u3_u0_n95, u0_u3_u0_n96, u0_u3_u0_n97, u0_u3_u0_n98, u0_u3_u0_n99, u0_u3_u1_n100, u0_u3_u1_n101, u0_u3_u1_n102, u0_u3_u1_n103, 
       u0_u3_u1_n104, u0_u3_u1_n105, u0_u3_u1_n106, u0_u3_u1_n107, u0_u3_u1_n108, u0_u3_u1_n109, u0_u3_u1_n110, u0_u3_u1_n111, u0_u3_u1_n112, 
       u0_u3_u1_n113, u0_u3_u1_n114, u0_u3_u1_n115, u0_u3_u1_n116, u0_u3_u1_n117, u0_u3_u1_n118, u0_u3_u1_n119, u0_u3_u1_n120, u0_u3_u1_n121, 
       u0_u3_u1_n122, u0_u3_u1_n123, u0_u3_u1_n124, u0_u3_u1_n125, u0_u3_u1_n126, u0_u3_u1_n127, u0_u3_u1_n128, u0_u3_u1_n129, u0_u3_u1_n130, 
       u0_u3_u1_n131, u0_u3_u1_n132, u0_u3_u1_n133, u0_u3_u1_n134, u0_u3_u1_n135, u0_u3_u1_n136, u0_u3_u1_n137, u0_u3_u1_n138, u0_u3_u1_n139, 
       u0_u3_u1_n140, u0_u3_u1_n141, u0_u3_u1_n142, u0_u3_u1_n143, u0_u3_u1_n144, u0_u3_u1_n145, u0_u3_u1_n146, u0_u3_u1_n147, u0_u3_u1_n148, 
       u0_u3_u1_n149, u0_u3_u1_n150, u0_u3_u1_n151, u0_u3_u1_n152, u0_u3_u1_n153, u0_u3_u1_n154, u0_u3_u1_n155, u0_u3_u1_n156, u0_u3_u1_n157, 
       u0_u3_u1_n158, u0_u3_u1_n159, u0_u3_u1_n160, u0_u3_u1_n161, u0_u3_u1_n162, u0_u3_u1_n163, u0_u3_u1_n164, u0_u3_u1_n165, u0_u3_u1_n166, 
       u0_u3_u1_n167, u0_u3_u1_n168, u0_u3_u1_n169, u0_u3_u1_n170, u0_u3_u1_n171, u0_u3_u1_n172, u0_u3_u1_n173, u0_u3_u1_n174, u0_u3_u1_n175, 
       u0_u3_u1_n176, u0_u3_u1_n177, u0_u3_u1_n178, u0_u3_u1_n179, u0_u3_u1_n180, u0_u3_u1_n181, u0_u3_u1_n182, u0_u3_u1_n183, u0_u3_u1_n184, 
       u0_u3_u1_n185, u0_u3_u1_n186, u0_u3_u1_n187, u0_u3_u1_n188, u0_u3_u1_n95, u0_u3_u1_n96, u0_u3_u1_n97, u0_u3_u1_n98, u0_u3_u1_n99, 
       u0_u3_u2_n100, u0_u3_u2_n101, u0_u3_u2_n102, u0_u3_u2_n103, u0_u3_u2_n104, u0_u3_u2_n105, u0_u3_u2_n106, u0_u3_u2_n107, u0_u3_u2_n108, 
       u0_u3_u2_n109, u0_u3_u2_n110, u0_u3_u2_n111, u0_u3_u2_n112, u0_u3_u2_n113, u0_u3_u2_n114, u0_u3_u2_n115, u0_u3_u2_n116, u0_u3_u2_n117, 
       u0_u3_u2_n118, u0_u3_u2_n119, u0_u3_u2_n120, u0_u3_u2_n121, u0_u3_u2_n122, u0_u3_u2_n123, u0_u3_u2_n124, u0_u3_u2_n125, u0_u3_u2_n126, 
       u0_u3_u2_n127, u0_u3_u2_n128, u0_u3_u2_n129, u0_u3_u2_n130, u0_u3_u2_n131, u0_u3_u2_n132, u0_u3_u2_n133, u0_u3_u2_n134, u0_u3_u2_n135, 
       u0_u3_u2_n136, u0_u3_u2_n137, u0_u3_u2_n138, u0_u3_u2_n139, u0_u3_u2_n140, u0_u3_u2_n141, u0_u3_u2_n142, u0_u3_u2_n143, u0_u3_u2_n144, 
       u0_u3_u2_n145, u0_u3_u2_n146, u0_u3_u2_n147, u0_u3_u2_n148, u0_u3_u2_n149, u0_u3_u2_n150, u0_u3_u2_n151, u0_u3_u2_n152, u0_u3_u2_n153, 
       u0_u3_u2_n154, u0_u3_u2_n155, u0_u3_u2_n156, u0_u3_u2_n157, u0_u3_u2_n158, u0_u3_u2_n159, u0_u3_u2_n160, u0_u3_u2_n161, u0_u3_u2_n162, 
       u0_u3_u2_n163, u0_u3_u2_n164, u0_u3_u2_n165, u0_u3_u2_n166, u0_u3_u2_n167, u0_u3_u2_n168, u0_u3_u2_n169, u0_u3_u2_n170, u0_u3_u2_n171, 
       u0_u3_u2_n172, u0_u3_u2_n173, u0_u3_u2_n174, u0_u3_u2_n175, u0_u3_u2_n176, u0_u3_u2_n177, u0_u3_u2_n178, u0_u3_u2_n179, u0_u3_u2_n180, 
       u0_u3_u2_n181, u0_u3_u2_n182, u0_u3_u2_n183, u0_u3_u2_n184, u0_u3_u2_n185, u0_u3_u2_n186, u0_u3_u2_n187, u0_u3_u2_n188, u0_u3_u2_n95, 
       u0_u3_u2_n96, u0_u3_u2_n97, u0_u3_u2_n98, u0_u3_u2_n99, u0_u5_X_11, u0_u5_X_13, u0_u5_X_18, u0_u5_X_20, u0_u5_X_21, 
       u0_u5_X_23, u0_u5_X_25, u0_u5_u1_n100, u0_u5_u1_n101, u0_u5_u1_n102, u0_u5_u1_n103, u0_u5_u1_n104, u0_u5_u1_n105, u0_u5_u1_n106, 
       u0_u5_u1_n107, u0_u5_u1_n108, u0_u5_u1_n109, u0_u5_u1_n110, u0_u5_u1_n111, u0_u5_u1_n112, u0_u5_u1_n113, u0_u5_u1_n114, u0_u5_u1_n115, 
       u0_u5_u1_n116, u0_u5_u1_n117, u0_u5_u1_n118, u0_u5_u1_n119, u0_u5_u1_n120, u0_u5_u1_n121, u0_u5_u1_n122, u0_u5_u1_n123, u0_u5_u1_n124, 
       u0_u5_u1_n125, u0_u5_u1_n126, u0_u5_u1_n127, u0_u5_u1_n128, u0_u5_u1_n129, u0_u5_u1_n130, u0_u5_u1_n131, u0_u5_u1_n132, u0_u5_u1_n133, 
       u0_u5_u1_n134, u0_u5_u1_n135, u0_u5_u1_n136, u0_u5_u1_n137, u0_u5_u1_n138, u0_u5_u1_n139, u0_u5_u1_n140, u0_u5_u1_n141, u0_u5_u1_n142, 
       u0_u5_u1_n143, u0_u5_u1_n144, u0_u5_u1_n145, u0_u5_u1_n146, u0_u5_u1_n147, u0_u5_u1_n148, u0_u5_u1_n149, u0_u5_u1_n150, u0_u5_u1_n151, 
       u0_u5_u1_n152, u0_u5_u1_n153, u0_u5_u1_n154, u0_u5_u1_n155, u0_u5_u1_n156, u0_u5_u1_n157, u0_u5_u1_n158, u0_u5_u1_n159, u0_u5_u1_n160, 
       u0_u5_u1_n161, u0_u5_u1_n162, u0_u5_u1_n163, u0_u5_u1_n164, u0_u5_u1_n165, u0_u5_u1_n166, u0_u5_u1_n167, u0_u5_u1_n168, u0_u5_u1_n169, 
       u0_u5_u1_n170, u0_u5_u1_n171, u0_u5_u1_n172, u0_u5_u1_n173, u0_u5_u1_n174, u0_u5_u1_n175, u0_u5_u1_n176, u0_u5_u1_n177, u0_u5_u1_n178, 
       u0_u5_u1_n179, u0_u5_u1_n180, u0_u5_u1_n181, u0_u5_u1_n182, u0_u5_u1_n183, u0_u5_u1_n184, u0_u5_u1_n185, u0_u5_u1_n186, u0_u5_u1_n187, 
       u0_u5_u1_n188, u0_u5_u1_n95, u0_u5_u1_n96, u0_u5_u1_n97, u0_u5_u1_n98, u0_u5_u1_n99, u0_u5_u2_n100, u0_u5_u2_n101, u0_u5_u2_n102, 
       u0_u5_u2_n103, u0_u5_u2_n104, u0_u5_u2_n105, u0_u5_u2_n106, u0_u5_u2_n107, u0_u5_u2_n108, u0_u5_u2_n109, u0_u5_u2_n110, u0_u5_u2_n111, 
       u0_u5_u2_n112, u0_u5_u2_n113, u0_u5_u2_n114, u0_u5_u2_n115, u0_u5_u2_n116, u0_u5_u2_n117, u0_u5_u2_n118, u0_u5_u2_n119, u0_u5_u2_n120, 
       u0_u5_u2_n121, u0_u5_u2_n122, u0_u5_u2_n123, u0_u5_u2_n124, u0_u5_u2_n125, u0_u5_u2_n126, u0_u5_u2_n127, u0_u5_u2_n128, u0_u5_u2_n129, 
       u0_u5_u2_n130, u0_u5_u2_n131, u0_u5_u2_n132, u0_u5_u2_n133, u0_u5_u2_n134, u0_u5_u2_n135, u0_u5_u2_n136, u0_u5_u2_n137, u0_u5_u2_n138, 
       u0_u5_u2_n139, u0_u5_u2_n140, u0_u5_u2_n141, u0_u5_u2_n142, u0_u5_u2_n143, u0_u5_u2_n144, u0_u5_u2_n145, u0_u5_u2_n146, u0_u5_u2_n147, 
       u0_u5_u2_n148, u0_u5_u2_n149, u0_u5_u2_n150, u0_u5_u2_n151, u0_u5_u2_n152, u0_u5_u2_n153, u0_u5_u2_n154, u0_u5_u2_n155, u0_u5_u2_n156, 
       u0_u5_u2_n157, u0_u5_u2_n158, u0_u5_u2_n159, u0_u5_u2_n160, u0_u5_u2_n161, u0_u5_u2_n162, u0_u5_u2_n163, u0_u5_u2_n164, u0_u5_u2_n165, 
       u0_u5_u2_n166, u0_u5_u2_n167, u0_u5_u2_n168, u0_u5_u2_n169, u0_u5_u2_n170, u0_u5_u2_n171, u0_u5_u2_n172, u0_u5_u2_n173, u0_u5_u2_n174, 
       u0_u5_u2_n175, u0_u5_u2_n176, u0_u5_u2_n177, u0_u5_u2_n178, u0_u5_u2_n179, u0_u5_u2_n180, u0_u5_u2_n181, u0_u5_u2_n182, u0_u5_u2_n183, 
       u0_u5_u2_n184, u0_u5_u2_n185, u0_u5_u2_n186, u0_u5_u2_n187, u0_u5_u2_n188, u0_u5_u2_n95, u0_u5_u2_n96, u0_u5_u2_n97, u0_u5_u2_n98, 
       u0_u5_u2_n99, u0_u5_u3_n100, u0_u5_u3_n101, u0_u5_u3_n102, u0_u5_u3_n103, u0_u5_u3_n104, u0_u5_u3_n105, u0_u5_u3_n106, u0_u5_u3_n107, 
       u0_u5_u3_n108, u0_u5_u3_n109, u0_u5_u3_n110, u0_u5_u3_n111, u0_u5_u3_n112, u0_u5_u3_n113, u0_u5_u3_n114, u0_u5_u3_n115, u0_u5_u3_n116, 
       u0_u5_u3_n117, u0_u5_u3_n118, u0_u5_u3_n119, u0_u5_u3_n120, u0_u5_u3_n121, u0_u5_u3_n122, u0_u5_u3_n123, u0_u5_u3_n124, u0_u5_u3_n125, 
       u0_u5_u3_n126, u0_u5_u3_n127, u0_u5_u3_n128, u0_u5_u3_n129, u0_u5_u3_n130, u0_u5_u3_n131, u0_u5_u3_n132, u0_u5_u3_n133, u0_u5_u3_n134, 
       u0_u5_u3_n135, u0_u5_u3_n136, u0_u5_u3_n137, u0_u5_u3_n138, u0_u5_u3_n139, u0_u5_u3_n140, u0_u5_u3_n141, u0_u5_u3_n142, u0_u5_u3_n143, 
       u0_u5_u3_n144, u0_u5_u3_n145, u0_u5_u3_n146, u0_u5_u3_n147, u0_u5_u3_n148, u0_u5_u3_n149, u0_u5_u3_n150, u0_u5_u3_n151, u0_u5_u3_n152, 
       u0_u5_u3_n153, u0_u5_u3_n154, u0_u5_u3_n155, u0_u5_u3_n156, u0_u5_u3_n157, u0_u5_u3_n158, u0_u5_u3_n159, u0_u5_u3_n160, u0_u5_u3_n161, 
       u0_u5_u3_n162, u0_u5_u3_n163, u0_u5_u3_n164, u0_u5_u3_n165, u0_u5_u3_n166, u0_u5_u3_n167, u0_u5_u3_n168, u0_u5_u3_n169, u0_u5_u3_n170, 
       u0_u5_u3_n171, u0_u5_u3_n172, u0_u5_u3_n173, u0_u5_u3_n174, u0_u5_u3_n175, u0_u5_u3_n176, u0_u5_u3_n177, u0_u5_u3_n178, u0_u5_u3_n179, 
       u0_u5_u3_n180, u0_u5_u3_n181, u0_u5_u3_n182, u0_u5_u3_n183, u0_u5_u3_n184, u0_u5_u3_n185, u0_u5_u3_n186, u0_u5_u3_n94, u0_u5_u3_n95, 
       u0_u5_u3_n96, u0_u5_u3_n97, u0_u5_u3_n98, u0_u5_u3_n99, u0_u5_u4_n100, u0_u5_u4_n101, u0_u5_u4_n102, u0_u5_u4_n103, u0_u5_u4_n104, 
       u0_u5_u4_n105, u0_u5_u4_n106, u0_u5_u4_n107, u0_u5_u4_n108, u0_u5_u4_n109, u0_u5_u4_n110, u0_u5_u4_n111, u0_u5_u4_n112, u0_u5_u4_n113, 
       u0_u5_u4_n114, u0_u5_u4_n115, u0_u5_u4_n116, u0_u5_u4_n117, u0_u5_u4_n118, u0_u5_u4_n119, u0_u5_u4_n120, u0_u5_u4_n121, u0_u5_u4_n122, 
       u0_u5_u4_n123, u0_u5_u4_n124, u0_u5_u4_n125, u0_u5_u4_n126, u0_u5_u4_n127, u0_u5_u4_n128, u0_u5_u4_n129, u0_u5_u4_n130, u0_u5_u4_n131, 
       u0_u5_u4_n132, u0_u5_u4_n133, u0_u5_u4_n134, u0_u5_u4_n135, u0_u5_u4_n136, u0_u5_u4_n137, u0_u5_u4_n138, u0_u5_u4_n139, u0_u5_u4_n140, 
       u0_u5_u4_n141, u0_u5_u4_n142, u0_u5_u4_n143, u0_u5_u4_n144, u0_u5_u4_n145, u0_u5_u4_n146, u0_u5_u4_n147, u0_u5_u4_n148, u0_u5_u4_n149, 
       u0_u5_u4_n150, u0_u5_u4_n151, u0_u5_u4_n152, u0_u5_u4_n153, u0_u5_u4_n154, u0_u5_u4_n155, u0_u5_u4_n156, u0_u5_u4_n157, u0_u5_u4_n158, 
       u0_u5_u4_n159, u0_u5_u4_n160, u0_u5_u4_n161, u0_u5_u4_n162, u0_u5_u4_n163, u0_u5_u4_n164, u0_u5_u4_n165, u0_u5_u4_n166, u0_u5_u4_n167, 
       u0_u5_u4_n168, u0_u5_u4_n169, u0_u5_u4_n170, u0_u5_u4_n171, u0_u5_u4_n172, u0_u5_u4_n173, u0_u5_u4_n174, u0_u5_u4_n175, u0_u5_u4_n176, 
       u0_u5_u4_n177, u0_u5_u4_n178, u0_u5_u4_n179, u0_u5_u4_n180, u0_u5_u4_n181, u0_u5_u4_n182, u0_u5_u4_n183, u0_u5_u4_n184, u0_u5_u4_n185, 
       u0_u5_u4_n186, u0_u5_u4_n94, u0_u5_u4_n95, u0_u5_u4_n96, u0_u5_u4_n97, u0_u5_u4_n98, u0_u5_u4_n99, u0_u7_X_19, u0_u7_X_20, 
       u0_u7_X_21, u0_u7_X_23, u0_u7_X_24, u0_u7_X_25, u0_u7_X_26, u0_u7_X_27, u0_u7_X_29, u0_u7_X_30, u0_u7_X_31, 
       u0_u7_X_32, u0_u7_X_34, u0_u7_X_35, u0_u7_X_43, u0_u7_X_44, u0_u7_X_47, u0_u7_X_48, u0_u7_u3_n100, u0_u7_u3_n101, 
       u0_u7_u3_n102, u0_u7_u3_n103, u0_u7_u3_n104, u0_u7_u3_n105, u0_u7_u3_n106, u0_u7_u3_n107, u0_u7_u3_n108, u0_u7_u3_n109, u0_u7_u3_n110, 
       u0_u7_u3_n111, u0_u7_u3_n112, u0_u7_u3_n113, u0_u7_u3_n114, u0_u7_u3_n115, u0_u7_u3_n116, u0_u7_u3_n117, u0_u7_u3_n118, u0_u7_u3_n119, 
       u0_u7_u3_n120, u0_u7_u3_n121, u0_u7_u3_n122, u0_u7_u3_n123, u0_u7_u3_n124, u0_u7_u3_n125, u0_u7_u3_n126, u0_u7_u3_n127, u0_u7_u3_n128, 
       u0_u7_u3_n129, u0_u7_u3_n130, u0_u7_u3_n131, u0_u7_u3_n132, u0_u7_u3_n133, u0_u7_u3_n134, u0_u7_u3_n135, u0_u7_u3_n136, u0_u7_u3_n137, 
       u0_u7_u3_n138, u0_u7_u3_n139, u0_u7_u3_n140, u0_u7_u3_n141, u0_u7_u3_n142, u0_u7_u3_n143, u0_u7_u3_n144, u0_u7_u3_n145, u0_u7_u3_n146, 
       u0_u7_u3_n147, u0_u7_u3_n148, u0_u7_u3_n149, u0_u7_u3_n150, u0_u7_u3_n151, u0_u7_u3_n152, u0_u7_u3_n153, u0_u7_u3_n154, u0_u7_u3_n155, 
       u0_u7_u3_n156, u0_u7_u3_n157, u0_u7_u3_n158, u0_u7_u3_n159, u0_u7_u3_n160, u0_u7_u3_n161, u0_u7_u3_n162, u0_u7_u3_n163, u0_u7_u3_n164, 
       u0_u7_u3_n165, u0_u7_u3_n166, u0_u7_u3_n167, u0_u7_u3_n168, u0_u7_u3_n169, u0_u7_u3_n170, u0_u7_u3_n171, u0_u7_u3_n172, u0_u7_u3_n173, 
       u0_u7_u3_n174, u0_u7_u3_n175, u0_u7_u3_n176, u0_u7_u3_n177, u0_u7_u3_n178, u0_u7_u3_n179, u0_u7_u3_n180, u0_u7_u3_n181, u0_u7_u3_n182, 
       u0_u7_u3_n183, u0_u7_u3_n184, u0_u7_u3_n185, u0_u7_u3_n186, u0_u7_u3_n94, u0_u7_u3_n95, u0_u7_u3_n96, u0_u7_u3_n97, u0_u7_u3_n98, 
       u0_u7_u3_n99, u0_u7_u4_n100, u0_u7_u4_n101, u0_u7_u4_n102, u0_u7_u4_n103, u0_u7_u4_n104, u0_u7_u4_n105, u0_u7_u4_n106, u0_u7_u4_n107, 
       u0_u7_u4_n108, u0_u7_u4_n109, u0_u7_u4_n110, u0_u7_u4_n111, u0_u7_u4_n112, u0_u7_u4_n113, u0_u7_u4_n114, u0_u7_u4_n115, u0_u7_u4_n116, 
       u0_u7_u4_n117, u0_u7_u4_n118, u0_u7_u4_n119, u0_u7_u4_n120, u0_u7_u4_n121, u0_u7_u4_n122, u0_u7_u4_n123, u0_u7_u4_n124, u0_u7_u4_n125, 
       u0_u7_u4_n126, u0_u7_u4_n127, u0_u7_u4_n128, u0_u7_u4_n129, u0_u7_u4_n130, u0_u7_u4_n131, u0_u7_u4_n132, u0_u7_u4_n133, u0_u7_u4_n134, 
       u0_u7_u4_n135, u0_u7_u4_n136, u0_u7_u4_n137, u0_u7_u4_n138, u0_u7_u4_n139, u0_u7_u4_n140, u0_u7_u4_n141, u0_u7_u4_n142, u0_u7_u4_n143, 
       u0_u7_u4_n144, u0_u7_u4_n145, u0_u7_u4_n146, u0_u7_u4_n147, u0_u7_u4_n148, u0_u7_u4_n149, u0_u7_u4_n150, u0_u7_u4_n151, u0_u7_u4_n152, 
       u0_u7_u4_n153, u0_u7_u4_n154, u0_u7_u4_n155, u0_u7_u4_n156, u0_u7_u4_n157, u0_u7_u4_n158, u0_u7_u4_n159, u0_u7_u4_n160, u0_u7_u4_n161, 
       u0_u7_u4_n162, u0_u7_u4_n163, u0_u7_u4_n164, u0_u7_u4_n165, u0_u7_u4_n166, u0_u7_u4_n167, u0_u7_u4_n168, u0_u7_u4_n169, u0_u7_u4_n170, 
       u0_u7_u4_n171, u0_u7_u4_n172, u0_u7_u4_n173, u0_u7_u4_n174, u0_u7_u4_n175, u0_u7_u4_n176, u0_u7_u4_n177, u0_u7_u4_n178, u0_u7_u4_n179, 
       u0_u7_u4_n180, u0_u7_u4_n181, u0_u7_u4_n182, u0_u7_u4_n183, u0_u7_u4_n184, u0_u7_u4_n185, u0_u7_u4_n186, u0_u7_u4_n94, u0_u7_u4_n95, 
       u0_u7_u4_n96, u0_u7_u4_n97, u0_u7_u4_n98, u0_u7_u4_n99, u0_u7_u5_n100, u0_u7_u5_n101, u0_u7_u5_n102, u0_u7_u5_n103, u0_u7_u5_n104, 
       u0_u7_u5_n105, u0_u7_u5_n106, u0_u7_u5_n107, u0_u7_u5_n108, u0_u7_u5_n109, u0_u7_u5_n110, u0_u7_u5_n111, u0_u7_u5_n112, u0_u7_u5_n113, 
       u0_u7_u5_n114, u0_u7_u5_n115, u0_u7_u5_n116, u0_u7_u5_n117, u0_u7_u5_n118, u0_u7_u5_n119, u0_u7_u5_n120, u0_u7_u5_n121, u0_u7_u5_n122, 
       u0_u7_u5_n123, u0_u7_u5_n124, u0_u7_u5_n125, u0_u7_u5_n126, u0_u7_u5_n127, u0_u7_u5_n128, u0_u7_u5_n129, u0_u7_u5_n130, u0_u7_u5_n131, 
       u0_u7_u5_n132, u0_u7_u5_n133, u0_u7_u5_n134, u0_u7_u5_n135, u0_u7_u5_n136, u0_u7_u5_n137, u0_u7_u5_n138, u0_u7_u5_n139, u0_u7_u5_n140, 
       u0_u7_u5_n141, u0_u7_u5_n142, u0_u7_u5_n143, u0_u7_u5_n144, u0_u7_u5_n145, u0_u7_u5_n146, u0_u7_u5_n147, u0_u7_u5_n148, u0_u7_u5_n149, 
       u0_u7_u5_n150, u0_u7_u5_n151, u0_u7_u5_n152, u0_u7_u5_n153, u0_u7_u5_n154, u0_u7_u5_n155, u0_u7_u5_n156, u0_u7_u5_n157, u0_u7_u5_n158, 
       u0_u7_u5_n159, u0_u7_u5_n160, u0_u7_u5_n161, u0_u7_u5_n162, u0_u7_u5_n163, u0_u7_u5_n164, u0_u7_u5_n165, u0_u7_u5_n166, u0_u7_u5_n167, 
       u0_u7_u5_n168, u0_u7_u5_n169, u0_u7_u5_n170, u0_u7_u5_n171, u0_u7_u5_n172, u0_u7_u5_n173, u0_u7_u5_n174, u0_u7_u5_n175, u0_u7_u5_n176, 
       u0_u7_u5_n177, u0_u7_u5_n178, u0_u7_u5_n179, u0_u7_u5_n180, u0_u7_u5_n181, u0_u7_u5_n182, u0_u7_u5_n183, u0_u7_u5_n184, u0_u7_u5_n185, 
       u0_u7_u5_n186, u0_u7_u5_n187, u0_u7_u5_n188, u0_u7_u5_n189, u0_u7_u5_n190, u0_u7_u5_n191, u0_u7_u5_n192, u0_u7_u5_n193, u0_u7_u5_n194, 
       u0_u7_u5_n195, u0_u7_u5_n196, u0_u7_u5_n99, u0_u7_u7_n100, u0_u7_u7_n101, u0_u7_u7_n102, u0_u7_u7_n103, u0_u7_u7_n104, u0_u7_u7_n105, 
       u0_u7_u7_n106, u0_u7_u7_n107, u0_u7_u7_n108, u0_u7_u7_n109, u0_u7_u7_n110, u0_u7_u7_n111, u0_u7_u7_n112, u0_u7_u7_n113, u0_u7_u7_n114, 
       u0_u7_u7_n115, u0_u7_u7_n116, u0_u7_u7_n117, u0_u7_u7_n118, u0_u7_u7_n119, u0_u7_u7_n120, u0_u7_u7_n121, u0_u7_u7_n122, u0_u7_u7_n123, 
       u0_u7_u7_n124, u0_u7_u7_n125, u0_u7_u7_n126, u0_u7_u7_n127, u0_u7_u7_n128, u0_u7_u7_n129, u0_u7_u7_n130, u0_u7_u7_n131, u0_u7_u7_n132, 
       u0_u7_u7_n133, u0_u7_u7_n134, u0_u7_u7_n135, u0_u7_u7_n136, u0_u7_u7_n137, u0_u7_u7_n138, u0_u7_u7_n139, u0_u7_u7_n140, u0_u7_u7_n141, 
       u0_u7_u7_n142, u0_u7_u7_n143, u0_u7_u7_n144, u0_u7_u7_n145, u0_u7_u7_n146, u0_u7_u7_n147, u0_u7_u7_n148, u0_u7_u7_n149, u0_u7_u7_n150, 
       u0_u7_u7_n151, u0_u7_u7_n152, u0_u7_u7_n153, u0_u7_u7_n154, u0_u7_u7_n155, u0_u7_u7_n156, u0_u7_u7_n157, u0_u7_u7_n158, u0_u7_u7_n159, 
       u0_u7_u7_n160, u0_u7_u7_n161, u0_u7_u7_n162, u0_u7_u7_n163, u0_u7_u7_n164, u0_u7_u7_n165, u0_u7_u7_n166, u0_u7_u7_n167, u0_u7_u7_n168, 
       u0_u7_u7_n169, u0_u7_u7_n170, u0_u7_u7_n171, u0_u7_u7_n172, u0_u7_u7_n173, u0_u7_u7_n174, u0_u7_u7_n175, u0_u7_u7_n176, u0_u7_u7_n177, 
       u0_u7_u7_n178, u0_u7_u7_n179, u0_u7_u7_n180, u0_u7_u7_n91, u0_u7_u7_n92, u0_u7_u7_n93, u0_u7_u7_n94, u0_u7_u7_n95, u0_u7_u7_n96, 
       u0_u7_u7_n97, u0_u7_u7_n98, u0_u7_u7_n99, u0_uk_n693, u0_uk_n700, u0_uk_n706, u0_uk_n709, u0_uk_n714, u0_uk_n745, 
       u0_uk_n752, u0_uk_n753, u0_uk_n821, u0_uk_n822, u0_uk_n836, u0_uk_n837, u0_uk_n838, u0_uk_n870, u0_uk_n872, 
       u0_uk_n873, u0_uk_n874, u0_uk_n876, u0_uk_n877, u0_uk_n882, u0_uk_n883, u0_uk_n903, u0_uk_n908, u0_uk_n909, 
       u0_uk_n910, u0_uk_n929, u0_uk_n930, u0_uk_n941, u0_uk_n943, u0_uk_n952, u0_uk_n958, u0_uk_n959, u0_uk_n996, 
       u0_uk_n997, u1_K10_22, u1_K11_12, u1_K11_14, u1_K11_8, u1_K12_15, u1_K12_3, u1_K12_4, u1_K13_21, 
       u1_K13_22, u1_K13_6, u1_K1_22, u1_K6_10, u1_K6_2, u1_K6_21, u1_K6_4, u1_K6_9, u1_K9_10, 
       u1_K9_11, u1_K9_9, u1_u0_X_21, u1_u0_X_22, u1_u0_X_3, u1_u0_X_4, u1_u0_u0_n100, u1_u0_u0_n101, u1_u0_u0_n102, 
       u1_u0_u0_n103, u1_u0_u0_n104, u1_u0_u0_n105, u1_u0_u0_n106, u1_u0_u0_n107, u1_u0_u0_n108, u1_u0_u0_n109, u1_u0_u0_n110, u1_u0_u0_n111, 
       u1_u0_u0_n112, u1_u0_u0_n113, u1_u0_u0_n114, u1_u0_u0_n115, u1_u0_u0_n116, u1_u0_u0_n117, u1_u0_u0_n118, u1_u0_u0_n119, u1_u0_u0_n120, 
       u1_u0_u0_n121, u1_u0_u0_n122, u1_u0_u0_n123, u1_u0_u0_n124, u1_u0_u0_n125, u1_u0_u0_n126, u1_u0_u0_n127, u1_u0_u0_n128, u1_u0_u0_n129, 
       u1_u0_u0_n130, u1_u0_u0_n131, u1_u0_u0_n132, u1_u0_u0_n133, u1_u0_u0_n134, u1_u0_u0_n135, u1_u0_u0_n136, u1_u0_u0_n137, u1_u0_u0_n138, 
       u1_u0_u0_n139, u1_u0_u0_n140, u1_u0_u0_n141, u1_u0_u0_n142, u1_u0_u0_n143, u1_u0_u0_n144, u1_u0_u0_n145, u1_u0_u0_n146, u1_u0_u0_n147, 
       u1_u0_u0_n148, u1_u0_u0_n149, u1_u0_u0_n150, u1_u0_u0_n151, u1_u0_u0_n152, u1_u0_u0_n153, u1_u0_u0_n154, u1_u0_u0_n155, u1_u0_u0_n156, 
       u1_u0_u0_n157, u1_u0_u0_n158, u1_u0_u0_n159, u1_u0_u0_n160, u1_u0_u0_n161, u1_u0_u0_n162, u1_u0_u0_n163, u1_u0_u0_n164, u1_u0_u0_n165, 
       u1_u0_u0_n166, u1_u0_u0_n167, u1_u0_u0_n168, u1_u0_u0_n169, u1_u0_u0_n170, u1_u0_u0_n171, u1_u0_u0_n172, u1_u0_u0_n173, u1_u0_u0_n174, 
       u1_u0_u0_n88, u1_u0_u0_n89, u1_u0_u0_n90, u1_u0_u0_n91, u1_u0_u0_n92, u1_u0_u0_n93, u1_u0_u0_n94, u1_u0_u0_n95, u1_u0_u0_n96, 
       u1_u0_u0_n97, u1_u0_u0_n98, u1_u0_u0_n99, u1_u0_u3_n100, u1_u0_u3_n101, u1_u0_u3_n102, u1_u0_u3_n103, u1_u0_u3_n104, u1_u0_u3_n105, 
       u1_u0_u3_n106, u1_u0_u3_n107, u1_u0_u3_n108, u1_u0_u3_n109, u1_u0_u3_n110, u1_u0_u3_n111, u1_u0_u3_n112, u1_u0_u3_n113, u1_u0_u3_n114, 
       u1_u0_u3_n115, u1_u0_u3_n116, u1_u0_u3_n117, u1_u0_u3_n118, u1_u0_u3_n119, u1_u0_u3_n120, u1_u0_u3_n121, u1_u0_u3_n122, u1_u0_u3_n123, 
       u1_u0_u3_n124, u1_u0_u3_n125, u1_u0_u3_n126, u1_u0_u3_n127, u1_u0_u3_n128, u1_u0_u3_n129, u1_u0_u3_n130, u1_u0_u3_n131, u1_u0_u3_n132, 
       u1_u0_u3_n133, u1_u0_u3_n134, u1_u0_u3_n135, u1_u0_u3_n136, u1_u0_u3_n137, u1_u0_u3_n138, u1_u0_u3_n139, u1_u0_u3_n140, u1_u0_u3_n141, 
       u1_u0_u3_n142, u1_u0_u3_n143, u1_u0_u3_n144, u1_u0_u3_n145, u1_u0_u3_n146, u1_u0_u3_n147, u1_u0_u3_n148, u1_u0_u3_n149, u1_u0_u3_n150, 
       u1_u0_u3_n151, u1_u0_u3_n152, u1_u0_u3_n153, u1_u0_u3_n154, u1_u0_u3_n155, u1_u0_u3_n156, u1_u0_u3_n157, u1_u0_u3_n158, u1_u0_u3_n159, 
       u1_u0_u3_n160, u1_u0_u3_n161, u1_u0_u3_n162, u1_u0_u3_n163, u1_u0_u3_n164, u1_u0_u3_n165, u1_u0_u3_n166, u1_u0_u3_n167, u1_u0_u3_n168, 
       u1_u0_u3_n169, u1_u0_u3_n170, u1_u0_u3_n171, u1_u0_u3_n172, u1_u0_u3_n173, u1_u0_u3_n174, u1_u0_u3_n175, u1_u0_u3_n176, u1_u0_u3_n177, 
       u1_u0_u3_n178, u1_u0_u3_n179, u1_u0_u3_n180, u1_u0_u3_n181, u1_u0_u3_n182, u1_u0_u3_n183, u1_u0_u3_n184, u1_u0_u3_n185, u1_u0_u3_n186, 
       u1_u0_u3_n94, u1_u0_u3_n95, u1_u0_u3_n96, u1_u0_u3_n97, u1_u0_u3_n98, u1_u0_u3_n99, u1_u10_X_10, u1_u10_X_11, u1_u10_X_12, 
       u1_u10_X_13, u1_u10_X_14, u1_u10_X_15, u1_u10_X_16, u1_u10_X_8, u1_u10_X_9, u1_u10_u1_n100, u1_u10_u1_n101, u1_u10_u1_n102, 
       u1_u10_u1_n103, u1_u10_u1_n104, u1_u10_u1_n105, u1_u10_u1_n106, u1_u10_u1_n107, u1_u10_u1_n108, u1_u10_u1_n109, u1_u10_u1_n110, u1_u10_u1_n111, 
       u1_u10_u1_n112, u1_u10_u1_n113, u1_u10_u1_n114, u1_u10_u1_n115, u1_u10_u1_n116, u1_u10_u1_n117, u1_u10_u1_n118, u1_u10_u1_n119, u1_u10_u1_n120, 
       u1_u10_u1_n121, u1_u10_u1_n122, u1_u10_u1_n123, u1_u10_u1_n124, u1_u10_u1_n125, u1_u10_u1_n126, u1_u10_u1_n127, u1_u10_u1_n128, u1_u10_u1_n129, 
       u1_u10_u1_n130, u1_u10_u1_n131, u1_u10_u1_n132, u1_u10_u1_n133, u1_u10_u1_n134, u1_u10_u1_n135, u1_u10_u1_n136, u1_u10_u1_n137, u1_u10_u1_n138, 
       u1_u10_u1_n139, u1_u10_u1_n140, u1_u10_u1_n141, u1_u10_u1_n142, u1_u10_u1_n143, u1_u10_u1_n144, u1_u10_u1_n145, u1_u10_u1_n146, u1_u10_u1_n147, 
       u1_u10_u1_n148, u1_u10_u1_n149, u1_u10_u1_n150, u1_u10_u1_n151, u1_u10_u1_n152, u1_u10_u1_n153, u1_u10_u1_n154, u1_u10_u1_n155, u1_u10_u1_n156, 
       u1_u10_u1_n157, u1_u10_u1_n158, u1_u10_u1_n159, u1_u10_u1_n160, u1_u10_u1_n161, u1_u10_u1_n162, u1_u10_u1_n163, u1_u10_u1_n164, u1_u10_u1_n165, 
       u1_u10_u1_n166, u1_u10_u1_n167, u1_u10_u1_n168, u1_u10_u1_n169, u1_u10_u1_n170, u1_u10_u1_n171, u1_u10_u1_n172, u1_u10_u1_n173, u1_u10_u1_n174, 
       u1_u10_u1_n175, u1_u10_u1_n176, u1_u10_u1_n177, u1_u10_u1_n178, u1_u10_u1_n179, u1_u10_u1_n180, u1_u10_u1_n181, u1_u10_u1_n182, u1_u10_u1_n183, 
       u1_u10_u1_n184, u1_u10_u1_n185, u1_u10_u1_n186, u1_u10_u1_n187, u1_u10_u1_n188, u1_u10_u1_n95, u1_u10_u1_n96, u1_u10_u1_n97, u1_u10_u1_n98, 
       u1_u10_u1_n99, u1_u10_u2_n100, u1_u10_u2_n101, u1_u10_u2_n102, u1_u10_u2_n103, u1_u10_u2_n104, u1_u10_u2_n105, u1_u10_u2_n106, u1_u10_u2_n107, 
       u1_u10_u2_n108, u1_u10_u2_n109, u1_u10_u2_n110, u1_u10_u2_n111, u1_u10_u2_n112, u1_u10_u2_n113, u1_u10_u2_n114, u1_u10_u2_n115, u1_u10_u2_n116, 
       u1_u10_u2_n117, u1_u10_u2_n118, u1_u10_u2_n119, u1_u10_u2_n120, u1_u10_u2_n121, u1_u10_u2_n122, u1_u10_u2_n123, u1_u10_u2_n124, u1_u10_u2_n125, 
       u1_u10_u2_n126, u1_u10_u2_n127, u1_u10_u2_n128, u1_u10_u2_n129, u1_u10_u2_n130, u1_u10_u2_n131, u1_u10_u2_n132, u1_u10_u2_n133, u1_u10_u2_n134, 
       u1_u10_u2_n135, u1_u10_u2_n136, u1_u10_u2_n137, u1_u10_u2_n138, u1_u10_u2_n139, u1_u10_u2_n140, u1_u10_u2_n141, u1_u10_u2_n142, u1_u10_u2_n143, 
       u1_u10_u2_n144, u1_u10_u2_n145, u1_u10_u2_n146, u1_u10_u2_n147, u1_u10_u2_n148, u1_u10_u2_n149, u1_u10_u2_n150, u1_u10_u2_n151, u1_u10_u2_n152, 
       u1_u10_u2_n153, u1_u10_u2_n154, u1_u10_u2_n155, u1_u10_u2_n156, u1_u10_u2_n157, u1_u10_u2_n158, u1_u10_u2_n159, u1_u10_u2_n160, u1_u10_u2_n161, 
       u1_u10_u2_n162, u1_u10_u2_n163, u1_u10_u2_n164, u1_u10_u2_n165, u1_u10_u2_n166, u1_u10_u2_n167, u1_u10_u2_n168, u1_u10_u2_n169, u1_u10_u2_n170, 
       u1_u10_u2_n171, u1_u10_u2_n172, u1_u10_u2_n173, u1_u10_u2_n174, u1_u10_u2_n175, u1_u10_u2_n176, u1_u10_u2_n177, u1_u10_u2_n178, u1_u10_u2_n179, 
       u1_u10_u2_n180, u1_u10_u2_n181, u1_u10_u2_n182, u1_u10_u2_n183, u1_u10_u2_n184, u1_u10_u2_n185, u1_u10_u2_n186, u1_u10_u2_n187, u1_u10_u2_n188, 
       u1_u10_u2_n95, u1_u10_u2_n96, u1_u10_u2_n97, u1_u10_u2_n98, u1_u10_u2_n99, u1_u11_X_10, u1_u11_X_11, u1_u11_X_12, u1_u11_X_13, 
       u1_u11_X_14, u1_u11_X_15, u1_u11_X_16, u1_u11_X_3, u1_u11_X_4, u1_u11_X_5, u1_u11_X_7, u1_u11_X_9, u1_u11_u0_n100, 
       u1_u11_u0_n101, u1_u11_u0_n102, u1_u11_u0_n103, u1_u11_u0_n104, u1_u11_u0_n105, u1_u11_u0_n106, u1_u11_u0_n107, u1_u11_u0_n108, u1_u11_u0_n109, 
       u1_u11_u0_n110, u1_u11_u0_n111, u1_u11_u0_n112, u1_u11_u0_n113, u1_u11_u0_n114, u1_u11_u0_n115, u1_u11_u0_n116, u1_u11_u0_n117, u1_u11_u0_n118, 
       u1_u11_u0_n119, u1_u11_u0_n120, u1_u11_u0_n121, u1_u11_u0_n122, u1_u11_u0_n123, u1_u11_u0_n124, u1_u11_u0_n125, u1_u11_u0_n126, u1_u11_u0_n127, 
       u1_u11_u0_n128, u1_u11_u0_n129, u1_u11_u0_n130, u1_u11_u0_n131, u1_u11_u0_n132, u1_u11_u0_n133, u1_u11_u0_n134, u1_u11_u0_n135, u1_u11_u0_n136, 
       u1_u11_u0_n137, u1_u11_u0_n138, u1_u11_u0_n139, u1_u11_u0_n140, u1_u11_u0_n141, u1_u11_u0_n142, u1_u11_u0_n143, u1_u11_u0_n144, u1_u11_u0_n145, 
       u1_u11_u0_n146, u1_u11_u0_n147, u1_u11_u0_n148, u1_u11_u0_n149, u1_u11_u0_n150, u1_u11_u0_n151, u1_u11_u0_n152, u1_u11_u0_n153, u1_u11_u0_n154, 
       u1_u11_u0_n155, u1_u11_u0_n156, u1_u11_u0_n157, u1_u11_u0_n158, u1_u11_u0_n159, u1_u11_u0_n160, u1_u11_u0_n161, u1_u11_u0_n162, u1_u11_u0_n163, 
       u1_u11_u0_n164, u1_u11_u0_n165, u1_u11_u0_n166, u1_u11_u0_n167, u1_u11_u0_n168, u1_u11_u0_n169, u1_u11_u0_n170, u1_u11_u0_n171, u1_u11_u0_n172, 
       u1_u11_u0_n173, u1_u11_u0_n174, u1_u11_u0_n88, u1_u11_u0_n89, u1_u11_u0_n90, u1_u11_u0_n91, u1_u11_u0_n92, u1_u11_u0_n93, u1_u11_u0_n94, 
       u1_u11_u0_n95, u1_u11_u0_n96, u1_u11_u0_n97, u1_u11_u0_n98, u1_u11_u0_n99, u1_u11_u1_n100, u1_u11_u1_n101, u1_u11_u1_n102, u1_u11_u1_n103, 
       u1_u11_u1_n104, u1_u11_u1_n105, u1_u11_u1_n106, u1_u11_u1_n107, u1_u11_u1_n108, u1_u11_u1_n109, u1_u11_u1_n110, u1_u11_u1_n111, u1_u11_u1_n112, 
       u1_u11_u1_n113, u1_u11_u1_n114, u1_u11_u1_n115, u1_u11_u1_n116, u1_u11_u1_n117, u1_u11_u1_n118, u1_u11_u1_n119, u1_u11_u1_n120, u1_u11_u1_n121, 
       u1_u11_u1_n122, u1_u11_u1_n123, u1_u11_u1_n124, u1_u11_u1_n125, u1_u11_u1_n126, u1_u11_u1_n127, u1_u11_u1_n128, u1_u11_u1_n129, u1_u11_u1_n130, 
       u1_u11_u1_n131, u1_u11_u1_n132, u1_u11_u1_n133, u1_u11_u1_n134, u1_u11_u1_n135, u1_u11_u1_n136, u1_u11_u1_n137, u1_u11_u1_n138, u1_u11_u1_n139, 
       u1_u11_u1_n140, u1_u11_u1_n141, u1_u11_u1_n142, u1_u11_u1_n143, u1_u11_u1_n144, u1_u11_u1_n145, u1_u11_u1_n146, u1_u11_u1_n147, u1_u11_u1_n148, 
       u1_u11_u1_n149, u1_u11_u1_n150, u1_u11_u1_n151, u1_u11_u1_n152, u1_u11_u1_n153, u1_u11_u1_n154, u1_u11_u1_n155, u1_u11_u1_n156, u1_u11_u1_n157, 
       u1_u11_u1_n158, u1_u11_u1_n159, u1_u11_u1_n160, u1_u11_u1_n161, u1_u11_u1_n162, u1_u11_u1_n163, u1_u11_u1_n164, u1_u11_u1_n165, u1_u11_u1_n166, 
       u1_u11_u1_n167, u1_u11_u1_n168, u1_u11_u1_n169, u1_u11_u1_n170, u1_u11_u1_n171, u1_u11_u1_n172, u1_u11_u1_n173, u1_u11_u1_n174, u1_u11_u1_n175, 
       u1_u11_u1_n176, u1_u11_u1_n177, u1_u11_u1_n178, u1_u11_u1_n179, u1_u11_u1_n180, u1_u11_u1_n181, u1_u11_u1_n182, u1_u11_u1_n183, u1_u11_u1_n184, 
       u1_u11_u1_n185, u1_u11_u1_n186, u1_u11_u1_n187, u1_u11_u1_n188, u1_u11_u1_n95, u1_u11_u1_n96, u1_u11_u1_n97, u1_u11_u1_n98, u1_u11_u1_n99, 
       u1_u11_u2_n100, u1_u11_u2_n101, u1_u11_u2_n102, u1_u11_u2_n103, u1_u11_u2_n104, u1_u11_u2_n105, u1_u11_u2_n106, u1_u11_u2_n107, u1_u11_u2_n108, 
       u1_u11_u2_n109, u1_u11_u2_n110, u1_u11_u2_n111, u1_u11_u2_n112, u1_u11_u2_n113, u1_u11_u2_n114, u1_u11_u2_n115, u1_u11_u2_n116, u1_u11_u2_n117, 
       u1_u11_u2_n118, u1_u11_u2_n119, u1_u11_u2_n120, u1_u11_u2_n121, u1_u11_u2_n122, u1_u11_u2_n123, u1_u11_u2_n124, u1_u11_u2_n125, u1_u11_u2_n126, 
       u1_u11_u2_n127, u1_u11_u2_n128, u1_u11_u2_n129, u1_u11_u2_n130, u1_u11_u2_n131, u1_u11_u2_n132, u1_u11_u2_n133, u1_u11_u2_n134, u1_u11_u2_n135, 
       u1_u11_u2_n136, u1_u11_u2_n137, u1_u11_u2_n138, u1_u11_u2_n139, u1_u11_u2_n140, u1_u11_u2_n141, u1_u11_u2_n142, u1_u11_u2_n143, u1_u11_u2_n144, 
       u1_u11_u2_n145, u1_u11_u2_n146, u1_u11_u2_n147, u1_u11_u2_n148, u1_u11_u2_n149, u1_u11_u2_n150, u1_u11_u2_n151, u1_u11_u2_n152, u1_u11_u2_n153, 
       u1_u11_u2_n154, u1_u11_u2_n155, u1_u11_u2_n156, u1_u11_u2_n157, u1_u11_u2_n158, u1_u11_u2_n159, u1_u11_u2_n160, u1_u11_u2_n161, u1_u11_u2_n162, 
       u1_u11_u2_n163, u1_u11_u2_n164, u1_u11_u2_n165, u1_u11_u2_n166, u1_u11_u2_n167, u1_u11_u2_n168, u1_u11_u2_n169, u1_u11_u2_n170, u1_u11_u2_n171, 
       u1_u11_u2_n172, u1_u11_u2_n173, u1_u11_u2_n174, u1_u11_u2_n175, u1_u11_u2_n176, u1_u11_u2_n177, u1_u11_u2_n178, u1_u11_u2_n179, u1_u11_u2_n180, 
       u1_u11_u2_n181, u1_u11_u2_n182, u1_u11_u2_n183, u1_u11_u2_n184, u1_u11_u2_n185, u1_u11_u2_n186, u1_u11_u2_n187, u1_u11_u2_n188, u1_u11_u2_n95, 
       u1_u11_u2_n96, u1_u11_u2_n97, u1_u11_u2_n98, u1_u11_u2_n99, u1_u12_X_1, u1_u12_X_21, u1_u12_X_22, u1_u12_X_24, u1_u12_X_26, 
       u1_u12_X_27, u1_u12_X_28, u1_u12_X_3, u1_u12_X_4, u1_u12_X_45, u1_u12_X_46, u1_u12_X_47, u1_u12_X_6, u1_u12_u0_n100, 
       u1_u12_u0_n101, u1_u12_u0_n102, u1_u12_u0_n103, u1_u12_u0_n104, u1_u12_u0_n105, u1_u12_u0_n106, u1_u12_u0_n107, u1_u12_u0_n108, u1_u12_u0_n109, 
       u1_u12_u0_n110, u1_u12_u0_n111, u1_u12_u0_n112, u1_u12_u0_n113, u1_u12_u0_n114, u1_u12_u0_n115, u1_u12_u0_n116, u1_u12_u0_n117, u1_u12_u0_n118, 
       u1_u12_u0_n119, u1_u12_u0_n120, u1_u12_u0_n121, u1_u12_u0_n122, u1_u12_u0_n123, u1_u12_u0_n124, u1_u12_u0_n125, u1_u12_u0_n126, u1_u12_u0_n127, 
       u1_u12_u0_n128, u1_u12_u0_n129, u1_u12_u0_n130, u1_u12_u0_n131, u1_u12_u0_n132, u1_u12_u0_n133, u1_u12_u0_n134, u1_u12_u0_n135, u1_u12_u0_n136, 
       u1_u12_u0_n137, u1_u12_u0_n138, u1_u12_u0_n139, u1_u12_u0_n140, u1_u12_u0_n141, u1_u12_u0_n142, u1_u12_u0_n143, u1_u12_u0_n144, u1_u12_u0_n145, 
       u1_u12_u0_n146, u1_u12_u0_n147, u1_u12_u0_n148, u1_u12_u0_n149, u1_u12_u0_n150, u1_u12_u0_n151, u1_u12_u0_n152, u1_u12_u0_n153, u1_u12_u0_n154, 
       u1_u12_u0_n155, u1_u12_u0_n156, u1_u12_u0_n157, u1_u12_u0_n158, u1_u12_u0_n159, u1_u12_u0_n160, u1_u12_u0_n161, u1_u12_u0_n162, u1_u12_u0_n163, 
       u1_u12_u0_n164, u1_u12_u0_n165, u1_u12_u0_n166, u1_u12_u0_n167, u1_u12_u0_n168, u1_u12_u0_n169, u1_u12_u0_n170, u1_u12_u0_n171, u1_u12_u0_n172, 
       u1_u12_u0_n173, u1_u12_u0_n174, u1_u12_u0_n88, u1_u12_u0_n89, u1_u12_u0_n90, u1_u12_u0_n91, u1_u12_u0_n92, u1_u12_u0_n93, u1_u12_u0_n94, 
       u1_u12_u0_n95, u1_u12_u0_n96, u1_u12_u0_n97, u1_u12_u0_n98, u1_u12_u0_n99, u1_u12_u3_n100, u1_u12_u3_n101, u1_u12_u3_n102, u1_u12_u3_n103, 
       u1_u12_u3_n104, u1_u12_u3_n105, u1_u12_u3_n106, u1_u12_u3_n107, u1_u12_u3_n108, u1_u12_u3_n109, u1_u12_u3_n110, u1_u12_u3_n111, u1_u12_u3_n112, 
       u1_u12_u3_n113, u1_u12_u3_n114, u1_u12_u3_n115, u1_u12_u3_n116, u1_u12_u3_n117, u1_u12_u3_n118, u1_u12_u3_n119, u1_u12_u3_n120, u1_u12_u3_n121, 
       u1_u12_u3_n122, u1_u12_u3_n123, u1_u12_u3_n124, u1_u12_u3_n125, u1_u12_u3_n126, u1_u12_u3_n127, u1_u12_u3_n128, u1_u12_u3_n129, u1_u12_u3_n130, 
       u1_u12_u3_n131, u1_u12_u3_n132, u1_u12_u3_n133, u1_u12_u3_n134, u1_u12_u3_n135, u1_u12_u3_n136, u1_u12_u3_n137, u1_u12_u3_n138, u1_u12_u3_n139, 
       u1_u12_u3_n140, u1_u12_u3_n141, u1_u12_u3_n142, u1_u12_u3_n143, u1_u12_u3_n144, u1_u12_u3_n145, u1_u12_u3_n146, u1_u12_u3_n147, u1_u12_u3_n148, 
       u1_u12_u3_n149, u1_u12_u3_n150, u1_u12_u3_n151, u1_u12_u3_n152, u1_u12_u3_n153, u1_u12_u3_n154, u1_u12_u3_n155, u1_u12_u3_n156, u1_u12_u3_n157, 
       u1_u12_u3_n158, u1_u12_u3_n159, u1_u12_u3_n160, u1_u12_u3_n161, u1_u12_u3_n162, u1_u12_u3_n163, u1_u12_u3_n164, u1_u12_u3_n165, u1_u12_u3_n166, 
       u1_u12_u3_n167, u1_u12_u3_n168, u1_u12_u3_n169, u1_u12_u3_n170, u1_u12_u3_n171, u1_u12_u3_n172, u1_u12_u3_n173, u1_u12_u3_n174, u1_u12_u3_n175, 
       u1_u12_u3_n176, u1_u12_u3_n177, u1_u12_u3_n178, u1_u12_u3_n179, u1_u12_u3_n180, u1_u12_u3_n181, u1_u12_u3_n182, u1_u12_u3_n183, u1_u12_u3_n184, 
       u1_u12_u3_n185, u1_u12_u3_n186, u1_u12_u3_n94, u1_u12_u3_n95, u1_u12_u3_n96, u1_u12_u3_n97, u1_u12_u3_n98, u1_u12_u3_n99, u1_u12_u4_n100, 
       u1_u12_u4_n101, u1_u12_u4_n102, u1_u12_u4_n103, u1_u12_u4_n104, u1_u12_u4_n105, u1_u12_u4_n106, u1_u12_u4_n107, u1_u12_u4_n108, u1_u12_u4_n109, 
       u1_u12_u4_n110, u1_u12_u4_n111, u1_u12_u4_n112, u1_u12_u4_n113, u1_u12_u4_n114, u1_u12_u4_n115, u1_u12_u4_n116, u1_u12_u4_n117, u1_u12_u4_n118, 
       u1_u12_u4_n119, u1_u12_u4_n120, u1_u12_u4_n121, u1_u12_u4_n122, u1_u12_u4_n123, u1_u12_u4_n124, u1_u12_u4_n125, u1_u12_u4_n126, u1_u12_u4_n127, 
       u1_u12_u4_n128, u1_u12_u4_n129, u1_u12_u4_n130, u1_u12_u4_n131, u1_u12_u4_n132, u1_u12_u4_n133, u1_u12_u4_n134, u1_u12_u4_n135, u1_u12_u4_n136, 
       u1_u12_u4_n137, u1_u12_u4_n138, u1_u12_u4_n139, u1_u12_u4_n140, u1_u12_u4_n141, u1_u12_u4_n142, u1_u12_u4_n143, u1_u12_u4_n144, u1_u12_u4_n145, 
       u1_u12_u4_n146, u1_u12_u4_n147, u1_u12_u4_n148, u1_u12_u4_n149, u1_u12_u4_n150, u1_u12_u4_n151, u1_u12_u4_n152, u1_u12_u4_n153, u1_u12_u4_n154, 
       u1_u12_u4_n155, u1_u12_u4_n156, u1_u12_u4_n157, u1_u12_u4_n158, u1_u12_u4_n159, u1_u12_u4_n160, u1_u12_u4_n161, u1_u12_u4_n162, u1_u12_u4_n163, 
       u1_u12_u4_n164, u1_u12_u4_n165, u1_u12_u4_n166, u1_u12_u4_n167, u1_u12_u4_n168, u1_u12_u4_n169, u1_u12_u4_n170, u1_u12_u4_n171, u1_u12_u4_n172, 
       u1_u12_u4_n173, u1_u12_u4_n174, u1_u12_u4_n175, u1_u12_u4_n176, u1_u12_u4_n177, u1_u12_u4_n178, u1_u12_u4_n179, u1_u12_u4_n180, u1_u12_u4_n181, 
       u1_u12_u4_n182, u1_u12_u4_n183, u1_u12_u4_n184, u1_u12_u4_n185, u1_u12_u4_n186, u1_u12_u4_n94, u1_u12_u4_n95, u1_u12_u4_n96, u1_u12_u4_n97, 
       u1_u12_u4_n98, u1_u12_u4_n99, u1_u12_u7_n100, u1_u12_u7_n101, u1_u12_u7_n102, u1_u12_u7_n103, u1_u12_u7_n104, u1_u12_u7_n105, u1_u12_u7_n106, 
       u1_u12_u7_n107, u1_u12_u7_n108, u1_u12_u7_n109, u1_u12_u7_n110, u1_u12_u7_n111, u1_u12_u7_n112, u1_u12_u7_n113, u1_u12_u7_n114, u1_u12_u7_n115, 
       u1_u12_u7_n116, u1_u12_u7_n117, u1_u12_u7_n118, u1_u12_u7_n119, u1_u12_u7_n120, u1_u12_u7_n121, u1_u12_u7_n122, u1_u12_u7_n123, u1_u12_u7_n124, 
       u1_u12_u7_n125, u1_u12_u7_n126, u1_u12_u7_n127, u1_u12_u7_n128, u1_u12_u7_n129, u1_u12_u7_n130, u1_u12_u7_n131, u1_u12_u7_n132, u1_u12_u7_n133, 
       u1_u12_u7_n134, u1_u12_u7_n135, u1_u12_u7_n136, u1_u12_u7_n137, u1_u12_u7_n138, u1_u12_u7_n139, u1_u12_u7_n140, u1_u12_u7_n141, u1_u12_u7_n142, 
       u1_u12_u7_n143, u1_u12_u7_n144, u1_u12_u7_n145, u1_u12_u7_n146, u1_u12_u7_n147, u1_u12_u7_n148, u1_u12_u7_n149, u1_u12_u7_n150, u1_u12_u7_n151, 
       u1_u12_u7_n152, u1_u12_u7_n153, u1_u12_u7_n154, u1_u12_u7_n155, u1_u12_u7_n156, u1_u12_u7_n157, u1_u12_u7_n158, u1_u12_u7_n159, u1_u12_u7_n160, 
       u1_u12_u7_n161, u1_u12_u7_n162, u1_u12_u7_n163, u1_u12_u7_n164, u1_u12_u7_n165, u1_u12_u7_n166, u1_u12_u7_n167, u1_u12_u7_n168, u1_u12_u7_n169, 
       u1_u12_u7_n170, u1_u12_u7_n171, u1_u12_u7_n172, u1_u12_u7_n173, u1_u12_u7_n174, u1_u12_u7_n175, u1_u12_u7_n176, u1_u12_u7_n177, u1_u12_u7_n178, 
       u1_u12_u7_n179, u1_u12_u7_n180, u1_u12_u7_n91, u1_u12_u7_n92, u1_u12_u7_n93, u1_u12_u7_n94, u1_u12_u7_n95, u1_u12_u7_n96, u1_u12_u7_n97, 
       u1_u12_u7_n98, u1_u12_u7_n99, u1_u14_X_14, u1_u14_X_15, u1_u14_X_16, u1_u14_X_17, u1_u14_X_18, u1_u14_X_19, u1_u14_X_20, 
       u1_u14_X_21, u1_u14_X_22, u1_u14_u2_n100, u1_u14_u2_n101, u1_u14_u2_n102, u1_u14_u2_n103, u1_u14_u2_n104, u1_u14_u2_n105, u1_u14_u2_n106, 
       u1_u14_u2_n107, u1_u14_u2_n108, u1_u14_u2_n109, u1_u14_u2_n110, u1_u14_u2_n111, u1_u14_u2_n112, u1_u14_u2_n113, u1_u14_u2_n114, u1_u14_u2_n115, 
       u1_u14_u2_n116, u1_u14_u2_n117, u1_u14_u2_n118, u1_u14_u2_n119, u1_u14_u2_n120, u1_u14_u2_n121, u1_u14_u2_n122, u1_u14_u2_n123, u1_u14_u2_n124, 
       u1_u14_u2_n125, u1_u14_u2_n126, u1_u14_u2_n127, u1_u14_u2_n128, u1_u14_u2_n129, u1_u14_u2_n130, u1_u14_u2_n131, u1_u14_u2_n132, u1_u14_u2_n133, 
       u1_u14_u2_n134, u1_u14_u2_n135, u1_u14_u2_n136, u1_u14_u2_n137, u1_u14_u2_n138, u1_u14_u2_n139, u1_u14_u2_n140, u1_u14_u2_n141, u1_u14_u2_n142, 
       u1_u14_u2_n143, u1_u14_u2_n144, u1_u14_u2_n145, u1_u14_u2_n146, u1_u14_u2_n147, u1_u14_u2_n148, u1_u14_u2_n149, u1_u14_u2_n150, u1_u14_u2_n151, 
       u1_u14_u2_n152, u1_u14_u2_n153, u1_u14_u2_n154, u1_u14_u2_n155, u1_u14_u2_n156, u1_u14_u2_n157, u1_u14_u2_n158, u1_u14_u2_n159, u1_u14_u2_n160, 
       u1_u14_u2_n161, u1_u14_u2_n162, u1_u14_u2_n163, u1_u14_u2_n164, u1_u14_u2_n165, u1_u14_u2_n166, u1_u14_u2_n167, u1_u14_u2_n168, u1_u14_u2_n169, 
       u1_u14_u2_n170, u1_u14_u2_n171, u1_u14_u2_n172, u1_u14_u2_n173, u1_u14_u2_n174, u1_u14_u2_n175, u1_u14_u2_n176, u1_u14_u2_n177, u1_u14_u2_n178, 
       u1_u14_u2_n179, u1_u14_u2_n180, u1_u14_u2_n181, u1_u14_u2_n182, u1_u14_u2_n183, u1_u14_u2_n184, u1_u14_u2_n185, u1_u14_u2_n186, u1_u14_u2_n187, 
       u1_u14_u2_n188, u1_u14_u2_n95, u1_u14_u2_n96, u1_u14_u2_n97, u1_u14_u2_n98, u1_u14_u2_n99, u1_u14_u3_n100, u1_u14_u3_n101, u1_u14_u3_n102, 
       u1_u14_u3_n103, u1_u14_u3_n104, u1_u14_u3_n105, u1_u14_u3_n106, u1_u14_u3_n107, u1_u14_u3_n108, u1_u14_u3_n109, u1_u14_u3_n110, u1_u14_u3_n111, 
       u1_u14_u3_n112, u1_u14_u3_n113, u1_u14_u3_n114, u1_u14_u3_n115, u1_u14_u3_n116, u1_u14_u3_n117, u1_u14_u3_n118, u1_u14_u3_n119, u1_u14_u3_n120, 
       u1_u14_u3_n121, u1_u14_u3_n122, u1_u14_u3_n123, u1_u14_u3_n124, u1_u14_u3_n125, u1_u14_u3_n126, u1_u14_u3_n127, u1_u14_u3_n128, u1_u14_u3_n129, 
       u1_u14_u3_n130, u1_u14_u3_n131, u1_u14_u3_n132, u1_u14_u3_n133, u1_u14_u3_n134, u1_u14_u3_n135, u1_u14_u3_n136, u1_u14_u3_n137, u1_u14_u3_n138, 
       u1_u14_u3_n139, u1_u14_u3_n140, u1_u14_u3_n141, u1_u14_u3_n142, u1_u14_u3_n143, u1_u14_u3_n144, u1_u14_u3_n145, u1_u14_u3_n146, u1_u14_u3_n147, 
       u1_u14_u3_n148, u1_u14_u3_n149, u1_u14_u3_n150, u1_u14_u3_n151, u1_u14_u3_n152, u1_u14_u3_n153, u1_u14_u3_n154, u1_u14_u3_n155, u1_u14_u3_n156, 
       u1_u14_u3_n157, u1_u14_u3_n158, u1_u14_u3_n159, u1_u14_u3_n160, u1_u14_u3_n161, u1_u14_u3_n162, u1_u14_u3_n163, u1_u14_u3_n164, u1_u14_u3_n165, 
       u1_u14_u3_n166, u1_u14_u3_n167, u1_u14_u3_n168, u1_u14_u3_n169, u1_u14_u3_n170, u1_u14_u3_n171, u1_u14_u3_n172, u1_u14_u3_n173, u1_u14_u3_n174, 
       u1_u14_u3_n175, u1_u14_u3_n176, u1_u14_u3_n177, u1_u14_u3_n178, u1_u14_u3_n179, u1_u14_u3_n180, u1_u14_u3_n181, u1_u14_u3_n182, u1_u14_u3_n183, 
       u1_u14_u3_n184, u1_u14_u3_n185, u1_u14_u3_n186, u1_u14_u3_n94, u1_u14_u3_n95, u1_u14_u3_n96, u1_u14_u3_n97, u1_u14_u3_n98, u1_u14_u3_n99, 
       u1_u15_X_10, u1_u15_X_3, u1_u15_X_4, u1_u15_X_6, u1_u15_X_8, u1_u15_X_9, u1_u15_u0_n100, u1_u15_u0_n101, u1_u15_u0_n102, 
       u1_u15_u0_n103, u1_u15_u0_n104, u1_u15_u0_n105, u1_u15_u0_n106, u1_u15_u0_n107, u1_u15_u0_n108, u1_u15_u0_n109, u1_u15_u0_n110, u1_u15_u0_n111, 
       u1_u15_u0_n112, u1_u15_u0_n113, u1_u15_u0_n114, u1_u15_u0_n115, u1_u15_u0_n116, u1_u15_u0_n117, u1_u15_u0_n118, u1_u15_u0_n119, u1_u15_u0_n120, 
       u1_u15_u0_n121, u1_u15_u0_n122, u1_u15_u0_n123, u1_u15_u0_n124, u1_u15_u0_n125, u1_u15_u0_n126, u1_u15_u0_n127, u1_u15_u0_n128, u1_u15_u0_n129, 
       u1_u15_u0_n130, u1_u15_u0_n131, u1_u15_u0_n132, u1_u15_u0_n133, u1_u15_u0_n134, u1_u15_u0_n135, u1_u15_u0_n136, u1_u15_u0_n137, u1_u15_u0_n138, 
       u1_u15_u0_n139, u1_u15_u0_n140, u1_u15_u0_n141, u1_u15_u0_n142, u1_u15_u0_n143, u1_u15_u0_n144, u1_u15_u0_n145, u1_u15_u0_n146, u1_u15_u0_n147, 
       u1_u15_u0_n148, u1_u15_u0_n149, u1_u15_u0_n150, u1_u15_u0_n151, u1_u15_u0_n152, u1_u15_u0_n153, u1_u15_u0_n154, u1_u15_u0_n155, u1_u15_u0_n156, 
       u1_u15_u0_n157, u1_u15_u0_n158, u1_u15_u0_n159, u1_u15_u0_n160, u1_u15_u0_n161, u1_u15_u0_n162, u1_u15_u0_n163, u1_u15_u0_n164, u1_u15_u0_n165, 
       u1_u15_u0_n166, u1_u15_u0_n167, u1_u15_u0_n168, u1_u15_u0_n169, u1_u15_u0_n170, u1_u15_u0_n171, u1_u15_u0_n172, u1_u15_u0_n173, u1_u15_u0_n174, 
       u1_u15_u0_n88, u1_u15_u0_n89, u1_u15_u0_n90, u1_u15_u0_n91, u1_u15_u0_n92, u1_u15_u0_n93, u1_u15_u0_n94, u1_u15_u0_n95, u1_u15_u0_n96, 
       u1_u15_u0_n97, u1_u15_u0_n98, u1_u15_u0_n99, u1_u15_u1_n100, u1_u15_u1_n101, u1_u15_u1_n102, u1_u15_u1_n103, u1_u15_u1_n104, u1_u15_u1_n105, 
       u1_u15_u1_n106, u1_u15_u1_n107, u1_u15_u1_n108, u1_u15_u1_n109, u1_u15_u1_n110, u1_u15_u1_n111, u1_u15_u1_n112, u1_u15_u1_n113, u1_u15_u1_n114, 
       u1_u15_u1_n115, u1_u15_u1_n116, u1_u15_u1_n117, u1_u15_u1_n118, u1_u15_u1_n119, u1_u15_u1_n120, u1_u15_u1_n121, u1_u15_u1_n122, u1_u15_u1_n123, 
       u1_u15_u1_n124, u1_u15_u1_n125, u1_u15_u1_n126, u1_u15_u1_n127, u1_u15_u1_n128, u1_u15_u1_n129, u1_u15_u1_n130, u1_u15_u1_n131, u1_u15_u1_n132, 
       u1_u15_u1_n133, u1_u15_u1_n134, u1_u15_u1_n135, u1_u15_u1_n136, u1_u15_u1_n137, u1_u15_u1_n138, u1_u15_u1_n139, u1_u15_u1_n140, u1_u15_u1_n141, 
       u1_u15_u1_n142, u1_u15_u1_n143, u1_u15_u1_n144, u1_u15_u1_n145, u1_u15_u1_n146, u1_u15_u1_n147, u1_u15_u1_n148, u1_u15_u1_n149, u1_u15_u1_n150, 
       u1_u15_u1_n151, u1_u15_u1_n152, u1_u15_u1_n153, u1_u15_u1_n154, u1_u15_u1_n155, u1_u15_u1_n156, u1_u15_u1_n157, u1_u15_u1_n158, u1_u15_u1_n159, 
       u1_u15_u1_n160, u1_u15_u1_n161, u1_u15_u1_n162, u1_u15_u1_n163, u1_u15_u1_n164, u1_u15_u1_n165, u1_u15_u1_n166, u1_u15_u1_n167, u1_u15_u1_n168, 
       u1_u15_u1_n169, u1_u15_u1_n170, u1_u15_u1_n171, u1_u15_u1_n172, u1_u15_u1_n173, u1_u15_u1_n174, u1_u15_u1_n175, u1_u15_u1_n176, u1_u15_u1_n177, 
       u1_u15_u1_n178, u1_u15_u1_n179, u1_u15_u1_n180, u1_u15_u1_n181, u1_u15_u1_n182, u1_u15_u1_n183, u1_u15_u1_n184, u1_u15_u1_n185, u1_u15_u1_n186, 
       u1_u15_u1_n187, u1_u15_u1_n188, u1_u15_u1_n95, u1_u15_u1_n96, u1_u15_u1_n97, u1_u15_u1_n98, u1_u15_u1_n99, u1_u1_X_33, u1_u1_X_34, 
       u1_u1_u5_n100, u1_u1_u5_n101, u1_u1_u5_n102, u1_u1_u5_n103, u1_u1_u5_n104, u1_u1_u5_n105, u1_u1_u5_n106, u1_u1_u5_n107, u1_u1_u5_n108, 
       u1_u1_u5_n109, u1_u1_u5_n110, u1_u1_u5_n111, u1_u1_u5_n112, u1_u1_u5_n113, u1_u1_u5_n114, u1_u1_u5_n115, u1_u1_u5_n116, u1_u1_u5_n117, 
       u1_u1_u5_n118, u1_u1_u5_n119, u1_u1_u5_n120, u1_u1_u5_n121, u1_u1_u5_n122, u1_u1_u5_n123, u1_u1_u5_n124, u1_u1_u5_n125, u1_u1_u5_n126, 
       u1_u1_u5_n127, u1_u1_u5_n128, u1_u1_u5_n129, u1_u1_u5_n130, u1_u1_u5_n131, u1_u1_u5_n132, u1_u1_u5_n133, u1_u1_u5_n134, u1_u1_u5_n135, 
       u1_u1_u5_n136, u1_u1_u5_n137, u1_u1_u5_n138, u1_u1_u5_n139, u1_u1_u5_n140, u1_u1_u5_n141, u1_u1_u5_n142, u1_u1_u5_n143, u1_u1_u5_n144, 
       u1_u1_u5_n145, u1_u1_u5_n146, u1_u1_u5_n147, u1_u1_u5_n148, u1_u1_u5_n149, u1_u1_u5_n150, u1_u1_u5_n151, u1_u1_u5_n152, u1_u1_u5_n153, 
       u1_u1_u5_n154, u1_u1_u5_n155, u1_u1_u5_n156, u1_u1_u5_n157, u1_u1_u5_n158, u1_u1_u5_n159, u1_u1_u5_n160, u1_u1_u5_n161, u1_u1_u5_n162, 
       u1_u1_u5_n163, u1_u1_u5_n164, u1_u1_u5_n165, u1_u1_u5_n166, u1_u1_u5_n167, u1_u1_u5_n168, u1_u1_u5_n169, u1_u1_u5_n170, u1_u1_u5_n171, 
       u1_u1_u5_n172, u1_u1_u5_n173, u1_u1_u5_n174, u1_u1_u5_n175, u1_u1_u5_n176, u1_u1_u5_n177, u1_u1_u5_n178, u1_u1_u5_n179, u1_u1_u5_n180, 
       u1_u1_u5_n181, u1_u1_u5_n182, u1_u1_u5_n183, u1_u1_u5_n184, u1_u1_u5_n185, u1_u1_u5_n186, u1_u1_u5_n187, u1_u1_u5_n188, u1_u1_u5_n189, 
       u1_u1_u5_n190, u1_u1_u5_n191, u1_u1_u5_n192, u1_u1_u5_n193, u1_u1_u5_n194, u1_u1_u5_n195, u1_u1_u5_n196, u1_u1_u5_n99, u1_u2_X_10, 
       u1_u2_X_3, u1_u2_X_4, u1_u2_X_5, u1_u2_X_7, u1_u2_X_9, u1_u2_u0_n100, u1_u2_u0_n101, u1_u2_u0_n102, u1_u2_u0_n103, 
       u1_u2_u0_n104, u1_u2_u0_n105, u1_u2_u0_n106, u1_u2_u0_n107, u1_u2_u0_n108, u1_u2_u0_n109, u1_u2_u0_n110, u1_u2_u0_n111, u1_u2_u0_n112, 
       u1_u2_u0_n113, u1_u2_u0_n114, u1_u2_u0_n115, u1_u2_u0_n116, u1_u2_u0_n117, u1_u2_u0_n118, u1_u2_u0_n119, u1_u2_u0_n120, u1_u2_u0_n121, 
       u1_u2_u0_n122, u1_u2_u0_n123, u1_u2_u0_n124, u1_u2_u0_n125, u1_u2_u0_n126, u1_u2_u0_n127, u1_u2_u0_n128, u1_u2_u0_n129, u1_u2_u0_n130, 
       u1_u2_u0_n131, u1_u2_u0_n132, u1_u2_u0_n133, u1_u2_u0_n134, u1_u2_u0_n135, u1_u2_u0_n136, u1_u2_u0_n137, u1_u2_u0_n138, u1_u2_u0_n139, 
       u1_u2_u0_n140, u1_u2_u0_n141, u1_u2_u0_n142, u1_u2_u0_n143, u1_u2_u0_n144, u1_u2_u0_n145, u1_u2_u0_n146, u1_u2_u0_n147, u1_u2_u0_n148, 
       u1_u2_u0_n149, u1_u2_u0_n150, u1_u2_u0_n151, u1_u2_u0_n152, u1_u2_u0_n153, u1_u2_u0_n154, u1_u2_u0_n155, u1_u2_u0_n156, u1_u2_u0_n157, 
       u1_u2_u0_n158, u1_u2_u0_n159, u1_u2_u0_n160, u1_u2_u0_n161, u1_u2_u0_n162, u1_u2_u0_n163, u1_u2_u0_n164, u1_u2_u0_n165, u1_u2_u0_n166, 
       u1_u2_u0_n167, u1_u2_u0_n168, u1_u2_u0_n169, u1_u2_u0_n170, u1_u2_u0_n171, u1_u2_u0_n172, u1_u2_u0_n173, u1_u2_u0_n174, u1_u2_u0_n88, 
       u1_u2_u0_n89, u1_u2_u0_n90, u1_u2_u0_n91, u1_u2_u0_n92, u1_u2_u0_n93, u1_u2_u0_n94, u1_u2_u0_n95, u1_u2_u0_n96, u1_u2_u0_n97, 
       u1_u2_u0_n98, u1_u2_u0_n99, u1_u2_u1_n100, u1_u2_u1_n101, u1_u2_u1_n102, u1_u2_u1_n103, u1_u2_u1_n104, u1_u2_u1_n105, u1_u2_u1_n106, 
       u1_u2_u1_n107, u1_u2_u1_n108, u1_u2_u1_n109, u1_u2_u1_n110, u1_u2_u1_n111, u1_u2_u1_n112, u1_u2_u1_n113, u1_u2_u1_n114, u1_u2_u1_n115, 
       u1_u2_u1_n116, u1_u2_u1_n117, u1_u2_u1_n118, u1_u2_u1_n119, u1_u2_u1_n120, u1_u2_u1_n121, u1_u2_u1_n122, u1_u2_u1_n123, u1_u2_u1_n124, 
       u1_u2_u1_n125, u1_u2_u1_n126, u1_u2_u1_n127, u1_u2_u1_n128, u1_u2_u1_n129, u1_u2_u1_n130, u1_u2_u1_n131, u1_u2_u1_n132, u1_u2_u1_n133, 
       u1_u2_u1_n134, u1_u2_u1_n135, u1_u2_u1_n136, u1_u2_u1_n137, u1_u2_u1_n138, u1_u2_u1_n139, u1_u2_u1_n140, u1_u2_u1_n141, u1_u2_u1_n142, 
       u1_u2_u1_n143, u1_u2_u1_n144, u1_u2_u1_n145, u1_u2_u1_n146, u1_u2_u1_n147, u1_u2_u1_n148, u1_u2_u1_n149, u1_u2_u1_n150, u1_u2_u1_n151, 
       u1_u2_u1_n152, u1_u2_u1_n153, u1_u2_u1_n154, u1_u2_u1_n155, u1_u2_u1_n156, u1_u2_u1_n157, u1_u2_u1_n158, u1_u2_u1_n159, u1_u2_u1_n160, 
       u1_u2_u1_n161, u1_u2_u1_n162, u1_u2_u1_n163, u1_u2_u1_n164, u1_u2_u1_n165, u1_u2_u1_n166, u1_u2_u1_n167, u1_u2_u1_n168, u1_u2_u1_n169, 
       u1_u2_u1_n170, u1_u2_u1_n171, u1_u2_u1_n172, u1_u2_u1_n173, u1_u2_u1_n174, u1_u2_u1_n175, u1_u2_u1_n176, u1_u2_u1_n177, u1_u2_u1_n178, 
       u1_u2_u1_n179, u1_u2_u1_n180, u1_u2_u1_n181, u1_u2_u1_n182, u1_u2_u1_n183, u1_u2_u1_n184, u1_u2_u1_n185, u1_u2_u1_n186, u1_u2_u1_n187, 
       u1_u2_u1_n188, u1_u2_u1_n95, u1_u2_u1_n96, u1_u2_u1_n97, u1_u2_u1_n98, u1_u2_u1_n99, u1_u3_X_45, u1_u3_X_46, u1_u3_u7_n100, 
       u1_u3_u7_n101, u1_u3_u7_n102, u1_u3_u7_n103, u1_u3_u7_n104, u1_u3_u7_n105, u1_u3_u7_n106, u1_u3_u7_n107, u1_u3_u7_n108, u1_u3_u7_n109, 
       u1_u3_u7_n110, u1_u3_u7_n111, u1_u3_u7_n112, u1_u3_u7_n113, u1_u3_u7_n114, u1_u3_u7_n115, u1_u3_u7_n116, u1_u3_u7_n117, u1_u3_u7_n118, 
       u1_u3_u7_n119, u1_u3_u7_n120, u1_u3_u7_n121, u1_u3_u7_n122, u1_u3_u7_n123, u1_u3_u7_n124, u1_u3_u7_n125, u1_u3_u7_n126, u1_u3_u7_n127, 
       u1_u3_u7_n128, u1_u3_u7_n129, u1_u3_u7_n130, u1_u3_u7_n131, u1_u3_u7_n132, u1_u3_u7_n133, u1_u3_u7_n134, u1_u3_u7_n135, u1_u3_u7_n136, 
       u1_u3_u7_n137, u1_u3_u7_n138, u1_u3_u7_n139, u1_u3_u7_n140, u1_u3_u7_n141, u1_u3_u7_n142, u1_u3_u7_n143, u1_u3_u7_n144, u1_u3_u7_n145, 
       u1_u3_u7_n146, u1_u3_u7_n147, u1_u3_u7_n148, u1_u3_u7_n149, u1_u3_u7_n150, u1_u3_u7_n151, u1_u3_u7_n152, u1_u3_u7_n153, u1_u3_u7_n154, 
       u1_u3_u7_n155, u1_u3_u7_n156, u1_u3_u7_n157, u1_u3_u7_n158, u1_u3_u7_n159, u1_u3_u7_n160, u1_u3_u7_n161, u1_u3_u7_n162, u1_u3_u7_n163, 
       u1_u3_u7_n164, u1_u3_u7_n165, u1_u3_u7_n166, u1_u3_u7_n167, u1_u3_u7_n168, u1_u3_u7_n169, u1_u3_u7_n170, u1_u3_u7_n171, u1_u3_u7_n172, 
       u1_u3_u7_n173, u1_u3_u7_n174, u1_u3_u7_n175, u1_u3_u7_n176, u1_u3_u7_n177, u1_u3_u7_n178, u1_u3_u7_n179, u1_u3_u7_n180, u1_u3_u7_n91, 
       u1_u3_u7_n92, u1_u3_u7_n93, u1_u3_u7_n94, u1_u3_u7_n95, u1_u3_u7_n96, u1_u3_u7_n97, u1_u3_u7_n98, u1_u3_u7_n99, u1_u4_X_10, 
       u1_u4_X_9, u1_u4_u1_n100, u1_u4_u1_n101, u1_u4_u1_n102, u1_u4_u1_n103, u1_u4_u1_n104, u1_u4_u1_n105, u1_u4_u1_n106, u1_u4_u1_n107, 
       u1_u4_u1_n108, u1_u4_u1_n109, u1_u4_u1_n110, u1_u4_u1_n111, u1_u4_u1_n112, u1_u4_u1_n113, u1_u4_u1_n114, u1_u4_u1_n115, u1_u4_u1_n116, 
       u1_u4_u1_n117, u1_u4_u1_n118, u1_u4_u1_n119, u1_u4_u1_n120, u1_u4_u1_n121, u1_u4_u1_n122, u1_u4_u1_n123, u1_u4_u1_n124, u1_u4_u1_n125, 
       u1_u4_u1_n126, u1_u4_u1_n127, u1_u4_u1_n128, u1_u4_u1_n129, u1_u4_u1_n130, u1_u4_u1_n131, u1_u4_u1_n132, u1_u4_u1_n133, u1_u4_u1_n134, 
       u1_u4_u1_n135, u1_u4_u1_n136, u1_u4_u1_n137, u1_u4_u1_n138, u1_u4_u1_n139, u1_u4_u1_n140, u1_u4_u1_n141, u1_u4_u1_n142, u1_u4_u1_n143, 
       u1_u4_u1_n144, u1_u4_u1_n145, u1_u4_u1_n146, u1_u4_u1_n147, u1_u4_u1_n148, u1_u4_u1_n149, u1_u4_u1_n150, u1_u4_u1_n151, u1_u4_u1_n152, 
       u1_u4_u1_n153, u1_u4_u1_n154, u1_u4_u1_n155, u1_u4_u1_n156, u1_u4_u1_n157, u1_u4_u1_n158, u1_u4_u1_n159, u1_u4_u1_n160, u1_u4_u1_n161, 
       u1_u4_u1_n162, u1_u4_u1_n163, u1_u4_u1_n164, u1_u4_u1_n165, u1_u4_u1_n166, u1_u4_u1_n167, u1_u4_u1_n168, u1_u4_u1_n169, u1_u4_u1_n170, 
       u1_u4_u1_n171, u1_u4_u1_n172, u1_u4_u1_n173, u1_u4_u1_n174, u1_u4_u1_n175, u1_u4_u1_n176, u1_u4_u1_n177, u1_u4_u1_n178, u1_u4_u1_n179, 
       u1_u4_u1_n180, u1_u4_u1_n181, u1_u4_u1_n182, u1_u4_u1_n183, u1_u4_u1_n184, u1_u4_u1_n185, u1_u4_u1_n186, u1_u4_u1_n187, u1_u4_u1_n188, 
       u1_u4_u1_n95, u1_u4_u1_n96, u1_u4_u1_n97, u1_u4_u1_n98, u1_u4_u1_n99, u1_u5_X_1, u1_u5_X_10, u1_u5_X_2, u1_u5_X_21, 
       u1_u5_X_22, u1_u5_X_3, u1_u5_X_33, u1_u5_X_34, u1_u5_X_35, u1_u5_X_36, u1_u5_X_37, u1_u5_X_38, u1_u5_X_39, 
       u1_u5_X_4, u1_u5_X_40, u1_u5_X_41, u1_u5_X_42, u1_u5_X_43, u1_u5_X_44, u1_u5_X_45, u1_u5_X_46, u1_u5_X_47, 
       u1_u5_X_48, u1_u5_X_6, u1_u5_X_8, u1_u5_X_9, u1_u5_u0_n100, u1_u5_u0_n101, u1_u5_u0_n102, u1_u5_u0_n103, u1_u5_u0_n104, 
       u1_u5_u0_n105, u1_u5_u0_n106, u1_u5_u0_n107, u1_u5_u0_n108, u1_u5_u0_n109, u1_u5_u0_n110, u1_u5_u0_n111, u1_u5_u0_n112, u1_u5_u0_n113, 
       u1_u5_u0_n114, u1_u5_u0_n115, u1_u5_u0_n116, u1_u5_u0_n117, u1_u5_u0_n118, u1_u5_u0_n119, u1_u5_u0_n120, u1_u5_u0_n121, u1_u5_u0_n122, 
       u1_u5_u0_n123, u1_u5_u0_n124, u1_u5_u0_n125, u1_u5_u0_n126, u1_u5_u0_n127, u1_u5_u0_n128, u1_u5_u0_n129, u1_u5_u0_n130, u1_u5_u0_n131, 
       u1_u5_u0_n132, u1_u5_u0_n133, u1_u5_u0_n134, u1_u5_u0_n135, u1_u5_u0_n136, u1_u5_u0_n137, u1_u5_u0_n138, u1_u5_u0_n139, u1_u5_u0_n140, 
       u1_u5_u0_n141, u1_u5_u0_n142, u1_u5_u0_n143, u1_u5_u0_n144, u1_u5_u0_n145, u1_u5_u0_n146, u1_u5_u0_n147, u1_u5_u0_n148, u1_u5_u0_n149, 
       u1_u5_u0_n150, u1_u5_u0_n151, u1_u5_u0_n152, u1_u5_u0_n153, u1_u5_u0_n154, u1_u5_u0_n155, u1_u5_u0_n156, u1_u5_u0_n157, u1_u5_u0_n158, 
       u1_u5_u0_n159, u1_u5_u0_n160, u1_u5_u0_n161, u1_u5_u0_n162, u1_u5_u0_n163, u1_u5_u0_n164, u1_u5_u0_n165, u1_u5_u0_n166, u1_u5_u0_n167, 
       u1_u5_u0_n168, u1_u5_u0_n169, u1_u5_u0_n170, u1_u5_u0_n171, u1_u5_u0_n172, u1_u5_u0_n173, u1_u5_u0_n174, u1_u5_u0_n88, u1_u5_u0_n89, 
       u1_u5_u0_n90, u1_u5_u0_n91, u1_u5_u0_n92, u1_u5_u0_n93, u1_u5_u0_n94, u1_u5_u0_n95, u1_u5_u0_n96, u1_u5_u0_n97, u1_u5_u0_n98, 
       u1_u5_u0_n99, u1_u5_u1_n100, u1_u5_u1_n101, u1_u5_u1_n102, u1_u5_u1_n103, u1_u5_u1_n104, u1_u5_u1_n105, u1_u5_u1_n106, u1_u5_u1_n107, 
       u1_u5_u1_n108, u1_u5_u1_n109, u1_u5_u1_n110, u1_u5_u1_n111, u1_u5_u1_n112, u1_u5_u1_n113, u1_u5_u1_n114, u1_u5_u1_n115, u1_u5_u1_n116, 
       u1_u5_u1_n117, u1_u5_u1_n118, u1_u5_u1_n119, u1_u5_u1_n120, u1_u5_u1_n121, u1_u5_u1_n122, u1_u5_u1_n123, u1_u5_u1_n124, u1_u5_u1_n125, 
       u1_u5_u1_n126, u1_u5_u1_n127, u1_u5_u1_n128, u1_u5_u1_n129, u1_u5_u1_n130, u1_u5_u1_n131, u1_u5_u1_n132, u1_u5_u1_n133, u1_u5_u1_n134, 
       u1_u5_u1_n135, u1_u5_u1_n136, u1_u5_u1_n137, u1_u5_u1_n138, u1_u5_u1_n139, u1_u5_u1_n140, u1_u5_u1_n141, u1_u5_u1_n142, u1_u5_u1_n143, 
       u1_u5_u1_n144, u1_u5_u1_n145, u1_u5_u1_n146, u1_u5_u1_n147, u1_u5_u1_n148, u1_u5_u1_n149, u1_u5_u1_n150, u1_u5_u1_n151, u1_u5_u1_n152, 
       u1_u5_u1_n153, u1_u5_u1_n154, u1_u5_u1_n155, u1_u5_u1_n156, u1_u5_u1_n157, u1_u5_u1_n158, u1_u5_u1_n159, u1_u5_u1_n160, u1_u5_u1_n161, 
       u1_u5_u1_n162, u1_u5_u1_n163, u1_u5_u1_n164, u1_u5_u1_n165, u1_u5_u1_n166, u1_u5_u1_n167, u1_u5_u1_n168, u1_u5_u1_n169, u1_u5_u1_n170, 
       u1_u5_u1_n171, u1_u5_u1_n172, u1_u5_u1_n173, u1_u5_u1_n174, u1_u5_u1_n175, u1_u5_u1_n176, u1_u5_u1_n177, u1_u5_u1_n178, u1_u5_u1_n179, 
       u1_u5_u1_n180, u1_u5_u1_n181, u1_u5_u1_n182, u1_u5_u1_n183, u1_u5_u1_n184, u1_u5_u1_n185, u1_u5_u1_n186, u1_u5_u1_n187, u1_u5_u1_n188, 
       u1_u5_u1_n95, u1_u5_u1_n96, u1_u5_u1_n97, u1_u5_u1_n98, u1_u5_u1_n99, u1_u5_u3_n100, u1_u5_u3_n101, u1_u5_u3_n102, u1_u5_u3_n103, 
       u1_u5_u3_n104, u1_u5_u3_n105, u1_u5_u3_n106, u1_u5_u3_n107, u1_u5_u3_n108, u1_u5_u3_n109, u1_u5_u3_n110, u1_u5_u3_n111, u1_u5_u3_n112, 
       u1_u5_u3_n113, u1_u5_u3_n114, u1_u5_u3_n115, u1_u5_u3_n116, u1_u5_u3_n117, u1_u5_u3_n118, u1_u5_u3_n119, u1_u5_u3_n120, u1_u5_u3_n121, 
       u1_u5_u3_n122, u1_u5_u3_n123, u1_u5_u3_n124, u1_u5_u3_n125, u1_u5_u3_n126, u1_u5_u3_n127, u1_u5_u3_n128, u1_u5_u3_n129, u1_u5_u3_n130, 
       u1_u5_u3_n131, u1_u5_u3_n132, u1_u5_u3_n133, u1_u5_u3_n134, u1_u5_u3_n135, u1_u5_u3_n136, u1_u5_u3_n137, u1_u5_u3_n138, u1_u5_u3_n139, 
       u1_u5_u3_n140, u1_u5_u3_n141, u1_u5_u3_n142, u1_u5_u3_n143, u1_u5_u3_n144, u1_u5_u3_n145, u1_u5_u3_n146, u1_u5_u3_n147, u1_u5_u3_n148, 
       u1_u5_u3_n149, u1_u5_u3_n150, u1_u5_u3_n151, u1_u5_u3_n152, u1_u5_u3_n153, u1_u5_u3_n154, u1_u5_u3_n155, u1_u5_u3_n156, u1_u5_u3_n157, 
       u1_u5_u3_n158, u1_u5_u3_n159, u1_u5_u3_n160, u1_u5_u3_n161, u1_u5_u3_n162, u1_u5_u3_n163, u1_u5_u3_n164, u1_u5_u3_n165, u1_u5_u3_n166, 
       u1_u5_u3_n167, u1_u5_u3_n168, u1_u5_u3_n169, u1_u5_u3_n170, u1_u5_u3_n171, u1_u5_u3_n172, u1_u5_u3_n173, u1_u5_u3_n174, u1_u5_u3_n175, 
       u1_u5_u3_n176, u1_u5_u3_n177, u1_u5_u3_n178, u1_u5_u3_n179, u1_u5_u3_n180, u1_u5_u3_n181, u1_u5_u3_n182, u1_u5_u3_n183, u1_u5_u3_n184, 
       u1_u5_u3_n185, u1_u5_u3_n186, u1_u5_u3_n94, u1_u5_u3_n95, u1_u5_u3_n96, u1_u5_u3_n97, u1_u5_u3_n98, u1_u5_u3_n99, u1_u5_u5_n100, 
       u1_u5_u5_n101, u1_u5_u5_n102, u1_u5_u5_n103, u1_u5_u5_n104, u1_u5_u5_n105, u1_u5_u5_n106, u1_u5_u5_n107, u1_u5_u5_n108, u1_u5_u5_n109, 
       u1_u5_u5_n110, u1_u5_u5_n111, u1_u5_u5_n112, u1_u5_u5_n113, u1_u5_u5_n114, u1_u5_u5_n115, u1_u5_u5_n116, u1_u5_u5_n117, u1_u5_u5_n118, 
       u1_u5_u5_n119, u1_u5_u5_n120, u1_u5_u5_n121, u1_u5_u5_n122, u1_u5_u5_n123, u1_u5_u5_n124, u1_u5_u5_n125, u1_u5_u5_n126, u1_u5_u5_n127, 
       u1_u5_u5_n128, u1_u5_u5_n129, u1_u5_u5_n130, u1_u5_u5_n131, u1_u5_u5_n132, u1_u5_u5_n133, u1_u5_u5_n134, u1_u5_u5_n135, u1_u5_u5_n136, 
       u1_u5_u5_n137, u1_u5_u5_n138, u1_u5_u5_n139, u1_u5_u5_n140, u1_u5_u5_n141, u1_u5_u5_n142, u1_u5_u5_n143, u1_u5_u5_n144, u1_u5_u5_n145, 
       u1_u5_u5_n146, u1_u5_u5_n147, u1_u5_u5_n148, u1_u5_u5_n149, u1_u5_u5_n150, u1_u5_u5_n151, u1_u5_u5_n152, u1_u5_u5_n153, u1_u5_u5_n154, 
       u1_u5_u5_n155, u1_u5_u5_n156, u1_u5_u5_n157, u1_u5_u5_n158, u1_u5_u5_n159, u1_u5_u5_n160, u1_u5_u5_n161, u1_u5_u5_n162, u1_u5_u5_n163, 
       u1_u5_u5_n164, u1_u5_u5_n165, u1_u5_u5_n166, u1_u5_u5_n167, u1_u5_u5_n168, u1_u5_u5_n169, u1_u5_u5_n170, u1_u5_u5_n171, u1_u5_u5_n172, 
       u1_u5_u5_n173, u1_u5_u5_n174, u1_u5_u5_n175, u1_u5_u5_n176, u1_u5_u5_n177, u1_u5_u5_n178, u1_u5_u5_n179, u1_u5_u5_n180, u1_u5_u5_n181, 
       u1_u5_u5_n182, u1_u5_u5_n183, u1_u5_u5_n184, u1_u5_u5_n185, u1_u5_u5_n186, u1_u5_u5_n187, u1_u5_u5_n188, u1_u5_u5_n189, u1_u5_u5_n190, 
       u1_u5_u5_n191, u1_u5_u5_n192, u1_u5_u5_n193, u1_u5_u5_n194, u1_u5_u5_n195, u1_u5_u5_n196, u1_u5_u5_n99, u1_u5_u6_n100, u1_u5_u6_n101, 
       u1_u5_u6_n102, u1_u5_u6_n103, u1_u5_u6_n104, u1_u5_u6_n105, u1_u5_u6_n106, u1_u5_u6_n107, u1_u5_u6_n108, u1_u5_u6_n109, u1_u5_u6_n110, 
       u1_u5_u6_n111, u1_u5_u6_n112, u1_u5_u6_n113, u1_u5_u6_n114, u1_u5_u6_n115, u1_u5_u6_n116, u1_u5_u6_n117, u1_u5_u6_n118, u1_u5_u6_n119, 
       u1_u5_u6_n120, u1_u5_u6_n121, u1_u5_u6_n122, u1_u5_u6_n123, u1_u5_u6_n124, u1_u5_u6_n125, u1_u5_u6_n126, u1_u5_u6_n127, u1_u5_u6_n128, 
       u1_u5_u6_n129, u1_u5_u6_n130, u1_u5_u6_n131, u1_u5_u6_n132, u1_u5_u6_n133, u1_u5_u6_n134, u1_u5_u6_n135, u1_u5_u6_n136, u1_u5_u6_n137, 
       u1_u5_u6_n138, u1_u5_u6_n139, u1_u5_u6_n140, u1_u5_u6_n141, u1_u5_u6_n142, u1_u5_u6_n143, u1_u5_u6_n144, u1_u5_u6_n145, u1_u5_u6_n146, 
       u1_u5_u6_n147, u1_u5_u6_n148, u1_u5_u6_n149, u1_u5_u6_n150, u1_u5_u6_n151, u1_u5_u6_n152, u1_u5_u6_n153, u1_u5_u6_n154, u1_u5_u6_n155, 
       u1_u5_u6_n156, u1_u5_u6_n157, u1_u5_u6_n158, u1_u5_u6_n159, u1_u5_u6_n160, u1_u5_u6_n161, u1_u5_u6_n162, u1_u5_u6_n163, u1_u5_u6_n164, 
       u1_u5_u6_n165, u1_u5_u6_n166, u1_u5_u6_n167, u1_u5_u6_n168, u1_u5_u6_n169, u1_u5_u6_n170, u1_u5_u6_n171, u1_u5_u6_n172, u1_u5_u6_n173, 
       u1_u5_u6_n174, u1_u5_u6_n88, u1_u5_u6_n89, u1_u5_u6_n90, u1_u5_u6_n91, u1_u5_u6_n92, u1_u5_u6_n93, u1_u5_u6_n94, u1_u5_u6_n95, 
       u1_u5_u6_n96, u1_u5_u6_n97, u1_u5_u6_n98, u1_u5_u6_n99, u1_u5_u7_n100, u1_u5_u7_n101, u1_u5_u7_n102, u1_u5_u7_n103, u1_u5_u7_n104, 
       u1_u5_u7_n105, u1_u5_u7_n106, u1_u5_u7_n107, u1_u5_u7_n108, u1_u5_u7_n109, u1_u5_u7_n110, u1_u5_u7_n111, u1_u5_u7_n112, u1_u5_u7_n113, 
       u1_u5_u7_n114, u1_u5_u7_n115, u1_u5_u7_n116, u1_u5_u7_n117, u1_u5_u7_n118, u1_u5_u7_n119, u1_u5_u7_n120, u1_u5_u7_n121, u1_u5_u7_n122, 
       u1_u5_u7_n123, u1_u5_u7_n124, u1_u5_u7_n125, u1_u5_u7_n126, u1_u5_u7_n127, u1_u5_u7_n128, u1_u5_u7_n129, u1_u5_u7_n130, u1_u5_u7_n131, 
       u1_u5_u7_n132, u1_u5_u7_n133, u1_u5_u7_n134, u1_u5_u7_n135, u1_u5_u7_n136, u1_u5_u7_n137, u1_u5_u7_n138, u1_u5_u7_n139, u1_u5_u7_n140, 
       u1_u5_u7_n141, u1_u5_u7_n142, u1_u5_u7_n143, u1_u5_u7_n144, u1_u5_u7_n145, u1_u5_u7_n146, u1_u5_u7_n147, u1_u5_u7_n148, u1_u5_u7_n149, 
       u1_u5_u7_n150, u1_u5_u7_n151, u1_u5_u7_n152, u1_u5_u7_n153, u1_u5_u7_n154, u1_u5_u7_n155, u1_u5_u7_n156, u1_u5_u7_n157, u1_u5_u7_n158, 
       u1_u5_u7_n159, u1_u5_u7_n160, u1_u5_u7_n161, u1_u5_u7_n162, u1_u5_u7_n163, u1_u5_u7_n164, u1_u5_u7_n165, u1_u5_u7_n166, u1_u5_u7_n167, 
       u1_u5_u7_n168, u1_u5_u7_n169, u1_u5_u7_n170, u1_u5_u7_n171, u1_u5_u7_n172, u1_u5_u7_n173, u1_u5_u7_n174, u1_u5_u7_n175, u1_u5_u7_n176, 
       u1_u5_u7_n177, u1_u5_u7_n178, u1_u5_u7_n179, u1_u5_u7_n180, u1_u5_u7_n91, u1_u5_u7_n92, u1_u5_u7_n93, u1_u5_u7_n94, u1_u5_u7_n95, 
       u1_u5_u7_n96, u1_u5_u7_n97, u1_u5_u7_n98, u1_u5_u7_n99, u1_u7_X_45, u1_u7_X_46, u1_u7_u7_n100, u1_u7_u7_n101, u1_u7_u7_n102, 
       u1_u7_u7_n103, u1_u7_u7_n104, u1_u7_u7_n105, u1_u7_u7_n106, u1_u7_u7_n107, u1_u7_u7_n108, u1_u7_u7_n109, u1_u7_u7_n110, u1_u7_u7_n111, 
       u1_u7_u7_n112, u1_u7_u7_n113, u1_u7_u7_n114, u1_u7_u7_n115, u1_u7_u7_n116, u1_u7_u7_n117, u1_u7_u7_n118, u1_u7_u7_n119, u1_u7_u7_n120, 
       u1_u7_u7_n121, u1_u7_u7_n122, u1_u7_u7_n123, u1_u7_u7_n124, u1_u7_u7_n125, u1_u7_u7_n126, u1_u7_u7_n127, u1_u7_u7_n128, u1_u7_u7_n129, 
       u1_u7_u7_n130, u1_u7_u7_n131, u1_u7_u7_n132, u1_u7_u7_n133, u1_u7_u7_n134, u1_u7_u7_n135, u1_u7_u7_n136, u1_u7_u7_n137, u1_u7_u7_n138, 
       u1_u7_u7_n139, u1_u7_u7_n140, u1_u7_u7_n141, u1_u7_u7_n142, u1_u7_u7_n143, u1_u7_u7_n144, u1_u7_u7_n145, u1_u7_u7_n146, u1_u7_u7_n147, 
       u1_u7_u7_n148, u1_u7_u7_n149, u1_u7_u7_n150, u1_u7_u7_n151, u1_u7_u7_n152, u1_u7_u7_n153, u1_u7_u7_n154, u1_u7_u7_n155, u1_u7_u7_n156, 
       u1_u7_u7_n157, u1_u7_u7_n158, u1_u7_u7_n159, u1_u7_u7_n160, u1_u7_u7_n161, u1_u7_u7_n162, u1_u7_u7_n163, u1_u7_u7_n164, u1_u7_u7_n165, 
       u1_u7_u7_n166, u1_u7_u7_n167, u1_u7_u7_n168, u1_u7_u7_n169, u1_u7_u7_n170, u1_u7_u7_n171, u1_u7_u7_n172, u1_u7_u7_n173, u1_u7_u7_n174, 
       u1_u7_u7_n175, u1_u7_u7_n176, u1_u7_u7_n177, u1_u7_u7_n178, u1_u7_u7_n179, u1_u7_u7_n180, u1_u7_u7_n91, u1_u7_u7_n92, u1_u7_u7_n93, 
       u1_u7_u7_n94, u1_u7_u7_n95, u1_u7_u7_n96, u1_u7_u7_n97, u1_u7_u7_n98, u1_u7_u7_n99, u1_u8_X_10, u1_u8_X_11, u1_u8_X_9, 
       u1_u8_u1_n100, u1_u8_u1_n101, u1_u8_u1_n102, u1_u8_u1_n103, u1_u8_u1_n104, u1_u8_u1_n105, u1_u8_u1_n106, u1_u8_u1_n107, u1_u8_u1_n108, 
       u1_u8_u1_n109, u1_u8_u1_n110, u1_u8_u1_n111, u1_u8_u1_n112, u1_u8_u1_n113, u1_u8_u1_n114, u1_u8_u1_n115, u1_u8_u1_n116, u1_u8_u1_n117, 
       u1_u8_u1_n118, u1_u8_u1_n119, u1_u8_u1_n120, u1_u8_u1_n121, u1_u8_u1_n122, u1_u8_u1_n123, u1_u8_u1_n124, u1_u8_u1_n125, u1_u8_u1_n126, 
       u1_u8_u1_n127, u1_u8_u1_n128, u1_u8_u1_n129, u1_u8_u1_n130, u1_u8_u1_n131, u1_u8_u1_n132, u1_u8_u1_n133, u1_u8_u1_n134, u1_u8_u1_n135, 
       u1_u8_u1_n136, u1_u8_u1_n137, u1_u8_u1_n138, u1_u8_u1_n139, u1_u8_u1_n140, u1_u8_u1_n141, u1_u8_u1_n142, u1_u8_u1_n143, u1_u8_u1_n144, 
       u1_u8_u1_n145, u1_u8_u1_n146, u1_u8_u1_n147, u1_u8_u1_n148, u1_u8_u1_n149, u1_u8_u1_n150, u1_u8_u1_n151, u1_u8_u1_n152, u1_u8_u1_n153, 
       u1_u8_u1_n154, u1_u8_u1_n155, u1_u8_u1_n156, u1_u8_u1_n157, u1_u8_u1_n158, u1_u8_u1_n159, u1_u8_u1_n160, u1_u8_u1_n161, u1_u8_u1_n162, 
       u1_u8_u1_n163, u1_u8_u1_n164, u1_u8_u1_n165, u1_u8_u1_n166, u1_u8_u1_n167, u1_u8_u1_n168, u1_u8_u1_n169, u1_u8_u1_n170, u1_u8_u1_n171, 
       u1_u8_u1_n172, u1_u8_u1_n173, u1_u8_u1_n174, u1_u8_u1_n175, u1_u8_u1_n176, u1_u8_u1_n177, u1_u8_u1_n178, u1_u8_u1_n179, u1_u8_u1_n180, 
       u1_u8_u1_n181, u1_u8_u1_n182, u1_u8_u1_n183, u1_u8_u1_n184, u1_u8_u1_n185, u1_u8_u1_n186, u1_u8_u1_n187, u1_u8_u1_n188, u1_u8_u1_n95, 
       u1_u8_u1_n96, u1_u8_u1_n97, u1_u8_u1_n98, u1_u8_u1_n99, u1_u9_X_15, u1_u9_X_16, u1_u9_X_17, u1_u9_X_18, u1_u9_X_19, 
       u1_u9_X_20, u1_u9_X_21, u1_u9_X_22, u1_u9_X_45, u1_u9_X_46, u1_u9_u2_n100, u1_u9_u2_n101, u1_u9_u2_n102, u1_u9_u2_n103, 
       u1_u9_u2_n104, u1_u9_u2_n105, u1_u9_u2_n106, u1_u9_u2_n107, u1_u9_u2_n108, u1_u9_u2_n109, u1_u9_u2_n110, u1_u9_u2_n111, u1_u9_u2_n112, 
       u1_u9_u2_n113, u1_u9_u2_n114, u1_u9_u2_n115, u1_u9_u2_n116, u1_u9_u2_n117, u1_u9_u2_n118, u1_u9_u2_n119, u1_u9_u2_n120, u1_u9_u2_n121, 
       u1_u9_u2_n122, u1_u9_u2_n123, u1_u9_u2_n124, u1_u9_u2_n125, u1_u9_u2_n126, u1_u9_u2_n127, u1_u9_u2_n128, u1_u9_u2_n129, u1_u9_u2_n130, 
       u1_u9_u2_n131, u1_u9_u2_n132, u1_u9_u2_n133, u1_u9_u2_n134, u1_u9_u2_n135, u1_u9_u2_n136, u1_u9_u2_n137, u1_u9_u2_n138, u1_u9_u2_n139, 
       u1_u9_u2_n140, u1_u9_u2_n141, u1_u9_u2_n142, u1_u9_u2_n143, u1_u9_u2_n144, u1_u9_u2_n145, u1_u9_u2_n146, u1_u9_u2_n147, u1_u9_u2_n148, 
       u1_u9_u2_n149, u1_u9_u2_n150, u1_u9_u2_n151, u1_u9_u2_n152, u1_u9_u2_n153, u1_u9_u2_n154, u1_u9_u2_n155, u1_u9_u2_n156, u1_u9_u2_n157, 
       u1_u9_u2_n158, u1_u9_u2_n159, u1_u9_u2_n160, u1_u9_u2_n161, u1_u9_u2_n162, u1_u9_u2_n163, u1_u9_u2_n164, u1_u9_u2_n165, u1_u9_u2_n166, 
       u1_u9_u2_n167, u1_u9_u2_n168, u1_u9_u2_n169, u1_u9_u2_n170, u1_u9_u2_n171, u1_u9_u2_n172, u1_u9_u2_n173, u1_u9_u2_n174, u1_u9_u2_n175, 
       u1_u9_u2_n176, u1_u9_u2_n177, u1_u9_u2_n178, u1_u9_u2_n179, u1_u9_u2_n180, u1_u9_u2_n181, u1_u9_u2_n182, u1_u9_u2_n183, u1_u9_u2_n184, 
       u1_u9_u2_n185, u1_u9_u2_n186, u1_u9_u2_n187, u1_u9_u2_n188, u1_u9_u2_n95, u1_u9_u2_n96, u1_u9_u2_n97, u1_u9_u2_n98, u1_u9_u2_n99, 
       u1_u9_u3_n100, u1_u9_u3_n101, u1_u9_u3_n102, u1_u9_u3_n103, u1_u9_u3_n104, u1_u9_u3_n105, u1_u9_u3_n106, u1_u9_u3_n107, u1_u9_u3_n108, 
       u1_u9_u3_n109, u1_u9_u3_n110, u1_u9_u3_n111, u1_u9_u3_n112, u1_u9_u3_n113, u1_u9_u3_n114, u1_u9_u3_n115, u1_u9_u3_n116, u1_u9_u3_n117, 
       u1_u9_u3_n118, u1_u9_u3_n119, u1_u9_u3_n120, u1_u9_u3_n121, u1_u9_u3_n122, u1_u9_u3_n123, u1_u9_u3_n124, u1_u9_u3_n125, u1_u9_u3_n126, 
       u1_u9_u3_n127, u1_u9_u3_n128, u1_u9_u3_n129, u1_u9_u3_n130, u1_u9_u3_n131, u1_u9_u3_n132, u1_u9_u3_n133, u1_u9_u3_n134, u1_u9_u3_n135, 
       u1_u9_u3_n136, u1_u9_u3_n137, u1_u9_u3_n138, u1_u9_u3_n139, u1_u9_u3_n140, u1_u9_u3_n141, u1_u9_u3_n142, u1_u9_u3_n143, u1_u9_u3_n144, 
       u1_u9_u3_n145, u1_u9_u3_n146, u1_u9_u3_n147, u1_u9_u3_n148, u1_u9_u3_n149, u1_u9_u3_n150, u1_u9_u3_n151, u1_u9_u3_n152, u1_u9_u3_n153, 
       u1_u9_u3_n154, u1_u9_u3_n155, u1_u9_u3_n156, u1_u9_u3_n157, u1_u9_u3_n158, u1_u9_u3_n159, u1_u9_u3_n160, u1_u9_u3_n161, u1_u9_u3_n162, 
       u1_u9_u3_n163, u1_u9_u3_n164, u1_u9_u3_n165, u1_u9_u3_n166, u1_u9_u3_n167, u1_u9_u3_n168, u1_u9_u3_n169, u1_u9_u3_n170, u1_u9_u3_n171, 
       u1_u9_u3_n172, u1_u9_u3_n173, u1_u9_u3_n174, u1_u9_u3_n175, u1_u9_u3_n176, u1_u9_u3_n177, u1_u9_u3_n178, u1_u9_u3_n179, u1_u9_u3_n180, 
       u1_u9_u3_n181, u1_u9_u3_n182, u1_u9_u3_n183, u1_u9_u3_n184, u1_u9_u3_n185, u1_u9_u3_n186, u1_u9_u3_n94, u1_u9_u3_n95, u1_u9_u3_n96, 
       u1_u9_u3_n97, u1_u9_u3_n98, u1_u9_u3_n99, u1_u9_u7_n100, u1_u9_u7_n101, u1_u9_u7_n102, u1_u9_u7_n103, u1_u9_u7_n104, u1_u9_u7_n105, 
       u1_u9_u7_n106, u1_u9_u7_n107, u1_u9_u7_n108, u1_u9_u7_n109, u1_u9_u7_n110, u1_u9_u7_n111, u1_u9_u7_n112, u1_u9_u7_n113, u1_u9_u7_n114, 
       u1_u9_u7_n115, u1_u9_u7_n116, u1_u9_u7_n117, u1_u9_u7_n118, u1_u9_u7_n119, u1_u9_u7_n120, u1_u9_u7_n121, u1_u9_u7_n122, u1_u9_u7_n123, 
       u1_u9_u7_n124, u1_u9_u7_n125, u1_u9_u7_n126, u1_u9_u7_n127, u1_u9_u7_n128, u1_u9_u7_n129, u1_u9_u7_n130, u1_u9_u7_n131, u1_u9_u7_n132, 
       u1_u9_u7_n133, u1_u9_u7_n134, u1_u9_u7_n135, u1_u9_u7_n136, u1_u9_u7_n137, u1_u9_u7_n138, u1_u9_u7_n139, u1_u9_u7_n140, u1_u9_u7_n141, 
       u1_u9_u7_n142, u1_u9_u7_n143, u1_u9_u7_n144, u1_u9_u7_n145, u1_u9_u7_n146, u1_u9_u7_n147, u1_u9_u7_n148, u1_u9_u7_n149, u1_u9_u7_n150, 
       u1_u9_u7_n151, u1_u9_u7_n152, u1_u9_u7_n153, u1_u9_u7_n154, u1_u9_u7_n155, u1_u9_u7_n156, u1_u9_u7_n157, u1_u9_u7_n158, u1_u9_u7_n159, 
       u1_u9_u7_n160, u1_u9_u7_n161, u1_u9_u7_n162, u1_u9_u7_n163, u1_u9_u7_n164, u1_u9_u7_n165, u1_u9_u7_n166, u1_u9_u7_n167, u1_u9_u7_n168, 
       u1_u9_u7_n169, u1_u9_u7_n170, u1_u9_u7_n171, u1_u9_u7_n172, u1_u9_u7_n173, u1_u9_u7_n174, u1_u9_u7_n175, u1_u9_u7_n176, u1_u9_u7_n177, 
       u1_u9_u7_n178, u1_u9_u7_n179, u1_u9_u7_n180, u1_u9_u7_n91, u1_u9_u7_n92, u1_u9_u7_n93, u1_u9_u7_n94, u1_u9_u7_n95, u1_u9_u7_n96, 
       u1_u9_u7_n97, u1_u9_u7_n98, u1_u9_u7_n99, u2_K10_31, u2_K10_33, u2_K10_35, u2_K15_26, u2_K15_27, u2_K15_33, 
       u2_K15_36, u2_K1_25, u2_K1_26, u2_K1_27, u2_K1_29, u2_K1_31, u2_K1_32, u2_K1_33, u2_K1_35, 
       u2_K1_36, u2_K1_38, u2_K1_39, u2_K1_41, u2_K1_42, u2_K1_44, u2_K1_47, u2_K1_48, u2_u0_X_25, 
       u2_u0_X_26, u2_u0_X_27, u2_u0_X_29, u2_u0_X_30, u2_u0_X_31, u2_u0_X_32, u2_u0_X_33, u2_u0_X_35, u2_u0_X_36, 
       u2_u0_X_37, u2_u0_X_38, u2_u0_X_39, u2_u0_X_41, u2_u0_X_42, u2_u0_X_43, u2_u0_X_44, u2_u0_X_47, u2_u0_X_48, 
       u2_u0_u4_n100, u2_u0_u4_n101, u2_u0_u4_n102, u2_u0_u4_n103, u2_u0_u4_n104, u2_u0_u4_n105, u2_u0_u4_n106, u2_u0_u4_n107, u2_u0_u4_n108, 
       u2_u0_u4_n109, u2_u0_u4_n110, u2_u0_u4_n111, u2_u0_u4_n112, u2_u0_u4_n113, u2_u0_u4_n114, u2_u0_u4_n115, u2_u0_u4_n116, u2_u0_u4_n117, 
       u2_u0_u4_n118, u2_u0_u4_n119, u2_u0_u4_n120, u2_u0_u4_n121, u2_u0_u4_n122, u2_u0_u4_n123, u2_u0_u4_n124, u2_u0_u4_n125, u2_u0_u4_n126, 
       u2_u0_u4_n127, u2_u0_u4_n128, u2_u0_u4_n129, u2_u0_u4_n130, u2_u0_u4_n131, u2_u0_u4_n132, u2_u0_u4_n133, u2_u0_u4_n134, u2_u0_u4_n135, 
       u2_u0_u4_n136, u2_u0_u4_n137, u2_u0_u4_n138, u2_u0_u4_n139, u2_u0_u4_n140, u2_u0_u4_n141, u2_u0_u4_n142, u2_u0_u4_n143, u2_u0_u4_n144, 
       u2_u0_u4_n145, u2_u0_u4_n146, u2_u0_u4_n147, u2_u0_u4_n148, u2_u0_u4_n149, u2_u0_u4_n150, u2_u0_u4_n151, u2_u0_u4_n152, u2_u0_u4_n153, 
       u2_u0_u4_n154, u2_u0_u4_n155, u2_u0_u4_n156, u2_u0_u4_n157, u2_u0_u4_n158, u2_u0_u4_n159, u2_u0_u4_n160, u2_u0_u4_n161, u2_u0_u4_n162, 
       u2_u0_u4_n163, u2_u0_u4_n164, u2_u0_u4_n165, u2_u0_u4_n166, u2_u0_u4_n167, u2_u0_u4_n168, u2_u0_u4_n169, u2_u0_u4_n170, u2_u0_u4_n171, 
       u2_u0_u4_n172, u2_u0_u4_n173, u2_u0_u4_n174, u2_u0_u4_n175, u2_u0_u4_n176, u2_u0_u4_n177, u2_u0_u4_n178, u2_u0_u4_n179, u2_u0_u4_n180, 
       u2_u0_u4_n181, u2_u0_u4_n182, u2_u0_u4_n183, u2_u0_u4_n184, u2_u0_u4_n185, u2_u0_u4_n186, u2_u0_u4_n94, u2_u0_u4_n95, u2_u0_u4_n96, 
       u2_u0_u4_n97, u2_u0_u4_n98, u2_u0_u4_n99, u2_u0_u5_n100, u2_u0_u5_n101, u2_u0_u5_n102, u2_u0_u5_n103, u2_u0_u5_n104, u2_u0_u5_n105, 
       u2_u0_u5_n106, u2_u0_u5_n107, u2_u0_u5_n108, u2_u0_u5_n109, u2_u0_u5_n110, u2_u0_u5_n111, u2_u0_u5_n112, u2_u0_u5_n113, u2_u0_u5_n114, 
       u2_u0_u5_n115, u2_u0_u5_n116, u2_u0_u5_n117, u2_u0_u5_n118, u2_u0_u5_n119, u2_u0_u5_n120, u2_u0_u5_n121, u2_u0_u5_n122, u2_u0_u5_n123, 
       u2_u0_u5_n124, u2_u0_u5_n125, u2_u0_u5_n126, u2_u0_u5_n127, u2_u0_u5_n128, u2_u0_u5_n129, u2_u0_u5_n130, u2_u0_u5_n131, u2_u0_u5_n132, 
       u2_u0_u5_n133, u2_u0_u5_n134, u2_u0_u5_n135, u2_u0_u5_n136, u2_u0_u5_n137, u2_u0_u5_n138, u2_u0_u5_n139, u2_u0_u5_n140, u2_u0_u5_n141, 
       u2_u0_u5_n142, u2_u0_u5_n143, u2_u0_u5_n144, u2_u0_u5_n145, u2_u0_u5_n146, u2_u0_u5_n147, u2_u0_u5_n148, u2_u0_u5_n149, u2_u0_u5_n150, 
       u2_u0_u5_n151, u2_u0_u5_n152, u2_u0_u5_n153, u2_u0_u5_n154, u2_u0_u5_n155, u2_u0_u5_n156, u2_u0_u5_n157, u2_u0_u5_n158, u2_u0_u5_n159, 
       u2_u0_u5_n160, u2_u0_u5_n161, u2_u0_u5_n162, u2_u0_u5_n163, u2_u0_u5_n164, u2_u0_u5_n165, u2_u0_u5_n166, u2_u0_u5_n167, u2_u0_u5_n168, 
       u2_u0_u5_n169, u2_u0_u5_n170, u2_u0_u5_n171, u2_u0_u5_n172, u2_u0_u5_n173, u2_u0_u5_n174, u2_u0_u5_n175, u2_u0_u5_n176, u2_u0_u5_n177, 
       u2_u0_u5_n178, u2_u0_u5_n179, u2_u0_u5_n180, u2_u0_u5_n181, u2_u0_u5_n182, u2_u0_u5_n183, u2_u0_u5_n184, u2_u0_u5_n185, u2_u0_u5_n186, 
       u2_u0_u5_n187, u2_u0_u5_n188, u2_u0_u5_n189, u2_u0_u5_n190, u2_u0_u5_n191, u2_u0_u5_n192, u2_u0_u5_n193, u2_u0_u5_n194, u2_u0_u5_n195, 
       u2_u0_u5_n196, u2_u0_u5_n99, u2_u0_u6_n100, u2_u0_u6_n101, u2_u0_u6_n102, u2_u0_u6_n103, u2_u0_u6_n104, u2_u0_u6_n105, u2_u0_u6_n106, 
       u2_u0_u6_n107, u2_u0_u6_n108, u2_u0_u6_n109, u2_u0_u6_n110, u2_u0_u6_n111, u2_u0_u6_n112, u2_u0_u6_n113, u2_u0_u6_n114, u2_u0_u6_n115, 
       u2_u0_u6_n116, u2_u0_u6_n117, u2_u0_u6_n118, u2_u0_u6_n119, u2_u0_u6_n120, u2_u0_u6_n121, u2_u0_u6_n122, u2_u0_u6_n123, u2_u0_u6_n124, 
       u2_u0_u6_n125, u2_u0_u6_n126, u2_u0_u6_n127, u2_u0_u6_n128, u2_u0_u6_n129, u2_u0_u6_n130, u2_u0_u6_n131, u2_u0_u6_n132, u2_u0_u6_n133, 
       u2_u0_u6_n134, u2_u0_u6_n135, u2_u0_u6_n136, u2_u0_u6_n137, u2_u0_u6_n138, u2_u0_u6_n139, u2_u0_u6_n140, u2_u0_u6_n141, u2_u0_u6_n142, 
       u2_u0_u6_n143, u2_u0_u6_n144, u2_u0_u6_n145, u2_u0_u6_n146, u2_u0_u6_n147, u2_u0_u6_n148, u2_u0_u6_n149, u2_u0_u6_n150, u2_u0_u6_n151, 
       u2_u0_u6_n152, u2_u0_u6_n153, u2_u0_u6_n154, u2_u0_u6_n155, u2_u0_u6_n156, u2_u0_u6_n157, u2_u0_u6_n158, u2_u0_u6_n159, u2_u0_u6_n160, 
       u2_u0_u6_n161, u2_u0_u6_n162, u2_u0_u6_n163, u2_u0_u6_n164, u2_u0_u6_n165, u2_u0_u6_n166, u2_u0_u6_n167, u2_u0_u6_n168, u2_u0_u6_n169, 
       u2_u0_u6_n170, u2_u0_u6_n171, u2_u0_u6_n172, u2_u0_u6_n173, u2_u0_u6_n174, u2_u0_u6_n88, u2_u0_u6_n89, u2_u0_u6_n90, u2_u0_u6_n91, 
       u2_u0_u6_n92, u2_u0_u6_n93, u2_u0_u6_n94, u2_u0_u6_n95, u2_u0_u6_n96, u2_u0_u6_n97, u2_u0_u6_n98, u2_u0_u6_n99, u2_u0_u7_n100, 
       u2_u0_u7_n101, u2_u0_u7_n102, u2_u0_u7_n103, u2_u0_u7_n104, u2_u0_u7_n105, u2_u0_u7_n106, u2_u0_u7_n107, u2_u0_u7_n108, u2_u0_u7_n109, 
       u2_u0_u7_n110, u2_u0_u7_n111, u2_u0_u7_n112, u2_u0_u7_n113, u2_u0_u7_n114, u2_u0_u7_n115, u2_u0_u7_n116, u2_u0_u7_n117, u2_u0_u7_n118, 
       u2_u0_u7_n119, u2_u0_u7_n120, u2_u0_u7_n121, u2_u0_u7_n122, u2_u0_u7_n123, u2_u0_u7_n124, u2_u0_u7_n125, u2_u0_u7_n126, u2_u0_u7_n127, 
       u2_u0_u7_n128, u2_u0_u7_n129, u2_u0_u7_n130, u2_u0_u7_n131, u2_u0_u7_n132, u2_u0_u7_n133, u2_u0_u7_n134, u2_u0_u7_n135, u2_u0_u7_n136, 
       u2_u0_u7_n137, u2_u0_u7_n138, u2_u0_u7_n139, u2_u0_u7_n140, u2_u0_u7_n141, u2_u0_u7_n142, u2_u0_u7_n143, u2_u0_u7_n144, u2_u0_u7_n145, 
       u2_u0_u7_n146, u2_u0_u7_n147, u2_u0_u7_n148, u2_u0_u7_n149, u2_u0_u7_n150, u2_u0_u7_n151, u2_u0_u7_n152, u2_u0_u7_n153, u2_u0_u7_n154, 
       u2_u0_u7_n155, u2_u0_u7_n156, u2_u0_u7_n157, u2_u0_u7_n158, u2_u0_u7_n159, u2_u0_u7_n160, u2_u0_u7_n161, u2_u0_u7_n162, u2_u0_u7_n163, 
       u2_u0_u7_n164, u2_u0_u7_n165, u2_u0_u7_n166, u2_u0_u7_n167, u2_u0_u7_n168, u2_u0_u7_n169, u2_u0_u7_n170, u2_u0_u7_n171, u2_u0_u7_n172, 
       u2_u0_u7_n173, u2_u0_u7_n174, u2_u0_u7_n175, u2_u0_u7_n176, u2_u0_u7_n177, u2_u0_u7_n178, u2_u0_u7_n179, u2_u0_u7_n180, u2_u0_u7_n91, 
       u2_u0_u7_n92, u2_u0_u7_n93, u2_u0_u7_n94, u2_u0_u7_n95, u2_u0_u7_n96, u2_u0_u7_n97, u2_u0_u7_n98, u2_u0_u7_n99, u2_u14_X_26, 
       u2_u14_X_27, u2_u14_X_29, u2_u14_X_31, u2_u14_X_33, u2_u14_X_35, u2_u14_X_36, u2_u14_u4_n100, u2_u14_u4_n101, u2_u14_u4_n102, 
       u2_u14_u4_n103, u2_u14_u4_n104, u2_u14_u4_n105, u2_u14_u4_n106, u2_u14_u4_n107, u2_u14_u4_n108, u2_u14_u4_n109, u2_u14_u4_n110, u2_u14_u4_n111, 
       u2_u14_u4_n112, u2_u14_u4_n113, u2_u14_u4_n114, u2_u14_u4_n115, u2_u14_u4_n116, u2_u14_u4_n117, u2_u14_u4_n118, u2_u14_u4_n119, u2_u14_u4_n120, 
       u2_u14_u4_n121, u2_u14_u4_n122, u2_u14_u4_n123, u2_u14_u4_n124, u2_u14_u4_n125, u2_u14_u4_n126, u2_u14_u4_n127, u2_u14_u4_n128, u2_u14_u4_n129, 
       u2_u14_u4_n130, u2_u14_u4_n131, u2_u14_u4_n132, u2_u14_u4_n133, u2_u14_u4_n134, u2_u14_u4_n135, u2_u14_u4_n136, u2_u14_u4_n137, u2_u14_u4_n138, 
       u2_u14_u4_n139, u2_u14_u4_n140, u2_u14_u4_n141, u2_u14_u4_n142, u2_u14_u4_n143, u2_u14_u4_n144, u2_u14_u4_n145, u2_u14_u4_n146, u2_u14_u4_n147, 
       u2_u14_u4_n148, u2_u14_u4_n149, u2_u14_u4_n150, u2_u14_u4_n151, u2_u14_u4_n152, u2_u14_u4_n153, u2_u14_u4_n154, u2_u14_u4_n155, u2_u14_u4_n156, 
       u2_u14_u4_n157, u2_u14_u4_n158, u2_u14_u4_n159, u2_u14_u4_n160, u2_u14_u4_n161, u2_u14_u4_n162, u2_u14_u4_n163, u2_u14_u4_n164, u2_u14_u4_n165, 
       u2_u14_u4_n166, u2_u14_u4_n167, u2_u14_u4_n168, u2_u14_u4_n169, u2_u14_u4_n170, u2_u14_u4_n171, u2_u14_u4_n172, u2_u14_u4_n173, u2_u14_u4_n174, 
       u2_u14_u4_n175, u2_u14_u4_n176, u2_u14_u4_n177, u2_u14_u4_n178, u2_u14_u4_n179, u2_u14_u4_n180, u2_u14_u4_n181, u2_u14_u4_n182, u2_u14_u4_n183, 
       u2_u14_u4_n184, u2_u14_u4_n185, u2_u14_u4_n186, u2_u14_u4_n94, u2_u14_u4_n95, u2_u14_u4_n96, u2_u14_u4_n97, u2_u14_u4_n98, u2_u14_u4_n99, 
       u2_u14_u5_n100, u2_u14_u5_n101, u2_u14_u5_n102, u2_u14_u5_n103, u2_u14_u5_n104, u2_u14_u5_n105, u2_u14_u5_n106, u2_u14_u5_n107, u2_u14_u5_n108, 
       u2_u14_u5_n109, u2_u14_u5_n110, u2_u14_u5_n111, u2_u14_u5_n112, u2_u14_u5_n113, u2_u14_u5_n114, u2_u14_u5_n115, u2_u14_u5_n116, u2_u14_u5_n117, 
       u2_u14_u5_n118, u2_u14_u5_n119, u2_u14_u5_n120, u2_u14_u5_n121, u2_u14_u5_n122, u2_u14_u5_n123, u2_u14_u5_n124, u2_u14_u5_n125, u2_u14_u5_n126, 
       u2_u14_u5_n127, u2_u14_u5_n128, u2_u14_u5_n129, u2_u14_u5_n130, u2_u14_u5_n131, u2_u14_u5_n132, u2_u14_u5_n133, u2_u14_u5_n134, u2_u14_u5_n135, 
       u2_u14_u5_n136, u2_u14_u5_n137, u2_u14_u5_n138, u2_u14_u5_n139, u2_u14_u5_n140, u2_u14_u5_n141, u2_u14_u5_n142, u2_u14_u5_n143, u2_u14_u5_n144, 
       u2_u14_u5_n145, u2_u14_u5_n146, u2_u14_u5_n147, u2_u14_u5_n148, u2_u14_u5_n149, u2_u14_u5_n150, u2_u14_u5_n151, u2_u14_u5_n152, u2_u14_u5_n153, 
       u2_u14_u5_n154, u2_u14_u5_n155, u2_u14_u5_n156, u2_u14_u5_n157, u2_u14_u5_n158, u2_u14_u5_n159, u2_u14_u5_n160, u2_u14_u5_n161, u2_u14_u5_n162, 
       u2_u14_u5_n163, u2_u14_u5_n164, u2_u14_u5_n165, u2_u14_u5_n166, u2_u14_u5_n167, u2_u14_u5_n168, u2_u14_u5_n169, u2_u14_u5_n170, u2_u14_u5_n171, 
       u2_u14_u5_n172, u2_u14_u5_n173, u2_u14_u5_n174, u2_u14_u5_n175, u2_u14_u5_n176, u2_u14_u5_n177, u2_u14_u5_n178, u2_u14_u5_n179, u2_u14_u5_n180, 
       u2_u14_u5_n181, u2_u14_u5_n182, u2_u14_u5_n183, u2_u14_u5_n184, u2_u14_u5_n185, u2_u14_u5_n186, u2_u14_u5_n187, u2_u14_u5_n188, u2_u14_u5_n189, 
       u2_u14_u5_n190, u2_u14_u5_n191, u2_u14_u5_n192, u2_u14_u5_n193, u2_u14_u5_n194, u2_u14_u5_n195, u2_u14_u5_n196, u2_u14_u5_n99, u2_u9_X_31, 
       u2_u9_X_33, u2_u9_X_35, u2_u9_X_36, u2_u9_u5_n100, u2_u9_u5_n101, u2_u9_u5_n102, u2_u9_u5_n103, u2_u9_u5_n104, u2_u9_u5_n105, 
       u2_u9_u5_n106, u2_u9_u5_n107, u2_u9_u5_n108, u2_u9_u5_n109, u2_u9_u5_n110, u2_u9_u5_n111, u2_u9_u5_n112, u2_u9_u5_n113, u2_u9_u5_n114, 
       u2_u9_u5_n115, u2_u9_u5_n116, u2_u9_u5_n117, u2_u9_u5_n118, u2_u9_u5_n119, u2_u9_u5_n120, u2_u9_u5_n121, u2_u9_u5_n122, u2_u9_u5_n123, 
       u2_u9_u5_n124, u2_u9_u5_n125, u2_u9_u5_n126, u2_u9_u5_n127, u2_u9_u5_n128, u2_u9_u5_n129, u2_u9_u5_n130, u2_u9_u5_n131, u2_u9_u5_n132, 
       u2_u9_u5_n133, u2_u9_u5_n134, u2_u9_u5_n135, u2_u9_u5_n136, u2_u9_u5_n137, u2_u9_u5_n138, u2_u9_u5_n139, u2_u9_u5_n140, u2_u9_u5_n141, 
       u2_u9_u5_n142, u2_u9_u5_n143, u2_u9_u5_n144, u2_u9_u5_n145, u2_u9_u5_n146, u2_u9_u5_n147, u2_u9_u5_n148, u2_u9_u5_n149, u2_u9_u5_n150, 
       u2_u9_u5_n151, u2_u9_u5_n152, u2_u9_u5_n153, u2_u9_u5_n154, u2_u9_u5_n155, u2_u9_u5_n156, u2_u9_u5_n157, u2_u9_u5_n158, u2_u9_u5_n159, 
       u2_u9_u5_n160, u2_u9_u5_n161, u2_u9_u5_n162, u2_u9_u5_n163, u2_u9_u5_n164, u2_u9_u5_n165, u2_u9_u5_n166, u2_u9_u5_n167, u2_u9_u5_n168, 
       u2_u9_u5_n169, u2_u9_u5_n170, u2_u9_u5_n171, u2_u9_u5_n172, u2_u9_u5_n173, u2_u9_u5_n174, u2_u9_u5_n175, u2_u9_u5_n176, u2_u9_u5_n177, 
       u2_u9_u5_n178, u2_u9_u5_n179, u2_u9_u5_n180, u2_u9_u5_n181, u2_u9_u5_n182, u2_u9_u5_n183, u2_u9_u5_n184, u2_u9_u5_n185, u2_u9_u5_n186, 
       u2_u9_u5_n187, u2_u9_u5_n188, u2_u9_u5_n189, u2_u9_u5_n190, u2_u9_u5_n191, u2_u9_u5_n192, u2_u9_u5_n193, u2_u9_u5_n194, u2_u9_u5_n195, 
       u2_u9_u5_n196, u2_u9_u5_n99, u2_uk_n1147, u2_uk_n1151, u2_uk_n1157, u2_uk_n1158, u2_uk_n1165, u2_uk_n291, u2_uk_n294, 
       u2_uk_n297, u2_uk_n975, u2_uk_n976, u2_uk_n977, u2_uk_n980, u2_uk_n981, u2_uk_n982, u2_uk_n985, u2_uk_n987, 
        u2_uk_n989;
  XOR2_X1 u0_u0_U11 (.B( u0_K1_44 ) , .A( u0_desIn_r_33 ) , .Z( u0_u0_X_44 ) );
  XOR2_X1 u0_u0_U12 (.B( u0_K1_43 ) , .A( u0_desIn_r_25 ) , .Z( u0_u0_X_43 ) );
  XOR2_X1 u0_u0_U13 (.B( u0_K1_42 ) , .A( u0_desIn_r_33 ) , .Z( u0_u0_X_42 ) );
  XOR2_X1 u0_u0_U14 (.B( u0_K1_41 ) , .A( u0_desIn_r_25 ) , .Z( u0_u0_X_41 ) );
  XOR2_X1 u0_u0_U18 (.B( u0_K1_38 ) , .A( u0_desIn_r_1 ) , .Z( u0_u0_X_38 ) );
  XOR2_X1 u0_u0_U19 (.B( u0_K1_37 ) , .A( u0_desIn_r_59 ) , .Z( u0_u0_X_37 ) );
  XOR2_X1 u0_u0_U20 (.B( u0_K1_36 ) , .A( u0_desIn_r_1 ) , .Z( u0_u0_X_36 ) );
  XOR2_X1 u0_u0_U21 (.B( u0_K1_35 ) , .A( u0_desIn_r_59 ) , .Z( u0_u0_X_35 ) );
  XOR2_X1 u0_u0_U22 (.B( u0_K1_34 ) , .A( u0_desIn_r_51 ) , .Z( u0_u0_X_34 ) );
  XOR2_X1 u0_u0_U25 (.B( u0_K1_31 ) , .A( u0_desIn_r_27 ) , .Z( u0_u0_X_31 ) );
  XOR2_X1 u0_u0_U28 (.B( u0_K1_29 ) , .A( u0_desIn_r_27 ) , .Z( u0_u0_X_29 ) );
  XOR2_X1 u0_u0_U30 (.B( u0_K1_27 ) , .A( u0_desIn_r_11 ) , .Z( u0_u0_X_27 ) );
  XOR2_X1 u0_u0_U31 (.B( u0_K1_26 ) , .A( u0_desIn_r_3 ) , .Z( u0_u0_X_26 ) );
  XOR2_X1 u0_u0_U7 (.B( u0_K1_48 ) , .A( u0_desIn_r_7 ) , .Z( u0_u0_X_48 ) );
  XOR2_X1 u0_u0_U8 (.B( u0_K1_47 ) , .A( u0_desIn_r_57 ) , .Z( u0_u0_X_47 ) );
  OAI22_X1 u0_u0_u4_U10 (.A2( u0_u0_u4_n16 ) , .A1( u0_u0_u4_n32 ) , .B1( u0_u0_u4_n34 ) , .ZN( u0_u0_u4_n50 ) , .B2( u0_u0_u4_n52 ) );
  AND3_X1 u0_u0_u4_U11 (.A1( u0_u0_u4_n30 ) , .A3( u0_u0_u4_n42 ) , .ZN( u0_u0_u4_n52 ) , .A2( u0_u0_u4_n53 ) );
  NAND2_X1 u0_u0_u4_U12 (.A1( u0_u0_u4_n14 ) , .A2( u0_u0_u4_n17 ) , .ZN( u0_u0_u4_n55 ) );
  AOI21_X1 u0_u0_u4_U13 (.A( u0_u0_u4_n17 ) , .ZN( u0_u0_u4_n25 ) , .B1( u0_u0_u4_n26 ) , .B2( u0_u0_u4_n27 ) );
  AOI21_X1 u0_u0_u4_U14 (.A( u0_u0_u4_n13 ) , .B1( u0_u0_u4_n3 ) , .B2( u0_u0_u4_n44 ) , .ZN( u0_u0_u4_n80 ) );
  AOI21_X1 u0_u0_u4_U15 (.A( u0_u0_u4_n13 ) , .ZN( u0_u0_u4_n24 ) , .B1( u0_u0_u4_n28 ) , .B2( u0_u0_u4_n29 ) );
  AOI21_X1 u0_u0_u4_U16 (.ZN( u0_u0_u4_n22 ) , .B1( u0_u0_u4_n32 ) , .B2( u0_u0_u4_n33 ) , .A( u0_u0_u4_n34 ) );
  AOI21_X1 u0_u0_u4_U17 (.ZN( u0_u0_u4_n23 ) , .B1( u0_u0_u4_n3 ) , .B2( u0_u0_u4_n30 ) , .A( u0_u0_u4_n31 ) );
  INV_X1 u0_u0_u4_U18 (.ZN( u0_u0_u4_n17 ) , .A( u0_u0_u4_n49 ) );
  AND2_X1 u0_u0_u4_U19 (.A1( u0_u0_u4_n27 ) , .ZN( u0_u0_u4_n32 ) , .A2( u0_u0_u4_n67 ) );
  INV_X1 u0_u0_u4_U20 (.ZN( u0_u0_u4_n12 ) , .A( u0_u0_u4_n31 ) );
  NAND2_X1 u0_u0_u4_U21 (.A1( u0_u0_u4_n40 ) , .ZN( u0_u0_u4_n56 ) , .A2( u0_u0_u4_n69 ) );
  NAND2_X1 u0_u0_u4_U22 (.ZN( u0_u0_u4_n57 ) , .A2( u0_u0_u4_n67 ) , .A1( u0_u0_u4_n68 ) );
  NAND2_X1 u0_u0_u4_U23 (.A1( u0_u0_u4_n39 ) , .A2( u0_u0_u4_n69 ) , .ZN( u0_u0_u4_n70 ) );
  NAND2_X1 u0_u0_u4_U24 (.A2( u0_u0_u4_n39 ) , .A1( u0_u0_u4_n53 ) , .ZN( u0_u0_u4_n58 ) );
  AND3_X1 u0_u0_u4_U25 (.ZN( u0_u0_u4_n26 ) , .A3( u0_u0_u4_n33 ) , .A2( u0_u0_u4_n44 ) , .A1( u0_u0_u4_n68 ) );
  AND2_X1 u0_u0_u4_U26 (.ZN( u0_u0_u4_n28 ) , .A2( u0_u0_u4_n40 ) , .A1( u0_u0_u4_n42 ) );
  OR3_X1 u0_u0_u4_U27 (.ZN( u0_u0_u4_n51 ) , .A1( u0_u0_u4_n71 ) , .A2( u0_u0_u4_n72 ) , .A3( u0_u0_u4_n73 ) );
  AOI21_X1 u0_u0_u4_U28 (.B1( u0_u0_u4_n13 ) , .B2( u0_u0_u4_n14 ) , .ZN( u0_u0_u4_n71 ) , .A( u0_u0_u4_n74 ) );
  AOI21_X1 u0_u0_u4_U29 (.A( u0_u0_u4_n31 ) , .B1( u0_u0_u4_n41 ) , .B2( u0_u0_u4_n42 ) , .ZN( u0_u0_u4_n72 ) );
  NOR2_X1 u0_u0_u4_U3 (.A2( u0_u0_u4_n5 ) , .A1( u0_u0_u4_n6 ) , .ZN( u0_u0_u4_n66 ) );
  OAI22_X1 u0_u0_u4_U30 (.A1( u0_u0_u4_n16 ) , .B2( u0_u0_u4_n17 ) , .B1( u0_u0_u4_n27 ) , .A2( u0_u0_u4_n66 ) , .ZN( u0_u0_u4_n73 ) );
  INV_X1 u0_u0_u4_U31 (.A( u0_u0_u4_n29 ) , .ZN( u0_u0_u4_n5 ) );
  INV_X1 u0_u0_u4_U32 (.ZN( u0_u0_u4_n6 ) , .A( u0_u0_u4_n91 ) );
  INV_X1 u0_u0_u4_U33 (.A( u0_u0_u4_n43 ) , .ZN( u0_u0_u4_n8 ) );
  INV_X1 u0_u0_u4_U34 (.A( u0_u0_u4_n30 ) , .ZN( u0_u0_u4_n9 ) );
  NAND2_X1 u0_u0_u4_U35 (.A2( u0_u0_u4_n33 ) , .ZN( u0_u0_u4_n90 ) , .A1( u0_u0_u4_n91 ) );
  INV_X1 u0_u0_u4_U36 (.ZN( u0_u0_u4_n1 ) , .A( u0_u0_u4_n92 ) );
  OAI221_X1 u0_u0_u4_U37 (.C2( u0_u0_u4_n14 ) , .B2( u0_u0_u4_n16 ) , .B1( u0_u0_u4_n29 ) , .C1( u0_u0_u4_n53 ) , .ZN( u0_u0_u4_n92 ) , .A( u0_u0_u4_n93 ) );
  AOI222_X1 u0_u0_u4_U38 (.C2( u0_u0_u4_n12 ) , .B1( u0_u0_u4_n2 ) , .A1( u0_u0_u4_n49 ) , .B2( u0_u0_u4_n55 ) , .C1( u0_u0_u4_n6 ) , .A2( u0_u0_u4_n8 ) , .ZN( u0_u0_u4_n93 ) );
  INV_X1 u0_u0_u4_U39 (.ZN( u0_u0_u4_n2 ) , .A( u0_u0_u4_n74 ) );
  INV_X1 u0_u0_u4_U4 (.ZN( u0_u0_u4_n3 ) , .A( u0_u0_u4_n70 ) );
  INV_X1 u0_u0_u4_U40 (.ZN( u0_u0_u4_n4 ) , .A( u0_u0_u4_n44 ) );
  NOR2_X1 u0_u0_u4_U41 (.A2( u0_u0_u4_n18 ) , .A1( u0_u0_u4_n19 ) , .ZN( u0_u0_u4_n49 ) );
  NOR2_X1 u0_u0_u4_U42 (.ZN( u0_u0_u4_n34 ) , .A2( u0_u0_u4_n35 ) , .A1( u0_u0_u4_n37 ) );
  NOR2_X1 u0_u0_u4_U43 (.ZN( u0_u0_u4_n31 ) , .A1( u0_u0_u4_n49 ) , .A2( u0_u0_u4_n59 ) );
  AOI22_X1 u0_u0_u4_U44 (.A2( u0_u0_u4_n15 ) , .B1( u0_u0_u4_n59 ) , .ZN( u0_u0_u4_n63 ) , .A1( u0_u0_u4_n64 ) , .B2( u0_u0_u4_n65 ) );
  INV_X1 u0_u0_u4_U45 (.ZN( u0_u0_u4_n15 ) , .A( u0_u0_u4_n34 ) );
  NAND2_X1 u0_u0_u4_U46 (.A1( u0_u0_u4_n26 ) , .ZN( u0_u0_u4_n64 ) , .A2( u0_u0_u4_n67 ) );
  AOI22_X1 u0_u0_u4_U47 (.A1( u0_u0_u4_n37 ) , .ZN( u0_u0_u4_n47 ) , .A2( u0_u0_u4_n54 ) , .B2( u0_u0_u4_n55 ) , .B1( u0_u0_u4_n8 ) );
  NAND2_X1 u0_u0_u4_U48 (.A1( u0_u0_u4_n33 ) , .A2( u0_u0_u4_n41 ) , .ZN( u0_u0_u4_n54 ) );
  NAND2_X1 u0_u0_u4_U49 (.ZN( u0_u0_u4_n33 ) , .A1( u0_u0_u4_n84 ) , .A2( u0_u0_u4_n89 ) );
  NOR4_X1 u0_u0_u4_U5 (.ZN( u0_u0_u4_n77 ) , .A1( u0_u0_u4_n78 ) , .A2( u0_u0_u4_n79 ) , .A3( u0_u0_u4_n80 ) , .A4( u0_u0_u4_n81 ) );
  NAND2_X1 u0_u0_u4_U50 (.ZN( u0_u0_u4_n29 ) , .A1( u0_u0_u4_n86 ) , .A2( u0_u0_u4_n88 ) );
  AOI21_X1 u0_u0_u4_U51 (.B2( u0_u0_u4_n37 ) , .A( u0_u0_u4_n51 ) , .ZN( u0_u0_u4_n60 ) , .B1( u0_u0_u4_n7 ) );
  INV_X1 u0_u0_u4_U52 (.A( u0_u0_u4_n27 ) , .ZN( u0_u0_u4_n7 ) );
  NAND2_X1 u0_u0_u4_U53 (.ZN( u0_u0_u4_n41 ) , .A1( u0_u0_u4_n82 ) , .A2( u0_u0_u4_n83 ) );
  NAND2_X1 u0_u0_u4_U54 (.ZN( u0_u0_u4_n27 ) , .A1( u0_u0_u4_n85 ) , .A2( u0_u0_u4_n86 ) );
  NAND2_X1 u0_u0_u4_U55 (.ZN( u0_u0_u4_n53 ) , .A2( u0_u0_u4_n88 ) , .A1( u0_u0_u4_n89 ) );
  NAND2_X1 u0_u0_u4_U56 (.ZN( u0_u0_u4_n44 ) , .A2( u0_u0_u4_n83 ) , .A1( u0_u0_u4_n84 ) );
  NAND2_X1 u0_u0_u4_U57 (.ZN( u0_u0_u4_n42 ) , .A2( u0_u0_u4_n82 ) , .A1( u0_u0_u4_n89 ) );
  NAND2_X1 u0_u0_u4_U58 (.ZN( u0_u0_u4_n67 ) , .A2( u0_u0_u4_n82 ) , .A1( u0_u0_u4_n87 ) );
  NAND2_X1 u0_u0_u4_U59 (.ZN( u0_u0_u4_n39 ) , .A2( u0_u0_u4_n83 ) , .A1( u0_u0_u4_n85 ) );
  AOI21_X1 u0_u0_u4_U6 (.A( u0_u0_u4_n17 ) , .B1( u0_u0_u4_n29 ) , .B2( u0_u0_u4_n41 ) , .ZN( u0_u0_u4_n81 ) );
  NAND2_X1 u0_u0_u4_U60 (.ZN( u0_u0_u4_n30 ) , .A1( u0_u0_u4_n84 ) , .A2( u0_u0_u4_n87 ) );
  INV_X1 u0_u0_u4_U61 (.ZN( u0_u0_u4_n14 ) , .A( u0_u0_u4_n37 ) );
  INV_X1 u0_u0_u4_U62 (.ZN( u0_u0_u4_n16 ) , .A( u0_u0_u4_n35 ) );
  NAND2_X1 u0_u0_u4_U63 (.ZN( u0_u0_u4_n69 ) , .A1( u0_u0_u4_n87 ) , .A2( u0_u0_u4_n88 ) );
  NAND2_X1 u0_u0_u4_U64 (.ZN( u0_u0_u4_n43 ) , .A1( u0_u0_u4_n85 ) , .A2( u0_u0_u4_n87 ) );
  NAND2_X1 u0_u0_u4_U65 (.A1( u0_u0_u4_n82 ) , .A2( u0_u0_u4_n86 ) , .ZN( u0_u0_u4_n91 ) );
  INV_X1 u0_u0_u4_U66 (.ZN( u0_u0_u4_n13 ) , .A( u0_u0_u4_n59 ) );
  NAND2_X1 u0_u0_u4_U67 (.ZN( u0_u0_u4_n68 ) , .A2( u0_u0_u4_n85 ) , .A1( u0_u0_u4_n89 ) );
  NAND2_X1 u0_u0_u4_U68 (.ZN( u0_u0_u4_n40 ) , .A1( u0_u0_u4_n84 ) , .A2( u0_u0_u4_n86 ) );
  NAND2_X1 u0_u0_u4_U69 (.ZN( u0_u0_u4_n74 ) , .A2( u0_u0_u4_n83 ) , .A1( u0_u0_u4_n88 ) );
  AOI21_X1 u0_u0_u4_U7 (.A( u0_u0_u4_n31 ) , .B1( u0_u0_u4_n32 ) , .B2( u0_u0_u4_n53 ) , .ZN( u0_u0_u4_n79 ) );
  NOR2_X1 u0_u0_u4_U70 (.A2( u0_u0_X_28 ) , .A1( u0_u0_u4_n19 ) , .ZN( u0_u0_u4_n37 ) );
  NOR2_X1 u0_u0_u4_U71 (.A2( u0_u0_X_29 ) , .A1( u0_u0_u4_n18 ) , .ZN( u0_u0_u4_n35 ) );
  NOR2_X1 u0_u0_u4_U72 (.A2( u0_u0_X_30 ) , .A1( u0_u0_u4_n11 ) , .ZN( u0_u0_u4_n82 ) );
  NOR2_X1 u0_u0_u4_U73 (.A2( u0_u0_X_26 ) , .A1( u0_u0_u4_n10 ) , .ZN( u0_u0_u4_n87 ) );
  NOR2_X1 u0_u0_u4_U74 (.A2( u0_u0_X_28 ) , .A1( u0_u0_X_29 ) , .ZN( u0_u0_u4_n59 ) );
  NOR2_X1 u0_u0_u4_U75 (.A2( u0_u0_X_27 ) , .A1( u0_u0_X_30 ) , .ZN( u0_u0_u4_n85 ) );
  NOR2_X1 u0_u0_u4_U76 (.A2( u0_u0_X_25 ) , .A1( u0_u0_X_26 ) , .ZN( u0_u0_u4_n89 ) );
  AND2_X1 u0_u0_u4_U77 (.A2( u0_u0_X_25 ) , .A1( u0_u0_X_26 ) , .ZN( u0_u0_u4_n83 ) );
  AND2_X1 u0_u0_u4_U78 (.A1( u0_u0_X_30 ) , .A2( u0_u0_u4_n11 ) , .ZN( u0_u0_u4_n88 ) );
  AND2_X1 u0_u0_u4_U79 (.A1( u0_u0_X_26 ) , .A2( u0_u0_u4_n10 ) , .ZN( u0_u0_u4_n86 ) );
  AOI21_X1 u0_u0_u4_U8 (.B1( u0_u0_u4_n28 ) , .B2( u0_u0_u4_n3 ) , .A( u0_u0_u4_n34 ) , .ZN( u0_u0_u4_n78 ) );
  AND2_X1 u0_u0_u4_U80 (.A1( u0_u0_X_27 ) , .A2( u0_u0_X_30 ) , .ZN( u0_u0_u4_n84 ) );
  INV_X1 u0_u0_u4_U81 (.A( u0_u0_X_28 ) , .ZN( u0_u0_u4_n18 ) );
  INV_X1 u0_u0_u4_U82 (.A( u0_u0_X_29 ) , .ZN( u0_u0_u4_n19 ) );
  INV_X1 u0_u0_u4_U83 (.A( u0_u0_X_25 ) , .ZN( u0_u0_u4_n10 ) );
  INV_X1 u0_u0_u4_U84 (.A( u0_u0_X_27 ) , .ZN( u0_u0_u4_n11 ) );
  NAND4_X1 u0_u0_u4_U85 (.ZN( u0_out0_25 ) , .A1( u0_u0_u4_n45 ) , .A2( u0_u0_u4_n46 ) , .A3( u0_u0_u4_n47 ) , .A4( u0_u0_u4_n48 ) );
  OAI21_X1 u0_u0_u4_U86 (.ZN( u0_u0_u4_n45 ) , .B1( u0_u0_u4_n57 ) , .B2( u0_u0_u4_n58 ) , .A( u0_u0_u4_n59 ) );
  OAI21_X1 u0_u0_u4_U87 (.A( u0_u0_u4_n12 ) , .B1( u0_u0_u4_n4 ) , .ZN( u0_u0_u4_n46 ) , .B2( u0_u0_u4_n56 ) );
  NAND4_X1 u0_u0_u4_U88 (.ZN( u0_out0_14 ) , .A1( u0_u0_u4_n60 ) , .A2( u0_u0_u4_n61 ) , .A3( u0_u0_u4_n62 ) , .A4( u0_u0_u4_n63 ) );
  AOI22_X1 u0_u0_u4_U89 (.A2( u0_u0_u4_n12 ) , .B1( u0_u0_u4_n35 ) , .A1( u0_u0_u4_n58 ) , .ZN( u0_u0_u4_n61 ) , .B2( u0_u0_u4_n70 ) );
  AOI211_X1 u0_u0_u4_U9 (.ZN( u0_u0_u4_n48 ) , .C2( u0_u0_u4_n49 ) , .C1( u0_u0_u4_n5 ) , .A( u0_u0_u4_n50 ) , .B( u0_u0_u4_n51 ) );
  AOI22_X1 u0_u0_u4_U90 (.B1( u0_u0_u4_n49 ) , .A2( u0_u0_u4_n55 ) , .B2( u0_u0_u4_n56 ) , .ZN( u0_u0_u4_n62 ) , .A1( u0_u0_u4_n9 ) );
  NAND4_X1 u0_u0_u4_U91 (.ZN( u0_out0_8 ) , .A1( u0_u0_u4_n1 ) , .A2( u0_u0_u4_n75 ) , .A3( u0_u0_u4_n76 ) , .A4( u0_u0_u4_n77 ) );
  NAND2_X1 u0_u0_u4_U92 (.A1( u0_u0_u4_n37 ) , .A2( u0_u0_u4_n57 ) , .ZN( u0_u0_u4_n75 ) );
  AOI22_X1 u0_u0_u4_U93 (.A1( u0_u0_u4_n35 ) , .B2( u0_u0_u4_n55 ) , .ZN( u0_u0_u4_n76 ) , .B1( u0_u0_u4_n9 ) , .A2( u0_u0_u4_n90 ) );
  AOI22_X1 u0_u0_u4_U94 (.ZN( u0_u0_u4_n20 ) , .A1( u0_u0_u4_n35 ) , .A2( u0_u0_u4_n36 ) , .B1( u0_u0_u4_n37 ) , .B2( u0_u0_u4_n38 ) );
  NOR4_X1 u0_u0_u4_U95 (.ZN( u0_u0_u4_n21 ) , .A1( u0_u0_u4_n22 ) , .A2( u0_u0_u4_n23 ) , .A3( u0_u0_u4_n24 ) , .A4( u0_u0_u4_n25 ) );
  NAND3_X1 u0_u0_u4_U96 (.ZN( u0_out0_3 ) , .A2( u0_u0_u4_n1 ) , .A1( u0_u0_u4_n20 ) , .A3( u0_u0_u4_n21 ) );
  NAND3_X1 u0_u0_u4_U97 (.ZN( u0_u0_u4_n38 ) , .A1( u0_u0_u4_n39 ) , .A2( u0_u0_u4_n40 ) , .A3( u0_u0_u4_n41 ) );
  NAND3_X1 u0_u0_u4_U98 (.ZN( u0_u0_u4_n36 ) , .A1( u0_u0_u4_n42 ) , .A2( u0_u0_u4_n43 ) , .A3( u0_u0_u4_n44 ) );
  NAND3_X1 u0_u0_u4_U99 (.A1( u0_u0_u4_n33 ) , .A2( u0_u0_u4_n43 ) , .ZN( u0_u0_u4_n65 ) , .A3( u0_u0_u4_n66 ) );
  INV_X1 u0_u0_u5_U10 (.ZN( u0_u0_u5_n20 ) , .A( u0_u0_u5_n76 ) );
  AOI222_X1 u0_u0_u5_U100 (.A2( u0_u0_u5_n18 ) , .C2( u0_u0_u5_n19 ) , .B2( u0_u0_u5_n23 ) , .C1( u0_u0_u5_n49 ) , .A1( u0_u0_u5_n66 ) , .ZN( u0_u0_u5_n84 ) , .B1( u0_u0_u5_n98 ) );
  NAND4_X1 u0_u0_u5_U101 (.ZN( u0_out0_29 ) , .A1( u0_u0_u5_n1 ) , .A2( u0_u0_u5_n29 ) , .A3( u0_u0_u5_n67 ) , .A4( u0_u0_u5_n68 ) );
  AOI221_X1 u0_u0_u5_U102 (.C1( u0_u0_u5_n13 ) , .B1( u0_u0_u5_n21 ) , .B2( u0_u0_u5_n38 ) , .C2( u0_u0_u5_n65 ) , .ZN( u0_u0_u5_n68 ) , .A( u0_u0_u5_n69 ) );
  AOI222_X1 u0_u0_u5_U103 (.B2( u0_u0_u5_n18 ) , .C2( u0_u0_u5_n22 ) , .C1( u0_u0_u5_n3 ) , .B1( u0_u0_u5_n50 ) , .A2( u0_u0_u5_n51 ) , .ZN( u0_u0_u5_n67 ) , .A1( u0_u0_u5_n9 ) );
  NAND3_X1 u0_u0_u5_U104 (.A1( u0_u0_u5_n36 ) , .A3( u0_u0_u5_n39 ) , .A2( u0_u0_u5_n43 ) , .ZN( u0_u0_u5_n98 ) );
  NOR2_X1 u0_u0_u5_U11 (.A1( u0_u0_u5_n20 ) , .A2( u0_u0_u5_n24 ) , .ZN( u0_u0_u5_n37 ) );
  INV_X1 u0_u0_u5_U12 (.ZN( u0_u0_u5_n23 ) , .A( u0_u0_u5_n47 ) );
  AOI21_X1 u0_u0_u5_U13 (.ZN( u0_u0_u5_n35 ) , .B2( u0_u0_u5_n36 ) , .A( u0_u0_u5_n37 ) , .B1( u0_u0_u5_n5 ) );
  INV_X1 u0_u0_u5_U14 (.A( u0_u0_u5_n38 ) , .ZN( u0_u0_u5_n5 ) );
  AOI21_X1 u0_u0_u5_U15 (.ZN( u0_u0_u5_n34 ) , .B1( u0_u0_u5_n39 ) , .B2( u0_u0_u5_n40 ) , .A( u0_u0_u5_n41 ) );
  AOI21_X1 u0_u0_u5_U16 (.A( u0_u0_u5_n47 ) , .ZN( u0_u0_u5_n56 ) , .B1( u0_u0_u5_n57 ) , .B2( u0_u0_u5_n58 ) );
  OAI21_X1 u0_u0_u5_U17 (.ZN( u0_u0_u5_n55 ) , .B1( u0_u0_u5_n62 ) , .B2( u0_u0_u5_n63 ) , .A( u0_u0_u5_n64 ) );
  OAI21_X1 u0_u0_u5_U18 (.A( u0_u0_u5_n24 ) , .B2( u0_u0_u5_n50 ) , .ZN( u0_u0_u5_n64 ) , .B1( u0_u0_u5_n9 ) );
  NAND2_X1 u0_u0_u5_U19 (.ZN( u0_u0_u5_n60 ) , .A1( u0_u0_u5_n74 ) , .A2( u0_u0_u5_n78 ) );
  INV_X1 u0_u0_u5_U20 (.ZN( u0_u0_u5_n3 ) , .A( u0_u0_u5_n42 ) );
  NAND2_X1 u0_u0_u5_U21 (.A2( u0_u0_u5_n25 ) , .ZN( u0_u0_u5_n65 ) , .A1( u0_u0_u5_n76 ) );
  NAND2_X1 u0_u0_u5_U22 (.A1( u0_u0_u5_n43 ) , .ZN( u0_u0_u5_n61 ) , .A2( u0_u0_u5_n75 ) );
  NAND2_X1 u0_u0_u5_U23 (.ZN( u0_u0_u5_n38 ) , .A1( u0_u0_u5_n77 ) , .A2( u0_u0_u5_n78 ) );
  INV_X1 u0_u0_u5_U24 (.ZN( u0_u0_u5_n22 ) , .A( u0_u0_u5_n41 ) );
  INV_X1 u0_u0_u5_U25 (.A( u0_u0_u5_n39 ) , .ZN( u0_u0_u5_n9 ) );
  INV_X1 u0_u0_u5_U26 (.ZN( u0_u0_u5_n18 ) , .A( u0_u0_u5_n45 ) );
  INV_X1 u0_u0_u5_U27 (.ZN( u0_u0_u5_n15 ) , .A( u0_u0_u5_n57 ) );
  INV_X1 u0_u0_u5_U28 (.ZN( u0_u0_u5_n14 ) , .A( u0_u0_u5_n46 ) );
  INV_X1 u0_u0_u5_U29 (.ZN( u0_u0_u5_n12 ) , .A( u0_u0_u5_n74 ) );
  NOR2_X1 u0_u0_u5_U3 (.A1( u0_u0_u5_n14 ) , .ZN( u0_u0_u5_n63 ) , .A2( u0_u0_u5_n7 ) );
  INV_X1 u0_u0_u5_U30 (.ZN( u0_u0_u5_n13 ) , .A( u0_u0_u5_n36 ) );
  INV_X1 u0_u0_u5_U31 (.A( u0_u0_u5_n58 ) , .ZN( u0_u0_u5_n8 ) );
  INV_X1 u0_u0_u5_U32 (.A( u0_u0_u5_n40 ) , .ZN( u0_u0_u5_n7 ) );
  INV_X1 u0_u0_u5_U33 (.ZN( u0_u0_u5_n4 ) , .A( u0_u0_u5_n77 ) );
  NAND2_X1 u0_u0_u5_U34 (.A2( u0_u0_u5_n42 ) , .A1( u0_u0_u5_n57 ) , .ZN( u0_u0_u5_n86 ) );
  NOR2_X1 u0_u0_u5_U35 (.A2( u0_u0_u5_n17 ) , .A1( u0_u0_u5_n27 ) , .ZN( u0_u0_u5_n97 ) );
  INV_X1 u0_u0_u5_U36 (.ZN( u0_u0_u5_n1 ) , .A( u0_u0_u5_n80 ) );
  OAI221_X1 u0_u0_u5_U37 (.B1( u0_u0_u5_n25 ) , .C2( u0_u0_u5_n39 ) , .C1( u0_u0_u5_n44 ) , .B2( u0_u0_u5_n78 ) , .ZN( u0_u0_u5_n80 ) , .A( u0_u0_u5_n81 ) );
  AOI222_X1 u0_u0_u5_U38 (.B1( u0_u0_u5_n10 ) , .C2( u0_u0_u5_n20 ) , .A2( u0_u0_u5_n23 ) , .A1( u0_u0_u5_n4 ) , .C1( u0_u0_u5_n49 ) , .B2( u0_u0_u5_n52 ) , .ZN( u0_u0_u5_n81 ) );
  INV_X1 u0_u0_u5_U39 (.ZN( u0_u0_u5_n10 ) , .A( u0_u0_u5_n82 ) );
  INV_X1 u0_u0_u5_U4 (.A( u0_u0_u5_n59 ) , .ZN( u0_u0_u5_n6 ) );
  AOI22_X1 u0_u0_u5_U40 (.A1( u0_u0_u5_n12 ) , .B1( u0_u0_u5_n23 ) , .ZN( u0_u0_u5_n28 ) , .A2( u0_u0_u5_n51 ) , .B2( u0_u0_u5_n66 ) );
  NOR2_X1 u0_u0_u5_U41 (.A2( u0_u0_u5_n24 ) , .ZN( u0_u0_u5_n47 ) , .A1( u0_u0_u5_n51 ) );
  AOI21_X1 u0_u0_u5_U42 (.B1( u0_u0_u5_n11 ) , .ZN( u0_u0_u5_n29 ) , .B2( u0_u0_u5_n52 ) , .A( u0_u0_u5_n79 ) );
  INV_X1 u0_u0_u5_U43 (.ZN( u0_u0_u5_n11 ) , .A( u0_u0_u5_n75 ) );
  NOR2_X1 u0_u0_u5_U44 (.A2( u0_u0_u5_n21 ) , .ZN( u0_u0_u5_n45 ) , .A1( u0_u0_u5_n51 ) );
  NOR2_X1 u0_u0_u5_U45 (.A2( u0_u0_u5_n44 ) , .ZN( u0_u0_u5_n79 ) , .A1( u0_u0_u5_n82 ) );
  NOR2_X1 u0_u0_u5_U46 (.A1( u0_u0_u5_n23 ) , .ZN( u0_u0_u5_n41 ) , .A2( u0_u0_u5_n52 ) );
  NOR2_X1 u0_u0_u5_U47 (.A1( u0_u0_u5_n21 ) , .A2( u0_u0_u5_n52 ) , .ZN( u0_u0_u5_n76 ) );
  AOI22_X1 u0_u0_u5_U48 (.B2( u0_u0_u5_n22 ) , .B1( u0_u0_u5_n4 ) , .A1( u0_u0_u5_n52 ) , .A2( u0_u0_u5_n60 ) , .ZN( u0_u0_u5_n83 ) );
  OAI211_X1 u0_u0_u5_U49 (.ZN( u0_u0_u5_n69 ) , .C1( u0_u0_u5_n70 ) , .C2( u0_u0_u5_n71 ) , .A( u0_u0_u5_n72 ) , .B( u0_u0_u5_n73 ) );
  OAI21_X1 u0_u0_u5_U5 (.A( u0_u0_u5_n20 ) , .ZN( u0_u0_u5_n59 ) , .B1( u0_u0_u5_n60 ) , .B2( u0_u0_u5_n61 ) );
  NOR3_X1 u0_u0_u5_U50 (.A2( u0_u0_u5_n15 ) , .A3( u0_u0_u5_n49 ) , .A1( u0_u0_u5_n61 ) , .ZN( u0_u0_u5_n70 ) );
  OAI21_X1 u0_u0_u5_U51 (.B2( u0_u0_u5_n14 ) , .A( u0_u0_u5_n20 ) , .ZN( u0_u0_u5_n73 ) , .B1( u0_u0_u5_n8 ) );
  OAI21_X1 u0_u0_u5_U52 (.B2( u0_u0_u5_n12 ) , .A( u0_u0_u5_n23 ) , .B1( u0_u0_u5_n7 ) , .ZN( u0_u0_u5_n72 ) );
  AOI21_X1 u0_u0_u5_U53 (.ZN( u0_u0_u5_n33 ) , .B1( u0_u0_u5_n42 ) , .B2( u0_u0_u5_n43 ) , .A( u0_u0_u5_n44 ) );
  AOI21_X1 u0_u0_u5_U54 (.A( u0_u0_u5_n44 ) , .B2( u0_u0_u5_n58 ) , .B1( u0_u0_u5_n75 ) , .ZN( u0_u0_u5_n87 ) );
  INV_X1 u0_u0_u5_U55 (.ZN( u0_u0_u5_n21 ) , .A( u0_u0_u5_n44 ) );
  INV_X1 u0_u0_u5_U56 (.ZN( u0_u0_u5_n24 ) , .A( u0_u0_u5_n71 ) );
  AND2_X1 u0_u0_u5_U57 (.ZN( u0_u0_u5_n50 ) , .A1( u0_u0_u5_n90 ) , .A2( u0_u0_u5_n93 ) );
  AND2_X1 u0_u0_u5_U58 (.ZN( u0_u0_u5_n49 ) , .A1( u0_u0_u5_n89 ) , .A2( u0_u0_u5_n93 ) );
  NAND2_X1 u0_u0_u5_U59 (.ZN( u0_u0_u5_n39 ) , .A2( u0_u0_u5_n91 ) , .A1( u0_u0_u5_n92 ) );
  INV_X1 u0_u0_u5_U6 (.ZN( u0_u0_u5_n19 ) , .A( u0_u0_u5_n62 ) );
  NAND2_X1 u0_u0_u5_U60 (.ZN( u0_u0_u5_n58 ) , .A1( u0_u0_u5_n88 ) , .A2( u0_u0_u5_n89 ) );
  NAND2_X1 u0_u0_u5_U61 (.ZN( u0_u0_u5_n78 ) , .A2( u0_u0_u5_n89 ) , .A1( u0_u0_u5_n91 ) );
  NAND2_X1 u0_u0_u5_U62 (.ZN( u0_u0_u5_n57 ) , .A1( u0_u0_u5_n92 ) , .A2( u0_u0_u5_n94 ) );
  NAND2_X1 u0_u0_u5_U63 (.ZN( u0_u0_u5_n42 ) , .A1( u0_u0_u5_n92 ) , .A2( u0_u0_u5_n93 ) );
  NAND2_X1 u0_u0_u5_U64 (.ZN( u0_u0_u5_n75 ) , .A1( u0_u0_u5_n90 ) , .A2( u0_u0_u5_n91 ) );
  NAND2_X1 u0_u0_u5_U65 (.ZN( u0_u0_u5_n82 ) , .A1( u0_u0_u5_n91 ) , .A2( u0_u0_u5_n97 ) );
  NAND2_X1 u0_u0_u5_U66 (.ZN( u0_u0_u5_n36 ) , .A1( u0_u0_u5_n94 ) , .A2( u0_u0_u5_n97 ) );
  NAND2_X1 u0_u0_u5_U67 (.ZN( u0_u0_u5_n43 ) , .A2( u0_u0_u5_n88 ) , .A1( u0_u0_u5_n92 ) );
  INV_X1 u0_u0_u5_U68 (.ZN( u0_u0_u5_n25 ) , .A( u0_u0_u5_n51 ) );
  NAND2_X1 u0_u0_u5_U69 (.ZN( u0_u0_u5_n74 ) , .A2( u0_u0_u5_n89 ) , .A1( u0_u0_u5_n94 ) );
  OAI22_X1 u0_u0_u5_U7 (.ZN( u0_u0_u5_n32 ) , .A1( u0_u0_u5_n45 ) , .A2( u0_u0_u5_n46 ) , .B1( u0_u0_u5_n47 ) , .B2( u0_u0_u5_n48 ) );
  NAND2_X1 u0_u0_u5_U70 (.ZN( u0_u0_u5_n46 ) , .A1( u0_u0_u5_n90 ) , .A2( u0_u0_u5_n94 ) );
  NAND2_X1 u0_u0_u5_U71 (.ZN( u0_u0_u5_n77 ) , .A1( u0_u0_u5_n88 ) , .A2( u0_u0_u5_n90 ) );
  NAND2_X1 u0_u0_u5_U72 (.ZN( u0_u0_u5_n40 ) , .A1( u0_u0_u5_n88 ) , .A2( u0_u0_u5_n97 ) );
  AND2_X1 u0_u0_u5_U73 (.ZN( u0_u0_u5_n66 ) , .A1( u0_u0_u5_n93 ) , .A2( u0_u0_u5_n97 ) );
  INV_X1 u0_u0_u5_U74 (.ZN( u0_u0_u5_n2 ) , .A( u0_u0_u5_n95 ) );
  OAI221_X1 u0_u0_u5_U75 (.B2( u0_u0_u5_n37 ) , .B1( u0_u0_u5_n63 ) , .C1( u0_u0_u5_n71 ) , .C2( u0_u0_u5_n82 ) , .ZN( u0_u0_u5_n95 ) , .A( u0_u0_u5_n96 ) );
  OAI21_X1 u0_u0_u5_U76 (.B2( u0_u0_u5_n50 ) , .A( u0_u0_u5_n51 ) , .B1( u0_u0_u5_n60 ) , .ZN( u0_u0_u5_n96 ) );
  NOR2_X1 u0_u0_u5_U77 (.A2( u0_u0_X_34 ) , .A1( u0_u0_X_35 ) , .ZN( u0_u0_u5_n52 ) );
  NOR2_X1 u0_u0_u5_U78 (.A2( u0_u0_X_34 ) , .A1( u0_u0_u5_n26 ) , .ZN( u0_u0_u5_n51 ) );
  NOR2_X1 u0_u0_u5_U79 (.A2( u0_u0_X_31 ) , .A1( u0_u0_X_32 ) , .ZN( u0_u0_u5_n94 ) );
  NOR3_X1 u0_u0_u5_U8 (.A3( u0_u0_u5_n3 ) , .ZN( u0_u0_u5_n48 ) , .A1( u0_u0_u5_n49 ) , .A2( u0_u0_u5_n50 ) );
  NOR2_X1 u0_u0_u5_U80 (.A2( u0_u0_X_36 ) , .A1( u0_u0_u5_n17 ) , .ZN( u0_u0_u5_n92 ) );
  NOR2_X1 u0_u0_u5_U81 (.A2( u0_u0_X_33 ) , .A1( u0_u0_u5_n27 ) , .ZN( u0_u0_u5_n89 ) );
  NOR2_X1 u0_u0_u5_U82 (.A2( u0_u0_X_33 ) , .A1( u0_u0_X_36 ) , .ZN( u0_u0_u5_n90 ) );
  NOR2_X1 u0_u0_u5_U83 (.A2( u0_u0_X_31 ) , .A1( u0_u0_u5_n16 ) , .ZN( u0_u0_u5_n93 ) );
  NAND2_X1 u0_u0_u5_U84 (.A2( u0_u0_X_34 ) , .A1( u0_u0_X_35 ) , .ZN( u0_u0_u5_n44 ) );
  NAND2_X1 u0_u0_u5_U85 (.A1( u0_u0_X_34 ) , .A2( u0_u0_u5_n26 ) , .ZN( u0_u0_u5_n71 ) );
  AND2_X1 u0_u0_u5_U86 (.A1( u0_u0_X_31 ) , .A2( u0_u0_X_32 ) , .ZN( u0_u0_u5_n91 ) );
  AND2_X1 u0_u0_u5_U87 (.A1( u0_u0_X_31 ) , .A2( u0_u0_u5_n16 ) , .ZN( u0_u0_u5_n88 ) );
  INV_X1 u0_u0_u5_U88 (.A( u0_u0_X_33 ) , .ZN( u0_u0_u5_n17 ) );
  INV_X1 u0_u0_u5_U89 (.A( u0_u0_X_35 ) , .ZN( u0_u0_u5_n26 ) );
  NOR2_X1 u0_u0_u5_U9 (.A2( u0_u0_u5_n21 ) , .A1( u0_u0_u5_n24 ) , .ZN( u0_u0_u5_n62 ) );
  INV_X1 u0_u0_u5_U90 (.A( u0_u0_X_36 ) , .ZN( u0_u0_u5_n27 ) );
  INV_X1 u0_u0_u5_U91 (.A( u0_u0_X_32 ) , .ZN( u0_u0_u5_n16 ) );
  NAND4_X1 u0_u0_u5_U92 (.ZN( u0_out0_19 ) , .A1( u0_u0_u5_n28 ) , .A2( u0_u0_u5_n29 ) , .A3( u0_u0_u5_n30 ) , .A4( u0_u0_u5_n31 ) );
  AOI22_X1 u0_u0_u5_U93 (.B1( u0_u0_u5_n15 ) , .ZN( u0_u0_u5_n30 ) , .A2( u0_u0_u5_n51 ) , .B2( u0_u0_u5_n52 ) , .A1( u0_u0_u5_n8 ) );
  NOR4_X1 u0_u0_u5_U94 (.ZN( u0_u0_u5_n31 ) , .A1( u0_u0_u5_n32 ) , .A2( u0_u0_u5_n33 ) , .A3( u0_u0_u5_n34 ) , .A4( u0_u0_u5_n35 ) );
  NAND4_X1 u0_u0_u5_U95 (.ZN( u0_out0_11 ) , .A1( u0_u0_u5_n1 ) , .A2( u0_u0_u5_n28 ) , .A3( u0_u0_u5_n53 ) , .A4( u0_u0_u5_n54 ) );
  AOI22_X1 u0_u0_u5_U96 (.B1( u0_u0_u5_n13 ) , .A1( u0_u0_u5_n3 ) , .B2( u0_u0_u5_n52 ) , .ZN( u0_u0_u5_n53 ) , .A2( u0_u0_u5_n65 ) );
  NOR3_X1 u0_u0_u5_U97 (.ZN( u0_u0_u5_n54 ) , .A1( u0_u0_u5_n55 ) , .A3( u0_u0_u5_n56 ) , .A2( u0_u0_u5_n6 ) );
  NAND4_X1 u0_u0_u5_U98 (.ZN( u0_out0_4 ) , .A3( u0_u0_u5_n2 ) , .A1( u0_u0_u5_n83 ) , .A2( u0_u0_u5_n84 ) , .A4( u0_u0_u5_n85 ) );
  AOI211_X1 u0_u0_u5_U99 (.C2( u0_u0_u5_n20 ) , .B( u0_u0_u5_n79 ) , .ZN( u0_u0_u5_n85 ) , .C1( u0_u0_u5_n86 ) , .A( u0_u0_u5_n87 ) );
  AOI22_X1 u0_u0_u6_U10 (.B2( u0_u0_u6_n14 ) , .A2( u0_u0_u6_n24 ) , .B1( u0_u0_u6_n5 ) , .A1( u0_u0_u6_n8 ) , .ZN( u0_u0_u6_n86 ) );
  AOI21_X1 u0_u0_u6_U11 (.A( u0_u0_u6_n17 ) , .B2( u0_u0_u6_n43 ) , .B1( u0_u0_u6_n68 ) , .ZN( u0_u0_u6_n87 ) );
  AOI21_X1 u0_u0_u6_U12 (.A( u0_u0_u6_n17 ) , .ZN( u0_u0_u6_n26 ) , .B1( u0_u0_u6_n27 ) , .B2( u0_u0_u6_n28 ) );
  AOI21_X1 u0_u0_u6_U13 (.B1( u0_u0_u6_n11 ) , .B2( u0_u0_u6_n16 ) , .A( u0_u0_u6_n33 ) , .ZN( u0_u0_u6_n69 ) );
  INV_X1 u0_u0_u6_U14 (.ZN( u0_u0_u6_n14 ) , .A( u0_u0_u6_n20 ) );
  INV_X1 u0_u0_u6_U15 (.ZN( u0_u0_u6_n11 ) , .A( u0_u0_u6_n47 ) );
  NAND2_X1 u0_u0_u6_U16 (.A2( u0_u0_u6_n46 ) , .A1( u0_u0_u6_n53 ) , .ZN( u0_u0_u6_n65 ) );
  NAND2_X1 u0_u0_u6_U17 (.A1( u0_u0_u6_n27 ) , .A2( u0_u0_u6_n29 ) , .ZN( u0_u0_u6_n51 ) );
  INV_X1 u0_u0_u6_U18 (.ZN( u0_u0_u6_n4 ) , .A( u0_u0_u6_n43 ) );
  AND2_X1 u0_u0_u6_U19 (.A2( u0_u0_u6_n28 ) , .ZN( u0_u0_u6_n45 ) , .A1( u0_u0_u6_n75 ) );
  INV_X1 u0_u0_u6_U20 (.ZN( u0_u0_u6_n2 ) , .A( u0_u0_u6_n48 ) );
  INV_X1 u0_u0_u6_U21 (.A( u0_u0_u6_n54 ) , .ZN( u0_u0_u6_n8 ) );
  INV_X1 u0_u0_u6_U22 (.ZN( u0_u0_u6_n6 ) , .A( u0_u0_u6_n75 ) );
  INV_X1 u0_u0_u6_U23 (.ZN( u0_u0_u6_n5 ) , .A( u0_u0_u6_n52 ) );
  INV_X1 u0_u0_u6_U24 (.A( u0_u0_u6_n62 ) , .ZN( u0_u0_u6_n7 ) );
  AND2_X1 u0_u0_u6_U25 (.ZN( u0_u0_u6_n42 ) , .A2( u0_u0_u6_n56 ) , .A1( u0_u0_u6_n68 ) );
  AND2_X1 u0_u0_u6_U26 (.ZN( u0_u0_u6_n44 ) , .A1( u0_u0_u6_n53 ) , .A2( u0_u0_u6_n54 ) );
  AND3_X1 u0_u0_u6_U27 (.A3( u0_u0_u6_n30 ) , .A1( u0_u0_u6_n43 ) , .A2( u0_u0_u6_n48 ) , .ZN( u0_u0_u6_n55 ) );
  INV_X1 u0_u0_u6_U28 (.ZN( u0_u0_u6_n12 ) , .A( u0_u0_u6_n29 ) );
  AOI222_X1 u0_u0_u6_U29 (.C2( u0_u0_u6_n16 ) , .B2( u0_u0_u6_n24 ) , .A2( u0_u0_u6_n49 ) , .A1( u0_u0_u6_n57 ) , .B1( u0_u0_u6_n6 ) , .ZN( u0_u0_u6_n61 ) , .C1( u0_u0_u6_n7 ) );
  INV_X1 u0_u0_u6_U3 (.A( u0_u0_u6_n65 ) , .ZN( u0_u0_u6_n9 ) );
  NOR2_X1 u0_u0_u6_U30 (.A2( u0_u0_u6_n10 ) , .A1( u0_u0_u6_n13 ) , .ZN( u0_u0_u6_n77 ) );
  AOI211_X1 u0_u0_u6_U31 (.C2( u0_u0_u6_n24 ) , .ZN( u0_u0_u6_n38 ) , .C1( u0_u0_u6_n39 ) , .A( u0_u0_u6_n40 ) , .B( u0_u0_u6_n41 ) );
  AOI21_X1 u0_u0_u6_U32 (.A( u0_u0_u6_n17 ) , .ZN( u0_u0_u6_n41 ) , .B1( u0_u0_u6_n42 ) , .B2( u0_u0_u6_n43 ) );
  NAND4_X1 u0_u0_u6_U33 (.ZN( u0_u0_u6_n39 ) , .A1( u0_u0_u6_n45 ) , .A2( u0_u0_u6_n46 ) , .A3( u0_u0_u6_n47 ) , .A4( u0_u0_u6_n48 ) );
  AOI21_X1 u0_u0_u6_U34 (.B2( u0_u0_u6_n29 ) , .A( u0_u0_u6_n31 ) , .ZN( u0_u0_u6_n40 ) , .B1( u0_u0_u6_n44 ) );
  NAND2_X1 u0_u0_u6_U35 (.A2( u0_u0_u6_n17 ) , .ZN( u0_u0_u6_n24 ) , .A1( u0_u0_u6_n31 ) );
  NAND2_X1 u0_u0_u6_U36 (.ZN( u0_u0_u6_n43 ) , .A2( u0_u0_u6_n78 ) , .A1( u0_u0_u6_n84 ) );
  AOI22_X1 u0_u0_u6_U37 (.A2( u0_u0_u6_n14 ) , .ZN( u0_u0_u6_n60 ) , .A1( u0_u0_u6_n63 ) , .B1( u0_u0_u6_n64 ) , .B2( u0_u0_u6_n65 ) );
  NAND4_X1 u0_u0_u6_U38 (.A2( u0_u0_u6_n28 ) , .A4( u0_u0_u6_n43 ) , .ZN( u0_u0_u6_n63 ) , .A3( u0_u0_u6_n66 ) , .A1( u0_u0_u6_n9 ) );
  NOR2_X1 u0_u0_u6_U39 (.A2( u0_u0_u6_n2 ) , .A1( u0_u0_u6_n5 ) , .ZN( u0_u0_u6_n66 ) );
  INV_X1 u0_u0_u6_U4 (.ZN( u0_u0_u6_n1 ) , .A( u0_u0_u6_n33 ) );
  NOR2_X1 u0_u0_u6_U40 (.A1( u0_u0_u6_n15 ) , .ZN( u0_u0_u6_n20 ) , .A2( u0_u0_u6_n49 ) );
  NAND2_X1 u0_u0_u6_U41 (.ZN( u0_u0_u6_n29 ) , .A1( u0_u0_u6_n76 ) , .A2( u0_u0_u6_n81 ) );
  AOI21_X1 u0_u0_u6_U42 (.ZN( u0_u0_u6_n25 ) , .B1( u0_u0_u6_n29 ) , .B2( u0_u0_u6_n30 ) , .A( u0_u0_u6_n31 ) );
  INV_X1 u0_u0_u6_U43 (.ZN( u0_u0_u6_n17 ) , .A( u0_u0_u6_n64 ) );
  NAND2_X1 u0_u0_u6_U44 (.ZN( u0_u0_u6_n48 ) , .A2( u0_u0_u6_n83 ) , .A1( u0_u0_u6_n84 ) );
  NAND2_X1 u0_u0_u6_U45 (.ZN( u0_u0_u6_n46 ) , .A1( u0_u0_u6_n79 ) , .A2( u0_u0_u6_n80 ) );
  INV_X1 u0_u0_u6_U46 (.ZN( u0_u0_u6_n16 ) , .A( u0_u0_u6_n31 ) );
  NAND2_X1 u0_u0_u6_U47 (.ZN( u0_u0_u6_n30 ) , .A1( u0_u0_u6_n77 ) , .A2( u0_u0_u6_n78 ) );
  NAND2_X1 u0_u0_u6_U48 (.ZN( u0_u0_u6_n27 ) , .A1( u0_u0_u6_n81 ) , .A2( u0_u0_u6_n83 ) );
  NAND2_X1 u0_u0_u6_U49 (.A1( u0_u0_u6_n31 ) , .A2( u0_u0_u6_n36 ) , .ZN( u0_u0_u6_n67 ) );
  NAND2_X1 u0_u0_u6_U5 (.ZN( u0_u0_u6_n23 ) , .A2( u0_u0_u6_n32 ) , .A1( u0_u0_u6_n9 ) );
  NAND2_X1 u0_u0_u6_U50 (.ZN( u0_u0_u6_n54 ) , .A1( u0_u0_u6_n78 ) , .A2( u0_u0_u6_n80 ) );
  NAND2_X1 u0_u0_u6_U51 (.ZN( u0_u0_u6_n68 ) , .A1( u0_u0_u6_n80 ) , .A2( u0_u0_u6_n83 ) );
  AND2_X1 u0_u0_u6_U52 (.ZN( u0_u0_u6_n57 ) , .A1( u0_u0_u6_n76 ) , .A2( u0_u0_u6_n84 ) );
  NAND2_X1 u0_u0_u6_U53 (.ZN( u0_u0_u6_n28 ) , .A1( u0_u0_u6_n76 ) , .A2( u0_u0_u6_n77 ) );
  NAND2_X1 u0_u0_u6_U54 (.ZN( u0_u0_u6_n47 ) , .A2( u0_u0_u6_n79 ) , .A1( u0_u0_u6_n81 ) );
  NAND2_X1 u0_u0_u6_U55 (.ZN( u0_u0_u6_n56 ) , .A1( u0_u0_u6_n76 ) , .A2( u0_u0_u6_n80 ) );
  NAND2_X1 u0_u0_u6_U56 (.ZN( u0_u0_u6_n52 ) , .A1( u0_u0_u6_n79 ) , .A2( u0_u0_u6_n84 ) );
  NAND2_X1 u0_u0_u6_U57 (.ZN( u0_u0_u6_n75 ) , .A1( u0_u0_u6_n77 ) , .A2( u0_u0_u6_n83 ) );
  NAND2_X1 u0_u0_u6_U58 (.ZN( u0_u0_u6_n53 ) , .A2( u0_u0_u6_n78 ) , .A1( u0_u0_u6_n81 ) );
  INV_X1 u0_u0_u6_U59 (.ZN( u0_u0_u6_n15 ) , .A( u0_u0_u6_n36 ) );
  AOI22_X1 u0_u0_u6_U6 (.A2( u0_u0_u6_n14 ) , .B1( u0_u0_u6_n15 ) , .ZN( u0_u0_u6_n72 ) , .A1( u0_u0_u6_n73 ) , .B2( u0_u0_u6_n74 ) );
  NAND2_X1 u0_u0_u6_U60 (.ZN( u0_u0_u6_n62 ) , .A2( u0_u0_u6_n77 ) , .A1( u0_u0_u6_n79 ) );
  NOR2_X1 u0_u0_u6_U61 (.A2( u0_u0_X_40 ) , .A1( u0_u0_X_41 ) , .ZN( u0_u0_u6_n49 ) );
  NOR2_X1 u0_u0_u6_U62 (.A2( u0_u0_X_39 ) , .A1( u0_u0_X_42 ) , .ZN( u0_u0_u6_n83 ) );
  NOR2_X1 u0_u0_u6_U63 (.A2( u0_u0_X_39 ) , .A1( u0_u0_u6_n19 ) , .ZN( u0_u0_u6_n78 ) );
  NOR2_X1 u0_u0_u6_U64 (.A2( u0_u0_X_38 ) , .A1( u0_u0_u6_n10 ) , .ZN( u0_u0_u6_n80 ) );
  NOR2_X1 u0_u0_u6_U65 (.A2( u0_u0_X_41 ) , .A1( u0_u0_u6_n18 ) , .ZN( u0_u0_u6_n64 ) );
  NOR2_X1 u0_u0_u6_U66 (.A2( u0_u0_X_37 ) , .A1( u0_u0_u6_n13 ) , .ZN( u0_u0_u6_n81 ) );
  NOR2_X1 u0_u0_u6_U67 (.A2( u0_u0_X_37 ) , .A1( u0_u0_X_38 ) , .ZN( u0_u0_u6_n84 ) );
  NAND2_X1 u0_u0_u6_U68 (.A1( u0_u0_X_41 ) , .A2( u0_u0_u6_n18 ) , .ZN( u0_u0_u6_n31 ) );
  NAND2_X1 u0_u0_u6_U69 (.A2( u0_u0_X_40 ) , .A1( u0_u0_X_41 ) , .ZN( u0_u0_u6_n36 ) );
  NOR2_X1 u0_u0_u6_U7 (.ZN( u0_u0_u6_n32 ) , .A1( u0_u0_u6_n57 ) , .A2( u0_u0_u6_n7 ) );
  AND2_X1 u0_u0_u6_U70 (.A1( u0_u0_X_39 ) , .A2( u0_u0_u6_n19 ) , .ZN( u0_u0_u6_n79 ) );
  AND2_X1 u0_u0_u6_U71 (.A1( u0_u0_X_39 ) , .A2( u0_u0_X_42 ) , .ZN( u0_u0_u6_n76 ) );
  INV_X1 u0_u0_u6_U72 (.A( u0_u0_X_40 ) , .ZN( u0_u0_u6_n18 ) );
  INV_X1 u0_u0_u6_U73 (.A( u0_u0_X_37 ) , .ZN( u0_u0_u6_n10 ) );
  INV_X1 u0_u0_u6_U74 (.A( u0_u0_X_38 ) , .ZN( u0_u0_u6_n13 ) );
  INV_X1 u0_u0_u6_U75 (.A( u0_u0_X_42 ) , .ZN( u0_u0_u6_n19 ) );
  NAND4_X1 u0_u0_u6_U76 (.ZN( u0_out0_12 ) , .A1( u0_u0_u6_n58 ) , .A2( u0_u0_u6_n59 ) , .A3( u0_u0_u6_n60 ) , .A4( u0_u0_u6_n61 ) );
  OAI22_X1 u0_u0_u6_U77 (.A2( u0_u0_u6_n11 ) , .B1( u0_u0_u6_n49 ) , .ZN( u0_u0_u6_n59 ) , .B2( u0_u0_u6_n64 ) , .A1( u0_u0_u6_n8 ) );
  OAI21_X1 u0_u0_u6_U78 (.B1( u0_u0_u6_n12 ) , .B2( u0_u0_u6_n34 ) , .ZN( u0_u0_u6_n58 ) , .A( u0_u0_u6_n67 ) );
  NAND4_X1 u0_u0_u6_U79 (.ZN( u0_out0_32 ) , .A1( u0_u0_u6_n69 ) , .A2( u0_u0_u6_n70 ) , .A3( u0_u0_u6_n71 ) , .A4( u0_u0_u6_n72 ) );
  OAI21_X1 u0_u0_u6_U8 (.A( u0_u0_u6_n16 ) , .B2( u0_u0_u6_n2 ) , .B1( u0_u0_u6_n6 ) , .ZN( u0_u0_u6_n85 ) );
  AOI22_X1 u0_u0_u6_U80 (.B1( u0_u0_u6_n4 ) , .B2( u0_u0_u6_n49 ) , .A1( u0_u0_u6_n57 ) , .A2( u0_u0_u6_n67 ) , .ZN( u0_u0_u6_n70 ) );
  AOI22_X1 u0_u0_u6_U81 (.B2( u0_u0_u6_n24 ) , .B1( u0_u0_u6_n51 ) , .A1( u0_u0_u6_n64 ) , .ZN( u0_u0_u6_n71 ) , .A2( u0_u0_u6_n82 ) );
  OAI211_X1 u0_u0_u6_U82 (.ZN( u0_out0_7 ) , .A( u0_u0_u6_n1 ) , .C1( u0_u0_u6_n20 ) , .C2( u0_u0_u6_n21 ) , .B( u0_u0_u6_n22 ) );
  NOR3_X1 u0_u0_u6_U83 (.A3( u0_u0_u6_n11 ) , .ZN( u0_u0_u6_n21 ) , .A1( u0_u0_u6_n34 ) , .A2( u0_u0_u6_n4 ) );
  AOI211_X1 u0_u0_u6_U84 (.ZN( u0_u0_u6_n22 ) , .C1( u0_u0_u6_n23 ) , .C2( u0_u0_u6_n24 ) , .A( u0_u0_u6_n25 ) , .B( u0_u0_u6_n26 ) );
  OAI211_X1 u0_u0_u6_U85 (.ZN( u0_out0_22 ) , .C1( u0_u0_u6_n35 ) , .C2( u0_u0_u6_n36 ) , .A( u0_u0_u6_n37 ) , .B( u0_u0_u6_n38 ) );
  AOI22_X1 u0_u0_u6_U86 (.B2( u0_u0_u6_n14 ) , .ZN( u0_u0_u6_n37 ) , .A1( u0_u0_u6_n49 ) , .A2( u0_u0_u6_n50 ) , .B1( u0_u0_u6_n51 ) );
  AND4_X1 u0_u0_u6_U87 (.A2( u0_u0_u6_n32 ) , .ZN( u0_u0_u6_n35 ) , .A4( u0_u0_u6_n46 ) , .A1( u0_u0_u6_n55 ) , .A3( u0_u0_u6_n56 ) );
  NAND3_X1 u0_u0_u6_U88 (.A3( u0_u0_u6_n44 ) , .A1( u0_u0_u6_n45 ) , .ZN( u0_u0_u6_n50 ) , .A2( u0_u0_u6_n52 ) );
  NAND3_X1 u0_u0_u6_U89 (.A2( u0_u0_u6_n27 ) , .A1( u0_u0_u6_n30 ) , .ZN( u0_u0_u6_n34 ) , .A3( u0_u0_u6_n42 ) );
  INV_X1 u0_u0_u6_U9 (.ZN( u0_u0_u6_n3 ) , .A( u0_u0_u6_n87 ) );
  NAND3_X1 u0_u0_u6_U90 (.A1( u0_u0_u6_n48 ) , .A2( u0_u0_u6_n54 ) , .A3( u0_u0_u6_n68 ) , .ZN( u0_u0_u6_n74 ) );
  NAND3_X1 u0_u0_u6_U91 (.A2( u0_u0_u6_n30 ) , .A3( u0_u0_u6_n45 ) , .ZN( u0_u0_u6_n73 ) , .A1( u0_u0_u6_n9 ) );
  NAND3_X1 u0_u0_u6_U92 (.A2( u0_u0_u6_n52 ) , .A1( u0_u0_u6_n56 ) , .A3( u0_u0_u6_n62 ) , .ZN( u0_u0_u6_n82 ) );
  NAND3_X1 u0_u0_u6_U93 (.A2( u0_u0_u6_n3 ) , .ZN( u0_u0_u6_n33 ) , .A1( u0_u0_u6_n85 ) , .A3( u0_u0_u6_n86 ) );
  OAI21_X1 u0_u0_u7_U10 (.B1( u0_u0_u7_n13 ) , .A( u0_u0_u7_n20 ) , .B2( u0_u0_u7_n8 ) , .ZN( u0_u0_u7_n90 ) );
  AOI211_X1 u0_u0_u7_U11 (.B( u0_u0_u7_n1 ) , .C1( u0_u0_u7_n4 ) , .C2( u0_u0_u7_n55 ) , .ZN( u0_u0_u7_n63 ) , .A( u0_u0_u7_n64 ) );
  OAI22_X1 u0_u0_u7_U12 (.B2( u0_u0_u7_n19 ) , .A1( u0_u0_u7_n44 ) , .A2( u0_u0_u7_n48 ) , .ZN( u0_u0_u7_n64 ) , .B1( u0_u0_u7_n66 ) );
  INV_X1 u0_u0_u7_U13 (.ZN( u0_u0_u7_n1 ) , .A( u0_u0_u7_n65 ) );
  NOR3_X1 u0_u0_u7_U14 (.A1( u0_u0_u7_n12 ) , .A2( u0_u0_u7_n13 ) , .A3( u0_u0_u7_n36 ) , .ZN( u0_u0_u7_n66 ) );
  INV_X1 u0_u0_u7_U15 (.A( u0_u0_u7_n48 ) , .ZN( u0_u0_u7_n5 ) );
  NOR3_X1 u0_u0_u7_U16 (.A3( u0_u0_u7_n10 ) , .ZN( u0_u0_u7_n45 ) , .A1( u0_u0_u7_n46 ) , .A2( u0_u0_u7_n47 ) );
  NOR2_X1 u0_u0_u7_U17 (.ZN( u0_u0_u7_n28 ) , .A2( u0_u0_u7_n47 ) , .A1( u0_u0_u7_n51 ) );
  AOI21_X1 u0_u0_u7_U18 (.A( u0_u0_u7_n17 ) , .B1( u0_u0_u7_n54 ) , .B2( u0_u0_u7_n69 ) , .ZN( u0_u0_u7_n77 ) );
  AOI21_X1 u0_u0_u7_U19 (.A( u0_u0_u7_n19 ) , .B2( u0_u0_u7_n35 ) , .B1( u0_u0_u7_n48 ) , .ZN( u0_u0_u7_n75 ) );
  AOI21_X1 u0_u0_u7_U20 (.B2( u0_u0_u7_n53 ) , .B1( u0_u0_u7_n6 ) , .ZN( u0_u0_u7_n74 ) , .A( u0_u0_u7_n80 ) );
  INV_X1 u0_u0_u7_U21 (.ZN( u0_u0_u7_n16 ) , .A( u0_u0_u7_n80 ) );
  NOR2_X1 u0_u0_u7_U22 (.A1( u0_u0_u7_n12 ) , .A2( u0_u0_u7_n47 ) , .ZN( u0_u0_u7_n70 ) );
  INV_X1 u0_u0_u7_U23 (.ZN( u0_u0_u7_n10 ) , .A( u0_u0_u7_n43 ) );
  INV_X1 u0_u0_u7_U24 (.ZN( u0_u0_u7_n4 ) , .A( u0_u0_u7_n50 ) );
  INV_X1 u0_u0_u7_U25 (.ZN( u0_u0_u7_n7 ) , .A( u0_u0_u7_n71 ) );
  NAND2_X1 u0_u0_u7_U26 (.ZN( u0_u0_u7_n32 ) , .A2( u0_u0_u7_n49 ) , .A1( u0_u0_u7_n52 ) );
  NAND2_X1 u0_u0_u7_U27 (.ZN( u0_u0_u7_n51 ) , .A2( u0_u0_u7_n57 ) , .A1( u0_u0_u7_n68 ) );
  INV_X1 u0_u0_u7_U28 (.A( u0_u0_u7_n69 ) , .ZN( u0_u0_u7_n8 ) );
  INV_X1 u0_u0_u7_U29 (.ZN( u0_u0_u7_n13 ) , .A( u0_u0_u7_n53 ) );
  OAI21_X1 u0_u0_u7_U3 (.B2( u0_u0_u7_n10 ) , .A( u0_u0_u7_n16 ) , .ZN( u0_u0_u7_n22 ) , .B1( u0_u0_u7_n7 ) );
  INV_X1 u0_u0_u7_U30 (.ZN( u0_u0_u7_n12 ) , .A( u0_u0_u7_n33 ) );
  INV_X1 u0_u0_u7_U31 (.ZN( u0_u0_u7_n2 ) , .A( u0_u0_u7_n54 ) );
  INV_X1 u0_u0_u7_U32 (.A( u0_u0_u7_n28 ) , .ZN( u0_u0_u7_n9 ) );
  NOR2_X1 u0_u0_u7_U33 (.A1( u0_u0_u7_n25 ) , .A2( u0_u0_u7_n31 ) , .ZN( u0_u0_u7_n80 ) );
  AOI211_X1 u0_u0_u7_U34 (.C1( u0_u0_u7_n25 ) , .ZN( u0_u0_u7_n39 ) , .C2( u0_u0_u7_n40 ) , .A( u0_u0_u7_n41 ) , .B( u0_u0_u7_n42 ) );
  NAND4_X1 u0_u0_u7_U35 (.A4( u0_u0_u7_n34 ) , .ZN( u0_u0_u7_n40 ) , .A1( u0_u0_u7_n52 ) , .A2( u0_u0_u7_n53 ) , .A3( u0_u0_u7_n54 ) );
  AOI21_X1 u0_u0_u7_U36 (.B2( u0_u0_u7_n35 ) , .ZN( u0_u0_u7_n42 ) , .B1( u0_u0_u7_n43 ) , .A( u0_u0_u7_n44 ) );
  OAI22_X1 u0_u0_u7_U37 (.A2( u0_u0_u7_n17 ) , .B2( u0_u0_u7_n19 ) , .A1( u0_u0_u7_n28 ) , .ZN( u0_u0_u7_n41 ) , .B1( u0_u0_u7_n45 ) );
  INV_X1 u0_u0_u7_U38 (.ZN( u0_u0_u7_n20 ) , .A( u0_u0_u7_n56 ) );
  AOI21_X1 u0_u0_u7_U39 (.B1( u0_u0_u7_n16 ) , .B2( u0_u0_u7_n4 ) , .ZN( u0_u0_u7_n58 ) , .A( u0_u0_u7_n84 ) );
  INV_X1 u0_u0_u7_U4 (.A( u0_u0_u7_n32 ) , .ZN( u0_u0_u7_n6 ) );
  AOI21_X1 u0_u0_u7_U40 (.A( u0_u0_u7_n56 ) , .B1( u0_u0_u7_n57 ) , .B2( u0_u0_u7_n68 ) , .ZN( u0_u0_u7_n84 ) );
  INV_X1 u0_u0_u7_U41 (.ZN( u0_u0_u7_n19 ) , .A( u0_u0_u7_n29 ) );
  AOI22_X1 u0_u0_u7_U42 (.B2( u0_u0_u7_n16 ) , .A1( u0_u0_u7_n25 ) , .B1( u0_u0_u7_n51 ) , .ZN( u0_u0_u7_n62 ) , .A2( u0_u0_u7_n67 ) );
  NAND2_X1 u0_u0_u7_U43 (.A1( u0_u0_u7_n6 ) , .ZN( u0_u0_u7_n67 ) , .A2( u0_u0_u7_n69 ) );
  NOR2_X1 u0_u0_u7_U44 (.A2( u0_u0_u7_n20 ) , .A1( u0_u0_u7_n31 ) , .ZN( u0_u0_u7_n44 ) );
  AND2_X1 u0_u0_u7_U45 (.ZN( u0_u0_u7_n36 ) , .A1( u0_u0_u7_n82 ) , .A2( u0_u0_u7_n83 ) );
  AOI21_X1 u0_u0_u7_U46 (.B1( u0_u0_u7_n34 ) , .A( u0_u0_u7_n56 ) , .B2( u0_u0_u7_n71 ) , .ZN( u0_u0_u7_n76 ) );
  NAND2_X1 u0_u0_u7_U47 (.ZN( u0_u0_u7_n35 ) , .A2( u0_u0_u7_n83 ) , .A1( u0_u0_u7_n86 ) );
  NAND2_X1 u0_u0_u7_U48 (.ZN( u0_u0_u7_n34 ) , .A2( u0_u0_u7_n78 ) , .A1( u0_u0_u7_n88 ) );
  NAND2_X1 u0_u0_u7_U49 (.ZN( u0_u0_u7_n54 ) , .A1( u0_u0_u7_n78 ) , .A2( u0_u0_u7_n82 ) );
  INV_X1 u0_u0_u7_U5 (.A( u0_u0_u7_n27 ) , .ZN( u0_u0_u7_n3 ) );
  NAND2_X1 u0_u0_u7_U50 (.ZN( u0_u0_u7_n48 ) , .A1( u0_u0_u7_n78 ) , .A2( u0_u0_u7_n79 ) );
  OR2_X1 u0_u0_u7_U51 (.A1( u0_u0_u7_n25 ) , .A2( u0_u0_u7_n29 ) , .ZN( u0_u0_u7_n55 ) );
  NAND2_X1 u0_u0_u7_U52 (.ZN( u0_u0_u7_n69 ) , .A1( u0_u0_u7_n82 ) , .A2( u0_u0_u7_n85 ) );
  NAND2_X1 u0_u0_u7_U53 (.ZN( u0_u0_u7_n53 ) , .A2( u0_u0_u7_n79 ) , .A1( u0_u0_u7_n83 ) );
  NAND2_X1 u0_u0_u7_U54 (.ZN( u0_u0_u7_n68 ) , .A1( u0_u0_u7_n81 ) , .A2( u0_u0_u7_n88 ) );
  NAND2_X1 u0_u0_u7_U55 (.ZN( u0_u0_u7_n71 ) , .A2( u0_u0_u7_n85 ) , .A1( u0_u0_u7_n86 ) );
  INV_X1 u0_u0_u7_U56 (.ZN( u0_u0_u7_n17 ) , .A( u0_u0_u7_n31 ) );
  AND2_X1 u0_u0_u7_U57 (.ZN( u0_u0_u7_n47 ) , .A2( u0_u0_u7_n83 ) , .A1( u0_u0_u7_n88 ) );
  NAND2_X1 u0_u0_u7_U58 (.ZN( u0_u0_u7_n57 ) , .A2( u0_u0_u7_n79 ) , .A1( u0_u0_u7_n85 ) );
  NAND2_X1 u0_u0_u7_U59 (.ZN( u0_u0_u7_n52 ) , .A2( u0_u0_u7_n79 ) , .A1( u0_u0_u7_n81 ) );
  AOI211_X1 u0_u0_u7_U6 (.C2( u0_u0_u7_n10 ) , .C1( u0_u0_u7_n20 ) , .A( u0_u0_u7_n26 ) , .ZN( u0_u0_u7_n65 ) , .B( u0_u0_u7_n87 ) );
  NAND2_X1 u0_u0_u7_U60 (.ZN( u0_u0_u7_n50 ) , .A2( u0_u0_u7_n78 ) , .A1( u0_u0_u7_n86 ) );
  NAND2_X1 u0_u0_u7_U61 (.ZN( u0_u0_u7_n43 ) , .A1( u0_u0_u7_n81 ) , .A2( u0_u0_u7_n82 ) );
  NAND2_X1 u0_u0_u7_U62 (.ZN( u0_u0_u7_n49 ) , .A2( u0_u0_u7_n85 ) , .A1( u0_u0_u7_n88 ) );
  NAND2_X1 u0_u0_u7_U63 (.ZN( u0_u0_u7_n33 ) , .A1( u0_u0_u7_n81 ) , .A2( u0_u0_u7_n86 ) );
  NOR2_X1 u0_u0_u7_U64 (.A2( u0_u0_X_47 ) , .A1( u0_u0_u7_n18 ) , .ZN( u0_u0_u7_n31 ) );
  NOR2_X1 u0_u0_u7_U65 (.A2( u0_u0_X_43 ) , .A1( u0_u0_X_44 ) , .ZN( u0_u0_u7_n78 ) );
  NOR2_X1 u0_u0_u7_U66 (.A2( u0_u0_X_48 ) , .A1( u0_u0_u7_n15 ) , .ZN( u0_u0_u7_n86 ) );
  NOR2_X1 u0_u0_u7_U67 (.A2( u0_u0_X_45 ) , .A1( u0_u0_X_48 ) , .ZN( u0_u0_u7_n82 ) );
  NOR2_X1 u0_u0_u7_U68 (.A2( u0_u0_X_44 ) , .A1( u0_u0_u7_n14 ) , .ZN( u0_u0_u7_n83 ) );
  NOR2_X1 u0_u0_u7_U69 (.A2( u0_u0_X_46 ) , .A1( u0_u0_X_47 ) , .ZN( u0_u0_u7_n29 ) );
  OAI222_X1 u0_u0_u7_U7 (.B1( u0_u0_u7_n17 ) , .A2( u0_u0_u7_n19 ) , .C1( u0_u0_u7_n35 ) , .A1( u0_u0_u7_n68 ) , .B2( u0_u0_u7_n70 ) , .C2( u0_u0_u7_n80 ) , .ZN( u0_u0_u7_n87 ) );
  NAND2_X1 u0_u0_u7_U70 (.A2( u0_u0_X_46 ) , .A1( u0_u0_X_47 ) , .ZN( u0_u0_u7_n56 ) );
  AND2_X1 u0_u0_u7_U71 (.A1( u0_u0_X_47 ) , .A2( u0_u0_u7_n18 ) , .ZN( u0_u0_u7_n25 ) );
  AND2_X1 u0_u0_u7_U72 (.A2( u0_u0_X_45 ) , .A1( u0_u0_X_48 ) , .ZN( u0_u0_u7_n79 ) );
  AND2_X1 u0_u0_u7_U73 (.A2( u0_u0_X_43 ) , .A1( u0_u0_X_44 ) , .ZN( u0_u0_u7_n85 ) );
  AND2_X1 u0_u0_u7_U74 (.A1( u0_u0_X_44 ) , .A2( u0_u0_u7_n14 ) , .ZN( u0_u0_u7_n81 ) );
  AND2_X1 u0_u0_u7_U75 (.A1( u0_u0_X_48 ) , .A2( u0_u0_u7_n15 ) , .ZN( u0_u0_u7_n88 ) );
  INV_X1 u0_u0_u7_U76 (.A( u0_u0_X_46 ) , .ZN( u0_u0_u7_n18 ) );
  INV_X1 u0_u0_u7_U77 (.A( u0_u0_X_45 ) , .ZN( u0_u0_u7_n15 ) );
  NAND4_X1 u0_u0_u7_U78 (.ZN( u0_out0_27 ) , .A1( u0_u0_u7_n60 ) , .A2( u0_u0_u7_n61 ) , .A3( u0_u0_u7_n62 ) , .A4( u0_u0_u7_n63 ) );
  OAI21_X1 u0_u0_u7_U79 (.A( u0_u0_u7_n31 ) , .B2( u0_u0_u7_n36 ) , .ZN( u0_u0_u7_n60 ) , .B1( u0_u0_u7_n7 ) );
  OAI221_X1 u0_u0_u7_U8 (.B2( u0_u0_u7_n19 ) , .ZN( u0_u0_u7_n26 ) , .C2( u0_u0_u7_n34 ) , .C1( u0_u0_u7_n80 ) , .B1( u0_u0_u7_n89 ) , .A( u0_u0_u7_n90 ) );
  OAI21_X1 u0_u0_u7_U80 (.B2( u0_u0_u7_n11 ) , .B1( u0_u0_u7_n2 ) , .A( u0_u0_u7_n20 ) , .ZN( u0_u0_u7_n61 ) );
  NAND4_X1 u0_u0_u7_U81 (.ZN( u0_out0_21 ) , .A1( u0_u0_u7_n21 ) , .A2( u0_u0_u7_n22 ) , .A3( u0_u0_u7_n23 ) , .A4( u0_u0_u7_n24 ) );
  OAI21_X1 u0_u0_u7_U82 (.A( u0_u0_u7_n20 ) , .ZN( u0_u0_u7_n21 ) , .B1( u0_u0_u7_n36 ) , .B2( u0_u0_u7_n4 ) );
  AOI22_X1 u0_u0_u7_U83 (.ZN( u0_u0_u7_n23 ) , .A1( u0_u0_u7_n29 ) , .A2( u0_u0_u7_n30 ) , .B1( u0_u0_u7_n31 ) , .B2( u0_u0_u7_n32 ) );
  NAND4_X1 u0_u0_u7_U84 (.ZN( u0_out0_5 ) , .A2( u0_u0_u7_n58 ) , .A1( u0_u0_u7_n65 ) , .A3( u0_u0_u7_n72 ) , .A4( u0_u0_u7_n73 ) );
  AOI22_X1 u0_u0_u7_U85 (.A1( u0_u0_u7_n10 ) , .B1( u0_u0_u7_n25 ) , .B2( u0_u0_u7_n36 ) , .A2( u0_u0_u7_n55 ) , .ZN( u0_u0_u7_n72 ) );
  NOR4_X1 u0_u0_u7_U86 (.ZN( u0_u0_u7_n73 ) , .A1( u0_u0_u7_n74 ) , .A2( u0_u0_u7_n75 ) , .A3( u0_u0_u7_n76 ) , .A4( u0_u0_u7_n77 ) );
  NAND4_X1 u0_u0_u7_U87 (.ZN( u0_out0_15 ) , .A1( u0_u0_u7_n3 ) , .A2( u0_u0_u7_n37 ) , .A3( u0_u0_u7_n38 ) , .A4( u0_u0_u7_n39 ) );
  OR2_X1 u0_u0_u7_U88 (.ZN( u0_u0_u7_n37 ) , .A1( u0_u0_u7_n52 ) , .A2( u0_u0_u7_n56 ) );
  AOI22_X1 u0_u0_u7_U89 (.B2( u0_u0_u7_n16 ) , .ZN( u0_u0_u7_n38 ) , .A2( u0_u0_u7_n55 ) , .A1( u0_u0_u7_n7 ) , .B1( u0_u0_u7_n8 ) );
  AND3_X1 u0_u0_u7_U9 (.A1( u0_u0_u7_n49 ) , .A2( u0_u0_u7_n54 ) , .A3( u0_u0_u7_n71 ) , .ZN( u0_u0_u7_n89 ) );
  INV_X1 u0_u0_u7_U90 (.A( u0_u0_X_43 ) , .ZN( u0_u0_u7_n14 ) );
  AOI211_X1 u0_u0_u7_U91 (.ZN( u0_u0_u7_n24 ) , .C1( u0_u0_u7_n25 ) , .A( u0_u0_u7_n26 ) , .B( u0_u0_u7_n27 ) , .C2( u0_u0_u7_n9 ) );
  OAI211_X1 u0_u0_u7_U92 (.C1( u0_u0_u7_n19 ) , .ZN( u0_u0_u7_n27 ) , .C2( u0_u0_u7_n57 ) , .A( u0_u0_u7_n58 ) , .B( u0_u0_u7_n59 ) );
  AOI222_X1 u0_u0_u7_U93 (.B2( u0_u0_u7_n11 ) , .A2( u0_u0_u7_n16 ) , .B1( u0_u0_u7_n20 ) , .C1( u0_u0_u7_n36 ) , .A1( u0_u0_u7_n5 ) , .C2( u0_u0_u7_n55 ) , .ZN( u0_u0_u7_n59 ) );
  INV_X1 u0_u0_u7_U94 (.ZN( u0_u0_u7_n11 ) , .A( u0_u0_u7_n70 ) );
  NAND3_X1 u0_u0_u7_U95 (.ZN( u0_u0_u7_n30 ) , .A1( u0_u0_u7_n33 ) , .A2( u0_u0_u7_n34 ) , .A3( u0_u0_u7_n35 ) );
  NAND3_X1 u0_u0_u7_U96 (.ZN( u0_u0_u7_n46 ) , .A1( u0_u0_u7_n48 ) , .A2( u0_u0_u7_n49 ) , .A3( u0_u0_u7_n50 ) );
  XOR2_X1 u0_u10_U33 (.B( u0_K11_24 ) , .A( u0_R9_17 ) , .Z( u0_u10_X_24 ) );
  XOR2_X1 u0_u10_U34 (.B( u0_K11_23 ) , .A( u0_R9_16 ) , .Z( u0_u10_X_23 ) );
  XOR2_X1 u0_u10_U35 (.B( u0_K11_22 ) , .A( u0_R9_15 ) , .Z( u0_u10_X_22 ) );
  XOR2_X1 u0_u10_U37 (.B( u0_K11_20 ) , .A( u0_R9_13 ) , .Z( u0_u10_X_20 ) );
  XOR2_X1 u0_u10_U39 (.B( u0_K11_19 ) , .A( u0_R9_12 ) , .Z( u0_u10_X_19 ) );
  XOR2_X1 u0_u10_U40 (.B( u0_K11_18 ) , .A( u0_R9_13 ) , .Z( u0_u10_X_18 ) );
  XOR2_X1 u0_u10_U41 (.B( u0_K11_17 ) , .A( u0_R9_12 ) , .Z( u0_u10_X_17 ) );
  XOR2_X1 u0_u10_U42 (.B( u0_K11_16 ) , .A( u0_R9_11 ) , .Z( u0_u10_X_16 ) );
  XOR2_X1 u0_u10_U43 (.B( u0_K11_15 ) , .A( u0_R9_10 ) , .Z( u0_u10_X_15 ) );
  XOR2_X1 u0_u10_U44 (.B( u0_K11_14 ) , .A( u0_R9_9 ) , .Z( u0_u10_X_14 ) );
  XOR2_X1 u0_u10_U45 (.B( u0_K11_13 ) , .A( u0_R9_8 ) , .Z( u0_u10_X_13 ) );
  OAI22_X1 u0_u10_u2_U10 (.ZN( u0_u10_u2_n109 ) , .A2( u0_u10_u2_n113 ) , .B2( u0_u10_u2_n133 ) , .B1( u0_u10_u2_n167 ) , .A1( u0_u10_u2_n168 ) );
  NAND3_X1 u0_u10_u2_U100 (.A2( u0_u10_u2_n100 ) , .A1( u0_u10_u2_n104 ) , .A3( u0_u10_u2_n138 ) , .ZN( u0_u10_u2_n98 ) );
  OAI22_X1 u0_u10_u2_U11 (.B1( u0_u10_u2_n151 ) , .A2( u0_u10_u2_n152 ) , .A1( u0_u10_u2_n153 ) , .ZN( u0_u10_u2_n160 ) , .B2( u0_u10_u2_n168 ) );
  NOR3_X1 u0_u10_u2_U12 (.A1( u0_u10_u2_n150 ) , .ZN( u0_u10_u2_n151 ) , .A3( u0_u10_u2_n175 ) , .A2( u0_u10_u2_n188 ) );
  AOI21_X1 u0_u10_u2_U13 (.ZN( u0_u10_u2_n144 ) , .B2( u0_u10_u2_n155 ) , .A( u0_u10_u2_n172 ) , .B1( u0_u10_u2_n185 ) );
  AOI21_X1 u0_u10_u2_U14 (.B2( u0_u10_u2_n143 ) , .ZN( u0_u10_u2_n145 ) , .B1( u0_u10_u2_n152 ) , .A( u0_u10_u2_n171 ) );
  AOI21_X1 u0_u10_u2_U15 (.B2( u0_u10_u2_n120 ) , .B1( u0_u10_u2_n121 ) , .ZN( u0_u10_u2_n126 ) , .A( u0_u10_u2_n167 ) );
  INV_X1 u0_u10_u2_U16 (.A( u0_u10_u2_n156 ) , .ZN( u0_u10_u2_n171 ) );
  INV_X1 u0_u10_u2_U17 (.A( u0_u10_u2_n120 ) , .ZN( u0_u10_u2_n188 ) );
  NAND2_X1 u0_u10_u2_U18 (.A2( u0_u10_u2_n122 ) , .ZN( u0_u10_u2_n150 ) , .A1( u0_u10_u2_n152 ) );
  INV_X1 u0_u10_u2_U19 (.A( u0_u10_u2_n153 ) , .ZN( u0_u10_u2_n170 ) );
  INV_X1 u0_u10_u2_U20 (.A( u0_u10_u2_n137 ) , .ZN( u0_u10_u2_n173 ) );
  NAND2_X1 u0_u10_u2_U21 (.A1( u0_u10_u2_n132 ) , .A2( u0_u10_u2_n139 ) , .ZN( u0_u10_u2_n157 ) );
  INV_X1 u0_u10_u2_U22 (.A( u0_u10_u2_n113 ) , .ZN( u0_u10_u2_n178 ) );
  INV_X1 u0_u10_u2_U23 (.A( u0_u10_u2_n139 ) , .ZN( u0_u10_u2_n175 ) );
  INV_X1 u0_u10_u2_U24 (.A( u0_u10_u2_n155 ) , .ZN( u0_u10_u2_n181 ) );
  INV_X1 u0_u10_u2_U25 (.A( u0_u10_u2_n119 ) , .ZN( u0_u10_u2_n177 ) );
  INV_X1 u0_u10_u2_U26 (.A( u0_u10_u2_n116 ) , .ZN( u0_u10_u2_n180 ) );
  INV_X1 u0_u10_u2_U27 (.A( u0_u10_u2_n131 ) , .ZN( u0_u10_u2_n179 ) );
  INV_X1 u0_u10_u2_U28 (.A( u0_u10_u2_n154 ) , .ZN( u0_u10_u2_n176 ) );
  NAND2_X1 u0_u10_u2_U29 (.A2( u0_u10_u2_n116 ) , .A1( u0_u10_u2_n117 ) , .ZN( u0_u10_u2_n118 ) );
  NOR2_X1 u0_u10_u2_U3 (.ZN( u0_u10_u2_n121 ) , .A2( u0_u10_u2_n177 ) , .A1( u0_u10_u2_n180 ) );
  INV_X1 u0_u10_u2_U30 (.A( u0_u10_u2_n132 ) , .ZN( u0_u10_u2_n182 ) );
  INV_X1 u0_u10_u2_U31 (.A( u0_u10_u2_n158 ) , .ZN( u0_u10_u2_n183 ) );
  OAI21_X1 u0_u10_u2_U32 (.A( u0_u10_u2_n156 ) , .B1( u0_u10_u2_n157 ) , .ZN( u0_u10_u2_n158 ) , .B2( u0_u10_u2_n179 ) );
  NOR2_X1 u0_u10_u2_U33 (.ZN( u0_u10_u2_n156 ) , .A1( u0_u10_u2_n166 ) , .A2( u0_u10_u2_n169 ) );
  NOR2_X1 u0_u10_u2_U34 (.A2( u0_u10_u2_n114 ) , .ZN( u0_u10_u2_n137 ) , .A1( u0_u10_u2_n140 ) );
  NOR2_X1 u0_u10_u2_U35 (.A2( u0_u10_u2_n138 ) , .ZN( u0_u10_u2_n153 ) , .A1( u0_u10_u2_n156 ) );
  AOI211_X1 u0_u10_u2_U36 (.ZN( u0_u10_u2_n130 ) , .C1( u0_u10_u2_n138 ) , .C2( u0_u10_u2_n179 ) , .B( u0_u10_u2_n96 ) , .A( u0_u10_u2_n97 ) );
  OAI22_X1 u0_u10_u2_U37 (.B1( u0_u10_u2_n133 ) , .A2( u0_u10_u2_n137 ) , .A1( u0_u10_u2_n152 ) , .B2( u0_u10_u2_n168 ) , .ZN( u0_u10_u2_n97 ) );
  OAI221_X1 u0_u10_u2_U38 (.B1( u0_u10_u2_n113 ) , .C1( u0_u10_u2_n132 ) , .A( u0_u10_u2_n149 ) , .B2( u0_u10_u2_n171 ) , .C2( u0_u10_u2_n172 ) , .ZN( u0_u10_u2_n96 ) );
  OAI221_X1 u0_u10_u2_U39 (.A( u0_u10_u2_n115 ) , .C2( u0_u10_u2_n123 ) , .B2( u0_u10_u2_n143 ) , .B1( u0_u10_u2_n153 ) , .ZN( u0_u10_u2_n163 ) , .C1( u0_u10_u2_n168 ) );
  INV_X1 u0_u10_u2_U4 (.A( u0_u10_u2_n134 ) , .ZN( u0_u10_u2_n185 ) );
  OAI21_X1 u0_u10_u2_U40 (.A( u0_u10_u2_n114 ) , .ZN( u0_u10_u2_n115 ) , .B1( u0_u10_u2_n176 ) , .B2( u0_u10_u2_n178 ) );
  OAI221_X1 u0_u10_u2_U41 (.A( u0_u10_u2_n135 ) , .B2( u0_u10_u2_n136 ) , .B1( u0_u10_u2_n137 ) , .ZN( u0_u10_u2_n162 ) , .C2( u0_u10_u2_n167 ) , .C1( u0_u10_u2_n185 ) );
  AND3_X1 u0_u10_u2_U42 (.A3( u0_u10_u2_n131 ) , .A2( u0_u10_u2_n132 ) , .A1( u0_u10_u2_n133 ) , .ZN( u0_u10_u2_n136 ) );
  AOI22_X1 u0_u10_u2_U43 (.ZN( u0_u10_u2_n135 ) , .B1( u0_u10_u2_n140 ) , .A1( u0_u10_u2_n156 ) , .B2( u0_u10_u2_n180 ) , .A2( u0_u10_u2_n188 ) );
  AOI21_X1 u0_u10_u2_U44 (.ZN( u0_u10_u2_n149 ) , .B1( u0_u10_u2_n173 ) , .B2( u0_u10_u2_n188 ) , .A( u0_u10_u2_n95 ) );
  AND3_X1 u0_u10_u2_U45 (.A2( u0_u10_u2_n100 ) , .A1( u0_u10_u2_n104 ) , .A3( u0_u10_u2_n156 ) , .ZN( u0_u10_u2_n95 ) );
  OAI21_X1 u0_u10_u2_U46 (.A( u0_u10_u2_n141 ) , .B2( u0_u10_u2_n142 ) , .ZN( u0_u10_u2_n146 ) , .B1( u0_u10_u2_n153 ) );
  OAI21_X1 u0_u10_u2_U47 (.A( u0_u10_u2_n140 ) , .ZN( u0_u10_u2_n141 ) , .B1( u0_u10_u2_n176 ) , .B2( u0_u10_u2_n177 ) );
  NOR3_X1 u0_u10_u2_U48 (.ZN( u0_u10_u2_n142 ) , .A3( u0_u10_u2_n175 ) , .A2( u0_u10_u2_n178 ) , .A1( u0_u10_u2_n181 ) );
  OAI21_X1 u0_u10_u2_U49 (.A( u0_u10_u2_n101 ) , .B2( u0_u10_u2_n121 ) , .B1( u0_u10_u2_n153 ) , .ZN( u0_u10_u2_n164 ) );
  INV_X1 u0_u10_u2_U5 (.A( u0_u10_u2_n150 ) , .ZN( u0_u10_u2_n184 ) );
  NAND2_X1 u0_u10_u2_U50 (.A2( u0_u10_u2_n100 ) , .A1( u0_u10_u2_n107 ) , .ZN( u0_u10_u2_n155 ) );
  NAND2_X1 u0_u10_u2_U51 (.A2( u0_u10_u2_n105 ) , .A1( u0_u10_u2_n108 ) , .ZN( u0_u10_u2_n143 ) );
  NAND2_X1 u0_u10_u2_U52 (.A1( u0_u10_u2_n104 ) , .A2( u0_u10_u2_n106 ) , .ZN( u0_u10_u2_n152 ) );
  NAND2_X1 u0_u10_u2_U53 (.A1( u0_u10_u2_n100 ) , .A2( u0_u10_u2_n105 ) , .ZN( u0_u10_u2_n132 ) );
  INV_X1 u0_u10_u2_U54 (.A( u0_u10_u2_n140 ) , .ZN( u0_u10_u2_n168 ) );
  INV_X1 u0_u10_u2_U55 (.A( u0_u10_u2_n138 ) , .ZN( u0_u10_u2_n167 ) );
  NAND2_X1 u0_u10_u2_U56 (.A1( u0_u10_u2_n102 ) , .A2( u0_u10_u2_n106 ) , .ZN( u0_u10_u2_n113 ) );
  NAND2_X1 u0_u10_u2_U57 (.A1( u0_u10_u2_n106 ) , .A2( u0_u10_u2_n107 ) , .ZN( u0_u10_u2_n131 ) );
  NAND2_X1 u0_u10_u2_U58 (.A1( u0_u10_u2_n103 ) , .A2( u0_u10_u2_n107 ) , .ZN( u0_u10_u2_n139 ) );
  NAND2_X1 u0_u10_u2_U59 (.A1( u0_u10_u2_n103 ) , .A2( u0_u10_u2_n105 ) , .ZN( u0_u10_u2_n133 ) );
  NOR4_X1 u0_u10_u2_U6 (.A4( u0_u10_u2_n124 ) , .A3( u0_u10_u2_n125 ) , .A2( u0_u10_u2_n126 ) , .A1( u0_u10_u2_n127 ) , .ZN( u0_u10_u2_n128 ) );
  NAND2_X1 u0_u10_u2_U60 (.A1( u0_u10_u2_n102 ) , .A2( u0_u10_u2_n103 ) , .ZN( u0_u10_u2_n154 ) );
  NAND2_X1 u0_u10_u2_U61 (.A2( u0_u10_u2_n103 ) , .A1( u0_u10_u2_n104 ) , .ZN( u0_u10_u2_n119 ) );
  NAND2_X1 u0_u10_u2_U62 (.A2( u0_u10_u2_n107 ) , .A1( u0_u10_u2_n108 ) , .ZN( u0_u10_u2_n123 ) );
  NAND2_X1 u0_u10_u2_U63 (.A1( u0_u10_u2_n104 ) , .A2( u0_u10_u2_n108 ) , .ZN( u0_u10_u2_n122 ) );
  INV_X1 u0_u10_u2_U64 (.A( u0_u10_u2_n114 ) , .ZN( u0_u10_u2_n172 ) );
  NAND2_X1 u0_u10_u2_U65 (.A2( u0_u10_u2_n100 ) , .A1( u0_u10_u2_n102 ) , .ZN( u0_u10_u2_n116 ) );
  NAND2_X1 u0_u10_u2_U66 (.A1( u0_u10_u2_n102 ) , .A2( u0_u10_u2_n108 ) , .ZN( u0_u10_u2_n120 ) );
  NAND2_X1 u0_u10_u2_U67 (.A2( u0_u10_u2_n105 ) , .A1( u0_u10_u2_n106 ) , .ZN( u0_u10_u2_n117 ) );
  INV_X1 u0_u10_u2_U68 (.ZN( u0_u10_u2_n187 ) , .A( u0_u10_u2_n99 ) );
  OAI21_X1 u0_u10_u2_U69 (.B1( u0_u10_u2_n137 ) , .B2( u0_u10_u2_n143 ) , .A( u0_u10_u2_n98 ) , .ZN( u0_u10_u2_n99 ) );
  AOI21_X1 u0_u10_u2_U7 (.ZN( u0_u10_u2_n124 ) , .B1( u0_u10_u2_n131 ) , .B2( u0_u10_u2_n143 ) , .A( u0_u10_u2_n172 ) );
  NOR2_X1 u0_u10_u2_U70 (.A2( u0_u10_X_16 ) , .ZN( u0_u10_u2_n140 ) , .A1( u0_u10_u2_n166 ) );
  NOR2_X1 u0_u10_u2_U71 (.A2( u0_u10_X_13 ) , .A1( u0_u10_X_14 ) , .ZN( u0_u10_u2_n100 ) );
  NOR2_X1 u0_u10_u2_U72 (.A2( u0_u10_X_16 ) , .A1( u0_u10_X_17 ) , .ZN( u0_u10_u2_n138 ) );
  NOR2_X1 u0_u10_u2_U73 (.A2( u0_u10_X_15 ) , .A1( u0_u10_X_18 ) , .ZN( u0_u10_u2_n104 ) );
  NOR2_X1 u0_u10_u2_U74 (.A2( u0_u10_X_14 ) , .ZN( u0_u10_u2_n103 ) , .A1( u0_u10_u2_n174 ) );
  NOR2_X1 u0_u10_u2_U75 (.A2( u0_u10_X_15 ) , .ZN( u0_u10_u2_n102 ) , .A1( u0_u10_u2_n165 ) );
  NOR2_X1 u0_u10_u2_U76 (.A2( u0_u10_X_17 ) , .ZN( u0_u10_u2_n114 ) , .A1( u0_u10_u2_n169 ) );
  AND2_X1 u0_u10_u2_U77 (.A1( u0_u10_X_15 ) , .ZN( u0_u10_u2_n105 ) , .A2( u0_u10_u2_n165 ) );
  AND2_X1 u0_u10_u2_U78 (.A2( u0_u10_X_15 ) , .A1( u0_u10_X_18 ) , .ZN( u0_u10_u2_n107 ) );
  AND2_X1 u0_u10_u2_U79 (.A1( u0_u10_X_14 ) , .ZN( u0_u10_u2_n106 ) , .A2( u0_u10_u2_n174 ) );
  AOI21_X1 u0_u10_u2_U8 (.B2( u0_u10_u2_n119 ) , .ZN( u0_u10_u2_n127 ) , .A( u0_u10_u2_n137 ) , .B1( u0_u10_u2_n155 ) );
  AND2_X1 u0_u10_u2_U80 (.A1( u0_u10_X_13 ) , .A2( u0_u10_X_14 ) , .ZN( u0_u10_u2_n108 ) );
  INV_X1 u0_u10_u2_U81 (.A( u0_u10_X_16 ) , .ZN( u0_u10_u2_n169 ) );
  INV_X1 u0_u10_u2_U82 (.A( u0_u10_X_17 ) , .ZN( u0_u10_u2_n166 ) );
  INV_X1 u0_u10_u2_U83 (.A( u0_u10_X_13 ) , .ZN( u0_u10_u2_n174 ) );
  INV_X1 u0_u10_u2_U84 (.A( u0_u10_X_18 ) , .ZN( u0_u10_u2_n165 ) );
  NAND4_X1 u0_u10_u2_U85 (.ZN( u0_out10_30 ) , .A4( u0_u10_u2_n147 ) , .A3( u0_u10_u2_n148 ) , .A2( u0_u10_u2_n149 ) , .A1( u0_u10_u2_n187 ) );
  NOR3_X1 u0_u10_u2_U86 (.A3( u0_u10_u2_n144 ) , .A2( u0_u10_u2_n145 ) , .A1( u0_u10_u2_n146 ) , .ZN( u0_u10_u2_n147 ) );
  AOI21_X1 u0_u10_u2_U87 (.B2( u0_u10_u2_n138 ) , .ZN( u0_u10_u2_n148 ) , .A( u0_u10_u2_n162 ) , .B1( u0_u10_u2_n182 ) );
  NAND4_X1 u0_u10_u2_U88 (.ZN( u0_out10_24 ) , .A4( u0_u10_u2_n111 ) , .A3( u0_u10_u2_n112 ) , .A1( u0_u10_u2_n130 ) , .A2( u0_u10_u2_n187 ) );
  AOI221_X1 u0_u10_u2_U89 (.A( u0_u10_u2_n109 ) , .B1( u0_u10_u2_n110 ) , .ZN( u0_u10_u2_n111 ) , .C1( u0_u10_u2_n134 ) , .C2( u0_u10_u2_n170 ) , .B2( u0_u10_u2_n173 ) );
  AOI21_X1 u0_u10_u2_U9 (.B2( u0_u10_u2_n123 ) , .ZN( u0_u10_u2_n125 ) , .A( u0_u10_u2_n171 ) , .B1( u0_u10_u2_n184 ) );
  AOI21_X1 u0_u10_u2_U90 (.ZN( u0_u10_u2_n112 ) , .B2( u0_u10_u2_n156 ) , .A( u0_u10_u2_n164 ) , .B1( u0_u10_u2_n181 ) );
  NAND4_X1 u0_u10_u2_U91 (.ZN( u0_out10_16 ) , .A4( u0_u10_u2_n128 ) , .A3( u0_u10_u2_n129 ) , .A1( u0_u10_u2_n130 ) , .A2( u0_u10_u2_n186 ) );
  AOI22_X1 u0_u10_u2_U92 (.A2( u0_u10_u2_n118 ) , .ZN( u0_u10_u2_n129 ) , .A1( u0_u10_u2_n140 ) , .B1( u0_u10_u2_n157 ) , .B2( u0_u10_u2_n170 ) );
  INV_X1 u0_u10_u2_U93 (.A( u0_u10_u2_n163 ) , .ZN( u0_u10_u2_n186 ) );
  OR4_X1 u0_u10_u2_U94 (.ZN( u0_out10_6 ) , .A4( u0_u10_u2_n161 ) , .A3( u0_u10_u2_n162 ) , .A2( u0_u10_u2_n163 ) , .A1( u0_u10_u2_n164 ) );
  OR3_X1 u0_u10_u2_U95 (.A2( u0_u10_u2_n159 ) , .A1( u0_u10_u2_n160 ) , .ZN( u0_u10_u2_n161 ) , .A3( u0_u10_u2_n183 ) );
  AOI21_X1 u0_u10_u2_U96 (.B2( u0_u10_u2_n154 ) , .B1( u0_u10_u2_n155 ) , .ZN( u0_u10_u2_n159 ) , .A( u0_u10_u2_n167 ) );
  NAND3_X1 u0_u10_u2_U97 (.A2( u0_u10_u2_n117 ) , .A1( u0_u10_u2_n122 ) , .A3( u0_u10_u2_n123 ) , .ZN( u0_u10_u2_n134 ) );
  NAND3_X1 u0_u10_u2_U98 (.ZN( u0_u10_u2_n110 ) , .A2( u0_u10_u2_n131 ) , .A3( u0_u10_u2_n139 ) , .A1( u0_u10_u2_n154 ) );
  NAND3_X1 u0_u10_u2_U99 (.A2( u0_u10_u2_n100 ) , .ZN( u0_u10_u2_n101 ) , .A1( u0_u10_u2_n104 ) , .A3( u0_u10_u2_n114 ) );
  OAI22_X1 u0_u10_u3_U10 (.B1( u0_u10_u3_n113 ) , .A2( u0_u10_u3_n135 ) , .A1( u0_u10_u3_n150 ) , .B2( u0_u10_u3_n164 ) , .ZN( u0_u10_u3_n98 ) );
  OAI211_X1 u0_u10_u3_U11 (.B( u0_u10_u3_n106 ) , .ZN( u0_u10_u3_n119 ) , .C2( u0_u10_u3_n128 ) , .C1( u0_u10_u3_n167 ) , .A( u0_u10_u3_n181 ) );
  AOI221_X1 u0_u10_u3_U12 (.C1( u0_u10_u3_n105 ) , .ZN( u0_u10_u3_n106 ) , .A( u0_u10_u3_n131 ) , .B2( u0_u10_u3_n132 ) , .C2( u0_u10_u3_n133 ) , .B1( u0_u10_u3_n169 ) );
  INV_X1 u0_u10_u3_U13 (.ZN( u0_u10_u3_n181 ) , .A( u0_u10_u3_n98 ) );
  NAND2_X1 u0_u10_u3_U14 (.ZN( u0_u10_u3_n105 ) , .A2( u0_u10_u3_n130 ) , .A1( u0_u10_u3_n155 ) );
  AOI22_X1 u0_u10_u3_U15 (.B1( u0_u10_u3_n115 ) , .A2( u0_u10_u3_n116 ) , .ZN( u0_u10_u3_n123 ) , .B2( u0_u10_u3_n133 ) , .A1( u0_u10_u3_n169 ) );
  NAND2_X1 u0_u10_u3_U16 (.ZN( u0_u10_u3_n116 ) , .A2( u0_u10_u3_n151 ) , .A1( u0_u10_u3_n182 ) );
  NOR2_X1 u0_u10_u3_U17 (.ZN( u0_u10_u3_n126 ) , .A2( u0_u10_u3_n150 ) , .A1( u0_u10_u3_n164 ) );
  AOI21_X1 u0_u10_u3_U18 (.ZN( u0_u10_u3_n112 ) , .B2( u0_u10_u3_n146 ) , .B1( u0_u10_u3_n155 ) , .A( u0_u10_u3_n167 ) );
  NAND2_X1 u0_u10_u3_U19 (.A1( u0_u10_u3_n135 ) , .ZN( u0_u10_u3_n142 ) , .A2( u0_u10_u3_n164 ) );
  NAND2_X1 u0_u10_u3_U20 (.ZN( u0_u10_u3_n132 ) , .A2( u0_u10_u3_n152 ) , .A1( u0_u10_u3_n156 ) );
  AND2_X1 u0_u10_u3_U21 (.A2( u0_u10_u3_n113 ) , .A1( u0_u10_u3_n114 ) , .ZN( u0_u10_u3_n151 ) );
  INV_X1 u0_u10_u3_U22 (.A( u0_u10_u3_n133 ) , .ZN( u0_u10_u3_n165 ) );
  INV_X1 u0_u10_u3_U23 (.A( u0_u10_u3_n135 ) , .ZN( u0_u10_u3_n170 ) );
  NAND2_X1 u0_u10_u3_U24 (.A1( u0_u10_u3_n107 ) , .A2( u0_u10_u3_n108 ) , .ZN( u0_u10_u3_n140 ) );
  NAND2_X1 u0_u10_u3_U25 (.ZN( u0_u10_u3_n117 ) , .A1( u0_u10_u3_n124 ) , .A2( u0_u10_u3_n148 ) );
  NAND2_X1 u0_u10_u3_U26 (.ZN( u0_u10_u3_n143 ) , .A1( u0_u10_u3_n165 ) , .A2( u0_u10_u3_n167 ) );
  INV_X1 u0_u10_u3_U27 (.A( u0_u10_u3_n130 ) , .ZN( u0_u10_u3_n177 ) );
  INV_X1 u0_u10_u3_U28 (.A( u0_u10_u3_n128 ) , .ZN( u0_u10_u3_n176 ) );
  INV_X1 u0_u10_u3_U29 (.A( u0_u10_u3_n155 ) , .ZN( u0_u10_u3_n174 ) );
  INV_X1 u0_u10_u3_U3 (.A( u0_u10_u3_n129 ) , .ZN( u0_u10_u3_n183 ) );
  INV_X1 u0_u10_u3_U30 (.A( u0_u10_u3_n139 ) , .ZN( u0_u10_u3_n185 ) );
  NOR2_X1 u0_u10_u3_U31 (.ZN( u0_u10_u3_n135 ) , .A2( u0_u10_u3_n141 ) , .A1( u0_u10_u3_n169 ) );
  OAI222_X1 u0_u10_u3_U32 (.C2( u0_u10_u3_n107 ) , .A2( u0_u10_u3_n108 ) , .B1( u0_u10_u3_n135 ) , .ZN( u0_u10_u3_n138 ) , .B2( u0_u10_u3_n146 ) , .C1( u0_u10_u3_n154 ) , .A1( u0_u10_u3_n164 ) );
  NOR4_X1 u0_u10_u3_U33 (.A4( u0_u10_u3_n157 ) , .A3( u0_u10_u3_n158 ) , .A2( u0_u10_u3_n159 ) , .A1( u0_u10_u3_n160 ) , .ZN( u0_u10_u3_n161 ) );
  AOI21_X1 u0_u10_u3_U34 (.B2( u0_u10_u3_n152 ) , .B1( u0_u10_u3_n153 ) , .ZN( u0_u10_u3_n158 ) , .A( u0_u10_u3_n164 ) );
  AOI21_X1 u0_u10_u3_U35 (.A( u0_u10_u3_n154 ) , .B2( u0_u10_u3_n155 ) , .B1( u0_u10_u3_n156 ) , .ZN( u0_u10_u3_n157 ) );
  AOI21_X1 u0_u10_u3_U36 (.A( u0_u10_u3_n149 ) , .B2( u0_u10_u3_n150 ) , .B1( u0_u10_u3_n151 ) , .ZN( u0_u10_u3_n159 ) );
  AOI211_X1 u0_u10_u3_U37 (.ZN( u0_u10_u3_n109 ) , .A( u0_u10_u3_n119 ) , .C2( u0_u10_u3_n129 ) , .B( u0_u10_u3_n138 ) , .C1( u0_u10_u3_n141 ) );
  AOI211_X1 u0_u10_u3_U38 (.B( u0_u10_u3_n119 ) , .A( u0_u10_u3_n120 ) , .C2( u0_u10_u3_n121 ) , .ZN( u0_u10_u3_n122 ) , .C1( u0_u10_u3_n179 ) );
  INV_X1 u0_u10_u3_U39 (.A( u0_u10_u3_n156 ) , .ZN( u0_u10_u3_n179 ) );
  INV_X1 u0_u10_u3_U4 (.A( u0_u10_u3_n140 ) , .ZN( u0_u10_u3_n182 ) );
  OAI22_X1 u0_u10_u3_U40 (.B1( u0_u10_u3_n118 ) , .ZN( u0_u10_u3_n120 ) , .A1( u0_u10_u3_n135 ) , .B2( u0_u10_u3_n154 ) , .A2( u0_u10_u3_n178 ) );
  AND3_X1 u0_u10_u3_U41 (.ZN( u0_u10_u3_n118 ) , .A2( u0_u10_u3_n124 ) , .A1( u0_u10_u3_n144 ) , .A3( u0_u10_u3_n152 ) );
  INV_X1 u0_u10_u3_U42 (.A( u0_u10_u3_n121 ) , .ZN( u0_u10_u3_n164 ) );
  NAND2_X1 u0_u10_u3_U43 (.ZN( u0_u10_u3_n133 ) , .A1( u0_u10_u3_n154 ) , .A2( u0_u10_u3_n164 ) );
  OAI211_X1 u0_u10_u3_U44 (.B( u0_u10_u3_n127 ) , .ZN( u0_u10_u3_n139 ) , .C1( u0_u10_u3_n150 ) , .C2( u0_u10_u3_n154 ) , .A( u0_u10_u3_n184 ) );
  INV_X1 u0_u10_u3_U45 (.A( u0_u10_u3_n125 ) , .ZN( u0_u10_u3_n184 ) );
  AOI221_X1 u0_u10_u3_U46 (.A( u0_u10_u3_n126 ) , .ZN( u0_u10_u3_n127 ) , .C2( u0_u10_u3_n132 ) , .C1( u0_u10_u3_n169 ) , .B2( u0_u10_u3_n170 ) , .B1( u0_u10_u3_n174 ) );
  OAI22_X1 u0_u10_u3_U47 (.A1( u0_u10_u3_n124 ) , .ZN( u0_u10_u3_n125 ) , .B2( u0_u10_u3_n145 ) , .A2( u0_u10_u3_n165 ) , .B1( u0_u10_u3_n167 ) );
  NOR2_X1 u0_u10_u3_U48 (.A1( u0_u10_u3_n113 ) , .ZN( u0_u10_u3_n131 ) , .A2( u0_u10_u3_n154 ) );
  NAND2_X1 u0_u10_u3_U49 (.A1( u0_u10_u3_n103 ) , .ZN( u0_u10_u3_n150 ) , .A2( u0_u10_u3_n99 ) );
  INV_X1 u0_u10_u3_U5 (.A( u0_u10_u3_n117 ) , .ZN( u0_u10_u3_n178 ) );
  NAND2_X1 u0_u10_u3_U50 (.A2( u0_u10_u3_n102 ) , .ZN( u0_u10_u3_n155 ) , .A1( u0_u10_u3_n97 ) );
  INV_X1 u0_u10_u3_U51 (.A( u0_u10_u3_n141 ) , .ZN( u0_u10_u3_n167 ) );
  AOI21_X1 u0_u10_u3_U52 (.B2( u0_u10_u3_n114 ) , .B1( u0_u10_u3_n146 ) , .A( u0_u10_u3_n154 ) , .ZN( u0_u10_u3_n94 ) );
  AOI21_X1 u0_u10_u3_U53 (.ZN( u0_u10_u3_n110 ) , .B2( u0_u10_u3_n142 ) , .B1( u0_u10_u3_n186 ) , .A( u0_u10_u3_n95 ) );
  INV_X1 u0_u10_u3_U54 (.A( u0_u10_u3_n145 ) , .ZN( u0_u10_u3_n186 ) );
  AOI21_X1 u0_u10_u3_U55 (.B1( u0_u10_u3_n124 ) , .A( u0_u10_u3_n149 ) , .B2( u0_u10_u3_n155 ) , .ZN( u0_u10_u3_n95 ) );
  INV_X1 u0_u10_u3_U56 (.A( u0_u10_u3_n149 ) , .ZN( u0_u10_u3_n169 ) );
  NAND2_X1 u0_u10_u3_U57 (.ZN( u0_u10_u3_n124 ) , .A1( u0_u10_u3_n96 ) , .A2( u0_u10_u3_n97 ) );
  NAND2_X1 u0_u10_u3_U58 (.A2( u0_u10_u3_n100 ) , .ZN( u0_u10_u3_n146 ) , .A1( u0_u10_u3_n96 ) );
  NAND2_X1 u0_u10_u3_U59 (.A1( u0_u10_u3_n101 ) , .ZN( u0_u10_u3_n145 ) , .A2( u0_u10_u3_n99 ) );
  AOI221_X1 u0_u10_u3_U6 (.A( u0_u10_u3_n131 ) , .C2( u0_u10_u3_n132 ) , .C1( u0_u10_u3_n133 ) , .ZN( u0_u10_u3_n134 ) , .B1( u0_u10_u3_n143 ) , .B2( u0_u10_u3_n177 ) );
  NAND2_X1 u0_u10_u3_U60 (.A1( u0_u10_u3_n100 ) , .ZN( u0_u10_u3_n156 ) , .A2( u0_u10_u3_n99 ) );
  NAND2_X1 u0_u10_u3_U61 (.A2( u0_u10_u3_n101 ) , .A1( u0_u10_u3_n104 ) , .ZN( u0_u10_u3_n148 ) );
  NAND2_X1 u0_u10_u3_U62 (.A1( u0_u10_u3_n100 ) , .A2( u0_u10_u3_n102 ) , .ZN( u0_u10_u3_n128 ) );
  NAND2_X1 u0_u10_u3_U63 (.A2( u0_u10_u3_n101 ) , .A1( u0_u10_u3_n102 ) , .ZN( u0_u10_u3_n152 ) );
  NAND2_X1 u0_u10_u3_U64 (.A2( u0_u10_u3_n101 ) , .ZN( u0_u10_u3_n114 ) , .A1( u0_u10_u3_n96 ) );
  NAND2_X1 u0_u10_u3_U65 (.ZN( u0_u10_u3_n107 ) , .A1( u0_u10_u3_n97 ) , .A2( u0_u10_u3_n99 ) );
  NAND2_X1 u0_u10_u3_U66 (.A2( u0_u10_u3_n100 ) , .A1( u0_u10_u3_n104 ) , .ZN( u0_u10_u3_n113 ) );
  NAND2_X1 u0_u10_u3_U67 (.A1( u0_u10_u3_n104 ) , .ZN( u0_u10_u3_n153 ) , .A2( u0_u10_u3_n97 ) );
  NAND2_X1 u0_u10_u3_U68 (.A2( u0_u10_u3_n103 ) , .A1( u0_u10_u3_n104 ) , .ZN( u0_u10_u3_n130 ) );
  NAND2_X1 u0_u10_u3_U69 (.A2( u0_u10_u3_n103 ) , .ZN( u0_u10_u3_n144 ) , .A1( u0_u10_u3_n96 ) );
  OAI22_X1 u0_u10_u3_U7 (.B2( u0_u10_u3_n147 ) , .A2( u0_u10_u3_n148 ) , .ZN( u0_u10_u3_n160 ) , .B1( u0_u10_u3_n165 ) , .A1( u0_u10_u3_n168 ) );
  NAND2_X1 u0_u10_u3_U70 (.A1( u0_u10_u3_n102 ) , .A2( u0_u10_u3_n103 ) , .ZN( u0_u10_u3_n108 ) );
  NOR2_X1 u0_u10_u3_U71 (.A2( u0_u10_X_19 ) , .A1( u0_u10_X_20 ) , .ZN( u0_u10_u3_n99 ) );
  NOR2_X1 u0_u10_u3_U72 (.A2( u0_u10_X_21 ) , .A1( u0_u10_X_24 ) , .ZN( u0_u10_u3_n103 ) );
  NOR2_X1 u0_u10_u3_U73 (.A2( u0_u10_X_24 ) , .A1( u0_u10_u3_n171 ) , .ZN( u0_u10_u3_n97 ) );
  NOR2_X1 u0_u10_u3_U74 (.A2( u0_u10_X_23 ) , .ZN( u0_u10_u3_n141 ) , .A1( u0_u10_u3_n166 ) );
  NOR2_X1 u0_u10_u3_U75 (.A2( u0_u10_X_19 ) , .A1( u0_u10_u3_n172 ) , .ZN( u0_u10_u3_n96 ) );
  NAND2_X1 u0_u10_u3_U76 (.A1( u0_u10_X_22 ) , .A2( u0_u10_X_23 ) , .ZN( u0_u10_u3_n154 ) );
  NAND2_X1 u0_u10_u3_U77 (.A1( u0_u10_X_23 ) , .ZN( u0_u10_u3_n149 ) , .A2( u0_u10_u3_n166 ) );
  NOR2_X1 u0_u10_u3_U78 (.A2( u0_u10_X_22 ) , .A1( u0_u10_X_23 ) , .ZN( u0_u10_u3_n121 ) );
  AND2_X1 u0_u10_u3_U79 (.A1( u0_u10_X_24 ) , .ZN( u0_u10_u3_n101 ) , .A2( u0_u10_u3_n171 ) );
  AND3_X1 u0_u10_u3_U8 (.A3( u0_u10_u3_n144 ) , .A2( u0_u10_u3_n145 ) , .A1( u0_u10_u3_n146 ) , .ZN( u0_u10_u3_n147 ) );
  AND2_X1 u0_u10_u3_U80 (.A1( u0_u10_X_19 ) , .ZN( u0_u10_u3_n102 ) , .A2( u0_u10_u3_n172 ) );
  AND2_X1 u0_u10_u3_U81 (.A1( u0_u10_X_21 ) , .A2( u0_u10_X_24 ) , .ZN( u0_u10_u3_n100 ) );
  AND2_X1 u0_u10_u3_U82 (.A2( u0_u10_X_19 ) , .A1( u0_u10_X_20 ) , .ZN( u0_u10_u3_n104 ) );
  INV_X1 u0_u10_u3_U83 (.A( u0_u10_X_22 ) , .ZN( u0_u10_u3_n166 ) );
  INV_X1 u0_u10_u3_U84 (.A( u0_u10_X_21 ) , .ZN( u0_u10_u3_n171 ) );
  INV_X1 u0_u10_u3_U85 (.A( u0_u10_X_20 ) , .ZN( u0_u10_u3_n172 ) );
  OR4_X1 u0_u10_u3_U86 (.ZN( u0_out10_10 ) , .A4( u0_u10_u3_n136 ) , .A3( u0_u10_u3_n137 ) , .A1( u0_u10_u3_n138 ) , .A2( u0_u10_u3_n139 ) );
  OAI222_X1 u0_u10_u3_U87 (.C1( u0_u10_u3_n128 ) , .ZN( u0_u10_u3_n137 ) , .B1( u0_u10_u3_n148 ) , .A2( u0_u10_u3_n150 ) , .B2( u0_u10_u3_n154 ) , .C2( u0_u10_u3_n164 ) , .A1( u0_u10_u3_n167 ) );
  OAI221_X1 u0_u10_u3_U88 (.A( u0_u10_u3_n134 ) , .B2( u0_u10_u3_n135 ) , .ZN( u0_u10_u3_n136 ) , .C1( u0_u10_u3_n149 ) , .B1( u0_u10_u3_n151 ) , .C2( u0_u10_u3_n183 ) );
  NAND4_X1 u0_u10_u3_U89 (.ZN( u0_out10_26 ) , .A4( u0_u10_u3_n109 ) , .A3( u0_u10_u3_n110 ) , .A2( u0_u10_u3_n111 ) , .A1( u0_u10_u3_n173 ) );
  INV_X1 u0_u10_u3_U9 (.A( u0_u10_u3_n143 ) , .ZN( u0_u10_u3_n168 ) );
  INV_X1 u0_u10_u3_U90 (.ZN( u0_u10_u3_n173 ) , .A( u0_u10_u3_n94 ) );
  OAI21_X1 u0_u10_u3_U91 (.ZN( u0_u10_u3_n111 ) , .B2( u0_u10_u3_n117 ) , .A( u0_u10_u3_n133 ) , .B1( u0_u10_u3_n176 ) );
  NAND4_X1 u0_u10_u3_U92 (.ZN( u0_out10_20 ) , .A4( u0_u10_u3_n122 ) , .A3( u0_u10_u3_n123 ) , .A1( u0_u10_u3_n175 ) , .A2( u0_u10_u3_n180 ) );
  INV_X1 u0_u10_u3_U93 (.A( u0_u10_u3_n126 ) , .ZN( u0_u10_u3_n180 ) );
  INV_X1 u0_u10_u3_U94 (.A( u0_u10_u3_n112 ) , .ZN( u0_u10_u3_n175 ) );
  NAND4_X1 u0_u10_u3_U95 (.ZN( u0_out10_1 ) , .A4( u0_u10_u3_n161 ) , .A3( u0_u10_u3_n162 ) , .A2( u0_u10_u3_n163 ) , .A1( u0_u10_u3_n185 ) );
  NAND2_X1 u0_u10_u3_U96 (.ZN( u0_u10_u3_n163 ) , .A2( u0_u10_u3_n170 ) , .A1( u0_u10_u3_n176 ) );
  AOI22_X1 u0_u10_u3_U97 (.B2( u0_u10_u3_n140 ) , .B1( u0_u10_u3_n141 ) , .A2( u0_u10_u3_n142 ) , .ZN( u0_u10_u3_n162 ) , .A1( u0_u10_u3_n177 ) );
  NAND3_X1 u0_u10_u3_U98 (.A1( u0_u10_u3_n114 ) , .ZN( u0_u10_u3_n115 ) , .A2( u0_u10_u3_n145 ) , .A3( u0_u10_u3_n153 ) );
  NAND3_X1 u0_u10_u3_U99 (.ZN( u0_u10_u3_n129 ) , .A2( u0_u10_u3_n144 ) , .A1( u0_u10_u3_n153 ) , .A3( u0_u10_u3_n182 ) );
  XOR2_X1 u0_u12_U1 (.B( u0_K13_9 ) , .A( u0_R11_6 ) , .Z( u0_u12_X_9 ) );
  XOR2_X1 u0_u12_U12 (.B( u0_K13_43 ) , .A( u0_R11_28 ) , .Z( u0_u12_X_43 ) );
  XOR2_X1 u0_u12_U2 (.B( u0_K13_8 ) , .A( u0_R11_5 ) , .Z( u0_u12_X_8 ) );
  XOR2_X1 u0_u12_U3 (.B( u0_K13_7 ) , .A( u0_R11_4 ) , .Z( u0_u12_X_7 ) );
  XOR2_X1 u0_u12_U38 (.B( u0_K13_1 ) , .A( u0_R11_32 ) , .Z( u0_u12_X_1 ) );
  XOR2_X1 u0_u12_U4 (.B( u0_K13_6 ) , .A( u0_R11_5 ) , .Z( u0_u12_X_6 ) );
  XOR2_X1 u0_u12_U46 (.B( u0_K13_12 ) , .A( u0_R11_9 ) , .Z( u0_u12_X_12 ) );
  XOR2_X1 u0_u12_U47 (.B( u0_K13_11 ) , .A( u0_R11_8 ) , .Z( u0_u12_X_11 ) );
  XOR2_X1 u0_u12_U48 (.B( u0_K13_10 ) , .A( u0_R11_7 ) , .Z( u0_u12_X_10 ) );
  XOR2_X1 u0_u12_U5 (.B( u0_K13_5 ) , .A( u0_R11_4 ) , .Z( u0_u12_X_5 ) );
  XOR2_X1 u0_u12_U6 (.B( u0_K13_4 ) , .A( u0_R11_3 ) , .Z( u0_u12_X_4 ) );
  XOR2_X1 u0_u12_U8 (.B( u0_K13_47 ) , .A( u0_R11_32 ) , .Z( u0_u12_X_47 ) );
  NAND2_X1 u0_u12_u0_U10 (.ZN( u0_u12_u0_n113 ) , .A1( u0_u12_u0_n139 ) , .A2( u0_u12_u0_n149 ) );
  AND3_X1 u0_u12_u0_U11 (.A2( u0_u12_u0_n112 ) , .ZN( u0_u12_u0_n127 ) , .A3( u0_u12_u0_n130 ) , .A1( u0_u12_u0_n148 ) );
  AND2_X1 u0_u12_u0_U12 (.ZN( u0_u12_u0_n107 ) , .A1( u0_u12_u0_n130 ) , .A2( u0_u12_u0_n140 ) );
  AND2_X1 u0_u12_u0_U13 (.A2( u0_u12_u0_n129 ) , .A1( u0_u12_u0_n130 ) , .ZN( u0_u12_u0_n151 ) );
  AND2_X1 u0_u12_u0_U14 (.A1( u0_u12_u0_n108 ) , .A2( u0_u12_u0_n125 ) , .ZN( u0_u12_u0_n145 ) );
  INV_X1 u0_u12_u0_U15 (.A( u0_u12_u0_n143 ) , .ZN( u0_u12_u0_n173 ) );
  NOR2_X1 u0_u12_u0_U16 (.A2( u0_u12_u0_n136 ) , .ZN( u0_u12_u0_n147 ) , .A1( u0_u12_u0_n160 ) );
  AOI21_X1 u0_u12_u0_U17 (.B1( u0_u12_u0_n103 ) , .ZN( u0_u12_u0_n132 ) , .A( u0_u12_u0_n165 ) , .B2( u0_u12_u0_n93 ) );
  INV_X1 u0_u12_u0_U18 (.A( u0_u12_u0_n142 ) , .ZN( u0_u12_u0_n165 ) );
  OAI22_X1 u0_u12_u0_U19 (.B1( u0_u12_u0_n131 ) , .A1( u0_u12_u0_n144 ) , .B2( u0_u12_u0_n147 ) , .A2( u0_u12_u0_n90 ) , .ZN( u0_u12_u0_n91 ) );
  AND3_X1 u0_u12_u0_U20 (.A3( u0_u12_u0_n121 ) , .A2( u0_u12_u0_n125 ) , .A1( u0_u12_u0_n148 ) , .ZN( u0_u12_u0_n90 ) );
  OAI22_X1 u0_u12_u0_U21 (.B1( u0_u12_u0_n125 ) , .ZN( u0_u12_u0_n126 ) , .A1( u0_u12_u0_n138 ) , .A2( u0_u12_u0_n146 ) , .B2( u0_u12_u0_n147 ) );
  INV_X1 u0_u12_u0_U22 (.A( u0_u12_u0_n136 ) , .ZN( u0_u12_u0_n161 ) );
  AOI22_X1 u0_u12_u0_U23 (.B2( u0_u12_u0_n109 ) , .A2( u0_u12_u0_n110 ) , .ZN( u0_u12_u0_n111 ) , .B1( u0_u12_u0_n118 ) , .A1( u0_u12_u0_n160 ) );
  NAND2_X1 u0_u12_u0_U24 (.A2( u0_u12_u0_n103 ) , .ZN( u0_u12_u0_n140 ) , .A1( u0_u12_u0_n94 ) );
  NAND2_X1 u0_u12_u0_U25 (.A2( u0_u12_u0_n102 ) , .A1( u0_u12_u0_n103 ) , .ZN( u0_u12_u0_n149 ) );
  INV_X1 u0_u12_u0_U26 (.A( u0_u12_u0_n118 ) , .ZN( u0_u12_u0_n158 ) );
  NAND2_X1 u0_u12_u0_U27 (.A2( u0_u12_u0_n100 ) , .ZN( u0_u12_u0_n131 ) , .A1( u0_u12_u0_n92 ) );
  NAND2_X1 u0_u12_u0_U28 (.ZN( u0_u12_u0_n108 ) , .A1( u0_u12_u0_n92 ) , .A2( u0_u12_u0_n94 ) );
  AOI21_X1 u0_u12_u0_U29 (.ZN( u0_u12_u0_n104 ) , .B1( u0_u12_u0_n107 ) , .B2( u0_u12_u0_n141 ) , .A( u0_u12_u0_n144 ) );
  INV_X1 u0_u12_u0_U3 (.A( u0_u12_u0_n113 ) , .ZN( u0_u12_u0_n166 ) );
  AOI21_X1 u0_u12_u0_U30 (.ZN( u0_u12_u0_n116 ) , .B2( u0_u12_u0_n142 ) , .A( u0_u12_u0_n144 ) , .B1( u0_u12_u0_n166 ) );
  AOI21_X1 u0_u12_u0_U31 (.B1( u0_u12_u0_n127 ) , .B2( u0_u12_u0_n129 ) , .A( u0_u12_u0_n138 ) , .ZN( u0_u12_u0_n96 ) );
  NAND2_X1 u0_u12_u0_U32 (.A2( u0_u12_u0_n102 ) , .ZN( u0_u12_u0_n114 ) , .A1( u0_u12_u0_n92 ) );
  NOR2_X1 u0_u12_u0_U33 (.A1( u0_u12_u0_n120 ) , .ZN( u0_u12_u0_n143 ) , .A2( u0_u12_u0_n167 ) );
  OAI221_X1 u0_u12_u0_U34 (.C1( u0_u12_u0_n112 ) , .ZN( u0_u12_u0_n120 ) , .B1( u0_u12_u0_n138 ) , .B2( u0_u12_u0_n141 ) , .C2( u0_u12_u0_n147 ) , .A( u0_u12_u0_n172 ) );
  AOI211_X1 u0_u12_u0_U35 (.B( u0_u12_u0_n115 ) , .A( u0_u12_u0_n116 ) , .C2( u0_u12_u0_n117 ) , .C1( u0_u12_u0_n118 ) , .ZN( u0_u12_u0_n119 ) );
  NAND2_X1 u0_u12_u0_U36 (.A1( u0_u12_u0_n100 ) , .A2( u0_u12_u0_n103 ) , .ZN( u0_u12_u0_n125 ) );
  NAND2_X1 u0_u12_u0_U37 (.A1( u0_u12_u0_n101 ) , .A2( u0_u12_u0_n102 ) , .ZN( u0_u12_u0_n150 ) );
  INV_X1 u0_u12_u0_U38 (.A( u0_u12_u0_n138 ) , .ZN( u0_u12_u0_n160 ) );
  NAND2_X1 u0_u12_u0_U39 (.A2( u0_u12_u0_n100 ) , .A1( u0_u12_u0_n101 ) , .ZN( u0_u12_u0_n139 ) );
  AOI21_X1 u0_u12_u0_U4 (.B1( u0_u12_u0_n114 ) , .ZN( u0_u12_u0_n115 ) , .B2( u0_u12_u0_n129 ) , .A( u0_u12_u0_n161 ) );
  NAND2_X1 u0_u12_u0_U40 (.A1( u0_u12_u0_n101 ) , .ZN( u0_u12_u0_n130 ) , .A2( u0_u12_u0_n94 ) );
  NAND2_X1 u0_u12_u0_U41 (.ZN( u0_u12_u0_n112 ) , .A2( u0_u12_u0_n92 ) , .A1( u0_u12_u0_n93 ) );
  INV_X1 u0_u12_u0_U42 (.ZN( u0_u12_u0_n172 ) , .A( u0_u12_u0_n88 ) );
  OAI222_X1 u0_u12_u0_U43 (.C1( u0_u12_u0_n108 ) , .A1( u0_u12_u0_n125 ) , .B2( u0_u12_u0_n128 ) , .B1( u0_u12_u0_n144 ) , .A2( u0_u12_u0_n158 ) , .C2( u0_u12_u0_n161 ) , .ZN( u0_u12_u0_n88 ) );
  NAND2_X1 u0_u12_u0_U44 (.A2( u0_u12_u0_n101 ) , .ZN( u0_u12_u0_n121 ) , .A1( u0_u12_u0_n93 ) );
  OR3_X1 u0_u12_u0_U45 (.A3( u0_u12_u0_n152 ) , .A2( u0_u12_u0_n153 ) , .A1( u0_u12_u0_n154 ) , .ZN( u0_u12_u0_n155 ) );
  AOI21_X1 u0_u12_u0_U46 (.A( u0_u12_u0_n144 ) , .B2( u0_u12_u0_n145 ) , .B1( u0_u12_u0_n146 ) , .ZN( u0_u12_u0_n154 ) );
  AOI21_X1 u0_u12_u0_U47 (.B2( u0_u12_u0_n150 ) , .B1( u0_u12_u0_n151 ) , .ZN( u0_u12_u0_n152 ) , .A( u0_u12_u0_n158 ) );
  AOI21_X1 u0_u12_u0_U48 (.A( u0_u12_u0_n147 ) , .B2( u0_u12_u0_n148 ) , .B1( u0_u12_u0_n149 ) , .ZN( u0_u12_u0_n153 ) );
  INV_X1 u0_u12_u0_U49 (.ZN( u0_u12_u0_n171 ) , .A( u0_u12_u0_n99 ) );
  AOI21_X1 u0_u12_u0_U5 (.B2( u0_u12_u0_n131 ) , .ZN( u0_u12_u0_n134 ) , .B1( u0_u12_u0_n151 ) , .A( u0_u12_u0_n158 ) );
  OAI211_X1 u0_u12_u0_U50 (.C2( u0_u12_u0_n140 ) , .C1( u0_u12_u0_n161 ) , .A( u0_u12_u0_n169 ) , .B( u0_u12_u0_n98 ) , .ZN( u0_u12_u0_n99 ) );
  INV_X1 u0_u12_u0_U51 (.ZN( u0_u12_u0_n169 ) , .A( u0_u12_u0_n91 ) );
  AOI211_X1 u0_u12_u0_U52 (.C1( u0_u12_u0_n118 ) , .A( u0_u12_u0_n123 ) , .B( u0_u12_u0_n96 ) , .C2( u0_u12_u0_n97 ) , .ZN( u0_u12_u0_n98 ) );
  NOR2_X1 u0_u12_u0_U53 (.A2( u0_u12_X_4 ) , .A1( u0_u12_X_5 ) , .ZN( u0_u12_u0_n118 ) );
  NOR2_X1 u0_u12_u0_U54 (.A2( u0_u12_X_1 ) , .ZN( u0_u12_u0_n101 ) , .A1( u0_u12_u0_n163 ) );
  NOR2_X1 u0_u12_u0_U55 (.A2( u0_u12_X_6 ) , .ZN( u0_u12_u0_n100 ) , .A1( u0_u12_u0_n162 ) );
  NAND2_X1 u0_u12_u0_U56 (.A2( u0_u12_X_4 ) , .A1( u0_u12_X_5 ) , .ZN( u0_u12_u0_n144 ) );
  NOR2_X1 u0_u12_u0_U57 (.A2( u0_u12_X_5 ) , .ZN( u0_u12_u0_n136 ) , .A1( u0_u12_u0_n159 ) );
  NAND2_X1 u0_u12_u0_U58 (.A1( u0_u12_X_5 ) , .ZN( u0_u12_u0_n138 ) , .A2( u0_u12_u0_n159 ) );
  AND2_X1 u0_u12_u0_U59 (.A2( u0_u12_X_3 ) , .A1( u0_u12_X_6 ) , .ZN( u0_u12_u0_n102 ) );
  NOR2_X1 u0_u12_u0_U6 (.A1( u0_u12_u0_n108 ) , .ZN( u0_u12_u0_n123 ) , .A2( u0_u12_u0_n158 ) );
  AND2_X1 u0_u12_u0_U60 (.A1( u0_u12_X_6 ) , .A2( u0_u12_u0_n162 ) , .ZN( u0_u12_u0_n93 ) );
  INV_X1 u0_u12_u0_U61 (.A( u0_u12_X_4 ) , .ZN( u0_u12_u0_n159 ) );
  INV_X1 u0_u12_u0_U62 (.A( u0_u12_X_3 ) , .ZN( u0_u12_u0_n162 ) );
  INV_X1 u0_u12_u0_U63 (.A( u0_u12_u0_n126 ) , .ZN( u0_u12_u0_n168 ) );
  AOI211_X1 u0_u12_u0_U64 (.B( u0_u12_u0_n133 ) , .A( u0_u12_u0_n134 ) , .C2( u0_u12_u0_n135 ) , .C1( u0_u12_u0_n136 ) , .ZN( u0_u12_u0_n137 ) );
  OR4_X1 u0_u12_u0_U65 (.ZN( u0_out12_17 ) , .A4( u0_u12_u0_n122 ) , .A2( u0_u12_u0_n123 ) , .A1( u0_u12_u0_n124 ) , .A3( u0_u12_u0_n170 ) );
  AOI21_X1 u0_u12_u0_U66 (.B2( u0_u12_u0_n107 ) , .ZN( u0_u12_u0_n124 ) , .B1( u0_u12_u0_n128 ) , .A( u0_u12_u0_n161 ) );
  INV_X1 u0_u12_u0_U67 (.A( u0_u12_u0_n111 ) , .ZN( u0_u12_u0_n170 ) );
  OR4_X1 u0_u12_u0_U68 (.ZN( u0_out12_31 ) , .A4( u0_u12_u0_n155 ) , .A2( u0_u12_u0_n156 ) , .A1( u0_u12_u0_n157 ) , .A3( u0_u12_u0_n173 ) );
  AOI21_X1 u0_u12_u0_U69 (.A( u0_u12_u0_n138 ) , .B2( u0_u12_u0_n139 ) , .B1( u0_u12_u0_n140 ) , .ZN( u0_u12_u0_n157 ) );
  OAI21_X1 u0_u12_u0_U7 (.B1( u0_u12_u0_n150 ) , .B2( u0_u12_u0_n158 ) , .A( u0_u12_u0_n172 ) , .ZN( u0_u12_u0_n89 ) );
  AOI21_X1 u0_u12_u0_U70 (.B2( u0_u12_u0_n141 ) , .B1( u0_u12_u0_n142 ) , .ZN( u0_u12_u0_n156 ) , .A( u0_u12_u0_n161 ) );
  INV_X1 u0_u12_u0_U71 (.ZN( u0_u12_u0_n174 ) , .A( u0_u12_u0_n89 ) );
  AOI211_X1 u0_u12_u0_U72 (.B( u0_u12_u0_n104 ) , .A( u0_u12_u0_n105 ) , .ZN( u0_u12_u0_n106 ) , .C2( u0_u12_u0_n113 ) , .C1( u0_u12_u0_n160 ) );
  AND2_X1 u0_u12_u0_U73 (.A2( u0_u12_X_1 ) , .A1( u0_u12_X_2 ) , .ZN( u0_u12_u0_n95 ) );
  INV_X1 u0_u12_u0_U74 (.A( u0_u12_X_1 ) , .ZN( u0_u12_u0_n164 ) );
  NOR2_X1 u0_u12_u0_U75 (.A2( u0_u12_X_3 ) , .A1( u0_u12_X_6 ) , .ZN( u0_u12_u0_n94 ) );
  OAI221_X1 u0_u12_u0_U76 (.C1( u0_u12_u0_n121 ) , .ZN( u0_u12_u0_n122 ) , .B2( u0_u12_u0_n127 ) , .A( u0_u12_u0_n143 ) , .B1( u0_u12_u0_n144 ) , .C2( u0_u12_u0_n147 ) );
  AOI21_X1 u0_u12_u0_U77 (.B1( u0_u12_u0_n132 ) , .ZN( u0_u12_u0_n133 ) , .A( u0_u12_u0_n144 ) , .B2( u0_u12_u0_n166 ) );
  OAI22_X1 u0_u12_u0_U78 (.ZN( u0_u12_u0_n105 ) , .A2( u0_u12_u0_n132 ) , .B1( u0_u12_u0_n146 ) , .A1( u0_u12_u0_n147 ) , .B2( u0_u12_u0_n161 ) );
  NAND2_X1 u0_u12_u0_U79 (.ZN( u0_u12_u0_n110 ) , .A2( u0_u12_u0_n132 ) , .A1( u0_u12_u0_n145 ) );
  AND2_X1 u0_u12_u0_U8 (.A1( u0_u12_u0_n114 ) , .A2( u0_u12_u0_n121 ) , .ZN( u0_u12_u0_n146 ) );
  INV_X1 u0_u12_u0_U80 (.A( u0_u12_u0_n119 ) , .ZN( u0_u12_u0_n167 ) );
  NAND2_X1 u0_u12_u0_U81 (.ZN( u0_u12_u0_n148 ) , .A1( u0_u12_u0_n93 ) , .A2( u0_u12_u0_n95 ) );
  NAND2_X1 u0_u12_u0_U82 (.A1( u0_u12_u0_n100 ) , .ZN( u0_u12_u0_n129 ) , .A2( u0_u12_u0_n95 ) );
  NAND2_X1 u0_u12_u0_U83 (.A1( u0_u12_u0_n102 ) , .ZN( u0_u12_u0_n128 ) , .A2( u0_u12_u0_n95 ) );
  NOR2_X1 u0_u12_u0_U84 (.A2( u0_u12_X_1 ) , .A1( u0_u12_X_2 ) , .ZN( u0_u12_u0_n92 ) );
  NAND2_X1 u0_u12_u0_U85 (.ZN( u0_u12_u0_n142 ) , .A1( u0_u12_u0_n94 ) , .A2( u0_u12_u0_n95 ) );
  NOR2_X1 u0_u12_u0_U86 (.A2( u0_u12_X_2 ) , .ZN( u0_u12_u0_n103 ) , .A1( u0_u12_u0_n164 ) );
  INV_X1 u0_u12_u0_U87 (.A( u0_u12_X_2 ) , .ZN( u0_u12_u0_n163 ) );
  NAND3_X1 u0_u12_u0_U88 (.ZN( u0_out12_23 ) , .A3( u0_u12_u0_n137 ) , .A1( u0_u12_u0_n168 ) , .A2( u0_u12_u0_n171 ) );
  NAND3_X1 u0_u12_u0_U89 (.A3( u0_u12_u0_n127 ) , .A2( u0_u12_u0_n128 ) , .ZN( u0_u12_u0_n135 ) , .A1( u0_u12_u0_n150 ) );
  AND2_X1 u0_u12_u0_U9 (.A1( u0_u12_u0_n131 ) , .ZN( u0_u12_u0_n141 ) , .A2( u0_u12_u0_n150 ) );
  NAND3_X1 u0_u12_u0_U90 (.ZN( u0_u12_u0_n117 ) , .A3( u0_u12_u0_n132 ) , .A2( u0_u12_u0_n139 ) , .A1( u0_u12_u0_n148 ) );
  NAND3_X1 u0_u12_u0_U91 (.ZN( u0_u12_u0_n109 ) , .A2( u0_u12_u0_n114 ) , .A3( u0_u12_u0_n140 ) , .A1( u0_u12_u0_n149 ) );
  NAND3_X1 u0_u12_u0_U92 (.ZN( u0_out12_9 ) , .A3( u0_u12_u0_n106 ) , .A2( u0_u12_u0_n171 ) , .A1( u0_u12_u0_n174 ) );
  NAND3_X1 u0_u12_u0_U93 (.A2( u0_u12_u0_n128 ) , .A1( u0_u12_u0_n132 ) , .A3( u0_u12_u0_n146 ) , .ZN( u0_u12_u0_n97 ) );
  NOR2_X1 u0_u12_u1_U10 (.A1( u0_u12_u1_n112 ) , .A2( u0_u12_u1_n116 ) , .ZN( u0_u12_u1_n118 ) );
  NAND3_X1 u0_u12_u1_U100 (.ZN( u0_u12_u1_n113 ) , .A1( u0_u12_u1_n120 ) , .A3( u0_u12_u1_n133 ) , .A2( u0_u12_u1_n155 ) );
  OAI21_X1 u0_u12_u1_U11 (.ZN( u0_u12_u1_n101 ) , .B1( u0_u12_u1_n141 ) , .A( u0_u12_u1_n146 ) , .B2( u0_u12_u1_n183 ) );
  AOI21_X1 u0_u12_u1_U12 (.B2( u0_u12_u1_n155 ) , .B1( u0_u12_u1_n156 ) , .ZN( u0_u12_u1_n157 ) , .A( u0_u12_u1_n174 ) );
  OR4_X1 u0_u12_u1_U13 (.A4( u0_u12_u1_n106 ) , .A3( u0_u12_u1_n107 ) , .ZN( u0_u12_u1_n108 ) , .A1( u0_u12_u1_n117 ) , .A2( u0_u12_u1_n184 ) );
  AOI21_X1 u0_u12_u1_U14 (.ZN( u0_u12_u1_n106 ) , .A( u0_u12_u1_n112 ) , .B1( u0_u12_u1_n154 ) , .B2( u0_u12_u1_n156 ) );
  INV_X1 u0_u12_u1_U15 (.A( u0_u12_u1_n101 ) , .ZN( u0_u12_u1_n184 ) );
  AOI21_X1 u0_u12_u1_U16 (.ZN( u0_u12_u1_n107 ) , .B1( u0_u12_u1_n134 ) , .B2( u0_u12_u1_n149 ) , .A( u0_u12_u1_n174 ) );
  NAND2_X1 u0_u12_u1_U17 (.ZN( u0_u12_u1_n140 ) , .A2( u0_u12_u1_n150 ) , .A1( u0_u12_u1_n155 ) );
  NAND2_X1 u0_u12_u1_U18 (.A1( u0_u12_u1_n131 ) , .ZN( u0_u12_u1_n147 ) , .A2( u0_u12_u1_n153 ) );
  INV_X1 u0_u12_u1_U19 (.A( u0_u12_u1_n139 ) , .ZN( u0_u12_u1_n174 ) );
  INV_X1 u0_u12_u1_U20 (.A( u0_u12_u1_n112 ) , .ZN( u0_u12_u1_n171 ) );
  NAND2_X1 u0_u12_u1_U21 (.ZN( u0_u12_u1_n141 ) , .A1( u0_u12_u1_n153 ) , .A2( u0_u12_u1_n156 ) );
  AND2_X1 u0_u12_u1_U22 (.A1( u0_u12_u1_n123 ) , .ZN( u0_u12_u1_n134 ) , .A2( u0_u12_u1_n161 ) );
  NAND2_X1 u0_u12_u1_U23 (.A2( u0_u12_u1_n115 ) , .A1( u0_u12_u1_n116 ) , .ZN( u0_u12_u1_n148 ) );
  NAND2_X1 u0_u12_u1_U24 (.A2( u0_u12_u1_n133 ) , .A1( u0_u12_u1_n135 ) , .ZN( u0_u12_u1_n159 ) );
  NAND2_X1 u0_u12_u1_U25 (.A2( u0_u12_u1_n115 ) , .A1( u0_u12_u1_n120 ) , .ZN( u0_u12_u1_n132 ) );
  INV_X1 u0_u12_u1_U26 (.A( u0_u12_u1_n154 ) , .ZN( u0_u12_u1_n178 ) );
  INV_X1 u0_u12_u1_U27 (.A( u0_u12_u1_n151 ) , .ZN( u0_u12_u1_n183 ) );
  AND2_X1 u0_u12_u1_U28 (.A1( u0_u12_u1_n129 ) , .A2( u0_u12_u1_n133 ) , .ZN( u0_u12_u1_n149 ) );
  INV_X1 u0_u12_u1_U29 (.A( u0_u12_u1_n131 ) , .ZN( u0_u12_u1_n180 ) );
  INV_X1 u0_u12_u1_U3 (.A( u0_u12_u1_n159 ) , .ZN( u0_u12_u1_n182 ) );
  AOI221_X1 u0_u12_u1_U30 (.B1( u0_u12_u1_n140 ) , .ZN( u0_u12_u1_n167 ) , .B2( u0_u12_u1_n172 ) , .C2( u0_u12_u1_n175 ) , .C1( u0_u12_u1_n178 ) , .A( u0_u12_u1_n188 ) );
  INV_X1 u0_u12_u1_U31 (.ZN( u0_u12_u1_n188 ) , .A( u0_u12_u1_n97 ) );
  AOI211_X1 u0_u12_u1_U32 (.A( u0_u12_u1_n118 ) , .C1( u0_u12_u1_n132 ) , .C2( u0_u12_u1_n139 ) , .B( u0_u12_u1_n96 ) , .ZN( u0_u12_u1_n97 ) );
  AOI21_X1 u0_u12_u1_U33 (.B2( u0_u12_u1_n121 ) , .B1( u0_u12_u1_n135 ) , .A( u0_u12_u1_n152 ) , .ZN( u0_u12_u1_n96 ) );
  OAI221_X1 u0_u12_u1_U34 (.A( u0_u12_u1_n119 ) , .C2( u0_u12_u1_n129 ) , .ZN( u0_u12_u1_n138 ) , .B2( u0_u12_u1_n152 ) , .C1( u0_u12_u1_n174 ) , .B1( u0_u12_u1_n187 ) );
  INV_X1 u0_u12_u1_U35 (.A( u0_u12_u1_n148 ) , .ZN( u0_u12_u1_n187 ) );
  AOI211_X1 u0_u12_u1_U36 (.B( u0_u12_u1_n117 ) , .A( u0_u12_u1_n118 ) , .ZN( u0_u12_u1_n119 ) , .C2( u0_u12_u1_n146 ) , .C1( u0_u12_u1_n159 ) );
  NOR2_X1 u0_u12_u1_U37 (.A1( u0_u12_u1_n168 ) , .A2( u0_u12_u1_n176 ) , .ZN( u0_u12_u1_n98 ) );
  AOI211_X1 u0_u12_u1_U38 (.B( u0_u12_u1_n162 ) , .A( u0_u12_u1_n163 ) , .C2( u0_u12_u1_n164 ) , .ZN( u0_u12_u1_n165 ) , .C1( u0_u12_u1_n171 ) );
  AOI21_X1 u0_u12_u1_U39 (.A( u0_u12_u1_n160 ) , .B2( u0_u12_u1_n161 ) , .ZN( u0_u12_u1_n162 ) , .B1( u0_u12_u1_n182 ) );
  AOI221_X1 u0_u12_u1_U4 (.A( u0_u12_u1_n138 ) , .C2( u0_u12_u1_n139 ) , .C1( u0_u12_u1_n140 ) , .B2( u0_u12_u1_n141 ) , .ZN( u0_u12_u1_n142 ) , .B1( u0_u12_u1_n175 ) );
  OR2_X1 u0_u12_u1_U40 (.A2( u0_u12_u1_n157 ) , .A1( u0_u12_u1_n158 ) , .ZN( u0_u12_u1_n163 ) );
  NAND2_X1 u0_u12_u1_U41 (.A1( u0_u12_u1_n128 ) , .ZN( u0_u12_u1_n146 ) , .A2( u0_u12_u1_n160 ) );
  NAND2_X1 u0_u12_u1_U42 (.A2( u0_u12_u1_n112 ) , .ZN( u0_u12_u1_n139 ) , .A1( u0_u12_u1_n152 ) );
  NAND2_X1 u0_u12_u1_U43 (.A1( u0_u12_u1_n105 ) , .ZN( u0_u12_u1_n156 ) , .A2( u0_u12_u1_n99 ) );
  NOR2_X1 u0_u12_u1_U44 (.ZN( u0_u12_u1_n117 ) , .A1( u0_u12_u1_n121 ) , .A2( u0_u12_u1_n160 ) );
  OAI21_X1 u0_u12_u1_U45 (.B2( u0_u12_u1_n123 ) , .ZN( u0_u12_u1_n145 ) , .B1( u0_u12_u1_n160 ) , .A( u0_u12_u1_n185 ) );
  INV_X1 u0_u12_u1_U46 (.A( u0_u12_u1_n122 ) , .ZN( u0_u12_u1_n185 ) );
  AOI21_X1 u0_u12_u1_U47 (.B2( u0_u12_u1_n120 ) , .B1( u0_u12_u1_n121 ) , .ZN( u0_u12_u1_n122 ) , .A( u0_u12_u1_n128 ) );
  AOI21_X1 u0_u12_u1_U48 (.A( u0_u12_u1_n128 ) , .B2( u0_u12_u1_n129 ) , .ZN( u0_u12_u1_n130 ) , .B1( u0_u12_u1_n150 ) );
  NAND2_X1 u0_u12_u1_U49 (.ZN( u0_u12_u1_n112 ) , .A1( u0_u12_u1_n169 ) , .A2( u0_u12_u1_n170 ) );
  AOI211_X1 u0_u12_u1_U5 (.ZN( u0_u12_u1_n124 ) , .A( u0_u12_u1_n138 ) , .C2( u0_u12_u1_n139 ) , .B( u0_u12_u1_n145 ) , .C1( u0_u12_u1_n147 ) );
  NAND2_X1 u0_u12_u1_U50 (.ZN( u0_u12_u1_n129 ) , .A2( u0_u12_u1_n95 ) , .A1( u0_u12_u1_n98 ) );
  NAND2_X1 u0_u12_u1_U51 (.A1( u0_u12_u1_n102 ) , .ZN( u0_u12_u1_n154 ) , .A2( u0_u12_u1_n99 ) );
  NAND2_X1 u0_u12_u1_U52 (.A2( u0_u12_u1_n100 ) , .ZN( u0_u12_u1_n135 ) , .A1( u0_u12_u1_n99 ) );
  AOI21_X1 u0_u12_u1_U53 (.A( u0_u12_u1_n152 ) , .B2( u0_u12_u1_n153 ) , .B1( u0_u12_u1_n154 ) , .ZN( u0_u12_u1_n158 ) );
  INV_X1 u0_u12_u1_U54 (.A( u0_u12_u1_n160 ) , .ZN( u0_u12_u1_n175 ) );
  NAND2_X1 u0_u12_u1_U55 (.A1( u0_u12_u1_n100 ) , .ZN( u0_u12_u1_n116 ) , .A2( u0_u12_u1_n95 ) );
  NAND2_X1 u0_u12_u1_U56 (.A1( u0_u12_u1_n102 ) , .ZN( u0_u12_u1_n131 ) , .A2( u0_u12_u1_n95 ) );
  NAND2_X1 u0_u12_u1_U57 (.A2( u0_u12_u1_n104 ) , .ZN( u0_u12_u1_n121 ) , .A1( u0_u12_u1_n98 ) );
  NAND2_X1 u0_u12_u1_U58 (.A1( u0_u12_u1_n103 ) , .ZN( u0_u12_u1_n153 ) , .A2( u0_u12_u1_n98 ) );
  NAND2_X1 u0_u12_u1_U59 (.A2( u0_u12_u1_n104 ) , .A1( u0_u12_u1_n105 ) , .ZN( u0_u12_u1_n133 ) );
  AOI22_X1 u0_u12_u1_U6 (.B2( u0_u12_u1_n113 ) , .A2( u0_u12_u1_n114 ) , .ZN( u0_u12_u1_n125 ) , .A1( u0_u12_u1_n171 ) , .B1( u0_u12_u1_n173 ) );
  NAND2_X1 u0_u12_u1_U60 (.ZN( u0_u12_u1_n150 ) , .A2( u0_u12_u1_n98 ) , .A1( u0_u12_u1_n99 ) );
  NAND2_X1 u0_u12_u1_U61 (.A1( u0_u12_u1_n105 ) , .ZN( u0_u12_u1_n155 ) , .A2( u0_u12_u1_n95 ) );
  OAI21_X1 u0_u12_u1_U62 (.ZN( u0_u12_u1_n109 ) , .B1( u0_u12_u1_n129 ) , .B2( u0_u12_u1_n160 ) , .A( u0_u12_u1_n167 ) );
  NAND2_X1 u0_u12_u1_U63 (.A2( u0_u12_u1_n100 ) , .A1( u0_u12_u1_n103 ) , .ZN( u0_u12_u1_n120 ) );
  NAND2_X1 u0_u12_u1_U64 (.A1( u0_u12_u1_n102 ) , .A2( u0_u12_u1_n104 ) , .ZN( u0_u12_u1_n115 ) );
  NAND2_X1 u0_u12_u1_U65 (.A2( u0_u12_u1_n100 ) , .A1( u0_u12_u1_n104 ) , .ZN( u0_u12_u1_n151 ) );
  NAND2_X1 u0_u12_u1_U66 (.A2( u0_u12_u1_n103 ) , .A1( u0_u12_u1_n105 ) , .ZN( u0_u12_u1_n161 ) );
  INV_X1 u0_u12_u1_U67 (.A( u0_u12_u1_n152 ) , .ZN( u0_u12_u1_n173 ) );
  INV_X1 u0_u12_u1_U68 (.A( u0_u12_u1_n128 ) , .ZN( u0_u12_u1_n172 ) );
  NAND2_X1 u0_u12_u1_U69 (.A2( u0_u12_u1_n102 ) , .A1( u0_u12_u1_n103 ) , .ZN( u0_u12_u1_n123 ) );
  NAND2_X1 u0_u12_u1_U7 (.ZN( u0_u12_u1_n114 ) , .A1( u0_u12_u1_n134 ) , .A2( u0_u12_u1_n156 ) );
  NOR2_X1 u0_u12_u1_U70 (.A2( u0_u12_X_7 ) , .A1( u0_u12_X_8 ) , .ZN( u0_u12_u1_n95 ) );
  NOR2_X1 u0_u12_u1_U71 (.A1( u0_u12_X_12 ) , .A2( u0_u12_X_9 ) , .ZN( u0_u12_u1_n100 ) );
  NOR2_X1 u0_u12_u1_U72 (.A2( u0_u12_X_8 ) , .A1( u0_u12_u1_n177 ) , .ZN( u0_u12_u1_n99 ) );
  NOR2_X1 u0_u12_u1_U73 (.A2( u0_u12_X_12 ) , .ZN( u0_u12_u1_n102 ) , .A1( u0_u12_u1_n176 ) );
  NOR2_X1 u0_u12_u1_U74 (.A2( u0_u12_X_9 ) , .ZN( u0_u12_u1_n105 ) , .A1( u0_u12_u1_n168 ) );
  NAND2_X1 u0_u12_u1_U75 (.A1( u0_u12_X_10 ) , .ZN( u0_u12_u1_n160 ) , .A2( u0_u12_u1_n169 ) );
  NAND2_X1 u0_u12_u1_U76 (.A2( u0_u12_X_10 ) , .A1( u0_u12_X_11 ) , .ZN( u0_u12_u1_n152 ) );
  NAND2_X1 u0_u12_u1_U77 (.A1( u0_u12_X_11 ) , .ZN( u0_u12_u1_n128 ) , .A2( u0_u12_u1_n170 ) );
  AND2_X1 u0_u12_u1_U78 (.A2( u0_u12_X_7 ) , .A1( u0_u12_X_8 ) , .ZN( u0_u12_u1_n104 ) );
  AND2_X1 u0_u12_u1_U79 (.A1( u0_u12_X_8 ) , .ZN( u0_u12_u1_n103 ) , .A2( u0_u12_u1_n177 ) );
  AOI22_X1 u0_u12_u1_U8 (.B2( u0_u12_u1_n136 ) , .A2( u0_u12_u1_n137 ) , .ZN( u0_u12_u1_n143 ) , .A1( u0_u12_u1_n171 ) , .B1( u0_u12_u1_n173 ) );
  INV_X1 u0_u12_u1_U80 (.A( u0_u12_X_10 ) , .ZN( u0_u12_u1_n170 ) );
  INV_X1 u0_u12_u1_U81 (.A( u0_u12_X_9 ) , .ZN( u0_u12_u1_n176 ) );
  INV_X1 u0_u12_u1_U82 (.A( u0_u12_X_11 ) , .ZN( u0_u12_u1_n169 ) );
  INV_X1 u0_u12_u1_U83 (.A( u0_u12_X_12 ) , .ZN( u0_u12_u1_n168 ) );
  INV_X1 u0_u12_u1_U84 (.A( u0_u12_X_7 ) , .ZN( u0_u12_u1_n177 ) );
  NAND4_X1 u0_u12_u1_U85 (.ZN( u0_out12_28 ) , .A4( u0_u12_u1_n124 ) , .A3( u0_u12_u1_n125 ) , .A2( u0_u12_u1_n126 ) , .A1( u0_u12_u1_n127 ) );
  OAI21_X1 u0_u12_u1_U86 (.ZN( u0_u12_u1_n127 ) , .B2( u0_u12_u1_n139 ) , .B1( u0_u12_u1_n175 ) , .A( u0_u12_u1_n183 ) );
  OAI21_X1 u0_u12_u1_U87 (.ZN( u0_u12_u1_n126 ) , .B2( u0_u12_u1_n140 ) , .A( u0_u12_u1_n146 ) , .B1( u0_u12_u1_n178 ) );
  NAND4_X1 u0_u12_u1_U88 (.ZN( u0_out12_18 ) , .A4( u0_u12_u1_n165 ) , .A3( u0_u12_u1_n166 ) , .A1( u0_u12_u1_n167 ) , .A2( u0_u12_u1_n186 ) );
  AOI22_X1 u0_u12_u1_U89 (.B2( u0_u12_u1_n146 ) , .B1( u0_u12_u1_n147 ) , .A2( u0_u12_u1_n148 ) , .ZN( u0_u12_u1_n166 ) , .A1( u0_u12_u1_n172 ) );
  INV_X1 u0_u12_u1_U9 (.A( u0_u12_u1_n147 ) , .ZN( u0_u12_u1_n181 ) );
  INV_X1 u0_u12_u1_U90 (.A( u0_u12_u1_n145 ) , .ZN( u0_u12_u1_n186 ) );
  NAND4_X1 u0_u12_u1_U91 (.ZN( u0_out12_2 ) , .A4( u0_u12_u1_n142 ) , .A3( u0_u12_u1_n143 ) , .A2( u0_u12_u1_n144 ) , .A1( u0_u12_u1_n179 ) );
  OAI21_X1 u0_u12_u1_U92 (.B2( u0_u12_u1_n132 ) , .ZN( u0_u12_u1_n144 ) , .A( u0_u12_u1_n146 ) , .B1( u0_u12_u1_n180 ) );
  INV_X1 u0_u12_u1_U93 (.A( u0_u12_u1_n130 ) , .ZN( u0_u12_u1_n179 ) );
  OR4_X1 u0_u12_u1_U94 (.ZN( u0_out12_13 ) , .A4( u0_u12_u1_n108 ) , .A3( u0_u12_u1_n109 ) , .A2( u0_u12_u1_n110 ) , .A1( u0_u12_u1_n111 ) );
  AOI21_X1 u0_u12_u1_U95 (.ZN( u0_u12_u1_n111 ) , .A( u0_u12_u1_n128 ) , .B2( u0_u12_u1_n131 ) , .B1( u0_u12_u1_n135 ) );
  AOI21_X1 u0_u12_u1_U96 (.ZN( u0_u12_u1_n110 ) , .A( u0_u12_u1_n116 ) , .B1( u0_u12_u1_n152 ) , .B2( u0_u12_u1_n160 ) );
  NAND3_X1 u0_u12_u1_U97 (.A3( u0_u12_u1_n149 ) , .A2( u0_u12_u1_n150 ) , .A1( u0_u12_u1_n151 ) , .ZN( u0_u12_u1_n164 ) );
  NAND3_X1 u0_u12_u1_U98 (.A3( u0_u12_u1_n134 ) , .A2( u0_u12_u1_n135 ) , .ZN( u0_u12_u1_n136 ) , .A1( u0_u12_u1_n151 ) );
  NAND3_X1 u0_u12_u1_U99 (.A1( u0_u12_u1_n133 ) , .ZN( u0_u12_u1_n137 ) , .A2( u0_u12_u1_n154 ) , .A3( u0_u12_u1_n181 ) );
  AND3_X1 u0_u12_u7_U10 (.A3( u0_u12_u7_n110 ) , .A2( u0_u12_u7_n127 ) , .A1( u0_u12_u7_n132 ) , .ZN( u0_u12_u7_n92 ) );
  OAI21_X1 u0_u12_u7_U11 (.A( u0_u12_u7_n161 ) , .B1( u0_u12_u7_n168 ) , .B2( u0_u12_u7_n173 ) , .ZN( u0_u12_u7_n91 ) );
  AOI211_X1 u0_u12_u7_U12 (.A( u0_u12_u7_n117 ) , .ZN( u0_u12_u7_n118 ) , .C2( u0_u12_u7_n126 ) , .C1( u0_u12_u7_n177 ) , .B( u0_u12_u7_n180 ) );
  OAI22_X1 u0_u12_u7_U13 (.B1( u0_u12_u7_n115 ) , .ZN( u0_u12_u7_n117 ) , .A2( u0_u12_u7_n133 ) , .A1( u0_u12_u7_n137 ) , .B2( u0_u12_u7_n162 ) );
  INV_X1 u0_u12_u7_U14 (.A( u0_u12_u7_n116 ) , .ZN( u0_u12_u7_n180 ) );
  NOR3_X1 u0_u12_u7_U15 (.ZN( u0_u12_u7_n115 ) , .A3( u0_u12_u7_n145 ) , .A2( u0_u12_u7_n168 ) , .A1( u0_u12_u7_n169 ) );
  OAI211_X1 u0_u12_u7_U16 (.B( u0_u12_u7_n122 ) , .A( u0_u12_u7_n123 ) , .C2( u0_u12_u7_n124 ) , .ZN( u0_u12_u7_n154 ) , .C1( u0_u12_u7_n162 ) );
  AOI222_X1 u0_u12_u7_U17 (.ZN( u0_u12_u7_n122 ) , .C2( u0_u12_u7_n126 ) , .C1( u0_u12_u7_n145 ) , .B1( u0_u12_u7_n161 ) , .A2( u0_u12_u7_n165 ) , .B2( u0_u12_u7_n170 ) , .A1( u0_u12_u7_n176 ) );
  INV_X1 u0_u12_u7_U18 (.A( u0_u12_u7_n133 ) , .ZN( u0_u12_u7_n176 ) );
  NOR3_X1 u0_u12_u7_U19 (.A2( u0_u12_u7_n134 ) , .A1( u0_u12_u7_n135 ) , .ZN( u0_u12_u7_n136 ) , .A3( u0_u12_u7_n171 ) );
  NOR2_X1 u0_u12_u7_U20 (.A1( u0_u12_u7_n130 ) , .A2( u0_u12_u7_n134 ) , .ZN( u0_u12_u7_n153 ) );
  INV_X1 u0_u12_u7_U21 (.A( u0_u12_u7_n101 ) , .ZN( u0_u12_u7_n165 ) );
  NOR2_X1 u0_u12_u7_U22 (.ZN( u0_u12_u7_n111 ) , .A2( u0_u12_u7_n134 ) , .A1( u0_u12_u7_n169 ) );
  AOI21_X1 u0_u12_u7_U23 (.ZN( u0_u12_u7_n104 ) , .B2( u0_u12_u7_n112 ) , .B1( u0_u12_u7_n127 ) , .A( u0_u12_u7_n164 ) );
  AOI21_X1 u0_u12_u7_U24 (.ZN( u0_u12_u7_n106 ) , .B1( u0_u12_u7_n133 ) , .B2( u0_u12_u7_n146 ) , .A( u0_u12_u7_n162 ) );
  AOI21_X1 u0_u12_u7_U25 (.A( u0_u12_u7_n101 ) , .ZN( u0_u12_u7_n107 ) , .B2( u0_u12_u7_n128 ) , .B1( u0_u12_u7_n175 ) );
  INV_X1 u0_u12_u7_U26 (.A( u0_u12_u7_n138 ) , .ZN( u0_u12_u7_n171 ) );
  INV_X1 u0_u12_u7_U27 (.A( u0_u12_u7_n131 ) , .ZN( u0_u12_u7_n177 ) );
  INV_X1 u0_u12_u7_U28 (.A( u0_u12_u7_n110 ) , .ZN( u0_u12_u7_n174 ) );
  NAND2_X1 u0_u12_u7_U29 (.A1( u0_u12_u7_n129 ) , .A2( u0_u12_u7_n132 ) , .ZN( u0_u12_u7_n149 ) );
  OAI21_X1 u0_u12_u7_U3 (.ZN( u0_u12_u7_n159 ) , .A( u0_u12_u7_n165 ) , .B2( u0_u12_u7_n171 ) , .B1( u0_u12_u7_n174 ) );
  NAND2_X1 u0_u12_u7_U30 (.A1( u0_u12_u7_n113 ) , .A2( u0_u12_u7_n124 ) , .ZN( u0_u12_u7_n130 ) );
  INV_X1 u0_u12_u7_U31 (.A( u0_u12_u7_n112 ) , .ZN( u0_u12_u7_n173 ) );
  INV_X1 u0_u12_u7_U32 (.A( u0_u12_u7_n128 ) , .ZN( u0_u12_u7_n168 ) );
  INV_X1 u0_u12_u7_U33 (.A( u0_u12_u7_n148 ) , .ZN( u0_u12_u7_n169 ) );
  INV_X1 u0_u12_u7_U34 (.A( u0_u12_u7_n127 ) , .ZN( u0_u12_u7_n179 ) );
  NOR2_X1 u0_u12_u7_U35 (.ZN( u0_u12_u7_n101 ) , .A2( u0_u12_u7_n150 ) , .A1( u0_u12_u7_n156 ) );
  AOI211_X1 u0_u12_u7_U36 (.B( u0_u12_u7_n154 ) , .A( u0_u12_u7_n155 ) , .C1( u0_u12_u7_n156 ) , .ZN( u0_u12_u7_n157 ) , .C2( u0_u12_u7_n172 ) );
  INV_X1 u0_u12_u7_U37 (.A( u0_u12_u7_n153 ) , .ZN( u0_u12_u7_n172 ) );
  AOI211_X1 u0_u12_u7_U38 (.B( u0_u12_u7_n139 ) , .A( u0_u12_u7_n140 ) , .C2( u0_u12_u7_n141 ) , .ZN( u0_u12_u7_n142 ) , .C1( u0_u12_u7_n156 ) );
  NAND4_X1 u0_u12_u7_U39 (.A3( u0_u12_u7_n127 ) , .A2( u0_u12_u7_n128 ) , .A1( u0_u12_u7_n129 ) , .ZN( u0_u12_u7_n141 ) , .A4( u0_u12_u7_n147 ) );
  INV_X1 u0_u12_u7_U4 (.A( u0_u12_u7_n111 ) , .ZN( u0_u12_u7_n170 ) );
  AOI21_X1 u0_u12_u7_U40 (.A( u0_u12_u7_n137 ) , .B1( u0_u12_u7_n138 ) , .ZN( u0_u12_u7_n139 ) , .B2( u0_u12_u7_n146 ) );
  OAI22_X1 u0_u12_u7_U41 (.B1( u0_u12_u7_n136 ) , .ZN( u0_u12_u7_n140 ) , .A1( u0_u12_u7_n153 ) , .B2( u0_u12_u7_n162 ) , .A2( u0_u12_u7_n164 ) );
  AOI21_X1 u0_u12_u7_U42 (.ZN( u0_u12_u7_n123 ) , .B1( u0_u12_u7_n165 ) , .B2( u0_u12_u7_n177 ) , .A( u0_u12_u7_n97 ) );
  AOI21_X1 u0_u12_u7_U43 (.B2( u0_u12_u7_n113 ) , .B1( u0_u12_u7_n124 ) , .A( u0_u12_u7_n125 ) , .ZN( u0_u12_u7_n97 ) );
  INV_X1 u0_u12_u7_U44 (.A( u0_u12_u7_n125 ) , .ZN( u0_u12_u7_n161 ) );
  INV_X1 u0_u12_u7_U45 (.A( u0_u12_u7_n152 ) , .ZN( u0_u12_u7_n162 ) );
  AOI22_X1 u0_u12_u7_U46 (.A2( u0_u12_u7_n114 ) , .ZN( u0_u12_u7_n119 ) , .B1( u0_u12_u7_n130 ) , .A1( u0_u12_u7_n156 ) , .B2( u0_u12_u7_n165 ) );
  NAND2_X1 u0_u12_u7_U47 (.A2( u0_u12_u7_n112 ) , .ZN( u0_u12_u7_n114 ) , .A1( u0_u12_u7_n175 ) );
  AND2_X1 u0_u12_u7_U48 (.ZN( u0_u12_u7_n145 ) , .A2( u0_u12_u7_n98 ) , .A1( u0_u12_u7_n99 ) );
  NOR2_X1 u0_u12_u7_U49 (.ZN( u0_u12_u7_n137 ) , .A1( u0_u12_u7_n150 ) , .A2( u0_u12_u7_n161 ) );
  INV_X1 u0_u12_u7_U5 (.A( u0_u12_u7_n149 ) , .ZN( u0_u12_u7_n175 ) );
  AOI21_X1 u0_u12_u7_U50 (.ZN( u0_u12_u7_n105 ) , .B2( u0_u12_u7_n110 ) , .A( u0_u12_u7_n125 ) , .B1( u0_u12_u7_n147 ) );
  NAND2_X1 u0_u12_u7_U51 (.ZN( u0_u12_u7_n146 ) , .A1( u0_u12_u7_n95 ) , .A2( u0_u12_u7_n98 ) );
  NAND2_X1 u0_u12_u7_U52 (.A2( u0_u12_u7_n103 ) , .ZN( u0_u12_u7_n147 ) , .A1( u0_u12_u7_n93 ) );
  NAND2_X1 u0_u12_u7_U53 (.A1( u0_u12_u7_n103 ) , .ZN( u0_u12_u7_n127 ) , .A2( u0_u12_u7_n99 ) );
  OR2_X1 u0_u12_u7_U54 (.ZN( u0_u12_u7_n126 ) , .A2( u0_u12_u7_n152 ) , .A1( u0_u12_u7_n156 ) );
  NAND2_X1 u0_u12_u7_U55 (.A2( u0_u12_u7_n102 ) , .A1( u0_u12_u7_n103 ) , .ZN( u0_u12_u7_n133 ) );
  NAND2_X1 u0_u12_u7_U56 (.ZN( u0_u12_u7_n112 ) , .A2( u0_u12_u7_n96 ) , .A1( u0_u12_u7_n99 ) );
  NAND2_X1 u0_u12_u7_U57 (.A2( u0_u12_u7_n102 ) , .ZN( u0_u12_u7_n128 ) , .A1( u0_u12_u7_n98 ) );
  NAND2_X1 u0_u12_u7_U58 (.A1( u0_u12_u7_n100 ) , .ZN( u0_u12_u7_n113 ) , .A2( u0_u12_u7_n93 ) );
  NAND2_X1 u0_u12_u7_U59 (.A2( u0_u12_u7_n102 ) , .ZN( u0_u12_u7_n124 ) , .A1( u0_u12_u7_n96 ) );
  INV_X1 u0_u12_u7_U6 (.A( u0_u12_u7_n154 ) , .ZN( u0_u12_u7_n178 ) );
  NAND2_X1 u0_u12_u7_U60 (.ZN( u0_u12_u7_n110 ) , .A1( u0_u12_u7_n95 ) , .A2( u0_u12_u7_n96 ) );
  INV_X1 u0_u12_u7_U61 (.A( u0_u12_u7_n150 ) , .ZN( u0_u12_u7_n164 ) );
  AND2_X1 u0_u12_u7_U62 (.ZN( u0_u12_u7_n134 ) , .A1( u0_u12_u7_n93 ) , .A2( u0_u12_u7_n98 ) );
  NAND2_X1 u0_u12_u7_U63 (.A1( u0_u12_u7_n100 ) , .A2( u0_u12_u7_n102 ) , .ZN( u0_u12_u7_n129 ) );
  NAND2_X1 u0_u12_u7_U64 (.A2( u0_u12_u7_n103 ) , .ZN( u0_u12_u7_n131 ) , .A1( u0_u12_u7_n95 ) );
  NAND2_X1 u0_u12_u7_U65 (.A1( u0_u12_u7_n100 ) , .ZN( u0_u12_u7_n138 ) , .A2( u0_u12_u7_n99 ) );
  NAND2_X1 u0_u12_u7_U66 (.ZN( u0_u12_u7_n132 ) , .A1( u0_u12_u7_n93 ) , .A2( u0_u12_u7_n96 ) );
  NAND2_X1 u0_u12_u7_U67 (.A1( u0_u12_u7_n100 ) , .ZN( u0_u12_u7_n148 ) , .A2( u0_u12_u7_n95 ) );
  NOR2_X1 u0_u12_u7_U68 (.A2( u0_u12_X_47 ) , .ZN( u0_u12_u7_n150 ) , .A1( u0_u12_u7_n163 ) );
  NOR2_X1 u0_u12_u7_U69 (.A2( u0_u12_X_43 ) , .A1( u0_u12_X_44 ) , .ZN( u0_u12_u7_n103 ) );
  AOI211_X1 u0_u12_u7_U7 (.ZN( u0_u12_u7_n116 ) , .A( u0_u12_u7_n155 ) , .C1( u0_u12_u7_n161 ) , .C2( u0_u12_u7_n171 ) , .B( u0_u12_u7_n94 ) );
  NOR2_X1 u0_u12_u7_U70 (.A2( u0_u12_X_48 ) , .A1( u0_u12_u7_n166 ) , .ZN( u0_u12_u7_n95 ) );
  NOR2_X1 u0_u12_u7_U71 (.A2( u0_u12_X_45 ) , .A1( u0_u12_X_48 ) , .ZN( u0_u12_u7_n99 ) );
  NOR2_X1 u0_u12_u7_U72 (.A2( u0_u12_X_44 ) , .A1( u0_u12_u7_n167 ) , .ZN( u0_u12_u7_n98 ) );
  NOR2_X1 u0_u12_u7_U73 (.A2( u0_u12_X_46 ) , .A1( u0_u12_X_47 ) , .ZN( u0_u12_u7_n152 ) );
  AND2_X1 u0_u12_u7_U74 (.A1( u0_u12_X_47 ) , .ZN( u0_u12_u7_n156 ) , .A2( u0_u12_u7_n163 ) );
  NAND2_X1 u0_u12_u7_U75 (.A2( u0_u12_X_46 ) , .A1( u0_u12_X_47 ) , .ZN( u0_u12_u7_n125 ) );
  AND2_X1 u0_u12_u7_U76 (.A2( u0_u12_X_45 ) , .A1( u0_u12_X_48 ) , .ZN( u0_u12_u7_n102 ) );
  AND2_X1 u0_u12_u7_U77 (.A2( u0_u12_X_43 ) , .A1( u0_u12_X_44 ) , .ZN( u0_u12_u7_n96 ) );
  AND2_X1 u0_u12_u7_U78 (.A1( u0_u12_X_44 ) , .ZN( u0_u12_u7_n100 ) , .A2( u0_u12_u7_n167 ) );
  AND2_X1 u0_u12_u7_U79 (.A1( u0_u12_X_48 ) , .A2( u0_u12_u7_n166 ) , .ZN( u0_u12_u7_n93 ) );
  OAI222_X1 u0_u12_u7_U8 (.C2( u0_u12_u7_n101 ) , .B2( u0_u12_u7_n111 ) , .A1( u0_u12_u7_n113 ) , .C1( u0_u12_u7_n146 ) , .A2( u0_u12_u7_n162 ) , .B1( u0_u12_u7_n164 ) , .ZN( u0_u12_u7_n94 ) );
  INV_X1 u0_u12_u7_U80 (.A( u0_u12_X_46 ) , .ZN( u0_u12_u7_n163 ) );
  INV_X1 u0_u12_u7_U81 (.A( u0_u12_X_43 ) , .ZN( u0_u12_u7_n167 ) );
  INV_X1 u0_u12_u7_U82 (.A( u0_u12_X_45 ) , .ZN( u0_u12_u7_n166 ) );
  NAND4_X1 u0_u12_u7_U83 (.ZN( u0_out12_27 ) , .A4( u0_u12_u7_n118 ) , .A3( u0_u12_u7_n119 ) , .A2( u0_u12_u7_n120 ) , .A1( u0_u12_u7_n121 ) );
  OAI21_X1 u0_u12_u7_U84 (.ZN( u0_u12_u7_n121 ) , .B2( u0_u12_u7_n145 ) , .A( u0_u12_u7_n150 ) , .B1( u0_u12_u7_n174 ) );
  OAI21_X1 u0_u12_u7_U85 (.ZN( u0_u12_u7_n120 ) , .A( u0_u12_u7_n161 ) , .B2( u0_u12_u7_n170 ) , .B1( u0_u12_u7_n179 ) );
  NAND4_X1 u0_u12_u7_U86 (.ZN( u0_out12_21 ) , .A4( u0_u12_u7_n157 ) , .A3( u0_u12_u7_n158 ) , .A2( u0_u12_u7_n159 ) , .A1( u0_u12_u7_n160 ) );
  OAI21_X1 u0_u12_u7_U87 (.B1( u0_u12_u7_n145 ) , .ZN( u0_u12_u7_n160 ) , .A( u0_u12_u7_n161 ) , .B2( u0_u12_u7_n177 ) );
  AOI22_X1 u0_u12_u7_U88 (.B2( u0_u12_u7_n149 ) , .B1( u0_u12_u7_n150 ) , .A2( u0_u12_u7_n151 ) , .A1( u0_u12_u7_n152 ) , .ZN( u0_u12_u7_n158 ) );
  NAND4_X1 u0_u12_u7_U89 (.ZN( u0_out12_15 ) , .A4( u0_u12_u7_n142 ) , .A3( u0_u12_u7_n143 ) , .A2( u0_u12_u7_n144 ) , .A1( u0_u12_u7_n178 ) );
  OAI221_X1 u0_u12_u7_U9 (.C1( u0_u12_u7_n101 ) , .C2( u0_u12_u7_n147 ) , .ZN( u0_u12_u7_n155 ) , .B2( u0_u12_u7_n162 ) , .A( u0_u12_u7_n91 ) , .B1( u0_u12_u7_n92 ) );
  OR2_X1 u0_u12_u7_U90 (.A2( u0_u12_u7_n125 ) , .A1( u0_u12_u7_n129 ) , .ZN( u0_u12_u7_n144 ) );
  AOI22_X1 u0_u12_u7_U91 (.A2( u0_u12_u7_n126 ) , .ZN( u0_u12_u7_n143 ) , .B2( u0_u12_u7_n165 ) , .B1( u0_u12_u7_n173 ) , .A1( u0_u12_u7_n174 ) );
  NAND4_X1 u0_u12_u7_U92 (.ZN( u0_out12_5 ) , .A4( u0_u12_u7_n108 ) , .A3( u0_u12_u7_n109 ) , .A1( u0_u12_u7_n116 ) , .A2( u0_u12_u7_n123 ) );
  AOI22_X1 u0_u12_u7_U93 (.ZN( u0_u12_u7_n109 ) , .A2( u0_u12_u7_n126 ) , .B2( u0_u12_u7_n145 ) , .B1( u0_u12_u7_n156 ) , .A1( u0_u12_u7_n171 ) );
  NOR4_X1 u0_u12_u7_U94 (.A4( u0_u12_u7_n104 ) , .A3( u0_u12_u7_n105 ) , .A2( u0_u12_u7_n106 ) , .A1( u0_u12_u7_n107 ) , .ZN( u0_u12_u7_n108 ) );
  NAND3_X1 u0_u12_u7_U95 (.A3( u0_u12_u7_n146 ) , .A2( u0_u12_u7_n147 ) , .A1( u0_u12_u7_n148 ) , .ZN( u0_u12_u7_n151 ) );
  NAND3_X1 u0_u12_u7_U96 (.A3( u0_u12_u7_n131 ) , .A2( u0_u12_u7_n132 ) , .A1( u0_u12_u7_n133 ) , .ZN( u0_u12_u7_n135 ) );
  XOR2_X1 u0_u13_U10 (.B( u0_K14_45 ) , .A( u0_R12_30 ) , .Z( u0_u13_X_45 ) );
  XOR2_X1 u0_u13_U11 (.B( u0_K14_44 ) , .A( u0_R12_29 ) , .Z( u0_u13_X_44 ) );
  XOR2_X1 u0_u13_U12 (.B( u0_K14_43 ) , .A( u0_R12_28 ) , .Z( u0_u13_X_43 ) );
  XOR2_X1 u0_u13_U13 (.B( u0_K14_42 ) , .A( u0_R12_29 ) , .Z( u0_u13_X_42 ) );
  XOR2_X1 u0_u13_U14 (.B( u0_K14_41 ) , .A( u0_R12_28 ) , .Z( u0_u13_X_41 ) );
  XOR2_X1 u0_u13_U17 (.B( u0_K14_39 ) , .A( u0_R12_26 ) , .Z( u0_u13_X_39 ) );
  XOR2_X1 u0_u13_U18 (.B( u0_K14_38 ) , .A( u0_R12_25 ) , .Z( u0_u13_X_38 ) );
  XOR2_X1 u0_u13_U19 (.B( u0_K14_37 ) , .A( u0_R12_24 ) , .Z( u0_u13_X_37 ) );
  XOR2_X1 u0_u13_U20 (.B( u0_K14_36 ) , .A( u0_R12_25 ) , .Z( u0_u13_X_36 ) );
  XOR2_X1 u0_u13_U21 (.B( u0_K14_35 ) , .A( u0_R12_24 ) , .Z( u0_u13_X_35 ) );
  XOR2_X1 u0_u13_U22 (.B( u0_K14_34 ) , .A( u0_R12_23 ) , .Z( u0_u13_X_34 ) );
  XOR2_X1 u0_u13_U23 (.B( u0_K14_33 ) , .A( u0_R12_22 ) , .Z( u0_u13_X_33 ) );
  XOR2_X1 u0_u13_U24 (.B( u0_K14_32 ) , .A( u0_R12_21 ) , .Z( u0_u13_X_32 ) );
  XOR2_X1 u0_u13_U25 (.B( u0_K14_31 ) , .A( u0_R12_20 ) , .Z( u0_u13_X_31 ) );
  XOR2_X1 u0_u13_U7 (.B( u0_K14_48 ) , .A( u0_R12_1 ) , .Z( u0_u13_X_48 ) );
  XOR2_X1 u0_u13_U8 (.B( u0_K14_47 ) , .A( u0_R12_32 ) , .Z( u0_u13_X_47 ) );
  INV_X1 u0_u13_u5_U10 (.A( u0_u13_u5_n121 ) , .ZN( u0_u13_u5_n177 ) );
  NOR3_X1 u0_u13_u5_U100 (.A3( u0_u13_u5_n141 ) , .A1( u0_u13_u5_n142 ) , .ZN( u0_u13_u5_n143 ) , .A2( u0_u13_u5_n191 ) );
  NAND4_X1 u0_u13_u5_U101 (.ZN( u0_out13_4 ) , .A4( u0_u13_u5_n112 ) , .A2( u0_u13_u5_n113 ) , .A1( u0_u13_u5_n114 ) , .A3( u0_u13_u5_n195 ) );
  AOI211_X1 u0_u13_u5_U102 (.A( u0_u13_u5_n110 ) , .C1( u0_u13_u5_n111 ) , .ZN( u0_u13_u5_n112 ) , .B( u0_u13_u5_n118 ) , .C2( u0_u13_u5_n177 ) );
  AOI222_X1 u0_u13_u5_U103 (.ZN( u0_u13_u5_n113 ) , .A1( u0_u13_u5_n131 ) , .C1( u0_u13_u5_n148 ) , .B2( u0_u13_u5_n174 ) , .C2( u0_u13_u5_n178 ) , .A2( u0_u13_u5_n179 ) , .B1( u0_u13_u5_n99 ) );
  NAND3_X1 u0_u13_u5_U104 (.A2( u0_u13_u5_n154 ) , .A3( u0_u13_u5_n158 ) , .A1( u0_u13_u5_n161 ) , .ZN( u0_u13_u5_n99 ) );
  NOR2_X1 u0_u13_u5_U11 (.ZN( u0_u13_u5_n160 ) , .A2( u0_u13_u5_n173 ) , .A1( u0_u13_u5_n177 ) );
  INV_X1 u0_u13_u5_U12 (.A( u0_u13_u5_n150 ) , .ZN( u0_u13_u5_n174 ) );
  AOI21_X1 u0_u13_u5_U13 (.A( u0_u13_u5_n160 ) , .B2( u0_u13_u5_n161 ) , .ZN( u0_u13_u5_n162 ) , .B1( u0_u13_u5_n192 ) );
  INV_X1 u0_u13_u5_U14 (.A( u0_u13_u5_n159 ) , .ZN( u0_u13_u5_n192 ) );
  AOI21_X1 u0_u13_u5_U15 (.A( u0_u13_u5_n156 ) , .B2( u0_u13_u5_n157 ) , .B1( u0_u13_u5_n158 ) , .ZN( u0_u13_u5_n163 ) );
  AOI21_X1 u0_u13_u5_U16 (.B2( u0_u13_u5_n139 ) , .B1( u0_u13_u5_n140 ) , .ZN( u0_u13_u5_n141 ) , .A( u0_u13_u5_n150 ) );
  OAI21_X1 u0_u13_u5_U17 (.A( u0_u13_u5_n133 ) , .B2( u0_u13_u5_n134 ) , .B1( u0_u13_u5_n135 ) , .ZN( u0_u13_u5_n142 ) );
  OAI21_X1 u0_u13_u5_U18 (.ZN( u0_u13_u5_n133 ) , .B2( u0_u13_u5_n147 ) , .A( u0_u13_u5_n173 ) , .B1( u0_u13_u5_n188 ) );
  NAND2_X1 u0_u13_u5_U19 (.A2( u0_u13_u5_n119 ) , .A1( u0_u13_u5_n123 ) , .ZN( u0_u13_u5_n137 ) );
  INV_X1 u0_u13_u5_U20 (.A( u0_u13_u5_n155 ) , .ZN( u0_u13_u5_n194 ) );
  NAND2_X1 u0_u13_u5_U21 (.A1( u0_u13_u5_n121 ) , .ZN( u0_u13_u5_n132 ) , .A2( u0_u13_u5_n172 ) );
  NAND2_X1 u0_u13_u5_U22 (.A2( u0_u13_u5_n122 ) , .ZN( u0_u13_u5_n136 ) , .A1( u0_u13_u5_n154 ) );
  NAND2_X1 u0_u13_u5_U23 (.A2( u0_u13_u5_n119 ) , .A1( u0_u13_u5_n120 ) , .ZN( u0_u13_u5_n159 ) );
  INV_X1 u0_u13_u5_U24 (.A( u0_u13_u5_n156 ) , .ZN( u0_u13_u5_n175 ) );
  INV_X1 u0_u13_u5_U25 (.A( u0_u13_u5_n158 ) , .ZN( u0_u13_u5_n188 ) );
  INV_X1 u0_u13_u5_U26 (.A( u0_u13_u5_n152 ) , .ZN( u0_u13_u5_n179 ) );
  INV_X1 u0_u13_u5_U27 (.A( u0_u13_u5_n140 ) , .ZN( u0_u13_u5_n182 ) );
  INV_X1 u0_u13_u5_U28 (.A( u0_u13_u5_n151 ) , .ZN( u0_u13_u5_n183 ) );
  INV_X1 u0_u13_u5_U29 (.A( u0_u13_u5_n123 ) , .ZN( u0_u13_u5_n185 ) );
  NOR2_X1 u0_u13_u5_U3 (.ZN( u0_u13_u5_n134 ) , .A1( u0_u13_u5_n183 ) , .A2( u0_u13_u5_n190 ) );
  INV_X1 u0_u13_u5_U30 (.A( u0_u13_u5_n161 ) , .ZN( u0_u13_u5_n184 ) );
  INV_X1 u0_u13_u5_U31 (.A( u0_u13_u5_n139 ) , .ZN( u0_u13_u5_n189 ) );
  INV_X1 u0_u13_u5_U32 (.A( u0_u13_u5_n157 ) , .ZN( u0_u13_u5_n190 ) );
  INV_X1 u0_u13_u5_U33 (.A( u0_u13_u5_n120 ) , .ZN( u0_u13_u5_n193 ) );
  NAND2_X1 u0_u13_u5_U34 (.ZN( u0_u13_u5_n111 ) , .A1( u0_u13_u5_n140 ) , .A2( u0_u13_u5_n155 ) );
  INV_X1 u0_u13_u5_U35 (.A( u0_u13_u5_n117 ) , .ZN( u0_u13_u5_n196 ) );
  OAI221_X1 u0_u13_u5_U36 (.A( u0_u13_u5_n116 ) , .ZN( u0_u13_u5_n117 ) , .B2( u0_u13_u5_n119 ) , .C1( u0_u13_u5_n153 ) , .C2( u0_u13_u5_n158 ) , .B1( u0_u13_u5_n172 ) );
  AOI222_X1 u0_u13_u5_U37 (.ZN( u0_u13_u5_n116 ) , .B2( u0_u13_u5_n145 ) , .C1( u0_u13_u5_n148 ) , .A2( u0_u13_u5_n174 ) , .C2( u0_u13_u5_n177 ) , .B1( u0_u13_u5_n187 ) , .A1( u0_u13_u5_n193 ) );
  INV_X1 u0_u13_u5_U38 (.A( u0_u13_u5_n115 ) , .ZN( u0_u13_u5_n187 ) );
  NOR2_X1 u0_u13_u5_U39 (.ZN( u0_u13_u5_n100 ) , .A1( u0_u13_u5_n170 ) , .A2( u0_u13_u5_n180 ) );
  INV_X1 u0_u13_u5_U4 (.A( u0_u13_u5_n138 ) , .ZN( u0_u13_u5_n191 ) );
  AOI22_X1 u0_u13_u5_U40 (.B2( u0_u13_u5_n131 ) , .A2( u0_u13_u5_n146 ) , .ZN( u0_u13_u5_n169 ) , .B1( u0_u13_u5_n174 ) , .A1( u0_u13_u5_n185 ) );
  NOR2_X1 u0_u13_u5_U41 (.A1( u0_u13_u5_n146 ) , .ZN( u0_u13_u5_n150 ) , .A2( u0_u13_u5_n173 ) );
  AOI21_X1 u0_u13_u5_U42 (.A( u0_u13_u5_n118 ) , .B2( u0_u13_u5_n145 ) , .ZN( u0_u13_u5_n168 ) , .B1( u0_u13_u5_n186 ) );
  INV_X1 u0_u13_u5_U43 (.A( u0_u13_u5_n122 ) , .ZN( u0_u13_u5_n186 ) );
  NOR2_X1 u0_u13_u5_U44 (.A1( u0_u13_u5_n146 ) , .ZN( u0_u13_u5_n152 ) , .A2( u0_u13_u5_n176 ) );
  NOR2_X1 u0_u13_u5_U45 (.A1( u0_u13_u5_n115 ) , .ZN( u0_u13_u5_n118 ) , .A2( u0_u13_u5_n153 ) );
  NOR2_X1 u0_u13_u5_U46 (.A2( u0_u13_u5_n145 ) , .ZN( u0_u13_u5_n156 ) , .A1( u0_u13_u5_n174 ) );
  NOR2_X1 u0_u13_u5_U47 (.ZN( u0_u13_u5_n121 ) , .A2( u0_u13_u5_n145 ) , .A1( u0_u13_u5_n176 ) );
  AOI22_X1 u0_u13_u5_U48 (.ZN( u0_u13_u5_n114 ) , .A2( u0_u13_u5_n137 ) , .A1( u0_u13_u5_n145 ) , .B2( u0_u13_u5_n175 ) , .B1( u0_u13_u5_n193 ) );
  OAI211_X1 u0_u13_u5_U49 (.B( u0_u13_u5_n124 ) , .A( u0_u13_u5_n125 ) , .C2( u0_u13_u5_n126 ) , .C1( u0_u13_u5_n127 ) , .ZN( u0_u13_u5_n128 ) );
  OAI21_X1 u0_u13_u5_U5 (.B2( u0_u13_u5_n136 ) , .B1( u0_u13_u5_n137 ) , .ZN( u0_u13_u5_n138 ) , .A( u0_u13_u5_n177 ) );
  NOR3_X1 u0_u13_u5_U50 (.ZN( u0_u13_u5_n127 ) , .A1( u0_u13_u5_n136 ) , .A3( u0_u13_u5_n148 ) , .A2( u0_u13_u5_n182 ) );
  OAI21_X1 u0_u13_u5_U51 (.ZN( u0_u13_u5_n124 ) , .A( u0_u13_u5_n177 ) , .B2( u0_u13_u5_n183 ) , .B1( u0_u13_u5_n189 ) );
  OAI21_X1 u0_u13_u5_U52 (.ZN( u0_u13_u5_n125 ) , .A( u0_u13_u5_n174 ) , .B2( u0_u13_u5_n185 ) , .B1( u0_u13_u5_n190 ) );
  AOI21_X1 u0_u13_u5_U53 (.A( u0_u13_u5_n153 ) , .B2( u0_u13_u5_n154 ) , .B1( u0_u13_u5_n155 ) , .ZN( u0_u13_u5_n164 ) );
  AOI21_X1 u0_u13_u5_U54 (.ZN( u0_u13_u5_n110 ) , .B1( u0_u13_u5_n122 ) , .B2( u0_u13_u5_n139 ) , .A( u0_u13_u5_n153 ) );
  INV_X1 u0_u13_u5_U55 (.A( u0_u13_u5_n153 ) , .ZN( u0_u13_u5_n176 ) );
  INV_X1 u0_u13_u5_U56 (.A( u0_u13_u5_n126 ) , .ZN( u0_u13_u5_n173 ) );
  AND2_X1 u0_u13_u5_U57 (.A2( u0_u13_u5_n104 ) , .A1( u0_u13_u5_n107 ) , .ZN( u0_u13_u5_n147 ) );
  AND2_X1 u0_u13_u5_U58 (.A2( u0_u13_u5_n104 ) , .A1( u0_u13_u5_n108 ) , .ZN( u0_u13_u5_n148 ) );
  NAND2_X1 u0_u13_u5_U59 (.A1( u0_u13_u5_n105 ) , .A2( u0_u13_u5_n106 ) , .ZN( u0_u13_u5_n158 ) );
  INV_X1 u0_u13_u5_U6 (.A( u0_u13_u5_n135 ) , .ZN( u0_u13_u5_n178 ) );
  NAND2_X1 u0_u13_u5_U60 (.A2( u0_u13_u5_n108 ) , .A1( u0_u13_u5_n109 ) , .ZN( u0_u13_u5_n139 ) );
  NAND2_X1 u0_u13_u5_U61 (.A1( u0_u13_u5_n106 ) , .A2( u0_u13_u5_n108 ) , .ZN( u0_u13_u5_n119 ) );
  NAND2_X1 u0_u13_u5_U62 (.A2( u0_u13_u5_n103 ) , .A1( u0_u13_u5_n105 ) , .ZN( u0_u13_u5_n140 ) );
  NAND2_X1 u0_u13_u5_U63 (.A2( u0_u13_u5_n104 ) , .A1( u0_u13_u5_n105 ) , .ZN( u0_u13_u5_n155 ) );
  NAND2_X1 u0_u13_u5_U64 (.A2( u0_u13_u5_n106 ) , .A1( u0_u13_u5_n107 ) , .ZN( u0_u13_u5_n122 ) );
  NAND2_X1 u0_u13_u5_U65 (.A2( u0_u13_u5_n100 ) , .A1( u0_u13_u5_n106 ) , .ZN( u0_u13_u5_n115 ) );
  NAND2_X1 u0_u13_u5_U66 (.A2( u0_u13_u5_n100 ) , .A1( u0_u13_u5_n103 ) , .ZN( u0_u13_u5_n161 ) );
  NAND2_X1 u0_u13_u5_U67 (.A1( u0_u13_u5_n105 ) , .A2( u0_u13_u5_n109 ) , .ZN( u0_u13_u5_n154 ) );
  INV_X1 u0_u13_u5_U68 (.A( u0_u13_u5_n146 ) , .ZN( u0_u13_u5_n172 ) );
  NAND2_X1 u0_u13_u5_U69 (.A1( u0_u13_u5_n103 ) , .A2( u0_u13_u5_n108 ) , .ZN( u0_u13_u5_n123 ) );
  OAI22_X1 u0_u13_u5_U7 (.B2( u0_u13_u5_n149 ) , .B1( u0_u13_u5_n150 ) , .A2( u0_u13_u5_n151 ) , .A1( u0_u13_u5_n152 ) , .ZN( u0_u13_u5_n165 ) );
  NAND2_X1 u0_u13_u5_U70 (.A2( u0_u13_u5_n103 ) , .A1( u0_u13_u5_n107 ) , .ZN( u0_u13_u5_n151 ) );
  NAND2_X1 u0_u13_u5_U71 (.A2( u0_u13_u5_n107 ) , .A1( u0_u13_u5_n109 ) , .ZN( u0_u13_u5_n120 ) );
  NAND2_X1 u0_u13_u5_U72 (.A2( u0_u13_u5_n100 ) , .A1( u0_u13_u5_n109 ) , .ZN( u0_u13_u5_n157 ) );
  AND2_X1 u0_u13_u5_U73 (.A2( u0_u13_u5_n100 ) , .A1( u0_u13_u5_n104 ) , .ZN( u0_u13_u5_n131 ) );
  INV_X1 u0_u13_u5_U74 (.A( u0_u13_u5_n102 ) , .ZN( u0_u13_u5_n195 ) );
  OAI221_X1 u0_u13_u5_U75 (.A( u0_u13_u5_n101 ) , .ZN( u0_u13_u5_n102 ) , .C2( u0_u13_u5_n115 ) , .C1( u0_u13_u5_n126 ) , .B1( u0_u13_u5_n134 ) , .B2( u0_u13_u5_n160 ) );
  OAI21_X1 u0_u13_u5_U76 (.ZN( u0_u13_u5_n101 ) , .B1( u0_u13_u5_n137 ) , .A( u0_u13_u5_n146 ) , .B2( u0_u13_u5_n147 ) );
  NOR2_X1 u0_u13_u5_U77 (.A2( u0_u13_X_34 ) , .A1( u0_u13_X_35 ) , .ZN( u0_u13_u5_n145 ) );
  NOR2_X1 u0_u13_u5_U78 (.A2( u0_u13_X_34 ) , .ZN( u0_u13_u5_n146 ) , .A1( u0_u13_u5_n171 ) );
  NOR2_X1 u0_u13_u5_U79 (.A2( u0_u13_X_31 ) , .A1( u0_u13_X_32 ) , .ZN( u0_u13_u5_n103 ) );
  NOR3_X1 u0_u13_u5_U8 (.A2( u0_u13_u5_n147 ) , .A1( u0_u13_u5_n148 ) , .ZN( u0_u13_u5_n149 ) , .A3( u0_u13_u5_n194 ) );
  NOR2_X1 u0_u13_u5_U80 (.A2( u0_u13_X_36 ) , .ZN( u0_u13_u5_n105 ) , .A1( u0_u13_u5_n180 ) );
  NOR2_X1 u0_u13_u5_U81 (.A2( u0_u13_X_33 ) , .ZN( u0_u13_u5_n108 ) , .A1( u0_u13_u5_n170 ) );
  NOR2_X1 u0_u13_u5_U82 (.A2( u0_u13_X_33 ) , .A1( u0_u13_X_36 ) , .ZN( u0_u13_u5_n107 ) );
  NOR2_X1 u0_u13_u5_U83 (.A2( u0_u13_X_31 ) , .ZN( u0_u13_u5_n104 ) , .A1( u0_u13_u5_n181 ) );
  NAND2_X1 u0_u13_u5_U84 (.A2( u0_u13_X_34 ) , .A1( u0_u13_X_35 ) , .ZN( u0_u13_u5_n153 ) );
  NAND2_X1 u0_u13_u5_U85 (.A1( u0_u13_X_34 ) , .ZN( u0_u13_u5_n126 ) , .A2( u0_u13_u5_n171 ) );
  AND2_X1 u0_u13_u5_U86 (.A1( u0_u13_X_31 ) , .A2( u0_u13_X_32 ) , .ZN( u0_u13_u5_n106 ) );
  AND2_X1 u0_u13_u5_U87 (.A1( u0_u13_X_31 ) , .ZN( u0_u13_u5_n109 ) , .A2( u0_u13_u5_n181 ) );
  INV_X1 u0_u13_u5_U88 (.A( u0_u13_X_33 ) , .ZN( u0_u13_u5_n180 ) );
  INV_X1 u0_u13_u5_U89 (.A( u0_u13_X_35 ) , .ZN( u0_u13_u5_n171 ) );
  NOR2_X1 u0_u13_u5_U9 (.ZN( u0_u13_u5_n135 ) , .A1( u0_u13_u5_n173 ) , .A2( u0_u13_u5_n176 ) );
  INV_X1 u0_u13_u5_U90 (.A( u0_u13_X_36 ) , .ZN( u0_u13_u5_n170 ) );
  INV_X1 u0_u13_u5_U91 (.A( u0_u13_X_32 ) , .ZN( u0_u13_u5_n181 ) );
  NAND4_X1 u0_u13_u5_U92 (.ZN( u0_out13_29 ) , .A4( u0_u13_u5_n129 ) , .A3( u0_u13_u5_n130 ) , .A2( u0_u13_u5_n168 ) , .A1( u0_u13_u5_n196 ) );
  AOI221_X1 u0_u13_u5_U93 (.A( u0_u13_u5_n128 ) , .ZN( u0_u13_u5_n129 ) , .C2( u0_u13_u5_n132 ) , .B2( u0_u13_u5_n159 ) , .B1( u0_u13_u5_n176 ) , .C1( u0_u13_u5_n184 ) );
  AOI222_X1 u0_u13_u5_U94 (.ZN( u0_u13_u5_n130 ) , .A2( u0_u13_u5_n146 ) , .B1( u0_u13_u5_n147 ) , .C2( u0_u13_u5_n175 ) , .B2( u0_u13_u5_n179 ) , .A1( u0_u13_u5_n188 ) , .C1( u0_u13_u5_n194 ) );
  NAND4_X1 u0_u13_u5_U95 (.ZN( u0_out13_19 ) , .A4( u0_u13_u5_n166 ) , .A3( u0_u13_u5_n167 ) , .A2( u0_u13_u5_n168 ) , .A1( u0_u13_u5_n169 ) );
  AOI22_X1 u0_u13_u5_U96 (.B2( u0_u13_u5_n145 ) , .A2( u0_u13_u5_n146 ) , .ZN( u0_u13_u5_n167 ) , .B1( u0_u13_u5_n182 ) , .A1( u0_u13_u5_n189 ) );
  NOR4_X1 u0_u13_u5_U97 (.A4( u0_u13_u5_n162 ) , .A3( u0_u13_u5_n163 ) , .A2( u0_u13_u5_n164 ) , .A1( u0_u13_u5_n165 ) , .ZN( u0_u13_u5_n166 ) );
  NAND4_X1 u0_u13_u5_U98 (.ZN( u0_out13_11 ) , .A4( u0_u13_u5_n143 ) , .A3( u0_u13_u5_n144 ) , .A2( u0_u13_u5_n169 ) , .A1( u0_u13_u5_n196 ) );
  AOI22_X1 u0_u13_u5_U99 (.A2( u0_u13_u5_n132 ) , .ZN( u0_u13_u5_n144 ) , .B2( u0_u13_u5_n145 ) , .B1( u0_u13_u5_n184 ) , .A1( u0_u13_u5_n194 ) );
  AOI22_X1 u0_u13_u6_U10 (.A2( u0_u13_u6_n151 ) , .B2( u0_u13_u6_n161 ) , .A1( u0_u13_u6_n167 ) , .B1( u0_u13_u6_n170 ) , .ZN( u0_u13_u6_n89 ) );
  AOI21_X1 u0_u13_u6_U11 (.B1( u0_u13_u6_n107 ) , .B2( u0_u13_u6_n132 ) , .A( u0_u13_u6_n158 ) , .ZN( u0_u13_u6_n88 ) );
  AOI21_X1 u0_u13_u6_U12 (.B2( u0_u13_u6_n147 ) , .B1( u0_u13_u6_n148 ) , .ZN( u0_u13_u6_n149 ) , .A( u0_u13_u6_n158 ) );
  AOI21_X1 u0_u13_u6_U13 (.ZN( u0_u13_u6_n106 ) , .A( u0_u13_u6_n142 ) , .B2( u0_u13_u6_n159 ) , .B1( u0_u13_u6_n164 ) );
  INV_X1 u0_u13_u6_U14 (.A( u0_u13_u6_n155 ) , .ZN( u0_u13_u6_n161 ) );
  INV_X1 u0_u13_u6_U15 (.A( u0_u13_u6_n128 ) , .ZN( u0_u13_u6_n164 ) );
  NAND2_X1 u0_u13_u6_U16 (.ZN( u0_u13_u6_n110 ) , .A1( u0_u13_u6_n122 ) , .A2( u0_u13_u6_n129 ) );
  NAND2_X1 u0_u13_u6_U17 (.ZN( u0_u13_u6_n124 ) , .A2( u0_u13_u6_n146 ) , .A1( u0_u13_u6_n148 ) );
  INV_X1 u0_u13_u6_U18 (.A( u0_u13_u6_n132 ) , .ZN( u0_u13_u6_n171 ) );
  AND2_X1 u0_u13_u6_U19 (.A1( u0_u13_u6_n100 ) , .ZN( u0_u13_u6_n130 ) , .A2( u0_u13_u6_n147 ) );
  INV_X1 u0_u13_u6_U20 (.A( u0_u13_u6_n127 ) , .ZN( u0_u13_u6_n173 ) );
  INV_X1 u0_u13_u6_U21 (.A( u0_u13_u6_n121 ) , .ZN( u0_u13_u6_n167 ) );
  INV_X1 u0_u13_u6_U22 (.A( u0_u13_u6_n100 ) , .ZN( u0_u13_u6_n169 ) );
  INV_X1 u0_u13_u6_U23 (.A( u0_u13_u6_n123 ) , .ZN( u0_u13_u6_n170 ) );
  INV_X1 u0_u13_u6_U24 (.A( u0_u13_u6_n113 ) , .ZN( u0_u13_u6_n168 ) );
  AND2_X1 u0_u13_u6_U25 (.A1( u0_u13_u6_n107 ) , .A2( u0_u13_u6_n119 ) , .ZN( u0_u13_u6_n133 ) );
  AND2_X1 u0_u13_u6_U26 (.A2( u0_u13_u6_n121 ) , .A1( u0_u13_u6_n122 ) , .ZN( u0_u13_u6_n131 ) );
  AND3_X1 u0_u13_u6_U27 (.ZN( u0_u13_u6_n120 ) , .A2( u0_u13_u6_n127 ) , .A1( u0_u13_u6_n132 ) , .A3( u0_u13_u6_n145 ) );
  INV_X1 u0_u13_u6_U28 (.A( u0_u13_u6_n146 ) , .ZN( u0_u13_u6_n163 ) );
  AOI222_X1 u0_u13_u6_U29 (.ZN( u0_u13_u6_n114 ) , .A1( u0_u13_u6_n118 ) , .A2( u0_u13_u6_n126 ) , .B2( u0_u13_u6_n151 ) , .C2( u0_u13_u6_n159 ) , .C1( u0_u13_u6_n168 ) , .B1( u0_u13_u6_n169 ) );
  INV_X1 u0_u13_u6_U3 (.A( u0_u13_u6_n110 ) , .ZN( u0_u13_u6_n166 ) );
  NOR2_X1 u0_u13_u6_U30 (.A1( u0_u13_u6_n162 ) , .A2( u0_u13_u6_n165 ) , .ZN( u0_u13_u6_n98 ) );
  AOI211_X1 u0_u13_u6_U31 (.B( u0_u13_u6_n134 ) , .A( u0_u13_u6_n135 ) , .C1( u0_u13_u6_n136 ) , .ZN( u0_u13_u6_n137 ) , .C2( u0_u13_u6_n151 ) );
  AOI21_X1 u0_u13_u6_U32 (.B2( u0_u13_u6_n132 ) , .B1( u0_u13_u6_n133 ) , .ZN( u0_u13_u6_n134 ) , .A( u0_u13_u6_n158 ) );
  AOI21_X1 u0_u13_u6_U33 (.B1( u0_u13_u6_n131 ) , .ZN( u0_u13_u6_n135 ) , .A( u0_u13_u6_n144 ) , .B2( u0_u13_u6_n146 ) );
  NAND4_X1 u0_u13_u6_U34 (.A4( u0_u13_u6_n127 ) , .A3( u0_u13_u6_n128 ) , .A2( u0_u13_u6_n129 ) , .A1( u0_u13_u6_n130 ) , .ZN( u0_u13_u6_n136 ) );
  NAND2_X1 u0_u13_u6_U35 (.A1( u0_u13_u6_n144 ) , .ZN( u0_u13_u6_n151 ) , .A2( u0_u13_u6_n158 ) );
  NAND2_X1 u0_u13_u6_U36 (.ZN( u0_u13_u6_n132 ) , .A1( u0_u13_u6_n91 ) , .A2( u0_u13_u6_n97 ) );
  AOI22_X1 u0_u13_u6_U37 (.B2( u0_u13_u6_n110 ) , .B1( u0_u13_u6_n111 ) , .A1( u0_u13_u6_n112 ) , .ZN( u0_u13_u6_n115 ) , .A2( u0_u13_u6_n161 ) );
  NAND4_X1 u0_u13_u6_U38 (.A3( u0_u13_u6_n109 ) , .ZN( u0_u13_u6_n112 ) , .A4( u0_u13_u6_n132 ) , .A2( u0_u13_u6_n147 ) , .A1( u0_u13_u6_n166 ) );
  NOR2_X1 u0_u13_u6_U39 (.ZN( u0_u13_u6_n109 ) , .A1( u0_u13_u6_n170 ) , .A2( u0_u13_u6_n173 ) );
  INV_X1 u0_u13_u6_U4 (.A( u0_u13_u6_n142 ) , .ZN( u0_u13_u6_n174 ) );
  NOR2_X1 u0_u13_u6_U40 (.A2( u0_u13_u6_n126 ) , .ZN( u0_u13_u6_n155 ) , .A1( u0_u13_u6_n160 ) );
  NAND2_X1 u0_u13_u6_U41 (.ZN( u0_u13_u6_n146 ) , .A2( u0_u13_u6_n94 ) , .A1( u0_u13_u6_n99 ) );
  AOI21_X1 u0_u13_u6_U42 (.A( u0_u13_u6_n144 ) , .B2( u0_u13_u6_n145 ) , .B1( u0_u13_u6_n146 ) , .ZN( u0_u13_u6_n150 ) );
  INV_X1 u0_u13_u6_U43 (.A( u0_u13_u6_n111 ) , .ZN( u0_u13_u6_n158 ) );
  NAND2_X1 u0_u13_u6_U44 (.ZN( u0_u13_u6_n127 ) , .A1( u0_u13_u6_n91 ) , .A2( u0_u13_u6_n92 ) );
  NAND2_X1 u0_u13_u6_U45 (.ZN( u0_u13_u6_n129 ) , .A2( u0_u13_u6_n95 ) , .A1( u0_u13_u6_n96 ) );
  INV_X1 u0_u13_u6_U46 (.A( u0_u13_u6_n144 ) , .ZN( u0_u13_u6_n159 ) );
  NAND2_X1 u0_u13_u6_U47 (.ZN( u0_u13_u6_n145 ) , .A2( u0_u13_u6_n97 ) , .A1( u0_u13_u6_n98 ) );
  NAND2_X1 u0_u13_u6_U48 (.ZN( u0_u13_u6_n148 ) , .A2( u0_u13_u6_n92 ) , .A1( u0_u13_u6_n94 ) );
  NAND2_X1 u0_u13_u6_U49 (.ZN( u0_u13_u6_n108 ) , .A2( u0_u13_u6_n139 ) , .A1( u0_u13_u6_n144 ) );
  NAND2_X1 u0_u13_u6_U5 (.A2( u0_u13_u6_n143 ) , .ZN( u0_u13_u6_n152 ) , .A1( u0_u13_u6_n166 ) );
  NAND2_X1 u0_u13_u6_U50 (.ZN( u0_u13_u6_n121 ) , .A2( u0_u13_u6_n95 ) , .A1( u0_u13_u6_n97 ) );
  NAND2_X1 u0_u13_u6_U51 (.ZN( u0_u13_u6_n107 ) , .A2( u0_u13_u6_n92 ) , .A1( u0_u13_u6_n95 ) );
  AND2_X1 u0_u13_u6_U52 (.ZN( u0_u13_u6_n118 ) , .A2( u0_u13_u6_n91 ) , .A1( u0_u13_u6_n99 ) );
  NAND2_X1 u0_u13_u6_U53 (.ZN( u0_u13_u6_n147 ) , .A2( u0_u13_u6_n98 ) , .A1( u0_u13_u6_n99 ) );
  NAND2_X1 u0_u13_u6_U54 (.ZN( u0_u13_u6_n128 ) , .A1( u0_u13_u6_n94 ) , .A2( u0_u13_u6_n96 ) );
  NAND2_X1 u0_u13_u6_U55 (.ZN( u0_u13_u6_n119 ) , .A2( u0_u13_u6_n95 ) , .A1( u0_u13_u6_n99 ) );
  NAND2_X1 u0_u13_u6_U56 (.ZN( u0_u13_u6_n123 ) , .A2( u0_u13_u6_n91 ) , .A1( u0_u13_u6_n96 ) );
  NAND2_X1 u0_u13_u6_U57 (.ZN( u0_u13_u6_n100 ) , .A2( u0_u13_u6_n92 ) , .A1( u0_u13_u6_n98 ) );
  NAND2_X1 u0_u13_u6_U58 (.ZN( u0_u13_u6_n122 ) , .A1( u0_u13_u6_n94 ) , .A2( u0_u13_u6_n97 ) );
  INV_X1 u0_u13_u6_U59 (.A( u0_u13_u6_n139 ) , .ZN( u0_u13_u6_n160 ) );
  AOI22_X1 u0_u13_u6_U6 (.B2( u0_u13_u6_n101 ) , .A1( u0_u13_u6_n102 ) , .ZN( u0_u13_u6_n103 ) , .B1( u0_u13_u6_n160 ) , .A2( u0_u13_u6_n161 ) );
  NAND2_X1 u0_u13_u6_U60 (.ZN( u0_u13_u6_n113 ) , .A1( u0_u13_u6_n96 ) , .A2( u0_u13_u6_n98 ) );
  NOR2_X1 u0_u13_u6_U61 (.A2( u0_u13_X_40 ) , .A1( u0_u13_X_41 ) , .ZN( u0_u13_u6_n126 ) );
  NOR2_X1 u0_u13_u6_U62 (.A2( u0_u13_X_39 ) , .A1( u0_u13_X_42 ) , .ZN( u0_u13_u6_n92 ) );
  NOR2_X1 u0_u13_u6_U63 (.A2( u0_u13_X_39 ) , .A1( u0_u13_u6_n156 ) , .ZN( u0_u13_u6_n97 ) );
  NOR2_X1 u0_u13_u6_U64 (.A2( u0_u13_X_38 ) , .A1( u0_u13_u6_n165 ) , .ZN( u0_u13_u6_n95 ) );
  NOR2_X1 u0_u13_u6_U65 (.A2( u0_u13_X_41 ) , .ZN( u0_u13_u6_n111 ) , .A1( u0_u13_u6_n157 ) );
  NOR2_X1 u0_u13_u6_U66 (.A2( u0_u13_X_37 ) , .A1( u0_u13_u6_n162 ) , .ZN( u0_u13_u6_n94 ) );
  NOR2_X1 u0_u13_u6_U67 (.A2( u0_u13_X_37 ) , .A1( u0_u13_X_38 ) , .ZN( u0_u13_u6_n91 ) );
  NAND2_X1 u0_u13_u6_U68 (.A1( u0_u13_X_41 ) , .ZN( u0_u13_u6_n144 ) , .A2( u0_u13_u6_n157 ) );
  NAND2_X1 u0_u13_u6_U69 (.A2( u0_u13_X_40 ) , .A1( u0_u13_X_41 ) , .ZN( u0_u13_u6_n139 ) );
  NOR2_X1 u0_u13_u6_U7 (.A1( u0_u13_u6_n118 ) , .ZN( u0_u13_u6_n143 ) , .A2( u0_u13_u6_n168 ) );
  AND2_X1 u0_u13_u6_U70 (.A1( u0_u13_X_39 ) , .A2( u0_u13_u6_n156 ) , .ZN( u0_u13_u6_n96 ) );
  AND2_X1 u0_u13_u6_U71 (.A1( u0_u13_X_39 ) , .A2( u0_u13_X_42 ) , .ZN( u0_u13_u6_n99 ) );
  INV_X1 u0_u13_u6_U72 (.A( u0_u13_X_40 ) , .ZN( u0_u13_u6_n157 ) );
  INV_X1 u0_u13_u6_U73 (.A( u0_u13_X_37 ) , .ZN( u0_u13_u6_n165 ) );
  INV_X1 u0_u13_u6_U74 (.A( u0_u13_X_38 ) , .ZN( u0_u13_u6_n162 ) );
  INV_X1 u0_u13_u6_U75 (.A( u0_u13_X_42 ) , .ZN( u0_u13_u6_n156 ) );
  NAND4_X1 u0_u13_u6_U76 (.ZN( u0_out13_32 ) , .A4( u0_u13_u6_n103 ) , .A3( u0_u13_u6_n104 ) , .A2( u0_u13_u6_n105 ) , .A1( u0_u13_u6_n106 ) );
  AOI22_X1 u0_u13_u6_U77 (.ZN( u0_u13_u6_n105 ) , .A2( u0_u13_u6_n108 ) , .A1( u0_u13_u6_n118 ) , .B2( u0_u13_u6_n126 ) , .B1( u0_u13_u6_n171 ) );
  AOI22_X1 u0_u13_u6_U78 (.ZN( u0_u13_u6_n104 ) , .A1( u0_u13_u6_n111 ) , .B1( u0_u13_u6_n124 ) , .B2( u0_u13_u6_n151 ) , .A2( u0_u13_u6_n93 ) );
  NAND4_X1 u0_u13_u6_U79 (.ZN( u0_out13_12 ) , .A4( u0_u13_u6_n114 ) , .A3( u0_u13_u6_n115 ) , .A2( u0_u13_u6_n116 ) , .A1( u0_u13_u6_n117 ) );
  OAI21_X1 u0_u13_u6_U8 (.A( u0_u13_u6_n159 ) , .B1( u0_u13_u6_n169 ) , .B2( u0_u13_u6_n173 ) , .ZN( u0_u13_u6_n90 ) );
  OAI22_X1 u0_u13_u6_U80 (.B2( u0_u13_u6_n111 ) , .ZN( u0_u13_u6_n116 ) , .B1( u0_u13_u6_n126 ) , .A2( u0_u13_u6_n164 ) , .A1( u0_u13_u6_n167 ) );
  OAI21_X1 u0_u13_u6_U81 (.A( u0_u13_u6_n108 ) , .ZN( u0_u13_u6_n117 ) , .B2( u0_u13_u6_n141 ) , .B1( u0_u13_u6_n163 ) );
  OAI211_X1 u0_u13_u6_U82 (.ZN( u0_out13_7 ) , .B( u0_u13_u6_n153 ) , .C2( u0_u13_u6_n154 ) , .C1( u0_u13_u6_n155 ) , .A( u0_u13_u6_n174 ) );
  NOR3_X1 u0_u13_u6_U83 (.A1( u0_u13_u6_n141 ) , .ZN( u0_u13_u6_n154 ) , .A3( u0_u13_u6_n164 ) , .A2( u0_u13_u6_n171 ) );
  AOI211_X1 u0_u13_u6_U84 (.B( u0_u13_u6_n149 ) , .A( u0_u13_u6_n150 ) , .C2( u0_u13_u6_n151 ) , .C1( u0_u13_u6_n152 ) , .ZN( u0_u13_u6_n153 ) );
  OAI211_X1 u0_u13_u6_U85 (.ZN( u0_out13_22 ) , .B( u0_u13_u6_n137 ) , .A( u0_u13_u6_n138 ) , .C2( u0_u13_u6_n139 ) , .C1( u0_u13_u6_n140 ) );
  AOI22_X1 u0_u13_u6_U86 (.B1( u0_u13_u6_n124 ) , .A2( u0_u13_u6_n125 ) , .A1( u0_u13_u6_n126 ) , .ZN( u0_u13_u6_n138 ) , .B2( u0_u13_u6_n161 ) );
  AND4_X1 u0_u13_u6_U87 (.A3( u0_u13_u6_n119 ) , .A1( u0_u13_u6_n120 ) , .A4( u0_u13_u6_n129 ) , .ZN( u0_u13_u6_n140 ) , .A2( u0_u13_u6_n143 ) );
  NAND3_X1 u0_u13_u6_U88 (.A2( u0_u13_u6_n123 ) , .ZN( u0_u13_u6_n125 ) , .A1( u0_u13_u6_n130 ) , .A3( u0_u13_u6_n131 ) );
  NAND3_X1 u0_u13_u6_U89 (.A3( u0_u13_u6_n133 ) , .ZN( u0_u13_u6_n141 ) , .A1( u0_u13_u6_n145 ) , .A2( u0_u13_u6_n148 ) );
  INV_X1 u0_u13_u6_U9 (.ZN( u0_u13_u6_n172 ) , .A( u0_u13_u6_n88 ) );
  NAND3_X1 u0_u13_u6_U90 (.ZN( u0_u13_u6_n101 ) , .A3( u0_u13_u6_n107 ) , .A2( u0_u13_u6_n121 ) , .A1( u0_u13_u6_n127 ) );
  NAND3_X1 u0_u13_u6_U91 (.ZN( u0_u13_u6_n102 ) , .A3( u0_u13_u6_n130 ) , .A2( u0_u13_u6_n145 ) , .A1( u0_u13_u6_n166 ) );
  NAND3_X1 u0_u13_u6_U92 (.A3( u0_u13_u6_n113 ) , .A1( u0_u13_u6_n119 ) , .A2( u0_u13_u6_n123 ) , .ZN( u0_u13_u6_n93 ) );
  NAND3_X1 u0_u13_u6_U93 (.ZN( u0_u13_u6_n142 ) , .A2( u0_u13_u6_n172 ) , .A3( u0_u13_u6_n89 ) , .A1( u0_u13_u6_n90 ) );
  AND3_X1 u0_u13_u7_U10 (.A3( u0_u13_u7_n110 ) , .A2( u0_u13_u7_n127 ) , .A1( u0_u13_u7_n132 ) , .ZN( u0_u13_u7_n92 ) );
  OAI21_X1 u0_u13_u7_U11 (.A( u0_u13_u7_n161 ) , .B1( u0_u13_u7_n168 ) , .B2( u0_u13_u7_n173 ) , .ZN( u0_u13_u7_n91 ) );
  AOI211_X1 u0_u13_u7_U12 (.A( u0_u13_u7_n117 ) , .ZN( u0_u13_u7_n118 ) , .C2( u0_u13_u7_n126 ) , .C1( u0_u13_u7_n177 ) , .B( u0_u13_u7_n180 ) );
  OAI22_X1 u0_u13_u7_U13 (.B1( u0_u13_u7_n115 ) , .ZN( u0_u13_u7_n117 ) , .A2( u0_u13_u7_n133 ) , .A1( u0_u13_u7_n137 ) , .B2( u0_u13_u7_n162 ) );
  INV_X1 u0_u13_u7_U14 (.A( u0_u13_u7_n116 ) , .ZN( u0_u13_u7_n180 ) );
  NOR3_X1 u0_u13_u7_U15 (.ZN( u0_u13_u7_n115 ) , .A3( u0_u13_u7_n145 ) , .A2( u0_u13_u7_n168 ) , .A1( u0_u13_u7_n169 ) );
  OAI211_X1 u0_u13_u7_U16 (.B( u0_u13_u7_n122 ) , .A( u0_u13_u7_n123 ) , .C2( u0_u13_u7_n124 ) , .ZN( u0_u13_u7_n154 ) , .C1( u0_u13_u7_n162 ) );
  AOI222_X1 u0_u13_u7_U17 (.ZN( u0_u13_u7_n122 ) , .C2( u0_u13_u7_n126 ) , .C1( u0_u13_u7_n145 ) , .B1( u0_u13_u7_n161 ) , .A2( u0_u13_u7_n165 ) , .B2( u0_u13_u7_n170 ) , .A1( u0_u13_u7_n176 ) );
  INV_X1 u0_u13_u7_U18 (.A( u0_u13_u7_n133 ) , .ZN( u0_u13_u7_n176 ) );
  NOR3_X1 u0_u13_u7_U19 (.A2( u0_u13_u7_n134 ) , .A1( u0_u13_u7_n135 ) , .ZN( u0_u13_u7_n136 ) , .A3( u0_u13_u7_n171 ) );
  NOR2_X1 u0_u13_u7_U20 (.A1( u0_u13_u7_n130 ) , .A2( u0_u13_u7_n134 ) , .ZN( u0_u13_u7_n153 ) );
  INV_X1 u0_u13_u7_U21 (.A( u0_u13_u7_n101 ) , .ZN( u0_u13_u7_n165 ) );
  NOR2_X1 u0_u13_u7_U22 (.ZN( u0_u13_u7_n111 ) , .A2( u0_u13_u7_n134 ) , .A1( u0_u13_u7_n169 ) );
  AOI21_X1 u0_u13_u7_U23 (.ZN( u0_u13_u7_n104 ) , .B2( u0_u13_u7_n112 ) , .B1( u0_u13_u7_n127 ) , .A( u0_u13_u7_n164 ) );
  AOI21_X1 u0_u13_u7_U24 (.ZN( u0_u13_u7_n106 ) , .B1( u0_u13_u7_n133 ) , .B2( u0_u13_u7_n146 ) , .A( u0_u13_u7_n162 ) );
  AOI21_X1 u0_u13_u7_U25 (.A( u0_u13_u7_n101 ) , .ZN( u0_u13_u7_n107 ) , .B2( u0_u13_u7_n128 ) , .B1( u0_u13_u7_n175 ) );
  INV_X1 u0_u13_u7_U26 (.A( u0_u13_u7_n138 ) , .ZN( u0_u13_u7_n171 ) );
  INV_X1 u0_u13_u7_U27 (.A( u0_u13_u7_n131 ) , .ZN( u0_u13_u7_n177 ) );
  INV_X1 u0_u13_u7_U28 (.A( u0_u13_u7_n110 ) , .ZN( u0_u13_u7_n174 ) );
  NAND2_X1 u0_u13_u7_U29 (.A1( u0_u13_u7_n129 ) , .A2( u0_u13_u7_n132 ) , .ZN( u0_u13_u7_n149 ) );
  OAI21_X1 u0_u13_u7_U3 (.ZN( u0_u13_u7_n159 ) , .A( u0_u13_u7_n165 ) , .B2( u0_u13_u7_n171 ) , .B1( u0_u13_u7_n174 ) );
  NAND2_X1 u0_u13_u7_U30 (.A1( u0_u13_u7_n113 ) , .A2( u0_u13_u7_n124 ) , .ZN( u0_u13_u7_n130 ) );
  INV_X1 u0_u13_u7_U31 (.A( u0_u13_u7_n112 ) , .ZN( u0_u13_u7_n173 ) );
  INV_X1 u0_u13_u7_U32 (.A( u0_u13_u7_n128 ) , .ZN( u0_u13_u7_n168 ) );
  INV_X1 u0_u13_u7_U33 (.A( u0_u13_u7_n148 ) , .ZN( u0_u13_u7_n169 ) );
  INV_X1 u0_u13_u7_U34 (.A( u0_u13_u7_n127 ) , .ZN( u0_u13_u7_n179 ) );
  NOR2_X1 u0_u13_u7_U35 (.ZN( u0_u13_u7_n101 ) , .A2( u0_u13_u7_n150 ) , .A1( u0_u13_u7_n156 ) );
  AOI211_X1 u0_u13_u7_U36 (.B( u0_u13_u7_n154 ) , .A( u0_u13_u7_n155 ) , .C1( u0_u13_u7_n156 ) , .ZN( u0_u13_u7_n157 ) , .C2( u0_u13_u7_n172 ) );
  INV_X1 u0_u13_u7_U37 (.A( u0_u13_u7_n153 ) , .ZN( u0_u13_u7_n172 ) );
  AOI211_X1 u0_u13_u7_U38 (.B( u0_u13_u7_n139 ) , .A( u0_u13_u7_n140 ) , .C2( u0_u13_u7_n141 ) , .ZN( u0_u13_u7_n142 ) , .C1( u0_u13_u7_n156 ) );
  NAND4_X1 u0_u13_u7_U39 (.A3( u0_u13_u7_n127 ) , .A2( u0_u13_u7_n128 ) , .A1( u0_u13_u7_n129 ) , .ZN( u0_u13_u7_n141 ) , .A4( u0_u13_u7_n147 ) );
  INV_X1 u0_u13_u7_U4 (.A( u0_u13_u7_n111 ) , .ZN( u0_u13_u7_n170 ) );
  AOI21_X1 u0_u13_u7_U40 (.A( u0_u13_u7_n137 ) , .B1( u0_u13_u7_n138 ) , .ZN( u0_u13_u7_n139 ) , .B2( u0_u13_u7_n146 ) );
  OAI22_X1 u0_u13_u7_U41 (.B1( u0_u13_u7_n136 ) , .ZN( u0_u13_u7_n140 ) , .A1( u0_u13_u7_n153 ) , .B2( u0_u13_u7_n162 ) , .A2( u0_u13_u7_n164 ) );
  AOI21_X1 u0_u13_u7_U42 (.ZN( u0_u13_u7_n123 ) , .B1( u0_u13_u7_n165 ) , .B2( u0_u13_u7_n177 ) , .A( u0_u13_u7_n97 ) );
  AOI21_X1 u0_u13_u7_U43 (.B2( u0_u13_u7_n113 ) , .B1( u0_u13_u7_n124 ) , .A( u0_u13_u7_n125 ) , .ZN( u0_u13_u7_n97 ) );
  INV_X1 u0_u13_u7_U44 (.A( u0_u13_u7_n125 ) , .ZN( u0_u13_u7_n161 ) );
  INV_X1 u0_u13_u7_U45 (.A( u0_u13_u7_n152 ) , .ZN( u0_u13_u7_n162 ) );
  AOI22_X1 u0_u13_u7_U46 (.A2( u0_u13_u7_n114 ) , .ZN( u0_u13_u7_n119 ) , .B1( u0_u13_u7_n130 ) , .A1( u0_u13_u7_n156 ) , .B2( u0_u13_u7_n165 ) );
  NAND2_X1 u0_u13_u7_U47 (.A2( u0_u13_u7_n112 ) , .ZN( u0_u13_u7_n114 ) , .A1( u0_u13_u7_n175 ) );
  AND2_X1 u0_u13_u7_U48 (.ZN( u0_u13_u7_n145 ) , .A2( u0_u13_u7_n98 ) , .A1( u0_u13_u7_n99 ) );
  NOR2_X1 u0_u13_u7_U49 (.ZN( u0_u13_u7_n137 ) , .A1( u0_u13_u7_n150 ) , .A2( u0_u13_u7_n161 ) );
  INV_X1 u0_u13_u7_U5 (.A( u0_u13_u7_n149 ) , .ZN( u0_u13_u7_n175 ) );
  AOI21_X1 u0_u13_u7_U50 (.ZN( u0_u13_u7_n105 ) , .B2( u0_u13_u7_n110 ) , .A( u0_u13_u7_n125 ) , .B1( u0_u13_u7_n147 ) );
  NAND2_X1 u0_u13_u7_U51 (.ZN( u0_u13_u7_n146 ) , .A1( u0_u13_u7_n95 ) , .A2( u0_u13_u7_n98 ) );
  NAND2_X1 u0_u13_u7_U52 (.A2( u0_u13_u7_n103 ) , .ZN( u0_u13_u7_n147 ) , .A1( u0_u13_u7_n93 ) );
  NAND2_X1 u0_u13_u7_U53 (.A1( u0_u13_u7_n103 ) , .ZN( u0_u13_u7_n127 ) , .A2( u0_u13_u7_n99 ) );
  OR2_X1 u0_u13_u7_U54 (.ZN( u0_u13_u7_n126 ) , .A2( u0_u13_u7_n152 ) , .A1( u0_u13_u7_n156 ) );
  NAND2_X1 u0_u13_u7_U55 (.A2( u0_u13_u7_n102 ) , .A1( u0_u13_u7_n103 ) , .ZN( u0_u13_u7_n133 ) );
  NAND2_X1 u0_u13_u7_U56 (.ZN( u0_u13_u7_n112 ) , .A2( u0_u13_u7_n96 ) , .A1( u0_u13_u7_n99 ) );
  NAND2_X1 u0_u13_u7_U57 (.A2( u0_u13_u7_n102 ) , .ZN( u0_u13_u7_n128 ) , .A1( u0_u13_u7_n98 ) );
  NAND2_X1 u0_u13_u7_U58 (.A1( u0_u13_u7_n100 ) , .ZN( u0_u13_u7_n113 ) , .A2( u0_u13_u7_n93 ) );
  NAND2_X1 u0_u13_u7_U59 (.A2( u0_u13_u7_n102 ) , .ZN( u0_u13_u7_n124 ) , .A1( u0_u13_u7_n96 ) );
  INV_X1 u0_u13_u7_U6 (.A( u0_u13_u7_n154 ) , .ZN( u0_u13_u7_n178 ) );
  NAND2_X1 u0_u13_u7_U60 (.ZN( u0_u13_u7_n110 ) , .A1( u0_u13_u7_n95 ) , .A2( u0_u13_u7_n96 ) );
  INV_X1 u0_u13_u7_U61 (.A( u0_u13_u7_n150 ) , .ZN( u0_u13_u7_n164 ) );
  AND2_X1 u0_u13_u7_U62 (.ZN( u0_u13_u7_n134 ) , .A1( u0_u13_u7_n93 ) , .A2( u0_u13_u7_n98 ) );
  NAND2_X1 u0_u13_u7_U63 (.A1( u0_u13_u7_n100 ) , .A2( u0_u13_u7_n102 ) , .ZN( u0_u13_u7_n129 ) );
  NAND2_X1 u0_u13_u7_U64 (.A2( u0_u13_u7_n103 ) , .ZN( u0_u13_u7_n131 ) , .A1( u0_u13_u7_n95 ) );
  NAND2_X1 u0_u13_u7_U65 (.A1( u0_u13_u7_n100 ) , .ZN( u0_u13_u7_n138 ) , .A2( u0_u13_u7_n99 ) );
  NAND2_X1 u0_u13_u7_U66 (.ZN( u0_u13_u7_n132 ) , .A1( u0_u13_u7_n93 ) , .A2( u0_u13_u7_n96 ) );
  NAND2_X1 u0_u13_u7_U67 (.A1( u0_u13_u7_n100 ) , .ZN( u0_u13_u7_n148 ) , .A2( u0_u13_u7_n95 ) );
  NOR2_X1 u0_u13_u7_U68 (.A2( u0_u13_X_47 ) , .ZN( u0_u13_u7_n150 ) , .A1( u0_u13_u7_n163 ) );
  NOR2_X1 u0_u13_u7_U69 (.A2( u0_u13_X_43 ) , .A1( u0_u13_X_44 ) , .ZN( u0_u13_u7_n103 ) );
  AOI211_X1 u0_u13_u7_U7 (.ZN( u0_u13_u7_n116 ) , .A( u0_u13_u7_n155 ) , .C1( u0_u13_u7_n161 ) , .C2( u0_u13_u7_n171 ) , .B( u0_u13_u7_n94 ) );
  NOR2_X1 u0_u13_u7_U70 (.A2( u0_u13_X_48 ) , .A1( u0_u13_u7_n166 ) , .ZN( u0_u13_u7_n95 ) );
  NOR2_X1 u0_u13_u7_U71 (.A2( u0_u13_X_45 ) , .A1( u0_u13_X_48 ) , .ZN( u0_u13_u7_n99 ) );
  NOR2_X1 u0_u13_u7_U72 (.A2( u0_u13_X_44 ) , .A1( u0_u13_u7_n167 ) , .ZN( u0_u13_u7_n98 ) );
  NOR2_X1 u0_u13_u7_U73 (.A2( u0_u13_X_46 ) , .A1( u0_u13_X_47 ) , .ZN( u0_u13_u7_n152 ) );
  AND2_X1 u0_u13_u7_U74 (.A1( u0_u13_X_47 ) , .ZN( u0_u13_u7_n156 ) , .A2( u0_u13_u7_n163 ) );
  NAND2_X1 u0_u13_u7_U75 (.A2( u0_u13_X_46 ) , .A1( u0_u13_X_47 ) , .ZN( u0_u13_u7_n125 ) );
  AND2_X1 u0_u13_u7_U76 (.A2( u0_u13_X_45 ) , .A1( u0_u13_X_48 ) , .ZN( u0_u13_u7_n102 ) );
  AND2_X1 u0_u13_u7_U77 (.A2( u0_u13_X_43 ) , .A1( u0_u13_X_44 ) , .ZN( u0_u13_u7_n96 ) );
  AND2_X1 u0_u13_u7_U78 (.A1( u0_u13_X_44 ) , .ZN( u0_u13_u7_n100 ) , .A2( u0_u13_u7_n167 ) );
  AND2_X1 u0_u13_u7_U79 (.A1( u0_u13_X_48 ) , .A2( u0_u13_u7_n166 ) , .ZN( u0_u13_u7_n93 ) );
  OAI222_X1 u0_u13_u7_U8 (.C2( u0_u13_u7_n101 ) , .B2( u0_u13_u7_n111 ) , .A1( u0_u13_u7_n113 ) , .C1( u0_u13_u7_n146 ) , .A2( u0_u13_u7_n162 ) , .B1( u0_u13_u7_n164 ) , .ZN( u0_u13_u7_n94 ) );
  INV_X1 u0_u13_u7_U80 (.A( u0_u13_X_46 ) , .ZN( u0_u13_u7_n163 ) );
  INV_X1 u0_u13_u7_U81 (.A( u0_u13_X_43 ) , .ZN( u0_u13_u7_n167 ) );
  INV_X1 u0_u13_u7_U82 (.A( u0_u13_X_45 ) , .ZN( u0_u13_u7_n166 ) );
  NAND4_X1 u0_u13_u7_U83 (.ZN( u0_out13_27 ) , .A4( u0_u13_u7_n118 ) , .A3( u0_u13_u7_n119 ) , .A2( u0_u13_u7_n120 ) , .A1( u0_u13_u7_n121 ) );
  OAI21_X1 u0_u13_u7_U84 (.ZN( u0_u13_u7_n121 ) , .B2( u0_u13_u7_n145 ) , .A( u0_u13_u7_n150 ) , .B1( u0_u13_u7_n174 ) );
  OAI21_X1 u0_u13_u7_U85 (.ZN( u0_u13_u7_n120 ) , .A( u0_u13_u7_n161 ) , .B2( u0_u13_u7_n170 ) , .B1( u0_u13_u7_n179 ) );
  NAND4_X1 u0_u13_u7_U86 (.ZN( u0_out13_21 ) , .A4( u0_u13_u7_n157 ) , .A3( u0_u13_u7_n158 ) , .A2( u0_u13_u7_n159 ) , .A1( u0_u13_u7_n160 ) );
  OAI21_X1 u0_u13_u7_U87 (.B1( u0_u13_u7_n145 ) , .ZN( u0_u13_u7_n160 ) , .A( u0_u13_u7_n161 ) , .B2( u0_u13_u7_n177 ) );
  AOI22_X1 u0_u13_u7_U88 (.B2( u0_u13_u7_n149 ) , .B1( u0_u13_u7_n150 ) , .A2( u0_u13_u7_n151 ) , .A1( u0_u13_u7_n152 ) , .ZN( u0_u13_u7_n158 ) );
  NAND4_X1 u0_u13_u7_U89 (.ZN( u0_out13_15 ) , .A4( u0_u13_u7_n142 ) , .A3( u0_u13_u7_n143 ) , .A2( u0_u13_u7_n144 ) , .A1( u0_u13_u7_n178 ) );
  OAI221_X1 u0_u13_u7_U9 (.C1( u0_u13_u7_n101 ) , .C2( u0_u13_u7_n147 ) , .ZN( u0_u13_u7_n155 ) , .B2( u0_u13_u7_n162 ) , .A( u0_u13_u7_n91 ) , .B1( u0_u13_u7_n92 ) );
  OR2_X1 u0_u13_u7_U90 (.A2( u0_u13_u7_n125 ) , .A1( u0_u13_u7_n129 ) , .ZN( u0_u13_u7_n144 ) );
  AOI22_X1 u0_u13_u7_U91 (.A2( u0_u13_u7_n126 ) , .ZN( u0_u13_u7_n143 ) , .B2( u0_u13_u7_n165 ) , .B1( u0_u13_u7_n173 ) , .A1( u0_u13_u7_n174 ) );
  NAND4_X1 u0_u13_u7_U92 (.ZN( u0_out13_5 ) , .A4( u0_u13_u7_n108 ) , .A3( u0_u13_u7_n109 ) , .A1( u0_u13_u7_n116 ) , .A2( u0_u13_u7_n123 ) );
  AOI22_X1 u0_u13_u7_U93 (.ZN( u0_u13_u7_n109 ) , .A2( u0_u13_u7_n126 ) , .B2( u0_u13_u7_n145 ) , .B1( u0_u13_u7_n156 ) , .A1( u0_u13_u7_n171 ) );
  NOR4_X1 u0_u13_u7_U94 (.A4( u0_u13_u7_n104 ) , .A3( u0_u13_u7_n105 ) , .A2( u0_u13_u7_n106 ) , .A1( u0_u13_u7_n107 ) , .ZN( u0_u13_u7_n108 ) );
  NAND3_X1 u0_u13_u7_U95 (.A3( u0_u13_u7_n146 ) , .A2( u0_u13_u7_n147 ) , .A1( u0_u13_u7_n148 ) , .ZN( u0_u13_u7_n151 ) );
  NAND3_X1 u0_u13_u7_U96 (.A3( u0_u13_u7_n131 ) , .A2( u0_u13_u7_n132 ) , .A1( u0_u13_u7_n133 ) , .ZN( u0_u13_u7_n135 ) );
  XOR2_X1 u0_u15_U1 (.A( u0_FP_38 ) , .B( u0_K16_9 ) , .Z( u0_u15_X_9 ) );
  XOR2_X1 u0_u15_U16 (.A( u0_FP_34 ) , .B( u0_K16_3 ) , .Z( u0_u15_X_3 ) );
  XOR2_X1 u0_u15_U2 (.A( u0_FP_37 ) , .B( u0_K16_8 ) , .Z( u0_u15_X_8 ) );
  XOR2_X1 u0_u15_U27 (.A( u0_FP_33 ) , .B( u0_K16_2 ) , .Z( u0_u15_X_2 ) );
  XOR2_X1 u0_u15_U3 (.A( u0_FP_36 ) , .B( u0_K16_7 ) , .Z( u0_u15_X_7 ) );
  XOR2_X1 u0_u15_U33 (.A( u0_FP_49 ) , .B( u0_K16_24 ) , .Z( u0_u15_X_24 ) );
  XOR2_X1 u0_u15_U34 (.A( u0_FP_48 ) , .B( u0_K16_23 ) , .Z( u0_u15_X_23 ) );
  XOR2_X1 u0_u15_U37 (.A( u0_FP_45 ) , .B( u0_K16_20 ) , .Z( u0_u15_X_20 ) );
  XOR2_X1 u0_u15_U38 (.A( u0_FP_64 ) , .B( u0_K16_1 ) , .Z( u0_u15_X_1 ) );
  XOR2_X1 u0_u15_U4 (.A( u0_FP_37 ) , .B( u0_K16_6 ) , .Z( u0_u15_X_6 ) );
  XOR2_X1 u0_u15_U40 (.A( u0_FP_45 ) , .B( u0_K16_18 ) , .Z( u0_u15_X_18 ) );
  XOR2_X1 u0_u15_U42 (.A( u0_FP_43 ) , .B( u0_K16_16 ) , .Z( u0_u15_X_16 ) );
  XOR2_X1 u0_u15_U43 (.A( u0_FP_42 ) , .B( u0_K16_15 ) , .Z( u0_u15_X_15 ) );
  XOR2_X1 u0_u15_U44 (.A( u0_FP_41 ) , .B( u0_K16_14 ) , .Z( u0_u15_X_14 ) );
  XOR2_X1 u0_u15_U45 (.A( u0_FP_40 ) , .B( u0_K16_13 ) , .Z( u0_u15_X_13 ) );
  XOR2_X1 u0_u15_U46 (.A( u0_FP_41 ) , .B( u0_K16_12 ) , .Z( u0_u15_X_12 ) );
  XOR2_X1 u0_u15_U47 (.A( u0_FP_40 ) , .B( u0_K16_11 ) , .Z( u0_u15_X_11 ) );
  XOR2_X1 u0_u15_U48 (.A( u0_FP_39 ) , .B( u0_K16_10 ) , .Z( u0_u15_X_10 ) );
  XOR2_X1 u0_u15_U5 (.A( u0_FP_36 ) , .B( u0_K16_5 ) , .Z( u0_u15_X_5 ) );
  AND3_X1 u0_u15_u0_U10 (.A2( u0_u15_u0_n112 ) , .ZN( u0_u15_u0_n127 ) , .A3( u0_u15_u0_n130 ) , .A1( u0_u15_u0_n148 ) );
  NAND2_X1 u0_u15_u0_U11 (.ZN( u0_u15_u0_n113 ) , .A1( u0_u15_u0_n139 ) , .A2( u0_u15_u0_n149 ) );
  AND2_X1 u0_u15_u0_U12 (.ZN( u0_u15_u0_n107 ) , .A1( u0_u15_u0_n130 ) , .A2( u0_u15_u0_n140 ) );
  AND2_X1 u0_u15_u0_U13 (.A2( u0_u15_u0_n129 ) , .A1( u0_u15_u0_n130 ) , .ZN( u0_u15_u0_n151 ) );
  AND2_X1 u0_u15_u0_U14 (.A1( u0_u15_u0_n108 ) , .A2( u0_u15_u0_n125 ) , .ZN( u0_u15_u0_n145 ) );
  INV_X1 u0_u15_u0_U15 (.A( u0_u15_u0_n143 ) , .ZN( u0_u15_u0_n173 ) );
  NOR2_X1 u0_u15_u0_U16 (.A2( u0_u15_u0_n136 ) , .ZN( u0_u15_u0_n147 ) , .A1( u0_u15_u0_n160 ) );
  AOI21_X1 u0_u15_u0_U17 (.B1( u0_u15_u0_n103 ) , .ZN( u0_u15_u0_n132 ) , .A( u0_u15_u0_n165 ) , .B2( u0_u15_u0_n93 ) );
  INV_X1 u0_u15_u0_U18 (.A( u0_u15_u0_n142 ) , .ZN( u0_u15_u0_n165 ) );
  OAI221_X1 u0_u15_u0_U19 (.C1( u0_u15_u0_n121 ) , .ZN( u0_u15_u0_n122 ) , .B2( u0_u15_u0_n127 ) , .A( u0_u15_u0_n143 ) , .B1( u0_u15_u0_n144 ) , .C2( u0_u15_u0_n147 ) );
  OAI22_X1 u0_u15_u0_U20 (.B1( u0_u15_u0_n131 ) , .A1( u0_u15_u0_n144 ) , .B2( u0_u15_u0_n147 ) , .A2( u0_u15_u0_n90 ) , .ZN( u0_u15_u0_n91 ) );
  AND3_X1 u0_u15_u0_U21 (.A3( u0_u15_u0_n121 ) , .A2( u0_u15_u0_n125 ) , .A1( u0_u15_u0_n148 ) , .ZN( u0_u15_u0_n90 ) );
  OAI22_X1 u0_u15_u0_U22 (.B1( u0_u15_u0_n125 ) , .ZN( u0_u15_u0_n126 ) , .A1( u0_u15_u0_n138 ) , .A2( u0_u15_u0_n146 ) , .B2( u0_u15_u0_n147 ) );
  NOR2_X1 u0_u15_u0_U23 (.A1( u0_u15_u0_n163 ) , .A2( u0_u15_u0_n164 ) , .ZN( u0_u15_u0_n95 ) );
  INV_X1 u0_u15_u0_U24 (.A( u0_u15_u0_n136 ) , .ZN( u0_u15_u0_n161 ) );
  NOR2_X1 u0_u15_u0_U25 (.A1( u0_u15_u0_n120 ) , .ZN( u0_u15_u0_n143 ) , .A2( u0_u15_u0_n167 ) );
  OAI221_X1 u0_u15_u0_U26 (.C1( u0_u15_u0_n112 ) , .ZN( u0_u15_u0_n120 ) , .B1( u0_u15_u0_n138 ) , .B2( u0_u15_u0_n141 ) , .C2( u0_u15_u0_n147 ) , .A( u0_u15_u0_n172 ) );
  AOI211_X1 u0_u15_u0_U27 (.B( u0_u15_u0_n115 ) , .A( u0_u15_u0_n116 ) , .C2( u0_u15_u0_n117 ) , .C1( u0_u15_u0_n118 ) , .ZN( u0_u15_u0_n119 ) );
  AOI22_X1 u0_u15_u0_U28 (.B2( u0_u15_u0_n109 ) , .A2( u0_u15_u0_n110 ) , .ZN( u0_u15_u0_n111 ) , .B1( u0_u15_u0_n118 ) , .A1( u0_u15_u0_n160 ) );
  NAND2_X1 u0_u15_u0_U29 (.A2( u0_u15_u0_n102 ) , .A1( u0_u15_u0_n103 ) , .ZN( u0_u15_u0_n149 ) );
  INV_X1 u0_u15_u0_U3 (.A( u0_u15_u0_n113 ) , .ZN( u0_u15_u0_n166 ) );
  INV_X1 u0_u15_u0_U30 (.A( u0_u15_u0_n118 ) , .ZN( u0_u15_u0_n158 ) );
  NAND2_X1 u0_u15_u0_U31 (.A2( u0_u15_u0_n100 ) , .ZN( u0_u15_u0_n131 ) , .A1( u0_u15_u0_n92 ) );
  NAND2_X1 u0_u15_u0_U32 (.ZN( u0_u15_u0_n108 ) , .A1( u0_u15_u0_n92 ) , .A2( u0_u15_u0_n94 ) );
  AOI21_X1 u0_u15_u0_U33 (.ZN( u0_u15_u0_n104 ) , .B1( u0_u15_u0_n107 ) , .B2( u0_u15_u0_n141 ) , .A( u0_u15_u0_n144 ) );
  AOI21_X1 u0_u15_u0_U34 (.B1( u0_u15_u0_n127 ) , .B2( u0_u15_u0_n129 ) , .A( u0_u15_u0_n138 ) , .ZN( u0_u15_u0_n96 ) );
  NAND2_X1 u0_u15_u0_U35 (.A2( u0_u15_u0_n102 ) , .ZN( u0_u15_u0_n114 ) , .A1( u0_u15_u0_n92 ) );
  AOI21_X1 u0_u15_u0_U36 (.ZN( u0_u15_u0_n116 ) , .B2( u0_u15_u0_n142 ) , .A( u0_u15_u0_n144 ) , .B1( u0_u15_u0_n166 ) );
  NAND2_X1 u0_u15_u0_U37 (.A2( u0_u15_u0_n103 ) , .ZN( u0_u15_u0_n140 ) , .A1( u0_u15_u0_n94 ) );
  NAND2_X1 u0_u15_u0_U38 (.A1( u0_u15_u0_n100 ) , .A2( u0_u15_u0_n103 ) , .ZN( u0_u15_u0_n125 ) );
  NAND2_X1 u0_u15_u0_U39 (.A1( u0_u15_u0_n101 ) , .A2( u0_u15_u0_n102 ) , .ZN( u0_u15_u0_n150 ) );
  AOI21_X1 u0_u15_u0_U4 (.B1( u0_u15_u0_n114 ) , .ZN( u0_u15_u0_n115 ) , .B2( u0_u15_u0_n129 ) , .A( u0_u15_u0_n161 ) );
  INV_X1 u0_u15_u0_U40 (.A( u0_u15_u0_n138 ) , .ZN( u0_u15_u0_n160 ) );
  NAND2_X1 u0_u15_u0_U41 (.A2( u0_u15_u0_n100 ) , .A1( u0_u15_u0_n101 ) , .ZN( u0_u15_u0_n139 ) );
  NAND2_X1 u0_u15_u0_U42 (.ZN( u0_u15_u0_n112 ) , .A2( u0_u15_u0_n92 ) , .A1( u0_u15_u0_n93 ) );
  NAND2_X1 u0_u15_u0_U43 (.A1( u0_u15_u0_n101 ) , .ZN( u0_u15_u0_n130 ) , .A2( u0_u15_u0_n94 ) );
  NAND2_X1 u0_u15_u0_U44 (.A2( u0_u15_u0_n101 ) , .ZN( u0_u15_u0_n121 ) , .A1( u0_u15_u0_n93 ) );
  INV_X1 u0_u15_u0_U45 (.ZN( u0_u15_u0_n172 ) , .A( u0_u15_u0_n88 ) );
  OAI222_X1 u0_u15_u0_U46 (.C1( u0_u15_u0_n108 ) , .A1( u0_u15_u0_n125 ) , .B2( u0_u15_u0_n128 ) , .B1( u0_u15_u0_n144 ) , .A2( u0_u15_u0_n158 ) , .C2( u0_u15_u0_n161 ) , .ZN( u0_u15_u0_n88 ) );
  OR3_X1 u0_u15_u0_U47 (.A3( u0_u15_u0_n152 ) , .A2( u0_u15_u0_n153 ) , .A1( u0_u15_u0_n154 ) , .ZN( u0_u15_u0_n155 ) );
  AOI21_X1 u0_u15_u0_U48 (.B2( u0_u15_u0_n150 ) , .B1( u0_u15_u0_n151 ) , .ZN( u0_u15_u0_n152 ) , .A( u0_u15_u0_n158 ) );
  AOI21_X1 u0_u15_u0_U49 (.A( u0_u15_u0_n144 ) , .B2( u0_u15_u0_n145 ) , .B1( u0_u15_u0_n146 ) , .ZN( u0_u15_u0_n154 ) );
  AOI21_X1 u0_u15_u0_U5 (.B2( u0_u15_u0_n131 ) , .ZN( u0_u15_u0_n134 ) , .B1( u0_u15_u0_n151 ) , .A( u0_u15_u0_n158 ) );
  AOI21_X1 u0_u15_u0_U50 (.A( u0_u15_u0_n147 ) , .B2( u0_u15_u0_n148 ) , .B1( u0_u15_u0_n149 ) , .ZN( u0_u15_u0_n153 ) );
  INV_X1 u0_u15_u0_U51 (.ZN( u0_u15_u0_n171 ) , .A( u0_u15_u0_n99 ) );
  OAI211_X1 u0_u15_u0_U52 (.C2( u0_u15_u0_n140 ) , .C1( u0_u15_u0_n161 ) , .A( u0_u15_u0_n169 ) , .B( u0_u15_u0_n98 ) , .ZN( u0_u15_u0_n99 ) );
  AOI211_X1 u0_u15_u0_U53 (.C1( u0_u15_u0_n118 ) , .A( u0_u15_u0_n123 ) , .B( u0_u15_u0_n96 ) , .C2( u0_u15_u0_n97 ) , .ZN( u0_u15_u0_n98 ) );
  INV_X1 u0_u15_u0_U54 (.ZN( u0_u15_u0_n169 ) , .A( u0_u15_u0_n91 ) );
  NOR2_X1 u0_u15_u0_U55 (.A2( u0_u15_X_4 ) , .A1( u0_u15_X_5 ) , .ZN( u0_u15_u0_n118 ) );
  NOR2_X1 u0_u15_u0_U56 (.A2( u0_u15_X_1 ) , .ZN( u0_u15_u0_n101 ) , .A1( u0_u15_u0_n163 ) );
  NOR2_X1 u0_u15_u0_U57 (.A2( u0_u15_X_3 ) , .A1( u0_u15_X_6 ) , .ZN( u0_u15_u0_n94 ) );
  NOR2_X1 u0_u15_u0_U58 (.A2( u0_u15_X_6 ) , .ZN( u0_u15_u0_n100 ) , .A1( u0_u15_u0_n162 ) );
  NAND2_X1 u0_u15_u0_U59 (.A2( u0_u15_X_4 ) , .A1( u0_u15_X_5 ) , .ZN( u0_u15_u0_n144 ) );
  NOR2_X1 u0_u15_u0_U6 (.A1( u0_u15_u0_n108 ) , .ZN( u0_u15_u0_n123 ) , .A2( u0_u15_u0_n158 ) );
  NOR2_X1 u0_u15_u0_U60 (.A2( u0_u15_X_5 ) , .ZN( u0_u15_u0_n136 ) , .A1( u0_u15_u0_n159 ) );
  NAND2_X1 u0_u15_u0_U61 (.A1( u0_u15_X_5 ) , .ZN( u0_u15_u0_n138 ) , .A2( u0_u15_u0_n159 ) );
  AND2_X1 u0_u15_u0_U62 (.A2( u0_u15_X_3 ) , .A1( u0_u15_X_6 ) , .ZN( u0_u15_u0_n102 ) );
  AND2_X1 u0_u15_u0_U63 (.A1( u0_u15_X_6 ) , .A2( u0_u15_u0_n162 ) , .ZN( u0_u15_u0_n93 ) );
  INV_X1 u0_u15_u0_U64 (.A( u0_u15_X_4 ) , .ZN( u0_u15_u0_n159 ) );
  INV_X1 u0_u15_u0_U65 (.A( u0_u15_X_1 ) , .ZN( u0_u15_u0_n164 ) );
  INV_X1 u0_u15_u0_U66 (.A( u0_u15_X_3 ) , .ZN( u0_u15_u0_n162 ) );
  INV_X1 u0_u15_u0_U67 (.A( u0_u15_u0_n126 ) , .ZN( u0_u15_u0_n168 ) );
  AOI211_X1 u0_u15_u0_U68 (.B( u0_u15_u0_n133 ) , .A( u0_u15_u0_n134 ) , .C2( u0_u15_u0_n135 ) , .C1( u0_u15_u0_n136 ) , .ZN( u0_u15_u0_n137 ) );
  INV_X1 u0_u15_u0_U69 (.ZN( u0_u15_u0_n174 ) , .A( u0_u15_u0_n89 ) );
  OAI21_X1 u0_u15_u0_U7 (.B1( u0_u15_u0_n150 ) , .B2( u0_u15_u0_n158 ) , .A( u0_u15_u0_n172 ) , .ZN( u0_u15_u0_n89 ) );
  AOI211_X1 u0_u15_u0_U70 (.B( u0_u15_u0_n104 ) , .A( u0_u15_u0_n105 ) , .ZN( u0_u15_u0_n106 ) , .C2( u0_u15_u0_n113 ) , .C1( u0_u15_u0_n160 ) );
  OR4_X1 u0_u15_u0_U71 (.ZN( u0_out15_17 ) , .A4( u0_u15_u0_n122 ) , .A2( u0_u15_u0_n123 ) , .A1( u0_u15_u0_n124 ) , .A3( u0_u15_u0_n170 ) );
  AOI21_X1 u0_u15_u0_U72 (.B2( u0_u15_u0_n107 ) , .ZN( u0_u15_u0_n124 ) , .B1( u0_u15_u0_n128 ) , .A( u0_u15_u0_n161 ) );
  INV_X1 u0_u15_u0_U73 (.A( u0_u15_u0_n111 ) , .ZN( u0_u15_u0_n170 ) );
  OR4_X1 u0_u15_u0_U74 (.ZN( u0_out15_31 ) , .A4( u0_u15_u0_n155 ) , .A2( u0_u15_u0_n156 ) , .A1( u0_u15_u0_n157 ) , .A3( u0_u15_u0_n173 ) );
  AOI21_X1 u0_u15_u0_U75 (.A( u0_u15_u0_n138 ) , .B2( u0_u15_u0_n139 ) , .B1( u0_u15_u0_n140 ) , .ZN( u0_u15_u0_n157 ) );
  AOI21_X1 u0_u15_u0_U76 (.B2( u0_u15_u0_n141 ) , .B1( u0_u15_u0_n142 ) , .ZN( u0_u15_u0_n156 ) , .A( u0_u15_u0_n161 ) );
  AOI21_X1 u0_u15_u0_U77 (.B1( u0_u15_u0_n132 ) , .ZN( u0_u15_u0_n133 ) , .A( u0_u15_u0_n144 ) , .B2( u0_u15_u0_n166 ) );
  OAI22_X1 u0_u15_u0_U78 (.ZN( u0_u15_u0_n105 ) , .A2( u0_u15_u0_n132 ) , .B1( u0_u15_u0_n146 ) , .A1( u0_u15_u0_n147 ) , .B2( u0_u15_u0_n161 ) );
  NAND2_X1 u0_u15_u0_U79 (.ZN( u0_u15_u0_n110 ) , .A2( u0_u15_u0_n132 ) , .A1( u0_u15_u0_n145 ) );
  AND2_X1 u0_u15_u0_U8 (.A1( u0_u15_u0_n114 ) , .A2( u0_u15_u0_n121 ) , .ZN( u0_u15_u0_n146 ) );
  INV_X1 u0_u15_u0_U80 (.A( u0_u15_u0_n119 ) , .ZN( u0_u15_u0_n167 ) );
  NAND2_X1 u0_u15_u0_U81 (.ZN( u0_u15_u0_n148 ) , .A1( u0_u15_u0_n93 ) , .A2( u0_u15_u0_n95 ) );
  NAND2_X1 u0_u15_u0_U82 (.A1( u0_u15_u0_n100 ) , .ZN( u0_u15_u0_n129 ) , .A2( u0_u15_u0_n95 ) );
  NAND2_X1 u0_u15_u0_U83 (.A1( u0_u15_u0_n102 ) , .ZN( u0_u15_u0_n128 ) , .A2( u0_u15_u0_n95 ) );
  NOR2_X1 u0_u15_u0_U84 (.A2( u0_u15_X_1 ) , .A1( u0_u15_X_2 ) , .ZN( u0_u15_u0_n92 ) );
  NAND2_X1 u0_u15_u0_U85 (.ZN( u0_u15_u0_n142 ) , .A1( u0_u15_u0_n94 ) , .A2( u0_u15_u0_n95 ) );
  NOR2_X1 u0_u15_u0_U86 (.A2( u0_u15_X_2 ) , .ZN( u0_u15_u0_n103 ) , .A1( u0_u15_u0_n164 ) );
  INV_X1 u0_u15_u0_U87 (.A( u0_u15_X_2 ) , .ZN( u0_u15_u0_n163 ) );
  NAND3_X1 u0_u15_u0_U88 (.ZN( u0_out15_23 ) , .A3( u0_u15_u0_n137 ) , .A1( u0_u15_u0_n168 ) , .A2( u0_u15_u0_n171 ) );
  NAND3_X1 u0_u15_u0_U89 (.A3( u0_u15_u0_n127 ) , .A2( u0_u15_u0_n128 ) , .ZN( u0_u15_u0_n135 ) , .A1( u0_u15_u0_n150 ) );
  AND2_X1 u0_u15_u0_U9 (.A1( u0_u15_u0_n131 ) , .ZN( u0_u15_u0_n141 ) , .A2( u0_u15_u0_n150 ) );
  NAND3_X1 u0_u15_u0_U90 (.ZN( u0_u15_u0_n117 ) , .A3( u0_u15_u0_n132 ) , .A2( u0_u15_u0_n139 ) , .A1( u0_u15_u0_n148 ) );
  NAND3_X1 u0_u15_u0_U91 (.ZN( u0_u15_u0_n109 ) , .A2( u0_u15_u0_n114 ) , .A3( u0_u15_u0_n140 ) , .A1( u0_u15_u0_n149 ) );
  NAND3_X1 u0_u15_u0_U92 (.ZN( u0_out15_9 ) , .A3( u0_u15_u0_n106 ) , .A2( u0_u15_u0_n171 ) , .A1( u0_u15_u0_n174 ) );
  NAND3_X1 u0_u15_u0_U93 (.A2( u0_u15_u0_n128 ) , .A1( u0_u15_u0_n132 ) , .A3( u0_u15_u0_n146 ) , .ZN( u0_u15_u0_n97 ) );
  NOR2_X1 u0_u15_u1_U10 (.A1( u0_u15_u1_n112 ) , .A2( u0_u15_u1_n116 ) , .ZN( u0_u15_u1_n118 ) );
  NAND3_X1 u0_u15_u1_U100 (.ZN( u0_u15_u1_n113 ) , .A1( u0_u15_u1_n120 ) , .A3( u0_u15_u1_n133 ) , .A2( u0_u15_u1_n155 ) );
  OAI21_X1 u0_u15_u1_U11 (.ZN( u0_u15_u1_n101 ) , .B1( u0_u15_u1_n141 ) , .A( u0_u15_u1_n146 ) , .B2( u0_u15_u1_n183 ) );
  AOI21_X1 u0_u15_u1_U12 (.B2( u0_u15_u1_n155 ) , .B1( u0_u15_u1_n156 ) , .ZN( u0_u15_u1_n157 ) , .A( u0_u15_u1_n174 ) );
  NAND2_X1 u0_u15_u1_U13 (.ZN( u0_u15_u1_n140 ) , .A2( u0_u15_u1_n150 ) , .A1( u0_u15_u1_n155 ) );
  NAND2_X1 u0_u15_u1_U14 (.A1( u0_u15_u1_n131 ) , .ZN( u0_u15_u1_n147 ) , .A2( u0_u15_u1_n153 ) );
  INV_X1 u0_u15_u1_U15 (.A( u0_u15_u1_n139 ) , .ZN( u0_u15_u1_n174 ) );
  OR4_X1 u0_u15_u1_U16 (.A4( u0_u15_u1_n106 ) , .A3( u0_u15_u1_n107 ) , .ZN( u0_u15_u1_n108 ) , .A1( u0_u15_u1_n117 ) , .A2( u0_u15_u1_n184 ) );
  AOI21_X1 u0_u15_u1_U17 (.ZN( u0_u15_u1_n106 ) , .A( u0_u15_u1_n112 ) , .B1( u0_u15_u1_n154 ) , .B2( u0_u15_u1_n156 ) );
  AOI21_X1 u0_u15_u1_U18 (.ZN( u0_u15_u1_n107 ) , .B1( u0_u15_u1_n134 ) , .B2( u0_u15_u1_n149 ) , .A( u0_u15_u1_n174 ) );
  INV_X1 u0_u15_u1_U19 (.A( u0_u15_u1_n101 ) , .ZN( u0_u15_u1_n184 ) );
  INV_X1 u0_u15_u1_U20 (.A( u0_u15_u1_n112 ) , .ZN( u0_u15_u1_n171 ) );
  NAND2_X1 u0_u15_u1_U21 (.ZN( u0_u15_u1_n141 ) , .A1( u0_u15_u1_n153 ) , .A2( u0_u15_u1_n156 ) );
  AND2_X1 u0_u15_u1_U22 (.A1( u0_u15_u1_n123 ) , .ZN( u0_u15_u1_n134 ) , .A2( u0_u15_u1_n161 ) );
  NAND2_X1 u0_u15_u1_U23 (.A2( u0_u15_u1_n115 ) , .A1( u0_u15_u1_n116 ) , .ZN( u0_u15_u1_n148 ) );
  NAND2_X1 u0_u15_u1_U24 (.A2( u0_u15_u1_n133 ) , .A1( u0_u15_u1_n135 ) , .ZN( u0_u15_u1_n159 ) );
  NAND2_X1 u0_u15_u1_U25 (.A2( u0_u15_u1_n115 ) , .A1( u0_u15_u1_n120 ) , .ZN( u0_u15_u1_n132 ) );
  INV_X1 u0_u15_u1_U26 (.A( u0_u15_u1_n154 ) , .ZN( u0_u15_u1_n178 ) );
  INV_X1 u0_u15_u1_U27 (.A( u0_u15_u1_n151 ) , .ZN( u0_u15_u1_n183 ) );
  AND2_X1 u0_u15_u1_U28 (.A1( u0_u15_u1_n129 ) , .A2( u0_u15_u1_n133 ) , .ZN( u0_u15_u1_n149 ) );
  INV_X1 u0_u15_u1_U29 (.A( u0_u15_u1_n131 ) , .ZN( u0_u15_u1_n180 ) );
  INV_X1 u0_u15_u1_U3 (.A( u0_u15_u1_n159 ) , .ZN( u0_u15_u1_n182 ) );
  OAI221_X1 u0_u15_u1_U30 (.A( u0_u15_u1_n119 ) , .C2( u0_u15_u1_n129 ) , .ZN( u0_u15_u1_n138 ) , .B2( u0_u15_u1_n152 ) , .C1( u0_u15_u1_n174 ) , .B1( u0_u15_u1_n187 ) );
  INV_X1 u0_u15_u1_U31 (.A( u0_u15_u1_n148 ) , .ZN( u0_u15_u1_n187 ) );
  AOI211_X1 u0_u15_u1_U32 (.B( u0_u15_u1_n117 ) , .A( u0_u15_u1_n118 ) , .ZN( u0_u15_u1_n119 ) , .C2( u0_u15_u1_n146 ) , .C1( u0_u15_u1_n159 ) );
  NOR2_X1 u0_u15_u1_U33 (.A1( u0_u15_u1_n168 ) , .A2( u0_u15_u1_n176 ) , .ZN( u0_u15_u1_n98 ) );
  AOI211_X1 u0_u15_u1_U34 (.B( u0_u15_u1_n162 ) , .A( u0_u15_u1_n163 ) , .C2( u0_u15_u1_n164 ) , .ZN( u0_u15_u1_n165 ) , .C1( u0_u15_u1_n171 ) );
  AOI21_X1 u0_u15_u1_U35 (.A( u0_u15_u1_n160 ) , .B2( u0_u15_u1_n161 ) , .ZN( u0_u15_u1_n162 ) , .B1( u0_u15_u1_n182 ) );
  OR2_X1 u0_u15_u1_U36 (.A2( u0_u15_u1_n157 ) , .A1( u0_u15_u1_n158 ) , .ZN( u0_u15_u1_n163 ) );
  NAND2_X1 u0_u15_u1_U37 (.A1( u0_u15_u1_n128 ) , .ZN( u0_u15_u1_n146 ) , .A2( u0_u15_u1_n160 ) );
  NAND2_X1 u0_u15_u1_U38 (.A2( u0_u15_u1_n112 ) , .ZN( u0_u15_u1_n139 ) , .A1( u0_u15_u1_n152 ) );
  NAND2_X1 u0_u15_u1_U39 (.A1( u0_u15_u1_n105 ) , .ZN( u0_u15_u1_n156 ) , .A2( u0_u15_u1_n99 ) );
  AOI221_X1 u0_u15_u1_U4 (.A( u0_u15_u1_n138 ) , .C2( u0_u15_u1_n139 ) , .C1( u0_u15_u1_n140 ) , .B2( u0_u15_u1_n141 ) , .ZN( u0_u15_u1_n142 ) , .B1( u0_u15_u1_n175 ) );
  AOI221_X1 u0_u15_u1_U40 (.B1( u0_u15_u1_n140 ) , .ZN( u0_u15_u1_n167 ) , .B2( u0_u15_u1_n172 ) , .C2( u0_u15_u1_n175 ) , .C1( u0_u15_u1_n178 ) , .A( u0_u15_u1_n188 ) );
  INV_X1 u0_u15_u1_U41 (.ZN( u0_u15_u1_n188 ) , .A( u0_u15_u1_n97 ) );
  AOI211_X1 u0_u15_u1_U42 (.A( u0_u15_u1_n118 ) , .C1( u0_u15_u1_n132 ) , .C2( u0_u15_u1_n139 ) , .B( u0_u15_u1_n96 ) , .ZN( u0_u15_u1_n97 ) );
  AOI21_X1 u0_u15_u1_U43 (.B2( u0_u15_u1_n121 ) , .B1( u0_u15_u1_n135 ) , .A( u0_u15_u1_n152 ) , .ZN( u0_u15_u1_n96 ) );
  NOR2_X1 u0_u15_u1_U44 (.ZN( u0_u15_u1_n117 ) , .A1( u0_u15_u1_n121 ) , .A2( u0_u15_u1_n160 ) );
  AOI21_X1 u0_u15_u1_U45 (.A( u0_u15_u1_n128 ) , .B2( u0_u15_u1_n129 ) , .ZN( u0_u15_u1_n130 ) , .B1( u0_u15_u1_n150 ) );
  OAI21_X1 u0_u15_u1_U46 (.B2( u0_u15_u1_n123 ) , .ZN( u0_u15_u1_n145 ) , .B1( u0_u15_u1_n160 ) , .A( u0_u15_u1_n185 ) );
  INV_X1 u0_u15_u1_U47 (.A( u0_u15_u1_n122 ) , .ZN( u0_u15_u1_n185 ) );
  AOI21_X1 u0_u15_u1_U48 (.B2( u0_u15_u1_n120 ) , .B1( u0_u15_u1_n121 ) , .ZN( u0_u15_u1_n122 ) , .A( u0_u15_u1_n128 ) );
  NAND2_X1 u0_u15_u1_U49 (.ZN( u0_u15_u1_n112 ) , .A1( u0_u15_u1_n169 ) , .A2( u0_u15_u1_n170 ) );
  AOI211_X1 u0_u15_u1_U5 (.ZN( u0_u15_u1_n124 ) , .A( u0_u15_u1_n138 ) , .C2( u0_u15_u1_n139 ) , .B( u0_u15_u1_n145 ) , .C1( u0_u15_u1_n147 ) );
  NAND2_X1 u0_u15_u1_U50 (.ZN( u0_u15_u1_n129 ) , .A2( u0_u15_u1_n95 ) , .A1( u0_u15_u1_n98 ) );
  NAND2_X1 u0_u15_u1_U51 (.A1( u0_u15_u1_n102 ) , .ZN( u0_u15_u1_n154 ) , .A2( u0_u15_u1_n99 ) );
  NAND2_X1 u0_u15_u1_U52 (.A2( u0_u15_u1_n100 ) , .ZN( u0_u15_u1_n135 ) , .A1( u0_u15_u1_n99 ) );
  AOI21_X1 u0_u15_u1_U53 (.A( u0_u15_u1_n152 ) , .B2( u0_u15_u1_n153 ) , .B1( u0_u15_u1_n154 ) , .ZN( u0_u15_u1_n158 ) );
  INV_X1 u0_u15_u1_U54 (.A( u0_u15_u1_n160 ) , .ZN( u0_u15_u1_n175 ) );
  NAND2_X1 u0_u15_u1_U55 (.A1( u0_u15_u1_n100 ) , .ZN( u0_u15_u1_n116 ) , .A2( u0_u15_u1_n95 ) );
  NAND2_X1 u0_u15_u1_U56 (.A1( u0_u15_u1_n102 ) , .ZN( u0_u15_u1_n131 ) , .A2( u0_u15_u1_n95 ) );
  NAND2_X1 u0_u15_u1_U57 (.A2( u0_u15_u1_n104 ) , .ZN( u0_u15_u1_n121 ) , .A1( u0_u15_u1_n98 ) );
  NAND2_X1 u0_u15_u1_U58 (.A1( u0_u15_u1_n103 ) , .ZN( u0_u15_u1_n153 ) , .A2( u0_u15_u1_n98 ) );
  NAND2_X1 u0_u15_u1_U59 (.A2( u0_u15_u1_n104 ) , .A1( u0_u15_u1_n105 ) , .ZN( u0_u15_u1_n133 ) );
  AOI22_X1 u0_u15_u1_U6 (.B2( u0_u15_u1_n136 ) , .A2( u0_u15_u1_n137 ) , .ZN( u0_u15_u1_n143 ) , .A1( u0_u15_u1_n171 ) , .B1( u0_u15_u1_n173 ) );
  NAND2_X1 u0_u15_u1_U60 (.ZN( u0_u15_u1_n150 ) , .A2( u0_u15_u1_n98 ) , .A1( u0_u15_u1_n99 ) );
  NAND2_X1 u0_u15_u1_U61 (.A1( u0_u15_u1_n105 ) , .ZN( u0_u15_u1_n155 ) , .A2( u0_u15_u1_n95 ) );
  OAI21_X1 u0_u15_u1_U62 (.ZN( u0_u15_u1_n109 ) , .B1( u0_u15_u1_n129 ) , .B2( u0_u15_u1_n160 ) , .A( u0_u15_u1_n167 ) );
  NAND2_X1 u0_u15_u1_U63 (.A2( u0_u15_u1_n100 ) , .A1( u0_u15_u1_n103 ) , .ZN( u0_u15_u1_n120 ) );
  NAND2_X1 u0_u15_u1_U64 (.A1( u0_u15_u1_n102 ) , .A2( u0_u15_u1_n104 ) , .ZN( u0_u15_u1_n115 ) );
  NAND2_X1 u0_u15_u1_U65 (.A2( u0_u15_u1_n100 ) , .A1( u0_u15_u1_n104 ) , .ZN( u0_u15_u1_n151 ) );
  NAND2_X1 u0_u15_u1_U66 (.A2( u0_u15_u1_n103 ) , .A1( u0_u15_u1_n105 ) , .ZN( u0_u15_u1_n161 ) );
  INV_X1 u0_u15_u1_U67 (.A( u0_u15_u1_n152 ) , .ZN( u0_u15_u1_n173 ) );
  INV_X1 u0_u15_u1_U68 (.A( u0_u15_u1_n128 ) , .ZN( u0_u15_u1_n172 ) );
  NAND2_X1 u0_u15_u1_U69 (.A2( u0_u15_u1_n102 ) , .A1( u0_u15_u1_n103 ) , .ZN( u0_u15_u1_n123 ) );
  INV_X1 u0_u15_u1_U7 (.A( u0_u15_u1_n147 ) , .ZN( u0_u15_u1_n181 ) );
  NOR2_X1 u0_u15_u1_U70 (.A2( u0_u15_X_7 ) , .A1( u0_u15_X_8 ) , .ZN( u0_u15_u1_n95 ) );
  NOR2_X1 u0_u15_u1_U71 (.A1( u0_u15_X_12 ) , .A2( u0_u15_X_9 ) , .ZN( u0_u15_u1_n100 ) );
  NOR2_X1 u0_u15_u1_U72 (.A2( u0_u15_X_8 ) , .A1( u0_u15_u1_n177 ) , .ZN( u0_u15_u1_n99 ) );
  NOR2_X1 u0_u15_u1_U73 (.A2( u0_u15_X_12 ) , .ZN( u0_u15_u1_n102 ) , .A1( u0_u15_u1_n176 ) );
  NOR2_X1 u0_u15_u1_U74 (.A2( u0_u15_X_9 ) , .ZN( u0_u15_u1_n105 ) , .A1( u0_u15_u1_n168 ) );
  NAND2_X1 u0_u15_u1_U75 (.A1( u0_u15_X_10 ) , .ZN( u0_u15_u1_n160 ) , .A2( u0_u15_u1_n169 ) );
  NAND2_X1 u0_u15_u1_U76 (.A2( u0_u15_X_10 ) , .A1( u0_u15_X_11 ) , .ZN( u0_u15_u1_n152 ) );
  NAND2_X1 u0_u15_u1_U77 (.A1( u0_u15_X_11 ) , .ZN( u0_u15_u1_n128 ) , .A2( u0_u15_u1_n170 ) );
  AND2_X1 u0_u15_u1_U78 (.A2( u0_u15_X_7 ) , .A1( u0_u15_X_8 ) , .ZN( u0_u15_u1_n104 ) );
  AND2_X1 u0_u15_u1_U79 (.A1( u0_u15_X_8 ) , .ZN( u0_u15_u1_n103 ) , .A2( u0_u15_u1_n177 ) );
  AOI22_X1 u0_u15_u1_U8 (.B2( u0_u15_u1_n113 ) , .A2( u0_u15_u1_n114 ) , .ZN( u0_u15_u1_n125 ) , .A1( u0_u15_u1_n171 ) , .B1( u0_u15_u1_n173 ) );
  INV_X1 u0_u15_u1_U80 (.A( u0_u15_X_10 ) , .ZN( u0_u15_u1_n170 ) );
  INV_X1 u0_u15_u1_U81 (.A( u0_u15_X_9 ) , .ZN( u0_u15_u1_n176 ) );
  INV_X1 u0_u15_u1_U82 (.A( u0_u15_X_11 ) , .ZN( u0_u15_u1_n169 ) );
  INV_X1 u0_u15_u1_U83 (.A( u0_u15_X_12 ) , .ZN( u0_u15_u1_n168 ) );
  INV_X1 u0_u15_u1_U84 (.A( u0_u15_X_7 ) , .ZN( u0_u15_u1_n177 ) );
  NAND4_X1 u0_u15_u1_U85 (.ZN( u0_out15_18 ) , .A4( u0_u15_u1_n165 ) , .A3( u0_u15_u1_n166 ) , .A1( u0_u15_u1_n167 ) , .A2( u0_u15_u1_n186 ) );
  AOI22_X1 u0_u15_u1_U86 (.B2( u0_u15_u1_n146 ) , .B1( u0_u15_u1_n147 ) , .A2( u0_u15_u1_n148 ) , .ZN( u0_u15_u1_n166 ) , .A1( u0_u15_u1_n172 ) );
  INV_X1 u0_u15_u1_U87 (.A( u0_u15_u1_n145 ) , .ZN( u0_u15_u1_n186 ) );
  NAND4_X1 u0_u15_u1_U88 (.ZN( u0_out15_2 ) , .A4( u0_u15_u1_n142 ) , .A3( u0_u15_u1_n143 ) , .A2( u0_u15_u1_n144 ) , .A1( u0_u15_u1_n179 ) );
  OAI21_X1 u0_u15_u1_U89 (.B2( u0_u15_u1_n132 ) , .ZN( u0_u15_u1_n144 ) , .A( u0_u15_u1_n146 ) , .B1( u0_u15_u1_n180 ) );
  NAND2_X1 u0_u15_u1_U9 (.ZN( u0_u15_u1_n114 ) , .A1( u0_u15_u1_n134 ) , .A2( u0_u15_u1_n156 ) );
  INV_X1 u0_u15_u1_U90 (.A( u0_u15_u1_n130 ) , .ZN( u0_u15_u1_n179 ) );
  NAND4_X1 u0_u15_u1_U91 (.ZN( u0_out15_28 ) , .A4( u0_u15_u1_n124 ) , .A3( u0_u15_u1_n125 ) , .A2( u0_u15_u1_n126 ) , .A1( u0_u15_u1_n127 ) );
  OAI21_X1 u0_u15_u1_U92 (.ZN( u0_u15_u1_n127 ) , .B2( u0_u15_u1_n139 ) , .B1( u0_u15_u1_n175 ) , .A( u0_u15_u1_n183 ) );
  OAI21_X1 u0_u15_u1_U93 (.ZN( u0_u15_u1_n126 ) , .B2( u0_u15_u1_n140 ) , .A( u0_u15_u1_n146 ) , .B1( u0_u15_u1_n178 ) );
  OR4_X1 u0_u15_u1_U94 (.ZN( u0_out15_13 ) , .A4( u0_u15_u1_n108 ) , .A3( u0_u15_u1_n109 ) , .A2( u0_u15_u1_n110 ) , .A1( u0_u15_u1_n111 ) );
  AOI21_X1 u0_u15_u1_U95 (.ZN( u0_u15_u1_n111 ) , .A( u0_u15_u1_n128 ) , .B2( u0_u15_u1_n131 ) , .B1( u0_u15_u1_n135 ) );
  AOI21_X1 u0_u15_u1_U96 (.ZN( u0_u15_u1_n110 ) , .A( u0_u15_u1_n116 ) , .B1( u0_u15_u1_n152 ) , .B2( u0_u15_u1_n160 ) );
  NAND3_X1 u0_u15_u1_U97 (.A3( u0_u15_u1_n149 ) , .A2( u0_u15_u1_n150 ) , .A1( u0_u15_u1_n151 ) , .ZN( u0_u15_u1_n164 ) );
  NAND3_X1 u0_u15_u1_U98 (.A3( u0_u15_u1_n134 ) , .A2( u0_u15_u1_n135 ) , .ZN( u0_u15_u1_n136 ) , .A1( u0_u15_u1_n151 ) );
  NAND3_X1 u0_u15_u1_U99 (.A1( u0_u15_u1_n133 ) , .ZN( u0_u15_u1_n137 ) , .A2( u0_u15_u1_n154 ) , .A3( u0_u15_u1_n181 ) );
  OAI22_X1 u0_u15_u2_U10 (.B1( u0_u15_u2_n151 ) , .A2( u0_u15_u2_n152 ) , .A1( u0_u15_u2_n153 ) , .ZN( u0_u15_u2_n160 ) , .B2( u0_u15_u2_n168 ) );
  NAND3_X1 u0_u15_u2_U100 (.A2( u0_u15_u2_n100 ) , .A1( u0_u15_u2_n104 ) , .A3( u0_u15_u2_n138 ) , .ZN( u0_u15_u2_n98 ) );
  NOR3_X1 u0_u15_u2_U11 (.A1( u0_u15_u2_n150 ) , .ZN( u0_u15_u2_n151 ) , .A3( u0_u15_u2_n175 ) , .A2( u0_u15_u2_n188 ) );
  AOI21_X1 u0_u15_u2_U12 (.B2( u0_u15_u2_n123 ) , .ZN( u0_u15_u2_n125 ) , .A( u0_u15_u2_n171 ) , .B1( u0_u15_u2_n184 ) );
  INV_X1 u0_u15_u2_U13 (.A( u0_u15_u2_n150 ) , .ZN( u0_u15_u2_n184 ) );
  AOI21_X1 u0_u15_u2_U14 (.ZN( u0_u15_u2_n144 ) , .B2( u0_u15_u2_n155 ) , .A( u0_u15_u2_n172 ) , .B1( u0_u15_u2_n185 ) );
  AOI21_X1 u0_u15_u2_U15 (.B2( u0_u15_u2_n143 ) , .ZN( u0_u15_u2_n145 ) , .B1( u0_u15_u2_n152 ) , .A( u0_u15_u2_n171 ) );
  INV_X1 u0_u15_u2_U16 (.A( u0_u15_u2_n156 ) , .ZN( u0_u15_u2_n171 ) );
  INV_X1 u0_u15_u2_U17 (.A( u0_u15_u2_n120 ) , .ZN( u0_u15_u2_n188 ) );
  NAND2_X1 u0_u15_u2_U18 (.A2( u0_u15_u2_n122 ) , .ZN( u0_u15_u2_n150 ) , .A1( u0_u15_u2_n152 ) );
  INV_X1 u0_u15_u2_U19 (.A( u0_u15_u2_n153 ) , .ZN( u0_u15_u2_n170 ) );
  INV_X1 u0_u15_u2_U20 (.A( u0_u15_u2_n137 ) , .ZN( u0_u15_u2_n173 ) );
  NAND2_X1 u0_u15_u2_U21 (.A1( u0_u15_u2_n132 ) , .A2( u0_u15_u2_n139 ) , .ZN( u0_u15_u2_n157 ) );
  INV_X1 u0_u15_u2_U22 (.A( u0_u15_u2_n113 ) , .ZN( u0_u15_u2_n178 ) );
  INV_X1 u0_u15_u2_U23 (.A( u0_u15_u2_n139 ) , .ZN( u0_u15_u2_n175 ) );
  INV_X1 u0_u15_u2_U24 (.A( u0_u15_u2_n155 ) , .ZN( u0_u15_u2_n181 ) );
  INV_X1 u0_u15_u2_U25 (.A( u0_u15_u2_n119 ) , .ZN( u0_u15_u2_n177 ) );
  INV_X1 u0_u15_u2_U26 (.A( u0_u15_u2_n116 ) , .ZN( u0_u15_u2_n180 ) );
  INV_X1 u0_u15_u2_U27 (.A( u0_u15_u2_n131 ) , .ZN( u0_u15_u2_n179 ) );
  INV_X1 u0_u15_u2_U28 (.A( u0_u15_u2_n154 ) , .ZN( u0_u15_u2_n176 ) );
  NAND2_X1 u0_u15_u2_U29 (.A2( u0_u15_u2_n116 ) , .A1( u0_u15_u2_n117 ) , .ZN( u0_u15_u2_n118 ) );
  NOR2_X1 u0_u15_u2_U3 (.ZN( u0_u15_u2_n121 ) , .A2( u0_u15_u2_n177 ) , .A1( u0_u15_u2_n180 ) );
  INV_X1 u0_u15_u2_U30 (.A( u0_u15_u2_n132 ) , .ZN( u0_u15_u2_n182 ) );
  INV_X1 u0_u15_u2_U31 (.A( u0_u15_u2_n158 ) , .ZN( u0_u15_u2_n183 ) );
  OAI21_X1 u0_u15_u2_U32 (.A( u0_u15_u2_n156 ) , .B1( u0_u15_u2_n157 ) , .ZN( u0_u15_u2_n158 ) , .B2( u0_u15_u2_n179 ) );
  NOR2_X1 u0_u15_u2_U33 (.ZN( u0_u15_u2_n156 ) , .A1( u0_u15_u2_n166 ) , .A2( u0_u15_u2_n169 ) );
  NOR2_X1 u0_u15_u2_U34 (.A2( u0_u15_u2_n114 ) , .ZN( u0_u15_u2_n137 ) , .A1( u0_u15_u2_n140 ) );
  NOR2_X1 u0_u15_u2_U35 (.A2( u0_u15_u2_n138 ) , .ZN( u0_u15_u2_n153 ) , .A1( u0_u15_u2_n156 ) );
  AOI211_X1 u0_u15_u2_U36 (.ZN( u0_u15_u2_n130 ) , .C1( u0_u15_u2_n138 ) , .C2( u0_u15_u2_n179 ) , .B( u0_u15_u2_n96 ) , .A( u0_u15_u2_n97 ) );
  OAI22_X1 u0_u15_u2_U37 (.B1( u0_u15_u2_n133 ) , .A2( u0_u15_u2_n137 ) , .A1( u0_u15_u2_n152 ) , .B2( u0_u15_u2_n168 ) , .ZN( u0_u15_u2_n97 ) );
  OAI221_X1 u0_u15_u2_U38 (.B1( u0_u15_u2_n113 ) , .C1( u0_u15_u2_n132 ) , .A( u0_u15_u2_n149 ) , .B2( u0_u15_u2_n171 ) , .C2( u0_u15_u2_n172 ) , .ZN( u0_u15_u2_n96 ) );
  OAI221_X1 u0_u15_u2_U39 (.A( u0_u15_u2_n115 ) , .C2( u0_u15_u2_n123 ) , .B2( u0_u15_u2_n143 ) , .B1( u0_u15_u2_n153 ) , .ZN( u0_u15_u2_n163 ) , .C1( u0_u15_u2_n168 ) );
  INV_X1 u0_u15_u2_U4 (.A( u0_u15_u2_n134 ) , .ZN( u0_u15_u2_n185 ) );
  OAI21_X1 u0_u15_u2_U40 (.A( u0_u15_u2_n114 ) , .ZN( u0_u15_u2_n115 ) , .B1( u0_u15_u2_n176 ) , .B2( u0_u15_u2_n178 ) );
  OAI221_X1 u0_u15_u2_U41 (.A( u0_u15_u2_n135 ) , .B2( u0_u15_u2_n136 ) , .B1( u0_u15_u2_n137 ) , .ZN( u0_u15_u2_n162 ) , .C2( u0_u15_u2_n167 ) , .C1( u0_u15_u2_n185 ) );
  AND3_X1 u0_u15_u2_U42 (.A3( u0_u15_u2_n131 ) , .A2( u0_u15_u2_n132 ) , .A1( u0_u15_u2_n133 ) , .ZN( u0_u15_u2_n136 ) );
  AOI22_X1 u0_u15_u2_U43 (.ZN( u0_u15_u2_n135 ) , .B1( u0_u15_u2_n140 ) , .A1( u0_u15_u2_n156 ) , .B2( u0_u15_u2_n180 ) , .A2( u0_u15_u2_n188 ) );
  AOI21_X1 u0_u15_u2_U44 (.ZN( u0_u15_u2_n149 ) , .B1( u0_u15_u2_n173 ) , .B2( u0_u15_u2_n188 ) , .A( u0_u15_u2_n95 ) );
  AND3_X1 u0_u15_u2_U45 (.A2( u0_u15_u2_n100 ) , .A1( u0_u15_u2_n104 ) , .A3( u0_u15_u2_n156 ) , .ZN( u0_u15_u2_n95 ) );
  OAI21_X1 u0_u15_u2_U46 (.A( u0_u15_u2_n141 ) , .B2( u0_u15_u2_n142 ) , .ZN( u0_u15_u2_n146 ) , .B1( u0_u15_u2_n153 ) );
  OAI21_X1 u0_u15_u2_U47 (.A( u0_u15_u2_n140 ) , .ZN( u0_u15_u2_n141 ) , .B1( u0_u15_u2_n176 ) , .B2( u0_u15_u2_n177 ) );
  NOR3_X1 u0_u15_u2_U48 (.ZN( u0_u15_u2_n142 ) , .A3( u0_u15_u2_n175 ) , .A2( u0_u15_u2_n178 ) , .A1( u0_u15_u2_n181 ) );
  OAI21_X1 u0_u15_u2_U49 (.A( u0_u15_u2_n101 ) , .B2( u0_u15_u2_n121 ) , .B1( u0_u15_u2_n153 ) , .ZN( u0_u15_u2_n164 ) );
  NOR4_X1 u0_u15_u2_U5 (.A4( u0_u15_u2_n124 ) , .A3( u0_u15_u2_n125 ) , .A2( u0_u15_u2_n126 ) , .A1( u0_u15_u2_n127 ) , .ZN( u0_u15_u2_n128 ) );
  NAND2_X1 u0_u15_u2_U50 (.A2( u0_u15_u2_n100 ) , .A1( u0_u15_u2_n107 ) , .ZN( u0_u15_u2_n155 ) );
  NAND2_X1 u0_u15_u2_U51 (.A2( u0_u15_u2_n105 ) , .A1( u0_u15_u2_n108 ) , .ZN( u0_u15_u2_n143 ) );
  NAND2_X1 u0_u15_u2_U52 (.A1( u0_u15_u2_n104 ) , .A2( u0_u15_u2_n106 ) , .ZN( u0_u15_u2_n152 ) );
  NAND2_X1 u0_u15_u2_U53 (.A1( u0_u15_u2_n100 ) , .A2( u0_u15_u2_n105 ) , .ZN( u0_u15_u2_n132 ) );
  INV_X1 u0_u15_u2_U54 (.A( u0_u15_u2_n140 ) , .ZN( u0_u15_u2_n168 ) );
  INV_X1 u0_u15_u2_U55 (.A( u0_u15_u2_n138 ) , .ZN( u0_u15_u2_n167 ) );
  INV_X1 u0_u15_u2_U56 (.ZN( u0_u15_u2_n187 ) , .A( u0_u15_u2_n99 ) );
  OAI21_X1 u0_u15_u2_U57 (.B1( u0_u15_u2_n137 ) , .B2( u0_u15_u2_n143 ) , .A( u0_u15_u2_n98 ) , .ZN( u0_u15_u2_n99 ) );
  NAND2_X1 u0_u15_u2_U58 (.A1( u0_u15_u2_n102 ) , .A2( u0_u15_u2_n106 ) , .ZN( u0_u15_u2_n113 ) );
  NAND2_X1 u0_u15_u2_U59 (.A1( u0_u15_u2_n106 ) , .A2( u0_u15_u2_n107 ) , .ZN( u0_u15_u2_n131 ) );
  AOI21_X1 u0_u15_u2_U6 (.B2( u0_u15_u2_n119 ) , .ZN( u0_u15_u2_n127 ) , .A( u0_u15_u2_n137 ) , .B1( u0_u15_u2_n155 ) );
  NAND2_X1 u0_u15_u2_U60 (.A1( u0_u15_u2_n103 ) , .A2( u0_u15_u2_n107 ) , .ZN( u0_u15_u2_n139 ) );
  NAND2_X1 u0_u15_u2_U61 (.A1( u0_u15_u2_n103 ) , .A2( u0_u15_u2_n105 ) , .ZN( u0_u15_u2_n133 ) );
  NAND2_X1 u0_u15_u2_U62 (.A1( u0_u15_u2_n102 ) , .A2( u0_u15_u2_n103 ) , .ZN( u0_u15_u2_n154 ) );
  NAND2_X1 u0_u15_u2_U63 (.A2( u0_u15_u2_n103 ) , .A1( u0_u15_u2_n104 ) , .ZN( u0_u15_u2_n119 ) );
  NAND2_X1 u0_u15_u2_U64 (.A2( u0_u15_u2_n107 ) , .A1( u0_u15_u2_n108 ) , .ZN( u0_u15_u2_n123 ) );
  NAND2_X1 u0_u15_u2_U65 (.A1( u0_u15_u2_n104 ) , .A2( u0_u15_u2_n108 ) , .ZN( u0_u15_u2_n122 ) );
  INV_X1 u0_u15_u2_U66 (.A( u0_u15_u2_n114 ) , .ZN( u0_u15_u2_n172 ) );
  NAND2_X1 u0_u15_u2_U67 (.A2( u0_u15_u2_n100 ) , .A1( u0_u15_u2_n102 ) , .ZN( u0_u15_u2_n116 ) );
  NAND2_X1 u0_u15_u2_U68 (.A1( u0_u15_u2_n102 ) , .A2( u0_u15_u2_n108 ) , .ZN( u0_u15_u2_n120 ) );
  NAND2_X1 u0_u15_u2_U69 (.A2( u0_u15_u2_n105 ) , .A1( u0_u15_u2_n106 ) , .ZN( u0_u15_u2_n117 ) );
  AOI21_X1 u0_u15_u2_U7 (.ZN( u0_u15_u2_n124 ) , .B1( u0_u15_u2_n131 ) , .B2( u0_u15_u2_n143 ) , .A( u0_u15_u2_n172 ) );
  NOR2_X1 u0_u15_u2_U70 (.A2( u0_u15_X_16 ) , .ZN( u0_u15_u2_n140 ) , .A1( u0_u15_u2_n166 ) );
  NOR2_X1 u0_u15_u2_U71 (.A2( u0_u15_X_13 ) , .A1( u0_u15_X_14 ) , .ZN( u0_u15_u2_n100 ) );
  NOR2_X1 u0_u15_u2_U72 (.A2( u0_u15_X_16 ) , .A1( u0_u15_X_17 ) , .ZN( u0_u15_u2_n138 ) );
  NOR2_X1 u0_u15_u2_U73 (.A2( u0_u15_X_15 ) , .A1( u0_u15_X_18 ) , .ZN( u0_u15_u2_n104 ) );
  NOR2_X1 u0_u15_u2_U74 (.A2( u0_u15_X_14 ) , .ZN( u0_u15_u2_n103 ) , .A1( u0_u15_u2_n174 ) );
  NOR2_X1 u0_u15_u2_U75 (.A2( u0_u15_X_15 ) , .ZN( u0_u15_u2_n102 ) , .A1( u0_u15_u2_n165 ) );
  NOR2_X1 u0_u15_u2_U76 (.A2( u0_u15_X_17 ) , .ZN( u0_u15_u2_n114 ) , .A1( u0_u15_u2_n169 ) );
  AND2_X1 u0_u15_u2_U77 (.A1( u0_u15_X_15 ) , .ZN( u0_u15_u2_n105 ) , .A2( u0_u15_u2_n165 ) );
  AND2_X1 u0_u15_u2_U78 (.A2( u0_u15_X_15 ) , .A1( u0_u15_X_18 ) , .ZN( u0_u15_u2_n107 ) );
  AND2_X1 u0_u15_u2_U79 (.A1( u0_u15_X_14 ) , .ZN( u0_u15_u2_n106 ) , .A2( u0_u15_u2_n174 ) );
  AOI21_X1 u0_u15_u2_U8 (.B2( u0_u15_u2_n120 ) , .B1( u0_u15_u2_n121 ) , .ZN( u0_u15_u2_n126 ) , .A( u0_u15_u2_n167 ) );
  AND2_X1 u0_u15_u2_U80 (.A1( u0_u15_X_13 ) , .A2( u0_u15_X_14 ) , .ZN( u0_u15_u2_n108 ) );
  INV_X1 u0_u15_u2_U81 (.A( u0_u15_X_16 ) , .ZN( u0_u15_u2_n169 ) );
  INV_X1 u0_u15_u2_U82 (.A( u0_u15_X_17 ) , .ZN( u0_u15_u2_n166 ) );
  INV_X1 u0_u15_u2_U83 (.A( u0_u15_X_13 ) , .ZN( u0_u15_u2_n174 ) );
  INV_X1 u0_u15_u2_U84 (.A( u0_u15_X_18 ) , .ZN( u0_u15_u2_n165 ) );
  NAND4_X1 u0_u15_u2_U85 (.ZN( u0_out15_30 ) , .A4( u0_u15_u2_n147 ) , .A3( u0_u15_u2_n148 ) , .A2( u0_u15_u2_n149 ) , .A1( u0_u15_u2_n187 ) );
  NOR3_X1 u0_u15_u2_U86 (.A3( u0_u15_u2_n144 ) , .A2( u0_u15_u2_n145 ) , .A1( u0_u15_u2_n146 ) , .ZN( u0_u15_u2_n147 ) );
  AOI21_X1 u0_u15_u2_U87 (.B2( u0_u15_u2_n138 ) , .ZN( u0_u15_u2_n148 ) , .A( u0_u15_u2_n162 ) , .B1( u0_u15_u2_n182 ) );
  NAND4_X1 u0_u15_u2_U88 (.ZN( u0_out15_24 ) , .A4( u0_u15_u2_n111 ) , .A3( u0_u15_u2_n112 ) , .A1( u0_u15_u2_n130 ) , .A2( u0_u15_u2_n187 ) );
  AOI221_X1 u0_u15_u2_U89 (.A( u0_u15_u2_n109 ) , .B1( u0_u15_u2_n110 ) , .ZN( u0_u15_u2_n111 ) , .C1( u0_u15_u2_n134 ) , .C2( u0_u15_u2_n170 ) , .B2( u0_u15_u2_n173 ) );
  OAI22_X1 u0_u15_u2_U9 (.ZN( u0_u15_u2_n109 ) , .A2( u0_u15_u2_n113 ) , .B2( u0_u15_u2_n133 ) , .B1( u0_u15_u2_n167 ) , .A1( u0_u15_u2_n168 ) );
  AOI21_X1 u0_u15_u2_U90 (.ZN( u0_u15_u2_n112 ) , .B2( u0_u15_u2_n156 ) , .A( u0_u15_u2_n164 ) , .B1( u0_u15_u2_n181 ) );
  NAND4_X1 u0_u15_u2_U91 (.ZN( u0_out15_16 ) , .A4( u0_u15_u2_n128 ) , .A3( u0_u15_u2_n129 ) , .A1( u0_u15_u2_n130 ) , .A2( u0_u15_u2_n186 ) );
  AOI22_X1 u0_u15_u2_U92 (.A2( u0_u15_u2_n118 ) , .ZN( u0_u15_u2_n129 ) , .A1( u0_u15_u2_n140 ) , .B1( u0_u15_u2_n157 ) , .B2( u0_u15_u2_n170 ) );
  INV_X1 u0_u15_u2_U93 (.A( u0_u15_u2_n163 ) , .ZN( u0_u15_u2_n186 ) );
  OR4_X1 u0_u15_u2_U94 (.ZN( u0_out15_6 ) , .A4( u0_u15_u2_n161 ) , .A3( u0_u15_u2_n162 ) , .A2( u0_u15_u2_n163 ) , .A1( u0_u15_u2_n164 ) );
  OR3_X1 u0_u15_u2_U95 (.A2( u0_u15_u2_n159 ) , .A1( u0_u15_u2_n160 ) , .ZN( u0_u15_u2_n161 ) , .A3( u0_u15_u2_n183 ) );
  AOI21_X1 u0_u15_u2_U96 (.B2( u0_u15_u2_n154 ) , .B1( u0_u15_u2_n155 ) , .ZN( u0_u15_u2_n159 ) , .A( u0_u15_u2_n167 ) );
  NAND3_X1 u0_u15_u2_U97 (.A2( u0_u15_u2_n117 ) , .A1( u0_u15_u2_n122 ) , .A3( u0_u15_u2_n123 ) , .ZN( u0_u15_u2_n134 ) );
  NAND3_X1 u0_u15_u2_U98 (.ZN( u0_u15_u2_n110 ) , .A2( u0_u15_u2_n131 ) , .A3( u0_u15_u2_n139 ) , .A1( u0_u15_u2_n154 ) );
  NAND3_X1 u0_u15_u2_U99 (.A2( u0_u15_u2_n100 ) , .ZN( u0_u15_u2_n101 ) , .A1( u0_u15_u2_n104 ) , .A3( u0_u15_u2_n114 ) );
  OAI22_X1 u0_u15_u3_U10 (.B1( u0_u15_u3_n113 ) , .A2( u0_u15_u3_n135 ) , .A1( u0_u15_u3_n150 ) , .B2( u0_u15_u3_n164 ) , .ZN( u0_u15_u3_n98 ) );
  OAI211_X1 u0_u15_u3_U11 (.B( u0_u15_u3_n106 ) , .ZN( u0_u15_u3_n119 ) , .C2( u0_u15_u3_n128 ) , .C1( u0_u15_u3_n167 ) , .A( u0_u15_u3_n181 ) );
  AOI221_X1 u0_u15_u3_U12 (.C1( u0_u15_u3_n105 ) , .ZN( u0_u15_u3_n106 ) , .A( u0_u15_u3_n131 ) , .B2( u0_u15_u3_n132 ) , .C2( u0_u15_u3_n133 ) , .B1( u0_u15_u3_n169 ) );
  INV_X1 u0_u15_u3_U13 (.ZN( u0_u15_u3_n181 ) , .A( u0_u15_u3_n98 ) );
  NAND2_X1 u0_u15_u3_U14 (.ZN( u0_u15_u3_n105 ) , .A2( u0_u15_u3_n130 ) , .A1( u0_u15_u3_n155 ) );
  AOI22_X1 u0_u15_u3_U15 (.B1( u0_u15_u3_n115 ) , .A2( u0_u15_u3_n116 ) , .ZN( u0_u15_u3_n123 ) , .B2( u0_u15_u3_n133 ) , .A1( u0_u15_u3_n169 ) );
  NAND2_X1 u0_u15_u3_U16 (.ZN( u0_u15_u3_n116 ) , .A2( u0_u15_u3_n151 ) , .A1( u0_u15_u3_n182 ) );
  NOR2_X1 u0_u15_u3_U17 (.ZN( u0_u15_u3_n126 ) , .A2( u0_u15_u3_n150 ) , .A1( u0_u15_u3_n164 ) );
  AOI21_X1 u0_u15_u3_U18 (.ZN( u0_u15_u3_n112 ) , .B2( u0_u15_u3_n146 ) , .B1( u0_u15_u3_n155 ) , .A( u0_u15_u3_n167 ) );
  NAND2_X1 u0_u15_u3_U19 (.A1( u0_u15_u3_n135 ) , .ZN( u0_u15_u3_n142 ) , .A2( u0_u15_u3_n164 ) );
  NAND2_X1 u0_u15_u3_U20 (.ZN( u0_u15_u3_n132 ) , .A2( u0_u15_u3_n152 ) , .A1( u0_u15_u3_n156 ) );
  AND2_X1 u0_u15_u3_U21 (.A2( u0_u15_u3_n113 ) , .A1( u0_u15_u3_n114 ) , .ZN( u0_u15_u3_n151 ) );
  INV_X1 u0_u15_u3_U22 (.A( u0_u15_u3_n133 ) , .ZN( u0_u15_u3_n165 ) );
  INV_X1 u0_u15_u3_U23 (.A( u0_u15_u3_n135 ) , .ZN( u0_u15_u3_n170 ) );
  NAND2_X1 u0_u15_u3_U24 (.A1( u0_u15_u3_n107 ) , .A2( u0_u15_u3_n108 ) , .ZN( u0_u15_u3_n140 ) );
  NAND2_X1 u0_u15_u3_U25 (.ZN( u0_u15_u3_n117 ) , .A1( u0_u15_u3_n124 ) , .A2( u0_u15_u3_n148 ) );
  NAND2_X1 u0_u15_u3_U26 (.ZN( u0_u15_u3_n143 ) , .A1( u0_u15_u3_n165 ) , .A2( u0_u15_u3_n167 ) );
  INV_X1 u0_u15_u3_U27 (.A( u0_u15_u3_n130 ) , .ZN( u0_u15_u3_n177 ) );
  INV_X1 u0_u15_u3_U28 (.A( u0_u15_u3_n128 ) , .ZN( u0_u15_u3_n176 ) );
  INV_X1 u0_u15_u3_U29 (.A( u0_u15_u3_n155 ) , .ZN( u0_u15_u3_n174 ) );
  INV_X1 u0_u15_u3_U3 (.A( u0_u15_u3_n129 ) , .ZN( u0_u15_u3_n183 ) );
  INV_X1 u0_u15_u3_U30 (.A( u0_u15_u3_n139 ) , .ZN( u0_u15_u3_n185 ) );
  NOR2_X1 u0_u15_u3_U31 (.ZN( u0_u15_u3_n135 ) , .A2( u0_u15_u3_n141 ) , .A1( u0_u15_u3_n169 ) );
  OAI222_X1 u0_u15_u3_U32 (.C2( u0_u15_u3_n107 ) , .A2( u0_u15_u3_n108 ) , .B1( u0_u15_u3_n135 ) , .ZN( u0_u15_u3_n138 ) , .B2( u0_u15_u3_n146 ) , .C1( u0_u15_u3_n154 ) , .A1( u0_u15_u3_n164 ) );
  NOR4_X1 u0_u15_u3_U33 (.A4( u0_u15_u3_n157 ) , .A3( u0_u15_u3_n158 ) , .A2( u0_u15_u3_n159 ) , .A1( u0_u15_u3_n160 ) , .ZN( u0_u15_u3_n161 ) );
  AOI21_X1 u0_u15_u3_U34 (.B2( u0_u15_u3_n152 ) , .B1( u0_u15_u3_n153 ) , .ZN( u0_u15_u3_n158 ) , .A( u0_u15_u3_n164 ) );
  AOI21_X1 u0_u15_u3_U35 (.A( u0_u15_u3_n154 ) , .B2( u0_u15_u3_n155 ) , .B1( u0_u15_u3_n156 ) , .ZN( u0_u15_u3_n157 ) );
  AOI21_X1 u0_u15_u3_U36 (.A( u0_u15_u3_n149 ) , .B2( u0_u15_u3_n150 ) , .B1( u0_u15_u3_n151 ) , .ZN( u0_u15_u3_n159 ) );
  AOI211_X1 u0_u15_u3_U37 (.ZN( u0_u15_u3_n109 ) , .A( u0_u15_u3_n119 ) , .C2( u0_u15_u3_n129 ) , .B( u0_u15_u3_n138 ) , .C1( u0_u15_u3_n141 ) );
  AOI211_X1 u0_u15_u3_U38 (.B( u0_u15_u3_n119 ) , .A( u0_u15_u3_n120 ) , .C2( u0_u15_u3_n121 ) , .ZN( u0_u15_u3_n122 ) , .C1( u0_u15_u3_n179 ) );
  INV_X1 u0_u15_u3_U39 (.A( u0_u15_u3_n156 ) , .ZN( u0_u15_u3_n179 ) );
  INV_X1 u0_u15_u3_U4 (.A( u0_u15_u3_n140 ) , .ZN( u0_u15_u3_n182 ) );
  OAI22_X1 u0_u15_u3_U40 (.B1( u0_u15_u3_n118 ) , .ZN( u0_u15_u3_n120 ) , .A1( u0_u15_u3_n135 ) , .B2( u0_u15_u3_n154 ) , .A2( u0_u15_u3_n178 ) );
  AND3_X1 u0_u15_u3_U41 (.ZN( u0_u15_u3_n118 ) , .A2( u0_u15_u3_n124 ) , .A1( u0_u15_u3_n144 ) , .A3( u0_u15_u3_n152 ) );
  INV_X1 u0_u15_u3_U42 (.A( u0_u15_u3_n121 ) , .ZN( u0_u15_u3_n164 ) );
  NAND2_X1 u0_u15_u3_U43 (.ZN( u0_u15_u3_n133 ) , .A1( u0_u15_u3_n154 ) , .A2( u0_u15_u3_n164 ) );
  OAI211_X1 u0_u15_u3_U44 (.B( u0_u15_u3_n127 ) , .ZN( u0_u15_u3_n139 ) , .C1( u0_u15_u3_n150 ) , .C2( u0_u15_u3_n154 ) , .A( u0_u15_u3_n184 ) );
  INV_X1 u0_u15_u3_U45 (.A( u0_u15_u3_n125 ) , .ZN( u0_u15_u3_n184 ) );
  AOI221_X1 u0_u15_u3_U46 (.A( u0_u15_u3_n126 ) , .ZN( u0_u15_u3_n127 ) , .C2( u0_u15_u3_n132 ) , .C1( u0_u15_u3_n169 ) , .B2( u0_u15_u3_n170 ) , .B1( u0_u15_u3_n174 ) );
  OAI22_X1 u0_u15_u3_U47 (.A1( u0_u15_u3_n124 ) , .ZN( u0_u15_u3_n125 ) , .B2( u0_u15_u3_n145 ) , .A2( u0_u15_u3_n165 ) , .B1( u0_u15_u3_n167 ) );
  NOR2_X1 u0_u15_u3_U48 (.A1( u0_u15_u3_n113 ) , .ZN( u0_u15_u3_n131 ) , .A2( u0_u15_u3_n154 ) );
  NAND2_X1 u0_u15_u3_U49 (.A1( u0_u15_u3_n103 ) , .ZN( u0_u15_u3_n150 ) , .A2( u0_u15_u3_n99 ) );
  INV_X1 u0_u15_u3_U5 (.A( u0_u15_u3_n117 ) , .ZN( u0_u15_u3_n178 ) );
  NAND2_X1 u0_u15_u3_U50 (.A2( u0_u15_u3_n102 ) , .ZN( u0_u15_u3_n155 ) , .A1( u0_u15_u3_n97 ) );
  INV_X1 u0_u15_u3_U51 (.A( u0_u15_u3_n141 ) , .ZN( u0_u15_u3_n167 ) );
  AOI21_X1 u0_u15_u3_U52 (.B2( u0_u15_u3_n114 ) , .B1( u0_u15_u3_n146 ) , .A( u0_u15_u3_n154 ) , .ZN( u0_u15_u3_n94 ) );
  AOI21_X1 u0_u15_u3_U53 (.ZN( u0_u15_u3_n110 ) , .B2( u0_u15_u3_n142 ) , .B1( u0_u15_u3_n186 ) , .A( u0_u15_u3_n95 ) );
  INV_X1 u0_u15_u3_U54 (.A( u0_u15_u3_n145 ) , .ZN( u0_u15_u3_n186 ) );
  AOI21_X1 u0_u15_u3_U55 (.B1( u0_u15_u3_n124 ) , .A( u0_u15_u3_n149 ) , .B2( u0_u15_u3_n155 ) , .ZN( u0_u15_u3_n95 ) );
  INV_X1 u0_u15_u3_U56 (.A( u0_u15_u3_n149 ) , .ZN( u0_u15_u3_n169 ) );
  NAND2_X1 u0_u15_u3_U57 (.ZN( u0_u15_u3_n124 ) , .A1( u0_u15_u3_n96 ) , .A2( u0_u15_u3_n97 ) );
  NAND2_X1 u0_u15_u3_U58 (.A2( u0_u15_u3_n100 ) , .ZN( u0_u15_u3_n146 ) , .A1( u0_u15_u3_n96 ) );
  NAND2_X1 u0_u15_u3_U59 (.A1( u0_u15_u3_n101 ) , .ZN( u0_u15_u3_n145 ) , .A2( u0_u15_u3_n99 ) );
  AOI221_X1 u0_u15_u3_U6 (.A( u0_u15_u3_n131 ) , .C2( u0_u15_u3_n132 ) , .C1( u0_u15_u3_n133 ) , .ZN( u0_u15_u3_n134 ) , .B1( u0_u15_u3_n143 ) , .B2( u0_u15_u3_n177 ) );
  NAND2_X1 u0_u15_u3_U60 (.A1( u0_u15_u3_n100 ) , .ZN( u0_u15_u3_n156 ) , .A2( u0_u15_u3_n99 ) );
  NAND2_X1 u0_u15_u3_U61 (.A2( u0_u15_u3_n101 ) , .A1( u0_u15_u3_n104 ) , .ZN( u0_u15_u3_n148 ) );
  NAND2_X1 u0_u15_u3_U62 (.A1( u0_u15_u3_n100 ) , .A2( u0_u15_u3_n102 ) , .ZN( u0_u15_u3_n128 ) );
  NAND2_X1 u0_u15_u3_U63 (.A2( u0_u15_u3_n101 ) , .A1( u0_u15_u3_n102 ) , .ZN( u0_u15_u3_n152 ) );
  NAND2_X1 u0_u15_u3_U64 (.A2( u0_u15_u3_n101 ) , .ZN( u0_u15_u3_n114 ) , .A1( u0_u15_u3_n96 ) );
  NAND2_X1 u0_u15_u3_U65 (.ZN( u0_u15_u3_n107 ) , .A1( u0_u15_u3_n97 ) , .A2( u0_u15_u3_n99 ) );
  NAND2_X1 u0_u15_u3_U66 (.A2( u0_u15_u3_n100 ) , .A1( u0_u15_u3_n104 ) , .ZN( u0_u15_u3_n113 ) );
  NAND2_X1 u0_u15_u3_U67 (.A1( u0_u15_u3_n104 ) , .ZN( u0_u15_u3_n153 ) , .A2( u0_u15_u3_n97 ) );
  NAND2_X1 u0_u15_u3_U68 (.A2( u0_u15_u3_n103 ) , .A1( u0_u15_u3_n104 ) , .ZN( u0_u15_u3_n130 ) );
  NAND2_X1 u0_u15_u3_U69 (.A2( u0_u15_u3_n103 ) , .ZN( u0_u15_u3_n144 ) , .A1( u0_u15_u3_n96 ) );
  OAI22_X1 u0_u15_u3_U7 (.B2( u0_u15_u3_n147 ) , .A2( u0_u15_u3_n148 ) , .ZN( u0_u15_u3_n160 ) , .B1( u0_u15_u3_n165 ) , .A1( u0_u15_u3_n168 ) );
  NAND2_X1 u0_u15_u3_U70 (.A1( u0_u15_u3_n102 ) , .A2( u0_u15_u3_n103 ) , .ZN( u0_u15_u3_n108 ) );
  NOR2_X1 u0_u15_u3_U71 (.A2( u0_u15_X_19 ) , .A1( u0_u15_X_20 ) , .ZN( u0_u15_u3_n99 ) );
  NOR2_X1 u0_u15_u3_U72 (.A2( u0_u15_X_21 ) , .A1( u0_u15_X_24 ) , .ZN( u0_u15_u3_n103 ) );
  NOR2_X1 u0_u15_u3_U73 (.A2( u0_u15_X_24 ) , .A1( u0_u15_u3_n171 ) , .ZN( u0_u15_u3_n97 ) );
  NOR2_X1 u0_u15_u3_U74 (.A2( u0_u15_X_23 ) , .ZN( u0_u15_u3_n141 ) , .A1( u0_u15_u3_n166 ) );
  NOR2_X1 u0_u15_u3_U75 (.A2( u0_u15_X_19 ) , .A1( u0_u15_u3_n172 ) , .ZN( u0_u15_u3_n96 ) );
  NAND2_X1 u0_u15_u3_U76 (.A1( u0_u15_X_22 ) , .A2( u0_u15_X_23 ) , .ZN( u0_u15_u3_n154 ) );
  NAND2_X1 u0_u15_u3_U77 (.A1( u0_u15_X_23 ) , .ZN( u0_u15_u3_n149 ) , .A2( u0_u15_u3_n166 ) );
  NOR2_X1 u0_u15_u3_U78 (.A2( u0_u15_X_22 ) , .A1( u0_u15_X_23 ) , .ZN( u0_u15_u3_n121 ) );
  AND2_X1 u0_u15_u3_U79 (.A1( u0_u15_X_24 ) , .ZN( u0_u15_u3_n101 ) , .A2( u0_u15_u3_n171 ) );
  AND3_X1 u0_u15_u3_U8 (.A3( u0_u15_u3_n144 ) , .A2( u0_u15_u3_n145 ) , .A1( u0_u15_u3_n146 ) , .ZN( u0_u15_u3_n147 ) );
  AND2_X1 u0_u15_u3_U80 (.A1( u0_u15_X_19 ) , .ZN( u0_u15_u3_n102 ) , .A2( u0_u15_u3_n172 ) );
  AND2_X1 u0_u15_u3_U81 (.A1( u0_u15_X_21 ) , .A2( u0_u15_X_24 ) , .ZN( u0_u15_u3_n100 ) );
  AND2_X1 u0_u15_u3_U82 (.A2( u0_u15_X_19 ) , .A1( u0_u15_X_20 ) , .ZN( u0_u15_u3_n104 ) );
  INV_X1 u0_u15_u3_U83 (.A( u0_u15_X_22 ) , .ZN( u0_u15_u3_n166 ) );
  INV_X1 u0_u15_u3_U84 (.A( u0_u15_X_21 ) , .ZN( u0_u15_u3_n171 ) );
  INV_X1 u0_u15_u3_U85 (.A( u0_u15_X_20 ) , .ZN( u0_u15_u3_n172 ) );
  OR4_X1 u0_u15_u3_U86 (.ZN( u0_out15_10 ) , .A4( u0_u15_u3_n136 ) , .A3( u0_u15_u3_n137 ) , .A1( u0_u15_u3_n138 ) , .A2( u0_u15_u3_n139 ) );
  OAI222_X1 u0_u15_u3_U87 (.C1( u0_u15_u3_n128 ) , .ZN( u0_u15_u3_n137 ) , .B1( u0_u15_u3_n148 ) , .A2( u0_u15_u3_n150 ) , .B2( u0_u15_u3_n154 ) , .C2( u0_u15_u3_n164 ) , .A1( u0_u15_u3_n167 ) );
  OAI221_X1 u0_u15_u3_U88 (.A( u0_u15_u3_n134 ) , .B2( u0_u15_u3_n135 ) , .ZN( u0_u15_u3_n136 ) , .C1( u0_u15_u3_n149 ) , .B1( u0_u15_u3_n151 ) , .C2( u0_u15_u3_n183 ) );
  NAND4_X1 u0_u15_u3_U89 (.ZN( u0_out15_26 ) , .A4( u0_u15_u3_n109 ) , .A3( u0_u15_u3_n110 ) , .A2( u0_u15_u3_n111 ) , .A1( u0_u15_u3_n173 ) );
  INV_X1 u0_u15_u3_U9 (.A( u0_u15_u3_n143 ) , .ZN( u0_u15_u3_n168 ) );
  INV_X1 u0_u15_u3_U90 (.ZN( u0_u15_u3_n173 ) , .A( u0_u15_u3_n94 ) );
  OAI21_X1 u0_u15_u3_U91 (.ZN( u0_u15_u3_n111 ) , .B2( u0_u15_u3_n117 ) , .A( u0_u15_u3_n133 ) , .B1( u0_u15_u3_n176 ) );
  NAND4_X1 u0_u15_u3_U92 (.ZN( u0_out15_20 ) , .A4( u0_u15_u3_n122 ) , .A3( u0_u15_u3_n123 ) , .A1( u0_u15_u3_n175 ) , .A2( u0_u15_u3_n180 ) );
  INV_X1 u0_u15_u3_U93 (.A( u0_u15_u3_n126 ) , .ZN( u0_u15_u3_n180 ) );
  INV_X1 u0_u15_u3_U94 (.A( u0_u15_u3_n112 ) , .ZN( u0_u15_u3_n175 ) );
  NAND4_X1 u0_u15_u3_U95 (.ZN( u0_out15_1 ) , .A4( u0_u15_u3_n161 ) , .A3( u0_u15_u3_n162 ) , .A2( u0_u15_u3_n163 ) , .A1( u0_u15_u3_n185 ) );
  NAND2_X1 u0_u15_u3_U96 (.ZN( u0_u15_u3_n163 ) , .A2( u0_u15_u3_n170 ) , .A1( u0_u15_u3_n176 ) );
  AOI22_X1 u0_u15_u3_U97 (.B2( u0_u15_u3_n140 ) , .B1( u0_u15_u3_n141 ) , .A2( u0_u15_u3_n142 ) , .ZN( u0_u15_u3_n162 ) , .A1( u0_u15_u3_n177 ) );
  NAND3_X1 u0_u15_u3_U98 (.A1( u0_u15_u3_n114 ) , .ZN( u0_u15_u3_n115 ) , .A2( u0_u15_u3_n145 ) , .A3( u0_u15_u3_n153 ) );
  NAND3_X1 u0_u15_u3_U99 (.ZN( u0_u15_u3_n129 ) , .A2( u0_u15_u3_n144 ) , .A1( u0_u15_u3_n153 ) , .A3( u0_u15_u3_n182 ) );
  XOR2_X1 u0_u1_U2 (.B( u0_K2_8 ) , .A( u0_R0_5 ) , .Z( u0_u1_X_8 ) );
  XOR2_X1 u0_u1_U3 (.B( u0_K2_7 ) , .A( u0_R0_4 ) , .Z( u0_u1_X_7 ) );
  XOR2_X1 u0_u1_U4 (.B( u0_K2_6 ) , .A( u0_R0_5 ) , .Z( u0_u1_X_6 ) );
  XOR2_X1 u0_u1_U5 (.B( u0_K2_5 ) , .A( u0_R0_4 ) , .Z( u0_u1_X_5 ) );
  AND3_X1 u0_u1_u0_U10 (.A2( u0_u1_u0_n112 ) , .ZN( u0_u1_u0_n127 ) , .A3( u0_u1_u0_n130 ) , .A1( u0_u1_u0_n148 ) );
  NAND2_X1 u0_u1_u0_U11 (.ZN( u0_u1_u0_n113 ) , .A1( u0_u1_u0_n139 ) , .A2( u0_u1_u0_n149 ) );
  AND2_X1 u0_u1_u0_U12 (.ZN( u0_u1_u0_n107 ) , .A1( u0_u1_u0_n130 ) , .A2( u0_u1_u0_n140 ) );
  AND2_X1 u0_u1_u0_U13 (.A2( u0_u1_u0_n129 ) , .A1( u0_u1_u0_n130 ) , .ZN( u0_u1_u0_n151 ) );
  AND2_X1 u0_u1_u0_U14 (.A1( u0_u1_u0_n108 ) , .A2( u0_u1_u0_n125 ) , .ZN( u0_u1_u0_n145 ) );
  INV_X1 u0_u1_u0_U15 (.A( u0_u1_u0_n143 ) , .ZN( u0_u1_u0_n173 ) );
  NOR2_X1 u0_u1_u0_U16 (.A2( u0_u1_u0_n136 ) , .ZN( u0_u1_u0_n147 ) , .A1( u0_u1_u0_n160 ) );
  NOR2_X1 u0_u1_u0_U17 (.A1( u0_u1_u0_n163 ) , .A2( u0_u1_u0_n164 ) , .ZN( u0_u1_u0_n95 ) );
  AOI21_X1 u0_u1_u0_U18 (.B1( u0_u1_u0_n103 ) , .ZN( u0_u1_u0_n132 ) , .A( u0_u1_u0_n165 ) , .B2( u0_u1_u0_n93 ) );
  INV_X1 u0_u1_u0_U19 (.A( u0_u1_u0_n142 ) , .ZN( u0_u1_u0_n165 ) );
  OAI221_X1 u0_u1_u0_U20 (.C1( u0_u1_u0_n121 ) , .ZN( u0_u1_u0_n122 ) , .B2( u0_u1_u0_n127 ) , .A( u0_u1_u0_n143 ) , .B1( u0_u1_u0_n144 ) , .C2( u0_u1_u0_n147 ) );
  OAI22_X1 u0_u1_u0_U21 (.B1( u0_u1_u0_n125 ) , .ZN( u0_u1_u0_n126 ) , .A1( u0_u1_u0_n138 ) , .A2( u0_u1_u0_n146 ) , .B2( u0_u1_u0_n147 ) );
  OAI22_X1 u0_u1_u0_U22 (.B1( u0_u1_u0_n131 ) , .A1( u0_u1_u0_n144 ) , .B2( u0_u1_u0_n147 ) , .A2( u0_u1_u0_n90 ) , .ZN( u0_u1_u0_n91 ) );
  AND3_X1 u0_u1_u0_U23 (.A3( u0_u1_u0_n121 ) , .A2( u0_u1_u0_n125 ) , .A1( u0_u1_u0_n148 ) , .ZN( u0_u1_u0_n90 ) );
  INV_X1 u0_u1_u0_U24 (.A( u0_u1_u0_n136 ) , .ZN( u0_u1_u0_n161 ) );
  NOR2_X1 u0_u1_u0_U25 (.A1( u0_u1_u0_n120 ) , .ZN( u0_u1_u0_n143 ) , .A2( u0_u1_u0_n167 ) );
  OAI221_X1 u0_u1_u0_U26 (.C1( u0_u1_u0_n112 ) , .ZN( u0_u1_u0_n120 ) , .B1( u0_u1_u0_n138 ) , .B2( u0_u1_u0_n141 ) , .C2( u0_u1_u0_n147 ) , .A( u0_u1_u0_n172 ) );
  AOI211_X1 u0_u1_u0_U27 (.B( u0_u1_u0_n115 ) , .A( u0_u1_u0_n116 ) , .C2( u0_u1_u0_n117 ) , .C1( u0_u1_u0_n118 ) , .ZN( u0_u1_u0_n119 ) );
  AOI22_X1 u0_u1_u0_U28 (.B2( u0_u1_u0_n109 ) , .A2( u0_u1_u0_n110 ) , .ZN( u0_u1_u0_n111 ) , .B1( u0_u1_u0_n118 ) , .A1( u0_u1_u0_n160 ) );
  INV_X1 u0_u1_u0_U29 (.A( u0_u1_u0_n118 ) , .ZN( u0_u1_u0_n158 ) );
  INV_X1 u0_u1_u0_U3 (.A( u0_u1_u0_n113 ) , .ZN( u0_u1_u0_n166 ) );
  AOI21_X1 u0_u1_u0_U30 (.ZN( u0_u1_u0_n104 ) , .B1( u0_u1_u0_n107 ) , .B2( u0_u1_u0_n141 ) , .A( u0_u1_u0_n144 ) );
  AOI21_X1 u0_u1_u0_U31 (.B1( u0_u1_u0_n127 ) , .B2( u0_u1_u0_n129 ) , .A( u0_u1_u0_n138 ) , .ZN( u0_u1_u0_n96 ) );
  AOI21_X1 u0_u1_u0_U32 (.ZN( u0_u1_u0_n116 ) , .B2( u0_u1_u0_n142 ) , .A( u0_u1_u0_n144 ) , .B1( u0_u1_u0_n166 ) );
  NAND2_X1 u0_u1_u0_U33 (.A1( u0_u1_u0_n100 ) , .A2( u0_u1_u0_n103 ) , .ZN( u0_u1_u0_n125 ) );
  NAND2_X1 u0_u1_u0_U34 (.A2( u0_u1_u0_n103 ) , .ZN( u0_u1_u0_n140 ) , .A1( u0_u1_u0_n94 ) );
  NAND2_X1 u0_u1_u0_U35 (.A1( u0_u1_u0_n101 ) , .A2( u0_u1_u0_n102 ) , .ZN( u0_u1_u0_n150 ) );
  INV_X1 u0_u1_u0_U36 (.A( u0_u1_u0_n138 ) , .ZN( u0_u1_u0_n160 ) );
  NAND2_X1 u0_u1_u0_U37 (.ZN( u0_u1_u0_n142 ) , .A1( u0_u1_u0_n94 ) , .A2( u0_u1_u0_n95 ) );
  NAND2_X1 u0_u1_u0_U38 (.A1( u0_u1_u0_n102 ) , .ZN( u0_u1_u0_n128 ) , .A2( u0_u1_u0_n95 ) );
  NAND2_X1 u0_u1_u0_U39 (.A2( u0_u1_u0_n102 ) , .A1( u0_u1_u0_n103 ) , .ZN( u0_u1_u0_n149 ) );
  AOI21_X1 u0_u1_u0_U4 (.B1( u0_u1_u0_n114 ) , .ZN( u0_u1_u0_n115 ) , .B2( u0_u1_u0_n129 ) , .A( u0_u1_u0_n161 ) );
  NAND2_X1 u0_u1_u0_U40 (.A1( u0_u1_u0_n100 ) , .ZN( u0_u1_u0_n129 ) , .A2( u0_u1_u0_n95 ) );
  NAND2_X1 u0_u1_u0_U41 (.A2( u0_u1_u0_n100 ) , .A1( u0_u1_u0_n101 ) , .ZN( u0_u1_u0_n139 ) );
  NAND2_X1 u0_u1_u0_U42 (.A2( u0_u1_u0_n100 ) , .ZN( u0_u1_u0_n131 ) , .A1( u0_u1_u0_n92 ) );
  NAND2_X1 u0_u1_u0_U43 (.ZN( u0_u1_u0_n108 ) , .A1( u0_u1_u0_n92 ) , .A2( u0_u1_u0_n94 ) );
  NAND2_X1 u0_u1_u0_U44 (.ZN( u0_u1_u0_n148 ) , .A1( u0_u1_u0_n93 ) , .A2( u0_u1_u0_n95 ) );
  NAND2_X1 u0_u1_u0_U45 (.A2( u0_u1_u0_n102 ) , .ZN( u0_u1_u0_n114 ) , .A1( u0_u1_u0_n92 ) );
  NAND2_X1 u0_u1_u0_U46 (.A1( u0_u1_u0_n101 ) , .ZN( u0_u1_u0_n130 ) , .A2( u0_u1_u0_n94 ) );
  NAND2_X1 u0_u1_u0_U47 (.A2( u0_u1_u0_n101 ) , .ZN( u0_u1_u0_n121 ) , .A1( u0_u1_u0_n93 ) );
  INV_X1 u0_u1_u0_U48 (.ZN( u0_u1_u0_n172 ) , .A( u0_u1_u0_n88 ) );
  OAI222_X1 u0_u1_u0_U49 (.C1( u0_u1_u0_n108 ) , .A1( u0_u1_u0_n125 ) , .B2( u0_u1_u0_n128 ) , .B1( u0_u1_u0_n144 ) , .A2( u0_u1_u0_n158 ) , .C2( u0_u1_u0_n161 ) , .ZN( u0_u1_u0_n88 ) );
  AOI21_X1 u0_u1_u0_U5 (.B2( u0_u1_u0_n131 ) , .ZN( u0_u1_u0_n134 ) , .B1( u0_u1_u0_n151 ) , .A( u0_u1_u0_n158 ) );
  NAND2_X1 u0_u1_u0_U50 (.ZN( u0_u1_u0_n112 ) , .A2( u0_u1_u0_n92 ) , .A1( u0_u1_u0_n93 ) );
  OR3_X1 u0_u1_u0_U51 (.A3( u0_u1_u0_n152 ) , .A2( u0_u1_u0_n153 ) , .A1( u0_u1_u0_n154 ) , .ZN( u0_u1_u0_n155 ) );
  AOI21_X1 u0_u1_u0_U52 (.B2( u0_u1_u0_n150 ) , .B1( u0_u1_u0_n151 ) , .ZN( u0_u1_u0_n152 ) , .A( u0_u1_u0_n158 ) );
  AOI21_X1 u0_u1_u0_U53 (.A( u0_u1_u0_n144 ) , .B2( u0_u1_u0_n145 ) , .B1( u0_u1_u0_n146 ) , .ZN( u0_u1_u0_n154 ) );
  AOI21_X1 u0_u1_u0_U54 (.A( u0_u1_u0_n147 ) , .B2( u0_u1_u0_n148 ) , .B1( u0_u1_u0_n149 ) , .ZN( u0_u1_u0_n153 ) );
  INV_X1 u0_u1_u0_U55 (.ZN( u0_u1_u0_n171 ) , .A( u0_u1_u0_n99 ) );
  OAI211_X1 u0_u1_u0_U56 (.C2( u0_u1_u0_n140 ) , .C1( u0_u1_u0_n161 ) , .A( u0_u1_u0_n169 ) , .B( u0_u1_u0_n98 ) , .ZN( u0_u1_u0_n99 ) );
  INV_X1 u0_u1_u0_U57 (.ZN( u0_u1_u0_n169 ) , .A( u0_u1_u0_n91 ) );
  AOI211_X1 u0_u1_u0_U58 (.C1( u0_u1_u0_n118 ) , .A( u0_u1_u0_n123 ) , .B( u0_u1_u0_n96 ) , .C2( u0_u1_u0_n97 ) , .ZN( u0_u1_u0_n98 ) );
  NOR2_X1 u0_u1_u0_U59 (.A2( u0_u1_X_2 ) , .ZN( u0_u1_u0_n103 ) , .A1( u0_u1_u0_n164 ) );
  NOR2_X1 u0_u1_u0_U6 (.A1( u0_u1_u0_n108 ) , .ZN( u0_u1_u0_n123 ) , .A2( u0_u1_u0_n158 ) );
  NOR2_X1 u0_u1_u0_U60 (.A2( u0_u1_X_3 ) , .A1( u0_u1_X_6 ) , .ZN( u0_u1_u0_n94 ) );
  NOR2_X1 u0_u1_u0_U61 (.A2( u0_u1_X_6 ) , .ZN( u0_u1_u0_n100 ) , .A1( u0_u1_u0_n162 ) );
  NOR2_X1 u0_u1_u0_U62 (.A2( u0_u1_X_4 ) , .A1( u0_u1_X_5 ) , .ZN( u0_u1_u0_n118 ) );
  NOR2_X1 u0_u1_u0_U63 (.A2( u0_u1_X_1 ) , .A1( u0_u1_X_2 ) , .ZN( u0_u1_u0_n92 ) );
  NOR2_X1 u0_u1_u0_U64 (.A2( u0_u1_X_1 ) , .ZN( u0_u1_u0_n101 ) , .A1( u0_u1_u0_n163 ) );
  NAND2_X1 u0_u1_u0_U65 (.A2( u0_u1_X_4 ) , .A1( u0_u1_X_5 ) , .ZN( u0_u1_u0_n144 ) );
  NOR2_X1 u0_u1_u0_U66 (.A2( u0_u1_X_5 ) , .ZN( u0_u1_u0_n136 ) , .A1( u0_u1_u0_n159 ) );
  NAND2_X1 u0_u1_u0_U67 (.A1( u0_u1_X_5 ) , .ZN( u0_u1_u0_n138 ) , .A2( u0_u1_u0_n159 ) );
  AND2_X1 u0_u1_u0_U68 (.A2( u0_u1_X_3 ) , .A1( u0_u1_X_6 ) , .ZN( u0_u1_u0_n102 ) );
  AND2_X1 u0_u1_u0_U69 (.A1( u0_u1_X_6 ) , .A2( u0_u1_u0_n162 ) , .ZN( u0_u1_u0_n93 ) );
  OAI21_X1 u0_u1_u0_U7 (.B1( u0_u1_u0_n150 ) , .B2( u0_u1_u0_n158 ) , .A( u0_u1_u0_n172 ) , .ZN( u0_u1_u0_n89 ) );
  INV_X1 u0_u1_u0_U70 (.A( u0_u1_X_4 ) , .ZN( u0_u1_u0_n159 ) );
  INV_X1 u0_u1_u0_U71 (.A( u0_u1_X_1 ) , .ZN( u0_u1_u0_n164 ) );
  INV_X1 u0_u1_u0_U72 (.A( u0_u1_X_2 ) , .ZN( u0_u1_u0_n163 ) );
  INV_X1 u0_u1_u0_U73 (.A( u0_u1_X_3 ) , .ZN( u0_u1_u0_n162 ) );
  INV_X1 u0_u1_u0_U74 (.ZN( u0_u1_u0_n174 ) , .A( u0_u1_u0_n89 ) );
  AOI211_X1 u0_u1_u0_U75 (.B( u0_u1_u0_n104 ) , .A( u0_u1_u0_n105 ) , .ZN( u0_u1_u0_n106 ) , .C2( u0_u1_u0_n113 ) , .C1( u0_u1_u0_n160 ) );
  INV_X1 u0_u1_u0_U76 (.A( u0_u1_u0_n126 ) , .ZN( u0_u1_u0_n168 ) );
  AOI211_X1 u0_u1_u0_U77 (.B( u0_u1_u0_n133 ) , .A( u0_u1_u0_n134 ) , .C2( u0_u1_u0_n135 ) , .C1( u0_u1_u0_n136 ) , .ZN( u0_u1_u0_n137 ) );
  OR4_X1 u0_u1_u0_U78 (.ZN( u0_out1_31 ) , .A4( u0_u1_u0_n155 ) , .A2( u0_u1_u0_n156 ) , .A1( u0_u1_u0_n157 ) , .A3( u0_u1_u0_n173 ) );
  AOI21_X1 u0_u1_u0_U79 (.A( u0_u1_u0_n138 ) , .B2( u0_u1_u0_n139 ) , .B1( u0_u1_u0_n140 ) , .ZN( u0_u1_u0_n157 ) );
  AND2_X1 u0_u1_u0_U8 (.A1( u0_u1_u0_n114 ) , .A2( u0_u1_u0_n121 ) , .ZN( u0_u1_u0_n146 ) );
  AOI21_X1 u0_u1_u0_U80 (.B2( u0_u1_u0_n141 ) , .B1( u0_u1_u0_n142 ) , .ZN( u0_u1_u0_n156 ) , .A( u0_u1_u0_n161 ) );
  OR4_X1 u0_u1_u0_U81 (.ZN( u0_out1_17 ) , .A4( u0_u1_u0_n122 ) , .A2( u0_u1_u0_n123 ) , .A1( u0_u1_u0_n124 ) , .A3( u0_u1_u0_n170 ) );
  AOI21_X1 u0_u1_u0_U82 (.B2( u0_u1_u0_n107 ) , .ZN( u0_u1_u0_n124 ) , .B1( u0_u1_u0_n128 ) , .A( u0_u1_u0_n161 ) );
  INV_X1 u0_u1_u0_U83 (.A( u0_u1_u0_n111 ) , .ZN( u0_u1_u0_n170 ) );
  AOI21_X1 u0_u1_u0_U84 (.B1( u0_u1_u0_n132 ) , .ZN( u0_u1_u0_n133 ) , .A( u0_u1_u0_n144 ) , .B2( u0_u1_u0_n166 ) );
  OAI22_X1 u0_u1_u0_U85 (.ZN( u0_u1_u0_n105 ) , .A2( u0_u1_u0_n132 ) , .B1( u0_u1_u0_n146 ) , .A1( u0_u1_u0_n147 ) , .B2( u0_u1_u0_n161 ) );
  NAND2_X1 u0_u1_u0_U86 (.ZN( u0_u1_u0_n110 ) , .A2( u0_u1_u0_n132 ) , .A1( u0_u1_u0_n145 ) );
  INV_X1 u0_u1_u0_U87 (.A( u0_u1_u0_n119 ) , .ZN( u0_u1_u0_n167 ) );
  NAND3_X1 u0_u1_u0_U88 (.ZN( u0_out1_23 ) , .A3( u0_u1_u0_n137 ) , .A1( u0_u1_u0_n168 ) , .A2( u0_u1_u0_n171 ) );
  NAND3_X1 u0_u1_u0_U89 (.A3( u0_u1_u0_n127 ) , .A2( u0_u1_u0_n128 ) , .ZN( u0_u1_u0_n135 ) , .A1( u0_u1_u0_n150 ) );
  AND2_X1 u0_u1_u0_U9 (.A1( u0_u1_u0_n131 ) , .ZN( u0_u1_u0_n141 ) , .A2( u0_u1_u0_n150 ) );
  NAND3_X1 u0_u1_u0_U90 (.ZN( u0_u1_u0_n117 ) , .A3( u0_u1_u0_n132 ) , .A2( u0_u1_u0_n139 ) , .A1( u0_u1_u0_n148 ) );
  NAND3_X1 u0_u1_u0_U91 (.ZN( u0_u1_u0_n109 ) , .A2( u0_u1_u0_n114 ) , .A3( u0_u1_u0_n140 ) , .A1( u0_u1_u0_n149 ) );
  NAND3_X1 u0_u1_u0_U92 (.ZN( u0_out1_9 ) , .A3( u0_u1_u0_n106 ) , .A2( u0_u1_u0_n171 ) , .A1( u0_u1_u0_n174 ) );
  NAND3_X1 u0_u1_u0_U93 (.A2( u0_u1_u0_n128 ) , .A1( u0_u1_u0_n132 ) , .A3( u0_u1_u0_n146 ) , .ZN( u0_u1_u0_n97 ) );
  NOR2_X1 u0_u1_u1_U10 (.A1( u0_u1_u1_n112 ) , .A2( u0_u1_u1_n116 ) , .ZN( u0_u1_u1_n118 ) );
  NAND3_X1 u0_u1_u1_U100 (.ZN( u0_u1_u1_n113 ) , .A1( u0_u1_u1_n120 ) , .A3( u0_u1_u1_n133 ) , .A2( u0_u1_u1_n155 ) );
  OAI21_X1 u0_u1_u1_U11 (.ZN( u0_u1_u1_n101 ) , .B1( u0_u1_u1_n141 ) , .A( u0_u1_u1_n146 ) , .B2( u0_u1_u1_n183 ) );
  AOI21_X1 u0_u1_u1_U12 (.B2( u0_u1_u1_n155 ) , .B1( u0_u1_u1_n156 ) , .ZN( u0_u1_u1_n157 ) , .A( u0_u1_u1_n174 ) );
  OR4_X1 u0_u1_u1_U13 (.A4( u0_u1_u1_n106 ) , .A3( u0_u1_u1_n107 ) , .ZN( u0_u1_u1_n108 ) , .A1( u0_u1_u1_n117 ) , .A2( u0_u1_u1_n184 ) );
  AOI21_X1 u0_u1_u1_U14 (.ZN( u0_u1_u1_n106 ) , .A( u0_u1_u1_n112 ) , .B1( u0_u1_u1_n154 ) , .B2( u0_u1_u1_n156 ) );
  INV_X1 u0_u1_u1_U15 (.A( u0_u1_u1_n101 ) , .ZN( u0_u1_u1_n184 ) );
  AOI21_X1 u0_u1_u1_U16 (.ZN( u0_u1_u1_n107 ) , .B1( u0_u1_u1_n134 ) , .B2( u0_u1_u1_n149 ) , .A( u0_u1_u1_n174 ) );
  NAND2_X1 u0_u1_u1_U17 (.ZN( u0_u1_u1_n140 ) , .A2( u0_u1_u1_n150 ) , .A1( u0_u1_u1_n155 ) );
  NAND2_X1 u0_u1_u1_U18 (.A1( u0_u1_u1_n131 ) , .ZN( u0_u1_u1_n147 ) , .A2( u0_u1_u1_n153 ) );
  INV_X1 u0_u1_u1_U19 (.A( u0_u1_u1_n139 ) , .ZN( u0_u1_u1_n174 ) );
  INV_X1 u0_u1_u1_U20 (.A( u0_u1_u1_n112 ) , .ZN( u0_u1_u1_n171 ) );
  NAND2_X1 u0_u1_u1_U21 (.ZN( u0_u1_u1_n141 ) , .A1( u0_u1_u1_n153 ) , .A2( u0_u1_u1_n156 ) );
  AND2_X1 u0_u1_u1_U22 (.A1( u0_u1_u1_n123 ) , .ZN( u0_u1_u1_n134 ) , .A2( u0_u1_u1_n161 ) );
  NAND2_X1 u0_u1_u1_U23 (.A2( u0_u1_u1_n115 ) , .A1( u0_u1_u1_n116 ) , .ZN( u0_u1_u1_n148 ) );
  NAND2_X1 u0_u1_u1_U24 (.A2( u0_u1_u1_n133 ) , .A1( u0_u1_u1_n135 ) , .ZN( u0_u1_u1_n159 ) );
  NAND2_X1 u0_u1_u1_U25 (.A2( u0_u1_u1_n115 ) , .A1( u0_u1_u1_n120 ) , .ZN( u0_u1_u1_n132 ) );
  INV_X1 u0_u1_u1_U26 (.A( u0_u1_u1_n154 ) , .ZN( u0_u1_u1_n178 ) );
  INV_X1 u0_u1_u1_U27 (.A( u0_u1_u1_n151 ) , .ZN( u0_u1_u1_n183 ) );
  AND2_X1 u0_u1_u1_U28 (.A1( u0_u1_u1_n129 ) , .A2( u0_u1_u1_n133 ) , .ZN( u0_u1_u1_n149 ) );
  INV_X1 u0_u1_u1_U29 (.A( u0_u1_u1_n131 ) , .ZN( u0_u1_u1_n180 ) );
  INV_X1 u0_u1_u1_U3 (.A( u0_u1_u1_n159 ) , .ZN( u0_u1_u1_n182 ) );
  AOI221_X1 u0_u1_u1_U30 (.B1( u0_u1_u1_n140 ) , .ZN( u0_u1_u1_n167 ) , .B2( u0_u1_u1_n172 ) , .C2( u0_u1_u1_n175 ) , .C1( u0_u1_u1_n178 ) , .A( u0_u1_u1_n188 ) );
  INV_X1 u0_u1_u1_U31 (.ZN( u0_u1_u1_n188 ) , .A( u0_u1_u1_n97 ) );
  AOI211_X1 u0_u1_u1_U32 (.A( u0_u1_u1_n118 ) , .C1( u0_u1_u1_n132 ) , .C2( u0_u1_u1_n139 ) , .B( u0_u1_u1_n96 ) , .ZN( u0_u1_u1_n97 ) );
  AOI21_X1 u0_u1_u1_U33 (.B2( u0_u1_u1_n121 ) , .B1( u0_u1_u1_n135 ) , .A( u0_u1_u1_n152 ) , .ZN( u0_u1_u1_n96 ) );
  OAI221_X1 u0_u1_u1_U34 (.A( u0_u1_u1_n119 ) , .C2( u0_u1_u1_n129 ) , .ZN( u0_u1_u1_n138 ) , .B2( u0_u1_u1_n152 ) , .C1( u0_u1_u1_n174 ) , .B1( u0_u1_u1_n187 ) );
  INV_X1 u0_u1_u1_U35 (.A( u0_u1_u1_n148 ) , .ZN( u0_u1_u1_n187 ) );
  AOI211_X1 u0_u1_u1_U36 (.B( u0_u1_u1_n117 ) , .A( u0_u1_u1_n118 ) , .ZN( u0_u1_u1_n119 ) , .C2( u0_u1_u1_n146 ) , .C1( u0_u1_u1_n159 ) );
  NOR2_X1 u0_u1_u1_U37 (.A1( u0_u1_u1_n168 ) , .A2( u0_u1_u1_n176 ) , .ZN( u0_u1_u1_n98 ) );
  AOI211_X1 u0_u1_u1_U38 (.B( u0_u1_u1_n162 ) , .A( u0_u1_u1_n163 ) , .C2( u0_u1_u1_n164 ) , .ZN( u0_u1_u1_n165 ) , .C1( u0_u1_u1_n171 ) );
  AOI21_X1 u0_u1_u1_U39 (.A( u0_u1_u1_n160 ) , .B2( u0_u1_u1_n161 ) , .ZN( u0_u1_u1_n162 ) , .B1( u0_u1_u1_n182 ) );
  AOI221_X1 u0_u1_u1_U4 (.A( u0_u1_u1_n138 ) , .C2( u0_u1_u1_n139 ) , .C1( u0_u1_u1_n140 ) , .B2( u0_u1_u1_n141 ) , .ZN( u0_u1_u1_n142 ) , .B1( u0_u1_u1_n175 ) );
  OR2_X1 u0_u1_u1_U40 (.A2( u0_u1_u1_n157 ) , .A1( u0_u1_u1_n158 ) , .ZN( u0_u1_u1_n163 ) );
  OAI21_X1 u0_u1_u1_U41 (.B2( u0_u1_u1_n123 ) , .ZN( u0_u1_u1_n145 ) , .B1( u0_u1_u1_n160 ) , .A( u0_u1_u1_n185 ) );
  INV_X1 u0_u1_u1_U42 (.A( u0_u1_u1_n122 ) , .ZN( u0_u1_u1_n185 ) );
  AOI21_X1 u0_u1_u1_U43 (.B2( u0_u1_u1_n120 ) , .B1( u0_u1_u1_n121 ) , .ZN( u0_u1_u1_n122 ) , .A( u0_u1_u1_n128 ) );
  NAND2_X1 u0_u1_u1_U44 (.A1( u0_u1_u1_n128 ) , .ZN( u0_u1_u1_n146 ) , .A2( u0_u1_u1_n160 ) );
  NAND2_X1 u0_u1_u1_U45 (.A2( u0_u1_u1_n112 ) , .ZN( u0_u1_u1_n139 ) , .A1( u0_u1_u1_n152 ) );
  NAND2_X1 u0_u1_u1_U46 (.A1( u0_u1_u1_n105 ) , .ZN( u0_u1_u1_n156 ) , .A2( u0_u1_u1_n99 ) );
  NOR2_X1 u0_u1_u1_U47 (.ZN( u0_u1_u1_n117 ) , .A1( u0_u1_u1_n121 ) , .A2( u0_u1_u1_n160 ) );
  AOI21_X1 u0_u1_u1_U48 (.A( u0_u1_u1_n128 ) , .B2( u0_u1_u1_n129 ) , .ZN( u0_u1_u1_n130 ) , .B1( u0_u1_u1_n150 ) );
  NAND2_X1 u0_u1_u1_U49 (.ZN( u0_u1_u1_n112 ) , .A1( u0_u1_u1_n169 ) , .A2( u0_u1_u1_n170 ) );
  AOI211_X1 u0_u1_u1_U5 (.ZN( u0_u1_u1_n124 ) , .A( u0_u1_u1_n138 ) , .C2( u0_u1_u1_n139 ) , .B( u0_u1_u1_n145 ) , .C1( u0_u1_u1_n147 ) );
  NAND2_X1 u0_u1_u1_U50 (.ZN( u0_u1_u1_n129 ) , .A2( u0_u1_u1_n95 ) , .A1( u0_u1_u1_n98 ) );
  NAND2_X1 u0_u1_u1_U51 (.A1( u0_u1_u1_n102 ) , .ZN( u0_u1_u1_n154 ) , .A2( u0_u1_u1_n99 ) );
  NAND2_X1 u0_u1_u1_U52 (.A2( u0_u1_u1_n100 ) , .ZN( u0_u1_u1_n135 ) , .A1( u0_u1_u1_n99 ) );
  AOI21_X1 u0_u1_u1_U53 (.A( u0_u1_u1_n152 ) , .B2( u0_u1_u1_n153 ) , .B1( u0_u1_u1_n154 ) , .ZN( u0_u1_u1_n158 ) );
  INV_X1 u0_u1_u1_U54 (.A( u0_u1_u1_n160 ) , .ZN( u0_u1_u1_n175 ) );
  NAND2_X1 u0_u1_u1_U55 (.A1( u0_u1_u1_n100 ) , .ZN( u0_u1_u1_n116 ) , .A2( u0_u1_u1_n95 ) );
  NAND2_X1 u0_u1_u1_U56 (.A1( u0_u1_u1_n102 ) , .ZN( u0_u1_u1_n131 ) , .A2( u0_u1_u1_n95 ) );
  NAND2_X1 u0_u1_u1_U57 (.A2( u0_u1_u1_n104 ) , .ZN( u0_u1_u1_n121 ) , .A1( u0_u1_u1_n98 ) );
  NAND2_X1 u0_u1_u1_U58 (.A1( u0_u1_u1_n103 ) , .ZN( u0_u1_u1_n153 ) , .A2( u0_u1_u1_n98 ) );
  NAND2_X1 u0_u1_u1_U59 (.A2( u0_u1_u1_n104 ) , .A1( u0_u1_u1_n105 ) , .ZN( u0_u1_u1_n133 ) );
  AOI22_X1 u0_u1_u1_U6 (.B2( u0_u1_u1_n113 ) , .A2( u0_u1_u1_n114 ) , .ZN( u0_u1_u1_n125 ) , .A1( u0_u1_u1_n171 ) , .B1( u0_u1_u1_n173 ) );
  NAND2_X1 u0_u1_u1_U60 (.ZN( u0_u1_u1_n150 ) , .A2( u0_u1_u1_n98 ) , .A1( u0_u1_u1_n99 ) );
  NAND2_X1 u0_u1_u1_U61 (.A1( u0_u1_u1_n105 ) , .ZN( u0_u1_u1_n155 ) , .A2( u0_u1_u1_n95 ) );
  OAI21_X1 u0_u1_u1_U62 (.ZN( u0_u1_u1_n109 ) , .B1( u0_u1_u1_n129 ) , .B2( u0_u1_u1_n160 ) , .A( u0_u1_u1_n167 ) );
  NAND2_X1 u0_u1_u1_U63 (.A2( u0_u1_u1_n100 ) , .A1( u0_u1_u1_n103 ) , .ZN( u0_u1_u1_n120 ) );
  NAND2_X1 u0_u1_u1_U64 (.A1( u0_u1_u1_n102 ) , .A2( u0_u1_u1_n104 ) , .ZN( u0_u1_u1_n115 ) );
  NAND2_X1 u0_u1_u1_U65 (.A2( u0_u1_u1_n100 ) , .A1( u0_u1_u1_n104 ) , .ZN( u0_u1_u1_n151 ) );
  NAND2_X1 u0_u1_u1_U66 (.A2( u0_u1_u1_n103 ) , .A1( u0_u1_u1_n105 ) , .ZN( u0_u1_u1_n161 ) );
  INV_X1 u0_u1_u1_U67 (.A( u0_u1_u1_n152 ) , .ZN( u0_u1_u1_n173 ) );
  INV_X1 u0_u1_u1_U68 (.A( u0_u1_u1_n128 ) , .ZN( u0_u1_u1_n172 ) );
  NAND2_X1 u0_u1_u1_U69 (.A2( u0_u1_u1_n102 ) , .A1( u0_u1_u1_n103 ) , .ZN( u0_u1_u1_n123 ) );
  NAND2_X1 u0_u1_u1_U7 (.ZN( u0_u1_u1_n114 ) , .A1( u0_u1_u1_n134 ) , .A2( u0_u1_u1_n156 ) );
  NOR2_X1 u0_u1_u1_U70 (.A2( u0_u1_X_7 ) , .A1( u0_u1_X_8 ) , .ZN( u0_u1_u1_n95 ) );
  NOR2_X1 u0_u1_u1_U71 (.A1( u0_u1_X_12 ) , .A2( u0_u1_X_9 ) , .ZN( u0_u1_u1_n100 ) );
  NOR2_X1 u0_u1_u1_U72 (.A2( u0_u1_X_8 ) , .A1( u0_u1_u1_n177 ) , .ZN( u0_u1_u1_n99 ) );
  NOR2_X1 u0_u1_u1_U73 (.A2( u0_u1_X_12 ) , .ZN( u0_u1_u1_n102 ) , .A1( u0_u1_u1_n176 ) );
  NOR2_X1 u0_u1_u1_U74 (.A2( u0_u1_X_9 ) , .ZN( u0_u1_u1_n105 ) , .A1( u0_u1_u1_n168 ) );
  NAND2_X1 u0_u1_u1_U75 (.A1( u0_u1_X_10 ) , .ZN( u0_u1_u1_n160 ) , .A2( u0_u1_u1_n169 ) );
  NAND2_X1 u0_u1_u1_U76 (.A2( u0_u1_X_10 ) , .A1( u0_u1_X_11 ) , .ZN( u0_u1_u1_n152 ) );
  NAND2_X1 u0_u1_u1_U77 (.A1( u0_u1_X_11 ) , .ZN( u0_u1_u1_n128 ) , .A2( u0_u1_u1_n170 ) );
  AND2_X1 u0_u1_u1_U78 (.A2( u0_u1_X_7 ) , .A1( u0_u1_X_8 ) , .ZN( u0_u1_u1_n104 ) );
  AND2_X1 u0_u1_u1_U79 (.A1( u0_u1_X_8 ) , .ZN( u0_u1_u1_n103 ) , .A2( u0_u1_u1_n177 ) );
  AOI22_X1 u0_u1_u1_U8 (.B2( u0_u1_u1_n136 ) , .A2( u0_u1_u1_n137 ) , .ZN( u0_u1_u1_n143 ) , .A1( u0_u1_u1_n171 ) , .B1( u0_u1_u1_n173 ) );
  INV_X1 u0_u1_u1_U80 (.A( u0_u1_X_10 ) , .ZN( u0_u1_u1_n170 ) );
  INV_X1 u0_u1_u1_U81 (.A( u0_u1_X_9 ) , .ZN( u0_u1_u1_n176 ) );
  INV_X1 u0_u1_u1_U82 (.A( u0_u1_X_11 ) , .ZN( u0_u1_u1_n169 ) );
  INV_X1 u0_u1_u1_U83 (.A( u0_u1_X_12 ) , .ZN( u0_u1_u1_n168 ) );
  INV_X1 u0_u1_u1_U84 (.A( u0_u1_X_7 ) , .ZN( u0_u1_u1_n177 ) );
  NAND4_X1 u0_u1_u1_U85 (.ZN( u0_out1_28 ) , .A4( u0_u1_u1_n124 ) , .A3( u0_u1_u1_n125 ) , .A2( u0_u1_u1_n126 ) , .A1( u0_u1_u1_n127 ) );
  OAI21_X1 u0_u1_u1_U86 (.ZN( u0_u1_u1_n127 ) , .B2( u0_u1_u1_n139 ) , .B1( u0_u1_u1_n175 ) , .A( u0_u1_u1_n183 ) );
  OAI21_X1 u0_u1_u1_U87 (.ZN( u0_u1_u1_n126 ) , .B2( u0_u1_u1_n140 ) , .A( u0_u1_u1_n146 ) , .B1( u0_u1_u1_n178 ) );
  NAND4_X1 u0_u1_u1_U88 (.ZN( u0_out1_18 ) , .A4( u0_u1_u1_n165 ) , .A3( u0_u1_u1_n166 ) , .A1( u0_u1_u1_n167 ) , .A2( u0_u1_u1_n186 ) );
  AOI22_X1 u0_u1_u1_U89 (.B2( u0_u1_u1_n146 ) , .B1( u0_u1_u1_n147 ) , .A2( u0_u1_u1_n148 ) , .ZN( u0_u1_u1_n166 ) , .A1( u0_u1_u1_n172 ) );
  INV_X1 u0_u1_u1_U9 (.A( u0_u1_u1_n147 ) , .ZN( u0_u1_u1_n181 ) );
  INV_X1 u0_u1_u1_U90 (.A( u0_u1_u1_n145 ) , .ZN( u0_u1_u1_n186 ) );
  NAND4_X1 u0_u1_u1_U91 (.ZN( u0_out1_2 ) , .A4( u0_u1_u1_n142 ) , .A3( u0_u1_u1_n143 ) , .A2( u0_u1_u1_n144 ) , .A1( u0_u1_u1_n179 ) );
  INV_X1 u0_u1_u1_U92 (.A( u0_u1_u1_n130 ) , .ZN( u0_u1_u1_n179 ) );
  OAI21_X1 u0_u1_u1_U93 (.B2( u0_u1_u1_n132 ) , .ZN( u0_u1_u1_n144 ) , .A( u0_u1_u1_n146 ) , .B1( u0_u1_u1_n180 ) );
  OR4_X1 u0_u1_u1_U94 (.ZN( u0_out1_13 ) , .A4( u0_u1_u1_n108 ) , .A3( u0_u1_u1_n109 ) , .A2( u0_u1_u1_n110 ) , .A1( u0_u1_u1_n111 ) );
  AOI21_X1 u0_u1_u1_U95 (.ZN( u0_u1_u1_n111 ) , .A( u0_u1_u1_n128 ) , .B2( u0_u1_u1_n131 ) , .B1( u0_u1_u1_n135 ) );
  AOI21_X1 u0_u1_u1_U96 (.ZN( u0_u1_u1_n110 ) , .A( u0_u1_u1_n116 ) , .B1( u0_u1_u1_n152 ) , .B2( u0_u1_u1_n160 ) );
  NAND3_X1 u0_u1_u1_U97 (.A3( u0_u1_u1_n149 ) , .A2( u0_u1_u1_n150 ) , .A1( u0_u1_u1_n151 ) , .ZN( u0_u1_u1_n164 ) );
  NAND3_X1 u0_u1_u1_U98 (.A3( u0_u1_u1_n134 ) , .A2( u0_u1_u1_n135 ) , .ZN( u0_u1_u1_n136 ) , .A1( u0_u1_u1_n151 ) );
  NAND3_X1 u0_u1_u1_U99 (.A1( u0_u1_u1_n133 ) , .ZN( u0_u1_u1_n137 ) , .A2( u0_u1_u1_n154 ) , .A3( u0_u1_u1_n181 ) );
  XOR2_X1 u0_u3_U1 (.B( u0_K4_9 ) , .A( u0_R2_6 ) , .Z( u0_u3_X_9 ) );
  XOR2_X1 u0_u3_U27 (.B( u0_K4_2 ) , .A( u0_R2_1 ) , .Z( u0_u3_X_2 ) );
  XOR2_X1 u0_u3_U3 (.B( u0_K4_7 ) , .A( u0_R2_4 ) , .Z( u0_u3_X_7 ) );
  XOR2_X1 u0_u3_U38 (.B( u0_K4_1 ) , .A( u0_R2_32 ) , .Z( u0_u3_X_1 ) );
  XOR2_X1 u0_u3_U40 (.B( u0_K4_18 ) , .A( u0_R2_13 ) , .Z( u0_u3_X_18 ) );
  XOR2_X1 u0_u3_U41 (.B( u0_K4_17 ) , .A( u0_R2_12 ) , .Z( u0_u3_X_17 ) );
  XOR2_X1 u0_u3_U42 (.B( u0_K4_16 ) , .A( u0_R2_11 ) , .Z( u0_u3_X_16 ) );
  XOR2_X1 u0_u3_U43 (.B( u0_K4_15 ) , .A( u0_R2_10 ) , .Z( u0_u3_X_15 ) );
  XOR2_X1 u0_u3_U44 (.B( u0_K4_14 ) , .A( u0_R2_9 ) , .Z( u0_u3_X_14 ) );
  XOR2_X1 u0_u3_U45 (.B( u0_K4_13 ) , .A( u0_R2_8 ) , .Z( u0_u3_X_13 ) );
  XOR2_X1 u0_u3_U46 (.B( u0_K4_12 ) , .A( u0_R2_9 ) , .Z( u0_u3_X_12 ) );
  XOR2_X1 u0_u3_U47 (.B( u0_K4_11 ) , .A( u0_R2_8 ) , .Z( u0_u3_X_11 ) );
  XOR2_X1 u0_u3_U48 (.B( u0_K4_10 ) , .A( u0_R2_7 ) , .Z( u0_u3_X_10 ) );
  XOR2_X1 u0_u3_U5 (.B( u0_K4_5 ) , .A( u0_R2_4 ) , .Z( u0_u3_X_5 ) );
  XOR2_X1 u0_u3_U6 (.B( u0_K4_4 ) , .A( u0_R2_3 ) , .Z( u0_u3_X_4 ) );
  AND2_X1 u0_u3_u0_U10 (.A1( u0_u3_u0_n133 ) , .ZN( u0_u3_u0_n143 ) , .A2( u0_u3_u0_n152 ) );
  AND2_X1 u0_u3_u0_U11 (.ZN( u0_u3_u0_n109 ) , .A1( u0_u3_u0_n132 ) , .A2( u0_u3_u0_n142 ) );
  AND2_X1 u0_u3_u0_U12 (.A2( u0_u3_u0_n131 ) , .A1( u0_u3_u0_n132 ) , .ZN( u0_u3_u0_n153 ) );
  AND2_X1 u0_u3_u0_U13 (.A1( u0_u3_u0_n110 ) , .A2( u0_u3_u0_n127 ) , .ZN( u0_u3_u0_n147 ) );
  INV_X1 u0_u3_u0_U14 (.A( u0_u3_u0_n145 ) , .ZN( u0_u3_u0_n175 ) );
  NOR2_X1 u0_u3_u0_U15 (.A2( u0_u3_u0_n138 ) , .ZN( u0_u3_u0_n149 ) , .A1( u0_u3_u0_n162 ) );
  AOI21_X1 u0_u3_u0_U16 (.B1( u0_u3_u0_n105 ) , .ZN( u0_u3_u0_n134 ) , .A( u0_u3_u0_n167 ) , .B2( u0_u3_u0_n95 ) );
  OAI22_X1 u0_u3_u0_U17 (.B1( u0_u3_u0_n133 ) , .A1( u0_u3_u0_n146 ) , .B2( u0_u3_u0_n149 ) , .A2( u0_u3_u0_n92 ) , .ZN( u0_u3_u0_n93 ) );
  AND3_X1 u0_u3_u0_U18 (.A3( u0_u3_u0_n123 ) , .A2( u0_u3_u0_n127 ) , .A1( u0_u3_u0_n150 ) , .ZN( u0_u3_u0_n92 ) );
  OAI22_X1 u0_u3_u0_U19 (.B1( u0_u3_u0_n127 ) , .ZN( u0_u3_u0_n128 ) , .A1( u0_u3_u0_n140 ) , .A2( u0_u3_u0_n148 ) , .B2( u0_u3_u0_n149 ) );
  NOR2_X1 u0_u3_u0_U20 (.A1( u0_u3_u0_n165 ) , .A2( u0_u3_u0_n166 ) , .ZN( u0_u3_u0_n97 ) );
  AOI22_X1 u0_u3_u0_U21 (.B2( u0_u3_u0_n111 ) , .A2( u0_u3_u0_n112 ) , .ZN( u0_u3_u0_n113 ) , .B1( u0_u3_u0_n120 ) , .A1( u0_u3_u0_n162 ) );
  NAND2_X1 u0_u3_u0_U22 (.A2( u0_u3_u0_n104 ) , .A1( u0_u3_u0_n105 ) , .ZN( u0_u3_u0_n151 ) );
  INV_X1 u0_u3_u0_U23 (.A( u0_u3_u0_n138 ) , .ZN( u0_u3_u0_n163 ) );
  INV_X1 u0_u3_u0_U24 (.A( u0_u3_u0_n120 ) , .ZN( u0_u3_u0_n160 ) );
  NAND2_X1 u0_u3_u0_U25 (.A2( u0_u3_u0_n102 ) , .ZN( u0_u3_u0_n133 ) , .A1( u0_u3_u0_n94 ) );
  NAND2_X1 u0_u3_u0_U26 (.ZN( u0_u3_u0_n110 ) , .A1( u0_u3_u0_n94 ) , .A2( u0_u3_u0_n96 ) );
  AOI21_X1 u0_u3_u0_U27 (.ZN( u0_u3_u0_n106 ) , .B1( u0_u3_u0_n109 ) , .B2( u0_u3_u0_n143 ) , .A( u0_u3_u0_n146 ) );
  AOI21_X1 u0_u3_u0_U28 (.B1( u0_u3_u0_n129 ) , .B2( u0_u3_u0_n131 ) , .A( u0_u3_u0_n140 ) , .ZN( u0_u3_u0_n98 ) );
  NAND2_X1 u0_u3_u0_U29 (.A2( u0_u3_u0_n104 ) , .ZN( u0_u3_u0_n116 ) , .A1( u0_u3_u0_n94 ) );
  INV_X1 u0_u3_u0_U3 (.A( u0_u3_u0_n115 ) , .ZN( u0_u3_u0_n168 ) );
  NOR2_X1 u0_u3_u0_U30 (.A1( u0_u3_u0_n122 ) , .ZN( u0_u3_u0_n145 ) , .A2( u0_u3_u0_n169 ) );
  OAI221_X1 u0_u3_u0_U31 (.C1( u0_u3_u0_n114 ) , .ZN( u0_u3_u0_n122 ) , .B1( u0_u3_u0_n140 ) , .B2( u0_u3_u0_n143 ) , .C2( u0_u3_u0_n149 ) , .A( u0_u3_u0_n174 ) );
  AOI211_X1 u0_u3_u0_U32 (.B( u0_u3_u0_n117 ) , .A( u0_u3_u0_n118 ) , .C2( u0_u3_u0_n119 ) , .C1( u0_u3_u0_n120 ) , .ZN( u0_u3_u0_n121 ) );
  NAND2_X1 u0_u3_u0_U33 (.A2( u0_u3_u0_n105 ) , .ZN( u0_u3_u0_n142 ) , .A1( u0_u3_u0_n96 ) );
  NAND2_X1 u0_u3_u0_U34 (.A1( u0_u3_u0_n102 ) , .A2( u0_u3_u0_n105 ) , .ZN( u0_u3_u0_n127 ) );
  NAND2_X1 u0_u3_u0_U35 (.A1( u0_u3_u0_n103 ) , .A2( u0_u3_u0_n104 ) , .ZN( u0_u3_u0_n152 ) );
  INV_X1 u0_u3_u0_U36 (.A( u0_u3_u0_n140 ) , .ZN( u0_u3_u0_n162 ) );
  NAND2_X1 u0_u3_u0_U37 (.A2( u0_u3_u0_n102 ) , .A1( u0_u3_u0_n103 ) , .ZN( u0_u3_u0_n141 ) );
  NAND2_X1 u0_u3_u0_U38 (.ZN( u0_u3_u0_n114 ) , .A2( u0_u3_u0_n94 ) , .A1( u0_u3_u0_n95 ) );
  NAND2_X1 u0_u3_u0_U39 (.A1( u0_u3_u0_n103 ) , .ZN( u0_u3_u0_n132 ) , .A2( u0_u3_u0_n96 ) );
  AOI21_X1 u0_u3_u0_U4 (.B1( u0_u3_u0_n116 ) , .ZN( u0_u3_u0_n117 ) , .B2( u0_u3_u0_n131 ) , .A( u0_u3_u0_n163 ) );
  INV_X1 u0_u3_u0_U40 (.ZN( u0_u3_u0_n174 ) , .A( u0_u3_u0_n90 ) );
  OAI222_X1 u0_u3_u0_U41 (.C1( u0_u3_u0_n110 ) , .A1( u0_u3_u0_n127 ) , .B2( u0_u3_u0_n130 ) , .B1( u0_u3_u0_n146 ) , .A2( u0_u3_u0_n160 ) , .C2( u0_u3_u0_n163 ) , .ZN( u0_u3_u0_n90 ) );
  OR3_X1 u0_u3_u0_U42 (.A3( u0_u3_u0_n154 ) , .A2( u0_u3_u0_n155 ) , .A1( u0_u3_u0_n156 ) , .ZN( u0_u3_u0_n157 ) );
  AOI21_X1 u0_u3_u0_U43 (.A( u0_u3_u0_n146 ) , .B2( u0_u3_u0_n147 ) , .B1( u0_u3_u0_n148 ) , .ZN( u0_u3_u0_n156 ) );
  AOI21_X1 u0_u3_u0_U44 (.B2( u0_u3_u0_n152 ) , .B1( u0_u3_u0_n153 ) , .ZN( u0_u3_u0_n154 ) , .A( u0_u3_u0_n160 ) );
  AOI21_X1 u0_u3_u0_U45 (.A( u0_u3_u0_n149 ) , .B2( u0_u3_u0_n150 ) , .B1( u0_u3_u0_n151 ) , .ZN( u0_u3_u0_n155 ) );
  INV_X1 u0_u3_u0_U46 (.A( u0_u3_u0_n101 ) , .ZN( u0_u3_u0_n173 ) );
  OAI211_X1 u0_u3_u0_U47 (.B( u0_u3_u0_n100 ) , .ZN( u0_u3_u0_n101 ) , .C2( u0_u3_u0_n142 ) , .C1( u0_u3_u0_n163 ) , .A( u0_u3_u0_n171 ) );
  INV_X1 u0_u3_u0_U48 (.ZN( u0_u3_u0_n171 ) , .A( u0_u3_u0_n93 ) );
  AOI211_X1 u0_u3_u0_U49 (.ZN( u0_u3_u0_n100 ) , .C1( u0_u3_u0_n120 ) , .A( u0_u3_u0_n125 ) , .B( u0_u3_u0_n98 ) , .C2( u0_u3_u0_n99 ) );
  AOI21_X1 u0_u3_u0_U5 (.B2( u0_u3_u0_n133 ) , .ZN( u0_u3_u0_n136 ) , .B1( u0_u3_u0_n153 ) , .A( u0_u3_u0_n160 ) );
  NOR2_X1 u0_u3_u0_U50 (.A2( u0_u3_X_4 ) , .A1( u0_u3_X_5 ) , .ZN( u0_u3_u0_n120 ) );
  NOR2_X1 u0_u3_u0_U51 (.A2( u0_u3_X_3 ) , .A1( u0_u3_X_6 ) , .ZN( u0_u3_u0_n96 ) );
  NOR2_X1 u0_u3_u0_U52 (.A2( u0_u3_X_6 ) , .ZN( u0_u3_u0_n102 ) , .A1( u0_u3_u0_n164 ) );
  NOR2_X1 u0_u3_u0_U53 (.A2( u0_u3_X_1 ) , .ZN( u0_u3_u0_n103 ) , .A1( u0_u3_u0_n165 ) );
  NAND2_X1 u0_u3_u0_U54 (.A2( u0_u3_X_4 ) , .A1( u0_u3_X_5 ) , .ZN( u0_u3_u0_n146 ) );
  NOR2_X1 u0_u3_u0_U55 (.A2( u0_u3_X_5 ) , .ZN( u0_u3_u0_n138 ) , .A1( u0_u3_u0_n161 ) );
  NAND2_X1 u0_u3_u0_U56 (.A1( u0_u3_X_5 ) , .ZN( u0_u3_u0_n140 ) , .A2( u0_u3_u0_n161 ) );
  AND2_X1 u0_u3_u0_U57 (.A2( u0_u3_X_3 ) , .A1( u0_u3_X_6 ) , .ZN( u0_u3_u0_n104 ) );
  AND2_X1 u0_u3_u0_U58 (.A1( u0_u3_X_6 ) , .A2( u0_u3_u0_n164 ) , .ZN( u0_u3_u0_n95 ) );
  INV_X1 u0_u3_u0_U59 (.A( u0_u3_X_4 ) , .ZN( u0_u3_u0_n161 ) );
  NOR2_X1 u0_u3_u0_U6 (.A1( u0_u3_u0_n110 ) , .ZN( u0_u3_u0_n125 ) , .A2( u0_u3_u0_n160 ) );
  INV_X1 u0_u3_u0_U60 (.A( u0_u3_X_1 ) , .ZN( u0_u3_u0_n166 ) );
  INV_X1 u0_u3_u0_U61 (.A( u0_u3_X_3 ) , .ZN( u0_u3_u0_n164 ) );
  INV_X1 u0_u3_u0_U62 (.A( u0_u3_u0_n128 ) , .ZN( u0_u3_u0_n170 ) );
  AOI211_X1 u0_u3_u0_U63 (.B( u0_u3_u0_n135 ) , .A( u0_u3_u0_n136 ) , .C2( u0_u3_u0_n137 ) , .C1( u0_u3_u0_n138 ) , .ZN( u0_u3_u0_n139 ) );
  OR4_X1 u0_u3_u0_U64 (.ZN( u0_out3_31 ) , .A4( u0_u3_u0_n157 ) , .A2( u0_u3_u0_n158 ) , .A1( u0_u3_u0_n159 ) , .A3( u0_u3_u0_n175 ) );
  AOI21_X1 u0_u3_u0_U65 (.A( u0_u3_u0_n140 ) , .B2( u0_u3_u0_n141 ) , .B1( u0_u3_u0_n142 ) , .ZN( u0_u3_u0_n159 ) );
  OR4_X1 u0_u3_u0_U66 (.ZN( u0_out3_17 ) , .A4( u0_u3_u0_n124 ) , .A2( u0_u3_u0_n125 ) , .A1( u0_u3_u0_n126 ) , .A3( u0_u3_u0_n172 ) );
  AOI21_X1 u0_u3_u0_U67 (.B2( u0_u3_u0_n109 ) , .ZN( u0_u3_u0_n126 ) , .B1( u0_u3_u0_n130 ) , .A( u0_u3_u0_n163 ) );
  INV_X1 u0_u3_u0_U68 (.A( u0_u3_u0_n113 ) , .ZN( u0_u3_u0_n172 ) );
  INV_X1 u0_u3_u0_U69 (.ZN( u0_u3_u0_n176 ) , .A( u0_u3_u0_n91 ) );
  OAI21_X1 u0_u3_u0_U7 (.B1( u0_u3_u0_n152 ) , .B2( u0_u3_u0_n160 ) , .A( u0_u3_u0_n174 ) , .ZN( u0_u3_u0_n91 ) );
  AOI211_X1 u0_u3_u0_U70 (.B( u0_u3_u0_n106 ) , .A( u0_u3_u0_n107 ) , .ZN( u0_u3_u0_n108 ) , .C2( u0_u3_u0_n115 ) , .C1( u0_u3_u0_n162 ) );
  AOI21_X1 u0_u3_u0_U71 (.B2( u0_u3_u0_n143 ) , .B1( u0_u3_u0_n144 ) , .ZN( u0_u3_u0_n158 ) , .A( u0_u3_u0_n163 ) );
  AOI21_X1 u0_u3_u0_U72 (.ZN( u0_u3_u0_n118 ) , .B2( u0_u3_u0_n144 ) , .A( u0_u3_u0_n146 ) , .B1( u0_u3_u0_n168 ) );
  INV_X1 u0_u3_u0_U73 (.A( u0_u3_u0_n144 ) , .ZN( u0_u3_u0_n167 ) );
  NOR2_X1 u0_u3_u0_U74 (.A2( u0_u3_X_1 ) , .A1( u0_u3_X_2 ) , .ZN( u0_u3_u0_n94 ) );
  NOR2_X1 u0_u3_u0_U75 (.A2( u0_u3_X_2 ) , .ZN( u0_u3_u0_n105 ) , .A1( u0_u3_u0_n166 ) );
  INV_X1 u0_u3_u0_U76 (.A( u0_u3_X_2 ) , .ZN( u0_u3_u0_n165 ) );
  OR2_X1 u0_u3_u0_U77 (.A2( u0_u3_u0_n129 ) , .A1( u0_u3_u0_n146 ) , .ZN( u0_u3_u0_n88 ) );
  OR2_X1 u0_u3_u0_U78 (.A1( u0_u3_u0_n123 ) , .A2( u0_u3_u0_n149 ) , .ZN( u0_u3_u0_n89 ) );
  NAND3_X1 u0_u3_u0_U79 (.ZN( u0_u3_u0_n124 ) , .A3( u0_u3_u0_n145 ) , .A1( u0_u3_u0_n88 ) , .A2( u0_u3_u0_n89 ) );
  AND2_X1 u0_u3_u0_U8 (.A1( u0_u3_u0_n116 ) , .A2( u0_u3_u0_n123 ) , .ZN( u0_u3_u0_n148 ) );
  AND3_X1 u0_u3_u0_U80 (.A2( u0_u3_u0_n114 ) , .ZN( u0_u3_u0_n129 ) , .A3( u0_u3_u0_n132 ) , .A1( u0_u3_u0_n150 ) );
  NAND2_X1 u0_u3_u0_U81 (.A2( u0_u3_u0_n103 ) , .ZN( u0_u3_u0_n123 ) , .A1( u0_u3_u0_n95 ) );
  AOI21_X1 u0_u3_u0_U82 (.B1( u0_u3_u0_n134 ) , .ZN( u0_u3_u0_n135 ) , .A( u0_u3_u0_n146 ) , .B2( u0_u3_u0_n168 ) );
  OAI22_X1 u0_u3_u0_U83 (.ZN( u0_u3_u0_n107 ) , .A2( u0_u3_u0_n134 ) , .B1( u0_u3_u0_n148 ) , .A1( u0_u3_u0_n149 ) , .B2( u0_u3_u0_n163 ) );
  NAND2_X1 u0_u3_u0_U84 (.ZN( u0_u3_u0_n112 ) , .A2( u0_u3_u0_n134 ) , .A1( u0_u3_u0_n147 ) );
  INV_X1 u0_u3_u0_U85 (.A( u0_u3_u0_n121 ) , .ZN( u0_u3_u0_n169 ) );
  NAND2_X1 u0_u3_u0_U86 (.ZN( u0_u3_u0_n150 ) , .A1( u0_u3_u0_n95 ) , .A2( u0_u3_u0_n97 ) );
  NAND2_X1 u0_u3_u0_U87 (.A1( u0_u3_u0_n102 ) , .ZN( u0_u3_u0_n131 ) , .A2( u0_u3_u0_n97 ) );
  NAND3_X1 u0_u3_u0_U88 (.ZN( u0_out3_23 ) , .A3( u0_u3_u0_n139 ) , .A1( u0_u3_u0_n170 ) , .A2( u0_u3_u0_n173 ) );
  NAND3_X1 u0_u3_u0_U89 (.A3( u0_u3_u0_n129 ) , .A2( u0_u3_u0_n130 ) , .ZN( u0_u3_u0_n137 ) , .A1( u0_u3_u0_n152 ) );
  NAND2_X1 u0_u3_u0_U9 (.ZN( u0_u3_u0_n115 ) , .A1( u0_u3_u0_n141 ) , .A2( u0_u3_u0_n151 ) );
  NAND3_X1 u0_u3_u0_U90 (.ZN( u0_u3_u0_n119 ) , .A3( u0_u3_u0_n134 ) , .A2( u0_u3_u0_n141 ) , .A1( u0_u3_u0_n150 ) );
  NAND3_X1 u0_u3_u0_U91 (.ZN( u0_u3_u0_n111 ) , .A2( u0_u3_u0_n116 ) , .A3( u0_u3_u0_n142 ) , .A1( u0_u3_u0_n151 ) );
  NAND3_X1 u0_u3_u0_U92 (.ZN( u0_out3_9 ) , .A3( u0_u3_u0_n108 ) , .A2( u0_u3_u0_n173 ) , .A1( u0_u3_u0_n176 ) );
  NAND3_X1 u0_u3_u0_U93 (.A2( u0_u3_u0_n130 ) , .A1( u0_u3_u0_n134 ) , .A3( u0_u3_u0_n148 ) , .ZN( u0_u3_u0_n99 ) );
  NAND2_X1 u0_u3_u0_U94 (.A1( u0_u3_u0_n104 ) , .ZN( u0_u3_u0_n130 ) , .A2( u0_u3_u0_n97 ) );
  NAND2_X1 u0_u3_u0_U95 (.ZN( u0_u3_u0_n144 ) , .A1( u0_u3_u0_n96 ) , .A2( u0_u3_u0_n97 ) );
  NOR2_X1 u0_u3_u1_U10 (.A1( u0_u3_u1_n112 ) , .A2( u0_u3_u1_n116 ) , .ZN( u0_u3_u1_n118 ) );
  NAND3_X1 u0_u3_u1_U100 (.ZN( u0_u3_u1_n113 ) , .A1( u0_u3_u1_n120 ) , .A3( u0_u3_u1_n133 ) , .A2( u0_u3_u1_n155 ) );
  OAI21_X1 u0_u3_u1_U11 (.ZN( u0_u3_u1_n101 ) , .B1( u0_u3_u1_n141 ) , .A( u0_u3_u1_n146 ) , .B2( u0_u3_u1_n183 ) );
  AOI21_X1 u0_u3_u1_U12 (.B2( u0_u3_u1_n155 ) , .B1( u0_u3_u1_n156 ) , .ZN( u0_u3_u1_n157 ) , .A( u0_u3_u1_n174 ) );
  NAND2_X1 u0_u3_u1_U13 (.ZN( u0_u3_u1_n140 ) , .A2( u0_u3_u1_n150 ) , .A1( u0_u3_u1_n155 ) );
  NAND2_X1 u0_u3_u1_U14 (.A1( u0_u3_u1_n131 ) , .ZN( u0_u3_u1_n147 ) , .A2( u0_u3_u1_n153 ) );
  INV_X1 u0_u3_u1_U15 (.A( u0_u3_u1_n139 ) , .ZN( u0_u3_u1_n174 ) );
  OR4_X1 u0_u3_u1_U16 (.A4( u0_u3_u1_n106 ) , .A3( u0_u3_u1_n107 ) , .ZN( u0_u3_u1_n108 ) , .A1( u0_u3_u1_n117 ) , .A2( u0_u3_u1_n184 ) );
  AOI21_X1 u0_u3_u1_U17 (.ZN( u0_u3_u1_n106 ) , .A( u0_u3_u1_n112 ) , .B1( u0_u3_u1_n154 ) , .B2( u0_u3_u1_n156 ) );
  INV_X1 u0_u3_u1_U18 (.A( u0_u3_u1_n101 ) , .ZN( u0_u3_u1_n184 ) );
  AOI21_X1 u0_u3_u1_U19 (.ZN( u0_u3_u1_n107 ) , .B1( u0_u3_u1_n134 ) , .B2( u0_u3_u1_n149 ) , .A( u0_u3_u1_n174 ) );
  INV_X1 u0_u3_u1_U20 (.A( u0_u3_u1_n112 ) , .ZN( u0_u3_u1_n171 ) );
  NAND2_X1 u0_u3_u1_U21 (.ZN( u0_u3_u1_n141 ) , .A1( u0_u3_u1_n153 ) , .A2( u0_u3_u1_n156 ) );
  AND2_X1 u0_u3_u1_U22 (.A1( u0_u3_u1_n123 ) , .ZN( u0_u3_u1_n134 ) , .A2( u0_u3_u1_n161 ) );
  NAND2_X1 u0_u3_u1_U23 (.A2( u0_u3_u1_n115 ) , .A1( u0_u3_u1_n116 ) , .ZN( u0_u3_u1_n148 ) );
  NAND2_X1 u0_u3_u1_U24 (.A2( u0_u3_u1_n133 ) , .A1( u0_u3_u1_n135 ) , .ZN( u0_u3_u1_n159 ) );
  NAND2_X1 u0_u3_u1_U25 (.A2( u0_u3_u1_n115 ) , .A1( u0_u3_u1_n120 ) , .ZN( u0_u3_u1_n132 ) );
  INV_X1 u0_u3_u1_U26 (.A( u0_u3_u1_n154 ) , .ZN( u0_u3_u1_n178 ) );
  INV_X1 u0_u3_u1_U27 (.A( u0_u3_u1_n151 ) , .ZN( u0_u3_u1_n183 ) );
  AND2_X1 u0_u3_u1_U28 (.A1( u0_u3_u1_n129 ) , .A2( u0_u3_u1_n133 ) , .ZN( u0_u3_u1_n149 ) );
  INV_X1 u0_u3_u1_U29 (.A( u0_u3_u1_n131 ) , .ZN( u0_u3_u1_n180 ) );
  INV_X1 u0_u3_u1_U3 (.A( u0_u3_u1_n159 ) , .ZN( u0_u3_u1_n182 ) );
  AOI221_X1 u0_u3_u1_U30 (.B1( u0_u3_u1_n140 ) , .ZN( u0_u3_u1_n167 ) , .B2( u0_u3_u1_n172 ) , .C2( u0_u3_u1_n175 ) , .C1( u0_u3_u1_n178 ) , .A( u0_u3_u1_n188 ) );
  INV_X1 u0_u3_u1_U31 (.ZN( u0_u3_u1_n188 ) , .A( u0_u3_u1_n97 ) );
  AOI211_X1 u0_u3_u1_U32 (.A( u0_u3_u1_n118 ) , .C1( u0_u3_u1_n132 ) , .C2( u0_u3_u1_n139 ) , .B( u0_u3_u1_n96 ) , .ZN( u0_u3_u1_n97 ) );
  AOI21_X1 u0_u3_u1_U33 (.B2( u0_u3_u1_n121 ) , .B1( u0_u3_u1_n135 ) , .A( u0_u3_u1_n152 ) , .ZN( u0_u3_u1_n96 ) );
  OAI221_X1 u0_u3_u1_U34 (.A( u0_u3_u1_n119 ) , .C2( u0_u3_u1_n129 ) , .ZN( u0_u3_u1_n138 ) , .B2( u0_u3_u1_n152 ) , .C1( u0_u3_u1_n174 ) , .B1( u0_u3_u1_n187 ) );
  INV_X1 u0_u3_u1_U35 (.A( u0_u3_u1_n148 ) , .ZN( u0_u3_u1_n187 ) );
  AOI211_X1 u0_u3_u1_U36 (.B( u0_u3_u1_n117 ) , .A( u0_u3_u1_n118 ) , .ZN( u0_u3_u1_n119 ) , .C2( u0_u3_u1_n146 ) , .C1( u0_u3_u1_n159 ) );
  NOR2_X1 u0_u3_u1_U37 (.A1( u0_u3_u1_n168 ) , .A2( u0_u3_u1_n176 ) , .ZN( u0_u3_u1_n98 ) );
  NAND2_X1 u0_u3_u1_U38 (.A1( u0_u3_u1_n128 ) , .ZN( u0_u3_u1_n146 ) , .A2( u0_u3_u1_n160 ) );
  NAND2_X1 u0_u3_u1_U39 (.A2( u0_u3_u1_n112 ) , .ZN( u0_u3_u1_n139 ) , .A1( u0_u3_u1_n152 ) );
  AOI221_X1 u0_u3_u1_U4 (.A( u0_u3_u1_n138 ) , .C2( u0_u3_u1_n139 ) , .C1( u0_u3_u1_n140 ) , .B2( u0_u3_u1_n141 ) , .ZN( u0_u3_u1_n142 ) , .B1( u0_u3_u1_n175 ) );
  NAND2_X1 u0_u3_u1_U40 (.A1( u0_u3_u1_n105 ) , .ZN( u0_u3_u1_n156 ) , .A2( u0_u3_u1_n99 ) );
  NOR2_X1 u0_u3_u1_U41 (.ZN( u0_u3_u1_n117 ) , .A1( u0_u3_u1_n121 ) , .A2( u0_u3_u1_n160 ) );
  OAI21_X1 u0_u3_u1_U42 (.B2( u0_u3_u1_n123 ) , .ZN( u0_u3_u1_n145 ) , .B1( u0_u3_u1_n160 ) , .A( u0_u3_u1_n185 ) );
  INV_X1 u0_u3_u1_U43 (.A( u0_u3_u1_n122 ) , .ZN( u0_u3_u1_n185 ) );
  AOI21_X1 u0_u3_u1_U44 (.B2( u0_u3_u1_n120 ) , .B1( u0_u3_u1_n121 ) , .ZN( u0_u3_u1_n122 ) , .A( u0_u3_u1_n128 ) );
  AOI21_X1 u0_u3_u1_U45 (.A( u0_u3_u1_n128 ) , .B2( u0_u3_u1_n129 ) , .ZN( u0_u3_u1_n130 ) , .B1( u0_u3_u1_n150 ) );
  NAND2_X1 u0_u3_u1_U46 (.ZN( u0_u3_u1_n112 ) , .A1( u0_u3_u1_n169 ) , .A2( u0_u3_u1_n170 ) );
  NAND2_X1 u0_u3_u1_U47 (.ZN( u0_u3_u1_n129 ) , .A2( u0_u3_u1_n95 ) , .A1( u0_u3_u1_n98 ) );
  NAND2_X1 u0_u3_u1_U48 (.A1( u0_u3_u1_n102 ) , .ZN( u0_u3_u1_n154 ) , .A2( u0_u3_u1_n99 ) );
  NAND2_X1 u0_u3_u1_U49 (.A2( u0_u3_u1_n100 ) , .ZN( u0_u3_u1_n135 ) , .A1( u0_u3_u1_n99 ) );
  AOI211_X1 u0_u3_u1_U5 (.ZN( u0_u3_u1_n124 ) , .A( u0_u3_u1_n138 ) , .C2( u0_u3_u1_n139 ) , .B( u0_u3_u1_n145 ) , .C1( u0_u3_u1_n147 ) );
  AOI21_X1 u0_u3_u1_U50 (.A( u0_u3_u1_n152 ) , .B2( u0_u3_u1_n153 ) , .B1( u0_u3_u1_n154 ) , .ZN( u0_u3_u1_n158 ) );
  INV_X1 u0_u3_u1_U51 (.A( u0_u3_u1_n160 ) , .ZN( u0_u3_u1_n175 ) );
  NAND2_X1 u0_u3_u1_U52 (.A1( u0_u3_u1_n100 ) , .ZN( u0_u3_u1_n116 ) , .A2( u0_u3_u1_n95 ) );
  NAND2_X1 u0_u3_u1_U53 (.A1( u0_u3_u1_n102 ) , .ZN( u0_u3_u1_n131 ) , .A2( u0_u3_u1_n95 ) );
  NAND2_X1 u0_u3_u1_U54 (.A2( u0_u3_u1_n104 ) , .ZN( u0_u3_u1_n121 ) , .A1( u0_u3_u1_n98 ) );
  NAND2_X1 u0_u3_u1_U55 (.A1( u0_u3_u1_n103 ) , .ZN( u0_u3_u1_n153 ) , .A2( u0_u3_u1_n98 ) );
  NAND2_X1 u0_u3_u1_U56 (.A2( u0_u3_u1_n104 ) , .A1( u0_u3_u1_n105 ) , .ZN( u0_u3_u1_n133 ) );
  NAND2_X1 u0_u3_u1_U57 (.ZN( u0_u3_u1_n150 ) , .A2( u0_u3_u1_n98 ) , .A1( u0_u3_u1_n99 ) );
  NAND2_X1 u0_u3_u1_U58 (.A1( u0_u3_u1_n105 ) , .ZN( u0_u3_u1_n155 ) , .A2( u0_u3_u1_n95 ) );
  OAI21_X1 u0_u3_u1_U59 (.ZN( u0_u3_u1_n109 ) , .B1( u0_u3_u1_n129 ) , .B2( u0_u3_u1_n160 ) , .A( u0_u3_u1_n167 ) );
  AOI22_X1 u0_u3_u1_U6 (.B2( u0_u3_u1_n113 ) , .A2( u0_u3_u1_n114 ) , .ZN( u0_u3_u1_n125 ) , .A1( u0_u3_u1_n171 ) , .B1( u0_u3_u1_n173 ) );
  NAND2_X1 u0_u3_u1_U60 (.A2( u0_u3_u1_n100 ) , .A1( u0_u3_u1_n103 ) , .ZN( u0_u3_u1_n120 ) );
  NAND2_X1 u0_u3_u1_U61 (.A1( u0_u3_u1_n102 ) , .A2( u0_u3_u1_n104 ) , .ZN( u0_u3_u1_n115 ) );
  NAND2_X1 u0_u3_u1_U62 (.A2( u0_u3_u1_n100 ) , .A1( u0_u3_u1_n104 ) , .ZN( u0_u3_u1_n151 ) );
  NAND2_X1 u0_u3_u1_U63 (.A2( u0_u3_u1_n103 ) , .A1( u0_u3_u1_n105 ) , .ZN( u0_u3_u1_n161 ) );
  INV_X1 u0_u3_u1_U64 (.A( u0_u3_u1_n152 ) , .ZN( u0_u3_u1_n173 ) );
  INV_X1 u0_u3_u1_U65 (.A( u0_u3_u1_n128 ) , .ZN( u0_u3_u1_n172 ) );
  NAND2_X1 u0_u3_u1_U66 (.A2( u0_u3_u1_n102 ) , .A1( u0_u3_u1_n103 ) , .ZN( u0_u3_u1_n123 ) );
  AOI211_X1 u0_u3_u1_U67 (.B( u0_u3_u1_n162 ) , .A( u0_u3_u1_n163 ) , .C2( u0_u3_u1_n164 ) , .ZN( u0_u3_u1_n165 ) , .C1( u0_u3_u1_n171 ) );
  AOI21_X1 u0_u3_u1_U68 (.A( u0_u3_u1_n160 ) , .B2( u0_u3_u1_n161 ) , .ZN( u0_u3_u1_n162 ) , .B1( u0_u3_u1_n182 ) );
  OR2_X1 u0_u3_u1_U69 (.A2( u0_u3_u1_n157 ) , .A1( u0_u3_u1_n158 ) , .ZN( u0_u3_u1_n163 ) );
  NAND2_X1 u0_u3_u1_U7 (.ZN( u0_u3_u1_n114 ) , .A1( u0_u3_u1_n134 ) , .A2( u0_u3_u1_n156 ) );
  NOR2_X1 u0_u3_u1_U70 (.A2( u0_u3_X_7 ) , .A1( u0_u3_X_8 ) , .ZN( u0_u3_u1_n95 ) );
  NOR2_X1 u0_u3_u1_U71 (.A1( u0_u3_X_12 ) , .A2( u0_u3_X_9 ) , .ZN( u0_u3_u1_n100 ) );
  NOR2_X1 u0_u3_u1_U72 (.A2( u0_u3_X_8 ) , .A1( u0_u3_u1_n177 ) , .ZN( u0_u3_u1_n99 ) );
  NOR2_X1 u0_u3_u1_U73 (.A2( u0_u3_X_12 ) , .ZN( u0_u3_u1_n102 ) , .A1( u0_u3_u1_n176 ) );
  NOR2_X1 u0_u3_u1_U74 (.A2( u0_u3_X_9 ) , .ZN( u0_u3_u1_n105 ) , .A1( u0_u3_u1_n168 ) );
  NAND2_X1 u0_u3_u1_U75 (.A1( u0_u3_X_10 ) , .ZN( u0_u3_u1_n160 ) , .A2( u0_u3_u1_n169 ) );
  NAND2_X1 u0_u3_u1_U76 (.A2( u0_u3_X_10 ) , .A1( u0_u3_X_11 ) , .ZN( u0_u3_u1_n152 ) );
  NAND2_X1 u0_u3_u1_U77 (.A1( u0_u3_X_11 ) , .ZN( u0_u3_u1_n128 ) , .A2( u0_u3_u1_n170 ) );
  AND2_X1 u0_u3_u1_U78 (.A2( u0_u3_X_7 ) , .A1( u0_u3_X_8 ) , .ZN( u0_u3_u1_n104 ) );
  AND2_X1 u0_u3_u1_U79 (.A1( u0_u3_X_8 ) , .ZN( u0_u3_u1_n103 ) , .A2( u0_u3_u1_n177 ) );
  AOI22_X1 u0_u3_u1_U8 (.B2( u0_u3_u1_n136 ) , .A2( u0_u3_u1_n137 ) , .ZN( u0_u3_u1_n143 ) , .A1( u0_u3_u1_n171 ) , .B1( u0_u3_u1_n173 ) );
  INV_X1 u0_u3_u1_U80 (.A( u0_u3_X_10 ) , .ZN( u0_u3_u1_n170 ) );
  INV_X1 u0_u3_u1_U81 (.A( u0_u3_X_9 ) , .ZN( u0_u3_u1_n176 ) );
  INV_X1 u0_u3_u1_U82 (.A( u0_u3_X_11 ) , .ZN( u0_u3_u1_n169 ) );
  INV_X1 u0_u3_u1_U83 (.A( u0_u3_X_12 ) , .ZN( u0_u3_u1_n168 ) );
  INV_X1 u0_u3_u1_U84 (.A( u0_u3_X_7 ) , .ZN( u0_u3_u1_n177 ) );
  NAND4_X1 u0_u3_u1_U85 (.ZN( u0_out3_28 ) , .A4( u0_u3_u1_n124 ) , .A3( u0_u3_u1_n125 ) , .A2( u0_u3_u1_n126 ) , .A1( u0_u3_u1_n127 ) );
  OAI21_X1 u0_u3_u1_U86 (.ZN( u0_u3_u1_n127 ) , .B2( u0_u3_u1_n139 ) , .B1( u0_u3_u1_n175 ) , .A( u0_u3_u1_n183 ) );
  OAI21_X1 u0_u3_u1_U87 (.ZN( u0_u3_u1_n126 ) , .B2( u0_u3_u1_n140 ) , .A( u0_u3_u1_n146 ) , .B1( u0_u3_u1_n178 ) );
  NAND4_X1 u0_u3_u1_U88 (.ZN( u0_out3_18 ) , .A4( u0_u3_u1_n165 ) , .A3( u0_u3_u1_n166 ) , .A1( u0_u3_u1_n167 ) , .A2( u0_u3_u1_n186 ) );
  AOI22_X1 u0_u3_u1_U89 (.B2( u0_u3_u1_n146 ) , .B1( u0_u3_u1_n147 ) , .A2( u0_u3_u1_n148 ) , .ZN( u0_u3_u1_n166 ) , .A1( u0_u3_u1_n172 ) );
  INV_X1 u0_u3_u1_U9 (.A( u0_u3_u1_n147 ) , .ZN( u0_u3_u1_n181 ) );
  INV_X1 u0_u3_u1_U90 (.A( u0_u3_u1_n145 ) , .ZN( u0_u3_u1_n186 ) );
  NAND4_X1 u0_u3_u1_U91 (.ZN( u0_out3_2 ) , .A4( u0_u3_u1_n142 ) , .A3( u0_u3_u1_n143 ) , .A2( u0_u3_u1_n144 ) , .A1( u0_u3_u1_n179 ) );
  INV_X1 u0_u3_u1_U92 (.A( u0_u3_u1_n130 ) , .ZN( u0_u3_u1_n179 ) );
  OAI21_X1 u0_u3_u1_U93 (.B2( u0_u3_u1_n132 ) , .ZN( u0_u3_u1_n144 ) , .A( u0_u3_u1_n146 ) , .B1( u0_u3_u1_n180 ) );
  OR4_X1 u0_u3_u1_U94 (.ZN( u0_out3_13 ) , .A4( u0_u3_u1_n108 ) , .A3( u0_u3_u1_n109 ) , .A2( u0_u3_u1_n110 ) , .A1( u0_u3_u1_n111 ) );
  AOI21_X1 u0_u3_u1_U95 (.ZN( u0_u3_u1_n111 ) , .A( u0_u3_u1_n128 ) , .B2( u0_u3_u1_n131 ) , .B1( u0_u3_u1_n135 ) );
  AOI21_X1 u0_u3_u1_U96 (.ZN( u0_u3_u1_n110 ) , .A( u0_u3_u1_n116 ) , .B1( u0_u3_u1_n152 ) , .B2( u0_u3_u1_n160 ) );
  NAND3_X1 u0_u3_u1_U97 (.A3( u0_u3_u1_n149 ) , .A2( u0_u3_u1_n150 ) , .A1( u0_u3_u1_n151 ) , .ZN( u0_u3_u1_n164 ) );
  NAND3_X1 u0_u3_u1_U98 (.A3( u0_u3_u1_n134 ) , .A2( u0_u3_u1_n135 ) , .ZN( u0_u3_u1_n136 ) , .A1( u0_u3_u1_n151 ) );
  NAND3_X1 u0_u3_u1_U99 (.A1( u0_u3_u1_n133 ) , .ZN( u0_u3_u1_n137 ) , .A2( u0_u3_u1_n154 ) , .A3( u0_u3_u1_n181 ) );
  OAI22_X1 u0_u3_u2_U10 (.B1( u0_u3_u2_n151 ) , .A2( u0_u3_u2_n152 ) , .A1( u0_u3_u2_n153 ) , .ZN( u0_u3_u2_n160 ) , .B2( u0_u3_u2_n168 ) );
  NAND3_X1 u0_u3_u2_U100 (.A2( u0_u3_u2_n100 ) , .A1( u0_u3_u2_n104 ) , .A3( u0_u3_u2_n138 ) , .ZN( u0_u3_u2_n98 ) );
  NOR3_X1 u0_u3_u2_U11 (.A1( u0_u3_u2_n150 ) , .ZN( u0_u3_u2_n151 ) , .A3( u0_u3_u2_n175 ) , .A2( u0_u3_u2_n188 ) );
  AOI21_X1 u0_u3_u2_U12 (.B2( u0_u3_u2_n123 ) , .ZN( u0_u3_u2_n125 ) , .A( u0_u3_u2_n171 ) , .B1( u0_u3_u2_n184 ) );
  INV_X1 u0_u3_u2_U13 (.A( u0_u3_u2_n150 ) , .ZN( u0_u3_u2_n184 ) );
  AOI21_X1 u0_u3_u2_U14 (.ZN( u0_u3_u2_n144 ) , .B2( u0_u3_u2_n155 ) , .A( u0_u3_u2_n172 ) , .B1( u0_u3_u2_n185 ) );
  AOI21_X1 u0_u3_u2_U15 (.B2( u0_u3_u2_n143 ) , .ZN( u0_u3_u2_n145 ) , .B1( u0_u3_u2_n152 ) , .A( u0_u3_u2_n171 ) );
  INV_X1 u0_u3_u2_U16 (.A( u0_u3_u2_n156 ) , .ZN( u0_u3_u2_n171 ) );
  INV_X1 u0_u3_u2_U17 (.A( u0_u3_u2_n120 ) , .ZN( u0_u3_u2_n188 ) );
  NAND2_X1 u0_u3_u2_U18 (.A2( u0_u3_u2_n122 ) , .ZN( u0_u3_u2_n150 ) , .A1( u0_u3_u2_n152 ) );
  INV_X1 u0_u3_u2_U19 (.A( u0_u3_u2_n153 ) , .ZN( u0_u3_u2_n170 ) );
  INV_X1 u0_u3_u2_U20 (.A( u0_u3_u2_n137 ) , .ZN( u0_u3_u2_n173 ) );
  NAND2_X1 u0_u3_u2_U21 (.A1( u0_u3_u2_n132 ) , .A2( u0_u3_u2_n139 ) , .ZN( u0_u3_u2_n157 ) );
  INV_X1 u0_u3_u2_U22 (.A( u0_u3_u2_n113 ) , .ZN( u0_u3_u2_n178 ) );
  INV_X1 u0_u3_u2_U23 (.A( u0_u3_u2_n139 ) , .ZN( u0_u3_u2_n175 ) );
  INV_X1 u0_u3_u2_U24 (.A( u0_u3_u2_n155 ) , .ZN( u0_u3_u2_n181 ) );
  INV_X1 u0_u3_u2_U25 (.A( u0_u3_u2_n119 ) , .ZN( u0_u3_u2_n177 ) );
  INV_X1 u0_u3_u2_U26 (.A( u0_u3_u2_n116 ) , .ZN( u0_u3_u2_n180 ) );
  INV_X1 u0_u3_u2_U27 (.A( u0_u3_u2_n131 ) , .ZN( u0_u3_u2_n179 ) );
  INV_X1 u0_u3_u2_U28 (.A( u0_u3_u2_n154 ) , .ZN( u0_u3_u2_n176 ) );
  NAND2_X1 u0_u3_u2_U29 (.A2( u0_u3_u2_n116 ) , .A1( u0_u3_u2_n117 ) , .ZN( u0_u3_u2_n118 ) );
  NOR2_X1 u0_u3_u2_U3 (.ZN( u0_u3_u2_n121 ) , .A2( u0_u3_u2_n177 ) , .A1( u0_u3_u2_n180 ) );
  INV_X1 u0_u3_u2_U30 (.A( u0_u3_u2_n132 ) , .ZN( u0_u3_u2_n182 ) );
  INV_X1 u0_u3_u2_U31 (.A( u0_u3_u2_n158 ) , .ZN( u0_u3_u2_n183 ) );
  OAI21_X1 u0_u3_u2_U32 (.A( u0_u3_u2_n156 ) , .B1( u0_u3_u2_n157 ) , .ZN( u0_u3_u2_n158 ) , .B2( u0_u3_u2_n179 ) );
  NOR2_X1 u0_u3_u2_U33 (.ZN( u0_u3_u2_n156 ) , .A1( u0_u3_u2_n166 ) , .A2( u0_u3_u2_n169 ) );
  NOR2_X1 u0_u3_u2_U34 (.A2( u0_u3_u2_n114 ) , .ZN( u0_u3_u2_n137 ) , .A1( u0_u3_u2_n140 ) );
  NOR2_X1 u0_u3_u2_U35 (.A2( u0_u3_u2_n138 ) , .ZN( u0_u3_u2_n153 ) , .A1( u0_u3_u2_n156 ) );
  AOI211_X1 u0_u3_u2_U36 (.ZN( u0_u3_u2_n130 ) , .C1( u0_u3_u2_n138 ) , .C2( u0_u3_u2_n179 ) , .B( u0_u3_u2_n96 ) , .A( u0_u3_u2_n97 ) );
  OAI22_X1 u0_u3_u2_U37 (.B1( u0_u3_u2_n133 ) , .A2( u0_u3_u2_n137 ) , .A1( u0_u3_u2_n152 ) , .B2( u0_u3_u2_n168 ) , .ZN( u0_u3_u2_n97 ) );
  OAI221_X1 u0_u3_u2_U38 (.B1( u0_u3_u2_n113 ) , .C1( u0_u3_u2_n132 ) , .A( u0_u3_u2_n149 ) , .B2( u0_u3_u2_n171 ) , .C2( u0_u3_u2_n172 ) , .ZN( u0_u3_u2_n96 ) );
  OAI221_X1 u0_u3_u2_U39 (.A( u0_u3_u2_n115 ) , .C2( u0_u3_u2_n123 ) , .B2( u0_u3_u2_n143 ) , .B1( u0_u3_u2_n153 ) , .ZN( u0_u3_u2_n163 ) , .C1( u0_u3_u2_n168 ) );
  INV_X1 u0_u3_u2_U4 (.A( u0_u3_u2_n134 ) , .ZN( u0_u3_u2_n185 ) );
  OAI21_X1 u0_u3_u2_U40 (.A( u0_u3_u2_n114 ) , .ZN( u0_u3_u2_n115 ) , .B1( u0_u3_u2_n176 ) , .B2( u0_u3_u2_n178 ) );
  OAI221_X1 u0_u3_u2_U41 (.A( u0_u3_u2_n135 ) , .B2( u0_u3_u2_n136 ) , .B1( u0_u3_u2_n137 ) , .ZN( u0_u3_u2_n162 ) , .C2( u0_u3_u2_n167 ) , .C1( u0_u3_u2_n185 ) );
  AND3_X1 u0_u3_u2_U42 (.A3( u0_u3_u2_n131 ) , .A2( u0_u3_u2_n132 ) , .A1( u0_u3_u2_n133 ) , .ZN( u0_u3_u2_n136 ) );
  AOI22_X1 u0_u3_u2_U43 (.ZN( u0_u3_u2_n135 ) , .B1( u0_u3_u2_n140 ) , .A1( u0_u3_u2_n156 ) , .B2( u0_u3_u2_n180 ) , .A2( u0_u3_u2_n188 ) );
  AOI21_X1 u0_u3_u2_U44 (.ZN( u0_u3_u2_n149 ) , .B1( u0_u3_u2_n173 ) , .B2( u0_u3_u2_n188 ) , .A( u0_u3_u2_n95 ) );
  AND3_X1 u0_u3_u2_U45 (.A2( u0_u3_u2_n100 ) , .A1( u0_u3_u2_n104 ) , .A3( u0_u3_u2_n156 ) , .ZN( u0_u3_u2_n95 ) );
  OAI21_X1 u0_u3_u2_U46 (.A( u0_u3_u2_n141 ) , .B2( u0_u3_u2_n142 ) , .ZN( u0_u3_u2_n146 ) , .B1( u0_u3_u2_n153 ) );
  OAI21_X1 u0_u3_u2_U47 (.A( u0_u3_u2_n140 ) , .ZN( u0_u3_u2_n141 ) , .B1( u0_u3_u2_n176 ) , .B2( u0_u3_u2_n177 ) );
  NOR3_X1 u0_u3_u2_U48 (.ZN( u0_u3_u2_n142 ) , .A3( u0_u3_u2_n175 ) , .A2( u0_u3_u2_n178 ) , .A1( u0_u3_u2_n181 ) );
  OAI21_X1 u0_u3_u2_U49 (.A( u0_u3_u2_n101 ) , .B2( u0_u3_u2_n121 ) , .B1( u0_u3_u2_n153 ) , .ZN( u0_u3_u2_n164 ) );
  NOR4_X1 u0_u3_u2_U5 (.A4( u0_u3_u2_n124 ) , .A3( u0_u3_u2_n125 ) , .A2( u0_u3_u2_n126 ) , .A1( u0_u3_u2_n127 ) , .ZN( u0_u3_u2_n128 ) );
  NAND2_X1 u0_u3_u2_U50 (.A2( u0_u3_u2_n100 ) , .A1( u0_u3_u2_n107 ) , .ZN( u0_u3_u2_n155 ) );
  NAND2_X1 u0_u3_u2_U51 (.A2( u0_u3_u2_n105 ) , .A1( u0_u3_u2_n108 ) , .ZN( u0_u3_u2_n143 ) );
  NAND2_X1 u0_u3_u2_U52 (.A1( u0_u3_u2_n104 ) , .A2( u0_u3_u2_n106 ) , .ZN( u0_u3_u2_n152 ) );
  NAND2_X1 u0_u3_u2_U53 (.A1( u0_u3_u2_n100 ) , .A2( u0_u3_u2_n105 ) , .ZN( u0_u3_u2_n132 ) );
  INV_X1 u0_u3_u2_U54 (.A( u0_u3_u2_n140 ) , .ZN( u0_u3_u2_n168 ) );
  INV_X1 u0_u3_u2_U55 (.A( u0_u3_u2_n138 ) , .ZN( u0_u3_u2_n167 ) );
  INV_X1 u0_u3_u2_U56 (.ZN( u0_u3_u2_n187 ) , .A( u0_u3_u2_n99 ) );
  OAI21_X1 u0_u3_u2_U57 (.B1( u0_u3_u2_n137 ) , .B2( u0_u3_u2_n143 ) , .A( u0_u3_u2_n98 ) , .ZN( u0_u3_u2_n99 ) );
  NAND2_X1 u0_u3_u2_U58 (.A1( u0_u3_u2_n102 ) , .A2( u0_u3_u2_n106 ) , .ZN( u0_u3_u2_n113 ) );
  NAND2_X1 u0_u3_u2_U59 (.A1( u0_u3_u2_n106 ) , .A2( u0_u3_u2_n107 ) , .ZN( u0_u3_u2_n131 ) );
  AOI21_X1 u0_u3_u2_U6 (.B2( u0_u3_u2_n119 ) , .ZN( u0_u3_u2_n127 ) , .A( u0_u3_u2_n137 ) , .B1( u0_u3_u2_n155 ) );
  NAND2_X1 u0_u3_u2_U60 (.A1( u0_u3_u2_n103 ) , .A2( u0_u3_u2_n107 ) , .ZN( u0_u3_u2_n139 ) );
  NAND2_X1 u0_u3_u2_U61 (.A1( u0_u3_u2_n103 ) , .A2( u0_u3_u2_n105 ) , .ZN( u0_u3_u2_n133 ) );
  NAND2_X1 u0_u3_u2_U62 (.A1( u0_u3_u2_n102 ) , .A2( u0_u3_u2_n103 ) , .ZN( u0_u3_u2_n154 ) );
  NAND2_X1 u0_u3_u2_U63 (.A2( u0_u3_u2_n103 ) , .A1( u0_u3_u2_n104 ) , .ZN( u0_u3_u2_n119 ) );
  NAND2_X1 u0_u3_u2_U64 (.A2( u0_u3_u2_n107 ) , .A1( u0_u3_u2_n108 ) , .ZN( u0_u3_u2_n123 ) );
  NAND2_X1 u0_u3_u2_U65 (.A1( u0_u3_u2_n104 ) , .A2( u0_u3_u2_n108 ) , .ZN( u0_u3_u2_n122 ) );
  INV_X1 u0_u3_u2_U66 (.A( u0_u3_u2_n114 ) , .ZN( u0_u3_u2_n172 ) );
  NAND2_X1 u0_u3_u2_U67 (.A2( u0_u3_u2_n100 ) , .A1( u0_u3_u2_n102 ) , .ZN( u0_u3_u2_n116 ) );
  NAND2_X1 u0_u3_u2_U68 (.A1( u0_u3_u2_n102 ) , .A2( u0_u3_u2_n108 ) , .ZN( u0_u3_u2_n120 ) );
  NAND2_X1 u0_u3_u2_U69 (.A2( u0_u3_u2_n105 ) , .A1( u0_u3_u2_n106 ) , .ZN( u0_u3_u2_n117 ) );
  AOI21_X1 u0_u3_u2_U7 (.ZN( u0_u3_u2_n124 ) , .B1( u0_u3_u2_n131 ) , .B2( u0_u3_u2_n143 ) , .A( u0_u3_u2_n172 ) );
  NOR2_X1 u0_u3_u2_U70 (.A2( u0_u3_X_16 ) , .ZN( u0_u3_u2_n140 ) , .A1( u0_u3_u2_n166 ) );
  NOR2_X1 u0_u3_u2_U71 (.A2( u0_u3_X_13 ) , .A1( u0_u3_X_14 ) , .ZN( u0_u3_u2_n100 ) );
  NOR2_X1 u0_u3_u2_U72 (.A2( u0_u3_X_16 ) , .A1( u0_u3_X_17 ) , .ZN( u0_u3_u2_n138 ) );
  NOR2_X1 u0_u3_u2_U73 (.A2( u0_u3_X_15 ) , .A1( u0_u3_X_18 ) , .ZN( u0_u3_u2_n104 ) );
  NOR2_X1 u0_u3_u2_U74 (.A2( u0_u3_X_14 ) , .ZN( u0_u3_u2_n103 ) , .A1( u0_u3_u2_n174 ) );
  NOR2_X1 u0_u3_u2_U75 (.A2( u0_u3_X_15 ) , .ZN( u0_u3_u2_n102 ) , .A1( u0_u3_u2_n165 ) );
  NOR2_X1 u0_u3_u2_U76 (.A2( u0_u3_X_17 ) , .ZN( u0_u3_u2_n114 ) , .A1( u0_u3_u2_n169 ) );
  AND2_X1 u0_u3_u2_U77 (.A1( u0_u3_X_15 ) , .ZN( u0_u3_u2_n105 ) , .A2( u0_u3_u2_n165 ) );
  AND2_X1 u0_u3_u2_U78 (.A2( u0_u3_X_15 ) , .A1( u0_u3_X_18 ) , .ZN( u0_u3_u2_n107 ) );
  AND2_X1 u0_u3_u2_U79 (.A1( u0_u3_X_14 ) , .ZN( u0_u3_u2_n106 ) , .A2( u0_u3_u2_n174 ) );
  AOI21_X1 u0_u3_u2_U8 (.B2( u0_u3_u2_n120 ) , .B1( u0_u3_u2_n121 ) , .ZN( u0_u3_u2_n126 ) , .A( u0_u3_u2_n167 ) );
  AND2_X1 u0_u3_u2_U80 (.A1( u0_u3_X_13 ) , .A2( u0_u3_X_14 ) , .ZN( u0_u3_u2_n108 ) );
  INV_X1 u0_u3_u2_U81 (.A( u0_u3_X_16 ) , .ZN( u0_u3_u2_n169 ) );
  INV_X1 u0_u3_u2_U82 (.A( u0_u3_X_17 ) , .ZN( u0_u3_u2_n166 ) );
  INV_X1 u0_u3_u2_U83 (.A( u0_u3_X_13 ) , .ZN( u0_u3_u2_n174 ) );
  INV_X1 u0_u3_u2_U84 (.A( u0_u3_X_18 ) , .ZN( u0_u3_u2_n165 ) );
  NAND4_X1 u0_u3_u2_U85 (.ZN( u0_out3_24 ) , .A4( u0_u3_u2_n111 ) , .A3( u0_u3_u2_n112 ) , .A1( u0_u3_u2_n130 ) , .A2( u0_u3_u2_n187 ) );
  AOI221_X1 u0_u3_u2_U86 (.A( u0_u3_u2_n109 ) , .B1( u0_u3_u2_n110 ) , .ZN( u0_u3_u2_n111 ) , .C1( u0_u3_u2_n134 ) , .C2( u0_u3_u2_n170 ) , .B2( u0_u3_u2_n173 ) );
  AOI21_X1 u0_u3_u2_U87 (.ZN( u0_u3_u2_n112 ) , .B2( u0_u3_u2_n156 ) , .A( u0_u3_u2_n164 ) , .B1( u0_u3_u2_n181 ) );
  NAND4_X1 u0_u3_u2_U88 (.ZN( u0_out3_16 ) , .A4( u0_u3_u2_n128 ) , .A3( u0_u3_u2_n129 ) , .A1( u0_u3_u2_n130 ) , .A2( u0_u3_u2_n186 ) );
  AOI22_X1 u0_u3_u2_U89 (.A2( u0_u3_u2_n118 ) , .ZN( u0_u3_u2_n129 ) , .A1( u0_u3_u2_n140 ) , .B1( u0_u3_u2_n157 ) , .B2( u0_u3_u2_n170 ) );
  OAI22_X1 u0_u3_u2_U9 (.ZN( u0_u3_u2_n109 ) , .A2( u0_u3_u2_n113 ) , .B2( u0_u3_u2_n133 ) , .B1( u0_u3_u2_n167 ) , .A1( u0_u3_u2_n168 ) );
  INV_X1 u0_u3_u2_U90 (.A( u0_u3_u2_n163 ) , .ZN( u0_u3_u2_n186 ) );
  NAND4_X1 u0_u3_u2_U91 (.ZN( u0_out3_30 ) , .A4( u0_u3_u2_n147 ) , .A3( u0_u3_u2_n148 ) , .A2( u0_u3_u2_n149 ) , .A1( u0_u3_u2_n187 ) );
  AOI21_X1 u0_u3_u2_U92 (.B2( u0_u3_u2_n138 ) , .ZN( u0_u3_u2_n148 ) , .A( u0_u3_u2_n162 ) , .B1( u0_u3_u2_n182 ) );
  NOR3_X1 u0_u3_u2_U93 (.A3( u0_u3_u2_n144 ) , .A2( u0_u3_u2_n145 ) , .A1( u0_u3_u2_n146 ) , .ZN( u0_u3_u2_n147 ) );
  OR4_X1 u0_u3_u2_U94 (.ZN( u0_out3_6 ) , .A4( u0_u3_u2_n161 ) , .A3( u0_u3_u2_n162 ) , .A2( u0_u3_u2_n163 ) , .A1( u0_u3_u2_n164 ) );
  OR3_X1 u0_u3_u2_U95 (.A2( u0_u3_u2_n159 ) , .A1( u0_u3_u2_n160 ) , .ZN( u0_u3_u2_n161 ) , .A3( u0_u3_u2_n183 ) );
  AOI21_X1 u0_u3_u2_U96 (.B2( u0_u3_u2_n154 ) , .B1( u0_u3_u2_n155 ) , .ZN( u0_u3_u2_n159 ) , .A( u0_u3_u2_n167 ) );
  NAND3_X1 u0_u3_u2_U97 (.A2( u0_u3_u2_n117 ) , .A1( u0_u3_u2_n122 ) , .A3( u0_u3_u2_n123 ) , .ZN( u0_u3_u2_n134 ) );
  NAND3_X1 u0_u3_u2_U98 (.ZN( u0_u3_u2_n110 ) , .A2( u0_u3_u2_n131 ) , .A3( u0_u3_u2_n139 ) , .A1( u0_u3_u2_n154 ) );
  NAND3_X1 u0_u3_u2_U99 (.A2( u0_u3_u2_n100 ) , .ZN( u0_u3_u2_n101 ) , .A1( u0_u3_u2_n104 ) , .A3( u0_u3_u2_n114 ) );
  XOR2_X1 u0_u5_U32 (.B( u0_K6_25 ) , .A( u0_R4_16 ) , .Z( u0_u5_X_25 ) );
  XOR2_X1 u0_u5_U34 (.B( u0_K6_23 ) , .A( u0_R4_16 ) , .Z( u0_u5_X_23 ) );
  XOR2_X1 u0_u5_U36 (.B( u0_K6_21 ) , .A( u0_R4_14 ) , .Z( u0_u5_X_21 ) );
  XOR2_X1 u0_u5_U37 (.B( u0_K6_20 ) , .A( u0_R4_13 ) , .Z( u0_u5_X_20 ) );
  XOR2_X1 u0_u5_U40 (.B( u0_K6_18 ) , .A( u0_R4_13 ) , .Z( u0_u5_X_18 ) );
  XOR2_X1 u0_u5_U45 (.B( u0_K6_13 ) , .A( u0_R4_8 ) , .Z( u0_u5_X_13 ) );
  XOR2_X1 u0_u5_U47 (.B( u0_K6_11 ) , .A( u0_R4_8 ) , .Z( u0_u5_X_11 ) );
  NOR2_X1 u0_u5_u1_U10 (.A1( u0_u5_u1_n112 ) , .A2( u0_u5_u1_n116 ) , .ZN( u0_u5_u1_n118 ) );
  NAND3_X1 u0_u5_u1_U100 (.ZN( u0_u5_u1_n113 ) , .A1( u0_u5_u1_n120 ) , .A3( u0_u5_u1_n133 ) , .A2( u0_u5_u1_n155 ) );
  OAI21_X1 u0_u5_u1_U11 (.ZN( u0_u5_u1_n101 ) , .B1( u0_u5_u1_n141 ) , .A( u0_u5_u1_n146 ) , .B2( u0_u5_u1_n183 ) );
  AOI21_X1 u0_u5_u1_U12 (.B2( u0_u5_u1_n155 ) , .B1( u0_u5_u1_n156 ) , .ZN( u0_u5_u1_n157 ) , .A( u0_u5_u1_n174 ) );
  NAND2_X1 u0_u5_u1_U13 (.ZN( u0_u5_u1_n140 ) , .A2( u0_u5_u1_n150 ) , .A1( u0_u5_u1_n155 ) );
  NAND2_X1 u0_u5_u1_U14 (.A1( u0_u5_u1_n131 ) , .ZN( u0_u5_u1_n147 ) , .A2( u0_u5_u1_n153 ) );
  INV_X1 u0_u5_u1_U15 (.A( u0_u5_u1_n139 ) , .ZN( u0_u5_u1_n174 ) );
  OR4_X1 u0_u5_u1_U16 (.A4( u0_u5_u1_n106 ) , .A3( u0_u5_u1_n107 ) , .ZN( u0_u5_u1_n108 ) , .A1( u0_u5_u1_n117 ) , .A2( u0_u5_u1_n184 ) );
  AOI21_X1 u0_u5_u1_U17 (.ZN( u0_u5_u1_n106 ) , .A( u0_u5_u1_n112 ) , .B1( u0_u5_u1_n154 ) , .B2( u0_u5_u1_n156 ) );
  INV_X1 u0_u5_u1_U18 (.A( u0_u5_u1_n101 ) , .ZN( u0_u5_u1_n184 ) );
  AOI21_X1 u0_u5_u1_U19 (.ZN( u0_u5_u1_n107 ) , .B1( u0_u5_u1_n134 ) , .B2( u0_u5_u1_n149 ) , .A( u0_u5_u1_n174 ) );
  INV_X1 u0_u5_u1_U20 (.A( u0_u5_u1_n112 ) , .ZN( u0_u5_u1_n171 ) );
  NAND2_X1 u0_u5_u1_U21 (.ZN( u0_u5_u1_n141 ) , .A1( u0_u5_u1_n153 ) , .A2( u0_u5_u1_n156 ) );
  AND2_X1 u0_u5_u1_U22 (.A1( u0_u5_u1_n123 ) , .ZN( u0_u5_u1_n134 ) , .A2( u0_u5_u1_n161 ) );
  NAND2_X1 u0_u5_u1_U23 (.A2( u0_u5_u1_n115 ) , .A1( u0_u5_u1_n116 ) , .ZN( u0_u5_u1_n148 ) );
  NAND2_X1 u0_u5_u1_U24 (.A2( u0_u5_u1_n133 ) , .A1( u0_u5_u1_n135 ) , .ZN( u0_u5_u1_n159 ) );
  NAND2_X1 u0_u5_u1_U25 (.A2( u0_u5_u1_n115 ) , .A1( u0_u5_u1_n120 ) , .ZN( u0_u5_u1_n132 ) );
  INV_X1 u0_u5_u1_U26 (.A( u0_u5_u1_n154 ) , .ZN( u0_u5_u1_n178 ) );
  INV_X1 u0_u5_u1_U27 (.A( u0_u5_u1_n151 ) , .ZN( u0_u5_u1_n183 ) );
  AND2_X1 u0_u5_u1_U28 (.A1( u0_u5_u1_n129 ) , .A2( u0_u5_u1_n133 ) , .ZN( u0_u5_u1_n149 ) );
  INV_X1 u0_u5_u1_U29 (.A( u0_u5_u1_n131 ) , .ZN( u0_u5_u1_n180 ) );
  INV_X1 u0_u5_u1_U3 (.A( u0_u5_u1_n159 ) , .ZN( u0_u5_u1_n182 ) );
  OAI221_X1 u0_u5_u1_U30 (.A( u0_u5_u1_n119 ) , .C2( u0_u5_u1_n129 ) , .ZN( u0_u5_u1_n138 ) , .B2( u0_u5_u1_n152 ) , .C1( u0_u5_u1_n174 ) , .B1( u0_u5_u1_n187 ) );
  INV_X1 u0_u5_u1_U31 (.A( u0_u5_u1_n148 ) , .ZN( u0_u5_u1_n187 ) );
  AOI211_X1 u0_u5_u1_U32 (.B( u0_u5_u1_n117 ) , .A( u0_u5_u1_n118 ) , .ZN( u0_u5_u1_n119 ) , .C2( u0_u5_u1_n146 ) , .C1( u0_u5_u1_n159 ) );
  NOR2_X1 u0_u5_u1_U33 (.A1( u0_u5_u1_n168 ) , .A2( u0_u5_u1_n176 ) , .ZN( u0_u5_u1_n98 ) );
  OAI21_X1 u0_u5_u1_U34 (.B2( u0_u5_u1_n123 ) , .ZN( u0_u5_u1_n145 ) , .B1( u0_u5_u1_n160 ) , .A( u0_u5_u1_n185 ) );
  INV_X1 u0_u5_u1_U35 (.A( u0_u5_u1_n122 ) , .ZN( u0_u5_u1_n185 ) );
  AOI21_X1 u0_u5_u1_U36 (.B2( u0_u5_u1_n120 ) , .B1( u0_u5_u1_n121 ) , .ZN( u0_u5_u1_n122 ) , .A( u0_u5_u1_n128 ) );
  NAND2_X1 u0_u5_u1_U37 (.A1( u0_u5_u1_n128 ) , .ZN( u0_u5_u1_n146 ) , .A2( u0_u5_u1_n160 ) );
  NAND2_X1 u0_u5_u1_U38 (.A2( u0_u5_u1_n112 ) , .ZN( u0_u5_u1_n139 ) , .A1( u0_u5_u1_n152 ) );
  NAND2_X1 u0_u5_u1_U39 (.A1( u0_u5_u1_n105 ) , .ZN( u0_u5_u1_n156 ) , .A2( u0_u5_u1_n99 ) );
  AOI221_X1 u0_u5_u1_U4 (.A( u0_u5_u1_n138 ) , .C2( u0_u5_u1_n139 ) , .C1( u0_u5_u1_n140 ) , .B2( u0_u5_u1_n141 ) , .ZN( u0_u5_u1_n142 ) , .B1( u0_u5_u1_n175 ) );
  AOI221_X1 u0_u5_u1_U40 (.B1( u0_u5_u1_n140 ) , .ZN( u0_u5_u1_n167 ) , .B2( u0_u5_u1_n172 ) , .C2( u0_u5_u1_n175 ) , .C1( u0_u5_u1_n178 ) , .A( u0_u5_u1_n188 ) );
  INV_X1 u0_u5_u1_U41 (.ZN( u0_u5_u1_n188 ) , .A( u0_u5_u1_n97 ) );
  AOI211_X1 u0_u5_u1_U42 (.A( u0_u5_u1_n118 ) , .C1( u0_u5_u1_n132 ) , .C2( u0_u5_u1_n139 ) , .B( u0_u5_u1_n96 ) , .ZN( u0_u5_u1_n97 ) );
  AOI21_X1 u0_u5_u1_U43 (.B2( u0_u5_u1_n121 ) , .B1( u0_u5_u1_n135 ) , .A( u0_u5_u1_n152 ) , .ZN( u0_u5_u1_n96 ) );
  NOR2_X1 u0_u5_u1_U44 (.ZN( u0_u5_u1_n117 ) , .A1( u0_u5_u1_n121 ) , .A2( u0_u5_u1_n160 ) );
  AOI21_X1 u0_u5_u1_U45 (.A( u0_u5_u1_n128 ) , .B2( u0_u5_u1_n129 ) , .ZN( u0_u5_u1_n130 ) , .B1( u0_u5_u1_n150 ) );
  NAND2_X1 u0_u5_u1_U46 (.ZN( u0_u5_u1_n112 ) , .A1( u0_u5_u1_n169 ) , .A2( u0_u5_u1_n170 ) );
  NAND2_X1 u0_u5_u1_U47 (.ZN( u0_u5_u1_n129 ) , .A2( u0_u5_u1_n95 ) , .A1( u0_u5_u1_n98 ) );
  NAND2_X1 u0_u5_u1_U48 (.A1( u0_u5_u1_n102 ) , .ZN( u0_u5_u1_n154 ) , .A2( u0_u5_u1_n99 ) );
  NAND2_X1 u0_u5_u1_U49 (.A2( u0_u5_u1_n100 ) , .ZN( u0_u5_u1_n135 ) , .A1( u0_u5_u1_n99 ) );
  AOI211_X1 u0_u5_u1_U5 (.ZN( u0_u5_u1_n124 ) , .A( u0_u5_u1_n138 ) , .C2( u0_u5_u1_n139 ) , .B( u0_u5_u1_n145 ) , .C1( u0_u5_u1_n147 ) );
  AOI21_X1 u0_u5_u1_U50 (.A( u0_u5_u1_n152 ) , .B2( u0_u5_u1_n153 ) , .B1( u0_u5_u1_n154 ) , .ZN( u0_u5_u1_n158 ) );
  INV_X1 u0_u5_u1_U51 (.A( u0_u5_u1_n160 ) , .ZN( u0_u5_u1_n175 ) );
  NAND2_X1 u0_u5_u1_U52 (.A1( u0_u5_u1_n100 ) , .ZN( u0_u5_u1_n116 ) , .A2( u0_u5_u1_n95 ) );
  NAND2_X1 u0_u5_u1_U53 (.A1( u0_u5_u1_n102 ) , .ZN( u0_u5_u1_n131 ) , .A2( u0_u5_u1_n95 ) );
  NAND2_X1 u0_u5_u1_U54 (.A2( u0_u5_u1_n104 ) , .ZN( u0_u5_u1_n121 ) , .A1( u0_u5_u1_n98 ) );
  NAND2_X1 u0_u5_u1_U55 (.A1( u0_u5_u1_n103 ) , .ZN( u0_u5_u1_n153 ) , .A2( u0_u5_u1_n98 ) );
  NAND2_X1 u0_u5_u1_U56 (.A2( u0_u5_u1_n104 ) , .A1( u0_u5_u1_n105 ) , .ZN( u0_u5_u1_n133 ) );
  NAND2_X1 u0_u5_u1_U57 (.ZN( u0_u5_u1_n150 ) , .A2( u0_u5_u1_n98 ) , .A1( u0_u5_u1_n99 ) );
  NAND2_X1 u0_u5_u1_U58 (.A1( u0_u5_u1_n105 ) , .ZN( u0_u5_u1_n155 ) , .A2( u0_u5_u1_n95 ) );
  OAI21_X1 u0_u5_u1_U59 (.ZN( u0_u5_u1_n109 ) , .B1( u0_u5_u1_n129 ) , .B2( u0_u5_u1_n160 ) , .A( u0_u5_u1_n167 ) );
  AOI22_X1 u0_u5_u1_U6 (.B2( u0_u5_u1_n136 ) , .A2( u0_u5_u1_n137 ) , .ZN( u0_u5_u1_n143 ) , .A1( u0_u5_u1_n171 ) , .B1( u0_u5_u1_n173 ) );
  NAND2_X1 u0_u5_u1_U60 (.A2( u0_u5_u1_n100 ) , .A1( u0_u5_u1_n103 ) , .ZN( u0_u5_u1_n120 ) );
  NAND2_X1 u0_u5_u1_U61 (.A1( u0_u5_u1_n102 ) , .A2( u0_u5_u1_n104 ) , .ZN( u0_u5_u1_n115 ) );
  NAND2_X1 u0_u5_u1_U62 (.A2( u0_u5_u1_n100 ) , .A1( u0_u5_u1_n104 ) , .ZN( u0_u5_u1_n151 ) );
  NAND2_X1 u0_u5_u1_U63 (.A2( u0_u5_u1_n103 ) , .A1( u0_u5_u1_n105 ) , .ZN( u0_u5_u1_n161 ) );
  INV_X1 u0_u5_u1_U64 (.A( u0_u5_u1_n152 ) , .ZN( u0_u5_u1_n173 ) );
  INV_X1 u0_u5_u1_U65 (.A( u0_u5_u1_n128 ) , .ZN( u0_u5_u1_n172 ) );
  NAND2_X1 u0_u5_u1_U66 (.A2( u0_u5_u1_n102 ) , .A1( u0_u5_u1_n103 ) , .ZN( u0_u5_u1_n123 ) );
  AOI211_X1 u0_u5_u1_U67 (.B( u0_u5_u1_n162 ) , .A( u0_u5_u1_n163 ) , .C2( u0_u5_u1_n164 ) , .ZN( u0_u5_u1_n165 ) , .C1( u0_u5_u1_n171 ) );
  AOI21_X1 u0_u5_u1_U68 (.A( u0_u5_u1_n160 ) , .B2( u0_u5_u1_n161 ) , .ZN( u0_u5_u1_n162 ) , .B1( u0_u5_u1_n182 ) );
  OR2_X1 u0_u5_u1_U69 (.A2( u0_u5_u1_n157 ) , .A1( u0_u5_u1_n158 ) , .ZN( u0_u5_u1_n163 ) );
  INV_X1 u0_u5_u1_U7 (.A( u0_u5_u1_n147 ) , .ZN( u0_u5_u1_n181 ) );
  NOR2_X1 u0_u5_u1_U70 (.A2( u0_u5_X_7 ) , .A1( u0_u5_X_8 ) , .ZN( u0_u5_u1_n95 ) );
  NOR2_X1 u0_u5_u1_U71 (.A1( u0_u5_X_12 ) , .A2( u0_u5_X_9 ) , .ZN( u0_u5_u1_n100 ) );
  NOR2_X1 u0_u5_u1_U72 (.A2( u0_u5_X_8 ) , .A1( u0_u5_u1_n177 ) , .ZN( u0_u5_u1_n99 ) );
  NOR2_X1 u0_u5_u1_U73 (.A2( u0_u5_X_12 ) , .ZN( u0_u5_u1_n102 ) , .A1( u0_u5_u1_n176 ) );
  NOR2_X1 u0_u5_u1_U74 (.A2( u0_u5_X_9 ) , .ZN( u0_u5_u1_n105 ) , .A1( u0_u5_u1_n168 ) );
  NAND2_X1 u0_u5_u1_U75 (.A1( u0_u5_X_10 ) , .ZN( u0_u5_u1_n160 ) , .A2( u0_u5_u1_n169 ) );
  NAND2_X1 u0_u5_u1_U76 (.A2( u0_u5_X_10 ) , .A1( u0_u5_X_11 ) , .ZN( u0_u5_u1_n152 ) );
  NAND2_X1 u0_u5_u1_U77 (.A1( u0_u5_X_11 ) , .ZN( u0_u5_u1_n128 ) , .A2( u0_u5_u1_n170 ) );
  AND2_X1 u0_u5_u1_U78 (.A2( u0_u5_X_7 ) , .A1( u0_u5_X_8 ) , .ZN( u0_u5_u1_n104 ) );
  AND2_X1 u0_u5_u1_U79 (.A1( u0_u5_X_8 ) , .ZN( u0_u5_u1_n103 ) , .A2( u0_u5_u1_n177 ) );
  AOI22_X1 u0_u5_u1_U8 (.B2( u0_u5_u1_n113 ) , .A2( u0_u5_u1_n114 ) , .ZN( u0_u5_u1_n125 ) , .A1( u0_u5_u1_n171 ) , .B1( u0_u5_u1_n173 ) );
  INV_X1 u0_u5_u1_U80 (.A( u0_u5_X_10 ) , .ZN( u0_u5_u1_n170 ) );
  INV_X1 u0_u5_u1_U81 (.A( u0_u5_X_9 ) , .ZN( u0_u5_u1_n176 ) );
  INV_X1 u0_u5_u1_U82 (.A( u0_u5_X_11 ) , .ZN( u0_u5_u1_n169 ) );
  INV_X1 u0_u5_u1_U83 (.A( u0_u5_X_12 ) , .ZN( u0_u5_u1_n168 ) );
  INV_X1 u0_u5_u1_U84 (.A( u0_u5_X_7 ) , .ZN( u0_u5_u1_n177 ) );
  NAND4_X1 u0_u5_u1_U85 (.ZN( u0_out5_28 ) , .A4( u0_u5_u1_n124 ) , .A3( u0_u5_u1_n125 ) , .A2( u0_u5_u1_n126 ) , .A1( u0_u5_u1_n127 ) );
  OAI21_X1 u0_u5_u1_U86 (.ZN( u0_u5_u1_n127 ) , .B2( u0_u5_u1_n139 ) , .B1( u0_u5_u1_n175 ) , .A( u0_u5_u1_n183 ) );
  OAI21_X1 u0_u5_u1_U87 (.ZN( u0_u5_u1_n126 ) , .B2( u0_u5_u1_n140 ) , .A( u0_u5_u1_n146 ) , .B1( u0_u5_u1_n178 ) );
  NAND4_X1 u0_u5_u1_U88 (.ZN( u0_out5_18 ) , .A4( u0_u5_u1_n165 ) , .A3( u0_u5_u1_n166 ) , .A1( u0_u5_u1_n167 ) , .A2( u0_u5_u1_n186 ) );
  AOI22_X1 u0_u5_u1_U89 (.B2( u0_u5_u1_n146 ) , .B1( u0_u5_u1_n147 ) , .A2( u0_u5_u1_n148 ) , .ZN( u0_u5_u1_n166 ) , .A1( u0_u5_u1_n172 ) );
  NAND2_X1 u0_u5_u1_U9 (.ZN( u0_u5_u1_n114 ) , .A1( u0_u5_u1_n134 ) , .A2( u0_u5_u1_n156 ) );
  INV_X1 u0_u5_u1_U90 (.A( u0_u5_u1_n145 ) , .ZN( u0_u5_u1_n186 ) );
  NAND4_X1 u0_u5_u1_U91 (.ZN( u0_out5_2 ) , .A4( u0_u5_u1_n142 ) , .A3( u0_u5_u1_n143 ) , .A2( u0_u5_u1_n144 ) , .A1( u0_u5_u1_n179 ) );
  OAI21_X1 u0_u5_u1_U92 (.B2( u0_u5_u1_n132 ) , .ZN( u0_u5_u1_n144 ) , .A( u0_u5_u1_n146 ) , .B1( u0_u5_u1_n180 ) );
  INV_X1 u0_u5_u1_U93 (.A( u0_u5_u1_n130 ) , .ZN( u0_u5_u1_n179 ) );
  OR4_X1 u0_u5_u1_U94 (.ZN( u0_out5_13 ) , .A4( u0_u5_u1_n108 ) , .A3( u0_u5_u1_n109 ) , .A2( u0_u5_u1_n110 ) , .A1( u0_u5_u1_n111 ) );
  AOI21_X1 u0_u5_u1_U95 (.ZN( u0_u5_u1_n110 ) , .A( u0_u5_u1_n116 ) , .B1( u0_u5_u1_n152 ) , .B2( u0_u5_u1_n160 ) );
  AOI21_X1 u0_u5_u1_U96 (.ZN( u0_u5_u1_n111 ) , .A( u0_u5_u1_n128 ) , .B2( u0_u5_u1_n131 ) , .B1( u0_u5_u1_n135 ) );
  NAND3_X1 u0_u5_u1_U97 (.A3( u0_u5_u1_n149 ) , .A2( u0_u5_u1_n150 ) , .A1( u0_u5_u1_n151 ) , .ZN( u0_u5_u1_n164 ) );
  NAND3_X1 u0_u5_u1_U98 (.A3( u0_u5_u1_n134 ) , .A2( u0_u5_u1_n135 ) , .ZN( u0_u5_u1_n136 ) , .A1( u0_u5_u1_n151 ) );
  NAND3_X1 u0_u5_u1_U99 (.A1( u0_u5_u1_n133 ) , .ZN( u0_u5_u1_n137 ) , .A2( u0_u5_u1_n154 ) , .A3( u0_u5_u1_n181 ) );
  OAI22_X1 u0_u5_u2_U10 (.ZN( u0_u5_u2_n109 ) , .A2( u0_u5_u2_n113 ) , .B2( u0_u5_u2_n133 ) , .B1( u0_u5_u2_n167 ) , .A1( u0_u5_u2_n168 ) );
  NAND3_X1 u0_u5_u2_U100 (.A2( u0_u5_u2_n100 ) , .A1( u0_u5_u2_n104 ) , .A3( u0_u5_u2_n138 ) , .ZN( u0_u5_u2_n98 ) );
  OAI22_X1 u0_u5_u2_U11 (.B1( u0_u5_u2_n151 ) , .A2( u0_u5_u2_n152 ) , .A1( u0_u5_u2_n153 ) , .ZN( u0_u5_u2_n160 ) , .B2( u0_u5_u2_n168 ) );
  NOR3_X1 u0_u5_u2_U12 (.A1( u0_u5_u2_n150 ) , .ZN( u0_u5_u2_n151 ) , .A3( u0_u5_u2_n175 ) , .A2( u0_u5_u2_n188 ) );
  AOI21_X1 u0_u5_u2_U13 (.ZN( u0_u5_u2_n144 ) , .B2( u0_u5_u2_n155 ) , .A( u0_u5_u2_n172 ) , .B1( u0_u5_u2_n185 ) );
  AOI21_X1 u0_u5_u2_U14 (.B2( u0_u5_u2_n143 ) , .ZN( u0_u5_u2_n145 ) , .B1( u0_u5_u2_n152 ) , .A( u0_u5_u2_n171 ) );
  AOI21_X1 u0_u5_u2_U15 (.B2( u0_u5_u2_n120 ) , .B1( u0_u5_u2_n121 ) , .ZN( u0_u5_u2_n126 ) , .A( u0_u5_u2_n167 ) );
  INV_X1 u0_u5_u2_U16 (.A( u0_u5_u2_n156 ) , .ZN( u0_u5_u2_n171 ) );
  INV_X1 u0_u5_u2_U17 (.A( u0_u5_u2_n120 ) , .ZN( u0_u5_u2_n188 ) );
  NAND2_X1 u0_u5_u2_U18 (.A2( u0_u5_u2_n122 ) , .ZN( u0_u5_u2_n150 ) , .A1( u0_u5_u2_n152 ) );
  INV_X1 u0_u5_u2_U19 (.A( u0_u5_u2_n153 ) , .ZN( u0_u5_u2_n170 ) );
  INV_X1 u0_u5_u2_U20 (.A( u0_u5_u2_n137 ) , .ZN( u0_u5_u2_n173 ) );
  NAND2_X1 u0_u5_u2_U21 (.A1( u0_u5_u2_n132 ) , .A2( u0_u5_u2_n139 ) , .ZN( u0_u5_u2_n157 ) );
  INV_X1 u0_u5_u2_U22 (.A( u0_u5_u2_n113 ) , .ZN( u0_u5_u2_n178 ) );
  INV_X1 u0_u5_u2_U23 (.A( u0_u5_u2_n139 ) , .ZN( u0_u5_u2_n175 ) );
  INV_X1 u0_u5_u2_U24 (.A( u0_u5_u2_n155 ) , .ZN( u0_u5_u2_n181 ) );
  INV_X1 u0_u5_u2_U25 (.A( u0_u5_u2_n119 ) , .ZN( u0_u5_u2_n177 ) );
  INV_X1 u0_u5_u2_U26 (.A( u0_u5_u2_n116 ) , .ZN( u0_u5_u2_n180 ) );
  INV_X1 u0_u5_u2_U27 (.A( u0_u5_u2_n131 ) , .ZN( u0_u5_u2_n179 ) );
  INV_X1 u0_u5_u2_U28 (.A( u0_u5_u2_n154 ) , .ZN( u0_u5_u2_n176 ) );
  NAND2_X1 u0_u5_u2_U29 (.A2( u0_u5_u2_n116 ) , .A1( u0_u5_u2_n117 ) , .ZN( u0_u5_u2_n118 ) );
  NOR2_X1 u0_u5_u2_U3 (.ZN( u0_u5_u2_n121 ) , .A2( u0_u5_u2_n177 ) , .A1( u0_u5_u2_n180 ) );
  INV_X1 u0_u5_u2_U30 (.A( u0_u5_u2_n132 ) , .ZN( u0_u5_u2_n182 ) );
  INV_X1 u0_u5_u2_U31 (.A( u0_u5_u2_n158 ) , .ZN( u0_u5_u2_n183 ) );
  OAI21_X1 u0_u5_u2_U32 (.A( u0_u5_u2_n156 ) , .B1( u0_u5_u2_n157 ) , .ZN( u0_u5_u2_n158 ) , .B2( u0_u5_u2_n179 ) );
  NOR2_X1 u0_u5_u2_U33 (.ZN( u0_u5_u2_n156 ) , .A1( u0_u5_u2_n166 ) , .A2( u0_u5_u2_n169 ) );
  NOR2_X1 u0_u5_u2_U34 (.A2( u0_u5_u2_n114 ) , .ZN( u0_u5_u2_n137 ) , .A1( u0_u5_u2_n140 ) );
  NOR2_X1 u0_u5_u2_U35 (.A2( u0_u5_u2_n138 ) , .ZN( u0_u5_u2_n153 ) , .A1( u0_u5_u2_n156 ) );
  AOI211_X1 u0_u5_u2_U36 (.ZN( u0_u5_u2_n130 ) , .C1( u0_u5_u2_n138 ) , .C2( u0_u5_u2_n179 ) , .B( u0_u5_u2_n96 ) , .A( u0_u5_u2_n97 ) );
  OAI22_X1 u0_u5_u2_U37 (.B1( u0_u5_u2_n133 ) , .A2( u0_u5_u2_n137 ) , .A1( u0_u5_u2_n152 ) , .B2( u0_u5_u2_n168 ) , .ZN( u0_u5_u2_n97 ) );
  OAI221_X1 u0_u5_u2_U38 (.B1( u0_u5_u2_n113 ) , .C1( u0_u5_u2_n132 ) , .A( u0_u5_u2_n149 ) , .B2( u0_u5_u2_n171 ) , .C2( u0_u5_u2_n172 ) , .ZN( u0_u5_u2_n96 ) );
  OAI221_X1 u0_u5_u2_U39 (.A( u0_u5_u2_n115 ) , .C2( u0_u5_u2_n123 ) , .B2( u0_u5_u2_n143 ) , .B1( u0_u5_u2_n153 ) , .ZN( u0_u5_u2_n163 ) , .C1( u0_u5_u2_n168 ) );
  INV_X1 u0_u5_u2_U4 (.A( u0_u5_u2_n134 ) , .ZN( u0_u5_u2_n185 ) );
  OAI21_X1 u0_u5_u2_U40 (.A( u0_u5_u2_n114 ) , .ZN( u0_u5_u2_n115 ) , .B1( u0_u5_u2_n176 ) , .B2( u0_u5_u2_n178 ) );
  OAI221_X1 u0_u5_u2_U41 (.A( u0_u5_u2_n135 ) , .B2( u0_u5_u2_n136 ) , .B1( u0_u5_u2_n137 ) , .ZN( u0_u5_u2_n162 ) , .C2( u0_u5_u2_n167 ) , .C1( u0_u5_u2_n185 ) );
  AND3_X1 u0_u5_u2_U42 (.A3( u0_u5_u2_n131 ) , .A2( u0_u5_u2_n132 ) , .A1( u0_u5_u2_n133 ) , .ZN( u0_u5_u2_n136 ) );
  AOI22_X1 u0_u5_u2_U43 (.ZN( u0_u5_u2_n135 ) , .B1( u0_u5_u2_n140 ) , .A1( u0_u5_u2_n156 ) , .B2( u0_u5_u2_n180 ) , .A2( u0_u5_u2_n188 ) );
  AOI21_X1 u0_u5_u2_U44 (.ZN( u0_u5_u2_n149 ) , .B1( u0_u5_u2_n173 ) , .B2( u0_u5_u2_n188 ) , .A( u0_u5_u2_n95 ) );
  AND3_X1 u0_u5_u2_U45 (.A2( u0_u5_u2_n100 ) , .A1( u0_u5_u2_n104 ) , .A3( u0_u5_u2_n156 ) , .ZN( u0_u5_u2_n95 ) );
  OAI21_X1 u0_u5_u2_U46 (.A( u0_u5_u2_n141 ) , .B2( u0_u5_u2_n142 ) , .ZN( u0_u5_u2_n146 ) , .B1( u0_u5_u2_n153 ) );
  OAI21_X1 u0_u5_u2_U47 (.A( u0_u5_u2_n140 ) , .ZN( u0_u5_u2_n141 ) , .B1( u0_u5_u2_n176 ) , .B2( u0_u5_u2_n177 ) );
  NOR3_X1 u0_u5_u2_U48 (.ZN( u0_u5_u2_n142 ) , .A3( u0_u5_u2_n175 ) , .A2( u0_u5_u2_n178 ) , .A1( u0_u5_u2_n181 ) );
  OAI21_X1 u0_u5_u2_U49 (.A( u0_u5_u2_n101 ) , .B2( u0_u5_u2_n121 ) , .B1( u0_u5_u2_n153 ) , .ZN( u0_u5_u2_n164 ) );
  INV_X1 u0_u5_u2_U5 (.A( u0_u5_u2_n150 ) , .ZN( u0_u5_u2_n184 ) );
  NAND2_X1 u0_u5_u2_U50 (.A2( u0_u5_u2_n100 ) , .A1( u0_u5_u2_n107 ) , .ZN( u0_u5_u2_n155 ) );
  NAND2_X1 u0_u5_u2_U51 (.A2( u0_u5_u2_n105 ) , .A1( u0_u5_u2_n108 ) , .ZN( u0_u5_u2_n143 ) );
  NAND2_X1 u0_u5_u2_U52 (.A1( u0_u5_u2_n104 ) , .A2( u0_u5_u2_n106 ) , .ZN( u0_u5_u2_n152 ) );
  NAND2_X1 u0_u5_u2_U53 (.A1( u0_u5_u2_n100 ) , .A2( u0_u5_u2_n105 ) , .ZN( u0_u5_u2_n132 ) );
  INV_X1 u0_u5_u2_U54 (.A( u0_u5_u2_n140 ) , .ZN( u0_u5_u2_n168 ) );
  INV_X1 u0_u5_u2_U55 (.A( u0_u5_u2_n138 ) , .ZN( u0_u5_u2_n167 ) );
  NAND2_X1 u0_u5_u2_U56 (.A1( u0_u5_u2_n102 ) , .A2( u0_u5_u2_n106 ) , .ZN( u0_u5_u2_n113 ) );
  NAND2_X1 u0_u5_u2_U57 (.A1( u0_u5_u2_n106 ) , .A2( u0_u5_u2_n107 ) , .ZN( u0_u5_u2_n131 ) );
  NAND2_X1 u0_u5_u2_U58 (.A1( u0_u5_u2_n103 ) , .A2( u0_u5_u2_n107 ) , .ZN( u0_u5_u2_n139 ) );
  NAND2_X1 u0_u5_u2_U59 (.A1( u0_u5_u2_n103 ) , .A2( u0_u5_u2_n105 ) , .ZN( u0_u5_u2_n133 ) );
  NOR4_X1 u0_u5_u2_U6 (.A4( u0_u5_u2_n124 ) , .A3( u0_u5_u2_n125 ) , .A2( u0_u5_u2_n126 ) , .A1( u0_u5_u2_n127 ) , .ZN( u0_u5_u2_n128 ) );
  NAND2_X1 u0_u5_u2_U60 (.A1( u0_u5_u2_n102 ) , .A2( u0_u5_u2_n103 ) , .ZN( u0_u5_u2_n154 ) );
  NAND2_X1 u0_u5_u2_U61 (.A2( u0_u5_u2_n103 ) , .A1( u0_u5_u2_n104 ) , .ZN( u0_u5_u2_n119 ) );
  NAND2_X1 u0_u5_u2_U62 (.A2( u0_u5_u2_n107 ) , .A1( u0_u5_u2_n108 ) , .ZN( u0_u5_u2_n123 ) );
  NAND2_X1 u0_u5_u2_U63 (.A1( u0_u5_u2_n104 ) , .A2( u0_u5_u2_n108 ) , .ZN( u0_u5_u2_n122 ) );
  INV_X1 u0_u5_u2_U64 (.A( u0_u5_u2_n114 ) , .ZN( u0_u5_u2_n172 ) );
  NAND2_X1 u0_u5_u2_U65 (.A2( u0_u5_u2_n100 ) , .A1( u0_u5_u2_n102 ) , .ZN( u0_u5_u2_n116 ) );
  NAND2_X1 u0_u5_u2_U66 (.A1( u0_u5_u2_n102 ) , .A2( u0_u5_u2_n108 ) , .ZN( u0_u5_u2_n120 ) );
  NAND2_X1 u0_u5_u2_U67 (.A2( u0_u5_u2_n105 ) , .A1( u0_u5_u2_n106 ) , .ZN( u0_u5_u2_n117 ) );
  INV_X1 u0_u5_u2_U68 (.ZN( u0_u5_u2_n187 ) , .A( u0_u5_u2_n99 ) );
  OAI21_X1 u0_u5_u2_U69 (.B1( u0_u5_u2_n137 ) , .B2( u0_u5_u2_n143 ) , .A( u0_u5_u2_n98 ) , .ZN( u0_u5_u2_n99 ) );
  AOI21_X1 u0_u5_u2_U7 (.B2( u0_u5_u2_n119 ) , .ZN( u0_u5_u2_n127 ) , .A( u0_u5_u2_n137 ) , .B1( u0_u5_u2_n155 ) );
  NOR2_X1 u0_u5_u2_U70 (.A2( u0_u5_X_16 ) , .ZN( u0_u5_u2_n140 ) , .A1( u0_u5_u2_n166 ) );
  NOR2_X1 u0_u5_u2_U71 (.A2( u0_u5_X_13 ) , .A1( u0_u5_X_14 ) , .ZN( u0_u5_u2_n100 ) );
  NOR2_X1 u0_u5_u2_U72 (.A2( u0_u5_X_16 ) , .A1( u0_u5_X_17 ) , .ZN( u0_u5_u2_n138 ) );
  NOR2_X1 u0_u5_u2_U73 (.A2( u0_u5_X_15 ) , .A1( u0_u5_X_18 ) , .ZN( u0_u5_u2_n104 ) );
  NOR2_X1 u0_u5_u2_U74 (.A2( u0_u5_X_14 ) , .ZN( u0_u5_u2_n103 ) , .A1( u0_u5_u2_n174 ) );
  NOR2_X1 u0_u5_u2_U75 (.A2( u0_u5_X_15 ) , .ZN( u0_u5_u2_n102 ) , .A1( u0_u5_u2_n165 ) );
  NOR2_X1 u0_u5_u2_U76 (.A2( u0_u5_X_17 ) , .ZN( u0_u5_u2_n114 ) , .A1( u0_u5_u2_n169 ) );
  AND2_X1 u0_u5_u2_U77 (.A1( u0_u5_X_15 ) , .ZN( u0_u5_u2_n105 ) , .A2( u0_u5_u2_n165 ) );
  AND2_X1 u0_u5_u2_U78 (.A2( u0_u5_X_15 ) , .A1( u0_u5_X_18 ) , .ZN( u0_u5_u2_n107 ) );
  AND2_X1 u0_u5_u2_U79 (.A1( u0_u5_X_14 ) , .ZN( u0_u5_u2_n106 ) , .A2( u0_u5_u2_n174 ) );
  AOI21_X1 u0_u5_u2_U8 (.ZN( u0_u5_u2_n124 ) , .B1( u0_u5_u2_n131 ) , .B2( u0_u5_u2_n143 ) , .A( u0_u5_u2_n172 ) );
  AND2_X1 u0_u5_u2_U80 (.A1( u0_u5_X_13 ) , .A2( u0_u5_X_14 ) , .ZN( u0_u5_u2_n108 ) );
  INV_X1 u0_u5_u2_U81 (.A( u0_u5_X_16 ) , .ZN( u0_u5_u2_n169 ) );
  INV_X1 u0_u5_u2_U82 (.A( u0_u5_X_17 ) , .ZN( u0_u5_u2_n166 ) );
  INV_X1 u0_u5_u2_U83 (.A( u0_u5_X_13 ) , .ZN( u0_u5_u2_n174 ) );
  INV_X1 u0_u5_u2_U84 (.A( u0_u5_X_18 ) , .ZN( u0_u5_u2_n165 ) );
  NAND4_X1 u0_u5_u2_U85 (.ZN( u0_out5_30 ) , .A4( u0_u5_u2_n147 ) , .A3( u0_u5_u2_n148 ) , .A2( u0_u5_u2_n149 ) , .A1( u0_u5_u2_n187 ) );
  NOR3_X1 u0_u5_u2_U86 (.A3( u0_u5_u2_n144 ) , .A2( u0_u5_u2_n145 ) , .A1( u0_u5_u2_n146 ) , .ZN( u0_u5_u2_n147 ) );
  AOI21_X1 u0_u5_u2_U87 (.B2( u0_u5_u2_n138 ) , .ZN( u0_u5_u2_n148 ) , .A( u0_u5_u2_n162 ) , .B1( u0_u5_u2_n182 ) );
  NAND4_X1 u0_u5_u2_U88 (.ZN( u0_out5_24 ) , .A4( u0_u5_u2_n111 ) , .A3( u0_u5_u2_n112 ) , .A1( u0_u5_u2_n130 ) , .A2( u0_u5_u2_n187 ) );
  AOI221_X1 u0_u5_u2_U89 (.A( u0_u5_u2_n109 ) , .B1( u0_u5_u2_n110 ) , .ZN( u0_u5_u2_n111 ) , .C1( u0_u5_u2_n134 ) , .C2( u0_u5_u2_n170 ) , .B2( u0_u5_u2_n173 ) );
  AOI21_X1 u0_u5_u2_U9 (.B2( u0_u5_u2_n123 ) , .ZN( u0_u5_u2_n125 ) , .A( u0_u5_u2_n171 ) , .B1( u0_u5_u2_n184 ) );
  AOI21_X1 u0_u5_u2_U90 (.ZN( u0_u5_u2_n112 ) , .B2( u0_u5_u2_n156 ) , .A( u0_u5_u2_n164 ) , .B1( u0_u5_u2_n181 ) );
  NAND4_X1 u0_u5_u2_U91 (.ZN( u0_out5_16 ) , .A4( u0_u5_u2_n128 ) , .A3( u0_u5_u2_n129 ) , .A1( u0_u5_u2_n130 ) , .A2( u0_u5_u2_n186 ) );
  AOI22_X1 u0_u5_u2_U92 (.A2( u0_u5_u2_n118 ) , .ZN( u0_u5_u2_n129 ) , .A1( u0_u5_u2_n140 ) , .B1( u0_u5_u2_n157 ) , .B2( u0_u5_u2_n170 ) );
  INV_X1 u0_u5_u2_U93 (.A( u0_u5_u2_n163 ) , .ZN( u0_u5_u2_n186 ) );
  OR4_X1 u0_u5_u2_U94 (.ZN( u0_out5_6 ) , .A4( u0_u5_u2_n161 ) , .A3( u0_u5_u2_n162 ) , .A2( u0_u5_u2_n163 ) , .A1( u0_u5_u2_n164 ) );
  OR3_X1 u0_u5_u2_U95 (.A2( u0_u5_u2_n159 ) , .A1( u0_u5_u2_n160 ) , .ZN( u0_u5_u2_n161 ) , .A3( u0_u5_u2_n183 ) );
  AOI21_X1 u0_u5_u2_U96 (.B2( u0_u5_u2_n154 ) , .B1( u0_u5_u2_n155 ) , .ZN( u0_u5_u2_n159 ) , .A( u0_u5_u2_n167 ) );
  NAND3_X1 u0_u5_u2_U97 (.A2( u0_u5_u2_n117 ) , .A1( u0_u5_u2_n122 ) , .A3( u0_u5_u2_n123 ) , .ZN( u0_u5_u2_n134 ) );
  NAND3_X1 u0_u5_u2_U98 (.ZN( u0_u5_u2_n110 ) , .A2( u0_u5_u2_n131 ) , .A3( u0_u5_u2_n139 ) , .A1( u0_u5_u2_n154 ) );
  NAND3_X1 u0_u5_u2_U99 (.A2( u0_u5_u2_n100 ) , .ZN( u0_u5_u2_n101 ) , .A1( u0_u5_u2_n104 ) , .A3( u0_u5_u2_n114 ) );
  OAI22_X1 u0_u5_u3_U10 (.B1( u0_u5_u3_n113 ) , .A2( u0_u5_u3_n135 ) , .A1( u0_u5_u3_n150 ) , .B2( u0_u5_u3_n164 ) , .ZN( u0_u5_u3_n98 ) );
  OAI211_X1 u0_u5_u3_U11 (.B( u0_u5_u3_n106 ) , .ZN( u0_u5_u3_n119 ) , .C2( u0_u5_u3_n128 ) , .C1( u0_u5_u3_n167 ) , .A( u0_u5_u3_n181 ) );
  AOI221_X1 u0_u5_u3_U12 (.C1( u0_u5_u3_n105 ) , .ZN( u0_u5_u3_n106 ) , .A( u0_u5_u3_n131 ) , .B2( u0_u5_u3_n132 ) , .C2( u0_u5_u3_n133 ) , .B1( u0_u5_u3_n169 ) );
  INV_X1 u0_u5_u3_U13 (.ZN( u0_u5_u3_n181 ) , .A( u0_u5_u3_n98 ) );
  NAND2_X1 u0_u5_u3_U14 (.ZN( u0_u5_u3_n105 ) , .A2( u0_u5_u3_n130 ) , .A1( u0_u5_u3_n155 ) );
  AOI22_X1 u0_u5_u3_U15 (.B1( u0_u5_u3_n115 ) , .A2( u0_u5_u3_n116 ) , .ZN( u0_u5_u3_n123 ) , .B2( u0_u5_u3_n133 ) , .A1( u0_u5_u3_n169 ) );
  NAND2_X1 u0_u5_u3_U16 (.ZN( u0_u5_u3_n116 ) , .A2( u0_u5_u3_n151 ) , .A1( u0_u5_u3_n182 ) );
  NOR2_X1 u0_u5_u3_U17 (.ZN( u0_u5_u3_n126 ) , .A2( u0_u5_u3_n150 ) , .A1( u0_u5_u3_n164 ) );
  AOI21_X1 u0_u5_u3_U18 (.ZN( u0_u5_u3_n112 ) , .B2( u0_u5_u3_n146 ) , .B1( u0_u5_u3_n155 ) , .A( u0_u5_u3_n167 ) );
  NAND2_X1 u0_u5_u3_U19 (.A1( u0_u5_u3_n135 ) , .ZN( u0_u5_u3_n142 ) , .A2( u0_u5_u3_n164 ) );
  NAND2_X1 u0_u5_u3_U20 (.ZN( u0_u5_u3_n132 ) , .A2( u0_u5_u3_n152 ) , .A1( u0_u5_u3_n156 ) );
  AND2_X1 u0_u5_u3_U21 (.A2( u0_u5_u3_n113 ) , .A1( u0_u5_u3_n114 ) , .ZN( u0_u5_u3_n151 ) );
  INV_X1 u0_u5_u3_U22 (.A( u0_u5_u3_n133 ) , .ZN( u0_u5_u3_n165 ) );
  INV_X1 u0_u5_u3_U23 (.A( u0_u5_u3_n135 ) , .ZN( u0_u5_u3_n170 ) );
  NAND2_X1 u0_u5_u3_U24 (.A1( u0_u5_u3_n107 ) , .A2( u0_u5_u3_n108 ) , .ZN( u0_u5_u3_n140 ) );
  NAND2_X1 u0_u5_u3_U25 (.ZN( u0_u5_u3_n117 ) , .A1( u0_u5_u3_n124 ) , .A2( u0_u5_u3_n148 ) );
  NAND2_X1 u0_u5_u3_U26 (.ZN( u0_u5_u3_n143 ) , .A1( u0_u5_u3_n165 ) , .A2( u0_u5_u3_n167 ) );
  INV_X1 u0_u5_u3_U27 (.A( u0_u5_u3_n130 ) , .ZN( u0_u5_u3_n177 ) );
  INV_X1 u0_u5_u3_U28 (.A( u0_u5_u3_n128 ) , .ZN( u0_u5_u3_n176 ) );
  INV_X1 u0_u5_u3_U29 (.A( u0_u5_u3_n155 ) , .ZN( u0_u5_u3_n174 ) );
  INV_X1 u0_u5_u3_U3 (.A( u0_u5_u3_n129 ) , .ZN( u0_u5_u3_n183 ) );
  INV_X1 u0_u5_u3_U30 (.A( u0_u5_u3_n139 ) , .ZN( u0_u5_u3_n185 ) );
  NOR2_X1 u0_u5_u3_U31 (.ZN( u0_u5_u3_n135 ) , .A2( u0_u5_u3_n141 ) , .A1( u0_u5_u3_n169 ) );
  OAI222_X1 u0_u5_u3_U32 (.C2( u0_u5_u3_n107 ) , .A2( u0_u5_u3_n108 ) , .B1( u0_u5_u3_n135 ) , .ZN( u0_u5_u3_n138 ) , .B2( u0_u5_u3_n146 ) , .C1( u0_u5_u3_n154 ) , .A1( u0_u5_u3_n164 ) );
  NOR4_X1 u0_u5_u3_U33 (.A4( u0_u5_u3_n157 ) , .A3( u0_u5_u3_n158 ) , .A2( u0_u5_u3_n159 ) , .A1( u0_u5_u3_n160 ) , .ZN( u0_u5_u3_n161 ) );
  AOI21_X1 u0_u5_u3_U34 (.B2( u0_u5_u3_n152 ) , .B1( u0_u5_u3_n153 ) , .ZN( u0_u5_u3_n158 ) , .A( u0_u5_u3_n164 ) );
  AOI21_X1 u0_u5_u3_U35 (.A( u0_u5_u3_n154 ) , .B2( u0_u5_u3_n155 ) , .B1( u0_u5_u3_n156 ) , .ZN( u0_u5_u3_n157 ) );
  AOI21_X1 u0_u5_u3_U36 (.A( u0_u5_u3_n149 ) , .B2( u0_u5_u3_n150 ) , .B1( u0_u5_u3_n151 ) , .ZN( u0_u5_u3_n159 ) );
  AOI211_X1 u0_u5_u3_U37 (.ZN( u0_u5_u3_n109 ) , .A( u0_u5_u3_n119 ) , .C2( u0_u5_u3_n129 ) , .B( u0_u5_u3_n138 ) , .C1( u0_u5_u3_n141 ) );
  AOI211_X1 u0_u5_u3_U38 (.B( u0_u5_u3_n119 ) , .A( u0_u5_u3_n120 ) , .C2( u0_u5_u3_n121 ) , .ZN( u0_u5_u3_n122 ) , .C1( u0_u5_u3_n179 ) );
  INV_X1 u0_u5_u3_U39 (.A( u0_u5_u3_n156 ) , .ZN( u0_u5_u3_n179 ) );
  INV_X1 u0_u5_u3_U4 (.A( u0_u5_u3_n140 ) , .ZN( u0_u5_u3_n182 ) );
  OAI22_X1 u0_u5_u3_U40 (.B1( u0_u5_u3_n118 ) , .ZN( u0_u5_u3_n120 ) , .A1( u0_u5_u3_n135 ) , .B2( u0_u5_u3_n154 ) , .A2( u0_u5_u3_n178 ) );
  AND3_X1 u0_u5_u3_U41 (.ZN( u0_u5_u3_n118 ) , .A2( u0_u5_u3_n124 ) , .A1( u0_u5_u3_n144 ) , .A3( u0_u5_u3_n152 ) );
  INV_X1 u0_u5_u3_U42 (.A( u0_u5_u3_n121 ) , .ZN( u0_u5_u3_n164 ) );
  NAND2_X1 u0_u5_u3_U43 (.ZN( u0_u5_u3_n133 ) , .A1( u0_u5_u3_n154 ) , .A2( u0_u5_u3_n164 ) );
  OAI211_X1 u0_u5_u3_U44 (.B( u0_u5_u3_n127 ) , .ZN( u0_u5_u3_n139 ) , .C1( u0_u5_u3_n150 ) , .C2( u0_u5_u3_n154 ) , .A( u0_u5_u3_n184 ) );
  INV_X1 u0_u5_u3_U45 (.A( u0_u5_u3_n125 ) , .ZN( u0_u5_u3_n184 ) );
  AOI221_X1 u0_u5_u3_U46 (.A( u0_u5_u3_n126 ) , .ZN( u0_u5_u3_n127 ) , .C2( u0_u5_u3_n132 ) , .C1( u0_u5_u3_n169 ) , .B2( u0_u5_u3_n170 ) , .B1( u0_u5_u3_n174 ) );
  OAI22_X1 u0_u5_u3_U47 (.A1( u0_u5_u3_n124 ) , .ZN( u0_u5_u3_n125 ) , .B2( u0_u5_u3_n145 ) , .A2( u0_u5_u3_n165 ) , .B1( u0_u5_u3_n167 ) );
  NOR2_X1 u0_u5_u3_U48 (.A1( u0_u5_u3_n113 ) , .ZN( u0_u5_u3_n131 ) , .A2( u0_u5_u3_n154 ) );
  NAND2_X1 u0_u5_u3_U49 (.A1( u0_u5_u3_n103 ) , .ZN( u0_u5_u3_n150 ) , .A2( u0_u5_u3_n99 ) );
  INV_X1 u0_u5_u3_U5 (.A( u0_u5_u3_n117 ) , .ZN( u0_u5_u3_n178 ) );
  NAND2_X1 u0_u5_u3_U50 (.A2( u0_u5_u3_n102 ) , .ZN( u0_u5_u3_n155 ) , .A1( u0_u5_u3_n97 ) );
  INV_X1 u0_u5_u3_U51 (.A( u0_u5_u3_n141 ) , .ZN( u0_u5_u3_n167 ) );
  AOI21_X1 u0_u5_u3_U52 (.B2( u0_u5_u3_n114 ) , .B1( u0_u5_u3_n146 ) , .A( u0_u5_u3_n154 ) , .ZN( u0_u5_u3_n94 ) );
  AOI21_X1 u0_u5_u3_U53 (.ZN( u0_u5_u3_n110 ) , .B2( u0_u5_u3_n142 ) , .B1( u0_u5_u3_n186 ) , .A( u0_u5_u3_n95 ) );
  INV_X1 u0_u5_u3_U54 (.A( u0_u5_u3_n145 ) , .ZN( u0_u5_u3_n186 ) );
  AOI21_X1 u0_u5_u3_U55 (.B1( u0_u5_u3_n124 ) , .A( u0_u5_u3_n149 ) , .B2( u0_u5_u3_n155 ) , .ZN( u0_u5_u3_n95 ) );
  INV_X1 u0_u5_u3_U56 (.A( u0_u5_u3_n149 ) , .ZN( u0_u5_u3_n169 ) );
  NAND2_X1 u0_u5_u3_U57 (.ZN( u0_u5_u3_n124 ) , .A1( u0_u5_u3_n96 ) , .A2( u0_u5_u3_n97 ) );
  NAND2_X1 u0_u5_u3_U58 (.A2( u0_u5_u3_n100 ) , .ZN( u0_u5_u3_n146 ) , .A1( u0_u5_u3_n96 ) );
  NAND2_X1 u0_u5_u3_U59 (.A1( u0_u5_u3_n101 ) , .ZN( u0_u5_u3_n145 ) , .A2( u0_u5_u3_n99 ) );
  AOI221_X1 u0_u5_u3_U6 (.A( u0_u5_u3_n131 ) , .C2( u0_u5_u3_n132 ) , .C1( u0_u5_u3_n133 ) , .ZN( u0_u5_u3_n134 ) , .B1( u0_u5_u3_n143 ) , .B2( u0_u5_u3_n177 ) );
  NAND2_X1 u0_u5_u3_U60 (.A1( u0_u5_u3_n100 ) , .ZN( u0_u5_u3_n156 ) , .A2( u0_u5_u3_n99 ) );
  NAND2_X1 u0_u5_u3_U61 (.A2( u0_u5_u3_n101 ) , .A1( u0_u5_u3_n104 ) , .ZN( u0_u5_u3_n148 ) );
  NAND2_X1 u0_u5_u3_U62 (.A1( u0_u5_u3_n100 ) , .A2( u0_u5_u3_n102 ) , .ZN( u0_u5_u3_n128 ) );
  NAND2_X1 u0_u5_u3_U63 (.A2( u0_u5_u3_n101 ) , .A1( u0_u5_u3_n102 ) , .ZN( u0_u5_u3_n152 ) );
  NAND2_X1 u0_u5_u3_U64 (.A2( u0_u5_u3_n101 ) , .ZN( u0_u5_u3_n114 ) , .A1( u0_u5_u3_n96 ) );
  NAND2_X1 u0_u5_u3_U65 (.ZN( u0_u5_u3_n107 ) , .A1( u0_u5_u3_n97 ) , .A2( u0_u5_u3_n99 ) );
  NAND2_X1 u0_u5_u3_U66 (.A2( u0_u5_u3_n100 ) , .A1( u0_u5_u3_n104 ) , .ZN( u0_u5_u3_n113 ) );
  NAND2_X1 u0_u5_u3_U67 (.A1( u0_u5_u3_n104 ) , .ZN( u0_u5_u3_n153 ) , .A2( u0_u5_u3_n97 ) );
  NAND2_X1 u0_u5_u3_U68 (.A2( u0_u5_u3_n103 ) , .A1( u0_u5_u3_n104 ) , .ZN( u0_u5_u3_n130 ) );
  NAND2_X1 u0_u5_u3_U69 (.A2( u0_u5_u3_n103 ) , .ZN( u0_u5_u3_n144 ) , .A1( u0_u5_u3_n96 ) );
  OAI22_X1 u0_u5_u3_U7 (.B2( u0_u5_u3_n147 ) , .A2( u0_u5_u3_n148 ) , .ZN( u0_u5_u3_n160 ) , .B1( u0_u5_u3_n165 ) , .A1( u0_u5_u3_n168 ) );
  NAND2_X1 u0_u5_u3_U70 (.A1( u0_u5_u3_n102 ) , .A2( u0_u5_u3_n103 ) , .ZN( u0_u5_u3_n108 ) );
  NOR2_X1 u0_u5_u3_U71 (.A2( u0_u5_X_19 ) , .A1( u0_u5_X_20 ) , .ZN( u0_u5_u3_n99 ) );
  NOR2_X1 u0_u5_u3_U72 (.A2( u0_u5_X_21 ) , .A1( u0_u5_X_24 ) , .ZN( u0_u5_u3_n103 ) );
  NOR2_X1 u0_u5_u3_U73 (.A2( u0_u5_X_24 ) , .A1( u0_u5_u3_n171 ) , .ZN( u0_u5_u3_n97 ) );
  NOR2_X1 u0_u5_u3_U74 (.A2( u0_u5_X_23 ) , .ZN( u0_u5_u3_n141 ) , .A1( u0_u5_u3_n166 ) );
  NOR2_X1 u0_u5_u3_U75 (.A2( u0_u5_X_19 ) , .A1( u0_u5_u3_n172 ) , .ZN( u0_u5_u3_n96 ) );
  NAND2_X1 u0_u5_u3_U76 (.A1( u0_u5_X_22 ) , .A2( u0_u5_X_23 ) , .ZN( u0_u5_u3_n154 ) );
  NAND2_X1 u0_u5_u3_U77 (.A1( u0_u5_X_23 ) , .ZN( u0_u5_u3_n149 ) , .A2( u0_u5_u3_n166 ) );
  NOR2_X1 u0_u5_u3_U78 (.A2( u0_u5_X_22 ) , .A1( u0_u5_X_23 ) , .ZN( u0_u5_u3_n121 ) );
  AND2_X1 u0_u5_u3_U79 (.A1( u0_u5_X_24 ) , .ZN( u0_u5_u3_n101 ) , .A2( u0_u5_u3_n171 ) );
  AND3_X1 u0_u5_u3_U8 (.A3( u0_u5_u3_n144 ) , .A2( u0_u5_u3_n145 ) , .A1( u0_u5_u3_n146 ) , .ZN( u0_u5_u3_n147 ) );
  AND2_X1 u0_u5_u3_U80 (.A1( u0_u5_X_19 ) , .ZN( u0_u5_u3_n102 ) , .A2( u0_u5_u3_n172 ) );
  AND2_X1 u0_u5_u3_U81 (.A1( u0_u5_X_21 ) , .A2( u0_u5_X_24 ) , .ZN( u0_u5_u3_n100 ) );
  AND2_X1 u0_u5_u3_U82 (.A2( u0_u5_X_19 ) , .A1( u0_u5_X_20 ) , .ZN( u0_u5_u3_n104 ) );
  INV_X1 u0_u5_u3_U83 (.A( u0_u5_X_22 ) , .ZN( u0_u5_u3_n166 ) );
  INV_X1 u0_u5_u3_U84 (.A( u0_u5_X_21 ) , .ZN( u0_u5_u3_n171 ) );
  INV_X1 u0_u5_u3_U85 (.A( u0_u5_X_20 ) , .ZN( u0_u5_u3_n172 ) );
  NAND4_X1 u0_u5_u3_U86 (.ZN( u0_out5_26 ) , .A4( u0_u5_u3_n109 ) , .A3( u0_u5_u3_n110 ) , .A2( u0_u5_u3_n111 ) , .A1( u0_u5_u3_n173 ) );
  INV_X1 u0_u5_u3_U87 (.ZN( u0_u5_u3_n173 ) , .A( u0_u5_u3_n94 ) );
  OAI21_X1 u0_u5_u3_U88 (.ZN( u0_u5_u3_n111 ) , .B2( u0_u5_u3_n117 ) , .A( u0_u5_u3_n133 ) , .B1( u0_u5_u3_n176 ) );
  NAND4_X1 u0_u5_u3_U89 (.ZN( u0_out5_20 ) , .A4( u0_u5_u3_n122 ) , .A3( u0_u5_u3_n123 ) , .A1( u0_u5_u3_n175 ) , .A2( u0_u5_u3_n180 ) );
  INV_X1 u0_u5_u3_U9 (.A( u0_u5_u3_n143 ) , .ZN( u0_u5_u3_n168 ) );
  INV_X1 u0_u5_u3_U90 (.A( u0_u5_u3_n126 ) , .ZN( u0_u5_u3_n180 ) );
  INV_X1 u0_u5_u3_U91 (.A( u0_u5_u3_n112 ) , .ZN( u0_u5_u3_n175 ) );
  NAND4_X1 u0_u5_u3_U92 (.ZN( u0_out5_1 ) , .A4( u0_u5_u3_n161 ) , .A3( u0_u5_u3_n162 ) , .A2( u0_u5_u3_n163 ) , .A1( u0_u5_u3_n185 ) );
  NAND2_X1 u0_u5_u3_U93 (.ZN( u0_u5_u3_n163 ) , .A2( u0_u5_u3_n170 ) , .A1( u0_u5_u3_n176 ) );
  AOI22_X1 u0_u5_u3_U94 (.B2( u0_u5_u3_n140 ) , .B1( u0_u5_u3_n141 ) , .A2( u0_u5_u3_n142 ) , .ZN( u0_u5_u3_n162 ) , .A1( u0_u5_u3_n177 ) );
  OR4_X1 u0_u5_u3_U95 (.ZN( u0_out5_10 ) , .A4( u0_u5_u3_n136 ) , .A3( u0_u5_u3_n137 ) , .A1( u0_u5_u3_n138 ) , .A2( u0_u5_u3_n139 ) );
  OAI222_X1 u0_u5_u3_U96 (.C1( u0_u5_u3_n128 ) , .ZN( u0_u5_u3_n137 ) , .B1( u0_u5_u3_n148 ) , .A2( u0_u5_u3_n150 ) , .B2( u0_u5_u3_n154 ) , .C2( u0_u5_u3_n164 ) , .A1( u0_u5_u3_n167 ) );
  OAI221_X1 u0_u5_u3_U97 (.A( u0_u5_u3_n134 ) , .B2( u0_u5_u3_n135 ) , .ZN( u0_u5_u3_n136 ) , .C1( u0_u5_u3_n149 ) , .B1( u0_u5_u3_n151 ) , .C2( u0_u5_u3_n183 ) );
  NAND3_X1 u0_u5_u3_U98 (.A1( u0_u5_u3_n114 ) , .ZN( u0_u5_u3_n115 ) , .A2( u0_u5_u3_n145 ) , .A3( u0_u5_u3_n153 ) );
  NAND3_X1 u0_u5_u3_U99 (.ZN( u0_u5_u3_n129 ) , .A2( u0_u5_u3_n144 ) , .A1( u0_u5_u3_n153 ) , .A3( u0_u5_u3_n182 ) );
  OAI22_X1 u0_u5_u4_U10 (.B2( u0_u5_u4_n135 ) , .ZN( u0_u5_u4_n137 ) , .B1( u0_u5_u4_n153 ) , .A1( u0_u5_u4_n155 ) , .A2( u0_u5_u4_n171 ) );
  AND3_X1 u0_u5_u4_U11 (.A2( u0_u5_u4_n134 ) , .ZN( u0_u5_u4_n135 ) , .A3( u0_u5_u4_n145 ) , .A1( u0_u5_u4_n157 ) );
  NAND2_X1 u0_u5_u4_U12 (.ZN( u0_u5_u4_n132 ) , .A2( u0_u5_u4_n170 ) , .A1( u0_u5_u4_n173 ) );
  AOI21_X1 u0_u5_u4_U13 (.B2( u0_u5_u4_n160 ) , .B1( u0_u5_u4_n161 ) , .ZN( u0_u5_u4_n162 ) , .A( u0_u5_u4_n170 ) );
  AOI21_X1 u0_u5_u4_U14 (.ZN( u0_u5_u4_n107 ) , .B2( u0_u5_u4_n143 ) , .A( u0_u5_u4_n174 ) , .B1( u0_u5_u4_n184 ) );
  AOI21_X1 u0_u5_u4_U15 (.B2( u0_u5_u4_n158 ) , .B1( u0_u5_u4_n159 ) , .ZN( u0_u5_u4_n163 ) , .A( u0_u5_u4_n174 ) );
  AOI21_X1 u0_u5_u4_U16 (.A( u0_u5_u4_n153 ) , .B2( u0_u5_u4_n154 ) , .B1( u0_u5_u4_n155 ) , .ZN( u0_u5_u4_n165 ) );
  AOI21_X1 u0_u5_u4_U17 (.A( u0_u5_u4_n156 ) , .B2( u0_u5_u4_n157 ) , .ZN( u0_u5_u4_n164 ) , .B1( u0_u5_u4_n184 ) );
  INV_X1 u0_u5_u4_U18 (.A( u0_u5_u4_n138 ) , .ZN( u0_u5_u4_n170 ) );
  AND2_X1 u0_u5_u4_U19 (.A2( u0_u5_u4_n120 ) , .ZN( u0_u5_u4_n155 ) , .A1( u0_u5_u4_n160 ) );
  INV_X1 u0_u5_u4_U20 (.A( u0_u5_u4_n156 ) , .ZN( u0_u5_u4_n175 ) );
  NAND2_X1 u0_u5_u4_U21 (.A2( u0_u5_u4_n118 ) , .ZN( u0_u5_u4_n131 ) , .A1( u0_u5_u4_n147 ) );
  NAND2_X1 u0_u5_u4_U22 (.A1( u0_u5_u4_n119 ) , .A2( u0_u5_u4_n120 ) , .ZN( u0_u5_u4_n130 ) );
  NAND2_X1 u0_u5_u4_U23 (.ZN( u0_u5_u4_n117 ) , .A2( u0_u5_u4_n118 ) , .A1( u0_u5_u4_n148 ) );
  NAND2_X1 u0_u5_u4_U24 (.ZN( u0_u5_u4_n129 ) , .A1( u0_u5_u4_n134 ) , .A2( u0_u5_u4_n148 ) );
  AND3_X1 u0_u5_u4_U25 (.A1( u0_u5_u4_n119 ) , .A2( u0_u5_u4_n143 ) , .A3( u0_u5_u4_n154 ) , .ZN( u0_u5_u4_n161 ) );
  AND2_X1 u0_u5_u4_U26 (.A1( u0_u5_u4_n145 ) , .A2( u0_u5_u4_n147 ) , .ZN( u0_u5_u4_n159 ) );
  OR3_X1 u0_u5_u4_U27 (.A3( u0_u5_u4_n114 ) , .A2( u0_u5_u4_n115 ) , .A1( u0_u5_u4_n116 ) , .ZN( u0_u5_u4_n136 ) );
  AOI21_X1 u0_u5_u4_U28 (.A( u0_u5_u4_n113 ) , .ZN( u0_u5_u4_n116 ) , .B2( u0_u5_u4_n173 ) , .B1( u0_u5_u4_n174 ) );
  AOI21_X1 u0_u5_u4_U29 (.ZN( u0_u5_u4_n115 ) , .B2( u0_u5_u4_n145 ) , .B1( u0_u5_u4_n146 ) , .A( u0_u5_u4_n156 ) );
  NOR2_X1 u0_u5_u4_U3 (.ZN( u0_u5_u4_n121 ) , .A1( u0_u5_u4_n181 ) , .A2( u0_u5_u4_n182 ) );
  OAI22_X1 u0_u5_u4_U30 (.ZN( u0_u5_u4_n114 ) , .A2( u0_u5_u4_n121 ) , .B1( u0_u5_u4_n160 ) , .B2( u0_u5_u4_n170 ) , .A1( u0_u5_u4_n171 ) );
  INV_X1 u0_u5_u4_U31 (.A( u0_u5_u4_n158 ) , .ZN( u0_u5_u4_n182 ) );
  INV_X1 u0_u5_u4_U32 (.ZN( u0_u5_u4_n181 ) , .A( u0_u5_u4_n96 ) );
  INV_X1 u0_u5_u4_U33 (.A( u0_u5_u4_n144 ) , .ZN( u0_u5_u4_n179 ) );
  INV_X1 u0_u5_u4_U34 (.A( u0_u5_u4_n157 ) , .ZN( u0_u5_u4_n178 ) );
  NAND2_X1 u0_u5_u4_U35 (.A2( u0_u5_u4_n154 ) , .A1( u0_u5_u4_n96 ) , .ZN( u0_u5_u4_n97 ) );
  INV_X1 u0_u5_u4_U36 (.ZN( u0_u5_u4_n186 ) , .A( u0_u5_u4_n95 ) );
  OAI221_X1 u0_u5_u4_U37 (.C1( u0_u5_u4_n134 ) , .B1( u0_u5_u4_n158 ) , .B2( u0_u5_u4_n171 ) , .C2( u0_u5_u4_n173 ) , .A( u0_u5_u4_n94 ) , .ZN( u0_u5_u4_n95 ) );
  AOI222_X1 u0_u5_u4_U38 (.B2( u0_u5_u4_n132 ) , .A1( u0_u5_u4_n138 ) , .C2( u0_u5_u4_n175 ) , .A2( u0_u5_u4_n179 ) , .C1( u0_u5_u4_n181 ) , .B1( u0_u5_u4_n185 ) , .ZN( u0_u5_u4_n94 ) );
  INV_X1 u0_u5_u4_U39 (.A( u0_u5_u4_n113 ) , .ZN( u0_u5_u4_n185 ) );
  INV_X1 u0_u5_u4_U4 (.A( u0_u5_u4_n117 ) , .ZN( u0_u5_u4_n184 ) );
  INV_X1 u0_u5_u4_U40 (.A( u0_u5_u4_n143 ) , .ZN( u0_u5_u4_n183 ) );
  NOR2_X1 u0_u5_u4_U41 (.ZN( u0_u5_u4_n138 ) , .A1( u0_u5_u4_n168 ) , .A2( u0_u5_u4_n169 ) );
  NOR2_X1 u0_u5_u4_U42 (.A1( u0_u5_u4_n150 ) , .A2( u0_u5_u4_n152 ) , .ZN( u0_u5_u4_n153 ) );
  NOR2_X1 u0_u5_u4_U43 (.A2( u0_u5_u4_n128 ) , .A1( u0_u5_u4_n138 ) , .ZN( u0_u5_u4_n156 ) );
  AOI22_X1 u0_u5_u4_U44 (.B2( u0_u5_u4_n122 ) , .A1( u0_u5_u4_n123 ) , .ZN( u0_u5_u4_n124 ) , .B1( u0_u5_u4_n128 ) , .A2( u0_u5_u4_n172 ) );
  INV_X1 u0_u5_u4_U45 (.A( u0_u5_u4_n153 ) , .ZN( u0_u5_u4_n172 ) );
  NAND2_X1 u0_u5_u4_U46 (.A2( u0_u5_u4_n120 ) , .ZN( u0_u5_u4_n123 ) , .A1( u0_u5_u4_n161 ) );
  AOI22_X1 u0_u5_u4_U47 (.B2( u0_u5_u4_n132 ) , .A2( u0_u5_u4_n133 ) , .ZN( u0_u5_u4_n140 ) , .A1( u0_u5_u4_n150 ) , .B1( u0_u5_u4_n179 ) );
  NAND2_X1 u0_u5_u4_U48 (.ZN( u0_u5_u4_n133 ) , .A2( u0_u5_u4_n146 ) , .A1( u0_u5_u4_n154 ) );
  NAND2_X1 u0_u5_u4_U49 (.A1( u0_u5_u4_n103 ) , .ZN( u0_u5_u4_n154 ) , .A2( u0_u5_u4_n98 ) );
  NOR4_X1 u0_u5_u4_U5 (.A4( u0_u5_u4_n106 ) , .A3( u0_u5_u4_n107 ) , .A2( u0_u5_u4_n108 ) , .A1( u0_u5_u4_n109 ) , .ZN( u0_u5_u4_n110 ) );
  NAND2_X1 u0_u5_u4_U50 (.A1( u0_u5_u4_n101 ) , .ZN( u0_u5_u4_n158 ) , .A2( u0_u5_u4_n99 ) );
  AOI21_X1 u0_u5_u4_U51 (.ZN( u0_u5_u4_n127 ) , .A( u0_u5_u4_n136 ) , .B2( u0_u5_u4_n150 ) , .B1( u0_u5_u4_n180 ) );
  INV_X1 u0_u5_u4_U52 (.A( u0_u5_u4_n160 ) , .ZN( u0_u5_u4_n180 ) );
  NAND2_X1 u0_u5_u4_U53 (.A2( u0_u5_u4_n104 ) , .A1( u0_u5_u4_n105 ) , .ZN( u0_u5_u4_n146 ) );
  NAND2_X1 u0_u5_u4_U54 (.A2( u0_u5_u4_n101 ) , .A1( u0_u5_u4_n102 ) , .ZN( u0_u5_u4_n160 ) );
  NAND2_X1 u0_u5_u4_U55 (.ZN( u0_u5_u4_n134 ) , .A1( u0_u5_u4_n98 ) , .A2( u0_u5_u4_n99 ) );
  NAND2_X1 u0_u5_u4_U56 (.A1( u0_u5_u4_n103 ) , .A2( u0_u5_u4_n104 ) , .ZN( u0_u5_u4_n143 ) );
  NAND2_X1 u0_u5_u4_U57 (.A2( u0_u5_u4_n105 ) , .ZN( u0_u5_u4_n145 ) , .A1( u0_u5_u4_n98 ) );
  NAND2_X1 u0_u5_u4_U58 (.A1( u0_u5_u4_n100 ) , .A2( u0_u5_u4_n105 ) , .ZN( u0_u5_u4_n120 ) );
  NAND2_X1 u0_u5_u4_U59 (.A1( u0_u5_u4_n102 ) , .A2( u0_u5_u4_n104 ) , .ZN( u0_u5_u4_n148 ) );
  AOI21_X1 u0_u5_u4_U6 (.ZN( u0_u5_u4_n106 ) , .B2( u0_u5_u4_n146 ) , .B1( u0_u5_u4_n158 ) , .A( u0_u5_u4_n170 ) );
  NAND2_X1 u0_u5_u4_U60 (.A2( u0_u5_u4_n100 ) , .A1( u0_u5_u4_n103 ) , .ZN( u0_u5_u4_n157 ) );
  INV_X1 u0_u5_u4_U61 (.A( u0_u5_u4_n150 ) , .ZN( u0_u5_u4_n173 ) );
  INV_X1 u0_u5_u4_U62 (.A( u0_u5_u4_n152 ) , .ZN( u0_u5_u4_n171 ) );
  NAND2_X1 u0_u5_u4_U63 (.A1( u0_u5_u4_n100 ) , .ZN( u0_u5_u4_n118 ) , .A2( u0_u5_u4_n99 ) );
  NAND2_X1 u0_u5_u4_U64 (.A2( u0_u5_u4_n100 ) , .A1( u0_u5_u4_n102 ) , .ZN( u0_u5_u4_n144 ) );
  NAND2_X1 u0_u5_u4_U65 (.A2( u0_u5_u4_n101 ) , .A1( u0_u5_u4_n105 ) , .ZN( u0_u5_u4_n96 ) );
  INV_X1 u0_u5_u4_U66 (.A( u0_u5_u4_n128 ) , .ZN( u0_u5_u4_n174 ) );
  NAND2_X1 u0_u5_u4_U67 (.A2( u0_u5_u4_n102 ) , .ZN( u0_u5_u4_n119 ) , .A1( u0_u5_u4_n98 ) );
  NAND2_X1 u0_u5_u4_U68 (.A2( u0_u5_u4_n101 ) , .A1( u0_u5_u4_n103 ) , .ZN( u0_u5_u4_n147 ) );
  NAND2_X1 u0_u5_u4_U69 (.A2( u0_u5_u4_n104 ) , .ZN( u0_u5_u4_n113 ) , .A1( u0_u5_u4_n99 ) );
  AOI21_X1 u0_u5_u4_U7 (.ZN( u0_u5_u4_n108 ) , .B2( u0_u5_u4_n134 ) , .B1( u0_u5_u4_n155 ) , .A( u0_u5_u4_n156 ) );
  NOR2_X1 u0_u5_u4_U70 (.A2( u0_u5_X_28 ) , .ZN( u0_u5_u4_n150 ) , .A1( u0_u5_u4_n168 ) );
  NOR2_X1 u0_u5_u4_U71 (.A2( u0_u5_X_29 ) , .ZN( u0_u5_u4_n152 ) , .A1( u0_u5_u4_n169 ) );
  NOR2_X1 u0_u5_u4_U72 (.A2( u0_u5_X_30 ) , .ZN( u0_u5_u4_n105 ) , .A1( u0_u5_u4_n176 ) );
  NOR2_X1 u0_u5_u4_U73 (.A2( u0_u5_X_26 ) , .ZN( u0_u5_u4_n100 ) , .A1( u0_u5_u4_n177 ) );
  NOR2_X1 u0_u5_u4_U74 (.A2( u0_u5_X_28 ) , .A1( u0_u5_X_29 ) , .ZN( u0_u5_u4_n128 ) );
  NOR2_X1 u0_u5_u4_U75 (.A2( u0_u5_X_27 ) , .A1( u0_u5_X_30 ) , .ZN( u0_u5_u4_n102 ) );
  NOR2_X1 u0_u5_u4_U76 (.A2( u0_u5_X_25 ) , .A1( u0_u5_X_26 ) , .ZN( u0_u5_u4_n98 ) );
  AND2_X1 u0_u5_u4_U77 (.A2( u0_u5_X_25 ) , .A1( u0_u5_X_26 ) , .ZN( u0_u5_u4_n104 ) );
  AND2_X1 u0_u5_u4_U78 (.A1( u0_u5_X_30 ) , .A2( u0_u5_u4_n176 ) , .ZN( u0_u5_u4_n99 ) );
  AND2_X1 u0_u5_u4_U79 (.A1( u0_u5_X_26 ) , .ZN( u0_u5_u4_n101 ) , .A2( u0_u5_u4_n177 ) );
  AOI21_X1 u0_u5_u4_U8 (.ZN( u0_u5_u4_n109 ) , .A( u0_u5_u4_n153 ) , .B1( u0_u5_u4_n159 ) , .B2( u0_u5_u4_n184 ) );
  AND2_X1 u0_u5_u4_U80 (.A1( u0_u5_X_27 ) , .A2( u0_u5_X_30 ) , .ZN( u0_u5_u4_n103 ) );
  INV_X1 u0_u5_u4_U81 (.A( u0_u5_X_28 ) , .ZN( u0_u5_u4_n169 ) );
  INV_X1 u0_u5_u4_U82 (.A( u0_u5_X_29 ) , .ZN( u0_u5_u4_n168 ) );
  INV_X1 u0_u5_u4_U83 (.A( u0_u5_X_25 ) , .ZN( u0_u5_u4_n177 ) );
  INV_X1 u0_u5_u4_U84 (.A( u0_u5_X_27 ) , .ZN( u0_u5_u4_n176 ) );
  NAND4_X1 u0_u5_u4_U85 (.ZN( u0_out5_25 ) , .A4( u0_u5_u4_n139 ) , .A3( u0_u5_u4_n140 ) , .A2( u0_u5_u4_n141 ) , .A1( u0_u5_u4_n142 ) );
  OAI21_X1 u0_u5_u4_U86 (.A( u0_u5_u4_n128 ) , .B2( u0_u5_u4_n129 ) , .B1( u0_u5_u4_n130 ) , .ZN( u0_u5_u4_n142 ) );
  OAI21_X1 u0_u5_u4_U87 (.B2( u0_u5_u4_n131 ) , .ZN( u0_u5_u4_n141 ) , .A( u0_u5_u4_n175 ) , .B1( u0_u5_u4_n183 ) );
  NAND4_X1 u0_u5_u4_U88 (.ZN( u0_out5_14 ) , .A4( u0_u5_u4_n124 ) , .A3( u0_u5_u4_n125 ) , .A2( u0_u5_u4_n126 ) , .A1( u0_u5_u4_n127 ) );
  AOI22_X1 u0_u5_u4_U89 (.B2( u0_u5_u4_n117 ) , .ZN( u0_u5_u4_n126 ) , .A1( u0_u5_u4_n129 ) , .B1( u0_u5_u4_n152 ) , .A2( u0_u5_u4_n175 ) );
  AOI211_X1 u0_u5_u4_U9 (.B( u0_u5_u4_n136 ) , .A( u0_u5_u4_n137 ) , .C2( u0_u5_u4_n138 ) , .ZN( u0_u5_u4_n139 ) , .C1( u0_u5_u4_n182 ) );
  AOI22_X1 u0_u5_u4_U90 (.ZN( u0_u5_u4_n125 ) , .B2( u0_u5_u4_n131 ) , .A2( u0_u5_u4_n132 ) , .B1( u0_u5_u4_n138 ) , .A1( u0_u5_u4_n178 ) );
  NAND4_X1 u0_u5_u4_U91 (.ZN( u0_out5_8 ) , .A4( u0_u5_u4_n110 ) , .A3( u0_u5_u4_n111 ) , .A2( u0_u5_u4_n112 ) , .A1( u0_u5_u4_n186 ) );
  NAND2_X1 u0_u5_u4_U92 (.ZN( u0_u5_u4_n112 ) , .A2( u0_u5_u4_n130 ) , .A1( u0_u5_u4_n150 ) );
  AOI22_X1 u0_u5_u4_U93 (.ZN( u0_u5_u4_n111 ) , .B2( u0_u5_u4_n132 ) , .A1( u0_u5_u4_n152 ) , .B1( u0_u5_u4_n178 ) , .A2( u0_u5_u4_n97 ) );
  AOI22_X1 u0_u5_u4_U94 (.B2( u0_u5_u4_n149 ) , .B1( u0_u5_u4_n150 ) , .A2( u0_u5_u4_n151 ) , .A1( u0_u5_u4_n152 ) , .ZN( u0_u5_u4_n167 ) );
  NOR4_X1 u0_u5_u4_U95 (.A4( u0_u5_u4_n162 ) , .A3( u0_u5_u4_n163 ) , .A2( u0_u5_u4_n164 ) , .A1( u0_u5_u4_n165 ) , .ZN( u0_u5_u4_n166 ) );
  NAND3_X1 u0_u5_u4_U96 (.ZN( u0_out5_3 ) , .A3( u0_u5_u4_n166 ) , .A1( u0_u5_u4_n167 ) , .A2( u0_u5_u4_n186 ) );
  NAND3_X1 u0_u5_u4_U97 (.A3( u0_u5_u4_n146 ) , .A2( u0_u5_u4_n147 ) , .A1( u0_u5_u4_n148 ) , .ZN( u0_u5_u4_n149 ) );
  NAND3_X1 u0_u5_u4_U98 (.A3( u0_u5_u4_n143 ) , .A2( u0_u5_u4_n144 ) , .A1( u0_u5_u4_n145 ) , .ZN( u0_u5_u4_n151 ) );
  NAND3_X1 u0_u5_u4_U99 (.A3( u0_u5_u4_n121 ) , .ZN( u0_u5_u4_n122 ) , .A2( u0_u5_u4_n144 ) , .A1( u0_u5_u4_n154 ) );
  XOR2_X1 u0_u7_U11 (.B( u0_K8_44 ) , .A( u0_R6_29 ) , .Z( u0_u7_X_44 ) );
  XOR2_X1 u0_u7_U12 (.B( u0_K8_43 ) , .A( u0_R6_28 ) , .Z( u0_u7_X_43 ) );
  XOR2_X1 u0_u7_U21 (.B( u0_K8_35 ) , .A( u0_R6_24 ) , .Z( u0_u7_X_35 ) );
  XOR2_X1 u0_u7_U22 (.B( u0_K8_34 ) , .A( u0_R6_23 ) , .Z( u0_u7_X_34 ) );
  XOR2_X1 u0_u7_U24 (.B( u0_K8_32 ) , .A( u0_R6_21 ) , .Z( u0_u7_X_32 ) );
  XOR2_X1 u0_u7_U25 (.B( u0_K8_31 ) , .A( u0_R6_20 ) , .Z( u0_u7_X_31 ) );
  XOR2_X1 u0_u7_U26 (.B( u0_K8_30 ) , .A( u0_R6_21 ) , .Z( u0_u7_X_30 ) );
  XOR2_X1 u0_u7_U28 (.B( u0_K8_29 ) , .A( u0_R6_20 ) , .Z( u0_u7_X_29 ) );
  XOR2_X1 u0_u7_U30 (.B( u0_K8_27 ) , .A( u0_R6_18 ) , .Z( u0_u7_X_27 ) );
  XOR2_X1 u0_u7_U31 (.B( u0_K8_26 ) , .A( u0_R6_17 ) , .Z( u0_u7_X_26 ) );
  XOR2_X1 u0_u7_U32 (.B( u0_K8_25 ) , .A( u0_R6_16 ) , .Z( u0_u7_X_25 ) );
  XOR2_X1 u0_u7_U33 (.B( u0_K8_24 ) , .A( u0_R6_17 ) , .Z( u0_u7_X_24 ) );
  XOR2_X1 u0_u7_U34 (.B( u0_K8_23 ) , .A( u0_R6_16 ) , .Z( u0_u7_X_23 ) );
  XOR2_X1 u0_u7_U36 (.B( u0_K8_21 ) , .A( u0_R6_14 ) , .Z( u0_u7_X_21 ) );
  XOR2_X1 u0_u7_U37 (.B( u0_K8_20 ) , .A( u0_R6_13 ) , .Z( u0_u7_X_20 ) );
  XOR2_X1 u0_u7_U39 (.B( u0_K8_19 ) , .A( u0_R6_12 ) , .Z( u0_u7_X_19 ) );
  XOR2_X1 u0_u7_U7 (.B( u0_K8_48 ) , .A( u0_R6_1 ) , .Z( u0_u7_X_48 ) );
  XOR2_X1 u0_u7_U8 (.B( u0_K8_47 ) , .A( u0_R6_32 ) , .Z( u0_u7_X_47 ) );
  OAI22_X1 u0_u7_u3_U10 (.B1( u0_u7_u3_n113 ) , .A2( u0_u7_u3_n135 ) , .A1( u0_u7_u3_n150 ) , .B2( u0_u7_u3_n164 ) , .ZN( u0_u7_u3_n98 ) );
  OAI211_X1 u0_u7_u3_U11 (.B( u0_u7_u3_n106 ) , .ZN( u0_u7_u3_n119 ) , .C2( u0_u7_u3_n128 ) , .C1( u0_u7_u3_n167 ) , .A( u0_u7_u3_n181 ) );
  AOI221_X1 u0_u7_u3_U12 (.C1( u0_u7_u3_n105 ) , .ZN( u0_u7_u3_n106 ) , .A( u0_u7_u3_n131 ) , .B2( u0_u7_u3_n132 ) , .C2( u0_u7_u3_n133 ) , .B1( u0_u7_u3_n169 ) );
  INV_X1 u0_u7_u3_U13 (.ZN( u0_u7_u3_n181 ) , .A( u0_u7_u3_n98 ) );
  NAND2_X1 u0_u7_u3_U14 (.ZN( u0_u7_u3_n105 ) , .A2( u0_u7_u3_n130 ) , .A1( u0_u7_u3_n155 ) );
  AOI22_X1 u0_u7_u3_U15 (.B1( u0_u7_u3_n115 ) , .A2( u0_u7_u3_n116 ) , .ZN( u0_u7_u3_n123 ) , .B2( u0_u7_u3_n133 ) , .A1( u0_u7_u3_n169 ) );
  NAND2_X1 u0_u7_u3_U16 (.ZN( u0_u7_u3_n116 ) , .A2( u0_u7_u3_n151 ) , .A1( u0_u7_u3_n182 ) );
  NOR2_X1 u0_u7_u3_U17 (.ZN( u0_u7_u3_n126 ) , .A2( u0_u7_u3_n150 ) , .A1( u0_u7_u3_n164 ) );
  AOI21_X1 u0_u7_u3_U18 (.ZN( u0_u7_u3_n112 ) , .B2( u0_u7_u3_n146 ) , .B1( u0_u7_u3_n155 ) , .A( u0_u7_u3_n167 ) );
  NAND2_X1 u0_u7_u3_U19 (.A1( u0_u7_u3_n135 ) , .ZN( u0_u7_u3_n142 ) , .A2( u0_u7_u3_n164 ) );
  NAND2_X1 u0_u7_u3_U20 (.ZN( u0_u7_u3_n132 ) , .A2( u0_u7_u3_n152 ) , .A1( u0_u7_u3_n156 ) );
  AND2_X1 u0_u7_u3_U21 (.A2( u0_u7_u3_n113 ) , .A1( u0_u7_u3_n114 ) , .ZN( u0_u7_u3_n151 ) );
  INV_X1 u0_u7_u3_U22 (.A( u0_u7_u3_n133 ) , .ZN( u0_u7_u3_n165 ) );
  INV_X1 u0_u7_u3_U23 (.A( u0_u7_u3_n135 ) , .ZN( u0_u7_u3_n170 ) );
  NAND2_X1 u0_u7_u3_U24 (.A1( u0_u7_u3_n107 ) , .A2( u0_u7_u3_n108 ) , .ZN( u0_u7_u3_n140 ) );
  NAND2_X1 u0_u7_u3_U25 (.ZN( u0_u7_u3_n117 ) , .A1( u0_u7_u3_n124 ) , .A2( u0_u7_u3_n148 ) );
  NAND2_X1 u0_u7_u3_U26 (.ZN( u0_u7_u3_n143 ) , .A1( u0_u7_u3_n165 ) , .A2( u0_u7_u3_n167 ) );
  INV_X1 u0_u7_u3_U27 (.A( u0_u7_u3_n130 ) , .ZN( u0_u7_u3_n177 ) );
  INV_X1 u0_u7_u3_U28 (.A( u0_u7_u3_n128 ) , .ZN( u0_u7_u3_n176 ) );
  INV_X1 u0_u7_u3_U29 (.A( u0_u7_u3_n155 ) , .ZN( u0_u7_u3_n174 ) );
  INV_X1 u0_u7_u3_U3 (.A( u0_u7_u3_n129 ) , .ZN( u0_u7_u3_n183 ) );
  INV_X1 u0_u7_u3_U30 (.A( u0_u7_u3_n139 ) , .ZN( u0_u7_u3_n185 ) );
  NOR2_X1 u0_u7_u3_U31 (.ZN( u0_u7_u3_n135 ) , .A2( u0_u7_u3_n141 ) , .A1( u0_u7_u3_n169 ) );
  OAI222_X1 u0_u7_u3_U32 (.C2( u0_u7_u3_n107 ) , .A2( u0_u7_u3_n108 ) , .B1( u0_u7_u3_n135 ) , .ZN( u0_u7_u3_n138 ) , .B2( u0_u7_u3_n146 ) , .C1( u0_u7_u3_n154 ) , .A1( u0_u7_u3_n164 ) );
  NOR4_X1 u0_u7_u3_U33 (.A4( u0_u7_u3_n157 ) , .A3( u0_u7_u3_n158 ) , .A2( u0_u7_u3_n159 ) , .A1( u0_u7_u3_n160 ) , .ZN( u0_u7_u3_n161 ) );
  AOI21_X1 u0_u7_u3_U34 (.B2( u0_u7_u3_n152 ) , .B1( u0_u7_u3_n153 ) , .ZN( u0_u7_u3_n158 ) , .A( u0_u7_u3_n164 ) );
  AOI21_X1 u0_u7_u3_U35 (.A( u0_u7_u3_n154 ) , .B2( u0_u7_u3_n155 ) , .B1( u0_u7_u3_n156 ) , .ZN( u0_u7_u3_n157 ) );
  AOI21_X1 u0_u7_u3_U36 (.A( u0_u7_u3_n149 ) , .B2( u0_u7_u3_n150 ) , .B1( u0_u7_u3_n151 ) , .ZN( u0_u7_u3_n159 ) );
  AOI211_X1 u0_u7_u3_U37 (.ZN( u0_u7_u3_n109 ) , .A( u0_u7_u3_n119 ) , .C2( u0_u7_u3_n129 ) , .B( u0_u7_u3_n138 ) , .C1( u0_u7_u3_n141 ) );
  AOI211_X1 u0_u7_u3_U38 (.B( u0_u7_u3_n119 ) , .A( u0_u7_u3_n120 ) , .C2( u0_u7_u3_n121 ) , .ZN( u0_u7_u3_n122 ) , .C1( u0_u7_u3_n179 ) );
  INV_X1 u0_u7_u3_U39 (.A( u0_u7_u3_n156 ) , .ZN( u0_u7_u3_n179 ) );
  INV_X1 u0_u7_u3_U4 (.A( u0_u7_u3_n140 ) , .ZN( u0_u7_u3_n182 ) );
  OAI22_X1 u0_u7_u3_U40 (.B1( u0_u7_u3_n118 ) , .ZN( u0_u7_u3_n120 ) , .A1( u0_u7_u3_n135 ) , .B2( u0_u7_u3_n154 ) , .A2( u0_u7_u3_n178 ) );
  AND3_X1 u0_u7_u3_U41 (.ZN( u0_u7_u3_n118 ) , .A2( u0_u7_u3_n124 ) , .A1( u0_u7_u3_n144 ) , .A3( u0_u7_u3_n152 ) );
  INV_X1 u0_u7_u3_U42 (.A( u0_u7_u3_n121 ) , .ZN( u0_u7_u3_n164 ) );
  NAND2_X1 u0_u7_u3_U43 (.ZN( u0_u7_u3_n133 ) , .A1( u0_u7_u3_n154 ) , .A2( u0_u7_u3_n164 ) );
  OAI211_X1 u0_u7_u3_U44 (.B( u0_u7_u3_n127 ) , .ZN( u0_u7_u3_n139 ) , .C1( u0_u7_u3_n150 ) , .C2( u0_u7_u3_n154 ) , .A( u0_u7_u3_n184 ) );
  INV_X1 u0_u7_u3_U45 (.A( u0_u7_u3_n125 ) , .ZN( u0_u7_u3_n184 ) );
  AOI221_X1 u0_u7_u3_U46 (.A( u0_u7_u3_n126 ) , .ZN( u0_u7_u3_n127 ) , .C2( u0_u7_u3_n132 ) , .C1( u0_u7_u3_n169 ) , .B2( u0_u7_u3_n170 ) , .B1( u0_u7_u3_n174 ) );
  OAI22_X1 u0_u7_u3_U47 (.A1( u0_u7_u3_n124 ) , .ZN( u0_u7_u3_n125 ) , .B2( u0_u7_u3_n145 ) , .A2( u0_u7_u3_n165 ) , .B1( u0_u7_u3_n167 ) );
  NOR2_X1 u0_u7_u3_U48 (.A1( u0_u7_u3_n113 ) , .ZN( u0_u7_u3_n131 ) , .A2( u0_u7_u3_n154 ) );
  NAND2_X1 u0_u7_u3_U49 (.A1( u0_u7_u3_n103 ) , .ZN( u0_u7_u3_n150 ) , .A2( u0_u7_u3_n99 ) );
  INV_X1 u0_u7_u3_U5 (.A( u0_u7_u3_n117 ) , .ZN( u0_u7_u3_n178 ) );
  NAND2_X1 u0_u7_u3_U50 (.A2( u0_u7_u3_n102 ) , .ZN( u0_u7_u3_n155 ) , .A1( u0_u7_u3_n97 ) );
  INV_X1 u0_u7_u3_U51 (.A( u0_u7_u3_n141 ) , .ZN( u0_u7_u3_n167 ) );
  AOI21_X1 u0_u7_u3_U52 (.B2( u0_u7_u3_n114 ) , .B1( u0_u7_u3_n146 ) , .A( u0_u7_u3_n154 ) , .ZN( u0_u7_u3_n94 ) );
  AOI21_X1 u0_u7_u3_U53 (.ZN( u0_u7_u3_n110 ) , .B2( u0_u7_u3_n142 ) , .B1( u0_u7_u3_n186 ) , .A( u0_u7_u3_n95 ) );
  INV_X1 u0_u7_u3_U54 (.A( u0_u7_u3_n145 ) , .ZN( u0_u7_u3_n186 ) );
  AOI21_X1 u0_u7_u3_U55 (.B1( u0_u7_u3_n124 ) , .A( u0_u7_u3_n149 ) , .B2( u0_u7_u3_n155 ) , .ZN( u0_u7_u3_n95 ) );
  INV_X1 u0_u7_u3_U56 (.A( u0_u7_u3_n149 ) , .ZN( u0_u7_u3_n169 ) );
  NAND2_X1 u0_u7_u3_U57 (.ZN( u0_u7_u3_n124 ) , .A1( u0_u7_u3_n96 ) , .A2( u0_u7_u3_n97 ) );
  NAND2_X1 u0_u7_u3_U58 (.A2( u0_u7_u3_n100 ) , .ZN( u0_u7_u3_n146 ) , .A1( u0_u7_u3_n96 ) );
  NAND2_X1 u0_u7_u3_U59 (.A1( u0_u7_u3_n101 ) , .ZN( u0_u7_u3_n145 ) , .A2( u0_u7_u3_n99 ) );
  AOI221_X1 u0_u7_u3_U6 (.A( u0_u7_u3_n131 ) , .C2( u0_u7_u3_n132 ) , .C1( u0_u7_u3_n133 ) , .ZN( u0_u7_u3_n134 ) , .B1( u0_u7_u3_n143 ) , .B2( u0_u7_u3_n177 ) );
  NAND2_X1 u0_u7_u3_U60 (.A1( u0_u7_u3_n100 ) , .ZN( u0_u7_u3_n156 ) , .A2( u0_u7_u3_n99 ) );
  NAND2_X1 u0_u7_u3_U61 (.A2( u0_u7_u3_n101 ) , .A1( u0_u7_u3_n104 ) , .ZN( u0_u7_u3_n148 ) );
  NAND2_X1 u0_u7_u3_U62 (.A1( u0_u7_u3_n100 ) , .A2( u0_u7_u3_n102 ) , .ZN( u0_u7_u3_n128 ) );
  NAND2_X1 u0_u7_u3_U63 (.A2( u0_u7_u3_n101 ) , .A1( u0_u7_u3_n102 ) , .ZN( u0_u7_u3_n152 ) );
  NAND2_X1 u0_u7_u3_U64 (.A2( u0_u7_u3_n101 ) , .ZN( u0_u7_u3_n114 ) , .A1( u0_u7_u3_n96 ) );
  NAND2_X1 u0_u7_u3_U65 (.ZN( u0_u7_u3_n107 ) , .A1( u0_u7_u3_n97 ) , .A2( u0_u7_u3_n99 ) );
  NAND2_X1 u0_u7_u3_U66 (.A2( u0_u7_u3_n100 ) , .A1( u0_u7_u3_n104 ) , .ZN( u0_u7_u3_n113 ) );
  NAND2_X1 u0_u7_u3_U67 (.A1( u0_u7_u3_n104 ) , .ZN( u0_u7_u3_n153 ) , .A2( u0_u7_u3_n97 ) );
  NAND2_X1 u0_u7_u3_U68 (.A2( u0_u7_u3_n103 ) , .A1( u0_u7_u3_n104 ) , .ZN( u0_u7_u3_n130 ) );
  NAND2_X1 u0_u7_u3_U69 (.A2( u0_u7_u3_n103 ) , .ZN( u0_u7_u3_n144 ) , .A1( u0_u7_u3_n96 ) );
  OAI22_X1 u0_u7_u3_U7 (.B2( u0_u7_u3_n147 ) , .A2( u0_u7_u3_n148 ) , .ZN( u0_u7_u3_n160 ) , .B1( u0_u7_u3_n165 ) , .A1( u0_u7_u3_n168 ) );
  NAND2_X1 u0_u7_u3_U70 (.A1( u0_u7_u3_n102 ) , .A2( u0_u7_u3_n103 ) , .ZN( u0_u7_u3_n108 ) );
  NOR2_X1 u0_u7_u3_U71 (.A2( u0_u7_X_19 ) , .A1( u0_u7_X_20 ) , .ZN( u0_u7_u3_n99 ) );
  NOR2_X1 u0_u7_u3_U72 (.A2( u0_u7_X_21 ) , .A1( u0_u7_X_24 ) , .ZN( u0_u7_u3_n103 ) );
  NOR2_X1 u0_u7_u3_U73 (.A2( u0_u7_X_24 ) , .A1( u0_u7_u3_n171 ) , .ZN( u0_u7_u3_n97 ) );
  NOR2_X1 u0_u7_u3_U74 (.A2( u0_u7_X_23 ) , .ZN( u0_u7_u3_n141 ) , .A1( u0_u7_u3_n166 ) );
  NOR2_X1 u0_u7_u3_U75 (.A2( u0_u7_X_19 ) , .A1( u0_u7_u3_n172 ) , .ZN( u0_u7_u3_n96 ) );
  NAND2_X1 u0_u7_u3_U76 (.A1( u0_u7_X_22 ) , .A2( u0_u7_X_23 ) , .ZN( u0_u7_u3_n154 ) );
  NAND2_X1 u0_u7_u3_U77 (.A1( u0_u7_X_23 ) , .ZN( u0_u7_u3_n149 ) , .A2( u0_u7_u3_n166 ) );
  NOR2_X1 u0_u7_u3_U78 (.A2( u0_u7_X_22 ) , .A1( u0_u7_X_23 ) , .ZN( u0_u7_u3_n121 ) );
  AND2_X1 u0_u7_u3_U79 (.A1( u0_u7_X_24 ) , .ZN( u0_u7_u3_n101 ) , .A2( u0_u7_u3_n171 ) );
  AND3_X1 u0_u7_u3_U8 (.A3( u0_u7_u3_n144 ) , .A2( u0_u7_u3_n145 ) , .A1( u0_u7_u3_n146 ) , .ZN( u0_u7_u3_n147 ) );
  AND2_X1 u0_u7_u3_U80 (.A1( u0_u7_X_19 ) , .ZN( u0_u7_u3_n102 ) , .A2( u0_u7_u3_n172 ) );
  AND2_X1 u0_u7_u3_U81 (.A1( u0_u7_X_21 ) , .A2( u0_u7_X_24 ) , .ZN( u0_u7_u3_n100 ) );
  AND2_X1 u0_u7_u3_U82 (.A2( u0_u7_X_19 ) , .A1( u0_u7_X_20 ) , .ZN( u0_u7_u3_n104 ) );
  INV_X1 u0_u7_u3_U83 (.A( u0_u7_X_22 ) , .ZN( u0_u7_u3_n166 ) );
  INV_X1 u0_u7_u3_U84 (.A( u0_u7_X_21 ) , .ZN( u0_u7_u3_n171 ) );
  INV_X1 u0_u7_u3_U85 (.A( u0_u7_X_20 ) , .ZN( u0_u7_u3_n172 ) );
  OR4_X1 u0_u7_u3_U86 (.ZN( u0_out7_10 ) , .A4( u0_u7_u3_n136 ) , .A3( u0_u7_u3_n137 ) , .A1( u0_u7_u3_n138 ) , .A2( u0_u7_u3_n139 ) );
  OAI222_X1 u0_u7_u3_U87 (.C1( u0_u7_u3_n128 ) , .ZN( u0_u7_u3_n137 ) , .B1( u0_u7_u3_n148 ) , .A2( u0_u7_u3_n150 ) , .B2( u0_u7_u3_n154 ) , .C2( u0_u7_u3_n164 ) , .A1( u0_u7_u3_n167 ) );
  OAI221_X1 u0_u7_u3_U88 (.A( u0_u7_u3_n134 ) , .B2( u0_u7_u3_n135 ) , .ZN( u0_u7_u3_n136 ) , .C1( u0_u7_u3_n149 ) , .B1( u0_u7_u3_n151 ) , .C2( u0_u7_u3_n183 ) );
  NAND4_X1 u0_u7_u3_U89 (.ZN( u0_out7_26 ) , .A4( u0_u7_u3_n109 ) , .A3( u0_u7_u3_n110 ) , .A2( u0_u7_u3_n111 ) , .A1( u0_u7_u3_n173 ) );
  INV_X1 u0_u7_u3_U9 (.A( u0_u7_u3_n143 ) , .ZN( u0_u7_u3_n168 ) );
  INV_X1 u0_u7_u3_U90 (.ZN( u0_u7_u3_n173 ) , .A( u0_u7_u3_n94 ) );
  OAI21_X1 u0_u7_u3_U91 (.ZN( u0_u7_u3_n111 ) , .B2( u0_u7_u3_n117 ) , .A( u0_u7_u3_n133 ) , .B1( u0_u7_u3_n176 ) );
  NAND4_X1 u0_u7_u3_U92 (.ZN( u0_out7_20 ) , .A4( u0_u7_u3_n122 ) , .A3( u0_u7_u3_n123 ) , .A1( u0_u7_u3_n175 ) , .A2( u0_u7_u3_n180 ) );
  INV_X1 u0_u7_u3_U93 (.A( u0_u7_u3_n126 ) , .ZN( u0_u7_u3_n180 ) );
  INV_X1 u0_u7_u3_U94 (.A( u0_u7_u3_n112 ) , .ZN( u0_u7_u3_n175 ) );
  NAND4_X1 u0_u7_u3_U95 (.ZN( u0_out7_1 ) , .A4( u0_u7_u3_n161 ) , .A3( u0_u7_u3_n162 ) , .A2( u0_u7_u3_n163 ) , .A1( u0_u7_u3_n185 ) );
  NAND2_X1 u0_u7_u3_U96 (.ZN( u0_u7_u3_n163 ) , .A2( u0_u7_u3_n170 ) , .A1( u0_u7_u3_n176 ) );
  AOI22_X1 u0_u7_u3_U97 (.B2( u0_u7_u3_n140 ) , .B1( u0_u7_u3_n141 ) , .A2( u0_u7_u3_n142 ) , .ZN( u0_u7_u3_n162 ) , .A1( u0_u7_u3_n177 ) );
  NAND3_X1 u0_u7_u3_U98 (.A1( u0_u7_u3_n114 ) , .ZN( u0_u7_u3_n115 ) , .A2( u0_u7_u3_n145 ) , .A3( u0_u7_u3_n153 ) );
  NAND3_X1 u0_u7_u3_U99 (.ZN( u0_u7_u3_n129 ) , .A2( u0_u7_u3_n144 ) , .A1( u0_u7_u3_n153 ) , .A3( u0_u7_u3_n182 ) );
  OAI22_X1 u0_u7_u4_U10 (.B2( u0_u7_u4_n135 ) , .ZN( u0_u7_u4_n137 ) , .B1( u0_u7_u4_n153 ) , .A1( u0_u7_u4_n155 ) , .A2( u0_u7_u4_n171 ) );
  AND3_X1 u0_u7_u4_U11 (.A2( u0_u7_u4_n134 ) , .ZN( u0_u7_u4_n135 ) , .A3( u0_u7_u4_n145 ) , .A1( u0_u7_u4_n157 ) );
  OR3_X1 u0_u7_u4_U12 (.A3( u0_u7_u4_n114 ) , .A2( u0_u7_u4_n115 ) , .A1( u0_u7_u4_n116 ) , .ZN( u0_u7_u4_n136 ) );
  AOI21_X1 u0_u7_u4_U13 (.A( u0_u7_u4_n113 ) , .ZN( u0_u7_u4_n116 ) , .B2( u0_u7_u4_n173 ) , .B1( u0_u7_u4_n174 ) );
  AOI21_X1 u0_u7_u4_U14 (.ZN( u0_u7_u4_n115 ) , .B2( u0_u7_u4_n145 ) , .B1( u0_u7_u4_n146 ) , .A( u0_u7_u4_n156 ) );
  OAI22_X1 u0_u7_u4_U15 (.ZN( u0_u7_u4_n114 ) , .A2( u0_u7_u4_n121 ) , .B1( u0_u7_u4_n160 ) , .B2( u0_u7_u4_n170 ) , .A1( u0_u7_u4_n171 ) );
  NAND2_X1 u0_u7_u4_U16 (.ZN( u0_u7_u4_n132 ) , .A2( u0_u7_u4_n170 ) , .A1( u0_u7_u4_n173 ) );
  AOI21_X1 u0_u7_u4_U17 (.B2( u0_u7_u4_n160 ) , .B1( u0_u7_u4_n161 ) , .ZN( u0_u7_u4_n162 ) , .A( u0_u7_u4_n170 ) );
  AOI21_X1 u0_u7_u4_U18 (.ZN( u0_u7_u4_n107 ) , .B2( u0_u7_u4_n143 ) , .A( u0_u7_u4_n174 ) , .B1( u0_u7_u4_n184 ) );
  AOI21_X1 u0_u7_u4_U19 (.B2( u0_u7_u4_n158 ) , .B1( u0_u7_u4_n159 ) , .ZN( u0_u7_u4_n163 ) , .A( u0_u7_u4_n174 ) );
  AOI21_X1 u0_u7_u4_U20 (.A( u0_u7_u4_n153 ) , .B2( u0_u7_u4_n154 ) , .B1( u0_u7_u4_n155 ) , .ZN( u0_u7_u4_n165 ) );
  AOI21_X1 u0_u7_u4_U21 (.A( u0_u7_u4_n156 ) , .B2( u0_u7_u4_n157 ) , .ZN( u0_u7_u4_n164 ) , .B1( u0_u7_u4_n184 ) );
  INV_X1 u0_u7_u4_U22 (.A( u0_u7_u4_n138 ) , .ZN( u0_u7_u4_n170 ) );
  AND2_X1 u0_u7_u4_U23 (.A2( u0_u7_u4_n120 ) , .ZN( u0_u7_u4_n155 ) , .A1( u0_u7_u4_n160 ) );
  INV_X1 u0_u7_u4_U24 (.A( u0_u7_u4_n156 ) , .ZN( u0_u7_u4_n175 ) );
  NAND2_X1 u0_u7_u4_U25 (.A2( u0_u7_u4_n118 ) , .ZN( u0_u7_u4_n131 ) , .A1( u0_u7_u4_n147 ) );
  NAND2_X1 u0_u7_u4_U26 (.A1( u0_u7_u4_n119 ) , .A2( u0_u7_u4_n120 ) , .ZN( u0_u7_u4_n130 ) );
  NAND2_X1 u0_u7_u4_U27 (.ZN( u0_u7_u4_n117 ) , .A2( u0_u7_u4_n118 ) , .A1( u0_u7_u4_n148 ) );
  NAND2_X1 u0_u7_u4_U28 (.ZN( u0_u7_u4_n129 ) , .A1( u0_u7_u4_n134 ) , .A2( u0_u7_u4_n148 ) );
  AND3_X1 u0_u7_u4_U29 (.A1( u0_u7_u4_n119 ) , .A2( u0_u7_u4_n143 ) , .A3( u0_u7_u4_n154 ) , .ZN( u0_u7_u4_n161 ) );
  NOR2_X1 u0_u7_u4_U3 (.ZN( u0_u7_u4_n121 ) , .A1( u0_u7_u4_n181 ) , .A2( u0_u7_u4_n182 ) );
  AND2_X1 u0_u7_u4_U30 (.A1( u0_u7_u4_n145 ) , .A2( u0_u7_u4_n147 ) , .ZN( u0_u7_u4_n159 ) );
  INV_X1 u0_u7_u4_U31 (.A( u0_u7_u4_n158 ) , .ZN( u0_u7_u4_n182 ) );
  INV_X1 u0_u7_u4_U32 (.ZN( u0_u7_u4_n181 ) , .A( u0_u7_u4_n96 ) );
  INV_X1 u0_u7_u4_U33 (.A( u0_u7_u4_n144 ) , .ZN( u0_u7_u4_n179 ) );
  INV_X1 u0_u7_u4_U34 (.A( u0_u7_u4_n157 ) , .ZN( u0_u7_u4_n178 ) );
  NAND2_X1 u0_u7_u4_U35 (.A2( u0_u7_u4_n154 ) , .A1( u0_u7_u4_n96 ) , .ZN( u0_u7_u4_n97 ) );
  INV_X1 u0_u7_u4_U36 (.ZN( u0_u7_u4_n186 ) , .A( u0_u7_u4_n95 ) );
  OAI221_X1 u0_u7_u4_U37 (.C1( u0_u7_u4_n134 ) , .B1( u0_u7_u4_n158 ) , .B2( u0_u7_u4_n171 ) , .C2( u0_u7_u4_n173 ) , .A( u0_u7_u4_n94 ) , .ZN( u0_u7_u4_n95 ) );
  AOI222_X1 u0_u7_u4_U38 (.B2( u0_u7_u4_n132 ) , .A1( u0_u7_u4_n138 ) , .C2( u0_u7_u4_n175 ) , .A2( u0_u7_u4_n179 ) , .C1( u0_u7_u4_n181 ) , .B1( u0_u7_u4_n185 ) , .ZN( u0_u7_u4_n94 ) );
  INV_X1 u0_u7_u4_U39 (.A( u0_u7_u4_n113 ) , .ZN( u0_u7_u4_n185 ) );
  INV_X1 u0_u7_u4_U4 (.A( u0_u7_u4_n117 ) , .ZN( u0_u7_u4_n184 ) );
  INV_X1 u0_u7_u4_U40 (.A( u0_u7_u4_n143 ) , .ZN( u0_u7_u4_n183 ) );
  NOR2_X1 u0_u7_u4_U41 (.ZN( u0_u7_u4_n138 ) , .A1( u0_u7_u4_n168 ) , .A2( u0_u7_u4_n169 ) );
  NOR2_X1 u0_u7_u4_U42 (.A1( u0_u7_u4_n150 ) , .A2( u0_u7_u4_n152 ) , .ZN( u0_u7_u4_n153 ) );
  NOR2_X1 u0_u7_u4_U43 (.A2( u0_u7_u4_n128 ) , .A1( u0_u7_u4_n138 ) , .ZN( u0_u7_u4_n156 ) );
  AOI22_X1 u0_u7_u4_U44 (.B2( u0_u7_u4_n122 ) , .A1( u0_u7_u4_n123 ) , .ZN( u0_u7_u4_n124 ) , .B1( u0_u7_u4_n128 ) , .A2( u0_u7_u4_n172 ) );
  NAND2_X1 u0_u7_u4_U45 (.A2( u0_u7_u4_n120 ) , .ZN( u0_u7_u4_n123 ) , .A1( u0_u7_u4_n161 ) );
  INV_X1 u0_u7_u4_U46 (.A( u0_u7_u4_n153 ) , .ZN( u0_u7_u4_n172 ) );
  AOI22_X1 u0_u7_u4_U47 (.B2( u0_u7_u4_n132 ) , .A2( u0_u7_u4_n133 ) , .ZN( u0_u7_u4_n140 ) , .A1( u0_u7_u4_n150 ) , .B1( u0_u7_u4_n179 ) );
  NAND2_X1 u0_u7_u4_U48 (.ZN( u0_u7_u4_n133 ) , .A2( u0_u7_u4_n146 ) , .A1( u0_u7_u4_n154 ) );
  NAND2_X1 u0_u7_u4_U49 (.A1( u0_u7_u4_n103 ) , .ZN( u0_u7_u4_n154 ) , .A2( u0_u7_u4_n98 ) );
  NOR4_X1 u0_u7_u4_U5 (.A4( u0_u7_u4_n106 ) , .A3( u0_u7_u4_n107 ) , .A2( u0_u7_u4_n108 ) , .A1( u0_u7_u4_n109 ) , .ZN( u0_u7_u4_n110 ) );
  NAND2_X1 u0_u7_u4_U50 (.A1( u0_u7_u4_n101 ) , .ZN( u0_u7_u4_n158 ) , .A2( u0_u7_u4_n99 ) );
  AOI21_X1 u0_u7_u4_U51 (.ZN( u0_u7_u4_n127 ) , .A( u0_u7_u4_n136 ) , .B2( u0_u7_u4_n150 ) , .B1( u0_u7_u4_n180 ) );
  INV_X1 u0_u7_u4_U52 (.A( u0_u7_u4_n160 ) , .ZN( u0_u7_u4_n180 ) );
  NAND2_X1 u0_u7_u4_U53 (.A2( u0_u7_u4_n104 ) , .A1( u0_u7_u4_n105 ) , .ZN( u0_u7_u4_n146 ) );
  NAND2_X1 u0_u7_u4_U54 (.A2( u0_u7_u4_n101 ) , .A1( u0_u7_u4_n102 ) , .ZN( u0_u7_u4_n160 ) );
  NAND2_X1 u0_u7_u4_U55 (.ZN( u0_u7_u4_n134 ) , .A1( u0_u7_u4_n98 ) , .A2( u0_u7_u4_n99 ) );
  NAND2_X1 u0_u7_u4_U56 (.A1( u0_u7_u4_n103 ) , .A2( u0_u7_u4_n104 ) , .ZN( u0_u7_u4_n143 ) );
  NAND2_X1 u0_u7_u4_U57 (.A2( u0_u7_u4_n105 ) , .ZN( u0_u7_u4_n145 ) , .A1( u0_u7_u4_n98 ) );
  NAND2_X1 u0_u7_u4_U58 (.A1( u0_u7_u4_n100 ) , .A2( u0_u7_u4_n105 ) , .ZN( u0_u7_u4_n120 ) );
  NAND2_X1 u0_u7_u4_U59 (.A1( u0_u7_u4_n102 ) , .A2( u0_u7_u4_n104 ) , .ZN( u0_u7_u4_n148 ) );
  AOI21_X1 u0_u7_u4_U6 (.ZN( u0_u7_u4_n106 ) , .B2( u0_u7_u4_n146 ) , .B1( u0_u7_u4_n158 ) , .A( u0_u7_u4_n170 ) );
  NAND2_X1 u0_u7_u4_U60 (.A2( u0_u7_u4_n100 ) , .A1( u0_u7_u4_n103 ) , .ZN( u0_u7_u4_n157 ) );
  INV_X1 u0_u7_u4_U61 (.A( u0_u7_u4_n150 ) , .ZN( u0_u7_u4_n173 ) );
  INV_X1 u0_u7_u4_U62 (.A( u0_u7_u4_n152 ) , .ZN( u0_u7_u4_n171 ) );
  NAND2_X1 u0_u7_u4_U63 (.A1( u0_u7_u4_n100 ) , .ZN( u0_u7_u4_n118 ) , .A2( u0_u7_u4_n99 ) );
  NAND2_X1 u0_u7_u4_U64 (.A2( u0_u7_u4_n100 ) , .A1( u0_u7_u4_n102 ) , .ZN( u0_u7_u4_n144 ) );
  NAND2_X1 u0_u7_u4_U65 (.A2( u0_u7_u4_n101 ) , .A1( u0_u7_u4_n105 ) , .ZN( u0_u7_u4_n96 ) );
  INV_X1 u0_u7_u4_U66 (.A( u0_u7_u4_n128 ) , .ZN( u0_u7_u4_n174 ) );
  NAND2_X1 u0_u7_u4_U67 (.A2( u0_u7_u4_n102 ) , .ZN( u0_u7_u4_n119 ) , .A1( u0_u7_u4_n98 ) );
  NAND2_X1 u0_u7_u4_U68 (.A2( u0_u7_u4_n101 ) , .A1( u0_u7_u4_n103 ) , .ZN( u0_u7_u4_n147 ) );
  NAND2_X1 u0_u7_u4_U69 (.A2( u0_u7_u4_n104 ) , .ZN( u0_u7_u4_n113 ) , .A1( u0_u7_u4_n99 ) );
  AOI21_X1 u0_u7_u4_U7 (.ZN( u0_u7_u4_n108 ) , .B2( u0_u7_u4_n134 ) , .B1( u0_u7_u4_n155 ) , .A( u0_u7_u4_n156 ) );
  NOR2_X1 u0_u7_u4_U70 (.A2( u0_u7_X_28 ) , .ZN( u0_u7_u4_n150 ) , .A1( u0_u7_u4_n168 ) );
  NOR2_X1 u0_u7_u4_U71 (.A2( u0_u7_X_29 ) , .ZN( u0_u7_u4_n152 ) , .A1( u0_u7_u4_n169 ) );
  NOR2_X1 u0_u7_u4_U72 (.A2( u0_u7_X_26 ) , .ZN( u0_u7_u4_n100 ) , .A1( u0_u7_u4_n177 ) );
  NOR2_X1 u0_u7_u4_U73 (.A2( u0_u7_X_30 ) , .ZN( u0_u7_u4_n105 ) , .A1( u0_u7_u4_n176 ) );
  NOR2_X1 u0_u7_u4_U74 (.A2( u0_u7_X_28 ) , .A1( u0_u7_X_29 ) , .ZN( u0_u7_u4_n128 ) );
  NOR2_X1 u0_u7_u4_U75 (.A2( u0_u7_X_25 ) , .A1( u0_u7_X_26 ) , .ZN( u0_u7_u4_n98 ) );
  NOR2_X1 u0_u7_u4_U76 (.A2( u0_u7_X_27 ) , .A1( u0_u7_X_30 ) , .ZN( u0_u7_u4_n102 ) );
  AND2_X1 u0_u7_u4_U77 (.A2( u0_u7_X_25 ) , .A1( u0_u7_X_26 ) , .ZN( u0_u7_u4_n104 ) );
  AND2_X1 u0_u7_u4_U78 (.A1( u0_u7_X_30 ) , .A2( u0_u7_u4_n176 ) , .ZN( u0_u7_u4_n99 ) );
  AND2_X1 u0_u7_u4_U79 (.A1( u0_u7_X_26 ) , .ZN( u0_u7_u4_n101 ) , .A2( u0_u7_u4_n177 ) );
  AOI21_X1 u0_u7_u4_U8 (.ZN( u0_u7_u4_n109 ) , .A( u0_u7_u4_n153 ) , .B1( u0_u7_u4_n159 ) , .B2( u0_u7_u4_n184 ) );
  AND2_X1 u0_u7_u4_U80 (.A1( u0_u7_X_27 ) , .A2( u0_u7_X_30 ) , .ZN( u0_u7_u4_n103 ) );
  INV_X1 u0_u7_u4_U81 (.A( u0_u7_X_28 ) , .ZN( u0_u7_u4_n169 ) );
  INV_X1 u0_u7_u4_U82 (.A( u0_u7_X_29 ) , .ZN( u0_u7_u4_n168 ) );
  INV_X1 u0_u7_u4_U83 (.A( u0_u7_X_25 ) , .ZN( u0_u7_u4_n177 ) );
  INV_X1 u0_u7_u4_U84 (.A( u0_u7_X_27 ) , .ZN( u0_u7_u4_n176 ) );
  NAND4_X1 u0_u7_u4_U85 (.ZN( u0_out7_25 ) , .A4( u0_u7_u4_n139 ) , .A3( u0_u7_u4_n140 ) , .A2( u0_u7_u4_n141 ) , .A1( u0_u7_u4_n142 ) );
  OAI21_X1 u0_u7_u4_U86 (.A( u0_u7_u4_n128 ) , .B2( u0_u7_u4_n129 ) , .B1( u0_u7_u4_n130 ) , .ZN( u0_u7_u4_n142 ) );
  OAI21_X1 u0_u7_u4_U87 (.B2( u0_u7_u4_n131 ) , .ZN( u0_u7_u4_n141 ) , .A( u0_u7_u4_n175 ) , .B1( u0_u7_u4_n183 ) );
  NAND4_X1 u0_u7_u4_U88 (.ZN( u0_out7_14 ) , .A4( u0_u7_u4_n124 ) , .A3( u0_u7_u4_n125 ) , .A2( u0_u7_u4_n126 ) , .A1( u0_u7_u4_n127 ) );
  AOI22_X1 u0_u7_u4_U89 (.B2( u0_u7_u4_n117 ) , .ZN( u0_u7_u4_n126 ) , .A1( u0_u7_u4_n129 ) , .B1( u0_u7_u4_n152 ) , .A2( u0_u7_u4_n175 ) );
  AOI211_X1 u0_u7_u4_U9 (.B( u0_u7_u4_n136 ) , .A( u0_u7_u4_n137 ) , .C2( u0_u7_u4_n138 ) , .ZN( u0_u7_u4_n139 ) , .C1( u0_u7_u4_n182 ) );
  AOI22_X1 u0_u7_u4_U90 (.ZN( u0_u7_u4_n125 ) , .B2( u0_u7_u4_n131 ) , .A2( u0_u7_u4_n132 ) , .B1( u0_u7_u4_n138 ) , .A1( u0_u7_u4_n178 ) );
  NAND4_X1 u0_u7_u4_U91 (.ZN( u0_out7_8 ) , .A4( u0_u7_u4_n110 ) , .A3( u0_u7_u4_n111 ) , .A2( u0_u7_u4_n112 ) , .A1( u0_u7_u4_n186 ) );
  NAND2_X1 u0_u7_u4_U92 (.ZN( u0_u7_u4_n112 ) , .A2( u0_u7_u4_n130 ) , .A1( u0_u7_u4_n150 ) );
  AOI22_X1 u0_u7_u4_U93 (.ZN( u0_u7_u4_n111 ) , .B2( u0_u7_u4_n132 ) , .A1( u0_u7_u4_n152 ) , .B1( u0_u7_u4_n178 ) , .A2( u0_u7_u4_n97 ) );
  AOI22_X1 u0_u7_u4_U94 (.B2( u0_u7_u4_n149 ) , .B1( u0_u7_u4_n150 ) , .A2( u0_u7_u4_n151 ) , .A1( u0_u7_u4_n152 ) , .ZN( u0_u7_u4_n167 ) );
  NOR4_X1 u0_u7_u4_U95 (.A4( u0_u7_u4_n162 ) , .A3( u0_u7_u4_n163 ) , .A2( u0_u7_u4_n164 ) , .A1( u0_u7_u4_n165 ) , .ZN( u0_u7_u4_n166 ) );
  NAND3_X1 u0_u7_u4_U96 (.ZN( u0_out7_3 ) , .A3( u0_u7_u4_n166 ) , .A1( u0_u7_u4_n167 ) , .A2( u0_u7_u4_n186 ) );
  NAND3_X1 u0_u7_u4_U97 (.A3( u0_u7_u4_n146 ) , .A2( u0_u7_u4_n147 ) , .A1( u0_u7_u4_n148 ) , .ZN( u0_u7_u4_n149 ) );
  NAND3_X1 u0_u7_u4_U98 (.A3( u0_u7_u4_n143 ) , .A2( u0_u7_u4_n144 ) , .A1( u0_u7_u4_n145 ) , .ZN( u0_u7_u4_n151 ) );
  NAND3_X1 u0_u7_u4_U99 (.A3( u0_u7_u4_n121 ) , .ZN( u0_u7_u4_n122 ) , .A2( u0_u7_u4_n144 ) , .A1( u0_u7_u4_n154 ) );
  INV_X1 u0_u7_u5_U10 (.A( u0_u7_u5_n121 ) , .ZN( u0_u7_u5_n177 ) );
  NOR3_X1 u0_u7_u5_U100 (.A3( u0_u7_u5_n141 ) , .A1( u0_u7_u5_n142 ) , .ZN( u0_u7_u5_n143 ) , .A2( u0_u7_u5_n191 ) );
  NAND4_X1 u0_u7_u5_U101 (.ZN( u0_out7_4 ) , .A4( u0_u7_u5_n112 ) , .A2( u0_u7_u5_n113 ) , .A1( u0_u7_u5_n114 ) , .A3( u0_u7_u5_n195 ) );
  AOI211_X1 u0_u7_u5_U102 (.A( u0_u7_u5_n110 ) , .C1( u0_u7_u5_n111 ) , .ZN( u0_u7_u5_n112 ) , .B( u0_u7_u5_n118 ) , .C2( u0_u7_u5_n177 ) );
  AOI222_X1 u0_u7_u5_U103 (.ZN( u0_u7_u5_n113 ) , .A1( u0_u7_u5_n131 ) , .C1( u0_u7_u5_n148 ) , .B2( u0_u7_u5_n174 ) , .C2( u0_u7_u5_n178 ) , .A2( u0_u7_u5_n179 ) , .B1( u0_u7_u5_n99 ) );
  NAND3_X1 u0_u7_u5_U104 (.A2( u0_u7_u5_n154 ) , .A3( u0_u7_u5_n158 ) , .A1( u0_u7_u5_n161 ) , .ZN( u0_u7_u5_n99 ) );
  NOR2_X1 u0_u7_u5_U11 (.ZN( u0_u7_u5_n160 ) , .A2( u0_u7_u5_n173 ) , .A1( u0_u7_u5_n177 ) );
  INV_X1 u0_u7_u5_U12 (.A( u0_u7_u5_n150 ) , .ZN( u0_u7_u5_n174 ) );
  AOI21_X1 u0_u7_u5_U13 (.A( u0_u7_u5_n160 ) , .B2( u0_u7_u5_n161 ) , .ZN( u0_u7_u5_n162 ) , .B1( u0_u7_u5_n192 ) );
  INV_X1 u0_u7_u5_U14 (.A( u0_u7_u5_n159 ) , .ZN( u0_u7_u5_n192 ) );
  AOI21_X1 u0_u7_u5_U15 (.A( u0_u7_u5_n156 ) , .B2( u0_u7_u5_n157 ) , .B1( u0_u7_u5_n158 ) , .ZN( u0_u7_u5_n163 ) );
  AOI21_X1 u0_u7_u5_U16 (.B2( u0_u7_u5_n139 ) , .B1( u0_u7_u5_n140 ) , .ZN( u0_u7_u5_n141 ) , .A( u0_u7_u5_n150 ) );
  OAI21_X1 u0_u7_u5_U17 (.A( u0_u7_u5_n133 ) , .B2( u0_u7_u5_n134 ) , .B1( u0_u7_u5_n135 ) , .ZN( u0_u7_u5_n142 ) );
  OAI21_X1 u0_u7_u5_U18 (.ZN( u0_u7_u5_n133 ) , .B2( u0_u7_u5_n147 ) , .A( u0_u7_u5_n173 ) , .B1( u0_u7_u5_n188 ) );
  NAND2_X1 u0_u7_u5_U19 (.A2( u0_u7_u5_n119 ) , .A1( u0_u7_u5_n123 ) , .ZN( u0_u7_u5_n137 ) );
  INV_X1 u0_u7_u5_U20 (.A( u0_u7_u5_n155 ) , .ZN( u0_u7_u5_n194 ) );
  NAND2_X1 u0_u7_u5_U21 (.A1( u0_u7_u5_n121 ) , .ZN( u0_u7_u5_n132 ) , .A2( u0_u7_u5_n172 ) );
  NAND2_X1 u0_u7_u5_U22 (.A2( u0_u7_u5_n122 ) , .ZN( u0_u7_u5_n136 ) , .A1( u0_u7_u5_n154 ) );
  NAND2_X1 u0_u7_u5_U23 (.A2( u0_u7_u5_n119 ) , .A1( u0_u7_u5_n120 ) , .ZN( u0_u7_u5_n159 ) );
  INV_X1 u0_u7_u5_U24 (.A( u0_u7_u5_n156 ) , .ZN( u0_u7_u5_n175 ) );
  INV_X1 u0_u7_u5_U25 (.A( u0_u7_u5_n158 ) , .ZN( u0_u7_u5_n188 ) );
  INV_X1 u0_u7_u5_U26 (.A( u0_u7_u5_n152 ) , .ZN( u0_u7_u5_n179 ) );
  INV_X1 u0_u7_u5_U27 (.A( u0_u7_u5_n140 ) , .ZN( u0_u7_u5_n182 ) );
  INV_X1 u0_u7_u5_U28 (.A( u0_u7_u5_n151 ) , .ZN( u0_u7_u5_n183 ) );
  INV_X1 u0_u7_u5_U29 (.A( u0_u7_u5_n123 ) , .ZN( u0_u7_u5_n185 ) );
  NOR2_X1 u0_u7_u5_U3 (.ZN( u0_u7_u5_n134 ) , .A1( u0_u7_u5_n183 ) , .A2( u0_u7_u5_n190 ) );
  INV_X1 u0_u7_u5_U30 (.A( u0_u7_u5_n161 ) , .ZN( u0_u7_u5_n184 ) );
  INV_X1 u0_u7_u5_U31 (.A( u0_u7_u5_n139 ) , .ZN( u0_u7_u5_n189 ) );
  INV_X1 u0_u7_u5_U32 (.A( u0_u7_u5_n157 ) , .ZN( u0_u7_u5_n190 ) );
  INV_X1 u0_u7_u5_U33 (.A( u0_u7_u5_n120 ) , .ZN( u0_u7_u5_n193 ) );
  NAND2_X1 u0_u7_u5_U34 (.ZN( u0_u7_u5_n111 ) , .A1( u0_u7_u5_n140 ) , .A2( u0_u7_u5_n155 ) );
  NOR2_X1 u0_u7_u5_U35 (.ZN( u0_u7_u5_n100 ) , .A1( u0_u7_u5_n170 ) , .A2( u0_u7_u5_n180 ) );
  INV_X1 u0_u7_u5_U36 (.A( u0_u7_u5_n117 ) , .ZN( u0_u7_u5_n196 ) );
  OAI221_X1 u0_u7_u5_U37 (.A( u0_u7_u5_n116 ) , .ZN( u0_u7_u5_n117 ) , .B2( u0_u7_u5_n119 ) , .C1( u0_u7_u5_n153 ) , .C2( u0_u7_u5_n158 ) , .B1( u0_u7_u5_n172 ) );
  AOI222_X1 u0_u7_u5_U38 (.ZN( u0_u7_u5_n116 ) , .B2( u0_u7_u5_n145 ) , .C1( u0_u7_u5_n148 ) , .A2( u0_u7_u5_n174 ) , .C2( u0_u7_u5_n177 ) , .B1( u0_u7_u5_n187 ) , .A1( u0_u7_u5_n193 ) );
  INV_X1 u0_u7_u5_U39 (.A( u0_u7_u5_n115 ) , .ZN( u0_u7_u5_n187 ) );
  INV_X1 u0_u7_u5_U4 (.A( u0_u7_u5_n138 ) , .ZN( u0_u7_u5_n191 ) );
  AOI22_X1 u0_u7_u5_U40 (.B2( u0_u7_u5_n131 ) , .A2( u0_u7_u5_n146 ) , .ZN( u0_u7_u5_n169 ) , .B1( u0_u7_u5_n174 ) , .A1( u0_u7_u5_n185 ) );
  NOR2_X1 u0_u7_u5_U41 (.A1( u0_u7_u5_n146 ) , .ZN( u0_u7_u5_n150 ) , .A2( u0_u7_u5_n173 ) );
  AOI21_X1 u0_u7_u5_U42 (.A( u0_u7_u5_n118 ) , .B2( u0_u7_u5_n145 ) , .ZN( u0_u7_u5_n168 ) , .B1( u0_u7_u5_n186 ) );
  INV_X1 u0_u7_u5_U43 (.A( u0_u7_u5_n122 ) , .ZN( u0_u7_u5_n186 ) );
  NOR2_X1 u0_u7_u5_U44 (.A1( u0_u7_u5_n146 ) , .ZN( u0_u7_u5_n152 ) , .A2( u0_u7_u5_n176 ) );
  NOR2_X1 u0_u7_u5_U45 (.A1( u0_u7_u5_n115 ) , .ZN( u0_u7_u5_n118 ) , .A2( u0_u7_u5_n153 ) );
  NOR2_X1 u0_u7_u5_U46 (.A2( u0_u7_u5_n145 ) , .ZN( u0_u7_u5_n156 ) , .A1( u0_u7_u5_n174 ) );
  NOR2_X1 u0_u7_u5_U47 (.ZN( u0_u7_u5_n121 ) , .A2( u0_u7_u5_n145 ) , .A1( u0_u7_u5_n176 ) );
  AOI22_X1 u0_u7_u5_U48 (.ZN( u0_u7_u5_n114 ) , .A2( u0_u7_u5_n137 ) , .A1( u0_u7_u5_n145 ) , .B2( u0_u7_u5_n175 ) , .B1( u0_u7_u5_n193 ) );
  OAI211_X1 u0_u7_u5_U49 (.B( u0_u7_u5_n124 ) , .A( u0_u7_u5_n125 ) , .C2( u0_u7_u5_n126 ) , .C1( u0_u7_u5_n127 ) , .ZN( u0_u7_u5_n128 ) );
  OAI21_X1 u0_u7_u5_U5 (.B2( u0_u7_u5_n136 ) , .B1( u0_u7_u5_n137 ) , .ZN( u0_u7_u5_n138 ) , .A( u0_u7_u5_n177 ) );
  NOR3_X1 u0_u7_u5_U50 (.ZN( u0_u7_u5_n127 ) , .A1( u0_u7_u5_n136 ) , .A3( u0_u7_u5_n148 ) , .A2( u0_u7_u5_n182 ) );
  OAI21_X1 u0_u7_u5_U51 (.ZN( u0_u7_u5_n124 ) , .A( u0_u7_u5_n177 ) , .B2( u0_u7_u5_n183 ) , .B1( u0_u7_u5_n189 ) );
  OAI21_X1 u0_u7_u5_U52 (.ZN( u0_u7_u5_n125 ) , .A( u0_u7_u5_n174 ) , .B2( u0_u7_u5_n185 ) , .B1( u0_u7_u5_n190 ) );
  AOI21_X1 u0_u7_u5_U53 (.A( u0_u7_u5_n153 ) , .B2( u0_u7_u5_n154 ) , .B1( u0_u7_u5_n155 ) , .ZN( u0_u7_u5_n164 ) );
  AOI21_X1 u0_u7_u5_U54 (.ZN( u0_u7_u5_n110 ) , .B1( u0_u7_u5_n122 ) , .B2( u0_u7_u5_n139 ) , .A( u0_u7_u5_n153 ) );
  INV_X1 u0_u7_u5_U55 (.A( u0_u7_u5_n153 ) , .ZN( u0_u7_u5_n176 ) );
  INV_X1 u0_u7_u5_U56 (.A( u0_u7_u5_n126 ) , .ZN( u0_u7_u5_n173 ) );
  AND2_X1 u0_u7_u5_U57 (.A2( u0_u7_u5_n104 ) , .A1( u0_u7_u5_n107 ) , .ZN( u0_u7_u5_n147 ) );
  AND2_X1 u0_u7_u5_U58 (.A2( u0_u7_u5_n104 ) , .A1( u0_u7_u5_n108 ) , .ZN( u0_u7_u5_n148 ) );
  NAND2_X1 u0_u7_u5_U59 (.A1( u0_u7_u5_n105 ) , .A2( u0_u7_u5_n106 ) , .ZN( u0_u7_u5_n158 ) );
  INV_X1 u0_u7_u5_U6 (.A( u0_u7_u5_n135 ) , .ZN( u0_u7_u5_n178 ) );
  NAND2_X1 u0_u7_u5_U60 (.A2( u0_u7_u5_n108 ) , .A1( u0_u7_u5_n109 ) , .ZN( u0_u7_u5_n139 ) );
  NAND2_X1 u0_u7_u5_U61 (.A1( u0_u7_u5_n106 ) , .A2( u0_u7_u5_n108 ) , .ZN( u0_u7_u5_n119 ) );
  NAND2_X1 u0_u7_u5_U62 (.A2( u0_u7_u5_n103 ) , .A1( u0_u7_u5_n105 ) , .ZN( u0_u7_u5_n140 ) );
  NAND2_X1 u0_u7_u5_U63 (.A2( u0_u7_u5_n104 ) , .A1( u0_u7_u5_n105 ) , .ZN( u0_u7_u5_n155 ) );
  NAND2_X1 u0_u7_u5_U64 (.A2( u0_u7_u5_n106 ) , .A1( u0_u7_u5_n107 ) , .ZN( u0_u7_u5_n122 ) );
  NAND2_X1 u0_u7_u5_U65 (.A2( u0_u7_u5_n100 ) , .A1( u0_u7_u5_n106 ) , .ZN( u0_u7_u5_n115 ) );
  NAND2_X1 u0_u7_u5_U66 (.A2( u0_u7_u5_n100 ) , .A1( u0_u7_u5_n103 ) , .ZN( u0_u7_u5_n161 ) );
  NAND2_X1 u0_u7_u5_U67 (.A1( u0_u7_u5_n105 ) , .A2( u0_u7_u5_n109 ) , .ZN( u0_u7_u5_n154 ) );
  INV_X1 u0_u7_u5_U68 (.A( u0_u7_u5_n146 ) , .ZN( u0_u7_u5_n172 ) );
  NAND2_X1 u0_u7_u5_U69 (.A1( u0_u7_u5_n103 ) , .A2( u0_u7_u5_n108 ) , .ZN( u0_u7_u5_n123 ) );
  OAI22_X1 u0_u7_u5_U7 (.B2( u0_u7_u5_n149 ) , .B1( u0_u7_u5_n150 ) , .A2( u0_u7_u5_n151 ) , .A1( u0_u7_u5_n152 ) , .ZN( u0_u7_u5_n165 ) );
  NAND2_X1 u0_u7_u5_U70 (.A2( u0_u7_u5_n103 ) , .A1( u0_u7_u5_n107 ) , .ZN( u0_u7_u5_n151 ) );
  NAND2_X1 u0_u7_u5_U71 (.A2( u0_u7_u5_n107 ) , .A1( u0_u7_u5_n109 ) , .ZN( u0_u7_u5_n120 ) );
  NAND2_X1 u0_u7_u5_U72 (.A2( u0_u7_u5_n100 ) , .A1( u0_u7_u5_n109 ) , .ZN( u0_u7_u5_n157 ) );
  AND2_X1 u0_u7_u5_U73 (.A2( u0_u7_u5_n100 ) , .A1( u0_u7_u5_n104 ) , .ZN( u0_u7_u5_n131 ) );
  INV_X1 u0_u7_u5_U74 (.A( u0_u7_u5_n102 ) , .ZN( u0_u7_u5_n195 ) );
  OAI221_X1 u0_u7_u5_U75 (.A( u0_u7_u5_n101 ) , .ZN( u0_u7_u5_n102 ) , .C2( u0_u7_u5_n115 ) , .C1( u0_u7_u5_n126 ) , .B1( u0_u7_u5_n134 ) , .B2( u0_u7_u5_n160 ) );
  OAI21_X1 u0_u7_u5_U76 (.ZN( u0_u7_u5_n101 ) , .B1( u0_u7_u5_n137 ) , .A( u0_u7_u5_n146 ) , .B2( u0_u7_u5_n147 ) );
  NOR2_X1 u0_u7_u5_U77 (.A2( u0_u7_X_34 ) , .A1( u0_u7_X_35 ) , .ZN( u0_u7_u5_n145 ) );
  NOR2_X1 u0_u7_u5_U78 (.A2( u0_u7_X_34 ) , .ZN( u0_u7_u5_n146 ) , .A1( u0_u7_u5_n171 ) );
  NOR2_X1 u0_u7_u5_U79 (.A2( u0_u7_X_31 ) , .A1( u0_u7_X_32 ) , .ZN( u0_u7_u5_n103 ) );
  NOR3_X1 u0_u7_u5_U8 (.A2( u0_u7_u5_n147 ) , .A1( u0_u7_u5_n148 ) , .ZN( u0_u7_u5_n149 ) , .A3( u0_u7_u5_n194 ) );
  NOR2_X1 u0_u7_u5_U80 (.A2( u0_u7_X_36 ) , .ZN( u0_u7_u5_n105 ) , .A1( u0_u7_u5_n180 ) );
  NOR2_X1 u0_u7_u5_U81 (.A2( u0_u7_X_33 ) , .ZN( u0_u7_u5_n108 ) , .A1( u0_u7_u5_n170 ) );
  NOR2_X1 u0_u7_u5_U82 (.A2( u0_u7_X_33 ) , .A1( u0_u7_X_36 ) , .ZN( u0_u7_u5_n107 ) );
  NOR2_X1 u0_u7_u5_U83 (.A2( u0_u7_X_31 ) , .ZN( u0_u7_u5_n104 ) , .A1( u0_u7_u5_n181 ) );
  NAND2_X1 u0_u7_u5_U84 (.A2( u0_u7_X_34 ) , .A1( u0_u7_X_35 ) , .ZN( u0_u7_u5_n153 ) );
  NAND2_X1 u0_u7_u5_U85 (.A1( u0_u7_X_34 ) , .ZN( u0_u7_u5_n126 ) , .A2( u0_u7_u5_n171 ) );
  AND2_X1 u0_u7_u5_U86 (.A1( u0_u7_X_31 ) , .A2( u0_u7_X_32 ) , .ZN( u0_u7_u5_n106 ) );
  AND2_X1 u0_u7_u5_U87 (.A1( u0_u7_X_31 ) , .ZN( u0_u7_u5_n109 ) , .A2( u0_u7_u5_n181 ) );
  INV_X1 u0_u7_u5_U88 (.A( u0_u7_X_33 ) , .ZN( u0_u7_u5_n180 ) );
  INV_X1 u0_u7_u5_U89 (.A( u0_u7_X_35 ) , .ZN( u0_u7_u5_n171 ) );
  NOR2_X1 u0_u7_u5_U9 (.ZN( u0_u7_u5_n135 ) , .A1( u0_u7_u5_n173 ) , .A2( u0_u7_u5_n176 ) );
  INV_X1 u0_u7_u5_U90 (.A( u0_u7_X_36 ) , .ZN( u0_u7_u5_n170 ) );
  INV_X1 u0_u7_u5_U91 (.A( u0_u7_X_32 ) , .ZN( u0_u7_u5_n181 ) );
  NAND4_X1 u0_u7_u5_U92 (.ZN( u0_out7_29 ) , .A4( u0_u7_u5_n129 ) , .A3( u0_u7_u5_n130 ) , .A2( u0_u7_u5_n168 ) , .A1( u0_u7_u5_n196 ) );
  AOI221_X1 u0_u7_u5_U93 (.A( u0_u7_u5_n128 ) , .ZN( u0_u7_u5_n129 ) , .C2( u0_u7_u5_n132 ) , .B2( u0_u7_u5_n159 ) , .B1( u0_u7_u5_n176 ) , .C1( u0_u7_u5_n184 ) );
  AOI222_X1 u0_u7_u5_U94 (.ZN( u0_u7_u5_n130 ) , .A2( u0_u7_u5_n146 ) , .B1( u0_u7_u5_n147 ) , .C2( u0_u7_u5_n175 ) , .B2( u0_u7_u5_n179 ) , .A1( u0_u7_u5_n188 ) , .C1( u0_u7_u5_n194 ) );
  NAND4_X1 u0_u7_u5_U95 (.ZN( u0_out7_19 ) , .A4( u0_u7_u5_n166 ) , .A3( u0_u7_u5_n167 ) , .A2( u0_u7_u5_n168 ) , .A1( u0_u7_u5_n169 ) );
  AOI22_X1 u0_u7_u5_U96 (.B2( u0_u7_u5_n145 ) , .A2( u0_u7_u5_n146 ) , .ZN( u0_u7_u5_n167 ) , .B1( u0_u7_u5_n182 ) , .A1( u0_u7_u5_n189 ) );
  NOR4_X1 u0_u7_u5_U97 (.A4( u0_u7_u5_n162 ) , .A3( u0_u7_u5_n163 ) , .A2( u0_u7_u5_n164 ) , .A1( u0_u7_u5_n165 ) , .ZN( u0_u7_u5_n166 ) );
  NAND4_X1 u0_u7_u5_U98 (.ZN( u0_out7_11 ) , .A4( u0_u7_u5_n143 ) , .A3( u0_u7_u5_n144 ) , .A2( u0_u7_u5_n169 ) , .A1( u0_u7_u5_n196 ) );
  AOI22_X1 u0_u7_u5_U99 (.A2( u0_u7_u5_n132 ) , .ZN( u0_u7_u5_n144 ) , .B2( u0_u7_u5_n145 ) , .B1( u0_u7_u5_n184 ) , .A1( u0_u7_u5_n194 ) );
  OAI221_X1 u0_u7_u7_U10 (.C1( u0_u7_u7_n101 ) , .C2( u0_u7_u7_n147 ) , .ZN( u0_u7_u7_n155 ) , .B2( u0_u7_u7_n162 ) , .A( u0_u7_u7_n91 ) , .B1( u0_u7_u7_n92 ) );
  AND3_X1 u0_u7_u7_U11 (.A3( u0_u7_u7_n110 ) , .A2( u0_u7_u7_n127 ) , .A1( u0_u7_u7_n132 ) , .ZN( u0_u7_u7_n92 ) );
  OAI21_X1 u0_u7_u7_U12 (.A( u0_u7_u7_n161 ) , .B1( u0_u7_u7_n168 ) , .B2( u0_u7_u7_n173 ) , .ZN( u0_u7_u7_n91 ) );
  AOI211_X1 u0_u7_u7_U13 (.A( u0_u7_u7_n117 ) , .ZN( u0_u7_u7_n118 ) , .C2( u0_u7_u7_n126 ) , .C1( u0_u7_u7_n177 ) , .B( u0_u7_u7_n180 ) );
  OAI22_X1 u0_u7_u7_U14 (.B1( u0_u7_u7_n115 ) , .ZN( u0_u7_u7_n117 ) , .A2( u0_u7_u7_n133 ) , .A1( u0_u7_u7_n137 ) , .B2( u0_u7_u7_n162 ) );
  INV_X1 u0_u7_u7_U15 (.A( u0_u7_u7_n116 ) , .ZN( u0_u7_u7_n180 ) );
  NOR3_X1 u0_u7_u7_U16 (.ZN( u0_u7_u7_n115 ) , .A3( u0_u7_u7_n145 ) , .A2( u0_u7_u7_n168 ) , .A1( u0_u7_u7_n169 ) );
  NOR3_X1 u0_u7_u7_U17 (.A2( u0_u7_u7_n134 ) , .A1( u0_u7_u7_n135 ) , .ZN( u0_u7_u7_n136 ) , .A3( u0_u7_u7_n171 ) );
  NOR2_X1 u0_u7_u7_U18 (.A1( u0_u7_u7_n130 ) , .A2( u0_u7_u7_n134 ) , .ZN( u0_u7_u7_n153 ) );
  NOR2_X1 u0_u7_u7_U19 (.ZN( u0_u7_u7_n111 ) , .A2( u0_u7_u7_n134 ) , .A1( u0_u7_u7_n169 ) );
  AOI21_X1 u0_u7_u7_U20 (.ZN( u0_u7_u7_n104 ) , .B2( u0_u7_u7_n112 ) , .B1( u0_u7_u7_n127 ) , .A( u0_u7_u7_n164 ) );
  AOI21_X1 u0_u7_u7_U21 (.ZN( u0_u7_u7_n106 ) , .B1( u0_u7_u7_n133 ) , .B2( u0_u7_u7_n146 ) , .A( u0_u7_u7_n162 ) );
  AOI21_X1 u0_u7_u7_U22 (.A( u0_u7_u7_n101 ) , .ZN( u0_u7_u7_n107 ) , .B2( u0_u7_u7_n128 ) , .B1( u0_u7_u7_n175 ) );
  INV_X1 u0_u7_u7_U23 (.A( u0_u7_u7_n101 ) , .ZN( u0_u7_u7_n165 ) );
  INV_X1 u0_u7_u7_U24 (.A( u0_u7_u7_n138 ) , .ZN( u0_u7_u7_n171 ) );
  INV_X1 u0_u7_u7_U25 (.A( u0_u7_u7_n131 ) , .ZN( u0_u7_u7_n177 ) );
  INV_X1 u0_u7_u7_U26 (.A( u0_u7_u7_n110 ) , .ZN( u0_u7_u7_n174 ) );
  NAND2_X1 u0_u7_u7_U27 (.A1( u0_u7_u7_n129 ) , .A2( u0_u7_u7_n132 ) , .ZN( u0_u7_u7_n149 ) );
  NAND2_X1 u0_u7_u7_U28 (.A1( u0_u7_u7_n113 ) , .A2( u0_u7_u7_n124 ) , .ZN( u0_u7_u7_n130 ) );
  INV_X1 u0_u7_u7_U29 (.A( u0_u7_u7_n128 ) , .ZN( u0_u7_u7_n168 ) );
  OAI21_X1 u0_u7_u7_U3 (.ZN( u0_u7_u7_n159 ) , .A( u0_u7_u7_n165 ) , .B2( u0_u7_u7_n171 ) , .B1( u0_u7_u7_n174 ) );
  INV_X1 u0_u7_u7_U30 (.A( u0_u7_u7_n148 ) , .ZN( u0_u7_u7_n169 ) );
  INV_X1 u0_u7_u7_U31 (.A( u0_u7_u7_n112 ) , .ZN( u0_u7_u7_n173 ) );
  INV_X1 u0_u7_u7_U32 (.A( u0_u7_u7_n127 ) , .ZN( u0_u7_u7_n179 ) );
  NOR2_X1 u0_u7_u7_U33 (.ZN( u0_u7_u7_n101 ) , .A2( u0_u7_u7_n150 ) , .A1( u0_u7_u7_n156 ) );
  AOI211_X1 u0_u7_u7_U34 (.B( u0_u7_u7_n154 ) , .A( u0_u7_u7_n155 ) , .C1( u0_u7_u7_n156 ) , .ZN( u0_u7_u7_n157 ) , .C2( u0_u7_u7_n172 ) );
  INV_X1 u0_u7_u7_U35 (.A( u0_u7_u7_n153 ) , .ZN( u0_u7_u7_n172 ) );
  AOI211_X1 u0_u7_u7_U36 (.B( u0_u7_u7_n139 ) , .A( u0_u7_u7_n140 ) , .C2( u0_u7_u7_n141 ) , .ZN( u0_u7_u7_n142 ) , .C1( u0_u7_u7_n156 ) );
  NAND4_X1 u0_u7_u7_U37 (.A3( u0_u7_u7_n127 ) , .A2( u0_u7_u7_n128 ) , .A1( u0_u7_u7_n129 ) , .ZN( u0_u7_u7_n141 ) , .A4( u0_u7_u7_n147 ) );
  AOI21_X1 u0_u7_u7_U38 (.A( u0_u7_u7_n137 ) , .B1( u0_u7_u7_n138 ) , .ZN( u0_u7_u7_n139 ) , .B2( u0_u7_u7_n146 ) );
  OAI22_X1 u0_u7_u7_U39 (.B1( u0_u7_u7_n136 ) , .ZN( u0_u7_u7_n140 ) , .A1( u0_u7_u7_n153 ) , .B2( u0_u7_u7_n162 ) , .A2( u0_u7_u7_n164 ) );
  INV_X1 u0_u7_u7_U4 (.A( u0_u7_u7_n149 ) , .ZN( u0_u7_u7_n175 ) );
  INV_X1 u0_u7_u7_U40 (.A( u0_u7_u7_n125 ) , .ZN( u0_u7_u7_n161 ) );
  AOI21_X1 u0_u7_u7_U41 (.ZN( u0_u7_u7_n123 ) , .B1( u0_u7_u7_n165 ) , .B2( u0_u7_u7_n177 ) , .A( u0_u7_u7_n97 ) );
  AOI21_X1 u0_u7_u7_U42 (.B2( u0_u7_u7_n113 ) , .B1( u0_u7_u7_n124 ) , .A( u0_u7_u7_n125 ) , .ZN( u0_u7_u7_n97 ) );
  INV_X1 u0_u7_u7_U43 (.A( u0_u7_u7_n152 ) , .ZN( u0_u7_u7_n162 ) );
  AOI22_X1 u0_u7_u7_U44 (.A2( u0_u7_u7_n114 ) , .ZN( u0_u7_u7_n119 ) , .B1( u0_u7_u7_n130 ) , .A1( u0_u7_u7_n156 ) , .B2( u0_u7_u7_n165 ) );
  NAND2_X1 u0_u7_u7_U45 (.A2( u0_u7_u7_n112 ) , .ZN( u0_u7_u7_n114 ) , .A1( u0_u7_u7_n175 ) );
  NOR2_X1 u0_u7_u7_U46 (.ZN( u0_u7_u7_n137 ) , .A1( u0_u7_u7_n150 ) , .A2( u0_u7_u7_n161 ) );
  AND2_X1 u0_u7_u7_U47 (.ZN( u0_u7_u7_n145 ) , .A2( u0_u7_u7_n98 ) , .A1( u0_u7_u7_n99 ) );
  AOI21_X1 u0_u7_u7_U48 (.ZN( u0_u7_u7_n105 ) , .B2( u0_u7_u7_n110 ) , .A( u0_u7_u7_n125 ) , .B1( u0_u7_u7_n147 ) );
  NAND2_X1 u0_u7_u7_U49 (.ZN( u0_u7_u7_n146 ) , .A1( u0_u7_u7_n95 ) , .A2( u0_u7_u7_n98 ) );
  INV_X1 u0_u7_u7_U5 (.A( u0_u7_u7_n154 ) , .ZN( u0_u7_u7_n178 ) );
  NAND2_X1 u0_u7_u7_U50 (.A2( u0_u7_u7_n103 ) , .ZN( u0_u7_u7_n147 ) , .A1( u0_u7_u7_n93 ) );
  NAND2_X1 u0_u7_u7_U51 (.A1( u0_u7_u7_n103 ) , .ZN( u0_u7_u7_n127 ) , .A2( u0_u7_u7_n99 ) );
  NAND2_X1 u0_u7_u7_U52 (.A2( u0_u7_u7_n102 ) , .A1( u0_u7_u7_n103 ) , .ZN( u0_u7_u7_n133 ) );
  OR2_X1 u0_u7_u7_U53 (.ZN( u0_u7_u7_n126 ) , .A2( u0_u7_u7_n152 ) , .A1( u0_u7_u7_n156 ) );
  NAND2_X1 u0_u7_u7_U54 (.ZN( u0_u7_u7_n112 ) , .A2( u0_u7_u7_n96 ) , .A1( u0_u7_u7_n99 ) );
  NAND2_X1 u0_u7_u7_U55 (.A2( u0_u7_u7_n102 ) , .ZN( u0_u7_u7_n128 ) , .A1( u0_u7_u7_n98 ) );
  INV_X1 u0_u7_u7_U56 (.A( u0_u7_u7_n150 ) , .ZN( u0_u7_u7_n164 ) );
  AND2_X1 u0_u7_u7_U57 (.ZN( u0_u7_u7_n134 ) , .A1( u0_u7_u7_n93 ) , .A2( u0_u7_u7_n98 ) );
  NAND2_X1 u0_u7_u7_U58 (.ZN( u0_u7_u7_n110 ) , .A1( u0_u7_u7_n95 ) , .A2( u0_u7_u7_n96 ) );
  NAND2_X1 u0_u7_u7_U59 (.A2( u0_u7_u7_n102 ) , .ZN( u0_u7_u7_n124 ) , .A1( u0_u7_u7_n96 ) );
  INV_X1 u0_u7_u7_U6 (.A( u0_u7_u7_n111 ) , .ZN( u0_u7_u7_n170 ) );
  NAND2_X1 u0_u7_u7_U60 (.ZN( u0_u7_u7_n132 ) , .A1( u0_u7_u7_n93 ) , .A2( u0_u7_u7_n96 ) );
  NAND2_X1 u0_u7_u7_U61 (.A2( u0_u7_u7_n103 ) , .ZN( u0_u7_u7_n131 ) , .A1( u0_u7_u7_n95 ) );
  NOR2_X1 u0_u7_u7_U62 (.A2( u0_u7_X_47 ) , .ZN( u0_u7_u7_n150 ) , .A1( u0_u7_u7_n163 ) );
  NOR2_X1 u0_u7_u7_U63 (.A2( u0_u7_X_43 ) , .A1( u0_u7_X_44 ) , .ZN( u0_u7_u7_n103 ) );
  NOR2_X1 u0_u7_u7_U64 (.A2( u0_u7_X_48 ) , .A1( u0_u7_u7_n166 ) , .ZN( u0_u7_u7_n95 ) );
  NOR2_X1 u0_u7_u7_U65 (.A2( u0_u7_X_44 ) , .A1( u0_u7_u7_n167 ) , .ZN( u0_u7_u7_n98 ) );
  NOR2_X1 u0_u7_u7_U66 (.A2( u0_u7_X_45 ) , .A1( u0_u7_X_48 ) , .ZN( u0_u7_u7_n99 ) );
  NOR2_X1 u0_u7_u7_U67 (.A2( u0_u7_X_46 ) , .A1( u0_u7_X_47 ) , .ZN( u0_u7_u7_n152 ) );
  AND2_X1 u0_u7_u7_U68 (.A1( u0_u7_X_47 ) , .ZN( u0_u7_u7_n156 ) , .A2( u0_u7_u7_n163 ) );
  NAND2_X1 u0_u7_u7_U69 (.A2( u0_u7_X_46 ) , .A1( u0_u7_X_47 ) , .ZN( u0_u7_u7_n125 ) );
  AOI211_X1 u0_u7_u7_U7 (.ZN( u0_u7_u7_n116 ) , .A( u0_u7_u7_n155 ) , .C1( u0_u7_u7_n161 ) , .C2( u0_u7_u7_n171 ) , .B( u0_u7_u7_n94 ) );
  AND2_X1 u0_u7_u7_U70 (.A2( u0_u7_X_43 ) , .A1( u0_u7_X_44 ) , .ZN( u0_u7_u7_n96 ) );
  AND2_X1 u0_u7_u7_U71 (.A2( u0_u7_X_45 ) , .A1( u0_u7_X_48 ) , .ZN( u0_u7_u7_n102 ) );
  AND2_X1 u0_u7_u7_U72 (.A1( u0_u7_X_48 ) , .A2( u0_u7_u7_n166 ) , .ZN( u0_u7_u7_n93 ) );
  INV_X1 u0_u7_u7_U73 (.A( u0_u7_X_46 ) , .ZN( u0_u7_u7_n163 ) );
  AND2_X1 u0_u7_u7_U74 (.A1( u0_u7_X_44 ) , .ZN( u0_u7_u7_n100 ) , .A2( u0_u7_u7_n167 ) );
  INV_X1 u0_u7_u7_U75 (.A( u0_u7_X_45 ) , .ZN( u0_u7_u7_n166 ) );
  INV_X1 u0_u7_u7_U76 (.A( u0_u7_X_43 ) , .ZN( u0_u7_u7_n167 ) );
  NAND4_X1 u0_u7_u7_U77 (.ZN( u0_out7_5 ) , .A4( u0_u7_u7_n108 ) , .A3( u0_u7_u7_n109 ) , .A1( u0_u7_u7_n116 ) , .A2( u0_u7_u7_n123 ) );
  AOI22_X1 u0_u7_u7_U78 (.ZN( u0_u7_u7_n109 ) , .A2( u0_u7_u7_n126 ) , .B2( u0_u7_u7_n145 ) , .B1( u0_u7_u7_n156 ) , .A1( u0_u7_u7_n171 ) );
  NOR4_X1 u0_u7_u7_U79 (.A4( u0_u7_u7_n104 ) , .A3( u0_u7_u7_n105 ) , .A2( u0_u7_u7_n106 ) , .A1( u0_u7_u7_n107 ) , .ZN( u0_u7_u7_n108 ) );
  OAI222_X1 u0_u7_u7_U8 (.C2( u0_u7_u7_n101 ) , .B2( u0_u7_u7_n111 ) , .A1( u0_u7_u7_n113 ) , .C1( u0_u7_u7_n146 ) , .A2( u0_u7_u7_n162 ) , .B1( u0_u7_u7_n164 ) , .ZN( u0_u7_u7_n94 ) );
  NAND4_X1 u0_u7_u7_U80 (.ZN( u0_out7_27 ) , .A4( u0_u7_u7_n118 ) , .A3( u0_u7_u7_n119 ) , .A2( u0_u7_u7_n120 ) , .A1( u0_u7_u7_n121 ) );
  OAI21_X1 u0_u7_u7_U81 (.ZN( u0_u7_u7_n121 ) , .B2( u0_u7_u7_n145 ) , .A( u0_u7_u7_n150 ) , .B1( u0_u7_u7_n174 ) );
  OAI21_X1 u0_u7_u7_U82 (.ZN( u0_u7_u7_n120 ) , .A( u0_u7_u7_n161 ) , .B2( u0_u7_u7_n170 ) , .B1( u0_u7_u7_n179 ) );
  NAND4_X1 u0_u7_u7_U83 (.ZN( u0_out7_21 ) , .A4( u0_u7_u7_n157 ) , .A3( u0_u7_u7_n158 ) , .A2( u0_u7_u7_n159 ) , .A1( u0_u7_u7_n160 ) );
  OAI21_X1 u0_u7_u7_U84 (.B1( u0_u7_u7_n145 ) , .ZN( u0_u7_u7_n160 ) , .A( u0_u7_u7_n161 ) , .B2( u0_u7_u7_n177 ) );
  AOI22_X1 u0_u7_u7_U85 (.B2( u0_u7_u7_n149 ) , .B1( u0_u7_u7_n150 ) , .A2( u0_u7_u7_n151 ) , .A1( u0_u7_u7_n152 ) , .ZN( u0_u7_u7_n158 ) );
  NAND4_X1 u0_u7_u7_U86 (.ZN( u0_out7_15 ) , .A4( u0_u7_u7_n142 ) , .A3( u0_u7_u7_n143 ) , .A2( u0_u7_u7_n144 ) , .A1( u0_u7_u7_n178 ) );
  OR2_X1 u0_u7_u7_U87 (.A2( u0_u7_u7_n125 ) , .A1( u0_u7_u7_n129 ) , .ZN( u0_u7_u7_n144 ) );
  AOI22_X1 u0_u7_u7_U88 (.A2( u0_u7_u7_n126 ) , .ZN( u0_u7_u7_n143 ) , .B2( u0_u7_u7_n165 ) , .B1( u0_u7_u7_n173 ) , .A1( u0_u7_u7_n174 ) );
  NAND2_X1 u0_u7_u7_U89 (.A1( u0_u7_u7_n100 ) , .ZN( u0_u7_u7_n148 ) , .A2( u0_u7_u7_n95 ) );
  INV_X1 u0_u7_u7_U9 (.A( u0_u7_u7_n133 ) , .ZN( u0_u7_u7_n176 ) );
  NAND2_X1 u0_u7_u7_U90 (.A1( u0_u7_u7_n100 ) , .ZN( u0_u7_u7_n113 ) , .A2( u0_u7_u7_n93 ) );
  NAND2_X1 u0_u7_u7_U91 (.A1( u0_u7_u7_n100 ) , .ZN( u0_u7_u7_n138 ) , .A2( u0_u7_u7_n99 ) );
  NAND2_X1 u0_u7_u7_U92 (.A1( u0_u7_u7_n100 ) , .A2( u0_u7_u7_n102 ) , .ZN( u0_u7_u7_n129 ) );
  OAI211_X1 u0_u7_u7_U93 (.B( u0_u7_u7_n122 ) , .A( u0_u7_u7_n123 ) , .C2( u0_u7_u7_n124 ) , .ZN( u0_u7_u7_n154 ) , .C1( u0_u7_u7_n162 ) );
  AOI222_X1 u0_u7_u7_U94 (.ZN( u0_u7_u7_n122 ) , .C2( u0_u7_u7_n126 ) , .C1( u0_u7_u7_n145 ) , .B1( u0_u7_u7_n161 ) , .A2( u0_u7_u7_n165 ) , .B2( u0_u7_u7_n170 ) , .A1( u0_u7_u7_n176 ) );
  NAND3_X1 u0_u7_u7_U95 (.A3( u0_u7_u7_n146 ) , .A2( u0_u7_u7_n147 ) , .A1( u0_u7_u7_n148 ) , .ZN( u0_u7_u7_n151 ) );
  NAND3_X1 u0_u7_u7_U96 (.A3( u0_u7_u7_n131 ) , .A2( u0_u7_u7_n132 ) , .A1( u0_u7_u7_n133 ) , .ZN( u0_u7_u7_n135 ) );
  INV_X1 u0_uk_U10 (.A( u0_uk_n252 ) , .ZN( u0_uk_n31 ) );
  OAI21_X1 u0_uk_U1014 (.ZN( u0_K1_37 ) , .B1( u0_uk_n129 ) , .B2( u0_uk_n714 ) , .A( u0_uk_n876 ) );
  NAND2_X1 u0_uk_U1015 (.A1( u0_key_r_50 ) , .A2( u0_uk_n17 ) , .ZN( u0_uk_n876 ) );
  OAI21_X1 u0_uk_U1020 (.ZN( u0_K14_44 ) , .B1( u0_uk_n163 ) , .B2( u0_uk_n81 ) , .A( u0_uk_n930 ) );
  NAND2_X1 u0_uk_U1021 (.A1( u0_uk_K_r12_15 ) , .A2( u0_uk_n203 ) , .ZN( u0_uk_n930 ) );
  OAI21_X1 u0_uk_U104 (.ZN( u0_K4_5 ) , .B1( u0_uk_n10 ) , .B2( u0_uk_n502 ) , .A( u0_uk_n821 ) );
  NAND2_X1 u0_uk_U105 (.A1( u0_uk_K_r2_53 ) , .ZN( u0_uk_n821 ) , .A2( u0_uk_n99 ) );
  INV_X1 u0_uk_U1062 (.A( u0_key_r_9 ) , .ZN( u0_uk_n709 ) );
  INV_X1 u0_uk_U1067 (.A( u0_key_r_23 ) , .ZN( u0_uk_n700 ) );
  INV_X1 u0_uk_U1069 (.A( u0_key_r_30 ) , .ZN( u0_uk_n693 ) );
  INV_X1 u0_uk_U1074 (.A( u0_key_r_37 ) , .ZN( u0_uk_n687 ) );
  INV_X1 u0_uk_U1077 (.A( u0_key_r_16 ) , .ZN( u0_uk_n706 ) );
  INV_X1 u0_uk_U1080 (.A( u0_key_r_2 ) , .ZN( u0_uk_n714 ) );
  OAI21_X1 u0_uk_U1089 (.ZN( u0_K16_14 ) , .B1( u0_uk_n252 ) , .B2( u0_uk_n653 ) , .A( u0_uk_n908 ) );
  OAI22_X1 u0_uk_U109 (.ZN( u0_K14_41 ) , .A1( u0_uk_n230 ) , .B2( u0_uk_n77 ) , .A2( u0_uk_n82 ) , .B1( u0_uk_n93 ) );
  NAND2_X1 u0_uk_U1090 (.A1( u0_uk_K_r14_18 ) , .A2( u0_uk_n207 ) , .ZN( u0_uk_n908 ) );
  INV_X1 u0_uk_U1107 (.ZN( u0_K1_41 ) , .A( u0_uk_n874 ) );
  AOI22_X1 u0_uk_U1108 (.B2( u0_key_r_35 ) , .A2( u0_key_r_42 ) , .B1( u0_uk_n145 ) , .A1( u0_uk_n251 ) , .ZN( u0_uk_n874 ) );
  INV_X1 u0_uk_U1119 (.ZN( u0_K2_7 ) , .A( u0_uk_n855 ) );
  OAI22_X1 u0_uk_U113 (.ZN( u0_K13_47 ) , .B2( u0_uk_n106 ) , .B1( u0_uk_n252 ) , .A2( u0_uk_n96 ) , .A1( u0_uk_n99 ) );
  INV_X1 u0_uk_U1135 (.ZN( u0_K4_2 ) , .A( u0_uk_n828 ) );
  INV_X1 u0_uk_U1143 (.ZN( u0_K13_12 ) , .A( u0_uk_n958 ) );
  AOI22_X1 u0_uk_U1144 (.B2( u0_uk_K_r11_34 ) , .A2( u0_uk_K_r11_54 ) , .A1( u0_uk_n11 ) , .B1( u0_uk_n217 ) , .ZN( u0_uk_n958 ) );
  INV_X1 u0_uk_U1159 (.ZN( u0_K13_6 ) , .A( u0_uk_n940 ) );
  OAI22_X1 u0_uk_U118 (.ZN( u0_K8_47 ) , .A1( u0_uk_n257 ) , .B1( u0_uk_n27 ) , .A2( u0_uk_n321 ) , .B2( u0_uk_n327 ) );
  OAI22_X1 u0_uk_U127 (.ZN( u0_K4_15 ) , .A1( u0_uk_n242 ) , .A2( u0_uk_n502 ) , .B2( u0_uk_n530 ) , .B1( u0_uk_n83 ) );
  INV_X1 u0_uk_U13 (.A( u0_uk_n252 ) , .ZN( u0_uk_n60 ) );
  OAI22_X1 u0_uk_U139 (.ZN( u0_K11_15 ) , .A1( u0_uk_n147 ) , .A2( u0_uk_n197 ) , .B2( u0_uk_n212 ) , .B1( u0_uk_n93 ) );
  OAI22_X1 u0_uk_U145 (.ZN( u0_K16_15 ) , .B1( u0_uk_n17 ) , .A1( u0_uk_n187 ) , .A2( u0_uk_n645 ) , .B2( u0_uk_n652 ) );
  INV_X1 u0_uk_U151 (.ZN( u0_K11_19 ) , .A( u0_uk_n1000 ) );
  INV_X1 u0_uk_U16 (.ZN( u0_uk_n110 ) , .A( u0_uk_n222 ) );
  OAI21_X1 u0_uk_U173 (.ZN( u0_K8_30 ) , .B1( u0_uk_n250 ) , .B2( u0_uk_n333 ) , .A( u0_uk_n753 ) );
  NAND2_X1 u0_uk_U174 (.A1( u0_uk_K_r6_29 ) , .A2( u0_uk_n207 ) , .ZN( u0_uk_n753 ) );
  INV_X1 u0_uk_U180 (.ZN( u0_K11_14 ) , .A( u0_uk_n1002 ) );
  INV_X1 u0_uk_U213 (.A( u0_key_r_14 ) , .ZN( u0_uk_n707 ) );
  OAI22_X1 u0_uk_U215 (.ZN( u0_K8_31 ) , .A1( u0_uk_n102 ) , .B1( u0_uk_n223 ) , .A2( u0_uk_n321 ) , .B2( u0_uk_n359 ) );
  OAI22_X1 u0_uk_U234 (.ZN( u0_K14_31 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n240 ) , .A2( u0_uk_n55 ) , .B2( u0_uk_n61 ) );
  OAI22_X1 u0_uk_U237 (.ZN( u0_K14_39 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n163 ) , .A2( u0_uk_n52 ) , .B2( u0_uk_n56 ) );
  OAI21_X1 u0_uk_U247 (.ZN( u0_K8_44 ) , .B1( u0_uk_n117 ) , .B2( u0_uk_n320 ) , .A( u0_uk_n745 ) );
  NAND2_X1 u0_uk_U248 (.A1( u0_uk_K_r6_0 ) , .A2( u0_uk_n11 ) , .ZN( u0_uk_n745 ) );
  OAI22_X1 u0_uk_U249 (.ZN( u0_K8_48 ) , .A1( u0_uk_n100 ) , .B1( u0_uk_n223 ) , .B2( u0_uk_n347 ) , .A2( u0_uk_n354 ) );
  INV_X1 u0_uk_U250 (.ZN( u0_K1_48 ) , .A( u0_uk_n870 ) );
  AOI22_X1 u0_uk_U251 (.B2( u0_key_r_21 ) , .A2( u0_key_r_28 ) , .B1( u0_uk_n145 ) , .A1( u0_uk_n213 ) , .ZN( u0_uk_n870 ) );
  INV_X1 u0_uk_U252 (.ZN( u0_K1_44 ) , .A( u0_uk_n872 ) );
  AOI22_X1 u0_uk_U253 (.B2( u0_key_r_36 ) , .A2( u0_key_r_43 ) , .B1( u0_uk_n145 ) , .A1( u0_uk_n223 ) , .ZN( u0_uk_n872 ) );
  OAI22_X1 u0_uk_U254 (.ZN( u0_K14_48 ) , .B1( u0_uk_n128 ) , .A1( u0_uk_n230 ) , .A2( u0_uk_n52 ) , .B2( u0_uk_n90 ) );
  OAI22_X1 u0_uk_U277 (.ZN( u0_K16_6 ) , .B1( u0_uk_n145 ) , .A1( u0_uk_n155 ) , .A2( u0_uk_n639 ) , .B2( u0_uk_n644 ) );
  BUF_X1 u0_uk_U28 (.Z( u0_uk_n147 ) , .A( u0_uk_n250 ) );
  INV_X1 u0_uk_U297 (.ZN( u0_K1_26 ) , .A( u0_uk_n883 ) );
  AOI22_X1 u0_uk_U298 (.B2( u0_key_r_31 ) , .A2( u0_key_r_51 ) , .A1( u0_uk_n146 ) , .B1( u0_uk_n207 ) , .ZN( u0_uk_n883 ) );
  BUF_X1 u0_uk_U31 (.Z( u0_uk_n155 ) , .A( u0_uk_n223 ) );
  OAI22_X1 u0_uk_U318 (.ZN( u0_K8_26 ) , .A1( u0_uk_n102 ) , .B1( u0_uk_n222 ) , .B2( u0_uk_n348 ) , .A2( u0_uk_n355 ) );
  BUF_X1 u0_uk_U34 (.Z( u0_uk_n164 ) , .A( u0_uk_n214 ) );
  INV_X1 u0_uk_U345 (.ZN( u0_K4_4 ) , .A( u0_uk_n822 ) );
  AOI22_X1 u0_uk_U346 (.B2( u0_uk_K_r2_13 ) , .A2( u0_uk_K_r2_18 ) , .B1( u0_uk_n203 ) , .ZN( u0_uk_n822 ) , .A1( u0_uk_n94 ) );
  BUF_X1 u0_uk_U40 (.Z( u0_uk_n230 ) , .A( u0_uk_n257 ) );
  OAI22_X1 u0_uk_U401 (.ZN( u0_K4_16 ) , .B1( u0_uk_n128 ) , .A1( u0_uk_n238 ) , .A2( u0_uk_n525 ) , .B2( u0_uk_n529 ) );
  OAI22_X1 u0_uk_U406 (.ZN( u0_K13_9 ) , .A2( u0_uk_n115 ) , .B2( u0_uk_n127 ) , .A1( u0_uk_n230 ) , .B1( u0_uk_n93 ) );
  BUF_X1 u0_uk_U42 (.Z( u0_uk_n238 ) , .A( u0_uk_n252 ) );
  OAI22_X1 u0_uk_U421 (.ZN( u0_K4_9 ) , .A1( u0_uk_n146 ) , .B1( u0_uk_n217 ) , .A2( u0_uk_n519 ) , .B2( u0_uk_n529 ) );
  OAI22_X1 u0_uk_U429 (.ZN( u0_K16_9 ) , .B1( u0_uk_n141 ) , .A1( u0_uk_n187 ) , .A2( u0_uk_n630 ) , .B2( u0_uk_n637 ) );
  OAI22_X1 u0_uk_U430 (.ZN( u0_K16_16 ) , .B1( u0_uk_n17 ) , .A1( u0_uk_n187 ) , .A2( u0_uk_n644 ) , .B2( u0_uk_n651 ) );
  OAI22_X1 u0_uk_U444 (.ZN( u0_K14_33 ) , .A1( u0_uk_n230 ) , .A2( u0_uk_n55 ) , .B2( u0_uk_n73 ) , .B1( u0_uk_n94 ) );
  OAI22_X1 u0_uk_U451 (.ZN( u0_K14_37 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n231 ) , .A2( u0_uk_n67 ) , .B2( u0_uk_n73 ) );
  OAI22_X1 u0_uk_U469 (.ZN( u0_K1_29 ) , .A1( u0_uk_n142 ) , .B1( u0_uk_n188 ) , .A2( u0_uk_n700 ) , .B2( u0_uk_n706 ) );
  BUF_X1 u0_uk_U48 (.Z( u0_uk_n222 ) , .A( u0_uk_n250 ) );
  BUF_X1 u0_uk_U49 (.Z( u0_uk_n231 ) , .A( u0_uk_n250 ) );
  INV_X1 u0_uk_U506 (.ZN( u0_K8_29 ) , .A( u0_uk_n755 ) );
  INV_X1 u0_uk_U508 (.ZN( u0_K11_17 ) , .A( u0_uk_n1001 ) );
  OAI21_X1 u0_uk_U513 (.ZN( u0_K4_17 ) , .B1( u0_uk_n250 ) , .B2( u0_uk_n519 ) , .A( u0_uk_n838 ) );
  NAND2_X1 u0_uk_U514 (.A1( u0_uk_K_r2_27 ) , .A2( u0_uk_n208 ) , .ZN( u0_uk_n838 ) );
  BUF_X1 u0_uk_U52 (.Z( u0_uk_n207 ) , .A( u0_uk_n217 ) );
  OAI22_X1 u0_uk_U526 (.ZN( u0_K4_12 ) , .A1( u0_uk_n10 ) , .B1( u0_uk_n161 ) , .A2( u0_uk_n497 ) , .B2( u0_uk_n517 ) );
  OAI22_X1 u0_uk_U531 (.ZN( u0_K1_36 ) , .A1( u0_uk_n128 ) , .B1( u0_uk_n188 ) , .A2( u0_uk_n693 ) , .B2( u0_uk_n700 ) );
  OAI21_X1 u0_uk_U532 (.ZN( u0_K16_12 ) , .B1( u0_uk_n252 ) , .B2( u0_uk_n660 ) , .A( u0_uk_n910 ) );
  NAND2_X1 u0_uk_U533 (.A1( u0_uk_K_r14_12 ) , .A2( u0_uk_n207 ) , .ZN( u0_uk_n910 ) );
  OAI22_X1 u0_uk_U545 (.ZN( u0_K14_36 ) , .A1( u0_uk_n230 ) , .A2( u0_uk_n50 ) , .B2( u0_uk_n88 ) , .B1( u0_uk_n93 ) );
  OAI22_X1 u0_uk_U549 (.ZN( u0_K1_38 ) , .A1( u0_uk_n118 ) , .B1( u0_uk_n188 ) , .A2( u0_uk_n687 ) , .B2( u0_uk_n693 ) );
  BUF_X1 u0_uk_U55 (.A( u0_uk_n250 ) , .Z( u0_uk_n252 ) );
  BUF_X1 u0_uk_U56 (.Z( u0_uk_n250 ) , .A( u0_uk_n257 ) );
  OAI22_X1 u0_uk_U571 (.ZN( u0_K16_10 ) , .A1( u0_uk_n155 ) , .B1( u0_uk_n17 ) , .A2( u0_uk_n636 ) , .B2( u0_uk_n639 ) );
  INV_X1 u0_uk_U577 (.ZN( u0_K13_10 ) , .A( u0_uk_n960 ) );
  INV_X1 u0_uk_U584 (.ZN( u0_K4_10 ) , .A( u0_uk_n839 ) );
  INV_X1 u0_uk_U592 (.ZN( u0_K11_22 ) , .A( u0_uk_n997 ) );
  AOI22_X1 u0_uk_U593 (.B2( u0_uk_K_r9_13 ) , .A2( u0_uk_K_r9_19 ) , .B1( u0_uk_n146 ) , .A1( u0_uk_n251 ) , .ZN( u0_uk_n997 ) );
  OAI22_X1 u0_uk_U605 (.ZN( u0_K8_35 ) , .A1( u0_uk_n242 ) , .B1( u0_uk_n31 ) , .A2( u0_uk_n341 ) , .B2( u0_uk_n347 ) );
  INV_X1 u0_uk_U612 (.ZN( u0_K14_35 ) , .A( u0_uk_n933 ) );
  INV_X1 u0_uk_U62 (.ZN( u0_K8_34 ) , .A( u0_uk_n752 ) );
  INV_X1 u0_uk_U620 (.ZN( u0_K1_35 ) , .A( u0_uk_n877 ) );
  AOI22_X1 u0_uk_U621 (.B2( u0_key_r_28 ) , .A2( u0_key_r_35 ) , .B1( u0_uk_n146 ) , .A1( u0_uk_n161 ) , .ZN( u0_uk_n877 ) );
  INV_X1 u0_uk_U628 (.ZN( u0_K13_11 ) , .A( u0_uk_n959 ) );
  AOI22_X1 u0_uk_U629 (.B2( u0_uk_K_r11_17 ) , .A2( u0_uk_K_r11_54 ) , .B1( u0_uk_n129 ) , .A1( u0_uk_n240 ) , .ZN( u0_uk_n959 ) );
  AOI22_X1 u0_uk_U63 (.B2( u0_uk_K_r6_14 ) , .A2( u0_uk_K_r6_21 ) , .A1( u0_uk_n141 ) , .B1( u0_uk_n202 ) , .ZN( u0_uk_n752 ) );
  INV_X1 u0_uk_U65 (.ZN( u0_K14_34 ) , .A( u0_uk_n934 ) );
  OAI22_X1 u0_uk_U650 (.ZN( u0_K14_43 ) , .B1( u0_uk_n203 ) , .A2( u0_uk_n56 ) , .B2( u0_uk_n59 ) , .A1( u0_uk_n60 ) );
  OAI21_X1 u0_uk_U662 (.ZN( u0_K14_45 ) , .B1( u0_uk_n217 ) , .B2( u0_uk_n58 ) , .A( u0_uk_n929 ) );
  NAND2_X1 u0_uk_U663 (.A1( u0_uk_K_r12_16 ) , .A2( u0_uk_n252 ) , .ZN( u0_uk_n929 ) );
  OAI21_X1 u0_uk_U664 (.ZN( u0_K13_43 ) , .B1( u0_uk_n252 ) , .A( u0_uk_n943 ) , .B2( u0_uk_n96 ) );
  NAND2_X1 u0_uk_U665 (.A1( u0_uk_K_r11_29 ) , .A2( u0_uk_n207 ) , .ZN( u0_uk_n943 ) );
  OAI22_X1 u0_uk_U677 (.ZN( u0_K16_3 ) , .B1( u0_uk_n102 ) , .A1( u0_uk_n187 ) , .A2( u0_uk_n652 ) , .B2( u0_uk_n660 ) );
  OAI22_X1 u0_uk_U684 (.ZN( u0_K4_7 ) , .B1( u0_uk_n202 ) , .B2( u0_uk_n531 ) , .A2( u0_uk_n535 ) , .A1( u0_uk_n99 ) );
  OAI22_X1 u0_uk_U685 (.ZN( u0_K16_7 ) , .B1( u0_uk_n117 ) , .A1( u0_uk_n155 ) , .A2( u0_uk_n651 ) , .B2( u0_uk_n659 ) );
  INV_X1 u0_uk_U697 (.ZN( u0_K8_43 ) , .A( u0_uk_n746 ) );
  OAI22_X1 u0_uk_U701 (.ZN( u0_K8_25 ) , .A1( u0_uk_n161 ) , .A2( u0_uk_n320 ) , .B2( u0_uk_n325 ) , .B1( u0_uk_n60 ) );
  INV_X1 u0_uk_U704 (.ZN( u0_K13_7 ) , .A( u0_uk_n939 ) );
  OAI22_X1 u0_uk_U718 (.ZN( u0_K8_32 ) , .A1( u0_uk_n213 ) , .B1( u0_uk_n27 ) , .A2( u0_uk_n325 ) , .B2( u0_uk_n332 ) );
  OAI22_X1 u0_uk_U724 (.ZN( u0_K14_32 ) , .A1( u0_uk_n164 ) , .A2( u0_uk_n51 ) , .B2( u0_uk_n89 ) , .B1( u0_uk_n94 ) );
  OAI22_X1 u0_uk_U74 (.ZN( u0_K16_23 ) , .A1( u0_uk_n164 ) , .A2( u0_uk_n640 ) , .B2( u0_uk_n645 ) , .B1( u0_uk_n92 ) );
  INV_X1 u0_uk_U742 (.ZN( u0_K1_42 ) , .A( u0_uk_n873 ) );
  AOI22_X1 u0_uk_U743 (.B2( u0_key_r_31 ) , .A2( u0_key_r_38 ) , .B1( u0_uk_n145 ) , .A1( u0_uk_n251 ) , .ZN( u0_uk_n873 ) );
  OAI22_X1 u0_uk_U749 (.ZN( u0_K8_27 ) , .B1( u0_uk_n128 ) , .A1( u0_uk_n257 ) , .A2( u0_uk_n354 ) , .B2( u0_uk_n359 ) );
  OAI21_X1 u0_uk_U75 (.ZN( u0_K11_23 ) , .B2( u0_uk_n190 ) , .B1( u0_uk_n250 ) , .A( u0_uk_n996 ) );
  OAI22_X1 u0_uk_U752 (.ZN( u0_K11_13 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n164 ) , .A2( u0_uk_n196 ) , .B2( u0_uk_n200 ) );
  NAND2_X1 u0_uk_U76 (.A1( u0_uk_K_r9_27 ) , .A2( u0_uk_n202 ) , .ZN( u0_uk_n996 ) );
  OAI22_X1 u0_uk_U772 (.ZN( u0_K4_13 ) , .B1( u0_uk_n240 ) , .B2( u0_uk_n530 ) , .A2( u0_uk_n534 ) , .A1( u0_uk_n60 ) );
  INV_X1 u0_uk_U786 (.ZN( u0_K6_21 ) , .A( u0_uk_n797 ) );
  OAI21_X1 u0_uk_U788 (.ZN( u0_K16_13 ) , .B1( u0_uk_n147 ) , .B2( u0_uk_n631 ) , .A( u0_uk_n909 ) );
  NAND2_X1 u0_uk_U789 (.A1( u0_uk_K_r14_46 ) , .A2( u0_uk_n208 ) , .ZN( u0_uk_n909 ) );
  INV_X1 u0_uk_U794 (.ZN( u0_K1_27 ) , .A( u0_uk_n882 ) );
  AOI22_X1 u0_uk_U795 (.B2( u0_key_r_14 ) , .A2( u0_key_r_21 ) , .B1( u0_uk_n146 ) , .A1( u0_uk_n238 ) , .ZN( u0_uk_n882 ) );
  OAI22_X1 u0_uk_U798 (.ZN( u0_K16_1 ) , .A1( u0_uk_n155 ) , .B1( u0_uk_n17 ) , .A2( u0_uk_n637 ) , .B2( u0_uk_n640 ) );
  OAI21_X1 u0_uk_U802 (.ZN( u0_K4_1 ) , .B1( u0_uk_n252 ) , .B2( u0_uk_n535 ) , .A( u0_uk_n836 ) );
  NAND2_X1 u0_uk_U803 (.A1( u0_uk_K_r2_25 ) , .A2( u0_uk_n207 ) , .ZN( u0_uk_n836 ) );
  OAI21_X1 u0_uk_U804 (.ZN( u0_K4_18 ) , .B2( u0_uk_n510 ) , .A( u0_uk_n837 ) , .B1( u0_uk_n92 ) );
  NAND2_X1 u0_uk_U805 (.A1( u0_uk_K_r2_20 ) , .A2( u0_uk_n31 ) , .ZN( u0_uk_n837 ) );
  OAI22_X1 u0_uk_U822 (.ZN( u0_K16_20 ) , .A1( u0_uk_n155 ) , .B1( u0_uk_n17 ) , .A2( u0_uk_n629 ) , .B2( u0_uk_n636 ) );
  OAI22_X1 u0_uk_U824 (.ZN( u0_K8_20 ) , .B1( u0_uk_n110 ) , .A1( u0_uk_n213 ) , .A2( u0_uk_n331 ) , .B2( u0_uk_n337 ) );
  INV_X1 u0_uk_U827 (.ZN( u0_K6_18 ) , .A( u0_uk_n799 ) );
  INV_X1 u0_uk_U829 (.ZN( u0_K11_20 ) , .A( u0_uk_n999 ) );
  OAI21_X1 u0_uk_U835 (.ZN( u0_K13_1 ) , .B2( u0_uk_n131 ) , .B1( u0_uk_n31 ) , .A( u0_uk_n952 ) );
  NAND2_X1 u0_uk_U836 (.A1( u0_uk_K_r11_25 ) , .A2( u0_uk_n11 ) , .ZN( u0_uk_n952 ) );
  OAI22_X1 u0_uk_U843 (.ZN( u0_K1_43 ) , .B1( u0_uk_n109 ) , .A1( u0_uk_n164 ) , .B2( u0_uk_n706 ) , .A2( u0_uk_n709 ) );
  OAI21_X1 u0_uk_U860 (.ZN( u0_K16_2 ) , .B1( u0_uk_n128 ) , .B2( u0_uk_n668 ) , .A( u0_uk_n903 ) );
  NAND2_X1 u0_uk_U861 (.A1( u0_uk_K_r14_11 ) , .A2( u0_uk_n118 ) , .ZN( u0_uk_n903 ) );
  OAI22_X1 u0_uk_U884 (.ZN( u0_K4_11 ) , .B1( u0_uk_n117 ) , .A1( u0_uk_n164 ) , .A2( u0_uk_n497 ) , .B2( u0_uk_n525 ) );
  INV_X1 u0_uk_U9 (.A( u0_uk_n147 ) , .ZN( u0_uk_n17 ) );
  OAI22_X1 u0_uk_U909 (.ZN( u0_K8_21 ) , .B1( u0_uk_n102 ) , .A1( u0_uk_n257 ) , .A2( u0_uk_n330 ) , .B2( u0_uk_n336 ) );
  OAI22_X1 u0_uk_U914 (.ZN( u0_K4_14 ) , .A1( u0_uk_n164 ) , .A2( u0_uk_n510 ) , .B2( u0_uk_n536 ) , .B1( u0_uk_n99 ) );
  OAI22_X1 u0_uk_U933 (.ZN( u0_K11_16 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n182 ) , .A2( u0_uk_n190 ) , .B2( u0_uk_n196 ) );
  OAI22_X1 u0_uk_U94 (.ZN( u0_K16_5 ) , .A1( u0_uk_n118 ) , .B1( u0_uk_n187 ) , .B2( u0_uk_n664 ) , .A2( u0_uk_n667 ) );
  OAI22_X1 u0_uk_U942 (.ZN( u0_K11_24 ) , .A1( u0_uk_n109 ) , .A2( u0_uk_n201 ) , .B2( u0_uk_n206 ) , .B1( u0_uk_n222 ) );
  OAI22_X1 u0_uk_U944 (.ZN( u0_K8_24 ) , .A1( u0_uk_n102 ) , .B1( u0_uk_n213 ) , .A2( u0_uk_n318 ) , .B2( u0_uk_n358 ) );
  OAI22_X1 u0_uk_U947 (.ZN( u0_K14_47 ) , .A1( u0_uk_n17 ) , .B1( u0_uk_n231 ) , .A2( u0_uk_n58 ) , .B2( u0_uk_n68 ) );
  OAI22_X1 u0_uk_U952 (.ZN( u0_K13_4 ) , .A1( u0_uk_n117 ) , .A2( u0_uk_n121 ) , .B2( u0_uk_n126 ) , .B1( u0_uk_n214 ) );
  OAI22_X1 u0_uk_U959 (.ZN( u0_K11_18 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n214 ) , .A2( u0_uk_n215 ) , .B2( u0_uk_n221 ) );
  OAI22_X1 u0_uk_U966 (.ZN( u0_K14_38 ) , .A1( u0_uk_n141 ) , .B1( u0_uk_n250 ) , .B2( u0_uk_n65 ) , .A2( u0_uk_n81 ) );
  INV_X1 u0_uk_U98 (.ZN( u0_K13_5 ) , .A( u0_uk_n941 ) );
  OAI22_X1 u0_uk_U988 (.ZN( u0_K6_25 ) , .A1( u0_uk_n102 ) , .B1( u0_uk_n214 ) , .A2( u0_uk_n418 ) , .B2( u0_uk_n434 ) );
  AOI22_X1 u0_uk_U99 (.B2( u0_uk_K_r11_48 ) , .A2( u0_uk_K_r11_53 ) , .B1( u0_uk_n141 ) , .A1( u0_uk_n220 ) , .ZN( u0_uk_n941 ) );
  OAI22_X1 u0_uk_U991 (.ZN( u0_K1_34 ) , .A1( u0_uk_n118 ) , .B1( u0_uk_n188 ) , .A2( u0_uk_n709 ) , .B2( u0_uk_n714 ) );
  XOR2_X1 u1_u0_U16 (.B( u1_K1_3 ) , .A( u1_desIn_r_15 ) , .Z( u1_u0_X_3 ) );
  XOR2_X1 u1_u0_U35 (.B( u1_K1_22 ) , .A( u1_desIn_r_53 ) , .Z( u1_u0_X_22 ) );
  XOR2_X1 u1_u0_U36 (.B( u1_K1_21 ) , .A( u1_desIn_r_45 ) , .Z( u1_u0_X_21 ) );
  XOR2_X1 u1_u0_U6 (.B( u1_K1_4 ) , .A( u1_desIn_r_23 ) , .Z( u1_u0_X_4 ) );
  NAND2_X1 u1_u0_u0_U10 (.ZN( u1_u0_u0_n113 ) , .A1( u1_u0_u0_n139 ) , .A2( u1_u0_u0_n149 ) );
  AND3_X1 u1_u0_u0_U11 (.A2( u1_u0_u0_n112 ) , .ZN( u1_u0_u0_n127 ) , .A3( u1_u0_u0_n130 ) , .A1( u1_u0_u0_n148 ) );
  AND2_X1 u1_u0_u0_U12 (.ZN( u1_u0_u0_n107 ) , .A1( u1_u0_u0_n130 ) , .A2( u1_u0_u0_n140 ) );
  AND2_X1 u1_u0_u0_U13 (.A2( u1_u0_u0_n129 ) , .A1( u1_u0_u0_n130 ) , .ZN( u1_u0_u0_n151 ) );
  AND2_X1 u1_u0_u0_U14 (.A1( u1_u0_u0_n108 ) , .A2( u1_u0_u0_n125 ) , .ZN( u1_u0_u0_n145 ) );
  INV_X1 u1_u0_u0_U15 (.A( u1_u0_u0_n143 ) , .ZN( u1_u0_u0_n173 ) );
  NOR2_X1 u1_u0_u0_U16 (.A2( u1_u0_u0_n136 ) , .ZN( u1_u0_u0_n147 ) , .A1( u1_u0_u0_n160 ) );
  INV_X1 u1_u0_u0_U17 (.ZN( u1_u0_u0_n172 ) , .A( u1_u0_u0_n88 ) );
  OAI222_X1 u1_u0_u0_U18 (.C1( u1_u0_u0_n108 ) , .A1( u1_u0_u0_n125 ) , .B2( u1_u0_u0_n128 ) , .B1( u1_u0_u0_n144 ) , .A2( u1_u0_u0_n158 ) , .C2( u1_u0_u0_n161 ) , .ZN( u1_u0_u0_n88 ) );
  AOI21_X1 u1_u0_u0_U19 (.B1( u1_u0_u0_n103 ) , .ZN( u1_u0_u0_n132 ) , .A( u1_u0_u0_n165 ) , .B2( u1_u0_u0_n93 ) );
  INV_X1 u1_u0_u0_U20 (.A( u1_u0_u0_n142 ) , .ZN( u1_u0_u0_n165 ) );
  OAI22_X1 u1_u0_u0_U21 (.B1( u1_u0_u0_n125 ) , .ZN( u1_u0_u0_n126 ) , .A1( u1_u0_u0_n138 ) , .A2( u1_u0_u0_n146 ) , .B2( u1_u0_u0_n147 ) );
  OAI22_X1 u1_u0_u0_U22 (.B1( u1_u0_u0_n131 ) , .A1( u1_u0_u0_n144 ) , .B2( u1_u0_u0_n147 ) , .A2( u1_u0_u0_n90 ) , .ZN( u1_u0_u0_n91 ) );
  AND3_X1 u1_u0_u0_U23 (.A3( u1_u0_u0_n121 ) , .A2( u1_u0_u0_n125 ) , .A1( u1_u0_u0_n148 ) , .ZN( u1_u0_u0_n90 ) );
  INV_X1 u1_u0_u0_U24 (.A( u1_u0_u0_n136 ) , .ZN( u1_u0_u0_n161 ) );
  AOI22_X1 u1_u0_u0_U25 (.B2( u1_u0_u0_n109 ) , .A2( u1_u0_u0_n110 ) , .ZN( u1_u0_u0_n111 ) , .B1( u1_u0_u0_n118 ) , .A1( u1_u0_u0_n160 ) );
  INV_X1 u1_u0_u0_U26 (.A( u1_u0_u0_n118 ) , .ZN( u1_u0_u0_n158 ) );
  AOI21_X1 u1_u0_u0_U27 (.B1( u1_u0_u0_n127 ) , .B2( u1_u0_u0_n129 ) , .A( u1_u0_u0_n138 ) , .ZN( u1_u0_u0_n96 ) );
  AOI21_X1 u1_u0_u0_U28 (.ZN( u1_u0_u0_n104 ) , .B1( u1_u0_u0_n107 ) , .B2( u1_u0_u0_n141 ) , .A( u1_u0_u0_n144 ) );
  NAND2_X1 u1_u0_u0_U29 (.A1( u1_u0_u0_n100 ) , .A2( u1_u0_u0_n103 ) , .ZN( u1_u0_u0_n125 ) );
  INV_X1 u1_u0_u0_U3 (.A( u1_u0_u0_n113 ) , .ZN( u1_u0_u0_n166 ) );
  NAND2_X1 u1_u0_u0_U30 (.A2( u1_u0_u0_n100 ) , .ZN( u1_u0_u0_n131 ) , .A1( u1_u0_u0_n92 ) );
  NAND2_X1 u1_u0_u0_U31 (.A2( u1_u0_u0_n102 ) , .ZN( u1_u0_u0_n114 ) , .A1( u1_u0_u0_n92 ) );
  NOR2_X1 u1_u0_u0_U32 (.A1( u1_u0_u0_n120 ) , .ZN( u1_u0_u0_n143 ) , .A2( u1_u0_u0_n167 ) );
  OAI221_X1 u1_u0_u0_U33 (.C1( u1_u0_u0_n112 ) , .ZN( u1_u0_u0_n120 ) , .B1( u1_u0_u0_n138 ) , .B2( u1_u0_u0_n141 ) , .C2( u1_u0_u0_n147 ) , .A( u1_u0_u0_n172 ) );
  AOI21_X1 u1_u0_u0_U34 (.ZN( u1_u0_u0_n116 ) , .B2( u1_u0_u0_n142 ) , .A( u1_u0_u0_n144 ) , .B1( u1_u0_u0_n166 ) );
  INV_X1 u1_u0_u0_U35 (.A( u1_u0_u0_n138 ) , .ZN( u1_u0_u0_n160 ) );
  NAND2_X1 u1_u0_u0_U36 (.A2( u1_u0_u0_n102 ) , .A1( u1_u0_u0_n103 ) , .ZN( u1_u0_u0_n149 ) );
  NAND2_X1 u1_u0_u0_U37 (.ZN( u1_u0_u0_n112 ) , .A2( u1_u0_u0_n92 ) , .A1( u1_u0_u0_n93 ) );
  OR3_X1 u1_u0_u0_U38 (.A3( u1_u0_u0_n152 ) , .A2( u1_u0_u0_n153 ) , .A1( u1_u0_u0_n154 ) , .ZN( u1_u0_u0_n155 ) );
  AOI21_X1 u1_u0_u0_U39 (.B2( u1_u0_u0_n150 ) , .B1( u1_u0_u0_n151 ) , .ZN( u1_u0_u0_n152 ) , .A( u1_u0_u0_n158 ) );
  NOR2_X1 u1_u0_u0_U4 (.A1( u1_u0_u0_n108 ) , .ZN( u1_u0_u0_n123 ) , .A2( u1_u0_u0_n158 ) );
  AOI21_X1 u1_u0_u0_U40 (.A( u1_u0_u0_n144 ) , .B2( u1_u0_u0_n145 ) , .B1( u1_u0_u0_n146 ) , .ZN( u1_u0_u0_n154 ) );
  AOI21_X1 u1_u0_u0_U41 (.A( u1_u0_u0_n147 ) , .B2( u1_u0_u0_n148 ) , .B1( u1_u0_u0_n149 ) , .ZN( u1_u0_u0_n153 ) );
  INV_X1 u1_u0_u0_U42 (.ZN( u1_u0_u0_n171 ) , .A( u1_u0_u0_n99 ) );
  OAI211_X1 u1_u0_u0_U43 (.C2( u1_u0_u0_n140 ) , .C1( u1_u0_u0_n161 ) , .A( u1_u0_u0_n169 ) , .B( u1_u0_u0_n98 ) , .ZN( u1_u0_u0_n99 ) );
  AOI211_X1 u1_u0_u0_U44 (.C1( u1_u0_u0_n118 ) , .A( u1_u0_u0_n123 ) , .B( u1_u0_u0_n96 ) , .C2( u1_u0_u0_n97 ) , .ZN( u1_u0_u0_n98 ) );
  INV_X1 u1_u0_u0_U45 (.ZN( u1_u0_u0_n169 ) , .A( u1_u0_u0_n91 ) );
  NOR2_X1 u1_u0_u0_U46 (.A2( u1_u0_X_2 ) , .ZN( u1_u0_u0_n103 ) , .A1( u1_u0_u0_n164 ) );
  NOR2_X1 u1_u0_u0_U47 (.A2( u1_u0_X_4 ) , .A1( u1_u0_X_5 ) , .ZN( u1_u0_u0_n118 ) );
  NAND2_X1 u1_u0_u0_U48 (.A2( u1_u0_X_4 ) , .A1( u1_u0_X_5 ) , .ZN( u1_u0_u0_n144 ) );
  NOR2_X1 u1_u0_u0_U49 (.A2( u1_u0_X_5 ) , .ZN( u1_u0_u0_n136 ) , .A1( u1_u0_u0_n159 ) );
  AOI21_X1 u1_u0_u0_U5 (.B2( u1_u0_u0_n131 ) , .ZN( u1_u0_u0_n134 ) , .B1( u1_u0_u0_n151 ) , .A( u1_u0_u0_n158 ) );
  NAND2_X1 u1_u0_u0_U50 (.A1( u1_u0_X_5 ) , .ZN( u1_u0_u0_n138 ) , .A2( u1_u0_u0_n159 ) );
  AND2_X1 u1_u0_u0_U51 (.A2( u1_u0_X_3 ) , .A1( u1_u0_X_6 ) , .ZN( u1_u0_u0_n102 ) );
  AND2_X1 u1_u0_u0_U52 (.A1( u1_u0_X_6 ) , .A2( u1_u0_u0_n162 ) , .ZN( u1_u0_u0_n93 ) );
  INV_X1 u1_u0_u0_U53 (.A( u1_u0_X_4 ) , .ZN( u1_u0_u0_n159 ) );
  INV_X1 u1_u0_u0_U54 (.A( u1_u0_X_2 ) , .ZN( u1_u0_u0_n163 ) );
  INV_X1 u1_u0_u0_U55 (.A( u1_u0_X_3 ) , .ZN( u1_u0_u0_n162 ) );
  INV_X1 u1_u0_u0_U56 (.A( u1_u0_u0_n126 ) , .ZN( u1_u0_u0_n168 ) );
  AOI211_X1 u1_u0_u0_U57 (.B( u1_u0_u0_n133 ) , .A( u1_u0_u0_n134 ) , .C2( u1_u0_u0_n135 ) , .C1( u1_u0_u0_n136 ) , .ZN( u1_u0_u0_n137 ) );
  OR4_X1 u1_u0_u0_U58 (.ZN( u1_out0_17 ) , .A4( u1_u0_u0_n122 ) , .A2( u1_u0_u0_n123 ) , .A1( u1_u0_u0_n124 ) , .A3( u1_u0_u0_n170 ) );
  AOI21_X1 u1_u0_u0_U59 (.B2( u1_u0_u0_n107 ) , .ZN( u1_u0_u0_n124 ) , .B1( u1_u0_u0_n128 ) , .A( u1_u0_u0_n161 ) );
  OAI21_X1 u1_u0_u0_U6 (.B1( u1_u0_u0_n150 ) , .B2( u1_u0_u0_n158 ) , .A( u1_u0_u0_n172 ) , .ZN( u1_u0_u0_n89 ) );
  INV_X1 u1_u0_u0_U60 (.A( u1_u0_u0_n111 ) , .ZN( u1_u0_u0_n170 ) );
  OR4_X1 u1_u0_u0_U61 (.ZN( u1_out0_31 ) , .A4( u1_u0_u0_n155 ) , .A2( u1_u0_u0_n156 ) , .A1( u1_u0_u0_n157 ) , .A3( u1_u0_u0_n173 ) );
  AOI21_X1 u1_u0_u0_U62 (.A( u1_u0_u0_n138 ) , .B2( u1_u0_u0_n139 ) , .B1( u1_u0_u0_n140 ) , .ZN( u1_u0_u0_n157 ) );
  AOI21_X1 u1_u0_u0_U63 (.B2( u1_u0_u0_n141 ) , .B1( u1_u0_u0_n142 ) , .ZN( u1_u0_u0_n156 ) , .A( u1_u0_u0_n161 ) );
  INV_X1 u1_u0_u0_U64 (.ZN( u1_u0_u0_n174 ) , .A( u1_u0_u0_n89 ) );
  AOI211_X1 u1_u0_u0_U65 (.B( u1_u0_u0_n104 ) , .A( u1_u0_u0_n105 ) , .ZN( u1_u0_u0_n106 ) , .C2( u1_u0_u0_n113 ) , .C1( u1_u0_u0_n160 ) );
  AOI211_X1 u1_u0_u0_U66 (.B( u1_u0_u0_n115 ) , .A( u1_u0_u0_n116 ) , .C2( u1_u0_u0_n117 ) , .C1( u1_u0_u0_n118 ) , .ZN( u1_u0_u0_n119 ) );
  NAND2_X1 u1_u0_u0_U67 (.A2( u1_u0_u0_n101 ) , .ZN( u1_u0_u0_n121 ) , .A1( u1_u0_u0_n93 ) );
  NAND2_X1 u1_u0_u0_U68 (.A1( u1_u0_u0_n101 ) , .A2( u1_u0_u0_n102 ) , .ZN( u1_u0_u0_n150 ) );
  NOR2_X1 u1_u0_u0_U69 (.A2( u1_u0_X_1 ) , .A1( u1_u0_X_2 ) , .ZN( u1_u0_u0_n92 ) );
  AOI21_X1 u1_u0_u0_U7 (.B1( u1_u0_u0_n114 ) , .ZN( u1_u0_u0_n115 ) , .B2( u1_u0_u0_n129 ) , .A( u1_u0_u0_n161 ) );
  NAND2_X1 u1_u0_u0_U70 (.A2( u1_u0_u0_n100 ) , .A1( u1_u0_u0_n101 ) , .ZN( u1_u0_u0_n139 ) );
  NOR2_X1 u1_u0_u0_U71 (.A2( u1_u0_X_1 ) , .ZN( u1_u0_u0_n101 ) , .A1( u1_u0_u0_n163 ) );
  INV_X1 u1_u0_u0_U72 (.A( u1_u0_X_1 ) , .ZN( u1_u0_u0_n164 ) );
  NAND2_X1 u1_u0_u0_U73 (.A1( u1_u0_u0_n102 ) , .ZN( u1_u0_u0_n128 ) , .A2( u1_u0_u0_n95 ) );
  NAND2_X1 u1_u0_u0_U74 (.A1( u1_u0_u0_n100 ) , .ZN( u1_u0_u0_n129 ) , .A2( u1_u0_u0_n95 ) );
  NAND2_X1 u1_u0_u0_U75 (.ZN( u1_u0_u0_n148 ) , .A1( u1_u0_u0_n93 ) , .A2( u1_u0_u0_n95 ) );
  OAI221_X1 u1_u0_u0_U76 (.C1( u1_u0_u0_n121 ) , .ZN( u1_u0_u0_n122 ) , .B2( u1_u0_u0_n127 ) , .A( u1_u0_u0_n143 ) , .B1( u1_u0_u0_n144 ) , .C2( u1_u0_u0_n147 ) );
  NOR2_X1 u1_u0_u0_U77 (.A1( u1_u0_u0_n163 ) , .A2( u1_u0_u0_n164 ) , .ZN( u1_u0_u0_n95 ) );
  AOI21_X1 u1_u0_u0_U78 (.B1( u1_u0_u0_n132 ) , .ZN( u1_u0_u0_n133 ) , .A( u1_u0_u0_n144 ) , .B2( u1_u0_u0_n166 ) );
  OAI22_X1 u1_u0_u0_U79 (.ZN( u1_u0_u0_n105 ) , .A2( u1_u0_u0_n132 ) , .B1( u1_u0_u0_n146 ) , .A1( u1_u0_u0_n147 ) , .B2( u1_u0_u0_n161 ) );
  AND2_X1 u1_u0_u0_U8 (.A1( u1_u0_u0_n114 ) , .A2( u1_u0_u0_n121 ) , .ZN( u1_u0_u0_n146 ) );
  NAND2_X1 u1_u0_u0_U80 (.ZN( u1_u0_u0_n110 ) , .A2( u1_u0_u0_n132 ) , .A1( u1_u0_u0_n145 ) );
  INV_X1 u1_u0_u0_U81 (.A( u1_u0_u0_n119 ) , .ZN( u1_u0_u0_n167 ) );
  NAND2_X1 u1_u0_u0_U82 (.A2( u1_u0_u0_n103 ) , .ZN( u1_u0_u0_n140 ) , .A1( u1_u0_u0_n94 ) );
  NAND2_X1 u1_u0_u0_U83 (.A1( u1_u0_u0_n101 ) , .ZN( u1_u0_u0_n130 ) , .A2( u1_u0_u0_n94 ) );
  NAND2_X1 u1_u0_u0_U84 (.ZN( u1_u0_u0_n108 ) , .A1( u1_u0_u0_n92 ) , .A2( u1_u0_u0_n94 ) );
  NAND2_X1 u1_u0_u0_U85 (.ZN( u1_u0_u0_n142 ) , .A1( u1_u0_u0_n94 ) , .A2( u1_u0_u0_n95 ) );
  NOR2_X1 u1_u0_u0_U86 (.A2( u1_u0_X_6 ) , .ZN( u1_u0_u0_n100 ) , .A1( u1_u0_u0_n162 ) );
  NOR2_X1 u1_u0_u0_U87 (.A2( u1_u0_X_3 ) , .A1( u1_u0_X_6 ) , .ZN( u1_u0_u0_n94 ) );
  NAND3_X1 u1_u0_u0_U88 (.ZN( u1_out0_23 ) , .A3( u1_u0_u0_n137 ) , .A1( u1_u0_u0_n168 ) , .A2( u1_u0_u0_n171 ) );
  NAND3_X1 u1_u0_u0_U89 (.A3( u1_u0_u0_n127 ) , .A2( u1_u0_u0_n128 ) , .ZN( u1_u0_u0_n135 ) , .A1( u1_u0_u0_n150 ) );
  AND2_X1 u1_u0_u0_U9 (.A1( u1_u0_u0_n131 ) , .ZN( u1_u0_u0_n141 ) , .A2( u1_u0_u0_n150 ) );
  NAND3_X1 u1_u0_u0_U90 (.ZN( u1_u0_u0_n117 ) , .A3( u1_u0_u0_n132 ) , .A2( u1_u0_u0_n139 ) , .A1( u1_u0_u0_n148 ) );
  NAND3_X1 u1_u0_u0_U91 (.ZN( u1_u0_u0_n109 ) , .A2( u1_u0_u0_n114 ) , .A3( u1_u0_u0_n140 ) , .A1( u1_u0_u0_n149 ) );
  NAND3_X1 u1_u0_u0_U92 (.ZN( u1_out0_9 ) , .A3( u1_u0_u0_n106 ) , .A2( u1_u0_u0_n171 ) , .A1( u1_u0_u0_n174 ) );
  NAND3_X1 u1_u0_u0_U93 (.A2( u1_u0_u0_n128 ) , .A1( u1_u0_u0_n132 ) , .A3( u1_u0_u0_n146 ) , .ZN( u1_u0_u0_n97 ) );
  OAI22_X1 u1_u0_u3_U10 (.B1( u1_u0_u3_n113 ) , .A2( u1_u0_u3_n135 ) , .A1( u1_u0_u3_n150 ) , .B2( u1_u0_u3_n164 ) , .ZN( u1_u0_u3_n98 ) );
  OAI211_X1 u1_u0_u3_U11 (.B( u1_u0_u3_n106 ) , .ZN( u1_u0_u3_n119 ) , .C2( u1_u0_u3_n128 ) , .C1( u1_u0_u3_n167 ) , .A( u1_u0_u3_n181 ) );
  AOI221_X1 u1_u0_u3_U12 (.C1( u1_u0_u3_n105 ) , .ZN( u1_u0_u3_n106 ) , .A( u1_u0_u3_n131 ) , .B2( u1_u0_u3_n132 ) , .C2( u1_u0_u3_n133 ) , .B1( u1_u0_u3_n169 ) );
  INV_X1 u1_u0_u3_U13 (.ZN( u1_u0_u3_n181 ) , .A( u1_u0_u3_n98 ) );
  NAND2_X1 u1_u0_u3_U14 (.ZN( u1_u0_u3_n105 ) , .A2( u1_u0_u3_n130 ) , .A1( u1_u0_u3_n155 ) );
  AOI22_X1 u1_u0_u3_U15 (.B1( u1_u0_u3_n115 ) , .A2( u1_u0_u3_n116 ) , .ZN( u1_u0_u3_n123 ) , .B2( u1_u0_u3_n133 ) , .A1( u1_u0_u3_n169 ) );
  NAND2_X1 u1_u0_u3_U16 (.ZN( u1_u0_u3_n116 ) , .A2( u1_u0_u3_n151 ) , .A1( u1_u0_u3_n182 ) );
  NOR2_X1 u1_u0_u3_U17 (.ZN( u1_u0_u3_n126 ) , .A2( u1_u0_u3_n150 ) , .A1( u1_u0_u3_n164 ) );
  AOI21_X1 u1_u0_u3_U18 (.ZN( u1_u0_u3_n112 ) , .B2( u1_u0_u3_n146 ) , .B1( u1_u0_u3_n155 ) , .A( u1_u0_u3_n167 ) );
  NAND2_X1 u1_u0_u3_U19 (.A1( u1_u0_u3_n135 ) , .ZN( u1_u0_u3_n142 ) , .A2( u1_u0_u3_n164 ) );
  NAND2_X1 u1_u0_u3_U20 (.ZN( u1_u0_u3_n132 ) , .A2( u1_u0_u3_n152 ) , .A1( u1_u0_u3_n156 ) );
  INV_X1 u1_u0_u3_U21 (.A( u1_u0_u3_n133 ) , .ZN( u1_u0_u3_n165 ) );
  AND2_X1 u1_u0_u3_U22 (.A2( u1_u0_u3_n113 ) , .A1( u1_u0_u3_n114 ) , .ZN( u1_u0_u3_n151 ) );
  INV_X1 u1_u0_u3_U23 (.A( u1_u0_u3_n135 ) , .ZN( u1_u0_u3_n170 ) );
  NAND2_X1 u1_u0_u3_U24 (.A1( u1_u0_u3_n107 ) , .A2( u1_u0_u3_n108 ) , .ZN( u1_u0_u3_n140 ) );
  NAND2_X1 u1_u0_u3_U25 (.ZN( u1_u0_u3_n117 ) , .A1( u1_u0_u3_n124 ) , .A2( u1_u0_u3_n148 ) );
  NAND2_X1 u1_u0_u3_U26 (.ZN( u1_u0_u3_n143 ) , .A1( u1_u0_u3_n165 ) , .A2( u1_u0_u3_n167 ) );
  INV_X1 u1_u0_u3_U27 (.A( u1_u0_u3_n130 ) , .ZN( u1_u0_u3_n177 ) );
  INV_X1 u1_u0_u3_U28 (.A( u1_u0_u3_n128 ) , .ZN( u1_u0_u3_n176 ) );
  INV_X1 u1_u0_u3_U29 (.A( u1_u0_u3_n155 ) , .ZN( u1_u0_u3_n174 ) );
  INV_X1 u1_u0_u3_U3 (.A( u1_u0_u3_n140 ) , .ZN( u1_u0_u3_n182 ) );
  INV_X1 u1_u0_u3_U30 (.A( u1_u0_u3_n139 ) , .ZN( u1_u0_u3_n185 ) );
  NOR2_X1 u1_u0_u3_U31 (.ZN( u1_u0_u3_n135 ) , .A2( u1_u0_u3_n141 ) , .A1( u1_u0_u3_n169 ) );
  OAI222_X1 u1_u0_u3_U32 (.C2( u1_u0_u3_n107 ) , .A2( u1_u0_u3_n108 ) , .B1( u1_u0_u3_n135 ) , .ZN( u1_u0_u3_n138 ) , .B2( u1_u0_u3_n146 ) , .C1( u1_u0_u3_n154 ) , .A1( u1_u0_u3_n164 ) );
  NOR4_X1 u1_u0_u3_U33 (.A4( u1_u0_u3_n157 ) , .A3( u1_u0_u3_n158 ) , .A2( u1_u0_u3_n159 ) , .A1( u1_u0_u3_n160 ) , .ZN( u1_u0_u3_n161 ) );
  AOI21_X1 u1_u0_u3_U34 (.B2( u1_u0_u3_n152 ) , .B1( u1_u0_u3_n153 ) , .ZN( u1_u0_u3_n158 ) , .A( u1_u0_u3_n164 ) );
  AOI21_X1 u1_u0_u3_U35 (.A( u1_u0_u3_n154 ) , .B2( u1_u0_u3_n155 ) , .B1( u1_u0_u3_n156 ) , .ZN( u1_u0_u3_n157 ) );
  AOI21_X1 u1_u0_u3_U36 (.A( u1_u0_u3_n149 ) , .B2( u1_u0_u3_n150 ) , .B1( u1_u0_u3_n151 ) , .ZN( u1_u0_u3_n159 ) );
  OAI211_X1 u1_u0_u3_U37 (.B( u1_u0_u3_n127 ) , .ZN( u1_u0_u3_n139 ) , .C1( u1_u0_u3_n150 ) , .C2( u1_u0_u3_n154 ) , .A( u1_u0_u3_n184 ) );
  INV_X1 u1_u0_u3_U38 (.A( u1_u0_u3_n125 ) , .ZN( u1_u0_u3_n184 ) );
  AOI221_X1 u1_u0_u3_U39 (.A( u1_u0_u3_n126 ) , .ZN( u1_u0_u3_n127 ) , .C2( u1_u0_u3_n132 ) , .C1( u1_u0_u3_n169 ) , .B2( u1_u0_u3_n170 ) , .B1( u1_u0_u3_n174 ) );
  INV_X1 u1_u0_u3_U4 (.A( u1_u0_u3_n129 ) , .ZN( u1_u0_u3_n183 ) );
  OAI22_X1 u1_u0_u3_U40 (.A1( u1_u0_u3_n124 ) , .ZN( u1_u0_u3_n125 ) , .B2( u1_u0_u3_n145 ) , .A2( u1_u0_u3_n165 ) , .B1( u1_u0_u3_n167 ) );
  AOI211_X1 u1_u0_u3_U41 (.ZN( u1_u0_u3_n109 ) , .A( u1_u0_u3_n119 ) , .C2( u1_u0_u3_n129 ) , .B( u1_u0_u3_n138 ) , .C1( u1_u0_u3_n141 ) );
  AOI211_X1 u1_u0_u3_U42 (.B( u1_u0_u3_n119 ) , .A( u1_u0_u3_n120 ) , .C2( u1_u0_u3_n121 ) , .ZN( u1_u0_u3_n122 ) , .C1( u1_u0_u3_n179 ) );
  INV_X1 u1_u0_u3_U43 (.A( u1_u0_u3_n156 ) , .ZN( u1_u0_u3_n179 ) );
  OAI22_X1 u1_u0_u3_U44 (.B1( u1_u0_u3_n118 ) , .ZN( u1_u0_u3_n120 ) , .A1( u1_u0_u3_n135 ) , .B2( u1_u0_u3_n154 ) , .A2( u1_u0_u3_n178 ) );
  AND3_X1 u1_u0_u3_U45 (.ZN( u1_u0_u3_n118 ) , .A2( u1_u0_u3_n124 ) , .A1( u1_u0_u3_n144 ) , .A3( u1_u0_u3_n152 ) );
  INV_X1 u1_u0_u3_U46 (.A( u1_u0_u3_n121 ) , .ZN( u1_u0_u3_n164 ) );
  NAND2_X1 u1_u0_u3_U47 (.ZN( u1_u0_u3_n133 ) , .A1( u1_u0_u3_n154 ) , .A2( u1_u0_u3_n164 ) );
  NOR2_X1 u1_u0_u3_U48 (.A1( u1_u0_u3_n113 ) , .ZN( u1_u0_u3_n131 ) , .A2( u1_u0_u3_n154 ) );
  NAND2_X1 u1_u0_u3_U49 (.A1( u1_u0_u3_n103 ) , .ZN( u1_u0_u3_n150 ) , .A2( u1_u0_u3_n99 ) );
  INV_X1 u1_u0_u3_U5 (.A( u1_u0_u3_n117 ) , .ZN( u1_u0_u3_n178 ) );
  NAND2_X1 u1_u0_u3_U50 (.A2( u1_u0_u3_n102 ) , .ZN( u1_u0_u3_n155 ) , .A1( u1_u0_u3_n97 ) );
  INV_X1 u1_u0_u3_U51 (.A( u1_u0_u3_n141 ) , .ZN( u1_u0_u3_n167 ) );
  AOI21_X1 u1_u0_u3_U52 (.B2( u1_u0_u3_n114 ) , .B1( u1_u0_u3_n146 ) , .A( u1_u0_u3_n154 ) , .ZN( u1_u0_u3_n94 ) );
  AOI21_X1 u1_u0_u3_U53 (.ZN( u1_u0_u3_n110 ) , .B2( u1_u0_u3_n142 ) , .B1( u1_u0_u3_n186 ) , .A( u1_u0_u3_n95 ) );
  INV_X1 u1_u0_u3_U54 (.A( u1_u0_u3_n145 ) , .ZN( u1_u0_u3_n186 ) );
  AOI21_X1 u1_u0_u3_U55 (.B1( u1_u0_u3_n124 ) , .A( u1_u0_u3_n149 ) , .B2( u1_u0_u3_n155 ) , .ZN( u1_u0_u3_n95 ) );
  INV_X1 u1_u0_u3_U56 (.A( u1_u0_u3_n149 ) , .ZN( u1_u0_u3_n169 ) );
  NAND2_X1 u1_u0_u3_U57 (.ZN( u1_u0_u3_n124 ) , .A1( u1_u0_u3_n96 ) , .A2( u1_u0_u3_n97 ) );
  NAND2_X1 u1_u0_u3_U58 (.A2( u1_u0_u3_n100 ) , .ZN( u1_u0_u3_n146 ) , .A1( u1_u0_u3_n96 ) );
  NAND2_X1 u1_u0_u3_U59 (.A1( u1_u0_u3_n101 ) , .ZN( u1_u0_u3_n145 ) , .A2( u1_u0_u3_n99 ) );
  AOI221_X1 u1_u0_u3_U6 (.A( u1_u0_u3_n131 ) , .C2( u1_u0_u3_n132 ) , .C1( u1_u0_u3_n133 ) , .ZN( u1_u0_u3_n134 ) , .B1( u1_u0_u3_n143 ) , .B2( u1_u0_u3_n177 ) );
  NAND2_X1 u1_u0_u3_U60 (.A1( u1_u0_u3_n100 ) , .ZN( u1_u0_u3_n156 ) , .A2( u1_u0_u3_n99 ) );
  NAND2_X1 u1_u0_u3_U61 (.A2( u1_u0_u3_n101 ) , .A1( u1_u0_u3_n104 ) , .ZN( u1_u0_u3_n148 ) );
  NAND2_X1 u1_u0_u3_U62 (.A1( u1_u0_u3_n100 ) , .A2( u1_u0_u3_n102 ) , .ZN( u1_u0_u3_n128 ) );
  NAND2_X1 u1_u0_u3_U63 (.A2( u1_u0_u3_n101 ) , .A1( u1_u0_u3_n102 ) , .ZN( u1_u0_u3_n152 ) );
  NAND2_X1 u1_u0_u3_U64 (.A2( u1_u0_u3_n101 ) , .ZN( u1_u0_u3_n114 ) , .A1( u1_u0_u3_n96 ) );
  NAND2_X1 u1_u0_u3_U65 (.ZN( u1_u0_u3_n107 ) , .A1( u1_u0_u3_n97 ) , .A2( u1_u0_u3_n99 ) );
  NAND2_X1 u1_u0_u3_U66 (.A2( u1_u0_u3_n100 ) , .A1( u1_u0_u3_n104 ) , .ZN( u1_u0_u3_n113 ) );
  NAND2_X1 u1_u0_u3_U67 (.A1( u1_u0_u3_n104 ) , .ZN( u1_u0_u3_n153 ) , .A2( u1_u0_u3_n97 ) );
  NAND2_X1 u1_u0_u3_U68 (.A2( u1_u0_u3_n103 ) , .A1( u1_u0_u3_n104 ) , .ZN( u1_u0_u3_n130 ) );
  NAND2_X1 u1_u0_u3_U69 (.A2( u1_u0_u3_n103 ) , .ZN( u1_u0_u3_n144 ) , .A1( u1_u0_u3_n96 ) );
  OAI22_X1 u1_u0_u3_U7 (.B2( u1_u0_u3_n147 ) , .A2( u1_u0_u3_n148 ) , .ZN( u1_u0_u3_n160 ) , .B1( u1_u0_u3_n165 ) , .A1( u1_u0_u3_n168 ) );
  NAND2_X1 u1_u0_u3_U70 (.A1( u1_u0_u3_n102 ) , .A2( u1_u0_u3_n103 ) , .ZN( u1_u0_u3_n108 ) );
  NOR2_X1 u1_u0_u3_U71 (.A2( u1_u0_X_19 ) , .A1( u1_u0_X_20 ) , .ZN( u1_u0_u3_n99 ) );
  NOR2_X1 u1_u0_u3_U72 (.A2( u1_u0_X_21 ) , .A1( u1_u0_X_24 ) , .ZN( u1_u0_u3_n103 ) );
  NOR2_X1 u1_u0_u3_U73 (.A2( u1_u0_X_24 ) , .A1( u1_u0_u3_n171 ) , .ZN( u1_u0_u3_n97 ) );
  NOR2_X1 u1_u0_u3_U74 (.A2( u1_u0_X_23 ) , .ZN( u1_u0_u3_n141 ) , .A1( u1_u0_u3_n166 ) );
  NOR2_X1 u1_u0_u3_U75 (.A2( u1_u0_X_19 ) , .A1( u1_u0_u3_n172 ) , .ZN( u1_u0_u3_n96 ) );
  NAND2_X1 u1_u0_u3_U76 (.A1( u1_u0_X_22 ) , .A2( u1_u0_X_23 ) , .ZN( u1_u0_u3_n154 ) );
  NAND2_X1 u1_u0_u3_U77 (.A1( u1_u0_X_23 ) , .ZN( u1_u0_u3_n149 ) , .A2( u1_u0_u3_n166 ) );
  NOR2_X1 u1_u0_u3_U78 (.A2( u1_u0_X_22 ) , .A1( u1_u0_X_23 ) , .ZN( u1_u0_u3_n121 ) );
  AND2_X1 u1_u0_u3_U79 (.A1( u1_u0_X_24 ) , .ZN( u1_u0_u3_n101 ) , .A2( u1_u0_u3_n171 ) );
  AND3_X1 u1_u0_u3_U8 (.A3( u1_u0_u3_n144 ) , .A2( u1_u0_u3_n145 ) , .A1( u1_u0_u3_n146 ) , .ZN( u1_u0_u3_n147 ) );
  AND2_X1 u1_u0_u3_U80 (.A1( u1_u0_X_19 ) , .ZN( u1_u0_u3_n102 ) , .A2( u1_u0_u3_n172 ) );
  AND2_X1 u1_u0_u3_U81 (.A1( u1_u0_X_21 ) , .A2( u1_u0_X_24 ) , .ZN( u1_u0_u3_n100 ) );
  AND2_X1 u1_u0_u3_U82 (.A2( u1_u0_X_19 ) , .A1( u1_u0_X_20 ) , .ZN( u1_u0_u3_n104 ) );
  INV_X1 u1_u0_u3_U83 (.A( u1_u0_X_22 ) , .ZN( u1_u0_u3_n166 ) );
  INV_X1 u1_u0_u3_U84 (.A( u1_u0_X_21 ) , .ZN( u1_u0_u3_n171 ) );
  INV_X1 u1_u0_u3_U85 (.A( u1_u0_X_20 ) , .ZN( u1_u0_u3_n172 ) );
  NAND4_X1 u1_u0_u3_U86 (.ZN( u1_out0_26 ) , .A4( u1_u0_u3_n109 ) , .A3( u1_u0_u3_n110 ) , .A2( u1_u0_u3_n111 ) , .A1( u1_u0_u3_n173 ) );
  INV_X1 u1_u0_u3_U87 (.ZN( u1_u0_u3_n173 ) , .A( u1_u0_u3_n94 ) );
  OAI21_X1 u1_u0_u3_U88 (.ZN( u1_u0_u3_n111 ) , .B2( u1_u0_u3_n117 ) , .A( u1_u0_u3_n133 ) , .B1( u1_u0_u3_n176 ) );
  NAND4_X1 u1_u0_u3_U89 (.ZN( u1_out0_20 ) , .A4( u1_u0_u3_n122 ) , .A3( u1_u0_u3_n123 ) , .A1( u1_u0_u3_n175 ) , .A2( u1_u0_u3_n180 ) );
  INV_X1 u1_u0_u3_U9 (.A( u1_u0_u3_n143 ) , .ZN( u1_u0_u3_n168 ) );
  INV_X1 u1_u0_u3_U90 (.A( u1_u0_u3_n126 ) , .ZN( u1_u0_u3_n180 ) );
  INV_X1 u1_u0_u3_U91 (.A( u1_u0_u3_n112 ) , .ZN( u1_u0_u3_n175 ) );
  NAND4_X1 u1_u0_u3_U92 (.ZN( u1_out0_1 ) , .A4( u1_u0_u3_n161 ) , .A3( u1_u0_u3_n162 ) , .A2( u1_u0_u3_n163 ) , .A1( u1_u0_u3_n185 ) );
  NAND2_X1 u1_u0_u3_U93 (.ZN( u1_u0_u3_n163 ) , .A2( u1_u0_u3_n170 ) , .A1( u1_u0_u3_n176 ) );
  AOI22_X1 u1_u0_u3_U94 (.B2( u1_u0_u3_n140 ) , .B1( u1_u0_u3_n141 ) , .A2( u1_u0_u3_n142 ) , .ZN( u1_u0_u3_n162 ) , .A1( u1_u0_u3_n177 ) );
  OR4_X1 u1_u0_u3_U95 (.ZN( u1_out0_10 ) , .A4( u1_u0_u3_n136 ) , .A3( u1_u0_u3_n137 ) , .A1( u1_u0_u3_n138 ) , .A2( u1_u0_u3_n139 ) );
  OAI222_X1 u1_u0_u3_U96 (.C1( u1_u0_u3_n128 ) , .ZN( u1_u0_u3_n137 ) , .B1( u1_u0_u3_n148 ) , .A2( u1_u0_u3_n150 ) , .B2( u1_u0_u3_n154 ) , .C2( u1_u0_u3_n164 ) , .A1( u1_u0_u3_n167 ) );
  OAI221_X1 u1_u0_u3_U97 (.A( u1_u0_u3_n134 ) , .B2( u1_u0_u3_n135 ) , .ZN( u1_u0_u3_n136 ) , .C1( u1_u0_u3_n149 ) , .B1( u1_u0_u3_n151 ) , .C2( u1_u0_u3_n183 ) );
  NAND3_X1 u1_u0_u3_U98 (.A1( u1_u0_u3_n114 ) , .ZN( u1_u0_u3_n115 ) , .A2( u1_u0_u3_n145 ) , .A3( u1_u0_u3_n153 ) );
  NAND3_X1 u1_u0_u3_U99 (.ZN( u1_u0_u3_n129 ) , .A2( u1_u0_u3_n144 ) , .A1( u1_u0_u3_n153 ) , .A3( u1_u0_u3_n182 ) );
  XOR2_X1 u1_u10_U1 (.B( u1_K11_9 ) , .A( u1_R9_6 ) , .Z( u1_u10_X_9 ) );
  XOR2_X1 u1_u10_U2 (.B( u1_K11_8 ) , .A( u1_R9_5 ) , .Z( u1_u10_X_8 ) );
  XOR2_X1 u1_u10_U42 (.B( u1_K11_16 ) , .A( u1_R9_11 ) , .Z( u1_u10_X_16 ) );
  XOR2_X1 u1_u10_U43 (.B( u1_K11_15 ) , .A( u1_R9_10 ) , .Z( u1_u10_X_15 ) );
  XOR2_X1 u1_u10_U44 (.B( u1_K11_14 ) , .A( u1_R9_9 ) , .Z( u1_u10_X_14 ) );
  XOR2_X1 u1_u10_U45 (.B( u1_K11_13 ) , .A( u1_R9_8 ) , .Z( u1_u10_X_13 ) );
  XOR2_X1 u1_u10_U46 (.B( u1_K11_12 ) , .A( u1_R9_9 ) , .Z( u1_u10_X_12 ) );
  XOR2_X1 u1_u10_U47 (.B( u1_K11_11 ) , .A( u1_R9_8 ) , .Z( u1_u10_X_11 ) );
  XOR2_X1 u1_u10_U48 (.B( u1_K11_10 ) , .A( u1_R9_7 ) , .Z( u1_u10_X_10 ) );
  AOI21_X1 u1_u10_u1_U10 (.B2( u1_u10_u1_n155 ) , .B1( u1_u10_u1_n156 ) , .ZN( u1_u10_u1_n157 ) , .A( u1_u10_u1_n174 ) );
  NAND3_X1 u1_u10_u1_U100 (.ZN( u1_u10_u1_n113 ) , .A1( u1_u10_u1_n120 ) , .A3( u1_u10_u1_n133 ) , .A2( u1_u10_u1_n155 ) );
  NAND2_X1 u1_u10_u1_U11 (.ZN( u1_u10_u1_n140 ) , .A2( u1_u10_u1_n150 ) , .A1( u1_u10_u1_n155 ) );
  NAND2_X1 u1_u10_u1_U12 (.A1( u1_u10_u1_n131 ) , .ZN( u1_u10_u1_n147 ) , .A2( u1_u10_u1_n153 ) );
  AOI22_X1 u1_u10_u1_U13 (.B2( u1_u10_u1_n136 ) , .A2( u1_u10_u1_n137 ) , .ZN( u1_u10_u1_n143 ) , .A1( u1_u10_u1_n171 ) , .B1( u1_u10_u1_n173 ) );
  INV_X1 u1_u10_u1_U14 (.A( u1_u10_u1_n147 ) , .ZN( u1_u10_u1_n181 ) );
  INV_X1 u1_u10_u1_U15 (.A( u1_u10_u1_n139 ) , .ZN( u1_u10_u1_n174 ) );
  OR4_X1 u1_u10_u1_U16 (.A4( u1_u10_u1_n106 ) , .A3( u1_u10_u1_n107 ) , .ZN( u1_u10_u1_n108 ) , .A1( u1_u10_u1_n117 ) , .A2( u1_u10_u1_n184 ) );
  AOI21_X1 u1_u10_u1_U17 (.ZN( u1_u10_u1_n106 ) , .A( u1_u10_u1_n112 ) , .B1( u1_u10_u1_n154 ) , .B2( u1_u10_u1_n156 ) );
  AOI21_X1 u1_u10_u1_U18 (.ZN( u1_u10_u1_n107 ) , .B1( u1_u10_u1_n134 ) , .B2( u1_u10_u1_n149 ) , .A( u1_u10_u1_n174 ) );
  INV_X1 u1_u10_u1_U19 (.A( u1_u10_u1_n101 ) , .ZN( u1_u10_u1_n184 ) );
  INV_X1 u1_u10_u1_U20 (.A( u1_u10_u1_n112 ) , .ZN( u1_u10_u1_n171 ) );
  NAND2_X1 u1_u10_u1_U21 (.ZN( u1_u10_u1_n141 ) , .A1( u1_u10_u1_n153 ) , .A2( u1_u10_u1_n156 ) );
  AND2_X1 u1_u10_u1_U22 (.A1( u1_u10_u1_n123 ) , .ZN( u1_u10_u1_n134 ) , .A2( u1_u10_u1_n161 ) );
  NAND2_X1 u1_u10_u1_U23 (.A2( u1_u10_u1_n115 ) , .A1( u1_u10_u1_n116 ) , .ZN( u1_u10_u1_n148 ) );
  NAND2_X1 u1_u10_u1_U24 (.A2( u1_u10_u1_n133 ) , .A1( u1_u10_u1_n135 ) , .ZN( u1_u10_u1_n159 ) );
  NAND2_X1 u1_u10_u1_U25 (.A2( u1_u10_u1_n115 ) , .A1( u1_u10_u1_n120 ) , .ZN( u1_u10_u1_n132 ) );
  INV_X1 u1_u10_u1_U26 (.A( u1_u10_u1_n154 ) , .ZN( u1_u10_u1_n178 ) );
  INV_X1 u1_u10_u1_U27 (.A( u1_u10_u1_n151 ) , .ZN( u1_u10_u1_n183 ) );
  AND2_X1 u1_u10_u1_U28 (.A1( u1_u10_u1_n129 ) , .A2( u1_u10_u1_n133 ) , .ZN( u1_u10_u1_n149 ) );
  INV_X1 u1_u10_u1_U29 (.A( u1_u10_u1_n131 ) , .ZN( u1_u10_u1_n180 ) );
  INV_X1 u1_u10_u1_U3 (.A( u1_u10_u1_n159 ) , .ZN( u1_u10_u1_n182 ) );
  OAI221_X1 u1_u10_u1_U30 (.A( u1_u10_u1_n119 ) , .C2( u1_u10_u1_n129 ) , .ZN( u1_u10_u1_n138 ) , .B2( u1_u10_u1_n152 ) , .C1( u1_u10_u1_n174 ) , .B1( u1_u10_u1_n187 ) );
  INV_X1 u1_u10_u1_U31 (.A( u1_u10_u1_n148 ) , .ZN( u1_u10_u1_n187 ) );
  AOI211_X1 u1_u10_u1_U32 (.B( u1_u10_u1_n117 ) , .A( u1_u10_u1_n118 ) , .ZN( u1_u10_u1_n119 ) , .C2( u1_u10_u1_n146 ) , .C1( u1_u10_u1_n159 ) );
  NOR2_X1 u1_u10_u1_U33 (.A1( u1_u10_u1_n168 ) , .A2( u1_u10_u1_n176 ) , .ZN( u1_u10_u1_n98 ) );
  AOI211_X1 u1_u10_u1_U34 (.B( u1_u10_u1_n162 ) , .A( u1_u10_u1_n163 ) , .C2( u1_u10_u1_n164 ) , .ZN( u1_u10_u1_n165 ) , .C1( u1_u10_u1_n171 ) );
  AOI21_X1 u1_u10_u1_U35 (.A( u1_u10_u1_n160 ) , .B2( u1_u10_u1_n161 ) , .ZN( u1_u10_u1_n162 ) , .B1( u1_u10_u1_n182 ) );
  OR2_X1 u1_u10_u1_U36 (.A2( u1_u10_u1_n157 ) , .A1( u1_u10_u1_n158 ) , .ZN( u1_u10_u1_n163 ) );
  OAI21_X1 u1_u10_u1_U37 (.B2( u1_u10_u1_n123 ) , .ZN( u1_u10_u1_n145 ) , .B1( u1_u10_u1_n160 ) , .A( u1_u10_u1_n185 ) );
  INV_X1 u1_u10_u1_U38 (.A( u1_u10_u1_n122 ) , .ZN( u1_u10_u1_n185 ) );
  AOI21_X1 u1_u10_u1_U39 (.B2( u1_u10_u1_n120 ) , .B1( u1_u10_u1_n121 ) , .ZN( u1_u10_u1_n122 ) , .A( u1_u10_u1_n128 ) );
  AOI221_X1 u1_u10_u1_U4 (.A( u1_u10_u1_n138 ) , .C2( u1_u10_u1_n139 ) , .C1( u1_u10_u1_n140 ) , .B2( u1_u10_u1_n141 ) , .ZN( u1_u10_u1_n142 ) , .B1( u1_u10_u1_n175 ) );
  NAND2_X1 u1_u10_u1_U40 (.A1( u1_u10_u1_n128 ) , .ZN( u1_u10_u1_n146 ) , .A2( u1_u10_u1_n160 ) );
  NAND2_X1 u1_u10_u1_U41 (.A2( u1_u10_u1_n112 ) , .ZN( u1_u10_u1_n139 ) , .A1( u1_u10_u1_n152 ) );
  NAND2_X1 u1_u10_u1_U42 (.A1( u1_u10_u1_n105 ) , .ZN( u1_u10_u1_n156 ) , .A2( u1_u10_u1_n99 ) );
  AOI221_X1 u1_u10_u1_U43 (.B1( u1_u10_u1_n140 ) , .ZN( u1_u10_u1_n167 ) , .B2( u1_u10_u1_n172 ) , .C2( u1_u10_u1_n175 ) , .C1( u1_u10_u1_n178 ) , .A( u1_u10_u1_n188 ) );
  INV_X1 u1_u10_u1_U44 (.ZN( u1_u10_u1_n188 ) , .A( u1_u10_u1_n97 ) );
  AOI211_X1 u1_u10_u1_U45 (.A( u1_u10_u1_n118 ) , .C1( u1_u10_u1_n132 ) , .C2( u1_u10_u1_n139 ) , .B( u1_u10_u1_n96 ) , .ZN( u1_u10_u1_n97 ) );
  AOI21_X1 u1_u10_u1_U46 (.B2( u1_u10_u1_n121 ) , .B1( u1_u10_u1_n135 ) , .A( u1_u10_u1_n152 ) , .ZN( u1_u10_u1_n96 ) );
  NOR2_X1 u1_u10_u1_U47 (.ZN( u1_u10_u1_n117 ) , .A1( u1_u10_u1_n121 ) , .A2( u1_u10_u1_n160 ) );
  AOI21_X1 u1_u10_u1_U48 (.A( u1_u10_u1_n128 ) , .B2( u1_u10_u1_n129 ) , .ZN( u1_u10_u1_n130 ) , .B1( u1_u10_u1_n150 ) );
  NAND2_X1 u1_u10_u1_U49 (.ZN( u1_u10_u1_n112 ) , .A1( u1_u10_u1_n169 ) , .A2( u1_u10_u1_n170 ) );
  AOI211_X1 u1_u10_u1_U5 (.ZN( u1_u10_u1_n124 ) , .A( u1_u10_u1_n138 ) , .C2( u1_u10_u1_n139 ) , .B( u1_u10_u1_n145 ) , .C1( u1_u10_u1_n147 ) );
  NAND2_X1 u1_u10_u1_U50 (.ZN( u1_u10_u1_n129 ) , .A2( u1_u10_u1_n95 ) , .A1( u1_u10_u1_n98 ) );
  NAND2_X1 u1_u10_u1_U51 (.A1( u1_u10_u1_n102 ) , .ZN( u1_u10_u1_n154 ) , .A2( u1_u10_u1_n99 ) );
  NAND2_X1 u1_u10_u1_U52 (.A2( u1_u10_u1_n100 ) , .ZN( u1_u10_u1_n135 ) , .A1( u1_u10_u1_n99 ) );
  AOI21_X1 u1_u10_u1_U53 (.A( u1_u10_u1_n152 ) , .B2( u1_u10_u1_n153 ) , .B1( u1_u10_u1_n154 ) , .ZN( u1_u10_u1_n158 ) );
  INV_X1 u1_u10_u1_U54 (.A( u1_u10_u1_n160 ) , .ZN( u1_u10_u1_n175 ) );
  NAND2_X1 u1_u10_u1_U55 (.A1( u1_u10_u1_n100 ) , .ZN( u1_u10_u1_n116 ) , .A2( u1_u10_u1_n95 ) );
  NAND2_X1 u1_u10_u1_U56 (.A1( u1_u10_u1_n102 ) , .ZN( u1_u10_u1_n131 ) , .A2( u1_u10_u1_n95 ) );
  NAND2_X1 u1_u10_u1_U57 (.A2( u1_u10_u1_n104 ) , .ZN( u1_u10_u1_n121 ) , .A1( u1_u10_u1_n98 ) );
  NAND2_X1 u1_u10_u1_U58 (.A1( u1_u10_u1_n103 ) , .ZN( u1_u10_u1_n153 ) , .A2( u1_u10_u1_n98 ) );
  NAND2_X1 u1_u10_u1_U59 (.A2( u1_u10_u1_n104 ) , .A1( u1_u10_u1_n105 ) , .ZN( u1_u10_u1_n133 ) );
  AOI22_X1 u1_u10_u1_U6 (.B2( u1_u10_u1_n113 ) , .A2( u1_u10_u1_n114 ) , .ZN( u1_u10_u1_n125 ) , .A1( u1_u10_u1_n171 ) , .B1( u1_u10_u1_n173 ) );
  NAND2_X1 u1_u10_u1_U60 (.ZN( u1_u10_u1_n150 ) , .A2( u1_u10_u1_n98 ) , .A1( u1_u10_u1_n99 ) );
  NAND2_X1 u1_u10_u1_U61 (.A1( u1_u10_u1_n105 ) , .ZN( u1_u10_u1_n155 ) , .A2( u1_u10_u1_n95 ) );
  OAI21_X1 u1_u10_u1_U62 (.ZN( u1_u10_u1_n109 ) , .B1( u1_u10_u1_n129 ) , .B2( u1_u10_u1_n160 ) , .A( u1_u10_u1_n167 ) );
  NAND2_X1 u1_u10_u1_U63 (.A2( u1_u10_u1_n100 ) , .A1( u1_u10_u1_n103 ) , .ZN( u1_u10_u1_n120 ) );
  NAND2_X1 u1_u10_u1_U64 (.A1( u1_u10_u1_n102 ) , .A2( u1_u10_u1_n104 ) , .ZN( u1_u10_u1_n115 ) );
  NAND2_X1 u1_u10_u1_U65 (.A2( u1_u10_u1_n100 ) , .A1( u1_u10_u1_n104 ) , .ZN( u1_u10_u1_n151 ) );
  NAND2_X1 u1_u10_u1_U66 (.A2( u1_u10_u1_n103 ) , .A1( u1_u10_u1_n105 ) , .ZN( u1_u10_u1_n161 ) );
  INV_X1 u1_u10_u1_U67 (.A( u1_u10_u1_n152 ) , .ZN( u1_u10_u1_n173 ) );
  INV_X1 u1_u10_u1_U68 (.A( u1_u10_u1_n128 ) , .ZN( u1_u10_u1_n172 ) );
  NAND2_X1 u1_u10_u1_U69 (.A2( u1_u10_u1_n102 ) , .A1( u1_u10_u1_n103 ) , .ZN( u1_u10_u1_n123 ) );
  NAND2_X1 u1_u10_u1_U7 (.ZN( u1_u10_u1_n114 ) , .A1( u1_u10_u1_n134 ) , .A2( u1_u10_u1_n156 ) );
  NOR2_X1 u1_u10_u1_U70 (.A2( u1_u10_X_7 ) , .A1( u1_u10_X_8 ) , .ZN( u1_u10_u1_n95 ) );
  NOR2_X1 u1_u10_u1_U71 (.A1( u1_u10_X_12 ) , .A2( u1_u10_X_9 ) , .ZN( u1_u10_u1_n100 ) );
  NOR2_X1 u1_u10_u1_U72 (.A2( u1_u10_X_8 ) , .A1( u1_u10_u1_n177 ) , .ZN( u1_u10_u1_n99 ) );
  NOR2_X1 u1_u10_u1_U73 (.A2( u1_u10_X_12 ) , .ZN( u1_u10_u1_n102 ) , .A1( u1_u10_u1_n176 ) );
  NOR2_X1 u1_u10_u1_U74 (.A2( u1_u10_X_9 ) , .ZN( u1_u10_u1_n105 ) , .A1( u1_u10_u1_n168 ) );
  NAND2_X1 u1_u10_u1_U75 (.A1( u1_u10_X_10 ) , .ZN( u1_u10_u1_n160 ) , .A2( u1_u10_u1_n169 ) );
  NAND2_X1 u1_u10_u1_U76 (.A2( u1_u10_X_10 ) , .A1( u1_u10_X_11 ) , .ZN( u1_u10_u1_n152 ) );
  NAND2_X1 u1_u10_u1_U77 (.A1( u1_u10_X_11 ) , .ZN( u1_u10_u1_n128 ) , .A2( u1_u10_u1_n170 ) );
  AND2_X1 u1_u10_u1_U78 (.A2( u1_u10_X_7 ) , .A1( u1_u10_X_8 ) , .ZN( u1_u10_u1_n104 ) );
  AND2_X1 u1_u10_u1_U79 (.A1( u1_u10_X_8 ) , .ZN( u1_u10_u1_n103 ) , .A2( u1_u10_u1_n177 ) );
  NOR2_X1 u1_u10_u1_U8 (.A1( u1_u10_u1_n112 ) , .A2( u1_u10_u1_n116 ) , .ZN( u1_u10_u1_n118 ) );
  INV_X1 u1_u10_u1_U80 (.A( u1_u10_X_10 ) , .ZN( u1_u10_u1_n170 ) );
  INV_X1 u1_u10_u1_U81 (.A( u1_u10_X_9 ) , .ZN( u1_u10_u1_n176 ) );
  INV_X1 u1_u10_u1_U82 (.A( u1_u10_X_11 ) , .ZN( u1_u10_u1_n169 ) );
  INV_X1 u1_u10_u1_U83 (.A( u1_u10_X_12 ) , .ZN( u1_u10_u1_n168 ) );
  INV_X1 u1_u10_u1_U84 (.A( u1_u10_X_7 ) , .ZN( u1_u10_u1_n177 ) );
  NAND4_X1 u1_u10_u1_U85 (.ZN( u1_out10_18 ) , .A4( u1_u10_u1_n165 ) , .A3( u1_u10_u1_n166 ) , .A1( u1_u10_u1_n167 ) , .A2( u1_u10_u1_n186 ) );
  AOI22_X1 u1_u10_u1_U86 (.B2( u1_u10_u1_n146 ) , .B1( u1_u10_u1_n147 ) , .A2( u1_u10_u1_n148 ) , .ZN( u1_u10_u1_n166 ) , .A1( u1_u10_u1_n172 ) );
  INV_X1 u1_u10_u1_U87 (.A( u1_u10_u1_n145 ) , .ZN( u1_u10_u1_n186 ) );
  NAND4_X1 u1_u10_u1_U88 (.ZN( u1_out10_2 ) , .A4( u1_u10_u1_n142 ) , .A3( u1_u10_u1_n143 ) , .A2( u1_u10_u1_n144 ) , .A1( u1_u10_u1_n179 ) );
  OAI21_X1 u1_u10_u1_U89 (.B2( u1_u10_u1_n132 ) , .ZN( u1_u10_u1_n144 ) , .A( u1_u10_u1_n146 ) , .B1( u1_u10_u1_n180 ) );
  OAI21_X1 u1_u10_u1_U9 (.ZN( u1_u10_u1_n101 ) , .B1( u1_u10_u1_n141 ) , .A( u1_u10_u1_n146 ) , .B2( u1_u10_u1_n183 ) );
  INV_X1 u1_u10_u1_U90 (.A( u1_u10_u1_n130 ) , .ZN( u1_u10_u1_n179 ) );
  OR4_X1 u1_u10_u1_U91 (.ZN( u1_out10_13 ) , .A4( u1_u10_u1_n108 ) , .A3( u1_u10_u1_n109 ) , .A2( u1_u10_u1_n110 ) , .A1( u1_u10_u1_n111 ) );
  AOI21_X1 u1_u10_u1_U92 (.ZN( u1_u10_u1_n111 ) , .A( u1_u10_u1_n128 ) , .B2( u1_u10_u1_n131 ) , .B1( u1_u10_u1_n135 ) );
  AOI21_X1 u1_u10_u1_U93 (.ZN( u1_u10_u1_n110 ) , .A( u1_u10_u1_n116 ) , .B1( u1_u10_u1_n152 ) , .B2( u1_u10_u1_n160 ) );
  NAND4_X1 u1_u10_u1_U94 (.ZN( u1_out10_28 ) , .A4( u1_u10_u1_n124 ) , .A3( u1_u10_u1_n125 ) , .A2( u1_u10_u1_n126 ) , .A1( u1_u10_u1_n127 ) );
  OAI21_X1 u1_u10_u1_U95 (.ZN( u1_u10_u1_n127 ) , .B2( u1_u10_u1_n139 ) , .B1( u1_u10_u1_n175 ) , .A( u1_u10_u1_n183 ) );
  OAI21_X1 u1_u10_u1_U96 (.ZN( u1_u10_u1_n126 ) , .B2( u1_u10_u1_n140 ) , .A( u1_u10_u1_n146 ) , .B1( u1_u10_u1_n178 ) );
  NAND3_X1 u1_u10_u1_U97 (.A3( u1_u10_u1_n149 ) , .A2( u1_u10_u1_n150 ) , .A1( u1_u10_u1_n151 ) , .ZN( u1_u10_u1_n164 ) );
  NAND3_X1 u1_u10_u1_U98 (.A3( u1_u10_u1_n134 ) , .A2( u1_u10_u1_n135 ) , .ZN( u1_u10_u1_n136 ) , .A1( u1_u10_u1_n151 ) );
  NAND3_X1 u1_u10_u1_U99 (.A1( u1_u10_u1_n133 ) , .ZN( u1_u10_u1_n137 ) , .A2( u1_u10_u1_n154 ) , .A3( u1_u10_u1_n181 ) );
  OAI22_X1 u1_u10_u2_U10 (.ZN( u1_u10_u2_n109 ) , .A2( u1_u10_u2_n113 ) , .B2( u1_u10_u2_n133 ) , .B1( u1_u10_u2_n167 ) , .A1( u1_u10_u2_n168 ) );
  NAND3_X1 u1_u10_u2_U100 (.A2( u1_u10_u2_n100 ) , .A1( u1_u10_u2_n104 ) , .A3( u1_u10_u2_n138 ) , .ZN( u1_u10_u2_n98 ) );
  OAI22_X1 u1_u10_u2_U11 (.B1( u1_u10_u2_n151 ) , .A2( u1_u10_u2_n152 ) , .A1( u1_u10_u2_n153 ) , .ZN( u1_u10_u2_n160 ) , .B2( u1_u10_u2_n168 ) );
  NOR3_X1 u1_u10_u2_U12 (.A1( u1_u10_u2_n150 ) , .ZN( u1_u10_u2_n151 ) , .A3( u1_u10_u2_n175 ) , .A2( u1_u10_u2_n188 ) );
  AOI21_X1 u1_u10_u2_U13 (.ZN( u1_u10_u2_n144 ) , .B2( u1_u10_u2_n155 ) , .A( u1_u10_u2_n172 ) , .B1( u1_u10_u2_n185 ) );
  AOI21_X1 u1_u10_u2_U14 (.B2( u1_u10_u2_n143 ) , .ZN( u1_u10_u2_n145 ) , .B1( u1_u10_u2_n152 ) , .A( u1_u10_u2_n171 ) );
  AOI21_X1 u1_u10_u2_U15 (.B2( u1_u10_u2_n120 ) , .B1( u1_u10_u2_n121 ) , .ZN( u1_u10_u2_n126 ) , .A( u1_u10_u2_n167 ) );
  INV_X1 u1_u10_u2_U16 (.A( u1_u10_u2_n156 ) , .ZN( u1_u10_u2_n171 ) );
  INV_X1 u1_u10_u2_U17 (.A( u1_u10_u2_n120 ) , .ZN( u1_u10_u2_n188 ) );
  NAND2_X1 u1_u10_u2_U18 (.A2( u1_u10_u2_n122 ) , .ZN( u1_u10_u2_n150 ) , .A1( u1_u10_u2_n152 ) );
  INV_X1 u1_u10_u2_U19 (.A( u1_u10_u2_n153 ) , .ZN( u1_u10_u2_n170 ) );
  INV_X1 u1_u10_u2_U20 (.A( u1_u10_u2_n137 ) , .ZN( u1_u10_u2_n173 ) );
  NAND2_X1 u1_u10_u2_U21 (.A1( u1_u10_u2_n132 ) , .A2( u1_u10_u2_n139 ) , .ZN( u1_u10_u2_n157 ) );
  INV_X1 u1_u10_u2_U22 (.A( u1_u10_u2_n113 ) , .ZN( u1_u10_u2_n178 ) );
  INV_X1 u1_u10_u2_U23 (.A( u1_u10_u2_n139 ) , .ZN( u1_u10_u2_n175 ) );
  INV_X1 u1_u10_u2_U24 (.A( u1_u10_u2_n155 ) , .ZN( u1_u10_u2_n181 ) );
  INV_X1 u1_u10_u2_U25 (.A( u1_u10_u2_n119 ) , .ZN( u1_u10_u2_n177 ) );
  INV_X1 u1_u10_u2_U26 (.A( u1_u10_u2_n116 ) , .ZN( u1_u10_u2_n180 ) );
  INV_X1 u1_u10_u2_U27 (.A( u1_u10_u2_n131 ) , .ZN( u1_u10_u2_n179 ) );
  INV_X1 u1_u10_u2_U28 (.A( u1_u10_u2_n154 ) , .ZN( u1_u10_u2_n176 ) );
  NAND2_X1 u1_u10_u2_U29 (.A2( u1_u10_u2_n116 ) , .A1( u1_u10_u2_n117 ) , .ZN( u1_u10_u2_n118 ) );
  NOR2_X1 u1_u10_u2_U3 (.ZN( u1_u10_u2_n121 ) , .A2( u1_u10_u2_n177 ) , .A1( u1_u10_u2_n180 ) );
  INV_X1 u1_u10_u2_U30 (.A( u1_u10_u2_n132 ) , .ZN( u1_u10_u2_n182 ) );
  INV_X1 u1_u10_u2_U31 (.A( u1_u10_u2_n158 ) , .ZN( u1_u10_u2_n183 ) );
  OAI21_X1 u1_u10_u2_U32 (.A( u1_u10_u2_n156 ) , .B1( u1_u10_u2_n157 ) , .ZN( u1_u10_u2_n158 ) , .B2( u1_u10_u2_n179 ) );
  NOR2_X1 u1_u10_u2_U33 (.ZN( u1_u10_u2_n156 ) , .A1( u1_u10_u2_n166 ) , .A2( u1_u10_u2_n169 ) );
  NOR2_X1 u1_u10_u2_U34 (.A2( u1_u10_u2_n114 ) , .ZN( u1_u10_u2_n137 ) , .A1( u1_u10_u2_n140 ) );
  NOR2_X1 u1_u10_u2_U35 (.A2( u1_u10_u2_n138 ) , .ZN( u1_u10_u2_n153 ) , .A1( u1_u10_u2_n156 ) );
  AOI211_X1 u1_u10_u2_U36 (.ZN( u1_u10_u2_n130 ) , .C1( u1_u10_u2_n138 ) , .C2( u1_u10_u2_n179 ) , .B( u1_u10_u2_n96 ) , .A( u1_u10_u2_n97 ) );
  OAI22_X1 u1_u10_u2_U37 (.B1( u1_u10_u2_n133 ) , .A2( u1_u10_u2_n137 ) , .A1( u1_u10_u2_n152 ) , .B2( u1_u10_u2_n168 ) , .ZN( u1_u10_u2_n97 ) );
  OAI221_X1 u1_u10_u2_U38 (.B1( u1_u10_u2_n113 ) , .C1( u1_u10_u2_n132 ) , .A( u1_u10_u2_n149 ) , .B2( u1_u10_u2_n171 ) , .C2( u1_u10_u2_n172 ) , .ZN( u1_u10_u2_n96 ) );
  OAI221_X1 u1_u10_u2_U39 (.A( u1_u10_u2_n115 ) , .C2( u1_u10_u2_n123 ) , .B2( u1_u10_u2_n143 ) , .B1( u1_u10_u2_n153 ) , .ZN( u1_u10_u2_n163 ) , .C1( u1_u10_u2_n168 ) );
  INV_X1 u1_u10_u2_U4 (.A( u1_u10_u2_n134 ) , .ZN( u1_u10_u2_n185 ) );
  OAI21_X1 u1_u10_u2_U40 (.A( u1_u10_u2_n114 ) , .ZN( u1_u10_u2_n115 ) , .B1( u1_u10_u2_n176 ) , .B2( u1_u10_u2_n178 ) );
  OAI221_X1 u1_u10_u2_U41 (.A( u1_u10_u2_n135 ) , .B2( u1_u10_u2_n136 ) , .B1( u1_u10_u2_n137 ) , .ZN( u1_u10_u2_n162 ) , .C2( u1_u10_u2_n167 ) , .C1( u1_u10_u2_n185 ) );
  AND3_X1 u1_u10_u2_U42 (.A3( u1_u10_u2_n131 ) , .A2( u1_u10_u2_n132 ) , .A1( u1_u10_u2_n133 ) , .ZN( u1_u10_u2_n136 ) );
  AOI22_X1 u1_u10_u2_U43 (.ZN( u1_u10_u2_n135 ) , .B1( u1_u10_u2_n140 ) , .A1( u1_u10_u2_n156 ) , .B2( u1_u10_u2_n180 ) , .A2( u1_u10_u2_n188 ) );
  AOI21_X1 u1_u10_u2_U44 (.ZN( u1_u10_u2_n149 ) , .B1( u1_u10_u2_n173 ) , .B2( u1_u10_u2_n188 ) , .A( u1_u10_u2_n95 ) );
  AND3_X1 u1_u10_u2_U45 (.A2( u1_u10_u2_n100 ) , .A1( u1_u10_u2_n104 ) , .A3( u1_u10_u2_n156 ) , .ZN( u1_u10_u2_n95 ) );
  OAI21_X1 u1_u10_u2_U46 (.A( u1_u10_u2_n101 ) , .B2( u1_u10_u2_n121 ) , .B1( u1_u10_u2_n153 ) , .ZN( u1_u10_u2_n164 ) );
  NAND2_X1 u1_u10_u2_U47 (.A2( u1_u10_u2_n100 ) , .A1( u1_u10_u2_n107 ) , .ZN( u1_u10_u2_n155 ) );
  NAND2_X1 u1_u10_u2_U48 (.A2( u1_u10_u2_n105 ) , .A1( u1_u10_u2_n108 ) , .ZN( u1_u10_u2_n143 ) );
  NAND2_X1 u1_u10_u2_U49 (.A1( u1_u10_u2_n104 ) , .A2( u1_u10_u2_n106 ) , .ZN( u1_u10_u2_n152 ) );
  INV_X1 u1_u10_u2_U5 (.A( u1_u10_u2_n150 ) , .ZN( u1_u10_u2_n184 ) );
  NAND2_X1 u1_u10_u2_U50 (.A1( u1_u10_u2_n100 ) , .A2( u1_u10_u2_n105 ) , .ZN( u1_u10_u2_n132 ) );
  INV_X1 u1_u10_u2_U51 (.A( u1_u10_u2_n140 ) , .ZN( u1_u10_u2_n168 ) );
  INV_X1 u1_u10_u2_U52 (.A( u1_u10_u2_n138 ) , .ZN( u1_u10_u2_n167 ) );
  OAI21_X1 u1_u10_u2_U53 (.A( u1_u10_u2_n141 ) , .B2( u1_u10_u2_n142 ) , .ZN( u1_u10_u2_n146 ) , .B1( u1_u10_u2_n153 ) );
  OAI21_X1 u1_u10_u2_U54 (.A( u1_u10_u2_n140 ) , .ZN( u1_u10_u2_n141 ) , .B1( u1_u10_u2_n176 ) , .B2( u1_u10_u2_n177 ) );
  NOR3_X1 u1_u10_u2_U55 (.ZN( u1_u10_u2_n142 ) , .A3( u1_u10_u2_n175 ) , .A2( u1_u10_u2_n178 ) , .A1( u1_u10_u2_n181 ) );
  NAND2_X1 u1_u10_u2_U56 (.A1( u1_u10_u2_n102 ) , .A2( u1_u10_u2_n106 ) , .ZN( u1_u10_u2_n113 ) );
  NAND2_X1 u1_u10_u2_U57 (.A1( u1_u10_u2_n106 ) , .A2( u1_u10_u2_n107 ) , .ZN( u1_u10_u2_n131 ) );
  NAND2_X1 u1_u10_u2_U58 (.A1( u1_u10_u2_n103 ) , .A2( u1_u10_u2_n107 ) , .ZN( u1_u10_u2_n139 ) );
  NAND2_X1 u1_u10_u2_U59 (.A1( u1_u10_u2_n103 ) , .A2( u1_u10_u2_n105 ) , .ZN( u1_u10_u2_n133 ) );
  NOR4_X1 u1_u10_u2_U6 (.A4( u1_u10_u2_n124 ) , .A3( u1_u10_u2_n125 ) , .A2( u1_u10_u2_n126 ) , .A1( u1_u10_u2_n127 ) , .ZN( u1_u10_u2_n128 ) );
  NAND2_X1 u1_u10_u2_U60 (.A1( u1_u10_u2_n102 ) , .A2( u1_u10_u2_n103 ) , .ZN( u1_u10_u2_n154 ) );
  NAND2_X1 u1_u10_u2_U61 (.A2( u1_u10_u2_n103 ) , .A1( u1_u10_u2_n104 ) , .ZN( u1_u10_u2_n119 ) );
  NAND2_X1 u1_u10_u2_U62 (.A2( u1_u10_u2_n107 ) , .A1( u1_u10_u2_n108 ) , .ZN( u1_u10_u2_n123 ) );
  NAND2_X1 u1_u10_u2_U63 (.A1( u1_u10_u2_n104 ) , .A2( u1_u10_u2_n108 ) , .ZN( u1_u10_u2_n122 ) );
  INV_X1 u1_u10_u2_U64 (.A( u1_u10_u2_n114 ) , .ZN( u1_u10_u2_n172 ) );
  NAND2_X1 u1_u10_u2_U65 (.A2( u1_u10_u2_n100 ) , .A1( u1_u10_u2_n102 ) , .ZN( u1_u10_u2_n116 ) );
  NAND2_X1 u1_u10_u2_U66 (.A1( u1_u10_u2_n102 ) , .A2( u1_u10_u2_n108 ) , .ZN( u1_u10_u2_n120 ) );
  NAND2_X1 u1_u10_u2_U67 (.A2( u1_u10_u2_n105 ) , .A1( u1_u10_u2_n106 ) , .ZN( u1_u10_u2_n117 ) );
  INV_X1 u1_u10_u2_U68 (.ZN( u1_u10_u2_n187 ) , .A( u1_u10_u2_n99 ) );
  OAI21_X1 u1_u10_u2_U69 (.B1( u1_u10_u2_n137 ) , .B2( u1_u10_u2_n143 ) , .A( u1_u10_u2_n98 ) , .ZN( u1_u10_u2_n99 ) );
  AOI21_X1 u1_u10_u2_U7 (.ZN( u1_u10_u2_n124 ) , .B1( u1_u10_u2_n131 ) , .B2( u1_u10_u2_n143 ) , .A( u1_u10_u2_n172 ) );
  NOR2_X1 u1_u10_u2_U70 (.A2( u1_u10_X_16 ) , .ZN( u1_u10_u2_n140 ) , .A1( u1_u10_u2_n166 ) );
  NOR2_X1 u1_u10_u2_U71 (.A2( u1_u10_X_13 ) , .A1( u1_u10_X_14 ) , .ZN( u1_u10_u2_n100 ) );
  NOR2_X1 u1_u10_u2_U72 (.A2( u1_u10_X_16 ) , .A1( u1_u10_X_17 ) , .ZN( u1_u10_u2_n138 ) );
  NOR2_X1 u1_u10_u2_U73 (.A2( u1_u10_X_15 ) , .A1( u1_u10_X_18 ) , .ZN( u1_u10_u2_n104 ) );
  NOR2_X1 u1_u10_u2_U74 (.A2( u1_u10_X_14 ) , .ZN( u1_u10_u2_n103 ) , .A1( u1_u10_u2_n174 ) );
  NOR2_X1 u1_u10_u2_U75 (.A2( u1_u10_X_15 ) , .ZN( u1_u10_u2_n102 ) , .A1( u1_u10_u2_n165 ) );
  NOR2_X1 u1_u10_u2_U76 (.A2( u1_u10_X_17 ) , .ZN( u1_u10_u2_n114 ) , .A1( u1_u10_u2_n169 ) );
  AND2_X1 u1_u10_u2_U77 (.A1( u1_u10_X_15 ) , .ZN( u1_u10_u2_n105 ) , .A2( u1_u10_u2_n165 ) );
  AND2_X1 u1_u10_u2_U78 (.A2( u1_u10_X_15 ) , .A1( u1_u10_X_18 ) , .ZN( u1_u10_u2_n107 ) );
  AND2_X1 u1_u10_u2_U79 (.A1( u1_u10_X_14 ) , .ZN( u1_u10_u2_n106 ) , .A2( u1_u10_u2_n174 ) );
  AOI21_X1 u1_u10_u2_U8 (.B2( u1_u10_u2_n119 ) , .ZN( u1_u10_u2_n127 ) , .A( u1_u10_u2_n137 ) , .B1( u1_u10_u2_n155 ) );
  AND2_X1 u1_u10_u2_U80 (.A1( u1_u10_X_13 ) , .A2( u1_u10_X_14 ) , .ZN( u1_u10_u2_n108 ) );
  INV_X1 u1_u10_u2_U81 (.A( u1_u10_X_16 ) , .ZN( u1_u10_u2_n169 ) );
  INV_X1 u1_u10_u2_U82 (.A( u1_u10_X_17 ) , .ZN( u1_u10_u2_n166 ) );
  INV_X1 u1_u10_u2_U83 (.A( u1_u10_X_13 ) , .ZN( u1_u10_u2_n174 ) );
  INV_X1 u1_u10_u2_U84 (.A( u1_u10_X_18 ) , .ZN( u1_u10_u2_n165 ) );
  NAND4_X1 u1_u10_u2_U85 (.ZN( u1_out10_30 ) , .A4( u1_u10_u2_n147 ) , .A3( u1_u10_u2_n148 ) , .A2( u1_u10_u2_n149 ) , .A1( u1_u10_u2_n187 ) );
  NOR3_X1 u1_u10_u2_U86 (.A3( u1_u10_u2_n144 ) , .A2( u1_u10_u2_n145 ) , .A1( u1_u10_u2_n146 ) , .ZN( u1_u10_u2_n147 ) );
  AOI21_X1 u1_u10_u2_U87 (.B2( u1_u10_u2_n138 ) , .ZN( u1_u10_u2_n148 ) , .A( u1_u10_u2_n162 ) , .B1( u1_u10_u2_n182 ) );
  NAND4_X1 u1_u10_u2_U88 (.ZN( u1_out10_24 ) , .A4( u1_u10_u2_n111 ) , .A3( u1_u10_u2_n112 ) , .A1( u1_u10_u2_n130 ) , .A2( u1_u10_u2_n187 ) );
  AOI221_X1 u1_u10_u2_U89 (.A( u1_u10_u2_n109 ) , .B1( u1_u10_u2_n110 ) , .ZN( u1_u10_u2_n111 ) , .C1( u1_u10_u2_n134 ) , .C2( u1_u10_u2_n170 ) , .B2( u1_u10_u2_n173 ) );
  AOI21_X1 u1_u10_u2_U9 (.B2( u1_u10_u2_n123 ) , .ZN( u1_u10_u2_n125 ) , .A( u1_u10_u2_n171 ) , .B1( u1_u10_u2_n184 ) );
  AOI21_X1 u1_u10_u2_U90 (.ZN( u1_u10_u2_n112 ) , .B2( u1_u10_u2_n156 ) , .A( u1_u10_u2_n164 ) , .B1( u1_u10_u2_n181 ) );
  NAND4_X1 u1_u10_u2_U91 (.ZN( u1_out10_16 ) , .A4( u1_u10_u2_n128 ) , .A3( u1_u10_u2_n129 ) , .A1( u1_u10_u2_n130 ) , .A2( u1_u10_u2_n186 ) );
  AOI22_X1 u1_u10_u2_U92 (.A2( u1_u10_u2_n118 ) , .ZN( u1_u10_u2_n129 ) , .A1( u1_u10_u2_n140 ) , .B1( u1_u10_u2_n157 ) , .B2( u1_u10_u2_n170 ) );
  INV_X1 u1_u10_u2_U93 (.A( u1_u10_u2_n163 ) , .ZN( u1_u10_u2_n186 ) );
  OR4_X1 u1_u10_u2_U94 (.ZN( u1_out10_6 ) , .A4( u1_u10_u2_n161 ) , .A3( u1_u10_u2_n162 ) , .A2( u1_u10_u2_n163 ) , .A1( u1_u10_u2_n164 ) );
  OR3_X1 u1_u10_u2_U95 (.A2( u1_u10_u2_n159 ) , .A1( u1_u10_u2_n160 ) , .ZN( u1_u10_u2_n161 ) , .A3( u1_u10_u2_n183 ) );
  AOI21_X1 u1_u10_u2_U96 (.B2( u1_u10_u2_n154 ) , .B1( u1_u10_u2_n155 ) , .ZN( u1_u10_u2_n159 ) , .A( u1_u10_u2_n167 ) );
  NAND3_X1 u1_u10_u2_U97 (.A2( u1_u10_u2_n117 ) , .A1( u1_u10_u2_n122 ) , .A3( u1_u10_u2_n123 ) , .ZN( u1_u10_u2_n134 ) );
  NAND3_X1 u1_u10_u2_U98 (.ZN( u1_u10_u2_n110 ) , .A2( u1_u10_u2_n131 ) , .A3( u1_u10_u2_n139 ) , .A1( u1_u10_u2_n154 ) );
  NAND3_X1 u1_u10_u2_U99 (.A2( u1_u10_u2_n100 ) , .ZN( u1_u10_u2_n101 ) , .A1( u1_u10_u2_n104 ) , .A3( u1_u10_u2_n114 ) );
  XOR2_X1 u1_u11_U1 (.B( u1_K12_9 ) , .A( u1_R10_6 ) , .Z( u1_u11_X_9 ) );
  XOR2_X1 u1_u11_U16 (.B( u1_K12_3 ) , .A( u1_R10_2 ) , .Z( u1_u11_X_3 ) );
  XOR2_X1 u1_u11_U3 (.B( u1_K12_7 ) , .A( u1_R10_4 ) , .Z( u1_u11_X_7 ) );
  XOR2_X1 u1_u11_U42 (.B( u1_K12_16 ) , .A( u1_R10_11 ) , .Z( u1_u11_X_16 ) );
  XOR2_X1 u1_u11_U43 (.B( u1_K12_15 ) , .A( u1_R10_10 ) , .Z( u1_u11_X_15 ) );
  XOR2_X1 u1_u11_U44 (.B( u1_K12_14 ) , .A( u1_R10_9 ) , .Z( u1_u11_X_14 ) );
  XOR2_X1 u1_u11_U45 (.B( u1_K12_13 ) , .A( u1_R10_8 ) , .Z( u1_u11_X_13 ) );
  XOR2_X1 u1_u11_U46 (.B( u1_K12_12 ) , .A( u1_R10_9 ) , .Z( u1_u11_X_12 ) );
  XOR2_X1 u1_u11_U47 (.B( u1_K12_11 ) , .A( u1_R10_8 ) , .Z( u1_u11_X_11 ) );
  XOR2_X1 u1_u11_U48 (.B( u1_K12_10 ) , .A( u1_R10_7 ) , .Z( u1_u11_X_10 ) );
  XOR2_X1 u1_u11_U5 (.B( u1_K12_5 ) , .A( u1_R10_4 ) , .Z( u1_u11_X_5 ) );
  XOR2_X1 u1_u11_U6 (.B( u1_K12_4 ) , .A( u1_R10_3 ) , .Z( u1_u11_X_4 ) );
  NAND2_X1 u1_u11_u0_U10 (.ZN( u1_u11_u0_n113 ) , .A1( u1_u11_u0_n139 ) , .A2( u1_u11_u0_n149 ) );
  AND3_X1 u1_u11_u0_U11 (.A2( u1_u11_u0_n112 ) , .ZN( u1_u11_u0_n127 ) , .A3( u1_u11_u0_n130 ) , .A1( u1_u11_u0_n148 ) );
  AND2_X1 u1_u11_u0_U12 (.ZN( u1_u11_u0_n107 ) , .A1( u1_u11_u0_n130 ) , .A2( u1_u11_u0_n140 ) );
  AND2_X1 u1_u11_u0_U13 (.A2( u1_u11_u0_n129 ) , .A1( u1_u11_u0_n130 ) , .ZN( u1_u11_u0_n151 ) );
  AND2_X1 u1_u11_u0_U14 (.A1( u1_u11_u0_n108 ) , .A2( u1_u11_u0_n125 ) , .ZN( u1_u11_u0_n145 ) );
  INV_X1 u1_u11_u0_U15 (.A( u1_u11_u0_n143 ) , .ZN( u1_u11_u0_n173 ) );
  NOR2_X1 u1_u11_u0_U16 (.A2( u1_u11_u0_n136 ) , .ZN( u1_u11_u0_n147 ) , .A1( u1_u11_u0_n160 ) );
  OAI22_X1 u1_u11_u0_U17 (.B1( u1_u11_u0_n131 ) , .A1( u1_u11_u0_n144 ) , .B2( u1_u11_u0_n147 ) , .A2( u1_u11_u0_n90 ) , .ZN( u1_u11_u0_n91 ) );
  AND3_X1 u1_u11_u0_U18 (.A3( u1_u11_u0_n121 ) , .A2( u1_u11_u0_n125 ) , .A1( u1_u11_u0_n148 ) , .ZN( u1_u11_u0_n90 ) );
  OAI22_X1 u1_u11_u0_U19 (.B1( u1_u11_u0_n125 ) , .ZN( u1_u11_u0_n126 ) , .A1( u1_u11_u0_n138 ) , .A2( u1_u11_u0_n146 ) , .B2( u1_u11_u0_n147 ) );
  NOR2_X1 u1_u11_u0_U20 (.A1( u1_u11_u0_n163 ) , .A2( u1_u11_u0_n164 ) , .ZN( u1_u11_u0_n95 ) );
  NAND2_X1 u1_u11_u0_U21 (.A1( u1_u11_u0_n101 ) , .A2( u1_u11_u0_n102 ) , .ZN( u1_u11_u0_n150 ) );
  AOI22_X1 u1_u11_u0_U22 (.B2( u1_u11_u0_n109 ) , .A2( u1_u11_u0_n110 ) , .ZN( u1_u11_u0_n111 ) , .B1( u1_u11_u0_n118 ) , .A1( u1_u11_u0_n160 ) );
  INV_X1 u1_u11_u0_U23 (.A( u1_u11_u0_n136 ) , .ZN( u1_u11_u0_n161 ) );
  INV_X1 u1_u11_u0_U24 (.A( u1_u11_u0_n118 ) , .ZN( u1_u11_u0_n158 ) );
  NAND2_X1 u1_u11_u0_U25 (.A2( u1_u11_u0_n100 ) , .A1( u1_u11_u0_n101 ) , .ZN( u1_u11_u0_n139 ) );
  NAND2_X1 u1_u11_u0_U26 (.A2( u1_u11_u0_n100 ) , .ZN( u1_u11_u0_n131 ) , .A1( u1_u11_u0_n92 ) );
  NAND2_X1 u1_u11_u0_U27 (.ZN( u1_u11_u0_n108 ) , .A1( u1_u11_u0_n92 ) , .A2( u1_u11_u0_n94 ) );
  AOI21_X1 u1_u11_u0_U28 (.ZN( u1_u11_u0_n104 ) , .B1( u1_u11_u0_n107 ) , .B2( u1_u11_u0_n141 ) , .A( u1_u11_u0_n144 ) );
  AOI21_X1 u1_u11_u0_U29 (.B1( u1_u11_u0_n127 ) , .B2( u1_u11_u0_n129 ) , .A( u1_u11_u0_n138 ) , .ZN( u1_u11_u0_n96 ) );
  INV_X1 u1_u11_u0_U3 (.A( u1_u11_u0_n113 ) , .ZN( u1_u11_u0_n166 ) );
  NAND2_X1 u1_u11_u0_U30 (.A2( u1_u11_u0_n102 ) , .ZN( u1_u11_u0_n114 ) , .A1( u1_u11_u0_n92 ) );
  NAND2_X1 u1_u11_u0_U31 (.A1( u1_u11_u0_n101 ) , .ZN( u1_u11_u0_n130 ) , .A2( u1_u11_u0_n94 ) );
  NOR2_X1 u1_u11_u0_U32 (.A1( u1_u11_u0_n120 ) , .ZN( u1_u11_u0_n143 ) , .A2( u1_u11_u0_n167 ) );
  OAI221_X1 u1_u11_u0_U33 (.C1( u1_u11_u0_n112 ) , .ZN( u1_u11_u0_n120 ) , .B1( u1_u11_u0_n138 ) , .B2( u1_u11_u0_n141 ) , .C2( u1_u11_u0_n147 ) , .A( u1_u11_u0_n172 ) );
  AOI211_X1 u1_u11_u0_U34 (.B( u1_u11_u0_n115 ) , .A( u1_u11_u0_n116 ) , .C2( u1_u11_u0_n117 ) , .C1( u1_u11_u0_n118 ) , .ZN( u1_u11_u0_n119 ) );
  NAND2_X1 u1_u11_u0_U35 (.A1( u1_u11_u0_n100 ) , .A2( u1_u11_u0_n103 ) , .ZN( u1_u11_u0_n125 ) );
  NAND2_X1 u1_u11_u0_U36 (.A2( u1_u11_u0_n103 ) , .ZN( u1_u11_u0_n140 ) , .A1( u1_u11_u0_n94 ) );
  INV_X1 u1_u11_u0_U37 (.A( u1_u11_u0_n138 ) , .ZN( u1_u11_u0_n160 ) );
  NAND2_X1 u1_u11_u0_U38 (.A2( u1_u11_u0_n102 ) , .A1( u1_u11_u0_n103 ) , .ZN( u1_u11_u0_n149 ) );
  NAND2_X1 u1_u11_u0_U39 (.A2( u1_u11_u0_n101 ) , .ZN( u1_u11_u0_n121 ) , .A1( u1_u11_u0_n93 ) );
  AOI21_X1 u1_u11_u0_U4 (.B1( u1_u11_u0_n114 ) , .ZN( u1_u11_u0_n115 ) , .B2( u1_u11_u0_n129 ) , .A( u1_u11_u0_n161 ) );
  NAND2_X1 u1_u11_u0_U40 (.ZN( u1_u11_u0_n112 ) , .A2( u1_u11_u0_n92 ) , .A1( u1_u11_u0_n93 ) );
  INV_X1 u1_u11_u0_U41 (.ZN( u1_u11_u0_n172 ) , .A( u1_u11_u0_n88 ) );
  OAI222_X1 u1_u11_u0_U42 (.C1( u1_u11_u0_n108 ) , .A1( u1_u11_u0_n125 ) , .B2( u1_u11_u0_n128 ) , .B1( u1_u11_u0_n144 ) , .A2( u1_u11_u0_n158 ) , .C2( u1_u11_u0_n161 ) , .ZN( u1_u11_u0_n88 ) );
  AOI21_X1 u1_u11_u0_U43 (.B1( u1_u11_u0_n103 ) , .ZN( u1_u11_u0_n132 ) , .A( u1_u11_u0_n165 ) , .B2( u1_u11_u0_n93 ) );
  OR3_X1 u1_u11_u0_U44 (.A3( u1_u11_u0_n152 ) , .A2( u1_u11_u0_n153 ) , .A1( u1_u11_u0_n154 ) , .ZN( u1_u11_u0_n155 ) );
  AOI21_X1 u1_u11_u0_U45 (.A( u1_u11_u0_n144 ) , .B2( u1_u11_u0_n145 ) , .B1( u1_u11_u0_n146 ) , .ZN( u1_u11_u0_n154 ) );
  AOI21_X1 u1_u11_u0_U46 (.B2( u1_u11_u0_n150 ) , .B1( u1_u11_u0_n151 ) , .ZN( u1_u11_u0_n152 ) , .A( u1_u11_u0_n158 ) );
  AOI21_X1 u1_u11_u0_U47 (.A( u1_u11_u0_n147 ) , .B2( u1_u11_u0_n148 ) , .B1( u1_u11_u0_n149 ) , .ZN( u1_u11_u0_n153 ) );
  INV_X1 u1_u11_u0_U48 (.ZN( u1_u11_u0_n171 ) , .A( u1_u11_u0_n99 ) );
  OAI211_X1 u1_u11_u0_U49 (.C2( u1_u11_u0_n140 ) , .C1( u1_u11_u0_n161 ) , .A( u1_u11_u0_n169 ) , .B( u1_u11_u0_n98 ) , .ZN( u1_u11_u0_n99 ) );
  AOI21_X1 u1_u11_u0_U5 (.B2( u1_u11_u0_n131 ) , .ZN( u1_u11_u0_n134 ) , .B1( u1_u11_u0_n151 ) , .A( u1_u11_u0_n158 ) );
  AOI211_X1 u1_u11_u0_U50 (.C1( u1_u11_u0_n118 ) , .A( u1_u11_u0_n123 ) , .B( u1_u11_u0_n96 ) , .C2( u1_u11_u0_n97 ) , .ZN( u1_u11_u0_n98 ) );
  INV_X1 u1_u11_u0_U51 (.ZN( u1_u11_u0_n169 ) , .A( u1_u11_u0_n91 ) );
  NOR2_X1 u1_u11_u0_U52 (.A2( u1_u11_X_2 ) , .ZN( u1_u11_u0_n103 ) , .A1( u1_u11_u0_n164 ) );
  NOR2_X1 u1_u11_u0_U53 (.A2( u1_u11_X_4 ) , .A1( u1_u11_X_5 ) , .ZN( u1_u11_u0_n118 ) );
  NOR2_X1 u1_u11_u0_U54 (.A2( u1_u11_X_3 ) , .A1( u1_u11_X_6 ) , .ZN( u1_u11_u0_n94 ) );
  NOR2_X1 u1_u11_u0_U55 (.A2( u1_u11_X_6 ) , .ZN( u1_u11_u0_n100 ) , .A1( u1_u11_u0_n162 ) );
  NAND2_X1 u1_u11_u0_U56 (.A2( u1_u11_X_4 ) , .A1( u1_u11_X_5 ) , .ZN( u1_u11_u0_n144 ) );
  NOR2_X1 u1_u11_u0_U57 (.A2( u1_u11_X_5 ) , .ZN( u1_u11_u0_n136 ) , .A1( u1_u11_u0_n159 ) );
  NAND2_X1 u1_u11_u0_U58 (.A1( u1_u11_X_5 ) , .ZN( u1_u11_u0_n138 ) , .A2( u1_u11_u0_n159 ) );
  AND2_X1 u1_u11_u0_U59 (.A2( u1_u11_X_3 ) , .A1( u1_u11_X_6 ) , .ZN( u1_u11_u0_n102 ) );
  NOR2_X1 u1_u11_u0_U6 (.A1( u1_u11_u0_n108 ) , .ZN( u1_u11_u0_n123 ) , .A2( u1_u11_u0_n158 ) );
  AND2_X1 u1_u11_u0_U60 (.A1( u1_u11_X_6 ) , .A2( u1_u11_u0_n162 ) , .ZN( u1_u11_u0_n93 ) );
  INV_X1 u1_u11_u0_U61 (.A( u1_u11_X_4 ) , .ZN( u1_u11_u0_n159 ) );
  INV_X1 u1_u11_u0_U62 (.A( u1_u11_X_3 ) , .ZN( u1_u11_u0_n162 ) );
  INV_X1 u1_u11_u0_U63 (.A( u1_u11_X_2 ) , .ZN( u1_u11_u0_n163 ) );
  AOI211_X1 u1_u11_u0_U64 (.B( u1_u11_u0_n133 ) , .A( u1_u11_u0_n134 ) , .C2( u1_u11_u0_n135 ) , .C1( u1_u11_u0_n136 ) , .ZN( u1_u11_u0_n137 ) );
  INV_X1 u1_u11_u0_U65 (.A( u1_u11_u0_n126 ) , .ZN( u1_u11_u0_n168 ) );
  OR4_X1 u1_u11_u0_U66 (.ZN( u1_out11_17 ) , .A4( u1_u11_u0_n122 ) , .A2( u1_u11_u0_n123 ) , .A1( u1_u11_u0_n124 ) , .A3( u1_u11_u0_n170 ) );
  AOI21_X1 u1_u11_u0_U67 (.B2( u1_u11_u0_n107 ) , .ZN( u1_u11_u0_n124 ) , .B1( u1_u11_u0_n128 ) , .A( u1_u11_u0_n161 ) );
  INV_X1 u1_u11_u0_U68 (.A( u1_u11_u0_n111 ) , .ZN( u1_u11_u0_n170 ) );
  OR4_X1 u1_u11_u0_U69 (.ZN( u1_out11_31 ) , .A4( u1_u11_u0_n155 ) , .A2( u1_u11_u0_n156 ) , .A1( u1_u11_u0_n157 ) , .A3( u1_u11_u0_n173 ) );
  OAI21_X1 u1_u11_u0_U7 (.B1( u1_u11_u0_n150 ) , .B2( u1_u11_u0_n158 ) , .A( u1_u11_u0_n172 ) , .ZN( u1_u11_u0_n89 ) );
  AOI21_X1 u1_u11_u0_U70 (.A( u1_u11_u0_n138 ) , .B2( u1_u11_u0_n139 ) , .B1( u1_u11_u0_n140 ) , .ZN( u1_u11_u0_n157 ) );
  INV_X1 u1_u11_u0_U71 (.ZN( u1_u11_u0_n174 ) , .A( u1_u11_u0_n89 ) );
  AOI211_X1 u1_u11_u0_U72 (.B( u1_u11_u0_n104 ) , .A( u1_u11_u0_n105 ) , .ZN( u1_u11_u0_n106 ) , .C2( u1_u11_u0_n113 ) , .C1( u1_u11_u0_n160 ) );
  AOI21_X1 u1_u11_u0_U73 (.B2( u1_u11_u0_n141 ) , .B1( u1_u11_u0_n142 ) , .ZN( u1_u11_u0_n156 ) , .A( u1_u11_u0_n161 ) );
  AOI21_X1 u1_u11_u0_U74 (.ZN( u1_u11_u0_n116 ) , .B2( u1_u11_u0_n142 ) , .A( u1_u11_u0_n144 ) , .B1( u1_u11_u0_n166 ) );
  INV_X1 u1_u11_u0_U75 (.A( u1_u11_u0_n142 ) , .ZN( u1_u11_u0_n165 ) );
  NOR2_X1 u1_u11_u0_U76 (.A2( u1_u11_X_1 ) , .A1( u1_u11_X_2 ) , .ZN( u1_u11_u0_n92 ) );
  NOR2_X1 u1_u11_u0_U77 (.A2( u1_u11_X_1 ) , .ZN( u1_u11_u0_n101 ) , .A1( u1_u11_u0_n163 ) );
  INV_X1 u1_u11_u0_U78 (.A( u1_u11_X_1 ) , .ZN( u1_u11_u0_n164 ) );
  OAI221_X1 u1_u11_u0_U79 (.C1( u1_u11_u0_n121 ) , .ZN( u1_u11_u0_n122 ) , .B2( u1_u11_u0_n127 ) , .A( u1_u11_u0_n143 ) , .B1( u1_u11_u0_n144 ) , .C2( u1_u11_u0_n147 ) );
  AND2_X1 u1_u11_u0_U8 (.A1( u1_u11_u0_n114 ) , .A2( u1_u11_u0_n121 ) , .ZN( u1_u11_u0_n146 ) );
  AOI21_X1 u1_u11_u0_U80 (.B1( u1_u11_u0_n132 ) , .ZN( u1_u11_u0_n133 ) , .A( u1_u11_u0_n144 ) , .B2( u1_u11_u0_n166 ) );
  OAI22_X1 u1_u11_u0_U81 (.ZN( u1_u11_u0_n105 ) , .A2( u1_u11_u0_n132 ) , .B1( u1_u11_u0_n146 ) , .A1( u1_u11_u0_n147 ) , .B2( u1_u11_u0_n161 ) );
  NAND2_X1 u1_u11_u0_U82 (.ZN( u1_u11_u0_n110 ) , .A2( u1_u11_u0_n132 ) , .A1( u1_u11_u0_n145 ) );
  INV_X1 u1_u11_u0_U83 (.A( u1_u11_u0_n119 ) , .ZN( u1_u11_u0_n167 ) );
  NAND2_X1 u1_u11_u0_U84 (.ZN( u1_u11_u0_n148 ) , .A1( u1_u11_u0_n93 ) , .A2( u1_u11_u0_n95 ) );
  NAND2_X1 u1_u11_u0_U85 (.A1( u1_u11_u0_n100 ) , .ZN( u1_u11_u0_n129 ) , .A2( u1_u11_u0_n95 ) );
  NAND2_X1 u1_u11_u0_U86 (.A1( u1_u11_u0_n102 ) , .ZN( u1_u11_u0_n128 ) , .A2( u1_u11_u0_n95 ) );
  NAND2_X1 u1_u11_u0_U87 (.ZN( u1_u11_u0_n142 ) , .A1( u1_u11_u0_n94 ) , .A2( u1_u11_u0_n95 ) );
  NAND3_X1 u1_u11_u0_U88 (.ZN( u1_out11_23 ) , .A3( u1_u11_u0_n137 ) , .A1( u1_u11_u0_n168 ) , .A2( u1_u11_u0_n171 ) );
  NAND3_X1 u1_u11_u0_U89 (.A3( u1_u11_u0_n127 ) , .A2( u1_u11_u0_n128 ) , .ZN( u1_u11_u0_n135 ) , .A1( u1_u11_u0_n150 ) );
  AND2_X1 u1_u11_u0_U9 (.A1( u1_u11_u0_n131 ) , .ZN( u1_u11_u0_n141 ) , .A2( u1_u11_u0_n150 ) );
  NAND3_X1 u1_u11_u0_U90 (.ZN( u1_u11_u0_n117 ) , .A3( u1_u11_u0_n132 ) , .A2( u1_u11_u0_n139 ) , .A1( u1_u11_u0_n148 ) );
  NAND3_X1 u1_u11_u0_U91 (.ZN( u1_u11_u0_n109 ) , .A2( u1_u11_u0_n114 ) , .A3( u1_u11_u0_n140 ) , .A1( u1_u11_u0_n149 ) );
  NAND3_X1 u1_u11_u0_U92 (.ZN( u1_out11_9 ) , .A3( u1_u11_u0_n106 ) , .A2( u1_u11_u0_n171 ) , .A1( u1_u11_u0_n174 ) );
  NAND3_X1 u1_u11_u0_U93 (.A2( u1_u11_u0_n128 ) , .A1( u1_u11_u0_n132 ) , .A3( u1_u11_u0_n146 ) , .ZN( u1_u11_u0_n97 ) );
  NOR2_X1 u1_u11_u1_U10 (.A1( u1_u11_u1_n112 ) , .A2( u1_u11_u1_n116 ) , .ZN( u1_u11_u1_n118 ) );
  NAND3_X1 u1_u11_u1_U100 (.ZN( u1_u11_u1_n113 ) , .A1( u1_u11_u1_n120 ) , .A3( u1_u11_u1_n133 ) , .A2( u1_u11_u1_n155 ) );
  OAI21_X1 u1_u11_u1_U11 (.ZN( u1_u11_u1_n101 ) , .B1( u1_u11_u1_n141 ) , .A( u1_u11_u1_n146 ) , .B2( u1_u11_u1_n183 ) );
  AOI21_X1 u1_u11_u1_U12 (.B2( u1_u11_u1_n155 ) , .B1( u1_u11_u1_n156 ) , .ZN( u1_u11_u1_n157 ) , .A( u1_u11_u1_n174 ) );
  NAND2_X1 u1_u11_u1_U13 (.ZN( u1_u11_u1_n140 ) , .A2( u1_u11_u1_n150 ) , .A1( u1_u11_u1_n155 ) );
  NAND2_X1 u1_u11_u1_U14 (.A1( u1_u11_u1_n131 ) , .ZN( u1_u11_u1_n147 ) , .A2( u1_u11_u1_n153 ) );
  INV_X1 u1_u11_u1_U15 (.A( u1_u11_u1_n139 ) , .ZN( u1_u11_u1_n174 ) );
  OR4_X1 u1_u11_u1_U16 (.A4( u1_u11_u1_n106 ) , .A3( u1_u11_u1_n107 ) , .ZN( u1_u11_u1_n108 ) , .A1( u1_u11_u1_n117 ) , .A2( u1_u11_u1_n184 ) );
  AOI21_X1 u1_u11_u1_U17 (.ZN( u1_u11_u1_n106 ) , .A( u1_u11_u1_n112 ) , .B1( u1_u11_u1_n154 ) , .B2( u1_u11_u1_n156 ) );
  AOI21_X1 u1_u11_u1_U18 (.ZN( u1_u11_u1_n107 ) , .B1( u1_u11_u1_n134 ) , .B2( u1_u11_u1_n149 ) , .A( u1_u11_u1_n174 ) );
  INV_X1 u1_u11_u1_U19 (.A( u1_u11_u1_n101 ) , .ZN( u1_u11_u1_n184 ) );
  INV_X1 u1_u11_u1_U20 (.A( u1_u11_u1_n112 ) , .ZN( u1_u11_u1_n171 ) );
  NAND2_X1 u1_u11_u1_U21 (.ZN( u1_u11_u1_n141 ) , .A1( u1_u11_u1_n153 ) , .A2( u1_u11_u1_n156 ) );
  AND2_X1 u1_u11_u1_U22 (.A1( u1_u11_u1_n123 ) , .ZN( u1_u11_u1_n134 ) , .A2( u1_u11_u1_n161 ) );
  NAND2_X1 u1_u11_u1_U23 (.A2( u1_u11_u1_n115 ) , .A1( u1_u11_u1_n116 ) , .ZN( u1_u11_u1_n148 ) );
  NAND2_X1 u1_u11_u1_U24 (.A2( u1_u11_u1_n133 ) , .A1( u1_u11_u1_n135 ) , .ZN( u1_u11_u1_n159 ) );
  NAND2_X1 u1_u11_u1_U25 (.A2( u1_u11_u1_n115 ) , .A1( u1_u11_u1_n120 ) , .ZN( u1_u11_u1_n132 ) );
  INV_X1 u1_u11_u1_U26 (.A( u1_u11_u1_n154 ) , .ZN( u1_u11_u1_n178 ) );
  INV_X1 u1_u11_u1_U27 (.A( u1_u11_u1_n151 ) , .ZN( u1_u11_u1_n183 ) );
  AND2_X1 u1_u11_u1_U28 (.A1( u1_u11_u1_n129 ) , .A2( u1_u11_u1_n133 ) , .ZN( u1_u11_u1_n149 ) );
  INV_X1 u1_u11_u1_U29 (.A( u1_u11_u1_n131 ) , .ZN( u1_u11_u1_n180 ) );
  INV_X1 u1_u11_u1_U3 (.A( u1_u11_u1_n159 ) , .ZN( u1_u11_u1_n182 ) );
  OAI221_X1 u1_u11_u1_U30 (.A( u1_u11_u1_n119 ) , .C2( u1_u11_u1_n129 ) , .ZN( u1_u11_u1_n138 ) , .B2( u1_u11_u1_n152 ) , .C1( u1_u11_u1_n174 ) , .B1( u1_u11_u1_n187 ) );
  INV_X1 u1_u11_u1_U31 (.A( u1_u11_u1_n148 ) , .ZN( u1_u11_u1_n187 ) );
  AOI211_X1 u1_u11_u1_U32 (.B( u1_u11_u1_n117 ) , .A( u1_u11_u1_n118 ) , .ZN( u1_u11_u1_n119 ) , .C2( u1_u11_u1_n146 ) , .C1( u1_u11_u1_n159 ) );
  NOR2_X1 u1_u11_u1_U33 (.A1( u1_u11_u1_n168 ) , .A2( u1_u11_u1_n176 ) , .ZN( u1_u11_u1_n98 ) );
  AOI211_X1 u1_u11_u1_U34 (.B( u1_u11_u1_n162 ) , .A( u1_u11_u1_n163 ) , .C2( u1_u11_u1_n164 ) , .ZN( u1_u11_u1_n165 ) , .C1( u1_u11_u1_n171 ) );
  AOI21_X1 u1_u11_u1_U35 (.A( u1_u11_u1_n160 ) , .B2( u1_u11_u1_n161 ) , .ZN( u1_u11_u1_n162 ) , .B1( u1_u11_u1_n182 ) );
  OR2_X1 u1_u11_u1_U36 (.A2( u1_u11_u1_n157 ) , .A1( u1_u11_u1_n158 ) , .ZN( u1_u11_u1_n163 ) );
  NAND2_X1 u1_u11_u1_U37 (.A1( u1_u11_u1_n128 ) , .ZN( u1_u11_u1_n146 ) , .A2( u1_u11_u1_n160 ) );
  NAND2_X1 u1_u11_u1_U38 (.A2( u1_u11_u1_n112 ) , .ZN( u1_u11_u1_n139 ) , .A1( u1_u11_u1_n152 ) );
  NAND2_X1 u1_u11_u1_U39 (.A1( u1_u11_u1_n105 ) , .ZN( u1_u11_u1_n156 ) , .A2( u1_u11_u1_n99 ) );
  AOI221_X1 u1_u11_u1_U4 (.A( u1_u11_u1_n138 ) , .C2( u1_u11_u1_n139 ) , .C1( u1_u11_u1_n140 ) , .B2( u1_u11_u1_n141 ) , .ZN( u1_u11_u1_n142 ) , .B1( u1_u11_u1_n175 ) );
  AOI221_X1 u1_u11_u1_U40 (.B1( u1_u11_u1_n140 ) , .ZN( u1_u11_u1_n167 ) , .B2( u1_u11_u1_n172 ) , .C2( u1_u11_u1_n175 ) , .C1( u1_u11_u1_n178 ) , .A( u1_u11_u1_n188 ) );
  INV_X1 u1_u11_u1_U41 (.ZN( u1_u11_u1_n188 ) , .A( u1_u11_u1_n97 ) );
  AOI211_X1 u1_u11_u1_U42 (.A( u1_u11_u1_n118 ) , .C1( u1_u11_u1_n132 ) , .C2( u1_u11_u1_n139 ) , .B( u1_u11_u1_n96 ) , .ZN( u1_u11_u1_n97 ) );
  AOI21_X1 u1_u11_u1_U43 (.B2( u1_u11_u1_n121 ) , .B1( u1_u11_u1_n135 ) , .A( u1_u11_u1_n152 ) , .ZN( u1_u11_u1_n96 ) );
  NOR2_X1 u1_u11_u1_U44 (.ZN( u1_u11_u1_n117 ) , .A1( u1_u11_u1_n121 ) , .A2( u1_u11_u1_n160 ) );
  OAI21_X1 u1_u11_u1_U45 (.B2( u1_u11_u1_n123 ) , .ZN( u1_u11_u1_n145 ) , .B1( u1_u11_u1_n160 ) , .A( u1_u11_u1_n185 ) );
  INV_X1 u1_u11_u1_U46 (.A( u1_u11_u1_n122 ) , .ZN( u1_u11_u1_n185 ) );
  AOI21_X1 u1_u11_u1_U47 (.B2( u1_u11_u1_n120 ) , .B1( u1_u11_u1_n121 ) , .ZN( u1_u11_u1_n122 ) , .A( u1_u11_u1_n128 ) );
  AOI21_X1 u1_u11_u1_U48 (.A( u1_u11_u1_n128 ) , .B2( u1_u11_u1_n129 ) , .ZN( u1_u11_u1_n130 ) , .B1( u1_u11_u1_n150 ) );
  NAND2_X1 u1_u11_u1_U49 (.ZN( u1_u11_u1_n112 ) , .A1( u1_u11_u1_n169 ) , .A2( u1_u11_u1_n170 ) );
  AOI211_X1 u1_u11_u1_U5 (.ZN( u1_u11_u1_n124 ) , .A( u1_u11_u1_n138 ) , .C2( u1_u11_u1_n139 ) , .B( u1_u11_u1_n145 ) , .C1( u1_u11_u1_n147 ) );
  NAND2_X1 u1_u11_u1_U50 (.ZN( u1_u11_u1_n129 ) , .A2( u1_u11_u1_n95 ) , .A1( u1_u11_u1_n98 ) );
  NAND2_X1 u1_u11_u1_U51 (.A1( u1_u11_u1_n102 ) , .ZN( u1_u11_u1_n154 ) , .A2( u1_u11_u1_n99 ) );
  NAND2_X1 u1_u11_u1_U52 (.A2( u1_u11_u1_n100 ) , .ZN( u1_u11_u1_n135 ) , .A1( u1_u11_u1_n99 ) );
  AOI21_X1 u1_u11_u1_U53 (.A( u1_u11_u1_n152 ) , .B2( u1_u11_u1_n153 ) , .B1( u1_u11_u1_n154 ) , .ZN( u1_u11_u1_n158 ) );
  INV_X1 u1_u11_u1_U54 (.A( u1_u11_u1_n160 ) , .ZN( u1_u11_u1_n175 ) );
  NAND2_X1 u1_u11_u1_U55 (.A1( u1_u11_u1_n100 ) , .ZN( u1_u11_u1_n116 ) , .A2( u1_u11_u1_n95 ) );
  NAND2_X1 u1_u11_u1_U56 (.A1( u1_u11_u1_n102 ) , .ZN( u1_u11_u1_n131 ) , .A2( u1_u11_u1_n95 ) );
  NAND2_X1 u1_u11_u1_U57 (.A2( u1_u11_u1_n104 ) , .ZN( u1_u11_u1_n121 ) , .A1( u1_u11_u1_n98 ) );
  NAND2_X1 u1_u11_u1_U58 (.A1( u1_u11_u1_n103 ) , .ZN( u1_u11_u1_n153 ) , .A2( u1_u11_u1_n98 ) );
  NAND2_X1 u1_u11_u1_U59 (.A2( u1_u11_u1_n104 ) , .A1( u1_u11_u1_n105 ) , .ZN( u1_u11_u1_n133 ) );
  AOI22_X1 u1_u11_u1_U6 (.B2( u1_u11_u1_n113 ) , .A2( u1_u11_u1_n114 ) , .ZN( u1_u11_u1_n125 ) , .A1( u1_u11_u1_n171 ) , .B1( u1_u11_u1_n173 ) );
  NAND2_X1 u1_u11_u1_U60 (.ZN( u1_u11_u1_n150 ) , .A2( u1_u11_u1_n98 ) , .A1( u1_u11_u1_n99 ) );
  NAND2_X1 u1_u11_u1_U61 (.A1( u1_u11_u1_n105 ) , .ZN( u1_u11_u1_n155 ) , .A2( u1_u11_u1_n95 ) );
  OAI21_X1 u1_u11_u1_U62 (.ZN( u1_u11_u1_n109 ) , .B1( u1_u11_u1_n129 ) , .B2( u1_u11_u1_n160 ) , .A( u1_u11_u1_n167 ) );
  NAND2_X1 u1_u11_u1_U63 (.A2( u1_u11_u1_n100 ) , .A1( u1_u11_u1_n103 ) , .ZN( u1_u11_u1_n120 ) );
  NAND2_X1 u1_u11_u1_U64 (.A1( u1_u11_u1_n102 ) , .A2( u1_u11_u1_n104 ) , .ZN( u1_u11_u1_n115 ) );
  NAND2_X1 u1_u11_u1_U65 (.A2( u1_u11_u1_n100 ) , .A1( u1_u11_u1_n104 ) , .ZN( u1_u11_u1_n151 ) );
  NAND2_X1 u1_u11_u1_U66 (.A2( u1_u11_u1_n103 ) , .A1( u1_u11_u1_n105 ) , .ZN( u1_u11_u1_n161 ) );
  INV_X1 u1_u11_u1_U67 (.A( u1_u11_u1_n152 ) , .ZN( u1_u11_u1_n173 ) );
  INV_X1 u1_u11_u1_U68 (.A( u1_u11_u1_n128 ) , .ZN( u1_u11_u1_n172 ) );
  NAND2_X1 u1_u11_u1_U69 (.A2( u1_u11_u1_n102 ) , .A1( u1_u11_u1_n103 ) , .ZN( u1_u11_u1_n123 ) );
  NAND2_X1 u1_u11_u1_U7 (.ZN( u1_u11_u1_n114 ) , .A1( u1_u11_u1_n134 ) , .A2( u1_u11_u1_n156 ) );
  NOR2_X1 u1_u11_u1_U70 (.A2( u1_u11_X_7 ) , .A1( u1_u11_X_8 ) , .ZN( u1_u11_u1_n95 ) );
  NOR2_X1 u1_u11_u1_U71 (.A1( u1_u11_X_12 ) , .A2( u1_u11_X_9 ) , .ZN( u1_u11_u1_n100 ) );
  NOR2_X1 u1_u11_u1_U72 (.A2( u1_u11_X_8 ) , .A1( u1_u11_u1_n177 ) , .ZN( u1_u11_u1_n99 ) );
  NOR2_X1 u1_u11_u1_U73 (.A2( u1_u11_X_12 ) , .ZN( u1_u11_u1_n102 ) , .A1( u1_u11_u1_n176 ) );
  NOR2_X1 u1_u11_u1_U74 (.A2( u1_u11_X_9 ) , .ZN( u1_u11_u1_n105 ) , .A1( u1_u11_u1_n168 ) );
  NAND2_X1 u1_u11_u1_U75 (.A1( u1_u11_X_10 ) , .ZN( u1_u11_u1_n160 ) , .A2( u1_u11_u1_n169 ) );
  NAND2_X1 u1_u11_u1_U76 (.A2( u1_u11_X_10 ) , .A1( u1_u11_X_11 ) , .ZN( u1_u11_u1_n152 ) );
  NAND2_X1 u1_u11_u1_U77 (.A1( u1_u11_X_11 ) , .ZN( u1_u11_u1_n128 ) , .A2( u1_u11_u1_n170 ) );
  AND2_X1 u1_u11_u1_U78 (.A2( u1_u11_X_7 ) , .A1( u1_u11_X_8 ) , .ZN( u1_u11_u1_n104 ) );
  AND2_X1 u1_u11_u1_U79 (.A1( u1_u11_X_8 ) , .ZN( u1_u11_u1_n103 ) , .A2( u1_u11_u1_n177 ) );
  AOI22_X1 u1_u11_u1_U8 (.B2( u1_u11_u1_n136 ) , .A2( u1_u11_u1_n137 ) , .ZN( u1_u11_u1_n143 ) , .A1( u1_u11_u1_n171 ) , .B1( u1_u11_u1_n173 ) );
  INV_X1 u1_u11_u1_U80 (.A( u1_u11_X_10 ) , .ZN( u1_u11_u1_n170 ) );
  INV_X1 u1_u11_u1_U81 (.A( u1_u11_X_9 ) , .ZN( u1_u11_u1_n176 ) );
  INV_X1 u1_u11_u1_U82 (.A( u1_u11_X_11 ) , .ZN( u1_u11_u1_n169 ) );
  INV_X1 u1_u11_u1_U83 (.A( u1_u11_X_12 ) , .ZN( u1_u11_u1_n168 ) );
  INV_X1 u1_u11_u1_U84 (.A( u1_u11_X_7 ) , .ZN( u1_u11_u1_n177 ) );
  NAND4_X1 u1_u11_u1_U85 (.ZN( u1_out11_18 ) , .A4( u1_u11_u1_n165 ) , .A3( u1_u11_u1_n166 ) , .A1( u1_u11_u1_n167 ) , .A2( u1_u11_u1_n186 ) );
  AOI22_X1 u1_u11_u1_U86 (.B2( u1_u11_u1_n146 ) , .B1( u1_u11_u1_n147 ) , .A2( u1_u11_u1_n148 ) , .ZN( u1_u11_u1_n166 ) , .A1( u1_u11_u1_n172 ) );
  INV_X1 u1_u11_u1_U87 (.A( u1_u11_u1_n145 ) , .ZN( u1_u11_u1_n186 ) );
  NAND4_X1 u1_u11_u1_U88 (.ZN( u1_out11_2 ) , .A4( u1_u11_u1_n142 ) , .A3( u1_u11_u1_n143 ) , .A2( u1_u11_u1_n144 ) , .A1( u1_u11_u1_n179 ) );
  OAI21_X1 u1_u11_u1_U89 (.B2( u1_u11_u1_n132 ) , .ZN( u1_u11_u1_n144 ) , .A( u1_u11_u1_n146 ) , .B1( u1_u11_u1_n180 ) );
  INV_X1 u1_u11_u1_U9 (.A( u1_u11_u1_n147 ) , .ZN( u1_u11_u1_n181 ) );
  INV_X1 u1_u11_u1_U90 (.A( u1_u11_u1_n130 ) , .ZN( u1_u11_u1_n179 ) );
  NAND4_X1 u1_u11_u1_U91 (.ZN( u1_out11_28 ) , .A4( u1_u11_u1_n124 ) , .A3( u1_u11_u1_n125 ) , .A2( u1_u11_u1_n126 ) , .A1( u1_u11_u1_n127 ) );
  OAI21_X1 u1_u11_u1_U92 (.ZN( u1_u11_u1_n127 ) , .B2( u1_u11_u1_n139 ) , .B1( u1_u11_u1_n175 ) , .A( u1_u11_u1_n183 ) );
  OAI21_X1 u1_u11_u1_U93 (.ZN( u1_u11_u1_n126 ) , .B2( u1_u11_u1_n140 ) , .A( u1_u11_u1_n146 ) , .B1( u1_u11_u1_n178 ) );
  OR4_X1 u1_u11_u1_U94 (.ZN( u1_out11_13 ) , .A4( u1_u11_u1_n108 ) , .A3( u1_u11_u1_n109 ) , .A2( u1_u11_u1_n110 ) , .A1( u1_u11_u1_n111 ) );
  AOI21_X1 u1_u11_u1_U95 (.ZN( u1_u11_u1_n111 ) , .A( u1_u11_u1_n128 ) , .B2( u1_u11_u1_n131 ) , .B1( u1_u11_u1_n135 ) );
  AOI21_X1 u1_u11_u1_U96 (.ZN( u1_u11_u1_n110 ) , .A( u1_u11_u1_n116 ) , .B1( u1_u11_u1_n152 ) , .B2( u1_u11_u1_n160 ) );
  NAND3_X1 u1_u11_u1_U97 (.A3( u1_u11_u1_n149 ) , .A2( u1_u11_u1_n150 ) , .A1( u1_u11_u1_n151 ) , .ZN( u1_u11_u1_n164 ) );
  NAND3_X1 u1_u11_u1_U98 (.A3( u1_u11_u1_n134 ) , .A2( u1_u11_u1_n135 ) , .ZN( u1_u11_u1_n136 ) , .A1( u1_u11_u1_n151 ) );
  NAND3_X1 u1_u11_u1_U99 (.A1( u1_u11_u1_n133 ) , .ZN( u1_u11_u1_n137 ) , .A2( u1_u11_u1_n154 ) , .A3( u1_u11_u1_n181 ) );
  OAI22_X1 u1_u11_u2_U10 (.ZN( u1_u11_u2_n109 ) , .A2( u1_u11_u2_n113 ) , .B2( u1_u11_u2_n133 ) , .B1( u1_u11_u2_n167 ) , .A1( u1_u11_u2_n168 ) );
  NAND3_X1 u1_u11_u2_U100 (.A2( u1_u11_u2_n100 ) , .A1( u1_u11_u2_n104 ) , .A3( u1_u11_u2_n138 ) , .ZN( u1_u11_u2_n98 ) );
  OAI22_X1 u1_u11_u2_U11 (.B1( u1_u11_u2_n151 ) , .A2( u1_u11_u2_n152 ) , .A1( u1_u11_u2_n153 ) , .ZN( u1_u11_u2_n160 ) , .B2( u1_u11_u2_n168 ) );
  NOR3_X1 u1_u11_u2_U12 (.A1( u1_u11_u2_n150 ) , .ZN( u1_u11_u2_n151 ) , .A3( u1_u11_u2_n175 ) , .A2( u1_u11_u2_n188 ) );
  AOI21_X1 u1_u11_u2_U13 (.ZN( u1_u11_u2_n144 ) , .B2( u1_u11_u2_n155 ) , .A( u1_u11_u2_n172 ) , .B1( u1_u11_u2_n185 ) );
  AOI21_X1 u1_u11_u2_U14 (.B2( u1_u11_u2_n143 ) , .ZN( u1_u11_u2_n145 ) , .B1( u1_u11_u2_n152 ) , .A( u1_u11_u2_n171 ) );
  AOI21_X1 u1_u11_u2_U15 (.B2( u1_u11_u2_n120 ) , .B1( u1_u11_u2_n121 ) , .ZN( u1_u11_u2_n126 ) , .A( u1_u11_u2_n167 ) );
  INV_X1 u1_u11_u2_U16 (.A( u1_u11_u2_n156 ) , .ZN( u1_u11_u2_n171 ) );
  INV_X1 u1_u11_u2_U17 (.A( u1_u11_u2_n120 ) , .ZN( u1_u11_u2_n188 ) );
  NAND2_X1 u1_u11_u2_U18 (.A2( u1_u11_u2_n122 ) , .ZN( u1_u11_u2_n150 ) , .A1( u1_u11_u2_n152 ) );
  INV_X1 u1_u11_u2_U19 (.A( u1_u11_u2_n153 ) , .ZN( u1_u11_u2_n170 ) );
  INV_X1 u1_u11_u2_U20 (.A( u1_u11_u2_n137 ) , .ZN( u1_u11_u2_n173 ) );
  NAND2_X1 u1_u11_u2_U21 (.A1( u1_u11_u2_n132 ) , .A2( u1_u11_u2_n139 ) , .ZN( u1_u11_u2_n157 ) );
  INV_X1 u1_u11_u2_U22 (.A( u1_u11_u2_n113 ) , .ZN( u1_u11_u2_n178 ) );
  INV_X1 u1_u11_u2_U23 (.A( u1_u11_u2_n139 ) , .ZN( u1_u11_u2_n175 ) );
  INV_X1 u1_u11_u2_U24 (.A( u1_u11_u2_n155 ) , .ZN( u1_u11_u2_n181 ) );
  INV_X1 u1_u11_u2_U25 (.A( u1_u11_u2_n119 ) , .ZN( u1_u11_u2_n177 ) );
  INV_X1 u1_u11_u2_U26 (.A( u1_u11_u2_n116 ) , .ZN( u1_u11_u2_n180 ) );
  INV_X1 u1_u11_u2_U27 (.A( u1_u11_u2_n131 ) , .ZN( u1_u11_u2_n179 ) );
  INV_X1 u1_u11_u2_U28 (.A( u1_u11_u2_n154 ) , .ZN( u1_u11_u2_n176 ) );
  NAND2_X1 u1_u11_u2_U29 (.A2( u1_u11_u2_n116 ) , .A1( u1_u11_u2_n117 ) , .ZN( u1_u11_u2_n118 ) );
  NOR2_X1 u1_u11_u2_U3 (.ZN( u1_u11_u2_n121 ) , .A2( u1_u11_u2_n177 ) , .A1( u1_u11_u2_n180 ) );
  INV_X1 u1_u11_u2_U30 (.A( u1_u11_u2_n132 ) , .ZN( u1_u11_u2_n182 ) );
  INV_X1 u1_u11_u2_U31 (.A( u1_u11_u2_n158 ) , .ZN( u1_u11_u2_n183 ) );
  OAI21_X1 u1_u11_u2_U32 (.A( u1_u11_u2_n156 ) , .B1( u1_u11_u2_n157 ) , .ZN( u1_u11_u2_n158 ) , .B2( u1_u11_u2_n179 ) );
  NOR2_X1 u1_u11_u2_U33 (.ZN( u1_u11_u2_n156 ) , .A1( u1_u11_u2_n166 ) , .A2( u1_u11_u2_n169 ) );
  NOR2_X1 u1_u11_u2_U34 (.A2( u1_u11_u2_n114 ) , .ZN( u1_u11_u2_n137 ) , .A1( u1_u11_u2_n140 ) );
  NOR2_X1 u1_u11_u2_U35 (.A2( u1_u11_u2_n138 ) , .ZN( u1_u11_u2_n153 ) , .A1( u1_u11_u2_n156 ) );
  AOI211_X1 u1_u11_u2_U36 (.ZN( u1_u11_u2_n130 ) , .C1( u1_u11_u2_n138 ) , .C2( u1_u11_u2_n179 ) , .B( u1_u11_u2_n96 ) , .A( u1_u11_u2_n97 ) );
  OAI22_X1 u1_u11_u2_U37 (.B1( u1_u11_u2_n133 ) , .A2( u1_u11_u2_n137 ) , .A1( u1_u11_u2_n152 ) , .B2( u1_u11_u2_n168 ) , .ZN( u1_u11_u2_n97 ) );
  OAI221_X1 u1_u11_u2_U38 (.B1( u1_u11_u2_n113 ) , .C1( u1_u11_u2_n132 ) , .A( u1_u11_u2_n149 ) , .B2( u1_u11_u2_n171 ) , .C2( u1_u11_u2_n172 ) , .ZN( u1_u11_u2_n96 ) );
  OAI221_X1 u1_u11_u2_U39 (.A( u1_u11_u2_n115 ) , .C2( u1_u11_u2_n123 ) , .B2( u1_u11_u2_n143 ) , .B1( u1_u11_u2_n153 ) , .ZN( u1_u11_u2_n163 ) , .C1( u1_u11_u2_n168 ) );
  INV_X1 u1_u11_u2_U4 (.A( u1_u11_u2_n134 ) , .ZN( u1_u11_u2_n185 ) );
  OAI21_X1 u1_u11_u2_U40 (.A( u1_u11_u2_n114 ) , .ZN( u1_u11_u2_n115 ) , .B1( u1_u11_u2_n176 ) , .B2( u1_u11_u2_n178 ) );
  OAI221_X1 u1_u11_u2_U41 (.A( u1_u11_u2_n135 ) , .B2( u1_u11_u2_n136 ) , .B1( u1_u11_u2_n137 ) , .ZN( u1_u11_u2_n162 ) , .C2( u1_u11_u2_n167 ) , .C1( u1_u11_u2_n185 ) );
  AND3_X1 u1_u11_u2_U42 (.A3( u1_u11_u2_n131 ) , .A2( u1_u11_u2_n132 ) , .A1( u1_u11_u2_n133 ) , .ZN( u1_u11_u2_n136 ) );
  AOI22_X1 u1_u11_u2_U43 (.ZN( u1_u11_u2_n135 ) , .B1( u1_u11_u2_n140 ) , .A1( u1_u11_u2_n156 ) , .B2( u1_u11_u2_n180 ) , .A2( u1_u11_u2_n188 ) );
  AOI21_X1 u1_u11_u2_U44 (.ZN( u1_u11_u2_n149 ) , .B1( u1_u11_u2_n173 ) , .B2( u1_u11_u2_n188 ) , .A( u1_u11_u2_n95 ) );
  AND3_X1 u1_u11_u2_U45 (.A2( u1_u11_u2_n100 ) , .A1( u1_u11_u2_n104 ) , .A3( u1_u11_u2_n156 ) , .ZN( u1_u11_u2_n95 ) );
  OAI21_X1 u1_u11_u2_U46 (.A( u1_u11_u2_n101 ) , .B2( u1_u11_u2_n121 ) , .B1( u1_u11_u2_n153 ) , .ZN( u1_u11_u2_n164 ) );
  NAND2_X1 u1_u11_u2_U47 (.A2( u1_u11_u2_n100 ) , .A1( u1_u11_u2_n107 ) , .ZN( u1_u11_u2_n155 ) );
  NAND2_X1 u1_u11_u2_U48 (.A2( u1_u11_u2_n105 ) , .A1( u1_u11_u2_n108 ) , .ZN( u1_u11_u2_n143 ) );
  NAND2_X1 u1_u11_u2_U49 (.A1( u1_u11_u2_n104 ) , .A2( u1_u11_u2_n106 ) , .ZN( u1_u11_u2_n152 ) );
  INV_X1 u1_u11_u2_U5 (.A( u1_u11_u2_n150 ) , .ZN( u1_u11_u2_n184 ) );
  NAND2_X1 u1_u11_u2_U50 (.A1( u1_u11_u2_n100 ) , .A2( u1_u11_u2_n105 ) , .ZN( u1_u11_u2_n132 ) );
  INV_X1 u1_u11_u2_U51 (.A( u1_u11_u2_n140 ) , .ZN( u1_u11_u2_n168 ) );
  INV_X1 u1_u11_u2_U52 (.A( u1_u11_u2_n138 ) , .ZN( u1_u11_u2_n167 ) );
  OAI21_X1 u1_u11_u2_U53 (.A( u1_u11_u2_n141 ) , .B2( u1_u11_u2_n142 ) , .ZN( u1_u11_u2_n146 ) , .B1( u1_u11_u2_n153 ) );
  OAI21_X1 u1_u11_u2_U54 (.A( u1_u11_u2_n140 ) , .ZN( u1_u11_u2_n141 ) , .B1( u1_u11_u2_n176 ) , .B2( u1_u11_u2_n177 ) );
  NOR3_X1 u1_u11_u2_U55 (.ZN( u1_u11_u2_n142 ) , .A3( u1_u11_u2_n175 ) , .A2( u1_u11_u2_n178 ) , .A1( u1_u11_u2_n181 ) );
  INV_X1 u1_u11_u2_U56 (.ZN( u1_u11_u2_n187 ) , .A( u1_u11_u2_n99 ) );
  OAI21_X1 u1_u11_u2_U57 (.B1( u1_u11_u2_n137 ) , .B2( u1_u11_u2_n143 ) , .A( u1_u11_u2_n98 ) , .ZN( u1_u11_u2_n99 ) );
  NAND2_X1 u1_u11_u2_U58 (.A1( u1_u11_u2_n102 ) , .A2( u1_u11_u2_n106 ) , .ZN( u1_u11_u2_n113 ) );
  NAND2_X1 u1_u11_u2_U59 (.A1( u1_u11_u2_n106 ) , .A2( u1_u11_u2_n107 ) , .ZN( u1_u11_u2_n131 ) );
  NOR4_X1 u1_u11_u2_U6 (.A4( u1_u11_u2_n124 ) , .A3( u1_u11_u2_n125 ) , .A2( u1_u11_u2_n126 ) , .A1( u1_u11_u2_n127 ) , .ZN( u1_u11_u2_n128 ) );
  NAND2_X1 u1_u11_u2_U60 (.A1( u1_u11_u2_n103 ) , .A2( u1_u11_u2_n107 ) , .ZN( u1_u11_u2_n139 ) );
  NAND2_X1 u1_u11_u2_U61 (.A1( u1_u11_u2_n103 ) , .A2( u1_u11_u2_n105 ) , .ZN( u1_u11_u2_n133 ) );
  NAND2_X1 u1_u11_u2_U62 (.A1( u1_u11_u2_n102 ) , .A2( u1_u11_u2_n103 ) , .ZN( u1_u11_u2_n154 ) );
  NAND2_X1 u1_u11_u2_U63 (.A2( u1_u11_u2_n103 ) , .A1( u1_u11_u2_n104 ) , .ZN( u1_u11_u2_n119 ) );
  NAND2_X1 u1_u11_u2_U64 (.A2( u1_u11_u2_n107 ) , .A1( u1_u11_u2_n108 ) , .ZN( u1_u11_u2_n123 ) );
  NAND2_X1 u1_u11_u2_U65 (.A1( u1_u11_u2_n104 ) , .A2( u1_u11_u2_n108 ) , .ZN( u1_u11_u2_n122 ) );
  INV_X1 u1_u11_u2_U66 (.A( u1_u11_u2_n114 ) , .ZN( u1_u11_u2_n172 ) );
  NAND2_X1 u1_u11_u2_U67 (.A2( u1_u11_u2_n100 ) , .A1( u1_u11_u2_n102 ) , .ZN( u1_u11_u2_n116 ) );
  NAND2_X1 u1_u11_u2_U68 (.A1( u1_u11_u2_n102 ) , .A2( u1_u11_u2_n108 ) , .ZN( u1_u11_u2_n120 ) );
  NAND2_X1 u1_u11_u2_U69 (.A2( u1_u11_u2_n105 ) , .A1( u1_u11_u2_n106 ) , .ZN( u1_u11_u2_n117 ) );
  AOI21_X1 u1_u11_u2_U7 (.ZN( u1_u11_u2_n124 ) , .B1( u1_u11_u2_n131 ) , .B2( u1_u11_u2_n143 ) , .A( u1_u11_u2_n172 ) );
  NOR2_X1 u1_u11_u2_U70 (.A2( u1_u11_X_16 ) , .ZN( u1_u11_u2_n140 ) , .A1( u1_u11_u2_n166 ) );
  NOR2_X1 u1_u11_u2_U71 (.A2( u1_u11_X_13 ) , .A1( u1_u11_X_14 ) , .ZN( u1_u11_u2_n100 ) );
  NOR2_X1 u1_u11_u2_U72 (.A2( u1_u11_X_16 ) , .A1( u1_u11_X_17 ) , .ZN( u1_u11_u2_n138 ) );
  NOR2_X1 u1_u11_u2_U73 (.A2( u1_u11_X_15 ) , .A1( u1_u11_X_18 ) , .ZN( u1_u11_u2_n104 ) );
  NOR2_X1 u1_u11_u2_U74 (.A2( u1_u11_X_14 ) , .ZN( u1_u11_u2_n103 ) , .A1( u1_u11_u2_n174 ) );
  NOR2_X1 u1_u11_u2_U75 (.A2( u1_u11_X_15 ) , .ZN( u1_u11_u2_n102 ) , .A1( u1_u11_u2_n165 ) );
  NOR2_X1 u1_u11_u2_U76 (.A2( u1_u11_X_17 ) , .ZN( u1_u11_u2_n114 ) , .A1( u1_u11_u2_n169 ) );
  AND2_X1 u1_u11_u2_U77 (.A1( u1_u11_X_15 ) , .ZN( u1_u11_u2_n105 ) , .A2( u1_u11_u2_n165 ) );
  AND2_X1 u1_u11_u2_U78 (.A2( u1_u11_X_15 ) , .A1( u1_u11_X_18 ) , .ZN( u1_u11_u2_n107 ) );
  AND2_X1 u1_u11_u2_U79 (.A1( u1_u11_X_14 ) , .ZN( u1_u11_u2_n106 ) , .A2( u1_u11_u2_n174 ) );
  AOI21_X1 u1_u11_u2_U8 (.B2( u1_u11_u2_n119 ) , .ZN( u1_u11_u2_n127 ) , .A( u1_u11_u2_n137 ) , .B1( u1_u11_u2_n155 ) );
  AND2_X1 u1_u11_u2_U80 (.A1( u1_u11_X_13 ) , .A2( u1_u11_X_14 ) , .ZN( u1_u11_u2_n108 ) );
  INV_X1 u1_u11_u2_U81 (.A( u1_u11_X_16 ) , .ZN( u1_u11_u2_n169 ) );
  INV_X1 u1_u11_u2_U82 (.A( u1_u11_X_17 ) , .ZN( u1_u11_u2_n166 ) );
  INV_X1 u1_u11_u2_U83 (.A( u1_u11_X_13 ) , .ZN( u1_u11_u2_n174 ) );
  INV_X1 u1_u11_u2_U84 (.A( u1_u11_X_18 ) , .ZN( u1_u11_u2_n165 ) );
  NAND4_X1 u1_u11_u2_U85 (.ZN( u1_out11_30 ) , .A4( u1_u11_u2_n147 ) , .A3( u1_u11_u2_n148 ) , .A2( u1_u11_u2_n149 ) , .A1( u1_u11_u2_n187 ) );
  NOR3_X1 u1_u11_u2_U86 (.A3( u1_u11_u2_n144 ) , .A2( u1_u11_u2_n145 ) , .A1( u1_u11_u2_n146 ) , .ZN( u1_u11_u2_n147 ) );
  AOI21_X1 u1_u11_u2_U87 (.B2( u1_u11_u2_n138 ) , .ZN( u1_u11_u2_n148 ) , .A( u1_u11_u2_n162 ) , .B1( u1_u11_u2_n182 ) );
  NAND4_X1 u1_u11_u2_U88 (.ZN( u1_out11_24 ) , .A4( u1_u11_u2_n111 ) , .A3( u1_u11_u2_n112 ) , .A1( u1_u11_u2_n130 ) , .A2( u1_u11_u2_n187 ) );
  AOI221_X1 u1_u11_u2_U89 (.A( u1_u11_u2_n109 ) , .B1( u1_u11_u2_n110 ) , .ZN( u1_u11_u2_n111 ) , .C1( u1_u11_u2_n134 ) , .C2( u1_u11_u2_n170 ) , .B2( u1_u11_u2_n173 ) );
  AOI21_X1 u1_u11_u2_U9 (.B2( u1_u11_u2_n123 ) , .ZN( u1_u11_u2_n125 ) , .A( u1_u11_u2_n171 ) , .B1( u1_u11_u2_n184 ) );
  AOI21_X1 u1_u11_u2_U90 (.ZN( u1_u11_u2_n112 ) , .B2( u1_u11_u2_n156 ) , .A( u1_u11_u2_n164 ) , .B1( u1_u11_u2_n181 ) );
  NAND4_X1 u1_u11_u2_U91 (.ZN( u1_out11_16 ) , .A4( u1_u11_u2_n128 ) , .A3( u1_u11_u2_n129 ) , .A1( u1_u11_u2_n130 ) , .A2( u1_u11_u2_n186 ) );
  AOI22_X1 u1_u11_u2_U92 (.A2( u1_u11_u2_n118 ) , .ZN( u1_u11_u2_n129 ) , .A1( u1_u11_u2_n140 ) , .B1( u1_u11_u2_n157 ) , .B2( u1_u11_u2_n170 ) );
  INV_X1 u1_u11_u2_U93 (.A( u1_u11_u2_n163 ) , .ZN( u1_u11_u2_n186 ) );
  OR4_X1 u1_u11_u2_U94 (.ZN( u1_out11_6 ) , .A4( u1_u11_u2_n161 ) , .A3( u1_u11_u2_n162 ) , .A2( u1_u11_u2_n163 ) , .A1( u1_u11_u2_n164 ) );
  OR3_X1 u1_u11_u2_U95 (.A2( u1_u11_u2_n159 ) , .A1( u1_u11_u2_n160 ) , .ZN( u1_u11_u2_n161 ) , .A3( u1_u11_u2_n183 ) );
  AOI21_X1 u1_u11_u2_U96 (.B2( u1_u11_u2_n154 ) , .B1( u1_u11_u2_n155 ) , .ZN( u1_u11_u2_n159 ) , .A( u1_u11_u2_n167 ) );
  NAND3_X1 u1_u11_u2_U97 (.A2( u1_u11_u2_n117 ) , .A1( u1_u11_u2_n122 ) , .A3( u1_u11_u2_n123 ) , .ZN( u1_u11_u2_n134 ) );
  NAND3_X1 u1_u11_u2_U98 (.ZN( u1_u11_u2_n110 ) , .A2( u1_u11_u2_n131 ) , .A3( u1_u11_u2_n139 ) , .A1( u1_u11_u2_n154 ) );
  NAND3_X1 u1_u11_u2_U99 (.A2( u1_u11_u2_n100 ) , .ZN( u1_u11_u2_n101 ) , .A1( u1_u11_u2_n104 ) , .A3( u1_u11_u2_n114 ) );
  XOR2_X1 u1_u12_U10 (.B( u1_K13_45 ) , .A( u1_R11_30 ) , .Z( u1_u12_X_45 ) );
  XOR2_X1 u1_u12_U16 (.B( u1_K13_3 ) , .A( u1_R11_2 ) , .Z( u1_u12_X_3 ) );
  XOR2_X1 u1_u12_U29 (.B( u1_K13_28 ) , .A( u1_R11_19 ) , .Z( u1_u12_X_28 ) );
  XOR2_X1 u1_u12_U30 (.B( u1_K13_27 ) , .A( u1_R11_18 ) , .Z( u1_u12_X_27 ) );
  XOR2_X1 u1_u12_U31 (.B( u1_K13_26 ) , .A( u1_R11_17 ) , .Z( u1_u12_X_26 ) );
  XOR2_X1 u1_u12_U33 (.B( u1_K13_24 ) , .A( u1_R11_17 ) , .Z( u1_u12_X_24 ) );
  XOR2_X1 u1_u12_U35 (.B( u1_K13_22 ) , .A( u1_R11_15 ) , .Z( u1_u12_X_22 ) );
  XOR2_X1 u1_u12_U36 (.B( u1_K13_21 ) , .A( u1_R11_14 ) , .Z( u1_u12_X_21 ) );
  XOR2_X1 u1_u12_U38 (.B( u1_K13_1 ) , .A( u1_R11_32 ) , .Z( u1_u12_X_1 ) );
  XOR2_X1 u1_u12_U4 (.B( u1_K13_6 ) , .A( u1_R11_5 ) , .Z( u1_u12_X_6 ) );
  XOR2_X1 u1_u12_U6 (.B( u1_K13_4 ) , .A( u1_R11_3 ) , .Z( u1_u12_X_4 ) );
  XOR2_X1 u1_u12_U8 (.B( u1_K13_47 ) , .A( u1_R11_32 ) , .Z( u1_u12_X_47 ) );
  XOR2_X1 u1_u12_U9 (.B( u1_K13_46 ) , .A( u1_R11_31 ) , .Z( u1_u12_X_46 ) );
  NAND2_X1 u1_u12_u0_U10 (.ZN( u1_u12_u0_n113 ) , .A1( u1_u12_u0_n139 ) , .A2( u1_u12_u0_n149 ) );
  AND3_X1 u1_u12_u0_U11 (.A2( u1_u12_u0_n112 ) , .ZN( u1_u12_u0_n127 ) , .A3( u1_u12_u0_n130 ) , .A1( u1_u12_u0_n148 ) );
  AND2_X1 u1_u12_u0_U12 (.ZN( u1_u12_u0_n107 ) , .A1( u1_u12_u0_n130 ) , .A2( u1_u12_u0_n140 ) );
  AND2_X1 u1_u12_u0_U13 (.A2( u1_u12_u0_n129 ) , .A1( u1_u12_u0_n130 ) , .ZN( u1_u12_u0_n151 ) );
  AND2_X1 u1_u12_u0_U14 (.A1( u1_u12_u0_n108 ) , .A2( u1_u12_u0_n125 ) , .ZN( u1_u12_u0_n145 ) );
  INV_X1 u1_u12_u0_U15 (.A( u1_u12_u0_n143 ) , .ZN( u1_u12_u0_n173 ) );
  NOR2_X1 u1_u12_u0_U16 (.A2( u1_u12_u0_n136 ) , .ZN( u1_u12_u0_n147 ) , .A1( u1_u12_u0_n160 ) );
  AOI21_X1 u1_u12_u0_U17 (.B1( u1_u12_u0_n103 ) , .ZN( u1_u12_u0_n132 ) , .A( u1_u12_u0_n165 ) , .B2( u1_u12_u0_n93 ) );
  INV_X1 u1_u12_u0_U18 (.A( u1_u12_u0_n142 ) , .ZN( u1_u12_u0_n165 ) );
  OAI22_X1 u1_u12_u0_U19 (.B1( u1_u12_u0_n131 ) , .A1( u1_u12_u0_n144 ) , .B2( u1_u12_u0_n147 ) , .A2( u1_u12_u0_n90 ) , .ZN( u1_u12_u0_n91 ) );
  AND3_X1 u1_u12_u0_U20 (.A3( u1_u12_u0_n121 ) , .A2( u1_u12_u0_n125 ) , .A1( u1_u12_u0_n148 ) , .ZN( u1_u12_u0_n90 ) );
  OAI22_X1 u1_u12_u0_U21 (.B1( u1_u12_u0_n125 ) , .ZN( u1_u12_u0_n126 ) , .A1( u1_u12_u0_n138 ) , .A2( u1_u12_u0_n146 ) , .B2( u1_u12_u0_n147 ) );
  INV_X1 u1_u12_u0_U22 (.A( u1_u12_u0_n136 ) , .ZN( u1_u12_u0_n161 ) );
  AOI22_X1 u1_u12_u0_U23 (.B2( u1_u12_u0_n109 ) , .A2( u1_u12_u0_n110 ) , .ZN( u1_u12_u0_n111 ) , .B1( u1_u12_u0_n118 ) , .A1( u1_u12_u0_n160 ) );
  NAND2_X1 u1_u12_u0_U24 (.A2( u1_u12_u0_n103 ) , .ZN( u1_u12_u0_n140 ) , .A1( u1_u12_u0_n94 ) );
  NAND2_X1 u1_u12_u0_U25 (.A2( u1_u12_u0_n102 ) , .A1( u1_u12_u0_n103 ) , .ZN( u1_u12_u0_n149 ) );
  INV_X1 u1_u12_u0_U26 (.A( u1_u12_u0_n118 ) , .ZN( u1_u12_u0_n158 ) );
  NAND2_X1 u1_u12_u0_U27 (.A2( u1_u12_u0_n100 ) , .ZN( u1_u12_u0_n131 ) , .A1( u1_u12_u0_n92 ) );
  NAND2_X1 u1_u12_u0_U28 (.ZN( u1_u12_u0_n108 ) , .A1( u1_u12_u0_n92 ) , .A2( u1_u12_u0_n94 ) );
  AOI21_X1 u1_u12_u0_U29 (.ZN( u1_u12_u0_n104 ) , .B1( u1_u12_u0_n107 ) , .B2( u1_u12_u0_n141 ) , .A( u1_u12_u0_n144 ) );
  INV_X1 u1_u12_u0_U3 (.A( u1_u12_u0_n113 ) , .ZN( u1_u12_u0_n166 ) );
  AOI21_X1 u1_u12_u0_U30 (.ZN( u1_u12_u0_n116 ) , .B2( u1_u12_u0_n142 ) , .A( u1_u12_u0_n144 ) , .B1( u1_u12_u0_n166 ) );
  AOI21_X1 u1_u12_u0_U31 (.B1( u1_u12_u0_n127 ) , .B2( u1_u12_u0_n129 ) , .A( u1_u12_u0_n138 ) , .ZN( u1_u12_u0_n96 ) );
  NAND2_X1 u1_u12_u0_U32 (.A2( u1_u12_u0_n102 ) , .ZN( u1_u12_u0_n114 ) , .A1( u1_u12_u0_n92 ) );
  NOR2_X1 u1_u12_u0_U33 (.A1( u1_u12_u0_n120 ) , .ZN( u1_u12_u0_n143 ) , .A2( u1_u12_u0_n167 ) );
  OAI221_X1 u1_u12_u0_U34 (.C1( u1_u12_u0_n112 ) , .ZN( u1_u12_u0_n120 ) , .B1( u1_u12_u0_n138 ) , .B2( u1_u12_u0_n141 ) , .C2( u1_u12_u0_n147 ) , .A( u1_u12_u0_n172 ) );
  AOI211_X1 u1_u12_u0_U35 (.B( u1_u12_u0_n115 ) , .A( u1_u12_u0_n116 ) , .C2( u1_u12_u0_n117 ) , .C1( u1_u12_u0_n118 ) , .ZN( u1_u12_u0_n119 ) );
  NAND2_X1 u1_u12_u0_U36 (.A1( u1_u12_u0_n100 ) , .A2( u1_u12_u0_n103 ) , .ZN( u1_u12_u0_n125 ) );
  NAND2_X1 u1_u12_u0_U37 (.A1( u1_u12_u0_n101 ) , .A2( u1_u12_u0_n102 ) , .ZN( u1_u12_u0_n150 ) );
  INV_X1 u1_u12_u0_U38 (.A( u1_u12_u0_n138 ) , .ZN( u1_u12_u0_n160 ) );
  NAND2_X1 u1_u12_u0_U39 (.A2( u1_u12_u0_n100 ) , .A1( u1_u12_u0_n101 ) , .ZN( u1_u12_u0_n139 ) );
  AOI21_X1 u1_u12_u0_U4 (.B1( u1_u12_u0_n114 ) , .ZN( u1_u12_u0_n115 ) , .B2( u1_u12_u0_n129 ) , .A( u1_u12_u0_n161 ) );
  NAND2_X1 u1_u12_u0_U40 (.A1( u1_u12_u0_n101 ) , .ZN( u1_u12_u0_n130 ) , .A2( u1_u12_u0_n94 ) );
  NAND2_X1 u1_u12_u0_U41 (.ZN( u1_u12_u0_n112 ) , .A2( u1_u12_u0_n92 ) , .A1( u1_u12_u0_n93 ) );
  INV_X1 u1_u12_u0_U42 (.ZN( u1_u12_u0_n172 ) , .A( u1_u12_u0_n88 ) );
  OAI222_X1 u1_u12_u0_U43 (.C1( u1_u12_u0_n108 ) , .A1( u1_u12_u0_n125 ) , .B2( u1_u12_u0_n128 ) , .B1( u1_u12_u0_n144 ) , .A2( u1_u12_u0_n158 ) , .C2( u1_u12_u0_n161 ) , .ZN( u1_u12_u0_n88 ) );
  NAND2_X1 u1_u12_u0_U44 (.A2( u1_u12_u0_n101 ) , .ZN( u1_u12_u0_n121 ) , .A1( u1_u12_u0_n93 ) );
  OR3_X1 u1_u12_u0_U45 (.A3( u1_u12_u0_n152 ) , .A2( u1_u12_u0_n153 ) , .A1( u1_u12_u0_n154 ) , .ZN( u1_u12_u0_n155 ) );
  AOI21_X1 u1_u12_u0_U46 (.B2( u1_u12_u0_n150 ) , .B1( u1_u12_u0_n151 ) , .ZN( u1_u12_u0_n152 ) , .A( u1_u12_u0_n158 ) );
  AOI21_X1 u1_u12_u0_U47 (.A( u1_u12_u0_n144 ) , .B2( u1_u12_u0_n145 ) , .B1( u1_u12_u0_n146 ) , .ZN( u1_u12_u0_n154 ) );
  AOI21_X1 u1_u12_u0_U48 (.A( u1_u12_u0_n147 ) , .B2( u1_u12_u0_n148 ) , .B1( u1_u12_u0_n149 ) , .ZN( u1_u12_u0_n153 ) );
  INV_X1 u1_u12_u0_U49 (.ZN( u1_u12_u0_n171 ) , .A( u1_u12_u0_n99 ) );
  AOI21_X1 u1_u12_u0_U5 (.B2( u1_u12_u0_n131 ) , .ZN( u1_u12_u0_n134 ) , .B1( u1_u12_u0_n151 ) , .A( u1_u12_u0_n158 ) );
  OAI211_X1 u1_u12_u0_U50 (.C2( u1_u12_u0_n140 ) , .C1( u1_u12_u0_n161 ) , .A( u1_u12_u0_n169 ) , .B( u1_u12_u0_n98 ) , .ZN( u1_u12_u0_n99 ) );
  INV_X1 u1_u12_u0_U51 (.ZN( u1_u12_u0_n169 ) , .A( u1_u12_u0_n91 ) );
  AOI211_X1 u1_u12_u0_U52 (.C1( u1_u12_u0_n118 ) , .A( u1_u12_u0_n123 ) , .B( u1_u12_u0_n96 ) , .C2( u1_u12_u0_n97 ) , .ZN( u1_u12_u0_n98 ) );
  NOR2_X1 u1_u12_u0_U53 (.A2( u1_u12_X_4 ) , .A1( u1_u12_X_5 ) , .ZN( u1_u12_u0_n118 ) );
  NOR2_X1 u1_u12_u0_U54 (.A2( u1_u12_X_1 ) , .ZN( u1_u12_u0_n101 ) , .A1( u1_u12_u0_n163 ) );
  NOR2_X1 u1_u12_u0_U55 (.A2( u1_u12_X_6 ) , .ZN( u1_u12_u0_n100 ) , .A1( u1_u12_u0_n162 ) );
  NAND2_X1 u1_u12_u0_U56 (.A2( u1_u12_X_4 ) , .A1( u1_u12_X_5 ) , .ZN( u1_u12_u0_n144 ) );
  NOR2_X1 u1_u12_u0_U57 (.A2( u1_u12_X_5 ) , .ZN( u1_u12_u0_n136 ) , .A1( u1_u12_u0_n159 ) );
  NAND2_X1 u1_u12_u0_U58 (.A1( u1_u12_X_5 ) , .ZN( u1_u12_u0_n138 ) , .A2( u1_u12_u0_n159 ) );
  AND2_X1 u1_u12_u0_U59 (.A2( u1_u12_X_3 ) , .A1( u1_u12_X_6 ) , .ZN( u1_u12_u0_n102 ) );
  NOR2_X1 u1_u12_u0_U6 (.A1( u1_u12_u0_n108 ) , .ZN( u1_u12_u0_n123 ) , .A2( u1_u12_u0_n158 ) );
  AND2_X1 u1_u12_u0_U60 (.A1( u1_u12_X_6 ) , .A2( u1_u12_u0_n162 ) , .ZN( u1_u12_u0_n93 ) );
  INV_X1 u1_u12_u0_U61 (.A( u1_u12_X_4 ) , .ZN( u1_u12_u0_n159 ) );
  INV_X1 u1_u12_u0_U62 (.A( u1_u12_X_1 ) , .ZN( u1_u12_u0_n164 ) );
  INV_X1 u1_u12_u0_U63 (.A( u1_u12_X_3 ) , .ZN( u1_u12_u0_n162 ) );
  OR4_X1 u1_u12_u0_U64 (.ZN( u1_out12_17 ) , .A4( u1_u12_u0_n122 ) , .A2( u1_u12_u0_n123 ) , .A1( u1_u12_u0_n124 ) , .A3( u1_u12_u0_n170 ) );
  AOI21_X1 u1_u12_u0_U65 (.B2( u1_u12_u0_n107 ) , .ZN( u1_u12_u0_n124 ) , .B1( u1_u12_u0_n128 ) , .A( u1_u12_u0_n161 ) );
  INV_X1 u1_u12_u0_U66 (.A( u1_u12_u0_n111 ) , .ZN( u1_u12_u0_n170 ) );
  OR4_X1 u1_u12_u0_U67 (.ZN( u1_out12_31 ) , .A4( u1_u12_u0_n155 ) , .A2( u1_u12_u0_n156 ) , .A1( u1_u12_u0_n157 ) , .A3( u1_u12_u0_n173 ) );
  AOI21_X1 u1_u12_u0_U68 (.A( u1_u12_u0_n138 ) , .B2( u1_u12_u0_n139 ) , .B1( u1_u12_u0_n140 ) , .ZN( u1_u12_u0_n157 ) );
  AOI21_X1 u1_u12_u0_U69 (.B2( u1_u12_u0_n141 ) , .B1( u1_u12_u0_n142 ) , .ZN( u1_u12_u0_n156 ) , .A( u1_u12_u0_n161 ) );
  OAI21_X1 u1_u12_u0_U7 (.B1( u1_u12_u0_n150 ) , .B2( u1_u12_u0_n158 ) , .A( u1_u12_u0_n172 ) , .ZN( u1_u12_u0_n89 ) );
  INV_X1 u1_u12_u0_U70 (.ZN( u1_u12_u0_n174 ) , .A( u1_u12_u0_n89 ) );
  AOI211_X1 u1_u12_u0_U71 (.B( u1_u12_u0_n104 ) , .A( u1_u12_u0_n105 ) , .ZN( u1_u12_u0_n106 ) , .C2( u1_u12_u0_n113 ) , .C1( u1_u12_u0_n160 ) );
  INV_X1 u1_u12_u0_U72 (.A( u1_u12_u0_n126 ) , .ZN( u1_u12_u0_n168 ) );
  AOI211_X1 u1_u12_u0_U73 (.B( u1_u12_u0_n133 ) , .A( u1_u12_u0_n134 ) , .C2( u1_u12_u0_n135 ) , .C1( u1_u12_u0_n136 ) , .ZN( u1_u12_u0_n137 ) );
  NOR2_X1 u1_u12_u0_U74 (.A1( u1_u12_u0_n163 ) , .A2( u1_u12_u0_n164 ) , .ZN( u1_u12_u0_n95 ) );
  NOR2_X1 u1_u12_u0_U75 (.A2( u1_u12_X_3 ) , .A1( u1_u12_X_6 ) , .ZN( u1_u12_u0_n94 ) );
  OAI221_X1 u1_u12_u0_U76 (.C1( u1_u12_u0_n121 ) , .ZN( u1_u12_u0_n122 ) , .B2( u1_u12_u0_n127 ) , .A( u1_u12_u0_n143 ) , .B1( u1_u12_u0_n144 ) , .C2( u1_u12_u0_n147 ) );
  AOI21_X1 u1_u12_u0_U77 (.B1( u1_u12_u0_n132 ) , .ZN( u1_u12_u0_n133 ) , .A( u1_u12_u0_n144 ) , .B2( u1_u12_u0_n166 ) );
  OAI22_X1 u1_u12_u0_U78 (.ZN( u1_u12_u0_n105 ) , .A2( u1_u12_u0_n132 ) , .B1( u1_u12_u0_n146 ) , .A1( u1_u12_u0_n147 ) , .B2( u1_u12_u0_n161 ) );
  NAND2_X1 u1_u12_u0_U79 (.ZN( u1_u12_u0_n110 ) , .A2( u1_u12_u0_n132 ) , .A1( u1_u12_u0_n145 ) );
  AND2_X1 u1_u12_u0_U8 (.A1( u1_u12_u0_n114 ) , .A2( u1_u12_u0_n121 ) , .ZN( u1_u12_u0_n146 ) );
  INV_X1 u1_u12_u0_U80 (.A( u1_u12_u0_n119 ) , .ZN( u1_u12_u0_n167 ) );
  NAND2_X1 u1_u12_u0_U81 (.ZN( u1_u12_u0_n148 ) , .A1( u1_u12_u0_n93 ) , .A2( u1_u12_u0_n95 ) );
  NAND2_X1 u1_u12_u0_U82 (.A1( u1_u12_u0_n100 ) , .ZN( u1_u12_u0_n129 ) , .A2( u1_u12_u0_n95 ) );
  NAND2_X1 u1_u12_u0_U83 (.A1( u1_u12_u0_n102 ) , .ZN( u1_u12_u0_n128 ) , .A2( u1_u12_u0_n95 ) );
  NOR2_X1 u1_u12_u0_U84 (.A2( u1_u12_X_1 ) , .A1( u1_u12_X_2 ) , .ZN( u1_u12_u0_n92 ) );
  NAND2_X1 u1_u12_u0_U85 (.ZN( u1_u12_u0_n142 ) , .A1( u1_u12_u0_n94 ) , .A2( u1_u12_u0_n95 ) );
  NOR2_X1 u1_u12_u0_U86 (.A2( u1_u12_X_2 ) , .ZN( u1_u12_u0_n103 ) , .A1( u1_u12_u0_n164 ) );
  INV_X1 u1_u12_u0_U87 (.A( u1_u12_X_2 ) , .ZN( u1_u12_u0_n163 ) );
  NAND3_X1 u1_u12_u0_U88 (.ZN( u1_out12_23 ) , .A3( u1_u12_u0_n137 ) , .A1( u1_u12_u0_n168 ) , .A2( u1_u12_u0_n171 ) );
  NAND3_X1 u1_u12_u0_U89 (.A3( u1_u12_u0_n127 ) , .A2( u1_u12_u0_n128 ) , .ZN( u1_u12_u0_n135 ) , .A1( u1_u12_u0_n150 ) );
  AND2_X1 u1_u12_u0_U9 (.A1( u1_u12_u0_n131 ) , .ZN( u1_u12_u0_n141 ) , .A2( u1_u12_u0_n150 ) );
  NAND3_X1 u1_u12_u0_U90 (.ZN( u1_u12_u0_n117 ) , .A3( u1_u12_u0_n132 ) , .A2( u1_u12_u0_n139 ) , .A1( u1_u12_u0_n148 ) );
  NAND3_X1 u1_u12_u0_U91 (.ZN( u1_u12_u0_n109 ) , .A2( u1_u12_u0_n114 ) , .A3( u1_u12_u0_n140 ) , .A1( u1_u12_u0_n149 ) );
  NAND3_X1 u1_u12_u0_U92 (.ZN( u1_out12_9 ) , .A3( u1_u12_u0_n106 ) , .A2( u1_u12_u0_n171 ) , .A1( u1_u12_u0_n174 ) );
  NAND3_X1 u1_u12_u0_U93 (.A2( u1_u12_u0_n128 ) , .A1( u1_u12_u0_n132 ) , .A3( u1_u12_u0_n146 ) , .ZN( u1_u12_u0_n97 ) );
  OAI22_X1 u1_u12_u3_U10 (.B1( u1_u12_u3_n113 ) , .A2( u1_u12_u3_n135 ) , .A1( u1_u12_u3_n150 ) , .B2( u1_u12_u3_n164 ) , .ZN( u1_u12_u3_n98 ) );
  OAI211_X1 u1_u12_u3_U11 (.B( u1_u12_u3_n106 ) , .ZN( u1_u12_u3_n119 ) , .C2( u1_u12_u3_n128 ) , .C1( u1_u12_u3_n167 ) , .A( u1_u12_u3_n181 ) );
  AOI221_X1 u1_u12_u3_U12 (.C1( u1_u12_u3_n105 ) , .ZN( u1_u12_u3_n106 ) , .A( u1_u12_u3_n131 ) , .B2( u1_u12_u3_n132 ) , .C2( u1_u12_u3_n133 ) , .B1( u1_u12_u3_n169 ) );
  INV_X1 u1_u12_u3_U13 (.ZN( u1_u12_u3_n181 ) , .A( u1_u12_u3_n98 ) );
  NAND2_X1 u1_u12_u3_U14 (.ZN( u1_u12_u3_n105 ) , .A2( u1_u12_u3_n130 ) , .A1( u1_u12_u3_n155 ) );
  AOI22_X1 u1_u12_u3_U15 (.B1( u1_u12_u3_n115 ) , .A2( u1_u12_u3_n116 ) , .ZN( u1_u12_u3_n123 ) , .B2( u1_u12_u3_n133 ) , .A1( u1_u12_u3_n169 ) );
  NAND2_X1 u1_u12_u3_U16 (.ZN( u1_u12_u3_n116 ) , .A2( u1_u12_u3_n151 ) , .A1( u1_u12_u3_n182 ) );
  NOR2_X1 u1_u12_u3_U17 (.ZN( u1_u12_u3_n126 ) , .A2( u1_u12_u3_n150 ) , .A1( u1_u12_u3_n164 ) );
  AOI21_X1 u1_u12_u3_U18 (.ZN( u1_u12_u3_n112 ) , .B2( u1_u12_u3_n146 ) , .B1( u1_u12_u3_n155 ) , .A( u1_u12_u3_n167 ) );
  NAND2_X1 u1_u12_u3_U19 (.A1( u1_u12_u3_n135 ) , .ZN( u1_u12_u3_n142 ) , .A2( u1_u12_u3_n164 ) );
  NAND2_X1 u1_u12_u3_U20 (.ZN( u1_u12_u3_n132 ) , .A2( u1_u12_u3_n152 ) , .A1( u1_u12_u3_n156 ) );
  AND2_X1 u1_u12_u3_U21 (.A2( u1_u12_u3_n113 ) , .A1( u1_u12_u3_n114 ) , .ZN( u1_u12_u3_n151 ) );
  INV_X1 u1_u12_u3_U22 (.A( u1_u12_u3_n133 ) , .ZN( u1_u12_u3_n165 ) );
  INV_X1 u1_u12_u3_U23 (.A( u1_u12_u3_n135 ) , .ZN( u1_u12_u3_n170 ) );
  NAND2_X1 u1_u12_u3_U24 (.A1( u1_u12_u3_n107 ) , .A2( u1_u12_u3_n108 ) , .ZN( u1_u12_u3_n140 ) );
  NAND2_X1 u1_u12_u3_U25 (.ZN( u1_u12_u3_n117 ) , .A1( u1_u12_u3_n124 ) , .A2( u1_u12_u3_n148 ) );
  NAND2_X1 u1_u12_u3_U26 (.ZN( u1_u12_u3_n143 ) , .A1( u1_u12_u3_n165 ) , .A2( u1_u12_u3_n167 ) );
  INV_X1 u1_u12_u3_U27 (.A( u1_u12_u3_n130 ) , .ZN( u1_u12_u3_n177 ) );
  INV_X1 u1_u12_u3_U28 (.A( u1_u12_u3_n128 ) , .ZN( u1_u12_u3_n176 ) );
  INV_X1 u1_u12_u3_U29 (.A( u1_u12_u3_n155 ) , .ZN( u1_u12_u3_n174 ) );
  INV_X1 u1_u12_u3_U3 (.A( u1_u12_u3_n129 ) , .ZN( u1_u12_u3_n183 ) );
  INV_X1 u1_u12_u3_U30 (.A( u1_u12_u3_n139 ) , .ZN( u1_u12_u3_n185 ) );
  NOR2_X1 u1_u12_u3_U31 (.ZN( u1_u12_u3_n135 ) , .A2( u1_u12_u3_n141 ) , .A1( u1_u12_u3_n169 ) );
  OAI222_X1 u1_u12_u3_U32 (.C2( u1_u12_u3_n107 ) , .A2( u1_u12_u3_n108 ) , .B1( u1_u12_u3_n135 ) , .ZN( u1_u12_u3_n138 ) , .B2( u1_u12_u3_n146 ) , .C1( u1_u12_u3_n154 ) , .A1( u1_u12_u3_n164 ) );
  NOR4_X1 u1_u12_u3_U33 (.A4( u1_u12_u3_n157 ) , .A3( u1_u12_u3_n158 ) , .A2( u1_u12_u3_n159 ) , .A1( u1_u12_u3_n160 ) , .ZN( u1_u12_u3_n161 ) );
  AOI21_X1 u1_u12_u3_U34 (.B2( u1_u12_u3_n152 ) , .B1( u1_u12_u3_n153 ) , .ZN( u1_u12_u3_n158 ) , .A( u1_u12_u3_n164 ) );
  AOI21_X1 u1_u12_u3_U35 (.A( u1_u12_u3_n154 ) , .B2( u1_u12_u3_n155 ) , .B1( u1_u12_u3_n156 ) , .ZN( u1_u12_u3_n157 ) );
  AOI21_X1 u1_u12_u3_U36 (.A( u1_u12_u3_n149 ) , .B2( u1_u12_u3_n150 ) , .B1( u1_u12_u3_n151 ) , .ZN( u1_u12_u3_n159 ) );
  AOI211_X1 u1_u12_u3_U37 (.ZN( u1_u12_u3_n109 ) , .A( u1_u12_u3_n119 ) , .C2( u1_u12_u3_n129 ) , .B( u1_u12_u3_n138 ) , .C1( u1_u12_u3_n141 ) );
  AOI211_X1 u1_u12_u3_U38 (.B( u1_u12_u3_n119 ) , .A( u1_u12_u3_n120 ) , .C2( u1_u12_u3_n121 ) , .ZN( u1_u12_u3_n122 ) , .C1( u1_u12_u3_n179 ) );
  INV_X1 u1_u12_u3_U39 (.A( u1_u12_u3_n156 ) , .ZN( u1_u12_u3_n179 ) );
  INV_X1 u1_u12_u3_U4 (.A( u1_u12_u3_n140 ) , .ZN( u1_u12_u3_n182 ) );
  OAI22_X1 u1_u12_u3_U40 (.B1( u1_u12_u3_n118 ) , .ZN( u1_u12_u3_n120 ) , .A1( u1_u12_u3_n135 ) , .B2( u1_u12_u3_n154 ) , .A2( u1_u12_u3_n178 ) );
  AND3_X1 u1_u12_u3_U41 (.ZN( u1_u12_u3_n118 ) , .A2( u1_u12_u3_n124 ) , .A1( u1_u12_u3_n144 ) , .A3( u1_u12_u3_n152 ) );
  INV_X1 u1_u12_u3_U42 (.A( u1_u12_u3_n121 ) , .ZN( u1_u12_u3_n164 ) );
  NAND2_X1 u1_u12_u3_U43 (.ZN( u1_u12_u3_n133 ) , .A1( u1_u12_u3_n154 ) , .A2( u1_u12_u3_n164 ) );
  OAI211_X1 u1_u12_u3_U44 (.B( u1_u12_u3_n127 ) , .ZN( u1_u12_u3_n139 ) , .C1( u1_u12_u3_n150 ) , .C2( u1_u12_u3_n154 ) , .A( u1_u12_u3_n184 ) );
  INV_X1 u1_u12_u3_U45 (.A( u1_u12_u3_n125 ) , .ZN( u1_u12_u3_n184 ) );
  AOI221_X1 u1_u12_u3_U46 (.A( u1_u12_u3_n126 ) , .ZN( u1_u12_u3_n127 ) , .C2( u1_u12_u3_n132 ) , .C1( u1_u12_u3_n169 ) , .B2( u1_u12_u3_n170 ) , .B1( u1_u12_u3_n174 ) );
  OAI22_X1 u1_u12_u3_U47 (.A1( u1_u12_u3_n124 ) , .ZN( u1_u12_u3_n125 ) , .B2( u1_u12_u3_n145 ) , .A2( u1_u12_u3_n165 ) , .B1( u1_u12_u3_n167 ) );
  NOR2_X1 u1_u12_u3_U48 (.A1( u1_u12_u3_n113 ) , .ZN( u1_u12_u3_n131 ) , .A2( u1_u12_u3_n154 ) );
  NAND2_X1 u1_u12_u3_U49 (.A1( u1_u12_u3_n103 ) , .ZN( u1_u12_u3_n150 ) , .A2( u1_u12_u3_n99 ) );
  INV_X1 u1_u12_u3_U5 (.A( u1_u12_u3_n117 ) , .ZN( u1_u12_u3_n178 ) );
  NAND2_X1 u1_u12_u3_U50 (.A2( u1_u12_u3_n102 ) , .ZN( u1_u12_u3_n155 ) , .A1( u1_u12_u3_n97 ) );
  INV_X1 u1_u12_u3_U51 (.A( u1_u12_u3_n141 ) , .ZN( u1_u12_u3_n167 ) );
  AOI21_X1 u1_u12_u3_U52 (.B2( u1_u12_u3_n114 ) , .B1( u1_u12_u3_n146 ) , .A( u1_u12_u3_n154 ) , .ZN( u1_u12_u3_n94 ) );
  AOI21_X1 u1_u12_u3_U53 (.ZN( u1_u12_u3_n110 ) , .B2( u1_u12_u3_n142 ) , .B1( u1_u12_u3_n186 ) , .A( u1_u12_u3_n95 ) );
  INV_X1 u1_u12_u3_U54 (.A( u1_u12_u3_n145 ) , .ZN( u1_u12_u3_n186 ) );
  AOI21_X1 u1_u12_u3_U55 (.B1( u1_u12_u3_n124 ) , .A( u1_u12_u3_n149 ) , .B2( u1_u12_u3_n155 ) , .ZN( u1_u12_u3_n95 ) );
  INV_X1 u1_u12_u3_U56 (.A( u1_u12_u3_n149 ) , .ZN( u1_u12_u3_n169 ) );
  NAND2_X1 u1_u12_u3_U57 (.ZN( u1_u12_u3_n124 ) , .A1( u1_u12_u3_n96 ) , .A2( u1_u12_u3_n97 ) );
  NAND2_X1 u1_u12_u3_U58 (.A2( u1_u12_u3_n100 ) , .ZN( u1_u12_u3_n146 ) , .A1( u1_u12_u3_n96 ) );
  NAND2_X1 u1_u12_u3_U59 (.A1( u1_u12_u3_n101 ) , .ZN( u1_u12_u3_n145 ) , .A2( u1_u12_u3_n99 ) );
  AOI221_X1 u1_u12_u3_U6 (.A( u1_u12_u3_n131 ) , .C2( u1_u12_u3_n132 ) , .C1( u1_u12_u3_n133 ) , .ZN( u1_u12_u3_n134 ) , .B1( u1_u12_u3_n143 ) , .B2( u1_u12_u3_n177 ) );
  NAND2_X1 u1_u12_u3_U60 (.A1( u1_u12_u3_n100 ) , .ZN( u1_u12_u3_n156 ) , .A2( u1_u12_u3_n99 ) );
  NAND2_X1 u1_u12_u3_U61 (.A2( u1_u12_u3_n101 ) , .A1( u1_u12_u3_n104 ) , .ZN( u1_u12_u3_n148 ) );
  NAND2_X1 u1_u12_u3_U62 (.A1( u1_u12_u3_n100 ) , .A2( u1_u12_u3_n102 ) , .ZN( u1_u12_u3_n128 ) );
  NAND2_X1 u1_u12_u3_U63 (.A2( u1_u12_u3_n101 ) , .A1( u1_u12_u3_n102 ) , .ZN( u1_u12_u3_n152 ) );
  NAND2_X1 u1_u12_u3_U64 (.A2( u1_u12_u3_n101 ) , .ZN( u1_u12_u3_n114 ) , .A1( u1_u12_u3_n96 ) );
  NAND2_X1 u1_u12_u3_U65 (.ZN( u1_u12_u3_n107 ) , .A1( u1_u12_u3_n97 ) , .A2( u1_u12_u3_n99 ) );
  NAND2_X1 u1_u12_u3_U66 (.A2( u1_u12_u3_n100 ) , .A1( u1_u12_u3_n104 ) , .ZN( u1_u12_u3_n113 ) );
  NAND2_X1 u1_u12_u3_U67 (.A1( u1_u12_u3_n104 ) , .ZN( u1_u12_u3_n153 ) , .A2( u1_u12_u3_n97 ) );
  NAND2_X1 u1_u12_u3_U68 (.A2( u1_u12_u3_n103 ) , .A1( u1_u12_u3_n104 ) , .ZN( u1_u12_u3_n130 ) );
  NAND2_X1 u1_u12_u3_U69 (.A2( u1_u12_u3_n103 ) , .ZN( u1_u12_u3_n144 ) , .A1( u1_u12_u3_n96 ) );
  OAI22_X1 u1_u12_u3_U7 (.B2( u1_u12_u3_n147 ) , .A2( u1_u12_u3_n148 ) , .ZN( u1_u12_u3_n160 ) , .B1( u1_u12_u3_n165 ) , .A1( u1_u12_u3_n168 ) );
  NAND2_X1 u1_u12_u3_U70 (.A1( u1_u12_u3_n102 ) , .A2( u1_u12_u3_n103 ) , .ZN( u1_u12_u3_n108 ) );
  NOR2_X1 u1_u12_u3_U71 (.A2( u1_u12_X_19 ) , .A1( u1_u12_X_20 ) , .ZN( u1_u12_u3_n99 ) );
  NOR2_X1 u1_u12_u3_U72 (.A2( u1_u12_X_21 ) , .A1( u1_u12_X_24 ) , .ZN( u1_u12_u3_n103 ) );
  NOR2_X1 u1_u12_u3_U73 (.A2( u1_u12_X_24 ) , .A1( u1_u12_u3_n171 ) , .ZN( u1_u12_u3_n97 ) );
  NOR2_X1 u1_u12_u3_U74 (.A2( u1_u12_X_23 ) , .ZN( u1_u12_u3_n141 ) , .A1( u1_u12_u3_n166 ) );
  NOR2_X1 u1_u12_u3_U75 (.A2( u1_u12_X_19 ) , .A1( u1_u12_u3_n172 ) , .ZN( u1_u12_u3_n96 ) );
  NAND2_X1 u1_u12_u3_U76 (.A1( u1_u12_X_22 ) , .A2( u1_u12_X_23 ) , .ZN( u1_u12_u3_n154 ) );
  NAND2_X1 u1_u12_u3_U77 (.A1( u1_u12_X_23 ) , .ZN( u1_u12_u3_n149 ) , .A2( u1_u12_u3_n166 ) );
  NOR2_X1 u1_u12_u3_U78 (.A2( u1_u12_X_22 ) , .A1( u1_u12_X_23 ) , .ZN( u1_u12_u3_n121 ) );
  AND2_X1 u1_u12_u3_U79 (.A1( u1_u12_X_24 ) , .ZN( u1_u12_u3_n101 ) , .A2( u1_u12_u3_n171 ) );
  AND3_X1 u1_u12_u3_U8 (.A3( u1_u12_u3_n144 ) , .A2( u1_u12_u3_n145 ) , .A1( u1_u12_u3_n146 ) , .ZN( u1_u12_u3_n147 ) );
  AND2_X1 u1_u12_u3_U80 (.A1( u1_u12_X_19 ) , .ZN( u1_u12_u3_n102 ) , .A2( u1_u12_u3_n172 ) );
  AND2_X1 u1_u12_u3_U81 (.A1( u1_u12_X_21 ) , .A2( u1_u12_X_24 ) , .ZN( u1_u12_u3_n100 ) );
  AND2_X1 u1_u12_u3_U82 (.A2( u1_u12_X_19 ) , .A1( u1_u12_X_20 ) , .ZN( u1_u12_u3_n104 ) );
  INV_X1 u1_u12_u3_U83 (.A( u1_u12_X_22 ) , .ZN( u1_u12_u3_n166 ) );
  INV_X1 u1_u12_u3_U84 (.A( u1_u12_X_21 ) , .ZN( u1_u12_u3_n171 ) );
  INV_X1 u1_u12_u3_U85 (.A( u1_u12_X_20 ) , .ZN( u1_u12_u3_n172 ) );
  NAND4_X1 u1_u12_u3_U86 (.ZN( u1_out12_26 ) , .A4( u1_u12_u3_n109 ) , .A3( u1_u12_u3_n110 ) , .A2( u1_u12_u3_n111 ) , .A1( u1_u12_u3_n173 ) );
  INV_X1 u1_u12_u3_U87 (.ZN( u1_u12_u3_n173 ) , .A( u1_u12_u3_n94 ) );
  OAI21_X1 u1_u12_u3_U88 (.ZN( u1_u12_u3_n111 ) , .B2( u1_u12_u3_n117 ) , .A( u1_u12_u3_n133 ) , .B1( u1_u12_u3_n176 ) );
  NAND4_X1 u1_u12_u3_U89 (.ZN( u1_out12_20 ) , .A4( u1_u12_u3_n122 ) , .A3( u1_u12_u3_n123 ) , .A1( u1_u12_u3_n175 ) , .A2( u1_u12_u3_n180 ) );
  INV_X1 u1_u12_u3_U9 (.A( u1_u12_u3_n143 ) , .ZN( u1_u12_u3_n168 ) );
  INV_X1 u1_u12_u3_U90 (.A( u1_u12_u3_n126 ) , .ZN( u1_u12_u3_n180 ) );
  INV_X1 u1_u12_u3_U91 (.A( u1_u12_u3_n112 ) , .ZN( u1_u12_u3_n175 ) );
  NAND4_X1 u1_u12_u3_U92 (.ZN( u1_out12_1 ) , .A4( u1_u12_u3_n161 ) , .A3( u1_u12_u3_n162 ) , .A2( u1_u12_u3_n163 ) , .A1( u1_u12_u3_n185 ) );
  NAND2_X1 u1_u12_u3_U93 (.ZN( u1_u12_u3_n163 ) , .A2( u1_u12_u3_n170 ) , .A1( u1_u12_u3_n176 ) );
  AOI22_X1 u1_u12_u3_U94 (.B2( u1_u12_u3_n140 ) , .B1( u1_u12_u3_n141 ) , .A2( u1_u12_u3_n142 ) , .ZN( u1_u12_u3_n162 ) , .A1( u1_u12_u3_n177 ) );
  OR4_X1 u1_u12_u3_U95 (.ZN( u1_out12_10 ) , .A4( u1_u12_u3_n136 ) , .A3( u1_u12_u3_n137 ) , .A1( u1_u12_u3_n138 ) , .A2( u1_u12_u3_n139 ) );
  OAI222_X1 u1_u12_u3_U96 (.C1( u1_u12_u3_n128 ) , .ZN( u1_u12_u3_n137 ) , .B1( u1_u12_u3_n148 ) , .A2( u1_u12_u3_n150 ) , .B2( u1_u12_u3_n154 ) , .C2( u1_u12_u3_n164 ) , .A1( u1_u12_u3_n167 ) );
  OAI221_X1 u1_u12_u3_U97 (.A( u1_u12_u3_n134 ) , .B2( u1_u12_u3_n135 ) , .ZN( u1_u12_u3_n136 ) , .C1( u1_u12_u3_n149 ) , .B1( u1_u12_u3_n151 ) , .C2( u1_u12_u3_n183 ) );
  NAND3_X1 u1_u12_u3_U98 (.A1( u1_u12_u3_n114 ) , .ZN( u1_u12_u3_n115 ) , .A2( u1_u12_u3_n145 ) , .A3( u1_u12_u3_n153 ) );
  NAND3_X1 u1_u12_u3_U99 (.ZN( u1_u12_u3_n129 ) , .A2( u1_u12_u3_n144 ) , .A1( u1_u12_u3_n153 ) , .A3( u1_u12_u3_n182 ) );
  OAI22_X1 u1_u12_u4_U10 (.B2( u1_u12_u4_n135 ) , .ZN( u1_u12_u4_n137 ) , .B1( u1_u12_u4_n153 ) , .A1( u1_u12_u4_n155 ) , .A2( u1_u12_u4_n171 ) );
  AND3_X1 u1_u12_u4_U11 (.A2( u1_u12_u4_n134 ) , .ZN( u1_u12_u4_n135 ) , .A3( u1_u12_u4_n145 ) , .A1( u1_u12_u4_n157 ) );
  NAND2_X1 u1_u12_u4_U12 (.ZN( u1_u12_u4_n132 ) , .A2( u1_u12_u4_n170 ) , .A1( u1_u12_u4_n173 ) );
  AOI21_X1 u1_u12_u4_U13 (.B2( u1_u12_u4_n160 ) , .B1( u1_u12_u4_n161 ) , .ZN( u1_u12_u4_n162 ) , .A( u1_u12_u4_n170 ) );
  AOI21_X1 u1_u12_u4_U14 (.ZN( u1_u12_u4_n107 ) , .B2( u1_u12_u4_n143 ) , .A( u1_u12_u4_n174 ) , .B1( u1_u12_u4_n184 ) );
  AOI21_X1 u1_u12_u4_U15 (.B2( u1_u12_u4_n158 ) , .B1( u1_u12_u4_n159 ) , .ZN( u1_u12_u4_n163 ) , .A( u1_u12_u4_n174 ) );
  AOI21_X1 u1_u12_u4_U16 (.A( u1_u12_u4_n153 ) , .B2( u1_u12_u4_n154 ) , .B1( u1_u12_u4_n155 ) , .ZN( u1_u12_u4_n165 ) );
  AOI21_X1 u1_u12_u4_U17 (.A( u1_u12_u4_n156 ) , .B2( u1_u12_u4_n157 ) , .ZN( u1_u12_u4_n164 ) , .B1( u1_u12_u4_n184 ) );
  INV_X1 u1_u12_u4_U18 (.A( u1_u12_u4_n138 ) , .ZN( u1_u12_u4_n170 ) );
  AND2_X1 u1_u12_u4_U19 (.A2( u1_u12_u4_n120 ) , .ZN( u1_u12_u4_n155 ) , .A1( u1_u12_u4_n160 ) );
  INV_X1 u1_u12_u4_U20 (.A( u1_u12_u4_n156 ) , .ZN( u1_u12_u4_n175 ) );
  NAND2_X1 u1_u12_u4_U21 (.A2( u1_u12_u4_n118 ) , .ZN( u1_u12_u4_n131 ) , .A1( u1_u12_u4_n147 ) );
  NAND2_X1 u1_u12_u4_U22 (.A1( u1_u12_u4_n119 ) , .A2( u1_u12_u4_n120 ) , .ZN( u1_u12_u4_n130 ) );
  NAND2_X1 u1_u12_u4_U23 (.ZN( u1_u12_u4_n117 ) , .A2( u1_u12_u4_n118 ) , .A1( u1_u12_u4_n148 ) );
  NAND2_X1 u1_u12_u4_U24 (.ZN( u1_u12_u4_n129 ) , .A1( u1_u12_u4_n134 ) , .A2( u1_u12_u4_n148 ) );
  AND3_X1 u1_u12_u4_U25 (.A1( u1_u12_u4_n119 ) , .A2( u1_u12_u4_n143 ) , .A3( u1_u12_u4_n154 ) , .ZN( u1_u12_u4_n161 ) );
  AND2_X1 u1_u12_u4_U26 (.A1( u1_u12_u4_n145 ) , .A2( u1_u12_u4_n147 ) , .ZN( u1_u12_u4_n159 ) );
  OR3_X1 u1_u12_u4_U27 (.A3( u1_u12_u4_n114 ) , .A2( u1_u12_u4_n115 ) , .A1( u1_u12_u4_n116 ) , .ZN( u1_u12_u4_n136 ) );
  AOI21_X1 u1_u12_u4_U28 (.A( u1_u12_u4_n113 ) , .ZN( u1_u12_u4_n116 ) , .B2( u1_u12_u4_n173 ) , .B1( u1_u12_u4_n174 ) );
  AOI21_X1 u1_u12_u4_U29 (.ZN( u1_u12_u4_n115 ) , .B2( u1_u12_u4_n145 ) , .B1( u1_u12_u4_n146 ) , .A( u1_u12_u4_n156 ) );
  NOR2_X1 u1_u12_u4_U3 (.ZN( u1_u12_u4_n121 ) , .A1( u1_u12_u4_n181 ) , .A2( u1_u12_u4_n182 ) );
  OAI22_X1 u1_u12_u4_U30 (.ZN( u1_u12_u4_n114 ) , .A2( u1_u12_u4_n121 ) , .B1( u1_u12_u4_n160 ) , .B2( u1_u12_u4_n170 ) , .A1( u1_u12_u4_n171 ) );
  INV_X1 u1_u12_u4_U31 (.A( u1_u12_u4_n158 ) , .ZN( u1_u12_u4_n182 ) );
  INV_X1 u1_u12_u4_U32 (.ZN( u1_u12_u4_n181 ) , .A( u1_u12_u4_n96 ) );
  INV_X1 u1_u12_u4_U33 (.A( u1_u12_u4_n144 ) , .ZN( u1_u12_u4_n179 ) );
  INV_X1 u1_u12_u4_U34 (.A( u1_u12_u4_n157 ) , .ZN( u1_u12_u4_n178 ) );
  NAND2_X1 u1_u12_u4_U35 (.A2( u1_u12_u4_n154 ) , .A1( u1_u12_u4_n96 ) , .ZN( u1_u12_u4_n97 ) );
  INV_X1 u1_u12_u4_U36 (.ZN( u1_u12_u4_n186 ) , .A( u1_u12_u4_n95 ) );
  OAI221_X1 u1_u12_u4_U37 (.C1( u1_u12_u4_n134 ) , .B1( u1_u12_u4_n158 ) , .B2( u1_u12_u4_n171 ) , .C2( u1_u12_u4_n173 ) , .A( u1_u12_u4_n94 ) , .ZN( u1_u12_u4_n95 ) );
  AOI222_X1 u1_u12_u4_U38 (.B2( u1_u12_u4_n132 ) , .A1( u1_u12_u4_n138 ) , .C2( u1_u12_u4_n175 ) , .A2( u1_u12_u4_n179 ) , .C1( u1_u12_u4_n181 ) , .B1( u1_u12_u4_n185 ) , .ZN( u1_u12_u4_n94 ) );
  INV_X1 u1_u12_u4_U39 (.A( u1_u12_u4_n113 ) , .ZN( u1_u12_u4_n185 ) );
  INV_X1 u1_u12_u4_U4 (.A( u1_u12_u4_n117 ) , .ZN( u1_u12_u4_n184 ) );
  INV_X1 u1_u12_u4_U40 (.A( u1_u12_u4_n143 ) , .ZN( u1_u12_u4_n183 ) );
  NOR2_X1 u1_u12_u4_U41 (.ZN( u1_u12_u4_n138 ) , .A1( u1_u12_u4_n168 ) , .A2( u1_u12_u4_n169 ) );
  NOR2_X1 u1_u12_u4_U42 (.A1( u1_u12_u4_n150 ) , .A2( u1_u12_u4_n152 ) , .ZN( u1_u12_u4_n153 ) );
  NOR2_X1 u1_u12_u4_U43 (.A2( u1_u12_u4_n128 ) , .A1( u1_u12_u4_n138 ) , .ZN( u1_u12_u4_n156 ) );
  AOI22_X1 u1_u12_u4_U44 (.B2( u1_u12_u4_n122 ) , .A1( u1_u12_u4_n123 ) , .ZN( u1_u12_u4_n124 ) , .B1( u1_u12_u4_n128 ) , .A2( u1_u12_u4_n172 ) );
  INV_X1 u1_u12_u4_U45 (.A( u1_u12_u4_n153 ) , .ZN( u1_u12_u4_n172 ) );
  NAND2_X1 u1_u12_u4_U46 (.A2( u1_u12_u4_n120 ) , .ZN( u1_u12_u4_n123 ) , .A1( u1_u12_u4_n161 ) );
  AOI22_X1 u1_u12_u4_U47 (.B2( u1_u12_u4_n132 ) , .A2( u1_u12_u4_n133 ) , .ZN( u1_u12_u4_n140 ) , .A1( u1_u12_u4_n150 ) , .B1( u1_u12_u4_n179 ) );
  NAND2_X1 u1_u12_u4_U48 (.ZN( u1_u12_u4_n133 ) , .A2( u1_u12_u4_n146 ) , .A1( u1_u12_u4_n154 ) );
  NAND2_X1 u1_u12_u4_U49 (.A1( u1_u12_u4_n103 ) , .ZN( u1_u12_u4_n154 ) , .A2( u1_u12_u4_n98 ) );
  NOR4_X1 u1_u12_u4_U5 (.A4( u1_u12_u4_n106 ) , .A3( u1_u12_u4_n107 ) , .A2( u1_u12_u4_n108 ) , .A1( u1_u12_u4_n109 ) , .ZN( u1_u12_u4_n110 ) );
  NAND2_X1 u1_u12_u4_U50 (.A1( u1_u12_u4_n101 ) , .ZN( u1_u12_u4_n158 ) , .A2( u1_u12_u4_n99 ) );
  AOI21_X1 u1_u12_u4_U51 (.ZN( u1_u12_u4_n127 ) , .A( u1_u12_u4_n136 ) , .B2( u1_u12_u4_n150 ) , .B1( u1_u12_u4_n180 ) );
  INV_X1 u1_u12_u4_U52 (.A( u1_u12_u4_n160 ) , .ZN( u1_u12_u4_n180 ) );
  NAND2_X1 u1_u12_u4_U53 (.A2( u1_u12_u4_n104 ) , .A1( u1_u12_u4_n105 ) , .ZN( u1_u12_u4_n146 ) );
  NAND2_X1 u1_u12_u4_U54 (.A2( u1_u12_u4_n101 ) , .A1( u1_u12_u4_n102 ) , .ZN( u1_u12_u4_n160 ) );
  NAND2_X1 u1_u12_u4_U55 (.ZN( u1_u12_u4_n134 ) , .A1( u1_u12_u4_n98 ) , .A2( u1_u12_u4_n99 ) );
  NAND2_X1 u1_u12_u4_U56 (.A1( u1_u12_u4_n103 ) , .A2( u1_u12_u4_n104 ) , .ZN( u1_u12_u4_n143 ) );
  NAND2_X1 u1_u12_u4_U57 (.A2( u1_u12_u4_n105 ) , .ZN( u1_u12_u4_n145 ) , .A1( u1_u12_u4_n98 ) );
  NAND2_X1 u1_u12_u4_U58 (.A1( u1_u12_u4_n100 ) , .A2( u1_u12_u4_n105 ) , .ZN( u1_u12_u4_n120 ) );
  NAND2_X1 u1_u12_u4_U59 (.A1( u1_u12_u4_n102 ) , .A2( u1_u12_u4_n104 ) , .ZN( u1_u12_u4_n148 ) );
  AOI21_X1 u1_u12_u4_U6 (.ZN( u1_u12_u4_n106 ) , .B2( u1_u12_u4_n146 ) , .B1( u1_u12_u4_n158 ) , .A( u1_u12_u4_n170 ) );
  NAND2_X1 u1_u12_u4_U60 (.A2( u1_u12_u4_n100 ) , .A1( u1_u12_u4_n103 ) , .ZN( u1_u12_u4_n157 ) );
  INV_X1 u1_u12_u4_U61 (.A( u1_u12_u4_n150 ) , .ZN( u1_u12_u4_n173 ) );
  INV_X1 u1_u12_u4_U62 (.A( u1_u12_u4_n152 ) , .ZN( u1_u12_u4_n171 ) );
  NAND2_X1 u1_u12_u4_U63 (.A1( u1_u12_u4_n100 ) , .ZN( u1_u12_u4_n118 ) , .A2( u1_u12_u4_n99 ) );
  NAND2_X1 u1_u12_u4_U64 (.A2( u1_u12_u4_n100 ) , .A1( u1_u12_u4_n102 ) , .ZN( u1_u12_u4_n144 ) );
  NAND2_X1 u1_u12_u4_U65 (.A2( u1_u12_u4_n101 ) , .A1( u1_u12_u4_n105 ) , .ZN( u1_u12_u4_n96 ) );
  INV_X1 u1_u12_u4_U66 (.A( u1_u12_u4_n128 ) , .ZN( u1_u12_u4_n174 ) );
  NAND2_X1 u1_u12_u4_U67 (.A2( u1_u12_u4_n102 ) , .ZN( u1_u12_u4_n119 ) , .A1( u1_u12_u4_n98 ) );
  NAND2_X1 u1_u12_u4_U68 (.A2( u1_u12_u4_n101 ) , .A1( u1_u12_u4_n103 ) , .ZN( u1_u12_u4_n147 ) );
  NAND2_X1 u1_u12_u4_U69 (.A2( u1_u12_u4_n104 ) , .ZN( u1_u12_u4_n113 ) , .A1( u1_u12_u4_n99 ) );
  AOI21_X1 u1_u12_u4_U7 (.ZN( u1_u12_u4_n108 ) , .B2( u1_u12_u4_n134 ) , .B1( u1_u12_u4_n155 ) , .A( u1_u12_u4_n156 ) );
  NOR2_X1 u1_u12_u4_U70 (.A2( u1_u12_X_28 ) , .ZN( u1_u12_u4_n150 ) , .A1( u1_u12_u4_n168 ) );
  NOR2_X1 u1_u12_u4_U71 (.A2( u1_u12_X_29 ) , .ZN( u1_u12_u4_n152 ) , .A1( u1_u12_u4_n169 ) );
  NOR2_X1 u1_u12_u4_U72 (.A2( u1_u12_X_30 ) , .ZN( u1_u12_u4_n105 ) , .A1( u1_u12_u4_n176 ) );
  NOR2_X1 u1_u12_u4_U73 (.A2( u1_u12_X_26 ) , .ZN( u1_u12_u4_n100 ) , .A1( u1_u12_u4_n177 ) );
  NOR2_X1 u1_u12_u4_U74 (.A2( u1_u12_X_28 ) , .A1( u1_u12_X_29 ) , .ZN( u1_u12_u4_n128 ) );
  NOR2_X1 u1_u12_u4_U75 (.A2( u1_u12_X_27 ) , .A1( u1_u12_X_30 ) , .ZN( u1_u12_u4_n102 ) );
  NOR2_X1 u1_u12_u4_U76 (.A2( u1_u12_X_25 ) , .A1( u1_u12_X_26 ) , .ZN( u1_u12_u4_n98 ) );
  AND2_X1 u1_u12_u4_U77 (.A2( u1_u12_X_25 ) , .A1( u1_u12_X_26 ) , .ZN( u1_u12_u4_n104 ) );
  AND2_X1 u1_u12_u4_U78 (.A1( u1_u12_X_30 ) , .A2( u1_u12_u4_n176 ) , .ZN( u1_u12_u4_n99 ) );
  AND2_X1 u1_u12_u4_U79 (.A1( u1_u12_X_26 ) , .ZN( u1_u12_u4_n101 ) , .A2( u1_u12_u4_n177 ) );
  AOI21_X1 u1_u12_u4_U8 (.ZN( u1_u12_u4_n109 ) , .A( u1_u12_u4_n153 ) , .B1( u1_u12_u4_n159 ) , .B2( u1_u12_u4_n184 ) );
  AND2_X1 u1_u12_u4_U80 (.A1( u1_u12_X_27 ) , .A2( u1_u12_X_30 ) , .ZN( u1_u12_u4_n103 ) );
  INV_X1 u1_u12_u4_U81 (.A( u1_u12_X_28 ) , .ZN( u1_u12_u4_n169 ) );
  INV_X1 u1_u12_u4_U82 (.A( u1_u12_X_29 ) , .ZN( u1_u12_u4_n168 ) );
  INV_X1 u1_u12_u4_U83 (.A( u1_u12_X_25 ) , .ZN( u1_u12_u4_n177 ) );
  INV_X1 u1_u12_u4_U84 (.A( u1_u12_X_27 ) , .ZN( u1_u12_u4_n176 ) );
  NAND4_X1 u1_u12_u4_U85 (.ZN( u1_out12_25 ) , .A4( u1_u12_u4_n139 ) , .A3( u1_u12_u4_n140 ) , .A2( u1_u12_u4_n141 ) , .A1( u1_u12_u4_n142 ) );
  OAI21_X1 u1_u12_u4_U86 (.A( u1_u12_u4_n128 ) , .B2( u1_u12_u4_n129 ) , .B1( u1_u12_u4_n130 ) , .ZN( u1_u12_u4_n142 ) );
  OAI21_X1 u1_u12_u4_U87 (.B2( u1_u12_u4_n131 ) , .ZN( u1_u12_u4_n141 ) , .A( u1_u12_u4_n175 ) , .B1( u1_u12_u4_n183 ) );
  NAND4_X1 u1_u12_u4_U88 (.ZN( u1_out12_14 ) , .A4( u1_u12_u4_n124 ) , .A3( u1_u12_u4_n125 ) , .A2( u1_u12_u4_n126 ) , .A1( u1_u12_u4_n127 ) );
  AOI22_X1 u1_u12_u4_U89 (.B2( u1_u12_u4_n117 ) , .ZN( u1_u12_u4_n126 ) , .A1( u1_u12_u4_n129 ) , .B1( u1_u12_u4_n152 ) , .A2( u1_u12_u4_n175 ) );
  AOI211_X1 u1_u12_u4_U9 (.B( u1_u12_u4_n136 ) , .A( u1_u12_u4_n137 ) , .C2( u1_u12_u4_n138 ) , .ZN( u1_u12_u4_n139 ) , .C1( u1_u12_u4_n182 ) );
  AOI22_X1 u1_u12_u4_U90 (.ZN( u1_u12_u4_n125 ) , .B2( u1_u12_u4_n131 ) , .A2( u1_u12_u4_n132 ) , .B1( u1_u12_u4_n138 ) , .A1( u1_u12_u4_n178 ) );
  NAND4_X1 u1_u12_u4_U91 (.ZN( u1_out12_8 ) , .A4( u1_u12_u4_n110 ) , .A3( u1_u12_u4_n111 ) , .A2( u1_u12_u4_n112 ) , .A1( u1_u12_u4_n186 ) );
  NAND2_X1 u1_u12_u4_U92 (.ZN( u1_u12_u4_n112 ) , .A2( u1_u12_u4_n130 ) , .A1( u1_u12_u4_n150 ) );
  AOI22_X1 u1_u12_u4_U93 (.ZN( u1_u12_u4_n111 ) , .B2( u1_u12_u4_n132 ) , .A1( u1_u12_u4_n152 ) , .B1( u1_u12_u4_n178 ) , .A2( u1_u12_u4_n97 ) );
  AOI22_X1 u1_u12_u4_U94 (.B2( u1_u12_u4_n149 ) , .B1( u1_u12_u4_n150 ) , .A2( u1_u12_u4_n151 ) , .A1( u1_u12_u4_n152 ) , .ZN( u1_u12_u4_n167 ) );
  NOR4_X1 u1_u12_u4_U95 (.A4( u1_u12_u4_n162 ) , .A3( u1_u12_u4_n163 ) , .A2( u1_u12_u4_n164 ) , .A1( u1_u12_u4_n165 ) , .ZN( u1_u12_u4_n166 ) );
  NAND3_X1 u1_u12_u4_U96 (.ZN( u1_out12_3 ) , .A3( u1_u12_u4_n166 ) , .A1( u1_u12_u4_n167 ) , .A2( u1_u12_u4_n186 ) );
  NAND3_X1 u1_u12_u4_U97 (.A3( u1_u12_u4_n146 ) , .A2( u1_u12_u4_n147 ) , .A1( u1_u12_u4_n148 ) , .ZN( u1_u12_u4_n149 ) );
  NAND3_X1 u1_u12_u4_U98 (.A3( u1_u12_u4_n143 ) , .A2( u1_u12_u4_n144 ) , .A1( u1_u12_u4_n145 ) , .ZN( u1_u12_u4_n151 ) );
  NAND3_X1 u1_u12_u4_U99 (.A3( u1_u12_u4_n121 ) , .ZN( u1_u12_u4_n122 ) , .A2( u1_u12_u4_n144 ) , .A1( u1_u12_u4_n154 ) );
  AND3_X1 u1_u12_u7_U10 (.A3( u1_u12_u7_n110 ) , .A2( u1_u12_u7_n127 ) , .A1( u1_u12_u7_n132 ) , .ZN( u1_u12_u7_n92 ) );
  OAI21_X1 u1_u12_u7_U11 (.A( u1_u12_u7_n161 ) , .B1( u1_u12_u7_n168 ) , .B2( u1_u12_u7_n173 ) , .ZN( u1_u12_u7_n91 ) );
  AOI211_X1 u1_u12_u7_U12 (.A( u1_u12_u7_n117 ) , .ZN( u1_u12_u7_n118 ) , .C2( u1_u12_u7_n126 ) , .C1( u1_u12_u7_n177 ) , .B( u1_u12_u7_n180 ) );
  OAI22_X1 u1_u12_u7_U13 (.B1( u1_u12_u7_n115 ) , .ZN( u1_u12_u7_n117 ) , .A2( u1_u12_u7_n133 ) , .A1( u1_u12_u7_n137 ) , .B2( u1_u12_u7_n162 ) );
  INV_X1 u1_u12_u7_U14 (.A( u1_u12_u7_n116 ) , .ZN( u1_u12_u7_n180 ) );
  NOR3_X1 u1_u12_u7_U15 (.ZN( u1_u12_u7_n115 ) , .A3( u1_u12_u7_n145 ) , .A2( u1_u12_u7_n168 ) , .A1( u1_u12_u7_n169 ) );
  OAI211_X1 u1_u12_u7_U16 (.B( u1_u12_u7_n122 ) , .A( u1_u12_u7_n123 ) , .C2( u1_u12_u7_n124 ) , .ZN( u1_u12_u7_n154 ) , .C1( u1_u12_u7_n162 ) );
  AOI222_X1 u1_u12_u7_U17 (.ZN( u1_u12_u7_n122 ) , .C2( u1_u12_u7_n126 ) , .C1( u1_u12_u7_n145 ) , .B1( u1_u12_u7_n161 ) , .A2( u1_u12_u7_n165 ) , .B2( u1_u12_u7_n170 ) , .A1( u1_u12_u7_n176 ) );
  INV_X1 u1_u12_u7_U18 (.A( u1_u12_u7_n133 ) , .ZN( u1_u12_u7_n176 ) );
  NOR3_X1 u1_u12_u7_U19 (.A2( u1_u12_u7_n134 ) , .A1( u1_u12_u7_n135 ) , .ZN( u1_u12_u7_n136 ) , .A3( u1_u12_u7_n171 ) );
  NOR2_X1 u1_u12_u7_U20 (.A1( u1_u12_u7_n130 ) , .A2( u1_u12_u7_n134 ) , .ZN( u1_u12_u7_n153 ) );
  INV_X1 u1_u12_u7_U21 (.A( u1_u12_u7_n101 ) , .ZN( u1_u12_u7_n165 ) );
  NOR2_X1 u1_u12_u7_U22 (.ZN( u1_u12_u7_n111 ) , .A2( u1_u12_u7_n134 ) , .A1( u1_u12_u7_n169 ) );
  AOI21_X1 u1_u12_u7_U23 (.ZN( u1_u12_u7_n104 ) , .B2( u1_u12_u7_n112 ) , .B1( u1_u12_u7_n127 ) , .A( u1_u12_u7_n164 ) );
  AOI21_X1 u1_u12_u7_U24 (.ZN( u1_u12_u7_n106 ) , .B1( u1_u12_u7_n133 ) , .B2( u1_u12_u7_n146 ) , .A( u1_u12_u7_n162 ) );
  AOI21_X1 u1_u12_u7_U25 (.A( u1_u12_u7_n101 ) , .ZN( u1_u12_u7_n107 ) , .B2( u1_u12_u7_n128 ) , .B1( u1_u12_u7_n175 ) );
  INV_X1 u1_u12_u7_U26 (.A( u1_u12_u7_n138 ) , .ZN( u1_u12_u7_n171 ) );
  INV_X1 u1_u12_u7_U27 (.A( u1_u12_u7_n131 ) , .ZN( u1_u12_u7_n177 ) );
  INV_X1 u1_u12_u7_U28 (.A( u1_u12_u7_n110 ) , .ZN( u1_u12_u7_n174 ) );
  NAND2_X1 u1_u12_u7_U29 (.A1( u1_u12_u7_n129 ) , .A2( u1_u12_u7_n132 ) , .ZN( u1_u12_u7_n149 ) );
  OAI21_X1 u1_u12_u7_U3 (.ZN( u1_u12_u7_n159 ) , .A( u1_u12_u7_n165 ) , .B2( u1_u12_u7_n171 ) , .B1( u1_u12_u7_n174 ) );
  NAND2_X1 u1_u12_u7_U30 (.A1( u1_u12_u7_n113 ) , .A2( u1_u12_u7_n124 ) , .ZN( u1_u12_u7_n130 ) );
  INV_X1 u1_u12_u7_U31 (.A( u1_u12_u7_n112 ) , .ZN( u1_u12_u7_n173 ) );
  INV_X1 u1_u12_u7_U32 (.A( u1_u12_u7_n128 ) , .ZN( u1_u12_u7_n168 ) );
  INV_X1 u1_u12_u7_U33 (.A( u1_u12_u7_n148 ) , .ZN( u1_u12_u7_n169 ) );
  INV_X1 u1_u12_u7_U34 (.A( u1_u12_u7_n127 ) , .ZN( u1_u12_u7_n179 ) );
  NOR2_X1 u1_u12_u7_U35 (.ZN( u1_u12_u7_n101 ) , .A2( u1_u12_u7_n150 ) , .A1( u1_u12_u7_n156 ) );
  AOI211_X1 u1_u12_u7_U36 (.B( u1_u12_u7_n154 ) , .A( u1_u12_u7_n155 ) , .C1( u1_u12_u7_n156 ) , .ZN( u1_u12_u7_n157 ) , .C2( u1_u12_u7_n172 ) );
  INV_X1 u1_u12_u7_U37 (.A( u1_u12_u7_n153 ) , .ZN( u1_u12_u7_n172 ) );
  AOI211_X1 u1_u12_u7_U38 (.B( u1_u12_u7_n139 ) , .A( u1_u12_u7_n140 ) , .C2( u1_u12_u7_n141 ) , .ZN( u1_u12_u7_n142 ) , .C1( u1_u12_u7_n156 ) );
  NAND4_X1 u1_u12_u7_U39 (.A3( u1_u12_u7_n127 ) , .A2( u1_u12_u7_n128 ) , .A1( u1_u12_u7_n129 ) , .ZN( u1_u12_u7_n141 ) , .A4( u1_u12_u7_n147 ) );
  INV_X1 u1_u12_u7_U4 (.A( u1_u12_u7_n111 ) , .ZN( u1_u12_u7_n170 ) );
  AOI21_X1 u1_u12_u7_U40 (.A( u1_u12_u7_n137 ) , .B1( u1_u12_u7_n138 ) , .ZN( u1_u12_u7_n139 ) , .B2( u1_u12_u7_n146 ) );
  OAI22_X1 u1_u12_u7_U41 (.B1( u1_u12_u7_n136 ) , .ZN( u1_u12_u7_n140 ) , .A1( u1_u12_u7_n153 ) , .B2( u1_u12_u7_n162 ) , .A2( u1_u12_u7_n164 ) );
  AOI21_X1 u1_u12_u7_U42 (.ZN( u1_u12_u7_n123 ) , .B1( u1_u12_u7_n165 ) , .B2( u1_u12_u7_n177 ) , .A( u1_u12_u7_n97 ) );
  AOI21_X1 u1_u12_u7_U43 (.B2( u1_u12_u7_n113 ) , .B1( u1_u12_u7_n124 ) , .A( u1_u12_u7_n125 ) , .ZN( u1_u12_u7_n97 ) );
  INV_X1 u1_u12_u7_U44 (.A( u1_u12_u7_n125 ) , .ZN( u1_u12_u7_n161 ) );
  INV_X1 u1_u12_u7_U45 (.A( u1_u12_u7_n152 ) , .ZN( u1_u12_u7_n162 ) );
  AOI22_X1 u1_u12_u7_U46 (.A2( u1_u12_u7_n114 ) , .ZN( u1_u12_u7_n119 ) , .B1( u1_u12_u7_n130 ) , .A1( u1_u12_u7_n156 ) , .B2( u1_u12_u7_n165 ) );
  NAND2_X1 u1_u12_u7_U47 (.A2( u1_u12_u7_n112 ) , .ZN( u1_u12_u7_n114 ) , .A1( u1_u12_u7_n175 ) );
  AND2_X1 u1_u12_u7_U48 (.ZN( u1_u12_u7_n145 ) , .A2( u1_u12_u7_n98 ) , .A1( u1_u12_u7_n99 ) );
  NOR2_X1 u1_u12_u7_U49 (.ZN( u1_u12_u7_n137 ) , .A1( u1_u12_u7_n150 ) , .A2( u1_u12_u7_n161 ) );
  INV_X1 u1_u12_u7_U5 (.A( u1_u12_u7_n149 ) , .ZN( u1_u12_u7_n175 ) );
  AOI21_X1 u1_u12_u7_U50 (.ZN( u1_u12_u7_n105 ) , .B2( u1_u12_u7_n110 ) , .A( u1_u12_u7_n125 ) , .B1( u1_u12_u7_n147 ) );
  NAND2_X1 u1_u12_u7_U51 (.ZN( u1_u12_u7_n146 ) , .A1( u1_u12_u7_n95 ) , .A2( u1_u12_u7_n98 ) );
  NAND2_X1 u1_u12_u7_U52 (.A2( u1_u12_u7_n103 ) , .ZN( u1_u12_u7_n147 ) , .A1( u1_u12_u7_n93 ) );
  NAND2_X1 u1_u12_u7_U53 (.A1( u1_u12_u7_n103 ) , .ZN( u1_u12_u7_n127 ) , .A2( u1_u12_u7_n99 ) );
  OR2_X1 u1_u12_u7_U54 (.ZN( u1_u12_u7_n126 ) , .A2( u1_u12_u7_n152 ) , .A1( u1_u12_u7_n156 ) );
  NAND2_X1 u1_u12_u7_U55 (.A2( u1_u12_u7_n102 ) , .A1( u1_u12_u7_n103 ) , .ZN( u1_u12_u7_n133 ) );
  NAND2_X1 u1_u12_u7_U56 (.ZN( u1_u12_u7_n112 ) , .A2( u1_u12_u7_n96 ) , .A1( u1_u12_u7_n99 ) );
  NAND2_X1 u1_u12_u7_U57 (.A2( u1_u12_u7_n102 ) , .ZN( u1_u12_u7_n128 ) , .A1( u1_u12_u7_n98 ) );
  NAND2_X1 u1_u12_u7_U58 (.A1( u1_u12_u7_n100 ) , .ZN( u1_u12_u7_n113 ) , .A2( u1_u12_u7_n93 ) );
  NAND2_X1 u1_u12_u7_U59 (.A2( u1_u12_u7_n102 ) , .ZN( u1_u12_u7_n124 ) , .A1( u1_u12_u7_n96 ) );
  INV_X1 u1_u12_u7_U6 (.A( u1_u12_u7_n154 ) , .ZN( u1_u12_u7_n178 ) );
  NAND2_X1 u1_u12_u7_U60 (.ZN( u1_u12_u7_n110 ) , .A1( u1_u12_u7_n95 ) , .A2( u1_u12_u7_n96 ) );
  INV_X1 u1_u12_u7_U61 (.A( u1_u12_u7_n150 ) , .ZN( u1_u12_u7_n164 ) );
  AND2_X1 u1_u12_u7_U62 (.ZN( u1_u12_u7_n134 ) , .A1( u1_u12_u7_n93 ) , .A2( u1_u12_u7_n98 ) );
  NAND2_X1 u1_u12_u7_U63 (.A1( u1_u12_u7_n100 ) , .A2( u1_u12_u7_n102 ) , .ZN( u1_u12_u7_n129 ) );
  NAND2_X1 u1_u12_u7_U64 (.A2( u1_u12_u7_n103 ) , .ZN( u1_u12_u7_n131 ) , .A1( u1_u12_u7_n95 ) );
  NAND2_X1 u1_u12_u7_U65 (.A1( u1_u12_u7_n100 ) , .ZN( u1_u12_u7_n138 ) , .A2( u1_u12_u7_n99 ) );
  NAND2_X1 u1_u12_u7_U66 (.ZN( u1_u12_u7_n132 ) , .A1( u1_u12_u7_n93 ) , .A2( u1_u12_u7_n96 ) );
  NAND2_X1 u1_u12_u7_U67 (.A1( u1_u12_u7_n100 ) , .ZN( u1_u12_u7_n148 ) , .A2( u1_u12_u7_n95 ) );
  NOR2_X1 u1_u12_u7_U68 (.A2( u1_u12_X_47 ) , .ZN( u1_u12_u7_n150 ) , .A1( u1_u12_u7_n163 ) );
  NOR2_X1 u1_u12_u7_U69 (.A2( u1_u12_X_43 ) , .A1( u1_u12_X_44 ) , .ZN( u1_u12_u7_n103 ) );
  AOI211_X1 u1_u12_u7_U7 (.ZN( u1_u12_u7_n116 ) , .A( u1_u12_u7_n155 ) , .C1( u1_u12_u7_n161 ) , .C2( u1_u12_u7_n171 ) , .B( u1_u12_u7_n94 ) );
  NOR2_X1 u1_u12_u7_U70 (.A2( u1_u12_X_48 ) , .A1( u1_u12_u7_n166 ) , .ZN( u1_u12_u7_n95 ) );
  NOR2_X1 u1_u12_u7_U71 (.A2( u1_u12_X_45 ) , .A1( u1_u12_X_48 ) , .ZN( u1_u12_u7_n99 ) );
  NOR2_X1 u1_u12_u7_U72 (.A2( u1_u12_X_44 ) , .A1( u1_u12_u7_n167 ) , .ZN( u1_u12_u7_n98 ) );
  NOR2_X1 u1_u12_u7_U73 (.A2( u1_u12_X_46 ) , .A1( u1_u12_X_47 ) , .ZN( u1_u12_u7_n152 ) );
  AND2_X1 u1_u12_u7_U74 (.A1( u1_u12_X_47 ) , .ZN( u1_u12_u7_n156 ) , .A2( u1_u12_u7_n163 ) );
  NAND2_X1 u1_u12_u7_U75 (.A2( u1_u12_X_46 ) , .A1( u1_u12_X_47 ) , .ZN( u1_u12_u7_n125 ) );
  AND2_X1 u1_u12_u7_U76 (.A2( u1_u12_X_45 ) , .A1( u1_u12_X_48 ) , .ZN( u1_u12_u7_n102 ) );
  AND2_X1 u1_u12_u7_U77 (.A2( u1_u12_X_43 ) , .A1( u1_u12_X_44 ) , .ZN( u1_u12_u7_n96 ) );
  AND2_X1 u1_u12_u7_U78 (.A1( u1_u12_X_44 ) , .ZN( u1_u12_u7_n100 ) , .A2( u1_u12_u7_n167 ) );
  AND2_X1 u1_u12_u7_U79 (.A1( u1_u12_X_48 ) , .A2( u1_u12_u7_n166 ) , .ZN( u1_u12_u7_n93 ) );
  OAI222_X1 u1_u12_u7_U8 (.C2( u1_u12_u7_n101 ) , .B2( u1_u12_u7_n111 ) , .A1( u1_u12_u7_n113 ) , .C1( u1_u12_u7_n146 ) , .A2( u1_u12_u7_n162 ) , .B1( u1_u12_u7_n164 ) , .ZN( u1_u12_u7_n94 ) );
  INV_X1 u1_u12_u7_U80 (.A( u1_u12_X_46 ) , .ZN( u1_u12_u7_n163 ) );
  INV_X1 u1_u12_u7_U81 (.A( u1_u12_X_43 ) , .ZN( u1_u12_u7_n167 ) );
  INV_X1 u1_u12_u7_U82 (.A( u1_u12_X_45 ) , .ZN( u1_u12_u7_n166 ) );
  NAND4_X1 u1_u12_u7_U83 (.ZN( u1_out12_5 ) , .A4( u1_u12_u7_n108 ) , .A3( u1_u12_u7_n109 ) , .A1( u1_u12_u7_n116 ) , .A2( u1_u12_u7_n123 ) );
  AOI22_X1 u1_u12_u7_U84 (.ZN( u1_u12_u7_n109 ) , .A2( u1_u12_u7_n126 ) , .B2( u1_u12_u7_n145 ) , .B1( u1_u12_u7_n156 ) , .A1( u1_u12_u7_n171 ) );
  NOR4_X1 u1_u12_u7_U85 (.A4( u1_u12_u7_n104 ) , .A3( u1_u12_u7_n105 ) , .A2( u1_u12_u7_n106 ) , .A1( u1_u12_u7_n107 ) , .ZN( u1_u12_u7_n108 ) );
  NAND4_X1 u1_u12_u7_U86 (.ZN( u1_out12_27 ) , .A4( u1_u12_u7_n118 ) , .A3( u1_u12_u7_n119 ) , .A2( u1_u12_u7_n120 ) , .A1( u1_u12_u7_n121 ) );
  OAI21_X1 u1_u12_u7_U87 (.ZN( u1_u12_u7_n121 ) , .B2( u1_u12_u7_n145 ) , .A( u1_u12_u7_n150 ) , .B1( u1_u12_u7_n174 ) );
  OAI21_X1 u1_u12_u7_U88 (.ZN( u1_u12_u7_n120 ) , .A( u1_u12_u7_n161 ) , .B2( u1_u12_u7_n170 ) , .B1( u1_u12_u7_n179 ) );
  NAND4_X1 u1_u12_u7_U89 (.ZN( u1_out12_21 ) , .A4( u1_u12_u7_n157 ) , .A3( u1_u12_u7_n158 ) , .A2( u1_u12_u7_n159 ) , .A1( u1_u12_u7_n160 ) );
  OAI221_X1 u1_u12_u7_U9 (.C1( u1_u12_u7_n101 ) , .C2( u1_u12_u7_n147 ) , .ZN( u1_u12_u7_n155 ) , .B2( u1_u12_u7_n162 ) , .A( u1_u12_u7_n91 ) , .B1( u1_u12_u7_n92 ) );
  OAI21_X1 u1_u12_u7_U90 (.B1( u1_u12_u7_n145 ) , .ZN( u1_u12_u7_n160 ) , .A( u1_u12_u7_n161 ) , .B2( u1_u12_u7_n177 ) );
  AOI22_X1 u1_u12_u7_U91 (.B2( u1_u12_u7_n149 ) , .B1( u1_u12_u7_n150 ) , .A2( u1_u12_u7_n151 ) , .A1( u1_u12_u7_n152 ) , .ZN( u1_u12_u7_n158 ) );
  NAND4_X1 u1_u12_u7_U92 (.ZN( u1_out12_15 ) , .A4( u1_u12_u7_n142 ) , .A3( u1_u12_u7_n143 ) , .A2( u1_u12_u7_n144 ) , .A1( u1_u12_u7_n178 ) );
  OR2_X1 u1_u12_u7_U93 (.A2( u1_u12_u7_n125 ) , .A1( u1_u12_u7_n129 ) , .ZN( u1_u12_u7_n144 ) );
  AOI22_X1 u1_u12_u7_U94 (.A2( u1_u12_u7_n126 ) , .ZN( u1_u12_u7_n143 ) , .B2( u1_u12_u7_n165 ) , .B1( u1_u12_u7_n173 ) , .A1( u1_u12_u7_n174 ) );
  NAND3_X1 u1_u12_u7_U95 (.A3( u1_u12_u7_n146 ) , .A2( u1_u12_u7_n147 ) , .A1( u1_u12_u7_n148 ) , .ZN( u1_u12_u7_n151 ) );
  NAND3_X1 u1_u12_u7_U96 (.A3( u1_u12_u7_n131 ) , .A2( u1_u12_u7_n132 ) , .A1( u1_u12_u7_n133 ) , .ZN( u1_u12_u7_n135 ) );
  XOR2_X1 u1_u14_U35 (.B( u1_K15_22 ) , .A( u1_R13_15 ) , .Z( u1_u14_X_22 ) );
  XOR2_X1 u1_u14_U36 (.B( u1_K15_21 ) , .A( u1_R13_14 ) , .Z( u1_u14_X_21 ) );
  XOR2_X1 u1_u14_U37 (.B( u1_K15_20 ) , .A( u1_R13_13 ) , .Z( u1_u14_X_20 ) );
  XOR2_X1 u1_u14_U39 (.B( u1_K15_19 ) , .A( u1_R13_12 ) , .Z( u1_u14_X_19 ) );
  XOR2_X1 u1_u14_U40 (.B( u1_K15_18 ) , .A( u1_R13_13 ) , .Z( u1_u14_X_18 ) );
  XOR2_X1 u1_u14_U41 (.B( u1_K15_17 ) , .A( u1_R13_12 ) , .Z( u1_u14_X_17 ) );
  XOR2_X1 u1_u14_U42 (.B( u1_K15_16 ) , .A( u1_R13_11 ) , .Z( u1_u14_X_16 ) );
  XOR2_X1 u1_u14_U43 (.B( u1_K15_15 ) , .A( u1_R13_10 ) , .Z( u1_u14_X_15 ) );
  XOR2_X1 u1_u14_U44 (.B( u1_K15_14 ) , .A( u1_R13_9 ) , .Z( u1_u14_X_14 ) );
  OAI22_X1 u1_u14_u2_U10 (.ZN( u1_u14_u2_n109 ) , .A2( u1_u14_u2_n113 ) , .B2( u1_u14_u2_n133 ) , .B1( u1_u14_u2_n167 ) , .A1( u1_u14_u2_n168 ) );
  NAND3_X1 u1_u14_u2_U100 (.A2( u1_u14_u2_n100 ) , .A1( u1_u14_u2_n104 ) , .A3( u1_u14_u2_n138 ) , .ZN( u1_u14_u2_n98 ) );
  OAI22_X1 u1_u14_u2_U11 (.B1( u1_u14_u2_n151 ) , .A2( u1_u14_u2_n152 ) , .A1( u1_u14_u2_n153 ) , .ZN( u1_u14_u2_n160 ) , .B2( u1_u14_u2_n168 ) );
  NOR3_X1 u1_u14_u2_U12 (.A1( u1_u14_u2_n150 ) , .ZN( u1_u14_u2_n151 ) , .A3( u1_u14_u2_n175 ) , .A2( u1_u14_u2_n188 ) );
  AOI21_X1 u1_u14_u2_U13 (.ZN( u1_u14_u2_n144 ) , .B2( u1_u14_u2_n155 ) , .A( u1_u14_u2_n172 ) , .B1( u1_u14_u2_n185 ) );
  AOI21_X1 u1_u14_u2_U14 (.B2( u1_u14_u2_n143 ) , .ZN( u1_u14_u2_n145 ) , .B1( u1_u14_u2_n152 ) , .A( u1_u14_u2_n171 ) );
  AOI21_X1 u1_u14_u2_U15 (.B2( u1_u14_u2_n120 ) , .B1( u1_u14_u2_n121 ) , .ZN( u1_u14_u2_n126 ) , .A( u1_u14_u2_n167 ) );
  INV_X1 u1_u14_u2_U16 (.A( u1_u14_u2_n156 ) , .ZN( u1_u14_u2_n171 ) );
  INV_X1 u1_u14_u2_U17 (.A( u1_u14_u2_n120 ) , .ZN( u1_u14_u2_n188 ) );
  NAND2_X1 u1_u14_u2_U18 (.A2( u1_u14_u2_n122 ) , .ZN( u1_u14_u2_n150 ) , .A1( u1_u14_u2_n152 ) );
  INV_X1 u1_u14_u2_U19 (.A( u1_u14_u2_n153 ) , .ZN( u1_u14_u2_n170 ) );
  INV_X1 u1_u14_u2_U20 (.A( u1_u14_u2_n137 ) , .ZN( u1_u14_u2_n173 ) );
  NAND2_X1 u1_u14_u2_U21 (.A1( u1_u14_u2_n132 ) , .A2( u1_u14_u2_n139 ) , .ZN( u1_u14_u2_n157 ) );
  INV_X1 u1_u14_u2_U22 (.A( u1_u14_u2_n113 ) , .ZN( u1_u14_u2_n178 ) );
  INV_X1 u1_u14_u2_U23 (.A( u1_u14_u2_n139 ) , .ZN( u1_u14_u2_n175 ) );
  INV_X1 u1_u14_u2_U24 (.A( u1_u14_u2_n155 ) , .ZN( u1_u14_u2_n181 ) );
  INV_X1 u1_u14_u2_U25 (.A( u1_u14_u2_n119 ) , .ZN( u1_u14_u2_n177 ) );
  INV_X1 u1_u14_u2_U26 (.A( u1_u14_u2_n116 ) , .ZN( u1_u14_u2_n180 ) );
  INV_X1 u1_u14_u2_U27 (.A( u1_u14_u2_n131 ) , .ZN( u1_u14_u2_n179 ) );
  INV_X1 u1_u14_u2_U28 (.A( u1_u14_u2_n154 ) , .ZN( u1_u14_u2_n176 ) );
  NAND2_X1 u1_u14_u2_U29 (.A2( u1_u14_u2_n116 ) , .A1( u1_u14_u2_n117 ) , .ZN( u1_u14_u2_n118 ) );
  NOR2_X1 u1_u14_u2_U3 (.ZN( u1_u14_u2_n121 ) , .A2( u1_u14_u2_n177 ) , .A1( u1_u14_u2_n180 ) );
  INV_X1 u1_u14_u2_U30 (.A( u1_u14_u2_n132 ) , .ZN( u1_u14_u2_n182 ) );
  INV_X1 u1_u14_u2_U31 (.A( u1_u14_u2_n158 ) , .ZN( u1_u14_u2_n183 ) );
  OAI21_X1 u1_u14_u2_U32 (.A( u1_u14_u2_n156 ) , .B1( u1_u14_u2_n157 ) , .ZN( u1_u14_u2_n158 ) , .B2( u1_u14_u2_n179 ) );
  NOR2_X1 u1_u14_u2_U33 (.ZN( u1_u14_u2_n156 ) , .A1( u1_u14_u2_n166 ) , .A2( u1_u14_u2_n169 ) );
  NOR2_X1 u1_u14_u2_U34 (.A2( u1_u14_u2_n114 ) , .ZN( u1_u14_u2_n137 ) , .A1( u1_u14_u2_n140 ) );
  NOR2_X1 u1_u14_u2_U35 (.A2( u1_u14_u2_n138 ) , .ZN( u1_u14_u2_n153 ) , .A1( u1_u14_u2_n156 ) );
  AOI211_X1 u1_u14_u2_U36 (.ZN( u1_u14_u2_n130 ) , .C1( u1_u14_u2_n138 ) , .C2( u1_u14_u2_n179 ) , .B( u1_u14_u2_n96 ) , .A( u1_u14_u2_n97 ) );
  OAI22_X1 u1_u14_u2_U37 (.B1( u1_u14_u2_n133 ) , .A2( u1_u14_u2_n137 ) , .A1( u1_u14_u2_n152 ) , .B2( u1_u14_u2_n168 ) , .ZN( u1_u14_u2_n97 ) );
  OAI221_X1 u1_u14_u2_U38 (.B1( u1_u14_u2_n113 ) , .C1( u1_u14_u2_n132 ) , .A( u1_u14_u2_n149 ) , .B2( u1_u14_u2_n171 ) , .C2( u1_u14_u2_n172 ) , .ZN( u1_u14_u2_n96 ) );
  OAI221_X1 u1_u14_u2_U39 (.A( u1_u14_u2_n115 ) , .C2( u1_u14_u2_n123 ) , .B2( u1_u14_u2_n143 ) , .B1( u1_u14_u2_n153 ) , .ZN( u1_u14_u2_n163 ) , .C1( u1_u14_u2_n168 ) );
  INV_X1 u1_u14_u2_U4 (.A( u1_u14_u2_n134 ) , .ZN( u1_u14_u2_n185 ) );
  OAI21_X1 u1_u14_u2_U40 (.A( u1_u14_u2_n114 ) , .ZN( u1_u14_u2_n115 ) , .B1( u1_u14_u2_n176 ) , .B2( u1_u14_u2_n178 ) );
  OAI221_X1 u1_u14_u2_U41 (.A( u1_u14_u2_n135 ) , .B2( u1_u14_u2_n136 ) , .B1( u1_u14_u2_n137 ) , .ZN( u1_u14_u2_n162 ) , .C2( u1_u14_u2_n167 ) , .C1( u1_u14_u2_n185 ) );
  AND3_X1 u1_u14_u2_U42 (.A3( u1_u14_u2_n131 ) , .A2( u1_u14_u2_n132 ) , .A1( u1_u14_u2_n133 ) , .ZN( u1_u14_u2_n136 ) );
  AOI22_X1 u1_u14_u2_U43 (.ZN( u1_u14_u2_n135 ) , .B1( u1_u14_u2_n140 ) , .A1( u1_u14_u2_n156 ) , .B2( u1_u14_u2_n180 ) , .A2( u1_u14_u2_n188 ) );
  AOI21_X1 u1_u14_u2_U44 (.ZN( u1_u14_u2_n149 ) , .B1( u1_u14_u2_n173 ) , .B2( u1_u14_u2_n188 ) , .A( u1_u14_u2_n95 ) );
  AND3_X1 u1_u14_u2_U45 (.A2( u1_u14_u2_n100 ) , .A1( u1_u14_u2_n104 ) , .A3( u1_u14_u2_n156 ) , .ZN( u1_u14_u2_n95 ) );
  OAI21_X1 u1_u14_u2_U46 (.A( u1_u14_u2_n101 ) , .B2( u1_u14_u2_n121 ) , .B1( u1_u14_u2_n153 ) , .ZN( u1_u14_u2_n164 ) );
  NAND2_X1 u1_u14_u2_U47 (.A2( u1_u14_u2_n100 ) , .A1( u1_u14_u2_n107 ) , .ZN( u1_u14_u2_n155 ) );
  NAND2_X1 u1_u14_u2_U48 (.A2( u1_u14_u2_n105 ) , .A1( u1_u14_u2_n108 ) , .ZN( u1_u14_u2_n143 ) );
  NAND2_X1 u1_u14_u2_U49 (.A1( u1_u14_u2_n104 ) , .A2( u1_u14_u2_n106 ) , .ZN( u1_u14_u2_n152 ) );
  INV_X1 u1_u14_u2_U5 (.A( u1_u14_u2_n150 ) , .ZN( u1_u14_u2_n184 ) );
  NAND2_X1 u1_u14_u2_U50 (.A1( u1_u14_u2_n100 ) , .A2( u1_u14_u2_n105 ) , .ZN( u1_u14_u2_n132 ) );
  INV_X1 u1_u14_u2_U51 (.A( u1_u14_u2_n140 ) , .ZN( u1_u14_u2_n168 ) );
  INV_X1 u1_u14_u2_U52 (.A( u1_u14_u2_n138 ) , .ZN( u1_u14_u2_n167 ) );
  OAI21_X1 u1_u14_u2_U53 (.A( u1_u14_u2_n141 ) , .B2( u1_u14_u2_n142 ) , .ZN( u1_u14_u2_n146 ) , .B1( u1_u14_u2_n153 ) );
  OAI21_X1 u1_u14_u2_U54 (.A( u1_u14_u2_n140 ) , .ZN( u1_u14_u2_n141 ) , .B1( u1_u14_u2_n176 ) , .B2( u1_u14_u2_n177 ) );
  NOR3_X1 u1_u14_u2_U55 (.ZN( u1_u14_u2_n142 ) , .A3( u1_u14_u2_n175 ) , .A2( u1_u14_u2_n178 ) , .A1( u1_u14_u2_n181 ) );
  INV_X1 u1_u14_u2_U56 (.ZN( u1_u14_u2_n187 ) , .A( u1_u14_u2_n99 ) );
  OAI21_X1 u1_u14_u2_U57 (.B1( u1_u14_u2_n137 ) , .B2( u1_u14_u2_n143 ) , .A( u1_u14_u2_n98 ) , .ZN( u1_u14_u2_n99 ) );
  NAND2_X1 u1_u14_u2_U58 (.A1( u1_u14_u2_n102 ) , .A2( u1_u14_u2_n106 ) , .ZN( u1_u14_u2_n113 ) );
  NAND2_X1 u1_u14_u2_U59 (.A1( u1_u14_u2_n106 ) , .A2( u1_u14_u2_n107 ) , .ZN( u1_u14_u2_n131 ) );
  NOR4_X1 u1_u14_u2_U6 (.A4( u1_u14_u2_n124 ) , .A3( u1_u14_u2_n125 ) , .A2( u1_u14_u2_n126 ) , .A1( u1_u14_u2_n127 ) , .ZN( u1_u14_u2_n128 ) );
  NAND2_X1 u1_u14_u2_U60 (.A1( u1_u14_u2_n103 ) , .A2( u1_u14_u2_n107 ) , .ZN( u1_u14_u2_n139 ) );
  NAND2_X1 u1_u14_u2_U61 (.A1( u1_u14_u2_n103 ) , .A2( u1_u14_u2_n105 ) , .ZN( u1_u14_u2_n133 ) );
  NAND2_X1 u1_u14_u2_U62 (.A1( u1_u14_u2_n102 ) , .A2( u1_u14_u2_n103 ) , .ZN( u1_u14_u2_n154 ) );
  NAND2_X1 u1_u14_u2_U63 (.A2( u1_u14_u2_n103 ) , .A1( u1_u14_u2_n104 ) , .ZN( u1_u14_u2_n119 ) );
  NAND2_X1 u1_u14_u2_U64 (.A2( u1_u14_u2_n107 ) , .A1( u1_u14_u2_n108 ) , .ZN( u1_u14_u2_n123 ) );
  NAND2_X1 u1_u14_u2_U65 (.A1( u1_u14_u2_n104 ) , .A2( u1_u14_u2_n108 ) , .ZN( u1_u14_u2_n122 ) );
  INV_X1 u1_u14_u2_U66 (.A( u1_u14_u2_n114 ) , .ZN( u1_u14_u2_n172 ) );
  NAND2_X1 u1_u14_u2_U67 (.A2( u1_u14_u2_n100 ) , .A1( u1_u14_u2_n102 ) , .ZN( u1_u14_u2_n116 ) );
  NAND2_X1 u1_u14_u2_U68 (.A1( u1_u14_u2_n102 ) , .A2( u1_u14_u2_n108 ) , .ZN( u1_u14_u2_n120 ) );
  NAND2_X1 u1_u14_u2_U69 (.A2( u1_u14_u2_n105 ) , .A1( u1_u14_u2_n106 ) , .ZN( u1_u14_u2_n117 ) );
  AOI21_X1 u1_u14_u2_U7 (.B2( u1_u14_u2_n119 ) , .ZN( u1_u14_u2_n127 ) , .A( u1_u14_u2_n137 ) , .B1( u1_u14_u2_n155 ) );
  NOR2_X1 u1_u14_u2_U70 (.A2( u1_u14_X_16 ) , .ZN( u1_u14_u2_n140 ) , .A1( u1_u14_u2_n166 ) );
  NOR2_X1 u1_u14_u2_U71 (.A2( u1_u14_X_13 ) , .A1( u1_u14_X_14 ) , .ZN( u1_u14_u2_n100 ) );
  NOR2_X1 u1_u14_u2_U72 (.A2( u1_u14_X_16 ) , .A1( u1_u14_X_17 ) , .ZN( u1_u14_u2_n138 ) );
  NOR2_X1 u1_u14_u2_U73 (.A2( u1_u14_X_15 ) , .A1( u1_u14_X_18 ) , .ZN( u1_u14_u2_n104 ) );
  NOR2_X1 u1_u14_u2_U74 (.A2( u1_u14_X_14 ) , .ZN( u1_u14_u2_n103 ) , .A1( u1_u14_u2_n174 ) );
  NOR2_X1 u1_u14_u2_U75 (.A2( u1_u14_X_15 ) , .ZN( u1_u14_u2_n102 ) , .A1( u1_u14_u2_n165 ) );
  NOR2_X1 u1_u14_u2_U76 (.A2( u1_u14_X_17 ) , .ZN( u1_u14_u2_n114 ) , .A1( u1_u14_u2_n169 ) );
  AND2_X1 u1_u14_u2_U77 (.A1( u1_u14_X_15 ) , .ZN( u1_u14_u2_n105 ) , .A2( u1_u14_u2_n165 ) );
  AND2_X1 u1_u14_u2_U78 (.A2( u1_u14_X_15 ) , .A1( u1_u14_X_18 ) , .ZN( u1_u14_u2_n107 ) );
  AND2_X1 u1_u14_u2_U79 (.A1( u1_u14_X_14 ) , .ZN( u1_u14_u2_n106 ) , .A2( u1_u14_u2_n174 ) );
  AOI21_X1 u1_u14_u2_U8 (.ZN( u1_u14_u2_n124 ) , .B1( u1_u14_u2_n131 ) , .B2( u1_u14_u2_n143 ) , .A( u1_u14_u2_n172 ) );
  AND2_X1 u1_u14_u2_U80 (.A1( u1_u14_X_13 ) , .A2( u1_u14_X_14 ) , .ZN( u1_u14_u2_n108 ) );
  INV_X1 u1_u14_u2_U81 (.A( u1_u14_X_16 ) , .ZN( u1_u14_u2_n169 ) );
  INV_X1 u1_u14_u2_U82 (.A( u1_u14_X_17 ) , .ZN( u1_u14_u2_n166 ) );
  INV_X1 u1_u14_u2_U83 (.A( u1_u14_X_13 ) , .ZN( u1_u14_u2_n174 ) );
  INV_X1 u1_u14_u2_U84 (.A( u1_u14_X_18 ) , .ZN( u1_u14_u2_n165 ) );
  NAND4_X1 u1_u14_u2_U85 (.ZN( u1_out14_30 ) , .A4( u1_u14_u2_n147 ) , .A3( u1_u14_u2_n148 ) , .A2( u1_u14_u2_n149 ) , .A1( u1_u14_u2_n187 ) );
  NOR3_X1 u1_u14_u2_U86 (.A3( u1_u14_u2_n144 ) , .A2( u1_u14_u2_n145 ) , .A1( u1_u14_u2_n146 ) , .ZN( u1_u14_u2_n147 ) );
  AOI21_X1 u1_u14_u2_U87 (.B2( u1_u14_u2_n138 ) , .ZN( u1_u14_u2_n148 ) , .A( u1_u14_u2_n162 ) , .B1( u1_u14_u2_n182 ) );
  NAND4_X1 u1_u14_u2_U88 (.ZN( u1_out14_24 ) , .A4( u1_u14_u2_n111 ) , .A3( u1_u14_u2_n112 ) , .A1( u1_u14_u2_n130 ) , .A2( u1_u14_u2_n187 ) );
  AOI221_X1 u1_u14_u2_U89 (.A( u1_u14_u2_n109 ) , .B1( u1_u14_u2_n110 ) , .ZN( u1_u14_u2_n111 ) , .C1( u1_u14_u2_n134 ) , .C2( u1_u14_u2_n170 ) , .B2( u1_u14_u2_n173 ) );
  AOI21_X1 u1_u14_u2_U9 (.B2( u1_u14_u2_n123 ) , .ZN( u1_u14_u2_n125 ) , .A( u1_u14_u2_n171 ) , .B1( u1_u14_u2_n184 ) );
  AOI21_X1 u1_u14_u2_U90 (.ZN( u1_u14_u2_n112 ) , .B2( u1_u14_u2_n156 ) , .A( u1_u14_u2_n164 ) , .B1( u1_u14_u2_n181 ) );
  NAND4_X1 u1_u14_u2_U91 (.ZN( u1_out14_16 ) , .A4( u1_u14_u2_n128 ) , .A3( u1_u14_u2_n129 ) , .A1( u1_u14_u2_n130 ) , .A2( u1_u14_u2_n186 ) );
  AOI22_X1 u1_u14_u2_U92 (.A2( u1_u14_u2_n118 ) , .ZN( u1_u14_u2_n129 ) , .A1( u1_u14_u2_n140 ) , .B1( u1_u14_u2_n157 ) , .B2( u1_u14_u2_n170 ) );
  INV_X1 u1_u14_u2_U93 (.A( u1_u14_u2_n163 ) , .ZN( u1_u14_u2_n186 ) );
  OR4_X1 u1_u14_u2_U94 (.ZN( u1_out14_6 ) , .A4( u1_u14_u2_n161 ) , .A3( u1_u14_u2_n162 ) , .A2( u1_u14_u2_n163 ) , .A1( u1_u14_u2_n164 ) );
  OR3_X1 u1_u14_u2_U95 (.A2( u1_u14_u2_n159 ) , .A1( u1_u14_u2_n160 ) , .ZN( u1_u14_u2_n161 ) , .A3( u1_u14_u2_n183 ) );
  AOI21_X1 u1_u14_u2_U96 (.B2( u1_u14_u2_n154 ) , .B1( u1_u14_u2_n155 ) , .ZN( u1_u14_u2_n159 ) , .A( u1_u14_u2_n167 ) );
  NAND3_X1 u1_u14_u2_U97 (.A2( u1_u14_u2_n117 ) , .A1( u1_u14_u2_n122 ) , .A3( u1_u14_u2_n123 ) , .ZN( u1_u14_u2_n134 ) );
  NAND3_X1 u1_u14_u2_U98 (.ZN( u1_u14_u2_n110 ) , .A2( u1_u14_u2_n131 ) , .A3( u1_u14_u2_n139 ) , .A1( u1_u14_u2_n154 ) );
  NAND3_X1 u1_u14_u2_U99 (.A2( u1_u14_u2_n100 ) , .ZN( u1_u14_u2_n101 ) , .A1( u1_u14_u2_n104 ) , .A3( u1_u14_u2_n114 ) );
  OAI22_X1 u1_u14_u3_U10 (.B1( u1_u14_u3_n113 ) , .A2( u1_u14_u3_n135 ) , .A1( u1_u14_u3_n150 ) , .B2( u1_u14_u3_n164 ) , .ZN( u1_u14_u3_n98 ) );
  OAI211_X1 u1_u14_u3_U11 (.B( u1_u14_u3_n106 ) , .ZN( u1_u14_u3_n119 ) , .C2( u1_u14_u3_n128 ) , .C1( u1_u14_u3_n167 ) , .A( u1_u14_u3_n181 ) );
  AOI221_X1 u1_u14_u3_U12 (.C1( u1_u14_u3_n105 ) , .ZN( u1_u14_u3_n106 ) , .A( u1_u14_u3_n131 ) , .B2( u1_u14_u3_n132 ) , .C2( u1_u14_u3_n133 ) , .B1( u1_u14_u3_n169 ) );
  INV_X1 u1_u14_u3_U13 (.ZN( u1_u14_u3_n181 ) , .A( u1_u14_u3_n98 ) );
  NAND2_X1 u1_u14_u3_U14 (.ZN( u1_u14_u3_n105 ) , .A2( u1_u14_u3_n130 ) , .A1( u1_u14_u3_n155 ) );
  AOI22_X1 u1_u14_u3_U15 (.B1( u1_u14_u3_n115 ) , .A2( u1_u14_u3_n116 ) , .ZN( u1_u14_u3_n123 ) , .B2( u1_u14_u3_n133 ) , .A1( u1_u14_u3_n169 ) );
  NAND2_X1 u1_u14_u3_U16 (.ZN( u1_u14_u3_n116 ) , .A2( u1_u14_u3_n151 ) , .A1( u1_u14_u3_n182 ) );
  NOR2_X1 u1_u14_u3_U17 (.ZN( u1_u14_u3_n126 ) , .A2( u1_u14_u3_n150 ) , .A1( u1_u14_u3_n164 ) );
  AOI21_X1 u1_u14_u3_U18 (.ZN( u1_u14_u3_n112 ) , .B2( u1_u14_u3_n146 ) , .B1( u1_u14_u3_n155 ) , .A( u1_u14_u3_n167 ) );
  NAND2_X1 u1_u14_u3_U19 (.A1( u1_u14_u3_n135 ) , .ZN( u1_u14_u3_n142 ) , .A2( u1_u14_u3_n164 ) );
  NAND2_X1 u1_u14_u3_U20 (.ZN( u1_u14_u3_n132 ) , .A2( u1_u14_u3_n152 ) , .A1( u1_u14_u3_n156 ) );
  AND2_X1 u1_u14_u3_U21 (.A2( u1_u14_u3_n113 ) , .A1( u1_u14_u3_n114 ) , .ZN( u1_u14_u3_n151 ) );
  INV_X1 u1_u14_u3_U22 (.A( u1_u14_u3_n133 ) , .ZN( u1_u14_u3_n165 ) );
  INV_X1 u1_u14_u3_U23 (.A( u1_u14_u3_n135 ) , .ZN( u1_u14_u3_n170 ) );
  NAND2_X1 u1_u14_u3_U24 (.A1( u1_u14_u3_n107 ) , .A2( u1_u14_u3_n108 ) , .ZN( u1_u14_u3_n140 ) );
  NAND2_X1 u1_u14_u3_U25 (.ZN( u1_u14_u3_n117 ) , .A1( u1_u14_u3_n124 ) , .A2( u1_u14_u3_n148 ) );
  NAND2_X1 u1_u14_u3_U26 (.ZN( u1_u14_u3_n143 ) , .A1( u1_u14_u3_n165 ) , .A2( u1_u14_u3_n167 ) );
  INV_X1 u1_u14_u3_U27 (.A( u1_u14_u3_n130 ) , .ZN( u1_u14_u3_n177 ) );
  INV_X1 u1_u14_u3_U28 (.A( u1_u14_u3_n128 ) , .ZN( u1_u14_u3_n176 ) );
  INV_X1 u1_u14_u3_U29 (.A( u1_u14_u3_n155 ) , .ZN( u1_u14_u3_n174 ) );
  INV_X1 u1_u14_u3_U3 (.A( u1_u14_u3_n129 ) , .ZN( u1_u14_u3_n183 ) );
  INV_X1 u1_u14_u3_U30 (.A( u1_u14_u3_n139 ) , .ZN( u1_u14_u3_n185 ) );
  NOR2_X1 u1_u14_u3_U31 (.ZN( u1_u14_u3_n135 ) , .A2( u1_u14_u3_n141 ) , .A1( u1_u14_u3_n169 ) );
  OAI222_X1 u1_u14_u3_U32 (.C2( u1_u14_u3_n107 ) , .A2( u1_u14_u3_n108 ) , .B1( u1_u14_u3_n135 ) , .ZN( u1_u14_u3_n138 ) , .B2( u1_u14_u3_n146 ) , .C1( u1_u14_u3_n154 ) , .A1( u1_u14_u3_n164 ) );
  NOR4_X1 u1_u14_u3_U33 (.A4( u1_u14_u3_n157 ) , .A3( u1_u14_u3_n158 ) , .A2( u1_u14_u3_n159 ) , .A1( u1_u14_u3_n160 ) , .ZN( u1_u14_u3_n161 ) );
  AOI21_X1 u1_u14_u3_U34 (.B2( u1_u14_u3_n152 ) , .B1( u1_u14_u3_n153 ) , .ZN( u1_u14_u3_n158 ) , .A( u1_u14_u3_n164 ) );
  AOI21_X1 u1_u14_u3_U35 (.A( u1_u14_u3_n154 ) , .B2( u1_u14_u3_n155 ) , .B1( u1_u14_u3_n156 ) , .ZN( u1_u14_u3_n157 ) );
  AOI21_X1 u1_u14_u3_U36 (.A( u1_u14_u3_n149 ) , .B2( u1_u14_u3_n150 ) , .B1( u1_u14_u3_n151 ) , .ZN( u1_u14_u3_n159 ) );
  AOI211_X1 u1_u14_u3_U37 (.ZN( u1_u14_u3_n109 ) , .A( u1_u14_u3_n119 ) , .C2( u1_u14_u3_n129 ) , .B( u1_u14_u3_n138 ) , .C1( u1_u14_u3_n141 ) );
  AOI211_X1 u1_u14_u3_U38 (.B( u1_u14_u3_n119 ) , .A( u1_u14_u3_n120 ) , .C2( u1_u14_u3_n121 ) , .ZN( u1_u14_u3_n122 ) , .C1( u1_u14_u3_n179 ) );
  INV_X1 u1_u14_u3_U39 (.A( u1_u14_u3_n156 ) , .ZN( u1_u14_u3_n179 ) );
  INV_X1 u1_u14_u3_U4 (.A( u1_u14_u3_n140 ) , .ZN( u1_u14_u3_n182 ) );
  OAI22_X1 u1_u14_u3_U40 (.B1( u1_u14_u3_n118 ) , .ZN( u1_u14_u3_n120 ) , .A1( u1_u14_u3_n135 ) , .B2( u1_u14_u3_n154 ) , .A2( u1_u14_u3_n178 ) );
  AND3_X1 u1_u14_u3_U41 (.ZN( u1_u14_u3_n118 ) , .A2( u1_u14_u3_n124 ) , .A1( u1_u14_u3_n144 ) , .A3( u1_u14_u3_n152 ) );
  INV_X1 u1_u14_u3_U42 (.A( u1_u14_u3_n121 ) , .ZN( u1_u14_u3_n164 ) );
  NAND2_X1 u1_u14_u3_U43 (.ZN( u1_u14_u3_n133 ) , .A1( u1_u14_u3_n154 ) , .A2( u1_u14_u3_n164 ) );
  OAI211_X1 u1_u14_u3_U44 (.B( u1_u14_u3_n127 ) , .ZN( u1_u14_u3_n139 ) , .C1( u1_u14_u3_n150 ) , .C2( u1_u14_u3_n154 ) , .A( u1_u14_u3_n184 ) );
  INV_X1 u1_u14_u3_U45 (.A( u1_u14_u3_n125 ) , .ZN( u1_u14_u3_n184 ) );
  AOI221_X1 u1_u14_u3_U46 (.A( u1_u14_u3_n126 ) , .ZN( u1_u14_u3_n127 ) , .C2( u1_u14_u3_n132 ) , .C1( u1_u14_u3_n169 ) , .B2( u1_u14_u3_n170 ) , .B1( u1_u14_u3_n174 ) );
  OAI22_X1 u1_u14_u3_U47 (.A1( u1_u14_u3_n124 ) , .ZN( u1_u14_u3_n125 ) , .B2( u1_u14_u3_n145 ) , .A2( u1_u14_u3_n165 ) , .B1( u1_u14_u3_n167 ) );
  NOR2_X1 u1_u14_u3_U48 (.A1( u1_u14_u3_n113 ) , .ZN( u1_u14_u3_n131 ) , .A2( u1_u14_u3_n154 ) );
  NAND2_X1 u1_u14_u3_U49 (.A1( u1_u14_u3_n103 ) , .ZN( u1_u14_u3_n150 ) , .A2( u1_u14_u3_n99 ) );
  INV_X1 u1_u14_u3_U5 (.A( u1_u14_u3_n117 ) , .ZN( u1_u14_u3_n178 ) );
  NAND2_X1 u1_u14_u3_U50 (.A2( u1_u14_u3_n102 ) , .ZN( u1_u14_u3_n155 ) , .A1( u1_u14_u3_n97 ) );
  INV_X1 u1_u14_u3_U51 (.A( u1_u14_u3_n141 ) , .ZN( u1_u14_u3_n167 ) );
  AOI21_X1 u1_u14_u3_U52 (.B2( u1_u14_u3_n114 ) , .B1( u1_u14_u3_n146 ) , .A( u1_u14_u3_n154 ) , .ZN( u1_u14_u3_n94 ) );
  AOI21_X1 u1_u14_u3_U53 (.ZN( u1_u14_u3_n110 ) , .B2( u1_u14_u3_n142 ) , .B1( u1_u14_u3_n186 ) , .A( u1_u14_u3_n95 ) );
  INV_X1 u1_u14_u3_U54 (.A( u1_u14_u3_n145 ) , .ZN( u1_u14_u3_n186 ) );
  AOI21_X1 u1_u14_u3_U55 (.B1( u1_u14_u3_n124 ) , .A( u1_u14_u3_n149 ) , .B2( u1_u14_u3_n155 ) , .ZN( u1_u14_u3_n95 ) );
  INV_X1 u1_u14_u3_U56 (.A( u1_u14_u3_n149 ) , .ZN( u1_u14_u3_n169 ) );
  NAND2_X1 u1_u14_u3_U57 (.ZN( u1_u14_u3_n124 ) , .A1( u1_u14_u3_n96 ) , .A2( u1_u14_u3_n97 ) );
  NAND2_X1 u1_u14_u3_U58 (.A2( u1_u14_u3_n100 ) , .ZN( u1_u14_u3_n146 ) , .A1( u1_u14_u3_n96 ) );
  NAND2_X1 u1_u14_u3_U59 (.A1( u1_u14_u3_n101 ) , .ZN( u1_u14_u3_n145 ) , .A2( u1_u14_u3_n99 ) );
  AOI221_X1 u1_u14_u3_U6 (.A( u1_u14_u3_n131 ) , .C2( u1_u14_u3_n132 ) , .C1( u1_u14_u3_n133 ) , .ZN( u1_u14_u3_n134 ) , .B1( u1_u14_u3_n143 ) , .B2( u1_u14_u3_n177 ) );
  NAND2_X1 u1_u14_u3_U60 (.A1( u1_u14_u3_n100 ) , .ZN( u1_u14_u3_n156 ) , .A2( u1_u14_u3_n99 ) );
  NAND2_X1 u1_u14_u3_U61 (.A2( u1_u14_u3_n101 ) , .A1( u1_u14_u3_n104 ) , .ZN( u1_u14_u3_n148 ) );
  NAND2_X1 u1_u14_u3_U62 (.A1( u1_u14_u3_n100 ) , .A2( u1_u14_u3_n102 ) , .ZN( u1_u14_u3_n128 ) );
  NAND2_X1 u1_u14_u3_U63 (.A2( u1_u14_u3_n101 ) , .A1( u1_u14_u3_n102 ) , .ZN( u1_u14_u3_n152 ) );
  NAND2_X1 u1_u14_u3_U64 (.A2( u1_u14_u3_n101 ) , .ZN( u1_u14_u3_n114 ) , .A1( u1_u14_u3_n96 ) );
  NAND2_X1 u1_u14_u3_U65 (.ZN( u1_u14_u3_n107 ) , .A1( u1_u14_u3_n97 ) , .A2( u1_u14_u3_n99 ) );
  NAND2_X1 u1_u14_u3_U66 (.A2( u1_u14_u3_n100 ) , .A1( u1_u14_u3_n104 ) , .ZN( u1_u14_u3_n113 ) );
  NAND2_X1 u1_u14_u3_U67 (.A1( u1_u14_u3_n104 ) , .ZN( u1_u14_u3_n153 ) , .A2( u1_u14_u3_n97 ) );
  NAND2_X1 u1_u14_u3_U68 (.A2( u1_u14_u3_n103 ) , .A1( u1_u14_u3_n104 ) , .ZN( u1_u14_u3_n130 ) );
  NAND2_X1 u1_u14_u3_U69 (.A2( u1_u14_u3_n103 ) , .ZN( u1_u14_u3_n144 ) , .A1( u1_u14_u3_n96 ) );
  OAI22_X1 u1_u14_u3_U7 (.B2( u1_u14_u3_n147 ) , .A2( u1_u14_u3_n148 ) , .ZN( u1_u14_u3_n160 ) , .B1( u1_u14_u3_n165 ) , .A1( u1_u14_u3_n168 ) );
  NAND2_X1 u1_u14_u3_U70 (.A1( u1_u14_u3_n102 ) , .A2( u1_u14_u3_n103 ) , .ZN( u1_u14_u3_n108 ) );
  NOR2_X1 u1_u14_u3_U71 (.A2( u1_u14_X_19 ) , .A1( u1_u14_X_20 ) , .ZN( u1_u14_u3_n99 ) );
  NOR2_X1 u1_u14_u3_U72 (.A2( u1_u14_X_21 ) , .A1( u1_u14_X_24 ) , .ZN( u1_u14_u3_n103 ) );
  NOR2_X1 u1_u14_u3_U73 (.A2( u1_u14_X_24 ) , .A1( u1_u14_u3_n171 ) , .ZN( u1_u14_u3_n97 ) );
  NOR2_X1 u1_u14_u3_U74 (.A2( u1_u14_X_23 ) , .ZN( u1_u14_u3_n141 ) , .A1( u1_u14_u3_n166 ) );
  NOR2_X1 u1_u14_u3_U75 (.A2( u1_u14_X_19 ) , .A1( u1_u14_u3_n172 ) , .ZN( u1_u14_u3_n96 ) );
  NAND2_X1 u1_u14_u3_U76 (.A1( u1_u14_X_22 ) , .A2( u1_u14_X_23 ) , .ZN( u1_u14_u3_n154 ) );
  NAND2_X1 u1_u14_u3_U77 (.A1( u1_u14_X_23 ) , .ZN( u1_u14_u3_n149 ) , .A2( u1_u14_u3_n166 ) );
  NOR2_X1 u1_u14_u3_U78 (.A2( u1_u14_X_22 ) , .A1( u1_u14_X_23 ) , .ZN( u1_u14_u3_n121 ) );
  AND2_X1 u1_u14_u3_U79 (.A1( u1_u14_X_24 ) , .ZN( u1_u14_u3_n101 ) , .A2( u1_u14_u3_n171 ) );
  AND3_X1 u1_u14_u3_U8 (.A3( u1_u14_u3_n144 ) , .A2( u1_u14_u3_n145 ) , .A1( u1_u14_u3_n146 ) , .ZN( u1_u14_u3_n147 ) );
  AND2_X1 u1_u14_u3_U80 (.A1( u1_u14_X_19 ) , .ZN( u1_u14_u3_n102 ) , .A2( u1_u14_u3_n172 ) );
  AND2_X1 u1_u14_u3_U81 (.A1( u1_u14_X_21 ) , .A2( u1_u14_X_24 ) , .ZN( u1_u14_u3_n100 ) );
  AND2_X1 u1_u14_u3_U82 (.A2( u1_u14_X_19 ) , .A1( u1_u14_X_20 ) , .ZN( u1_u14_u3_n104 ) );
  INV_X1 u1_u14_u3_U83 (.A( u1_u14_X_22 ) , .ZN( u1_u14_u3_n166 ) );
  INV_X1 u1_u14_u3_U84 (.A( u1_u14_X_21 ) , .ZN( u1_u14_u3_n171 ) );
  INV_X1 u1_u14_u3_U85 (.A( u1_u14_X_20 ) , .ZN( u1_u14_u3_n172 ) );
  NAND4_X1 u1_u14_u3_U86 (.ZN( u1_out14_26 ) , .A4( u1_u14_u3_n109 ) , .A3( u1_u14_u3_n110 ) , .A2( u1_u14_u3_n111 ) , .A1( u1_u14_u3_n173 ) );
  INV_X1 u1_u14_u3_U87 (.ZN( u1_u14_u3_n173 ) , .A( u1_u14_u3_n94 ) );
  OAI21_X1 u1_u14_u3_U88 (.ZN( u1_u14_u3_n111 ) , .B2( u1_u14_u3_n117 ) , .A( u1_u14_u3_n133 ) , .B1( u1_u14_u3_n176 ) );
  NAND4_X1 u1_u14_u3_U89 (.ZN( u1_out14_20 ) , .A4( u1_u14_u3_n122 ) , .A3( u1_u14_u3_n123 ) , .A1( u1_u14_u3_n175 ) , .A2( u1_u14_u3_n180 ) );
  INV_X1 u1_u14_u3_U9 (.A( u1_u14_u3_n143 ) , .ZN( u1_u14_u3_n168 ) );
  INV_X1 u1_u14_u3_U90 (.A( u1_u14_u3_n126 ) , .ZN( u1_u14_u3_n180 ) );
  INV_X1 u1_u14_u3_U91 (.A( u1_u14_u3_n112 ) , .ZN( u1_u14_u3_n175 ) );
  NAND4_X1 u1_u14_u3_U92 (.ZN( u1_out14_1 ) , .A4( u1_u14_u3_n161 ) , .A3( u1_u14_u3_n162 ) , .A2( u1_u14_u3_n163 ) , .A1( u1_u14_u3_n185 ) );
  NAND2_X1 u1_u14_u3_U93 (.ZN( u1_u14_u3_n163 ) , .A2( u1_u14_u3_n170 ) , .A1( u1_u14_u3_n176 ) );
  AOI22_X1 u1_u14_u3_U94 (.B2( u1_u14_u3_n140 ) , .B1( u1_u14_u3_n141 ) , .A2( u1_u14_u3_n142 ) , .ZN( u1_u14_u3_n162 ) , .A1( u1_u14_u3_n177 ) );
  OR4_X1 u1_u14_u3_U95 (.ZN( u1_out14_10 ) , .A4( u1_u14_u3_n136 ) , .A3( u1_u14_u3_n137 ) , .A1( u1_u14_u3_n138 ) , .A2( u1_u14_u3_n139 ) );
  OAI222_X1 u1_u14_u3_U96 (.C1( u1_u14_u3_n128 ) , .ZN( u1_u14_u3_n137 ) , .B1( u1_u14_u3_n148 ) , .A2( u1_u14_u3_n150 ) , .B2( u1_u14_u3_n154 ) , .C2( u1_u14_u3_n164 ) , .A1( u1_u14_u3_n167 ) );
  OAI221_X1 u1_u14_u3_U97 (.A( u1_u14_u3_n134 ) , .B2( u1_u14_u3_n135 ) , .ZN( u1_u14_u3_n136 ) , .C1( u1_u14_u3_n149 ) , .B1( u1_u14_u3_n151 ) , .C2( u1_u14_u3_n183 ) );
  NAND3_X1 u1_u14_u3_U98 (.A1( u1_u14_u3_n114 ) , .ZN( u1_u14_u3_n115 ) , .A2( u1_u14_u3_n145 ) , .A3( u1_u14_u3_n153 ) );
  NAND3_X1 u1_u14_u3_U99 (.ZN( u1_u14_u3_n129 ) , .A2( u1_u14_u3_n144 ) , .A1( u1_u14_u3_n153 ) , .A3( u1_u14_u3_n182 ) );
  XOR2_X1 u1_u15_U1 (.A( u1_FP_38 ) , .B( u1_K16_9 ) , .Z( u1_u15_X_9 ) );
  XOR2_X1 u1_u15_U16 (.A( u1_FP_34 ) , .B( u1_K16_3 ) , .Z( u1_u15_X_3 ) );
  XOR2_X1 u1_u15_U2 (.A( u1_FP_37 ) , .B( u1_K16_8 ) , .Z( u1_u15_X_8 ) );
  XOR2_X1 u1_u15_U4 (.A( u1_FP_37 ) , .B( u1_K16_6 ) , .Z( u1_u15_X_6 ) );
  XOR2_X1 u1_u15_U48 (.A( u1_FP_39 ) , .B( u1_K16_10 ) , .Z( u1_u15_X_10 ) );
  XOR2_X1 u1_u15_U6 (.A( u1_FP_35 ) , .B( u1_K16_4 ) , .Z( u1_u15_X_4 ) );
  AND3_X1 u1_u15_u0_U10 (.A2( u1_u15_u0_n112 ) , .ZN( u1_u15_u0_n127 ) , .A3( u1_u15_u0_n130 ) , .A1( u1_u15_u0_n148 ) );
  NAND2_X1 u1_u15_u0_U11 (.ZN( u1_u15_u0_n113 ) , .A1( u1_u15_u0_n139 ) , .A2( u1_u15_u0_n149 ) );
  AND2_X1 u1_u15_u0_U12 (.ZN( u1_u15_u0_n107 ) , .A1( u1_u15_u0_n130 ) , .A2( u1_u15_u0_n140 ) );
  AND2_X1 u1_u15_u0_U13 (.A2( u1_u15_u0_n129 ) , .A1( u1_u15_u0_n130 ) , .ZN( u1_u15_u0_n151 ) );
  AND2_X1 u1_u15_u0_U14 (.A1( u1_u15_u0_n108 ) , .A2( u1_u15_u0_n125 ) , .ZN( u1_u15_u0_n145 ) );
  INV_X1 u1_u15_u0_U15 (.A( u1_u15_u0_n143 ) , .ZN( u1_u15_u0_n173 ) );
  NOR2_X1 u1_u15_u0_U16 (.A2( u1_u15_u0_n136 ) , .ZN( u1_u15_u0_n147 ) , .A1( u1_u15_u0_n160 ) );
  AOI21_X1 u1_u15_u0_U17 (.B1( u1_u15_u0_n103 ) , .ZN( u1_u15_u0_n132 ) , .A( u1_u15_u0_n165 ) , .B2( u1_u15_u0_n93 ) );
  INV_X1 u1_u15_u0_U18 (.A( u1_u15_u0_n142 ) , .ZN( u1_u15_u0_n165 ) );
  OAI221_X1 u1_u15_u0_U19 (.C1( u1_u15_u0_n121 ) , .ZN( u1_u15_u0_n122 ) , .B2( u1_u15_u0_n127 ) , .A( u1_u15_u0_n143 ) , .B1( u1_u15_u0_n144 ) , .C2( u1_u15_u0_n147 ) );
  OAI22_X1 u1_u15_u0_U20 (.B1( u1_u15_u0_n131 ) , .A1( u1_u15_u0_n144 ) , .B2( u1_u15_u0_n147 ) , .A2( u1_u15_u0_n90 ) , .ZN( u1_u15_u0_n91 ) );
  AND3_X1 u1_u15_u0_U21 (.A3( u1_u15_u0_n121 ) , .A2( u1_u15_u0_n125 ) , .A1( u1_u15_u0_n148 ) , .ZN( u1_u15_u0_n90 ) );
  OAI22_X1 u1_u15_u0_U22 (.B1( u1_u15_u0_n125 ) , .ZN( u1_u15_u0_n126 ) , .A1( u1_u15_u0_n138 ) , .A2( u1_u15_u0_n146 ) , .B2( u1_u15_u0_n147 ) );
  NOR2_X1 u1_u15_u0_U23 (.A1( u1_u15_u0_n163 ) , .A2( u1_u15_u0_n164 ) , .ZN( u1_u15_u0_n95 ) );
  INV_X1 u1_u15_u0_U24 (.A( u1_u15_u0_n136 ) , .ZN( u1_u15_u0_n161 ) );
  NOR2_X1 u1_u15_u0_U25 (.A1( u1_u15_u0_n120 ) , .ZN( u1_u15_u0_n143 ) , .A2( u1_u15_u0_n167 ) );
  OAI221_X1 u1_u15_u0_U26 (.C1( u1_u15_u0_n112 ) , .ZN( u1_u15_u0_n120 ) , .B1( u1_u15_u0_n138 ) , .B2( u1_u15_u0_n141 ) , .C2( u1_u15_u0_n147 ) , .A( u1_u15_u0_n172 ) );
  AOI211_X1 u1_u15_u0_U27 (.B( u1_u15_u0_n115 ) , .A( u1_u15_u0_n116 ) , .C2( u1_u15_u0_n117 ) , .C1( u1_u15_u0_n118 ) , .ZN( u1_u15_u0_n119 ) );
  AOI22_X1 u1_u15_u0_U28 (.B2( u1_u15_u0_n109 ) , .A2( u1_u15_u0_n110 ) , .ZN( u1_u15_u0_n111 ) , .B1( u1_u15_u0_n118 ) , .A1( u1_u15_u0_n160 ) );
  NAND2_X1 u1_u15_u0_U29 (.A2( u1_u15_u0_n102 ) , .A1( u1_u15_u0_n103 ) , .ZN( u1_u15_u0_n149 ) );
  INV_X1 u1_u15_u0_U3 (.A( u1_u15_u0_n113 ) , .ZN( u1_u15_u0_n166 ) );
  INV_X1 u1_u15_u0_U30 (.A( u1_u15_u0_n118 ) , .ZN( u1_u15_u0_n158 ) );
  NAND2_X1 u1_u15_u0_U31 (.A2( u1_u15_u0_n100 ) , .ZN( u1_u15_u0_n131 ) , .A1( u1_u15_u0_n92 ) );
  NAND2_X1 u1_u15_u0_U32 (.ZN( u1_u15_u0_n108 ) , .A1( u1_u15_u0_n92 ) , .A2( u1_u15_u0_n94 ) );
  AOI21_X1 u1_u15_u0_U33 (.ZN( u1_u15_u0_n104 ) , .B1( u1_u15_u0_n107 ) , .B2( u1_u15_u0_n141 ) , .A( u1_u15_u0_n144 ) );
  AOI21_X1 u1_u15_u0_U34 (.B1( u1_u15_u0_n127 ) , .B2( u1_u15_u0_n129 ) , .A( u1_u15_u0_n138 ) , .ZN( u1_u15_u0_n96 ) );
  NAND2_X1 u1_u15_u0_U35 (.A2( u1_u15_u0_n102 ) , .ZN( u1_u15_u0_n114 ) , .A1( u1_u15_u0_n92 ) );
  AOI21_X1 u1_u15_u0_U36 (.ZN( u1_u15_u0_n116 ) , .B2( u1_u15_u0_n142 ) , .A( u1_u15_u0_n144 ) , .B1( u1_u15_u0_n166 ) );
  NAND2_X1 u1_u15_u0_U37 (.A2( u1_u15_u0_n103 ) , .ZN( u1_u15_u0_n140 ) , .A1( u1_u15_u0_n94 ) );
  NAND2_X1 u1_u15_u0_U38 (.A1( u1_u15_u0_n100 ) , .A2( u1_u15_u0_n103 ) , .ZN( u1_u15_u0_n125 ) );
  NAND2_X1 u1_u15_u0_U39 (.A1( u1_u15_u0_n101 ) , .A2( u1_u15_u0_n102 ) , .ZN( u1_u15_u0_n150 ) );
  AOI21_X1 u1_u15_u0_U4 (.B1( u1_u15_u0_n114 ) , .ZN( u1_u15_u0_n115 ) , .B2( u1_u15_u0_n129 ) , .A( u1_u15_u0_n161 ) );
  INV_X1 u1_u15_u0_U40 (.A( u1_u15_u0_n138 ) , .ZN( u1_u15_u0_n160 ) );
  NAND2_X1 u1_u15_u0_U41 (.A2( u1_u15_u0_n100 ) , .A1( u1_u15_u0_n101 ) , .ZN( u1_u15_u0_n139 ) );
  NAND2_X1 u1_u15_u0_U42 (.ZN( u1_u15_u0_n112 ) , .A2( u1_u15_u0_n92 ) , .A1( u1_u15_u0_n93 ) );
  NAND2_X1 u1_u15_u0_U43 (.A1( u1_u15_u0_n101 ) , .ZN( u1_u15_u0_n130 ) , .A2( u1_u15_u0_n94 ) );
  NAND2_X1 u1_u15_u0_U44 (.A2( u1_u15_u0_n101 ) , .ZN( u1_u15_u0_n121 ) , .A1( u1_u15_u0_n93 ) );
  INV_X1 u1_u15_u0_U45 (.ZN( u1_u15_u0_n172 ) , .A( u1_u15_u0_n88 ) );
  OAI222_X1 u1_u15_u0_U46 (.C1( u1_u15_u0_n108 ) , .A1( u1_u15_u0_n125 ) , .B2( u1_u15_u0_n128 ) , .B1( u1_u15_u0_n144 ) , .A2( u1_u15_u0_n158 ) , .C2( u1_u15_u0_n161 ) , .ZN( u1_u15_u0_n88 ) );
  OR3_X1 u1_u15_u0_U47 (.A3( u1_u15_u0_n152 ) , .A2( u1_u15_u0_n153 ) , .A1( u1_u15_u0_n154 ) , .ZN( u1_u15_u0_n155 ) );
  AOI21_X1 u1_u15_u0_U48 (.B2( u1_u15_u0_n150 ) , .B1( u1_u15_u0_n151 ) , .ZN( u1_u15_u0_n152 ) , .A( u1_u15_u0_n158 ) );
  AOI21_X1 u1_u15_u0_U49 (.A( u1_u15_u0_n144 ) , .B2( u1_u15_u0_n145 ) , .B1( u1_u15_u0_n146 ) , .ZN( u1_u15_u0_n154 ) );
  AOI21_X1 u1_u15_u0_U5 (.B2( u1_u15_u0_n131 ) , .ZN( u1_u15_u0_n134 ) , .B1( u1_u15_u0_n151 ) , .A( u1_u15_u0_n158 ) );
  AOI21_X1 u1_u15_u0_U50 (.A( u1_u15_u0_n147 ) , .B2( u1_u15_u0_n148 ) , .B1( u1_u15_u0_n149 ) , .ZN( u1_u15_u0_n153 ) );
  INV_X1 u1_u15_u0_U51 (.ZN( u1_u15_u0_n171 ) , .A( u1_u15_u0_n99 ) );
  OAI211_X1 u1_u15_u0_U52 (.C2( u1_u15_u0_n140 ) , .C1( u1_u15_u0_n161 ) , .A( u1_u15_u0_n169 ) , .B( u1_u15_u0_n98 ) , .ZN( u1_u15_u0_n99 ) );
  AOI211_X1 u1_u15_u0_U53 (.C1( u1_u15_u0_n118 ) , .A( u1_u15_u0_n123 ) , .B( u1_u15_u0_n96 ) , .C2( u1_u15_u0_n97 ) , .ZN( u1_u15_u0_n98 ) );
  INV_X1 u1_u15_u0_U54 (.ZN( u1_u15_u0_n169 ) , .A( u1_u15_u0_n91 ) );
  NOR2_X1 u1_u15_u0_U55 (.A2( u1_u15_X_4 ) , .A1( u1_u15_X_5 ) , .ZN( u1_u15_u0_n118 ) );
  NOR2_X1 u1_u15_u0_U56 (.A2( u1_u15_X_1 ) , .ZN( u1_u15_u0_n101 ) , .A1( u1_u15_u0_n163 ) );
  NOR2_X1 u1_u15_u0_U57 (.A2( u1_u15_X_3 ) , .A1( u1_u15_X_6 ) , .ZN( u1_u15_u0_n94 ) );
  NOR2_X1 u1_u15_u0_U58 (.A2( u1_u15_X_6 ) , .ZN( u1_u15_u0_n100 ) , .A1( u1_u15_u0_n162 ) );
  NAND2_X1 u1_u15_u0_U59 (.A2( u1_u15_X_4 ) , .A1( u1_u15_X_5 ) , .ZN( u1_u15_u0_n144 ) );
  NOR2_X1 u1_u15_u0_U6 (.A1( u1_u15_u0_n108 ) , .ZN( u1_u15_u0_n123 ) , .A2( u1_u15_u0_n158 ) );
  NOR2_X1 u1_u15_u0_U60 (.A2( u1_u15_X_5 ) , .ZN( u1_u15_u0_n136 ) , .A1( u1_u15_u0_n159 ) );
  NAND2_X1 u1_u15_u0_U61 (.A1( u1_u15_X_5 ) , .ZN( u1_u15_u0_n138 ) , .A2( u1_u15_u0_n159 ) );
  AND2_X1 u1_u15_u0_U62 (.A2( u1_u15_X_3 ) , .A1( u1_u15_X_6 ) , .ZN( u1_u15_u0_n102 ) );
  AND2_X1 u1_u15_u0_U63 (.A1( u1_u15_X_6 ) , .A2( u1_u15_u0_n162 ) , .ZN( u1_u15_u0_n93 ) );
  INV_X1 u1_u15_u0_U64 (.A( u1_u15_X_4 ) , .ZN( u1_u15_u0_n159 ) );
  INV_X1 u1_u15_u0_U65 (.A( u1_u15_X_1 ) , .ZN( u1_u15_u0_n164 ) );
  INV_X1 u1_u15_u0_U66 (.A( u1_u15_X_3 ) , .ZN( u1_u15_u0_n162 ) );
  INV_X1 u1_u15_u0_U67 (.A( u1_u15_u0_n126 ) , .ZN( u1_u15_u0_n168 ) );
  AOI211_X1 u1_u15_u0_U68 (.B( u1_u15_u0_n133 ) , .A( u1_u15_u0_n134 ) , .C2( u1_u15_u0_n135 ) , .C1( u1_u15_u0_n136 ) , .ZN( u1_u15_u0_n137 ) );
  INV_X1 u1_u15_u0_U69 (.ZN( u1_u15_u0_n174 ) , .A( u1_u15_u0_n89 ) );
  OAI21_X1 u1_u15_u0_U7 (.B1( u1_u15_u0_n150 ) , .B2( u1_u15_u0_n158 ) , .A( u1_u15_u0_n172 ) , .ZN( u1_u15_u0_n89 ) );
  AOI211_X1 u1_u15_u0_U70 (.B( u1_u15_u0_n104 ) , .A( u1_u15_u0_n105 ) , .ZN( u1_u15_u0_n106 ) , .C2( u1_u15_u0_n113 ) , .C1( u1_u15_u0_n160 ) );
  OR4_X1 u1_u15_u0_U71 (.ZN( u1_out15_17 ) , .A4( u1_u15_u0_n122 ) , .A2( u1_u15_u0_n123 ) , .A1( u1_u15_u0_n124 ) , .A3( u1_u15_u0_n170 ) );
  AOI21_X1 u1_u15_u0_U72 (.B2( u1_u15_u0_n107 ) , .ZN( u1_u15_u0_n124 ) , .B1( u1_u15_u0_n128 ) , .A( u1_u15_u0_n161 ) );
  INV_X1 u1_u15_u0_U73 (.A( u1_u15_u0_n111 ) , .ZN( u1_u15_u0_n170 ) );
  OR4_X1 u1_u15_u0_U74 (.ZN( u1_out15_31 ) , .A4( u1_u15_u0_n155 ) , .A2( u1_u15_u0_n156 ) , .A1( u1_u15_u0_n157 ) , .A3( u1_u15_u0_n173 ) );
  AOI21_X1 u1_u15_u0_U75 (.A( u1_u15_u0_n138 ) , .B2( u1_u15_u0_n139 ) , .B1( u1_u15_u0_n140 ) , .ZN( u1_u15_u0_n157 ) );
  AOI21_X1 u1_u15_u0_U76 (.B2( u1_u15_u0_n141 ) , .B1( u1_u15_u0_n142 ) , .ZN( u1_u15_u0_n156 ) , .A( u1_u15_u0_n161 ) );
  AOI21_X1 u1_u15_u0_U77 (.B1( u1_u15_u0_n132 ) , .ZN( u1_u15_u0_n133 ) , .A( u1_u15_u0_n144 ) , .B2( u1_u15_u0_n166 ) );
  OAI22_X1 u1_u15_u0_U78 (.ZN( u1_u15_u0_n105 ) , .A2( u1_u15_u0_n132 ) , .B1( u1_u15_u0_n146 ) , .A1( u1_u15_u0_n147 ) , .B2( u1_u15_u0_n161 ) );
  NAND2_X1 u1_u15_u0_U79 (.ZN( u1_u15_u0_n110 ) , .A2( u1_u15_u0_n132 ) , .A1( u1_u15_u0_n145 ) );
  AND2_X1 u1_u15_u0_U8 (.A1( u1_u15_u0_n114 ) , .A2( u1_u15_u0_n121 ) , .ZN( u1_u15_u0_n146 ) );
  INV_X1 u1_u15_u0_U80 (.A( u1_u15_u0_n119 ) , .ZN( u1_u15_u0_n167 ) );
  NAND2_X1 u1_u15_u0_U81 (.ZN( u1_u15_u0_n148 ) , .A1( u1_u15_u0_n93 ) , .A2( u1_u15_u0_n95 ) );
  NAND2_X1 u1_u15_u0_U82 (.A1( u1_u15_u0_n100 ) , .ZN( u1_u15_u0_n129 ) , .A2( u1_u15_u0_n95 ) );
  NAND2_X1 u1_u15_u0_U83 (.A1( u1_u15_u0_n102 ) , .ZN( u1_u15_u0_n128 ) , .A2( u1_u15_u0_n95 ) );
  NOR2_X1 u1_u15_u0_U84 (.A2( u1_u15_X_1 ) , .A1( u1_u15_X_2 ) , .ZN( u1_u15_u0_n92 ) );
  NAND2_X1 u1_u15_u0_U85 (.ZN( u1_u15_u0_n142 ) , .A1( u1_u15_u0_n94 ) , .A2( u1_u15_u0_n95 ) );
  NOR2_X1 u1_u15_u0_U86 (.A2( u1_u15_X_2 ) , .ZN( u1_u15_u0_n103 ) , .A1( u1_u15_u0_n164 ) );
  INV_X1 u1_u15_u0_U87 (.A( u1_u15_X_2 ) , .ZN( u1_u15_u0_n163 ) );
  NAND3_X1 u1_u15_u0_U88 (.ZN( u1_out15_23 ) , .A3( u1_u15_u0_n137 ) , .A1( u1_u15_u0_n168 ) , .A2( u1_u15_u0_n171 ) );
  NAND3_X1 u1_u15_u0_U89 (.A3( u1_u15_u0_n127 ) , .A2( u1_u15_u0_n128 ) , .ZN( u1_u15_u0_n135 ) , .A1( u1_u15_u0_n150 ) );
  AND2_X1 u1_u15_u0_U9 (.A1( u1_u15_u0_n131 ) , .ZN( u1_u15_u0_n141 ) , .A2( u1_u15_u0_n150 ) );
  NAND3_X1 u1_u15_u0_U90 (.ZN( u1_u15_u0_n117 ) , .A3( u1_u15_u0_n132 ) , .A2( u1_u15_u0_n139 ) , .A1( u1_u15_u0_n148 ) );
  NAND3_X1 u1_u15_u0_U91 (.ZN( u1_u15_u0_n109 ) , .A2( u1_u15_u0_n114 ) , .A3( u1_u15_u0_n140 ) , .A1( u1_u15_u0_n149 ) );
  NAND3_X1 u1_u15_u0_U92 (.ZN( u1_out15_9 ) , .A3( u1_u15_u0_n106 ) , .A2( u1_u15_u0_n171 ) , .A1( u1_u15_u0_n174 ) );
  NAND3_X1 u1_u15_u0_U93 (.A2( u1_u15_u0_n128 ) , .A1( u1_u15_u0_n132 ) , .A3( u1_u15_u0_n146 ) , .ZN( u1_u15_u0_n97 ) );
  AOI21_X1 u1_u15_u1_U10 (.B2( u1_u15_u1_n155 ) , .B1( u1_u15_u1_n156 ) , .ZN( u1_u15_u1_n157 ) , .A( u1_u15_u1_n174 ) );
  NAND3_X1 u1_u15_u1_U100 (.ZN( u1_u15_u1_n113 ) , .A1( u1_u15_u1_n120 ) , .A3( u1_u15_u1_n133 ) , .A2( u1_u15_u1_n155 ) );
  NAND2_X1 u1_u15_u1_U11 (.ZN( u1_u15_u1_n140 ) , .A2( u1_u15_u1_n150 ) , .A1( u1_u15_u1_n155 ) );
  NAND2_X1 u1_u15_u1_U12 (.A1( u1_u15_u1_n131 ) , .ZN( u1_u15_u1_n147 ) , .A2( u1_u15_u1_n153 ) );
  INV_X1 u1_u15_u1_U13 (.A( u1_u15_u1_n139 ) , .ZN( u1_u15_u1_n174 ) );
  OR4_X1 u1_u15_u1_U14 (.A4( u1_u15_u1_n106 ) , .A3( u1_u15_u1_n107 ) , .ZN( u1_u15_u1_n108 ) , .A1( u1_u15_u1_n117 ) , .A2( u1_u15_u1_n184 ) );
  AOI21_X1 u1_u15_u1_U15 (.ZN( u1_u15_u1_n106 ) , .A( u1_u15_u1_n112 ) , .B1( u1_u15_u1_n154 ) , .B2( u1_u15_u1_n156 ) );
  AOI21_X1 u1_u15_u1_U16 (.ZN( u1_u15_u1_n107 ) , .B1( u1_u15_u1_n134 ) , .B2( u1_u15_u1_n149 ) , .A( u1_u15_u1_n174 ) );
  INV_X1 u1_u15_u1_U17 (.A( u1_u15_u1_n101 ) , .ZN( u1_u15_u1_n184 ) );
  INV_X1 u1_u15_u1_U18 (.A( u1_u15_u1_n112 ) , .ZN( u1_u15_u1_n171 ) );
  NAND2_X1 u1_u15_u1_U19 (.ZN( u1_u15_u1_n141 ) , .A1( u1_u15_u1_n153 ) , .A2( u1_u15_u1_n156 ) );
  AND2_X1 u1_u15_u1_U20 (.A1( u1_u15_u1_n123 ) , .ZN( u1_u15_u1_n134 ) , .A2( u1_u15_u1_n161 ) );
  NAND2_X1 u1_u15_u1_U21 (.A2( u1_u15_u1_n115 ) , .A1( u1_u15_u1_n116 ) , .ZN( u1_u15_u1_n148 ) );
  NAND2_X1 u1_u15_u1_U22 (.A2( u1_u15_u1_n133 ) , .A1( u1_u15_u1_n135 ) , .ZN( u1_u15_u1_n159 ) );
  NAND2_X1 u1_u15_u1_U23 (.A2( u1_u15_u1_n115 ) , .A1( u1_u15_u1_n120 ) , .ZN( u1_u15_u1_n132 ) );
  INV_X1 u1_u15_u1_U24 (.A( u1_u15_u1_n154 ) , .ZN( u1_u15_u1_n178 ) );
  AOI22_X1 u1_u15_u1_U25 (.B2( u1_u15_u1_n113 ) , .A2( u1_u15_u1_n114 ) , .ZN( u1_u15_u1_n125 ) , .A1( u1_u15_u1_n171 ) , .B1( u1_u15_u1_n173 ) );
  NAND2_X1 u1_u15_u1_U26 (.ZN( u1_u15_u1_n114 ) , .A1( u1_u15_u1_n134 ) , .A2( u1_u15_u1_n156 ) );
  INV_X1 u1_u15_u1_U27 (.A( u1_u15_u1_n151 ) , .ZN( u1_u15_u1_n183 ) );
  AND2_X1 u1_u15_u1_U28 (.A1( u1_u15_u1_n129 ) , .A2( u1_u15_u1_n133 ) , .ZN( u1_u15_u1_n149 ) );
  INV_X1 u1_u15_u1_U29 (.A( u1_u15_u1_n131 ) , .ZN( u1_u15_u1_n180 ) );
  INV_X1 u1_u15_u1_U3 (.A( u1_u15_u1_n159 ) , .ZN( u1_u15_u1_n182 ) );
  OAI221_X1 u1_u15_u1_U30 (.A( u1_u15_u1_n119 ) , .C2( u1_u15_u1_n129 ) , .ZN( u1_u15_u1_n138 ) , .B2( u1_u15_u1_n152 ) , .C1( u1_u15_u1_n174 ) , .B1( u1_u15_u1_n187 ) );
  INV_X1 u1_u15_u1_U31 (.A( u1_u15_u1_n148 ) , .ZN( u1_u15_u1_n187 ) );
  AOI211_X1 u1_u15_u1_U32 (.B( u1_u15_u1_n117 ) , .A( u1_u15_u1_n118 ) , .ZN( u1_u15_u1_n119 ) , .C2( u1_u15_u1_n146 ) , .C1( u1_u15_u1_n159 ) );
  NOR2_X1 u1_u15_u1_U33 (.A1( u1_u15_u1_n168 ) , .A2( u1_u15_u1_n176 ) , .ZN( u1_u15_u1_n98 ) );
  AOI211_X1 u1_u15_u1_U34 (.B( u1_u15_u1_n162 ) , .A( u1_u15_u1_n163 ) , .C2( u1_u15_u1_n164 ) , .ZN( u1_u15_u1_n165 ) , .C1( u1_u15_u1_n171 ) );
  AOI21_X1 u1_u15_u1_U35 (.A( u1_u15_u1_n160 ) , .B2( u1_u15_u1_n161 ) , .ZN( u1_u15_u1_n162 ) , .B1( u1_u15_u1_n182 ) );
  OR2_X1 u1_u15_u1_U36 (.A2( u1_u15_u1_n157 ) , .A1( u1_u15_u1_n158 ) , .ZN( u1_u15_u1_n163 ) );
  NAND2_X1 u1_u15_u1_U37 (.A1( u1_u15_u1_n128 ) , .ZN( u1_u15_u1_n146 ) , .A2( u1_u15_u1_n160 ) );
  NAND2_X1 u1_u15_u1_U38 (.A2( u1_u15_u1_n112 ) , .ZN( u1_u15_u1_n139 ) , .A1( u1_u15_u1_n152 ) );
  NAND2_X1 u1_u15_u1_U39 (.A1( u1_u15_u1_n105 ) , .ZN( u1_u15_u1_n156 ) , .A2( u1_u15_u1_n99 ) );
  AOI221_X1 u1_u15_u1_U4 (.A( u1_u15_u1_n138 ) , .C2( u1_u15_u1_n139 ) , .C1( u1_u15_u1_n140 ) , .B2( u1_u15_u1_n141 ) , .ZN( u1_u15_u1_n142 ) , .B1( u1_u15_u1_n175 ) );
  AOI221_X1 u1_u15_u1_U40 (.B1( u1_u15_u1_n140 ) , .ZN( u1_u15_u1_n167 ) , .B2( u1_u15_u1_n172 ) , .C2( u1_u15_u1_n175 ) , .C1( u1_u15_u1_n178 ) , .A( u1_u15_u1_n188 ) );
  INV_X1 u1_u15_u1_U41 (.ZN( u1_u15_u1_n188 ) , .A( u1_u15_u1_n97 ) );
  AOI211_X1 u1_u15_u1_U42 (.A( u1_u15_u1_n118 ) , .C1( u1_u15_u1_n132 ) , .C2( u1_u15_u1_n139 ) , .B( u1_u15_u1_n96 ) , .ZN( u1_u15_u1_n97 ) );
  AOI21_X1 u1_u15_u1_U43 (.B2( u1_u15_u1_n121 ) , .B1( u1_u15_u1_n135 ) , .A( u1_u15_u1_n152 ) , .ZN( u1_u15_u1_n96 ) );
  NOR2_X1 u1_u15_u1_U44 (.ZN( u1_u15_u1_n117 ) , .A1( u1_u15_u1_n121 ) , .A2( u1_u15_u1_n160 ) );
  AOI21_X1 u1_u15_u1_U45 (.A( u1_u15_u1_n128 ) , .B2( u1_u15_u1_n129 ) , .ZN( u1_u15_u1_n130 ) , .B1( u1_u15_u1_n150 ) );
  OAI21_X1 u1_u15_u1_U46 (.B2( u1_u15_u1_n123 ) , .ZN( u1_u15_u1_n145 ) , .B1( u1_u15_u1_n160 ) , .A( u1_u15_u1_n185 ) );
  INV_X1 u1_u15_u1_U47 (.A( u1_u15_u1_n122 ) , .ZN( u1_u15_u1_n185 ) );
  AOI21_X1 u1_u15_u1_U48 (.B2( u1_u15_u1_n120 ) , .B1( u1_u15_u1_n121 ) , .ZN( u1_u15_u1_n122 ) , .A( u1_u15_u1_n128 ) );
  NAND2_X1 u1_u15_u1_U49 (.ZN( u1_u15_u1_n112 ) , .A1( u1_u15_u1_n169 ) , .A2( u1_u15_u1_n170 ) );
  AOI211_X1 u1_u15_u1_U5 (.ZN( u1_u15_u1_n124 ) , .A( u1_u15_u1_n138 ) , .C2( u1_u15_u1_n139 ) , .B( u1_u15_u1_n145 ) , .C1( u1_u15_u1_n147 ) );
  NAND2_X1 u1_u15_u1_U50 (.ZN( u1_u15_u1_n129 ) , .A2( u1_u15_u1_n95 ) , .A1( u1_u15_u1_n98 ) );
  NAND2_X1 u1_u15_u1_U51 (.A1( u1_u15_u1_n102 ) , .ZN( u1_u15_u1_n154 ) , .A2( u1_u15_u1_n99 ) );
  NAND2_X1 u1_u15_u1_U52 (.A2( u1_u15_u1_n100 ) , .ZN( u1_u15_u1_n135 ) , .A1( u1_u15_u1_n99 ) );
  AOI21_X1 u1_u15_u1_U53 (.A( u1_u15_u1_n152 ) , .B2( u1_u15_u1_n153 ) , .B1( u1_u15_u1_n154 ) , .ZN( u1_u15_u1_n158 ) );
  INV_X1 u1_u15_u1_U54 (.A( u1_u15_u1_n160 ) , .ZN( u1_u15_u1_n175 ) );
  NAND2_X1 u1_u15_u1_U55 (.A1( u1_u15_u1_n100 ) , .ZN( u1_u15_u1_n116 ) , .A2( u1_u15_u1_n95 ) );
  NAND2_X1 u1_u15_u1_U56 (.A1( u1_u15_u1_n102 ) , .ZN( u1_u15_u1_n131 ) , .A2( u1_u15_u1_n95 ) );
  NAND2_X1 u1_u15_u1_U57 (.A2( u1_u15_u1_n104 ) , .ZN( u1_u15_u1_n121 ) , .A1( u1_u15_u1_n98 ) );
  NAND2_X1 u1_u15_u1_U58 (.A1( u1_u15_u1_n103 ) , .ZN( u1_u15_u1_n153 ) , .A2( u1_u15_u1_n98 ) );
  NAND2_X1 u1_u15_u1_U59 (.A2( u1_u15_u1_n104 ) , .A1( u1_u15_u1_n105 ) , .ZN( u1_u15_u1_n133 ) );
  AOI22_X1 u1_u15_u1_U6 (.B2( u1_u15_u1_n136 ) , .A2( u1_u15_u1_n137 ) , .ZN( u1_u15_u1_n143 ) , .A1( u1_u15_u1_n171 ) , .B1( u1_u15_u1_n173 ) );
  NAND2_X1 u1_u15_u1_U60 (.ZN( u1_u15_u1_n150 ) , .A2( u1_u15_u1_n98 ) , .A1( u1_u15_u1_n99 ) );
  NAND2_X1 u1_u15_u1_U61 (.A1( u1_u15_u1_n105 ) , .ZN( u1_u15_u1_n155 ) , .A2( u1_u15_u1_n95 ) );
  OAI21_X1 u1_u15_u1_U62 (.ZN( u1_u15_u1_n109 ) , .B1( u1_u15_u1_n129 ) , .B2( u1_u15_u1_n160 ) , .A( u1_u15_u1_n167 ) );
  NAND2_X1 u1_u15_u1_U63 (.A2( u1_u15_u1_n100 ) , .A1( u1_u15_u1_n103 ) , .ZN( u1_u15_u1_n120 ) );
  NAND2_X1 u1_u15_u1_U64 (.A1( u1_u15_u1_n102 ) , .A2( u1_u15_u1_n104 ) , .ZN( u1_u15_u1_n115 ) );
  NAND2_X1 u1_u15_u1_U65 (.A2( u1_u15_u1_n100 ) , .A1( u1_u15_u1_n104 ) , .ZN( u1_u15_u1_n151 ) );
  NAND2_X1 u1_u15_u1_U66 (.A2( u1_u15_u1_n103 ) , .A1( u1_u15_u1_n105 ) , .ZN( u1_u15_u1_n161 ) );
  INV_X1 u1_u15_u1_U67 (.A( u1_u15_u1_n152 ) , .ZN( u1_u15_u1_n173 ) );
  INV_X1 u1_u15_u1_U68 (.A( u1_u15_u1_n128 ) , .ZN( u1_u15_u1_n172 ) );
  NAND2_X1 u1_u15_u1_U69 (.A2( u1_u15_u1_n102 ) , .A1( u1_u15_u1_n103 ) , .ZN( u1_u15_u1_n123 ) );
  INV_X1 u1_u15_u1_U7 (.A( u1_u15_u1_n147 ) , .ZN( u1_u15_u1_n181 ) );
  NOR2_X1 u1_u15_u1_U70 (.A2( u1_u15_X_7 ) , .A1( u1_u15_X_8 ) , .ZN( u1_u15_u1_n95 ) );
  NOR2_X1 u1_u15_u1_U71 (.A1( u1_u15_X_12 ) , .A2( u1_u15_X_9 ) , .ZN( u1_u15_u1_n100 ) );
  NOR2_X1 u1_u15_u1_U72 (.A2( u1_u15_X_8 ) , .A1( u1_u15_u1_n177 ) , .ZN( u1_u15_u1_n99 ) );
  NOR2_X1 u1_u15_u1_U73 (.A2( u1_u15_X_12 ) , .ZN( u1_u15_u1_n102 ) , .A1( u1_u15_u1_n176 ) );
  NOR2_X1 u1_u15_u1_U74 (.A2( u1_u15_X_9 ) , .ZN( u1_u15_u1_n105 ) , .A1( u1_u15_u1_n168 ) );
  NAND2_X1 u1_u15_u1_U75 (.A1( u1_u15_X_10 ) , .ZN( u1_u15_u1_n160 ) , .A2( u1_u15_u1_n169 ) );
  NAND2_X1 u1_u15_u1_U76 (.A2( u1_u15_X_10 ) , .A1( u1_u15_X_11 ) , .ZN( u1_u15_u1_n152 ) );
  NAND2_X1 u1_u15_u1_U77 (.A1( u1_u15_X_11 ) , .ZN( u1_u15_u1_n128 ) , .A2( u1_u15_u1_n170 ) );
  AND2_X1 u1_u15_u1_U78 (.A2( u1_u15_X_7 ) , .A1( u1_u15_X_8 ) , .ZN( u1_u15_u1_n104 ) );
  AND2_X1 u1_u15_u1_U79 (.A1( u1_u15_X_8 ) , .ZN( u1_u15_u1_n103 ) , .A2( u1_u15_u1_n177 ) );
  NOR2_X1 u1_u15_u1_U8 (.A1( u1_u15_u1_n112 ) , .A2( u1_u15_u1_n116 ) , .ZN( u1_u15_u1_n118 ) );
  INV_X1 u1_u15_u1_U80 (.A( u1_u15_X_10 ) , .ZN( u1_u15_u1_n170 ) );
  INV_X1 u1_u15_u1_U81 (.A( u1_u15_X_9 ) , .ZN( u1_u15_u1_n176 ) );
  INV_X1 u1_u15_u1_U82 (.A( u1_u15_X_11 ) , .ZN( u1_u15_u1_n169 ) );
  INV_X1 u1_u15_u1_U83 (.A( u1_u15_X_12 ) , .ZN( u1_u15_u1_n168 ) );
  INV_X1 u1_u15_u1_U84 (.A( u1_u15_X_7 ) , .ZN( u1_u15_u1_n177 ) );
  NAND4_X1 u1_u15_u1_U85 (.ZN( u1_out15_18 ) , .A4( u1_u15_u1_n165 ) , .A3( u1_u15_u1_n166 ) , .A1( u1_u15_u1_n167 ) , .A2( u1_u15_u1_n186 ) );
  AOI22_X1 u1_u15_u1_U86 (.B2( u1_u15_u1_n146 ) , .B1( u1_u15_u1_n147 ) , .A2( u1_u15_u1_n148 ) , .ZN( u1_u15_u1_n166 ) , .A1( u1_u15_u1_n172 ) );
  INV_X1 u1_u15_u1_U87 (.A( u1_u15_u1_n145 ) , .ZN( u1_u15_u1_n186 ) );
  NAND4_X1 u1_u15_u1_U88 (.ZN( u1_out15_2 ) , .A4( u1_u15_u1_n142 ) , .A3( u1_u15_u1_n143 ) , .A2( u1_u15_u1_n144 ) , .A1( u1_u15_u1_n179 ) );
  OAI21_X1 u1_u15_u1_U89 (.B2( u1_u15_u1_n132 ) , .ZN( u1_u15_u1_n144 ) , .A( u1_u15_u1_n146 ) , .B1( u1_u15_u1_n180 ) );
  OAI21_X1 u1_u15_u1_U9 (.ZN( u1_u15_u1_n101 ) , .B1( u1_u15_u1_n141 ) , .A( u1_u15_u1_n146 ) , .B2( u1_u15_u1_n183 ) );
  INV_X1 u1_u15_u1_U90 (.A( u1_u15_u1_n130 ) , .ZN( u1_u15_u1_n179 ) );
  NAND4_X1 u1_u15_u1_U91 (.ZN( u1_out15_28 ) , .A4( u1_u15_u1_n124 ) , .A3( u1_u15_u1_n125 ) , .A2( u1_u15_u1_n126 ) , .A1( u1_u15_u1_n127 ) );
  OAI21_X1 u1_u15_u1_U92 (.ZN( u1_u15_u1_n127 ) , .B2( u1_u15_u1_n139 ) , .B1( u1_u15_u1_n175 ) , .A( u1_u15_u1_n183 ) );
  OAI21_X1 u1_u15_u1_U93 (.ZN( u1_u15_u1_n126 ) , .B2( u1_u15_u1_n140 ) , .A( u1_u15_u1_n146 ) , .B1( u1_u15_u1_n178 ) );
  OR4_X1 u1_u15_u1_U94 (.ZN( u1_out15_13 ) , .A4( u1_u15_u1_n108 ) , .A3( u1_u15_u1_n109 ) , .A2( u1_u15_u1_n110 ) , .A1( u1_u15_u1_n111 ) );
  AOI21_X1 u1_u15_u1_U95 (.ZN( u1_u15_u1_n111 ) , .A( u1_u15_u1_n128 ) , .B2( u1_u15_u1_n131 ) , .B1( u1_u15_u1_n135 ) );
  AOI21_X1 u1_u15_u1_U96 (.ZN( u1_u15_u1_n110 ) , .A( u1_u15_u1_n116 ) , .B1( u1_u15_u1_n152 ) , .B2( u1_u15_u1_n160 ) );
  NAND3_X1 u1_u15_u1_U97 (.A3( u1_u15_u1_n149 ) , .A2( u1_u15_u1_n150 ) , .A1( u1_u15_u1_n151 ) , .ZN( u1_u15_u1_n164 ) );
  NAND3_X1 u1_u15_u1_U98 (.A3( u1_u15_u1_n134 ) , .A2( u1_u15_u1_n135 ) , .ZN( u1_u15_u1_n136 ) , .A1( u1_u15_u1_n151 ) );
  NAND3_X1 u1_u15_u1_U99 (.A1( u1_u15_u1_n133 ) , .ZN( u1_u15_u1_n137 ) , .A2( u1_u15_u1_n154 ) , .A3( u1_u15_u1_n181 ) );
  XOR2_X1 u1_u1_U22 (.B( u1_K2_34 ) , .A( u1_R0_23 ) , .Z( u1_u1_X_34 ) );
  XOR2_X1 u1_u1_U23 (.B( u1_K2_33 ) , .A( u1_R0_22 ) , .Z( u1_u1_X_33 ) );
  INV_X1 u1_u1_u5_U10 (.A( u1_u1_u5_n121 ) , .ZN( u1_u1_u5_n177 ) );
  NOR3_X1 u1_u1_u5_U100 (.A3( u1_u1_u5_n141 ) , .A1( u1_u1_u5_n142 ) , .ZN( u1_u1_u5_n143 ) , .A2( u1_u1_u5_n191 ) );
  NAND4_X1 u1_u1_u5_U101 (.ZN( u1_out1_4 ) , .A4( u1_u1_u5_n112 ) , .A2( u1_u1_u5_n113 ) , .A1( u1_u1_u5_n114 ) , .A3( u1_u1_u5_n195 ) );
  AOI211_X1 u1_u1_u5_U102 (.A( u1_u1_u5_n110 ) , .C1( u1_u1_u5_n111 ) , .ZN( u1_u1_u5_n112 ) , .B( u1_u1_u5_n118 ) , .C2( u1_u1_u5_n177 ) );
  AOI222_X1 u1_u1_u5_U103 (.ZN( u1_u1_u5_n113 ) , .A1( u1_u1_u5_n131 ) , .C1( u1_u1_u5_n148 ) , .B2( u1_u1_u5_n174 ) , .C2( u1_u1_u5_n178 ) , .A2( u1_u1_u5_n179 ) , .B1( u1_u1_u5_n99 ) );
  NAND3_X1 u1_u1_u5_U104 (.A2( u1_u1_u5_n154 ) , .A3( u1_u1_u5_n158 ) , .A1( u1_u1_u5_n161 ) , .ZN( u1_u1_u5_n99 ) );
  NOR2_X1 u1_u1_u5_U11 (.ZN( u1_u1_u5_n160 ) , .A2( u1_u1_u5_n173 ) , .A1( u1_u1_u5_n177 ) );
  INV_X1 u1_u1_u5_U12 (.A( u1_u1_u5_n150 ) , .ZN( u1_u1_u5_n174 ) );
  AOI21_X1 u1_u1_u5_U13 (.A( u1_u1_u5_n160 ) , .B2( u1_u1_u5_n161 ) , .ZN( u1_u1_u5_n162 ) , .B1( u1_u1_u5_n192 ) );
  INV_X1 u1_u1_u5_U14 (.A( u1_u1_u5_n159 ) , .ZN( u1_u1_u5_n192 ) );
  AOI21_X1 u1_u1_u5_U15 (.A( u1_u1_u5_n156 ) , .B2( u1_u1_u5_n157 ) , .B1( u1_u1_u5_n158 ) , .ZN( u1_u1_u5_n163 ) );
  AOI21_X1 u1_u1_u5_U16 (.B2( u1_u1_u5_n139 ) , .B1( u1_u1_u5_n140 ) , .ZN( u1_u1_u5_n141 ) , .A( u1_u1_u5_n150 ) );
  OAI21_X1 u1_u1_u5_U17 (.A( u1_u1_u5_n133 ) , .B2( u1_u1_u5_n134 ) , .B1( u1_u1_u5_n135 ) , .ZN( u1_u1_u5_n142 ) );
  OAI21_X1 u1_u1_u5_U18 (.ZN( u1_u1_u5_n133 ) , .B2( u1_u1_u5_n147 ) , .A( u1_u1_u5_n173 ) , .B1( u1_u1_u5_n188 ) );
  NAND2_X1 u1_u1_u5_U19 (.A2( u1_u1_u5_n119 ) , .A1( u1_u1_u5_n123 ) , .ZN( u1_u1_u5_n137 ) );
  INV_X1 u1_u1_u5_U20 (.A( u1_u1_u5_n155 ) , .ZN( u1_u1_u5_n194 ) );
  NAND2_X1 u1_u1_u5_U21 (.A1( u1_u1_u5_n121 ) , .ZN( u1_u1_u5_n132 ) , .A2( u1_u1_u5_n172 ) );
  NAND2_X1 u1_u1_u5_U22 (.A2( u1_u1_u5_n122 ) , .ZN( u1_u1_u5_n136 ) , .A1( u1_u1_u5_n154 ) );
  NAND2_X1 u1_u1_u5_U23 (.A2( u1_u1_u5_n119 ) , .A1( u1_u1_u5_n120 ) , .ZN( u1_u1_u5_n159 ) );
  INV_X1 u1_u1_u5_U24 (.A( u1_u1_u5_n156 ) , .ZN( u1_u1_u5_n175 ) );
  INV_X1 u1_u1_u5_U25 (.A( u1_u1_u5_n158 ) , .ZN( u1_u1_u5_n188 ) );
  INV_X1 u1_u1_u5_U26 (.A( u1_u1_u5_n152 ) , .ZN( u1_u1_u5_n179 ) );
  INV_X1 u1_u1_u5_U27 (.A( u1_u1_u5_n140 ) , .ZN( u1_u1_u5_n182 ) );
  INV_X1 u1_u1_u5_U28 (.A( u1_u1_u5_n151 ) , .ZN( u1_u1_u5_n183 ) );
  INV_X1 u1_u1_u5_U29 (.A( u1_u1_u5_n123 ) , .ZN( u1_u1_u5_n185 ) );
  NOR2_X1 u1_u1_u5_U3 (.ZN( u1_u1_u5_n134 ) , .A1( u1_u1_u5_n183 ) , .A2( u1_u1_u5_n190 ) );
  INV_X1 u1_u1_u5_U30 (.A( u1_u1_u5_n161 ) , .ZN( u1_u1_u5_n184 ) );
  INV_X1 u1_u1_u5_U31 (.A( u1_u1_u5_n139 ) , .ZN( u1_u1_u5_n189 ) );
  INV_X1 u1_u1_u5_U32 (.A( u1_u1_u5_n157 ) , .ZN( u1_u1_u5_n190 ) );
  INV_X1 u1_u1_u5_U33 (.A( u1_u1_u5_n120 ) , .ZN( u1_u1_u5_n193 ) );
  NAND2_X1 u1_u1_u5_U34 (.ZN( u1_u1_u5_n111 ) , .A1( u1_u1_u5_n140 ) , .A2( u1_u1_u5_n155 ) );
  INV_X1 u1_u1_u5_U35 (.A( u1_u1_u5_n117 ) , .ZN( u1_u1_u5_n196 ) );
  OAI221_X1 u1_u1_u5_U36 (.A( u1_u1_u5_n116 ) , .ZN( u1_u1_u5_n117 ) , .B2( u1_u1_u5_n119 ) , .C1( u1_u1_u5_n153 ) , .C2( u1_u1_u5_n158 ) , .B1( u1_u1_u5_n172 ) );
  AOI222_X1 u1_u1_u5_U37 (.ZN( u1_u1_u5_n116 ) , .B2( u1_u1_u5_n145 ) , .C1( u1_u1_u5_n148 ) , .A2( u1_u1_u5_n174 ) , .C2( u1_u1_u5_n177 ) , .B1( u1_u1_u5_n187 ) , .A1( u1_u1_u5_n193 ) );
  INV_X1 u1_u1_u5_U38 (.A( u1_u1_u5_n115 ) , .ZN( u1_u1_u5_n187 ) );
  NOR2_X1 u1_u1_u5_U39 (.ZN( u1_u1_u5_n100 ) , .A1( u1_u1_u5_n170 ) , .A2( u1_u1_u5_n180 ) );
  INV_X1 u1_u1_u5_U4 (.A( u1_u1_u5_n138 ) , .ZN( u1_u1_u5_n191 ) );
  AOI22_X1 u1_u1_u5_U40 (.B2( u1_u1_u5_n131 ) , .A2( u1_u1_u5_n146 ) , .ZN( u1_u1_u5_n169 ) , .B1( u1_u1_u5_n174 ) , .A1( u1_u1_u5_n185 ) );
  NOR2_X1 u1_u1_u5_U41 (.A1( u1_u1_u5_n146 ) , .ZN( u1_u1_u5_n150 ) , .A2( u1_u1_u5_n173 ) );
  AOI21_X1 u1_u1_u5_U42 (.A( u1_u1_u5_n118 ) , .B2( u1_u1_u5_n145 ) , .ZN( u1_u1_u5_n168 ) , .B1( u1_u1_u5_n186 ) );
  INV_X1 u1_u1_u5_U43 (.A( u1_u1_u5_n122 ) , .ZN( u1_u1_u5_n186 ) );
  NOR2_X1 u1_u1_u5_U44 (.A1( u1_u1_u5_n146 ) , .ZN( u1_u1_u5_n152 ) , .A2( u1_u1_u5_n176 ) );
  NOR2_X1 u1_u1_u5_U45 (.A1( u1_u1_u5_n115 ) , .ZN( u1_u1_u5_n118 ) , .A2( u1_u1_u5_n153 ) );
  NOR2_X1 u1_u1_u5_U46 (.A2( u1_u1_u5_n145 ) , .ZN( u1_u1_u5_n156 ) , .A1( u1_u1_u5_n174 ) );
  NOR2_X1 u1_u1_u5_U47 (.ZN( u1_u1_u5_n121 ) , .A2( u1_u1_u5_n145 ) , .A1( u1_u1_u5_n176 ) );
  AOI22_X1 u1_u1_u5_U48 (.ZN( u1_u1_u5_n114 ) , .A2( u1_u1_u5_n137 ) , .A1( u1_u1_u5_n145 ) , .B2( u1_u1_u5_n175 ) , .B1( u1_u1_u5_n193 ) );
  OAI211_X1 u1_u1_u5_U49 (.B( u1_u1_u5_n124 ) , .A( u1_u1_u5_n125 ) , .C2( u1_u1_u5_n126 ) , .C1( u1_u1_u5_n127 ) , .ZN( u1_u1_u5_n128 ) );
  OAI21_X1 u1_u1_u5_U5 (.B2( u1_u1_u5_n136 ) , .B1( u1_u1_u5_n137 ) , .ZN( u1_u1_u5_n138 ) , .A( u1_u1_u5_n177 ) );
  OAI21_X1 u1_u1_u5_U50 (.ZN( u1_u1_u5_n124 ) , .A( u1_u1_u5_n177 ) , .B2( u1_u1_u5_n183 ) , .B1( u1_u1_u5_n189 ) );
  NOR3_X1 u1_u1_u5_U51 (.ZN( u1_u1_u5_n127 ) , .A1( u1_u1_u5_n136 ) , .A3( u1_u1_u5_n148 ) , .A2( u1_u1_u5_n182 ) );
  OAI21_X1 u1_u1_u5_U52 (.ZN( u1_u1_u5_n125 ) , .A( u1_u1_u5_n174 ) , .B2( u1_u1_u5_n185 ) , .B1( u1_u1_u5_n190 ) );
  AOI21_X1 u1_u1_u5_U53 (.A( u1_u1_u5_n153 ) , .B2( u1_u1_u5_n154 ) , .B1( u1_u1_u5_n155 ) , .ZN( u1_u1_u5_n164 ) );
  AOI21_X1 u1_u1_u5_U54 (.ZN( u1_u1_u5_n110 ) , .B1( u1_u1_u5_n122 ) , .B2( u1_u1_u5_n139 ) , .A( u1_u1_u5_n153 ) );
  INV_X1 u1_u1_u5_U55 (.A( u1_u1_u5_n153 ) , .ZN( u1_u1_u5_n176 ) );
  INV_X1 u1_u1_u5_U56 (.A( u1_u1_u5_n126 ) , .ZN( u1_u1_u5_n173 ) );
  AND2_X1 u1_u1_u5_U57 (.A2( u1_u1_u5_n104 ) , .A1( u1_u1_u5_n107 ) , .ZN( u1_u1_u5_n147 ) );
  AND2_X1 u1_u1_u5_U58 (.A2( u1_u1_u5_n104 ) , .A1( u1_u1_u5_n108 ) , .ZN( u1_u1_u5_n148 ) );
  NAND2_X1 u1_u1_u5_U59 (.A1( u1_u1_u5_n105 ) , .A2( u1_u1_u5_n106 ) , .ZN( u1_u1_u5_n158 ) );
  INV_X1 u1_u1_u5_U6 (.A( u1_u1_u5_n135 ) , .ZN( u1_u1_u5_n178 ) );
  NAND2_X1 u1_u1_u5_U60 (.A2( u1_u1_u5_n108 ) , .A1( u1_u1_u5_n109 ) , .ZN( u1_u1_u5_n139 ) );
  NAND2_X1 u1_u1_u5_U61 (.A1( u1_u1_u5_n106 ) , .A2( u1_u1_u5_n108 ) , .ZN( u1_u1_u5_n119 ) );
  NAND2_X1 u1_u1_u5_U62 (.A2( u1_u1_u5_n103 ) , .A1( u1_u1_u5_n105 ) , .ZN( u1_u1_u5_n140 ) );
  NAND2_X1 u1_u1_u5_U63 (.A2( u1_u1_u5_n104 ) , .A1( u1_u1_u5_n105 ) , .ZN( u1_u1_u5_n155 ) );
  NAND2_X1 u1_u1_u5_U64 (.A2( u1_u1_u5_n106 ) , .A1( u1_u1_u5_n107 ) , .ZN( u1_u1_u5_n122 ) );
  NAND2_X1 u1_u1_u5_U65 (.A2( u1_u1_u5_n100 ) , .A1( u1_u1_u5_n106 ) , .ZN( u1_u1_u5_n115 ) );
  NAND2_X1 u1_u1_u5_U66 (.A2( u1_u1_u5_n100 ) , .A1( u1_u1_u5_n103 ) , .ZN( u1_u1_u5_n161 ) );
  NAND2_X1 u1_u1_u5_U67 (.A1( u1_u1_u5_n105 ) , .A2( u1_u1_u5_n109 ) , .ZN( u1_u1_u5_n154 ) );
  INV_X1 u1_u1_u5_U68 (.A( u1_u1_u5_n146 ) , .ZN( u1_u1_u5_n172 ) );
  NAND2_X1 u1_u1_u5_U69 (.A1( u1_u1_u5_n103 ) , .A2( u1_u1_u5_n108 ) , .ZN( u1_u1_u5_n123 ) );
  OAI22_X1 u1_u1_u5_U7 (.B2( u1_u1_u5_n149 ) , .B1( u1_u1_u5_n150 ) , .A2( u1_u1_u5_n151 ) , .A1( u1_u1_u5_n152 ) , .ZN( u1_u1_u5_n165 ) );
  NAND2_X1 u1_u1_u5_U70 (.A2( u1_u1_u5_n103 ) , .A1( u1_u1_u5_n107 ) , .ZN( u1_u1_u5_n151 ) );
  NAND2_X1 u1_u1_u5_U71 (.A2( u1_u1_u5_n107 ) , .A1( u1_u1_u5_n109 ) , .ZN( u1_u1_u5_n120 ) );
  NAND2_X1 u1_u1_u5_U72 (.A2( u1_u1_u5_n100 ) , .A1( u1_u1_u5_n109 ) , .ZN( u1_u1_u5_n157 ) );
  AND2_X1 u1_u1_u5_U73 (.A2( u1_u1_u5_n100 ) , .A1( u1_u1_u5_n104 ) , .ZN( u1_u1_u5_n131 ) );
  INV_X1 u1_u1_u5_U74 (.A( u1_u1_u5_n102 ) , .ZN( u1_u1_u5_n195 ) );
  OAI221_X1 u1_u1_u5_U75 (.A( u1_u1_u5_n101 ) , .ZN( u1_u1_u5_n102 ) , .C2( u1_u1_u5_n115 ) , .C1( u1_u1_u5_n126 ) , .B1( u1_u1_u5_n134 ) , .B2( u1_u1_u5_n160 ) );
  OAI21_X1 u1_u1_u5_U76 (.ZN( u1_u1_u5_n101 ) , .B1( u1_u1_u5_n137 ) , .A( u1_u1_u5_n146 ) , .B2( u1_u1_u5_n147 ) );
  NOR2_X1 u1_u1_u5_U77 (.A2( u1_u1_X_34 ) , .A1( u1_u1_X_35 ) , .ZN( u1_u1_u5_n145 ) );
  NOR2_X1 u1_u1_u5_U78 (.A2( u1_u1_X_34 ) , .ZN( u1_u1_u5_n146 ) , .A1( u1_u1_u5_n171 ) );
  NOR2_X1 u1_u1_u5_U79 (.A2( u1_u1_X_31 ) , .A1( u1_u1_X_32 ) , .ZN( u1_u1_u5_n103 ) );
  NOR3_X1 u1_u1_u5_U8 (.A2( u1_u1_u5_n147 ) , .A1( u1_u1_u5_n148 ) , .ZN( u1_u1_u5_n149 ) , .A3( u1_u1_u5_n194 ) );
  NOR2_X1 u1_u1_u5_U80 (.A2( u1_u1_X_36 ) , .ZN( u1_u1_u5_n105 ) , .A1( u1_u1_u5_n180 ) );
  NOR2_X1 u1_u1_u5_U81 (.A2( u1_u1_X_33 ) , .ZN( u1_u1_u5_n108 ) , .A1( u1_u1_u5_n170 ) );
  NOR2_X1 u1_u1_u5_U82 (.A2( u1_u1_X_33 ) , .A1( u1_u1_X_36 ) , .ZN( u1_u1_u5_n107 ) );
  NOR2_X1 u1_u1_u5_U83 (.A2( u1_u1_X_31 ) , .ZN( u1_u1_u5_n104 ) , .A1( u1_u1_u5_n181 ) );
  NAND2_X1 u1_u1_u5_U84 (.A2( u1_u1_X_34 ) , .A1( u1_u1_X_35 ) , .ZN( u1_u1_u5_n153 ) );
  NAND2_X1 u1_u1_u5_U85 (.A1( u1_u1_X_34 ) , .ZN( u1_u1_u5_n126 ) , .A2( u1_u1_u5_n171 ) );
  AND2_X1 u1_u1_u5_U86 (.A1( u1_u1_X_31 ) , .A2( u1_u1_X_32 ) , .ZN( u1_u1_u5_n106 ) );
  AND2_X1 u1_u1_u5_U87 (.A1( u1_u1_X_31 ) , .ZN( u1_u1_u5_n109 ) , .A2( u1_u1_u5_n181 ) );
  INV_X1 u1_u1_u5_U88 (.A( u1_u1_X_33 ) , .ZN( u1_u1_u5_n180 ) );
  INV_X1 u1_u1_u5_U89 (.A( u1_u1_X_35 ) , .ZN( u1_u1_u5_n171 ) );
  NOR2_X1 u1_u1_u5_U9 (.ZN( u1_u1_u5_n135 ) , .A1( u1_u1_u5_n173 ) , .A2( u1_u1_u5_n176 ) );
  INV_X1 u1_u1_u5_U90 (.A( u1_u1_X_36 ) , .ZN( u1_u1_u5_n170 ) );
  INV_X1 u1_u1_u5_U91 (.A( u1_u1_X_32 ) , .ZN( u1_u1_u5_n181 ) );
  NAND4_X1 u1_u1_u5_U92 (.ZN( u1_out1_29 ) , .A4( u1_u1_u5_n129 ) , .A3( u1_u1_u5_n130 ) , .A2( u1_u1_u5_n168 ) , .A1( u1_u1_u5_n196 ) );
  AOI221_X1 u1_u1_u5_U93 (.A( u1_u1_u5_n128 ) , .ZN( u1_u1_u5_n129 ) , .C2( u1_u1_u5_n132 ) , .B2( u1_u1_u5_n159 ) , .B1( u1_u1_u5_n176 ) , .C1( u1_u1_u5_n184 ) );
  AOI222_X1 u1_u1_u5_U94 (.ZN( u1_u1_u5_n130 ) , .A2( u1_u1_u5_n146 ) , .B1( u1_u1_u5_n147 ) , .C2( u1_u1_u5_n175 ) , .B2( u1_u1_u5_n179 ) , .A1( u1_u1_u5_n188 ) , .C1( u1_u1_u5_n194 ) );
  NAND4_X1 u1_u1_u5_U95 (.ZN( u1_out1_19 ) , .A4( u1_u1_u5_n166 ) , .A3( u1_u1_u5_n167 ) , .A2( u1_u1_u5_n168 ) , .A1( u1_u1_u5_n169 ) );
  AOI22_X1 u1_u1_u5_U96 (.B2( u1_u1_u5_n145 ) , .A2( u1_u1_u5_n146 ) , .ZN( u1_u1_u5_n167 ) , .B1( u1_u1_u5_n182 ) , .A1( u1_u1_u5_n189 ) );
  NOR4_X1 u1_u1_u5_U97 (.A4( u1_u1_u5_n162 ) , .A3( u1_u1_u5_n163 ) , .A2( u1_u1_u5_n164 ) , .A1( u1_u1_u5_n165 ) , .ZN( u1_u1_u5_n166 ) );
  NAND4_X1 u1_u1_u5_U98 (.ZN( u1_out1_11 ) , .A4( u1_u1_u5_n143 ) , .A3( u1_u1_u5_n144 ) , .A2( u1_u1_u5_n169 ) , .A1( u1_u1_u5_n196 ) );
  AOI22_X1 u1_u1_u5_U99 (.A2( u1_u1_u5_n132 ) , .ZN( u1_u1_u5_n144 ) , .B2( u1_u1_u5_n145 ) , .B1( u1_u1_u5_n184 ) , .A1( u1_u1_u5_n194 ) );
  XOR2_X1 u1_u2_U1 (.B( u1_K3_9 ) , .A( u1_R1_6 ) , .Z( u1_u2_X_9 ) );
  XOR2_X1 u1_u2_U16 (.B( u1_K3_3 ) , .A( u1_R1_2 ) , .Z( u1_u2_X_3 ) );
  XOR2_X1 u1_u2_U3 (.B( u1_K3_7 ) , .A( u1_R1_4 ) , .Z( u1_u2_X_7 ) );
  XOR2_X1 u1_u2_U48 (.B( u1_K3_10 ) , .A( u1_R1_7 ) , .Z( u1_u2_X_10 ) );
  XOR2_X1 u1_u2_U5 (.B( u1_K3_5 ) , .A( u1_R1_4 ) , .Z( u1_u2_X_5 ) );
  XOR2_X1 u1_u2_U6 (.B( u1_K3_4 ) , .A( u1_R1_3 ) , .Z( u1_u2_X_4 ) );
  AND3_X1 u1_u2_u0_U10 (.A2( u1_u2_u0_n112 ) , .ZN( u1_u2_u0_n127 ) , .A3( u1_u2_u0_n130 ) , .A1( u1_u2_u0_n148 ) );
  NAND2_X1 u1_u2_u0_U11 (.ZN( u1_u2_u0_n113 ) , .A1( u1_u2_u0_n139 ) , .A2( u1_u2_u0_n149 ) );
  AND2_X1 u1_u2_u0_U12 (.ZN( u1_u2_u0_n107 ) , .A1( u1_u2_u0_n130 ) , .A2( u1_u2_u0_n140 ) );
  AND2_X1 u1_u2_u0_U13 (.A2( u1_u2_u0_n129 ) , .A1( u1_u2_u0_n130 ) , .ZN( u1_u2_u0_n151 ) );
  AND2_X1 u1_u2_u0_U14 (.A1( u1_u2_u0_n108 ) , .A2( u1_u2_u0_n125 ) , .ZN( u1_u2_u0_n145 ) );
  INV_X1 u1_u2_u0_U15 (.A( u1_u2_u0_n143 ) , .ZN( u1_u2_u0_n173 ) );
  NOR2_X1 u1_u2_u0_U16 (.A2( u1_u2_u0_n136 ) , .ZN( u1_u2_u0_n147 ) , .A1( u1_u2_u0_n160 ) );
  INV_X1 u1_u2_u0_U17 (.ZN( u1_u2_u0_n172 ) , .A( u1_u2_u0_n88 ) );
  OAI222_X1 u1_u2_u0_U18 (.C1( u1_u2_u0_n108 ) , .A1( u1_u2_u0_n125 ) , .B2( u1_u2_u0_n128 ) , .B1( u1_u2_u0_n144 ) , .A2( u1_u2_u0_n158 ) , .C2( u1_u2_u0_n161 ) , .ZN( u1_u2_u0_n88 ) );
  NOR2_X1 u1_u2_u0_U19 (.A1( u1_u2_u0_n163 ) , .A2( u1_u2_u0_n164 ) , .ZN( u1_u2_u0_n95 ) );
  AOI21_X1 u1_u2_u0_U20 (.B1( u1_u2_u0_n103 ) , .ZN( u1_u2_u0_n132 ) , .A( u1_u2_u0_n165 ) , .B2( u1_u2_u0_n93 ) );
  INV_X1 u1_u2_u0_U21 (.A( u1_u2_u0_n142 ) , .ZN( u1_u2_u0_n165 ) );
  OAI221_X1 u1_u2_u0_U22 (.C1( u1_u2_u0_n121 ) , .ZN( u1_u2_u0_n122 ) , .B2( u1_u2_u0_n127 ) , .A( u1_u2_u0_n143 ) , .B1( u1_u2_u0_n144 ) , .C2( u1_u2_u0_n147 ) );
  OAI22_X1 u1_u2_u0_U23 (.B1( u1_u2_u0_n125 ) , .ZN( u1_u2_u0_n126 ) , .A1( u1_u2_u0_n138 ) , .A2( u1_u2_u0_n146 ) , .B2( u1_u2_u0_n147 ) );
  OAI22_X1 u1_u2_u0_U24 (.B1( u1_u2_u0_n131 ) , .A1( u1_u2_u0_n144 ) , .B2( u1_u2_u0_n147 ) , .A2( u1_u2_u0_n90 ) , .ZN( u1_u2_u0_n91 ) );
  AND3_X1 u1_u2_u0_U25 (.A3( u1_u2_u0_n121 ) , .A2( u1_u2_u0_n125 ) , .A1( u1_u2_u0_n148 ) , .ZN( u1_u2_u0_n90 ) );
  INV_X1 u1_u2_u0_U26 (.A( u1_u2_u0_n136 ) , .ZN( u1_u2_u0_n161 ) );
  NOR2_X1 u1_u2_u0_U27 (.A1( u1_u2_u0_n120 ) , .ZN( u1_u2_u0_n143 ) , .A2( u1_u2_u0_n167 ) );
  OAI221_X1 u1_u2_u0_U28 (.C1( u1_u2_u0_n112 ) , .ZN( u1_u2_u0_n120 ) , .B1( u1_u2_u0_n138 ) , .B2( u1_u2_u0_n141 ) , .C2( u1_u2_u0_n147 ) , .A( u1_u2_u0_n172 ) );
  AOI211_X1 u1_u2_u0_U29 (.B( u1_u2_u0_n115 ) , .A( u1_u2_u0_n116 ) , .C2( u1_u2_u0_n117 ) , .C1( u1_u2_u0_n118 ) , .ZN( u1_u2_u0_n119 ) );
  INV_X1 u1_u2_u0_U3 (.A( u1_u2_u0_n113 ) , .ZN( u1_u2_u0_n166 ) );
  AOI22_X1 u1_u2_u0_U30 (.B2( u1_u2_u0_n109 ) , .A2( u1_u2_u0_n110 ) , .ZN( u1_u2_u0_n111 ) , .B1( u1_u2_u0_n118 ) , .A1( u1_u2_u0_n160 ) );
  INV_X1 u1_u2_u0_U31 (.A( u1_u2_u0_n118 ) , .ZN( u1_u2_u0_n158 ) );
  AOI21_X1 u1_u2_u0_U32 (.ZN( u1_u2_u0_n104 ) , .B1( u1_u2_u0_n107 ) , .B2( u1_u2_u0_n141 ) , .A( u1_u2_u0_n144 ) );
  AOI21_X1 u1_u2_u0_U33 (.B1( u1_u2_u0_n127 ) , .B2( u1_u2_u0_n129 ) , .A( u1_u2_u0_n138 ) , .ZN( u1_u2_u0_n96 ) );
  AOI21_X1 u1_u2_u0_U34 (.ZN( u1_u2_u0_n116 ) , .B2( u1_u2_u0_n142 ) , .A( u1_u2_u0_n144 ) , .B1( u1_u2_u0_n166 ) );
  NAND2_X1 u1_u2_u0_U35 (.A1( u1_u2_u0_n100 ) , .A2( u1_u2_u0_n103 ) , .ZN( u1_u2_u0_n125 ) );
  NAND2_X1 u1_u2_u0_U36 (.A1( u1_u2_u0_n101 ) , .A2( u1_u2_u0_n102 ) , .ZN( u1_u2_u0_n150 ) );
  INV_X1 u1_u2_u0_U37 (.A( u1_u2_u0_n138 ) , .ZN( u1_u2_u0_n160 ) );
  NAND2_X1 u1_u2_u0_U38 (.A1( u1_u2_u0_n102 ) , .ZN( u1_u2_u0_n128 ) , .A2( u1_u2_u0_n95 ) );
  NAND2_X1 u1_u2_u0_U39 (.A1( u1_u2_u0_n100 ) , .ZN( u1_u2_u0_n129 ) , .A2( u1_u2_u0_n95 ) );
  AOI21_X1 u1_u2_u0_U4 (.B1( u1_u2_u0_n114 ) , .ZN( u1_u2_u0_n115 ) , .B2( u1_u2_u0_n129 ) , .A( u1_u2_u0_n161 ) );
  NAND2_X1 u1_u2_u0_U40 (.A2( u1_u2_u0_n100 ) , .ZN( u1_u2_u0_n131 ) , .A1( u1_u2_u0_n92 ) );
  NAND2_X1 u1_u2_u0_U41 (.A2( u1_u2_u0_n100 ) , .A1( u1_u2_u0_n101 ) , .ZN( u1_u2_u0_n139 ) );
  NAND2_X1 u1_u2_u0_U42 (.ZN( u1_u2_u0_n148 ) , .A1( u1_u2_u0_n93 ) , .A2( u1_u2_u0_n95 ) );
  NAND2_X1 u1_u2_u0_U43 (.A2( u1_u2_u0_n102 ) , .A1( u1_u2_u0_n103 ) , .ZN( u1_u2_u0_n149 ) );
  NAND2_X1 u1_u2_u0_U44 (.A2( u1_u2_u0_n102 ) , .ZN( u1_u2_u0_n114 ) , .A1( u1_u2_u0_n92 ) );
  NAND2_X1 u1_u2_u0_U45 (.A2( u1_u2_u0_n101 ) , .ZN( u1_u2_u0_n121 ) , .A1( u1_u2_u0_n93 ) );
  NAND2_X1 u1_u2_u0_U46 (.ZN( u1_u2_u0_n112 ) , .A2( u1_u2_u0_n92 ) , .A1( u1_u2_u0_n93 ) );
  OR3_X1 u1_u2_u0_U47 (.A3( u1_u2_u0_n152 ) , .A2( u1_u2_u0_n153 ) , .A1( u1_u2_u0_n154 ) , .ZN( u1_u2_u0_n155 ) );
  AOI21_X1 u1_u2_u0_U48 (.B2( u1_u2_u0_n150 ) , .B1( u1_u2_u0_n151 ) , .ZN( u1_u2_u0_n152 ) , .A( u1_u2_u0_n158 ) );
  AOI21_X1 u1_u2_u0_U49 (.A( u1_u2_u0_n144 ) , .B2( u1_u2_u0_n145 ) , .B1( u1_u2_u0_n146 ) , .ZN( u1_u2_u0_n154 ) );
  AOI21_X1 u1_u2_u0_U5 (.B2( u1_u2_u0_n131 ) , .ZN( u1_u2_u0_n134 ) , .B1( u1_u2_u0_n151 ) , .A( u1_u2_u0_n158 ) );
  AOI21_X1 u1_u2_u0_U50 (.A( u1_u2_u0_n147 ) , .B2( u1_u2_u0_n148 ) , .B1( u1_u2_u0_n149 ) , .ZN( u1_u2_u0_n153 ) );
  INV_X1 u1_u2_u0_U51 (.ZN( u1_u2_u0_n171 ) , .A( u1_u2_u0_n99 ) );
  OAI211_X1 u1_u2_u0_U52 (.C2( u1_u2_u0_n140 ) , .C1( u1_u2_u0_n161 ) , .A( u1_u2_u0_n169 ) , .B( u1_u2_u0_n98 ) , .ZN( u1_u2_u0_n99 ) );
  AOI211_X1 u1_u2_u0_U53 (.C1( u1_u2_u0_n118 ) , .A( u1_u2_u0_n123 ) , .B( u1_u2_u0_n96 ) , .C2( u1_u2_u0_n97 ) , .ZN( u1_u2_u0_n98 ) );
  INV_X1 u1_u2_u0_U54 (.ZN( u1_u2_u0_n169 ) , .A( u1_u2_u0_n91 ) );
  NOR2_X1 u1_u2_u0_U55 (.A2( u1_u2_X_6 ) , .ZN( u1_u2_u0_n100 ) , .A1( u1_u2_u0_n162 ) );
  NOR2_X1 u1_u2_u0_U56 (.A2( u1_u2_X_4 ) , .A1( u1_u2_X_5 ) , .ZN( u1_u2_u0_n118 ) );
  NOR2_X1 u1_u2_u0_U57 (.A2( u1_u2_X_2 ) , .ZN( u1_u2_u0_n103 ) , .A1( u1_u2_u0_n164 ) );
  NOR2_X1 u1_u2_u0_U58 (.A2( u1_u2_X_1 ) , .A1( u1_u2_X_2 ) , .ZN( u1_u2_u0_n92 ) );
  NOR2_X1 u1_u2_u0_U59 (.A2( u1_u2_X_1 ) , .ZN( u1_u2_u0_n101 ) , .A1( u1_u2_u0_n163 ) );
  NOR2_X1 u1_u2_u0_U6 (.A1( u1_u2_u0_n108 ) , .ZN( u1_u2_u0_n123 ) , .A2( u1_u2_u0_n158 ) );
  NAND2_X1 u1_u2_u0_U60 (.A2( u1_u2_X_4 ) , .A1( u1_u2_X_5 ) , .ZN( u1_u2_u0_n144 ) );
  NOR2_X1 u1_u2_u0_U61 (.A2( u1_u2_X_5 ) , .ZN( u1_u2_u0_n136 ) , .A1( u1_u2_u0_n159 ) );
  NAND2_X1 u1_u2_u0_U62 (.A1( u1_u2_X_5 ) , .ZN( u1_u2_u0_n138 ) , .A2( u1_u2_u0_n159 ) );
  AND2_X1 u1_u2_u0_U63 (.A2( u1_u2_X_3 ) , .A1( u1_u2_X_6 ) , .ZN( u1_u2_u0_n102 ) );
  AND2_X1 u1_u2_u0_U64 (.A1( u1_u2_X_6 ) , .A2( u1_u2_u0_n162 ) , .ZN( u1_u2_u0_n93 ) );
  INV_X1 u1_u2_u0_U65 (.A( u1_u2_X_4 ) , .ZN( u1_u2_u0_n159 ) );
  INV_X1 u1_u2_u0_U66 (.A( u1_u2_X_1 ) , .ZN( u1_u2_u0_n164 ) );
  INV_X1 u1_u2_u0_U67 (.A( u1_u2_X_2 ) , .ZN( u1_u2_u0_n163 ) );
  INV_X1 u1_u2_u0_U68 (.ZN( u1_u2_u0_n174 ) , .A( u1_u2_u0_n89 ) );
  AOI211_X1 u1_u2_u0_U69 (.B( u1_u2_u0_n104 ) , .A( u1_u2_u0_n105 ) , .ZN( u1_u2_u0_n106 ) , .C2( u1_u2_u0_n113 ) , .C1( u1_u2_u0_n160 ) );
  OAI21_X1 u1_u2_u0_U7 (.B1( u1_u2_u0_n150 ) , .B2( u1_u2_u0_n158 ) , .A( u1_u2_u0_n172 ) , .ZN( u1_u2_u0_n89 ) );
  OR4_X1 u1_u2_u0_U70 (.ZN( u1_out2_17 ) , .A4( u1_u2_u0_n122 ) , .A2( u1_u2_u0_n123 ) , .A1( u1_u2_u0_n124 ) , .A3( u1_u2_u0_n170 ) );
  AOI21_X1 u1_u2_u0_U71 (.B2( u1_u2_u0_n107 ) , .ZN( u1_u2_u0_n124 ) , .B1( u1_u2_u0_n128 ) , .A( u1_u2_u0_n161 ) );
  INV_X1 u1_u2_u0_U72 (.A( u1_u2_u0_n111 ) , .ZN( u1_u2_u0_n170 ) );
  OR4_X1 u1_u2_u0_U73 (.ZN( u1_out2_31 ) , .A4( u1_u2_u0_n155 ) , .A2( u1_u2_u0_n156 ) , .A1( u1_u2_u0_n157 ) , .A3( u1_u2_u0_n173 ) );
  AOI21_X1 u1_u2_u0_U74 (.A( u1_u2_u0_n138 ) , .B2( u1_u2_u0_n139 ) , .B1( u1_u2_u0_n140 ) , .ZN( u1_u2_u0_n157 ) );
  AOI21_X1 u1_u2_u0_U75 (.B2( u1_u2_u0_n141 ) , .B1( u1_u2_u0_n142 ) , .ZN( u1_u2_u0_n156 ) , .A( u1_u2_u0_n161 ) );
  INV_X1 u1_u2_u0_U76 (.A( u1_u2_u0_n126 ) , .ZN( u1_u2_u0_n168 ) );
  AOI211_X1 u1_u2_u0_U77 (.B( u1_u2_u0_n133 ) , .A( u1_u2_u0_n134 ) , .C2( u1_u2_u0_n135 ) , .C1( u1_u2_u0_n136 ) , .ZN( u1_u2_u0_n137 ) );
  AOI21_X1 u1_u2_u0_U78 (.B1( u1_u2_u0_n132 ) , .ZN( u1_u2_u0_n133 ) , .A( u1_u2_u0_n144 ) , .B2( u1_u2_u0_n166 ) );
  OAI22_X1 u1_u2_u0_U79 (.ZN( u1_u2_u0_n105 ) , .A2( u1_u2_u0_n132 ) , .B1( u1_u2_u0_n146 ) , .A1( u1_u2_u0_n147 ) , .B2( u1_u2_u0_n161 ) );
  AND2_X1 u1_u2_u0_U8 (.A1( u1_u2_u0_n114 ) , .A2( u1_u2_u0_n121 ) , .ZN( u1_u2_u0_n146 ) );
  NAND2_X1 u1_u2_u0_U80 (.ZN( u1_u2_u0_n110 ) , .A2( u1_u2_u0_n132 ) , .A1( u1_u2_u0_n145 ) );
  INV_X1 u1_u2_u0_U81 (.A( u1_u2_u0_n119 ) , .ZN( u1_u2_u0_n167 ) );
  NAND2_X1 u1_u2_u0_U82 (.A2( u1_u2_u0_n103 ) , .ZN( u1_u2_u0_n140 ) , .A1( u1_u2_u0_n94 ) );
  NAND2_X1 u1_u2_u0_U83 (.A1( u1_u2_u0_n101 ) , .ZN( u1_u2_u0_n130 ) , .A2( u1_u2_u0_n94 ) );
  NAND2_X1 u1_u2_u0_U84 (.ZN( u1_u2_u0_n108 ) , .A1( u1_u2_u0_n92 ) , .A2( u1_u2_u0_n94 ) );
  NAND2_X1 u1_u2_u0_U85 (.ZN( u1_u2_u0_n142 ) , .A1( u1_u2_u0_n94 ) , .A2( u1_u2_u0_n95 ) );
  INV_X1 u1_u2_u0_U86 (.A( u1_u2_X_3 ) , .ZN( u1_u2_u0_n162 ) );
  NOR2_X1 u1_u2_u0_U87 (.A2( u1_u2_X_3 ) , .A1( u1_u2_X_6 ) , .ZN( u1_u2_u0_n94 ) );
  NAND3_X1 u1_u2_u0_U88 (.ZN( u1_out2_23 ) , .A3( u1_u2_u0_n137 ) , .A1( u1_u2_u0_n168 ) , .A2( u1_u2_u0_n171 ) );
  NAND3_X1 u1_u2_u0_U89 (.A3( u1_u2_u0_n127 ) , .A2( u1_u2_u0_n128 ) , .ZN( u1_u2_u0_n135 ) , .A1( u1_u2_u0_n150 ) );
  AND2_X1 u1_u2_u0_U9 (.A1( u1_u2_u0_n131 ) , .ZN( u1_u2_u0_n141 ) , .A2( u1_u2_u0_n150 ) );
  NAND3_X1 u1_u2_u0_U90 (.ZN( u1_u2_u0_n117 ) , .A3( u1_u2_u0_n132 ) , .A2( u1_u2_u0_n139 ) , .A1( u1_u2_u0_n148 ) );
  NAND3_X1 u1_u2_u0_U91 (.ZN( u1_u2_u0_n109 ) , .A2( u1_u2_u0_n114 ) , .A3( u1_u2_u0_n140 ) , .A1( u1_u2_u0_n149 ) );
  NAND3_X1 u1_u2_u0_U92 (.ZN( u1_out2_9 ) , .A3( u1_u2_u0_n106 ) , .A2( u1_u2_u0_n171 ) , .A1( u1_u2_u0_n174 ) );
  NAND3_X1 u1_u2_u0_U93 (.A2( u1_u2_u0_n128 ) , .A1( u1_u2_u0_n132 ) , .A3( u1_u2_u0_n146 ) , .ZN( u1_u2_u0_n97 ) );
  NOR2_X1 u1_u2_u1_U10 (.A1( u1_u2_u1_n112 ) , .A2( u1_u2_u1_n116 ) , .ZN( u1_u2_u1_n118 ) );
  NAND3_X1 u1_u2_u1_U100 (.ZN( u1_u2_u1_n113 ) , .A1( u1_u2_u1_n120 ) , .A3( u1_u2_u1_n133 ) , .A2( u1_u2_u1_n155 ) );
  OAI21_X1 u1_u2_u1_U11 (.ZN( u1_u2_u1_n101 ) , .B1( u1_u2_u1_n141 ) , .A( u1_u2_u1_n146 ) , .B2( u1_u2_u1_n183 ) );
  AOI21_X1 u1_u2_u1_U12 (.B2( u1_u2_u1_n155 ) , .B1( u1_u2_u1_n156 ) , .ZN( u1_u2_u1_n157 ) , .A( u1_u2_u1_n174 ) );
  OR4_X1 u1_u2_u1_U13 (.A4( u1_u2_u1_n106 ) , .A3( u1_u2_u1_n107 ) , .ZN( u1_u2_u1_n108 ) , .A1( u1_u2_u1_n117 ) , .A2( u1_u2_u1_n184 ) );
  AOI21_X1 u1_u2_u1_U14 (.ZN( u1_u2_u1_n106 ) , .A( u1_u2_u1_n112 ) , .B1( u1_u2_u1_n154 ) , .B2( u1_u2_u1_n156 ) );
  INV_X1 u1_u2_u1_U15 (.A( u1_u2_u1_n101 ) , .ZN( u1_u2_u1_n184 ) );
  AOI21_X1 u1_u2_u1_U16 (.ZN( u1_u2_u1_n107 ) , .B1( u1_u2_u1_n134 ) , .B2( u1_u2_u1_n149 ) , .A( u1_u2_u1_n174 ) );
  NAND2_X1 u1_u2_u1_U17 (.ZN( u1_u2_u1_n140 ) , .A2( u1_u2_u1_n150 ) , .A1( u1_u2_u1_n155 ) );
  NAND2_X1 u1_u2_u1_U18 (.A1( u1_u2_u1_n131 ) , .ZN( u1_u2_u1_n147 ) , .A2( u1_u2_u1_n153 ) );
  INV_X1 u1_u2_u1_U19 (.A( u1_u2_u1_n139 ) , .ZN( u1_u2_u1_n174 ) );
  INV_X1 u1_u2_u1_U20 (.A( u1_u2_u1_n112 ) , .ZN( u1_u2_u1_n171 ) );
  NAND2_X1 u1_u2_u1_U21 (.ZN( u1_u2_u1_n141 ) , .A1( u1_u2_u1_n153 ) , .A2( u1_u2_u1_n156 ) );
  AND2_X1 u1_u2_u1_U22 (.A1( u1_u2_u1_n123 ) , .ZN( u1_u2_u1_n134 ) , .A2( u1_u2_u1_n161 ) );
  NAND2_X1 u1_u2_u1_U23 (.A2( u1_u2_u1_n115 ) , .A1( u1_u2_u1_n116 ) , .ZN( u1_u2_u1_n148 ) );
  NAND2_X1 u1_u2_u1_U24 (.A2( u1_u2_u1_n133 ) , .A1( u1_u2_u1_n135 ) , .ZN( u1_u2_u1_n159 ) );
  NAND2_X1 u1_u2_u1_U25 (.A2( u1_u2_u1_n115 ) , .A1( u1_u2_u1_n120 ) , .ZN( u1_u2_u1_n132 ) );
  INV_X1 u1_u2_u1_U26 (.A( u1_u2_u1_n154 ) , .ZN( u1_u2_u1_n178 ) );
  INV_X1 u1_u2_u1_U27 (.A( u1_u2_u1_n151 ) , .ZN( u1_u2_u1_n183 ) );
  AND2_X1 u1_u2_u1_U28 (.A1( u1_u2_u1_n129 ) , .A2( u1_u2_u1_n133 ) , .ZN( u1_u2_u1_n149 ) );
  INV_X1 u1_u2_u1_U29 (.A( u1_u2_u1_n131 ) , .ZN( u1_u2_u1_n180 ) );
  INV_X1 u1_u2_u1_U3 (.A( u1_u2_u1_n159 ) , .ZN( u1_u2_u1_n182 ) );
  OAI221_X1 u1_u2_u1_U30 (.A( u1_u2_u1_n119 ) , .C2( u1_u2_u1_n129 ) , .ZN( u1_u2_u1_n138 ) , .B2( u1_u2_u1_n152 ) , .C1( u1_u2_u1_n174 ) , .B1( u1_u2_u1_n187 ) );
  INV_X1 u1_u2_u1_U31 (.A( u1_u2_u1_n148 ) , .ZN( u1_u2_u1_n187 ) );
  AOI211_X1 u1_u2_u1_U32 (.B( u1_u2_u1_n117 ) , .A( u1_u2_u1_n118 ) , .ZN( u1_u2_u1_n119 ) , .C2( u1_u2_u1_n146 ) , .C1( u1_u2_u1_n159 ) );
  NOR2_X1 u1_u2_u1_U33 (.A1( u1_u2_u1_n168 ) , .A2( u1_u2_u1_n176 ) , .ZN( u1_u2_u1_n98 ) );
  AOI211_X1 u1_u2_u1_U34 (.B( u1_u2_u1_n162 ) , .A( u1_u2_u1_n163 ) , .C2( u1_u2_u1_n164 ) , .ZN( u1_u2_u1_n165 ) , .C1( u1_u2_u1_n171 ) );
  AOI21_X1 u1_u2_u1_U35 (.A( u1_u2_u1_n160 ) , .B2( u1_u2_u1_n161 ) , .ZN( u1_u2_u1_n162 ) , .B1( u1_u2_u1_n182 ) );
  OR2_X1 u1_u2_u1_U36 (.A2( u1_u2_u1_n157 ) , .A1( u1_u2_u1_n158 ) , .ZN( u1_u2_u1_n163 ) );
  OAI21_X1 u1_u2_u1_U37 (.B2( u1_u2_u1_n123 ) , .ZN( u1_u2_u1_n145 ) , .B1( u1_u2_u1_n160 ) , .A( u1_u2_u1_n185 ) );
  INV_X1 u1_u2_u1_U38 (.A( u1_u2_u1_n122 ) , .ZN( u1_u2_u1_n185 ) );
  AOI21_X1 u1_u2_u1_U39 (.B2( u1_u2_u1_n120 ) , .B1( u1_u2_u1_n121 ) , .ZN( u1_u2_u1_n122 ) , .A( u1_u2_u1_n128 ) );
  AOI221_X1 u1_u2_u1_U4 (.A( u1_u2_u1_n138 ) , .C2( u1_u2_u1_n139 ) , .C1( u1_u2_u1_n140 ) , .B2( u1_u2_u1_n141 ) , .ZN( u1_u2_u1_n142 ) , .B1( u1_u2_u1_n175 ) );
  NAND2_X1 u1_u2_u1_U40 (.A1( u1_u2_u1_n128 ) , .ZN( u1_u2_u1_n146 ) , .A2( u1_u2_u1_n160 ) );
  NAND2_X1 u1_u2_u1_U41 (.A2( u1_u2_u1_n112 ) , .ZN( u1_u2_u1_n139 ) , .A1( u1_u2_u1_n152 ) );
  NAND2_X1 u1_u2_u1_U42 (.A1( u1_u2_u1_n105 ) , .ZN( u1_u2_u1_n156 ) , .A2( u1_u2_u1_n99 ) );
  AOI221_X1 u1_u2_u1_U43 (.B1( u1_u2_u1_n140 ) , .ZN( u1_u2_u1_n167 ) , .B2( u1_u2_u1_n172 ) , .C2( u1_u2_u1_n175 ) , .C1( u1_u2_u1_n178 ) , .A( u1_u2_u1_n188 ) );
  INV_X1 u1_u2_u1_U44 (.ZN( u1_u2_u1_n188 ) , .A( u1_u2_u1_n97 ) );
  AOI211_X1 u1_u2_u1_U45 (.A( u1_u2_u1_n118 ) , .C1( u1_u2_u1_n132 ) , .C2( u1_u2_u1_n139 ) , .B( u1_u2_u1_n96 ) , .ZN( u1_u2_u1_n97 ) );
  AOI21_X1 u1_u2_u1_U46 (.B2( u1_u2_u1_n121 ) , .B1( u1_u2_u1_n135 ) , .A( u1_u2_u1_n152 ) , .ZN( u1_u2_u1_n96 ) );
  NOR2_X1 u1_u2_u1_U47 (.ZN( u1_u2_u1_n117 ) , .A1( u1_u2_u1_n121 ) , .A2( u1_u2_u1_n160 ) );
  AOI21_X1 u1_u2_u1_U48 (.A( u1_u2_u1_n128 ) , .B2( u1_u2_u1_n129 ) , .ZN( u1_u2_u1_n130 ) , .B1( u1_u2_u1_n150 ) );
  NAND2_X1 u1_u2_u1_U49 (.ZN( u1_u2_u1_n112 ) , .A1( u1_u2_u1_n169 ) , .A2( u1_u2_u1_n170 ) );
  AOI211_X1 u1_u2_u1_U5 (.ZN( u1_u2_u1_n124 ) , .A( u1_u2_u1_n138 ) , .C2( u1_u2_u1_n139 ) , .B( u1_u2_u1_n145 ) , .C1( u1_u2_u1_n147 ) );
  NAND2_X1 u1_u2_u1_U50 (.ZN( u1_u2_u1_n129 ) , .A2( u1_u2_u1_n95 ) , .A1( u1_u2_u1_n98 ) );
  NAND2_X1 u1_u2_u1_U51 (.A1( u1_u2_u1_n102 ) , .ZN( u1_u2_u1_n154 ) , .A2( u1_u2_u1_n99 ) );
  NAND2_X1 u1_u2_u1_U52 (.A2( u1_u2_u1_n100 ) , .ZN( u1_u2_u1_n135 ) , .A1( u1_u2_u1_n99 ) );
  AOI21_X1 u1_u2_u1_U53 (.A( u1_u2_u1_n152 ) , .B2( u1_u2_u1_n153 ) , .B1( u1_u2_u1_n154 ) , .ZN( u1_u2_u1_n158 ) );
  INV_X1 u1_u2_u1_U54 (.A( u1_u2_u1_n160 ) , .ZN( u1_u2_u1_n175 ) );
  NAND2_X1 u1_u2_u1_U55 (.A1( u1_u2_u1_n100 ) , .ZN( u1_u2_u1_n116 ) , .A2( u1_u2_u1_n95 ) );
  NAND2_X1 u1_u2_u1_U56 (.A1( u1_u2_u1_n102 ) , .ZN( u1_u2_u1_n131 ) , .A2( u1_u2_u1_n95 ) );
  NAND2_X1 u1_u2_u1_U57 (.A2( u1_u2_u1_n104 ) , .ZN( u1_u2_u1_n121 ) , .A1( u1_u2_u1_n98 ) );
  NAND2_X1 u1_u2_u1_U58 (.A1( u1_u2_u1_n103 ) , .ZN( u1_u2_u1_n153 ) , .A2( u1_u2_u1_n98 ) );
  NAND2_X1 u1_u2_u1_U59 (.A2( u1_u2_u1_n104 ) , .A1( u1_u2_u1_n105 ) , .ZN( u1_u2_u1_n133 ) );
  AOI22_X1 u1_u2_u1_U6 (.B2( u1_u2_u1_n113 ) , .A2( u1_u2_u1_n114 ) , .ZN( u1_u2_u1_n125 ) , .A1( u1_u2_u1_n171 ) , .B1( u1_u2_u1_n173 ) );
  NAND2_X1 u1_u2_u1_U60 (.ZN( u1_u2_u1_n150 ) , .A2( u1_u2_u1_n98 ) , .A1( u1_u2_u1_n99 ) );
  NAND2_X1 u1_u2_u1_U61 (.A1( u1_u2_u1_n105 ) , .ZN( u1_u2_u1_n155 ) , .A2( u1_u2_u1_n95 ) );
  OAI21_X1 u1_u2_u1_U62 (.ZN( u1_u2_u1_n109 ) , .B1( u1_u2_u1_n129 ) , .B2( u1_u2_u1_n160 ) , .A( u1_u2_u1_n167 ) );
  NAND2_X1 u1_u2_u1_U63 (.A2( u1_u2_u1_n100 ) , .A1( u1_u2_u1_n103 ) , .ZN( u1_u2_u1_n120 ) );
  NAND2_X1 u1_u2_u1_U64 (.A1( u1_u2_u1_n102 ) , .A2( u1_u2_u1_n104 ) , .ZN( u1_u2_u1_n115 ) );
  NAND2_X1 u1_u2_u1_U65 (.A2( u1_u2_u1_n100 ) , .A1( u1_u2_u1_n104 ) , .ZN( u1_u2_u1_n151 ) );
  NAND2_X1 u1_u2_u1_U66 (.A2( u1_u2_u1_n103 ) , .A1( u1_u2_u1_n105 ) , .ZN( u1_u2_u1_n161 ) );
  INV_X1 u1_u2_u1_U67 (.A( u1_u2_u1_n152 ) , .ZN( u1_u2_u1_n173 ) );
  INV_X1 u1_u2_u1_U68 (.A( u1_u2_u1_n128 ) , .ZN( u1_u2_u1_n172 ) );
  NAND2_X1 u1_u2_u1_U69 (.A2( u1_u2_u1_n102 ) , .A1( u1_u2_u1_n103 ) , .ZN( u1_u2_u1_n123 ) );
  NAND2_X1 u1_u2_u1_U7 (.ZN( u1_u2_u1_n114 ) , .A1( u1_u2_u1_n134 ) , .A2( u1_u2_u1_n156 ) );
  NOR2_X1 u1_u2_u1_U70 (.A2( u1_u2_X_7 ) , .A1( u1_u2_X_8 ) , .ZN( u1_u2_u1_n95 ) );
  NOR2_X1 u1_u2_u1_U71 (.A1( u1_u2_X_12 ) , .A2( u1_u2_X_9 ) , .ZN( u1_u2_u1_n100 ) );
  NOR2_X1 u1_u2_u1_U72 (.A2( u1_u2_X_8 ) , .A1( u1_u2_u1_n177 ) , .ZN( u1_u2_u1_n99 ) );
  NOR2_X1 u1_u2_u1_U73 (.A2( u1_u2_X_12 ) , .ZN( u1_u2_u1_n102 ) , .A1( u1_u2_u1_n176 ) );
  NOR2_X1 u1_u2_u1_U74 (.A2( u1_u2_X_9 ) , .ZN( u1_u2_u1_n105 ) , .A1( u1_u2_u1_n168 ) );
  NAND2_X1 u1_u2_u1_U75 (.A1( u1_u2_X_10 ) , .ZN( u1_u2_u1_n160 ) , .A2( u1_u2_u1_n169 ) );
  NAND2_X1 u1_u2_u1_U76 (.A2( u1_u2_X_10 ) , .A1( u1_u2_X_11 ) , .ZN( u1_u2_u1_n152 ) );
  NAND2_X1 u1_u2_u1_U77 (.A1( u1_u2_X_11 ) , .ZN( u1_u2_u1_n128 ) , .A2( u1_u2_u1_n170 ) );
  AND2_X1 u1_u2_u1_U78 (.A2( u1_u2_X_7 ) , .A1( u1_u2_X_8 ) , .ZN( u1_u2_u1_n104 ) );
  AND2_X1 u1_u2_u1_U79 (.A1( u1_u2_X_8 ) , .ZN( u1_u2_u1_n103 ) , .A2( u1_u2_u1_n177 ) );
  AOI22_X1 u1_u2_u1_U8 (.B2( u1_u2_u1_n136 ) , .A2( u1_u2_u1_n137 ) , .ZN( u1_u2_u1_n143 ) , .A1( u1_u2_u1_n171 ) , .B1( u1_u2_u1_n173 ) );
  INV_X1 u1_u2_u1_U80 (.A( u1_u2_X_10 ) , .ZN( u1_u2_u1_n170 ) );
  INV_X1 u1_u2_u1_U81 (.A( u1_u2_X_9 ) , .ZN( u1_u2_u1_n176 ) );
  INV_X1 u1_u2_u1_U82 (.A( u1_u2_X_11 ) , .ZN( u1_u2_u1_n169 ) );
  INV_X1 u1_u2_u1_U83 (.A( u1_u2_X_12 ) , .ZN( u1_u2_u1_n168 ) );
  INV_X1 u1_u2_u1_U84 (.A( u1_u2_X_7 ) , .ZN( u1_u2_u1_n177 ) );
  NAND4_X1 u1_u2_u1_U85 (.ZN( u1_out2_18 ) , .A4( u1_u2_u1_n165 ) , .A3( u1_u2_u1_n166 ) , .A1( u1_u2_u1_n167 ) , .A2( u1_u2_u1_n186 ) );
  AOI22_X1 u1_u2_u1_U86 (.B2( u1_u2_u1_n146 ) , .B1( u1_u2_u1_n147 ) , .A2( u1_u2_u1_n148 ) , .ZN( u1_u2_u1_n166 ) , .A1( u1_u2_u1_n172 ) );
  INV_X1 u1_u2_u1_U87 (.A( u1_u2_u1_n145 ) , .ZN( u1_u2_u1_n186 ) );
  NAND4_X1 u1_u2_u1_U88 (.ZN( u1_out2_2 ) , .A4( u1_u2_u1_n142 ) , .A3( u1_u2_u1_n143 ) , .A2( u1_u2_u1_n144 ) , .A1( u1_u2_u1_n179 ) );
  OAI21_X1 u1_u2_u1_U89 (.B2( u1_u2_u1_n132 ) , .ZN( u1_u2_u1_n144 ) , .A( u1_u2_u1_n146 ) , .B1( u1_u2_u1_n180 ) );
  INV_X1 u1_u2_u1_U9 (.A( u1_u2_u1_n147 ) , .ZN( u1_u2_u1_n181 ) );
  INV_X1 u1_u2_u1_U90 (.A( u1_u2_u1_n130 ) , .ZN( u1_u2_u1_n179 ) );
  NAND4_X1 u1_u2_u1_U91 (.ZN( u1_out2_28 ) , .A4( u1_u2_u1_n124 ) , .A3( u1_u2_u1_n125 ) , .A2( u1_u2_u1_n126 ) , .A1( u1_u2_u1_n127 ) );
  OAI21_X1 u1_u2_u1_U92 (.ZN( u1_u2_u1_n127 ) , .B2( u1_u2_u1_n139 ) , .B1( u1_u2_u1_n175 ) , .A( u1_u2_u1_n183 ) );
  OAI21_X1 u1_u2_u1_U93 (.ZN( u1_u2_u1_n126 ) , .B2( u1_u2_u1_n140 ) , .A( u1_u2_u1_n146 ) , .B1( u1_u2_u1_n178 ) );
  OR4_X1 u1_u2_u1_U94 (.ZN( u1_out2_13 ) , .A4( u1_u2_u1_n108 ) , .A3( u1_u2_u1_n109 ) , .A2( u1_u2_u1_n110 ) , .A1( u1_u2_u1_n111 ) );
  AOI21_X1 u1_u2_u1_U95 (.ZN( u1_u2_u1_n111 ) , .A( u1_u2_u1_n128 ) , .B2( u1_u2_u1_n131 ) , .B1( u1_u2_u1_n135 ) );
  AOI21_X1 u1_u2_u1_U96 (.ZN( u1_u2_u1_n110 ) , .A( u1_u2_u1_n116 ) , .B1( u1_u2_u1_n152 ) , .B2( u1_u2_u1_n160 ) );
  NAND3_X1 u1_u2_u1_U97 (.A3( u1_u2_u1_n149 ) , .A2( u1_u2_u1_n150 ) , .A1( u1_u2_u1_n151 ) , .ZN( u1_u2_u1_n164 ) );
  NAND3_X1 u1_u2_u1_U98 (.A3( u1_u2_u1_n134 ) , .A2( u1_u2_u1_n135 ) , .ZN( u1_u2_u1_n136 ) , .A1( u1_u2_u1_n151 ) );
  NAND3_X1 u1_u2_u1_U99 (.A1( u1_u2_u1_n133 ) , .ZN( u1_u2_u1_n137 ) , .A2( u1_u2_u1_n154 ) , .A3( u1_u2_u1_n181 ) );
  XOR2_X1 u1_u3_U10 (.B( u1_K4_45 ) , .A( u1_R2_30 ) , .Z( u1_u3_X_45 ) );
  XOR2_X1 u1_u3_U9 (.B( u1_K4_46 ) , .A( u1_R2_31 ) , .Z( u1_u3_X_46 ) );
  AND3_X1 u1_u3_u7_U10 (.A3( u1_u3_u7_n110 ) , .A2( u1_u3_u7_n127 ) , .A1( u1_u3_u7_n132 ) , .ZN( u1_u3_u7_n92 ) );
  OAI21_X1 u1_u3_u7_U11 (.A( u1_u3_u7_n161 ) , .B1( u1_u3_u7_n168 ) , .B2( u1_u3_u7_n173 ) , .ZN( u1_u3_u7_n91 ) );
  AOI211_X1 u1_u3_u7_U12 (.A( u1_u3_u7_n117 ) , .ZN( u1_u3_u7_n118 ) , .C2( u1_u3_u7_n126 ) , .C1( u1_u3_u7_n177 ) , .B( u1_u3_u7_n180 ) );
  OAI22_X1 u1_u3_u7_U13 (.B1( u1_u3_u7_n115 ) , .ZN( u1_u3_u7_n117 ) , .A2( u1_u3_u7_n133 ) , .A1( u1_u3_u7_n137 ) , .B2( u1_u3_u7_n162 ) );
  INV_X1 u1_u3_u7_U14 (.A( u1_u3_u7_n116 ) , .ZN( u1_u3_u7_n180 ) );
  NOR3_X1 u1_u3_u7_U15 (.ZN( u1_u3_u7_n115 ) , .A3( u1_u3_u7_n145 ) , .A2( u1_u3_u7_n168 ) , .A1( u1_u3_u7_n169 ) );
  OAI211_X1 u1_u3_u7_U16 (.B( u1_u3_u7_n122 ) , .A( u1_u3_u7_n123 ) , .C2( u1_u3_u7_n124 ) , .ZN( u1_u3_u7_n154 ) , .C1( u1_u3_u7_n162 ) );
  AOI222_X1 u1_u3_u7_U17 (.ZN( u1_u3_u7_n122 ) , .C2( u1_u3_u7_n126 ) , .C1( u1_u3_u7_n145 ) , .B1( u1_u3_u7_n161 ) , .A2( u1_u3_u7_n165 ) , .B2( u1_u3_u7_n170 ) , .A1( u1_u3_u7_n176 ) );
  INV_X1 u1_u3_u7_U18 (.A( u1_u3_u7_n133 ) , .ZN( u1_u3_u7_n176 ) );
  NOR3_X1 u1_u3_u7_U19 (.A2( u1_u3_u7_n134 ) , .A1( u1_u3_u7_n135 ) , .ZN( u1_u3_u7_n136 ) , .A3( u1_u3_u7_n171 ) );
  NOR2_X1 u1_u3_u7_U20 (.A1( u1_u3_u7_n130 ) , .A2( u1_u3_u7_n134 ) , .ZN( u1_u3_u7_n153 ) );
  INV_X1 u1_u3_u7_U21 (.A( u1_u3_u7_n101 ) , .ZN( u1_u3_u7_n165 ) );
  NOR2_X1 u1_u3_u7_U22 (.ZN( u1_u3_u7_n111 ) , .A2( u1_u3_u7_n134 ) , .A1( u1_u3_u7_n169 ) );
  AOI21_X1 u1_u3_u7_U23 (.ZN( u1_u3_u7_n104 ) , .B2( u1_u3_u7_n112 ) , .B1( u1_u3_u7_n127 ) , .A( u1_u3_u7_n164 ) );
  AOI21_X1 u1_u3_u7_U24 (.ZN( u1_u3_u7_n106 ) , .B1( u1_u3_u7_n133 ) , .B2( u1_u3_u7_n146 ) , .A( u1_u3_u7_n162 ) );
  AOI21_X1 u1_u3_u7_U25 (.A( u1_u3_u7_n101 ) , .ZN( u1_u3_u7_n107 ) , .B2( u1_u3_u7_n128 ) , .B1( u1_u3_u7_n175 ) );
  INV_X1 u1_u3_u7_U26 (.A( u1_u3_u7_n138 ) , .ZN( u1_u3_u7_n171 ) );
  INV_X1 u1_u3_u7_U27 (.A( u1_u3_u7_n131 ) , .ZN( u1_u3_u7_n177 ) );
  INV_X1 u1_u3_u7_U28 (.A( u1_u3_u7_n110 ) , .ZN( u1_u3_u7_n174 ) );
  NAND2_X1 u1_u3_u7_U29 (.A1( u1_u3_u7_n129 ) , .A2( u1_u3_u7_n132 ) , .ZN( u1_u3_u7_n149 ) );
  OAI21_X1 u1_u3_u7_U3 (.ZN( u1_u3_u7_n159 ) , .A( u1_u3_u7_n165 ) , .B2( u1_u3_u7_n171 ) , .B1( u1_u3_u7_n174 ) );
  NAND2_X1 u1_u3_u7_U30 (.A1( u1_u3_u7_n113 ) , .A2( u1_u3_u7_n124 ) , .ZN( u1_u3_u7_n130 ) );
  INV_X1 u1_u3_u7_U31 (.A( u1_u3_u7_n112 ) , .ZN( u1_u3_u7_n173 ) );
  INV_X1 u1_u3_u7_U32 (.A( u1_u3_u7_n128 ) , .ZN( u1_u3_u7_n168 ) );
  INV_X1 u1_u3_u7_U33 (.A( u1_u3_u7_n148 ) , .ZN( u1_u3_u7_n169 ) );
  INV_X1 u1_u3_u7_U34 (.A( u1_u3_u7_n127 ) , .ZN( u1_u3_u7_n179 ) );
  NOR2_X1 u1_u3_u7_U35 (.ZN( u1_u3_u7_n101 ) , .A2( u1_u3_u7_n150 ) , .A1( u1_u3_u7_n156 ) );
  AOI211_X1 u1_u3_u7_U36 (.B( u1_u3_u7_n154 ) , .A( u1_u3_u7_n155 ) , .C1( u1_u3_u7_n156 ) , .ZN( u1_u3_u7_n157 ) , .C2( u1_u3_u7_n172 ) );
  INV_X1 u1_u3_u7_U37 (.A( u1_u3_u7_n153 ) , .ZN( u1_u3_u7_n172 ) );
  AOI211_X1 u1_u3_u7_U38 (.B( u1_u3_u7_n139 ) , .A( u1_u3_u7_n140 ) , .C2( u1_u3_u7_n141 ) , .ZN( u1_u3_u7_n142 ) , .C1( u1_u3_u7_n156 ) );
  NAND4_X1 u1_u3_u7_U39 (.A3( u1_u3_u7_n127 ) , .A2( u1_u3_u7_n128 ) , .A1( u1_u3_u7_n129 ) , .ZN( u1_u3_u7_n141 ) , .A4( u1_u3_u7_n147 ) );
  INV_X1 u1_u3_u7_U4 (.A( u1_u3_u7_n111 ) , .ZN( u1_u3_u7_n170 ) );
  AOI21_X1 u1_u3_u7_U40 (.A( u1_u3_u7_n137 ) , .B1( u1_u3_u7_n138 ) , .ZN( u1_u3_u7_n139 ) , .B2( u1_u3_u7_n146 ) );
  OAI22_X1 u1_u3_u7_U41 (.B1( u1_u3_u7_n136 ) , .ZN( u1_u3_u7_n140 ) , .A1( u1_u3_u7_n153 ) , .B2( u1_u3_u7_n162 ) , .A2( u1_u3_u7_n164 ) );
  AOI21_X1 u1_u3_u7_U42 (.ZN( u1_u3_u7_n123 ) , .B1( u1_u3_u7_n165 ) , .B2( u1_u3_u7_n177 ) , .A( u1_u3_u7_n97 ) );
  AOI21_X1 u1_u3_u7_U43 (.B2( u1_u3_u7_n113 ) , .B1( u1_u3_u7_n124 ) , .A( u1_u3_u7_n125 ) , .ZN( u1_u3_u7_n97 ) );
  INV_X1 u1_u3_u7_U44 (.A( u1_u3_u7_n125 ) , .ZN( u1_u3_u7_n161 ) );
  INV_X1 u1_u3_u7_U45 (.A( u1_u3_u7_n152 ) , .ZN( u1_u3_u7_n162 ) );
  AOI22_X1 u1_u3_u7_U46 (.A2( u1_u3_u7_n114 ) , .ZN( u1_u3_u7_n119 ) , .B1( u1_u3_u7_n130 ) , .A1( u1_u3_u7_n156 ) , .B2( u1_u3_u7_n165 ) );
  NAND2_X1 u1_u3_u7_U47 (.A2( u1_u3_u7_n112 ) , .ZN( u1_u3_u7_n114 ) , .A1( u1_u3_u7_n175 ) );
  AND2_X1 u1_u3_u7_U48 (.ZN( u1_u3_u7_n145 ) , .A2( u1_u3_u7_n98 ) , .A1( u1_u3_u7_n99 ) );
  NOR2_X1 u1_u3_u7_U49 (.ZN( u1_u3_u7_n137 ) , .A1( u1_u3_u7_n150 ) , .A2( u1_u3_u7_n161 ) );
  INV_X1 u1_u3_u7_U5 (.A( u1_u3_u7_n149 ) , .ZN( u1_u3_u7_n175 ) );
  AOI21_X1 u1_u3_u7_U50 (.ZN( u1_u3_u7_n105 ) , .B2( u1_u3_u7_n110 ) , .A( u1_u3_u7_n125 ) , .B1( u1_u3_u7_n147 ) );
  NAND2_X1 u1_u3_u7_U51 (.ZN( u1_u3_u7_n146 ) , .A1( u1_u3_u7_n95 ) , .A2( u1_u3_u7_n98 ) );
  NAND2_X1 u1_u3_u7_U52 (.A2( u1_u3_u7_n103 ) , .ZN( u1_u3_u7_n147 ) , .A1( u1_u3_u7_n93 ) );
  NAND2_X1 u1_u3_u7_U53 (.A1( u1_u3_u7_n103 ) , .ZN( u1_u3_u7_n127 ) , .A2( u1_u3_u7_n99 ) );
  OR2_X1 u1_u3_u7_U54 (.ZN( u1_u3_u7_n126 ) , .A2( u1_u3_u7_n152 ) , .A1( u1_u3_u7_n156 ) );
  NAND2_X1 u1_u3_u7_U55 (.A2( u1_u3_u7_n102 ) , .A1( u1_u3_u7_n103 ) , .ZN( u1_u3_u7_n133 ) );
  NAND2_X1 u1_u3_u7_U56 (.ZN( u1_u3_u7_n112 ) , .A2( u1_u3_u7_n96 ) , .A1( u1_u3_u7_n99 ) );
  NAND2_X1 u1_u3_u7_U57 (.A2( u1_u3_u7_n102 ) , .ZN( u1_u3_u7_n128 ) , .A1( u1_u3_u7_n98 ) );
  NAND2_X1 u1_u3_u7_U58 (.A1( u1_u3_u7_n100 ) , .ZN( u1_u3_u7_n113 ) , .A2( u1_u3_u7_n93 ) );
  NAND2_X1 u1_u3_u7_U59 (.A2( u1_u3_u7_n102 ) , .ZN( u1_u3_u7_n124 ) , .A1( u1_u3_u7_n96 ) );
  INV_X1 u1_u3_u7_U6 (.A( u1_u3_u7_n154 ) , .ZN( u1_u3_u7_n178 ) );
  NAND2_X1 u1_u3_u7_U60 (.ZN( u1_u3_u7_n110 ) , .A1( u1_u3_u7_n95 ) , .A2( u1_u3_u7_n96 ) );
  INV_X1 u1_u3_u7_U61 (.A( u1_u3_u7_n150 ) , .ZN( u1_u3_u7_n164 ) );
  AND2_X1 u1_u3_u7_U62 (.ZN( u1_u3_u7_n134 ) , .A1( u1_u3_u7_n93 ) , .A2( u1_u3_u7_n98 ) );
  NAND2_X1 u1_u3_u7_U63 (.A1( u1_u3_u7_n100 ) , .A2( u1_u3_u7_n102 ) , .ZN( u1_u3_u7_n129 ) );
  NAND2_X1 u1_u3_u7_U64 (.A2( u1_u3_u7_n103 ) , .ZN( u1_u3_u7_n131 ) , .A1( u1_u3_u7_n95 ) );
  NAND2_X1 u1_u3_u7_U65 (.A1( u1_u3_u7_n100 ) , .ZN( u1_u3_u7_n138 ) , .A2( u1_u3_u7_n99 ) );
  NAND2_X1 u1_u3_u7_U66 (.ZN( u1_u3_u7_n132 ) , .A1( u1_u3_u7_n93 ) , .A2( u1_u3_u7_n96 ) );
  NAND2_X1 u1_u3_u7_U67 (.A1( u1_u3_u7_n100 ) , .ZN( u1_u3_u7_n148 ) , .A2( u1_u3_u7_n95 ) );
  NOR2_X1 u1_u3_u7_U68 (.A2( u1_u3_X_47 ) , .ZN( u1_u3_u7_n150 ) , .A1( u1_u3_u7_n163 ) );
  NOR2_X1 u1_u3_u7_U69 (.A2( u1_u3_X_43 ) , .A1( u1_u3_X_44 ) , .ZN( u1_u3_u7_n103 ) );
  AOI211_X1 u1_u3_u7_U7 (.ZN( u1_u3_u7_n116 ) , .A( u1_u3_u7_n155 ) , .C1( u1_u3_u7_n161 ) , .C2( u1_u3_u7_n171 ) , .B( u1_u3_u7_n94 ) );
  NOR2_X1 u1_u3_u7_U70 (.A2( u1_u3_X_48 ) , .A1( u1_u3_u7_n166 ) , .ZN( u1_u3_u7_n95 ) );
  NOR2_X1 u1_u3_u7_U71 (.A2( u1_u3_X_45 ) , .A1( u1_u3_X_48 ) , .ZN( u1_u3_u7_n99 ) );
  NOR2_X1 u1_u3_u7_U72 (.A2( u1_u3_X_44 ) , .A1( u1_u3_u7_n167 ) , .ZN( u1_u3_u7_n98 ) );
  NOR2_X1 u1_u3_u7_U73 (.A2( u1_u3_X_46 ) , .A1( u1_u3_X_47 ) , .ZN( u1_u3_u7_n152 ) );
  AND2_X1 u1_u3_u7_U74 (.A1( u1_u3_X_47 ) , .ZN( u1_u3_u7_n156 ) , .A2( u1_u3_u7_n163 ) );
  NAND2_X1 u1_u3_u7_U75 (.A2( u1_u3_X_46 ) , .A1( u1_u3_X_47 ) , .ZN( u1_u3_u7_n125 ) );
  AND2_X1 u1_u3_u7_U76 (.A2( u1_u3_X_45 ) , .A1( u1_u3_X_48 ) , .ZN( u1_u3_u7_n102 ) );
  AND2_X1 u1_u3_u7_U77 (.A2( u1_u3_X_43 ) , .A1( u1_u3_X_44 ) , .ZN( u1_u3_u7_n96 ) );
  AND2_X1 u1_u3_u7_U78 (.A1( u1_u3_X_44 ) , .ZN( u1_u3_u7_n100 ) , .A2( u1_u3_u7_n167 ) );
  AND2_X1 u1_u3_u7_U79 (.A1( u1_u3_X_48 ) , .A2( u1_u3_u7_n166 ) , .ZN( u1_u3_u7_n93 ) );
  OAI222_X1 u1_u3_u7_U8 (.C2( u1_u3_u7_n101 ) , .B2( u1_u3_u7_n111 ) , .A1( u1_u3_u7_n113 ) , .C1( u1_u3_u7_n146 ) , .A2( u1_u3_u7_n162 ) , .B1( u1_u3_u7_n164 ) , .ZN( u1_u3_u7_n94 ) );
  INV_X1 u1_u3_u7_U80 (.A( u1_u3_X_46 ) , .ZN( u1_u3_u7_n163 ) );
  INV_X1 u1_u3_u7_U81 (.A( u1_u3_X_43 ) , .ZN( u1_u3_u7_n167 ) );
  INV_X1 u1_u3_u7_U82 (.A( u1_u3_X_45 ) , .ZN( u1_u3_u7_n166 ) );
  NAND4_X1 u1_u3_u7_U83 (.ZN( u1_out3_5 ) , .A4( u1_u3_u7_n108 ) , .A3( u1_u3_u7_n109 ) , .A1( u1_u3_u7_n116 ) , .A2( u1_u3_u7_n123 ) );
  AOI22_X1 u1_u3_u7_U84 (.ZN( u1_u3_u7_n109 ) , .A2( u1_u3_u7_n126 ) , .B2( u1_u3_u7_n145 ) , .B1( u1_u3_u7_n156 ) , .A1( u1_u3_u7_n171 ) );
  NOR4_X1 u1_u3_u7_U85 (.A4( u1_u3_u7_n104 ) , .A3( u1_u3_u7_n105 ) , .A2( u1_u3_u7_n106 ) , .A1( u1_u3_u7_n107 ) , .ZN( u1_u3_u7_n108 ) );
  NAND4_X1 u1_u3_u7_U86 (.ZN( u1_out3_27 ) , .A4( u1_u3_u7_n118 ) , .A3( u1_u3_u7_n119 ) , .A2( u1_u3_u7_n120 ) , .A1( u1_u3_u7_n121 ) );
  OAI21_X1 u1_u3_u7_U87 (.ZN( u1_u3_u7_n121 ) , .B2( u1_u3_u7_n145 ) , .A( u1_u3_u7_n150 ) , .B1( u1_u3_u7_n174 ) );
  OAI21_X1 u1_u3_u7_U88 (.ZN( u1_u3_u7_n120 ) , .A( u1_u3_u7_n161 ) , .B2( u1_u3_u7_n170 ) , .B1( u1_u3_u7_n179 ) );
  NAND4_X1 u1_u3_u7_U89 (.ZN( u1_out3_21 ) , .A4( u1_u3_u7_n157 ) , .A3( u1_u3_u7_n158 ) , .A2( u1_u3_u7_n159 ) , .A1( u1_u3_u7_n160 ) );
  OAI221_X1 u1_u3_u7_U9 (.C1( u1_u3_u7_n101 ) , .C2( u1_u3_u7_n147 ) , .ZN( u1_u3_u7_n155 ) , .B2( u1_u3_u7_n162 ) , .A( u1_u3_u7_n91 ) , .B1( u1_u3_u7_n92 ) );
  OAI21_X1 u1_u3_u7_U90 (.B1( u1_u3_u7_n145 ) , .ZN( u1_u3_u7_n160 ) , .A( u1_u3_u7_n161 ) , .B2( u1_u3_u7_n177 ) );
  AOI22_X1 u1_u3_u7_U91 (.B2( u1_u3_u7_n149 ) , .B1( u1_u3_u7_n150 ) , .A2( u1_u3_u7_n151 ) , .A1( u1_u3_u7_n152 ) , .ZN( u1_u3_u7_n158 ) );
  NAND4_X1 u1_u3_u7_U92 (.ZN( u1_out3_15 ) , .A4( u1_u3_u7_n142 ) , .A3( u1_u3_u7_n143 ) , .A2( u1_u3_u7_n144 ) , .A1( u1_u3_u7_n178 ) );
  OR2_X1 u1_u3_u7_U93 (.A2( u1_u3_u7_n125 ) , .A1( u1_u3_u7_n129 ) , .ZN( u1_u3_u7_n144 ) );
  AOI22_X1 u1_u3_u7_U94 (.A2( u1_u3_u7_n126 ) , .ZN( u1_u3_u7_n143 ) , .B2( u1_u3_u7_n165 ) , .B1( u1_u3_u7_n173 ) , .A1( u1_u3_u7_n174 ) );
  NAND3_X1 u1_u3_u7_U95 (.A3( u1_u3_u7_n146 ) , .A2( u1_u3_u7_n147 ) , .A1( u1_u3_u7_n148 ) , .ZN( u1_u3_u7_n151 ) );
  NAND3_X1 u1_u3_u7_U96 (.A3( u1_u3_u7_n131 ) , .A2( u1_u3_u7_n132 ) , .A1( u1_u3_u7_n133 ) , .ZN( u1_u3_u7_n135 ) );
  XOR2_X1 u1_u4_U1 (.B( u1_K5_9 ) , .A( u1_R3_6 ) , .Z( u1_u4_X_9 ) );
  XOR2_X1 u1_u4_U48 (.B( u1_K5_10 ) , .A( u1_R3_7 ) , .Z( u1_u4_X_10 ) );
  NOR2_X1 u1_u4_u1_U10 (.A1( u1_u4_u1_n112 ) , .A2( u1_u4_u1_n116 ) , .ZN( u1_u4_u1_n118 ) );
  NAND3_X1 u1_u4_u1_U100 (.ZN( u1_u4_u1_n113 ) , .A1( u1_u4_u1_n120 ) , .A3( u1_u4_u1_n133 ) , .A2( u1_u4_u1_n155 ) );
  OAI21_X1 u1_u4_u1_U11 (.ZN( u1_u4_u1_n101 ) , .B1( u1_u4_u1_n141 ) , .A( u1_u4_u1_n146 ) , .B2( u1_u4_u1_n183 ) );
  AOI21_X1 u1_u4_u1_U12 (.B2( u1_u4_u1_n155 ) , .B1( u1_u4_u1_n156 ) , .ZN( u1_u4_u1_n157 ) , .A( u1_u4_u1_n174 ) );
  NAND2_X1 u1_u4_u1_U13 (.ZN( u1_u4_u1_n140 ) , .A2( u1_u4_u1_n150 ) , .A1( u1_u4_u1_n155 ) );
  NAND2_X1 u1_u4_u1_U14 (.A1( u1_u4_u1_n131 ) , .ZN( u1_u4_u1_n147 ) , .A2( u1_u4_u1_n153 ) );
  INV_X1 u1_u4_u1_U15 (.A( u1_u4_u1_n139 ) , .ZN( u1_u4_u1_n174 ) );
  OR4_X1 u1_u4_u1_U16 (.A4( u1_u4_u1_n106 ) , .A3( u1_u4_u1_n107 ) , .ZN( u1_u4_u1_n108 ) , .A1( u1_u4_u1_n117 ) , .A2( u1_u4_u1_n184 ) );
  AOI21_X1 u1_u4_u1_U17 (.ZN( u1_u4_u1_n106 ) , .A( u1_u4_u1_n112 ) , .B1( u1_u4_u1_n154 ) , .B2( u1_u4_u1_n156 ) );
  AOI21_X1 u1_u4_u1_U18 (.ZN( u1_u4_u1_n107 ) , .B1( u1_u4_u1_n134 ) , .B2( u1_u4_u1_n149 ) , .A( u1_u4_u1_n174 ) );
  INV_X1 u1_u4_u1_U19 (.A( u1_u4_u1_n101 ) , .ZN( u1_u4_u1_n184 ) );
  INV_X1 u1_u4_u1_U20 (.A( u1_u4_u1_n112 ) , .ZN( u1_u4_u1_n171 ) );
  NAND2_X1 u1_u4_u1_U21 (.ZN( u1_u4_u1_n141 ) , .A1( u1_u4_u1_n153 ) , .A2( u1_u4_u1_n156 ) );
  AND2_X1 u1_u4_u1_U22 (.A1( u1_u4_u1_n123 ) , .ZN( u1_u4_u1_n134 ) , .A2( u1_u4_u1_n161 ) );
  NAND2_X1 u1_u4_u1_U23 (.A2( u1_u4_u1_n115 ) , .A1( u1_u4_u1_n116 ) , .ZN( u1_u4_u1_n148 ) );
  NAND2_X1 u1_u4_u1_U24 (.A2( u1_u4_u1_n133 ) , .A1( u1_u4_u1_n135 ) , .ZN( u1_u4_u1_n159 ) );
  NAND2_X1 u1_u4_u1_U25 (.A2( u1_u4_u1_n115 ) , .A1( u1_u4_u1_n120 ) , .ZN( u1_u4_u1_n132 ) );
  INV_X1 u1_u4_u1_U26 (.A( u1_u4_u1_n154 ) , .ZN( u1_u4_u1_n178 ) );
  INV_X1 u1_u4_u1_U27 (.A( u1_u4_u1_n151 ) , .ZN( u1_u4_u1_n183 ) );
  AND2_X1 u1_u4_u1_U28 (.A1( u1_u4_u1_n129 ) , .A2( u1_u4_u1_n133 ) , .ZN( u1_u4_u1_n149 ) );
  INV_X1 u1_u4_u1_U29 (.A( u1_u4_u1_n131 ) , .ZN( u1_u4_u1_n180 ) );
  INV_X1 u1_u4_u1_U3 (.A( u1_u4_u1_n159 ) , .ZN( u1_u4_u1_n182 ) );
  OAI221_X1 u1_u4_u1_U30 (.A( u1_u4_u1_n119 ) , .C2( u1_u4_u1_n129 ) , .ZN( u1_u4_u1_n138 ) , .B2( u1_u4_u1_n152 ) , .C1( u1_u4_u1_n174 ) , .B1( u1_u4_u1_n187 ) );
  INV_X1 u1_u4_u1_U31 (.A( u1_u4_u1_n148 ) , .ZN( u1_u4_u1_n187 ) );
  AOI211_X1 u1_u4_u1_U32 (.B( u1_u4_u1_n117 ) , .A( u1_u4_u1_n118 ) , .ZN( u1_u4_u1_n119 ) , .C2( u1_u4_u1_n146 ) , .C1( u1_u4_u1_n159 ) );
  NOR2_X1 u1_u4_u1_U33 (.A1( u1_u4_u1_n168 ) , .A2( u1_u4_u1_n176 ) , .ZN( u1_u4_u1_n98 ) );
  AOI211_X1 u1_u4_u1_U34 (.B( u1_u4_u1_n162 ) , .A( u1_u4_u1_n163 ) , .C2( u1_u4_u1_n164 ) , .ZN( u1_u4_u1_n165 ) , .C1( u1_u4_u1_n171 ) );
  AOI21_X1 u1_u4_u1_U35 (.A( u1_u4_u1_n160 ) , .B2( u1_u4_u1_n161 ) , .ZN( u1_u4_u1_n162 ) , .B1( u1_u4_u1_n182 ) );
  OR2_X1 u1_u4_u1_U36 (.A2( u1_u4_u1_n157 ) , .A1( u1_u4_u1_n158 ) , .ZN( u1_u4_u1_n163 ) );
  NAND2_X1 u1_u4_u1_U37 (.A1( u1_u4_u1_n128 ) , .ZN( u1_u4_u1_n146 ) , .A2( u1_u4_u1_n160 ) );
  NAND2_X1 u1_u4_u1_U38 (.A2( u1_u4_u1_n112 ) , .ZN( u1_u4_u1_n139 ) , .A1( u1_u4_u1_n152 ) );
  NAND2_X1 u1_u4_u1_U39 (.A1( u1_u4_u1_n105 ) , .ZN( u1_u4_u1_n156 ) , .A2( u1_u4_u1_n99 ) );
  AOI221_X1 u1_u4_u1_U4 (.A( u1_u4_u1_n138 ) , .C2( u1_u4_u1_n139 ) , .C1( u1_u4_u1_n140 ) , .B2( u1_u4_u1_n141 ) , .ZN( u1_u4_u1_n142 ) , .B1( u1_u4_u1_n175 ) );
  AOI221_X1 u1_u4_u1_U40 (.B1( u1_u4_u1_n140 ) , .ZN( u1_u4_u1_n167 ) , .B2( u1_u4_u1_n172 ) , .C2( u1_u4_u1_n175 ) , .C1( u1_u4_u1_n178 ) , .A( u1_u4_u1_n188 ) );
  INV_X1 u1_u4_u1_U41 (.ZN( u1_u4_u1_n188 ) , .A( u1_u4_u1_n97 ) );
  AOI211_X1 u1_u4_u1_U42 (.A( u1_u4_u1_n118 ) , .C1( u1_u4_u1_n132 ) , .C2( u1_u4_u1_n139 ) , .B( u1_u4_u1_n96 ) , .ZN( u1_u4_u1_n97 ) );
  AOI21_X1 u1_u4_u1_U43 (.B2( u1_u4_u1_n121 ) , .B1( u1_u4_u1_n135 ) , .A( u1_u4_u1_n152 ) , .ZN( u1_u4_u1_n96 ) );
  NOR2_X1 u1_u4_u1_U44 (.ZN( u1_u4_u1_n117 ) , .A1( u1_u4_u1_n121 ) , .A2( u1_u4_u1_n160 ) );
  OAI21_X1 u1_u4_u1_U45 (.B2( u1_u4_u1_n123 ) , .ZN( u1_u4_u1_n145 ) , .B1( u1_u4_u1_n160 ) , .A( u1_u4_u1_n185 ) );
  INV_X1 u1_u4_u1_U46 (.A( u1_u4_u1_n122 ) , .ZN( u1_u4_u1_n185 ) );
  AOI21_X1 u1_u4_u1_U47 (.B2( u1_u4_u1_n120 ) , .B1( u1_u4_u1_n121 ) , .ZN( u1_u4_u1_n122 ) , .A( u1_u4_u1_n128 ) );
  AOI21_X1 u1_u4_u1_U48 (.A( u1_u4_u1_n128 ) , .B2( u1_u4_u1_n129 ) , .ZN( u1_u4_u1_n130 ) , .B1( u1_u4_u1_n150 ) );
  NAND2_X1 u1_u4_u1_U49 (.ZN( u1_u4_u1_n112 ) , .A1( u1_u4_u1_n169 ) , .A2( u1_u4_u1_n170 ) );
  AOI211_X1 u1_u4_u1_U5 (.ZN( u1_u4_u1_n124 ) , .A( u1_u4_u1_n138 ) , .C2( u1_u4_u1_n139 ) , .B( u1_u4_u1_n145 ) , .C1( u1_u4_u1_n147 ) );
  NAND2_X1 u1_u4_u1_U50 (.ZN( u1_u4_u1_n129 ) , .A2( u1_u4_u1_n95 ) , .A1( u1_u4_u1_n98 ) );
  NAND2_X1 u1_u4_u1_U51 (.A1( u1_u4_u1_n102 ) , .ZN( u1_u4_u1_n154 ) , .A2( u1_u4_u1_n99 ) );
  NAND2_X1 u1_u4_u1_U52 (.A2( u1_u4_u1_n100 ) , .ZN( u1_u4_u1_n135 ) , .A1( u1_u4_u1_n99 ) );
  AOI21_X1 u1_u4_u1_U53 (.A( u1_u4_u1_n152 ) , .B2( u1_u4_u1_n153 ) , .B1( u1_u4_u1_n154 ) , .ZN( u1_u4_u1_n158 ) );
  INV_X1 u1_u4_u1_U54 (.A( u1_u4_u1_n160 ) , .ZN( u1_u4_u1_n175 ) );
  NAND2_X1 u1_u4_u1_U55 (.A1( u1_u4_u1_n100 ) , .ZN( u1_u4_u1_n116 ) , .A2( u1_u4_u1_n95 ) );
  NAND2_X1 u1_u4_u1_U56 (.A1( u1_u4_u1_n102 ) , .ZN( u1_u4_u1_n131 ) , .A2( u1_u4_u1_n95 ) );
  NAND2_X1 u1_u4_u1_U57 (.A2( u1_u4_u1_n104 ) , .ZN( u1_u4_u1_n121 ) , .A1( u1_u4_u1_n98 ) );
  NAND2_X1 u1_u4_u1_U58 (.A1( u1_u4_u1_n103 ) , .ZN( u1_u4_u1_n153 ) , .A2( u1_u4_u1_n98 ) );
  NAND2_X1 u1_u4_u1_U59 (.A2( u1_u4_u1_n104 ) , .A1( u1_u4_u1_n105 ) , .ZN( u1_u4_u1_n133 ) );
  AOI22_X1 u1_u4_u1_U6 (.B2( u1_u4_u1_n113 ) , .A2( u1_u4_u1_n114 ) , .ZN( u1_u4_u1_n125 ) , .A1( u1_u4_u1_n171 ) , .B1( u1_u4_u1_n173 ) );
  NAND2_X1 u1_u4_u1_U60 (.ZN( u1_u4_u1_n150 ) , .A2( u1_u4_u1_n98 ) , .A1( u1_u4_u1_n99 ) );
  NAND2_X1 u1_u4_u1_U61 (.A1( u1_u4_u1_n105 ) , .ZN( u1_u4_u1_n155 ) , .A2( u1_u4_u1_n95 ) );
  OAI21_X1 u1_u4_u1_U62 (.ZN( u1_u4_u1_n109 ) , .B1( u1_u4_u1_n129 ) , .B2( u1_u4_u1_n160 ) , .A( u1_u4_u1_n167 ) );
  NAND2_X1 u1_u4_u1_U63 (.A2( u1_u4_u1_n100 ) , .A1( u1_u4_u1_n103 ) , .ZN( u1_u4_u1_n120 ) );
  NAND2_X1 u1_u4_u1_U64 (.A1( u1_u4_u1_n102 ) , .A2( u1_u4_u1_n104 ) , .ZN( u1_u4_u1_n115 ) );
  NAND2_X1 u1_u4_u1_U65 (.A2( u1_u4_u1_n100 ) , .A1( u1_u4_u1_n104 ) , .ZN( u1_u4_u1_n151 ) );
  NAND2_X1 u1_u4_u1_U66 (.A2( u1_u4_u1_n103 ) , .A1( u1_u4_u1_n105 ) , .ZN( u1_u4_u1_n161 ) );
  INV_X1 u1_u4_u1_U67 (.A( u1_u4_u1_n152 ) , .ZN( u1_u4_u1_n173 ) );
  INV_X1 u1_u4_u1_U68 (.A( u1_u4_u1_n128 ) , .ZN( u1_u4_u1_n172 ) );
  NAND2_X1 u1_u4_u1_U69 (.A2( u1_u4_u1_n102 ) , .A1( u1_u4_u1_n103 ) , .ZN( u1_u4_u1_n123 ) );
  NAND2_X1 u1_u4_u1_U7 (.ZN( u1_u4_u1_n114 ) , .A1( u1_u4_u1_n134 ) , .A2( u1_u4_u1_n156 ) );
  NOR2_X1 u1_u4_u1_U70 (.A2( u1_u4_X_7 ) , .A1( u1_u4_X_8 ) , .ZN( u1_u4_u1_n95 ) );
  NOR2_X1 u1_u4_u1_U71 (.A1( u1_u4_X_12 ) , .A2( u1_u4_X_9 ) , .ZN( u1_u4_u1_n100 ) );
  NOR2_X1 u1_u4_u1_U72 (.A2( u1_u4_X_8 ) , .A1( u1_u4_u1_n177 ) , .ZN( u1_u4_u1_n99 ) );
  NOR2_X1 u1_u4_u1_U73 (.A2( u1_u4_X_12 ) , .ZN( u1_u4_u1_n102 ) , .A1( u1_u4_u1_n176 ) );
  NOR2_X1 u1_u4_u1_U74 (.A2( u1_u4_X_9 ) , .ZN( u1_u4_u1_n105 ) , .A1( u1_u4_u1_n168 ) );
  NAND2_X1 u1_u4_u1_U75 (.A1( u1_u4_X_10 ) , .ZN( u1_u4_u1_n160 ) , .A2( u1_u4_u1_n169 ) );
  NAND2_X1 u1_u4_u1_U76 (.A2( u1_u4_X_10 ) , .A1( u1_u4_X_11 ) , .ZN( u1_u4_u1_n152 ) );
  NAND2_X1 u1_u4_u1_U77 (.A1( u1_u4_X_11 ) , .ZN( u1_u4_u1_n128 ) , .A2( u1_u4_u1_n170 ) );
  AND2_X1 u1_u4_u1_U78 (.A2( u1_u4_X_7 ) , .A1( u1_u4_X_8 ) , .ZN( u1_u4_u1_n104 ) );
  AND2_X1 u1_u4_u1_U79 (.A1( u1_u4_X_8 ) , .ZN( u1_u4_u1_n103 ) , .A2( u1_u4_u1_n177 ) );
  AOI22_X1 u1_u4_u1_U8 (.B2( u1_u4_u1_n136 ) , .A2( u1_u4_u1_n137 ) , .ZN( u1_u4_u1_n143 ) , .A1( u1_u4_u1_n171 ) , .B1( u1_u4_u1_n173 ) );
  INV_X1 u1_u4_u1_U80 (.A( u1_u4_X_10 ) , .ZN( u1_u4_u1_n170 ) );
  INV_X1 u1_u4_u1_U81 (.A( u1_u4_X_9 ) , .ZN( u1_u4_u1_n176 ) );
  INV_X1 u1_u4_u1_U82 (.A( u1_u4_X_11 ) , .ZN( u1_u4_u1_n169 ) );
  INV_X1 u1_u4_u1_U83 (.A( u1_u4_X_12 ) , .ZN( u1_u4_u1_n168 ) );
  INV_X1 u1_u4_u1_U84 (.A( u1_u4_X_7 ) , .ZN( u1_u4_u1_n177 ) );
  NAND4_X1 u1_u4_u1_U85 (.ZN( u1_out4_18 ) , .A4( u1_u4_u1_n165 ) , .A3( u1_u4_u1_n166 ) , .A1( u1_u4_u1_n167 ) , .A2( u1_u4_u1_n186 ) );
  AOI22_X1 u1_u4_u1_U86 (.B2( u1_u4_u1_n146 ) , .B1( u1_u4_u1_n147 ) , .A2( u1_u4_u1_n148 ) , .ZN( u1_u4_u1_n166 ) , .A1( u1_u4_u1_n172 ) );
  INV_X1 u1_u4_u1_U87 (.A( u1_u4_u1_n145 ) , .ZN( u1_u4_u1_n186 ) );
  NAND4_X1 u1_u4_u1_U88 (.ZN( u1_out4_2 ) , .A4( u1_u4_u1_n142 ) , .A3( u1_u4_u1_n143 ) , .A2( u1_u4_u1_n144 ) , .A1( u1_u4_u1_n179 ) );
  OAI21_X1 u1_u4_u1_U89 (.B2( u1_u4_u1_n132 ) , .ZN( u1_u4_u1_n144 ) , .A( u1_u4_u1_n146 ) , .B1( u1_u4_u1_n180 ) );
  INV_X1 u1_u4_u1_U9 (.A( u1_u4_u1_n147 ) , .ZN( u1_u4_u1_n181 ) );
  INV_X1 u1_u4_u1_U90 (.A( u1_u4_u1_n130 ) , .ZN( u1_u4_u1_n179 ) );
  NAND4_X1 u1_u4_u1_U91 (.ZN( u1_out4_28 ) , .A4( u1_u4_u1_n124 ) , .A3( u1_u4_u1_n125 ) , .A2( u1_u4_u1_n126 ) , .A1( u1_u4_u1_n127 ) );
  OAI21_X1 u1_u4_u1_U92 (.ZN( u1_u4_u1_n127 ) , .B2( u1_u4_u1_n139 ) , .B1( u1_u4_u1_n175 ) , .A( u1_u4_u1_n183 ) );
  OAI21_X1 u1_u4_u1_U93 (.ZN( u1_u4_u1_n126 ) , .B2( u1_u4_u1_n140 ) , .A( u1_u4_u1_n146 ) , .B1( u1_u4_u1_n178 ) );
  OR4_X1 u1_u4_u1_U94 (.ZN( u1_out4_13 ) , .A4( u1_u4_u1_n108 ) , .A3( u1_u4_u1_n109 ) , .A2( u1_u4_u1_n110 ) , .A1( u1_u4_u1_n111 ) );
  AOI21_X1 u1_u4_u1_U95 (.ZN( u1_u4_u1_n111 ) , .A( u1_u4_u1_n128 ) , .B2( u1_u4_u1_n131 ) , .B1( u1_u4_u1_n135 ) );
  AOI21_X1 u1_u4_u1_U96 (.ZN( u1_u4_u1_n110 ) , .A( u1_u4_u1_n116 ) , .B1( u1_u4_u1_n152 ) , .B2( u1_u4_u1_n160 ) );
  NAND3_X1 u1_u4_u1_U97 (.A3( u1_u4_u1_n149 ) , .A2( u1_u4_u1_n150 ) , .A1( u1_u4_u1_n151 ) , .ZN( u1_u4_u1_n164 ) );
  NAND3_X1 u1_u4_u1_U98 (.A3( u1_u4_u1_n134 ) , .A2( u1_u4_u1_n135 ) , .ZN( u1_u4_u1_n136 ) , .A1( u1_u4_u1_n151 ) );
  NAND3_X1 u1_u4_u1_U99 (.A1( u1_u4_u1_n133 ) , .ZN( u1_u4_u1_n137 ) , .A2( u1_u4_u1_n154 ) , .A3( u1_u4_u1_n181 ) );
  XOR2_X1 u1_u5_U1 (.B( u1_K6_9 ) , .A( u1_R4_6 ) , .Z( u1_u5_X_9 ) );
  XOR2_X1 u1_u5_U10 (.B( u1_K6_45 ) , .A( u1_R4_30 ) , .Z( u1_u5_X_45 ) );
  XOR2_X1 u1_u5_U11 (.B( u1_K6_44 ) , .A( u1_R4_29 ) , .Z( u1_u5_X_44 ) );
  XOR2_X1 u1_u5_U12 (.B( u1_K6_43 ) , .A( u1_R4_28 ) , .Z( u1_u5_X_43 ) );
  XOR2_X1 u1_u5_U13 (.B( u1_K6_42 ) , .A( u1_R4_29 ) , .Z( u1_u5_X_42 ) );
  XOR2_X1 u1_u5_U14 (.B( u1_K6_41 ) , .A( u1_R4_28 ) , .Z( u1_u5_X_41 ) );
  XOR2_X1 u1_u5_U15 (.B( u1_K6_40 ) , .A( u1_R4_27 ) , .Z( u1_u5_X_40 ) );
  XOR2_X1 u1_u5_U16 (.B( u1_K6_3 ) , .A( u1_R4_2 ) , .Z( u1_u5_X_3 ) );
  XOR2_X1 u1_u5_U17 (.B( u1_K6_39 ) , .A( u1_R4_26 ) , .Z( u1_u5_X_39 ) );
  XOR2_X1 u1_u5_U18 (.B( u1_K6_38 ) , .A( u1_R4_25 ) , .Z( u1_u5_X_38 ) );
  XOR2_X1 u1_u5_U19 (.B( u1_K6_37 ) , .A( u1_R4_24 ) , .Z( u1_u5_X_37 ) );
  XOR2_X1 u1_u5_U2 (.B( u1_K6_8 ) , .A( u1_R4_5 ) , .Z( u1_u5_X_8 ) );
  XOR2_X1 u1_u5_U20 (.B( u1_K6_36 ) , .A( u1_R4_25 ) , .Z( u1_u5_X_36 ) );
  XOR2_X1 u1_u5_U21 (.B( u1_K6_35 ) , .A( u1_R4_24 ) , .Z( u1_u5_X_35 ) );
  XOR2_X1 u1_u5_U22 (.B( u1_K6_34 ) , .A( u1_R4_23 ) , .Z( u1_u5_X_34 ) );
  XOR2_X1 u1_u5_U23 (.B( u1_K6_33 ) , .A( u1_R4_22 ) , .Z( u1_u5_X_33 ) );
  XOR2_X1 u1_u5_U27 (.B( u1_K6_2 ) , .A( u1_R4_1 ) , .Z( u1_u5_X_2 ) );
  XOR2_X1 u1_u5_U35 (.B( u1_K6_22 ) , .A( u1_R4_15 ) , .Z( u1_u5_X_22 ) );
  XOR2_X1 u1_u5_U36 (.B( u1_K6_21 ) , .A( u1_R4_14 ) , .Z( u1_u5_X_21 ) );
  XOR2_X1 u1_u5_U38 (.B( u1_K6_1 ) , .A( u1_R4_32 ) , .Z( u1_u5_X_1 ) );
  XOR2_X1 u1_u5_U4 (.B( u1_K6_6 ) , .A( u1_R4_5 ) , .Z( u1_u5_X_6 ) );
  XOR2_X1 u1_u5_U48 (.B( u1_K6_10 ) , .A( u1_R4_7 ) , .Z( u1_u5_X_10 ) );
  XOR2_X1 u1_u5_U6 (.B( u1_K6_4 ) , .A( u1_R4_3 ) , .Z( u1_u5_X_4 ) );
  XOR2_X1 u1_u5_U7 (.B( u1_K6_48 ) , .A( u1_R4_1 ) , .Z( u1_u5_X_48 ) );
  XOR2_X1 u1_u5_U8 (.B( u1_K6_47 ) , .A( u1_R4_32 ) , .Z( u1_u5_X_47 ) );
  XOR2_X1 u1_u5_U9 (.B( u1_K6_46 ) , .A( u1_R4_31 ) , .Z( u1_u5_X_46 ) );
  NAND2_X1 u1_u5_u0_U10 (.ZN( u1_u5_u0_n113 ) , .A1( u1_u5_u0_n139 ) , .A2( u1_u5_u0_n149 ) );
  AND3_X1 u1_u5_u0_U11 (.A2( u1_u5_u0_n112 ) , .ZN( u1_u5_u0_n127 ) , .A3( u1_u5_u0_n130 ) , .A1( u1_u5_u0_n148 ) );
  AND2_X1 u1_u5_u0_U12 (.ZN( u1_u5_u0_n107 ) , .A1( u1_u5_u0_n130 ) , .A2( u1_u5_u0_n140 ) );
  AND2_X1 u1_u5_u0_U13 (.A2( u1_u5_u0_n129 ) , .A1( u1_u5_u0_n130 ) , .ZN( u1_u5_u0_n151 ) );
  AND2_X1 u1_u5_u0_U14 (.A1( u1_u5_u0_n108 ) , .A2( u1_u5_u0_n125 ) , .ZN( u1_u5_u0_n145 ) );
  INV_X1 u1_u5_u0_U15 (.A( u1_u5_u0_n143 ) , .ZN( u1_u5_u0_n173 ) );
  NOR2_X1 u1_u5_u0_U16 (.A2( u1_u5_u0_n136 ) , .ZN( u1_u5_u0_n147 ) , .A1( u1_u5_u0_n160 ) );
  AOI21_X1 u1_u5_u0_U17 (.B1( u1_u5_u0_n103 ) , .ZN( u1_u5_u0_n132 ) , .A( u1_u5_u0_n165 ) , .B2( u1_u5_u0_n93 ) );
  INV_X1 u1_u5_u0_U18 (.A( u1_u5_u0_n142 ) , .ZN( u1_u5_u0_n165 ) );
  OAI22_X1 u1_u5_u0_U19 (.B1( u1_u5_u0_n131 ) , .A1( u1_u5_u0_n144 ) , .B2( u1_u5_u0_n147 ) , .A2( u1_u5_u0_n90 ) , .ZN( u1_u5_u0_n91 ) );
  AND3_X1 u1_u5_u0_U20 (.A3( u1_u5_u0_n121 ) , .A2( u1_u5_u0_n125 ) , .A1( u1_u5_u0_n148 ) , .ZN( u1_u5_u0_n90 ) );
  OAI22_X1 u1_u5_u0_U21 (.B1( u1_u5_u0_n125 ) , .ZN( u1_u5_u0_n126 ) , .A1( u1_u5_u0_n138 ) , .A2( u1_u5_u0_n146 ) , .B2( u1_u5_u0_n147 ) );
  NOR2_X1 u1_u5_u0_U22 (.A1( u1_u5_u0_n163 ) , .A2( u1_u5_u0_n164 ) , .ZN( u1_u5_u0_n95 ) );
  INV_X1 u1_u5_u0_U23 (.A( u1_u5_u0_n136 ) , .ZN( u1_u5_u0_n161 ) );
  AOI22_X1 u1_u5_u0_U24 (.B2( u1_u5_u0_n109 ) , .A2( u1_u5_u0_n110 ) , .ZN( u1_u5_u0_n111 ) , .B1( u1_u5_u0_n118 ) , .A1( u1_u5_u0_n160 ) );
  NAND2_X1 u1_u5_u0_U25 (.A2( u1_u5_u0_n102 ) , .A1( u1_u5_u0_n103 ) , .ZN( u1_u5_u0_n149 ) );
  INV_X1 u1_u5_u0_U26 (.A( u1_u5_u0_n118 ) , .ZN( u1_u5_u0_n158 ) );
  NAND2_X1 u1_u5_u0_U27 (.A2( u1_u5_u0_n100 ) , .ZN( u1_u5_u0_n131 ) , .A1( u1_u5_u0_n92 ) );
  NAND2_X1 u1_u5_u0_U28 (.ZN( u1_u5_u0_n108 ) , .A1( u1_u5_u0_n92 ) , .A2( u1_u5_u0_n94 ) );
  AOI21_X1 u1_u5_u0_U29 (.ZN( u1_u5_u0_n104 ) , .B1( u1_u5_u0_n107 ) , .B2( u1_u5_u0_n141 ) , .A( u1_u5_u0_n144 ) );
  INV_X1 u1_u5_u0_U3 (.A( u1_u5_u0_n113 ) , .ZN( u1_u5_u0_n166 ) );
  AOI21_X1 u1_u5_u0_U30 (.B1( u1_u5_u0_n127 ) , .B2( u1_u5_u0_n129 ) , .A( u1_u5_u0_n138 ) , .ZN( u1_u5_u0_n96 ) );
  NAND2_X1 u1_u5_u0_U31 (.A2( u1_u5_u0_n102 ) , .ZN( u1_u5_u0_n114 ) , .A1( u1_u5_u0_n92 ) );
  AOI21_X1 u1_u5_u0_U32 (.ZN( u1_u5_u0_n116 ) , .B2( u1_u5_u0_n142 ) , .A( u1_u5_u0_n144 ) , .B1( u1_u5_u0_n166 ) );
  NOR2_X1 u1_u5_u0_U33 (.A1( u1_u5_u0_n120 ) , .ZN( u1_u5_u0_n143 ) , .A2( u1_u5_u0_n167 ) );
  OAI221_X1 u1_u5_u0_U34 (.C1( u1_u5_u0_n112 ) , .ZN( u1_u5_u0_n120 ) , .B1( u1_u5_u0_n138 ) , .B2( u1_u5_u0_n141 ) , .C2( u1_u5_u0_n147 ) , .A( u1_u5_u0_n172 ) );
  AOI211_X1 u1_u5_u0_U35 (.B( u1_u5_u0_n115 ) , .A( u1_u5_u0_n116 ) , .C2( u1_u5_u0_n117 ) , .C1( u1_u5_u0_n118 ) , .ZN( u1_u5_u0_n119 ) );
  NAND2_X1 u1_u5_u0_U36 (.A2( u1_u5_u0_n103 ) , .ZN( u1_u5_u0_n140 ) , .A1( u1_u5_u0_n94 ) );
  NAND2_X1 u1_u5_u0_U37 (.A1( u1_u5_u0_n100 ) , .A2( u1_u5_u0_n103 ) , .ZN( u1_u5_u0_n125 ) );
  NAND2_X1 u1_u5_u0_U38 (.A1( u1_u5_u0_n101 ) , .A2( u1_u5_u0_n102 ) , .ZN( u1_u5_u0_n150 ) );
  INV_X1 u1_u5_u0_U39 (.A( u1_u5_u0_n138 ) , .ZN( u1_u5_u0_n160 ) );
  AOI21_X1 u1_u5_u0_U4 (.B1( u1_u5_u0_n114 ) , .ZN( u1_u5_u0_n115 ) , .B2( u1_u5_u0_n129 ) , .A( u1_u5_u0_n161 ) );
  NAND2_X1 u1_u5_u0_U40 (.A2( u1_u5_u0_n100 ) , .A1( u1_u5_u0_n101 ) , .ZN( u1_u5_u0_n139 ) );
  NAND2_X1 u1_u5_u0_U41 (.ZN( u1_u5_u0_n112 ) , .A2( u1_u5_u0_n92 ) , .A1( u1_u5_u0_n93 ) );
  NAND2_X1 u1_u5_u0_U42 (.A1( u1_u5_u0_n101 ) , .ZN( u1_u5_u0_n130 ) , .A2( u1_u5_u0_n94 ) );
  INV_X1 u1_u5_u0_U43 (.ZN( u1_u5_u0_n172 ) , .A( u1_u5_u0_n88 ) );
  OAI222_X1 u1_u5_u0_U44 (.C1( u1_u5_u0_n108 ) , .A1( u1_u5_u0_n125 ) , .B2( u1_u5_u0_n128 ) , .B1( u1_u5_u0_n144 ) , .A2( u1_u5_u0_n158 ) , .C2( u1_u5_u0_n161 ) , .ZN( u1_u5_u0_n88 ) );
  NAND2_X1 u1_u5_u0_U45 (.A2( u1_u5_u0_n101 ) , .ZN( u1_u5_u0_n121 ) , .A1( u1_u5_u0_n93 ) );
  OR3_X1 u1_u5_u0_U46 (.A3( u1_u5_u0_n152 ) , .A2( u1_u5_u0_n153 ) , .A1( u1_u5_u0_n154 ) , .ZN( u1_u5_u0_n155 ) );
  AOI21_X1 u1_u5_u0_U47 (.A( u1_u5_u0_n144 ) , .B2( u1_u5_u0_n145 ) , .B1( u1_u5_u0_n146 ) , .ZN( u1_u5_u0_n154 ) );
  AOI21_X1 u1_u5_u0_U48 (.B2( u1_u5_u0_n150 ) , .B1( u1_u5_u0_n151 ) , .ZN( u1_u5_u0_n152 ) , .A( u1_u5_u0_n158 ) );
  AOI21_X1 u1_u5_u0_U49 (.A( u1_u5_u0_n147 ) , .B2( u1_u5_u0_n148 ) , .B1( u1_u5_u0_n149 ) , .ZN( u1_u5_u0_n153 ) );
  AOI21_X1 u1_u5_u0_U5 (.B2( u1_u5_u0_n131 ) , .ZN( u1_u5_u0_n134 ) , .B1( u1_u5_u0_n151 ) , .A( u1_u5_u0_n158 ) );
  INV_X1 u1_u5_u0_U50 (.ZN( u1_u5_u0_n171 ) , .A( u1_u5_u0_n99 ) );
  OAI211_X1 u1_u5_u0_U51 (.C2( u1_u5_u0_n140 ) , .C1( u1_u5_u0_n161 ) , .A( u1_u5_u0_n169 ) , .B( u1_u5_u0_n98 ) , .ZN( u1_u5_u0_n99 ) );
  INV_X1 u1_u5_u0_U52 (.ZN( u1_u5_u0_n169 ) , .A( u1_u5_u0_n91 ) );
  AOI211_X1 u1_u5_u0_U53 (.C1( u1_u5_u0_n118 ) , .A( u1_u5_u0_n123 ) , .B( u1_u5_u0_n96 ) , .C2( u1_u5_u0_n97 ) , .ZN( u1_u5_u0_n98 ) );
  NOR2_X1 u1_u5_u0_U54 (.A2( u1_u5_X_4 ) , .A1( u1_u5_X_5 ) , .ZN( u1_u5_u0_n118 ) );
  NOR2_X1 u1_u5_u0_U55 (.A2( u1_u5_X_1 ) , .ZN( u1_u5_u0_n101 ) , .A1( u1_u5_u0_n163 ) );
  NOR2_X1 u1_u5_u0_U56 (.A2( u1_u5_X_3 ) , .A1( u1_u5_X_6 ) , .ZN( u1_u5_u0_n94 ) );
  NOR2_X1 u1_u5_u0_U57 (.A2( u1_u5_X_6 ) , .ZN( u1_u5_u0_n100 ) , .A1( u1_u5_u0_n162 ) );
  NAND2_X1 u1_u5_u0_U58 (.A2( u1_u5_X_4 ) , .A1( u1_u5_X_5 ) , .ZN( u1_u5_u0_n144 ) );
  NOR2_X1 u1_u5_u0_U59 (.A2( u1_u5_X_5 ) , .ZN( u1_u5_u0_n136 ) , .A1( u1_u5_u0_n159 ) );
  NOR2_X1 u1_u5_u0_U6 (.A1( u1_u5_u0_n108 ) , .ZN( u1_u5_u0_n123 ) , .A2( u1_u5_u0_n158 ) );
  NAND2_X1 u1_u5_u0_U60 (.A1( u1_u5_X_5 ) , .ZN( u1_u5_u0_n138 ) , .A2( u1_u5_u0_n159 ) );
  AND2_X1 u1_u5_u0_U61 (.A2( u1_u5_X_3 ) , .A1( u1_u5_X_6 ) , .ZN( u1_u5_u0_n102 ) );
  AND2_X1 u1_u5_u0_U62 (.A1( u1_u5_X_6 ) , .A2( u1_u5_u0_n162 ) , .ZN( u1_u5_u0_n93 ) );
  INV_X1 u1_u5_u0_U63 (.A( u1_u5_X_4 ) , .ZN( u1_u5_u0_n159 ) );
  INV_X1 u1_u5_u0_U64 (.A( u1_u5_X_1 ) , .ZN( u1_u5_u0_n164 ) );
  INV_X1 u1_u5_u0_U65 (.A( u1_u5_X_3 ) , .ZN( u1_u5_u0_n162 ) );
  INV_X1 u1_u5_u0_U66 (.A( u1_u5_u0_n126 ) , .ZN( u1_u5_u0_n168 ) );
  AOI211_X1 u1_u5_u0_U67 (.B( u1_u5_u0_n133 ) , .A( u1_u5_u0_n134 ) , .C2( u1_u5_u0_n135 ) , .C1( u1_u5_u0_n136 ) , .ZN( u1_u5_u0_n137 ) );
  OR4_X1 u1_u5_u0_U68 (.ZN( u1_out5_17 ) , .A1( u1_u5_u0_n122 ) , .A2( u1_u5_u0_n123 ) , .A4( u1_u5_u0_n124 ) , .A3( u1_u5_u0_n170 ) );
  AOI21_X1 u1_u5_u0_U69 (.B2( u1_u5_u0_n107 ) , .ZN( u1_u5_u0_n124 ) , .B1( u1_u5_u0_n128 ) , .A( u1_u5_u0_n161 ) );
  OAI21_X1 u1_u5_u0_U7 (.B1( u1_u5_u0_n150 ) , .B2( u1_u5_u0_n158 ) , .A( u1_u5_u0_n172 ) , .ZN( u1_u5_u0_n89 ) );
  INV_X1 u1_u5_u0_U70 (.A( u1_u5_u0_n111 ) , .ZN( u1_u5_u0_n170 ) );
  OR4_X1 u1_u5_u0_U71 (.ZN( u1_out5_31 ) , .A4( u1_u5_u0_n155 ) , .A2( u1_u5_u0_n156 ) , .A1( u1_u5_u0_n157 ) , .A3( u1_u5_u0_n173 ) );
  AOI21_X1 u1_u5_u0_U72 (.A( u1_u5_u0_n138 ) , .B2( u1_u5_u0_n139 ) , .B1( u1_u5_u0_n140 ) , .ZN( u1_u5_u0_n157 ) );
  AOI21_X1 u1_u5_u0_U73 (.B2( u1_u5_u0_n141 ) , .B1( u1_u5_u0_n142 ) , .ZN( u1_u5_u0_n156 ) , .A( u1_u5_u0_n161 ) );
  INV_X1 u1_u5_u0_U74 (.ZN( u1_u5_u0_n174 ) , .A( u1_u5_u0_n89 ) );
  AOI211_X1 u1_u5_u0_U75 (.B( u1_u5_u0_n104 ) , .A( u1_u5_u0_n105 ) , .ZN( u1_u5_u0_n106 ) , .C2( u1_u5_u0_n113 ) , .C1( u1_u5_u0_n160 ) );
  OAI221_X1 u1_u5_u0_U76 (.C1( u1_u5_u0_n121 ) , .ZN( u1_u5_u0_n122 ) , .B2( u1_u5_u0_n127 ) , .A( u1_u5_u0_n143 ) , .B1( u1_u5_u0_n144 ) , .C2( u1_u5_u0_n147 ) );
  AOI21_X1 u1_u5_u0_U77 (.B1( u1_u5_u0_n132 ) , .ZN( u1_u5_u0_n133 ) , .A( u1_u5_u0_n144 ) , .B2( u1_u5_u0_n166 ) );
  OAI22_X1 u1_u5_u0_U78 (.ZN( u1_u5_u0_n105 ) , .A2( u1_u5_u0_n132 ) , .B1( u1_u5_u0_n146 ) , .A1( u1_u5_u0_n147 ) , .B2( u1_u5_u0_n161 ) );
  NAND2_X1 u1_u5_u0_U79 (.ZN( u1_u5_u0_n110 ) , .A2( u1_u5_u0_n132 ) , .A1( u1_u5_u0_n145 ) );
  AND2_X1 u1_u5_u0_U8 (.A1( u1_u5_u0_n114 ) , .A2( u1_u5_u0_n121 ) , .ZN( u1_u5_u0_n146 ) );
  INV_X1 u1_u5_u0_U80 (.A( u1_u5_u0_n119 ) , .ZN( u1_u5_u0_n167 ) );
  NAND2_X1 u1_u5_u0_U81 (.ZN( u1_u5_u0_n148 ) , .A1( u1_u5_u0_n93 ) , .A2( u1_u5_u0_n95 ) );
  NAND2_X1 u1_u5_u0_U82 (.A1( u1_u5_u0_n100 ) , .ZN( u1_u5_u0_n129 ) , .A2( u1_u5_u0_n95 ) );
  NAND2_X1 u1_u5_u0_U83 (.A1( u1_u5_u0_n102 ) , .ZN( u1_u5_u0_n128 ) , .A2( u1_u5_u0_n95 ) );
  NOR2_X1 u1_u5_u0_U84 (.A2( u1_u5_X_1 ) , .A1( u1_u5_X_2 ) , .ZN( u1_u5_u0_n92 ) );
  NAND2_X1 u1_u5_u0_U85 (.ZN( u1_u5_u0_n142 ) , .A1( u1_u5_u0_n94 ) , .A2( u1_u5_u0_n95 ) );
  NOR2_X1 u1_u5_u0_U86 (.A2( u1_u5_X_2 ) , .ZN( u1_u5_u0_n103 ) , .A1( u1_u5_u0_n164 ) );
  INV_X1 u1_u5_u0_U87 (.A( u1_u5_X_2 ) , .ZN( u1_u5_u0_n163 ) );
  NAND3_X1 u1_u5_u0_U88 (.ZN( u1_out5_23 ) , .A3( u1_u5_u0_n137 ) , .A1( u1_u5_u0_n168 ) , .A2( u1_u5_u0_n171 ) );
  NAND3_X1 u1_u5_u0_U89 (.A3( u1_u5_u0_n127 ) , .A2( u1_u5_u0_n128 ) , .ZN( u1_u5_u0_n135 ) , .A1( u1_u5_u0_n150 ) );
  AND2_X1 u1_u5_u0_U9 (.A1( u1_u5_u0_n131 ) , .ZN( u1_u5_u0_n141 ) , .A2( u1_u5_u0_n150 ) );
  NAND3_X1 u1_u5_u0_U90 (.ZN( u1_u5_u0_n117 ) , .A3( u1_u5_u0_n132 ) , .A2( u1_u5_u0_n139 ) , .A1( u1_u5_u0_n148 ) );
  NAND3_X1 u1_u5_u0_U91 (.ZN( u1_u5_u0_n109 ) , .A2( u1_u5_u0_n114 ) , .A3( u1_u5_u0_n140 ) , .A1( u1_u5_u0_n149 ) );
  NAND3_X1 u1_u5_u0_U92 (.ZN( u1_out5_9 ) , .A3( u1_u5_u0_n106 ) , .A2( u1_u5_u0_n171 ) , .A1( u1_u5_u0_n174 ) );
  NAND3_X1 u1_u5_u0_U93 (.A2( u1_u5_u0_n128 ) , .A1( u1_u5_u0_n132 ) , .A3( u1_u5_u0_n146 ) , .ZN( u1_u5_u0_n97 ) );
  AOI21_X1 u1_u5_u1_U10 (.B2( u1_u5_u1_n155 ) , .B1( u1_u5_u1_n156 ) , .ZN( u1_u5_u1_n157 ) , .A( u1_u5_u1_n174 ) );
  NAND3_X1 u1_u5_u1_U100 (.ZN( u1_u5_u1_n113 ) , .A1( u1_u5_u1_n120 ) , .A3( u1_u5_u1_n133 ) , .A2( u1_u5_u1_n155 ) );
  NAND2_X1 u1_u5_u1_U11 (.ZN( u1_u5_u1_n140 ) , .A2( u1_u5_u1_n150 ) , .A1( u1_u5_u1_n155 ) );
  NAND2_X1 u1_u5_u1_U12 (.A1( u1_u5_u1_n131 ) , .ZN( u1_u5_u1_n147 ) , .A2( u1_u5_u1_n153 ) );
  INV_X1 u1_u5_u1_U13 (.A( u1_u5_u1_n139 ) , .ZN( u1_u5_u1_n174 ) );
  OR4_X1 u1_u5_u1_U14 (.A4( u1_u5_u1_n106 ) , .A3( u1_u5_u1_n107 ) , .ZN( u1_u5_u1_n108 ) , .A1( u1_u5_u1_n117 ) , .A2( u1_u5_u1_n184 ) );
  AOI21_X1 u1_u5_u1_U15 (.ZN( u1_u5_u1_n106 ) , .A( u1_u5_u1_n112 ) , .B1( u1_u5_u1_n154 ) , .B2( u1_u5_u1_n156 ) );
  INV_X1 u1_u5_u1_U16 (.A( u1_u5_u1_n101 ) , .ZN( u1_u5_u1_n184 ) );
  AOI21_X1 u1_u5_u1_U17 (.ZN( u1_u5_u1_n107 ) , .B1( u1_u5_u1_n134 ) , .B2( u1_u5_u1_n149 ) , .A( u1_u5_u1_n174 ) );
  INV_X1 u1_u5_u1_U18 (.A( u1_u5_u1_n112 ) , .ZN( u1_u5_u1_n171 ) );
  NAND2_X1 u1_u5_u1_U19 (.ZN( u1_u5_u1_n141 ) , .A1( u1_u5_u1_n153 ) , .A2( u1_u5_u1_n156 ) );
  AND2_X1 u1_u5_u1_U20 (.A1( u1_u5_u1_n123 ) , .ZN( u1_u5_u1_n134 ) , .A2( u1_u5_u1_n161 ) );
  NAND2_X1 u1_u5_u1_U21 (.A2( u1_u5_u1_n115 ) , .A1( u1_u5_u1_n116 ) , .ZN( u1_u5_u1_n148 ) );
  NAND2_X1 u1_u5_u1_U22 (.A2( u1_u5_u1_n133 ) , .A1( u1_u5_u1_n135 ) , .ZN( u1_u5_u1_n159 ) );
  NAND2_X1 u1_u5_u1_U23 (.A2( u1_u5_u1_n115 ) , .A1( u1_u5_u1_n120 ) , .ZN( u1_u5_u1_n132 ) );
  INV_X1 u1_u5_u1_U24 (.A( u1_u5_u1_n154 ) , .ZN( u1_u5_u1_n178 ) );
  AOI22_X1 u1_u5_u1_U25 (.B2( u1_u5_u1_n113 ) , .A2( u1_u5_u1_n114 ) , .ZN( u1_u5_u1_n125 ) , .A1( u1_u5_u1_n171 ) , .B1( u1_u5_u1_n173 ) );
  NAND2_X1 u1_u5_u1_U26 (.ZN( u1_u5_u1_n114 ) , .A1( u1_u5_u1_n134 ) , .A2( u1_u5_u1_n156 ) );
  INV_X1 u1_u5_u1_U27 (.A( u1_u5_u1_n151 ) , .ZN( u1_u5_u1_n183 ) );
  AND2_X1 u1_u5_u1_U28 (.A1( u1_u5_u1_n129 ) , .A2( u1_u5_u1_n133 ) , .ZN( u1_u5_u1_n149 ) );
  INV_X1 u1_u5_u1_U29 (.A( u1_u5_u1_n131 ) , .ZN( u1_u5_u1_n180 ) );
  INV_X1 u1_u5_u1_U3 (.A( u1_u5_u1_n159 ) , .ZN( u1_u5_u1_n182 ) );
  OAI221_X1 u1_u5_u1_U30 (.A( u1_u5_u1_n119 ) , .C2( u1_u5_u1_n129 ) , .ZN( u1_u5_u1_n138 ) , .B2( u1_u5_u1_n152 ) , .C1( u1_u5_u1_n174 ) , .B1( u1_u5_u1_n187 ) );
  INV_X1 u1_u5_u1_U31 (.A( u1_u5_u1_n148 ) , .ZN( u1_u5_u1_n187 ) );
  AOI211_X1 u1_u5_u1_U32 (.B( u1_u5_u1_n117 ) , .A( u1_u5_u1_n118 ) , .ZN( u1_u5_u1_n119 ) , .C2( u1_u5_u1_n146 ) , .C1( u1_u5_u1_n159 ) );
  NOR2_X1 u1_u5_u1_U33 (.A1( u1_u5_u1_n168 ) , .A2( u1_u5_u1_n176 ) , .ZN( u1_u5_u1_n98 ) );
  AOI211_X1 u1_u5_u1_U34 (.B( u1_u5_u1_n162 ) , .A( u1_u5_u1_n163 ) , .C2( u1_u5_u1_n164 ) , .ZN( u1_u5_u1_n165 ) , .C1( u1_u5_u1_n171 ) );
  AOI21_X1 u1_u5_u1_U35 (.A( u1_u5_u1_n160 ) , .B2( u1_u5_u1_n161 ) , .ZN( u1_u5_u1_n162 ) , .B1( u1_u5_u1_n182 ) );
  OR2_X1 u1_u5_u1_U36 (.A2( u1_u5_u1_n157 ) , .A1( u1_u5_u1_n158 ) , .ZN( u1_u5_u1_n163 ) );
  OAI21_X1 u1_u5_u1_U37 (.B2( u1_u5_u1_n123 ) , .ZN( u1_u5_u1_n145 ) , .B1( u1_u5_u1_n160 ) , .A( u1_u5_u1_n185 ) );
  INV_X1 u1_u5_u1_U38 (.A( u1_u5_u1_n122 ) , .ZN( u1_u5_u1_n185 ) );
  AOI21_X1 u1_u5_u1_U39 (.B2( u1_u5_u1_n120 ) , .B1( u1_u5_u1_n121 ) , .ZN( u1_u5_u1_n122 ) , .A( u1_u5_u1_n128 ) );
  AOI221_X1 u1_u5_u1_U4 (.A( u1_u5_u1_n138 ) , .C2( u1_u5_u1_n139 ) , .C1( u1_u5_u1_n140 ) , .B2( u1_u5_u1_n141 ) , .ZN( u1_u5_u1_n142 ) , .B1( u1_u5_u1_n175 ) );
  NAND2_X1 u1_u5_u1_U40 (.A1( u1_u5_u1_n128 ) , .ZN( u1_u5_u1_n146 ) , .A2( u1_u5_u1_n160 ) );
  NAND2_X1 u1_u5_u1_U41 (.A2( u1_u5_u1_n112 ) , .ZN( u1_u5_u1_n139 ) , .A1( u1_u5_u1_n152 ) );
  NAND2_X1 u1_u5_u1_U42 (.A1( u1_u5_u1_n105 ) , .ZN( u1_u5_u1_n156 ) , .A2( u1_u5_u1_n99 ) );
  AOI221_X1 u1_u5_u1_U43 (.B1( u1_u5_u1_n140 ) , .ZN( u1_u5_u1_n167 ) , .B2( u1_u5_u1_n172 ) , .C2( u1_u5_u1_n175 ) , .C1( u1_u5_u1_n178 ) , .A( u1_u5_u1_n188 ) );
  INV_X1 u1_u5_u1_U44 (.ZN( u1_u5_u1_n188 ) , .A( u1_u5_u1_n97 ) );
  AOI211_X1 u1_u5_u1_U45 (.A( u1_u5_u1_n118 ) , .C1( u1_u5_u1_n132 ) , .C2( u1_u5_u1_n139 ) , .B( u1_u5_u1_n96 ) , .ZN( u1_u5_u1_n97 ) );
  AOI21_X1 u1_u5_u1_U46 (.B2( u1_u5_u1_n121 ) , .B1( u1_u5_u1_n135 ) , .A( u1_u5_u1_n152 ) , .ZN( u1_u5_u1_n96 ) );
  NOR2_X1 u1_u5_u1_U47 (.ZN( u1_u5_u1_n117 ) , .A1( u1_u5_u1_n121 ) , .A2( u1_u5_u1_n160 ) );
  AOI21_X1 u1_u5_u1_U48 (.A( u1_u5_u1_n128 ) , .B2( u1_u5_u1_n129 ) , .ZN( u1_u5_u1_n130 ) , .B1( u1_u5_u1_n150 ) );
  NAND2_X1 u1_u5_u1_U49 (.ZN( u1_u5_u1_n112 ) , .A1( u1_u5_u1_n169 ) , .A2( u1_u5_u1_n170 ) );
  AOI211_X1 u1_u5_u1_U5 (.ZN( u1_u5_u1_n124 ) , .A( u1_u5_u1_n138 ) , .C2( u1_u5_u1_n139 ) , .B( u1_u5_u1_n145 ) , .C1( u1_u5_u1_n147 ) );
  NAND2_X1 u1_u5_u1_U50 (.ZN( u1_u5_u1_n129 ) , .A2( u1_u5_u1_n95 ) , .A1( u1_u5_u1_n98 ) );
  NAND2_X1 u1_u5_u1_U51 (.A1( u1_u5_u1_n102 ) , .ZN( u1_u5_u1_n154 ) , .A2( u1_u5_u1_n99 ) );
  NAND2_X1 u1_u5_u1_U52 (.A2( u1_u5_u1_n100 ) , .ZN( u1_u5_u1_n135 ) , .A1( u1_u5_u1_n99 ) );
  AOI21_X1 u1_u5_u1_U53 (.A( u1_u5_u1_n152 ) , .B2( u1_u5_u1_n153 ) , .B1( u1_u5_u1_n154 ) , .ZN( u1_u5_u1_n158 ) );
  INV_X1 u1_u5_u1_U54 (.A( u1_u5_u1_n160 ) , .ZN( u1_u5_u1_n175 ) );
  NAND2_X1 u1_u5_u1_U55 (.A1( u1_u5_u1_n100 ) , .ZN( u1_u5_u1_n116 ) , .A2( u1_u5_u1_n95 ) );
  NAND2_X1 u1_u5_u1_U56 (.A1( u1_u5_u1_n102 ) , .ZN( u1_u5_u1_n131 ) , .A2( u1_u5_u1_n95 ) );
  NAND2_X1 u1_u5_u1_U57 (.A2( u1_u5_u1_n104 ) , .ZN( u1_u5_u1_n121 ) , .A1( u1_u5_u1_n98 ) );
  NAND2_X1 u1_u5_u1_U58 (.A1( u1_u5_u1_n103 ) , .ZN( u1_u5_u1_n153 ) , .A2( u1_u5_u1_n98 ) );
  NAND2_X1 u1_u5_u1_U59 (.A2( u1_u5_u1_n104 ) , .A1( u1_u5_u1_n105 ) , .ZN( u1_u5_u1_n133 ) );
  AOI22_X1 u1_u5_u1_U6 (.B2( u1_u5_u1_n136 ) , .A2( u1_u5_u1_n137 ) , .ZN( u1_u5_u1_n143 ) , .A1( u1_u5_u1_n171 ) , .B1( u1_u5_u1_n173 ) );
  NAND2_X1 u1_u5_u1_U60 (.ZN( u1_u5_u1_n150 ) , .A2( u1_u5_u1_n98 ) , .A1( u1_u5_u1_n99 ) );
  NAND2_X1 u1_u5_u1_U61 (.A1( u1_u5_u1_n105 ) , .ZN( u1_u5_u1_n155 ) , .A2( u1_u5_u1_n95 ) );
  OAI21_X1 u1_u5_u1_U62 (.ZN( u1_u5_u1_n109 ) , .B1( u1_u5_u1_n129 ) , .B2( u1_u5_u1_n160 ) , .A( u1_u5_u1_n167 ) );
  NAND2_X1 u1_u5_u1_U63 (.A2( u1_u5_u1_n100 ) , .A1( u1_u5_u1_n103 ) , .ZN( u1_u5_u1_n120 ) );
  NAND2_X1 u1_u5_u1_U64 (.A1( u1_u5_u1_n102 ) , .A2( u1_u5_u1_n104 ) , .ZN( u1_u5_u1_n115 ) );
  NAND2_X1 u1_u5_u1_U65 (.A2( u1_u5_u1_n100 ) , .A1( u1_u5_u1_n104 ) , .ZN( u1_u5_u1_n151 ) );
  NAND2_X1 u1_u5_u1_U66 (.A2( u1_u5_u1_n103 ) , .A1( u1_u5_u1_n105 ) , .ZN( u1_u5_u1_n161 ) );
  INV_X1 u1_u5_u1_U67 (.A( u1_u5_u1_n152 ) , .ZN( u1_u5_u1_n173 ) );
  INV_X1 u1_u5_u1_U68 (.A( u1_u5_u1_n128 ) , .ZN( u1_u5_u1_n172 ) );
  NAND2_X1 u1_u5_u1_U69 (.A2( u1_u5_u1_n102 ) , .A1( u1_u5_u1_n103 ) , .ZN( u1_u5_u1_n123 ) );
  INV_X1 u1_u5_u1_U7 (.A( u1_u5_u1_n147 ) , .ZN( u1_u5_u1_n181 ) );
  NOR2_X1 u1_u5_u1_U70 (.A2( u1_u5_X_7 ) , .A1( u1_u5_X_8 ) , .ZN( u1_u5_u1_n95 ) );
  NOR2_X1 u1_u5_u1_U71 (.A1( u1_u5_X_12 ) , .A2( u1_u5_X_9 ) , .ZN( u1_u5_u1_n100 ) );
  NOR2_X1 u1_u5_u1_U72 (.A2( u1_u5_X_8 ) , .A1( u1_u5_u1_n177 ) , .ZN( u1_u5_u1_n99 ) );
  NOR2_X1 u1_u5_u1_U73 (.A2( u1_u5_X_12 ) , .ZN( u1_u5_u1_n102 ) , .A1( u1_u5_u1_n176 ) );
  NOR2_X1 u1_u5_u1_U74 (.A2( u1_u5_X_9 ) , .ZN( u1_u5_u1_n105 ) , .A1( u1_u5_u1_n168 ) );
  NAND2_X1 u1_u5_u1_U75 (.A1( u1_u5_X_10 ) , .ZN( u1_u5_u1_n160 ) , .A2( u1_u5_u1_n169 ) );
  NAND2_X1 u1_u5_u1_U76 (.A2( u1_u5_X_10 ) , .A1( u1_u5_X_11 ) , .ZN( u1_u5_u1_n152 ) );
  NAND2_X1 u1_u5_u1_U77 (.A1( u1_u5_X_11 ) , .ZN( u1_u5_u1_n128 ) , .A2( u1_u5_u1_n170 ) );
  AND2_X1 u1_u5_u1_U78 (.A2( u1_u5_X_7 ) , .A1( u1_u5_X_8 ) , .ZN( u1_u5_u1_n104 ) );
  AND2_X1 u1_u5_u1_U79 (.A1( u1_u5_X_8 ) , .ZN( u1_u5_u1_n103 ) , .A2( u1_u5_u1_n177 ) );
  NOR2_X1 u1_u5_u1_U8 (.A1( u1_u5_u1_n112 ) , .A2( u1_u5_u1_n116 ) , .ZN( u1_u5_u1_n118 ) );
  INV_X1 u1_u5_u1_U80 (.A( u1_u5_X_10 ) , .ZN( u1_u5_u1_n170 ) );
  INV_X1 u1_u5_u1_U81 (.A( u1_u5_X_9 ) , .ZN( u1_u5_u1_n176 ) );
  INV_X1 u1_u5_u1_U82 (.A( u1_u5_X_11 ) , .ZN( u1_u5_u1_n169 ) );
  INV_X1 u1_u5_u1_U83 (.A( u1_u5_X_12 ) , .ZN( u1_u5_u1_n168 ) );
  INV_X1 u1_u5_u1_U84 (.A( u1_u5_X_7 ) , .ZN( u1_u5_u1_n177 ) );
  NAND4_X1 u1_u5_u1_U85 (.ZN( u1_out5_18 ) , .A4( u1_u5_u1_n165 ) , .A3( u1_u5_u1_n166 ) , .A1( u1_u5_u1_n167 ) , .A2( u1_u5_u1_n186 ) );
  AOI22_X1 u1_u5_u1_U86 (.B2( u1_u5_u1_n146 ) , .B1( u1_u5_u1_n147 ) , .A2( u1_u5_u1_n148 ) , .ZN( u1_u5_u1_n166 ) , .A1( u1_u5_u1_n172 ) );
  INV_X1 u1_u5_u1_U87 (.A( u1_u5_u1_n145 ) , .ZN( u1_u5_u1_n186 ) );
  OR4_X1 u1_u5_u1_U88 (.ZN( u1_out5_13 ) , .A4( u1_u5_u1_n108 ) , .A3( u1_u5_u1_n109 ) , .A2( u1_u5_u1_n110 ) , .A1( u1_u5_u1_n111 ) );
  AOI21_X1 u1_u5_u1_U89 (.ZN( u1_u5_u1_n110 ) , .A( u1_u5_u1_n116 ) , .B1( u1_u5_u1_n152 ) , .B2( u1_u5_u1_n160 ) );
  OAI21_X1 u1_u5_u1_U9 (.ZN( u1_u5_u1_n101 ) , .B1( u1_u5_u1_n141 ) , .A( u1_u5_u1_n146 ) , .B2( u1_u5_u1_n183 ) );
  AOI21_X1 u1_u5_u1_U90 (.ZN( u1_u5_u1_n111 ) , .A( u1_u5_u1_n128 ) , .B2( u1_u5_u1_n131 ) , .B1( u1_u5_u1_n135 ) );
  NAND4_X1 u1_u5_u1_U91 (.ZN( u1_out5_2 ) , .A4( u1_u5_u1_n142 ) , .A3( u1_u5_u1_n143 ) , .A2( u1_u5_u1_n144 ) , .A1( u1_u5_u1_n179 ) );
  OAI21_X1 u1_u5_u1_U92 (.B2( u1_u5_u1_n132 ) , .ZN( u1_u5_u1_n144 ) , .A( u1_u5_u1_n146 ) , .B1( u1_u5_u1_n180 ) );
  INV_X1 u1_u5_u1_U93 (.A( u1_u5_u1_n130 ) , .ZN( u1_u5_u1_n179 ) );
  NAND4_X1 u1_u5_u1_U94 (.ZN( u1_out5_28 ) , .A4( u1_u5_u1_n124 ) , .A3( u1_u5_u1_n125 ) , .A2( u1_u5_u1_n126 ) , .A1( u1_u5_u1_n127 ) );
  OAI21_X1 u1_u5_u1_U95 (.ZN( u1_u5_u1_n127 ) , .B2( u1_u5_u1_n139 ) , .B1( u1_u5_u1_n175 ) , .A( u1_u5_u1_n183 ) );
  OAI21_X1 u1_u5_u1_U96 (.ZN( u1_u5_u1_n126 ) , .B2( u1_u5_u1_n140 ) , .A( u1_u5_u1_n146 ) , .B1( u1_u5_u1_n178 ) );
  NAND3_X1 u1_u5_u1_U97 (.A3( u1_u5_u1_n149 ) , .A2( u1_u5_u1_n150 ) , .A1( u1_u5_u1_n151 ) , .ZN( u1_u5_u1_n164 ) );
  NAND3_X1 u1_u5_u1_U98 (.A3( u1_u5_u1_n134 ) , .A2( u1_u5_u1_n135 ) , .ZN( u1_u5_u1_n136 ) , .A1( u1_u5_u1_n151 ) );
  NAND3_X1 u1_u5_u1_U99 (.A1( u1_u5_u1_n133 ) , .ZN( u1_u5_u1_n137 ) , .A2( u1_u5_u1_n154 ) , .A3( u1_u5_u1_n181 ) );
  OAI22_X1 u1_u5_u3_U10 (.B1( u1_u5_u3_n113 ) , .A2( u1_u5_u3_n135 ) , .A1( u1_u5_u3_n150 ) , .B2( u1_u5_u3_n164 ) , .ZN( u1_u5_u3_n98 ) );
  OAI211_X1 u1_u5_u3_U11 (.B( u1_u5_u3_n106 ) , .ZN( u1_u5_u3_n119 ) , .C2( u1_u5_u3_n128 ) , .C1( u1_u5_u3_n167 ) , .A( u1_u5_u3_n181 ) );
  AOI221_X1 u1_u5_u3_U12 (.C1( u1_u5_u3_n105 ) , .ZN( u1_u5_u3_n106 ) , .A( u1_u5_u3_n131 ) , .B2( u1_u5_u3_n132 ) , .C2( u1_u5_u3_n133 ) , .B1( u1_u5_u3_n169 ) );
  INV_X1 u1_u5_u3_U13 (.ZN( u1_u5_u3_n181 ) , .A( u1_u5_u3_n98 ) );
  NAND2_X1 u1_u5_u3_U14 (.ZN( u1_u5_u3_n105 ) , .A2( u1_u5_u3_n130 ) , .A1( u1_u5_u3_n155 ) );
  AOI22_X1 u1_u5_u3_U15 (.B1( u1_u5_u3_n115 ) , .A2( u1_u5_u3_n116 ) , .ZN( u1_u5_u3_n123 ) , .B2( u1_u5_u3_n133 ) , .A1( u1_u5_u3_n169 ) );
  NAND2_X1 u1_u5_u3_U16 (.ZN( u1_u5_u3_n116 ) , .A2( u1_u5_u3_n151 ) , .A1( u1_u5_u3_n182 ) );
  NOR2_X1 u1_u5_u3_U17 (.ZN( u1_u5_u3_n126 ) , .A2( u1_u5_u3_n150 ) , .A1( u1_u5_u3_n164 ) );
  AOI21_X1 u1_u5_u3_U18 (.ZN( u1_u5_u3_n112 ) , .B2( u1_u5_u3_n146 ) , .B1( u1_u5_u3_n155 ) , .A( u1_u5_u3_n167 ) );
  NAND2_X1 u1_u5_u3_U19 (.A1( u1_u5_u3_n135 ) , .ZN( u1_u5_u3_n142 ) , .A2( u1_u5_u3_n164 ) );
  NAND2_X1 u1_u5_u3_U20 (.ZN( u1_u5_u3_n132 ) , .A2( u1_u5_u3_n152 ) , .A1( u1_u5_u3_n156 ) );
  AND2_X1 u1_u5_u3_U21 (.A2( u1_u5_u3_n113 ) , .A1( u1_u5_u3_n114 ) , .ZN( u1_u5_u3_n151 ) );
  INV_X1 u1_u5_u3_U22 (.A( u1_u5_u3_n133 ) , .ZN( u1_u5_u3_n165 ) );
  INV_X1 u1_u5_u3_U23 (.A( u1_u5_u3_n135 ) , .ZN( u1_u5_u3_n170 ) );
  NAND2_X1 u1_u5_u3_U24 (.A1( u1_u5_u3_n107 ) , .A2( u1_u5_u3_n108 ) , .ZN( u1_u5_u3_n140 ) );
  NAND2_X1 u1_u5_u3_U25 (.ZN( u1_u5_u3_n117 ) , .A1( u1_u5_u3_n124 ) , .A2( u1_u5_u3_n148 ) );
  NAND2_X1 u1_u5_u3_U26 (.ZN( u1_u5_u3_n143 ) , .A1( u1_u5_u3_n165 ) , .A2( u1_u5_u3_n167 ) );
  INV_X1 u1_u5_u3_U27 (.A( u1_u5_u3_n130 ) , .ZN( u1_u5_u3_n177 ) );
  INV_X1 u1_u5_u3_U28 (.A( u1_u5_u3_n128 ) , .ZN( u1_u5_u3_n176 ) );
  INV_X1 u1_u5_u3_U29 (.A( u1_u5_u3_n155 ) , .ZN( u1_u5_u3_n174 ) );
  INV_X1 u1_u5_u3_U3 (.A( u1_u5_u3_n129 ) , .ZN( u1_u5_u3_n183 ) );
  INV_X1 u1_u5_u3_U30 (.A( u1_u5_u3_n139 ) , .ZN( u1_u5_u3_n185 ) );
  NOR2_X1 u1_u5_u3_U31 (.ZN( u1_u5_u3_n135 ) , .A2( u1_u5_u3_n141 ) , .A1( u1_u5_u3_n169 ) );
  OAI222_X1 u1_u5_u3_U32 (.C2( u1_u5_u3_n107 ) , .A2( u1_u5_u3_n108 ) , .B1( u1_u5_u3_n135 ) , .ZN( u1_u5_u3_n138 ) , .B2( u1_u5_u3_n146 ) , .C1( u1_u5_u3_n154 ) , .A1( u1_u5_u3_n164 ) );
  NOR4_X1 u1_u5_u3_U33 (.A4( u1_u5_u3_n157 ) , .A3( u1_u5_u3_n158 ) , .A2( u1_u5_u3_n159 ) , .A1( u1_u5_u3_n160 ) , .ZN( u1_u5_u3_n161 ) );
  AOI21_X1 u1_u5_u3_U34 (.B2( u1_u5_u3_n152 ) , .B1( u1_u5_u3_n153 ) , .ZN( u1_u5_u3_n158 ) , .A( u1_u5_u3_n164 ) );
  AOI21_X1 u1_u5_u3_U35 (.A( u1_u5_u3_n154 ) , .B2( u1_u5_u3_n155 ) , .B1( u1_u5_u3_n156 ) , .ZN( u1_u5_u3_n157 ) );
  AOI21_X1 u1_u5_u3_U36 (.A( u1_u5_u3_n149 ) , .B2( u1_u5_u3_n150 ) , .B1( u1_u5_u3_n151 ) , .ZN( u1_u5_u3_n159 ) );
  AOI211_X1 u1_u5_u3_U37 (.ZN( u1_u5_u3_n109 ) , .A( u1_u5_u3_n119 ) , .C2( u1_u5_u3_n129 ) , .B( u1_u5_u3_n138 ) , .C1( u1_u5_u3_n141 ) );
  AOI211_X1 u1_u5_u3_U38 (.B( u1_u5_u3_n119 ) , .A( u1_u5_u3_n120 ) , .C2( u1_u5_u3_n121 ) , .ZN( u1_u5_u3_n122 ) , .C1( u1_u5_u3_n179 ) );
  INV_X1 u1_u5_u3_U39 (.A( u1_u5_u3_n156 ) , .ZN( u1_u5_u3_n179 ) );
  INV_X1 u1_u5_u3_U4 (.A( u1_u5_u3_n140 ) , .ZN( u1_u5_u3_n182 ) );
  OAI22_X1 u1_u5_u3_U40 (.B1( u1_u5_u3_n118 ) , .ZN( u1_u5_u3_n120 ) , .A1( u1_u5_u3_n135 ) , .B2( u1_u5_u3_n154 ) , .A2( u1_u5_u3_n178 ) );
  AND3_X1 u1_u5_u3_U41 (.ZN( u1_u5_u3_n118 ) , .A2( u1_u5_u3_n124 ) , .A1( u1_u5_u3_n144 ) , .A3( u1_u5_u3_n152 ) );
  INV_X1 u1_u5_u3_U42 (.A( u1_u5_u3_n121 ) , .ZN( u1_u5_u3_n164 ) );
  NAND2_X1 u1_u5_u3_U43 (.ZN( u1_u5_u3_n133 ) , .A1( u1_u5_u3_n154 ) , .A2( u1_u5_u3_n164 ) );
  OAI211_X1 u1_u5_u3_U44 (.B( u1_u5_u3_n127 ) , .ZN( u1_u5_u3_n139 ) , .C1( u1_u5_u3_n150 ) , .C2( u1_u5_u3_n154 ) , .A( u1_u5_u3_n184 ) );
  INV_X1 u1_u5_u3_U45 (.A( u1_u5_u3_n125 ) , .ZN( u1_u5_u3_n184 ) );
  AOI221_X1 u1_u5_u3_U46 (.A( u1_u5_u3_n126 ) , .ZN( u1_u5_u3_n127 ) , .C2( u1_u5_u3_n132 ) , .C1( u1_u5_u3_n169 ) , .B2( u1_u5_u3_n170 ) , .B1( u1_u5_u3_n174 ) );
  OAI22_X1 u1_u5_u3_U47 (.A1( u1_u5_u3_n124 ) , .ZN( u1_u5_u3_n125 ) , .B2( u1_u5_u3_n145 ) , .A2( u1_u5_u3_n165 ) , .B1( u1_u5_u3_n167 ) );
  NOR2_X1 u1_u5_u3_U48 (.A1( u1_u5_u3_n113 ) , .ZN( u1_u5_u3_n131 ) , .A2( u1_u5_u3_n154 ) );
  NAND2_X1 u1_u5_u3_U49 (.A1( u1_u5_u3_n103 ) , .ZN( u1_u5_u3_n150 ) , .A2( u1_u5_u3_n99 ) );
  INV_X1 u1_u5_u3_U5 (.A( u1_u5_u3_n117 ) , .ZN( u1_u5_u3_n178 ) );
  NAND2_X1 u1_u5_u3_U50 (.A2( u1_u5_u3_n102 ) , .ZN( u1_u5_u3_n155 ) , .A1( u1_u5_u3_n97 ) );
  INV_X1 u1_u5_u3_U51 (.A( u1_u5_u3_n141 ) , .ZN( u1_u5_u3_n167 ) );
  AOI21_X1 u1_u5_u3_U52 (.B2( u1_u5_u3_n114 ) , .B1( u1_u5_u3_n146 ) , .A( u1_u5_u3_n154 ) , .ZN( u1_u5_u3_n94 ) );
  AOI21_X1 u1_u5_u3_U53 (.ZN( u1_u5_u3_n110 ) , .B2( u1_u5_u3_n142 ) , .B1( u1_u5_u3_n186 ) , .A( u1_u5_u3_n95 ) );
  INV_X1 u1_u5_u3_U54 (.A( u1_u5_u3_n145 ) , .ZN( u1_u5_u3_n186 ) );
  AOI21_X1 u1_u5_u3_U55 (.B1( u1_u5_u3_n124 ) , .A( u1_u5_u3_n149 ) , .B2( u1_u5_u3_n155 ) , .ZN( u1_u5_u3_n95 ) );
  INV_X1 u1_u5_u3_U56 (.A( u1_u5_u3_n149 ) , .ZN( u1_u5_u3_n169 ) );
  NAND2_X1 u1_u5_u3_U57 (.ZN( u1_u5_u3_n124 ) , .A1( u1_u5_u3_n96 ) , .A2( u1_u5_u3_n97 ) );
  NAND2_X1 u1_u5_u3_U58 (.A2( u1_u5_u3_n100 ) , .ZN( u1_u5_u3_n146 ) , .A1( u1_u5_u3_n96 ) );
  NAND2_X1 u1_u5_u3_U59 (.A1( u1_u5_u3_n101 ) , .ZN( u1_u5_u3_n145 ) , .A2( u1_u5_u3_n99 ) );
  AOI221_X1 u1_u5_u3_U6 (.A( u1_u5_u3_n131 ) , .C2( u1_u5_u3_n132 ) , .C1( u1_u5_u3_n133 ) , .ZN( u1_u5_u3_n134 ) , .B1( u1_u5_u3_n143 ) , .B2( u1_u5_u3_n177 ) );
  NAND2_X1 u1_u5_u3_U60 (.A1( u1_u5_u3_n100 ) , .ZN( u1_u5_u3_n156 ) , .A2( u1_u5_u3_n99 ) );
  NAND2_X1 u1_u5_u3_U61 (.A2( u1_u5_u3_n101 ) , .A1( u1_u5_u3_n104 ) , .ZN( u1_u5_u3_n148 ) );
  NAND2_X1 u1_u5_u3_U62 (.A1( u1_u5_u3_n100 ) , .A2( u1_u5_u3_n102 ) , .ZN( u1_u5_u3_n128 ) );
  NAND2_X1 u1_u5_u3_U63 (.A2( u1_u5_u3_n101 ) , .A1( u1_u5_u3_n102 ) , .ZN( u1_u5_u3_n152 ) );
  NAND2_X1 u1_u5_u3_U64 (.A2( u1_u5_u3_n101 ) , .ZN( u1_u5_u3_n114 ) , .A1( u1_u5_u3_n96 ) );
  NAND2_X1 u1_u5_u3_U65 (.ZN( u1_u5_u3_n107 ) , .A1( u1_u5_u3_n97 ) , .A2( u1_u5_u3_n99 ) );
  NAND2_X1 u1_u5_u3_U66 (.A2( u1_u5_u3_n100 ) , .A1( u1_u5_u3_n104 ) , .ZN( u1_u5_u3_n113 ) );
  NAND2_X1 u1_u5_u3_U67 (.A1( u1_u5_u3_n104 ) , .ZN( u1_u5_u3_n153 ) , .A2( u1_u5_u3_n97 ) );
  NAND2_X1 u1_u5_u3_U68 (.A2( u1_u5_u3_n103 ) , .A1( u1_u5_u3_n104 ) , .ZN( u1_u5_u3_n130 ) );
  NAND2_X1 u1_u5_u3_U69 (.A2( u1_u5_u3_n103 ) , .ZN( u1_u5_u3_n144 ) , .A1( u1_u5_u3_n96 ) );
  OAI22_X1 u1_u5_u3_U7 (.B2( u1_u5_u3_n147 ) , .A2( u1_u5_u3_n148 ) , .ZN( u1_u5_u3_n160 ) , .B1( u1_u5_u3_n165 ) , .A1( u1_u5_u3_n168 ) );
  NAND2_X1 u1_u5_u3_U70 (.A1( u1_u5_u3_n102 ) , .A2( u1_u5_u3_n103 ) , .ZN( u1_u5_u3_n108 ) );
  NOR2_X1 u1_u5_u3_U71 (.A2( u1_u5_X_19 ) , .A1( u1_u5_X_20 ) , .ZN( u1_u5_u3_n99 ) );
  NOR2_X1 u1_u5_u3_U72 (.A2( u1_u5_X_21 ) , .A1( u1_u5_X_24 ) , .ZN( u1_u5_u3_n103 ) );
  NOR2_X1 u1_u5_u3_U73 (.A2( u1_u5_X_24 ) , .A1( u1_u5_u3_n171 ) , .ZN( u1_u5_u3_n97 ) );
  NOR2_X1 u1_u5_u3_U74 (.A2( u1_u5_X_23 ) , .ZN( u1_u5_u3_n141 ) , .A1( u1_u5_u3_n166 ) );
  NOR2_X1 u1_u5_u3_U75 (.A2( u1_u5_X_19 ) , .A1( u1_u5_u3_n172 ) , .ZN( u1_u5_u3_n96 ) );
  NAND2_X1 u1_u5_u3_U76 (.A1( u1_u5_X_22 ) , .A2( u1_u5_X_23 ) , .ZN( u1_u5_u3_n154 ) );
  NAND2_X1 u1_u5_u3_U77 (.A1( u1_u5_X_23 ) , .ZN( u1_u5_u3_n149 ) , .A2( u1_u5_u3_n166 ) );
  NOR2_X1 u1_u5_u3_U78 (.A2( u1_u5_X_22 ) , .A1( u1_u5_X_23 ) , .ZN( u1_u5_u3_n121 ) );
  AND2_X1 u1_u5_u3_U79 (.A1( u1_u5_X_24 ) , .ZN( u1_u5_u3_n101 ) , .A2( u1_u5_u3_n171 ) );
  AND3_X1 u1_u5_u3_U8 (.A3( u1_u5_u3_n144 ) , .A2( u1_u5_u3_n145 ) , .A1( u1_u5_u3_n146 ) , .ZN( u1_u5_u3_n147 ) );
  AND2_X1 u1_u5_u3_U80 (.A1( u1_u5_X_19 ) , .ZN( u1_u5_u3_n102 ) , .A2( u1_u5_u3_n172 ) );
  AND2_X1 u1_u5_u3_U81 (.A1( u1_u5_X_21 ) , .A2( u1_u5_X_24 ) , .ZN( u1_u5_u3_n100 ) );
  AND2_X1 u1_u5_u3_U82 (.A2( u1_u5_X_19 ) , .A1( u1_u5_X_20 ) , .ZN( u1_u5_u3_n104 ) );
  INV_X1 u1_u5_u3_U83 (.A( u1_u5_X_22 ) , .ZN( u1_u5_u3_n166 ) );
  INV_X1 u1_u5_u3_U84 (.A( u1_u5_X_21 ) , .ZN( u1_u5_u3_n171 ) );
  INV_X1 u1_u5_u3_U85 (.A( u1_u5_X_20 ) , .ZN( u1_u5_u3_n172 ) );
  NAND4_X1 u1_u5_u3_U86 (.ZN( u1_out5_26 ) , .A4( u1_u5_u3_n109 ) , .A3( u1_u5_u3_n110 ) , .A2( u1_u5_u3_n111 ) , .A1( u1_u5_u3_n173 ) );
  INV_X1 u1_u5_u3_U87 (.ZN( u1_u5_u3_n173 ) , .A( u1_u5_u3_n94 ) );
  OAI21_X1 u1_u5_u3_U88 (.ZN( u1_u5_u3_n111 ) , .B2( u1_u5_u3_n117 ) , .A( u1_u5_u3_n133 ) , .B1( u1_u5_u3_n176 ) );
  NAND4_X1 u1_u5_u3_U89 (.ZN( u1_out5_20 ) , .A4( u1_u5_u3_n122 ) , .A3( u1_u5_u3_n123 ) , .A1( u1_u5_u3_n175 ) , .A2( u1_u5_u3_n180 ) );
  INV_X1 u1_u5_u3_U9 (.A( u1_u5_u3_n143 ) , .ZN( u1_u5_u3_n168 ) );
  INV_X1 u1_u5_u3_U90 (.A( u1_u5_u3_n126 ) , .ZN( u1_u5_u3_n180 ) );
  INV_X1 u1_u5_u3_U91 (.A( u1_u5_u3_n112 ) , .ZN( u1_u5_u3_n175 ) );
  OR4_X1 u1_u5_u3_U92 (.ZN( u1_out5_10 ) , .A4( u1_u5_u3_n136 ) , .A3( u1_u5_u3_n137 ) , .A1( u1_u5_u3_n138 ) , .A2( u1_u5_u3_n139 ) );
  OAI222_X1 u1_u5_u3_U93 (.C1( u1_u5_u3_n128 ) , .ZN( u1_u5_u3_n137 ) , .B1( u1_u5_u3_n148 ) , .A2( u1_u5_u3_n150 ) , .B2( u1_u5_u3_n154 ) , .C2( u1_u5_u3_n164 ) , .A1( u1_u5_u3_n167 ) );
  OAI221_X1 u1_u5_u3_U94 (.A( u1_u5_u3_n134 ) , .B2( u1_u5_u3_n135 ) , .ZN( u1_u5_u3_n136 ) , .C1( u1_u5_u3_n149 ) , .B1( u1_u5_u3_n151 ) , .C2( u1_u5_u3_n183 ) );
  NAND4_X1 u1_u5_u3_U95 (.ZN( u1_out5_1 ) , .A4( u1_u5_u3_n161 ) , .A3( u1_u5_u3_n162 ) , .A2( u1_u5_u3_n163 ) , .A1( u1_u5_u3_n185 ) );
  NAND2_X1 u1_u5_u3_U96 (.ZN( u1_u5_u3_n163 ) , .A2( u1_u5_u3_n170 ) , .A1( u1_u5_u3_n176 ) );
  AOI22_X1 u1_u5_u3_U97 (.B2( u1_u5_u3_n140 ) , .B1( u1_u5_u3_n141 ) , .A2( u1_u5_u3_n142 ) , .ZN( u1_u5_u3_n162 ) , .A1( u1_u5_u3_n177 ) );
  NAND3_X1 u1_u5_u3_U98 (.A1( u1_u5_u3_n114 ) , .ZN( u1_u5_u3_n115 ) , .A2( u1_u5_u3_n145 ) , .A3( u1_u5_u3_n153 ) );
  NAND3_X1 u1_u5_u3_U99 (.ZN( u1_u5_u3_n129 ) , .A2( u1_u5_u3_n144 ) , .A1( u1_u5_u3_n153 ) , .A3( u1_u5_u3_n182 ) );
  INV_X1 u1_u5_u5_U10 (.A( u1_u5_u5_n121 ) , .ZN( u1_u5_u5_n177 ) );
  NOR3_X1 u1_u5_u5_U100 (.A3( u1_u5_u5_n141 ) , .A1( u1_u5_u5_n142 ) , .ZN( u1_u5_u5_n143 ) , .A2( u1_u5_u5_n191 ) );
  NAND4_X1 u1_u5_u5_U101 (.ZN( u1_out5_4 ) , .A4( u1_u5_u5_n112 ) , .A2( u1_u5_u5_n113 ) , .A1( u1_u5_u5_n114 ) , .A3( u1_u5_u5_n195 ) );
  AOI211_X1 u1_u5_u5_U102 (.A( u1_u5_u5_n110 ) , .C1( u1_u5_u5_n111 ) , .ZN( u1_u5_u5_n112 ) , .B( u1_u5_u5_n118 ) , .C2( u1_u5_u5_n177 ) );
  AOI222_X1 u1_u5_u5_U103 (.ZN( u1_u5_u5_n113 ) , .A1( u1_u5_u5_n131 ) , .C1( u1_u5_u5_n148 ) , .B2( u1_u5_u5_n174 ) , .C2( u1_u5_u5_n178 ) , .A2( u1_u5_u5_n179 ) , .B1( u1_u5_u5_n99 ) );
  NAND3_X1 u1_u5_u5_U104 (.A2( u1_u5_u5_n154 ) , .A3( u1_u5_u5_n158 ) , .A1( u1_u5_u5_n161 ) , .ZN( u1_u5_u5_n99 ) );
  NOR2_X1 u1_u5_u5_U11 (.ZN( u1_u5_u5_n160 ) , .A2( u1_u5_u5_n173 ) , .A1( u1_u5_u5_n177 ) );
  INV_X1 u1_u5_u5_U12 (.A( u1_u5_u5_n150 ) , .ZN( u1_u5_u5_n174 ) );
  AOI21_X1 u1_u5_u5_U13 (.A( u1_u5_u5_n160 ) , .B2( u1_u5_u5_n161 ) , .ZN( u1_u5_u5_n162 ) , .B1( u1_u5_u5_n192 ) );
  INV_X1 u1_u5_u5_U14 (.A( u1_u5_u5_n159 ) , .ZN( u1_u5_u5_n192 ) );
  AOI21_X1 u1_u5_u5_U15 (.A( u1_u5_u5_n156 ) , .B2( u1_u5_u5_n157 ) , .B1( u1_u5_u5_n158 ) , .ZN( u1_u5_u5_n163 ) );
  AOI21_X1 u1_u5_u5_U16 (.B2( u1_u5_u5_n139 ) , .B1( u1_u5_u5_n140 ) , .ZN( u1_u5_u5_n141 ) , .A( u1_u5_u5_n150 ) );
  OAI21_X1 u1_u5_u5_U17 (.A( u1_u5_u5_n133 ) , .B2( u1_u5_u5_n134 ) , .B1( u1_u5_u5_n135 ) , .ZN( u1_u5_u5_n142 ) );
  OAI21_X1 u1_u5_u5_U18 (.ZN( u1_u5_u5_n133 ) , .B2( u1_u5_u5_n147 ) , .A( u1_u5_u5_n173 ) , .B1( u1_u5_u5_n188 ) );
  NAND2_X1 u1_u5_u5_U19 (.A2( u1_u5_u5_n119 ) , .A1( u1_u5_u5_n123 ) , .ZN( u1_u5_u5_n137 ) );
  INV_X1 u1_u5_u5_U20 (.A( u1_u5_u5_n155 ) , .ZN( u1_u5_u5_n194 ) );
  NAND2_X1 u1_u5_u5_U21 (.A1( u1_u5_u5_n121 ) , .ZN( u1_u5_u5_n132 ) , .A2( u1_u5_u5_n172 ) );
  NAND2_X1 u1_u5_u5_U22 (.A2( u1_u5_u5_n122 ) , .ZN( u1_u5_u5_n136 ) , .A1( u1_u5_u5_n154 ) );
  NAND2_X1 u1_u5_u5_U23 (.A2( u1_u5_u5_n119 ) , .A1( u1_u5_u5_n120 ) , .ZN( u1_u5_u5_n159 ) );
  INV_X1 u1_u5_u5_U24 (.A( u1_u5_u5_n156 ) , .ZN( u1_u5_u5_n175 ) );
  INV_X1 u1_u5_u5_U25 (.A( u1_u5_u5_n158 ) , .ZN( u1_u5_u5_n188 ) );
  INV_X1 u1_u5_u5_U26 (.A( u1_u5_u5_n152 ) , .ZN( u1_u5_u5_n179 ) );
  INV_X1 u1_u5_u5_U27 (.A( u1_u5_u5_n140 ) , .ZN( u1_u5_u5_n182 ) );
  INV_X1 u1_u5_u5_U28 (.A( u1_u5_u5_n151 ) , .ZN( u1_u5_u5_n183 ) );
  INV_X1 u1_u5_u5_U29 (.A( u1_u5_u5_n123 ) , .ZN( u1_u5_u5_n185 ) );
  NOR2_X1 u1_u5_u5_U3 (.ZN( u1_u5_u5_n134 ) , .A1( u1_u5_u5_n183 ) , .A2( u1_u5_u5_n190 ) );
  INV_X1 u1_u5_u5_U30 (.A( u1_u5_u5_n161 ) , .ZN( u1_u5_u5_n184 ) );
  INV_X1 u1_u5_u5_U31 (.A( u1_u5_u5_n139 ) , .ZN( u1_u5_u5_n189 ) );
  INV_X1 u1_u5_u5_U32 (.A( u1_u5_u5_n157 ) , .ZN( u1_u5_u5_n190 ) );
  INV_X1 u1_u5_u5_U33 (.A( u1_u5_u5_n120 ) , .ZN( u1_u5_u5_n193 ) );
  NAND2_X1 u1_u5_u5_U34 (.ZN( u1_u5_u5_n111 ) , .A1( u1_u5_u5_n140 ) , .A2( u1_u5_u5_n155 ) );
  NOR2_X1 u1_u5_u5_U35 (.ZN( u1_u5_u5_n100 ) , .A1( u1_u5_u5_n170 ) , .A2( u1_u5_u5_n180 ) );
  INV_X1 u1_u5_u5_U36 (.A( u1_u5_u5_n117 ) , .ZN( u1_u5_u5_n196 ) );
  OAI221_X1 u1_u5_u5_U37 (.A( u1_u5_u5_n116 ) , .ZN( u1_u5_u5_n117 ) , .B2( u1_u5_u5_n119 ) , .C1( u1_u5_u5_n153 ) , .C2( u1_u5_u5_n158 ) , .B1( u1_u5_u5_n172 ) );
  AOI222_X1 u1_u5_u5_U38 (.ZN( u1_u5_u5_n116 ) , .B2( u1_u5_u5_n145 ) , .C1( u1_u5_u5_n148 ) , .A2( u1_u5_u5_n174 ) , .C2( u1_u5_u5_n177 ) , .B1( u1_u5_u5_n187 ) , .A1( u1_u5_u5_n193 ) );
  INV_X1 u1_u5_u5_U39 (.A( u1_u5_u5_n115 ) , .ZN( u1_u5_u5_n187 ) );
  INV_X1 u1_u5_u5_U4 (.A( u1_u5_u5_n138 ) , .ZN( u1_u5_u5_n191 ) );
  AOI22_X1 u1_u5_u5_U40 (.B2( u1_u5_u5_n131 ) , .A2( u1_u5_u5_n146 ) , .ZN( u1_u5_u5_n169 ) , .B1( u1_u5_u5_n174 ) , .A1( u1_u5_u5_n185 ) );
  NOR2_X1 u1_u5_u5_U41 (.A1( u1_u5_u5_n146 ) , .ZN( u1_u5_u5_n150 ) , .A2( u1_u5_u5_n173 ) );
  AOI21_X1 u1_u5_u5_U42 (.A( u1_u5_u5_n118 ) , .B2( u1_u5_u5_n145 ) , .ZN( u1_u5_u5_n168 ) , .B1( u1_u5_u5_n186 ) );
  INV_X1 u1_u5_u5_U43 (.A( u1_u5_u5_n122 ) , .ZN( u1_u5_u5_n186 ) );
  NOR2_X1 u1_u5_u5_U44 (.A1( u1_u5_u5_n146 ) , .ZN( u1_u5_u5_n152 ) , .A2( u1_u5_u5_n176 ) );
  NOR2_X1 u1_u5_u5_U45 (.A1( u1_u5_u5_n115 ) , .ZN( u1_u5_u5_n118 ) , .A2( u1_u5_u5_n153 ) );
  NOR2_X1 u1_u5_u5_U46 (.A2( u1_u5_u5_n145 ) , .ZN( u1_u5_u5_n156 ) , .A1( u1_u5_u5_n174 ) );
  NOR2_X1 u1_u5_u5_U47 (.ZN( u1_u5_u5_n121 ) , .A2( u1_u5_u5_n145 ) , .A1( u1_u5_u5_n176 ) );
  AOI22_X1 u1_u5_u5_U48 (.ZN( u1_u5_u5_n114 ) , .A2( u1_u5_u5_n137 ) , .A1( u1_u5_u5_n145 ) , .B2( u1_u5_u5_n175 ) , .B1( u1_u5_u5_n193 ) );
  OAI211_X1 u1_u5_u5_U49 (.B( u1_u5_u5_n124 ) , .A( u1_u5_u5_n125 ) , .C2( u1_u5_u5_n126 ) , .C1( u1_u5_u5_n127 ) , .ZN( u1_u5_u5_n128 ) );
  OAI21_X1 u1_u5_u5_U5 (.B2( u1_u5_u5_n136 ) , .B1( u1_u5_u5_n137 ) , .ZN( u1_u5_u5_n138 ) , .A( u1_u5_u5_n177 ) );
  NOR3_X1 u1_u5_u5_U50 (.ZN( u1_u5_u5_n127 ) , .A1( u1_u5_u5_n136 ) , .A3( u1_u5_u5_n148 ) , .A2( u1_u5_u5_n182 ) );
  OAI21_X1 u1_u5_u5_U51 (.ZN( u1_u5_u5_n124 ) , .A( u1_u5_u5_n177 ) , .B2( u1_u5_u5_n183 ) , .B1( u1_u5_u5_n189 ) );
  OAI21_X1 u1_u5_u5_U52 (.ZN( u1_u5_u5_n125 ) , .A( u1_u5_u5_n174 ) , .B2( u1_u5_u5_n185 ) , .B1( u1_u5_u5_n190 ) );
  AOI21_X1 u1_u5_u5_U53 (.A( u1_u5_u5_n153 ) , .B2( u1_u5_u5_n154 ) , .B1( u1_u5_u5_n155 ) , .ZN( u1_u5_u5_n164 ) );
  AOI21_X1 u1_u5_u5_U54 (.ZN( u1_u5_u5_n110 ) , .B1( u1_u5_u5_n122 ) , .B2( u1_u5_u5_n139 ) , .A( u1_u5_u5_n153 ) );
  INV_X1 u1_u5_u5_U55 (.A( u1_u5_u5_n153 ) , .ZN( u1_u5_u5_n176 ) );
  INV_X1 u1_u5_u5_U56 (.A( u1_u5_u5_n126 ) , .ZN( u1_u5_u5_n173 ) );
  AND2_X1 u1_u5_u5_U57 (.A2( u1_u5_u5_n104 ) , .A1( u1_u5_u5_n107 ) , .ZN( u1_u5_u5_n147 ) );
  AND2_X1 u1_u5_u5_U58 (.A2( u1_u5_u5_n104 ) , .A1( u1_u5_u5_n108 ) , .ZN( u1_u5_u5_n148 ) );
  NAND2_X1 u1_u5_u5_U59 (.A1( u1_u5_u5_n105 ) , .A2( u1_u5_u5_n106 ) , .ZN( u1_u5_u5_n158 ) );
  INV_X1 u1_u5_u5_U6 (.A( u1_u5_u5_n135 ) , .ZN( u1_u5_u5_n178 ) );
  NAND2_X1 u1_u5_u5_U60 (.A2( u1_u5_u5_n108 ) , .A1( u1_u5_u5_n109 ) , .ZN( u1_u5_u5_n139 ) );
  NAND2_X1 u1_u5_u5_U61 (.A1( u1_u5_u5_n106 ) , .A2( u1_u5_u5_n108 ) , .ZN( u1_u5_u5_n119 ) );
  NAND2_X1 u1_u5_u5_U62 (.A2( u1_u5_u5_n103 ) , .A1( u1_u5_u5_n105 ) , .ZN( u1_u5_u5_n140 ) );
  NAND2_X1 u1_u5_u5_U63 (.A2( u1_u5_u5_n104 ) , .A1( u1_u5_u5_n105 ) , .ZN( u1_u5_u5_n155 ) );
  NAND2_X1 u1_u5_u5_U64 (.A2( u1_u5_u5_n106 ) , .A1( u1_u5_u5_n107 ) , .ZN( u1_u5_u5_n122 ) );
  NAND2_X1 u1_u5_u5_U65 (.A2( u1_u5_u5_n100 ) , .A1( u1_u5_u5_n106 ) , .ZN( u1_u5_u5_n115 ) );
  NAND2_X1 u1_u5_u5_U66 (.A2( u1_u5_u5_n100 ) , .A1( u1_u5_u5_n103 ) , .ZN( u1_u5_u5_n161 ) );
  NAND2_X1 u1_u5_u5_U67 (.A1( u1_u5_u5_n105 ) , .A2( u1_u5_u5_n109 ) , .ZN( u1_u5_u5_n154 ) );
  INV_X1 u1_u5_u5_U68 (.A( u1_u5_u5_n146 ) , .ZN( u1_u5_u5_n172 ) );
  NAND2_X1 u1_u5_u5_U69 (.A1( u1_u5_u5_n103 ) , .A2( u1_u5_u5_n108 ) , .ZN( u1_u5_u5_n123 ) );
  OAI22_X1 u1_u5_u5_U7 (.B2( u1_u5_u5_n149 ) , .B1( u1_u5_u5_n150 ) , .A2( u1_u5_u5_n151 ) , .A1( u1_u5_u5_n152 ) , .ZN( u1_u5_u5_n165 ) );
  NAND2_X1 u1_u5_u5_U70 (.A2( u1_u5_u5_n103 ) , .A1( u1_u5_u5_n107 ) , .ZN( u1_u5_u5_n151 ) );
  NAND2_X1 u1_u5_u5_U71 (.A2( u1_u5_u5_n107 ) , .A1( u1_u5_u5_n109 ) , .ZN( u1_u5_u5_n120 ) );
  NAND2_X1 u1_u5_u5_U72 (.A2( u1_u5_u5_n100 ) , .A1( u1_u5_u5_n109 ) , .ZN( u1_u5_u5_n157 ) );
  AND2_X1 u1_u5_u5_U73 (.A2( u1_u5_u5_n100 ) , .A1( u1_u5_u5_n104 ) , .ZN( u1_u5_u5_n131 ) );
  INV_X1 u1_u5_u5_U74 (.A( u1_u5_u5_n102 ) , .ZN( u1_u5_u5_n195 ) );
  OAI221_X1 u1_u5_u5_U75 (.A( u1_u5_u5_n101 ) , .ZN( u1_u5_u5_n102 ) , .C2( u1_u5_u5_n115 ) , .C1( u1_u5_u5_n126 ) , .B1( u1_u5_u5_n134 ) , .B2( u1_u5_u5_n160 ) );
  OAI21_X1 u1_u5_u5_U76 (.ZN( u1_u5_u5_n101 ) , .B1( u1_u5_u5_n137 ) , .A( u1_u5_u5_n146 ) , .B2( u1_u5_u5_n147 ) );
  NOR2_X1 u1_u5_u5_U77 (.A2( u1_u5_X_34 ) , .A1( u1_u5_X_35 ) , .ZN( u1_u5_u5_n145 ) );
  NOR2_X1 u1_u5_u5_U78 (.A2( u1_u5_X_34 ) , .ZN( u1_u5_u5_n146 ) , .A1( u1_u5_u5_n171 ) );
  NOR2_X1 u1_u5_u5_U79 (.A2( u1_u5_X_31 ) , .A1( u1_u5_X_32 ) , .ZN( u1_u5_u5_n103 ) );
  NOR3_X1 u1_u5_u5_U8 (.A2( u1_u5_u5_n147 ) , .A1( u1_u5_u5_n148 ) , .ZN( u1_u5_u5_n149 ) , .A3( u1_u5_u5_n194 ) );
  NOR2_X1 u1_u5_u5_U80 (.A2( u1_u5_X_36 ) , .ZN( u1_u5_u5_n105 ) , .A1( u1_u5_u5_n180 ) );
  NOR2_X1 u1_u5_u5_U81 (.A2( u1_u5_X_33 ) , .ZN( u1_u5_u5_n108 ) , .A1( u1_u5_u5_n170 ) );
  NOR2_X1 u1_u5_u5_U82 (.A2( u1_u5_X_33 ) , .A1( u1_u5_X_36 ) , .ZN( u1_u5_u5_n107 ) );
  NOR2_X1 u1_u5_u5_U83 (.A2( u1_u5_X_31 ) , .ZN( u1_u5_u5_n104 ) , .A1( u1_u5_u5_n181 ) );
  NAND2_X1 u1_u5_u5_U84 (.A2( u1_u5_X_34 ) , .A1( u1_u5_X_35 ) , .ZN( u1_u5_u5_n153 ) );
  NAND2_X1 u1_u5_u5_U85 (.A1( u1_u5_X_34 ) , .ZN( u1_u5_u5_n126 ) , .A2( u1_u5_u5_n171 ) );
  AND2_X1 u1_u5_u5_U86 (.A1( u1_u5_X_31 ) , .A2( u1_u5_X_32 ) , .ZN( u1_u5_u5_n106 ) );
  AND2_X1 u1_u5_u5_U87 (.A1( u1_u5_X_31 ) , .ZN( u1_u5_u5_n109 ) , .A2( u1_u5_u5_n181 ) );
  INV_X1 u1_u5_u5_U88 (.A( u1_u5_X_33 ) , .ZN( u1_u5_u5_n180 ) );
  INV_X1 u1_u5_u5_U89 (.A( u1_u5_X_35 ) , .ZN( u1_u5_u5_n171 ) );
  NOR2_X1 u1_u5_u5_U9 (.ZN( u1_u5_u5_n135 ) , .A1( u1_u5_u5_n173 ) , .A2( u1_u5_u5_n176 ) );
  INV_X1 u1_u5_u5_U90 (.A( u1_u5_X_36 ) , .ZN( u1_u5_u5_n170 ) );
  INV_X1 u1_u5_u5_U91 (.A( u1_u5_X_32 ) , .ZN( u1_u5_u5_n181 ) );
  NAND4_X1 u1_u5_u5_U92 (.ZN( u1_out5_29 ) , .A4( u1_u5_u5_n129 ) , .A3( u1_u5_u5_n130 ) , .A2( u1_u5_u5_n168 ) , .A1( u1_u5_u5_n196 ) );
  AOI221_X1 u1_u5_u5_U93 (.A( u1_u5_u5_n128 ) , .ZN( u1_u5_u5_n129 ) , .C2( u1_u5_u5_n132 ) , .B2( u1_u5_u5_n159 ) , .B1( u1_u5_u5_n176 ) , .C1( u1_u5_u5_n184 ) );
  AOI222_X1 u1_u5_u5_U94 (.ZN( u1_u5_u5_n130 ) , .A2( u1_u5_u5_n146 ) , .B1( u1_u5_u5_n147 ) , .C2( u1_u5_u5_n175 ) , .B2( u1_u5_u5_n179 ) , .A1( u1_u5_u5_n188 ) , .C1( u1_u5_u5_n194 ) );
  NAND4_X1 u1_u5_u5_U95 (.ZN( u1_out5_19 ) , .A4( u1_u5_u5_n166 ) , .A3( u1_u5_u5_n167 ) , .A2( u1_u5_u5_n168 ) , .A1( u1_u5_u5_n169 ) );
  AOI22_X1 u1_u5_u5_U96 (.B2( u1_u5_u5_n145 ) , .A2( u1_u5_u5_n146 ) , .ZN( u1_u5_u5_n167 ) , .B1( u1_u5_u5_n182 ) , .A1( u1_u5_u5_n189 ) );
  NOR4_X1 u1_u5_u5_U97 (.A4( u1_u5_u5_n162 ) , .A3( u1_u5_u5_n163 ) , .A2( u1_u5_u5_n164 ) , .A1( u1_u5_u5_n165 ) , .ZN( u1_u5_u5_n166 ) );
  NAND4_X1 u1_u5_u5_U98 (.ZN( u1_out5_11 ) , .A4( u1_u5_u5_n143 ) , .A3( u1_u5_u5_n144 ) , .A2( u1_u5_u5_n169 ) , .A1( u1_u5_u5_n196 ) );
  AOI22_X1 u1_u5_u5_U99 (.A2( u1_u5_u5_n132 ) , .ZN( u1_u5_u5_n144 ) , .B2( u1_u5_u5_n145 ) , .B1( u1_u5_u5_n184 ) , .A1( u1_u5_u5_n194 ) );
  OAI21_X1 u1_u5_u6_U10 (.A( u1_u5_u6_n159 ) , .B1( u1_u5_u6_n169 ) , .B2( u1_u5_u6_n173 ) , .ZN( u1_u5_u6_n90 ) );
  INV_X1 u1_u5_u6_U11 (.ZN( u1_u5_u6_n172 ) , .A( u1_u5_u6_n88 ) );
  AOI22_X1 u1_u5_u6_U12 (.A2( u1_u5_u6_n151 ) , .B2( u1_u5_u6_n161 ) , .A1( u1_u5_u6_n167 ) , .B1( u1_u5_u6_n170 ) , .ZN( u1_u5_u6_n89 ) );
  AOI21_X1 u1_u5_u6_U13 (.ZN( u1_u5_u6_n106 ) , .A( u1_u5_u6_n142 ) , .B2( u1_u5_u6_n159 ) , .B1( u1_u5_u6_n164 ) );
  INV_X1 u1_u5_u6_U14 (.A( u1_u5_u6_n155 ) , .ZN( u1_u5_u6_n161 ) );
  INV_X1 u1_u5_u6_U15 (.A( u1_u5_u6_n128 ) , .ZN( u1_u5_u6_n164 ) );
  NAND2_X1 u1_u5_u6_U16 (.ZN( u1_u5_u6_n110 ) , .A1( u1_u5_u6_n122 ) , .A2( u1_u5_u6_n129 ) );
  NAND2_X1 u1_u5_u6_U17 (.ZN( u1_u5_u6_n124 ) , .A2( u1_u5_u6_n146 ) , .A1( u1_u5_u6_n148 ) );
  INV_X1 u1_u5_u6_U18 (.A( u1_u5_u6_n132 ) , .ZN( u1_u5_u6_n171 ) );
  AND2_X1 u1_u5_u6_U19 (.A1( u1_u5_u6_n100 ) , .ZN( u1_u5_u6_n130 ) , .A2( u1_u5_u6_n147 ) );
  INV_X1 u1_u5_u6_U20 (.A( u1_u5_u6_n127 ) , .ZN( u1_u5_u6_n173 ) );
  INV_X1 u1_u5_u6_U21 (.A( u1_u5_u6_n121 ) , .ZN( u1_u5_u6_n167 ) );
  INV_X1 u1_u5_u6_U22 (.A( u1_u5_u6_n100 ) , .ZN( u1_u5_u6_n169 ) );
  INV_X1 u1_u5_u6_U23 (.A( u1_u5_u6_n123 ) , .ZN( u1_u5_u6_n170 ) );
  INV_X1 u1_u5_u6_U24 (.A( u1_u5_u6_n113 ) , .ZN( u1_u5_u6_n168 ) );
  AND2_X1 u1_u5_u6_U25 (.A1( u1_u5_u6_n107 ) , .A2( u1_u5_u6_n119 ) , .ZN( u1_u5_u6_n133 ) );
  AND2_X1 u1_u5_u6_U26 (.A2( u1_u5_u6_n121 ) , .A1( u1_u5_u6_n122 ) , .ZN( u1_u5_u6_n131 ) );
  AND3_X1 u1_u5_u6_U27 (.ZN( u1_u5_u6_n120 ) , .A2( u1_u5_u6_n127 ) , .A1( u1_u5_u6_n132 ) , .A3( u1_u5_u6_n145 ) );
  INV_X1 u1_u5_u6_U28 (.A( u1_u5_u6_n146 ) , .ZN( u1_u5_u6_n163 ) );
  AOI222_X1 u1_u5_u6_U29 (.ZN( u1_u5_u6_n114 ) , .A1( u1_u5_u6_n118 ) , .A2( u1_u5_u6_n126 ) , .B2( u1_u5_u6_n151 ) , .C2( u1_u5_u6_n159 ) , .C1( u1_u5_u6_n168 ) , .B1( u1_u5_u6_n169 ) );
  INV_X1 u1_u5_u6_U3 (.A( u1_u5_u6_n110 ) , .ZN( u1_u5_u6_n166 ) );
  NOR2_X1 u1_u5_u6_U30 (.A1( u1_u5_u6_n162 ) , .A2( u1_u5_u6_n165 ) , .ZN( u1_u5_u6_n98 ) );
  NAND2_X1 u1_u5_u6_U31 (.A1( u1_u5_u6_n144 ) , .ZN( u1_u5_u6_n151 ) , .A2( u1_u5_u6_n158 ) );
  NAND2_X1 u1_u5_u6_U32 (.ZN( u1_u5_u6_n132 ) , .A1( u1_u5_u6_n91 ) , .A2( u1_u5_u6_n97 ) );
  NOR2_X1 u1_u5_u6_U33 (.A2( u1_u5_u6_n126 ) , .ZN( u1_u5_u6_n155 ) , .A1( u1_u5_u6_n160 ) );
  NAND2_X1 u1_u5_u6_U34 (.ZN( u1_u5_u6_n146 ) , .A2( u1_u5_u6_n94 ) , .A1( u1_u5_u6_n99 ) );
  AOI21_X1 u1_u5_u6_U35 (.A( u1_u5_u6_n144 ) , .B2( u1_u5_u6_n145 ) , .B1( u1_u5_u6_n146 ) , .ZN( u1_u5_u6_n150 ) );
  INV_X1 u1_u5_u6_U36 (.A( u1_u5_u6_n111 ) , .ZN( u1_u5_u6_n158 ) );
  NAND2_X1 u1_u5_u6_U37 (.ZN( u1_u5_u6_n127 ) , .A1( u1_u5_u6_n91 ) , .A2( u1_u5_u6_n92 ) );
  NAND2_X1 u1_u5_u6_U38 (.ZN( u1_u5_u6_n129 ) , .A2( u1_u5_u6_n95 ) , .A1( u1_u5_u6_n96 ) );
  INV_X1 u1_u5_u6_U39 (.A( u1_u5_u6_n144 ) , .ZN( u1_u5_u6_n159 ) );
  INV_X1 u1_u5_u6_U4 (.A( u1_u5_u6_n142 ) , .ZN( u1_u5_u6_n174 ) );
  NAND2_X1 u1_u5_u6_U40 (.ZN( u1_u5_u6_n145 ) , .A2( u1_u5_u6_n97 ) , .A1( u1_u5_u6_n98 ) );
  NAND2_X1 u1_u5_u6_U41 (.ZN( u1_u5_u6_n148 ) , .A2( u1_u5_u6_n92 ) , .A1( u1_u5_u6_n94 ) );
  NAND2_X1 u1_u5_u6_U42 (.ZN( u1_u5_u6_n108 ) , .A2( u1_u5_u6_n139 ) , .A1( u1_u5_u6_n144 ) );
  NAND2_X1 u1_u5_u6_U43 (.ZN( u1_u5_u6_n121 ) , .A2( u1_u5_u6_n95 ) , .A1( u1_u5_u6_n97 ) );
  NAND2_X1 u1_u5_u6_U44 (.ZN( u1_u5_u6_n107 ) , .A2( u1_u5_u6_n92 ) , .A1( u1_u5_u6_n95 ) );
  AND2_X1 u1_u5_u6_U45 (.ZN( u1_u5_u6_n118 ) , .A2( u1_u5_u6_n91 ) , .A1( u1_u5_u6_n99 ) );
  AOI22_X1 u1_u5_u6_U46 (.B2( u1_u5_u6_n110 ) , .B1( u1_u5_u6_n111 ) , .A1( u1_u5_u6_n112 ) , .ZN( u1_u5_u6_n115 ) , .A2( u1_u5_u6_n161 ) );
  NAND4_X1 u1_u5_u6_U47 (.A3( u1_u5_u6_n109 ) , .ZN( u1_u5_u6_n112 ) , .A4( u1_u5_u6_n132 ) , .A2( u1_u5_u6_n147 ) , .A1( u1_u5_u6_n166 ) );
  NOR2_X1 u1_u5_u6_U48 (.ZN( u1_u5_u6_n109 ) , .A1( u1_u5_u6_n170 ) , .A2( u1_u5_u6_n173 ) );
  NAND2_X1 u1_u5_u6_U49 (.ZN( u1_u5_u6_n147 ) , .A2( u1_u5_u6_n98 ) , .A1( u1_u5_u6_n99 ) );
  NAND2_X1 u1_u5_u6_U5 (.A2( u1_u5_u6_n143 ) , .ZN( u1_u5_u6_n152 ) , .A1( u1_u5_u6_n166 ) );
  NAND2_X1 u1_u5_u6_U50 (.ZN( u1_u5_u6_n128 ) , .A1( u1_u5_u6_n94 ) , .A2( u1_u5_u6_n96 ) );
  AOI211_X1 u1_u5_u6_U51 (.B( u1_u5_u6_n134 ) , .A( u1_u5_u6_n135 ) , .C1( u1_u5_u6_n136 ) , .ZN( u1_u5_u6_n137 ) , .C2( u1_u5_u6_n151 ) );
  AOI21_X1 u1_u5_u6_U52 (.B2( u1_u5_u6_n132 ) , .B1( u1_u5_u6_n133 ) , .ZN( u1_u5_u6_n134 ) , .A( u1_u5_u6_n158 ) );
  AOI21_X1 u1_u5_u6_U53 (.B1( u1_u5_u6_n131 ) , .ZN( u1_u5_u6_n135 ) , .A( u1_u5_u6_n144 ) , .B2( u1_u5_u6_n146 ) );
  NAND4_X1 u1_u5_u6_U54 (.A4( u1_u5_u6_n127 ) , .A3( u1_u5_u6_n128 ) , .A2( u1_u5_u6_n129 ) , .A1( u1_u5_u6_n130 ) , .ZN( u1_u5_u6_n136 ) );
  NAND2_X1 u1_u5_u6_U55 (.ZN( u1_u5_u6_n119 ) , .A2( u1_u5_u6_n95 ) , .A1( u1_u5_u6_n99 ) );
  NAND2_X1 u1_u5_u6_U56 (.ZN( u1_u5_u6_n123 ) , .A2( u1_u5_u6_n91 ) , .A1( u1_u5_u6_n96 ) );
  NAND2_X1 u1_u5_u6_U57 (.ZN( u1_u5_u6_n100 ) , .A2( u1_u5_u6_n92 ) , .A1( u1_u5_u6_n98 ) );
  NAND2_X1 u1_u5_u6_U58 (.ZN( u1_u5_u6_n122 ) , .A1( u1_u5_u6_n94 ) , .A2( u1_u5_u6_n97 ) );
  INV_X1 u1_u5_u6_U59 (.A( u1_u5_u6_n139 ) , .ZN( u1_u5_u6_n160 ) );
  AOI22_X1 u1_u5_u6_U6 (.B2( u1_u5_u6_n101 ) , .A1( u1_u5_u6_n102 ) , .ZN( u1_u5_u6_n103 ) , .B1( u1_u5_u6_n160 ) , .A2( u1_u5_u6_n161 ) );
  NAND2_X1 u1_u5_u6_U60 (.ZN( u1_u5_u6_n113 ) , .A1( u1_u5_u6_n96 ) , .A2( u1_u5_u6_n98 ) );
  NOR2_X1 u1_u5_u6_U61 (.A2( u1_u5_X_40 ) , .A1( u1_u5_X_41 ) , .ZN( u1_u5_u6_n126 ) );
  NOR2_X1 u1_u5_u6_U62 (.A2( u1_u5_X_39 ) , .A1( u1_u5_X_42 ) , .ZN( u1_u5_u6_n92 ) );
  NOR2_X1 u1_u5_u6_U63 (.A2( u1_u5_X_39 ) , .A1( u1_u5_u6_n156 ) , .ZN( u1_u5_u6_n97 ) );
  NOR2_X1 u1_u5_u6_U64 (.A2( u1_u5_X_38 ) , .A1( u1_u5_u6_n165 ) , .ZN( u1_u5_u6_n95 ) );
  NOR2_X1 u1_u5_u6_U65 (.A2( u1_u5_X_41 ) , .ZN( u1_u5_u6_n111 ) , .A1( u1_u5_u6_n157 ) );
  NOR2_X1 u1_u5_u6_U66 (.A2( u1_u5_X_37 ) , .A1( u1_u5_u6_n162 ) , .ZN( u1_u5_u6_n94 ) );
  NOR2_X1 u1_u5_u6_U67 (.A2( u1_u5_X_37 ) , .A1( u1_u5_X_38 ) , .ZN( u1_u5_u6_n91 ) );
  NAND2_X1 u1_u5_u6_U68 (.A1( u1_u5_X_41 ) , .ZN( u1_u5_u6_n144 ) , .A2( u1_u5_u6_n157 ) );
  NAND2_X1 u1_u5_u6_U69 (.A2( u1_u5_X_40 ) , .A1( u1_u5_X_41 ) , .ZN( u1_u5_u6_n139 ) );
  NOR2_X1 u1_u5_u6_U7 (.A1( u1_u5_u6_n118 ) , .ZN( u1_u5_u6_n143 ) , .A2( u1_u5_u6_n168 ) );
  AND2_X1 u1_u5_u6_U70 (.A1( u1_u5_X_39 ) , .A2( u1_u5_u6_n156 ) , .ZN( u1_u5_u6_n96 ) );
  AND2_X1 u1_u5_u6_U71 (.A1( u1_u5_X_39 ) , .A2( u1_u5_X_42 ) , .ZN( u1_u5_u6_n99 ) );
  INV_X1 u1_u5_u6_U72 (.A( u1_u5_X_40 ) , .ZN( u1_u5_u6_n157 ) );
  INV_X1 u1_u5_u6_U73 (.A( u1_u5_X_37 ) , .ZN( u1_u5_u6_n165 ) );
  INV_X1 u1_u5_u6_U74 (.A( u1_u5_X_38 ) , .ZN( u1_u5_u6_n162 ) );
  INV_X1 u1_u5_u6_U75 (.A( u1_u5_X_42 ) , .ZN( u1_u5_u6_n156 ) );
  NAND4_X1 u1_u5_u6_U76 (.ZN( u1_out5_32 ) , .A4( u1_u5_u6_n103 ) , .A3( u1_u5_u6_n104 ) , .A2( u1_u5_u6_n105 ) , .A1( u1_u5_u6_n106 ) );
  AOI22_X1 u1_u5_u6_U77 (.ZN( u1_u5_u6_n105 ) , .A2( u1_u5_u6_n108 ) , .A1( u1_u5_u6_n118 ) , .B2( u1_u5_u6_n126 ) , .B1( u1_u5_u6_n171 ) );
  AOI22_X1 u1_u5_u6_U78 (.ZN( u1_u5_u6_n104 ) , .A1( u1_u5_u6_n111 ) , .B1( u1_u5_u6_n124 ) , .B2( u1_u5_u6_n151 ) , .A2( u1_u5_u6_n93 ) );
  NAND4_X1 u1_u5_u6_U79 (.ZN( u1_out5_12 ) , .A4( u1_u5_u6_n114 ) , .A3( u1_u5_u6_n115 ) , .A2( u1_u5_u6_n116 ) , .A1( u1_u5_u6_n117 ) );
  AOI21_X1 u1_u5_u6_U8 (.B1( u1_u5_u6_n107 ) , .B2( u1_u5_u6_n132 ) , .A( u1_u5_u6_n158 ) , .ZN( u1_u5_u6_n88 ) );
  OAI22_X1 u1_u5_u6_U80 (.B2( u1_u5_u6_n111 ) , .ZN( u1_u5_u6_n116 ) , .B1( u1_u5_u6_n126 ) , .A2( u1_u5_u6_n164 ) , .A1( u1_u5_u6_n167 ) );
  OAI21_X1 u1_u5_u6_U81 (.A( u1_u5_u6_n108 ) , .ZN( u1_u5_u6_n117 ) , .B2( u1_u5_u6_n141 ) , .B1( u1_u5_u6_n163 ) );
  OAI211_X1 u1_u5_u6_U82 (.ZN( u1_out5_7 ) , .B( u1_u5_u6_n153 ) , .C2( u1_u5_u6_n154 ) , .C1( u1_u5_u6_n155 ) , .A( u1_u5_u6_n174 ) );
  NOR3_X1 u1_u5_u6_U83 (.A1( u1_u5_u6_n141 ) , .ZN( u1_u5_u6_n154 ) , .A3( u1_u5_u6_n164 ) , .A2( u1_u5_u6_n171 ) );
  AOI211_X1 u1_u5_u6_U84 (.B( u1_u5_u6_n149 ) , .A( u1_u5_u6_n150 ) , .C2( u1_u5_u6_n151 ) , .C1( u1_u5_u6_n152 ) , .ZN( u1_u5_u6_n153 ) );
  OAI211_X1 u1_u5_u6_U85 (.ZN( u1_out5_22 ) , .B( u1_u5_u6_n137 ) , .A( u1_u5_u6_n138 ) , .C2( u1_u5_u6_n139 ) , .C1( u1_u5_u6_n140 ) );
  AOI22_X1 u1_u5_u6_U86 (.B1( u1_u5_u6_n124 ) , .A2( u1_u5_u6_n125 ) , .A1( u1_u5_u6_n126 ) , .ZN( u1_u5_u6_n138 ) , .B2( u1_u5_u6_n161 ) );
  AND4_X1 u1_u5_u6_U87 (.A3( u1_u5_u6_n119 ) , .A1( u1_u5_u6_n120 ) , .A4( u1_u5_u6_n129 ) , .ZN( u1_u5_u6_n140 ) , .A2( u1_u5_u6_n143 ) );
  NAND3_X1 u1_u5_u6_U88 (.A2( u1_u5_u6_n123 ) , .ZN( u1_u5_u6_n125 ) , .A1( u1_u5_u6_n130 ) , .A3( u1_u5_u6_n131 ) );
  NAND3_X1 u1_u5_u6_U89 (.A3( u1_u5_u6_n133 ) , .ZN( u1_u5_u6_n141 ) , .A1( u1_u5_u6_n145 ) , .A2( u1_u5_u6_n148 ) );
  AOI21_X1 u1_u5_u6_U9 (.B2( u1_u5_u6_n147 ) , .B1( u1_u5_u6_n148 ) , .ZN( u1_u5_u6_n149 ) , .A( u1_u5_u6_n158 ) );
  NAND3_X1 u1_u5_u6_U90 (.ZN( u1_u5_u6_n101 ) , .A3( u1_u5_u6_n107 ) , .A2( u1_u5_u6_n121 ) , .A1( u1_u5_u6_n127 ) );
  NAND3_X1 u1_u5_u6_U91 (.ZN( u1_u5_u6_n102 ) , .A3( u1_u5_u6_n130 ) , .A2( u1_u5_u6_n145 ) , .A1( u1_u5_u6_n166 ) );
  NAND3_X1 u1_u5_u6_U92 (.A3( u1_u5_u6_n113 ) , .A1( u1_u5_u6_n119 ) , .A2( u1_u5_u6_n123 ) , .ZN( u1_u5_u6_n93 ) );
  NAND3_X1 u1_u5_u6_U93 (.ZN( u1_u5_u6_n142 ) , .A2( u1_u5_u6_n172 ) , .A3( u1_u5_u6_n89 ) , .A1( u1_u5_u6_n90 ) );
  AND3_X1 u1_u5_u7_U10 (.A3( u1_u5_u7_n110 ) , .A2( u1_u5_u7_n127 ) , .A1( u1_u5_u7_n132 ) , .ZN( u1_u5_u7_n92 ) );
  OAI21_X1 u1_u5_u7_U11 (.A( u1_u5_u7_n161 ) , .B1( u1_u5_u7_n168 ) , .B2( u1_u5_u7_n173 ) , .ZN( u1_u5_u7_n91 ) );
  AOI211_X1 u1_u5_u7_U12 (.A( u1_u5_u7_n117 ) , .ZN( u1_u5_u7_n118 ) , .C2( u1_u5_u7_n126 ) , .C1( u1_u5_u7_n177 ) , .B( u1_u5_u7_n180 ) );
  OAI22_X1 u1_u5_u7_U13 (.B1( u1_u5_u7_n115 ) , .ZN( u1_u5_u7_n117 ) , .A2( u1_u5_u7_n133 ) , .A1( u1_u5_u7_n137 ) , .B2( u1_u5_u7_n162 ) );
  INV_X1 u1_u5_u7_U14 (.A( u1_u5_u7_n116 ) , .ZN( u1_u5_u7_n180 ) );
  NOR3_X1 u1_u5_u7_U15 (.ZN( u1_u5_u7_n115 ) , .A3( u1_u5_u7_n145 ) , .A2( u1_u5_u7_n168 ) , .A1( u1_u5_u7_n169 ) );
  OAI211_X1 u1_u5_u7_U16 (.B( u1_u5_u7_n122 ) , .A( u1_u5_u7_n123 ) , .C2( u1_u5_u7_n124 ) , .ZN( u1_u5_u7_n154 ) , .C1( u1_u5_u7_n162 ) );
  AOI222_X1 u1_u5_u7_U17 (.ZN( u1_u5_u7_n122 ) , .C2( u1_u5_u7_n126 ) , .C1( u1_u5_u7_n145 ) , .B1( u1_u5_u7_n161 ) , .A2( u1_u5_u7_n165 ) , .B2( u1_u5_u7_n170 ) , .A1( u1_u5_u7_n176 ) );
  INV_X1 u1_u5_u7_U18 (.A( u1_u5_u7_n133 ) , .ZN( u1_u5_u7_n176 ) );
  NOR3_X1 u1_u5_u7_U19 (.A2( u1_u5_u7_n134 ) , .A1( u1_u5_u7_n135 ) , .ZN( u1_u5_u7_n136 ) , .A3( u1_u5_u7_n171 ) );
  NOR2_X1 u1_u5_u7_U20 (.A1( u1_u5_u7_n130 ) , .A2( u1_u5_u7_n134 ) , .ZN( u1_u5_u7_n153 ) );
  INV_X1 u1_u5_u7_U21 (.A( u1_u5_u7_n101 ) , .ZN( u1_u5_u7_n165 ) );
  NOR2_X1 u1_u5_u7_U22 (.ZN( u1_u5_u7_n111 ) , .A2( u1_u5_u7_n134 ) , .A1( u1_u5_u7_n169 ) );
  AOI21_X1 u1_u5_u7_U23 (.ZN( u1_u5_u7_n104 ) , .B2( u1_u5_u7_n112 ) , .B1( u1_u5_u7_n127 ) , .A( u1_u5_u7_n164 ) );
  AOI21_X1 u1_u5_u7_U24 (.ZN( u1_u5_u7_n106 ) , .B1( u1_u5_u7_n133 ) , .B2( u1_u5_u7_n146 ) , .A( u1_u5_u7_n162 ) );
  AOI21_X1 u1_u5_u7_U25 (.A( u1_u5_u7_n101 ) , .ZN( u1_u5_u7_n107 ) , .B2( u1_u5_u7_n128 ) , .B1( u1_u5_u7_n175 ) );
  INV_X1 u1_u5_u7_U26 (.A( u1_u5_u7_n138 ) , .ZN( u1_u5_u7_n171 ) );
  INV_X1 u1_u5_u7_U27 (.A( u1_u5_u7_n131 ) , .ZN( u1_u5_u7_n177 ) );
  INV_X1 u1_u5_u7_U28 (.A( u1_u5_u7_n110 ) , .ZN( u1_u5_u7_n174 ) );
  NAND2_X1 u1_u5_u7_U29 (.A1( u1_u5_u7_n129 ) , .A2( u1_u5_u7_n132 ) , .ZN( u1_u5_u7_n149 ) );
  OAI21_X1 u1_u5_u7_U3 (.ZN( u1_u5_u7_n159 ) , .A( u1_u5_u7_n165 ) , .B2( u1_u5_u7_n171 ) , .B1( u1_u5_u7_n174 ) );
  NAND2_X1 u1_u5_u7_U30 (.A1( u1_u5_u7_n113 ) , .A2( u1_u5_u7_n124 ) , .ZN( u1_u5_u7_n130 ) );
  INV_X1 u1_u5_u7_U31 (.A( u1_u5_u7_n112 ) , .ZN( u1_u5_u7_n173 ) );
  INV_X1 u1_u5_u7_U32 (.A( u1_u5_u7_n128 ) , .ZN( u1_u5_u7_n168 ) );
  INV_X1 u1_u5_u7_U33 (.A( u1_u5_u7_n148 ) , .ZN( u1_u5_u7_n169 ) );
  INV_X1 u1_u5_u7_U34 (.A( u1_u5_u7_n127 ) , .ZN( u1_u5_u7_n179 ) );
  NOR2_X1 u1_u5_u7_U35 (.ZN( u1_u5_u7_n101 ) , .A2( u1_u5_u7_n150 ) , .A1( u1_u5_u7_n156 ) );
  AOI211_X1 u1_u5_u7_U36 (.B( u1_u5_u7_n154 ) , .A( u1_u5_u7_n155 ) , .C1( u1_u5_u7_n156 ) , .ZN( u1_u5_u7_n157 ) , .C2( u1_u5_u7_n172 ) );
  INV_X1 u1_u5_u7_U37 (.A( u1_u5_u7_n153 ) , .ZN( u1_u5_u7_n172 ) );
  AOI211_X1 u1_u5_u7_U38 (.B( u1_u5_u7_n139 ) , .A( u1_u5_u7_n140 ) , .C2( u1_u5_u7_n141 ) , .ZN( u1_u5_u7_n142 ) , .C1( u1_u5_u7_n156 ) );
  NAND4_X1 u1_u5_u7_U39 (.A3( u1_u5_u7_n127 ) , .A2( u1_u5_u7_n128 ) , .A1( u1_u5_u7_n129 ) , .ZN( u1_u5_u7_n141 ) , .A4( u1_u5_u7_n147 ) );
  INV_X1 u1_u5_u7_U4 (.A( u1_u5_u7_n111 ) , .ZN( u1_u5_u7_n170 ) );
  AOI21_X1 u1_u5_u7_U40 (.A( u1_u5_u7_n137 ) , .B1( u1_u5_u7_n138 ) , .ZN( u1_u5_u7_n139 ) , .B2( u1_u5_u7_n146 ) );
  OAI22_X1 u1_u5_u7_U41 (.B1( u1_u5_u7_n136 ) , .ZN( u1_u5_u7_n140 ) , .A1( u1_u5_u7_n153 ) , .B2( u1_u5_u7_n162 ) , .A2( u1_u5_u7_n164 ) );
  AOI21_X1 u1_u5_u7_U42 (.ZN( u1_u5_u7_n123 ) , .B1( u1_u5_u7_n165 ) , .B2( u1_u5_u7_n177 ) , .A( u1_u5_u7_n97 ) );
  AOI21_X1 u1_u5_u7_U43 (.B2( u1_u5_u7_n113 ) , .B1( u1_u5_u7_n124 ) , .A( u1_u5_u7_n125 ) , .ZN( u1_u5_u7_n97 ) );
  INV_X1 u1_u5_u7_U44 (.A( u1_u5_u7_n125 ) , .ZN( u1_u5_u7_n161 ) );
  INV_X1 u1_u5_u7_U45 (.A( u1_u5_u7_n152 ) , .ZN( u1_u5_u7_n162 ) );
  AOI22_X1 u1_u5_u7_U46 (.A2( u1_u5_u7_n114 ) , .ZN( u1_u5_u7_n119 ) , .B1( u1_u5_u7_n130 ) , .A1( u1_u5_u7_n156 ) , .B2( u1_u5_u7_n165 ) );
  NAND2_X1 u1_u5_u7_U47 (.A2( u1_u5_u7_n112 ) , .ZN( u1_u5_u7_n114 ) , .A1( u1_u5_u7_n175 ) );
  AND2_X1 u1_u5_u7_U48 (.ZN( u1_u5_u7_n145 ) , .A2( u1_u5_u7_n98 ) , .A1( u1_u5_u7_n99 ) );
  NOR2_X1 u1_u5_u7_U49 (.ZN( u1_u5_u7_n137 ) , .A1( u1_u5_u7_n150 ) , .A2( u1_u5_u7_n161 ) );
  INV_X1 u1_u5_u7_U5 (.A( u1_u5_u7_n149 ) , .ZN( u1_u5_u7_n175 ) );
  AOI21_X1 u1_u5_u7_U50 (.ZN( u1_u5_u7_n105 ) , .B2( u1_u5_u7_n110 ) , .A( u1_u5_u7_n125 ) , .B1( u1_u5_u7_n147 ) );
  NAND2_X1 u1_u5_u7_U51 (.ZN( u1_u5_u7_n146 ) , .A1( u1_u5_u7_n95 ) , .A2( u1_u5_u7_n98 ) );
  NAND2_X1 u1_u5_u7_U52 (.A2( u1_u5_u7_n103 ) , .ZN( u1_u5_u7_n147 ) , .A1( u1_u5_u7_n93 ) );
  NAND2_X1 u1_u5_u7_U53 (.A1( u1_u5_u7_n103 ) , .ZN( u1_u5_u7_n127 ) , .A2( u1_u5_u7_n99 ) );
  OR2_X1 u1_u5_u7_U54 (.ZN( u1_u5_u7_n126 ) , .A2( u1_u5_u7_n152 ) , .A1( u1_u5_u7_n156 ) );
  NAND2_X1 u1_u5_u7_U55 (.A2( u1_u5_u7_n102 ) , .A1( u1_u5_u7_n103 ) , .ZN( u1_u5_u7_n133 ) );
  NAND2_X1 u1_u5_u7_U56 (.ZN( u1_u5_u7_n112 ) , .A2( u1_u5_u7_n96 ) , .A1( u1_u5_u7_n99 ) );
  NAND2_X1 u1_u5_u7_U57 (.A2( u1_u5_u7_n102 ) , .ZN( u1_u5_u7_n128 ) , .A1( u1_u5_u7_n98 ) );
  NAND2_X1 u1_u5_u7_U58 (.A1( u1_u5_u7_n100 ) , .ZN( u1_u5_u7_n113 ) , .A2( u1_u5_u7_n93 ) );
  NAND2_X1 u1_u5_u7_U59 (.A2( u1_u5_u7_n102 ) , .ZN( u1_u5_u7_n124 ) , .A1( u1_u5_u7_n96 ) );
  INV_X1 u1_u5_u7_U6 (.A( u1_u5_u7_n154 ) , .ZN( u1_u5_u7_n178 ) );
  NAND2_X1 u1_u5_u7_U60 (.ZN( u1_u5_u7_n110 ) , .A1( u1_u5_u7_n95 ) , .A2( u1_u5_u7_n96 ) );
  INV_X1 u1_u5_u7_U61 (.A( u1_u5_u7_n150 ) , .ZN( u1_u5_u7_n164 ) );
  AND2_X1 u1_u5_u7_U62 (.ZN( u1_u5_u7_n134 ) , .A1( u1_u5_u7_n93 ) , .A2( u1_u5_u7_n98 ) );
  NAND2_X1 u1_u5_u7_U63 (.A1( u1_u5_u7_n100 ) , .A2( u1_u5_u7_n102 ) , .ZN( u1_u5_u7_n129 ) );
  NAND2_X1 u1_u5_u7_U64 (.A2( u1_u5_u7_n103 ) , .ZN( u1_u5_u7_n131 ) , .A1( u1_u5_u7_n95 ) );
  NAND2_X1 u1_u5_u7_U65 (.A1( u1_u5_u7_n100 ) , .ZN( u1_u5_u7_n138 ) , .A2( u1_u5_u7_n99 ) );
  NAND2_X1 u1_u5_u7_U66 (.ZN( u1_u5_u7_n132 ) , .A1( u1_u5_u7_n93 ) , .A2( u1_u5_u7_n96 ) );
  NAND2_X1 u1_u5_u7_U67 (.A1( u1_u5_u7_n100 ) , .ZN( u1_u5_u7_n148 ) , .A2( u1_u5_u7_n95 ) );
  NOR2_X1 u1_u5_u7_U68 (.A2( u1_u5_X_47 ) , .ZN( u1_u5_u7_n150 ) , .A1( u1_u5_u7_n163 ) );
  NOR2_X1 u1_u5_u7_U69 (.A2( u1_u5_X_43 ) , .A1( u1_u5_X_44 ) , .ZN( u1_u5_u7_n103 ) );
  AOI211_X1 u1_u5_u7_U7 (.ZN( u1_u5_u7_n116 ) , .A( u1_u5_u7_n155 ) , .C1( u1_u5_u7_n161 ) , .C2( u1_u5_u7_n171 ) , .B( u1_u5_u7_n94 ) );
  NOR2_X1 u1_u5_u7_U70 (.A2( u1_u5_X_48 ) , .A1( u1_u5_u7_n166 ) , .ZN( u1_u5_u7_n95 ) );
  NOR2_X1 u1_u5_u7_U71 (.A2( u1_u5_X_45 ) , .A1( u1_u5_X_48 ) , .ZN( u1_u5_u7_n99 ) );
  NOR2_X1 u1_u5_u7_U72 (.A2( u1_u5_X_44 ) , .A1( u1_u5_u7_n167 ) , .ZN( u1_u5_u7_n98 ) );
  NOR2_X1 u1_u5_u7_U73 (.A2( u1_u5_X_46 ) , .A1( u1_u5_X_47 ) , .ZN( u1_u5_u7_n152 ) );
  AND2_X1 u1_u5_u7_U74 (.A1( u1_u5_X_47 ) , .ZN( u1_u5_u7_n156 ) , .A2( u1_u5_u7_n163 ) );
  NAND2_X1 u1_u5_u7_U75 (.A2( u1_u5_X_46 ) , .A1( u1_u5_X_47 ) , .ZN( u1_u5_u7_n125 ) );
  AND2_X1 u1_u5_u7_U76 (.A2( u1_u5_X_45 ) , .A1( u1_u5_X_48 ) , .ZN( u1_u5_u7_n102 ) );
  AND2_X1 u1_u5_u7_U77 (.A2( u1_u5_X_43 ) , .A1( u1_u5_X_44 ) , .ZN( u1_u5_u7_n96 ) );
  AND2_X1 u1_u5_u7_U78 (.A1( u1_u5_X_44 ) , .ZN( u1_u5_u7_n100 ) , .A2( u1_u5_u7_n167 ) );
  AND2_X1 u1_u5_u7_U79 (.A1( u1_u5_X_48 ) , .A2( u1_u5_u7_n166 ) , .ZN( u1_u5_u7_n93 ) );
  OAI222_X1 u1_u5_u7_U8 (.C2( u1_u5_u7_n101 ) , .B2( u1_u5_u7_n111 ) , .A1( u1_u5_u7_n113 ) , .C1( u1_u5_u7_n146 ) , .A2( u1_u5_u7_n162 ) , .B1( u1_u5_u7_n164 ) , .ZN( u1_u5_u7_n94 ) );
  INV_X1 u1_u5_u7_U80 (.A( u1_u5_X_46 ) , .ZN( u1_u5_u7_n163 ) );
  INV_X1 u1_u5_u7_U81 (.A( u1_u5_X_43 ) , .ZN( u1_u5_u7_n167 ) );
  INV_X1 u1_u5_u7_U82 (.A( u1_u5_X_45 ) , .ZN( u1_u5_u7_n166 ) );
  NAND4_X1 u1_u5_u7_U83 (.ZN( u1_out5_5 ) , .A4( u1_u5_u7_n108 ) , .A3( u1_u5_u7_n109 ) , .A1( u1_u5_u7_n116 ) , .A2( u1_u5_u7_n123 ) );
  AOI22_X1 u1_u5_u7_U84 (.ZN( u1_u5_u7_n109 ) , .A2( u1_u5_u7_n126 ) , .B2( u1_u5_u7_n145 ) , .B1( u1_u5_u7_n156 ) , .A1( u1_u5_u7_n171 ) );
  NOR4_X1 u1_u5_u7_U85 (.A4( u1_u5_u7_n104 ) , .A3( u1_u5_u7_n105 ) , .A2( u1_u5_u7_n106 ) , .A1( u1_u5_u7_n107 ) , .ZN( u1_u5_u7_n108 ) );
  NAND4_X1 u1_u5_u7_U86 (.ZN( u1_out5_27 ) , .A4( u1_u5_u7_n118 ) , .A3( u1_u5_u7_n119 ) , .A2( u1_u5_u7_n120 ) , .A1( u1_u5_u7_n121 ) );
  OAI21_X1 u1_u5_u7_U87 (.ZN( u1_u5_u7_n121 ) , .B2( u1_u5_u7_n145 ) , .A( u1_u5_u7_n150 ) , .B1( u1_u5_u7_n174 ) );
  OAI21_X1 u1_u5_u7_U88 (.ZN( u1_u5_u7_n120 ) , .A( u1_u5_u7_n161 ) , .B2( u1_u5_u7_n170 ) , .B1( u1_u5_u7_n179 ) );
  NAND4_X1 u1_u5_u7_U89 (.ZN( u1_out5_21 ) , .A4( u1_u5_u7_n157 ) , .A3( u1_u5_u7_n158 ) , .A2( u1_u5_u7_n159 ) , .A1( u1_u5_u7_n160 ) );
  OAI221_X1 u1_u5_u7_U9 (.C1( u1_u5_u7_n101 ) , .C2( u1_u5_u7_n147 ) , .ZN( u1_u5_u7_n155 ) , .B2( u1_u5_u7_n162 ) , .A( u1_u5_u7_n91 ) , .B1( u1_u5_u7_n92 ) );
  OAI21_X1 u1_u5_u7_U90 (.B1( u1_u5_u7_n145 ) , .ZN( u1_u5_u7_n160 ) , .A( u1_u5_u7_n161 ) , .B2( u1_u5_u7_n177 ) );
  AOI22_X1 u1_u5_u7_U91 (.B2( u1_u5_u7_n149 ) , .B1( u1_u5_u7_n150 ) , .A2( u1_u5_u7_n151 ) , .A1( u1_u5_u7_n152 ) , .ZN( u1_u5_u7_n158 ) );
  NAND4_X1 u1_u5_u7_U92 (.ZN( u1_out5_15 ) , .A4( u1_u5_u7_n142 ) , .A3( u1_u5_u7_n143 ) , .A2( u1_u5_u7_n144 ) , .A1( u1_u5_u7_n178 ) );
  OR2_X1 u1_u5_u7_U93 (.A2( u1_u5_u7_n125 ) , .A1( u1_u5_u7_n129 ) , .ZN( u1_u5_u7_n144 ) );
  AOI22_X1 u1_u5_u7_U94 (.A2( u1_u5_u7_n126 ) , .ZN( u1_u5_u7_n143 ) , .B2( u1_u5_u7_n165 ) , .B1( u1_u5_u7_n173 ) , .A1( u1_u5_u7_n174 ) );
  NAND3_X1 u1_u5_u7_U95 (.A3( u1_u5_u7_n146 ) , .A2( u1_u5_u7_n147 ) , .A1( u1_u5_u7_n148 ) , .ZN( u1_u5_u7_n151 ) );
  NAND3_X1 u1_u5_u7_U96 (.A3( u1_u5_u7_n131 ) , .A2( u1_u5_u7_n132 ) , .A1( u1_u5_u7_n133 ) , .ZN( u1_u5_u7_n135 ) );
  XOR2_X1 u1_u7_U10 (.B( u1_K8_45 ) , .A( u1_R6_30 ) , .Z( u1_u7_X_45 ) );
  XOR2_X1 u1_u7_U9 (.B( u1_K8_46 ) , .A( u1_R6_31 ) , .Z( u1_u7_X_46 ) );
  OAI221_X1 u1_u7_u7_U10 (.C1( u1_u7_u7_n101 ) , .C2( u1_u7_u7_n147 ) , .ZN( u1_u7_u7_n155 ) , .B2( u1_u7_u7_n162 ) , .A( u1_u7_u7_n91 ) , .B1( u1_u7_u7_n92 ) );
  AND3_X1 u1_u7_u7_U11 (.A3( u1_u7_u7_n110 ) , .A2( u1_u7_u7_n127 ) , .A1( u1_u7_u7_n132 ) , .ZN( u1_u7_u7_n92 ) );
  OAI21_X1 u1_u7_u7_U12 (.A( u1_u7_u7_n161 ) , .B1( u1_u7_u7_n168 ) , .B2( u1_u7_u7_n173 ) , .ZN( u1_u7_u7_n91 ) );
  AOI211_X1 u1_u7_u7_U13 (.A( u1_u7_u7_n117 ) , .ZN( u1_u7_u7_n118 ) , .C2( u1_u7_u7_n126 ) , .C1( u1_u7_u7_n177 ) , .B( u1_u7_u7_n180 ) );
  OAI22_X1 u1_u7_u7_U14 (.B1( u1_u7_u7_n115 ) , .ZN( u1_u7_u7_n117 ) , .A2( u1_u7_u7_n133 ) , .A1( u1_u7_u7_n137 ) , .B2( u1_u7_u7_n162 ) );
  INV_X1 u1_u7_u7_U15 (.A( u1_u7_u7_n116 ) , .ZN( u1_u7_u7_n180 ) );
  NOR3_X1 u1_u7_u7_U16 (.ZN( u1_u7_u7_n115 ) , .A3( u1_u7_u7_n145 ) , .A2( u1_u7_u7_n168 ) , .A1( u1_u7_u7_n169 ) );
  NOR3_X1 u1_u7_u7_U17 (.A2( u1_u7_u7_n134 ) , .A1( u1_u7_u7_n135 ) , .ZN( u1_u7_u7_n136 ) , .A3( u1_u7_u7_n171 ) );
  NOR2_X1 u1_u7_u7_U18 (.A1( u1_u7_u7_n130 ) , .A2( u1_u7_u7_n134 ) , .ZN( u1_u7_u7_n153 ) );
  NOR2_X1 u1_u7_u7_U19 (.ZN( u1_u7_u7_n111 ) , .A2( u1_u7_u7_n134 ) , .A1( u1_u7_u7_n169 ) );
  AOI21_X1 u1_u7_u7_U20 (.ZN( u1_u7_u7_n104 ) , .B2( u1_u7_u7_n112 ) , .B1( u1_u7_u7_n127 ) , .A( u1_u7_u7_n164 ) );
  AOI21_X1 u1_u7_u7_U21 (.ZN( u1_u7_u7_n106 ) , .B1( u1_u7_u7_n133 ) , .B2( u1_u7_u7_n146 ) , .A( u1_u7_u7_n162 ) );
  AOI21_X1 u1_u7_u7_U22 (.A( u1_u7_u7_n101 ) , .ZN( u1_u7_u7_n107 ) , .B2( u1_u7_u7_n128 ) , .B1( u1_u7_u7_n175 ) );
  INV_X1 u1_u7_u7_U23 (.A( u1_u7_u7_n101 ) , .ZN( u1_u7_u7_n165 ) );
  INV_X1 u1_u7_u7_U24 (.A( u1_u7_u7_n138 ) , .ZN( u1_u7_u7_n171 ) );
  INV_X1 u1_u7_u7_U25 (.A( u1_u7_u7_n131 ) , .ZN( u1_u7_u7_n177 ) );
  INV_X1 u1_u7_u7_U26 (.A( u1_u7_u7_n110 ) , .ZN( u1_u7_u7_n174 ) );
  NAND2_X1 u1_u7_u7_U27 (.A1( u1_u7_u7_n129 ) , .A2( u1_u7_u7_n132 ) , .ZN( u1_u7_u7_n149 ) );
  NAND2_X1 u1_u7_u7_U28 (.A1( u1_u7_u7_n113 ) , .A2( u1_u7_u7_n124 ) , .ZN( u1_u7_u7_n130 ) );
  INV_X1 u1_u7_u7_U29 (.A( u1_u7_u7_n128 ) , .ZN( u1_u7_u7_n168 ) );
  OAI21_X1 u1_u7_u7_U3 (.ZN( u1_u7_u7_n159 ) , .A( u1_u7_u7_n165 ) , .B2( u1_u7_u7_n171 ) , .B1( u1_u7_u7_n174 ) );
  INV_X1 u1_u7_u7_U30 (.A( u1_u7_u7_n148 ) , .ZN( u1_u7_u7_n169 ) );
  INV_X1 u1_u7_u7_U31 (.A( u1_u7_u7_n112 ) , .ZN( u1_u7_u7_n173 ) );
  INV_X1 u1_u7_u7_U32 (.A( u1_u7_u7_n127 ) , .ZN( u1_u7_u7_n179 ) );
  NOR2_X1 u1_u7_u7_U33 (.ZN( u1_u7_u7_n101 ) , .A2( u1_u7_u7_n150 ) , .A1( u1_u7_u7_n156 ) );
  AOI211_X1 u1_u7_u7_U34 (.B( u1_u7_u7_n154 ) , .A( u1_u7_u7_n155 ) , .C1( u1_u7_u7_n156 ) , .ZN( u1_u7_u7_n157 ) , .C2( u1_u7_u7_n172 ) );
  INV_X1 u1_u7_u7_U35 (.A( u1_u7_u7_n153 ) , .ZN( u1_u7_u7_n172 ) );
  AOI211_X1 u1_u7_u7_U36 (.B( u1_u7_u7_n139 ) , .A( u1_u7_u7_n140 ) , .C2( u1_u7_u7_n141 ) , .ZN( u1_u7_u7_n142 ) , .C1( u1_u7_u7_n156 ) );
  NAND4_X1 u1_u7_u7_U37 (.A3( u1_u7_u7_n127 ) , .A2( u1_u7_u7_n128 ) , .A1( u1_u7_u7_n129 ) , .ZN( u1_u7_u7_n141 ) , .A4( u1_u7_u7_n147 ) );
  AOI21_X1 u1_u7_u7_U38 (.A( u1_u7_u7_n137 ) , .B1( u1_u7_u7_n138 ) , .ZN( u1_u7_u7_n139 ) , .B2( u1_u7_u7_n146 ) );
  OAI22_X1 u1_u7_u7_U39 (.B1( u1_u7_u7_n136 ) , .ZN( u1_u7_u7_n140 ) , .A1( u1_u7_u7_n153 ) , .B2( u1_u7_u7_n162 ) , .A2( u1_u7_u7_n164 ) );
  INV_X1 u1_u7_u7_U4 (.A( u1_u7_u7_n149 ) , .ZN( u1_u7_u7_n175 ) );
  INV_X1 u1_u7_u7_U40 (.A( u1_u7_u7_n125 ) , .ZN( u1_u7_u7_n161 ) );
  AOI21_X1 u1_u7_u7_U41 (.ZN( u1_u7_u7_n123 ) , .B1( u1_u7_u7_n165 ) , .B2( u1_u7_u7_n177 ) , .A( u1_u7_u7_n97 ) );
  AOI21_X1 u1_u7_u7_U42 (.B2( u1_u7_u7_n113 ) , .B1( u1_u7_u7_n124 ) , .A( u1_u7_u7_n125 ) , .ZN( u1_u7_u7_n97 ) );
  INV_X1 u1_u7_u7_U43 (.A( u1_u7_u7_n152 ) , .ZN( u1_u7_u7_n162 ) );
  AOI22_X1 u1_u7_u7_U44 (.A2( u1_u7_u7_n114 ) , .ZN( u1_u7_u7_n119 ) , .B1( u1_u7_u7_n130 ) , .A1( u1_u7_u7_n156 ) , .B2( u1_u7_u7_n165 ) );
  NAND2_X1 u1_u7_u7_U45 (.A2( u1_u7_u7_n112 ) , .ZN( u1_u7_u7_n114 ) , .A1( u1_u7_u7_n175 ) );
  NOR2_X1 u1_u7_u7_U46 (.ZN( u1_u7_u7_n137 ) , .A1( u1_u7_u7_n150 ) , .A2( u1_u7_u7_n161 ) );
  AND2_X1 u1_u7_u7_U47 (.ZN( u1_u7_u7_n145 ) , .A2( u1_u7_u7_n98 ) , .A1( u1_u7_u7_n99 ) );
  AOI21_X1 u1_u7_u7_U48 (.ZN( u1_u7_u7_n105 ) , .B2( u1_u7_u7_n110 ) , .A( u1_u7_u7_n125 ) , .B1( u1_u7_u7_n147 ) );
  NAND2_X1 u1_u7_u7_U49 (.ZN( u1_u7_u7_n146 ) , .A1( u1_u7_u7_n95 ) , .A2( u1_u7_u7_n98 ) );
  INV_X1 u1_u7_u7_U5 (.A( u1_u7_u7_n154 ) , .ZN( u1_u7_u7_n178 ) );
  NAND2_X1 u1_u7_u7_U50 (.A2( u1_u7_u7_n103 ) , .ZN( u1_u7_u7_n147 ) , .A1( u1_u7_u7_n93 ) );
  NAND2_X1 u1_u7_u7_U51 (.A1( u1_u7_u7_n103 ) , .ZN( u1_u7_u7_n127 ) , .A2( u1_u7_u7_n99 ) );
  NAND2_X1 u1_u7_u7_U52 (.A2( u1_u7_u7_n102 ) , .A1( u1_u7_u7_n103 ) , .ZN( u1_u7_u7_n133 ) );
  OR2_X1 u1_u7_u7_U53 (.ZN( u1_u7_u7_n126 ) , .A2( u1_u7_u7_n152 ) , .A1( u1_u7_u7_n156 ) );
  NAND2_X1 u1_u7_u7_U54 (.ZN( u1_u7_u7_n112 ) , .A2( u1_u7_u7_n96 ) , .A1( u1_u7_u7_n99 ) );
  NAND2_X1 u1_u7_u7_U55 (.A2( u1_u7_u7_n102 ) , .ZN( u1_u7_u7_n128 ) , .A1( u1_u7_u7_n98 ) );
  INV_X1 u1_u7_u7_U56 (.A( u1_u7_u7_n150 ) , .ZN( u1_u7_u7_n164 ) );
  AND2_X1 u1_u7_u7_U57 (.ZN( u1_u7_u7_n134 ) , .A1( u1_u7_u7_n93 ) , .A2( u1_u7_u7_n98 ) );
  NAND2_X1 u1_u7_u7_U58 (.ZN( u1_u7_u7_n110 ) , .A1( u1_u7_u7_n95 ) , .A2( u1_u7_u7_n96 ) );
  NAND2_X1 u1_u7_u7_U59 (.A2( u1_u7_u7_n102 ) , .ZN( u1_u7_u7_n124 ) , .A1( u1_u7_u7_n96 ) );
  INV_X1 u1_u7_u7_U6 (.A( u1_u7_u7_n111 ) , .ZN( u1_u7_u7_n170 ) );
  NAND2_X1 u1_u7_u7_U60 (.ZN( u1_u7_u7_n132 ) , .A1( u1_u7_u7_n93 ) , .A2( u1_u7_u7_n96 ) );
  NAND2_X1 u1_u7_u7_U61 (.A2( u1_u7_u7_n103 ) , .ZN( u1_u7_u7_n131 ) , .A1( u1_u7_u7_n95 ) );
  NOR2_X1 u1_u7_u7_U62 (.A2( u1_u7_X_47 ) , .ZN( u1_u7_u7_n150 ) , .A1( u1_u7_u7_n163 ) );
  NOR2_X1 u1_u7_u7_U63 (.A2( u1_u7_X_43 ) , .A1( u1_u7_X_44 ) , .ZN( u1_u7_u7_n103 ) );
  NOR2_X1 u1_u7_u7_U64 (.A2( u1_u7_X_48 ) , .A1( u1_u7_u7_n166 ) , .ZN( u1_u7_u7_n95 ) );
  NOR2_X1 u1_u7_u7_U65 (.A2( u1_u7_X_44 ) , .A1( u1_u7_u7_n167 ) , .ZN( u1_u7_u7_n98 ) );
  NOR2_X1 u1_u7_u7_U66 (.A2( u1_u7_X_45 ) , .A1( u1_u7_X_48 ) , .ZN( u1_u7_u7_n99 ) );
  NOR2_X1 u1_u7_u7_U67 (.A2( u1_u7_X_46 ) , .A1( u1_u7_X_47 ) , .ZN( u1_u7_u7_n152 ) );
  AND2_X1 u1_u7_u7_U68 (.A1( u1_u7_X_47 ) , .ZN( u1_u7_u7_n156 ) , .A2( u1_u7_u7_n163 ) );
  NAND2_X1 u1_u7_u7_U69 (.A2( u1_u7_X_46 ) , .A1( u1_u7_X_47 ) , .ZN( u1_u7_u7_n125 ) );
  AOI211_X1 u1_u7_u7_U7 (.ZN( u1_u7_u7_n116 ) , .A( u1_u7_u7_n155 ) , .C1( u1_u7_u7_n161 ) , .C2( u1_u7_u7_n171 ) , .B( u1_u7_u7_n94 ) );
  AND2_X1 u1_u7_u7_U70 (.A2( u1_u7_X_43 ) , .A1( u1_u7_X_44 ) , .ZN( u1_u7_u7_n96 ) );
  AND2_X1 u1_u7_u7_U71 (.A2( u1_u7_X_45 ) , .A1( u1_u7_X_48 ) , .ZN( u1_u7_u7_n102 ) );
  AND2_X1 u1_u7_u7_U72 (.A1( u1_u7_X_48 ) , .A2( u1_u7_u7_n166 ) , .ZN( u1_u7_u7_n93 ) );
  INV_X1 u1_u7_u7_U73 (.A( u1_u7_X_46 ) , .ZN( u1_u7_u7_n163 ) );
  AND2_X1 u1_u7_u7_U74 (.A1( u1_u7_X_44 ) , .ZN( u1_u7_u7_n100 ) , .A2( u1_u7_u7_n167 ) );
  INV_X1 u1_u7_u7_U75 (.A( u1_u7_X_45 ) , .ZN( u1_u7_u7_n166 ) );
  INV_X1 u1_u7_u7_U76 (.A( u1_u7_X_43 ) , .ZN( u1_u7_u7_n167 ) );
  NAND4_X1 u1_u7_u7_U77 (.ZN( u1_out7_5 ) , .A4( u1_u7_u7_n108 ) , .A3( u1_u7_u7_n109 ) , .A1( u1_u7_u7_n116 ) , .A2( u1_u7_u7_n123 ) );
  AOI22_X1 u1_u7_u7_U78 (.ZN( u1_u7_u7_n109 ) , .A2( u1_u7_u7_n126 ) , .B2( u1_u7_u7_n145 ) , .B1( u1_u7_u7_n156 ) , .A1( u1_u7_u7_n171 ) );
  NOR4_X1 u1_u7_u7_U79 (.A4( u1_u7_u7_n104 ) , .A3( u1_u7_u7_n105 ) , .A2( u1_u7_u7_n106 ) , .A1( u1_u7_u7_n107 ) , .ZN( u1_u7_u7_n108 ) );
  OAI222_X1 u1_u7_u7_U8 (.C2( u1_u7_u7_n101 ) , .B2( u1_u7_u7_n111 ) , .A1( u1_u7_u7_n113 ) , .C1( u1_u7_u7_n146 ) , .A2( u1_u7_u7_n162 ) , .B1( u1_u7_u7_n164 ) , .ZN( u1_u7_u7_n94 ) );
  NAND4_X1 u1_u7_u7_U80 (.ZN( u1_out7_27 ) , .A4( u1_u7_u7_n118 ) , .A3( u1_u7_u7_n119 ) , .A2( u1_u7_u7_n120 ) , .A1( u1_u7_u7_n121 ) );
  OAI21_X1 u1_u7_u7_U81 (.ZN( u1_u7_u7_n121 ) , .B2( u1_u7_u7_n145 ) , .A( u1_u7_u7_n150 ) , .B1( u1_u7_u7_n174 ) );
  OAI21_X1 u1_u7_u7_U82 (.ZN( u1_u7_u7_n120 ) , .A( u1_u7_u7_n161 ) , .B2( u1_u7_u7_n170 ) , .B1( u1_u7_u7_n179 ) );
  NAND4_X1 u1_u7_u7_U83 (.ZN( u1_out7_21 ) , .A4( u1_u7_u7_n157 ) , .A3( u1_u7_u7_n158 ) , .A2( u1_u7_u7_n159 ) , .A1( u1_u7_u7_n160 ) );
  OAI21_X1 u1_u7_u7_U84 (.B1( u1_u7_u7_n145 ) , .ZN( u1_u7_u7_n160 ) , .A( u1_u7_u7_n161 ) , .B2( u1_u7_u7_n177 ) );
  AOI22_X1 u1_u7_u7_U85 (.B2( u1_u7_u7_n149 ) , .B1( u1_u7_u7_n150 ) , .A2( u1_u7_u7_n151 ) , .A1( u1_u7_u7_n152 ) , .ZN( u1_u7_u7_n158 ) );
  NAND4_X1 u1_u7_u7_U86 (.ZN( u1_out7_15 ) , .A4( u1_u7_u7_n142 ) , .A3( u1_u7_u7_n143 ) , .A2( u1_u7_u7_n144 ) , .A1( u1_u7_u7_n178 ) );
  OR2_X1 u1_u7_u7_U87 (.A2( u1_u7_u7_n125 ) , .A1( u1_u7_u7_n129 ) , .ZN( u1_u7_u7_n144 ) );
  AOI22_X1 u1_u7_u7_U88 (.A2( u1_u7_u7_n126 ) , .ZN( u1_u7_u7_n143 ) , .B2( u1_u7_u7_n165 ) , .B1( u1_u7_u7_n173 ) , .A1( u1_u7_u7_n174 ) );
  NAND2_X1 u1_u7_u7_U89 (.A1( u1_u7_u7_n100 ) , .ZN( u1_u7_u7_n148 ) , .A2( u1_u7_u7_n95 ) );
  INV_X1 u1_u7_u7_U9 (.A( u1_u7_u7_n133 ) , .ZN( u1_u7_u7_n176 ) );
  NAND2_X1 u1_u7_u7_U90 (.A1( u1_u7_u7_n100 ) , .ZN( u1_u7_u7_n113 ) , .A2( u1_u7_u7_n93 ) );
  NAND2_X1 u1_u7_u7_U91 (.A1( u1_u7_u7_n100 ) , .ZN( u1_u7_u7_n138 ) , .A2( u1_u7_u7_n99 ) );
  NAND2_X1 u1_u7_u7_U92 (.A1( u1_u7_u7_n100 ) , .A2( u1_u7_u7_n102 ) , .ZN( u1_u7_u7_n129 ) );
  OAI211_X1 u1_u7_u7_U93 (.B( u1_u7_u7_n122 ) , .A( u1_u7_u7_n123 ) , .C2( u1_u7_u7_n124 ) , .ZN( u1_u7_u7_n154 ) , .C1( u1_u7_u7_n162 ) );
  AOI222_X1 u1_u7_u7_U94 (.ZN( u1_u7_u7_n122 ) , .C2( u1_u7_u7_n126 ) , .C1( u1_u7_u7_n145 ) , .B1( u1_u7_u7_n161 ) , .A2( u1_u7_u7_n165 ) , .B2( u1_u7_u7_n170 ) , .A1( u1_u7_u7_n176 ) );
  NAND3_X1 u1_u7_u7_U95 (.A3( u1_u7_u7_n146 ) , .A2( u1_u7_u7_n147 ) , .A1( u1_u7_u7_n148 ) , .ZN( u1_u7_u7_n151 ) );
  NAND3_X1 u1_u7_u7_U96 (.A3( u1_u7_u7_n131 ) , .A2( u1_u7_u7_n132 ) , .A1( u1_u7_u7_n133 ) , .ZN( u1_u7_u7_n135 ) );
  XOR2_X1 u1_u8_U1 (.B( u1_K9_9 ) , .A( u1_R7_6 ) , .Z( u1_u8_X_9 ) );
  XOR2_X1 u1_u8_U47 (.B( u1_K9_11 ) , .A( u1_R7_8 ) , .Z( u1_u8_X_11 ) );
  XOR2_X1 u1_u8_U48 (.B( u1_K9_10 ) , .A( u1_R7_7 ) , .Z( u1_u8_X_10 ) );
  AOI21_X1 u1_u8_u1_U10 (.B2( u1_u8_u1_n155 ) , .B1( u1_u8_u1_n156 ) , .ZN( u1_u8_u1_n157 ) , .A( u1_u8_u1_n174 ) );
  NAND3_X1 u1_u8_u1_U100 (.ZN( u1_u8_u1_n113 ) , .A1( u1_u8_u1_n120 ) , .A3( u1_u8_u1_n133 ) , .A2( u1_u8_u1_n155 ) );
  NAND2_X1 u1_u8_u1_U11 (.ZN( u1_u8_u1_n140 ) , .A2( u1_u8_u1_n150 ) , .A1( u1_u8_u1_n155 ) );
  NAND2_X1 u1_u8_u1_U12 (.A1( u1_u8_u1_n131 ) , .ZN( u1_u8_u1_n147 ) , .A2( u1_u8_u1_n153 ) );
  AOI22_X1 u1_u8_u1_U13 (.B2( u1_u8_u1_n136 ) , .A2( u1_u8_u1_n137 ) , .ZN( u1_u8_u1_n143 ) , .A1( u1_u8_u1_n171 ) , .B1( u1_u8_u1_n173 ) );
  INV_X1 u1_u8_u1_U14 (.A( u1_u8_u1_n147 ) , .ZN( u1_u8_u1_n181 ) );
  INV_X1 u1_u8_u1_U15 (.A( u1_u8_u1_n139 ) , .ZN( u1_u8_u1_n174 ) );
  INV_X1 u1_u8_u1_U16 (.A( u1_u8_u1_n112 ) , .ZN( u1_u8_u1_n171 ) );
  NAND2_X1 u1_u8_u1_U17 (.ZN( u1_u8_u1_n141 ) , .A1( u1_u8_u1_n153 ) , .A2( u1_u8_u1_n156 ) );
  AND2_X1 u1_u8_u1_U18 (.A1( u1_u8_u1_n123 ) , .ZN( u1_u8_u1_n134 ) , .A2( u1_u8_u1_n161 ) );
  NAND2_X1 u1_u8_u1_U19 (.A2( u1_u8_u1_n115 ) , .A1( u1_u8_u1_n116 ) , .ZN( u1_u8_u1_n148 ) );
  NAND2_X1 u1_u8_u1_U20 (.A2( u1_u8_u1_n133 ) , .A1( u1_u8_u1_n135 ) , .ZN( u1_u8_u1_n159 ) );
  NAND2_X1 u1_u8_u1_U21 (.A2( u1_u8_u1_n115 ) , .A1( u1_u8_u1_n120 ) , .ZN( u1_u8_u1_n132 ) );
  INV_X1 u1_u8_u1_U22 (.A( u1_u8_u1_n154 ) , .ZN( u1_u8_u1_n178 ) );
  INV_X1 u1_u8_u1_U23 (.A( u1_u8_u1_n151 ) , .ZN( u1_u8_u1_n183 ) );
  AND2_X1 u1_u8_u1_U24 (.A1( u1_u8_u1_n129 ) , .A2( u1_u8_u1_n133 ) , .ZN( u1_u8_u1_n149 ) );
  INV_X1 u1_u8_u1_U25 (.A( u1_u8_u1_n131 ) , .ZN( u1_u8_u1_n180 ) );
  OR4_X1 u1_u8_u1_U26 (.A4( u1_u8_u1_n106 ) , .A3( u1_u8_u1_n107 ) , .ZN( u1_u8_u1_n108 ) , .A1( u1_u8_u1_n117 ) , .A2( u1_u8_u1_n184 ) );
  AOI21_X1 u1_u8_u1_U27 (.ZN( u1_u8_u1_n106 ) , .A( u1_u8_u1_n112 ) , .B1( u1_u8_u1_n154 ) , .B2( u1_u8_u1_n156 ) );
  AOI21_X1 u1_u8_u1_U28 (.ZN( u1_u8_u1_n107 ) , .B1( u1_u8_u1_n134 ) , .B2( u1_u8_u1_n149 ) , .A( u1_u8_u1_n174 ) );
  INV_X1 u1_u8_u1_U29 (.A( u1_u8_u1_n101 ) , .ZN( u1_u8_u1_n184 ) );
  INV_X1 u1_u8_u1_U3 (.A( u1_u8_u1_n159 ) , .ZN( u1_u8_u1_n182 ) );
  AOI221_X1 u1_u8_u1_U30 (.B1( u1_u8_u1_n140 ) , .ZN( u1_u8_u1_n167 ) , .B2( u1_u8_u1_n172 ) , .C2( u1_u8_u1_n175 ) , .C1( u1_u8_u1_n178 ) , .A( u1_u8_u1_n188 ) );
  INV_X1 u1_u8_u1_U31 (.ZN( u1_u8_u1_n188 ) , .A( u1_u8_u1_n97 ) );
  AOI211_X1 u1_u8_u1_U32 (.A( u1_u8_u1_n118 ) , .C1( u1_u8_u1_n132 ) , .C2( u1_u8_u1_n139 ) , .B( u1_u8_u1_n96 ) , .ZN( u1_u8_u1_n97 ) );
  AOI21_X1 u1_u8_u1_U33 (.B2( u1_u8_u1_n121 ) , .B1( u1_u8_u1_n135 ) , .A( u1_u8_u1_n152 ) , .ZN( u1_u8_u1_n96 ) );
  OAI221_X1 u1_u8_u1_U34 (.A( u1_u8_u1_n119 ) , .C2( u1_u8_u1_n129 ) , .ZN( u1_u8_u1_n138 ) , .B2( u1_u8_u1_n152 ) , .C1( u1_u8_u1_n174 ) , .B1( u1_u8_u1_n187 ) );
  INV_X1 u1_u8_u1_U35 (.A( u1_u8_u1_n148 ) , .ZN( u1_u8_u1_n187 ) );
  AOI211_X1 u1_u8_u1_U36 (.B( u1_u8_u1_n117 ) , .A( u1_u8_u1_n118 ) , .ZN( u1_u8_u1_n119 ) , .C2( u1_u8_u1_n146 ) , .C1( u1_u8_u1_n159 ) );
  NOR2_X1 u1_u8_u1_U37 (.A1( u1_u8_u1_n168 ) , .A2( u1_u8_u1_n176 ) , .ZN( u1_u8_u1_n98 ) );
  AOI211_X1 u1_u8_u1_U38 (.B( u1_u8_u1_n162 ) , .A( u1_u8_u1_n163 ) , .C2( u1_u8_u1_n164 ) , .ZN( u1_u8_u1_n165 ) , .C1( u1_u8_u1_n171 ) );
  AOI21_X1 u1_u8_u1_U39 (.A( u1_u8_u1_n160 ) , .B2( u1_u8_u1_n161 ) , .ZN( u1_u8_u1_n162 ) , .B1( u1_u8_u1_n182 ) );
  AOI221_X1 u1_u8_u1_U4 (.A( u1_u8_u1_n138 ) , .C2( u1_u8_u1_n139 ) , .C1( u1_u8_u1_n140 ) , .B2( u1_u8_u1_n141 ) , .ZN( u1_u8_u1_n142 ) , .B1( u1_u8_u1_n175 ) );
  OR2_X1 u1_u8_u1_U40 (.A2( u1_u8_u1_n157 ) , .A1( u1_u8_u1_n158 ) , .ZN( u1_u8_u1_n163 ) );
  NAND2_X1 u1_u8_u1_U41 (.A1( u1_u8_u1_n128 ) , .ZN( u1_u8_u1_n146 ) , .A2( u1_u8_u1_n160 ) );
  NAND2_X1 u1_u8_u1_U42 (.A2( u1_u8_u1_n112 ) , .ZN( u1_u8_u1_n139 ) , .A1( u1_u8_u1_n152 ) );
  NAND2_X1 u1_u8_u1_U43 (.A1( u1_u8_u1_n105 ) , .ZN( u1_u8_u1_n156 ) , .A2( u1_u8_u1_n99 ) );
  NOR2_X1 u1_u8_u1_U44 (.ZN( u1_u8_u1_n117 ) , .A1( u1_u8_u1_n121 ) , .A2( u1_u8_u1_n160 ) );
  OAI21_X1 u1_u8_u1_U45 (.B2( u1_u8_u1_n123 ) , .ZN( u1_u8_u1_n145 ) , .B1( u1_u8_u1_n160 ) , .A( u1_u8_u1_n185 ) );
  INV_X1 u1_u8_u1_U46 (.A( u1_u8_u1_n122 ) , .ZN( u1_u8_u1_n185 ) );
  AOI21_X1 u1_u8_u1_U47 (.B2( u1_u8_u1_n120 ) , .B1( u1_u8_u1_n121 ) , .ZN( u1_u8_u1_n122 ) , .A( u1_u8_u1_n128 ) );
  AOI21_X1 u1_u8_u1_U48 (.A( u1_u8_u1_n128 ) , .B2( u1_u8_u1_n129 ) , .ZN( u1_u8_u1_n130 ) , .B1( u1_u8_u1_n150 ) );
  NAND2_X1 u1_u8_u1_U49 (.ZN( u1_u8_u1_n112 ) , .A1( u1_u8_u1_n169 ) , .A2( u1_u8_u1_n170 ) );
  AOI211_X1 u1_u8_u1_U5 (.ZN( u1_u8_u1_n124 ) , .A( u1_u8_u1_n138 ) , .C2( u1_u8_u1_n139 ) , .B( u1_u8_u1_n145 ) , .C1( u1_u8_u1_n147 ) );
  NAND2_X1 u1_u8_u1_U50 (.ZN( u1_u8_u1_n129 ) , .A2( u1_u8_u1_n95 ) , .A1( u1_u8_u1_n98 ) );
  NAND2_X1 u1_u8_u1_U51 (.A1( u1_u8_u1_n102 ) , .ZN( u1_u8_u1_n154 ) , .A2( u1_u8_u1_n99 ) );
  NAND2_X1 u1_u8_u1_U52 (.A2( u1_u8_u1_n100 ) , .ZN( u1_u8_u1_n135 ) , .A1( u1_u8_u1_n99 ) );
  AOI21_X1 u1_u8_u1_U53 (.A( u1_u8_u1_n152 ) , .B2( u1_u8_u1_n153 ) , .B1( u1_u8_u1_n154 ) , .ZN( u1_u8_u1_n158 ) );
  INV_X1 u1_u8_u1_U54 (.A( u1_u8_u1_n160 ) , .ZN( u1_u8_u1_n175 ) );
  NAND2_X1 u1_u8_u1_U55 (.A1( u1_u8_u1_n100 ) , .ZN( u1_u8_u1_n116 ) , .A2( u1_u8_u1_n95 ) );
  NAND2_X1 u1_u8_u1_U56 (.A1( u1_u8_u1_n102 ) , .ZN( u1_u8_u1_n131 ) , .A2( u1_u8_u1_n95 ) );
  NAND2_X1 u1_u8_u1_U57 (.A2( u1_u8_u1_n104 ) , .ZN( u1_u8_u1_n121 ) , .A1( u1_u8_u1_n98 ) );
  NAND2_X1 u1_u8_u1_U58 (.A1( u1_u8_u1_n103 ) , .ZN( u1_u8_u1_n153 ) , .A2( u1_u8_u1_n98 ) );
  NAND2_X1 u1_u8_u1_U59 (.A2( u1_u8_u1_n104 ) , .A1( u1_u8_u1_n105 ) , .ZN( u1_u8_u1_n133 ) );
  AOI22_X1 u1_u8_u1_U6 (.B2( u1_u8_u1_n113 ) , .A2( u1_u8_u1_n114 ) , .ZN( u1_u8_u1_n125 ) , .A1( u1_u8_u1_n171 ) , .B1( u1_u8_u1_n173 ) );
  NAND2_X1 u1_u8_u1_U60 (.ZN( u1_u8_u1_n150 ) , .A2( u1_u8_u1_n98 ) , .A1( u1_u8_u1_n99 ) );
  NAND2_X1 u1_u8_u1_U61 (.A1( u1_u8_u1_n105 ) , .ZN( u1_u8_u1_n155 ) , .A2( u1_u8_u1_n95 ) );
  OAI21_X1 u1_u8_u1_U62 (.ZN( u1_u8_u1_n109 ) , .B1( u1_u8_u1_n129 ) , .B2( u1_u8_u1_n160 ) , .A( u1_u8_u1_n167 ) );
  NAND2_X1 u1_u8_u1_U63 (.A2( u1_u8_u1_n100 ) , .A1( u1_u8_u1_n103 ) , .ZN( u1_u8_u1_n120 ) );
  NAND2_X1 u1_u8_u1_U64 (.A1( u1_u8_u1_n102 ) , .A2( u1_u8_u1_n104 ) , .ZN( u1_u8_u1_n115 ) );
  NAND2_X1 u1_u8_u1_U65 (.A2( u1_u8_u1_n100 ) , .A1( u1_u8_u1_n104 ) , .ZN( u1_u8_u1_n151 ) );
  NAND2_X1 u1_u8_u1_U66 (.A2( u1_u8_u1_n103 ) , .A1( u1_u8_u1_n105 ) , .ZN( u1_u8_u1_n161 ) );
  INV_X1 u1_u8_u1_U67 (.A( u1_u8_u1_n152 ) , .ZN( u1_u8_u1_n173 ) );
  INV_X1 u1_u8_u1_U68 (.A( u1_u8_u1_n128 ) , .ZN( u1_u8_u1_n172 ) );
  NAND2_X1 u1_u8_u1_U69 (.A2( u1_u8_u1_n102 ) , .A1( u1_u8_u1_n103 ) , .ZN( u1_u8_u1_n123 ) );
  NAND2_X1 u1_u8_u1_U7 (.ZN( u1_u8_u1_n114 ) , .A1( u1_u8_u1_n134 ) , .A2( u1_u8_u1_n156 ) );
  NOR2_X1 u1_u8_u1_U70 (.A2( u1_u8_X_7 ) , .A1( u1_u8_X_8 ) , .ZN( u1_u8_u1_n95 ) );
  NOR2_X1 u1_u8_u1_U71 (.A1( u1_u8_X_12 ) , .A2( u1_u8_X_9 ) , .ZN( u1_u8_u1_n100 ) );
  NOR2_X1 u1_u8_u1_U72 (.A2( u1_u8_X_8 ) , .A1( u1_u8_u1_n177 ) , .ZN( u1_u8_u1_n99 ) );
  NOR2_X1 u1_u8_u1_U73 (.A2( u1_u8_X_12 ) , .ZN( u1_u8_u1_n102 ) , .A1( u1_u8_u1_n176 ) );
  NOR2_X1 u1_u8_u1_U74 (.A2( u1_u8_X_9 ) , .ZN( u1_u8_u1_n105 ) , .A1( u1_u8_u1_n168 ) );
  NAND2_X1 u1_u8_u1_U75 (.A1( u1_u8_X_10 ) , .ZN( u1_u8_u1_n160 ) , .A2( u1_u8_u1_n169 ) );
  NAND2_X1 u1_u8_u1_U76 (.A2( u1_u8_X_10 ) , .A1( u1_u8_X_11 ) , .ZN( u1_u8_u1_n152 ) );
  NAND2_X1 u1_u8_u1_U77 (.A1( u1_u8_X_11 ) , .ZN( u1_u8_u1_n128 ) , .A2( u1_u8_u1_n170 ) );
  AND2_X1 u1_u8_u1_U78 (.A2( u1_u8_X_7 ) , .A1( u1_u8_X_8 ) , .ZN( u1_u8_u1_n104 ) );
  AND2_X1 u1_u8_u1_U79 (.A1( u1_u8_X_8 ) , .ZN( u1_u8_u1_n103 ) , .A2( u1_u8_u1_n177 ) );
  NOR2_X1 u1_u8_u1_U8 (.A1( u1_u8_u1_n112 ) , .A2( u1_u8_u1_n116 ) , .ZN( u1_u8_u1_n118 ) );
  INV_X1 u1_u8_u1_U80 (.A( u1_u8_X_10 ) , .ZN( u1_u8_u1_n170 ) );
  INV_X1 u1_u8_u1_U81 (.A( u1_u8_X_9 ) , .ZN( u1_u8_u1_n176 ) );
  INV_X1 u1_u8_u1_U82 (.A( u1_u8_X_11 ) , .ZN( u1_u8_u1_n169 ) );
  INV_X1 u1_u8_u1_U83 (.A( u1_u8_X_12 ) , .ZN( u1_u8_u1_n168 ) );
  INV_X1 u1_u8_u1_U84 (.A( u1_u8_X_7 ) , .ZN( u1_u8_u1_n177 ) );
  NAND4_X1 u1_u8_u1_U85 (.ZN( u1_out8_28 ) , .A4( u1_u8_u1_n124 ) , .A3( u1_u8_u1_n125 ) , .A2( u1_u8_u1_n126 ) , .A1( u1_u8_u1_n127 ) );
  OAI21_X1 u1_u8_u1_U86 (.ZN( u1_u8_u1_n127 ) , .B2( u1_u8_u1_n139 ) , .B1( u1_u8_u1_n175 ) , .A( u1_u8_u1_n183 ) );
  OAI21_X1 u1_u8_u1_U87 (.ZN( u1_u8_u1_n126 ) , .B2( u1_u8_u1_n140 ) , .A( u1_u8_u1_n146 ) , .B1( u1_u8_u1_n178 ) );
  NAND4_X1 u1_u8_u1_U88 (.ZN( u1_out8_18 ) , .A4( u1_u8_u1_n165 ) , .A3( u1_u8_u1_n166 ) , .A1( u1_u8_u1_n167 ) , .A2( u1_u8_u1_n186 ) );
  AOI22_X1 u1_u8_u1_U89 (.B2( u1_u8_u1_n146 ) , .B1( u1_u8_u1_n147 ) , .A2( u1_u8_u1_n148 ) , .ZN( u1_u8_u1_n166 ) , .A1( u1_u8_u1_n172 ) );
  OAI21_X1 u1_u8_u1_U9 (.ZN( u1_u8_u1_n101 ) , .B1( u1_u8_u1_n141 ) , .A( u1_u8_u1_n146 ) , .B2( u1_u8_u1_n183 ) );
  INV_X1 u1_u8_u1_U90 (.A( u1_u8_u1_n145 ) , .ZN( u1_u8_u1_n186 ) );
  NAND4_X1 u1_u8_u1_U91 (.ZN( u1_out8_2 ) , .A4( u1_u8_u1_n142 ) , .A3( u1_u8_u1_n143 ) , .A2( u1_u8_u1_n144 ) , .A1( u1_u8_u1_n179 ) );
  OAI21_X1 u1_u8_u1_U92 (.B2( u1_u8_u1_n132 ) , .ZN( u1_u8_u1_n144 ) , .A( u1_u8_u1_n146 ) , .B1( u1_u8_u1_n180 ) );
  INV_X1 u1_u8_u1_U93 (.A( u1_u8_u1_n130 ) , .ZN( u1_u8_u1_n179 ) );
  OR4_X1 u1_u8_u1_U94 (.ZN( u1_out8_13 ) , .A4( u1_u8_u1_n108 ) , .A3( u1_u8_u1_n109 ) , .A2( u1_u8_u1_n110 ) , .A1( u1_u8_u1_n111 ) );
  AOI21_X1 u1_u8_u1_U95 (.ZN( u1_u8_u1_n111 ) , .A( u1_u8_u1_n128 ) , .B2( u1_u8_u1_n131 ) , .B1( u1_u8_u1_n135 ) );
  AOI21_X1 u1_u8_u1_U96 (.ZN( u1_u8_u1_n110 ) , .A( u1_u8_u1_n116 ) , .B1( u1_u8_u1_n152 ) , .B2( u1_u8_u1_n160 ) );
  NAND3_X1 u1_u8_u1_U97 (.A3( u1_u8_u1_n149 ) , .A2( u1_u8_u1_n150 ) , .A1( u1_u8_u1_n151 ) , .ZN( u1_u8_u1_n164 ) );
  NAND3_X1 u1_u8_u1_U98 (.A3( u1_u8_u1_n134 ) , .A2( u1_u8_u1_n135 ) , .ZN( u1_u8_u1_n136 ) , .A1( u1_u8_u1_n151 ) );
  NAND3_X1 u1_u8_u1_U99 (.A1( u1_u8_u1_n133 ) , .ZN( u1_u8_u1_n137 ) , .A2( u1_u8_u1_n154 ) , .A3( u1_u8_u1_n181 ) );
  XOR2_X1 u1_u9_U10 (.B( u1_K10_45 ) , .A( u1_R8_30 ) , .Z( u1_u9_X_45 ) );
  XOR2_X1 u1_u9_U35 (.B( u1_K10_22 ) , .A( u1_R8_15 ) , .Z( u1_u9_X_22 ) );
  XOR2_X1 u1_u9_U36 (.B( u1_K10_21 ) , .A( u1_R8_14 ) , .Z( u1_u9_X_21 ) );
  XOR2_X1 u1_u9_U37 (.B( u1_K10_20 ) , .A( u1_R8_13 ) , .Z( u1_u9_X_20 ) );
  XOR2_X1 u1_u9_U39 (.B( u1_K10_19 ) , .A( u1_R8_12 ) , .Z( u1_u9_X_19 ) );
  XOR2_X1 u1_u9_U40 (.B( u1_K10_18 ) , .A( u1_R8_13 ) , .Z( u1_u9_X_18 ) );
  XOR2_X1 u1_u9_U41 (.B( u1_K10_17 ) , .A( u1_R8_12 ) , .Z( u1_u9_X_17 ) );
  XOR2_X1 u1_u9_U42 (.B( u1_K10_16 ) , .A( u1_R8_11 ) , .Z( u1_u9_X_16 ) );
  XOR2_X1 u1_u9_U43 (.B( u1_K10_15 ) , .A( u1_R8_10 ) , .Z( u1_u9_X_15 ) );
  XOR2_X1 u1_u9_U9 (.B( u1_K10_46 ) , .A( u1_R8_31 ) , .Z( u1_u9_X_46 ) );
  OAI22_X1 u1_u9_u2_U10 (.B1( u1_u9_u2_n151 ) , .A2( u1_u9_u2_n152 ) , .A1( u1_u9_u2_n153 ) , .ZN( u1_u9_u2_n160 ) , .B2( u1_u9_u2_n168 ) );
  NAND3_X1 u1_u9_u2_U100 (.A2( u1_u9_u2_n100 ) , .A1( u1_u9_u2_n104 ) , .A3( u1_u9_u2_n138 ) , .ZN( u1_u9_u2_n98 ) );
  NOR3_X1 u1_u9_u2_U11 (.A1( u1_u9_u2_n150 ) , .ZN( u1_u9_u2_n151 ) , .A3( u1_u9_u2_n175 ) , .A2( u1_u9_u2_n188 ) );
  AOI21_X1 u1_u9_u2_U12 (.B2( u1_u9_u2_n123 ) , .ZN( u1_u9_u2_n125 ) , .A( u1_u9_u2_n171 ) , .B1( u1_u9_u2_n184 ) );
  INV_X1 u1_u9_u2_U13 (.A( u1_u9_u2_n150 ) , .ZN( u1_u9_u2_n184 ) );
  AOI21_X1 u1_u9_u2_U14 (.ZN( u1_u9_u2_n144 ) , .B2( u1_u9_u2_n155 ) , .A( u1_u9_u2_n172 ) , .B1( u1_u9_u2_n185 ) );
  AOI21_X1 u1_u9_u2_U15 (.B2( u1_u9_u2_n143 ) , .ZN( u1_u9_u2_n145 ) , .B1( u1_u9_u2_n152 ) , .A( u1_u9_u2_n171 ) );
  INV_X1 u1_u9_u2_U16 (.A( u1_u9_u2_n156 ) , .ZN( u1_u9_u2_n171 ) );
  INV_X1 u1_u9_u2_U17 (.A( u1_u9_u2_n120 ) , .ZN( u1_u9_u2_n188 ) );
  NAND2_X1 u1_u9_u2_U18 (.A2( u1_u9_u2_n122 ) , .ZN( u1_u9_u2_n150 ) , .A1( u1_u9_u2_n152 ) );
  INV_X1 u1_u9_u2_U19 (.A( u1_u9_u2_n153 ) , .ZN( u1_u9_u2_n170 ) );
  INV_X1 u1_u9_u2_U20 (.A( u1_u9_u2_n137 ) , .ZN( u1_u9_u2_n173 ) );
  NAND2_X1 u1_u9_u2_U21 (.A1( u1_u9_u2_n132 ) , .A2( u1_u9_u2_n139 ) , .ZN( u1_u9_u2_n157 ) );
  INV_X1 u1_u9_u2_U22 (.A( u1_u9_u2_n113 ) , .ZN( u1_u9_u2_n178 ) );
  INV_X1 u1_u9_u2_U23 (.A( u1_u9_u2_n139 ) , .ZN( u1_u9_u2_n175 ) );
  INV_X1 u1_u9_u2_U24 (.A( u1_u9_u2_n155 ) , .ZN( u1_u9_u2_n181 ) );
  INV_X1 u1_u9_u2_U25 (.A( u1_u9_u2_n119 ) , .ZN( u1_u9_u2_n177 ) );
  INV_X1 u1_u9_u2_U26 (.A( u1_u9_u2_n116 ) , .ZN( u1_u9_u2_n180 ) );
  INV_X1 u1_u9_u2_U27 (.A( u1_u9_u2_n131 ) , .ZN( u1_u9_u2_n179 ) );
  INV_X1 u1_u9_u2_U28 (.A( u1_u9_u2_n154 ) , .ZN( u1_u9_u2_n176 ) );
  NAND2_X1 u1_u9_u2_U29 (.A2( u1_u9_u2_n116 ) , .A1( u1_u9_u2_n117 ) , .ZN( u1_u9_u2_n118 ) );
  NOR2_X1 u1_u9_u2_U3 (.ZN( u1_u9_u2_n121 ) , .A2( u1_u9_u2_n177 ) , .A1( u1_u9_u2_n180 ) );
  INV_X1 u1_u9_u2_U30 (.A( u1_u9_u2_n132 ) , .ZN( u1_u9_u2_n182 ) );
  INV_X1 u1_u9_u2_U31 (.A( u1_u9_u2_n158 ) , .ZN( u1_u9_u2_n183 ) );
  OAI21_X1 u1_u9_u2_U32 (.A( u1_u9_u2_n156 ) , .B1( u1_u9_u2_n157 ) , .ZN( u1_u9_u2_n158 ) , .B2( u1_u9_u2_n179 ) );
  NOR2_X1 u1_u9_u2_U33 (.ZN( u1_u9_u2_n156 ) , .A1( u1_u9_u2_n166 ) , .A2( u1_u9_u2_n169 ) );
  NOR2_X1 u1_u9_u2_U34 (.A2( u1_u9_u2_n114 ) , .ZN( u1_u9_u2_n137 ) , .A1( u1_u9_u2_n140 ) );
  NOR2_X1 u1_u9_u2_U35 (.A2( u1_u9_u2_n138 ) , .ZN( u1_u9_u2_n153 ) , .A1( u1_u9_u2_n156 ) );
  AOI211_X1 u1_u9_u2_U36 (.ZN( u1_u9_u2_n130 ) , .C1( u1_u9_u2_n138 ) , .C2( u1_u9_u2_n179 ) , .B( u1_u9_u2_n96 ) , .A( u1_u9_u2_n97 ) );
  OAI22_X1 u1_u9_u2_U37 (.B1( u1_u9_u2_n133 ) , .A2( u1_u9_u2_n137 ) , .A1( u1_u9_u2_n152 ) , .B2( u1_u9_u2_n168 ) , .ZN( u1_u9_u2_n97 ) );
  OAI221_X1 u1_u9_u2_U38 (.B1( u1_u9_u2_n113 ) , .C1( u1_u9_u2_n132 ) , .A( u1_u9_u2_n149 ) , .B2( u1_u9_u2_n171 ) , .C2( u1_u9_u2_n172 ) , .ZN( u1_u9_u2_n96 ) );
  OAI221_X1 u1_u9_u2_U39 (.A( u1_u9_u2_n115 ) , .C2( u1_u9_u2_n123 ) , .B2( u1_u9_u2_n143 ) , .B1( u1_u9_u2_n153 ) , .ZN( u1_u9_u2_n163 ) , .C1( u1_u9_u2_n168 ) );
  INV_X1 u1_u9_u2_U4 (.A( u1_u9_u2_n134 ) , .ZN( u1_u9_u2_n185 ) );
  OAI21_X1 u1_u9_u2_U40 (.A( u1_u9_u2_n114 ) , .ZN( u1_u9_u2_n115 ) , .B1( u1_u9_u2_n176 ) , .B2( u1_u9_u2_n178 ) );
  OAI221_X1 u1_u9_u2_U41 (.A( u1_u9_u2_n135 ) , .B2( u1_u9_u2_n136 ) , .B1( u1_u9_u2_n137 ) , .ZN( u1_u9_u2_n162 ) , .C2( u1_u9_u2_n167 ) , .C1( u1_u9_u2_n185 ) );
  AND3_X1 u1_u9_u2_U42 (.A3( u1_u9_u2_n131 ) , .A2( u1_u9_u2_n132 ) , .A1( u1_u9_u2_n133 ) , .ZN( u1_u9_u2_n136 ) );
  AOI22_X1 u1_u9_u2_U43 (.ZN( u1_u9_u2_n135 ) , .B1( u1_u9_u2_n140 ) , .A1( u1_u9_u2_n156 ) , .B2( u1_u9_u2_n180 ) , .A2( u1_u9_u2_n188 ) );
  AOI21_X1 u1_u9_u2_U44 (.ZN( u1_u9_u2_n149 ) , .B1( u1_u9_u2_n173 ) , .B2( u1_u9_u2_n188 ) , .A( u1_u9_u2_n95 ) );
  AND3_X1 u1_u9_u2_U45 (.A2( u1_u9_u2_n100 ) , .A1( u1_u9_u2_n104 ) , .A3( u1_u9_u2_n156 ) , .ZN( u1_u9_u2_n95 ) );
  OAI21_X1 u1_u9_u2_U46 (.A( u1_u9_u2_n101 ) , .B2( u1_u9_u2_n121 ) , .B1( u1_u9_u2_n153 ) , .ZN( u1_u9_u2_n164 ) );
  NAND2_X1 u1_u9_u2_U47 (.A2( u1_u9_u2_n100 ) , .A1( u1_u9_u2_n107 ) , .ZN( u1_u9_u2_n155 ) );
  NAND2_X1 u1_u9_u2_U48 (.A2( u1_u9_u2_n105 ) , .A1( u1_u9_u2_n108 ) , .ZN( u1_u9_u2_n143 ) );
  NAND2_X1 u1_u9_u2_U49 (.A1( u1_u9_u2_n104 ) , .A2( u1_u9_u2_n106 ) , .ZN( u1_u9_u2_n152 ) );
  NOR4_X1 u1_u9_u2_U5 (.A4( u1_u9_u2_n124 ) , .A3( u1_u9_u2_n125 ) , .A2( u1_u9_u2_n126 ) , .A1( u1_u9_u2_n127 ) , .ZN( u1_u9_u2_n128 ) );
  NAND2_X1 u1_u9_u2_U50 (.A1( u1_u9_u2_n100 ) , .A2( u1_u9_u2_n105 ) , .ZN( u1_u9_u2_n132 ) );
  INV_X1 u1_u9_u2_U51 (.A( u1_u9_u2_n140 ) , .ZN( u1_u9_u2_n168 ) );
  INV_X1 u1_u9_u2_U52 (.A( u1_u9_u2_n138 ) , .ZN( u1_u9_u2_n167 ) );
  OAI21_X1 u1_u9_u2_U53 (.A( u1_u9_u2_n141 ) , .B2( u1_u9_u2_n142 ) , .ZN( u1_u9_u2_n146 ) , .B1( u1_u9_u2_n153 ) );
  OAI21_X1 u1_u9_u2_U54 (.A( u1_u9_u2_n140 ) , .ZN( u1_u9_u2_n141 ) , .B1( u1_u9_u2_n176 ) , .B2( u1_u9_u2_n177 ) );
  NOR3_X1 u1_u9_u2_U55 (.ZN( u1_u9_u2_n142 ) , .A3( u1_u9_u2_n175 ) , .A2( u1_u9_u2_n178 ) , .A1( u1_u9_u2_n181 ) );
  NAND2_X1 u1_u9_u2_U56 (.A1( u1_u9_u2_n102 ) , .A2( u1_u9_u2_n106 ) , .ZN( u1_u9_u2_n113 ) );
  NAND2_X1 u1_u9_u2_U57 (.A1( u1_u9_u2_n106 ) , .A2( u1_u9_u2_n107 ) , .ZN( u1_u9_u2_n131 ) );
  NAND2_X1 u1_u9_u2_U58 (.A1( u1_u9_u2_n103 ) , .A2( u1_u9_u2_n107 ) , .ZN( u1_u9_u2_n139 ) );
  NAND2_X1 u1_u9_u2_U59 (.A1( u1_u9_u2_n103 ) , .A2( u1_u9_u2_n105 ) , .ZN( u1_u9_u2_n133 ) );
  AOI21_X1 u1_u9_u2_U6 (.B2( u1_u9_u2_n119 ) , .ZN( u1_u9_u2_n127 ) , .A( u1_u9_u2_n137 ) , .B1( u1_u9_u2_n155 ) );
  NAND2_X1 u1_u9_u2_U60 (.A1( u1_u9_u2_n102 ) , .A2( u1_u9_u2_n103 ) , .ZN( u1_u9_u2_n154 ) );
  NAND2_X1 u1_u9_u2_U61 (.A2( u1_u9_u2_n103 ) , .A1( u1_u9_u2_n104 ) , .ZN( u1_u9_u2_n119 ) );
  NAND2_X1 u1_u9_u2_U62 (.A2( u1_u9_u2_n107 ) , .A1( u1_u9_u2_n108 ) , .ZN( u1_u9_u2_n123 ) );
  NAND2_X1 u1_u9_u2_U63 (.A1( u1_u9_u2_n104 ) , .A2( u1_u9_u2_n108 ) , .ZN( u1_u9_u2_n122 ) );
  INV_X1 u1_u9_u2_U64 (.A( u1_u9_u2_n114 ) , .ZN( u1_u9_u2_n172 ) );
  NAND2_X1 u1_u9_u2_U65 (.A2( u1_u9_u2_n100 ) , .A1( u1_u9_u2_n102 ) , .ZN( u1_u9_u2_n116 ) );
  NAND2_X1 u1_u9_u2_U66 (.A1( u1_u9_u2_n102 ) , .A2( u1_u9_u2_n108 ) , .ZN( u1_u9_u2_n120 ) );
  NAND2_X1 u1_u9_u2_U67 (.A2( u1_u9_u2_n105 ) , .A1( u1_u9_u2_n106 ) , .ZN( u1_u9_u2_n117 ) );
  INV_X1 u1_u9_u2_U68 (.ZN( u1_u9_u2_n187 ) , .A( u1_u9_u2_n99 ) );
  OAI21_X1 u1_u9_u2_U69 (.B1( u1_u9_u2_n137 ) , .B2( u1_u9_u2_n143 ) , .A( u1_u9_u2_n98 ) , .ZN( u1_u9_u2_n99 ) );
  AOI21_X1 u1_u9_u2_U7 (.ZN( u1_u9_u2_n124 ) , .B1( u1_u9_u2_n131 ) , .B2( u1_u9_u2_n143 ) , .A( u1_u9_u2_n172 ) );
  NOR2_X1 u1_u9_u2_U70 (.A2( u1_u9_X_16 ) , .ZN( u1_u9_u2_n140 ) , .A1( u1_u9_u2_n166 ) );
  NOR2_X1 u1_u9_u2_U71 (.A2( u1_u9_X_13 ) , .A1( u1_u9_X_14 ) , .ZN( u1_u9_u2_n100 ) );
  NOR2_X1 u1_u9_u2_U72 (.A2( u1_u9_X_16 ) , .A1( u1_u9_X_17 ) , .ZN( u1_u9_u2_n138 ) );
  NOR2_X1 u1_u9_u2_U73 (.A2( u1_u9_X_15 ) , .A1( u1_u9_X_18 ) , .ZN( u1_u9_u2_n104 ) );
  NOR2_X1 u1_u9_u2_U74 (.A2( u1_u9_X_14 ) , .ZN( u1_u9_u2_n103 ) , .A1( u1_u9_u2_n174 ) );
  NOR2_X1 u1_u9_u2_U75 (.A2( u1_u9_X_15 ) , .ZN( u1_u9_u2_n102 ) , .A1( u1_u9_u2_n165 ) );
  NOR2_X1 u1_u9_u2_U76 (.A2( u1_u9_X_17 ) , .ZN( u1_u9_u2_n114 ) , .A1( u1_u9_u2_n169 ) );
  AND2_X1 u1_u9_u2_U77 (.A1( u1_u9_X_15 ) , .ZN( u1_u9_u2_n105 ) , .A2( u1_u9_u2_n165 ) );
  AND2_X1 u1_u9_u2_U78 (.A2( u1_u9_X_15 ) , .A1( u1_u9_X_18 ) , .ZN( u1_u9_u2_n107 ) );
  AND2_X1 u1_u9_u2_U79 (.A1( u1_u9_X_14 ) , .ZN( u1_u9_u2_n106 ) , .A2( u1_u9_u2_n174 ) );
  AOI21_X1 u1_u9_u2_U8 (.B2( u1_u9_u2_n120 ) , .B1( u1_u9_u2_n121 ) , .ZN( u1_u9_u2_n126 ) , .A( u1_u9_u2_n167 ) );
  AND2_X1 u1_u9_u2_U80 (.A1( u1_u9_X_13 ) , .A2( u1_u9_X_14 ) , .ZN( u1_u9_u2_n108 ) );
  INV_X1 u1_u9_u2_U81 (.A( u1_u9_X_16 ) , .ZN( u1_u9_u2_n169 ) );
  INV_X1 u1_u9_u2_U82 (.A( u1_u9_X_17 ) , .ZN( u1_u9_u2_n166 ) );
  INV_X1 u1_u9_u2_U83 (.A( u1_u9_X_13 ) , .ZN( u1_u9_u2_n174 ) );
  INV_X1 u1_u9_u2_U84 (.A( u1_u9_X_18 ) , .ZN( u1_u9_u2_n165 ) );
  NAND4_X1 u1_u9_u2_U85 (.ZN( u1_out9_24 ) , .A4( u1_u9_u2_n111 ) , .A3( u1_u9_u2_n112 ) , .A1( u1_u9_u2_n130 ) , .A2( u1_u9_u2_n187 ) );
  AOI221_X1 u1_u9_u2_U86 (.A( u1_u9_u2_n109 ) , .B1( u1_u9_u2_n110 ) , .ZN( u1_u9_u2_n111 ) , .C1( u1_u9_u2_n134 ) , .C2( u1_u9_u2_n170 ) , .B2( u1_u9_u2_n173 ) );
  AOI21_X1 u1_u9_u2_U87 (.ZN( u1_u9_u2_n112 ) , .B2( u1_u9_u2_n156 ) , .A( u1_u9_u2_n164 ) , .B1( u1_u9_u2_n181 ) );
  NAND4_X1 u1_u9_u2_U88 (.ZN( u1_out9_16 ) , .A4( u1_u9_u2_n128 ) , .A3( u1_u9_u2_n129 ) , .A1( u1_u9_u2_n130 ) , .A2( u1_u9_u2_n186 ) );
  AOI22_X1 u1_u9_u2_U89 (.A2( u1_u9_u2_n118 ) , .ZN( u1_u9_u2_n129 ) , .A1( u1_u9_u2_n140 ) , .B1( u1_u9_u2_n157 ) , .B2( u1_u9_u2_n170 ) );
  OAI22_X1 u1_u9_u2_U9 (.ZN( u1_u9_u2_n109 ) , .A2( u1_u9_u2_n113 ) , .B2( u1_u9_u2_n133 ) , .B1( u1_u9_u2_n167 ) , .A1( u1_u9_u2_n168 ) );
  INV_X1 u1_u9_u2_U90 (.A( u1_u9_u2_n163 ) , .ZN( u1_u9_u2_n186 ) );
  NAND4_X1 u1_u9_u2_U91 (.ZN( u1_out9_30 ) , .A4( u1_u9_u2_n147 ) , .A3( u1_u9_u2_n148 ) , .A2( u1_u9_u2_n149 ) , .A1( u1_u9_u2_n187 ) );
  AOI21_X1 u1_u9_u2_U92 (.B2( u1_u9_u2_n138 ) , .ZN( u1_u9_u2_n148 ) , .A( u1_u9_u2_n162 ) , .B1( u1_u9_u2_n182 ) );
  NOR3_X1 u1_u9_u2_U93 (.A3( u1_u9_u2_n144 ) , .A2( u1_u9_u2_n145 ) , .A1( u1_u9_u2_n146 ) , .ZN( u1_u9_u2_n147 ) );
  OR4_X1 u1_u9_u2_U94 (.ZN( u1_out9_6 ) , .A4( u1_u9_u2_n161 ) , .A3( u1_u9_u2_n162 ) , .A2( u1_u9_u2_n163 ) , .A1( u1_u9_u2_n164 ) );
  OR3_X1 u1_u9_u2_U95 (.A2( u1_u9_u2_n159 ) , .A1( u1_u9_u2_n160 ) , .ZN( u1_u9_u2_n161 ) , .A3( u1_u9_u2_n183 ) );
  AOI21_X1 u1_u9_u2_U96 (.B2( u1_u9_u2_n154 ) , .B1( u1_u9_u2_n155 ) , .ZN( u1_u9_u2_n159 ) , .A( u1_u9_u2_n167 ) );
  NAND3_X1 u1_u9_u2_U97 (.A2( u1_u9_u2_n117 ) , .A1( u1_u9_u2_n122 ) , .A3( u1_u9_u2_n123 ) , .ZN( u1_u9_u2_n134 ) );
  NAND3_X1 u1_u9_u2_U98 (.ZN( u1_u9_u2_n110 ) , .A2( u1_u9_u2_n131 ) , .A3( u1_u9_u2_n139 ) , .A1( u1_u9_u2_n154 ) );
  NAND3_X1 u1_u9_u2_U99 (.A2( u1_u9_u2_n100 ) , .ZN( u1_u9_u2_n101 ) , .A1( u1_u9_u2_n104 ) , .A3( u1_u9_u2_n114 ) );
  OAI22_X1 u1_u9_u3_U10 (.B1( u1_u9_u3_n113 ) , .A2( u1_u9_u3_n135 ) , .A1( u1_u9_u3_n150 ) , .B2( u1_u9_u3_n164 ) , .ZN( u1_u9_u3_n98 ) );
  OAI211_X1 u1_u9_u3_U11 (.B( u1_u9_u3_n106 ) , .ZN( u1_u9_u3_n119 ) , .C2( u1_u9_u3_n128 ) , .C1( u1_u9_u3_n167 ) , .A( u1_u9_u3_n181 ) );
  AOI221_X1 u1_u9_u3_U12 (.C1( u1_u9_u3_n105 ) , .ZN( u1_u9_u3_n106 ) , .A( u1_u9_u3_n131 ) , .B2( u1_u9_u3_n132 ) , .C2( u1_u9_u3_n133 ) , .B1( u1_u9_u3_n169 ) );
  INV_X1 u1_u9_u3_U13 (.ZN( u1_u9_u3_n181 ) , .A( u1_u9_u3_n98 ) );
  NAND2_X1 u1_u9_u3_U14 (.ZN( u1_u9_u3_n105 ) , .A2( u1_u9_u3_n130 ) , .A1( u1_u9_u3_n155 ) );
  AOI22_X1 u1_u9_u3_U15 (.B1( u1_u9_u3_n115 ) , .A2( u1_u9_u3_n116 ) , .ZN( u1_u9_u3_n123 ) , .B2( u1_u9_u3_n133 ) , .A1( u1_u9_u3_n169 ) );
  NAND2_X1 u1_u9_u3_U16 (.ZN( u1_u9_u3_n116 ) , .A2( u1_u9_u3_n151 ) , .A1( u1_u9_u3_n182 ) );
  NOR2_X1 u1_u9_u3_U17 (.ZN( u1_u9_u3_n126 ) , .A2( u1_u9_u3_n150 ) , .A1( u1_u9_u3_n164 ) );
  AOI21_X1 u1_u9_u3_U18 (.ZN( u1_u9_u3_n112 ) , .B2( u1_u9_u3_n146 ) , .B1( u1_u9_u3_n155 ) , .A( u1_u9_u3_n167 ) );
  NAND2_X1 u1_u9_u3_U19 (.A1( u1_u9_u3_n135 ) , .ZN( u1_u9_u3_n142 ) , .A2( u1_u9_u3_n164 ) );
  NAND2_X1 u1_u9_u3_U20 (.ZN( u1_u9_u3_n132 ) , .A2( u1_u9_u3_n152 ) , .A1( u1_u9_u3_n156 ) );
  AND2_X1 u1_u9_u3_U21 (.A2( u1_u9_u3_n113 ) , .A1( u1_u9_u3_n114 ) , .ZN( u1_u9_u3_n151 ) );
  INV_X1 u1_u9_u3_U22 (.A( u1_u9_u3_n133 ) , .ZN( u1_u9_u3_n165 ) );
  INV_X1 u1_u9_u3_U23 (.A( u1_u9_u3_n135 ) , .ZN( u1_u9_u3_n170 ) );
  NAND2_X1 u1_u9_u3_U24 (.A1( u1_u9_u3_n107 ) , .A2( u1_u9_u3_n108 ) , .ZN( u1_u9_u3_n140 ) );
  NAND2_X1 u1_u9_u3_U25 (.ZN( u1_u9_u3_n117 ) , .A1( u1_u9_u3_n124 ) , .A2( u1_u9_u3_n148 ) );
  NAND2_X1 u1_u9_u3_U26 (.ZN( u1_u9_u3_n143 ) , .A1( u1_u9_u3_n165 ) , .A2( u1_u9_u3_n167 ) );
  INV_X1 u1_u9_u3_U27 (.A( u1_u9_u3_n130 ) , .ZN( u1_u9_u3_n177 ) );
  INV_X1 u1_u9_u3_U28 (.A( u1_u9_u3_n128 ) , .ZN( u1_u9_u3_n176 ) );
  INV_X1 u1_u9_u3_U29 (.A( u1_u9_u3_n155 ) , .ZN( u1_u9_u3_n174 ) );
  INV_X1 u1_u9_u3_U3 (.A( u1_u9_u3_n129 ) , .ZN( u1_u9_u3_n183 ) );
  INV_X1 u1_u9_u3_U30 (.A( u1_u9_u3_n139 ) , .ZN( u1_u9_u3_n185 ) );
  NOR2_X1 u1_u9_u3_U31 (.ZN( u1_u9_u3_n135 ) , .A2( u1_u9_u3_n141 ) , .A1( u1_u9_u3_n169 ) );
  OAI222_X1 u1_u9_u3_U32 (.C2( u1_u9_u3_n107 ) , .A2( u1_u9_u3_n108 ) , .B1( u1_u9_u3_n135 ) , .ZN( u1_u9_u3_n138 ) , .B2( u1_u9_u3_n146 ) , .C1( u1_u9_u3_n154 ) , .A1( u1_u9_u3_n164 ) );
  NOR4_X1 u1_u9_u3_U33 (.A4( u1_u9_u3_n157 ) , .A3( u1_u9_u3_n158 ) , .A2( u1_u9_u3_n159 ) , .A1( u1_u9_u3_n160 ) , .ZN( u1_u9_u3_n161 ) );
  AOI21_X1 u1_u9_u3_U34 (.B2( u1_u9_u3_n152 ) , .B1( u1_u9_u3_n153 ) , .ZN( u1_u9_u3_n158 ) , .A( u1_u9_u3_n164 ) );
  AOI21_X1 u1_u9_u3_U35 (.A( u1_u9_u3_n154 ) , .B2( u1_u9_u3_n155 ) , .B1( u1_u9_u3_n156 ) , .ZN( u1_u9_u3_n157 ) );
  AOI21_X1 u1_u9_u3_U36 (.A( u1_u9_u3_n149 ) , .B2( u1_u9_u3_n150 ) , .B1( u1_u9_u3_n151 ) , .ZN( u1_u9_u3_n159 ) );
  AOI211_X1 u1_u9_u3_U37 (.ZN( u1_u9_u3_n109 ) , .A( u1_u9_u3_n119 ) , .C2( u1_u9_u3_n129 ) , .B( u1_u9_u3_n138 ) , .C1( u1_u9_u3_n141 ) );
  AOI211_X1 u1_u9_u3_U38 (.B( u1_u9_u3_n119 ) , .A( u1_u9_u3_n120 ) , .C2( u1_u9_u3_n121 ) , .ZN( u1_u9_u3_n122 ) , .C1( u1_u9_u3_n179 ) );
  INV_X1 u1_u9_u3_U39 (.A( u1_u9_u3_n156 ) , .ZN( u1_u9_u3_n179 ) );
  INV_X1 u1_u9_u3_U4 (.A( u1_u9_u3_n140 ) , .ZN( u1_u9_u3_n182 ) );
  OAI22_X1 u1_u9_u3_U40 (.B1( u1_u9_u3_n118 ) , .ZN( u1_u9_u3_n120 ) , .A1( u1_u9_u3_n135 ) , .B2( u1_u9_u3_n154 ) , .A2( u1_u9_u3_n178 ) );
  AND3_X1 u1_u9_u3_U41 (.ZN( u1_u9_u3_n118 ) , .A2( u1_u9_u3_n124 ) , .A1( u1_u9_u3_n144 ) , .A3( u1_u9_u3_n152 ) );
  INV_X1 u1_u9_u3_U42 (.A( u1_u9_u3_n121 ) , .ZN( u1_u9_u3_n164 ) );
  NAND2_X1 u1_u9_u3_U43 (.ZN( u1_u9_u3_n133 ) , .A1( u1_u9_u3_n154 ) , .A2( u1_u9_u3_n164 ) );
  OAI211_X1 u1_u9_u3_U44 (.B( u1_u9_u3_n127 ) , .ZN( u1_u9_u3_n139 ) , .C1( u1_u9_u3_n150 ) , .C2( u1_u9_u3_n154 ) , .A( u1_u9_u3_n184 ) );
  INV_X1 u1_u9_u3_U45 (.A( u1_u9_u3_n125 ) , .ZN( u1_u9_u3_n184 ) );
  AOI221_X1 u1_u9_u3_U46 (.A( u1_u9_u3_n126 ) , .ZN( u1_u9_u3_n127 ) , .C2( u1_u9_u3_n132 ) , .C1( u1_u9_u3_n169 ) , .B2( u1_u9_u3_n170 ) , .B1( u1_u9_u3_n174 ) );
  OAI22_X1 u1_u9_u3_U47 (.A1( u1_u9_u3_n124 ) , .ZN( u1_u9_u3_n125 ) , .B2( u1_u9_u3_n145 ) , .A2( u1_u9_u3_n165 ) , .B1( u1_u9_u3_n167 ) );
  NOR2_X1 u1_u9_u3_U48 (.A1( u1_u9_u3_n113 ) , .ZN( u1_u9_u3_n131 ) , .A2( u1_u9_u3_n154 ) );
  NAND2_X1 u1_u9_u3_U49 (.A1( u1_u9_u3_n103 ) , .ZN( u1_u9_u3_n150 ) , .A2( u1_u9_u3_n99 ) );
  INV_X1 u1_u9_u3_U5 (.A( u1_u9_u3_n117 ) , .ZN( u1_u9_u3_n178 ) );
  NAND2_X1 u1_u9_u3_U50 (.A2( u1_u9_u3_n102 ) , .ZN( u1_u9_u3_n155 ) , .A1( u1_u9_u3_n97 ) );
  INV_X1 u1_u9_u3_U51 (.A( u1_u9_u3_n141 ) , .ZN( u1_u9_u3_n167 ) );
  AOI21_X1 u1_u9_u3_U52 (.B2( u1_u9_u3_n114 ) , .B1( u1_u9_u3_n146 ) , .A( u1_u9_u3_n154 ) , .ZN( u1_u9_u3_n94 ) );
  AOI21_X1 u1_u9_u3_U53 (.ZN( u1_u9_u3_n110 ) , .B2( u1_u9_u3_n142 ) , .B1( u1_u9_u3_n186 ) , .A( u1_u9_u3_n95 ) );
  INV_X1 u1_u9_u3_U54 (.A( u1_u9_u3_n145 ) , .ZN( u1_u9_u3_n186 ) );
  AOI21_X1 u1_u9_u3_U55 (.B1( u1_u9_u3_n124 ) , .A( u1_u9_u3_n149 ) , .B2( u1_u9_u3_n155 ) , .ZN( u1_u9_u3_n95 ) );
  INV_X1 u1_u9_u3_U56 (.A( u1_u9_u3_n149 ) , .ZN( u1_u9_u3_n169 ) );
  NAND2_X1 u1_u9_u3_U57 (.ZN( u1_u9_u3_n124 ) , .A1( u1_u9_u3_n96 ) , .A2( u1_u9_u3_n97 ) );
  NAND2_X1 u1_u9_u3_U58 (.A2( u1_u9_u3_n100 ) , .ZN( u1_u9_u3_n146 ) , .A1( u1_u9_u3_n96 ) );
  NAND2_X1 u1_u9_u3_U59 (.A1( u1_u9_u3_n101 ) , .ZN( u1_u9_u3_n145 ) , .A2( u1_u9_u3_n99 ) );
  AOI221_X1 u1_u9_u3_U6 (.A( u1_u9_u3_n131 ) , .C2( u1_u9_u3_n132 ) , .C1( u1_u9_u3_n133 ) , .ZN( u1_u9_u3_n134 ) , .B1( u1_u9_u3_n143 ) , .B2( u1_u9_u3_n177 ) );
  NAND2_X1 u1_u9_u3_U60 (.A1( u1_u9_u3_n100 ) , .ZN( u1_u9_u3_n156 ) , .A2( u1_u9_u3_n99 ) );
  NAND2_X1 u1_u9_u3_U61 (.A2( u1_u9_u3_n101 ) , .A1( u1_u9_u3_n104 ) , .ZN( u1_u9_u3_n148 ) );
  NAND2_X1 u1_u9_u3_U62 (.A1( u1_u9_u3_n100 ) , .A2( u1_u9_u3_n102 ) , .ZN( u1_u9_u3_n128 ) );
  NAND2_X1 u1_u9_u3_U63 (.A2( u1_u9_u3_n101 ) , .A1( u1_u9_u3_n102 ) , .ZN( u1_u9_u3_n152 ) );
  NAND2_X1 u1_u9_u3_U64 (.A2( u1_u9_u3_n101 ) , .ZN( u1_u9_u3_n114 ) , .A1( u1_u9_u3_n96 ) );
  NAND2_X1 u1_u9_u3_U65 (.ZN( u1_u9_u3_n107 ) , .A1( u1_u9_u3_n97 ) , .A2( u1_u9_u3_n99 ) );
  NAND2_X1 u1_u9_u3_U66 (.A2( u1_u9_u3_n100 ) , .A1( u1_u9_u3_n104 ) , .ZN( u1_u9_u3_n113 ) );
  NAND2_X1 u1_u9_u3_U67 (.A1( u1_u9_u3_n104 ) , .ZN( u1_u9_u3_n153 ) , .A2( u1_u9_u3_n97 ) );
  NAND2_X1 u1_u9_u3_U68 (.A2( u1_u9_u3_n103 ) , .A1( u1_u9_u3_n104 ) , .ZN( u1_u9_u3_n130 ) );
  NAND2_X1 u1_u9_u3_U69 (.A2( u1_u9_u3_n103 ) , .ZN( u1_u9_u3_n144 ) , .A1( u1_u9_u3_n96 ) );
  OAI22_X1 u1_u9_u3_U7 (.B2( u1_u9_u3_n147 ) , .A2( u1_u9_u3_n148 ) , .ZN( u1_u9_u3_n160 ) , .B1( u1_u9_u3_n165 ) , .A1( u1_u9_u3_n168 ) );
  NAND2_X1 u1_u9_u3_U70 (.A1( u1_u9_u3_n102 ) , .A2( u1_u9_u3_n103 ) , .ZN( u1_u9_u3_n108 ) );
  NOR2_X1 u1_u9_u3_U71 (.A2( u1_u9_X_19 ) , .A1( u1_u9_X_20 ) , .ZN( u1_u9_u3_n99 ) );
  NOR2_X1 u1_u9_u3_U72 (.A2( u1_u9_X_21 ) , .A1( u1_u9_X_24 ) , .ZN( u1_u9_u3_n103 ) );
  NOR2_X1 u1_u9_u3_U73 (.A2( u1_u9_X_24 ) , .A1( u1_u9_u3_n171 ) , .ZN( u1_u9_u3_n97 ) );
  NOR2_X1 u1_u9_u3_U74 (.A2( u1_u9_X_23 ) , .ZN( u1_u9_u3_n141 ) , .A1( u1_u9_u3_n166 ) );
  NOR2_X1 u1_u9_u3_U75 (.A2( u1_u9_X_19 ) , .A1( u1_u9_u3_n172 ) , .ZN( u1_u9_u3_n96 ) );
  NAND2_X1 u1_u9_u3_U76 (.A1( u1_u9_X_22 ) , .A2( u1_u9_X_23 ) , .ZN( u1_u9_u3_n154 ) );
  NAND2_X1 u1_u9_u3_U77 (.A1( u1_u9_X_23 ) , .ZN( u1_u9_u3_n149 ) , .A2( u1_u9_u3_n166 ) );
  NOR2_X1 u1_u9_u3_U78 (.A2( u1_u9_X_22 ) , .A1( u1_u9_X_23 ) , .ZN( u1_u9_u3_n121 ) );
  AND2_X1 u1_u9_u3_U79 (.A1( u1_u9_X_24 ) , .ZN( u1_u9_u3_n101 ) , .A2( u1_u9_u3_n171 ) );
  AND3_X1 u1_u9_u3_U8 (.A3( u1_u9_u3_n144 ) , .A2( u1_u9_u3_n145 ) , .A1( u1_u9_u3_n146 ) , .ZN( u1_u9_u3_n147 ) );
  AND2_X1 u1_u9_u3_U80 (.A1( u1_u9_X_19 ) , .ZN( u1_u9_u3_n102 ) , .A2( u1_u9_u3_n172 ) );
  AND2_X1 u1_u9_u3_U81 (.A1( u1_u9_X_21 ) , .A2( u1_u9_X_24 ) , .ZN( u1_u9_u3_n100 ) );
  AND2_X1 u1_u9_u3_U82 (.A2( u1_u9_X_19 ) , .A1( u1_u9_X_20 ) , .ZN( u1_u9_u3_n104 ) );
  INV_X1 u1_u9_u3_U83 (.A( u1_u9_X_22 ) , .ZN( u1_u9_u3_n166 ) );
  INV_X1 u1_u9_u3_U84 (.A( u1_u9_X_21 ) , .ZN( u1_u9_u3_n171 ) );
  INV_X1 u1_u9_u3_U85 (.A( u1_u9_X_20 ) , .ZN( u1_u9_u3_n172 ) );
  OR4_X1 u1_u9_u3_U86 (.ZN( u1_out9_10 ) , .A4( u1_u9_u3_n136 ) , .A3( u1_u9_u3_n137 ) , .A1( u1_u9_u3_n138 ) , .A2( u1_u9_u3_n139 ) );
  OAI222_X1 u1_u9_u3_U87 (.C1( u1_u9_u3_n128 ) , .ZN( u1_u9_u3_n137 ) , .B1( u1_u9_u3_n148 ) , .A2( u1_u9_u3_n150 ) , .B2( u1_u9_u3_n154 ) , .C2( u1_u9_u3_n164 ) , .A1( u1_u9_u3_n167 ) );
  OAI221_X1 u1_u9_u3_U88 (.A( u1_u9_u3_n134 ) , .B2( u1_u9_u3_n135 ) , .ZN( u1_u9_u3_n136 ) , .C1( u1_u9_u3_n149 ) , .B1( u1_u9_u3_n151 ) , .C2( u1_u9_u3_n183 ) );
  NAND4_X1 u1_u9_u3_U89 (.ZN( u1_out9_26 ) , .A4( u1_u9_u3_n109 ) , .A3( u1_u9_u3_n110 ) , .A2( u1_u9_u3_n111 ) , .A1( u1_u9_u3_n173 ) );
  INV_X1 u1_u9_u3_U9 (.A( u1_u9_u3_n143 ) , .ZN( u1_u9_u3_n168 ) );
  INV_X1 u1_u9_u3_U90 (.ZN( u1_u9_u3_n173 ) , .A( u1_u9_u3_n94 ) );
  OAI21_X1 u1_u9_u3_U91 (.ZN( u1_u9_u3_n111 ) , .B2( u1_u9_u3_n117 ) , .A( u1_u9_u3_n133 ) , .B1( u1_u9_u3_n176 ) );
  NAND4_X1 u1_u9_u3_U92 (.ZN( u1_out9_20 ) , .A4( u1_u9_u3_n122 ) , .A3( u1_u9_u3_n123 ) , .A1( u1_u9_u3_n175 ) , .A2( u1_u9_u3_n180 ) );
  INV_X1 u1_u9_u3_U93 (.A( u1_u9_u3_n126 ) , .ZN( u1_u9_u3_n180 ) );
  INV_X1 u1_u9_u3_U94 (.A( u1_u9_u3_n112 ) , .ZN( u1_u9_u3_n175 ) );
  NAND4_X1 u1_u9_u3_U95 (.ZN( u1_out9_1 ) , .A4( u1_u9_u3_n161 ) , .A3( u1_u9_u3_n162 ) , .A2( u1_u9_u3_n163 ) , .A1( u1_u9_u3_n185 ) );
  NAND2_X1 u1_u9_u3_U96 (.ZN( u1_u9_u3_n163 ) , .A2( u1_u9_u3_n170 ) , .A1( u1_u9_u3_n176 ) );
  AOI22_X1 u1_u9_u3_U97 (.B2( u1_u9_u3_n140 ) , .B1( u1_u9_u3_n141 ) , .A2( u1_u9_u3_n142 ) , .ZN( u1_u9_u3_n162 ) , .A1( u1_u9_u3_n177 ) );
  NAND3_X1 u1_u9_u3_U98 (.A1( u1_u9_u3_n114 ) , .ZN( u1_u9_u3_n115 ) , .A2( u1_u9_u3_n145 ) , .A3( u1_u9_u3_n153 ) );
  NAND3_X1 u1_u9_u3_U99 (.ZN( u1_u9_u3_n129 ) , .A2( u1_u9_u3_n144 ) , .A1( u1_u9_u3_n153 ) , .A3( u1_u9_u3_n182 ) );
  AND3_X1 u1_u9_u7_U10 (.A3( u1_u9_u7_n110 ) , .A2( u1_u9_u7_n127 ) , .A1( u1_u9_u7_n132 ) , .ZN( u1_u9_u7_n92 ) );
  OAI21_X1 u1_u9_u7_U11 (.A( u1_u9_u7_n161 ) , .B1( u1_u9_u7_n168 ) , .B2( u1_u9_u7_n173 ) , .ZN( u1_u9_u7_n91 ) );
  AOI211_X1 u1_u9_u7_U12 (.A( u1_u9_u7_n117 ) , .ZN( u1_u9_u7_n118 ) , .C2( u1_u9_u7_n126 ) , .C1( u1_u9_u7_n177 ) , .B( u1_u9_u7_n180 ) );
  OAI22_X1 u1_u9_u7_U13 (.B1( u1_u9_u7_n115 ) , .ZN( u1_u9_u7_n117 ) , .A2( u1_u9_u7_n133 ) , .A1( u1_u9_u7_n137 ) , .B2( u1_u9_u7_n162 ) );
  INV_X1 u1_u9_u7_U14 (.A( u1_u9_u7_n116 ) , .ZN( u1_u9_u7_n180 ) );
  NOR3_X1 u1_u9_u7_U15 (.ZN( u1_u9_u7_n115 ) , .A3( u1_u9_u7_n145 ) , .A2( u1_u9_u7_n168 ) , .A1( u1_u9_u7_n169 ) );
  OAI211_X1 u1_u9_u7_U16 (.B( u1_u9_u7_n122 ) , .A( u1_u9_u7_n123 ) , .C2( u1_u9_u7_n124 ) , .ZN( u1_u9_u7_n154 ) , .C1( u1_u9_u7_n162 ) );
  AOI222_X1 u1_u9_u7_U17 (.ZN( u1_u9_u7_n122 ) , .C2( u1_u9_u7_n126 ) , .C1( u1_u9_u7_n145 ) , .B1( u1_u9_u7_n161 ) , .A2( u1_u9_u7_n165 ) , .B2( u1_u9_u7_n170 ) , .A1( u1_u9_u7_n176 ) );
  INV_X1 u1_u9_u7_U18 (.A( u1_u9_u7_n133 ) , .ZN( u1_u9_u7_n176 ) );
  NOR3_X1 u1_u9_u7_U19 (.A2( u1_u9_u7_n134 ) , .A1( u1_u9_u7_n135 ) , .ZN( u1_u9_u7_n136 ) , .A3( u1_u9_u7_n171 ) );
  NOR2_X1 u1_u9_u7_U20 (.A1( u1_u9_u7_n130 ) , .A2( u1_u9_u7_n134 ) , .ZN( u1_u9_u7_n153 ) );
  INV_X1 u1_u9_u7_U21 (.A( u1_u9_u7_n101 ) , .ZN( u1_u9_u7_n165 ) );
  NOR2_X1 u1_u9_u7_U22 (.ZN( u1_u9_u7_n111 ) , .A2( u1_u9_u7_n134 ) , .A1( u1_u9_u7_n169 ) );
  AOI21_X1 u1_u9_u7_U23 (.ZN( u1_u9_u7_n104 ) , .B2( u1_u9_u7_n112 ) , .B1( u1_u9_u7_n127 ) , .A( u1_u9_u7_n164 ) );
  AOI21_X1 u1_u9_u7_U24 (.ZN( u1_u9_u7_n106 ) , .B1( u1_u9_u7_n133 ) , .B2( u1_u9_u7_n146 ) , .A( u1_u9_u7_n162 ) );
  AOI21_X1 u1_u9_u7_U25 (.A( u1_u9_u7_n101 ) , .ZN( u1_u9_u7_n107 ) , .B2( u1_u9_u7_n128 ) , .B1( u1_u9_u7_n175 ) );
  INV_X1 u1_u9_u7_U26 (.A( u1_u9_u7_n138 ) , .ZN( u1_u9_u7_n171 ) );
  INV_X1 u1_u9_u7_U27 (.A( u1_u9_u7_n131 ) , .ZN( u1_u9_u7_n177 ) );
  INV_X1 u1_u9_u7_U28 (.A( u1_u9_u7_n110 ) , .ZN( u1_u9_u7_n174 ) );
  NAND2_X1 u1_u9_u7_U29 (.A1( u1_u9_u7_n129 ) , .A2( u1_u9_u7_n132 ) , .ZN( u1_u9_u7_n149 ) );
  OAI21_X1 u1_u9_u7_U3 (.ZN( u1_u9_u7_n159 ) , .A( u1_u9_u7_n165 ) , .B2( u1_u9_u7_n171 ) , .B1( u1_u9_u7_n174 ) );
  NAND2_X1 u1_u9_u7_U30 (.A1( u1_u9_u7_n113 ) , .A2( u1_u9_u7_n124 ) , .ZN( u1_u9_u7_n130 ) );
  INV_X1 u1_u9_u7_U31 (.A( u1_u9_u7_n112 ) , .ZN( u1_u9_u7_n173 ) );
  INV_X1 u1_u9_u7_U32 (.A( u1_u9_u7_n128 ) , .ZN( u1_u9_u7_n168 ) );
  INV_X1 u1_u9_u7_U33 (.A( u1_u9_u7_n148 ) , .ZN( u1_u9_u7_n169 ) );
  INV_X1 u1_u9_u7_U34 (.A( u1_u9_u7_n127 ) , .ZN( u1_u9_u7_n179 ) );
  NOR2_X1 u1_u9_u7_U35 (.ZN( u1_u9_u7_n101 ) , .A2( u1_u9_u7_n150 ) , .A1( u1_u9_u7_n156 ) );
  AOI211_X1 u1_u9_u7_U36 (.B( u1_u9_u7_n154 ) , .A( u1_u9_u7_n155 ) , .C1( u1_u9_u7_n156 ) , .ZN( u1_u9_u7_n157 ) , .C2( u1_u9_u7_n172 ) );
  INV_X1 u1_u9_u7_U37 (.A( u1_u9_u7_n153 ) , .ZN( u1_u9_u7_n172 ) );
  AOI211_X1 u1_u9_u7_U38 (.B( u1_u9_u7_n139 ) , .A( u1_u9_u7_n140 ) , .C2( u1_u9_u7_n141 ) , .ZN( u1_u9_u7_n142 ) , .C1( u1_u9_u7_n156 ) );
  NAND4_X1 u1_u9_u7_U39 (.A3( u1_u9_u7_n127 ) , .A2( u1_u9_u7_n128 ) , .A1( u1_u9_u7_n129 ) , .ZN( u1_u9_u7_n141 ) , .A4( u1_u9_u7_n147 ) );
  INV_X1 u1_u9_u7_U4 (.A( u1_u9_u7_n111 ) , .ZN( u1_u9_u7_n170 ) );
  AOI21_X1 u1_u9_u7_U40 (.A( u1_u9_u7_n137 ) , .B1( u1_u9_u7_n138 ) , .ZN( u1_u9_u7_n139 ) , .B2( u1_u9_u7_n146 ) );
  OAI22_X1 u1_u9_u7_U41 (.B1( u1_u9_u7_n136 ) , .ZN( u1_u9_u7_n140 ) , .A1( u1_u9_u7_n153 ) , .B2( u1_u9_u7_n162 ) , .A2( u1_u9_u7_n164 ) );
  AOI21_X1 u1_u9_u7_U42 (.ZN( u1_u9_u7_n123 ) , .B1( u1_u9_u7_n165 ) , .B2( u1_u9_u7_n177 ) , .A( u1_u9_u7_n97 ) );
  AOI21_X1 u1_u9_u7_U43 (.B2( u1_u9_u7_n113 ) , .B1( u1_u9_u7_n124 ) , .A( u1_u9_u7_n125 ) , .ZN( u1_u9_u7_n97 ) );
  INV_X1 u1_u9_u7_U44 (.A( u1_u9_u7_n125 ) , .ZN( u1_u9_u7_n161 ) );
  INV_X1 u1_u9_u7_U45 (.A( u1_u9_u7_n152 ) , .ZN( u1_u9_u7_n162 ) );
  AOI22_X1 u1_u9_u7_U46 (.A2( u1_u9_u7_n114 ) , .ZN( u1_u9_u7_n119 ) , .B1( u1_u9_u7_n130 ) , .A1( u1_u9_u7_n156 ) , .B2( u1_u9_u7_n165 ) );
  NAND2_X1 u1_u9_u7_U47 (.A2( u1_u9_u7_n112 ) , .ZN( u1_u9_u7_n114 ) , .A1( u1_u9_u7_n175 ) );
  AND2_X1 u1_u9_u7_U48 (.ZN( u1_u9_u7_n145 ) , .A2( u1_u9_u7_n98 ) , .A1( u1_u9_u7_n99 ) );
  NOR2_X1 u1_u9_u7_U49 (.ZN( u1_u9_u7_n137 ) , .A1( u1_u9_u7_n150 ) , .A2( u1_u9_u7_n161 ) );
  INV_X1 u1_u9_u7_U5 (.A( u1_u9_u7_n149 ) , .ZN( u1_u9_u7_n175 ) );
  AOI21_X1 u1_u9_u7_U50 (.ZN( u1_u9_u7_n105 ) , .B2( u1_u9_u7_n110 ) , .A( u1_u9_u7_n125 ) , .B1( u1_u9_u7_n147 ) );
  NAND2_X1 u1_u9_u7_U51 (.ZN( u1_u9_u7_n146 ) , .A1( u1_u9_u7_n95 ) , .A2( u1_u9_u7_n98 ) );
  NAND2_X1 u1_u9_u7_U52 (.A2( u1_u9_u7_n103 ) , .ZN( u1_u9_u7_n147 ) , .A1( u1_u9_u7_n93 ) );
  NAND2_X1 u1_u9_u7_U53 (.A1( u1_u9_u7_n103 ) , .ZN( u1_u9_u7_n127 ) , .A2( u1_u9_u7_n99 ) );
  OR2_X1 u1_u9_u7_U54 (.ZN( u1_u9_u7_n126 ) , .A2( u1_u9_u7_n152 ) , .A1( u1_u9_u7_n156 ) );
  NAND2_X1 u1_u9_u7_U55 (.A2( u1_u9_u7_n102 ) , .A1( u1_u9_u7_n103 ) , .ZN( u1_u9_u7_n133 ) );
  NAND2_X1 u1_u9_u7_U56 (.ZN( u1_u9_u7_n112 ) , .A2( u1_u9_u7_n96 ) , .A1( u1_u9_u7_n99 ) );
  NAND2_X1 u1_u9_u7_U57 (.A2( u1_u9_u7_n102 ) , .ZN( u1_u9_u7_n128 ) , .A1( u1_u9_u7_n98 ) );
  NAND2_X1 u1_u9_u7_U58 (.A1( u1_u9_u7_n100 ) , .ZN( u1_u9_u7_n113 ) , .A2( u1_u9_u7_n93 ) );
  NAND2_X1 u1_u9_u7_U59 (.A2( u1_u9_u7_n102 ) , .ZN( u1_u9_u7_n124 ) , .A1( u1_u9_u7_n96 ) );
  INV_X1 u1_u9_u7_U6 (.A( u1_u9_u7_n154 ) , .ZN( u1_u9_u7_n178 ) );
  NAND2_X1 u1_u9_u7_U60 (.ZN( u1_u9_u7_n110 ) , .A1( u1_u9_u7_n95 ) , .A2( u1_u9_u7_n96 ) );
  INV_X1 u1_u9_u7_U61 (.A( u1_u9_u7_n150 ) , .ZN( u1_u9_u7_n164 ) );
  AND2_X1 u1_u9_u7_U62 (.ZN( u1_u9_u7_n134 ) , .A1( u1_u9_u7_n93 ) , .A2( u1_u9_u7_n98 ) );
  NAND2_X1 u1_u9_u7_U63 (.A1( u1_u9_u7_n100 ) , .A2( u1_u9_u7_n102 ) , .ZN( u1_u9_u7_n129 ) );
  NAND2_X1 u1_u9_u7_U64 (.A2( u1_u9_u7_n103 ) , .ZN( u1_u9_u7_n131 ) , .A1( u1_u9_u7_n95 ) );
  NAND2_X1 u1_u9_u7_U65 (.A1( u1_u9_u7_n100 ) , .ZN( u1_u9_u7_n138 ) , .A2( u1_u9_u7_n99 ) );
  NAND2_X1 u1_u9_u7_U66 (.ZN( u1_u9_u7_n132 ) , .A1( u1_u9_u7_n93 ) , .A2( u1_u9_u7_n96 ) );
  NAND2_X1 u1_u9_u7_U67 (.A1( u1_u9_u7_n100 ) , .ZN( u1_u9_u7_n148 ) , .A2( u1_u9_u7_n95 ) );
  NOR2_X1 u1_u9_u7_U68 (.A2( u1_u9_X_47 ) , .ZN( u1_u9_u7_n150 ) , .A1( u1_u9_u7_n163 ) );
  NOR2_X1 u1_u9_u7_U69 (.A2( u1_u9_X_43 ) , .A1( u1_u9_X_44 ) , .ZN( u1_u9_u7_n103 ) );
  AOI211_X1 u1_u9_u7_U7 (.ZN( u1_u9_u7_n116 ) , .A( u1_u9_u7_n155 ) , .C1( u1_u9_u7_n161 ) , .C2( u1_u9_u7_n171 ) , .B( u1_u9_u7_n94 ) );
  NOR2_X1 u1_u9_u7_U70 (.A2( u1_u9_X_48 ) , .A1( u1_u9_u7_n166 ) , .ZN( u1_u9_u7_n95 ) );
  NOR2_X1 u1_u9_u7_U71 (.A2( u1_u9_X_45 ) , .A1( u1_u9_X_48 ) , .ZN( u1_u9_u7_n99 ) );
  NOR2_X1 u1_u9_u7_U72 (.A2( u1_u9_X_44 ) , .A1( u1_u9_u7_n167 ) , .ZN( u1_u9_u7_n98 ) );
  NOR2_X1 u1_u9_u7_U73 (.A2( u1_u9_X_46 ) , .A1( u1_u9_X_47 ) , .ZN( u1_u9_u7_n152 ) );
  AND2_X1 u1_u9_u7_U74 (.A1( u1_u9_X_47 ) , .ZN( u1_u9_u7_n156 ) , .A2( u1_u9_u7_n163 ) );
  NAND2_X1 u1_u9_u7_U75 (.A2( u1_u9_X_46 ) , .A1( u1_u9_X_47 ) , .ZN( u1_u9_u7_n125 ) );
  AND2_X1 u1_u9_u7_U76 (.A2( u1_u9_X_45 ) , .A1( u1_u9_X_48 ) , .ZN( u1_u9_u7_n102 ) );
  AND2_X1 u1_u9_u7_U77 (.A2( u1_u9_X_43 ) , .A1( u1_u9_X_44 ) , .ZN( u1_u9_u7_n96 ) );
  AND2_X1 u1_u9_u7_U78 (.A1( u1_u9_X_44 ) , .ZN( u1_u9_u7_n100 ) , .A2( u1_u9_u7_n167 ) );
  AND2_X1 u1_u9_u7_U79 (.A1( u1_u9_X_48 ) , .A2( u1_u9_u7_n166 ) , .ZN( u1_u9_u7_n93 ) );
  OAI222_X1 u1_u9_u7_U8 (.C2( u1_u9_u7_n101 ) , .B2( u1_u9_u7_n111 ) , .A1( u1_u9_u7_n113 ) , .C1( u1_u9_u7_n146 ) , .A2( u1_u9_u7_n162 ) , .B1( u1_u9_u7_n164 ) , .ZN( u1_u9_u7_n94 ) );
  INV_X1 u1_u9_u7_U80 (.A( u1_u9_X_46 ) , .ZN( u1_u9_u7_n163 ) );
  INV_X1 u1_u9_u7_U81 (.A( u1_u9_X_43 ) , .ZN( u1_u9_u7_n167 ) );
  INV_X1 u1_u9_u7_U82 (.A( u1_u9_X_45 ) , .ZN( u1_u9_u7_n166 ) );
  NAND4_X1 u1_u9_u7_U83 (.ZN( u1_out9_5 ) , .A4( u1_u9_u7_n108 ) , .A3( u1_u9_u7_n109 ) , .A1( u1_u9_u7_n116 ) , .A2( u1_u9_u7_n123 ) );
  AOI22_X1 u1_u9_u7_U84 (.ZN( u1_u9_u7_n109 ) , .A2( u1_u9_u7_n126 ) , .B2( u1_u9_u7_n145 ) , .B1( u1_u9_u7_n156 ) , .A1( u1_u9_u7_n171 ) );
  NOR4_X1 u1_u9_u7_U85 (.A4( u1_u9_u7_n104 ) , .A3( u1_u9_u7_n105 ) , .A2( u1_u9_u7_n106 ) , .A1( u1_u9_u7_n107 ) , .ZN( u1_u9_u7_n108 ) );
  NAND4_X1 u1_u9_u7_U86 (.ZN( u1_out9_27 ) , .A4( u1_u9_u7_n118 ) , .A3( u1_u9_u7_n119 ) , .A2( u1_u9_u7_n120 ) , .A1( u1_u9_u7_n121 ) );
  OAI21_X1 u1_u9_u7_U87 (.ZN( u1_u9_u7_n121 ) , .B2( u1_u9_u7_n145 ) , .A( u1_u9_u7_n150 ) , .B1( u1_u9_u7_n174 ) );
  OAI21_X1 u1_u9_u7_U88 (.ZN( u1_u9_u7_n120 ) , .A( u1_u9_u7_n161 ) , .B2( u1_u9_u7_n170 ) , .B1( u1_u9_u7_n179 ) );
  NAND4_X1 u1_u9_u7_U89 (.ZN( u1_out9_21 ) , .A4( u1_u9_u7_n157 ) , .A3( u1_u9_u7_n158 ) , .A2( u1_u9_u7_n159 ) , .A1( u1_u9_u7_n160 ) );
  OAI221_X1 u1_u9_u7_U9 (.C1( u1_u9_u7_n101 ) , .C2( u1_u9_u7_n147 ) , .ZN( u1_u9_u7_n155 ) , .B2( u1_u9_u7_n162 ) , .A( u1_u9_u7_n91 ) , .B1( u1_u9_u7_n92 ) );
  OAI21_X1 u1_u9_u7_U90 (.B1( u1_u9_u7_n145 ) , .ZN( u1_u9_u7_n160 ) , .A( u1_u9_u7_n161 ) , .B2( u1_u9_u7_n177 ) );
  AOI22_X1 u1_u9_u7_U91 (.B2( u1_u9_u7_n149 ) , .B1( u1_u9_u7_n150 ) , .A2( u1_u9_u7_n151 ) , .A1( u1_u9_u7_n152 ) , .ZN( u1_u9_u7_n158 ) );
  NAND4_X1 u1_u9_u7_U92 (.ZN( u1_out9_15 ) , .A4( u1_u9_u7_n142 ) , .A3( u1_u9_u7_n143 ) , .A2( u1_u9_u7_n144 ) , .A1( u1_u9_u7_n178 ) );
  OR2_X1 u1_u9_u7_U93 (.A2( u1_u9_u7_n125 ) , .A1( u1_u9_u7_n129 ) , .ZN( u1_u9_u7_n144 ) );
  AOI22_X1 u1_u9_u7_U94 (.A2( u1_u9_u7_n126 ) , .ZN( u1_u9_u7_n143 ) , .B2( u1_u9_u7_n165 ) , .B1( u1_u9_u7_n173 ) , .A1( u1_u9_u7_n174 ) );
  NAND3_X1 u1_u9_u7_U95 (.A3( u1_u9_u7_n146 ) , .A2( u1_u9_u7_n147 ) , .A1( u1_u9_u7_n148 ) , .ZN( u1_u9_u7_n151 ) );
  NAND3_X1 u1_u9_u7_U96 (.A3( u1_u9_u7_n131 ) , .A2( u1_u9_u7_n132 ) , .A1( u1_u9_u7_n133 ) , .ZN( u1_u9_u7_n135 ) );
  INV_X1 u1_uk_U1119 (.ZN( u1_K9_11 ) , .A( u1_uk_n1148 ) );
  INV_X1 u1_uk_U1129 (.ZN( u1_K11_8 ) , .A( u1_uk_n501 ) );
  INV_X1 u1_uk_U1131 (.ZN( u1_K11_12 ) , .A( u1_uk_n379 ) );
  INV_X1 u1_uk_U1155 (.ZN( u1_K6_2 ) , .A( u1_uk_n1096 ) );
  INV_X1 u1_uk_U1172 (.ZN( u1_K13_6 ) , .A( u1_uk_n949 ) );
  INV_X1 u1_uk_U144 (.ZN( u1_K12_15 ) , .A( u1_uk_n504 ) );
  INV_X1 u1_uk_U190 (.ZN( u1_K11_14 ) , .A( u1_uk_n382 ) );
  INV_X1 u1_uk_U351 (.ZN( u1_K6_4 ) , .A( u1_uk_n1101 ) );
  INV_X1 u1_uk_U359 (.ZN( u1_K12_4 ) , .A( u1_uk_n656 ) );
  INV_X1 u1_uk_U447 (.ZN( u1_K9_9 ) , .A( u1_uk_n1171 ) );
  INV_X1 u1_uk_U449 (.ZN( u1_K6_9 ) , .A( u1_uk_n1104 ) );
  INV_X1 u1_uk_U587 (.ZN( u1_K9_10 ) , .A( u1_uk_n1147 ) );
  INV_X1 u1_uk_U590 (.ZN( u1_K6_10 ) , .A( u1_uk_n1088 ) );
  INV_X1 u1_uk_U599 (.ZN( u1_K13_22 ) , .A( u1_uk_n692 ) );
  INV_X1 u1_uk_U603 (.ZN( u1_K10_22 ) , .A( u1_uk_n312 ) );
  INV_X1 u1_uk_U610 (.ZN( u1_K1_22 ) , .A( u1_uk_n1004 ) );
  INV_X1 u1_uk_U703 (.ZN( u1_K12_3 ) , .A( u1_uk_n601 ) );
  INV_X1 u1_uk_U783 (.ZN( u1_K13_21 ) , .A( u1_uk_n689 ) );
  INV_X1 u1_uk_U785 (.ZN( u1_K6_21 ) , .A( u1_uk_n1092 ) );
  XOR2_X1 u2_u0_U11 (.B( u2_K1_44 ) , .A( u2_desIn_r_33 ) , .Z( u2_u0_X_44 ) );
  XOR2_X1 u2_u0_U12 (.B( u2_K1_43 ) , .A( u2_desIn_r_25 ) , .Z( u2_u0_X_43 ) );
  XOR2_X1 u2_u0_U13 (.B( u2_K1_42 ) , .A( u2_desIn_r_33 ) , .Z( u2_u0_X_42 ) );
  XOR2_X1 u2_u0_U14 (.B( u2_K1_41 ) , .A( u2_desIn_r_25 ) , .Z( u2_u0_X_41 ) );
  XOR2_X1 u2_u0_U17 (.B( u2_K1_39 ) , .A( u2_desIn_r_9 ) , .Z( u2_u0_X_39 ) );
  XOR2_X1 u2_u0_U18 (.B( u2_K1_38 ) , .A( u2_desIn_r_1 ) , .Z( u2_u0_X_38 ) );
  XOR2_X1 u2_u0_U19 (.B( u2_K1_37 ) , .A( u2_desIn_r_59 ) , .Z( u2_u0_X_37 ) );
  XOR2_X1 u2_u0_U20 (.B( u2_K1_36 ) , .A( u2_desIn_r_1 ) , .Z( u2_u0_X_36 ) );
  XOR2_X1 u2_u0_U21 (.B( u2_K1_35 ) , .A( u2_desIn_r_59 ) , .Z( u2_u0_X_35 ) );
  XOR2_X1 u2_u0_U23 (.B( u2_K1_33 ) , .A( u2_desIn_r_43 ) , .Z( u2_u0_X_33 ) );
  XOR2_X1 u2_u0_U24 (.B( u2_K1_32 ) , .A( u2_desIn_r_35 ) , .Z( u2_u0_X_32 ) );
  XOR2_X1 u2_u0_U25 (.B( u2_K1_31 ) , .A( u2_desIn_r_27 ) , .Z( u2_u0_X_31 ) );
  XOR2_X1 u2_u0_U26 (.B( u2_K1_30 ) , .A( u2_desIn_r_35 ) , .Z( u2_u0_X_30 ) );
  XOR2_X1 u2_u0_U28 (.B( u2_K1_29 ) , .A( u2_desIn_r_27 ) , .Z( u2_u0_X_29 ) );
  XOR2_X1 u2_u0_U30 (.B( u2_K1_27 ) , .A( u2_desIn_r_11 ) , .Z( u2_u0_X_27 ) );
  XOR2_X1 u2_u0_U31 (.B( u2_K1_26 ) , .A( u2_desIn_r_3 ) , .Z( u2_u0_X_26 ) );
  XOR2_X1 u2_u0_U32 (.B( u2_K1_25 ) , .A( u2_desIn_r_61 ) , .Z( u2_u0_X_25 ) );
  XOR2_X1 u2_u0_U7 (.B( u2_K1_48 ) , .A( u2_desIn_r_7 ) , .Z( u2_u0_X_48 ) );
  XOR2_X1 u2_u0_U8 (.B( u2_K1_47 ) , .A( u2_desIn_r_57 ) , .Z( u2_u0_X_47 ) );
  OAI22_X1 u2_u0_u4_U10 (.B2( u2_u0_u4_n135 ) , .ZN( u2_u0_u4_n137 ) , .B1( u2_u0_u4_n153 ) , .A1( u2_u0_u4_n155 ) , .A2( u2_u0_u4_n171 ) );
  AND3_X1 u2_u0_u4_U11 (.A2( u2_u0_u4_n134 ) , .ZN( u2_u0_u4_n135 ) , .A3( u2_u0_u4_n145 ) , .A1( u2_u0_u4_n157 ) );
  NAND2_X1 u2_u0_u4_U12 (.ZN( u2_u0_u4_n132 ) , .A2( u2_u0_u4_n170 ) , .A1( u2_u0_u4_n173 ) );
  AOI21_X1 u2_u0_u4_U13 (.B2( u2_u0_u4_n160 ) , .B1( u2_u0_u4_n161 ) , .ZN( u2_u0_u4_n162 ) , .A( u2_u0_u4_n170 ) );
  AOI21_X1 u2_u0_u4_U14 (.ZN( u2_u0_u4_n107 ) , .B2( u2_u0_u4_n143 ) , .A( u2_u0_u4_n174 ) , .B1( u2_u0_u4_n184 ) );
  AOI21_X1 u2_u0_u4_U15 (.B2( u2_u0_u4_n158 ) , .B1( u2_u0_u4_n159 ) , .ZN( u2_u0_u4_n163 ) , .A( u2_u0_u4_n174 ) );
  AOI21_X1 u2_u0_u4_U16 (.A( u2_u0_u4_n153 ) , .B2( u2_u0_u4_n154 ) , .B1( u2_u0_u4_n155 ) , .ZN( u2_u0_u4_n165 ) );
  AOI21_X1 u2_u0_u4_U17 (.A( u2_u0_u4_n156 ) , .B2( u2_u0_u4_n157 ) , .ZN( u2_u0_u4_n164 ) , .B1( u2_u0_u4_n184 ) );
  INV_X1 u2_u0_u4_U18 (.A( u2_u0_u4_n138 ) , .ZN( u2_u0_u4_n170 ) );
  AND2_X1 u2_u0_u4_U19 (.A2( u2_u0_u4_n120 ) , .ZN( u2_u0_u4_n155 ) , .A1( u2_u0_u4_n160 ) );
  INV_X1 u2_u0_u4_U20 (.A( u2_u0_u4_n156 ) , .ZN( u2_u0_u4_n175 ) );
  NAND2_X1 u2_u0_u4_U21 (.A2( u2_u0_u4_n118 ) , .ZN( u2_u0_u4_n131 ) , .A1( u2_u0_u4_n147 ) );
  NAND2_X1 u2_u0_u4_U22 (.A1( u2_u0_u4_n119 ) , .A2( u2_u0_u4_n120 ) , .ZN( u2_u0_u4_n130 ) );
  NAND2_X1 u2_u0_u4_U23 (.ZN( u2_u0_u4_n117 ) , .A2( u2_u0_u4_n118 ) , .A1( u2_u0_u4_n148 ) );
  NAND2_X1 u2_u0_u4_U24 (.ZN( u2_u0_u4_n129 ) , .A1( u2_u0_u4_n134 ) , .A2( u2_u0_u4_n148 ) );
  AND3_X1 u2_u0_u4_U25 (.A1( u2_u0_u4_n119 ) , .A2( u2_u0_u4_n143 ) , .A3( u2_u0_u4_n154 ) , .ZN( u2_u0_u4_n161 ) );
  AND2_X1 u2_u0_u4_U26 (.A1( u2_u0_u4_n145 ) , .A2( u2_u0_u4_n147 ) , .ZN( u2_u0_u4_n159 ) );
  OR3_X1 u2_u0_u4_U27 (.A3( u2_u0_u4_n114 ) , .A2( u2_u0_u4_n115 ) , .A1( u2_u0_u4_n116 ) , .ZN( u2_u0_u4_n136 ) );
  AOI21_X1 u2_u0_u4_U28 (.A( u2_u0_u4_n113 ) , .ZN( u2_u0_u4_n116 ) , .B2( u2_u0_u4_n173 ) , .B1( u2_u0_u4_n174 ) );
  AOI21_X1 u2_u0_u4_U29 (.ZN( u2_u0_u4_n115 ) , .B2( u2_u0_u4_n145 ) , .B1( u2_u0_u4_n146 ) , .A( u2_u0_u4_n156 ) );
  NOR2_X1 u2_u0_u4_U3 (.ZN( u2_u0_u4_n121 ) , .A1( u2_u0_u4_n181 ) , .A2( u2_u0_u4_n182 ) );
  OAI22_X1 u2_u0_u4_U30 (.ZN( u2_u0_u4_n114 ) , .A2( u2_u0_u4_n121 ) , .B1( u2_u0_u4_n160 ) , .B2( u2_u0_u4_n170 ) , .A1( u2_u0_u4_n171 ) );
  INV_X1 u2_u0_u4_U31 (.A( u2_u0_u4_n158 ) , .ZN( u2_u0_u4_n182 ) );
  INV_X1 u2_u0_u4_U32 (.ZN( u2_u0_u4_n181 ) , .A( u2_u0_u4_n96 ) );
  INV_X1 u2_u0_u4_U33 (.A( u2_u0_u4_n144 ) , .ZN( u2_u0_u4_n179 ) );
  INV_X1 u2_u0_u4_U34 (.A( u2_u0_u4_n157 ) , .ZN( u2_u0_u4_n178 ) );
  NAND2_X1 u2_u0_u4_U35 (.A2( u2_u0_u4_n154 ) , .A1( u2_u0_u4_n96 ) , .ZN( u2_u0_u4_n97 ) );
  INV_X1 u2_u0_u4_U36 (.ZN( u2_u0_u4_n186 ) , .A( u2_u0_u4_n95 ) );
  OAI221_X1 u2_u0_u4_U37 (.C1( u2_u0_u4_n134 ) , .B1( u2_u0_u4_n158 ) , .B2( u2_u0_u4_n171 ) , .C2( u2_u0_u4_n173 ) , .A( u2_u0_u4_n94 ) , .ZN( u2_u0_u4_n95 ) );
  AOI222_X1 u2_u0_u4_U38 (.B2( u2_u0_u4_n132 ) , .A1( u2_u0_u4_n138 ) , .C2( u2_u0_u4_n175 ) , .A2( u2_u0_u4_n179 ) , .C1( u2_u0_u4_n181 ) , .B1( u2_u0_u4_n185 ) , .ZN( u2_u0_u4_n94 ) );
  INV_X1 u2_u0_u4_U39 (.A( u2_u0_u4_n113 ) , .ZN( u2_u0_u4_n185 ) );
  INV_X1 u2_u0_u4_U4 (.A( u2_u0_u4_n117 ) , .ZN( u2_u0_u4_n184 ) );
  INV_X1 u2_u0_u4_U40 (.A( u2_u0_u4_n143 ) , .ZN( u2_u0_u4_n183 ) );
  NOR2_X1 u2_u0_u4_U41 (.ZN( u2_u0_u4_n138 ) , .A1( u2_u0_u4_n168 ) , .A2( u2_u0_u4_n169 ) );
  NOR2_X1 u2_u0_u4_U42 (.A1( u2_u0_u4_n150 ) , .A2( u2_u0_u4_n152 ) , .ZN( u2_u0_u4_n153 ) );
  NOR2_X1 u2_u0_u4_U43 (.A2( u2_u0_u4_n128 ) , .A1( u2_u0_u4_n138 ) , .ZN( u2_u0_u4_n156 ) );
  AOI22_X1 u2_u0_u4_U44 (.B2( u2_u0_u4_n122 ) , .A1( u2_u0_u4_n123 ) , .ZN( u2_u0_u4_n124 ) , .B1( u2_u0_u4_n128 ) , .A2( u2_u0_u4_n172 ) );
  INV_X1 u2_u0_u4_U45 (.A( u2_u0_u4_n153 ) , .ZN( u2_u0_u4_n172 ) );
  NAND2_X1 u2_u0_u4_U46 (.A2( u2_u0_u4_n120 ) , .ZN( u2_u0_u4_n123 ) , .A1( u2_u0_u4_n161 ) );
  AOI22_X1 u2_u0_u4_U47 (.B2( u2_u0_u4_n132 ) , .A2( u2_u0_u4_n133 ) , .ZN( u2_u0_u4_n140 ) , .A1( u2_u0_u4_n150 ) , .B1( u2_u0_u4_n179 ) );
  NAND2_X1 u2_u0_u4_U48 (.ZN( u2_u0_u4_n133 ) , .A2( u2_u0_u4_n146 ) , .A1( u2_u0_u4_n154 ) );
  NAND2_X1 u2_u0_u4_U49 (.A1( u2_u0_u4_n103 ) , .ZN( u2_u0_u4_n154 ) , .A2( u2_u0_u4_n98 ) );
  NOR4_X1 u2_u0_u4_U5 (.A4( u2_u0_u4_n106 ) , .A3( u2_u0_u4_n107 ) , .A2( u2_u0_u4_n108 ) , .A1( u2_u0_u4_n109 ) , .ZN( u2_u0_u4_n110 ) );
  NAND2_X1 u2_u0_u4_U50 (.A1( u2_u0_u4_n101 ) , .ZN( u2_u0_u4_n158 ) , .A2( u2_u0_u4_n99 ) );
  AOI21_X1 u2_u0_u4_U51 (.ZN( u2_u0_u4_n127 ) , .A( u2_u0_u4_n136 ) , .B2( u2_u0_u4_n150 ) , .B1( u2_u0_u4_n180 ) );
  INV_X1 u2_u0_u4_U52 (.A( u2_u0_u4_n160 ) , .ZN( u2_u0_u4_n180 ) );
  NAND2_X1 u2_u0_u4_U53 (.A2( u2_u0_u4_n104 ) , .A1( u2_u0_u4_n105 ) , .ZN( u2_u0_u4_n146 ) );
  NAND2_X1 u2_u0_u4_U54 (.A2( u2_u0_u4_n101 ) , .A1( u2_u0_u4_n102 ) , .ZN( u2_u0_u4_n160 ) );
  NAND2_X1 u2_u0_u4_U55 (.ZN( u2_u0_u4_n134 ) , .A1( u2_u0_u4_n98 ) , .A2( u2_u0_u4_n99 ) );
  NAND2_X1 u2_u0_u4_U56 (.A1( u2_u0_u4_n103 ) , .A2( u2_u0_u4_n104 ) , .ZN( u2_u0_u4_n143 ) );
  NAND2_X1 u2_u0_u4_U57 (.A2( u2_u0_u4_n105 ) , .ZN( u2_u0_u4_n145 ) , .A1( u2_u0_u4_n98 ) );
  NAND2_X1 u2_u0_u4_U58 (.A1( u2_u0_u4_n100 ) , .A2( u2_u0_u4_n105 ) , .ZN( u2_u0_u4_n120 ) );
  NAND2_X1 u2_u0_u4_U59 (.A1( u2_u0_u4_n102 ) , .A2( u2_u0_u4_n104 ) , .ZN( u2_u0_u4_n148 ) );
  AOI21_X1 u2_u0_u4_U6 (.ZN( u2_u0_u4_n106 ) , .B2( u2_u0_u4_n146 ) , .B1( u2_u0_u4_n158 ) , .A( u2_u0_u4_n170 ) );
  NAND2_X1 u2_u0_u4_U60 (.A2( u2_u0_u4_n100 ) , .A1( u2_u0_u4_n103 ) , .ZN( u2_u0_u4_n157 ) );
  INV_X1 u2_u0_u4_U61 (.A( u2_u0_u4_n150 ) , .ZN( u2_u0_u4_n173 ) );
  INV_X1 u2_u0_u4_U62 (.A( u2_u0_u4_n152 ) , .ZN( u2_u0_u4_n171 ) );
  NAND2_X1 u2_u0_u4_U63 (.A1( u2_u0_u4_n100 ) , .ZN( u2_u0_u4_n118 ) , .A2( u2_u0_u4_n99 ) );
  NAND2_X1 u2_u0_u4_U64 (.A2( u2_u0_u4_n100 ) , .A1( u2_u0_u4_n102 ) , .ZN( u2_u0_u4_n144 ) );
  NAND2_X1 u2_u0_u4_U65 (.A2( u2_u0_u4_n101 ) , .A1( u2_u0_u4_n105 ) , .ZN( u2_u0_u4_n96 ) );
  INV_X1 u2_u0_u4_U66 (.A( u2_u0_u4_n128 ) , .ZN( u2_u0_u4_n174 ) );
  NAND2_X1 u2_u0_u4_U67 (.A2( u2_u0_u4_n102 ) , .ZN( u2_u0_u4_n119 ) , .A1( u2_u0_u4_n98 ) );
  NAND2_X1 u2_u0_u4_U68 (.A2( u2_u0_u4_n101 ) , .A1( u2_u0_u4_n103 ) , .ZN( u2_u0_u4_n147 ) );
  NAND2_X1 u2_u0_u4_U69 (.A2( u2_u0_u4_n104 ) , .ZN( u2_u0_u4_n113 ) , .A1( u2_u0_u4_n99 ) );
  AOI21_X1 u2_u0_u4_U7 (.ZN( u2_u0_u4_n108 ) , .B2( u2_u0_u4_n134 ) , .B1( u2_u0_u4_n155 ) , .A( u2_u0_u4_n156 ) );
  NOR2_X1 u2_u0_u4_U70 (.A2( u2_u0_X_28 ) , .ZN( u2_u0_u4_n150 ) , .A1( u2_u0_u4_n168 ) );
  NOR2_X1 u2_u0_u4_U71 (.A2( u2_u0_X_29 ) , .ZN( u2_u0_u4_n152 ) , .A1( u2_u0_u4_n169 ) );
  NOR2_X1 u2_u0_u4_U72 (.A2( u2_u0_X_30 ) , .ZN( u2_u0_u4_n105 ) , .A1( u2_u0_u4_n176 ) );
  NOR2_X1 u2_u0_u4_U73 (.A2( u2_u0_X_26 ) , .ZN( u2_u0_u4_n100 ) , .A1( u2_u0_u4_n177 ) );
  NOR2_X1 u2_u0_u4_U74 (.A2( u2_u0_X_28 ) , .A1( u2_u0_X_29 ) , .ZN( u2_u0_u4_n128 ) );
  NOR2_X1 u2_u0_u4_U75 (.A2( u2_u0_X_27 ) , .A1( u2_u0_X_30 ) , .ZN( u2_u0_u4_n102 ) );
  NOR2_X1 u2_u0_u4_U76 (.A2( u2_u0_X_25 ) , .A1( u2_u0_X_26 ) , .ZN( u2_u0_u4_n98 ) );
  AND2_X1 u2_u0_u4_U77 (.A2( u2_u0_X_25 ) , .A1( u2_u0_X_26 ) , .ZN( u2_u0_u4_n104 ) );
  AND2_X1 u2_u0_u4_U78 (.A1( u2_u0_X_30 ) , .A2( u2_u0_u4_n176 ) , .ZN( u2_u0_u4_n99 ) );
  AND2_X1 u2_u0_u4_U79 (.A1( u2_u0_X_26 ) , .ZN( u2_u0_u4_n101 ) , .A2( u2_u0_u4_n177 ) );
  AOI21_X1 u2_u0_u4_U8 (.ZN( u2_u0_u4_n109 ) , .A( u2_u0_u4_n153 ) , .B1( u2_u0_u4_n159 ) , .B2( u2_u0_u4_n184 ) );
  AND2_X1 u2_u0_u4_U80 (.A1( u2_u0_X_27 ) , .A2( u2_u0_X_30 ) , .ZN( u2_u0_u4_n103 ) );
  INV_X1 u2_u0_u4_U81 (.A( u2_u0_X_28 ) , .ZN( u2_u0_u4_n169 ) );
  INV_X1 u2_u0_u4_U82 (.A( u2_u0_X_29 ) , .ZN( u2_u0_u4_n168 ) );
  INV_X1 u2_u0_u4_U83 (.A( u2_u0_X_25 ) , .ZN( u2_u0_u4_n177 ) );
  INV_X1 u2_u0_u4_U84 (.A( u2_u0_X_27 ) , .ZN( u2_u0_u4_n176 ) );
  NAND4_X1 u2_u0_u4_U85 (.ZN( u2_out0_25 ) , .A4( u2_u0_u4_n139 ) , .A3( u2_u0_u4_n140 ) , .A2( u2_u0_u4_n141 ) , .A1( u2_u0_u4_n142 ) );
  OAI21_X1 u2_u0_u4_U86 (.A( u2_u0_u4_n128 ) , .B2( u2_u0_u4_n129 ) , .B1( u2_u0_u4_n130 ) , .ZN( u2_u0_u4_n142 ) );
  OAI21_X1 u2_u0_u4_U87 (.B2( u2_u0_u4_n131 ) , .ZN( u2_u0_u4_n141 ) , .A( u2_u0_u4_n175 ) , .B1( u2_u0_u4_n183 ) );
  NAND4_X1 u2_u0_u4_U88 (.ZN( u2_out0_14 ) , .A4( u2_u0_u4_n124 ) , .A3( u2_u0_u4_n125 ) , .A2( u2_u0_u4_n126 ) , .A1( u2_u0_u4_n127 ) );
  AOI22_X1 u2_u0_u4_U89 (.B2( u2_u0_u4_n117 ) , .ZN( u2_u0_u4_n126 ) , .A1( u2_u0_u4_n129 ) , .B1( u2_u0_u4_n152 ) , .A2( u2_u0_u4_n175 ) );
  AOI211_X1 u2_u0_u4_U9 (.B( u2_u0_u4_n136 ) , .A( u2_u0_u4_n137 ) , .C2( u2_u0_u4_n138 ) , .ZN( u2_u0_u4_n139 ) , .C1( u2_u0_u4_n182 ) );
  AOI22_X1 u2_u0_u4_U90 (.ZN( u2_u0_u4_n125 ) , .B2( u2_u0_u4_n131 ) , .A2( u2_u0_u4_n132 ) , .B1( u2_u0_u4_n138 ) , .A1( u2_u0_u4_n178 ) );
  NAND4_X1 u2_u0_u4_U91 (.ZN( u2_out0_8 ) , .A4( u2_u0_u4_n110 ) , .A3( u2_u0_u4_n111 ) , .A2( u2_u0_u4_n112 ) , .A1( u2_u0_u4_n186 ) );
  NAND2_X1 u2_u0_u4_U92 (.ZN( u2_u0_u4_n112 ) , .A2( u2_u0_u4_n130 ) , .A1( u2_u0_u4_n150 ) );
  AOI22_X1 u2_u0_u4_U93 (.ZN( u2_u0_u4_n111 ) , .B2( u2_u0_u4_n132 ) , .A1( u2_u0_u4_n152 ) , .B1( u2_u0_u4_n178 ) , .A2( u2_u0_u4_n97 ) );
  AOI22_X1 u2_u0_u4_U94 (.B2( u2_u0_u4_n149 ) , .B1( u2_u0_u4_n150 ) , .A2( u2_u0_u4_n151 ) , .A1( u2_u0_u4_n152 ) , .ZN( u2_u0_u4_n167 ) );
  NOR4_X1 u2_u0_u4_U95 (.A4( u2_u0_u4_n162 ) , .A3( u2_u0_u4_n163 ) , .A2( u2_u0_u4_n164 ) , .A1( u2_u0_u4_n165 ) , .ZN( u2_u0_u4_n166 ) );
  NAND3_X1 u2_u0_u4_U96 (.ZN( u2_out0_3 ) , .A3( u2_u0_u4_n166 ) , .A1( u2_u0_u4_n167 ) , .A2( u2_u0_u4_n186 ) );
  NAND3_X1 u2_u0_u4_U97 (.A3( u2_u0_u4_n146 ) , .A2( u2_u0_u4_n147 ) , .A1( u2_u0_u4_n148 ) , .ZN( u2_u0_u4_n149 ) );
  NAND3_X1 u2_u0_u4_U98 (.A3( u2_u0_u4_n143 ) , .A2( u2_u0_u4_n144 ) , .A1( u2_u0_u4_n145 ) , .ZN( u2_u0_u4_n151 ) );
  NAND3_X1 u2_u0_u4_U99 (.A3( u2_u0_u4_n121 ) , .ZN( u2_u0_u4_n122 ) , .A2( u2_u0_u4_n144 ) , .A1( u2_u0_u4_n154 ) );
  INV_X1 u2_u0_u5_U10 (.A( u2_u0_u5_n121 ) , .ZN( u2_u0_u5_n177 ) );
  NOR3_X1 u2_u0_u5_U100 (.A3( u2_u0_u5_n141 ) , .A1( u2_u0_u5_n142 ) , .ZN( u2_u0_u5_n143 ) , .A2( u2_u0_u5_n191 ) );
  NAND4_X1 u2_u0_u5_U101 (.ZN( u2_out0_4 ) , .A4( u2_u0_u5_n112 ) , .A2( u2_u0_u5_n113 ) , .A1( u2_u0_u5_n114 ) , .A3( u2_u0_u5_n195 ) );
  AOI211_X1 u2_u0_u5_U102 (.A( u2_u0_u5_n110 ) , .C1( u2_u0_u5_n111 ) , .ZN( u2_u0_u5_n112 ) , .B( u2_u0_u5_n118 ) , .C2( u2_u0_u5_n177 ) );
  AOI222_X1 u2_u0_u5_U103 (.ZN( u2_u0_u5_n113 ) , .A1( u2_u0_u5_n131 ) , .C1( u2_u0_u5_n148 ) , .B2( u2_u0_u5_n174 ) , .C2( u2_u0_u5_n178 ) , .A2( u2_u0_u5_n179 ) , .B1( u2_u0_u5_n99 ) );
  NAND3_X1 u2_u0_u5_U104 (.A2( u2_u0_u5_n154 ) , .A3( u2_u0_u5_n158 ) , .A1( u2_u0_u5_n161 ) , .ZN( u2_u0_u5_n99 ) );
  NOR2_X1 u2_u0_u5_U11 (.ZN( u2_u0_u5_n160 ) , .A2( u2_u0_u5_n173 ) , .A1( u2_u0_u5_n177 ) );
  INV_X1 u2_u0_u5_U12 (.A( u2_u0_u5_n150 ) , .ZN( u2_u0_u5_n174 ) );
  AOI21_X1 u2_u0_u5_U13 (.A( u2_u0_u5_n160 ) , .B2( u2_u0_u5_n161 ) , .ZN( u2_u0_u5_n162 ) , .B1( u2_u0_u5_n192 ) );
  INV_X1 u2_u0_u5_U14 (.A( u2_u0_u5_n159 ) , .ZN( u2_u0_u5_n192 ) );
  AOI21_X1 u2_u0_u5_U15 (.A( u2_u0_u5_n156 ) , .B2( u2_u0_u5_n157 ) , .B1( u2_u0_u5_n158 ) , .ZN( u2_u0_u5_n163 ) );
  AOI21_X1 u2_u0_u5_U16 (.B2( u2_u0_u5_n139 ) , .B1( u2_u0_u5_n140 ) , .ZN( u2_u0_u5_n141 ) , .A( u2_u0_u5_n150 ) );
  OAI21_X1 u2_u0_u5_U17 (.A( u2_u0_u5_n133 ) , .B2( u2_u0_u5_n134 ) , .B1( u2_u0_u5_n135 ) , .ZN( u2_u0_u5_n142 ) );
  OAI21_X1 u2_u0_u5_U18 (.ZN( u2_u0_u5_n133 ) , .B2( u2_u0_u5_n147 ) , .A( u2_u0_u5_n173 ) , .B1( u2_u0_u5_n188 ) );
  NAND2_X1 u2_u0_u5_U19 (.A2( u2_u0_u5_n119 ) , .A1( u2_u0_u5_n123 ) , .ZN( u2_u0_u5_n137 ) );
  INV_X1 u2_u0_u5_U20 (.A( u2_u0_u5_n155 ) , .ZN( u2_u0_u5_n194 ) );
  NAND2_X1 u2_u0_u5_U21 (.A1( u2_u0_u5_n121 ) , .ZN( u2_u0_u5_n132 ) , .A2( u2_u0_u5_n172 ) );
  NAND2_X1 u2_u0_u5_U22 (.A2( u2_u0_u5_n122 ) , .ZN( u2_u0_u5_n136 ) , .A1( u2_u0_u5_n154 ) );
  NAND2_X1 u2_u0_u5_U23 (.A2( u2_u0_u5_n119 ) , .A1( u2_u0_u5_n120 ) , .ZN( u2_u0_u5_n159 ) );
  INV_X1 u2_u0_u5_U24 (.A( u2_u0_u5_n156 ) , .ZN( u2_u0_u5_n175 ) );
  INV_X1 u2_u0_u5_U25 (.A( u2_u0_u5_n158 ) , .ZN( u2_u0_u5_n188 ) );
  INV_X1 u2_u0_u5_U26 (.A( u2_u0_u5_n152 ) , .ZN( u2_u0_u5_n179 ) );
  INV_X1 u2_u0_u5_U27 (.A( u2_u0_u5_n140 ) , .ZN( u2_u0_u5_n182 ) );
  INV_X1 u2_u0_u5_U28 (.A( u2_u0_u5_n151 ) , .ZN( u2_u0_u5_n183 ) );
  INV_X1 u2_u0_u5_U29 (.A( u2_u0_u5_n123 ) , .ZN( u2_u0_u5_n185 ) );
  NOR2_X1 u2_u0_u5_U3 (.ZN( u2_u0_u5_n134 ) , .A1( u2_u0_u5_n183 ) , .A2( u2_u0_u5_n190 ) );
  INV_X1 u2_u0_u5_U30 (.A( u2_u0_u5_n161 ) , .ZN( u2_u0_u5_n184 ) );
  INV_X1 u2_u0_u5_U31 (.A( u2_u0_u5_n139 ) , .ZN( u2_u0_u5_n189 ) );
  INV_X1 u2_u0_u5_U32 (.A( u2_u0_u5_n157 ) , .ZN( u2_u0_u5_n190 ) );
  INV_X1 u2_u0_u5_U33 (.A( u2_u0_u5_n120 ) , .ZN( u2_u0_u5_n193 ) );
  NAND2_X1 u2_u0_u5_U34 (.ZN( u2_u0_u5_n111 ) , .A1( u2_u0_u5_n140 ) , .A2( u2_u0_u5_n155 ) );
  NOR2_X1 u2_u0_u5_U35 (.ZN( u2_u0_u5_n100 ) , .A1( u2_u0_u5_n170 ) , .A2( u2_u0_u5_n180 ) );
  INV_X1 u2_u0_u5_U36 (.A( u2_u0_u5_n117 ) , .ZN( u2_u0_u5_n196 ) );
  OAI221_X1 u2_u0_u5_U37 (.A( u2_u0_u5_n116 ) , .ZN( u2_u0_u5_n117 ) , .B2( u2_u0_u5_n119 ) , .C1( u2_u0_u5_n153 ) , .C2( u2_u0_u5_n158 ) , .B1( u2_u0_u5_n172 ) );
  AOI222_X1 u2_u0_u5_U38 (.ZN( u2_u0_u5_n116 ) , .B2( u2_u0_u5_n145 ) , .C1( u2_u0_u5_n148 ) , .A2( u2_u0_u5_n174 ) , .C2( u2_u0_u5_n177 ) , .B1( u2_u0_u5_n187 ) , .A1( u2_u0_u5_n193 ) );
  INV_X1 u2_u0_u5_U39 (.A( u2_u0_u5_n115 ) , .ZN( u2_u0_u5_n187 ) );
  INV_X1 u2_u0_u5_U4 (.A( u2_u0_u5_n138 ) , .ZN( u2_u0_u5_n191 ) );
  AOI22_X1 u2_u0_u5_U40 (.B2( u2_u0_u5_n131 ) , .A2( u2_u0_u5_n146 ) , .ZN( u2_u0_u5_n169 ) , .B1( u2_u0_u5_n174 ) , .A1( u2_u0_u5_n185 ) );
  NOR2_X1 u2_u0_u5_U41 (.A1( u2_u0_u5_n146 ) , .ZN( u2_u0_u5_n150 ) , .A2( u2_u0_u5_n173 ) );
  AOI21_X1 u2_u0_u5_U42 (.A( u2_u0_u5_n118 ) , .B2( u2_u0_u5_n145 ) , .ZN( u2_u0_u5_n168 ) , .B1( u2_u0_u5_n186 ) );
  INV_X1 u2_u0_u5_U43 (.A( u2_u0_u5_n122 ) , .ZN( u2_u0_u5_n186 ) );
  NOR2_X1 u2_u0_u5_U44 (.A1( u2_u0_u5_n146 ) , .ZN( u2_u0_u5_n152 ) , .A2( u2_u0_u5_n176 ) );
  NOR2_X1 u2_u0_u5_U45 (.A1( u2_u0_u5_n115 ) , .ZN( u2_u0_u5_n118 ) , .A2( u2_u0_u5_n153 ) );
  NOR2_X1 u2_u0_u5_U46 (.A2( u2_u0_u5_n145 ) , .ZN( u2_u0_u5_n156 ) , .A1( u2_u0_u5_n174 ) );
  NOR2_X1 u2_u0_u5_U47 (.ZN( u2_u0_u5_n121 ) , .A2( u2_u0_u5_n145 ) , .A1( u2_u0_u5_n176 ) );
  AOI22_X1 u2_u0_u5_U48 (.ZN( u2_u0_u5_n114 ) , .A2( u2_u0_u5_n137 ) , .A1( u2_u0_u5_n145 ) , .B2( u2_u0_u5_n175 ) , .B1( u2_u0_u5_n193 ) );
  OAI211_X1 u2_u0_u5_U49 (.B( u2_u0_u5_n124 ) , .A( u2_u0_u5_n125 ) , .C2( u2_u0_u5_n126 ) , .C1( u2_u0_u5_n127 ) , .ZN( u2_u0_u5_n128 ) );
  OAI21_X1 u2_u0_u5_U5 (.B2( u2_u0_u5_n136 ) , .B1( u2_u0_u5_n137 ) , .ZN( u2_u0_u5_n138 ) , .A( u2_u0_u5_n177 ) );
  NOR3_X1 u2_u0_u5_U50 (.ZN( u2_u0_u5_n127 ) , .A1( u2_u0_u5_n136 ) , .A3( u2_u0_u5_n148 ) , .A2( u2_u0_u5_n182 ) );
  OAI21_X1 u2_u0_u5_U51 (.ZN( u2_u0_u5_n124 ) , .A( u2_u0_u5_n177 ) , .B2( u2_u0_u5_n183 ) , .B1( u2_u0_u5_n189 ) );
  OAI21_X1 u2_u0_u5_U52 (.ZN( u2_u0_u5_n125 ) , .A( u2_u0_u5_n174 ) , .B2( u2_u0_u5_n185 ) , .B1( u2_u0_u5_n190 ) );
  AOI21_X1 u2_u0_u5_U53 (.A( u2_u0_u5_n153 ) , .B2( u2_u0_u5_n154 ) , .B1( u2_u0_u5_n155 ) , .ZN( u2_u0_u5_n164 ) );
  AOI21_X1 u2_u0_u5_U54 (.ZN( u2_u0_u5_n110 ) , .B1( u2_u0_u5_n122 ) , .B2( u2_u0_u5_n139 ) , .A( u2_u0_u5_n153 ) );
  INV_X1 u2_u0_u5_U55 (.A( u2_u0_u5_n153 ) , .ZN( u2_u0_u5_n176 ) );
  INV_X1 u2_u0_u5_U56 (.A( u2_u0_u5_n126 ) , .ZN( u2_u0_u5_n173 ) );
  AND2_X1 u2_u0_u5_U57 (.A2( u2_u0_u5_n104 ) , .A1( u2_u0_u5_n107 ) , .ZN( u2_u0_u5_n147 ) );
  AND2_X1 u2_u0_u5_U58 (.A2( u2_u0_u5_n104 ) , .A1( u2_u0_u5_n108 ) , .ZN( u2_u0_u5_n148 ) );
  NAND2_X1 u2_u0_u5_U59 (.A1( u2_u0_u5_n105 ) , .A2( u2_u0_u5_n106 ) , .ZN( u2_u0_u5_n158 ) );
  INV_X1 u2_u0_u5_U6 (.A( u2_u0_u5_n135 ) , .ZN( u2_u0_u5_n178 ) );
  NAND2_X1 u2_u0_u5_U60 (.A2( u2_u0_u5_n108 ) , .A1( u2_u0_u5_n109 ) , .ZN( u2_u0_u5_n139 ) );
  NAND2_X1 u2_u0_u5_U61 (.A1( u2_u0_u5_n106 ) , .A2( u2_u0_u5_n108 ) , .ZN( u2_u0_u5_n119 ) );
  NAND2_X1 u2_u0_u5_U62 (.A2( u2_u0_u5_n103 ) , .A1( u2_u0_u5_n105 ) , .ZN( u2_u0_u5_n140 ) );
  NAND2_X1 u2_u0_u5_U63 (.A2( u2_u0_u5_n104 ) , .A1( u2_u0_u5_n105 ) , .ZN( u2_u0_u5_n155 ) );
  NAND2_X1 u2_u0_u5_U64 (.A2( u2_u0_u5_n106 ) , .A1( u2_u0_u5_n107 ) , .ZN( u2_u0_u5_n122 ) );
  NAND2_X1 u2_u0_u5_U65 (.A2( u2_u0_u5_n100 ) , .A1( u2_u0_u5_n106 ) , .ZN( u2_u0_u5_n115 ) );
  NAND2_X1 u2_u0_u5_U66 (.A2( u2_u0_u5_n100 ) , .A1( u2_u0_u5_n103 ) , .ZN( u2_u0_u5_n161 ) );
  NAND2_X1 u2_u0_u5_U67 (.A1( u2_u0_u5_n105 ) , .A2( u2_u0_u5_n109 ) , .ZN( u2_u0_u5_n154 ) );
  INV_X1 u2_u0_u5_U68 (.A( u2_u0_u5_n146 ) , .ZN( u2_u0_u5_n172 ) );
  NAND2_X1 u2_u0_u5_U69 (.A1( u2_u0_u5_n103 ) , .A2( u2_u0_u5_n108 ) , .ZN( u2_u0_u5_n123 ) );
  OAI22_X1 u2_u0_u5_U7 (.B2( u2_u0_u5_n149 ) , .B1( u2_u0_u5_n150 ) , .A2( u2_u0_u5_n151 ) , .A1( u2_u0_u5_n152 ) , .ZN( u2_u0_u5_n165 ) );
  NAND2_X1 u2_u0_u5_U70 (.A2( u2_u0_u5_n103 ) , .A1( u2_u0_u5_n107 ) , .ZN( u2_u0_u5_n151 ) );
  NAND2_X1 u2_u0_u5_U71 (.A2( u2_u0_u5_n107 ) , .A1( u2_u0_u5_n109 ) , .ZN( u2_u0_u5_n120 ) );
  NAND2_X1 u2_u0_u5_U72 (.A2( u2_u0_u5_n100 ) , .A1( u2_u0_u5_n109 ) , .ZN( u2_u0_u5_n157 ) );
  AND2_X1 u2_u0_u5_U73 (.A2( u2_u0_u5_n100 ) , .A1( u2_u0_u5_n104 ) , .ZN( u2_u0_u5_n131 ) );
  INV_X1 u2_u0_u5_U74 (.A( u2_u0_u5_n102 ) , .ZN( u2_u0_u5_n195 ) );
  OAI221_X1 u2_u0_u5_U75 (.A( u2_u0_u5_n101 ) , .ZN( u2_u0_u5_n102 ) , .C2( u2_u0_u5_n115 ) , .C1( u2_u0_u5_n126 ) , .B1( u2_u0_u5_n134 ) , .B2( u2_u0_u5_n160 ) );
  OAI21_X1 u2_u0_u5_U76 (.ZN( u2_u0_u5_n101 ) , .B1( u2_u0_u5_n137 ) , .A( u2_u0_u5_n146 ) , .B2( u2_u0_u5_n147 ) );
  NOR2_X1 u2_u0_u5_U77 (.A2( u2_u0_X_34 ) , .A1( u2_u0_X_35 ) , .ZN( u2_u0_u5_n145 ) );
  NOR2_X1 u2_u0_u5_U78 (.A2( u2_u0_X_34 ) , .ZN( u2_u0_u5_n146 ) , .A1( u2_u0_u5_n171 ) );
  NOR2_X1 u2_u0_u5_U79 (.A2( u2_u0_X_31 ) , .A1( u2_u0_X_32 ) , .ZN( u2_u0_u5_n103 ) );
  NOR3_X1 u2_u0_u5_U8 (.A2( u2_u0_u5_n147 ) , .A1( u2_u0_u5_n148 ) , .ZN( u2_u0_u5_n149 ) , .A3( u2_u0_u5_n194 ) );
  NOR2_X1 u2_u0_u5_U80 (.A2( u2_u0_X_36 ) , .ZN( u2_u0_u5_n105 ) , .A1( u2_u0_u5_n180 ) );
  NOR2_X1 u2_u0_u5_U81 (.A2( u2_u0_X_33 ) , .ZN( u2_u0_u5_n108 ) , .A1( u2_u0_u5_n170 ) );
  NOR2_X1 u2_u0_u5_U82 (.A2( u2_u0_X_33 ) , .A1( u2_u0_X_36 ) , .ZN( u2_u0_u5_n107 ) );
  NOR2_X1 u2_u0_u5_U83 (.A2( u2_u0_X_31 ) , .ZN( u2_u0_u5_n104 ) , .A1( u2_u0_u5_n181 ) );
  NAND2_X1 u2_u0_u5_U84 (.A2( u2_u0_X_34 ) , .A1( u2_u0_X_35 ) , .ZN( u2_u0_u5_n153 ) );
  NAND2_X1 u2_u0_u5_U85 (.A1( u2_u0_X_34 ) , .ZN( u2_u0_u5_n126 ) , .A2( u2_u0_u5_n171 ) );
  AND2_X1 u2_u0_u5_U86 (.A1( u2_u0_X_31 ) , .A2( u2_u0_X_32 ) , .ZN( u2_u0_u5_n106 ) );
  AND2_X1 u2_u0_u5_U87 (.A1( u2_u0_X_31 ) , .ZN( u2_u0_u5_n109 ) , .A2( u2_u0_u5_n181 ) );
  INV_X1 u2_u0_u5_U88 (.A( u2_u0_X_33 ) , .ZN( u2_u0_u5_n180 ) );
  INV_X1 u2_u0_u5_U89 (.A( u2_u0_X_35 ) , .ZN( u2_u0_u5_n171 ) );
  NOR2_X1 u2_u0_u5_U9 (.ZN( u2_u0_u5_n135 ) , .A1( u2_u0_u5_n173 ) , .A2( u2_u0_u5_n176 ) );
  INV_X1 u2_u0_u5_U90 (.A( u2_u0_X_36 ) , .ZN( u2_u0_u5_n170 ) );
  INV_X1 u2_u0_u5_U91 (.A( u2_u0_X_32 ) , .ZN( u2_u0_u5_n181 ) );
  NAND4_X1 u2_u0_u5_U92 (.ZN( u2_out0_29 ) , .A4( u2_u0_u5_n129 ) , .A3( u2_u0_u5_n130 ) , .A2( u2_u0_u5_n168 ) , .A1( u2_u0_u5_n196 ) );
  AOI221_X1 u2_u0_u5_U93 (.A( u2_u0_u5_n128 ) , .ZN( u2_u0_u5_n129 ) , .C2( u2_u0_u5_n132 ) , .B2( u2_u0_u5_n159 ) , .B1( u2_u0_u5_n176 ) , .C1( u2_u0_u5_n184 ) );
  AOI222_X1 u2_u0_u5_U94 (.ZN( u2_u0_u5_n130 ) , .A2( u2_u0_u5_n146 ) , .B1( u2_u0_u5_n147 ) , .C2( u2_u0_u5_n175 ) , .B2( u2_u0_u5_n179 ) , .A1( u2_u0_u5_n188 ) , .C1( u2_u0_u5_n194 ) );
  NAND4_X1 u2_u0_u5_U95 (.ZN( u2_out0_19 ) , .A4( u2_u0_u5_n166 ) , .A3( u2_u0_u5_n167 ) , .A2( u2_u0_u5_n168 ) , .A1( u2_u0_u5_n169 ) );
  AOI22_X1 u2_u0_u5_U96 (.B2( u2_u0_u5_n145 ) , .A2( u2_u0_u5_n146 ) , .ZN( u2_u0_u5_n167 ) , .B1( u2_u0_u5_n182 ) , .A1( u2_u0_u5_n189 ) );
  NOR4_X1 u2_u0_u5_U97 (.A4( u2_u0_u5_n162 ) , .A3( u2_u0_u5_n163 ) , .A2( u2_u0_u5_n164 ) , .A1( u2_u0_u5_n165 ) , .ZN( u2_u0_u5_n166 ) );
  NAND4_X1 u2_u0_u5_U98 (.ZN( u2_out0_11 ) , .A4( u2_u0_u5_n143 ) , .A3( u2_u0_u5_n144 ) , .A2( u2_u0_u5_n169 ) , .A1( u2_u0_u5_n196 ) );
  AOI22_X1 u2_u0_u5_U99 (.A2( u2_u0_u5_n132 ) , .ZN( u2_u0_u5_n144 ) , .B2( u2_u0_u5_n145 ) , .B1( u2_u0_u5_n184 ) , .A1( u2_u0_u5_n194 ) );
  AOI22_X1 u2_u0_u6_U10 (.A2( u2_u0_u6_n151 ) , .B2( u2_u0_u6_n161 ) , .A1( u2_u0_u6_n167 ) , .B1( u2_u0_u6_n170 ) , .ZN( u2_u0_u6_n89 ) );
  AOI21_X1 u2_u0_u6_U11 (.B1( u2_u0_u6_n107 ) , .B2( u2_u0_u6_n132 ) , .A( u2_u0_u6_n158 ) , .ZN( u2_u0_u6_n88 ) );
  AOI21_X1 u2_u0_u6_U12 (.B2( u2_u0_u6_n147 ) , .B1( u2_u0_u6_n148 ) , .ZN( u2_u0_u6_n149 ) , .A( u2_u0_u6_n158 ) );
  AOI21_X1 u2_u0_u6_U13 (.ZN( u2_u0_u6_n106 ) , .A( u2_u0_u6_n142 ) , .B2( u2_u0_u6_n159 ) , .B1( u2_u0_u6_n164 ) );
  INV_X1 u2_u0_u6_U14 (.A( u2_u0_u6_n155 ) , .ZN( u2_u0_u6_n161 ) );
  INV_X1 u2_u0_u6_U15 (.A( u2_u0_u6_n128 ) , .ZN( u2_u0_u6_n164 ) );
  NAND2_X1 u2_u0_u6_U16 (.ZN( u2_u0_u6_n110 ) , .A1( u2_u0_u6_n122 ) , .A2( u2_u0_u6_n129 ) );
  NAND2_X1 u2_u0_u6_U17 (.ZN( u2_u0_u6_n124 ) , .A2( u2_u0_u6_n146 ) , .A1( u2_u0_u6_n148 ) );
  INV_X1 u2_u0_u6_U18 (.A( u2_u0_u6_n132 ) , .ZN( u2_u0_u6_n171 ) );
  AND2_X1 u2_u0_u6_U19 (.A1( u2_u0_u6_n100 ) , .ZN( u2_u0_u6_n130 ) , .A2( u2_u0_u6_n147 ) );
  INV_X1 u2_u0_u6_U20 (.A( u2_u0_u6_n127 ) , .ZN( u2_u0_u6_n173 ) );
  INV_X1 u2_u0_u6_U21 (.A( u2_u0_u6_n121 ) , .ZN( u2_u0_u6_n167 ) );
  INV_X1 u2_u0_u6_U22 (.A( u2_u0_u6_n100 ) , .ZN( u2_u0_u6_n169 ) );
  INV_X1 u2_u0_u6_U23 (.A( u2_u0_u6_n123 ) , .ZN( u2_u0_u6_n170 ) );
  INV_X1 u2_u0_u6_U24 (.A( u2_u0_u6_n113 ) , .ZN( u2_u0_u6_n168 ) );
  AND2_X1 u2_u0_u6_U25 (.A1( u2_u0_u6_n107 ) , .A2( u2_u0_u6_n119 ) , .ZN( u2_u0_u6_n133 ) );
  AND2_X1 u2_u0_u6_U26 (.A2( u2_u0_u6_n121 ) , .A1( u2_u0_u6_n122 ) , .ZN( u2_u0_u6_n131 ) );
  AND3_X1 u2_u0_u6_U27 (.ZN( u2_u0_u6_n120 ) , .A2( u2_u0_u6_n127 ) , .A1( u2_u0_u6_n132 ) , .A3( u2_u0_u6_n145 ) );
  INV_X1 u2_u0_u6_U28 (.A( u2_u0_u6_n146 ) , .ZN( u2_u0_u6_n163 ) );
  AOI222_X1 u2_u0_u6_U29 (.ZN( u2_u0_u6_n114 ) , .A1( u2_u0_u6_n118 ) , .A2( u2_u0_u6_n126 ) , .B2( u2_u0_u6_n151 ) , .C2( u2_u0_u6_n159 ) , .C1( u2_u0_u6_n168 ) , .B1( u2_u0_u6_n169 ) );
  INV_X1 u2_u0_u6_U3 (.A( u2_u0_u6_n110 ) , .ZN( u2_u0_u6_n166 ) );
  NOR2_X1 u2_u0_u6_U30 (.A1( u2_u0_u6_n162 ) , .A2( u2_u0_u6_n165 ) , .ZN( u2_u0_u6_n98 ) );
  AOI211_X1 u2_u0_u6_U31 (.B( u2_u0_u6_n134 ) , .A( u2_u0_u6_n135 ) , .C1( u2_u0_u6_n136 ) , .ZN( u2_u0_u6_n137 ) , .C2( u2_u0_u6_n151 ) );
  AOI21_X1 u2_u0_u6_U32 (.B2( u2_u0_u6_n132 ) , .B1( u2_u0_u6_n133 ) , .ZN( u2_u0_u6_n134 ) , .A( u2_u0_u6_n158 ) );
  NAND4_X1 u2_u0_u6_U33 (.A4( u2_u0_u6_n127 ) , .A3( u2_u0_u6_n128 ) , .A2( u2_u0_u6_n129 ) , .A1( u2_u0_u6_n130 ) , .ZN( u2_u0_u6_n136 ) );
  AOI21_X1 u2_u0_u6_U34 (.B1( u2_u0_u6_n131 ) , .ZN( u2_u0_u6_n135 ) , .A( u2_u0_u6_n144 ) , .B2( u2_u0_u6_n146 ) );
  NAND2_X1 u2_u0_u6_U35 (.A1( u2_u0_u6_n144 ) , .ZN( u2_u0_u6_n151 ) , .A2( u2_u0_u6_n158 ) );
  NAND2_X1 u2_u0_u6_U36 (.ZN( u2_u0_u6_n132 ) , .A1( u2_u0_u6_n91 ) , .A2( u2_u0_u6_n97 ) );
  AOI22_X1 u2_u0_u6_U37 (.B2( u2_u0_u6_n110 ) , .B1( u2_u0_u6_n111 ) , .A1( u2_u0_u6_n112 ) , .ZN( u2_u0_u6_n115 ) , .A2( u2_u0_u6_n161 ) );
  NAND4_X1 u2_u0_u6_U38 (.A3( u2_u0_u6_n109 ) , .ZN( u2_u0_u6_n112 ) , .A4( u2_u0_u6_n132 ) , .A2( u2_u0_u6_n147 ) , .A1( u2_u0_u6_n166 ) );
  NOR2_X1 u2_u0_u6_U39 (.ZN( u2_u0_u6_n109 ) , .A1( u2_u0_u6_n170 ) , .A2( u2_u0_u6_n173 ) );
  INV_X1 u2_u0_u6_U4 (.A( u2_u0_u6_n142 ) , .ZN( u2_u0_u6_n174 ) );
  NOR2_X1 u2_u0_u6_U40 (.A2( u2_u0_u6_n126 ) , .ZN( u2_u0_u6_n155 ) , .A1( u2_u0_u6_n160 ) );
  NAND2_X1 u2_u0_u6_U41 (.ZN( u2_u0_u6_n146 ) , .A2( u2_u0_u6_n94 ) , .A1( u2_u0_u6_n99 ) );
  AOI21_X1 u2_u0_u6_U42 (.A( u2_u0_u6_n144 ) , .B2( u2_u0_u6_n145 ) , .B1( u2_u0_u6_n146 ) , .ZN( u2_u0_u6_n150 ) );
  INV_X1 u2_u0_u6_U43 (.A( u2_u0_u6_n111 ) , .ZN( u2_u0_u6_n158 ) );
  NAND2_X1 u2_u0_u6_U44 (.ZN( u2_u0_u6_n127 ) , .A1( u2_u0_u6_n91 ) , .A2( u2_u0_u6_n92 ) );
  NAND2_X1 u2_u0_u6_U45 (.ZN( u2_u0_u6_n129 ) , .A2( u2_u0_u6_n95 ) , .A1( u2_u0_u6_n96 ) );
  INV_X1 u2_u0_u6_U46 (.A( u2_u0_u6_n144 ) , .ZN( u2_u0_u6_n159 ) );
  NAND2_X1 u2_u0_u6_U47 (.ZN( u2_u0_u6_n145 ) , .A2( u2_u0_u6_n97 ) , .A1( u2_u0_u6_n98 ) );
  NAND2_X1 u2_u0_u6_U48 (.ZN( u2_u0_u6_n148 ) , .A2( u2_u0_u6_n92 ) , .A1( u2_u0_u6_n94 ) );
  NAND2_X1 u2_u0_u6_U49 (.ZN( u2_u0_u6_n108 ) , .A2( u2_u0_u6_n139 ) , .A1( u2_u0_u6_n144 ) );
  NAND2_X1 u2_u0_u6_U5 (.A2( u2_u0_u6_n143 ) , .ZN( u2_u0_u6_n152 ) , .A1( u2_u0_u6_n166 ) );
  NAND2_X1 u2_u0_u6_U50 (.ZN( u2_u0_u6_n121 ) , .A2( u2_u0_u6_n95 ) , .A1( u2_u0_u6_n97 ) );
  NAND2_X1 u2_u0_u6_U51 (.ZN( u2_u0_u6_n107 ) , .A2( u2_u0_u6_n92 ) , .A1( u2_u0_u6_n95 ) );
  AND2_X1 u2_u0_u6_U52 (.ZN( u2_u0_u6_n118 ) , .A2( u2_u0_u6_n91 ) , .A1( u2_u0_u6_n99 ) );
  NAND2_X1 u2_u0_u6_U53 (.ZN( u2_u0_u6_n147 ) , .A2( u2_u0_u6_n98 ) , .A1( u2_u0_u6_n99 ) );
  NAND2_X1 u2_u0_u6_U54 (.ZN( u2_u0_u6_n128 ) , .A1( u2_u0_u6_n94 ) , .A2( u2_u0_u6_n96 ) );
  NAND2_X1 u2_u0_u6_U55 (.ZN( u2_u0_u6_n119 ) , .A2( u2_u0_u6_n95 ) , .A1( u2_u0_u6_n99 ) );
  NAND2_X1 u2_u0_u6_U56 (.ZN( u2_u0_u6_n123 ) , .A2( u2_u0_u6_n91 ) , .A1( u2_u0_u6_n96 ) );
  NAND2_X1 u2_u0_u6_U57 (.ZN( u2_u0_u6_n100 ) , .A2( u2_u0_u6_n92 ) , .A1( u2_u0_u6_n98 ) );
  NAND2_X1 u2_u0_u6_U58 (.ZN( u2_u0_u6_n122 ) , .A1( u2_u0_u6_n94 ) , .A2( u2_u0_u6_n97 ) );
  INV_X1 u2_u0_u6_U59 (.A( u2_u0_u6_n139 ) , .ZN( u2_u0_u6_n160 ) );
  AOI22_X1 u2_u0_u6_U6 (.B2( u2_u0_u6_n101 ) , .A1( u2_u0_u6_n102 ) , .ZN( u2_u0_u6_n103 ) , .B1( u2_u0_u6_n160 ) , .A2( u2_u0_u6_n161 ) );
  NAND2_X1 u2_u0_u6_U60 (.ZN( u2_u0_u6_n113 ) , .A1( u2_u0_u6_n96 ) , .A2( u2_u0_u6_n98 ) );
  NOR2_X1 u2_u0_u6_U61 (.A2( u2_u0_X_40 ) , .A1( u2_u0_X_41 ) , .ZN( u2_u0_u6_n126 ) );
  NOR2_X1 u2_u0_u6_U62 (.A2( u2_u0_X_39 ) , .A1( u2_u0_X_42 ) , .ZN( u2_u0_u6_n92 ) );
  NOR2_X1 u2_u0_u6_U63 (.A2( u2_u0_X_39 ) , .A1( u2_u0_u6_n156 ) , .ZN( u2_u0_u6_n97 ) );
  NOR2_X1 u2_u0_u6_U64 (.A2( u2_u0_X_38 ) , .A1( u2_u0_u6_n165 ) , .ZN( u2_u0_u6_n95 ) );
  NOR2_X1 u2_u0_u6_U65 (.A2( u2_u0_X_41 ) , .ZN( u2_u0_u6_n111 ) , .A1( u2_u0_u6_n157 ) );
  NOR2_X1 u2_u0_u6_U66 (.A2( u2_u0_X_37 ) , .A1( u2_u0_u6_n162 ) , .ZN( u2_u0_u6_n94 ) );
  NOR2_X1 u2_u0_u6_U67 (.A2( u2_u0_X_37 ) , .A1( u2_u0_X_38 ) , .ZN( u2_u0_u6_n91 ) );
  NAND2_X1 u2_u0_u6_U68 (.A1( u2_u0_X_41 ) , .ZN( u2_u0_u6_n144 ) , .A2( u2_u0_u6_n157 ) );
  NAND2_X1 u2_u0_u6_U69 (.A2( u2_u0_X_40 ) , .A1( u2_u0_X_41 ) , .ZN( u2_u0_u6_n139 ) );
  NOR2_X1 u2_u0_u6_U7 (.A1( u2_u0_u6_n118 ) , .ZN( u2_u0_u6_n143 ) , .A2( u2_u0_u6_n168 ) );
  AND2_X1 u2_u0_u6_U70 (.A1( u2_u0_X_39 ) , .A2( u2_u0_u6_n156 ) , .ZN( u2_u0_u6_n96 ) );
  AND2_X1 u2_u0_u6_U71 (.A1( u2_u0_X_39 ) , .A2( u2_u0_X_42 ) , .ZN( u2_u0_u6_n99 ) );
  INV_X1 u2_u0_u6_U72 (.A( u2_u0_X_40 ) , .ZN( u2_u0_u6_n157 ) );
  INV_X1 u2_u0_u6_U73 (.A( u2_u0_X_37 ) , .ZN( u2_u0_u6_n165 ) );
  INV_X1 u2_u0_u6_U74 (.A( u2_u0_X_38 ) , .ZN( u2_u0_u6_n162 ) );
  INV_X1 u2_u0_u6_U75 (.A( u2_u0_X_42 ) , .ZN( u2_u0_u6_n156 ) );
  NAND4_X1 u2_u0_u6_U76 (.ZN( u2_out0_32 ) , .A4( u2_u0_u6_n103 ) , .A3( u2_u0_u6_n104 ) , .A2( u2_u0_u6_n105 ) , .A1( u2_u0_u6_n106 ) );
  AOI22_X1 u2_u0_u6_U77 (.ZN( u2_u0_u6_n105 ) , .A2( u2_u0_u6_n108 ) , .A1( u2_u0_u6_n118 ) , .B2( u2_u0_u6_n126 ) , .B1( u2_u0_u6_n171 ) );
  AOI22_X1 u2_u0_u6_U78 (.ZN( u2_u0_u6_n104 ) , .A1( u2_u0_u6_n111 ) , .B1( u2_u0_u6_n124 ) , .B2( u2_u0_u6_n151 ) , .A2( u2_u0_u6_n93 ) );
  NAND4_X1 u2_u0_u6_U79 (.ZN( u2_out0_12 ) , .A4( u2_u0_u6_n114 ) , .A3( u2_u0_u6_n115 ) , .A2( u2_u0_u6_n116 ) , .A1( u2_u0_u6_n117 ) );
  OAI21_X1 u2_u0_u6_U8 (.A( u2_u0_u6_n159 ) , .B1( u2_u0_u6_n169 ) , .B2( u2_u0_u6_n173 ) , .ZN( u2_u0_u6_n90 ) );
  OAI22_X1 u2_u0_u6_U80 (.B2( u2_u0_u6_n111 ) , .ZN( u2_u0_u6_n116 ) , .B1( u2_u0_u6_n126 ) , .A2( u2_u0_u6_n164 ) , .A1( u2_u0_u6_n167 ) );
  OAI21_X1 u2_u0_u6_U81 (.A( u2_u0_u6_n108 ) , .ZN( u2_u0_u6_n117 ) , .B2( u2_u0_u6_n141 ) , .B1( u2_u0_u6_n163 ) );
  OAI211_X1 u2_u0_u6_U82 (.ZN( u2_out0_7 ) , .B( u2_u0_u6_n153 ) , .C2( u2_u0_u6_n154 ) , .C1( u2_u0_u6_n155 ) , .A( u2_u0_u6_n174 ) );
  NOR3_X1 u2_u0_u6_U83 (.A1( u2_u0_u6_n141 ) , .ZN( u2_u0_u6_n154 ) , .A3( u2_u0_u6_n164 ) , .A2( u2_u0_u6_n171 ) );
  AOI211_X1 u2_u0_u6_U84 (.B( u2_u0_u6_n149 ) , .A( u2_u0_u6_n150 ) , .C2( u2_u0_u6_n151 ) , .C1( u2_u0_u6_n152 ) , .ZN( u2_u0_u6_n153 ) );
  OAI211_X1 u2_u0_u6_U85 (.ZN( u2_out0_22 ) , .B( u2_u0_u6_n137 ) , .A( u2_u0_u6_n138 ) , .C2( u2_u0_u6_n139 ) , .C1( u2_u0_u6_n140 ) );
  AOI22_X1 u2_u0_u6_U86 (.B1( u2_u0_u6_n124 ) , .A2( u2_u0_u6_n125 ) , .A1( u2_u0_u6_n126 ) , .ZN( u2_u0_u6_n138 ) , .B2( u2_u0_u6_n161 ) );
  AND4_X1 u2_u0_u6_U87 (.A3( u2_u0_u6_n119 ) , .A1( u2_u0_u6_n120 ) , .A4( u2_u0_u6_n129 ) , .ZN( u2_u0_u6_n140 ) , .A2( u2_u0_u6_n143 ) );
  NAND3_X1 u2_u0_u6_U88 (.A2( u2_u0_u6_n123 ) , .ZN( u2_u0_u6_n125 ) , .A1( u2_u0_u6_n130 ) , .A3( u2_u0_u6_n131 ) );
  NAND3_X1 u2_u0_u6_U89 (.A3( u2_u0_u6_n133 ) , .ZN( u2_u0_u6_n141 ) , .A1( u2_u0_u6_n145 ) , .A2( u2_u0_u6_n148 ) );
  INV_X1 u2_u0_u6_U9 (.ZN( u2_u0_u6_n172 ) , .A( u2_u0_u6_n88 ) );
  NAND3_X1 u2_u0_u6_U90 (.ZN( u2_u0_u6_n101 ) , .A3( u2_u0_u6_n107 ) , .A2( u2_u0_u6_n121 ) , .A1( u2_u0_u6_n127 ) );
  NAND3_X1 u2_u0_u6_U91 (.ZN( u2_u0_u6_n102 ) , .A3( u2_u0_u6_n130 ) , .A2( u2_u0_u6_n145 ) , .A1( u2_u0_u6_n166 ) );
  NAND3_X1 u2_u0_u6_U92 (.A3( u2_u0_u6_n113 ) , .A1( u2_u0_u6_n119 ) , .A2( u2_u0_u6_n123 ) , .ZN( u2_u0_u6_n93 ) );
  NAND3_X1 u2_u0_u6_U93 (.ZN( u2_u0_u6_n142 ) , .A2( u2_u0_u6_n172 ) , .A3( u2_u0_u6_n89 ) , .A1( u2_u0_u6_n90 ) );
  INV_X1 u2_u0_u7_U10 (.A( u2_u0_u7_n133 ) , .ZN( u2_u0_u7_n176 ) );
  OAI221_X1 u2_u0_u7_U11 (.C1( u2_u0_u7_n101 ) , .C2( u2_u0_u7_n147 ) , .ZN( u2_u0_u7_n155 ) , .B2( u2_u0_u7_n162 ) , .A( u2_u0_u7_n91 ) , .B1( u2_u0_u7_n92 ) );
  AND3_X1 u2_u0_u7_U12 (.A3( u2_u0_u7_n110 ) , .A2( u2_u0_u7_n127 ) , .A1( u2_u0_u7_n132 ) , .ZN( u2_u0_u7_n92 ) );
  OAI21_X1 u2_u0_u7_U13 (.A( u2_u0_u7_n161 ) , .B1( u2_u0_u7_n168 ) , .B2( u2_u0_u7_n173 ) , .ZN( u2_u0_u7_n91 ) );
  AOI211_X1 u2_u0_u7_U14 (.A( u2_u0_u7_n117 ) , .ZN( u2_u0_u7_n118 ) , .C2( u2_u0_u7_n126 ) , .C1( u2_u0_u7_n177 ) , .B( u2_u0_u7_n180 ) );
  OAI22_X1 u2_u0_u7_U15 (.B1( u2_u0_u7_n115 ) , .ZN( u2_u0_u7_n117 ) , .A2( u2_u0_u7_n133 ) , .A1( u2_u0_u7_n137 ) , .B2( u2_u0_u7_n162 ) );
  INV_X1 u2_u0_u7_U16 (.A( u2_u0_u7_n116 ) , .ZN( u2_u0_u7_n180 ) );
  NOR3_X1 u2_u0_u7_U17 (.ZN( u2_u0_u7_n115 ) , .A3( u2_u0_u7_n145 ) , .A2( u2_u0_u7_n168 ) , .A1( u2_u0_u7_n169 ) );
  NOR3_X1 u2_u0_u7_U18 (.A2( u2_u0_u7_n134 ) , .A1( u2_u0_u7_n135 ) , .ZN( u2_u0_u7_n136 ) , .A3( u2_u0_u7_n171 ) );
  NOR2_X1 u2_u0_u7_U19 (.A1( u2_u0_u7_n130 ) , .A2( u2_u0_u7_n134 ) , .ZN( u2_u0_u7_n153 ) );
  INV_X1 u2_u0_u7_U20 (.A( u2_u0_u7_n101 ) , .ZN( u2_u0_u7_n165 ) );
  NOR2_X1 u2_u0_u7_U21 (.ZN( u2_u0_u7_n111 ) , .A2( u2_u0_u7_n134 ) , .A1( u2_u0_u7_n169 ) );
  AOI21_X1 u2_u0_u7_U22 (.ZN( u2_u0_u7_n104 ) , .B2( u2_u0_u7_n112 ) , .B1( u2_u0_u7_n127 ) , .A( u2_u0_u7_n164 ) );
  AOI21_X1 u2_u0_u7_U23 (.ZN( u2_u0_u7_n106 ) , .B1( u2_u0_u7_n133 ) , .B2( u2_u0_u7_n146 ) , .A( u2_u0_u7_n162 ) );
  AOI21_X1 u2_u0_u7_U24 (.A( u2_u0_u7_n101 ) , .ZN( u2_u0_u7_n107 ) , .B2( u2_u0_u7_n128 ) , .B1( u2_u0_u7_n175 ) );
  INV_X1 u2_u0_u7_U25 (.A( u2_u0_u7_n138 ) , .ZN( u2_u0_u7_n171 ) );
  INV_X1 u2_u0_u7_U26 (.A( u2_u0_u7_n131 ) , .ZN( u2_u0_u7_n177 ) );
  INV_X1 u2_u0_u7_U27 (.A( u2_u0_u7_n110 ) , .ZN( u2_u0_u7_n174 ) );
  NAND2_X1 u2_u0_u7_U28 (.A1( u2_u0_u7_n129 ) , .A2( u2_u0_u7_n132 ) , .ZN( u2_u0_u7_n149 ) );
  NAND2_X1 u2_u0_u7_U29 (.A1( u2_u0_u7_n113 ) , .A2( u2_u0_u7_n124 ) , .ZN( u2_u0_u7_n130 ) );
  OAI21_X1 u2_u0_u7_U3 (.ZN( u2_u0_u7_n159 ) , .A( u2_u0_u7_n165 ) , .B2( u2_u0_u7_n171 ) , .B1( u2_u0_u7_n174 ) );
  INV_X1 u2_u0_u7_U30 (.A( u2_u0_u7_n112 ) , .ZN( u2_u0_u7_n173 ) );
  INV_X1 u2_u0_u7_U31 (.A( u2_u0_u7_n128 ) , .ZN( u2_u0_u7_n168 ) );
  INV_X1 u2_u0_u7_U32 (.A( u2_u0_u7_n148 ) , .ZN( u2_u0_u7_n169 ) );
  INV_X1 u2_u0_u7_U33 (.A( u2_u0_u7_n127 ) , .ZN( u2_u0_u7_n179 ) );
  NOR2_X1 u2_u0_u7_U34 (.ZN( u2_u0_u7_n101 ) , .A2( u2_u0_u7_n150 ) , .A1( u2_u0_u7_n156 ) );
  AOI211_X1 u2_u0_u7_U35 (.B( u2_u0_u7_n139 ) , .A( u2_u0_u7_n140 ) , .C2( u2_u0_u7_n141 ) , .ZN( u2_u0_u7_n142 ) , .C1( u2_u0_u7_n156 ) );
  NAND4_X1 u2_u0_u7_U36 (.A3( u2_u0_u7_n127 ) , .A2( u2_u0_u7_n128 ) , .A1( u2_u0_u7_n129 ) , .ZN( u2_u0_u7_n141 ) , .A4( u2_u0_u7_n147 ) );
  AOI21_X1 u2_u0_u7_U37 (.A( u2_u0_u7_n137 ) , .B1( u2_u0_u7_n138 ) , .ZN( u2_u0_u7_n139 ) , .B2( u2_u0_u7_n146 ) );
  OAI22_X1 u2_u0_u7_U38 (.B1( u2_u0_u7_n136 ) , .ZN( u2_u0_u7_n140 ) , .A1( u2_u0_u7_n153 ) , .B2( u2_u0_u7_n162 ) , .A2( u2_u0_u7_n164 ) );
  AOI211_X1 u2_u0_u7_U39 (.B( u2_u0_u7_n154 ) , .A( u2_u0_u7_n155 ) , .C1( u2_u0_u7_n156 ) , .ZN( u2_u0_u7_n157 ) , .C2( u2_u0_u7_n172 ) );
  INV_X1 u2_u0_u7_U4 (.A( u2_u0_u7_n111 ) , .ZN( u2_u0_u7_n170 ) );
  INV_X1 u2_u0_u7_U40 (.A( u2_u0_u7_n153 ) , .ZN( u2_u0_u7_n172 ) );
  INV_X1 u2_u0_u7_U41 (.A( u2_u0_u7_n125 ) , .ZN( u2_u0_u7_n161 ) );
  NAND2_X1 u2_u0_u7_U42 (.A2( u2_u0_u7_n102 ) , .A1( u2_u0_u7_n103 ) , .ZN( u2_u0_u7_n133 ) );
  NAND2_X1 u2_u0_u7_U43 (.A1( u2_u0_u7_n103 ) , .ZN( u2_u0_u7_n127 ) , .A2( u2_u0_u7_n99 ) );
  AOI21_X1 u2_u0_u7_U44 (.ZN( u2_u0_u7_n123 ) , .B1( u2_u0_u7_n165 ) , .B2( u2_u0_u7_n177 ) , .A( u2_u0_u7_n97 ) );
  AOI21_X1 u2_u0_u7_U45 (.B2( u2_u0_u7_n113 ) , .B1( u2_u0_u7_n124 ) , .A( u2_u0_u7_n125 ) , .ZN( u2_u0_u7_n97 ) );
  INV_X1 u2_u0_u7_U46 (.A( u2_u0_u7_n152 ) , .ZN( u2_u0_u7_n162 ) );
  AND2_X1 u2_u0_u7_U47 (.ZN( u2_u0_u7_n145 ) , .A2( u2_u0_u7_n98 ) , .A1( u2_u0_u7_n99 ) );
  NOR2_X1 u2_u0_u7_U48 (.ZN( u2_u0_u7_n137 ) , .A1( u2_u0_u7_n150 ) , .A2( u2_u0_u7_n161 ) );
  AOI21_X1 u2_u0_u7_U49 (.ZN( u2_u0_u7_n105 ) , .B2( u2_u0_u7_n110 ) , .A( u2_u0_u7_n125 ) , .B1( u2_u0_u7_n147 ) );
  INV_X1 u2_u0_u7_U5 (.A( u2_u0_u7_n154 ) , .ZN( u2_u0_u7_n178 ) );
  NAND2_X1 u2_u0_u7_U50 (.A2( u2_u0_u7_n103 ) , .ZN( u2_u0_u7_n147 ) , .A1( u2_u0_u7_n93 ) );
  NAND2_X1 u2_u0_u7_U51 (.ZN( u2_u0_u7_n146 ) , .A1( u2_u0_u7_n95 ) , .A2( u2_u0_u7_n98 ) );
  OR2_X1 u2_u0_u7_U52 (.ZN( u2_u0_u7_n126 ) , .A2( u2_u0_u7_n152 ) , .A1( u2_u0_u7_n156 ) );
  NAND2_X1 u2_u0_u7_U53 (.ZN( u2_u0_u7_n112 ) , .A2( u2_u0_u7_n96 ) , .A1( u2_u0_u7_n99 ) );
  NAND2_X1 u2_u0_u7_U54 (.A2( u2_u0_u7_n102 ) , .ZN( u2_u0_u7_n128 ) , .A1( u2_u0_u7_n98 ) );
  NAND2_X1 u2_u0_u7_U55 (.A1( u2_u0_u7_n100 ) , .ZN( u2_u0_u7_n113 ) , .A2( u2_u0_u7_n93 ) );
  NAND2_X1 u2_u0_u7_U56 (.ZN( u2_u0_u7_n110 ) , .A1( u2_u0_u7_n95 ) , .A2( u2_u0_u7_n96 ) );
  INV_X1 u2_u0_u7_U57 (.A( u2_u0_u7_n150 ) , .ZN( u2_u0_u7_n164 ) );
  AND2_X1 u2_u0_u7_U58 (.ZN( u2_u0_u7_n134 ) , .A1( u2_u0_u7_n93 ) , .A2( u2_u0_u7_n98 ) );
  NAND2_X1 u2_u0_u7_U59 (.A2( u2_u0_u7_n103 ) , .ZN( u2_u0_u7_n131 ) , .A1( u2_u0_u7_n95 ) );
  INV_X1 u2_u0_u7_U6 (.A( u2_u0_u7_n149 ) , .ZN( u2_u0_u7_n175 ) );
  NAND2_X1 u2_u0_u7_U60 (.A2( u2_u0_u7_n102 ) , .ZN( u2_u0_u7_n124 ) , .A1( u2_u0_u7_n96 ) );
  NAND2_X1 u2_u0_u7_U61 (.A1( u2_u0_u7_n100 ) , .A2( u2_u0_u7_n102 ) , .ZN( u2_u0_u7_n129 ) );
  NAND2_X1 u2_u0_u7_U62 (.A1( u2_u0_u7_n100 ) , .ZN( u2_u0_u7_n138 ) , .A2( u2_u0_u7_n99 ) );
  NAND2_X1 u2_u0_u7_U63 (.ZN( u2_u0_u7_n132 ) , .A1( u2_u0_u7_n93 ) , .A2( u2_u0_u7_n96 ) );
  NAND2_X1 u2_u0_u7_U64 (.A1( u2_u0_u7_n100 ) , .ZN( u2_u0_u7_n148 ) , .A2( u2_u0_u7_n95 ) );
  AOI22_X1 u2_u0_u7_U65 (.A2( u2_u0_u7_n114 ) , .ZN( u2_u0_u7_n119 ) , .B1( u2_u0_u7_n130 ) , .A1( u2_u0_u7_n156 ) , .B2( u2_u0_u7_n165 ) );
  NAND2_X1 u2_u0_u7_U66 (.A2( u2_u0_u7_n112 ) , .ZN( u2_u0_u7_n114 ) , .A1( u2_u0_u7_n175 ) );
  NOR2_X1 u2_u0_u7_U67 (.A2( u2_u0_X_47 ) , .ZN( u2_u0_u7_n150 ) , .A1( u2_u0_u7_n163 ) );
  NOR2_X1 u2_u0_u7_U68 (.A2( u2_u0_X_48 ) , .A1( u2_u0_u7_n166 ) , .ZN( u2_u0_u7_n95 ) );
  NOR2_X1 u2_u0_u7_U69 (.A2( u2_u0_X_45 ) , .A1( u2_u0_X_48 ) , .ZN( u2_u0_u7_n99 ) );
  AOI211_X1 u2_u0_u7_U7 (.ZN( u2_u0_u7_n116 ) , .A( u2_u0_u7_n155 ) , .C1( u2_u0_u7_n161 ) , .C2( u2_u0_u7_n171 ) , .B( u2_u0_u7_n94 ) );
  NOR2_X1 u2_u0_u7_U70 (.A2( u2_u0_X_44 ) , .A1( u2_u0_u7_n167 ) , .ZN( u2_u0_u7_n98 ) );
  NOR2_X1 u2_u0_u7_U71 (.A2( u2_u0_X_46 ) , .A1( u2_u0_X_47 ) , .ZN( u2_u0_u7_n152 ) );
  AND2_X1 u2_u0_u7_U72 (.A1( u2_u0_X_47 ) , .ZN( u2_u0_u7_n156 ) , .A2( u2_u0_u7_n163 ) );
  NAND2_X1 u2_u0_u7_U73 (.A2( u2_u0_X_46 ) , .A1( u2_u0_X_47 ) , .ZN( u2_u0_u7_n125 ) );
  AND2_X1 u2_u0_u7_U74 (.A2( u2_u0_X_45 ) , .A1( u2_u0_X_48 ) , .ZN( u2_u0_u7_n102 ) );
  AND2_X1 u2_u0_u7_U75 (.A2( u2_u0_X_43 ) , .A1( u2_u0_X_44 ) , .ZN( u2_u0_u7_n96 ) );
  AND2_X1 u2_u0_u7_U76 (.A1( u2_u0_X_44 ) , .ZN( u2_u0_u7_n100 ) , .A2( u2_u0_u7_n167 ) );
  AND2_X1 u2_u0_u7_U77 (.A1( u2_u0_X_48 ) , .A2( u2_u0_u7_n166 ) , .ZN( u2_u0_u7_n93 ) );
  INV_X1 u2_u0_u7_U78 (.A( u2_u0_X_46 ) , .ZN( u2_u0_u7_n163 ) );
  INV_X1 u2_u0_u7_U79 (.A( u2_u0_X_45 ) , .ZN( u2_u0_u7_n166 ) );
  OAI222_X1 u2_u0_u7_U8 (.C2( u2_u0_u7_n101 ) , .B2( u2_u0_u7_n111 ) , .A1( u2_u0_u7_n113 ) , .C1( u2_u0_u7_n146 ) , .A2( u2_u0_u7_n162 ) , .B1( u2_u0_u7_n164 ) , .ZN( u2_u0_u7_n94 ) );
  OAI21_X1 u2_u0_u7_U80 (.B1( u2_u0_u7_n145 ) , .ZN( u2_u0_u7_n160 ) , .A( u2_u0_u7_n161 ) , .B2( u2_u0_u7_n177 ) );
  AOI22_X1 u2_u0_u7_U81 (.B2( u2_u0_u7_n149 ) , .B1( u2_u0_u7_n150 ) , .A2( u2_u0_u7_n151 ) , .A1( u2_u0_u7_n152 ) , .ZN( u2_u0_u7_n158 ) );
  NAND4_X1 u2_u0_u7_U82 (.ZN( u2_out0_27 ) , .A4( u2_u0_u7_n118 ) , .A3( u2_u0_u7_n119 ) , .A2( u2_u0_u7_n120 ) , .A1( u2_u0_u7_n121 ) );
  OAI21_X1 u2_u0_u7_U83 (.ZN( u2_u0_u7_n121 ) , .B2( u2_u0_u7_n145 ) , .A( u2_u0_u7_n150 ) , .B1( u2_u0_u7_n174 ) );
  OAI21_X1 u2_u0_u7_U84 (.ZN( u2_u0_u7_n120 ) , .A( u2_u0_u7_n161 ) , .B2( u2_u0_u7_n170 ) , .B1( u2_u0_u7_n179 ) );
  NAND4_X1 u2_u0_u7_U85 (.ZN( u2_out0_15 ) , .A4( u2_u0_u7_n142 ) , .A3( u2_u0_u7_n143 ) , .A2( u2_u0_u7_n144 ) , .A1( u2_u0_u7_n178 ) );
  OR2_X1 u2_u0_u7_U86 (.A2( u2_u0_u7_n125 ) , .A1( u2_u0_u7_n129 ) , .ZN( u2_u0_u7_n144 ) );
  AOI22_X1 u2_u0_u7_U87 (.A2( u2_u0_u7_n126 ) , .ZN( u2_u0_u7_n143 ) , .B2( u2_u0_u7_n165 ) , .B1( u2_u0_u7_n173 ) , .A1( u2_u0_u7_n174 ) );
  NAND4_X1 u2_u0_u7_U88 (.ZN( u2_out0_5 ) , .A4( u2_u0_u7_n108 ) , .A3( u2_u0_u7_n109 ) , .A1( u2_u0_u7_n116 ) , .A2( u2_u0_u7_n123 ) );
  AOI22_X1 u2_u0_u7_U89 (.ZN( u2_u0_u7_n109 ) , .A2( u2_u0_u7_n126 ) , .B2( u2_u0_u7_n145 ) , .B1( u2_u0_u7_n156 ) , .A1( u2_u0_u7_n171 ) );
  AOI222_X1 u2_u0_u7_U9 (.ZN( u2_u0_u7_n122 ) , .C2( u2_u0_u7_n126 ) , .C1( u2_u0_u7_n145 ) , .B1( u2_u0_u7_n161 ) , .A2( u2_u0_u7_n165 ) , .B2( u2_u0_u7_n170 ) , .A1( u2_u0_u7_n176 ) );
  NOR4_X1 u2_u0_u7_U90 (.A4( u2_u0_u7_n104 ) , .A3( u2_u0_u7_n105 ) , .A2( u2_u0_u7_n106 ) , .A1( u2_u0_u7_n107 ) , .ZN( u2_u0_u7_n108 ) );
  NAND4_X1 u2_u0_u7_U91 (.ZN( u2_out0_21 ) , .A4( u2_u0_u7_n157 ) , .A3( u2_u0_u7_n158 ) , .A2( u2_u0_u7_n159 ) , .A1( u2_u0_u7_n160 ) );
  OAI211_X1 u2_u0_u7_U92 (.B( u2_u0_u7_n122 ) , .A( u2_u0_u7_n123 ) , .C2( u2_u0_u7_n124 ) , .ZN( u2_u0_u7_n154 ) , .C1( u2_u0_u7_n162 ) );
  NOR2_X1 u2_u0_u7_U93 (.A2( u2_u0_X_43 ) , .A1( u2_u0_X_44 ) , .ZN( u2_u0_u7_n103 ) );
  INV_X1 u2_u0_u7_U94 (.A( u2_u0_X_43 ) , .ZN( u2_u0_u7_n167 ) );
  NAND3_X1 u2_u0_u7_U95 (.A3( u2_u0_u7_n146 ) , .A2( u2_u0_u7_n147 ) , .A1( u2_u0_u7_n148 ) , .ZN( u2_u0_u7_n151 ) );
  NAND3_X1 u2_u0_u7_U96 (.A3( u2_u0_u7_n131 ) , .A2( u2_u0_u7_n132 ) , .A1( u2_u0_u7_n133 ) , .ZN( u2_u0_u7_n135 ) );
  XOR2_X1 u2_u14_U20 (.B( u2_K15_36 ) , .A( u2_R13_25 ) , .Z( u2_u14_X_36 ) );
  XOR2_X1 u2_u14_U21 (.B( u2_K15_35 ) , .A( u2_R13_24 ) , .Z( u2_u14_X_35 ) );
  XOR2_X1 u2_u14_U23 (.B( u2_K15_33 ) , .A( u2_R13_22 ) , .Z( u2_u14_X_33 ) );
  XOR2_X1 u2_u14_U25 (.B( u2_K15_31 ) , .A( u2_R13_20 ) , .Z( u2_u14_X_31 ) );
  XOR2_X1 u2_u14_U28 (.B( u2_K15_29 ) , .A( u2_R13_20 ) , .Z( u2_u14_X_29 ) );
  XOR2_X1 u2_u14_U30 (.B( u2_K15_27 ) , .A( u2_R13_18 ) , .Z( u2_u14_X_27 ) );
  XOR2_X1 u2_u14_U31 (.B( u2_K15_26 ) , .A( u2_R13_17 ) , .Z( u2_u14_X_26 ) );
  OAI22_X1 u2_u14_u4_U10 (.B2( u2_u14_u4_n135 ) , .ZN( u2_u14_u4_n137 ) , .B1( u2_u14_u4_n153 ) , .A1( u2_u14_u4_n155 ) , .A2( u2_u14_u4_n171 ) );
  AND3_X1 u2_u14_u4_U11 (.A2( u2_u14_u4_n134 ) , .ZN( u2_u14_u4_n135 ) , .A3( u2_u14_u4_n145 ) , .A1( u2_u14_u4_n157 ) );
  NAND2_X1 u2_u14_u4_U12 (.ZN( u2_u14_u4_n132 ) , .A2( u2_u14_u4_n170 ) , .A1( u2_u14_u4_n173 ) );
  AOI21_X1 u2_u14_u4_U13 (.B2( u2_u14_u4_n160 ) , .B1( u2_u14_u4_n161 ) , .ZN( u2_u14_u4_n162 ) , .A( u2_u14_u4_n170 ) );
  AOI21_X1 u2_u14_u4_U14 (.ZN( u2_u14_u4_n107 ) , .B2( u2_u14_u4_n143 ) , .A( u2_u14_u4_n174 ) , .B1( u2_u14_u4_n184 ) );
  AOI21_X1 u2_u14_u4_U15 (.B2( u2_u14_u4_n158 ) , .B1( u2_u14_u4_n159 ) , .ZN( u2_u14_u4_n163 ) , .A( u2_u14_u4_n174 ) );
  AOI21_X1 u2_u14_u4_U16 (.A( u2_u14_u4_n153 ) , .B2( u2_u14_u4_n154 ) , .B1( u2_u14_u4_n155 ) , .ZN( u2_u14_u4_n165 ) );
  AOI21_X1 u2_u14_u4_U17 (.A( u2_u14_u4_n156 ) , .B2( u2_u14_u4_n157 ) , .ZN( u2_u14_u4_n164 ) , .B1( u2_u14_u4_n184 ) );
  INV_X1 u2_u14_u4_U18 (.A( u2_u14_u4_n138 ) , .ZN( u2_u14_u4_n170 ) );
  AND2_X1 u2_u14_u4_U19 (.A2( u2_u14_u4_n120 ) , .ZN( u2_u14_u4_n155 ) , .A1( u2_u14_u4_n160 ) );
  INV_X1 u2_u14_u4_U20 (.A( u2_u14_u4_n156 ) , .ZN( u2_u14_u4_n175 ) );
  NAND2_X1 u2_u14_u4_U21 (.A2( u2_u14_u4_n118 ) , .ZN( u2_u14_u4_n131 ) , .A1( u2_u14_u4_n147 ) );
  NAND2_X1 u2_u14_u4_U22 (.A1( u2_u14_u4_n119 ) , .A2( u2_u14_u4_n120 ) , .ZN( u2_u14_u4_n130 ) );
  NAND2_X1 u2_u14_u4_U23 (.ZN( u2_u14_u4_n117 ) , .A2( u2_u14_u4_n118 ) , .A1( u2_u14_u4_n148 ) );
  NAND2_X1 u2_u14_u4_U24 (.ZN( u2_u14_u4_n129 ) , .A1( u2_u14_u4_n134 ) , .A2( u2_u14_u4_n148 ) );
  AND3_X1 u2_u14_u4_U25 (.A1( u2_u14_u4_n119 ) , .A2( u2_u14_u4_n143 ) , .A3( u2_u14_u4_n154 ) , .ZN( u2_u14_u4_n161 ) );
  AND2_X1 u2_u14_u4_U26 (.A1( u2_u14_u4_n145 ) , .A2( u2_u14_u4_n147 ) , .ZN( u2_u14_u4_n159 ) );
  OR3_X1 u2_u14_u4_U27 (.A3( u2_u14_u4_n114 ) , .A2( u2_u14_u4_n115 ) , .A1( u2_u14_u4_n116 ) , .ZN( u2_u14_u4_n136 ) );
  AOI21_X1 u2_u14_u4_U28 (.A( u2_u14_u4_n113 ) , .ZN( u2_u14_u4_n116 ) , .B2( u2_u14_u4_n173 ) , .B1( u2_u14_u4_n174 ) );
  AOI21_X1 u2_u14_u4_U29 (.ZN( u2_u14_u4_n115 ) , .B2( u2_u14_u4_n145 ) , .B1( u2_u14_u4_n146 ) , .A( u2_u14_u4_n156 ) );
  NOR2_X1 u2_u14_u4_U3 (.ZN( u2_u14_u4_n121 ) , .A1( u2_u14_u4_n181 ) , .A2( u2_u14_u4_n182 ) );
  OAI22_X1 u2_u14_u4_U30 (.ZN( u2_u14_u4_n114 ) , .A2( u2_u14_u4_n121 ) , .B1( u2_u14_u4_n160 ) , .B2( u2_u14_u4_n170 ) , .A1( u2_u14_u4_n171 ) );
  INV_X1 u2_u14_u4_U31 (.A( u2_u14_u4_n158 ) , .ZN( u2_u14_u4_n182 ) );
  INV_X1 u2_u14_u4_U32 (.ZN( u2_u14_u4_n181 ) , .A( u2_u14_u4_n96 ) );
  INV_X1 u2_u14_u4_U33 (.A( u2_u14_u4_n144 ) , .ZN( u2_u14_u4_n179 ) );
  INV_X1 u2_u14_u4_U34 (.A( u2_u14_u4_n157 ) , .ZN( u2_u14_u4_n178 ) );
  NAND2_X1 u2_u14_u4_U35 (.A2( u2_u14_u4_n154 ) , .A1( u2_u14_u4_n96 ) , .ZN( u2_u14_u4_n97 ) );
  INV_X1 u2_u14_u4_U36 (.ZN( u2_u14_u4_n186 ) , .A( u2_u14_u4_n95 ) );
  OAI221_X1 u2_u14_u4_U37 (.C1( u2_u14_u4_n134 ) , .B1( u2_u14_u4_n158 ) , .B2( u2_u14_u4_n171 ) , .C2( u2_u14_u4_n173 ) , .A( u2_u14_u4_n94 ) , .ZN( u2_u14_u4_n95 ) );
  AOI222_X1 u2_u14_u4_U38 (.B2( u2_u14_u4_n132 ) , .A1( u2_u14_u4_n138 ) , .C2( u2_u14_u4_n175 ) , .A2( u2_u14_u4_n179 ) , .C1( u2_u14_u4_n181 ) , .B1( u2_u14_u4_n185 ) , .ZN( u2_u14_u4_n94 ) );
  INV_X1 u2_u14_u4_U39 (.A( u2_u14_u4_n113 ) , .ZN( u2_u14_u4_n185 ) );
  INV_X1 u2_u14_u4_U4 (.A( u2_u14_u4_n117 ) , .ZN( u2_u14_u4_n184 ) );
  INV_X1 u2_u14_u4_U40 (.A( u2_u14_u4_n143 ) , .ZN( u2_u14_u4_n183 ) );
  NOR2_X1 u2_u14_u4_U41 (.ZN( u2_u14_u4_n138 ) , .A1( u2_u14_u4_n168 ) , .A2( u2_u14_u4_n169 ) );
  NOR2_X1 u2_u14_u4_U42 (.A1( u2_u14_u4_n150 ) , .A2( u2_u14_u4_n152 ) , .ZN( u2_u14_u4_n153 ) );
  NOR2_X1 u2_u14_u4_U43 (.A2( u2_u14_u4_n128 ) , .A1( u2_u14_u4_n138 ) , .ZN( u2_u14_u4_n156 ) );
  AOI22_X1 u2_u14_u4_U44 (.B2( u2_u14_u4_n122 ) , .A1( u2_u14_u4_n123 ) , .ZN( u2_u14_u4_n124 ) , .B1( u2_u14_u4_n128 ) , .A2( u2_u14_u4_n172 ) );
  INV_X1 u2_u14_u4_U45 (.A( u2_u14_u4_n153 ) , .ZN( u2_u14_u4_n172 ) );
  NAND2_X1 u2_u14_u4_U46 (.A2( u2_u14_u4_n120 ) , .ZN( u2_u14_u4_n123 ) , .A1( u2_u14_u4_n161 ) );
  AOI22_X1 u2_u14_u4_U47 (.B2( u2_u14_u4_n132 ) , .A2( u2_u14_u4_n133 ) , .ZN( u2_u14_u4_n140 ) , .A1( u2_u14_u4_n150 ) , .B1( u2_u14_u4_n179 ) );
  NAND2_X1 u2_u14_u4_U48 (.ZN( u2_u14_u4_n133 ) , .A2( u2_u14_u4_n146 ) , .A1( u2_u14_u4_n154 ) );
  NAND2_X1 u2_u14_u4_U49 (.A1( u2_u14_u4_n103 ) , .ZN( u2_u14_u4_n154 ) , .A2( u2_u14_u4_n98 ) );
  NOR4_X1 u2_u14_u4_U5 (.A4( u2_u14_u4_n106 ) , .A3( u2_u14_u4_n107 ) , .A2( u2_u14_u4_n108 ) , .A1( u2_u14_u4_n109 ) , .ZN( u2_u14_u4_n110 ) );
  NAND2_X1 u2_u14_u4_U50 (.A1( u2_u14_u4_n101 ) , .ZN( u2_u14_u4_n158 ) , .A2( u2_u14_u4_n99 ) );
  AOI21_X1 u2_u14_u4_U51 (.ZN( u2_u14_u4_n127 ) , .A( u2_u14_u4_n136 ) , .B2( u2_u14_u4_n150 ) , .B1( u2_u14_u4_n180 ) );
  INV_X1 u2_u14_u4_U52 (.A( u2_u14_u4_n160 ) , .ZN( u2_u14_u4_n180 ) );
  NAND2_X1 u2_u14_u4_U53 (.A2( u2_u14_u4_n104 ) , .A1( u2_u14_u4_n105 ) , .ZN( u2_u14_u4_n146 ) );
  NAND2_X1 u2_u14_u4_U54 (.A2( u2_u14_u4_n101 ) , .A1( u2_u14_u4_n102 ) , .ZN( u2_u14_u4_n160 ) );
  NAND2_X1 u2_u14_u4_U55 (.ZN( u2_u14_u4_n134 ) , .A1( u2_u14_u4_n98 ) , .A2( u2_u14_u4_n99 ) );
  NAND2_X1 u2_u14_u4_U56 (.A1( u2_u14_u4_n103 ) , .A2( u2_u14_u4_n104 ) , .ZN( u2_u14_u4_n143 ) );
  NAND2_X1 u2_u14_u4_U57 (.A2( u2_u14_u4_n105 ) , .ZN( u2_u14_u4_n145 ) , .A1( u2_u14_u4_n98 ) );
  NAND2_X1 u2_u14_u4_U58 (.A1( u2_u14_u4_n100 ) , .A2( u2_u14_u4_n105 ) , .ZN( u2_u14_u4_n120 ) );
  NAND2_X1 u2_u14_u4_U59 (.A1( u2_u14_u4_n102 ) , .A2( u2_u14_u4_n104 ) , .ZN( u2_u14_u4_n148 ) );
  AOI21_X1 u2_u14_u4_U6 (.ZN( u2_u14_u4_n106 ) , .B2( u2_u14_u4_n146 ) , .B1( u2_u14_u4_n158 ) , .A( u2_u14_u4_n170 ) );
  NAND2_X1 u2_u14_u4_U60 (.A2( u2_u14_u4_n100 ) , .A1( u2_u14_u4_n103 ) , .ZN( u2_u14_u4_n157 ) );
  INV_X1 u2_u14_u4_U61 (.A( u2_u14_u4_n150 ) , .ZN( u2_u14_u4_n173 ) );
  INV_X1 u2_u14_u4_U62 (.A( u2_u14_u4_n152 ) , .ZN( u2_u14_u4_n171 ) );
  NAND2_X1 u2_u14_u4_U63 (.A1( u2_u14_u4_n100 ) , .ZN( u2_u14_u4_n118 ) , .A2( u2_u14_u4_n99 ) );
  NAND2_X1 u2_u14_u4_U64 (.A2( u2_u14_u4_n100 ) , .A1( u2_u14_u4_n102 ) , .ZN( u2_u14_u4_n144 ) );
  NAND2_X1 u2_u14_u4_U65 (.A2( u2_u14_u4_n101 ) , .A1( u2_u14_u4_n105 ) , .ZN( u2_u14_u4_n96 ) );
  INV_X1 u2_u14_u4_U66 (.A( u2_u14_u4_n128 ) , .ZN( u2_u14_u4_n174 ) );
  NAND2_X1 u2_u14_u4_U67 (.A2( u2_u14_u4_n102 ) , .ZN( u2_u14_u4_n119 ) , .A1( u2_u14_u4_n98 ) );
  NAND2_X1 u2_u14_u4_U68 (.A2( u2_u14_u4_n101 ) , .A1( u2_u14_u4_n103 ) , .ZN( u2_u14_u4_n147 ) );
  NAND2_X1 u2_u14_u4_U69 (.A2( u2_u14_u4_n104 ) , .ZN( u2_u14_u4_n113 ) , .A1( u2_u14_u4_n99 ) );
  AOI21_X1 u2_u14_u4_U7 (.ZN( u2_u14_u4_n108 ) , .B2( u2_u14_u4_n134 ) , .B1( u2_u14_u4_n155 ) , .A( u2_u14_u4_n156 ) );
  NOR2_X1 u2_u14_u4_U70 (.A2( u2_u14_X_28 ) , .ZN( u2_u14_u4_n150 ) , .A1( u2_u14_u4_n168 ) );
  NOR2_X1 u2_u14_u4_U71 (.A2( u2_u14_X_29 ) , .ZN( u2_u14_u4_n152 ) , .A1( u2_u14_u4_n169 ) );
  NOR2_X1 u2_u14_u4_U72 (.A2( u2_u14_X_30 ) , .ZN( u2_u14_u4_n105 ) , .A1( u2_u14_u4_n176 ) );
  NOR2_X1 u2_u14_u4_U73 (.A2( u2_u14_X_26 ) , .ZN( u2_u14_u4_n100 ) , .A1( u2_u14_u4_n177 ) );
  NOR2_X1 u2_u14_u4_U74 (.A2( u2_u14_X_28 ) , .A1( u2_u14_X_29 ) , .ZN( u2_u14_u4_n128 ) );
  NOR2_X1 u2_u14_u4_U75 (.A2( u2_u14_X_27 ) , .A1( u2_u14_X_30 ) , .ZN( u2_u14_u4_n102 ) );
  NOR2_X1 u2_u14_u4_U76 (.A2( u2_u14_X_25 ) , .A1( u2_u14_X_26 ) , .ZN( u2_u14_u4_n98 ) );
  AND2_X1 u2_u14_u4_U77 (.A2( u2_u14_X_25 ) , .A1( u2_u14_X_26 ) , .ZN( u2_u14_u4_n104 ) );
  AND2_X1 u2_u14_u4_U78 (.A1( u2_u14_X_30 ) , .A2( u2_u14_u4_n176 ) , .ZN( u2_u14_u4_n99 ) );
  AND2_X1 u2_u14_u4_U79 (.A1( u2_u14_X_26 ) , .ZN( u2_u14_u4_n101 ) , .A2( u2_u14_u4_n177 ) );
  AOI21_X1 u2_u14_u4_U8 (.ZN( u2_u14_u4_n109 ) , .A( u2_u14_u4_n153 ) , .B1( u2_u14_u4_n159 ) , .B2( u2_u14_u4_n184 ) );
  AND2_X1 u2_u14_u4_U80 (.A1( u2_u14_X_27 ) , .A2( u2_u14_X_30 ) , .ZN( u2_u14_u4_n103 ) );
  INV_X1 u2_u14_u4_U81 (.A( u2_u14_X_28 ) , .ZN( u2_u14_u4_n169 ) );
  INV_X1 u2_u14_u4_U82 (.A( u2_u14_X_29 ) , .ZN( u2_u14_u4_n168 ) );
  INV_X1 u2_u14_u4_U83 (.A( u2_u14_X_25 ) , .ZN( u2_u14_u4_n177 ) );
  INV_X1 u2_u14_u4_U84 (.A( u2_u14_X_27 ) , .ZN( u2_u14_u4_n176 ) );
  NAND4_X1 u2_u14_u4_U85 (.ZN( u2_out14_25 ) , .A4( u2_u14_u4_n139 ) , .A3( u2_u14_u4_n140 ) , .A2( u2_u14_u4_n141 ) , .A1( u2_u14_u4_n142 ) );
  OAI21_X1 u2_u14_u4_U86 (.A( u2_u14_u4_n128 ) , .B2( u2_u14_u4_n129 ) , .B1( u2_u14_u4_n130 ) , .ZN( u2_u14_u4_n142 ) );
  OAI21_X1 u2_u14_u4_U87 (.B2( u2_u14_u4_n131 ) , .ZN( u2_u14_u4_n141 ) , .A( u2_u14_u4_n175 ) , .B1( u2_u14_u4_n183 ) );
  NAND4_X1 u2_u14_u4_U88 (.ZN( u2_out14_14 ) , .A4( u2_u14_u4_n124 ) , .A3( u2_u14_u4_n125 ) , .A2( u2_u14_u4_n126 ) , .A1( u2_u14_u4_n127 ) );
  AOI22_X1 u2_u14_u4_U89 (.B2( u2_u14_u4_n117 ) , .ZN( u2_u14_u4_n126 ) , .A1( u2_u14_u4_n129 ) , .B1( u2_u14_u4_n152 ) , .A2( u2_u14_u4_n175 ) );
  AOI211_X1 u2_u14_u4_U9 (.B( u2_u14_u4_n136 ) , .A( u2_u14_u4_n137 ) , .C2( u2_u14_u4_n138 ) , .ZN( u2_u14_u4_n139 ) , .C1( u2_u14_u4_n182 ) );
  AOI22_X1 u2_u14_u4_U90 (.ZN( u2_u14_u4_n125 ) , .B2( u2_u14_u4_n131 ) , .A2( u2_u14_u4_n132 ) , .B1( u2_u14_u4_n138 ) , .A1( u2_u14_u4_n178 ) );
  NAND4_X1 u2_u14_u4_U91 (.ZN( u2_out14_8 ) , .A4( u2_u14_u4_n110 ) , .A3( u2_u14_u4_n111 ) , .A2( u2_u14_u4_n112 ) , .A1( u2_u14_u4_n186 ) );
  NAND2_X1 u2_u14_u4_U92 (.ZN( u2_u14_u4_n112 ) , .A2( u2_u14_u4_n130 ) , .A1( u2_u14_u4_n150 ) );
  AOI22_X1 u2_u14_u4_U93 (.ZN( u2_u14_u4_n111 ) , .B2( u2_u14_u4_n132 ) , .A1( u2_u14_u4_n152 ) , .B1( u2_u14_u4_n178 ) , .A2( u2_u14_u4_n97 ) );
  AOI22_X1 u2_u14_u4_U94 (.B2( u2_u14_u4_n149 ) , .B1( u2_u14_u4_n150 ) , .A2( u2_u14_u4_n151 ) , .A1( u2_u14_u4_n152 ) , .ZN( u2_u14_u4_n167 ) );
  NOR4_X1 u2_u14_u4_U95 (.A4( u2_u14_u4_n162 ) , .A3( u2_u14_u4_n163 ) , .A2( u2_u14_u4_n164 ) , .A1( u2_u14_u4_n165 ) , .ZN( u2_u14_u4_n166 ) );
  NAND3_X1 u2_u14_u4_U96 (.ZN( u2_out14_3 ) , .A3( u2_u14_u4_n166 ) , .A1( u2_u14_u4_n167 ) , .A2( u2_u14_u4_n186 ) );
  NAND3_X1 u2_u14_u4_U97 (.A3( u2_u14_u4_n146 ) , .A2( u2_u14_u4_n147 ) , .A1( u2_u14_u4_n148 ) , .ZN( u2_u14_u4_n149 ) );
  NAND3_X1 u2_u14_u4_U98 (.A3( u2_u14_u4_n143 ) , .A2( u2_u14_u4_n144 ) , .A1( u2_u14_u4_n145 ) , .ZN( u2_u14_u4_n151 ) );
  NAND3_X1 u2_u14_u4_U99 (.A3( u2_u14_u4_n121 ) , .ZN( u2_u14_u4_n122 ) , .A2( u2_u14_u4_n144 ) , .A1( u2_u14_u4_n154 ) );
  INV_X1 u2_u14_u5_U10 (.A( u2_u14_u5_n121 ) , .ZN( u2_u14_u5_n177 ) );
  NOR3_X1 u2_u14_u5_U100 (.A3( u2_u14_u5_n141 ) , .A1( u2_u14_u5_n142 ) , .ZN( u2_u14_u5_n143 ) , .A2( u2_u14_u5_n191 ) );
  NAND4_X1 u2_u14_u5_U101 (.ZN( u2_out14_4 ) , .A4( u2_u14_u5_n112 ) , .A2( u2_u14_u5_n113 ) , .A1( u2_u14_u5_n114 ) , .A3( u2_u14_u5_n195 ) );
  AOI211_X1 u2_u14_u5_U102 (.A( u2_u14_u5_n110 ) , .C1( u2_u14_u5_n111 ) , .ZN( u2_u14_u5_n112 ) , .B( u2_u14_u5_n118 ) , .C2( u2_u14_u5_n177 ) );
  AOI222_X1 u2_u14_u5_U103 (.ZN( u2_u14_u5_n113 ) , .A1( u2_u14_u5_n131 ) , .C1( u2_u14_u5_n148 ) , .B2( u2_u14_u5_n174 ) , .C2( u2_u14_u5_n178 ) , .A2( u2_u14_u5_n179 ) , .B1( u2_u14_u5_n99 ) );
  NAND3_X1 u2_u14_u5_U104 (.A2( u2_u14_u5_n154 ) , .A3( u2_u14_u5_n158 ) , .A1( u2_u14_u5_n161 ) , .ZN( u2_u14_u5_n99 ) );
  NOR2_X1 u2_u14_u5_U11 (.ZN( u2_u14_u5_n160 ) , .A2( u2_u14_u5_n173 ) , .A1( u2_u14_u5_n177 ) );
  INV_X1 u2_u14_u5_U12 (.A( u2_u14_u5_n150 ) , .ZN( u2_u14_u5_n174 ) );
  AOI21_X1 u2_u14_u5_U13 (.A( u2_u14_u5_n160 ) , .B2( u2_u14_u5_n161 ) , .ZN( u2_u14_u5_n162 ) , .B1( u2_u14_u5_n192 ) );
  INV_X1 u2_u14_u5_U14 (.A( u2_u14_u5_n159 ) , .ZN( u2_u14_u5_n192 ) );
  AOI21_X1 u2_u14_u5_U15 (.A( u2_u14_u5_n156 ) , .B2( u2_u14_u5_n157 ) , .B1( u2_u14_u5_n158 ) , .ZN( u2_u14_u5_n163 ) );
  AOI21_X1 u2_u14_u5_U16 (.B2( u2_u14_u5_n139 ) , .B1( u2_u14_u5_n140 ) , .ZN( u2_u14_u5_n141 ) , .A( u2_u14_u5_n150 ) );
  OAI21_X1 u2_u14_u5_U17 (.A( u2_u14_u5_n133 ) , .B2( u2_u14_u5_n134 ) , .B1( u2_u14_u5_n135 ) , .ZN( u2_u14_u5_n142 ) );
  OAI21_X1 u2_u14_u5_U18 (.ZN( u2_u14_u5_n133 ) , .B2( u2_u14_u5_n147 ) , .A( u2_u14_u5_n173 ) , .B1( u2_u14_u5_n188 ) );
  NAND2_X1 u2_u14_u5_U19 (.A2( u2_u14_u5_n119 ) , .A1( u2_u14_u5_n123 ) , .ZN( u2_u14_u5_n137 ) );
  INV_X1 u2_u14_u5_U20 (.A( u2_u14_u5_n155 ) , .ZN( u2_u14_u5_n194 ) );
  NAND2_X1 u2_u14_u5_U21 (.A1( u2_u14_u5_n121 ) , .ZN( u2_u14_u5_n132 ) , .A2( u2_u14_u5_n172 ) );
  NAND2_X1 u2_u14_u5_U22 (.A2( u2_u14_u5_n122 ) , .ZN( u2_u14_u5_n136 ) , .A1( u2_u14_u5_n154 ) );
  NAND2_X1 u2_u14_u5_U23 (.A2( u2_u14_u5_n119 ) , .A1( u2_u14_u5_n120 ) , .ZN( u2_u14_u5_n159 ) );
  INV_X1 u2_u14_u5_U24 (.A( u2_u14_u5_n156 ) , .ZN( u2_u14_u5_n175 ) );
  INV_X1 u2_u14_u5_U25 (.A( u2_u14_u5_n158 ) , .ZN( u2_u14_u5_n188 ) );
  INV_X1 u2_u14_u5_U26 (.A( u2_u14_u5_n152 ) , .ZN( u2_u14_u5_n179 ) );
  INV_X1 u2_u14_u5_U27 (.A( u2_u14_u5_n140 ) , .ZN( u2_u14_u5_n182 ) );
  INV_X1 u2_u14_u5_U28 (.A( u2_u14_u5_n151 ) , .ZN( u2_u14_u5_n183 ) );
  INV_X1 u2_u14_u5_U29 (.A( u2_u14_u5_n123 ) , .ZN( u2_u14_u5_n185 ) );
  NOR2_X1 u2_u14_u5_U3 (.ZN( u2_u14_u5_n134 ) , .A1( u2_u14_u5_n183 ) , .A2( u2_u14_u5_n190 ) );
  INV_X1 u2_u14_u5_U30 (.A( u2_u14_u5_n161 ) , .ZN( u2_u14_u5_n184 ) );
  INV_X1 u2_u14_u5_U31 (.A( u2_u14_u5_n139 ) , .ZN( u2_u14_u5_n189 ) );
  INV_X1 u2_u14_u5_U32 (.A( u2_u14_u5_n157 ) , .ZN( u2_u14_u5_n190 ) );
  INV_X1 u2_u14_u5_U33 (.A( u2_u14_u5_n120 ) , .ZN( u2_u14_u5_n193 ) );
  NAND2_X1 u2_u14_u5_U34 (.ZN( u2_u14_u5_n111 ) , .A1( u2_u14_u5_n140 ) , .A2( u2_u14_u5_n155 ) );
  INV_X1 u2_u14_u5_U35 (.A( u2_u14_u5_n117 ) , .ZN( u2_u14_u5_n196 ) );
  OAI221_X1 u2_u14_u5_U36 (.A( u2_u14_u5_n116 ) , .ZN( u2_u14_u5_n117 ) , .B2( u2_u14_u5_n119 ) , .C1( u2_u14_u5_n153 ) , .C2( u2_u14_u5_n158 ) , .B1( u2_u14_u5_n172 ) );
  AOI222_X1 u2_u14_u5_U37 (.ZN( u2_u14_u5_n116 ) , .B2( u2_u14_u5_n145 ) , .C1( u2_u14_u5_n148 ) , .A2( u2_u14_u5_n174 ) , .C2( u2_u14_u5_n177 ) , .B1( u2_u14_u5_n187 ) , .A1( u2_u14_u5_n193 ) );
  INV_X1 u2_u14_u5_U38 (.A( u2_u14_u5_n115 ) , .ZN( u2_u14_u5_n187 ) );
  NOR2_X1 u2_u14_u5_U39 (.ZN( u2_u14_u5_n100 ) , .A1( u2_u14_u5_n170 ) , .A2( u2_u14_u5_n180 ) );
  INV_X1 u2_u14_u5_U4 (.A( u2_u14_u5_n138 ) , .ZN( u2_u14_u5_n191 ) );
  AOI22_X1 u2_u14_u5_U40 (.B2( u2_u14_u5_n131 ) , .A2( u2_u14_u5_n146 ) , .ZN( u2_u14_u5_n169 ) , .B1( u2_u14_u5_n174 ) , .A1( u2_u14_u5_n185 ) );
  NOR2_X1 u2_u14_u5_U41 (.A1( u2_u14_u5_n146 ) , .ZN( u2_u14_u5_n150 ) , .A2( u2_u14_u5_n173 ) );
  AOI21_X1 u2_u14_u5_U42 (.A( u2_u14_u5_n118 ) , .B2( u2_u14_u5_n145 ) , .ZN( u2_u14_u5_n168 ) , .B1( u2_u14_u5_n186 ) );
  INV_X1 u2_u14_u5_U43 (.A( u2_u14_u5_n122 ) , .ZN( u2_u14_u5_n186 ) );
  NOR2_X1 u2_u14_u5_U44 (.A1( u2_u14_u5_n146 ) , .ZN( u2_u14_u5_n152 ) , .A2( u2_u14_u5_n176 ) );
  NOR2_X1 u2_u14_u5_U45 (.A1( u2_u14_u5_n115 ) , .ZN( u2_u14_u5_n118 ) , .A2( u2_u14_u5_n153 ) );
  NOR2_X1 u2_u14_u5_U46 (.A2( u2_u14_u5_n145 ) , .ZN( u2_u14_u5_n156 ) , .A1( u2_u14_u5_n174 ) );
  NOR2_X1 u2_u14_u5_U47 (.ZN( u2_u14_u5_n121 ) , .A2( u2_u14_u5_n145 ) , .A1( u2_u14_u5_n176 ) );
  AOI22_X1 u2_u14_u5_U48 (.ZN( u2_u14_u5_n114 ) , .A2( u2_u14_u5_n137 ) , .A1( u2_u14_u5_n145 ) , .B2( u2_u14_u5_n175 ) , .B1( u2_u14_u5_n193 ) );
  OAI211_X1 u2_u14_u5_U49 (.B( u2_u14_u5_n124 ) , .A( u2_u14_u5_n125 ) , .C2( u2_u14_u5_n126 ) , .C1( u2_u14_u5_n127 ) , .ZN( u2_u14_u5_n128 ) );
  OAI21_X1 u2_u14_u5_U5 (.B2( u2_u14_u5_n136 ) , .B1( u2_u14_u5_n137 ) , .ZN( u2_u14_u5_n138 ) , .A( u2_u14_u5_n177 ) );
  NOR3_X1 u2_u14_u5_U50 (.ZN( u2_u14_u5_n127 ) , .A1( u2_u14_u5_n136 ) , .A3( u2_u14_u5_n148 ) , .A2( u2_u14_u5_n182 ) );
  OAI21_X1 u2_u14_u5_U51 (.ZN( u2_u14_u5_n124 ) , .A( u2_u14_u5_n177 ) , .B2( u2_u14_u5_n183 ) , .B1( u2_u14_u5_n189 ) );
  OAI21_X1 u2_u14_u5_U52 (.ZN( u2_u14_u5_n125 ) , .A( u2_u14_u5_n174 ) , .B2( u2_u14_u5_n185 ) , .B1( u2_u14_u5_n190 ) );
  AOI21_X1 u2_u14_u5_U53 (.A( u2_u14_u5_n153 ) , .B2( u2_u14_u5_n154 ) , .B1( u2_u14_u5_n155 ) , .ZN( u2_u14_u5_n164 ) );
  AOI21_X1 u2_u14_u5_U54 (.ZN( u2_u14_u5_n110 ) , .B1( u2_u14_u5_n122 ) , .B2( u2_u14_u5_n139 ) , .A( u2_u14_u5_n153 ) );
  INV_X1 u2_u14_u5_U55 (.A( u2_u14_u5_n153 ) , .ZN( u2_u14_u5_n176 ) );
  INV_X1 u2_u14_u5_U56 (.A( u2_u14_u5_n126 ) , .ZN( u2_u14_u5_n173 ) );
  AND2_X1 u2_u14_u5_U57 (.A2( u2_u14_u5_n104 ) , .A1( u2_u14_u5_n107 ) , .ZN( u2_u14_u5_n147 ) );
  AND2_X1 u2_u14_u5_U58 (.A2( u2_u14_u5_n104 ) , .A1( u2_u14_u5_n108 ) , .ZN( u2_u14_u5_n148 ) );
  NAND2_X1 u2_u14_u5_U59 (.A1( u2_u14_u5_n105 ) , .A2( u2_u14_u5_n106 ) , .ZN( u2_u14_u5_n158 ) );
  INV_X1 u2_u14_u5_U6 (.A( u2_u14_u5_n135 ) , .ZN( u2_u14_u5_n178 ) );
  NAND2_X1 u2_u14_u5_U60 (.A2( u2_u14_u5_n108 ) , .A1( u2_u14_u5_n109 ) , .ZN( u2_u14_u5_n139 ) );
  NAND2_X1 u2_u14_u5_U61 (.A1( u2_u14_u5_n106 ) , .A2( u2_u14_u5_n108 ) , .ZN( u2_u14_u5_n119 ) );
  NAND2_X1 u2_u14_u5_U62 (.A2( u2_u14_u5_n103 ) , .A1( u2_u14_u5_n105 ) , .ZN( u2_u14_u5_n140 ) );
  NAND2_X1 u2_u14_u5_U63 (.A2( u2_u14_u5_n104 ) , .A1( u2_u14_u5_n105 ) , .ZN( u2_u14_u5_n155 ) );
  NAND2_X1 u2_u14_u5_U64 (.A2( u2_u14_u5_n106 ) , .A1( u2_u14_u5_n107 ) , .ZN( u2_u14_u5_n122 ) );
  NAND2_X1 u2_u14_u5_U65 (.A2( u2_u14_u5_n100 ) , .A1( u2_u14_u5_n106 ) , .ZN( u2_u14_u5_n115 ) );
  NAND2_X1 u2_u14_u5_U66 (.A2( u2_u14_u5_n100 ) , .A1( u2_u14_u5_n103 ) , .ZN( u2_u14_u5_n161 ) );
  NAND2_X1 u2_u14_u5_U67 (.A1( u2_u14_u5_n105 ) , .A2( u2_u14_u5_n109 ) , .ZN( u2_u14_u5_n154 ) );
  INV_X1 u2_u14_u5_U68 (.A( u2_u14_u5_n146 ) , .ZN( u2_u14_u5_n172 ) );
  NAND2_X1 u2_u14_u5_U69 (.A1( u2_u14_u5_n103 ) , .A2( u2_u14_u5_n108 ) , .ZN( u2_u14_u5_n123 ) );
  OAI22_X1 u2_u14_u5_U7 (.B2( u2_u14_u5_n149 ) , .B1( u2_u14_u5_n150 ) , .A2( u2_u14_u5_n151 ) , .A1( u2_u14_u5_n152 ) , .ZN( u2_u14_u5_n165 ) );
  NAND2_X1 u2_u14_u5_U70 (.A2( u2_u14_u5_n103 ) , .A1( u2_u14_u5_n107 ) , .ZN( u2_u14_u5_n151 ) );
  NAND2_X1 u2_u14_u5_U71 (.A2( u2_u14_u5_n107 ) , .A1( u2_u14_u5_n109 ) , .ZN( u2_u14_u5_n120 ) );
  NAND2_X1 u2_u14_u5_U72 (.A2( u2_u14_u5_n100 ) , .A1( u2_u14_u5_n109 ) , .ZN( u2_u14_u5_n157 ) );
  AND2_X1 u2_u14_u5_U73 (.A2( u2_u14_u5_n100 ) , .A1( u2_u14_u5_n104 ) , .ZN( u2_u14_u5_n131 ) );
  INV_X1 u2_u14_u5_U74 (.A( u2_u14_u5_n102 ) , .ZN( u2_u14_u5_n195 ) );
  OAI221_X1 u2_u14_u5_U75 (.A( u2_u14_u5_n101 ) , .ZN( u2_u14_u5_n102 ) , .C2( u2_u14_u5_n115 ) , .C1( u2_u14_u5_n126 ) , .B1( u2_u14_u5_n134 ) , .B2( u2_u14_u5_n160 ) );
  OAI21_X1 u2_u14_u5_U76 (.ZN( u2_u14_u5_n101 ) , .B1( u2_u14_u5_n137 ) , .A( u2_u14_u5_n146 ) , .B2( u2_u14_u5_n147 ) );
  NOR2_X1 u2_u14_u5_U77 (.A2( u2_u14_X_34 ) , .A1( u2_u14_X_35 ) , .ZN( u2_u14_u5_n145 ) );
  NOR2_X1 u2_u14_u5_U78 (.A2( u2_u14_X_34 ) , .ZN( u2_u14_u5_n146 ) , .A1( u2_u14_u5_n171 ) );
  NOR2_X1 u2_u14_u5_U79 (.A2( u2_u14_X_31 ) , .A1( u2_u14_X_32 ) , .ZN( u2_u14_u5_n103 ) );
  NOR3_X1 u2_u14_u5_U8 (.A2( u2_u14_u5_n147 ) , .A1( u2_u14_u5_n148 ) , .ZN( u2_u14_u5_n149 ) , .A3( u2_u14_u5_n194 ) );
  NOR2_X1 u2_u14_u5_U80 (.A2( u2_u14_X_36 ) , .ZN( u2_u14_u5_n105 ) , .A1( u2_u14_u5_n180 ) );
  NOR2_X1 u2_u14_u5_U81 (.A2( u2_u14_X_33 ) , .ZN( u2_u14_u5_n108 ) , .A1( u2_u14_u5_n170 ) );
  NOR2_X1 u2_u14_u5_U82 (.A2( u2_u14_X_33 ) , .A1( u2_u14_X_36 ) , .ZN( u2_u14_u5_n107 ) );
  NOR2_X1 u2_u14_u5_U83 (.A2( u2_u14_X_31 ) , .ZN( u2_u14_u5_n104 ) , .A1( u2_u14_u5_n181 ) );
  NAND2_X1 u2_u14_u5_U84 (.A2( u2_u14_X_34 ) , .A1( u2_u14_X_35 ) , .ZN( u2_u14_u5_n153 ) );
  NAND2_X1 u2_u14_u5_U85 (.A1( u2_u14_X_34 ) , .ZN( u2_u14_u5_n126 ) , .A2( u2_u14_u5_n171 ) );
  AND2_X1 u2_u14_u5_U86 (.A1( u2_u14_X_31 ) , .A2( u2_u14_X_32 ) , .ZN( u2_u14_u5_n106 ) );
  AND2_X1 u2_u14_u5_U87 (.A1( u2_u14_X_31 ) , .ZN( u2_u14_u5_n109 ) , .A2( u2_u14_u5_n181 ) );
  INV_X1 u2_u14_u5_U88 (.A( u2_u14_X_33 ) , .ZN( u2_u14_u5_n180 ) );
  INV_X1 u2_u14_u5_U89 (.A( u2_u14_X_35 ) , .ZN( u2_u14_u5_n171 ) );
  NOR2_X1 u2_u14_u5_U9 (.ZN( u2_u14_u5_n135 ) , .A1( u2_u14_u5_n173 ) , .A2( u2_u14_u5_n176 ) );
  INV_X1 u2_u14_u5_U90 (.A( u2_u14_X_36 ) , .ZN( u2_u14_u5_n170 ) );
  INV_X1 u2_u14_u5_U91 (.A( u2_u14_X_32 ) , .ZN( u2_u14_u5_n181 ) );
  NAND4_X1 u2_u14_u5_U92 (.ZN( u2_out14_29 ) , .A4( u2_u14_u5_n129 ) , .A3( u2_u14_u5_n130 ) , .A2( u2_u14_u5_n168 ) , .A1( u2_u14_u5_n196 ) );
  AOI221_X1 u2_u14_u5_U93 (.A( u2_u14_u5_n128 ) , .ZN( u2_u14_u5_n129 ) , .C2( u2_u14_u5_n132 ) , .B2( u2_u14_u5_n159 ) , .B1( u2_u14_u5_n176 ) , .C1( u2_u14_u5_n184 ) );
  AOI222_X1 u2_u14_u5_U94 (.ZN( u2_u14_u5_n130 ) , .A2( u2_u14_u5_n146 ) , .B1( u2_u14_u5_n147 ) , .C2( u2_u14_u5_n175 ) , .B2( u2_u14_u5_n179 ) , .A1( u2_u14_u5_n188 ) , .C1( u2_u14_u5_n194 ) );
  NAND4_X1 u2_u14_u5_U95 (.ZN( u2_out14_19 ) , .A4( u2_u14_u5_n166 ) , .A3( u2_u14_u5_n167 ) , .A2( u2_u14_u5_n168 ) , .A1( u2_u14_u5_n169 ) );
  AOI22_X1 u2_u14_u5_U96 (.B2( u2_u14_u5_n145 ) , .A2( u2_u14_u5_n146 ) , .ZN( u2_u14_u5_n167 ) , .B1( u2_u14_u5_n182 ) , .A1( u2_u14_u5_n189 ) );
  NOR4_X1 u2_u14_u5_U97 (.A4( u2_u14_u5_n162 ) , .A3( u2_u14_u5_n163 ) , .A2( u2_u14_u5_n164 ) , .A1( u2_u14_u5_n165 ) , .ZN( u2_u14_u5_n166 ) );
  NAND4_X1 u2_u14_u5_U98 (.ZN( u2_out14_11 ) , .A4( u2_u14_u5_n143 ) , .A3( u2_u14_u5_n144 ) , .A2( u2_u14_u5_n169 ) , .A1( u2_u14_u5_n196 ) );
  AOI22_X1 u2_u14_u5_U99 (.A2( u2_u14_u5_n132 ) , .ZN( u2_u14_u5_n144 ) , .B2( u2_u14_u5_n145 ) , .B1( u2_u14_u5_n184 ) , .A1( u2_u14_u5_n194 ) );
  XOR2_X1 u2_u9_U20 (.B( u2_K10_36 ) , .A( u2_R8_25 ) , .Z( u2_u9_X_36 ) );
  XOR2_X1 u2_u9_U21 (.B( u2_K10_35 ) , .A( u2_R8_24 ) , .Z( u2_u9_X_35 ) );
  XOR2_X1 u2_u9_U23 (.B( u2_K10_33 ) , .A( u2_R8_22 ) , .Z( u2_u9_X_33 ) );
  XOR2_X1 u2_u9_U25 (.B( u2_K10_31 ) , .A( u2_R8_20 ) , .Z( u2_u9_X_31 ) );
  NOR2_X1 u2_u9_u5_U10 (.ZN( u2_u9_u5_n135 ) , .A1( u2_u9_u5_n173 ) , .A2( u2_u9_u5_n176 ) );
  NOR3_X1 u2_u9_u5_U100 (.A3( u2_u9_u5_n141 ) , .A1( u2_u9_u5_n142 ) , .ZN( u2_u9_u5_n143 ) , .A2( u2_u9_u5_n191 ) );
  NAND4_X1 u2_u9_u5_U101 (.ZN( u2_out9_4 ) , .A4( u2_u9_u5_n112 ) , .A2( u2_u9_u5_n113 ) , .A1( u2_u9_u5_n114 ) , .A3( u2_u9_u5_n195 ) );
  AOI211_X1 u2_u9_u5_U102 (.A( u2_u9_u5_n110 ) , .C1( u2_u9_u5_n111 ) , .ZN( u2_u9_u5_n112 ) , .B( u2_u9_u5_n118 ) , .C2( u2_u9_u5_n177 ) );
  INV_X1 u2_u9_u5_U103 (.A( u2_u9_u5_n102 ) , .ZN( u2_u9_u5_n195 ) );
  NAND3_X1 u2_u9_u5_U104 (.A2( u2_u9_u5_n154 ) , .A3( u2_u9_u5_n158 ) , .A1( u2_u9_u5_n161 ) , .ZN( u2_u9_u5_n99 ) );
  INV_X1 u2_u9_u5_U11 (.A( u2_u9_u5_n121 ) , .ZN( u2_u9_u5_n177 ) );
  NOR2_X1 u2_u9_u5_U12 (.ZN( u2_u9_u5_n160 ) , .A2( u2_u9_u5_n173 ) , .A1( u2_u9_u5_n177 ) );
  INV_X1 u2_u9_u5_U13 (.A( u2_u9_u5_n150 ) , .ZN( u2_u9_u5_n174 ) );
  AOI21_X1 u2_u9_u5_U14 (.A( u2_u9_u5_n160 ) , .B2( u2_u9_u5_n161 ) , .ZN( u2_u9_u5_n162 ) , .B1( u2_u9_u5_n192 ) );
  INV_X1 u2_u9_u5_U15 (.A( u2_u9_u5_n159 ) , .ZN( u2_u9_u5_n192 ) );
  AOI21_X1 u2_u9_u5_U16 (.A( u2_u9_u5_n156 ) , .B2( u2_u9_u5_n157 ) , .B1( u2_u9_u5_n158 ) , .ZN( u2_u9_u5_n163 ) );
  AOI21_X1 u2_u9_u5_U17 (.B2( u2_u9_u5_n139 ) , .B1( u2_u9_u5_n140 ) , .ZN( u2_u9_u5_n141 ) , .A( u2_u9_u5_n150 ) );
  OAI21_X1 u2_u9_u5_U18 (.A( u2_u9_u5_n133 ) , .B2( u2_u9_u5_n134 ) , .B1( u2_u9_u5_n135 ) , .ZN( u2_u9_u5_n142 ) );
  OAI21_X1 u2_u9_u5_U19 (.ZN( u2_u9_u5_n133 ) , .B2( u2_u9_u5_n147 ) , .A( u2_u9_u5_n173 ) , .B1( u2_u9_u5_n188 ) );
  NAND2_X1 u2_u9_u5_U20 (.A2( u2_u9_u5_n119 ) , .A1( u2_u9_u5_n123 ) , .ZN( u2_u9_u5_n137 ) );
  INV_X1 u2_u9_u5_U21 (.A( u2_u9_u5_n155 ) , .ZN( u2_u9_u5_n194 ) );
  NAND2_X1 u2_u9_u5_U22 (.A1( u2_u9_u5_n121 ) , .ZN( u2_u9_u5_n132 ) , .A2( u2_u9_u5_n172 ) );
  NAND2_X1 u2_u9_u5_U23 (.A2( u2_u9_u5_n122 ) , .ZN( u2_u9_u5_n136 ) , .A1( u2_u9_u5_n154 ) );
  NAND2_X1 u2_u9_u5_U24 (.A2( u2_u9_u5_n119 ) , .A1( u2_u9_u5_n120 ) , .ZN( u2_u9_u5_n159 ) );
  INV_X1 u2_u9_u5_U25 (.A( u2_u9_u5_n156 ) , .ZN( u2_u9_u5_n175 ) );
  INV_X1 u2_u9_u5_U26 (.A( u2_u9_u5_n158 ) , .ZN( u2_u9_u5_n188 ) );
  INV_X1 u2_u9_u5_U27 (.A( u2_u9_u5_n152 ) , .ZN( u2_u9_u5_n179 ) );
  INV_X1 u2_u9_u5_U28 (.A( u2_u9_u5_n140 ) , .ZN( u2_u9_u5_n182 ) );
  INV_X1 u2_u9_u5_U29 (.A( u2_u9_u5_n151 ) , .ZN( u2_u9_u5_n183 ) );
  NOR2_X1 u2_u9_u5_U3 (.ZN( u2_u9_u5_n134 ) , .A1( u2_u9_u5_n183 ) , .A2( u2_u9_u5_n190 ) );
  INV_X1 u2_u9_u5_U30 (.A( u2_u9_u5_n123 ) , .ZN( u2_u9_u5_n185 ) );
  INV_X1 u2_u9_u5_U31 (.A( u2_u9_u5_n161 ) , .ZN( u2_u9_u5_n184 ) );
  INV_X1 u2_u9_u5_U32 (.A( u2_u9_u5_n139 ) , .ZN( u2_u9_u5_n189 ) );
  INV_X1 u2_u9_u5_U33 (.A( u2_u9_u5_n157 ) , .ZN( u2_u9_u5_n190 ) );
  INV_X1 u2_u9_u5_U34 (.A( u2_u9_u5_n120 ) , .ZN( u2_u9_u5_n193 ) );
  NAND2_X1 u2_u9_u5_U35 (.ZN( u2_u9_u5_n111 ) , .A1( u2_u9_u5_n140 ) , .A2( u2_u9_u5_n155 ) );
  NOR2_X1 u2_u9_u5_U36 (.ZN( u2_u9_u5_n100 ) , .A1( u2_u9_u5_n170 ) , .A2( u2_u9_u5_n180 ) );
  INV_X1 u2_u9_u5_U37 (.A( u2_u9_u5_n117 ) , .ZN( u2_u9_u5_n196 ) );
  OAI221_X1 u2_u9_u5_U38 (.A( u2_u9_u5_n116 ) , .ZN( u2_u9_u5_n117 ) , .B2( u2_u9_u5_n119 ) , .C1( u2_u9_u5_n153 ) , .C2( u2_u9_u5_n158 ) , .B1( u2_u9_u5_n172 ) );
  AOI222_X1 u2_u9_u5_U39 (.ZN( u2_u9_u5_n116 ) , .B2( u2_u9_u5_n145 ) , .C1( u2_u9_u5_n148 ) , .A2( u2_u9_u5_n174 ) , .C2( u2_u9_u5_n177 ) , .B1( u2_u9_u5_n187 ) , .A1( u2_u9_u5_n193 ) );
  INV_X1 u2_u9_u5_U4 (.A( u2_u9_u5_n138 ) , .ZN( u2_u9_u5_n191 ) );
  INV_X1 u2_u9_u5_U40 (.A( u2_u9_u5_n115 ) , .ZN( u2_u9_u5_n187 ) );
  OAI221_X1 u2_u9_u5_U41 (.A( u2_u9_u5_n101 ) , .ZN( u2_u9_u5_n102 ) , .C2( u2_u9_u5_n115 ) , .C1( u2_u9_u5_n126 ) , .B1( u2_u9_u5_n134 ) , .B2( u2_u9_u5_n160 ) );
  OAI21_X1 u2_u9_u5_U42 (.ZN( u2_u9_u5_n101 ) , .B1( u2_u9_u5_n137 ) , .A( u2_u9_u5_n146 ) , .B2( u2_u9_u5_n147 ) );
  AOI22_X1 u2_u9_u5_U43 (.B2( u2_u9_u5_n131 ) , .A2( u2_u9_u5_n146 ) , .ZN( u2_u9_u5_n169 ) , .B1( u2_u9_u5_n174 ) , .A1( u2_u9_u5_n185 ) );
  NOR2_X1 u2_u9_u5_U44 (.A1( u2_u9_u5_n146 ) , .ZN( u2_u9_u5_n150 ) , .A2( u2_u9_u5_n173 ) );
  AOI21_X1 u2_u9_u5_U45 (.A( u2_u9_u5_n118 ) , .B2( u2_u9_u5_n145 ) , .ZN( u2_u9_u5_n168 ) , .B1( u2_u9_u5_n186 ) );
  INV_X1 u2_u9_u5_U46 (.A( u2_u9_u5_n122 ) , .ZN( u2_u9_u5_n186 ) );
  NOR2_X1 u2_u9_u5_U47 (.A1( u2_u9_u5_n146 ) , .ZN( u2_u9_u5_n152 ) , .A2( u2_u9_u5_n176 ) );
  NOR2_X1 u2_u9_u5_U48 (.A1( u2_u9_u5_n115 ) , .ZN( u2_u9_u5_n118 ) , .A2( u2_u9_u5_n153 ) );
  NOR2_X1 u2_u9_u5_U49 (.A2( u2_u9_u5_n145 ) , .ZN( u2_u9_u5_n156 ) , .A1( u2_u9_u5_n174 ) );
  OAI21_X1 u2_u9_u5_U5 (.B2( u2_u9_u5_n136 ) , .B1( u2_u9_u5_n137 ) , .ZN( u2_u9_u5_n138 ) , .A( u2_u9_u5_n177 ) );
  NOR2_X1 u2_u9_u5_U50 (.ZN( u2_u9_u5_n121 ) , .A2( u2_u9_u5_n145 ) , .A1( u2_u9_u5_n176 ) );
  AOI22_X1 u2_u9_u5_U51 (.ZN( u2_u9_u5_n114 ) , .A2( u2_u9_u5_n137 ) , .A1( u2_u9_u5_n145 ) , .B2( u2_u9_u5_n175 ) , .B1( u2_u9_u5_n193 ) );
  OAI211_X1 u2_u9_u5_U52 (.B( u2_u9_u5_n124 ) , .A( u2_u9_u5_n125 ) , .C2( u2_u9_u5_n126 ) , .C1( u2_u9_u5_n127 ) , .ZN( u2_u9_u5_n128 ) );
  NOR3_X1 u2_u9_u5_U53 (.ZN( u2_u9_u5_n127 ) , .A1( u2_u9_u5_n136 ) , .A3( u2_u9_u5_n148 ) , .A2( u2_u9_u5_n182 ) );
  OAI21_X1 u2_u9_u5_U54 (.ZN( u2_u9_u5_n124 ) , .A( u2_u9_u5_n177 ) , .B2( u2_u9_u5_n183 ) , .B1( u2_u9_u5_n189 ) );
  OAI21_X1 u2_u9_u5_U55 (.ZN( u2_u9_u5_n125 ) , .A( u2_u9_u5_n174 ) , .B2( u2_u9_u5_n185 ) , .B1( u2_u9_u5_n190 ) );
  AOI21_X1 u2_u9_u5_U56 (.A( u2_u9_u5_n153 ) , .B2( u2_u9_u5_n154 ) , .B1( u2_u9_u5_n155 ) , .ZN( u2_u9_u5_n164 ) );
  AOI21_X1 u2_u9_u5_U57 (.ZN( u2_u9_u5_n110 ) , .B1( u2_u9_u5_n122 ) , .B2( u2_u9_u5_n139 ) , .A( u2_u9_u5_n153 ) );
  INV_X1 u2_u9_u5_U58 (.A( u2_u9_u5_n153 ) , .ZN( u2_u9_u5_n176 ) );
  INV_X1 u2_u9_u5_U59 (.A( u2_u9_u5_n126 ) , .ZN( u2_u9_u5_n173 ) );
  AOI222_X1 u2_u9_u5_U6 (.ZN( u2_u9_u5_n113 ) , .A1( u2_u9_u5_n131 ) , .C1( u2_u9_u5_n148 ) , .B2( u2_u9_u5_n174 ) , .C2( u2_u9_u5_n178 ) , .A2( u2_u9_u5_n179 ) , .B1( u2_u9_u5_n99 ) );
  AND2_X1 u2_u9_u5_U60 (.A2( u2_u9_u5_n104 ) , .A1( u2_u9_u5_n107 ) , .ZN( u2_u9_u5_n147 ) );
  AND2_X1 u2_u9_u5_U61 (.A2( u2_u9_u5_n104 ) , .A1( u2_u9_u5_n108 ) , .ZN( u2_u9_u5_n148 ) );
  NAND2_X1 u2_u9_u5_U62 (.A1( u2_u9_u5_n105 ) , .A2( u2_u9_u5_n106 ) , .ZN( u2_u9_u5_n158 ) );
  NAND2_X1 u2_u9_u5_U63 (.A2( u2_u9_u5_n108 ) , .A1( u2_u9_u5_n109 ) , .ZN( u2_u9_u5_n139 ) );
  NAND2_X1 u2_u9_u5_U64 (.A1( u2_u9_u5_n106 ) , .A2( u2_u9_u5_n108 ) , .ZN( u2_u9_u5_n119 ) );
  NAND2_X1 u2_u9_u5_U65 (.A2( u2_u9_u5_n103 ) , .A1( u2_u9_u5_n105 ) , .ZN( u2_u9_u5_n140 ) );
  NAND2_X1 u2_u9_u5_U66 (.A2( u2_u9_u5_n104 ) , .A1( u2_u9_u5_n105 ) , .ZN( u2_u9_u5_n155 ) );
  NAND2_X1 u2_u9_u5_U67 (.A2( u2_u9_u5_n106 ) , .A1( u2_u9_u5_n107 ) , .ZN( u2_u9_u5_n122 ) );
  NAND2_X1 u2_u9_u5_U68 (.A2( u2_u9_u5_n100 ) , .A1( u2_u9_u5_n106 ) , .ZN( u2_u9_u5_n115 ) );
  NAND2_X1 u2_u9_u5_U69 (.A2( u2_u9_u5_n100 ) , .A1( u2_u9_u5_n103 ) , .ZN( u2_u9_u5_n161 ) );
  INV_X1 u2_u9_u5_U7 (.A( u2_u9_u5_n135 ) , .ZN( u2_u9_u5_n178 ) );
  NAND2_X1 u2_u9_u5_U70 (.A1( u2_u9_u5_n105 ) , .A2( u2_u9_u5_n109 ) , .ZN( u2_u9_u5_n154 ) );
  INV_X1 u2_u9_u5_U71 (.A( u2_u9_u5_n146 ) , .ZN( u2_u9_u5_n172 ) );
  NAND2_X1 u2_u9_u5_U72 (.A1( u2_u9_u5_n103 ) , .A2( u2_u9_u5_n108 ) , .ZN( u2_u9_u5_n123 ) );
  NAND2_X1 u2_u9_u5_U73 (.A2( u2_u9_u5_n103 ) , .A1( u2_u9_u5_n107 ) , .ZN( u2_u9_u5_n151 ) );
  NAND2_X1 u2_u9_u5_U74 (.A2( u2_u9_u5_n107 ) , .A1( u2_u9_u5_n109 ) , .ZN( u2_u9_u5_n120 ) );
  NAND2_X1 u2_u9_u5_U75 (.A2( u2_u9_u5_n100 ) , .A1( u2_u9_u5_n109 ) , .ZN( u2_u9_u5_n157 ) );
  AND2_X1 u2_u9_u5_U76 (.A2( u2_u9_u5_n100 ) , .A1( u2_u9_u5_n104 ) , .ZN( u2_u9_u5_n131 ) );
  NOR2_X1 u2_u9_u5_U77 (.A2( u2_u9_X_34 ) , .A1( u2_u9_X_35 ) , .ZN( u2_u9_u5_n145 ) );
  NOR2_X1 u2_u9_u5_U78 (.A2( u2_u9_X_34 ) , .ZN( u2_u9_u5_n146 ) , .A1( u2_u9_u5_n171 ) );
  NOR2_X1 u2_u9_u5_U79 (.A2( u2_u9_X_31 ) , .A1( u2_u9_X_32 ) , .ZN( u2_u9_u5_n103 ) );
  OAI22_X1 u2_u9_u5_U8 (.B2( u2_u9_u5_n149 ) , .B1( u2_u9_u5_n150 ) , .A2( u2_u9_u5_n151 ) , .A1( u2_u9_u5_n152 ) , .ZN( u2_u9_u5_n165 ) );
  NOR2_X1 u2_u9_u5_U80 (.A2( u2_u9_X_36 ) , .ZN( u2_u9_u5_n105 ) , .A1( u2_u9_u5_n180 ) );
  NOR2_X1 u2_u9_u5_U81 (.A2( u2_u9_X_33 ) , .ZN( u2_u9_u5_n108 ) , .A1( u2_u9_u5_n170 ) );
  NOR2_X1 u2_u9_u5_U82 (.A2( u2_u9_X_33 ) , .A1( u2_u9_X_36 ) , .ZN( u2_u9_u5_n107 ) );
  NOR2_X1 u2_u9_u5_U83 (.A2( u2_u9_X_31 ) , .ZN( u2_u9_u5_n104 ) , .A1( u2_u9_u5_n181 ) );
  NAND2_X1 u2_u9_u5_U84 (.A2( u2_u9_X_34 ) , .A1( u2_u9_X_35 ) , .ZN( u2_u9_u5_n153 ) );
  NAND2_X1 u2_u9_u5_U85 (.A1( u2_u9_X_34 ) , .ZN( u2_u9_u5_n126 ) , .A2( u2_u9_u5_n171 ) );
  AND2_X1 u2_u9_u5_U86 (.A1( u2_u9_X_31 ) , .A2( u2_u9_X_32 ) , .ZN( u2_u9_u5_n106 ) );
  AND2_X1 u2_u9_u5_U87 (.A1( u2_u9_X_31 ) , .ZN( u2_u9_u5_n109 ) , .A2( u2_u9_u5_n181 ) );
  INV_X1 u2_u9_u5_U88 (.A( u2_u9_X_33 ) , .ZN( u2_u9_u5_n180 ) );
  INV_X1 u2_u9_u5_U89 (.A( u2_u9_X_35 ) , .ZN( u2_u9_u5_n171 ) );
  NOR3_X1 u2_u9_u5_U9 (.A2( u2_u9_u5_n147 ) , .A1( u2_u9_u5_n148 ) , .ZN( u2_u9_u5_n149 ) , .A3( u2_u9_u5_n194 ) );
  INV_X1 u2_u9_u5_U90 (.A( u2_u9_X_36 ) , .ZN( u2_u9_u5_n170 ) );
  INV_X1 u2_u9_u5_U91 (.A( u2_u9_X_32 ) , .ZN( u2_u9_u5_n181 ) );
  NAND4_X1 u2_u9_u5_U92 (.ZN( u2_out9_29 ) , .A4( u2_u9_u5_n129 ) , .A3( u2_u9_u5_n130 ) , .A2( u2_u9_u5_n168 ) , .A1( u2_u9_u5_n196 ) );
  AOI221_X1 u2_u9_u5_U93 (.A( u2_u9_u5_n128 ) , .ZN( u2_u9_u5_n129 ) , .C2( u2_u9_u5_n132 ) , .B2( u2_u9_u5_n159 ) , .B1( u2_u9_u5_n176 ) , .C1( u2_u9_u5_n184 ) );
  AOI222_X1 u2_u9_u5_U94 (.ZN( u2_u9_u5_n130 ) , .A2( u2_u9_u5_n146 ) , .B1( u2_u9_u5_n147 ) , .C2( u2_u9_u5_n175 ) , .B2( u2_u9_u5_n179 ) , .A1( u2_u9_u5_n188 ) , .C1( u2_u9_u5_n194 ) );
  NAND4_X1 u2_u9_u5_U95 (.ZN( u2_out9_19 ) , .A4( u2_u9_u5_n166 ) , .A3( u2_u9_u5_n167 ) , .A2( u2_u9_u5_n168 ) , .A1( u2_u9_u5_n169 ) );
  AOI22_X1 u2_u9_u5_U96 (.B2( u2_u9_u5_n145 ) , .A2( u2_u9_u5_n146 ) , .ZN( u2_u9_u5_n167 ) , .B1( u2_u9_u5_n182 ) , .A1( u2_u9_u5_n189 ) );
  NOR4_X1 u2_u9_u5_U97 (.A4( u2_u9_u5_n162 ) , .A3( u2_u9_u5_n163 ) , .A2( u2_u9_u5_n164 ) , .A1( u2_u9_u5_n165 ) , .ZN( u2_u9_u5_n166 ) );
  NAND4_X1 u2_u9_u5_U98 (.ZN( u2_out9_11 ) , .A4( u2_u9_u5_n143 ) , .A3( u2_u9_u5_n144 ) , .A2( u2_u9_u5_n169 ) , .A1( u2_u9_u5_n196 ) );
  AOI22_X1 u2_u9_u5_U99 (.A2( u2_u9_u5_n132 ) , .ZN( u2_u9_u5_n144 ) , .B2( u2_u9_u5_n145 ) , .B1( u2_u9_u5_n184 ) , .A1( u2_u9_u5_n194 ) );
  INV_X1 u2_uk_U1044 (.A( u2_key_r_7 ) , .ZN( u2_uk_n1147 ) );
  INV_X1 u2_uk_U1047 (.A( u2_key_r_23 ) , .ZN( u2_uk_n1158 ) );
  INV_X1 u2_uk_U1049 (.A( u2_key_r_30 ) , .ZN( u2_uk_n1165 ) );
  INV_X1 u2_uk_U1055 (.A( u2_key_r_37 ) , .ZN( u2_uk_n1171 ) );
  INV_X1 u2_uk_U1057 (.A( u2_key_r_0 ) , .ZN( u2_uk_n1142 ) );
  INV_X1 u2_uk_U1058 (.A( u2_key_r_16 ) , .ZN( u2_uk_n1152 ) );
  INV_X1 u2_uk_U1092 (.ZN( u2_K1_41 ) , .A( u2_uk_n985 ) );
  AOI22_X1 u2_uk_U1093 (.B2( u2_key_r_35 ) , .A2( u2_key_r_42 ) , .A1( u2_uk_n162 ) , .B1( u2_uk_n60 ) , .ZN( u2_uk_n985 ) );
  INV_X1 u2_uk_U1118 (.ZN( u2_K1_32 ) , .A( u2_uk_n980 ) );
  AOI22_X1 u2_uk_U1119 (.B2( u2_key_r_22 ) , .A2( u2_key_r_29 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n163 ) , .ZN( u2_uk_n980 ) );
  OAI22_X1 u2_uk_U211 (.ZN( u2_K1_31 ) , .A2( u2_uk_n1147 ) , .B2( u2_uk_n1151 ) , .A1( u2_uk_n208 ) , .B1( u2_uk_n31 ) );
  INV_X1 u2_uk_U212 (.A( u2_key_r_14 ) , .ZN( u2_uk_n1151 ) );
  OAI21_X1 u2_uk_U225 (.ZN( u2_K10_31 ) , .B2( u2_uk_n1615 ) , .B1( u2_uk_n164 ) , .A( u2_uk_n291 ) );
  NAND2_X1 u2_uk_U226 (.A1( u2_uk_K_r8_16 ) , .A2( u2_uk_n155 ) , .ZN( u2_uk_n291 ) );
  OAI21_X1 u2_uk_U232 (.ZN( u2_K1_39 ) , .B2( u2_uk_n1157 ) , .B1( u2_uk_n63 ) , .A( u2_uk_n984 ) );
  INV_X1 u2_uk_U234 (.A( u2_key_r_22 ) , .ZN( u2_uk_n1157 ) );
  INV_X1 u2_uk_U247 (.ZN( u2_K1_48 ) , .A( u2_uk_n989 ) );
  AOI22_X1 u2_uk_U248 (.B2( u2_key_r_21 ) , .A2( u2_key_r_28 ) , .B1( u2_uk_n100 ) , .A1( u2_uk_n217 ) , .ZN( u2_uk_n989 ) );
  INV_X1 u2_uk_U298 (.ZN( u2_K1_26 ) , .A( u2_uk_n976 ) );
  AOI22_X1 u2_uk_U299 (.B2( u2_key_r_31 ) , .A2( u2_key_r_51 ) , .A1( u2_uk_n118 ) , .B1( u2_uk_n217 ) , .ZN( u2_uk_n976 ) );
  INV_X1 u2_uk_U305 (.ZN( u2_K15_26 ) , .A( u2_uk_n939 ) );
  OAI21_X1 u2_uk_U362 (.ZN( u2_K15_33 ) , .B1( u2_uk_n109 ) , .B2( u2_uk_n1840 ) , .A( u2_uk_n942 ) );
  INV_X1 u2_uk_U446 (.ZN( u2_K10_33 ) , .A( u2_uk_n294 ) );
  AOI22_X1 u2_uk_U447 (.B2( u2_uk_K_r8_22 ) , .A2( u2_uk_K_r8_42 ) , .A1( u2_uk_n117 ) , .B1( u2_uk_n217 ) , .ZN( u2_uk_n294 ) );
  INV_X1 u2_uk_U448 (.ZN( u2_K1_33 ) , .A( u2_uk_n981 ) );
  AOI22_X1 u2_uk_U449 (.B2( u2_key_r_44 ) , .A2( u2_key_r_51 ) , .B1( u2_uk_n100 ) , .A1( u2_uk_n163 ) , .ZN( u2_uk_n981 ) );
  OAI22_X1 u2_uk_U472 (.ZN( u2_K1_29 ) , .B2( u2_uk_n1152 ) , .A2( u2_uk_n1158 ) , .B1( u2_uk_n182 ) , .A1( u2_uk_n94 ) );
  OAI22_X1 u2_uk_U533 (.ZN( u2_K1_36 ) , .B2( u2_uk_n1158 ) , .A2( u2_uk_n1165 ) , .B1( u2_uk_n222 ) , .A1( u2_uk_n94 ) );
  OAI22_X1 u2_uk_U548 (.ZN( u2_K15_36 ) , .B2( u2_uk_n1826 ) , .A2( u2_uk_n1840 ) , .A1( u2_uk_n222 ) , .B1( u2_uk_n92 ) );
  OAI22_X1 u2_uk_U553 (.ZN( u2_K1_38 ) , .A1( u2_uk_n10 ) , .B2( u2_uk_n1165 ) , .A2( u2_uk_n1171 ) , .B1( u2_uk_n203 ) );
  INV_X1 u2_uk_U614 (.ZN( u2_K10_35 ) , .A( u2_uk_n297 ) );
  AOI22_X1 u2_uk_U615 (.B2( u2_uk_K_r8_2 ) , .A2( u2_uk_K_r8_37 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n238 ) , .ZN( u2_uk_n297 ) );
  INV_X1 u2_uk_U621 (.ZN( u2_K1_35 ) , .A( u2_uk_n982 ) );
  AOI22_X1 u2_uk_U622 (.B2( u2_key_r_28 ) , .A2( u2_key_r_35 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n207 ) , .ZN( u2_uk_n982 ) );
  INV_X1 u2_uk_U644 (.ZN( u2_K1_44 ) , .A( u2_uk_n987 ) );
  AOI22_X1 u2_uk_U645 (.B2( u2_key_r_36 ) , .A2( u2_key_r_43 ) , .B1( u2_uk_n102 ) , .A1( u2_uk_n182 ) , .ZN( u2_uk_n987 ) );
  INV_X1 u2_uk_U650 (.A( u2_key_r_44 ) , .ZN( u2_uk_n1178 ) );
  INV_X1 u2_uk_U703 (.ZN( u2_K1_25 ) , .A( u2_uk_n975 ) );
  AOI22_X1 u2_uk_U704 (.B2( u2_key_r_29 ) , .A2( u2_key_r_36 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n162 ) , .ZN( u2_uk_n975 ) );
  INV_X1 u2_uk_U739 (.ZN( u2_K1_42 ) , .A( u2_uk_n986 ) );
  OAI22_X1 u2_uk_U767 (.ZN( u2_K15_27 ) , .A2( u2_uk_n1817 ) , .B2( u2_uk_n1835 ) , .B1( u2_uk_n222 ) , .A1( u2_uk_n99 ) );
  INV_X1 u2_uk_U791 (.ZN( u2_K1_27 ) , .A( u2_uk_n977 ) );
  AOI22_X1 u2_uk_U792 (.B2( u2_key_r_14 ) , .A2( u2_key_r_21 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n162 ) , .ZN( u2_uk_n977 ) );
  OAI22_X1 u2_uk_U966 (.ZN( u2_K1_47 ) , .B2( u2_uk_n1142 ) , .A2( u2_uk_n1147 ) , .B1( u2_uk_n142 ) , .A1( u2_uk_n99 ) );
endmodule

