module des_des_die_1 ( u0_K12_34, u0_K12_35, u0_K12_36, u0_K4_43, u0_K4_48, u0_K6_11, u0_K6_13, u0_K6_16, u0_K6_19, 
       u0_K6_20, u0_K6_22, u0_K6_23, u0_K6_24, u0_K8_1, u0_K8_11, u0_K8_19, u0_K8_28, u0_K8_33, 
       u0_K8_36, u0_K8_45, u0_L0_1, u0_L0_10, u0_L0_20, u0_L0_26, u0_L10_11, u0_L10_17, u0_L10_19, 
       u0_L10_23, u0_L10_29, u0_L10_31, u0_L10_4, u0_L10_9, u0_L1_14, u0_L1_25, u0_L1_3, u0_L1_8, 
       u0_L2_12, u0_L2_15, u0_L2_21, u0_L2_22, u0_L2_27, u0_L2_32, u0_L2_5, u0_L2_7, u0_L4_1, 
       u0_L4_10, u0_L4_11, u0_L4_13, u0_L4_15, u0_L4_16, u0_L4_17, u0_L4_18, u0_L4_19, u0_L4_2, 
       u0_L4_20, u0_L4_21, u0_L4_23, u0_L4_24, u0_L4_26, u0_L4_27, u0_L4_28, u0_L4_29, u0_L4_30, 
       u0_L4_31, u0_L4_4, u0_L4_5, u0_L4_6, u0_L4_9, u0_L6_1, u0_L6_10, u0_L6_11, u0_L6_12, 
       u0_L6_13, u0_L6_14, u0_L6_15, u0_L6_16, u0_L6_17, u0_L6_18, u0_L6_19, u0_L6_2, u0_L6_20, 
       u0_L6_21, u0_L6_22, u0_L6_23, u0_L6_24, u0_L6_25, u0_L6_26, u0_L6_27, u0_L6_28, u0_L6_29, 
       u0_L6_3, u0_L6_30, u0_L6_31, u0_L6_32, u0_L6_4, u0_L6_5, u0_L6_6, u0_L6_7, u0_L6_8, 
       u0_L6_9, u0_R0_12, u0_R0_13, u0_R0_14, u0_R0_15, u0_R0_16, u0_R0_17, u0_R10_1, u0_R10_2, 
       u0_R10_20, u0_R10_21, u0_R10_22, u0_R10_23, u0_R10_24, u0_R10_25, u0_R10_3, u0_R10_32, u0_R10_4, 
       u0_R10_5, u0_R1_16, u0_R1_17, u0_R1_18, u0_R1_19, u0_R1_20, u0_R1_21, u0_R2_1, u0_R2_24, 
       u0_R2_25, u0_R2_26, u0_R2_27, u0_R2_28, u0_R2_29, u0_R2_30, u0_R2_31, u0_R2_32, u0_R4_1, 
       u0_R4_10, u0_R4_11, u0_R4_12, u0_R4_13, u0_R4_14, u0_R4_15, u0_R4_16, u0_R4_17, u0_R4_2, 
       u0_R4_20, u0_R4_21, u0_R4_22, u0_R4_23, u0_R4_24, u0_R4_25, u0_R4_28, u0_R4_29, u0_R4_3, 
       u0_R4_30, u0_R4_31, u0_R4_32, u0_R4_4, u0_R4_5, u0_R4_6, u0_R4_7, u0_R4_8, u0_R4_9, 
       u0_R6_1, u0_R6_10, u0_R6_11, u0_R6_12, u0_R6_13, u0_R6_14, u0_R6_15, u0_R6_16, u0_R6_17, 
       u0_R6_18, u0_R6_19, u0_R6_2, u0_R6_20, u0_R6_21, u0_R6_22, u0_R6_23, u0_R6_24, u0_R6_25, 
       u0_R6_26, u0_R6_27, u0_R6_28, u0_R6_29, u0_R6_3, u0_R6_30, u0_R6_31, u0_R6_32, u0_R6_4, 
       u0_R6_5, u0_R6_6, u0_R6_7, u0_R6_8, u0_R6_9, u0_key_r_10, u0_key_r_45, u0_key_r_46, u0_uk_K_r0_11, 
       u0_uk_K_r0_47, u0_uk_K_r10_10, u0_uk_K_r10_14, u0_uk_K_r10_16, u0_uk_K_r10_18, u0_uk_K_r10_19, u0_uk_K_r10_23, u0_uk_K_r10_27, u0_uk_K_r10_28, 
       u0_uk_K_r10_39, u0_uk_K_r10_44, u0_uk_K_r10_48, u0_uk_K_r11_28, u0_uk_K_r11_8, u0_uk_K_r1_36, u0_uk_K_r1_42, u0_uk_K_r1_44, u0_uk_K_r2_50, 
       u0_uk_K_r3_4, u0_uk_K_r4_11, u0_uk_K_r4_23, u0_uk_K_r4_3, u0_uk_K_r4_33, u0_uk_K_r4_4, u0_uk_K_r4_41, u0_uk_K_r4_47, u0_uk_K_r4_48, 
       u0_uk_K_r4_49, u0_uk_K_r4_5, u0_uk_K_r4_54, u0_uk_K_r4_55, u0_uk_K_r5_13, u0_uk_K_r6_0, u0_uk_K_r6_10, u0_uk_K_r6_14, u0_uk_K_r6_19, 
       u0_uk_K_r6_21, u0_uk_K_r6_22, u0_uk_K_r6_26, u0_uk_K_r6_27, u0_uk_K_r6_29, u0_uk_K_r6_3, u0_uk_K_r6_31, u0_uk_K_r6_34, u0_uk_K_r6_37, 
       u0_uk_K_r6_46, u0_uk_K_r6_53, u0_uk_K_r6_7, u0_uk_K_r8_21, u0_uk_K_r8_43, u0_uk_n10, u0_uk_n100, u0_uk_n109, u0_uk_n110, 
       u0_uk_n118, u0_uk_n128, u0_uk_n140, u0_uk_n142, u0_uk_n146, u0_uk_n147, u0_uk_n148, u0_uk_n150, u0_uk_n156, 
       u0_uk_n161, u0_uk_n163, u0_uk_n164, u0_uk_n172, u0_uk_n173, u0_uk_n176, u0_uk_n177, u0_uk_n188, u0_uk_n191, 
       u0_uk_n203, u0_uk_n207, u0_uk_n208, u0_uk_n209, u0_uk_n214, u0_uk_n217, u0_uk_n220, u0_uk_n222, u0_uk_n230, 
       u0_uk_n231, u0_uk_n238, u0_uk_n240, u0_uk_n250, u0_uk_n251, u0_uk_n252, u0_uk_n257, u0_uk_n31, u0_uk_n318, 
       u0_uk_n320, u0_uk_n321, u0_uk_n322, u0_uk_n323, u0_uk_n324, u0_uk_n325, u0_uk_n326, u0_uk_n327, u0_uk_n328, 
       u0_uk_n329, u0_uk_n330, u0_uk_n331, u0_uk_n332, u0_uk_n333, u0_uk_n336, u0_uk_n337, u0_uk_n339, u0_uk_n340, 
       u0_uk_n341, u0_uk_n343, u0_uk_n344, u0_uk_n345, u0_uk_n347, u0_uk_n348, u0_uk_n350, u0_uk_n351, u0_uk_n352, 
       u0_uk_n354, u0_uk_n355, u0_uk_n356, u0_uk_n357, u0_uk_n358, u0_uk_n359, u0_uk_n410, u0_uk_n411, u0_uk_n412, 
       u0_uk_n414, u0_uk_n417, u0_uk_n418, u0_uk_n419, u0_uk_n423, u0_uk_n424, u0_uk_n425, u0_uk_n426, u0_uk_n427, 
       u0_uk_n428, u0_uk_n429, u0_uk_n430, u0_uk_n432, u0_uk_n433, u0_uk_n434, u0_uk_n435, u0_uk_n436, u0_uk_n439, 
       u0_uk_n440, u0_uk_n441, u0_uk_n442, u0_uk_n445, u0_uk_n447, u0_uk_n448, u0_uk_n450, u0_uk_n498, u0_uk_n499, 
       u0_uk_n505, u0_uk_n506, u0_uk_n508, u0_uk_n513, u0_uk_n514, u0_uk_n516, u0_uk_n521, u0_uk_n522, u0_uk_n527, 
       u0_uk_n528, u0_uk_n537, u0_uk_n538, u0_uk_n539, u0_uk_n543, u0_uk_n544, u0_uk_n545, u0_uk_n555, u0_uk_n559, 
       u0_uk_n560, u0_uk_n570, u0_uk_n575, u0_uk_n579, u0_uk_n589, u0_uk_n596, u0_uk_n598, u0_uk_n609, u0_uk_n610, 
       u0_uk_n615, u0_uk_n620, u0_uk_n624, u0_uk_n625, u0_uk_n63, u0_uk_n746, u0_uk_n748, u0_uk_n755, u0_uk_n759, 
       u0_uk_n785, u0_uk_n786, u0_uk_n793, u0_uk_n799, u0_uk_n83, u0_uk_n92, u0_uk_n93, u0_uk_n963, u1_FP_42, 
       u1_FP_43, u1_FP_54, u1_FP_55, u1_K10_10, u1_K10_11, u1_K10_13, u1_K10_14, u1_K10_15, u1_K10_16, 
       u1_K10_17, u1_K10_18, u1_K10_19, u1_K10_20, u1_K10_21, u1_K10_34, u1_K10_36, u1_K12_39, u1_K12_40, 
       u1_K12_45, u1_K12_46, u1_K15_21, u1_K15_22, u1_K16_15, u1_K16_16, u1_K16_33, u1_K1_28, u1_K1_29, 
       u1_K1_31, u1_K1_34, u1_K2_9, u1_K3_10, u1_K3_9, u1_K4_39, u1_K4_40, u1_K4_9, u1_K6_45, 
       u1_K6_46, u1_K7_10, u1_K7_45, u1_K7_9, u1_K8_45, u1_K8_46, u1_K9_3, u1_K9_4, u1_L0_13, 
       u1_L0_18, u1_L0_2, u1_L0_28, u1_L10_12, u1_L10_15, u1_L10_21, u1_L10_22, u1_L10_27, u1_L10_32, 
       u1_L10_5, u1_L10_7, u1_L13_1, u1_L13_10, u1_L13_20, u1_L13_26, u1_L14_11, u1_L14_16, u1_L14_19, 
       u1_L14_24, u1_L14_29, u1_L14_30, u1_L14_4, u1_L14_6, u1_L1_13, u1_L1_18, u1_L1_2, u1_L1_28, 
       u1_L2_12, u1_L2_13, u1_L2_18, u1_L2_2, u1_L2_22, u1_L2_28, u1_L2_32, u1_L2_7, u1_L4_15, 
       u1_L4_21, u1_L4_27, u1_L4_5, u1_L5_13, u1_L5_15, u1_L5_18, u1_L5_2, u1_L5_21, u1_L5_27, 
       u1_L5_28, u1_L5_5, u1_L6_15, u1_L6_21, u1_L6_27, u1_L6_5, u1_L7_17, u1_L7_23, u1_L7_31, 
       u1_L7_9, u1_L8_1, u1_L8_10, u1_L8_11, u1_L8_12, u1_L8_13, u1_L8_16, u1_L8_18, u1_L8_19, 
       u1_L8_2, u1_L8_20, u1_L8_22, u1_L8_24, u1_L8_26, u1_L8_28, u1_L8_29, u1_L8_30, u1_L8_32, 
       u1_L8_4, u1_L8_6, u1_L8_7, u1_R0_6, u1_R0_7, u1_R10_26, u1_R10_27, u1_R10_30, u1_R10_31, 
       u1_R13_14, u1_R13_15, u1_R1_6, u1_R1_7, u1_R2_26, u1_R2_27, u1_R2_6, u1_R2_7, u1_R4_30, 
       u1_R4_31, u1_R5_30, u1_R5_31, u1_R5_6, u1_R5_7, u1_R6_30, u1_R6_31, u1_R7_2, u1_R7_3, 
       u1_R8_10, u1_R8_11, u1_R8_12, u1_R8_13, u1_R8_14, u1_R8_15, u1_R8_22, u1_R8_23, u1_R8_24, 
       u1_R8_25, u1_R8_26, u1_R8_27, u1_R8_6, u1_R8_7, u1_R8_8, u1_R8_9, u1_desIn_r_0, u1_desIn_r_11, 
       u1_desIn_r_18, u1_desIn_r_19, u1_desIn_r_20, u1_desIn_r_22, u1_desIn_r_27, u1_desIn_r_30, u1_desIn_r_32, u1_desIn_r_43, u1_desIn_r_44, 
       u1_desIn_r_51, u1_desIn_r_62, u1_u0_X_25, u1_u0_X_26, u1_u0_X_30, u1_u0_X_32, u1_u0_X_35, u1_u0_X_36, u1_u11_X_37, 
       u1_u11_X_38, u1_u11_X_41, u1_u11_X_42, u1_u11_X_43, u1_u11_X_44, u1_u11_X_47, u1_u11_X_48, u1_u14_X_19, u1_u14_X_20, 
       u1_u14_X_23, u1_u14_X_24, u1_u15_X_13, u1_u15_X_14, u1_u15_X_17, u1_u15_X_18, u1_u15_X_31, u1_u15_X_32, u1_u15_X_35, 
       u1_u15_X_36, u1_u1_X_11, u1_u1_X_12, u1_u1_X_7, u1_u1_X_8, u1_u2_X_11, u1_u2_X_12, u1_u2_X_7, u1_u2_X_8, 
       u1_u3_X_11, u1_u3_X_12, u1_u3_X_37, u1_u3_X_38, u1_u3_X_41, u1_u3_X_42, u1_u3_X_7, u1_u3_X_8, u1_u5_X_43, 
       u1_u5_X_44, u1_u5_X_47, u1_u5_X_48, u1_u6_X_11, u1_u6_X_12, u1_u6_X_43, u1_u6_X_44, u1_u6_X_47, u1_u6_X_48, 
       u1_u6_X_7, u1_u6_X_8, u1_u7_X_43, u1_u7_X_44, u1_u7_X_47, u1_u7_X_48, u1_u8_X_1, u1_u8_X_2, u1_u8_X_5, 
       u1_u8_X_6, u1_u9_X_23, u1_u9_X_24, u1_u9_X_31, u1_u9_X_32, u1_u9_X_41, u1_u9_X_42, u1_u9_X_7, u1_u9_X_8, 
       u1_uk_n1007, u1_uk_n1011, u1_uk_n1021, u1_uk_n1050, u1_uk_n1124, u1_uk_n299, u1_uk_n312, u1_uk_n349, u1_uk_n353, 
       u1_uk_n366, u1_uk_n369, u1_uk_n373, u1_uk_n375, u1_uk_n376, u1_uk_n988, u2_K2_1, u2_K2_43, u2_K2_44, 
       u2_K2_45, u2_K2_46, u2_K2_47, u2_K2_48, u2_L0_15, u2_L0_17, u2_L0_21, u2_L0_23, u2_L0_27, 
       u2_L0_31, u2_L0_5, u2_L0_9, u2_R0_1, u2_R0_2, u2_R0_28, u2_R0_29, u2_R0_3, u2_R0_30, 
       u2_R0_31, u2_R0_32, u2_R0_4, u2_R0_5, u2_uk_n10, u2_uk_n1238, u2_uk_n1239, u2_uk_n1243, u2_uk_n1244, 
       u2_uk_n1247, u2_uk_n1249, u2_uk_n1254, u2_uk_n1267, u2_uk_n1270, u2_uk_n1275, u2_uk_n129, u2_uk_n142, u2_uk_n213, 
       u2_uk_n220, u2_uk_n31, u2_uk_n83, u2_uk_n99, u0_N100, u0_N102, u0_N107, u0_N110, u0_N116, u0_N117, u0_N122, u0_N127, u0_N160, 
        u0_N161, u0_N163, u0_N164, u0_N165, u0_N168, u0_N169, u0_N170, u0_N172, u0_N174, 
        u0_N175, u0_N176, u0_N177, u0_N178, u0_N179, u0_N180, u0_N182, u0_N183, u0_N185, 
        u0_N186, u0_N187, u0_N188, u0_N189, u0_N190, u0_N224, u0_N225, u0_N226, u0_N227, 
        u0_N228, u0_N229, u0_N230, u0_N231, u0_N232, u0_N233, u0_N234, u0_N235, u0_N236, 
        u0_N237, u0_N238, u0_N239, u0_N240, u0_N241, u0_N242, u0_N243, u0_N244, u0_N245, 
        u0_N246, u0_N247, u0_N248, u0_N249, u0_N250, u0_N251, u0_N252, u0_N253, u0_N254, 
        u0_N255, u0_N32, u0_N355, u0_N360, u0_N362, u0_N368, u0_N370, u0_N374, u0_N380, 
        u0_N382, u0_N41, u0_N51, u0_N57, u0_N66, u0_N71, u0_N77, u0_N88, u0_uk_n1010, 
        u0_uk_n1016, u0_uk_n102, u0_uk_n11, u0_uk_n117, u0_uk_n141, u0_uk_n145, u0_uk_n162, u0_uk_n182, u0_uk_n202, 
        u0_uk_n213, u0_uk_n223, u0_uk_n242, u0_uk_n27, u0_uk_n60, u0_uk_n777, u0_uk_n798, u0_uk_n804, u0_uk_n848, 
        u0_uk_n880, u0_uk_n888, u0_uk_n890, u0_uk_n942, u0_uk_n945, u0_uk_n961, u0_uk_n969, u1_FP_11, u1_FP_16, 
        u1_FP_19, u1_FP_24, u1_FP_29, u1_FP_30, u1_FP_4, u1_FP_6, u1_N10, u1_N102, u1_N107, 
        u1_N108, u1_N113, u1_N117, u1_N123, u1_N127, u1_N13, u1_N164, u1_N174, u1_N18, 
        u1_N180, u1_N186, u1_N193, u1_N196, u1_N2, u1_N204, u1_N206, u1_N209, u1_N212, 
        u1_N218, u1_N219, u1_N228, u1_N238, u1_N24, u1_N244, u1_N250, u1_N264, u1_N272, 
        u1_N278, u1_N28, u1_N286, u1_N288, u1_N289, u1_N291, u1_N293, u1_N294, u1_N297, 
        u1_N298, u1_N299, u1_N3, u1_N300, u1_N303, u1_N305, u1_N306, u1_N307, u1_N309, 
        u1_N311, u1_N313, u1_N315, u1_N316, u1_N317, u1_N319, u1_N33, u1_N356, u1_N358, 
        u1_N363, u1_N366, u1_N372, u1_N373, u1_N378, u1_N383, u1_N44, u1_N448, u1_N457, 
        u1_N467, u1_N473, u1_N49, u1_N59, u1_N65, u1_N7, u1_N76, u1_N81, u1_N91, 
        u1_N97, u2_N36, u2_N40, u2_N46, u2_N48, u2_N52, u2_N54, u2_N58, u2_N62 );
  input u0_K12_34, u0_K12_35, u0_K12_36, u0_K4_43, u0_K4_48, u0_K6_11, u0_K6_13, u0_K6_16, u0_K6_19, 
        u0_K6_20, u0_K6_22, u0_K6_23, u0_K6_24, u0_K8_1, u0_K8_11, u0_K8_19, u0_K8_28, u0_K8_33, 
        u0_K8_36, u0_K8_45, u0_L0_1, u0_L0_10, u0_L0_20, u0_L0_26, u0_L10_11, u0_L10_17, u0_L10_19, 
        u0_L10_23, u0_L10_29, u0_L10_31, u0_L10_4, u0_L10_9, u0_L1_14, u0_L1_25, u0_L1_3, u0_L1_8, 
        u0_L2_12, u0_L2_15, u0_L2_21, u0_L2_22, u0_L2_27, u0_L2_32, u0_L2_5, u0_L2_7, u0_L4_1, 
        u0_L4_10, u0_L4_11, u0_L4_13, u0_L4_15, u0_L4_16, u0_L4_17, u0_L4_18, u0_L4_19, u0_L4_2, 
        u0_L4_20, u0_L4_21, u0_L4_23, u0_L4_24, u0_L4_26, u0_L4_27, u0_L4_28, u0_L4_29, u0_L4_30, 
        u0_L4_31, u0_L4_4, u0_L4_5, u0_L4_6, u0_L4_9, u0_L6_1, u0_L6_10, u0_L6_11, u0_L6_12, 
        u0_L6_13, u0_L6_14, u0_L6_15, u0_L6_16, u0_L6_17, u0_L6_18, u0_L6_19, u0_L6_2, u0_L6_20, 
        u0_L6_21, u0_L6_22, u0_L6_23, u0_L6_24, u0_L6_25, u0_L6_26, u0_L6_27, u0_L6_28, u0_L6_29, 
        u0_L6_3, u0_L6_30, u0_L6_31, u0_L6_32, u0_L6_4, u0_L6_5, u0_L6_6, u0_L6_7, u0_L6_8, 
        u0_L6_9, u0_R0_12, u0_R0_13, u0_R0_14, u0_R0_15, u0_R0_16, u0_R0_17, u0_R10_1, u0_R10_2, 
        u0_R10_20, u0_R10_21, u0_R10_22, u0_R10_23, u0_R10_24, u0_R10_25, u0_R10_3, u0_R10_32, u0_R10_4, 
        u0_R10_5, u0_R1_16, u0_R1_17, u0_R1_18, u0_R1_19, u0_R1_20, u0_R1_21, u0_R2_1, u0_R2_24, 
        u0_R2_25, u0_R2_26, u0_R2_27, u0_R2_28, u0_R2_29, u0_R2_30, u0_R2_31, u0_R2_32, u0_R4_1, 
        u0_R4_10, u0_R4_11, u0_R4_12, u0_R4_13, u0_R4_14, u0_R4_15, u0_R4_16, u0_R4_17, u0_R4_2, 
        u0_R4_20, u0_R4_21, u0_R4_22, u0_R4_23, u0_R4_24, u0_R4_25, u0_R4_28, u0_R4_29, u0_R4_3, 
        u0_R4_30, u0_R4_31, u0_R4_32, u0_R4_4, u0_R4_5, u0_R4_6, u0_R4_7, u0_R4_8, u0_R4_9, 
        u0_R6_1, u0_R6_10, u0_R6_11, u0_R6_12, u0_R6_13, u0_R6_14, u0_R6_15, u0_R6_16, u0_R6_17, 
        u0_R6_18, u0_R6_19, u0_R6_2, u0_R6_20, u0_R6_21, u0_R6_22, u0_R6_23, u0_R6_24, u0_R6_25, 
        u0_R6_26, u0_R6_27, u0_R6_28, u0_R6_29, u0_R6_3, u0_R6_30, u0_R6_31, u0_R6_32, u0_R6_4, 
        u0_R6_5, u0_R6_6, u0_R6_7, u0_R6_8, u0_R6_9, u0_key_r_10, u0_key_r_45, u0_key_r_46, u0_uk_K_r0_11, 
        u0_uk_K_r0_47, u0_uk_K_r10_10, u0_uk_K_r10_14, u0_uk_K_r10_16, u0_uk_K_r10_18, u0_uk_K_r10_19, u0_uk_K_r10_23, u0_uk_K_r10_27, u0_uk_K_r10_28, 
        u0_uk_K_r10_39, u0_uk_K_r10_44, u0_uk_K_r10_48, u0_uk_K_r11_28, u0_uk_K_r11_8, u0_uk_K_r1_36, u0_uk_K_r1_42, u0_uk_K_r1_44, u0_uk_K_r2_50, 
        u0_uk_K_r3_4, u0_uk_K_r4_11, u0_uk_K_r4_23, u0_uk_K_r4_3, u0_uk_K_r4_33, u0_uk_K_r4_4, u0_uk_K_r4_41, u0_uk_K_r4_47, u0_uk_K_r4_48, 
        u0_uk_K_r4_49, u0_uk_K_r4_5, u0_uk_K_r4_54, u0_uk_K_r4_55, u0_uk_K_r5_13, u0_uk_K_r6_0, u0_uk_K_r6_10, u0_uk_K_r6_14, u0_uk_K_r6_19, 
        u0_uk_K_r6_21, u0_uk_K_r6_22, u0_uk_K_r6_26, u0_uk_K_r6_27, u0_uk_K_r6_29, u0_uk_K_r6_3, u0_uk_K_r6_31, u0_uk_K_r6_34, u0_uk_K_r6_37, 
        u0_uk_K_r6_46, u0_uk_K_r6_53, u0_uk_K_r6_7, u0_uk_K_r8_21, u0_uk_K_r8_43, u0_uk_n10, u0_uk_n100, u0_uk_n109, u0_uk_n110, 
        u0_uk_n118, u0_uk_n128, u0_uk_n140, u0_uk_n142, u0_uk_n146, u0_uk_n147, u0_uk_n148, u0_uk_n150, u0_uk_n156, 
        u0_uk_n161, u0_uk_n163, u0_uk_n164, u0_uk_n172, u0_uk_n173, u0_uk_n176, u0_uk_n177, u0_uk_n188, u0_uk_n191, 
        u0_uk_n203, u0_uk_n207, u0_uk_n208, u0_uk_n209, u0_uk_n214, u0_uk_n217, u0_uk_n220, u0_uk_n222, u0_uk_n230, 
        u0_uk_n231, u0_uk_n238, u0_uk_n240, u0_uk_n250, u0_uk_n251, u0_uk_n252, u0_uk_n257, u0_uk_n31, u0_uk_n318, 
        u0_uk_n320, u0_uk_n321, u0_uk_n322, u0_uk_n323, u0_uk_n324, u0_uk_n325, u0_uk_n326, u0_uk_n327, u0_uk_n328, 
        u0_uk_n329, u0_uk_n330, u0_uk_n331, u0_uk_n332, u0_uk_n333, u0_uk_n336, u0_uk_n337, u0_uk_n339, u0_uk_n340, 
        u0_uk_n341, u0_uk_n343, u0_uk_n344, u0_uk_n345, u0_uk_n347, u0_uk_n348, u0_uk_n350, u0_uk_n351, u0_uk_n352, 
        u0_uk_n354, u0_uk_n355, u0_uk_n356, u0_uk_n357, u0_uk_n358, u0_uk_n359, u0_uk_n410, u0_uk_n411, u0_uk_n412, 
        u0_uk_n414, u0_uk_n417, u0_uk_n418, u0_uk_n419, u0_uk_n423, u0_uk_n424, u0_uk_n425, u0_uk_n426, u0_uk_n427, 
        u0_uk_n428, u0_uk_n429, u0_uk_n430, u0_uk_n432, u0_uk_n433, u0_uk_n434, u0_uk_n435, u0_uk_n436, u0_uk_n439, 
        u0_uk_n440, u0_uk_n441, u0_uk_n442, u0_uk_n445, u0_uk_n447, u0_uk_n448, u0_uk_n450, u0_uk_n498, u0_uk_n499, 
        u0_uk_n505, u0_uk_n506, u0_uk_n508, u0_uk_n513, u0_uk_n514, u0_uk_n516, u0_uk_n521, u0_uk_n522, u0_uk_n527, 
        u0_uk_n528, u0_uk_n537, u0_uk_n538, u0_uk_n539, u0_uk_n543, u0_uk_n544, u0_uk_n545, u0_uk_n555, u0_uk_n559, 
        u0_uk_n560, u0_uk_n570, u0_uk_n575, u0_uk_n579, u0_uk_n589, u0_uk_n596, u0_uk_n598, u0_uk_n609, u0_uk_n610, 
        u0_uk_n615, u0_uk_n620, u0_uk_n624, u0_uk_n625, u0_uk_n63, u0_uk_n746, u0_uk_n748, u0_uk_n755, u0_uk_n759, 
        u0_uk_n785, u0_uk_n786, u0_uk_n793, u0_uk_n799, u0_uk_n83, u0_uk_n92, u0_uk_n93, u0_uk_n963, u1_FP_42, 
        u1_FP_43, u1_FP_54, u1_FP_55, u1_K10_10, u1_K10_11, u1_K10_13, u1_K10_14, u1_K10_15, u1_K10_16, 
        u1_K10_17, u1_K10_18, u1_K10_19, u1_K10_20, u1_K10_21, u1_K10_34, u1_K10_36, u1_K12_39, u1_K12_40, 
        u1_K12_45, u1_K12_46, u1_K15_21, u1_K15_22, u1_K16_15, u1_K16_16, u1_K16_33, u1_K1_28, u1_K1_29, 
        u1_K1_31, u1_K1_34, u1_K2_9, u1_K3_10, u1_K3_9, u1_K4_39, u1_K4_40, u1_K4_9, u1_K6_45, 
        u1_K6_46, u1_K7_10, u1_K7_45, u1_K7_9, u1_K8_45, u1_K8_46, u1_K9_3, u1_K9_4, u1_L0_13, 
        u1_L0_18, u1_L0_2, u1_L0_28, u1_L10_12, u1_L10_15, u1_L10_21, u1_L10_22, u1_L10_27, u1_L10_32, 
        u1_L10_5, u1_L10_7, u1_L13_1, u1_L13_10, u1_L13_20, u1_L13_26, u1_L14_11, u1_L14_16, u1_L14_19, 
        u1_L14_24, u1_L14_29, u1_L14_30, u1_L14_4, u1_L14_6, u1_L1_13, u1_L1_18, u1_L1_2, u1_L1_28, 
        u1_L2_12, u1_L2_13, u1_L2_18, u1_L2_2, u1_L2_22, u1_L2_28, u1_L2_32, u1_L2_7, u1_L4_15, 
        u1_L4_21, u1_L4_27, u1_L4_5, u1_L5_13, u1_L5_15, u1_L5_18, u1_L5_2, u1_L5_21, u1_L5_27, 
        u1_L5_28, u1_L5_5, u1_L6_15, u1_L6_21, u1_L6_27, u1_L6_5, u1_L7_17, u1_L7_23, u1_L7_31, 
        u1_L7_9, u1_L8_1, u1_L8_10, u1_L8_11, u1_L8_12, u1_L8_13, u1_L8_16, u1_L8_18, u1_L8_19, 
        u1_L8_2, u1_L8_20, u1_L8_22, u1_L8_24, u1_L8_26, u1_L8_28, u1_L8_29, u1_L8_30, u1_L8_32, 
        u1_L8_4, u1_L8_6, u1_L8_7, u1_R0_6, u1_R0_7, u1_R10_26, u1_R10_27, u1_R10_30, u1_R10_31, 
        u1_R13_14, u1_R13_15, u1_R1_6, u1_R1_7, u1_R2_26, u1_R2_27, u1_R2_6, u1_R2_7, u1_R4_30, 
        u1_R4_31, u1_R5_30, u1_R5_31, u1_R5_6, u1_R5_7, u1_R6_30, u1_R6_31, u1_R7_2, u1_R7_3, 
        u1_R8_10, u1_R8_11, u1_R8_12, u1_R8_13, u1_R8_14, u1_R8_15, u1_R8_22, u1_R8_23, u1_R8_24, 
        u1_R8_25, u1_R8_26, u1_R8_27, u1_R8_6, u1_R8_7, u1_R8_8, u1_R8_9, u1_desIn_r_0, u1_desIn_r_11, 
        u1_desIn_r_18, u1_desIn_r_19, u1_desIn_r_20, u1_desIn_r_22, u1_desIn_r_27, u1_desIn_r_30, u1_desIn_r_32, u1_desIn_r_43, u1_desIn_r_44, 
        u1_desIn_r_51, u1_desIn_r_62, u1_u0_X_25, u1_u0_X_26, u1_u0_X_30, u1_u0_X_32, u1_u0_X_35, u1_u0_X_36, u1_u11_X_37, 
        u1_u11_X_38, u1_u11_X_41, u1_u11_X_42, u1_u11_X_43, u1_u11_X_44, u1_u11_X_47, u1_u11_X_48, u1_u14_X_19, u1_u14_X_20, 
        u1_u14_X_23, u1_u14_X_24, u1_u15_X_13, u1_u15_X_14, u1_u15_X_17, u1_u15_X_18, u1_u15_X_31, u1_u15_X_32, u1_u15_X_35, 
        u1_u15_X_36, u1_u1_X_11, u1_u1_X_12, u1_u1_X_7, u1_u1_X_8, u1_u2_X_11, u1_u2_X_12, u1_u2_X_7, u1_u2_X_8, 
        u1_u3_X_11, u1_u3_X_12, u1_u3_X_37, u1_u3_X_38, u1_u3_X_41, u1_u3_X_42, u1_u3_X_7, u1_u3_X_8, u1_u5_X_43, 
        u1_u5_X_44, u1_u5_X_47, u1_u5_X_48, u1_u6_X_11, u1_u6_X_12, u1_u6_X_43, u1_u6_X_44, u1_u6_X_47, u1_u6_X_48, 
        u1_u6_X_7, u1_u6_X_8, u1_u7_X_43, u1_u7_X_44, u1_u7_X_47, u1_u7_X_48, u1_u8_X_1, u1_u8_X_2, u1_u8_X_5, 
        u1_u8_X_6, u1_u9_X_23, u1_u9_X_24, u1_u9_X_31, u1_u9_X_32, u1_u9_X_41, u1_u9_X_42, u1_u9_X_7, u1_u9_X_8, 
        u1_uk_n1007, u1_uk_n1011, u1_uk_n1021, u1_uk_n1050, u1_uk_n1124, u1_uk_n299, u1_uk_n312, u1_uk_n349, u1_uk_n353, 
        u1_uk_n366, u1_uk_n369, u1_uk_n373, u1_uk_n375, u1_uk_n376, u1_uk_n988, u2_K2_1, u2_K2_43, u2_K2_44, 
        u2_K2_45, u2_K2_46, u2_K2_47, u2_K2_48, u2_L0_15, u2_L0_17, u2_L0_21, u2_L0_23, u2_L0_27, 
        u2_L0_31, u2_L0_5, u2_L0_9, u2_R0_1, u2_R0_2, u2_R0_28, u2_R0_29, u2_R0_3, u2_R0_30, 
        u2_R0_31, u2_R0_32, u2_R0_4, u2_R0_5, u2_uk_n10, u2_uk_n1238, u2_uk_n1239, u2_uk_n1243, u2_uk_n1244, 
        u2_uk_n1247, u2_uk_n1249, u2_uk_n1254, u2_uk_n1267, u2_uk_n1270, u2_uk_n1275, u2_uk_n129, u2_uk_n142, u2_uk_n213, 
        u2_uk_n220, u2_uk_n31, u2_uk_n83, u2_uk_n99;
  output u0_N100, u0_N102, u0_N107, u0_N110, u0_N116, u0_N117, u0_N122, u0_N127, u0_N160, 
        u0_N161, u0_N163, u0_N164, u0_N165, u0_N168, u0_N169, u0_N170, u0_N172, u0_N174, 
        u0_N175, u0_N176, u0_N177, u0_N178, u0_N179, u0_N180, u0_N182, u0_N183, u0_N185, 
        u0_N186, u0_N187, u0_N188, u0_N189, u0_N190, u0_N224, u0_N225, u0_N226, u0_N227, 
        u0_N228, u0_N229, u0_N230, u0_N231, u0_N232, u0_N233, u0_N234, u0_N235, u0_N236, 
        u0_N237, u0_N238, u0_N239, u0_N240, u0_N241, u0_N242, u0_N243, u0_N244, u0_N245, 
        u0_N246, u0_N247, u0_N248, u0_N249, u0_N250, u0_N251, u0_N252, u0_N253, u0_N254, 
        u0_N255, u0_N32, u0_N355, u0_N360, u0_N362, u0_N368, u0_N370, u0_N374, u0_N380, 
        u0_N382, u0_N41, u0_N51, u0_N57, u0_N66, u0_N71, u0_N77, u0_N88, u0_uk_n1010, 
        u0_uk_n1016, u0_uk_n102, u0_uk_n11, u0_uk_n117, u0_uk_n141, u0_uk_n145, u0_uk_n162, u0_uk_n182, u0_uk_n202, 
        u0_uk_n213, u0_uk_n223, u0_uk_n242, u0_uk_n27, u0_uk_n60, u0_uk_n777, u0_uk_n798, u0_uk_n804, u0_uk_n848, 
        u0_uk_n880, u0_uk_n888, u0_uk_n890, u0_uk_n942, u0_uk_n945, u0_uk_n961, u0_uk_n969, u1_FP_11, u1_FP_16, 
        u1_FP_19, u1_FP_24, u1_FP_29, u1_FP_30, u1_FP_4, u1_FP_6, u1_N10, u1_N102, u1_N107, 
        u1_N108, u1_N113, u1_N117, u1_N123, u1_N127, u1_N13, u1_N164, u1_N174, u1_N18, 
        u1_N180, u1_N186, u1_N193, u1_N196, u1_N2, u1_N204, u1_N206, u1_N209, u1_N212, 
        u1_N218, u1_N219, u1_N228, u1_N238, u1_N24, u1_N244, u1_N250, u1_N264, u1_N272, 
        u1_N278, u1_N28, u1_N286, u1_N288, u1_N289, u1_N291, u1_N293, u1_N294, u1_N297, 
        u1_N298, u1_N299, u1_N3, u1_N300, u1_N303, u1_N305, u1_N306, u1_N307, u1_N309, 
        u1_N311, u1_N313, u1_N315, u1_N316, u1_N317, u1_N319, u1_N33, u1_N356, u1_N358, 
        u1_N363, u1_N366, u1_N372, u1_N373, u1_N378, u1_N383, u1_N44, u1_N448, u1_N457, 
        u1_N467, u1_N473, u1_N49, u1_N59, u1_N65, u1_N7, u1_N76, u1_N81, u1_N91, 
        u1_N97, u2_N36, u2_N40, u2_N46, u2_N48, u2_N52, u2_N54, u2_N58, u2_N62;
  wire u0_K12_1, u0_K12_2, u0_K12_3, u0_K12_31, u0_K12_32, u0_K12_33, u0_K12_4, u0_K12_5, u0_K12_6, 
       u0_K2_19, u0_K2_20, u0_K2_21, u0_K2_22, u0_K2_23, u0_K2_24, u0_K3_25, u0_K3_26, u0_K3_27, 
       u0_K3_28, u0_K3_29, u0_K3_30, u0_K4_37, u0_K4_38, u0_K4_39, u0_K4_40, u0_K4_41, u0_K4_42, 
       u0_K4_44, u0_K4_45, u0_K4_46, u0_K4_47, u0_K6_1, u0_K6_10, u0_K6_12, u0_K6_14, u0_K6_15, 
       u0_K6_17, u0_K6_18, u0_K6_2, u0_K6_21, u0_K6_3, u0_K6_31, u0_K6_32, u0_K6_33, u0_K6_34, 
       u0_K6_35, u0_K6_36, u0_K6_4, u0_K6_43, u0_K6_44, u0_K6_45, u0_K6_46, u0_K6_47, u0_K6_48, 
       u0_K6_5, u0_K6_6, u0_K6_7, u0_K6_8, u0_K6_9, u0_K8_10, u0_K8_12, u0_K8_13, u0_K8_14, 
       u0_K8_15, u0_K8_16, u0_K8_17, u0_K8_18, u0_K8_2, u0_K8_20, u0_K8_21, u0_K8_22, u0_K8_23, 
       u0_K8_24, u0_K8_25, u0_K8_26, u0_K8_27, u0_K8_29, u0_K8_3, u0_K8_30, u0_K8_31, u0_K8_32, 
       u0_K8_34, u0_K8_35, u0_K8_37, u0_K8_38, u0_K8_39, u0_K8_4, u0_K8_40, u0_K8_41, u0_K8_42, 
       u0_K8_43, u0_K8_44, u0_K8_46, u0_K8_47, u0_K8_48, u0_K8_5, u0_K8_6, u0_K8_7, u0_K8_8, 
       u0_K8_9, u0_out11_11, u0_out11_17, u0_out11_19, u0_out11_23, u0_out11_29, u0_out11_31, u0_out11_4, u0_out11_9, 
       u0_out1_1, u0_out1_10, u0_out1_20, u0_out1_26, u0_out2_14, u0_out2_25, u0_out2_3, u0_out2_8, u0_out3_12, 
       u0_out3_15, u0_out3_21, u0_out3_22, u0_out3_27, u0_out3_32, u0_out3_5, u0_out3_7, u0_out5_1, u0_out5_10, 
       u0_out5_11, u0_out5_13, u0_out5_15, u0_out5_16, u0_out5_17, u0_out5_18, u0_out5_19, u0_out5_2, u0_out5_20, 
       u0_out5_21, u0_out5_23, u0_out5_24, u0_out5_26, u0_out5_27, u0_out5_28, u0_out5_29, u0_out5_30, u0_out5_31, 
       u0_out5_4, u0_out5_5, u0_out5_6, u0_out5_9, u0_out7_1, u0_out7_10, u0_out7_11, u0_out7_12, u0_out7_13, 
       u0_out7_14, u0_out7_15, u0_out7_16, u0_out7_17, u0_out7_18, u0_out7_19, u0_out7_2, u0_out7_20, u0_out7_21, 
       u0_out7_22, u0_out7_23, u0_out7_24, u0_out7_25, u0_out7_26, u0_out7_27, u0_out7_28, u0_out7_29, u0_out7_3, 
       u0_out7_30, u0_out7_31, u0_out7_32, u0_out7_4, u0_out7_5, u0_out7_6, u0_out7_7, u0_out7_8, u0_out7_9, 
       u0_u11_X_1, u0_u11_X_2, u0_u11_X_3, u0_u11_X_31, u0_u11_X_32, u0_u11_X_33, u0_u11_X_34, u0_u11_X_35, u0_u11_X_36, 
       u0_u11_X_4, u0_u11_X_5, u0_u11_X_6, u0_u11_u0_n100, u0_u11_u0_n101, u0_u11_u0_n102, u0_u11_u0_n103, u0_u11_u0_n104, u0_u11_u0_n105, 
       u0_u11_u0_n106, u0_u11_u0_n107, u0_u11_u0_n108, u0_u11_u0_n109, u0_u11_u0_n110, u0_u11_u0_n111, u0_u11_u0_n112, u0_u11_u0_n113, u0_u11_u0_n114, 
       u0_u11_u0_n115, u0_u11_u0_n116, u0_u11_u0_n117, u0_u11_u0_n118, u0_u11_u0_n119, u0_u11_u0_n120, u0_u11_u0_n121, u0_u11_u0_n122, u0_u11_u0_n123, 
       u0_u11_u0_n124, u0_u11_u0_n125, u0_u11_u0_n126, u0_u11_u0_n127, u0_u11_u0_n128, u0_u11_u0_n129, u0_u11_u0_n130, u0_u11_u0_n131, u0_u11_u0_n132, 
       u0_u11_u0_n133, u0_u11_u0_n134, u0_u11_u0_n135, u0_u11_u0_n136, u0_u11_u0_n137, u0_u11_u0_n138, u0_u11_u0_n139, u0_u11_u0_n140, u0_u11_u0_n141, 
       u0_u11_u0_n142, u0_u11_u0_n143, u0_u11_u0_n144, u0_u11_u0_n145, u0_u11_u0_n146, u0_u11_u0_n147, u0_u11_u0_n148, u0_u11_u0_n149, u0_u11_u0_n150, 
       u0_u11_u0_n151, u0_u11_u0_n152, u0_u11_u0_n153, u0_u11_u0_n154, u0_u11_u0_n155, u0_u11_u0_n156, u0_u11_u0_n157, u0_u11_u0_n158, u0_u11_u0_n159, 
       u0_u11_u0_n160, u0_u11_u0_n161, u0_u11_u0_n162, u0_u11_u0_n163, u0_u11_u0_n164, u0_u11_u0_n165, u0_u11_u0_n166, u0_u11_u0_n167, u0_u11_u0_n168, 
       u0_u11_u0_n169, u0_u11_u0_n170, u0_u11_u0_n171, u0_u11_u0_n172, u0_u11_u0_n173, u0_u11_u0_n174, u0_u11_u0_n88, u0_u11_u0_n89, u0_u11_u0_n90, 
       u0_u11_u0_n91, u0_u11_u0_n92, u0_u11_u0_n93, u0_u11_u0_n94, u0_u11_u0_n95, u0_u11_u0_n96, u0_u11_u0_n97, u0_u11_u0_n98, u0_u11_u0_n99, 
       u0_u11_u5_n100, u0_u11_u5_n101, u0_u11_u5_n102, u0_u11_u5_n103, u0_u11_u5_n104, u0_u11_u5_n105, u0_u11_u5_n106, u0_u11_u5_n107, u0_u11_u5_n108, 
       u0_u11_u5_n109, u0_u11_u5_n110, u0_u11_u5_n111, u0_u11_u5_n112, u0_u11_u5_n113, u0_u11_u5_n114, u0_u11_u5_n115, u0_u11_u5_n116, u0_u11_u5_n117, 
       u0_u11_u5_n118, u0_u11_u5_n119, u0_u11_u5_n120, u0_u11_u5_n121, u0_u11_u5_n122, u0_u11_u5_n123, u0_u11_u5_n124, u0_u11_u5_n125, u0_u11_u5_n126, 
       u0_u11_u5_n127, u0_u11_u5_n128, u0_u11_u5_n129, u0_u11_u5_n130, u0_u11_u5_n131, u0_u11_u5_n132, u0_u11_u5_n133, u0_u11_u5_n134, u0_u11_u5_n135, 
       u0_u11_u5_n136, u0_u11_u5_n137, u0_u11_u5_n138, u0_u11_u5_n139, u0_u11_u5_n140, u0_u11_u5_n141, u0_u11_u5_n142, u0_u11_u5_n143, u0_u11_u5_n144, 
       u0_u11_u5_n145, u0_u11_u5_n146, u0_u11_u5_n147, u0_u11_u5_n148, u0_u11_u5_n149, u0_u11_u5_n150, u0_u11_u5_n151, u0_u11_u5_n152, u0_u11_u5_n153, 
       u0_u11_u5_n154, u0_u11_u5_n155, u0_u11_u5_n156, u0_u11_u5_n157, u0_u11_u5_n158, u0_u11_u5_n159, u0_u11_u5_n160, u0_u11_u5_n161, u0_u11_u5_n162, 
       u0_u11_u5_n163, u0_u11_u5_n164, u0_u11_u5_n165, u0_u11_u5_n166, u0_u11_u5_n167, u0_u11_u5_n168, u0_u11_u5_n169, u0_u11_u5_n170, u0_u11_u5_n171, 
       u0_u11_u5_n172, u0_u11_u5_n173, u0_u11_u5_n174, u0_u11_u5_n175, u0_u11_u5_n176, u0_u11_u5_n177, u0_u11_u5_n178, u0_u11_u5_n179, u0_u11_u5_n180, 
       u0_u11_u5_n181, u0_u11_u5_n182, u0_u11_u5_n183, u0_u11_u5_n184, u0_u11_u5_n185, u0_u11_u5_n186, u0_u11_u5_n187, u0_u11_u5_n188, u0_u11_u5_n189, 
       u0_u11_u5_n190, u0_u11_u5_n191, u0_u11_u5_n192, u0_u11_u5_n193, u0_u11_u5_n194, u0_u11_u5_n195, u0_u11_u5_n196, u0_u11_u5_n99, u0_u1_X_19, 
       u0_u1_X_20, u0_u1_X_21, u0_u1_X_22, u0_u1_X_23, u0_u1_X_24, u0_u1_u3_n100, u0_u1_u3_n101, u0_u1_u3_n102, u0_u1_u3_n103, 
       u0_u1_u3_n104, u0_u1_u3_n105, u0_u1_u3_n106, u0_u1_u3_n107, u0_u1_u3_n108, u0_u1_u3_n109, u0_u1_u3_n110, u0_u1_u3_n111, u0_u1_u3_n112, 
       u0_u1_u3_n113, u0_u1_u3_n114, u0_u1_u3_n115, u0_u1_u3_n116, u0_u1_u3_n117, u0_u1_u3_n118, u0_u1_u3_n119, u0_u1_u3_n120, u0_u1_u3_n121, 
       u0_u1_u3_n122, u0_u1_u3_n123, u0_u1_u3_n124, u0_u1_u3_n125, u0_u1_u3_n126, u0_u1_u3_n127, u0_u1_u3_n128, u0_u1_u3_n129, u0_u1_u3_n130, 
       u0_u1_u3_n131, u0_u1_u3_n132, u0_u1_u3_n133, u0_u1_u3_n134, u0_u1_u3_n135, u0_u1_u3_n136, u0_u1_u3_n137, u0_u1_u3_n138, u0_u1_u3_n139, 
       u0_u1_u3_n140, u0_u1_u3_n141, u0_u1_u3_n142, u0_u1_u3_n143, u0_u1_u3_n144, u0_u1_u3_n145, u0_u1_u3_n146, u0_u1_u3_n147, u0_u1_u3_n148, 
       u0_u1_u3_n149, u0_u1_u3_n150, u0_u1_u3_n151, u0_u1_u3_n152, u0_u1_u3_n153, u0_u1_u3_n154, u0_u1_u3_n155, u0_u1_u3_n156, u0_u1_u3_n157, 
       u0_u1_u3_n158, u0_u1_u3_n159, u0_u1_u3_n160, u0_u1_u3_n161, u0_u1_u3_n162, u0_u1_u3_n163, u0_u1_u3_n164, u0_u1_u3_n165, u0_u1_u3_n166, 
       u0_u1_u3_n167, u0_u1_u3_n168, u0_u1_u3_n169, u0_u1_u3_n170, u0_u1_u3_n171, u0_u1_u3_n172, u0_u1_u3_n173, u0_u1_u3_n174, u0_u1_u3_n175, 
       u0_u1_u3_n176, u0_u1_u3_n177, u0_u1_u3_n178, u0_u1_u3_n179, u0_u1_u3_n180, u0_u1_u3_n181, u0_u1_u3_n182, u0_u1_u3_n183, u0_u1_u3_n184, 
       u0_u1_u3_n185, u0_u1_u3_n186, u0_u1_u3_n94, u0_u1_u3_n95, u0_u1_u3_n96, u0_u1_u3_n97, u0_u1_u3_n98, u0_u1_u3_n99, u0_u2_X_25, 
       u0_u2_X_26, u0_u2_X_27, u0_u2_X_28, u0_u2_X_29, u0_u2_X_30, u0_u2_u4_n100, u0_u2_u4_n101, u0_u2_u4_n102, u0_u2_u4_n103, 
       u0_u2_u4_n104, u0_u2_u4_n105, u0_u2_u4_n106, u0_u2_u4_n107, u0_u2_u4_n108, u0_u2_u4_n109, u0_u2_u4_n110, u0_u2_u4_n111, u0_u2_u4_n112, 
       u0_u2_u4_n113, u0_u2_u4_n114, u0_u2_u4_n115, u0_u2_u4_n116, u0_u2_u4_n117, u0_u2_u4_n118, u0_u2_u4_n119, u0_u2_u4_n120, u0_u2_u4_n121, 
       u0_u2_u4_n122, u0_u2_u4_n123, u0_u2_u4_n124, u0_u2_u4_n125, u0_u2_u4_n126, u0_u2_u4_n127, u0_u2_u4_n128, u0_u2_u4_n129, u0_u2_u4_n130, 
       u0_u2_u4_n131, u0_u2_u4_n132, u0_u2_u4_n133, u0_u2_u4_n134, u0_u2_u4_n135, u0_u2_u4_n136, u0_u2_u4_n137, u0_u2_u4_n138, u0_u2_u4_n139, 
       u0_u2_u4_n140, u0_u2_u4_n141, u0_u2_u4_n142, u0_u2_u4_n143, u0_u2_u4_n144, u0_u2_u4_n145, u0_u2_u4_n146, u0_u2_u4_n147, u0_u2_u4_n148, 
       u0_u2_u4_n149, u0_u2_u4_n150, u0_u2_u4_n151, u0_u2_u4_n152, u0_u2_u4_n153, u0_u2_u4_n154, u0_u2_u4_n155, u0_u2_u4_n156, u0_u2_u4_n157, 
       u0_u2_u4_n158, u0_u2_u4_n159, u0_u2_u4_n160, u0_u2_u4_n161, u0_u2_u4_n162, u0_u2_u4_n163, u0_u2_u4_n164, u0_u2_u4_n165, u0_u2_u4_n166, 
       u0_u2_u4_n167, u0_u2_u4_n168, u0_u2_u4_n169, u0_u2_u4_n170, u0_u2_u4_n171, u0_u2_u4_n172, u0_u2_u4_n173, u0_u2_u4_n174, u0_u2_u4_n175, 
       u0_u2_u4_n176, u0_u2_u4_n177, u0_u2_u4_n178, u0_u2_u4_n179, u0_u2_u4_n180, u0_u2_u4_n181, u0_u2_u4_n182, u0_u2_u4_n183, u0_u2_u4_n184, 
       u0_u2_u4_n185, u0_u2_u4_n186, u0_u2_u4_n94, u0_u2_u4_n95, u0_u2_u4_n96, u0_u2_u4_n97, u0_u2_u4_n98, u0_u2_u4_n99, u0_u3_X_37, 
       u0_u3_X_38, u0_u3_X_39, u0_u3_X_40, u0_u3_X_41, u0_u3_X_42, u0_u3_X_43, u0_u3_X_44, u0_u3_X_45, u0_u3_X_46, 
       u0_u3_X_47, u0_u3_X_48, u0_u3_u6_n100, u0_u3_u6_n101, u0_u3_u6_n102, u0_u3_u6_n103, u0_u3_u6_n104, u0_u3_u6_n105, u0_u3_u6_n106, 
       u0_u3_u6_n107, u0_u3_u6_n108, u0_u3_u6_n109, u0_u3_u6_n110, u0_u3_u6_n111, u0_u3_u6_n112, u0_u3_u6_n113, u0_u3_u6_n114, u0_u3_u6_n115, 
       u0_u3_u6_n116, u0_u3_u6_n117, u0_u3_u6_n118, u0_u3_u6_n119, u0_u3_u6_n120, u0_u3_u6_n121, u0_u3_u6_n122, u0_u3_u6_n123, u0_u3_u6_n124, 
       u0_u3_u6_n125, u0_u3_u6_n126, u0_u3_u6_n127, u0_u3_u6_n128, u0_u3_u6_n129, u0_u3_u6_n130, u0_u3_u6_n131, u0_u3_u6_n132, u0_u3_u6_n133, 
       u0_u3_u6_n134, u0_u3_u6_n135, u0_u3_u6_n136, u0_u3_u6_n137, u0_u3_u6_n138, u0_u3_u6_n139, u0_u3_u6_n140, u0_u3_u6_n141, u0_u3_u6_n142, 
       u0_u3_u6_n143, u0_u3_u6_n144, u0_u3_u6_n145, u0_u3_u6_n146, u0_u3_u6_n147, u0_u3_u6_n148, u0_u3_u6_n149, u0_u3_u6_n150, u0_u3_u6_n151, 
       u0_u3_u6_n152, u0_u3_u6_n153, u0_u3_u6_n154, u0_u3_u6_n155, u0_u3_u6_n156, u0_u3_u6_n157, u0_u3_u6_n158, u0_u3_u6_n159, u0_u3_u6_n160, 
       u0_u3_u6_n161, u0_u3_u6_n162, u0_u3_u6_n163, u0_u3_u6_n164, u0_u3_u6_n165, u0_u3_u6_n166, u0_u3_u6_n167, u0_u3_u6_n168, u0_u3_u6_n169, 
       u0_u3_u6_n170, u0_u3_u6_n171, u0_u3_u6_n172, u0_u3_u6_n173, u0_u3_u6_n174, u0_u3_u6_n88, u0_u3_u6_n89, u0_u3_u6_n90, u0_u3_u6_n91, 
       u0_u3_u6_n92, u0_u3_u6_n93, u0_u3_u6_n94, u0_u3_u6_n95, u0_u3_u6_n96, u0_u3_u6_n97, u0_u3_u6_n98, u0_u3_u6_n99, u0_u3_u7_n100, 
       u0_u3_u7_n101, u0_u3_u7_n102, u0_u3_u7_n103, u0_u3_u7_n104, u0_u3_u7_n105, u0_u3_u7_n106, u0_u3_u7_n107, u0_u3_u7_n108, u0_u3_u7_n109, 
       u0_u3_u7_n110, u0_u3_u7_n111, u0_u3_u7_n112, u0_u3_u7_n113, u0_u3_u7_n114, u0_u3_u7_n115, u0_u3_u7_n116, u0_u3_u7_n117, u0_u3_u7_n118, 
       u0_u3_u7_n119, u0_u3_u7_n120, u0_u3_u7_n121, u0_u3_u7_n122, u0_u3_u7_n123, u0_u3_u7_n124, u0_u3_u7_n125, u0_u3_u7_n126, u0_u3_u7_n127, 
       u0_u3_u7_n128, u0_u3_u7_n129, u0_u3_u7_n130, u0_u3_u7_n131, u0_u3_u7_n132, u0_u3_u7_n133, u0_u3_u7_n134, u0_u3_u7_n135, u0_u3_u7_n136, 
       u0_u3_u7_n137, u0_u3_u7_n138, u0_u3_u7_n139, u0_u3_u7_n140, u0_u3_u7_n141, u0_u3_u7_n142, u0_u3_u7_n143, u0_u3_u7_n144, u0_u3_u7_n145, 
       u0_u3_u7_n146, u0_u3_u7_n147, u0_u3_u7_n148, u0_u3_u7_n149, u0_u3_u7_n150, u0_u3_u7_n151, u0_u3_u7_n152, u0_u3_u7_n153, u0_u3_u7_n154, 
       u0_u3_u7_n155, u0_u3_u7_n156, u0_u3_u7_n157, u0_u3_u7_n158, u0_u3_u7_n159, u0_u3_u7_n160, u0_u3_u7_n161, u0_u3_u7_n162, u0_u3_u7_n163, 
       u0_u3_u7_n164, u0_u3_u7_n165, u0_u3_u7_n166, u0_u3_u7_n167, u0_u3_u7_n168, u0_u3_u7_n169, u0_u3_u7_n170, u0_u3_u7_n171, u0_u3_u7_n172, 
       u0_u3_u7_n173, u0_u3_u7_n174, u0_u3_u7_n175, u0_u3_u7_n176, u0_u3_u7_n177, u0_u3_u7_n178, u0_u3_u7_n179, u0_u3_u7_n180, u0_u3_u7_n91, 
       u0_u3_u7_n92, u0_u3_u7_n93, u0_u3_u7_n94, u0_u3_u7_n95, u0_u3_u7_n96, u0_u3_u7_n97, u0_u3_u7_n98, u0_u3_u7_n99, u0_u5_X_1, 
       u0_u5_X_10, u0_u5_X_11, u0_u5_X_12, u0_u5_X_13, u0_u5_X_14, u0_u5_X_15, u0_u5_X_16, u0_u5_X_17, u0_u5_X_18, 
       u0_u5_X_19, u0_u5_X_2, u0_u5_X_20, u0_u5_X_21, u0_u5_X_22, u0_u5_X_23, u0_u5_X_24, u0_u5_X_3, u0_u5_X_31, 
       u0_u5_X_32, u0_u5_X_33, u0_u5_X_34, u0_u5_X_35, u0_u5_X_36, u0_u5_X_4, u0_u5_X_43, u0_u5_X_44, u0_u5_X_45, 
       u0_u5_X_46, u0_u5_X_47, u0_u5_X_48, u0_u5_X_5, u0_u5_X_6, u0_u5_X_7, u0_u5_X_8, u0_u5_X_9, u0_u5_u0_n100, 
       u0_u5_u0_n101, u0_u5_u0_n102, u0_u5_u0_n103, u0_u5_u0_n104, u0_u5_u0_n105, u0_u5_u0_n106, u0_u5_u0_n107, u0_u5_u0_n108, u0_u5_u0_n109, 
       u0_u5_u0_n110, u0_u5_u0_n111, u0_u5_u0_n112, u0_u5_u0_n113, u0_u5_u0_n114, u0_u5_u0_n115, u0_u5_u0_n116, u0_u5_u0_n117, u0_u5_u0_n118, 
       u0_u5_u0_n119, u0_u5_u0_n120, u0_u5_u0_n121, u0_u5_u0_n122, u0_u5_u0_n123, u0_u5_u0_n124, u0_u5_u0_n125, u0_u5_u0_n126, u0_u5_u0_n127, 
       u0_u5_u0_n128, u0_u5_u0_n129, u0_u5_u0_n130, u0_u5_u0_n131, u0_u5_u0_n132, u0_u5_u0_n133, u0_u5_u0_n134, u0_u5_u0_n135, u0_u5_u0_n136, 
       u0_u5_u0_n137, u0_u5_u0_n138, u0_u5_u0_n139, u0_u5_u0_n140, u0_u5_u0_n141, u0_u5_u0_n142, u0_u5_u0_n143, u0_u5_u0_n144, u0_u5_u0_n145, 
       u0_u5_u0_n146, u0_u5_u0_n147, u0_u5_u0_n148, u0_u5_u0_n149, u0_u5_u0_n150, u0_u5_u0_n151, u0_u5_u0_n152, u0_u5_u0_n153, u0_u5_u0_n154, 
       u0_u5_u0_n155, u0_u5_u0_n156, u0_u5_u0_n157, u0_u5_u0_n158, u0_u5_u0_n159, u0_u5_u0_n160, u0_u5_u0_n161, u0_u5_u0_n162, u0_u5_u0_n163, 
       u0_u5_u0_n164, u0_u5_u0_n165, u0_u5_u0_n166, u0_u5_u0_n167, u0_u5_u0_n168, u0_u5_u0_n169, u0_u5_u0_n170, u0_u5_u0_n171, u0_u5_u0_n172, 
       u0_u5_u0_n173, u0_u5_u0_n174, u0_u5_u0_n88, u0_u5_u0_n89, u0_u5_u0_n90, u0_u5_u0_n91, u0_u5_u0_n92, u0_u5_u0_n93, u0_u5_u0_n94, 
       u0_u5_u0_n95, u0_u5_u0_n96, u0_u5_u0_n97, u0_u5_u0_n98, u0_u5_u0_n99, u0_u5_u1_n100, u0_u5_u1_n101, u0_u5_u1_n102, u0_u5_u1_n103, 
       u0_u5_u1_n104, u0_u5_u1_n105, u0_u5_u1_n106, u0_u5_u1_n107, u0_u5_u1_n108, u0_u5_u1_n109, u0_u5_u1_n110, u0_u5_u1_n111, u0_u5_u1_n112, 
       u0_u5_u1_n113, u0_u5_u1_n114, u0_u5_u1_n115, u0_u5_u1_n116, u0_u5_u1_n117, u0_u5_u1_n118, u0_u5_u1_n119, u0_u5_u1_n120, u0_u5_u1_n121, 
       u0_u5_u1_n122, u0_u5_u1_n123, u0_u5_u1_n124, u0_u5_u1_n125, u0_u5_u1_n126, u0_u5_u1_n127, u0_u5_u1_n128, u0_u5_u1_n129, u0_u5_u1_n130, 
       u0_u5_u1_n131, u0_u5_u1_n132, u0_u5_u1_n133, u0_u5_u1_n134, u0_u5_u1_n135, u0_u5_u1_n136, u0_u5_u1_n137, u0_u5_u1_n138, u0_u5_u1_n139, 
       u0_u5_u1_n140, u0_u5_u1_n141, u0_u5_u1_n142, u0_u5_u1_n143, u0_u5_u1_n144, u0_u5_u1_n145, u0_u5_u1_n146, u0_u5_u1_n147, u0_u5_u1_n148, 
       u0_u5_u1_n149, u0_u5_u1_n150, u0_u5_u1_n151, u0_u5_u1_n152, u0_u5_u1_n153, u0_u5_u1_n154, u0_u5_u1_n155, u0_u5_u1_n156, u0_u5_u1_n157, 
       u0_u5_u1_n158, u0_u5_u1_n159, u0_u5_u1_n160, u0_u5_u1_n161, u0_u5_u1_n162, u0_u5_u1_n163, u0_u5_u1_n164, u0_u5_u1_n165, u0_u5_u1_n166, 
       u0_u5_u1_n167, u0_u5_u1_n168, u0_u5_u1_n169, u0_u5_u1_n170, u0_u5_u1_n171, u0_u5_u1_n172, u0_u5_u1_n173, u0_u5_u1_n174, u0_u5_u1_n175, 
       u0_u5_u1_n176, u0_u5_u1_n177, u0_u5_u1_n178, u0_u5_u1_n179, u0_u5_u1_n180, u0_u5_u1_n181, u0_u5_u1_n182, u0_u5_u1_n183, u0_u5_u1_n184, 
       u0_u5_u1_n185, u0_u5_u1_n186, u0_u5_u1_n187, u0_u5_u1_n188, u0_u5_u1_n95, u0_u5_u1_n96, u0_u5_u1_n97, u0_u5_u1_n98, u0_u5_u1_n99, 
       u0_u5_u2_n100, u0_u5_u2_n101, u0_u5_u2_n102, u0_u5_u2_n103, u0_u5_u2_n104, u0_u5_u2_n105, u0_u5_u2_n106, u0_u5_u2_n107, u0_u5_u2_n108, 
       u0_u5_u2_n109, u0_u5_u2_n110, u0_u5_u2_n111, u0_u5_u2_n112, u0_u5_u2_n113, u0_u5_u2_n114, u0_u5_u2_n115, u0_u5_u2_n116, u0_u5_u2_n117, 
       u0_u5_u2_n118, u0_u5_u2_n119, u0_u5_u2_n120, u0_u5_u2_n121, u0_u5_u2_n122, u0_u5_u2_n123, u0_u5_u2_n124, u0_u5_u2_n125, u0_u5_u2_n126, 
       u0_u5_u2_n127, u0_u5_u2_n128, u0_u5_u2_n129, u0_u5_u2_n130, u0_u5_u2_n131, u0_u5_u2_n132, u0_u5_u2_n133, u0_u5_u2_n134, u0_u5_u2_n135, 
       u0_u5_u2_n136, u0_u5_u2_n137, u0_u5_u2_n138, u0_u5_u2_n139, u0_u5_u2_n140, u0_u5_u2_n141, u0_u5_u2_n142, u0_u5_u2_n143, u0_u5_u2_n144, 
       u0_u5_u2_n145, u0_u5_u2_n146, u0_u5_u2_n147, u0_u5_u2_n148, u0_u5_u2_n149, u0_u5_u2_n150, u0_u5_u2_n151, u0_u5_u2_n152, u0_u5_u2_n153, 
       u0_u5_u2_n154, u0_u5_u2_n155, u0_u5_u2_n156, u0_u5_u2_n157, u0_u5_u2_n158, u0_u5_u2_n159, u0_u5_u2_n160, u0_u5_u2_n161, u0_u5_u2_n162, 
       u0_u5_u2_n163, u0_u5_u2_n164, u0_u5_u2_n165, u0_u5_u2_n166, u0_u5_u2_n167, u0_u5_u2_n168, u0_u5_u2_n169, u0_u5_u2_n170, u0_u5_u2_n171, 
       u0_u5_u2_n172, u0_u5_u2_n173, u0_u5_u2_n174, u0_u5_u2_n175, u0_u5_u2_n176, u0_u5_u2_n177, u0_u5_u2_n178, u0_u5_u2_n179, u0_u5_u2_n180, 
       u0_u5_u2_n181, u0_u5_u2_n182, u0_u5_u2_n183, u0_u5_u2_n184, u0_u5_u2_n185, u0_u5_u2_n186, u0_u5_u2_n187, u0_u5_u2_n188, u0_u5_u2_n95, 
       u0_u5_u2_n96, u0_u5_u2_n97, u0_u5_u2_n98, u0_u5_u2_n99, u0_u5_u3_n100, u0_u5_u3_n101, u0_u5_u3_n102, u0_u5_u3_n103, u0_u5_u3_n104, 
       u0_u5_u3_n105, u0_u5_u3_n106, u0_u5_u3_n107, u0_u5_u3_n108, u0_u5_u3_n109, u0_u5_u3_n110, u0_u5_u3_n111, u0_u5_u3_n112, u0_u5_u3_n113, 
       u0_u5_u3_n114, u0_u5_u3_n115, u0_u5_u3_n116, u0_u5_u3_n117, u0_u5_u3_n118, u0_u5_u3_n119, u0_u5_u3_n120, u0_u5_u3_n121, u0_u5_u3_n122, 
       u0_u5_u3_n123, u0_u5_u3_n124, u0_u5_u3_n125, u0_u5_u3_n126, u0_u5_u3_n127, u0_u5_u3_n128, u0_u5_u3_n129, u0_u5_u3_n130, u0_u5_u3_n131, 
       u0_u5_u3_n132, u0_u5_u3_n133, u0_u5_u3_n134, u0_u5_u3_n135, u0_u5_u3_n136, u0_u5_u3_n137, u0_u5_u3_n138, u0_u5_u3_n139, u0_u5_u3_n140, 
       u0_u5_u3_n141, u0_u5_u3_n142, u0_u5_u3_n143, u0_u5_u3_n144, u0_u5_u3_n145, u0_u5_u3_n146, u0_u5_u3_n147, u0_u5_u3_n148, u0_u5_u3_n149, 
       u0_u5_u3_n150, u0_u5_u3_n151, u0_u5_u3_n152, u0_u5_u3_n153, u0_u5_u3_n154, u0_u5_u3_n155, u0_u5_u3_n156, u0_u5_u3_n157, u0_u5_u3_n158, 
       u0_u5_u3_n159, u0_u5_u3_n160, u0_u5_u3_n161, u0_u5_u3_n162, u0_u5_u3_n163, u0_u5_u3_n164, u0_u5_u3_n165, u0_u5_u3_n166, u0_u5_u3_n167, 
       u0_u5_u3_n168, u0_u5_u3_n169, u0_u5_u3_n170, u0_u5_u3_n171, u0_u5_u3_n172, u0_u5_u3_n173, u0_u5_u3_n174, u0_u5_u3_n175, u0_u5_u3_n176, 
       u0_u5_u3_n177, u0_u5_u3_n178, u0_u5_u3_n179, u0_u5_u3_n180, u0_u5_u3_n181, u0_u5_u3_n182, u0_u5_u3_n183, u0_u5_u3_n184, u0_u5_u3_n185, 
       u0_u5_u3_n186, u0_u5_u3_n94, u0_u5_u3_n95, u0_u5_u3_n96, u0_u5_u3_n97, u0_u5_u3_n98, u0_u5_u3_n99, u0_u5_u5_n100, u0_u5_u5_n101, 
       u0_u5_u5_n102, u0_u5_u5_n103, u0_u5_u5_n104, u0_u5_u5_n105, u0_u5_u5_n106, u0_u5_u5_n107, u0_u5_u5_n108, u0_u5_u5_n109, u0_u5_u5_n110, 
       u0_u5_u5_n111, u0_u5_u5_n112, u0_u5_u5_n113, u0_u5_u5_n114, u0_u5_u5_n115, u0_u5_u5_n116, u0_u5_u5_n117, u0_u5_u5_n118, u0_u5_u5_n119, 
       u0_u5_u5_n120, u0_u5_u5_n121, u0_u5_u5_n122, u0_u5_u5_n123, u0_u5_u5_n124, u0_u5_u5_n125, u0_u5_u5_n126, u0_u5_u5_n127, u0_u5_u5_n128, 
       u0_u5_u5_n129, u0_u5_u5_n130, u0_u5_u5_n131, u0_u5_u5_n132, u0_u5_u5_n133, u0_u5_u5_n134, u0_u5_u5_n135, u0_u5_u5_n136, u0_u5_u5_n137, 
       u0_u5_u5_n138, u0_u5_u5_n139, u0_u5_u5_n140, u0_u5_u5_n141, u0_u5_u5_n142, u0_u5_u5_n143, u0_u5_u5_n144, u0_u5_u5_n145, u0_u5_u5_n146, 
       u0_u5_u5_n147, u0_u5_u5_n148, u0_u5_u5_n149, u0_u5_u5_n150, u0_u5_u5_n151, u0_u5_u5_n152, u0_u5_u5_n153, u0_u5_u5_n154, u0_u5_u5_n155, 
       u0_u5_u5_n156, u0_u5_u5_n157, u0_u5_u5_n158, u0_u5_u5_n159, u0_u5_u5_n160, u0_u5_u5_n161, u0_u5_u5_n162, u0_u5_u5_n163, u0_u5_u5_n164, 
       u0_u5_u5_n165, u0_u5_u5_n166, u0_u5_u5_n167, u0_u5_u5_n168, u0_u5_u5_n169, u0_u5_u5_n170, u0_u5_u5_n171, u0_u5_u5_n172, u0_u5_u5_n173, 
       u0_u5_u5_n174, u0_u5_u5_n175, u0_u5_u5_n176, u0_u5_u5_n177, u0_u5_u5_n178, u0_u5_u5_n179, u0_u5_u5_n180, u0_u5_u5_n181, u0_u5_u5_n182, 
       u0_u5_u5_n183, u0_u5_u5_n184, u0_u5_u5_n185, u0_u5_u5_n186, u0_u5_u5_n187, u0_u5_u5_n188, u0_u5_u5_n189, u0_u5_u5_n190, u0_u5_u5_n191, 
       u0_u5_u5_n192, u0_u5_u5_n193, u0_u5_u5_n194, u0_u5_u5_n195, u0_u5_u5_n196, u0_u5_u5_n99, u0_u5_u7_n100, u0_u5_u7_n101, u0_u5_u7_n102, 
       u0_u5_u7_n103, u0_u5_u7_n104, u0_u5_u7_n105, u0_u5_u7_n106, u0_u5_u7_n107, u0_u5_u7_n108, u0_u5_u7_n109, u0_u5_u7_n110, u0_u5_u7_n111, 
       u0_u5_u7_n112, u0_u5_u7_n113, u0_u5_u7_n114, u0_u5_u7_n115, u0_u5_u7_n116, u0_u5_u7_n117, u0_u5_u7_n118, u0_u5_u7_n119, u0_u5_u7_n120, 
       u0_u5_u7_n121, u0_u5_u7_n122, u0_u5_u7_n123, u0_u5_u7_n124, u0_u5_u7_n125, u0_u5_u7_n126, u0_u5_u7_n127, u0_u5_u7_n128, u0_u5_u7_n129, 
       u0_u5_u7_n130, u0_u5_u7_n131, u0_u5_u7_n132, u0_u5_u7_n133, u0_u5_u7_n134, u0_u5_u7_n135, u0_u5_u7_n136, u0_u5_u7_n137, u0_u5_u7_n138, 
       u0_u5_u7_n139, u0_u5_u7_n140, u0_u5_u7_n141, u0_u5_u7_n142, u0_u5_u7_n143, u0_u5_u7_n144, u0_u5_u7_n145, u0_u5_u7_n146, u0_u5_u7_n147, 
       u0_u5_u7_n148, u0_u5_u7_n149, u0_u5_u7_n150, u0_u5_u7_n151, u0_u5_u7_n152, u0_u5_u7_n153, u0_u5_u7_n154, u0_u5_u7_n155, u0_u5_u7_n156, 
       u0_u5_u7_n157, u0_u5_u7_n158, u0_u5_u7_n159, u0_u5_u7_n160, u0_u5_u7_n161, u0_u5_u7_n162, u0_u5_u7_n163, u0_u5_u7_n164, u0_u5_u7_n165, 
       u0_u5_u7_n166, u0_u5_u7_n167, u0_u5_u7_n168, u0_u5_u7_n169, u0_u5_u7_n170, u0_u5_u7_n171, u0_u5_u7_n172, u0_u5_u7_n173, u0_u5_u7_n174, 
       u0_u5_u7_n175, u0_u5_u7_n176, u0_u5_u7_n177, u0_u5_u7_n178, u0_u5_u7_n179, u0_u5_u7_n180, u0_u5_u7_n91, u0_u5_u7_n92, u0_u5_u7_n93, 
       u0_u5_u7_n94, u0_u5_u7_n95, u0_u5_u7_n96, u0_u5_u7_n97, u0_u5_u7_n98, u0_u5_u7_n99, u0_u7_X_1, u0_u7_X_10, u0_u7_X_11, 
       u0_u7_X_12, u0_u7_X_13, u0_u7_X_14, u0_u7_X_15, u0_u7_X_16, u0_u7_X_17, u0_u7_X_18, u0_u7_X_19, u0_u7_X_2, 
       u0_u7_X_20, u0_u7_X_21, u0_u7_X_22, u0_u7_X_23, u0_u7_X_24, u0_u7_X_25, u0_u7_X_26, u0_u7_X_27, u0_u7_X_28, 
       u0_u7_X_29, u0_u7_X_3, u0_u7_X_30, u0_u7_X_31, u0_u7_X_32, u0_u7_X_33, u0_u7_X_34, u0_u7_X_35, u0_u7_X_36, 
       u0_u7_X_37, u0_u7_X_38, u0_u7_X_39, u0_u7_X_4, u0_u7_X_40, u0_u7_X_41, u0_u7_X_42, u0_u7_X_43, u0_u7_X_44, 
       u0_u7_X_45, u0_u7_X_46, u0_u7_X_47, u0_u7_X_48, u0_u7_X_5, u0_u7_X_6, u0_u7_X_7, u0_u7_X_8, u0_u7_X_9, 
       u0_u7_u0_n100, u0_u7_u0_n101, u0_u7_u0_n102, u0_u7_u0_n103, u0_u7_u0_n104, u0_u7_u0_n105, u0_u7_u0_n106, u0_u7_u0_n107, u0_u7_u0_n108, 
       u0_u7_u0_n109, u0_u7_u0_n110, u0_u7_u0_n111, u0_u7_u0_n112, u0_u7_u0_n113, u0_u7_u0_n114, u0_u7_u0_n115, u0_u7_u0_n116, u0_u7_u0_n117, 
       u0_u7_u0_n118, u0_u7_u0_n119, u0_u7_u0_n120, u0_u7_u0_n121, u0_u7_u0_n122, u0_u7_u0_n123, u0_u7_u0_n124, u0_u7_u0_n125, u0_u7_u0_n126, 
       u0_u7_u0_n127, u0_u7_u0_n128, u0_u7_u0_n129, u0_u7_u0_n130, u0_u7_u0_n131, u0_u7_u0_n132, u0_u7_u0_n133, u0_u7_u0_n134, u0_u7_u0_n135, 
       u0_u7_u0_n136, u0_u7_u0_n137, u0_u7_u0_n138, u0_u7_u0_n139, u0_u7_u0_n140, u0_u7_u0_n141, u0_u7_u0_n142, u0_u7_u0_n143, u0_u7_u0_n144, 
       u0_u7_u0_n145, u0_u7_u0_n146, u0_u7_u0_n147, u0_u7_u0_n148, u0_u7_u0_n149, u0_u7_u0_n150, u0_u7_u0_n151, u0_u7_u0_n152, u0_u7_u0_n153, 
       u0_u7_u0_n154, u0_u7_u0_n155, u0_u7_u0_n156, u0_u7_u0_n157, u0_u7_u0_n158, u0_u7_u0_n159, u0_u7_u0_n160, u0_u7_u0_n161, u0_u7_u0_n162, 
       u0_u7_u0_n163, u0_u7_u0_n164, u0_u7_u0_n165, u0_u7_u0_n166, u0_u7_u0_n167, u0_u7_u0_n168, u0_u7_u0_n169, u0_u7_u0_n170, u0_u7_u0_n171, 
       u0_u7_u0_n172, u0_u7_u0_n173, u0_u7_u0_n174, u0_u7_u0_n88, u0_u7_u0_n89, u0_u7_u0_n90, u0_u7_u0_n91, u0_u7_u0_n92, u0_u7_u0_n93, 
       u0_u7_u0_n94, u0_u7_u0_n95, u0_u7_u0_n96, u0_u7_u0_n97, u0_u7_u0_n98, u0_u7_u0_n99, u0_u7_u1_n100, u0_u7_u1_n101, u0_u7_u1_n102, 
       u0_u7_u1_n103, u0_u7_u1_n104, u0_u7_u1_n105, u0_u7_u1_n106, u0_u7_u1_n107, u0_u7_u1_n108, u0_u7_u1_n109, u0_u7_u1_n110, u0_u7_u1_n111, 
       u0_u7_u1_n112, u0_u7_u1_n113, u0_u7_u1_n114, u0_u7_u1_n115, u0_u7_u1_n116, u0_u7_u1_n117, u0_u7_u1_n118, u0_u7_u1_n119, u0_u7_u1_n120, 
       u0_u7_u1_n121, u0_u7_u1_n122, u0_u7_u1_n123, u0_u7_u1_n124, u0_u7_u1_n125, u0_u7_u1_n126, u0_u7_u1_n127, u0_u7_u1_n128, u0_u7_u1_n129, 
       u0_u7_u1_n130, u0_u7_u1_n131, u0_u7_u1_n132, u0_u7_u1_n133, u0_u7_u1_n134, u0_u7_u1_n135, u0_u7_u1_n136, u0_u7_u1_n137, u0_u7_u1_n138, 
       u0_u7_u1_n139, u0_u7_u1_n140, u0_u7_u1_n141, u0_u7_u1_n142, u0_u7_u1_n143, u0_u7_u1_n144, u0_u7_u1_n145, u0_u7_u1_n146, u0_u7_u1_n147, 
       u0_u7_u1_n148, u0_u7_u1_n149, u0_u7_u1_n150, u0_u7_u1_n151, u0_u7_u1_n152, u0_u7_u1_n153, u0_u7_u1_n154, u0_u7_u1_n155, u0_u7_u1_n156, 
       u0_u7_u1_n157, u0_u7_u1_n158, u0_u7_u1_n159, u0_u7_u1_n160, u0_u7_u1_n161, u0_u7_u1_n162, u0_u7_u1_n163, u0_u7_u1_n164, u0_u7_u1_n165, 
       u0_u7_u1_n166, u0_u7_u1_n167, u0_u7_u1_n168, u0_u7_u1_n169, u0_u7_u1_n170, u0_u7_u1_n171, u0_u7_u1_n172, u0_u7_u1_n173, u0_u7_u1_n174, 
       u0_u7_u1_n175, u0_u7_u1_n176, u0_u7_u1_n177, u0_u7_u1_n178, u0_u7_u1_n179, u0_u7_u1_n180, u0_u7_u1_n181, u0_u7_u1_n182, u0_u7_u1_n183, 
       u0_u7_u1_n184, u0_u7_u1_n185, u0_u7_u1_n186, u0_u7_u1_n187, u0_u7_u1_n188, u0_u7_u1_n95, u0_u7_u1_n96, u0_u7_u1_n97, u0_u7_u1_n98, 
       u0_u7_u1_n99, u0_u7_u2_n100, u0_u7_u2_n101, u0_u7_u2_n102, u0_u7_u2_n103, u0_u7_u2_n104, u0_u7_u2_n105, u0_u7_u2_n106, u0_u7_u2_n107, 
       u0_u7_u2_n108, u0_u7_u2_n109, u0_u7_u2_n110, u0_u7_u2_n111, u0_u7_u2_n112, u0_u7_u2_n113, u0_u7_u2_n114, u0_u7_u2_n115, u0_u7_u2_n116, 
       u0_u7_u2_n117, u0_u7_u2_n118, u0_u7_u2_n119, u0_u7_u2_n120, u0_u7_u2_n121, u0_u7_u2_n122, u0_u7_u2_n123, u0_u7_u2_n124, u0_u7_u2_n125, 
       u0_u7_u2_n126, u0_u7_u2_n127, u0_u7_u2_n128, u0_u7_u2_n129, u0_u7_u2_n130, u0_u7_u2_n131, u0_u7_u2_n132, u0_u7_u2_n133, u0_u7_u2_n134, 
       u0_u7_u2_n135, u0_u7_u2_n136, u0_u7_u2_n137, u0_u7_u2_n138, u0_u7_u2_n139, u0_u7_u2_n140, u0_u7_u2_n141, u0_u7_u2_n142, u0_u7_u2_n143, 
       u0_u7_u2_n144, u0_u7_u2_n145, u0_u7_u2_n146, u0_u7_u2_n147, u0_u7_u2_n148, u0_u7_u2_n149, u0_u7_u2_n150, u0_u7_u2_n151, u0_u7_u2_n152, 
       u0_u7_u2_n153, u0_u7_u2_n154, u0_u7_u2_n155, u0_u7_u2_n156, u0_u7_u2_n157, u0_u7_u2_n158, u0_u7_u2_n159, u0_u7_u2_n160, u0_u7_u2_n161, 
       u0_u7_u2_n162, u0_u7_u2_n163, u0_u7_u2_n164, u0_u7_u2_n165, u0_u7_u2_n166, u0_u7_u2_n167, u0_u7_u2_n168, u0_u7_u2_n169, u0_u7_u2_n170, 
       u0_u7_u2_n171, u0_u7_u2_n172, u0_u7_u2_n173, u0_u7_u2_n174, u0_u7_u2_n175, u0_u7_u2_n176, u0_u7_u2_n177, u0_u7_u2_n178, u0_u7_u2_n179, 
       u0_u7_u2_n180, u0_u7_u2_n181, u0_u7_u2_n182, u0_u7_u2_n183, u0_u7_u2_n184, u0_u7_u2_n185, u0_u7_u2_n186, u0_u7_u2_n187, u0_u7_u2_n188, 
       u0_u7_u2_n95, u0_u7_u2_n96, u0_u7_u2_n97, u0_u7_u2_n98, u0_u7_u2_n99, u0_u7_u3_n100, u0_u7_u3_n101, u0_u7_u3_n102, u0_u7_u3_n103, 
       u0_u7_u3_n104, u0_u7_u3_n105, u0_u7_u3_n106, u0_u7_u3_n107, u0_u7_u3_n108, u0_u7_u3_n109, u0_u7_u3_n110, u0_u7_u3_n111, u0_u7_u3_n112, 
       u0_u7_u3_n113, u0_u7_u3_n114, u0_u7_u3_n115, u0_u7_u3_n116, u0_u7_u3_n117, u0_u7_u3_n118, u0_u7_u3_n119, u0_u7_u3_n120, u0_u7_u3_n121, 
       u0_u7_u3_n122, u0_u7_u3_n123, u0_u7_u3_n124, u0_u7_u3_n125, u0_u7_u3_n126, u0_u7_u3_n127, u0_u7_u3_n128, u0_u7_u3_n129, u0_u7_u3_n130, 
       u0_u7_u3_n131, u0_u7_u3_n132, u0_u7_u3_n133, u0_u7_u3_n134, u0_u7_u3_n135, u0_u7_u3_n136, u0_u7_u3_n137, u0_u7_u3_n138, u0_u7_u3_n139, 
       u0_u7_u3_n140, u0_u7_u3_n141, u0_u7_u3_n142, u0_u7_u3_n143, u0_u7_u3_n144, u0_u7_u3_n145, u0_u7_u3_n146, u0_u7_u3_n147, u0_u7_u3_n148, 
       u0_u7_u3_n149, u0_u7_u3_n150, u0_u7_u3_n151, u0_u7_u3_n152, u0_u7_u3_n153, u0_u7_u3_n154, u0_u7_u3_n155, u0_u7_u3_n156, u0_u7_u3_n157, 
       u0_u7_u3_n158, u0_u7_u3_n159, u0_u7_u3_n160, u0_u7_u3_n161, u0_u7_u3_n162, u0_u7_u3_n163, u0_u7_u3_n164, u0_u7_u3_n165, u0_u7_u3_n166, 
       u0_u7_u3_n167, u0_u7_u3_n168, u0_u7_u3_n169, u0_u7_u3_n170, u0_u7_u3_n171, u0_u7_u3_n172, u0_u7_u3_n173, u0_u7_u3_n174, u0_u7_u3_n175, 
       u0_u7_u3_n176, u0_u7_u3_n177, u0_u7_u3_n178, u0_u7_u3_n179, u0_u7_u3_n180, u0_u7_u3_n181, u0_u7_u3_n182, u0_u7_u3_n183, u0_u7_u3_n184, 
       u0_u7_u3_n185, u0_u7_u3_n186, u0_u7_u3_n94, u0_u7_u3_n95, u0_u7_u3_n96, u0_u7_u3_n97, u0_u7_u3_n98, u0_u7_u3_n99, u0_u7_u4_n100, 
       u0_u7_u4_n101, u0_u7_u4_n102, u0_u7_u4_n103, u0_u7_u4_n104, u0_u7_u4_n105, u0_u7_u4_n106, u0_u7_u4_n107, u0_u7_u4_n108, u0_u7_u4_n109, 
       u0_u7_u4_n110, u0_u7_u4_n111, u0_u7_u4_n112, u0_u7_u4_n113, u0_u7_u4_n114, u0_u7_u4_n115, u0_u7_u4_n116, u0_u7_u4_n117, u0_u7_u4_n118, 
       u0_u7_u4_n119, u0_u7_u4_n120, u0_u7_u4_n121, u0_u7_u4_n122, u0_u7_u4_n123, u0_u7_u4_n124, u0_u7_u4_n125, u0_u7_u4_n126, u0_u7_u4_n127, 
       u0_u7_u4_n128, u0_u7_u4_n129, u0_u7_u4_n130, u0_u7_u4_n131, u0_u7_u4_n132, u0_u7_u4_n133, u0_u7_u4_n134, u0_u7_u4_n135, u0_u7_u4_n136, 
       u0_u7_u4_n137, u0_u7_u4_n138, u0_u7_u4_n139, u0_u7_u4_n140, u0_u7_u4_n141, u0_u7_u4_n142, u0_u7_u4_n143, u0_u7_u4_n144, u0_u7_u4_n145, 
       u0_u7_u4_n146, u0_u7_u4_n147, u0_u7_u4_n148, u0_u7_u4_n149, u0_u7_u4_n150, u0_u7_u4_n151, u0_u7_u4_n152, u0_u7_u4_n153, u0_u7_u4_n154, 
       u0_u7_u4_n155, u0_u7_u4_n156, u0_u7_u4_n157, u0_u7_u4_n158, u0_u7_u4_n159, u0_u7_u4_n160, u0_u7_u4_n161, u0_u7_u4_n162, u0_u7_u4_n163, 
       u0_u7_u4_n164, u0_u7_u4_n165, u0_u7_u4_n166, u0_u7_u4_n167, u0_u7_u4_n168, u0_u7_u4_n169, u0_u7_u4_n170, u0_u7_u4_n171, u0_u7_u4_n172, 
       u0_u7_u4_n173, u0_u7_u4_n174, u0_u7_u4_n175, u0_u7_u4_n176, u0_u7_u4_n177, u0_u7_u4_n178, u0_u7_u4_n179, u0_u7_u4_n180, u0_u7_u4_n181, 
       u0_u7_u4_n182, u0_u7_u4_n183, u0_u7_u4_n184, u0_u7_u4_n185, u0_u7_u4_n186, u0_u7_u4_n94, u0_u7_u4_n95, u0_u7_u4_n96, u0_u7_u4_n97, 
       u0_u7_u4_n98, u0_u7_u4_n99, u0_u7_u5_n100, u0_u7_u5_n101, u0_u7_u5_n102, u0_u7_u5_n103, u0_u7_u5_n104, u0_u7_u5_n105, u0_u7_u5_n106, 
       u0_u7_u5_n107, u0_u7_u5_n108, u0_u7_u5_n109, u0_u7_u5_n110, u0_u7_u5_n111, u0_u7_u5_n112, u0_u7_u5_n113, u0_u7_u5_n114, u0_u7_u5_n115, 
       u0_u7_u5_n116, u0_u7_u5_n117, u0_u7_u5_n118, u0_u7_u5_n119, u0_u7_u5_n120, u0_u7_u5_n121, u0_u7_u5_n122, u0_u7_u5_n123, u0_u7_u5_n124, 
       u0_u7_u5_n125, u0_u7_u5_n126, u0_u7_u5_n127, u0_u7_u5_n128, u0_u7_u5_n129, u0_u7_u5_n130, u0_u7_u5_n131, u0_u7_u5_n132, u0_u7_u5_n133, 
       u0_u7_u5_n134, u0_u7_u5_n135, u0_u7_u5_n136, u0_u7_u5_n137, u0_u7_u5_n138, u0_u7_u5_n139, u0_u7_u5_n140, u0_u7_u5_n141, u0_u7_u5_n142, 
       u0_u7_u5_n143, u0_u7_u5_n144, u0_u7_u5_n145, u0_u7_u5_n146, u0_u7_u5_n147, u0_u7_u5_n148, u0_u7_u5_n149, u0_u7_u5_n150, u0_u7_u5_n151, 
       u0_u7_u5_n152, u0_u7_u5_n153, u0_u7_u5_n154, u0_u7_u5_n155, u0_u7_u5_n156, u0_u7_u5_n157, u0_u7_u5_n158, u0_u7_u5_n159, u0_u7_u5_n160, 
       u0_u7_u5_n161, u0_u7_u5_n162, u0_u7_u5_n163, u0_u7_u5_n164, u0_u7_u5_n165, u0_u7_u5_n166, u0_u7_u5_n167, u0_u7_u5_n168, u0_u7_u5_n169, 
       u0_u7_u5_n170, u0_u7_u5_n171, u0_u7_u5_n172, u0_u7_u5_n173, u0_u7_u5_n174, u0_u7_u5_n175, u0_u7_u5_n176, u0_u7_u5_n177, u0_u7_u5_n178, 
       u0_u7_u5_n179, u0_u7_u5_n180, u0_u7_u5_n181, u0_u7_u5_n182, u0_u7_u5_n183, u0_u7_u5_n184, u0_u7_u5_n185, u0_u7_u5_n186, u0_u7_u5_n187, 
       u0_u7_u5_n188, u0_u7_u5_n189, u0_u7_u5_n190, u0_u7_u5_n191, u0_u7_u5_n192, u0_u7_u5_n193, u0_u7_u5_n194, u0_u7_u5_n195, u0_u7_u5_n196, 
       u0_u7_u5_n99, u0_u7_u6_n100, u0_u7_u6_n101, u0_u7_u6_n102, u0_u7_u6_n103, u0_u7_u6_n104, u0_u7_u6_n105, u0_u7_u6_n106, u0_u7_u6_n107, 
       u0_u7_u6_n108, u0_u7_u6_n109, u0_u7_u6_n110, u0_u7_u6_n111, u0_u7_u6_n112, u0_u7_u6_n113, u0_u7_u6_n114, u0_u7_u6_n115, u0_u7_u6_n116, 
       u0_u7_u6_n117, u0_u7_u6_n118, u0_u7_u6_n119, u0_u7_u6_n120, u0_u7_u6_n121, u0_u7_u6_n122, u0_u7_u6_n123, u0_u7_u6_n124, u0_u7_u6_n125, 
       u0_u7_u6_n126, u0_u7_u6_n127, u0_u7_u6_n128, u0_u7_u6_n129, u0_u7_u6_n130, u0_u7_u6_n131, u0_u7_u6_n132, u0_u7_u6_n133, u0_u7_u6_n134, 
       u0_u7_u6_n135, u0_u7_u6_n136, u0_u7_u6_n137, u0_u7_u6_n138, u0_u7_u6_n139, u0_u7_u6_n140, u0_u7_u6_n141, u0_u7_u6_n142, u0_u7_u6_n143, 
       u0_u7_u6_n144, u0_u7_u6_n145, u0_u7_u6_n146, u0_u7_u6_n147, u0_u7_u6_n148, u0_u7_u6_n149, u0_u7_u6_n150, u0_u7_u6_n151, u0_u7_u6_n152, 
       u0_u7_u6_n153, u0_u7_u6_n154, u0_u7_u6_n155, u0_u7_u6_n156, u0_u7_u6_n157, u0_u7_u6_n158, u0_u7_u6_n159, u0_u7_u6_n160, u0_u7_u6_n161, 
       u0_u7_u6_n162, u0_u7_u6_n163, u0_u7_u6_n164, u0_u7_u6_n165, u0_u7_u6_n166, u0_u7_u6_n167, u0_u7_u6_n168, u0_u7_u6_n169, u0_u7_u6_n170, 
       u0_u7_u6_n171, u0_u7_u6_n172, u0_u7_u6_n173, u0_u7_u6_n174, u0_u7_u6_n88, u0_u7_u6_n89, u0_u7_u6_n90, u0_u7_u6_n91, u0_u7_u6_n92, 
       u0_u7_u6_n93, u0_u7_u6_n94, u0_u7_u6_n95, u0_u7_u6_n96, u0_u7_u6_n97, u0_u7_u6_n98, u0_u7_u6_n99, u0_u7_u7_n100, u0_u7_u7_n101, 
       u0_u7_u7_n102, u0_u7_u7_n103, u0_u7_u7_n104, u0_u7_u7_n105, u0_u7_u7_n106, u0_u7_u7_n107, u0_u7_u7_n108, u0_u7_u7_n109, u0_u7_u7_n110, 
       u0_u7_u7_n111, u0_u7_u7_n112, u0_u7_u7_n113, u0_u7_u7_n114, u0_u7_u7_n115, u0_u7_u7_n116, u0_u7_u7_n117, u0_u7_u7_n118, u0_u7_u7_n119, 
       u0_u7_u7_n120, u0_u7_u7_n121, u0_u7_u7_n122, u0_u7_u7_n123, u0_u7_u7_n124, u0_u7_u7_n125, u0_u7_u7_n126, u0_u7_u7_n127, u0_u7_u7_n128, 
       u0_u7_u7_n129, u0_u7_u7_n130, u0_u7_u7_n131, u0_u7_u7_n132, u0_u7_u7_n133, u0_u7_u7_n134, u0_u7_u7_n135, u0_u7_u7_n136, u0_u7_u7_n137, 
       u0_u7_u7_n138, u0_u7_u7_n139, u0_u7_u7_n140, u0_u7_u7_n141, u0_u7_u7_n142, u0_u7_u7_n143, u0_u7_u7_n144, u0_u7_u7_n145, u0_u7_u7_n146, 
       u0_u7_u7_n147, u0_u7_u7_n148, u0_u7_u7_n149, u0_u7_u7_n150, u0_u7_u7_n151, u0_u7_u7_n152, u0_u7_u7_n153, u0_u7_u7_n154, u0_u7_u7_n155, 
       u0_u7_u7_n156, u0_u7_u7_n157, u0_u7_u7_n158, u0_u7_u7_n159, u0_u7_u7_n160, u0_u7_u7_n161, u0_u7_u7_n162, u0_u7_u7_n163, u0_u7_u7_n164, 
       u0_u7_u7_n165, u0_u7_u7_n166, u0_u7_u7_n167, u0_u7_u7_n168, u0_u7_u7_n169, u0_u7_u7_n170, u0_u7_u7_n171, u0_u7_u7_n172, u0_u7_u7_n173, 
       u0_u7_u7_n174, u0_u7_u7_n175, u0_u7_u7_n176, u0_u7_u7_n177, u0_u7_u7_n178, u0_u7_u7_n179, u0_u7_u7_n180, u0_u7_u7_n91, u0_u7_u7_n92, 
       u0_u7_u7_n93, u0_u7_u7_n94, u0_u7_u7_n95, u0_u7_u7_n96, u0_u7_u7_n97, u0_u7_u7_n98, u0_u7_u7_n99, u0_uk_n743, u0_uk_n744, 
       u0_uk_n745, u0_uk_n747, u0_uk_n749, u0_uk_n750, u0_uk_n751, u0_uk_n752, u0_uk_n753, u0_uk_n754, u0_uk_n757, 
       u0_uk_n758, u0_uk_n760, u0_uk_n761, u0_uk_n787, u0_uk_n788, u0_uk_n789, u0_uk_n792, u0_uk_n797, u0_uk_n800, 
       u0_uk_n801, u0_uk_n825, u0_uk_n849, u0_uk_n850, u0_uk_n864, u0_uk_n962, u0_uk_n968, u0_uk_n971, u0_uk_n972, 
       u0_uk_n973, u0_uk_n978, u1_K10_12, u1_K10_22, u1_K10_33, u1_K10_35, u1_K10_37, u1_K10_38, u1_K10_39, 
       u1_K10_40, u1_K10_9, u1_K16_34, u1_K1_27, u1_K1_33, u1_K2_10, u1_K4_10, u1_K7_46, u1_out0_11, 
       u1_out0_14, u1_out0_19, u1_out0_25, u1_out0_29, u1_out0_3, u1_out0_4, u1_out0_8, u1_out11_12, u1_out11_15, 
       u1_out11_21, u1_out11_22, u1_out11_27, u1_out11_32, u1_out11_5, u1_out11_7, u1_out14_1, u1_out14_10, u1_out14_20, 
       u1_out14_26, u1_out15_11, u1_out15_16, u1_out15_19, u1_out15_24, u1_out15_29, u1_out15_30, u1_out15_4, u1_out15_6, 
       u1_out1_13, u1_out1_18, u1_out1_2, u1_out1_28, u1_out2_13, u1_out2_18, u1_out2_2, u1_out2_28, u1_out3_12, 
       u1_out3_13, u1_out3_18, u1_out3_2, u1_out3_22, u1_out3_28, u1_out3_32, u1_out3_7, u1_out5_15, u1_out5_21, 
       u1_out5_27, u1_out5_5, u1_out6_13, u1_out6_15, u1_out6_18, u1_out6_2, u1_out6_21, u1_out6_27, u1_out6_28, 
       u1_out6_5, u1_out7_15, u1_out7_21, u1_out7_27, u1_out7_5, u1_out8_17, u1_out8_23, u1_out8_31, u1_out8_9, 
       u1_out9_1, u1_out9_10, u1_out9_11, u1_out9_12, u1_out9_13, u1_out9_16, u1_out9_18, u1_out9_19, u1_out9_2, 
       u1_out9_20, u1_out9_22, u1_out9_24, u1_out9_26, u1_out9_28, u1_out9_29, u1_out9_30, u1_out9_32, u1_out9_4, 
       u1_out9_6, u1_out9_7, u1_u0_X_27, u1_u0_X_28, u1_u0_X_29, u1_u0_X_31, u1_u0_X_33, u1_u0_X_34, u1_u0_u4_n100, 
       u1_u0_u4_n101, u1_u0_u4_n102, u1_u0_u4_n103, u1_u0_u4_n104, u1_u0_u4_n105, u1_u0_u4_n106, u1_u0_u4_n107, u1_u0_u4_n108, u1_u0_u4_n109, 
       u1_u0_u4_n110, u1_u0_u4_n111, u1_u0_u4_n112, u1_u0_u4_n113, u1_u0_u4_n114, u1_u0_u4_n115, u1_u0_u4_n116, u1_u0_u4_n117, u1_u0_u4_n118, 
       u1_u0_u4_n119, u1_u0_u4_n120, u1_u0_u4_n121, u1_u0_u4_n122, u1_u0_u4_n123, u1_u0_u4_n124, u1_u0_u4_n125, u1_u0_u4_n126, u1_u0_u4_n127, 
       u1_u0_u4_n128, u1_u0_u4_n129, u1_u0_u4_n130, u1_u0_u4_n131, u1_u0_u4_n132, u1_u0_u4_n133, u1_u0_u4_n134, u1_u0_u4_n135, u1_u0_u4_n136, 
       u1_u0_u4_n137, u1_u0_u4_n138, u1_u0_u4_n139, u1_u0_u4_n140, u1_u0_u4_n141, u1_u0_u4_n142, u1_u0_u4_n143, u1_u0_u4_n144, u1_u0_u4_n145, 
       u1_u0_u4_n146, u1_u0_u4_n147, u1_u0_u4_n148, u1_u0_u4_n149, u1_u0_u4_n150, u1_u0_u4_n151, u1_u0_u4_n152, u1_u0_u4_n153, u1_u0_u4_n154, 
       u1_u0_u4_n155, u1_u0_u4_n156, u1_u0_u4_n157, u1_u0_u4_n158, u1_u0_u4_n159, u1_u0_u4_n160, u1_u0_u4_n161, u1_u0_u4_n162, u1_u0_u4_n163, 
       u1_u0_u4_n164, u1_u0_u4_n165, u1_u0_u4_n166, u1_u0_u4_n167, u1_u0_u4_n168, u1_u0_u4_n169, u1_u0_u4_n170, u1_u0_u4_n171, u1_u0_u4_n172, 
       u1_u0_u4_n173, u1_u0_u4_n174, u1_u0_u4_n175, u1_u0_u4_n176, u1_u0_u4_n177, u1_u0_u4_n178, u1_u0_u4_n179, u1_u0_u4_n180, u1_u0_u4_n181, 
       u1_u0_u4_n182, u1_u0_u4_n183, u1_u0_u4_n184, u1_u0_u4_n185, u1_u0_u4_n186, u1_u0_u4_n94, u1_u0_u4_n95, u1_u0_u4_n96, u1_u0_u4_n97, 
       u1_u0_u4_n98, u1_u0_u4_n99, u1_u0_u5_n100, u1_u0_u5_n101, u1_u0_u5_n102, u1_u0_u5_n103, u1_u0_u5_n104, u1_u0_u5_n105, u1_u0_u5_n106, 
       u1_u0_u5_n107, u1_u0_u5_n108, u1_u0_u5_n109, u1_u0_u5_n110, u1_u0_u5_n111, u1_u0_u5_n112, u1_u0_u5_n113, u1_u0_u5_n114, u1_u0_u5_n115, 
       u1_u0_u5_n116, u1_u0_u5_n117, u1_u0_u5_n118, u1_u0_u5_n119, u1_u0_u5_n120, u1_u0_u5_n121, u1_u0_u5_n122, u1_u0_u5_n123, u1_u0_u5_n124, 
       u1_u0_u5_n125, u1_u0_u5_n126, u1_u0_u5_n127, u1_u0_u5_n128, u1_u0_u5_n129, u1_u0_u5_n130, u1_u0_u5_n131, u1_u0_u5_n132, u1_u0_u5_n133, 
       u1_u0_u5_n134, u1_u0_u5_n135, u1_u0_u5_n136, u1_u0_u5_n137, u1_u0_u5_n138, u1_u0_u5_n139, u1_u0_u5_n140, u1_u0_u5_n141, u1_u0_u5_n142, 
       u1_u0_u5_n143, u1_u0_u5_n144, u1_u0_u5_n145, u1_u0_u5_n146, u1_u0_u5_n147, u1_u0_u5_n148, u1_u0_u5_n149, u1_u0_u5_n150, u1_u0_u5_n151, 
       u1_u0_u5_n152, u1_u0_u5_n153, u1_u0_u5_n154, u1_u0_u5_n155, u1_u0_u5_n156, u1_u0_u5_n157, u1_u0_u5_n158, u1_u0_u5_n159, u1_u0_u5_n160, 
       u1_u0_u5_n161, u1_u0_u5_n162, u1_u0_u5_n163, u1_u0_u5_n164, u1_u0_u5_n165, u1_u0_u5_n166, u1_u0_u5_n167, u1_u0_u5_n168, u1_u0_u5_n169, 
       u1_u0_u5_n170, u1_u0_u5_n171, u1_u0_u5_n172, u1_u0_u5_n173, u1_u0_u5_n174, u1_u0_u5_n175, u1_u0_u5_n176, u1_u0_u5_n177, u1_u0_u5_n178, 
       u1_u0_u5_n179, u1_u0_u5_n180, u1_u0_u5_n181, u1_u0_u5_n182, u1_u0_u5_n183, u1_u0_u5_n184, u1_u0_u5_n185, u1_u0_u5_n186, u1_u0_u5_n187, 
       u1_u0_u5_n188, u1_u0_u5_n189, u1_u0_u5_n190, u1_u0_u5_n191, u1_u0_u5_n192, u1_u0_u5_n193, u1_u0_u5_n194, u1_u0_u5_n195, u1_u0_u5_n196, 
       u1_u0_u5_n99, u1_u11_X_39, u1_u11_X_40, u1_u11_X_45, u1_u11_X_46, u1_u11_u6_n100, u1_u11_u6_n101, u1_u11_u6_n102, u1_u11_u6_n103, 
       u1_u11_u6_n104, u1_u11_u6_n105, u1_u11_u6_n106, u1_u11_u6_n107, u1_u11_u6_n108, u1_u11_u6_n109, u1_u11_u6_n110, u1_u11_u6_n111, u1_u11_u6_n112, 
       u1_u11_u6_n113, u1_u11_u6_n114, u1_u11_u6_n115, u1_u11_u6_n116, u1_u11_u6_n117, u1_u11_u6_n118, u1_u11_u6_n119, u1_u11_u6_n120, u1_u11_u6_n121, 
       u1_u11_u6_n122, u1_u11_u6_n123, u1_u11_u6_n124, u1_u11_u6_n125, u1_u11_u6_n126, u1_u11_u6_n127, u1_u11_u6_n128, u1_u11_u6_n129, u1_u11_u6_n130, 
       u1_u11_u6_n131, u1_u11_u6_n132, u1_u11_u6_n133, u1_u11_u6_n134, u1_u11_u6_n135, u1_u11_u6_n136, u1_u11_u6_n137, u1_u11_u6_n138, u1_u11_u6_n139, 
       u1_u11_u6_n140, u1_u11_u6_n141, u1_u11_u6_n142, u1_u11_u6_n143, u1_u11_u6_n144, u1_u11_u6_n145, u1_u11_u6_n146, u1_u11_u6_n147, u1_u11_u6_n148, 
       u1_u11_u6_n149, u1_u11_u6_n150, u1_u11_u6_n151, u1_u11_u6_n152, u1_u11_u6_n153, u1_u11_u6_n154, u1_u11_u6_n155, u1_u11_u6_n156, u1_u11_u6_n157, 
       u1_u11_u6_n158, u1_u11_u6_n159, u1_u11_u6_n160, u1_u11_u6_n161, u1_u11_u6_n162, u1_u11_u6_n163, u1_u11_u6_n164, u1_u11_u6_n165, u1_u11_u6_n166, 
       u1_u11_u6_n167, u1_u11_u6_n168, u1_u11_u6_n169, u1_u11_u6_n170, u1_u11_u6_n171, u1_u11_u6_n172, u1_u11_u6_n173, u1_u11_u6_n174, u1_u11_u6_n88, 
       u1_u11_u6_n89, u1_u11_u6_n90, u1_u11_u6_n91, u1_u11_u6_n92, u1_u11_u6_n93, u1_u11_u6_n94, u1_u11_u6_n95, u1_u11_u6_n96, u1_u11_u6_n97, 
       u1_u11_u6_n98, u1_u11_u6_n99, u1_u11_u7_n100, u1_u11_u7_n101, u1_u11_u7_n102, u1_u11_u7_n103, u1_u11_u7_n104, u1_u11_u7_n105, u1_u11_u7_n106, 
       u1_u11_u7_n107, u1_u11_u7_n108, u1_u11_u7_n109, u1_u11_u7_n110, u1_u11_u7_n111, u1_u11_u7_n112, u1_u11_u7_n113, u1_u11_u7_n114, u1_u11_u7_n115, 
       u1_u11_u7_n116, u1_u11_u7_n117, u1_u11_u7_n118, u1_u11_u7_n119, u1_u11_u7_n120, u1_u11_u7_n121, u1_u11_u7_n122, u1_u11_u7_n123, u1_u11_u7_n124, 
       u1_u11_u7_n125, u1_u11_u7_n126, u1_u11_u7_n127, u1_u11_u7_n128, u1_u11_u7_n129, u1_u11_u7_n130, u1_u11_u7_n131, u1_u11_u7_n132, u1_u11_u7_n133, 
       u1_u11_u7_n134, u1_u11_u7_n135, u1_u11_u7_n136, u1_u11_u7_n137, u1_u11_u7_n138, u1_u11_u7_n139, u1_u11_u7_n140, u1_u11_u7_n141, u1_u11_u7_n142, 
       u1_u11_u7_n143, u1_u11_u7_n144, u1_u11_u7_n145, u1_u11_u7_n146, u1_u11_u7_n147, u1_u11_u7_n148, u1_u11_u7_n149, u1_u11_u7_n150, u1_u11_u7_n151, 
       u1_u11_u7_n152, u1_u11_u7_n153, u1_u11_u7_n154, u1_u11_u7_n155, u1_u11_u7_n156, u1_u11_u7_n157, u1_u11_u7_n158, u1_u11_u7_n159, u1_u11_u7_n160, 
       u1_u11_u7_n161, u1_u11_u7_n162, u1_u11_u7_n163, u1_u11_u7_n164, u1_u11_u7_n165, u1_u11_u7_n166, u1_u11_u7_n167, u1_u11_u7_n168, u1_u11_u7_n169, 
       u1_u11_u7_n170, u1_u11_u7_n171, u1_u11_u7_n172, u1_u11_u7_n173, u1_u11_u7_n174, u1_u11_u7_n175, u1_u11_u7_n176, u1_u11_u7_n177, u1_u11_u7_n178, 
       u1_u11_u7_n179, u1_u11_u7_n180, u1_u11_u7_n91, u1_u11_u7_n92, u1_u11_u7_n93, u1_u11_u7_n94, u1_u11_u7_n95, u1_u11_u7_n96, u1_u11_u7_n97, 
       u1_u11_u7_n98, u1_u11_u7_n99, u1_u14_X_21, u1_u14_X_22, u1_u14_u3_n100, u1_u14_u3_n101, u1_u14_u3_n102, u1_u14_u3_n103, u1_u14_u3_n104, 
       u1_u14_u3_n105, u1_u14_u3_n106, u1_u14_u3_n107, u1_u14_u3_n108, u1_u14_u3_n109, u1_u14_u3_n110, u1_u14_u3_n111, u1_u14_u3_n112, u1_u14_u3_n113, 
       u1_u14_u3_n114, u1_u14_u3_n115, u1_u14_u3_n116, u1_u14_u3_n117, u1_u14_u3_n118, u1_u14_u3_n119, u1_u14_u3_n120, u1_u14_u3_n121, u1_u14_u3_n122, 
       u1_u14_u3_n123, u1_u14_u3_n124, u1_u14_u3_n125, u1_u14_u3_n126, u1_u14_u3_n127, u1_u14_u3_n128, u1_u14_u3_n129, u1_u14_u3_n130, u1_u14_u3_n131, 
       u1_u14_u3_n132, u1_u14_u3_n133, u1_u14_u3_n134, u1_u14_u3_n135, u1_u14_u3_n136, u1_u14_u3_n137, u1_u14_u3_n138, u1_u14_u3_n139, u1_u14_u3_n140, 
       u1_u14_u3_n141, u1_u14_u3_n142, u1_u14_u3_n143, u1_u14_u3_n144, u1_u14_u3_n145, u1_u14_u3_n146, u1_u14_u3_n147, u1_u14_u3_n148, u1_u14_u3_n149, 
       u1_u14_u3_n150, u1_u14_u3_n151, u1_u14_u3_n152, u1_u14_u3_n153, u1_u14_u3_n154, u1_u14_u3_n155, u1_u14_u3_n156, u1_u14_u3_n157, u1_u14_u3_n158, 
       u1_u14_u3_n159, u1_u14_u3_n160, u1_u14_u3_n161, u1_u14_u3_n162, u1_u14_u3_n163, u1_u14_u3_n164, u1_u14_u3_n165, u1_u14_u3_n166, u1_u14_u3_n167, 
       u1_u14_u3_n168, u1_u14_u3_n169, u1_u14_u3_n170, u1_u14_u3_n171, u1_u14_u3_n172, u1_u14_u3_n173, u1_u14_u3_n174, u1_u14_u3_n175, u1_u14_u3_n176, 
       u1_u14_u3_n177, u1_u14_u3_n178, u1_u14_u3_n179, u1_u14_u3_n180, u1_u14_u3_n181, u1_u14_u3_n182, u1_u14_u3_n183, u1_u14_u3_n184, u1_u14_u3_n185, 
       u1_u14_u3_n186, u1_u14_u3_n94, u1_u14_u3_n95, u1_u14_u3_n96, u1_u14_u3_n97, u1_u14_u3_n98, u1_u14_u3_n99, u1_u15_X_15, u1_u15_X_16, 
       u1_u15_X_33, u1_u15_X_34, u1_u15_u2_n100, u1_u15_u2_n101, u1_u15_u2_n102, u1_u15_u2_n103, u1_u15_u2_n104, u1_u15_u2_n105, u1_u15_u2_n106, 
       u1_u15_u2_n107, u1_u15_u2_n108, u1_u15_u2_n109, u1_u15_u2_n110, u1_u15_u2_n111, u1_u15_u2_n112, u1_u15_u2_n113, u1_u15_u2_n114, u1_u15_u2_n115, 
       u1_u15_u2_n116, u1_u15_u2_n117, u1_u15_u2_n118, u1_u15_u2_n119, u1_u15_u2_n120, u1_u15_u2_n121, u1_u15_u2_n122, u1_u15_u2_n123, u1_u15_u2_n124, 
       u1_u15_u2_n125, u1_u15_u2_n126, u1_u15_u2_n127, u1_u15_u2_n128, u1_u15_u2_n129, u1_u15_u2_n130, u1_u15_u2_n131, u1_u15_u2_n132, u1_u15_u2_n133, 
       u1_u15_u2_n134, u1_u15_u2_n135, u1_u15_u2_n136, u1_u15_u2_n137, u1_u15_u2_n138, u1_u15_u2_n139, u1_u15_u2_n140, u1_u15_u2_n141, u1_u15_u2_n142, 
       u1_u15_u2_n143, u1_u15_u2_n144, u1_u15_u2_n145, u1_u15_u2_n146, u1_u15_u2_n147, u1_u15_u2_n148, u1_u15_u2_n149, u1_u15_u2_n150, u1_u15_u2_n151, 
       u1_u15_u2_n152, u1_u15_u2_n153, u1_u15_u2_n154, u1_u15_u2_n155, u1_u15_u2_n156, u1_u15_u2_n157, u1_u15_u2_n158, u1_u15_u2_n159, u1_u15_u2_n160, 
       u1_u15_u2_n161, u1_u15_u2_n162, u1_u15_u2_n163, u1_u15_u2_n164, u1_u15_u2_n165, u1_u15_u2_n166, u1_u15_u2_n167, u1_u15_u2_n168, u1_u15_u2_n169, 
       u1_u15_u2_n170, u1_u15_u2_n171, u1_u15_u2_n172, u1_u15_u2_n173, u1_u15_u2_n174, u1_u15_u2_n175, u1_u15_u2_n176, u1_u15_u2_n177, u1_u15_u2_n178, 
       u1_u15_u2_n179, u1_u15_u2_n180, u1_u15_u2_n181, u1_u15_u2_n182, u1_u15_u2_n183, u1_u15_u2_n184, u1_u15_u2_n185, u1_u15_u2_n186, u1_u15_u2_n187, 
       u1_u15_u2_n188, u1_u15_u2_n95, u1_u15_u2_n96, u1_u15_u2_n97, u1_u15_u2_n98, u1_u15_u2_n99, u1_u15_u5_n100, u1_u15_u5_n101, u1_u15_u5_n102, 
       u1_u15_u5_n103, u1_u15_u5_n104, u1_u15_u5_n105, u1_u15_u5_n106, u1_u15_u5_n107, u1_u15_u5_n108, u1_u15_u5_n109, u1_u15_u5_n110, u1_u15_u5_n111, 
       u1_u15_u5_n112, u1_u15_u5_n113, u1_u15_u5_n114, u1_u15_u5_n115, u1_u15_u5_n116, u1_u15_u5_n117, u1_u15_u5_n118, u1_u15_u5_n119, u1_u15_u5_n120, 
       u1_u15_u5_n121, u1_u15_u5_n122, u1_u15_u5_n123, u1_u15_u5_n124, u1_u15_u5_n125, u1_u15_u5_n126, u1_u15_u5_n127, u1_u15_u5_n128, u1_u15_u5_n129, 
       u1_u15_u5_n130, u1_u15_u5_n131, u1_u15_u5_n132, u1_u15_u5_n133, u1_u15_u5_n134, u1_u15_u5_n135, u1_u15_u5_n136, u1_u15_u5_n137, u1_u15_u5_n138, 
       u1_u15_u5_n139, u1_u15_u5_n140, u1_u15_u5_n141, u1_u15_u5_n142, u1_u15_u5_n143, u1_u15_u5_n144, u1_u15_u5_n145, u1_u15_u5_n146, u1_u15_u5_n147, 
       u1_u15_u5_n148, u1_u15_u5_n149, u1_u15_u5_n150, u1_u15_u5_n151, u1_u15_u5_n152, u1_u15_u5_n153, u1_u15_u5_n154, u1_u15_u5_n155, u1_u15_u5_n156, 
       u1_u15_u5_n157, u1_u15_u5_n158, u1_u15_u5_n159, u1_u15_u5_n160, u1_u15_u5_n161, u1_u15_u5_n162, u1_u15_u5_n163, u1_u15_u5_n164, u1_u15_u5_n165, 
       u1_u15_u5_n166, u1_u15_u5_n167, u1_u15_u5_n168, u1_u15_u5_n169, u1_u15_u5_n170, u1_u15_u5_n171, u1_u15_u5_n172, u1_u15_u5_n173, u1_u15_u5_n174, 
       u1_u15_u5_n175, u1_u15_u5_n176, u1_u15_u5_n177, u1_u15_u5_n178, u1_u15_u5_n179, u1_u15_u5_n180, u1_u15_u5_n181, u1_u15_u5_n182, u1_u15_u5_n183, 
       u1_u15_u5_n184, u1_u15_u5_n185, u1_u15_u5_n186, u1_u15_u5_n187, u1_u15_u5_n188, u1_u15_u5_n189, u1_u15_u5_n190, u1_u15_u5_n191, u1_u15_u5_n192, 
       u1_u15_u5_n193, u1_u15_u5_n194, u1_u15_u5_n195, u1_u15_u5_n196, u1_u15_u5_n99, u1_u1_X_10, u1_u1_X_9, u1_u1_u1_n100, u1_u1_u1_n101, 
       u1_u1_u1_n102, u1_u1_u1_n103, u1_u1_u1_n104, u1_u1_u1_n105, u1_u1_u1_n106, u1_u1_u1_n107, u1_u1_u1_n108, u1_u1_u1_n109, u1_u1_u1_n110, 
       u1_u1_u1_n111, u1_u1_u1_n112, u1_u1_u1_n113, u1_u1_u1_n114, u1_u1_u1_n115, u1_u1_u1_n116, u1_u1_u1_n117, u1_u1_u1_n118, u1_u1_u1_n119, 
       u1_u1_u1_n120, u1_u1_u1_n121, u1_u1_u1_n122, u1_u1_u1_n123, u1_u1_u1_n124, u1_u1_u1_n125, u1_u1_u1_n126, u1_u1_u1_n127, u1_u1_u1_n128, 
       u1_u1_u1_n129, u1_u1_u1_n130, u1_u1_u1_n131, u1_u1_u1_n132, u1_u1_u1_n133, u1_u1_u1_n134, u1_u1_u1_n135, u1_u1_u1_n136, u1_u1_u1_n137, 
       u1_u1_u1_n138, u1_u1_u1_n139, u1_u1_u1_n140, u1_u1_u1_n141, u1_u1_u1_n142, u1_u1_u1_n143, u1_u1_u1_n144, u1_u1_u1_n145, u1_u1_u1_n146, 
       u1_u1_u1_n147, u1_u1_u1_n148, u1_u1_u1_n149, u1_u1_u1_n150, u1_u1_u1_n151, u1_u1_u1_n152, u1_u1_u1_n153, u1_u1_u1_n154, u1_u1_u1_n155, 
       u1_u1_u1_n156, u1_u1_u1_n157, u1_u1_u1_n158, u1_u1_u1_n159, u1_u1_u1_n160, u1_u1_u1_n161, u1_u1_u1_n162, u1_u1_u1_n163, u1_u1_u1_n164, 
       u1_u1_u1_n165, u1_u1_u1_n166, u1_u1_u1_n167, u1_u1_u1_n168, u1_u1_u1_n169, u1_u1_u1_n170, u1_u1_u1_n171, u1_u1_u1_n172, u1_u1_u1_n173, 
       u1_u1_u1_n174, u1_u1_u1_n175, u1_u1_u1_n176, u1_u1_u1_n177, u1_u1_u1_n178, u1_u1_u1_n179, u1_u1_u1_n180, u1_u1_u1_n181, u1_u1_u1_n182, 
       u1_u1_u1_n183, u1_u1_u1_n184, u1_u1_u1_n185, u1_u1_u1_n186, u1_u1_u1_n187, u1_u1_u1_n188, u1_u1_u1_n95, u1_u1_u1_n96, u1_u1_u1_n97, 
       u1_u1_u1_n98, u1_u1_u1_n99, u1_u2_X_10, u1_u2_X_9, u1_u2_u1_n100, u1_u2_u1_n101, u1_u2_u1_n102, u1_u2_u1_n103, u1_u2_u1_n104, 
       u1_u2_u1_n105, u1_u2_u1_n106, u1_u2_u1_n107, u1_u2_u1_n108, u1_u2_u1_n109, u1_u2_u1_n110, u1_u2_u1_n111, u1_u2_u1_n112, u1_u2_u1_n113, 
       u1_u2_u1_n114, u1_u2_u1_n115, u1_u2_u1_n116, u1_u2_u1_n117, u1_u2_u1_n118, u1_u2_u1_n119, u1_u2_u1_n120, u1_u2_u1_n121, u1_u2_u1_n122, 
       u1_u2_u1_n123, u1_u2_u1_n124, u1_u2_u1_n125, u1_u2_u1_n126, u1_u2_u1_n127, u1_u2_u1_n128, u1_u2_u1_n129, u1_u2_u1_n130, u1_u2_u1_n131, 
       u1_u2_u1_n132, u1_u2_u1_n133, u1_u2_u1_n134, u1_u2_u1_n135, u1_u2_u1_n136, u1_u2_u1_n137, u1_u2_u1_n138, u1_u2_u1_n139, u1_u2_u1_n140, 
       u1_u2_u1_n141, u1_u2_u1_n142, u1_u2_u1_n143, u1_u2_u1_n144, u1_u2_u1_n145, u1_u2_u1_n146, u1_u2_u1_n147, u1_u2_u1_n148, u1_u2_u1_n149, 
       u1_u2_u1_n150, u1_u2_u1_n151, u1_u2_u1_n152, u1_u2_u1_n153, u1_u2_u1_n154, u1_u2_u1_n155, u1_u2_u1_n156, u1_u2_u1_n157, u1_u2_u1_n158, 
       u1_u2_u1_n159, u1_u2_u1_n160, u1_u2_u1_n161, u1_u2_u1_n162, u1_u2_u1_n163, u1_u2_u1_n164, u1_u2_u1_n165, u1_u2_u1_n166, u1_u2_u1_n167, 
       u1_u2_u1_n168, u1_u2_u1_n169, u1_u2_u1_n170, u1_u2_u1_n171, u1_u2_u1_n172, u1_u2_u1_n173, u1_u2_u1_n174, u1_u2_u1_n175, u1_u2_u1_n176, 
       u1_u2_u1_n177, u1_u2_u1_n178, u1_u2_u1_n179, u1_u2_u1_n180, u1_u2_u1_n181, u1_u2_u1_n182, u1_u2_u1_n183, u1_u2_u1_n184, u1_u2_u1_n185, 
       u1_u2_u1_n186, u1_u2_u1_n187, u1_u2_u1_n188, u1_u2_u1_n95, u1_u2_u1_n96, u1_u2_u1_n97, u1_u2_u1_n98, u1_u2_u1_n99, u1_u3_X_10, 
       u1_u3_X_39, u1_u3_X_40, u1_u3_X_9, u1_u3_u1_n100, u1_u3_u1_n101, u1_u3_u1_n102, u1_u3_u1_n103, u1_u3_u1_n104, u1_u3_u1_n105, 
       u1_u3_u1_n106, u1_u3_u1_n107, u1_u3_u1_n108, u1_u3_u1_n109, u1_u3_u1_n110, u1_u3_u1_n111, u1_u3_u1_n112, u1_u3_u1_n113, u1_u3_u1_n114, 
       u1_u3_u1_n115, u1_u3_u1_n116, u1_u3_u1_n117, u1_u3_u1_n118, u1_u3_u1_n119, u1_u3_u1_n120, u1_u3_u1_n121, u1_u3_u1_n122, u1_u3_u1_n123, 
       u1_u3_u1_n124, u1_u3_u1_n125, u1_u3_u1_n126, u1_u3_u1_n127, u1_u3_u1_n128, u1_u3_u1_n129, u1_u3_u1_n130, u1_u3_u1_n131, u1_u3_u1_n132, 
       u1_u3_u1_n133, u1_u3_u1_n134, u1_u3_u1_n135, u1_u3_u1_n136, u1_u3_u1_n137, u1_u3_u1_n138, u1_u3_u1_n139, u1_u3_u1_n140, u1_u3_u1_n141, 
       u1_u3_u1_n142, u1_u3_u1_n143, u1_u3_u1_n144, u1_u3_u1_n145, u1_u3_u1_n146, u1_u3_u1_n147, u1_u3_u1_n148, u1_u3_u1_n149, u1_u3_u1_n150, 
       u1_u3_u1_n151, u1_u3_u1_n152, u1_u3_u1_n153, u1_u3_u1_n154, u1_u3_u1_n155, u1_u3_u1_n156, u1_u3_u1_n157, u1_u3_u1_n158, u1_u3_u1_n159, 
       u1_u3_u1_n160, u1_u3_u1_n161, u1_u3_u1_n162, u1_u3_u1_n163, u1_u3_u1_n164, u1_u3_u1_n165, u1_u3_u1_n166, u1_u3_u1_n167, u1_u3_u1_n168, 
       u1_u3_u1_n169, u1_u3_u1_n170, u1_u3_u1_n171, u1_u3_u1_n172, u1_u3_u1_n173, u1_u3_u1_n174, u1_u3_u1_n175, u1_u3_u1_n176, u1_u3_u1_n177, 
       u1_u3_u1_n178, u1_u3_u1_n179, u1_u3_u1_n180, u1_u3_u1_n181, u1_u3_u1_n182, u1_u3_u1_n183, u1_u3_u1_n184, u1_u3_u1_n185, u1_u3_u1_n186, 
       u1_u3_u1_n187, u1_u3_u1_n188, u1_u3_u1_n95, u1_u3_u1_n96, u1_u3_u1_n97, u1_u3_u1_n98, u1_u3_u1_n99, u1_u3_u6_n100, u1_u3_u6_n101, 
       u1_u3_u6_n102, u1_u3_u6_n103, u1_u3_u6_n104, u1_u3_u6_n105, u1_u3_u6_n106, u1_u3_u6_n107, u1_u3_u6_n108, u1_u3_u6_n109, u1_u3_u6_n110, 
       u1_u3_u6_n111, u1_u3_u6_n112, u1_u3_u6_n113, u1_u3_u6_n114, u1_u3_u6_n115, u1_u3_u6_n116, u1_u3_u6_n117, u1_u3_u6_n118, u1_u3_u6_n119, 
       u1_u3_u6_n120, u1_u3_u6_n121, u1_u3_u6_n122, u1_u3_u6_n123, u1_u3_u6_n124, u1_u3_u6_n125, u1_u3_u6_n126, u1_u3_u6_n127, u1_u3_u6_n128, 
       u1_u3_u6_n129, u1_u3_u6_n130, u1_u3_u6_n131, u1_u3_u6_n132, u1_u3_u6_n133, u1_u3_u6_n134, u1_u3_u6_n135, u1_u3_u6_n136, u1_u3_u6_n137, 
       u1_u3_u6_n138, u1_u3_u6_n139, u1_u3_u6_n140, u1_u3_u6_n141, u1_u3_u6_n142, u1_u3_u6_n143, u1_u3_u6_n144, u1_u3_u6_n145, u1_u3_u6_n146, 
       u1_u3_u6_n147, u1_u3_u6_n148, u1_u3_u6_n149, u1_u3_u6_n150, u1_u3_u6_n151, u1_u3_u6_n152, u1_u3_u6_n153, u1_u3_u6_n154, u1_u3_u6_n155, 
       u1_u3_u6_n156, u1_u3_u6_n157, u1_u3_u6_n158, u1_u3_u6_n159, u1_u3_u6_n160, u1_u3_u6_n161, u1_u3_u6_n162, u1_u3_u6_n163, u1_u3_u6_n164, 
       u1_u3_u6_n165, u1_u3_u6_n166, u1_u3_u6_n167, u1_u3_u6_n168, u1_u3_u6_n169, u1_u3_u6_n170, u1_u3_u6_n171, u1_u3_u6_n172, u1_u3_u6_n173, 
       u1_u3_u6_n174, u1_u3_u6_n88, u1_u3_u6_n89, u1_u3_u6_n90, u1_u3_u6_n91, u1_u3_u6_n92, u1_u3_u6_n93, u1_u3_u6_n94, u1_u3_u6_n95, 
       u1_u3_u6_n96, u1_u3_u6_n97, u1_u3_u6_n98, u1_u3_u6_n99, u1_u5_X_45, u1_u5_X_46, u1_u5_u7_n100, u1_u5_u7_n101, u1_u5_u7_n102, 
       u1_u5_u7_n103, u1_u5_u7_n104, u1_u5_u7_n105, u1_u5_u7_n106, u1_u5_u7_n107, u1_u5_u7_n108, u1_u5_u7_n109, u1_u5_u7_n110, u1_u5_u7_n111, 
       u1_u5_u7_n112, u1_u5_u7_n113, u1_u5_u7_n114, u1_u5_u7_n115, u1_u5_u7_n116, u1_u5_u7_n117, u1_u5_u7_n118, u1_u5_u7_n119, u1_u5_u7_n120, 
       u1_u5_u7_n121, u1_u5_u7_n122, u1_u5_u7_n123, u1_u5_u7_n124, u1_u5_u7_n125, u1_u5_u7_n126, u1_u5_u7_n127, u1_u5_u7_n128, u1_u5_u7_n129, 
       u1_u5_u7_n130, u1_u5_u7_n131, u1_u5_u7_n132, u1_u5_u7_n133, u1_u5_u7_n134, u1_u5_u7_n135, u1_u5_u7_n136, u1_u5_u7_n137, u1_u5_u7_n138, 
       u1_u5_u7_n139, u1_u5_u7_n140, u1_u5_u7_n141, u1_u5_u7_n142, u1_u5_u7_n143, u1_u5_u7_n144, u1_u5_u7_n145, u1_u5_u7_n146, u1_u5_u7_n147, 
       u1_u5_u7_n148, u1_u5_u7_n149, u1_u5_u7_n150, u1_u5_u7_n151, u1_u5_u7_n152, u1_u5_u7_n153, u1_u5_u7_n154, u1_u5_u7_n155, u1_u5_u7_n156, 
       u1_u5_u7_n157, u1_u5_u7_n158, u1_u5_u7_n159, u1_u5_u7_n160, u1_u5_u7_n161, u1_u5_u7_n162, u1_u5_u7_n163, u1_u5_u7_n164, u1_u5_u7_n165, 
       u1_u5_u7_n166, u1_u5_u7_n167, u1_u5_u7_n168, u1_u5_u7_n169, u1_u5_u7_n170, u1_u5_u7_n171, u1_u5_u7_n172, u1_u5_u7_n173, u1_u5_u7_n174, 
       u1_u5_u7_n175, u1_u5_u7_n176, u1_u5_u7_n177, u1_u5_u7_n178, u1_u5_u7_n179, u1_u5_u7_n180, u1_u5_u7_n91, u1_u5_u7_n92, u1_u5_u7_n93, 
       u1_u5_u7_n94, u1_u5_u7_n95, u1_u5_u7_n96, u1_u5_u7_n97, u1_u5_u7_n98, u1_u5_u7_n99, u1_u6_X_10, u1_u6_X_45, u1_u6_X_46, 
       u1_u6_X_9, u1_u6_u1_n100, u1_u6_u1_n101, u1_u6_u1_n102, u1_u6_u1_n103, u1_u6_u1_n104, u1_u6_u1_n105, u1_u6_u1_n106, u1_u6_u1_n107, 
       u1_u6_u1_n108, u1_u6_u1_n109, u1_u6_u1_n110, u1_u6_u1_n111, u1_u6_u1_n112, u1_u6_u1_n113, u1_u6_u1_n114, u1_u6_u1_n115, u1_u6_u1_n116, 
       u1_u6_u1_n117, u1_u6_u1_n118, u1_u6_u1_n119, u1_u6_u1_n120, u1_u6_u1_n121, u1_u6_u1_n122, u1_u6_u1_n123, u1_u6_u1_n124, u1_u6_u1_n125, 
       u1_u6_u1_n126, u1_u6_u1_n127, u1_u6_u1_n128, u1_u6_u1_n129, u1_u6_u1_n130, u1_u6_u1_n131, u1_u6_u1_n132, u1_u6_u1_n133, u1_u6_u1_n134, 
       u1_u6_u1_n135, u1_u6_u1_n136, u1_u6_u1_n137, u1_u6_u1_n138, u1_u6_u1_n139, u1_u6_u1_n140, u1_u6_u1_n141, u1_u6_u1_n142, u1_u6_u1_n143, 
       u1_u6_u1_n144, u1_u6_u1_n145, u1_u6_u1_n146, u1_u6_u1_n147, u1_u6_u1_n148, u1_u6_u1_n149, u1_u6_u1_n150, u1_u6_u1_n151, u1_u6_u1_n152, 
       u1_u6_u1_n153, u1_u6_u1_n154, u1_u6_u1_n155, u1_u6_u1_n156, u1_u6_u1_n157, u1_u6_u1_n158, u1_u6_u1_n159, u1_u6_u1_n160, u1_u6_u1_n161, 
       u1_u6_u1_n162, u1_u6_u1_n163, u1_u6_u1_n164, u1_u6_u1_n165, u1_u6_u1_n166, u1_u6_u1_n167, u1_u6_u1_n168, u1_u6_u1_n169, u1_u6_u1_n170, 
       u1_u6_u1_n171, u1_u6_u1_n172, u1_u6_u1_n173, u1_u6_u1_n174, u1_u6_u1_n175, u1_u6_u1_n176, u1_u6_u1_n177, u1_u6_u1_n178, u1_u6_u1_n179, 
       u1_u6_u1_n180, u1_u6_u1_n181, u1_u6_u1_n182, u1_u6_u1_n183, u1_u6_u1_n184, u1_u6_u1_n185, u1_u6_u1_n186, u1_u6_u1_n187, u1_u6_u1_n188, 
       u1_u6_u1_n95, u1_u6_u1_n96, u1_u6_u1_n97, u1_u6_u1_n98, u1_u6_u1_n99, u1_u6_u7_n100, u1_u6_u7_n101, u1_u6_u7_n102, u1_u6_u7_n103, 
       u1_u6_u7_n104, u1_u6_u7_n105, u1_u6_u7_n106, u1_u6_u7_n107, u1_u6_u7_n108, u1_u6_u7_n109, u1_u6_u7_n110, u1_u6_u7_n111, u1_u6_u7_n112, 
       u1_u6_u7_n113, u1_u6_u7_n114, u1_u6_u7_n115, u1_u6_u7_n116, u1_u6_u7_n117, u1_u6_u7_n118, u1_u6_u7_n119, u1_u6_u7_n120, u1_u6_u7_n121, 
       u1_u6_u7_n122, u1_u6_u7_n123, u1_u6_u7_n124, u1_u6_u7_n125, u1_u6_u7_n126, u1_u6_u7_n127, u1_u6_u7_n128, u1_u6_u7_n129, u1_u6_u7_n130, 
       u1_u6_u7_n131, u1_u6_u7_n132, u1_u6_u7_n133, u1_u6_u7_n134, u1_u6_u7_n135, u1_u6_u7_n136, u1_u6_u7_n137, u1_u6_u7_n138, u1_u6_u7_n139, 
       u1_u6_u7_n140, u1_u6_u7_n141, u1_u6_u7_n142, u1_u6_u7_n143, u1_u6_u7_n144, u1_u6_u7_n145, u1_u6_u7_n146, u1_u6_u7_n147, u1_u6_u7_n148, 
       u1_u6_u7_n149, u1_u6_u7_n150, u1_u6_u7_n151, u1_u6_u7_n152, u1_u6_u7_n153, u1_u6_u7_n154, u1_u6_u7_n155, u1_u6_u7_n156, u1_u6_u7_n157, 
       u1_u6_u7_n158, u1_u6_u7_n159, u1_u6_u7_n160, u1_u6_u7_n161, u1_u6_u7_n162, u1_u6_u7_n163, u1_u6_u7_n164, u1_u6_u7_n165, u1_u6_u7_n166, 
       u1_u6_u7_n167, u1_u6_u7_n168, u1_u6_u7_n169, u1_u6_u7_n170, u1_u6_u7_n171, u1_u6_u7_n172, u1_u6_u7_n173, u1_u6_u7_n174, u1_u6_u7_n175, 
       u1_u6_u7_n176, u1_u6_u7_n177, u1_u6_u7_n178, u1_u6_u7_n179, u1_u6_u7_n180, u1_u6_u7_n91, u1_u6_u7_n92, u1_u6_u7_n93, u1_u6_u7_n94, 
       u1_u6_u7_n95, u1_u6_u7_n96, u1_u6_u7_n97, u1_u6_u7_n98, u1_u6_u7_n99, u1_u7_X_45, u1_u7_X_46, u1_u7_u7_n100, u1_u7_u7_n101, 
       u1_u7_u7_n102, u1_u7_u7_n103, u1_u7_u7_n104, u1_u7_u7_n105, u1_u7_u7_n106, u1_u7_u7_n107, u1_u7_u7_n108, u1_u7_u7_n109, u1_u7_u7_n110, 
       u1_u7_u7_n111, u1_u7_u7_n112, u1_u7_u7_n113, u1_u7_u7_n114, u1_u7_u7_n115, u1_u7_u7_n116, u1_u7_u7_n117, u1_u7_u7_n118, u1_u7_u7_n119, 
       u1_u7_u7_n120, u1_u7_u7_n121, u1_u7_u7_n122, u1_u7_u7_n123, u1_u7_u7_n124, u1_u7_u7_n125, u1_u7_u7_n126, u1_u7_u7_n127, u1_u7_u7_n128, 
       u1_u7_u7_n129, u1_u7_u7_n130, u1_u7_u7_n131, u1_u7_u7_n132, u1_u7_u7_n133, u1_u7_u7_n134, u1_u7_u7_n135, u1_u7_u7_n136, u1_u7_u7_n137, 
       u1_u7_u7_n138, u1_u7_u7_n139, u1_u7_u7_n140, u1_u7_u7_n141, u1_u7_u7_n142, u1_u7_u7_n143, u1_u7_u7_n144, u1_u7_u7_n145, u1_u7_u7_n146, 
       u1_u7_u7_n147, u1_u7_u7_n148, u1_u7_u7_n149, u1_u7_u7_n150, u1_u7_u7_n151, u1_u7_u7_n152, u1_u7_u7_n153, u1_u7_u7_n154, u1_u7_u7_n155, 
       u1_u7_u7_n156, u1_u7_u7_n157, u1_u7_u7_n158, u1_u7_u7_n159, u1_u7_u7_n160, u1_u7_u7_n161, u1_u7_u7_n162, u1_u7_u7_n163, u1_u7_u7_n164, 
       u1_u7_u7_n165, u1_u7_u7_n166, u1_u7_u7_n167, u1_u7_u7_n168, u1_u7_u7_n169, u1_u7_u7_n170, u1_u7_u7_n171, u1_u7_u7_n172, u1_u7_u7_n173, 
       u1_u7_u7_n174, u1_u7_u7_n175, u1_u7_u7_n176, u1_u7_u7_n177, u1_u7_u7_n178, u1_u7_u7_n179, u1_u7_u7_n180, u1_u7_u7_n91, u1_u7_u7_n92, 
       u1_u7_u7_n93, u1_u7_u7_n94, u1_u7_u7_n95, u1_u7_u7_n96, u1_u7_u7_n97, u1_u7_u7_n98, u1_u7_u7_n99, u1_u8_X_3, u1_u8_X_4, 
       u1_u8_u0_n100, u1_u8_u0_n101, u1_u8_u0_n102, u1_u8_u0_n103, u1_u8_u0_n104, u1_u8_u0_n105, u1_u8_u0_n106, u1_u8_u0_n107, u1_u8_u0_n108, 
       u1_u8_u0_n109, u1_u8_u0_n110, u1_u8_u0_n111, u1_u8_u0_n112, u1_u8_u0_n113, u1_u8_u0_n114, u1_u8_u0_n115, u1_u8_u0_n116, u1_u8_u0_n117, 
       u1_u8_u0_n118, u1_u8_u0_n119, u1_u8_u0_n120, u1_u8_u0_n121, u1_u8_u0_n122, u1_u8_u0_n123, u1_u8_u0_n124, u1_u8_u0_n125, u1_u8_u0_n126, 
       u1_u8_u0_n127, u1_u8_u0_n128, u1_u8_u0_n129, u1_u8_u0_n130, u1_u8_u0_n131, u1_u8_u0_n132, u1_u8_u0_n133, u1_u8_u0_n134, u1_u8_u0_n135, 
       u1_u8_u0_n136, u1_u8_u0_n137, u1_u8_u0_n138, u1_u8_u0_n139, u1_u8_u0_n140, u1_u8_u0_n141, u1_u8_u0_n142, u1_u8_u0_n143, u1_u8_u0_n144, 
       u1_u8_u0_n145, u1_u8_u0_n146, u1_u8_u0_n147, u1_u8_u0_n148, u1_u8_u0_n149, u1_u8_u0_n150, u1_u8_u0_n151, u1_u8_u0_n152, u1_u8_u0_n153, 
       u1_u8_u0_n154, u1_u8_u0_n155, u1_u8_u0_n156, u1_u8_u0_n157, u1_u8_u0_n158, u1_u8_u0_n159, u1_u8_u0_n160, u1_u8_u0_n161, u1_u8_u0_n162, 
       u1_u8_u0_n163, u1_u8_u0_n164, u1_u8_u0_n165, u1_u8_u0_n166, u1_u8_u0_n167, u1_u8_u0_n168, u1_u8_u0_n169, u1_u8_u0_n170, u1_u8_u0_n171, 
       u1_u8_u0_n172, u1_u8_u0_n173, u1_u8_u0_n174, u1_u8_u0_n88, u1_u8_u0_n89, u1_u8_u0_n90, u1_u8_u0_n91, u1_u8_u0_n92, u1_u8_u0_n93, 
       u1_u8_u0_n94, u1_u8_u0_n95, u1_u8_u0_n96, u1_u8_u0_n97, u1_u8_u0_n98, u1_u8_u0_n99, u1_u9_X_10, u1_u9_X_11, u1_u9_X_12, 
       u1_u9_X_13, u1_u9_X_14, u1_u9_X_15, u1_u9_X_16, u1_u9_X_17, u1_u9_X_18, u1_u9_X_19, u1_u9_X_20, u1_u9_X_21, 
       u1_u9_X_22, u1_u9_X_33, u1_u9_X_34, u1_u9_X_35, u1_u9_X_36, u1_u9_X_37, u1_u9_X_38, u1_u9_X_39, u1_u9_X_40, 
       u1_u9_X_9, u1_u9_u1_n100, u1_u9_u1_n101, u1_u9_u1_n102, u1_u9_u1_n103, u1_u9_u1_n104, u1_u9_u1_n105, u1_u9_u1_n106, u1_u9_u1_n107, 
       u1_u9_u1_n108, u1_u9_u1_n109, u1_u9_u1_n110, u1_u9_u1_n111, u1_u9_u1_n112, u1_u9_u1_n113, u1_u9_u1_n114, u1_u9_u1_n115, u1_u9_u1_n116, 
       u1_u9_u1_n117, u1_u9_u1_n118, u1_u9_u1_n119, u1_u9_u1_n120, u1_u9_u1_n121, u1_u9_u1_n122, u1_u9_u1_n123, u1_u9_u1_n124, u1_u9_u1_n125, 
       u1_u9_u1_n126, u1_u9_u1_n127, u1_u9_u1_n128, u1_u9_u1_n129, u1_u9_u1_n130, u1_u9_u1_n131, u1_u9_u1_n132, u1_u9_u1_n133, u1_u9_u1_n134, 
       u1_u9_u1_n135, u1_u9_u1_n136, u1_u9_u1_n137, u1_u9_u1_n138, u1_u9_u1_n139, u1_u9_u1_n140, u1_u9_u1_n141, u1_u9_u1_n142, u1_u9_u1_n143, 
       u1_u9_u1_n144, u1_u9_u1_n145, u1_u9_u1_n146, u1_u9_u1_n147, u1_u9_u1_n148, u1_u9_u1_n149, u1_u9_u1_n150, u1_u9_u1_n151, u1_u9_u1_n152, 
       u1_u9_u1_n153, u1_u9_u1_n154, u1_u9_u1_n155, u1_u9_u1_n156, u1_u9_u1_n157, u1_u9_u1_n158, u1_u9_u1_n159, u1_u9_u1_n160, u1_u9_u1_n161, 
       u1_u9_u1_n162, u1_u9_u1_n163, u1_u9_u1_n164, u1_u9_u1_n165, u1_u9_u1_n166, u1_u9_u1_n167, u1_u9_u1_n168, u1_u9_u1_n169, u1_u9_u1_n170, 
       u1_u9_u1_n171, u1_u9_u1_n172, u1_u9_u1_n173, u1_u9_u1_n174, u1_u9_u1_n175, u1_u9_u1_n176, u1_u9_u1_n177, u1_u9_u1_n178, u1_u9_u1_n179, 
       u1_u9_u1_n180, u1_u9_u1_n181, u1_u9_u1_n182, u1_u9_u1_n183, u1_u9_u1_n184, u1_u9_u1_n185, u1_u9_u1_n186, u1_u9_u1_n187, u1_u9_u1_n188, 
       u1_u9_u1_n95, u1_u9_u1_n96, u1_u9_u1_n97, u1_u9_u1_n98, u1_u9_u1_n99, u1_u9_u2_n100, u1_u9_u2_n101, u1_u9_u2_n102, u1_u9_u2_n103, 
       u1_u9_u2_n104, u1_u9_u2_n105, u1_u9_u2_n106, u1_u9_u2_n107, u1_u9_u2_n108, u1_u9_u2_n109, u1_u9_u2_n110, u1_u9_u2_n111, u1_u9_u2_n112, 
       u1_u9_u2_n113, u1_u9_u2_n114, u1_u9_u2_n115, u1_u9_u2_n116, u1_u9_u2_n117, u1_u9_u2_n118, u1_u9_u2_n119, u1_u9_u2_n120, u1_u9_u2_n121, 
       u1_u9_u2_n122, u1_u9_u2_n123, u1_u9_u2_n124, u1_u9_u2_n125, u1_u9_u2_n126, u1_u9_u2_n127, u1_u9_u2_n128, u1_u9_u2_n129, u1_u9_u2_n130, 
       u1_u9_u2_n131, u1_u9_u2_n132, u1_u9_u2_n133, u1_u9_u2_n134, u1_u9_u2_n135, u1_u9_u2_n136, u1_u9_u2_n137, u1_u9_u2_n138, u1_u9_u2_n139, 
       u1_u9_u2_n140, u1_u9_u2_n141, u1_u9_u2_n142, u1_u9_u2_n143, u1_u9_u2_n144, u1_u9_u2_n145, u1_u9_u2_n146, u1_u9_u2_n147, u1_u9_u2_n148, 
       u1_u9_u2_n149, u1_u9_u2_n150, u1_u9_u2_n151, u1_u9_u2_n152, u1_u9_u2_n153, u1_u9_u2_n154, u1_u9_u2_n155, u1_u9_u2_n156, u1_u9_u2_n157, 
       u1_u9_u2_n158, u1_u9_u2_n159, u1_u9_u2_n160, u1_u9_u2_n161, u1_u9_u2_n162, u1_u9_u2_n163, u1_u9_u2_n164, u1_u9_u2_n165, u1_u9_u2_n166, 
       u1_u9_u2_n167, u1_u9_u2_n168, u1_u9_u2_n169, u1_u9_u2_n170, u1_u9_u2_n171, u1_u9_u2_n172, u1_u9_u2_n173, u1_u9_u2_n174, u1_u9_u2_n175, 
       u1_u9_u2_n176, u1_u9_u2_n177, u1_u9_u2_n178, u1_u9_u2_n179, u1_u9_u2_n180, u1_u9_u2_n181, u1_u9_u2_n182, u1_u9_u2_n183, u1_u9_u2_n184, 
       u1_u9_u2_n185, u1_u9_u2_n186, u1_u9_u2_n187, u1_u9_u2_n188, u1_u9_u2_n95, u1_u9_u2_n96, u1_u9_u2_n97, u1_u9_u2_n98, u1_u9_u2_n99, 
       u1_u9_u3_n100, u1_u9_u3_n101, u1_u9_u3_n102, u1_u9_u3_n103, u1_u9_u3_n104, u1_u9_u3_n105, u1_u9_u3_n106, u1_u9_u3_n107, u1_u9_u3_n108, 
       u1_u9_u3_n109, u1_u9_u3_n110, u1_u9_u3_n111, u1_u9_u3_n112, u1_u9_u3_n113, u1_u9_u3_n114, u1_u9_u3_n115, u1_u9_u3_n116, u1_u9_u3_n117, 
       u1_u9_u3_n118, u1_u9_u3_n119, u1_u9_u3_n120, u1_u9_u3_n121, u1_u9_u3_n122, u1_u9_u3_n123, u1_u9_u3_n124, u1_u9_u3_n125, u1_u9_u3_n126, 
       u1_u9_u3_n127, u1_u9_u3_n128, u1_u9_u3_n129, u1_u9_u3_n130, u1_u9_u3_n131, u1_u9_u3_n132, u1_u9_u3_n133, u1_u9_u3_n134, u1_u9_u3_n135, 
       u1_u9_u3_n136, u1_u9_u3_n137, u1_u9_u3_n138, u1_u9_u3_n139, u1_u9_u3_n140, u1_u9_u3_n141, u1_u9_u3_n142, u1_u9_u3_n143, u1_u9_u3_n144, 
       u1_u9_u3_n145, u1_u9_u3_n146, u1_u9_u3_n147, u1_u9_u3_n148, u1_u9_u3_n149, u1_u9_u3_n150, u1_u9_u3_n151, u1_u9_u3_n152, u1_u9_u3_n153, 
       u1_u9_u3_n154, u1_u9_u3_n155, u1_u9_u3_n156, u1_u9_u3_n157, u1_u9_u3_n158, u1_u9_u3_n159, u1_u9_u3_n160, u1_u9_u3_n161, u1_u9_u3_n162, 
       u1_u9_u3_n163, u1_u9_u3_n164, u1_u9_u3_n165, u1_u9_u3_n166, u1_u9_u3_n167, u1_u9_u3_n168, u1_u9_u3_n169, u1_u9_u3_n170, u1_u9_u3_n171, 
       u1_u9_u3_n172, u1_u9_u3_n173, u1_u9_u3_n174, u1_u9_u3_n175, u1_u9_u3_n176, u1_u9_u3_n177, u1_u9_u3_n178, u1_u9_u3_n179, u1_u9_u3_n180, 
       u1_u9_u3_n181, u1_u9_u3_n182, u1_u9_u3_n183, u1_u9_u3_n184, u1_u9_u3_n185, u1_u9_u3_n186, u1_u9_u3_n94, u1_u9_u3_n95, u1_u9_u3_n96, 
       u1_u9_u3_n97, u1_u9_u3_n98, u1_u9_u3_n99, u1_u9_u5_n100, u1_u9_u5_n101, u1_u9_u5_n102, u1_u9_u5_n103, u1_u9_u5_n104, u1_u9_u5_n105, 
       u1_u9_u5_n106, u1_u9_u5_n107, u1_u9_u5_n108, u1_u9_u5_n109, u1_u9_u5_n110, u1_u9_u5_n111, u1_u9_u5_n112, u1_u9_u5_n113, u1_u9_u5_n114, 
       u1_u9_u5_n115, u1_u9_u5_n116, u1_u9_u5_n117, u1_u9_u5_n118, u1_u9_u5_n119, u1_u9_u5_n120, u1_u9_u5_n121, u1_u9_u5_n122, u1_u9_u5_n123, 
       u1_u9_u5_n124, u1_u9_u5_n125, u1_u9_u5_n126, u1_u9_u5_n127, u1_u9_u5_n128, u1_u9_u5_n129, u1_u9_u5_n130, u1_u9_u5_n131, u1_u9_u5_n132, 
       u1_u9_u5_n133, u1_u9_u5_n134, u1_u9_u5_n135, u1_u9_u5_n136, u1_u9_u5_n137, u1_u9_u5_n138, u1_u9_u5_n139, u1_u9_u5_n140, u1_u9_u5_n141, 
       u1_u9_u5_n142, u1_u9_u5_n143, u1_u9_u5_n144, u1_u9_u5_n145, u1_u9_u5_n146, u1_u9_u5_n147, u1_u9_u5_n148, u1_u9_u5_n149, u1_u9_u5_n150, 
       u1_u9_u5_n151, u1_u9_u5_n152, u1_u9_u5_n153, u1_u9_u5_n154, u1_u9_u5_n155, u1_u9_u5_n156, u1_u9_u5_n157, u1_u9_u5_n158, u1_u9_u5_n159, 
       u1_u9_u5_n160, u1_u9_u5_n161, u1_u9_u5_n162, u1_u9_u5_n163, u1_u9_u5_n164, u1_u9_u5_n165, u1_u9_u5_n166, u1_u9_u5_n167, u1_u9_u5_n168, 
       u1_u9_u5_n169, u1_u9_u5_n170, u1_u9_u5_n171, u1_u9_u5_n172, u1_u9_u5_n173, u1_u9_u5_n174, u1_u9_u5_n175, u1_u9_u5_n176, u1_u9_u5_n177, 
       u1_u9_u5_n178, u1_u9_u5_n179, u1_u9_u5_n180, u1_u9_u5_n181, u1_u9_u5_n182, u1_u9_u5_n183, u1_u9_u5_n184, u1_u9_u5_n185, u1_u9_u5_n186, 
       u1_u9_u5_n187, u1_u9_u5_n188, u1_u9_u5_n189, u1_u9_u5_n190, u1_u9_u5_n191, u1_u9_u5_n192, u1_u9_u5_n193, u1_u9_u5_n194, u1_u9_u5_n195, 
       u1_u9_u5_n196, u1_u9_u5_n99, u1_u9_u6_n100, u1_u9_u6_n101, u1_u9_u6_n102, u1_u9_u6_n103, u1_u9_u6_n104, u1_u9_u6_n105, u1_u9_u6_n106, 
       u1_u9_u6_n107, u1_u9_u6_n108, u1_u9_u6_n109, u1_u9_u6_n110, u1_u9_u6_n111, u1_u9_u6_n112, u1_u9_u6_n113, u1_u9_u6_n114, u1_u9_u6_n115, 
       u1_u9_u6_n116, u1_u9_u6_n117, u1_u9_u6_n118, u1_u9_u6_n119, u1_u9_u6_n120, u1_u9_u6_n121, u1_u9_u6_n122, u1_u9_u6_n123, u1_u9_u6_n124, 
       u1_u9_u6_n125, u1_u9_u6_n126, u1_u9_u6_n127, u1_u9_u6_n128, u1_u9_u6_n129, u1_u9_u6_n130, u1_u9_u6_n131, u1_u9_u6_n132, u1_u9_u6_n133, 
       u1_u9_u6_n134, u1_u9_u6_n135, u1_u9_u6_n136, u1_u9_u6_n137, u1_u9_u6_n138, u1_u9_u6_n139, u1_u9_u6_n140, u1_u9_u6_n141, u1_u9_u6_n142, 
       u1_u9_u6_n143, u1_u9_u6_n144, u1_u9_u6_n145, u1_u9_u6_n146, u1_u9_u6_n147, u1_u9_u6_n148, u1_u9_u6_n149, u1_u9_u6_n150, u1_u9_u6_n151, 
       u1_u9_u6_n152, u1_u9_u6_n153, u1_u9_u6_n154, u1_u9_u6_n155, u1_u9_u6_n156, u1_u9_u6_n157, u1_u9_u6_n158, u1_u9_u6_n159, u1_u9_u6_n160, 
       u1_u9_u6_n161, u1_u9_u6_n162, u1_u9_u6_n163, u1_u9_u6_n164, u1_u9_u6_n165, u1_u9_u6_n166, u1_u9_u6_n167, u1_u9_u6_n168, u1_u9_u6_n169, 
       u1_u9_u6_n170, u1_u9_u6_n171, u1_u9_u6_n172, u1_u9_u6_n173, u1_u9_u6_n174, u1_u9_u6_n88, u1_u9_u6_n89, u1_u9_u6_n90, u1_u9_u6_n91, 
       u1_u9_u6_n92, u1_u9_u6_n93, u1_u9_u6_n94, u1_u9_u6_n95, u1_u9_u6_n96, u1_u9_u6_n97, u1_u9_u6_n98, u1_u9_u6_n99, u2_K2_2, 
       u2_K2_3, u2_K2_4, u2_K2_5, u2_K2_6, u2_out1_15, u2_out1_17, u2_out1_21, u2_out1_23, u2_out1_27, 
       u2_out1_31, u2_out1_5, u2_out1_9, u2_u1_X_1, u2_u1_X_2, u2_u1_X_3, u2_u1_X_4, u2_u1_X_43, u2_u1_X_44, 
       u2_u1_X_45, u2_u1_X_46, u2_u1_X_47, u2_u1_X_48, u2_u1_X_5, u2_u1_X_6, u2_u1_u0_n100, u2_u1_u0_n101, u2_u1_u0_n102, 
       u2_u1_u0_n103, u2_u1_u0_n104, u2_u1_u0_n105, u2_u1_u0_n106, u2_u1_u0_n107, u2_u1_u0_n108, u2_u1_u0_n109, u2_u1_u0_n110, u2_u1_u0_n111, 
       u2_u1_u0_n112, u2_u1_u0_n113, u2_u1_u0_n114, u2_u1_u0_n115, u2_u1_u0_n116, u2_u1_u0_n117, u2_u1_u0_n118, u2_u1_u0_n119, u2_u1_u0_n120, 
       u2_u1_u0_n121, u2_u1_u0_n122, u2_u1_u0_n123, u2_u1_u0_n124, u2_u1_u0_n125, u2_u1_u0_n126, u2_u1_u0_n127, u2_u1_u0_n128, u2_u1_u0_n129, 
       u2_u1_u0_n130, u2_u1_u0_n131, u2_u1_u0_n132, u2_u1_u0_n133, u2_u1_u0_n134, u2_u1_u0_n135, u2_u1_u0_n136, u2_u1_u0_n137, u2_u1_u0_n138, 
       u2_u1_u0_n139, u2_u1_u0_n140, u2_u1_u0_n141, u2_u1_u0_n142, u2_u1_u0_n143, u2_u1_u0_n144, u2_u1_u0_n145, u2_u1_u0_n146, u2_u1_u0_n147, 
       u2_u1_u0_n148, u2_u1_u0_n149, u2_u1_u0_n150, u2_u1_u0_n151, u2_u1_u0_n152, u2_u1_u0_n153, u2_u1_u0_n154, u2_u1_u0_n155, u2_u1_u0_n156, 
       u2_u1_u0_n157, u2_u1_u0_n158, u2_u1_u0_n159, u2_u1_u0_n160, u2_u1_u0_n161, u2_u1_u0_n162, u2_u1_u0_n163, u2_u1_u0_n164, u2_u1_u0_n165, 
       u2_u1_u0_n166, u2_u1_u0_n167, u2_u1_u0_n168, u2_u1_u0_n169, u2_u1_u0_n170, u2_u1_u0_n171, u2_u1_u0_n172, u2_u1_u0_n173, u2_u1_u0_n174, 
       u2_u1_u0_n88, u2_u1_u0_n89, u2_u1_u0_n90, u2_u1_u0_n91, u2_u1_u0_n92, u2_u1_u0_n93, u2_u1_u0_n94, u2_u1_u0_n95, u2_u1_u0_n96, 
       u2_u1_u0_n97, u2_u1_u0_n98, u2_u1_u0_n99, u2_u1_u7_n100, u2_u1_u7_n101, u2_u1_u7_n102, u2_u1_u7_n103, u2_u1_u7_n104, u2_u1_u7_n105, 
       u2_u1_u7_n106, u2_u1_u7_n107, u2_u1_u7_n108, u2_u1_u7_n109, u2_u1_u7_n110, u2_u1_u7_n111, u2_u1_u7_n112, u2_u1_u7_n113, u2_u1_u7_n114, 
       u2_u1_u7_n115, u2_u1_u7_n116, u2_u1_u7_n117, u2_u1_u7_n118, u2_u1_u7_n119, u2_u1_u7_n120, u2_u1_u7_n121, u2_u1_u7_n122, u2_u1_u7_n123, 
       u2_u1_u7_n124, u2_u1_u7_n125, u2_u1_u7_n126, u2_u1_u7_n127, u2_u1_u7_n128, u2_u1_u7_n129, u2_u1_u7_n130, u2_u1_u7_n131, u2_u1_u7_n132, 
       u2_u1_u7_n133, u2_u1_u7_n134, u2_u1_u7_n135, u2_u1_u7_n136, u2_u1_u7_n137, u2_u1_u7_n138, u2_u1_u7_n139, u2_u1_u7_n140, u2_u1_u7_n141, 
       u2_u1_u7_n142, u2_u1_u7_n143, u2_u1_u7_n144, u2_u1_u7_n145, u2_u1_u7_n146, u2_u1_u7_n147, u2_u1_u7_n148, u2_u1_u7_n149, u2_u1_u7_n150, 
       u2_u1_u7_n151, u2_u1_u7_n152, u2_u1_u7_n153, u2_u1_u7_n154, u2_u1_u7_n155, u2_u1_u7_n156, u2_u1_u7_n157, u2_u1_u7_n158, u2_u1_u7_n159, 
       u2_u1_u7_n160, u2_u1_u7_n161, u2_u1_u7_n162, u2_u1_u7_n163, u2_u1_u7_n164, u2_u1_u7_n165, u2_u1_u7_n166, u2_u1_u7_n167, u2_u1_u7_n168, 
       u2_u1_u7_n169, u2_u1_u7_n170, u2_u1_u7_n171, u2_u1_u7_n172, u2_u1_u7_n173, u2_u1_u7_n174, u2_u1_u7_n175, u2_u1_u7_n176, u2_u1_u7_n177, 
       u2_u1_u7_n178, u2_u1_u7_n179, u2_u1_u7_n180, u2_u1_u7_n91, u2_u1_u7_n92, u2_u1_u7_n93, u2_u1_u7_n94, u2_u1_u7_n95, u2_u1_u7_n96, 
       u2_u1_u7_n97, u2_u1_u7_n98,  u2_u1_u7_n99;
  XOR2_X1 u0_U136 (.B( u0_L0_10 ) , .Z( u0_N41 ) , .A( u0_out1_10 ) );
  XOR2_X1 u0_U15 (.B( u0_L1_25 ) , .Z( u0_N88 ) , .A( u0_out2_25 ) );
  XOR2_X1 u0_U167 (.B( u0_L10_31 ) , .Z( u0_N382 ) , .A( u0_out11_31 ) );
  XOR2_X1 u0_U169 (.B( u0_L10_29 ) , .Z( u0_N380 ) , .A( u0_out11_29 ) );
  XOR2_X1 u0_U176 (.B( u0_L10_23 ) , .Z( u0_N374 ) , .A( u0_out11_23 ) );
  XOR2_X1 u0_U180 (.B( u0_L10_19 ) , .Z( u0_N370 ) , .A( u0_out11_19 ) );
  XOR2_X1 u0_U183 (.B( u0_L10_17 ) , .Z( u0_N368 ) , .A( u0_out11_17 ) );
  XOR2_X1 u0_U189 (.B( u0_L10_11 ) , .Z( u0_N362 ) , .A( u0_out11_11 ) );
  XOR2_X1 u0_U191 (.B( u0_L10_9 ) , .Z( u0_N360 ) , .A( u0_out11_9 ) );
  XOR2_X1 u0_U197 (.B( u0_L10_4 ) , .Z( u0_N355 ) , .A( u0_out11_4 ) );
  XOR2_X1 u0_U236 (.B( u0_L0_1 ) , .Z( u0_N32 ) , .A( u0_out1_1 ) );
  XOR2_X1 u0_U27 (.B( u0_L1_14 ) , .Z( u0_N77 ) , .A( u0_out2_14 ) );
  XOR2_X1 u0_U308 (.B( u0_L6_32 ) , .Z( u0_N255 ) , .A( u0_out7_32 ) );
  XOR2_X1 u0_U309 (.B( u0_L6_31 ) , .Z( u0_N254 ) , .A( u0_out7_31 ) );
  XOR2_X1 u0_U310 (.B( u0_L6_30 ) , .Z( u0_N253 ) , .A( u0_out7_30 ) );
  XOR2_X1 u0_U311 (.B( u0_L6_29 ) , .Z( u0_N252 ) , .A( u0_out7_29 ) );
  XOR2_X1 u0_U312 (.B( u0_L6_28 ) , .Z( u0_N251 ) , .A( u0_out7_28 ) );
  XOR2_X1 u0_U313 (.B( u0_L6_27 ) , .Z( u0_N250 ) , .A( u0_out7_27 ) );
  XOR2_X1 u0_U315 (.B( u0_L6_26 ) , .Z( u0_N249 ) , .A( u0_out7_26 ) );
  XOR2_X1 u0_U316 (.B( u0_L6_25 ) , .Z( u0_N248 ) , .A( u0_out7_25 ) );
  XOR2_X1 u0_U317 (.B( u0_L6_24 ) , .Z( u0_N247 ) , .A( u0_out7_24 ) );
  XOR2_X1 u0_U318 (.B( u0_L6_23 ) , .Z( u0_N246 ) , .A( u0_out7_23 ) );
  XOR2_X1 u0_U319 (.B( u0_L6_22 ) , .Z( u0_N245 ) , .A( u0_out7_22 ) );
  XOR2_X1 u0_U320 (.B( u0_L6_21 ) , .Z( u0_N244 ) , .A( u0_out7_21 ) );
  XOR2_X1 u0_U321 (.B( u0_L6_20 ) , .Z( u0_N243 ) , .A( u0_out7_20 ) );
  XOR2_X1 u0_U322 (.B( u0_L6_19 ) , .Z( u0_N242 ) , .A( u0_out7_19 ) );
  XOR2_X1 u0_U323 (.B( u0_L6_18 ) , .Z( u0_N241 ) , .A( u0_out7_18 ) );
  XOR2_X1 u0_U324 (.B( u0_L6_17 ) , .Z( u0_N240 ) , .A( u0_out7_17 ) );
  XOR2_X1 u0_U326 (.B( u0_L6_16 ) , .Z( u0_N239 ) , .A( u0_out7_16 ) );
  XOR2_X1 u0_U327 (.B( u0_L6_15 ) , .Z( u0_N238 ) , .A( u0_out7_15 ) );
  XOR2_X1 u0_U328 (.B( u0_L6_14 ) , .Z( u0_N237 ) , .A( u0_out7_14 ) );
  XOR2_X1 u0_U329 (.B( u0_L6_13 ) , .Z( u0_N236 ) , .A( u0_out7_13 ) );
  XOR2_X1 u0_U33 (.B( u0_L1_8 ) , .Z( u0_N71 ) , .A( u0_out2_8 ) );
  XOR2_X1 u0_U330 (.B( u0_L6_12 ) , .Z( u0_N235 ) , .A( u0_out7_12 ) );
  XOR2_X1 u0_U331 (.B( u0_L6_11 ) , .Z( u0_N234 ) , .A( u0_out7_11 ) );
  XOR2_X1 u0_U332 (.B( u0_L6_10 ) , .Z( u0_N233 ) , .A( u0_out7_10 ) );
  XOR2_X1 u0_U333 (.B( u0_L6_9 ) , .Z( u0_N232 ) , .A( u0_out7_9 ) );
  XOR2_X1 u0_U334 (.B( u0_L6_8 ) , .Z( u0_N231 ) , .A( u0_out7_8 ) );
  XOR2_X1 u0_U335 (.B( u0_L6_7 ) , .Z( u0_N230 ) , .A( u0_out7_7 ) );
  XOR2_X1 u0_U337 (.B( u0_L6_6 ) , .Z( u0_N229 ) , .A( u0_out7_6 ) );
  XOR2_X1 u0_U338 (.B( u0_L6_5 ) , .Z( u0_N228 ) , .A( u0_out7_5 ) );
  XOR2_X1 u0_U339 (.B( u0_L6_4 ) , .Z( u0_N227 ) , .A( u0_out7_4 ) );
  XOR2_X1 u0_U340 (.B( u0_L6_3 ) , .Z( u0_N226 ) , .A( u0_out7_3 ) );
  XOR2_X1 u0_U341 (.B( u0_L6_2 ) , .Z( u0_N225 ) , .A( u0_out7_2 ) );
  XOR2_X1 u0_U342 (.B( u0_L6_1 ) , .Z( u0_N224 ) , .A( u0_out7_1 ) );
  XOR2_X1 u0_U380 (.B( u0_L4_31 ) , .Z( u0_N190 ) , .A( u0_out5_31 ) );
  XOR2_X1 u0_U382 (.B( u0_L4_30 ) , .Z( u0_N189 ) , .A( u0_out5_30 ) );
  XOR2_X1 u0_U383 (.B( u0_L4_29 ) , .Z( u0_N188 ) , .A( u0_out5_29 ) );
  XOR2_X1 u0_U384 (.B( u0_L4_28 ) , .Z( u0_N187 ) , .A( u0_out5_28 ) );
  XOR2_X1 u0_U385 (.B( u0_L4_27 ) , .Z( u0_N186 ) , .A( u0_out5_27 ) );
  XOR2_X1 u0_U386 (.B( u0_L4_26 ) , .Z( u0_N185 ) , .A( u0_out5_26 ) );
  XOR2_X1 u0_U388 (.B( u0_L4_24 ) , .Z( u0_N183 ) , .A( u0_out5_24 ) );
  XOR2_X1 u0_U389 (.B( u0_L4_23 ) , .Z( u0_N182 ) , .A( u0_out5_23 ) );
  XOR2_X1 u0_U39 (.B( u0_L1_3 ) , .Z( u0_N66 ) , .A( u0_out2_3 ) );
  XOR2_X1 u0_U391 (.B( u0_L4_21 ) , .Z( u0_N180 ) , .A( u0_out5_21 ) );
  XOR2_X1 u0_U393 (.B( u0_L4_20 ) , .Z( u0_N179 ) , .A( u0_out5_20 ) );
  XOR2_X1 u0_U394 (.B( u0_L4_19 ) , .Z( u0_N178 ) , .A( u0_out5_19 ) );
  XOR2_X1 u0_U395 (.B( u0_L4_18 ) , .Z( u0_N177 ) , .A( u0_out5_18 ) );
  XOR2_X1 u0_U396 (.B( u0_L4_17 ) , .Z( u0_N176 ) , .A( u0_out5_17 ) );
  XOR2_X1 u0_U397 (.B( u0_L4_16 ) , .Z( u0_N175 ) , .A( u0_out5_16 ) );
  XOR2_X1 u0_U398 (.B( u0_L4_15 ) , .Z( u0_N174 ) , .A( u0_out5_15 ) );
  XOR2_X1 u0_U400 (.B( u0_L4_13 ) , .Z( u0_N172 ) , .A( u0_out5_13 ) );
  XOR2_X1 u0_U402 (.B( u0_L4_11 ) , .Z( u0_N170 ) , .A( u0_out5_11 ) );
  XOR2_X1 u0_U404 (.B( u0_L4_10 ) , .Z( u0_N169 ) , .A( u0_out5_10 ) );
  XOR2_X1 u0_U405 (.B( u0_L4_9 ) , .Z( u0_N168 ) , .A( u0_out5_9 ) );
  XOR2_X1 u0_U408 (.B( u0_L4_6 ) , .Z( u0_N165 ) , .A( u0_out5_6 ) );
  XOR2_X1 u0_U409 (.B( u0_L4_5 ) , .Z( u0_N164 ) , .A( u0_out5_5 ) );
  XOR2_X1 u0_U410 (.B( u0_L4_4 ) , .Z( u0_N163 ) , .A( u0_out5_4 ) );
  XOR2_X1 u0_U412 (.B( u0_L4_2 ) , .Z( u0_N161 ) , .A( u0_out5_2 ) );
  XOR2_X1 u0_U413 (.B( u0_L4_1 ) , .Z( u0_N160 ) , .A( u0_out5_1 ) );
  XOR2_X1 u0_U450 (.B( u0_L2_32 ) , .Z( u0_N127 ) , .A( u0_out3_32 ) );
  XOR2_X1 u0_U455 (.B( u0_L2_27 ) , .Z( u0_N122 ) , .A( u0_out3_27 ) );
  XOR2_X1 u0_U461 (.B( u0_L2_22 ) , .Z( u0_N117 ) , .A( u0_out3_22 ) );
  XOR2_X1 u0_U462 (.B( u0_L2_21 ) , .Z( u0_N116 ) , .A( u0_out3_21 ) );
  XOR2_X1 u0_U468 (.B( u0_L2_15 ) , .Z( u0_N110 ) , .A( u0_out3_15 ) );
  XOR2_X1 u0_U472 (.B( u0_L2_12 ) , .Z( u0_N107 ) , .A( u0_out3_12 ) );
  XOR2_X1 u0_U477 (.B( u0_L2_7 ) , .Z( u0_N102 ) , .A( u0_out3_7 ) );
  XOR2_X1 u0_U479 (.B( u0_L2_5 ) , .Z( u0_N100 ) , .A( u0_out3_5 ) );
  XOR2_X1 u0_U49 (.B( u0_L0_26 ) , .Z( u0_N57 ) , .A( u0_out1_26 ) );
  XOR2_X1 u0_U55 (.B( u0_L0_20 ) , .Z( u0_N51 ) , .A( u0_out1_20 ) );
  XOR2_X1 u0_u11_U16 (.B( u0_K12_3 ) , .A( u0_R10_2 ) , .Z( u0_u11_X_3 ) );
  XOR2_X1 u0_u11_U20 (.B( u0_K12_36 ) , .A( u0_R10_25 ) , .Z( u0_u11_X_36 ) );
  XOR2_X1 u0_u11_U21 (.B( u0_K12_35 ) , .A( u0_R10_24 ) , .Z( u0_u11_X_35 ) );
  XOR2_X1 u0_u11_U22 (.B( u0_K12_34 ) , .A( u0_R10_23 ) , .Z( u0_u11_X_34 ) );
  XOR2_X1 u0_u11_U23 (.B( u0_K12_33 ) , .A( u0_R10_22 ) , .Z( u0_u11_X_33 ) );
  XOR2_X1 u0_u11_U24 (.B( u0_K12_32 ) , .A( u0_R10_21 ) , .Z( u0_u11_X_32 ) );
  XOR2_X1 u0_u11_U25 (.B( u0_K12_31 ) , .A( u0_R10_20 ) , .Z( u0_u11_X_31 ) );
  XOR2_X1 u0_u11_U27 (.B( u0_K12_2 ) , .A( u0_R10_1 ) , .Z( u0_u11_X_2 ) );
  XOR2_X1 u0_u11_U38 (.B( u0_K12_1 ) , .A( u0_R10_32 ) , .Z( u0_u11_X_1 ) );
  XOR2_X1 u0_u11_U4 (.B( u0_K12_6 ) , .A( u0_R10_5 ) , .Z( u0_u11_X_6 ) );
  XOR2_X1 u0_u11_U5 (.B( u0_K12_5 ) , .A( u0_R10_4 ) , .Z( u0_u11_X_5 ) );
  XOR2_X1 u0_u11_U6 (.B( u0_K12_4 ) , .A( u0_R10_3 ) , .Z( u0_u11_X_4 ) );
  AND3_X1 u0_u11_u0_U10 (.A2( u0_u11_u0_n112 ) , .ZN( u0_u11_u0_n127 ) , .A3( u0_u11_u0_n130 ) , .A1( u0_u11_u0_n148 ) );
  NAND2_X1 u0_u11_u0_U11 (.ZN( u0_u11_u0_n113 ) , .A1( u0_u11_u0_n139 ) , .A2( u0_u11_u0_n149 ) );
  AND2_X1 u0_u11_u0_U12 (.ZN( u0_u11_u0_n107 ) , .A1( u0_u11_u0_n130 ) , .A2( u0_u11_u0_n140 ) );
  AND2_X1 u0_u11_u0_U13 (.A2( u0_u11_u0_n129 ) , .A1( u0_u11_u0_n130 ) , .ZN( u0_u11_u0_n151 ) );
  AND2_X1 u0_u11_u0_U14 (.A1( u0_u11_u0_n108 ) , .A2( u0_u11_u0_n125 ) , .ZN( u0_u11_u0_n145 ) );
  INV_X1 u0_u11_u0_U15 (.A( u0_u11_u0_n143 ) , .ZN( u0_u11_u0_n173 ) );
  NOR2_X1 u0_u11_u0_U16 (.A2( u0_u11_u0_n136 ) , .ZN( u0_u11_u0_n147 ) , .A1( u0_u11_u0_n160 ) );
  AOI21_X1 u0_u11_u0_U17 (.B1( u0_u11_u0_n103 ) , .ZN( u0_u11_u0_n132 ) , .A( u0_u11_u0_n165 ) , .B2( u0_u11_u0_n93 ) );
  INV_X1 u0_u11_u0_U18 (.A( u0_u11_u0_n142 ) , .ZN( u0_u11_u0_n165 ) );
  OAI22_X1 u0_u11_u0_U19 (.B1( u0_u11_u0_n125 ) , .ZN( u0_u11_u0_n126 ) , .A1( u0_u11_u0_n138 ) , .A2( u0_u11_u0_n146 ) , .B2( u0_u11_u0_n147 ) );
  OAI22_X1 u0_u11_u0_U20 (.B1( u0_u11_u0_n131 ) , .A1( u0_u11_u0_n144 ) , .B2( u0_u11_u0_n147 ) , .A2( u0_u11_u0_n90 ) , .ZN( u0_u11_u0_n91 ) );
  AND3_X1 u0_u11_u0_U21 (.A3( u0_u11_u0_n121 ) , .A2( u0_u11_u0_n125 ) , .A1( u0_u11_u0_n148 ) , .ZN( u0_u11_u0_n90 ) );
  INV_X1 u0_u11_u0_U22 (.A( u0_u11_u0_n136 ) , .ZN( u0_u11_u0_n161 ) );
  AOI22_X1 u0_u11_u0_U23 (.B2( u0_u11_u0_n109 ) , .A2( u0_u11_u0_n110 ) , .ZN( u0_u11_u0_n111 ) , .B1( u0_u11_u0_n118 ) , .A1( u0_u11_u0_n160 ) );
  NAND2_X1 u0_u11_u0_U24 (.A1( u0_u11_u0_n100 ) , .A2( u0_u11_u0_n103 ) , .ZN( u0_u11_u0_n125 ) );
  INV_X1 u0_u11_u0_U25 (.A( u0_u11_u0_n118 ) , .ZN( u0_u11_u0_n158 ) );
  AOI21_X1 u0_u11_u0_U26 (.B1( u0_u11_u0_n127 ) , .B2( u0_u11_u0_n129 ) , .A( u0_u11_u0_n138 ) , .ZN( u0_u11_u0_n96 ) );
  AOI21_X1 u0_u11_u0_U27 (.ZN( u0_u11_u0_n104 ) , .B1( u0_u11_u0_n107 ) , .B2( u0_u11_u0_n141 ) , .A( u0_u11_u0_n144 ) );
  AOI21_X1 u0_u11_u0_U28 (.ZN( u0_u11_u0_n116 ) , .B2( u0_u11_u0_n142 ) , .A( u0_u11_u0_n144 ) , .B1( u0_u11_u0_n166 ) );
  NOR2_X1 u0_u11_u0_U29 (.A1( u0_u11_u0_n120 ) , .ZN( u0_u11_u0_n143 ) , .A2( u0_u11_u0_n167 ) );
  INV_X1 u0_u11_u0_U3 (.A( u0_u11_u0_n113 ) , .ZN( u0_u11_u0_n166 ) );
  OAI221_X1 u0_u11_u0_U30 (.C1( u0_u11_u0_n112 ) , .ZN( u0_u11_u0_n120 ) , .B1( u0_u11_u0_n138 ) , .B2( u0_u11_u0_n141 ) , .C2( u0_u11_u0_n147 ) , .A( u0_u11_u0_n172 ) );
  AOI211_X1 u0_u11_u0_U31 (.B( u0_u11_u0_n115 ) , .A( u0_u11_u0_n116 ) , .C2( u0_u11_u0_n117 ) , .C1( u0_u11_u0_n118 ) , .ZN( u0_u11_u0_n119 ) );
  NAND2_X1 u0_u11_u0_U32 (.A2( u0_u11_u0_n103 ) , .ZN( u0_u11_u0_n140 ) , .A1( u0_u11_u0_n94 ) );
  NAND2_X1 u0_u11_u0_U33 (.A1( u0_u11_u0_n101 ) , .A2( u0_u11_u0_n102 ) , .ZN( u0_u11_u0_n150 ) );
  INV_X1 u0_u11_u0_U34 (.A( u0_u11_u0_n138 ) , .ZN( u0_u11_u0_n160 ) );
  NAND2_X1 u0_u11_u0_U35 (.A2( u0_u11_u0_n100 ) , .A1( u0_u11_u0_n101 ) , .ZN( u0_u11_u0_n139 ) );
  NAND2_X1 u0_u11_u0_U36 (.A2( u0_u11_u0_n100 ) , .ZN( u0_u11_u0_n131 ) , .A1( u0_u11_u0_n92 ) );
  NAND2_X1 u0_u11_u0_U37 (.A2( u0_u11_u0_n102 ) , .A1( u0_u11_u0_n103 ) , .ZN( u0_u11_u0_n149 ) );
  NAND2_X1 u0_u11_u0_U38 (.ZN( u0_u11_u0_n108 ) , .A1( u0_u11_u0_n92 ) , .A2( u0_u11_u0_n94 ) );
  NAND2_X1 u0_u11_u0_U39 (.A2( u0_u11_u0_n102 ) , .ZN( u0_u11_u0_n114 ) , .A1( u0_u11_u0_n92 ) );
  AOI21_X1 u0_u11_u0_U4 (.B1( u0_u11_u0_n114 ) , .ZN( u0_u11_u0_n115 ) , .B2( u0_u11_u0_n129 ) , .A( u0_u11_u0_n161 ) );
  NAND2_X1 u0_u11_u0_U40 (.A1( u0_u11_u0_n101 ) , .ZN( u0_u11_u0_n130 ) , .A2( u0_u11_u0_n94 ) );
  INV_X1 u0_u11_u0_U41 (.ZN( u0_u11_u0_n172 ) , .A( u0_u11_u0_n88 ) );
  OAI222_X1 u0_u11_u0_U42 (.C1( u0_u11_u0_n108 ) , .A1( u0_u11_u0_n125 ) , .B2( u0_u11_u0_n128 ) , .B1( u0_u11_u0_n144 ) , .A2( u0_u11_u0_n158 ) , .C2( u0_u11_u0_n161 ) , .ZN( u0_u11_u0_n88 ) );
  NAND2_X1 u0_u11_u0_U43 (.ZN( u0_u11_u0_n112 ) , .A2( u0_u11_u0_n92 ) , .A1( u0_u11_u0_n93 ) );
  NAND2_X1 u0_u11_u0_U44 (.A2( u0_u11_u0_n101 ) , .ZN( u0_u11_u0_n121 ) , .A1( u0_u11_u0_n93 ) );
  OR3_X1 u0_u11_u0_U45 (.A3( u0_u11_u0_n152 ) , .A2( u0_u11_u0_n153 ) , .A1( u0_u11_u0_n154 ) , .ZN( u0_u11_u0_n155 ) );
  AOI21_X1 u0_u11_u0_U46 (.A( u0_u11_u0_n144 ) , .B2( u0_u11_u0_n145 ) , .B1( u0_u11_u0_n146 ) , .ZN( u0_u11_u0_n154 ) );
  AOI21_X1 u0_u11_u0_U47 (.B2( u0_u11_u0_n150 ) , .B1( u0_u11_u0_n151 ) , .ZN( u0_u11_u0_n152 ) , .A( u0_u11_u0_n158 ) );
  AOI21_X1 u0_u11_u0_U48 (.A( u0_u11_u0_n147 ) , .B2( u0_u11_u0_n148 ) , .B1( u0_u11_u0_n149 ) , .ZN( u0_u11_u0_n153 ) );
  INV_X1 u0_u11_u0_U49 (.ZN( u0_u11_u0_n171 ) , .A( u0_u11_u0_n99 ) );
  AOI21_X1 u0_u11_u0_U5 (.B2( u0_u11_u0_n131 ) , .ZN( u0_u11_u0_n134 ) , .B1( u0_u11_u0_n151 ) , .A( u0_u11_u0_n158 ) );
  OAI211_X1 u0_u11_u0_U50 (.C2( u0_u11_u0_n140 ) , .C1( u0_u11_u0_n161 ) , .A( u0_u11_u0_n169 ) , .B( u0_u11_u0_n98 ) , .ZN( u0_u11_u0_n99 ) );
  AOI211_X1 u0_u11_u0_U51 (.C1( u0_u11_u0_n118 ) , .A( u0_u11_u0_n123 ) , .B( u0_u11_u0_n96 ) , .C2( u0_u11_u0_n97 ) , .ZN( u0_u11_u0_n98 ) );
  INV_X1 u0_u11_u0_U52 (.ZN( u0_u11_u0_n169 ) , .A( u0_u11_u0_n91 ) );
  NOR2_X1 u0_u11_u0_U53 (.A2( u0_u11_X_2 ) , .ZN( u0_u11_u0_n103 ) , .A1( u0_u11_u0_n164 ) );
  NOR2_X1 u0_u11_u0_U54 (.A2( u0_u11_X_4 ) , .A1( u0_u11_X_5 ) , .ZN( u0_u11_u0_n118 ) );
  NOR2_X1 u0_u11_u0_U55 (.A2( u0_u11_X_1 ) , .A1( u0_u11_X_2 ) , .ZN( u0_u11_u0_n92 ) );
  NOR2_X1 u0_u11_u0_U56 (.A2( u0_u11_X_1 ) , .ZN( u0_u11_u0_n101 ) , .A1( u0_u11_u0_n163 ) );
  NOR2_X1 u0_u11_u0_U57 (.A2( u0_u11_X_3 ) , .A1( u0_u11_X_6 ) , .ZN( u0_u11_u0_n94 ) );
  NAND2_X1 u0_u11_u0_U58 (.A2( u0_u11_X_4 ) , .A1( u0_u11_X_5 ) , .ZN( u0_u11_u0_n144 ) );
  NOR2_X1 u0_u11_u0_U59 (.A2( u0_u11_X_5 ) , .ZN( u0_u11_u0_n136 ) , .A1( u0_u11_u0_n159 ) );
  NOR2_X1 u0_u11_u0_U6 (.A1( u0_u11_u0_n108 ) , .ZN( u0_u11_u0_n123 ) , .A2( u0_u11_u0_n158 ) );
  NAND2_X1 u0_u11_u0_U60 (.A1( u0_u11_X_5 ) , .ZN( u0_u11_u0_n138 ) , .A2( u0_u11_u0_n159 ) );
  AND2_X1 u0_u11_u0_U61 (.A2( u0_u11_X_3 ) , .A1( u0_u11_X_6 ) , .ZN( u0_u11_u0_n102 ) );
  AND2_X1 u0_u11_u0_U62 (.A1( u0_u11_X_6 ) , .A2( u0_u11_u0_n162 ) , .ZN( u0_u11_u0_n93 ) );
  INV_X1 u0_u11_u0_U63 (.A( u0_u11_X_4 ) , .ZN( u0_u11_u0_n159 ) );
  INV_X1 u0_u11_u0_U64 (.A( u0_u11_X_2 ) , .ZN( u0_u11_u0_n163 ) );
  INV_X1 u0_u11_u0_U65 (.A( u0_u11_X_1 ) , .ZN( u0_u11_u0_n164 ) );
  INV_X1 u0_u11_u0_U66 (.A( u0_u11_u0_n126 ) , .ZN( u0_u11_u0_n168 ) );
  AOI211_X1 u0_u11_u0_U67 (.B( u0_u11_u0_n133 ) , .A( u0_u11_u0_n134 ) , .C2( u0_u11_u0_n135 ) , .C1( u0_u11_u0_n136 ) , .ZN( u0_u11_u0_n137 ) );
  OR4_X1 u0_u11_u0_U68 (.ZN( u0_out11_17 ) , .A4( u0_u11_u0_n122 ) , .A2( u0_u11_u0_n123 ) , .A1( u0_u11_u0_n124 ) , .A3( u0_u11_u0_n170 ) );
  AOI21_X1 u0_u11_u0_U69 (.B2( u0_u11_u0_n107 ) , .ZN( u0_u11_u0_n124 ) , .B1( u0_u11_u0_n128 ) , .A( u0_u11_u0_n161 ) );
  OAI21_X1 u0_u11_u0_U7 (.B1( u0_u11_u0_n150 ) , .B2( u0_u11_u0_n158 ) , .A( u0_u11_u0_n172 ) , .ZN( u0_u11_u0_n89 ) );
  INV_X1 u0_u11_u0_U70 (.A( u0_u11_u0_n111 ) , .ZN( u0_u11_u0_n170 ) );
  OR4_X1 u0_u11_u0_U71 (.ZN( u0_out11_31 ) , .A4( u0_u11_u0_n155 ) , .A2( u0_u11_u0_n156 ) , .A1( u0_u11_u0_n157 ) , .A3( u0_u11_u0_n173 ) );
  AOI21_X1 u0_u11_u0_U72 (.A( u0_u11_u0_n138 ) , .B2( u0_u11_u0_n139 ) , .B1( u0_u11_u0_n140 ) , .ZN( u0_u11_u0_n157 ) );
  AOI21_X1 u0_u11_u0_U73 (.B2( u0_u11_u0_n141 ) , .B1( u0_u11_u0_n142 ) , .ZN( u0_u11_u0_n156 ) , .A( u0_u11_u0_n161 ) );
  INV_X1 u0_u11_u0_U74 (.ZN( u0_u11_u0_n174 ) , .A( u0_u11_u0_n89 ) );
  AOI211_X1 u0_u11_u0_U75 (.B( u0_u11_u0_n104 ) , .A( u0_u11_u0_n105 ) , .ZN( u0_u11_u0_n106 ) , .C2( u0_u11_u0_n113 ) , .C1( u0_u11_u0_n160 ) );
  NOR2_X1 u0_u11_u0_U76 (.A2( u0_u11_X_6 ) , .ZN( u0_u11_u0_n100 ) , .A1( u0_u11_u0_n162 ) );
  INV_X1 u0_u11_u0_U77 (.A( u0_u11_X_3 ) , .ZN( u0_u11_u0_n162 ) );
  NOR2_X1 u0_u11_u0_U78 (.A1( u0_u11_u0_n163 ) , .A2( u0_u11_u0_n164 ) , .ZN( u0_u11_u0_n95 ) );
  OAI221_X1 u0_u11_u0_U79 (.C1( u0_u11_u0_n121 ) , .ZN( u0_u11_u0_n122 ) , .B2( u0_u11_u0_n127 ) , .A( u0_u11_u0_n143 ) , .B1( u0_u11_u0_n144 ) , .C2( u0_u11_u0_n147 ) );
  AND2_X1 u0_u11_u0_U8 (.A1( u0_u11_u0_n114 ) , .A2( u0_u11_u0_n121 ) , .ZN( u0_u11_u0_n146 ) );
  AOI21_X1 u0_u11_u0_U80 (.B1( u0_u11_u0_n132 ) , .ZN( u0_u11_u0_n133 ) , .A( u0_u11_u0_n144 ) , .B2( u0_u11_u0_n166 ) );
  OAI22_X1 u0_u11_u0_U81 (.ZN( u0_u11_u0_n105 ) , .A2( u0_u11_u0_n132 ) , .B1( u0_u11_u0_n146 ) , .A1( u0_u11_u0_n147 ) , .B2( u0_u11_u0_n161 ) );
  NAND2_X1 u0_u11_u0_U82 (.ZN( u0_u11_u0_n110 ) , .A2( u0_u11_u0_n132 ) , .A1( u0_u11_u0_n145 ) );
  INV_X1 u0_u11_u0_U83 (.A( u0_u11_u0_n119 ) , .ZN( u0_u11_u0_n167 ) );
  NAND2_X1 u0_u11_u0_U84 (.ZN( u0_u11_u0_n148 ) , .A1( u0_u11_u0_n93 ) , .A2( u0_u11_u0_n95 ) );
  NAND2_X1 u0_u11_u0_U85 (.A1( u0_u11_u0_n100 ) , .ZN( u0_u11_u0_n129 ) , .A2( u0_u11_u0_n95 ) );
  NAND2_X1 u0_u11_u0_U86 (.A1( u0_u11_u0_n102 ) , .ZN( u0_u11_u0_n128 ) , .A2( u0_u11_u0_n95 ) );
  NAND2_X1 u0_u11_u0_U87 (.ZN( u0_u11_u0_n142 ) , .A1( u0_u11_u0_n94 ) , .A2( u0_u11_u0_n95 ) );
  NAND3_X1 u0_u11_u0_U88 (.ZN( u0_out11_23 ) , .A3( u0_u11_u0_n137 ) , .A1( u0_u11_u0_n168 ) , .A2( u0_u11_u0_n171 ) );
  NAND3_X1 u0_u11_u0_U89 (.A3( u0_u11_u0_n127 ) , .A2( u0_u11_u0_n128 ) , .ZN( u0_u11_u0_n135 ) , .A1( u0_u11_u0_n150 ) );
  AND2_X1 u0_u11_u0_U9 (.A1( u0_u11_u0_n131 ) , .ZN( u0_u11_u0_n141 ) , .A2( u0_u11_u0_n150 ) );
  NAND3_X1 u0_u11_u0_U90 (.ZN( u0_u11_u0_n117 ) , .A3( u0_u11_u0_n132 ) , .A2( u0_u11_u0_n139 ) , .A1( u0_u11_u0_n148 ) );
  NAND3_X1 u0_u11_u0_U91 (.ZN( u0_u11_u0_n109 ) , .A2( u0_u11_u0_n114 ) , .A3( u0_u11_u0_n140 ) , .A1( u0_u11_u0_n149 ) );
  NAND3_X1 u0_u11_u0_U92 (.ZN( u0_out11_9 ) , .A3( u0_u11_u0_n106 ) , .A2( u0_u11_u0_n171 ) , .A1( u0_u11_u0_n174 ) );
  NAND3_X1 u0_u11_u0_U93 (.A2( u0_u11_u0_n128 ) , .A1( u0_u11_u0_n132 ) , .A3( u0_u11_u0_n146 ) , .ZN( u0_u11_u0_n97 ) );
  INV_X1 u0_u11_u5_U10 (.A( u0_u11_u5_n121 ) , .ZN( u0_u11_u5_n177 ) );
  NOR3_X1 u0_u11_u5_U100 (.A3( u0_u11_u5_n141 ) , .A1( u0_u11_u5_n142 ) , .ZN( u0_u11_u5_n143 ) , .A2( u0_u11_u5_n191 ) );
  NAND4_X1 u0_u11_u5_U101 (.ZN( u0_out11_4 ) , .A4( u0_u11_u5_n112 ) , .A2( u0_u11_u5_n113 ) , .A1( u0_u11_u5_n114 ) , .A3( u0_u11_u5_n195 ) );
  AOI211_X1 u0_u11_u5_U102 (.A( u0_u11_u5_n110 ) , .C1( u0_u11_u5_n111 ) , .ZN( u0_u11_u5_n112 ) , .B( u0_u11_u5_n118 ) , .C2( u0_u11_u5_n177 ) );
  AOI222_X1 u0_u11_u5_U103 (.ZN( u0_u11_u5_n113 ) , .A1( u0_u11_u5_n131 ) , .C1( u0_u11_u5_n148 ) , .B2( u0_u11_u5_n174 ) , .C2( u0_u11_u5_n178 ) , .A2( u0_u11_u5_n179 ) , .B1( u0_u11_u5_n99 ) );
  NAND3_X1 u0_u11_u5_U104 (.A2( u0_u11_u5_n154 ) , .A3( u0_u11_u5_n158 ) , .A1( u0_u11_u5_n161 ) , .ZN( u0_u11_u5_n99 ) );
  NOR2_X1 u0_u11_u5_U11 (.ZN( u0_u11_u5_n160 ) , .A2( u0_u11_u5_n173 ) , .A1( u0_u11_u5_n177 ) );
  INV_X1 u0_u11_u5_U12 (.A( u0_u11_u5_n150 ) , .ZN( u0_u11_u5_n174 ) );
  AOI21_X1 u0_u11_u5_U13 (.A( u0_u11_u5_n160 ) , .B2( u0_u11_u5_n161 ) , .ZN( u0_u11_u5_n162 ) , .B1( u0_u11_u5_n192 ) );
  INV_X1 u0_u11_u5_U14 (.A( u0_u11_u5_n159 ) , .ZN( u0_u11_u5_n192 ) );
  AOI21_X1 u0_u11_u5_U15 (.A( u0_u11_u5_n156 ) , .B2( u0_u11_u5_n157 ) , .B1( u0_u11_u5_n158 ) , .ZN( u0_u11_u5_n163 ) );
  AOI21_X1 u0_u11_u5_U16 (.B2( u0_u11_u5_n139 ) , .B1( u0_u11_u5_n140 ) , .ZN( u0_u11_u5_n141 ) , .A( u0_u11_u5_n150 ) );
  OAI21_X1 u0_u11_u5_U17 (.A( u0_u11_u5_n133 ) , .B2( u0_u11_u5_n134 ) , .B1( u0_u11_u5_n135 ) , .ZN( u0_u11_u5_n142 ) );
  OAI21_X1 u0_u11_u5_U18 (.ZN( u0_u11_u5_n133 ) , .B2( u0_u11_u5_n147 ) , .A( u0_u11_u5_n173 ) , .B1( u0_u11_u5_n188 ) );
  NAND2_X1 u0_u11_u5_U19 (.A2( u0_u11_u5_n119 ) , .A1( u0_u11_u5_n123 ) , .ZN( u0_u11_u5_n137 ) );
  INV_X1 u0_u11_u5_U20 (.A( u0_u11_u5_n155 ) , .ZN( u0_u11_u5_n194 ) );
  NAND2_X1 u0_u11_u5_U21 (.A1( u0_u11_u5_n121 ) , .ZN( u0_u11_u5_n132 ) , .A2( u0_u11_u5_n172 ) );
  NAND2_X1 u0_u11_u5_U22 (.A2( u0_u11_u5_n122 ) , .ZN( u0_u11_u5_n136 ) , .A1( u0_u11_u5_n154 ) );
  NAND2_X1 u0_u11_u5_U23 (.A2( u0_u11_u5_n119 ) , .A1( u0_u11_u5_n120 ) , .ZN( u0_u11_u5_n159 ) );
  INV_X1 u0_u11_u5_U24 (.A( u0_u11_u5_n156 ) , .ZN( u0_u11_u5_n175 ) );
  INV_X1 u0_u11_u5_U25 (.A( u0_u11_u5_n158 ) , .ZN( u0_u11_u5_n188 ) );
  INV_X1 u0_u11_u5_U26 (.A( u0_u11_u5_n152 ) , .ZN( u0_u11_u5_n179 ) );
  INV_X1 u0_u11_u5_U27 (.A( u0_u11_u5_n140 ) , .ZN( u0_u11_u5_n182 ) );
  INV_X1 u0_u11_u5_U28 (.A( u0_u11_u5_n151 ) , .ZN( u0_u11_u5_n183 ) );
  INV_X1 u0_u11_u5_U29 (.A( u0_u11_u5_n123 ) , .ZN( u0_u11_u5_n185 ) );
  NOR2_X1 u0_u11_u5_U3 (.ZN( u0_u11_u5_n134 ) , .A1( u0_u11_u5_n183 ) , .A2( u0_u11_u5_n190 ) );
  INV_X1 u0_u11_u5_U30 (.A( u0_u11_u5_n161 ) , .ZN( u0_u11_u5_n184 ) );
  INV_X1 u0_u11_u5_U31 (.A( u0_u11_u5_n139 ) , .ZN( u0_u11_u5_n189 ) );
  INV_X1 u0_u11_u5_U32 (.A( u0_u11_u5_n157 ) , .ZN( u0_u11_u5_n190 ) );
  INV_X1 u0_u11_u5_U33 (.A( u0_u11_u5_n120 ) , .ZN( u0_u11_u5_n193 ) );
  NAND2_X1 u0_u11_u5_U34 (.ZN( u0_u11_u5_n111 ) , .A1( u0_u11_u5_n140 ) , .A2( u0_u11_u5_n155 ) );
  NOR2_X1 u0_u11_u5_U35 (.ZN( u0_u11_u5_n100 ) , .A1( u0_u11_u5_n170 ) , .A2( u0_u11_u5_n180 ) );
  INV_X1 u0_u11_u5_U36 (.A( u0_u11_u5_n117 ) , .ZN( u0_u11_u5_n196 ) );
  OAI221_X1 u0_u11_u5_U37 (.A( u0_u11_u5_n116 ) , .ZN( u0_u11_u5_n117 ) , .B2( u0_u11_u5_n119 ) , .C1( u0_u11_u5_n153 ) , .C2( u0_u11_u5_n158 ) , .B1( u0_u11_u5_n172 ) );
  AOI222_X1 u0_u11_u5_U38 (.ZN( u0_u11_u5_n116 ) , .B2( u0_u11_u5_n145 ) , .C1( u0_u11_u5_n148 ) , .A2( u0_u11_u5_n174 ) , .C2( u0_u11_u5_n177 ) , .B1( u0_u11_u5_n187 ) , .A1( u0_u11_u5_n193 ) );
  INV_X1 u0_u11_u5_U39 (.A( u0_u11_u5_n115 ) , .ZN( u0_u11_u5_n187 ) );
  INV_X1 u0_u11_u5_U4 (.A( u0_u11_u5_n138 ) , .ZN( u0_u11_u5_n191 ) );
  AOI22_X1 u0_u11_u5_U40 (.B2( u0_u11_u5_n131 ) , .A2( u0_u11_u5_n146 ) , .ZN( u0_u11_u5_n169 ) , .B1( u0_u11_u5_n174 ) , .A1( u0_u11_u5_n185 ) );
  NOR2_X1 u0_u11_u5_U41 (.A1( u0_u11_u5_n146 ) , .ZN( u0_u11_u5_n150 ) , .A2( u0_u11_u5_n173 ) );
  AOI21_X1 u0_u11_u5_U42 (.A( u0_u11_u5_n118 ) , .B2( u0_u11_u5_n145 ) , .ZN( u0_u11_u5_n168 ) , .B1( u0_u11_u5_n186 ) );
  INV_X1 u0_u11_u5_U43 (.A( u0_u11_u5_n122 ) , .ZN( u0_u11_u5_n186 ) );
  NOR2_X1 u0_u11_u5_U44 (.A1( u0_u11_u5_n146 ) , .ZN( u0_u11_u5_n152 ) , .A2( u0_u11_u5_n176 ) );
  NOR2_X1 u0_u11_u5_U45 (.A1( u0_u11_u5_n115 ) , .ZN( u0_u11_u5_n118 ) , .A2( u0_u11_u5_n153 ) );
  NOR2_X1 u0_u11_u5_U46 (.A2( u0_u11_u5_n145 ) , .ZN( u0_u11_u5_n156 ) , .A1( u0_u11_u5_n174 ) );
  NOR2_X1 u0_u11_u5_U47 (.ZN( u0_u11_u5_n121 ) , .A2( u0_u11_u5_n145 ) , .A1( u0_u11_u5_n176 ) );
  AOI22_X1 u0_u11_u5_U48 (.ZN( u0_u11_u5_n114 ) , .A2( u0_u11_u5_n137 ) , .A1( u0_u11_u5_n145 ) , .B2( u0_u11_u5_n175 ) , .B1( u0_u11_u5_n193 ) );
  OAI211_X1 u0_u11_u5_U49 (.B( u0_u11_u5_n124 ) , .A( u0_u11_u5_n125 ) , .C2( u0_u11_u5_n126 ) , .C1( u0_u11_u5_n127 ) , .ZN( u0_u11_u5_n128 ) );
  OAI21_X1 u0_u11_u5_U5 (.B2( u0_u11_u5_n136 ) , .B1( u0_u11_u5_n137 ) , .ZN( u0_u11_u5_n138 ) , .A( u0_u11_u5_n177 ) );
  OAI21_X1 u0_u11_u5_U50 (.ZN( u0_u11_u5_n124 ) , .A( u0_u11_u5_n177 ) , .B2( u0_u11_u5_n183 ) , .B1( u0_u11_u5_n189 ) );
  NOR3_X1 u0_u11_u5_U51 (.ZN( u0_u11_u5_n127 ) , .A1( u0_u11_u5_n136 ) , .A3( u0_u11_u5_n148 ) , .A2( u0_u11_u5_n182 ) );
  OAI21_X1 u0_u11_u5_U52 (.ZN( u0_u11_u5_n125 ) , .A( u0_u11_u5_n174 ) , .B2( u0_u11_u5_n185 ) , .B1( u0_u11_u5_n190 ) );
  AOI21_X1 u0_u11_u5_U53 (.A( u0_u11_u5_n153 ) , .B2( u0_u11_u5_n154 ) , .B1( u0_u11_u5_n155 ) , .ZN( u0_u11_u5_n164 ) );
  AOI21_X1 u0_u11_u5_U54 (.ZN( u0_u11_u5_n110 ) , .B1( u0_u11_u5_n122 ) , .B2( u0_u11_u5_n139 ) , .A( u0_u11_u5_n153 ) );
  INV_X1 u0_u11_u5_U55 (.A( u0_u11_u5_n153 ) , .ZN( u0_u11_u5_n176 ) );
  INV_X1 u0_u11_u5_U56 (.A( u0_u11_u5_n126 ) , .ZN( u0_u11_u5_n173 ) );
  AND2_X1 u0_u11_u5_U57 (.A2( u0_u11_u5_n104 ) , .A1( u0_u11_u5_n107 ) , .ZN( u0_u11_u5_n147 ) );
  AND2_X1 u0_u11_u5_U58 (.A2( u0_u11_u5_n104 ) , .A1( u0_u11_u5_n108 ) , .ZN( u0_u11_u5_n148 ) );
  NAND2_X1 u0_u11_u5_U59 (.A1( u0_u11_u5_n105 ) , .A2( u0_u11_u5_n106 ) , .ZN( u0_u11_u5_n158 ) );
  INV_X1 u0_u11_u5_U6 (.A( u0_u11_u5_n135 ) , .ZN( u0_u11_u5_n178 ) );
  NAND2_X1 u0_u11_u5_U60 (.A2( u0_u11_u5_n108 ) , .A1( u0_u11_u5_n109 ) , .ZN( u0_u11_u5_n139 ) );
  NAND2_X1 u0_u11_u5_U61 (.A1( u0_u11_u5_n106 ) , .A2( u0_u11_u5_n108 ) , .ZN( u0_u11_u5_n119 ) );
  NAND2_X1 u0_u11_u5_U62 (.A2( u0_u11_u5_n103 ) , .A1( u0_u11_u5_n105 ) , .ZN( u0_u11_u5_n140 ) );
  NAND2_X1 u0_u11_u5_U63 (.A2( u0_u11_u5_n104 ) , .A1( u0_u11_u5_n105 ) , .ZN( u0_u11_u5_n155 ) );
  NAND2_X1 u0_u11_u5_U64 (.A2( u0_u11_u5_n106 ) , .A1( u0_u11_u5_n107 ) , .ZN( u0_u11_u5_n122 ) );
  NAND2_X1 u0_u11_u5_U65 (.A2( u0_u11_u5_n100 ) , .A1( u0_u11_u5_n106 ) , .ZN( u0_u11_u5_n115 ) );
  NAND2_X1 u0_u11_u5_U66 (.A2( u0_u11_u5_n100 ) , .A1( u0_u11_u5_n103 ) , .ZN( u0_u11_u5_n161 ) );
  NAND2_X1 u0_u11_u5_U67 (.A1( u0_u11_u5_n105 ) , .A2( u0_u11_u5_n109 ) , .ZN( u0_u11_u5_n154 ) );
  INV_X1 u0_u11_u5_U68 (.A( u0_u11_u5_n146 ) , .ZN( u0_u11_u5_n172 ) );
  NAND2_X1 u0_u11_u5_U69 (.A1( u0_u11_u5_n103 ) , .A2( u0_u11_u5_n108 ) , .ZN( u0_u11_u5_n123 ) );
  OAI22_X1 u0_u11_u5_U7 (.B2( u0_u11_u5_n149 ) , .B1( u0_u11_u5_n150 ) , .A2( u0_u11_u5_n151 ) , .A1( u0_u11_u5_n152 ) , .ZN( u0_u11_u5_n165 ) );
  NAND2_X1 u0_u11_u5_U70 (.A2( u0_u11_u5_n103 ) , .A1( u0_u11_u5_n107 ) , .ZN( u0_u11_u5_n151 ) );
  NAND2_X1 u0_u11_u5_U71 (.A2( u0_u11_u5_n107 ) , .A1( u0_u11_u5_n109 ) , .ZN( u0_u11_u5_n120 ) );
  NAND2_X1 u0_u11_u5_U72 (.A2( u0_u11_u5_n100 ) , .A1( u0_u11_u5_n109 ) , .ZN( u0_u11_u5_n157 ) );
  AND2_X1 u0_u11_u5_U73 (.A2( u0_u11_u5_n100 ) , .A1( u0_u11_u5_n104 ) , .ZN( u0_u11_u5_n131 ) );
  INV_X1 u0_u11_u5_U74 (.A( u0_u11_u5_n102 ) , .ZN( u0_u11_u5_n195 ) );
  OAI221_X1 u0_u11_u5_U75 (.A( u0_u11_u5_n101 ) , .ZN( u0_u11_u5_n102 ) , .C2( u0_u11_u5_n115 ) , .C1( u0_u11_u5_n126 ) , .B1( u0_u11_u5_n134 ) , .B2( u0_u11_u5_n160 ) );
  OAI21_X1 u0_u11_u5_U76 (.ZN( u0_u11_u5_n101 ) , .B1( u0_u11_u5_n137 ) , .A( u0_u11_u5_n146 ) , .B2( u0_u11_u5_n147 ) );
  NOR2_X1 u0_u11_u5_U77 (.A2( u0_u11_X_34 ) , .A1( u0_u11_X_35 ) , .ZN( u0_u11_u5_n145 ) );
  NOR2_X1 u0_u11_u5_U78 (.A2( u0_u11_X_34 ) , .ZN( u0_u11_u5_n146 ) , .A1( u0_u11_u5_n171 ) );
  NOR2_X1 u0_u11_u5_U79 (.A2( u0_u11_X_31 ) , .A1( u0_u11_X_32 ) , .ZN( u0_u11_u5_n103 ) );
  NOR3_X1 u0_u11_u5_U8 (.A2( u0_u11_u5_n147 ) , .A1( u0_u11_u5_n148 ) , .ZN( u0_u11_u5_n149 ) , .A3( u0_u11_u5_n194 ) );
  NOR2_X1 u0_u11_u5_U80 (.A2( u0_u11_X_36 ) , .ZN( u0_u11_u5_n105 ) , .A1( u0_u11_u5_n180 ) );
  NOR2_X1 u0_u11_u5_U81 (.A2( u0_u11_X_33 ) , .ZN( u0_u11_u5_n108 ) , .A1( u0_u11_u5_n170 ) );
  NOR2_X1 u0_u11_u5_U82 (.A2( u0_u11_X_33 ) , .A1( u0_u11_X_36 ) , .ZN( u0_u11_u5_n107 ) );
  NOR2_X1 u0_u11_u5_U83 (.A2( u0_u11_X_31 ) , .ZN( u0_u11_u5_n104 ) , .A1( u0_u11_u5_n181 ) );
  NAND2_X1 u0_u11_u5_U84 (.A2( u0_u11_X_34 ) , .A1( u0_u11_X_35 ) , .ZN( u0_u11_u5_n153 ) );
  NAND2_X1 u0_u11_u5_U85 (.A1( u0_u11_X_34 ) , .ZN( u0_u11_u5_n126 ) , .A2( u0_u11_u5_n171 ) );
  AND2_X1 u0_u11_u5_U86 (.A1( u0_u11_X_31 ) , .A2( u0_u11_X_32 ) , .ZN( u0_u11_u5_n106 ) );
  AND2_X1 u0_u11_u5_U87 (.A1( u0_u11_X_31 ) , .ZN( u0_u11_u5_n109 ) , .A2( u0_u11_u5_n181 ) );
  INV_X1 u0_u11_u5_U88 (.A( u0_u11_X_33 ) , .ZN( u0_u11_u5_n180 ) );
  INV_X1 u0_u11_u5_U89 (.A( u0_u11_X_35 ) , .ZN( u0_u11_u5_n171 ) );
  NOR2_X1 u0_u11_u5_U9 (.ZN( u0_u11_u5_n135 ) , .A1( u0_u11_u5_n173 ) , .A2( u0_u11_u5_n176 ) );
  INV_X1 u0_u11_u5_U90 (.A( u0_u11_X_36 ) , .ZN( u0_u11_u5_n170 ) );
  INV_X1 u0_u11_u5_U91 (.A( u0_u11_X_32 ) , .ZN( u0_u11_u5_n181 ) );
  NAND4_X1 u0_u11_u5_U92 (.ZN( u0_out11_29 ) , .A4( u0_u11_u5_n129 ) , .A3( u0_u11_u5_n130 ) , .A2( u0_u11_u5_n168 ) , .A1( u0_u11_u5_n196 ) );
  AOI221_X1 u0_u11_u5_U93 (.A( u0_u11_u5_n128 ) , .ZN( u0_u11_u5_n129 ) , .C2( u0_u11_u5_n132 ) , .B2( u0_u11_u5_n159 ) , .B1( u0_u11_u5_n176 ) , .C1( u0_u11_u5_n184 ) );
  AOI222_X1 u0_u11_u5_U94 (.ZN( u0_u11_u5_n130 ) , .A2( u0_u11_u5_n146 ) , .B1( u0_u11_u5_n147 ) , .C2( u0_u11_u5_n175 ) , .B2( u0_u11_u5_n179 ) , .A1( u0_u11_u5_n188 ) , .C1( u0_u11_u5_n194 ) );
  NAND4_X1 u0_u11_u5_U95 (.ZN( u0_out11_19 ) , .A4( u0_u11_u5_n166 ) , .A3( u0_u11_u5_n167 ) , .A2( u0_u11_u5_n168 ) , .A1( u0_u11_u5_n169 ) );
  AOI22_X1 u0_u11_u5_U96 (.B2( u0_u11_u5_n145 ) , .A2( u0_u11_u5_n146 ) , .ZN( u0_u11_u5_n167 ) , .B1( u0_u11_u5_n182 ) , .A1( u0_u11_u5_n189 ) );
  NOR4_X1 u0_u11_u5_U97 (.A4( u0_u11_u5_n162 ) , .A3( u0_u11_u5_n163 ) , .A2( u0_u11_u5_n164 ) , .A1( u0_u11_u5_n165 ) , .ZN( u0_u11_u5_n166 ) );
  NAND4_X1 u0_u11_u5_U98 (.ZN( u0_out11_11 ) , .A4( u0_u11_u5_n143 ) , .A3( u0_u11_u5_n144 ) , .A2( u0_u11_u5_n169 ) , .A1( u0_u11_u5_n196 ) );
  AOI22_X1 u0_u11_u5_U99 (.A2( u0_u11_u5_n132 ) , .ZN( u0_u11_u5_n144 ) , .B2( u0_u11_u5_n145 ) , .B1( u0_u11_u5_n184 ) , .A1( u0_u11_u5_n194 ) );
  XOR2_X1 u0_u1_U33 (.B( u0_K2_24 ) , .A( u0_R0_17 ) , .Z( u0_u1_X_24 ) );
  XOR2_X1 u0_u1_U34 (.B( u0_K2_23 ) , .A( u0_R0_16 ) , .Z( u0_u1_X_23 ) );
  XOR2_X1 u0_u1_U35 (.B( u0_K2_22 ) , .A( u0_R0_15 ) , .Z( u0_u1_X_22 ) );
  XOR2_X1 u0_u1_U36 (.B( u0_K2_21 ) , .A( u0_R0_14 ) , .Z( u0_u1_X_21 ) );
  XOR2_X1 u0_u1_U37 (.B( u0_K2_20 ) , .A( u0_R0_13 ) , .Z( u0_u1_X_20 ) );
  XOR2_X1 u0_u1_U39 (.B( u0_K2_19 ) , .A( u0_R0_12 ) , .Z( u0_u1_X_19 ) );
  OAI22_X1 u0_u1_u3_U10 (.B1( u0_u1_u3_n113 ) , .A2( u0_u1_u3_n135 ) , .A1( u0_u1_u3_n150 ) , .B2( u0_u1_u3_n164 ) , .ZN( u0_u1_u3_n98 ) );
  OAI211_X1 u0_u1_u3_U11 (.B( u0_u1_u3_n106 ) , .ZN( u0_u1_u3_n119 ) , .C2( u0_u1_u3_n128 ) , .C1( u0_u1_u3_n167 ) , .A( u0_u1_u3_n181 ) );
  AOI221_X1 u0_u1_u3_U12 (.C1( u0_u1_u3_n105 ) , .ZN( u0_u1_u3_n106 ) , .A( u0_u1_u3_n131 ) , .B2( u0_u1_u3_n132 ) , .C2( u0_u1_u3_n133 ) , .B1( u0_u1_u3_n169 ) );
  INV_X1 u0_u1_u3_U13 (.ZN( u0_u1_u3_n181 ) , .A( u0_u1_u3_n98 ) );
  NAND2_X1 u0_u1_u3_U14 (.ZN( u0_u1_u3_n105 ) , .A2( u0_u1_u3_n130 ) , .A1( u0_u1_u3_n155 ) );
  AOI22_X1 u0_u1_u3_U15 (.B1( u0_u1_u3_n115 ) , .A2( u0_u1_u3_n116 ) , .ZN( u0_u1_u3_n123 ) , .B2( u0_u1_u3_n133 ) , .A1( u0_u1_u3_n169 ) );
  NAND2_X1 u0_u1_u3_U16 (.ZN( u0_u1_u3_n116 ) , .A2( u0_u1_u3_n151 ) , .A1( u0_u1_u3_n182 ) );
  NOR2_X1 u0_u1_u3_U17 (.ZN( u0_u1_u3_n126 ) , .A2( u0_u1_u3_n150 ) , .A1( u0_u1_u3_n164 ) );
  AOI21_X1 u0_u1_u3_U18 (.ZN( u0_u1_u3_n112 ) , .B2( u0_u1_u3_n146 ) , .B1( u0_u1_u3_n155 ) , .A( u0_u1_u3_n167 ) );
  NAND2_X1 u0_u1_u3_U19 (.A1( u0_u1_u3_n135 ) , .ZN( u0_u1_u3_n142 ) , .A2( u0_u1_u3_n164 ) );
  NAND2_X1 u0_u1_u3_U20 (.ZN( u0_u1_u3_n132 ) , .A2( u0_u1_u3_n152 ) , .A1( u0_u1_u3_n156 ) );
  AND2_X1 u0_u1_u3_U21 (.A2( u0_u1_u3_n113 ) , .A1( u0_u1_u3_n114 ) , .ZN( u0_u1_u3_n151 ) );
  INV_X1 u0_u1_u3_U22 (.A( u0_u1_u3_n133 ) , .ZN( u0_u1_u3_n165 ) );
  INV_X1 u0_u1_u3_U23 (.A( u0_u1_u3_n135 ) , .ZN( u0_u1_u3_n170 ) );
  NAND2_X1 u0_u1_u3_U24 (.A1( u0_u1_u3_n107 ) , .A2( u0_u1_u3_n108 ) , .ZN( u0_u1_u3_n140 ) );
  NAND2_X1 u0_u1_u3_U25 (.ZN( u0_u1_u3_n117 ) , .A1( u0_u1_u3_n124 ) , .A2( u0_u1_u3_n148 ) );
  NAND2_X1 u0_u1_u3_U26 (.ZN( u0_u1_u3_n143 ) , .A1( u0_u1_u3_n165 ) , .A2( u0_u1_u3_n167 ) );
  INV_X1 u0_u1_u3_U27 (.A( u0_u1_u3_n130 ) , .ZN( u0_u1_u3_n177 ) );
  INV_X1 u0_u1_u3_U28 (.A( u0_u1_u3_n128 ) , .ZN( u0_u1_u3_n176 ) );
  INV_X1 u0_u1_u3_U29 (.A( u0_u1_u3_n155 ) , .ZN( u0_u1_u3_n174 ) );
  INV_X1 u0_u1_u3_U3 (.A( u0_u1_u3_n129 ) , .ZN( u0_u1_u3_n183 ) );
  INV_X1 u0_u1_u3_U30 (.A( u0_u1_u3_n139 ) , .ZN( u0_u1_u3_n185 ) );
  NOR2_X1 u0_u1_u3_U31 (.ZN( u0_u1_u3_n135 ) , .A2( u0_u1_u3_n141 ) , .A1( u0_u1_u3_n169 ) );
  OAI222_X1 u0_u1_u3_U32 (.C2( u0_u1_u3_n107 ) , .A2( u0_u1_u3_n108 ) , .B1( u0_u1_u3_n135 ) , .ZN( u0_u1_u3_n138 ) , .B2( u0_u1_u3_n146 ) , .C1( u0_u1_u3_n154 ) , .A1( u0_u1_u3_n164 ) );
  NOR4_X1 u0_u1_u3_U33 (.A4( u0_u1_u3_n157 ) , .A3( u0_u1_u3_n158 ) , .A2( u0_u1_u3_n159 ) , .A1( u0_u1_u3_n160 ) , .ZN( u0_u1_u3_n161 ) );
  AOI21_X1 u0_u1_u3_U34 (.B2( u0_u1_u3_n152 ) , .B1( u0_u1_u3_n153 ) , .ZN( u0_u1_u3_n158 ) , .A( u0_u1_u3_n164 ) );
  AOI21_X1 u0_u1_u3_U35 (.A( u0_u1_u3_n154 ) , .B2( u0_u1_u3_n155 ) , .B1( u0_u1_u3_n156 ) , .ZN( u0_u1_u3_n157 ) );
  AOI21_X1 u0_u1_u3_U36 (.A( u0_u1_u3_n149 ) , .B2( u0_u1_u3_n150 ) , .B1( u0_u1_u3_n151 ) , .ZN( u0_u1_u3_n159 ) );
  AOI211_X1 u0_u1_u3_U37 (.ZN( u0_u1_u3_n109 ) , .A( u0_u1_u3_n119 ) , .C2( u0_u1_u3_n129 ) , .B( u0_u1_u3_n138 ) , .C1( u0_u1_u3_n141 ) );
  AOI211_X1 u0_u1_u3_U38 (.B( u0_u1_u3_n119 ) , .A( u0_u1_u3_n120 ) , .C2( u0_u1_u3_n121 ) , .ZN( u0_u1_u3_n122 ) , .C1( u0_u1_u3_n179 ) );
  INV_X1 u0_u1_u3_U39 (.A( u0_u1_u3_n156 ) , .ZN( u0_u1_u3_n179 ) );
  INV_X1 u0_u1_u3_U4 (.A( u0_u1_u3_n140 ) , .ZN( u0_u1_u3_n182 ) );
  OAI22_X1 u0_u1_u3_U40 (.B1( u0_u1_u3_n118 ) , .ZN( u0_u1_u3_n120 ) , .A1( u0_u1_u3_n135 ) , .B2( u0_u1_u3_n154 ) , .A2( u0_u1_u3_n178 ) );
  AND3_X1 u0_u1_u3_U41 (.ZN( u0_u1_u3_n118 ) , .A2( u0_u1_u3_n124 ) , .A1( u0_u1_u3_n144 ) , .A3( u0_u1_u3_n152 ) );
  INV_X1 u0_u1_u3_U42 (.A( u0_u1_u3_n121 ) , .ZN( u0_u1_u3_n164 ) );
  NAND2_X1 u0_u1_u3_U43 (.ZN( u0_u1_u3_n133 ) , .A1( u0_u1_u3_n154 ) , .A2( u0_u1_u3_n164 ) );
  OAI211_X1 u0_u1_u3_U44 (.B( u0_u1_u3_n127 ) , .ZN( u0_u1_u3_n139 ) , .C1( u0_u1_u3_n150 ) , .C2( u0_u1_u3_n154 ) , .A( u0_u1_u3_n184 ) );
  INV_X1 u0_u1_u3_U45 (.A( u0_u1_u3_n125 ) , .ZN( u0_u1_u3_n184 ) );
  AOI221_X1 u0_u1_u3_U46 (.A( u0_u1_u3_n126 ) , .ZN( u0_u1_u3_n127 ) , .C2( u0_u1_u3_n132 ) , .C1( u0_u1_u3_n169 ) , .B2( u0_u1_u3_n170 ) , .B1( u0_u1_u3_n174 ) );
  OAI22_X1 u0_u1_u3_U47 (.A1( u0_u1_u3_n124 ) , .ZN( u0_u1_u3_n125 ) , .B2( u0_u1_u3_n145 ) , .A2( u0_u1_u3_n165 ) , .B1( u0_u1_u3_n167 ) );
  NOR2_X1 u0_u1_u3_U48 (.A1( u0_u1_u3_n113 ) , .ZN( u0_u1_u3_n131 ) , .A2( u0_u1_u3_n154 ) );
  NAND2_X1 u0_u1_u3_U49 (.A1( u0_u1_u3_n103 ) , .ZN( u0_u1_u3_n150 ) , .A2( u0_u1_u3_n99 ) );
  INV_X1 u0_u1_u3_U5 (.A( u0_u1_u3_n117 ) , .ZN( u0_u1_u3_n178 ) );
  NAND2_X1 u0_u1_u3_U50 (.A2( u0_u1_u3_n102 ) , .ZN( u0_u1_u3_n155 ) , .A1( u0_u1_u3_n97 ) );
  INV_X1 u0_u1_u3_U51 (.A( u0_u1_u3_n141 ) , .ZN( u0_u1_u3_n167 ) );
  AOI21_X1 u0_u1_u3_U52 (.B2( u0_u1_u3_n114 ) , .B1( u0_u1_u3_n146 ) , .A( u0_u1_u3_n154 ) , .ZN( u0_u1_u3_n94 ) );
  AOI21_X1 u0_u1_u3_U53 (.ZN( u0_u1_u3_n110 ) , .B2( u0_u1_u3_n142 ) , .B1( u0_u1_u3_n186 ) , .A( u0_u1_u3_n95 ) );
  INV_X1 u0_u1_u3_U54 (.A( u0_u1_u3_n145 ) , .ZN( u0_u1_u3_n186 ) );
  AOI21_X1 u0_u1_u3_U55 (.B1( u0_u1_u3_n124 ) , .A( u0_u1_u3_n149 ) , .B2( u0_u1_u3_n155 ) , .ZN( u0_u1_u3_n95 ) );
  INV_X1 u0_u1_u3_U56 (.A( u0_u1_u3_n149 ) , .ZN( u0_u1_u3_n169 ) );
  NAND2_X1 u0_u1_u3_U57 (.ZN( u0_u1_u3_n124 ) , .A1( u0_u1_u3_n96 ) , .A2( u0_u1_u3_n97 ) );
  NAND2_X1 u0_u1_u3_U58 (.A2( u0_u1_u3_n100 ) , .ZN( u0_u1_u3_n146 ) , .A1( u0_u1_u3_n96 ) );
  NAND2_X1 u0_u1_u3_U59 (.A1( u0_u1_u3_n101 ) , .ZN( u0_u1_u3_n145 ) , .A2( u0_u1_u3_n99 ) );
  AOI221_X1 u0_u1_u3_U6 (.A( u0_u1_u3_n131 ) , .C2( u0_u1_u3_n132 ) , .C1( u0_u1_u3_n133 ) , .ZN( u0_u1_u3_n134 ) , .B1( u0_u1_u3_n143 ) , .B2( u0_u1_u3_n177 ) );
  NAND2_X1 u0_u1_u3_U60 (.A1( u0_u1_u3_n100 ) , .ZN( u0_u1_u3_n156 ) , .A2( u0_u1_u3_n99 ) );
  NAND2_X1 u0_u1_u3_U61 (.A2( u0_u1_u3_n101 ) , .A1( u0_u1_u3_n104 ) , .ZN( u0_u1_u3_n148 ) );
  NAND2_X1 u0_u1_u3_U62 (.A1( u0_u1_u3_n100 ) , .A2( u0_u1_u3_n102 ) , .ZN( u0_u1_u3_n128 ) );
  NAND2_X1 u0_u1_u3_U63 (.A2( u0_u1_u3_n101 ) , .A1( u0_u1_u3_n102 ) , .ZN( u0_u1_u3_n152 ) );
  NAND2_X1 u0_u1_u3_U64 (.A2( u0_u1_u3_n101 ) , .ZN( u0_u1_u3_n114 ) , .A1( u0_u1_u3_n96 ) );
  NAND2_X1 u0_u1_u3_U65 (.ZN( u0_u1_u3_n107 ) , .A1( u0_u1_u3_n97 ) , .A2( u0_u1_u3_n99 ) );
  NAND2_X1 u0_u1_u3_U66 (.A2( u0_u1_u3_n100 ) , .A1( u0_u1_u3_n104 ) , .ZN( u0_u1_u3_n113 ) );
  NAND2_X1 u0_u1_u3_U67 (.A1( u0_u1_u3_n104 ) , .ZN( u0_u1_u3_n153 ) , .A2( u0_u1_u3_n97 ) );
  NAND2_X1 u0_u1_u3_U68 (.A2( u0_u1_u3_n103 ) , .A1( u0_u1_u3_n104 ) , .ZN( u0_u1_u3_n130 ) );
  NAND2_X1 u0_u1_u3_U69 (.A2( u0_u1_u3_n103 ) , .ZN( u0_u1_u3_n144 ) , .A1( u0_u1_u3_n96 ) );
  OAI22_X1 u0_u1_u3_U7 (.B2( u0_u1_u3_n147 ) , .A2( u0_u1_u3_n148 ) , .ZN( u0_u1_u3_n160 ) , .B1( u0_u1_u3_n165 ) , .A1( u0_u1_u3_n168 ) );
  NAND2_X1 u0_u1_u3_U70 (.A1( u0_u1_u3_n102 ) , .A2( u0_u1_u3_n103 ) , .ZN( u0_u1_u3_n108 ) );
  NOR2_X1 u0_u1_u3_U71 (.A2( u0_u1_X_19 ) , .A1( u0_u1_X_20 ) , .ZN( u0_u1_u3_n99 ) );
  NOR2_X1 u0_u1_u3_U72 (.A2( u0_u1_X_21 ) , .A1( u0_u1_X_24 ) , .ZN( u0_u1_u3_n103 ) );
  NOR2_X1 u0_u1_u3_U73 (.A2( u0_u1_X_24 ) , .A1( u0_u1_u3_n171 ) , .ZN( u0_u1_u3_n97 ) );
  NOR2_X1 u0_u1_u3_U74 (.A2( u0_u1_X_23 ) , .ZN( u0_u1_u3_n141 ) , .A1( u0_u1_u3_n166 ) );
  NOR2_X1 u0_u1_u3_U75 (.A2( u0_u1_X_19 ) , .A1( u0_u1_u3_n172 ) , .ZN( u0_u1_u3_n96 ) );
  NAND2_X1 u0_u1_u3_U76 (.A1( u0_u1_X_22 ) , .A2( u0_u1_X_23 ) , .ZN( u0_u1_u3_n154 ) );
  NAND2_X1 u0_u1_u3_U77 (.A1( u0_u1_X_23 ) , .ZN( u0_u1_u3_n149 ) , .A2( u0_u1_u3_n166 ) );
  NOR2_X1 u0_u1_u3_U78 (.A2( u0_u1_X_22 ) , .A1( u0_u1_X_23 ) , .ZN( u0_u1_u3_n121 ) );
  AND2_X1 u0_u1_u3_U79 (.A1( u0_u1_X_24 ) , .ZN( u0_u1_u3_n101 ) , .A2( u0_u1_u3_n171 ) );
  AND3_X1 u0_u1_u3_U8 (.A3( u0_u1_u3_n144 ) , .A2( u0_u1_u3_n145 ) , .A1( u0_u1_u3_n146 ) , .ZN( u0_u1_u3_n147 ) );
  AND2_X1 u0_u1_u3_U80 (.A1( u0_u1_X_19 ) , .ZN( u0_u1_u3_n102 ) , .A2( u0_u1_u3_n172 ) );
  AND2_X1 u0_u1_u3_U81 (.A1( u0_u1_X_21 ) , .A2( u0_u1_X_24 ) , .ZN( u0_u1_u3_n100 ) );
  AND2_X1 u0_u1_u3_U82 (.A2( u0_u1_X_19 ) , .A1( u0_u1_X_20 ) , .ZN( u0_u1_u3_n104 ) );
  INV_X1 u0_u1_u3_U83 (.A( u0_u1_X_22 ) , .ZN( u0_u1_u3_n166 ) );
  INV_X1 u0_u1_u3_U84 (.A( u0_u1_X_21 ) , .ZN( u0_u1_u3_n171 ) );
  INV_X1 u0_u1_u3_U85 (.A( u0_u1_X_20 ) , .ZN( u0_u1_u3_n172 ) );
  OR4_X1 u0_u1_u3_U86 (.ZN( u0_out1_10 ) , .A4( u0_u1_u3_n136 ) , .A3( u0_u1_u3_n137 ) , .A1( u0_u1_u3_n138 ) , .A2( u0_u1_u3_n139 ) );
  OAI222_X1 u0_u1_u3_U87 (.C1( u0_u1_u3_n128 ) , .ZN( u0_u1_u3_n137 ) , .B1( u0_u1_u3_n148 ) , .A2( u0_u1_u3_n150 ) , .B2( u0_u1_u3_n154 ) , .C2( u0_u1_u3_n164 ) , .A1( u0_u1_u3_n167 ) );
  OAI221_X1 u0_u1_u3_U88 (.A( u0_u1_u3_n134 ) , .B2( u0_u1_u3_n135 ) , .ZN( u0_u1_u3_n136 ) , .C1( u0_u1_u3_n149 ) , .B1( u0_u1_u3_n151 ) , .C2( u0_u1_u3_n183 ) );
  NAND4_X1 u0_u1_u3_U89 (.ZN( u0_out1_26 ) , .A4( u0_u1_u3_n109 ) , .A3( u0_u1_u3_n110 ) , .A2( u0_u1_u3_n111 ) , .A1( u0_u1_u3_n173 ) );
  INV_X1 u0_u1_u3_U9 (.A( u0_u1_u3_n143 ) , .ZN( u0_u1_u3_n168 ) );
  INV_X1 u0_u1_u3_U90 (.ZN( u0_u1_u3_n173 ) , .A( u0_u1_u3_n94 ) );
  OAI21_X1 u0_u1_u3_U91 (.ZN( u0_u1_u3_n111 ) , .B2( u0_u1_u3_n117 ) , .A( u0_u1_u3_n133 ) , .B1( u0_u1_u3_n176 ) );
  NAND4_X1 u0_u1_u3_U92 (.ZN( u0_out1_20 ) , .A4( u0_u1_u3_n122 ) , .A3( u0_u1_u3_n123 ) , .A1( u0_u1_u3_n175 ) , .A2( u0_u1_u3_n180 ) );
  INV_X1 u0_u1_u3_U93 (.A( u0_u1_u3_n112 ) , .ZN( u0_u1_u3_n175 ) );
  INV_X1 u0_u1_u3_U94 (.A( u0_u1_u3_n126 ) , .ZN( u0_u1_u3_n180 ) );
  NAND4_X1 u0_u1_u3_U95 (.ZN( u0_out1_1 ) , .A4( u0_u1_u3_n161 ) , .A3( u0_u1_u3_n162 ) , .A2( u0_u1_u3_n163 ) , .A1( u0_u1_u3_n185 ) );
  NAND2_X1 u0_u1_u3_U96 (.ZN( u0_u1_u3_n163 ) , .A2( u0_u1_u3_n170 ) , .A1( u0_u1_u3_n176 ) );
  AOI22_X1 u0_u1_u3_U97 (.B2( u0_u1_u3_n140 ) , .B1( u0_u1_u3_n141 ) , .A2( u0_u1_u3_n142 ) , .ZN( u0_u1_u3_n162 ) , .A1( u0_u1_u3_n177 ) );
  NAND3_X1 u0_u1_u3_U98 (.A1( u0_u1_u3_n114 ) , .ZN( u0_u1_u3_n115 ) , .A2( u0_u1_u3_n145 ) , .A3( u0_u1_u3_n153 ) );
  NAND3_X1 u0_u1_u3_U99 (.ZN( u0_u1_u3_n129 ) , .A2( u0_u1_u3_n144 ) , .A1( u0_u1_u3_n153 ) , .A3( u0_u1_u3_n182 ) );
  XOR2_X1 u0_u2_U26 (.B( u0_K3_30 ) , .A( u0_R1_21 ) , .Z( u0_u2_X_30 ) );
  XOR2_X1 u0_u2_U28 (.B( u0_K3_29 ) , .A( u0_R1_20 ) , .Z( u0_u2_X_29 ) );
  XOR2_X1 u0_u2_U29 (.B( u0_K3_28 ) , .A( u0_R1_19 ) , .Z( u0_u2_X_28 ) );
  XOR2_X1 u0_u2_U30 (.B( u0_K3_27 ) , .A( u0_R1_18 ) , .Z( u0_u2_X_27 ) );
  XOR2_X1 u0_u2_U31 (.B( u0_K3_26 ) , .A( u0_R1_17 ) , .Z( u0_u2_X_26 ) );
  XOR2_X1 u0_u2_U32 (.B( u0_K3_25 ) , .A( u0_R1_16 ) , .Z( u0_u2_X_25 ) );
  OAI22_X1 u0_u2_u4_U10 (.B2( u0_u2_u4_n135 ) , .ZN( u0_u2_u4_n137 ) , .B1( u0_u2_u4_n153 ) , .A1( u0_u2_u4_n155 ) , .A2( u0_u2_u4_n171 ) );
  AND3_X1 u0_u2_u4_U11 (.A2( u0_u2_u4_n134 ) , .ZN( u0_u2_u4_n135 ) , .A3( u0_u2_u4_n145 ) , .A1( u0_u2_u4_n157 ) );
  NAND2_X1 u0_u2_u4_U12 (.ZN( u0_u2_u4_n132 ) , .A2( u0_u2_u4_n170 ) , .A1( u0_u2_u4_n173 ) );
  AOI21_X1 u0_u2_u4_U13 (.B2( u0_u2_u4_n160 ) , .B1( u0_u2_u4_n161 ) , .ZN( u0_u2_u4_n162 ) , .A( u0_u2_u4_n170 ) );
  AOI21_X1 u0_u2_u4_U14 (.ZN( u0_u2_u4_n107 ) , .B2( u0_u2_u4_n143 ) , .A( u0_u2_u4_n174 ) , .B1( u0_u2_u4_n184 ) );
  AOI21_X1 u0_u2_u4_U15 (.B2( u0_u2_u4_n158 ) , .B1( u0_u2_u4_n159 ) , .ZN( u0_u2_u4_n163 ) , .A( u0_u2_u4_n174 ) );
  AOI21_X1 u0_u2_u4_U16 (.A( u0_u2_u4_n153 ) , .B2( u0_u2_u4_n154 ) , .B1( u0_u2_u4_n155 ) , .ZN( u0_u2_u4_n165 ) );
  AOI21_X1 u0_u2_u4_U17 (.A( u0_u2_u4_n156 ) , .B2( u0_u2_u4_n157 ) , .ZN( u0_u2_u4_n164 ) , .B1( u0_u2_u4_n184 ) );
  INV_X1 u0_u2_u4_U18 (.A( u0_u2_u4_n138 ) , .ZN( u0_u2_u4_n170 ) );
  AND2_X1 u0_u2_u4_U19 (.A2( u0_u2_u4_n120 ) , .ZN( u0_u2_u4_n155 ) , .A1( u0_u2_u4_n160 ) );
  INV_X1 u0_u2_u4_U20 (.A( u0_u2_u4_n156 ) , .ZN( u0_u2_u4_n175 ) );
  NAND2_X1 u0_u2_u4_U21 (.A2( u0_u2_u4_n118 ) , .ZN( u0_u2_u4_n131 ) , .A1( u0_u2_u4_n147 ) );
  NAND2_X1 u0_u2_u4_U22 (.A1( u0_u2_u4_n119 ) , .A2( u0_u2_u4_n120 ) , .ZN( u0_u2_u4_n130 ) );
  NAND2_X1 u0_u2_u4_U23 (.ZN( u0_u2_u4_n117 ) , .A2( u0_u2_u4_n118 ) , .A1( u0_u2_u4_n148 ) );
  NAND2_X1 u0_u2_u4_U24 (.ZN( u0_u2_u4_n129 ) , .A1( u0_u2_u4_n134 ) , .A2( u0_u2_u4_n148 ) );
  AND3_X1 u0_u2_u4_U25 (.A1( u0_u2_u4_n119 ) , .A2( u0_u2_u4_n143 ) , .A3( u0_u2_u4_n154 ) , .ZN( u0_u2_u4_n161 ) );
  AND2_X1 u0_u2_u4_U26 (.A1( u0_u2_u4_n145 ) , .A2( u0_u2_u4_n147 ) , .ZN( u0_u2_u4_n159 ) );
  OR3_X1 u0_u2_u4_U27 (.A3( u0_u2_u4_n114 ) , .A2( u0_u2_u4_n115 ) , .A1( u0_u2_u4_n116 ) , .ZN( u0_u2_u4_n136 ) );
  AOI21_X1 u0_u2_u4_U28 (.A( u0_u2_u4_n113 ) , .ZN( u0_u2_u4_n116 ) , .B2( u0_u2_u4_n173 ) , .B1( u0_u2_u4_n174 ) );
  AOI21_X1 u0_u2_u4_U29 (.ZN( u0_u2_u4_n115 ) , .B2( u0_u2_u4_n145 ) , .B1( u0_u2_u4_n146 ) , .A( u0_u2_u4_n156 ) );
  NOR2_X1 u0_u2_u4_U3 (.ZN( u0_u2_u4_n121 ) , .A1( u0_u2_u4_n181 ) , .A2( u0_u2_u4_n182 ) );
  OAI22_X1 u0_u2_u4_U30 (.ZN( u0_u2_u4_n114 ) , .A2( u0_u2_u4_n121 ) , .B1( u0_u2_u4_n160 ) , .B2( u0_u2_u4_n170 ) , .A1( u0_u2_u4_n171 ) );
  INV_X1 u0_u2_u4_U31 (.A( u0_u2_u4_n158 ) , .ZN( u0_u2_u4_n182 ) );
  INV_X1 u0_u2_u4_U32 (.ZN( u0_u2_u4_n181 ) , .A( u0_u2_u4_n96 ) );
  INV_X1 u0_u2_u4_U33 (.A( u0_u2_u4_n144 ) , .ZN( u0_u2_u4_n179 ) );
  INV_X1 u0_u2_u4_U34 (.A( u0_u2_u4_n157 ) , .ZN( u0_u2_u4_n178 ) );
  NAND2_X1 u0_u2_u4_U35 (.A2( u0_u2_u4_n154 ) , .A1( u0_u2_u4_n96 ) , .ZN( u0_u2_u4_n97 ) );
  INV_X1 u0_u2_u4_U36 (.ZN( u0_u2_u4_n186 ) , .A( u0_u2_u4_n95 ) );
  OAI221_X1 u0_u2_u4_U37 (.C1( u0_u2_u4_n134 ) , .B1( u0_u2_u4_n158 ) , .B2( u0_u2_u4_n171 ) , .C2( u0_u2_u4_n173 ) , .A( u0_u2_u4_n94 ) , .ZN( u0_u2_u4_n95 ) );
  AOI222_X1 u0_u2_u4_U38 (.B2( u0_u2_u4_n132 ) , .A1( u0_u2_u4_n138 ) , .C2( u0_u2_u4_n175 ) , .A2( u0_u2_u4_n179 ) , .C1( u0_u2_u4_n181 ) , .B1( u0_u2_u4_n185 ) , .ZN( u0_u2_u4_n94 ) );
  INV_X1 u0_u2_u4_U39 (.A( u0_u2_u4_n113 ) , .ZN( u0_u2_u4_n185 ) );
  INV_X1 u0_u2_u4_U4 (.A( u0_u2_u4_n117 ) , .ZN( u0_u2_u4_n184 ) );
  INV_X1 u0_u2_u4_U40 (.A( u0_u2_u4_n143 ) , .ZN( u0_u2_u4_n183 ) );
  NOR2_X1 u0_u2_u4_U41 (.ZN( u0_u2_u4_n138 ) , .A1( u0_u2_u4_n168 ) , .A2( u0_u2_u4_n169 ) );
  NOR2_X1 u0_u2_u4_U42 (.A1( u0_u2_u4_n150 ) , .A2( u0_u2_u4_n152 ) , .ZN( u0_u2_u4_n153 ) );
  NOR2_X1 u0_u2_u4_U43 (.A2( u0_u2_u4_n128 ) , .A1( u0_u2_u4_n138 ) , .ZN( u0_u2_u4_n156 ) );
  AOI22_X1 u0_u2_u4_U44 (.B2( u0_u2_u4_n122 ) , .A1( u0_u2_u4_n123 ) , .ZN( u0_u2_u4_n124 ) , .B1( u0_u2_u4_n128 ) , .A2( u0_u2_u4_n172 ) );
  INV_X1 u0_u2_u4_U45 (.A( u0_u2_u4_n153 ) , .ZN( u0_u2_u4_n172 ) );
  NAND2_X1 u0_u2_u4_U46 (.A2( u0_u2_u4_n120 ) , .ZN( u0_u2_u4_n123 ) , .A1( u0_u2_u4_n161 ) );
  AOI22_X1 u0_u2_u4_U47 (.B2( u0_u2_u4_n132 ) , .A2( u0_u2_u4_n133 ) , .ZN( u0_u2_u4_n140 ) , .A1( u0_u2_u4_n150 ) , .B1( u0_u2_u4_n179 ) );
  NAND2_X1 u0_u2_u4_U48 (.ZN( u0_u2_u4_n133 ) , .A2( u0_u2_u4_n146 ) , .A1( u0_u2_u4_n154 ) );
  NAND2_X1 u0_u2_u4_U49 (.A1( u0_u2_u4_n103 ) , .ZN( u0_u2_u4_n154 ) , .A2( u0_u2_u4_n98 ) );
  NOR4_X1 u0_u2_u4_U5 (.A4( u0_u2_u4_n106 ) , .A3( u0_u2_u4_n107 ) , .A2( u0_u2_u4_n108 ) , .A1( u0_u2_u4_n109 ) , .ZN( u0_u2_u4_n110 ) );
  NAND2_X1 u0_u2_u4_U50 (.A1( u0_u2_u4_n101 ) , .ZN( u0_u2_u4_n158 ) , .A2( u0_u2_u4_n99 ) );
  AOI21_X1 u0_u2_u4_U51 (.ZN( u0_u2_u4_n127 ) , .A( u0_u2_u4_n136 ) , .B2( u0_u2_u4_n150 ) , .B1( u0_u2_u4_n180 ) );
  INV_X1 u0_u2_u4_U52 (.A( u0_u2_u4_n160 ) , .ZN( u0_u2_u4_n180 ) );
  NAND2_X1 u0_u2_u4_U53 (.A2( u0_u2_u4_n104 ) , .A1( u0_u2_u4_n105 ) , .ZN( u0_u2_u4_n146 ) );
  NAND2_X1 u0_u2_u4_U54 (.A2( u0_u2_u4_n101 ) , .A1( u0_u2_u4_n102 ) , .ZN( u0_u2_u4_n160 ) );
  NAND2_X1 u0_u2_u4_U55 (.ZN( u0_u2_u4_n134 ) , .A1( u0_u2_u4_n98 ) , .A2( u0_u2_u4_n99 ) );
  NAND2_X1 u0_u2_u4_U56 (.A1( u0_u2_u4_n103 ) , .A2( u0_u2_u4_n104 ) , .ZN( u0_u2_u4_n143 ) );
  NAND2_X1 u0_u2_u4_U57 (.A2( u0_u2_u4_n105 ) , .ZN( u0_u2_u4_n145 ) , .A1( u0_u2_u4_n98 ) );
  NAND2_X1 u0_u2_u4_U58 (.A1( u0_u2_u4_n100 ) , .A2( u0_u2_u4_n105 ) , .ZN( u0_u2_u4_n120 ) );
  NAND2_X1 u0_u2_u4_U59 (.A1( u0_u2_u4_n102 ) , .A2( u0_u2_u4_n104 ) , .ZN( u0_u2_u4_n148 ) );
  AOI21_X1 u0_u2_u4_U6 (.ZN( u0_u2_u4_n106 ) , .B2( u0_u2_u4_n146 ) , .B1( u0_u2_u4_n158 ) , .A( u0_u2_u4_n170 ) );
  NAND2_X1 u0_u2_u4_U60 (.A2( u0_u2_u4_n100 ) , .A1( u0_u2_u4_n103 ) , .ZN( u0_u2_u4_n157 ) );
  INV_X1 u0_u2_u4_U61 (.A( u0_u2_u4_n150 ) , .ZN( u0_u2_u4_n173 ) );
  INV_X1 u0_u2_u4_U62 (.A( u0_u2_u4_n152 ) , .ZN( u0_u2_u4_n171 ) );
  NAND2_X1 u0_u2_u4_U63 (.A1( u0_u2_u4_n100 ) , .ZN( u0_u2_u4_n118 ) , .A2( u0_u2_u4_n99 ) );
  NAND2_X1 u0_u2_u4_U64 (.A2( u0_u2_u4_n100 ) , .A1( u0_u2_u4_n102 ) , .ZN( u0_u2_u4_n144 ) );
  NAND2_X1 u0_u2_u4_U65 (.A2( u0_u2_u4_n101 ) , .A1( u0_u2_u4_n105 ) , .ZN( u0_u2_u4_n96 ) );
  INV_X1 u0_u2_u4_U66 (.A( u0_u2_u4_n128 ) , .ZN( u0_u2_u4_n174 ) );
  NAND2_X1 u0_u2_u4_U67 (.A2( u0_u2_u4_n102 ) , .ZN( u0_u2_u4_n119 ) , .A1( u0_u2_u4_n98 ) );
  NAND2_X1 u0_u2_u4_U68 (.A2( u0_u2_u4_n101 ) , .A1( u0_u2_u4_n103 ) , .ZN( u0_u2_u4_n147 ) );
  NAND2_X1 u0_u2_u4_U69 (.A2( u0_u2_u4_n104 ) , .ZN( u0_u2_u4_n113 ) , .A1( u0_u2_u4_n99 ) );
  AOI21_X1 u0_u2_u4_U7 (.ZN( u0_u2_u4_n108 ) , .B2( u0_u2_u4_n134 ) , .B1( u0_u2_u4_n155 ) , .A( u0_u2_u4_n156 ) );
  NOR2_X1 u0_u2_u4_U70 (.A2( u0_u2_X_28 ) , .ZN( u0_u2_u4_n150 ) , .A1( u0_u2_u4_n168 ) );
  NOR2_X1 u0_u2_u4_U71 (.A2( u0_u2_X_29 ) , .ZN( u0_u2_u4_n152 ) , .A1( u0_u2_u4_n169 ) );
  NOR2_X1 u0_u2_u4_U72 (.A2( u0_u2_X_30 ) , .ZN( u0_u2_u4_n105 ) , .A1( u0_u2_u4_n176 ) );
  NOR2_X1 u0_u2_u4_U73 (.A2( u0_u2_X_26 ) , .ZN( u0_u2_u4_n100 ) , .A1( u0_u2_u4_n177 ) );
  NOR2_X1 u0_u2_u4_U74 (.A2( u0_u2_X_28 ) , .A1( u0_u2_X_29 ) , .ZN( u0_u2_u4_n128 ) );
  NOR2_X1 u0_u2_u4_U75 (.A2( u0_u2_X_27 ) , .A1( u0_u2_X_30 ) , .ZN( u0_u2_u4_n102 ) );
  NOR2_X1 u0_u2_u4_U76 (.A2( u0_u2_X_25 ) , .A1( u0_u2_X_26 ) , .ZN( u0_u2_u4_n98 ) );
  AND2_X1 u0_u2_u4_U77 (.A2( u0_u2_X_25 ) , .A1( u0_u2_X_26 ) , .ZN( u0_u2_u4_n104 ) );
  AND2_X1 u0_u2_u4_U78 (.A1( u0_u2_X_30 ) , .A2( u0_u2_u4_n176 ) , .ZN( u0_u2_u4_n99 ) );
  AND2_X1 u0_u2_u4_U79 (.A1( u0_u2_X_26 ) , .ZN( u0_u2_u4_n101 ) , .A2( u0_u2_u4_n177 ) );
  AOI21_X1 u0_u2_u4_U8 (.ZN( u0_u2_u4_n109 ) , .A( u0_u2_u4_n153 ) , .B1( u0_u2_u4_n159 ) , .B2( u0_u2_u4_n184 ) );
  AND2_X1 u0_u2_u4_U80 (.A1( u0_u2_X_27 ) , .A2( u0_u2_X_30 ) , .ZN( u0_u2_u4_n103 ) );
  INV_X1 u0_u2_u4_U81 (.A( u0_u2_X_28 ) , .ZN( u0_u2_u4_n169 ) );
  INV_X1 u0_u2_u4_U82 (.A( u0_u2_X_29 ) , .ZN( u0_u2_u4_n168 ) );
  INV_X1 u0_u2_u4_U83 (.A( u0_u2_X_25 ) , .ZN( u0_u2_u4_n177 ) );
  INV_X1 u0_u2_u4_U84 (.A( u0_u2_X_27 ) , .ZN( u0_u2_u4_n176 ) );
  NAND4_X1 u0_u2_u4_U85 (.ZN( u0_out2_25 ) , .A4( u0_u2_u4_n139 ) , .A3( u0_u2_u4_n140 ) , .A2( u0_u2_u4_n141 ) , .A1( u0_u2_u4_n142 ) );
  OAI21_X1 u0_u2_u4_U86 (.A( u0_u2_u4_n128 ) , .B2( u0_u2_u4_n129 ) , .B1( u0_u2_u4_n130 ) , .ZN( u0_u2_u4_n142 ) );
  OAI21_X1 u0_u2_u4_U87 (.B2( u0_u2_u4_n131 ) , .ZN( u0_u2_u4_n141 ) , .A( u0_u2_u4_n175 ) , .B1( u0_u2_u4_n183 ) );
  NAND4_X1 u0_u2_u4_U88 (.ZN( u0_out2_14 ) , .A4( u0_u2_u4_n124 ) , .A3( u0_u2_u4_n125 ) , .A2( u0_u2_u4_n126 ) , .A1( u0_u2_u4_n127 ) );
  AOI22_X1 u0_u2_u4_U89 (.B2( u0_u2_u4_n117 ) , .ZN( u0_u2_u4_n126 ) , .A1( u0_u2_u4_n129 ) , .B1( u0_u2_u4_n152 ) , .A2( u0_u2_u4_n175 ) );
  AOI211_X1 u0_u2_u4_U9 (.B( u0_u2_u4_n136 ) , .A( u0_u2_u4_n137 ) , .C2( u0_u2_u4_n138 ) , .ZN( u0_u2_u4_n139 ) , .C1( u0_u2_u4_n182 ) );
  AOI22_X1 u0_u2_u4_U90 (.ZN( u0_u2_u4_n125 ) , .B2( u0_u2_u4_n131 ) , .A2( u0_u2_u4_n132 ) , .B1( u0_u2_u4_n138 ) , .A1( u0_u2_u4_n178 ) );
  NAND4_X1 u0_u2_u4_U91 (.ZN( u0_out2_8 ) , .A4( u0_u2_u4_n110 ) , .A3( u0_u2_u4_n111 ) , .A2( u0_u2_u4_n112 ) , .A1( u0_u2_u4_n186 ) );
  NAND2_X1 u0_u2_u4_U92 (.ZN( u0_u2_u4_n112 ) , .A2( u0_u2_u4_n130 ) , .A1( u0_u2_u4_n150 ) );
  AOI22_X1 u0_u2_u4_U93 (.ZN( u0_u2_u4_n111 ) , .B2( u0_u2_u4_n132 ) , .A1( u0_u2_u4_n152 ) , .B1( u0_u2_u4_n178 ) , .A2( u0_u2_u4_n97 ) );
  AOI22_X1 u0_u2_u4_U94 (.B2( u0_u2_u4_n149 ) , .B1( u0_u2_u4_n150 ) , .A2( u0_u2_u4_n151 ) , .A1( u0_u2_u4_n152 ) , .ZN( u0_u2_u4_n167 ) );
  NOR4_X1 u0_u2_u4_U95 (.A4( u0_u2_u4_n162 ) , .A3( u0_u2_u4_n163 ) , .A2( u0_u2_u4_n164 ) , .A1( u0_u2_u4_n165 ) , .ZN( u0_u2_u4_n166 ) );
  NAND3_X1 u0_u2_u4_U96 (.ZN( u0_out2_3 ) , .A3( u0_u2_u4_n166 ) , .A1( u0_u2_u4_n167 ) , .A2( u0_u2_u4_n186 ) );
  NAND3_X1 u0_u2_u4_U97 (.A3( u0_u2_u4_n146 ) , .A2( u0_u2_u4_n147 ) , .A1( u0_u2_u4_n148 ) , .ZN( u0_u2_u4_n149 ) );
  NAND3_X1 u0_u2_u4_U98 (.A3( u0_u2_u4_n143 ) , .A2( u0_u2_u4_n144 ) , .A1( u0_u2_u4_n145 ) , .ZN( u0_u2_u4_n151 ) );
  NAND3_X1 u0_u2_u4_U99 (.A3( u0_u2_u4_n121 ) , .ZN( u0_u2_u4_n122 ) , .A2( u0_u2_u4_n144 ) , .A1( u0_u2_u4_n154 ) );
  XOR2_X1 u0_u3_U10 (.B( u0_K4_45 ) , .A( u0_R2_30 ) , .Z( u0_u3_X_45 ) );
  XOR2_X1 u0_u3_U11 (.B( u0_K4_44 ) , .A( u0_R2_29 ) , .Z( u0_u3_X_44 ) );
  XOR2_X1 u0_u3_U12 (.B( u0_K4_43 ) , .A( u0_R2_28 ) , .Z( u0_u3_X_43 ) );
  XOR2_X1 u0_u3_U13 (.B( u0_K4_42 ) , .A( u0_R2_29 ) , .Z( u0_u3_X_42 ) );
  XOR2_X1 u0_u3_U14 (.B( u0_K4_41 ) , .A( u0_R2_28 ) , .Z( u0_u3_X_41 ) );
  XOR2_X1 u0_u3_U15 (.B( u0_K4_40 ) , .A( u0_R2_27 ) , .Z( u0_u3_X_40 ) );
  XOR2_X1 u0_u3_U17 (.B( u0_K4_39 ) , .A( u0_R2_26 ) , .Z( u0_u3_X_39 ) );
  XOR2_X1 u0_u3_U18 (.B( u0_K4_38 ) , .A( u0_R2_25 ) , .Z( u0_u3_X_38 ) );
  XOR2_X1 u0_u3_U19 (.B( u0_K4_37 ) , .A( u0_R2_24 ) , .Z( u0_u3_X_37 ) );
  XOR2_X1 u0_u3_U7 (.B( u0_K4_48 ) , .A( u0_R2_1 ) , .Z( u0_u3_X_48 ) );
  XOR2_X1 u0_u3_U8 (.B( u0_K4_47 ) , .A( u0_R2_32 ) , .Z( u0_u3_X_47 ) );
  XOR2_X1 u0_u3_U9 (.B( u0_K4_46 ) , .A( u0_R2_31 ) , .Z( u0_u3_X_46 ) );
  INV_X1 u0_u3_u6_U10 (.ZN( u0_u3_u6_n172 ) , .A( u0_u3_u6_n88 ) );
  OAI21_X1 u0_u3_u6_U11 (.A( u0_u3_u6_n159 ) , .B1( u0_u3_u6_n169 ) , .B2( u0_u3_u6_n173 ) , .ZN( u0_u3_u6_n90 ) );
  AOI22_X1 u0_u3_u6_U12 (.A2( u0_u3_u6_n151 ) , .B2( u0_u3_u6_n161 ) , .A1( u0_u3_u6_n167 ) , .B1( u0_u3_u6_n170 ) , .ZN( u0_u3_u6_n89 ) );
  AOI21_X1 u0_u3_u6_U13 (.ZN( u0_u3_u6_n106 ) , .A( u0_u3_u6_n142 ) , .B2( u0_u3_u6_n159 ) , .B1( u0_u3_u6_n164 ) );
  INV_X1 u0_u3_u6_U14 (.A( u0_u3_u6_n155 ) , .ZN( u0_u3_u6_n161 ) );
  INV_X1 u0_u3_u6_U15 (.A( u0_u3_u6_n128 ) , .ZN( u0_u3_u6_n164 ) );
  NAND2_X1 u0_u3_u6_U16 (.ZN( u0_u3_u6_n110 ) , .A1( u0_u3_u6_n122 ) , .A2( u0_u3_u6_n129 ) );
  NAND2_X1 u0_u3_u6_U17 (.ZN( u0_u3_u6_n124 ) , .A2( u0_u3_u6_n146 ) , .A1( u0_u3_u6_n148 ) );
  INV_X1 u0_u3_u6_U18 (.A( u0_u3_u6_n132 ) , .ZN( u0_u3_u6_n171 ) );
  AND2_X1 u0_u3_u6_U19 (.A1( u0_u3_u6_n100 ) , .ZN( u0_u3_u6_n130 ) , .A2( u0_u3_u6_n147 ) );
  INV_X1 u0_u3_u6_U20 (.A( u0_u3_u6_n127 ) , .ZN( u0_u3_u6_n173 ) );
  INV_X1 u0_u3_u6_U21 (.A( u0_u3_u6_n121 ) , .ZN( u0_u3_u6_n167 ) );
  INV_X1 u0_u3_u6_U22 (.A( u0_u3_u6_n100 ) , .ZN( u0_u3_u6_n169 ) );
  INV_X1 u0_u3_u6_U23 (.A( u0_u3_u6_n123 ) , .ZN( u0_u3_u6_n170 ) );
  INV_X1 u0_u3_u6_U24 (.A( u0_u3_u6_n113 ) , .ZN( u0_u3_u6_n168 ) );
  AND2_X1 u0_u3_u6_U25 (.A1( u0_u3_u6_n107 ) , .A2( u0_u3_u6_n119 ) , .ZN( u0_u3_u6_n133 ) );
  AND2_X1 u0_u3_u6_U26 (.A2( u0_u3_u6_n121 ) , .A1( u0_u3_u6_n122 ) , .ZN( u0_u3_u6_n131 ) );
  AND3_X1 u0_u3_u6_U27 (.ZN( u0_u3_u6_n120 ) , .A2( u0_u3_u6_n127 ) , .A1( u0_u3_u6_n132 ) , .A3( u0_u3_u6_n145 ) );
  INV_X1 u0_u3_u6_U28 (.A( u0_u3_u6_n146 ) , .ZN( u0_u3_u6_n163 ) );
  AOI222_X1 u0_u3_u6_U29 (.ZN( u0_u3_u6_n114 ) , .A1( u0_u3_u6_n118 ) , .A2( u0_u3_u6_n126 ) , .B2( u0_u3_u6_n151 ) , .C2( u0_u3_u6_n159 ) , .C1( u0_u3_u6_n168 ) , .B1( u0_u3_u6_n169 ) );
  INV_X1 u0_u3_u6_U3 (.A( u0_u3_u6_n110 ) , .ZN( u0_u3_u6_n166 ) );
  NOR2_X1 u0_u3_u6_U30 (.A1( u0_u3_u6_n162 ) , .A2( u0_u3_u6_n165 ) , .ZN( u0_u3_u6_n98 ) );
  NAND2_X1 u0_u3_u6_U31 (.A1( u0_u3_u6_n144 ) , .ZN( u0_u3_u6_n151 ) , .A2( u0_u3_u6_n158 ) );
  NAND2_X1 u0_u3_u6_U32 (.ZN( u0_u3_u6_n132 ) , .A1( u0_u3_u6_n91 ) , .A2( u0_u3_u6_n97 ) );
  AOI22_X1 u0_u3_u6_U33 (.B2( u0_u3_u6_n110 ) , .B1( u0_u3_u6_n111 ) , .A1( u0_u3_u6_n112 ) , .ZN( u0_u3_u6_n115 ) , .A2( u0_u3_u6_n161 ) );
  NAND4_X1 u0_u3_u6_U34 (.A3( u0_u3_u6_n109 ) , .ZN( u0_u3_u6_n112 ) , .A4( u0_u3_u6_n132 ) , .A2( u0_u3_u6_n147 ) , .A1( u0_u3_u6_n166 ) );
  NOR2_X1 u0_u3_u6_U35 (.ZN( u0_u3_u6_n109 ) , .A1( u0_u3_u6_n170 ) , .A2( u0_u3_u6_n173 ) );
  NOR2_X1 u0_u3_u6_U36 (.A2( u0_u3_u6_n126 ) , .ZN( u0_u3_u6_n155 ) , .A1( u0_u3_u6_n160 ) );
  NAND2_X1 u0_u3_u6_U37 (.ZN( u0_u3_u6_n146 ) , .A2( u0_u3_u6_n94 ) , .A1( u0_u3_u6_n99 ) );
  AOI21_X1 u0_u3_u6_U38 (.A( u0_u3_u6_n144 ) , .B2( u0_u3_u6_n145 ) , .B1( u0_u3_u6_n146 ) , .ZN( u0_u3_u6_n150 ) );
  AOI211_X1 u0_u3_u6_U39 (.B( u0_u3_u6_n134 ) , .A( u0_u3_u6_n135 ) , .C1( u0_u3_u6_n136 ) , .ZN( u0_u3_u6_n137 ) , .C2( u0_u3_u6_n151 ) );
  INV_X1 u0_u3_u6_U4 (.A( u0_u3_u6_n142 ) , .ZN( u0_u3_u6_n174 ) );
  AOI21_X1 u0_u3_u6_U40 (.B2( u0_u3_u6_n132 ) , .B1( u0_u3_u6_n133 ) , .ZN( u0_u3_u6_n134 ) , .A( u0_u3_u6_n158 ) );
  NAND4_X1 u0_u3_u6_U41 (.A4( u0_u3_u6_n127 ) , .A3( u0_u3_u6_n128 ) , .A2( u0_u3_u6_n129 ) , .A1( u0_u3_u6_n130 ) , .ZN( u0_u3_u6_n136 ) );
  AOI21_X1 u0_u3_u6_U42 (.B1( u0_u3_u6_n131 ) , .ZN( u0_u3_u6_n135 ) , .A( u0_u3_u6_n144 ) , .B2( u0_u3_u6_n146 ) );
  INV_X1 u0_u3_u6_U43 (.A( u0_u3_u6_n111 ) , .ZN( u0_u3_u6_n158 ) );
  NAND2_X1 u0_u3_u6_U44 (.ZN( u0_u3_u6_n127 ) , .A1( u0_u3_u6_n91 ) , .A2( u0_u3_u6_n92 ) );
  NAND2_X1 u0_u3_u6_U45 (.ZN( u0_u3_u6_n129 ) , .A2( u0_u3_u6_n95 ) , .A1( u0_u3_u6_n96 ) );
  INV_X1 u0_u3_u6_U46 (.A( u0_u3_u6_n144 ) , .ZN( u0_u3_u6_n159 ) );
  NAND2_X1 u0_u3_u6_U47 (.ZN( u0_u3_u6_n145 ) , .A2( u0_u3_u6_n97 ) , .A1( u0_u3_u6_n98 ) );
  NAND2_X1 u0_u3_u6_U48 (.ZN( u0_u3_u6_n148 ) , .A2( u0_u3_u6_n92 ) , .A1( u0_u3_u6_n94 ) );
  NAND2_X1 u0_u3_u6_U49 (.ZN( u0_u3_u6_n108 ) , .A2( u0_u3_u6_n139 ) , .A1( u0_u3_u6_n144 ) );
  NAND2_X1 u0_u3_u6_U5 (.A2( u0_u3_u6_n143 ) , .ZN( u0_u3_u6_n152 ) , .A1( u0_u3_u6_n166 ) );
  NAND2_X1 u0_u3_u6_U50 (.ZN( u0_u3_u6_n121 ) , .A2( u0_u3_u6_n95 ) , .A1( u0_u3_u6_n97 ) );
  NAND2_X1 u0_u3_u6_U51 (.ZN( u0_u3_u6_n107 ) , .A2( u0_u3_u6_n92 ) , .A1( u0_u3_u6_n95 ) );
  AND2_X1 u0_u3_u6_U52 (.ZN( u0_u3_u6_n118 ) , .A2( u0_u3_u6_n91 ) , .A1( u0_u3_u6_n99 ) );
  NAND2_X1 u0_u3_u6_U53 (.ZN( u0_u3_u6_n147 ) , .A2( u0_u3_u6_n98 ) , .A1( u0_u3_u6_n99 ) );
  NAND2_X1 u0_u3_u6_U54 (.ZN( u0_u3_u6_n128 ) , .A1( u0_u3_u6_n94 ) , .A2( u0_u3_u6_n96 ) );
  NAND2_X1 u0_u3_u6_U55 (.ZN( u0_u3_u6_n119 ) , .A2( u0_u3_u6_n95 ) , .A1( u0_u3_u6_n99 ) );
  NAND2_X1 u0_u3_u6_U56 (.ZN( u0_u3_u6_n123 ) , .A2( u0_u3_u6_n91 ) , .A1( u0_u3_u6_n96 ) );
  NAND2_X1 u0_u3_u6_U57 (.ZN( u0_u3_u6_n100 ) , .A2( u0_u3_u6_n92 ) , .A1( u0_u3_u6_n98 ) );
  NAND2_X1 u0_u3_u6_U58 (.ZN( u0_u3_u6_n122 ) , .A1( u0_u3_u6_n94 ) , .A2( u0_u3_u6_n97 ) );
  INV_X1 u0_u3_u6_U59 (.A( u0_u3_u6_n139 ) , .ZN( u0_u3_u6_n160 ) );
  AOI22_X1 u0_u3_u6_U6 (.B2( u0_u3_u6_n101 ) , .A1( u0_u3_u6_n102 ) , .ZN( u0_u3_u6_n103 ) , .B1( u0_u3_u6_n160 ) , .A2( u0_u3_u6_n161 ) );
  NAND2_X1 u0_u3_u6_U60 (.ZN( u0_u3_u6_n113 ) , .A1( u0_u3_u6_n96 ) , .A2( u0_u3_u6_n98 ) );
  NOR2_X1 u0_u3_u6_U61 (.A2( u0_u3_X_40 ) , .A1( u0_u3_X_41 ) , .ZN( u0_u3_u6_n126 ) );
  NOR2_X1 u0_u3_u6_U62 (.A2( u0_u3_X_39 ) , .A1( u0_u3_X_42 ) , .ZN( u0_u3_u6_n92 ) );
  NOR2_X1 u0_u3_u6_U63 (.A2( u0_u3_X_39 ) , .A1( u0_u3_u6_n156 ) , .ZN( u0_u3_u6_n97 ) );
  NOR2_X1 u0_u3_u6_U64 (.A2( u0_u3_X_38 ) , .A1( u0_u3_u6_n165 ) , .ZN( u0_u3_u6_n95 ) );
  NOR2_X1 u0_u3_u6_U65 (.A2( u0_u3_X_41 ) , .ZN( u0_u3_u6_n111 ) , .A1( u0_u3_u6_n157 ) );
  NOR2_X1 u0_u3_u6_U66 (.A2( u0_u3_X_37 ) , .A1( u0_u3_u6_n162 ) , .ZN( u0_u3_u6_n94 ) );
  NOR2_X1 u0_u3_u6_U67 (.A2( u0_u3_X_37 ) , .A1( u0_u3_X_38 ) , .ZN( u0_u3_u6_n91 ) );
  NAND2_X1 u0_u3_u6_U68 (.A1( u0_u3_X_41 ) , .ZN( u0_u3_u6_n144 ) , .A2( u0_u3_u6_n157 ) );
  NAND2_X1 u0_u3_u6_U69 (.A2( u0_u3_X_40 ) , .A1( u0_u3_X_41 ) , .ZN( u0_u3_u6_n139 ) );
  NOR2_X1 u0_u3_u6_U7 (.A1( u0_u3_u6_n118 ) , .ZN( u0_u3_u6_n143 ) , .A2( u0_u3_u6_n168 ) );
  AND2_X1 u0_u3_u6_U70 (.A1( u0_u3_X_39 ) , .A2( u0_u3_u6_n156 ) , .ZN( u0_u3_u6_n96 ) );
  AND2_X1 u0_u3_u6_U71 (.A1( u0_u3_X_39 ) , .A2( u0_u3_X_42 ) , .ZN( u0_u3_u6_n99 ) );
  INV_X1 u0_u3_u6_U72 (.A( u0_u3_X_40 ) , .ZN( u0_u3_u6_n157 ) );
  INV_X1 u0_u3_u6_U73 (.A( u0_u3_X_37 ) , .ZN( u0_u3_u6_n165 ) );
  INV_X1 u0_u3_u6_U74 (.A( u0_u3_X_38 ) , .ZN( u0_u3_u6_n162 ) );
  INV_X1 u0_u3_u6_U75 (.A( u0_u3_X_42 ) , .ZN( u0_u3_u6_n156 ) );
  NAND4_X1 u0_u3_u6_U76 (.ZN( u0_out3_32 ) , .A4( u0_u3_u6_n103 ) , .A3( u0_u3_u6_n104 ) , .A2( u0_u3_u6_n105 ) , .A1( u0_u3_u6_n106 ) );
  AOI22_X1 u0_u3_u6_U77 (.ZN( u0_u3_u6_n105 ) , .A2( u0_u3_u6_n108 ) , .A1( u0_u3_u6_n118 ) , .B2( u0_u3_u6_n126 ) , .B1( u0_u3_u6_n171 ) );
  AOI22_X1 u0_u3_u6_U78 (.ZN( u0_u3_u6_n104 ) , .A1( u0_u3_u6_n111 ) , .B1( u0_u3_u6_n124 ) , .B2( u0_u3_u6_n151 ) , .A2( u0_u3_u6_n93 ) );
  NAND4_X1 u0_u3_u6_U79 (.ZN( u0_out3_12 ) , .A4( u0_u3_u6_n114 ) , .A3( u0_u3_u6_n115 ) , .A2( u0_u3_u6_n116 ) , .A1( u0_u3_u6_n117 ) );
  AOI21_X1 u0_u3_u6_U8 (.B1( u0_u3_u6_n107 ) , .B2( u0_u3_u6_n132 ) , .A( u0_u3_u6_n158 ) , .ZN( u0_u3_u6_n88 ) );
  OAI22_X1 u0_u3_u6_U80 (.B2( u0_u3_u6_n111 ) , .ZN( u0_u3_u6_n116 ) , .B1( u0_u3_u6_n126 ) , .A2( u0_u3_u6_n164 ) , .A1( u0_u3_u6_n167 ) );
  OAI21_X1 u0_u3_u6_U81 (.A( u0_u3_u6_n108 ) , .ZN( u0_u3_u6_n117 ) , .B2( u0_u3_u6_n141 ) , .B1( u0_u3_u6_n163 ) );
  OAI211_X1 u0_u3_u6_U82 (.ZN( u0_out3_22 ) , .B( u0_u3_u6_n137 ) , .A( u0_u3_u6_n138 ) , .C2( u0_u3_u6_n139 ) , .C1( u0_u3_u6_n140 ) );
  AOI22_X1 u0_u3_u6_U83 (.B1( u0_u3_u6_n124 ) , .A2( u0_u3_u6_n125 ) , .A1( u0_u3_u6_n126 ) , .ZN( u0_u3_u6_n138 ) , .B2( u0_u3_u6_n161 ) );
  AND4_X1 u0_u3_u6_U84 (.A3( u0_u3_u6_n119 ) , .A1( u0_u3_u6_n120 ) , .A4( u0_u3_u6_n129 ) , .ZN( u0_u3_u6_n140 ) , .A2( u0_u3_u6_n143 ) );
  OAI211_X1 u0_u3_u6_U85 (.ZN( u0_out3_7 ) , .B( u0_u3_u6_n153 ) , .C2( u0_u3_u6_n154 ) , .C1( u0_u3_u6_n155 ) , .A( u0_u3_u6_n174 ) );
  NOR3_X1 u0_u3_u6_U86 (.A1( u0_u3_u6_n141 ) , .ZN( u0_u3_u6_n154 ) , .A3( u0_u3_u6_n164 ) , .A2( u0_u3_u6_n171 ) );
  AOI211_X1 u0_u3_u6_U87 (.B( u0_u3_u6_n149 ) , .A( u0_u3_u6_n150 ) , .C2( u0_u3_u6_n151 ) , .C1( u0_u3_u6_n152 ) , .ZN( u0_u3_u6_n153 ) );
  NAND3_X1 u0_u3_u6_U88 (.A2( u0_u3_u6_n123 ) , .ZN( u0_u3_u6_n125 ) , .A1( u0_u3_u6_n130 ) , .A3( u0_u3_u6_n131 ) );
  NAND3_X1 u0_u3_u6_U89 (.A3( u0_u3_u6_n133 ) , .ZN( u0_u3_u6_n141 ) , .A1( u0_u3_u6_n145 ) , .A2( u0_u3_u6_n148 ) );
  AOI21_X1 u0_u3_u6_U9 (.B2( u0_u3_u6_n147 ) , .B1( u0_u3_u6_n148 ) , .ZN( u0_u3_u6_n149 ) , .A( u0_u3_u6_n158 ) );
  NAND3_X1 u0_u3_u6_U90 (.ZN( u0_u3_u6_n101 ) , .A3( u0_u3_u6_n107 ) , .A2( u0_u3_u6_n121 ) , .A1( u0_u3_u6_n127 ) );
  NAND3_X1 u0_u3_u6_U91 (.ZN( u0_u3_u6_n102 ) , .A3( u0_u3_u6_n130 ) , .A2( u0_u3_u6_n145 ) , .A1( u0_u3_u6_n166 ) );
  NAND3_X1 u0_u3_u6_U92 (.A3( u0_u3_u6_n113 ) , .A1( u0_u3_u6_n119 ) , .A2( u0_u3_u6_n123 ) , .ZN( u0_u3_u6_n93 ) );
  NAND3_X1 u0_u3_u6_U93 (.ZN( u0_u3_u6_n142 ) , .A2( u0_u3_u6_n172 ) , .A3( u0_u3_u6_n89 ) , .A1( u0_u3_u6_n90 ) );
  AND3_X1 u0_u3_u7_U10 (.A3( u0_u3_u7_n110 ) , .A2( u0_u3_u7_n127 ) , .A1( u0_u3_u7_n132 ) , .ZN( u0_u3_u7_n92 ) );
  OAI21_X1 u0_u3_u7_U11 (.A( u0_u3_u7_n161 ) , .B1( u0_u3_u7_n168 ) , .B2( u0_u3_u7_n173 ) , .ZN( u0_u3_u7_n91 ) );
  AOI211_X1 u0_u3_u7_U12 (.A( u0_u3_u7_n117 ) , .ZN( u0_u3_u7_n118 ) , .C2( u0_u3_u7_n126 ) , .C1( u0_u3_u7_n177 ) , .B( u0_u3_u7_n180 ) );
  OAI22_X1 u0_u3_u7_U13 (.B1( u0_u3_u7_n115 ) , .ZN( u0_u3_u7_n117 ) , .A2( u0_u3_u7_n133 ) , .A1( u0_u3_u7_n137 ) , .B2( u0_u3_u7_n162 ) );
  INV_X1 u0_u3_u7_U14 (.A( u0_u3_u7_n116 ) , .ZN( u0_u3_u7_n180 ) );
  NOR3_X1 u0_u3_u7_U15 (.ZN( u0_u3_u7_n115 ) , .A3( u0_u3_u7_n145 ) , .A2( u0_u3_u7_n168 ) , .A1( u0_u3_u7_n169 ) );
  OAI211_X1 u0_u3_u7_U16 (.B( u0_u3_u7_n122 ) , .A( u0_u3_u7_n123 ) , .C2( u0_u3_u7_n124 ) , .ZN( u0_u3_u7_n154 ) , .C1( u0_u3_u7_n162 ) );
  AOI222_X1 u0_u3_u7_U17 (.ZN( u0_u3_u7_n122 ) , .C2( u0_u3_u7_n126 ) , .C1( u0_u3_u7_n145 ) , .B1( u0_u3_u7_n161 ) , .A2( u0_u3_u7_n165 ) , .B2( u0_u3_u7_n170 ) , .A1( u0_u3_u7_n176 ) );
  INV_X1 u0_u3_u7_U18 (.A( u0_u3_u7_n133 ) , .ZN( u0_u3_u7_n176 ) );
  NOR3_X1 u0_u3_u7_U19 (.A2( u0_u3_u7_n134 ) , .A1( u0_u3_u7_n135 ) , .ZN( u0_u3_u7_n136 ) , .A3( u0_u3_u7_n171 ) );
  NOR2_X1 u0_u3_u7_U20 (.A1( u0_u3_u7_n130 ) , .A2( u0_u3_u7_n134 ) , .ZN( u0_u3_u7_n153 ) );
  INV_X1 u0_u3_u7_U21 (.A( u0_u3_u7_n101 ) , .ZN( u0_u3_u7_n165 ) );
  NOR2_X1 u0_u3_u7_U22 (.ZN( u0_u3_u7_n111 ) , .A2( u0_u3_u7_n134 ) , .A1( u0_u3_u7_n169 ) );
  AOI21_X1 u0_u3_u7_U23 (.ZN( u0_u3_u7_n104 ) , .B2( u0_u3_u7_n112 ) , .B1( u0_u3_u7_n127 ) , .A( u0_u3_u7_n164 ) );
  AOI21_X1 u0_u3_u7_U24 (.ZN( u0_u3_u7_n106 ) , .B1( u0_u3_u7_n133 ) , .B2( u0_u3_u7_n146 ) , .A( u0_u3_u7_n162 ) );
  AOI21_X1 u0_u3_u7_U25 (.A( u0_u3_u7_n101 ) , .ZN( u0_u3_u7_n107 ) , .B2( u0_u3_u7_n128 ) , .B1( u0_u3_u7_n175 ) );
  INV_X1 u0_u3_u7_U26 (.A( u0_u3_u7_n138 ) , .ZN( u0_u3_u7_n171 ) );
  INV_X1 u0_u3_u7_U27 (.A( u0_u3_u7_n131 ) , .ZN( u0_u3_u7_n177 ) );
  INV_X1 u0_u3_u7_U28 (.A( u0_u3_u7_n110 ) , .ZN( u0_u3_u7_n174 ) );
  NAND2_X1 u0_u3_u7_U29 (.A1( u0_u3_u7_n129 ) , .A2( u0_u3_u7_n132 ) , .ZN( u0_u3_u7_n149 ) );
  OAI21_X1 u0_u3_u7_U3 (.ZN( u0_u3_u7_n159 ) , .A( u0_u3_u7_n165 ) , .B2( u0_u3_u7_n171 ) , .B1( u0_u3_u7_n174 ) );
  NAND2_X1 u0_u3_u7_U30 (.A1( u0_u3_u7_n113 ) , .A2( u0_u3_u7_n124 ) , .ZN( u0_u3_u7_n130 ) );
  INV_X1 u0_u3_u7_U31 (.A( u0_u3_u7_n112 ) , .ZN( u0_u3_u7_n173 ) );
  INV_X1 u0_u3_u7_U32 (.A( u0_u3_u7_n128 ) , .ZN( u0_u3_u7_n168 ) );
  INV_X1 u0_u3_u7_U33 (.A( u0_u3_u7_n148 ) , .ZN( u0_u3_u7_n169 ) );
  INV_X1 u0_u3_u7_U34 (.A( u0_u3_u7_n127 ) , .ZN( u0_u3_u7_n179 ) );
  NOR2_X1 u0_u3_u7_U35 (.ZN( u0_u3_u7_n101 ) , .A2( u0_u3_u7_n150 ) , .A1( u0_u3_u7_n156 ) );
  AOI211_X1 u0_u3_u7_U36 (.B( u0_u3_u7_n154 ) , .A( u0_u3_u7_n155 ) , .C1( u0_u3_u7_n156 ) , .ZN( u0_u3_u7_n157 ) , .C2( u0_u3_u7_n172 ) );
  INV_X1 u0_u3_u7_U37 (.A( u0_u3_u7_n153 ) , .ZN( u0_u3_u7_n172 ) );
  AOI211_X1 u0_u3_u7_U38 (.B( u0_u3_u7_n139 ) , .A( u0_u3_u7_n140 ) , .C2( u0_u3_u7_n141 ) , .ZN( u0_u3_u7_n142 ) , .C1( u0_u3_u7_n156 ) );
  NAND4_X1 u0_u3_u7_U39 (.A3( u0_u3_u7_n127 ) , .A2( u0_u3_u7_n128 ) , .A1( u0_u3_u7_n129 ) , .ZN( u0_u3_u7_n141 ) , .A4( u0_u3_u7_n147 ) );
  INV_X1 u0_u3_u7_U4 (.A( u0_u3_u7_n111 ) , .ZN( u0_u3_u7_n170 ) );
  AOI21_X1 u0_u3_u7_U40 (.A( u0_u3_u7_n137 ) , .B1( u0_u3_u7_n138 ) , .ZN( u0_u3_u7_n139 ) , .B2( u0_u3_u7_n146 ) );
  OAI22_X1 u0_u3_u7_U41 (.B1( u0_u3_u7_n136 ) , .ZN( u0_u3_u7_n140 ) , .A1( u0_u3_u7_n153 ) , .B2( u0_u3_u7_n162 ) , .A2( u0_u3_u7_n164 ) );
  AOI21_X1 u0_u3_u7_U42 (.ZN( u0_u3_u7_n123 ) , .B1( u0_u3_u7_n165 ) , .B2( u0_u3_u7_n177 ) , .A( u0_u3_u7_n97 ) );
  AOI21_X1 u0_u3_u7_U43 (.B2( u0_u3_u7_n113 ) , .B1( u0_u3_u7_n124 ) , .A( u0_u3_u7_n125 ) , .ZN( u0_u3_u7_n97 ) );
  INV_X1 u0_u3_u7_U44 (.A( u0_u3_u7_n125 ) , .ZN( u0_u3_u7_n161 ) );
  INV_X1 u0_u3_u7_U45 (.A( u0_u3_u7_n152 ) , .ZN( u0_u3_u7_n162 ) );
  AOI22_X1 u0_u3_u7_U46 (.A2( u0_u3_u7_n114 ) , .ZN( u0_u3_u7_n119 ) , .B1( u0_u3_u7_n130 ) , .A1( u0_u3_u7_n156 ) , .B2( u0_u3_u7_n165 ) );
  NAND2_X1 u0_u3_u7_U47 (.A2( u0_u3_u7_n112 ) , .ZN( u0_u3_u7_n114 ) , .A1( u0_u3_u7_n175 ) );
  AND2_X1 u0_u3_u7_U48 (.ZN( u0_u3_u7_n145 ) , .A2( u0_u3_u7_n98 ) , .A1( u0_u3_u7_n99 ) );
  NOR2_X1 u0_u3_u7_U49 (.ZN( u0_u3_u7_n137 ) , .A1( u0_u3_u7_n150 ) , .A2( u0_u3_u7_n161 ) );
  INV_X1 u0_u3_u7_U5 (.A( u0_u3_u7_n149 ) , .ZN( u0_u3_u7_n175 ) );
  AOI21_X1 u0_u3_u7_U50 (.ZN( u0_u3_u7_n105 ) , .B2( u0_u3_u7_n110 ) , .A( u0_u3_u7_n125 ) , .B1( u0_u3_u7_n147 ) );
  NAND2_X1 u0_u3_u7_U51 (.ZN( u0_u3_u7_n146 ) , .A1( u0_u3_u7_n95 ) , .A2( u0_u3_u7_n98 ) );
  NAND2_X1 u0_u3_u7_U52 (.A2( u0_u3_u7_n103 ) , .ZN( u0_u3_u7_n147 ) , .A1( u0_u3_u7_n93 ) );
  NAND2_X1 u0_u3_u7_U53 (.A1( u0_u3_u7_n103 ) , .ZN( u0_u3_u7_n127 ) , .A2( u0_u3_u7_n99 ) );
  OR2_X1 u0_u3_u7_U54 (.ZN( u0_u3_u7_n126 ) , .A2( u0_u3_u7_n152 ) , .A1( u0_u3_u7_n156 ) );
  NAND2_X1 u0_u3_u7_U55 (.A2( u0_u3_u7_n102 ) , .A1( u0_u3_u7_n103 ) , .ZN( u0_u3_u7_n133 ) );
  NAND2_X1 u0_u3_u7_U56 (.ZN( u0_u3_u7_n112 ) , .A2( u0_u3_u7_n96 ) , .A1( u0_u3_u7_n99 ) );
  NAND2_X1 u0_u3_u7_U57 (.A2( u0_u3_u7_n102 ) , .ZN( u0_u3_u7_n128 ) , .A1( u0_u3_u7_n98 ) );
  NAND2_X1 u0_u3_u7_U58 (.A1( u0_u3_u7_n100 ) , .ZN( u0_u3_u7_n113 ) , .A2( u0_u3_u7_n93 ) );
  NAND2_X1 u0_u3_u7_U59 (.A2( u0_u3_u7_n102 ) , .ZN( u0_u3_u7_n124 ) , .A1( u0_u3_u7_n96 ) );
  INV_X1 u0_u3_u7_U6 (.A( u0_u3_u7_n154 ) , .ZN( u0_u3_u7_n178 ) );
  NAND2_X1 u0_u3_u7_U60 (.ZN( u0_u3_u7_n110 ) , .A1( u0_u3_u7_n95 ) , .A2( u0_u3_u7_n96 ) );
  INV_X1 u0_u3_u7_U61 (.A( u0_u3_u7_n150 ) , .ZN( u0_u3_u7_n164 ) );
  AND2_X1 u0_u3_u7_U62 (.ZN( u0_u3_u7_n134 ) , .A1( u0_u3_u7_n93 ) , .A2( u0_u3_u7_n98 ) );
  NAND2_X1 u0_u3_u7_U63 (.A1( u0_u3_u7_n100 ) , .A2( u0_u3_u7_n102 ) , .ZN( u0_u3_u7_n129 ) );
  NAND2_X1 u0_u3_u7_U64 (.A2( u0_u3_u7_n103 ) , .ZN( u0_u3_u7_n131 ) , .A1( u0_u3_u7_n95 ) );
  NAND2_X1 u0_u3_u7_U65 (.A1( u0_u3_u7_n100 ) , .ZN( u0_u3_u7_n138 ) , .A2( u0_u3_u7_n99 ) );
  NAND2_X1 u0_u3_u7_U66 (.ZN( u0_u3_u7_n132 ) , .A1( u0_u3_u7_n93 ) , .A2( u0_u3_u7_n96 ) );
  NAND2_X1 u0_u3_u7_U67 (.A1( u0_u3_u7_n100 ) , .ZN( u0_u3_u7_n148 ) , .A2( u0_u3_u7_n95 ) );
  NOR2_X1 u0_u3_u7_U68 (.A2( u0_u3_X_47 ) , .ZN( u0_u3_u7_n150 ) , .A1( u0_u3_u7_n163 ) );
  NOR2_X1 u0_u3_u7_U69 (.A2( u0_u3_X_43 ) , .A1( u0_u3_X_44 ) , .ZN( u0_u3_u7_n103 ) );
  AOI211_X1 u0_u3_u7_U7 (.ZN( u0_u3_u7_n116 ) , .A( u0_u3_u7_n155 ) , .C1( u0_u3_u7_n161 ) , .C2( u0_u3_u7_n171 ) , .B( u0_u3_u7_n94 ) );
  NOR2_X1 u0_u3_u7_U70 (.A2( u0_u3_X_48 ) , .A1( u0_u3_u7_n166 ) , .ZN( u0_u3_u7_n95 ) );
  NOR2_X1 u0_u3_u7_U71 (.A2( u0_u3_X_45 ) , .A1( u0_u3_X_48 ) , .ZN( u0_u3_u7_n99 ) );
  NOR2_X1 u0_u3_u7_U72 (.A2( u0_u3_X_44 ) , .A1( u0_u3_u7_n167 ) , .ZN( u0_u3_u7_n98 ) );
  NOR2_X1 u0_u3_u7_U73 (.A2( u0_u3_X_46 ) , .A1( u0_u3_X_47 ) , .ZN( u0_u3_u7_n152 ) );
  AND2_X1 u0_u3_u7_U74 (.A1( u0_u3_X_47 ) , .ZN( u0_u3_u7_n156 ) , .A2( u0_u3_u7_n163 ) );
  NAND2_X1 u0_u3_u7_U75 (.A2( u0_u3_X_46 ) , .A1( u0_u3_X_47 ) , .ZN( u0_u3_u7_n125 ) );
  AND2_X1 u0_u3_u7_U76 (.A2( u0_u3_X_45 ) , .A1( u0_u3_X_48 ) , .ZN( u0_u3_u7_n102 ) );
  AND2_X1 u0_u3_u7_U77 (.A2( u0_u3_X_43 ) , .A1( u0_u3_X_44 ) , .ZN( u0_u3_u7_n96 ) );
  AND2_X1 u0_u3_u7_U78 (.A1( u0_u3_X_44 ) , .ZN( u0_u3_u7_n100 ) , .A2( u0_u3_u7_n167 ) );
  AND2_X1 u0_u3_u7_U79 (.A1( u0_u3_X_48 ) , .A2( u0_u3_u7_n166 ) , .ZN( u0_u3_u7_n93 ) );
  OAI222_X1 u0_u3_u7_U8 (.C2( u0_u3_u7_n101 ) , .B2( u0_u3_u7_n111 ) , .A1( u0_u3_u7_n113 ) , .C1( u0_u3_u7_n146 ) , .A2( u0_u3_u7_n162 ) , .B1( u0_u3_u7_n164 ) , .ZN( u0_u3_u7_n94 ) );
  INV_X1 u0_u3_u7_U80 (.A( u0_u3_X_46 ) , .ZN( u0_u3_u7_n163 ) );
  INV_X1 u0_u3_u7_U81 (.A( u0_u3_X_43 ) , .ZN( u0_u3_u7_n167 ) );
  INV_X1 u0_u3_u7_U82 (.A( u0_u3_X_45 ) , .ZN( u0_u3_u7_n166 ) );
  NAND4_X1 u0_u3_u7_U83 (.ZN( u0_out3_5 ) , .A4( u0_u3_u7_n108 ) , .A3( u0_u3_u7_n109 ) , .A1( u0_u3_u7_n116 ) , .A2( u0_u3_u7_n123 ) );
  AOI22_X1 u0_u3_u7_U84 (.ZN( u0_u3_u7_n109 ) , .A2( u0_u3_u7_n126 ) , .B2( u0_u3_u7_n145 ) , .B1( u0_u3_u7_n156 ) , .A1( u0_u3_u7_n171 ) );
  NOR4_X1 u0_u3_u7_U85 (.A4( u0_u3_u7_n104 ) , .A3( u0_u3_u7_n105 ) , .A2( u0_u3_u7_n106 ) , .A1( u0_u3_u7_n107 ) , .ZN( u0_u3_u7_n108 ) );
  NAND4_X1 u0_u3_u7_U86 (.ZN( u0_out3_27 ) , .A4( u0_u3_u7_n118 ) , .A3( u0_u3_u7_n119 ) , .A2( u0_u3_u7_n120 ) , .A1( u0_u3_u7_n121 ) );
  OAI21_X1 u0_u3_u7_U87 (.ZN( u0_u3_u7_n121 ) , .B2( u0_u3_u7_n145 ) , .A( u0_u3_u7_n150 ) , .B1( u0_u3_u7_n174 ) );
  OAI21_X1 u0_u3_u7_U88 (.ZN( u0_u3_u7_n120 ) , .A( u0_u3_u7_n161 ) , .B2( u0_u3_u7_n170 ) , .B1( u0_u3_u7_n179 ) );
  NAND4_X1 u0_u3_u7_U89 (.ZN( u0_out3_21 ) , .A4( u0_u3_u7_n157 ) , .A3( u0_u3_u7_n158 ) , .A2( u0_u3_u7_n159 ) , .A1( u0_u3_u7_n160 ) );
  OAI221_X1 u0_u3_u7_U9 (.C1( u0_u3_u7_n101 ) , .C2( u0_u3_u7_n147 ) , .ZN( u0_u3_u7_n155 ) , .B2( u0_u3_u7_n162 ) , .A( u0_u3_u7_n91 ) , .B1( u0_u3_u7_n92 ) );
  OAI21_X1 u0_u3_u7_U90 (.B1( u0_u3_u7_n145 ) , .ZN( u0_u3_u7_n160 ) , .A( u0_u3_u7_n161 ) , .B2( u0_u3_u7_n177 ) );
  AOI22_X1 u0_u3_u7_U91 (.B2( u0_u3_u7_n149 ) , .B1( u0_u3_u7_n150 ) , .A2( u0_u3_u7_n151 ) , .A1( u0_u3_u7_n152 ) , .ZN( u0_u3_u7_n158 ) );
  NAND4_X1 u0_u3_u7_U92 (.ZN( u0_out3_15 ) , .A4( u0_u3_u7_n142 ) , .A3( u0_u3_u7_n143 ) , .A2( u0_u3_u7_n144 ) , .A1( u0_u3_u7_n178 ) );
  OR2_X1 u0_u3_u7_U93 (.A2( u0_u3_u7_n125 ) , .A1( u0_u3_u7_n129 ) , .ZN( u0_u3_u7_n144 ) );
  AOI22_X1 u0_u3_u7_U94 (.A2( u0_u3_u7_n126 ) , .ZN( u0_u3_u7_n143 ) , .B2( u0_u3_u7_n165 ) , .B1( u0_u3_u7_n173 ) , .A1( u0_u3_u7_n174 ) );
  NAND3_X1 u0_u3_u7_U95 (.A3( u0_u3_u7_n146 ) , .A2( u0_u3_u7_n147 ) , .A1( u0_u3_u7_n148 ) , .ZN( u0_u3_u7_n151 ) );
  NAND3_X1 u0_u3_u7_U96 (.A3( u0_u3_u7_n131 ) , .A2( u0_u3_u7_n132 ) , .A1( u0_u3_u7_n133 ) , .ZN( u0_u3_u7_n135 ) );
  XOR2_X1 u0_u5_U1 (.B( u0_K6_9 ) , .A( u0_R4_6 ) , .Z( u0_u5_X_9 ) );
  XOR2_X1 u0_u5_U10 (.B( u0_K6_45 ) , .A( u0_R4_30 ) , .Z( u0_u5_X_45 ) );
  XOR2_X1 u0_u5_U11 (.B( u0_K6_44 ) , .A( u0_R4_29 ) , .Z( u0_u5_X_44 ) );
  XOR2_X1 u0_u5_U12 (.B( u0_K6_43 ) , .A( u0_R4_28 ) , .Z( u0_u5_X_43 ) );
  XOR2_X1 u0_u5_U16 (.B( u0_K6_3 ) , .A( u0_R4_2 ) , .Z( u0_u5_X_3 ) );
  XOR2_X1 u0_u5_U2 (.B( u0_K6_8 ) , .A( u0_R4_5 ) , .Z( u0_u5_X_8 ) );
  XOR2_X1 u0_u5_U20 (.B( u0_K6_36 ) , .A( u0_R4_25 ) , .Z( u0_u5_X_36 ) );
  XOR2_X1 u0_u5_U21 (.B( u0_K6_35 ) , .A( u0_R4_24 ) , .Z( u0_u5_X_35 ) );
  XOR2_X1 u0_u5_U22 (.B( u0_K6_34 ) , .A( u0_R4_23 ) , .Z( u0_u5_X_34 ) );
  XOR2_X1 u0_u5_U23 (.B( u0_K6_33 ) , .A( u0_R4_22 ) , .Z( u0_u5_X_33 ) );
  XOR2_X1 u0_u5_U24 (.B( u0_K6_32 ) , .A( u0_R4_21 ) , .Z( u0_u5_X_32 ) );
  XOR2_X1 u0_u5_U25 (.B( u0_K6_31 ) , .A( u0_R4_20 ) , .Z( u0_u5_X_31 ) );
  XOR2_X1 u0_u5_U27 (.B( u0_K6_2 ) , .A( u0_R4_1 ) , .Z( u0_u5_X_2 ) );
  XOR2_X1 u0_u5_U3 (.B( u0_K6_7 ) , .A( u0_R4_4 ) , .Z( u0_u5_X_7 ) );
  XOR2_X1 u0_u5_U33 (.B( u0_K6_24 ) , .A( u0_R4_17 ) , .Z( u0_u5_X_24 ) );
  XOR2_X1 u0_u5_U34 (.B( u0_K6_23 ) , .A( u0_R4_16 ) , .Z( u0_u5_X_23 ) );
  XOR2_X1 u0_u5_U35 (.B( u0_K6_22 ) , .A( u0_R4_15 ) , .Z( u0_u5_X_22 ) );
  XOR2_X1 u0_u5_U36 (.B( u0_K6_21 ) , .A( u0_R4_14 ) , .Z( u0_u5_X_21 ) );
  XOR2_X1 u0_u5_U37 (.B( u0_K6_20 ) , .A( u0_R4_13 ) , .Z( u0_u5_X_20 ) );
  XOR2_X1 u0_u5_U38 (.B( u0_K6_1 ) , .A( u0_R4_32 ) , .Z( u0_u5_X_1 ) );
  XOR2_X1 u0_u5_U39 (.B( u0_K6_19 ) , .A( u0_R4_12 ) , .Z( u0_u5_X_19 ) );
  XOR2_X1 u0_u5_U4 (.B( u0_K6_6 ) , .A( u0_R4_5 ) , .Z( u0_u5_X_6 ) );
  XOR2_X1 u0_u5_U40 (.B( u0_K6_18 ) , .A( u0_R4_13 ) , .Z( u0_u5_X_18 ) );
  XOR2_X1 u0_u5_U41 (.B( u0_K6_17 ) , .A( u0_R4_12 ) , .Z( u0_u5_X_17 ) );
  XOR2_X1 u0_u5_U42 (.B( u0_K6_16 ) , .A( u0_R4_11 ) , .Z( u0_u5_X_16 ) );
  XOR2_X1 u0_u5_U43 (.B( u0_K6_15 ) , .A( u0_R4_10 ) , .Z( u0_u5_X_15 ) );
  XOR2_X1 u0_u5_U44 (.B( u0_K6_14 ) , .A( u0_R4_9 ) , .Z( u0_u5_X_14 ) );
  XOR2_X1 u0_u5_U45 (.B( u0_K6_13 ) , .A( u0_R4_8 ) , .Z( u0_u5_X_13 ) );
  XOR2_X1 u0_u5_U46 (.B( u0_K6_12 ) , .A( u0_R4_9 ) , .Z( u0_u5_X_12 ) );
  XOR2_X1 u0_u5_U47 (.B( u0_K6_11 ) , .A( u0_R4_8 ) , .Z( u0_u5_X_11 ) );
  XOR2_X1 u0_u5_U48 (.B( u0_K6_10 ) , .A( u0_R4_7 ) , .Z( u0_u5_X_10 ) );
  XOR2_X1 u0_u5_U5 (.B( u0_K6_5 ) , .A( u0_R4_4 ) , .Z( u0_u5_X_5 ) );
  XOR2_X1 u0_u5_U6 (.B( u0_K6_4 ) , .A( u0_R4_3 ) , .Z( u0_u5_X_4 ) );
  XOR2_X1 u0_u5_U7 (.B( u0_K6_48 ) , .A( u0_R4_1 ) , .Z( u0_u5_X_48 ) );
  XOR2_X1 u0_u5_U8 (.B( u0_K6_47 ) , .A( u0_R4_32 ) , .Z( u0_u5_X_47 ) );
  XOR2_X1 u0_u5_U9 (.B( u0_K6_46 ) , .A( u0_R4_31 ) , .Z( u0_u5_X_46 ) );
  AND2_X1 u0_u5_u0_U10 (.A1( u0_u5_u0_n131 ) , .ZN( u0_u5_u0_n141 ) , .A2( u0_u5_u0_n150 ) );
  AND3_X1 u0_u5_u0_U11 (.A2( u0_u5_u0_n112 ) , .ZN( u0_u5_u0_n127 ) , .A3( u0_u5_u0_n130 ) , .A1( u0_u5_u0_n148 ) );
  AND2_X1 u0_u5_u0_U12 (.ZN( u0_u5_u0_n107 ) , .A1( u0_u5_u0_n130 ) , .A2( u0_u5_u0_n140 ) );
  AND2_X1 u0_u5_u0_U13 (.A2( u0_u5_u0_n129 ) , .A1( u0_u5_u0_n130 ) , .ZN( u0_u5_u0_n151 ) );
  AND2_X1 u0_u5_u0_U14 (.A1( u0_u5_u0_n108 ) , .A2( u0_u5_u0_n125 ) , .ZN( u0_u5_u0_n145 ) );
  INV_X1 u0_u5_u0_U15 (.A( u0_u5_u0_n143 ) , .ZN( u0_u5_u0_n173 ) );
  NOR2_X1 u0_u5_u0_U16 (.A2( u0_u5_u0_n136 ) , .ZN( u0_u5_u0_n147 ) , .A1( u0_u5_u0_n160 ) );
  AOI21_X1 u0_u5_u0_U17 (.B1( u0_u5_u0_n103 ) , .ZN( u0_u5_u0_n132 ) , .A( u0_u5_u0_n165 ) , .B2( u0_u5_u0_n93 ) );
  OAI22_X1 u0_u5_u0_U18 (.B1( u0_u5_u0_n131 ) , .A1( u0_u5_u0_n144 ) , .B2( u0_u5_u0_n147 ) , .A2( u0_u5_u0_n90 ) , .ZN( u0_u5_u0_n91 ) );
  AND3_X1 u0_u5_u0_U19 (.A3( u0_u5_u0_n121 ) , .A2( u0_u5_u0_n125 ) , .A1( u0_u5_u0_n148 ) , .ZN( u0_u5_u0_n90 ) );
  OAI22_X1 u0_u5_u0_U20 (.B1( u0_u5_u0_n125 ) , .ZN( u0_u5_u0_n126 ) , .A1( u0_u5_u0_n138 ) , .A2( u0_u5_u0_n146 ) , .B2( u0_u5_u0_n147 ) );
  NOR2_X1 u0_u5_u0_U21 (.A1( u0_u5_u0_n163 ) , .A2( u0_u5_u0_n164 ) , .ZN( u0_u5_u0_n95 ) );
  AOI22_X1 u0_u5_u0_U22 (.B2( u0_u5_u0_n109 ) , .A2( u0_u5_u0_n110 ) , .ZN( u0_u5_u0_n111 ) , .B1( u0_u5_u0_n118 ) , .A1( u0_u5_u0_n160 ) );
  NAND2_X1 u0_u5_u0_U23 (.A2( u0_u5_u0_n102 ) , .A1( u0_u5_u0_n103 ) , .ZN( u0_u5_u0_n149 ) );
  INV_X1 u0_u5_u0_U24 (.A( u0_u5_u0_n136 ) , .ZN( u0_u5_u0_n161 ) );
  INV_X1 u0_u5_u0_U25 (.A( u0_u5_u0_n118 ) , .ZN( u0_u5_u0_n158 ) );
  NAND2_X1 u0_u5_u0_U26 (.A2( u0_u5_u0_n100 ) , .ZN( u0_u5_u0_n131 ) , .A1( u0_u5_u0_n92 ) );
  NAND2_X1 u0_u5_u0_U27 (.ZN( u0_u5_u0_n108 ) , .A1( u0_u5_u0_n92 ) , .A2( u0_u5_u0_n94 ) );
  AOI21_X1 u0_u5_u0_U28 (.ZN( u0_u5_u0_n104 ) , .B1( u0_u5_u0_n107 ) , .B2( u0_u5_u0_n141 ) , .A( u0_u5_u0_n144 ) );
  AOI21_X1 u0_u5_u0_U29 (.B1( u0_u5_u0_n127 ) , .B2( u0_u5_u0_n129 ) , .A( u0_u5_u0_n138 ) , .ZN( u0_u5_u0_n96 ) );
  INV_X1 u0_u5_u0_U3 (.A( u0_u5_u0_n113 ) , .ZN( u0_u5_u0_n166 ) );
  NAND2_X1 u0_u5_u0_U30 (.A2( u0_u5_u0_n102 ) , .ZN( u0_u5_u0_n114 ) , .A1( u0_u5_u0_n92 ) );
  NOR2_X1 u0_u5_u0_U31 (.A1( u0_u5_u0_n120 ) , .ZN( u0_u5_u0_n143 ) , .A2( u0_u5_u0_n167 ) );
  OAI221_X1 u0_u5_u0_U32 (.C1( u0_u5_u0_n112 ) , .ZN( u0_u5_u0_n120 ) , .B1( u0_u5_u0_n138 ) , .B2( u0_u5_u0_n141 ) , .C2( u0_u5_u0_n147 ) , .A( u0_u5_u0_n172 ) );
  AOI211_X1 u0_u5_u0_U33 (.B( u0_u5_u0_n115 ) , .A( u0_u5_u0_n116 ) , .C2( u0_u5_u0_n117 ) , .C1( u0_u5_u0_n118 ) , .ZN( u0_u5_u0_n119 ) );
  NAND2_X1 u0_u5_u0_U34 (.A2( u0_u5_u0_n103 ) , .ZN( u0_u5_u0_n140 ) , .A1( u0_u5_u0_n94 ) );
  NAND2_X1 u0_u5_u0_U35 (.A1( u0_u5_u0_n100 ) , .A2( u0_u5_u0_n103 ) , .ZN( u0_u5_u0_n125 ) );
  NAND2_X1 u0_u5_u0_U36 (.A1( u0_u5_u0_n101 ) , .A2( u0_u5_u0_n102 ) , .ZN( u0_u5_u0_n150 ) );
  INV_X1 u0_u5_u0_U37 (.A( u0_u5_u0_n138 ) , .ZN( u0_u5_u0_n160 ) );
  NAND2_X1 u0_u5_u0_U38 (.A2( u0_u5_u0_n100 ) , .A1( u0_u5_u0_n101 ) , .ZN( u0_u5_u0_n139 ) );
  NAND2_X1 u0_u5_u0_U39 (.ZN( u0_u5_u0_n112 ) , .A2( u0_u5_u0_n92 ) , .A1( u0_u5_u0_n93 ) );
  AOI21_X1 u0_u5_u0_U4 (.B1( u0_u5_u0_n114 ) , .ZN( u0_u5_u0_n115 ) , .B2( u0_u5_u0_n129 ) , .A( u0_u5_u0_n161 ) );
  NAND2_X1 u0_u5_u0_U40 (.A1( u0_u5_u0_n101 ) , .ZN( u0_u5_u0_n130 ) , .A2( u0_u5_u0_n94 ) );
  INV_X1 u0_u5_u0_U41 (.ZN( u0_u5_u0_n172 ) , .A( u0_u5_u0_n88 ) );
  OAI222_X1 u0_u5_u0_U42 (.C1( u0_u5_u0_n108 ) , .A1( u0_u5_u0_n125 ) , .B2( u0_u5_u0_n128 ) , .B1( u0_u5_u0_n144 ) , .A2( u0_u5_u0_n158 ) , .C2( u0_u5_u0_n161 ) , .ZN( u0_u5_u0_n88 ) );
  NAND2_X1 u0_u5_u0_U43 (.A2( u0_u5_u0_n101 ) , .ZN( u0_u5_u0_n121 ) , .A1( u0_u5_u0_n93 ) );
  OR3_X1 u0_u5_u0_U44 (.A3( u0_u5_u0_n152 ) , .A2( u0_u5_u0_n153 ) , .A1( u0_u5_u0_n154 ) , .ZN( u0_u5_u0_n155 ) );
  AOI21_X1 u0_u5_u0_U45 (.A( u0_u5_u0_n144 ) , .B2( u0_u5_u0_n145 ) , .B1( u0_u5_u0_n146 ) , .ZN( u0_u5_u0_n154 ) );
  AOI21_X1 u0_u5_u0_U46 (.B2( u0_u5_u0_n150 ) , .B1( u0_u5_u0_n151 ) , .ZN( u0_u5_u0_n152 ) , .A( u0_u5_u0_n158 ) );
  AOI21_X1 u0_u5_u0_U47 (.A( u0_u5_u0_n147 ) , .B2( u0_u5_u0_n148 ) , .B1( u0_u5_u0_n149 ) , .ZN( u0_u5_u0_n153 ) );
  INV_X1 u0_u5_u0_U48 (.ZN( u0_u5_u0_n171 ) , .A( u0_u5_u0_n99 ) );
  OAI211_X1 u0_u5_u0_U49 (.C2( u0_u5_u0_n140 ) , .C1( u0_u5_u0_n161 ) , .A( u0_u5_u0_n169 ) , .B( u0_u5_u0_n98 ) , .ZN( u0_u5_u0_n99 ) );
  AOI21_X1 u0_u5_u0_U5 (.B2( u0_u5_u0_n131 ) , .ZN( u0_u5_u0_n134 ) , .B1( u0_u5_u0_n151 ) , .A( u0_u5_u0_n158 ) );
  AOI211_X1 u0_u5_u0_U50 (.C1( u0_u5_u0_n118 ) , .A( u0_u5_u0_n123 ) , .B( u0_u5_u0_n96 ) , .C2( u0_u5_u0_n97 ) , .ZN( u0_u5_u0_n98 ) );
  INV_X1 u0_u5_u0_U51 (.ZN( u0_u5_u0_n169 ) , .A( u0_u5_u0_n91 ) );
  NOR2_X1 u0_u5_u0_U52 (.A2( u0_u5_X_4 ) , .A1( u0_u5_X_5 ) , .ZN( u0_u5_u0_n118 ) );
  NOR2_X1 u0_u5_u0_U53 (.A2( u0_u5_X_1 ) , .ZN( u0_u5_u0_n101 ) , .A1( u0_u5_u0_n163 ) );
  NOR2_X1 u0_u5_u0_U54 (.A2( u0_u5_X_3 ) , .A1( u0_u5_X_6 ) , .ZN( u0_u5_u0_n94 ) );
  NOR2_X1 u0_u5_u0_U55 (.A2( u0_u5_X_6 ) , .ZN( u0_u5_u0_n100 ) , .A1( u0_u5_u0_n162 ) );
  NAND2_X1 u0_u5_u0_U56 (.A2( u0_u5_X_4 ) , .A1( u0_u5_X_5 ) , .ZN( u0_u5_u0_n144 ) );
  NOR2_X1 u0_u5_u0_U57 (.A2( u0_u5_X_5 ) , .ZN( u0_u5_u0_n136 ) , .A1( u0_u5_u0_n159 ) );
  NAND2_X1 u0_u5_u0_U58 (.A1( u0_u5_X_5 ) , .ZN( u0_u5_u0_n138 ) , .A2( u0_u5_u0_n159 ) );
  AND2_X1 u0_u5_u0_U59 (.A2( u0_u5_X_3 ) , .A1( u0_u5_X_6 ) , .ZN( u0_u5_u0_n102 ) );
  NOR2_X1 u0_u5_u0_U6 (.A1( u0_u5_u0_n108 ) , .ZN( u0_u5_u0_n123 ) , .A2( u0_u5_u0_n158 ) );
  AND2_X1 u0_u5_u0_U60 (.A1( u0_u5_X_6 ) , .A2( u0_u5_u0_n162 ) , .ZN( u0_u5_u0_n93 ) );
  INV_X1 u0_u5_u0_U61 (.A( u0_u5_X_4 ) , .ZN( u0_u5_u0_n159 ) );
  INV_X1 u0_u5_u0_U62 (.A( u0_u5_X_1 ) , .ZN( u0_u5_u0_n164 ) );
  INV_X1 u0_u5_u0_U63 (.A( u0_u5_X_3 ) , .ZN( u0_u5_u0_n162 ) );
  AOI211_X1 u0_u5_u0_U64 (.B( u0_u5_u0_n133 ) , .A( u0_u5_u0_n134 ) , .C2( u0_u5_u0_n135 ) , .C1( u0_u5_u0_n136 ) , .ZN( u0_u5_u0_n137 ) );
  INV_X1 u0_u5_u0_U65 (.A( u0_u5_u0_n126 ) , .ZN( u0_u5_u0_n168 ) );
  OR4_X1 u0_u5_u0_U66 (.ZN( u0_out5_17 ) , .A4( u0_u5_u0_n122 ) , .A2( u0_u5_u0_n123 ) , .A1( u0_u5_u0_n124 ) , .A3( u0_u5_u0_n170 ) );
  AOI21_X1 u0_u5_u0_U67 (.B2( u0_u5_u0_n107 ) , .ZN( u0_u5_u0_n124 ) , .B1( u0_u5_u0_n128 ) , .A( u0_u5_u0_n161 ) );
  INV_X1 u0_u5_u0_U68 (.A( u0_u5_u0_n111 ) , .ZN( u0_u5_u0_n170 ) );
  OR4_X1 u0_u5_u0_U69 (.ZN( u0_out5_31 ) , .A4( u0_u5_u0_n155 ) , .A2( u0_u5_u0_n156 ) , .A1( u0_u5_u0_n157 ) , .A3( u0_u5_u0_n173 ) );
  OAI21_X1 u0_u5_u0_U7 (.B1( u0_u5_u0_n150 ) , .B2( u0_u5_u0_n158 ) , .A( u0_u5_u0_n172 ) , .ZN( u0_u5_u0_n89 ) );
  AOI21_X1 u0_u5_u0_U70 (.A( u0_u5_u0_n138 ) , .B2( u0_u5_u0_n139 ) , .B1( u0_u5_u0_n140 ) , .ZN( u0_u5_u0_n157 ) );
  INV_X1 u0_u5_u0_U71 (.ZN( u0_u5_u0_n174 ) , .A( u0_u5_u0_n89 ) );
  AOI211_X1 u0_u5_u0_U72 (.B( u0_u5_u0_n104 ) , .A( u0_u5_u0_n105 ) , .ZN( u0_u5_u0_n106 ) , .C2( u0_u5_u0_n113 ) , .C1( u0_u5_u0_n160 ) );
  INV_X1 u0_u5_u0_U73 (.A( u0_u5_u0_n142 ) , .ZN( u0_u5_u0_n165 ) );
  AOI21_X1 u0_u5_u0_U74 (.ZN( u0_u5_u0_n116 ) , .B2( u0_u5_u0_n142 ) , .A( u0_u5_u0_n144 ) , .B1( u0_u5_u0_n166 ) );
  AOI21_X1 u0_u5_u0_U75 (.B2( u0_u5_u0_n141 ) , .B1( u0_u5_u0_n142 ) , .ZN( u0_u5_u0_n156 ) , .A( u0_u5_u0_n161 ) );
  OAI221_X1 u0_u5_u0_U76 (.C1( u0_u5_u0_n121 ) , .ZN( u0_u5_u0_n122 ) , .B2( u0_u5_u0_n127 ) , .A( u0_u5_u0_n143 ) , .B1( u0_u5_u0_n144 ) , .C2( u0_u5_u0_n147 ) );
  AOI21_X1 u0_u5_u0_U77 (.B1( u0_u5_u0_n132 ) , .ZN( u0_u5_u0_n133 ) , .A( u0_u5_u0_n144 ) , .B2( u0_u5_u0_n166 ) );
  OAI22_X1 u0_u5_u0_U78 (.ZN( u0_u5_u0_n105 ) , .A2( u0_u5_u0_n132 ) , .B1( u0_u5_u0_n146 ) , .A1( u0_u5_u0_n147 ) , .B2( u0_u5_u0_n161 ) );
  NAND2_X1 u0_u5_u0_U79 (.ZN( u0_u5_u0_n110 ) , .A2( u0_u5_u0_n132 ) , .A1( u0_u5_u0_n145 ) );
  AND2_X1 u0_u5_u0_U8 (.A1( u0_u5_u0_n114 ) , .A2( u0_u5_u0_n121 ) , .ZN( u0_u5_u0_n146 ) );
  INV_X1 u0_u5_u0_U80 (.A( u0_u5_u0_n119 ) , .ZN( u0_u5_u0_n167 ) );
  NAND2_X1 u0_u5_u0_U81 (.ZN( u0_u5_u0_n148 ) , .A1( u0_u5_u0_n93 ) , .A2( u0_u5_u0_n95 ) );
  NAND2_X1 u0_u5_u0_U82 (.A1( u0_u5_u0_n100 ) , .ZN( u0_u5_u0_n129 ) , .A2( u0_u5_u0_n95 ) );
  NAND2_X1 u0_u5_u0_U83 (.A1( u0_u5_u0_n102 ) , .ZN( u0_u5_u0_n128 ) , .A2( u0_u5_u0_n95 ) );
  NOR2_X1 u0_u5_u0_U84 (.A2( u0_u5_X_1 ) , .A1( u0_u5_X_2 ) , .ZN( u0_u5_u0_n92 ) );
  NAND2_X1 u0_u5_u0_U85 (.ZN( u0_u5_u0_n142 ) , .A1( u0_u5_u0_n94 ) , .A2( u0_u5_u0_n95 ) );
  NOR2_X1 u0_u5_u0_U86 (.A2( u0_u5_X_2 ) , .ZN( u0_u5_u0_n103 ) , .A1( u0_u5_u0_n164 ) );
  INV_X1 u0_u5_u0_U87 (.A( u0_u5_X_2 ) , .ZN( u0_u5_u0_n163 ) );
  NAND3_X1 u0_u5_u0_U88 (.ZN( u0_out5_23 ) , .A3( u0_u5_u0_n137 ) , .A1( u0_u5_u0_n168 ) , .A2( u0_u5_u0_n171 ) );
  NAND3_X1 u0_u5_u0_U89 (.A3( u0_u5_u0_n127 ) , .A2( u0_u5_u0_n128 ) , .ZN( u0_u5_u0_n135 ) , .A1( u0_u5_u0_n150 ) );
  NAND2_X1 u0_u5_u0_U9 (.ZN( u0_u5_u0_n113 ) , .A1( u0_u5_u0_n139 ) , .A2( u0_u5_u0_n149 ) );
  NAND3_X1 u0_u5_u0_U90 (.ZN( u0_u5_u0_n117 ) , .A3( u0_u5_u0_n132 ) , .A2( u0_u5_u0_n139 ) , .A1( u0_u5_u0_n148 ) );
  NAND3_X1 u0_u5_u0_U91 (.ZN( u0_u5_u0_n109 ) , .A2( u0_u5_u0_n114 ) , .A3( u0_u5_u0_n140 ) , .A1( u0_u5_u0_n149 ) );
  NAND3_X1 u0_u5_u0_U92 (.ZN( u0_out5_9 ) , .A3( u0_u5_u0_n106 ) , .A2( u0_u5_u0_n171 ) , .A1( u0_u5_u0_n174 ) );
  NAND3_X1 u0_u5_u0_U93 (.A2( u0_u5_u0_n128 ) , .A1( u0_u5_u0_n132 ) , .A3( u0_u5_u0_n146 ) , .ZN( u0_u5_u0_n97 ) );
  NOR2_X1 u0_u5_u1_U10 (.A1( u0_u5_u1_n112 ) , .A2( u0_u5_u1_n116 ) , .ZN( u0_u5_u1_n118 ) );
  NAND3_X1 u0_u5_u1_U100 (.ZN( u0_u5_u1_n113 ) , .A1( u0_u5_u1_n120 ) , .A3( u0_u5_u1_n133 ) , .A2( u0_u5_u1_n155 ) );
  OAI21_X1 u0_u5_u1_U11 (.ZN( u0_u5_u1_n101 ) , .B1( u0_u5_u1_n141 ) , .A( u0_u5_u1_n146 ) , .B2( u0_u5_u1_n183 ) );
  AOI21_X1 u0_u5_u1_U12 (.B2( u0_u5_u1_n155 ) , .B1( u0_u5_u1_n156 ) , .ZN( u0_u5_u1_n157 ) , .A( u0_u5_u1_n174 ) );
  NAND2_X1 u0_u5_u1_U13 (.ZN( u0_u5_u1_n140 ) , .A2( u0_u5_u1_n150 ) , .A1( u0_u5_u1_n155 ) );
  NAND2_X1 u0_u5_u1_U14 (.A1( u0_u5_u1_n131 ) , .ZN( u0_u5_u1_n147 ) , .A2( u0_u5_u1_n153 ) );
  INV_X1 u0_u5_u1_U15 (.A( u0_u5_u1_n139 ) , .ZN( u0_u5_u1_n174 ) );
  OR4_X1 u0_u5_u1_U16 (.A4( u0_u5_u1_n106 ) , .A3( u0_u5_u1_n107 ) , .ZN( u0_u5_u1_n108 ) , .A1( u0_u5_u1_n117 ) , .A2( u0_u5_u1_n184 ) );
  AOI21_X1 u0_u5_u1_U17 (.ZN( u0_u5_u1_n106 ) , .A( u0_u5_u1_n112 ) , .B1( u0_u5_u1_n154 ) , .B2( u0_u5_u1_n156 ) );
  INV_X1 u0_u5_u1_U18 (.A( u0_u5_u1_n101 ) , .ZN( u0_u5_u1_n184 ) );
  AOI21_X1 u0_u5_u1_U19 (.ZN( u0_u5_u1_n107 ) , .B1( u0_u5_u1_n134 ) , .B2( u0_u5_u1_n149 ) , .A( u0_u5_u1_n174 ) );
  INV_X1 u0_u5_u1_U20 (.A( u0_u5_u1_n112 ) , .ZN( u0_u5_u1_n171 ) );
  NAND2_X1 u0_u5_u1_U21 (.ZN( u0_u5_u1_n141 ) , .A1( u0_u5_u1_n153 ) , .A2( u0_u5_u1_n156 ) );
  AND2_X1 u0_u5_u1_U22 (.A1( u0_u5_u1_n123 ) , .ZN( u0_u5_u1_n134 ) , .A2( u0_u5_u1_n161 ) );
  NAND2_X1 u0_u5_u1_U23 (.A2( u0_u5_u1_n115 ) , .A1( u0_u5_u1_n116 ) , .ZN( u0_u5_u1_n148 ) );
  NAND2_X1 u0_u5_u1_U24 (.A2( u0_u5_u1_n133 ) , .A1( u0_u5_u1_n135 ) , .ZN( u0_u5_u1_n159 ) );
  NAND2_X1 u0_u5_u1_U25 (.A2( u0_u5_u1_n115 ) , .A1( u0_u5_u1_n120 ) , .ZN( u0_u5_u1_n132 ) );
  INV_X1 u0_u5_u1_U26 (.A( u0_u5_u1_n154 ) , .ZN( u0_u5_u1_n178 ) );
  INV_X1 u0_u5_u1_U27 (.A( u0_u5_u1_n151 ) , .ZN( u0_u5_u1_n183 ) );
  AND2_X1 u0_u5_u1_U28 (.A1( u0_u5_u1_n129 ) , .A2( u0_u5_u1_n133 ) , .ZN( u0_u5_u1_n149 ) );
  INV_X1 u0_u5_u1_U29 (.A( u0_u5_u1_n131 ) , .ZN( u0_u5_u1_n180 ) );
  INV_X1 u0_u5_u1_U3 (.A( u0_u5_u1_n159 ) , .ZN( u0_u5_u1_n182 ) );
  OAI221_X1 u0_u5_u1_U30 (.A( u0_u5_u1_n119 ) , .C2( u0_u5_u1_n129 ) , .ZN( u0_u5_u1_n138 ) , .B2( u0_u5_u1_n152 ) , .C1( u0_u5_u1_n174 ) , .B1( u0_u5_u1_n187 ) );
  INV_X1 u0_u5_u1_U31 (.A( u0_u5_u1_n148 ) , .ZN( u0_u5_u1_n187 ) );
  AOI211_X1 u0_u5_u1_U32 (.B( u0_u5_u1_n117 ) , .A( u0_u5_u1_n118 ) , .ZN( u0_u5_u1_n119 ) , .C2( u0_u5_u1_n146 ) , .C1( u0_u5_u1_n159 ) );
  NOR2_X1 u0_u5_u1_U33 (.A1( u0_u5_u1_n168 ) , .A2( u0_u5_u1_n176 ) , .ZN( u0_u5_u1_n98 ) );
  OAI21_X1 u0_u5_u1_U34 (.B2( u0_u5_u1_n123 ) , .ZN( u0_u5_u1_n145 ) , .B1( u0_u5_u1_n160 ) , .A( u0_u5_u1_n185 ) );
  INV_X1 u0_u5_u1_U35 (.A( u0_u5_u1_n122 ) , .ZN( u0_u5_u1_n185 ) );
  AOI21_X1 u0_u5_u1_U36 (.B2( u0_u5_u1_n120 ) , .B1( u0_u5_u1_n121 ) , .ZN( u0_u5_u1_n122 ) , .A( u0_u5_u1_n128 ) );
  NAND2_X1 u0_u5_u1_U37 (.A1( u0_u5_u1_n128 ) , .ZN( u0_u5_u1_n146 ) , .A2( u0_u5_u1_n160 ) );
  NAND2_X1 u0_u5_u1_U38 (.A2( u0_u5_u1_n112 ) , .ZN( u0_u5_u1_n139 ) , .A1( u0_u5_u1_n152 ) );
  NAND2_X1 u0_u5_u1_U39 (.A1( u0_u5_u1_n105 ) , .ZN( u0_u5_u1_n156 ) , .A2( u0_u5_u1_n99 ) );
  AOI221_X1 u0_u5_u1_U4 (.A( u0_u5_u1_n138 ) , .C2( u0_u5_u1_n139 ) , .C1( u0_u5_u1_n140 ) , .B2( u0_u5_u1_n141 ) , .ZN( u0_u5_u1_n142 ) , .B1( u0_u5_u1_n175 ) );
  AOI221_X1 u0_u5_u1_U40 (.B1( u0_u5_u1_n140 ) , .ZN( u0_u5_u1_n167 ) , .B2( u0_u5_u1_n172 ) , .C2( u0_u5_u1_n175 ) , .C1( u0_u5_u1_n178 ) , .A( u0_u5_u1_n188 ) );
  INV_X1 u0_u5_u1_U41 (.ZN( u0_u5_u1_n188 ) , .A( u0_u5_u1_n97 ) );
  AOI211_X1 u0_u5_u1_U42 (.A( u0_u5_u1_n118 ) , .C1( u0_u5_u1_n132 ) , .C2( u0_u5_u1_n139 ) , .B( u0_u5_u1_n96 ) , .ZN( u0_u5_u1_n97 ) );
  AOI21_X1 u0_u5_u1_U43 (.B2( u0_u5_u1_n121 ) , .B1( u0_u5_u1_n135 ) , .A( u0_u5_u1_n152 ) , .ZN( u0_u5_u1_n96 ) );
  NOR2_X1 u0_u5_u1_U44 (.ZN( u0_u5_u1_n117 ) , .A1( u0_u5_u1_n121 ) , .A2( u0_u5_u1_n160 ) );
  AOI21_X1 u0_u5_u1_U45 (.A( u0_u5_u1_n128 ) , .B2( u0_u5_u1_n129 ) , .ZN( u0_u5_u1_n130 ) , .B1( u0_u5_u1_n150 ) );
  NAND2_X1 u0_u5_u1_U46 (.ZN( u0_u5_u1_n112 ) , .A1( u0_u5_u1_n169 ) , .A2( u0_u5_u1_n170 ) );
  NAND2_X1 u0_u5_u1_U47 (.ZN( u0_u5_u1_n129 ) , .A2( u0_u5_u1_n95 ) , .A1( u0_u5_u1_n98 ) );
  NAND2_X1 u0_u5_u1_U48 (.A1( u0_u5_u1_n102 ) , .ZN( u0_u5_u1_n154 ) , .A2( u0_u5_u1_n99 ) );
  NAND2_X1 u0_u5_u1_U49 (.A2( u0_u5_u1_n100 ) , .ZN( u0_u5_u1_n135 ) , .A1( u0_u5_u1_n99 ) );
  AOI211_X1 u0_u5_u1_U5 (.ZN( u0_u5_u1_n124 ) , .A( u0_u5_u1_n138 ) , .C2( u0_u5_u1_n139 ) , .B( u0_u5_u1_n145 ) , .C1( u0_u5_u1_n147 ) );
  AOI21_X1 u0_u5_u1_U50 (.A( u0_u5_u1_n152 ) , .B2( u0_u5_u1_n153 ) , .B1( u0_u5_u1_n154 ) , .ZN( u0_u5_u1_n158 ) );
  INV_X1 u0_u5_u1_U51 (.A( u0_u5_u1_n160 ) , .ZN( u0_u5_u1_n175 ) );
  NAND2_X1 u0_u5_u1_U52 (.A1( u0_u5_u1_n100 ) , .ZN( u0_u5_u1_n116 ) , .A2( u0_u5_u1_n95 ) );
  NAND2_X1 u0_u5_u1_U53 (.A1( u0_u5_u1_n102 ) , .ZN( u0_u5_u1_n131 ) , .A2( u0_u5_u1_n95 ) );
  NAND2_X1 u0_u5_u1_U54 (.A2( u0_u5_u1_n104 ) , .ZN( u0_u5_u1_n121 ) , .A1( u0_u5_u1_n98 ) );
  NAND2_X1 u0_u5_u1_U55 (.A1( u0_u5_u1_n103 ) , .ZN( u0_u5_u1_n153 ) , .A2( u0_u5_u1_n98 ) );
  NAND2_X1 u0_u5_u1_U56 (.A2( u0_u5_u1_n104 ) , .A1( u0_u5_u1_n105 ) , .ZN( u0_u5_u1_n133 ) );
  NAND2_X1 u0_u5_u1_U57 (.ZN( u0_u5_u1_n150 ) , .A2( u0_u5_u1_n98 ) , .A1( u0_u5_u1_n99 ) );
  NAND2_X1 u0_u5_u1_U58 (.A1( u0_u5_u1_n105 ) , .ZN( u0_u5_u1_n155 ) , .A2( u0_u5_u1_n95 ) );
  OAI21_X1 u0_u5_u1_U59 (.ZN( u0_u5_u1_n109 ) , .B1( u0_u5_u1_n129 ) , .B2( u0_u5_u1_n160 ) , .A( u0_u5_u1_n167 ) );
  AOI22_X1 u0_u5_u1_U6 (.B2( u0_u5_u1_n136 ) , .A2( u0_u5_u1_n137 ) , .ZN( u0_u5_u1_n143 ) , .A1( u0_u5_u1_n171 ) , .B1( u0_u5_u1_n173 ) );
  NAND2_X1 u0_u5_u1_U60 (.A2( u0_u5_u1_n100 ) , .A1( u0_u5_u1_n103 ) , .ZN( u0_u5_u1_n120 ) );
  NAND2_X1 u0_u5_u1_U61 (.A1( u0_u5_u1_n102 ) , .A2( u0_u5_u1_n104 ) , .ZN( u0_u5_u1_n115 ) );
  NAND2_X1 u0_u5_u1_U62 (.A2( u0_u5_u1_n100 ) , .A1( u0_u5_u1_n104 ) , .ZN( u0_u5_u1_n151 ) );
  NAND2_X1 u0_u5_u1_U63 (.A2( u0_u5_u1_n103 ) , .A1( u0_u5_u1_n105 ) , .ZN( u0_u5_u1_n161 ) );
  INV_X1 u0_u5_u1_U64 (.A( u0_u5_u1_n152 ) , .ZN( u0_u5_u1_n173 ) );
  INV_X1 u0_u5_u1_U65 (.A( u0_u5_u1_n128 ) , .ZN( u0_u5_u1_n172 ) );
  NAND2_X1 u0_u5_u1_U66 (.A2( u0_u5_u1_n102 ) , .A1( u0_u5_u1_n103 ) , .ZN( u0_u5_u1_n123 ) );
  AOI211_X1 u0_u5_u1_U67 (.B( u0_u5_u1_n162 ) , .A( u0_u5_u1_n163 ) , .C2( u0_u5_u1_n164 ) , .ZN( u0_u5_u1_n165 ) , .C1( u0_u5_u1_n171 ) );
  AOI21_X1 u0_u5_u1_U68 (.A( u0_u5_u1_n160 ) , .B2( u0_u5_u1_n161 ) , .ZN( u0_u5_u1_n162 ) , .B1( u0_u5_u1_n182 ) );
  OR2_X1 u0_u5_u1_U69 (.A2( u0_u5_u1_n157 ) , .A1( u0_u5_u1_n158 ) , .ZN( u0_u5_u1_n163 ) );
  INV_X1 u0_u5_u1_U7 (.A( u0_u5_u1_n147 ) , .ZN( u0_u5_u1_n181 ) );
  NOR2_X1 u0_u5_u1_U70 (.A2( u0_u5_X_7 ) , .A1( u0_u5_X_8 ) , .ZN( u0_u5_u1_n95 ) );
  NOR2_X1 u0_u5_u1_U71 (.A1( u0_u5_X_12 ) , .A2( u0_u5_X_9 ) , .ZN( u0_u5_u1_n100 ) );
  NOR2_X1 u0_u5_u1_U72 (.A2( u0_u5_X_8 ) , .A1( u0_u5_u1_n177 ) , .ZN( u0_u5_u1_n99 ) );
  NOR2_X1 u0_u5_u1_U73 (.A2( u0_u5_X_12 ) , .ZN( u0_u5_u1_n102 ) , .A1( u0_u5_u1_n176 ) );
  NOR2_X1 u0_u5_u1_U74 (.A2( u0_u5_X_9 ) , .ZN( u0_u5_u1_n105 ) , .A1( u0_u5_u1_n168 ) );
  NAND2_X1 u0_u5_u1_U75 (.A1( u0_u5_X_10 ) , .ZN( u0_u5_u1_n160 ) , .A2( u0_u5_u1_n169 ) );
  NAND2_X1 u0_u5_u1_U76 (.A2( u0_u5_X_10 ) , .A1( u0_u5_X_11 ) , .ZN( u0_u5_u1_n152 ) );
  NAND2_X1 u0_u5_u1_U77 (.A1( u0_u5_X_11 ) , .ZN( u0_u5_u1_n128 ) , .A2( u0_u5_u1_n170 ) );
  AND2_X1 u0_u5_u1_U78 (.A2( u0_u5_X_7 ) , .A1( u0_u5_X_8 ) , .ZN( u0_u5_u1_n104 ) );
  AND2_X1 u0_u5_u1_U79 (.A1( u0_u5_X_8 ) , .ZN( u0_u5_u1_n103 ) , .A2( u0_u5_u1_n177 ) );
  AOI22_X1 u0_u5_u1_U8 (.B2( u0_u5_u1_n113 ) , .A2( u0_u5_u1_n114 ) , .ZN( u0_u5_u1_n125 ) , .A1( u0_u5_u1_n171 ) , .B1( u0_u5_u1_n173 ) );
  INV_X1 u0_u5_u1_U80 (.A( u0_u5_X_10 ) , .ZN( u0_u5_u1_n170 ) );
  INV_X1 u0_u5_u1_U81 (.A( u0_u5_X_9 ) , .ZN( u0_u5_u1_n176 ) );
  INV_X1 u0_u5_u1_U82 (.A( u0_u5_X_11 ) , .ZN( u0_u5_u1_n169 ) );
  INV_X1 u0_u5_u1_U83 (.A( u0_u5_X_12 ) , .ZN( u0_u5_u1_n168 ) );
  INV_X1 u0_u5_u1_U84 (.A( u0_u5_X_7 ) , .ZN( u0_u5_u1_n177 ) );
  NAND4_X1 u0_u5_u1_U85 (.ZN( u0_out5_28 ) , .A4( u0_u5_u1_n124 ) , .A3( u0_u5_u1_n125 ) , .A2( u0_u5_u1_n126 ) , .A1( u0_u5_u1_n127 ) );
  OAI21_X1 u0_u5_u1_U86 (.ZN( u0_u5_u1_n127 ) , .B2( u0_u5_u1_n139 ) , .B1( u0_u5_u1_n175 ) , .A( u0_u5_u1_n183 ) );
  OAI21_X1 u0_u5_u1_U87 (.ZN( u0_u5_u1_n126 ) , .B2( u0_u5_u1_n140 ) , .A( u0_u5_u1_n146 ) , .B1( u0_u5_u1_n178 ) );
  NAND4_X1 u0_u5_u1_U88 (.ZN( u0_out5_18 ) , .A4( u0_u5_u1_n165 ) , .A3( u0_u5_u1_n166 ) , .A1( u0_u5_u1_n167 ) , .A2( u0_u5_u1_n186 ) );
  AOI22_X1 u0_u5_u1_U89 (.B2( u0_u5_u1_n146 ) , .B1( u0_u5_u1_n147 ) , .A2( u0_u5_u1_n148 ) , .ZN( u0_u5_u1_n166 ) , .A1( u0_u5_u1_n172 ) );
  NAND2_X1 u0_u5_u1_U9 (.ZN( u0_u5_u1_n114 ) , .A1( u0_u5_u1_n134 ) , .A2( u0_u5_u1_n156 ) );
  INV_X1 u0_u5_u1_U90 (.A( u0_u5_u1_n145 ) , .ZN( u0_u5_u1_n186 ) );
  NAND4_X1 u0_u5_u1_U91 (.ZN( u0_out5_2 ) , .A4( u0_u5_u1_n142 ) , .A3( u0_u5_u1_n143 ) , .A2( u0_u5_u1_n144 ) , .A1( u0_u5_u1_n179 ) );
  OAI21_X1 u0_u5_u1_U92 (.B2( u0_u5_u1_n132 ) , .ZN( u0_u5_u1_n144 ) , .A( u0_u5_u1_n146 ) , .B1( u0_u5_u1_n180 ) );
  INV_X1 u0_u5_u1_U93 (.A( u0_u5_u1_n130 ) , .ZN( u0_u5_u1_n179 ) );
  OR4_X1 u0_u5_u1_U94 (.ZN( u0_out5_13 ) , .A4( u0_u5_u1_n108 ) , .A3( u0_u5_u1_n109 ) , .A2( u0_u5_u1_n110 ) , .A1( u0_u5_u1_n111 ) );
  AOI21_X1 u0_u5_u1_U95 (.ZN( u0_u5_u1_n110 ) , .A( u0_u5_u1_n116 ) , .B1( u0_u5_u1_n152 ) , .B2( u0_u5_u1_n160 ) );
  AOI21_X1 u0_u5_u1_U96 (.ZN( u0_u5_u1_n111 ) , .A( u0_u5_u1_n128 ) , .B2( u0_u5_u1_n131 ) , .B1( u0_u5_u1_n135 ) );
  NAND3_X1 u0_u5_u1_U97 (.A3( u0_u5_u1_n149 ) , .A2( u0_u5_u1_n150 ) , .A1( u0_u5_u1_n151 ) , .ZN( u0_u5_u1_n164 ) );
  NAND3_X1 u0_u5_u1_U98 (.A3( u0_u5_u1_n134 ) , .A2( u0_u5_u1_n135 ) , .ZN( u0_u5_u1_n136 ) , .A1( u0_u5_u1_n151 ) );
  NAND3_X1 u0_u5_u1_U99 (.A1( u0_u5_u1_n133 ) , .ZN( u0_u5_u1_n137 ) , .A2( u0_u5_u1_n154 ) , .A3( u0_u5_u1_n181 ) );
  OAI22_X1 u0_u5_u2_U10 (.ZN( u0_u5_u2_n109 ) , .A2( u0_u5_u2_n113 ) , .B2( u0_u5_u2_n133 ) , .B1( u0_u5_u2_n167 ) , .A1( u0_u5_u2_n168 ) );
  NAND3_X1 u0_u5_u2_U100 (.A2( u0_u5_u2_n100 ) , .A1( u0_u5_u2_n104 ) , .A3( u0_u5_u2_n138 ) , .ZN( u0_u5_u2_n98 ) );
  OAI22_X1 u0_u5_u2_U11 (.B1( u0_u5_u2_n151 ) , .A2( u0_u5_u2_n152 ) , .A1( u0_u5_u2_n153 ) , .ZN( u0_u5_u2_n160 ) , .B2( u0_u5_u2_n168 ) );
  NOR3_X1 u0_u5_u2_U12 (.A1( u0_u5_u2_n150 ) , .ZN( u0_u5_u2_n151 ) , .A3( u0_u5_u2_n175 ) , .A2( u0_u5_u2_n188 ) );
  AOI21_X1 u0_u5_u2_U13 (.ZN( u0_u5_u2_n144 ) , .B2( u0_u5_u2_n155 ) , .A( u0_u5_u2_n172 ) , .B1( u0_u5_u2_n185 ) );
  AOI21_X1 u0_u5_u2_U14 (.B2( u0_u5_u2_n143 ) , .ZN( u0_u5_u2_n145 ) , .B1( u0_u5_u2_n152 ) , .A( u0_u5_u2_n171 ) );
  AOI21_X1 u0_u5_u2_U15 (.B2( u0_u5_u2_n120 ) , .B1( u0_u5_u2_n121 ) , .ZN( u0_u5_u2_n126 ) , .A( u0_u5_u2_n167 ) );
  INV_X1 u0_u5_u2_U16 (.A( u0_u5_u2_n156 ) , .ZN( u0_u5_u2_n171 ) );
  INV_X1 u0_u5_u2_U17 (.A( u0_u5_u2_n120 ) , .ZN( u0_u5_u2_n188 ) );
  NAND2_X1 u0_u5_u2_U18 (.A2( u0_u5_u2_n122 ) , .ZN( u0_u5_u2_n150 ) , .A1( u0_u5_u2_n152 ) );
  INV_X1 u0_u5_u2_U19 (.A( u0_u5_u2_n153 ) , .ZN( u0_u5_u2_n170 ) );
  INV_X1 u0_u5_u2_U20 (.A( u0_u5_u2_n137 ) , .ZN( u0_u5_u2_n173 ) );
  NAND2_X1 u0_u5_u2_U21 (.A1( u0_u5_u2_n132 ) , .A2( u0_u5_u2_n139 ) , .ZN( u0_u5_u2_n157 ) );
  INV_X1 u0_u5_u2_U22 (.A( u0_u5_u2_n113 ) , .ZN( u0_u5_u2_n178 ) );
  INV_X1 u0_u5_u2_U23 (.A( u0_u5_u2_n139 ) , .ZN( u0_u5_u2_n175 ) );
  INV_X1 u0_u5_u2_U24 (.A( u0_u5_u2_n155 ) , .ZN( u0_u5_u2_n181 ) );
  INV_X1 u0_u5_u2_U25 (.A( u0_u5_u2_n119 ) , .ZN( u0_u5_u2_n177 ) );
  INV_X1 u0_u5_u2_U26 (.A( u0_u5_u2_n116 ) , .ZN( u0_u5_u2_n180 ) );
  INV_X1 u0_u5_u2_U27 (.A( u0_u5_u2_n131 ) , .ZN( u0_u5_u2_n179 ) );
  INV_X1 u0_u5_u2_U28 (.A( u0_u5_u2_n154 ) , .ZN( u0_u5_u2_n176 ) );
  NAND2_X1 u0_u5_u2_U29 (.A2( u0_u5_u2_n116 ) , .A1( u0_u5_u2_n117 ) , .ZN( u0_u5_u2_n118 ) );
  NOR2_X1 u0_u5_u2_U3 (.ZN( u0_u5_u2_n121 ) , .A2( u0_u5_u2_n177 ) , .A1( u0_u5_u2_n180 ) );
  INV_X1 u0_u5_u2_U30 (.A( u0_u5_u2_n132 ) , .ZN( u0_u5_u2_n182 ) );
  INV_X1 u0_u5_u2_U31 (.A( u0_u5_u2_n158 ) , .ZN( u0_u5_u2_n183 ) );
  OAI21_X1 u0_u5_u2_U32 (.A( u0_u5_u2_n156 ) , .B1( u0_u5_u2_n157 ) , .ZN( u0_u5_u2_n158 ) , .B2( u0_u5_u2_n179 ) );
  NOR2_X1 u0_u5_u2_U33 (.ZN( u0_u5_u2_n156 ) , .A1( u0_u5_u2_n166 ) , .A2( u0_u5_u2_n169 ) );
  NOR2_X1 u0_u5_u2_U34 (.A2( u0_u5_u2_n114 ) , .ZN( u0_u5_u2_n137 ) , .A1( u0_u5_u2_n140 ) );
  NOR2_X1 u0_u5_u2_U35 (.A2( u0_u5_u2_n138 ) , .ZN( u0_u5_u2_n153 ) , .A1( u0_u5_u2_n156 ) );
  AOI211_X1 u0_u5_u2_U36 (.ZN( u0_u5_u2_n130 ) , .C1( u0_u5_u2_n138 ) , .C2( u0_u5_u2_n179 ) , .B( u0_u5_u2_n96 ) , .A( u0_u5_u2_n97 ) );
  OAI22_X1 u0_u5_u2_U37 (.B1( u0_u5_u2_n133 ) , .A2( u0_u5_u2_n137 ) , .A1( u0_u5_u2_n152 ) , .B2( u0_u5_u2_n168 ) , .ZN( u0_u5_u2_n97 ) );
  OAI221_X1 u0_u5_u2_U38 (.B1( u0_u5_u2_n113 ) , .C1( u0_u5_u2_n132 ) , .A( u0_u5_u2_n149 ) , .B2( u0_u5_u2_n171 ) , .C2( u0_u5_u2_n172 ) , .ZN( u0_u5_u2_n96 ) );
  OAI221_X1 u0_u5_u2_U39 (.A( u0_u5_u2_n115 ) , .C2( u0_u5_u2_n123 ) , .B2( u0_u5_u2_n143 ) , .B1( u0_u5_u2_n153 ) , .ZN( u0_u5_u2_n163 ) , .C1( u0_u5_u2_n168 ) );
  INV_X1 u0_u5_u2_U4 (.A( u0_u5_u2_n134 ) , .ZN( u0_u5_u2_n185 ) );
  OAI21_X1 u0_u5_u2_U40 (.A( u0_u5_u2_n114 ) , .ZN( u0_u5_u2_n115 ) , .B1( u0_u5_u2_n176 ) , .B2( u0_u5_u2_n178 ) );
  OAI221_X1 u0_u5_u2_U41 (.A( u0_u5_u2_n135 ) , .B2( u0_u5_u2_n136 ) , .B1( u0_u5_u2_n137 ) , .ZN( u0_u5_u2_n162 ) , .C2( u0_u5_u2_n167 ) , .C1( u0_u5_u2_n185 ) );
  AND3_X1 u0_u5_u2_U42 (.A3( u0_u5_u2_n131 ) , .A2( u0_u5_u2_n132 ) , .A1( u0_u5_u2_n133 ) , .ZN( u0_u5_u2_n136 ) );
  AOI22_X1 u0_u5_u2_U43 (.ZN( u0_u5_u2_n135 ) , .B1( u0_u5_u2_n140 ) , .A1( u0_u5_u2_n156 ) , .B2( u0_u5_u2_n180 ) , .A2( u0_u5_u2_n188 ) );
  AOI21_X1 u0_u5_u2_U44 (.ZN( u0_u5_u2_n149 ) , .B1( u0_u5_u2_n173 ) , .B2( u0_u5_u2_n188 ) , .A( u0_u5_u2_n95 ) );
  AND3_X1 u0_u5_u2_U45 (.A2( u0_u5_u2_n100 ) , .A1( u0_u5_u2_n104 ) , .A3( u0_u5_u2_n156 ) , .ZN( u0_u5_u2_n95 ) );
  OAI21_X1 u0_u5_u2_U46 (.A( u0_u5_u2_n141 ) , .B2( u0_u5_u2_n142 ) , .ZN( u0_u5_u2_n146 ) , .B1( u0_u5_u2_n153 ) );
  OAI21_X1 u0_u5_u2_U47 (.A( u0_u5_u2_n140 ) , .ZN( u0_u5_u2_n141 ) , .B1( u0_u5_u2_n176 ) , .B2( u0_u5_u2_n177 ) );
  NOR3_X1 u0_u5_u2_U48 (.ZN( u0_u5_u2_n142 ) , .A3( u0_u5_u2_n175 ) , .A2( u0_u5_u2_n178 ) , .A1( u0_u5_u2_n181 ) );
  OAI21_X1 u0_u5_u2_U49 (.A( u0_u5_u2_n101 ) , .B2( u0_u5_u2_n121 ) , .B1( u0_u5_u2_n153 ) , .ZN( u0_u5_u2_n164 ) );
  INV_X1 u0_u5_u2_U5 (.A( u0_u5_u2_n150 ) , .ZN( u0_u5_u2_n184 ) );
  NAND2_X1 u0_u5_u2_U50 (.A2( u0_u5_u2_n100 ) , .A1( u0_u5_u2_n107 ) , .ZN( u0_u5_u2_n155 ) );
  NAND2_X1 u0_u5_u2_U51 (.A2( u0_u5_u2_n105 ) , .A1( u0_u5_u2_n108 ) , .ZN( u0_u5_u2_n143 ) );
  NAND2_X1 u0_u5_u2_U52 (.A1( u0_u5_u2_n104 ) , .A2( u0_u5_u2_n106 ) , .ZN( u0_u5_u2_n152 ) );
  NAND2_X1 u0_u5_u2_U53 (.A1( u0_u5_u2_n100 ) , .A2( u0_u5_u2_n105 ) , .ZN( u0_u5_u2_n132 ) );
  INV_X1 u0_u5_u2_U54 (.A( u0_u5_u2_n140 ) , .ZN( u0_u5_u2_n168 ) );
  INV_X1 u0_u5_u2_U55 (.A( u0_u5_u2_n138 ) , .ZN( u0_u5_u2_n167 ) );
  NAND2_X1 u0_u5_u2_U56 (.A1( u0_u5_u2_n102 ) , .A2( u0_u5_u2_n106 ) , .ZN( u0_u5_u2_n113 ) );
  NAND2_X1 u0_u5_u2_U57 (.A1( u0_u5_u2_n106 ) , .A2( u0_u5_u2_n107 ) , .ZN( u0_u5_u2_n131 ) );
  NAND2_X1 u0_u5_u2_U58 (.A1( u0_u5_u2_n103 ) , .A2( u0_u5_u2_n107 ) , .ZN( u0_u5_u2_n139 ) );
  NAND2_X1 u0_u5_u2_U59 (.A1( u0_u5_u2_n103 ) , .A2( u0_u5_u2_n105 ) , .ZN( u0_u5_u2_n133 ) );
  NOR4_X1 u0_u5_u2_U6 (.A4( u0_u5_u2_n124 ) , .A3( u0_u5_u2_n125 ) , .A2( u0_u5_u2_n126 ) , .A1( u0_u5_u2_n127 ) , .ZN( u0_u5_u2_n128 ) );
  NAND2_X1 u0_u5_u2_U60 (.A1( u0_u5_u2_n102 ) , .A2( u0_u5_u2_n103 ) , .ZN( u0_u5_u2_n154 ) );
  NAND2_X1 u0_u5_u2_U61 (.A2( u0_u5_u2_n103 ) , .A1( u0_u5_u2_n104 ) , .ZN( u0_u5_u2_n119 ) );
  NAND2_X1 u0_u5_u2_U62 (.A2( u0_u5_u2_n107 ) , .A1( u0_u5_u2_n108 ) , .ZN( u0_u5_u2_n123 ) );
  NAND2_X1 u0_u5_u2_U63 (.A1( u0_u5_u2_n104 ) , .A2( u0_u5_u2_n108 ) , .ZN( u0_u5_u2_n122 ) );
  INV_X1 u0_u5_u2_U64 (.A( u0_u5_u2_n114 ) , .ZN( u0_u5_u2_n172 ) );
  NAND2_X1 u0_u5_u2_U65 (.A2( u0_u5_u2_n100 ) , .A1( u0_u5_u2_n102 ) , .ZN( u0_u5_u2_n116 ) );
  NAND2_X1 u0_u5_u2_U66 (.A1( u0_u5_u2_n102 ) , .A2( u0_u5_u2_n108 ) , .ZN( u0_u5_u2_n120 ) );
  NAND2_X1 u0_u5_u2_U67 (.A2( u0_u5_u2_n105 ) , .A1( u0_u5_u2_n106 ) , .ZN( u0_u5_u2_n117 ) );
  INV_X1 u0_u5_u2_U68 (.ZN( u0_u5_u2_n187 ) , .A( u0_u5_u2_n99 ) );
  OAI21_X1 u0_u5_u2_U69 (.B1( u0_u5_u2_n137 ) , .B2( u0_u5_u2_n143 ) , .A( u0_u5_u2_n98 ) , .ZN( u0_u5_u2_n99 ) );
  AOI21_X1 u0_u5_u2_U7 (.B2( u0_u5_u2_n119 ) , .ZN( u0_u5_u2_n127 ) , .A( u0_u5_u2_n137 ) , .B1( u0_u5_u2_n155 ) );
  NOR2_X1 u0_u5_u2_U70 (.A2( u0_u5_X_16 ) , .ZN( u0_u5_u2_n140 ) , .A1( u0_u5_u2_n166 ) );
  NOR2_X1 u0_u5_u2_U71 (.A2( u0_u5_X_13 ) , .A1( u0_u5_X_14 ) , .ZN( u0_u5_u2_n100 ) );
  NOR2_X1 u0_u5_u2_U72 (.A2( u0_u5_X_16 ) , .A1( u0_u5_X_17 ) , .ZN( u0_u5_u2_n138 ) );
  NOR2_X1 u0_u5_u2_U73 (.A2( u0_u5_X_15 ) , .A1( u0_u5_X_18 ) , .ZN( u0_u5_u2_n104 ) );
  NOR2_X1 u0_u5_u2_U74 (.A2( u0_u5_X_14 ) , .ZN( u0_u5_u2_n103 ) , .A1( u0_u5_u2_n174 ) );
  NOR2_X1 u0_u5_u2_U75 (.A2( u0_u5_X_15 ) , .ZN( u0_u5_u2_n102 ) , .A1( u0_u5_u2_n165 ) );
  NOR2_X1 u0_u5_u2_U76 (.A2( u0_u5_X_17 ) , .ZN( u0_u5_u2_n114 ) , .A1( u0_u5_u2_n169 ) );
  AND2_X1 u0_u5_u2_U77 (.A1( u0_u5_X_15 ) , .ZN( u0_u5_u2_n105 ) , .A2( u0_u5_u2_n165 ) );
  AND2_X1 u0_u5_u2_U78 (.A2( u0_u5_X_15 ) , .A1( u0_u5_X_18 ) , .ZN( u0_u5_u2_n107 ) );
  AND2_X1 u0_u5_u2_U79 (.A1( u0_u5_X_14 ) , .ZN( u0_u5_u2_n106 ) , .A2( u0_u5_u2_n174 ) );
  AOI21_X1 u0_u5_u2_U8 (.ZN( u0_u5_u2_n124 ) , .B1( u0_u5_u2_n131 ) , .B2( u0_u5_u2_n143 ) , .A( u0_u5_u2_n172 ) );
  AND2_X1 u0_u5_u2_U80 (.A1( u0_u5_X_13 ) , .A2( u0_u5_X_14 ) , .ZN( u0_u5_u2_n108 ) );
  INV_X1 u0_u5_u2_U81 (.A( u0_u5_X_16 ) , .ZN( u0_u5_u2_n169 ) );
  INV_X1 u0_u5_u2_U82 (.A( u0_u5_X_17 ) , .ZN( u0_u5_u2_n166 ) );
  INV_X1 u0_u5_u2_U83 (.A( u0_u5_X_13 ) , .ZN( u0_u5_u2_n174 ) );
  INV_X1 u0_u5_u2_U84 (.A( u0_u5_X_18 ) , .ZN( u0_u5_u2_n165 ) );
  NAND4_X1 u0_u5_u2_U85 (.ZN( u0_out5_30 ) , .A4( u0_u5_u2_n147 ) , .A3( u0_u5_u2_n148 ) , .A2( u0_u5_u2_n149 ) , .A1( u0_u5_u2_n187 ) );
  NOR3_X1 u0_u5_u2_U86 (.A3( u0_u5_u2_n144 ) , .A2( u0_u5_u2_n145 ) , .A1( u0_u5_u2_n146 ) , .ZN( u0_u5_u2_n147 ) );
  AOI21_X1 u0_u5_u2_U87 (.B2( u0_u5_u2_n138 ) , .ZN( u0_u5_u2_n148 ) , .A( u0_u5_u2_n162 ) , .B1( u0_u5_u2_n182 ) );
  NAND4_X1 u0_u5_u2_U88 (.ZN( u0_out5_24 ) , .A4( u0_u5_u2_n111 ) , .A3( u0_u5_u2_n112 ) , .A1( u0_u5_u2_n130 ) , .A2( u0_u5_u2_n187 ) );
  AOI221_X1 u0_u5_u2_U89 (.A( u0_u5_u2_n109 ) , .B1( u0_u5_u2_n110 ) , .ZN( u0_u5_u2_n111 ) , .C1( u0_u5_u2_n134 ) , .C2( u0_u5_u2_n170 ) , .B2( u0_u5_u2_n173 ) );
  AOI21_X1 u0_u5_u2_U9 (.B2( u0_u5_u2_n123 ) , .ZN( u0_u5_u2_n125 ) , .A( u0_u5_u2_n171 ) , .B1( u0_u5_u2_n184 ) );
  AOI21_X1 u0_u5_u2_U90 (.ZN( u0_u5_u2_n112 ) , .B2( u0_u5_u2_n156 ) , .A( u0_u5_u2_n164 ) , .B1( u0_u5_u2_n181 ) );
  NAND4_X1 u0_u5_u2_U91 (.ZN( u0_out5_16 ) , .A4( u0_u5_u2_n128 ) , .A3( u0_u5_u2_n129 ) , .A1( u0_u5_u2_n130 ) , .A2( u0_u5_u2_n186 ) );
  AOI22_X1 u0_u5_u2_U92 (.A2( u0_u5_u2_n118 ) , .ZN( u0_u5_u2_n129 ) , .A1( u0_u5_u2_n140 ) , .B1( u0_u5_u2_n157 ) , .B2( u0_u5_u2_n170 ) );
  INV_X1 u0_u5_u2_U93 (.A( u0_u5_u2_n163 ) , .ZN( u0_u5_u2_n186 ) );
  OR4_X1 u0_u5_u2_U94 (.ZN( u0_out5_6 ) , .A4( u0_u5_u2_n161 ) , .A3( u0_u5_u2_n162 ) , .A2( u0_u5_u2_n163 ) , .A1( u0_u5_u2_n164 ) );
  OR3_X1 u0_u5_u2_U95 (.A2( u0_u5_u2_n159 ) , .A1( u0_u5_u2_n160 ) , .ZN( u0_u5_u2_n161 ) , .A3( u0_u5_u2_n183 ) );
  AOI21_X1 u0_u5_u2_U96 (.B2( u0_u5_u2_n154 ) , .B1( u0_u5_u2_n155 ) , .ZN( u0_u5_u2_n159 ) , .A( u0_u5_u2_n167 ) );
  NAND3_X1 u0_u5_u2_U97 (.A2( u0_u5_u2_n117 ) , .A1( u0_u5_u2_n122 ) , .A3( u0_u5_u2_n123 ) , .ZN( u0_u5_u2_n134 ) );
  NAND3_X1 u0_u5_u2_U98 (.ZN( u0_u5_u2_n110 ) , .A2( u0_u5_u2_n131 ) , .A3( u0_u5_u2_n139 ) , .A1( u0_u5_u2_n154 ) );
  NAND3_X1 u0_u5_u2_U99 (.A2( u0_u5_u2_n100 ) , .ZN( u0_u5_u2_n101 ) , .A1( u0_u5_u2_n104 ) , .A3( u0_u5_u2_n114 ) );
  OAI22_X1 u0_u5_u3_U10 (.B1( u0_u5_u3_n113 ) , .A2( u0_u5_u3_n135 ) , .A1( u0_u5_u3_n150 ) , .B2( u0_u5_u3_n164 ) , .ZN( u0_u5_u3_n98 ) );
  OAI211_X1 u0_u5_u3_U11 (.B( u0_u5_u3_n106 ) , .ZN( u0_u5_u3_n119 ) , .C2( u0_u5_u3_n128 ) , .C1( u0_u5_u3_n167 ) , .A( u0_u5_u3_n181 ) );
  AOI221_X1 u0_u5_u3_U12 (.C1( u0_u5_u3_n105 ) , .ZN( u0_u5_u3_n106 ) , .A( u0_u5_u3_n131 ) , .B2( u0_u5_u3_n132 ) , .C2( u0_u5_u3_n133 ) , .B1( u0_u5_u3_n169 ) );
  INV_X1 u0_u5_u3_U13 (.ZN( u0_u5_u3_n181 ) , .A( u0_u5_u3_n98 ) );
  NAND2_X1 u0_u5_u3_U14 (.ZN( u0_u5_u3_n105 ) , .A2( u0_u5_u3_n130 ) , .A1( u0_u5_u3_n155 ) );
  AOI22_X1 u0_u5_u3_U15 (.B1( u0_u5_u3_n115 ) , .A2( u0_u5_u3_n116 ) , .ZN( u0_u5_u3_n123 ) , .B2( u0_u5_u3_n133 ) , .A1( u0_u5_u3_n169 ) );
  NAND2_X1 u0_u5_u3_U16 (.ZN( u0_u5_u3_n116 ) , .A2( u0_u5_u3_n151 ) , .A1( u0_u5_u3_n182 ) );
  NOR2_X1 u0_u5_u3_U17 (.ZN( u0_u5_u3_n126 ) , .A2( u0_u5_u3_n150 ) , .A1( u0_u5_u3_n164 ) );
  AOI21_X1 u0_u5_u3_U18 (.ZN( u0_u5_u3_n112 ) , .B2( u0_u5_u3_n146 ) , .B1( u0_u5_u3_n155 ) , .A( u0_u5_u3_n167 ) );
  NAND2_X1 u0_u5_u3_U19 (.A1( u0_u5_u3_n135 ) , .ZN( u0_u5_u3_n142 ) , .A2( u0_u5_u3_n164 ) );
  NAND2_X1 u0_u5_u3_U20 (.ZN( u0_u5_u3_n132 ) , .A2( u0_u5_u3_n152 ) , .A1( u0_u5_u3_n156 ) );
  AND2_X1 u0_u5_u3_U21 (.A2( u0_u5_u3_n113 ) , .A1( u0_u5_u3_n114 ) , .ZN( u0_u5_u3_n151 ) );
  INV_X1 u0_u5_u3_U22 (.A( u0_u5_u3_n133 ) , .ZN( u0_u5_u3_n165 ) );
  INV_X1 u0_u5_u3_U23 (.A( u0_u5_u3_n135 ) , .ZN( u0_u5_u3_n170 ) );
  NAND2_X1 u0_u5_u3_U24 (.A1( u0_u5_u3_n107 ) , .A2( u0_u5_u3_n108 ) , .ZN( u0_u5_u3_n140 ) );
  NAND2_X1 u0_u5_u3_U25 (.ZN( u0_u5_u3_n117 ) , .A1( u0_u5_u3_n124 ) , .A2( u0_u5_u3_n148 ) );
  NAND2_X1 u0_u5_u3_U26 (.ZN( u0_u5_u3_n143 ) , .A1( u0_u5_u3_n165 ) , .A2( u0_u5_u3_n167 ) );
  INV_X1 u0_u5_u3_U27 (.A( u0_u5_u3_n130 ) , .ZN( u0_u5_u3_n177 ) );
  INV_X1 u0_u5_u3_U28 (.A( u0_u5_u3_n128 ) , .ZN( u0_u5_u3_n176 ) );
  INV_X1 u0_u5_u3_U29 (.A( u0_u5_u3_n155 ) , .ZN( u0_u5_u3_n174 ) );
  INV_X1 u0_u5_u3_U3 (.A( u0_u5_u3_n129 ) , .ZN( u0_u5_u3_n183 ) );
  INV_X1 u0_u5_u3_U30 (.A( u0_u5_u3_n139 ) , .ZN( u0_u5_u3_n185 ) );
  NOR2_X1 u0_u5_u3_U31 (.ZN( u0_u5_u3_n135 ) , .A2( u0_u5_u3_n141 ) , .A1( u0_u5_u3_n169 ) );
  OAI222_X1 u0_u5_u3_U32 (.C2( u0_u5_u3_n107 ) , .A2( u0_u5_u3_n108 ) , .B1( u0_u5_u3_n135 ) , .ZN( u0_u5_u3_n138 ) , .B2( u0_u5_u3_n146 ) , .C1( u0_u5_u3_n154 ) , .A1( u0_u5_u3_n164 ) );
  NOR4_X1 u0_u5_u3_U33 (.A4( u0_u5_u3_n157 ) , .A3( u0_u5_u3_n158 ) , .A2( u0_u5_u3_n159 ) , .A1( u0_u5_u3_n160 ) , .ZN( u0_u5_u3_n161 ) );
  AOI21_X1 u0_u5_u3_U34 (.B2( u0_u5_u3_n152 ) , .B1( u0_u5_u3_n153 ) , .ZN( u0_u5_u3_n158 ) , .A( u0_u5_u3_n164 ) );
  AOI21_X1 u0_u5_u3_U35 (.A( u0_u5_u3_n154 ) , .B2( u0_u5_u3_n155 ) , .B1( u0_u5_u3_n156 ) , .ZN( u0_u5_u3_n157 ) );
  AOI21_X1 u0_u5_u3_U36 (.A( u0_u5_u3_n149 ) , .B2( u0_u5_u3_n150 ) , .B1( u0_u5_u3_n151 ) , .ZN( u0_u5_u3_n159 ) );
  AOI211_X1 u0_u5_u3_U37 (.ZN( u0_u5_u3_n109 ) , .A( u0_u5_u3_n119 ) , .C2( u0_u5_u3_n129 ) , .B( u0_u5_u3_n138 ) , .C1( u0_u5_u3_n141 ) );
  AOI211_X1 u0_u5_u3_U38 (.B( u0_u5_u3_n119 ) , .A( u0_u5_u3_n120 ) , .C2( u0_u5_u3_n121 ) , .ZN( u0_u5_u3_n122 ) , .C1( u0_u5_u3_n179 ) );
  INV_X1 u0_u5_u3_U39 (.A( u0_u5_u3_n156 ) , .ZN( u0_u5_u3_n179 ) );
  INV_X1 u0_u5_u3_U4 (.A( u0_u5_u3_n140 ) , .ZN( u0_u5_u3_n182 ) );
  OAI22_X1 u0_u5_u3_U40 (.B1( u0_u5_u3_n118 ) , .ZN( u0_u5_u3_n120 ) , .A1( u0_u5_u3_n135 ) , .B2( u0_u5_u3_n154 ) , .A2( u0_u5_u3_n178 ) );
  AND3_X1 u0_u5_u3_U41 (.ZN( u0_u5_u3_n118 ) , .A2( u0_u5_u3_n124 ) , .A1( u0_u5_u3_n144 ) , .A3( u0_u5_u3_n152 ) );
  INV_X1 u0_u5_u3_U42 (.A( u0_u5_u3_n121 ) , .ZN( u0_u5_u3_n164 ) );
  NAND2_X1 u0_u5_u3_U43 (.ZN( u0_u5_u3_n133 ) , .A1( u0_u5_u3_n154 ) , .A2( u0_u5_u3_n164 ) );
  OAI211_X1 u0_u5_u3_U44 (.B( u0_u5_u3_n127 ) , .ZN( u0_u5_u3_n139 ) , .C1( u0_u5_u3_n150 ) , .C2( u0_u5_u3_n154 ) , .A( u0_u5_u3_n184 ) );
  INV_X1 u0_u5_u3_U45 (.A( u0_u5_u3_n125 ) , .ZN( u0_u5_u3_n184 ) );
  AOI221_X1 u0_u5_u3_U46 (.A( u0_u5_u3_n126 ) , .ZN( u0_u5_u3_n127 ) , .C2( u0_u5_u3_n132 ) , .C1( u0_u5_u3_n169 ) , .B2( u0_u5_u3_n170 ) , .B1( u0_u5_u3_n174 ) );
  OAI22_X1 u0_u5_u3_U47 (.A1( u0_u5_u3_n124 ) , .ZN( u0_u5_u3_n125 ) , .B2( u0_u5_u3_n145 ) , .A2( u0_u5_u3_n165 ) , .B1( u0_u5_u3_n167 ) );
  NOR2_X1 u0_u5_u3_U48 (.A1( u0_u5_u3_n113 ) , .ZN( u0_u5_u3_n131 ) , .A2( u0_u5_u3_n154 ) );
  NAND2_X1 u0_u5_u3_U49 (.A1( u0_u5_u3_n103 ) , .ZN( u0_u5_u3_n150 ) , .A2( u0_u5_u3_n99 ) );
  INV_X1 u0_u5_u3_U5 (.A( u0_u5_u3_n117 ) , .ZN( u0_u5_u3_n178 ) );
  NAND2_X1 u0_u5_u3_U50 (.A2( u0_u5_u3_n102 ) , .ZN( u0_u5_u3_n155 ) , .A1( u0_u5_u3_n97 ) );
  INV_X1 u0_u5_u3_U51 (.A( u0_u5_u3_n141 ) , .ZN( u0_u5_u3_n167 ) );
  AOI21_X1 u0_u5_u3_U52 (.B2( u0_u5_u3_n114 ) , .B1( u0_u5_u3_n146 ) , .A( u0_u5_u3_n154 ) , .ZN( u0_u5_u3_n94 ) );
  AOI21_X1 u0_u5_u3_U53 (.ZN( u0_u5_u3_n110 ) , .B2( u0_u5_u3_n142 ) , .B1( u0_u5_u3_n186 ) , .A( u0_u5_u3_n95 ) );
  INV_X1 u0_u5_u3_U54 (.A( u0_u5_u3_n145 ) , .ZN( u0_u5_u3_n186 ) );
  AOI21_X1 u0_u5_u3_U55 (.B1( u0_u5_u3_n124 ) , .A( u0_u5_u3_n149 ) , .B2( u0_u5_u3_n155 ) , .ZN( u0_u5_u3_n95 ) );
  INV_X1 u0_u5_u3_U56 (.A( u0_u5_u3_n149 ) , .ZN( u0_u5_u3_n169 ) );
  NAND2_X1 u0_u5_u3_U57 (.ZN( u0_u5_u3_n124 ) , .A1( u0_u5_u3_n96 ) , .A2( u0_u5_u3_n97 ) );
  NAND2_X1 u0_u5_u3_U58 (.A2( u0_u5_u3_n100 ) , .ZN( u0_u5_u3_n146 ) , .A1( u0_u5_u3_n96 ) );
  NAND2_X1 u0_u5_u3_U59 (.A1( u0_u5_u3_n101 ) , .ZN( u0_u5_u3_n145 ) , .A2( u0_u5_u3_n99 ) );
  AOI221_X1 u0_u5_u3_U6 (.A( u0_u5_u3_n131 ) , .C2( u0_u5_u3_n132 ) , .C1( u0_u5_u3_n133 ) , .ZN( u0_u5_u3_n134 ) , .B1( u0_u5_u3_n143 ) , .B2( u0_u5_u3_n177 ) );
  NAND2_X1 u0_u5_u3_U60 (.A1( u0_u5_u3_n100 ) , .ZN( u0_u5_u3_n156 ) , .A2( u0_u5_u3_n99 ) );
  NAND2_X1 u0_u5_u3_U61 (.A2( u0_u5_u3_n101 ) , .A1( u0_u5_u3_n104 ) , .ZN( u0_u5_u3_n148 ) );
  NAND2_X1 u0_u5_u3_U62 (.A1( u0_u5_u3_n100 ) , .A2( u0_u5_u3_n102 ) , .ZN( u0_u5_u3_n128 ) );
  NAND2_X1 u0_u5_u3_U63 (.A2( u0_u5_u3_n101 ) , .A1( u0_u5_u3_n102 ) , .ZN( u0_u5_u3_n152 ) );
  NAND2_X1 u0_u5_u3_U64 (.A2( u0_u5_u3_n101 ) , .ZN( u0_u5_u3_n114 ) , .A1( u0_u5_u3_n96 ) );
  NAND2_X1 u0_u5_u3_U65 (.ZN( u0_u5_u3_n107 ) , .A1( u0_u5_u3_n97 ) , .A2( u0_u5_u3_n99 ) );
  NAND2_X1 u0_u5_u3_U66 (.A2( u0_u5_u3_n100 ) , .A1( u0_u5_u3_n104 ) , .ZN( u0_u5_u3_n113 ) );
  NAND2_X1 u0_u5_u3_U67 (.A1( u0_u5_u3_n104 ) , .ZN( u0_u5_u3_n153 ) , .A2( u0_u5_u3_n97 ) );
  NAND2_X1 u0_u5_u3_U68 (.A2( u0_u5_u3_n103 ) , .A1( u0_u5_u3_n104 ) , .ZN( u0_u5_u3_n130 ) );
  NAND2_X1 u0_u5_u3_U69 (.A2( u0_u5_u3_n103 ) , .ZN( u0_u5_u3_n144 ) , .A1( u0_u5_u3_n96 ) );
  OAI22_X1 u0_u5_u3_U7 (.B2( u0_u5_u3_n147 ) , .A2( u0_u5_u3_n148 ) , .ZN( u0_u5_u3_n160 ) , .B1( u0_u5_u3_n165 ) , .A1( u0_u5_u3_n168 ) );
  NAND2_X1 u0_u5_u3_U70 (.A1( u0_u5_u3_n102 ) , .A2( u0_u5_u3_n103 ) , .ZN( u0_u5_u3_n108 ) );
  NOR2_X1 u0_u5_u3_U71 (.A2( u0_u5_X_19 ) , .A1( u0_u5_X_20 ) , .ZN( u0_u5_u3_n99 ) );
  NOR2_X1 u0_u5_u3_U72 (.A2( u0_u5_X_21 ) , .A1( u0_u5_X_24 ) , .ZN( u0_u5_u3_n103 ) );
  NOR2_X1 u0_u5_u3_U73 (.A2( u0_u5_X_24 ) , .A1( u0_u5_u3_n171 ) , .ZN( u0_u5_u3_n97 ) );
  NOR2_X1 u0_u5_u3_U74 (.A2( u0_u5_X_23 ) , .ZN( u0_u5_u3_n141 ) , .A1( u0_u5_u3_n166 ) );
  NOR2_X1 u0_u5_u3_U75 (.A2( u0_u5_X_19 ) , .A1( u0_u5_u3_n172 ) , .ZN( u0_u5_u3_n96 ) );
  NAND2_X1 u0_u5_u3_U76 (.A1( u0_u5_X_22 ) , .A2( u0_u5_X_23 ) , .ZN( u0_u5_u3_n154 ) );
  NAND2_X1 u0_u5_u3_U77 (.A1( u0_u5_X_23 ) , .ZN( u0_u5_u3_n149 ) , .A2( u0_u5_u3_n166 ) );
  NOR2_X1 u0_u5_u3_U78 (.A2( u0_u5_X_22 ) , .A1( u0_u5_X_23 ) , .ZN( u0_u5_u3_n121 ) );
  AND2_X1 u0_u5_u3_U79 (.A1( u0_u5_X_24 ) , .ZN( u0_u5_u3_n101 ) , .A2( u0_u5_u3_n171 ) );
  AND3_X1 u0_u5_u3_U8 (.A3( u0_u5_u3_n144 ) , .A2( u0_u5_u3_n145 ) , .A1( u0_u5_u3_n146 ) , .ZN( u0_u5_u3_n147 ) );
  AND2_X1 u0_u5_u3_U80 (.A1( u0_u5_X_19 ) , .ZN( u0_u5_u3_n102 ) , .A2( u0_u5_u3_n172 ) );
  AND2_X1 u0_u5_u3_U81 (.A1( u0_u5_X_21 ) , .A2( u0_u5_X_24 ) , .ZN( u0_u5_u3_n100 ) );
  AND2_X1 u0_u5_u3_U82 (.A2( u0_u5_X_19 ) , .A1( u0_u5_X_20 ) , .ZN( u0_u5_u3_n104 ) );
  INV_X1 u0_u5_u3_U83 (.A( u0_u5_X_22 ) , .ZN( u0_u5_u3_n166 ) );
  INV_X1 u0_u5_u3_U84 (.A( u0_u5_X_21 ) , .ZN( u0_u5_u3_n171 ) );
  INV_X1 u0_u5_u3_U85 (.A( u0_u5_X_20 ) , .ZN( u0_u5_u3_n172 ) );
  NAND4_X1 u0_u5_u3_U86 (.ZN( u0_out5_26 ) , .A4( u0_u5_u3_n109 ) , .A3( u0_u5_u3_n110 ) , .A2( u0_u5_u3_n111 ) , .A1( u0_u5_u3_n173 ) );
  INV_X1 u0_u5_u3_U87 (.ZN( u0_u5_u3_n173 ) , .A( u0_u5_u3_n94 ) );
  OAI21_X1 u0_u5_u3_U88 (.ZN( u0_u5_u3_n111 ) , .B2( u0_u5_u3_n117 ) , .A( u0_u5_u3_n133 ) , .B1( u0_u5_u3_n176 ) );
  NAND4_X1 u0_u5_u3_U89 (.ZN( u0_out5_20 ) , .A4( u0_u5_u3_n122 ) , .A3( u0_u5_u3_n123 ) , .A1( u0_u5_u3_n175 ) , .A2( u0_u5_u3_n180 ) );
  INV_X1 u0_u5_u3_U9 (.A( u0_u5_u3_n143 ) , .ZN( u0_u5_u3_n168 ) );
  INV_X1 u0_u5_u3_U90 (.A( u0_u5_u3_n126 ) , .ZN( u0_u5_u3_n180 ) );
  INV_X1 u0_u5_u3_U91 (.A( u0_u5_u3_n112 ) , .ZN( u0_u5_u3_n175 ) );
  NAND4_X1 u0_u5_u3_U92 (.ZN( u0_out5_1 ) , .A4( u0_u5_u3_n161 ) , .A3( u0_u5_u3_n162 ) , .A2( u0_u5_u3_n163 ) , .A1( u0_u5_u3_n185 ) );
  NAND2_X1 u0_u5_u3_U93 (.ZN( u0_u5_u3_n163 ) , .A2( u0_u5_u3_n170 ) , .A1( u0_u5_u3_n176 ) );
  AOI22_X1 u0_u5_u3_U94 (.B2( u0_u5_u3_n140 ) , .B1( u0_u5_u3_n141 ) , .A2( u0_u5_u3_n142 ) , .ZN( u0_u5_u3_n162 ) , .A1( u0_u5_u3_n177 ) );
  OR4_X1 u0_u5_u3_U95 (.ZN( u0_out5_10 ) , .A4( u0_u5_u3_n136 ) , .A3( u0_u5_u3_n137 ) , .A1( u0_u5_u3_n138 ) , .A2( u0_u5_u3_n139 ) );
  OAI222_X1 u0_u5_u3_U96 (.C1( u0_u5_u3_n128 ) , .ZN( u0_u5_u3_n137 ) , .B1( u0_u5_u3_n148 ) , .A2( u0_u5_u3_n150 ) , .B2( u0_u5_u3_n154 ) , .C2( u0_u5_u3_n164 ) , .A1( u0_u5_u3_n167 ) );
  OAI221_X1 u0_u5_u3_U97 (.A( u0_u5_u3_n134 ) , .B2( u0_u5_u3_n135 ) , .ZN( u0_u5_u3_n136 ) , .C1( u0_u5_u3_n149 ) , .B1( u0_u5_u3_n151 ) , .C2( u0_u5_u3_n183 ) );
  NAND3_X1 u0_u5_u3_U98 (.A1( u0_u5_u3_n114 ) , .ZN( u0_u5_u3_n115 ) , .A2( u0_u5_u3_n145 ) , .A3( u0_u5_u3_n153 ) );
  NAND3_X1 u0_u5_u3_U99 (.ZN( u0_u5_u3_n129 ) , .A2( u0_u5_u3_n144 ) , .A1( u0_u5_u3_n153 ) , .A3( u0_u5_u3_n182 ) );
  INV_X1 u0_u5_u5_U10 (.A( u0_u5_u5_n121 ) , .ZN( u0_u5_u5_n177 ) );
  NOR3_X1 u0_u5_u5_U100 (.A3( u0_u5_u5_n141 ) , .A1( u0_u5_u5_n142 ) , .ZN( u0_u5_u5_n143 ) , .A2( u0_u5_u5_n191 ) );
  NAND4_X1 u0_u5_u5_U101 (.ZN( u0_out5_4 ) , .A4( u0_u5_u5_n112 ) , .A2( u0_u5_u5_n113 ) , .A1( u0_u5_u5_n114 ) , .A3( u0_u5_u5_n195 ) );
  AOI211_X1 u0_u5_u5_U102 (.A( u0_u5_u5_n110 ) , .C1( u0_u5_u5_n111 ) , .ZN( u0_u5_u5_n112 ) , .B( u0_u5_u5_n118 ) , .C2( u0_u5_u5_n177 ) );
  AOI222_X1 u0_u5_u5_U103 (.ZN( u0_u5_u5_n113 ) , .A1( u0_u5_u5_n131 ) , .C1( u0_u5_u5_n148 ) , .B2( u0_u5_u5_n174 ) , .C2( u0_u5_u5_n178 ) , .A2( u0_u5_u5_n179 ) , .B1( u0_u5_u5_n99 ) );
  NAND3_X1 u0_u5_u5_U104 (.A2( u0_u5_u5_n154 ) , .A3( u0_u5_u5_n158 ) , .A1( u0_u5_u5_n161 ) , .ZN( u0_u5_u5_n99 ) );
  NOR2_X1 u0_u5_u5_U11 (.ZN( u0_u5_u5_n160 ) , .A2( u0_u5_u5_n173 ) , .A1( u0_u5_u5_n177 ) );
  INV_X1 u0_u5_u5_U12 (.A( u0_u5_u5_n150 ) , .ZN( u0_u5_u5_n174 ) );
  AOI21_X1 u0_u5_u5_U13 (.A( u0_u5_u5_n160 ) , .B2( u0_u5_u5_n161 ) , .ZN( u0_u5_u5_n162 ) , .B1( u0_u5_u5_n192 ) );
  INV_X1 u0_u5_u5_U14 (.A( u0_u5_u5_n159 ) , .ZN( u0_u5_u5_n192 ) );
  AOI21_X1 u0_u5_u5_U15 (.A( u0_u5_u5_n156 ) , .B2( u0_u5_u5_n157 ) , .B1( u0_u5_u5_n158 ) , .ZN( u0_u5_u5_n163 ) );
  AOI21_X1 u0_u5_u5_U16 (.B2( u0_u5_u5_n139 ) , .B1( u0_u5_u5_n140 ) , .ZN( u0_u5_u5_n141 ) , .A( u0_u5_u5_n150 ) );
  OAI21_X1 u0_u5_u5_U17 (.A( u0_u5_u5_n133 ) , .B2( u0_u5_u5_n134 ) , .B1( u0_u5_u5_n135 ) , .ZN( u0_u5_u5_n142 ) );
  OAI21_X1 u0_u5_u5_U18 (.ZN( u0_u5_u5_n133 ) , .B2( u0_u5_u5_n147 ) , .A( u0_u5_u5_n173 ) , .B1( u0_u5_u5_n188 ) );
  NAND2_X1 u0_u5_u5_U19 (.A2( u0_u5_u5_n119 ) , .A1( u0_u5_u5_n123 ) , .ZN( u0_u5_u5_n137 ) );
  INV_X1 u0_u5_u5_U20 (.A( u0_u5_u5_n155 ) , .ZN( u0_u5_u5_n194 ) );
  NAND2_X1 u0_u5_u5_U21 (.A1( u0_u5_u5_n121 ) , .ZN( u0_u5_u5_n132 ) , .A2( u0_u5_u5_n172 ) );
  NAND2_X1 u0_u5_u5_U22 (.A2( u0_u5_u5_n122 ) , .ZN( u0_u5_u5_n136 ) , .A1( u0_u5_u5_n154 ) );
  NAND2_X1 u0_u5_u5_U23 (.A2( u0_u5_u5_n119 ) , .A1( u0_u5_u5_n120 ) , .ZN( u0_u5_u5_n159 ) );
  INV_X1 u0_u5_u5_U24 (.A( u0_u5_u5_n156 ) , .ZN( u0_u5_u5_n175 ) );
  INV_X1 u0_u5_u5_U25 (.A( u0_u5_u5_n158 ) , .ZN( u0_u5_u5_n188 ) );
  INV_X1 u0_u5_u5_U26 (.A( u0_u5_u5_n152 ) , .ZN( u0_u5_u5_n179 ) );
  INV_X1 u0_u5_u5_U27 (.A( u0_u5_u5_n140 ) , .ZN( u0_u5_u5_n182 ) );
  INV_X1 u0_u5_u5_U28 (.A( u0_u5_u5_n151 ) , .ZN( u0_u5_u5_n183 ) );
  INV_X1 u0_u5_u5_U29 (.A( u0_u5_u5_n123 ) , .ZN( u0_u5_u5_n185 ) );
  NOR2_X1 u0_u5_u5_U3 (.ZN( u0_u5_u5_n134 ) , .A1( u0_u5_u5_n183 ) , .A2( u0_u5_u5_n190 ) );
  INV_X1 u0_u5_u5_U30 (.A( u0_u5_u5_n161 ) , .ZN( u0_u5_u5_n184 ) );
  INV_X1 u0_u5_u5_U31 (.A( u0_u5_u5_n139 ) , .ZN( u0_u5_u5_n189 ) );
  INV_X1 u0_u5_u5_U32 (.A( u0_u5_u5_n157 ) , .ZN( u0_u5_u5_n190 ) );
  INV_X1 u0_u5_u5_U33 (.A( u0_u5_u5_n120 ) , .ZN( u0_u5_u5_n193 ) );
  NAND2_X1 u0_u5_u5_U34 (.ZN( u0_u5_u5_n111 ) , .A1( u0_u5_u5_n140 ) , .A2( u0_u5_u5_n155 ) );
  NOR2_X1 u0_u5_u5_U35 (.ZN( u0_u5_u5_n100 ) , .A1( u0_u5_u5_n170 ) , .A2( u0_u5_u5_n180 ) );
  INV_X1 u0_u5_u5_U36 (.A( u0_u5_u5_n117 ) , .ZN( u0_u5_u5_n196 ) );
  OAI221_X1 u0_u5_u5_U37 (.A( u0_u5_u5_n116 ) , .ZN( u0_u5_u5_n117 ) , .B2( u0_u5_u5_n119 ) , .C1( u0_u5_u5_n153 ) , .C2( u0_u5_u5_n158 ) , .B1( u0_u5_u5_n172 ) );
  AOI222_X1 u0_u5_u5_U38 (.ZN( u0_u5_u5_n116 ) , .B2( u0_u5_u5_n145 ) , .C1( u0_u5_u5_n148 ) , .A2( u0_u5_u5_n174 ) , .C2( u0_u5_u5_n177 ) , .B1( u0_u5_u5_n187 ) , .A1( u0_u5_u5_n193 ) );
  INV_X1 u0_u5_u5_U39 (.A( u0_u5_u5_n115 ) , .ZN( u0_u5_u5_n187 ) );
  INV_X1 u0_u5_u5_U4 (.A( u0_u5_u5_n138 ) , .ZN( u0_u5_u5_n191 ) );
  AOI22_X1 u0_u5_u5_U40 (.B2( u0_u5_u5_n131 ) , .A2( u0_u5_u5_n146 ) , .ZN( u0_u5_u5_n169 ) , .B1( u0_u5_u5_n174 ) , .A1( u0_u5_u5_n185 ) );
  NOR2_X1 u0_u5_u5_U41 (.A1( u0_u5_u5_n146 ) , .ZN( u0_u5_u5_n150 ) , .A2( u0_u5_u5_n173 ) );
  AOI21_X1 u0_u5_u5_U42 (.A( u0_u5_u5_n118 ) , .B2( u0_u5_u5_n145 ) , .ZN( u0_u5_u5_n168 ) , .B1( u0_u5_u5_n186 ) );
  INV_X1 u0_u5_u5_U43 (.A( u0_u5_u5_n122 ) , .ZN( u0_u5_u5_n186 ) );
  NOR2_X1 u0_u5_u5_U44 (.A1( u0_u5_u5_n146 ) , .ZN( u0_u5_u5_n152 ) , .A2( u0_u5_u5_n176 ) );
  NOR2_X1 u0_u5_u5_U45 (.A1( u0_u5_u5_n115 ) , .ZN( u0_u5_u5_n118 ) , .A2( u0_u5_u5_n153 ) );
  NOR2_X1 u0_u5_u5_U46 (.A2( u0_u5_u5_n145 ) , .ZN( u0_u5_u5_n156 ) , .A1( u0_u5_u5_n174 ) );
  NOR2_X1 u0_u5_u5_U47 (.ZN( u0_u5_u5_n121 ) , .A2( u0_u5_u5_n145 ) , .A1( u0_u5_u5_n176 ) );
  AOI22_X1 u0_u5_u5_U48 (.ZN( u0_u5_u5_n114 ) , .A2( u0_u5_u5_n137 ) , .A1( u0_u5_u5_n145 ) , .B2( u0_u5_u5_n175 ) , .B1( u0_u5_u5_n193 ) );
  OAI211_X1 u0_u5_u5_U49 (.B( u0_u5_u5_n124 ) , .A( u0_u5_u5_n125 ) , .C2( u0_u5_u5_n126 ) , .C1( u0_u5_u5_n127 ) , .ZN( u0_u5_u5_n128 ) );
  OAI21_X1 u0_u5_u5_U5 (.B2( u0_u5_u5_n136 ) , .B1( u0_u5_u5_n137 ) , .ZN( u0_u5_u5_n138 ) , .A( u0_u5_u5_n177 ) );
  NOR3_X1 u0_u5_u5_U50 (.ZN( u0_u5_u5_n127 ) , .A1( u0_u5_u5_n136 ) , .A3( u0_u5_u5_n148 ) , .A2( u0_u5_u5_n182 ) );
  OAI21_X1 u0_u5_u5_U51 (.ZN( u0_u5_u5_n124 ) , .A( u0_u5_u5_n177 ) , .B2( u0_u5_u5_n183 ) , .B1( u0_u5_u5_n189 ) );
  OAI21_X1 u0_u5_u5_U52 (.ZN( u0_u5_u5_n125 ) , .A( u0_u5_u5_n174 ) , .B2( u0_u5_u5_n185 ) , .B1( u0_u5_u5_n190 ) );
  AOI21_X1 u0_u5_u5_U53 (.A( u0_u5_u5_n153 ) , .B2( u0_u5_u5_n154 ) , .B1( u0_u5_u5_n155 ) , .ZN( u0_u5_u5_n164 ) );
  AOI21_X1 u0_u5_u5_U54 (.ZN( u0_u5_u5_n110 ) , .B1( u0_u5_u5_n122 ) , .B2( u0_u5_u5_n139 ) , .A( u0_u5_u5_n153 ) );
  INV_X1 u0_u5_u5_U55 (.A( u0_u5_u5_n153 ) , .ZN( u0_u5_u5_n176 ) );
  INV_X1 u0_u5_u5_U56 (.A( u0_u5_u5_n126 ) , .ZN( u0_u5_u5_n173 ) );
  AND2_X1 u0_u5_u5_U57 (.A2( u0_u5_u5_n104 ) , .A1( u0_u5_u5_n107 ) , .ZN( u0_u5_u5_n147 ) );
  AND2_X1 u0_u5_u5_U58 (.A2( u0_u5_u5_n104 ) , .A1( u0_u5_u5_n108 ) , .ZN( u0_u5_u5_n148 ) );
  NAND2_X1 u0_u5_u5_U59 (.A1( u0_u5_u5_n105 ) , .A2( u0_u5_u5_n106 ) , .ZN( u0_u5_u5_n158 ) );
  INV_X1 u0_u5_u5_U6 (.A( u0_u5_u5_n135 ) , .ZN( u0_u5_u5_n178 ) );
  NAND2_X1 u0_u5_u5_U60 (.A2( u0_u5_u5_n108 ) , .A1( u0_u5_u5_n109 ) , .ZN( u0_u5_u5_n139 ) );
  NAND2_X1 u0_u5_u5_U61 (.A1( u0_u5_u5_n106 ) , .A2( u0_u5_u5_n108 ) , .ZN( u0_u5_u5_n119 ) );
  NAND2_X1 u0_u5_u5_U62 (.A2( u0_u5_u5_n103 ) , .A1( u0_u5_u5_n105 ) , .ZN( u0_u5_u5_n140 ) );
  NAND2_X1 u0_u5_u5_U63 (.A2( u0_u5_u5_n104 ) , .A1( u0_u5_u5_n105 ) , .ZN( u0_u5_u5_n155 ) );
  NAND2_X1 u0_u5_u5_U64 (.A2( u0_u5_u5_n106 ) , .A1( u0_u5_u5_n107 ) , .ZN( u0_u5_u5_n122 ) );
  NAND2_X1 u0_u5_u5_U65 (.A2( u0_u5_u5_n100 ) , .A1( u0_u5_u5_n106 ) , .ZN( u0_u5_u5_n115 ) );
  NAND2_X1 u0_u5_u5_U66 (.A2( u0_u5_u5_n100 ) , .A1( u0_u5_u5_n103 ) , .ZN( u0_u5_u5_n161 ) );
  NAND2_X1 u0_u5_u5_U67 (.A1( u0_u5_u5_n105 ) , .A2( u0_u5_u5_n109 ) , .ZN( u0_u5_u5_n154 ) );
  INV_X1 u0_u5_u5_U68 (.A( u0_u5_u5_n146 ) , .ZN( u0_u5_u5_n172 ) );
  NAND2_X1 u0_u5_u5_U69 (.A1( u0_u5_u5_n103 ) , .A2( u0_u5_u5_n108 ) , .ZN( u0_u5_u5_n123 ) );
  OAI22_X1 u0_u5_u5_U7 (.B2( u0_u5_u5_n149 ) , .B1( u0_u5_u5_n150 ) , .A2( u0_u5_u5_n151 ) , .A1( u0_u5_u5_n152 ) , .ZN( u0_u5_u5_n165 ) );
  NAND2_X1 u0_u5_u5_U70 (.A2( u0_u5_u5_n103 ) , .A1( u0_u5_u5_n107 ) , .ZN( u0_u5_u5_n151 ) );
  NAND2_X1 u0_u5_u5_U71 (.A2( u0_u5_u5_n107 ) , .A1( u0_u5_u5_n109 ) , .ZN( u0_u5_u5_n120 ) );
  NAND2_X1 u0_u5_u5_U72 (.A2( u0_u5_u5_n100 ) , .A1( u0_u5_u5_n109 ) , .ZN( u0_u5_u5_n157 ) );
  AND2_X1 u0_u5_u5_U73 (.A2( u0_u5_u5_n100 ) , .A1( u0_u5_u5_n104 ) , .ZN( u0_u5_u5_n131 ) );
  INV_X1 u0_u5_u5_U74 (.A( u0_u5_u5_n102 ) , .ZN( u0_u5_u5_n195 ) );
  OAI221_X1 u0_u5_u5_U75 (.A( u0_u5_u5_n101 ) , .ZN( u0_u5_u5_n102 ) , .C2( u0_u5_u5_n115 ) , .C1( u0_u5_u5_n126 ) , .B1( u0_u5_u5_n134 ) , .B2( u0_u5_u5_n160 ) );
  OAI21_X1 u0_u5_u5_U76 (.ZN( u0_u5_u5_n101 ) , .B1( u0_u5_u5_n137 ) , .A( u0_u5_u5_n146 ) , .B2( u0_u5_u5_n147 ) );
  NOR2_X1 u0_u5_u5_U77 (.A2( u0_u5_X_34 ) , .A1( u0_u5_X_35 ) , .ZN( u0_u5_u5_n145 ) );
  NOR2_X1 u0_u5_u5_U78 (.A2( u0_u5_X_34 ) , .ZN( u0_u5_u5_n146 ) , .A1( u0_u5_u5_n171 ) );
  NOR2_X1 u0_u5_u5_U79 (.A2( u0_u5_X_31 ) , .A1( u0_u5_X_32 ) , .ZN( u0_u5_u5_n103 ) );
  NOR3_X1 u0_u5_u5_U8 (.A2( u0_u5_u5_n147 ) , .A1( u0_u5_u5_n148 ) , .ZN( u0_u5_u5_n149 ) , .A3( u0_u5_u5_n194 ) );
  NOR2_X1 u0_u5_u5_U80 (.A2( u0_u5_X_36 ) , .ZN( u0_u5_u5_n105 ) , .A1( u0_u5_u5_n180 ) );
  NOR2_X1 u0_u5_u5_U81 (.A2( u0_u5_X_33 ) , .ZN( u0_u5_u5_n108 ) , .A1( u0_u5_u5_n170 ) );
  NOR2_X1 u0_u5_u5_U82 (.A2( u0_u5_X_33 ) , .A1( u0_u5_X_36 ) , .ZN( u0_u5_u5_n107 ) );
  NOR2_X1 u0_u5_u5_U83 (.A2( u0_u5_X_31 ) , .ZN( u0_u5_u5_n104 ) , .A1( u0_u5_u5_n181 ) );
  NAND2_X1 u0_u5_u5_U84 (.A2( u0_u5_X_34 ) , .A1( u0_u5_X_35 ) , .ZN( u0_u5_u5_n153 ) );
  NAND2_X1 u0_u5_u5_U85 (.A1( u0_u5_X_34 ) , .ZN( u0_u5_u5_n126 ) , .A2( u0_u5_u5_n171 ) );
  AND2_X1 u0_u5_u5_U86 (.A1( u0_u5_X_31 ) , .A2( u0_u5_X_32 ) , .ZN( u0_u5_u5_n106 ) );
  AND2_X1 u0_u5_u5_U87 (.A1( u0_u5_X_31 ) , .ZN( u0_u5_u5_n109 ) , .A2( u0_u5_u5_n181 ) );
  INV_X1 u0_u5_u5_U88 (.A( u0_u5_X_33 ) , .ZN( u0_u5_u5_n180 ) );
  INV_X1 u0_u5_u5_U89 (.A( u0_u5_X_35 ) , .ZN( u0_u5_u5_n171 ) );
  NOR2_X1 u0_u5_u5_U9 (.ZN( u0_u5_u5_n135 ) , .A1( u0_u5_u5_n173 ) , .A2( u0_u5_u5_n176 ) );
  INV_X1 u0_u5_u5_U90 (.A( u0_u5_X_36 ) , .ZN( u0_u5_u5_n170 ) );
  INV_X1 u0_u5_u5_U91 (.A( u0_u5_X_32 ) , .ZN( u0_u5_u5_n181 ) );
  NAND4_X1 u0_u5_u5_U92 (.ZN( u0_out5_29 ) , .A4( u0_u5_u5_n129 ) , .A3( u0_u5_u5_n130 ) , .A2( u0_u5_u5_n168 ) , .A1( u0_u5_u5_n196 ) );
  AOI221_X1 u0_u5_u5_U93 (.A( u0_u5_u5_n128 ) , .ZN( u0_u5_u5_n129 ) , .C2( u0_u5_u5_n132 ) , .B2( u0_u5_u5_n159 ) , .B1( u0_u5_u5_n176 ) , .C1( u0_u5_u5_n184 ) );
  AOI222_X1 u0_u5_u5_U94 (.ZN( u0_u5_u5_n130 ) , .A2( u0_u5_u5_n146 ) , .B1( u0_u5_u5_n147 ) , .C2( u0_u5_u5_n175 ) , .B2( u0_u5_u5_n179 ) , .A1( u0_u5_u5_n188 ) , .C1( u0_u5_u5_n194 ) );
  NAND4_X1 u0_u5_u5_U95 (.ZN( u0_out5_19 ) , .A4( u0_u5_u5_n166 ) , .A3( u0_u5_u5_n167 ) , .A2( u0_u5_u5_n168 ) , .A1( u0_u5_u5_n169 ) );
  AOI22_X1 u0_u5_u5_U96 (.B2( u0_u5_u5_n145 ) , .A2( u0_u5_u5_n146 ) , .ZN( u0_u5_u5_n167 ) , .B1( u0_u5_u5_n182 ) , .A1( u0_u5_u5_n189 ) );
  NOR4_X1 u0_u5_u5_U97 (.A4( u0_u5_u5_n162 ) , .A3( u0_u5_u5_n163 ) , .A2( u0_u5_u5_n164 ) , .A1( u0_u5_u5_n165 ) , .ZN( u0_u5_u5_n166 ) );
  NAND4_X1 u0_u5_u5_U98 (.ZN( u0_out5_11 ) , .A4( u0_u5_u5_n143 ) , .A3( u0_u5_u5_n144 ) , .A2( u0_u5_u5_n169 ) , .A1( u0_u5_u5_n196 ) );
  AOI22_X1 u0_u5_u5_U99 (.A2( u0_u5_u5_n132 ) , .ZN( u0_u5_u5_n144 ) , .B2( u0_u5_u5_n145 ) , .B1( u0_u5_u5_n184 ) , .A1( u0_u5_u5_n194 ) );
  AND3_X1 u0_u5_u7_U10 (.A3( u0_u5_u7_n110 ) , .A2( u0_u5_u7_n127 ) , .A1( u0_u5_u7_n132 ) , .ZN( u0_u5_u7_n92 ) );
  OAI21_X1 u0_u5_u7_U11 (.A( u0_u5_u7_n161 ) , .B1( u0_u5_u7_n168 ) , .B2( u0_u5_u7_n173 ) , .ZN( u0_u5_u7_n91 ) );
  AOI211_X1 u0_u5_u7_U12 (.A( u0_u5_u7_n117 ) , .ZN( u0_u5_u7_n118 ) , .C2( u0_u5_u7_n126 ) , .C1( u0_u5_u7_n177 ) , .B( u0_u5_u7_n180 ) );
  OAI22_X1 u0_u5_u7_U13 (.B1( u0_u5_u7_n115 ) , .ZN( u0_u5_u7_n117 ) , .A2( u0_u5_u7_n133 ) , .A1( u0_u5_u7_n137 ) , .B2( u0_u5_u7_n162 ) );
  INV_X1 u0_u5_u7_U14 (.A( u0_u5_u7_n116 ) , .ZN( u0_u5_u7_n180 ) );
  NOR3_X1 u0_u5_u7_U15 (.ZN( u0_u5_u7_n115 ) , .A3( u0_u5_u7_n145 ) , .A2( u0_u5_u7_n168 ) , .A1( u0_u5_u7_n169 ) );
  OAI211_X1 u0_u5_u7_U16 (.B( u0_u5_u7_n122 ) , .A( u0_u5_u7_n123 ) , .C2( u0_u5_u7_n124 ) , .ZN( u0_u5_u7_n154 ) , .C1( u0_u5_u7_n162 ) );
  AOI222_X1 u0_u5_u7_U17 (.ZN( u0_u5_u7_n122 ) , .C2( u0_u5_u7_n126 ) , .C1( u0_u5_u7_n145 ) , .B1( u0_u5_u7_n161 ) , .A2( u0_u5_u7_n165 ) , .B2( u0_u5_u7_n170 ) , .A1( u0_u5_u7_n176 ) );
  INV_X1 u0_u5_u7_U18 (.A( u0_u5_u7_n133 ) , .ZN( u0_u5_u7_n176 ) );
  NOR3_X1 u0_u5_u7_U19 (.A2( u0_u5_u7_n134 ) , .A1( u0_u5_u7_n135 ) , .ZN( u0_u5_u7_n136 ) , .A3( u0_u5_u7_n171 ) );
  NOR2_X1 u0_u5_u7_U20 (.A1( u0_u5_u7_n130 ) , .A2( u0_u5_u7_n134 ) , .ZN( u0_u5_u7_n153 ) );
  INV_X1 u0_u5_u7_U21 (.A( u0_u5_u7_n101 ) , .ZN( u0_u5_u7_n165 ) );
  NOR2_X1 u0_u5_u7_U22 (.ZN( u0_u5_u7_n111 ) , .A2( u0_u5_u7_n134 ) , .A1( u0_u5_u7_n169 ) );
  AOI21_X1 u0_u5_u7_U23 (.ZN( u0_u5_u7_n104 ) , .B2( u0_u5_u7_n112 ) , .B1( u0_u5_u7_n127 ) , .A( u0_u5_u7_n164 ) );
  AOI21_X1 u0_u5_u7_U24 (.ZN( u0_u5_u7_n106 ) , .B1( u0_u5_u7_n133 ) , .B2( u0_u5_u7_n146 ) , .A( u0_u5_u7_n162 ) );
  AOI21_X1 u0_u5_u7_U25 (.A( u0_u5_u7_n101 ) , .ZN( u0_u5_u7_n107 ) , .B2( u0_u5_u7_n128 ) , .B1( u0_u5_u7_n175 ) );
  INV_X1 u0_u5_u7_U26 (.A( u0_u5_u7_n138 ) , .ZN( u0_u5_u7_n171 ) );
  INV_X1 u0_u5_u7_U27 (.A( u0_u5_u7_n131 ) , .ZN( u0_u5_u7_n177 ) );
  INV_X1 u0_u5_u7_U28 (.A( u0_u5_u7_n110 ) , .ZN( u0_u5_u7_n174 ) );
  NAND2_X1 u0_u5_u7_U29 (.A1( u0_u5_u7_n129 ) , .A2( u0_u5_u7_n132 ) , .ZN( u0_u5_u7_n149 ) );
  OAI21_X1 u0_u5_u7_U3 (.ZN( u0_u5_u7_n159 ) , .A( u0_u5_u7_n165 ) , .B2( u0_u5_u7_n171 ) , .B1( u0_u5_u7_n174 ) );
  NAND2_X1 u0_u5_u7_U30 (.A1( u0_u5_u7_n113 ) , .A2( u0_u5_u7_n124 ) , .ZN( u0_u5_u7_n130 ) );
  INV_X1 u0_u5_u7_U31 (.A( u0_u5_u7_n112 ) , .ZN( u0_u5_u7_n173 ) );
  INV_X1 u0_u5_u7_U32 (.A( u0_u5_u7_n128 ) , .ZN( u0_u5_u7_n168 ) );
  INV_X1 u0_u5_u7_U33 (.A( u0_u5_u7_n148 ) , .ZN( u0_u5_u7_n169 ) );
  INV_X1 u0_u5_u7_U34 (.A( u0_u5_u7_n127 ) , .ZN( u0_u5_u7_n179 ) );
  NOR2_X1 u0_u5_u7_U35 (.ZN( u0_u5_u7_n101 ) , .A2( u0_u5_u7_n150 ) , .A1( u0_u5_u7_n156 ) );
  AOI211_X1 u0_u5_u7_U36 (.B( u0_u5_u7_n154 ) , .A( u0_u5_u7_n155 ) , .C1( u0_u5_u7_n156 ) , .ZN( u0_u5_u7_n157 ) , .C2( u0_u5_u7_n172 ) );
  INV_X1 u0_u5_u7_U37 (.A( u0_u5_u7_n153 ) , .ZN( u0_u5_u7_n172 ) );
  AOI211_X1 u0_u5_u7_U38 (.B( u0_u5_u7_n139 ) , .A( u0_u5_u7_n140 ) , .C2( u0_u5_u7_n141 ) , .ZN( u0_u5_u7_n142 ) , .C1( u0_u5_u7_n156 ) );
  NAND4_X1 u0_u5_u7_U39 (.A3( u0_u5_u7_n127 ) , .A2( u0_u5_u7_n128 ) , .A1( u0_u5_u7_n129 ) , .ZN( u0_u5_u7_n141 ) , .A4( u0_u5_u7_n147 ) );
  INV_X1 u0_u5_u7_U4 (.A( u0_u5_u7_n111 ) , .ZN( u0_u5_u7_n170 ) );
  AOI21_X1 u0_u5_u7_U40 (.A( u0_u5_u7_n137 ) , .B1( u0_u5_u7_n138 ) , .ZN( u0_u5_u7_n139 ) , .B2( u0_u5_u7_n146 ) );
  OAI22_X1 u0_u5_u7_U41 (.B1( u0_u5_u7_n136 ) , .ZN( u0_u5_u7_n140 ) , .A1( u0_u5_u7_n153 ) , .B2( u0_u5_u7_n162 ) , .A2( u0_u5_u7_n164 ) );
  AOI21_X1 u0_u5_u7_U42 (.ZN( u0_u5_u7_n123 ) , .B1( u0_u5_u7_n165 ) , .B2( u0_u5_u7_n177 ) , .A( u0_u5_u7_n97 ) );
  AOI21_X1 u0_u5_u7_U43 (.B2( u0_u5_u7_n113 ) , .B1( u0_u5_u7_n124 ) , .A( u0_u5_u7_n125 ) , .ZN( u0_u5_u7_n97 ) );
  INV_X1 u0_u5_u7_U44 (.A( u0_u5_u7_n125 ) , .ZN( u0_u5_u7_n161 ) );
  INV_X1 u0_u5_u7_U45 (.A( u0_u5_u7_n152 ) , .ZN( u0_u5_u7_n162 ) );
  AOI22_X1 u0_u5_u7_U46 (.A2( u0_u5_u7_n114 ) , .ZN( u0_u5_u7_n119 ) , .B1( u0_u5_u7_n130 ) , .A1( u0_u5_u7_n156 ) , .B2( u0_u5_u7_n165 ) );
  NAND2_X1 u0_u5_u7_U47 (.A2( u0_u5_u7_n112 ) , .ZN( u0_u5_u7_n114 ) , .A1( u0_u5_u7_n175 ) );
  AND2_X1 u0_u5_u7_U48 (.ZN( u0_u5_u7_n145 ) , .A2( u0_u5_u7_n98 ) , .A1( u0_u5_u7_n99 ) );
  NOR2_X1 u0_u5_u7_U49 (.ZN( u0_u5_u7_n137 ) , .A1( u0_u5_u7_n150 ) , .A2( u0_u5_u7_n161 ) );
  INV_X1 u0_u5_u7_U5 (.A( u0_u5_u7_n149 ) , .ZN( u0_u5_u7_n175 ) );
  AOI21_X1 u0_u5_u7_U50 (.ZN( u0_u5_u7_n105 ) , .B2( u0_u5_u7_n110 ) , .A( u0_u5_u7_n125 ) , .B1( u0_u5_u7_n147 ) );
  NAND2_X1 u0_u5_u7_U51 (.ZN( u0_u5_u7_n146 ) , .A1( u0_u5_u7_n95 ) , .A2( u0_u5_u7_n98 ) );
  NAND2_X1 u0_u5_u7_U52 (.A2( u0_u5_u7_n103 ) , .ZN( u0_u5_u7_n147 ) , .A1( u0_u5_u7_n93 ) );
  NAND2_X1 u0_u5_u7_U53 (.A1( u0_u5_u7_n103 ) , .ZN( u0_u5_u7_n127 ) , .A2( u0_u5_u7_n99 ) );
  OR2_X1 u0_u5_u7_U54 (.ZN( u0_u5_u7_n126 ) , .A2( u0_u5_u7_n152 ) , .A1( u0_u5_u7_n156 ) );
  NAND2_X1 u0_u5_u7_U55 (.A2( u0_u5_u7_n102 ) , .A1( u0_u5_u7_n103 ) , .ZN( u0_u5_u7_n133 ) );
  NAND2_X1 u0_u5_u7_U56 (.ZN( u0_u5_u7_n112 ) , .A2( u0_u5_u7_n96 ) , .A1( u0_u5_u7_n99 ) );
  NAND2_X1 u0_u5_u7_U57 (.A2( u0_u5_u7_n102 ) , .ZN( u0_u5_u7_n128 ) , .A1( u0_u5_u7_n98 ) );
  NAND2_X1 u0_u5_u7_U58 (.A1( u0_u5_u7_n100 ) , .ZN( u0_u5_u7_n113 ) , .A2( u0_u5_u7_n93 ) );
  NAND2_X1 u0_u5_u7_U59 (.A2( u0_u5_u7_n102 ) , .ZN( u0_u5_u7_n124 ) , .A1( u0_u5_u7_n96 ) );
  INV_X1 u0_u5_u7_U6 (.A( u0_u5_u7_n154 ) , .ZN( u0_u5_u7_n178 ) );
  NAND2_X1 u0_u5_u7_U60 (.ZN( u0_u5_u7_n110 ) , .A1( u0_u5_u7_n95 ) , .A2( u0_u5_u7_n96 ) );
  INV_X1 u0_u5_u7_U61 (.A( u0_u5_u7_n150 ) , .ZN( u0_u5_u7_n164 ) );
  AND2_X1 u0_u5_u7_U62 (.ZN( u0_u5_u7_n134 ) , .A1( u0_u5_u7_n93 ) , .A2( u0_u5_u7_n98 ) );
  NAND2_X1 u0_u5_u7_U63 (.A1( u0_u5_u7_n100 ) , .A2( u0_u5_u7_n102 ) , .ZN( u0_u5_u7_n129 ) );
  NAND2_X1 u0_u5_u7_U64 (.A2( u0_u5_u7_n103 ) , .ZN( u0_u5_u7_n131 ) , .A1( u0_u5_u7_n95 ) );
  NAND2_X1 u0_u5_u7_U65 (.A1( u0_u5_u7_n100 ) , .ZN( u0_u5_u7_n138 ) , .A2( u0_u5_u7_n99 ) );
  NAND2_X1 u0_u5_u7_U66 (.ZN( u0_u5_u7_n132 ) , .A1( u0_u5_u7_n93 ) , .A2( u0_u5_u7_n96 ) );
  NAND2_X1 u0_u5_u7_U67 (.A1( u0_u5_u7_n100 ) , .ZN( u0_u5_u7_n148 ) , .A2( u0_u5_u7_n95 ) );
  NOR2_X1 u0_u5_u7_U68 (.A2( u0_u5_X_47 ) , .ZN( u0_u5_u7_n150 ) , .A1( u0_u5_u7_n163 ) );
  NOR2_X1 u0_u5_u7_U69 (.A2( u0_u5_X_43 ) , .A1( u0_u5_X_44 ) , .ZN( u0_u5_u7_n103 ) );
  AOI211_X1 u0_u5_u7_U7 (.ZN( u0_u5_u7_n116 ) , .A( u0_u5_u7_n155 ) , .C1( u0_u5_u7_n161 ) , .C2( u0_u5_u7_n171 ) , .B( u0_u5_u7_n94 ) );
  NOR2_X1 u0_u5_u7_U70 (.A2( u0_u5_X_48 ) , .A1( u0_u5_u7_n166 ) , .ZN( u0_u5_u7_n95 ) );
  NOR2_X1 u0_u5_u7_U71 (.A2( u0_u5_X_45 ) , .A1( u0_u5_X_48 ) , .ZN( u0_u5_u7_n99 ) );
  NOR2_X1 u0_u5_u7_U72 (.A2( u0_u5_X_44 ) , .A1( u0_u5_u7_n167 ) , .ZN( u0_u5_u7_n98 ) );
  NOR2_X1 u0_u5_u7_U73 (.A2( u0_u5_X_46 ) , .A1( u0_u5_X_47 ) , .ZN( u0_u5_u7_n152 ) );
  AND2_X1 u0_u5_u7_U74 (.A1( u0_u5_X_47 ) , .ZN( u0_u5_u7_n156 ) , .A2( u0_u5_u7_n163 ) );
  NAND2_X1 u0_u5_u7_U75 (.A2( u0_u5_X_46 ) , .A1( u0_u5_X_47 ) , .ZN( u0_u5_u7_n125 ) );
  AND2_X1 u0_u5_u7_U76 (.A2( u0_u5_X_45 ) , .A1( u0_u5_X_48 ) , .ZN( u0_u5_u7_n102 ) );
  AND2_X1 u0_u5_u7_U77 (.A2( u0_u5_X_43 ) , .A1( u0_u5_X_44 ) , .ZN( u0_u5_u7_n96 ) );
  AND2_X1 u0_u5_u7_U78 (.A1( u0_u5_X_44 ) , .ZN( u0_u5_u7_n100 ) , .A2( u0_u5_u7_n167 ) );
  AND2_X1 u0_u5_u7_U79 (.A1( u0_u5_X_48 ) , .A2( u0_u5_u7_n166 ) , .ZN( u0_u5_u7_n93 ) );
  OAI222_X1 u0_u5_u7_U8 (.C2( u0_u5_u7_n101 ) , .B2( u0_u5_u7_n111 ) , .A1( u0_u5_u7_n113 ) , .C1( u0_u5_u7_n146 ) , .A2( u0_u5_u7_n162 ) , .B1( u0_u5_u7_n164 ) , .ZN( u0_u5_u7_n94 ) );
  INV_X1 u0_u5_u7_U80 (.A( u0_u5_X_46 ) , .ZN( u0_u5_u7_n163 ) );
  INV_X1 u0_u5_u7_U81 (.A( u0_u5_X_43 ) , .ZN( u0_u5_u7_n167 ) );
  INV_X1 u0_u5_u7_U82 (.A( u0_u5_X_45 ) , .ZN( u0_u5_u7_n166 ) );
  NAND4_X1 u0_u5_u7_U83 (.ZN( u0_out5_27 ) , .A4( u0_u5_u7_n118 ) , .A3( u0_u5_u7_n119 ) , .A2( u0_u5_u7_n120 ) , .A1( u0_u5_u7_n121 ) );
  OAI21_X1 u0_u5_u7_U84 (.ZN( u0_u5_u7_n121 ) , .B2( u0_u5_u7_n145 ) , .A( u0_u5_u7_n150 ) , .B1( u0_u5_u7_n174 ) );
  OAI21_X1 u0_u5_u7_U85 (.ZN( u0_u5_u7_n120 ) , .A( u0_u5_u7_n161 ) , .B2( u0_u5_u7_n170 ) , .B1( u0_u5_u7_n179 ) );
  NAND4_X1 u0_u5_u7_U86 (.ZN( u0_out5_21 ) , .A4( u0_u5_u7_n157 ) , .A3( u0_u5_u7_n158 ) , .A2( u0_u5_u7_n159 ) , .A1( u0_u5_u7_n160 ) );
  OAI21_X1 u0_u5_u7_U87 (.B1( u0_u5_u7_n145 ) , .ZN( u0_u5_u7_n160 ) , .A( u0_u5_u7_n161 ) , .B2( u0_u5_u7_n177 ) );
  AOI22_X1 u0_u5_u7_U88 (.B2( u0_u5_u7_n149 ) , .B1( u0_u5_u7_n150 ) , .A2( u0_u5_u7_n151 ) , .A1( u0_u5_u7_n152 ) , .ZN( u0_u5_u7_n158 ) );
  NAND4_X1 u0_u5_u7_U89 (.ZN( u0_out5_15 ) , .A4( u0_u5_u7_n142 ) , .A3( u0_u5_u7_n143 ) , .A2( u0_u5_u7_n144 ) , .A1( u0_u5_u7_n178 ) );
  OAI221_X1 u0_u5_u7_U9 (.C1( u0_u5_u7_n101 ) , .C2( u0_u5_u7_n147 ) , .ZN( u0_u5_u7_n155 ) , .B2( u0_u5_u7_n162 ) , .A( u0_u5_u7_n91 ) , .B1( u0_u5_u7_n92 ) );
  OR2_X1 u0_u5_u7_U90 (.A2( u0_u5_u7_n125 ) , .A1( u0_u5_u7_n129 ) , .ZN( u0_u5_u7_n144 ) );
  AOI22_X1 u0_u5_u7_U91 (.A2( u0_u5_u7_n126 ) , .ZN( u0_u5_u7_n143 ) , .B2( u0_u5_u7_n165 ) , .B1( u0_u5_u7_n173 ) , .A1( u0_u5_u7_n174 ) );
  NAND4_X1 u0_u5_u7_U92 (.ZN( u0_out5_5 ) , .A4( u0_u5_u7_n108 ) , .A3( u0_u5_u7_n109 ) , .A1( u0_u5_u7_n116 ) , .A2( u0_u5_u7_n123 ) );
  AOI22_X1 u0_u5_u7_U93 (.ZN( u0_u5_u7_n109 ) , .A2( u0_u5_u7_n126 ) , .B2( u0_u5_u7_n145 ) , .B1( u0_u5_u7_n156 ) , .A1( u0_u5_u7_n171 ) );
  NOR4_X1 u0_u5_u7_U94 (.A4( u0_u5_u7_n104 ) , .A3( u0_u5_u7_n105 ) , .A2( u0_u5_u7_n106 ) , .A1( u0_u5_u7_n107 ) , .ZN( u0_u5_u7_n108 ) );
  NAND3_X1 u0_u5_u7_U95 (.A3( u0_u5_u7_n146 ) , .A2( u0_u5_u7_n147 ) , .A1( u0_u5_u7_n148 ) , .ZN( u0_u5_u7_n151 ) );
  NAND3_X1 u0_u5_u7_U96 (.A3( u0_u5_u7_n131 ) , .A2( u0_u5_u7_n132 ) , .A1( u0_u5_u7_n133 ) , .ZN( u0_u5_u7_n135 ) );
  XOR2_X1 u0_u7_U1 (.B( u0_K8_9 ) , .A( u0_R6_6 ) , .Z( u0_u7_X_9 ) );
  XOR2_X1 u0_u7_U10 (.B( u0_K8_45 ) , .A( u0_R6_30 ) , .Z( u0_u7_X_45 ) );
  XOR2_X1 u0_u7_U11 (.B( u0_K8_44 ) , .A( u0_R6_29 ) , .Z( u0_u7_X_44 ) );
  XOR2_X1 u0_u7_U12 (.B( u0_K8_43 ) , .A( u0_R6_28 ) , .Z( u0_u7_X_43 ) );
  XOR2_X1 u0_u7_U13 (.B( u0_K8_42 ) , .A( u0_R6_29 ) , .Z( u0_u7_X_42 ) );
  XOR2_X1 u0_u7_U14 (.B( u0_K8_41 ) , .A( u0_R6_28 ) , .Z( u0_u7_X_41 ) );
  XOR2_X1 u0_u7_U15 (.B( u0_K8_40 ) , .A( u0_R6_27 ) , .Z( u0_u7_X_40 ) );
  XOR2_X1 u0_u7_U16 (.B( u0_K8_3 ) , .A( u0_R6_2 ) , .Z( u0_u7_X_3 ) );
  XOR2_X1 u0_u7_U17 (.B( u0_K8_39 ) , .A( u0_R6_26 ) , .Z( u0_u7_X_39 ) );
  XOR2_X1 u0_u7_U18 (.B( u0_K8_38 ) , .A( u0_R6_25 ) , .Z( u0_u7_X_38 ) );
  XOR2_X1 u0_u7_U19 (.B( u0_K8_37 ) , .A( u0_R6_24 ) , .Z( u0_u7_X_37 ) );
  XOR2_X1 u0_u7_U2 (.B( u0_K8_8 ) , .A( u0_R6_5 ) , .Z( u0_u7_X_8 ) );
  XOR2_X1 u0_u7_U20 (.B( u0_K8_36 ) , .A( u0_R6_25 ) , .Z( u0_u7_X_36 ) );
  XOR2_X1 u0_u7_U21 (.B( u0_K8_35 ) , .A( u0_R6_24 ) , .Z( u0_u7_X_35 ) );
  XOR2_X1 u0_u7_U22 (.B( u0_K8_34 ) , .A( u0_R6_23 ) , .Z( u0_u7_X_34 ) );
  XOR2_X1 u0_u7_U23 (.B( u0_K8_33 ) , .A( u0_R6_22 ) , .Z( u0_u7_X_33 ) );
  XOR2_X1 u0_u7_U24 (.B( u0_K8_32 ) , .A( u0_R6_21 ) , .Z( u0_u7_X_32 ) );
  XOR2_X1 u0_u7_U25 (.B( u0_K8_31 ) , .A( u0_R6_20 ) , .Z( u0_u7_X_31 ) );
  XOR2_X1 u0_u7_U26 (.B( u0_K8_30 ) , .A( u0_R6_21 ) , .Z( u0_u7_X_30 ) );
  XOR2_X1 u0_u7_U27 (.B( u0_K8_2 ) , .A( u0_R6_1 ) , .Z( u0_u7_X_2 ) );
  XOR2_X1 u0_u7_U28 (.B( u0_K8_29 ) , .A( u0_R6_20 ) , .Z( u0_u7_X_29 ) );
  XOR2_X1 u0_u7_U29 (.B( u0_K8_28 ) , .A( u0_R6_19 ) , .Z( u0_u7_X_28 ) );
  XOR2_X1 u0_u7_U3 (.B( u0_K8_7 ) , .A( u0_R6_4 ) , .Z( u0_u7_X_7 ) );
  XOR2_X1 u0_u7_U30 (.B( u0_K8_27 ) , .A( u0_R6_18 ) , .Z( u0_u7_X_27 ) );
  XOR2_X1 u0_u7_U31 (.B( u0_K8_26 ) , .A( u0_R6_17 ) , .Z( u0_u7_X_26 ) );
  XOR2_X1 u0_u7_U32 (.B( u0_K8_25 ) , .A( u0_R6_16 ) , .Z( u0_u7_X_25 ) );
  XOR2_X1 u0_u7_U33 (.B( u0_K8_24 ) , .A( u0_R6_17 ) , .Z( u0_u7_X_24 ) );
  XOR2_X1 u0_u7_U34 (.B( u0_K8_23 ) , .A( u0_R6_16 ) , .Z( u0_u7_X_23 ) );
  XOR2_X1 u0_u7_U35 (.B( u0_K8_22 ) , .A( u0_R6_15 ) , .Z( u0_u7_X_22 ) );
  XOR2_X1 u0_u7_U36 (.B( u0_K8_21 ) , .A( u0_R6_14 ) , .Z( u0_u7_X_21 ) );
  XOR2_X1 u0_u7_U37 (.B( u0_K8_20 ) , .A( u0_R6_13 ) , .Z( u0_u7_X_20 ) );
  XOR2_X1 u0_u7_U38 (.B( u0_K8_1 ) , .A( u0_R6_32 ) , .Z( u0_u7_X_1 ) );
  XOR2_X1 u0_u7_U39 (.B( u0_K8_19 ) , .A( u0_R6_12 ) , .Z( u0_u7_X_19 ) );
  XOR2_X1 u0_u7_U4 (.B( u0_K8_6 ) , .A( u0_R6_5 ) , .Z( u0_u7_X_6 ) );
  XOR2_X1 u0_u7_U40 (.B( u0_K8_18 ) , .A( u0_R6_13 ) , .Z( u0_u7_X_18 ) );
  XOR2_X1 u0_u7_U41 (.B( u0_K8_17 ) , .A( u0_R6_12 ) , .Z( u0_u7_X_17 ) );
  XOR2_X1 u0_u7_U42 (.B( u0_K8_16 ) , .A( u0_R6_11 ) , .Z( u0_u7_X_16 ) );
  XOR2_X1 u0_u7_U43 (.B( u0_K8_15 ) , .A( u0_R6_10 ) , .Z( u0_u7_X_15 ) );
  XOR2_X1 u0_u7_U44 (.B( u0_K8_14 ) , .A( u0_R6_9 ) , .Z( u0_u7_X_14 ) );
  XOR2_X1 u0_u7_U45 (.B( u0_K8_13 ) , .A( u0_R6_8 ) , .Z( u0_u7_X_13 ) );
  XOR2_X1 u0_u7_U46 (.B( u0_K8_12 ) , .A( u0_R6_9 ) , .Z( u0_u7_X_12 ) );
  XOR2_X1 u0_u7_U47 (.B( u0_K8_11 ) , .A( u0_R6_8 ) , .Z( u0_u7_X_11 ) );
  XOR2_X1 u0_u7_U48 (.B( u0_K8_10 ) , .A( u0_R6_7 ) , .Z( u0_u7_X_10 ) );
  XOR2_X1 u0_u7_U5 (.B( u0_K8_5 ) , .A( u0_R6_4 ) , .Z( u0_u7_X_5 ) );
  XOR2_X1 u0_u7_U6 (.B( u0_K8_4 ) , .A( u0_R6_3 ) , .Z( u0_u7_X_4 ) );
  XOR2_X1 u0_u7_U7 (.B( u0_K8_48 ) , .A( u0_R6_1 ) , .Z( u0_u7_X_48 ) );
  XOR2_X1 u0_u7_U8 (.B( u0_K8_47 ) , .A( u0_R6_32 ) , .Z( u0_u7_X_47 ) );
  XOR2_X1 u0_u7_U9 (.B( u0_K8_46 ) , .A( u0_R6_31 ) , .Z( u0_u7_X_46 ) );
  AND3_X1 u0_u7_u0_U10 (.A2( u0_u7_u0_n112 ) , .ZN( u0_u7_u0_n127 ) , .A3( u0_u7_u0_n130 ) , .A1( u0_u7_u0_n148 ) );
  NAND2_X1 u0_u7_u0_U11 (.ZN( u0_u7_u0_n113 ) , .A1( u0_u7_u0_n139 ) , .A2( u0_u7_u0_n149 ) );
  AND2_X1 u0_u7_u0_U12 (.ZN( u0_u7_u0_n107 ) , .A1( u0_u7_u0_n130 ) , .A2( u0_u7_u0_n140 ) );
  AND2_X1 u0_u7_u0_U13 (.A2( u0_u7_u0_n129 ) , .A1( u0_u7_u0_n130 ) , .ZN( u0_u7_u0_n151 ) );
  AND2_X1 u0_u7_u0_U14 (.A1( u0_u7_u0_n108 ) , .A2( u0_u7_u0_n125 ) , .ZN( u0_u7_u0_n145 ) );
  INV_X1 u0_u7_u0_U15 (.A( u0_u7_u0_n143 ) , .ZN( u0_u7_u0_n173 ) );
  NOR2_X1 u0_u7_u0_U16 (.A2( u0_u7_u0_n136 ) , .ZN( u0_u7_u0_n147 ) , .A1( u0_u7_u0_n160 ) );
  INV_X1 u0_u7_u0_U17 (.ZN( u0_u7_u0_n172 ) , .A( u0_u7_u0_n88 ) );
  OAI222_X1 u0_u7_u0_U18 (.C1( u0_u7_u0_n108 ) , .A1( u0_u7_u0_n125 ) , .B2( u0_u7_u0_n128 ) , .B1( u0_u7_u0_n144 ) , .A2( u0_u7_u0_n158 ) , .C2( u0_u7_u0_n161 ) , .ZN( u0_u7_u0_n88 ) );
  NOR2_X1 u0_u7_u0_U19 (.A1( u0_u7_u0_n163 ) , .A2( u0_u7_u0_n164 ) , .ZN( u0_u7_u0_n95 ) );
  AOI21_X1 u0_u7_u0_U20 (.B1( u0_u7_u0_n103 ) , .ZN( u0_u7_u0_n132 ) , .A( u0_u7_u0_n165 ) , .B2( u0_u7_u0_n93 ) );
  INV_X1 u0_u7_u0_U21 (.A( u0_u7_u0_n142 ) , .ZN( u0_u7_u0_n165 ) );
  OAI22_X1 u0_u7_u0_U22 (.B1( u0_u7_u0_n125 ) , .ZN( u0_u7_u0_n126 ) , .A1( u0_u7_u0_n138 ) , .A2( u0_u7_u0_n146 ) , .B2( u0_u7_u0_n147 ) );
  OAI22_X1 u0_u7_u0_U23 (.B1( u0_u7_u0_n131 ) , .A1( u0_u7_u0_n144 ) , .B2( u0_u7_u0_n147 ) , .A2( u0_u7_u0_n90 ) , .ZN( u0_u7_u0_n91 ) );
  AND3_X1 u0_u7_u0_U24 (.A3( u0_u7_u0_n121 ) , .A2( u0_u7_u0_n125 ) , .A1( u0_u7_u0_n148 ) , .ZN( u0_u7_u0_n90 ) );
  NAND2_X1 u0_u7_u0_U25 (.A1( u0_u7_u0_n100 ) , .A2( u0_u7_u0_n103 ) , .ZN( u0_u7_u0_n125 ) );
  INV_X1 u0_u7_u0_U26 (.A( u0_u7_u0_n136 ) , .ZN( u0_u7_u0_n161 ) );
  AOI22_X1 u0_u7_u0_U27 (.B2( u0_u7_u0_n109 ) , .A2( u0_u7_u0_n110 ) , .ZN( u0_u7_u0_n111 ) , .B1( u0_u7_u0_n118 ) , .A1( u0_u7_u0_n160 ) );
  NAND2_X1 u0_u7_u0_U28 (.A1( u0_u7_u0_n100 ) , .ZN( u0_u7_u0_n129 ) , .A2( u0_u7_u0_n95 ) );
  INV_X1 u0_u7_u0_U29 (.A( u0_u7_u0_n118 ) , .ZN( u0_u7_u0_n158 ) );
  INV_X1 u0_u7_u0_U3 (.A( u0_u7_u0_n113 ) , .ZN( u0_u7_u0_n166 ) );
  AOI21_X1 u0_u7_u0_U30 (.ZN( u0_u7_u0_n104 ) , .B1( u0_u7_u0_n107 ) , .B2( u0_u7_u0_n141 ) , .A( u0_u7_u0_n144 ) );
  AOI21_X1 u0_u7_u0_U31 (.B1( u0_u7_u0_n127 ) , .B2( u0_u7_u0_n129 ) , .A( u0_u7_u0_n138 ) , .ZN( u0_u7_u0_n96 ) );
  AOI21_X1 u0_u7_u0_U32 (.ZN( u0_u7_u0_n116 ) , .B2( u0_u7_u0_n142 ) , .A( u0_u7_u0_n144 ) , .B1( u0_u7_u0_n166 ) );
  NOR2_X1 u0_u7_u0_U33 (.A1( u0_u7_u0_n120 ) , .ZN( u0_u7_u0_n143 ) , .A2( u0_u7_u0_n167 ) );
  OAI221_X1 u0_u7_u0_U34 (.C1( u0_u7_u0_n112 ) , .ZN( u0_u7_u0_n120 ) , .B1( u0_u7_u0_n138 ) , .B2( u0_u7_u0_n141 ) , .C2( u0_u7_u0_n147 ) , .A( u0_u7_u0_n172 ) );
  AOI211_X1 u0_u7_u0_U35 (.B( u0_u7_u0_n115 ) , .A( u0_u7_u0_n116 ) , .C2( u0_u7_u0_n117 ) , .C1( u0_u7_u0_n118 ) , .ZN( u0_u7_u0_n119 ) );
  NAND2_X1 u0_u7_u0_U36 (.A2( u0_u7_u0_n100 ) , .A1( u0_u7_u0_n101 ) , .ZN( u0_u7_u0_n139 ) );
  NAND2_X1 u0_u7_u0_U37 (.A2( u0_u7_u0_n100 ) , .ZN( u0_u7_u0_n131 ) , .A1( u0_u7_u0_n92 ) );
  NAND2_X1 u0_u7_u0_U38 (.A1( u0_u7_u0_n101 ) , .A2( u0_u7_u0_n102 ) , .ZN( u0_u7_u0_n150 ) );
  INV_X1 u0_u7_u0_U39 (.A( u0_u7_u0_n138 ) , .ZN( u0_u7_u0_n160 ) );
  AOI21_X1 u0_u7_u0_U4 (.B1( u0_u7_u0_n114 ) , .ZN( u0_u7_u0_n115 ) , .B2( u0_u7_u0_n129 ) , .A( u0_u7_u0_n161 ) );
  NAND2_X1 u0_u7_u0_U40 (.A1( u0_u7_u0_n102 ) , .ZN( u0_u7_u0_n128 ) , .A2( u0_u7_u0_n95 ) );
  NAND2_X1 u0_u7_u0_U41 (.ZN( u0_u7_u0_n148 ) , .A1( u0_u7_u0_n93 ) , .A2( u0_u7_u0_n95 ) );
  NAND2_X1 u0_u7_u0_U42 (.A2( u0_u7_u0_n102 ) , .A1( u0_u7_u0_n103 ) , .ZN( u0_u7_u0_n149 ) );
  NAND2_X1 u0_u7_u0_U43 (.A2( u0_u7_u0_n102 ) , .ZN( u0_u7_u0_n114 ) , .A1( u0_u7_u0_n92 ) );
  NAND2_X1 u0_u7_u0_U44 (.A2( u0_u7_u0_n101 ) , .ZN( u0_u7_u0_n121 ) , .A1( u0_u7_u0_n93 ) );
  NAND2_X1 u0_u7_u0_U45 (.ZN( u0_u7_u0_n112 ) , .A2( u0_u7_u0_n92 ) , .A1( u0_u7_u0_n93 ) );
  OR3_X1 u0_u7_u0_U46 (.A3( u0_u7_u0_n152 ) , .A2( u0_u7_u0_n153 ) , .A1( u0_u7_u0_n154 ) , .ZN( u0_u7_u0_n155 ) );
  AOI21_X1 u0_u7_u0_U47 (.A( u0_u7_u0_n144 ) , .B2( u0_u7_u0_n145 ) , .B1( u0_u7_u0_n146 ) , .ZN( u0_u7_u0_n154 ) );
  AOI21_X1 u0_u7_u0_U48 (.B2( u0_u7_u0_n150 ) , .B1( u0_u7_u0_n151 ) , .ZN( u0_u7_u0_n152 ) , .A( u0_u7_u0_n158 ) );
  AOI21_X1 u0_u7_u0_U49 (.A( u0_u7_u0_n147 ) , .B2( u0_u7_u0_n148 ) , .B1( u0_u7_u0_n149 ) , .ZN( u0_u7_u0_n153 ) );
  AOI21_X1 u0_u7_u0_U5 (.B2( u0_u7_u0_n131 ) , .ZN( u0_u7_u0_n134 ) , .B1( u0_u7_u0_n151 ) , .A( u0_u7_u0_n158 ) );
  INV_X1 u0_u7_u0_U50 (.ZN( u0_u7_u0_n171 ) , .A( u0_u7_u0_n99 ) );
  OAI211_X1 u0_u7_u0_U51 (.C2( u0_u7_u0_n140 ) , .C1( u0_u7_u0_n161 ) , .A( u0_u7_u0_n169 ) , .B( u0_u7_u0_n98 ) , .ZN( u0_u7_u0_n99 ) );
  INV_X1 u0_u7_u0_U52 (.ZN( u0_u7_u0_n169 ) , .A( u0_u7_u0_n91 ) );
  AOI211_X1 u0_u7_u0_U53 (.C1( u0_u7_u0_n118 ) , .A( u0_u7_u0_n123 ) , .B( u0_u7_u0_n96 ) , .C2( u0_u7_u0_n97 ) , .ZN( u0_u7_u0_n98 ) );
  NOR2_X1 u0_u7_u0_U54 (.A2( u0_u7_X_4 ) , .A1( u0_u7_X_5 ) , .ZN( u0_u7_u0_n118 ) );
  NOR2_X1 u0_u7_u0_U55 (.A2( u0_u7_X_2 ) , .ZN( u0_u7_u0_n103 ) , .A1( u0_u7_u0_n164 ) );
  NOR2_X1 u0_u7_u0_U56 (.A2( u0_u7_X_1 ) , .A1( u0_u7_X_2 ) , .ZN( u0_u7_u0_n92 ) );
  NOR2_X1 u0_u7_u0_U57 (.A2( u0_u7_X_1 ) , .ZN( u0_u7_u0_n101 ) , .A1( u0_u7_u0_n163 ) );
  NAND2_X1 u0_u7_u0_U58 (.A2( u0_u7_X_4 ) , .A1( u0_u7_X_5 ) , .ZN( u0_u7_u0_n144 ) );
  NOR2_X1 u0_u7_u0_U59 (.A2( u0_u7_X_5 ) , .ZN( u0_u7_u0_n136 ) , .A1( u0_u7_u0_n159 ) );
  NOR2_X1 u0_u7_u0_U6 (.A1( u0_u7_u0_n108 ) , .ZN( u0_u7_u0_n123 ) , .A2( u0_u7_u0_n158 ) );
  NAND2_X1 u0_u7_u0_U60 (.A1( u0_u7_X_5 ) , .ZN( u0_u7_u0_n138 ) , .A2( u0_u7_u0_n159 ) );
  NOR2_X1 u0_u7_u0_U61 (.A2( u0_u7_X_3 ) , .A1( u0_u7_X_6 ) , .ZN( u0_u7_u0_n94 ) );
  AND2_X1 u0_u7_u0_U62 (.A2( u0_u7_X_3 ) , .A1( u0_u7_X_6 ) , .ZN( u0_u7_u0_n102 ) );
  AND2_X1 u0_u7_u0_U63 (.A1( u0_u7_X_6 ) , .A2( u0_u7_u0_n162 ) , .ZN( u0_u7_u0_n93 ) );
  INV_X1 u0_u7_u0_U64 (.A( u0_u7_X_4 ) , .ZN( u0_u7_u0_n159 ) );
  INV_X1 u0_u7_u0_U65 (.A( u0_u7_X_1 ) , .ZN( u0_u7_u0_n164 ) );
  INV_X1 u0_u7_u0_U66 (.A( u0_u7_X_2 ) , .ZN( u0_u7_u0_n163 ) );
  INV_X1 u0_u7_u0_U67 (.A( u0_u7_u0_n126 ) , .ZN( u0_u7_u0_n168 ) );
  AOI211_X1 u0_u7_u0_U68 (.B( u0_u7_u0_n133 ) , .A( u0_u7_u0_n134 ) , .C2( u0_u7_u0_n135 ) , .C1( u0_u7_u0_n136 ) , .ZN( u0_u7_u0_n137 ) );
  OR4_X1 u0_u7_u0_U69 (.ZN( u0_out7_17 ) , .A4( u0_u7_u0_n122 ) , .A2( u0_u7_u0_n123 ) , .A1( u0_u7_u0_n124 ) , .A3( u0_u7_u0_n170 ) );
  OAI21_X1 u0_u7_u0_U7 (.B1( u0_u7_u0_n150 ) , .B2( u0_u7_u0_n158 ) , .A( u0_u7_u0_n172 ) , .ZN( u0_u7_u0_n89 ) );
  AOI21_X1 u0_u7_u0_U70 (.B2( u0_u7_u0_n107 ) , .ZN( u0_u7_u0_n124 ) , .B1( u0_u7_u0_n128 ) , .A( u0_u7_u0_n161 ) );
  INV_X1 u0_u7_u0_U71 (.A( u0_u7_u0_n111 ) , .ZN( u0_u7_u0_n170 ) );
  OR4_X1 u0_u7_u0_U72 (.ZN( u0_out7_31 ) , .A4( u0_u7_u0_n155 ) , .A2( u0_u7_u0_n156 ) , .A1( u0_u7_u0_n157 ) , .A3( u0_u7_u0_n173 ) );
  AOI21_X1 u0_u7_u0_U73 (.A( u0_u7_u0_n138 ) , .B2( u0_u7_u0_n139 ) , .B1( u0_u7_u0_n140 ) , .ZN( u0_u7_u0_n157 ) );
  AOI21_X1 u0_u7_u0_U74 (.B2( u0_u7_u0_n141 ) , .B1( u0_u7_u0_n142 ) , .ZN( u0_u7_u0_n156 ) , .A( u0_u7_u0_n161 ) );
  INV_X1 u0_u7_u0_U75 (.ZN( u0_u7_u0_n174 ) , .A( u0_u7_u0_n89 ) );
  AOI211_X1 u0_u7_u0_U76 (.B( u0_u7_u0_n104 ) , .A( u0_u7_u0_n105 ) , .ZN( u0_u7_u0_n106 ) , .C2( u0_u7_u0_n113 ) , .C1( u0_u7_u0_n160 ) );
  OAI221_X1 u0_u7_u0_U77 (.C1( u0_u7_u0_n121 ) , .ZN( u0_u7_u0_n122 ) , .B2( u0_u7_u0_n127 ) , .A( u0_u7_u0_n143 ) , .B1( u0_u7_u0_n144 ) , .C2( u0_u7_u0_n147 ) );
  NOR2_X1 u0_u7_u0_U78 (.A2( u0_u7_X_6 ) , .ZN( u0_u7_u0_n100 ) , .A1( u0_u7_u0_n162 ) );
  INV_X1 u0_u7_u0_U79 (.A( u0_u7_X_3 ) , .ZN( u0_u7_u0_n162 ) );
  AND2_X1 u0_u7_u0_U8 (.A1( u0_u7_u0_n114 ) , .A2( u0_u7_u0_n121 ) , .ZN( u0_u7_u0_n146 ) );
  AOI21_X1 u0_u7_u0_U80 (.B1( u0_u7_u0_n132 ) , .ZN( u0_u7_u0_n133 ) , .A( u0_u7_u0_n144 ) , .B2( u0_u7_u0_n166 ) );
  OAI22_X1 u0_u7_u0_U81 (.ZN( u0_u7_u0_n105 ) , .A2( u0_u7_u0_n132 ) , .B1( u0_u7_u0_n146 ) , .A1( u0_u7_u0_n147 ) , .B2( u0_u7_u0_n161 ) );
  NAND2_X1 u0_u7_u0_U82 (.ZN( u0_u7_u0_n110 ) , .A2( u0_u7_u0_n132 ) , .A1( u0_u7_u0_n145 ) );
  INV_X1 u0_u7_u0_U83 (.A( u0_u7_u0_n119 ) , .ZN( u0_u7_u0_n167 ) );
  NAND2_X1 u0_u7_u0_U84 (.A2( u0_u7_u0_n103 ) , .ZN( u0_u7_u0_n140 ) , .A1( u0_u7_u0_n94 ) );
  NAND2_X1 u0_u7_u0_U85 (.A1( u0_u7_u0_n101 ) , .ZN( u0_u7_u0_n130 ) , .A2( u0_u7_u0_n94 ) );
  NAND2_X1 u0_u7_u0_U86 (.ZN( u0_u7_u0_n108 ) , .A1( u0_u7_u0_n92 ) , .A2( u0_u7_u0_n94 ) );
  NAND2_X1 u0_u7_u0_U87 (.ZN( u0_u7_u0_n142 ) , .A1( u0_u7_u0_n94 ) , .A2( u0_u7_u0_n95 ) );
  NAND3_X1 u0_u7_u0_U88 (.ZN( u0_out7_23 ) , .A3( u0_u7_u0_n137 ) , .A1( u0_u7_u0_n168 ) , .A2( u0_u7_u0_n171 ) );
  NAND3_X1 u0_u7_u0_U89 (.A3( u0_u7_u0_n127 ) , .A2( u0_u7_u0_n128 ) , .ZN( u0_u7_u0_n135 ) , .A1( u0_u7_u0_n150 ) );
  AND2_X1 u0_u7_u0_U9 (.A1( u0_u7_u0_n131 ) , .ZN( u0_u7_u0_n141 ) , .A2( u0_u7_u0_n150 ) );
  NAND3_X1 u0_u7_u0_U90 (.ZN( u0_u7_u0_n117 ) , .A3( u0_u7_u0_n132 ) , .A2( u0_u7_u0_n139 ) , .A1( u0_u7_u0_n148 ) );
  NAND3_X1 u0_u7_u0_U91 (.ZN( u0_u7_u0_n109 ) , .A2( u0_u7_u0_n114 ) , .A3( u0_u7_u0_n140 ) , .A1( u0_u7_u0_n149 ) );
  NAND3_X1 u0_u7_u0_U92 (.ZN( u0_out7_9 ) , .A3( u0_u7_u0_n106 ) , .A2( u0_u7_u0_n171 ) , .A1( u0_u7_u0_n174 ) );
  NAND3_X1 u0_u7_u0_U93 (.A2( u0_u7_u0_n128 ) , .A1( u0_u7_u0_n132 ) , .A3( u0_u7_u0_n146 ) , .ZN( u0_u7_u0_n97 ) );
  AOI21_X1 u0_u7_u1_U10 (.B2( u0_u7_u1_n155 ) , .B1( u0_u7_u1_n156 ) , .ZN( u0_u7_u1_n157 ) , .A( u0_u7_u1_n174 ) );
  NAND3_X1 u0_u7_u1_U100 (.ZN( u0_u7_u1_n113 ) , .A1( u0_u7_u1_n120 ) , .A3( u0_u7_u1_n133 ) , .A2( u0_u7_u1_n155 ) );
  NAND2_X1 u0_u7_u1_U11 (.ZN( u0_u7_u1_n140 ) , .A2( u0_u7_u1_n150 ) , .A1( u0_u7_u1_n155 ) );
  NAND2_X1 u0_u7_u1_U12 (.A1( u0_u7_u1_n131 ) , .ZN( u0_u7_u1_n147 ) , .A2( u0_u7_u1_n153 ) );
  AOI22_X1 u0_u7_u1_U13 (.B2( u0_u7_u1_n136 ) , .A2( u0_u7_u1_n137 ) , .ZN( u0_u7_u1_n143 ) , .A1( u0_u7_u1_n171 ) , .B1( u0_u7_u1_n173 ) );
  INV_X1 u0_u7_u1_U14 (.A( u0_u7_u1_n147 ) , .ZN( u0_u7_u1_n181 ) );
  INV_X1 u0_u7_u1_U15 (.A( u0_u7_u1_n139 ) , .ZN( u0_u7_u1_n174 ) );
  OR4_X1 u0_u7_u1_U16 (.A4( u0_u7_u1_n106 ) , .A3( u0_u7_u1_n107 ) , .ZN( u0_u7_u1_n108 ) , .A1( u0_u7_u1_n117 ) , .A2( u0_u7_u1_n184 ) );
  AOI21_X1 u0_u7_u1_U17 (.ZN( u0_u7_u1_n106 ) , .A( u0_u7_u1_n112 ) , .B1( u0_u7_u1_n154 ) , .B2( u0_u7_u1_n156 ) );
  AOI21_X1 u0_u7_u1_U18 (.ZN( u0_u7_u1_n107 ) , .B1( u0_u7_u1_n134 ) , .B2( u0_u7_u1_n149 ) , .A( u0_u7_u1_n174 ) );
  INV_X1 u0_u7_u1_U19 (.A( u0_u7_u1_n101 ) , .ZN( u0_u7_u1_n184 ) );
  INV_X1 u0_u7_u1_U20 (.A( u0_u7_u1_n112 ) , .ZN( u0_u7_u1_n171 ) );
  NAND2_X1 u0_u7_u1_U21 (.ZN( u0_u7_u1_n141 ) , .A1( u0_u7_u1_n153 ) , .A2( u0_u7_u1_n156 ) );
  AND2_X1 u0_u7_u1_U22 (.A1( u0_u7_u1_n123 ) , .ZN( u0_u7_u1_n134 ) , .A2( u0_u7_u1_n161 ) );
  NAND2_X1 u0_u7_u1_U23 (.A2( u0_u7_u1_n115 ) , .A1( u0_u7_u1_n116 ) , .ZN( u0_u7_u1_n148 ) );
  NAND2_X1 u0_u7_u1_U24 (.A2( u0_u7_u1_n133 ) , .A1( u0_u7_u1_n135 ) , .ZN( u0_u7_u1_n159 ) );
  NAND2_X1 u0_u7_u1_U25 (.A2( u0_u7_u1_n115 ) , .A1( u0_u7_u1_n120 ) , .ZN( u0_u7_u1_n132 ) );
  INV_X1 u0_u7_u1_U26 (.A( u0_u7_u1_n154 ) , .ZN( u0_u7_u1_n178 ) );
  INV_X1 u0_u7_u1_U27 (.A( u0_u7_u1_n151 ) , .ZN( u0_u7_u1_n183 ) );
  AND2_X1 u0_u7_u1_U28 (.A1( u0_u7_u1_n129 ) , .A2( u0_u7_u1_n133 ) , .ZN( u0_u7_u1_n149 ) );
  INV_X1 u0_u7_u1_U29 (.A( u0_u7_u1_n131 ) , .ZN( u0_u7_u1_n180 ) );
  INV_X1 u0_u7_u1_U3 (.A( u0_u7_u1_n159 ) , .ZN( u0_u7_u1_n182 ) );
  OAI221_X1 u0_u7_u1_U30 (.A( u0_u7_u1_n119 ) , .C2( u0_u7_u1_n129 ) , .ZN( u0_u7_u1_n138 ) , .B2( u0_u7_u1_n152 ) , .C1( u0_u7_u1_n174 ) , .B1( u0_u7_u1_n187 ) );
  INV_X1 u0_u7_u1_U31 (.A( u0_u7_u1_n148 ) , .ZN( u0_u7_u1_n187 ) );
  AOI211_X1 u0_u7_u1_U32 (.B( u0_u7_u1_n117 ) , .A( u0_u7_u1_n118 ) , .ZN( u0_u7_u1_n119 ) , .C2( u0_u7_u1_n146 ) , .C1( u0_u7_u1_n159 ) );
  NOR2_X1 u0_u7_u1_U33 (.A1( u0_u7_u1_n168 ) , .A2( u0_u7_u1_n176 ) , .ZN( u0_u7_u1_n98 ) );
  AOI211_X1 u0_u7_u1_U34 (.B( u0_u7_u1_n162 ) , .A( u0_u7_u1_n163 ) , .C2( u0_u7_u1_n164 ) , .ZN( u0_u7_u1_n165 ) , .C1( u0_u7_u1_n171 ) );
  AOI21_X1 u0_u7_u1_U35 (.A( u0_u7_u1_n160 ) , .B2( u0_u7_u1_n161 ) , .ZN( u0_u7_u1_n162 ) , .B1( u0_u7_u1_n182 ) );
  OR2_X1 u0_u7_u1_U36 (.A2( u0_u7_u1_n157 ) , .A1( u0_u7_u1_n158 ) , .ZN( u0_u7_u1_n163 ) );
  NAND2_X1 u0_u7_u1_U37 (.A1( u0_u7_u1_n128 ) , .ZN( u0_u7_u1_n146 ) , .A2( u0_u7_u1_n160 ) );
  NAND2_X1 u0_u7_u1_U38 (.A2( u0_u7_u1_n112 ) , .ZN( u0_u7_u1_n139 ) , .A1( u0_u7_u1_n152 ) );
  NAND2_X1 u0_u7_u1_U39 (.A1( u0_u7_u1_n105 ) , .ZN( u0_u7_u1_n156 ) , .A2( u0_u7_u1_n99 ) );
  AOI221_X1 u0_u7_u1_U4 (.A( u0_u7_u1_n138 ) , .C2( u0_u7_u1_n139 ) , .C1( u0_u7_u1_n140 ) , .B2( u0_u7_u1_n141 ) , .ZN( u0_u7_u1_n142 ) , .B1( u0_u7_u1_n175 ) );
  AOI221_X1 u0_u7_u1_U40 (.B1( u0_u7_u1_n140 ) , .ZN( u0_u7_u1_n167 ) , .B2( u0_u7_u1_n172 ) , .C2( u0_u7_u1_n175 ) , .C1( u0_u7_u1_n178 ) , .A( u0_u7_u1_n188 ) );
  INV_X1 u0_u7_u1_U41 (.ZN( u0_u7_u1_n188 ) , .A( u0_u7_u1_n97 ) );
  AOI211_X1 u0_u7_u1_U42 (.A( u0_u7_u1_n118 ) , .C1( u0_u7_u1_n132 ) , .C2( u0_u7_u1_n139 ) , .B( u0_u7_u1_n96 ) , .ZN( u0_u7_u1_n97 ) );
  AOI21_X1 u0_u7_u1_U43 (.B2( u0_u7_u1_n121 ) , .B1( u0_u7_u1_n135 ) , .A( u0_u7_u1_n152 ) , .ZN( u0_u7_u1_n96 ) );
  NOR2_X1 u0_u7_u1_U44 (.ZN( u0_u7_u1_n117 ) , .A1( u0_u7_u1_n121 ) , .A2( u0_u7_u1_n160 ) );
  OAI21_X1 u0_u7_u1_U45 (.B2( u0_u7_u1_n123 ) , .ZN( u0_u7_u1_n145 ) , .B1( u0_u7_u1_n160 ) , .A( u0_u7_u1_n185 ) );
  INV_X1 u0_u7_u1_U46 (.A( u0_u7_u1_n122 ) , .ZN( u0_u7_u1_n185 ) );
  AOI21_X1 u0_u7_u1_U47 (.B2( u0_u7_u1_n120 ) , .B1( u0_u7_u1_n121 ) , .ZN( u0_u7_u1_n122 ) , .A( u0_u7_u1_n128 ) );
  AOI21_X1 u0_u7_u1_U48 (.A( u0_u7_u1_n128 ) , .B2( u0_u7_u1_n129 ) , .ZN( u0_u7_u1_n130 ) , .B1( u0_u7_u1_n150 ) );
  NAND2_X1 u0_u7_u1_U49 (.ZN( u0_u7_u1_n112 ) , .A1( u0_u7_u1_n169 ) , .A2( u0_u7_u1_n170 ) );
  AOI211_X1 u0_u7_u1_U5 (.ZN( u0_u7_u1_n124 ) , .A( u0_u7_u1_n138 ) , .C2( u0_u7_u1_n139 ) , .B( u0_u7_u1_n145 ) , .C1( u0_u7_u1_n147 ) );
  NAND2_X1 u0_u7_u1_U50 (.ZN( u0_u7_u1_n129 ) , .A2( u0_u7_u1_n95 ) , .A1( u0_u7_u1_n98 ) );
  NAND2_X1 u0_u7_u1_U51 (.A1( u0_u7_u1_n102 ) , .ZN( u0_u7_u1_n154 ) , .A2( u0_u7_u1_n99 ) );
  NAND2_X1 u0_u7_u1_U52 (.A2( u0_u7_u1_n100 ) , .ZN( u0_u7_u1_n135 ) , .A1( u0_u7_u1_n99 ) );
  AOI21_X1 u0_u7_u1_U53 (.A( u0_u7_u1_n152 ) , .B2( u0_u7_u1_n153 ) , .B1( u0_u7_u1_n154 ) , .ZN( u0_u7_u1_n158 ) );
  INV_X1 u0_u7_u1_U54 (.A( u0_u7_u1_n160 ) , .ZN( u0_u7_u1_n175 ) );
  NAND2_X1 u0_u7_u1_U55 (.A1( u0_u7_u1_n100 ) , .ZN( u0_u7_u1_n116 ) , .A2( u0_u7_u1_n95 ) );
  NAND2_X1 u0_u7_u1_U56 (.A1( u0_u7_u1_n102 ) , .ZN( u0_u7_u1_n131 ) , .A2( u0_u7_u1_n95 ) );
  NAND2_X1 u0_u7_u1_U57 (.A2( u0_u7_u1_n104 ) , .ZN( u0_u7_u1_n121 ) , .A1( u0_u7_u1_n98 ) );
  NAND2_X1 u0_u7_u1_U58 (.A1( u0_u7_u1_n103 ) , .ZN( u0_u7_u1_n153 ) , .A2( u0_u7_u1_n98 ) );
  NAND2_X1 u0_u7_u1_U59 (.A2( u0_u7_u1_n104 ) , .A1( u0_u7_u1_n105 ) , .ZN( u0_u7_u1_n133 ) );
  AOI22_X1 u0_u7_u1_U6 (.B2( u0_u7_u1_n113 ) , .A2( u0_u7_u1_n114 ) , .ZN( u0_u7_u1_n125 ) , .A1( u0_u7_u1_n171 ) , .B1( u0_u7_u1_n173 ) );
  NAND2_X1 u0_u7_u1_U60 (.ZN( u0_u7_u1_n150 ) , .A2( u0_u7_u1_n98 ) , .A1( u0_u7_u1_n99 ) );
  NAND2_X1 u0_u7_u1_U61 (.A1( u0_u7_u1_n105 ) , .ZN( u0_u7_u1_n155 ) , .A2( u0_u7_u1_n95 ) );
  OAI21_X1 u0_u7_u1_U62 (.ZN( u0_u7_u1_n109 ) , .B1( u0_u7_u1_n129 ) , .B2( u0_u7_u1_n160 ) , .A( u0_u7_u1_n167 ) );
  NAND2_X1 u0_u7_u1_U63 (.A2( u0_u7_u1_n100 ) , .A1( u0_u7_u1_n103 ) , .ZN( u0_u7_u1_n120 ) );
  NAND2_X1 u0_u7_u1_U64 (.A1( u0_u7_u1_n102 ) , .A2( u0_u7_u1_n104 ) , .ZN( u0_u7_u1_n115 ) );
  NAND2_X1 u0_u7_u1_U65 (.A2( u0_u7_u1_n100 ) , .A1( u0_u7_u1_n104 ) , .ZN( u0_u7_u1_n151 ) );
  NAND2_X1 u0_u7_u1_U66 (.A2( u0_u7_u1_n103 ) , .A1( u0_u7_u1_n105 ) , .ZN( u0_u7_u1_n161 ) );
  INV_X1 u0_u7_u1_U67 (.A( u0_u7_u1_n152 ) , .ZN( u0_u7_u1_n173 ) );
  INV_X1 u0_u7_u1_U68 (.A( u0_u7_u1_n128 ) , .ZN( u0_u7_u1_n172 ) );
  NAND2_X1 u0_u7_u1_U69 (.A2( u0_u7_u1_n102 ) , .A1( u0_u7_u1_n103 ) , .ZN( u0_u7_u1_n123 ) );
  NAND2_X1 u0_u7_u1_U7 (.ZN( u0_u7_u1_n114 ) , .A1( u0_u7_u1_n134 ) , .A2( u0_u7_u1_n156 ) );
  NOR2_X1 u0_u7_u1_U70 (.A2( u0_u7_X_7 ) , .A1( u0_u7_X_8 ) , .ZN( u0_u7_u1_n95 ) );
  NOR2_X1 u0_u7_u1_U71 (.A1( u0_u7_X_12 ) , .A2( u0_u7_X_9 ) , .ZN( u0_u7_u1_n100 ) );
  NOR2_X1 u0_u7_u1_U72 (.A2( u0_u7_X_8 ) , .A1( u0_u7_u1_n177 ) , .ZN( u0_u7_u1_n99 ) );
  NOR2_X1 u0_u7_u1_U73 (.A2( u0_u7_X_12 ) , .ZN( u0_u7_u1_n102 ) , .A1( u0_u7_u1_n176 ) );
  NOR2_X1 u0_u7_u1_U74 (.A2( u0_u7_X_9 ) , .ZN( u0_u7_u1_n105 ) , .A1( u0_u7_u1_n168 ) );
  NAND2_X1 u0_u7_u1_U75 (.A1( u0_u7_X_10 ) , .ZN( u0_u7_u1_n160 ) , .A2( u0_u7_u1_n169 ) );
  NAND2_X1 u0_u7_u1_U76 (.A2( u0_u7_X_10 ) , .A1( u0_u7_X_11 ) , .ZN( u0_u7_u1_n152 ) );
  NAND2_X1 u0_u7_u1_U77 (.A1( u0_u7_X_11 ) , .ZN( u0_u7_u1_n128 ) , .A2( u0_u7_u1_n170 ) );
  AND2_X1 u0_u7_u1_U78 (.A2( u0_u7_X_7 ) , .A1( u0_u7_X_8 ) , .ZN( u0_u7_u1_n104 ) );
  AND2_X1 u0_u7_u1_U79 (.A1( u0_u7_X_8 ) , .ZN( u0_u7_u1_n103 ) , .A2( u0_u7_u1_n177 ) );
  NOR2_X1 u0_u7_u1_U8 (.A1( u0_u7_u1_n112 ) , .A2( u0_u7_u1_n116 ) , .ZN( u0_u7_u1_n118 ) );
  INV_X1 u0_u7_u1_U80 (.A( u0_u7_X_10 ) , .ZN( u0_u7_u1_n170 ) );
  INV_X1 u0_u7_u1_U81 (.A( u0_u7_X_9 ) , .ZN( u0_u7_u1_n176 ) );
  INV_X1 u0_u7_u1_U82 (.A( u0_u7_X_11 ) , .ZN( u0_u7_u1_n169 ) );
  INV_X1 u0_u7_u1_U83 (.A( u0_u7_X_12 ) , .ZN( u0_u7_u1_n168 ) );
  INV_X1 u0_u7_u1_U84 (.A( u0_u7_X_7 ) , .ZN( u0_u7_u1_n177 ) );
  NAND4_X1 u0_u7_u1_U85 (.ZN( u0_out7_28 ) , .A4( u0_u7_u1_n124 ) , .A3( u0_u7_u1_n125 ) , .A2( u0_u7_u1_n126 ) , .A1( u0_u7_u1_n127 ) );
  OAI21_X1 u0_u7_u1_U86 (.ZN( u0_u7_u1_n127 ) , .B2( u0_u7_u1_n139 ) , .B1( u0_u7_u1_n175 ) , .A( u0_u7_u1_n183 ) );
  OAI21_X1 u0_u7_u1_U87 (.ZN( u0_u7_u1_n126 ) , .B2( u0_u7_u1_n140 ) , .A( u0_u7_u1_n146 ) , .B1( u0_u7_u1_n178 ) );
  NAND4_X1 u0_u7_u1_U88 (.ZN( u0_out7_18 ) , .A4( u0_u7_u1_n165 ) , .A3( u0_u7_u1_n166 ) , .A1( u0_u7_u1_n167 ) , .A2( u0_u7_u1_n186 ) );
  AOI22_X1 u0_u7_u1_U89 (.B2( u0_u7_u1_n146 ) , .B1( u0_u7_u1_n147 ) , .A2( u0_u7_u1_n148 ) , .ZN( u0_u7_u1_n166 ) , .A1( u0_u7_u1_n172 ) );
  OAI21_X1 u0_u7_u1_U9 (.ZN( u0_u7_u1_n101 ) , .B1( u0_u7_u1_n141 ) , .A( u0_u7_u1_n146 ) , .B2( u0_u7_u1_n183 ) );
  INV_X1 u0_u7_u1_U90 (.A( u0_u7_u1_n145 ) , .ZN( u0_u7_u1_n186 ) );
  NAND4_X1 u0_u7_u1_U91 (.ZN( u0_out7_2 ) , .A4( u0_u7_u1_n142 ) , .A3( u0_u7_u1_n143 ) , .A2( u0_u7_u1_n144 ) , .A1( u0_u7_u1_n179 ) );
  OAI21_X1 u0_u7_u1_U92 (.B2( u0_u7_u1_n132 ) , .ZN( u0_u7_u1_n144 ) , .A( u0_u7_u1_n146 ) , .B1( u0_u7_u1_n180 ) );
  INV_X1 u0_u7_u1_U93 (.A( u0_u7_u1_n130 ) , .ZN( u0_u7_u1_n179 ) );
  OR4_X1 u0_u7_u1_U94 (.ZN( u0_out7_13 ) , .A4( u0_u7_u1_n108 ) , .A3( u0_u7_u1_n109 ) , .A2( u0_u7_u1_n110 ) , .A1( u0_u7_u1_n111 ) );
  AOI21_X1 u0_u7_u1_U95 (.ZN( u0_u7_u1_n111 ) , .A( u0_u7_u1_n128 ) , .B2( u0_u7_u1_n131 ) , .B1( u0_u7_u1_n135 ) );
  AOI21_X1 u0_u7_u1_U96 (.ZN( u0_u7_u1_n110 ) , .A( u0_u7_u1_n116 ) , .B1( u0_u7_u1_n152 ) , .B2( u0_u7_u1_n160 ) );
  NAND3_X1 u0_u7_u1_U97 (.A3( u0_u7_u1_n149 ) , .A2( u0_u7_u1_n150 ) , .A1( u0_u7_u1_n151 ) , .ZN( u0_u7_u1_n164 ) );
  NAND3_X1 u0_u7_u1_U98 (.A3( u0_u7_u1_n134 ) , .A2( u0_u7_u1_n135 ) , .ZN( u0_u7_u1_n136 ) , .A1( u0_u7_u1_n151 ) );
  NAND3_X1 u0_u7_u1_U99 (.A1( u0_u7_u1_n133 ) , .ZN( u0_u7_u1_n137 ) , .A2( u0_u7_u1_n154 ) , .A3( u0_u7_u1_n181 ) );
  OAI22_X1 u0_u7_u2_U10 (.ZN( u0_u7_u2_n109 ) , .A2( u0_u7_u2_n113 ) , .B2( u0_u7_u2_n133 ) , .B1( u0_u7_u2_n167 ) , .A1( u0_u7_u2_n168 ) );
  NAND3_X1 u0_u7_u2_U100 (.A2( u0_u7_u2_n100 ) , .A1( u0_u7_u2_n104 ) , .A3( u0_u7_u2_n138 ) , .ZN( u0_u7_u2_n98 ) );
  OAI22_X1 u0_u7_u2_U11 (.B1( u0_u7_u2_n151 ) , .A2( u0_u7_u2_n152 ) , .A1( u0_u7_u2_n153 ) , .ZN( u0_u7_u2_n160 ) , .B2( u0_u7_u2_n168 ) );
  NOR3_X1 u0_u7_u2_U12 (.A1( u0_u7_u2_n150 ) , .ZN( u0_u7_u2_n151 ) , .A3( u0_u7_u2_n175 ) , .A2( u0_u7_u2_n188 ) );
  AOI21_X1 u0_u7_u2_U13 (.ZN( u0_u7_u2_n144 ) , .B2( u0_u7_u2_n155 ) , .A( u0_u7_u2_n172 ) , .B1( u0_u7_u2_n185 ) );
  AOI21_X1 u0_u7_u2_U14 (.B2( u0_u7_u2_n143 ) , .ZN( u0_u7_u2_n145 ) , .B1( u0_u7_u2_n152 ) , .A( u0_u7_u2_n171 ) );
  AOI21_X1 u0_u7_u2_U15 (.B2( u0_u7_u2_n120 ) , .B1( u0_u7_u2_n121 ) , .ZN( u0_u7_u2_n126 ) , .A( u0_u7_u2_n167 ) );
  INV_X1 u0_u7_u2_U16 (.A( u0_u7_u2_n156 ) , .ZN( u0_u7_u2_n171 ) );
  INV_X1 u0_u7_u2_U17 (.A( u0_u7_u2_n120 ) , .ZN( u0_u7_u2_n188 ) );
  NAND2_X1 u0_u7_u2_U18 (.A2( u0_u7_u2_n122 ) , .ZN( u0_u7_u2_n150 ) , .A1( u0_u7_u2_n152 ) );
  INV_X1 u0_u7_u2_U19 (.A( u0_u7_u2_n153 ) , .ZN( u0_u7_u2_n170 ) );
  INV_X1 u0_u7_u2_U20 (.A( u0_u7_u2_n137 ) , .ZN( u0_u7_u2_n173 ) );
  NAND2_X1 u0_u7_u2_U21 (.A1( u0_u7_u2_n132 ) , .A2( u0_u7_u2_n139 ) , .ZN( u0_u7_u2_n157 ) );
  INV_X1 u0_u7_u2_U22 (.A( u0_u7_u2_n113 ) , .ZN( u0_u7_u2_n178 ) );
  INV_X1 u0_u7_u2_U23 (.A( u0_u7_u2_n139 ) , .ZN( u0_u7_u2_n175 ) );
  INV_X1 u0_u7_u2_U24 (.A( u0_u7_u2_n155 ) , .ZN( u0_u7_u2_n181 ) );
  INV_X1 u0_u7_u2_U25 (.A( u0_u7_u2_n119 ) , .ZN( u0_u7_u2_n177 ) );
  INV_X1 u0_u7_u2_U26 (.A( u0_u7_u2_n116 ) , .ZN( u0_u7_u2_n180 ) );
  INV_X1 u0_u7_u2_U27 (.A( u0_u7_u2_n131 ) , .ZN( u0_u7_u2_n179 ) );
  INV_X1 u0_u7_u2_U28 (.A( u0_u7_u2_n154 ) , .ZN( u0_u7_u2_n176 ) );
  NAND2_X1 u0_u7_u2_U29 (.A2( u0_u7_u2_n116 ) , .A1( u0_u7_u2_n117 ) , .ZN( u0_u7_u2_n118 ) );
  NOR2_X1 u0_u7_u2_U3 (.ZN( u0_u7_u2_n121 ) , .A2( u0_u7_u2_n177 ) , .A1( u0_u7_u2_n180 ) );
  INV_X1 u0_u7_u2_U30 (.A( u0_u7_u2_n132 ) , .ZN( u0_u7_u2_n182 ) );
  INV_X1 u0_u7_u2_U31 (.A( u0_u7_u2_n158 ) , .ZN( u0_u7_u2_n183 ) );
  OAI21_X1 u0_u7_u2_U32 (.A( u0_u7_u2_n156 ) , .B1( u0_u7_u2_n157 ) , .ZN( u0_u7_u2_n158 ) , .B2( u0_u7_u2_n179 ) );
  NOR2_X1 u0_u7_u2_U33 (.ZN( u0_u7_u2_n156 ) , .A1( u0_u7_u2_n166 ) , .A2( u0_u7_u2_n169 ) );
  NOR2_X1 u0_u7_u2_U34 (.A2( u0_u7_u2_n114 ) , .ZN( u0_u7_u2_n137 ) , .A1( u0_u7_u2_n140 ) );
  NOR2_X1 u0_u7_u2_U35 (.A2( u0_u7_u2_n138 ) , .ZN( u0_u7_u2_n153 ) , .A1( u0_u7_u2_n156 ) );
  AOI211_X1 u0_u7_u2_U36 (.ZN( u0_u7_u2_n130 ) , .C1( u0_u7_u2_n138 ) , .C2( u0_u7_u2_n179 ) , .B( u0_u7_u2_n96 ) , .A( u0_u7_u2_n97 ) );
  OAI22_X1 u0_u7_u2_U37 (.B1( u0_u7_u2_n133 ) , .A2( u0_u7_u2_n137 ) , .A1( u0_u7_u2_n152 ) , .B2( u0_u7_u2_n168 ) , .ZN( u0_u7_u2_n97 ) );
  OAI221_X1 u0_u7_u2_U38 (.B1( u0_u7_u2_n113 ) , .C1( u0_u7_u2_n132 ) , .A( u0_u7_u2_n149 ) , .B2( u0_u7_u2_n171 ) , .C2( u0_u7_u2_n172 ) , .ZN( u0_u7_u2_n96 ) );
  OAI221_X1 u0_u7_u2_U39 (.A( u0_u7_u2_n115 ) , .C2( u0_u7_u2_n123 ) , .B2( u0_u7_u2_n143 ) , .B1( u0_u7_u2_n153 ) , .ZN( u0_u7_u2_n163 ) , .C1( u0_u7_u2_n168 ) );
  INV_X1 u0_u7_u2_U4 (.A( u0_u7_u2_n134 ) , .ZN( u0_u7_u2_n185 ) );
  OAI21_X1 u0_u7_u2_U40 (.A( u0_u7_u2_n114 ) , .ZN( u0_u7_u2_n115 ) , .B1( u0_u7_u2_n176 ) , .B2( u0_u7_u2_n178 ) );
  OAI221_X1 u0_u7_u2_U41 (.A( u0_u7_u2_n135 ) , .B2( u0_u7_u2_n136 ) , .B1( u0_u7_u2_n137 ) , .ZN( u0_u7_u2_n162 ) , .C2( u0_u7_u2_n167 ) , .C1( u0_u7_u2_n185 ) );
  AND3_X1 u0_u7_u2_U42 (.A3( u0_u7_u2_n131 ) , .A2( u0_u7_u2_n132 ) , .A1( u0_u7_u2_n133 ) , .ZN( u0_u7_u2_n136 ) );
  AOI22_X1 u0_u7_u2_U43 (.ZN( u0_u7_u2_n135 ) , .B1( u0_u7_u2_n140 ) , .A1( u0_u7_u2_n156 ) , .B2( u0_u7_u2_n180 ) , .A2( u0_u7_u2_n188 ) );
  AOI21_X1 u0_u7_u2_U44 (.ZN( u0_u7_u2_n149 ) , .B1( u0_u7_u2_n173 ) , .B2( u0_u7_u2_n188 ) , .A( u0_u7_u2_n95 ) );
  AND3_X1 u0_u7_u2_U45 (.A2( u0_u7_u2_n100 ) , .A1( u0_u7_u2_n104 ) , .A3( u0_u7_u2_n156 ) , .ZN( u0_u7_u2_n95 ) );
  OAI21_X1 u0_u7_u2_U46 (.A( u0_u7_u2_n101 ) , .B2( u0_u7_u2_n121 ) , .B1( u0_u7_u2_n153 ) , .ZN( u0_u7_u2_n164 ) );
  NAND2_X1 u0_u7_u2_U47 (.A2( u0_u7_u2_n100 ) , .A1( u0_u7_u2_n107 ) , .ZN( u0_u7_u2_n155 ) );
  NAND2_X1 u0_u7_u2_U48 (.A2( u0_u7_u2_n105 ) , .A1( u0_u7_u2_n108 ) , .ZN( u0_u7_u2_n143 ) );
  NAND2_X1 u0_u7_u2_U49 (.A1( u0_u7_u2_n104 ) , .A2( u0_u7_u2_n106 ) , .ZN( u0_u7_u2_n152 ) );
  INV_X1 u0_u7_u2_U5 (.A( u0_u7_u2_n150 ) , .ZN( u0_u7_u2_n184 ) );
  NAND2_X1 u0_u7_u2_U50 (.A1( u0_u7_u2_n100 ) , .A2( u0_u7_u2_n105 ) , .ZN( u0_u7_u2_n132 ) );
  INV_X1 u0_u7_u2_U51 (.A( u0_u7_u2_n140 ) , .ZN( u0_u7_u2_n168 ) );
  INV_X1 u0_u7_u2_U52 (.A( u0_u7_u2_n138 ) , .ZN( u0_u7_u2_n167 ) );
  OAI21_X1 u0_u7_u2_U53 (.A( u0_u7_u2_n141 ) , .B2( u0_u7_u2_n142 ) , .ZN( u0_u7_u2_n146 ) , .B1( u0_u7_u2_n153 ) );
  OAI21_X1 u0_u7_u2_U54 (.A( u0_u7_u2_n140 ) , .ZN( u0_u7_u2_n141 ) , .B1( u0_u7_u2_n176 ) , .B2( u0_u7_u2_n177 ) );
  NOR3_X1 u0_u7_u2_U55 (.ZN( u0_u7_u2_n142 ) , .A3( u0_u7_u2_n175 ) , .A2( u0_u7_u2_n178 ) , .A1( u0_u7_u2_n181 ) );
  INV_X1 u0_u7_u2_U56 (.ZN( u0_u7_u2_n187 ) , .A( u0_u7_u2_n99 ) );
  OAI21_X1 u0_u7_u2_U57 (.B1( u0_u7_u2_n137 ) , .B2( u0_u7_u2_n143 ) , .A( u0_u7_u2_n98 ) , .ZN( u0_u7_u2_n99 ) );
  NAND2_X1 u0_u7_u2_U58 (.A1( u0_u7_u2_n102 ) , .A2( u0_u7_u2_n106 ) , .ZN( u0_u7_u2_n113 ) );
  NAND2_X1 u0_u7_u2_U59 (.A1( u0_u7_u2_n106 ) , .A2( u0_u7_u2_n107 ) , .ZN( u0_u7_u2_n131 ) );
  NOR4_X1 u0_u7_u2_U6 (.A4( u0_u7_u2_n124 ) , .A3( u0_u7_u2_n125 ) , .A2( u0_u7_u2_n126 ) , .A1( u0_u7_u2_n127 ) , .ZN( u0_u7_u2_n128 ) );
  NAND2_X1 u0_u7_u2_U60 (.A1( u0_u7_u2_n103 ) , .A2( u0_u7_u2_n107 ) , .ZN( u0_u7_u2_n139 ) );
  NAND2_X1 u0_u7_u2_U61 (.A1( u0_u7_u2_n103 ) , .A2( u0_u7_u2_n105 ) , .ZN( u0_u7_u2_n133 ) );
  NAND2_X1 u0_u7_u2_U62 (.A1( u0_u7_u2_n102 ) , .A2( u0_u7_u2_n103 ) , .ZN( u0_u7_u2_n154 ) );
  NAND2_X1 u0_u7_u2_U63 (.A2( u0_u7_u2_n103 ) , .A1( u0_u7_u2_n104 ) , .ZN( u0_u7_u2_n119 ) );
  NAND2_X1 u0_u7_u2_U64 (.A2( u0_u7_u2_n107 ) , .A1( u0_u7_u2_n108 ) , .ZN( u0_u7_u2_n123 ) );
  NAND2_X1 u0_u7_u2_U65 (.A1( u0_u7_u2_n104 ) , .A2( u0_u7_u2_n108 ) , .ZN( u0_u7_u2_n122 ) );
  INV_X1 u0_u7_u2_U66 (.A( u0_u7_u2_n114 ) , .ZN( u0_u7_u2_n172 ) );
  NAND2_X1 u0_u7_u2_U67 (.A2( u0_u7_u2_n100 ) , .A1( u0_u7_u2_n102 ) , .ZN( u0_u7_u2_n116 ) );
  NAND2_X1 u0_u7_u2_U68 (.A1( u0_u7_u2_n102 ) , .A2( u0_u7_u2_n108 ) , .ZN( u0_u7_u2_n120 ) );
  NAND2_X1 u0_u7_u2_U69 (.A2( u0_u7_u2_n105 ) , .A1( u0_u7_u2_n106 ) , .ZN( u0_u7_u2_n117 ) );
  AOI21_X1 u0_u7_u2_U7 (.B2( u0_u7_u2_n119 ) , .ZN( u0_u7_u2_n127 ) , .A( u0_u7_u2_n137 ) , .B1( u0_u7_u2_n155 ) );
  NOR2_X1 u0_u7_u2_U70 (.A2( u0_u7_X_16 ) , .ZN( u0_u7_u2_n140 ) , .A1( u0_u7_u2_n166 ) );
  NOR2_X1 u0_u7_u2_U71 (.A2( u0_u7_X_13 ) , .A1( u0_u7_X_14 ) , .ZN( u0_u7_u2_n100 ) );
  NOR2_X1 u0_u7_u2_U72 (.A2( u0_u7_X_16 ) , .A1( u0_u7_X_17 ) , .ZN( u0_u7_u2_n138 ) );
  NOR2_X1 u0_u7_u2_U73 (.A2( u0_u7_X_15 ) , .A1( u0_u7_X_18 ) , .ZN( u0_u7_u2_n104 ) );
  NOR2_X1 u0_u7_u2_U74 (.A2( u0_u7_X_14 ) , .ZN( u0_u7_u2_n103 ) , .A1( u0_u7_u2_n174 ) );
  NOR2_X1 u0_u7_u2_U75 (.A2( u0_u7_X_15 ) , .ZN( u0_u7_u2_n102 ) , .A1( u0_u7_u2_n165 ) );
  NOR2_X1 u0_u7_u2_U76 (.A2( u0_u7_X_17 ) , .ZN( u0_u7_u2_n114 ) , .A1( u0_u7_u2_n169 ) );
  AND2_X1 u0_u7_u2_U77 (.A1( u0_u7_X_15 ) , .ZN( u0_u7_u2_n105 ) , .A2( u0_u7_u2_n165 ) );
  AND2_X1 u0_u7_u2_U78 (.A2( u0_u7_X_15 ) , .A1( u0_u7_X_18 ) , .ZN( u0_u7_u2_n107 ) );
  AND2_X1 u0_u7_u2_U79 (.A1( u0_u7_X_14 ) , .ZN( u0_u7_u2_n106 ) , .A2( u0_u7_u2_n174 ) );
  AOI21_X1 u0_u7_u2_U8 (.ZN( u0_u7_u2_n124 ) , .B1( u0_u7_u2_n131 ) , .B2( u0_u7_u2_n143 ) , .A( u0_u7_u2_n172 ) );
  AND2_X1 u0_u7_u2_U80 (.A1( u0_u7_X_13 ) , .A2( u0_u7_X_14 ) , .ZN( u0_u7_u2_n108 ) );
  INV_X1 u0_u7_u2_U81 (.A( u0_u7_X_16 ) , .ZN( u0_u7_u2_n169 ) );
  INV_X1 u0_u7_u2_U82 (.A( u0_u7_X_17 ) , .ZN( u0_u7_u2_n166 ) );
  INV_X1 u0_u7_u2_U83 (.A( u0_u7_X_13 ) , .ZN( u0_u7_u2_n174 ) );
  INV_X1 u0_u7_u2_U84 (.A( u0_u7_X_18 ) , .ZN( u0_u7_u2_n165 ) );
  NAND4_X1 u0_u7_u2_U85 (.ZN( u0_out7_30 ) , .A4( u0_u7_u2_n147 ) , .A3( u0_u7_u2_n148 ) , .A2( u0_u7_u2_n149 ) , .A1( u0_u7_u2_n187 ) );
  NOR3_X1 u0_u7_u2_U86 (.A3( u0_u7_u2_n144 ) , .A2( u0_u7_u2_n145 ) , .A1( u0_u7_u2_n146 ) , .ZN( u0_u7_u2_n147 ) );
  AOI21_X1 u0_u7_u2_U87 (.B2( u0_u7_u2_n138 ) , .ZN( u0_u7_u2_n148 ) , .A( u0_u7_u2_n162 ) , .B1( u0_u7_u2_n182 ) );
  NAND4_X1 u0_u7_u2_U88 (.ZN( u0_out7_24 ) , .A4( u0_u7_u2_n111 ) , .A3( u0_u7_u2_n112 ) , .A1( u0_u7_u2_n130 ) , .A2( u0_u7_u2_n187 ) );
  AOI221_X1 u0_u7_u2_U89 (.A( u0_u7_u2_n109 ) , .B1( u0_u7_u2_n110 ) , .ZN( u0_u7_u2_n111 ) , .C1( u0_u7_u2_n134 ) , .C2( u0_u7_u2_n170 ) , .B2( u0_u7_u2_n173 ) );
  AOI21_X1 u0_u7_u2_U9 (.B2( u0_u7_u2_n123 ) , .ZN( u0_u7_u2_n125 ) , .A( u0_u7_u2_n171 ) , .B1( u0_u7_u2_n184 ) );
  AOI21_X1 u0_u7_u2_U90 (.ZN( u0_u7_u2_n112 ) , .B2( u0_u7_u2_n156 ) , .A( u0_u7_u2_n164 ) , .B1( u0_u7_u2_n181 ) );
  NAND4_X1 u0_u7_u2_U91 (.ZN( u0_out7_16 ) , .A4( u0_u7_u2_n128 ) , .A3( u0_u7_u2_n129 ) , .A1( u0_u7_u2_n130 ) , .A2( u0_u7_u2_n186 ) );
  AOI22_X1 u0_u7_u2_U92 (.A2( u0_u7_u2_n118 ) , .ZN( u0_u7_u2_n129 ) , .A1( u0_u7_u2_n140 ) , .B1( u0_u7_u2_n157 ) , .B2( u0_u7_u2_n170 ) );
  INV_X1 u0_u7_u2_U93 (.A( u0_u7_u2_n163 ) , .ZN( u0_u7_u2_n186 ) );
  OR4_X1 u0_u7_u2_U94 (.ZN( u0_out7_6 ) , .A4( u0_u7_u2_n161 ) , .A3( u0_u7_u2_n162 ) , .A2( u0_u7_u2_n163 ) , .A1( u0_u7_u2_n164 ) );
  OR3_X1 u0_u7_u2_U95 (.A2( u0_u7_u2_n159 ) , .A1( u0_u7_u2_n160 ) , .ZN( u0_u7_u2_n161 ) , .A3( u0_u7_u2_n183 ) );
  AOI21_X1 u0_u7_u2_U96 (.B2( u0_u7_u2_n154 ) , .B1( u0_u7_u2_n155 ) , .ZN( u0_u7_u2_n159 ) , .A( u0_u7_u2_n167 ) );
  NAND3_X1 u0_u7_u2_U97 (.A2( u0_u7_u2_n117 ) , .A1( u0_u7_u2_n122 ) , .A3( u0_u7_u2_n123 ) , .ZN( u0_u7_u2_n134 ) );
  NAND3_X1 u0_u7_u2_U98 (.ZN( u0_u7_u2_n110 ) , .A2( u0_u7_u2_n131 ) , .A3( u0_u7_u2_n139 ) , .A1( u0_u7_u2_n154 ) );
  NAND3_X1 u0_u7_u2_U99 (.A2( u0_u7_u2_n100 ) , .ZN( u0_u7_u2_n101 ) , .A1( u0_u7_u2_n104 ) , .A3( u0_u7_u2_n114 ) );
  OAI22_X1 u0_u7_u3_U10 (.B1( u0_u7_u3_n113 ) , .A2( u0_u7_u3_n135 ) , .A1( u0_u7_u3_n150 ) , .B2( u0_u7_u3_n164 ) , .ZN( u0_u7_u3_n98 ) );
  OAI211_X1 u0_u7_u3_U11 (.B( u0_u7_u3_n106 ) , .ZN( u0_u7_u3_n119 ) , .C2( u0_u7_u3_n128 ) , .C1( u0_u7_u3_n167 ) , .A( u0_u7_u3_n181 ) );
  AOI221_X1 u0_u7_u3_U12 (.C1( u0_u7_u3_n105 ) , .ZN( u0_u7_u3_n106 ) , .A( u0_u7_u3_n131 ) , .B2( u0_u7_u3_n132 ) , .C2( u0_u7_u3_n133 ) , .B1( u0_u7_u3_n169 ) );
  INV_X1 u0_u7_u3_U13 (.ZN( u0_u7_u3_n181 ) , .A( u0_u7_u3_n98 ) );
  NAND2_X1 u0_u7_u3_U14 (.ZN( u0_u7_u3_n105 ) , .A2( u0_u7_u3_n130 ) , .A1( u0_u7_u3_n155 ) );
  AOI22_X1 u0_u7_u3_U15 (.B1( u0_u7_u3_n115 ) , .A2( u0_u7_u3_n116 ) , .ZN( u0_u7_u3_n123 ) , .B2( u0_u7_u3_n133 ) , .A1( u0_u7_u3_n169 ) );
  NAND2_X1 u0_u7_u3_U16 (.ZN( u0_u7_u3_n116 ) , .A2( u0_u7_u3_n151 ) , .A1( u0_u7_u3_n182 ) );
  NOR2_X1 u0_u7_u3_U17 (.ZN( u0_u7_u3_n126 ) , .A2( u0_u7_u3_n150 ) , .A1( u0_u7_u3_n164 ) );
  AOI21_X1 u0_u7_u3_U18 (.ZN( u0_u7_u3_n112 ) , .B2( u0_u7_u3_n146 ) , .B1( u0_u7_u3_n155 ) , .A( u0_u7_u3_n167 ) );
  NAND2_X1 u0_u7_u3_U19 (.A1( u0_u7_u3_n135 ) , .ZN( u0_u7_u3_n142 ) , .A2( u0_u7_u3_n164 ) );
  NAND2_X1 u0_u7_u3_U20 (.ZN( u0_u7_u3_n132 ) , .A2( u0_u7_u3_n152 ) , .A1( u0_u7_u3_n156 ) );
  AND2_X1 u0_u7_u3_U21 (.A2( u0_u7_u3_n113 ) , .A1( u0_u7_u3_n114 ) , .ZN( u0_u7_u3_n151 ) );
  INV_X1 u0_u7_u3_U22 (.A( u0_u7_u3_n133 ) , .ZN( u0_u7_u3_n165 ) );
  INV_X1 u0_u7_u3_U23 (.A( u0_u7_u3_n135 ) , .ZN( u0_u7_u3_n170 ) );
  NAND2_X1 u0_u7_u3_U24 (.A1( u0_u7_u3_n107 ) , .A2( u0_u7_u3_n108 ) , .ZN( u0_u7_u3_n140 ) );
  NAND2_X1 u0_u7_u3_U25 (.ZN( u0_u7_u3_n117 ) , .A1( u0_u7_u3_n124 ) , .A2( u0_u7_u3_n148 ) );
  NAND2_X1 u0_u7_u3_U26 (.ZN( u0_u7_u3_n143 ) , .A1( u0_u7_u3_n165 ) , .A2( u0_u7_u3_n167 ) );
  INV_X1 u0_u7_u3_U27 (.A( u0_u7_u3_n130 ) , .ZN( u0_u7_u3_n177 ) );
  INV_X1 u0_u7_u3_U28 (.A( u0_u7_u3_n128 ) , .ZN( u0_u7_u3_n176 ) );
  INV_X1 u0_u7_u3_U29 (.A( u0_u7_u3_n155 ) , .ZN( u0_u7_u3_n174 ) );
  INV_X1 u0_u7_u3_U3 (.A( u0_u7_u3_n129 ) , .ZN( u0_u7_u3_n183 ) );
  INV_X1 u0_u7_u3_U30 (.A( u0_u7_u3_n139 ) , .ZN( u0_u7_u3_n185 ) );
  NOR2_X1 u0_u7_u3_U31 (.ZN( u0_u7_u3_n135 ) , .A2( u0_u7_u3_n141 ) , .A1( u0_u7_u3_n169 ) );
  OAI222_X1 u0_u7_u3_U32 (.C2( u0_u7_u3_n107 ) , .A2( u0_u7_u3_n108 ) , .B1( u0_u7_u3_n135 ) , .ZN( u0_u7_u3_n138 ) , .B2( u0_u7_u3_n146 ) , .C1( u0_u7_u3_n154 ) , .A1( u0_u7_u3_n164 ) );
  NOR4_X1 u0_u7_u3_U33 (.A4( u0_u7_u3_n157 ) , .A3( u0_u7_u3_n158 ) , .A2( u0_u7_u3_n159 ) , .A1( u0_u7_u3_n160 ) , .ZN( u0_u7_u3_n161 ) );
  AOI21_X1 u0_u7_u3_U34 (.B2( u0_u7_u3_n152 ) , .B1( u0_u7_u3_n153 ) , .ZN( u0_u7_u3_n158 ) , .A( u0_u7_u3_n164 ) );
  AOI21_X1 u0_u7_u3_U35 (.A( u0_u7_u3_n154 ) , .B2( u0_u7_u3_n155 ) , .B1( u0_u7_u3_n156 ) , .ZN( u0_u7_u3_n157 ) );
  AOI21_X1 u0_u7_u3_U36 (.A( u0_u7_u3_n149 ) , .B2( u0_u7_u3_n150 ) , .B1( u0_u7_u3_n151 ) , .ZN( u0_u7_u3_n159 ) );
  AOI211_X1 u0_u7_u3_U37 (.ZN( u0_u7_u3_n109 ) , .A( u0_u7_u3_n119 ) , .C2( u0_u7_u3_n129 ) , .B( u0_u7_u3_n138 ) , .C1( u0_u7_u3_n141 ) );
  AOI211_X1 u0_u7_u3_U38 (.B( u0_u7_u3_n119 ) , .A( u0_u7_u3_n120 ) , .C2( u0_u7_u3_n121 ) , .ZN( u0_u7_u3_n122 ) , .C1( u0_u7_u3_n179 ) );
  INV_X1 u0_u7_u3_U39 (.A( u0_u7_u3_n156 ) , .ZN( u0_u7_u3_n179 ) );
  INV_X1 u0_u7_u3_U4 (.A( u0_u7_u3_n140 ) , .ZN( u0_u7_u3_n182 ) );
  OAI22_X1 u0_u7_u3_U40 (.B1( u0_u7_u3_n118 ) , .ZN( u0_u7_u3_n120 ) , .A1( u0_u7_u3_n135 ) , .B2( u0_u7_u3_n154 ) , .A2( u0_u7_u3_n178 ) );
  AND3_X1 u0_u7_u3_U41 (.ZN( u0_u7_u3_n118 ) , .A2( u0_u7_u3_n124 ) , .A1( u0_u7_u3_n144 ) , .A3( u0_u7_u3_n152 ) );
  INV_X1 u0_u7_u3_U42 (.A( u0_u7_u3_n121 ) , .ZN( u0_u7_u3_n164 ) );
  NAND2_X1 u0_u7_u3_U43 (.ZN( u0_u7_u3_n133 ) , .A1( u0_u7_u3_n154 ) , .A2( u0_u7_u3_n164 ) );
  OAI211_X1 u0_u7_u3_U44 (.B( u0_u7_u3_n127 ) , .ZN( u0_u7_u3_n139 ) , .C1( u0_u7_u3_n150 ) , .C2( u0_u7_u3_n154 ) , .A( u0_u7_u3_n184 ) );
  INV_X1 u0_u7_u3_U45 (.A( u0_u7_u3_n125 ) , .ZN( u0_u7_u3_n184 ) );
  AOI221_X1 u0_u7_u3_U46 (.A( u0_u7_u3_n126 ) , .ZN( u0_u7_u3_n127 ) , .C2( u0_u7_u3_n132 ) , .C1( u0_u7_u3_n169 ) , .B2( u0_u7_u3_n170 ) , .B1( u0_u7_u3_n174 ) );
  OAI22_X1 u0_u7_u3_U47 (.A1( u0_u7_u3_n124 ) , .ZN( u0_u7_u3_n125 ) , .B2( u0_u7_u3_n145 ) , .A2( u0_u7_u3_n165 ) , .B1( u0_u7_u3_n167 ) );
  NOR2_X1 u0_u7_u3_U48 (.A1( u0_u7_u3_n113 ) , .ZN( u0_u7_u3_n131 ) , .A2( u0_u7_u3_n154 ) );
  NAND2_X1 u0_u7_u3_U49 (.A1( u0_u7_u3_n103 ) , .ZN( u0_u7_u3_n150 ) , .A2( u0_u7_u3_n99 ) );
  INV_X1 u0_u7_u3_U5 (.A( u0_u7_u3_n117 ) , .ZN( u0_u7_u3_n178 ) );
  NAND2_X1 u0_u7_u3_U50 (.A2( u0_u7_u3_n102 ) , .ZN( u0_u7_u3_n155 ) , .A1( u0_u7_u3_n97 ) );
  INV_X1 u0_u7_u3_U51 (.A( u0_u7_u3_n141 ) , .ZN( u0_u7_u3_n167 ) );
  AOI21_X1 u0_u7_u3_U52 (.B2( u0_u7_u3_n114 ) , .B1( u0_u7_u3_n146 ) , .A( u0_u7_u3_n154 ) , .ZN( u0_u7_u3_n94 ) );
  AOI21_X1 u0_u7_u3_U53 (.ZN( u0_u7_u3_n110 ) , .B2( u0_u7_u3_n142 ) , .B1( u0_u7_u3_n186 ) , .A( u0_u7_u3_n95 ) );
  INV_X1 u0_u7_u3_U54 (.A( u0_u7_u3_n145 ) , .ZN( u0_u7_u3_n186 ) );
  AOI21_X1 u0_u7_u3_U55 (.B1( u0_u7_u3_n124 ) , .A( u0_u7_u3_n149 ) , .B2( u0_u7_u3_n155 ) , .ZN( u0_u7_u3_n95 ) );
  INV_X1 u0_u7_u3_U56 (.A( u0_u7_u3_n149 ) , .ZN( u0_u7_u3_n169 ) );
  NAND2_X1 u0_u7_u3_U57 (.ZN( u0_u7_u3_n124 ) , .A1( u0_u7_u3_n96 ) , .A2( u0_u7_u3_n97 ) );
  NAND2_X1 u0_u7_u3_U58 (.A2( u0_u7_u3_n100 ) , .ZN( u0_u7_u3_n146 ) , .A1( u0_u7_u3_n96 ) );
  NAND2_X1 u0_u7_u3_U59 (.A1( u0_u7_u3_n101 ) , .ZN( u0_u7_u3_n145 ) , .A2( u0_u7_u3_n99 ) );
  AOI221_X1 u0_u7_u3_U6 (.A( u0_u7_u3_n131 ) , .C2( u0_u7_u3_n132 ) , .C1( u0_u7_u3_n133 ) , .ZN( u0_u7_u3_n134 ) , .B1( u0_u7_u3_n143 ) , .B2( u0_u7_u3_n177 ) );
  NAND2_X1 u0_u7_u3_U60 (.A1( u0_u7_u3_n100 ) , .ZN( u0_u7_u3_n156 ) , .A2( u0_u7_u3_n99 ) );
  NAND2_X1 u0_u7_u3_U61 (.A2( u0_u7_u3_n101 ) , .A1( u0_u7_u3_n104 ) , .ZN( u0_u7_u3_n148 ) );
  NAND2_X1 u0_u7_u3_U62 (.A1( u0_u7_u3_n100 ) , .A2( u0_u7_u3_n102 ) , .ZN( u0_u7_u3_n128 ) );
  NAND2_X1 u0_u7_u3_U63 (.A2( u0_u7_u3_n101 ) , .A1( u0_u7_u3_n102 ) , .ZN( u0_u7_u3_n152 ) );
  NAND2_X1 u0_u7_u3_U64 (.A2( u0_u7_u3_n101 ) , .ZN( u0_u7_u3_n114 ) , .A1( u0_u7_u3_n96 ) );
  NAND2_X1 u0_u7_u3_U65 (.ZN( u0_u7_u3_n107 ) , .A1( u0_u7_u3_n97 ) , .A2( u0_u7_u3_n99 ) );
  NAND2_X1 u0_u7_u3_U66 (.A2( u0_u7_u3_n100 ) , .A1( u0_u7_u3_n104 ) , .ZN( u0_u7_u3_n113 ) );
  NAND2_X1 u0_u7_u3_U67 (.A1( u0_u7_u3_n104 ) , .ZN( u0_u7_u3_n153 ) , .A2( u0_u7_u3_n97 ) );
  NAND2_X1 u0_u7_u3_U68 (.A2( u0_u7_u3_n103 ) , .A1( u0_u7_u3_n104 ) , .ZN( u0_u7_u3_n130 ) );
  NAND2_X1 u0_u7_u3_U69 (.A2( u0_u7_u3_n103 ) , .ZN( u0_u7_u3_n144 ) , .A1( u0_u7_u3_n96 ) );
  OAI22_X1 u0_u7_u3_U7 (.B2( u0_u7_u3_n147 ) , .A2( u0_u7_u3_n148 ) , .ZN( u0_u7_u3_n160 ) , .B1( u0_u7_u3_n165 ) , .A1( u0_u7_u3_n168 ) );
  NAND2_X1 u0_u7_u3_U70 (.A1( u0_u7_u3_n102 ) , .A2( u0_u7_u3_n103 ) , .ZN( u0_u7_u3_n108 ) );
  NOR2_X1 u0_u7_u3_U71 (.A2( u0_u7_X_19 ) , .A1( u0_u7_X_20 ) , .ZN( u0_u7_u3_n99 ) );
  NOR2_X1 u0_u7_u3_U72 (.A2( u0_u7_X_21 ) , .A1( u0_u7_X_24 ) , .ZN( u0_u7_u3_n103 ) );
  NOR2_X1 u0_u7_u3_U73 (.A2( u0_u7_X_24 ) , .A1( u0_u7_u3_n171 ) , .ZN( u0_u7_u3_n97 ) );
  NOR2_X1 u0_u7_u3_U74 (.A2( u0_u7_X_23 ) , .ZN( u0_u7_u3_n141 ) , .A1( u0_u7_u3_n166 ) );
  NOR2_X1 u0_u7_u3_U75 (.A2( u0_u7_X_19 ) , .A1( u0_u7_u3_n172 ) , .ZN( u0_u7_u3_n96 ) );
  NAND2_X1 u0_u7_u3_U76 (.A1( u0_u7_X_22 ) , .A2( u0_u7_X_23 ) , .ZN( u0_u7_u3_n154 ) );
  NAND2_X1 u0_u7_u3_U77 (.A1( u0_u7_X_23 ) , .ZN( u0_u7_u3_n149 ) , .A2( u0_u7_u3_n166 ) );
  NOR2_X1 u0_u7_u3_U78 (.A2( u0_u7_X_22 ) , .A1( u0_u7_X_23 ) , .ZN( u0_u7_u3_n121 ) );
  AND2_X1 u0_u7_u3_U79 (.A1( u0_u7_X_24 ) , .ZN( u0_u7_u3_n101 ) , .A2( u0_u7_u3_n171 ) );
  AND3_X1 u0_u7_u3_U8 (.A3( u0_u7_u3_n144 ) , .A2( u0_u7_u3_n145 ) , .A1( u0_u7_u3_n146 ) , .ZN( u0_u7_u3_n147 ) );
  AND2_X1 u0_u7_u3_U80 (.A1( u0_u7_X_19 ) , .ZN( u0_u7_u3_n102 ) , .A2( u0_u7_u3_n172 ) );
  AND2_X1 u0_u7_u3_U81 (.A1( u0_u7_X_21 ) , .A2( u0_u7_X_24 ) , .ZN( u0_u7_u3_n100 ) );
  AND2_X1 u0_u7_u3_U82 (.A2( u0_u7_X_19 ) , .A1( u0_u7_X_20 ) , .ZN( u0_u7_u3_n104 ) );
  INV_X1 u0_u7_u3_U83 (.A( u0_u7_X_22 ) , .ZN( u0_u7_u3_n166 ) );
  INV_X1 u0_u7_u3_U84 (.A( u0_u7_X_21 ) , .ZN( u0_u7_u3_n171 ) );
  INV_X1 u0_u7_u3_U85 (.A( u0_u7_X_20 ) , .ZN( u0_u7_u3_n172 ) );
  OR4_X1 u0_u7_u3_U86 (.ZN( u0_out7_10 ) , .A4( u0_u7_u3_n136 ) , .A3( u0_u7_u3_n137 ) , .A1( u0_u7_u3_n138 ) , .A2( u0_u7_u3_n139 ) );
  OAI222_X1 u0_u7_u3_U87 (.C1( u0_u7_u3_n128 ) , .ZN( u0_u7_u3_n137 ) , .B1( u0_u7_u3_n148 ) , .A2( u0_u7_u3_n150 ) , .B2( u0_u7_u3_n154 ) , .C2( u0_u7_u3_n164 ) , .A1( u0_u7_u3_n167 ) );
  OAI221_X1 u0_u7_u3_U88 (.A( u0_u7_u3_n134 ) , .B2( u0_u7_u3_n135 ) , .ZN( u0_u7_u3_n136 ) , .C1( u0_u7_u3_n149 ) , .B1( u0_u7_u3_n151 ) , .C2( u0_u7_u3_n183 ) );
  NAND4_X1 u0_u7_u3_U89 (.ZN( u0_out7_26 ) , .A4( u0_u7_u3_n109 ) , .A3( u0_u7_u3_n110 ) , .A2( u0_u7_u3_n111 ) , .A1( u0_u7_u3_n173 ) );
  INV_X1 u0_u7_u3_U9 (.A( u0_u7_u3_n143 ) , .ZN( u0_u7_u3_n168 ) );
  INV_X1 u0_u7_u3_U90 (.ZN( u0_u7_u3_n173 ) , .A( u0_u7_u3_n94 ) );
  OAI21_X1 u0_u7_u3_U91 (.ZN( u0_u7_u3_n111 ) , .B2( u0_u7_u3_n117 ) , .A( u0_u7_u3_n133 ) , .B1( u0_u7_u3_n176 ) );
  NAND4_X1 u0_u7_u3_U92 (.ZN( u0_out7_20 ) , .A4( u0_u7_u3_n122 ) , .A3( u0_u7_u3_n123 ) , .A1( u0_u7_u3_n175 ) , .A2( u0_u7_u3_n180 ) );
  INV_X1 u0_u7_u3_U93 (.A( u0_u7_u3_n126 ) , .ZN( u0_u7_u3_n180 ) );
  INV_X1 u0_u7_u3_U94 (.A( u0_u7_u3_n112 ) , .ZN( u0_u7_u3_n175 ) );
  NAND4_X1 u0_u7_u3_U95 (.ZN( u0_out7_1 ) , .A4( u0_u7_u3_n161 ) , .A3( u0_u7_u3_n162 ) , .A2( u0_u7_u3_n163 ) , .A1( u0_u7_u3_n185 ) );
  NAND2_X1 u0_u7_u3_U96 (.ZN( u0_u7_u3_n163 ) , .A2( u0_u7_u3_n170 ) , .A1( u0_u7_u3_n176 ) );
  AOI22_X1 u0_u7_u3_U97 (.B2( u0_u7_u3_n140 ) , .B1( u0_u7_u3_n141 ) , .A2( u0_u7_u3_n142 ) , .ZN( u0_u7_u3_n162 ) , .A1( u0_u7_u3_n177 ) );
  NAND3_X1 u0_u7_u3_U98 (.A1( u0_u7_u3_n114 ) , .ZN( u0_u7_u3_n115 ) , .A2( u0_u7_u3_n145 ) , .A3( u0_u7_u3_n153 ) );
  NAND3_X1 u0_u7_u3_U99 (.ZN( u0_u7_u3_n129 ) , .A2( u0_u7_u3_n144 ) , .A1( u0_u7_u3_n153 ) , .A3( u0_u7_u3_n182 ) );
  OAI22_X1 u0_u7_u4_U10 (.B2( u0_u7_u4_n135 ) , .ZN( u0_u7_u4_n137 ) , .B1( u0_u7_u4_n153 ) , .A1( u0_u7_u4_n155 ) , .A2( u0_u7_u4_n171 ) );
  AND3_X1 u0_u7_u4_U11 (.A2( u0_u7_u4_n134 ) , .ZN( u0_u7_u4_n135 ) , .A3( u0_u7_u4_n145 ) , .A1( u0_u7_u4_n157 ) );
  OR3_X1 u0_u7_u4_U12 (.A3( u0_u7_u4_n114 ) , .A2( u0_u7_u4_n115 ) , .A1( u0_u7_u4_n116 ) , .ZN( u0_u7_u4_n136 ) );
  AOI21_X1 u0_u7_u4_U13 (.A( u0_u7_u4_n113 ) , .ZN( u0_u7_u4_n116 ) , .B2( u0_u7_u4_n173 ) , .B1( u0_u7_u4_n174 ) );
  AOI21_X1 u0_u7_u4_U14 (.ZN( u0_u7_u4_n115 ) , .B2( u0_u7_u4_n145 ) , .B1( u0_u7_u4_n146 ) , .A( u0_u7_u4_n156 ) );
  OAI22_X1 u0_u7_u4_U15 (.ZN( u0_u7_u4_n114 ) , .A2( u0_u7_u4_n121 ) , .B1( u0_u7_u4_n160 ) , .B2( u0_u7_u4_n170 ) , .A1( u0_u7_u4_n171 ) );
  NAND2_X1 u0_u7_u4_U16 (.ZN( u0_u7_u4_n132 ) , .A2( u0_u7_u4_n170 ) , .A1( u0_u7_u4_n173 ) );
  AOI21_X1 u0_u7_u4_U17 (.B2( u0_u7_u4_n160 ) , .B1( u0_u7_u4_n161 ) , .ZN( u0_u7_u4_n162 ) , .A( u0_u7_u4_n170 ) );
  AOI21_X1 u0_u7_u4_U18 (.ZN( u0_u7_u4_n107 ) , .B2( u0_u7_u4_n143 ) , .A( u0_u7_u4_n174 ) , .B1( u0_u7_u4_n184 ) );
  AOI21_X1 u0_u7_u4_U19 (.B2( u0_u7_u4_n158 ) , .B1( u0_u7_u4_n159 ) , .ZN( u0_u7_u4_n163 ) , .A( u0_u7_u4_n174 ) );
  AOI21_X1 u0_u7_u4_U20 (.A( u0_u7_u4_n153 ) , .B2( u0_u7_u4_n154 ) , .B1( u0_u7_u4_n155 ) , .ZN( u0_u7_u4_n165 ) );
  AOI21_X1 u0_u7_u4_U21 (.A( u0_u7_u4_n156 ) , .B2( u0_u7_u4_n157 ) , .ZN( u0_u7_u4_n164 ) , .B1( u0_u7_u4_n184 ) );
  INV_X1 u0_u7_u4_U22 (.A( u0_u7_u4_n138 ) , .ZN( u0_u7_u4_n170 ) );
  AND2_X1 u0_u7_u4_U23 (.A2( u0_u7_u4_n120 ) , .ZN( u0_u7_u4_n155 ) , .A1( u0_u7_u4_n160 ) );
  INV_X1 u0_u7_u4_U24 (.A( u0_u7_u4_n156 ) , .ZN( u0_u7_u4_n175 ) );
  NAND2_X1 u0_u7_u4_U25 (.A2( u0_u7_u4_n118 ) , .ZN( u0_u7_u4_n131 ) , .A1( u0_u7_u4_n147 ) );
  NAND2_X1 u0_u7_u4_U26 (.A1( u0_u7_u4_n119 ) , .A2( u0_u7_u4_n120 ) , .ZN( u0_u7_u4_n130 ) );
  NAND2_X1 u0_u7_u4_U27 (.ZN( u0_u7_u4_n117 ) , .A2( u0_u7_u4_n118 ) , .A1( u0_u7_u4_n148 ) );
  NAND2_X1 u0_u7_u4_U28 (.ZN( u0_u7_u4_n129 ) , .A1( u0_u7_u4_n134 ) , .A2( u0_u7_u4_n148 ) );
  AND3_X1 u0_u7_u4_U29 (.A1( u0_u7_u4_n119 ) , .A2( u0_u7_u4_n143 ) , .A3( u0_u7_u4_n154 ) , .ZN( u0_u7_u4_n161 ) );
  NOR2_X1 u0_u7_u4_U3 (.ZN( u0_u7_u4_n121 ) , .A1( u0_u7_u4_n181 ) , .A2( u0_u7_u4_n182 ) );
  AND2_X1 u0_u7_u4_U30 (.A1( u0_u7_u4_n145 ) , .A2( u0_u7_u4_n147 ) , .ZN( u0_u7_u4_n159 ) );
  INV_X1 u0_u7_u4_U31 (.A( u0_u7_u4_n158 ) , .ZN( u0_u7_u4_n182 ) );
  INV_X1 u0_u7_u4_U32 (.ZN( u0_u7_u4_n181 ) , .A( u0_u7_u4_n96 ) );
  INV_X1 u0_u7_u4_U33 (.A( u0_u7_u4_n144 ) , .ZN( u0_u7_u4_n179 ) );
  INV_X1 u0_u7_u4_U34 (.A( u0_u7_u4_n157 ) , .ZN( u0_u7_u4_n178 ) );
  NAND2_X1 u0_u7_u4_U35 (.A2( u0_u7_u4_n154 ) , .A1( u0_u7_u4_n96 ) , .ZN( u0_u7_u4_n97 ) );
  INV_X1 u0_u7_u4_U36 (.ZN( u0_u7_u4_n186 ) , .A( u0_u7_u4_n95 ) );
  OAI221_X1 u0_u7_u4_U37 (.C1( u0_u7_u4_n134 ) , .B1( u0_u7_u4_n158 ) , .B2( u0_u7_u4_n171 ) , .C2( u0_u7_u4_n173 ) , .A( u0_u7_u4_n94 ) , .ZN( u0_u7_u4_n95 ) );
  AOI222_X1 u0_u7_u4_U38 (.B2( u0_u7_u4_n132 ) , .A1( u0_u7_u4_n138 ) , .C2( u0_u7_u4_n175 ) , .A2( u0_u7_u4_n179 ) , .C1( u0_u7_u4_n181 ) , .B1( u0_u7_u4_n185 ) , .ZN( u0_u7_u4_n94 ) );
  INV_X1 u0_u7_u4_U39 (.A( u0_u7_u4_n113 ) , .ZN( u0_u7_u4_n185 ) );
  INV_X1 u0_u7_u4_U4 (.A( u0_u7_u4_n117 ) , .ZN( u0_u7_u4_n184 ) );
  INV_X1 u0_u7_u4_U40 (.A( u0_u7_u4_n143 ) , .ZN( u0_u7_u4_n183 ) );
  NOR2_X1 u0_u7_u4_U41 (.ZN( u0_u7_u4_n138 ) , .A1( u0_u7_u4_n168 ) , .A2( u0_u7_u4_n169 ) );
  NOR2_X1 u0_u7_u4_U42 (.A1( u0_u7_u4_n150 ) , .A2( u0_u7_u4_n152 ) , .ZN( u0_u7_u4_n153 ) );
  NOR2_X1 u0_u7_u4_U43 (.A2( u0_u7_u4_n128 ) , .A1( u0_u7_u4_n138 ) , .ZN( u0_u7_u4_n156 ) );
  AOI22_X1 u0_u7_u4_U44 (.B2( u0_u7_u4_n122 ) , .A1( u0_u7_u4_n123 ) , .ZN( u0_u7_u4_n124 ) , .B1( u0_u7_u4_n128 ) , .A2( u0_u7_u4_n172 ) );
  NAND2_X1 u0_u7_u4_U45 (.A2( u0_u7_u4_n120 ) , .ZN( u0_u7_u4_n123 ) , .A1( u0_u7_u4_n161 ) );
  INV_X1 u0_u7_u4_U46 (.A( u0_u7_u4_n153 ) , .ZN( u0_u7_u4_n172 ) );
  AOI22_X1 u0_u7_u4_U47 (.B2( u0_u7_u4_n132 ) , .A2( u0_u7_u4_n133 ) , .ZN( u0_u7_u4_n140 ) , .A1( u0_u7_u4_n150 ) , .B1( u0_u7_u4_n179 ) );
  NAND2_X1 u0_u7_u4_U48 (.ZN( u0_u7_u4_n133 ) , .A2( u0_u7_u4_n146 ) , .A1( u0_u7_u4_n154 ) );
  NAND2_X1 u0_u7_u4_U49 (.A1( u0_u7_u4_n103 ) , .ZN( u0_u7_u4_n154 ) , .A2( u0_u7_u4_n98 ) );
  NOR4_X1 u0_u7_u4_U5 (.A4( u0_u7_u4_n106 ) , .A3( u0_u7_u4_n107 ) , .A2( u0_u7_u4_n108 ) , .A1( u0_u7_u4_n109 ) , .ZN( u0_u7_u4_n110 ) );
  NAND2_X1 u0_u7_u4_U50 (.A1( u0_u7_u4_n101 ) , .ZN( u0_u7_u4_n158 ) , .A2( u0_u7_u4_n99 ) );
  AOI21_X1 u0_u7_u4_U51 (.ZN( u0_u7_u4_n127 ) , .A( u0_u7_u4_n136 ) , .B2( u0_u7_u4_n150 ) , .B1( u0_u7_u4_n180 ) );
  INV_X1 u0_u7_u4_U52 (.A( u0_u7_u4_n160 ) , .ZN( u0_u7_u4_n180 ) );
  NAND2_X1 u0_u7_u4_U53 (.A2( u0_u7_u4_n104 ) , .A1( u0_u7_u4_n105 ) , .ZN( u0_u7_u4_n146 ) );
  NAND2_X1 u0_u7_u4_U54 (.A2( u0_u7_u4_n101 ) , .A1( u0_u7_u4_n102 ) , .ZN( u0_u7_u4_n160 ) );
  NAND2_X1 u0_u7_u4_U55 (.ZN( u0_u7_u4_n134 ) , .A1( u0_u7_u4_n98 ) , .A2( u0_u7_u4_n99 ) );
  NAND2_X1 u0_u7_u4_U56 (.A1( u0_u7_u4_n103 ) , .A2( u0_u7_u4_n104 ) , .ZN( u0_u7_u4_n143 ) );
  NAND2_X1 u0_u7_u4_U57 (.A2( u0_u7_u4_n105 ) , .ZN( u0_u7_u4_n145 ) , .A1( u0_u7_u4_n98 ) );
  NAND2_X1 u0_u7_u4_U58 (.A1( u0_u7_u4_n100 ) , .A2( u0_u7_u4_n105 ) , .ZN( u0_u7_u4_n120 ) );
  NAND2_X1 u0_u7_u4_U59 (.A1( u0_u7_u4_n102 ) , .A2( u0_u7_u4_n104 ) , .ZN( u0_u7_u4_n148 ) );
  AOI21_X1 u0_u7_u4_U6 (.ZN( u0_u7_u4_n106 ) , .B2( u0_u7_u4_n146 ) , .B1( u0_u7_u4_n158 ) , .A( u0_u7_u4_n170 ) );
  NAND2_X1 u0_u7_u4_U60 (.A2( u0_u7_u4_n100 ) , .A1( u0_u7_u4_n103 ) , .ZN( u0_u7_u4_n157 ) );
  INV_X1 u0_u7_u4_U61 (.A( u0_u7_u4_n150 ) , .ZN( u0_u7_u4_n173 ) );
  INV_X1 u0_u7_u4_U62 (.A( u0_u7_u4_n152 ) , .ZN( u0_u7_u4_n171 ) );
  NAND2_X1 u0_u7_u4_U63 (.A1( u0_u7_u4_n100 ) , .ZN( u0_u7_u4_n118 ) , .A2( u0_u7_u4_n99 ) );
  NAND2_X1 u0_u7_u4_U64 (.A2( u0_u7_u4_n100 ) , .A1( u0_u7_u4_n102 ) , .ZN( u0_u7_u4_n144 ) );
  NAND2_X1 u0_u7_u4_U65 (.A2( u0_u7_u4_n101 ) , .A1( u0_u7_u4_n105 ) , .ZN( u0_u7_u4_n96 ) );
  INV_X1 u0_u7_u4_U66 (.A( u0_u7_u4_n128 ) , .ZN( u0_u7_u4_n174 ) );
  NAND2_X1 u0_u7_u4_U67 (.A2( u0_u7_u4_n102 ) , .ZN( u0_u7_u4_n119 ) , .A1( u0_u7_u4_n98 ) );
  NAND2_X1 u0_u7_u4_U68 (.A2( u0_u7_u4_n101 ) , .A1( u0_u7_u4_n103 ) , .ZN( u0_u7_u4_n147 ) );
  NAND2_X1 u0_u7_u4_U69 (.A2( u0_u7_u4_n104 ) , .ZN( u0_u7_u4_n113 ) , .A1( u0_u7_u4_n99 ) );
  AOI21_X1 u0_u7_u4_U7 (.ZN( u0_u7_u4_n108 ) , .B2( u0_u7_u4_n134 ) , .B1( u0_u7_u4_n155 ) , .A( u0_u7_u4_n156 ) );
  NOR2_X1 u0_u7_u4_U70 (.A2( u0_u7_X_28 ) , .ZN( u0_u7_u4_n150 ) , .A1( u0_u7_u4_n168 ) );
  NOR2_X1 u0_u7_u4_U71 (.A2( u0_u7_X_29 ) , .ZN( u0_u7_u4_n152 ) , .A1( u0_u7_u4_n169 ) );
  NOR2_X1 u0_u7_u4_U72 (.A2( u0_u7_X_26 ) , .ZN( u0_u7_u4_n100 ) , .A1( u0_u7_u4_n177 ) );
  NOR2_X1 u0_u7_u4_U73 (.A2( u0_u7_X_30 ) , .ZN( u0_u7_u4_n105 ) , .A1( u0_u7_u4_n176 ) );
  NOR2_X1 u0_u7_u4_U74 (.A2( u0_u7_X_28 ) , .A1( u0_u7_X_29 ) , .ZN( u0_u7_u4_n128 ) );
  NOR2_X1 u0_u7_u4_U75 (.A2( u0_u7_X_25 ) , .A1( u0_u7_X_26 ) , .ZN( u0_u7_u4_n98 ) );
  NOR2_X1 u0_u7_u4_U76 (.A2( u0_u7_X_27 ) , .A1( u0_u7_X_30 ) , .ZN( u0_u7_u4_n102 ) );
  AND2_X1 u0_u7_u4_U77 (.A2( u0_u7_X_25 ) , .A1( u0_u7_X_26 ) , .ZN( u0_u7_u4_n104 ) );
  AND2_X1 u0_u7_u4_U78 (.A1( u0_u7_X_30 ) , .A2( u0_u7_u4_n176 ) , .ZN( u0_u7_u4_n99 ) );
  AND2_X1 u0_u7_u4_U79 (.A1( u0_u7_X_26 ) , .ZN( u0_u7_u4_n101 ) , .A2( u0_u7_u4_n177 ) );
  AOI21_X1 u0_u7_u4_U8 (.ZN( u0_u7_u4_n109 ) , .A( u0_u7_u4_n153 ) , .B1( u0_u7_u4_n159 ) , .B2( u0_u7_u4_n184 ) );
  AND2_X1 u0_u7_u4_U80 (.A1( u0_u7_X_27 ) , .A2( u0_u7_X_30 ) , .ZN( u0_u7_u4_n103 ) );
  INV_X1 u0_u7_u4_U81 (.A( u0_u7_X_28 ) , .ZN( u0_u7_u4_n169 ) );
  INV_X1 u0_u7_u4_U82 (.A( u0_u7_X_29 ) , .ZN( u0_u7_u4_n168 ) );
  INV_X1 u0_u7_u4_U83 (.A( u0_u7_X_25 ) , .ZN( u0_u7_u4_n177 ) );
  INV_X1 u0_u7_u4_U84 (.A( u0_u7_X_27 ) , .ZN( u0_u7_u4_n176 ) );
  NAND4_X1 u0_u7_u4_U85 (.ZN( u0_out7_25 ) , .A4( u0_u7_u4_n139 ) , .A3( u0_u7_u4_n140 ) , .A2( u0_u7_u4_n141 ) , .A1( u0_u7_u4_n142 ) );
  OAI21_X1 u0_u7_u4_U86 (.A( u0_u7_u4_n128 ) , .B2( u0_u7_u4_n129 ) , .B1( u0_u7_u4_n130 ) , .ZN( u0_u7_u4_n142 ) );
  OAI21_X1 u0_u7_u4_U87 (.B2( u0_u7_u4_n131 ) , .ZN( u0_u7_u4_n141 ) , .A( u0_u7_u4_n175 ) , .B1( u0_u7_u4_n183 ) );
  NAND4_X1 u0_u7_u4_U88 (.ZN( u0_out7_14 ) , .A4( u0_u7_u4_n124 ) , .A3( u0_u7_u4_n125 ) , .A2( u0_u7_u4_n126 ) , .A1( u0_u7_u4_n127 ) );
  AOI22_X1 u0_u7_u4_U89 (.B2( u0_u7_u4_n117 ) , .ZN( u0_u7_u4_n126 ) , .A1( u0_u7_u4_n129 ) , .B1( u0_u7_u4_n152 ) , .A2( u0_u7_u4_n175 ) );
  AOI211_X1 u0_u7_u4_U9 (.B( u0_u7_u4_n136 ) , .A( u0_u7_u4_n137 ) , .C2( u0_u7_u4_n138 ) , .ZN( u0_u7_u4_n139 ) , .C1( u0_u7_u4_n182 ) );
  AOI22_X1 u0_u7_u4_U90 (.ZN( u0_u7_u4_n125 ) , .B2( u0_u7_u4_n131 ) , .A2( u0_u7_u4_n132 ) , .B1( u0_u7_u4_n138 ) , .A1( u0_u7_u4_n178 ) );
  NAND4_X1 u0_u7_u4_U91 (.ZN( u0_out7_8 ) , .A4( u0_u7_u4_n110 ) , .A3( u0_u7_u4_n111 ) , .A2( u0_u7_u4_n112 ) , .A1( u0_u7_u4_n186 ) );
  NAND2_X1 u0_u7_u4_U92 (.ZN( u0_u7_u4_n112 ) , .A2( u0_u7_u4_n130 ) , .A1( u0_u7_u4_n150 ) );
  AOI22_X1 u0_u7_u4_U93 (.ZN( u0_u7_u4_n111 ) , .B2( u0_u7_u4_n132 ) , .A1( u0_u7_u4_n152 ) , .B1( u0_u7_u4_n178 ) , .A2( u0_u7_u4_n97 ) );
  AOI22_X1 u0_u7_u4_U94 (.B2( u0_u7_u4_n149 ) , .B1( u0_u7_u4_n150 ) , .A2( u0_u7_u4_n151 ) , .A1( u0_u7_u4_n152 ) , .ZN( u0_u7_u4_n167 ) );
  NOR4_X1 u0_u7_u4_U95 (.A4( u0_u7_u4_n162 ) , .A3( u0_u7_u4_n163 ) , .A2( u0_u7_u4_n164 ) , .A1( u0_u7_u4_n165 ) , .ZN( u0_u7_u4_n166 ) );
  NAND3_X1 u0_u7_u4_U96 (.ZN( u0_out7_3 ) , .A3( u0_u7_u4_n166 ) , .A1( u0_u7_u4_n167 ) , .A2( u0_u7_u4_n186 ) );
  NAND3_X1 u0_u7_u4_U97 (.A3( u0_u7_u4_n146 ) , .A2( u0_u7_u4_n147 ) , .A1( u0_u7_u4_n148 ) , .ZN( u0_u7_u4_n149 ) );
  NAND3_X1 u0_u7_u4_U98 (.A3( u0_u7_u4_n143 ) , .A2( u0_u7_u4_n144 ) , .A1( u0_u7_u4_n145 ) , .ZN( u0_u7_u4_n151 ) );
  NAND3_X1 u0_u7_u4_U99 (.A3( u0_u7_u4_n121 ) , .ZN( u0_u7_u4_n122 ) , .A2( u0_u7_u4_n144 ) , .A1( u0_u7_u4_n154 ) );
  INV_X1 u0_u7_u5_U10 (.A( u0_u7_u5_n121 ) , .ZN( u0_u7_u5_n177 ) );
  NOR3_X1 u0_u7_u5_U100 (.A3( u0_u7_u5_n141 ) , .A1( u0_u7_u5_n142 ) , .ZN( u0_u7_u5_n143 ) , .A2( u0_u7_u5_n191 ) );
  NAND4_X1 u0_u7_u5_U101 (.ZN( u0_out7_4 ) , .A4( u0_u7_u5_n112 ) , .A2( u0_u7_u5_n113 ) , .A1( u0_u7_u5_n114 ) , .A3( u0_u7_u5_n195 ) );
  AOI211_X1 u0_u7_u5_U102 (.A( u0_u7_u5_n110 ) , .C1( u0_u7_u5_n111 ) , .ZN( u0_u7_u5_n112 ) , .B( u0_u7_u5_n118 ) , .C2( u0_u7_u5_n177 ) );
  AOI222_X1 u0_u7_u5_U103 (.ZN( u0_u7_u5_n113 ) , .A1( u0_u7_u5_n131 ) , .C1( u0_u7_u5_n148 ) , .B2( u0_u7_u5_n174 ) , .C2( u0_u7_u5_n178 ) , .A2( u0_u7_u5_n179 ) , .B1( u0_u7_u5_n99 ) );
  NAND3_X1 u0_u7_u5_U104 (.A2( u0_u7_u5_n154 ) , .A3( u0_u7_u5_n158 ) , .A1( u0_u7_u5_n161 ) , .ZN( u0_u7_u5_n99 ) );
  NOR2_X1 u0_u7_u5_U11 (.ZN( u0_u7_u5_n160 ) , .A2( u0_u7_u5_n173 ) , .A1( u0_u7_u5_n177 ) );
  INV_X1 u0_u7_u5_U12 (.A( u0_u7_u5_n150 ) , .ZN( u0_u7_u5_n174 ) );
  AOI21_X1 u0_u7_u5_U13 (.A( u0_u7_u5_n160 ) , .B2( u0_u7_u5_n161 ) , .ZN( u0_u7_u5_n162 ) , .B1( u0_u7_u5_n192 ) );
  INV_X1 u0_u7_u5_U14 (.A( u0_u7_u5_n159 ) , .ZN( u0_u7_u5_n192 ) );
  AOI21_X1 u0_u7_u5_U15 (.A( u0_u7_u5_n156 ) , .B2( u0_u7_u5_n157 ) , .B1( u0_u7_u5_n158 ) , .ZN( u0_u7_u5_n163 ) );
  AOI21_X1 u0_u7_u5_U16 (.B2( u0_u7_u5_n139 ) , .B1( u0_u7_u5_n140 ) , .ZN( u0_u7_u5_n141 ) , .A( u0_u7_u5_n150 ) );
  OAI21_X1 u0_u7_u5_U17 (.A( u0_u7_u5_n133 ) , .B2( u0_u7_u5_n134 ) , .B1( u0_u7_u5_n135 ) , .ZN( u0_u7_u5_n142 ) );
  OAI21_X1 u0_u7_u5_U18 (.ZN( u0_u7_u5_n133 ) , .B2( u0_u7_u5_n147 ) , .A( u0_u7_u5_n173 ) , .B1( u0_u7_u5_n188 ) );
  NAND2_X1 u0_u7_u5_U19 (.A2( u0_u7_u5_n119 ) , .A1( u0_u7_u5_n123 ) , .ZN( u0_u7_u5_n137 ) );
  INV_X1 u0_u7_u5_U20 (.A( u0_u7_u5_n155 ) , .ZN( u0_u7_u5_n194 ) );
  NAND2_X1 u0_u7_u5_U21 (.A1( u0_u7_u5_n121 ) , .ZN( u0_u7_u5_n132 ) , .A2( u0_u7_u5_n172 ) );
  NAND2_X1 u0_u7_u5_U22 (.A2( u0_u7_u5_n122 ) , .ZN( u0_u7_u5_n136 ) , .A1( u0_u7_u5_n154 ) );
  NAND2_X1 u0_u7_u5_U23 (.A2( u0_u7_u5_n119 ) , .A1( u0_u7_u5_n120 ) , .ZN( u0_u7_u5_n159 ) );
  INV_X1 u0_u7_u5_U24 (.A( u0_u7_u5_n156 ) , .ZN( u0_u7_u5_n175 ) );
  INV_X1 u0_u7_u5_U25 (.A( u0_u7_u5_n158 ) , .ZN( u0_u7_u5_n188 ) );
  INV_X1 u0_u7_u5_U26 (.A( u0_u7_u5_n152 ) , .ZN( u0_u7_u5_n179 ) );
  INV_X1 u0_u7_u5_U27 (.A( u0_u7_u5_n140 ) , .ZN( u0_u7_u5_n182 ) );
  INV_X1 u0_u7_u5_U28 (.A( u0_u7_u5_n151 ) , .ZN( u0_u7_u5_n183 ) );
  INV_X1 u0_u7_u5_U29 (.A( u0_u7_u5_n123 ) , .ZN( u0_u7_u5_n185 ) );
  NOR2_X1 u0_u7_u5_U3 (.ZN( u0_u7_u5_n134 ) , .A1( u0_u7_u5_n183 ) , .A2( u0_u7_u5_n190 ) );
  INV_X1 u0_u7_u5_U30 (.A( u0_u7_u5_n161 ) , .ZN( u0_u7_u5_n184 ) );
  INV_X1 u0_u7_u5_U31 (.A( u0_u7_u5_n139 ) , .ZN( u0_u7_u5_n189 ) );
  INV_X1 u0_u7_u5_U32 (.A( u0_u7_u5_n157 ) , .ZN( u0_u7_u5_n190 ) );
  INV_X1 u0_u7_u5_U33 (.A( u0_u7_u5_n120 ) , .ZN( u0_u7_u5_n193 ) );
  NAND2_X1 u0_u7_u5_U34 (.ZN( u0_u7_u5_n111 ) , .A1( u0_u7_u5_n140 ) , .A2( u0_u7_u5_n155 ) );
  NOR2_X1 u0_u7_u5_U35 (.ZN( u0_u7_u5_n100 ) , .A1( u0_u7_u5_n170 ) , .A2( u0_u7_u5_n180 ) );
  INV_X1 u0_u7_u5_U36 (.A( u0_u7_u5_n117 ) , .ZN( u0_u7_u5_n196 ) );
  OAI221_X1 u0_u7_u5_U37 (.A( u0_u7_u5_n116 ) , .ZN( u0_u7_u5_n117 ) , .B2( u0_u7_u5_n119 ) , .C1( u0_u7_u5_n153 ) , .C2( u0_u7_u5_n158 ) , .B1( u0_u7_u5_n172 ) );
  AOI222_X1 u0_u7_u5_U38 (.ZN( u0_u7_u5_n116 ) , .B2( u0_u7_u5_n145 ) , .C1( u0_u7_u5_n148 ) , .A2( u0_u7_u5_n174 ) , .C2( u0_u7_u5_n177 ) , .B1( u0_u7_u5_n187 ) , .A1( u0_u7_u5_n193 ) );
  INV_X1 u0_u7_u5_U39 (.A( u0_u7_u5_n115 ) , .ZN( u0_u7_u5_n187 ) );
  INV_X1 u0_u7_u5_U4 (.A( u0_u7_u5_n138 ) , .ZN( u0_u7_u5_n191 ) );
  AOI22_X1 u0_u7_u5_U40 (.B2( u0_u7_u5_n131 ) , .A2( u0_u7_u5_n146 ) , .ZN( u0_u7_u5_n169 ) , .B1( u0_u7_u5_n174 ) , .A1( u0_u7_u5_n185 ) );
  NOR2_X1 u0_u7_u5_U41 (.A1( u0_u7_u5_n146 ) , .ZN( u0_u7_u5_n150 ) , .A2( u0_u7_u5_n173 ) );
  AOI21_X1 u0_u7_u5_U42 (.A( u0_u7_u5_n118 ) , .B2( u0_u7_u5_n145 ) , .ZN( u0_u7_u5_n168 ) , .B1( u0_u7_u5_n186 ) );
  INV_X1 u0_u7_u5_U43 (.A( u0_u7_u5_n122 ) , .ZN( u0_u7_u5_n186 ) );
  NOR2_X1 u0_u7_u5_U44 (.A1( u0_u7_u5_n146 ) , .ZN( u0_u7_u5_n152 ) , .A2( u0_u7_u5_n176 ) );
  NOR2_X1 u0_u7_u5_U45 (.A1( u0_u7_u5_n115 ) , .ZN( u0_u7_u5_n118 ) , .A2( u0_u7_u5_n153 ) );
  NOR2_X1 u0_u7_u5_U46 (.A2( u0_u7_u5_n145 ) , .ZN( u0_u7_u5_n156 ) , .A1( u0_u7_u5_n174 ) );
  NOR2_X1 u0_u7_u5_U47 (.ZN( u0_u7_u5_n121 ) , .A2( u0_u7_u5_n145 ) , .A1( u0_u7_u5_n176 ) );
  AOI22_X1 u0_u7_u5_U48 (.ZN( u0_u7_u5_n114 ) , .A2( u0_u7_u5_n137 ) , .A1( u0_u7_u5_n145 ) , .B2( u0_u7_u5_n175 ) , .B1( u0_u7_u5_n193 ) );
  OAI211_X1 u0_u7_u5_U49 (.B( u0_u7_u5_n124 ) , .A( u0_u7_u5_n125 ) , .C2( u0_u7_u5_n126 ) , .C1( u0_u7_u5_n127 ) , .ZN( u0_u7_u5_n128 ) );
  OAI21_X1 u0_u7_u5_U5 (.B2( u0_u7_u5_n136 ) , .B1( u0_u7_u5_n137 ) , .ZN( u0_u7_u5_n138 ) , .A( u0_u7_u5_n177 ) );
  NOR3_X1 u0_u7_u5_U50 (.ZN( u0_u7_u5_n127 ) , .A1( u0_u7_u5_n136 ) , .A3( u0_u7_u5_n148 ) , .A2( u0_u7_u5_n182 ) );
  OAI21_X1 u0_u7_u5_U51 (.ZN( u0_u7_u5_n124 ) , .A( u0_u7_u5_n177 ) , .B2( u0_u7_u5_n183 ) , .B1( u0_u7_u5_n189 ) );
  OAI21_X1 u0_u7_u5_U52 (.ZN( u0_u7_u5_n125 ) , .A( u0_u7_u5_n174 ) , .B2( u0_u7_u5_n185 ) , .B1( u0_u7_u5_n190 ) );
  AOI21_X1 u0_u7_u5_U53 (.A( u0_u7_u5_n153 ) , .B2( u0_u7_u5_n154 ) , .B1( u0_u7_u5_n155 ) , .ZN( u0_u7_u5_n164 ) );
  AOI21_X1 u0_u7_u5_U54 (.ZN( u0_u7_u5_n110 ) , .B1( u0_u7_u5_n122 ) , .B2( u0_u7_u5_n139 ) , .A( u0_u7_u5_n153 ) );
  INV_X1 u0_u7_u5_U55 (.A( u0_u7_u5_n153 ) , .ZN( u0_u7_u5_n176 ) );
  INV_X1 u0_u7_u5_U56 (.A( u0_u7_u5_n126 ) , .ZN( u0_u7_u5_n173 ) );
  AND2_X1 u0_u7_u5_U57 (.A2( u0_u7_u5_n104 ) , .A1( u0_u7_u5_n107 ) , .ZN( u0_u7_u5_n147 ) );
  AND2_X1 u0_u7_u5_U58 (.A2( u0_u7_u5_n104 ) , .A1( u0_u7_u5_n108 ) , .ZN( u0_u7_u5_n148 ) );
  NAND2_X1 u0_u7_u5_U59 (.A1( u0_u7_u5_n105 ) , .A2( u0_u7_u5_n106 ) , .ZN( u0_u7_u5_n158 ) );
  INV_X1 u0_u7_u5_U6 (.A( u0_u7_u5_n135 ) , .ZN( u0_u7_u5_n178 ) );
  NAND2_X1 u0_u7_u5_U60 (.A2( u0_u7_u5_n108 ) , .A1( u0_u7_u5_n109 ) , .ZN( u0_u7_u5_n139 ) );
  NAND2_X1 u0_u7_u5_U61 (.A1( u0_u7_u5_n106 ) , .A2( u0_u7_u5_n108 ) , .ZN( u0_u7_u5_n119 ) );
  NAND2_X1 u0_u7_u5_U62 (.A2( u0_u7_u5_n103 ) , .A1( u0_u7_u5_n105 ) , .ZN( u0_u7_u5_n140 ) );
  NAND2_X1 u0_u7_u5_U63 (.A2( u0_u7_u5_n104 ) , .A1( u0_u7_u5_n105 ) , .ZN( u0_u7_u5_n155 ) );
  NAND2_X1 u0_u7_u5_U64 (.A2( u0_u7_u5_n106 ) , .A1( u0_u7_u5_n107 ) , .ZN( u0_u7_u5_n122 ) );
  NAND2_X1 u0_u7_u5_U65 (.A2( u0_u7_u5_n100 ) , .A1( u0_u7_u5_n106 ) , .ZN( u0_u7_u5_n115 ) );
  NAND2_X1 u0_u7_u5_U66 (.A2( u0_u7_u5_n100 ) , .A1( u0_u7_u5_n103 ) , .ZN( u0_u7_u5_n161 ) );
  NAND2_X1 u0_u7_u5_U67 (.A1( u0_u7_u5_n105 ) , .A2( u0_u7_u5_n109 ) , .ZN( u0_u7_u5_n154 ) );
  INV_X1 u0_u7_u5_U68 (.A( u0_u7_u5_n146 ) , .ZN( u0_u7_u5_n172 ) );
  NAND2_X1 u0_u7_u5_U69 (.A1( u0_u7_u5_n103 ) , .A2( u0_u7_u5_n108 ) , .ZN( u0_u7_u5_n123 ) );
  OAI22_X1 u0_u7_u5_U7 (.B2( u0_u7_u5_n149 ) , .B1( u0_u7_u5_n150 ) , .A2( u0_u7_u5_n151 ) , .A1( u0_u7_u5_n152 ) , .ZN( u0_u7_u5_n165 ) );
  NAND2_X1 u0_u7_u5_U70 (.A2( u0_u7_u5_n103 ) , .A1( u0_u7_u5_n107 ) , .ZN( u0_u7_u5_n151 ) );
  NAND2_X1 u0_u7_u5_U71 (.A2( u0_u7_u5_n107 ) , .A1( u0_u7_u5_n109 ) , .ZN( u0_u7_u5_n120 ) );
  NAND2_X1 u0_u7_u5_U72 (.A2( u0_u7_u5_n100 ) , .A1( u0_u7_u5_n109 ) , .ZN( u0_u7_u5_n157 ) );
  AND2_X1 u0_u7_u5_U73 (.A2( u0_u7_u5_n100 ) , .A1( u0_u7_u5_n104 ) , .ZN( u0_u7_u5_n131 ) );
  INV_X1 u0_u7_u5_U74 (.A( u0_u7_u5_n102 ) , .ZN( u0_u7_u5_n195 ) );
  OAI221_X1 u0_u7_u5_U75 (.A( u0_u7_u5_n101 ) , .ZN( u0_u7_u5_n102 ) , .C2( u0_u7_u5_n115 ) , .C1( u0_u7_u5_n126 ) , .B1( u0_u7_u5_n134 ) , .B2( u0_u7_u5_n160 ) );
  OAI21_X1 u0_u7_u5_U76 (.ZN( u0_u7_u5_n101 ) , .B1( u0_u7_u5_n137 ) , .A( u0_u7_u5_n146 ) , .B2( u0_u7_u5_n147 ) );
  NOR2_X1 u0_u7_u5_U77 (.A2( u0_u7_X_34 ) , .A1( u0_u7_X_35 ) , .ZN( u0_u7_u5_n145 ) );
  NOR2_X1 u0_u7_u5_U78 (.A2( u0_u7_X_34 ) , .ZN( u0_u7_u5_n146 ) , .A1( u0_u7_u5_n171 ) );
  NOR2_X1 u0_u7_u5_U79 (.A2( u0_u7_X_31 ) , .A1( u0_u7_X_32 ) , .ZN( u0_u7_u5_n103 ) );
  NOR3_X1 u0_u7_u5_U8 (.A2( u0_u7_u5_n147 ) , .A1( u0_u7_u5_n148 ) , .ZN( u0_u7_u5_n149 ) , .A3( u0_u7_u5_n194 ) );
  NOR2_X1 u0_u7_u5_U80 (.A2( u0_u7_X_36 ) , .ZN( u0_u7_u5_n105 ) , .A1( u0_u7_u5_n180 ) );
  NOR2_X1 u0_u7_u5_U81 (.A2( u0_u7_X_33 ) , .ZN( u0_u7_u5_n108 ) , .A1( u0_u7_u5_n170 ) );
  NOR2_X1 u0_u7_u5_U82 (.A2( u0_u7_X_33 ) , .A1( u0_u7_X_36 ) , .ZN( u0_u7_u5_n107 ) );
  NOR2_X1 u0_u7_u5_U83 (.A2( u0_u7_X_31 ) , .ZN( u0_u7_u5_n104 ) , .A1( u0_u7_u5_n181 ) );
  NAND2_X1 u0_u7_u5_U84 (.A2( u0_u7_X_34 ) , .A1( u0_u7_X_35 ) , .ZN( u0_u7_u5_n153 ) );
  NAND2_X1 u0_u7_u5_U85 (.A1( u0_u7_X_34 ) , .ZN( u0_u7_u5_n126 ) , .A2( u0_u7_u5_n171 ) );
  AND2_X1 u0_u7_u5_U86 (.A1( u0_u7_X_31 ) , .A2( u0_u7_X_32 ) , .ZN( u0_u7_u5_n106 ) );
  AND2_X1 u0_u7_u5_U87 (.A1( u0_u7_X_31 ) , .ZN( u0_u7_u5_n109 ) , .A2( u0_u7_u5_n181 ) );
  INV_X1 u0_u7_u5_U88 (.A( u0_u7_X_33 ) , .ZN( u0_u7_u5_n180 ) );
  INV_X1 u0_u7_u5_U89 (.A( u0_u7_X_35 ) , .ZN( u0_u7_u5_n171 ) );
  NOR2_X1 u0_u7_u5_U9 (.ZN( u0_u7_u5_n135 ) , .A1( u0_u7_u5_n173 ) , .A2( u0_u7_u5_n176 ) );
  INV_X1 u0_u7_u5_U90 (.A( u0_u7_X_36 ) , .ZN( u0_u7_u5_n170 ) );
  INV_X1 u0_u7_u5_U91 (.A( u0_u7_X_32 ) , .ZN( u0_u7_u5_n181 ) );
  NAND4_X1 u0_u7_u5_U92 (.ZN( u0_out7_29 ) , .A4( u0_u7_u5_n129 ) , .A3( u0_u7_u5_n130 ) , .A2( u0_u7_u5_n168 ) , .A1( u0_u7_u5_n196 ) );
  AOI221_X1 u0_u7_u5_U93 (.A( u0_u7_u5_n128 ) , .ZN( u0_u7_u5_n129 ) , .C2( u0_u7_u5_n132 ) , .B2( u0_u7_u5_n159 ) , .B1( u0_u7_u5_n176 ) , .C1( u0_u7_u5_n184 ) );
  AOI222_X1 u0_u7_u5_U94 (.ZN( u0_u7_u5_n130 ) , .A2( u0_u7_u5_n146 ) , .B1( u0_u7_u5_n147 ) , .C2( u0_u7_u5_n175 ) , .B2( u0_u7_u5_n179 ) , .A1( u0_u7_u5_n188 ) , .C1( u0_u7_u5_n194 ) );
  NAND4_X1 u0_u7_u5_U95 (.ZN( u0_out7_19 ) , .A4( u0_u7_u5_n166 ) , .A3( u0_u7_u5_n167 ) , .A2( u0_u7_u5_n168 ) , .A1( u0_u7_u5_n169 ) );
  AOI22_X1 u0_u7_u5_U96 (.B2( u0_u7_u5_n145 ) , .A2( u0_u7_u5_n146 ) , .ZN( u0_u7_u5_n167 ) , .B1( u0_u7_u5_n182 ) , .A1( u0_u7_u5_n189 ) );
  NOR4_X1 u0_u7_u5_U97 (.A4( u0_u7_u5_n162 ) , .A3( u0_u7_u5_n163 ) , .A2( u0_u7_u5_n164 ) , .A1( u0_u7_u5_n165 ) , .ZN( u0_u7_u5_n166 ) );
  NAND4_X1 u0_u7_u5_U98 (.ZN( u0_out7_11 ) , .A4( u0_u7_u5_n143 ) , .A3( u0_u7_u5_n144 ) , .A2( u0_u7_u5_n169 ) , .A1( u0_u7_u5_n196 ) );
  AOI22_X1 u0_u7_u5_U99 (.A2( u0_u7_u5_n132 ) , .ZN( u0_u7_u5_n144 ) , .B2( u0_u7_u5_n145 ) , .B1( u0_u7_u5_n184 ) , .A1( u0_u7_u5_n194 ) );
  INV_X1 u0_u7_u6_U10 (.ZN( u0_u7_u6_n172 ) , .A( u0_u7_u6_n88 ) );
  OAI21_X1 u0_u7_u6_U11 (.A( u0_u7_u6_n159 ) , .B1( u0_u7_u6_n169 ) , .B2( u0_u7_u6_n173 ) , .ZN( u0_u7_u6_n90 ) );
  AOI22_X1 u0_u7_u6_U12 (.A2( u0_u7_u6_n151 ) , .B2( u0_u7_u6_n161 ) , .A1( u0_u7_u6_n167 ) , .B1( u0_u7_u6_n170 ) , .ZN( u0_u7_u6_n89 ) );
  AOI21_X1 u0_u7_u6_U13 (.ZN( u0_u7_u6_n106 ) , .A( u0_u7_u6_n142 ) , .B2( u0_u7_u6_n159 ) , .B1( u0_u7_u6_n164 ) );
  INV_X1 u0_u7_u6_U14 (.A( u0_u7_u6_n155 ) , .ZN( u0_u7_u6_n161 ) );
  INV_X1 u0_u7_u6_U15 (.A( u0_u7_u6_n128 ) , .ZN( u0_u7_u6_n164 ) );
  NAND2_X1 u0_u7_u6_U16 (.ZN( u0_u7_u6_n110 ) , .A1( u0_u7_u6_n122 ) , .A2( u0_u7_u6_n129 ) );
  NAND2_X1 u0_u7_u6_U17 (.ZN( u0_u7_u6_n124 ) , .A2( u0_u7_u6_n146 ) , .A1( u0_u7_u6_n148 ) );
  INV_X1 u0_u7_u6_U18 (.A( u0_u7_u6_n132 ) , .ZN( u0_u7_u6_n171 ) );
  AND2_X1 u0_u7_u6_U19 (.A1( u0_u7_u6_n100 ) , .ZN( u0_u7_u6_n130 ) , .A2( u0_u7_u6_n147 ) );
  INV_X1 u0_u7_u6_U20 (.A( u0_u7_u6_n127 ) , .ZN( u0_u7_u6_n173 ) );
  INV_X1 u0_u7_u6_U21 (.A( u0_u7_u6_n121 ) , .ZN( u0_u7_u6_n167 ) );
  INV_X1 u0_u7_u6_U22 (.A( u0_u7_u6_n100 ) , .ZN( u0_u7_u6_n169 ) );
  INV_X1 u0_u7_u6_U23 (.A( u0_u7_u6_n123 ) , .ZN( u0_u7_u6_n170 ) );
  INV_X1 u0_u7_u6_U24 (.A( u0_u7_u6_n113 ) , .ZN( u0_u7_u6_n168 ) );
  AND2_X1 u0_u7_u6_U25 (.A1( u0_u7_u6_n107 ) , .A2( u0_u7_u6_n119 ) , .ZN( u0_u7_u6_n133 ) );
  AND2_X1 u0_u7_u6_U26 (.A2( u0_u7_u6_n121 ) , .A1( u0_u7_u6_n122 ) , .ZN( u0_u7_u6_n131 ) );
  AND3_X1 u0_u7_u6_U27 (.ZN( u0_u7_u6_n120 ) , .A2( u0_u7_u6_n127 ) , .A1( u0_u7_u6_n132 ) , .A3( u0_u7_u6_n145 ) );
  INV_X1 u0_u7_u6_U28 (.A( u0_u7_u6_n146 ) , .ZN( u0_u7_u6_n163 ) );
  AOI222_X1 u0_u7_u6_U29 (.ZN( u0_u7_u6_n114 ) , .A1( u0_u7_u6_n118 ) , .A2( u0_u7_u6_n126 ) , .B2( u0_u7_u6_n151 ) , .C2( u0_u7_u6_n159 ) , .C1( u0_u7_u6_n168 ) , .B1( u0_u7_u6_n169 ) );
  INV_X1 u0_u7_u6_U3 (.A( u0_u7_u6_n110 ) , .ZN( u0_u7_u6_n166 ) );
  NOR2_X1 u0_u7_u6_U30 (.A1( u0_u7_u6_n162 ) , .A2( u0_u7_u6_n165 ) , .ZN( u0_u7_u6_n98 ) );
  NAND2_X1 u0_u7_u6_U31 (.A1( u0_u7_u6_n144 ) , .ZN( u0_u7_u6_n151 ) , .A2( u0_u7_u6_n158 ) );
  NAND2_X1 u0_u7_u6_U32 (.ZN( u0_u7_u6_n132 ) , .A1( u0_u7_u6_n91 ) , .A2( u0_u7_u6_n97 ) );
  AOI22_X1 u0_u7_u6_U33 (.B2( u0_u7_u6_n110 ) , .B1( u0_u7_u6_n111 ) , .A1( u0_u7_u6_n112 ) , .ZN( u0_u7_u6_n115 ) , .A2( u0_u7_u6_n161 ) );
  NAND4_X1 u0_u7_u6_U34 (.A3( u0_u7_u6_n109 ) , .ZN( u0_u7_u6_n112 ) , .A4( u0_u7_u6_n132 ) , .A2( u0_u7_u6_n147 ) , .A1( u0_u7_u6_n166 ) );
  NOR2_X1 u0_u7_u6_U35 (.ZN( u0_u7_u6_n109 ) , .A1( u0_u7_u6_n170 ) , .A2( u0_u7_u6_n173 ) );
  NOR2_X1 u0_u7_u6_U36 (.A2( u0_u7_u6_n126 ) , .ZN( u0_u7_u6_n155 ) , .A1( u0_u7_u6_n160 ) );
  NAND2_X1 u0_u7_u6_U37 (.ZN( u0_u7_u6_n146 ) , .A2( u0_u7_u6_n94 ) , .A1( u0_u7_u6_n99 ) );
  AOI21_X1 u0_u7_u6_U38 (.A( u0_u7_u6_n144 ) , .B2( u0_u7_u6_n145 ) , .B1( u0_u7_u6_n146 ) , .ZN( u0_u7_u6_n150 ) );
  AOI211_X1 u0_u7_u6_U39 (.B( u0_u7_u6_n134 ) , .A( u0_u7_u6_n135 ) , .C1( u0_u7_u6_n136 ) , .ZN( u0_u7_u6_n137 ) , .C2( u0_u7_u6_n151 ) );
  INV_X1 u0_u7_u6_U4 (.A( u0_u7_u6_n142 ) , .ZN( u0_u7_u6_n174 ) );
  NAND4_X1 u0_u7_u6_U40 (.A4( u0_u7_u6_n127 ) , .A3( u0_u7_u6_n128 ) , .A2( u0_u7_u6_n129 ) , .A1( u0_u7_u6_n130 ) , .ZN( u0_u7_u6_n136 ) );
  AOI21_X1 u0_u7_u6_U41 (.B2( u0_u7_u6_n132 ) , .B1( u0_u7_u6_n133 ) , .ZN( u0_u7_u6_n134 ) , .A( u0_u7_u6_n158 ) );
  AOI21_X1 u0_u7_u6_U42 (.B1( u0_u7_u6_n131 ) , .ZN( u0_u7_u6_n135 ) , .A( u0_u7_u6_n144 ) , .B2( u0_u7_u6_n146 ) );
  INV_X1 u0_u7_u6_U43 (.A( u0_u7_u6_n111 ) , .ZN( u0_u7_u6_n158 ) );
  NAND2_X1 u0_u7_u6_U44 (.ZN( u0_u7_u6_n127 ) , .A1( u0_u7_u6_n91 ) , .A2( u0_u7_u6_n92 ) );
  NAND2_X1 u0_u7_u6_U45 (.ZN( u0_u7_u6_n129 ) , .A2( u0_u7_u6_n95 ) , .A1( u0_u7_u6_n96 ) );
  INV_X1 u0_u7_u6_U46 (.A( u0_u7_u6_n144 ) , .ZN( u0_u7_u6_n159 ) );
  NAND2_X1 u0_u7_u6_U47 (.ZN( u0_u7_u6_n145 ) , .A2( u0_u7_u6_n97 ) , .A1( u0_u7_u6_n98 ) );
  NAND2_X1 u0_u7_u6_U48 (.ZN( u0_u7_u6_n148 ) , .A2( u0_u7_u6_n92 ) , .A1( u0_u7_u6_n94 ) );
  NAND2_X1 u0_u7_u6_U49 (.ZN( u0_u7_u6_n108 ) , .A2( u0_u7_u6_n139 ) , .A1( u0_u7_u6_n144 ) );
  NAND2_X1 u0_u7_u6_U5 (.A2( u0_u7_u6_n143 ) , .ZN( u0_u7_u6_n152 ) , .A1( u0_u7_u6_n166 ) );
  NAND2_X1 u0_u7_u6_U50 (.ZN( u0_u7_u6_n121 ) , .A2( u0_u7_u6_n95 ) , .A1( u0_u7_u6_n97 ) );
  NAND2_X1 u0_u7_u6_U51 (.ZN( u0_u7_u6_n107 ) , .A2( u0_u7_u6_n92 ) , .A1( u0_u7_u6_n95 ) );
  AND2_X1 u0_u7_u6_U52 (.ZN( u0_u7_u6_n118 ) , .A2( u0_u7_u6_n91 ) , .A1( u0_u7_u6_n99 ) );
  NAND2_X1 u0_u7_u6_U53 (.ZN( u0_u7_u6_n147 ) , .A2( u0_u7_u6_n98 ) , .A1( u0_u7_u6_n99 ) );
  NAND2_X1 u0_u7_u6_U54 (.ZN( u0_u7_u6_n128 ) , .A1( u0_u7_u6_n94 ) , .A2( u0_u7_u6_n96 ) );
  NAND2_X1 u0_u7_u6_U55 (.ZN( u0_u7_u6_n119 ) , .A2( u0_u7_u6_n95 ) , .A1( u0_u7_u6_n99 ) );
  NAND2_X1 u0_u7_u6_U56 (.ZN( u0_u7_u6_n123 ) , .A2( u0_u7_u6_n91 ) , .A1( u0_u7_u6_n96 ) );
  NAND2_X1 u0_u7_u6_U57 (.ZN( u0_u7_u6_n100 ) , .A2( u0_u7_u6_n92 ) , .A1( u0_u7_u6_n98 ) );
  NAND2_X1 u0_u7_u6_U58 (.ZN( u0_u7_u6_n122 ) , .A1( u0_u7_u6_n94 ) , .A2( u0_u7_u6_n97 ) );
  INV_X1 u0_u7_u6_U59 (.A( u0_u7_u6_n139 ) , .ZN( u0_u7_u6_n160 ) );
  AOI22_X1 u0_u7_u6_U6 (.B2( u0_u7_u6_n101 ) , .A1( u0_u7_u6_n102 ) , .ZN( u0_u7_u6_n103 ) , .B1( u0_u7_u6_n160 ) , .A2( u0_u7_u6_n161 ) );
  NAND2_X1 u0_u7_u6_U60 (.ZN( u0_u7_u6_n113 ) , .A1( u0_u7_u6_n96 ) , .A2( u0_u7_u6_n98 ) );
  NOR2_X1 u0_u7_u6_U61 (.A2( u0_u7_X_40 ) , .A1( u0_u7_X_41 ) , .ZN( u0_u7_u6_n126 ) );
  NOR2_X1 u0_u7_u6_U62 (.A2( u0_u7_X_39 ) , .A1( u0_u7_X_42 ) , .ZN( u0_u7_u6_n92 ) );
  NOR2_X1 u0_u7_u6_U63 (.A2( u0_u7_X_39 ) , .A1( u0_u7_u6_n156 ) , .ZN( u0_u7_u6_n97 ) );
  NOR2_X1 u0_u7_u6_U64 (.A2( u0_u7_X_38 ) , .A1( u0_u7_u6_n165 ) , .ZN( u0_u7_u6_n95 ) );
  NOR2_X1 u0_u7_u6_U65 (.A2( u0_u7_X_41 ) , .ZN( u0_u7_u6_n111 ) , .A1( u0_u7_u6_n157 ) );
  NOR2_X1 u0_u7_u6_U66 (.A2( u0_u7_X_37 ) , .A1( u0_u7_u6_n162 ) , .ZN( u0_u7_u6_n94 ) );
  NOR2_X1 u0_u7_u6_U67 (.A2( u0_u7_X_37 ) , .A1( u0_u7_X_38 ) , .ZN( u0_u7_u6_n91 ) );
  NAND2_X1 u0_u7_u6_U68 (.A1( u0_u7_X_41 ) , .ZN( u0_u7_u6_n144 ) , .A2( u0_u7_u6_n157 ) );
  NAND2_X1 u0_u7_u6_U69 (.A2( u0_u7_X_40 ) , .A1( u0_u7_X_41 ) , .ZN( u0_u7_u6_n139 ) );
  NOR2_X1 u0_u7_u6_U7 (.A1( u0_u7_u6_n118 ) , .ZN( u0_u7_u6_n143 ) , .A2( u0_u7_u6_n168 ) );
  AND2_X1 u0_u7_u6_U70 (.A1( u0_u7_X_39 ) , .A2( u0_u7_u6_n156 ) , .ZN( u0_u7_u6_n96 ) );
  AND2_X1 u0_u7_u6_U71 (.A1( u0_u7_X_39 ) , .A2( u0_u7_X_42 ) , .ZN( u0_u7_u6_n99 ) );
  INV_X1 u0_u7_u6_U72 (.A( u0_u7_X_40 ) , .ZN( u0_u7_u6_n157 ) );
  INV_X1 u0_u7_u6_U73 (.A( u0_u7_X_37 ) , .ZN( u0_u7_u6_n165 ) );
  INV_X1 u0_u7_u6_U74 (.A( u0_u7_X_38 ) , .ZN( u0_u7_u6_n162 ) );
  INV_X1 u0_u7_u6_U75 (.A( u0_u7_X_42 ) , .ZN( u0_u7_u6_n156 ) );
  NAND4_X1 u0_u7_u6_U76 (.ZN( u0_out7_32 ) , .A4( u0_u7_u6_n103 ) , .A3( u0_u7_u6_n104 ) , .A2( u0_u7_u6_n105 ) , .A1( u0_u7_u6_n106 ) );
  AOI22_X1 u0_u7_u6_U77 (.ZN( u0_u7_u6_n105 ) , .A2( u0_u7_u6_n108 ) , .A1( u0_u7_u6_n118 ) , .B2( u0_u7_u6_n126 ) , .B1( u0_u7_u6_n171 ) );
  AOI22_X1 u0_u7_u6_U78 (.ZN( u0_u7_u6_n104 ) , .A1( u0_u7_u6_n111 ) , .B1( u0_u7_u6_n124 ) , .B2( u0_u7_u6_n151 ) , .A2( u0_u7_u6_n93 ) );
  NAND4_X1 u0_u7_u6_U79 (.ZN( u0_out7_12 ) , .A4( u0_u7_u6_n114 ) , .A3( u0_u7_u6_n115 ) , .A2( u0_u7_u6_n116 ) , .A1( u0_u7_u6_n117 ) );
  AOI21_X1 u0_u7_u6_U8 (.B1( u0_u7_u6_n107 ) , .B2( u0_u7_u6_n132 ) , .A( u0_u7_u6_n158 ) , .ZN( u0_u7_u6_n88 ) );
  OAI22_X1 u0_u7_u6_U80 (.B2( u0_u7_u6_n111 ) , .ZN( u0_u7_u6_n116 ) , .B1( u0_u7_u6_n126 ) , .A2( u0_u7_u6_n164 ) , .A1( u0_u7_u6_n167 ) );
  OAI21_X1 u0_u7_u6_U81 (.A( u0_u7_u6_n108 ) , .ZN( u0_u7_u6_n117 ) , .B2( u0_u7_u6_n141 ) , .B1( u0_u7_u6_n163 ) );
  OAI211_X1 u0_u7_u6_U82 (.ZN( u0_out7_22 ) , .B( u0_u7_u6_n137 ) , .A( u0_u7_u6_n138 ) , .C2( u0_u7_u6_n139 ) , .C1( u0_u7_u6_n140 ) );
  AOI22_X1 u0_u7_u6_U83 (.B1( u0_u7_u6_n124 ) , .A2( u0_u7_u6_n125 ) , .A1( u0_u7_u6_n126 ) , .ZN( u0_u7_u6_n138 ) , .B2( u0_u7_u6_n161 ) );
  AND4_X1 u0_u7_u6_U84 (.A3( u0_u7_u6_n119 ) , .A1( u0_u7_u6_n120 ) , .A4( u0_u7_u6_n129 ) , .ZN( u0_u7_u6_n140 ) , .A2( u0_u7_u6_n143 ) );
  OAI211_X1 u0_u7_u6_U85 (.ZN( u0_out7_7 ) , .B( u0_u7_u6_n153 ) , .C2( u0_u7_u6_n154 ) , .C1( u0_u7_u6_n155 ) , .A( u0_u7_u6_n174 ) );
  NOR3_X1 u0_u7_u6_U86 (.A1( u0_u7_u6_n141 ) , .ZN( u0_u7_u6_n154 ) , .A3( u0_u7_u6_n164 ) , .A2( u0_u7_u6_n171 ) );
  AOI211_X1 u0_u7_u6_U87 (.B( u0_u7_u6_n149 ) , .A( u0_u7_u6_n150 ) , .C2( u0_u7_u6_n151 ) , .C1( u0_u7_u6_n152 ) , .ZN( u0_u7_u6_n153 ) );
  NAND3_X1 u0_u7_u6_U88 (.A2( u0_u7_u6_n123 ) , .ZN( u0_u7_u6_n125 ) , .A1( u0_u7_u6_n130 ) , .A3( u0_u7_u6_n131 ) );
  NAND3_X1 u0_u7_u6_U89 (.A3( u0_u7_u6_n133 ) , .ZN( u0_u7_u6_n141 ) , .A1( u0_u7_u6_n145 ) , .A2( u0_u7_u6_n148 ) );
  AOI21_X1 u0_u7_u6_U9 (.B2( u0_u7_u6_n147 ) , .B1( u0_u7_u6_n148 ) , .ZN( u0_u7_u6_n149 ) , .A( u0_u7_u6_n158 ) );
  NAND3_X1 u0_u7_u6_U90 (.ZN( u0_u7_u6_n101 ) , .A3( u0_u7_u6_n107 ) , .A2( u0_u7_u6_n121 ) , .A1( u0_u7_u6_n127 ) );
  NAND3_X1 u0_u7_u6_U91 (.ZN( u0_u7_u6_n102 ) , .A3( u0_u7_u6_n130 ) , .A2( u0_u7_u6_n145 ) , .A1( u0_u7_u6_n166 ) );
  NAND3_X1 u0_u7_u6_U92 (.A3( u0_u7_u6_n113 ) , .A1( u0_u7_u6_n119 ) , .A2( u0_u7_u6_n123 ) , .ZN( u0_u7_u6_n93 ) );
  NAND3_X1 u0_u7_u6_U93 (.ZN( u0_u7_u6_n142 ) , .A2( u0_u7_u6_n172 ) , .A3( u0_u7_u6_n89 ) , .A1( u0_u7_u6_n90 ) );
  OAI221_X1 u0_u7_u7_U10 (.C1( u0_u7_u7_n101 ) , .C2( u0_u7_u7_n147 ) , .ZN( u0_u7_u7_n155 ) , .B2( u0_u7_u7_n162 ) , .A( u0_u7_u7_n91 ) , .B1( u0_u7_u7_n92 ) );
  AND3_X1 u0_u7_u7_U11 (.A3( u0_u7_u7_n110 ) , .A2( u0_u7_u7_n127 ) , .A1( u0_u7_u7_n132 ) , .ZN( u0_u7_u7_n92 ) );
  OAI21_X1 u0_u7_u7_U12 (.A( u0_u7_u7_n161 ) , .B1( u0_u7_u7_n168 ) , .B2( u0_u7_u7_n173 ) , .ZN( u0_u7_u7_n91 ) );
  AOI211_X1 u0_u7_u7_U13 (.A( u0_u7_u7_n117 ) , .ZN( u0_u7_u7_n118 ) , .C2( u0_u7_u7_n126 ) , .C1( u0_u7_u7_n177 ) , .B( u0_u7_u7_n180 ) );
  OAI22_X1 u0_u7_u7_U14 (.B1( u0_u7_u7_n115 ) , .ZN( u0_u7_u7_n117 ) , .A2( u0_u7_u7_n133 ) , .A1( u0_u7_u7_n137 ) , .B2( u0_u7_u7_n162 ) );
  INV_X1 u0_u7_u7_U15 (.A( u0_u7_u7_n116 ) , .ZN( u0_u7_u7_n180 ) );
  NOR3_X1 u0_u7_u7_U16 (.ZN( u0_u7_u7_n115 ) , .A3( u0_u7_u7_n145 ) , .A2( u0_u7_u7_n168 ) , .A1( u0_u7_u7_n169 ) );
  NOR3_X1 u0_u7_u7_U17 (.A2( u0_u7_u7_n134 ) , .A1( u0_u7_u7_n135 ) , .ZN( u0_u7_u7_n136 ) , .A3( u0_u7_u7_n171 ) );
  NOR2_X1 u0_u7_u7_U18 (.A1( u0_u7_u7_n130 ) , .A2( u0_u7_u7_n134 ) , .ZN( u0_u7_u7_n153 ) );
  NOR2_X1 u0_u7_u7_U19 (.ZN( u0_u7_u7_n111 ) , .A2( u0_u7_u7_n134 ) , .A1( u0_u7_u7_n169 ) );
  AOI21_X1 u0_u7_u7_U20 (.ZN( u0_u7_u7_n104 ) , .B2( u0_u7_u7_n112 ) , .B1( u0_u7_u7_n127 ) , .A( u0_u7_u7_n164 ) );
  AOI21_X1 u0_u7_u7_U21 (.ZN( u0_u7_u7_n106 ) , .B1( u0_u7_u7_n133 ) , .B2( u0_u7_u7_n146 ) , .A( u0_u7_u7_n162 ) );
  AOI21_X1 u0_u7_u7_U22 (.A( u0_u7_u7_n101 ) , .ZN( u0_u7_u7_n107 ) , .B2( u0_u7_u7_n128 ) , .B1( u0_u7_u7_n175 ) );
  INV_X1 u0_u7_u7_U23 (.A( u0_u7_u7_n101 ) , .ZN( u0_u7_u7_n165 ) );
  INV_X1 u0_u7_u7_U24 (.A( u0_u7_u7_n138 ) , .ZN( u0_u7_u7_n171 ) );
  INV_X1 u0_u7_u7_U25 (.A( u0_u7_u7_n131 ) , .ZN( u0_u7_u7_n177 ) );
  INV_X1 u0_u7_u7_U26 (.A( u0_u7_u7_n110 ) , .ZN( u0_u7_u7_n174 ) );
  NAND2_X1 u0_u7_u7_U27 (.A1( u0_u7_u7_n129 ) , .A2( u0_u7_u7_n132 ) , .ZN( u0_u7_u7_n149 ) );
  NAND2_X1 u0_u7_u7_U28 (.A1( u0_u7_u7_n113 ) , .A2( u0_u7_u7_n124 ) , .ZN( u0_u7_u7_n130 ) );
  INV_X1 u0_u7_u7_U29 (.A( u0_u7_u7_n128 ) , .ZN( u0_u7_u7_n168 ) );
  OAI21_X1 u0_u7_u7_U3 (.ZN( u0_u7_u7_n159 ) , .A( u0_u7_u7_n165 ) , .B2( u0_u7_u7_n171 ) , .B1( u0_u7_u7_n174 ) );
  INV_X1 u0_u7_u7_U30 (.A( u0_u7_u7_n148 ) , .ZN( u0_u7_u7_n169 ) );
  INV_X1 u0_u7_u7_U31 (.A( u0_u7_u7_n112 ) , .ZN( u0_u7_u7_n173 ) );
  INV_X1 u0_u7_u7_U32 (.A( u0_u7_u7_n127 ) , .ZN( u0_u7_u7_n179 ) );
  NOR2_X1 u0_u7_u7_U33 (.ZN( u0_u7_u7_n101 ) , .A2( u0_u7_u7_n150 ) , .A1( u0_u7_u7_n156 ) );
  AOI211_X1 u0_u7_u7_U34 (.B( u0_u7_u7_n154 ) , .A( u0_u7_u7_n155 ) , .C1( u0_u7_u7_n156 ) , .ZN( u0_u7_u7_n157 ) , .C2( u0_u7_u7_n172 ) );
  INV_X1 u0_u7_u7_U35 (.A( u0_u7_u7_n153 ) , .ZN( u0_u7_u7_n172 ) );
  AOI211_X1 u0_u7_u7_U36 (.B( u0_u7_u7_n139 ) , .A( u0_u7_u7_n140 ) , .C2( u0_u7_u7_n141 ) , .ZN( u0_u7_u7_n142 ) , .C1( u0_u7_u7_n156 ) );
  NAND4_X1 u0_u7_u7_U37 (.A3( u0_u7_u7_n127 ) , .A2( u0_u7_u7_n128 ) , .A1( u0_u7_u7_n129 ) , .ZN( u0_u7_u7_n141 ) , .A4( u0_u7_u7_n147 ) );
  AOI21_X1 u0_u7_u7_U38 (.A( u0_u7_u7_n137 ) , .B1( u0_u7_u7_n138 ) , .ZN( u0_u7_u7_n139 ) , .B2( u0_u7_u7_n146 ) );
  OAI22_X1 u0_u7_u7_U39 (.B1( u0_u7_u7_n136 ) , .ZN( u0_u7_u7_n140 ) , .A1( u0_u7_u7_n153 ) , .B2( u0_u7_u7_n162 ) , .A2( u0_u7_u7_n164 ) );
  INV_X1 u0_u7_u7_U4 (.A( u0_u7_u7_n149 ) , .ZN( u0_u7_u7_n175 ) );
  INV_X1 u0_u7_u7_U40 (.A( u0_u7_u7_n125 ) , .ZN( u0_u7_u7_n161 ) );
  AOI21_X1 u0_u7_u7_U41 (.ZN( u0_u7_u7_n123 ) , .B1( u0_u7_u7_n165 ) , .B2( u0_u7_u7_n177 ) , .A( u0_u7_u7_n97 ) );
  AOI21_X1 u0_u7_u7_U42 (.B2( u0_u7_u7_n113 ) , .B1( u0_u7_u7_n124 ) , .A( u0_u7_u7_n125 ) , .ZN( u0_u7_u7_n97 ) );
  INV_X1 u0_u7_u7_U43 (.A( u0_u7_u7_n152 ) , .ZN( u0_u7_u7_n162 ) );
  AOI22_X1 u0_u7_u7_U44 (.A2( u0_u7_u7_n114 ) , .ZN( u0_u7_u7_n119 ) , .B1( u0_u7_u7_n130 ) , .A1( u0_u7_u7_n156 ) , .B2( u0_u7_u7_n165 ) );
  NAND2_X1 u0_u7_u7_U45 (.A2( u0_u7_u7_n112 ) , .ZN( u0_u7_u7_n114 ) , .A1( u0_u7_u7_n175 ) );
  NOR2_X1 u0_u7_u7_U46 (.ZN( u0_u7_u7_n137 ) , .A1( u0_u7_u7_n150 ) , .A2( u0_u7_u7_n161 ) );
  AND2_X1 u0_u7_u7_U47 (.ZN( u0_u7_u7_n145 ) , .A2( u0_u7_u7_n98 ) , .A1( u0_u7_u7_n99 ) );
  AOI21_X1 u0_u7_u7_U48 (.ZN( u0_u7_u7_n105 ) , .B2( u0_u7_u7_n110 ) , .A( u0_u7_u7_n125 ) , .B1( u0_u7_u7_n147 ) );
  NAND2_X1 u0_u7_u7_U49 (.ZN( u0_u7_u7_n146 ) , .A1( u0_u7_u7_n95 ) , .A2( u0_u7_u7_n98 ) );
  INV_X1 u0_u7_u7_U5 (.A( u0_u7_u7_n154 ) , .ZN( u0_u7_u7_n178 ) );
  NAND2_X1 u0_u7_u7_U50 (.A2( u0_u7_u7_n103 ) , .ZN( u0_u7_u7_n147 ) , .A1( u0_u7_u7_n93 ) );
  NAND2_X1 u0_u7_u7_U51 (.A1( u0_u7_u7_n103 ) , .ZN( u0_u7_u7_n127 ) , .A2( u0_u7_u7_n99 ) );
  NAND2_X1 u0_u7_u7_U52 (.A2( u0_u7_u7_n102 ) , .A1( u0_u7_u7_n103 ) , .ZN( u0_u7_u7_n133 ) );
  OR2_X1 u0_u7_u7_U53 (.ZN( u0_u7_u7_n126 ) , .A2( u0_u7_u7_n152 ) , .A1( u0_u7_u7_n156 ) );
  NAND2_X1 u0_u7_u7_U54 (.ZN( u0_u7_u7_n112 ) , .A2( u0_u7_u7_n96 ) , .A1( u0_u7_u7_n99 ) );
  NAND2_X1 u0_u7_u7_U55 (.A2( u0_u7_u7_n102 ) , .ZN( u0_u7_u7_n128 ) , .A1( u0_u7_u7_n98 ) );
  INV_X1 u0_u7_u7_U56 (.A( u0_u7_u7_n150 ) , .ZN( u0_u7_u7_n164 ) );
  AND2_X1 u0_u7_u7_U57 (.ZN( u0_u7_u7_n134 ) , .A1( u0_u7_u7_n93 ) , .A2( u0_u7_u7_n98 ) );
  NAND2_X1 u0_u7_u7_U58 (.ZN( u0_u7_u7_n110 ) , .A1( u0_u7_u7_n95 ) , .A2( u0_u7_u7_n96 ) );
  NAND2_X1 u0_u7_u7_U59 (.A2( u0_u7_u7_n102 ) , .ZN( u0_u7_u7_n124 ) , .A1( u0_u7_u7_n96 ) );
  INV_X1 u0_u7_u7_U6 (.A( u0_u7_u7_n111 ) , .ZN( u0_u7_u7_n170 ) );
  NAND2_X1 u0_u7_u7_U60 (.ZN( u0_u7_u7_n132 ) , .A1( u0_u7_u7_n93 ) , .A2( u0_u7_u7_n96 ) );
  NAND2_X1 u0_u7_u7_U61 (.A2( u0_u7_u7_n103 ) , .ZN( u0_u7_u7_n131 ) , .A1( u0_u7_u7_n95 ) );
  NOR2_X1 u0_u7_u7_U62 (.A2( u0_u7_X_47 ) , .ZN( u0_u7_u7_n150 ) , .A1( u0_u7_u7_n163 ) );
  NOR2_X1 u0_u7_u7_U63 (.A2( u0_u7_X_43 ) , .A1( u0_u7_X_44 ) , .ZN( u0_u7_u7_n103 ) );
  NOR2_X1 u0_u7_u7_U64 (.A2( u0_u7_X_48 ) , .A1( u0_u7_u7_n166 ) , .ZN( u0_u7_u7_n95 ) );
  NOR2_X1 u0_u7_u7_U65 (.A2( u0_u7_X_44 ) , .A1( u0_u7_u7_n167 ) , .ZN( u0_u7_u7_n98 ) );
  NOR2_X1 u0_u7_u7_U66 (.A2( u0_u7_X_45 ) , .A1( u0_u7_X_48 ) , .ZN( u0_u7_u7_n99 ) );
  NOR2_X1 u0_u7_u7_U67 (.A2( u0_u7_X_46 ) , .A1( u0_u7_X_47 ) , .ZN( u0_u7_u7_n152 ) );
  AND2_X1 u0_u7_u7_U68 (.A1( u0_u7_X_47 ) , .ZN( u0_u7_u7_n156 ) , .A2( u0_u7_u7_n163 ) );
  NAND2_X1 u0_u7_u7_U69 (.A2( u0_u7_X_46 ) , .A1( u0_u7_X_47 ) , .ZN( u0_u7_u7_n125 ) );
  AOI211_X1 u0_u7_u7_U7 (.ZN( u0_u7_u7_n116 ) , .A( u0_u7_u7_n155 ) , .C1( u0_u7_u7_n161 ) , .C2( u0_u7_u7_n171 ) , .B( u0_u7_u7_n94 ) );
  AND2_X1 u0_u7_u7_U70 (.A2( u0_u7_X_43 ) , .A1( u0_u7_X_44 ) , .ZN( u0_u7_u7_n96 ) );
  AND2_X1 u0_u7_u7_U71 (.A2( u0_u7_X_45 ) , .A1( u0_u7_X_48 ) , .ZN( u0_u7_u7_n102 ) );
  AND2_X1 u0_u7_u7_U72 (.A1( u0_u7_X_48 ) , .A2( u0_u7_u7_n166 ) , .ZN( u0_u7_u7_n93 ) );
  INV_X1 u0_u7_u7_U73 (.A( u0_u7_X_46 ) , .ZN( u0_u7_u7_n163 ) );
  AND2_X1 u0_u7_u7_U74 (.A1( u0_u7_X_44 ) , .ZN( u0_u7_u7_n100 ) , .A2( u0_u7_u7_n167 ) );
  INV_X1 u0_u7_u7_U75 (.A( u0_u7_X_45 ) , .ZN( u0_u7_u7_n166 ) );
  INV_X1 u0_u7_u7_U76 (.A( u0_u7_X_43 ) , .ZN( u0_u7_u7_n167 ) );
  NAND4_X1 u0_u7_u7_U77 (.ZN( u0_out7_5 ) , .A4( u0_u7_u7_n108 ) , .A3( u0_u7_u7_n109 ) , .A1( u0_u7_u7_n116 ) , .A2( u0_u7_u7_n123 ) );
  AOI22_X1 u0_u7_u7_U78 (.ZN( u0_u7_u7_n109 ) , .A2( u0_u7_u7_n126 ) , .B2( u0_u7_u7_n145 ) , .B1( u0_u7_u7_n156 ) , .A1( u0_u7_u7_n171 ) );
  NOR4_X1 u0_u7_u7_U79 (.A4( u0_u7_u7_n104 ) , .A3( u0_u7_u7_n105 ) , .A2( u0_u7_u7_n106 ) , .A1( u0_u7_u7_n107 ) , .ZN( u0_u7_u7_n108 ) );
  OAI222_X1 u0_u7_u7_U8 (.C2( u0_u7_u7_n101 ) , .B2( u0_u7_u7_n111 ) , .A1( u0_u7_u7_n113 ) , .C1( u0_u7_u7_n146 ) , .A2( u0_u7_u7_n162 ) , .B1( u0_u7_u7_n164 ) , .ZN( u0_u7_u7_n94 ) );
  NAND4_X1 u0_u7_u7_U80 (.ZN( u0_out7_27 ) , .A4( u0_u7_u7_n118 ) , .A3( u0_u7_u7_n119 ) , .A2( u0_u7_u7_n120 ) , .A1( u0_u7_u7_n121 ) );
  OAI21_X1 u0_u7_u7_U81 (.ZN( u0_u7_u7_n121 ) , .B2( u0_u7_u7_n145 ) , .A( u0_u7_u7_n150 ) , .B1( u0_u7_u7_n174 ) );
  OAI21_X1 u0_u7_u7_U82 (.ZN( u0_u7_u7_n120 ) , .A( u0_u7_u7_n161 ) , .B2( u0_u7_u7_n170 ) , .B1( u0_u7_u7_n179 ) );
  NAND4_X1 u0_u7_u7_U83 (.ZN( u0_out7_21 ) , .A4( u0_u7_u7_n157 ) , .A3( u0_u7_u7_n158 ) , .A2( u0_u7_u7_n159 ) , .A1( u0_u7_u7_n160 ) );
  OAI21_X1 u0_u7_u7_U84 (.B1( u0_u7_u7_n145 ) , .ZN( u0_u7_u7_n160 ) , .A( u0_u7_u7_n161 ) , .B2( u0_u7_u7_n177 ) );
  AOI22_X1 u0_u7_u7_U85 (.B2( u0_u7_u7_n149 ) , .B1( u0_u7_u7_n150 ) , .A2( u0_u7_u7_n151 ) , .A1( u0_u7_u7_n152 ) , .ZN( u0_u7_u7_n158 ) );
  NAND4_X1 u0_u7_u7_U86 (.ZN( u0_out7_15 ) , .A4( u0_u7_u7_n142 ) , .A3( u0_u7_u7_n143 ) , .A2( u0_u7_u7_n144 ) , .A1( u0_u7_u7_n178 ) );
  OR2_X1 u0_u7_u7_U87 (.A2( u0_u7_u7_n125 ) , .A1( u0_u7_u7_n129 ) , .ZN( u0_u7_u7_n144 ) );
  AOI22_X1 u0_u7_u7_U88 (.A2( u0_u7_u7_n126 ) , .ZN( u0_u7_u7_n143 ) , .B2( u0_u7_u7_n165 ) , .B1( u0_u7_u7_n173 ) , .A1( u0_u7_u7_n174 ) );
  NAND2_X1 u0_u7_u7_U89 (.A1( u0_u7_u7_n100 ) , .ZN( u0_u7_u7_n148 ) , .A2( u0_u7_u7_n95 ) );
  INV_X1 u0_u7_u7_U9 (.A( u0_u7_u7_n133 ) , .ZN( u0_u7_u7_n176 ) );
  NAND2_X1 u0_u7_u7_U90 (.A1( u0_u7_u7_n100 ) , .ZN( u0_u7_u7_n113 ) , .A2( u0_u7_u7_n93 ) );
  NAND2_X1 u0_u7_u7_U91 (.A1( u0_u7_u7_n100 ) , .ZN( u0_u7_u7_n138 ) , .A2( u0_u7_u7_n99 ) );
  NAND2_X1 u0_u7_u7_U92 (.A1( u0_u7_u7_n100 ) , .A2( u0_u7_u7_n102 ) , .ZN( u0_u7_u7_n129 ) );
  OAI211_X1 u0_u7_u7_U93 (.B( u0_u7_u7_n122 ) , .A( u0_u7_u7_n123 ) , .C2( u0_u7_u7_n124 ) , .ZN( u0_u7_u7_n154 ) , .C1( u0_u7_u7_n162 ) );
  AOI222_X1 u0_u7_u7_U94 (.ZN( u0_u7_u7_n122 ) , .C2( u0_u7_u7_n126 ) , .C1( u0_u7_u7_n145 ) , .B1( u0_u7_u7_n161 ) , .A2( u0_u7_u7_n165 ) , .B2( u0_u7_u7_n170 ) , .A1( u0_u7_u7_n176 ) );
  NAND3_X1 u0_u7_u7_U95 (.A3( u0_u7_u7_n146 ) , .A2( u0_u7_u7_n147 ) , .A1( u0_u7_u7_n148 ) , .ZN( u0_u7_u7_n151 ) );
  NAND3_X1 u0_u7_u7_U96 (.A3( u0_u7_u7_n131 ) , .A2( u0_u7_u7_n132 ) , .A1( u0_u7_u7_n133 ) , .ZN( u0_u7_u7_n135 ) );
  OAI22_X1 u0_uk_U100 (.ZN( u0_K12_5 ) , .B2( u0_uk_n150 ) , .A2( u0_uk_n176 ) , .A1( u0_uk_n209 ) , .B1( u0_uk_n83 ) );
  OAI21_X1 u0_uk_U1002 (.ZN( u0_K8_4 ) , .B2( u0_uk_n351 ) , .A( u0_uk_n743 ) , .B1( u0_uk_n92 ) );
  NAND2_X1 u0_uk_U1003 (.A1( u0_uk_K_r6_19 ) , .A2( u0_uk_n11 ) , .ZN( u0_uk_n743 ) );
  NAND2_X1 u0_uk_U1009 (.A1( u0_key_r_46 ) , .A2( u0_uk_n60 ) , .ZN( u0_uk_n890 ) );
  NAND2_X1 u0_uk_U1011 (.A1( u0_key_r_10 ) , .A2( u0_uk_n27 ) , .ZN( u0_uk_n888 ) );
  OAI21_X1 u0_uk_U1024 (.ZN( u0_K8_46 ) , .B1( u0_uk_n250 ) , .B2( u0_uk_n326 ) , .A( u0_uk_n744 ) );
  NAND2_X1 u0_uk_U1025 (.A1( u0_uk_K_r6_37 ) , .A2( u0_uk_n203 ) , .ZN( u0_uk_n744 ) );
  OAI21_X1 u0_uk_U1032 (.ZN( u0_K8_41 ) , .B2( u0_uk_n341 ) , .B1( u0_uk_n63 ) , .A( u0_uk_n748 ) );
  OAI21_X1 u0_uk_U1054 (.ZN( u0_K8_42 ) , .B1( u0_uk_n31 ) , .B2( u0_uk_n348 ) , .A( u0_uk_n747 ) );
  NAND2_X1 u0_uk_U1055 (.A1( u0_uk_K_r6_22 ) , .A2( u0_uk_n10 ) , .ZN( u0_uk_n747 ) );
  OAI21_X1 u0_uk_U1058 (.ZN( u0_K4_38 ) , .B1( u0_uk_n27 ) , .B2( u0_uk_n505 ) , .A( u0_uk_n825 ) );
  NAND2_X1 u0_uk_U1059 (.A1( u0_uk_K_r2_50 ) , .A2( u0_uk_n63 ) , .ZN( u0_uk_n825 ) );
  OAI21_X1 u0_uk_U1087 (.ZN( u0_K8_14 ) , .B1( u0_uk_n250 ) , .B2( u0_uk_n329 ) , .A( u0_uk_n760 ) );
  NAND2_X1 u0_uk_U1088 (.A1( u0_uk_K_r6_34 ) , .A2( u0_uk_n202 ) , .ZN( u0_uk_n760 ) );
  OAI21_X1 u0_uk_U1095 (.ZN( u0_K8_39 ) , .B1( u0_uk_n191 ) , .B2( u0_uk_n332 ) , .A( u0_uk_n750 ) );
  NAND2_X1 u0_uk_U1096 (.A1( u0_uk_K_r6_31 ) , .A2( u0_uk_n208 ) , .ZN( u0_uk_n750 ) );
  INV_X1 u0_uk_U1113 (.ZN( u0_K8_12 ) , .A( u0_uk_n761 ) );
  AOI22_X1 u0_uk_U1114 (.B2( u0_uk_K_r6_3 ) , .A2( u0_uk_K_r6_53 ) , .B1( u0_uk_n142 ) , .A1( u0_uk_n162 ) , .ZN( u0_uk_n761 ) );
  INV_X1 u0_uk_U1117 (.ZN( u0_K12_4 ) , .A( u0_uk_n963 ) );
  INV_X1 u0_uk_U1145 (.ZN( u0_K8_15 ) , .A( u0_uk_n759 ) );
  INV_X1 u0_uk_U1156 (.ZN( u0_K6_2 ) , .A( u0_uk_n793 ) );
  INV_X1 u0_uk_U1158 (.ZN( u0_K8_3 ) , .A( u0_uk_n749 ) );
  AOI22_X1 u0_uk_U1160 (.B2( u0_uk_K_r10_39 ) , .A2( u0_uk_K_r10_48 ) , .B1( u0_uk_n11 ) , .A1( u0_uk_n213 ) , .ZN( u0_uk_n978 ) );
  INV_X1 u0_uk_U1161 (.ZN( u0_K12_1 ) , .A( u0_uk_n978 ) );
  OAI22_X1 u0_uk_U118 (.ZN( u0_K8_47 ) , .A1( u0_uk_n257 ) , .B1( u0_uk_n27 ) , .A2( u0_uk_n321 ) , .B2( u0_uk_n327 ) );
  OAI21_X1 u0_uk_U120 (.ZN( u0_K6_47 ) , .B1( u0_uk_n11 ) , .B2( u0_uk_n439 ) , .A( u0_uk_n789 ) );
  NAND2_X1 u0_uk_U121 (.A1( u0_uk_K_r4_23 ) , .ZN( u0_uk_n789 ) , .A2( u0_uk_n93 ) );
  OAI22_X1 u0_uk_U123 (.ZN( u0_K4_47 ) , .A1( u0_uk_n161 ) , .A2( u0_uk_n499 ) , .B2( u0_uk_n508 ) , .B1( u0_uk_n93 ) );
  INV_X1 u0_uk_U13 (.A( u0_uk_n252 ) , .ZN( u0_uk_n60 ) );
  NAND2_X1 u0_uk_U141 (.A1( u0_uk_K_r4_48 ) , .A2( u0_uk_n11 ) , .ZN( u0_uk_n798 ) );
  INV_X1 u0_uk_U159 (.ZN( u0_K2_19 ) , .A( u0_uk_n864 ) );
  AOI22_X1 u0_uk_U160 (.B2( u0_uk_K_r0_11 ) , .A2( u0_uk_K_r0_47 ) , .A1( u0_uk_n141 ) , .B1( u0_uk_n217 ) , .ZN( u0_uk_n864 ) );
  OAI21_X1 u0_uk_U173 (.ZN( u0_K8_30 ) , .B1( u0_uk_n250 ) , .B2( u0_uk_n333 ) , .A( u0_uk_n753 ) );
  NAND2_X1 u0_uk_U174 (.A1( u0_uk_K_r6_29 ) , .A2( u0_uk_n207 ) , .ZN( u0_uk_n753 ) );
  INV_X1 u0_uk_U18 (.ZN( u0_uk_n117 ) , .A( u0_uk_n182 ) );
  OAI22_X1 u0_uk_U186 (.ZN( u0_K6_14 ) , .A1( u0_uk_n102 ) , .B1( u0_uk_n164 ) , .B2( u0_uk_n442 ) , .A2( u0_uk_n448 ) );
  NAND2_X1 u0_uk_U194 (.A1( u0_uk_K_r11_28 ) , .A2( u0_uk_n11 ) , .ZN( u0_uk_n945 ) );
  NAND2_X1 u0_uk_U202 (.A1( u0_key_r_45 ) , .A2( u0_uk_n27 ) , .ZN( u0_uk_n880 ) );
  INV_X1 u0_uk_U21 (.ZN( u0_uk_n102 ) , .A( u0_uk_n162 ) );
  OAI22_X1 u0_uk_U215 (.ZN( u0_K8_31 ) , .A1( u0_uk_n102 ) , .B1( u0_uk_n223 ) , .A2( u0_uk_n321 ) , .B2( u0_uk_n359 ) );
  OAI21_X1 u0_uk_U216 (.ZN( u0_K12_31 ) , .B2( u0_uk_n173 ) , .B1( u0_uk_n250 ) , .A( u0_uk_n973 ) );
  NAND2_X1 u0_uk_U217 (.A1( u0_uk_K_r10_44 ) , .A2( u0_uk_n208 ) , .ZN( u0_uk_n973 ) );
  OAI22_X1 u0_uk_U228 (.ZN( u0_K6_31 ) , .A1( u0_uk_n182 ) , .A2( u0_uk_n428 ) , .B2( u0_uk_n433 ) , .B1( u0_uk_n60 ) );
  INV_X1 u0_uk_U24 (.ZN( u0_uk_n11 ) , .A( u0_uk_n242 ) );
  NAND2_X1 u0_uk_U240 (.A1( u0_uk_K_r10_16 ) , .A2( u0_uk_n11 ) , .ZN( u0_uk_n969 ) );
  OAI21_X1 u0_uk_U247 (.ZN( u0_K8_44 ) , .B1( u0_uk_n117 ) , .B2( u0_uk_n320 ) , .A( u0_uk_n745 ) );
  NAND2_X1 u0_uk_U248 (.A1( u0_uk_K_r6_0 ) , .A2( u0_uk_n11 ) , .ZN( u0_uk_n745 ) );
  OAI22_X1 u0_uk_U249 (.ZN( u0_K8_48 ) , .A1( u0_uk_n100 ) , .B1( u0_uk_n223 ) , .B2( u0_uk_n347 ) , .A2( u0_uk_n354 ) );
  NAND2_X1 u0_uk_U257 (.A1( u0_uk_K_r11_8 ) , .A2( u0_uk_n141 ) , .ZN( u0_uk_n942 ) );
  OAI22_X1 u0_uk_U268 (.ZN( u0_K6_44 ) , .A1( u0_uk_n109 ) , .B1( u0_uk_n231 ) , .A2( u0_uk_n412 ) , .B2( u0_uk_n430 ) );
  OAI22_X1 u0_uk_U269 (.ZN( u0_K6_48 ) , .A1( u0_uk_n242 ) , .A2( u0_uk_n418 ) , .B2( u0_uk_n425 ) , .B1( u0_uk_n60 ) );
  OAI22_X1 u0_uk_U272 (.ZN( u0_K4_44 ) , .A1( u0_uk_n141 ) , .B1( u0_uk_n202 ) , .A2( u0_uk_n521 ) , .B2( u0_uk_n538 ) );
  OAI22_X1 u0_uk_U279 (.ZN( u0_K6_6 ) , .A1( u0_uk_n162 ) , .A2( u0_uk_n410 ) , .B2( u0_uk_n414 ) , .B1( u0_uk_n60 ) );
  OAI21_X1 u0_uk_U280 (.ZN( u0_K6_8 ) , .B2( u0_uk_n442 ) , .B1( u0_uk_n63 ) , .A( u0_uk_n786 ) );
  OAI22_X1 u0_uk_U287 (.ZN( u0_K8_8 ) , .A1( u0_uk_n162 ) , .B1( u0_uk_n27 ) , .A2( u0_uk_n324 ) , .B2( u0_uk_n330 ) );
  BUF_X1 u0_uk_U29 (.Z( u0_uk_n162 ) , .A( u0_uk_n217 ) );
  OAI22_X1 u0_uk_U318 (.ZN( u0_K8_26 ) , .A1( u0_uk_n102 ) , .B1( u0_uk_n222 ) , .B2( u0_uk_n348 ) , .A2( u0_uk_n355 ) );
  OAI22_X1 u0_uk_U319 (.ZN( u0_K3_26 ) , .A1( u0_uk_n109 ) , .B1( u0_uk_n242 ) , .A2( u0_uk_n543 ) , .B2( u0_uk_n559 ) );
  OAI22_X1 u0_uk_U326 (.ZN( u0_K4_46 ) , .A1( u0_uk_n145 ) , .B1( u0_uk_n163 ) , .A2( u0_uk_n514 ) , .B2( u0_uk_n528 ) );
  INV_X1 u0_uk_U341 (.ZN( u0_K6_4 ) , .A( u0_uk_n788 ) );
  AOI22_X1 u0_uk_U342 (.B2( u0_uk_K_r4_41 ) , .A2( u0_uk_K_r4_47 ) , .A1( u0_uk_n142 ) , .B1( u0_uk_n202 ) , .ZN( u0_uk_n788 ) );
  NAND2_X1 u0_uk_U344 (.A1( u0_uk_K_r3_4 ) , .A2( u0_uk_n11 ) , .ZN( u0_uk_n804 ) );
  OAI22_X1 u0_uk_U363 (.ZN( u0_K8_40 ) , .A1( u0_uk_n162 ) , .B1( u0_uk_n27 ) , .A2( u0_uk_n327 ) , .B2( u0_uk_n333 ) );
  OAI22_X1 u0_uk_U365 (.ZN( u0_K4_40 ) , .B1( u0_uk_n145 ) , .A1( u0_uk_n182 ) , .A2( u0_uk_n506 ) , .B2( u0_uk_n516 ) );
  BUF_X1 u0_uk_U37 (.Z( u0_uk_n182 ) , .A( u0_uk_n214 ) );
  OAI22_X1 u0_uk_U378 (.ZN( u0_K3_28 ) , .A1( u0_uk_n209 ) , .A2( u0_uk_n555 ) , .B2( u0_uk_n560 ) , .B1( u0_uk_n63 ) );
  BUF_X1 u0_uk_U39 (.Z( u0_uk_n202 ) , .A( u0_uk_n208 ) );
  OAI22_X1 u0_uk_U396 (.ZN( u0_K8_16 ) , .A1( u0_uk_n213 ) , .A2( u0_uk_n344 ) , .B2( u0_uk_n352 ) , .B1( u0_uk_n63 ) );
  INV_X1 u0_uk_U4 (.ZN( u0_uk_n145 ) , .A( u0_uk_n242 ) );
  OAI22_X1 u0_uk_U409 (.ZN( u0_K8_9 ) , .A1( u0_uk_n100 ) , .B1( u0_uk_n162 ) , .B2( u0_uk_n350 ) , .A2( u0_uk_n356 ) );
  INV_X1 u0_uk_U414 (.ZN( u0_K8_37 ) , .A( u0_uk_n751 ) );
  AOI22_X1 u0_uk_U415 (.B2( u0_uk_K_r6_14 ) , .A2( u0_uk_K_r6_7 ) , .B1( u0_uk_n141 ) , .A1( u0_uk_n240 ) , .ZN( u0_uk_n751 ) );
  OAI21_X1 u0_uk_U441 (.ZN( u0_K12_33 ) , .B1( u0_uk_n10 ) , .B2( u0_uk_n140 ) , .A( u0_uk_n971 ) );
  NAND2_X1 u0_uk_U442 (.A1( u0_uk_K_r10_14 ) , .A2( u0_uk_n118 ) , .ZN( u0_uk_n971 ) );
  OAI22_X1 u0_uk_U448 (.ZN( u0_K6_33 ) , .A1( u0_uk_n213 ) , .A2( u0_uk_n425 ) , .B2( u0_uk_n430 ) , .B1( u0_uk_n60 ) );
  BUF_X1 u0_uk_U46 (.A( u0_uk_n162 ) , .Z( u0_uk_n223 ) );
  OAI22_X1 u0_uk_U463 (.ZN( u0_K4_37 ) , .A1( u0_uk_n141 ) , .B1( u0_uk_n251 ) , .A2( u0_uk_n513 ) , .B2( u0_uk_n527 ) );
  INV_X1 u0_uk_U464 (.ZN( u0_K6_9 ) , .A( u0_uk_n785 ) );
  NAND2_X1 u0_uk_U471 (.A1( u0_uk_K_r8_21 ) , .ZN( u0_uk_n1010 ) , .A2( u0_uk_n11 ) );
  OAI21_X1 u0_uk_U479 (.ZN( u0_K3_29 ) , .B1( u0_uk_n252 ) , .B2( u0_uk_n545 ) , .A( u0_uk_n849 ) );
  NAND2_X1 u0_uk_U480 (.A1( u0_uk_K_r1_44 ) , .A2( u0_uk_n220 ) , .ZN( u0_uk_n849 ) );
  OAI22_X1 u0_uk_U489 (.ZN( u0_K12_2 ) , .A1( u0_uk_n148 ) , .B2( u0_uk_n172 ) , .A2( u0_uk_n177 ) , .B1( u0_uk_n92 ) );
  OAI21_X1 u0_uk_U493 (.ZN( u0_K8_2 ) , .B2( u0_uk_n343 ) , .A( u0_uk_n754 ) , .B1( u0_uk_n83 ) );
  NAND2_X1 u0_uk_U494 (.A1( u0_uk_K_r6_27 ) , .A2( u0_uk_n11 ) , .ZN( u0_uk_n754 ) );
  INV_X1 u0_uk_U5 (.ZN( u0_uk_n141 ) , .A( u0_uk_n191 ) );
  BUF_X1 u0_uk_U50 (.A( u0_uk_n162 ) , .Z( u0_uk_n213 ) );
  INV_X1 u0_uk_U506 (.ZN( u0_K8_29 ) , .A( u0_uk_n755 ) );
  BUF_X1 u0_uk_U51 (.A( u0_uk_n161 ) , .Z( u0_uk_n242 ) );
  OAI21_X1 u0_uk_U510 (.ZN( u0_K8_17 ) , .B1( u0_uk_n252 ) , .B2( u0_uk_n336 ) , .A( u0_uk_n758 ) );
  NAND2_X1 u0_uk_U511 (.A1( u0_uk_K_r6_26 ) , .A2( u0_uk_n220 ) , .ZN( u0_uk_n758 ) );
  INV_X1 u0_uk_U542 (.ZN( u0_K6_17 ) , .A( u0_uk_n800 ) );
  AOI22_X1 u0_uk_U543 (.B2( u0_uk_K_r4_4 ) , .A2( u0_uk_K_r4_55 ) , .B1( u0_uk_n142 ) , .A1( u0_uk_n242 ) , .ZN( u0_uk_n800 ) );
  OAI22_X1 u0_uk_U581 (.ZN( u0_K8_10 ) , .A1( u0_uk_n223 ) , .B1( u0_uk_n31 ) , .A2( u0_uk_n337 ) , .B2( u0_uk_n339 ) );
  INV_X1 u0_uk_U582 (.ZN( u0_K6_10 ) , .A( u0_uk_n801 ) );
  AOI22_X1 u0_uk_U583 (.B2( u0_uk_K_r4_3 ) , .A2( u0_uk_K_r4_54 ) , .B1( u0_uk_n142 ) , .A1( u0_uk_n223 ) , .ZN( u0_uk_n801 ) );
  OAI22_X1 u0_uk_U598 (.ZN( u0_K8_22 ) , .A1( u0_uk_n257 ) , .A2( u0_uk_n323 ) , .B2( u0_uk_n329 ) , .B1( u0_uk_n92 ) );
  OAI22_X1 u0_uk_U605 (.ZN( u0_K8_35 ) , .A1( u0_uk_n242 ) , .B1( u0_uk_n31 ) , .A2( u0_uk_n341 ) , .B2( u0_uk_n347 ) );
  OAI22_X1 u0_uk_U618 (.ZN( u0_K6_35 ) , .A1( u0_uk_n242 ) , .A2( u0_uk_n412 ) , .B2( u0_uk_n419 ) , .B1( u0_uk_n60 ) );
  INV_X1 u0_uk_U62 (.ZN( u0_K8_34 ) , .A( u0_uk_n752 ) );
  AOI22_X1 u0_uk_U63 (.B2( u0_uk_K_r6_14 ) , .A2( u0_uk_K_r6_21 ) , .A1( u0_uk_n141 ) , .B1( u0_uk_n202 ) , .ZN( u0_uk_n752 ) );
  OAI21_X1 u0_uk_U645 (.ZN( u0_K12_6 ) , .B1( u0_uk_n147 ) , .B2( u0_uk_n156 ) , .A( u0_uk_n962 ) );
  NAND2_X1 u0_uk_U646 (.A1( u0_uk_K_r10_10 ) , .A2( u0_uk_n163 ) , .ZN( u0_uk_n962 ) );
  OAI21_X1 u0_uk_U68 (.ZN( u0_K6_34 ) , .B1( u0_uk_n118 ) , .B2( u0_uk_n417 ) , .A( u0_uk_n792 ) );
  NAND2_X1 u0_uk_U681 (.A1( u0_uk_K_r10_19 ) , .A2( u0_uk_n27 ) , .ZN( u0_uk_n961 ) );
  NAND2_X1 u0_uk_U69 (.A1( u0_uk_K_r4_49 ) , .ZN( u0_uk_n792 ) , .A2( u0_uk_n83 ) );
  INV_X1 u0_uk_U697 (.ZN( u0_K8_43 ) , .A( u0_uk_n746 ) );
  OAI21_X1 u0_uk_U699 (.ZN( u0_K6_7 ) , .B1( u0_uk_n252 ) , .B2( u0_uk_n423 ) , .A( u0_uk_n787 ) );
  INV_X1 u0_uk_U7 (.A( u0_uk_n147 ) , .ZN( u0_uk_n27 ) );
  NAND2_X1 u0_uk_U700 (.A1( u0_uk_K_r4_33 ) , .A2( u0_uk_n202 ) , .ZN( u0_uk_n787 ) );
  OAI22_X1 u0_uk_U701 (.ZN( u0_K8_25 ) , .A1( u0_uk_n161 ) , .A2( u0_uk_n320 ) , .B2( u0_uk_n325 ) , .B1( u0_uk_n60 ) );
  OAI22_X1 u0_uk_U718 (.ZN( u0_K8_32 ) , .A1( u0_uk_n213 ) , .B1( u0_uk_n27 ) , .A2( u0_uk_n325 ) , .B2( u0_uk_n332 ) );
  NAND2_X1 u0_uk_U72 (.A1( u0_uk_K_r1_36 ) , .A2( u0_uk_n11 ) , .ZN( u0_uk_n848 ) );
  OAI22_X1 u0_uk_U721 (.ZN( u0_K6_32 ) , .A1( u0_uk_n102 ) , .B1( u0_uk_n182 ) , .A2( u0_uk_n424 ) , .B2( u0_uk_n440 ) );
  OAI22_X1 u0_uk_U733 (.ZN( u0_K4_42 ) , .B1( u0_uk_n102 ) , .A1( u0_uk_n240 ) , .A2( u0_uk_n521 ) , .B2( u0_uk_n528 ) );
  INV_X1 u0_uk_U738 (.ZN( u0_K12_32 ) , .A( u0_uk_n972 ) );
  AOI22_X1 u0_uk_U739 (.B2( u0_uk_K_r10_23 ) , .A2( u0_uk_K_r10_28 ) , .A1( u0_uk_n251 ) , .B1( u0_uk_n60 ) , .ZN( u0_uk_n972 ) );
  NAND2_X1 u0_uk_U748 (.A1( u0_uk_K_r8_43 ) , .ZN( u0_uk_n1016 ) , .A2( u0_uk_n11 ) );
  OAI22_X1 u0_uk_U749 (.ZN( u0_K8_27 ) , .B1( u0_uk_n128 ) , .A1( u0_uk_n257 ) , .A2( u0_uk_n354 ) , .B2( u0_uk_n359 ) );
  OAI22_X1 u0_uk_U753 (.ZN( u0_K8_13 ) , .A1( u0_uk_n109 ) , .B1( u0_uk_n257 ) , .B2( u0_uk_n351 ) , .A2( u0_uk_n357 ) );
  OAI22_X1 u0_uk_U767 (.ZN( u0_K2_21 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n230 ) , .B2( u0_uk_n620 ) , .A2( u0_uk_n624 ) );
  OAI21_X1 u0_uk_U778 (.ZN( u0_K3_27 ) , .B1( u0_uk_n252 ) , .B2( u0_uk_n543 ) , .A( u0_uk_n850 ) );
  NAND2_X1 u0_uk_U779 (.A1( u0_uk_K_r1_42 ) , .A2( u0_uk_n220 ) , .ZN( u0_uk_n850 ) );
  INV_X1 u0_uk_U786 (.ZN( u0_K6_21 ) , .A( u0_uk_n797 ) );
  AOI22_X1 u0_uk_U787 (.B2( u0_uk_K_r4_11 ) , .A2( u0_uk_K_r4_5 ) , .B1( u0_uk_n142 ) , .A1( u0_uk_n220 ) , .ZN( u0_uk_n797 ) );
  OAI22_X1 u0_uk_U79 (.ZN( u0_K8_23 ) , .A1( u0_uk_n223 ) , .A2( u0_uk_n340 ) , .B2( u0_uk_n345 ) , .B1( u0_uk_n93 ) );
  OAI22_X1 u0_uk_U799 (.ZN( u0_K6_1 ) , .A1( u0_uk_n100 ) , .B1( u0_uk_n164 ) , .A2( u0_uk_n410 ) , .B2( u0_uk_n426 ) );
  OAI21_X1 u0_uk_U812 (.ZN( u0_K8_18 ) , .B2( u0_uk_n331 ) , .A( u0_uk_n757 ) , .B1( u0_uk_n93 ) );
  NAND2_X1 u0_uk_U813 (.A1( u0_uk_K_r6_46 ) , .A2( u0_uk_n10 ) , .ZN( u0_uk_n757 ) );
  OAI22_X1 u0_uk_U824 (.ZN( u0_K8_20 ) , .B1( u0_uk_n110 ) , .A1( u0_uk_n213 ) , .A2( u0_uk_n331 ) , .B2( u0_uk_n337 ) );
  INV_X1 u0_uk_U827 (.ZN( u0_K6_18 ) , .A( u0_uk_n799 ) );
  OAI22_X1 u0_uk_U83 (.ZN( u0_K2_23 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n231 ) , .A2( u0_uk_n589 ) , .B2( u0_uk_n610 ) );
  INV_X1 u0_uk_U844 (.ZN( u0_K12_3 ) , .A( u0_uk_n968 ) );
  AOI22_X1 u0_uk_U845 (.B2( u0_uk_K_r10_18 ) , .A2( u0_uk_K_r10_27 ) , .A1( u0_uk_n188 ) , .B1( u0_uk_n27 ) , .ZN( u0_uk_n968 ) );
  AOI22_X1 u0_uk_U846 (.B2( u0_uk_K_r6_10 ) , .A2( u0_uk_K_r6_3 ) , .B1( u0_uk_n141 ) , .A1( u0_uk_n161 ) , .ZN( u0_uk_n749 ) );
  OAI22_X1 u0_uk_U879 (.ZN( u0_K8_5 ) , .A1( u0_uk_n223 ) , .B1( u0_uk_n27 ) , .A2( u0_uk_n318 ) , .B2( u0_uk_n324 ) );
  OAI22_X1 u0_uk_U880 (.ZN( u0_K6_5 ) , .A1( u0_uk_n162 ) , .A2( u0_uk_n432 ) , .B2( u0_uk_n436 ) , .B1( u0_uk_n60 ) );
  OAI22_X1 u0_uk_U889 (.ZN( u0_K6_45 ) , .A1( u0_uk_n213 ) , .A2( u0_uk_n429 ) , .B2( u0_uk_n434 ) , .B1( u0_uk_n60 ) );
  OAI22_X1 u0_uk_U890 (.ZN( u0_K3_30 ) , .A1( u0_uk_n209 ) , .A2( u0_uk_n544 ) , .B2( u0_uk_n570 ) , .B1( u0_uk_n63 ) );
  OAI22_X1 u0_uk_U891 (.ZN( u0_K8_6 ) , .A1( u0_uk_n162 ) , .B1( u0_uk_n27 ) , .A2( u0_uk_n339 ) , .B2( u0_uk_n344 ) );
  OAI22_X1 u0_uk_U897 (.ZN( u0_K6_12 ) , .A1( u0_uk_n257 ) , .B2( u0_uk_n432 ) , .A2( u0_uk_n448 ) , .B1( u0_uk_n83 ) );
  OAI22_X1 u0_uk_U907 (.ZN( u0_K2_24 ) , .A1( u0_uk_n188 ) , .B2( u0_uk_n609 ) , .A2( u0_uk_n624 ) , .B1( u0_uk_n83 ) );
  OAI22_X1 u0_uk_U909 (.ZN( u0_K8_21 ) , .B1( u0_uk_n102 ) , .A1( u0_uk_n257 ) , .A2( u0_uk_n330 ) , .B2( u0_uk_n336 ) );
  OAI22_X1 u0_uk_U91 (.ZN( u0_K4_41 ) , .A1( u0_uk_n109 ) , .B1( u0_uk_n163 ) , .A2( u0_uk_n522 ) , .B2( u0_uk_n539 ) );
  OAI22_X1 u0_uk_U919 (.ZN( u0_K3_25 ) , .A1( u0_uk_n191 ) , .A2( u0_uk_n575 ) , .B2( u0_uk_n579 ) , .B1( u0_uk_n63 ) );
  OAI22_X1 u0_uk_U921 (.ZN( u0_K8_38 ) , .A1( u0_uk_n223 ) , .B1( u0_uk_n27 ) , .A2( u0_uk_n322 ) , .B2( u0_uk_n328 ) );
  OAI22_X1 u0_uk_U925 (.ZN( u0_K4_39 ) , .A1( u0_uk_n182 ) , .A2( u0_uk_n516 ) , .B2( u0_uk_n537 ) , .B1( u0_uk_n60 ) );
  OAI22_X1 u0_uk_U941 (.ZN( u0_K2_20 ) , .A1( u0_uk_n146 ) , .B1( u0_uk_n238 ) , .B2( u0_uk_n596 ) , .A2( u0_uk_n625 ) );
  OAI22_X1 u0_uk_U944 (.ZN( u0_K8_24 ) , .A1( u0_uk_n102 ) , .B1( u0_uk_n213 ) , .A2( u0_uk_n318 ) , .B2( u0_uk_n358 ) );
  OAI22_X1 u0_uk_U951 (.ZN( u0_K6_46 ) , .A1( u0_uk_n109 ) , .B1( u0_uk_n203 ) , .B2( u0_uk_n417 ) , .A2( u0_uk_n445 ) );
  OAI22_X1 u0_uk_U965 (.ZN( u0_K6_36 ) , .A1( u0_uk_n102 ) , .B1( u0_uk_n164 ) , .B2( u0_uk_n439 ) , .A2( u0_uk_n447 ) );
  OAI22_X1 u0_uk_U973 (.ZN( u0_K2_22 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n220 ) , .A2( u0_uk_n598 ) , .B2( u0_uk_n615 ) );
  OAI22_X1 u0_uk_U977 (.ZN( u0_K6_43 ) , .A1( u0_uk_n109 ) , .B1( u0_uk_n214 ) , .A2( u0_uk_n411 ) , .B2( u0_uk_n450 ) );
  OAI22_X1 u0_uk_U978 (.ZN( u0_K4_45 ) , .B1( u0_uk_n163 ) , .A1( u0_uk_n27 ) , .A2( u0_uk_n498 ) , .B2( u0_uk_n537 ) );
  OAI22_X1 u0_uk_U981 (.ZN( u0_K6_3 ) , .A1( u0_uk_n102 ) , .B1( u0_uk_n182 ) , .A2( u0_uk_n427 ) , .B2( u0_uk_n441 ) );
  OAI22_X1 u0_uk_U983 (.ZN( u0_K8_7 ) , .A1( u0_uk_n100 ) , .B1( u0_uk_n257 ) , .B2( u0_uk_n352 ) , .A2( u0_uk_n358 ) );
  OAI22_X1 u0_uk_U987 (.ZN( u0_K6_15 ) , .A1( u0_uk_n141 ) , .B1( u0_uk_n182 ) , .A2( u0_uk_n423 ) , .B2( u0_uk_n435 ) );
  NAND2_X1 u0_uk_U997 (.A1( u0_uk_K_r5_13 ) , .A2( u0_uk_n63 ) , .ZN( u0_uk_n777 ) );
  XOR2_X1 u1_U103 (.B( u1_L0_13 ) , .Z( u1_N44 ) , .A( u1_out1_13 ) );
  XOR2_X1 u1_U11 (.B( u1_L1_28 ) , .Z( u1_N91 ) , .A( u1_out2_28 ) );
  XOR2_X1 u1_U166 (.B( u1_L10_32 ) , .Z( u1_N383 ) , .A( u1_out11_32 ) );
  XOR2_X1 u1_U172 (.B( u1_L10_27 ) , .Z( u1_N378 ) , .A( u1_out11_27 ) );
  XOR2_X1 u1_U177 (.B( u1_L10_22 ) , .Z( u1_N373 ) , .A( u1_out11_22 ) );
  XOR2_X1 u1_U178 (.B( u1_L10_21 ) , .Z( u1_N372 ) , .A( u1_out11_21 ) );
  XOR2_X1 u1_U185 (.B( u1_L10_15 ) , .Z( u1_N366 ) , .A( u1_out11_15 ) );
  XOR2_X1 u1_U188 (.B( u1_L10_12 ) , .Z( u1_N363 ) , .A( u1_out11_12 ) );
  XOR2_X1 u1_U194 (.B( u1_L10_7 ) , .Z( u1_N358 ) , .A( u1_out11_7 ) );
  XOR2_X1 u1_U196 (.B( u1_L10_5 ) , .Z( u1_N356 ) , .A( u1_out11_5 ) );
  XOR2_X1 u1_U22 (.B( u1_L1_18 ) , .Z( u1_N81 ) , .A( u1_out2_18 ) );
  XOR2_X1 u1_U225 (.B( u1_L0_2 ) , .Z( u1_N33 ) , .A( u1_out1_2 ) );
  XOR2_X1 u1_U237 (.B( u1_L8_32 ) , .Z( u1_N319 ) , .A( u1_out9_32 ) );
  XOR2_X1 u1_U239 (.B( u1_L8_30 ) , .Z( u1_N317 ) , .A( u1_out9_30 ) );
  XOR2_X1 u1_U240 (.B( u1_L8_29 ) , .Z( u1_N316 ) , .A( u1_out9_29 ) );
  XOR2_X1 u1_U241 (.B( u1_L8_28 ) , .Z( u1_N315 ) , .A( u1_out9_28 ) );
  XOR2_X1 u1_U243 (.B( u1_L8_26 ) , .Z( u1_N313 ) , .A( u1_out9_26 ) );
  XOR2_X1 u1_U245 (.B( u1_L8_24 ) , .Z( u1_N311 ) , .A( u1_out9_24 ) );
  XOR2_X1 u1_U248 (.B( u1_L8_22 ) , .Z( u1_N309 ) , .A( u1_out9_22 ) );
  XOR2_X1 u1_U250 (.B( u1_L8_20 ) , .Z( u1_N307 ) , .A( u1_out9_20 ) );
  XOR2_X1 u1_U251 (.B( u1_L8_19 ) , .Z( u1_N306 ) , .A( u1_out9_19 ) );
  XOR2_X1 u1_U252 (.B( u1_L8_18 ) , .Z( u1_N305 ) , .A( u1_out9_18 ) );
  XOR2_X1 u1_U254 (.B( u1_L8_16 ) , .Z( u1_N303 ) , .A( u1_out9_16 ) );
  XOR2_X1 u1_U257 (.B( u1_L8_13 ) , .Z( u1_N300 ) , .A( u1_out9_13 ) );
  XOR2_X1 u1_U259 (.Z( u1_N3 ) , .B( u1_desIn_r_30 ) , .A( u1_out0_4 ) );
  XOR2_X1 u1_U260 (.B( u1_L8_12 ) , .Z( u1_N299 ) , .A( u1_out9_12 ) );
  XOR2_X1 u1_U261 (.B( u1_L8_11 ) , .Z( u1_N298 ) , .A( u1_out9_11 ) );
  XOR2_X1 u1_U262 (.B( u1_L8_10 ) , .Z( u1_N297 ) , .A( u1_out9_10 ) );
  XOR2_X1 u1_U265 (.B( u1_L8_7 ) , .Z( u1_N294 ) , .A( u1_out9_7 ) );
  XOR2_X1 u1_U266 (.B( u1_L8_6 ) , .Z( u1_N293 ) , .A( u1_out9_6 ) );
  XOR2_X1 u1_U268 (.B( u1_L8_4 ) , .Z( u1_N291 ) , .A( u1_out9_4 ) );
  XOR2_X1 u1_U271 (.B( u1_L8_2 ) , .Z( u1_N289 ) , .A( u1_out9_2 ) );
  XOR2_X1 u1_U272 (.B( u1_L8_1 ) , .Z( u1_N288 ) , .A( u1_out9_1 ) );
  XOR2_X1 u1_U274 (.B( u1_L7_31 ) , .Z( u1_N286 ) , .A( u1_out8_31 ) );
  XOR2_X1 u1_U28 (.B( u1_L1_13 ) , .Z( u1_N76 ) , .A( u1_out2_13 ) );
  XOR2_X1 u1_U281 (.Z( u1_N28 ) , .B( u1_desIn_r_32 ) , .A( u1_out0_29 ) );
  XOR2_X1 u1_U283 (.B( u1_L7_23 ) , .Z( u1_N278 ) , .A( u1_out8_23 ) );
  XOR2_X1 u1_U289 (.B( u1_L7_17 ) , .Z( u1_N272 ) , .A( u1_out8_17 ) );
  XOR2_X1 u1_U298 (.B( u1_L7_9 ) , .Z( u1_N264 ) , .A( u1_out8_9 ) );
  XOR2_X1 u1_U313 (.B( u1_L6_27 ) , .Z( u1_N250 ) , .A( u1_out7_27 ) );
  XOR2_X1 u1_U320 (.B( u1_L6_21 ) , .Z( u1_N244 ) , .A( u1_out7_21 ) );
  XOR2_X1 u1_U325 (.Z( u1_N24 ) , .B( u1_desIn_r_0 ) , .A( u1_out0_25 ) );
  XOR2_X1 u1_U327 (.B( u1_L6_15 ) , .Z( u1_N238 ) , .A( u1_out7_15 ) );
  XOR2_X1 u1_U338 (.B( u1_L6_5 ) , .Z( u1_N228 ) , .A( u1_out7_5 ) );
  XOR2_X1 u1_U348 (.B( u1_L5_28 ) , .Z( u1_N219 ) , .A( u1_out6_28 ) );
  XOR2_X1 u1_U349 (.B( u1_L5_27 ) , .Z( u1_N218 ) , .A( u1_out6_27 ) );
  XOR2_X1 u1_U35 (.Z( u1_N7 ) , .B( u1_desIn_r_62 ) , .A( u1_out0_8 ) );
  XOR2_X1 u1_U355 (.B( u1_L5_21 ) , .Z( u1_N212 ) , .A( u1_out6_21 ) );
  XOR2_X1 u1_U359 (.B( u1_L5_18 ) , .Z( u1_N209 ) , .A( u1_out6_18 ) );
  XOR2_X1 u1_U362 (.B( u1_L5_15 ) , .Z( u1_N206 ) , .A( u1_out6_15 ) );
  XOR2_X1 u1_U364 (.B( u1_L5_13 ) , .Z( u1_N204 ) , .A( u1_out6_13 ) );
  XOR2_X1 u1_U370 (.Z( u1_N2 ) , .B( u1_desIn_r_22 ) , .A( u1_out0_3 ) );
  XOR2_X1 u1_U374 (.B( u1_L5_5 ) , .Z( u1_N196 ) , .A( u1_out6_5 ) );
  XOR2_X1 u1_U377 (.B( u1_L5_2 ) , .Z( u1_N193 ) , .A( u1_out6_2 ) );
  XOR2_X1 u1_U385 (.B( u1_L4_27 ) , .Z( u1_N186 ) , .A( u1_out5_27 ) );
  XOR2_X1 u1_U391 (.B( u1_L4_21 ) , .Z( u1_N180 ) , .A( u1_out5_21 ) );
  XOR2_X1 u1_U392 (.Z( u1_N18 ) , .B( u1_desIn_r_18 ) , .A( u1_out0_19 ) );
  XOR2_X1 u1_U398 (.B( u1_L4_15 ) , .Z( u1_N174 ) , .A( u1_out5_15 ) );
  XOR2_X1 u1_U40 (.B( u1_L1_2 ) , .Z( u1_N65 ) , .A( u1_out2_2 ) );
  XOR2_X1 u1_U409 (.B( u1_L4_5 ) , .Z( u1_N164 ) , .A( u1_out5_5 ) );
  XOR2_X1 u1_U447 (.Z( u1_N13 ) , .B( u1_desIn_r_44 ) , .A( u1_out0_14 ) );
  XOR2_X1 u1_U450 (.B( u1_L2_32 ) , .Z( u1_N127 ) , .A( u1_out3_32 ) );
  XOR2_X1 u1_U454 (.B( u1_L2_28 ) , .Z( u1_N123 ) , .A( u1_out3_28 ) );
  XOR2_X1 u1_U461 (.B( u1_L2_22 ) , .Z( u1_N117 ) , .A( u1_out3_22 ) );
  XOR2_X1 u1_U465 (.B( u1_L2_18 ) , .Z( u1_N113 ) , .A( u1_out3_18 ) );
  XOR2_X1 u1_U47 (.B( u1_L0_28 ) , .Z( u1_N59 ) , .A( u1_out1_28 ) );
  XOR2_X1 u1_U471 (.B( u1_L2_13 ) , .Z( u1_N108 ) , .A( u1_out3_13 ) );
  XOR2_X1 u1_U472 (.B( u1_L2_12 ) , .Z( u1_N107 ) , .A( u1_out3_12 ) );
  XOR2_X1 u1_U477 (.B( u1_L2_7 ) , .Z( u1_N102 ) , .A( u1_out3_7 ) );
  XOR2_X1 u1_U480 (.Z( u1_N10 ) , .B( u1_desIn_r_20 ) , .A( u1_out0_11 ) );
  XOR2_X1 u1_U486 (.Z( u1_FP_6 ) , .B( u1_L14_6 ) , .A( u1_out15_6 ) );
  XOR2_X1 u1_U488 (.Z( u1_FP_4 ) , .B( u1_L14_4 ) , .A( u1_out15_4 ) );
  XOR2_X1 u1_U492 (.Z( u1_FP_30 ) , .B( u1_L14_30 ) , .A( u1_out15_30 ) );
  XOR2_X1 u1_U494 (.Z( u1_FP_29 ) , .B( u1_L14_29 ) , .A( u1_out15_29 ) );
  XOR2_X1 u1_U499 (.Z( u1_FP_24 ) , .B( u1_L14_24 ) , .A( u1_out15_24 ) );
  XOR2_X1 u1_U5 (.B( u1_L2_2 ) , .Z( u1_N97 ) , .A( u1_out3_2 ) );
  XOR2_X1 u1_U505 (.Z( u1_FP_19 ) , .B( u1_L14_19 ) , .A( u1_out15_19 ) );
  XOR2_X1 u1_U508 (.Z( u1_FP_16 ) , .B( u1_L14_16 ) , .A( u1_out15_16 ) );
  XOR2_X1 u1_U513 (.Z( u1_FP_11 ) , .B( u1_L14_11 ) , .A( u1_out15_11 ) );
  XOR2_X1 u1_U58 (.B( u1_L0_18 ) , .Z( u1_N49 ) , .A( u1_out1_18 ) );
  XOR2_X1 u1_U66 (.B( u1_L13_26 ) , .Z( u1_N473 ) , .A( u1_out14_26 ) );
  XOR2_X1 u1_U73 (.B( u1_L13_20 ) , .Z( u1_N467 ) , .A( u1_out14_20 ) );
  XOR2_X1 u1_U84 (.B( u1_L13_10 ) , .Z( u1_N457 ) , .A( u1_out14_10 ) );
  XOR2_X1 u1_U94 (.B( u1_L13_1 ) , .Z( u1_N448 ) , .A( u1_out14_1 ) );
  XOR2_X1 u1_u0_U22 (.B( u1_K1_34 ) , .A( u1_desIn_r_51 ) , .Z( u1_u0_X_34 ) );
  XOR2_X1 u1_u0_U23 (.B( u1_K1_33 ) , .A( u1_desIn_r_43 ) , .Z( u1_u0_X_33 ) );
  XOR2_X1 u1_u0_U25 (.B( u1_K1_31 ) , .A( u1_desIn_r_27 ) , .Z( u1_u0_X_31 ) );
  XOR2_X1 u1_u0_U28 (.B( u1_K1_29 ) , .A( u1_desIn_r_27 ) , .Z( u1_u0_X_29 ) );
  XOR2_X1 u1_u0_U29 (.B( u1_K1_28 ) , .A( u1_desIn_r_19 ) , .Z( u1_u0_X_28 ) );
  XOR2_X1 u1_u0_U30 (.B( u1_K1_27 ) , .A( u1_desIn_r_11 ) , .Z( u1_u0_X_27 ) );
  OAI22_X1 u1_u0_u4_U10 (.B2( u1_u0_u4_n135 ) , .ZN( u1_u0_u4_n137 ) , .B1( u1_u0_u4_n153 ) , .A1( u1_u0_u4_n155 ) , .A2( u1_u0_u4_n171 ) );
  AND3_X1 u1_u0_u4_U11 (.A2( u1_u0_u4_n134 ) , .ZN( u1_u0_u4_n135 ) , .A3( u1_u0_u4_n145 ) , .A1( u1_u0_u4_n157 ) );
  NAND2_X1 u1_u0_u4_U12 (.ZN( u1_u0_u4_n132 ) , .A2( u1_u0_u4_n170 ) , .A1( u1_u0_u4_n173 ) );
  AOI21_X1 u1_u0_u4_U13 (.B2( u1_u0_u4_n160 ) , .B1( u1_u0_u4_n161 ) , .ZN( u1_u0_u4_n162 ) , .A( u1_u0_u4_n170 ) );
  AOI21_X1 u1_u0_u4_U14 (.ZN( u1_u0_u4_n107 ) , .B2( u1_u0_u4_n143 ) , .A( u1_u0_u4_n174 ) , .B1( u1_u0_u4_n184 ) );
  AOI21_X1 u1_u0_u4_U15 (.B2( u1_u0_u4_n158 ) , .B1( u1_u0_u4_n159 ) , .ZN( u1_u0_u4_n163 ) , .A( u1_u0_u4_n174 ) );
  AOI21_X1 u1_u0_u4_U16 (.A( u1_u0_u4_n153 ) , .B2( u1_u0_u4_n154 ) , .B1( u1_u0_u4_n155 ) , .ZN( u1_u0_u4_n165 ) );
  AOI21_X1 u1_u0_u4_U17 (.A( u1_u0_u4_n156 ) , .B2( u1_u0_u4_n157 ) , .ZN( u1_u0_u4_n164 ) , .B1( u1_u0_u4_n184 ) );
  INV_X1 u1_u0_u4_U18 (.A( u1_u0_u4_n138 ) , .ZN( u1_u0_u4_n170 ) );
  AND2_X1 u1_u0_u4_U19 (.A2( u1_u0_u4_n120 ) , .ZN( u1_u0_u4_n155 ) , .A1( u1_u0_u4_n160 ) );
  INV_X1 u1_u0_u4_U20 (.A( u1_u0_u4_n156 ) , .ZN( u1_u0_u4_n175 ) );
  NAND2_X1 u1_u0_u4_U21 (.A2( u1_u0_u4_n118 ) , .ZN( u1_u0_u4_n131 ) , .A1( u1_u0_u4_n147 ) );
  NAND2_X1 u1_u0_u4_U22 (.A1( u1_u0_u4_n119 ) , .A2( u1_u0_u4_n120 ) , .ZN( u1_u0_u4_n130 ) );
  NAND2_X1 u1_u0_u4_U23 (.ZN( u1_u0_u4_n117 ) , .A2( u1_u0_u4_n118 ) , .A1( u1_u0_u4_n148 ) );
  NAND2_X1 u1_u0_u4_U24 (.ZN( u1_u0_u4_n129 ) , .A1( u1_u0_u4_n134 ) , .A2( u1_u0_u4_n148 ) );
  AND3_X1 u1_u0_u4_U25 (.A1( u1_u0_u4_n119 ) , .A2( u1_u0_u4_n143 ) , .A3( u1_u0_u4_n154 ) , .ZN( u1_u0_u4_n161 ) );
  AND2_X1 u1_u0_u4_U26 (.A1( u1_u0_u4_n145 ) , .A2( u1_u0_u4_n147 ) , .ZN( u1_u0_u4_n159 ) );
  OR3_X1 u1_u0_u4_U27 (.A3( u1_u0_u4_n114 ) , .A2( u1_u0_u4_n115 ) , .A1( u1_u0_u4_n116 ) , .ZN( u1_u0_u4_n136 ) );
  AOI21_X1 u1_u0_u4_U28 (.A( u1_u0_u4_n113 ) , .ZN( u1_u0_u4_n116 ) , .B2( u1_u0_u4_n173 ) , .B1( u1_u0_u4_n174 ) );
  AOI21_X1 u1_u0_u4_U29 (.ZN( u1_u0_u4_n115 ) , .B2( u1_u0_u4_n145 ) , .B1( u1_u0_u4_n146 ) , .A( u1_u0_u4_n156 ) );
  NOR2_X1 u1_u0_u4_U3 (.ZN( u1_u0_u4_n121 ) , .A1( u1_u0_u4_n181 ) , .A2( u1_u0_u4_n182 ) );
  OAI22_X1 u1_u0_u4_U30 (.ZN( u1_u0_u4_n114 ) , .A2( u1_u0_u4_n121 ) , .B1( u1_u0_u4_n160 ) , .B2( u1_u0_u4_n170 ) , .A1( u1_u0_u4_n171 ) );
  INV_X1 u1_u0_u4_U31 (.A( u1_u0_u4_n158 ) , .ZN( u1_u0_u4_n182 ) );
  INV_X1 u1_u0_u4_U32 (.ZN( u1_u0_u4_n181 ) , .A( u1_u0_u4_n96 ) );
  INV_X1 u1_u0_u4_U33 (.A( u1_u0_u4_n144 ) , .ZN( u1_u0_u4_n179 ) );
  INV_X1 u1_u0_u4_U34 (.A( u1_u0_u4_n157 ) , .ZN( u1_u0_u4_n178 ) );
  NAND2_X1 u1_u0_u4_U35 (.A2( u1_u0_u4_n154 ) , .A1( u1_u0_u4_n96 ) , .ZN( u1_u0_u4_n97 ) );
  INV_X1 u1_u0_u4_U36 (.ZN( u1_u0_u4_n186 ) , .A( u1_u0_u4_n95 ) );
  OAI221_X1 u1_u0_u4_U37 (.C1( u1_u0_u4_n134 ) , .B1( u1_u0_u4_n158 ) , .B2( u1_u0_u4_n171 ) , .C2( u1_u0_u4_n173 ) , .A( u1_u0_u4_n94 ) , .ZN( u1_u0_u4_n95 ) );
  AOI222_X1 u1_u0_u4_U38 (.B2( u1_u0_u4_n132 ) , .A1( u1_u0_u4_n138 ) , .C2( u1_u0_u4_n175 ) , .A2( u1_u0_u4_n179 ) , .C1( u1_u0_u4_n181 ) , .B1( u1_u0_u4_n185 ) , .ZN( u1_u0_u4_n94 ) );
  INV_X1 u1_u0_u4_U39 (.A( u1_u0_u4_n113 ) , .ZN( u1_u0_u4_n185 ) );
  INV_X1 u1_u0_u4_U4 (.A( u1_u0_u4_n117 ) , .ZN( u1_u0_u4_n184 ) );
  INV_X1 u1_u0_u4_U40 (.A( u1_u0_u4_n143 ) , .ZN( u1_u0_u4_n183 ) );
  NOR2_X1 u1_u0_u4_U41 (.ZN( u1_u0_u4_n138 ) , .A1( u1_u0_u4_n168 ) , .A2( u1_u0_u4_n169 ) );
  NOR2_X1 u1_u0_u4_U42 (.A1( u1_u0_u4_n150 ) , .A2( u1_u0_u4_n152 ) , .ZN( u1_u0_u4_n153 ) );
  NOR2_X1 u1_u0_u4_U43 (.A2( u1_u0_u4_n128 ) , .A1( u1_u0_u4_n138 ) , .ZN( u1_u0_u4_n156 ) );
  AOI22_X1 u1_u0_u4_U44 (.B2( u1_u0_u4_n122 ) , .A1( u1_u0_u4_n123 ) , .ZN( u1_u0_u4_n124 ) , .B1( u1_u0_u4_n128 ) , .A2( u1_u0_u4_n172 ) );
  INV_X1 u1_u0_u4_U45 (.A( u1_u0_u4_n153 ) , .ZN( u1_u0_u4_n172 ) );
  NAND2_X1 u1_u0_u4_U46 (.A2( u1_u0_u4_n120 ) , .ZN( u1_u0_u4_n123 ) , .A1( u1_u0_u4_n161 ) );
  AOI22_X1 u1_u0_u4_U47 (.B2( u1_u0_u4_n132 ) , .A2( u1_u0_u4_n133 ) , .ZN( u1_u0_u4_n140 ) , .A1( u1_u0_u4_n150 ) , .B1( u1_u0_u4_n179 ) );
  NAND2_X1 u1_u0_u4_U48 (.ZN( u1_u0_u4_n133 ) , .A2( u1_u0_u4_n146 ) , .A1( u1_u0_u4_n154 ) );
  NAND2_X1 u1_u0_u4_U49 (.A1( u1_u0_u4_n103 ) , .ZN( u1_u0_u4_n154 ) , .A2( u1_u0_u4_n98 ) );
  NOR4_X1 u1_u0_u4_U5 (.A4( u1_u0_u4_n106 ) , .A3( u1_u0_u4_n107 ) , .A2( u1_u0_u4_n108 ) , .A1( u1_u0_u4_n109 ) , .ZN( u1_u0_u4_n110 ) );
  NAND2_X1 u1_u0_u4_U50 (.A1( u1_u0_u4_n101 ) , .ZN( u1_u0_u4_n158 ) , .A2( u1_u0_u4_n99 ) );
  AOI21_X1 u1_u0_u4_U51 (.ZN( u1_u0_u4_n127 ) , .A( u1_u0_u4_n136 ) , .B2( u1_u0_u4_n150 ) , .B1( u1_u0_u4_n180 ) );
  INV_X1 u1_u0_u4_U52 (.A( u1_u0_u4_n160 ) , .ZN( u1_u0_u4_n180 ) );
  NAND2_X1 u1_u0_u4_U53 (.A2( u1_u0_u4_n104 ) , .A1( u1_u0_u4_n105 ) , .ZN( u1_u0_u4_n146 ) );
  NAND2_X1 u1_u0_u4_U54 (.A2( u1_u0_u4_n101 ) , .A1( u1_u0_u4_n102 ) , .ZN( u1_u0_u4_n160 ) );
  NAND2_X1 u1_u0_u4_U55 (.ZN( u1_u0_u4_n134 ) , .A1( u1_u0_u4_n98 ) , .A2( u1_u0_u4_n99 ) );
  NAND2_X1 u1_u0_u4_U56 (.A1( u1_u0_u4_n103 ) , .A2( u1_u0_u4_n104 ) , .ZN( u1_u0_u4_n143 ) );
  NAND2_X1 u1_u0_u4_U57 (.A2( u1_u0_u4_n105 ) , .ZN( u1_u0_u4_n145 ) , .A1( u1_u0_u4_n98 ) );
  NAND2_X1 u1_u0_u4_U58 (.A1( u1_u0_u4_n100 ) , .A2( u1_u0_u4_n105 ) , .ZN( u1_u0_u4_n120 ) );
  NAND2_X1 u1_u0_u4_U59 (.A1( u1_u0_u4_n102 ) , .A2( u1_u0_u4_n104 ) , .ZN( u1_u0_u4_n148 ) );
  AOI21_X1 u1_u0_u4_U6 (.ZN( u1_u0_u4_n106 ) , .B2( u1_u0_u4_n146 ) , .B1( u1_u0_u4_n158 ) , .A( u1_u0_u4_n170 ) );
  NAND2_X1 u1_u0_u4_U60 (.A2( u1_u0_u4_n100 ) , .A1( u1_u0_u4_n103 ) , .ZN( u1_u0_u4_n157 ) );
  INV_X1 u1_u0_u4_U61 (.A( u1_u0_u4_n150 ) , .ZN( u1_u0_u4_n173 ) );
  INV_X1 u1_u0_u4_U62 (.A( u1_u0_u4_n152 ) , .ZN( u1_u0_u4_n171 ) );
  NAND2_X1 u1_u0_u4_U63 (.A1( u1_u0_u4_n100 ) , .ZN( u1_u0_u4_n118 ) , .A2( u1_u0_u4_n99 ) );
  NAND2_X1 u1_u0_u4_U64 (.A2( u1_u0_u4_n100 ) , .A1( u1_u0_u4_n102 ) , .ZN( u1_u0_u4_n144 ) );
  NAND2_X1 u1_u0_u4_U65 (.A2( u1_u0_u4_n101 ) , .A1( u1_u0_u4_n105 ) , .ZN( u1_u0_u4_n96 ) );
  INV_X1 u1_u0_u4_U66 (.A( u1_u0_u4_n128 ) , .ZN( u1_u0_u4_n174 ) );
  NAND2_X1 u1_u0_u4_U67 (.A2( u1_u0_u4_n102 ) , .ZN( u1_u0_u4_n119 ) , .A1( u1_u0_u4_n98 ) );
  NAND2_X1 u1_u0_u4_U68 (.A2( u1_u0_u4_n101 ) , .A1( u1_u0_u4_n103 ) , .ZN( u1_u0_u4_n147 ) );
  NAND2_X1 u1_u0_u4_U69 (.A2( u1_u0_u4_n104 ) , .ZN( u1_u0_u4_n113 ) , .A1( u1_u0_u4_n99 ) );
  AOI21_X1 u1_u0_u4_U7 (.ZN( u1_u0_u4_n108 ) , .B2( u1_u0_u4_n134 ) , .B1( u1_u0_u4_n155 ) , .A( u1_u0_u4_n156 ) );
  NOR2_X1 u1_u0_u4_U70 (.A2( u1_u0_X_28 ) , .ZN( u1_u0_u4_n150 ) , .A1( u1_u0_u4_n168 ) );
  NOR2_X1 u1_u0_u4_U71 (.A2( u1_u0_X_29 ) , .ZN( u1_u0_u4_n152 ) , .A1( u1_u0_u4_n169 ) );
  NOR2_X1 u1_u0_u4_U72 (.A2( u1_u0_X_30 ) , .ZN( u1_u0_u4_n105 ) , .A1( u1_u0_u4_n176 ) );
  NOR2_X1 u1_u0_u4_U73 (.A2( u1_u0_X_26 ) , .ZN( u1_u0_u4_n100 ) , .A1( u1_u0_u4_n177 ) );
  NOR2_X1 u1_u0_u4_U74 (.A2( u1_u0_X_28 ) , .A1( u1_u0_X_29 ) , .ZN( u1_u0_u4_n128 ) );
  NOR2_X1 u1_u0_u4_U75 (.A2( u1_u0_X_27 ) , .A1( u1_u0_X_30 ) , .ZN( u1_u0_u4_n102 ) );
  NOR2_X1 u1_u0_u4_U76 (.A2( u1_u0_X_25 ) , .A1( u1_u0_X_26 ) , .ZN( u1_u0_u4_n98 ) );
  AND2_X1 u1_u0_u4_U77 (.A2( u1_u0_X_25 ) , .A1( u1_u0_X_26 ) , .ZN( u1_u0_u4_n104 ) );
  AND2_X1 u1_u0_u4_U78 (.A1( u1_u0_X_30 ) , .A2( u1_u0_u4_n176 ) , .ZN( u1_u0_u4_n99 ) );
  AND2_X1 u1_u0_u4_U79 (.A1( u1_u0_X_26 ) , .ZN( u1_u0_u4_n101 ) , .A2( u1_u0_u4_n177 ) );
  AOI21_X1 u1_u0_u4_U8 (.ZN( u1_u0_u4_n109 ) , .A( u1_u0_u4_n153 ) , .B1( u1_u0_u4_n159 ) , .B2( u1_u0_u4_n184 ) );
  AND2_X1 u1_u0_u4_U80 (.A1( u1_u0_X_27 ) , .A2( u1_u0_X_30 ) , .ZN( u1_u0_u4_n103 ) );
  INV_X1 u1_u0_u4_U81 (.A( u1_u0_X_28 ) , .ZN( u1_u0_u4_n169 ) );
  INV_X1 u1_u0_u4_U82 (.A( u1_u0_X_29 ) , .ZN( u1_u0_u4_n168 ) );
  INV_X1 u1_u0_u4_U83 (.A( u1_u0_X_25 ) , .ZN( u1_u0_u4_n177 ) );
  INV_X1 u1_u0_u4_U84 (.A( u1_u0_X_27 ) , .ZN( u1_u0_u4_n176 ) );
  NAND4_X1 u1_u0_u4_U85 (.ZN( u1_out0_25 ) , .A4( u1_u0_u4_n139 ) , .A3( u1_u0_u4_n140 ) , .A2( u1_u0_u4_n141 ) , .A1( u1_u0_u4_n142 ) );
  OAI21_X1 u1_u0_u4_U86 (.A( u1_u0_u4_n128 ) , .B2( u1_u0_u4_n129 ) , .B1( u1_u0_u4_n130 ) , .ZN( u1_u0_u4_n142 ) );
  OAI21_X1 u1_u0_u4_U87 (.B2( u1_u0_u4_n131 ) , .ZN( u1_u0_u4_n141 ) , .A( u1_u0_u4_n175 ) , .B1( u1_u0_u4_n183 ) );
  NAND4_X1 u1_u0_u4_U88 (.ZN( u1_out0_14 ) , .A4( u1_u0_u4_n124 ) , .A3( u1_u0_u4_n125 ) , .A2( u1_u0_u4_n126 ) , .A1( u1_u0_u4_n127 ) );
  AOI22_X1 u1_u0_u4_U89 (.B2( u1_u0_u4_n117 ) , .ZN( u1_u0_u4_n126 ) , .A1( u1_u0_u4_n129 ) , .B1( u1_u0_u4_n152 ) , .A2( u1_u0_u4_n175 ) );
  AOI211_X1 u1_u0_u4_U9 (.B( u1_u0_u4_n136 ) , .A( u1_u0_u4_n137 ) , .C2( u1_u0_u4_n138 ) , .ZN( u1_u0_u4_n139 ) , .C1( u1_u0_u4_n182 ) );
  AOI22_X1 u1_u0_u4_U90 (.ZN( u1_u0_u4_n125 ) , .B2( u1_u0_u4_n131 ) , .A2( u1_u0_u4_n132 ) , .B1( u1_u0_u4_n138 ) , .A1( u1_u0_u4_n178 ) );
  NAND4_X1 u1_u0_u4_U91 (.ZN( u1_out0_8 ) , .A4( u1_u0_u4_n110 ) , .A3( u1_u0_u4_n111 ) , .A2( u1_u0_u4_n112 ) , .A1( u1_u0_u4_n186 ) );
  NAND2_X1 u1_u0_u4_U92 (.ZN( u1_u0_u4_n112 ) , .A2( u1_u0_u4_n130 ) , .A1( u1_u0_u4_n150 ) );
  AOI22_X1 u1_u0_u4_U93 (.ZN( u1_u0_u4_n111 ) , .B2( u1_u0_u4_n132 ) , .A1( u1_u0_u4_n152 ) , .B1( u1_u0_u4_n178 ) , .A2( u1_u0_u4_n97 ) );
  AOI22_X1 u1_u0_u4_U94 (.B2( u1_u0_u4_n149 ) , .B1( u1_u0_u4_n150 ) , .A2( u1_u0_u4_n151 ) , .A1( u1_u0_u4_n152 ) , .ZN( u1_u0_u4_n167 ) );
  NOR4_X1 u1_u0_u4_U95 (.A4( u1_u0_u4_n162 ) , .A3( u1_u0_u4_n163 ) , .A2( u1_u0_u4_n164 ) , .A1( u1_u0_u4_n165 ) , .ZN( u1_u0_u4_n166 ) );
  NAND3_X1 u1_u0_u4_U96 (.ZN( u1_out0_3 ) , .A3( u1_u0_u4_n166 ) , .A1( u1_u0_u4_n167 ) , .A2( u1_u0_u4_n186 ) );
  NAND3_X1 u1_u0_u4_U97 (.A3( u1_u0_u4_n146 ) , .A2( u1_u0_u4_n147 ) , .A1( u1_u0_u4_n148 ) , .ZN( u1_u0_u4_n149 ) );
  NAND3_X1 u1_u0_u4_U98 (.A3( u1_u0_u4_n143 ) , .A2( u1_u0_u4_n144 ) , .A1( u1_u0_u4_n145 ) , .ZN( u1_u0_u4_n151 ) );
  NAND3_X1 u1_u0_u4_U99 (.A3( u1_u0_u4_n121 ) , .ZN( u1_u0_u4_n122 ) , .A2( u1_u0_u4_n144 ) , .A1( u1_u0_u4_n154 ) );
  INV_X1 u1_u0_u5_U10 (.A( u1_u0_u5_n121 ) , .ZN( u1_u0_u5_n177 ) );
  NOR3_X1 u1_u0_u5_U100 (.A3( u1_u0_u5_n141 ) , .A1( u1_u0_u5_n142 ) , .ZN( u1_u0_u5_n143 ) , .A2( u1_u0_u5_n191 ) );
  NAND4_X1 u1_u0_u5_U101 (.ZN( u1_out0_4 ) , .A4( u1_u0_u5_n112 ) , .A2( u1_u0_u5_n113 ) , .A1( u1_u0_u5_n114 ) , .A3( u1_u0_u5_n195 ) );
  AOI211_X1 u1_u0_u5_U102 (.A( u1_u0_u5_n110 ) , .C1( u1_u0_u5_n111 ) , .ZN( u1_u0_u5_n112 ) , .B( u1_u0_u5_n118 ) , .C2( u1_u0_u5_n177 ) );
  AOI222_X1 u1_u0_u5_U103 (.ZN( u1_u0_u5_n113 ) , .A1( u1_u0_u5_n131 ) , .C1( u1_u0_u5_n148 ) , .B2( u1_u0_u5_n174 ) , .C2( u1_u0_u5_n178 ) , .A2( u1_u0_u5_n179 ) , .B1( u1_u0_u5_n99 ) );
  NAND3_X1 u1_u0_u5_U104 (.A2( u1_u0_u5_n154 ) , .A3( u1_u0_u5_n158 ) , .A1( u1_u0_u5_n161 ) , .ZN( u1_u0_u5_n99 ) );
  NOR2_X1 u1_u0_u5_U11 (.ZN( u1_u0_u5_n160 ) , .A2( u1_u0_u5_n173 ) , .A1( u1_u0_u5_n177 ) );
  INV_X1 u1_u0_u5_U12 (.A( u1_u0_u5_n150 ) , .ZN( u1_u0_u5_n174 ) );
  AOI21_X1 u1_u0_u5_U13 (.A( u1_u0_u5_n160 ) , .B2( u1_u0_u5_n161 ) , .ZN( u1_u0_u5_n162 ) , .B1( u1_u0_u5_n192 ) );
  INV_X1 u1_u0_u5_U14 (.A( u1_u0_u5_n159 ) , .ZN( u1_u0_u5_n192 ) );
  AOI21_X1 u1_u0_u5_U15 (.A( u1_u0_u5_n156 ) , .B2( u1_u0_u5_n157 ) , .B1( u1_u0_u5_n158 ) , .ZN( u1_u0_u5_n163 ) );
  AOI21_X1 u1_u0_u5_U16 (.B2( u1_u0_u5_n139 ) , .B1( u1_u0_u5_n140 ) , .ZN( u1_u0_u5_n141 ) , .A( u1_u0_u5_n150 ) );
  OAI21_X1 u1_u0_u5_U17 (.A( u1_u0_u5_n133 ) , .B2( u1_u0_u5_n134 ) , .B1( u1_u0_u5_n135 ) , .ZN( u1_u0_u5_n142 ) );
  OAI21_X1 u1_u0_u5_U18 (.ZN( u1_u0_u5_n133 ) , .B2( u1_u0_u5_n147 ) , .A( u1_u0_u5_n173 ) , .B1( u1_u0_u5_n188 ) );
  NAND2_X1 u1_u0_u5_U19 (.A2( u1_u0_u5_n119 ) , .A1( u1_u0_u5_n123 ) , .ZN( u1_u0_u5_n137 ) );
  INV_X1 u1_u0_u5_U20 (.A( u1_u0_u5_n155 ) , .ZN( u1_u0_u5_n194 ) );
  NAND2_X1 u1_u0_u5_U21 (.A1( u1_u0_u5_n121 ) , .ZN( u1_u0_u5_n132 ) , .A2( u1_u0_u5_n172 ) );
  NAND2_X1 u1_u0_u5_U22 (.A2( u1_u0_u5_n122 ) , .ZN( u1_u0_u5_n136 ) , .A1( u1_u0_u5_n154 ) );
  NAND2_X1 u1_u0_u5_U23 (.A2( u1_u0_u5_n119 ) , .A1( u1_u0_u5_n120 ) , .ZN( u1_u0_u5_n159 ) );
  INV_X1 u1_u0_u5_U24 (.A( u1_u0_u5_n156 ) , .ZN( u1_u0_u5_n175 ) );
  INV_X1 u1_u0_u5_U25 (.A( u1_u0_u5_n158 ) , .ZN( u1_u0_u5_n188 ) );
  INV_X1 u1_u0_u5_U26 (.A( u1_u0_u5_n152 ) , .ZN( u1_u0_u5_n179 ) );
  INV_X1 u1_u0_u5_U27 (.A( u1_u0_u5_n140 ) , .ZN( u1_u0_u5_n182 ) );
  INV_X1 u1_u0_u5_U28 (.A( u1_u0_u5_n151 ) , .ZN( u1_u0_u5_n183 ) );
  INV_X1 u1_u0_u5_U29 (.A( u1_u0_u5_n123 ) , .ZN( u1_u0_u5_n185 ) );
  NOR2_X1 u1_u0_u5_U3 (.ZN( u1_u0_u5_n134 ) , .A1( u1_u0_u5_n183 ) , .A2( u1_u0_u5_n190 ) );
  INV_X1 u1_u0_u5_U30 (.A( u1_u0_u5_n161 ) , .ZN( u1_u0_u5_n184 ) );
  INV_X1 u1_u0_u5_U31 (.A( u1_u0_u5_n139 ) , .ZN( u1_u0_u5_n189 ) );
  INV_X1 u1_u0_u5_U32 (.A( u1_u0_u5_n157 ) , .ZN( u1_u0_u5_n190 ) );
  INV_X1 u1_u0_u5_U33 (.A( u1_u0_u5_n120 ) , .ZN( u1_u0_u5_n193 ) );
  NAND2_X1 u1_u0_u5_U34 (.ZN( u1_u0_u5_n111 ) , .A1( u1_u0_u5_n140 ) , .A2( u1_u0_u5_n155 ) );
  INV_X1 u1_u0_u5_U35 (.A( u1_u0_u5_n117 ) , .ZN( u1_u0_u5_n196 ) );
  OAI221_X1 u1_u0_u5_U36 (.A( u1_u0_u5_n116 ) , .ZN( u1_u0_u5_n117 ) , .B2( u1_u0_u5_n119 ) , .C1( u1_u0_u5_n153 ) , .C2( u1_u0_u5_n158 ) , .B1( u1_u0_u5_n172 ) );
  AOI222_X1 u1_u0_u5_U37 (.ZN( u1_u0_u5_n116 ) , .B2( u1_u0_u5_n145 ) , .C1( u1_u0_u5_n148 ) , .A2( u1_u0_u5_n174 ) , .C2( u1_u0_u5_n177 ) , .B1( u1_u0_u5_n187 ) , .A1( u1_u0_u5_n193 ) );
  INV_X1 u1_u0_u5_U38 (.A( u1_u0_u5_n115 ) , .ZN( u1_u0_u5_n187 ) );
  NOR2_X1 u1_u0_u5_U39 (.ZN( u1_u0_u5_n100 ) , .A1( u1_u0_u5_n170 ) , .A2( u1_u0_u5_n180 ) );
  INV_X1 u1_u0_u5_U4 (.A( u1_u0_u5_n138 ) , .ZN( u1_u0_u5_n191 ) );
  AOI22_X1 u1_u0_u5_U40 (.B2( u1_u0_u5_n131 ) , .A2( u1_u0_u5_n146 ) , .ZN( u1_u0_u5_n169 ) , .B1( u1_u0_u5_n174 ) , .A1( u1_u0_u5_n185 ) );
  NOR2_X1 u1_u0_u5_U41 (.A1( u1_u0_u5_n146 ) , .ZN( u1_u0_u5_n150 ) , .A2( u1_u0_u5_n173 ) );
  AOI21_X1 u1_u0_u5_U42 (.A( u1_u0_u5_n118 ) , .B2( u1_u0_u5_n145 ) , .ZN( u1_u0_u5_n168 ) , .B1( u1_u0_u5_n186 ) );
  INV_X1 u1_u0_u5_U43 (.A( u1_u0_u5_n122 ) , .ZN( u1_u0_u5_n186 ) );
  NOR2_X1 u1_u0_u5_U44 (.A1( u1_u0_u5_n146 ) , .ZN( u1_u0_u5_n152 ) , .A2( u1_u0_u5_n176 ) );
  NOR2_X1 u1_u0_u5_U45 (.A1( u1_u0_u5_n115 ) , .ZN( u1_u0_u5_n118 ) , .A2( u1_u0_u5_n153 ) );
  NOR2_X1 u1_u0_u5_U46 (.A2( u1_u0_u5_n145 ) , .ZN( u1_u0_u5_n156 ) , .A1( u1_u0_u5_n174 ) );
  NOR2_X1 u1_u0_u5_U47 (.ZN( u1_u0_u5_n121 ) , .A2( u1_u0_u5_n145 ) , .A1( u1_u0_u5_n176 ) );
  AOI22_X1 u1_u0_u5_U48 (.ZN( u1_u0_u5_n114 ) , .A2( u1_u0_u5_n137 ) , .A1( u1_u0_u5_n145 ) , .B2( u1_u0_u5_n175 ) , .B1( u1_u0_u5_n193 ) );
  OAI211_X1 u1_u0_u5_U49 (.B( u1_u0_u5_n124 ) , .A( u1_u0_u5_n125 ) , .C2( u1_u0_u5_n126 ) , .C1( u1_u0_u5_n127 ) , .ZN( u1_u0_u5_n128 ) );
  OAI21_X1 u1_u0_u5_U5 (.B2( u1_u0_u5_n136 ) , .B1( u1_u0_u5_n137 ) , .ZN( u1_u0_u5_n138 ) , .A( u1_u0_u5_n177 ) );
  NOR3_X1 u1_u0_u5_U50 (.ZN( u1_u0_u5_n127 ) , .A1( u1_u0_u5_n136 ) , .A3( u1_u0_u5_n148 ) , .A2( u1_u0_u5_n182 ) );
  OAI21_X1 u1_u0_u5_U51 (.ZN( u1_u0_u5_n124 ) , .A( u1_u0_u5_n177 ) , .B2( u1_u0_u5_n183 ) , .B1( u1_u0_u5_n189 ) );
  OAI21_X1 u1_u0_u5_U52 (.ZN( u1_u0_u5_n125 ) , .A( u1_u0_u5_n174 ) , .B2( u1_u0_u5_n185 ) , .B1( u1_u0_u5_n190 ) );
  AOI21_X1 u1_u0_u5_U53 (.A( u1_u0_u5_n153 ) , .B2( u1_u0_u5_n154 ) , .B1( u1_u0_u5_n155 ) , .ZN( u1_u0_u5_n164 ) );
  AOI21_X1 u1_u0_u5_U54 (.ZN( u1_u0_u5_n110 ) , .B1( u1_u0_u5_n122 ) , .B2( u1_u0_u5_n139 ) , .A( u1_u0_u5_n153 ) );
  INV_X1 u1_u0_u5_U55 (.A( u1_u0_u5_n153 ) , .ZN( u1_u0_u5_n176 ) );
  INV_X1 u1_u0_u5_U56 (.A( u1_u0_u5_n126 ) , .ZN( u1_u0_u5_n173 ) );
  AND2_X1 u1_u0_u5_U57 (.A2( u1_u0_u5_n104 ) , .A1( u1_u0_u5_n107 ) , .ZN( u1_u0_u5_n147 ) );
  AND2_X1 u1_u0_u5_U58 (.A2( u1_u0_u5_n104 ) , .A1( u1_u0_u5_n108 ) , .ZN( u1_u0_u5_n148 ) );
  NAND2_X1 u1_u0_u5_U59 (.A1( u1_u0_u5_n105 ) , .A2( u1_u0_u5_n106 ) , .ZN( u1_u0_u5_n158 ) );
  INV_X1 u1_u0_u5_U6 (.A( u1_u0_u5_n135 ) , .ZN( u1_u0_u5_n178 ) );
  NAND2_X1 u1_u0_u5_U60 (.A2( u1_u0_u5_n108 ) , .A1( u1_u0_u5_n109 ) , .ZN( u1_u0_u5_n139 ) );
  NAND2_X1 u1_u0_u5_U61 (.A1( u1_u0_u5_n106 ) , .A2( u1_u0_u5_n108 ) , .ZN( u1_u0_u5_n119 ) );
  NAND2_X1 u1_u0_u5_U62 (.A2( u1_u0_u5_n103 ) , .A1( u1_u0_u5_n105 ) , .ZN( u1_u0_u5_n140 ) );
  NAND2_X1 u1_u0_u5_U63 (.A2( u1_u0_u5_n104 ) , .A1( u1_u0_u5_n105 ) , .ZN( u1_u0_u5_n155 ) );
  NAND2_X1 u1_u0_u5_U64 (.A2( u1_u0_u5_n106 ) , .A1( u1_u0_u5_n107 ) , .ZN( u1_u0_u5_n122 ) );
  NAND2_X1 u1_u0_u5_U65 (.A2( u1_u0_u5_n100 ) , .A1( u1_u0_u5_n106 ) , .ZN( u1_u0_u5_n115 ) );
  NAND2_X1 u1_u0_u5_U66 (.A2( u1_u0_u5_n100 ) , .A1( u1_u0_u5_n103 ) , .ZN( u1_u0_u5_n161 ) );
  NAND2_X1 u1_u0_u5_U67 (.A1( u1_u0_u5_n105 ) , .A2( u1_u0_u5_n109 ) , .ZN( u1_u0_u5_n154 ) );
  INV_X1 u1_u0_u5_U68 (.A( u1_u0_u5_n146 ) , .ZN( u1_u0_u5_n172 ) );
  NAND2_X1 u1_u0_u5_U69 (.A1( u1_u0_u5_n103 ) , .A2( u1_u0_u5_n108 ) , .ZN( u1_u0_u5_n123 ) );
  OAI22_X1 u1_u0_u5_U7 (.B2( u1_u0_u5_n149 ) , .B1( u1_u0_u5_n150 ) , .A2( u1_u0_u5_n151 ) , .A1( u1_u0_u5_n152 ) , .ZN( u1_u0_u5_n165 ) );
  NAND2_X1 u1_u0_u5_U70 (.A2( u1_u0_u5_n103 ) , .A1( u1_u0_u5_n107 ) , .ZN( u1_u0_u5_n151 ) );
  NAND2_X1 u1_u0_u5_U71 (.A2( u1_u0_u5_n107 ) , .A1( u1_u0_u5_n109 ) , .ZN( u1_u0_u5_n120 ) );
  NAND2_X1 u1_u0_u5_U72 (.A2( u1_u0_u5_n100 ) , .A1( u1_u0_u5_n109 ) , .ZN( u1_u0_u5_n157 ) );
  AND2_X1 u1_u0_u5_U73 (.A2( u1_u0_u5_n100 ) , .A1( u1_u0_u5_n104 ) , .ZN( u1_u0_u5_n131 ) );
  INV_X1 u1_u0_u5_U74 (.A( u1_u0_u5_n102 ) , .ZN( u1_u0_u5_n195 ) );
  OAI221_X1 u1_u0_u5_U75 (.A( u1_u0_u5_n101 ) , .ZN( u1_u0_u5_n102 ) , .C2( u1_u0_u5_n115 ) , .C1( u1_u0_u5_n126 ) , .B1( u1_u0_u5_n134 ) , .B2( u1_u0_u5_n160 ) );
  OAI21_X1 u1_u0_u5_U76 (.ZN( u1_u0_u5_n101 ) , .B1( u1_u0_u5_n137 ) , .A( u1_u0_u5_n146 ) , .B2( u1_u0_u5_n147 ) );
  NOR2_X1 u1_u0_u5_U77 (.A2( u1_u0_X_34 ) , .A1( u1_u0_X_35 ) , .ZN( u1_u0_u5_n145 ) );
  NOR2_X1 u1_u0_u5_U78 (.A2( u1_u0_X_34 ) , .ZN( u1_u0_u5_n146 ) , .A1( u1_u0_u5_n171 ) );
  NOR2_X1 u1_u0_u5_U79 (.A2( u1_u0_X_31 ) , .A1( u1_u0_X_32 ) , .ZN( u1_u0_u5_n103 ) );
  NOR3_X1 u1_u0_u5_U8 (.A2( u1_u0_u5_n147 ) , .A1( u1_u0_u5_n148 ) , .ZN( u1_u0_u5_n149 ) , .A3( u1_u0_u5_n194 ) );
  NOR2_X1 u1_u0_u5_U80 (.A2( u1_u0_X_36 ) , .ZN( u1_u0_u5_n105 ) , .A1( u1_u0_u5_n180 ) );
  NOR2_X1 u1_u0_u5_U81 (.A2( u1_u0_X_33 ) , .ZN( u1_u0_u5_n108 ) , .A1( u1_u0_u5_n170 ) );
  NOR2_X1 u1_u0_u5_U82 (.A2( u1_u0_X_33 ) , .A1( u1_u0_X_36 ) , .ZN( u1_u0_u5_n107 ) );
  NOR2_X1 u1_u0_u5_U83 (.A2( u1_u0_X_31 ) , .ZN( u1_u0_u5_n104 ) , .A1( u1_u0_u5_n181 ) );
  NAND2_X1 u1_u0_u5_U84 (.A2( u1_u0_X_34 ) , .A1( u1_u0_X_35 ) , .ZN( u1_u0_u5_n153 ) );
  NAND2_X1 u1_u0_u5_U85 (.A1( u1_u0_X_34 ) , .ZN( u1_u0_u5_n126 ) , .A2( u1_u0_u5_n171 ) );
  AND2_X1 u1_u0_u5_U86 (.A1( u1_u0_X_31 ) , .A2( u1_u0_X_32 ) , .ZN( u1_u0_u5_n106 ) );
  AND2_X1 u1_u0_u5_U87 (.A1( u1_u0_X_31 ) , .ZN( u1_u0_u5_n109 ) , .A2( u1_u0_u5_n181 ) );
  INV_X1 u1_u0_u5_U88 (.A( u1_u0_X_33 ) , .ZN( u1_u0_u5_n180 ) );
  INV_X1 u1_u0_u5_U89 (.A( u1_u0_X_35 ) , .ZN( u1_u0_u5_n171 ) );
  NOR2_X1 u1_u0_u5_U9 (.ZN( u1_u0_u5_n135 ) , .A1( u1_u0_u5_n173 ) , .A2( u1_u0_u5_n176 ) );
  INV_X1 u1_u0_u5_U90 (.A( u1_u0_X_36 ) , .ZN( u1_u0_u5_n170 ) );
  INV_X1 u1_u0_u5_U91 (.A( u1_u0_X_32 ) , .ZN( u1_u0_u5_n181 ) );
  NAND4_X1 u1_u0_u5_U92 (.ZN( u1_out0_29 ) , .A4( u1_u0_u5_n129 ) , .A3( u1_u0_u5_n130 ) , .A2( u1_u0_u5_n168 ) , .A1( u1_u0_u5_n196 ) );
  AOI221_X1 u1_u0_u5_U93 (.A( u1_u0_u5_n128 ) , .ZN( u1_u0_u5_n129 ) , .C2( u1_u0_u5_n132 ) , .B2( u1_u0_u5_n159 ) , .B1( u1_u0_u5_n176 ) , .C1( u1_u0_u5_n184 ) );
  AOI222_X1 u1_u0_u5_U94 (.ZN( u1_u0_u5_n130 ) , .A2( u1_u0_u5_n146 ) , .B1( u1_u0_u5_n147 ) , .C2( u1_u0_u5_n175 ) , .B2( u1_u0_u5_n179 ) , .A1( u1_u0_u5_n188 ) , .C1( u1_u0_u5_n194 ) );
  NAND4_X1 u1_u0_u5_U95 (.ZN( u1_out0_19 ) , .A4( u1_u0_u5_n166 ) , .A3( u1_u0_u5_n167 ) , .A2( u1_u0_u5_n168 ) , .A1( u1_u0_u5_n169 ) );
  AOI22_X1 u1_u0_u5_U96 (.B2( u1_u0_u5_n145 ) , .A2( u1_u0_u5_n146 ) , .ZN( u1_u0_u5_n167 ) , .B1( u1_u0_u5_n182 ) , .A1( u1_u0_u5_n189 ) );
  NOR4_X1 u1_u0_u5_U97 (.A4( u1_u0_u5_n162 ) , .A3( u1_u0_u5_n163 ) , .A2( u1_u0_u5_n164 ) , .A1( u1_u0_u5_n165 ) , .ZN( u1_u0_u5_n166 ) );
  NAND4_X1 u1_u0_u5_U98 (.ZN( u1_out0_11 ) , .A4( u1_u0_u5_n143 ) , .A3( u1_u0_u5_n144 ) , .A2( u1_u0_u5_n169 ) , .A1( u1_u0_u5_n196 ) );
  AOI22_X1 u1_u0_u5_U99 (.A2( u1_u0_u5_n132 ) , .ZN( u1_u0_u5_n144 ) , .B2( u1_u0_u5_n145 ) , .B1( u1_u0_u5_n184 ) , .A1( u1_u0_u5_n194 ) );
  XOR2_X1 u1_u11_U10 (.B( u1_K12_45 ) , .A( u1_R10_30 ) , .Z( u1_u11_X_45 ) );
  XOR2_X1 u1_u11_U15 (.B( u1_K12_40 ) , .A( u1_R10_27 ) , .Z( u1_u11_X_40 ) );
  XOR2_X1 u1_u11_U17 (.B( u1_K12_39 ) , .A( u1_R10_26 ) , .Z( u1_u11_X_39 ) );
  XOR2_X1 u1_u11_U9 (.B( u1_K12_46 ) , .A( u1_R10_31 ) , .Z( u1_u11_X_46 ) );
  OAI21_X1 u1_u11_u6_U10 (.A( u1_u11_u6_n159 ) , .B1( u1_u11_u6_n169 ) , .B2( u1_u11_u6_n173 ) , .ZN( u1_u11_u6_n90 ) );
  INV_X1 u1_u11_u6_U11 (.ZN( u1_u11_u6_n172 ) , .A( u1_u11_u6_n88 ) );
  AOI22_X1 u1_u11_u6_U12 (.A2( u1_u11_u6_n151 ) , .B2( u1_u11_u6_n161 ) , .A1( u1_u11_u6_n167 ) , .B1( u1_u11_u6_n170 ) , .ZN( u1_u11_u6_n89 ) );
  AOI21_X1 u1_u11_u6_U13 (.ZN( u1_u11_u6_n106 ) , .A( u1_u11_u6_n142 ) , .B2( u1_u11_u6_n159 ) , .B1( u1_u11_u6_n164 ) );
  INV_X1 u1_u11_u6_U14 (.A( u1_u11_u6_n155 ) , .ZN( u1_u11_u6_n161 ) );
  INV_X1 u1_u11_u6_U15 (.A( u1_u11_u6_n128 ) , .ZN( u1_u11_u6_n164 ) );
  NAND2_X1 u1_u11_u6_U16 (.ZN( u1_u11_u6_n110 ) , .A1( u1_u11_u6_n122 ) , .A2( u1_u11_u6_n129 ) );
  NAND2_X1 u1_u11_u6_U17 (.ZN( u1_u11_u6_n124 ) , .A2( u1_u11_u6_n146 ) , .A1( u1_u11_u6_n148 ) );
  INV_X1 u1_u11_u6_U18 (.A( u1_u11_u6_n132 ) , .ZN( u1_u11_u6_n171 ) );
  AND2_X1 u1_u11_u6_U19 (.A1( u1_u11_u6_n100 ) , .ZN( u1_u11_u6_n130 ) , .A2( u1_u11_u6_n147 ) );
  INV_X1 u1_u11_u6_U20 (.A( u1_u11_u6_n127 ) , .ZN( u1_u11_u6_n173 ) );
  INV_X1 u1_u11_u6_U21 (.A( u1_u11_u6_n121 ) , .ZN( u1_u11_u6_n167 ) );
  INV_X1 u1_u11_u6_U22 (.A( u1_u11_u6_n100 ) , .ZN( u1_u11_u6_n169 ) );
  INV_X1 u1_u11_u6_U23 (.A( u1_u11_u6_n123 ) , .ZN( u1_u11_u6_n170 ) );
  INV_X1 u1_u11_u6_U24 (.A( u1_u11_u6_n113 ) , .ZN( u1_u11_u6_n168 ) );
  AND2_X1 u1_u11_u6_U25 (.A1( u1_u11_u6_n107 ) , .A2( u1_u11_u6_n119 ) , .ZN( u1_u11_u6_n133 ) );
  AND2_X1 u1_u11_u6_U26 (.A2( u1_u11_u6_n121 ) , .A1( u1_u11_u6_n122 ) , .ZN( u1_u11_u6_n131 ) );
  AND3_X1 u1_u11_u6_U27 (.ZN( u1_u11_u6_n120 ) , .A2( u1_u11_u6_n127 ) , .A1( u1_u11_u6_n132 ) , .A3( u1_u11_u6_n145 ) );
  INV_X1 u1_u11_u6_U28 (.A( u1_u11_u6_n146 ) , .ZN( u1_u11_u6_n163 ) );
  AOI222_X1 u1_u11_u6_U29 (.ZN( u1_u11_u6_n114 ) , .A1( u1_u11_u6_n118 ) , .A2( u1_u11_u6_n126 ) , .B2( u1_u11_u6_n151 ) , .C2( u1_u11_u6_n159 ) , .C1( u1_u11_u6_n168 ) , .B1( u1_u11_u6_n169 ) );
  INV_X1 u1_u11_u6_U3 (.A( u1_u11_u6_n110 ) , .ZN( u1_u11_u6_n166 ) );
  NOR2_X1 u1_u11_u6_U30 (.A1( u1_u11_u6_n162 ) , .A2( u1_u11_u6_n165 ) , .ZN( u1_u11_u6_n98 ) );
  NAND2_X1 u1_u11_u6_U31 (.A1( u1_u11_u6_n144 ) , .ZN( u1_u11_u6_n151 ) , .A2( u1_u11_u6_n158 ) );
  NAND2_X1 u1_u11_u6_U32 (.ZN( u1_u11_u6_n132 ) , .A1( u1_u11_u6_n91 ) , .A2( u1_u11_u6_n97 ) );
  AOI22_X1 u1_u11_u6_U33 (.B2( u1_u11_u6_n110 ) , .B1( u1_u11_u6_n111 ) , .A1( u1_u11_u6_n112 ) , .ZN( u1_u11_u6_n115 ) , .A2( u1_u11_u6_n161 ) );
  NAND4_X1 u1_u11_u6_U34 (.A3( u1_u11_u6_n109 ) , .ZN( u1_u11_u6_n112 ) , .A4( u1_u11_u6_n132 ) , .A2( u1_u11_u6_n147 ) , .A1( u1_u11_u6_n166 ) );
  NOR2_X1 u1_u11_u6_U35 (.ZN( u1_u11_u6_n109 ) , .A1( u1_u11_u6_n170 ) , .A2( u1_u11_u6_n173 ) );
  NOR2_X1 u1_u11_u6_U36 (.A2( u1_u11_u6_n126 ) , .ZN( u1_u11_u6_n155 ) , .A1( u1_u11_u6_n160 ) );
  NAND2_X1 u1_u11_u6_U37 (.ZN( u1_u11_u6_n146 ) , .A2( u1_u11_u6_n94 ) , .A1( u1_u11_u6_n99 ) );
  AOI21_X1 u1_u11_u6_U38 (.A( u1_u11_u6_n144 ) , .B2( u1_u11_u6_n145 ) , .B1( u1_u11_u6_n146 ) , .ZN( u1_u11_u6_n150 ) );
  AOI211_X1 u1_u11_u6_U39 (.B( u1_u11_u6_n134 ) , .A( u1_u11_u6_n135 ) , .C1( u1_u11_u6_n136 ) , .ZN( u1_u11_u6_n137 ) , .C2( u1_u11_u6_n151 ) );
  INV_X1 u1_u11_u6_U4 (.A( u1_u11_u6_n142 ) , .ZN( u1_u11_u6_n174 ) );
  NAND4_X1 u1_u11_u6_U40 (.A4( u1_u11_u6_n127 ) , .A3( u1_u11_u6_n128 ) , .A2( u1_u11_u6_n129 ) , .A1( u1_u11_u6_n130 ) , .ZN( u1_u11_u6_n136 ) );
  AOI21_X1 u1_u11_u6_U41 (.B2( u1_u11_u6_n132 ) , .B1( u1_u11_u6_n133 ) , .ZN( u1_u11_u6_n134 ) , .A( u1_u11_u6_n158 ) );
  AOI21_X1 u1_u11_u6_U42 (.B1( u1_u11_u6_n131 ) , .ZN( u1_u11_u6_n135 ) , .A( u1_u11_u6_n144 ) , .B2( u1_u11_u6_n146 ) );
  INV_X1 u1_u11_u6_U43 (.A( u1_u11_u6_n111 ) , .ZN( u1_u11_u6_n158 ) );
  NAND2_X1 u1_u11_u6_U44 (.ZN( u1_u11_u6_n127 ) , .A1( u1_u11_u6_n91 ) , .A2( u1_u11_u6_n92 ) );
  NAND2_X1 u1_u11_u6_U45 (.ZN( u1_u11_u6_n129 ) , .A2( u1_u11_u6_n95 ) , .A1( u1_u11_u6_n96 ) );
  INV_X1 u1_u11_u6_U46 (.A( u1_u11_u6_n144 ) , .ZN( u1_u11_u6_n159 ) );
  NAND2_X1 u1_u11_u6_U47 (.ZN( u1_u11_u6_n145 ) , .A2( u1_u11_u6_n97 ) , .A1( u1_u11_u6_n98 ) );
  NAND2_X1 u1_u11_u6_U48 (.ZN( u1_u11_u6_n148 ) , .A2( u1_u11_u6_n92 ) , .A1( u1_u11_u6_n94 ) );
  NAND2_X1 u1_u11_u6_U49 (.ZN( u1_u11_u6_n108 ) , .A2( u1_u11_u6_n139 ) , .A1( u1_u11_u6_n144 ) );
  NAND2_X1 u1_u11_u6_U5 (.A2( u1_u11_u6_n143 ) , .ZN( u1_u11_u6_n152 ) , .A1( u1_u11_u6_n166 ) );
  NAND2_X1 u1_u11_u6_U50 (.ZN( u1_u11_u6_n121 ) , .A2( u1_u11_u6_n95 ) , .A1( u1_u11_u6_n97 ) );
  NAND2_X1 u1_u11_u6_U51 (.ZN( u1_u11_u6_n107 ) , .A2( u1_u11_u6_n92 ) , .A1( u1_u11_u6_n95 ) );
  AND2_X1 u1_u11_u6_U52 (.ZN( u1_u11_u6_n118 ) , .A2( u1_u11_u6_n91 ) , .A1( u1_u11_u6_n99 ) );
  NAND2_X1 u1_u11_u6_U53 (.ZN( u1_u11_u6_n147 ) , .A2( u1_u11_u6_n98 ) , .A1( u1_u11_u6_n99 ) );
  NAND2_X1 u1_u11_u6_U54 (.ZN( u1_u11_u6_n128 ) , .A1( u1_u11_u6_n94 ) , .A2( u1_u11_u6_n96 ) );
  NAND2_X1 u1_u11_u6_U55 (.ZN( u1_u11_u6_n119 ) , .A2( u1_u11_u6_n95 ) , .A1( u1_u11_u6_n99 ) );
  NAND2_X1 u1_u11_u6_U56 (.ZN( u1_u11_u6_n123 ) , .A2( u1_u11_u6_n91 ) , .A1( u1_u11_u6_n96 ) );
  NAND2_X1 u1_u11_u6_U57 (.ZN( u1_u11_u6_n100 ) , .A2( u1_u11_u6_n92 ) , .A1( u1_u11_u6_n98 ) );
  NAND2_X1 u1_u11_u6_U58 (.ZN( u1_u11_u6_n122 ) , .A1( u1_u11_u6_n94 ) , .A2( u1_u11_u6_n97 ) );
  INV_X1 u1_u11_u6_U59 (.A( u1_u11_u6_n139 ) , .ZN( u1_u11_u6_n160 ) );
  AOI22_X1 u1_u11_u6_U6 (.B2( u1_u11_u6_n101 ) , .A1( u1_u11_u6_n102 ) , .ZN( u1_u11_u6_n103 ) , .B1( u1_u11_u6_n160 ) , .A2( u1_u11_u6_n161 ) );
  NAND2_X1 u1_u11_u6_U60 (.ZN( u1_u11_u6_n113 ) , .A1( u1_u11_u6_n96 ) , .A2( u1_u11_u6_n98 ) );
  NOR2_X1 u1_u11_u6_U61 (.A2( u1_u11_X_40 ) , .A1( u1_u11_X_41 ) , .ZN( u1_u11_u6_n126 ) );
  NOR2_X1 u1_u11_u6_U62 (.A2( u1_u11_X_39 ) , .A1( u1_u11_X_42 ) , .ZN( u1_u11_u6_n92 ) );
  NOR2_X1 u1_u11_u6_U63 (.A2( u1_u11_X_39 ) , .A1( u1_u11_u6_n156 ) , .ZN( u1_u11_u6_n97 ) );
  NOR2_X1 u1_u11_u6_U64 (.A2( u1_u11_X_38 ) , .A1( u1_u11_u6_n165 ) , .ZN( u1_u11_u6_n95 ) );
  NOR2_X1 u1_u11_u6_U65 (.A2( u1_u11_X_41 ) , .ZN( u1_u11_u6_n111 ) , .A1( u1_u11_u6_n157 ) );
  NOR2_X1 u1_u11_u6_U66 (.A2( u1_u11_X_37 ) , .A1( u1_u11_u6_n162 ) , .ZN( u1_u11_u6_n94 ) );
  NOR2_X1 u1_u11_u6_U67 (.A2( u1_u11_X_37 ) , .A1( u1_u11_X_38 ) , .ZN( u1_u11_u6_n91 ) );
  NAND2_X1 u1_u11_u6_U68 (.A1( u1_u11_X_41 ) , .ZN( u1_u11_u6_n144 ) , .A2( u1_u11_u6_n157 ) );
  NAND2_X1 u1_u11_u6_U69 (.A2( u1_u11_X_40 ) , .A1( u1_u11_X_41 ) , .ZN( u1_u11_u6_n139 ) );
  NOR2_X1 u1_u11_u6_U7 (.A1( u1_u11_u6_n118 ) , .ZN( u1_u11_u6_n143 ) , .A2( u1_u11_u6_n168 ) );
  AND2_X1 u1_u11_u6_U70 (.A1( u1_u11_X_39 ) , .A2( u1_u11_u6_n156 ) , .ZN( u1_u11_u6_n96 ) );
  AND2_X1 u1_u11_u6_U71 (.A1( u1_u11_X_39 ) , .A2( u1_u11_X_42 ) , .ZN( u1_u11_u6_n99 ) );
  INV_X1 u1_u11_u6_U72 (.A( u1_u11_X_40 ) , .ZN( u1_u11_u6_n157 ) );
  INV_X1 u1_u11_u6_U73 (.A( u1_u11_X_37 ) , .ZN( u1_u11_u6_n165 ) );
  INV_X1 u1_u11_u6_U74 (.A( u1_u11_X_38 ) , .ZN( u1_u11_u6_n162 ) );
  INV_X1 u1_u11_u6_U75 (.A( u1_u11_X_42 ) , .ZN( u1_u11_u6_n156 ) );
  NAND4_X1 u1_u11_u6_U76 (.ZN( u1_out11_32 ) , .A4( u1_u11_u6_n103 ) , .A3( u1_u11_u6_n104 ) , .A2( u1_u11_u6_n105 ) , .A1( u1_u11_u6_n106 ) );
  AOI22_X1 u1_u11_u6_U77 (.ZN( u1_u11_u6_n105 ) , .A2( u1_u11_u6_n108 ) , .A1( u1_u11_u6_n118 ) , .B2( u1_u11_u6_n126 ) , .B1( u1_u11_u6_n171 ) );
  AOI22_X1 u1_u11_u6_U78 (.ZN( u1_u11_u6_n104 ) , .A1( u1_u11_u6_n111 ) , .B1( u1_u11_u6_n124 ) , .B2( u1_u11_u6_n151 ) , .A2( u1_u11_u6_n93 ) );
  NAND4_X1 u1_u11_u6_U79 (.ZN( u1_out11_12 ) , .A4( u1_u11_u6_n114 ) , .A3( u1_u11_u6_n115 ) , .A2( u1_u11_u6_n116 ) , .A1( u1_u11_u6_n117 ) );
  AOI21_X1 u1_u11_u6_U8 (.B1( u1_u11_u6_n107 ) , .B2( u1_u11_u6_n132 ) , .A( u1_u11_u6_n158 ) , .ZN( u1_u11_u6_n88 ) );
  OAI22_X1 u1_u11_u6_U80 (.B2( u1_u11_u6_n111 ) , .ZN( u1_u11_u6_n116 ) , .B1( u1_u11_u6_n126 ) , .A2( u1_u11_u6_n164 ) , .A1( u1_u11_u6_n167 ) );
  OAI21_X1 u1_u11_u6_U81 (.A( u1_u11_u6_n108 ) , .ZN( u1_u11_u6_n117 ) , .B2( u1_u11_u6_n141 ) , .B1( u1_u11_u6_n163 ) );
  OAI211_X1 u1_u11_u6_U82 (.ZN( u1_out11_7 ) , .B( u1_u11_u6_n153 ) , .C2( u1_u11_u6_n154 ) , .C1( u1_u11_u6_n155 ) , .A( u1_u11_u6_n174 ) );
  NOR3_X1 u1_u11_u6_U83 (.A1( u1_u11_u6_n141 ) , .ZN( u1_u11_u6_n154 ) , .A3( u1_u11_u6_n164 ) , .A2( u1_u11_u6_n171 ) );
  AOI211_X1 u1_u11_u6_U84 (.B( u1_u11_u6_n149 ) , .A( u1_u11_u6_n150 ) , .C2( u1_u11_u6_n151 ) , .C1( u1_u11_u6_n152 ) , .ZN( u1_u11_u6_n153 ) );
  OAI211_X1 u1_u11_u6_U85 (.ZN( u1_out11_22 ) , .B( u1_u11_u6_n137 ) , .A( u1_u11_u6_n138 ) , .C2( u1_u11_u6_n139 ) , .C1( u1_u11_u6_n140 ) );
  AOI22_X1 u1_u11_u6_U86 (.B1( u1_u11_u6_n124 ) , .A2( u1_u11_u6_n125 ) , .A1( u1_u11_u6_n126 ) , .ZN( u1_u11_u6_n138 ) , .B2( u1_u11_u6_n161 ) );
  AND4_X1 u1_u11_u6_U87 (.A3( u1_u11_u6_n119 ) , .A1( u1_u11_u6_n120 ) , .A4( u1_u11_u6_n129 ) , .ZN( u1_u11_u6_n140 ) , .A2( u1_u11_u6_n143 ) );
  NAND3_X1 u1_u11_u6_U88 (.A2( u1_u11_u6_n123 ) , .ZN( u1_u11_u6_n125 ) , .A1( u1_u11_u6_n130 ) , .A3( u1_u11_u6_n131 ) );
  NAND3_X1 u1_u11_u6_U89 (.A3( u1_u11_u6_n133 ) , .ZN( u1_u11_u6_n141 ) , .A1( u1_u11_u6_n145 ) , .A2( u1_u11_u6_n148 ) );
  AOI21_X1 u1_u11_u6_U9 (.B2( u1_u11_u6_n147 ) , .B1( u1_u11_u6_n148 ) , .ZN( u1_u11_u6_n149 ) , .A( u1_u11_u6_n158 ) );
  NAND3_X1 u1_u11_u6_U90 (.ZN( u1_u11_u6_n101 ) , .A3( u1_u11_u6_n107 ) , .A2( u1_u11_u6_n121 ) , .A1( u1_u11_u6_n127 ) );
  NAND3_X1 u1_u11_u6_U91 (.ZN( u1_u11_u6_n102 ) , .A3( u1_u11_u6_n130 ) , .A2( u1_u11_u6_n145 ) , .A1( u1_u11_u6_n166 ) );
  NAND3_X1 u1_u11_u6_U92 (.A3( u1_u11_u6_n113 ) , .A1( u1_u11_u6_n119 ) , .A2( u1_u11_u6_n123 ) , .ZN( u1_u11_u6_n93 ) );
  NAND3_X1 u1_u11_u6_U93 (.ZN( u1_u11_u6_n142 ) , .A2( u1_u11_u6_n172 ) , .A3( u1_u11_u6_n89 ) , .A1( u1_u11_u6_n90 ) );
  AND3_X1 u1_u11_u7_U10 (.A3( u1_u11_u7_n110 ) , .A2( u1_u11_u7_n127 ) , .A1( u1_u11_u7_n132 ) , .ZN( u1_u11_u7_n92 ) );
  OAI21_X1 u1_u11_u7_U11 (.A( u1_u11_u7_n161 ) , .B1( u1_u11_u7_n168 ) , .B2( u1_u11_u7_n173 ) , .ZN( u1_u11_u7_n91 ) );
  AOI211_X1 u1_u11_u7_U12 (.A( u1_u11_u7_n117 ) , .ZN( u1_u11_u7_n118 ) , .C2( u1_u11_u7_n126 ) , .C1( u1_u11_u7_n177 ) , .B( u1_u11_u7_n180 ) );
  OAI22_X1 u1_u11_u7_U13 (.B1( u1_u11_u7_n115 ) , .ZN( u1_u11_u7_n117 ) , .A2( u1_u11_u7_n133 ) , .A1( u1_u11_u7_n137 ) , .B2( u1_u11_u7_n162 ) );
  INV_X1 u1_u11_u7_U14 (.A( u1_u11_u7_n116 ) , .ZN( u1_u11_u7_n180 ) );
  NOR3_X1 u1_u11_u7_U15 (.ZN( u1_u11_u7_n115 ) , .A3( u1_u11_u7_n145 ) , .A2( u1_u11_u7_n168 ) , .A1( u1_u11_u7_n169 ) );
  OAI211_X1 u1_u11_u7_U16 (.B( u1_u11_u7_n122 ) , .A( u1_u11_u7_n123 ) , .C2( u1_u11_u7_n124 ) , .ZN( u1_u11_u7_n154 ) , .C1( u1_u11_u7_n162 ) );
  AOI222_X1 u1_u11_u7_U17 (.ZN( u1_u11_u7_n122 ) , .C2( u1_u11_u7_n126 ) , .C1( u1_u11_u7_n145 ) , .B1( u1_u11_u7_n161 ) , .A2( u1_u11_u7_n165 ) , .B2( u1_u11_u7_n170 ) , .A1( u1_u11_u7_n176 ) );
  INV_X1 u1_u11_u7_U18 (.A( u1_u11_u7_n133 ) , .ZN( u1_u11_u7_n176 ) );
  NOR3_X1 u1_u11_u7_U19 (.A2( u1_u11_u7_n134 ) , .A1( u1_u11_u7_n135 ) , .ZN( u1_u11_u7_n136 ) , .A3( u1_u11_u7_n171 ) );
  NOR2_X1 u1_u11_u7_U20 (.A1( u1_u11_u7_n130 ) , .A2( u1_u11_u7_n134 ) , .ZN( u1_u11_u7_n153 ) );
  INV_X1 u1_u11_u7_U21 (.A( u1_u11_u7_n101 ) , .ZN( u1_u11_u7_n165 ) );
  NOR2_X1 u1_u11_u7_U22 (.ZN( u1_u11_u7_n111 ) , .A2( u1_u11_u7_n134 ) , .A1( u1_u11_u7_n169 ) );
  AOI21_X1 u1_u11_u7_U23 (.ZN( u1_u11_u7_n104 ) , .B2( u1_u11_u7_n112 ) , .B1( u1_u11_u7_n127 ) , .A( u1_u11_u7_n164 ) );
  AOI21_X1 u1_u11_u7_U24 (.ZN( u1_u11_u7_n106 ) , .B1( u1_u11_u7_n133 ) , .B2( u1_u11_u7_n146 ) , .A( u1_u11_u7_n162 ) );
  AOI21_X1 u1_u11_u7_U25 (.A( u1_u11_u7_n101 ) , .ZN( u1_u11_u7_n107 ) , .B2( u1_u11_u7_n128 ) , .B1( u1_u11_u7_n175 ) );
  INV_X1 u1_u11_u7_U26 (.A( u1_u11_u7_n138 ) , .ZN( u1_u11_u7_n171 ) );
  INV_X1 u1_u11_u7_U27 (.A( u1_u11_u7_n131 ) , .ZN( u1_u11_u7_n177 ) );
  INV_X1 u1_u11_u7_U28 (.A( u1_u11_u7_n110 ) , .ZN( u1_u11_u7_n174 ) );
  NAND2_X1 u1_u11_u7_U29 (.A1( u1_u11_u7_n129 ) , .A2( u1_u11_u7_n132 ) , .ZN( u1_u11_u7_n149 ) );
  OAI21_X1 u1_u11_u7_U3 (.ZN( u1_u11_u7_n159 ) , .A( u1_u11_u7_n165 ) , .B2( u1_u11_u7_n171 ) , .B1( u1_u11_u7_n174 ) );
  NAND2_X1 u1_u11_u7_U30 (.A1( u1_u11_u7_n113 ) , .A2( u1_u11_u7_n124 ) , .ZN( u1_u11_u7_n130 ) );
  INV_X1 u1_u11_u7_U31 (.A( u1_u11_u7_n112 ) , .ZN( u1_u11_u7_n173 ) );
  INV_X1 u1_u11_u7_U32 (.A( u1_u11_u7_n128 ) , .ZN( u1_u11_u7_n168 ) );
  INV_X1 u1_u11_u7_U33 (.A( u1_u11_u7_n148 ) , .ZN( u1_u11_u7_n169 ) );
  INV_X1 u1_u11_u7_U34 (.A( u1_u11_u7_n127 ) , .ZN( u1_u11_u7_n179 ) );
  NOR2_X1 u1_u11_u7_U35 (.ZN( u1_u11_u7_n101 ) , .A2( u1_u11_u7_n150 ) , .A1( u1_u11_u7_n156 ) );
  AOI211_X1 u1_u11_u7_U36 (.B( u1_u11_u7_n154 ) , .A( u1_u11_u7_n155 ) , .C1( u1_u11_u7_n156 ) , .ZN( u1_u11_u7_n157 ) , .C2( u1_u11_u7_n172 ) );
  INV_X1 u1_u11_u7_U37 (.A( u1_u11_u7_n153 ) , .ZN( u1_u11_u7_n172 ) );
  AOI211_X1 u1_u11_u7_U38 (.B( u1_u11_u7_n139 ) , .A( u1_u11_u7_n140 ) , .C2( u1_u11_u7_n141 ) , .ZN( u1_u11_u7_n142 ) , .C1( u1_u11_u7_n156 ) );
  AOI21_X1 u1_u11_u7_U39 (.A( u1_u11_u7_n137 ) , .B1( u1_u11_u7_n138 ) , .ZN( u1_u11_u7_n139 ) , .B2( u1_u11_u7_n146 ) );
  INV_X1 u1_u11_u7_U4 (.A( u1_u11_u7_n111 ) , .ZN( u1_u11_u7_n170 ) );
  NAND4_X1 u1_u11_u7_U40 (.A3( u1_u11_u7_n127 ) , .A2( u1_u11_u7_n128 ) , .A1( u1_u11_u7_n129 ) , .ZN( u1_u11_u7_n141 ) , .A4( u1_u11_u7_n147 ) );
  OAI22_X1 u1_u11_u7_U41 (.B1( u1_u11_u7_n136 ) , .ZN( u1_u11_u7_n140 ) , .A1( u1_u11_u7_n153 ) , .B2( u1_u11_u7_n162 ) , .A2( u1_u11_u7_n164 ) );
  AOI21_X1 u1_u11_u7_U42 (.ZN( u1_u11_u7_n123 ) , .B1( u1_u11_u7_n165 ) , .B2( u1_u11_u7_n177 ) , .A( u1_u11_u7_n97 ) );
  AOI21_X1 u1_u11_u7_U43 (.B2( u1_u11_u7_n113 ) , .B1( u1_u11_u7_n124 ) , .A( u1_u11_u7_n125 ) , .ZN( u1_u11_u7_n97 ) );
  INV_X1 u1_u11_u7_U44 (.A( u1_u11_u7_n125 ) , .ZN( u1_u11_u7_n161 ) );
  INV_X1 u1_u11_u7_U45 (.A( u1_u11_u7_n152 ) , .ZN( u1_u11_u7_n162 ) );
  AOI22_X1 u1_u11_u7_U46 (.A2( u1_u11_u7_n114 ) , .ZN( u1_u11_u7_n119 ) , .B1( u1_u11_u7_n130 ) , .A1( u1_u11_u7_n156 ) , .B2( u1_u11_u7_n165 ) );
  NAND2_X1 u1_u11_u7_U47 (.A2( u1_u11_u7_n112 ) , .ZN( u1_u11_u7_n114 ) , .A1( u1_u11_u7_n175 ) );
  AND2_X1 u1_u11_u7_U48 (.ZN( u1_u11_u7_n145 ) , .A2( u1_u11_u7_n98 ) , .A1( u1_u11_u7_n99 ) );
  NOR2_X1 u1_u11_u7_U49 (.ZN( u1_u11_u7_n137 ) , .A1( u1_u11_u7_n150 ) , .A2( u1_u11_u7_n161 ) );
  INV_X1 u1_u11_u7_U5 (.A( u1_u11_u7_n149 ) , .ZN( u1_u11_u7_n175 ) );
  AOI21_X1 u1_u11_u7_U50 (.ZN( u1_u11_u7_n105 ) , .B2( u1_u11_u7_n110 ) , .A( u1_u11_u7_n125 ) , .B1( u1_u11_u7_n147 ) );
  NAND2_X1 u1_u11_u7_U51 (.ZN( u1_u11_u7_n146 ) , .A1( u1_u11_u7_n95 ) , .A2( u1_u11_u7_n98 ) );
  NAND2_X1 u1_u11_u7_U52 (.A2( u1_u11_u7_n103 ) , .ZN( u1_u11_u7_n147 ) , .A1( u1_u11_u7_n93 ) );
  NAND2_X1 u1_u11_u7_U53 (.A1( u1_u11_u7_n103 ) , .ZN( u1_u11_u7_n127 ) , .A2( u1_u11_u7_n99 ) );
  OR2_X1 u1_u11_u7_U54 (.ZN( u1_u11_u7_n126 ) , .A2( u1_u11_u7_n152 ) , .A1( u1_u11_u7_n156 ) );
  NAND2_X1 u1_u11_u7_U55 (.A2( u1_u11_u7_n102 ) , .A1( u1_u11_u7_n103 ) , .ZN( u1_u11_u7_n133 ) );
  NAND2_X1 u1_u11_u7_U56 (.ZN( u1_u11_u7_n112 ) , .A2( u1_u11_u7_n96 ) , .A1( u1_u11_u7_n99 ) );
  NAND2_X1 u1_u11_u7_U57 (.A2( u1_u11_u7_n102 ) , .ZN( u1_u11_u7_n128 ) , .A1( u1_u11_u7_n98 ) );
  NAND2_X1 u1_u11_u7_U58 (.A1( u1_u11_u7_n100 ) , .ZN( u1_u11_u7_n113 ) , .A2( u1_u11_u7_n93 ) );
  NAND2_X1 u1_u11_u7_U59 (.A2( u1_u11_u7_n102 ) , .ZN( u1_u11_u7_n124 ) , .A1( u1_u11_u7_n96 ) );
  INV_X1 u1_u11_u7_U6 (.A( u1_u11_u7_n154 ) , .ZN( u1_u11_u7_n178 ) );
  NAND2_X1 u1_u11_u7_U60 (.ZN( u1_u11_u7_n110 ) , .A1( u1_u11_u7_n95 ) , .A2( u1_u11_u7_n96 ) );
  INV_X1 u1_u11_u7_U61 (.A( u1_u11_u7_n150 ) , .ZN( u1_u11_u7_n164 ) );
  AND2_X1 u1_u11_u7_U62 (.ZN( u1_u11_u7_n134 ) , .A1( u1_u11_u7_n93 ) , .A2( u1_u11_u7_n98 ) );
  NAND2_X1 u1_u11_u7_U63 (.A1( u1_u11_u7_n100 ) , .A2( u1_u11_u7_n102 ) , .ZN( u1_u11_u7_n129 ) );
  NAND2_X1 u1_u11_u7_U64 (.A2( u1_u11_u7_n103 ) , .ZN( u1_u11_u7_n131 ) , .A1( u1_u11_u7_n95 ) );
  NAND2_X1 u1_u11_u7_U65 (.A1( u1_u11_u7_n100 ) , .ZN( u1_u11_u7_n138 ) , .A2( u1_u11_u7_n99 ) );
  NAND2_X1 u1_u11_u7_U66 (.ZN( u1_u11_u7_n132 ) , .A1( u1_u11_u7_n93 ) , .A2( u1_u11_u7_n96 ) );
  NAND2_X1 u1_u11_u7_U67 (.A1( u1_u11_u7_n100 ) , .ZN( u1_u11_u7_n148 ) , .A2( u1_u11_u7_n95 ) );
  NOR2_X1 u1_u11_u7_U68 (.A2( u1_u11_X_47 ) , .ZN( u1_u11_u7_n150 ) , .A1( u1_u11_u7_n163 ) );
  NOR2_X1 u1_u11_u7_U69 (.A2( u1_u11_X_43 ) , .A1( u1_u11_X_44 ) , .ZN( u1_u11_u7_n103 ) );
  AOI211_X1 u1_u11_u7_U7 (.ZN( u1_u11_u7_n116 ) , .A( u1_u11_u7_n155 ) , .C1( u1_u11_u7_n161 ) , .C2( u1_u11_u7_n171 ) , .B( u1_u11_u7_n94 ) );
  NOR2_X1 u1_u11_u7_U70 (.A2( u1_u11_X_48 ) , .A1( u1_u11_u7_n166 ) , .ZN( u1_u11_u7_n95 ) );
  NOR2_X1 u1_u11_u7_U71 (.A2( u1_u11_X_45 ) , .A1( u1_u11_X_48 ) , .ZN( u1_u11_u7_n99 ) );
  NOR2_X1 u1_u11_u7_U72 (.A2( u1_u11_X_44 ) , .A1( u1_u11_u7_n167 ) , .ZN( u1_u11_u7_n98 ) );
  NOR2_X1 u1_u11_u7_U73 (.A2( u1_u11_X_46 ) , .A1( u1_u11_X_47 ) , .ZN( u1_u11_u7_n152 ) );
  AND2_X1 u1_u11_u7_U74 (.A1( u1_u11_X_47 ) , .ZN( u1_u11_u7_n156 ) , .A2( u1_u11_u7_n163 ) );
  NAND2_X1 u1_u11_u7_U75 (.A2( u1_u11_X_46 ) , .A1( u1_u11_X_47 ) , .ZN( u1_u11_u7_n125 ) );
  AND2_X1 u1_u11_u7_U76 (.A2( u1_u11_X_45 ) , .A1( u1_u11_X_48 ) , .ZN( u1_u11_u7_n102 ) );
  AND2_X1 u1_u11_u7_U77 (.A2( u1_u11_X_43 ) , .A1( u1_u11_X_44 ) , .ZN( u1_u11_u7_n96 ) );
  AND2_X1 u1_u11_u7_U78 (.A1( u1_u11_X_44 ) , .ZN( u1_u11_u7_n100 ) , .A2( u1_u11_u7_n167 ) );
  AND2_X1 u1_u11_u7_U79 (.A1( u1_u11_X_48 ) , .A2( u1_u11_u7_n166 ) , .ZN( u1_u11_u7_n93 ) );
  OAI222_X1 u1_u11_u7_U8 (.C2( u1_u11_u7_n101 ) , .B2( u1_u11_u7_n111 ) , .A1( u1_u11_u7_n113 ) , .C1( u1_u11_u7_n146 ) , .A2( u1_u11_u7_n162 ) , .B1( u1_u11_u7_n164 ) , .ZN( u1_u11_u7_n94 ) );
  INV_X1 u1_u11_u7_U80 (.A( u1_u11_X_46 ) , .ZN( u1_u11_u7_n163 ) );
  INV_X1 u1_u11_u7_U81 (.A( u1_u11_X_43 ) , .ZN( u1_u11_u7_n167 ) );
  INV_X1 u1_u11_u7_U82 (.A( u1_u11_X_45 ) , .ZN( u1_u11_u7_n166 ) );
  NAND4_X1 u1_u11_u7_U83 (.ZN( u1_out11_5 ) , .A4( u1_u11_u7_n108 ) , .A3( u1_u11_u7_n109 ) , .A1( u1_u11_u7_n116 ) , .A2( u1_u11_u7_n123 ) );
  AOI22_X1 u1_u11_u7_U84 (.ZN( u1_u11_u7_n109 ) , .A2( u1_u11_u7_n126 ) , .B2( u1_u11_u7_n145 ) , .B1( u1_u11_u7_n156 ) , .A1( u1_u11_u7_n171 ) );
  NOR4_X1 u1_u11_u7_U85 (.A4( u1_u11_u7_n104 ) , .A3( u1_u11_u7_n105 ) , .A2( u1_u11_u7_n106 ) , .A1( u1_u11_u7_n107 ) , .ZN( u1_u11_u7_n108 ) );
  NAND4_X1 u1_u11_u7_U86 (.ZN( u1_out11_27 ) , .A4( u1_u11_u7_n118 ) , .A3( u1_u11_u7_n119 ) , .A2( u1_u11_u7_n120 ) , .A1( u1_u11_u7_n121 ) );
  OAI21_X1 u1_u11_u7_U87 (.ZN( u1_u11_u7_n121 ) , .B2( u1_u11_u7_n145 ) , .A( u1_u11_u7_n150 ) , .B1( u1_u11_u7_n174 ) );
  OAI21_X1 u1_u11_u7_U88 (.ZN( u1_u11_u7_n120 ) , .A( u1_u11_u7_n161 ) , .B2( u1_u11_u7_n170 ) , .B1( u1_u11_u7_n179 ) );
  NAND4_X1 u1_u11_u7_U89 (.ZN( u1_out11_21 ) , .A4( u1_u11_u7_n157 ) , .A3( u1_u11_u7_n158 ) , .A2( u1_u11_u7_n159 ) , .A1( u1_u11_u7_n160 ) );
  OAI221_X1 u1_u11_u7_U9 (.C1( u1_u11_u7_n101 ) , .C2( u1_u11_u7_n147 ) , .ZN( u1_u11_u7_n155 ) , .B2( u1_u11_u7_n162 ) , .A( u1_u11_u7_n91 ) , .B1( u1_u11_u7_n92 ) );
  OAI21_X1 u1_u11_u7_U90 (.B1( u1_u11_u7_n145 ) , .ZN( u1_u11_u7_n160 ) , .A( u1_u11_u7_n161 ) , .B2( u1_u11_u7_n177 ) );
  AOI22_X1 u1_u11_u7_U91 (.B2( u1_u11_u7_n149 ) , .B1( u1_u11_u7_n150 ) , .A2( u1_u11_u7_n151 ) , .A1( u1_u11_u7_n152 ) , .ZN( u1_u11_u7_n158 ) );
  NAND4_X1 u1_u11_u7_U92 (.ZN( u1_out11_15 ) , .A4( u1_u11_u7_n142 ) , .A3( u1_u11_u7_n143 ) , .A2( u1_u11_u7_n144 ) , .A1( u1_u11_u7_n178 ) );
  OR2_X1 u1_u11_u7_U93 (.A2( u1_u11_u7_n125 ) , .A1( u1_u11_u7_n129 ) , .ZN( u1_u11_u7_n144 ) );
  AOI22_X1 u1_u11_u7_U94 (.A2( u1_u11_u7_n126 ) , .ZN( u1_u11_u7_n143 ) , .B2( u1_u11_u7_n165 ) , .B1( u1_u11_u7_n173 ) , .A1( u1_u11_u7_n174 ) );
  NAND3_X1 u1_u11_u7_U95 (.A3( u1_u11_u7_n146 ) , .A2( u1_u11_u7_n147 ) , .A1( u1_u11_u7_n148 ) , .ZN( u1_u11_u7_n151 ) );
  NAND3_X1 u1_u11_u7_U96 (.A3( u1_u11_u7_n131 ) , .A2( u1_u11_u7_n132 ) , .A1( u1_u11_u7_n133 ) , .ZN( u1_u11_u7_n135 ) );
  XOR2_X1 u1_u14_U35 (.B( u1_K15_22 ) , .A( u1_R13_15 ) , .Z( u1_u14_X_22 ) );
  XOR2_X1 u1_u14_U36 (.B( u1_K15_21 ) , .A( u1_R13_14 ) , .Z( u1_u14_X_21 ) );
  OAI22_X1 u1_u14_u3_U10 (.B1( u1_u14_u3_n113 ) , .A2( u1_u14_u3_n135 ) , .A1( u1_u14_u3_n150 ) , .B2( u1_u14_u3_n164 ) , .ZN( u1_u14_u3_n98 ) );
  OAI211_X1 u1_u14_u3_U11 (.B( u1_u14_u3_n106 ) , .ZN( u1_u14_u3_n119 ) , .C2( u1_u14_u3_n128 ) , .C1( u1_u14_u3_n167 ) , .A( u1_u14_u3_n181 ) );
  AOI221_X1 u1_u14_u3_U12 (.C1( u1_u14_u3_n105 ) , .ZN( u1_u14_u3_n106 ) , .A( u1_u14_u3_n131 ) , .B2( u1_u14_u3_n132 ) , .C2( u1_u14_u3_n133 ) , .B1( u1_u14_u3_n169 ) );
  INV_X1 u1_u14_u3_U13 (.ZN( u1_u14_u3_n181 ) , .A( u1_u14_u3_n98 ) );
  NAND2_X1 u1_u14_u3_U14 (.ZN( u1_u14_u3_n105 ) , .A2( u1_u14_u3_n130 ) , .A1( u1_u14_u3_n155 ) );
  AOI22_X1 u1_u14_u3_U15 (.B1( u1_u14_u3_n115 ) , .A2( u1_u14_u3_n116 ) , .ZN( u1_u14_u3_n123 ) , .B2( u1_u14_u3_n133 ) , .A1( u1_u14_u3_n169 ) );
  NAND2_X1 u1_u14_u3_U16 (.ZN( u1_u14_u3_n116 ) , .A2( u1_u14_u3_n151 ) , .A1( u1_u14_u3_n182 ) );
  NOR2_X1 u1_u14_u3_U17 (.ZN( u1_u14_u3_n126 ) , .A2( u1_u14_u3_n150 ) , .A1( u1_u14_u3_n164 ) );
  AOI21_X1 u1_u14_u3_U18 (.ZN( u1_u14_u3_n112 ) , .B2( u1_u14_u3_n146 ) , .B1( u1_u14_u3_n155 ) , .A( u1_u14_u3_n167 ) );
  NAND2_X1 u1_u14_u3_U19 (.A1( u1_u14_u3_n135 ) , .ZN( u1_u14_u3_n142 ) , .A2( u1_u14_u3_n164 ) );
  NAND2_X1 u1_u14_u3_U20 (.ZN( u1_u14_u3_n132 ) , .A2( u1_u14_u3_n152 ) , .A1( u1_u14_u3_n156 ) );
  AND2_X1 u1_u14_u3_U21 (.A2( u1_u14_u3_n113 ) , .A1( u1_u14_u3_n114 ) , .ZN( u1_u14_u3_n151 ) );
  INV_X1 u1_u14_u3_U22 (.A( u1_u14_u3_n133 ) , .ZN( u1_u14_u3_n165 ) );
  INV_X1 u1_u14_u3_U23 (.A( u1_u14_u3_n135 ) , .ZN( u1_u14_u3_n170 ) );
  NAND2_X1 u1_u14_u3_U24 (.A1( u1_u14_u3_n107 ) , .A2( u1_u14_u3_n108 ) , .ZN( u1_u14_u3_n140 ) );
  NAND2_X1 u1_u14_u3_U25 (.ZN( u1_u14_u3_n117 ) , .A1( u1_u14_u3_n124 ) , .A2( u1_u14_u3_n148 ) );
  NAND2_X1 u1_u14_u3_U26 (.ZN( u1_u14_u3_n143 ) , .A1( u1_u14_u3_n165 ) , .A2( u1_u14_u3_n167 ) );
  INV_X1 u1_u14_u3_U27 (.A( u1_u14_u3_n130 ) , .ZN( u1_u14_u3_n177 ) );
  INV_X1 u1_u14_u3_U28 (.A( u1_u14_u3_n128 ) , .ZN( u1_u14_u3_n176 ) );
  INV_X1 u1_u14_u3_U29 (.A( u1_u14_u3_n155 ) , .ZN( u1_u14_u3_n174 ) );
  INV_X1 u1_u14_u3_U3 (.A( u1_u14_u3_n129 ) , .ZN( u1_u14_u3_n183 ) );
  INV_X1 u1_u14_u3_U30 (.A( u1_u14_u3_n139 ) , .ZN( u1_u14_u3_n185 ) );
  NOR2_X1 u1_u14_u3_U31 (.ZN( u1_u14_u3_n135 ) , .A2( u1_u14_u3_n141 ) , .A1( u1_u14_u3_n169 ) );
  OAI222_X1 u1_u14_u3_U32 (.C2( u1_u14_u3_n107 ) , .A2( u1_u14_u3_n108 ) , .B1( u1_u14_u3_n135 ) , .ZN( u1_u14_u3_n138 ) , .B2( u1_u14_u3_n146 ) , .C1( u1_u14_u3_n154 ) , .A1( u1_u14_u3_n164 ) );
  NOR4_X1 u1_u14_u3_U33 (.A4( u1_u14_u3_n157 ) , .A3( u1_u14_u3_n158 ) , .A2( u1_u14_u3_n159 ) , .A1( u1_u14_u3_n160 ) , .ZN( u1_u14_u3_n161 ) );
  AOI21_X1 u1_u14_u3_U34 (.B2( u1_u14_u3_n152 ) , .B1( u1_u14_u3_n153 ) , .ZN( u1_u14_u3_n158 ) , .A( u1_u14_u3_n164 ) );
  AOI21_X1 u1_u14_u3_U35 (.A( u1_u14_u3_n154 ) , .B2( u1_u14_u3_n155 ) , .B1( u1_u14_u3_n156 ) , .ZN( u1_u14_u3_n157 ) );
  AOI21_X1 u1_u14_u3_U36 (.A( u1_u14_u3_n149 ) , .B2( u1_u14_u3_n150 ) , .B1( u1_u14_u3_n151 ) , .ZN( u1_u14_u3_n159 ) );
  AOI211_X1 u1_u14_u3_U37 (.ZN( u1_u14_u3_n109 ) , .A( u1_u14_u3_n119 ) , .C2( u1_u14_u3_n129 ) , .B( u1_u14_u3_n138 ) , .C1( u1_u14_u3_n141 ) );
  AOI211_X1 u1_u14_u3_U38 (.B( u1_u14_u3_n119 ) , .A( u1_u14_u3_n120 ) , .C2( u1_u14_u3_n121 ) , .ZN( u1_u14_u3_n122 ) , .C1( u1_u14_u3_n179 ) );
  INV_X1 u1_u14_u3_U39 (.A( u1_u14_u3_n156 ) , .ZN( u1_u14_u3_n179 ) );
  INV_X1 u1_u14_u3_U4 (.A( u1_u14_u3_n140 ) , .ZN( u1_u14_u3_n182 ) );
  OAI22_X1 u1_u14_u3_U40 (.B1( u1_u14_u3_n118 ) , .ZN( u1_u14_u3_n120 ) , .A1( u1_u14_u3_n135 ) , .B2( u1_u14_u3_n154 ) , .A2( u1_u14_u3_n178 ) );
  AND3_X1 u1_u14_u3_U41 (.ZN( u1_u14_u3_n118 ) , .A2( u1_u14_u3_n124 ) , .A1( u1_u14_u3_n144 ) , .A3( u1_u14_u3_n152 ) );
  INV_X1 u1_u14_u3_U42 (.A( u1_u14_u3_n121 ) , .ZN( u1_u14_u3_n164 ) );
  NAND2_X1 u1_u14_u3_U43 (.ZN( u1_u14_u3_n133 ) , .A1( u1_u14_u3_n154 ) , .A2( u1_u14_u3_n164 ) );
  OAI211_X1 u1_u14_u3_U44 (.B( u1_u14_u3_n127 ) , .ZN( u1_u14_u3_n139 ) , .C1( u1_u14_u3_n150 ) , .C2( u1_u14_u3_n154 ) , .A( u1_u14_u3_n184 ) );
  INV_X1 u1_u14_u3_U45 (.A( u1_u14_u3_n125 ) , .ZN( u1_u14_u3_n184 ) );
  AOI221_X1 u1_u14_u3_U46 (.A( u1_u14_u3_n126 ) , .ZN( u1_u14_u3_n127 ) , .C2( u1_u14_u3_n132 ) , .C1( u1_u14_u3_n169 ) , .B2( u1_u14_u3_n170 ) , .B1( u1_u14_u3_n174 ) );
  OAI22_X1 u1_u14_u3_U47 (.A1( u1_u14_u3_n124 ) , .ZN( u1_u14_u3_n125 ) , .B2( u1_u14_u3_n145 ) , .A2( u1_u14_u3_n165 ) , .B1( u1_u14_u3_n167 ) );
  NOR2_X1 u1_u14_u3_U48 (.A1( u1_u14_u3_n113 ) , .ZN( u1_u14_u3_n131 ) , .A2( u1_u14_u3_n154 ) );
  NAND2_X1 u1_u14_u3_U49 (.A1( u1_u14_u3_n103 ) , .ZN( u1_u14_u3_n150 ) , .A2( u1_u14_u3_n99 ) );
  INV_X1 u1_u14_u3_U5 (.A( u1_u14_u3_n117 ) , .ZN( u1_u14_u3_n178 ) );
  NAND2_X1 u1_u14_u3_U50 (.A2( u1_u14_u3_n102 ) , .ZN( u1_u14_u3_n155 ) , .A1( u1_u14_u3_n97 ) );
  INV_X1 u1_u14_u3_U51 (.A( u1_u14_u3_n141 ) , .ZN( u1_u14_u3_n167 ) );
  AOI21_X1 u1_u14_u3_U52 (.B2( u1_u14_u3_n114 ) , .B1( u1_u14_u3_n146 ) , .A( u1_u14_u3_n154 ) , .ZN( u1_u14_u3_n94 ) );
  AOI21_X1 u1_u14_u3_U53 (.ZN( u1_u14_u3_n110 ) , .B2( u1_u14_u3_n142 ) , .B1( u1_u14_u3_n186 ) , .A( u1_u14_u3_n95 ) );
  INV_X1 u1_u14_u3_U54 (.A( u1_u14_u3_n145 ) , .ZN( u1_u14_u3_n186 ) );
  AOI21_X1 u1_u14_u3_U55 (.B1( u1_u14_u3_n124 ) , .A( u1_u14_u3_n149 ) , .B2( u1_u14_u3_n155 ) , .ZN( u1_u14_u3_n95 ) );
  INV_X1 u1_u14_u3_U56 (.A( u1_u14_u3_n149 ) , .ZN( u1_u14_u3_n169 ) );
  NAND2_X1 u1_u14_u3_U57 (.ZN( u1_u14_u3_n124 ) , .A1( u1_u14_u3_n96 ) , .A2( u1_u14_u3_n97 ) );
  NAND2_X1 u1_u14_u3_U58 (.A2( u1_u14_u3_n100 ) , .ZN( u1_u14_u3_n146 ) , .A1( u1_u14_u3_n96 ) );
  NAND2_X1 u1_u14_u3_U59 (.A1( u1_u14_u3_n101 ) , .ZN( u1_u14_u3_n145 ) , .A2( u1_u14_u3_n99 ) );
  AOI221_X1 u1_u14_u3_U6 (.A( u1_u14_u3_n131 ) , .C2( u1_u14_u3_n132 ) , .C1( u1_u14_u3_n133 ) , .ZN( u1_u14_u3_n134 ) , .B1( u1_u14_u3_n143 ) , .B2( u1_u14_u3_n177 ) );
  NAND2_X1 u1_u14_u3_U60 (.A1( u1_u14_u3_n100 ) , .ZN( u1_u14_u3_n156 ) , .A2( u1_u14_u3_n99 ) );
  NAND2_X1 u1_u14_u3_U61 (.A2( u1_u14_u3_n101 ) , .A1( u1_u14_u3_n104 ) , .ZN( u1_u14_u3_n148 ) );
  NAND2_X1 u1_u14_u3_U62 (.A1( u1_u14_u3_n100 ) , .A2( u1_u14_u3_n102 ) , .ZN( u1_u14_u3_n128 ) );
  NAND2_X1 u1_u14_u3_U63 (.A2( u1_u14_u3_n101 ) , .A1( u1_u14_u3_n102 ) , .ZN( u1_u14_u3_n152 ) );
  NAND2_X1 u1_u14_u3_U64 (.A2( u1_u14_u3_n101 ) , .ZN( u1_u14_u3_n114 ) , .A1( u1_u14_u3_n96 ) );
  NAND2_X1 u1_u14_u3_U65 (.ZN( u1_u14_u3_n107 ) , .A1( u1_u14_u3_n97 ) , .A2( u1_u14_u3_n99 ) );
  NAND2_X1 u1_u14_u3_U66 (.A2( u1_u14_u3_n100 ) , .A1( u1_u14_u3_n104 ) , .ZN( u1_u14_u3_n113 ) );
  NAND2_X1 u1_u14_u3_U67 (.A1( u1_u14_u3_n104 ) , .ZN( u1_u14_u3_n153 ) , .A2( u1_u14_u3_n97 ) );
  NAND2_X1 u1_u14_u3_U68 (.A2( u1_u14_u3_n103 ) , .A1( u1_u14_u3_n104 ) , .ZN( u1_u14_u3_n130 ) );
  NAND2_X1 u1_u14_u3_U69 (.A2( u1_u14_u3_n103 ) , .ZN( u1_u14_u3_n144 ) , .A1( u1_u14_u3_n96 ) );
  OAI22_X1 u1_u14_u3_U7 (.B2( u1_u14_u3_n147 ) , .A2( u1_u14_u3_n148 ) , .ZN( u1_u14_u3_n160 ) , .B1( u1_u14_u3_n165 ) , .A1( u1_u14_u3_n168 ) );
  NAND2_X1 u1_u14_u3_U70 (.A1( u1_u14_u3_n102 ) , .A2( u1_u14_u3_n103 ) , .ZN( u1_u14_u3_n108 ) );
  NOR2_X1 u1_u14_u3_U71 (.A2( u1_u14_X_19 ) , .A1( u1_u14_X_20 ) , .ZN( u1_u14_u3_n99 ) );
  NOR2_X1 u1_u14_u3_U72 (.A2( u1_u14_X_21 ) , .A1( u1_u14_X_24 ) , .ZN( u1_u14_u3_n103 ) );
  NOR2_X1 u1_u14_u3_U73 (.A2( u1_u14_X_24 ) , .A1( u1_u14_u3_n171 ) , .ZN( u1_u14_u3_n97 ) );
  NOR2_X1 u1_u14_u3_U74 (.A2( u1_u14_X_23 ) , .ZN( u1_u14_u3_n141 ) , .A1( u1_u14_u3_n166 ) );
  NOR2_X1 u1_u14_u3_U75 (.A2( u1_u14_X_19 ) , .A1( u1_u14_u3_n172 ) , .ZN( u1_u14_u3_n96 ) );
  NAND2_X1 u1_u14_u3_U76 (.A1( u1_u14_X_22 ) , .A2( u1_u14_X_23 ) , .ZN( u1_u14_u3_n154 ) );
  NAND2_X1 u1_u14_u3_U77 (.A1( u1_u14_X_23 ) , .ZN( u1_u14_u3_n149 ) , .A2( u1_u14_u3_n166 ) );
  NOR2_X1 u1_u14_u3_U78 (.A2( u1_u14_X_22 ) , .A1( u1_u14_X_23 ) , .ZN( u1_u14_u3_n121 ) );
  AND2_X1 u1_u14_u3_U79 (.A1( u1_u14_X_24 ) , .ZN( u1_u14_u3_n101 ) , .A2( u1_u14_u3_n171 ) );
  AND3_X1 u1_u14_u3_U8 (.A3( u1_u14_u3_n144 ) , .A2( u1_u14_u3_n145 ) , .A1( u1_u14_u3_n146 ) , .ZN( u1_u14_u3_n147 ) );
  AND2_X1 u1_u14_u3_U80 (.A1( u1_u14_X_19 ) , .ZN( u1_u14_u3_n102 ) , .A2( u1_u14_u3_n172 ) );
  AND2_X1 u1_u14_u3_U81 (.A1( u1_u14_X_21 ) , .A2( u1_u14_X_24 ) , .ZN( u1_u14_u3_n100 ) );
  AND2_X1 u1_u14_u3_U82 (.A2( u1_u14_X_19 ) , .A1( u1_u14_X_20 ) , .ZN( u1_u14_u3_n104 ) );
  INV_X1 u1_u14_u3_U83 (.A( u1_u14_X_22 ) , .ZN( u1_u14_u3_n166 ) );
  INV_X1 u1_u14_u3_U84 (.A( u1_u14_X_21 ) , .ZN( u1_u14_u3_n171 ) );
  INV_X1 u1_u14_u3_U85 (.A( u1_u14_X_20 ) , .ZN( u1_u14_u3_n172 ) );
  NAND4_X1 u1_u14_u3_U86 (.ZN( u1_out14_26 ) , .A4( u1_u14_u3_n109 ) , .A3( u1_u14_u3_n110 ) , .A2( u1_u14_u3_n111 ) , .A1( u1_u14_u3_n173 ) );
  INV_X1 u1_u14_u3_U87 (.ZN( u1_u14_u3_n173 ) , .A( u1_u14_u3_n94 ) );
  OAI21_X1 u1_u14_u3_U88 (.ZN( u1_u14_u3_n111 ) , .B2( u1_u14_u3_n117 ) , .A( u1_u14_u3_n133 ) , .B1( u1_u14_u3_n176 ) );
  NAND4_X1 u1_u14_u3_U89 (.ZN( u1_out14_20 ) , .A4( u1_u14_u3_n122 ) , .A3( u1_u14_u3_n123 ) , .A1( u1_u14_u3_n175 ) , .A2( u1_u14_u3_n180 ) );
  INV_X1 u1_u14_u3_U9 (.A( u1_u14_u3_n143 ) , .ZN( u1_u14_u3_n168 ) );
  INV_X1 u1_u14_u3_U90 (.A( u1_u14_u3_n126 ) , .ZN( u1_u14_u3_n180 ) );
  INV_X1 u1_u14_u3_U91 (.A( u1_u14_u3_n112 ) , .ZN( u1_u14_u3_n175 ) );
  NAND4_X1 u1_u14_u3_U92 (.ZN( u1_out14_1 ) , .A4( u1_u14_u3_n161 ) , .A3( u1_u14_u3_n162 ) , .A2( u1_u14_u3_n163 ) , .A1( u1_u14_u3_n185 ) );
  NAND2_X1 u1_u14_u3_U93 (.ZN( u1_u14_u3_n163 ) , .A2( u1_u14_u3_n170 ) , .A1( u1_u14_u3_n176 ) );
  AOI22_X1 u1_u14_u3_U94 (.B2( u1_u14_u3_n140 ) , .B1( u1_u14_u3_n141 ) , .A2( u1_u14_u3_n142 ) , .ZN( u1_u14_u3_n162 ) , .A1( u1_u14_u3_n177 ) );
  OR4_X1 u1_u14_u3_U95 (.ZN( u1_out14_10 ) , .A4( u1_u14_u3_n136 ) , .A3( u1_u14_u3_n137 ) , .A1( u1_u14_u3_n138 ) , .A2( u1_u14_u3_n139 ) );
  OAI222_X1 u1_u14_u3_U96 (.C1( u1_u14_u3_n128 ) , .ZN( u1_u14_u3_n137 ) , .B1( u1_u14_u3_n148 ) , .A2( u1_u14_u3_n150 ) , .B2( u1_u14_u3_n154 ) , .C2( u1_u14_u3_n164 ) , .A1( u1_u14_u3_n167 ) );
  OAI221_X1 u1_u14_u3_U97 (.A( u1_u14_u3_n134 ) , .B2( u1_u14_u3_n135 ) , .ZN( u1_u14_u3_n136 ) , .C1( u1_u14_u3_n149 ) , .B1( u1_u14_u3_n151 ) , .C2( u1_u14_u3_n183 ) );
  NAND3_X1 u1_u14_u3_U98 (.A1( u1_u14_u3_n114 ) , .ZN( u1_u14_u3_n115 ) , .A2( u1_u14_u3_n145 ) , .A3( u1_u14_u3_n153 ) );
  NAND3_X1 u1_u14_u3_U99 (.ZN( u1_u14_u3_n129 ) , .A2( u1_u14_u3_n144 ) , .A1( u1_u14_u3_n153 ) , .A3( u1_u14_u3_n182 ) );
  XOR2_X1 u1_u15_U22 (.A( u1_FP_55 ) , .B( u1_K16_34 ) , .Z( u1_u15_X_34 ) );
  XOR2_X1 u1_u15_U23 (.A( u1_FP_54 ) , .B( u1_K16_33 ) , .Z( u1_u15_X_33 ) );
  XOR2_X1 u1_u15_U42 (.A( u1_FP_43 ) , .B( u1_K16_16 ) , .Z( u1_u15_X_16 ) );
  XOR2_X1 u1_u15_U43 (.A( u1_FP_42 ) , .B( u1_K16_15 ) , .Z( u1_u15_X_15 ) );
  OAI22_X1 u1_u15_u2_U10 (.B1( u1_u15_u2_n151 ) , .A2( u1_u15_u2_n152 ) , .A1( u1_u15_u2_n153 ) , .ZN( u1_u15_u2_n160 ) , .B2( u1_u15_u2_n168 ) );
  NAND3_X1 u1_u15_u2_U100 (.A2( u1_u15_u2_n100 ) , .A1( u1_u15_u2_n104 ) , .A3( u1_u15_u2_n138 ) , .ZN( u1_u15_u2_n98 ) );
  NOR3_X1 u1_u15_u2_U11 (.A1( u1_u15_u2_n150 ) , .ZN( u1_u15_u2_n151 ) , .A3( u1_u15_u2_n175 ) , .A2( u1_u15_u2_n188 ) );
  AOI21_X1 u1_u15_u2_U12 (.B2( u1_u15_u2_n123 ) , .ZN( u1_u15_u2_n125 ) , .A( u1_u15_u2_n171 ) , .B1( u1_u15_u2_n184 ) );
  INV_X1 u1_u15_u2_U13 (.A( u1_u15_u2_n150 ) , .ZN( u1_u15_u2_n184 ) );
  AOI21_X1 u1_u15_u2_U14 (.ZN( u1_u15_u2_n144 ) , .B2( u1_u15_u2_n155 ) , .A( u1_u15_u2_n172 ) , .B1( u1_u15_u2_n185 ) );
  AOI21_X1 u1_u15_u2_U15 (.B2( u1_u15_u2_n143 ) , .ZN( u1_u15_u2_n145 ) , .B1( u1_u15_u2_n152 ) , .A( u1_u15_u2_n171 ) );
  INV_X1 u1_u15_u2_U16 (.A( u1_u15_u2_n156 ) , .ZN( u1_u15_u2_n171 ) );
  INV_X1 u1_u15_u2_U17 (.A( u1_u15_u2_n120 ) , .ZN( u1_u15_u2_n188 ) );
  NAND2_X1 u1_u15_u2_U18 (.A2( u1_u15_u2_n122 ) , .ZN( u1_u15_u2_n150 ) , .A1( u1_u15_u2_n152 ) );
  INV_X1 u1_u15_u2_U19 (.A( u1_u15_u2_n153 ) , .ZN( u1_u15_u2_n170 ) );
  INV_X1 u1_u15_u2_U20 (.A( u1_u15_u2_n137 ) , .ZN( u1_u15_u2_n173 ) );
  NAND2_X1 u1_u15_u2_U21 (.A1( u1_u15_u2_n132 ) , .A2( u1_u15_u2_n139 ) , .ZN( u1_u15_u2_n157 ) );
  INV_X1 u1_u15_u2_U22 (.A( u1_u15_u2_n113 ) , .ZN( u1_u15_u2_n178 ) );
  INV_X1 u1_u15_u2_U23 (.A( u1_u15_u2_n139 ) , .ZN( u1_u15_u2_n175 ) );
  INV_X1 u1_u15_u2_U24 (.A( u1_u15_u2_n155 ) , .ZN( u1_u15_u2_n181 ) );
  INV_X1 u1_u15_u2_U25 (.A( u1_u15_u2_n119 ) , .ZN( u1_u15_u2_n177 ) );
  INV_X1 u1_u15_u2_U26 (.A( u1_u15_u2_n116 ) , .ZN( u1_u15_u2_n180 ) );
  INV_X1 u1_u15_u2_U27 (.A( u1_u15_u2_n131 ) , .ZN( u1_u15_u2_n179 ) );
  INV_X1 u1_u15_u2_U28 (.A( u1_u15_u2_n154 ) , .ZN( u1_u15_u2_n176 ) );
  NAND2_X1 u1_u15_u2_U29 (.A2( u1_u15_u2_n116 ) , .A1( u1_u15_u2_n117 ) , .ZN( u1_u15_u2_n118 ) );
  NOR2_X1 u1_u15_u2_U3 (.ZN( u1_u15_u2_n121 ) , .A2( u1_u15_u2_n177 ) , .A1( u1_u15_u2_n180 ) );
  INV_X1 u1_u15_u2_U30 (.A( u1_u15_u2_n132 ) , .ZN( u1_u15_u2_n182 ) );
  INV_X1 u1_u15_u2_U31 (.A( u1_u15_u2_n158 ) , .ZN( u1_u15_u2_n183 ) );
  OAI21_X1 u1_u15_u2_U32 (.A( u1_u15_u2_n156 ) , .B1( u1_u15_u2_n157 ) , .ZN( u1_u15_u2_n158 ) , .B2( u1_u15_u2_n179 ) );
  NOR2_X1 u1_u15_u2_U33 (.ZN( u1_u15_u2_n156 ) , .A1( u1_u15_u2_n166 ) , .A2( u1_u15_u2_n169 ) );
  NOR2_X1 u1_u15_u2_U34 (.A2( u1_u15_u2_n114 ) , .ZN( u1_u15_u2_n137 ) , .A1( u1_u15_u2_n140 ) );
  NOR2_X1 u1_u15_u2_U35 (.A2( u1_u15_u2_n138 ) , .ZN( u1_u15_u2_n153 ) , .A1( u1_u15_u2_n156 ) );
  AOI211_X1 u1_u15_u2_U36 (.ZN( u1_u15_u2_n130 ) , .C1( u1_u15_u2_n138 ) , .C2( u1_u15_u2_n179 ) , .B( u1_u15_u2_n96 ) , .A( u1_u15_u2_n97 ) );
  OAI22_X1 u1_u15_u2_U37 (.B1( u1_u15_u2_n133 ) , .A2( u1_u15_u2_n137 ) , .A1( u1_u15_u2_n152 ) , .B2( u1_u15_u2_n168 ) , .ZN( u1_u15_u2_n97 ) );
  OAI221_X1 u1_u15_u2_U38 (.B1( u1_u15_u2_n113 ) , .C1( u1_u15_u2_n132 ) , .A( u1_u15_u2_n149 ) , .B2( u1_u15_u2_n171 ) , .C2( u1_u15_u2_n172 ) , .ZN( u1_u15_u2_n96 ) );
  OAI221_X1 u1_u15_u2_U39 (.A( u1_u15_u2_n115 ) , .C2( u1_u15_u2_n123 ) , .B2( u1_u15_u2_n143 ) , .B1( u1_u15_u2_n153 ) , .ZN( u1_u15_u2_n163 ) , .C1( u1_u15_u2_n168 ) );
  INV_X1 u1_u15_u2_U4 (.A( u1_u15_u2_n134 ) , .ZN( u1_u15_u2_n185 ) );
  OAI21_X1 u1_u15_u2_U40 (.A( u1_u15_u2_n114 ) , .ZN( u1_u15_u2_n115 ) , .B1( u1_u15_u2_n176 ) , .B2( u1_u15_u2_n178 ) );
  OAI221_X1 u1_u15_u2_U41 (.A( u1_u15_u2_n135 ) , .B2( u1_u15_u2_n136 ) , .B1( u1_u15_u2_n137 ) , .ZN( u1_u15_u2_n162 ) , .C2( u1_u15_u2_n167 ) , .C1( u1_u15_u2_n185 ) );
  AND3_X1 u1_u15_u2_U42 (.A3( u1_u15_u2_n131 ) , .A2( u1_u15_u2_n132 ) , .A1( u1_u15_u2_n133 ) , .ZN( u1_u15_u2_n136 ) );
  AOI22_X1 u1_u15_u2_U43 (.ZN( u1_u15_u2_n135 ) , .B1( u1_u15_u2_n140 ) , .A1( u1_u15_u2_n156 ) , .B2( u1_u15_u2_n180 ) , .A2( u1_u15_u2_n188 ) );
  AOI21_X1 u1_u15_u2_U44 (.ZN( u1_u15_u2_n149 ) , .B1( u1_u15_u2_n173 ) , .B2( u1_u15_u2_n188 ) , .A( u1_u15_u2_n95 ) );
  AND3_X1 u1_u15_u2_U45 (.A2( u1_u15_u2_n100 ) , .A1( u1_u15_u2_n104 ) , .A3( u1_u15_u2_n156 ) , .ZN( u1_u15_u2_n95 ) );
  OAI21_X1 u1_u15_u2_U46 (.A( u1_u15_u2_n101 ) , .B2( u1_u15_u2_n121 ) , .B1( u1_u15_u2_n153 ) , .ZN( u1_u15_u2_n164 ) );
  NAND2_X1 u1_u15_u2_U47 (.A2( u1_u15_u2_n100 ) , .A1( u1_u15_u2_n107 ) , .ZN( u1_u15_u2_n155 ) );
  NAND2_X1 u1_u15_u2_U48 (.A2( u1_u15_u2_n105 ) , .A1( u1_u15_u2_n108 ) , .ZN( u1_u15_u2_n143 ) );
  NAND2_X1 u1_u15_u2_U49 (.A1( u1_u15_u2_n104 ) , .A2( u1_u15_u2_n106 ) , .ZN( u1_u15_u2_n152 ) );
  NOR4_X1 u1_u15_u2_U5 (.A4( u1_u15_u2_n124 ) , .A3( u1_u15_u2_n125 ) , .A2( u1_u15_u2_n126 ) , .A1( u1_u15_u2_n127 ) , .ZN( u1_u15_u2_n128 ) );
  NAND2_X1 u1_u15_u2_U50 (.A1( u1_u15_u2_n100 ) , .A2( u1_u15_u2_n105 ) , .ZN( u1_u15_u2_n132 ) );
  INV_X1 u1_u15_u2_U51 (.A( u1_u15_u2_n140 ) , .ZN( u1_u15_u2_n168 ) );
  INV_X1 u1_u15_u2_U52 (.A( u1_u15_u2_n138 ) , .ZN( u1_u15_u2_n167 ) );
  OAI21_X1 u1_u15_u2_U53 (.A( u1_u15_u2_n141 ) , .B2( u1_u15_u2_n142 ) , .ZN( u1_u15_u2_n146 ) , .B1( u1_u15_u2_n153 ) );
  OAI21_X1 u1_u15_u2_U54 (.A( u1_u15_u2_n140 ) , .ZN( u1_u15_u2_n141 ) , .B1( u1_u15_u2_n176 ) , .B2( u1_u15_u2_n177 ) );
  NOR3_X1 u1_u15_u2_U55 (.ZN( u1_u15_u2_n142 ) , .A3( u1_u15_u2_n175 ) , .A2( u1_u15_u2_n178 ) , .A1( u1_u15_u2_n181 ) );
  INV_X1 u1_u15_u2_U56 (.ZN( u1_u15_u2_n187 ) , .A( u1_u15_u2_n99 ) );
  OAI21_X1 u1_u15_u2_U57 (.B1( u1_u15_u2_n137 ) , .B2( u1_u15_u2_n143 ) , .A( u1_u15_u2_n98 ) , .ZN( u1_u15_u2_n99 ) );
  NAND2_X1 u1_u15_u2_U58 (.A1( u1_u15_u2_n102 ) , .A2( u1_u15_u2_n106 ) , .ZN( u1_u15_u2_n113 ) );
  NAND2_X1 u1_u15_u2_U59 (.A1( u1_u15_u2_n106 ) , .A2( u1_u15_u2_n107 ) , .ZN( u1_u15_u2_n131 ) );
  AOI21_X1 u1_u15_u2_U6 (.B2( u1_u15_u2_n119 ) , .ZN( u1_u15_u2_n127 ) , .A( u1_u15_u2_n137 ) , .B1( u1_u15_u2_n155 ) );
  NAND2_X1 u1_u15_u2_U60 (.A1( u1_u15_u2_n103 ) , .A2( u1_u15_u2_n107 ) , .ZN( u1_u15_u2_n139 ) );
  NAND2_X1 u1_u15_u2_U61 (.A1( u1_u15_u2_n103 ) , .A2( u1_u15_u2_n105 ) , .ZN( u1_u15_u2_n133 ) );
  NAND2_X1 u1_u15_u2_U62 (.A1( u1_u15_u2_n102 ) , .A2( u1_u15_u2_n103 ) , .ZN( u1_u15_u2_n154 ) );
  NAND2_X1 u1_u15_u2_U63 (.A2( u1_u15_u2_n103 ) , .A1( u1_u15_u2_n104 ) , .ZN( u1_u15_u2_n119 ) );
  NAND2_X1 u1_u15_u2_U64 (.A2( u1_u15_u2_n107 ) , .A1( u1_u15_u2_n108 ) , .ZN( u1_u15_u2_n123 ) );
  NAND2_X1 u1_u15_u2_U65 (.A1( u1_u15_u2_n104 ) , .A2( u1_u15_u2_n108 ) , .ZN( u1_u15_u2_n122 ) );
  INV_X1 u1_u15_u2_U66 (.A( u1_u15_u2_n114 ) , .ZN( u1_u15_u2_n172 ) );
  NAND2_X1 u1_u15_u2_U67 (.A2( u1_u15_u2_n100 ) , .A1( u1_u15_u2_n102 ) , .ZN( u1_u15_u2_n116 ) );
  NAND2_X1 u1_u15_u2_U68 (.A1( u1_u15_u2_n102 ) , .A2( u1_u15_u2_n108 ) , .ZN( u1_u15_u2_n120 ) );
  NAND2_X1 u1_u15_u2_U69 (.A2( u1_u15_u2_n105 ) , .A1( u1_u15_u2_n106 ) , .ZN( u1_u15_u2_n117 ) );
  AOI21_X1 u1_u15_u2_U7 (.ZN( u1_u15_u2_n124 ) , .B1( u1_u15_u2_n131 ) , .B2( u1_u15_u2_n143 ) , .A( u1_u15_u2_n172 ) );
  NOR2_X1 u1_u15_u2_U70 (.A2( u1_u15_X_16 ) , .ZN( u1_u15_u2_n140 ) , .A1( u1_u15_u2_n166 ) );
  NOR2_X1 u1_u15_u2_U71 (.A2( u1_u15_X_13 ) , .A1( u1_u15_X_14 ) , .ZN( u1_u15_u2_n100 ) );
  NOR2_X1 u1_u15_u2_U72 (.A2( u1_u15_X_16 ) , .A1( u1_u15_X_17 ) , .ZN( u1_u15_u2_n138 ) );
  NOR2_X1 u1_u15_u2_U73 (.A2( u1_u15_X_15 ) , .A1( u1_u15_X_18 ) , .ZN( u1_u15_u2_n104 ) );
  NOR2_X1 u1_u15_u2_U74 (.A2( u1_u15_X_14 ) , .ZN( u1_u15_u2_n103 ) , .A1( u1_u15_u2_n174 ) );
  NOR2_X1 u1_u15_u2_U75 (.A2( u1_u15_X_15 ) , .ZN( u1_u15_u2_n102 ) , .A1( u1_u15_u2_n165 ) );
  NOR2_X1 u1_u15_u2_U76 (.A2( u1_u15_X_17 ) , .ZN( u1_u15_u2_n114 ) , .A1( u1_u15_u2_n169 ) );
  AND2_X1 u1_u15_u2_U77 (.A1( u1_u15_X_15 ) , .ZN( u1_u15_u2_n105 ) , .A2( u1_u15_u2_n165 ) );
  AND2_X1 u1_u15_u2_U78 (.A2( u1_u15_X_15 ) , .A1( u1_u15_X_18 ) , .ZN( u1_u15_u2_n107 ) );
  AND2_X1 u1_u15_u2_U79 (.A1( u1_u15_X_14 ) , .ZN( u1_u15_u2_n106 ) , .A2( u1_u15_u2_n174 ) );
  AOI21_X1 u1_u15_u2_U8 (.B2( u1_u15_u2_n120 ) , .B1( u1_u15_u2_n121 ) , .ZN( u1_u15_u2_n126 ) , .A( u1_u15_u2_n167 ) );
  AND2_X1 u1_u15_u2_U80 (.A1( u1_u15_X_13 ) , .A2( u1_u15_X_14 ) , .ZN( u1_u15_u2_n108 ) );
  INV_X1 u1_u15_u2_U81 (.A( u1_u15_X_16 ) , .ZN( u1_u15_u2_n169 ) );
  INV_X1 u1_u15_u2_U82 (.A( u1_u15_X_17 ) , .ZN( u1_u15_u2_n166 ) );
  INV_X1 u1_u15_u2_U83 (.A( u1_u15_X_13 ) , .ZN( u1_u15_u2_n174 ) );
  INV_X1 u1_u15_u2_U84 (.A( u1_u15_X_18 ) , .ZN( u1_u15_u2_n165 ) );
  NAND4_X1 u1_u15_u2_U85 (.ZN( u1_out15_30 ) , .A4( u1_u15_u2_n147 ) , .A3( u1_u15_u2_n148 ) , .A2( u1_u15_u2_n149 ) , .A1( u1_u15_u2_n187 ) );
  NOR3_X1 u1_u15_u2_U86 (.A3( u1_u15_u2_n144 ) , .A2( u1_u15_u2_n145 ) , .A1( u1_u15_u2_n146 ) , .ZN( u1_u15_u2_n147 ) );
  AOI21_X1 u1_u15_u2_U87 (.B2( u1_u15_u2_n138 ) , .ZN( u1_u15_u2_n148 ) , .A( u1_u15_u2_n162 ) , .B1( u1_u15_u2_n182 ) );
  NAND4_X1 u1_u15_u2_U88 (.ZN( u1_out15_24 ) , .A4( u1_u15_u2_n111 ) , .A3( u1_u15_u2_n112 ) , .A1( u1_u15_u2_n130 ) , .A2( u1_u15_u2_n187 ) );
  AOI221_X1 u1_u15_u2_U89 (.A( u1_u15_u2_n109 ) , .B1( u1_u15_u2_n110 ) , .ZN( u1_u15_u2_n111 ) , .C1( u1_u15_u2_n134 ) , .C2( u1_u15_u2_n170 ) , .B2( u1_u15_u2_n173 ) );
  OAI22_X1 u1_u15_u2_U9 (.ZN( u1_u15_u2_n109 ) , .A2( u1_u15_u2_n113 ) , .B2( u1_u15_u2_n133 ) , .B1( u1_u15_u2_n167 ) , .A1( u1_u15_u2_n168 ) );
  AOI21_X1 u1_u15_u2_U90 (.ZN( u1_u15_u2_n112 ) , .B2( u1_u15_u2_n156 ) , .A( u1_u15_u2_n164 ) , .B1( u1_u15_u2_n181 ) );
  NAND4_X1 u1_u15_u2_U91 (.ZN( u1_out15_16 ) , .A4( u1_u15_u2_n128 ) , .A3( u1_u15_u2_n129 ) , .A1( u1_u15_u2_n130 ) , .A2( u1_u15_u2_n186 ) );
  AOI22_X1 u1_u15_u2_U92 (.A2( u1_u15_u2_n118 ) , .ZN( u1_u15_u2_n129 ) , .A1( u1_u15_u2_n140 ) , .B1( u1_u15_u2_n157 ) , .B2( u1_u15_u2_n170 ) );
  INV_X1 u1_u15_u2_U93 (.A( u1_u15_u2_n163 ) , .ZN( u1_u15_u2_n186 ) );
  OR4_X1 u1_u15_u2_U94 (.ZN( u1_out15_6 ) , .A4( u1_u15_u2_n161 ) , .A3( u1_u15_u2_n162 ) , .A2( u1_u15_u2_n163 ) , .A1( u1_u15_u2_n164 ) );
  OR3_X1 u1_u15_u2_U95 (.A2( u1_u15_u2_n159 ) , .A1( u1_u15_u2_n160 ) , .ZN( u1_u15_u2_n161 ) , .A3( u1_u15_u2_n183 ) );
  AOI21_X1 u1_u15_u2_U96 (.B2( u1_u15_u2_n154 ) , .B1( u1_u15_u2_n155 ) , .ZN( u1_u15_u2_n159 ) , .A( u1_u15_u2_n167 ) );
  NAND3_X1 u1_u15_u2_U97 (.A2( u1_u15_u2_n117 ) , .A1( u1_u15_u2_n122 ) , .A3( u1_u15_u2_n123 ) , .ZN( u1_u15_u2_n134 ) );
  NAND3_X1 u1_u15_u2_U98 (.ZN( u1_u15_u2_n110 ) , .A2( u1_u15_u2_n131 ) , .A3( u1_u15_u2_n139 ) , .A1( u1_u15_u2_n154 ) );
  NAND3_X1 u1_u15_u2_U99 (.A2( u1_u15_u2_n100 ) , .ZN( u1_u15_u2_n101 ) , .A1( u1_u15_u2_n104 ) , .A3( u1_u15_u2_n114 ) );
  INV_X1 u1_u15_u5_U10 (.A( u1_u15_u5_n121 ) , .ZN( u1_u15_u5_n177 ) );
  AOI222_X1 u1_u15_u5_U100 (.ZN( u1_u15_u5_n113 ) , .A1( u1_u15_u5_n131 ) , .C1( u1_u15_u5_n148 ) , .B2( u1_u15_u5_n174 ) , .C2( u1_u15_u5_n178 ) , .A2( u1_u15_u5_n179 ) , .B1( u1_u15_u5_n99 ) );
  NAND4_X1 u1_u15_u5_U101 (.ZN( u1_out15_29 ) , .A4( u1_u15_u5_n129 ) , .A3( u1_u15_u5_n130 ) , .A2( u1_u15_u5_n168 ) , .A1( u1_u15_u5_n196 ) );
  AOI221_X1 u1_u15_u5_U102 (.A( u1_u15_u5_n128 ) , .ZN( u1_u15_u5_n129 ) , .C2( u1_u15_u5_n132 ) , .B2( u1_u15_u5_n159 ) , .B1( u1_u15_u5_n176 ) , .C1( u1_u15_u5_n184 ) );
  AOI222_X1 u1_u15_u5_U103 (.ZN( u1_u15_u5_n130 ) , .A2( u1_u15_u5_n146 ) , .B1( u1_u15_u5_n147 ) , .C2( u1_u15_u5_n175 ) , .B2( u1_u15_u5_n179 ) , .A1( u1_u15_u5_n188 ) , .C1( u1_u15_u5_n194 ) );
  NAND3_X1 u1_u15_u5_U104 (.A2( u1_u15_u5_n154 ) , .A3( u1_u15_u5_n158 ) , .A1( u1_u15_u5_n161 ) , .ZN( u1_u15_u5_n99 ) );
  NOR2_X1 u1_u15_u5_U11 (.ZN( u1_u15_u5_n160 ) , .A2( u1_u15_u5_n173 ) , .A1( u1_u15_u5_n177 ) );
  INV_X1 u1_u15_u5_U12 (.A( u1_u15_u5_n150 ) , .ZN( u1_u15_u5_n174 ) );
  AOI21_X1 u1_u15_u5_U13 (.A( u1_u15_u5_n160 ) , .B2( u1_u15_u5_n161 ) , .ZN( u1_u15_u5_n162 ) , .B1( u1_u15_u5_n192 ) );
  INV_X1 u1_u15_u5_U14 (.A( u1_u15_u5_n159 ) , .ZN( u1_u15_u5_n192 ) );
  AOI21_X1 u1_u15_u5_U15 (.A( u1_u15_u5_n156 ) , .B2( u1_u15_u5_n157 ) , .B1( u1_u15_u5_n158 ) , .ZN( u1_u15_u5_n163 ) );
  AOI21_X1 u1_u15_u5_U16 (.B2( u1_u15_u5_n139 ) , .B1( u1_u15_u5_n140 ) , .ZN( u1_u15_u5_n141 ) , .A( u1_u15_u5_n150 ) );
  OAI21_X1 u1_u15_u5_U17 (.A( u1_u15_u5_n133 ) , .B2( u1_u15_u5_n134 ) , .B1( u1_u15_u5_n135 ) , .ZN( u1_u15_u5_n142 ) );
  OAI21_X1 u1_u15_u5_U18 (.ZN( u1_u15_u5_n133 ) , .B2( u1_u15_u5_n147 ) , .A( u1_u15_u5_n173 ) , .B1( u1_u15_u5_n188 ) );
  NAND2_X1 u1_u15_u5_U19 (.A2( u1_u15_u5_n119 ) , .A1( u1_u15_u5_n123 ) , .ZN( u1_u15_u5_n137 ) );
  INV_X1 u1_u15_u5_U20 (.A( u1_u15_u5_n155 ) , .ZN( u1_u15_u5_n194 ) );
  NAND2_X1 u1_u15_u5_U21 (.A1( u1_u15_u5_n121 ) , .ZN( u1_u15_u5_n132 ) , .A2( u1_u15_u5_n172 ) );
  NAND2_X1 u1_u15_u5_U22 (.A2( u1_u15_u5_n122 ) , .ZN( u1_u15_u5_n136 ) , .A1( u1_u15_u5_n154 ) );
  NAND2_X1 u1_u15_u5_U23 (.A2( u1_u15_u5_n119 ) , .A1( u1_u15_u5_n120 ) , .ZN( u1_u15_u5_n159 ) );
  INV_X1 u1_u15_u5_U24 (.A( u1_u15_u5_n156 ) , .ZN( u1_u15_u5_n175 ) );
  INV_X1 u1_u15_u5_U25 (.A( u1_u15_u5_n158 ) , .ZN( u1_u15_u5_n188 ) );
  INV_X1 u1_u15_u5_U26 (.A( u1_u15_u5_n152 ) , .ZN( u1_u15_u5_n179 ) );
  INV_X1 u1_u15_u5_U27 (.A( u1_u15_u5_n140 ) , .ZN( u1_u15_u5_n182 ) );
  INV_X1 u1_u15_u5_U28 (.A( u1_u15_u5_n151 ) , .ZN( u1_u15_u5_n183 ) );
  INV_X1 u1_u15_u5_U29 (.A( u1_u15_u5_n123 ) , .ZN( u1_u15_u5_n185 ) );
  NOR2_X1 u1_u15_u5_U3 (.ZN( u1_u15_u5_n134 ) , .A1( u1_u15_u5_n183 ) , .A2( u1_u15_u5_n190 ) );
  INV_X1 u1_u15_u5_U30 (.A( u1_u15_u5_n161 ) , .ZN( u1_u15_u5_n184 ) );
  INV_X1 u1_u15_u5_U31 (.A( u1_u15_u5_n139 ) , .ZN( u1_u15_u5_n189 ) );
  INV_X1 u1_u15_u5_U32 (.A( u1_u15_u5_n157 ) , .ZN( u1_u15_u5_n190 ) );
  INV_X1 u1_u15_u5_U33 (.A( u1_u15_u5_n120 ) , .ZN( u1_u15_u5_n193 ) );
  NAND2_X1 u1_u15_u5_U34 (.ZN( u1_u15_u5_n111 ) , .A1( u1_u15_u5_n140 ) , .A2( u1_u15_u5_n155 ) );
  NOR2_X1 u1_u15_u5_U35 (.ZN( u1_u15_u5_n100 ) , .A1( u1_u15_u5_n170 ) , .A2( u1_u15_u5_n180 ) );
  INV_X1 u1_u15_u5_U36 (.A( u1_u15_u5_n117 ) , .ZN( u1_u15_u5_n196 ) );
  OAI221_X1 u1_u15_u5_U37 (.A( u1_u15_u5_n116 ) , .ZN( u1_u15_u5_n117 ) , .B2( u1_u15_u5_n119 ) , .C1( u1_u15_u5_n153 ) , .C2( u1_u15_u5_n158 ) , .B1( u1_u15_u5_n172 ) );
  AOI222_X1 u1_u15_u5_U38 (.ZN( u1_u15_u5_n116 ) , .B2( u1_u15_u5_n145 ) , .C1( u1_u15_u5_n148 ) , .A2( u1_u15_u5_n174 ) , .C2( u1_u15_u5_n177 ) , .B1( u1_u15_u5_n187 ) , .A1( u1_u15_u5_n193 ) );
  INV_X1 u1_u15_u5_U39 (.A( u1_u15_u5_n115 ) , .ZN( u1_u15_u5_n187 ) );
  INV_X1 u1_u15_u5_U4 (.A( u1_u15_u5_n138 ) , .ZN( u1_u15_u5_n191 ) );
  AOI22_X1 u1_u15_u5_U40 (.B2( u1_u15_u5_n131 ) , .A2( u1_u15_u5_n146 ) , .ZN( u1_u15_u5_n169 ) , .B1( u1_u15_u5_n174 ) , .A1( u1_u15_u5_n185 ) );
  NOR2_X1 u1_u15_u5_U41 (.A1( u1_u15_u5_n146 ) , .ZN( u1_u15_u5_n150 ) , .A2( u1_u15_u5_n173 ) );
  AOI21_X1 u1_u15_u5_U42 (.A( u1_u15_u5_n118 ) , .B2( u1_u15_u5_n145 ) , .ZN( u1_u15_u5_n168 ) , .B1( u1_u15_u5_n186 ) );
  INV_X1 u1_u15_u5_U43 (.A( u1_u15_u5_n122 ) , .ZN( u1_u15_u5_n186 ) );
  NOR2_X1 u1_u15_u5_U44 (.A1( u1_u15_u5_n146 ) , .ZN( u1_u15_u5_n152 ) , .A2( u1_u15_u5_n176 ) );
  NOR2_X1 u1_u15_u5_U45 (.A1( u1_u15_u5_n115 ) , .ZN( u1_u15_u5_n118 ) , .A2( u1_u15_u5_n153 ) );
  NOR2_X1 u1_u15_u5_U46 (.A2( u1_u15_u5_n145 ) , .ZN( u1_u15_u5_n156 ) , .A1( u1_u15_u5_n174 ) );
  NOR2_X1 u1_u15_u5_U47 (.ZN( u1_u15_u5_n121 ) , .A2( u1_u15_u5_n145 ) , .A1( u1_u15_u5_n176 ) );
  AOI22_X1 u1_u15_u5_U48 (.ZN( u1_u15_u5_n114 ) , .A2( u1_u15_u5_n137 ) , .A1( u1_u15_u5_n145 ) , .B2( u1_u15_u5_n175 ) , .B1( u1_u15_u5_n193 ) );
  OAI211_X1 u1_u15_u5_U49 (.B( u1_u15_u5_n124 ) , .A( u1_u15_u5_n125 ) , .C2( u1_u15_u5_n126 ) , .C1( u1_u15_u5_n127 ) , .ZN( u1_u15_u5_n128 ) );
  OAI21_X1 u1_u15_u5_U5 (.B2( u1_u15_u5_n136 ) , .B1( u1_u15_u5_n137 ) , .ZN( u1_u15_u5_n138 ) , .A( u1_u15_u5_n177 ) );
  NOR3_X1 u1_u15_u5_U50 (.ZN( u1_u15_u5_n127 ) , .A1( u1_u15_u5_n136 ) , .A3( u1_u15_u5_n148 ) , .A2( u1_u15_u5_n182 ) );
  OAI21_X1 u1_u15_u5_U51 (.ZN( u1_u15_u5_n124 ) , .A( u1_u15_u5_n177 ) , .B2( u1_u15_u5_n183 ) , .B1( u1_u15_u5_n189 ) );
  OAI21_X1 u1_u15_u5_U52 (.ZN( u1_u15_u5_n125 ) , .A( u1_u15_u5_n174 ) , .B2( u1_u15_u5_n185 ) , .B1( u1_u15_u5_n190 ) );
  AOI21_X1 u1_u15_u5_U53 (.A( u1_u15_u5_n153 ) , .B2( u1_u15_u5_n154 ) , .B1( u1_u15_u5_n155 ) , .ZN( u1_u15_u5_n164 ) );
  AOI21_X1 u1_u15_u5_U54 (.ZN( u1_u15_u5_n110 ) , .B1( u1_u15_u5_n122 ) , .B2( u1_u15_u5_n139 ) , .A( u1_u15_u5_n153 ) );
  INV_X1 u1_u15_u5_U55 (.A( u1_u15_u5_n153 ) , .ZN( u1_u15_u5_n176 ) );
  INV_X1 u1_u15_u5_U56 (.A( u1_u15_u5_n126 ) , .ZN( u1_u15_u5_n173 ) );
  AND2_X1 u1_u15_u5_U57 (.A2( u1_u15_u5_n104 ) , .A1( u1_u15_u5_n107 ) , .ZN( u1_u15_u5_n147 ) );
  AND2_X1 u1_u15_u5_U58 (.A2( u1_u15_u5_n104 ) , .A1( u1_u15_u5_n108 ) , .ZN( u1_u15_u5_n148 ) );
  NAND2_X1 u1_u15_u5_U59 (.A1( u1_u15_u5_n105 ) , .A2( u1_u15_u5_n106 ) , .ZN( u1_u15_u5_n158 ) );
  INV_X1 u1_u15_u5_U6 (.A( u1_u15_u5_n135 ) , .ZN( u1_u15_u5_n178 ) );
  NAND2_X1 u1_u15_u5_U60 (.A2( u1_u15_u5_n108 ) , .A1( u1_u15_u5_n109 ) , .ZN( u1_u15_u5_n139 ) );
  NAND2_X1 u1_u15_u5_U61 (.A1( u1_u15_u5_n106 ) , .A2( u1_u15_u5_n108 ) , .ZN( u1_u15_u5_n119 ) );
  NAND2_X1 u1_u15_u5_U62 (.A2( u1_u15_u5_n103 ) , .A1( u1_u15_u5_n105 ) , .ZN( u1_u15_u5_n140 ) );
  NAND2_X1 u1_u15_u5_U63 (.A2( u1_u15_u5_n104 ) , .A1( u1_u15_u5_n105 ) , .ZN( u1_u15_u5_n155 ) );
  NAND2_X1 u1_u15_u5_U64 (.A2( u1_u15_u5_n106 ) , .A1( u1_u15_u5_n107 ) , .ZN( u1_u15_u5_n122 ) );
  NAND2_X1 u1_u15_u5_U65 (.A2( u1_u15_u5_n100 ) , .A1( u1_u15_u5_n106 ) , .ZN( u1_u15_u5_n115 ) );
  NAND2_X1 u1_u15_u5_U66 (.A2( u1_u15_u5_n100 ) , .A1( u1_u15_u5_n103 ) , .ZN( u1_u15_u5_n161 ) );
  NAND2_X1 u1_u15_u5_U67 (.A1( u1_u15_u5_n105 ) , .A2( u1_u15_u5_n109 ) , .ZN( u1_u15_u5_n154 ) );
  INV_X1 u1_u15_u5_U68 (.A( u1_u15_u5_n146 ) , .ZN( u1_u15_u5_n172 ) );
  NAND2_X1 u1_u15_u5_U69 (.A1( u1_u15_u5_n103 ) , .A2( u1_u15_u5_n108 ) , .ZN( u1_u15_u5_n123 ) );
  OAI22_X1 u1_u15_u5_U7 (.B2( u1_u15_u5_n149 ) , .B1( u1_u15_u5_n150 ) , .A2( u1_u15_u5_n151 ) , .A1( u1_u15_u5_n152 ) , .ZN( u1_u15_u5_n165 ) );
  NAND2_X1 u1_u15_u5_U70 (.A2( u1_u15_u5_n103 ) , .A1( u1_u15_u5_n107 ) , .ZN( u1_u15_u5_n151 ) );
  NAND2_X1 u1_u15_u5_U71 (.A2( u1_u15_u5_n107 ) , .A1( u1_u15_u5_n109 ) , .ZN( u1_u15_u5_n120 ) );
  NAND2_X1 u1_u15_u5_U72 (.A2( u1_u15_u5_n100 ) , .A1( u1_u15_u5_n109 ) , .ZN( u1_u15_u5_n157 ) );
  AND2_X1 u1_u15_u5_U73 (.A2( u1_u15_u5_n100 ) , .A1( u1_u15_u5_n104 ) , .ZN( u1_u15_u5_n131 ) );
  INV_X1 u1_u15_u5_U74 (.A( u1_u15_u5_n102 ) , .ZN( u1_u15_u5_n195 ) );
  OAI221_X1 u1_u15_u5_U75 (.A( u1_u15_u5_n101 ) , .ZN( u1_u15_u5_n102 ) , .C2( u1_u15_u5_n115 ) , .C1( u1_u15_u5_n126 ) , .B1( u1_u15_u5_n134 ) , .B2( u1_u15_u5_n160 ) );
  OAI21_X1 u1_u15_u5_U76 (.ZN( u1_u15_u5_n101 ) , .B1( u1_u15_u5_n137 ) , .A( u1_u15_u5_n146 ) , .B2( u1_u15_u5_n147 ) );
  NOR2_X1 u1_u15_u5_U77 (.A2( u1_u15_X_34 ) , .A1( u1_u15_X_35 ) , .ZN( u1_u15_u5_n145 ) );
  NOR2_X1 u1_u15_u5_U78 (.A2( u1_u15_X_34 ) , .ZN( u1_u15_u5_n146 ) , .A1( u1_u15_u5_n171 ) );
  NOR2_X1 u1_u15_u5_U79 (.A2( u1_u15_X_31 ) , .A1( u1_u15_X_32 ) , .ZN( u1_u15_u5_n103 ) );
  NOR3_X1 u1_u15_u5_U8 (.A2( u1_u15_u5_n147 ) , .A1( u1_u15_u5_n148 ) , .ZN( u1_u15_u5_n149 ) , .A3( u1_u15_u5_n194 ) );
  NOR2_X1 u1_u15_u5_U80 (.A2( u1_u15_X_36 ) , .ZN( u1_u15_u5_n105 ) , .A1( u1_u15_u5_n180 ) );
  NOR2_X1 u1_u15_u5_U81 (.A2( u1_u15_X_33 ) , .ZN( u1_u15_u5_n108 ) , .A1( u1_u15_u5_n170 ) );
  NOR2_X1 u1_u15_u5_U82 (.A2( u1_u15_X_33 ) , .A1( u1_u15_X_36 ) , .ZN( u1_u15_u5_n107 ) );
  NOR2_X1 u1_u15_u5_U83 (.A2( u1_u15_X_31 ) , .ZN( u1_u15_u5_n104 ) , .A1( u1_u15_u5_n181 ) );
  NAND2_X1 u1_u15_u5_U84 (.A2( u1_u15_X_34 ) , .A1( u1_u15_X_35 ) , .ZN( u1_u15_u5_n153 ) );
  NAND2_X1 u1_u15_u5_U85 (.A1( u1_u15_X_34 ) , .ZN( u1_u15_u5_n126 ) , .A2( u1_u15_u5_n171 ) );
  AND2_X1 u1_u15_u5_U86 (.A1( u1_u15_X_31 ) , .A2( u1_u15_X_32 ) , .ZN( u1_u15_u5_n106 ) );
  AND2_X1 u1_u15_u5_U87 (.A1( u1_u15_X_31 ) , .ZN( u1_u15_u5_n109 ) , .A2( u1_u15_u5_n181 ) );
  INV_X1 u1_u15_u5_U88 (.A( u1_u15_X_33 ) , .ZN( u1_u15_u5_n180 ) );
  INV_X1 u1_u15_u5_U89 (.A( u1_u15_X_35 ) , .ZN( u1_u15_u5_n171 ) );
  NOR2_X1 u1_u15_u5_U9 (.ZN( u1_u15_u5_n135 ) , .A1( u1_u15_u5_n173 ) , .A2( u1_u15_u5_n176 ) );
  INV_X1 u1_u15_u5_U90 (.A( u1_u15_X_36 ) , .ZN( u1_u15_u5_n170 ) );
  INV_X1 u1_u15_u5_U91 (.A( u1_u15_X_32 ) , .ZN( u1_u15_u5_n181 ) );
  NAND4_X1 u1_u15_u5_U92 (.ZN( u1_out15_19 ) , .A4( u1_u15_u5_n166 ) , .A3( u1_u15_u5_n167 ) , .A2( u1_u15_u5_n168 ) , .A1( u1_u15_u5_n169 ) );
  AOI22_X1 u1_u15_u5_U93 (.B2( u1_u15_u5_n145 ) , .A2( u1_u15_u5_n146 ) , .ZN( u1_u15_u5_n167 ) , .B1( u1_u15_u5_n182 ) , .A1( u1_u15_u5_n189 ) );
  NOR4_X1 u1_u15_u5_U94 (.A4( u1_u15_u5_n162 ) , .A3( u1_u15_u5_n163 ) , .A2( u1_u15_u5_n164 ) , .A1( u1_u15_u5_n165 ) , .ZN( u1_u15_u5_n166 ) );
  NAND4_X1 u1_u15_u5_U95 (.ZN( u1_out15_11 ) , .A4( u1_u15_u5_n143 ) , .A3( u1_u15_u5_n144 ) , .A2( u1_u15_u5_n169 ) , .A1( u1_u15_u5_n196 ) );
  AOI22_X1 u1_u15_u5_U96 (.A2( u1_u15_u5_n132 ) , .ZN( u1_u15_u5_n144 ) , .B2( u1_u15_u5_n145 ) , .B1( u1_u15_u5_n184 ) , .A1( u1_u15_u5_n194 ) );
  NOR3_X1 u1_u15_u5_U97 (.A3( u1_u15_u5_n141 ) , .A1( u1_u15_u5_n142 ) , .ZN( u1_u15_u5_n143 ) , .A2( u1_u15_u5_n191 ) );
  NAND4_X1 u1_u15_u5_U98 (.ZN( u1_out15_4 ) , .A4( u1_u15_u5_n112 ) , .A2( u1_u15_u5_n113 ) , .A1( u1_u15_u5_n114 ) , .A3( u1_u15_u5_n195 ) );
  AOI211_X1 u1_u15_u5_U99 (.A( u1_u15_u5_n110 ) , .C1( u1_u15_u5_n111 ) , .ZN( u1_u15_u5_n112 ) , .B( u1_u15_u5_n118 ) , .C2( u1_u15_u5_n177 ) );
  XOR2_X1 u1_u1_U1 (.B( u1_K2_9 ) , .A( u1_R0_6 ) , .Z( u1_u1_X_9 ) );
  XOR2_X1 u1_u1_U48 (.B( u1_K2_10 ) , .A( u1_R0_7 ) , .Z( u1_u1_X_10 ) );
  NOR2_X1 u1_u1_u1_U10 (.A1( u1_u1_u1_n112 ) , .A2( u1_u1_u1_n116 ) , .ZN( u1_u1_u1_n118 ) );
  NAND3_X1 u1_u1_u1_U100 (.ZN( u1_u1_u1_n113 ) , .A1( u1_u1_u1_n120 ) , .A3( u1_u1_u1_n133 ) , .A2( u1_u1_u1_n155 ) );
  OAI21_X1 u1_u1_u1_U11 (.ZN( u1_u1_u1_n101 ) , .B1( u1_u1_u1_n141 ) , .A( u1_u1_u1_n146 ) , .B2( u1_u1_u1_n183 ) );
  AOI21_X1 u1_u1_u1_U12 (.B2( u1_u1_u1_n155 ) , .B1( u1_u1_u1_n156 ) , .ZN( u1_u1_u1_n157 ) , .A( u1_u1_u1_n174 ) );
  NAND2_X1 u1_u1_u1_U13 (.ZN( u1_u1_u1_n140 ) , .A2( u1_u1_u1_n150 ) , .A1( u1_u1_u1_n155 ) );
  NAND2_X1 u1_u1_u1_U14 (.A1( u1_u1_u1_n131 ) , .ZN( u1_u1_u1_n147 ) , .A2( u1_u1_u1_n153 ) );
  INV_X1 u1_u1_u1_U15 (.A( u1_u1_u1_n139 ) , .ZN( u1_u1_u1_n174 ) );
  OR4_X1 u1_u1_u1_U16 (.A4( u1_u1_u1_n106 ) , .A3( u1_u1_u1_n107 ) , .ZN( u1_u1_u1_n108 ) , .A1( u1_u1_u1_n117 ) , .A2( u1_u1_u1_n184 ) );
  AOI21_X1 u1_u1_u1_U17 (.ZN( u1_u1_u1_n106 ) , .A( u1_u1_u1_n112 ) , .B1( u1_u1_u1_n154 ) , .B2( u1_u1_u1_n156 ) );
  INV_X1 u1_u1_u1_U18 (.A( u1_u1_u1_n101 ) , .ZN( u1_u1_u1_n184 ) );
  AOI21_X1 u1_u1_u1_U19 (.ZN( u1_u1_u1_n107 ) , .B1( u1_u1_u1_n134 ) , .B2( u1_u1_u1_n149 ) , .A( u1_u1_u1_n174 ) );
  INV_X1 u1_u1_u1_U20 (.A( u1_u1_u1_n112 ) , .ZN( u1_u1_u1_n171 ) );
  NAND2_X1 u1_u1_u1_U21 (.ZN( u1_u1_u1_n141 ) , .A1( u1_u1_u1_n153 ) , .A2( u1_u1_u1_n156 ) );
  AND2_X1 u1_u1_u1_U22 (.A1( u1_u1_u1_n123 ) , .ZN( u1_u1_u1_n134 ) , .A2( u1_u1_u1_n161 ) );
  NAND2_X1 u1_u1_u1_U23 (.A2( u1_u1_u1_n115 ) , .A1( u1_u1_u1_n116 ) , .ZN( u1_u1_u1_n148 ) );
  NAND2_X1 u1_u1_u1_U24 (.A2( u1_u1_u1_n133 ) , .A1( u1_u1_u1_n135 ) , .ZN( u1_u1_u1_n159 ) );
  NAND2_X1 u1_u1_u1_U25 (.A2( u1_u1_u1_n115 ) , .A1( u1_u1_u1_n120 ) , .ZN( u1_u1_u1_n132 ) );
  INV_X1 u1_u1_u1_U26 (.A( u1_u1_u1_n154 ) , .ZN( u1_u1_u1_n178 ) );
  INV_X1 u1_u1_u1_U27 (.A( u1_u1_u1_n151 ) , .ZN( u1_u1_u1_n183 ) );
  AND2_X1 u1_u1_u1_U28 (.A1( u1_u1_u1_n129 ) , .A2( u1_u1_u1_n133 ) , .ZN( u1_u1_u1_n149 ) );
  INV_X1 u1_u1_u1_U29 (.A( u1_u1_u1_n131 ) , .ZN( u1_u1_u1_n180 ) );
  INV_X1 u1_u1_u1_U3 (.A( u1_u1_u1_n159 ) , .ZN( u1_u1_u1_n182 ) );
  AOI221_X1 u1_u1_u1_U30 (.B1( u1_u1_u1_n140 ) , .ZN( u1_u1_u1_n167 ) , .B2( u1_u1_u1_n172 ) , .C2( u1_u1_u1_n175 ) , .C1( u1_u1_u1_n178 ) , .A( u1_u1_u1_n188 ) );
  INV_X1 u1_u1_u1_U31 (.ZN( u1_u1_u1_n188 ) , .A( u1_u1_u1_n97 ) );
  AOI211_X1 u1_u1_u1_U32 (.A( u1_u1_u1_n118 ) , .C1( u1_u1_u1_n132 ) , .C2( u1_u1_u1_n139 ) , .B( u1_u1_u1_n96 ) , .ZN( u1_u1_u1_n97 ) );
  AOI21_X1 u1_u1_u1_U33 (.B2( u1_u1_u1_n121 ) , .B1( u1_u1_u1_n135 ) , .A( u1_u1_u1_n152 ) , .ZN( u1_u1_u1_n96 ) );
  OAI221_X1 u1_u1_u1_U34 (.A( u1_u1_u1_n119 ) , .C2( u1_u1_u1_n129 ) , .ZN( u1_u1_u1_n138 ) , .B2( u1_u1_u1_n152 ) , .C1( u1_u1_u1_n174 ) , .B1( u1_u1_u1_n187 ) );
  INV_X1 u1_u1_u1_U35 (.A( u1_u1_u1_n148 ) , .ZN( u1_u1_u1_n187 ) );
  AOI211_X1 u1_u1_u1_U36 (.B( u1_u1_u1_n117 ) , .A( u1_u1_u1_n118 ) , .ZN( u1_u1_u1_n119 ) , .C2( u1_u1_u1_n146 ) , .C1( u1_u1_u1_n159 ) );
  NOR2_X1 u1_u1_u1_U37 (.A1( u1_u1_u1_n168 ) , .A2( u1_u1_u1_n176 ) , .ZN( u1_u1_u1_n98 ) );
  AOI211_X1 u1_u1_u1_U38 (.B( u1_u1_u1_n162 ) , .A( u1_u1_u1_n163 ) , .C2( u1_u1_u1_n164 ) , .ZN( u1_u1_u1_n165 ) , .C1( u1_u1_u1_n171 ) );
  AOI21_X1 u1_u1_u1_U39 (.A( u1_u1_u1_n160 ) , .B2( u1_u1_u1_n161 ) , .ZN( u1_u1_u1_n162 ) , .B1( u1_u1_u1_n182 ) );
  AOI221_X1 u1_u1_u1_U4 (.A( u1_u1_u1_n138 ) , .C2( u1_u1_u1_n139 ) , .C1( u1_u1_u1_n140 ) , .B2( u1_u1_u1_n141 ) , .ZN( u1_u1_u1_n142 ) , .B1( u1_u1_u1_n175 ) );
  OR2_X1 u1_u1_u1_U40 (.A2( u1_u1_u1_n157 ) , .A1( u1_u1_u1_n158 ) , .ZN( u1_u1_u1_n163 ) );
  OAI21_X1 u1_u1_u1_U41 (.B2( u1_u1_u1_n123 ) , .ZN( u1_u1_u1_n145 ) , .B1( u1_u1_u1_n160 ) , .A( u1_u1_u1_n185 ) );
  INV_X1 u1_u1_u1_U42 (.A( u1_u1_u1_n122 ) , .ZN( u1_u1_u1_n185 ) );
  AOI21_X1 u1_u1_u1_U43 (.B2( u1_u1_u1_n120 ) , .B1( u1_u1_u1_n121 ) , .ZN( u1_u1_u1_n122 ) , .A( u1_u1_u1_n128 ) );
  NAND2_X1 u1_u1_u1_U44 (.A1( u1_u1_u1_n128 ) , .ZN( u1_u1_u1_n146 ) , .A2( u1_u1_u1_n160 ) );
  NAND2_X1 u1_u1_u1_U45 (.A2( u1_u1_u1_n112 ) , .ZN( u1_u1_u1_n139 ) , .A1( u1_u1_u1_n152 ) );
  NAND2_X1 u1_u1_u1_U46 (.A1( u1_u1_u1_n105 ) , .ZN( u1_u1_u1_n156 ) , .A2( u1_u1_u1_n99 ) );
  NOR2_X1 u1_u1_u1_U47 (.ZN( u1_u1_u1_n117 ) , .A1( u1_u1_u1_n121 ) , .A2( u1_u1_u1_n160 ) );
  AOI21_X1 u1_u1_u1_U48 (.A( u1_u1_u1_n128 ) , .B2( u1_u1_u1_n129 ) , .ZN( u1_u1_u1_n130 ) , .B1( u1_u1_u1_n150 ) );
  NAND2_X1 u1_u1_u1_U49 (.ZN( u1_u1_u1_n112 ) , .A1( u1_u1_u1_n169 ) , .A2( u1_u1_u1_n170 ) );
  AOI211_X1 u1_u1_u1_U5 (.ZN( u1_u1_u1_n124 ) , .A( u1_u1_u1_n138 ) , .C2( u1_u1_u1_n139 ) , .B( u1_u1_u1_n145 ) , .C1( u1_u1_u1_n147 ) );
  NAND2_X1 u1_u1_u1_U50 (.ZN( u1_u1_u1_n129 ) , .A2( u1_u1_u1_n95 ) , .A1( u1_u1_u1_n98 ) );
  NAND2_X1 u1_u1_u1_U51 (.A1( u1_u1_u1_n102 ) , .ZN( u1_u1_u1_n154 ) , .A2( u1_u1_u1_n99 ) );
  NAND2_X1 u1_u1_u1_U52 (.A2( u1_u1_u1_n100 ) , .ZN( u1_u1_u1_n135 ) , .A1( u1_u1_u1_n99 ) );
  AOI21_X1 u1_u1_u1_U53 (.A( u1_u1_u1_n152 ) , .B2( u1_u1_u1_n153 ) , .B1( u1_u1_u1_n154 ) , .ZN( u1_u1_u1_n158 ) );
  INV_X1 u1_u1_u1_U54 (.A( u1_u1_u1_n160 ) , .ZN( u1_u1_u1_n175 ) );
  NAND2_X1 u1_u1_u1_U55 (.A1( u1_u1_u1_n100 ) , .ZN( u1_u1_u1_n116 ) , .A2( u1_u1_u1_n95 ) );
  NAND2_X1 u1_u1_u1_U56 (.A1( u1_u1_u1_n102 ) , .ZN( u1_u1_u1_n131 ) , .A2( u1_u1_u1_n95 ) );
  NAND2_X1 u1_u1_u1_U57 (.A2( u1_u1_u1_n104 ) , .ZN( u1_u1_u1_n121 ) , .A1( u1_u1_u1_n98 ) );
  NAND2_X1 u1_u1_u1_U58 (.A1( u1_u1_u1_n103 ) , .ZN( u1_u1_u1_n153 ) , .A2( u1_u1_u1_n98 ) );
  NAND2_X1 u1_u1_u1_U59 (.A2( u1_u1_u1_n104 ) , .A1( u1_u1_u1_n105 ) , .ZN( u1_u1_u1_n133 ) );
  AOI22_X1 u1_u1_u1_U6 (.B2( u1_u1_u1_n113 ) , .A2( u1_u1_u1_n114 ) , .ZN( u1_u1_u1_n125 ) , .A1( u1_u1_u1_n171 ) , .B1( u1_u1_u1_n173 ) );
  NAND2_X1 u1_u1_u1_U60 (.ZN( u1_u1_u1_n150 ) , .A2( u1_u1_u1_n98 ) , .A1( u1_u1_u1_n99 ) );
  NAND2_X1 u1_u1_u1_U61 (.A1( u1_u1_u1_n105 ) , .ZN( u1_u1_u1_n155 ) , .A2( u1_u1_u1_n95 ) );
  OAI21_X1 u1_u1_u1_U62 (.ZN( u1_u1_u1_n109 ) , .B1( u1_u1_u1_n129 ) , .B2( u1_u1_u1_n160 ) , .A( u1_u1_u1_n167 ) );
  NAND2_X1 u1_u1_u1_U63 (.A2( u1_u1_u1_n100 ) , .A1( u1_u1_u1_n103 ) , .ZN( u1_u1_u1_n120 ) );
  NAND2_X1 u1_u1_u1_U64 (.A1( u1_u1_u1_n102 ) , .A2( u1_u1_u1_n104 ) , .ZN( u1_u1_u1_n115 ) );
  NAND2_X1 u1_u1_u1_U65 (.A2( u1_u1_u1_n100 ) , .A1( u1_u1_u1_n104 ) , .ZN( u1_u1_u1_n151 ) );
  NAND2_X1 u1_u1_u1_U66 (.A2( u1_u1_u1_n103 ) , .A1( u1_u1_u1_n105 ) , .ZN( u1_u1_u1_n161 ) );
  INV_X1 u1_u1_u1_U67 (.A( u1_u1_u1_n152 ) , .ZN( u1_u1_u1_n173 ) );
  INV_X1 u1_u1_u1_U68 (.A( u1_u1_u1_n128 ) , .ZN( u1_u1_u1_n172 ) );
  NAND2_X1 u1_u1_u1_U69 (.A2( u1_u1_u1_n102 ) , .A1( u1_u1_u1_n103 ) , .ZN( u1_u1_u1_n123 ) );
  NAND2_X1 u1_u1_u1_U7 (.ZN( u1_u1_u1_n114 ) , .A1( u1_u1_u1_n134 ) , .A2( u1_u1_u1_n156 ) );
  NOR2_X1 u1_u1_u1_U70 (.A2( u1_u1_X_7 ) , .A1( u1_u1_X_8 ) , .ZN( u1_u1_u1_n95 ) );
  NOR2_X1 u1_u1_u1_U71 (.A1( u1_u1_X_12 ) , .A2( u1_u1_X_9 ) , .ZN( u1_u1_u1_n100 ) );
  NOR2_X1 u1_u1_u1_U72 (.A2( u1_u1_X_8 ) , .A1( u1_u1_u1_n177 ) , .ZN( u1_u1_u1_n99 ) );
  NOR2_X1 u1_u1_u1_U73 (.A2( u1_u1_X_12 ) , .ZN( u1_u1_u1_n102 ) , .A1( u1_u1_u1_n176 ) );
  NOR2_X1 u1_u1_u1_U74 (.A2( u1_u1_X_9 ) , .ZN( u1_u1_u1_n105 ) , .A1( u1_u1_u1_n168 ) );
  NAND2_X1 u1_u1_u1_U75 (.A1( u1_u1_X_10 ) , .ZN( u1_u1_u1_n160 ) , .A2( u1_u1_u1_n169 ) );
  NAND2_X1 u1_u1_u1_U76 (.A2( u1_u1_X_10 ) , .A1( u1_u1_X_11 ) , .ZN( u1_u1_u1_n152 ) );
  NAND2_X1 u1_u1_u1_U77 (.A1( u1_u1_X_11 ) , .ZN( u1_u1_u1_n128 ) , .A2( u1_u1_u1_n170 ) );
  AND2_X1 u1_u1_u1_U78 (.A2( u1_u1_X_7 ) , .A1( u1_u1_X_8 ) , .ZN( u1_u1_u1_n104 ) );
  AND2_X1 u1_u1_u1_U79 (.A1( u1_u1_X_8 ) , .ZN( u1_u1_u1_n103 ) , .A2( u1_u1_u1_n177 ) );
  AOI22_X1 u1_u1_u1_U8 (.B2( u1_u1_u1_n136 ) , .A2( u1_u1_u1_n137 ) , .ZN( u1_u1_u1_n143 ) , .A1( u1_u1_u1_n171 ) , .B1( u1_u1_u1_n173 ) );
  INV_X1 u1_u1_u1_U80 (.A( u1_u1_X_10 ) , .ZN( u1_u1_u1_n170 ) );
  INV_X1 u1_u1_u1_U81 (.A( u1_u1_X_9 ) , .ZN( u1_u1_u1_n176 ) );
  INV_X1 u1_u1_u1_U82 (.A( u1_u1_X_11 ) , .ZN( u1_u1_u1_n169 ) );
  INV_X1 u1_u1_u1_U83 (.A( u1_u1_X_12 ) , .ZN( u1_u1_u1_n168 ) );
  INV_X1 u1_u1_u1_U84 (.A( u1_u1_X_7 ) , .ZN( u1_u1_u1_n177 ) );
  NAND4_X1 u1_u1_u1_U85 (.ZN( u1_out1_28 ) , .A4( u1_u1_u1_n124 ) , .A3( u1_u1_u1_n125 ) , .A2( u1_u1_u1_n126 ) , .A1( u1_u1_u1_n127 ) );
  OAI21_X1 u1_u1_u1_U86 (.ZN( u1_u1_u1_n127 ) , .B2( u1_u1_u1_n139 ) , .B1( u1_u1_u1_n175 ) , .A( u1_u1_u1_n183 ) );
  OAI21_X1 u1_u1_u1_U87 (.ZN( u1_u1_u1_n126 ) , .B2( u1_u1_u1_n140 ) , .A( u1_u1_u1_n146 ) , .B1( u1_u1_u1_n178 ) );
  NAND4_X1 u1_u1_u1_U88 (.ZN( u1_out1_18 ) , .A4( u1_u1_u1_n165 ) , .A3( u1_u1_u1_n166 ) , .A1( u1_u1_u1_n167 ) , .A2( u1_u1_u1_n186 ) );
  AOI22_X1 u1_u1_u1_U89 (.B2( u1_u1_u1_n146 ) , .B1( u1_u1_u1_n147 ) , .A2( u1_u1_u1_n148 ) , .ZN( u1_u1_u1_n166 ) , .A1( u1_u1_u1_n172 ) );
  INV_X1 u1_u1_u1_U9 (.A( u1_u1_u1_n147 ) , .ZN( u1_u1_u1_n181 ) );
  INV_X1 u1_u1_u1_U90 (.A( u1_u1_u1_n145 ) , .ZN( u1_u1_u1_n186 ) );
  NAND4_X1 u1_u1_u1_U91 (.ZN( u1_out1_2 ) , .A4( u1_u1_u1_n142 ) , .A3( u1_u1_u1_n143 ) , .A2( u1_u1_u1_n144 ) , .A1( u1_u1_u1_n179 ) );
  INV_X1 u1_u1_u1_U92 (.A( u1_u1_u1_n130 ) , .ZN( u1_u1_u1_n179 ) );
  OAI21_X1 u1_u1_u1_U93 (.B2( u1_u1_u1_n132 ) , .ZN( u1_u1_u1_n144 ) , .A( u1_u1_u1_n146 ) , .B1( u1_u1_u1_n180 ) );
  OR4_X1 u1_u1_u1_U94 (.ZN( u1_out1_13 ) , .A4( u1_u1_u1_n108 ) , .A3( u1_u1_u1_n109 ) , .A2( u1_u1_u1_n110 ) , .A1( u1_u1_u1_n111 ) );
  AOI21_X1 u1_u1_u1_U95 (.ZN( u1_u1_u1_n111 ) , .A( u1_u1_u1_n128 ) , .B2( u1_u1_u1_n131 ) , .B1( u1_u1_u1_n135 ) );
  AOI21_X1 u1_u1_u1_U96 (.ZN( u1_u1_u1_n110 ) , .A( u1_u1_u1_n116 ) , .B1( u1_u1_u1_n152 ) , .B2( u1_u1_u1_n160 ) );
  NAND3_X1 u1_u1_u1_U97 (.A3( u1_u1_u1_n149 ) , .A2( u1_u1_u1_n150 ) , .A1( u1_u1_u1_n151 ) , .ZN( u1_u1_u1_n164 ) );
  NAND3_X1 u1_u1_u1_U98 (.A3( u1_u1_u1_n134 ) , .A2( u1_u1_u1_n135 ) , .ZN( u1_u1_u1_n136 ) , .A1( u1_u1_u1_n151 ) );
  NAND3_X1 u1_u1_u1_U99 (.A1( u1_u1_u1_n133 ) , .ZN( u1_u1_u1_n137 ) , .A2( u1_u1_u1_n154 ) , .A3( u1_u1_u1_n181 ) );
  XOR2_X1 u1_u2_U1 (.B( u1_K3_9 ) , .A( u1_R1_6 ) , .Z( u1_u2_X_9 ) );
  XOR2_X1 u1_u2_U48 (.B( u1_K3_10 ) , .A( u1_R1_7 ) , .Z( u1_u2_X_10 ) );
  NOR2_X1 u1_u2_u1_U10 (.A1( u1_u2_u1_n112 ) , .A2( u1_u2_u1_n116 ) , .ZN( u1_u2_u1_n118 ) );
  NAND3_X1 u1_u2_u1_U100 (.ZN( u1_u2_u1_n113 ) , .A1( u1_u2_u1_n120 ) , .A3( u1_u2_u1_n133 ) , .A2( u1_u2_u1_n155 ) );
  OAI21_X1 u1_u2_u1_U11 (.ZN( u1_u2_u1_n101 ) , .B1( u1_u2_u1_n141 ) , .A( u1_u2_u1_n146 ) , .B2( u1_u2_u1_n183 ) );
  AOI21_X1 u1_u2_u1_U12 (.B2( u1_u2_u1_n155 ) , .B1( u1_u2_u1_n156 ) , .ZN( u1_u2_u1_n157 ) , .A( u1_u2_u1_n174 ) );
  OR4_X1 u1_u2_u1_U13 (.A4( u1_u2_u1_n106 ) , .A3( u1_u2_u1_n107 ) , .ZN( u1_u2_u1_n108 ) , .A1( u1_u2_u1_n117 ) , .A2( u1_u2_u1_n184 ) );
  AOI21_X1 u1_u2_u1_U14 (.ZN( u1_u2_u1_n106 ) , .A( u1_u2_u1_n112 ) , .B1( u1_u2_u1_n154 ) , .B2( u1_u2_u1_n156 ) );
  INV_X1 u1_u2_u1_U15 (.A( u1_u2_u1_n101 ) , .ZN( u1_u2_u1_n184 ) );
  AOI21_X1 u1_u2_u1_U16 (.ZN( u1_u2_u1_n107 ) , .B1( u1_u2_u1_n134 ) , .B2( u1_u2_u1_n149 ) , .A( u1_u2_u1_n174 ) );
  NAND2_X1 u1_u2_u1_U17 (.ZN( u1_u2_u1_n140 ) , .A2( u1_u2_u1_n150 ) , .A1( u1_u2_u1_n155 ) );
  NAND2_X1 u1_u2_u1_U18 (.A1( u1_u2_u1_n131 ) , .ZN( u1_u2_u1_n147 ) , .A2( u1_u2_u1_n153 ) );
  INV_X1 u1_u2_u1_U19 (.A( u1_u2_u1_n139 ) , .ZN( u1_u2_u1_n174 ) );
  INV_X1 u1_u2_u1_U20 (.A( u1_u2_u1_n112 ) , .ZN( u1_u2_u1_n171 ) );
  NAND2_X1 u1_u2_u1_U21 (.ZN( u1_u2_u1_n141 ) , .A1( u1_u2_u1_n153 ) , .A2( u1_u2_u1_n156 ) );
  AND2_X1 u1_u2_u1_U22 (.A1( u1_u2_u1_n123 ) , .ZN( u1_u2_u1_n134 ) , .A2( u1_u2_u1_n161 ) );
  NAND2_X1 u1_u2_u1_U23 (.A2( u1_u2_u1_n115 ) , .A1( u1_u2_u1_n116 ) , .ZN( u1_u2_u1_n148 ) );
  NAND2_X1 u1_u2_u1_U24 (.A2( u1_u2_u1_n133 ) , .A1( u1_u2_u1_n135 ) , .ZN( u1_u2_u1_n159 ) );
  NAND2_X1 u1_u2_u1_U25 (.A2( u1_u2_u1_n115 ) , .A1( u1_u2_u1_n120 ) , .ZN( u1_u2_u1_n132 ) );
  INV_X1 u1_u2_u1_U26 (.A( u1_u2_u1_n154 ) , .ZN( u1_u2_u1_n178 ) );
  INV_X1 u1_u2_u1_U27 (.A( u1_u2_u1_n151 ) , .ZN( u1_u2_u1_n183 ) );
  AND2_X1 u1_u2_u1_U28 (.A1( u1_u2_u1_n129 ) , .A2( u1_u2_u1_n133 ) , .ZN( u1_u2_u1_n149 ) );
  INV_X1 u1_u2_u1_U29 (.A( u1_u2_u1_n131 ) , .ZN( u1_u2_u1_n180 ) );
  INV_X1 u1_u2_u1_U3 (.A( u1_u2_u1_n159 ) , .ZN( u1_u2_u1_n182 ) );
  OAI221_X1 u1_u2_u1_U30 (.A( u1_u2_u1_n119 ) , .C2( u1_u2_u1_n129 ) , .ZN( u1_u2_u1_n138 ) , .B2( u1_u2_u1_n152 ) , .C1( u1_u2_u1_n174 ) , .B1( u1_u2_u1_n187 ) );
  INV_X1 u1_u2_u1_U31 (.A( u1_u2_u1_n148 ) , .ZN( u1_u2_u1_n187 ) );
  AOI211_X1 u1_u2_u1_U32 (.B( u1_u2_u1_n117 ) , .A( u1_u2_u1_n118 ) , .ZN( u1_u2_u1_n119 ) , .C2( u1_u2_u1_n146 ) , .C1( u1_u2_u1_n159 ) );
  NOR2_X1 u1_u2_u1_U33 (.A1( u1_u2_u1_n168 ) , .A2( u1_u2_u1_n176 ) , .ZN( u1_u2_u1_n98 ) );
  AOI211_X1 u1_u2_u1_U34 (.B( u1_u2_u1_n162 ) , .A( u1_u2_u1_n163 ) , .C2( u1_u2_u1_n164 ) , .ZN( u1_u2_u1_n165 ) , .C1( u1_u2_u1_n171 ) );
  AOI21_X1 u1_u2_u1_U35 (.A( u1_u2_u1_n160 ) , .B2( u1_u2_u1_n161 ) , .ZN( u1_u2_u1_n162 ) , .B1( u1_u2_u1_n182 ) );
  OR2_X1 u1_u2_u1_U36 (.A2( u1_u2_u1_n157 ) , .A1( u1_u2_u1_n158 ) , .ZN( u1_u2_u1_n163 ) );
  OAI21_X1 u1_u2_u1_U37 (.B2( u1_u2_u1_n123 ) , .ZN( u1_u2_u1_n145 ) , .B1( u1_u2_u1_n160 ) , .A( u1_u2_u1_n185 ) );
  INV_X1 u1_u2_u1_U38 (.A( u1_u2_u1_n122 ) , .ZN( u1_u2_u1_n185 ) );
  AOI21_X1 u1_u2_u1_U39 (.B2( u1_u2_u1_n120 ) , .B1( u1_u2_u1_n121 ) , .ZN( u1_u2_u1_n122 ) , .A( u1_u2_u1_n128 ) );
  AOI221_X1 u1_u2_u1_U4 (.A( u1_u2_u1_n138 ) , .C2( u1_u2_u1_n139 ) , .C1( u1_u2_u1_n140 ) , .B2( u1_u2_u1_n141 ) , .ZN( u1_u2_u1_n142 ) , .B1( u1_u2_u1_n175 ) );
  NAND2_X1 u1_u2_u1_U40 (.A1( u1_u2_u1_n128 ) , .ZN( u1_u2_u1_n146 ) , .A2( u1_u2_u1_n160 ) );
  NAND2_X1 u1_u2_u1_U41 (.A2( u1_u2_u1_n112 ) , .ZN( u1_u2_u1_n139 ) , .A1( u1_u2_u1_n152 ) );
  NAND2_X1 u1_u2_u1_U42 (.A1( u1_u2_u1_n105 ) , .ZN( u1_u2_u1_n156 ) , .A2( u1_u2_u1_n99 ) );
  AOI221_X1 u1_u2_u1_U43 (.B1( u1_u2_u1_n140 ) , .ZN( u1_u2_u1_n167 ) , .B2( u1_u2_u1_n172 ) , .C2( u1_u2_u1_n175 ) , .C1( u1_u2_u1_n178 ) , .A( u1_u2_u1_n188 ) );
  INV_X1 u1_u2_u1_U44 (.ZN( u1_u2_u1_n188 ) , .A( u1_u2_u1_n97 ) );
  AOI211_X1 u1_u2_u1_U45 (.A( u1_u2_u1_n118 ) , .C1( u1_u2_u1_n132 ) , .C2( u1_u2_u1_n139 ) , .B( u1_u2_u1_n96 ) , .ZN( u1_u2_u1_n97 ) );
  AOI21_X1 u1_u2_u1_U46 (.B2( u1_u2_u1_n121 ) , .B1( u1_u2_u1_n135 ) , .A( u1_u2_u1_n152 ) , .ZN( u1_u2_u1_n96 ) );
  NOR2_X1 u1_u2_u1_U47 (.ZN( u1_u2_u1_n117 ) , .A1( u1_u2_u1_n121 ) , .A2( u1_u2_u1_n160 ) );
  AOI21_X1 u1_u2_u1_U48 (.A( u1_u2_u1_n128 ) , .B2( u1_u2_u1_n129 ) , .ZN( u1_u2_u1_n130 ) , .B1( u1_u2_u1_n150 ) );
  NAND2_X1 u1_u2_u1_U49 (.ZN( u1_u2_u1_n112 ) , .A1( u1_u2_u1_n169 ) , .A2( u1_u2_u1_n170 ) );
  AOI211_X1 u1_u2_u1_U5 (.ZN( u1_u2_u1_n124 ) , .A( u1_u2_u1_n138 ) , .C2( u1_u2_u1_n139 ) , .B( u1_u2_u1_n145 ) , .C1( u1_u2_u1_n147 ) );
  NAND2_X1 u1_u2_u1_U50 (.ZN( u1_u2_u1_n129 ) , .A2( u1_u2_u1_n95 ) , .A1( u1_u2_u1_n98 ) );
  NAND2_X1 u1_u2_u1_U51 (.A1( u1_u2_u1_n102 ) , .ZN( u1_u2_u1_n154 ) , .A2( u1_u2_u1_n99 ) );
  NAND2_X1 u1_u2_u1_U52 (.A2( u1_u2_u1_n100 ) , .ZN( u1_u2_u1_n135 ) , .A1( u1_u2_u1_n99 ) );
  AOI21_X1 u1_u2_u1_U53 (.A( u1_u2_u1_n152 ) , .B2( u1_u2_u1_n153 ) , .B1( u1_u2_u1_n154 ) , .ZN( u1_u2_u1_n158 ) );
  INV_X1 u1_u2_u1_U54 (.A( u1_u2_u1_n160 ) , .ZN( u1_u2_u1_n175 ) );
  NAND2_X1 u1_u2_u1_U55 (.A1( u1_u2_u1_n100 ) , .ZN( u1_u2_u1_n116 ) , .A2( u1_u2_u1_n95 ) );
  NAND2_X1 u1_u2_u1_U56 (.A1( u1_u2_u1_n102 ) , .ZN( u1_u2_u1_n131 ) , .A2( u1_u2_u1_n95 ) );
  NAND2_X1 u1_u2_u1_U57 (.A2( u1_u2_u1_n104 ) , .ZN( u1_u2_u1_n121 ) , .A1( u1_u2_u1_n98 ) );
  NAND2_X1 u1_u2_u1_U58 (.A1( u1_u2_u1_n103 ) , .ZN( u1_u2_u1_n153 ) , .A2( u1_u2_u1_n98 ) );
  NAND2_X1 u1_u2_u1_U59 (.A2( u1_u2_u1_n104 ) , .A1( u1_u2_u1_n105 ) , .ZN( u1_u2_u1_n133 ) );
  AOI22_X1 u1_u2_u1_U6 (.B2( u1_u2_u1_n113 ) , .A2( u1_u2_u1_n114 ) , .ZN( u1_u2_u1_n125 ) , .A1( u1_u2_u1_n171 ) , .B1( u1_u2_u1_n173 ) );
  NAND2_X1 u1_u2_u1_U60 (.ZN( u1_u2_u1_n150 ) , .A2( u1_u2_u1_n98 ) , .A1( u1_u2_u1_n99 ) );
  NAND2_X1 u1_u2_u1_U61 (.A1( u1_u2_u1_n105 ) , .ZN( u1_u2_u1_n155 ) , .A2( u1_u2_u1_n95 ) );
  OAI21_X1 u1_u2_u1_U62 (.ZN( u1_u2_u1_n109 ) , .B1( u1_u2_u1_n129 ) , .B2( u1_u2_u1_n160 ) , .A( u1_u2_u1_n167 ) );
  NAND2_X1 u1_u2_u1_U63 (.A2( u1_u2_u1_n100 ) , .A1( u1_u2_u1_n103 ) , .ZN( u1_u2_u1_n120 ) );
  NAND2_X1 u1_u2_u1_U64 (.A1( u1_u2_u1_n102 ) , .A2( u1_u2_u1_n104 ) , .ZN( u1_u2_u1_n115 ) );
  NAND2_X1 u1_u2_u1_U65 (.A2( u1_u2_u1_n100 ) , .A1( u1_u2_u1_n104 ) , .ZN( u1_u2_u1_n151 ) );
  NAND2_X1 u1_u2_u1_U66 (.A2( u1_u2_u1_n103 ) , .A1( u1_u2_u1_n105 ) , .ZN( u1_u2_u1_n161 ) );
  INV_X1 u1_u2_u1_U67 (.A( u1_u2_u1_n152 ) , .ZN( u1_u2_u1_n173 ) );
  INV_X1 u1_u2_u1_U68 (.A( u1_u2_u1_n128 ) , .ZN( u1_u2_u1_n172 ) );
  NAND2_X1 u1_u2_u1_U69 (.A2( u1_u2_u1_n102 ) , .A1( u1_u2_u1_n103 ) , .ZN( u1_u2_u1_n123 ) );
  NAND2_X1 u1_u2_u1_U7 (.ZN( u1_u2_u1_n114 ) , .A1( u1_u2_u1_n134 ) , .A2( u1_u2_u1_n156 ) );
  NOR2_X1 u1_u2_u1_U70 (.A2( u1_u2_X_7 ) , .A1( u1_u2_X_8 ) , .ZN( u1_u2_u1_n95 ) );
  NOR2_X1 u1_u2_u1_U71 (.A1( u1_u2_X_12 ) , .A2( u1_u2_X_9 ) , .ZN( u1_u2_u1_n100 ) );
  NOR2_X1 u1_u2_u1_U72 (.A2( u1_u2_X_8 ) , .A1( u1_u2_u1_n177 ) , .ZN( u1_u2_u1_n99 ) );
  NOR2_X1 u1_u2_u1_U73 (.A2( u1_u2_X_12 ) , .ZN( u1_u2_u1_n102 ) , .A1( u1_u2_u1_n176 ) );
  NOR2_X1 u1_u2_u1_U74 (.A2( u1_u2_X_9 ) , .ZN( u1_u2_u1_n105 ) , .A1( u1_u2_u1_n168 ) );
  NAND2_X1 u1_u2_u1_U75 (.A1( u1_u2_X_10 ) , .ZN( u1_u2_u1_n160 ) , .A2( u1_u2_u1_n169 ) );
  NAND2_X1 u1_u2_u1_U76 (.A2( u1_u2_X_10 ) , .A1( u1_u2_X_11 ) , .ZN( u1_u2_u1_n152 ) );
  NAND2_X1 u1_u2_u1_U77 (.A1( u1_u2_X_11 ) , .ZN( u1_u2_u1_n128 ) , .A2( u1_u2_u1_n170 ) );
  AND2_X1 u1_u2_u1_U78 (.A2( u1_u2_X_7 ) , .A1( u1_u2_X_8 ) , .ZN( u1_u2_u1_n104 ) );
  AND2_X1 u1_u2_u1_U79 (.A1( u1_u2_X_8 ) , .ZN( u1_u2_u1_n103 ) , .A2( u1_u2_u1_n177 ) );
  AOI22_X1 u1_u2_u1_U8 (.B2( u1_u2_u1_n136 ) , .A2( u1_u2_u1_n137 ) , .ZN( u1_u2_u1_n143 ) , .A1( u1_u2_u1_n171 ) , .B1( u1_u2_u1_n173 ) );
  INV_X1 u1_u2_u1_U80 (.A( u1_u2_X_10 ) , .ZN( u1_u2_u1_n170 ) );
  INV_X1 u1_u2_u1_U81 (.A( u1_u2_X_9 ) , .ZN( u1_u2_u1_n176 ) );
  INV_X1 u1_u2_u1_U82 (.A( u1_u2_X_11 ) , .ZN( u1_u2_u1_n169 ) );
  INV_X1 u1_u2_u1_U83 (.A( u1_u2_X_12 ) , .ZN( u1_u2_u1_n168 ) );
  INV_X1 u1_u2_u1_U84 (.A( u1_u2_X_7 ) , .ZN( u1_u2_u1_n177 ) );
  NAND4_X1 u1_u2_u1_U85 (.ZN( u1_out2_18 ) , .A4( u1_u2_u1_n165 ) , .A3( u1_u2_u1_n166 ) , .A1( u1_u2_u1_n167 ) , .A2( u1_u2_u1_n186 ) );
  AOI22_X1 u1_u2_u1_U86 (.B2( u1_u2_u1_n146 ) , .B1( u1_u2_u1_n147 ) , .A2( u1_u2_u1_n148 ) , .ZN( u1_u2_u1_n166 ) , .A1( u1_u2_u1_n172 ) );
  INV_X1 u1_u2_u1_U87 (.A( u1_u2_u1_n145 ) , .ZN( u1_u2_u1_n186 ) );
  NAND4_X1 u1_u2_u1_U88 (.ZN( u1_out2_2 ) , .A4( u1_u2_u1_n142 ) , .A3( u1_u2_u1_n143 ) , .A2( u1_u2_u1_n144 ) , .A1( u1_u2_u1_n179 ) );
  OAI21_X1 u1_u2_u1_U89 (.B2( u1_u2_u1_n132 ) , .ZN( u1_u2_u1_n144 ) , .A( u1_u2_u1_n146 ) , .B1( u1_u2_u1_n180 ) );
  INV_X1 u1_u2_u1_U9 (.A( u1_u2_u1_n147 ) , .ZN( u1_u2_u1_n181 ) );
  INV_X1 u1_u2_u1_U90 (.A( u1_u2_u1_n130 ) , .ZN( u1_u2_u1_n179 ) );
  NAND4_X1 u1_u2_u1_U91 (.ZN( u1_out2_28 ) , .A4( u1_u2_u1_n124 ) , .A3( u1_u2_u1_n125 ) , .A2( u1_u2_u1_n126 ) , .A1( u1_u2_u1_n127 ) );
  OAI21_X1 u1_u2_u1_U92 (.ZN( u1_u2_u1_n127 ) , .B2( u1_u2_u1_n139 ) , .B1( u1_u2_u1_n175 ) , .A( u1_u2_u1_n183 ) );
  OAI21_X1 u1_u2_u1_U93 (.ZN( u1_u2_u1_n126 ) , .B2( u1_u2_u1_n140 ) , .A( u1_u2_u1_n146 ) , .B1( u1_u2_u1_n178 ) );
  OR4_X1 u1_u2_u1_U94 (.ZN( u1_out2_13 ) , .A4( u1_u2_u1_n108 ) , .A3( u1_u2_u1_n109 ) , .A2( u1_u2_u1_n110 ) , .A1( u1_u2_u1_n111 ) );
  AOI21_X1 u1_u2_u1_U95 (.ZN( u1_u2_u1_n111 ) , .A( u1_u2_u1_n128 ) , .B2( u1_u2_u1_n131 ) , .B1( u1_u2_u1_n135 ) );
  AOI21_X1 u1_u2_u1_U96 (.ZN( u1_u2_u1_n110 ) , .A( u1_u2_u1_n116 ) , .B1( u1_u2_u1_n152 ) , .B2( u1_u2_u1_n160 ) );
  NAND3_X1 u1_u2_u1_U97 (.A3( u1_u2_u1_n149 ) , .A2( u1_u2_u1_n150 ) , .A1( u1_u2_u1_n151 ) , .ZN( u1_u2_u1_n164 ) );
  NAND3_X1 u1_u2_u1_U98 (.A3( u1_u2_u1_n134 ) , .A2( u1_u2_u1_n135 ) , .ZN( u1_u2_u1_n136 ) , .A1( u1_u2_u1_n151 ) );
  NAND3_X1 u1_u2_u1_U99 (.A1( u1_u2_u1_n133 ) , .ZN( u1_u2_u1_n137 ) , .A2( u1_u2_u1_n154 ) , .A3( u1_u2_u1_n181 ) );
  XOR2_X1 u1_u3_U1 (.B( u1_K4_9 ) , .A( u1_R2_6 ) , .Z( u1_u3_X_9 ) );
  XOR2_X1 u1_u3_U15 (.B( u1_K4_40 ) , .A( u1_R2_27 ) , .Z( u1_u3_X_40 ) );
  XOR2_X1 u1_u3_U17 (.B( u1_K4_39 ) , .A( u1_R2_26 ) , .Z( u1_u3_X_39 ) );
  XOR2_X1 u1_u3_U48 (.B( u1_K4_10 ) , .A( u1_R2_7 ) , .Z( u1_u3_X_10 ) );
  AOI21_X1 u1_u3_u1_U10 (.B2( u1_u3_u1_n155 ) , .B1( u1_u3_u1_n156 ) , .ZN( u1_u3_u1_n157 ) , .A( u1_u3_u1_n174 ) );
  NAND3_X1 u1_u3_u1_U100 (.ZN( u1_u3_u1_n113 ) , .A1( u1_u3_u1_n120 ) , .A3( u1_u3_u1_n133 ) , .A2( u1_u3_u1_n155 ) );
  NAND2_X1 u1_u3_u1_U11 (.ZN( u1_u3_u1_n140 ) , .A2( u1_u3_u1_n150 ) , .A1( u1_u3_u1_n155 ) );
  NAND2_X1 u1_u3_u1_U12 (.A1( u1_u3_u1_n131 ) , .ZN( u1_u3_u1_n147 ) , .A2( u1_u3_u1_n153 ) );
  INV_X1 u1_u3_u1_U13 (.A( u1_u3_u1_n139 ) , .ZN( u1_u3_u1_n174 ) );
  OR4_X1 u1_u3_u1_U14 (.A4( u1_u3_u1_n106 ) , .A3( u1_u3_u1_n107 ) , .ZN( u1_u3_u1_n108 ) , .A1( u1_u3_u1_n117 ) , .A2( u1_u3_u1_n184 ) );
  AOI21_X1 u1_u3_u1_U15 (.ZN( u1_u3_u1_n106 ) , .A( u1_u3_u1_n112 ) , .B1( u1_u3_u1_n154 ) , .B2( u1_u3_u1_n156 ) );
  INV_X1 u1_u3_u1_U16 (.A( u1_u3_u1_n101 ) , .ZN( u1_u3_u1_n184 ) );
  AOI21_X1 u1_u3_u1_U17 (.ZN( u1_u3_u1_n107 ) , .B1( u1_u3_u1_n134 ) , .B2( u1_u3_u1_n149 ) , .A( u1_u3_u1_n174 ) );
  INV_X1 u1_u3_u1_U18 (.A( u1_u3_u1_n112 ) , .ZN( u1_u3_u1_n171 ) );
  NAND2_X1 u1_u3_u1_U19 (.ZN( u1_u3_u1_n141 ) , .A1( u1_u3_u1_n153 ) , .A2( u1_u3_u1_n156 ) );
  AND2_X1 u1_u3_u1_U20 (.A1( u1_u3_u1_n123 ) , .ZN( u1_u3_u1_n134 ) , .A2( u1_u3_u1_n161 ) );
  NAND2_X1 u1_u3_u1_U21 (.A2( u1_u3_u1_n115 ) , .A1( u1_u3_u1_n116 ) , .ZN( u1_u3_u1_n148 ) );
  NAND2_X1 u1_u3_u1_U22 (.A2( u1_u3_u1_n133 ) , .A1( u1_u3_u1_n135 ) , .ZN( u1_u3_u1_n159 ) );
  NAND2_X1 u1_u3_u1_U23 (.A2( u1_u3_u1_n115 ) , .A1( u1_u3_u1_n120 ) , .ZN( u1_u3_u1_n132 ) );
  INV_X1 u1_u3_u1_U24 (.A( u1_u3_u1_n154 ) , .ZN( u1_u3_u1_n178 ) );
  AOI22_X1 u1_u3_u1_U25 (.B2( u1_u3_u1_n113 ) , .A2( u1_u3_u1_n114 ) , .ZN( u1_u3_u1_n125 ) , .A1( u1_u3_u1_n171 ) , .B1( u1_u3_u1_n173 ) );
  NAND2_X1 u1_u3_u1_U26 (.ZN( u1_u3_u1_n114 ) , .A1( u1_u3_u1_n134 ) , .A2( u1_u3_u1_n156 ) );
  INV_X1 u1_u3_u1_U27 (.A( u1_u3_u1_n151 ) , .ZN( u1_u3_u1_n183 ) );
  AND2_X1 u1_u3_u1_U28 (.A1( u1_u3_u1_n129 ) , .A2( u1_u3_u1_n133 ) , .ZN( u1_u3_u1_n149 ) );
  INV_X1 u1_u3_u1_U29 (.A( u1_u3_u1_n131 ) , .ZN( u1_u3_u1_n180 ) );
  INV_X1 u1_u3_u1_U3 (.A( u1_u3_u1_n159 ) , .ZN( u1_u3_u1_n182 ) );
  AOI221_X1 u1_u3_u1_U30 (.B1( u1_u3_u1_n140 ) , .ZN( u1_u3_u1_n167 ) , .B2( u1_u3_u1_n172 ) , .C2( u1_u3_u1_n175 ) , .C1( u1_u3_u1_n178 ) , .A( u1_u3_u1_n188 ) );
  INV_X1 u1_u3_u1_U31 (.ZN( u1_u3_u1_n188 ) , .A( u1_u3_u1_n97 ) );
  AOI211_X1 u1_u3_u1_U32 (.A( u1_u3_u1_n118 ) , .C1( u1_u3_u1_n132 ) , .C2( u1_u3_u1_n139 ) , .B( u1_u3_u1_n96 ) , .ZN( u1_u3_u1_n97 ) );
  AOI21_X1 u1_u3_u1_U33 (.B2( u1_u3_u1_n121 ) , .B1( u1_u3_u1_n135 ) , .A( u1_u3_u1_n152 ) , .ZN( u1_u3_u1_n96 ) );
  OAI221_X1 u1_u3_u1_U34 (.A( u1_u3_u1_n119 ) , .C2( u1_u3_u1_n129 ) , .ZN( u1_u3_u1_n138 ) , .B2( u1_u3_u1_n152 ) , .C1( u1_u3_u1_n174 ) , .B1( u1_u3_u1_n187 ) );
  INV_X1 u1_u3_u1_U35 (.A( u1_u3_u1_n148 ) , .ZN( u1_u3_u1_n187 ) );
  AOI211_X1 u1_u3_u1_U36 (.B( u1_u3_u1_n117 ) , .A( u1_u3_u1_n118 ) , .ZN( u1_u3_u1_n119 ) , .C2( u1_u3_u1_n146 ) , .C1( u1_u3_u1_n159 ) );
  NOR2_X1 u1_u3_u1_U37 (.A1( u1_u3_u1_n168 ) , .A2( u1_u3_u1_n176 ) , .ZN( u1_u3_u1_n98 ) );
  AOI211_X1 u1_u3_u1_U38 (.B( u1_u3_u1_n162 ) , .A( u1_u3_u1_n163 ) , .C2( u1_u3_u1_n164 ) , .ZN( u1_u3_u1_n165 ) , .C1( u1_u3_u1_n171 ) );
  AOI21_X1 u1_u3_u1_U39 (.A( u1_u3_u1_n160 ) , .B2( u1_u3_u1_n161 ) , .ZN( u1_u3_u1_n162 ) , .B1( u1_u3_u1_n182 ) );
  AOI221_X1 u1_u3_u1_U4 (.A( u1_u3_u1_n138 ) , .C2( u1_u3_u1_n139 ) , .C1( u1_u3_u1_n140 ) , .B2( u1_u3_u1_n141 ) , .ZN( u1_u3_u1_n142 ) , .B1( u1_u3_u1_n175 ) );
  OR2_X1 u1_u3_u1_U40 (.A2( u1_u3_u1_n157 ) , .A1( u1_u3_u1_n158 ) , .ZN( u1_u3_u1_n163 ) );
  NAND2_X1 u1_u3_u1_U41 (.A1( u1_u3_u1_n128 ) , .ZN( u1_u3_u1_n146 ) , .A2( u1_u3_u1_n160 ) );
  NAND2_X1 u1_u3_u1_U42 (.A2( u1_u3_u1_n112 ) , .ZN( u1_u3_u1_n139 ) , .A1( u1_u3_u1_n152 ) );
  NAND2_X1 u1_u3_u1_U43 (.A1( u1_u3_u1_n105 ) , .ZN( u1_u3_u1_n156 ) , .A2( u1_u3_u1_n99 ) );
  NOR2_X1 u1_u3_u1_U44 (.ZN( u1_u3_u1_n117 ) , .A1( u1_u3_u1_n121 ) , .A2( u1_u3_u1_n160 ) );
  OAI21_X1 u1_u3_u1_U45 (.B2( u1_u3_u1_n123 ) , .ZN( u1_u3_u1_n145 ) , .B1( u1_u3_u1_n160 ) , .A( u1_u3_u1_n185 ) );
  INV_X1 u1_u3_u1_U46 (.A( u1_u3_u1_n122 ) , .ZN( u1_u3_u1_n185 ) );
  AOI21_X1 u1_u3_u1_U47 (.B2( u1_u3_u1_n120 ) , .B1( u1_u3_u1_n121 ) , .ZN( u1_u3_u1_n122 ) , .A( u1_u3_u1_n128 ) );
  AOI21_X1 u1_u3_u1_U48 (.A( u1_u3_u1_n128 ) , .B2( u1_u3_u1_n129 ) , .ZN( u1_u3_u1_n130 ) , .B1( u1_u3_u1_n150 ) );
  NAND2_X1 u1_u3_u1_U49 (.ZN( u1_u3_u1_n112 ) , .A1( u1_u3_u1_n169 ) , .A2( u1_u3_u1_n170 ) );
  AOI211_X1 u1_u3_u1_U5 (.ZN( u1_u3_u1_n124 ) , .A( u1_u3_u1_n138 ) , .C2( u1_u3_u1_n139 ) , .B( u1_u3_u1_n145 ) , .C1( u1_u3_u1_n147 ) );
  NAND2_X1 u1_u3_u1_U50 (.ZN( u1_u3_u1_n129 ) , .A2( u1_u3_u1_n95 ) , .A1( u1_u3_u1_n98 ) );
  NAND2_X1 u1_u3_u1_U51 (.A1( u1_u3_u1_n102 ) , .ZN( u1_u3_u1_n154 ) , .A2( u1_u3_u1_n99 ) );
  NAND2_X1 u1_u3_u1_U52 (.A2( u1_u3_u1_n100 ) , .ZN( u1_u3_u1_n135 ) , .A1( u1_u3_u1_n99 ) );
  AOI21_X1 u1_u3_u1_U53 (.A( u1_u3_u1_n152 ) , .B2( u1_u3_u1_n153 ) , .B1( u1_u3_u1_n154 ) , .ZN( u1_u3_u1_n158 ) );
  INV_X1 u1_u3_u1_U54 (.A( u1_u3_u1_n160 ) , .ZN( u1_u3_u1_n175 ) );
  NAND2_X1 u1_u3_u1_U55 (.A1( u1_u3_u1_n100 ) , .ZN( u1_u3_u1_n116 ) , .A2( u1_u3_u1_n95 ) );
  NAND2_X1 u1_u3_u1_U56 (.A1( u1_u3_u1_n102 ) , .ZN( u1_u3_u1_n131 ) , .A2( u1_u3_u1_n95 ) );
  NAND2_X1 u1_u3_u1_U57 (.A2( u1_u3_u1_n104 ) , .ZN( u1_u3_u1_n121 ) , .A1( u1_u3_u1_n98 ) );
  NAND2_X1 u1_u3_u1_U58 (.A1( u1_u3_u1_n103 ) , .ZN( u1_u3_u1_n153 ) , .A2( u1_u3_u1_n98 ) );
  NAND2_X1 u1_u3_u1_U59 (.A2( u1_u3_u1_n104 ) , .A1( u1_u3_u1_n105 ) , .ZN( u1_u3_u1_n133 ) );
  AOI22_X1 u1_u3_u1_U6 (.B2( u1_u3_u1_n136 ) , .A2( u1_u3_u1_n137 ) , .ZN( u1_u3_u1_n143 ) , .A1( u1_u3_u1_n171 ) , .B1( u1_u3_u1_n173 ) );
  NAND2_X1 u1_u3_u1_U60 (.ZN( u1_u3_u1_n150 ) , .A2( u1_u3_u1_n98 ) , .A1( u1_u3_u1_n99 ) );
  NAND2_X1 u1_u3_u1_U61 (.A1( u1_u3_u1_n105 ) , .ZN( u1_u3_u1_n155 ) , .A2( u1_u3_u1_n95 ) );
  OAI21_X1 u1_u3_u1_U62 (.ZN( u1_u3_u1_n109 ) , .B1( u1_u3_u1_n129 ) , .B2( u1_u3_u1_n160 ) , .A( u1_u3_u1_n167 ) );
  NAND2_X1 u1_u3_u1_U63 (.A2( u1_u3_u1_n100 ) , .A1( u1_u3_u1_n103 ) , .ZN( u1_u3_u1_n120 ) );
  NAND2_X1 u1_u3_u1_U64 (.A1( u1_u3_u1_n102 ) , .A2( u1_u3_u1_n104 ) , .ZN( u1_u3_u1_n115 ) );
  NAND2_X1 u1_u3_u1_U65 (.A2( u1_u3_u1_n100 ) , .A1( u1_u3_u1_n104 ) , .ZN( u1_u3_u1_n151 ) );
  NAND2_X1 u1_u3_u1_U66 (.A2( u1_u3_u1_n103 ) , .A1( u1_u3_u1_n105 ) , .ZN( u1_u3_u1_n161 ) );
  INV_X1 u1_u3_u1_U67 (.A( u1_u3_u1_n152 ) , .ZN( u1_u3_u1_n173 ) );
  INV_X1 u1_u3_u1_U68 (.A( u1_u3_u1_n128 ) , .ZN( u1_u3_u1_n172 ) );
  NAND2_X1 u1_u3_u1_U69 (.A2( u1_u3_u1_n102 ) , .A1( u1_u3_u1_n103 ) , .ZN( u1_u3_u1_n123 ) );
  INV_X1 u1_u3_u1_U7 (.A( u1_u3_u1_n147 ) , .ZN( u1_u3_u1_n181 ) );
  NOR2_X1 u1_u3_u1_U70 (.A2( u1_u3_X_7 ) , .A1( u1_u3_X_8 ) , .ZN( u1_u3_u1_n95 ) );
  NOR2_X1 u1_u3_u1_U71 (.A1( u1_u3_X_12 ) , .A2( u1_u3_X_9 ) , .ZN( u1_u3_u1_n100 ) );
  NOR2_X1 u1_u3_u1_U72 (.A2( u1_u3_X_8 ) , .A1( u1_u3_u1_n177 ) , .ZN( u1_u3_u1_n99 ) );
  NOR2_X1 u1_u3_u1_U73 (.A2( u1_u3_X_12 ) , .ZN( u1_u3_u1_n102 ) , .A1( u1_u3_u1_n176 ) );
  NOR2_X1 u1_u3_u1_U74 (.A2( u1_u3_X_9 ) , .ZN( u1_u3_u1_n105 ) , .A1( u1_u3_u1_n168 ) );
  NAND2_X1 u1_u3_u1_U75 (.A1( u1_u3_X_10 ) , .ZN( u1_u3_u1_n160 ) , .A2( u1_u3_u1_n169 ) );
  NAND2_X1 u1_u3_u1_U76 (.A2( u1_u3_X_10 ) , .A1( u1_u3_X_11 ) , .ZN( u1_u3_u1_n152 ) );
  NAND2_X1 u1_u3_u1_U77 (.A1( u1_u3_X_11 ) , .ZN( u1_u3_u1_n128 ) , .A2( u1_u3_u1_n170 ) );
  AND2_X1 u1_u3_u1_U78 (.A2( u1_u3_X_7 ) , .A1( u1_u3_X_8 ) , .ZN( u1_u3_u1_n104 ) );
  AND2_X1 u1_u3_u1_U79 (.A1( u1_u3_X_8 ) , .ZN( u1_u3_u1_n103 ) , .A2( u1_u3_u1_n177 ) );
  NOR2_X1 u1_u3_u1_U8 (.A1( u1_u3_u1_n112 ) , .A2( u1_u3_u1_n116 ) , .ZN( u1_u3_u1_n118 ) );
  INV_X1 u1_u3_u1_U80 (.A( u1_u3_X_10 ) , .ZN( u1_u3_u1_n170 ) );
  INV_X1 u1_u3_u1_U81 (.A( u1_u3_X_9 ) , .ZN( u1_u3_u1_n176 ) );
  INV_X1 u1_u3_u1_U82 (.A( u1_u3_X_11 ) , .ZN( u1_u3_u1_n169 ) );
  INV_X1 u1_u3_u1_U83 (.A( u1_u3_X_12 ) , .ZN( u1_u3_u1_n168 ) );
  INV_X1 u1_u3_u1_U84 (.A( u1_u3_X_7 ) , .ZN( u1_u3_u1_n177 ) );
  NAND4_X1 u1_u3_u1_U85 (.ZN( u1_out3_18 ) , .A4( u1_u3_u1_n165 ) , .A3( u1_u3_u1_n166 ) , .A1( u1_u3_u1_n167 ) , .A2( u1_u3_u1_n186 ) );
  AOI22_X1 u1_u3_u1_U86 (.B2( u1_u3_u1_n146 ) , .B1( u1_u3_u1_n147 ) , .A2( u1_u3_u1_n148 ) , .ZN( u1_u3_u1_n166 ) , .A1( u1_u3_u1_n172 ) );
  INV_X1 u1_u3_u1_U87 (.A( u1_u3_u1_n145 ) , .ZN( u1_u3_u1_n186 ) );
  OR4_X1 u1_u3_u1_U88 (.ZN( u1_out3_13 ) , .A4( u1_u3_u1_n108 ) , .A3( u1_u3_u1_n109 ) , .A2( u1_u3_u1_n110 ) , .A1( u1_u3_u1_n111 ) );
  AOI21_X1 u1_u3_u1_U89 (.ZN( u1_u3_u1_n111 ) , .A( u1_u3_u1_n128 ) , .B2( u1_u3_u1_n131 ) , .B1( u1_u3_u1_n135 ) );
  OAI21_X1 u1_u3_u1_U9 (.ZN( u1_u3_u1_n101 ) , .B1( u1_u3_u1_n141 ) , .A( u1_u3_u1_n146 ) , .B2( u1_u3_u1_n183 ) );
  AOI21_X1 u1_u3_u1_U90 (.ZN( u1_u3_u1_n110 ) , .A( u1_u3_u1_n116 ) , .B1( u1_u3_u1_n152 ) , .B2( u1_u3_u1_n160 ) );
  NAND4_X1 u1_u3_u1_U91 (.ZN( u1_out3_2 ) , .A4( u1_u3_u1_n142 ) , .A3( u1_u3_u1_n143 ) , .A2( u1_u3_u1_n144 ) , .A1( u1_u3_u1_n179 ) );
  INV_X1 u1_u3_u1_U92 (.A( u1_u3_u1_n130 ) , .ZN( u1_u3_u1_n179 ) );
  OAI21_X1 u1_u3_u1_U93 (.B2( u1_u3_u1_n132 ) , .ZN( u1_u3_u1_n144 ) , .A( u1_u3_u1_n146 ) , .B1( u1_u3_u1_n180 ) );
  NAND4_X1 u1_u3_u1_U94 (.ZN( u1_out3_28 ) , .A4( u1_u3_u1_n124 ) , .A3( u1_u3_u1_n125 ) , .A2( u1_u3_u1_n126 ) , .A1( u1_u3_u1_n127 ) );
  OAI21_X1 u1_u3_u1_U95 (.ZN( u1_u3_u1_n127 ) , .B2( u1_u3_u1_n139 ) , .B1( u1_u3_u1_n175 ) , .A( u1_u3_u1_n183 ) );
  OAI21_X1 u1_u3_u1_U96 (.ZN( u1_u3_u1_n126 ) , .B2( u1_u3_u1_n140 ) , .A( u1_u3_u1_n146 ) , .B1( u1_u3_u1_n178 ) );
  NAND3_X1 u1_u3_u1_U97 (.A3( u1_u3_u1_n149 ) , .A2( u1_u3_u1_n150 ) , .A1( u1_u3_u1_n151 ) , .ZN( u1_u3_u1_n164 ) );
  NAND3_X1 u1_u3_u1_U98 (.A3( u1_u3_u1_n134 ) , .A2( u1_u3_u1_n135 ) , .ZN( u1_u3_u1_n136 ) , .A1( u1_u3_u1_n151 ) );
  NAND3_X1 u1_u3_u1_U99 (.A1( u1_u3_u1_n133 ) , .ZN( u1_u3_u1_n137 ) , .A2( u1_u3_u1_n154 ) , .A3( u1_u3_u1_n181 ) );
  INV_X1 u1_u3_u6_U10 (.ZN( u1_u3_u6_n172 ) , .A( u1_u3_u6_n88 ) );
  OAI21_X1 u1_u3_u6_U11 (.A( u1_u3_u6_n159 ) , .B1( u1_u3_u6_n169 ) , .B2( u1_u3_u6_n173 ) , .ZN( u1_u3_u6_n90 ) );
  AOI22_X1 u1_u3_u6_U12 (.A2( u1_u3_u6_n151 ) , .B2( u1_u3_u6_n161 ) , .A1( u1_u3_u6_n167 ) , .B1( u1_u3_u6_n170 ) , .ZN( u1_u3_u6_n89 ) );
  AOI21_X1 u1_u3_u6_U13 (.ZN( u1_u3_u6_n106 ) , .A( u1_u3_u6_n142 ) , .B2( u1_u3_u6_n159 ) , .B1( u1_u3_u6_n164 ) );
  INV_X1 u1_u3_u6_U14 (.A( u1_u3_u6_n155 ) , .ZN( u1_u3_u6_n161 ) );
  INV_X1 u1_u3_u6_U15 (.A( u1_u3_u6_n128 ) , .ZN( u1_u3_u6_n164 ) );
  NAND2_X1 u1_u3_u6_U16 (.ZN( u1_u3_u6_n110 ) , .A1( u1_u3_u6_n122 ) , .A2( u1_u3_u6_n129 ) );
  NAND2_X1 u1_u3_u6_U17 (.ZN( u1_u3_u6_n124 ) , .A2( u1_u3_u6_n146 ) , .A1( u1_u3_u6_n148 ) );
  INV_X1 u1_u3_u6_U18 (.A( u1_u3_u6_n132 ) , .ZN( u1_u3_u6_n171 ) );
  AND2_X1 u1_u3_u6_U19 (.A1( u1_u3_u6_n100 ) , .ZN( u1_u3_u6_n130 ) , .A2( u1_u3_u6_n147 ) );
  INV_X1 u1_u3_u6_U20 (.A( u1_u3_u6_n127 ) , .ZN( u1_u3_u6_n173 ) );
  INV_X1 u1_u3_u6_U21 (.A( u1_u3_u6_n121 ) , .ZN( u1_u3_u6_n167 ) );
  INV_X1 u1_u3_u6_U22 (.A( u1_u3_u6_n100 ) , .ZN( u1_u3_u6_n169 ) );
  INV_X1 u1_u3_u6_U23 (.A( u1_u3_u6_n123 ) , .ZN( u1_u3_u6_n170 ) );
  INV_X1 u1_u3_u6_U24 (.A( u1_u3_u6_n113 ) , .ZN( u1_u3_u6_n168 ) );
  AND2_X1 u1_u3_u6_U25 (.A1( u1_u3_u6_n107 ) , .A2( u1_u3_u6_n119 ) , .ZN( u1_u3_u6_n133 ) );
  AND2_X1 u1_u3_u6_U26 (.A2( u1_u3_u6_n121 ) , .A1( u1_u3_u6_n122 ) , .ZN( u1_u3_u6_n131 ) );
  AND3_X1 u1_u3_u6_U27 (.ZN( u1_u3_u6_n120 ) , .A2( u1_u3_u6_n127 ) , .A1( u1_u3_u6_n132 ) , .A3( u1_u3_u6_n145 ) );
  INV_X1 u1_u3_u6_U28 (.A( u1_u3_u6_n146 ) , .ZN( u1_u3_u6_n163 ) );
  AOI222_X1 u1_u3_u6_U29 (.ZN( u1_u3_u6_n114 ) , .A1( u1_u3_u6_n118 ) , .A2( u1_u3_u6_n126 ) , .B2( u1_u3_u6_n151 ) , .C2( u1_u3_u6_n159 ) , .C1( u1_u3_u6_n168 ) , .B1( u1_u3_u6_n169 ) );
  INV_X1 u1_u3_u6_U3 (.A( u1_u3_u6_n110 ) , .ZN( u1_u3_u6_n166 ) );
  NOR2_X1 u1_u3_u6_U30 (.A1( u1_u3_u6_n162 ) , .A2( u1_u3_u6_n165 ) , .ZN( u1_u3_u6_n98 ) );
  NAND2_X1 u1_u3_u6_U31 (.A1( u1_u3_u6_n144 ) , .ZN( u1_u3_u6_n151 ) , .A2( u1_u3_u6_n158 ) );
  NAND2_X1 u1_u3_u6_U32 (.ZN( u1_u3_u6_n132 ) , .A1( u1_u3_u6_n91 ) , .A2( u1_u3_u6_n97 ) );
  AOI22_X1 u1_u3_u6_U33 (.B2( u1_u3_u6_n110 ) , .B1( u1_u3_u6_n111 ) , .A1( u1_u3_u6_n112 ) , .ZN( u1_u3_u6_n115 ) , .A2( u1_u3_u6_n161 ) );
  NAND4_X1 u1_u3_u6_U34 (.A3( u1_u3_u6_n109 ) , .ZN( u1_u3_u6_n112 ) , .A4( u1_u3_u6_n132 ) , .A2( u1_u3_u6_n147 ) , .A1( u1_u3_u6_n166 ) );
  NOR2_X1 u1_u3_u6_U35 (.ZN( u1_u3_u6_n109 ) , .A1( u1_u3_u6_n170 ) , .A2( u1_u3_u6_n173 ) );
  NOR2_X1 u1_u3_u6_U36 (.A2( u1_u3_u6_n126 ) , .ZN( u1_u3_u6_n155 ) , .A1( u1_u3_u6_n160 ) );
  NAND2_X1 u1_u3_u6_U37 (.ZN( u1_u3_u6_n146 ) , .A2( u1_u3_u6_n94 ) , .A1( u1_u3_u6_n99 ) );
  AOI21_X1 u1_u3_u6_U38 (.A( u1_u3_u6_n144 ) , .B2( u1_u3_u6_n145 ) , .B1( u1_u3_u6_n146 ) , .ZN( u1_u3_u6_n150 ) );
  AOI211_X1 u1_u3_u6_U39 (.B( u1_u3_u6_n134 ) , .A( u1_u3_u6_n135 ) , .C1( u1_u3_u6_n136 ) , .ZN( u1_u3_u6_n137 ) , .C2( u1_u3_u6_n151 ) );
  INV_X1 u1_u3_u6_U4 (.A( u1_u3_u6_n142 ) , .ZN( u1_u3_u6_n174 ) );
  AOI21_X1 u1_u3_u6_U40 (.B2( u1_u3_u6_n132 ) , .B1( u1_u3_u6_n133 ) , .ZN( u1_u3_u6_n134 ) , .A( u1_u3_u6_n158 ) );
  NAND4_X1 u1_u3_u6_U41 (.A4( u1_u3_u6_n127 ) , .A3( u1_u3_u6_n128 ) , .A2( u1_u3_u6_n129 ) , .A1( u1_u3_u6_n130 ) , .ZN( u1_u3_u6_n136 ) );
  AOI21_X1 u1_u3_u6_U42 (.B1( u1_u3_u6_n131 ) , .ZN( u1_u3_u6_n135 ) , .A( u1_u3_u6_n144 ) , .B2( u1_u3_u6_n146 ) );
  INV_X1 u1_u3_u6_U43 (.A( u1_u3_u6_n111 ) , .ZN( u1_u3_u6_n158 ) );
  NAND2_X1 u1_u3_u6_U44 (.ZN( u1_u3_u6_n127 ) , .A1( u1_u3_u6_n91 ) , .A2( u1_u3_u6_n92 ) );
  NAND2_X1 u1_u3_u6_U45 (.ZN( u1_u3_u6_n129 ) , .A2( u1_u3_u6_n95 ) , .A1( u1_u3_u6_n96 ) );
  INV_X1 u1_u3_u6_U46 (.A( u1_u3_u6_n144 ) , .ZN( u1_u3_u6_n159 ) );
  NAND2_X1 u1_u3_u6_U47 (.ZN( u1_u3_u6_n145 ) , .A2( u1_u3_u6_n97 ) , .A1( u1_u3_u6_n98 ) );
  NAND2_X1 u1_u3_u6_U48 (.ZN( u1_u3_u6_n148 ) , .A2( u1_u3_u6_n92 ) , .A1( u1_u3_u6_n94 ) );
  NAND2_X1 u1_u3_u6_U49 (.ZN( u1_u3_u6_n108 ) , .A2( u1_u3_u6_n139 ) , .A1( u1_u3_u6_n144 ) );
  NAND2_X1 u1_u3_u6_U5 (.A2( u1_u3_u6_n143 ) , .ZN( u1_u3_u6_n152 ) , .A1( u1_u3_u6_n166 ) );
  NAND2_X1 u1_u3_u6_U50 (.ZN( u1_u3_u6_n121 ) , .A2( u1_u3_u6_n95 ) , .A1( u1_u3_u6_n97 ) );
  NAND2_X1 u1_u3_u6_U51 (.ZN( u1_u3_u6_n107 ) , .A2( u1_u3_u6_n92 ) , .A1( u1_u3_u6_n95 ) );
  AND2_X1 u1_u3_u6_U52 (.ZN( u1_u3_u6_n118 ) , .A2( u1_u3_u6_n91 ) , .A1( u1_u3_u6_n99 ) );
  NAND2_X1 u1_u3_u6_U53 (.ZN( u1_u3_u6_n147 ) , .A2( u1_u3_u6_n98 ) , .A1( u1_u3_u6_n99 ) );
  NAND2_X1 u1_u3_u6_U54 (.ZN( u1_u3_u6_n128 ) , .A1( u1_u3_u6_n94 ) , .A2( u1_u3_u6_n96 ) );
  NAND2_X1 u1_u3_u6_U55 (.ZN( u1_u3_u6_n119 ) , .A2( u1_u3_u6_n95 ) , .A1( u1_u3_u6_n99 ) );
  NAND2_X1 u1_u3_u6_U56 (.ZN( u1_u3_u6_n123 ) , .A2( u1_u3_u6_n91 ) , .A1( u1_u3_u6_n96 ) );
  NAND2_X1 u1_u3_u6_U57 (.ZN( u1_u3_u6_n100 ) , .A2( u1_u3_u6_n92 ) , .A1( u1_u3_u6_n98 ) );
  NAND2_X1 u1_u3_u6_U58 (.ZN( u1_u3_u6_n122 ) , .A1( u1_u3_u6_n94 ) , .A2( u1_u3_u6_n97 ) );
  INV_X1 u1_u3_u6_U59 (.A( u1_u3_u6_n139 ) , .ZN( u1_u3_u6_n160 ) );
  AOI22_X1 u1_u3_u6_U6 (.B2( u1_u3_u6_n101 ) , .A1( u1_u3_u6_n102 ) , .ZN( u1_u3_u6_n103 ) , .B1( u1_u3_u6_n160 ) , .A2( u1_u3_u6_n161 ) );
  NAND2_X1 u1_u3_u6_U60 (.ZN( u1_u3_u6_n113 ) , .A1( u1_u3_u6_n96 ) , .A2( u1_u3_u6_n98 ) );
  NOR2_X1 u1_u3_u6_U61 (.A2( u1_u3_X_40 ) , .A1( u1_u3_X_41 ) , .ZN( u1_u3_u6_n126 ) );
  NOR2_X1 u1_u3_u6_U62 (.A2( u1_u3_X_39 ) , .A1( u1_u3_X_42 ) , .ZN( u1_u3_u6_n92 ) );
  NOR2_X1 u1_u3_u6_U63 (.A2( u1_u3_X_39 ) , .A1( u1_u3_u6_n156 ) , .ZN( u1_u3_u6_n97 ) );
  NOR2_X1 u1_u3_u6_U64 (.A2( u1_u3_X_38 ) , .A1( u1_u3_u6_n165 ) , .ZN( u1_u3_u6_n95 ) );
  NOR2_X1 u1_u3_u6_U65 (.A2( u1_u3_X_41 ) , .ZN( u1_u3_u6_n111 ) , .A1( u1_u3_u6_n157 ) );
  NOR2_X1 u1_u3_u6_U66 (.A2( u1_u3_X_37 ) , .A1( u1_u3_u6_n162 ) , .ZN( u1_u3_u6_n94 ) );
  NOR2_X1 u1_u3_u6_U67 (.A2( u1_u3_X_37 ) , .A1( u1_u3_X_38 ) , .ZN( u1_u3_u6_n91 ) );
  NAND2_X1 u1_u3_u6_U68 (.A1( u1_u3_X_41 ) , .ZN( u1_u3_u6_n144 ) , .A2( u1_u3_u6_n157 ) );
  NAND2_X1 u1_u3_u6_U69 (.A2( u1_u3_X_40 ) , .A1( u1_u3_X_41 ) , .ZN( u1_u3_u6_n139 ) );
  NOR2_X1 u1_u3_u6_U7 (.A1( u1_u3_u6_n118 ) , .ZN( u1_u3_u6_n143 ) , .A2( u1_u3_u6_n168 ) );
  AND2_X1 u1_u3_u6_U70 (.A1( u1_u3_X_39 ) , .A2( u1_u3_u6_n156 ) , .ZN( u1_u3_u6_n96 ) );
  AND2_X1 u1_u3_u6_U71 (.A1( u1_u3_X_39 ) , .A2( u1_u3_X_42 ) , .ZN( u1_u3_u6_n99 ) );
  INV_X1 u1_u3_u6_U72 (.A( u1_u3_X_40 ) , .ZN( u1_u3_u6_n157 ) );
  INV_X1 u1_u3_u6_U73 (.A( u1_u3_X_37 ) , .ZN( u1_u3_u6_n165 ) );
  INV_X1 u1_u3_u6_U74 (.A( u1_u3_X_38 ) , .ZN( u1_u3_u6_n162 ) );
  INV_X1 u1_u3_u6_U75 (.A( u1_u3_X_42 ) , .ZN( u1_u3_u6_n156 ) );
  NAND4_X1 u1_u3_u6_U76 (.ZN( u1_out3_32 ) , .A4( u1_u3_u6_n103 ) , .A3( u1_u3_u6_n104 ) , .A2( u1_u3_u6_n105 ) , .A1( u1_u3_u6_n106 ) );
  AOI22_X1 u1_u3_u6_U77 (.ZN( u1_u3_u6_n105 ) , .A2( u1_u3_u6_n108 ) , .A1( u1_u3_u6_n118 ) , .B2( u1_u3_u6_n126 ) , .B1( u1_u3_u6_n171 ) );
  AOI22_X1 u1_u3_u6_U78 (.ZN( u1_u3_u6_n104 ) , .A1( u1_u3_u6_n111 ) , .B1( u1_u3_u6_n124 ) , .B2( u1_u3_u6_n151 ) , .A2( u1_u3_u6_n93 ) );
  NAND4_X1 u1_u3_u6_U79 (.ZN( u1_out3_12 ) , .A4( u1_u3_u6_n114 ) , .A3( u1_u3_u6_n115 ) , .A2( u1_u3_u6_n116 ) , .A1( u1_u3_u6_n117 ) );
  AOI21_X1 u1_u3_u6_U8 (.B1( u1_u3_u6_n107 ) , .B2( u1_u3_u6_n132 ) , .A( u1_u3_u6_n158 ) , .ZN( u1_u3_u6_n88 ) );
  OAI22_X1 u1_u3_u6_U80 (.B2( u1_u3_u6_n111 ) , .ZN( u1_u3_u6_n116 ) , .B1( u1_u3_u6_n126 ) , .A2( u1_u3_u6_n164 ) , .A1( u1_u3_u6_n167 ) );
  OAI21_X1 u1_u3_u6_U81 (.A( u1_u3_u6_n108 ) , .ZN( u1_u3_u6_n117 ) , .B2( u1_u3_u6_n141 ) , .B1( u1_u3_u6_n163 ) );
  OAI211_X1 u1_u3_u6_U82 (.ZN( u1_out3_22 ) , .B( u1_u3_u6_n137 ) , .A( u1_u3_u6_n138 ) , .C2( u1_u3_u6_n139 ) , .C1( u1_u3_u6_n140 ) );
  AOI22_X1 u1_u3_u6_U83 (.B1( u1_u3_u6_n124 ) , .A2( u1_u3_u6_n125 ) , .A1( u1_u3_u6_n126 ) , .ZN( u1_u3_u6_n138 ) , .B2( u1_u3_u6_n161 ) );
  AND4_X1 u1_u3_u6_U84 (.A3( u1_u3_u6_n119 ) , .A1( u1_u3_u6_n120 ) , .A4( u1_u3_u6_n129 ) , .ZN( u1_u3_u6_n140 ) , .A2( u1_u3_u6_n143 ) );
  OAI211_X1 u1_u3_u6_U85 (.ZN( u1_out3_7 ) , .B( u1_u3_u6_n153 ) , .C2( u1_u3_u6_n154 ) , .C1( u1_u3_u6_n155 ) , .A( u1_u3_u6_n174 ) );
  NOR3_X1 u1_u3_u6_U86 (.A1( u1_u3_u6_n141 ) , .ZN( u1_u3_u6_n154 ) , .A3( u1_u3_u6_n164 ) , .A2( u1_u3_u6_n171 ) );
  AOI211_X1 u1_u3_u6_U87 (.B( u1_u3_u6_n149 ) , .A( u1_u3_u6_n150 ) , .C2( u1_u3_u6_n151 ) , .C1( u1_u3_u6_n152 ) , .ZN( u1_u3_u6_n153 ) );
  NAND3_X1 u1_u3_u6_U88 (.A2( u1_u3_u6_n123 ) , .ZN( u1_u3_u6_n125 ) , .A1( u1_u3_u6_n130 ) , .A3( u1_u3_u6_n131 ) );
  NAND3_X1 u1_u3_u6_U89 (.A3( u1_u3_u6_n133 ) , .ZN( u1_u3_u6_n141 ) , .A1( u1_u3_u6_n145 ) , .A2( u1_u3_u6_n148 ) );
  AOI21_X1 u1_u3_u6_U9 (.B2( u1_u3_u6_n147 ) , .B1( u1_u3_u6_n148 ) , .ZN( u1_u3_u6_n149 ) , .A( u1_u3_u6_n158 ) );
  NAND3_X1 u1_u3_u6_U90 (.ZN( u1_u3_u6_n101 ) , .A3( u1_u3_u6_n107 ) , .A2( u1_u3_u6_n121 ) , .A1( u1_u3_u6_n127 ) );
  NAND3_X1 u1_u3_u6_U91 (.ZN( u1_u3_u6_n102 ) , .A3( u1_u3_u6_n130 ) , .A2( u1_u3_u6_n145 ) , .A1( u1_u3_u6_n166 ) );
  NAND3_X1 u1_u3_u6_U92 (.A3( u1_u3_u6_n113 ) , .A1( u1_u3_u6_n119 ) , .A2( u1_u3_u6_n123 ) , .ZN( u1_u3_u6_n93 ) );
  NAND3_X1 u1_u3_u6_U93 (.ZN( u1_u3_u6_n142 ) , .A2( u1_u3_u6_n172 ) , .A3( u1_u3_u6_n89 ) , .A1( u1_u3_u6_n90 ) );
  XOR2_X1 u1_u5_U10 (.B( u1_K6_45 ) , .A( u1_R4_30 ) , .Z( u1_u5_X_45 ) );
  XOR2_X1 u1_u5_U9 (.B( u1_K6_46 ) , .A( u1_R4_31 ) , .Z( u1_u5_X_46 ) );
  AND3_X1 u1_u5_u7_U10 (.A3( u1_u5_u7_n110 ) , .A2( u1_u5_u7_n127 ) , .A1( u1_u5_u7_n132 ) , .ZN( u1_u5_u7_n92 ) );
  OAI21_X1 u1_u5_u7_U11 (.A( u1_u5_u7_n161 ) , .B1( u1_u5_u7_n168 ) , .B2( u1_u5_u7_n173 ) , .ZN( u1_u5_u7_n91 ) );
  AOI211_X1 u1_u5_u7_U12 (.A( u1_u5_u7_n117 ) , .ZN( u1_u5_u7_n118 ) , .C2( u1_u5_u7_n126 ) , .C1( u1_u5_u7_n177 ) , .B( u1_u5_u7_n180 ) );
  OAI22_X1 u1_u5_u7_U13 (.B1( u1_u5_u7_n115 ) , .ZN( u1_u5_u7_n117 ) , .A2( u1_u5_u7_n133 ) , .A1( u1_u5_u7_n137 ) , .B2( u1_u5_u7_n162 ) );
  INV_X1 u1_u5_u7_U14 (.A( u1_u5_u7_n116 ) , .ZN( u1_u5_u7_n180 ) );
  NOR3_X1 u1_u5_u7_U15 (.ZN( u1_u5_u7_n115 ) , .A3( u1_u5_u7_n145 ) , .A2( u1_u5_u7_n168 ) , .A1( u1_u5_u7_n169 ) );
  OAI211_X1 u1_u5_u7_U16 (.B( u1_u5_u7_n122 ) , .A( u1_u5_u7_n123 ) , .C2( u1_u5_u7_n124 ) , .ZN( u1_u5_u7_n154 ) , .C1( u1_u5_u7_n162 ) );
  AOI222_X1 u1_u5_u7_U17 (.ZN( u1_u5_u7_n122 ) , .C2( u1_u5_u7_n126 ) , .C1( u1_u5_u7_n145 ) , .B1( u1_u5_u7_n161 ) , .A2( u1_u5_u7_n165 ) , .B2( u1_u5_u7_n170 ) , .A1( u1_u5_u7_n176 ) );
  INV_X1 u1_u5_u7_U18 (.A( u1_u5_u7_n133 ) , .ZN( u1_u5_u7_n176 ) );
  NOR3_X1 u1_u5_u7_U19 (.A2( u1_u5_u7_n134 ) , .A1( u1_u5_u7_n135 ) , .ZN( u1_u5_u7_n136 ) , .A3( u1_u5_u7_n171 ) );
  NOR2_X1 u1_u5_u7_U20 (.A1( u1_u5_u7_n130 ) , .A2( u1_u5_u7_n134 ) , .ZN( u1_u5_u7_n153 ) );
  INV_X1 u1_u5_u7_U21 (.A( u1_u5_u7_n101 ) , .ZN( u1_u5_u7_n165 ) );
  NOR2_X1 u1_u5_u7_U22 (.ZN( u1_u5_u7_n111 ) , .A2( u1_u5_u7_n134 ) , .A1( u1_u5_u7_n169 ) );
  AOI21_X1 u1_u5_u7_U23 (.ZN( u1_u5_u7_n104 ) , .B2( u1_u5_u7_n112 ) , .B1( u1_u5_u7_n127 ) , .A( u1_u5_u7_n164 ) );
  AOI21_X1 u1_u5_u7_U24 (.ZN( u1_u5_u7_n106 ) , .B1( u1_u5_u7_n133 ) , .B2( u1_u5_u7_n146 ) , .A( u1_u5_u7_n162 ) );
  AOI21_X1 u1_u5_u7_U25 (.A( u1_u5_u7_n101 ) , .ZN( u1_u5_u7_n107 ) , .B2( u1_u5_u7_n128 ) , .B1( u1_u5_u7_n175 ) );
  INV_X1 u1_u5_u7_U26 (.A( u1_u5_u7_n138 ) , .ZN( u1_u5_u7_n171 ) );
  INV_X1 u1_u5_u7_U27 (.A( u1_u5_u7_n131 ) , .ZN( u1_u5_u7_n177 ) );
  INV_X1 u1_u5_u7_U28 (.A( u1_u5_u7_n110 ) , .ZN( u1_u5_u7_n174 ) );
  NAND2_X1 u1_u5_u7_U29 (.A1( u1_u5_u7_n129 ) , .A2( u1_u5_u7_n132 ) , .ZN( u1_u5_u7_n149 ) );
  OAI21_X1 u1_u5_u7_U3 (.ZN( u1_u5_u7_n159 ) , .A( u1_u5_u7_n165 ) , .B2( u1_u5_u7_n171 ) , .B1( u1_u5_u7_n174 ) );
  NAND2_X1 u1_u5_u7_U30 (.A1( u1_u5_u7_n113 ) , .A2( u1_u5_u7_n124 ) , .ZN( u1_u5_u7_n130 ) );
  INV_X1 u1_u5_u7_U31 (.A( u1_u5_u7_n112 ) , .ZN( u1_u5_u7_n173 ) );
  INV_X1 u1_u5_u7_U32 (.A( u1_u5_u7_n128 ) , .ZN( u1_u5_u7_n168 ) );
  INV_X1 u1_u5_u7_U33 (.A( u1_u5_u7_n148 ) , .ZN( u1_u5_u7_n169 ) );
  INV_X1 u1_u5_u7_U34 (.A( u1_u5_u7_n127 ) , .ZN( u1_u5_u7_n179 ) );
  NOR2_X1 u1_u5_u7_U35 (.ZN( u1_u5_u7_n101 ) , .A2( u1_u5_u7_n150 ) , .A1( u1_u5_u7_n156 ) );
  AOI211_X1 u1_u5_u7_U36 (.B( u1_u5_u7_n154 ) , .A( u1_u5_u7_n155 ) , .C1( u1_u5_u7_n156 ) , .ZN( u1_u5_u7_n157 ) , .C2( u1_u5_u7_n172 ) );
  INV_X1 u1_u5_u7_U37 (.A( u1_u5_u7_n153 ) , .ZN( u1_u5_u7_n172 ) );
  AOI211_X1 u1_u5_u7_U38 (.B( u1_u5_u7_n139 ) , .A( u1_u5_u7_n140 ) , .C2( u1_u5_u7_n141 ) , .ZN( u1_u5_u7_n142 ) , .C1( u1_u5_u7_n156 ) );
  NAND4_X1 u1_u5_u7_U39 (.A3( u1_u5_u7_n127 ) , .A2( u1_u5_u7_n128 ) , .A1( u1_u5_u7_n129 ) , .ZN( u1_u5_u7_n141 ) , .A4( u1_u5_u7_n147 ) );
  INV_X1 u1_u5_u7_U4 (.A( u1_u5_u7_n111 ) , .ZN( u1_u5_u7_n170 ) );
  AOI21_X1 u1_u5_u7_U40 (.A( u1_u5_u7_n137 ) , .B1( u1_u5_u7_n138 ) , .ZN( u1_u5_u7_n139 ) , .B2( u1_u5_u7_n146 ) );
  OAI22_X1 u1_u5_u7_U41 (.B1( u1_u5_u7_n136 ) , .ZN( u1_u5_u7_n140 ) , .A1( u1_u5_u7_n153 ) , .B2( u1_u5_u7_n162 ) , .A2( u1_u5_u7_n164 ) );
  AOI21_X1 u1_u5_u7_U42 (.ZN( u1_u5_u7_n123 ) , .B1( u1_u5_u7_n165 ) , .B2( u1_u5_u7_n177 ) , .A( u1_u5_u7_n97 ) );
  AOI21_X1 u1_u5_u7_U43 (.B2( u1_u5_u7_n113 ) , .B1( u1_u5_u7_n124 ) , .A( u1_u5_u7_n125 ) , .ZN( u1_u5_u7_n97 ) );
  INV_X1 u1_u5_u7_U44 (.A( u1_u5_u7_n125 ) , .ZN( u1_u5_u7_n161 ) );
  INV_X1 u1_u5_u7_U45 (.A( u1_u5_u7_n152 ) , .ZN( u1_u5_u7_n162 ) );
  AOI22_X1 u1_u5_u7_U46 (.A2( u1_u5_u7_n114 ) , .ZN( u1_u5_u7_n119 ) , .B1( u1_u5_u7_n130 ) , .A1( u1_u5_u7_n156 ) , .B2( u1_u5_u7_n165 ) );
  NAND2_X1 u1_u5_u7_U47 (.A2( u1_u5_u7_n112 ) , .ZN( u1_u5_u7_n114 ) , .A1( u1_u5_u7_n175 ) );
  AND2_X1 u1_u5_u7_U48 (.ZN( u1_u5_u7_n145 ) , .A2( u1_u5_u7_n98 ) , .A1( u1_u5_u7_n99 ) );
  NOR2_X1 u1_u5_u7_U49 (.ZN( u1_u5_u7_n137 ) , .A1( u1_u5_u7_n150 ) , .A2( u1_u5_u7_n161 ) );
  INV_X1 u1_u5_u7_U5 (.A( u1_u5_u7_n149 ) , .ZN( u1_u5_u7_n175 ) );
  AOI21_X1 u1_u5_u7_U50 (.ZN( u1_u5_u7_n105 ) , .B2( u1_u5_u7_n110 ) , .A( u1_u5_u7_n125 ) , .B1( u1_u5_u7_n147 ) );
  NAND2_X1 u1_u5_u7_U51 (.ZN( u1_u5_u7_n146 ) , .A1( u1_u5_u7_n95 ) , .A2( u1_u5_u7_n98 ) );
  NAND2_X1 u1_u5_u7_U52 (.A2( u1_u5_u7_n103 ) , .ZN( u1_u5_u7_n147 ) , .A1( u1_u5_u7_n93 ) );
  NAND2_X1 u1_u5_u7_U53 (.A1( u1_u5_u7_n103 ) , .ZN( u1_u5_u7_n127 ) , .A2( u1_u5_u7_n99 ) );
  OR2_X1 u1_u5_u7_U54 (.ZN( u1_u5_u7_n126 ) , .A2( u1_u5_u7_n152 ) , .A1( u1_u5_u7_n156 ) );
  NAND2_X1 u1_u5_u7_U55 (.A2( u1_u5_u7_n102 ) , .A1( u1_u5_u7_n103 ) , .ZN( u1_u5_u7_n133 ) );
  NAND2_X1 u1_u5_u7_U56 (.ZN( u1_u5_u7_n112 ) , .A2( u1_u5_u7_n96 ) , .A1( u1_u5_u7_n99 ) );
  NAND2_X1 u1_u5_u7_U57 (.A2( u1_u5_u7_n102 ) , .ZN( u1_u5_u7_n128 ) , .A1( u1_u5_u7_n98 ) );
  NAND2_X1 u1_u5_u7_U58 (.A1( u1_u5_u7_n100 ) , .ZN( u1_u5_u7_n113 ) , .A2( u1_u5_u7_n93 ) );
  NAND2_X1 u1_u5_u7_U59 (.A2( u1_u5_u7_n102 ) , .ZN( u1_u5_u7_n124 ) , .A1( u1_u5_u7_n96 ) );
  INV_X1 u1_u5_u7_U6 (.A( u1_u5_u7_n154 ) , .ZN( u1_u5_u7_n178 ) );
  NAND2_X1 u1_u5_u7_U60 (.ZN( u1_u5_u7_n110 ) , .A1( u1_u5_u7_n95 ) , .A2( u1_u5_u7_n96 ) );
  INV_X1 u1_u5_u7_U61 (.A( u1_u5_u7_n150 ) , .ZN( u1_u5_u7_n164 ) );
  AND2_X1 u1_u5_u7_U62 (.ZN( u1_u5_u7_n134 ) , .A1( u1_u5_u7_n93 ) , .A2( u1_u5_u7_n98 ) );
  NAND2_X1 u1_u5_u7_U63 (.A1( u1_u5_u7_n100 ) , .A2( u1_u5_u7_n102 ) , .ZN( u1_u5_u7_n129 ) );
  NAND2_X1 u1_u5_u7_U64 (.A2( u1_u5_u7_n103 ) , .ZN( u1_u5_u7_n131 ) , .A1( u1_u5_u7_n95 ) );
  NAND2_X1 u1_u5_u7_U65 (.A1( u1_u5_u7_n100 ) , .ZN( u1_u5_u7_n138 ) , .A2( u1_u5_u7_n99 ) );
  NAND2_X1 u1_u5_u7_U66 (.ZN( u1_u5_u7_n132 ) , .A1( u1_u5_u7_n93 ) , .A2( u1_u5_u7_n96 ) );
  NAND2_X1 u1_u5_u7_U67 (.A1( u1_u5_u7_n100 ) , .ZN( u1_u5_u7_n148 ) , .A2( u1_u5_u7_n95 ) );
  NOR2_X1 u1_u5_u7_U68 (.A2( u1_u5_X_47 ) , .ZN( u1_u5_u7_n150 ) , .A1( u1_u5_u7_n163 ) );
  NOR2_X1 u1_u5_u7_U69 (.A2( u1_u5_X_43 ) , .A1( u1_u5_X_44 ) , .ZN( u1_u5_u7_n103 ) );
  AOI211_X1 u1_u5_u7_U7 (.ZN( u1_u5_u7_n116 ) , .A( u1_u5_u7_n155 ) , .C1( u1_u5_u7_n161 ) , .C2( u1_u5_u7_n171 ) , .B( u1_u5_u7_n94 ) );
  NOR2_X1 u1_u5_u7_U70 (.A2( u1_u5_X_48 ) , .A1( u1_u5_u7_n166 ) , .ZN( u1_u5_u7_n95 ) );
  NOR2_X1 u1_u5_u7_U71 (.A2( u1_u5_X_45 ) , .A1( u1_u5_X_48 ) , .ZN( u1_u5_u7_n99 ) );
  NOR2_X1 u1_u5_u7_U72 (.A2( u1_u5_X_44 ) , .A1( u1_u5_u7_n167 ) , .ZN( u1_u5_u7_n98 ) );
  NOR2_X1 u1_u5_u7_U73 (.A2( u1_u5_X_46 ) , .A1( u1_u5_X_47 ) , .ZN( u1_u5_u7_n152 ) );
  AND2_X1 u1_u5_u7_U74 (.A1( u1_u5_X_47 ) , .ZN( u1_u5_u7_n156 ) , .A2( u1_u5_u7_n163 ) );
  NAND2_X1 u1_u5_u7_U75 (.A2( u1_u5_X_46 ) , .A1( u1_u5_X_47 ) , .ZN( u1_u5_u7_n125 ) );
  AND2_X1 u1_u5_u7_U76 (.A2( u1_u5_X_45 ) , .A1( u1_u5_X_48 ) , .ZN( u1_u5_u7_n102 ) );
  AND2_X1 u1_u5_u7_U77 (.A2( u1_u5_X_43 ) , .A1( u1_u5_X_44 ) , .ZN( u1_u5_u7_n96 ) );
  AND2_X1 u1_u5_u7_U78 (.A1( u1_u5_X_44 ) , .ZN( u1_u5_u7_n100 ) , .A2( u1_u5_u7_n167 ) );
  AND2_X1 u1_u5_u7_U79 (.A1( u1_u5_X_48 ) , .A2( u1_u5_u7_n166 ) , .ZN( u1_u5_u7_n93 ) );
  OAI222_X1 u1_u5_u7_U8 (.C2( u1_u5_u7_n101 ) , .B2( u1_u5_u7_n111 ) , .A1( u1_u5_u7_n113 ) , .C1( u1_u5_u7_n146 ) , .A2( u1_u5_u7_n162 ) , .B1( u1_u5_u7_n164 ) , .ZN( u1_u5_u7_n94 ) );
  INV_X1 u1_u5_u7_U80 (.A( u1_u5_X_46 ) , .ZN( u1_u5_u7_n163 ) );
  INV_X1 u1_u5_u7_U81 (.A( u1_u5_X_43 ) , .ZN( u1_u5_u7_n167 ) );
  INV_X1 u1_u5_u7_U82 (.A( u1_u5_X_45 ) , .ZN( u1_u5_u7_n166 ) );
  NAND4_X1 u1_u5_u7_U83 (.ZN( u1_out5_5 ) , .A4( u1_u5_u7_n108 ) , .A3( u1_u5_u7_n109 ) , .A1( u1_u5_u7_n116 ) , .A2( u1_u5_u7_n123 ) );
  AOI22_X1 u1_u5_u7_U84 (.ZN( u1_u5_u7_n109 ) , .A2( u1_u5_u7_n126 ) , .B2( u1_u5_u7_n145 ) , .B1( u1_u5_u7_n156 ) , .A1( u1_u5_u7_n171 ) );
  NOR4_X1 u1_u5_u7_U85 (.A4( u1_u5_u7_n104 ) , .A3( u1_u5_u7_n105 ) , .A2( u1_u5_u7_n106 ) , .A1( u1_u5_u7_n107 ) , .ZN( u1_u5_u7_n108 ) );
  NAND4_X1 u1_u5_u7_U86 (.ZN( u1_out5_27 ) , .A4( u1_u5_u7_n118 ) , .A3( u1_u5_u7_n119 ) , .A2( u1_u5_u7_n120 ) , .A1( u1_u5_u7_n121 ) );
  OAI21_X1 u1_u5_u7_U87 (.ZN( u1_u5_u7_n121 ) , .B2( u1_u5_u7_n145 ) , .A( u1_u5_u7_n150 ) , .B1( u1_u5_u7_n174 ) );
  OAI21_X1 u1_u5_u7_U88 (.ZN( u1_u5_u7_n120 ) , .A( u1_u5_u7_n161 ) , .B2( u1_u5_u7_n170 ) , .B1( u1_u5_u7_n179 ) );
  NAND4_X1 u1_u5_u7_U89 (.ZN( u1_out5_21 ) , .A4( u1_u5_u7_n157 ) , .A3( u1_u5_u7_n158 ) , .A2( u1_u5_u7_n159 ) , .A1( u1_u5_u7_n160 ) );
  OAI221_X1 u1_u5_u7_U9 (.C1( u1_u5_u7_n101 ) , .C2( u1_u5_u7_n147 ) , .ZN( u1_u5_u7_n155 ) , .B2( u1_u5_u7_n162 ) , .A( u1_u5_u7_n91 ) , .B1( u1_u5_u7_n92 ) );
  OAI21_X1 u1_u5_u7_U90 (.B1( u1_u5_u7_n145 ) , .ZN( u1_u5_u7_n160 ) , .A( u1_u5_u7_n161 ) , .B2( u1_u5_u7_n177 ) );
  AOI22_X1 u1_u5_u7_U91 (.B2( u1_u5_u7_n149 ) , .B1( u1_u5_u7_n150 ) , .A2( u1_u5_u7_n151 ) , .A1( u1_u5_u7_n152 ) , .ZN( u1_u5_u7_n158 ) );
  NAND4_X1 u1_u5_u7_U92 (.ZN( u1_out5_15 ) , .A4( u1_u5_u7_n142 ) , .A3( u1_u5_u7_n143 ) , .A2( u1_u5_u7_n144 ) , .A1( u1_u5_u7_n178 ) );
  OR2_X1 u1_u5_u7_U93 (.A2( u1_u5_u7_n125 ) , .A1( u1_u5_u7_n129 ) , .ZN( u1_u5_u7_n144 ) );
  AOI22_X1 u1_u5_u7_U94 (.A2( u1_u5_u7_n126 ) , .ZN( u1_u5_u7_n143 ) , .B2( u1_u5_u7_n165 ) , .B1( u1_u5_u7_n173 ) , .A1( u1_u5_u7_n174 ) );
  NAND3_X1 u1_u5_u7_U95 (.A3( u1_u5_u7_n146 ) , .A2( u1_u5_u7_n147 ) , .A1( u1_u5_u7_n148 ) , .ZN( u1_u5_u7_n151 ) );
  NAND3_X1 u1_u5_u7_U96 (.A3( u1_u5_u7_n131 ) , .A2( u1_u5_u7_n132 ) , .A1( u1_u5_u7_n133 ) , .ZN( u1_u5_u7_n135 ) );
  XOR2_X1 u1_u6_U1 (.B( u1_K7_9 ) , .A( u1_R5_6 ) , .Z( u1_u6_X_9 ) );
  XOR2_X1 u1_u6_U10 (.B( u1_K7_45 ) , .A( u1_R5_30 ) , .Z( u1_u6_X_45 ) );
  XOR2_X1 u1_u6_U48 (.B( u1_K7_10 ) , .A( u1_R5_7 ) , .Z( u1_u6_X_10 ) );
  XOR2_X1 u1_u6_U9 (.B( u1_K7_46 ) , .A( u1_R5_31 ) , .Z( u1_u6_X_46 ) );
  NOR2_X1 u1_u6_u1_U10 (.A1( u1_u6_u1_n112 ) , .A2( u1_u6_u1_n116 ) , .ZN( u1_u6_u1_n118 ) );
  NAND3_X1 u1_u6_u1_U100 (.ZN( u1_u6_u1_n113 ) , .A1( u1_u6_u1_n120 ) , .A3( u1_u6_u1_n133 ) , .A2( u1_u6_u1_n155 ) );
  OAI21_X1 u1_u6_u1_U11 (.ZN( u1_u6_u1_n101 ) , .B1( u1_u6_u1_n141 ) , .A( u1_u6_u1_n146 ) , .B2( u1_u6_u1_n183 ) );
  AOI21_X1 u1_u6_u1_U12 (.B2( u1_u6_u1_n155 ) , .B1( u1_u6_u1_n156 ) , .ZN( u1_u6_u1_n157 ) , .A( u1_u6_u1_n174 ) );
  NAND2_X1 u1_u6_u1_U13 (.ZN( u1_u6_u1_n140 ) , .A2( u1_u6_u1_n150 ) , .A1( u1_u6_u1_n155 ) );
  NAND2_X1 u1_u6_u1_U14 (.A1( u1_u6_u1_n131 ) , .ZN( u1_u6_u1_n147 ) , .A2( u1_u6_u1_n153 ) );
  INV_X1 u1_u6_u1_U15 (.A( u1_u6_u1_n139 ) , .ZN( u1_u6_u1_n174 ) );
  OR4_X1 u1_u6_u1_U16 (.A4( u1_u6_u1_n106 ) , .A3( u1_u6_u1_n107 ) , .ZN( u1_u6_u1_n108 ) , .A1( u1_u6_u1_n117 ) , .A2( u1_u6_u1_n184 ) );
  AOI21_X1 u1_u6_u1_U17 (.ZN( u1_u6_u1_n106 ) , .A( u1_u6_u1_n112 ) , .B1( u1_u6_u1_n154 ) , .B2( u1_u6_u1_n156 ) );
  AOI21_X1 u1_u6_u1_U18 (.ZN( u1_u6_u1_n107 ) , .B1( u1_u6_u1_n134 ) , .B2( u1_u6_u1_n149 ) , .A( u1_u6_u1_n174 ) );
  INV_X1 u1_u6_u1_U19 (.A( u1_u6_u1_n101 ) , .ZN( u1_u6_u1_n184 ) );
  INV_X1 u1_u6_u1_U20 (.A( u1_u6_u1_n112 ) , .ZN( u1_u6_u1_n171 ) );
  NAND2_X1 u1_u6_u1_U21 (.ZN( u1_u6_u1_n141 ) , .A1( u1_u6_u1_n153 ) , .A2( u1_u6_u1_n156 ) );
  AND2_X1 u1_u6_u1_U22 (.A1( u1_u6_u1_n123 ) , .ZN( u1_u6_u1_n134 ) , .A2( u1_u6_u1_n161 ) );
  NAND2_X1 u1_u6_u1_U23 (.A2( u1_u6_u1_n115 ) , .A1( u1_u6_u1_n116 ) , .ZN( u1_u6_u1_n148 ) );
  NAND2_X1 u1_u6_u1_U24 (.A2( u1_u6_u1_n133 ) , .A1( u1_u6_u1_n135 ) , .ZN( u1_u6_u1_n159 ) );
  NAND2_X1 u1_u6_u1_U25 (.A2( u1_u6_u1_n115 ) , .A1( u1_u6_u1_n120 ) , .ZN( u1_u6_u1_n132 ) );
  INV_X1 u1_u6_u1_U26 (.A( u1_u6_u1_n154 ) , .ZN( u1_u6_u1_n178 ) );
  INV_X1 u1_u6_u1_U27 (.A( u1_u6_u1_n151 ) , .ZN( u1_u6_u1_n183 ) );
  AND2_X1 u1_u6_u1_U28 (.A1( u1_u6_u1_n129 ) , .A2( u1_u6_u1_n133 ) , .ZN( u1_u6_u1_n149 ) );
  INV_X1 u1_u6_u1_U29 (.A( u1_u6_u1_n131 ) , .ZN( u1_u6_u1_n180 ) );
  INV_X1 u1_u6_u1_U3 (.A( u1_u6_u1_n159 ) , .ZN( u1_u6_u1_n182 ) );
  AOI221_X1 u1_u6_u1_U30 (.B1( u1_u6_u1_n140 ) , .ZN( u1_u6_u1_n167 ) , .B2( u1_u6_u1_n172 ) , .C2( u1_u6_u1_n175 ) , .C1( u1_u6_u1_n178 ) , .A( u1_u6_u1_n188 ) );
  INV_X1 u1_u6_u1_U31 (.ZN( u1_u6_u1_n188 ) , .A( u1_u6_u1_n97 ) );
  AOI211_X1 u1_u6_u1_U32 (.A( u1_u6_u1_n118 ) , .C1( u1_u6_u1_n132 ) , .C2( u1_u6_u1_n139 ) , .B( u1_u6_u1_n96 ) , .ZN( u1_u6_u1_n97 ) );
  AOI21_X1 u1_u6_u1_U33 (.B2( u1_u6_u1_n121 ) , .B1( u1_u6_u1_n135 ) , .A( u1_u6_u1_n152 ) , .ZN( u1_u6_u1_n96 ) );
  OAI221_X1 u1_u6_u1_U34 (.A( u1_u6_u1_n119 ) , .C2( u1_u6_u1_n129 ) , .ZN( u1_u6_u1_n138 ) , .B2( u1_u6_u1_n152 ) , .C1( u1_u6_u1_n174 ) , .B1( u1_u6_u1_n187 ) );
  INV_X1 u1_u6_u1_U35 (.A( u1_u6_u1_n148 ) , .ZN( u1_u6_u1_n187 ) );
  AOI211_X1 u1_u6_u1_U36 (.B( u1_u6_u1_n117 ) , .A( u1_u6_u1_n118 ) , .ZN( u1_u6_u1_n119 ) , .C2( u1_u6_u1_n146 ) , .C1( u1_u6_u1_n159 ) );
  NOR2_X1 u1_u6_u1_U37 (.A1( u1_u6_u1_n168 ) , .A2( u1_u6_u1_n176 ) , .ZN( u1_u6_u1_n98 ) );
  AOI211_X1 u1_u6_u1_U38 (.B( u1_u6_u1_n162 ) , .A( u1_u6_u1_n163 ) , .C2( u1_u6_u1_n164 ) , .ZN( u1_u6_u1_n165 ) , .C1( u1_u6_u1_n171 ) );
  AOI21_X1 u1_u6_u1_U39 (.A( u1_u6_u1_n160 ) , .B2( u1_u6_u1_n161 ) , .ZN( u1_u6_u1_n162 ) , .B1( u1_u6_u1_n182 ) );
  AOI221_X1 u1_u6_u1_U4 (.A( u1_u6_u1_n138 ) , .C2( u1_u6_u1_n139 ) , .C1( u1_u6_u1_n140 ) , .B2( u1_u6_u1_n141 ) , .ZN( u1_u6_u1_n142 ) , .B1( u1_u6_u1_n175 ) );
  OR2_X1 u1_u6_u1_U40 (.A2( u1_u6_u1_n157 ) , .A1( u1_u6_u1_n158 ) , .ZN( u1_u6_u1_n163 ) );
  NAND2_X1 u1_u6_u1_U41 (.A1( u1_u6_u1_n128 ) , .ZN( u1_u6_u1_n146 ) , .A2( u1_u6_u1_n160 ) );
  NAND2_X1 u1_u6_u1_U42 (.A2( u1_u6_u1_n112 ) , .ZN( u1_u6_u1_n139 ) , .A1( u1_u6_u1_n152 ) );
  NAND2_X1 u1_u6_u1_U43 (.A1( u1_u6_u1_n105 ) , .ZN( u1_u6_u1_n156 ) , .A2( u1_u6_u1_n99 ) );
  NOR2_X1 u1_u6_u1_U44 (.ZN( u1_u6_u1_n117 ) , .A1( u1_u6_u1_n121 ) , .A2( u1_u6_u1_n160 ) );
  OAI21_X1 u1_u6_u1_U45 (.B2( u1_u6_u1_n123 ) , .ZN( u1_u6_u1_n145 ) , .B1( u1_u6_u1_n160 ) , .A( u1_u6_u1_n185 ) );
  INV_X1 u1_u6_u1_U46 (.A( u1_u6_u1_n122 ) , .ZN( u1_u6_u1_n185 ) );
  AOI21_X1 u1_u6_u1_U47 (.B2( u1_u6_u1_n120 ) , .B1( u1_u6_u1_n121 ) , .ZN( u1_u6_u1_n122 ) , .A( u1_u6_u1_n128 ) );
  AOI21_X1 u1_u6_u1_U48 (.A( u1_u6_u1_n128 ) , .B2( u1_u6_u1_n129 ) , .ZN( u1_u6_u1_n130 ) , .B1( u1_u6_u1_n150 ) );
  NAND2_X1 u1_u6_u1_U49 (.ZN( u1_u6_u1_n112 ) , .A1( u1_u6_u1_n169 ) , .A2( u1_u6_u1_n170 ) );
  AOI211_X1 u1_u6_u1_U5 (.ZN( u1_u6_u1_n124 ) , .A( u1_u6_u1_n138 ) , .C2( u1_u6_u1_n139 ) , .B( u1_u6_u1_n145 ) , .C1( u1_u6_u1_n147 ) );
  NAND2_X1 u1_u6_u1_U50 (.ZN( u1_u6_u1_n129 ) , .A2( u1_u6_u1_n95 ) , .A1( u1_u6_u1_n98 ) );
  NAND2_X1 u1_u6_u1_U51 (.A1( u1_u6_u1_n102 ) , .ZN( u1_u6_u1_n154 ) , .A2( u1_u6_u1_n99 ) );
  NAND2_X1 u1_u6_u1_U52 (.A2( u1_u6_u1_n100 ) , .ZN( u1_u6_u1_n135 ) , .A1( u1_u6_u1_n99 ) );
  AOI21_X1 u1_u6_u1_U53 (.A( u1_u6_u1_n152 ) , .B2( u1_u6_u1_n153 ) , .B1( u1_u6_u1_n154 ) , .ZN( u1_u6_u1_n158 ) );
  INV_X1 u1_u6_u1_U54 (.A( u1_u6_u1_n160 ) , .ZN( u1_u6_u1_n175 ) );
  NAND2_X1 u1_u6_u1_U55 (.A1( u1_u6_u1_n100 ) , .ZN( u1_u6_u1_n116 ) , .A2( u1_u6_u1_n95 ) );
  NAND2_X1 u1_u6_u1_U56 (.A1( u1_u6_u1_n102 ) , .ZN( u1_u6_u1_n131 ) , .A2( u1_u6_u1_n95 ) );
  NAND2_X1 u1_u6_u1_U57 (.A2( u1_u6_u1_n104 ) , .ZN( u1_u6_u1_n121 ) , .A1( u1_u6_u1_n98 ) );
  NAND2_X1 u1_u6_u1_U58 (.A1( u1_u6_u1_n103 ) , .ZN( u1_u6_u1_n153 ) , .A2( u1_u6_u1_n98 ) );
  NAND2_X1 u1_u6_u1_U59 (.A2( u1_u6_u1_n104 ) , .A1( u1_u6_u1_n105 ) , .ZN( u1_u6_u1_n133 ) );
  AOI22_X1 u1_u6_u1_U6 (.B2( u1_u6_u1_n113 ) , .A2( u1_u6_u1_n114 ) , .ZN( u1_u6_u1_n125 ) , .A1( u1_u6_u1_n171 ) , .B1( u1_u6_u1_n173 ) );
  NAND2_X1 u1_u6_u1_U60 (.ZN( u1_u6_u1_n150 ) , .A2( u1_u6_u1_n98 ) , .A1( u1_u6_u1_n99 ) );
  NAND2_X1 u1_u6_u1_U61 (.A1( u1_u6_u1_n105 ) , .ZN( u1_u6_u1_n155 ) , .A2( u1_u6_u1_n95 ) );
  OAI21_X1 u1_u6_u1_U62 (.ZN( u1_u6_u1_n109 ) , .B1( u1_u6_u1_n129 ) , .B2( u1_u6_u1_n160 ) , .A( u1_u6_u1_n167 ) );
  NAND2_X1 u1_u6_u1_U63 (.A2( u1_u6_u1_n100 ) , .A1( u1_u6_u1_n103 ) , .ZN( u1_u6_u1_n120 ) );
  NAND2_X1 u1_u6_u1_U64 (.A1( u1_u6_u1_n102 ) , .A2( u1_u6_u1_n104 ) , .ZN( u1_u6_u1_n115 ) );
  NAND2_X1 u1_u6_u1_U65 (.A2( u1_u6_u1_n100 ) , .A1( u1_u6_u1_n104 ) , .ZN( u1_u6_u1_n151 ) );
  NAND2_X1 u1_u6_u1_U66 (.A2( u1_u6_u1_n103 ) , .A1( u1_u6_u1_n105 ) , .ZN( u1_u6_u1_n161 ) );
  INV_X1 u1_u6_u1_U67 (.A( u1_u6_u1_n152 ) , .ZN( u1_u6_u1_n173 ) );
  INV_X1 u1_u6_u1_U68 (.A( u1_u6_u1_n128 ) , .ZN( u1_u6_u1_n172 ) );
  NAND2_X1 u1_u6_u1_U69 (.A2( u1_u6_u1_n102 ) , .A1( u1_u6_u1_n103 ) , .ZN( u1_u6_u1_n123 ) );
  NAND2_X1 u1_u6_u1_U7 (.ZN( u1_u6_u1_n114 ) , .A1( u1_u6_u1_n134 ) , .A2( u1_u6_u1_n156 ) );
  NOR2_X1 u1_u6_u1_U70 (.A2( u1_u6_X_7 ) , .A1( u1_u6_X_8 ) , .ZN( u1_u6_u1_n95 ) );
  NOR2_X1 u1_u6_u1_U71 (.A1( u1_u6_X_12 ) , .A2( u1_u6_X_9 ) , .ZN( u1_u6_u1_n100 ) );
  NOR2_X1 u1_u6_u1_U72 (.A2( u1_u6_X_8 ) , .A1( u1_u6_u1_n177 ) , .ZN( u1_u6_u1_n99 ) );
  NOR2_X1 u1_u6_u1_U73 (.A2( u1_u6_X_12 ) , .ZN( u1_u6_u1_n102 ) , .A1( u1_u6_u1_n176 ) );
  NOR2_X1 u1_u6_u1_U74 (.A2( u1_u6_X_9 ) , .ZN( u1_u6_u1_n105 ) , .A1( u1_u6_u1_n168 ) );
  NAND2_X1 u1_u6_u1_U75 (.A1( u1_u6_X_10 ) , .ZN( u1_u6_u1_n160 ) , .A2( u1_u6_u1_n169 ) );
  NAND2_X1 u1_u6_u1_U76 (.A2( u1_u6_X_10 ) , .A1( u1_u6_X_11 ) , .ZN( u1_u6_u1_n152 ) );
  NAND2_X1 u1_u6_u1_U77 (.A1( u1_u6_X_11 ) , .ZN( u1_u6_u1_n128 ) , .A2( u1_u6_u1_n170 ) );
  AND2_X1 u1_u6_u1_U78 (.A2( u1_u6_X_7 ) , .A1( u1_u6_X_8 ) , .ZN( u1_u6_u1_n104 ) );
  AND2_X1 u1_u6_u1_U79 (.A1( u1_u6_X_8 ) , .ZN( u1_u6_u1_n103 ) , .A2( u1_u6_u1_n177 ) );
  AOI22_X1 u1_u6_u1_U8 (.B2( u1_u6_u1_n136 ) , .A2( u1_u6_u1_n137 ) , .ZN( u1_u6_u1_n143 ) , .A1( u1_u6_u1_n171 ) , .B1( u1_u6_u1_n173 ) );
  INV_X1 u1_u6_u1_U80 (.A( u1_u6_X_10 ) , .ZN( u1_u6_u1_n170 ) );
  INV_X1 u1_u6_u1_U81 (.A( u1_u6_X_9 ) , .ZN( u1_u6_u1_n176 ) );
  INV_X1 u1_u6_u1_U82 (.A( u1_u6_X_11 ) , .ZN( u1_u6_u1_n169 ) );
  INV_X1 u1_u6_u1_U83 (.A( u1_u6_X_12 ) , .ZN( u1_u6_u1_n168 ) );
  INV_X1 u1_u6_u1_U84 (.A( u1_u6_X_7 ) , .ZN( u1_u6_u1_n177 ) );
  NAND4_X1 u1_u6_u1_U85 (.ZN( u1_out6_18 ) , .A4( u1_u6_u1_n165 ) , .A3( u1_u6_u1_n166 ) , .A1( u1_u6_u1_n167 ) , .A2( u1_u6_u1_n186 ) );
  AOI22_X1 u1_u6_u1_U86 (.B2( u1_u6_u1_n146 ) , .B1( u1_u6_u1_n147 ) , .A2( u1_u6_u1_n148 ) , .ZN( u1_u6_u1_n166 ) , .A1( u1_u6_u1_n172 ) );
  INV_X1 u1_u6_u1_U87 (.A( u1_u6_u1_n145 ) , .ZN( u1_u6_u1_n186 ) );
  NAND4_X1 u1_u6_u1_U88 (.ZN( u1_out6_2 ) , .A4( u1_u6_u1_n142 ) , .A3( u1_u6_u1_n143 ) , .A2( u1_u6_u1_n144 ) , .A1( u1_u6_u1_n179 ) );
  OAI21_X1 u1_u6_u1_U89 (.B2( u1_u6_u1_n132 ) , .ZN( u1_u6_u1_n144 ) , .A( u1_u6_u1_n146 ) , .B1( u1_u6_u1_n180 ) );
  INV_X1 u1_u6_u1_U9 (.A( u1_u6_u1_n147 ) , .ZN( u1_u6_u1_n181 ) );
  INV_X1 u1_u6_u1_U90 (.A( u1_u6_u1_n130 ) , .ZN( u1_u6_u1_n179 ) );
  NAND4_X1 u1_u6_u1_U91 (.ZN( u1_out6_28 ) , .A4( u1_u6_u1_n124 ) , .A3( u1_u6_u1_n125 ) , .A2( u1_u6_u1_n126 ) , .A1( u1_u6_u1_n127 ) );
  OAI21_X1 u1_u6_u1_U92 (.ZN( u1_u6_u1_n127 ) , .B2( u1_u6_u1_n139 ) , .B1( u1_u6_u1_n175 ) , .A( u1_u6_u1_n183 ) );
  OAI21_X1 u1_u6_u1_U93 (.ZN( u1_u6_u1_n126 ) , .B2( u1_u6_u1_n140 ) , .A( u1_u6_u1_n146 ) , .B1( u1_u6_u1_n178 ) );
  OR4_X1 u1_u6_u1_U94 (.ZN( u1_out6_13 ) , .A4( u1_u6_u1_n108 ) , .A3( u1_u6_u1_n109 ) , .A2( u1_u6_u1_n110 ) , .A1( u1_u6_u1_n111 ) );
  AOI21_X1 u1_u6_u1_U95 (.ZN( u1_u6_u1_n111 ) , .A( u1_u6_u1_n128 ) , .B2( u1_u6_u1_n131 ) , .B1( u1_u6_u1_n135 ) );
  AOI21_X1 u1_u6_u1_U96 (.ZN( u1_u6_u1_n110 ) , .A( u1_u6_u1_n116 ) , .B1( u1_u6_u1_n152 ) , .B2( u1_u6_u1_n160 ) );
  NAND3_X1 u1_u6_u1_U97 (.A3( u1_u6_u1_n149 ) , .A2( u1_u6_u1_n150 ) , .A1( u1_u6_u1_n151 ) , .ZN( u1_u6_u1_n164 ) );
  NAND3_X1 u1_u6_u1_U98 (.A3( u1_u6_u1_n134 ) , .A2( u1_u6_u1_n135 ) , .ZN( u1_u6_u1_n136 ) , .A1( u1_u6_u1_n151 ) );
  NAND3_X1 u1_u6_u1_U99 (.A1( u1_u6_u1_n133 ) , .ZN( u1_u6_u1_n137 ) , .A2( u1_u6_u1_n154 ) , .A3( u1_u6_u1_n181 ) );
  AND3_X1 u1_u6_u7_U10 (.A3( u1_u6_u7_n110 ) , .A2( u1_u6_u7_n127 ) , .A1( u1_u6_u7_n132 ) , .ZN( u1_u6_u7_n92 ) );
  OAI21_X1 u1_u6_u7_U11 (.A( u1_u6_u7_n161 ) , .B1( u1_u6_u7_n168 ) , .B2( u1_u6_u7_n173 ) , .ZN( u1_u6_u7_n91 ) );
  AOI211_X1 u1_u6_u7_U12 (.A( u1_u6_u7_n117 ) , .ZN( u1_u6_u7_n118 ) , .C2( u1_u6_u7_n126 ) , .C1( u1_u6_u7_n177 ) , .B( u1_u6_u7_n180 ) );
  OAI22_X1 u1_u6_u7_U13 (.B1( u1_u6_u7_n115 ) , .ZN( u1_u6_u7_n117 ) , .A2( u1_u6_u7_n133 ) , .A1( u1_u6_u7_n137 ) , .B2( u1_u6_u7_n162 ) );
  INV_X1 u1_u6_u7_U14 (.A( u1_u6_u7_n116 ) , .ZN( u1_u6_u7_n180 ) );
  NOR3_X1 u1_u6_u7_U15 (.ZN( u1_u6_u7_n115 ) , .A3( u1_u6_u7_n145 ) , .A2( u1_u6_u7_n168 ) , .A1( u1_u6_u7_n169 ) );
  OAI211_X1 u1_u6_u7_U16 (.B( u1_u6_u7_n122 ) , .A( u1_u6_u7_n123 ) , .C2( u1_u6_u7_n124 ) , .ZN( u1_u6_u7_n154 ) , .C1( u1_u6_u7_n162 ) );
  AOI222_X1 u1_u6_u7_U17 (.ZN( u1_u6_u7_n122 ) , .C2( u1_u6_u7_n126 ) , .C1( u1_u6_u7_n145 ) , .B1( u1_u6_u7_n161 ) , .A2( u1_u6_u7_n165 ) , .B2( u1_u6_u7_n170 ) , .A1( u1_u6_u7_n176 ) );
  INV_X1 u1_u6_u7_U18 (.A( u1_u6_u7_n133 ) , .ZN( u1_u6_u7_n176 ) );
  NOR3_X1 u1_u6_u7_U19 (.A2( u1_u6_u7_n134 ) , .A1( u1_u6_u7_n135 ) , .ZN( u1_u6_u7_n136 ) , .A3( u1_u6_u7_n171 ) );
  NOR2_X1 u1_u6_u7_U20 (.A1( u1_u6_u7_n130 ) , .A2( u1_u6_u7_n134 ) , .ZN( u1_u6_u7_n153 ) );
  INV_X1 u1_u6_u7_U21 (.A( u1_u6_u7_n101 ) , .ZN( u1_u6_u7_n165 ) );
  NOR2_X1 u1_u6_u7_U22 (.ZN( u1_u6_u7_n111 ) , .A2( u1_u6_u7_n134 ) , .A1( u1_u6_u7_n169 ) );
  AOI21_X1 u1_u6_u7_U23 (.ZN( u1_u6_u7_n104 ) , .B2( u1_u6_u7_n112 ) , .B1( u1_u6_u7_n127 ) , .A( u1_u6_u7_n164 ) );
  AOI21_X1 u1_u6_u7_U24 (.ZN( u1_u6_u7_n106 ) , .B1( u1_u6_u7_n133 ) , .B2( u1_u6_u7_n146 ) , .A( u1_u6_u7_n162 ) );
  AOI21_X1 u1_u6_u7_U25 (.A( u1_u6_u7_n101 ) , .ZN( u1_u6_u7_n107 ) , .B2( u1_u6_u7_n128 ) , .B1( u1_u6_u7_n175 ) );
  INV_X1 u1_u6_u7_U26 (.A( u1_u6_u7_n138 ) , .ZN( u1_u6_u7_n171 ) );
  INV_X1 u1_u6_u7_U27 (.A( u1_u6_u7_n131 ) , .ZN( u1_u6_u7_n177 ) );
  INV_X1 u1_u6_u7_U28 (.A( u1_u6_u7_n110 ) , .ZN( u1_u6_u7_n174 ) );
  NAND2_X1 u1_u6_u7_U29 (.A1( u1_u6_u7_n129 ) , .A2( u1_u6_u7_n132 ) , .ZN( u1_u6_u7_n149 ) );
  OAI21_X1 u1_u6_u7_U3 (.ZN( u1_u6_u7_n159 ) , .A( u1_u6_u7_n165 ) , .B2( u1_u6_u7_n171 ) , .B1( u1_u6_u7_n174 ) );
  NAND2_X1 u1_u6_u7_U30 (.A1( u1_u6_u7_n113 ) , .A2( u1_u6_u7_n124 ) , .ZN( u1_u6_u7_n130 ) );
  INV_X1 u1_u6_u7_U31 (.A( u1_u6_u7_n112 ) , .ZN( u1_u6_u7_n173 ) );
  INV_X1 u1_u6_u7_U32 (.A( u1_u6_u7_n128 ) , .ZN( u1_u6_u7_n168 ) );
  INV_X1 u1_u6_u7_U33 (.A( u1_u6_u7_n148 ) , .ZN( u1_u6_u7_n169 ) );
  INV_X1 u1_u6_u7_U34 (.A( u1_u6_u7_n127 ) , .ZN( u1_u6_u7_n179 ) );
  NOR2_X1 u1_u6_u7_U35 (.ZN( u1_u6_u7_n101 ) , .A2( u1_u6_u7_n150 ) , .A1( u1_u6_u7_n156 ) );
  AOI211_X1 u1_u6_u7_U36 (.B( u1_u6_u7_n154 ) , .A( u1_u6_u7_n155 ) , .C1( u1_u6_u7_n156 ) , .ZN( u1_u6_u7_n157 ) , .C2( u1_u6_u7_n172 ) );
  INV_X1 u1_u6_u7_U37 (.A( u1_u6_u7_n153 ) , .ZN( u1_u6_u7_n172 ) );
  AOI211_X1 u1_u6_u7_U38 (.B( u1_u6_u7_n139 ) , .A( u1_u6_u7_n140 ) , .C2( u1_u6_u7_n141 ) , .ZN( u1_u6_u7_n142 ) , .C1( u1_u6_u7_n156 ) );
  NAND4_X1 u1_u6_u7_U39 (.A3( u1_u6_u7_n127 ) , .A2( u1_u6_u7_n128 ) , .A1( u1_u6_u7_n129 ) , .ZN( u1_u6_u7_n141 ) , .A4( u1_u6_u7_n147 ) );
  INV_X1 u1_u6_u7_U4 (.A( u1_u6_u7_n111 ) , .ZN( u1_u6_u7_n170 ) );
  AOI21_X1 u1_u6_u7_U40 (.A( u1_u6_u7_n137 ) , .B1( u1_u6_u7_n138 ) , .ZN( u1_u6_u7_n139 ) , .B2( u1_u6_u7_n146 ) );
  OAI22_X1 u1_u6_u7_U41 (.B1( u1_u6_u7_n136 ) , .ZN( u1_u6_u7_n140 ) , .A1( u1_u6_u7_n153 ) , .B2( u1_u6_u7_n162 ) , .A2( u1_u6_u7_n164 ) );
  AOI21_X1 u1_u6_u7_U42 (.ZN( u1_u6_u7_n123 ) , .B1( u1_u6_u7_n165 ) , .B2( u1_u6_u7_n177 ) , .A( u1_u6_u7_n97 ) );
  AOI21_X1 u1_u6_u7_U43 (.B2( u1_u6_u7_n113 ) , .B1( u1_u6_u7_n124 ) , .A( u1_u6_u7_n125 ) , .ZN( u1_u6_u7_n97 ) );
  INV_X1 u1_u6_u7_U44 (.A( u1_u6_u7_n125 ) , .ZN( u1_u6_u7_n161 ) );
  INV_X1 u1_u6_u7_U45 (.A( u1_u6_u7_n152 ) , .ZN( u1_u6_u7_n162 ) );
  AOI22_X1 u1_u6_u7_U46 (.A2( u1_u6_u7_n114 ) , .ZN( u1_u6_u7_n119 ) , .B1( u1_u6_u7_n130 ) , .A1( u1_u6_u7_n156 ) , .B2( u1_u6_u7_n165 ) );
  NAND2_X1 u1_u6_u7_U47 (.A2( u1_u6_u7_n112 ) , .ZN( u1_u6_u7_n114 ) , .A1( u1_u6_u7_n175 ) );
  AND2_X1 u1_u6_u7_U48 (.ZN( u1_u6_u7_n145 ) , .A2( u1_u6_u7_n98 ) , .A1( u1_u6_u7_n99 ) );
  NOR2_X1 u1_u6_u7_U49 (.ZN( u1_u6_u7_n137 ) , .A1( u1_u6_u7_n150 ) , .A2( u1_u6_u7_n161 ) );
  INV_X1 u1_u6_u7_U5 (.A( u1_u6_u7_n149 ) , .ZN( u1_u6_u7_n175 ) );
  AOI21_X1 u1_u6_u7_U50 (.ZN( u1_u6_u7_n105 ) , .B2( u1_u6_u7_n110 ) , .A( u1_u6_u7_n125 ) , .B1( u1_u6_u7_n147 ) );
  NAND2_X1 u1_u6_u7_U51 (.ZN( u1_u6_u7_n146 ) , .A1( u1_u6_u7_n95 ) , .A2( u1_u6_u7_n98 ) );
  NAND2_X1 u1_u6_u7_U52 (.A2( u1_u6_u7_n103 ) , .ZN( u1_u6_u7_n147 ) , .A1( u1_u6_u7_n93 ) );
  NAND2_X1 u1_u6_u7_U53 (.A1( u1_u6_u7_n103 ) , .ZN( u1_u6_u7_n127 ) , .A2( u1_u6_u7_n99 ) );
  OR2_X1 u1_u6_u7_U54 (.ZN( u1_u6_u7_n126 ) , .A2( u1_u6_u7_n152 ) , .A1( u1_u6_u7_n156 ) );
  NAND2_X1 u1_u6_u7_U55 (.A2( u1_u6_u7_n102 ) , .A1( u1_u6_u7_n103 ) , .ZN( u1_u6_u7_n133 ) );
  NAND2_X1 u1_u6_u7_U56 (.ZN( u1_u6_u7_n112 ) , .A2( u1_u6_u7_n96 ) , .A1( u1_u6_u7_n99 ) );
  NAND2_X1 u1_u6_u7_U57 (.A2( u1_u6_u7_n102 ) , .ZN( u1_u6_u7_n128 ) , .A1( u1_u6_u7_n98 ) );
  NAND2_X1 u1_u6_u7_U58 (.A1( u1_u6_u7_n100 ) , .ZN( u1_u6_u7_n113 ) , .A2( u1_u6_u7_n93 ) );
  NAND2_X1 u1_u6_u7_U59 (.A2( u1_u6_u7_n102 ) , .ZN( u1_u6_u7_n124 ) , .A1( u1_u6_u7_n96 ) );
  INV_X1 u1_u6_u7_U6 (.A( u1_u6_u7_n154 ) , .ZN( u1_u6_u7_n178 ) );
  NAND2_X1 u1_u6_u7_U60 (.ZN( u1_u6_u7_n110 ) , .A1( u1_u6_u7_n95 ) , .A2( u1_u6_u7_n96 ) );
  INV_X1 u1_u6_u7_U61 (.A( u1_u6_u7_n150 ) , .ZN( u1_u6_u7_n164 ) );
  AND2_X1 u1_u6_u7_U62 (.ZN( u1_u6_u7_n134 ) , .A1( u1_u6_u7_n93 ) , .A2( u1_u6_u7_n98 ) );
  NAND2_X1 u1_u6_u7_U63 (.A1( u1_u6_u7_n100 ) , .A2( u1_u6_u7_n102 ) , .ZN( u1_u6_u7_n129 ) );
  NAND2_X1 u1_u6_u7_U64 (.A2( u1_u6_u7_n103 ) , .ZN( u1_u6_u7_n131 ) , .A1( u1_u6_u7_n95 ) );
  NAND2_X1 u1_u6_u7_U65 (.A1( u1_u6_u7_n100 ) , .ZN( u1_u6_u7_n138 ) , .A2( u1_u6_u7_n99 ) );
  NAND2_X1 u1_u6_u7_U66 (.ZN( u1_u6_u7_n132 ) , .A1( u1_u6_u7_n93 ) , .A2( u1_u6_u7_n96 ) );
  NAND2_X1 u1_u6_u7_U67 (.A1( u1_u6_u7_n100 ) , .ZN( u1_u6_u7_n148 ) , .A2( u1_u6_u7_n95 ) );
  NOR2_X1 u1_u6_u7_U68 (.A2( u1_u6_X_47 ) , .ZN( u1_u6_u7_n150 ) , .A1( u1_u6_u7_n163 ) );
  NOR2_X1 u1_u6_u7_U69 (.A2( u1_u6_X_43 ) , .A1( u1_u6_X_44 ) , .ZN( u1_u6_u7_n103 ) );
  AOI211_X1 u1_u6_u7_U7 (.ZN( u1_u6_u7_n116 ) , .A( u1_u6_u7_n155 ) , .C1( u1_u6_u7_n161 ) , .C2( u1_u6_u7_n171 ) , .B( u1_u6_u7_n94 ) );
  NOR2_X1 u1_u6_u7_U70 (.A2( u1_u6_X_48 ) , .A1( u1_u6_u7_n166 ) , .ZN( u1_u6_u7_n95 ) );
  NOR2_X1 u1_u6_u7_U71 (.A2( u1_u6_X_45 ) , .A1( u1_u6_X_48 ) , .ZN( u1_u6_u7_n99 ) );
  NOR2_X1 u1_u6_u7_U72 (.A2( u1_u6_X_44 ) , .A1( u1_u6_u7_n167 ) , .ZN( u1_u6_u7_n98 ) );
  NOR2_X1 u1_u6_u7_U73 (.A2( u1_u6_X_46 ) , .A1( u1_u6_X_47 ) , .ZN( u1_u6_u7_n152 ) );
  AND2_X1 u1_u6_u7_U74 (.A1( u1_u6_X_47 ) , .ZN( u1_u6_u7_n156 ) , .A2( u1_u6_u7_n163 ) );
  NAND2_X1 u1_u6_u7_U75 (.A2( u1_u6_X_46 ) , .A1( u1_u6_X_47 ) , .ZN( u1_u6_u7_n125 ) );
  AND2_X1 u1_u6_u7_U76 (.A2( u1_u6_X_45 ) , .A1( u1_u6_X_48 ) , .ZN( u1_u6_u7_n102 ) );
  AND2_X1 u1_u6_u7_U77 (.A2( u1_u6_X_43 ) , .A1( u1_u6_X_44 ) , .ZN( u1_u6_u7_n96 ) );
  AND2_X1 u1_u6_u7_U78 (.A1( u1_u6_X_44 ) , .ZN( u1_u6_u7_n100 ) , .A2( u1_u6_u7_n167 ) );
  AND2_X1 u1_u6_u7_U79 (.A1( u1_u6_X_48 ) , .A2( u1_u6_u7_n166 ) , .ZN( u1_u6_u7_n93 ) );
  OAI222_X1 u1_u6_u7_U8 (.C2( u1_u6_u7_n101 ) , .B2( u1_u6_u7_n111 ) , .A1( u1_u6_u7_n113 ) , .C1( u1_u6_u7_n146 ) , .A2( u1_u6_u7_n162 ) , .B1( u1_u6_u7_n164 ) , .ZN( u1_u6_u7_n94 ) );
  INV_X1 u1_u6_u7_U80 (.A( u1_u6_X_46 ) , .ZN( u1_u6_u7_n163 ) );
  INV_X1 u1_u6_u7_U81 (.A( u1_u6_X_43 ) , .ZN( u1_u6_u7_n167 ) );
  INV_X1 u1_u6_u7_U82 (.A( u1_u6_X_45 ) , .ZN( u1_u6_u7_n166 ) );
  NAND4_X1 u1_u6_u7_U83 (.ZN( u1_out6_5 ) , .A4( u1_u6_u7_n108 ) , .A3( u1_u6_u7_n109 ) , .A1( u1_u6_u7_n116 ) , .A2( u1_u6_u7_n123 ) );
  AOI22_X1 u1_u6_u7_U84 (.ZN( u1_u6_u7_n109 ) , .A2( u1_u6_u7_n126 ) , .B2( u1_u6_u7_n145 ) , .B1( u1_u6_u7_n156 ) , .A1( u1_u6_u7_n171 ) );
  NOR4_X1 u1_u6_u7_U85 (.A4( u1_u6_u7_n104 ) , .A3( u1_u6_u7_n105 ) , .A2( u1_u6_u7_n106 ) , .A1( u1_u6_u7_n107 ) , .ZN( u1_u6_u7_n108 ) );
  NAND4_X1 u1_u6_u7_U86 (.ZN( u1_out6_21 ) , .A4( u1_u6_u7_n157 ) , .A3( u1_u6_u7_n158 ) , .A2( u1_u6_u7_n159 ) , .A1( u1_u6_u7_n160 ) );
  OAI21_X1 u1_u6_u7_U87 (.B1( u1_u6_u7_n145 ) , .ZN( u1_u6_u7_n160 ) , .A( u1_u6_u7_n161 ) , .B2( u1_u6_u7_n177 ) );
  AOI22_X1 u1_u6_u7_U88 (.B2( u1_u6_u7_n149 ) , .B1( u1_u6_u7_n150 ) , .A2( u1_u6_u7_n151 ) , .A1( u1_u6_u7_n152 ) , .ZN( u1_u6_u7_n158 ) );
  NAND4_X1 u1_u6_u7_U89 (.ZN( u1_out6_15 ) , .A4( u1_u6_u7_n142 ) , .A3( u1_u6_u7_n143 ) , .A2( u1_u6_u7_n144 ) , .A1( u1_u6_u7_n178 ) );
  OAI221_X1 u1_u6_u7_U9 (.C1( u1_u6_u7_n101 ) , .C2( u1_u6_u7_n147 ) , .ZN( u1_u6_u7_n155 ) , .B2( u1_u6_u7_n162 ) , .A( u1_u6_u7_n91 ) , .B1( u1_u6_u7_n92 ) );
  OR2_X1 u1_u6_u7_U90 (.A2( u1_u6_u7_n125 ) , .A1( u1_u6_u7_n129 ) , .ZN( u1_u6_u7_n144 ) );
  AOI22_X1 u1_u6_u7_U91 (.A2( u1_u6_u7_n126 ) , .ZN( u1_u6_u7_n143 ) , .B2( u1_u6_u7_n165 ) , .B1( u1_u6_u7_n173 ) , .A1( u1_u6_u7_n174 ) );
  NAND4_X1 u1_u6_u7_U92 (.ZN( u1_out6_27 ) , .A4( u1_u6_u7_n118 ) , .A3( u1_u6_u7_n119 ) , .A2( u1_u6_u7_n120 ) , .A1( u1_u6_u7_n121 ) );
  OAI21_X1 u1_u6_u7_U93 (.ZN( u1_u6_u7_n121 ) , .B2( u1_u6_u7_n145 ) , .A( u1_u6_u7_n150 ) , .B1( u1_u6_u7_n174 ) );
  OAI21_X1 u1_u6_u7_U94 (.ZN( u1_u6_u7_n120 ) , .A( u1_u6_u7_n161 ) , .B2( u1_u6_u7_n170 ) , .B1( u1_u6_u7_n179 ) );
  NAND3_X1 u1_u6_u7_U95 (.A3( u1_u6_u7_n146 ) , .A2( u1_u6_u7_n147 ) , .A1( u1_u6_u7_n148 ) , .ZN( u1_u6_u7_n151 ) );
  NAND3_X1 u1_u6_u7_U96 (.A3( u1_u6_u7_n131 ) , .A2( u1_u6_u7_n132 ) , .A1( u1_u6_u7_n133 ) , .ZN( u1_u6_u7_n135 ) );
  XOR2_X1 u1_u7_U10 (.B( u1_K8_45 ) , .A( u1_R6_30 ) , .Z( u1_u7_X_45 ) );
  XOR2_X1 u1_u7_U9 (.B( u1_K8_46 ) , .A( u1_R6_31 ) , .Z( u1_u7_X_46 ) );
  OAI221_X1 u1_u7_u7_U10 (.C1( u1_u7_u7_n101 ) , .C2( u1_u7_u7_n147 ) , .ZN( u1_u7_u7_n155 ) , .B2( u1_u7_u7_n162 ) , .A( u1_u7_u7_n91 ) , .B1( u1_u7_u7_n92 ) );
  AND3_X1 u1_u7_u7_U11 (.A3( u1_u7_u7_n110 ) , .A2( u1_u7_u7_n127 ) , .A1( u1_u7_u7_n132 ) , .ZN( u1_u7_u7_n92 ) );
  OAI21_X1 u1_u7_u7_U12 (.A( u1_u7_u7_n161 ) , .B1( u1_u7_u7_n168 ) , .B2( u1_u7_u7_n173 ) , .ZN( u1_u7_u7_n91 ) );
  AOI211_X1 u1_u7_u7_U13 (.A( u1_u7_u7_n117 ) , .ZN( u1_u7_u7_n118 ) , .C2( u1_u7_u7_n126 ) , .C1( u1_u7_u7_n177 ) , .B( u1_u7_u7_n180 ) );
  OAI22_X1 u1_u7_u7_U14 (.B1( u1_u7_u7_n115 ) , .ZN( u1_u7_u7_n117 ) , .A2( u1_u7_u7_n133 ) , .A1( u1_u7_u7_n137 ) , .B2( u1_u7_u7_n162 ) );
  INV_X1 u1_u7_u7_U15 (.A( u1_u7_u7_n116 ) , .ZN( u1_u7_u7_n180 ) );
  NOR3_X1 u1_u7_u7_U16 (.ZN( u1_u7_u7_n115 ) , .A3( u1_u7_u7_n145 ) , .A2( u1_u7_u7_n168 ) , .A1( u1_u7_u7_n169 ) );
  NOR3_X1 u1_u7_u7_U17 (.A2( u1_u7_u7_n134 ) , .A1( u1_u7_u7_n135 ) , .ZN( u1_u7_u7_n136 ) , .A3( u1_u7_u7_n171 ) );
  NOR2_X1 u1_u7_u7_U18 (.A1( u1_u7_u7_n130 ) , .A2( u1_u7_u7_n134 ) , .ZN( u1_u7_u7_n153 ) );
  NOR2_X1 u1_u7_u7_U19 (.ZN( u1_u7_u7_n111 ) , .A2( u1_u7_u7_n134 ) , .A1( u1_u7_u7_n169 ) );
  AOI21_X1 u1_u7_u7_U20 (.ZN( u1_u7_u7_n104 ) , .B2( u1_u7_u7_n112 ) , .B1( u1_u7_u7_n127 ) , .A( u1_u7_u7_n164 ) );
  AOI21_X1 u1_u7_u7_U21 (.ZN( u1_u7_u7_n106 ) , .B1( u1_u7_u7_n133 ) , .B2( u1_u7_u7_n146 ) , .A( u1_u7_u7_n162 ) );
  AOI21_X1 u1_u7_u7_U22 (.A( u1_u7_u7_n101 ) , .ZN( u1_u7_u7_n107 ) , .B2( u1_u7_u7_n128 ) , .B1( u1_u7_u7_n175 ) );
  INV_X1 u1_u7_u7_U23 (.A( u1_u7_u7_n101 ) , .ZN( u1_u7_u7_n165 ) );
  INV_X1 u1_u7_u7_U24 (.A( u1_u7_u7_n138 ) , .ZN( u1_u7_u7_n171 ) );
  INV_X1 u1_u7_u7_U25 (.A( u1_u7_u7_n131 ) , .ZN( u1_u7_u7_n177 ) );
  INV_X1 u1_u7_u7_U26 (.A( u1_u7_u7_n110 ) , .ZN( u1_u7_u7_n174 ) );
  NAND2_X1 u1_u7_u7_U27 (.A1( u1_u7_u7_n129 ) , .A2( u1_u7_u7_n132 ) , .ZN( u1_u7_u7_n149 ) );
  NAND2_X1 u1_u7_u7_U28 (.A1( u1_u7_u7_n113 ) , .A2( u1_u7_u7_n124 ) , .ZN( u1_u7_u7_n130 ) );
  INV_X1 u1_u7_u7_U29 (.A( u1_u7_u7_n128 ) , .ZN( u1_u7_u7_n168 ) );
  OAI21_X1 u1_u7_u7_U3 (.ZN( u1_u7_u7_n159 ) , .A( u1_u7_u7_n165 ) , .B2( u1_u7_u7_n171 ) , .B1( u1_u7_u7_n174 ) );
  INV_X1 u1_u7_u7_U30 (.A( u1_u7_u7_n148 ) , .ZN( u1_u7_u7_n169 ) );
  INV_X1 u1_u7_u7_U31 (.A( u1_u7_u7_n112 ) , .ZN( u1_u7_u7_n173 ) );
  INV_X1 u1_u7_u7_U32 (.A( u1_u7_u7_n127 ) , .ZN( u1_u7_u7_n179 ) );
  NOR2_X1 u1_u7_u7_U33 (.ZN( u1_u7_u7_n101 ) , .A2( u1_u7_u7_n150 ) , .A1( u1_u7_u7_n156 ) );
  AOI211_X1 u1_u7_u7_U34 (.B( u1_u7_u7_n154 ) , .A( u1_u7_u7_n155 ) , .C1( u1_u7_u7_n156 ) , .ZN( u1_u7_u7_n157 ) , .C2( u1_u7_u7_n172 ) );
  INV_X1 u1_u7_u7_U35 (.A( u1_u7_u7_n153 ) , .ZN( u1_u7_u7_n172 ) );
  AOI211_X1 u1_u7_u7_U36 (.B( u1_u7_u7_n139 ) , .A( u1_u7_u7_n140 ) , .C2( u1_u7_u7_n141 ) , .ZN( u1_u7_u7_n142 ) , .C1( u1_u7_u7_n156 ) );
  NAND4_X1 u1_u7_u7_U37 (.A3( u1_u7_u7_n127 ) , .A2( u1_u7_u7_n128 ) , .A1( u1_u7_u7_n129 ) , .ZN( u1_u7_u7_n141 ) , .A4( u1_u7_u7_n147 ) );
  AOI21_X1 u1_u7_u7_U38 (.A( u1_u7_u7_n137 ) , .B1( u1_u7_u7_n138 ) , .ZN( u1_u7_u7_n139 ) , .B2( u1_u7_u7_n146 ) );
  OAI22_X1 u1_u7_u7_U39 (.B1( u1_u7_u7_n136 ) , .ZN( u1_u7_u7_n140 ) , .A1( u1_u7_u7_n153 ) , .B2( u1_u7_u7_n162 ) , .A2( u1_u7_u7_n164 ) );
  INV_X1 u1_u7_u7_U4 (.A( u1_u7_u7_n149 ) , .ZN( u1_u7_u7_n175 ) );
  INV_X1 u1_u7_u7_U40 (.A( u1_u7_u7_n125 ) , .ZN( u1_u7_u7_n161 ) );
  AOI21_X1 u1_u7_u7_U41 (.ZN( u1_u7_u7_n123 ) , .B1( u1_u7_u7_n165 ) , .B2( u1_u7_u7_n177 ) , .A( u1_u7_u7_n97 ) );
  AOI21_X1 u1_u7_u7_U42 (.B2( u1_u7_u7_n113 ) , .B1( u1_u7_u7_n124 ) , .A( u1_u7_u7_n125 ) , .ZN( u1_u7_u7_n97 ) );
  INV_X1 u1_u7_u7_U43 (.A( u1_u7_u7_n152 ) , .ZN( u1_u7_u7_n162 ) );
  AOI22_X1 u1_u7_u7_U44 (.A2( u1_u7_u7_n114 ) , .ZN( u1_u7_u7_n119 ) , .B1( u1_u7_u7_n130 ) , .A1( u1_u7_u7_n156 ) , .B2( u1_u7_u7_n165 ) );
  NAND2_X1 u1_u7_u7_U45 (.A2( u1_u7_u7_n112 ) , .ZN( u1_u7_u7_n114 ) , .A1( u1_u7_u7_n175 ) );
  NOR2_X1 u1_u7_u7_U46 (.ZN( u1_u7_u7_n137 ) , .A1( u1_u7_u7_n150 ) , .A2( u1_u7_u7_n161 ) );
  AND2_X1 u1_u7_u7_U47 (.ZN( u1_u7_u7_n145 ) , .A2( u1_u7_u7_n98 ) , .A1( u1_u7_u7_n99 ) );
  AOI21_X1 u1_u7_u7_U48 (.ZN( u1_u7_u7_n105 ) , .B2( u1_u7_u7_n110 ) , .A( u1_u7_u7_n125 ) , .B1( u1_u7_u7_n147 ) );
  NAND2_X1 u1_u7_u7_U49 (.ZN( u1_u7_u7_n146 ) , .A1( u1_u7_u7_n95 ) , .A2( u1_u7_u7_n98 ) );
  INV_X1 u1_u7_u7_U5 (.A( u1_u7_u7_n154 ) , .ZN( u1_u7_u7_n178 ) );
  NAND2_X1 u1_u7_u7_U50 (.A2( u1_u7_u7_n103 ) , .ZN( u1_u7_u7_n147 ) , .A1( u1_u7_u7_n93 ) );
  NAND2_X1 u1_u7_u7_U51 (.A1( u1_u7_u7_n103 ) , .ZN( u1_u7_u7_n127 ) , .A2( u1_u7_u7_n99 ) );
  NAND2_X1 u1_u7_u7_U52 (.A2( u1_u7_u7_n102 ) , .A1( u1_u7_u7_n103 ) , .ZN( u1_u7_u7_n133 ) );
  OR2_X1 u1_u7_u7_U53 (.ZN( u1_u7_u7_n126 ) , .A2( u1_u7_u7_n152 ) , .A1( u1_u7_u7_n156 ) );
  NAND2_X1 u1_u7_u7_U54 (.ZN( u1_u7_u7_n112 ) , .A2( u1_u7_u7_n96 ) , .A1( u1_u7_u7_n99 ) );
  NAND2_X1 u1_u7_u7_U55 (.A2( u1_u7_u7_n102 ) , .ZN( u1_u7_u7_n128 ) , .A1( u1_u7_u7_n98 ) );
  INV_X1 u1_u7_u7_U56 (.A( u1_u7_u7_n150 ) , .ZN( u1_u7_u7_n164 ) );
  AND2_X1 u1_u7_u7_U57 (.ZN( u1_u7_u7_n134 ) , .A1( u1_u7_u7_n93 ) , .A2( u1_u7_u7_n98 ) );
  NAND2_X1 u1_u7_u7_U58 (.ZN( u1_u7_u7_n110 ) , .A1( u1_u7_u7_n95 ) , .A2( u1_u7_u7_n96 ) );
  NAND2_X1 u1_u7_u7_U59 (.A2( u1_u7_u7_n102 ) , .ZN( u1_u7_u7_n124 ) , .A1( u1_u7_u7_n96 ) );
  INV_X1 u1_u7_u7_U6 (.A( u1_u7_u7_n111 ) , .ZN( u1_u7_u7_n170 ) );
  NAND2_X1 u1_u7_u7_U60 (.ZN( u1_u7_u7_n132 ) , .A1( u1_u7_u7_n93 ) , .A2( u1_u7_u7_n96 ) );
  NAND2_X1 u1_u7_u7_U61 (.A2( u1_u7_u7_n103 ) , .ZN( u1_u7_u7_n131 ) , .A1( u1_u7_u7_n95 ) );
  NOR2_X1 u1_u7_u7_U62 (.A2( u1_u7_X_47 ) , .ZN( u1_u7_u7_n150 ) , .A1( u1_u7_u7_n163 ) );
  NOR2_X1 u1_u7_u7_U63 (.A2( u1_u7_X_43 ) , .A1( u1_u7_X_44 ) , .ZN( u1_u7_u7_n103 ) );
  NOR2_X1 u1_u7_u7_U64 (.A2( u1_u7_X_48 ) , .A1( u1_u7_u7_n166 ) , .ZN( u1_u7_u7_n95 ) );
  NOR2_X1 u1_u7_u7_U65 (.A2( u1_u7_X_44 ) , .A1( u1_u7_u7_n167 ) , .ZN( u1_u7_u7_n98 ) );
  NOR2_X1 u1_u7_u7_U66 (.A2( u1_u7_X_45 ) , .A1( u1_u7_X_48 ) , .ZN( u1_u7_u7_n99 ) );
  NOR2_X1 u1_u7_u7_U67 (.A2( u1_u7_X_46 ) , .A1( u1_u7_X_47 ) , .ZN( u1_u7_u7_n152 ) );
  AND2_X1 u1_u7_u7_U68 (.A1( u1_u7_X_47 ) , .ZN( u1_u7_u7_n156 ) , .A2( u1_u7_u7_n163 ) );
  NAND2_X1 u1_u7_u7_U69 (.A2( u1_u7_X_46 ) , .A1( u1_u7_X_47 ) , .ZN( u1_u7_u7_n125 ) );
  AOI211_X1 u1_u7_u7_U7 (.ZN( u1_u7_u7_n116 ) , .A( u1_u7_u7_n155 ) , .C1( u1_u7_u7_n161 ) , .C2( u1_u7_u7_n171 ) , .B( u1_u7_u7_n94 ) );
  AND2_X1 u1_u7_u7_U70 (.A2( u1_u7_X_43 ) , .A1( u1_u7_X_44 ) , .ZN( u1_u7_u7_n96 ) );
  AND2_X1 u1_u7_u7_U71 (.A2( u1_u7_X_45 ) , .A1( u1_u7_X_48 ) , .ZN( u1_u7_u7_n102 ) );
  AND2_X1 u1_u7_u7_U72 (.A1( u1_u7_X_48 ) , .A2( u1_u7_u7_n166 ) , .ZN( u1_u7_u7_n93 ) );
  INV_X1 u1_u7_u7_U73 (.A( u1_u7_X_46 ) , .ZN( u1_u7_u7_n163 ) );
  AND2_X1 u1_u7_u7_U74 (.A1( u1_u7_X_44 ) , .ZN( u1_u7_u7_n100 ) , .A2( u1_u7_u7_n167 ) );
  INV_X1 u1_u7_u7_U75 (.A( u1_u7_X_45 ) , .ZN( u1_u7_u7_n166 ) );
  INV_X1 u1_u7_u7_U76 (.A( u1_u7_X_43 ) , .ZN( u1_u7_u7_n167 ) );
  NAND4_X1 u1_u7_u7_U77 (.ZN( u1_out7_5 ) , .A4( u1_u7_u7_n108 ) , .A3( u1_u7_u7_n109 ) , .A1( u1_u7_u7_n116 ) , .A2( u1_u7_u7_n123 ) );
  AOI22_X1 u1_u7_u7_U78 (.ZN( u1_u7_u7_n109 ) , .A2( u1_u7_u7_n126 ) , .B2( u1_u7_u7_n145 ) , .B1( u1_u7_u7_n156 ) , .A1( u1_u7_u7_n171 ) );
  NOR4_X1 u1_u7_u7_U79 (.A4( u1_u7_u7_n104 ) , .A3( u1_u7_u7_n105 ) , .A2( u1_u7_u7_n106 ) , .A1( u1_u7_u7_n107 ) , .ZN( u1_u7_u7_n108 ) );
  OAI222_X1 u1_u7_u7_U8 (.C2( u1_u7_u7_n101 ) , .B2( u1_u7_u7_n111 ) , .A1( u1_u7_u7_n113 ) , .C1( u1_u7_u7_n146 ) , .A2( u1_u7_u7_n162 ) , .B1( u1_u7_u7_n164 ) , .ZN( u1_u7_u7_n94 ) );
  NAND4_X1 u1_u7_u7_U80 (.ZN( u1_out7_27 ) , .A4( u1_u7_u7_n118 ) , .A3( u1_u7_u7_n119 ) , .A2( u1_u7_u7_n120 ) , .A1( u1_u7_u7_n121 ) );
  OAI21_X1 u1_u7_u7_U81 (.ZN( u1_u7_u7_n121 ) , .B2( u1_u7_u7_n145 ) , .A( u1_u7_u7_n150 ) , .B1( u1_u7_u7_n174 ) );
  OAI21_X1 u1_u7_u7_U82 (.ZN( u1_u7_u7_n120 ) , .A( u1_u7_u7_n161 ) , .B2( u1_u7_u7_n170 ) , .B1( u1_u7_u7_n179 ) );
  NAND4_X1 u1_u7_u7_U83 (.ZN( u1_out7_21 ) , .A4( u1_u7_u7_n157 ) , .A3( u1_u7_u7_n158 ) , .A2( u1_u7_u7_n159 ) , .A1( u1_u7_u7_n160 ) );
  OAI21_X1 u1_u7_u7_U84 (.B1( u1_u7_u7_n145 ) , .ZN( u1_u7_u7_n160 ) , .A( u1_u7_u7_n161 ) , .B2( u1_u7_u7_n177 ) );
  AOI22_X1 u1_u7_u7_U85 (.B2( u1_u7_u7_n149 ) , .B1( u1_u7_u7_n150 ) , .A2( u1_u7_u7_n151 ) , .A1( u1_u7_u7_n152 ) , .ZN( u1_u7_u7_n158 ) );
  NAND4_X1 u1_u7_u7_U86 (.ZN( u1_out7_15 ) , .A4( u1_u7_u7_n142 ) , .A3( u1_u7_u7_n143 ) , .A2( u1_u7_u7_n144 ) , .A1( u1_u7_u7_n178 ) );
  OR2_X1 u1_u7_u7_U87 (.A2( u1_u7_u7_n125 ) , .A1( u1_u7_u7_n129 ) , .ZN( u1_u7_u7_n144 ) );
  AOI22_X1 u1_u7_u7_U88 (.A2( u1_u7_u7_n126 ) , .ZN( u1_u7_u7_n143 ) , .B2( u1_u7_u7_n165 ) , .B1( u1_u7_u7_n173 ) , .A1( u1_u7_u7_n174 ) );
  NAND2_X1 u1_u7_u7_U89 (.A1( u1_u7_u7_n100 ) , .ZN( u1_u7_u7_n148 ) , .A2( u1_u7_u7_n95 ) );
  INV_X1 u1_u7_u7_U9 (.A( u1_u7_u7_n133 ) , .ZN( u1_u7_u7_n176 ) );
  NAND2_X1 u1_u7_u7_U90 (.A1( u1_u7_u7_n100 ) , .ZN( u1_u7_u7_n113 ) , .A2( u1_u7_u7_n93 ) );
  NAND2_X1 u1_u7_u7_U91 (.A1( u1_u7_u7_n100 ) , .ZN( u1_u7_u7_n138 ) , .A2( u1_u7_u7_n99 ) );
  NAND2_X1 u1_u7_u7_U92 (.A1( u1_u7_u7_n100 ) , .A2( u1_u7_u7_n102 ) , .ZN( u1_u7_u7_n129 ) );
  OAI211_X1 u1_u7_u7_U93 (.B( u1_u7_u7_n122 ) , .A( u1_u7_u7_n123 ) , .C2( u1_u7_u7_n124 ) , .ZN( u1_u7_u7_n154 ) , .C1( u1_u7_u7_n162 ) );
  AOI222_X1 u1_u7_u7_U94 (.ZN( u1_u7_u7_n122 ) , .C2( u1_u7_u7_n126 ) , .C1( u1_u7_u7_n145 ) , .B1( u1_u7_u7_n161 ) , .A2( u1_u7_u7_n165 ) , .B2( u1_u7_u7_n170 ) , .A1( u1_u7_u7_n176 ) );
  NAND3_X1 u1_u7_u7_U95 (.A3( u1_u7_u7_n146 ) , .A2( u1_u7_u7_n147 ) , .A1( u1_u7_u7_n148 ) , .ZN( u1_u7_u7_n151 ) );
  NAND3_X1 u1_u7_u7_U96 (.A3( u1_u7_u7_n131 ) , .A2( u1_u7_u7_n132 ) , .A1( u1_u7_u7_n133 ) , .ZN( u1_u7_u7_n135 ) );
  XOR2_X1 u1_u8_U16 (.B( u1_K9_3 ) , .A( u1_R7_2 ) , .Z( u1_u8_X_3 ) );
  XOR2_X1 u1_u8_U6 (.B( u1_K9_4 ) , .A( u1_R7_3 ) , .Z( u1_u8_X_4 ) );
  AND2_X1 u1_u8_u0_U10 (.A1( u1_u8_u0_n131 ) , .ZN( u1_u8_u0_n141 ) , .A2( u1_u8_u0_n150 ) );
  AND3_X1 u1_u8_u0_U11 (.A2( u1_u8_u0_n112 ) , .ZN( u1_u8_u0_n127 ) , .A3( u1_u8_u0_n130 ) , .A1( u1_u8_u0_n148 ) );
  AND2_X1 u1_u8_u0_U12 (.ZN( u1_u8_u0_n107 ) , .A1( u1_u8_u0_n130 ) , .A2( u1_u8_u0_n140 ) );
  AND2_X1 u1_u8_u0_U13 (.A2( u1_u8_u0_n129 ) , .A1( u1_u8_u0_n130 ) , .ZN( u1_u8_u0_n151 ) );
  AND2_X1 u1_u8_u0_U14 (.A1( u1_u8_u0_n108 ) , .A2( u1_u8_u0_n125 ) , .ZN( u1_u8_u0_n145 ) );
  INV_X1 u1_u8_u0_U15 (.A( u1_u8_u0_n143 ) , .ZN( u1_u8_u0_n173 ) );
  NOR2_X1 u1_u8_u0_U16 (.A2( u1_u8_u0_n136 ) , .ZN( u1_u8_u0_n147 ) , .A1( u1_u8_u0_n160 ) );
  AOI21_X1 u1_u8_u0_U17 (.B1( u1_u8_u0_n103 ) , .ZN( u1_u8_u0_n132 ) , .A( u1_u8_u0_n165 ) , .B2( u1_u8_u0_n93 ) );
  OAI22_X1 u1_u8_u0_U18 (.B1( u1_u8_u0_n131 ) , .A1( u1_u8_u0_n144 ) , .B2( u1_u8_u0_n147 ) , .A2( u1_u8_u0_n90 ) , .ZN( u1_u8_u0_n91 ) );
  AND3_X1 u1_u8_u0_U19 (.A3( u1_u8_u0_n121 ) , .A2( u1_u8_u0_n125 ) , .A1( u1_u8_u0_n148 ) , .ZN( u1_u8_u0_n90 ) );
  OAI22_X1 u1_u8_u0_U20 (.B1( u1_u8_u0_n125 ) , .ZN( u1_u8_u0_n126 ) , .A1( u1_u8_u0_n138 ) , .A2( u1_u8_u0_n146 ) , .B2( u1_u8_u0_n147 ) );
  NOR2_X1 u1_u8_u0_U21 (.A1( u1_u8_u0_n163 ) , .A2( u1_u8_u0_n164 ) , .ZN( u1_u8_u0_n95 ) );
  AOI22_X1 u1_u8_u0_U22 (.B2( u1_u8_u0_n109 ) , .A2( u1_u8_u0_n110 ) , .ZN( u1_u8_u0_n111 ) , .B1( u1_u8_u0_n118 ) , .A1( u1_u8_u0_n160 ) );
  NAND2_X1 u1_u8_u0_U23 (.A2( u1_u8_u0_n102 ) , .A1( u1_u8_u0_n103 ) , .ZN( u1_u8_u0_n149 ) );
  INV_X1 u1_u8_u0_U24 (.A( u1_u8_u0_n136 ) , .ZN( u1_u8_u0_n161 ) );
  INV_X1 u1_u8_u0_U25 (.A( u1_u8_u0_n118 ) , .ZN( u1_u8_u0_n158 ) );
  NAND2_X1 u1_u8_u0_U26 (.A2( u1_u8_u0_n100 ) , .ZN( u1_u8_u0_n131 ) , .A1( u1_u8_u0_n92 ) );
  NAND2_X1 u1_u8_u0_U27 (.ZN( u1_u8_u0_n108 ) , .A1( u1_u8_u0_n92 ) , .A2( u1_u8_u0_n94 ) );
  AOI21_X1 u1_u8_u0_U28 (.ZN( u1_u8_u0_n104 ) , .B1( u1_u8_u0_n107 ) , .B2( u1_u8_u0_n141 ) , .A( u1_u8_u0_n144 ) );
  AOI21_X1 u1_u8_u0_U29 (.B1( u1_u8_u0_n127 ) , .B2( u1_u8_u0_n129 ) , .A( u1_u8_u0_n138 ) , .ZN( u1_u8_u0_n96 ) );
  INV_X1 u1_u8_u0_U3 (.A( u1_u8_u0_n113 ) , .ZN( u1_u8_u0_n166 ) );
  NAND2_X1 u1_u8_u0_U30 (.A2( u1_u8_u0_n102 ) , .ZN( u1_u8_u0_n114 ) , .A1( u1_u8_u0_n92 ) );
  NOR2_X1 u1_u8_u0_U31 (.A1( u1_u8_u0_n120 ) , .ZN( u1_u8_u0_n143 ) , .A2( u1_u8_u0_n167 ) );
  OAI221_X1 u1_u8_u0_U32 (.C1( u1_u8_u0_n112 ) , .ZN( u1_u8_u0_n120 ) , .B1( u1_u8_u0_n138 ) , .B2( u1_u8_u0_n141 ) , .C2( u1_u8_u0_n147 ) , .A( u1_u8_u0_n172 ) );
  AOI211_X1 u1_u8_u0_U33 (.B( u1_u8_u0_n115 ) , .A( u1_u8_u0_n116 ) , .C2( u1_u8_u0_n117 ) , .C1( u1_u8_u0_n118 ) , .ZN( u1_u8_u0_n119 ) );
  NAND2_X1 u1_u8_u0_U34 (.A2( u1_u8_u0_n103 ) , .ZN( u1_u8_u0_n140 ) , .A1( u1_u8_u0_n94 ) );
  NAND2_X1 u1_u8_u0_U35 (.A1( u1_u8_u0_n100 ) , .A2( u1_u8_u0_n103 ) , .ZN( u1_u8_u0_n125 ) );
  NAND2_X1 u1_u8_u0_U36 (.A1( u1_u8_u0_n101 ) , .A2( u1_u8_u0_n102 ) , .ZN( u1_u8_u0_n150 ) );
  INV_X1 u1_u8_u0_U37 (.A( u1_u8_u0_n138 ) , .ZN( u1_u8_u0_n160 ) );
  NAND2_X1 u1_u8_u0_U38 (.A2( u1_u8_u0_n100 ) , .A1( u1_u8_u0_n101 ) , .ZN( u1_u8_u0_n139 ) );
  NAND2_X1 u1_u8_u0_U39 (.ZN( u1_u8_u0_n112 ) , .A2( u1_u8_u0_n92 ) , .A1( u1_u8_u0_n93 ) );
  AOI21_X1 u1_u8_u0_U4 (.B1( u1_u8_u0_n114 ) , .ZN( u1_u8_u0_n115 ) , .B2( u1_u8_u0_n129 ) , .A( u1_u8_u0_n161 ) );
  NAND2_X1 u1_u8_u0_U40 (.A1( u1_u8_u0_n101 ) , .ZN( u1_u8_u0_n130 ) , .A2( u1_u8_u0_n94 ) );
  INV_X1 u1_u8_u0_U41 (.ZN( u1_u8_u0_n172 ) , .A( u1_u8_u0_n88 ) );
  OAI222_X1 u1_u8_u0_U42 (.C1( u1_u8_u0_n108 ) , .A1( u1_u8_u0_n125 ) , .B2( u1_u8_u0_n128 ) , .B1( u1_u8_u0_n144 ) , .A2( u1_u8_u0_n158 ) , .C2( u1_u8_u0_n161 ) , .ZN( u1_u8_u0_n88 ) );
  NAND2_X1 u1_u8_u0_U43 (.A2( u1_u8_u0_n101 ) , .ZN( u1_u8_u0_n121 ) , .A1( u1_u8_u0_n93 ) );
  OR3_X1 u1_u8_u0_U44 (.A3( u1_u8_u0_n152 ) , .A2( u1_u8_u0_n153 ) , .A1( u1_u8_u0_n154 ) , .ZN( u1_u8_u0_n155 ) );
  AOI21_X1 u1_u8_u0_U45 (.A( u1_u8_u0_n144 ) , .B2( u1_u8_u0_n145 ) , .B1( u1_u8_u0_n146 ) , .ZN( u1_u8_u0_n154 ) );
  AOI21_X1 u1_u8_u0_U46 (.B2( u1_u8_u0_n150 ) , .B1( u1_u8_u0_n151 ) , .ZN( u1_u8_u0_n152 ) , .A( u1_u8_u0_n158 ) );
  AOI21_X1 u1_u8_u0_U47 (.A( u1_u8_u0_n147 ) , .B2( u1_u8_u0_n148 ) , .B1( u1_u8_u0_n149 ) , .ZN( u1_u8_u0_n153 ) );
  INV_X1 u1_u8_u0_U48 (.ZN( u1_u8_u0_n171 ) , .A( u1_u8_u0_n99 ) );
  OAI211_X1 u1_u8_u0_U49 (.C2( u1_u8_u0_n140 ) , .C1( u1_u8_u0_n161 ) , .A( u1_u8_u0_n169 ) , .B( u1_u8_u0_n98 ) , .ZN( u1_u8_u0_n99 ) );
  AOI21_X1 u1_u8_u0_U5 (.B2( u1_u8_u0_n131 ) , .ZN( u1_u8_u0_n134 ) , .B1( u1_u8_u0_n151 ) , .A( u1_u8_u0_n158 ) );
  INV_X1 u1_u8_u0_U50 (.ZN( u1_u8_u0_n169 ) , .A( u1_u8_u0_n91 ) );
  AOI211_X1 u1_u8_u0_U51 (.C1( u1_u8_u0_n118 ) , .A( u1_u8_u0_n123 ) , .B( u1_u8_u0_n96 ) , .C2( u1_u8_u0_n97 ) , .ZN( u1_u8_u0_n98 ) );
  NOR2_X1 u1_u8_u0_U52 (.A2( u1_u8_X_4 ) , .A1( u1_u8_X_5 ) , .ZN( u1_u8_u0_n118 ) );
  NOR2_X1 u1_u8_u0_U53 (.A2( u1_u8_X_1 ) , .ZN( u1_u8_u0_n101 ) , .A1( u1_u8_u0_n163 ) );
  NOR2_X1 u1_u8_u0_U54 (.A2( u1_u8_X_3 ) , .A1( u1_u8_X_6 ) , .ZN( u1_u8_u0_n94 ) );
  NOR2_X1 u1_u8_u0_U55 (.A2( u1_u8_X_6 ) , .ZN( u1_u8_u0_n100 ) , .A1( u1_u8_u0_n162 ) );
  NAND2_X1 u1_u8_u0_U56 (.A2( u1_u8_X_4 ) , .A1( u1_u8_X_5 ) , .ZN( u1_u8_u0_n144 ) );
  NOR2_X1 u1_u8_u0_U57 (.A2( u1_u8_X_5 ) , .ZN( u1_u8_u0_n136 ) , .A1( u1_u8_u0_n159 ) );
  NAND2_X1 u1_u8_u0_U58 (.A1( u1_u8_X_5 ) , .ZN( u1_u8_u0_n138 ) , .A2( u1_u8_u0_n159 ) );
  AND2_X1 u1_u8_u0_U59 (.A2( u1_u8_X_3 ) , .A1( u1_u8_X_6 ) , .ZN( u1_u8_u0_n102 ) );
  NOR2_X1 u1_u8_u0_U6 (.A1( u1_u8_u0_n108 ) , .ZN( u1_u8_u0_n123 ) , .A2( u1_u8_u0_n158 ) );
  AND2_X1 u1_u8_u0_U60 (.A1( u1_u8_X_6 ) , .A2( u1_u8_u0_n162 ) , .ZN( u1_u8_u0_n93 ) );
  INV_X1 u1_u8_u0_U61 (.A( u1_u8_X_4 ) , .ZN( u1_u8_u0_n159 ) );
  INV_X1 u1_u8_u0_U62 (.A( u1_u8_X_1 ) , .ZN( u1_u8_u0_n164 ) );
  INV_X1 u1_u8_u0_U63 (.A( u1_u8_X_3 ) , .ZN( u1_u8_u0_n162 ) );
  INV_X1 u1_u8_u0_U64 (.A( u1_u8_u0_n126 ) , .ZN( u1_u8_u0_n168 ) );
  AOI211_X1 u1_u8_u0_U65 (.B( u1_u8_u0_n133 ) , .A( u1_u8_u0_n134 ) , .C2( u1_u8_u0_n135 ) , .C1( u1_u8_u0_n136 ) , .ZN( u1_u8_u0_n137 ) );
  OR4_X1 u1_u8_u0_U66 (.ZN( u1_out8_17 ) , .A4( u1_u8_u0_n122 ) , .A2( u1_u8_u0_n123 ) , .A1( u1_u8_u0_n124 ) , .A3( u1_u8_u0_n170 ) );
  AOI21_X1 u1_u8_u0_U67 (.B2( u1_u8_u0_n107 ) , .ZN( u1_u8_u0_n124 ) , .B1( u1_u8_u0_n128 ) , .A( u1_u8_u0_n161 ) );
  INV_X1 u1_u8_u0_U68 (.A( u1_u8_u0_n111 ) , .ZN( u1_u8_u0_n170 ) );
  OR4_X1 u1_u8_u0_U69 (.ZN( u1_out8_31 ) , .A4( u1_u8_u0_n155 ) , .A2( u1_u8_u0_n156 ) , .A1( u1_u8_u0_n157 ) , .A3( u1_u8_u0_n173 ) );
  OAI21_X1 u1_u8_u0_U7 (.B1( u1_u8_u0_n150 ) , .B2( u1_u8_u0_n158 ) , .A( u1_u8_u0_n172 ) , .ZN( u1_u8_u0_n89 ) );
  AOI21_X1 u1_u8_u0_U70 (.A( u1_u8_u0_n138 ) , .B2( u1_u8_u0_n139 ) , .B1( u1_u8_u0_n140 ) , .ZN( u1_u8_u0_n157 ) );
  AOI211_X1 u1_u8_u0_U71 (.B( u1_u8_u0_n104 ) , .A( u1_u8_u0_n105 ) , .ZN( u1_u8_u0_n106 ) , .C2( u1_u8_u0_n113 ) , .C1( u1_u8_u0_n160 ) );
  INV_X1 u1_u8_u0_U72 (.ZN( u1_u8_u0_n174 ) , .A( u1_u8_u0_n89 ) );
  AOI21_X1 u1_u8_u0_U73 (.B2( u1_u8_u0_n141 ) , .B1( u1_u8_u0_n142 ) , .ZN( u1_u8_u0_n156 ) , .A( u1_u8_u0_n161 ) );
  AOI21_X1 u1_u8_u0_U74 (.ZN( u1_u8_u0_n116 ) , .B2( u1_u8_u0_n142 ) , .A( u1_u8_u0_n144 ) , .B1( u1_u8_u0_n166 ) );
  INV_X1 u1_u8_u0_U75 (.A( u1_u8_u0_n142 ) , .ZN( u1_u8_u0_n165 ) );
  NOR2_X1 u1_u8_u0_U76 (.A2( u1_u8_X_1 ) , .A1( u1_u8_X_2 ) , .ZN( u1_u8_u0_n92 ) );
  NOR2_X1 u1_u8_u0_U77 (.A2( u1_u8_X_2 ) , .ZN( u1_u8_u0_n103 ) , .A1( u1_u8_u0_n164 ) );
  INV_X1 u1_u8_u0_U78 (.A( u1_u8_X_2 ) , .ZN( u1_u8_u0_n163 ) );
  OAI221_X1 u1_u8_u0_U79 (.C1( u1_u8_u0_n121 ) , .ZN( u1_u8_u0_n122 ) , .B2( u1_u8_u0_n127 ) , .A( u1_u8_u0_n143 ) , .B1( u1_u8_u0_n144 ) , .C2( u1_u8_u0_n147 ) );
  AND2_X1 u1_u8_u0_U8 (.A1( u1_u8_u0_n114 ) , .A2( u1_u8_u0_n121 ) , .ZN( u1_u8_u0_n146 ) );
  AOI21_X1 u1_u8_u0_U80 (.B1( u1_u8_u0_n132 ) , .ZN( u1_u8_u0_n133 ) , .A( u1_u8_u0_n144 ) , .B2( u1_u8_u0_n166 ) );
  OAI22_X1 u1_u8_u0_U81 (.ZN( u1_u8_u0_n105 ) , .A2( u1_u8_u0_n132 ) , .B1( u1_u8_u0_n146 ) , .A1( u1_u8_u0_n147 ) , .B2( u1_u8_u0_n161 ) );
  NAND2_X1 u1_u8_u0_U82 (.ZN( u1_u8_u0_n110 ) , .A2( u1_u8_u0_n132 ) , .A1( u1_u8_u0_n145 ) );
  INV_X1 u1_u8_u0_U83 (.A( u1_u8_u0_n119 ) , .ZN( u1_u8_u0_n167 ) );
  NAND2_X1 u1_u8_u0_U84 (.ZN( u1_u8_u0_n148 ) , .A1( u1_u8_u0_n93 ) , .A2( u1_u8_u0_n95 ) );
  NAND2_X1 u1_u8_u0_U85 (.A1( u1_u8_u0_n100 ) , .ZN( u1_u8_u0_n129 ) , .A2( u1_u8_u0_n95 ) );
  NAND2_X1 u1_u8_u0_U86 (.A1( u1_u8_u0_n102 ) , .ZN( u1_u8_u0_n128 ) , .A2( u1_u8_u0_n95 ) );
  NAND2_X1 u1_u8_u0_U87 (.ZN( u1_u8_u0_n142 ) , .A1( u1_u8_u0_n94 ) , .A2( u1_u8_u0_n95 ) );
  NAND3_X1 u1_u8_u0_U88 (.ZN( u1_out8_23 ) , .A3( u1_u8_u0_n137 ) , .A1( u1_u8_u0_n168 ) , .A2( u1_u8_u0_n171 ) );
  NAND3_X1 u1_u8_u0_U89 (.A3( u1_u8_u0_n127 ) , .A2( u1_u8_u0_n128 ) , .ZN( u1_u8_u0_n135 ) , .A1( u1_u8_u0_n150 ) );
  NAND2_X1 u1_u8_u0_U9 (.ZN( u1_u8_u0_n113 ) , .A1( u1_u8_u0_n139 ) , .A2( u1_u8_u0_n149 ) );
  NAND3_X1 u1_u8_u0_U90 (.ZN( u1_u8_u0_n117 ) , .A3( u1_u8_u0_n132 ) , .A2( u1_u8_u0_n139 ) , .A1( u1_u8_u0_n148 ) );
  NAND3_X1 u1_u8_u0_U91 (.ZN( u1_u8_u0_n109 ) , .A2( u1_u8_u0_n114 ) , .A3( u1_u8_u0_n140 ) , .A1( u1_u8_u0_n149 ) );
  NAND3_X1 u1_u8_u0_U92 (.ZN( u1_out8_9 ) , .A3( u1_u8_u0_n106 ) , .A2( u1_u8_u0_n171 ) , .A1( u1_u8_u0_n174 ) );
  NAND3_X1 u1_u8_u0_U93 (.A2( u1_u8_u0_n128 ) , .A1( u1_u8_u0_n132 ) , .A3( u1_u8_u0_n146 ) , .ZN( u1_u8_u0_n97 ) );
  XOR2_X1 u1_u9_U1 (.B( u1_K10_9 ) , .A( u1_R8_6 ) , .Z( u1_u9_X_9 ) );
  XOR2_X1 u1_u9_U15 (.B( u1_K10_40 ) , .A( u1_R8_27 ) , .Z( u1_u9_X_40 ) );
  XOR2_X1 u1_u9_U17 (.B( u1_K10_39 ) , .A( u1_R8_26 ) , .Z( u1_u9_X_39 ) );
  XOR2_X1 u1_u9_U18 (.B( u1_K10_38 ) , .A( u1_R8_25 ) , .Z( u1_u9_X_38 ) );
  XOR2_X1 u1_u9_U19 (.B( u1_K10_37 ) , .A( u1_R8_24 ) , .Z( u1_u9_X_37 ) );
  XOR2_X1 u1_u9_U20 (.B( u1_K10_36 ) , .A( u1_R8_25 ) , .Z( u1_u9_X_36 ) );
  XOR2_X1 u1_u9_U21 (.B( u1_K10_35 ) , .A( u1_R8_24 ) , .Z( u1_u9_X_35 ) );
  XOR2_X1 u1_u9_U22 (.B( u1_K10_34 ) , .A( u1_R8_23 ) , .Z( u1_u9_X_34 ) );
  XOR2_X1 u1_u9_U23 (.B( u1_K10_33 ) , .A( u1_R8_22 ) , .Z( u1_u9_X_33 ) );
  XOR2_X1 u1_u9_U35 (.B( u1_K10_22 ) , .A( u1_R8_15 ) , .Z( u1_u9_X_22 ) );
  XOR2_X1 u1_u9_U36 (.B( u1_K10_21 ) , .A( u1_R8_14 ) , .Z( u1_u9_X_21 ) );
  XOR2_X1 u1_u9_U37 (.B( u1_K10_20 ) , .A( u1_R8_13 ) , .Z( u1_u9_X_20 ) );
  XOR2_X1 u1_u9_U39 (.B( u1_K10_19 ) , .A( u1_R8_12 ) , .Z( u1_u9_X_19 ) );
  XOR2_X1 u1_u9_U40 (.B( u1_K10_18 ) , .A( u1_R8_13 ) , .Z( u1_u9_X_18 ) );
  XOR2_X1 u1_u9_U41 (.B( u1_K10_17 ) , .A( u1_R8_12 ) , .Z( u1_u9_X_17 ) );
  XOR2_X1 u1_u9_U42 (.B( u1_K10_16 ) , .A( u1_R8_11 ) , .Z( u1_u9_X_16 ) );
  XOR2_X1 u1_u9_U43 (.B( u1_K10_15 ) , .A( u1_R8_10 ) , .Z( u1_u9_X_15 ) );
  XOR2_X1 u1_u9_U44 (.B( u1_K10_14 ) , .A( u1_R8_9 ) , .Z( u1_u9_X_14 ) );
  XOR2_X1 u1_u9_U45 (.B( u1_K10_13 ) , .A( u1_R8_8 ) , .Z( u1_u9_X_13 ) );
  XOR2_X1 u1_u9_U46 (.B( u1_K10_12 ) , .A( u1_R8_9 ) , .Z( u1_u9_X_12 ) );
  XOR2_X1 u1_u9_U47 (.B( u1_K10_11 ) , .A( u1_R8_8 ) , .Z( u1_u9_X_11 ) );
  XOR2_X1 u1_u9_U48 (.B( u1_K10_10 ) , .A( u1_R8_7 ) , .Z( u1_u9_X_10 ) );
  NOR2_X1 u1_u9_u1_U10 (.A1( u1_u9_u1_n112 ) , .A2( u1_u9_u1_n116 ) , .ZN( u1_u9_u1_n118 ) );
  NAND3_X1 u1_u9_u1_U100 (.ZN( u1_u9_u1_n113 ) , .A1( u1_u9_u1_n120 ) , .A3( u1_u9_u1_n133 ) , .A2( u1_u9_u1_n155 ) );
  OAI21_X1 u1_u9_u1_U11 (.ZN( u1_u9_u1_n101 ) , .B1( u1_u9_u1_n141 ) , .A( u1_u9_u1_n146 ) , .B2( u1_u9_u1_n183 ) );
  AOI21_X1 u1_u9_u1_U12 (.B2( u1_u9_u1_n155 ) , .B1( u1_u9_u1_n156 ) , .ZN( u1_u9_u1_n157 ) , .A( u1_u9_u1_n174 ) );
  NAND2_X1 u1_u9_u1_U13 (.ZN( u1_u9_u1_n140 ) , .A2( u1_u9_u1_n150 ) , .A1( u1_u9_u1_n155 ) );
  NAND2_X1 u1_u9_u1_U14 (.A1( u1_u9_u1_n131 ) , .ZN( u1_u9_u1_n147 ) , .A2( u1_u9_u1_n153 ) );
  INV_X1 u1_u9_u1_U15 (.A( u1_u9_u1_n139 ) , .ZN( u1_u9_u1_n174 ) );
  OR4_X1 u1_u9_u1_U16 (.A4( u1_u9_u1_n106 ) , .A3( u1_u9_u1_n107 ) , .ZN( u1_u9_u1_n108 ) , .A1( u1_u9_u1_n117 ) , .A2( u1_u9_u1_n184 ) );
  AOI21_X1 u1_u9_u1_U17 (.ZN( u1_u9_u1_n106 ) , .A( u1_u9_u1_n112 ) , .B1( u1_u9_u1_n154 ) , .B2( u1_u9_u1_n156 ) );
  AOI21_X1 u1_u9_u1_U18 (.ZN( u1_u9_u1_n107 ) , .B1( u1_u9_u1_n134 ) , .B2( u1_u9_u1_n149 ) , .A( u1_u9_u1_n174 ) );
  INV_X1 u1_u9_u1_U19 (.A( u1_u9_u1_n101 ) , .ZN( u1_u9_u1_n184 ) );
  INV_X1 u1_u9_u1_U20 (.A( u1_u9_u1_n112 ) , .ZN( u1_u9_u1_n171 ) );
  NAND2_X1 u1_u9_u1_U21 (.ZN( u1_u9_u1_n141 ) , .A1( u1_u9_u1_n153 ) , .A2( u1_u9_u1_n156 ) );
  AND2_X1 u1_u9_u1_U22 (.A1( u1_u9_u1_n123 ) , .ZN( u1_u9_u1_n134 ) , .A2( u1_u9_u1_n161 ) );
  NAND2_X1 u1_u9_u1_U23 (.A2( u1_u9_u1_n115 ) , .A1( u1_u9_u1_n116 ) , .ZN( u1_u9_u1_n148 ) );
  NAND2_X1 u1_u9_u1_U24 (.A2( u1_u9_u1_n133 ) , .A1( u1_u9_u1_n135 ) , .ZN( u1_u9_u1_n159 ) );
  NAND2_X1 u1_u9_u1_U25 (.A2( u1_u9_u1_n115 ) , .A1( u1_u9_u1_n120 ) , .ZN( u1_u9_u1_n132 ) );
  INV_X1 u1_u9_u1_U26 (.A( u1_u9_u1_n154 ) , .ZN( u1_u9_u1_n178 ) );
  INV_X1 u1_u9_u1_U27 (.A( u1_u9_u1_n151 ) , .ZN( u1_u9_u1_n183 ) );
  AND2_X1 u1_u9_u1_U28 (.A1( u1_u9_u1_n129 ) , .A2( u1_u9_u1_n133 ) , .ZN( u1_u9_u1_n149 ) );
  INV_X1 u1_u9_u1_U29 (.A( u1_u9_u1_n131 ) , .ZN( u1_u9_u1_n180 ) );
  INV_X1 u1_u9_u1_U3 (.A( u1_u9_u1_n159 ) , .ZN( u1_u9_u1_n182 ) );
  OAI221_X1 u1_u9_u1_U30 (.A( u1_u9_u1_n119 ) , .C2( u1_u9_u1_n129 ) , .ZN( u1_u9_u1_n138 ) , .B2( u1_u9_u1_n152 ) , .C1( u1_u9_u1_n174 ) , .B1( u1_u9_u1_n187 ) );
  INV_X1 u1_u9_u1_U31 (.A( u1_u9_u1_n148 ) , .ZN( u1_u9_u1_n187 ) );
  AOI211_X1 u1_u9_u1_U32 (.B( u1_u9_u1_n117 ) , .A( u1_u9_u1_n118 ) , .ZN( u1_u9_u1_n119 ) , .C2( u1_u9_u1_n146 ) , .C1( u1_u9_u1_n159 ) );
  NOR2_X1 u1_u9_u1_U33 (.A1( u1_u9_u1_n168 ) , .A2( u1_u9_u1_n176 ) , .ZN( u1_u9_u1_n98 ) );
  AOI211_X1 u1_u9_u1_U34 (.B( u1_u9_u1_n162 ) , .A( u1_u9_u1_n163 ) , .C2( u1_u9_u1_n164 ) , .ZN( u1_u9_u1_n165 ) , .C1( u1_u9_u1_n171 ) );
  AOI21_X1 u1_u9_u1_U35 (.A( u1_u9_u1_n160 ) , .B2( u1_u9_u1_n161 ) , .ZN( u1_u9_u1_n162 ) , .B1( u1_u9_u1_n182 ) );
  OR2_X1 u1_u9_u1_U36 (.A2( u1_u9_u1_n157 ) , .A1( u1_u9_u1_n158 ) , .ZN( u1_u9_u1_n163 ) );
  NAND2_X1 u1_u9_u1_U37 (.A1( u1_u9_u1_n128 ) , .ZN( u1_u9_u1_n146 ) , .A2( u1_u9_u1_n160 ) );
  NAND2_X1 u1_u9_u1_U38 (.A2( u1_u9_u1_n112 ) , .ZN( u1_u9_u1_n139 ) , .A1( u1_u9_u1_n152 ) );
  NAND2_X1 u1_u9_u1_U39 (.A1( u1_u9_u1_n105 ) , .ZN( u1_u9_u1_n156 ) , .A2( u1_u9_u1_n99 ) );
  AOI221_X1 u1_u9_u1_U4 (.A( u1_u9_u1_n138 ) , .C2( u1_u9_u1_n139 ) , .C1( u1_u9_u1_n140 ) , .B2( u1_u9_u1_n141 ) , .ZN( u1_u9_u1_n142 ) , .B1( u1_u9_u1_n175 ) );
  AOI221_X1 u1_u9_u1_U40 (.B1( u1_u9_u1_n140 ) , .ZN( u1_u9_u1_n167 ) , .B2( u1_u9_u1_n172 ) , .C2( u1_u9_u1_n175 ) , .C1( u1_u9_u1_n178 ) , .A( u1_u9_u1_n188 ) );
  INV_X1 u1_u9_u1_U41 (.ZN( u1_u9_u1_n188 ) , .A( u1_u9_u1_n97 ) );
  AOI211_X1 u1_u9_u1_U42 (.A( u1_u9_u1_n118 ) , .C1( u1_u9_u1_n132 ) , .C2( u1_u9_u1_n139 ) , .B( u1_u9_u1_n96 ) , .ZN( u1_u9_u1_n97 ) );
  AOI21_X1 u1_u9_u1_U43 (.B2( u1_u9_u1_n121 ) , .B1( u1_u9_u1_n135 ) , .A( u1_u9_u1_n152 ) , .ZN( u1_u9_u1_n96 ) );
  NOR2_X1 u1_u9_u1_U44 (.ZN( u1_u9_u1_n117 ) , .A1( u1_u9_u1_n121 ) , .A2( u1_u9_u1_n160 ) );
  OAI21_X1 u1_u9_u1_U45 (.B2( u1_u9_u1_n123 ) , .ZN( u1_u9_u1_n145 ) , .B1( u1_u9_u1_n160 ) , .A( u1_u9_u1_n185 ) );
  INV_X1 u1_u9_u1_U46 (.A( u1_u9_u1_n122 ) , .ZN( u1_u9_u1_n185 ) );
  AOI21_X1 u1_u9_u1_U47 (.B2( u1_u9_u1_n120 ) , .B1( u1_u9_u1_n121 ) , .ZN( u1_u9_u1_n122 ) , .A( u1_u9_u1_n128 ) );
  AOI21_X1 u1_u9_u1_U48 (.A( u1_u9_u1_n128 ) , .B2( u1_u9_u1_n129 ) , .ZN( u1_u9_u1_n130 ) , .B1( u1_u9_u1_n150 ) );
  NAND2_X1 u1_u9_u1_U49 (.ZN( u1_u9_u1_n112 ) , .A1( u1_u9_u1_n169 ) , .A2( u1_u9_u1_n170 ) );
  AOI211_X1 u1_u9_u1_U5 (.ZN( u1_u9_u1_n124 ) , .A( u1_u9_u1_n138 ) , .C2( u1_u9_u1_n139 ) , .B( u1_u9_u1_n145 ) , .C1( u1_u9_u1_n147 ) );
  NAND2_X1 u1_u9_u1_U50 (.ZN( u1_u9_u1_n129 ) , .A2( u1_u9_u1_n95 ) , .A1( u1_u9_u1_n98 ) );
  NAND2_X1 u1_u9_u1_U51 (.A1( u1_u9_u1_n102 ) , .ZN( u1_u9_u1_n154 ) , .A2( u1_u9_u1_n99 ) );
  NAND2_X1 u1_u9_u1_U52 (.A2( u1_u9_u1_n100 ) , .ZN( u1_u9_u1_n135 ) , .A1( u1_u9_u1_n99 ) );
  AOI21_X1 u1_u9_u1_U53 (.A( u1_u9_u1_n152 ) , .B2( u1_u9_u1_n153 ) , .B1( u1_u9_u1_n154 ) , .ZN( u1_u9_u1_n158 ) );
  INV_X1 u1_u9_u1_U54 (.A( u1_u9_u1_n160 ) , .ZN( u1_u9_u1_n175 ) );
  NAND2_X1 u1_u9_u1_U55 (.A1( u1_u9_u1_n100 ) , .ZN( u1_u9_u1_n116 ) , .A2( u1_u9_u1_n95 ) );
  NAND2_X1 u1_u9_u1_U56 (.A1( u1_u9_u1_n102 ) , .ZN( u1_u9_u1_n131 ) , .A2( u1_u9_u1_n95 ) );
  NAND2_X1 u1_u9_u1_U57 (.A2( u1_u9_u1_n104 ) , .ZN( u1_u9_u1_n121 ) , .A1( u1_u9_u1_n98 ) );
  NAND2_X1 u1_u9_u1_U58 (.A1( u1_u9_u1_n103 ) , .ZN( u1_u9_u1_n153 ) , .A2( u1_u9_u1_n98 ) );
  NAND2_X1 u1_u9_u1_U59 (.A2( u1_u9_u1_n104 ) , .A1( u1_u9_u1_n105 ) , .ZN( u1_u9_u1_n133 ) );
  AOI22_X1 u1_u9_u1_U6 (.B2( u1_u9_u1_n136 ) , .A2( u1_u9_u1_n137 ) , .ZN( u1_u9_u1_n143 ) , .A1( u1_u9_u1_n171 ) , .B1( u1_u9_u1_n173 ) );
  NAND2_X1 u1_u9_u1_U60 (.ZN( u1_u9_u1_n150 ) , .A2( u1_u9_u1_n98 ) , .A1( u1_u9_u1_n99 ) );
  NAND2_X1 u1_u9_u1_U61 (.A1( u1_u9_u1_n105 ) , .ZN( u1_u9_u1_n155 ) , .A2( u1_u9_u1_n95 ) );
  OAI21_X1 u1_u9_u1_U62 (.ZN( u1_u9_u1_n109 ) , .B1( u1_u9_u1_n129 ) , .B2( u1_u9_u1_n160 ) , .A( u1_u9_u1_n167 ) );
  NAND2_X1 u1_u9_u1_U63 (.A2( u1_u9_u1_n100 ) , .A1( u1_u9_u1_n103 ) , .ZN( u1_u9_u1_n120 ) );
  NAND2_X1 u1_u9_u1_U64 (.A1( u1_u9_u1_n102 ) , .A2( u1_u9_u1_n104 ) , .ZN( u1_u9_u1_n115 ) );
  NAND2_X1 u1_u9_u1_U65 (.A2( u1_u9_u1_n100 ) , .A1( u1_u9_u1_n104 ) , .ZN( u1_u9_u1_n151 ) );
  NAND2_X1 u1_u9_u1_U66 (.A2( u1_u9_u1_n103 ) , .A1( u1_u9_u1_n105 ) , .ZN( u1_u9_u1_n161 ) );
  INV_X1 u1_u9_u1_U67 (.A( u1_u9_u1_n152 ) , .ZN( u1_u9_u1_n173 ) );
  INV_X1 u1_u9_u1_U68 (.A( u1_u9_u1_n128 ) , .ZN( u1_u9_u1_n172 ) );
  NAND2_X1 u1_u9_u1_U69 (.A2( u1_u9_u1_n102 ) , .A1( u1_u9_u1_n103 ) , .ZN( u1_u9_u1_n123 ) );
  INV_X1 u1_u9_u1_U7 (.A( u1_u9_u1_n147 ) , .ZN( u1_u9_u1_n181 ) );
  NOR2_X1 u1_u9_u1_U70 (.A2( u1_u9_X_7 ) , .A1( u1_u9_X_8 ) , .ZN( u1_u9_u1_n95 ) );
  NOR2_X1 u1_u9_u1_U71 (.A1( u1_u9_X_12 ) , .A2( u1_u9_X_9 ) , .ZN( u1_u9_u1_n100 ) );
  NOR2_X1 u1_u9_u1_U72 (.A2( u1_u9_X_8 ) , .A1( u1_u9_u1_n177 ) , .ZN( u1_u9_u1_n99 ) );
  NOR2_X1 u1_u9_u1_U73 (.A2( u1_u9_X_12 ) , .ZN( u1_u9_u1_n102 ) , .A1( u1_u9_u1_n176 ) );
  NOR2_X1 u1_u9_u1_U74 (.A2( u1_u9_X_9 ) , .ZN( u1_u9_u1_n105 ) , .A1( u1_u9_u1_n168 ) );
  NAND2_X1 u1_u9_u1_U75 (.A1( u1_u9_X_10 ) , .ZN( u1_u9_u1_n160 ) , .A2( u1_u9_u1_n169 ) );
  NAND2_X1 u1_u9_u1_U76 (.A2( u1_u9_X_10 ) , .A1( u1_u9_X_11 ) , .ZN( u1_u9_u1_n152 ) );
  NAND2_X1 u1_u9_u1_U77 (.A1( u1_u9_X_11 ) , .ZN( u1_u9_u1_n128 ) , .A2( u1_u9_u1_n170 ) );
  AND2_X1 u1_u9_u1_U78 (.A2( u1_u9_X_7 ) , .A1( u1_u9_X_8 ) , .ZN( u1_u9_u1_n104 ) );
  AND2_X1 u1_u9_u1_U79 (.A1( u1_u9_X_8 ) , .ZN( u1_u9_u1_n103 ) , .A2( u1_u9_u1_n177 ) );
  AOI22_X1 u1_u9_u1_U8 (.B2( u1_u9_u1_n113 ) , .A2( u1_u9_u1_n114 ) , .ZN( u1_u9_u1_n125 ) , .A1( u1_u9_u1_n171 ) , .B1( u1_u9_u1_n173 ) );
  INV_X1 u1_u9_u1_U80 (.A( u1_u9_X_10 ) , .ZN( u1_u9_u1_n170 ) );
  INV_X1 u1_u9_u1_U81 (.A( u1_u9_X_9 ) , .ZN( u1_u9_u1_n176 ) );
  INV_X1 u1_u9_u1_U82 (.A( u1_u9_X_11 ) , .ZN( u1_u9_u1_n169 ) );
  INV_X1 u1_u9_u1_U83 (.A( u1_u9_X_12 ) , .ZN( u1_u9_u1_n168 ) );
  INV_X1 u1_u9_u1_U84 (.A( u1_u9_X_7 ) , .ZN( u1_u9_u1_n177 ) );
  NAND4_X1 u1_u9_u1_U85 (.ZN( u1_out9_18 ) , .A4( u1_u9_u1_n165 ) , .A3( u1_u9_u1_n166 ) , .A1( u1_u9_u1_n167 ) , .A2( u1_u9_u1_n186 ) );
  AOI22_X1 u1_u9_u1_U86 (.B2( u1_u9_u1_n146 ) , .B1( u1_u9_u1_n147 ) , .A2( u1_u9_u1_n148 ) , .ZN( u1_u9_u1_n166 ) , .A1( u1_u9_u1_n172 ) );
  INV_X1 u1_u9_u1_U87 (.A( u1_u9_u1_n145 ) , .ZN( u1_u9_u1_n186 ) );
  NAND4_X1 u1_u9_u1_U88 (.ZN( u1_out9_2 ) , .A4( u1_u9_u1_n142 ) , .A3( u1_u9_u1_n143 ) , .A2( u1_u9_u1_n144 ) , .A1( u1_u9_u1_n179 ) );
  OAI21_X1 u1_u9_u1_U89 (.B2( u1_u9_u1_n132 ) , .ZN( u1_u9_u1_n144 ) , .A( u1_u9_u1_n146 ) , .B1( u1_u9_u1_n180 ) );
  NAND2_X1 u1_u9_u1_U9 (.ZN( u1_u9_u1_n114 ) , .A1( u1_u9_u1_n134 ) , .A2( u1_u9_u1_n156 ) );
  INV_X1 u1_u9_u1_U90 (.A( u1_u9_u1_n130 ) , .ZN( u1_u9_u1_n179 ) );
  NAND4_X1 u1_u9_u1_U91 (.ZN( u1_out9_28 ) , .A4( u1_u9_u1_n124 ) , .A3( u1_u9_u1_n125 ) , .A2( u1_u9_u1_n126 ) , .A1( u1_u9_u1_n127 ) );
  OAI21_X1 u1_u9_u1_U92 (.ZN( u1_u9_u1_n127 ) , .B2( u1_u9_u1_n139 ) , .B1( u1_u9_u1_n175 ) , .A( u1_u9_u1_n183 ) );
  OAI21_X1 u1_u9_u1_U93 (.ZN( u1_u9_u1_n126 ) , .B2( u1_u9_u1_n140 ) , .A( u1_u9_u1_n146 ) , .B1( u1_u9_u1_n178 ) );
  OR4_X1 u1_u9_u1_U94 (.ZN( u1_out9_13 ) , .A4( u1_u9_u1_n108 ) , .A3( u1_u9_u1_n109 ) , .A2( u1_u9_u1_n110 ) , .A1( u1_u9_u1_n111 ) );
  AOI21_X1 u1_u9_u1_U95 (.ZN( u1_u9_u1_n110 ) , .A( u1_u9_u1_n116 ) , .B1( u1_u9_u1_n152 ) , .B2( u1_u9_u1_n160 ) );
  AOI21_X1 u1_u9_u1_U96 (.ZN( u1_u9_u1_n111 ) , .A( u1_u9_u1_n128 ) , .B2( u1_u9_u1_n131 ) , .B1( u1_u9_u1_n135 ) );
  NAND3_X1 u1_u9_u1_U97 (.A3( u1_u9_u1_n149 ) , .A2( u1_u9_u1_n150 ) , .A1( u1_u9_u1_n151 ) , .ZN( u1_u9_u1_n164 ) );
  NAND3_X1 u1_u9_u1_U98 (.A3( u1_u9_u1_n134 ) , .A2( u1_u9_u1_n135 ) , .ZN( u1_u9_u1_n136 ) , .A1( u1_u9_u1_n151 ) );
  NAND3_X1 u1_u9_u1_U99 (.A1( u1_u9_u1_n133 ) , .ZN( u1_u9_u1_n137 ) , .A2( u1_u9_u1_n154 ) , .A3( u1_u9_u1_n181 ) );
  OAI22_X1 u1_u9_u2_U10 (.B1( u1_u9_u2_n151 ) , .A2( u1_u9_u2_n152 ) , .A1( u1_u9_u2_n153 ) , .ZN( u1_u9_u2_n160 ) , .B2( u1_u9_u2_n168 ) );
  NAND3_X1 u1_u9_u2_U100 (.A2( u1_u9_u2_n100 ) , .A1( u1_u9_u2_n104 ) , .A3( u1_u9_u2_n138 ) , .ZN( u1_u9_u2_n98 ) );
  NOR3_X1 u1_u9_u2_U11 (.A1( u1_u9_u2_n150 ) , .ZN( u1_u9_u2_n151 ) , .A3( u1_u9_u2_n175 ) , .A2( u1_u9_u2_n188 ) );
  AOI21_X1 u1_u9_u2_U12 (.B2( u1_u9_u2_n123 ) , .ZN( u1_u9_u2_n125 ) , .A( u1_u9_u2_n171 ) , .B1( u1_u9_u2_n184 ) );
  INV_X1 u1_u9_u2_U13 (.A( u1_u9_u2_n150 ) , .ZN( u1_u9_u2_n184 ) );
  AOI21_X1 u1_u9_u2_U14 (.ZN( u1_u9_u2_n144 ) , .B2( u1_u9_u2_n155 ) , .A( u1_u9_u2_n172 ) , .B1( u1_u9_u2_n185 ) );
  AOI21_X1 u1_u9_u2_U15 (.B2( u1_u9_u2_n143 ) , .ZN( u1_u9_u2_n145 ) , .B1( u1_u9_u2_n152 ) , .A( u1_u9_u2_n171 ) );
  INV_X1 u1_u9_u2_U16 (.A( u1_u9_u2_n156 ) , .ZN( u1_u9_u2_n171 ) );
  INV_X1 u1_u9_u2_U17 (.A( u1_u9_u2_n120 ) , .ZN( u1_u9_u2_n188 ) );
  NAND2_X1 u1_u9_u2_U18 (.A2( u1_u9_u2_n122 ) , .ZN( u1_u9_u2_n150 ) , .A1( u1_u9_u2_n152 ) );
  INV_X1 u1_u9_u2_U19 (.A( u1_u9_u2_n153 ) , .ZN( u1_u9_u2_n170 ) );
  INV_X1 u1_u9_u2_U20 (.A( u1_u9_u2_n137 ) , .ZN( u1_u9_u2_n173 ) );
  NAND2_X1 u1_u9_u2_U21 (.A1( u1_u9_u2_n132 ) , .A2( u1_u9_u2_n139 ) , .ZN( u1_u9_u2_n157 ) );
  INV_X1 u1_u9_u2_U22 (.A( u1_u9_u2_n113 ) , .ZN( u1_u9_u2_n178 ) );
  INV_X1 u1_u9_u2_U23 (.A( u1_u9_u2_n139 ) , .ZN( u1_u9_u2_n175 ) );
  INV_X1 u1_u9_u2_U24 (.A( u1_u9_u2_n155 ) , .ZN( u1_u9_u2_n181 ) );
  INV_X1 u1_u9_u2_U25 (.A( u1_u9_u2_n119 ) , .ZN( u1_u9_u2_n177 ) );
  INV_X1 u1_u9_u2_U26 (.A( u1_u9_u2_n116 ) , .ZN( u1_u9_u2_n180 ) );
  INV_X1 u1_u9_u2_U27 (.A( u1_u9_u2_n131 ) , .ZN( u1_u9_u2_n179 ) );
  INV_X1 u1_u9_u2_U28 (.A( u1_u9_u2_n154 ) , .ZN( u1_u9_u2_n176 ) );
  NAND2_X1 u1_u9_u2_U29 (.A2( u1_u9_u2_n116 ) , .A1( u1_u9_u2_n117 ) , .ZN( u1_u9_u2_n118 ) );
  NOR2_X1 u1_u9_u2_U3 (.ZN( u1_u9_u2_n121 ) , .A2( u1_u9_u2_n177 ) , .A1( u1_u9_u2_n180 ) );
  INV_X1 u1_u9_u2_U30 (.A( u1_u9_u2_n132 ) , .ZN( u1_u9_u2_n182 ) );
  INV_X1 u1_u9_u2_U31 (.A( u1_u9_u2_n158 ) , .ZN( u1_u9_u2_n183 ) );
  OAI21_X1 u1_u9_u2_U32 (.A( u1_u9_u2_n156 ) , .B1( u1_u9_u2_n157 ) , .ZN( u1_u9_u2_n158 ) , .B2( u1_u9_u2_n179 ) );
  NOR2_X1 u1_u9_u2_U33 (.ZN( u1_u9_u2_n156 ) , .A1( u1_u9_u2_n166 ) , .A2( u1_u9_u2_n169 ) );
  NOR2_X1 u1_u9_u2_U34 (.A2( u1_u9_u2_n114 ) , .ZN( u1_u9_u2_n137 ) , .A1( u1_u9_u2_n140 ) );
  NOR2_X1 u1_u9_u2_U35 (.A2( u1_u9_u2_n138 ) , .ZN( u1_u9_u2_n153 ) , .A1( u1_u9_u2_n156 ) );
  AOI211_X1 u1_u9_u2_U36 (.ZN( u1_u9_u2_n130 ) , .C1( u1_u9_u2_n138 ) , .C2( u1_u9_u2_n179 ) , .B( u1_u9_u2_n96 ) , .A( u1_u9_u2_n97 ) );
  OAI22_X1 u1_u9_u2_U37 (.B1( u1_u9_u2_n133 ) , .A2( u1_u9_u2_n137 ) , .A1( u1_u9_u2_n152 ) , .B2( u1_u9_u2_n168 ) , .ZN( u1_u9_u2_n97 ) );
  OAI221_X1 u1_u9_u2_U38 (.B1( u1_u9_u2_n113 ) , .C1( u1_u9_u2_n132 ) , .A( u1_u9_u2_n149 ) , .B2( u1_u9_u2_n171 ) , .C2( u1_u9_u2_n172 ) , .ZN( u1_u9_u2_n96 ) );
  OAI221_X1 u1_u9_u2_U39 (.A( u1_u9_u2_n115 ) , .C2( u1_u9_u2_n123 ) , .B2( u1_u9_u2_n143 ) , .B1( u1_u9_u2_n153 ) , .ZN( u1_u9_u2_n163 ) , .C1( u1_u9_u2_n168 ) );
  INV_X1 u1_u9_u2_U4 (.A( u1_u9_u2_n134 ) , .ZN( u1_u9_u2_n185 ) );
  OAI21_X1 u1_u9_u2_U40 (.A( u1_u9_u2_n114 ) , .ZN( u1_u9_u2_n115 ) , .B1( u1_u9_u2_n176 ) , .B2( u1_u9_u2_n178 ) );
  OAI221_X1 u1_u9_u2_U41 (.A( u1_u9_u2_n135 ) , .B2( u1_u9_u2_n136 ) , .B1( u1_u9_u2_n137 ) , .ZN( u1_u9_u2_n162 ) , .C2( u1_u9_u2_n167 ) , .C1( u1_u9_u2_n185 ) );
  AND3_X1 u1_u9_u2_U42 (.A3( u1_u9_u2_n131 ) , .A2( u1_u9_u2_n132 ) , .A1( u1_u9_u2_n133 ) , .ZN( u1_u9_u2_n136 ) );
  AOI22_X1 u1_u9_u2_U43 (.ZN( u1_u9_u2_n135 ) , .B1( u1_u9_u2_n140 ) , .A1( u1_u9_u2_n156 ) , .B2( u1_u9_u2_n180 ) , .A2( u1_u9_u2_n188 ) );
  AOI21_X1 u1_u9_u2_U44 (.ZN( u1_u9_u2_n149 ) , .B1( u1_u9_u2_n173 ) , .B2( u1_u9_u2_n188 ) , .A( u1_u9_u2_n95 ) );
  AND3_X1 u1_u9_u2_U45 (.A2( u1_u9_u2_n100 ) , .A1( u1_u9_u2_n104 ) , .A3( u1_u9_u2_n156 ) , .ZN( u1_u9_u2_n95 ) );
  OAI21_X1 u1_u9_u2_U46 (.A( u1_u9_u2_n101 ) , .B2( u1_u9_u2_n121 ) , .B1( u1_u9_u2_n153 ) , .ZN( u1_u9_u2_n164 ) );
  NAND2_X1 u1_u9_u2_U47 (.A2( u1_u9_u2_n100 ) , .A1( u1_u9_u2_n107 ) , .ZN( u1_u9_u2_n155 ) );
  NAND2_X1 u1_u9_u2_U48 (.A2( u1_u9_u2_n105 ) , .A1( u1_u9_u2_n108 ) , .ZN( u1_u9_u2_n143 ) );
  NAND2_X1 u1_u9_u2_U49 (.A1( u1_u9_u2_n104 ) , .A2( u1_u9_u2_n106 ) , .ZN( u1_u9_u2_n152 ) );
  NOR4_X1 u1_u9_u2_U5 (.A4( u1_u9_u2_n124 ) , .A3( u1_u9_u2_n125 ) , .A2( u1_u9_u2_n126 ) , .A1( u1_u9_u2_n127 ) , .ZN( u1_u9_u2_n128 ) );
  NAND2_X1 u1_u9_u2_U50 (.A1( u1_u9_u2_n100 ) , .A2( u1_u9_u2_n105 ) , .ZN( u1_u9_u2_n132 ) );
  INV_X1 u1_u9_u2_U51 (.A( u1_u9_u2_n140 ) , .ZN( u1_u9_u2_n168 ) );
  INV_X1 u1_u9_u2_U52 (.A( u1_u9_u2_n138 ) , .ZN( u1_u9_u2_n167 ) );
  OAI21_X1 u1_u9_u2_U53 (.A( u1_u9_u2_n141 ) , .B2( u1_u9_u2_n142 ) , .ZN( u1_u9_u2_n146 ) , .B1( u1_u9_u2_n153 ) );
  OAI21_X1 u1_u9_u2_U54 (.A( u1_u9_u2_n140 ) , .ZN( u1_u9_u2_n141 ) , .B1( u1_u9_u2_n176 ) , .B2( u1_u9_u2_n177 ) );
  NOR3_X1 u1_u9_u2_U55 (.ZN( u1_u9_u2_n142 ) , .A3( u1_u9_u2_n175 ) , .A2( u1_u9_u2_n178 ) , .A1( u1_u9_u2_n181 ) );
  NAND2_X1 u1_u9_u2_U56 (.A1( u1_u9_u2_n102 ) , .A2( u1_u9_u2_n106 ) , .ZN( u1_u9_u2_n113 ) );
  NAND2_X1 u1_u9_u2_U57 (.A1( u1_u9_u2_n106 ) , .A2( u1_u9_u2_n107 ) , .ZN( u1_u9_u2_n131 ) );
  NAND2_X1 u1_u9_u2_U58 (.A1( u1_u9_u2_n103 ) , .A2( u1_u9_u2_n107 ) , .ZN( u1_u9_u2_n139 ) );
  NAND2_X1 u1_u9_u2_U59 (.A1( u1_u9_u2_n103 ) , .A2( u1_u9_u2_n105 ) , .ZN( u1_u9_u2_n133 ) );
  AOI21_X1 u1_u9_u2_U6 (.B2( u1_u9_u2_n119 ) , .ZN( u1_u9_u2_n127 ) , .A( u1_u9_u2_n137 ) , .B1( u1_u9_u2_n155 ) );
  NAND2_X1 u1_u9_u2_U60 (.A1( u1_u9_u2_n102 ) , .A2( u1_u9_u2_n103 ) , .ZN( u1_u9_u2_n154 ) );
  NAND2_X1 u1_u9_u2_U61 (.A2( u1_u9_u2_n103 ) , .A1( u1_u9_u2_n104 ) , .ZN( u1_u9_u2_n119 ) );
  NAND2_X1 u1_u9_u2_U62 (.A2( u1_u9_u2_n107 ) , .A1( u1_u9_u2_n108 ) , .ZN( u1_u9_u2_n123 ) );
  NAND2_X1 u1_u9_u2_U63 (.A1( u1_u9_u2_n104 ) , .A2( u1_u9_u2_n108 ) , .ZN( u1_u9_u2_n122 ) );
  INV_X1 u1_u9_u2_U64 (.A( u1_u9_u2_n114 ) , .ZN( u1_u9_u2_n172 ) );
  NAND2_X1 u1_u9_u2_U65 (.A2( u1_u9_u2_n100 ) , .A1( u1_u9_u2_n102 ) , .ZN( u1_u9_u2_n116 ) );
  NAND2_X1 u1_u9_u2_U66 (.A1( u1_u9_u2_n102 ) , .A2( u1_u9_u2_n108 ) , .ZN( u1_u9_u2_n120 ) );
  NAND2_X1 u1_u9_u2_U67 (.A2( u1_u9_u2_n105 ) , .A1( u1_u9_u2_n106 ) , .ZN( u1_u9_u2_n117 ) );
  INV_X1 u1_u9_u2_U68 (.ZN( u1_u9_u2_n187 ) , .A( u1_u9_u2_n99 ) );
  OAI21_X1 u1_u9_u2_U69 (.B1( u1_u9_u2_n137 ) , .B2( u1_u9_u2_n143 ) , .A( u1_u9_u2_n98 ) , .ZN( u1_u9_u2_n99 ) );
  AOI21_X1 u1_u9_u2_U7 (.ZN( u1_u9_u2_n124 ) , .B1( u1_u9_u2_n131 ) , .B2( u1_u9_u2_n143 ) , .A( u1_u9_u2_n172 ) );
  NOR2_X1 u1_u9_u2_U70 (.A2( u1_u9_X_16 ) , .ZN( u1_u9_u2_n140 ) , .A1( u1_u9_u2_n166 ) );
  NOR2_X1 u1_u9_u2_U71 (.A2( u1_u9_X_13 ) , .A1( u1_u9_X_14 ) , .ZN( u1_u9_u2_n100 ) );
  NOR2_X1 u1_u9_u2_U72 (.A2( u1_u9_X_16 ) , .A1( u1_u9_X_17 ) , .ZN( u1_u9_u2_n138 ) );
  NOR2_X1 u1_u9_u2_U73 (.A2( u1_u9_X_15 ) , .A1( u1_u9_X_18 ) , .ZN( u1_u9_u2_n104 ) );
  NOR2_X1 u1_u9_u2_U74 (.A2( u1_u9_X_14 ) , .ZN( u1_u9_u2_n103 ) , .A1( u1_u9_u2_n174 ) );
  NOR2_X1 u1_u9_u2_U75 (.A2( u1_u9_X_15 ) , .ZN( u1_u9_u2_n102 ) , .A1( u1_u9_u2_n165 ) );
  NOR2_X1 u1_u9_u2_U76 (.A2( u1_u9_X_17 ) , .ZN( u1_u9_u2_n114 ) , .A1( u1_u9_u2_n169 ) );
  AND2_X1 u1_u9_u2_U77 (.A1( u1_u9_X_15 ) , .ZN( u1_u9_u2_n105 ) , .A2( u1_u9_u2_n165 ) );
  AND2_X1 u1_u9_u2_U78 (.A2( u1_u9_X_15 ) , .A1( u1_u9_X_18 ) , .ZN( u1_u9_u2_n107 ) );
  AND2_X1 u1_u9_u2_U79 (.A1( u1_u9_X_14 ) , .ZN( u1_u9_u2_n106 ) , .A2( u1_u9_u2_n174 ) );
  AOI21_X1 u1_u9_u2_U8 (.B2( u1_u9_u2_n120 ) , .B1( u1_u9_u2_n121 ) , .ZN( u1_u9_u2_n126 ) , .A( u1_u9_u2_n167 ) );
  AND2_X1 u1_u9_u2_U80 (.A1( u1_u9_X_13 ) , .A2( u1_u9_X_14 ) , .ZN( u1_u9_u2_n108 ) );
  INV_X1 u1_u9_u2_U81 (.A( u1_u9_X_16 ) , .ZN( u1_u9_u2_n169 ) );
  INV_X1 u1_u9_u2_U82 (.A( u1_u9_X_17 ) , .ZN( u1_u9_u2_n166 ) );
  INV_X1 u1_u9_u2_U83 (.A( u1_u9_X_13 ) , .ZN( u1_u9_u2_n174 ) );
  INV_X1 u1_u9_u2_U84 (.A( u1_u9_X_18 ) , .ZN( u1_u9_u2_n165 ) );
  NAND4_X1 u1_u9_u2_U85 (.ZN( u1_out9_24 ) , .A4( u1_u9_u2_n111 ) , .A3( u1_u9_u2_n112 ) , .A1( u1_u9_u2_n130 ) , .A2( u1_u9_u2_n187 ) );
  AOI221_X1 u1_u9_u2_U86 (.A( u1_u9_u2_n109 ) , .B1( u1_u9_u2_n110 ) , .ZN( u1_u9_u2_n111 ) , .C1( u1_u9_u2_n134 ) , .C2( u1_u9_u2_n170 ) , .B2( u1_u9_u2_n173 ) );
  AOI21_X1 u1_u9_u2_U87 (.ZN( u1_u9_u2_n112 ) , .B2( u1_u9_u2_n156 ) , .A( u1_u9_u2_n164 ) , .B1( u1_u9_u2_n181 ) );
  NAND4_X1 u1_u9_u2_U88 (.ZN( u1_out9_16 ) , .A4( u1_u9_u2_n128 ) , .A3( u1_u9_u2_n129 ) , .A1( u1_u9_u2_n130 ) , .A2( u1_u9_u2_n186 ) );
  AOI22_X1 u1_u9_u2_U89 (.A2( u1_u9_u2_n118 ) , .ZN( u1_u9_u2_n129 ) , .A1( u1_u9_u2_n140 ) , .B1( u1_u9_u2_n157 ) , .B2( u1_u9_u2_n170 ) );
  OAI22_X1 u1_u9_u2_U9 (.ZN( u1_u9_u2_n109 ) , .A2( u1_u9_u2_n113 ) , .B2( u1_u9_u2_n133 ) , .B1( u1_u9_u2_n167 ) , .A1( u1_u9_u2_n168 ) );
  INV_X1 u1_u9_u2_U90 (.A( u1_u9_u2_n163 ) , .ZN( u1_u9_u2_n186 ) );
  NAND4_X1 u1_u9_u2_U91 (.ZN( u1_out9_30 ) , .A4( u1_u9_u2_n147 ) , .A3( u1_u9_u2_n148 ) , .A2( u1_u9_u2_n149 ) , .A1( u1_u9_u2_n187 ) );
  AOI21_X1 u1_u9_u2_U92 (.B2( u1_u9_u2_n138 ) , .ZN( u1_u9_u2_n148 ) , .A( u1_u9_u2_n162 ) , .B1( u1_u9_u2_n182 ) );
  NOR3_X1 u1_u9_u2_U93 (.A3( u1_u9_u2_n144 ) , .A2( u1_u9_u2_n145 ) , .A1( u1_u9_u2_n146 ) , .ZN( u1_u9_u2_n147 ) );
  OR4_X1 u1_u9_u2_U94 (.ZN( u1_out9_6 ) , .A4( u1_u9_u2_n161 ) , .A3( u1_u9_u2_n162 ) , .A2( u1_u9_u2_n163 ) , .A1( u1_u9_u2_n164 ) );
  OR3_X1 u1_u9_u2_U95 (.A2( u1_u9_u2_n159 ) , .A1( u1_u9_u2_n160 ) , .ZN( u1_u9_u2_n161 ) , .A3( u1_u9_u2_n183 ) );
  AOI21_X1 u1_u9_u2_U96 (.B2( u1_u9_u2_n154 ) , .B1( u1_u9_u2_n155 ) , .ZN( u1_u9_u2_n159 ) , .A( u1_u9_u2_n167 ) );
  NAND3_X1 u1_u9_u2_U97 (.A2( u1_u9_u2_n117 ) , .A1( u1_u9_u2_n122 ) , .A3( u1_u9_u2_n123 ) , .ZN( u1_u9_u2_n134 ) );
  NAND3_X1 u1_u9_u2_U98 (.ZN( u1_u9_u2_n110 ) , .A2( u1_u9_u2_n131 ) , .A3( u1_u9_u2_n139 ) , .A1( u1_u9_u2_n154 ) );
  NAND3_X1 u1_u9_u2_U99 (.A2( u1_u9_u2_n100 ) , .ZN( u1_u9_u2_n101 ) , .A1( u1_u9_u2_n104 ) , .A3( u1_u9_u2_n114 ) );
  OAI22_X1 u1_u9_u3_U10 (.B1( u1_u9_u3_n113 ) , .A2( u1_u9_u3_n135 ) , .A1( u1_u9_u3_n150 ) , .B2( u1_u9_u3_n164 ) , .ZN( u1_u9_u3_n98 ) );
  OAI211_X1 u1_u9_u3_U11 (.B( u1_u9_u3_n106 ) , .ZN( u1_u9_u3_n119 ) , .C2( u1_u9_u3_n128 ) , .C1( u1_u9_u3_n167 ) , .A( u1_u9_u3_n181 ) );
  AOI221_X1 u1_u9_u3_U12 (.C1( u1_u9_u3_n105 ) , .ZN( u1_u9_u3_n106 ) , .A( u1_u9_u3_n131 ) , .B2( u1_u9_u3_n132 ) , .C2( u1_u9_u3_n133 ) , .B1( u1_u9_u3_n169 ) );
  INV_X1 u1_u9_u3_U13 (.ZN( u1_u9_u3_n181 ) , .A( u1_u9_u3_n98 ) );
  NAND2_X1 u1_u9_u3_U14 (.ZN( u1_u9_u3_n105 ) , .A2( u1_u9_u3_n130 ) , .A1( u1_u9_u3_n155 ) );
  AOI22_X1 u1_u9_u3_U15 (.B1( u1_u9_u3_n115 ) , .A2( u1_u9_u3_n116 ) , .ZN( u1_u9_u3_n123 ) , .B2( u1_u9_u3_n133 ) , .A1( u1_u9_u3_n169 ) );
  NAND2_X1 u1_u9_u3_U16 (.ZN( u1_u9_u3_n116 ) , .A2( u1_u9_u3_n151 ) , .A1( u1_u9_u3_n182 ) );
  NOR2_X1 u1_u9_u3_U17 (.ZN( u1_u9_u3_n126 ) , .A2( u1_u9_u3_n150 ) , .A1( u1_u9_u3_n164 ) );
  AOI21_X1 u1_u9_u3_U18 (.ZN( u1_u9_u3_n112 ) , .B2( u1_u9_u3_n146 ) , .B1( u1_u9_u3_n155 ) , .A( u1_u9_u3_n167 ) );
  NAND2_X1 u1_u9_u3_U19 (.A1( u1_u9_u3_n135 ) , .ZN( u1_u9_u3_n142 ) , .A2( u1_u9_u3_n164 ) );
  NAND2_X1 u1_u9_u3_U20 (.ZN( u1_u9_u3_n132 ) , .A2( u1_u9_u3_n152 ) , .A1( u1_u9_u3_n156 ) );
  AND2_X1 u1_u9_u3_U21 (.A2( u1_u9_u3_n113 ) , .A1( u1_u9_u3_n114 ) , .ZN( u1_u9_u3_n151 ) );
  INV_X1 u1_u9_u3_U22 (.A( u1_u9_u3_n133 ) , .ZN( u1_u9_u3_n165 ) );
  INV_X1 u1_u9_u3_U23 (.A( u1_u9_u3_n135 ) , .ZN( u1_u9_u3_n170 ) );
  NAND2_X1 u1_u9_u3_U24 (.A1( u1_u9_u3_n107 ) , .A2( u1_u9_u3_n108 ) , .ZN( u1_u9_u3_n140 ) );
  NAND2_X1 u1_u9_u3_U25 (.ZN( u1_u9_u3_n117 ) , .A1( u1_u9_u3_n124 ) , .A2( u1_u9_u3_n148 ) );
  NAND2_X1 u1_u9_u3_U26 (.ZN( u1_u9_u3_n143 ) , .A1( u1_u9_u3_n165 ) , .A2( u1_u9_u3_n167 ) );
  INV_X1 u1_u9_u3_U27 (.A( u1_u9_u3_n130 ) , .ZN( u1_u9_u3_n177 ) );
  INV_X1 u1_u9_u3_U28 (.A( u1_u9_u3_n128 ) , .ZN( u1_u9_u3_n176 ) );
  INV_X1 u1_u9_u3_U29 (.A( u1_u9_u3_n155 ) , .ZN( u1_u9_u3_n174 ) );
  INV_X1 u1_u9_u3_U3 (.A( u1_u9_u3_n129 ) , .ZN( u1_u9_u3_n183 ) );
  INV_X1 u1_u9_u3_U30 (.A( u1_u9_u3_n139 ) , .ZN( u1_u9_u3_n185 ) );
  NOR2_X1 u1_u9_u3_U31 (.ZN( u1_u9_u3_n135 ) , .A2( u1_u9_u3_n141 ) , .A1( u1_u9_u3_n169 ) );
  OAI222_X1 u1_u9_u3_U32 (.C2( u1_u9_u3_n107 ) , .A2( u1_u9_u3_n108 ) , .B1( u1_u9_u3_n135 ) , .ZN( u1_u9_u3_n138 ) , .B2( u1_u9_u3_n146 ) , .C1( u1_u9_u3_n154 ) , .A1( u1_u9_u3_n164 ) );
  NOR4_X1 u1_u9_u3_U33 (.A4( u1_u9_u3_n157 ) , .A3( u1_u9_u3_n158 ) , .A2( u1_u9_u3_n159 ) , .A1( u1_u9_u3_n160 ) , .ZN( u1_u9_u3_n161 ) );
  AOI21_X1 u1_u9_u3_U34 (.B2( u1_u9_u3_n152 ) , .B1( u1_u9_u3_n153 ) , .ZN( u1_u9_u3_n158 ) , .A( u1_u9_u3_n164 ) );
  AOI21_X1 u1_u9_u3_U35 (.A( u1_u9_u3_n154 ) , .B2( u1_u9_u3_n155 ) , .B1( u1_u9_u3_n156 ) , .ZN( u1_u9_u3_n157 ) );
  AOI21_X1 u1_u9_u3_U36 (.A( u1_u9_u3_n149 ) , .B2( u1_u9_u3_n150 ) , .B1( u1_u9_u3_n151 ) , .ZN( u1_u9_u3_n159 ) );
  AOI211_X1 u1_u9_u3_U37 (.ZN( u1_u9_u3_n109 ) , .A( u1_u9_u3_n119 ) , .C2( u1_u9_u3_n129 ) , .B( u1_u9_u3_n138 ) , .C1( u1_u9_u3_n141 ) );
  AOI211_X1 u1_u9_u3_U38 (.B( u1_u9_u3_n119 ) , .A( u1_u9_u3_n120 ) , .C2( u1_u9_u3_n121 ) , .ZN( u1_u9_u3_n122 ) , .C1( u1_u9_u3_n179 ) );
  INV_X1 u1_u9_u3_U39 (.A( u1_u9_u3_n156 ) , .ZN( u1_u9_u3_n179 ) );
  INV_X1 u1_u9_u3_U4 (.A( u1_u9_u3_n140 ) , .ZN( u1_u9_u3_n182 ) );
  OAI22_X1 u1_u9_u3_U40 (.B1( u1_u9_u3_n118 ) , .ZN( u1_u9_u3_n120 ) , .A1( u1_u9_u3_n135 ) , .B2( u1_u9_u3_n154 ) , .A2( u1_u9_u3_n178 ) );
  AND3_X1 u1_u9_u3_U41 (.ZN( u1_u9_u3_n118 ) , .A2( u1_u9_u3_n124 ) , .A1( u1_u9_u3_n144 ) , .A3( u1_u9_u3_n152 ) );
  INV_X1 u1_u9_u3_U42 (.A( u1_u9_u3_n121 ) , .ZN( u1_u9_u3_n164 ) );
  NAND2_X1 u1_u9_u3_U43 (.ZN( u1_u9_u3_n133 ) , .A1( u1_u9_u3_n154 ) , .A2( u1_u9_u3_n164 ) );
  OAI211_X1 u1_u9_u3_U44 (.B( u1_u9_u3_n127 ) , .ZN( u1_u9_u3_n139 ) , .C1( u1_u9_u3_n150 ) , .C2( u1_u9_u3_n154 ) , .A( u1_u9_u3_n184 ) );
  INV_X1 u1_u9_u3_U45 (.A( u1_u9_u3_n125 ) , .ZN( u1_u9_u3_n184 ) );
  AOI221_X1 u1_u9_u3_U46 (.A( u1_u9_u3_n126 ) , .ZN( u1_u9_u3_n127 ) , .C2( u1_u9_u3_n132 ) , .C1( u1_u9_u3_n169 ) , .B2( u1_u9_u3_n170 ) , .B1( u1_u9_u3_n174 ) );
  OAI22_X1 u1_u9_u3_U47 (.A1( u1_u9_u3_n124 ) , .ZN( u1_u9_u3_n125 ) , .B2( u1_u9_u3_n145 ) , .A2( u1_u9_u3_n165 ) , .B1( u1_u9_u3_n167 ) );
  NOR2_X1 u1_u9_u3_U48 (.A1( u1_u9_u3_n113 ) , .ZN( u1_u9_u3_n131 ) , .A2( u1_u9_u3_n154 ) );
  NAND2_X1 u1_u9_u3_U49 (.A1( u1_u9_u3_n103 ) , .ZN( u1_u9_u3_n150 ) , .A2( u1_u9_u3_n99 ) );
  INV_X1 u1_u9_u3_U5 (.A( u1_u9_u3_n117 ) , .ZN( u1_u9_u3_n178 ) );
  NAND2_X1 u1_u9_u3_U50 (.A2( u1_u9_u3_n102 ) , .ZN( u1_u9_u3_n155 ) , .A1( u1_u9_u3_n97 ) );
  INV_X1 u1_u9_u3_U51 (.A( u1_u9_u3_n141 ) , .ZN( u1_u9_u3_n167 ) );
  AOI21_X1 u1_u9_u3_U52 (.B2( u1_u9_u3_n114 ) , .B1( u1_u9_u3_n146 ) , .A( u1_u9_u3_n154 ) , .ZN( u1_u9_u3_n94 ) );
  AOI21_X1 u1_u9_u3_U53 (.ZN( u1_u9_u3_n110 ) , .B2( u1_u9_u3_n142 ) , .B1( u1_u9_u3_n186 ) , .A( u1_u9_u3_n95 ) );
  INV_X1 u1_u9_u3_U54 (.A( u1_u9_u3_n145 ) , .ZN( u1_u9_u3_n186 ) );
  AOI21_X1 u1_u9_u3_U55 (.B1( u1_u9_u3_n124 ) , .A( u1_u9_u3_n149 ) , .B2( u1_u9_u3_n155 ) , .ZN( u1_u9_u3_n95 ) );
  INV_X1 u1_u9_u3_U56 (.A( u1_u9_u3_n149 ) , .ZN( u1_u9_u3_n169 ) );
  NAND2_X1 u1_u9_u3_U57 (.ZN( u1_u9_u3_n124 ) , .A1( u1_u9_u3_n96 ) , .A2( u1_u9_u3_n97 ) );
  NAND2_X1 u1_u9_u3_U58 (.A2( u1_u9_u3_n100 ) , .ZN( u1_u9_u3_n146 ) , .A1( u1_u9_u3_n96 ) );
  NAND2_X1 u1_u9_u3_U59 (.A1( u1_u9_u3_n101 ) , .ZN( u1_u9_u3_n145 ) , .A2( u1_u9_u3_n99 ) );
  AOI221_X1 u1_u9_u3_U6 (.A( u1_u9_u3_n131 ) , .C2( u1_u9_u3_n132 ) , .C1( u1_u9_u3_n133 ) , .ZN( u1_u9_u3_n134 ) , .B1( u1_u9_u3_n143 ) , .B2( u1_u9_u3_n177 ) );
  NAND2_X1 u1_u9_u3_U60 (.A1( u1_u9_u3_n100 ) , .ZN( u1_u9_u3_n156 ) , .A2( u1_u9_u3_n99 ) );
  NAND2_X1 u1_u9_u3_U61 (.A2( u1_u9_u3_n101 ) , .A1( u1_u9_u3_n104 ) , .ZN( u1_u9_u3_n148 ) );
  NAND2_X1 u1_u9_u3_U62 (.A1( u1_u9_u3_n100 ) , .A2( u1_u9_u3_n102 ) , .ZN( u1_u9_u3_n128 ) );
  NAND2_X1 u1_u9_u3_U63 (.A2( u1_u9_u3_n101 ) , .A1( u1_u9_u3_n102 ) , .ZN( u1_u9_u3_n152 ) );
  NAND2_X1 u1_u9_u3_U64 (.A2( u1_u9_u3_n101 ) , .ZN( u1_u9_u3_n114 ) , .A1( u1_u9_u3_n96 ) );
  NAND2_X1 u1_u9_u3_U65 (.ZN( u1_u9_u3_n107 ) , .A1( u1_u9_u3_n97 ) , .A2( u1_u9_u3_n99 ) );
  NAND2_X1 u1_u9_u3_U66 (.A2( u1_u9_u3_n100 ) , .A1( u1_u9_u3_n104 ) , .ZN( u1_u9_u3_n113 ) );
  NAND2_X1 u1_u9_u3_U67 (.A1( u1_u9_u3_n104 ) , .ZN( u1_u9_u3_n153 ) , .A2( u1_u9_u3_n97 ) );
  NAND2_X1 u1_u9_u3_U68 (.A2( u1_u9_u3_n103 ) , .A1( u1_u9_u3_n104 ) , .ZN( u1_u9_u3_n130 ) );
  NAND2_X1 u1_u9_u3_U69 (.A2( u1_u9_u3_n103 ) , .ZN( u1_u9_u3_n144 ) , .A1( u1_u9_u3_n96 ) );
  OAI22_X1 u1_u9_u3_U7 (.B2( u1_u9_u3_n147 ) , .A2( u1_u9_u3_n148 ) , .ZN( u1_u9_u3_n160 ) , .B1( u1_u9_u3_n165 ) , .A1( u1_u9_u3_n168 ) );
  NAND2_X1 u1_u9_u3_U70 (.A1( u1_u9_u3_n102 ) , .A2( u1_u9_u3_n103 ) , .ZN( u1_u9_u3_n108 ) );
  NOR2_X1 u1_u9_u3_U71 (.A2( u1_u9_X_19 ) , .A1( u1_u9_X_20 ) , .ZN( u1_u9_u3_n99 ) );
  NOR2_X1 u1_u9_u3_U72 (.A2( u1_u9_X_21 ) , .A1( u1_u9_X_24 ) , .ZN( u1_u9_u3_n103 ) );
  NOR2_X1 u1_u9_u3_U73 (.A2( u1_u9_X_24 ) , .A1( u1_u9_u3_n171 ) , .ZN( u1_u9_u3_n97 ) );
  NOR2_X1 u1_u9_u3_U74 (.A2( u1_u9_X_23 ) , .ZN( u1_u9_u3_n141 ) , .A1( u1_u9_u3_n166 ) );
  NOR2_X1 u1_u9_u3_U75 (.A2( u1_u9_X_19 ) , .A1( u1_u9_u3_n172 ) , .ZN( u1_u9_u3_n96 ) );
  NAND2_X1 u1_u9_u3_U76 (.A1( u1_u9_X_22 ) , .A2( u1_u9_X_23 ) , .ZN( u1_u9_u3_n154 ) );
  NAND2_X1 u1_u9_u3_U77 (.A1( u1_u9_X_23 ) , .ZN( u1_u9_u3_n149 ) , .A2( u1_u9_u3_n166 ) );
  NOR2_X1 u1_u9_u3_U78 (.A2( u1_u9_X_22 ) , .A1( u1_u9_X_23 ) , .ZN( u1_u9_u3_n121 ) );
  AND2_X1 u1_u9_u3_U79 (.A1( u1_u9_X_24 ) , .ZN( u1_u9_u3_n101 ) , .A2( u1_u9_u3_n171 ) );
  AND3_X1 u1_u9_u3_U8 (.A3( u1_u9_u3_n144 ) , .A2( u1_u9_u3_n145 ) , .A1( u1_u9_u3_n146 ) , .ZN( u1_u9_u3_n147 ) );
  AND2_X1 u1_u9_u3_U80 (.A1( u1_u9_X_19 ) , .ZN( u1_u9_u3_n102 ) , .A2( u1_u9_u3_n172 ) );
  AND2_X1 u1_u9_u3_U81 (.A1( u1_u9_X_21 ) , .A2( u1_u9_X_24 ) , .ZN( u1_u9_u3_n100 ) );
  AND2_X1 u1_u9_u3_U82 (.A2( u1_u9_X_19 ) , .A1( u1_u9_X_20 ) , .ZN( u1_u9_u3_n104 ) );
  INV_X1 u1_u9_u3_U83 (.A( u1_u9_X_22 ) , .ZN( u1_u9_u3_n166 ) );
  INV_X1 u1_u9_u3_U84 (.A( u1_u9_X_21 ) , .ZN( u1_u9_u3_n171 ) );
  INV_X1 u1_u9_u3_U85 (.A( u1_u9_X_20 ) , .ZN( u1_u9_u3_n172 ) );
  OR4_X1 u1_u9_u3_U86 (.ZN( u1_out9_10 ) , .A4( u1_u9_u3_n136 ) , .A3( u1_u9_u3_n137 ) , .A1( u1_u9_u3_n138 ) , .A2( u1_u9_u3_n139 ) );
  OAI222_X1 u1_u9_u3_U87 (.C1( u1_u9_u3_n128 ) , .ZN( u1_u9_u3_n137 ) , .B1( u1_u9_u3_n148 ) , .A2( u1_u9_u3_n150 ) , .B2( u1_u9_u3_n154 ) , .C2( u1_u9_u3_n164 ) , .A1( u1_u9_u3_n167 ) );
  OAI221_X1 u1_u9_u3_U88 (.A( u1_u9_u3_n134 ) , .B2( u1_u9_u3_n135 ) , .ZN( u1_u9_u3_n136 ) , .C1( u1_u9_u3_n149 ) , .B1( u1_u9_u3_n151 ) , .C2( u1_u9_u3_n183 ) );
  NAND4_X1 u1_u9_u3_U89 (.ZN( u1_out9_26 ) , .A4( u1_u9_u3_n109 ) , .A3( u1_u9_u3_n110 ) , .A2( u1_u9_u3_n111 ) , .A1( u1_u9_u3_n173 ) );
  INV_X1 u1_u9_u3_U9 (.A( u1_u9_u3_n143 ) , .ZN( u1_u9_u3_n168 ) );
  INV_X1 u1_u9_u3_U90 (.ZN( u1_u9_u3_n173 ) , .A( u1_u9_u3_n94 ) );
  OAI21_X1 u1_u9_u3_U91 (.ZN( u1_u9_u3_n111 ) , .B2( u1_u9_u3_n117 ) , .A( u1_u9_u3_n133 ) , .B1( u1_u9_u3_n176 ) );
  NAND4_X1 u1_u9_u3_U92 (.ZN( u1_out9_20 ) , .A4( u1_u9_u3_n122 ) , .A3( u1_u9_u3_n123 ) , .A1( u1_u9_u3_n175 ) , .A2( u1_u9_u3_n180 ) );
  INV_X1 u1_u9_u3_U93 (.A( u1_u9_u3_n126 ) , .ZN( u1_u9_u3_n180 ) );
  INV_X1 u1_u9_u3_U94 (.A( u1_u9_u3_n112 ) , .ZN( u1_u9_u3_n175 ) );
  NAND4_X1 u1_u9_u3_U95 (.ZN( u1_out9_1 ) , .A4( u1_u9_u3_n161 ) , .A3( u1_u9_u3_n162 ) , .A2( u1_u9_u3_n163 ) , .A1( u1_u9_u3_n185 ) );
  NAND2_X1 u1_u9_u3_U96 (.ZN( u1_u9_u3_n163 ) , .A2( u1_u9_u3_n170 ) , .A1( u1_u9_u3_n176 ) );
  AOI22_X1 u1_u9_u3_U97 (.B2( u1_u9_u3_n140 ) , .B1( u1_u9_u3_n141 ) , .A2( u1_u9_u3_n142 ) , .ZN( u1_u9_u3_n162 ) , .A1( u1_u9_u3_n177 ) );
  NAND3_X1 u1_u9_u3_U98 (.A1( u1_u9_u3_n114 ) , .ZN( u1_u9_u3_n115 ) , .A2( u1_u9_u3_n145 ) , .A3( u1_u9_u3_n153 ) );
  NAND3_X1 u1_u9_u3_U99 (.ZN( u1_u9_u3_n129 ) , .A2( u1_u9_u3_n144 ) , .A1( u1_u9_u3_n153 ) , .A3( u1_u9_u3_n182 ) );
  NOR2_X1 u1_u9_u5_U10 (.ZN( u1_u9_u5_n135 ) , .A1( u1_u9_u5_n173 ) , .A2( u1_u9_u5_n176 ) );
  NOR3_X1 u1_u9_u5_U100 (.A3( u1_u9_u5_n141 ) , .A1( u1_u9_u5_n142 ) , .ZN( u1_u9_u5_n143 ) , .A2( u1_u9_u5_n191 ) );
  NAND4_X1 u1_u9_u5_U101 (.ZN( u1_out9_4 ) , .A4( u1_u9_u5_n112 ) , .A2( u1_u9_u5_n113 ) , .A1( u1_u9_u5_n114 ) , .A3( u1_u9_u5_n195 ) );
  AOI211_X1 u1_u9_u5_U102 (.A( u1_u9_u5_n110 ) , .C1( u1_u9_u5_n111 ) , .ZN( u1_u9_u5_n112 ) , .B( u1_u9_u5_n118 ) , .C2( u1_u9_u5_n177 ) );
  INV_X1 u1_u9_u5_U103 (.A( u1_u9_u5_n102 ) , .ZN( u1_u9_u5_n195 ) );
  NAND3_X1 u1_u9_u5_U104 (.A2( u1_u9_u5_n154 ) , .A3( u1_u9_u5_n158 ) , .A1( u1_u9_u5_n161 ) , .ZN( u1_u9_u5_n99 ) );
  INV_X1 u1_u9_u5_U11 (.A( u1_u9_u5_n121 ) , .ZN( u1_u9_u5_n177 ) );
  NOR2_X1 u1_u9_u5_U12 (.ZN( u1_u9_u5_n160 ) , .A2( u1_u9_u5_n173 ) , .A1( u1_u9_u5_n177 ) );
  INV_X1 u1_u9_u5_U13 (.A( u1_u9_u5_n150 ) , .ZN( u1_u9_u5_n174 ) );
  AOI21_X1 u1_u9_u5_U14 (.A( u1_u9_u5_n160 ) , .B2( u1_u9_u5_n161 ) , .ZN( u1_u9_u5_n162 ) , .B1( u1_u9_u5_n192 ) );
  INV_X1 u1_u9_u5_U15 (.A( u1_u9_u5_n159 ) , .ZN( u1_u9_u5_n192 ) );
  AOI21_X1 u1_u9_u5_U16 (.A( u1_u9_u5_n156 ) , .B2( u1_u9_u5_n157 ) , .B1( u1_u9_u5_n158 ) , .ZN( u1_u9_u5_n163 ) );
  AOI21_X1 u1_u9_u5_U17 (.B2( u1_u9_u5_n139 ) , .B1( u1_u9_u5_n140 ) , .ZN( u1_u9_u5_n141 ) , .A( u1_u9_u5_n150 ) );
  OAI21_X1 u1_u9_u5_U18 (.A( u1_u9_u5_n133 ) , .B2( u1_u9_u5_n134 ) , .B1( u1_u9_u5_n135 ) , .ZN( u1_u9_u5_n142 ) );
  OAI21_X1 u1_u9_u5_U19 (.ZN( u1_u9_u5_n133 ) , .B2( u1_u9_u5_n147 ) , .A( u1_u9_u5_n173 ) , .B1( u1_u9_u5_n188 ) );
  NAND2_X1 u1_u9_u5_U20 (.A2( u1_u9_u5_n119 ) , .A1( u1_u9_u5_n123 ) , .ZN( u1_u9_u5_n137 ) );
  INV_X1 u1_u9_u5_U21 (.A( u1_u9_u5_n155 ) , .ZN( u1_u9_u5_n194 ) );
  NAND2_X1 u1_u9_u5_U22 (.A1( u1_u9_u5_n121 ) , .ZN( u1_u9_u5_n132 ) , .A2( u1_u9_u5_n172 ) );
  NAND2_X1 u1_u9_u5_U23 (.A2( u1_u9_u5_n122 ) , .ZN( u1_u9_u5_n136 ) , .A1( u1_u9_u5_n154 ) );
  NAND2_X1 u1_u9_u5_U24 (.A2( u1_u9_u5_n119 ) , .A1( u1_u9_u5_n120 ) , .ZN( u1_u9_u5_n159 ) );
  INV_X1 u1_u9_u5_U25 (.A( u1_u9_u5_n156 ) , .ZN( u1_u9_u5_n175 ) );
  INV_X1 u1_u9_u5_U26 (.A( u1_u9_u5_n158 ) , .ZN( u1_u9_u5_n188 ) );
  INV_X1 u1_u9_u5_U27 (.A( u1_u9_u5_n152 ) , .ZN( u1_u9_u5_n179 ) );
  INV_X1 u1_u9_u5_U28 (.A( u1_u9_u5_n140 ) , .ZN( u1_u9_u5_n182 ) );
  INV_X1 u1_u9_u5_U29 (.A( u1_u9_u5_n151 ) , .ZN( u1_u9_u5_n183 ) );
  NOR2_X1 u1_u9_u5_U3 (.ZN( u1_u9_u5_n134 ) , .A1( u1_u9_u5_n183 ) , .A2( u1_u9_u5_n190 ) );
  INV_X1 u1_u9_u5_U30 (.A( u1_u9_u5_n123 ) , .ZN( u1_u9_u5_n185 ) );
  INV_X1 u1_u9_u5_U31 (.A( u1_u9_u5_n161 ) , .ZN( u1_u9_u5_n184 ) );
  INV_X1 u1_u9_u5_U32 (.A( u1_u9_u5_n139 ) , .ZN( u1_u9_u5_n189 ) );
  INV_X1 u1_u9_u5_U33 (.A( u1_u9_u5_n157 ) , .ZN( u1_u9_u5_n190 ) );
  INV_X1 u1_u9_u5_U34 (.A( u1_u9_u5_n120 ) , .ZN( u1_u9_u5_n193 ) );
  NAND2_X1 u1_u9_u5_U35 (.ZN( u1_u9_u5_n111 ) , .A1( u1_u9_u5_n140 ) , .A2( u1_u9_u5_n155 ) );
  NOR2_X1 u1_u9_u5_U36 (.ZN( u1_u9_u5_n100 ) , .A1( u1_u9_u5_n170 ) , .A2( u1_u9_u5_n180 ) );
  INV_X1 u1_u9_u5_U37 (.A( u1_u9_u5_n117 ) , .ZN( u1_u9_u5_n196 ) );
  OAI221_X1 u1_u9_u5_U38 (.A( u1_u9_u5_n116 ) , .ZN( u1_u9_u5_n117 ) , .B2( u1_u9_u5_n119 ) , .C1( u1_u9_u5_n153 ) , .C2( u1_u9_u5_n158 ) , .B1( u1_u9_u5_n172 ) );
  AOI222_X1 u1_u9_u5_U39 (.ZN( u1_u9_u5_n116 ) , .B2( u1_u9_u5_n145 ) , .C1( u1_u9_u5_n148 ) , .A2( u1_u9_u5_n174 ) , .C2( u1_u9_u5_n177 ) , .B1( u1_u9_u5_n187 ) , .A1( u1_u9_u5_n193 ) );
  INV_X1 u1_u9_u5_U4 (.A( u1_u9_u5_n138 ) , .ZN( u1_u9_u5_n191 ) );
  INV_X1 u1_u9_u5_U40 (.A( u1_u9_u5_n115 ) , .ZN( u1_u9_u5_n187 ) );
  OAI221_X1 u1_u9_u5_U41 (.A( u1_u9_u5_n101 ) , .ZN( u1_u9_u5_n102 ) , .C2( u1_u9_u5_n115 ) , .C1( u1_u9_u5_n126 ) , .B1( u1_u9_u5_n134 ) , .B2( u1_u9_u5_n160 ) );
  OAI21_X1 u1_u9_u5_U42 (.ZN( u1_u9_u5_n101 ) , .B1( u1_u9_u5_n137 ) , .A( u1_u9_u5_n146 ) , .B2( u1_u9_u5_n147 ) );
  AOI22_X1 u1_u9_u5_U43 (.B2( u1_u9_u5_n131 ) , .A2( u1_u9_u5_n146 ) , .ZN( u1_u9_u5_n169 ) , .B1( u1_u9_u5_n174 ) , .A1( u1_u9_u5_n185 ) );
  NOR2_X1 u1_u9_u5_U44 (.A1( u1_u9_u5_n146 ) , .ZN( u1_u9_u5_n150 ) , .A2( u1_u9_u5_n173 ) );
  AOI21_X1 u1_u9_u5_U45 (.A( u1_u9_u5_n118 ) , .B2( u1_u9_u5_n145 ) , .ZN( u1_u9_u5_n168 ) , .B1( u1_u9_u5_n186 ) );
  INV_X1 u1_u9_u5_U46 (.A( u1_u9_u5_n122 ) , .ZN( u1_u9_u5_n186 ) );
  NOR2_X1 u1_u9_u5_U47 (.A1( u1_u9_u5_n146 ) , .ZN( u1_u9_u5_n152 ) , .A2( u1_u9_u5_n176 ) );
  NOR2_X1 u1_u9_u5_U48 (.A1( u1_u9_u5_n115 ) , .ZN( u1_u9_u5_n118 ) , .A2( u1_u9_u5_n153 ) );
  NOR2_X1 u1_u9_u5_U49 (.A2( u1_u9_u5_n145 ) , .ZN( u1_u9_u5_n156 ) , .A1( u1_u9_u5_n174 ) );
  OAI21_X1 u1_u9_u5_U5 (.B2( u1_u9_u5_n136 ) , .B1( u1_u9_u5_n137 ) , .ZN( u1_u9_u5_n138 ) , .A( u1_u9_u5_n177 ) );
  NOR2_X1 u1_u9_u5_U50 (.ZN( u1_u9_u5_n121 ) , .A2( u1_u9_u5_n145 ) , .A1( u1_u9_u5_n176 ) );
  AOI22_X1 u1_u9_u5_U51 (.ZN( u1_u9_u5_n114 ) , .A2( u1_u9_u5_n137 ) , .A1( u1_u9_u5_n145 ) , .B2( u1_u9_u5_n175 ) , .B1( u1_u9_u5_n193 ) );
  OAI211_X1 u1_u9_u5_U52 (.B( u1_u9_u5_n124 ) , .A( u1_u9_u5_n125 ) , .C2( u1_u9_u5_n126 ) , .C1( u1_u9_u5_n127 ) , .ZN( u1_u9_u5_n128 ) );
  NOR3_X1 u1_u9_u5_U53 (.ZN( u1_u9_u5_n127 ) , .A1( u1_u9_u5_n136 ) , .A3( u1_u9_u5_n148 ) , .A2( u1_u9_u5_n182 ) );
  OAI21_X1 u1_u9_u5_U54 (.ZN( u1_u9_u5_n124 ) , .A( u1_u9_u5_n177 ) , .B2( u1_u9_u5_n183 ) , .B1( u1_u9_u5_n189 ) );
  OAI21_X1 u1_u9_u5_U55 (.ZN( u1_u9_u5_n125 ) , .A( u1_u9_u5_n174 ) , .B2( u1_u9_u5_n185 ) , .B1( u1_u9_u5_n190 ) );
  AOI21_X1 u1_u9_u5_U56 (.A( u1_u9_u5_n153 ) , .B2( u1_u9_u5_n154 ) , .B1( u1_u9_u5_n155 ) , .ZN( u1_u9_u5_n164 ) );
  AOI21_X1 u1_u9_u5_U57 (.ZN( u1_u9_u5_n110 ) , .B1( u1_u9_u5_n122 ) , .B2( u1_u9_u5_n139 ) , .A( u1_u9_u5_n153 ) );
  INV_X1 u1_u9_u5_U58 (.A( u1_u9_u5_n153 ) , .ZN( u1_u9_u5_n176 ) );
  INV_X1 u1_u9_u5_U59 (.A( u1_u9_u5_n126 ) , .ZN( u1_u9_u5_n173 ) );
  AOI222_X1 u1_u9_u5_U6 (.ZN( u1_u9_u5_n113 ) , .A1( u1_u9_u5_n131 ) , .C1( u1_u9_u5_n148 ) , .B2( u1_u9_u5_n174 ) , .C2( u1_u9_u5_n178 ) , .A2( u1_u9_u5_n179 ) , .B1( u1_u9_u5_n99 ) );
  AND2_X1 u1_u9_u5_U60 (.A2( u1_u9_u5_n104 ) , .A1( u1_u9_u5_n107 ) , .ZN( u1_u9_u5_n147 ) );
  AND2_X1 u1_u9_u5_U61 (.A2( u1_u9_u5_n104 ) , .A1( u1_u9_u5_n108 ) , .ZN( u1_u9_u5_n148 ) );
  NAND2_X1 u1_u9_u5_U62 (.A1( u1_u9_u5_n105 ) , .A2( u1_u9_u5_n106 ) , .ZN( u1_u9_u5_n158 ) );
  NAND2_X1 u1_u9_u5_U63 (.A2( u1_u9_u5_n108 ) , .A1( u1_u9_u5_n109 ) , .ZN( u1_u9_u5_n139 ) );
  NAND2_X1 u1_u9_u5_U64 (.A1( u1_u9_u5_n106 ) , .A2( u1_u9_u5_n108 ) , .ZN( u1_u9_u5_n119 ) );
  NAND2_X1 u1_u9_u5_U65 (.A2( u1_u9_u5_n103 ) , .A1( u1_u9_u5_n105 ) , .ZN( u1_u9_u5_n140 ) );
  NAND2_X1 u1_u9_u5_U66 (.A2( u1_u9_u5_n104 ) , .A1( u1_u9_u5_n105 ) , .ZN( u1_u9_u5_n155 ) );
  NAND2_X1 u1_u9_u5_U67 (.A2( u1_u9_u5_n106 ) , .A1( u1_u9_u5_n107 ) , .ZN( u1_u9_u5_n122 ) );
  NAND2_X1 u1_u9_u5_U68 (.A2( u1_u9_u5_n100 ) , .A1( u1_u9_u5_n106 ) , .ZN( u1_u9_u5_n115 ) );
  NAND2_X1 u1_u9_u5_U69 (.A2( u1_u9_u5_n100 ) , .A1( u1_u9_u5_n103 ) , .ZN( u1_u9_u5_n161 ) );
  INV_X1 u1_u9_u5_U7 (.A( u1_u9_u5_n135 ) , .ZN( u1_u9_u5_n178 ) );
  NAND2_X1 u1_u9_u5_U70 (.A1( u1_u9_u5_n105 ) , .A2( u1_u9_u5_n109 ) , .ZN( u1_u9_u5_n154 ) );
  INV_X1 u1_u9_u5_U71 (.A( u1_u9_u5_n146 ) , .ZN( u1_u9_u5_n172 ) );
  NAND2_X1 u1_u9_u5_U72 (.A1( u1_u9_u5_n103 ) , .A2( u1_u9_u5_n108 ) , .ZN( u1_u9_u5_n123 ) );
  NAND2_X1 u1_u9_u5_U73 (.A2( u1_u9_u5_n103 ) , .A1( u1_u9_u5_n107 ) , .ZN( u1_u9_u5_n151 ) );
  NAND2_X1 u1_u9_u5_U74 (.A2( u1_u9_u5_n107 ) , .A1( u1_u9_u5_n109 ) , .ZN( u1_u9_u5_n120 ) );
  NAND2_X1 u1_u9_u5_U75 (.A2( u1_u9_u5_n100 ) , .A1( u1_u9_u5_n109 ) , .ZN( u1_u9_u5_n157 ) );
  AND2_X1 u1_u9_u5_U76 (.A2( u1_u9_u5_n100 ) , .A1( u1_u9_u5_n104 ) , .ZN( u1_u9_u5_n131 ) );
  NOR2_X1 u1_u9_u5_U77 (.A2( u1_u9_X_34 ) , .A1( u1_u9_X_35 ) , .ZN( u1_u9_u5_n145 ) );
  NOR2_X1 u1_u9_u5_U78 (.A2( u1_u9_X_34 ) , .ZN( u1_u9_u5_n146 ) , .A1( u1_u9_u5_n171 ) );
  NOR2_X1 u1_u9_u5_U79 (.A2( u1_u9_X_31 ) , .A1( u1_u9_X_32 ) , .ZN( u1_u9_u5_n103 ) );
  OAI22_X1 u1_u9_u5_U8 (.B2( u1_u9_u5_n149 ) , .B1( u1_u9_u5_n150 ) , .A2( u1_u9_u5_n151 ) , .A1( u1_u9_u5_n152 ) , .ZN( u1_u9_u5_n165 ) );
  NOR2_X1 u1_u9_u5_U80 (.A2( u1_u9_X_36 ) , .ZN( u1_u9_u5_n105 ) , .A1( u1_u9_u5_n180 ) );
  NOR2_X1 u1_u9_u5_U81 (.A2( u1_u9_X_33 ) , .ZN( u1_u9_u5_n108 ) , .A1( u1_u9_u5_n170 ) );
  NOR2_X1 u1_u9_u5_U82 (.A2( u1_u9_X_33 ) , .A1( u1_u9_X_36 ) , .ZN( u1_u9_u5_n107 ) );
  NOR2_X1 u1_u9_u5_U83 (.A2( u1_u9_X_31 ) , .ZN( u1_u9_u5_n104 ) , .A1( u1_u9_u5_n181 ) );
  NAND2_X1 u1_u9_u5_U84 (.A2( u1_u9_X_34 ) , .A1( u1_u9_X_35 ) , .ZN( u1_u9_u5_n153 ) );
  NAND2_X1 u1_u9_u5_U85 (.A1( u1_u9_X_34 ) , .ZN( u1_u9_u5_n126 ) , .A2( u1_u9_u5_n171 ) );
  AND2_X1 u1_u9_u5_U86 (.A1( u1_u9_X_31 ) , .A2( u1_u9_X_32 ) , .ZN( u1_u9_u5_n106 ) );
  AND2_X1 u1_u9_u5_U87 (.A1( u1_u9_X_31 ) , .ZN( u1_u9_u5_n109 ) , .A2( u1_u9_u5_n181 ) );
  INV_X1 u1_u9_u5_U88 (.A( u1_u9_X_33 ) , .ZN( u1_u9_u5_n180 ) );
  INV_X1 u1_u9_u5_U89 (.A( u1_u9_X_35 ) , .ZN( u1_u9_u5_n171 ) );
  NOR3_X1 u1_u9_u5_U9 (.A2( u1_u9_u5_n147 ) , .A1( u1_u9_u5_n148 ) , .ZN( u1_u9_u5_n149 ) , .A3( u1_u9_u5_n194 ) );
  INV_X1 u1_u9_u5_U90 (.A( u1_u9_X_36 ) , .ZN( u1_u9_u5_n170 ) );
  INV_X1 u1_u9_u5_U91 (.A( u1_u9_X_32 ) , .ZN( u1_u9_u5_n181 ) );
  NAND4_X1 u1_u9_u5_U92 (.ZN( u1_out9_29 ) , .A4( u1_u9_u5_n129 ) , .A3( u1_u9_u5_n130 ) , .A2( u1_u9_u5_n168 ) , .A1( u1_u9_u5_n196 ) );
  AOI221_X1 u1_u9_u5_U93 (.A( u1_u9_u5_n128 ) , .ZN( u1_u9_u5_n129 ) , .C2( u1_u9_u5_n132 ) , .B2( u1_u9_u5_n159 ) , .B1( u1_u9_u5_n176 ) , .C1( u1_u9_u5_n184 ) );
  AOI222_X1 u1_u9_u5_U94 (.ZN( u1_u9_u5_n130 ) , .A2( u1_u9_u5_n146 ) , .B1( u1_u9_u5_n147 ) , .C2( u1_u9_u5_n175 ) , .B2( u1_u9_u5_n179 ) , .A1( u1_u9_u5_n188 ) , .C1( u1_u9_u5_n194 ) );
  NAND4_X1 u1_u9_u5_U95 (.ZN( u1_out9_19 ) , .A4( u1_u9_u5_n166 ) , .A3( u1_u9_u5_n167 ) , .A2( u1_u9_u5_n168 ) , .A1( u1_u9_u5_n169 ) );
  AOI22_X1 u1_u9_u5_U96 (.B2( u1_u9_u5_n145 ) , .A2( u1_u9_u5_n146 ) , .ZN( u1_u9_u5_n167 ) , .B1( u1_u9_u5_n182 ) , .A1( u1_u9_u5_n189 ) );
  NOR4_X1 u1_u9_u5_U97 (.A4( u1_u9_u5_n162 ) , .A3( u1_u9_u5_n163 ) , .A2( u1_u9_u5_n164 ) , .A1( u1_u9_u5_n165 ) , .ZN( u1_u9_u5_n166 ) );
  NAND4_X1 u1_u9_u5_U98 (.ZN( u1_out9_11 ) , .A4( u1_u9_u5_n143 ) , .A3( u1_u9_u5_n144 ) , .A2( u1_u9_u5_n169 ) , .A1( u1_u9_u5_n196 ) );
  AOI22_X1 u1_u9_u5_U99 (.A2( u1_u9_u5_n132 ) , .ZN( u1_u9_u5_n144 ) , .B2( u1_u9_u5_n145 ) , .B1( u1_u9_u5_n184 ) , .A1( u1_u9_u5_n194 ) );
  AOI22_X1 u1_u9_u6_U10 (.A2( u1_u9_u6_n151 ) , .B2( u1_u9_u6_n161 ) , .A1( u1_u9_u6_n167 ) , .B1( u1_u9_u6_n170 ) , .ZN( u1_u9_u6_n89 ) );
  AOI21_X1 u1_u9_u6_U11 (.B1( u1_u9_u6_n107 ) , .B2( u1_u9_u6_n132 ) , .A( u1_u9_u6_n158 ) , .ZN( u1_u9_u6_n88 ) );
  AOI21_X1 u1_u9_u6_U12 (.B2( u1_u9_u6_n147 ) , .B1( u1_u9_u6_n148 ) , .ZN( u1_u9_u6_n149 ) , .A( u1_u9_u6_n158 ) );
  AOI21_X1 u1_u9_u6_U13 (.ZN( u1_u9_u6_n106 ) , .A( u1_u9_u6_n142 ) , .B2( u1_u9_u6_n159 ) , .B1( u1_u9_u6_n164 ) );
  INV_X1 u1_u9_u6_U14 (.A( u1_u9_u6_n155 ) , .ZN( u1_u9_u6_n161 ) );
  INV_X1 u1_u9_u6_U15 (.A( u1_u9_u6_n128 ) , .ZN( u1_u9_u6_n164 ) );
  NAND2_X1 u1_u9_u6_U16 (.ZN( u1_u9_u6_n110 ) , .A1( u1_u9_u6_n122 ) , .A2( u1_u9_u6_n129 ) );
  NAND2_X1 u1_u9_u6_U17 (.ZN( u1_u9_u6_n124 ) , .A2( u1_u9_u6_n146 ) , .A1( u1_u9_u6_n148 ) );
  INV_X1 u1_u9_u6_U18 (.A( u1_u9_u6_n132 ) , .ZN( u1_u9_u6_n171 ) );
  AND2_X1 u1_u9_u6_U19 (.A1( u1_u9_u6_n100 ) , .ZN( u1_u9_u6_n130 ) , .A2( u1_u9_u6_n147 ) );
  INV_X1 u1_u9_u6_U20 (.A( u1_u9_u6_n127 ) , .ZN( u1_u9_u6_n173 ) );
  INV_X1 u1_u9_u6_U21 (.A( u1_u9_u6_n121 ) , .ZN( u1_u9_u6_n167 ) );
  INV_X1 u1_u9_u6_U22 (.A( u1_u9_u6_n100 ) , .ZN( u1_u9_u6_n169 ) );
  INV_X1 u1_u9_u6_U23 (.A( u1_u9_u6_n123 ) , .ZN( u1_u9_u6_n170 ) );
  INV_X1 u1_u9_u6_U24 (.A( u1_u9_u6_n113 ) , .ZN( u1_u9_u6_n168 ) );
  AND2_X1 u1_u9_u6_U25 (.A1( u1_u9_u6_n107 ) , .A2( u1_u9_u6_n119 ) , .ZN( u1_u9_u6_n133 ) );
  AND2_X1 u1_u9_u6_U26 (.A2( u1_u9_u6_n121 ) , .A1( u1_u9_u6_n122 ) , .ZN( u1_u9_u6_n131 ) );
  AND3_X1 u1_u9_u6_U27 (.ZN( u1_u9_u6_n120 ) , .A2( u1_u9_u6_n127 ) , .A1( u1_u9_u6_n132 ) , .A3( u1_u9_u6_n145 ) );
  INV_X1 u1_u9_u6_U28 (.A( u1_u9_u6_n146 ) , .ZN( u1_u9_u6_n163 ) );
  AOI222_X1 u1_u9_u6_U29 (.ZN( u1_u9_u6_n114 ) , .A1( u1_u9_u6_n118 ) , .A2( u1_u9_u6_n126 ) , .B2( u1_u9_u6_n151 ) , .C2( u1_u9_u6_n159 ) , .C1( u1_u9_u6_n168 ) , .B1( u1_u9_u6_n169 ) );
  INV_X1 u1_u9_u6_U3 (.A( u1_u9_u6_n110 ) , .ZN( u1_u9_u6_n166 ) );
  NOR2_X1 u1_u9_u6_U30 (.A1( u1_u9_u6_n162 ) , .A2( u1_u9_u6_n165 ) , .ZN( u1_u9_u6_n98 ) );
  NAND2_X1 u1_u9_u6_U31 (.A1( u1_u9_u6_n144 ) , .ZN( u1_u9_u6_n151 ) , .A2( u1_u9_u6_n158 ) );
  NAND2_X1 u1_u9_u6_U32 (.ZN( u1_u9_u6_n132 ) , .A1( u1_u9_u6_n91 ) , .A2( u1_u9_u6_n97 ) );
  AOI22_X1 u1_u9_u6_U33 (.B2( u1_u9_u6_n110 ) , .B1( u1_u9_u6_n111 ) , .A1( u1_u9_u6_n112 ) , .ZN( u1_u9_u6_n115 ) , .A2( u1_u9_u6_n161 ) );
  NAND4_X1 u1_u9_u6_U34 (.A3( u1_u9_u6_n109 ) , .ZN( u1_u9_u6_n112 ) , .A4( u1_u9_u6_n132 ) , .A2( u1_u9_u6_n147 ) , .A1( u1_u9_u6_n166 ) );
  NOR2_X1 u1_u9_u6_U35 (.ZN( u1_u9_u6_n109 ) , .A1( u1_u9_u6_n170 ) , .A2( u1_u9_u6_n173 ) );
  NOR2_X1 u1_u9_u6_U36 (.A2( u1_u9_u6_n126 ) , .ZN( u1_u9_u6_n155 ) , .A1( u1_u9_u6_n160 ) );
  NAND2_X1 u1_u9_u6_U37 (.ZN( u1_u9_u6_n146 ) , .A2( u1_u9_u6_n94 ) , .A1( u1_u9_u6_n99 ) );
  AOI21_X1 u1_u9_u6_U38 (.A( u1_u9_u6_n144 ) , .B2( u1_u9_u6_n145 ) , .B1( u1_u9_u6_n146 ) , .ZN( u1_u9_u6_n150 ) );
  AOI211_X1 u1_u9_u6_U39 (.B( u1_u9_u6_n134 ) , .A( u1_u9_u6_n135 ) , .C1( u1_u9_u6_n136 ) , .ZN( u1_u9_u6_n137 ) , .C2( u1_u9_u6_n151 ) );
  INV_X1 u1_u9_u6_U4 (.A( u1_u9_u6_n142 ) , .ZN( u1_u9_u6_n174 ) );
  NAND4_X1 u1_u9_u6_U40 (.A4( u1_u9_u6_n127 ) , .A3( u1_u9_u6_n128 ) , .A2( u1_u9_u6_n129 ) , .A1( u1_u9_u6_n130 ) , .ZN( u1_u9_u6_n136 ) );
  AOI21_X1 u1_u9_u6_U41 (.B2( u1_u9_u6_n132 ) , .B1( u1_u9_u6_n133 ) , .ZN( u1_u9_u6_n134 ) , .A( u1_u9_u6_n158 ) );
  AOI21_X1 u1_u9_u6_U42 (.B1( u1_u9_u6_n131 ) , .ZN( u1_u9_u6_n135 ) , .A( u1_u9_u6_n144 ) , .B2( u1_u9_u6_n146 ) );
  INV_X1 u1_u9_u6_U43 (.A( u1_u9_u6_n111 ) , .ZN( u1_u9_u6_n158 ) );
  NAND2_X1 u1_u9_u6_U44 (.ZN( u1_u9_u6_n127 ) , .A1( u1_u9_u6_n91 ) , .A2( u1_u9_u6_n92 ) );
  NAND2_X1 u1_u9_u6_U45 (.ZN( u1_u9_u6_n129 ) , .A2( u1_u9_u6_n95 ) , .A1( u1_u9_u6_n96 ) );
  INV_X1 u1_u9_u6_U46 (.A( u1_u9_u6_n144 ) , .ZN( u1_u9_u6_n159 ) );
  NAND2_X1 u1_u9_u6_U47 (.ZN( u1_u9_u6_n145 ) , .A2( u1_u9_u6_n97 ) , .A1( u1_u9_u6_n98 ) );
  NAND2_X1 u1_u9_u6_U48 (.ZN( u1_u9_u6_n148 ) , .A2( u1_u9_u6_n92 ) , .A1( u1_u9_u6_n94 ) );
  NAND2_X1 u1_u9_u6_U49 (.ZN( u1_u9_u6_n108 ) , .A2( u1_u9_u6_n139 ) , .A1( u1_u9_u6_n144 ) );
  NAND2_X1 u1_u9_u6_U5 (.A2( u1_u9_u6_n143 ) , .ZN( u1_u9_u6_n152 ) , .A1( u1_u9_u6_n166 ) );
  NAND2_X1 u1_u9_u6_U50 (.ZN( u1_u9_u6_n121 ) , .A2( u1_u9_u6_n95 ) , .A1( u1_u9_u6_n97 ) );
  NAND2_X1 u1_u9_u6_U51 (.ZN( u1_u9_u6_n107 ) , .A2( u1_u9_u6_n92 ) , .A1( u1_u9_u6_n95 ) );
  AND2_X1 u1_u9_u6_U52 (.ZN( u1_u9_u6_n118 ) , .A2( u1_u9_u6_n91 ) , .A1( u1_u9_u6_n99 ) );
  NAND2_X1 u1_u9_u6_U53 (.ZN( u1_u9_u6_n147 ) , .A2( u1_u9_u6_n98 ) , .A1( u1_u9_u6_n99 ) );
  NAND2_X1 u1_u9_u6_U54 (.ZN( u1_u9_u6_n128 ) , .A1( u1_u9_u6_n94 ) , .A2( u1_u9_u6_n96 ) );
  NAND2_X1 u1_u9_u6_U55 (.ZN( u1_u9_u6_n119 ) , .A2( u1_u9_u6_n95 ) , .A1( u1_u9_u6_n99 ) );
  NAND2_X1 u1_u9_u6_U56 (.ZN( u1_u9_u6_n123 ) , .A2( u1_u9_u6_n91 ) , .A1( u1_u9_u6_n96 ) );
  NAND2_X1 u1_u9_u6_U57 (.ZN( u1_u9_u6_n100 ) , .A2( u1_u9_u6_n92 ) , .A1( u1_u9_u6_n98 ) );
  NAND2_X1 u1_u9_u6_U58 (.ZN( u1_u9_u6_n122 ) , .A1( u1_u9_u6_n94 ) , .A2( u1_u9_u6_n97 ) );
  INV_X1 u1_u9_u6_U59 (.A( u1_u9_u6_n139 ) , .ZN( u1_u9_u6_n160 ) );
  AOI22_X1 u1_u9_u6_U6 (.B2( u1_u9_u6_n101 ) , .A1( u1_u9_u6_n102 ) , .ZN( u1_u9_u6_n103 ) , .B1( u1_u9_u6_n160 ) , .A2( u1_u9_u6_n161 ) );
  NAND2_X1 u1_u9_u6_U60 (.ZN( u1_u9_u6_n113 ) , .A1( u1_u9_u6_n96 ) , .A2( u1_u9_u6_n98 ) );
  NOR2_X1 u1_u9_u6_U61 (.A2( u1_u9_X_40 ) , .A1( u1_u9_X_41 ) , .ZN( u1_u9_u6_n126 ) );
  NOR2_X1 u1_u9_u6_U62 (.A2( u1_u9_X_39 ) , .A1( u1_u9_X_42 ) , .ZN( u1_u9_u6_n92 ) );
  NOR2_X1 u1_u9_u6_U63 (.A2( u1_u9_X_39 ) , .A1( u1_u9_u6_n156 ) , .ZN( u1_u9_u6_n97 ) );
  NOR2_X1 u1_u9_u6_U64 (.A2( u1_u9_X_38 ) , .A1( u1_u9_u6_n165 ) , .ZN( u1_u9_u6_n95 ) );
  NOR2_X1 u1_u9_u6_U65 (.A2( u1_u9_X_41 ) , .ZN( u1_u9_u6_n111 ) , .A1( u1_u9_u6_n157 ) );
  NOR2_X1 u1_u9_u6_U66 (.A2( u1_u9_X_37 ) , .A1( u1_u9_u6_n162 ) , .ZN( u1_u9_u6_n94 ) );
  NOR2_X1 u1_u9_u6_U67 (.A2( u1_u9_X_37 ) , .A1( u1_u9_X_38 ) , .ZN( u1_u9_u6_n91 ) );
  NAND2_X1 u1_u9_u6_U68 (.A1( u1_u9_X_41 ) , .ZN( u1_u9_u6_n144 ) , .A2( u1_u9_u6_n157 ) );
  NAND2_X1 u1_u9_u6_U69 (.A2( u1_u9_X_40 ) , .A1( u1_u9_X_41 ) , .ZN( u1_u9_u6_n139 ) );
  NOR2_X1 u1_u9_u6_U7 (.A1( u1_u9_u6_n118 ) , .ZN( u1_u9_u6_n143 ) , .A2( u1_u9_u6_n168 ) );
  AND2_X1 u1_u9_u6_U70 (.A1( u1_u9_X_39 ) , .A2( u1_u9_u6_n156 ) , .ZN( u1_u9_u6_n96 ) );
  AND2_X1 u1_u9_u6_U71 (.A1( u1_u9_X_39 ) , .A2( u1_u9_X_42 ) , .ZN( u1_u9_u6_n99 ) );
  INV_X1 u1_u9_u6_U72 (.A( u1_u9_X_40 ) , .ZN( u1_u9_u6_n157 ) );
  INV_X1 u1_u9_u6_U73 (.A( u1_u9_X_37 ) , .ZN( u1_u9_u6_n165 ) );
  INV_X1 u1_u9_u6_U74 (.A( u1_u9_X_38 ) , .ZN( u1_u9_u6_n162 ) );
  INV_X1 u1_u9_u6_U75 (.A( u1_u9_X_42 ) , .ZN( u1_u9_u6_n156 ) );
  NAND4_X1 u1_u9_u6_U76 (.ZN( u1_out9_12 ) , .A4( u1_u9_u6_n114 ) , .A3( u1_u9_u6_n115 ) , .A2( u1_u9_u6_n116 ) , .A1( u1_u9_u6_n117 ) );
  OAI22_X1 u1_u9_u6_U77 (.B2( u1_u9_u6_n111 ) , .ZN( u1_u9_u6_n116 ) , .B1( u1_u9_u6_n126 ) , .A2( u1_u9_u6_n164 ) , .A1( u1_u9_u6_n167 ) );
  OAI21_X1 u1_u9_u6_U78 (.A( u1_u9_u6_n108 ) , .ZN( u1_u9_u6_n117 ) , .B2( u1_u9_u6_n141 ) , .B1( u1_u9_u6_n163 ) );
  NAND4_X1 u1_u9_u6_U79 (.ZN( u1_out9_32 ) , .A4( u1_u9_u6_n103 ) , .A3( u1_u9_u6_n104 ) , .A2( u1_u9_u6_n105 ) , .A1( u1_u9_u6_n106 ) );
  OAI21_X1 u1_u9_u6_U8 (.A( u1_u9_u6_n159 ) , .B1( u1_u9_u6_n169 ) , .B2( u1_u9_u6_n173 ) , .ZN( u1_u9_u6_n90 ) );
  AOI22_X1 u1_u9_u6_U80 (.ZN( u1_u9_u6_n105 ) , .A2( u1_u9_u6_n108 ) , .A1( u1_u9_u6_n118 ) , .B2( u1_u9_u6_n126 ) , .B1( u1_u9_u6_n171 ) );
  AOI22_X1 u1_u9_u6_U81 (.ZN( u1_u9_u6_n104 ) , .A1( u1_u9_u6_n111 ) , .B1( u1_u9_u6_n124 ) , .B2( u1_u9_u6_n151 ) , .A2( u1_u9_u6_n93 ) );
  OAI211_X1 u1_u9_u6_U82 (.ZN( u1_out9_7 ) , .B( u1_u9_u6_n153 ) , .C2( u1_u9_u6_n154 ) , .C1( u1_u9_u6_n155 ) , .A( u1_u9_u6_n174 ) );
  NOR3_X1 u1_u9_u6_U83 (.A1( u1_u9_u6_n141 ) , .ZN( u1_u9_u6_n154 ) , .A3( u1_u9_u6_n164 ) , .A2( u1_u9_u6_n171 ) );
  AOI211_X1 u1_u9_u6_U84 (.B( u1_u9_u6_n149 ) , .A( u1_u9_u6_n150 ) , .C2( u1_u9_u6_n151 ) , .C1( u1_u9_u6_n152 ) , .ZN( u1_u9_u6_n153 ) );
  OAI211_X1 u1_u9_u6_U85 (.ZN( u1_out9_22 ) , .B( u1_u9_u6_n137 ) , .A( u1_u9_u6_n138 ) , .C2( u1_u9_u6_n139 ) , .C1( u1_u9_u6_n140 ) );
  AOI22_X1 u1_u9_u6_U86 (.B1( u1_u9_u6_n124 ) , .A2( u1_u9_u6_n125 ) , .A1( u1_u9_u6_n126 ) , .ZN( u1_u9_u6_n138 ) , .B2( u1_u9_u6_n161 ) );
  AND4_X1 u1_u9_u6_U87 (.A3( u1_u9_u6_n119 ) , .A1( u1_u9_u6_n120 ) , .A4( u1_u9_u6_n129 ) , .ZN( u1_u9_u6_n140 ) , .A2( u1_u9_u6_n143 ) );
  NAND3_X1 u1_u9_u6_U88 (.A2( u1_u9_u6_n123 ) , .ZN( u1_u9_u6_n125 ) , .A1( u1_u9_u6_n130 ) , .A3( u1_u9_u6_n131 ) );
  NAND3_X1 u1_u9_u6_U89 (.A3( u1_u9_u6_n133 ) , .ZN( u1_u9_u6_n141 ) , .A1( u1_u9_u6_n145 ) , .A2( u1_u9_u6_n148 ) );
  INV_X1 u1_u9_u6_U9 (.ZN( u1_u9_u6_n172 ) , .A( u1_u9_u6_n88 ) );
  NAND3_X1 u1_u9_u6_U90 (.ZN( u1_u9_u6_n101 ) , .A3( u1_u9_u6_n107 ) , .A2( u1_u9_u6_n121 ) , .A1( u1_u9_u6_n127 ) );
  NAND3_X1 u1_u9_u6_U91 (.ZN( u1_u9_u6_n102 ) , .A3( u1_u9_u6_n130 ) , .A2( u1_u9_u6_n145 ) , .A1( u1_u9_u6_n166 ) );
  NAND3_X1 u1_u9_u6_U92 (.A3( u1_u9_u6_n113 ) , .A1( u1_u9_u6_n119 ) , .A2( u1_u9_u6_n123 ) , .ZN( u1_u9_u6_n93 ) );
  NAND3_X1 u1_u9_u6_U93 (.ZN( u1_u9_u6_n142 ) , .A2( u1_u9_u6_n172 ) , .A3( u1_u9_u6_n89 ) , .A1( u1_u9_u6_n90 ) );
  INV_X1 u1_uk_U1121 (.ZN( u1_K2_10 ) , .A( u1_uk_n1021 ) );
  INV_X1 u1_uk_U1157 (.ZN( u1_K10_12 ) , .A( u1_uk_n299 ) );
  INV_X1 u1_uk_U231 (.ZN( u1_K10_39 ) , .A( u1_uk_n373 ) );
  INV_X1 u1_uk_U369 (.ZN( u1_K7_46 ) , .A( u1_uk_n1124 ) );
  INV_X1 u1_uk_U371 (.ZN( u1_K10_40 ) , .A( u1_uk_n375 ) );
  INV_X1 u1_uk_U441 (.ZN( u1_K10_37 ) , .A( u1_uk_n366 ) );
  INV_X1 u1_uk_U445 (.ZN( u1_K10_9 ) , .A( u1_uk_n376 ) );
  INV_X1 u1_uk_U463 (.ZN( u1_K10_33 ) , .A( u1_uk_n349 ) );
  INV_X1 u1_uk_U465 (.ZN( u1_K1_33 ) , .A( u1_uk_n1011 ) );
  INV_X1 u1_uk_U574 (.ZN( u1_K10_38 ) , .A( u1_uk_n369 ) );
  INV_X1 u1_uk_U592 (.ZN( u1_K4_10 ) , .A( u1_uk_n1050 ) );
  INV_X1 u1_uk_U603 (.ZN( u1_K10_22 ) , .A( u1_uk_n312 ) );
  INV_X1 u1_uk_U622 (.ZN( u1_K10_35 ) , .A( u1_uk_n353 ) );
  INV_X1 u1_uk_U67 (.ZN( u1_K16_34 ) , .A( u1_uk_n988 ) );
  INV_X1 u1_uk_U798 (.ZN( u1_K1_27 ) , .A( u1_uk_n1007 ) );
  XOR2_X1 u2_U147 (.B( u2_L0_9 ) , .Z( u2_N40 ) , .A( u2_out1_9 ) );
  XOR2_X1 u2_U192 (.B( u2_L0_5 ) , .Z( u2_N36 ) , .A( u2_out1_5 ) );
  XOR2_X1 u2_U43 (.B( u2_L0_31 ) , .Z( u2_N62 ) , .A( u2_out1_31 ) );
  XOR2_X1 u2_U48 (.B( u2_L0_27 ) , .Z( u2_N58 ) , .A( u2_out1_27 ) );
  XOR2_X1 u2_U52 (.B( u2_L0_23 ) , .Z( u2_N54 ) , .A( u2_out1_23 ) );
  XOR2_X1 u2_U54 (.B( u2_L0_21 ) , .Z( u2_N52 ) , .A( u2_out1_21 ) );
  XOR2_X1 u2_U59 (.B( u2_L0_17 ) , .Z( u2_N48 ) , .A( u2_out1_17 ) );
  XOR2_X1 u2_U81 (.B( u2_L0_15 ) , .Z( u2_N46 ) , .A( u2_out1_15 ) );
  XOR2_X1 u2_u1_U10 (.B( u2_K2_45 ) , .A( u2_R0_30 ) , .Z( u2_u1_X_45 ) );
  XOR2_X1 u2_u1_U11 (.B( u2_K2_44 ) , .A( u2_R0_29 ) , .Z( u2_u1_X_44 ) );
  XOR2_X1 u2_u1_U12 (.B( u2_K2_43 ) , .A( u2_R0_28 ) , .Z( u2_u1_X_43 ) );
  XOR2_X1 u2_u1_U16 (.B( u2_K2_3 ) , .A( u2_R0_2 ) , .Z( u2_u1_X_3 ) );
  XOR2_X1 u2_u1_U27 (.B( u2_K2_2 ) , .A( u2_R0_1 ) , .Z( u2_u1_X_2 ) );
  XOR2_X1 u2_u1_U38 (.B( u2_K2_1 ) , .A( u2_R0_32 ) , .Z( u2_u1_X_1 ) );
  XOR2_X1 u2_u1_U4 (.B( u2_K2_6 ) , .A( u2_R0_5 ) , .Z( u2_u1_X_6 ) );
  XOR2_X1 u2_u1_U5 (.B( u2_K2_5 ) , .A( u2_R0_4 ) , .Z( u2_u1_X_5 ) );
  XOR2_X1 u2_u1_U6 (.B( u2_K2_4 ) , .A( u2_R0_3 ) , .Z( u2_u1_X_4 ) );
  XOR2_X1 u2_u1_U7 (.B( u2_K2_48 ) , .A( u2_R0_1 ) , .Z( u2_u1_X_48 ) );
  XOR2_X1 u2_u1_U8 (.B( u2_K2_47 ) , .A( u2_R0_32 ) , .Z( u2_u1_X_47 ) );
  XOR2_X1 u2_u1_U9 (.B( u2_K2_46 ) , .A( u2_R0_31 ) , .Z( u2_u1_X_46 ) );
  AND3_X1 u2_u1_u0_U10 (.A2( u2_u1_u0_n112 ) , .ZN( u2_u1_u0_n127 ) , .A3( u2_u1_u0_n130 ) , .A1( u2_u1_u0_n148 ) );
  NAND2_X1 u2_u1_u0_U11 (.ZN( u2_u1_u0_n113 ) , .A1( u2_u1_u0_n139 ) , .A2( u2_u1_u0_n149 ) );
  AND2_X1 u2_u1_u0_U12 (.ZN( u2_u1_u0_n107 ) , .A1( u2_u1_u0_n130 ) , .A2( u2_u1_u0_n140 ) );
  AND2_X1 u2_u1_u0_U13 (.A2( u2_u1_u0_n129 ) , .A1( u2_u1_u0_n130 ) , .ZN( u2_u1_u0_n151 ) );
  AND2_X1 u2_u1_u0_U14 (.A1( u2_u1_u0_n108 ) , .A2( u2_u1_u0_n125 ) , .ZN( u2_u1_u0_n145 ) );
  INV_X1 u2_u1_u0_U15 (.A( u2_u1_u0_n143 ) , .ZN( u2_u1_u0_n173 ) );
  NOR2_X1 u2_u1_u0_U16 (.A2( u2_u1_u0_n136 ) , .ZN( u2_u1_u0_n147 ) , .A1( u2_u1_u0_n160 ) );
  NOR2_X1 u2_u1_u0_U17 (.A1( u2_u1_u0_n163 ) , .A2( u2_u1_u0_n164 ) , .ZN( u2_u1_u0_n95 ) );
  AOI21_X1 u2_u1_u0_U18 (.B1( u2_u1_u0_n103 ) , .ZN( u2_u1_u0_n132 ) , .A( u2_u1_u0_n165 ) , .B2( u2_u1_u0_n93 ) );
  INV_X1 u2_u1_u0_U19 (.A( u2_u1_u0_n142 ) , .ZN( u2_u1_u0_n165 ) );
  OAI221_X1 u2_u1_u0_U20 (.C1( u2_u1_u0_n121 ) , .ZN( u2_u1_u0_n122 ) , .B2( u2_u1_u0_n127 ) , .A( u2_u1_u0_n143 ) , .B1( u2_u1_u0_n144 ) , .C2( u2_u1_u0_n147 ) );
  OAI22_X1 u2_u1_u0_U21 (.B1( u2_u1_u0_n125 ) , .ZN( u2_u1_u0_n126 ) , .A1( u2_u1_u0_n138 ) , .A2( u2_u1_u0_n146 ) , .B2( u2_u1_u0_n147 ) );
  OAI22_X1 u2_u1_u0_U22 (.B1( u2_u1_u0_n131 ) , .A1( u2_u1_u0_n144 ) , .B2( u2_u1_u0_n147 ) , .A2( u2_u1_u0_n90 ) , .ZN( u2_u1_u0_n91 ) );
  AND3_X1 u2_u1_u0_U23 (.A3( u2_u1_u0_n121 ) , .A2( u2_u1_u0_n125 ) , .A1( u2_u1_u0_n148 ) , .ZN( u2_u1_u0_n90 ) );
  NAND2_X1 u2_u1_u0_U24 (.A1( u2_u1_u0_n100 ) , .A2( u2_u1_u0_n103 ) , .ZN( u2_u1_u0_n125 ) );
  INV_X1 u2_u1_u0_U25 (.A( u2_u1_u0_n136 ) , .ZN( u2_u1_u0_n161 ) );
  NOR2_X1 u2_u1_u0_U26 (.A1( u2_u1_u0_n120 ) , .ZN( u2_u1_u0_n143 ) , .A2( u2_u1_u0_n167 ) );
  OAI221_X1 u2_u1_u0_U27 (.C1( u2_u1_u0_n112 ) , .ZN( u2_u1_u0_n120 ) , .B1( u2_u1_u0_n138 ) , .B2( u2_u1_u0_n141 ) , .C2( u2_u1_u0_n147 ) , .A( u2_u1_u0_n172 ) );
  AOI211_X1 u2_u1_u0_U28 (.B( u2_u1_u0_n115 ) , .A( u2_u1_u0_n116 ) , .C2( u2_u1_u0_n117 ) , .C1( u2_u1_u0_n118 ) , .ZN( u2_u1_u0_n119 ) );
  AOI22_X1 u2_u1_u0_U29 (.B2( u2_u1_u0_n109 ) , .A2( u2_u1_u0_n110 ) , .ZN( u2_u1_u0_n111 ) , .B1( u2_u1_u0_n118 ) , .A1( u2_u1_u0_n160 ) );
  INV_X1 u2_u1_u0_U3 (.A( u2_u1_u0_n113 ) , .ZN( u2_u1_u0_n166 ) );
  NAND2_X1 u2_u1_u0_U30 (.A1( u2_u1_u0_n100 ) , .ZN( u2_u1_u0_n129 ) , .A2( u2_u1_u0_n95 ) );
  INV_X1 u2_u1_u0_U31 (.A( u2_u1_u0_n118 ) , .ZN( u2_u1_u0_n158 ) );
  AOI21_X1 u2_u1_u0_U32 (.ZN( u2_u1_u0_n104 ) , .B1( u2_u1_u0_n107 ) , .B2( u2_u1_u0_n141 ) , .A( u2_u1_u0_n144 ) );
  AOI21_X1 u2_u1_u0_U33 (.B1( u2_u1_u0_n127 ) , .B2( u2_u1_u0_n129 ) , .A( u2_u1_u0_n138 ) , .ZN( u2_u1_u0_n96 ) );
  AOI21_X1 u2_u1_u0_U34 (.ZN( u2_u1_u0_n116 ) , .B2( u2_u1_u0_n142 ) , .A( u2_u1_u0_n144 ) , .B1( u2_u1_u0_n166 ) );
  NAND2_X1 u2_u1_u0_U35 (.A2( u2_u1_u0_n100 ) , .A1( u2_u1_u0_n101 ) , .ZN( u2_u1_u0_n139 ) );
  NAND2_X1 u2_u1_u0_U36 (.A2( u2_u1_u0_n100 ) , .ZN( u2_u1_u0_n131 ) , .A1( u2_u1_u0_n92 ) );
  NAND2_X1 u2_u1_u0_U37 (.A1( u2_u1_u0_n101 ) , .A2( u2_u1_u0_n102 ) , .ZN( u2_u1_u0_n150 ) );
  INV_X1 u2_u1_u0_U38 (.A( u2_u1_u0_n138 ) , .ZN( u2_u1_u0_n160 ) );
  NAND2_X1 u2_u1_u0_U39 (.A1( u2_u1_u0_n102 ) , .ZN( u2_u1_u0_n128 ) , .A2( u2_u1_u0_n95 ) );
  AOI21_X1 u2_u1_u0_U4 (.B1( u2_u1_u0_n114 ) , .ZN( u2_u1_u0_n115 ) , .B2( u2_u1_u0_n129 ) , .A( u2_u1_u0_n161 ) );
  NAND2_X1 u2_u1_u0_U40 (.ZN( u2_u1_u0_n148 ) , .A1( u2_u1_u0_n93 ) , .A2( u2_u1_u0_n95 ) );
  NAND2_X1 u2_u1_u0_U41 (.A2( u2_u1_u0_n102 ) , .A1( u2_u1_u0_n103 ) , .ZN( u2_u1_u0_n149 ) );
  NAND2_X1 u2_u1_u0_U42 (.A2( u2_u1_u0_n102 ) , .ZN( u2_u1_u0_n114 ) , .A1( u2_u1_u0_n92 ) );
  NAND2_X1 u2_u1_u0_U43 (.A2( u2_u1_u0_n101 ) , .ZN( u2_u1_u0_n121 ) , .A1( u2_u1_u0_n93 ) );
  INV_X1 u2_u1_u0_U44 (.ZN( u2_u1_u0_n172 ) , .A( u2_u1_u0_n88 ) );
  OAI222_X1 u2_u1_u0_U45 (.C1( u2_u1_u0_n108 ) , .A1( u2_u1_u0_n125 ) , .B2( u2_u1_u0_n128 ) , .B1( u2_u1_u0_n144 ) , .A2( u2_u1_u0_n158 ) , .C2( u2_u1_u0_n161 ) , .ZN( u2_u1_u0_n88 ) );
  NAND2_X1 u2_u1_u0_U46 (.ZN( u2_u1_u0_n112 ) , .A2( u2_u1_u0_n92 ) , .A1( u2_u1_u0_n93 ) );
  OR3_X1 u2_u1_u0_U47 (.A3( u2_u1_u0_n152 ) , .A2( u2_u1_u0_n153 ) , .A1( u2_u1_u0_n154 ) , .ZN( u2_u1_u0_n155 ) );
  AOI21_X1 u2_u1_u0_U48 (.B2( u2_u1_u0_n150 ) , .B1( u2_u1_u0_n151 ) , .ZN( u2_u1_u0_n152 ) , .A( u2_u1_u0_n158 ) );
  AOI21_X1 u2_u1_u0_U49 (.A( u2_u1_u0_n144 ) , .B2( u2_u1_u0_n145 ) , .B1( u2_u1_u0_n146 ) , .ZN( u2_u1_u0_n154 ) );
  AOI21_X1 u2_u1_u0_U5 (.B2( u2_u1_u0_n131 ) , .ZN( u2_u1_u0_n134 ) , .B1( u2_u1_u0_n151 ) , .A( u2_u1_u0_n158 ) );
  AOI21_X1 u2_u1_u0_U50 (.A( u2_u1_u0_n147 ) , .B2( u2_u1_u0_n148 ) , .B1( u2_u1_u0_n149 ) , .ZN( u2_u1_u0_n153 ) );
  INV_X1 u2_u1_u0_U51 (.ZN( u2_u1_u0_n171 ) , .A( u2_u1_u0_n99 ) );
  OAI211_X1 u2_u1_u0_U52 (.C2( u2_u1_u0_n140 ) , .C1( u2_u1_u0_n161 ) , .A( u2_u1_u0_n169 ) , .B( u2_u1_u0_n98 ) , .ZN( u2_u1_u0_n99 ) );
  AOI211_X1 u2_u1_u0_U53 (.C1( u2_u1_u0_n118 ) , .A( u2_u1_u0_n123 ) , .B( u2_u1_u0_n96 ) , .C2( u2_u1_u0_n97 ) , .ZN( u2_u1_u0_n98 ) );
  INV_X1 u2_u1_u0_U54 (.ZN( u2_u1_u0_n169 ) , .A( u2_u1_u0_n91 ) );
  NOR2_X1 u2_u1_u0_U55 (.A2( u2_u1_X_4 ) , .A1( u2_u1_X_5 ) , .ZN( u2_u1_u0_n118 ) );
  NOR2_X1 u2_u1_u0_U56 (.A2( u2_u1_X_2 ) , .ZN( u2_u1_u0_n103 ) , .A1( u2_u1_u0_n164 ) );
  NOR2_X1 u2_u1_u0_U57 (.A2( u2_u1_X_1 ) , .A1( u2_u1_X_2 ) , .ZN( u2_u1_u0_n92 ) );
  NOR2_X1 u2_u1_u0_U58 (.A2( u2_u1_X_1 ) , .ZN( u2_u1_u0_n101 ) , .A1( u2_u1_u0_n163 ) );
  NAND2_X1 u2_u1_u0_U59 (.A2( u2_u1_X_4 ) , .A1( u2_u1_X_5 ) , .ZN( u2_u1_u0_n144 ) );
  NOR2_X1 u2_u1_u0_U6 (.A1( u2_u1_u0_n108 ) , .ZN( u2_u1_u0_n123 ) , .A2( u2_u1_u0_n158 ) );
  NOR2_X1 u2_u1_u0_U60 (.A2( u2_u1_X_5 ) , .ZN( u2_u1_u0_n136 ) , .A1( u2_u1_u0_n159 ) );
  NAND2_X1 u2_u1_u0_U61 (.A1( u2_u1_X_5 ) , .ZN( u2_u1_u0_n138 ) , .A2( u2_u1_u0_n159 ) );
  AND2_X1 u2_u1_u0_U62 (.A2( u2_u1_X_3 ) , .A1( u2_u1_X_6 ) , .ZN( u2_u1_u0_n102 ) );
  AND2_X1 u2_u1_u0_U63 (.A1( u2_u1_X_6 ) , .A2( u2_u1_u0_n162 ) , .ZN( u2_u1_u0_n93 ) );
  INV_X1 u2_u1_u0_U64 (.A( u2_u1_X_4 ) , .ZN( u2_u1_u0_n159 ) );
  INV_X1 u2_u1_u0_U65 (.A( u2_u1_X_1 ) , .ZN( u2_u1_u0_n164 ) );
  INV_X1 u2_u1_u0_U66 (.A( u2_u1_X_2 ) , .ZN( u2_u1_u0_n163 ) );
  INV_X1 u2_u1_u0_U67 (.A( u2_u1_X_3 ) , .ZN( u2_u1_u0_n162 ) );
  INV_X1 u2_u1_u0_U68 (.A( u2_u1_u0_n126 ) , .ZN( u2_u1_u0_n168 ) );
  AOI211_X1 u2_u1_u0_U69 (.B( u2_u1_u0_n133 ) , .A( u2_u1_u0_n134 ) , .C2( u2_u1_u0_n135 ) , .C1( u2_u1_u0_n136 ) , .ZN( u2_u1_u0_n137 ) );
  OAI21_X1 u2_u1_u0_U7 (.B1( u2_u1_u0_n150 ) , .B2( u2_u1_u0_n158 ) , .A( u2_u1_u0_n172 ) , .ZN( u2_u1_u0_n89 ) );
  INV_X1 u2_u1_u0_U70 (.ZN( u2_u1_u0_n174 ) , .A( u2_u1_u0_n89 ) );
  AOI211_X1 u2_u1_u0_U71 (.B( u2_u1_u0_n104 ) , .A( u2_u1_u0_n105 ) , .ZN( u2_u1_u0_n106 ) , .C2( u2_u1_u0_n113 ) , .C1( u2_u1_u0_n160 ) );
  OR4_X1 u2_u1_u0_U72 (.ZN( u2_out1_17 ) , .A4( u2_u1_u0_n122 ) , .A2( u2_u1_u0_n123 ) , .A1( u2_u1_u0_n124 ) , .A3( u2_u1_u0_n170 ) );
  AOI21_X1 u2_u1_u0_U73 (.B2( u2_u1_u0_n107 ) , .ZN( u2_u1_u0_n124 ) , .B1( u2_u1_u0_n128 ) , .A( u2_u1_u0_n161 ) );
  INV_X1 u2_u1_u0_U74 (.A( u2_u1_u0_n111 ) , .ZN( u2_u1_u0_n170 ) );
  OR4_X1 u2_u1_u0_U75 (.ZN( u2_out1_31 ) , .A4( u2_u1_u0_n155 ) , .A2( u2_u1_u0_n156 ) , .A1( u2_u1_u0_n157 ) , .A3( u2_u1_u0_n173 ) );
  AOI21_X1 u2_u1_u0_U76 (.A( u2_u1_u0_n138 ) , .B2( u2_u1_u0_n139 ) , .B1( u2_u1_u0_n140 ) , .ZN( u2_u1_u0_n157 ) );
  AOI21_X1 u2_u1_u0_U77 (.B2( u2_u1_u0_n141 ) , .B1( u2_u1_u0_n142 ) , .ZN( u2_u1_u0_n156 ) , .A( u2_u1_u0_n161 ) );
  AOI21_X1 u2_u1_u0_U78 (.B1( u2_u1_u0_n132 ) , .ZN( u2_u1_u0_n133 ) , .A( u2_u1_u0_n144 ) , .B2( u2_u1_u0_n166 ) );
  OAI22_X1 u2_u1_u0_U79 (.ZN( u2_u1_u0_n105 ) , .A2( u2_u1_u0_n132 ) , .B1( u2_u1_u0_n146 ) , .A1( u2_u1_u0_n147 ) , .B2( u2_u1_u0_n161 ) );
  AND2_X1 u2_u1_u0_U8 (.A1( u2_u1_u0_n114 ) , .A2( u2_u1_u0_n121 ) , .ZN( u2_u1_u0_n146 ) );
  NAND2_X1 u2_u1_u0_U80 (.ZN( u2_u1_u0_n110 ) , .A2( u2_u1_u0_n132 ) , .A1( u2_u1_u0_n145 ) );
  INV_X1 u2_u1_u0_U81 (.A( u2_u1_u0_n119 ) , .ZN( u2_u1_u0_n167 ) );
  NAND2_X1 u2_u1_u0_U82 (.A2( u2_u1_u0_n103 ) , .ZN( u2_u1_u0_n140 ) , .A1( u2_u1_u0_n94 ) );
  NAND2_X1 u2_u1_u0_U83 (.A1( u2_u1_u0_n101 ) , .ZN( u2_u1_u0_n130 ) , .A2( u2_u1_u0_n94 ) );
  NAND2_X1 u2_u1_u0_U84 (.ZN( u2_u1_u0_n108 ) , .A1( u2_u1_u0_n92 ) , .A2( u2_u1_u0_n94 ) );
  NAND2_X1 u2_u1_u0_U85 (.ZN( u2_u1_u0_n142 ) , .A1( u2_u1_u0_n94 ) , .A2( u2_u1_u0_n95 ) );
  NOR2_X1 u2_u1_u0_U86 (.A2( u2_u1_X_6 ) , .ZN( u2_u1_u0_n100 ) , .A1( u2_u1_u0_n162 ) );
  NOR2_X1 u2_u1_u0_U87 (.A2( u2_u1_X_3 ) , .A1( u2_u1_X_6 ) , .ZN( u2_u1_u0_n94 ) );
  NAND3_X1 u2_u1_u0_U88 (.ZN( u2_out1_23 ) , .A3( u2_u1_u0_n137 ) , .A1( u2_u1_u0_n168 ) , .A2( u2_u1_u0_n171 ) );
  NAND3_X1 u2_u1_u0_U89 (.A3( u2_u1_u0_n127 ) , .A2( u2_u1_u0_n128 ) , .ZN( u2_u1_u0_n135 ) , .A1( u2_u1_u0_n150 ) );
  AND2_X1 u2_u1_u0_U9 (.A1( u2_u1_u0_n131 ) , .ZN( u2_u1_u0_n141 ) , .A2( u2_u1_u0_n150 ) );
  NAND3_X1 u2_u1_u0_U90 (.ZN( u2_u1_u0_n117 ) , .A3( u2_u1_u0_n132 ) , .A2( u2_u1_u0_n139 ) , .A1( u2_u1_u0_n148 ) );
  NAND3_X1 u2_u1_u0_U91 (.ZN( u2_u1_u0_n109 ) , .A2( u2_u1_u0_n114 ) , .A3( u2_u1_u0_n140 ) , .A1( u2_u1_u0_n149 ) );
  NAND3_X1 u2_u1_u0_U92 (.ZN( u2_out1_9 ) , .A3( u2_u1_u0_n106 ) , .A2( u2_u1_u0_n171 ) , .A1( u2_u1_u0_n174 ) );
  NAND3_X1 u2_u1_u0_U93 (.A2( u2_u1_u0_n128 ) , .A1( u2_u1_u0_n132 ) , .A3( u2_u1_u0_n146 ) , .ZN( u2_u1_u0_n97 ) );
  AND3_X1 u2_u1_u7_U10 (.A3( u2_u1_u7_n110 ) , .A2( u2_u1_u7_n127 ) , .A1( u2_u1_u7_n132 ) , .ZN( u2_u1_u7_n92 ) );
  OAI21_X1 u2_u1_u7_U11 (.A( u2_u1_u7_n161 ) , .B1( u2_u1_u7_n168 ) , .B2( u2_u1_u7_n173 ) , .ZN( u2_u1_u7_n91 ) );
  AOI211_X1 u2_u1_u7_U12 (.A( u2_u1_u7_n117 ) , .ZN( u2_u1_u7_n118 ) , .C2( u2_u1_u7_n126 ) , .C1( u2_u1_u7_n177 ) , .B( u2_u1_u7_n180 ) );
  OAI22_X1 u2_u1_u7_U13 (.B1( u2_u1_u7_n115 ) , .ZN( u2_u1_u7_n117 ) , .A2( u2_u1_u7_n133 ) , .A1( u2_u1_u7_n137 ) , .B2( u2_u1_u7_n162 ) );
  INV_X1 u2_u1_u7_U14 (.A( u2_u1_u7_n116 ) , .ZN( u2_u1_u7_n180 ) );
  NOR3_X1 u2_u1_u7_U15 (.ZN( u2_u1_u7_n115 ) , .A3( u2_u1_u7_n145 ) , .A2( u2_u1_u7_n168 ) , .A1( u2_u1_u7_n169 ) );
  OAI211_X1 u2_u1_u7_U16 (.B( u2_u1_u7_n122 ) , .A( u2_u1_u7_n123 ) , .C2( u2_u1_u7_n124 ) , .ZN( u2_u1_u7_n154 ) , .C1( u2_u1_u7_n162 ) );
  AOI222_X1 u2_u1_u7_U17 (.ZN( u2_u1_u7_n122 ) , .C2( u2_u1_u7_n126 ) , .C1( u2_u1_u7_n145 ) , .B1( u2_u1_u7_n161 ) , .A2( u2_u1_u7_n165 ) , .B2( u2_u1_u7_n170 ) , .A1( u2_u1_u7_n176 ) );
  INV_X1 u2_u1_u7_U18 (.A( u2_u1_u7_n133 ) , .ZN( u2_u1_u7_n176 ) );
  NOR3_X1 u2_u1_u7_U19 (.A2( u2_u1_u7_n134 ) , .A1( u2_u1_u7_n135 ) , .ZN( u2_u1_u7_n136 ) , .A3( u2_u1_u7_n171 ) );
  NOR2_X1 u2_u1_u7_U20 (.A1( u2_u1_u7_n130 ) , .A2( u2_u1_u7_n134 ) , .ZN( u2_u1_u7_n153 ) );
  INV_X1 u2_u1_u7_U21 (.A( u2_u1_u7_n101 ) , .ZN( u2_u1_u7_n165 ) );
  NOR2_X1 u2_u1_u7_U22 (.ZN( u2_u1_u7_n111 ) , .A2( u2_u1_u7_n134 ) , .A1( u2_u1_u7_n169 ) );
  AOI21_X1 u2_u1_u7_U23 (.ZN( u2_u1_u7_n104 ) , .B2( u2_u1_u7_n112 ) , .B1( u2_u1_u7_n127 ) , .A( u2_u1_u7_n164 ) );
  AOI21_X1 u2_u1_u7_U24 (.ZN( u2_u1_u7_n106 ) , .B1( u2_u1_u7_n133 ) , .B2( u2_u1_u7_n146 ) , .A( u2_u1_u7_n162 ) );
  AOI21_X1 u2_u1_u7_U25 (.A( u2_u1_u7_n101 ) , .ZN( u2_u1_u7_n107 ) , .B2( u2_u1_u7_n128 ) , .B1( u2_u1_u7_n175 ) );
  INV_X1 u2_u1_u7_U26 (.A( u2_u1_u7_n138 ) , .ZN( u2_u1_u7_n171 ) );
  INV_X1 u2_u1_u7_U27 (.A( u2_u1_u7_n131 ) , .ZN( u2_u1_u7_n177 ) );
  INV_X1 u2_u1_u7_U28 (.A( u2_u1_u7_n110 ) , .ZN( u2_u1_u7_n174 ) );
  NAND2_X1 u2_u1_u7_U29 (.A1( u2_u1_u7_n129 ) , .A2( u2_u1_u7_n132 ) , .ZN( u2_u1_u7_n149 ) );
  OAI21_X1 u2_u1_u7_U3 (.ZN( u2_u1_u7_n159 ) , .A( u2_u1_u7_n165 ) , .B2( u2_u1_u7_n171 ) , .B1( u2_u1_u7_n174 ) );
  NAND2_X1 u2_u1_u7_U30 (.A1( u2_u1_u7_n113 ) , .A2( u2_u1_u7_n124 ) , .ZN( u2_u1_u7_n130 ) );
  INV_X1 u2_u1_u7_U31 (.A( u2_u1_u7_n112 ) , .ZN( u2_u1_u7_n173 ) );
  INV_X1 u2_u1_u7_U32 (.A( u2_u1_u7_n128 ) , .ZN( u2_u1_u7_n168 ) );
  INV_X1 u2_u1_u7_U33 (.A( u2_u1_u7_n148 ) , .ZN( u2_u1_u7_n169 ) );
  INV_X1 u2_u1_u7_U34 (.A( u2_u1_u7_n127 ) , .ZN( u2_u1_u7_n179 ) );
  NOR2_X1 u2_u1_u7_U35 (.ZN( u2_u1_u7_n101 ) , .A2( u2_u1_u7_n150 ) , .A1( u2_u1_u7_n156 ) );
  AOI211_X1 u2_u1_u7_U36 (.B( u2_u1_u7_n154 ) , .A( u2_u1_u7_n155 ) , .C1( u2_u1_u7_n156 ) , .ZN( u2_u1_u7_n157 ) , .C2( u2_u1_u7_n172 ) );
  INV_X1 u2_u1_u7_U37 (.A( u2_u1_u7_n153 ) , .ZN( u2_u1_u7_n172 ) );
  AOI211_X1 u2_u1_u7_U38 (.B( u2_u1_u7_n139 ) , .A( u2_u1_u7_n140 ) , .C2( u2_u1_u7_n141 ) , .ZN( u2_u1_u7_n142 ) , .C1( u2_u1_u7_n156 ) );
  NAND4_X1 u2_u1_u7_U39 (.A3( u2_u1_u7_n127 ) , .A2( u2_u1_u7_n128 ) , .A1( u2_u1_u7_n129 ) , .ZN( u2_u1_u7_n141 ) , .A4( u2_u1_u7_n147 ) );
  INV_X1 u2_u1_u7_U4 (.A( u2_u1_u7_n111 ) , .ZN( u2_u1_u7_n170 ) );
  AOI21_X1 u2_u1_u7_U40 (.A( u2_u1_u7_n137 ) , .B1( u2_u1_u7_n138 ) , .ZN( u2_u1_u7_n139 ) , .B2( u2_u1_u7_n146 ) );
  OAI22_X1 u2_u1_u7_U41 (.B1( u2_u1_u7_n136 ) , .ZN( u2_u1_u7_n140 ) , .A1( u2_u1_u7_n153 ) , .B2( u2_u1_u7_n162 ) , .A2( u2_u1_u7_n164 ) );
  AOI21_X1 u2_u1_u7_U42 (.ZN( u2_u1_u7_n123 ) , .B1( u2_u1_u7_n165 ) , .B2( u2_u1_u7_n177 ) , .A( u2_u1_u7_n97 ) );
  AOI21_X1 u2_u1_u7_U43 (.B2( u2_u1_u7_n113 ) , .B1( u2_u1_u7_n124 ) , .A( u2_u1_u7_n125 ) , .ZN( u2_u1_u7_n97 ) );
  INV_X1 u2_u1_u7_U44 (.A( u2_u1_u7_n125 ) , .ZN( u2_u1_u7_n161 ) );
  INV_X1 u2_u1_u7_U45 (.A( u2_u1_u7_n152 ) , .ZN( u2_u1_u7_n162 ) );
  AOI22_X1 u2_u1_u7_U46 (.A2( u2_u1_u7_n114 ) , .ZN( u2_u1_u7_n119 ) , .B1( u2_u1_u7_n130 ) , .A1( u2_u1_u7_n156 ) , .B2( u2_u1_u7_n165 ) );
  NAND2_X1 u2_u1_u7_U47 (.A2( u2_u1_u7_n112 ) , .ZN( u2_u1_u7_n114 ) , .A1( u2_u1_u7_n175 ) );
  AND2_X1 u2_u1_u7_U48 (.ZN( u2_u1_u7_n145 ) , .A2( u2_u1_u7_n98 ) , .A1( u2_u1_u7_n99 ) );
  NOR2_X1 u2_u1_u7_U49 (.ZN( u2_u1_u7_n137 ) , .A1( u2_u1_u7_n150 ) , .A2( u2_u1_u7_n161 ) );
  INV_X1 u2_u1_u7_U5 (.A( u2_u1_u7_n149 ) , .ZN( u2_u1_u7_n175 ) );
  AOI21_X1 u2_u1_u7_U50 (.ZN( u2_u1_u7_n105 ) , .B2( u2_u1_u7_n110 ) , .A( u2_u1_u7_n125 ) , .B1( u2_u1_u7_n147 ) );
  NAND2_X1 u2_u1_u7_U51 (.ZN( u2_u1_u7_n146 ) , .A1( u2_u1_u7_n95 ) , .A2( u2_u1_u7_n98 ) );
  NAND2_X1 u2_u1_u7_U52 (.A2( u2_u1_u7_n103 ) , .ZN( u2_u1_u7_n147 ) , .A1( u2_u1_u7_n93 ) );
  NAND2_X1 u2_u1_u7_U53 (.A1( u2_u1_u7_n103 ) , .ZN( u2_u1_u7_n127 ) , .A2( u2_u1_u7_n99 ) );
  OR2_X1 u2_u1_u7_U54 (.ZN( u2_u1_u7_n126 ) , .A2( u2_u1_u7_n152 ) , .A1( u2_u1_u7_n156 ) );
  NAND2_X1 u2_u1_u7_U55 (.A2( u2_u1_u7_n102 ) , .A1( u2_u1_u7_n103 ) , .ZN( u2_u1_u7_n133 ) );
  NAND2_X1 u2_u1_u7_U56 (.ZN( u2_u1_u7_n112 ) , .A2( u2_u1_u7_n96 ) , .A1( u2_u1_u7_n99 ) );
  NAND2_X1 u2_u1_u7_U57 (.A2( u2_u1_u7_n102 ) , .ZN( u2_u1_u7_n128 ) , .A1( u2_u1_u7_n98 ) );
  NAND2_X1 u2_u1_u7_U58 (.A1( u2_u1_u7_n100 ) , .ZN( u2_u1_u7_n113 ) , .A2( u2_u1_u7_n93 ) );
  NAND2_X1 u2_u1_u7_U59 (.A2( u2_u1_u7_n102 ) , .ZN( u2_u1_u7_n124 ) , .A1( u2_u1_u7_n96 ) );
  INV_X1 u2_u1_u7_U6 (.A( u2_u1_u7_n154 ) , .ZN( u2_u1_u7_n178 ) );
  NAND2_X1 u2_u1_u7_U60 (.ZN( u2_u1_u7_n110 ) , .A1( u2_u1_u7_n95 ) , .A2( u2_u1_u7_n96 ) );
  INV_X1 u2_u1_u7_U61 (.A( u2_u1_u7_n150 ) , .ZN( u2_u1_u7_n164 ) );
  AND2_X1 u2_u1_u7_U62 (.ZN( u2_u1_u7_n134 ) , .A1( u2_u1_u7_n93 ) , .A2( u2_u1_u7_n98 ) );
  NAND2_X1 u2_u1_u7_U63 (.A1( u2_u1_u7_n100 ) , .A2( u2_u1_u7_n102 ) , .ZN( u2_u1_u7_n129 ) );
  NAND2_X1 u2_u1_u7_U64 (.A2( u2_u1_u7_n103 ) , .ZN( u2_u1_u7_n131 ) , .A1( u2_u1_u7_n95 ) );
  NAND2_X1 u2_u1_u7_U65 (.A1( u2_u1_u7_n100 ) , .ZN( u2_u1_u7_n138 ) , .A2( u2_u1_u7_n99 ) );
  NAND2_X1 u2_u1_u7_U66 (.ZN( u2_u1_u7_n132 ) , .A1( u2_u1_u7_n93 ) , .A2( u2_u1_u7_n96 ) );
  NAND2_X1 u2_u1_u7_U67 (.A1( u2_u1_u7_n100 ) , .ZN( u2_u1_u7_n148 ) , .A2( u2_u1_u7_n95 ) );
  NOR2_X1 u2_u1_u7_U68 (.A2( u2_u1_X_47 ) , .ZN( u2_u1_u7_n150 ) , .A1( u2_u1_u7_n163 ) );
  NOR2_X1 u2_u1_u7_U69 (.A2( u2_u1_X_43 ) , .A1( u2_u1_X_44 ) , .ZN( u2_u1_u7_n103 ) );
  AOI211_X1 u2_u1_u7_U7 (.ZN( u2_u1_u7_n116 ) , .A( u2_u1_u7_n155 ) , .C1( u2_u1_u7_n161 ) , .C2( u2_u1_u7_n171 ) , .B( u2_u1_u7_n94 ) );
  NOR2_X1 u2_u1_u7_U70 (.A2( u2_u1_X_48 ) , .A1( u2_u1_u7_n166 ) , .ZN( u2_u1_u7_n95 ) );
  NOR2_X1 u2_u1_u7_U71 (.A2( u2_u1_X_45 ) , .A1( u2_u1_X_48 ) , .ZN( u2_u1_u7_n99 ) );
  NOR2_X1 u2_u1_u7_U72 (.A2( u2_u1_X_44 ) , .A1( u2_u1_u7_n167 ) , .ZN( u2_u1_u7_n98 ) );
  NOR2_X1 u2_u1_u7_U73 (.A2( u2_u1_X_46 ) , .A1( u2_u1_X_47 ) , .ZN( u2_u1_u7_n152 ) );
  AND2_X1 u2_u1_u7_U74 (.A1( u2_u1_X_47 ) , .ZN( u2_u1_u7_n156 ) , .A2( u2_u1_u7_n163 ) );
  NAND2_X1 u2_u1_u7_U75 (.A2( u2_u1_X_46 ) , .A1( u2_u1_X_47 ) , .ZN( u2_u1_u7_n125 ) );
  AND2_X1 u2_u1_u7_U76 (.A2( u2_u1_X_45 ) , .A1( u2_u1_X_48 ) , .ZN( u2_u1_u7_n102 ) );
  AND2_X1 u2_u1_u7_U77 (.A2( u2_u1_X_43 ) , .A1( u2_u1_X_44 ) , .ZN( u2_u1_u7_n96 ) );
  AND2_X1 u2_u1_u7_U78 (.A1( u2_u1_X_44 ) , .ZN( u2_u1_u7_n100 ) , .A2( u2_u1_u7_n167 ) );
  AND2_X1 u2_u1_u7_U79 (.A1( u2_u1_X_48 ) , .A2( u2_u1_u7_n166 ) , .ZN( u2_u1_u7_n93 ) );
  OAI222_X1 u2_u1_u7_U8 (.C2( u2_u1_u7_n101 ) , .B2( u2_u1_u7_n111 ) , .A1( u2_u1_u7_n113 ) , .C1( u2_u1_u7_n146 ) , .A2( u2_u1_u7_n162 ) , .B1( u2_u1_u7_n164 ) , .ZN( u2_u1_u7_n94 ) );
  INV_X1 u2_u1_u7_U80 (.A( u2_u1_X_46 ) , .ZN( u2_u1_u7_n163 ) );
  INV_X1 u2_u1_u7_U81 (.A( u2_u1_X_43 ) , .ZN( u2_u1_u7_n167 ) );
  INV_X1 u2_u1_u7_U82 (.A( u2_u1_X_45 ) , .ZN( u2_u1_u7_n166 ) );
  NAND4_X1 u2_u1_u7_U83 (.ZN( u2_out1_27 ) , .A4( u2_u1_u7_n118 ) , .A3( u2_u1_u7_n119 ) , .A2( u2_u1_u7_n120 ) , .A1( u2_u1_u7_n121 ) );
  OAI21_X1 u2_u1_u7_U84 (.ZN( u2_u1_u7_n121 ) , .B2( u2_u1_u7_n145 ) , .A( u2_u1_u7_n150 ) , .B1( u2_u1_u7_n174 ) );
  OAI21_X1 u2_u1_u7_U85 (.ZN( u2_u1_u7_n120 ) , .A( u2_u1_u7_n161 ) , .B2( u2_u1_u7_n170 ) , .B1( u2_u1_u7_n179 ) );
  NAND4_X1 u2_u1_u7_U86 (.ZN( u2_out1_15 ) , .A4( u2_u1_u7_n142 ) , .A3( u2_u1_u7_n143 ) , .A2( u2_u1_u7_n144 ) , .A1( u2_u1_u7_n178 ) );
  OR2_X1 u2_u1_u7_U87 (.A2( u2_u1_u7_n125 ) , .A1( u2_u1_u7_n129 ) , .ZN( u2_u1_u7_n144 ) );
  AOI22_X1 u2_u1_u7_U88 (.A2( u2_u1_u7_n126 ) , .ZN( u2_u1_u7_n143 ) , .B2( u2_u1_u7_n165 ) , .B1( u2_u1_u7_n173 ) , .A1( u2_u1_u7_n174 ) );
  NAND4_X1 u2_u1_u7_U89 (.ZN( u2_out1_5 ) , .A4( u2_u1_u7_n108 ) , .A3( u2_u1_u7_n109 ) , .A1( u2_u1_u7_n116 ) , .A2( u2_u1_u7_n123 ) );
  OAI221_X1 u2_u1_u7_U9 (.C1( u2_u1_u7_n101 ) , .C2( u2_u1_u7_n147 ) , .ZN( u2_u1_u7_n155 ) , .B2( u2_u1_u7_n162 ) , .A( u2_u1_u7_n91 ) , .B1( u2_u1_u7_n92 ) );
  AOI22_X1 u2_u1_u7_U90 (.ZN( u2_u1_u7_n109 ) , .A2( u2_u1_u7_n126 ) , .B2( u2_u1_u7_n145 ) , .B1( u2_u1_u7_n156 ) , .A1( u2_u1_u7_n171 ) );
  NOR4_X1 u2_u1_u7_U91 (.A4( u2_u1_u7_n104 ) , .A3( u2_u1_u7_n105 ) , .A2( u2_u1_u7_n106 ) , .A1( u2_u1_u7_n107 ) , .ZN( u2_u1_u7_n108 ) );
  NAND4_X1 u2_u1_u7_U92 (.ZN( u2_out1_21 ) , .A4( u2_u1_u7_n157 ) , .A3( u2_u1_u7_n158 ) , .A2( u2_u1_u7_n159 ) , .A1( u2_u1_u7_n160 ) );
  OAI21_X1 u2_u1_u7_U93 (.B1( u2_u1_u7_n145 ) , .ZN( u2_u1_u7_n160 ) , .A( u2_u1_u7_n161 ) , .B2( u2_u1_u7_n177 ) );
  AOI22_X1 u2_u1_u7_U94 (.B2( u2_u1_u7_n149 ) , .B1( u2_u1_u7_n150 ) , .A2( u2_u1_u7_n151 ) , .A1( u2_u1_u7_n152 ) , .ZN( u2_u1_u7_n158 ) );
  NAND3_X1 u2_u1_u7_U95 (.A3( u2_u1_u7_n146 ) , .A2( u2_u1_u7_n147 ) , .A1( u2_u1_u7_n148 ) , .ZN( u2_u1_u7_n151 ) );
  NAND3_X1 u2_u1_u7_U96 (.A3( u2_u1_u7_n131 ) , .A2( u2_u1_u7_n132 ) , .A1( u2_u1_u7_n133 ) , .ZN( u2_u1_u7_n135 ) );
  OAI22_X1 u2_uk_U104 (.ZN( u2_K2_5 ) , .B1( u2_uk_n10 ) , .B2( u2_uk_n1244 ) , .A2( u2_uk_n1247 ) , .A1( u2_uk_n220 ) );
  OAI22_X1 u2_uk_U343 (.ZN( u2_K2_4 ) , .B1( u2_uk_n10 ) , .B2( u2_uk_n1238 ) , .A2( u2_uk_n1267 ) , .A1( u2_uk_n129 ) );
  OAI22_X1 u2_uk_U532 (.ZN( u2_K2_2 ) , .B2( u2_uk_n1243 ) , .A2( u2_uk_n1275 ) , .A1( u2_uk_n213 ) , .B1( u2_uk_n31 ) );
  OAI22_X1 u2_uk_U830 (.ZN( u2_K2_6 ) , .B2( u2_uk_n1249 ) , .A2( u2_uk_n1270 ) , .B1( u2_uk_n142 ) , .A1( u2_uk_n99 ) );
  OAI22_X1 u2_uk_U836 (.ZN( u2_K2_3 ) , .B2( u2_uk_n1239 ) , .A2( u2_uk_n1254 ) , .B1( u2_uk_n129 ) , .A1( u2_uk_n83 ) );
endmodule

