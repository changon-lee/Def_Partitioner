module aes_aes_die_18 ( sa10_0, sa10_1, sa10_2, sa10_3, sa10_4, sa10_5, sa10_6, sa10_7, sa13_sr_0, sa13_sr_1, sa13_sr_2, sa13_sr_3, sa13_sr_4, sa13_sr_5, sa13_sr_6, sa13_sr_7 );
  input sa10_0, sa10_1, sa10_2, sa10_3, sa10_4, sa10_5, sa10_6, sa10_7;
  output sa13_sr_0, sa13_sr_1, sa13_sr_2, sa13_sr_3, sa13_sr_4, sa13_sr_5, sa13_sr_6, sa13_sr_7;
  wire us10_n438, us10_n439, us10_n440, us10_n441, us10_n442, us10_n443, us10_n444, us10_n445, us10_n446, 
       us10_n447, us10_n448, us10_n449, us10_n450, us10_n451, us10_n452, us10_n453, us10_n454, us10_n455, 
       us10_n456, us10_n457, us10_n458, us10_n459, us10_n460, us10_n461, us10_n462, us10_n463, us10_n464, 
       us10_n465, us10_n466, us10_n467, us10_n468, us10_n469, us10_n470, us10_n471, us10_n472, us10_n473, 
       us10_n474, us10_n475, us10_n476, us10_n477, us10_n478, us10_n479, us10_n480, us10_n481, us10_n482, 
       us10_n483, us10_n484, us10_n485, us10_n486, us10_n487, us10_n488, us10_n489, us10_n490, us10_n491, 
       us10_n492, us10_n493, us10_n494, us10_n495, us10_n496, us10_n497, us10_n498, us10_n499, us10_n500, 
       us10_n501, us10_n502, us10_n503, us10_n504, us10_n505, us10_n506, us10_n507, us10_n508, us10_n509, 
       us10_n510, us10_n511, us10_n512, us10_n513, us10_n514, us10_n515, us10_n516, us10_n517, us10_n518, 
       us10_n519, us10_n520, us10_n521, us10_n522, us10_n523, us10_n524, us10_n525, us10_n526, us10_n527, 
       us10_n528, us10_n529, us10_n530, us10_n531, us10_n532, us10_n533, us10_n534, us10_n535, us10_n536, 
       us10_n537, us10_n538, us10_n539, us10_n540, us10_n541, us10_n542, us10_n543, us10_n544, us10_n545, 
       us10_n546, us10_n547, us10_n548, us10_n549, us10_n550, us10_n551, us10_n552, us10_n553, us10_n554, 
       us10_n555, us10_n556, us10_n557, us10_n558, us10_n559, us10_n560, us10_n561, us10_n562, us10_n563, 
       us10_n564, us10_n565, us10_n566, us10_n567, us10_n568, us10_n569, us10_n570, us10_n571, us10_n572, 
       us10_n573, us10_n574, us10_n575, us10_n576, us10_n577, us10_n578, us10_n579, us10_n580, us10_n581, 
       us10_n582, us10_n583, us10_n584, us10_n585, us10_n586, us10_n587, us10_n588, us10_n589, us10_n590, 
       us10_n591, us10_n592, us10_n593, us10_n594, us10_n595, us10_n596, us10_n597, us10_n598, us10_n599, 
       us10_n600, us10_n601, us10_n602, us10_n603, us10_n604, us10_n605, us10_n606, us10_n607, us10_n608, 
       us10_n609, us10_n610, us10_n611, us10_n612, us10_n613, us10_n614, us10_n615, us10_n616, us10_n617, 
       us10_n618, us10_n619, us10_n620, us10_n621, us10_n622, us10_n623, us10_n624, us10_n625, us10_n626, 
       us10_n627, us10_n628, us10_n629, us10_n630, us10_n631, us10_n632, us10_n633, us10_n634, us10_n635, 
       us10_n636, us10_n637, us10_n638, us10_n639, us10_n640, us10_n641, us10_n642, us10_n643, us10_n644, 
       us10_n645, us10_n646, us10_n647, us10_n648, us10_n649, us10_n650, us10_n651, us10_n652, us10_n653, 
       us10_n654, us10_n655, us10_n656, us10_n657, us10_n658, us10_n659, us10_n660, us10_n661, us10_n662, 
       us10_n663, us10_n664, us10_n665, us10_n666, us10_n667, us10_n668, us10_n669, us10_n670, us10_n671, 
       us10_n672, us10_n673, us10_n674, us10_n675, us10_n676, us10_n677, us10_n678, us10_n679, us10_n680, 
       us10_n681, us10_n682, us10_n683, us10_n684, us10_n685, us10_n686, us10_n687, us10_n688, us10_n689, 
       us10_n690, us10_n691, us10_n692, us10_n693, us10_n694, us10_n695, us10_n696, us10_n697, us10_n698, 
       us10_n699, us10_n700, us10_n701, us10_n702, us10_n703, us10_n704, us10_n705, us10_n706, us10_n707, 
       us10_n708, us10_n709, us10_n710, us10_n711, us10_n712, us10_n713, us10_n714, us10_n715, us10_n716, 
       us10_n717, us10_n718, us10_n719, us10_n720, us10_n721, us10_n722, us10_n723, us10_n724, us10_n725, 
       us10_n726, us10_n727, us10_n728, us10_n729, us10_n730, us10_n731, us10_n732, us10_n733, us10_n734, 
       us10_n735, us10_n736, us10_n737, us10_n738, us10_n739, us10_n740, us10_n741, us10_n742, us10_n743, 
       us10_n744, us10_n745, us10_n746, us10_n747, us10_n748, us10_n749, us10_n750, us10_n751, us10_n752, 
       us10_n753, us10_n754, us10_n755, us10_n756, us10_n757, us10_n758, us10_n759, us10_n760, us10_n761, 
       us10_n762, us10_n763, us10_n764, us10_n765, us10_n766, us10_n767, us10_n768, us10_n769, us10_n770, 
       us10_n771, us10_n772, us10_n773, us10_n774, us10_n775, us10_n776, us10_n777, us10_n778, us10_n779, 
       us10_n780, us10_n781, us10_n782, us10_n783, us10_n784, us10_n785, us10_n786, us10_n787, us10_n788, 
       us10_n789, us10_n790, us10_n791, us10_n792, us10_n793, us10_n794, us10_n795, us10_n796, us10_n797, 
       us10_n798, us10_n799, us10_n800, us10_n801, us10_n802, us10_n803, us10_n804, us10_n805, us10_n806, 
       us10_n807, us10_n808, us10_n809, us10_n810, us10_n811, us10_n812, us10_n813, us10_n814, us10_n815, 
       us10_n816, us10_n817, us10_n818, us10_n819, us10_n820, us10_n821, us10_n822, us10_n823, us10_n824, 
       us10_n825, us10_n826, us10_n827, us10_n828, us10_n829, us10_n830, us10_n831, us10_n832, us10_n833, 
       us10_n834, us10_n835, us10_n836, us10_n837, us10_n838, us10_n839, us10_n840, us10_n841, us10_n842, 
       us10_n843, us10_n844, us10_n845, us10_n846, us10_n847, us10_n848, us10_n849, us10_n850, us10_n851, 
       us10_n852, us10_n853, us10_n854, us10_n855, us10_n856, us10_n857, us10_n858, us10_n859, us10_n860, 
       us10_n861, us10_n862, us10_n863, us10_n864, us10_n865, us10_n866, us10_n867, us10_n868, us10_n869, 
       us10_n870, us10_n871, us10_n872, us10_n873, us10_n874, us10_n875,  us10_n876;
  NOR2_X1 us10_U10 (.A1( us10_n678 ) , .ZN( us10_n693 ) , .A2( us10_n807 ) );
  NOR3_X1 us10_U100 (.ZN( us10_n549 ) , .A2( us10_n651 ) , .A1( us10_n667 ) , .A3( us10_n771 ) );
  AOI211_X1 us10_U101 (.B( us10_n539 ) , .A( us10_n540 ) , .ZN( us10_n551 ) , .C2( us10_n839 ) , .C1( us10_n851 ) );
  NOR4_X1 us10_U102 (.A4( us10_n544 ) , .A3( us10_n545 ) , .A2( us10_n546 ) , .A1( us10_n547 ) , .ZN( us10_n548 ) );
  NOR4_X1 us10_U103 (.ZN( us10_n620 ) , .A1( us10_n656 ) , .A3( us10_n666 ) , .A4( us10_n682 ) , .A2( us10_n766 ) );
  NOR4_X1 us10_U104 (.A4( us10_n609 ) , .A3( us10_n610 ) , .A2( us10_n611 ) , .A1( us10_n612 ) , .ZN( us10_n619 ) );
  NOR4_X1 us10_U105 (.A4( us10_n614 ) , .A3( us10_n615 ) , .A2( us10_n616 ) , .A1( us10_n617 ) , .ZN( us10_n618 ) );
  NAND4_X1 us10_U106 (.A4( us10_n485 ) , .A3( us10_n486 ) , .A2( us10_n487 ) , .A1( us10_n488 ) , .ZN( us10_n778 ) );
  NOR4_X1 us10_U107 (.A4( us10_n484 ) , .ZN( us10_n487 ) , .A1( us10_n566 ) , .A2( us10_n581 ) , .A3( us10_n602 ) );
  NOR4_X1 us10_U108 (.ZN( us10_n486 ) , .A1( us10_n507 ) , .A2( us10_n519 ) , .A4( us10_n546 ) , .A3( us10_n611 ) );
  NOR4_X1 us10_U109 (.ZN( us10_n485 ) , .A2( us10_n533 ) , .A1( us10_n558 ) , .A3( us10_n631 ) , .A4( us10_n718 ) );
  INV_X1 us10_U11 (.A( us10_n680 ) , .ZN( us10_n840 ) );
  NAND4_X1 us10_U110 (.A4( us10_n691 ) , .A3( us10_n692 ) , .A1( us10_n693 ) , .ZN( us10_n776 ) , .A2( us10_n872 ) );
  AOI221_X1 us10_U111 (.A( us10_n681 ) , .ZN( us10_n692 ) , .B2( us10_n840 ) , .C1( us10_n842 ) , .C2( us10_n862 ) , .B1( us10_n865 ) );
  INV_X1 us10_U112 (.A( us10_n679 ) , .ZN( us10_n872 ) );
  NOR4_X1 us10_U113 (.A4( us10_n687 ) , .A3( us10_n688 ) , .A2( us10_n689 ) , .A1( us10_n690 ) , .ZN( us10_n691 ) );
  NAND4_X1 us10_U114 (.A4( us10_n473 ) , .A3( us10_n474 ) , .A2( us10_n475 ) , .A1( us10_n476 ) , .ZN( us10_n678 ) );
  NOR4_X1 us10_U115 (.A4( us10_n470 ) , .ZN( us10_n476 ) , .A3( us10_n556 ) , .A1( us10_n735 ) , .A2( us10_n755 ) );
  NOR4_X1 us10_U116 (.ZN( us10_n475 ) , .A1( us10_n531 ) , .A3( us10_n568 ) , .A4( us10_n600 ) , .A2( us10_n642 ) );
  NOR4_X1 us10_U117 (.ZN( us10_n474 ) , .A1( us10_n506 ) , .A3( us10_n544 ) , .A2( us10_n583 ) , .A4( us10_n716 ) );
  NAND4_X1 us10_U118 (.A4( us10_n719 ) , .A3( us10_n720 ) , .A2( us10_n721 ) , .ZN( us10_n741 ) , .A1( us10_n857 ) );
  INV_X1 us10_U119 (.A( us10_n709 ) , .ZN( us10_n857 ) );
  NOR4_X1 us10_U12 (.A4( us10_n445 ) , .A3( us10_n446 ) , .A2( us10_n516 ) , .A1( us10_n541 ) , .ZN( us10_n706 ) );
  NOR4_X1 us10_U120 (.A4( us10_n715 ) , .A3( us10_n716 ) , .A2( us10_n717 ) , .A1( us10_n718 ) , .ZN( us10_n719 ) );
  AOI221_X1 us10_U121 (.A( us10_n710 ) , .ZN( us10_n721 ) , .C2( us10_n844 ) , .B2( us10_n845 ) , .C1( us10_n861 ) , .B1( us10_n862 ) );
  NOR2_X1 us10_U122 (.ZN( us10_n789 ) , .A2( us10_n862 ) , .A1( us10_n868 ) );
  NOR2_X1 us10_U123 (.ZN( us10_n733 ) , .A2( us10_n832 ) , .A1( us10_n845 ) );
  NAND4_X1 us10_U124 (.A4( us10_n573 ) , .A3( us10_n574 ) , .A1( us10_n575 ) , .ZN( us10_n723 ) , .A2( us10_n874 ) );
  NOR4_X1 us10_U125 (.A4( us10_n569 ) , .A3( us10_n570 ) , .A2( us10_n571 ) , .A1( us10_n572 ) , .ZN( us10_n573 ) );
  AOI221_X1 us10_U126 (.A( us10_n564 ) , .C2( us10_n565 ) , .ZN( us10_n574 ) , .B2( us10_n845 ) , .B1( us10_n852 ) , .C1( us10_n853 ) );
  INV_X1 us10_U127 (.A( us10_n607 ) , .ZN( us10_n874 ) );
  NAND4_X1 us10_U128 (.A4( us10_n633 ) , .A3( us10_n634 ) , .A2( us10_n635 ) , .A1( us10_n636 ) , .ZN( us10_n743 ) );
  AOI211_X1 us10_U129 (.B( us10_n623 ) , .A( us10_n624 ) , .ZN( us10_n635 ) , .C2( us10_n836 ) , .C1( us10_n863 ) );
  OR3_X1 us10_U13 (.ZN( us10_n446 ) , .A1( us10_n528 ) , .A3( us10_n577 ) , .A2( us10_n875 ) );
  NOR4_X1 us10_U130 (.A4( us10_n629 ) , .A3( us10_n630 ) , .A2( us10_n631 ) , .A1( us10_n632 ) , .ZN( us10_n633 ) );
  NOR4_X1 us10_U131 (.A4( us10_n626 ) , .A3( us10_n627 ) , .A2( us10_n628 ) , .ZN( us10_n634 ) , .A1( us10_n664 ) );
  NAND4_X1 us10_U132 (.A4( us10_n493 ) , .A3( us10_n494 ) , .A1( us10_n495 ) , .ZN( us10_n802 ) , .A2( us10_n867 ) );
  AOI221_X1 us10_U133 (.A( us10_n489 ) , .ZN( us10_n494 ) , .B2( us10_n836 ) , .C2( us10_n841 ) , .C1( us10_n851 ) , .B1( us10_n860 ) );
  INV_X1 us10_U134 (.A( us10_n778 ) , .ZN( us10_n867 ) );
  NOR2_X1 us10_U135 (.ZN( us10_n495 ) , .A1( us10_n678 ) , .A2( us10_n694 ) );
  NOR2_X1 us10_U136 (.ZN( us10_n748 ) , .A1( us10_n861 ) , .A2( us10_n862 ) );
  NOR2_X1 us10_U137 (.ZN( us10_n647 ) , .A1( us10_n854 ) , .A2( us10_n868 ) );
  INV_X1 us10_U138 (.A( us10_n762 ) , .ZN( us10_n830 ) );
  OR4_X1 us10_U139 (.ZN( us10_n466 ) , .A4( us10_n518 ) , .A3( us10_n529 ) , .A2( us10_n578 ) , .A1( us10_n712 ) );
  OR4_X1 us10_U14 (.A4( us10_n442 ) , .A2( us10_n443 ) , .A1( us10_n444 ) , .ZN( us10_n445 ) , .A3( us10_n553 ) );
  OR4_X1 us10_U140 (.A4( us10_n566 ) , .A3( us10_n567 ) , .A2( us10_n568 ) , .ZN( us10_n572 ) , .A1( us10_n665 ) );
  OR4_X1 us10_U141 (.A4( us10_n518 ) , .A2( us10_n519 ) , .A1( us10_n520 ) , .ZN( us10_n522 ) , .A3( us10_n821 ) );
  OR4_X1 us10_U142 (.A4( us10_n682 ) , .A3( us10_n683 ) , .A2( us10_n684 ) , .A1( us10_n685 ) , .ZN( us10_n690 ) );
  OR4_X1 us10_U143 (.A4( us10_n580 ) , .A3( us10_n581 ) , .A2( us10_n582 ) , .A1( us10_n583 ) , .ZN( us10_n584 ) );
  NAND2_X1 us10_U144 (.ZN( us10_n613 ) , .A2( us10_n837 ) , .A1( us10_n873 ) );
  OR3_X1 us10_U145 (.A3( us10_n506 ) , .A2( us10_n507 ) , .A1( us10_n508 ) , .ZN( us10_n511 ) );
  INV_X1 us10_U146 (.A( us10_n672 ) , .ZN( us10_n859 ) );
  AOI21_X1 us10_U147 (.A( us10_n670 ) , .B1( us10_n671 ) , .ZN( us10_n672 ) , .B2( us10_n856 ) );
  INV_X1 us10_U148 (.A( us10_n754 ) , .ZN( us10_n869 ) );
  OAI21_X1 us10_U149 (.B1( us10_n753 ) , .ZN( us10_n754 ) , .A( us10_n845 ) , .B2( us10_n868 ) );
  INV_X1 us10_U15 (.A( us10_n613 ) , .ZN( us10_n875 ) );
  INV_X1 us10_U150 (.A( us10_n463 ) , .ZN( us10_n864 ) );
  OAI21_X1 us10_U151 (.ZN( us10_n463 ) , .B1( us10_n809 ) , .A( us10_n834 ) , .B2( us10_n851 ) );
  AOI222_X1 us10_U152 (.ZN( us10_n660 ) , .A2( us10_n839 ) , .B1( us10_n841 ) , .C2( us10_n845 ) , .A1( us10_n860 ) , .C1( us10_n863 ) , .B2( us10_n870 ) );
  INV_X1 us10_U153 (.A( us10_n647 ) , .ZN( us10_n870 ) );
  NAND2_X1 us10_U154 (.A1( us10_n447 ) , .A2( us10_n465 ) , .ZN( us10_n749 ) );
  OAI222_X1 us10_U155 (.B2( us10_n708 ) , .ZN( us10_n709 ) , .C2( us10_n724 ) , .B1( us10_n747 ) , .A1( us10_n806 ) , .C1( us10_n814 ) , .A2( us10_n815 ) );
  OAI222_X1 us10_U156 (.A2( us10_n669 ) , .ZN( us10_n674 ) , .B1( us10_n747 ) , .B2( us10_n784 ) , .C2( us10_n788 ) , .C1( us10_n815 ) , .A1( us10_n817 ) );
  OAI222_X1 us10_U157 (.ZN( us10_n617 ) , .B1( us10_n697 ) , .C1( us10_n724 ) , .C2( us10_n747 ) , .B2( us10_n786 ) , .A2( us10_n792 ) , .A1( us10_n816 ) );
  NOR4_X1 us10_U158 (.A2( us10_n491 ) , .A1( us10_n492 ) , .ZN( us10_n493 ) , .A3( us10_n580 ) , .A4( us10_n612 ) );
  OR4_X1 us10_U159 (.ZN( us10_n492 ) , .A4( us10_n534 ) , .A2( us10_n547 ) , .A1( us10_n559 ) , .A3( us10_n632 ) );
  INV_X1 us10_U16 (.A( us10_n749 ) , .ZN( us10_n863 ) );
  OAI22_X1 us10_U160 (.B1( us10_n490 ) , .ZN( us10_n491 ) , .A1( us10_n686 ) , .A2( us10_n763 ) , .B2( us10_n817 ) );
  NOR3_X1 us10_U161 (.ZN( us10_n490 ) , .A1( us10_n782 ) , .A2( us10_n850 ) , .A3( us10_n863 ) );
  INV_X1 us10_U162 (.A( us10_n730 ) , .ZN( us10_n839 ) );
  AOI221_X1 us10_U163 (.A( us10_n450 ) , .ZN( us10_n459 ) , .C2( us10_n753 ) , .B1( us10_n832 ) , .C1( us10_n842 ) , .B2( us10_n861 ) );
  AOI21_X1 us10_U164 (.ZN( us10_n450 ) , .B2( us10_n792 ) , .A( us10_n803 ) , .B1( us10_n815 ) );
  AOI221_X1 us10_U165 (.A( us10_n483 ) , .ZN( us10_n488 ) , .B1( us10_n831 ) , .C2( us10_n844 ) , .C1( us10_n852 ) , .B2( us10_n862 ) );
  OAI22_X1 us10_U166 (.ZN( us10_n483 ) , .A1( us10_n708 ) , .B2( us10_n785 ) , .A2( us10_n806 ) , .B1( us10_n812 ) );
  INV_X1 us10_U167 (.A( us10_n790 ) , .ZN( us10_n832 ) );
  NAND2_X1 us10_U168 (.A1( us10_n451 ) , .A2( us10_n453 ) , .ZN( us10_n762 ) );
  INV_X1 us10_U169 (.A( us10_n786 ) , .ZN( us10_n862 ) );
  AOI222_X1 us10_U17 (.ZN( us10_n605 ) , .B2( us10_n671 ) , .B1( us10_n753 ) , .C2( us10_n831 ) , .A1( us10_n833 ) , .A2( us10_n862 ) , .C1( us10_n863 ) );
  OAI221_X1 us10_U170 (.A( us10_n783 ) , .C2( us10_n784 ) , .B2( us10_n785 ) , .B1( us10_n786 ) , .ZN( us10_n796 ) , .C1( us10_n813 ) );
  AOI22_X1 us10_U171 (.A2( us10_n782 ) , .ZN( us10_n783 ) , .B2( us10_n831 ) , .A1( us10_n834 ) , .B1( us10_n863 ) );
  OAI221_X1 us10_U172 (.A( us10_n696 ) , .ZN( us10_n703 ) , .C2( us10_n784 ) , .C1( us10_n785 ) , .B1( us10_n786 ) , .B2( us10_n806 ) );
  AOI22_X1 us10_U173 (.ZN( us10_n696 ) , .A1( us10_n830 ) , .B2( us10_n843 ) , .A2( us10_n865 ) , .B1( us10_n868 ) );
  OAI221_X1 us10_U174 (.A( us10_n727 ) , .C2( us10_n728 ) , .B2( us10_n729 ) , .B1( us10_n730 ) , .ZN( us10_n737 ) , .C1( us10_n817 ) );
  AOI22_X1 us10_U175 (.ZN( us10_n727 ) , .B1( us10_n832 ) , .A2( us10_n838 ) , .A1( us10_n863 ) , .B2( us10_n866 ) );
  INV_X1 us10_U176 (.A( us10_n784 ) , .ZN( us10_n861 ) );
  OAI22_X1 us10_U177 (.ZN( us10_n710 ) , .A2( us10_n728 ) , .B2( us10_n729 ) , .A1( us10_n744 ) , .B1( us10_n813 ) );
  INV_X1 us10_U178 (.A( us10_n816 ) , .ZN( us10_n831 ) );
  INV_X1 us10_U179 (.A( us10_n788 ) , .ZN( us10_n845 ) );
  AOI222_X1 us10_U18 (.ZN( us10_n563 ) , .B1( us10_n830 ) , .C1( us10_n841 ) , .A2( us10_n843 ) , .A1( us10_n854 ) , .B2( us10_n863 ) , .C2( us10_n873 ) );
  OAI22_X1 us10_U180 (.ZN( us10_n588 ) , .A2( us10_n747 ) , .B2( us10_n762 ) , .A1( us10_n763 ) , .B1( us10_n784 ) );
  OAI22_X1 us10_U181 (.ZN( us10_n489 ) , .A1( us10_n724 ) , .B2( us10_n728 ) , .B1( us10_n730 ) , .A2( us10_n779 ) );
  OAI22_X1 us10_U182 (.ZN( us10_n624 ) , .B1( us10_n669 ) , .B2( us10_n747 ) , .A1( us10_n815 ) , .A2( us10_n816 ) );
  INV_X1 us10_U183 (.A( us10_n744 ) , .ZN( us10_n837 ) );
  OAI22_X1 us10_U184 (.ZN( us10_n681 ) , .A1( us10_n699 ) , .A2( us10_n730 ) , .B2( us10_n784 ) , .B1( us10_n817 ) );
  OAI22_X1 us10_U185 (.B2( us10_n779 ) , .B1( us10_n780 ) , .ZN( us10_n781 ) , .A2( us10_n814 ) , .A1( us10_n815 ) );
  OAI22_X1 us10_U186 (.A1( us10_n724 ) , .ZN( us10_n726 ) , .B2( us10_n750 ) , .B1( us10_n812 ) , .A2( us10_n816 ) );
  INV_X1 us10_U187 (.A( us10_n814 ) , .ZN( us10_n833 ) );
  OAI22_X1 us10_U188 (.B2( us10_n744 ) , .ZN( us10_n746 ) , .A2( us10_n762 ) , .B1( us10_n780 ) , .A1( us10_n792 ) );
  INV_X1 us10_U189 (.A( us10_n669 ) , .ZN( us10_n865 ) );
  NOR4_X1 us10_U19 (.ZN( us10_n473 ) , .A2( us10_n521 ) , .A4( us10_n594 ) , .A1( us10_n609 ) , .A3( us10_n629 ) );
  OAI22_X1 us10_U190 (.ZN( us10_n496 ) , .A2( us10_n744 ) , .A1( us10_n780 ) , .B1( us10_n791 ) , .B2( us10_n806 ) );
  INV_X1 us10_U191 (.A( us10_n750 ) , .ZN( us10_n842 ) );
  AOI211_X1 us10_U192 (.A( us10_n637 ) , .ZN( us10_n645 ) , .B( us10_n743 ) , .C2( us10_n839 ) , .C1( us10_n854 ) );
  OAI22_X1 us10_U193 (.ZN( us10_n637 ) , .A1( us10_n699 ) , .B2( us10_n728 ) , .A2( us10_n762 ) , .B1( us10_n816 ) );
  OAI22_X1 us10_U194 (.ZN( us10_n590 ) , .B1( us10_n730 ) , .B2( us10_n749 ) , .A2( us10_n786 ) , .A1( us10_n803 ) );
  OAI22_X1 us10_U195 (.ZN( us10_n695 ) , .A2( us10_n730 ) , .A1( us10_n780 ) , .B1( us10_n791 ) , .B2( us10_n817 ) );
  INV_X1 us10_U196 (.A( us10_n747 ) , .ZN( us10_n834 ) );
  NOR2_X1 us10_U197 (.A1( us10_n697 ) , .ZN( us10_n770 ) , .A2( us10_n815 ) );
  NOR2_X1 us10_U198 (.ZN( us10_n666 ) , .A1( us10_n728 ) , .A2( us10_n803 ) );
  NOR2_X1 us10_U199 (.ZN( us10_n594 ) , .A2( us10_n697 ) , .A1( us10_n728 ) );
  NOR4_X1 us10_U20 (.ZN( us10_n479 ) , .A1( us10_n520 ) , .A4( us10_n557 ) , .A3( us10_n582 ) , .A2( us10_n630 ) );
  NOR2_X1 us10_U200 (.ZN( us10_n600 ) , .A2( us10_n697 ) , .A1( us10_n784 ) );
  NOR2_X1 us10_U201 (.ZN( us10_n570 ) , .A1( us10_n728 ) , .A2( us10_n806 ) );
  NOR2_X1 us10_U202 (.ZN( us10_n532 ) , .A2( us10_n749 ) , .A1( us10_n750 ) );
  NOR2_X1 us10_U203 (.ZN( us10_n615 ) , .A1( us10_n785 ) , .A2( us10_n815 ) );
  NOR2_X1 us10_U204 (.ZN( us10_n629 ) , .A2( us10_n728 ) , .A1( us10_n785 ) );
  NOR2_X1 us10_U205 (.ZN( us10_n654 ) , .A1( us10_n728 ) , .A2( us10_n813 ) );
  NOR2_X1 us10_U206 (.ZN( us10_n546 ) , .A2( us10_n780 ) , .A1( us10_n814 ) );
  NOR2_X1 us10_U207 (.ZN( us10_n718 ) , .A2( us10_n724 ) , .A1( us10_n744 ) );
  NOR2_X1 us10_U208 (.ZN( us10_n577 ) , .A2( us10_n699 ) , .A1( us10_n814 ) );
  NOR2_X1 us10_U209 (.ZN( us10_n612 ) , .A1( us10_n779 ) , .A2( us10_n786 ) );
  NOR4_X1 us10_U21 (.A4( us10_n532 ) , .A3( us10_n533 ) , .A2( us10_n534 ) , .ZN( us10_n535 ) , .A1( us10_n820 ) );
  NOR2_X1 us10_U210 (.ZN( us10_n628 ) , .A2( us10_n669 ) , .A1( us10_n785 ) );
  NOR2_X1 us10_U211 (.ZN( us10_n610 ) , .A1( us10_n784 ) , .A2( us10_n816 ) );
  NOR2_X1 us10_U212 (.ZN( us10_n651 ) , .A1( us10_n784 ) , .A2( us10_n788 ) );
  NOR2_X1 us10_U213 (.ZN( us10_n531 ) , .A2( us10_n780 ) , .A1( us10_n816 ) );
  NOR2_X1 us10_U214 (.ZN( us10_n599 ) , .A2( us10_n791 ) , .A1( us10_n816 ) );
  INV_X1 us10_U215 (.A( us10_n728 ) , .ZN( us10_n852 ) );
  NOR2_X1 us10_U216 (.A2( us10_n708 ) , .A1( us10_n750 ) , .ZN( us10_n771 ) );
  NOR2_X1 us10_U217 (.A1( us10_n699 ) , .ZN( us10_n768 ) , .A2( us10_n813 ) );
  NOR2_X1 us10_U218 (.ZN( us10_n667 ) , .A1( us10_n750 ) , .A2( us10_n815 ) );
  NOR2_X1 us10_U219 (.ZN( us10_n541 ) , .A2( us10_n697 ) , .A1( us10_n699 ) );
  NOR4_X1 us10_U22 (.A4( us10_n541 ) , .A3( us10_n542 ) , .A2( us10_n543 ) , .ZN( us10_n550 ) , .A1( us10_n688 ) );
  NOR2_X1 us10_U220 (.ZN( us10_n508 ) , .A2( us10_n780 ) , .A1( us10_n785 ) );
  NOR2_X1 us10_U221 (.ZN( us10_n543 ) , .A2( us10_n708 ) , .A1( us10_n785 ) );
  NOR2_X1 us10_U222 (.ZN( us10_n555 ) , .A1( us10_n750 ) , .A2( us10_n791 ) );
  NOR2_X1 us10_U223 (.ZN( us10_n611 ) , .A2( us10_n780 ) , .A1( us10_n806 ) );
  NOR2_X1 us10_U224 (.ZN( us10_n664 ) , .A1( us10_n785 ) , .A2( us10_n791 ) );
  NOR2_X1 us10_U225 (.ZN( us10_n652 ) , .A1( us10_n669 ) , .A2( us10_n814 ) );
  NOR2_X1 us10_U226 (.A1( us10_n669 ) , .ZN( us10_n673 ) , .A2( us10_n744 ) );
  NOR2_X1 us10_U227 (.ZN( us10_n602 ) , .A1( us10_n669 ) , .A2( us10_n803 ) );
  NOR2_X1 us10_U228 (.A1( us10_n669 ) , .ZN( us10_n688 ) , .A2( us10_n816 ) );
  NOR2_X1 us10_U229 (.A2( us10_n744 ) , .ZN( us10_n769 ) , .A1( us10_n812 ) );
  AOI221_X1 us10_U23 (.A( us10_n713 ) , .B2( us10_n714 ) , .ZN( us10_n720 ) , .C1( us10_n832 ) , .B1( us10_n839 ) , .C2( us10_n863 ) );
  INV_X1 us10_U230 (.A( us10_n792 ) , .ZN( us10_n851 ) );
  NOR2_X1 us10_U231 (.A1( us10_n669 ) , .ZN( us10_n766 ) , .A2( us10_n813 ) );
  NOR2_X1 us10_U232 (.ZN( us10_n527 ) , .A1( us10_n669 ) , .A2( us10_n779 ) );
  NOR2_X1 us10_U233 (.A2( us10_n697 ) , .ZN( us10_n716 ) , .A1( us10_n792 ) );
  OAI22_X1 us10_U234 (.B1( us10_n440 ) , .ZN( us10_n444 ) , .A2( us10_n728 ) , .A1( us10_n744 ) , .B2( us10_n749 ) );
  NOR3_X1 us10_U235 (.ZN( us10_n440 ) , .A2( us10_n836 ) , .A3( us10_n837 ) , .A1( us10_n846 ) );
  NOR2_X1 us10_U236 (.ZN( us10_n601 ) , .A2( us10_n780 ) , .A1( us10_n803 ) );
  NOR2_X1 us10_U237 (.ZN( us10_n661 ) , .A1( us10_n729 ) , .A2( us10_n790 ) );
  NOR2_X1 us10_U238 (.ZN( us10_n631 ) , .A1( us10_n724 ) , .A2( us10_n813 ) );
  NOR2_X1 us10_U239 (.ZN( us10_n528 ) , .A2( us10_n724 ) , .A1( us10_n803 ) );
  OR2_X1 us10_U24 (.A2( us10_n711 ) , .A1( us10_n712 ) , .ZN( us10_n713 ) );
  NOR2_X1 us10_U240 (.ZN( us10_n509 ) , .A1( us10_n729 ) , .A2( us10_n779 ) );
  NOR2_X1 us10_U241 (.ZN( us10_n507 ) , .A1( us10_n812 ) , .A2( us10_n817 ) );
  NOR2_X1 us10_U242 (.ZN( us10_n662 ) , .A2( us10_n697 ) , .A1( us10_n729 ) );
  NOR2_X1 us10_U243 (.ZN( us10_n630 ) , .A1( us10_n747 ) , .A2( us10_n815 ) );
  NOR2_X1 us10_U244 (.ZN( us10_n554 ) , .A1( us10_n786 ) , .A2( us10_n813 ) );
  NOR2_X1 us10_U245 (.ZN( us10_n545 ) , .A1( us10_n749 ) , .A2( us10_n814 ) );
  NOR2_X1 us10_U246 (.ZN( us10_n557 ) , .A1( us10_n792 ) , .A2( us10_n814 ) );
  NOR2_X1 us10_U247 (.ZN( us10_n717 ) , .A2( us10_n744 ) , .A1( us10_n786 ) );
  NOR2_X1 us10_U248 (.ZN( us10_n544 ) , .A2( us10_n785 ) , .A1( us10_n792 ) );
  INV_X1 us10_U249 (.A( us10_n806 ) , .ZN( us10_n841 ) );
  NOR2_X1 us10_U25 (.ZN( us10_n680 ) , .A2( us10_n834 ) , .A1( us10_n839 ) );
  OAI21_X1 us10_U250 (.ZN( us10_n731 ) , .A( us10_n833 ) , .B2( us10_n852 ) , .B1( us10_n873 ) );
  NOR2_X1 us10_U251 (.A2( us10_n697 ) , .A1( us10_n780 ) , .ZN( us10_n820 ) );
  NOR2_X1 us10_U252 (.ZN( us10_n663 ) , .A1( us10_n729 ) , .A2( us10_n785 ) );
  OAI22_X1 us10_U253 (.B2( us10_n750 ) , .B1( us10_n751 ) , .A1( us10_n752 ) , .ZN( us10_n756 ) , .A2( us10_n806 ) );
  NOR2_X1 us10_U254 (.ZN( us10_n751 ) , .A2( us10_n852 ) , .A1( us10_n860 ) );
  NOR3_X1 us10_U255 (.ZN( us10_n752 ) , .A2( us10_n853 ) , .A1( us10_n863 ) , .A3( us10_n865 ) );
  NOR2_X1 us10_U256 (.ZN( us10_n656 ) , .A1( us10_n747 ) , .A2( us10_n780 ) );
  NOR2_X1 us10_U257 (.ZN( us10_n530 ) , .A2( us10_n744 ) , .A1( us10_n792 ) );
  NOR2_X1 us10_U258 (.ZN( us10_n506 ) , .A2( us10_n728 ) , .A1( us10_n762 ) );
  NOR2_X1 us10_U259 (.ZN( us10_n558 ) , .A1( us10_n708 ) , .A2( us10_n816 ) );
  NOR4_X1 us10_U26 (.A4( us10_n514 ) , .A3( us10_n515 ) , .A2( us10_n516 ) , .A1( us10_n517 ) , .ZN( us10_n524 ) );
  NOR2_X1 us10_U260 (.ZN( us10_n516 ) , .A1( us10_n708 ) , .A2( us10_n744 ) );
  NOR2_X1 us10_U261 (.ZN( us10_n614 ) , .A1( us10_n762 ) , .A2( us10_n812 ) );
  AOI21_X1 us10_U262 (.A( us10_n812 ) , .B2( us10_n813 ) , .B1( us10_n814 ) , .ZN( us10_n819 ) );
  NOR2_X1 us10_U263 (.A1( us10_n749 ) , .ZN( us10_n767 ) , .A2( us10_n803 ) );
  AOI21_X1 us10_U264 (.ZN( us10_n593 ) , .B1( us10_n750 ) , .A( us10_n792 ) , .B2( us10_n813 ) );
  NOR2_X1 us10_U265 (.A1( us10_n730 ) , .ZN( us10_n765 ) , .A2( us10_n786 ) );
  NOR2_X1 us10_U266 (.ZN( us10_n655 ) , .A1( us10_n790 ) , .A2( us10_n815 ) );
  NOR2_X1 us10_U267 (.ZN( us10_n701 ) , .A2( us10_n786 ) , .A1( us10_n817 ) );
  NOR2_X1 us10_U268 (.ZN( us10_n579 ) , .A2( us10_n708 ) , .A1( us10_n730 ) );
  NOR2_X1 us10_U269 (.ZN( us10_n533 ) , .A2( us10_n724 ) , .A1( us10_n730 ) );
  AOI222_X1 us10_U27 (.ZN( us10_n525 ) , .A1( us10_n834 ) , .B2( us10_n837 ) , .C1( us10_n844 ) , .C2( us10_n850 ) , .A2( us10_n852 ) , .B1( us10_n866 ) );
  NOR2_X1 us10_U270 (.ZN( us10_n668 ) , .A2( us10_n708 ) , .A1( us10_n790 ) );
  INV_X1 us10_U271 (.A( us10_n813 ) , .ZN( us10_n836 ) );
  NOR2_X1 us10_U272 (.ZN( us10_n521 ) , .A1( us10_n790 ) , .A2( us10_n812 ) );
  AOI21_X1 us10_U273 (.ZN( us10_n571 ) , .B2( us10_n697 ) , .B1( us10_n806 ) , .A( us10_n812 ) );
  INV_X1 us10_U274 (.A( us10_n763 ) , .ZN( us10_n866 ) );
  NOR2_X1 us10_U275 (.ZN( us10_n517 ) , .A1( us10_n708 ) , .A2( us10_n803 ) );
  AOI21_X1 us10_U276 (.A( us10_n815 ) , .B2( us10_n816 ) , .B1( us10_n817 ) , .ZN( us10_n818 ) );
  INV_X1 us10_U277 (.A( us10_n729 ) , .ZN( us10_n868 ) );
  NOR2_X1 us10_U278 (.ZN( us10_n542 ) , .A1( us10_n762 ) , .A2( us10_n791 ) );
  AOI21_X1 us10_U279 (.ZN( us10_n499 ) , .B1( us10_n680 ) , .A( us10_n812 ) , .B2( us10_n816 ) );
  NOR4_X1 us10_U28 (.A3( us10_n521 ) , .A1( us10_n522 ) , .ZN( us10_n523 ) , .A2( us10_n673 ) , .A4( us10_n769 ) );
  NOR2_X1 us10_U280 (.ZN( us10_n609 ) , .A2( us10_n724 ) , .A1( us10_n817 ) );
  NOR2_X1 us10_U281 (.ZN( us10_n642 ) , .A2( us10_n788 ) , .A1( us10_n791 ) );
  AOI21_X1 us10_U282 (.ZN( us10_n592 ) , .B1( us10_n728 ) , .B2( us10_n784 ) , .A( us10_n790 ) );
  NOR2_X1 us10_U283 (.ZN( us10_n653 ) , .A1( us10_n762 ) , .A2( us10_n786 ) );
  AOI21_X1 us10_U284 (.B1( us10_n625 ) , .ZN( us10_n627 ) , .A( us10_n763 ) , .B2( us10_n814 ) );
  AOI21_X1 us10_U285 (.ZN( us10_n478 ) , .B2( us10_n697 ) , .A( us10_n749 ) , .B1( us10_n779 ) );
  AOI21_X1 us10_U286 (.ZN( us10_n648 ) , .A( us10_n762 ) , .B2( us10_n784 ) , .B1( us10_n792 ) );
  AOI21_X1 us10_U287 (.ZN( us10_n623 ) , .B1( us10_n699 ) , .A( us10_n779 ) , .B2( us10_n784 ) );
  NOR2_X1 us10_U288 (.ZN( us10_n582 ) , .A1( us10_n744 ) , .A2( us10_n815 ) );
  NOR2_X1 us10_U289 (.A2( us10_n708 ) , .A1( us10_n762 ) , .ZN( us10_n794 ) );
  AOI221_X1 us10_U29 (.A( us10_n781 ) , .ZN( us10_n798 ) , .C2( us10_n837 ) , .B2( us10_n838 ) , .B1( us10_n865 ) , .C1( us10_n866 ) );
  NOR2_X1 us10_U290 (.ZN( us10_n553 ) , .A2( us10_n744 ) , .A1( us10_n784 ) );
  NOR2_X1 us10_U291 (.ZN( us10_n519 ) , .A2( us10_n699 ) , .A1( us10_n816 ) );
  AOI21_X1 us10_U292 (.ZN( us10_n626 ) , .B2( us10_n669 ) , .A( us10_n790 ) , .B1( us10_n791 ) );
  NOR2_X1 us10_U293 (.ZN( us10_n520 ) , .A2( us10_n708 ) , .A1( us10_n814 ) );
  AOI21_X1 us10_U294 (.ZN( us10_n477 ) , .A( us10_n669 ) , .B1( us10_n750 ) , .B2( us10_n806 ) );
  AOI21_X1 us10_U295 (.ZN( us10_n589 ) , .B2( us10_n699 ) , .B1( us10_n815 ) , .A( us10_n817 ) );
  AOI21_X1 us10_U296 (.ZN( us10_n510 ) , .B2( us10_n669 ) , .A( us10_n730 ) , .B1( us10_n815 ) );
  AOI21_X1 us10_U297 (.ZN( us10_n540 ) , .A( us10_n763 ) , .B2( us10_n779 ) , .B1( us10_n817 ) );
  AOI21_X1 us10_U298 (.ZN( us10_n515 ) , .A( us10_n729 ) , .B1( us10_n750 ) , .B2( us10_n803 ) );
  NOR2_X1 us10_U299 (.ZN( us10_n547 ) , .A1( us10_n699 ) , .A2( us10_n744 ) );
  NAND4_X1 us10_U3 (.ZN( sa13_sr_0 ) , .A4( us10_n501 ) , .A3( us10_n502 ) , .A2( us10_n503 ) , .A1( us10_n504 ) );
  NOR4_X1 us10_U30 (.A4( us10_n793 ) , .A3( us10_n794 ) , .A2( us10_n795 ) , .A1( us10_n796 ) , .ZN( us10_n797 ) );
  NOR2_X1 us10_U300 (.ZN( us10_n581 ) , .A1( us10_n669 ) , .A2( us10_n788 ) );
  AOI21_X1 us10_U301 (.ZN( us10_n539 ) , .B2( us10_n812 ) , .A( us10_n814 ) , .B1( us10_n815 ) );
  NOR2_X1 us10_U302 (.ZN( us10_n559 ) , .A2( us10_n791 ) , .A1( us10_n803 ) );
  AOI21_X1 us10_U303 (.ZN( us10_n498 ) , .A( us10_n724 ) , .B2( us10_n762 ) , .B1( us10_n814 ) );
  NAND2_X2 us10_U304 (.A2( us10_n461 ) , .A1( us10_n462 ) , .ZN( us10_n747 ) );
  AOI21_X1 us10_U305 (.B1( us10_n699 ) , .ZN( us10_n700 ) , .A( us10_n732 ) , .B2( us10_n763 ) );
  AOI21_X1 us10_U306 (.ZN( us10_n591 ) , .B2( us10_n763 ) , .A( us10_n785 ) , .B1( us10_n812 ) );
  AOI21_X1 us10_U307 (.ZN( us10_n640 ) , .B2( us10_n747 ) , .A( us10_n792 ) , .B1( us10_n803 ) );
  AOI21_X1 us10_U308 (.ZN( us10_n569 ) , .B1( us10_n750 ) , .B2( us10_n762 ) , .A( us10_n780 ) );
  NOR2_X1 us10_U309 (.ZN( us10_n683 ) , .A2( us10_n699 ) , .A1( us10_n803 ) );
  NOR4_X1 us10_U31 (.A4( us10_n776 ) , .A3( us10_n777 ) , .A1( us10_n778 ) , .ZN( us10_n799 ) , .A2( us10_n801 ) );
  NOR2_X1 us10_U310 (.ZN( us10_n665 ) , .A1( us10_n780 ) , .A2( us10_n813 ) );
  AOI21_X1 us10_U311 (.ZN( us10_n500 ) , .A( us10_n697 ) , .B1( us10_n708 ) , .B2( us10_n786 ) );
  NOR2_X1 us10_U312 (.ZN( us10_n685 ) , .A1( us10_n729 ) , .A2( us10_n816 ) );
  INV_X1 us10_U313 (.A( us10_n791 ) , .ZN( us10_n873 ) );
  AOI21_X1 us10_U314 (.ZN( us10_n649 ) , .B1( us10_n729 ) , .B2( us10_n763 ) , .A( us10_n813 ) );
  AOI21_X1 us10_U315 (.B1( us10_n686 ) , .ZN( us10_n687 ) , .A( us10_n728 ) , .B2( us10_n761 ) );
  INV_X1 us10_U316 (.A( us10_n699 ) , .ZN( us10_n853 ) );
  NOR2_X1 us10_U317 (.ZN( us10_n568 ) , .A1( us10_n729 ) , .A2( us10_n762 ) );
  NOR2_X1 us10_U318 (.ZN( us10_n578 ) , .A1( us10_n708 ) , .A2( us10_n813 ) );
  AOI21_X1 us10_U319 (.ZN( us10_n514 ) , .A( us10_n779 ) , .B2( us10_n792 ) , .B1( us10_n812 ) );
  NOR4_X1 us10_U32 (.A4( us10_n734 ) , .A3( us10_n735 ) , .A2( us10_n736 ) , .A1( us10_n737 ) , .ZN( us10_n738 ) );
  NOR2_X1 us10_U320 (.ZN( us10_n684 ) , .A1( us10_n791 ) , .A2( us10_n813 ) );
  NOR2_X1 us10_U321 (.ZN( us10_n580 ) , .A2( us10_n697 ) , .A1( us10_n791 ) );
  NOR2_X1 us10_U322 (.A2( us10_n813 ) , .A1( us10_n815 ) , .ZN( us10_n821 ) );
  NOR2_X1 us10_U323 (.ZN( us10_n566 ) , .A2( us10_n697 ) , .A1( us10_n763 ) );
  AOI21_X1 us10_U324 (.ZN( us10_n497 ) , .A( us10_n779 ) , .B2( us10_n791 ) , .B1( us10_n804 ) );
  AOI21_X1 us10_U325 (.ZN( us10_n564 ) , .B1( us10_n724 ) , .A( us10_n779 ) , .B2( us10_n791 ) );
  NOR2_X1 us10_U326 (.ZN( us10_n632 ) , .A2( us10_n697 ) , .A1( us10_n724 ) );
  NAND2_X2 us10_U327 (.A2( us10_n454 ) , .A1( us10_n472 ) , .ZN( us10_n779 ) );
  NOR2_X1 us10_U328 (.ZN( us10_n529 ) , .A1( us10_n708 ) , .A2( us10_n779 ) );
  AOI21_X1 us10_U329 (.ZN( us10_n639 ) , .B2( us10_n749 ) , .A( us10_n788 ) , .B1( us10_n812 ) );
  AOI211_X1 us10_U33 (.B( us10_n725 ) , .A( us10_n726 ) , .ZN( us10_n739 ) , .C1( us10_n843 ) , .C2( us10_n855 ) );
  AOI21_X1 us10_U330 (.ZN( us10_n689 ) , .B2( us10_n749 ) , .B1( us10_n763 ) , .A( us10_n806 ) );
  AOI21_X1 us10_U331 (.A( us10_n790 ) , .B2( us10_n791 ) , .B1( us10_n792 ) , .ZN( us10_n793 ) );
  AOI21_X1 us10_U332 (.A( us10_n733 ) , .ZN( us10_n734 ) , .B2( us10_n780 ) , .B1( us10_n792 ) );
  AOI21_X1 us10_U333 (.ZN( us10_n641 ) , .B1( us10_n680 ) , .A( us10_n791 ) , .B2( us10_n817 ) );
  NOR2_X1 us10_U334 (.ZN( us10_n583 ) , .A1( us10_n792 ) , .A2( us10_n817 ) );
  NOR2_X1 us10_U335 (.ZN( us10_n711 ) , .A1( us10_n762 ) , .A2( us10_n763 ) );
  NOR2_X1 us10_U336 (.ZN( us10_n534 ) , .A1( us10_n724 ) , .A2( us10_n788 ) );
  NOR2_X1 us10_U337 (.ZN( us10_n682 ) , .A2( us10_n708 ) , .A1( us10_n817 ) );
  INV_X1 us10_U338 (.A( us10_n697 ) , .ZN( us10_n838 ) );
  AOI21_X1 us10_U339 (.ZN( us10_n442 ) , .A( us10_n699 ) , .B1( us10_n733 ) , .B2( us10_n750 ) );
  NOR3_X1 us10_U34 (.A3( us10_n722 ) , .A1( us10_n723 ) , .ZN( us10_n740 ) , .A2( us10_n741 ) );
  NAND2_X2 us10_U340 (.A1( us10_n455 ) , .A2( us10_n462 ) , .ZN( us10_n750 ) );
  INV_X1 us10_U341 (.A( us10_n815 ) , .ZN( us10_n855 ) );
  OAI21_X1 us10_U342 (.A( us10_n613 ) , .ZN( us10_n616 ) , .B1( us10_n625 ) , .B2( us10_n784 ) );
  NAND2_X2 us10_U343 (.A1( us10_n462 ) , .A2( us10_n472 ) , .ZN( us10_n788 ) );
  OAI21_X1 us10_U344 (.A( us10_n698 ) , .ZN( us10_n702 ) , .B2( us10_n750 ) , .B1( us10_n804 ) );
  OAI21_X1 us10_U345 (.ZN( us10_n698 ) , .B2( us10_n833 ) , .B1( us10_n838 ) , .A( us10_n860 ) );
  INV_X1 us10_U346 (.A( us10_n785 ) , .ZN( us10_n846 ) );
  INV_X1 us10_U347 (.A( us10_n780 ) , .ZN( us10_n850 ) );
  OAI21_X1 us10_U348 (.A( us10_n787 ) , .B2( us10_n788 ) , .B1( us10_n789 ) , .ZN( us10_n795 ) );
  OAI21_X1 us10_U349 (.ZN( us10_n787 ) , .A( us10_n839 ) , .B1( us10_n863 ) , .B2( us10_n873 ) );
  NOR4_X1 us10_U35 (.A3( us10_n755 ) , .A2( us10_n756 ) , .A1( us10_n757 ) , .ZN( us10_n758 ) , .A4( us10_n869 ) );
  NAND2_X1 us10_U350 (.A1( us10_n729 ) , .A2( us10_n784 ) , .ZN( us10_n811 ) );
  NAND2_X1 us10_U351 (.ZN( us10_n671 ) , .A1( us10_n806 ) , .A2( us10_n816 ) );
  NAND2_X1 us10_U352 (.ZN( us10_n714 ) , .A1( us10_n728 ) , .A2( us10_n780 ) );
  AOI21_X1 us10_U353 (.ZN( us10_n443 ) , .B1( us10_n789 ) , .B2( us10_n791 ) , .A( us10_n814 ) );
  NOR2_X1 us10_U354 (.ZN( us10_n712 ) , .A2( us10_n724 ) , .A1( us10_n790 ) );
  NAND2_X1 us10_U355 (.A2( us10_n762 ) , .A1( us10_n806 ) , .ZN( us10_n810 ) );
  NAND2_X2 us10_U356 (.A1( us10_n454 ) , .A2( us10_n461 ) , .ZN( us10_n813 ) );
  NOR2_X1 us10_U357 (.ZN( us10_n470 ) , .A2( us10_n779 ) , .A1( us10_n815 ) );
  NAND2_X1 us10_U358 (.A1( us10_n699 ) , .A2( us10_n729 ) , .ZN( us10_n782 ) );
  NOR2_X1 us10_U359 (.ZN( us10_n526 ) , .A1( us10_n724 ) , .A2( us10_n750 ) );
  AOI211_X1 us10_U36 (.B( us10_n745 ) , .A( us10_n746 ) , .ZN( us10_n759 ) , .C1( us10_n832 ) , .C2( us10_n853 ) );
  NOR2_X1 us10_U360 (.ZN( us10_n518 ) , .A1( us10_n708 ) , .A2( us10_n788 ) );
  NAND2_X1 us10_U361 (.A2( us10_n749 ) , .A1( us10_n786 ) , .ZN( us10_n809 ) );
  INV_X1 us10_U362 (.A( us10_n817 ) , .ZN( us10_n844 ) );
  NAND2_X2 us10_U363 (.A1( us10_n451 ) , .A2( us10_n454 ) , .ZN( us10_n814 ) );
  INV_X1 us10_U364 (.A( us10_n724 ) , .ZN( us10_n856 ) );
  AND2_X1 us10_U365 (.ZN( us10_n732 ) , .A1( us10_n779 ) , .A2( us10_n785 ) );
  AOI221_X1 us10_U366 (.A( us10_n764 ) , .ZN( us10_n774 ) , .C2( us10_n810 ) , .B2( us10_n835 ) , .C1( us10_n855 ) , .B1( us10_n866 ) );
  AOI21_X1 us10_U367 (.B2( us10_n763 ) , .ZN( us10_n764 ) , .A( us10_n788 ) , .B1( us10_n792 ) );
  INV_X1 us10_U368 (.A( us10_n761 ) , .ZN( us10_n835 ) );
  NAND2_X1 us10_U369 (.A1( us10_n451 ) , .A2( us10_n471 ) , .ZN( us10_n816 ) );
  NOR3_X1 us10_U37 (.A3( us10_n741 ) , .A2( us10_n742 ) , .A1( us10_n743 ) , .ZN( us10_n760 ) );
  NAND2_X1 us10_U370 (.A2( us10_n441 ) , .A1( us10_n447 ) , .ZN( us10_n784 ) );
  NAND2_X1 us10_U371 (.A2( us10_n448 ) , .A1( us10_n460 ) , .ZN( us10_n728 ) );
  NAND2_X1 us10_U372 (.A1( us10_n453 ) , .A2( us10_n472 ) , .ZN( us10_n785 ) );
  NAND2_X1 us10_U373 (.A1( us10_n453 ) , .A2( us10_n461 ) , .ZN( us10_n744 ) );
  NAND2_X1 us10_U374 (.A1( us10_n452 ) , .A2( us10_n465 ) , .ZN( us10_n669 ) );
  NAND2_X1 us10_U375 (.A2( us10_n453 ) , .A1( us10_n455 ) , .ZN( us10_n806 ) );
  NAND2_X1 us10_U376 (.A1( us10_n441 ) , .A2( us10_n460 ) , .ZN( us10_n699 ) );
  NAND2_X1 us10_U377 (.A1( us10_n455 ) , .A2( us10_n471 ) , .ZN( us10_n803 ) );
  NAND2_X1 us10_U378 (.A2( us10_n464 ) , .A1( us10_n465 ) , .ZN( us10_n812 ) );
  NAND2_X1 us10_U379 (.A1( us10_n447 ) , .A2( us10_n448 ) , .ZN( us10_n786 ) );
  NAND4_X1 us10_U38 (.ZN( sa13_sr_3 ) , .A4( us10_n704 ) , .A3( us10_n705 ) , .A2( us10_n706 ) , .A1( us10_n707 ) );
  NAND2_X2 us10_U380 (.A2( us10_n461 ) , .A1( us10_n471 ) , .ZN( us10_n697 ) );
  NAND2_X1 us10_U381 (.A2( us10_n448 ) , .A1( us10_n452 ) , .ZN( us10_n729 ) );
  NAND2_X1 us10_U382 (.A2( us10_n449 ) , .A1( us10_n452 ) , .ZN( us10_n763 ) );
  NAND2_X1 us10_U383 (.A2( us10_n454 ) , .A1( us10_n455 ) , .ZN( us10_n730 ) );
  NOR2_X1 us10_U384 (.ZN( us10_n465 ) , .A2( us10_n847 ) , .A1( us10_n848 ) );
  NOR2_X1 us10_U385 (.ZN( us10_n453 ) , .A1( us10_n826 ) , .A2( us10_n827 ) );
  NOR2_X1 us10_U386 (.ZN( us10_n451 ) , .A1( us10_n828 ) , .A2( us10_n829 ) );
  NAND2_X1 us10_U387 (.A1( us10_n451 ) , .A2( us10_n462 ) , .ZN( us10_n790 ) );
  NAND2_X2 us10_U388 (.A2( us10_n448 ) , .A1( us10_n464 ) , .ZN( us10_n815 ) );
  NAND2_X2 us10_U389 (.A2( us10_n441 ) , .A1( us10_n452 ) , .ZN( us10_n791 ) );
  NOR4_X1 us10_U39 (.A4( us10_n700 ) , .A3( us10_n701 ) , .A2( us10_n702 ) , .A1( us10_n703 ) , .ZN( us10_n704 ) );
  NAND2_X2 us10_U390 (.A1( us10_n449 ) , .A2( us10_n464 ) , .ZN( us10_n724 ) );
  NAND2_X1 us10_U391 (.A1( us10_n447 ) , .A2( us10_n449 ) , .ZN( us10_n805 ) );
  NAND2_X2 us10_U392 (.A1( us10_n449 ) , .A2( us10_n460 ) , .ZN( us10_n792 ) );
  NAND2_X2 us10_U393 (.A1( us10_n441 ) , .A2( us10_n464 ) , .ZN( us10_n708 ) );
  NAND2_X2 us10_U394 (.A2( us10_n471 ) , .A1( us10_n472 ) , .ZN( us10_n817 ) );
  NAND2_X2 us10_U395 (.A2( us10_n460 ) , .A1( us10_n465 ) , .ZN( us10_n780 ) );
  NOR2_X1 us10_U396 (.ZN( us10_n447 ) , .A2( us10_n849 ) , .A1( us10_n858 ) );
  NOR2_X1 us10_U397 (.A2( sa10_6 ) , .A1( sa10_7 ) , .ZN( us10_n464 ) );
  NOR2_X1 us10_U398 (.A2( sa10_7 ) , .ZN( us10_n460 ) , .A1( us10_n849 ) );
  NOR2_X1 us10_U399 (.A2( sa10_4 ) , .ZN( us10_n449 ) , .A1( us10_n848 ) );
  NOR3_X1 us10_U4 (.ZN( us10_n598 ) , .A1( us10_n608 ) , .A3( us10_n723 ) , .A2( us10_n742 ) );
  AOI211_X1 us10_U40 (.B( us10_n694 ) , .A( us10_n695 ) , .ZN( us10_n705 ) , .C2( us10_n831 ) , .C1( us10_n851 ) );
  NOR2_X1 us10_U400 (.A2( sa10_4 ) , .A1( sa10_5 ) , .ZN( us10_n441 ) );
  NOR2_X1 us10_U401 (.A2( sa10_5 ) , .ZN( us10_n448 ) , .A1( us10_n847 ) );
  NOR2_X1 us10_U402 (.A2( sa10_1 ) , .ZN( us10_n471 ) , .A1( us10_n826 ) );
  NOR2_X1 us10_U403 (.A2( sa10_2 ) , .A1( sa10_3 ) , .ZN( us10_n472 ) );
  NOR2_X1 us10_U404 (.A2( sa10_6 ) , .ZN( us10_n452 ) , .A1( us10_n858 ) );
  NOR2_X1 us10_U405 (.A2( sa10_2 ) , .ZN( us10_n461 ) , .A1( us10_n829 ) );
  NOR2_X1 us10_U406 (.A2( sa10_3 ) , .ZN( us10_n455 ) , .A1( us10_n828 ) );
  INV_X1 us10_U407 (.A( sa10_6 ) , .ZN( us10_n849 ) );
  INV_X1 us10_U408 (.A( sa10_4 ) , .ZN( us10_n847 ) );
  INV_X1 us10_U409 (.A( sa10_3 ) , .ZN( us10_n829 ) );
  NOR2_X1 us10_U41 (.ZN( us10_n707 ) , .A2( us10_n776 ) , .A1( us10_n800 ) );
  INV_X1 us10_U410 (.A( sa10_2 ) , .ZN( us10_n828 ) );
  INV_X1 us10_U411 (.A( sa10_7 ) , .ZN( us10_n858 ) );
  INV_X1 us10_U412 (.A( sa10_5 ) , .ZN( us10_n848 ) );
  INV_X1 us10_U413 (.A( sa10_1 ) , .ZN( us10_n827 ) );
  INV_X1 us10_U414 (.A( sa10_0 ) , .ZN( us10_n826 ) );
  NOR2_X1 us10_U415 (.A2( sa10_0 ) , .A1( sa10_1 ) , .ZN( us10_n462 ) );
  NOR2_X1 us10_U416 (.A2( sa10_0 ) , .ZN( us10_n454 ) , .A1( us10_n827 ) );
  OAI222_X1 us10_U417 (.B2( us10_n747 ) , .B1( us10_n748 ) , .A2( us10_n749 ) , .ZN( us10_n757 ) , .C2( us10_n805 ) , .C1( us10_n814 ) , .A1( us10_n817 ) );
  OAI22_X1 us10_U418 (.B2( us10_n803 ) , .B1( us10_n804 ) , .A2( us10_n805 ) , .A1( us10_n806 ) , .ZN( us10_n808 ) );
  OAI21_X1 us10_U419 (.A( us10_n731 ) , .B1( us10_n732 ) , .ZN( us10_n736 ) , .B2( us10_n805 ) );
  NAND4_X1 us10_U42 (.ZN( sa13_sr_7 ) , .A4( us10_n822 ) , .A3( us10_n823 ) , .A2( us10_n824 ) , .A1( us10_n825 ) );
  OAI222_X1 us10_U420 (.ZN( us10_n505 ) , .C2( us10_n625 ) , .B2( us10_n647 ) , .B1( us10_n747 ) , .A2( us10_n748 ) , .C1( us10_n805 ) , .A1( us10_n806 ) );
  AOI21_X1 us10_U421 (.ZN( us10_n650 ) , .A( us10_n779 ) , .B1( us10_n792 ) , .B2( us10_n805 ) );
  INV_X1 us10_U422 (.A( us10_n805 ) , .ZN( us10_n860 ) );
  NOR2_X1 us10_U423 (.ZN( us10_n735 ) , .A2( us10_n803 ) , .A1( us10_n805 ) );
  NOR2_X1 us10_U424 (.ZN( us10_n484 ) , .A1( us10_n788 ) , .A2( us10_n805 ) );
  NOR2_X1 us10_U425 (.A2( us10_n744 ) , .ZN( us10_n755 ) , .A1( us10_n805 ) );
  NAND2_X1 us10_U426 (.ZN( us10_n753 ) , .A1( us10_n763 ) , .A2( us10_n805 ) );
  NOR2_X1 us10_U427 (.ZN( us10_n715 ) , .A1( us10_n805 ) , .A2( us10_n817 ) );
  NOR2_X1 us10_U428 (.ZN( us10_n567 ) , .A1( us10_n747 ) , .A2( us10_n805 ) );
  AOI21_X1 us10_U429 (.ZN( us10_n552 ) , .B1( us10_n669 ) , .A( us10_n697 ) , .B2( us10_n805 ) );
  NOR4_X1 us10_U43 (.A4( us10_n818 ) , .A3( us10_n819 ) , .A2( us10_n820 ) , .A1( us10_n821 ) , .ZN( us10_n822 ) );
  NOR2_X1 us10_U430 (.ZN( us10_n556 ) , .A1( us10_n762 ) , .A2( us10_n805 ) );
  NOR2_X1 us10_U431 (.ZN( us10_n670 ) , .A1( us10_n790 ) , .A2( us10_n805 ) );
  AND2_X1 us10_U432 (.ZN( us10_n438 ) , .A2( us10_n831 ) , .A1( us10_n854 ) );
  AND2_X1 us10_U433 (.ZN( us10_n439 ) , .A2( us10_n843 ) , .A1( us10_n861 ) );
  NOR3_X1 us10_U434 (.A1( us10_n438 ) , .A2( us10_n439 ) , .A3( us10_n576 ) , .ZN( us10_n587 ) );
  NAND4_X1 us10_U435 (.ZN( sa13_sr_2 ) , .A4( us10_n643 ) , .A3( us10_n644 ) , .A2( us10_n645 ) , .A1( us10_n646 ) );
  INV_X1 us10_U436 (.A( us10_n812 ) , .ZN( us10_n854 ) );
  NAND3_X1 us10_U437 (.ZN( sa13_sr_6 ) , .A3( us10_n797 ) , .A2( us10_n798 ) , .A1( us10_n799 ) );
  NAND3_X1 us10_U438 (.ZN( sa13_sr_5 ) , .A3( us10_n758 ) , .A2( us10_n759 ) , .A1( us10_n760 ) );
  NAND3_X1 us10_U439 (.ZN( sa13_sr_4 ) , .A3( us10_n738 ) , .A2( us10_n739 ) , .A1( us10_n740 ) );
  AOI222_X1 us10_U44 (.C2( us10_n809 ) , .B2( us10_n810 ) , .A2( us10_n811 ) , .ZN( us10_n823 ) , .C1( us10_n832 ) , .A1( us10_n839 ) , .B1( us10_n853 ) );
  NAND3_X1 us10_U440 (.A3( us10_n675 ) , .A2( us10_n676 ) , .A1( us10_n677 ) , .ZN( us10_n807 ) );
  NAND3_X1 us10_U441 (.ZN( us10_n638 ) , .A3( us10_n708 ) , .A2( us10_n724 ) , .A1( us10_n792 ) );
  NAND3_X1 us10_U442 (.A3( us10_n618 ) , .A2( us10_n619 ) , .A1( us10_n620 ) , .ZN( us10_n725 ) );
  NAND3_X1 us10_U443 (.A3( us10_n585 ) , .A2( us10_n586 ) , .A1( us10_n587 ) , .ZN( us10_n621 ) );
  NAND3_X1 us10_U444 (.ZN( us10_n565 ) , .A3( us10_n680 ) , .A2( us10_n750 ) , .A1( us10_n785 ) );
  NAND3_X1 us10_U445 (.A3( us10_n523 ) , .A2( us10_n524 ) , .A1( us10_n525 ) , .ZN( us10_n742 ) );
  NAND3_X1 us10_U446 (.A3( us10_n512 ) , .A1( us10_n513 ) , .ZN( us10_n608 ) , .A2( us10_n871 ) );
  NAND3_X1 us10_U447 (.A3( us10_n467 ) , .A2( us10_n468 ) , .A1( us10_n469 ) , .ZN( us10_n777 ) );
  INV_X1 us10_U448 (.A( us10_n803 ) , .ZN( us10_n843 ) );
  AOI21_X1 us10_U449 (.ZN( us10_n576 ) , .B2( us10_n724 ) , .B1( us10_n748 ) , .A( us10_n785 ) );
  AOI211_X1 us10_U45 (.B( us10_n807 ) , .A( us10_n808 ) , .ZN( us10_n824 ) , .C1( us10_n842 ) , .C2( us10_n850 ) );
  NOR4_X1 us10_U46 (.A4( us10_n498 ) , .A3( us10_n499 ) , .A2( us10_n500 ) , .ZN( us10_n501 ) , .A1( us10_n527 ) );
  AOI221_X1 us10_U47 (.A( us10_n497 ) , .ZN( us10_n502 ) , .B2( us10_n843 ) , .C1( us10_n846 ) , .C2( us10_n860 ) , .B1( us10_n862 ) );
  AOI211_X1 us10_U48 (.A( us10_n496 ) , .ZN( us10_n503 ) , .B( us10_n802 ) , .C2( us10_n839 ) , .C1( us10_n851 ) );
  NAND4_X1 us10_U49 (.ZN( sa13_sr_1 ) , .A4( us10_n595 ) , .A3( us10_n596 ) , .A2( us10_n597 ) , .A1( us10_n598 ) );
  NOR3_X1 us10_U5 (.A3( us10_n800 ) , .A2( us10_n801 ) , .A1( us10_n802 ) , .ZN( us10_n825 ) );
  NOR4_X1 us10_U50 (.A4( us10_n591 ) , .A3( us10_n592 ) , .A2( us10_n593 ) , .A1( us10_n594 ) , .ZN( us10_n595 ) );
  AOI211_X1 us10_U51 (.B( us10_n589 ) , .A( us10_n590 ) , .ZN( us10_n596 ) , .C2( us10_n811 ) , .C1( us10_n833 ) );
  AOI211_X1 us10_U52 (.A( us10_n588 ) , .ZN( us10_n597 ) , .B( us10_n621 ) , .C1( us10_n845 ) , .C2( us10_n855 ) );
  NOR2_X1 us10_U53 (.ZN( us10_n804 ) , .A1( us10_n854 ) , .A2( us10_n861 ) );
  NOR2_X1 us10_U54 (.ZN( us10_n625 ) , .A2( us10_n836 ) , .A1( us10_n839 ) );
  AOI222_X1 us10_U55 (.ZN( us10_n469 ) , .B1( us10_n832 ) , .A1( us10_n839 ) , .C1( us10_n842 ) , .C2( us10_n851 ) , .A2( us10_n855 ) , .B2( us10_n865 ) );
  NOR4_X1 us10_U56 (.A1( us10_n466 ) , .ZN( us10_n467 ) , .A4( us10_n542 ) , .A2( us10_n554 ) , .A3( us10_n614 ) );
  AOI221_X1 us10_U57 (.ZN( us10_n468 ) , .C2( us10_n714 ) , .B2( us10_n831 ) , .C1( us10_n845 ) , .B1( us10_n860 ) , .A( us10_n864 ) );
  NAND4_X1 us10_U58 (.A4( us10_n603 ) , .A3( us10_n604 ) , .A2( us10_n605 ) , .A1( us10_n606 ) , .ZN( us10_n722 ) );
  NOR3_X1 us10_U59 (.A1( us10_n599 ) , .ZN( us10_n604 ) , .A3( us10_n663 ) , .A2( us10_n770 ) );
  NOR3_X1 us10_U6 (.ZN( us10_n504 ) , .A2( us10_n679 ) , .A3( us10_n777 ) , .A1( us10_n876 ) );
  NOR4_X1 us10_U60 (.A3( us10_n600 ) , .A2( us10_n601 ) , .A1( us10_n602 ) , .ZN( us10_n603 ) , .A4( us10_n655 ) );
  AOI222_X1 us10_U61 (.ZN( us10_n606 ) , .A1( us10_n830 ) , .C2( us10_n837 ) , .B1( us10_n842 ) , .A2( us10_n856 ) , .B2( us10_n861 ) , .C1( us10_n868 ) );
  AOI222_X1 us10_U62 (.B2( us10_n638 ) , .ZN( us10_n644 ) , .B1( us10_n841 ) , .A1( us10_n842 ) , .C2( us10_n846 ) , .C1( us10_n863 ) , .A2( us10_n865 ) );
  NOR4_X1 us10_U63 (.A4( us10_n639 ) , .A3( us10_n640 ) , .A2( us10_n641 ) , .A1( us10_n642 ) , .ZN( us10_n643 ) );
  NOR3_X1 us10_U64 (.A2( us10_n607 ) , .A1( us10_n608 ) , .ZN( us10_n646 ) , .A3( us10_n722 ) );
  NAND4_X1 us10_U65 (.A4( us10_n657 ) , .A3( us10_n658 ) , .A2( us10_n659 ) , .A1( us10_n660 ) , .ZN( us10_n800 ) );
  NOR3_X1 us10_U66 (.A3( us10_n648 ) , .A2( us10_n649 ) , .A1( us10_n650 ) , .ZN( us10_n659 ) );
  NOR3_X1 us10_U67 (.A3( us10_n651 ) , .A2( us10_n652 ) , .A1( us10_n653 ) , .ZN( us10_n658 ) );
  NOR3_X1 us10_U68 (.A3( us10_n654 ) , .A2( us10_n655 ) , .A1( us10_n656 ) , .ZN( us10_n657 ) );
  NAND4_X1 us10_U69 (.A4( us10_n560 ) , .A3( us10_n561 ) , .A2( us10_n562 ) , .A1( us10_n563 ) , .ZN( us10_n607 ) );
  INV_X1 us10_U7 (.A( us10_n706 ) , .ZN( us10_n876 ) );
  NOR4_X1 us10_U70 (.A4( us10_n552 ) , .A3( us10_n553 ) , .A2( us10_n554 ) , .A1( us10_n555 ) , .ZN( us10_n562 ) );
  NOR4_X1 us10_U71 (.A4( us10_n556 ) , .A3( us10_n557 ) , .A2( us10_n558 ) , .A1( us10_n559 ) , .ZN( us10_n560 ) );
  NOR4_X1 us10_U72 (.ZN( us10_n561 ) , .A1( us10_n653 ) , .A3( us10_n661 ) , .A4( us10_n685 ) , .A2( us10_n768 ) );
  NAND4_X1 us10_U73 (.A4( us10_n772 ) , .A3( us10_n773 ) , .A2( us10_n774 ) , .A1( us10_n775 ) , .ZN( us10_n801 ) );
  NOR3_X1 us10_U74 (.A3( us10_n765 ) , .A2( us10_n766 ) , .A1( us10_n767 ) , .ZN( us10_n773 ) );
  NOR4_X1 us10_U75 (.A4( us10_n768 ) , .A3( us10_n769 ) , .A2( us10_n770 ) , .A1( us10_n771 ) , .ZN( us10_n772 ) );
  AOI222_X1 us10_U76 (.ZN( us10_n775 ) , .A1( us10_n830 ) , .C1( us10_n834 ) , .B2( us10_n841 ) , .A2( us10_n850 ) , .B1( us10_n861 ) , .C2( us10_n873 ) );
  NOR4_X1 us10_U77 (.A4( us10_n665 ) , .A3( us10_n666 ) , .A2( us10_n667 ) , .A1( us10_n668 ) , .ZN( us10_n676 ) );
  NOR4_X1 us10_U78 (.A4( us10_n661 ) , .A3( us10_n662 ) , .A2( us10_n663 ) , .A1( us10_n664 ) , .ZN( us10_n677 ) );
  NOR4_X1 us10_U79 (.A3( us10_n673 ) , .A1( us10_n674 ) , .ZN( us10_n675 ) , .A4( us10_n715 ) , .A2( us10_n859 ) );
  NOR3_X1 us10_U8 (.A3( us10_n621 ) , .A2( us10_n622 ) , .ZN( us10_n636 ) , .A1( us10_n725 ) );
  NOR2_X1 us10_U80 (.ZN( us10_n761 ) , .A1( us10_n833 ) , .A2( us10_n834 ) );
  NOR4_X1 us10_U81 (.A4( us10_n577 ) , .A3( us10_n578 ) , .A2( us10_n579 ) , .ZN( us10_n586 ) , .A1( us10_n683 ) );
  NOR4_X1 us10_U82 (.A1( us10_n584 ) , .ZN( us10_n585 ) , .A3( us10_n652 ) , .A2( us10_n662 ) , .A4( us10_n767 ) );
  AOI222_X1 us10_U83 (.ZN( us10_n513 ) , .C1( us10_n832 ) , .B2( us10_n837 ) , .A2( us10_n843 ) , .C2( us10_n862 ) , .B1( us10_n863 ) , .A1( us10_n866 ) );
  NOR4_X1 us10_U84 (.A4( us10_n509 ) , .A2( us10_n510 ) , .A1( us10_n511 ) , .ZN( us10_n512 ) , .A3( us10_n670 ) );
  INV_X1 us10_U85 (.A( us10_n505 ) , .ZN( us10_n871 ) );
  NAND4_X1 us10_U86 (.A4( us10_n456 ) , .A3( us10_n457 ) , .A2( us10_n458 ) , .A1( us10_n459 ) , .ZN( us10_n679 ) );
  NOR3_X1 us10_U87 (.ZN( us10_n457 ) , .A3( us10_n530 ) , .A1( us10_n555 ) , .A2( us10_n570 ) );
  NOR4_X1 us10_U88 (.ZN( us10_n458 ) , .A2( us10_n509 ) , .A1( us10_n599 ) , .A4( us10_n628 ) , .A3( us10_n711 ) );
  NOR4_X1 us10_U89 (.ZN( us10_n456 ) , .A2( us10_n517 ) , .A1( us10_n543 ) , .A3( us10_n579 ) , .A4( us10_n615 ) );
  NOR2_X1 us10_U9 (.ZN( us10_n575 ) , .A1( us10_n622 ) , .A2( us10_n745 ) );
  NAND4_X1 us10_U90 (.A4( us10_n535 ) , .A3( us10_n536 ) , .A2( us10_n537 ) , .A1( us10_n538 ) , .ZN( us10_n622 ) );
  NOR4_X1 us10_U91 (.A4( us10_n526 ) , .A2( us10_n527 ) , .A1( us10_n528 ) , .ZN( us10_n538 ) , .A3( us10_n701 ) );
  NOR4_X1 us10_U92 (.A1( us10_n531 ) , .ZN( us10_n536 ) , .A2( us10_n654 ) , .A4( us10_n668 ) , .A3( us10_n765 ) );
  NOR4_X1 us10_U93 (.A4( us10_n529 ) , .A3( us10_n530 ) , .ZN( us10_n537 ) , .A2( us10_n684 ) , .A1( us10_n794 ) );
  NOR2_X1 us10_U94 (.ZN( us10_n686 ) , .A1( us10_n831 ) , .A2( us10_n832 ) );
  NAND4_X1 us10_U95 (.A4( us10_n479 ) , .A3( us10_n480 ) , .A2( us10_n481 ) , .A1( us10_n482 ) , .ZN( us10_n694 ) );
  NOR3_X1 us10_U96 (.ZN( us10_n480 ) , .A2( us10_n508 ) , .A3( us10_n601 ) , .A1( us10_n610 ) );
  AOI211_X1 us10_U97 (.B( us10_n477 ) , .A( us10_n478 ) , .ZN( us10_n482 ) , .C2( us10_n833 ) , .C1( us10_n861 ) );
  NOR4_X1 us10_U98 (.ZN( us10_n481 ) , .A3( us10_n532 ) , .A4( us10_n545 ) , .A2( us10_n567 ) , .A1( us10_n717 ) );
  NAND4_X1 us10_U99 (.A4( us10_n548 ) , .A3( us10_n549 ) , .A2( us10_n550 ) , .A1( us10_n551 ) , .ZN( us10_n745 ) );
endmodule

