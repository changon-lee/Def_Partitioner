module aes_aes ( clk, key, ld, rst, text_in, done, text_out );
  input clk;
  input [127:0] key;
  input ld;
  input rst;
  input [127:0] text_in;
  output done;
  output [127:0] text_out;

  wire N100, N101, N102, N103, N104, N105, N114, N115, 
       N116, N117, N118, N119, N120, N121, N130, N131, N132, 
       N133, N134, N135, N136, N137, N146, N147, N148, N149, 
       N150, N151, N152, N153, N162, N163, N164, N165, N166, 
       N167, N168, N169, N178, N179, N180, N181, N182, N183, 
       N184, N185, N194, N195, N196, N197, N198, N199, N200, 
       N201, N210, N211, N212, N213, N214, N215, N216, N217, 
       N226, N227, N228, N229, N230, N231, N232, N233, N242, 
       N243, N244, N245, N246, N247, N248, N249, N258, N259, 
       N260, N261, N262, N263, N264, N265, N274, N275, N276, 
       N277, N278, N279, N280, N281, N34, N35, N36, N37, 
       N378, N379, N38, N382, N383, N384, N385, N39, N392, 
       N393, N394, N395, N398, N399, N40, N41, N415, N419, 
       N423, N441, N454, N455, N456, N457, N458, N459, N460, 
       N461, N463, N466, N467, N468, N469, N470, N471, N472, 
       N473, N474, N475, N476, N477, N478, N479, N480, N481, 
       N482, N483, N484, N485, N486, N487, N488, N489, N490, 
       N491, N492, N493, N494, N495, N496, N497, N498, N499, 
       N50, N500, N501, N502, N503, N504, N505, N51, N52, 
       N53, N54, N55, N56, N57, N66, N67, N68, N69, 
       N70, N71, N72, N73, N82, N83, N84, N85, N86, 
       N87, N88, N89, N98, N99, n1, n101, n103, n105, 
       n107, n109, n11, n1109, n111, n1114, n113, n115, n117, 
       n119, n121, n123, n125, n127, n129, n13, n131, n133, 
       n135, n137, n139, n141, n143, n145, n147, n149, n15, 
       n151, n153, n155, n157, n159, n161, n163, n165, n167, 
       n169, n17, n171, n173, n175, n177, n179, n181, n183, 
       n185, n187, n189, n19, n191, n193, n195, n197, n199, 
       n201, n203, n205, n207, n209, n21, n211, n213, n215, 
       n217, n219, n221, n223, n225, n227, n229, n23, n231, 
       n233, n235, n237, n239, n241, n243, n245, n247, n249, 
       n25, n251, n253, n255, n27, n29, n3, n31, n33, 
       n35, n37, n39, n41, n43, n45, n47, n49, n5, 
       n51, n53, n55, n57, n59, n61, n63, n65, n67, 
       n69, n7, n71, n73, n75, n77, n79, n81, n83, 
       n85, n87, n89, n9, n91, n93, n95, n97, n99, 
       sa00_0, sa00_1, sa00_2, sa00_3, sa00_4, sa00_5, sa00_6, sa00_7, sa00_sr_0, 
       sa00_sr_1, sa00_sr_2, sa00_sr_3, sa00_sr_4, sa00_sr_5, sa00_sr_6, sa00_sr_7, sa01_0, sa01_1, 
       sa01_2, sa01_3, sa01_4, sa01_5, sa01_6, sa01_7, sa01_sr_0, sa01_sr_1, sa01_sr_2, 
       sa01_sr_3, sa01_sr_4, sa01_sr_5, sa01_sr_6, sa01_sr_7, sa02_0, sa02_1, sa02_2, sa02_3, 
       sa02_4, sa02_5, sa02_6, sa02_7, sa02_sr_0, sa02_sr_1, sa02_sr_2, sa02_sr_3, sa02_sr_4, 
       sa02_sr_5, sa02_sr_6, sa02_sr_7, sa03_0, sa03_1, sa03_2, sa03_3, sa03_4, sa03_5, 
       sa03_6, sa03_7, sa03_sr_0, sa03_sr_1, sa03_sr_2, sa03_sr_3, sa03_sr_4, sa03_sr_5, sa03_sr_6, 
       sa03_sr_7, sa10_0, sa10_1, sa10_2, sa10_3, sa10_4, sa10_5, sa10_6, sa10_7, 
       sa10_sr_0, sa10_sr_1, sa10_sr_2, sa10_sr_3, sa10_sr_4, sa10_sr_5, sa10_sr_6, sa10_sr_7, sa11_0, 
       sa11_1, sa11_2, sa11_3, sa11_4, sa11_5, sa11_6, sa11_7, sa11_sr_0, sa11_sr_1, 
       sa11_sr_2, sa11_sr_3, sa11_sr_4, sa11_sr_5, sa11_sr_6, sa11_sr_7, sa12_0, sa12_1, sa12_2, 
       sa12_3, sa12_4, sa12_5, sa12_6, sa12_7, sa12_sr_0, sa12_sr_1, sa12_sr_2, sa12_sr_3, 
       sa12_sr_4, sa12_sr_5, sa12_sr_6, sa12_sr_7, sa13_0, sa13_1, sa13_2, sa13_3, sa13_4, 
       sa13_5, sa13_6, sa13_7, sa13_sr_0, sa13_sr_1, sa13_sr_2, sa13_sr_3, sa13_sr_4, sa13_sr_5, 
       sa13_sr_6, sa13_sr_7, sa20_0, sa20_1, sa20_2, sa20_3, sa20_4, sa20_5, sa20_6, 
       sa20_7, sa20_sr_0, sa20_sr_1, sa20_sr_2, sa20_sr_3, sa20_sr_4, sa20_sr_5, sa20_sr_6, sa20_sr_7, 
       sa21_0, sa21_1, sa21_2, sa21_3, sa21_4, sa21_5, sa21_6, sa21_7, sa21_sr_0, 
       sa21_sr_1, sa21_sr_2, sa21_sr_3, sa21_sr_4, sa21_sr_5, sa21_sr_6, sa21_sr_7, sa22_0, sa22_1, 
       sa22_2, sa22_3, sa22_4, sa22_5, sa22_6, sa22_7, sa22_sr_0, sa22_sr_1, sa22_sr_2, 
       sa22_sr_3, sa22_sr_4, sa22_sr_5, sa22_sr_6, sa22_sr_7, sa23_0, sa23_1, sa23_2, sa23_3, 
       sa23_4, sa23_5, sa23_6, sa23_7, sa23_sr_0, sa23_sr_1, sa23_sr_2, sa23_sr_3, sa23_sr_4, 
       sa23_sr_5, sa23_sr_6, sa23_sr_7, sa30_0, sa30_1, sa30_2, sa30_3, sa30_4, sa30_5, 
       sa30_6, sa30_7, sa30_sr_0, sa30_sr_1, sa30_sr_2, sa30_sr_3, sa30_sr_4, sa30_sr_5, sa30_sr_6, 
       sa30_sr_7, sa31_0, sa31_1, sa31_2, sa31_3, sa31_4, sa31_5, sa31_6, sa31_7, 
       sa31_sr_0, sa31_sr_1, sa31_sr_2, sa31_sr_3, sa31_sr_4, sa31_sr_5, sa31_sr_6, sa31_sr_7, sa32_0, 
       sa32_1, sa32_2, sa32_3, sa32_4, sa32_5, sa32_6, sa32_7, sa32_sr_0, sa32_sr_1, 
       sa32_sr_2, sa32_sr_3, sa32_sr_4, sa32_sr_5, sa32_sr_6, sa32_sr_7, sa33_0, sa33_1, sa33_2, 
       sa33_3, sa33_4, sa33_5, sa33_6, sa33_7, sa33_sr_0, sa33_sr_1, sa33_sr_2, sa33_sr_3, 
       sa33_sr_4, sa33_sr_5, sa33_sr_6, sa33_sr_7, u0_n104, u0_n106, u0_n107, u0_n109, u0_n113, 
       u0_n115, u0_n116, u0_n118, u0_n119, u0_n121, u0_n122, u0_n124, u0_n128, u0_n130, 
       u0_n134, u0_n136, u0_n137, u0_n139, u0_n15, u0_n152, u0_n154, u0_n158, u0_n160, 
       u0_n176, u0_n188, u0_n190, u0_n194, u0_n196, u0_n198, u0_n200, u0_n204, u0_n208, 
       u0_n210, u0_n220, u0_n224, u0_n250, u0_n254, u0_n258, u0_n264, u0_n268, u0_n27, 
       u0_n270, u0_n272, u0_n274, u0_n29, u0_n33, u0_n35, u0_n37, u0_n39, u0_n43, 
       u0_n47, u0_n49, u0_n59, u0_n63, u0_n88, u0_r0_N70, u0_r0_N71, u0_r0_N72, u0_r0_N73, 
       u0_r0_N74, u0_r0_N75, u0_r0_N76, u0_r0_N77, u0_r0_N78, u0_r0_N79, u0_r0_N80, u0_r0_N81, u0_r0_n12, 
       u0_r0_n18, u0_r0_n3, u0_r0_n6, u0_r0_n8, u0_r0_n9, u0_r0_rcnt_0, u0_r0_rcnt_1, u0_r0_rcnt_2, u0_rcon_24, 
       u0_subword_1, u0_subword_11, u0_subword_16, u0_subword_19, u0_subword_20, u0_subword_21, u0_subword_22, u0_subword_23, u0_subword_25, 
       u0_subword_26, u0_subword_27, u0_subword_28, u0_subword_29, u0_subword_3, u0_subword_30, u0_subword_31, u0_subword_4, u0_subword_5, 
       u0_subword_6, u0_subword_9, w0_0, w0_1, w0_10, w0_11, w0_12, w0_13, w0_14, 
       w0_15, w0_16, w0_17, w0_18, w0_19, w0_2, w0_20, w0_21, w0_22, 
       w0_23, w0_24, w0_25, w0_26, w0_27, w0_28, w0_29, w0_3, w0_30, 
       w0_31, w0_4, w0_5, w0_6, w0_7, w0_8, w0_9, w1_0, w1_1, 
       w1_10, w1_11, w1_12, w1_13, w1_14, w1_15, w1_16, w1_17, w1_18, 
       w1_19, w1_2, w1_20, w1_21, w1_22, w1_23, w1_24, w1_25, w1_26, 
       w1_27, w1_28, w1_29, w1_3, w1_30, w1_31, w1_4, w1_5, w1_6, 
       w1_7, w1_8, w1_9, w2_0, w2_1, w2_10, w2_11, w2_12, w2_13, 
       w2_14, w2_15, w2_16, w2_17, w2_18, w2_19, w2_2, w2_20, w2_21, 
       w2_22, w2_23, w2_24, w2_25, w2_26, w2_27, w2_28, w2_29, w2_3, 
       w2_30, w2_31, w2_4, w2_5, w2_6, w2_7, w2_8, w2_9, w3_0, 
       w3_1, w3_10, w3_11, w3_16, w3_17, w3_18, w3_19, w3_2, w3_20, 
       w3_21, w3_22, w3_23, w3_24, w3_25, w3_26, w3_27, w3_28, w3_29, 
       w3_3, w3_30, w3_31, w3_4, w3_5, w3_6, w3_7, w3_8, w3_9 ;

  aes_aes_die_0 u0 ( clk, key, ld, rst, text_in, done, text_out, N100, N101, N102, N103, N104, N105, N114, N115, 
      N116, N117, N118, N119, N120, N121, N130, N131, N132, 
      N133, N134, N135, N136, N137, N146, N147, N148, N149, 
      N150, N151, N152, N153, N162, N163, N164, N165, N166, 
      N167, N168, N169, N178, N179, N180, N181, N182, N183, 
      N184, N185, N194, N195, N196, N197, N198, N199, N200, 
      N201, N210, N211, N212, N213, N214, N215, N216, N217, 
      N226, N227, N228, N229, N230, N231, N232, N233, N242, 
      N243, N244, N245, N246, N247, N248, N249, N258, N259, 
      N260, N261, N262, N263, N264, N265, N274, N275, N276, 
      N277, N278, N279, N280, N281, N34, N35, N36, N37, 
      N378, N379, N38, N382, N383, N384, N385, N39, N392, 
      N393, N394, N395, N398, N399, N40, N41, N415, N419, 
      N423, N441, N454, N455, N456, N457, N458, N459, N460, 
      N461, N463, N466, N467, N468, N469, N470, N471, N472, 
      N473, N474, N475, N476, N477, N478, N479, N480, N481, 
      N482, N483, N484, N485, N486, N487, N488, N489, N490, 
      N491, N492, N493, N494, N495, N496, N497, N498, N499, 
      N50, N500, N501, N502, N503, N504, N505, N51, N52, 
      N53, N54, N55, N56, N57, N66, N67, N68, N69, 
      N70, N71, N72, N73, N82, N83, N84, N85, N86, 
      N87, N88, N89, N98, N99, sa00_sr_4, sa00_sr_5, sa01_sr_2, sa01_sr_3, 
      sa01_sr_4, sa01_sr_5, sa01_sr_6, sa01_sr_7, sa02_sr_0, sa02_sr_1, sa02_sr_4, sa02_sr_5, sa03_sr_0, 
      sa03_sr_1, sa03_sr_2, sa03_sr_3, sa03_sr_4, sa03_sr_5, sa03_sr_6, sa03_sr_7, sa10_sr_0, sa10_sr_1, 
      sa10_sr_3, sa10_sr_4, sa10_sr_5, sa10_sr_6, sa10_sr_7, sa11_sr_0, sa11_sr_1, sa11_sr_3, sa11_sr_4, 
      sa11_sr_5, sa11_sr_7, sa12_sr_0, sa12_sr_1, sa12_sr_2, sa12_sr_3, sa12_sr_4, sa12_sr_5, sa12_sr_6, 
      sa12_sr_7, sa13_sr_1, sa13_sr_2, sa13_sr_3, sa13_sr_4, sa13_sr_5, sa13_sr_6, sa13_sr_7, sa20_sr_0, 
      sa20_sr_1, sa20_sr_2, sa20_sr_3, sa20_sr_4, sa20_sr_5, sa20_sr_6, sa20_sr_7, sa21_sr_4, sa21_sr_5, 
      sa21_sr_6, sa21_sr_7, sa22_sr_0, sa22_sr_1, sa22_sr_3, u0_n104, u0_n106, u0_n107, u0_n109, 
      u0_n113, u0_n115, u0_n116, u0_n118, u0_n119, u0_n121, u0_n122, u0_n124, u0_n128, 
      u0_n130, u0_n134, u0_n136, u0_n137, u0_n139, u0_n15, u0_n152, u0_n154, u0_n158, 
      u0_n160, u0_n176, u0_n188, u0_n190, u0_n194, u0_n196, u0_n198, u0_n200, u0_n204, 
      u0_n208, u0_n210, u0_n220, u0_n224, u0_n27, u0_n29, u0_n33, u0_n35, u0_n37, 
      u0_n39, u0_n43, u0_n47, u0_n49, u0_n59, u0_n63, u0_n88, u0_r0_N70, u0_r0_N71, 
      u0_r0_N72, u0_r0_N73, u0_r0_N74, u0_r0_N75, u0_r0_N76, u0_r0_N77, u0_r0_N81, u0_r0_n12, u0_r0_n18, 
      u0_subword_1, u0_subword_11, u0_subword_16, u0_subword_19, u0_subword_20, u0_subword_21, u0_subword_22, u0_subword_23, u0_subword_25, 
      u0_subword_26, u0_subword_27, u0_subword_28, u0_subword_29, u0_subword_3, u0_subword_30, u0_subword_31, u0_subword_4, u0_subword_5, 
      u0_subword_6, u0_subword_9, n1, n101, n103, n105, n107, n109, n11, 
      n1109, n111, n1114, n113, n115, n117, n119, n121, n123, 
      n125, n127, n129, n13, n131, n133, n135, n137, n139, 
      n141, n143, n145, n147, n149, n15, n151, n153, n155, 
      n157, n159, n161, n163, n165, n167, n169, n17, n171, 
      n173, n175, n177, n179, n181, n183, n185, n187, n189, 
      n19, n191, n193, n195, n197, n199, n201, n203, n205, 
      n207, n209, n21, n211, n213, n215, n217, n219, n221, 
      n223, n225, n227, n229, n23, n231, n233, n235, n237, 
      n239, n241, n243, n245, n247, n249, n25, n251, n253, 
      n255, n27, n29, n3, n31, n33, n35, n37, n39, 
      n41, n43, n45, n47, n49, n5, n51, n53, n55, 
      n57, n59, n61, n63, n65, n67, n69, n7, n71, 
      n73, n75, n77, n79, n81, n83, n85, n87, n89, 
      n9, n91, n93, n95, n97, n99, sa00_0, sa00_1, sa00_2, 
      sa00_3, sa00_4, sa00_5, sa00_6, sa00_7, sa01_0, sa01_1, sa01_2, sa01_3, 
      sa01_4, sa01_5, sa01_6, sa01_7, sa02_0, sa02_1, sa02_2, sa02_3, sa02_4, 
      sa02_5, sa02_6, sa02_7, sa03_0, sa03_1, sa03_2, sa03_3, sa03_4, sa03_5, 
      sa03_6, sa03_7, sa10_0, sa10_1, sa10_2, sa10_3, sa10_4, sa10_5, sa10_6, 
      sa10_7, sa11_0, sa11_1, sa11_2, sa11_3, sa11_4, sa11_5, sa11_6, sa11_7, 
      sa12_0, sa12_1, sa12_2, sa12_3, sa12_4, sa12_5, sa12_6, sa12_7, sa13_0, 
      sa13_1, sa13_2, sa13_3, sa13_4, sa13_5, sa13_6, sa13_7, sa20_0, sa20_1, 
      sa20_2, sa20_3, sa20_4, sa20_5, sa20_6, sa20_7, sa21_0, sa21_1, sa21_2, 
      sa21_3, sa21_4, sa21_5, sa21_6, sa21_7, sa22_0, sa22_1, sa22_2, sa22_3, 
      sa22_4, sa22_5, sa22_6, sa22_7, sa23_0, sa23_1, sa23_2, sa23_3, sa23_4, 
      sa23_5, sa23_6, sa23_7, sa30_0, sa30_1, sa30_2, sa30_3, sa30_4, sa30_5, 
      sa30_6, sa30_7, sa31_0, sa31_1, sa31_2, sa31_3, sa31_4, sa31_5, sa31_6, 
      sa31_7, sa32_0, sa32_1, sa32_2, sa32_3, sa32_4, sa32_5, sa32_6, sa32_7, 
      sa33_0, sa33_1, sa33_2, sa33_3, sa33_4, sa33_5, sa33_6, sa33_7, u0_n250, 
      u0_n254, u0_n258, u0_n264, u0_n268, u0_n270, u0_n272, u0_n274, u0_r0_N78, u0_r0_N79, 
      u0_r0_N80, u0_r0_n3, u0_r0_n6, u0_r0_n8, u0_r0_n9, u0_r0_rcnt_0, u0_r0_rcnt_1, u0_r0_rcnt_2, u0_rcon_24, 
      w0_0, w0_1, w0_10, w0_11, w0_12, w0_13, w0_14, w0_15, w0_16, 
      w0_17, w0_18, w0_19, w0_2, w0_20, w0_21, w0_22, w0_23, w0_24, 
      w0_25, w0_26, w0_27, w0_28, w0_29, w0_3, w0_30, w0_31, w0_4, 
      w0_5, w0_6, w0_7, w0_8, w0_9, w1_0, w1_1, w1_10, w1_11, 
      w1_12, w1_13, w1_14, w1_15, w1_16, w1_17, w1_18, w1_19, w1_2, 
      w1_20, w1_21, w1_22, w1_23, w1_24, w1_25, w1_26, w1_27, w1_28, 
      w1_29, w1_3, w1_30, w1_31, w1_4, w1_5, w1_6, w1_7, w1_8, 
      w1_9, w2_0, w2_1, w2_10, w2_11, w2_12, w2_13, w2_14, w2_15, 
      w2_16, w2_17, w2_18, w2_19, w2_2, w2_20, w2_21, w2_22, w2_23, 
      w2_24, w2_25, w2_26, w2_27, w2_28, w2_29, w2_3, w2_30, w2_31, 
      w2_4, w2_5, w2_6, w2_7, w2_8, w2_9, w3_0, w3_1, w3_10, 
      w3_11, w3_16, w3_17, w3_18, w3_19, w3_2, w3_20, w3_21, w3_22, 
      w3_23, w3_24, w3_25, w3_26, w3_27, w3_28, w3_29, w3_3, w3_30, 
      w3_31, w3_4, w3_5, w3_6, w3_7, w3_8, w3_9 );
  aes_aes_die_1 u1 ( sa11_0, sa11_1, sa11_2, sa11_3, sa11_4, sa11_5, sa11_6, sa11_7, sa13_0, 
      sa13_1, sa13_2, sa13_3, sa13_4, sa13_5, sa13_6, sa13_7, sa10_sr_0, sa10_sr_1, 
      sa10_sr_2, sa10_sr_3, sa10_sr_4, sa10_sr_5, sa10_sr_6, sa10_sr_7, sa12_sr_0, sa12_sr_1, sa12_sr_2, 
      sa12_sr_3, sa12_sr_4, sa12_sr_5, sa12_sr_6, sa12_sr_7 );
  aes_aes_die_2 u2 ( sa01_0, sa01_1, sa01_2, sa01_3, sa01_4, sa01_5, sa01_6, sa01_7, sa02_0, 
      sa02_1, sa02_2, sa02_3, sa02_4, sa02_5, sa02_6, sa02_7, sa01_sr_0, sa01_sr_1, 
      sa01_sr_2, sa01_sr_3, sa01_sr_4, sa01_sr_5, sa01_sr_6, sa01_sr_7, sa02_sr_0, sa02_sr_1, sa02_sr_2, 
      sa02_sr_3, sa02_sr_4, sa02_sr_5, sa02_sr_6, sa02_sr_7 );
  aes_aes_die_3 u3 ( sa03_0, sa03_1, sa03_2, sa03_3, sa03_4, sa03_5, sa03_6, sa03_7, sa33_0, 
      sa33_1, sa33_2, sa33_3, sa33_4, sa33_5, sa33_6, sa33_7, sa03_sr_0, sa03_sr_1, 
      sa03_sr_2, sa03_sr_3, sa03_sr_4, sa03_sr_5, sa03_sr_6, sa03_sr_7, sa30_sr_0, sa30_sr_1, sa30_sr_2, 
      sa30_sr_3, sa30_sr_4, sa30_sr_5, sa30_sr_6, sa30_sr_7 );
  aes_aes_die_4 u4 ( sa20_0, sa20_1, sa20_2, sa20_3, sa20_4, sa20_5, sa20_6, sa20_7, sa31_0, 
      sa31_1, sa31_2, sa31_3, sa31_4, sa31_5, sa31_6, sa31_7, sa22_sr_0, sa22_sr_1, 
      sa22_sr_2, sa22_sr_3, sa22_sr_4, sa22_sr_5, sa22_sr_6, sa22_sr_7, sa32_sr_0, sa32_sr_1, sa32_sr_2, 
      sa32_sr_3, sa32_sr_4, sa32_sr_5, sa32_sr_6, sa32_sr_7 );
  aes_aes_die_5 u5 ( sa10_0, sa10_1, sa10_2, sa10_3, sa10_4, sa10_5, sa10_6, sa10_7, sa22_0, 
      sa22_1, sa22_2, sa22_3, sa22_4, sa22_5, sa22_6, sa22_7, sa13_sr_0, sa13_sr_1, 
      sa13_sr_2, sa13_sr_3, sa13_sr_4, sa13_sr_5, sa13_sr_6, sa13_sr_7, sa20_sr_0, sa20_sr_1, sa20_sr_2, 
      sa20_sr_3, sa20_sr_4, sa20_sr_5, sa20_sr_6, sa20_sr_7 );
  aes_aes_die_6 u6 ( sa12_0, sa12_1, sa12_2, sa12_3, sa12_4, sa12_5, sa12_6, sa12_7, sa21_0, 
      sa21_1, sa21_2, sa21_3, sa21_4, sa21_5, sa21_6, sa21_7, sa11_sr_0, sa11_sr_1, 
      sa11_sr_2, sa11_sr_3, sa11_sr_4, sa11_sr_5, sa11_sr_6, sa11_sr_7, sa23_sr_0, sa23_sr_1, sa23_sr_2, 
      sa23_sr_3, sa23_sr_4, sa23_sr_5, sa23_sr_6, sa23_sr_7 );
  aes_aes_die_7 u7 ( sa23_0, sa23_1, sa23_2, sa23_3, sa23_4, sa23_5, sa23_6, sa23_7, u0_rcon_24, 
      w0_24, w3_16, w3_17, w3_18, w3_19, w3_20, w3_21, w3_22, w3_23, 
      sa21_sr_0, sa21_sr_1, sa21_sr_2, sa21_sr_3, sa21_sr_4, sa21_sr_5, sa21_sr_6, sa21_sr_7, u0_n15, 
      u0_subword_25, u0_subword_26, u0_subword_27, u0_subword_28, u0_subword_29, u0_subword_30, u0_subword_31 );
  aes_aes_die_8 u8 ( n1, n101, n103, n105, n107, n109, n11, n1109, n111, 
      n1114, n113, n115, n117, n119, n121, n123, n125, n127, 
      n129, n13, n131, n133, n135, n137, n139, n141, n143, 
      n145, n147, n149, n15, n151, n153, n155, n157, n159, 
      n161, n163, n165, n167, n169, n17, n171, n173, n175, 
      n177, n179, n181, n183, n185, n187, n189, n19, n191, 
      n193, n195, n197, n199, n201, n203, n205, n207, n209, 
      n21, n211, n213, n215, n217, n219, n221, n223, n225, 
      n227, n229, n23, n231, n233, n235, n237, n239, n241, 
      n243, n245, n247, n249, n25, n251, n253, n255, n27, 
      n29, n3, n31, n33, n35, n37, n39, n41, n43, 
      n45, n47, n49, n5, n51, n53, n55, n57, n59, 
      n61, n63, n65, n67, n69, n7, n71, n73, n75, 
      n77, n79, n81, n83, n85, n87, n89, n9, n91, 
      n93, n95, n97, n99, sa00_sr_0, sa00_sr_1, sa00_sr_2, sa00_sr_3, sa00_sr_4, 
      sa00_sr_5, sa00_sr_6, sa00_sr_7, sa01_sr_0, sa01_sr_1, sa01_sr_2, sa01_sr_3, sa01_sr_4, sa01_sr_5, 
      sa01_sr_6, sa01_sr_7, sa02_sr_0, sa02_sr_1, sa02_sr_2, sa02_sr_3, sa02_sr_4, sa02_sr_5, sa02_sr_6, 
      sa02_sr_7, sa03_sr_0, sa03_sr_1, sa03_sr_2, sa03_sr_3, sa03_sr_4, sa03_sr_5, sa03_sr_6, sa03_sr_7, 
      sa10_sr_0, sa10_sr_1, sa10_sr_2, sa10_sr_3, sa10_sr_4, sa10_sr_5, sa10_sr_6, sa10_sr_7, sa11_sr_0, 
      sa11_sr_1, sa11_sr_2, sa11_sr_3, sa11_sr_4, sa11_sr_5, sa11_sr_6, sa11_sr_7, sa12_sr_0, sa12_sr_1, 
      sa12_sr_2, sa12_sr_3, sa12_sr_4, sa12_sr_5, sa12_sr_6, sa12_sr_7, sa13_sr_0, sa13_sr_1, sa13_sr_2, 
      sa13_sr_3, sa13_sr_4, sa13_sr_5, sa13_sr_6, sa13_sr_7, sa20_sr_0, sa20_sr_1, sa20_sr_2, sa20_sr_3, 
      sa20_sr_4, sa20_sr_5, sa20_sr_6, sa20_sr_7, sa21_sr_0, sa21_sr_1, sa21_sr_2, sa21_sr_3, sa21_sr_4, 
      sa21_sr_5, sa21_sr_6, sa21_sr_7, sa22_sr_0, sa22_sr_1, sa22_sr_2, sa22_sr_3, sa22_sr_4, sa22_sr_5, 
      sa22_sr_6, sa22_sr_7, sa23_sr_0, sa23_sr_1, sa23_sr_2, sa23_sr_3, sa23_sr_4, sa23_sr_5, sa23_sr_6, 
      sa23_sr_7, sa30_sr_0, sa30_sr_1, sa30_sr_2, sa30_sr_3, sa30_sr_4, sa30_sr_5, sa30_sr_6, sa30_sr_7, 
      sa31_sr_0, sa31_sr_1, sa31_sr_2, sa31_sr_3, sa31_sr_4, sa31_sr_5, sa31_sr_6, sa31_sr_7, sa32_sr_0, 
      sa32_sr_1, sa32_sr_2, sa32_sr_3, sa32_sr_4, sa32_sr_5, sa32_sr_6, sa32_sr_7, sa33_sr_0, sa33_sr_1, 
      sa33_sr_2, sa33_sr_3, sa33_sr_4, sa33_sr_5, sa33_sr_6, sa33_sr_7, u0_n15, u0_n250, u0_n254, 
      u0_n258, u0_n264, u0_n27, u0_n29, u0_n33, u0_n35, u0_n37, u0_n39, u0_n43, 
      u0_n47, u0_n49, u0_n59, u0_n63, u0_r0_N78, u0_r0_N79, u0_r0_N80, u0_r0_n3, u0_r0_n6, 
      u0_r0_n8, u0_r0_n9, u0_r0_rcnt_0, u0_r0_rcnt_1, u0_r0_rcnt_2, w0_0, w0_1, w0_10, w0_11, 
      w0_12, w0_13, w0_14, w0_15, w0_16, w0_17, w0_18, w0_19, w0_2, 
      w0_20, w0_21, w0_22, w0_23, w0_24, w0_25, w0_26, w0_27, w0_28, 
      w0_29, w0_3, w0_30, w0_31, w0_4, w0_5, w0_6, w0_7, w0_8, 
      w0_9, w1_0, w1_1, w1_10, w1_11, w1_12, w1_13, w1_14, w1_15, 
      w1_16, w1_17, w1_18, w1_19, w1_2, w1_20, w1_21, w1_22, w1_23, 
      w1_24, w1_25, w1_26, w1_27, w1_28, w1_29, w1_3, w1_30, w1_31, 
      w1_4, w1_5, w1_6, w1_7, w1_8, w1_9, w2_0, w2_1, w2_10, 
      w2_11, w2_12, w2_13, w2_14, w2_15, w2_16, w2_17, w2_18, w2_19, 
      w2_2, w2_20, w2_21, w2_22, w2_23, w2_24, w2_25, w2_26, w2_27, 
      w2_28, w2_29, w2_3, w2_30, w2_31, w2_4, w2_5, w2_6, w2_7, 
      w2_8, w2_9, w3_0, w3_1, w3_10, w3_11, w3_16, w3_17, w3_18, 
      w3_19, w3_2, w3_20, w3_21, w3_22, w3_23, w3_24, w3_25, w3_26, 
      w3_27, w3_28, w3_29, w3_3, w3_30, w3_31, w3_4, w3_5, w3_6, 
      w3_7, w3_8, w3_9, N100, N101, N102, N103, N104, N105, 
      N114, N115, N116, N117, N118, N119, N120, N121, N130, 
      N131, N132, N133, N134, N135, N136, N137, N146, N147, 
      N148, N149, N150, N151, N152, N153, N162, N163, N164, 
      N165, N166, N167, N168, N169, N178, N179, N180, N181, 
      N182, N183, N184, N185, N194, N195, N196, N197, N198, 
      N199, N200, N201, N210, N211, N212, N213, N214, N215, 
      N216, N217, N226, N227, N228, N229, N230, N231, N232, 
      N233, N242, N243, N244, N245, N246, N247, N248, N249, 
      N258, N259, N260, N261, N262, N263, N264, N265, N274, 
      N275, N276, N277, N278, N279, N280, N281, N34, N35, 
      N36, N37, N378, N379, N38, N382, N383, N384, N385, 
      N39, N392, N393, N394, N395, N398, N399, N40, N41, 
      N415, N419, N423, N441, N454, N455, N456, N457, N458, 
      N459, N460, N461, N463, N466, N467, N468, N469, N470, 
      N471, N472, N473, N474, N475, N476, N477, N478, N479, 
      N480, N481, N482, N483, N484, N485, N486, N487, N488, 
      N489, N490, N491, N492, N493, N494, N495, N496, N497, 
      N498, N499, N50, N500, N501, N502, N503, N504, N505, 
      N51, N52, N53, N54, N55, N56, N57, N66, N67, 
      N68, N69, N70, N71, N72, N73, N82, N83, N84, 
      N85, N86, N87, N88, N89, N98, N99, u0_n104, u0_n106, 
      u0_n107, u0_n109, u0_n113, u0_n115, u0_n116, u0_n118, u0_n119, u0_n121, u0_n122, 
      u0_n124, u0_n128, u0_n130, u0_n134, u0_n136, u0_n137, u0_n139, u0_n152, u0_n154, 
      u0_n158, u0_n160, u0_n176, u0_n188, u0_n190, u0_n194, u0_n196, u0_n198, u0_n200, 
      u0_n204, u0_n208, u0_n210, u0_n220, u0_n224, u0_n88, u0_r0_N70, u0_r0_N71, u0_r0_N72, 
      u0_r0_N73, u0_r0_N74, u0_r0_N75, u0_r0_N76, u0_r0_N77, u0_r0_N81, u0_r0_n12, u0_r0_n18 );
  aes_aes_die_9 u9 ( sa30_0, sa30_1, sa30_2, sa30_3, sa30_4, sa30_5, sa30_6, sa30_7, w0_0, 
      w0_2, w0_7, w3_24, w3_25, w3_26, w3_27, w3_28, w3_29, w3_30, 
      w3_31, sa31_sr_0, sa31_sr_1, sa31_sr_2, sa31_sr_3, sa31_sr_4, sa31_sr_5, sa31_sr_6, sa31_sr_7, 
      u0_n49, u0_n59, u0_n63, u0_subword_1, u0_subword_3, u0_subword_4, u0_subword_5, u0_subword_6 );
  aes_aes_die_10 u10 ( sa00_0, sa00_1, sa00_2, sa00_3, sa00_4, sa00_5, sa00_6, sa00_7, sa32_0, 
      sa32_1, sa32_2, sa32_3, sa32_4, sa32_5, sa32_6, sa32_7, sa00_sr_0, sa00_sr_1, 
      sa00_sr_2, sa00_sr_3, sa00_sr_4, sa00_sr_5, sa00_sr_6, sa00_sr_7, sa33_sr_0, sa33_sr_1, sa33_sr_2, 
      sa33_sr_3, sa33_sr_4, sa33_sr_5, sa33_sr_6, sa33_sr_7 );
  aes_aes_die_11 u11 ( u0_n268, u0_n270, u0_n272, u0_n274, w0_10, w0_12, w0_13, w0_14, w0_15, 
      w0_17, w0_18, w0_8, w3_0, w3_1, w3_10, w3_11, w3_2, w3_3, 
      w3_4, w3_5, w3_6, w3_7, w3_8, w3_9, u0_n27, u0_n29, u0_n33, 
      u0_n35, u0_n37, u0_n39, u0_n43, u0_n47, u0_subword_11, u0_subword_16, u0_subword_19, u0_subword_20, 
      u0_subword_21, u0_subword_22, u0_subword_23, u0_subword_9 );
endmodule
