module des_des_die_13 ( );
  input   output   wire endmodule

