module des_des ( clk, decrypt, desIn, key1, key2, key3, desOut );
  input clk;
  input decrypt;
  input [63:0] desIn;
  input [55:0] key1;
  input [55:0] key2;
  input [55:0] key3;
  output [63:0] desOut;

  wire n116, u0_FP_11, u0_FP_12, u0_FP_14, u0_FP_15, u0_FP_19, u0_FP_21, u0_FP_22, 
       u0_FP_25, u0_FP_27, u0_FP_29, u0_FP_3, u0_FP_32, u0_FP_33, u0_FP_34, u0_FP_36, u0_FP_37, 
       u0_FP_38, u0_FP_39, u0_FP_4, u0_FP_40, u0_FP_41, u0_FP_42, u0_FP_43, u0_FP_45, u0_FP_48, 
       u0_FP_49, u0_FP_5, u0_FP_50, u0_FP_51, u0_FP_52, u0_FP_53, u0_FP_54, u0_FP_55, u0_FP_56, 
       u0_FP_57, u0_FP_58, u0_FP_59, u0_FP_60, u0_FP_61, u0_FP_62, u0_FP_63, u0_FP_64, u0_FP_7, 
       u0_FP_8, u0_K10_10, u0_K10_13, u0_K10_14, u0_K10_18, u0_K10_19, u0_K10_20, u0_K10_25, u0_K10_32, 
       u0_K10_36, u0_K11_25, u0_K11_37, u0_K11_48, u0_K12_19, u0_K12_22, u0_K12_34, u0_K12_35, u0_K12_36, 
       u0_K12_39, u0_K12_40, u0_K12_48, u0_K12_7, u0_K12_9, u0_K13_30, u0_K13_36, u0_K13_38, u0_K13_8, 
       u0_K14_10, u0_K14_12, u0_K14_13, u0_K14_14, u0_K14_15, u0_K14_18, u0_K14_23, u0_K14_4, u0_K14_42, 
       u0_K14_9, u0_K15_18, u0_K15_47, u0_K16_11, u0_K16_18, u0_K16_24, u0_K16_26, u0_K16_38, u0_K16_8, 
       u0_K1_13, u0_K1_14, u0_K1_17, u0_K1_31, u0_K1_47, u0_K2_17, u0_K2_30, u0_K2_44, u0_K2_5, 
       u0_K2_6, u0_K2_8, u0_K3_12, u0_K3_13, u0_K3_14, u0_K3_17, u0_K3_18, u0_K3_19, u0_K3_23, 
       u0_K3_5, u0_K3_6, u0_K4_24, u0_K4_43, u0_K4_48, u0_K5_1, u0_K5_13, u0_K5_14, u0_K5_15, 
       u0_K5_16, u0_K5_18, u0_K5_19, u0_K5_23, u0_K5_24, u0_K5_26, u0_K5_28, u0_K5_3, u0_K5_31, 
       u0_K5_32, u0_K5_4, u0_K5_41, u0_K5_44, u0_K5_47, u0_K5_48, u0_K5_9, u0_K6_11, u0_K6_13, 
       u0_K6_20, u0_K6_23, u0_K7_2, u0_K7_23, u0_K8_1, u0_K8_11, u0_K8_13, u0_K8_19, u0_K8_23, 
       u0_K9_14, u0_K9_15, u0_K9_32, u0_K9_39, u0_K9_4, u0_K9_40, u0_K9_45, u0_K9_6, u0_L10_1, 
       u0_L10_10, u0_L10_11, u0_L10_12, u0_L10_13, u0_L10_14, u0_L10_15, u0_L10_16, u0_L10_17, u0_L10_18, 
       u0_L10_19, u0_L10_2, u0_L10_20, u0_L10_21, u0_L10_22, u0_L10_23, u0_L10_24, u0_L10_25, u0_L10_26, 
       u0_L10_27, u0_L10_28, u0_L10_29, u0_L10_3, u0_L10_30, u0_L10_31, u0_L10_32, u0_L10_4, u0_L10_5, 
       u0_L10_6, u0_L10_7, u0_L10_8, u0_L10_9, u0_L12_13, u0_L12_16, u0_L12_17, u0_L12_18, u0_L12_2, 
       u0_L12_23, u0_L12_24, u0_L12_28, u0_L12_30, u0_L12_31, u0_L12_6, u0_L12_9, u0_L13_1, u0_L13_10, 
       u0_L13_13, u0_L13_18, u0_L13_2, u0_L13_20, u0_L13_26, u0_L13_28, u0_L14_11, u0_L14_12, u0_L14_14, 
       u0_L14_15, u0_L14_19, u0_L14_21, u0_L14_22, u0_L14_25, u0_L14_27, u0_L14_29, u0_L14_3, u0_L14_32, 
       u0_L14_4, u0_L14_5, u0_L14_7, u0_L14_8, u0_L3_1, u0_L3_10, u0_L3_13, u0_L3_14, u0_L3_15, 
       u0_L3_16, u0_L3_17, u0_L3_18, u0_L3_2, u0_L3_20, u0_L3_21, u0_L3_23, u0_L3_24, u0_L3_25, 
       u0_L3_26, u0_L3_27, u0_L3_28, u0_L3_3, u0_L3_30, u0_L3_31, u0_L3_5, u0_L3_6, u0_L3_8, 
       u0_L3_9, u0_L7_1, u0_L7_10, u0_L7_11, u0_L7_12, u0_L7_13, u0_L7_14, u0_L7_15, u0_L7_16, 
       u0_L7_17, u0_L7_18, u0_L7_19, u0_L7_2, u0_L7_20, u0_L7_21, u0_L7_22, u0_L7_23, u0_L7_24, 
       u0_L7_25, u0_L7_26, u0_L7_27, u0_L7_28, u0_L7_29, u0_L7_3, u0_L7_30, u0_L7_31, u0_L7_32, 
       u0_L7_4, u0_L7_5, u0_L7_6, u0_L7_7, u0_L7_8, u0_L7_9, u0_L8_1, u0_L8_10, u0_L8_13, 
       u0_L8_16, u0_L8_17, u0_L8_18, u0_L8_2, u0_L8_20, u0_L8_23, u0_L8_24, u0_L8_26, u0_L8_28, 
       u0_L8_30, u0_L8_31, u0_L8_6, u0_L8_9, u0_N128, u0_N129, u0_N130, u0_N132, u0_N133, 
       u0_N135, u0_N136, u0_N137, u0_N140, u0_N141, u0_N142, u0_N143, u0_N144, u0_N145, 
       u0_N147, u0_N148, u0_N150, u0_N151, u0_N152, u0_N153, u0_N154, u0_N155, u0_N157, 
       u0_N158, u0_N256, u0_N257, u0_N258, u0_N259, u0_N260, u0_N261, u0_N262, u0_N263, 
       u0_N264, u0_N265, u0_N266, u0_N267, u0_N268, u0_N269, u0_N270, u0_N271, u0_N272, 
       u0_N273, u0_N274, u0_N275, u0_N276, u0_N277, u0_N278, u0_N279, u0_N280, u0_N281, 
       u0_N282, u0_N283, u0_N284, u0_N285, u0_N286, u0_N287, u0_N288, u0_N289, u0_N293, 
       u0_N296, u0_N297, u0_N300, u0_N303, u0_N304, u0_N305, u0_N307, u0_N310, u0_N311, 
       u0_N313, u0_N315, u0_N317, u0_N318, u0_N352, u0_N353, u0_N354, u0_N355, u0_N356, 
       u0_N357, u0_N358, u0_N359, u0_N360, u0_N361, u0_N362, u0_N363, u0_N364, u0_N365, 
       u0_N366, u0_N367, u0_N368, u0_N369, u0_N370, u0_N371, u0_N372, u0_N373, u0_N374, 
       u0_N375, u0_N376, u0_N377, u0_N378, u0_N379, u0_N380, u0_N381, u0_N382, u0_N383, 
       u0_N417, u0_N421, u0_N424, u0_N428, u0_N431, u0_N432, u0_N433, u0_N438, u0_N439, 
       u0_N443, u0_N445, u0_N446, u0_N448, u0_N449, u0_N457, u0_N460, u0_N465, u0_N467, 
       u0_N473, u0_N475, u0_R0_12, u0_R0_14, u0_R0_17, u0_R0_18, u0_R0_19, u0_R0_21, u0_R0_22, 
       u0_R0_25, u0_R0_27, u0_R0_28, u0_R0_29, u0_R0_4, u0_R0_5, u0_R10_1, u0_R10_10, u0_R10_11, 
       u0_R10_12, u0_R10_13, u0_R10_14, u0_R10_15, u0_R10_16, u0_R10_17, u0_R10_18, u0_R10_19, u0_R10_2, 
       u0_R10_20, u0_R10_21, u0_R10_22, u0_R10_23, u0_R10_24, u0_R10_25, u0_R10_26, u0_R10_27, u0_R10_28, 
       u0_R10_29, u0_R10_3, u0_R10_30, u0_R10_31, u0_R10_32, u0_R10_4, u0_R10_5, u0_R10_6, u0_R10_7, 
       u0_R10_8, u0_R10_9, u0_R11_10, u0_R11_11, u0_R11_12, u0_R11_13, u0_R11_14, u0_R11_15, u0_R11_16, 
       u0_R11_17, u0_R11_20, u0_R11_21, u0_R11_22, u0_R11_23, u0_R11_24, u0_R11_25, u0_R11_28, u0_R11_3, 
       u0_R11_32, u0_R11_4, u0_R11_5, u0_R11_6, u0_R11_7, u0_R11_8, u0_R11_9, u0_R12_1, u0_R12_10, 
       u0_R12_11, u0_R12_12, u0_R12_13, u0_R12_16, u0_R12_19, u0_R12_2, u0_R12_20, u0_R12_21, u0_R12_22, 
       u0_R12_23, u0_R12_24, u0_R12_25, u0_R12_26, u0_R12_28, u0_R12_29, u0_R12_3, u0_R12_30, u0_R12_32, 
       u0_R12_4, u0_R12_5, u0_R12_6, u0_R12_7, u0_R12_8, u0_R12_9, u0_R13_1, u0_R13_11, u0_R13_12, 
       u0_R13_13, u0_R13_14, u0_R13_15, u0_R13_16, u0_R13_17, u0_R13_18, u0_R13_19, u0_R13_2, u0_R13_20, 
       u0_R13_21, u0_R13_22, u0_R13_23, u0_R13_24, u0_R13_25, u0_R13_26, u0_R13_27, u0_R13_28, u0_R13_29, 
       u0_R13_3, u0_R13_30, u0_R13_31, u0_R13_32, u0_R13_4, u0_R13_5, u0_R13_6, u0_R13_7, u0_R13_8, 
       u0_R13_9, u0_R1_1, u0_R1_12, u0_R1_13, u0_R1_16, u0_R1_17, u0_R1_18, u0_R1_19, u0_R1_20, 
       u0_R1_21, u0_R1_22, u0_R1_24, u0_R1_25, u0_R1_26, u0_R1_27, u0_R1_28, u0_R1_29, u0_R1_3, 
       u0_R1_31, u0_R1_32, u0_R1_4, u0_R1_5, u0_R1_8, u0_R1_9, u0_R2_1, u0_R2_10, u0_R2_11, 
       u0_R2_12, u0_R2_13, u0_R2_14, u0_R2_15, u0_R2_16, u0_R2_17, u0_R2_20, u0_R2_21, u0_R2_22, 
       u0_R2_23, u0_R2_26, u0_R2_27, u0_R2_28, u0_R2_29, u0_R2_3, u0_R2_30, u0_R2_31, u0_R2_32, 
       u0_R2_4, u0_R2_6, u0_R2_7, u0_R2_8, u0_R2_9, u0_R3_1, u0_R3_10, u0_R3_11, u0_R3_12, 
       u0_R3_13, u0_R3_14, u0_R3_15, u0_R3_16, u0_R3_17, u0_R3_18, u0_R3_19, u0_R3_2, u0_R3_20, 
       u0_R3_21, u0_R3_22, u0_R3_24, u0_R3_27, u0_R3_28, u0_R3_29, u0_R3_3, u0_R3_30, u0_R3_31, 
       u0_R3_32, u0_R3_4, u0_R3_5, u0_R3_6, u0_R3_7, u0_R3_8, u0_R3_9, u0_R4_1, u0_R4_13, 
       u0_R4_14, u0_R4_16, u0_R4_22, u0_R4_24, u0_R4_29, u0_R4_30, u0_R4_8, u0_R5_1, u0_R5_11, 
       u0_R5_12, u0_R5_13, u0_R5_14, u0_R5_16, u0_R5_17, u0_R5_18, u0_R5_19, u0_R5_2, u0_R5_20, 
       u0_R5_21, u0_R5_22, u0_R5_23, u0_R5_24, u0_R5_25, u0_R5_26, u0_R5_27, u0_R5_28, u0_R5_29, 
       u0_R5_3, u0_R5_30, u0_R5_31, u0_R5_32, u0_R5_4, u0_R5_5, u0_R5_7, u0_R5_8, u0_R5_9, 
       u0_R6_1, u0_R6_10, u0_R6_11, u0_R6_12, u0_R6_13, u0_R6_14, u0_R6_16, u0_R6_17, u0_R6_18, 
       u0_R6_2, u0_R6_20, u0_R6_21, u0_R6_23, u0_R6_24, u0_R6_26, u0_R6_27, u0_R6_28, u0_R6_29, 
       u0_R6_32, u0_R6_4, u0_R6_5, u0_R6_7, u0_R6_8, u0_R6_9, u0_R7_1, u0_R7_10, u0_R7_11, 
       u0_R7_12, u0_R7_13, u0_R7_14, u0_R7_15, u0_R7_16, u0_R7_17, u0_R7_18, u0_R7_19, u0_R7_2, 
       u0_R7_20, u0_R7_21, u0_R7_22, u0_R7_23, u0_R7_24, u0_R7_25, u0_R7_26, u0_R7_27, u0_R7_28, 
       u0_R7_29, u0_R7_3, u0_R7_30, u0_R7_31, u0_R7_32, u0_R7_4, u0_R7_5, u0_R7_6, u0_R7_7, 
       u0_R7_8, u0_R7_9, u0_R8_1, u0_R8_10, u0_R8_11, u0_R8_12, u0_R8_13, u0_R8_14, u0_R8_15, 
       u0_R8_16, u0_R8_17, u0_R8_19, u0_R8_2, u0_R8_20, u0_R8_21, u0_R8_22, u0_R8_24, u0_R8_25, 
       u0_R8_27, u0_R8_29, u0_R8_3, u0_R8_30, u0_R8_32, u0_R8_4, u0_R8_5, u0_R8_6, u0_R8_7, 
       u0_R8_8, u0_R8_9, u0_R9_1, u0_R9_10, u0_R9_11, u0_R9_12, u0_R9_13, u0_R9_15, u0_R9_16, 
       u0_R9_17, u0_R9_18, u0_R9_19, u0_R9_2, u0_R9_20, u0_R9_21, u0_R9_22, u0_R9_23, u0_R9_24, 
       u0_R9_25, u0_R9_27, u0_R9_28, u0_R9_29, u0_R9_3, u0_R9_31, u0_R9_32, u0_R9_4, u0_R9_5, 
       u0_R9_6, u0_R9_7, u0_R9_8, u0_R9_9, u0_desIn_r_1, u0_desIn_r_11, u0_desIn_r_15, u0_desIn_r_25, u0_desIn_r_27, 
       u0_desIn_r_29, u0_desIn_r_3, u0_desIn_r_31, u0_desIn_r_33, u0_desIn_r_37, u0_desIn_r_39, u0_desIn_r_45, u0_desIn_r_47, u0_desIn_r_5, 
       u0_desIn_r_51, u0_desIn_r_53, u0_desIn_r_55, u0_desIn_r_57, u0_desIn_r_59, u0_desIn_r_63, u0_desIn_r_7, u0_key_r_11, u0_key_r_12, 
       u0_key_r_13, u0_key_r_14, u0_key_r_16, u0_key_r_17, u0_key_r_19, u0_key_r_2, u0_key_r_20, u0_key_r_21, u0_key_r_23, 
       u0_key_r_24, u0_key_r_25, u0_key_r_26, u0_key_r_27, u0_key_r_28, u0_key_r_30, u0_key_r_31, u0_key_r_32, u0_key_r_34, 
       u0_key_r_35, u0_key_r_36, u0_key_r_37, u0_key_r_38, u0_key_r_39, u0_key_r_4, u0_key_r_40, u0_key_r_41, u0_key_r_42, 
       u0_key_r_43, u0_key_r_47, u0_key_r_48, u0_key_r_5, u0_key_r_50, u0_key_r_51, u0_key_r_54, u0_key_r_55, u0_key_r_6, 
       u0_key_r_9, u0_out0_1, u0_out0_10, u0_out0_11, u0_out0_12, u0_out0_13, u0_out0_14, u0_out0_15, u0_out0_16, 
       u0_out0_17, u0_out0_18, u0_out0_19, u0_out0_2, u0_out0_20, u0_out0_21, u0_out0_22, u0_out0_23, u0_out0_24, 
       u0_out0_25, u0_out0_26, u0_out0_27, u0_out0_28, u0_out0_29, u0_out0_3, u0_out0_30, u0_out0_31, u0_out0_32, 
       u0_out0_4, u0_out0_5, u0_out0_6, u0_out0_7, u0_out0_8, u0_out0_9, u0_out10_1, u0_out10_10, u0_out10_11, 
       u0_out10_12, u0_out10_13, u0_out10_14, u0_out10_15, u0_out10_16, u0_out10_17, u0_out10_18, u0_out10_19, u0_out10_2, 
       u0_out10_20, u0_out10_21, u0_out10_22, u0_out10_23, u0_out10_24, u0_out10_25, u0_out10_26, u0_out10_27, u0_out10_28, 
       u0_out10_29, u0_out10_3, u0_out10_30, u0_out10_31, u0_out10_32, u0_out10_4, u0_out10_5, u0_out10_6, u0_out10_7, 
       u0_out10_8, u0_out10_9, u0_out12_1, u0_out12_10, u0_out12_11, u0_out12_12, u0_out12_13, u0_out12_14, u0_out12_15, 
       u0_out12_16, u0_out12_17, u0_out12_18, u0_out12_19, u0_out12_2, u0_out12_20, u0_out12_21, u0_out12_22, u0_out12_23, 
       u0_out12_24, u0_out12_25, u0_out12_26, u0_out12_27, u0_out12_28, u0_out12_29, u0_out12_3, u0_out12_30, u0_out12_31, 
       u0_out12_32, u0_out12_4, u0_out12_5, u0_out12_6, u0_out12_7, u0_out12_8, u0_out12_9, u0_out13_1, u0_out13_10, 
       u0_out13_11, u0_out13_12, u0_out13_14, u0_out13_15, u0_out13_19, u0_out13_20, u0_out13_21, u0_out13_22, u0_out13_25, 
       u0_out13_26, u0_out13_27, u0_out13_29, u0_out13_3, u0_out13_32, u0_out13_4, u0_out13_5, u0_out13_7, u0_out13_8, 
       u0_out14_11, u0_out14_12, u0_out14_14, u0_out14_15, u0_out14_16, u0_out14_17, u0_out14_19, u0_out14_21, u0_out14_22, 
       u0_out14_23, u0_out14_24, u0_out14_25, u0_out14_27, u0_out14_29, u0_out14_3, u0_out14_30, u0_out14_31, u0_out14_32, 
       u0_out14_4, u0_out14_5, u0_out14_6, u0_out14_7, u0_out14_8, u0_out14_9, u0_out15_1, u0_out15_10, u0_out15_13, 
       u0_out15_16, u0_out15_17, u0_out15_18, u0_out15_2, u0_out15_20, u0_out15_23, u0_out15_24, u0_out15_26, u0_out15_28, 
       u0_out15_30, u0_out15_31, u0_out15_6, u0_out15_9, u0_out1_1, u0_out1_10, u0_out1_11, u0_out1_12, u0_out1_13, 
       u0_out1_14, u0_out1_15, u0_out1_16, u0_out1_17, u0_out1_18, u0_out1_19, u0_out1_2, u0_out1_20, u0_out1_21, 
       u0_out1_22, u0_out1_23, u0_out1_24, u0_out1_25, u0_out1_26, u0_out1_27, u0_out1_28, u0_out1_29, u0_out1_3, 
       u0_out1_30, u0_out1_31, u0_out1_32, u0_out1_4, u0_out1_5, u0_out1_6, u0_out1_7, u0_out1_8, u0_out1_9, 
       u0_out2_1, u0_out2_10, u0_out2_11, u0_out2_12, u0_out2_13, u0_out2_14, u0_out2_15, u0_out2_16, u0_out2_17, 
       u0_out2_18, u0_out2_19, u0_out2_2, u0_out2_20, u0_out2_21, u0_out2_22, u0_out2_23, u0_out2_24, u0_out2_25, 
       u0_out2_26, u0_out2_27, u0_out2_28, u0_out2_29, u0_out2_3, u0_out2_30, u0_out2_31, u0_out2_32, u0_out2_4, 
       u0_out2_5, u0_out2_6, u0_out2_7, u0_out2_8, u0_out2_9, u0_out3_1, u0_out3_10, u0_out3_11, u0_out3_12, 
       u0_out3_13, u0_out3_14, u0_out3_15, u0_out3_16, u0_out3_17, u0_out3_18, u0_out3_19, u0_out3_2, u0_out3_20, 
       u0_out3_21, u0_out3_22, u0_out3_23, u0_out3_24, u0_out3_25, u0_out3_26, u0_out3_27, u0_out3_28, u0_out3_29, 
       u0_out3_3, u0_out3_30, u0_out3_31, u0_out3_32, u0_out3_4, u0_out3_5, u0_out3_6, u0_out3_7, u0_out3_8, 
       u0_out3_9, u0_out4_11, u0_out4_12, u0_out4_19, u0_out4_22, u0_out4_29, u0_out4_32, u0_out4_4, u0_out4_7, 
       u0_out5_1, u0_out5_10, u0_out5_11, u0_out5_12, u0_out5_13, u0_out5_14, u0_out5_15, u0_out5_16, u0_out5_17, 
       u0_out5_18, u0_out5_19, u0_out5_2, u0_out5_20, u0_out5_21, u0_out5_22, u0_out5_23, u0_out5_24, u0_out5_25, 
       u0_out5_26, u0_out5_27, u0_out5_28, u0_out5_29, u0_out5_3, u0_out5_30, u0_out5_31, u0_out5_32, u0_out5_4, 
       u0_out5_5, u0_out5_6, u0_out5_7, u0_out5_8, u0_out5_9, u0_out6_1, u0_out6_10, u0_out6_11, u0_out6_12, 
       u0_out6_13, u0_out6_14, u0_out6_15, u0_out6_16, u0_out6_17, u0_out6_18, u0_out6_19, u0_out6_2, u0_out6_20, 
       u0_out6_21, u0_out6_22, u0_out6_23, u0_out6_24, u0_out6_25, u0_out6_26, u0_out6_27, u0_out6_28, u0_out6_29, 
       u0_out6_3, u0_out6_30, u0_out6_31, u0_out6_32, u0_out6_4, u0_out6_5, u0_out6_6, u0_out6_7, u0_out6_8, 
       u0_out6_9, u0_out7_1, u0_out7_10, u0_out7_11, u0_out7_12, u0_out7_13, u0_out7_14, u0_out7_15, u0_out7_16, 
       u0_out7_17, u0_out7_18, u0_out7_19, u0_out7_2, u0_out7_20, u0_out7_21, u0_out7_22, u0_out7_23, u0_out7_24, 
       u0_out7_25, u0_out7_26, u0_out7_27, u0_out7_28, u0_out7_29, u0_out7_3, u0_out7_30, u0_out7_31, u0_out7_32, 
       u0_out7_4, u0_out7_5, u0_out7_6, u0_out7_7, u0_out7_8, u0_out7_9, u0_out9_11, u0_out9_12, u0_out9_14, 
       u0_out9_15, u0_out9_19, u0_out9_21, u0_out9_22, u0_out9_25, u0_out9_27, u0_out9_29, u0_out9_3, u0_out9_32, 
       u0_out9_4, u0_out9_5, u0_out9_7, u0_out9_8, u0_u0_X_15, u0_u0_X_16, u0_u0_X_23, u0_u0_X_25, u0_u0_X_28, 
       u0_u0_X_30, u0_u0_X_32, u0_u0_X_33, u0_u0_X_39, u0_u0_X_4, u0_u0_X_40, u0_u0_X_45, u0_u0_X_46, u0_u10_X_21, 
       u0_u10_X_39, u0_u10_X_45, u0_u12_X_2, u0_u12_X_27, u0_u12_X_28, u0_u12_X_3, u0_u12_X_39, u0_u12_X_40, u0_u12_X_42, 
       u0_u12_X_44, u0_u12_X_45, u0_u12_X_46, u0_u12_X_48, u0_u13_X_21, u0_u13_X_22, u0_u13_X_24, u0_u13_X_26, u0_u13_X_27, 
       u0_u13_X_40, u0_u13_X_46, u0_u14_X_15, u0_u15_X_17, u0_u15_X_19, u0_u15_X_21, u0_u15_X_22, u0_u15_X_4, u0_u1_X_1, 
       u0_u1_X_10, u0_u1_X_11, u0_u1_X_12, u0_u1_X_13, u0_u1_X_14, u0_u1_X_15, u0_u1_X_16, u0_u1_X_18, u0_u1_X_2, 
       u0_u1_X_20, u0_u1_X_22, u0_u1_X_23, u0_u1_X_25, u0_u1_X_29, u0_u1_X_3, u0_u1_X_31, u0_u1_X_34, u0_u1_X_35, 
       u0_u1_X_37, u0_u1_X_39, u0_u1_X_4, u0_u1_X_45, u0_u1_X_46, u0_u1_X_47, u0_u1_X_48, u0_u1_X_9, u0_u2_X_10, 
       u0_u2_X_15, u0_u2_X_16, u0_u2_X_21, u0_u2_X_22, u0_u2_X_3, u0_u2_X_34, u0_u2_X_45, u0_u2_X_9, u0_u3_X_27, 
       u0_u3_X_28, u0_u3_X_3, u0_u3_X_35, u0_u3_X_36, u0_u3_X_37, u0_u3_X_38, u0_u3_X_6, u0_u3_X_8, u0_u4_X_34, 
       u0_u4_X_36, u0_u4_X_38, u0_u4_X_39, u0_u5_X_1, u0_u5_X_10, u0_u5_X_12, u0_u5_X_14, u0_u5_X_15, u0_u5_X_16, 
       u0_u5_X_17, u0_u5_X_19, u0_u5_X_22, u0_u5_X_24, u0_u5_X_26, u0_u5_X_27, u0_u5_X_28, u0_u5_X_29, u0_u5_X_3, 
       u0_u5_X_30, u0_u5_X_31, u0_u5_X_32, u0_u5_X_34, u0_u5_X_36, u0_u5_X_38, u0_u5_X_39, u0_u5_X_4, u0_u5_X_40, 
       u0_u5_X_41, u0_u5_X_43, u0_u5_X_46, u0_u5_X_47, u0_u5_X_5, u0_u5_X_6, u0_u5_X_7, u0_u5_X_8, u0_u5_X_9, 
       u0_u6_X_15, u0_u6_X_22, u0_u6_X_9, u0_u7_X_22, u0_u7_X_28, u0_u7_X_33, u0_u7_X_36, u0_u7_X_38, u0_u7_X_4, 
       u0_u7_X_45, u0_u7_X_46, u0_u7_X_9, u0_u9_X_27, u0_u9_X_34, u0_u9_X_39, u0_u9_X_41, u0_u9_X_43, u0_u9_X_46, 
       u0_uk_K_r0_15, u0_uk_K_r0_2, u0_uk_K_r0_28, u0_uk_K_r0_31, u0_uk_K_r0_36, u0_uk_K_r0_49, u0_uk_K_r0_7, u0_uk_K_r10_10, u0_uk_K_r10_14, 
       u0_uk_K_r10_18, u0_uk_K_r10_23, u0_uk_K_r10_25, u0_uk_K_r10_27, u0_uk_K_r10_28, u0_uk_K_r10_32, u0_uk_K_r10_34, u0_uk_K_r10_37, u0_uk_K_r10_39, 
       u0_uk_K_r10_41, u0_uk_K_r10_42, u0_uk_K_r10_43, u0_uk_K_r10_44, u0_uk_K_r10_47, u0_uk_K_r10_48, u0_uk_K_r10_9, u0_uk_K_r11_11, u0_uk_K_r11_17, 
       u0_uk_K_r11_20, u0_uk_K_r11_25, u0_uk_K_r11_27, u0_uk_K_r11_29, u0_uk_K_r11_33, u0_uk_K_r11_34, u0_uk_K_r11_48, u0_uk_K_r11_53, u0_uk_K_r11_54, 
       u0_uk_K_r11_6, u0_uk_K_r12_10, u0_uk_K_r12_15, u0_uk_K_r12_16, u0_uk_K_r12_25, u0_uk_K_r12_33, u0_uk_K_r12_44, u0_uk_K_r12_47, u0_uk_K_r13_0, 
       u0_uk_K_r13_13, u0_uk_K_r13_17, u0_uk_K_r13_22, u0_uk_K_r13_25, u0_uk_K_r13_32, u0_uk_K_r13_35, u0_uk_K_r13_38, u0_uk_K_r13_4, u0_uk_K_r13_44, 
       u0_uk_K_r13_55, u0_uk_K_r14_11, u0_uk_K_r14_12, u0_uk_K_r14_15, u0_uk_K_r14_16, u0_uk_K_r14_18, u0_uk_K_r14_2, u0_uk_K_r14_43, u0_uk_K_r14_45, 
       u0_uk_K_r14_46, u0_uk_K_r14_50, u0_uk_K_r14_8, u0_uk_K_r14_9, u0_uk_K_r1_15, u0_uk_K_r1_21, u0_uk_K_r1_22, u0_uk_K_r1_42, u0_uk_K_r1_44, 
       u0_uk_K_r1_7, u0_uk_K_r2_13, u0_uk_K_r2_18, u0_uk_K_r2_20, u0_uk_K_r2_25, u0_uk_K_r2_27, u0_uk_K_r2_28, u0_uk_K_r2_33, u0_uk_K_r2_53, 
       u0_uk_K_r2_55, u0_uk_K_r3_10, u0_uk_K_r3_11, u0_uk_K_r3_14, u0_uk_K_r3_15, u0_uk_K_r3_19, u0_uk_K_r3_24, u0_uk_K_r3_35, u0_uk_K_r3_38, 
       u0_uk_K_r3_47, u0_uk_K_r3_9, u0_uk_K_r4_38, u0_uk_K_r5_10, u0_uk_K_r5_16, u0_uk_K_r5_17, u0_uk_K_r5_19, u0_uk_K_r5_32, u0_uk_K_r5_37, 
       u0_uk_K_r5_39, u0_uk_K_r5_4, u0_uk_K_r5_8, u0_uk_K_r6_0, u0_uk_K_r6_10, u0_uk_K_r6_14, u0_uk_K_r6_21, u0_uk_K_r6_22, u0_uk_K_r6_26, 
       u0_uk_K_r6_27, u0_uk_K_r6_29, u0_uk_K_r6_3, u0_uk_K_r6_31, u0_uk_K_r6_34, u0_uk_K_r6_46, u0_uk_K_r6_53, u0_uk_K_r6_7, u0_uk_K_r7_0, 
       u0_uk_K_r7_1, u0_uk_K_r7_13, u0_uk_K_r7_15, u0_uk_K_r7_2, u0_uk_K_r7_20, u0_uk_K_r7_22, u0_uk_K_r7_23, u0_uk_K_r7_24, u0_uk_K_r7_25, 
       u0_uk_K_r7_26, u0_uk_K_r7_27, u0_uk_K_r7_30, u0_uk_K_r7_32, u0_uk_K_r7_39, u0_uk_K_r7_48, u0_uk_K_r7_55, u0_uk_K_r7_6, u0_uk_K_r7_8, 
       u0_uk_K_r7_9, u0_uk_K_r8_13, u0_uk_K_r8_16, u0_uk_K_r8_17, u0_uk_K_r8_2, u0_uk_K_r8_22, u0_uk_K_r8_27, u0_uk_K_r8_32, u0_uk_K_r8_37, 
       u0_uk_K_r8_40, u0_uk_K_r8_41, u0_uk_K_r9_0, u0_uk_K_r9_1, u0_uk_K_r9_13, u0_uk_K_r9_19, u0_uk_K_r9_25, u0_uk_K_r9_27, u0_uk_K_r9_31, 
       u0_uk_K_r9_33, u0_uk_K_r9_35, u0_uk_K_r9_45, u0_uk_K_r9_49, u0_uk_K_r9_6, u0_uk_K_r9_9, u0_uk_n1, u0_uk_n10, u0_uk_n100, 
       u0_uk_n1000, u0_uk_n1001, u0_uk_n1002, u0_uk_n1004, u0_uk_n1008, u0_uk_n1009, u0_uk_n1012, u0_uk_n1019, u0_uk_n102, 
       u0_uk_n1020, u0_uk_n1021, u0_uk_n1024, u0_uk_n104, u0_uk_n106, u0_uk_n108, u0_uk_n109, u0_uk_n11, u0_uk_n110, 
       u0_uk_n112, u0_uk_n113, u0_uk_n115, u0_uk_n116, u0_uk_n117, u0_uk_n118, u0_uk_n12, u0_uk_n120, u0_uk_n121, 
       u0_uk_n122, u0_uk_n123, u0_uk_n124, u0_uk_n126, u0_uk_n127, u0_uk_n128, u0_uk_n129, u0_uk_n13, u0_uk_n130, 
       u0_uk_n131, u0_uk_n132, u0_uk_n135, u0_uk_n136, u0_uk_n137, u0_uk_n139, u0_uk_n14, u0_uk_n140, u0_uk_n141, 
       u0_uk_n142, u0_uk_n143, u0_uk_n144, u0_uk_n145, u0_uk_n146, u0_uk_n147, u0_uk_n148, u0_uk_n149, u0_uk_n15, 
       u0_uk_n150, u0_uk_n151, u0_uk_n152, u0_uk_n153, u0_uk_n154, u0_uk_n155, u0_uk_n156, u0_uk_n157, u0_uk_n159, 
       u0_uk_n16, u0_uk_n161, u0_uk_n162, u0_uk_n163, u0_uk_n164, u0_uk_n165, u0_uk_n166, u0_uk_n167, u0_uk_n168, 
       u0_uk_n169, u0_uk_n17, u0_uk_n170, u0_uk_n171, u0_uk_n172, u0_uk_n173, u0_uk_n174, u0_uk_n175, u0_uk_n176, 
       u0_uk_n177, u0_uk_n178, u0_uk_n179, u0_uk_n18, u0_uk_n180, u0_uk_n181, u0_uk_n182, u0_uk_n183, u0_uk_n184, 
       u0_uk_n185, u0_uk_n186, u0_uk_n187, u0_uk_n188, u0_uk_n189, u0_uk_n19, u0_uk_n190, u0_uk_n191, u0_uk_n193, 
       u0_uk_n194, u0_uk_n195, u0_uk_n196, u0_uk_n197, u0_uk_n198, u0_uk_n199, u0_uk_n20, u0_uk_n200, u0_uk_n201, 
       u0_uk_n202, u0_uk_n203, u0_uk_n204, u0_uk_n205, u0_uk_n206, u0_uk_n207, u0_uk_n208, u0_uk_n209, u0_uk_n21, 
       u0_uk_n210, u0_uk_n212, u0_uk_n213, u0_uk_n214, u0_uk_n215, u0_uk_n216, u0_uk_n217, u0_uk_n218, u0_uk_n219, 
       u0_uk_n22, u0_uk_n220, u0_uk_n221, u0_uk_n222, u0_uk_n223, u0_uk_n224, u0_uk_n225, u0_uk_n226, u0_uk_n227, 
       u0_uk_n228, u0_uk_n229, u0_uk_n23, u0_uk_n230, u0_uk_n231, u0_uk_n232, u0_uk_n233, u0_uk_n234, u0_uk_n235, 
       u0_uk_n238, u0_uk_n239, u0_uk_n24, u0_uk_n240, u0_uk_n241, u0_uk_n242, u0_uk_n243, u0_uk_n244, u0_uk_n245, 
       u0_uk_n246, u0_uk_n248, u0_uk_n249, u0_uk_n25, u0_uk_n250, u0_uk_n251, u0_uk_n252, u0_uk_n253, u0_uk_n254, 
       u0_uk_n255, u0_uk_n257, u0_uk_n258, u0_uk_n259, u0_uk_n26, u0_uk_n260, u0_uk_n261, u0_uk_n262, u0_uk_n263, 
       u0_uk_n264, u0_uk_n266, u0_uk_n267, u0_uk_n268, u0_uk_n269, u0_uk_n27, u0_uk_n272, u0_uk_n273, u0_uk_n274, 
       u0_uk_n275, u0_uk_n276, u0_uk_n278, u0_uk_n28, u0_uk_n280, u0_uk_n281, u0_uk_n282, u0_uk_n283, u0_uk_n285, 
       u0_uk_n288, u0_uk_n289, u0_uk_n29, u0_uk_n290, u0_uk_n293, u0_uk_n296, u0_uk_n3, u0_uk_n30, u0_uk_n300, 
       u0_uk_n303, u0_uk_n304, u0_uk_n307, u0_uk_n309, u0_uk_n31, u0_uk_n310, u0_uk_n311, u0_uk_n314, u0_uk_n315, 
       u0_uk_n316, u0_uk_n318, u0_uk_n32, u0_uk_n320, u0_uk_n321, u0_uk_n324, u0_uk_n325, u0_uk_n327, u0_uk_n329, 
       u0_uk_n33, u0_uk_n330, u0_uk_n331, u0_uk_n332, u0_uk_n333, u0_uk_n336, u0_uk_n337, u0_uk_n339, u0_uk_n34, 
       u0_uk_n341, u0_uk_n343, u0_uk_n344, u0_uk_n347, u0_uk_n348, u0_uk_n35, u0_uk_n352, u0_uk_n354, u0_uk_n355, 
       u0_uk_n358, u0_uk_n359, u0_uk_n36, u0_uk_n361, u0_uk_n362, u0_uk_n365, u0_uk_n367, u0_uk_n368, u0_uk_n37, 
       u0_uk_n370, u0_uk_n371, u0_uk_n372, u0_uk_n374, u0_uk_n378, u0_uk_n38, u0_uk_n380, u0_uk_n381, u0_uk_n383, 
       u0_uk_n384, u0_uk_n387, u0_uk_n388, u0_uk_n389, u0_uk_n39, u0_uk_n392, u0_uk_n393, u0_uk_n394, u0_uk_n396, 
       u0_uk_n398, u0_uk_n399, u0_uk_n4, u0_uk_n40, u0_uk_n400, u0_uk_n401, u0_uk_n402, u0_uk_n403, u0_uk_n405, 
       u0_uk_n406, u0_uk_n41, u0_uk_n412, u0_uk_n413, u0_uk_n418, u0_uk_n419, u0_uk_n42, u0_uk_n420, u0_uk_n425, 
       u0_uk_n429, u0_uk_n43, u0_uk_n430, u0_uk_n434, u0_uk_n44, u0_uk_n45, u0_uk_n451, u0_uk_n453, u0_uk_n455, 
       u0_uk_n457, u0_uk_n458, u0_uk_n459, u0_uk_n46, u0_uk_n462, u0_uk_n463, u0_uk_n464, u0_uk_n465, u0_uk_n466, 
       u0_uk_n471, u0_uk_n473, u0_uk_n475, u0_uk_n476, u0_uk_n479, u0_uk_n480, u0_uk_n481, u0_uk_n483, u0_uk_n484, 
       u0_uk_n485, u0_uk_n486, u0_uk_n488, u0_uk_n489, u0_uk_n490, u0_uk_n491, u0_uk_n493, u0_uk_n494, u0_uk_n497, 
       u0_uk_n498, u0_uk_n499, u0_uk_n5, u0_uk_n50, u0_uk_n502, u0_uk_n506, u0_uk_n508, u0_uk_n51, u0_uk_n510, 
       u0_uk_n511, u0_uk_n513, u0_uk_n514, u0_uk_n516, u0_uk_n517, u0_uk_n519, u0_uk_n52, u0_uk_n521, u0_uk_n522, 
       u0_uk_n523, u0_uk_n525, u0_uk_n528, u0_uk_n529, u0_uk_n53, u0_uk_n530, u0_uk_n531, u0_uk_n532, u0_uk_n534, 
       u0_uk_n535, u0_uk_n536, u0_uk_n537, u0_uk_n538, u0_uk_n539, u0_uk_n54, u0_uk_n543, u0_uk_n544, u0_uk_n545, 
       u0_uk_n546, u0_uk_n547, u0_uk_n549, u0_uk_n55, u0_uk_n550, u0_uk_n552, u0_uk_n553, u0_uk_n554, u0_uk_n555, 
       u0_uk_n557, u0_uk_n558, u0_uk_n559, u0_uk_n56, u0_uk_n560, u0_uk_n561, u0_uk_n562, u0_uk_n565, u0_uk_n566, 
       u0_uk_n568, u0_uk_n57, u0_uk_n570, u0_uk_n573, u0_uk_n574, u0_uk_n575, u0_uk_n578, u0_uk_n579, u0_uk_n58, 
       u0_uk_n580, u0_uk_n581, u0_uk_n584, u0_uk_n59, u0_uk_n592, u0_uk_n593, u0_uk_n599, u0_uk_n6, u0_uk_n60, 
       u0_uk_n600, u0_uk_n609, u0_uk_n61, u0_uk_n612, u0_uk_n616, u0_uk_n62, u0_uk_n620, u0_uk_n623, u0_uk_n624, 
       u0_uk_n629, u0_uk_n63, u0_uk_n630, u0_uk_n631, u0_uk_n632, u0_uk_n633, u0_uk_n635, u0_uk_n636, u0_uk_n637, 
       u0_uk_n638, u0_uk_n639, u0_uk_n64, u0_uk_n640, u0_uk_n641, u0_uk_n642, u0_uk_n643, u0_uk_n644, u0_uk_n645, 
       u0_uk_n647, u0_uk_n648, u0_uk_n649, u0_uk_n65, u0_uk_n650, u0_uk_n651, u0_uk_n652, u0_uk_n653, u0_uk_n655, 
       u0_uk_n657, u0_uk_n658, u0_uk_n659, u0_uk_n660, u0_uk_n663, u0_uk_n664, u0_uk_n666, u0_uk_n667, u0_uk_n668, 
       u0_uk_n669, u0_uk_n67, u0_uk_n670, u0_uk_n68, u0_uk_n684, u0_uk_n687, u0_uk_n69, u0_uk_n690, u0_uk_n696, 
       u0_uk_n697, u0_uk_n698, u0_uk_n7, u0_uk_n705, u0_uk_n707, u0_uk_n719, u0_uk_n72, u0_uk_n720, u0_uk_n725, 
       u0_uk_n726, u0_uk_n728, u0_uk_n73, u0_uk_n731, u0_uk_n732, u0_uk_n735, u0_uk_n736, u0_uk_n739, u0_uk_n740, 
       u0_uk_n746, u0_uk_n748, u0_uk_n75, u0_uk_n755, u0_uk_n759, u0_uk_n763, u0_uk_n765, u0_uk_n766, u0_uk_n768, 
       u0_uk_n77, u0_uk_n770, u0_uk_n771, u0_uk_n774, u0_uk_n775, u0_uk_n776, u0_uk_n78, u0_uk_n780, u0_uk_n783, 
       u0_uk_n793, u0_uk_n797, u0_uk_n799, u0_uk_n8, u0_uk_n80, u0_uk_n805, u0_uk_n81, u0_uk_n810, u0_uk_n813, 
       u0_uk_n815, u0_uk_n82, u0_uk_n826, u0_uk_n828, u0_uk_n829, u0_uk_n83, u0_uk_n831, u0_uk_n832, u0_uk_n834, 
       u0_uk_n839, u0_uk_n84, u0_uk_n85, u0_uk_n851, u0_uk_n855, u0_uk_n864, u0_uk_n87, u0_uk_n88, u0_uk_n89, 
       u0_uk_n897, u0_uk_n898, u0_uk_n9, u0_uk_n90, u0_uk_n904, u0_uk_n91, u0_uk_n915, u0_uk_n916, u0_uk_n917, 
       u0_uk_n918, u0_uk_n92, u0_uk_n93, u0_uk_n933, u0_uk_n934, u0_uk_n939, u0_uk_n94, u0_uk_n940, u0_uk_n948, 
       u0_uk_n949, u0_uk_n95, u0_uk_n950, u0_uk_n953, u0_uk_n96, u0_uk_n960, u0_uk_n963, u0_uk_n98, u0_uk_n981, 
       u0_uk_n982, u0_uk_n985, u0_uk_n99, u0_uk_n990, u0_uk_n992, u0_uk_n999, u1_FP_33, u1_FP_34, u1_FP_35, 
       u1_FP_36, u1_FP_37, u1_FP_38, u1_FP_39, u1_FP_40, u1_FP_41, u1_FP_42, u1_FP_43, u1_FP_44, 
       u1_FP_45, u1_FP_46, u1_FP_47, u1_FP_48, u1_FP_49, u1_FP_50, u1_FP_51, u1_FP_52, u1_FP_53, 
       u1_FP_54, u1_FP_55, u1_FP_56, u1_FP_57, u1_FP_58, u1_FP_59, u1_FP_60, u1_FP_61, u1_FP_62, 
       u1_FP_63, u1_FP_64, u1_K10_10, u1_K10_15, u1_K10_16, u1_K10_17, u1_K10_18, u1_K10_19, u1_K10_20, 
       u1_K10_21, u1_K10_27, u1_K10_28, u1_K10_34, u1_K10_45, u1_K10_46, u1_K11_1, u1_K11_10, u1_K11_11, 
       u1_K11_13, u1_K11_15, u1_K11_16, u1_K11_3, u1_K11_4, u1_K11_45, u1_K11_6, u1_K11_9, u1_K12_10, 
       u1_K12_11, u1_K12_12, u1_K12_13, u1_K12_14, u1_K12_16, u1_K12_33, u1_K12_34, u1_K12_36, u1_K12_38, 
       u1_K12_39, u1_K12_40, u1_K12_41, u1_K12_43, u1_K12_45, u1_K12_46, u1_K12_5, u1_K12_7, u1_K12_9, 
       u1_K13_1, u1_K13_24, u1_K13_26, u1_K13_27, u1_K13_28, u1_K13_3, u1_K13_33, u1_K13_34, u1_K13_35, 
       u1_K13_36, u1_K13_37, u1_K13_38, u1_K13_39, u1_K13_4, u1_K13_40, u1_K13_45, u1_K13_46, u1_K13_47, 
       u1_K13_8, u1_K13_9, u1_K14_10, u1_K14_12, u1_K14_14, u1_K14_15, u1_K14_16, u1_K14_21, u1_K14_22, 
       u1_K14_27, u1_K14_28, u1_K14_29, u1_K14_3, u1_K14_31, u1_K14_33, u1_K14_4, u1_K14_9, u1_K15_10, 
       u1_K15_12, u1_K15_14, u1_K15_15, u1_K15_16, u1_K15_17, u1_K15_18, u1_K15_19, u1_K15_20, u1_K15_21, 
       u1_K15_22, u1_K15_27, u1_K15_28, u1_K15_3, u1_K15_33, u1_K15_34, u1_K15_4, u1_K15_45, u1_K15_46, 
       u1_K15_5, u1_K15_6, u1_K15_7, u1_K15_9, u1_K16_10, u1_K16_15, u1_K16_16, u1_K16_21, u1_K16_22, 
       u1_K16_24, u1_K16_26, u1_K16_27, u1_K16_28, u1_K16_3, u1_K16_39, u1_K16_4, u1_K16_40, u1_K16_6, 
       u1_K16_8, u1_K16_9, u1_K1_12, u1_K1_14, u1_K1_15, u1_K1_16, u1_K1_21, u1_K1_3, u1_K1_34, 
       u1_K1_39, u1_K1_4, u1_K1_40, u1_K1_43, u1_K1_45, u1_K1_46, u1_K1_9, u1_K2_1, u1_K2_21, 
       u1_K2_22, u1_K2_3, u1_K2_33, u1_K2_34, u1_K2_39, u1_K2_4, u1_K2_40, u1_K2_45, u1_K2_46, 
       u1_K2_47, u1_K3_10, u1_K3_15, u1_K3_16, u1_K3_27, u1_K3_28, u1_K3_3, u1_K3_39, u1_K3_4, 
       u1_K3_40, u1_K3_5, u1_K3_7, u1_K3_9, u1_K4_15, u1_K4_16, u1_K4_17, u1_K4_18, u1_K4_19, 
       u1_K4_21, u1_K4_22, u1_K4_24, u1_K4_27, u1_K4_28, u1_K4_39, u1_K4_40, u1_K4_45, u1_K4_46, 
       u1_K4_9, u1_K5_10, u1_K5_15, u1_K5_16, u1_K5_18, u1_K5_21, u1_K5_23, u1_K5_24, u1_K5_25, 
       u1_K5_26, u1_K5_28, u1_K5_29, u1_K5_30, u1_K5_31, u1_K5_32, u1_K5_33, u1_K5_34, u1_K5_37, 
       u1_K5_38, u1_K5_39, u1_K5_40, u1_K5_41, u1_K5_45, u1_K5_46, u1_K5_9, u1_K6_1, u1_K6_22, 
       u1_K6_3, u1_K6_33, u1_K6_34, u1_K6_35, u1_K6_36, u1_K6_37, u1_K6_38, u1_K6_39, u1_K6_40, 
       u1_K6_41, u1_K6_42, u1_K6_43, u1_K6_44, u1_K6_45, u1_K6_46, u1_K6_47, u1_K6_48, u1_K6_6, 
       u1_K6_8, u1_K7_10, u1_K7_11, u1_K7_14, u1_K7_15, u1_K7_16, u1_K7_17, u1_K7_18, u1_K7_19, 
       u1_K7_21, u1_K7_22, u1_K7_23, u1_K7_26, u1_K7_28, u1_K7_29, u1_K7_3, u1_K7_30, u1_K7_31, 
       u1_K7_33, u1_K7_39, u1_K7_4, u1_K7_40, u1_K7_41, u1_K7_43, u1_K7_45, u1_K7_5, u1_K7_7, 
       u1_K7_9, u1_K8_10, u1_K8_11, u1_K8_13, u1_K8_14, u1_K8_16, u1_K8_18, u1_K8_20, u1_K8_21, 
       u1_K8_22, u1_K8_23, u1_K8_25, u1_K8_27, u1_K8_28, u1_K8_4, u1_K8_45, u1_K8_46, u1_K8_5, 
       u1_K8_6, u1_K8_7, u1_K8_8, u1_K8_9, u1_K9_13, u1_K9_15, u1_K9_16, u1_K9_17, u1_K9_21, 
       u1_K9_23, u1_K9_24, u1_K9_25, u1_K9_28, u1_K9_3, u1_K9_34, u1_K9_36, u1_K9_37, u1_K9_38, 
       u1_K9_39, u1_K9_4, u1_K9_40, u1_R0_1, u1_R0_10, u1_R0_11, u1_R0_12, u1_R0_13, u1_R0_14, 
       u1_R0_15, u1_R0_16, u1_R0_17, u1_R0_18, u1_R0_19, u1_R0_2, u1_R0_20, u1_R0_21, u1_R0_22, 
       u1_R0_23, u1_R0_24, u1_R0_25, u1_R0_26, u1_R0_27, u1_R0_28, u1_R0_29, u1_R0_3, u1_R0_30, 
       u1_R0_31, u1_R0_32, u1_R0_4, u1_R0_5, u1_R0_6, u1_R0_7, u1_R0_8, u1_R0_9, u1_R10_1, 
       u1_R10_10, u1_R10_11, u1_R10_12, u1_R10_13, u1_R10_14, u1_R10_15, u1_R10_16, u1_R10_17, u1_R10_18, 
       u1_R10_19, u1_R10_2, u1_R10_20, u1_R10_21, u1_R10_22, u1_R10_23, u1_R10_24, u1_R10_25, u1_R10_26, 
       u1_R10_27, u1_R10_28, u1_R10_29, u1_R10_3, u1_R10_30, u1_R10_31, u1_R10_32, u1_R10_4, u1_R10_5, 
       u1_R10_6, u1_R10_7, u1_R10_8, u1_R10_9, u1_R11_1, u1_R11_10, u1_R11_11, u1_R11_12, u1_R11_13, 
       u1_R11_14, u1_R11_15, u1_R11_16, u1_R11_17, u1_R11_18, u1_R11_19, u1_R11_2, u1_R11_20, u1_R11_21, 
       u1_R11_22, u1_R11_23, u1_R11_24, u1_R11_25, u1_R11_26, u1_R11_27, u1_R11_28, u1_R11_29, u1_R11_3, 
       u1_R11_30, u1_R11_31, u1_R11_32, u1_R11_4, u1_R11_5, u1_R11_6, u1_R11_7, u1_R11_8, u1_R11_9, 
       u1_R12_1, u1_R12_10, u1_R12_11, u1_R12_12, u1_R12_13, u1_R12_14, u1_R12_15, u1_R12_16, u1_R12_17, 
       u1_R12_18, u1_R12_19, u1_R12_2, u1_R12_20, u1_R12_21, u1_R12_22, u1_R12_23, u1_R12_24, u1_R12_25, 
       u1_R12_26, u1_R12_27, u1_R12_28, u1_R12_29, u1_R12_3, u1_R12_30, u1_R12_31, u1_R12_32, u1_R12_4, 
       u1_R12_5, u1_R12_6, u1_R12_7, u1_R12_8, u1_R12_9, u1_R13_1, u1_R13_10, u1_R13_11, u1_R13_12, 
       u1_R13_13, u1_R13_14, u1_R13_15, u1_R13_16, u1_R13_17, u1_R13_18, u1_R13_19, u1_R13_2, u1_R13_20, 
       u1_R13_21, u1_R13_22, u1_R13_23, u1_R13_24, u1_R13_25, u1_R13_26, u1_R13_27, u1_R13_28, u1_R13_29, 
       u1_R13_3, u1_R13_30, u1_R13_31, u1_R13_32, u1_R13_4, u1_R13_5, u1_R13_6, u1_R13_7, u1_R13_8, 
       u1_R13_9, u1_R1_1, u1_R1_10, u1_R1_11, u1_R1_12, u1_R1_13, u1_R1_14, u1_R1_15, u1_R1_16, 
       u1_R1_17, u1_R1_18, u1_R1_19, u1_R1_2, u1_R1_20, u1_R1_21, u1_R1_22, u1_R1_23, u1_R1_24, 
       u1_R1_25, u1_R1_26, u1_R1_27, u1_R1_28, u1_R1_29, u1_R1_3, u1_R1_30, u1_R1_31, u1_R1_32, 
       u1_R1_4, u1_R1_5, u1_R1_6, u1_R1_7, u1_R1_8, u1_R1_9, u1_R2_1, u1_R2_10, u1_R2_11, 
       u1_R2_12, u1_R2_13, u1_R2_14, u1_R2_15, u1_R2_16, u1_R2_17, u1_R2_18, u1_R2_19, u1_R2_2, 
       u1_R2_20, u1_R2_21, u1_R2_22, u1_R2_23, u1_R2_24, u1_R2_25, u1_R2_26, u1_R2_27, u1_R2_28, 
       u1_R2_29, u1_R2_3, u1_R2_30, u1_R2_31, u1_R2_32, u1_R2_4, u1_R2_5, u1_R2_6, u1_R2_7, 
       u1_R2_8, u1_R2_9, u1_R3_1, u1_R3_10, u1_R3_11, u1_R3_12, u1_R3_13, u1_R3_14, u1_R3_15, 
       u1_R3_16, u1_R3_17, u1_R3_18, u1_R3_19, u1_R3_2, u1_R3_20, u1_R3_21, u1_R3_22, u1_R3_23, 
       u1_R3_24, u1_R3_25, u1_R3_26, u1_R3_27, u1_R3_28, u1_R3_29, u1_R3_3, u1_R3_30, u1_R3_31, 
       u1_R3_32, u1_R3_4, u1_R3_5, u1_R3_6, u1_R3_7, u1_R3_8, u1_R3_9, u1_R4_1, u1_R4_10, 
       u1_R4_11, u1_R4_12, u1_R4_13, u1_R4_14, u1_R4_15, u1_R4_16, u1_R4_17, u1_R4_18, u1_R4_19, 
       u1_R4_2, u1_R4_20, u1_R4_21, u1_R4_22, u1_R4_23, u1_R4_24, u1_R4_25, u1_R4_26, u1_R4_27, 
       u1_R4_28, u1_R4_29, u1_R4_3, u1_R4_30, u1_R4_31, u1_R4_32, u1_R4_4, u1_R4_5, u1_R4_6, 
       u1_R4_7, u1_R4_8, u1_R4_9, u1_R5_1, u1_R5_10, u1_R5_11, u1_R5_12, u1_R5_13, u1_R5_14, 
       u1_R5_15, u1_R5_16, u1_R5_17, u1_R5_18, u1_R5_19, u1_R5_2, u1_R5_20, u1_R5_21, u1_R5_22, 
       u1_R5_23, u1_R5_24, u1_R5_25, u1_R5_26, u1_R5_27, u1_R5_28, u1_R5_29, u1_R5_3, u1_R5_30, 
       u1_R5_31, u1_R5_32, u1_R5_4, u1_R5_5, u1_R5_6, u1_R5_7, u1_R5_8, u1_R5_9, u1_R6_1, 
       u1_R6_10, u1_R6_11, u1_R6_12, u1_R6_13, u1_R6_14, u1_R6_15, u1_R6_16, u1_R6_17, u1_R6_18, 
       u1_R6_19, u1_R6_2, u1_R6_20, u1_R6_21, u1_R6_22, u1_R6_23, u1_R6_24, u1_R6_25, u1_R6_26, 
       u1_R6_27, u1_R6_28, u1_R6_29, u1_R6_3, u1_R6_30, u1_R6_31, u1_R6_32, u1_R6_4, u1_R6_5, 
       u1_R6_6, u1_R6_7, u1_R6_8, u1_R6_9, u1_R7_1, u1_R7_10, u1_R7_11, u1_R7_12, u1_R7_13, 
       u1_R7_14, u1_R7_15, u1_R7_16, u1_R7_17, u1_R7_18, u1_R7_19, u1_R7_2, u1_R7_20, u1_R7_21, 
       u1_R7_22, u1_R7_23, u1_R7_24, u1_R7_25, u1_R7_26, u1_R7_27, u1_R7_28, u1_R7_29, u1_R7_3, 
       u1_R7_30, u1_R7_31, u1_R7_32, u1_R7_4, u1_R7_5, u1_R7_6, u1_R7_7, u1_R7_8, u1_R7_9, 
       u1_R8_1, u1_R8_10, u1_R8_11, u1_R8_12, u1_R8_13, u1_R8_14, u1_R8_15, u1_R8_16, u1_R8_17, 
       u1_R8_18, u1_R8_19, u1_R8_2, u1_R8_20, u1_R8_21, u1_R8_22, u1_R8_23, u1_R8_24, u1_R8_25, 
       u1_R8_26, u1_R8_27, u1_R8_28, u1_R8_29, u1_R8_3, u1_R8_30, u1_R8_31, u1_R8_32, u1_R8_4, 
       u1_R8_5, u1_R8_6, u1_R8_7, u1_R8_8, u1_R8_9, u1_R9_1, u1_R9_10, u1_R9_11, u1_R9_12, 
       u1_R9_13, u1_R9_14, u1_R9_15, u1_R9_16, u1_R9_17, u1_R9_18, u1_R9_19, u1_R9_2, u1_R9_20, 
       u1_R9_21, u1_R9_22, u1_R9_23, u1_R9_24, u1_R9_25, u1_R9_26, u1_R9_27, u1_R9_28, u1_R9_29, 
       u1_R9_3, u1_R9_30, u1_R9_31, u1_R9_32, u1_R9_4, u1_R9_5, u1_R9_6, u1_R9_7, u1_R9_8, 
       u1_R9_9, u1_desIn_r_1, u1_desIn_r_11, u1_desIn_r_13, u1_desIn_r_15, u1_desIn_r_17, u1_desIn_r_19, u1_desIn_r_21, u1_desIn_r_23, 
       u1_desIn_r_25, u1_desIn_r_27, u1_desIn_r_29, u1_desIn_r_3, u1_desIn_r_31, u1_desIn_r_33, u1_desIn_r_35, u1_desIn_r_37, u1_desIn_r_39, 
       u1_desIn_r_41, u1_desIn_r_43, u1_desIn_r_45, u1_desIn_r_47, u1_desIn_r_49, u1_desIn_r_5, u1_desIn_r_51, u1_desIn_r_53, u1_desIn_r_55, 
       u1_desIn_r_57, u1_desIn_r_59, u1_desIn_r_61, u1_desIn_r_63, u1_desIn_r_7, u1_desIn_r_9, u1_key_r_0, u1_key_r_1, u1_key_r_10, 
       u1_key_r_11, u1_key_r_12, u1_key_r_13, u1_key_r_14, u1_key_r_15, u1_key_r_16, u1_key_r_17, u1_key_r_18, u1_key_r_19, 
       u1_key_r_2, u1_key_r_20, u1_key_r_21, u1_key_r_22, u1_key_r_23, u1_key_r_24, u1_key_r_25, u1_key_r_26, u1_key_r_27, 
       u1_key_r_28, u1_key_r_29, u1_key_r_3, u1_key_r_30, u1_key_r_31, u1_key_r_32, u1_key_r_33, u1_key_r_34, u1_key_r_35, 
       u1_key_r_36, u1_key_r_37, u1_key_r_38, u1_key_r_39, u1_key_r_4, u1_key_r_40, u1_key_r_41, u1_key_r_42, u1_key_r_43, 
       u1_key_r_44, u1_key_r_45, u1_key_r_46, u1_key_r_47, u1_key_r_48, u1_key_r_49, u1_key_r_5, u1_key_r_50, u1_key_r_51, 
       u1_key_r_52, u1_key_r_53, u1_key_r_54, u1_key_r_55, u1_key_r_6, u1_key_r_7, u1_key_r_8, u1_key_r_9, u1_out0_1, 
       u1_out0_10, u1_out0_11, u1_out0_12, u1_out0_13, u1_out0_14, u1_out0_15, u1_out0_16, u1_out0_17, u1_out0_18, 
       u1_out0_19, u1_out0_2, u1_out0_20, u1_out0_21, u1_out0_22, u1_out0_23, u1_out0_24, u1_out0_25, u1_out0_26, 
       u1_out0_27, u1_out0_28, u1_out0_29, u1_out0_3, u1_out0_30, u1_out0_31, u1_out0_32, u1_out0_4, u1_out0_5, 
       u1_out0_6, u1_out0_7, u1_out0_8, u1_out0_9, u1_out10_1, u1_out10_10, u1_out10_11, u1_out10_12, u1_out10_13, 
       u1_out10_14, u1_out10_15, u1_out10_16, u1_out10_17, u1_out10_18, u1_out10_19, u1_out10_2, u1_out10_20, u1_out10_21, 
       u1_out10_22, u1_out10_23, u1_out10_24, u1_out10_25, u1_out10_26, u1_out10_27, u1_out10_28, u1_out10_29, u1_out10_3, 
       u1_out10_30, u1_out10_31, u1_out10_32, u1_out10_4, u1_out10_5, u1_out10_6, u1_out10_7, u1_out10_8, u1_out10_9, 
       u1_out11_1, u1_out11_10, u1_out11_11, u1_out11_12, u1_out11_13, u1_out11_14, u1_out11_15, u1_out11_16, u1_out11_17, 
       u1_out11_18, u1_out11_19, u1_out11_2, u1_out11_20, u1_out11_21, u1_out11_22, u1_out11_23, u1_out11_24, u1_out11_25, 
       u1_out11_26, u1_out11_27, u1_out11_28, u1_out11_29, u1_out11_3, u1_out11_30, u1_out11_31, u1_out11_32, u1_out11_4, 
       u1_out11_5, u1_out11_6, u1_out11_7, u1_out11_8, u1_out11_9, u1_out12_1, u1_out12_10, u1_out12_11, u1_out12_12, 
       u1_out12_13, u1_out12_14, u1_out12_15, u1_out12_16, u1_out12_17, u1_out12_18, u1_out12_19, u1_out12_2, u1_out12_20, 
       u1_out12_21, u1_out12_22, u1_out12_23, u1_out12_24, u1_out12_25, u1_out12_26, u1_out12_27, u1_out12_28, u1_out12_29, 
       u1_out12_3, u1_out12_30, u1_out12_31, u1_out12_32, u1_out12_4, u1_out12_5, u1_out12_6, u1_out12_7, u1_out12_8, 
       u1_out12_9, u1_out13_1, u1_out13_10, u1_out13_11, u1_out13_12, u1_out13_13, u1_out13_14, u1_out13_15, u1_out13_16, 
       u1_out13_17, u1_out13_18, u1_out13_19, u1_out13_2, u1_out13_20, u1_out13_21, u1_out13_22, u1_out13_23, u1_out13_24, 
       u1_out13_25, u1_out13_26, u1_out13_27, u1_out13_28, u1_out13_29, u1_out13_3, u1_out13_30, u1_out13_31, u1_out13_32, 
       u1_out13_4, u1_out13_5, u1_out13_6, u1_out13_7, u1_out13_8, u1_out13_9, u1_out14_1, u1_out14_10, u1_out14_11, 
       u1_out14_12, u1_out14_13, u1_out14_14, u1_out14_15, u1_out14_16, u1_out14_17, u1_out14_18, u1_out14_19, u1_out14_2, 
       u1_out14_20, u1_out14_21, u1_out14_22, u1_out14_23, u1_out14_24, u1_out14_25, u1_out14_26, u1_out14_27, u1_out14_28, 
       u1_out14_29, u1_out14_3, u1_out14_30, u1_out14_31, u1_out14_32, u1_out14_4, u1_out14_5, u1_out14_6, u1_out14_7, 
       u1_out14_8, u1_out14_9, u1_out15_1, u1_out15_10, u1_out15_11, u1_out15_12, u1_out15_13, u1_out15_14, u1_out15_15, 
       u1_out15_16, u1_out15_17, u1_out15_18, u1_out15_19, u1_out15_2, u1_out15_20, u1_out15_21, u1_out15_22, u1_out15_23, 
       u1_out15_24, u1_out15_25, u1_out15_26, u1_out15_27, u1_out15_28, u1_out15_29, u1_out15_3, u1_out15_30, u1_out15_31, 
       u1_out15_32, u1_out15_4, u1_out15_5, u1_out15_6, u1_out15_7, u1_out15_8, u1_out15_9, u1_out1_1, u1_out1_10, 
       u1_out1_11, u1_out1_12, u1_out1_13, u1_out1_14, u1_out1_15, u1_out1_16, u1_out1_17, u1_out1_18, u1_out1_19, 
       u1_out1_2, u1_out1_20, u1_out1_21, u1_out1_22, u1_out1_23, u1_out1_24, u1_out1_25, u1_out1_26, u1_out1_27, 
       u1_out1_28, u1_out1_29, u1_out1_3, u1_out1_30, u1_out1_31, u1_out1_32, u1_out1_4, u1_out1_5, u1_out1_6, 
       u1_out1_7, u1_out1_8, u1_out1_9, u1_out2_1, u1_out2_10, u1_out2_11, u1_out2_12, u1_out2_13, u1_out2_14, 
       u1_out2_15, u1_out2_16, u1_out2_17, u1_out2_18, u1_out2_19, u1_out2_2, u1_out2_20, u1_out2_21, u1_out2_22, 
       u1_out2_23, u1_out2_24, u1_out2_25, u1_out2_26, u1_out2_27, u1_out2_28, u1_out2_29, u1_out2_3, u1_out2_30, 
       u1_out2_31, u1_out2_32, u1_out2_4, u1_out2_5, u1_out2_6, u1_out2_7, u1_out2_8, u1_out2_9, u1_out3_1, 
       u1_out3_10, u1_out3_11, u1_out3_12, u1_out3_13, u1_out3_14, u1_out3_15, u1_out3_16, u1_out3_17, u1_out3_18, 
       u1_out3_19, u1_out3_2, u1_out3_20, u1_out3_21, u1_out3_22, u1_out3_23, u1_out3_24, u1_out3_25, u1_out3_26, 
       u1_out3_27, u1_out3_28, u1_out3_29, u1_out3_3, u1_out3_30, u1_out3_31, u1_out3_32, u1_out3_4, u1_out3_5, 
       u1_out3_6, u1_out3_7, u1_out3_8, u1_out3_9, u1_out4_1, u1_out4_10, u1_out4_11, u1_out4_12, u1_out4_13, 
       u1_out4_14, u1_out4_15, u1_out4_16, u1_out4_17, u1_out4_18, u1_out4_19, u1_out4_2, u1_out4_20, u1_out4_21, 
       u1_out4_22, u1_out4_23, u1_out4_24, u1_out4_25, u1_out4_26, u1_out4_27, u1_out4_28, u1_out4_29, u1_out4_3, 
       u1_out4_30, u1_out4_31, u1_out4_32, u1_out4_4, u1_out4_5, u1_out4_6, u1_out4_7, u1_out4_8, u1_out4_9, 
       u1_out5_1, u1_out5_10, u1_out5_11, u1_out5_12, u1_out5_13, u1_out5_14, u1_out5_15, u1_out5_16, u1_out5_17, 
       u1_out5_18, u1_out5_19, u1_out5_2, u1_out5_20, u1_out5_21, u1_out5_22, u1_out5_23, u1_out5_24, u1_out5_25, 
       u1_out5_26, u1_out5_27, u1_out5_28, u1_out5_29, u1_out5_3, u1_out5_30, u1_out5_31, u1_out5_32, u1_out5_4, 
       u1_out5_5, u1_out5_6, u1_out5_7, u1_out5_8, u1_out5_9, u1_out6_1, u1_out6_10, u1_out6_11, u1_out6_12, 
       u1_out6_13, u1_out6_14, u1_out6_15, u1_out6_16, u1_out6_17, u1_out6_18, u1_out6_19, u1_out6_2, u1_out6_20, 
       u1_out6_21, u1_out6_22, u1_out6_23, u1_out6_24, u1_out6_25, u1_out6_26, u1_out6_27, u1_out6_28, u1_out6_29, 
       u1_out6_3, u1_out6_30, u1_out6_31, u1_out6_32, u1_out6_4, u1_out6_5, u1_out6_6, u1_out6_7, u1_out6_8, 
       u1_out6_9, u1_out7_1, u1_out7_10, u1_out7_11, u1_out7_12, u1_out7_13, u1_out7_14, u1_out7_15, u1_out7_16, 
       u1_out7_17, u1_out7_18, u1_out7_19, u1_out7_2, u1_out7_20, u1_out7_21, u1_out7_22, u1_out7_23, u1_out7_24, 
       u1_out7_25, u1_out7_26, u1_out7_27, u1_out7_28, u1_out7_29, u1_out7_3, u1_out7_30, u1_out7_31, u1_out7_32, 
       u1_out7_4, u1_out7_5, u1_out7_6, u1_out7_7, u1_out7_8, u1_out7_9, u1_out8_1, u1_out8_10, u1_out8_11, 
       u1_out8_12, u1_out8_13, u1_out8_14, u1_out8_15, u1_out8_16, u1_out8_17, u1_out8_18, u1_out8_19, u1_out8_2, 
       u1_out8_20, u1_out8_21, u1_out8_22, u1_out8_23, u1_out8_24, u1_out8_25, u1_out8_26, u1_out8_27, u1_out8_28, 
       u1_out8_29, u1_out8_3, u1_out8_30, u1_out8_31, u1_out8_32, u1_out8_4, u1_out8_5, u1_out8_6, u1_out8_7, 
       u1_out8_8, u1_out8_9, u1_out9_1, u1_out9_10, u1_out9_11, u1_out9_12, u1_out9_13, u1_out9_14, u1_out9_15, 
       u1_out9_16, u1_out9_17, u1_out9_18, u1_out9_19, u1_out9_2, u1_out9_20, u1_out9_21, u1_out9_22, u1_out9_23, 
       u1_out9_24, u1_out9_25, u1_out9_26, u1_out9_27, u1_out9_28, u1_out9_29, u1_out9_3, u1_out9_30, u1_out9_31, 
       u1_out9_32, u1_out9_4, u1_out9_5, u1_out9_6, u1_out9_7, u1_out9_8, u1_out9_9, u1_u0_X_1, u1_u0_X_11, 
       u1_u0_X_13, u1_u0_X_17, u1_u0_X_18, u1_u0_X_19, u1_u0_X_2, u1_u0_X_20, u1_u0_X_23, u1_u0_X_24, u1_u0_X_31, 
       u1_u0_X_32, u1_u0_X_35, u1_u0_X_36, u1_u0_X_37, u1_u0_X_38, u1_u0_X_47, u1_u0_X_48, u1_u0_X_5, u1_u0_X_6, 
       u1_u0_X_7, u1_u0_X_8, u1_u10_X_17, u1_u10_X_18, u1_u10_X_2, u1_u10_X_43, u1_u10_X_44, u1_u10_X_48, u1_u10_X_5, 
       u1_u10_X_7, u1_u11_X_1, u1_u11_X_17, u1_u11_X_18, u1_u11_X_2, u1_u11_X_31, u1_u11_X_32, u1_u11_X_35, u1_u11_X_37, 
       u1_u11_X_42, u1_u11_X_44, u1_u11_X_47, u1_u11_X_48, u1_u11_X_6, u1_u11_X_8, u1_u12_X_11, u1_u12_X_12, u1_u12_X_19, 
       u1_u12_X_2, u1_u12_X_20, u1_u12_X_23, u1_u12_X_25, u1_u12_X_29, u1_u12_X_30, u1_u12_X_31, u1_u12_X_32, u1_u12_X_41, 
       u1_u12_X_42, u1_u12_X_43, u1_u12_X_44, u1_u12_X_48, u1_u12_X_5, u1_u12_X_7, u1_u13_X_1, u1_u13_X_11, u1_u13_X_13, 
       u1_u13_X_17, u1_u13_X_18, u1_u13_X_19, u1_u13_X_2, u1_u13_X_20, u1_u13_X_23, u1_u13_X_24, u1_u13_X_25, u1_u13_X_26, 
       u1_u13_X_30, u1_u13_X_32, u1_u13_X_35, u1_u13_X_36, u1_u13_X_5, u1_u13_X_6, u1_u13_X_7, u1_u13_X_8, u1_u14_X_1, 
       u1_u14_X_11, u1_u14_X_13, u1_u14_X_2, u1_u14_X_23, u1_u14_X_24, u1_u14_X_25, u1_u14_X_26, u1_u14_X_29, u1_u14_X_30, 
       u1_u14_X_31, u1_u14_X_32, u1_u14_X_35, u1_u14_X_36, u1_u14_X_43, u1_u14_X_44, u1_u14_X_47, u1_u14_X_48, u1_u15_X_1, 
       u1_u15_X_11, u1_u15_X_12, u1_u15_X_13, u1_u15_X_14, u1_u15_X_17, u1_u15_X_18, u1_u15_X_19, u1_u15_X_2, u1_u15_X_20, 
       u1_u15_X_23, u1_u15_X_25, u1_u15_X_29, u1_u15_X_30, u1_u15_X_37, u1_u15_X_38, u1_u15_X_41, u1_u15_X_42, u1_u15_X_5, 
       u1_u15_X_7, u1_u1_X_19, u1_u1_X_2, u1_u1_X_20, u1_u1_X_23, u1_u1_X_24, u1_u1_X_25, u1_u1_X_26, u1_u1_X_29, 
       u1_u1_X_30, u1_u1_X_31, u1_u1_X_32, u1_u1_X_35, u1_u1_X_36, u1_u1_X_37, u1_u1_X_38, u1_u1_X_41, u1_u1_X_42, 
       u1_u1_X_43, u1_u1_X_44, u1_u1_X_48, u1_u1_X_5, u1_u1_X_6, u1_u2_X_1, u1_u2_X_11, u1_u2_X_12, u1_u2_X_13, 
       u1_u2_X_14, u1_u2_X_17, u1_u2_X_18, u1_u2_X_2, u1_u2_X_25, u1_u2_X_26, u1_u2_X_29, u1_u2_X_30, u1_u2_X_37, 
       u1_u2_X_38, u1_u2_X_41, u1_u2_X_42, u1_u2_X_6, u1_u2_X_8, u1_u3_X_11, u1_u3_X_12, u1_u3_X_13, u1_u3_X_14, 
       u1_u3_X_29, u1_u3_X_30, u1_u3_X_37, u1_u3_X_38, u1_u3_X_41, u1_u3_X_42, u1_u3_X_43, u1_u3_X_44, u1_u3_X_47, 
       u1_u3_X_48, u1_u3_X_7, u1_u3_X_8, u1_u4_X_11, u1_u4_X_12, u1_u4_X_13, u1_u4_X_14, u1_u4_X_17, u1_u4_X_19, 
       u1_u4_X_42, u1_u4_X_44, u1_u4_X_47, u1_u4_X_48, u1_u4_X_7, u1_u4_X_8, u1_u5_X_11, u1_u5_X_12, u1_u5_X_19, 
       u1_u5_X_20, u1_u5_X_23, u1_u5_X_24, u1_u5_X_31, u1_u5_X_32, u1_u5_X_5, u1_u5_X_7, u1_u6_X_1, u1_u6_X_2, 
       u1_u6_X_35, u1_u6_X_36, u1_u6_X_37, u1_u6_X_38, u1_u6_X_42, u1_u6_X_44, u1_u6_X_47, u1_u6_X_48, u1_u7_X_1, 
       u1_u7_X_17, u1_u7_X_19, u1_u7_X_2, u1_u7_X_24, u1_u7_X_26, u1_u7_X_29, u1_u7_X_30, u1_u7_X_43, u1_u7_X_44, 
       u1_u7_X_47, u1_u7_X_48, u1_u8_X_1, u1_u8_X_12, u1_u8_X_14, u1_u8_X_2, u1_u8_X_29, u1_u8_X_30, u1_u8_X_31, 
       u1_u8_X_32, u1_u8_X_41, u1_u8_X_42, u1_u8_X_5, u1_u8_X_6, u1_u8_X_7, u1_u8_X_8, u1_u9_X_11, u1_u9_X_12, 
       u1_u9_X_13, u1_u9_X_14, u1_u9_X_23, u1_u9_X_24, u1_u9_X_25, u1_u9_X_26, u1_u9_X_29, u1_u9_X_30, u1_u9_X_31, 
       u1_u9_X_32, u1_u9_X_35, u1_u9_X_36, u1_u9_X_43, u1_u9_X_44, u1_u9_X_47, u1_u9_X_48, u1_u9_X_7, u1_u9_X_8, 
       u1_uk_K_r0_11, u1_uk_K_r0_13, u1_uk_K_r0_15, u1_uk_K_r0_17, u1_uk_K_r0_19, u1_uk_K_r0_2, u1_uk_K_r0_22, u1_uk_K_r0_25, u1_uk_K_r0_28, 
       u1_uk_K_r0_31, u1_uk_K_r0_32, u1_uk_K_r0_34, u1_uk_K_r0_36, u1_uk_K_r0_47, u1_uk_K_r0_49, u1_uk_K_r0_52, u1_uk_K_r0_55, u1_uk_K_r0_7, 
       u1_uk_K_r10_10, u1_uk_K_r10_11, u1_uk_K_r10_14, u1_uk_K_r10_16, u1_uk_K_r10_18, u1_uk_K_r10_19, u1_uk_K_r10_23, u1_uk_K_r10_25, u1_uk_K_r10_27, 
       u1_uk_K_r10_28, u1_uk_K_r10_32, u1_uk_K_r10_34, u1_uk_K_r10_37, u1_uk_K_r10_39, u1_uk_K_r10_4, u1_uk_K_r10_41, u1_uk_K_r10_42, u1_uk_K_r10_43, 
       u1_uk_K_r10_44, u1_uk_K_r10_47, u1_uk_K_r10_48, u1_uk_K_r10_49, u1_uk_K_r10_52, u1_uk_K_r10_9, u1_uk_K_r11_10, u1_uk_K_r11_11, u1_uk_K_r11_17, 
       u1_uk_K_r11_19, u1_uk_K_r11_20, u1_uk_K_r11_21, u1_uk_K_r11_24, u1_uk_K_r11_25, u1_uk_K_r11_26, u1_uk_K_r11_27, u1_uk_K_r11_28, u1_uk_K_r11_29, 
       u1_uk_K_r11_33, u1_uk_K_r11_34, u1_uk_K_r11_39, u1_uk_K_r11_4, u1_uk_K_r11_46, u1_uk_K_r11_47, u1_uk_K_r11_48, u1_uk_K_r11_5, u1_uk_K_r11_53, 
       u1_uk_K_r11_54, u1_uk_K_r11_6, u1_uk_K_r11_7, u1_uk_K_r11_8, u1_uk_K_r12_1, u1_uk_K_r12_10, u1_uk_K_r12_15, u1_uk_K_r12_16, u1_uk_K_r12_18, 
       u1_uk_K_r12_21, u1_uk_K_r12_22, u1_uk_K_r12_25, u1_uk_K_r12_30, u1_uk_K_r12_33, u1_uk_K_r12_36, u1_uk_K_r12_41, u1_uk_K_r12_42, u1_uk_K_r12_44, 
       u1_uk_K_r12_47, u1_uk_K_r12_7, u1_uk_K_r13_0, u1_uk_K_r13_13, u1_uk_K_r13_17, u1_uk_K_r13_19, u1_uk_K_r13_2, u1_uk_K_r13_22, u1_uk_K_r13_23, 
       u1_uk_K_r13_25, u1_uk_K_r13_31, u1_uk_K_r13_32, u1_uk_K_r13_35, u1_uk_K_r13_36, u1_uk_K_r13_38, u1_uk_K_r13_4, u1_uk_K_r13_44, u1_uk_K_r13_55, 
       u1_uk_K_r14_10, u1_uk_K_r14_11, u1_uk_K_r14_12, u1_uk_K_r14_15, u1_uk_K_r14_16, u1_uk_K_r14_18, u1_uk_K_r14_2, u1_uk_K_r14_23, u1_uk_K_r14_3, 
       u1_uk_K_r14_38, u1_uk_K_r14_39, u1_uk_K_r14_42, u1_uk_K_r14_43, u1_uk_K_r14_45, u1_uk_K_r14_46, u1_uk_K_r14_5, u1_uk_K_r14_50, u1_uk_K_r14_8, 
       u1_uk_K_r14_9, u1_uk_K_r1_10, u1_uk_K_r1_15, u1_uk_K_r1_16, u1_uk_K_r1_17, u1_uk_K_r1_18, u1_uk_K_r1_21, u1_uk_K_r1_22, u1_uk_K_r1_33, 
       u1_uk_K_r1_36, u1_uk_K_r1_41, u1_uk_K_r1_42, u1_uk_K_r1_44, u1_uk_K_r1_47, u1_uk_K_r1_6, u1_uk_K_r1_7, u1_uk_K_r2_13, u1_uk_K_r2_16, 
       u1_uk_K_r2_18, u1_uk_K_r2_20, u1_uk_K_r2_21, u1_uk_K_r2_24, u1_uk_K_r2_25, u1_uk_K_r2_26, u1_uk_K_r2_27, u1_uk_K_r2_28, u1_uk_K_r2_29, 
       u1_uk_K_r2_31, u1_uk_K_r2_33, u1_uk_K_r2_36, u1_uk_K_r2_4, u1_uk_K_r2_41, u1_uk_K_r2_46, u1_uk_K_r2_47, u1_uk_K_r2_49, u1_uk_K_r2_50, 
       u1_uk_K_r2_53, u1_uk_K_r2_55, u1_uk_K_r2_6, u1_uk_K_r2_7, u1_uk_K_r3_10, u1_uk_K_r3_11, u1_uk_K_r3_14, u1_uk_K_r3_15, u1_uk_K_r3_16, 
       u1_uk_K_r3_19, u1_uk_K_r3_24, u1_uk_K_r3_29, u1_uk_K_r3_33, u1_uk_K_r3_34, u1_uk_K_r3_35, u1_uk_K_r3_38, u1_uk_K_r3_4, u1_uk_K_r3_43, 
       u1_uk_K_r3_44, u1_uk_K_r3_47, u1_uk_K_r3_51, u1_uk_K_r3_52, u1_uk_K_r3_9, u1_uk_K_r4_0, u1_uk_K_r4_11, u1_uk_K_r4_17, u1_uk_K_r4_18, 
       u1_uk_K_r4_23, u1_uk_K_r4_27, u1_uk_K_r4_3, u1_uk_K_r4_31, u1_uk_K_r4_33, u1_uk_K_r4_35, u1_uk_K_r4_38, u1_uk_K_r4_4, u1_uk_K_r4_41, 
       u1_uk_K_r4_47, u1_uk_K_r4_48, u1_uk_K_r4_49, u1_uk_K_r4_5, u1_uk_K_r4_54, u1_uk_K_r4_55, u1_uk_K_r5_0, u1_uk_K_r5_1, u1_uk_K_r5_10, 
       u1_uk_K_r5_13, u1_uk_K_r5_16, u1_uk_K_r5_17, u1_uk_K_r5_18, u1_uk_K_r5_19, u1_uk_K_r5_21, u1_uk_K_r5_23, u1_uk_K_r5_26, u1_uk_K_r5_31, 
       u1_uk_K_r5_32, u1_uk_K_r5_35, u1_uk_K_r5_36, u1_uk_K_r5_37, u1_uk_K_r5_39, u1_uk_K_r5_4, u1_uk_K_r5_40, u1_uk_K_r5_41, u1_uk_K_r5_43, 
       u1_uk_K_r5_48, u1_uk_K_r5_5, u1_uk_K_r5_51, u1_uk_K_r5_53, u1_uk_K_r5_7, u1_uk_K_r5_8, u1_uk_K_r6_0, u1_uk_K_r6_10, u1_uk_K_r6_14, 
       u1_uk_K_r6_17, u1_uk_K_r6_19, u1_uk_K_r6_21, u1_uk_K_r6_22, u1_uk_K_r6_26, u1_uk_K_r6_27, u1_uk_K_r6_28, u1_uk_K_r6_29, u1_uk_K_r6_3, 
       u1_uk_K_r6_30, u1_uk_K_r6_31, u1_uk_K_r6_34, u1_uk_K_r6_35, u1_uk_K_r6_37, u1_uk_K_r6_46, u1_uk_K_r6_51, u1_uk_K_r6_53, u1_uk_K_r6_55, 
       u1_uk_K_r6_7, u1_uk_K_r7_0, u1_uk_K_r7_1, u1_uk_K_r7_13, u1_uk_K_r7_15, u1_uk_K_r7_16, u1_uk_K_r7_2, u1_uk_K_r7_20, u1_uk_K_r7_22, 
       u1_uk_K_r7_23, u1_uk_K_r7_24, u1_uk_K_r7_25, u1_uk_K_r7_26, u1_uk_K_r7_27, u1_uk_K_r7_29, u1_uk_K_r7_30, u1_uk_K_r7_31, u1_uk_K_r7_32, 
       u1_uk_K_r7_34, u1_uk_K_r7_37, u1_uk_K_r7_39, u1_uk_K_r7_41, u1_uk_K_r7_46, u1_uk_K_r7_48, u1_uk_K_r7_5, u1_uk_K_r7_53, u1_uk_K_r7_55, 
       u1_uk_K_r7_6, u1_uk_K_r7_7, u1_uk_K_r7_8, u1_uk_K_r7_9, u1_uk_K_r8_10, u1_uk_K_r8_13, u1_uk_K_r8_16, u1_uk_K_r8_17, u1_uk_K_r8_19, 
       u1_uk_K_r8_2, u1_uk_K_r8_21, u1_uk_K_r8_22, u1_uk_K_r8_27, u1_uk_K_r8_28, u1_uk_K_r8_32, u1_uk_K_r8_37, u1_uk_K_r8_39, u1_uk_K_r8_40, 
       u1_uk_K_r8_41, u1_uk_K_r8_42, u1_uk_K_r8_43, u1_uk_K_r8_44, u1_uk_K_r8_48, u1_uk_K_r8_5, u1_uk_K_r8_51, u1_uk_K_r8_52, u1_uk_K_r8_8, 
       u1_uk_K_r9_0, u1_uk_K_r9_1, u1_uk_K_r9_10, u1_uk_K_r9_12, u1_uk_K_r9_13, u1_uk_K_r9_15, u1_uk_K_r9_18, u1_uk_K_r9_19, u1_uk_K_r9_22, 
       u1_uk_K_r9_23, u1_uk_K_r9_25, u1_uk_K_r9_27, u1_uk_K_r9_30, u1_uk_K_r9_31, u1_uk_K_r9_33, u1_uk_K_r9_35, u1_uk_K_r9_38, u1_uk_K_r9_4, 
       u1_uk_K_r9_45, u1_uk_K_r9_48, u1_uk_K_r9_49, u1_uk_K_r9_5, u1_uk_K_r9_54, u1_uk_K_r9_55, u1_uk_K_r9_6, u1_uk_K_r9_7, u1_uk_K_r9_9, 
       u1_uk_n1004, u1_uk_n1011, u1_uk_n1015, u1_uk_n1016, u1_uk_n1017, u1_uk_n1027, u1_uk_n1028, u1_uk_n1050, u1_uk_n1054, 
       u1_uk_n1056, u1_uk_n1057, u1_uk_n1058, u1_uk_n1073, u1_uk_n1074, u1_uk_n1076, u1_uk_n1079, u1_uk_n1080, u1_uk_n1083, 
       u1_uk_n1088, u1_uk_n1092, u1_uk_n1096, u1_uk_n1101, u1_uk_n1104, u1_uk_n1105, u1_uk_n1106, u1_uk_n1109, u1_uk_n1113, 
       u1_uk_n1114, u1_uk_n1115, u1_uk_n1118, u1_uk_n1119, u1_uk_n1124, u1_uk_n1125, u1_uk_n1126, u1_uk_n1128, u1_uk_n1130, 
       u1_uk_n1140, u1_uk_n1147, u1_uk_n1148, u1_uk_n1153, u1_uk_n1154, u1_uk_n1156, u1_uk_n1157, u1_uk_n1158, u1_uk_n1159, 
       u1_uk_n1162, u1_uk_n1163, u1_uk_n1171, u1_uk_n1218, u1_uk_n1219, u1_uk_n1220, u1_uk_n1221, u1_uk_n1222, u1_uk_n1224, 
       u1_uk_n1225, u1_uk_n1227, u1_uk_n1228, u1_uk_n1229, u1_uk_n1230, u1_uk_n1231, u1_uk_n1233, u1_uk_n1234, u1_uk_n1235, 
       u1_uk_n1236, u1_uk_n1237, u1_uk_n1238, u1_uk_n1239, u1_uk_n1240, u1_uk_n1241, u1_uk_n1242, u1_uk_n1243, u1_uk_n1244, 
       u1_uk_n1245, u1_uk_n1246, u1_uk_n1247, u1_uk_n1248, u1_uk_n1249, u1_uk_n1250, u1_uk_n1251, u1_uk_n1252, u1_uk_n1253, 
       u1_uk_n1255, u1_uk_n1256, u1_uk_n1257, u1_uk_n1258, u1_uk_n1259, u1_uk_n1260, u1_uk_n1261, u1_uk_n1262, u1_uk_n1263, 
       u1_uk_n1264, u1_uk_n1265, u1_uk_n1266, u1_uk_n1267, u1_uk_n1268, u1_uk_n1269, u1_uk_n1270, u1_uk_n1271, u1_uk_n1272, 
       u1_uk_n1273, u1_uk_n1274, u1_uk_n1275, u1_uk_n1276, u1_uk_n1277, u1_uk_n1278, u1_uk_n1279, u1_uk_n1281, u1_uk_n1282, 
       u1_uk_n1284, u1_uk_n1286, u1_uk_n1288, u1_uk_n1289, u1_uk_n1290, u1_uk_n1291, u1_uk_n1292, u1_uk_n1293, u1_uk_n1294, 
       u1_uk_n1295, u1_uk_n1296, u1_uk_n1297, u1_uk_n1299, u1_uk_n1300, u1_uk_n1303, u1_uk_n1304, u1_uk_n1305, u1_uk_n1307, 
       u1_uk_n1308, u1_uk_n1309, u1_uk_n1310, u1_uk_n1311, u1_uk_n1312, u1_uk_n1313, u1_uk_n1314, u1_uk_n1315, u1_uk_n1316, 
       u1_uk_n1317, u1_uk_n1318, u1_uk_n1319, u1_uk_n1320, u1_uk_n1321, u1_uk_n1322, u1_uk_n1323, u1_uk_n1324, u1_uk_n1325, 
       u1_uk_n1326, u1_uk_n1327, u1_uk_n1328, u1_uk_n1329, u1_uk_n1330, u1_uk_n1331, u1_uk_n1332, u1_uk_n1333, u1_uk_n1334, 
       u1_uk_n1335, u1_uk_n1336, u1_uk_n1338, u1_uk_n1339, u1_uk_n1340, u1_uk_n1341, u1_uk_n1342, u1_uk_n1343, u1_uk_n1344, 
       u1_uk_n1345, u1_uk_n1346, u1_uk_n1347, u1_uk_n1348, u1_uk_n1349, u1_uk_n1350, u1_uk_n1351, u1_uk_n1352, u1_uk_n1353, 
       u1_uk_n1354, u1_uk_n1355, u1_uk_n1356, u1_uk_n1357, u1_uk_n1358, u1_uk_n1359, u1_uk_n1360, u1_uk_n1361, u1_uk_n1363, 
       u1_uk_n1365, u1_uk_n1366, u1_uk_n1367, u1_uk_n1369, u1_uk_n1371, u1_uk_n1372, u1_uk_n1374, u1_uk_n1375, u1_uk_n1376, 
       u1_uk_n1377, u1_uk_n1378, u1_uk_n1380, u1_uk_n1381, u1_uk_n1382, u1_uk_n1383, u1_uk_n1386, u1_uk_n1389, u1_uk_n1390, 
       u1_uk_n1391, u1_uk_n1393, u1_uk_n1394, u1_uk_n1395, u1_uk_n1396, u1_uk_n1397, u1_uk_n1398, u1_uk_n1399, u1_uk_n1400, 
       u1_uk_n1401, u1_uk_n1402, u1_uk_n1403, u1_uk_n1404, u1_uk_n1405, u1_uk_n1406, u1_uk_n1407, u1_uk_n1408, u1_uk_n1409, 
       u1_uk_n1410, u1_uk_n1411, u1_uk_n1412, u1_uk_n1413, u1_uk_n1414, u1_uk_n1415, u1_uk_n1417, u1_uk_n1418, u1_uk_n1419, 
       u1_uk_n1422, u1_uk_n1423, u1_uk_n1424, u1_uk_n1425, u1_uk_n1426, u1_uk_n1427, u1_uk_n1429, u1_uk_n1430, u1_uk_n1431, 
       u1_uk_n1433, u1_uk_n1435, u1_uk_n1436, u1_uk_n1437, u1_uk_n1438, u1_uk_n1439, u1_uk_n1440, u1_uk_n1441, u1_uk_n1442, 
       u1_uk_n1443, u1_uk_n1444, u1_uk_n1446, u1_uk_n1447, u1_uk_n1448, u1_uk_n1449, u1_uk_n1450, u1_uk_n1452, u1_uk_n1453, 
       u1_uk_n1454, u1_uk_n1455, u1_uk_n1456, u1_uk_n1457, u1_uk_n1458, u1_uk_n1459, u1_uk_n1460, u1_uk_n1461, u1_uk_n1462, 
       u1_uk_n1463, u1_uk_n1464, u1_uk_n1465, u1_uk_n1466, u1_uk_n1468, u1_uk_n1469, u1_uk_n1470, u1_uk_n1471, u1_uk_n1472, 
       u1_uk_n1474, u1_uk_n1475, u1_uk_n1476, u1_uk_n1477, u1_uk_n1478, u1_uk_n1482, u1_uk_n1483, u1_uk_n1484, u1_uk_n1485, 
       u1_uk_n1486, u1_uk_n1487, u1_uk_n1488, u1_uk_n1489, u1_uk_n1490, u1_uk_n1491, u1_uk_n1492, u1_uk_n1494, u1_uk_n1495, 
       u1_uk_n1496, u1_uk_n1498, u1_uk_n1499, u1_uk_n1500, u1_uk_n1501, u1_uk_n1504, u1_uk_n1505, u1_uk_n1507, u1_uk_n1508, 
       u1_uk_n1510, u1_uk_n1514, u1_uk_n1516, u1_uk_n1517, u1_uk_n1518, u1_uk_n1520, u1_uk_n1521, u1_uk_n1523, u1_uk_n1524, 
       u1_uk_n1526, u1_uk_n1527, u1_uk_n1528, u1_uk_n1529, u1_uk_n1530, u1_uk_n1531, u1_uk_n1532, u1_uk_n1533, u1_uk_n1534, 
       u1_uk_n1536, u1_uk_n1537, u1_uk_n1538, u1_uk_n1540, u1_uk_n1541, u1_uk_n1543, u1_uk_n1544, u1_uk_n1545, u1_uk_n1547, 
       u1_uk_n1548, u1_uk_n1549, u1_uk_n1551, u1_uk_n1552, u1_uk_n1554, u1_uk_n1555, u1_uk_n1556, u1_uk_n1557, u1_uk_n1558, 
       u1_uk_n1559, u1_uk_n1560, u1_uk_n1561, u1_uk_n1562, u1_uk_n1563, u1_uk_n1564, u1_uk_n1565, u1_uk_n1566, u1_uk_n1567, 
       u1_uk_n1568, u1_uk_n1570, u1_uk_n1571, u1_uk_n1572, u1_uk_n1573, u1_uk_n1574, u1_uk_n1577, u1_uk_n1578, u1_uk_n1579, 
       u1_uk_n1581, u1_uk_n1584, u1_uk_n1585, u1_uk_n1586, u1_uk_n1588, u1_uk_n1592, u1_uk_n1593, u1_uk_n1595, u1_uk_n1598, 
       u1_uk_n1599, u1_uk_n1600, u1_uk_n1601, u1_uk_n1603, u1_uk_n1604, u1_uk_n1605, u1_uk_n1606, u1_uk_n1607, u1_uk_n1608, 
       u1_uk_n1610, u1_uk_n1612, u1_uk_n1613, u1_uk_n1614, u1_uk_n1615, u1_uk_n1616, u1_uk_n1618, u1_uk_n1619, u1_uk_n1620, 
       u1_uk_n1621, u1_uk_n1622, u1_uk_n1623, u1_uk_n1624, u1_uk_n1625, u1_uk_n1626, u1_uk_n1627, u1_uk_n1628, u1_uk_n1629, 
       u1_uk_n1630, u1_uk_n1632, u1_uk_n1633, u1_uk_n1634, u1_uk_n1635, u1_uk_n1639, u1_uk_n1640, u1_uk_n1641, u1_uk_n1642, 
       u1_uk_n1643, u1_uk_n1644, u1_uk_n1645, u1_uk_n1647, u1_uk_n1649, u1_uk_n1651, u1_uk_n1652, u1_uk_n1653, u1_uk_n1654, 
       u1_uk_n1655, u1_uk_n1656, u1_uk_n1659, u1_uk_n1660, u1_uk_n1661, u1_uk_n1662, u1_uk_n1663, u1_uk_n1664, u1_uk_n1667, 
       u1_uk_n1669, u1_uk_n1670, u1_uk_n1672, u1_uk_n1673, u1_uk_n1676, u1_uk_n1677, u1_uk_n1678, u1_uk_n1682, u1_uk_n1683, 
       u1_uk_n1684, u1_uk_n1687, u1_uk_n1688, u1_uk_n1689, u1_uk_n1690, u1_uk_n1691, u1_uk_n1692, u1_uk_n1693, u1_uk_n1694, 
       u1_uk_n1695, u1_uk_n1696, u1_uk_n1698, u1_uk_n1699, u1_uk_n1702, u1_uk_n1703, u1_uk_n1704, u1_uk_n1705, u1_uk_n1707, 
       u1_uk_n1708, u1_uk_n1709, u1_uk_n1710, u1_uk_n1711, u1_uk_n1712, u1_uk_n1713, u1_uk_n1714, u1_uk_n1715, u1_uk_n1716, 
       u1_uk_n1717, u1_uk_n1718, u1_uk_n1719, u1_uk_n1720, u1_uk_n1721, u1_uk_n1722, u1_uk_n1723, u1_uk_n1728, u1_uk_n1729, 
       u1_uk_n1730, u1_uk_n1731, u1_uk_n1732, u1_uk_n1734, u1_uk_n1735, u1_uk_n1736, u1_uk_n1737, u1_uk_n1738, u1_uk_n1739, 
       u1_uk_n1744, u1_uk_n1745, u1_uk_n1748, u1_uk_n1749, u1_uk_n1750, u1_uk_n1751, u1_uk_n1752, u1_uk_n1753, u1_uk_n1754, 
       u1_uk_n1755, u1_uk_n1756, u1_uk_n1757, u1_uk_n1758, u1_uk_n1761, u1_uk_n1762, u1_uk_n1763, u1_uk_n1764, u1_uk_n1765, 
       u1_uk_n1766, u1_uk_n1767, u1_uk_n1768, u1_uk_n1769, u1_uk_n1772, u1_uk_n1773, u1_uk_n1774, u1_uk_n1775, u1_uk_n1776, 
       u1_uk_n1777, u1_uk_n1780, u1_uk_n1781, u1_uk_n1782, u1_uk_n1783, u1_uk_n1784, u1_uk_n1785, u1_uk_n1787, u1_uk_n1790, 
       u1_uk_n1791, u1_uk_n1792, u1_uk_n1793, u1_uk_n1797, u1_uk_n1798, u1_uk_n1799, u1_uk_n1800, u1_uk_n1801, u1_uk_n1802, 
       u1_uk_n1803, u1_uk_n1804, u1_uk_n1806, u1_uk_n1807, u1_uk_n1808, u1_uk_n1809, u1_uk_n1810, u1_uk_n1811, u1_uk_n1812, 
       u1_uk_n1813, u1_uk_n1814, u1_uk_n1815, u1_uk_n1816, u1_uk_n1817, u1_uk_n1818, u1_uk_n1819, u1_uk_n1820, u1_uk_n1821, 
       u1_uk_n1822, u1_uk_n1823, u1_uk_n1824, u1_uk_n1826, u1_uk_n1827, u1_uk_n1829, u1_uk_n1830, u1_uk_n1831, u1_uk_n1832, 
       u1_uk_n1833, u1_uk_n1834, u1_uk_n1835, u1_uk_n1836, u1_uk_n1837, u1_uk_n1838, u1_uk_n1839, u1_uk_n1840, u1_uk_n1841, 
       u1_uk_n1842, u1_uk_n1843, u1_uk_n1844, u1_uk_n1845, u1_uk_n1846, u1_uk_n1847, u1_uk_n1848, u1_uk_n1849, u1_uk_n1850, 
       u1_uk_n1851, u1_uk_n1852, u1_uk_n1853, u1_uk_n1854, u1_uk_n1855, u1_uk_n1856, u1_uk_n1858, u1_uk_n1859, u1_uk_n1860, 
       u1_uk_n1862, u1_uk_n1863, u1_uk_n1864, u1_uk_n1865, u1_uk_n1866, u1_uk_n1867, u1_uk_n1868, u1_uk_n1869, u1_uk_n1870, 
       u1_uk_n1872, u1_uk_n1873, u1_uk_n1874, u1_uk_n1875, u1_uk_n1876, u1_uk_n1879, u1_uk_n1880, u1_uk_n1881, u1_uk_n1882, 
       u1_uk_n1883, u1_uk_n1884, u1_uk_n1885, u1_uk_n1886, u1_uk_n1887, u1_uk_n312, u1_uk_n349, u1_uk_n376, u1_uk_n379, 
       u1_uk_n382, u1_uk_n468, u1_uk_n472, u1_uk_n501, u1_uk_n504, u1_uk_n601, u1_uk_n656, u1_uk_n671, u1_uk_n689, 
       u1_uk_n692, u1_uk_n949, u1_uk_n955, u1_uk_n976, u1_uk_n996, u2_FP_11, u2_FP_12, u2_FP_15, u2_FP_19, 
       u2_FP_21, u2_FP_22, u2_FP_27, u2_FP_29, u2_FP_32, u2_FP_33, u2_FP_34, u2_FP_35, u2_FP_36, 
       u2_FP_37, u2_FP_4, u2_FP_40, u2_FP_41, u2_FP_42, u2_FP_44, u2_FP_46, u2_FP_47, u2_FP_48, 
       u2_FP_49, u2_FP_5, u2_FP_51, u2_FP_52, u2_FP_53, u2_FP_54, u2_FP_55, u2_FP_56, u2_FP_57, 
       u2_FP_58, u2_FP_59, u2_FP_60, u2_FP_61, u2_FP_62, u2_FP_63, u2_FP_64, u2_FP_7, u2_K10_11, 
       u2_K10_17, u2_K10_19, u2_K10_25, u2_K10_26, u2_K10_29, u2_K10_36, u2_K10_42, u2_K10_43, u2_K10_44, 
       u2_K10_5, u2_K10_6, u2_K11_11, u2_K11_13, u2_K11_18, u2_K11_29, u2_K11_37, u2_K11_38, u2_K11_42, 
       u2_K11_45, u2_K11_48, u2_K11_6, u2_K11_7, u2_K12_2, u2_K12_20, u2_K12_22, u2_K12_24, u2_K12_25, 
       u2_K12_26, u2_K12_41, u2_K12_46, u2_K12_47, u2_K12_48, u2_K12_8, u2_K13_14, u2_K13_20, u2_K13_25, 
       u2_K13_26, u2_K13_3, u2_K13_31, u2_K13_32, u2_K13_34, u2_K13_37, u2_K13_40, u2_K13_42, u2_K13_44, 
       u2_K13_45, u2_K13_46, u2_K13_47, u2_K13_8, u2_K14_10, u2_K14_11, u2_K14_12, u2_K14_13, u2_K14_14, 
       u2_K14_16, u2_K14_17, u2_K14_18, u2_K14_3, u2_K14_42, u2_K14_43, u2_K14_48, u2_K14_6, u2_K14_8, 
       u2_K15_1, u2_K15_13, u2_K15_16, u2_K15_18, u2_K15_2, u2_K15_20, u2_K15_29, u2_K15_31, u2_K15_35, 
       u2_K15_37, u2_K15_44, u2_K15_47, u2_K15_48, u2_K15_5, u2_K16_26, u2_K16_31, u2_K16_42, u2_K16_44, 
       u2_K16_47, u2_K16_5, u2_K16_6, u2_K16_8, u2_K1_19, u2_K1_24, u2_K1_30, u2_K1_37, u2_K1_43, 
       u2_K2_1, u2_K2_12, u2_K2_18, u2_K2_20, u2_K2_29, u2_K2_36, u2_K2_43, u2_K2_47, u2_K2_48, 
       u2_K3_13, u2_K3_19, u2_K3_23, u2_K3_26, u2_K3_35, u2_K3_48, u2_K4_13, u2_K4_14, u2_K4_18, 
       u2_K4_19, u2_K4_35, u2_K5_11, u2_K5_13, u2_K5_14, u2_K5_17, u2_K5_18, u2_K5_19, u2_K5_2, 
       u2_K5_29, u2_K5_30, u2_K5_31, u2_K5_32, u2_K5_41, u2_K5_44, u2_K5_48, u2_K5_5, u2_K5_6, 
       u2_K5_8, u2_K6_11, u2_K6_13, u2_K6_19, u2_K6_20, u2_K6_23, u2_K6_24, u2_K6_25, u2_K6_36, 
       u2_K6_48, u2_K6_5, u2_K6_6, u2_K6_8, u2_K7_26, u2_K7_35, u2_K7_37, u2_K7_38, u2_K7_43, 
       u2_K7_44, u2_K7_48, u2_K7_5, u2_K7_7, u2_K8_13, u2_K8_18, u2_K8_24, u2_K8_26, u2_K8_31, 
       u2_K8_41, u2_K8_42, u2_K8_45, u2_K8_5, u2_K8_8, u2_K9_12, u2_K9_14, u2_K9_23, u2_K9_25, 
       u2_K9_29, u2_K9_3, u2_K9_32, u2_K9_36, u2_K9_38, u2_K9_40, u2_K9_45, u2_K9_5, u2_L10_1, 
       u2_L10_10, u2_L10_15, u2_L10_16, u2_L10_17, u2_L10_20, u2_L10_21, u2_L10_23, u2_L10_24, u2_L10_26, 
       u2_L10_27, u2_L10_30, u2_L10_31, u2_L10_5, u2_L10_6, u2_L10_9, u2_L11_1, u2_L11_10, u2_L11_11, 
       u2_L11_12, u2_L11_13, u2_L11_14, u2_L11_15, u2_L11_16, u2_L11_17, u2_L11_18, u2_L11_19, u2_L11_2, 
       u2_L11_20, u2_L11_21, u2_L11_22, u2_L11_23, u2_L11_24, u2_L11_25, u2_L11_26, u2_L11_3, u2_L11_30, 
       u2_L11_31, u2_L11_32, u2_L11_4, u2_L11_5, u2_L11_6, u2_L11_7, u2_L11_8, u2_L11_9, u2_L12_13, 
       u2_L12_15, u2_L12_16, u2_L12_17, u2_L12_18, u2_L12_2, u2_L12_21, u2_L12_23, u2_L12_24, u2_L12_27, 
       u2_L12_28, u2_L12_30, u2_L12_31, u2_L12_5, u2_L12_6, u2_L12_9, u2_L13_13, u2_L13_16, u2_L13_18, 
       u2_L13_2, u2_L13_24, u2_L13_28, u2_L13_30, u2_L13_6, u2_L14_11, u2_L14_12, u2_L14_15, u2_L14_19, 
       u2_L14_21, u2_L14_22, u2_L14_27, u2_L14_29, u2_L14_32, u2_L14_4, u2_L14_5, u2_L14_7, u2_L6_11, 
       u2_L6_14, u2_L6_15, u2_L6_19, u2_L6_21, u2_L6_22, u2_L6_25, u2_L6_27, u2_L6_29, u2_L6_3, 
       u2_L6_32, u2_L6_4, u2_L6_5, u2_L6_7, u2_L6_8, u2_L7_11, u2_L7_12, u2_L7_15, u2_L7_17, 
       u2_L7_19, u2_L7_21, u2_L7_22, u2_L7_23, u2_L7_27, u2_L7_29, u2_L7_31, u2_L7_32, u2_L7_4, 
       u2_L7_5, u2_L7_7, u2_L7_9, u2_L9_12, u2_L9_14, u2_L9_15, u2_L9_21, u2_L9_22, u2_L9_25, 
       u2_L9_27, u2_L9_3, u2_L9_32, u2_L9_5, u2_L9_7, u2_L9_8, u2_N226, u2_N227, u2_N228, 
       u2_N230, u2_N231, u2_N234, u2_N237, u2_N238, u2_N242, u2_N244, u2_N245, u2_N248, 
       u2_N250, u2_N252, u2_N255, u2_N259, u2_N260, u2_N262, u2_N264, u2_N266, u2_N267, 
       u2_N270, u2_N272, u2_N274, u2_N276, u2_N277, u2_N278, u2_N282, u2_N284, u2_N286, 
       u2_N287, u2_N322, u2_N324, u2_N326, u2_N327, u2_N331, u2_N333, u2_N334, u2_N340, 
       u2_N341, u2_N344, u2_N346, u2_N351, u2_N352, u2_N356, u2_N357, u2_N360, u2_N361, 
       u2_N366, u2_N367, u2_N368, u2_N371, u2_N372, u2_N374, u2_N375, u2_N377, u2_N378, 
       u2_N381, u2_N382, u2_N384, u2_N385, u2_N386, u2_N387, u2_N388, u2_N389, u2_N390, 
       u2_N391, u2_N392, u2_N393, u2_N394, u2_N395, u2_N396, u2_N397, u2_N398, u2_N399, 
       u2_N400, u2_N401, u2_N402, u2_N403, u2_N404, u2_N405, u2_N406, u2_N407, u2_N408, 
       u2_N409, u2_N413, u2_N414, u2_N415, u2_N417, u2_N420, u2_N421, u2_N424, u2_N428, 
       u2_N430, u2_N431, u2_N432, u2_N433, u2_N436, u2_N438, u2_N439, u2_N442, u2_N443, 
       u2_N445, u2_N446, u2_N449, u2_N453, u2_N460, u2_N463, u2_N465, u2_N471, u2_N475, 
       u2_N477, u2_R0_1, u2_R0_10, u2_R0_12, u2_R0_13, u2_R0_14, u2_R0_15, u2_R0_17, u2_R0_18, 
       u2_R0_19, u2_R0_20, u2_R0_21, u2_R0_25, u2_R0_28, u2_R0_3, u2_R0_32, u2_R0_4, u2_R0_5, 
       u2_R0_6, u2_R0_7, u2_R0_8, u2_R0_9, u2_R10_1, u2_R10_10, u2_R10_11, u2_R10_12, u2_R10_13, 
       u2_R10_14, u2_R10_15, u2_R10_16, u2_R10_17, u2_R10_19, u2_R10_2, u2_R10_21, u2_R10_28, u2_R10_29, 
       u2_R10_3, u2_R10_30, u2_R10_31, u2_R10_32, u2_R10_4, u2_R10_5, u2_R10_7, u2_R10_8, u2_R10_9, 
       u2_R11_1, u2_R11_10, u2_R11_11, u2_R11_12, u2_R11_13, u2_R11_14, u2_R11_15, u2_R11_16, u2_R11_17, 
       u2_R11_18, u2_R11_19, u2_R11_2, u2_R11_20, u2_R11_21, u2_R11_22, u2_R11_23, u2_R11_24, u2_R11_25, 
       u2_R11_26, u2_R11_27, u2_R11_28, u2_R11_29, u2_R11_3, u2_R11_30, u2_R11_31, u2_R11_32, u2_R11_4, 
       u2_R11_5, u2_R11_6, u2_R11_7, u2_R11_8, u2_R11_9, u2_R12_1, u2_R12_10, u2_R12_11, u2_R12_12, 
       u2_R12_13, u2_R12_17, u2_R12_18, u2_R12_2, u2_R12_20, u2_R12_21, u2_R12_22, u2_R12_23, u2_R12_24, 
       u2_R12_25, u2_R12_27, u2_R12_28, u2_R12_29, u2_R12_3, u2_R12_30, u2_R12_31, u2_R12_32, u2_R12_4, 
       u2_R12_5, u2_R12_6, u2_R12_7, u2_R12_8, u2_R12_9, u2_R13_1, u2_R13_10, u2_R13_11, u2_R13_12, 
       u2_R13_13, u2_R13_17, u2_R13_18, u2_R13_20, u2_R13_22, u2_R13_24, u2_R13_25, u2_R13_27, u2_R13_28, 
       u2_R13_29, u2_R13_30, u2_R13_32, u2_R13_4, u2_R13_5, u2_R13_6, u2_R13_7, u2_R13_8, u2_R13_9, 
       u2_R1_1, u2_R1_12, u2_R1_16, u2_R1_17, u2_R1_19, u2_R1_20, u2_R1_22, u2_R1_24, u2_R1_25, 
       u2_R1_27, u2_R1_3, u2_R1_30, u2_R1_5, u2_R1_8, u2_R1_9, u2_R2_1, u2_R2_11, u2_R2_12, 
       u2_R2_13, u2_R2_16, u2_R2_17, u2_R2_2, u2_R2_20, u2_R2_21, u2_R2_24, u2_R2_28, u2_R2_3, 
       u2_R2_32, u2_R2_6, u2_R2_7, u2_R2_8, u2_R2_9, u2_R3_1, u2_R3_12, u2_R3_13, u2_R3_15, 
       u2_R3_18, u2_R3_20, u2_R3_21, u2_R3_24, u2_R3_28, u2_R3_29, u2_R3_3, u2_R3_30, u2_R3_4, 
       u2_R3_5, u2_R3_8, u2_R3_9, u2_R4_1, u2_R4_12, u2_R4_13, u2_R4_14, u2_R4_16, u2_R4_17, 
       u2_R4_19, u2_R4_20, u2_R4_24, u2_R4_25, u2_R4_26, u2_R4_28, u2_R4_29, u2_R4_4, u2_R4_5, 
       u2_R4_6, u2_R4_7, u2_R4_8, u2_R5_1, u2_R5_10, u2_R5_11, u2_R5_12, u2_R5_13, u2_R5_14, 
       u2_R5_16, u2_R5_17, u2_R5_18, u2_R5_21, u2_R5_23, u2_R5_24, u2_R5_25, u2_R5_26, u2_R5_28, 
       u2_R5_29, u2_R5_32, u2_R5_4, u2_R5_5, u2_R5_8, u2_R5_9, u2_R6_1, u2_R6_10, u2_R6_11, 
       u2_R6_12, u2_R6_13, u2_R6_15, u2_R6_16, u2_R6_17, u2_R6_18, u2_R6_19, u2_R6_2, u2_R6_20, 
       u2_R6_21, u2_R6_22, u2_R6_23, u2_R6_24, u2_R6_25, u2_R6_26, u2_R6_27, u2_R6_28, u2_R6_29, 
       u2_R6_30, u2_R6_31, u2_R6_32, u2_R6_4, u2_R6_5, u2_R6_6, u2_R6_7, u2_R6_8, u2_R6_9, 
       u2_R7_1, u2_R7_11, u2_R7_12, u2_R7_13, u2_R7_14, u2_R7_15, u2_R7_16, u2_R7_17, u2_R7_2, 
       u2_R7_20, u2_R7_21, u2_R7_22, u2_R7_23, u2_R7_24, u2_R7_25, u2_R7_26, u2_R7_27, u2_R7_28, 
       u2_R7_29, u2_R7_3, u2_R7_30, u2_R7_31, u2_R7_32, u2_R7_4, u2_R7_5, u2_R7_6, u2_R7_7, 
       u2_R7_8, u2_R7_9, u2_R8_1, u2_R8_12, u2_R8_13, u2_R8_15, u2_R8_16, u2_R8_17, u2_R8_18, 
       u2_R8_19, u2_R8_20, u2_R8_22, u2_R8_24, u2_R8_25, u2_R8_26, u2_R8_27, u2_R8_28, u2_R8_29, 
       u2_R8_32, u2_R8_4, u2_R8_5, u2_R8_6, u2_R8_8, u2_R8_9, u2_R9_1, u2_R9_12, u2_R9_13, 
       u2_R9_15, u2_R9_16, u2_R9_17, u2_R9_18, u2_R9_19, u2_R9_2, u2_R9_20, u2_R9_21, u2_R9_24, 
       u2_R9_25, u2_R9_26, u2_R9_27, u2_R9_28, u2_R9_29, u2_R9_30, u2_R9_31, u2_R9_32, u2_R9_4, 
       u2_R9_5, u2_R9_8, u2_R9_9, u2_desIn_r_1, u2_desIn_r_11, u2_desIn_r_15, u2_desIn_r_23, u2_desIn_r_25, u2_desIn_r_27, 
       u2_desIn_r_29, u2_desIn_r_3, u2_desIn_r_33, u2_desIn_r_35, u2_desIn_r_37, u2_desIn_r_39, u2_desIn_r_43, u2_desIn_r_45, u2_desIn_r_5, 
       u2_desIn_r_53, u2_desIn_r_55, u2_desIn_r_57, u2_desIn_r_59, u2_desIn_r_61, u2_desIn_r_63, u2_desIn_r_7, u2_desIn_r_9, u2_key_r_0, 
       u2_key_r_10, u2_key_r_11, u2_key_r_12, u2_key_r_14, u2_key_r_16, u2_key_r_17, u2_key_r_19, u2_key_r_21, u2_key_r_22, 
       u2_key_r_23, u2_key_r_24, u2_key_r_25, u2_key_r_26, u2_key_r_28, u2_key_r_29, u2_key_r_3, u2_key_r_30, u2_key_r_31, 
       u2_key_r_32, u2_key_r_33, u2_key_r_34, u2_key_r_35, u2_key_r_36, u2_key_r_37, u2_key_r_40, u2_key_r_41, u2_key_r_42, 
       u2_key_r_43, u2_key_r_44, u2_key_r_46, u2_key_r_47, u2_key_r_48, u2_key_r_51, u2_key_r_53, u2_key_r_55, u2_key_r_6, 
       u2_key_r_7, u2_out0_1, u2_out0_10, u2_out0_11, u2_out0_12, u2_out0_13, u2_out0_14, u2_out0_15, u2_out0_16, 
       u2_out0_17, u2_out0_18, u2_out0_19, u2_out0_2, u2_out0_20, u2_out0_21, u2_out0_22, u2_out0_23, u2_out0_24, 
       u2_out0_25, u2_out0_26, u2_out0_27, u2_out0_28, u2_out0_29, u2_out0_3, u2_out0_30, u2_out0_31, u2_out0_32, 
       u2_out0_4, u2_out0_5, u2_out0_6, u2_out0_7, u2_out0_8, u2_out0_9, u2_out10_1, u2_out10_10, u2_out10_11, 
       u2_out10_13, u2_out10_16, u2_out10_17, u2_out10_18, u2_out10_19, u2_out10_2, u2_out10_20, u2_out10_23, u2_out10_24, 
       u2_out10_26, u2_out10_28, u2_out10_29, u2_out10_30, u2_out10_31, u2_out10_4, u2_out10_6, u2_out10_9, u2_out11_11, 
       u2_out11_12, u2_out11_13, u2_out11_14, u2_out11_18, u2_out11_19, u2_out11_2, u2_out11_22, u2_out11_25, u2_out11_28, 
       u2_out11_29, u2_out11_3, u2_out11_32, u2_out11_4, u2_out11_7, u2_out11_8, u2_out12_27, u2_out12_28, u2_out12_29, 
       u2_out13_1, u2_out13_10, u2_out13_11, u2_out13_12, u2_out13_14, u2_out13_19, u2_out13_20, u2_out13_22, u2_out13_25, 
       u2_out13_26, u2_out13_29, u2_out13_3, u2_out13_32, u2_out13_4, u2_out13_7, u2_out13_8, u2_out14_1, u2_out14_10, 
       u2_out14_11, u2_out14_12, u2_out14_14, u2_out14_15, u2_out14_17, u2_out14_19, u2_out14_20, u2_out14_21, u2_out14_22, 
       u2_out14_23, u2_out14_25, u2_out14_26, u2_out14_27, u2_out14_29, u2_out14_3, u2_out14_31, u2_out14_32, u2_out14_4, 
       u2_out14_5, u2_out14_7, u2_out14_8, u2_out14_9, u2_out15_1, u2_out15_10, u2_out15_13, u2_out15_14, u2_out15_16, 
       u2_out15_17, u2_out15_18, u2_out15_2, u2_out15_20, u2_out15_23, u2_out15_24, u2_out15_25, u2_out15_26, u2_out15_28, 
       u2_out15_3, u2_out15_30, u2_out15_31, u2_out15_6, u2_out15_8, u2_out15_9, u2_out1_1, u2_out1_10, u2_out1_11, 
       u2_out1_12, u2_out1_13, u2_out1_14, u2_out1_15, u2_out1_16, u2_out1_17, u2_out1_18, u2_out1_19, u2_out1_2, 
       u2_out1_20, u2_out1_21, u2_out1_22, u2_out1_23, u2_out1_24, u2_out1_25, u2_out1_26, u2_out1_27, u2_out1_28, 
       u2_out1_29, u2_out1_3, u2_out1_30, u2_out1_31, u2_out1_32, u2_out1_4, u2_out1_5, u2_out1_6, u2_out1_7, 
       u2_out1_8, u2_out1_9, u2_out2_1, u2_out2_10, u2_out2_11, u2_out2_12, u2_out2_13, u2_out2_14, u2_out2_15, 
       u2_out2_16, u2_out2_17, u2_out2_18, u2_out2_19, u2_out2_2, u2_out2_20, u2_out2_21, u2_out2_22, u2_out2_23, 
       u2_out2_24, u2_out2_25, u2_out2_26, u2_out2_27, u2_out2_28, u2_out2_29, u2_out2_3, u2_out2_30, u2_out2_31, 
       u2_out2_32, u2_out2_4, u2_out2_5, u2_out2_6, u2_out2_7, u2_out2_8, u2_out2_9, u2_out3_1, u2_out3_10, 
       u2_out3_11, u2_out3_12, u2_out3_13, u2_out3_14, u2_out3_15, u2_out3_16, u2_out3_17, u2_out3_18, u2_out3_19, 
       u2_out3_2, u2_out3_20, u2_out3_21, u2_out3_22, u2_out3_23, u2_out3_24, u2_out3_25, u2_out3_26, u2_out3_27, 
       u2_out3_28, u2_out3_29, u2_out3_3, u2_out3_30, u2_out3_31, u2_out3_32, u2_out3_4, u2_out3_5, u2_out3_6, 
       u2_out3_7, u2_out3_8, u2_out3_9, u2_out4_1, u2_out4_10, u2_out4_11, u2_out4_12, u2_out4_13, u2_out4_14, 
       u2_out4_15, u2_out4_16, u2_out4_17, u2_out4_18, u2_out4_19, u2_out4_2, u2_out4_20, u2_out4_21, u2_out4_22, 
       u2_out4_23, u2_out4_24, u2_out4_25, u2_out4_26, u2_out4_27, u2_out4_28, u2_out4_29, u2_out4_3, u2_out4_30, 
       u2_out4_31, u2_out4_32, u2_out4_4, u2_out4_5, u2_out4_6, u2_out4_7, u2_out4_8, u2_out4_9, u2_out5_1, 
       u2_out5_10, u2_out5_11, u2_out5_12, u2_out5_13, u2_out5_14, u2_out5_15, u2_out5_16, u2_out5_17, u2_out5_18, 
       u2_out5_19, u2_out5_2, u2_out5_20, u2_out5_21, u2_out5_22, u2_out5_23, u2_out5_24, u2_out5_25, u2_out5_26, 
       u2_out5_27, u2_out5_28, u2_out5_29, u2_out5_3, u2_out5_30, u2_out5_31, u2_out5_32, u2_out5_4, u2_out5_5, 
       u2_out5_6, u2_out5_7, u2_out5_8, u2_out5_9, u2_out6_1, u2_out6_10, u2_out6_11, u2_out6_12, u2_out6_13, 
       u2_out6_14, u2_out6_15, u2_out6_16, u2_out6_17, u2_out6_18, u2_out6_19, u2_out6_2, u2_out6_20, u2_out6_21, 
       u2_out6_22, u2_out6_23, u2_out6_24, u2_out6_25, u2_out6_26, u2_out6_27, u2_out6_28, u2_out6_29, u2_out6_3, 
       u2_out6_30, u2_out6_31, u2_out6_32, u2_out6_4, u2_out6_5, u2_out6_6, u2_out6_7, u2_out6_8, u2_out6_9, 
       u2_out7_1, u2_out7_10, u2_out7_12, u2_out7_13, u2_out7_16, u2_out7_17, u2_out7_18, u2_out7_2, u2_out7_20, 
       u2_out7_23, u2_out7_24, u2_out7_26, u2_out7_28, u2_out7_30, u2_out7_31, u2_out7_6, u2_out7_9, u2_out8_1, 
       u2_out8_10, u2_out8_13, u2_out8_14, u2_out8_16, u2_out8_18, u2_out8_2, u2_out8_20, u2_out8_24, u2_out8_25, 
       u2_out8_26, u2_out8_28, u2_out8_3, u2_out8_30, u2_out8_6, u2_out8_8, u2_out9_1, u2_out9_10, u2_out9_11, 
       u2_out9_12, u2_out9_13, u2_out9_14, u2_out9_15, u2_out9_16, u2_out9_17, u2_out9_18, u2_out9_19, u2_out9_2, 
       u2_out9_20, u2_out9_21, u2_out9_22, u2_out9_23, u2_out9_24, u2_out9_25, u2_out9_26, u2_out9_27, u2_out9_28, 
       u2_out9_29, u2_out9_3, u2_out9_30, u2_out9_31, u2_out9_32, u2_out9_4, u2_out9_5, u2_out9_6, u2_out9_7, 
       u2_out9_8, u2_out9_9, u2_u0_X_15, u2_u0_X_16, u2_u0_X_28, u2_u0_X_34, u2_u0_X_40, u2_u0_X_45, u2_u0_X_46, 
       u2_u0_X_5, u2_u0_X_7, u2_u0_X_9, u2_u10_X_10, u2_u10_X_15, u2_u10_X_16, u2_u10_X_21, u2_u10_X_33, u2_u10_X_34, 
       u2_u10_X_4, u2_u10_X_9, u2_u11_X_27, u2_u11_X_29, u2_u11_X_31, u2_u11_X_33, u2_u11_X_34, u2_u11_X_35, u2_u11_X_36, 
       u2_u11_X_37, u2_u11_X_38, u2_u11_X_39, u2_u11_X_40, u2_u11_X_9, u2_u13_X_19, u2_u13_X_20, u2_u13_X_21, u2_u13_X_22, 
       u2_u13_X_23, u2_u13_X_25, u2_u13_X_28, u2_u13_X_39, u2_u14_X_21, u2_u14_X_22, u2_u14_X_23, u2_u14_X_25, u2_u14_X_28, 
       u2_u14_X_3, u2_u14_X_30, u2_u14_X_32, u2_u14_X_34, u2_u14_X_39, u2_u14_X_4, u2_u14_X_46, u2_u15_X_10, u2_u15_X_16, 
       u2_u15_X_18, u2_u15_X_20, u2_u15_X_27, u2_u15_X_9, u2_u1_X_16, u2_u1_X_23, u2_u1_X_25, u2_u1_X_3, u2_u1_X_33, 
       u2_u1_X_34, u2_u1_X_35, u2_u1_X_37, u2_u1_X_39, u2_u1_X_40, u2_u1_X_42, u2_u1_X_44, u2_u1_X_45, u2_u1_X_46, 
       u2_u2_X_1, u2_u2_X_10, u2_u2_X_15, u2_u2_X_16, u2_u2_X_18, u2_u2_X_20, u2_u2_X_21, u2_u2_X_22, u2_u2_X_27, 
       u2_u2_X_3, u2_u2_X_30, u2_u2_X_32, u2_u2_X_34, u2_u2_X_39, u2_u2_X_41, u2_u2_X_42, u2_u2_X_43, u2_u2_X_44, 
       u2_u2_X_46, u2_u2_X_47, u2_u2_X_5, u2_u2_X_7, u2_u2_X_9, u2_u3_X_15, u2_u3_X_21, u2_u3_X_22, u2_u3_X_27, 
       u2_u3_X_28, u2_u3_X_33, u2_u3_X_34, u2_u3_X_36, u2_u3_X_38, u2_u3_X_39, u2_u3_X_40, u2_u3_X_42, u2_u3_X_44, 
       u2_u3_X_45, u2_u3_X_46, u2_u3_X_5, u2_u3_X_6, u2_u3_X_7, u2_u3_X_8, u2_u4_X_1, u2_u4_X_10, u2_u4_X_15, 
       u2_u4_X_16, u2_u4_X_21, u2_u4_X_23, u2_u4_X_24, u2_u4_X_25, u2_u4_X_26, u2_u4_X_28, u2_u4_X_3, u2_u4_X_33, 
       u2_u4_X_34, u2_u4_X_36, u2_u4_X_38, u2_u4_X_39, u2_u4_X_40, u2_u4_X_46, u2_u4_X_47, u2_u4_X_9, u2_u5_X_1, 
       u2_u5_X_12, u2_u5_X_14, u2_u5_X_15, u2_u5_X_16, u2_u5_X_22, u2_u5_X_27, u2_u5_X_3, u2_u5_X_30, u2_u5_X_32, 
       u2_u5_X_33, u2_u5_X_34, u2_u5_X_4, u2_u5_X_40, u2_u5_X_45, u2_u5_X_46, u2_u5_X_47, u2_u6_X_10, u2_u6_X_22, 
       u2_u6_X_28, u2_u6_X_29, u2_u6_X_3, u2_u6_X_31, u2_u6_X_33, u2_u6_X_4, u2_u6_X_40, u2_u6_X_45, u2_u6_X_46, 
       u2_u6_X_9, u2_u7_X_21, u2_u7_X_4, u2_u8_X_15, u2_u8_X_27, u2_u8_X_28, u2_u9_X_10, u2_u9_X_15, u2_u9_X_16, 
       u2_u9_X_21, u2_u9_X_3, u2_u9_X_30, u2_u9_X_32, u2_u9_X_34, u2_u9_X_4, u2_u9_X_45, u2_u9_X_46, u2_uk_K_r0_11, 
       u2_uk_K_r0_15, u2_uk_K_r0_17, u2_uk_K_r0_25, u2_uk_K_r0_32, u2_uk_K_r0_36, u2_uk_K_r0_47, u2_uk_K_r0_49, u2_uk_K_r10_10, u2_uk_K_r10_25, 
       u2_uk_K_r10_27, u2_uk_K_r10_32, u2_uk_K_r10_34, u2_uk_K_r10_4, u2_uk_K_r10_41, u2_uk_K_r10_43, u2_uk_K_r11_10, u2_uk_K_r11_11, u2_uk_K_r11_19, 
       u2_uk_K_r11_20, u2_uk_K_r11_21, u2_uk_K_r11_24, u2_uk_K_r11_25, u2_uk_K_r11_26, u2_uk_K_r11_27, u2_uk_K_r11_28, u2_uk_K_r11_29, u2_uk_K_r11_39, 
       u2_uk_K_r11_47, u2_uk_K_r11_48, u2_uk_K_r11_53, u2_uk_K_r11_6, u2_uk_K_r12_10, u2_uk_K_r12_15, u2_uk_K_r12_16, u2_uk_K_r12_25, u2_uk_K_r12_33, 
       u2_uk_K_r12_41, u2_uk_K_r12_42, u2_uk_K_r13_19, u2_uk_K_r13_25, u2_uk_K_r13_32, u2_uk_K_r13_55, u2_uk_K_r14_10, u2_uk_K_r14_12, u2_uk_K_r14_15, 
       u2_uk_K_r14_16, u2_uk_K_r14_18, u2_uk_K_r14_2, u2_uk_K_r14_3, u2_uk_K_r14_45, u2_uk_K_r14_46, u2_uk_K_r14_50, u2_uk_K_r14_9, u2_uk_K_r1_16, 
       u2_uk_K_r1_21, u2_uk_K_r1_44, u2_uk_K_r2_13, u2_uk_K_r2_18, u2_uk_K_r2_25, u2_uk_K_r2_27, u2_uk_K_r2_28, u2_uk_K_r2_31, u2_uk_K_r2_36, 
       u2_uk_K_r2_49, u2_uk_K_r2_55, u2_uk_K_r3_11, u2_uk_K_r3_19, u2_uk_K_r3_4, u2_uk_K_r3_43, u2_uk_K_r3_9, u2_uk_K_r4_0, u2_uk_K_r4_11, 
       u2_uk_K_r4_17, u2_uk_K_r4_33, u2_uk_K_r4_35, u2_uk_K_r4_38, u2_uk_K_r4_4, u2_uk_K_r4_5, u2_uk_K_r4_55, u2_uk_K_r5_10, u2_uk_K_r5_19, 
       u2_uk_K_r5_41, u2_uk_K_r6_0, u2_uk_K_r6_10, u2_uk_K_r6_14, u2_uk_K_r6_26, u2_uk_K_r6_29, u2_uk_K_r6_3, u2_uk_K_r6_31, u2_uk_K_r6_34, 
       u2_uk_K_r6_37, u2_uk_K_r6_51, u2_uk_K_r6_53, u2_uk_K_r6_7, u2_uk_K_r7_0, u2_uk_K_r7_25, u2_uk_K_r7_26, u2_uk_K_r7_31, u2_uk_K_r7_32, 
       u2_uk_K_r7_37, u2_uk_K_r7_39, u2_uk_K_r7_46, u2_uk_K_r8_13, u2_uk_K_r8_16, u2_uk_K_r8_2, u2_uk_K_r8_22, u2_uk_K_r8_37, u2_uk_K_r8_40, 
       u2_uk_K_r8_41, u2_uk_K_r8_42, u2_uk_K_r8_43, u2_uk_K_r8_48, u2_uk_K_r9_10, u2_uk_K_r9_13, u2_uk_K_r9_15, u2_uk_K_r9_19, u2_uk_K_r9_23, 
       u2_uk_K_r9_25, u2_uk_K_r9_27, u2_uk_K_r9_31, u2_uk_K_r9_4, u2_uk_K_r9_48, u2_uk_K_r9_55, u2_uk_n10, u2_uk_n100, u2_uk_n1001, 
       u2_uk_n1004, u2_uk_n1008, u2_uk_n102, u2_uk_n1020, u2_uk_n1024, u2_uk_n1027, u2_uk_n1028, u2_uk_n1031, u2_uk_n1035, 
       u2_uk_n1036, u2_uk_n1043, u2_uk_n1044, u2_uk_n1046, u2_uk_n1049, u2_uk_n1053, u2_uk_n1058, u2_uk_n1069, u2_uk_n1074, 
       u2_uk_n1075, u2_uk_n1076, u2_uk_n1077, u2_uk_n1079, u2_uk_n1082, u2_uk_n1083, u2_uk_n1084, u2_uk_n1085, u2_uk_n1088, 
       u2_uk_n1089, u2_uk_n109, u2_uk_n1091, u2_uk_n1093, u2_uk_n1095, u2_uk_n1096, u2_uk_n1097, u2_uk_n11, u2_uk_n110, 
       u2_uk_n1100, u2_uk_n1104, u2_uk_n1105, u2_uk_n1107, u2_uk_n1113, u2_uk_n1118, u2_uk_n1120, u2_uk_n1124, u2_uk_n1125, 
       u2_uk_n1127, u2_uk_n1128, u2_uk_n1130, u2_uk_n1131, u2_uk_n1132, u2_uk_n1133, u2_uk_n1134, u2_uk_n1136, u2_uk_n1137, 
       u2_uk_n1140, u2_uk_n1141, u2_uk_n1142, u2_uk_n1145, u2_uk_n1146, u2_uk_n1152, u2_uk_n1161, u2_uk_n1167, u2_uk_n1168, 
       u2_uk_n117, u2_uk_n1171, u2_uk_n1178, u2_uk_n1179, u2_uk_n118, u2_uk_n1188, u2_uk_n1189, u2_uk_n1190, u2_uk_n1194, 
       u2_uk_n1197, u2_uk_n1198, u2_uk_n1199, u2_uk_n1200, u2_uk_n1201, u2_uk_n1203, u2_uk_n1204, u2_uk_n1205, u2_uk_n1206, 
       u2_uk_n1207, u2_uk_n1208, u2_uk_n1209, u2_uk_n1210, u2_uk_n1212, u2_uk_n1213, u2_uk_n1215, u2_uk_n1216, u2_uk_n1217, 
       u2_uk_n1218, u2_uk_n1220, u2_uk_n1221, u2_uk_n1223, u2_uk_n1225, u2_uk_n1226, u2_uk_n1227, u2_uk_n1228, u2_uk_n1230, 
       u2_uk_n1231, u2_uk_n1232, u2_uk_n1234, u2_uk_n1238, u2_uk_n1240, u2_uk_n1243, u2_uk_n1244, u2_uk_n1245, u2_uk_n1246, 
       u2_uk_n1247, u2_uk_n1249, u2_uk_n1259, u2_uk_n1260, u2_uk_n1261, u2_uk_n1265, u2_uk_n1267, u2_uk_n1270, u2_uk_n1275, 
       u2_uk_n1279, u2_uk_n128, u2_uk_n1280, u2_uk_n1282, u2_uk_n1283, u2_uk_n1284, u2_uk_n1285, u2_uk_n1287, u2_uk_n129, 
       u2_uk_n1292, u2_uk_n1293, u2_uk_n1296, u2_uk_n1298, u2_uk_n1300, u2_uk_n1301, u2_uk_n1303, u2_uk_n1305, u2_uk_n1306, 
       u2_uk_n1309, u2_uk_n1310, u2_uk_n1311, u2_uk_n1313, u2_uk_n1314, u2_uk_n1317, u2_uk_n1319, u2_uk_n1322, u2_uk_n1323, 
       u2_uk_n1325, u2_uk_n1326, u2_uk_n1329, u2_uk_n1331, u2_uk_n1333, u2_uk_n1336, u2_uk_n1339, u2_uk_n1341, u2_uk_n1345, 
       u2_uk_n1350, u2_uk_n1353, u2_uk_n1359, u2_uk_n1361, u2_uk_n1363, u2_uk_n1365, u2_uk_n1370, u2_uk_n1375, u2_uk_n1381, 
       u2_uk_n1382, u2_uk_n1403, u2_uk_n1405, u2_uk_n1408, u2_uk_n141, u2_uk_n1411, u2_uk_n1412, u2_uk_n1418, u2_uk_n142, 
       u2_uk_n1420, u2_uk_n1425, u2_uk_n1428, u2_uk_n1430, u2_uk_n1435, u2_uk_n1438, u2_uk_n1439, u2_uk_n1445, u2_uk_n1446, 
       u2_uk_n1447, u2_uk_n145, u2_uk_n1453, u2_uk_n1454, u2_uk_n1456, u2_uk_n1458, u2_uk_n146, u2_uk_n1460, u2_uk_n1462, 
       u2_uk_n1465, u2_uk_n1466, u2_uk_n147, u2_uk_n1470, u2_uk_n1475, u2_uk_n148, u2_uk_n1486, u2_uk_n1488, u2_uk_n1491, 
       u2_uk_n1493, u2_uk_n1494, u2_uk_n1496, u2_uk_n1497, u2_uk_n1498, u2_uk_n1499, u2_uk_n1500, u2_uk_n1502, u2_uk_n1503, 
       u2_uk_n1504, u2_uk_n1506, u2_uk_n1508, u2_uk_n1511, u2_uk_n1513, u2_uk_n1514, u2_uk_n1515, u2_uk_n1517, u2_uk_n1518, 
       u2_uk_n1519, u2_uk_n1521, u2_uk_n1522, u2_uk_n1524, u2_uk_n1525, u2_uk_n1526, u2_uk_n1527, u2_uk_n1529, u2_uk_n1530, 
       u2_uk_n1531, u2_uk_n1532, u2_uk_n1533, u2_uk_n1535, u2_uk_n1536, u2_uk_n1537, u2_uk_n1538, u2_uk_n1542, u2_uk_n1544, 
       u2_uk_n1548, u2_uk_n1549, u2_uk_n155, u2_uk_n1551, u2_uk_n1555, u2_uk_n1556, u2_uk_n1558, u2_uk_n1563, u2_uk_n1565, 
       u2_uk_n1568, u2_uk_n1570, u2_uk_n1571, u2_uk_n1573, u2_uk_n1576, u2_uk_n1577, u2_uk_n1580, u2_uk_n1583, u2_uk_n1585, 
       u2_uk_n1586, u2_uk_n1590, u2_uk_n1591, u2_uk_n1592, u2_uk_n1594, u2_uk_n1599, u2_uk_n1600, u2_uk_n1602, u2_uk_n1604, 
       u2_uk_n1605, u2_uk_n1609, u2_uk_n161, u2_uk_n1610, u2_uk_n1615, u2_uk_n1617, u2_uk_n162, u2_uk_n1622, u2_uk_n1624, 
       u2_uk_n1626, u2_uk_n1629, u2_uk_n163, u2_uk_n1631, u2_uk_n1632, u2_uk_n1634, u2_uk_n1639, u2_uk_n164, u2_uk_n1640, 
       u2_uk_n1642, u2_uk_n1643, u2_uk_n1647, u2_uk_n1652, u2_uk_n1653, u2_uk_n1654, u2_uk_n1657, u2_uk_n1658, u2_uk_n1660, 
       u2_uk_n1665, u2_uk_n1666, u2_uk_n1668, u2_uk_n1672, u2_uk_n1673, u2_uk_n1674, u2_uk_n1675, u2_uk_n1677, u2_uk_n1680, 
       u2_uk_n1681, u2_uk_n1682, u2_uk_n1683, u2_uk_n1684, u2_uk_n1687, u2_uk_n1688, u2_uk_n1689, u2_uk_n1693, u2_uk_n17, 
       u2_uk_n1702, u2_uk_n1707, u2_uk_n1708, u2_uk_n1709, u2_uk_n1720, u2_uk_n1721, u2_uk_n1723, u2_uk_n1724, u2_uk_n1725, 
       u2_uk_n1726, u2_uk_n1727, u2_uk_n1728, u2_uk_n1731, u2_uk_n1732, u2_uk_n1734, u2_uk_n1736, u2_uk_n1737, u2_uk_n1738, 
       u2_uk_n1742, u2_uk_n1743, u2_uk_n1744, u2_uk_n1745, u2_uk_n1746, u2_uk_n1747, u2_uk_n1750, u2_uk_n1753, u2_uk_n1755, 
       u2_uk_n1761, u2_uk_n1762, u2_uk_n1763, u2_uk_n1767, u2_uk_n1769, u2_uk_n1770, u2_uk_n1773, u2_uk_n1776, u2_uk_n1777, 
       u2_uk_n1778, u2_uk_n1781, u2_uk_n1782, u2_uk_n1783, u2_uk_n1785, u2_uk_n1786, u2_uk_n1788, u2_uk_n1789, u2_uk_n1790, 
       u2_uk_n1791, u2_uk_n1792, u2_uk_n1793, u2_uk_n1794, u2_uk_n1796, u2_uk_n1797, u2_uk_n1800, u2_uk_n1801, u2_uk_n1803, 
       u2_uk_n1805, u2_uk_n1807, u2_uk_n1808, u2_uk_n1809, u2_uk_n1811, u2_uk_n1814, u2_uk_n1815, u2_uk_n1816, u2_uk_n1817, 
       u2_uk_n182, u2_uk_n1821, u2_uk_n1823, u2_uk_n1826, u2_uk_n1832, u2_uk_n1833, u2_uk_n1834, u2_uk_n1835, u2_uk_n1837, 
       u2_uk_n1839, u2_uk_n1840, u2_uk_n1843, u2_uk_n1849, u2_uk_n1850, u2_uk_n1851, u2_uk_n1852, u2_uk_n1853, u2_uk_n1855, 
       u2_uk_n187, u2_uk_n188, u2_uk_n191, u2_uk_n202, u2_uk_n203, u2_uk_n207, u2_uk_n208, u2_uk_n209, u2_uk_n213, 
       u2_uk_n214, u2_uk_n217, u2_uk_n220, u2_uk_n222, u2_uk_n223, u2_uk_n230, u2_uk_n231, u2_uk_n238, u2_uk_n240, 
       u2_uk_n251, u2_uk_n257, u2_uk_n27, u2_uk_n299, u2_uk_n301, u2_uk_n305, u2_uk_n308, u2_uk_n31, u2_uk_n313, 
       u2_uk_n319, u2_uk_n363, u2_uk_n369, u2_uk_n373, u2_uk_n376, u2_uk_n379, u2_uk_n385, u2_uk_n407, u2_uk_n408, 
       u2_uk_n415, u2_uk_n421, u2_uk_n443, u2_uk_n456, u2_uk_n467, u2_uk_n500, u2_uk_n503, u2_uk_n504, u2_uk_n520, 
       u2_uk_n526, u2_uk_n551, u2_uk_n586, u2_uk_n60, u2_uk_n608, u2_uk_n63, u2_uk_n665, u2_uk_n677, u2_uk_n682, 
       u2_uk_n689, u2_uk_n692, u2_uk_n694, u2_uk_n702, u2_uk_n83, u2_uk_n92, u2_uk_n93, u2_uk_n931, u2_uk_n933, 
       u2_uk_n939, u2_uk_n94, u2_uk_n942, u2_uk_n943, u2_uk_n944, u2_uk_n946, u2_uk_n947, u2_uk_n948, u2_uk_n954, 
       u2_uk_n955, u2_uk_n956, u2_uk_n961, u2_uk_n967, u2_uk_n970, u2_uk_n972, u2_uk_n984, u2_uk_n986, u2_uk_n99, 
       u2_uk_n991, u2_uk_n994, u2_uk_n997 ;

  des_des_die_0 u0 ( clk, decrypt, desIn, key1, key2, key3, desOut, u0_FP_11, u0_FP_12, u0_FP_14, u0_FP_15, u0_FP_19, u0_FP_21, u0_FP_22, u0_FP_25, 
      u0_FP_27, u0_FP_29, u0_FP_3, u0_FP_32, u0_FP_4, u0_FP_5, u0_FP_7, u0_FP_8, u0_N128, 
      u0_N129, u0_N130, u0_N132, u0_N133, u0_N135, u0_N136, u0_N137, u0_N140, u0_N141, 
      u0_N142, u0_N143, u0_N144, u0_N145, u0_N147, u0_N148, u0_N150, u0_N151, u0_N152, 
      u0_N153, u0_N154, u0_N155, u0_N157, u0_N158, u0_N256, u0_N257, u0_N258, u0_N259, 
      u0_N260, u0_N261, u0_N262, u0_N263, u0_N264, u0_N265, u0_N266, u0_N267, u0_N268, 
      u0_N269, u0_N270, u0_N271, u0_N272, u0_N273, u0_N274, u0_N275, u0_N276, u0_N277, 
      u0_N278, u0_N279, u0_N280, u0_N281, u0_N282, u0_N283, u0_N284, u0_N285, u0_N286, 
      u0_N287, u0_N288, u0_N289, u0_N293, u0_N296, u0_N297, u0_N300, u0_N303, u0_N304, 
      u0_N305, u0_N307, u0_N310, u0_N311, u0_N313, u0_N315, u0_N317, u0_N318, u0_N352, 
      u0_N353, u0_N354, u0_N355, u0_N356, u0_N357, u0_N358, u0_N359, u0_N360, u0_N361, 
      u0_N362, u0_N363, u0_N364, u0_N365, u0_N366, u0_N367, u0_N368, u0_N369, u0_N370, 
      u0_N371, u0_N372, u0_N373, u0_N374, u0_N375, u0_N376, u0_N377, u0_N378, u0_N379, 
      u0_N380, u0_N381, u0_N382, u0_N383, u0_N417, u0_N421, u0_N424, u0_N428, u0_N431, 
      u0_N432, u0_N433, u0_N438, u0_N439, u0_N443, u0_N445, u0_N446, u0_N448, u0_N449, 
      u0_N457, u0_N460, u0_N465, u0_N467, u0_N473, u0_N475, u0_out0_1, u0_out0_10, u0_out0_11, 
      u0_out0_12, u0_out0_13, u0_out0_14, u0_out0_15, u0_out0_16, u0_out0_17, u0_out0_18, u0_out0_19, u0_out0_2, 
      u0_out0_20, u0_out0_21, u0_out0_22, u0_out0_23, u0_out0_24, u0_out0_25, u0_out0_26, u0_out0_27, u0_out0_28, 
      u0_out0_29, u0_out0_3, u0_out0_30, u0_out0_31, u0_out0_32, u0_out0_4, u0_out0_5, u0_out0_6, u0_out0_7, 
      u0_out0_8, u0_out0_9, u0_out10_1, u0_out10_10, u0_out10_11, u0_out10_12, u0_out10_13, u0_out10_14, u0_out10_15, 
      u0_out10_16, u0_out10_17, u0_out10_18, u0_out10_19, u0_out10_2, u0_out10_20, u0_out10_21, u0_out10_22, u0_out10_23, 
      u0_out10_24, u0_out10_25, u0_out10_26, u0_out10_27, u0_out10_28, u0_out10_29, u0_out10_3, u0_out10_30, u0_out10_31, 
      u0_out10_32, u0_out10_4, u0_out10_5, u0_out10_6, u0_out10_7, u0_out10_8, u0_out10_9, u0_out12_1, u0_out12_10, 
      u0_out12_11, u0_out12_12, u0_out12_13, u0_out12_14, u0_out12_15, u0_out12_16, u0_out12_17, u0_out12_18, u0_out12_19, 
      u0_out12_2, u0_out12_20, u0_out12_21, u0_out12_22, u0_out12_23, u0_out12_24, u0_out12_25, u0_out12_26, u0_out12_27, 
      u0_out12_28, u0_out12_29, u0_out12_3, u0_out12_30, u0_out12_31, u0_out12_32, u0_out12_4, u0_out12_5, u0_out12_6, 
      u0_out12_7, u0_out12_8, u0_out12_9, u0_out13_1, u0_out13_10, u0_out13_11, u0_out13_12, u0_out13_14, u0_out13_15, 
      u0_out13_19, u0_out13_20, u0_out13_21, u0_out13_22, u0_out13_25, u0_out13_26, u0_out13_27, u0_out13_29, u0_out13_3, 
      u0_out13_32, u0_out13_4, u0_out13_5, u0_out13_7, u0_out13_8, u0_out14_11, u0_out14_12, u0_out14_14, u0_out14_15, 
      u0_out14_16, u0_out14_17, u0_out14_19, u0_out14_21, u0_out14_22, u0_out14_23, u0_out14_24, u0_out14_25, u0_out14_27, 
      u0_out14_29, u0_out14_3, u0_out14_30, u0_out14_31, u0_out14_32, u0_out14_4, u0_out14_5, u0_out14_6, u0_out14_7, 
      u0_out14_8, u0_out14_9, u0_out15_1, u0_out15_10, u0_out15_13, u0_out15_16, u0_out15_17, u0_out15_18, u0_out15_2, 
      u0_out15_20, u0_out15_23, u0_out15_24, u0_out15_26, u0_out15_28, u0_out15_30, u0_out15_31, u0_out15_6, u0_out15_9, 
      u0_out1_1, u0_out1_10, u0_out1_11, u0_out1_12, u0_out1_13, u0_out1_14, u0_out1_15, u0_out1_16, u0_out1_17, 
      u0_out1_18, u0_out1_19, u0_out1_2, u0_out1_20, u0_out1_21, u0_out1_22, u0_out1_23, u0_out1_24, u0_out1_25, 
      u0_out1_26, u0_out1_27, u0_out1_28, u0_out1_29, u0_out1_3, u0_out1_30, u0_out1_31, u0_out1_32, u0_out1_4, 
      u0_out1_5, u0_out1_6, u0_out1_7, u0_out1_8, u0_out1_9, u0_out2_1, u0_out2_10, u0_out2_11, u0_out2_12, 
      u0_out2_13, u0_out2_14, u0_out2_15, u0_out2_16, u0_out2_17, u0_out2_18, u0_out2_19, u0_out2_2, u0_out2_20, 
      u0_out2_21, u0_out2_22, u0_out2_23, u0_out2_24, u0_out2_25, u0_out2_26, u0_out2_27, u0_out2_28, u0_out2_29, 
      u0_out2_3, u0_out2_30, u0_out2_31, u0_out2_32, u0_out2_4, u0_out2_5, u0_out2_6, u0_out2_7, u0_out2_8, 
      u0_out2_9, u0_out3_1, u0_out3_10, u0_out3_11, u0_out3_12, u0_out3_13, u0_out3_14, u0_out3_15, u0_out3_16, 
      u0_out3_17, u0_out3_18, u0_out3_19, u0_out3_2, u0_out3_20, u0_out3_21, u0_out3_22, u0_out3_23, u0_out3_24, 
      u0_out3_25, u0_out3_26, u0_out3_27, u0_out3_28, u0_out3_29, u0_out3_3, u0_out3_30, u0_out3_31, u0_out3_32, 
      u0_out3_4, u0_out3_5, u0_out3_6, u0_out3_7, u0_out3_8, u0_out3_9, u0_out4_11, u0_out4_12, u0_out4_19, 
      u0_out4_22, u0_out4_29, u0_out4_32, u0_out4_4, u0_out4_7, u0_out5_1, u0_out5_10, u0_out5_11, u0_out5_12, 
      u0_out5_13, u0_out5_14, u0_out5_15, u0_out5_16, u0_out5_17, u0_out5_18, u0_out5_19, u0_out5_2, u0_out5_20, 
      u0_out5_21, u0_out5_22, u0_out5_23, u0_out5_24, u0_out5_25, u0_out5_26, u0_out5_27, u0_out5_28, u0_out5_29, 
      u0_out5_3, u0_out5_30, u0_out5_31, u0_out5_32, u0_out5_4, u0_out5_5, u0_out5_6, u0_out5_7, u0_out5_8, 
      u0_out5_9, u0_out6_1, u0_out6_10, u0_out6_11, u0_out6_12, u0_out6_13, u0_out6_14, u0_out6_15, u0_out6_16, 
      u0_out6_17, u0_out6_18, u0_out6_19, u0_out6_2, u0_out6_20, u0_out6_21, u0_out6_22, u0_out6_23, u0_out6_24, 
      u0_out6_25, u0_out6_26, u0_out6_27, u0_out6_28, u0_out6_29, u0_out6_3, u0_out6_30, u0_out6_31, u0_out6_32, 
      u0_out6_4, u0_out6_5, u0_out6_6, u0_out6_7, u0_out6_8, u0_out6_9, u0_out7_1, u0_out7_10, u0_out7_11, 
      u0_out7_12, u0_out7_13, u0_out7_14, u0_out7_15, u0_out7_16, u0_out7_17, u0_out7_18, u0_out7_19, u0_out7_2, 
      u0_out7_20, u0_out7_21, u0_out7_22, u0_out7_23, u0_out7_24, u0_out7_25, u0_out7_26, u0_out7_27, u0_out7_28, 
      u0_out7_29, u0_out7_3, u0_out7_30, u0_out7_31, u0_out7_32, u0_out7_4, u0_out7_5, u0_out7_6, u0_out7_7, 
      u0_out7_8, u0_out7_9, u0_out9_11, u0_out9_12, u0_out9_14, u0_out9_15, u0_out9_19, u0_out9_21, u0_out9_22, 
      u0_out9_25, u0_out9_27, u0_out9_29, u0_out9_3, u0_out9_32, u0_out9_4, u0_out9_5, u0_out9_7, u0_out9_8, 
      u0_uk_n10, u0_uk_n100, u0_uk_n102, u0_uk_n109, u0_uk_n11, u0_uk_n110, u0_uk_n117, u0_uk_n118, u0_uk_n128, 
      u0_uk_n129, u0_uk_n141, u0_uk_n142, u0_uk_n145, u0_uk_n146, u0_uk_n147, u0_uk_n148, u0_uk_n155, u0_uk_n161, 
      u0_uk_n162, u0_uk_n163, u0_uk_n164, u0_uk_n17, u0_uk_n182, u0_uk_n187, u0_uk_n188, u0_uk_n191, u0_uk_n202, 
      u0_uk_n203, u0_uk_n207, u0_uk_n208, u0_uk_n209, u0_uk_n213, u0_uk_n214, u0_uk_n217, u0_uk_n220, u0_uk_n222, 
      u0_uk_n223, u0_uk_n230, u0_uk_n231, u0_uk_n238, u0_uk_n240, u0_uk_n242, u0_uk_n250, u0_uk_n251, u0_uk_n252, 
      u0_uk_n27, u0_uk_n31, u0_uk_n60, u0_uk_n63, u0_uk_n684, u0_uk_n687, u0_uk_n690, u0_uk_n696, u0_uk_n697, 
      u0_uk_n698, u0_uk_n705, u0_uk_n707, u0_uk_n83, u0_uk_n92, u0_uk_n93, u0_uk_n94, u0_uk_n99, u1_out0_1, 
      u1_out0_10, u1_out0_11, u1_out0_12, u1_out0_13, u1_out0_14, u1_out0_15, u1_out0_16, u1_out0_17, u1_out0_18, 
      u1_out0_19, u1_out0_2, u1_out0_20, u1_out0_21, u1_out0_22, u1_out0_23, u1_out0_24, u1_out0_25, u1_out0_26, 
      u1_out0_27, u1_out0_28, u1_out0_29, u1_out0_3, u1_out0_30, u1_out0_31, u1_out0_32, u1_out0_4, u1_out0_5, 
      u1_out0_6, u1_out0_7, u1_out0_8, u1_out0_9, u1_out10_1, u1_out10_10, u1_out10_11, u1_out10_12, u1_out10_13, 
      u1_out10_14, u1_out10_15, u1_out10_16, u1_out10_17, u1_out10_18, u1_out10_19, u1_out10_2, u1_out10_20, u1_out10_21, 
      u1_out10_22, u1_out10_23, u1_out10_24, u1_out10_25, u1_out10_26, u1_out10_27, u1_out10_28, u1_out10_29, u1_out10_3, 
      u1_out10_30, u1_out10_31, u1_out10_32, u1_out10_4, u1_out10_5, u1_out10_6, u1_out10_7, u1_out10_8, u1_out10_9, 
      u1_out11_1, u1_out11_10, u1_out11_11, u1_out11_12, u1_out11_13, u1_out11_14, u1_out11_15, u1_out11_16, u1_out11_17, 
      u1_out11_18, u1_out11_19, u1_out11_2, u1_out11_20, u1_out11_21, u1_out11_22, u1_out11_23, u1_out11_24, u1_out11_25, 
      u1_out11_26, u1_out11_27, u1_out11_28, u1_out11_29, u1_out11_3, u1_out11_30, u1_out11_31, u1_out11_32, u1_out11_4, 
      u1_out11_5, u1_out11_6, u1_out11_7, u1_out11_8, u1_out11_9, u1_out12_1, u1_out12_10, u1_out12_11, u1_out12_12, 
      u1_out12_13, u1_out12_14, u1_out12_15, u1_out12_16, u1_out12_17, u1_out12_18, u1_out12_19, u1_out12_2, u1_out12_20, 
      u1_out12_21, u1_out12_22, u1_out12_23, u1_out12_24, u1_out12_25, u1_out12_26, u1_out12_27, u1_out12_28, u1_out12_29, 
      u1_out12_3, u1_out12_30, u1_out12_31, u1_out12_32, u1_out12_4, u1_out12_5, u1_out12_6, u1_out12_7, u1_out12_8, 
      u1_out12_9, u1_out13_1, u1_out13_10, u1_out13_11, u1_out13_12, u1_out13_13, u1_out13_14, u1_out13_15, u1_out13_16, 
      u1_out13_17, u1_out13_18, u1_out13_19, u1_out13_2, u1_out13_20, u1_out13_21, u1_out13_22, u1_out13_23, u1_out13_24, 
      u1_out13_25, u1_out13_26, u1_out13_27, u1_out13_28, u1_out13_29, u1_out13_3, u1_out13_30, u1_out13_31, u1_out13_32, 
      u1_out13_4, u1_out13_5, u1_out13_6, u1_out13_7, u1_out13_8, u1_out13_9, u1_out14_1, u1_out14_10, u1_out14_11, 
      u1_out14_12, u1_out14_13, u1_out14_14, u1_out14_15, u1_out14_16, u1_out14_17, u1_out14_18, u1_out14_19, u1_out14_2, 
      u1_out14_20, u1_out14_21, u1_out14_22, u1_out14_23, u1_out14_24, u1_out14_25, u1_out14_26, u1_out14_27, u1_out14_28, 
      u1_out14_29, u1_out14_3, u1_out14_30, u1_out14_31, u1_out14_32, u1_out14_4, u1_out14_5, u1_out14_6, u1_out14_7, 
      u1_out14_8, u1_out14_9, u1_out15_1, u1_out15_10, u1_out15_11, u1_out15_12, u1_out15_13, u1_out15_14, u1_out15_15, 
      u1_out15_16, u1_out15_17, u1_out15_18, u1_out15_19, u1_out15_2, u1_out15_20, u1_out15_21, u1_out15_22, u1_out15_23, 
      u1_out15_24, u1_out15_25, u1_out15_26, u1_out15_27, u1_out15_28, u1_out15_29, u1_out15_3, u1_out15_30, u1_out15_31, 
      u1_out15_32, u1_out15_4, u1_out15_5, u1_out15_6, u1_out15_7, u1_out15_8, u1_out15_9, u1_out1_1, u1_out1_10, 
      u1_out1_11, u1_out1_12, u1_out1_13, u1_out1_14, u1_out1_15, u1_out1_16, u1_out1_17, u1_out1_18, u1_out1_19, 
      u1_out1_2, u1_out1_20, u1_out1_21, u1_out1_22, u1_out1_23, u1_out1_24, u1_out1_25, u1_out1_26, u1_out1_27, 
      u1_out1_28, u1_out1_29, u1_out1_3, u1_out1_30, u1_out1_31, u1_out1_32, u1_out1_4, u1_out1_5, u1_out1_6, 
      u1_out1_7, u1_out1_8, u1_out1_9, u1_out2_1, u1_out2_10, u1_out2_11, u1_out2_12, u1_out2_13, u1_out2_14, 
      u1_out2_15, u1_out2_16, u1_out2_17, u1_out2_18, u1_out2_19, u1_out2_2, u1_out2_20, u1_out2_21, u1_out2_22, 
      u1_out2_23, u1_out2_24, u1_out2_25, u1_out2_26, u1_out2_27, u1_out2_28, u1_out2_29, u1_out2_3, u1_out2_30, 
      u1_out2_31, u1_out2_32, u1_out2_4, u1_out2_5, u1_out2_6, u1_out2_7, u1_out2_8, u1_out2_9, u1_out3_1, 
      u1_out3_10, u1_out3_11, u1_out3_12, u1_out3_13, u1_out3_14, u1_out3_15, u1_out3_16, u1_out3_17, u1_out3_18, 
      u1_out3_19, u1_out3_2, u1_out3_20, u1_out3_21, u1_out3_22, u1_out3_23, u1_out3_24, u1_out3_25, u1_out3_26, 
      u1_out3_27, u1_out3_28, u1_out3_29, u1_out3_3, u1_out3_30, u1_out3_31, u1_out3_32, u1_out3_4, u1_out3_5, 
      u1_out3_6, u1_out3_7, u1_out3_8, u1_out3_9, u1_out4_1, u1_out4_10, u1_out4_11, u1_out4_12, u1_out4_13, 
      u1_out4_14, u1_out4_15, u1_out4_16, u1_out4_17, u1_out4_18, u1_out4_19, u1_out4_2, u1_out4_20, u1_out4_21, 
      u1_out4_22, u1_out4_23, u1_out4_24, u1_out4_25, u1_out4_26, u1_out4_27, u1_out4_28, u1_out4_29, u1_out4_3, 
      u1_out4_30, u1_out4_31, u1_out4_32, u1_out4_4, u1_out4_5, u1_out4_6, u1_out4_7, u1_out4_8, u1_out4_9, 
      u1_out5_1, u1_out5_10, u1_out5_11, u1_out5_12, u1_out5_13, u1_out5_14, u1_out5_15, u1_out5_16, u1_out5_17, 
      u1_out5_18, u1_out5_19, u1_out5_2, u1_out5_20, u1_out5_21, u1_out5_22, u1_out5_23, u1_out5_24, u1_out5_25, 
      u1_out5_26, u1_out5_27, u1_out5_28, u1_out5_29, u1_out5_3, u1_out5_30, u1_out5_31, u1_out5_32, u1_out5_4, 
      u1_out5_5, u1_out5_6, u1_out5_7, u1_out5_8, u1_out5_9, u1_out6_1, u1_out6_10, u1_out6_11, u1_out6_12, 
      u1_out6_13, u1_out6_14, u1_out6_15, u1_out6_16, u1_out6_17, u1_out6_18, u1_out6_19, u1_out6_2, u1_out6_20, 
      u1_out6_21, u1_out6_22, u1_out6_23, u1_out6_24, u1_out6_25, u1_out6_26, u1_out6_27, u1_out6_28, u1_out6_29, 
      u1_out6_3, u1_out6_30, u1_out6_31, u1_out6_32, u1_out6_4, u1_out6_5, u1_out6_6, u1_out6_7, u1_out6_8, 
      u1_out6_9, u1_out7_1, u1_out7_10, u1_out7_11, u1_out7_12, u1_out7_13, u1_out7_14, u1_out7_15, u1_out7_16, 
      u1_out7_17, u1_out7_18, u1_out7_19, u1_out7_2, u1_out7_20, u1_out7_21, u1_out7_22, u1_out7_23, u1_out7_24, 
      u1_out7_25, u1_out7_26, u1_out7_27, u1_out7_28, u1_out7_29, u1_out7_3, u1_out7_30, u1_out7_31, u1_out7_32, 
      u1_out7_4, u1_out7_5, u1_out7_6, u1_out7_7, u1_out7_8, u1_out7_9, u1_out8_1, u1_out8_10, u1_out8_11, 
      u1_out8_12, u1_out8_13, u1_out8_14, u1_out8_15, u1_out8_16, u1_out8_17, u1_out8_18, u1_out8_19, u1_out8_2, 
      u1_out8_20, u1_out8_21, u1_out8_22, u1_out8_23, u1_out8_24, u1_out8_25, u1_out8_26, u1_out8_27, u1_out8_28, 
      u1_out8_29, u1_out8_3, u1_out8_30, u1_out8_31, u1_out8_32, u1_out8_4, u1_out8_5, u1_out8_6, u1_out8_7, 
      u1_out8_8, u1_out8_9, u1_out9_1, u1_out9_10, u1_out9_11, u1_out9_12, u1_out9_13, u1_out9_14, u1_out9_15, 
      u1_out9_16, u1_out9_17, u1_out9_18, u1_out9_19, u1_out9_2, u1_out9_20, u1_out9_21, u1_out9_22, u1_out9_23, 
      u1_out9_24, u1_out9_25, u1_out9_26, u1_out9_27, u1_out9_28, u1_out9_29, u1_out9_3, u1_out9_30, u1_out9_31, 
      u1_out9_32, u1_out9_4, u1_out9_5, u1_out9_6, u1_out9_7, u1_out9_8, u1_out9_9, u2_FP_11, u2_FP_12, 
      u2_FP_15, u2_FP_19, u2_FP_21, u2_FP_22, u2_FP_27, u2_FP_29, u2_FP_32, u2_FP_4, u2_FP_5, 
      u2_FP_7, u2_N226, u2_N227, u2_N228, u2_N230, u2_N231, u2_N234, u2_N237, u2_N238, 
      u2_N242, u2_N244, u2_N245, u2_N248, u2_N250, u2_N252, u2_N255, u2_N259, u2_N260, 
      u2_N262, u2_N264, u2_N266, u2_N267, u2_N270, u2_N272, u2_N274, u2_N276, u2_N277, 
      u2_N278, u2_N282, u2_N284, u2_N286, u2_N287, u2_N322, u2_N324, u2_N326, u2_N327, 
      u2_N331, u2_N333, u2_N334, u2_N340, u2_N341, u2_N344, u2_N346, u2_N351, u2_N352, 
      u2_N356, u2_N357, u2_N360, u2_N361, u2_N366, u2_N367, u2_N368, u2_N371, u2_N372, 
      u2_N374, u2_N375, u2_N377, u2_N378, u2_N381, u2_N382, u2_N384, u2_N385, u2_N386, 
      u2_N387, u2_N388, u2_N389, u2_N390, u2_N391, u2_N392, u2_N393, u2_N394, u2_N395, 
      u2_N396, u2_N397, u2_N398, u2_N399, u2_N400, u2_N401, u2_N402, u2_N403, u2_N404, 
      u2_N405, u2_N406, u2_N407, u2_N408, u2_N409, u2_N413, u2_N414, u2_N415, u2_N417, 
      u2_N420, u2_N421, u2_N424, u2_N428, u2_N430, u2_N431, u2_N432, u2_N433, u2_N436, 
      u2_N438, u2_N439, u2_N442, u2_N443, u2_N445, u2_N446, u2_N449, u2_N453, u2_N460, 
      u2_N463, u2_N465, u2_N471, u2_N475, u2_N477, u2_out0_1, u2_out0_10, u2_out0_11, u2_out0_12, 
      u2_out0_13, u2_out0_14, u2_out0_15, u2_out0_16, u2_out0_17, u2_out0_18, u2_out0_19, u2_out0_2, u2_out0_20, 
      u2_out0_21, u2_out0_22, u2_out0_23, u2_out0_24, u2_out0_25, u2_out0_26, u2_out0_27, u2_out0_28, u2_out0_29, 
      u2_out0_3, u2_out0_30, u2_out0_31, u2_out0_32, u2_out0_4, u2_out0_5, u2_out0_6, u2_out0_7, u2_out0_8, 
      u2_out0_9, u2_out10_1, u2_out10_10, u2_out10_11, u2_out10_13, u2_out10_16, u2_out10_17, u2_out10_18, u2_out10_19, 
      u2_out10_2, u2_out10_20, u2_out10_23, u2_out10_24, u2_out10_26, u2_out10_28, u2_out10_29, u2_out10_30, u2_out10_31, 
      u2_out10_4, u2_out10_6, u2_out10_9, u2_out11_11, u2_out11_12, u2_out11_13, u2_out11_14, u2_out11_18, u2_out11_19, 
      u2_out11_2, u2_out11_22, u2_out11_25, u2_out11_28, u2_out11_29, u2_out11_3, u2_out11_32, u2_out11_4, u2_out11_7, 
      u2_out11_8, u2_out12_27, u2_out12_28, u2_out12_29, u2_out13_1, u2_out13_10, u2_out13_11, u2_out13_12, u2_out13_14, 
      u2_out13_19, u2_out13_20, u2_out13_22, u2_out13_25, u2_out13_26, u2_out13_29, u2_out13_3, u2_out13_32, u2_out13_4, 
      u2_out13_7, u2_out13_8, u2_out14_1, u2_out14_10, u2_out14_11, u2_out14_12, u2_out14_14, u2_out14_15, u2_out14_17, 
      u2_out14_19, u2_out14_20, u2_out14_21, u2_out14_22, u2_out14_23, u2_out14_25, u2_out14_26, u2_out14_27, u2_out14_29, 
      u2_out14_3, u2_out14_31, u2_out14_32, u2_out14_4, u2_out14_5, u2_out14_7, u2_out14_8, u2_out14_9, u2_out15_1, 
      u2_out15_10, u2_out15_13, u2_out15_14, u2_out15_16, u2_out15_17, u2_out15_18, u2_out15_2, u2_out15_20, u2_out15_23, 
      u2_out15_24, u2_out15_25, u2_out15_26, u2_out15_28, u2_out15_3, u2_out15_30, u2_out15_31, u2_out15_6, u2_out15_8, 
      u2_out15_9, u2_out1_1, u2_out1_10, u2_out1_11, u2_out1_12, u2_out1_13, u2_out1_14, u2_out1_15, u2_out1_16, 
      u2_out1_17, u2_out1_18, u2_out1_19, u2_out1_2, u2_out1_20, u2_out1_21, u2_out1_22, u2_out1_23, u2_out1_24, 
      u2_out1_25, u2_out1_26, u2_out1_27, u2_out1_28, u2_out1_29, u2_out1_3, u2_out1_30, u2_out1_31, u2_out1_32, 
      u2_out1_4, u2_out1_5, u2_out1_6, u2_out1_7, u2_out1_8, u2_out1_9, u2_out2_1, u2_out2_10, u2_out2_11, 
      u2_out2_12, u2_out2_13, u2_out2_14, u2_out2_15, u2_out2_16, u2_out2_17, u2_out2_18, u2_out2_19, u2_out2_2, 
      u2_out2_20, u2_out2_21, u2_out2_22, u2_out2_23, u2_out2_24, u2_out2_25, u2_out2_26, u2_out2_27, u2_out2_28, 
      u2_out2_29, u2_out2_3, u2_out2_30, u2_out2_31, u2_out2_32, u2_out2_4, u2_out2_5, u2_out2_6, u2_out2_7, 
      u2_out2_8, u2_out2_9, u2_out3_1, u2_out3_10, u2_out3_11, u2_out3_12, u2_out3_13, u2_out3_14, u2_out3_15, 
      u2_out3_16, u2_out3_17, u2_out3_18, u2_out3_19, u2_out3_2, u2_out3_20, u2_out3_21, u2_out3_22, u2_out3_23, 
      u2_out3_24, u2_out3_25, u2_out3_26, u2_out3_27, u2_out3_28, u2_out3_29, u2_out3_3, u2_out3_30, u2_out3_31, 
      u2_out3_32, u2_out3_4, u2_out3_5, u2_out3_6, u2_out3_7, u2_out3_8, u2_out3_9, u2_out4_1, u2_out4_10, 
      u2_out4_11, u2_out4_12, u2_out4_13, u2_out4_14, u2_out4_15, u2_out4_16, u2_out4_17, u2_out4_18, u2_out4_19, 
      u2_out4_2, u2_out4_20, u2_out4_21, u2_out4_22, u2_out4_23, u2_out4_24, u2_out4_25, u2_out4_26, u2_out4_27, 
      u2_out4_28, u2_out4_29, u2_out4_3, u2_out4_30, u2_out4_31, u2_out4_32, u2_out4_4, u2_out4_5, u2_out4_6, 
      u2_out4_7, u2_out4_8, u2_out4_9, u2_out5_1, u2_out5_10, u2_out5_11, u2_out5_12, u2_out5_13, u2_out5_14, 
      u2_out5_15, u2_out5_16, u2_out5_17, u2_out5_18, u2_out5_19, u2_out5_2, u2_out5_20, u2_out5_21, u2_out5_22, 
      u2_out5_23, u2_out5_24, u2_out5_25, u2_out5_26, u2_out5_27, u2_out5_28, u2_out5_29, u2_out5_3, u2_out5_30, 
      u2_out5_31, u2_out5_32, u2_out5_4, u2_out5_5, u2_out5_6, u2_out5_7, u2_out5_8, u2_out5_9, u2_out6_1, 
      u2_out6_10, u2_out6_11, u2_out6_12, u2_out6_13, u2_out6_14, u2_out6_15, u2_out6_16, u2_out6_17, u2_out6_18, 
      u2_out6_19, u2_out6_2, u2_out6_20, u2_out6_21, u2_out6_22, u2_out6_23, u2_out6_24, u2_out6_25, u2_out6_26, 
      u2_out6_27, u2_out6_28, u2_out6_29, u2_out6_3, u2_out6_30, u2_out6_31, u2_out6_32, u2_out6_4, u2_out6_5, 
      u2_out6_6, u2_out6_7, u2_out6_8, u2_out6_9, u2_out7_1, u2_out7_10, u2_out7_12, u2_out7_13, u2_out7_16, 
      u2_out7_17, u2_out7_18, u2_out7_2, u2_out7_20, u2_out7_23, u2_out7_24, u2_out7_26, u2_out7_28, u2_out7_30, 
      u2_out7_31, u2_out7_6, u2_out7_9, u2_out8_1, u2_out8_10, u2_out8_13, u2_out8_14, u2_out8_16, u2_out8_18, 
      u2_out8_2, u2_out8_20, u2_out8_24, u2_out8_25, u2_out8_26, u2_out8_28, u2_out8_3, u2_out8_30, u2_out8_6, 
      u2_out8_8, u2_out9_1, u2_out9_10, u2_out9_11, u2_out9_12, u2_out9_13, u2_out9_14, u2_out9_15, u2_out9_16, 
      u2_out9_17, u2_out9_18, u2_out9_19, u2_out9_2, u2_out9_20, u2_out9_21, u2_out9_22, u2_out9_23, u2_out9_24, 
      u2_out9_25, u2_out9_26, u2_out9_27, u2_out9_28, u2_out9_29, u2_out9_3, u2_out9_30, u2_out9_31, u2_out9_32, 
      u2_out9_4, u2_out9_5, u2_out9_6, u2_out9_7, u2_out9_8, u2_out9_9, u2_uk_n10, u2_uk_n100, u2_uk_n102, 
      u2_uk_n109, u2_uk_n11, u2_uk_n110, u2_uk_n1142, u2_uk_n1146, u2_uk_n1152, u2_uk_n1161, u2_uk_n1167, u2_uk_n1168, 
      u2_uk_n117, u2_uk_n1171, u2_uk_n1178, u2_uk_n1179, u2_uk_n118, u2_uk_n128, u2_uk_n129, u2_uk_n141, u2_uk_n142, 
      u2_uk_n145, u2_uk_n146, u2_uk_n147, u2_uk_n148, u2_uk_n155, u2_uk_n161, u2_uk_n162, u2_uk_n163, u2_uk_n164, 
      u2_uk_n17, u2_uk_n182, u2_uk_n187, u2_uk_n188, u2_uk_n191, u2_uk_n202, u2_uk_n203, u2_uk_n207, u2_uk_n208, 
      u2_uk_n209, u2_uk_n213, u2_uk_n214, u2_uk_n217, u2_uk_n220, u2_uk_n222, u2_uk_n223, u2_uk_n230, u2_uk_n231, 
      u2_uk_n27, u2_uk_n31, u2_uk_n60, u2_uk_n63, u2_uk_n83, u2_uk_n92, u2_uk_n93, u2_uk_n94, u2_uk_n99, 
      n116, u0_FP_33, u0_FP_34, u0_FP_36, u0_FP_37, u0_FP_38, u0_FP_39, u0_FP_40, u0_FP_41, 
      u0_FP_42, u0_FP_43, u0_FP_45, u0_FP_48, u0_FP_49, u0_FP_50, u0_FP_51, u0_FP_52, u0_FP_53, 
      u0_FP_54, u0_FP_55, u0_FP_56, u0_FP_57, u0_FP_58, u0_FP_59, u0_FP_60, u0_FP_61, u0_FP_62, 
      u0_FP_63, u0_FP_64, u0_K10_10, u0_K10_13, u0_K10_14, u0_K10_18, u0_K10_19, u0_K10_20, u0_K10_25, 
      u0_K10_32, u0_K10_36, u0_K11_25, u0_K11_37, u0_K11_48, u0_K12_19, u0_K12_22, u0_K12_34, u0_K12_35, 
      u0_K12_36, u0_K12_39, u0_K12_40, u0_K12_48, u0_K12_7, u0_K12_9, u0_K13_30, u0_K13_36, u0_K13_38, 
      u0_K13_8, u0_K14_10, u0_K14_12, u0_K14_13, u0_K14_14, u0_K14_15, u0_K14_18, u0_K14_23, u0_K14_4, 
      u0_K14_42, u0_K14_9, u0_K15_18, u0_K15_47, u0_K16_11, u0_K16_18, u0_K16_24, u0_K16_26, u0_K16_38, 
      u0_K16_8, u0_K1_13, u0_K1_14, u0_K1_17, u0_K1_31, u0_K1_47, u0_K2_17, u0_K2_30, u0_K2_44, 
      u0_K2_5, u0_K2_6, u0_K2_8, u0_K3_12, u0_K3_13, u0_K3_14, u0_K3_17, u0_K3_18, u0_K3_19, 
      u0_K3_23, u0_K3_5, u0_K3_6, u0_K4_24, u0_K4_43, u0_K4_48, u0_K5_1, u0_K5_13, u0_K5_14, 
      u0_K5_15, u0_K5_16, u0_K5_18, u0_K5_19, u0_K5_23, u0_K5_24, u0_K5_26, u0_K5_28, u0_K5_3, 
      u0_K5_31, u0_K5_32, u0_K5_4, u0_K5_41, u0_K5_44, u0_K5_47, u0_K5_48, u0_K5_9, u0_K6_11, 
      u0_K6_13, u0_K6_20, u0_K6_23, u0_K7_2, u0_K7_23, u0_K8_1, u0_K8_11, u0_K8_13, u0_K8_19, 
      u0_K8_23, u0_K9_14, u0_K9_15, u0_K9_32, u0_K9_39, u0_K9_4, u0_K9_40, u0_K9_45, u0_K9_6, 
      u0_L10_1, u0_L10_10, u0_L10_11, u0_L10_12, u0_L10_13, u0_L10_14, u0_L10_15, u0_L10_16, u0_L10_17, 
      u0_L10_18, u0_L10_19, u0_L10_2, u0_L10_20, u0_L10_21, u0_L10_22, u0_L10_23, u0_L10_24, u0_L10_25, 
      u0_L10_26, u0_L10_27, u0_L10_28, u0_L10_29, u0_L10_3, u0_L10_30, u0_L10_31, u0_L10_32, u0_L10_4, 
      u0_L10_5, u0_L10_6, u0_L10_7, u0_L10_8, u0_L10_9, u0_L12_13, u0_L12_16, u0_L12_17, u0_L12_18, 
      u0_L12_2, u0_L12_23, u0_L12_24, u0_L12_28, u0_L12_30, u0_L12_31, u0_L12_6, u0_L12_9, u0_L13_1, 
      u0_L13_10, u0_L13_13, u0_L13_18, u0_L13_2, u0_L13_20, u0_L13_26, u0_L13_28, u0_L14_11, u0_L14_12, 
      u0_L14_14, u0_L14_15, u0_L14_19, u0_L14_21, u0_L14_22, u0_L14_25, u0_L14_27, u0_L14_29, u0_L14_3, 
      u0_L14_32, u0_L14_4, u0_L14_5, u0_L14_7, u0_L14_8, u0_L3_1, u0_L3_10, u0_L3_13, u0_L3_14, 
      u0_L3_15, u0_L3_16, u0_L3_17, u0_L3_18, u0_L3_2, u0_L3_20, u0_L3_21, u0_L3_23, u0_L3_24, 
      u0_L3_25, u0_L3_26, u0_L3_27, u0_L3_28, u0_L3_3, u0_L3_30, u0_L3_31, u0_L3_5, u0_L3_6, 
      u0_L3_8, u0_L3_9, u0_L7_1, u0_L7_10, u0_L7_11, u0_L7_12, u0_L7_13, u0_L7_14, u0_L7_15, 
      u0_L7_16, u0_L7_17, u0_L7_18, u0_L7_19, u0_L7_2, u0_L7_20, u0_L7_21, u0_L7_22, u0_L7_23, 
      u0_L7_24, u0_L7_25, u0_L7_26, u0_L7_27, u0_L7_28, u0_L7_29, u0_L7_3, u0_L7_30, u0_L7_31, 
      u0_L7_32, u0_L7_4, u0_L7_5, u0_L7_6, u0_L7_7, u0_L7_8, u0_L7_9, u0_L8_1, u0_L8_10, 
      u0_L8_13, u0_L8_16, u0_L8_17, u0_L8_18, u0_L8_2, u0_L8_20, u0_L8_23, u0_L8_24, u0_L8_26, 
      u0_L8_28, u0_L8_30, u0_L8_31, u0_L8_6, u0_L8_9, u0_R0_12, u0_R0_14, u0_R0_17, u0_R0_18, 
      u0_R0_19, u0_R0_21, u0_R0_22, u0_R0_25, u0_R0_27, u0_R0_28, u0_R0_29, u0_R0_4, u0_R0_5, 
      u0_R10_1, u0_R10_10, u0_R10_11, u0_R10_12, u0_R10_13, u0_R10_14, u0_R10_15, u0_R10_16, u0_R10_17, 
      u0_R10_18, u0_R10_19, u0_R10_2, u0_R10_20, u0_R10_21, u0_R10_22, u0_R10_23, u0_R10_24, u0_R10_25, 
      u0_R10_26, u0_R10_27, u0_R10_28, u0_R10_29, u0_R10_3, u0_R10_30, u0_R10_31, u0_R10_32, u0_R10_4, 
      u0_R10_5, u0_R10_6, u0_R10_7, u0_R10_8, u0_R10_9, u0_R11_10, u0_R11_11, u0_R11_12, u0_R11_13, 
      u0_R11_14, u0_R11_15, u0_R11_16, u0_R11_17, u0_R11_20, u0_R11_21, u0_R11_22, u0_R11_23, u0_R11_24, 
      u0_R11_25, u0_R11_28, u0_R11_3, u0_R11_32, u0_R11_4, u0_R11_5, u0_R11_6, u0_R11_7, u0_R11_8, 
      u0_R11_9, u0_R12_1, u0_R12_10, u0_R12_11, u0_R12_12, u0_R12_13, u0_R12_16, u0_R12_19, u0_R12_2, 
      u0_R12_20, u0_R12_21, u0_R12_22, u0_R12_23, u0_R12_24, u0_R12_25, u0_R12_26, u0_R12_28, u0_R12_29, 
      u0_R12_3, u0_R12_30, u0_R12_32, u0_R12_4, u0_R12_5, u0_R12_6, u0_R12_7, u0_R12_8, u0_R12_9, 
      u0_R13_1, u0_R13_11, u0_R13_12, u0_R13_13, u0_R13_14, u0_R13_15, u0_R13_16, u0_R13_17, u0_R13_18, 
      u0_R13_19, u0_R13_2, u0_R13_20, u0_R13_21, u0_R13_22, u0_R13_23, u0_R13_24, u0_R13_25, u0_R13_26, 
      u0_R13_27, u0_R13_28, u0_R13_29, u0_R13_3, u0_R13_30, u0_R13_31, u0_R13_32, u0_R13_4, u0_R13_5, 
      u0_R13_6, u0_R13_7, u0_R13_8, u0_R13_9, u0_R1_1, u0_R1_12, u0_R1_13, u0_R1_16, u0_R1_17, 
      u0_R1_18, u0_R1_19, u0_R1_20, u0_R1_21, u0_R1_22, u0_R1_24, u0_R1_25, u0_R1_26, u0_R1_27, 
      u0_R1_28, u0_R1_29, u0_R1_3, u0_R1_31, u0_R1_32, u0_R1_4, u0_R1_5, u0_R1_8, u0_R1_9, 
      u0_R2_1, u0_R2_10, u0_R2_11, u0_R2_12, u0_R2_13, u0_R2_14, u0_R2_15, u0_R2_16, u0_R2_17, 
      u0_R2_20, u0_R2_21, u0_R2_22, u0_R2_23, u0_R2_26, u0_R2_27, u0_R2_28, u0_R2_29, u0_R2_3, 
      u0_R2_30, u0_R2_31, u0_R2_32, u0_R2_4, u0_R2_6, u0_R2_7, u0_R2_8, u0_R2_9, u0_R3_1, 
      u0_R3_10, u0_R3_11, u0_R3_12, u0_R3_13, u0_R3_14, u0_R3_15, u0_R3_16, u0_R3_17, u0_R3_18, 
      u0_R3_19, u0_R3_2, u0_R3_20, u0_R3_21, u0_R3_22, u0_R3_24, u0_R3_27, u0_R3_28, u0_R3_29, 
      u0_R3_3, u0_R3_30, u0_R3_31, u0_R3_32, u0_R3_4, u0_R3_5, u0_R3_6, u0_R3_7, u0_R3_8, 
      u0_R3_9, u0_R4_1, u0_R4_13, u0_R4_14, u0_R4_16, u0_R4_22, u0_R4_24, u0_R4_29, u0_R4_30, 
      u0_R4_8, u0_R5_1, u0_R5_11, u0_R5_12, u0_R5_13, u0_R5_14, u0_R5_16, u0_R5_17, u0_R5_18, 
      u0_R5_19, u0_R5_2, u0_R5_20, u0_R5_21, u0_R5_22, u0_R5_23, u0_R5_24, u0_R5_25, u0_R5_26, 
      u0_R5_27, u0_R5_28, u0_R5_29, u0_R5_3, u0_R5_30, u0_R5_31, u0_R5_32, u0_R5_4, u0_R5_5, 
      u0_R5_7, u0_R5_8, u0_R5_9, u0_R6_1, u0_R6_10, u0_R6_11, u0_R6_12, u0_R6_13, u0_R6_14, 
      u0_R6_16, u0_R6_17, u0_R6_18, u0_R6_2, u0_R6_20, u0_R6_21, u0_R6_23, u0_R6_24, u0_R6_26, 
      u0_R6_27, u0_R6_28, u0_R6_29, u0_R6_32, u0_R6_4, u0_R6_5, u0_R6_7, u0_R6_8, u0_R6_9, 
      u0_R7_1, u0_R7_10, u0_R7_11, u0_R7_12, u0_R7_13, u0_R7_14, u0_R7_15, u0_R7_16, u0_R7_17, 
      u0_R7_18, u0_R7_19, u0_R7_2, u0_R7_20, u0_R7_21, u0_R7_22, u0_R7_23, u0_R7_24, u0_R7_25, 
      u0_R7_26, u0_R7_27, u0_R7_28, u0_R7_29, u0_R7_3, u0_R7_30, u0_R7_31, u0_R7_32, u0_R7_4, 
      u0_R7_5, u0_R7_6, u0_R7_7, u0_R7_8, u0_R7_9, u0_R8_1, u0_R8_10, u0_R8_11, u0_R8_12, 
      u0_R8_13, u0_R8_14, u0_R8_15, u0_R8_16, u0_R8_17, u0_R8_19, u0_R8_2, u0_R8_20, u0_R8_21, 
      u0_R8_22, u0_R8_24, u0_R8_25, u0_R8_27, u0_R8_29, u0_R8_3, u0_R8_30, u0_R8_32, u0_R8_4, 
      u0_R8_5, u0_R8_6, u0_R8_7, u0_R8_8, u0_R8_9, u0_R9_1, u0_R9_10, u0_R9_11, u0_R9_12, 
      u0_R9_13, u0_R9_15, u0_R9_16, u0_R9_17, u0_R9_18, u0_R9_19, u0_R9_2, u0_R9_20, u0_R9_21, 
      u0_R9_22, u0_R9_23, u0_R9_24, u0_R9_25, u0_R9_27, u0_R9_28, u0_R9_29, u0_R9_3, u0_R9_31, 
      u0_R9_32, u0_R9_4, u0_R9_5, u0_R9_6, u0_R9_7, u0_R9_8, u0_R9_9, u0_desIn_r_1, u0_desIn_r_11, 
      u0_desIn_r_15, u0_desIn_r_25, u0_desIn_r_27, u0_desIn_r_29, u0_desIn_r_3, u0_desIn_r_31, u0_desIn_r_33, u0_desIn_r_37, u0_desIn_r_39, 
      u0_desIn_r_45, u0_desIn_r_47, u0_desIn_r_5, u0_desIn_r_51, u0_desIn_r_53, u0_desIn_r_55, u0_desIn_r_57, u0_desIn_r_59, u0_desIn_r_63, 
      u0_desIn_r_7, u0_key_r_11, u0_key_r_12, u0_key_r_13, u0_key_r_14, u0_key_r_16, u0_key_r_17, u0_key_r_19, u0_key_r_2, 
      u0_key_r_20, u0_key_r_21, u0_key_r_23, u0_key_r_24, u0_key_r_25, u0_key_r_26, u0_key_r_27, u0_key_r_28, u0_key_r_30, 
      u0_key_r_31, u0_key_r_32, u0_key_r_34, u0_key_r_35, u0_key_r_36, u0_key_r_37, u0_key_r_38, u0_key_r_39, u0_key_r_4, 
      u0_key_r_40, u0_key_r_41, u0_key_r_42, u0_key_r_43, u0_key_r_47, u0_key_r_48, u0_key_r_5, u0_key_r_50, u0_key_r_51, 
      u0_key_r_54, u0_key_r_55, u0_key_r_6, u0_key_r_9, u0_u0_X_15, u0_u0_X_16, u0_u0_X_23, u0_u0_X_25, u0_u0_X_28, 
      u0_u0_X_30, u0_u0_X_32, u0_u0_X_33, u0_u0_X_39, u0_u0_X_4, u0_u0_X_40, u0_u0_X_45, u0_u0_X_46, u0_u10_X_21, 
      u0_u10_X_39, u0_u10_X_45, u0_u12_X_2, u0_u12_X_27, u0_u12_X_28, u0_u12_X_3, u0_u12_X_39, u0_u12_X_40, u0_u12_X_42, 
      u0_u12_X_44, u0_u12_X_45, u0_u12_X_46, u0_u12_X_48, u0_u13_X_21, u0_u13_X_22, u0_u13_X_24, u0_u13_X_26, u0_u13_X_27, 
      u0_u13_X_40, u0_u13_X_46, u0_u14_X_15, u0_u15_X_17, u0_u15_X_19, u0_u15_X_21, u0_u15_X_22, u0_u15_X_4, u0_u1_X_1, 
      u0_u1_X_10, u0_u1_X_11, u0_u1_X_12, u0_u1_X_13, u0_u1_X_14, u0_u1_X_15, u0_u1_X_16, u0_u1_X_18, u0_u1_X_2, 
      u0_u1_X_20, u0_u1_X_22, u0_u1_X_23, u0_u1_X_25, u0_u1_X_29, u0_u1_X_3, u0_u1_X_31, u0_u1_X_34, u0_u1_X_35, 
      u0_u1_X_37, u0_u1_X_39, u0_u1_X_4, u0_u1_X_45, u0_u1_X_46, u0_u1_X_47, u0_u1_X_48, u0_u1_X_9, u0_u2_X_10, 
      u0_u2_X_15, u0_u2_X_16, u0_u2_X_21, u0_u2_X_22, u0_u2_X_3, u0_u2_X_34, u0_u2_X_45, u0_u2_X_9, u0_u3_X_27, 
      u0_u3_X_28, u0_u3_X_3, u0_u3_X_35, u0_u3_X_36, u0_u3_X_37, u0_u3_X_38, u0_u3_X_6, u0_u3_X_8, u0_u4_X_34, 
      u0_u4_X_36, u0_u4_X_38, u0_u4_X_39, u0_u5_X_1, u0_u5_X_10, u0_u5_X_12, u0_u5_X_14, u0_u5_X_15, u0_u5_X_16, 
      u0_u5_X_17, u0_u5_X_19, u0_u5_X_22, u0_u5_X_24, u0_u5_X_26, u0_u5_X_27, u0_u5_X_28, u0_u5_X_29, u0_u5_X_3, 
      u0_u5_X_30, u0_u5_X_31, u0_u5_X_32, u0_u5_X_34, u0_u5_X_36, u0_u5_X_38, u0_u5_X_39, u0_u5_X_4, u0_u5_X_40, 
      u0_u5_X_41, u0_u5_X_43, u0_u5_X_46, u0_u5_X_47, u0_u5_X_5, u0_u5_X_6, u0_u5_X_7, u0_u5_X_8, u0_u5_X_9, 
      u0_u6_X_15, u0_u6_X_22, u0_u6_X_9, u0_u7_X_22, u0_u7_X_28, u0_u7_X_33, u0_u7_X_36, u0_u7_X_38, u0_u7_X_4, 
      u0_u7_X_45, u0_u7_X_46, u0_u7_X_9, u0_u9_X_27, u0_u9_X_34, u0_u9_X_39, u0_u9_X_41, u0_u9_X_43, u0_u9_X_46, 
      u0_uk_K_r0_15, u0_uk_K_r0_2, u0_uk_K_r0_28, u0_uk_K_r0_31, u0_uk_K_r0_36, u0_uk_K_r0_49, u0_uk_K_r0_7, u0_uk_K_r10_10, u0_uk_K_r10_14, 
      u0_uk_K_r10_18, u0_uk_K_r10_23, u0_uk_K_r10_25, u0_uk_K_r10_27, u0_uk_K_r10_28, u0_uk_K_r10_32, u0_uk_K_r10_34, u0_uk_K_r10_37, u0_uk_K_r10_39, 
      u0_uk_K_r10_41, u0_uk_K_r10_42, u0_uk_K_r10_43, u0_uk_K_r10_44, u0_uk_K_r10_47, u0_uk_K_r10_48, u0_uk_K_r10_9, u0_uk_K_r11_11, u0_uk_K_r11_17, 
      u0_uk_K_r11_20, u0_uk_K_r11_25, u0_uk_K_r11_27, u0_uk_K_r11_29, u0_uk_K_r11_33, u0_uk_K_r11_34, u0_uk_K_r11_48, u0_uk_K_r11_53, u0_uk_K_r11_54, 
      u0_uk_K_r11_6, u0_uk_K_r12_10, u0_uk_K_r12_15, u0_uk_K_r12_16, u0_uk_K_r12_25, u0_uk_K_r12_33, u0_uk_K_r12_44, u0_uk_K_r12_47, u0_uk_K_r13_0, 
      u0_uk_K_r13_13, u0_uk_K_r13_17, u0_uk_K_r13_22, u0_uk_K_r13_25, u0_uk_K_r13_32, u0_uk_K_r13_35, u0_uk_K_r13_38, u0_uk_K_r13_4, u0_uk_K_r13_44, 
      u0_uk_K_r13_55, u0_uk_K_r14_11, u0_uk_K_r14_12, u0_uk_K_r14_15, u0_uk_K_r14_16, u0_uk_K_r14_18, u0_uk_K_r14_2, u0_uk_K_r14_43, u0_uk_K_r14_45, 
      u0_uk_K_r14_46, u0_uk_K_r14_50, u0_uk_K_r14_8, u0_uk_K_r14_9, u0_uk_K_r1_15, u0_uk_K_r1_21, u0_uk_K_r1_22, u0_uk_K_r1_42, u0_uk_K_r1_44, 
      u0_uk_K_r1_7, u0_uk_K_r2_13, u0_uk_K_r2_18, u0_uk_K_r2_20, u0_uk_K_r2_25, u0_uk_K_r2_27, u0_uk_K_r2_28, u0_uk_K_r2_33, u0_uk_K_r2_53, 
      u0_uk_K_r2_55, u0_uk_K_r3_10, u0_uk_K_r3_11, u0_uk_K_r3_14, u0_uk_K_r3_15, u0_uk_K_r3_19, u0_uk_K_r3_24, u0_uk_K_r3_35, u0_uk_K_r3_38, 
      u0_uk_K_r3_47, u0_uk_K_r3_9, u0_uk_K_r4_38, u0_uk_K_r5_10, u0_uk_K_r5_16, u0_uk_K_r5_17, u0_uk_K_r5_19, u0_uk_K_r5_32, u0_uk_K_r5_37, 
      u0_uk_K_r5_39, u0_uk_K_r5_4, u0_uk_K_r5_8, u0_uk_K_r6_0, u0_uk_K_r6_10, u0_uk_K_r6_14, u0_uk_K_r6_21, u0_uk_K_r6_22, u0_uk_K_r6_26, 
      u0_uk_K_r6_27, u0_uk_K_r6_29, u0_uk_K_r6_3, u0_uk_K_r6_31, u0_uk_K_r6_34, u0_uk_K_r6_46, u0_uk_K_r6_53, u0_uk_K_r6_7, u0_uk_K_r7_0, 
      u0_uk_K_r7_1, u0_uk_K_r7_13, u0_uk_K_r7_15, u0_uk_K_r7_2, u0_uk_K_r7_20, u0_uk_K_r7_22, u0_uk_K_r7_23, u0_uk_K_r7_24, u0_uk_K_r7_25, 
      u0_uk_K_r7_26, u0_uk_K_r7_27, u0_uk_K_r7_30, u0_uk_K_r7_32, u0_uk_K_r7_39, u0_uk_K_r7_48, u0_uk_K_r7_55, u0_uk_K_r7_6, u0_uk_K_r7_8, 
      u0_uk_K_r7_9, u0_uk_K_r8_13, u0_uk_K_r8_16, u0_uk_K_r8_17, u0_uk_K_r8_2, u0_uk_K_r8_22, u0_uk_K_r8_27, u0_uk_K_r8_32, u0_uk_K_r8_37, 
      u0_uk_K_r8_40, u0_uk_K_r8_41, u0_uk_K_r9_0, u0_uk_K_r9_1, u0_uk_K_r9_13, u0_uk_K_r9_19, u0_uk_K_r9_25, u0_uk_K_r9_27, u0_uk_K_r9_31, 
      u0_uk_K_r9_33, u0_uk_K_r9_35, u0_uk_K_r9_45, u0_uk_K_r9_49, u0_uk_K_r9_6, u0_uk_K_r9_9, u0_uk_n1, u0_uk_n1000, u0_uk_n1001, 
      u0_uk_n1002, u0_uk_n1004, u0_uk_n1008, u0_uk_n1009, u0_uk_n1012, u0_uk_n1019, u0_uk_n1020, u0_uk_n1021, u0_uk_n1024, 
      u0_uk_n104, u0_uk_n106, u0_uk_n108, u0_uk_n112, u0_uk_n113, u0_uk_n115, u0_uk_n116, u0_uk_n12, u0_uk_n120, 
      u0_uk_n121, u0_uk_n122, u0_uk_n123, u0_uk_n124, u0_uk_n126, u0_uk_n127, u0_uk_n13, u0_uk_n130, u0_uk_n131, 
      u0_uk_n132, u0_uk_n135, u0_uk_n136, u0_uk_n137, u0_uk_n139, u0_uk_n14, u0_uk_n140, u0_uk_n143, u0_uk_n144, 
      u0_uk_n149, u0_uk_n15, u0_uk_n150, u0_uk_n151, u0_uk_n152, u0_uk_n153, u0_uk_n154, u0_uk_n156, u0_uk_n157, 
      u0_uk_n159, u0_uk_n16, u0_uk_n165, u0_uk_n166, u0_uk_n167, u0_uk_n168, u0_uk_n169, u0_uk_n170, u0_uk_n171, 
      u0_uk_n172, u0_uk_n173, u0_uk_n174, u0_uk_n175, u0_uk_n176, u0_uk_n177, u0_uk_n178, u0_uk_n179, u0_uk_n18, 
      u0_uk_n180, u0_uk_n181, u0_uk_n183, u0_uk_n184, u0_uk_n185, u0_uk_n186, u0_uk_n189, u0_uk_n19, u0_uk_n190, 
      u0_uk_n193, u0_uk_n194, u0_uk_n195, u0_uk_n196, u0_uk_n197, u0_uk_n198, u0_uk_n199, u0_uk_n20, u0_uk_n200, 
      u0_uk_n201, u0_uk_n204, u0_uk_n205, u0_uk_n206, u0_uk_n21, u0_uk_n210, u0_uk_n212, u0_uk_n215, u0_uk_n216, 
      u0_uk_n218, u0_uk_n219, u0_uk_n22, u0_uk_n221, u0_uk_n224, u0_uk_n225, u0_uk_n226, u0_uk_n227, u0_uk_n228, 
      u0_uk_n229, u0_uk_n23, u0_uk_n232, u0_uk_n233, u0_uk_n234, u0_uk_n235, u0_uk_n239, u0_uk_n24, u0_uk_n241, 
      u0_uk_n243, u0_uk_n244, u0_uk_n245, u0_uk_n246, u0_uk_n248, u0_uk_n249, u0_uk_n25, u0_uk_n253, u0_uk_n254, 
      u0_uk_n255, u0_uk_n257, u0_uk_n258, u0_uk_n259, u0_uk_n26, u0_uk_n260, u0_uk_n261, u0_uk_n262, u0_uk_n263, 
      u0_uk_n264, u0_uk_n266, u0_uk_n267, u0_uk_n268, u0_uk_n269, u0_uk_n272, u0_uk_n273, u0_uk_n274, u0_uk_n275, 
      u0_uk_n276, u0_uk_n278, u0_uk_n28, u0_uk_n280, u0_uk_n281, u0_uk_n282, u0_uk_n283, u0_uk_n285, u0_uk_n288, 
      u0_uk_n289, u0_uk_n29, u0_uk_n290, u0_uk_n293, u0_uk_n296, u0_uk_n3, u0_uk_n30, u0_uk_n300, u0_uk_n303, 
      u0_uk_n304, u0_uk_n307, u0_uk_n309, u0_uk_n310, u0_uk_n311, u0_uk_n314, u0_uk_n315, u0_uk_n316, u0_uk_n318, 
      u0_uk_n32, u0_uk_n320, u0_uk_n321, u0_uk_n324, u0_uk_n325, u0_uk_n327, u0_uk_n329, u0_uk_n33, u0_uk_n330, 
      u0_uk_n331, u0_uk_n332, u0_uk_n333, u0_uk_n336, u0_uk_n337, u0_uk_n339, u0_uk_n34, u0_uk_n341, u0_uk_n343, 
      u0_uk_n344, u0_uk_n347, u0_uk_n348, u0_uk_n35, u0_uk_n352, u0_uk_n354, u0_uk_n355, u0_uk_n358, u0_uk_n359, 
      u0_uk_n36, u0_uk_n361, u0_uk_n362, u0_uk_n365, u0_uk_n367, u0_uk_n368, u0_uk_n37, u0_uk_n370, u0_uk_n371, 
      u0_uk_n372, u0_uk_n374, u0_uk_n378, u0_uk_n38, u0_uk_n380, u0_uk_n381, u0_uk_n383, u0_uk_n384, u0_uk_n387, 
      u0_uk_n388, u0_uk_n389, u0_uk_n39, u0_uk_n392, u0_uk_n393, u0_uk_n394, u0_uk_n396, u0_uk_n398, u0_uk_n399, 
      u0_uk_n4, u0_uk_n40, u0_uk_n400, u0_uk_n401, u0_uk_n402, u0_uk_n403, u0_uk_n405, u0_uk_n406, u0_uk_n41, 
      u0_uk_n412, u0_uk_n413, u0_uk_n418, u0_uk_n419, u0_uk_n42, u0_uk_n420, u0_uk_n425, u0_uk_n429, u0_uk_n43, 
      u0_uk_n430, u0_uk_n434, u0_uk_n44, u0_uk_n45, u0_uk_n451, u0_uk_n453, u0_uk_n455, u0_uk_n457, u0_uk_n458, 
      u0_uk_n459, u0_uk_n46, u0_uk_n462, u0_uk_n463, u0_uk_n464, u0_uk_n465, u0_uk_n466, u0_uk_n471, u0_uk_n473, 
      u0_uk_n475, u0_uk_n476, u0_uk_n479, u0_uk_n480, u0_uk_n481, u0_uk_n483, u0_uk_n484, u0_uk_n485, u0_uk_n486, 
      u0_uk_n488, u0_uk_n489, u0_uk_n490, u0_uk_n491, u0_uk_n493, u0_uk_n494, u0_uk_n497, u0_uk_n498, u0_uk_n499, 
      u0_uk_n5, u0_uk_n50, u0_uk_n502, u0_uk_n506, u0_uk_n508, u0_uk_n51, u0_uk_n510, u0_uk_n511, u0_uk_n513, 
      u0_uk_n514, u0_uk_n516, u0_uk_n517, u0_uk_n519, u0_uk_n52, u0_uk_n521, u0_uk_n522, u0_uk_n523, u0_uk_n525, 
      u0_uk_n528, u0_uk_n529, u0_uk_n53, u0_uk_n530, u0_uk_n531, u0_uk_n532, u0_uk_n534, u0_uk_n535, u0_uk_n536, 
      u0_uk_n537, u0_uk_n538, u0_uk_n539, u0_uk_n54, u0_uk_n543, u0_uk_n544, u0_uk_n545, u0_uk_n546, u0_uk_n547, 
      u0_uk_n549, u0_uk_n55, u0_uk_n550, u0_uk_n552, u0_uk_n553, u0_uk_n554, u0_uk_n555, u0_uk_n557, u0_uk_n558, 
      u0_uk_n559, u0_uk_n56, u0_uk_n560, u0_uk_n561, u0_uk_n562, u0_uk_n565, u0_uk_n566, u0_uk_n568, u0_uk_n57, 
      u0_uk_n570, u0_uk_n573, u0_uk_n574, u0_uk_n575, u0_uk_n578, u0_uk_n579, u0_uk_n58, u0_uk_n580, u0_uk_n581, 
      u0_uk_n584, u0_uk_n59, u0_uk_n592, u0_uk_n593, u0_uk_n599, u0_uk_n6, u0_uk_n600, u0_uk_n609, u0_uk_n61, 
      u0_uk_n612, u0_uk_n616, u0_uk_n62, u0_uk_n620, u0_uk_n623, u0_uk_n624, u0_uk_n629, u0_uk_n630, u0_uk_n631, 
      u0_uk_n632, u0_uk_n633, u0_uk_n635, u0_uk_n636, u0_uk_n637, u0_uk_n638, u0_uk_n639, u0_uk_n64, u0_uk_n640, 
      u0_uk_n641, u0_uk_n642, u0_uk_n643, u0_uk_n644, u0_uk_n645, u0_uk_n647, u0_uk_n648, u0_uk_n649, u0_uk_n65, 
      u0_uk_n650, u0_uk_n651, u0_uk_n652, u0_uk_n653, u0_uk_n655, u0_uk_n657, u0_uk_n658, u0_uk_n659, u0_uk_n660, 
      u0_uk_n663, u0_uk_n664, u0_uk_n666, u0_uk_n667, u0_uk_n668, u0_uk_n669, u0_uk_n67, u0_uk_n670, u0_uk_n68, 
      u0_uk_n69, u0_uk_n7, u0_uk_n719, u0_uk_n72, u0_uk_n720, u0_uk_n725, u0_uk_n726, u0_uk_n728, u0_uk_n73, 
      u0_uk_n731, u0_uk_n732, u0_uk_n735, u0_uk_n736, u0_uk_n739, u0_uk_n740, u0_uk_n746, u0_uk_n748, u0_uk_n75, 
      u0_uk_n755, u0_uk_n759, u0_uk_n763, u0_uk_n765, u0_uk_n766, u0_uk_n768, u0_uk_n77, u0_uk_n770, u0_uk_n771, 
      u0_uk_n774, u0_uk_n775, u0_uk_n776, u0_uk_n78, u0_uk_n780, u0_uk_n783, u0_uk_n793, u0_uk_n797, u0_uk_n799, 
      u0_uk_n8, u0_uk_n80, u0_uk_n805, u0_uk_n81, u0_uk_n810, u0_uk_n813, u0_uk_n815, u0_uk_n82, u0_uk_n826, 
      u0_uk_n828, u0_uk_n829, u0_uk_n831, u0_uk_n832, u0_uk_n834, u0_uk_n839, u0_uk_n84, u0_uk_n85, u0_uk_n851, 
      u0_uk_n855, u0_uk_n864, u0_uk_n87, u0_uk_n88, u0_uk_n89, u0_uk_n897, u0_uk_n898, u0_uk_n9, u0_uk_n90, 
      u0_uk_n904, u0_uk_n91, u0_uk_n915, u0_uk_n916, u0_uk_n917, u0_uk_n918, u0_uk_n933, u0_uk_n934, u0_uk_n939, 
      u0_uk_n940, u0_uk_n948, u0_uk_n949, u0_uk_n95, u0_uk_n950, u0_uk_n953, u0_uk_n96, u0_uk_n960, u0_uk_n963, 
      u0_uk_n98, u0_uk_n981, u0_uk_n982, u0_uk_n985, u0_uk_n990, u0_uk_n992, u0_uk_n999, u1_FP_33, u1_FP_34, 
      u1_FP_35, u1_FP_36, u1_FP_37, u1_FP_38, u1_FP_39, u1_FP_40, u1_FP_41, u1_FP_42, u1_FP_43, 
      u1_FP_44, u1_FP_45, u1_FP_46, u1_FP_47, u1_FP_48, u1_FP_49, u1_FP_50, u1_FP_51, u1_FP_52, 
      u1_FP_53, u1_FP_54, u1_FP_55, u1_FP_56, u1_FP_57, u1_FP_58, u1_FP_59, u1_FP_60, u1_FP_61, 
      u1_FP_62, u1_FP_63, u1_FP_64, u1_R0_1, u1_R0_10, u1_R0_11, u1_R0_12, u1_R0_13, u1_R0_14, 
      u1_R0_15, u1_R0_16, u1_R0_17, u1_R0_18, u1_R0_19, u1_R0_2, u1_R0_20, u1_R0_21, u1_R0_22, 
      u1_R0_23, u1_R0_24, u1_R0_25, u1_R0_26, u1_R0_27, u1_R0_28, u1_R0_29, u1_R0_3, u1_R0_30, 
      u1_R0_31, u1_R0_32, u1_R0_4, u1_R0_5, u1_R0_6, u1_R0_7, u1_R0_8, u1_R0_9, u1_R10_1, 
      u1_R10_10, u1_R10_11, u1_R10_12, u1_R10_13, u1_R10_14, u1_R10_15, u1_R10_16, u1_R10_17, u1_R10_18, 
      u1_R10_19, u1_R10_2, u1_R10_20, u1_R10_21, u1_R10_22, u1_R10_23, u1_R10_24, u1_R10_25, u1_R10_26, 
      u1_R10_27, u1_R10_28, u1_R10_29, u1_R10_3, u1_R10_30, u1_R10_31, u1_R10_32, u1_R10_4, u1_R10_5, 
      u1_R10_6, u1_R10_7, u1_R10_8, u1_R10_9, u1_R11_1, u1_R11_10, u1_R11_11, u1_R11_12, u1_R11_13, 
      u1_R11_14, u1_R11_15, u1_R11_16, u1_R11_17, u1_R11_18, u1_R11_19, u1_R11_2, u1_R11_20, u1_R11_21, 
      u1_R11_22, u1_R11_23, u1_R11_24, u1_R11_25, u1_R11_26, u1_R11_27, u1_R11_28, u1_R11_29, u1_R11_3, 
      u1_R11_30, u1_R11_31, u1_R11_32, u1_R11_4, u1_R11_5, u1_R11_6, u1_R11_7, u1_R11_8, u1_R11_9, 
      u1_R12_1, u1_R12_10, u1_R12_11, u1_R12_12, u1_R12_13, u1_R12_14, u1_R12_15, u1_R12_16, u1_R12_17, 
      u1_R12_18, u1_R12_19, u1_R12_2, u1_R12_20, u1_R12_21, u1_R12_22, u1_R12_23, u1_R12_24, u1_R12_25, 
      u1_R12_26, u1_R12_27, u1_R12_28, u1_R12_29, u1_R12_3, u1_R12_30, u1_R12_31, u1_R12_32, u1_R12_4, 
      u1_R12_5, u1_R12_6, u1_R12_7, u1_R12_8, u1_R12_9, u1_R13_1, u1_R13_10, u1_R13_11, u1_R13_12, 
      u1_R13_13, u1_R13_14, u1_R13_15, u1_R13_16, u1_R13_17, u1_R13_18, u1_R13_19, u1_R13_2, u1_R13_20, 
      u1_R13_21, u1_R13_22, u1_R13_23, u1_R13_24, u1_R13_25, u1_R13_26, u1_R13_27, u1_R13_28, u1_R13_29, 
      u1_R13_3, u1_R13_30, u1_R13_31, u1_R13_32, u1_R13_4, u1_R13_5, u1_R13_6, u1_R13_7, u1_R13_8, 
      u1_R13_9, u1_R1_1, u1_R1_10, u1_R1_11, u1_R1_12, u1_R1_13, u1_R1_14, u1_R1_15, u1_R1_16, 
      u1_R1_17, u1_R1_18, u1_R1_19, u1_R1_2, u1_R1_20, u1_R1_21, u1_R1_22, u1_R1_23, u1_R1_24, 
      u1_R1_25, u1_R1_26, u1_R1_27, u1_R1_28, u1_R1_29, u1_R1_3, u1_R1_30, u1_R1_31, u1_R1_32, 
      u1_R1_4, u1_R1_5, u1_R1_6, u1_R1_7, u1_R1_8, u1_R1_9, u1_R2_1, u1_R2_10, u1_R2_11, 
      u1_R2_12, u1_R2_13, u1_R2_14, u1_R2_15, u1_R2_16, u1_R2_17, u1_R2_18, u1_R2_19, u1_R2_2, 
      u1_R2_20, u1_R2_21, u1_R2_22, u1_R2_23, u1_R2_24, u1_R2_25, u1_R2_26, u1_R2_27, u1_R2_28, 
      u1_R2_29, u1_R2_3, u1_R2_30, u1_R2_31, u1_R2_32, u1_R2_4, u1_R2_5, u1_R2_6, u1_R2_7, 
      u1_R2_8, u1_R2_9, u1_R3_1, u1_R3_10, u1_R3_11, u1_R3_12, u1_R3_13, u1_R3_14, u1_R3_15, 
      u1_R3_16, u1_R3_17, u1_R3_18, u1_R3_19, u1_R3_2, u1_R3_20, u1_R3_21, u1_R3_22, u1_R3_23, 
      u1_R3_24, u1_R3_25, u1_R3_26, u1_R3_27, u1_R3_28, u1_R3_29, u1_R3_3, u1_R3_30, u1_R3_31, 
      u1_R3_32, u1_R3_4, u1_R3_5, u1_R3_6, u1_R3_7, u1_R3_8, u1_R3_9, u1_R4_1, u1_R4_10, 
      u1_R4_11, u1_R4_12, u1_R4_13, u1_R4_14, u1_R4_15, u1_R4_16, u1_R4_17, u1_R4_18, u1_R4_19, 
      u1_R4_2, u1_R4_20, u1_R4_21, u1_R4_22, u1_R4_23, u1_R4_24, u1_R4_25, u1_R4_26, u1_R4_27, 
      u1_R4_28, u1_R4_29, u1_R4_3, u1_R4_30, u1_R4_31, u1_R4_32, u1_R4_4, u1_R4_5, u1_R4_6, 
      u1_R4_7, u1_R4_8, u1_R4_9, u1_R5_1, u1_R5_10, u1_R5_11, u1_R5_12, u1_R5_13, u1_R5_14, 
      u1_R5_15, u1_R5_16, u1_R5_17, u1_R5_18, u1_R5_19, u1_R5_2, u1_R5_20, u1_R5_21, u1_R5_22, 
      u1_R5_23, u1_R5_24, u1_R5_25, u1_R5_26, u1_R5_27, u1_R5_28, u1_R5_29, u1_R5_3, u1_R5_30, 
      u1_R5_31, u1_R5_32, u1_R5_4, u1_R5_5, u1_R5_6, u1_R5_7, u1_R5_8, u1_R5_9, u1_R6_1, 
      u1_R6_10, u1_R6_11, u1_R6_12, u1_R6_13, u1_R6_14, u1_R6_15, u1_R6_16, u1_R6_17, u1_R6_18, 
      u1_R6_19, u1_R6_2, u1_R6_20, u1_R6_21, u1_R6_22, u1_R6_23, u1_R6_24, u1_R6_25, u1_R6_26, 
      u1_R6_27, u1_R6_28, u1_R6_29, u1_R6_3, u1_R6_30, u1_R6_31, u1_R6_32, u1_R6_4, u1_R6_5, 
      u1_R6_6, u1_R6_7, u1_R6_8, u1_R6_9, u1_R7_1, u1_R7_10, u1_R7_11, u1_R7_12, u1_R7_13, 
      u1_R7_14, u1_R7_15, u1_R7_16, u1_R7_17, u1_R7_18, u1_R7_19, u1_R7_2, u1_R7_20, u1_R7_21, 
      u1_R7_22, u1_R7_23, u1_R7_24, u1_R7_25, u1_R7_26, u1_R7_27, u1_R7_28, u1_R7_29, u1_R7_3, 
      u1_R7_30, u1_R7_31, u1_R7_32, u1_R7_4, u1_R7_5, u1_R7_6, u1_R7_7, u1_R7_8, u1_R7_9, 
      u1_R8_1, u1_R8_10, u1_R8_11, u1_R8_12, u1_R8_13, u1_R8_14, u1_R8_15, u1_R8_16, u1_R8_17, 
      u1_R8_18, u1_R8_19, u1_R8_2, u1_R8_20, u1_R8_21, u1_R8_22, u1_R8_23, u1_R8_24, u1_R8_25, 
      u1_R8_26, u1_R8_27, u1_R8_28, u1_R8_29, u1_R8_3, u1_R8_30, u1_R8_31, u1_R8_32, u1_R8_4, 
      u1_R8_5, u1_R8_6, u1_R8_7, u1_R8_8, u1_R8_9, u1_R9_1, u1_R9_10, u1_R9_11, u1_R9_12, 
      u1_R9_13, u1_R9_14, u1_R9_15, u1_R9_16, u1_R9_17, u1_R9_18, u1_R9_19, u1_R9_2, u1_R9_20, 
      u1_R9_21, u1_R9_22, u1_R9_23, u1_R9_24, u1_R9_25, u1_R9_26, u1_R9_27, u1_R9_28, u1_R9_29, 
      u1_R9_3, u1_R9_30, u1_R9_31, u1_R9_32, u1_R9_4, u1_R9_5, u1_R9_6, u1_R9_7, u1_R9_8, 
      u1_R9_9, u1_desIn_r_1, u1_desIn_r_11, u1_desIn_r_13, u1_desIn_r_15, u1_desIn_r_17, u1_desIn_r_19, u1_desIn_r_21, u1_desIn_r_23, 
      u1_desIn_r_25, u1_desIn_r_27, u1_desIn_r_29, u1_desIn_r_3, u1_desIn_r_31, u1_desIn_r_33, u1_desIn_r_35, u1_desIn_r_37, u1_desIn_r_39, 
      u1_desIn_r_41, u1_desIn_r_43, u1_desIn_r_45, u1_desIn_r_47, u1_desIn_r_49, u1_desIn_r_5, u1_desIn_r_51, u1_desIn_r_53, u1_desIn_r_55, 
      u1_desIn_r_57, u1_desIn_r_59, u1_desIn_r_61, u1_desIn_r_63, u1_desIn_r_7, u1_desIn_r_9, u1_key_r_0, u1_key_r_1, u1_key_r_10, 
      u1_key_r_11, u1_key_r_12, u1_key_r_13, u1_key_r_14, u1_key_r_15, u1_key_r_16, u1_key_r_17, u1_key_r_18, u1_key_r_19, 
      u1_key_r_2, u1_key_r_20, u1_key_r_21, u1_key_r_22, u1_key_r_23, u1_key_r_24, u1_key_r_25, u1_key_r_26, u1_key_r_27, 
      u1_key_r_28, u1_key_r_29, u1_key_r_3, u1_key_r_30, u1_key_r_31, u1_key_r_32, u1_key_r_33, u1_key_r_34, u1_key_r_35, 
      u1_key_r_36, u1_key_r_37, u1_key_r_38, u1_key_r_39, u1_key_r_4, u1_key_r_40, u1_key_r_41, u1_key_r_42, u1_key_r_43, 
      u1_key_r_44, u1_key_r_45, u1_key_r_46, u1_key_r_47, u1_key_r_48, u1_key_r_49, u1_key_r_5, u1_key_r_50, u1_key_r_51, 
      u1_key_r_52, u1_key_r_53, u1_key_r_54, u1_key_r_55, u1_key_r_6, u1_key_r_7, u1_key_r_8, u1_key_r_9, u1_uk_K_r0_11, 
      u1_uk_K_r0_13, u1_uk_K_r0_15, u1_uk_K_r0_17, u1_uk_K_r0_19, u1_uk_K_r0_2, u1_uk_K_r0_22, u1_uk_K_r0_25, u1_uk_K_r0_28, u1_uk_K_r0_31, 
      u1_uk_K_r0_32, u1_uk_K_r0_34, u1_uk_K_r0_36, u1_uk_K_r0_47, u1_uk_K_r0_49, u1_uk_K_r0_52, u1_uk_K_r0_55, u1_uk_K_r0_7, u1_uk_K_r10_10, 
      u1_uk_K_r10_11, u1_uk_K_r10_14, u1_uk_K_r10_16, u1_uk_K_r10_18, u1_uk_K_r10_19, u1_uk_K_r10_23, u1_uk_K_r10_25, u1_uk_K_r10_27, u1_uk_K_r10_28, 
      u1_uk_K_r10_32, u1_uk_K_r10_34, u1_uk_K_r10_37, u1_uk_K_r10_39, u1_uk_K_r10_4, u1_uk_K_r10_41, u1_uk_K_r10_42, u1_uk_K_r10_43, u1_uk_K_r10_44, 
      u1_uk_K_r10_47, u1_uk_K_r10_48, u1_uk_K_r10_49, u1_uk_K_r10_52, u1_uk_K_r10_9, u1_uk_K_r11_10, u1_uk_K_r11_11, u1_uk_K_r11_17, u1_uk_K_r11_19, 
      u1_uk_K_r11_20, u1_uk_K_r11_21, u1_uk_K_r11_24, u1_uk_K_r11_25, u1_uk_K_r11_26, u1_uk_K_r11_27, u1_uk_K_r11_28, u1_uk_K_r11_29, u1_uk_K_r11_33, 
      u1_uk_K_r11_34, u1_uk_K_r11_39, u1_uk_K_r11_4, u1_uk_K_r11_46, u1_uk_K_r11_47, u1_uk_K_r11_48, u1_uk_K_r11_5, u1_uk_K_r11_53, u1_uk_K_r11_54, 
      u1_uk_K_r11_6, u1_uk_K_r11_7, u1_uk_K_r11_8, u1_uk_K_r12_1, u1_uk_K_r12_10, u1_uk_K_r12_15, u1_uk_K_r12_16, u1_uk_K_r12_18, u1_uk_K_r12_21, 
      u1_uk_K_r12_22, u1_uk_K_r12_25, u1_uk_K_r12_30, u1_uk_K_r12_33, u1_uk_K_r12_36, u1_uk_K_r12_41, u1_uk_K_r12_42, u1_uk_K_r12_44, u1_uk_K_r12_47, 
      u1_uk_K_r12_7, u1_uk_K_r13_0, u1_uk_K_r13_13, u1_uk_K_r13_17, u1_uk_K_r13_19, u1_uk_K_r13_2, u1_uk_K_r13_22, u1_uk_K_r13_23, u1_uk_K_r13_25, 
      u1_uk_K_r13_31, u1_uk_K_r13_32, u1_uk_K_r13_35, u1_uk_K_r13_36, u1_uk_K_r13_38, u1_uk_K_r13_4, u1_uk_K_r13_44, u1_uk_K_r13_55, u1_uk_K_r14_10, 
      u1_uk_K_r14_11, u1_uk_K_r14_12, u1_uk_K_r14_15, u1_uk_K_r14_16, u1_uk_K_r14_18, u1_uk_K_r14_2, u1_uk_K_r14_23, u1_uk_K_r14_3, u1_uk_K_r14_38, 
      u1_uk_K_r14_39, u1_uk_K_r14_42, u1_uk_K_r14_43, u1_uk_K_r14_45, u1_uk_K_r14_46, u1_uk_K_r14_5, u1_uk_K_r14_50, u1_uk_K_r14_8, u1_uk_K_r14_9, 
      u1_uk_K_r1_10, u1_uk_K_r1_15, u1_uk_K_r1_16, u1_uk_K_r1_17, u1_uk_K_r1_18, u1_uk_K_r1_21, u1_uk_K_r1_22, u1_uk_K_r1_33, u1_uk_K_r1_36, 
      u1_uk_K_r1_41, u1_uk_K_r1_42, u1_uk_K_r1_44, u1_uk_K_r1_47, u1_uk_K_r1_6, u1_uk_K_r1_7, u1_uk_K_r2_13, u1_uk_K_r2_16, u1_uk_K_r2_18, 
      u1_uk_K_r2_20, u1_uk_K_r2_21, u1_uk_K_r2_24, u1_uk_K_r2_25, u1_uk_K_r2_26, u1_uk_K_r2_27, u1_uk_K_r2_28, u1_uk_K_r2_29, u1_uk_K_r2_31, 
      u1_uk_K_r2_33, u1_uk_K_r2_36, u1_uk_K_r2_4, u1_uk_K_r2_41, u1_uk_K_r2_46, u1_uk_K_r2_47, u1_uk_K_r2_49, u1_uk_K_r2_50, u1_uk_K_r2_53, 
      u1_uk_K_r2_55, u1_uk_K_r2_6, u1_uk_K_r2_7, u1_uk_K_r3_10, u1_uk_K_r3_11, u1_uk_K_r3_14, u1_uk_K_r3_15, u1_uk_K_r3_16, u1_uk_K_r3_19, 
      u1_uk_K_r3_24, u1_uk_K_r3_29, u1_uk_K_r3_33, u1_uk_K_r3_34, u1_uk_K_r3_35, u1_uk_K_r3_38, u1_uk_K_r3_4, u1_uk_K_r3_43, u1_uk_K_r3_44, 
      u1_uk_K_r3_47, u1_uk_K_r3_51, u1_uk_K_r3_52, u1_uk_K_r3_9, u1_uk_K_r4_0, u1_uk_K_r4_11, u1_uk_K_r4_17, u1_uk_K_r4_18, u1_uk_K_r4_23, 
      u1_uk_K_r4_27, u1_uk_K_r4_3, u1_uk_K_r4_31, u1_uk_K_r4_33, u1_uk_K_r4_35, u1_uk_K_r4_38, u1_uk_K_r4_4, u1_uk_K_r4_41, u1_uk_K_r4_47, 
      u1_uk_K_r4_48, u1_uk_K_r4_49, u1_uk_K_r4_5, u1_uk_K_r4_54, u1_uk_K_r4_55, u1_uk_K_r5_0, u1_uk_K_r5_1, u1_uk_K_r5_10, u1_uk_K_r5_13, 
      u1_uk_K_r5_16, u1_uk_K_r5_17, u1_uk_K_r5_18, u1_uk_K_r5_19, u1_uk_K_r5_21, u1_uk_K_r5_23, u1_uk_K_r5_26, u1_uk_K_r5_31, u1_uk_K_r5_32, 
      u1_uk_K_r5_35, u1_uk_K_r5_36, u1_uk_K_r5_37, u1_uk_K_r5_39, u1_uk_K_r5_4, u1_uk_K_r5_40, u1_uk_K_r5_41, u1_uk_K_r5_43, u1_uk_K_r5_48, 
      u1_uk_K_r5_5, u1_uk_K_r5_51, u1_uk_K_r5_53, u1_uk_K_r5_7, u1_uk_K_r5_8, u1_uk_K_r6_0, u1_uk_K_r6_10, u1_uk_K_r6_14, u1_uk_K_r6_17, 
      u1_uk_K_r6_19, u1_uk_K_r6_21, u1_uk_K_r6_22, u1_uk_K_r6_26, u1_uk_K_r6_27, u1_uk_K_r6_28, u1_uk_K_r6_29, u1_uk_K_r6_3, u1_uk_K_r6_30, 
      u1_uk_K_r6_31, u1_uk_K_r6_34, u1_uk_K_r6_35, u1_uk_K_r6_37, u1_uk_K_r6_46, u1_uk_K_r6_51, u1_uk_K_r6_53, u1_uk_K_r6_55, u1_uk_K_r6_7, 
      u1_uk_K_r7_0, u1_uk_K_r7_1, u1_uk_K_r7_13, u1_uk_K_r7_15, u1_uk_K_r7_16, u1_uk_K_r7_2, u1_uk_K_r7_20, u1_uk_K_r7_22, u1_uk_K_r7_23, 
      u1_uk_K_r7_24, u1_uk_K_r7_25, u1_uk_K_r7_26, u1_uk_K_r7_27, u1_uk_K_r7_29, u1_uk_K_r7_30, u1_uk_K_r7_31, u1_uk_K_r7_32, u1_uk_K_r7_34, 
      u1_uk_K_r7_37, u1_uk_K_r7_39, u1_uk_K_r7_41, u1_uk_K_r7_46, u1_uk_K_r7_48, u1_uk_K_r7_5, u1_uk_K_r7_53, u1_uk_K_r7_55, u1_uk_K_r7_6, 
      u1_uk_K_r7_7, u1_uk_K_r7_8, u1_uk_K_r7_9, u1_uk_K_r8_10, u1_uk_K_r8_13, u1_uk_K_r8_16, u1_uk_K_r8_17, u1_uk_K_r8_19, u1_uk_K_r8_2, 
      u1_uk_K_r8_21, u1_uk_K_r8_22, u1_uk_K_r8_27, u1_uk_K_r8_28, u1_uk_K_r8_32, u1_uk_K_r8_37, u1_uk_K_r8_39, u1_uk_K_r8_40, u1_uk_K_r8_41, 
      u1_uk_K_r8_42, u1_uk_K_r8_43, u1_uk_K_r8_44, u1_uk_K_r8_48, u1_uk_K_r8_5, u1_uk_K_r8_51, u1_uk_K_r8_52, u1_uk_K_r8_8, u1_uk_K_r9_0, 
      u1_uk_K_r9_1, u1_uk_K_r9_10, u1_uk_K_r9_12, u1_uk_K_r9_13, u1_uk_K_r9_15, u1_uk_K_r9_18, u1_uk_K_r9_19, u1_uk_K_r9_22, u1_uk_K_r9_23, 
      u1_uk_K_r9_25, u1_uk_K_r9_27, u1_uk_K_r9_30, u1_uk_K_r9_31, u1_uk_K_r9_33, u1_uk_K_r9_35, u1_uk_K_r9_38, u1_uk_K_r9_4, u1_uk_K_r9_45, 
      u1_uk_K_r9_48, u1_uk_K_r9_49, u1_uk_K_r9_5, u1_uk_K_r9_54, u1_uk_K_r9_55, u1_uk_K_r9_6, u1_uk_K_r9_7, u1_uk_K_r9_9, u1_uk_n1218, 
      u1_uk_n1219, u1_uk_n1220, u1_uk_n1221, u1_uk_n1222, u1_uk_n1224, u1_uk_n1225, u1_uk_n1227, u1_uk_n1228, u1_uk_n1229, 
      u1_uk_n1230, u1_uk_n1231, u1_uk_n1233, u1_uk_n1234, u1_uk_n1235, u1_uk_n1236, u1_uk_n1237, u1_uk_n1238, u1_uk_n1239, 
      u1_uk_n1240, u1_uk_n1241, u1_uk_n1242, u1_uk_n1243, u1_uk_n1244, u1_uk_n1245, u1_uk_n1246, u1_uk_n1247, u1_uk_n1248, 
      u1_uk_n1249, u1_uk_n1250, u1_uk_n1251, u1_uk_n1252, u1_uk_n1253, u1_uk_n1255, u1_uk_n1256, u1_uk_n1257, u1_uk_n1258, 
      u1_uk_n1259, u1_uk_n1260, u1_uk_n1261, u1_uk_n1262, u1_uk_n1263, u1_uk_n1264, u1_uk_n1265, u1_uk_n1266, u1_uk_n1267, 
      u1_uk_n1268, u1_uk_n1269, u1_uk_n1270, u1_uk_n1271, u1_uk_n1272, u1_uk_n1273, u1_uk_n1274, u1_uk_n1275, u1_uk_n1276, 
      u1_uk_n1277, u1_uk_n1278, u1_uk_n1279, u1_uk_n1281, u1_uk_n1282, u1_uk_n1284, u1_uk_n1286, u1_uk_n1288, u1_uk_n1289, 
      u1_uk_n1290, u1_uk_n1291, u1_uk_n1292, u1_uk_n1293, u1_uk_n1294, u1_uk_n1295, u1_uk_n1296, u1_uk_n1297, u1_uk_n1299, 
      u1_uk_n1300, u1_uk_n1303, u1_uk_n1304, u1_uk_n1305, u1_uk_n1307, u1_uk_n1308, u1_uk_n1309, u1_uk_n1310, u1_uk_n1311, 
      u1_uk_n1312, u1_uk_n1313, u1_uk_n1314, u1_uk_n1315, u1_uk_n1316, u1_uk_n1317, u1_uk_n1318, u1_uk_n1319, u1_uk_n1320, 
      u1_uk_n1321, u1_uk_n1322, u1_uk_n1323, u1_uk_n1324, u1_uk_n1325, u1_uk_n1326, u1_uk_n1327, u1_uk_n1328, u1_uk_n1329, 
      u1_uk_n1330, u1_uk_n1331, u1_uk_n1332, u1_uk_n1333, u1_uk_n1334, u1_uk_n1335, u1_uk_n1336, u1_uk_n1338, u1_uk_n1339, 
      u1_uk_n1340, u1_uk_n1341, u1_uk_n1342, u1_uk_n1343, u1_uk_n1344, u1_uk_n1345, u1_uk_n1346, u1_uk_n1347, u1_uk_n1348, 
      u1_uk_n1349, u1_uk_n1350, u1_uk_n1351, u1_uk_n1352, u1_uk_n1353, u1_uk_n1354, u1_uk_n1355, u1_uk_n1356, u1_uk_n1357, 
      u1_uk_n1358, u1_uk_n1359, u1_uk_n1360, u1_uk_n1361, u1_uk_n1363, u1_uk_n1365, u1_uk_n1366, u1_uk_n1367, u1_uk_n1369, 
      u1_uk_n1371, u1_uk_n1372, u1_uk_n1374, u1_uk_n1375, u1_uk_n1376, u1_uk_n1377, u1_uk_n1378, u1_uk_n1380, u1_uk_n1381, 
      u1_uk_n1382, u1_uk_n1383, u1_uk_n1386, u1_uk_n1389, u1_uk_n1390, u1_uk_n1391, u1_uk_n1393, u1_uk_n1394, u1_uk_n1395, 
      u1_uk_n1396, u1_uk_n1397, u1_uk_n1398, u1_uk_n1399, u1_uk_n1400, u1_uk_n1401, u1_uk_n1402, u1_uk_n1403, u1_uk_n1404, 
      u1_uk_n1405, u1_uk_n1406, u1_uk_n1407, u1_uk_n1408, u1_uk_n1409, u1_uk_n1410, u1_uk_n1411, u1_uk_n1412, u1_uk_n1413, 
      u1_uk_n1414, u1_uk_n1415, u1_uk_n1417, u1_uk_n1418, u1_uk_n1419, u1_uk_n1422, u1_uk_n1423, u1_uk_n1424, u1_uk_n1425, 
      u1_uk_n1426, u1_uk_n1427, u1_uk_n1429, u1_uk_n1430, u1_uk_n1431, u1_uk_n1433, u1_uk_n1435, u1_uk_n1436, u1_uk_n1437, 
      u1_uk_n1438, u1_uk_n1439, u1_uk_n1440, u1_uk_n1441, u1_uk_n1442, u1_uk_n1443, u1_uk_n1444, u1_uk_n1446, u1_uk_n1447, 
      u1_uk_n1448, u1_uk_n1449, u1_uk_n1450, u1_uk_n1452, u1_uk_n1453, u1_uk_n1454, u1_uk_n1455, u1_uk_n1456, u1_uk_n1457, 
      u1_uk_n1458, u1_uk_n1459, u1_uk_n1460, u1_uk_n1461, u1_uk_n1462, u1_uk_n1463, u1_uk_n1464, u1_uk_n1465, u1_uk_n1466, 
      u1_uk_n1468, u1_uk_n1469, u1_uk_n1470, u1_uk_n1471, u1_uk_n1472, u1_uk_n1474, u1_uk_n1475, u1_uk_n1476, u1_uk_n1477, 
      u1_uk_n1478, u1_uk_n1482, u1_uk_n1483, u1_uk_n1484, u1_uk_n1485, u1_uk_n1486, u1_uk_n1487, u1_uk_n1488, u1_uk_n1489, 
      u1_uk_n1490, u1_uk_n1491, u1_uk_n1492, u1_uk_n1494, u1_uk_n1495, u1_uk_n1496, u1_uk_n1498, u1_uk_n1499, u1_uk_n1500, 
      u1_uk_n1501, u1_uk_n1504, u1_uk_n1505, u1_uk_n1507, u1_uk_n1508, u1_uk_n1510, u1_uk_n1514, u1_uk_n1516, u1_uk_n1517, 
      u1_uk_n1518, u1_uk_n1520, u1_uk_n1521, u1_uk_n1523, u1_uk_n1524, u1_uk_n1526, u1_uk_n1527, u1_uk_n1528, u1_uk_n1529, 
      u1_uk_n1530, u1_uk_n1531, u1_uk_n1532, u1_uk_n1533, u1_uk_n1534, u1_uk_n1536, u1_uk_n1537, u1_uk_n1538, u1_uk_n1540, 
      u1_uk_n1541, u1_uk_n1543, u1_uk_n1544, u1_uk_n1545, u1_uk_n1547, u1_uk_n1548, u1_uk_n1549, u1_uk_n1551, u1_uk_n1552, 
      u1_uk_n1554, u1_uk_n1555, u1_uk_n1556, u1_uk_n1557, u1_uk_n1558, u1_uk_n1559, u1_uk_n1560, u1_uk_n1561, u1_uk_n1562, 
      u1_uk_n1563, u1_uk_n1564, u1_uk_n1565, u1_uk_n1566, u1_uk_n1567, u1_uk_n1568, u1_uk_n1570, u1_uk_n1571, u1_uk_n1572, 
      u1_uk_n1573, u1_uk_n1574, u1_uk_n1577, u1_uk_n1578, u1_uk_n1579, u1_uk_n1581, u1_uk_n1584, u1_uk_n1585, u1_uk_n1586, 
      u1_uk_n1588, u1_uk_n1592, u1_uk_n1593, u1_uk_n1595, u1_uk_n1598, u1_uk_n1599, u1_uk_n1600, u1_uk_n1601, u1_uk_n1603, 
      u1_uk_n1604, u1_uk_n1605, u1_uk_n1606, u1_uk_n1607, u1_uk_n1608, u1_uk_n1610, u1_uk_n1612, u1_uk_n1613, u1_uk_n1614, 
      u1_uk_n1615, u1_uk_n1616, u1_uk_n1618, u1_uk_n1619, u1_uk_n1620, u1_uk_n1621, u1_uk_n1622, u1_uk_n1623, u1_uk_n1624, 
      u1_uk_n1625, u1_uk_n1626, u1_uk_n1627, u1_uk_n1628, u1_uk_n1629, u1_uk_n1630, u1_uk_n1632, u1_uk_n1633, u1_uk_n1634, 
      u1_uk_n1635, u1_uk_n1639, u1_uk_n1640, u1_uk_n1641, u1_uk_n1642, u1_uk_n1643, u1_uk_n1644, u1_uk_n1645, u1_uk_n1647, 
      u1_uk_n1649, u1_uk_n1651, u1_uk_n1652, u1_uk_n1653, u1_uk_n1654, u1_uk_n1655, u1_uk_n1656, u1_uk_n1659, u1_uk_n1660, 
      u1_uk_n1661, u1_uk_n1662, u1_uk_n1663, u1_uk_n1664, u1_uk_n1667, u1_uk_n1669, u1_uk_n1670, u1_uk_n1672, u1_uk_n1673, 
      u1_uk_n1676, u1_uk_n1677, u1_uk_n1678, u1_uk_n1682, u1_uk_n1683, u1_uk_n1684, u1_uk_n1687, u1_uk_n1688, u1_uk_n1689, 
      u1_uk_n1690, u1_uk_n1691, u1_uk_n1692, u1_uk_n1693, u1_uk_n1694, u1_uk_n1695, u1_uk_n1696, u1_uk_n1698, u1_uk_n1699, 
      u1_uk_n1702, u1_uk_n1703, u1_uk_n1704, u1_uk_n1705, u1_uk_n1707, u1_uk_n1708, u1_uk_n1709, u1_uk_n1710, u1_uk_n1711, 
      u1_uk_n1712, u1_uk_n1713, u1_uk_n1714, u1_uk_n1715, u1_uk_n1716, u1_uk_n1717, u1_uk_n1718, u1_uk_n1719, u1_uk_n1720, 
      u1_uk_n1721, u1_uk_n1722, u1_uk_n1723, u1_uk_n1728, u1_uk_n1729, u1_uk_n1730, u1_uk_n1731, u1_uk_n1732, u1_uk_n1734, 
      u1_uk_n1735, u1_uk_n1736, u1_uk_n1737, u1_uk_n1738, u1_uk_n1739, u1_uk_n1744, u1_uk_n1745, u1_uk_n1748, u1_uk_n1749, 
      u1_uk_n1750, u1_uk_n1751, u1_uk_n1752, u1_uk_n1753, u1_uk_n1754, u1_uk_n1755, u1_uk_n1756, u1_uk_n1757, u1_uk_n1758, 
      u1_uk_n1761, u1_uk_n1762, u1_uk_n1763, u1_uk_n1764, u1_uk_n1765, u1_uk_n1766, u1_uk_n1767, u1_uk_n1768, u1_uk_n1769, 
      u1_uk_n1772, u1_uk_n1773, u1_uk_n1774, u1_uk_n1775, u1_uk_n1776, u1_uk_n1777, u1_uk_n1780, u1_uk_n1781, u1_uk_n1782, 
      u1_uk_n1783, u1_uk_n1784, u1_uk_n1785, u1_uk_n1787, u1_uk_n1790, u1_uk_n1791, u1_uk_n1792, u1_uk_n1793, u1_uk_n1797, 
      u1_uk_n1798, u1_uk_n1799, u1_uk_n1800, u1_uk_n1801, u1_uk_n1802, u1_uk_n1803, u1_uk_n1804, u1_uk_n1806, u1_uk_n1807, 
      u1_uk_n1808, u1_uk_n1809, u1_uk_n1810, u1_uk_n1811, u1_uk_n1812, u1_uk_n1813, u1_uk_n1814, u1_uk_n1815, u1_uk_n1816, 
      u1_uk_n1817, u1_uk_n1818, u1_uk_n1819, u1_uk_n1820, u1_uk_n1821, u1_uk_n1822, u1_uk_n1823, u1_uk_n1824, u1_uk_n1826, 
      u1_uk_n1827, u1_uk_n1829, u1_uk_n1830, u1_uk_n1831, u1_uk_n1832, u1_uk_n1833, u1_uk_n1834, u1_uk_n1835, u1_uk_n1836, 
      u1_uk_n1837, u1_uk_n1838, u1_uk_n1839, u1_uk_n1840, u1_uk_n1841, u1_uk_n1842, u1_uk_n1843, u1_uk_n1844, u1_uk_n1845, 
      u1_uk_n1846, u1_uk_n1847, u1_uk_n1848, u1_uk_n1849, u1_uk_n1850, u1_uk_n1851, u1_uk_n1852, u1_uk_n1853, u1_uk_n1854, 
      u1_uk_n1855, u1_uk_n1856, u1_uk_n1858, u1_uk_n1859, u1_uk_n1860, u1_uk_n1862, u1_uk_n1863, u1_uk_n1864, u1_uk_n1865, 
      u1_uk_n1866, u1_uk_n1867, u1_uk_n1868, u1_uk_n1869, u1_uk_n1870, u1_uk_n1872, u1_uk_n1873, u1_uk_n1874, u1_uk_n1875, 
      u1_uk_n1876, u1_uk_n1879, u1_uk_n1880, u1_uk_n1881, u1_uk_n1882, u1_uk_n1883, u1_uk_n1884, u1_uk_n1885, u1_uk_n1886, 
      u1_uk_n1887, u2_FP_33, u2_FP_34, u2_FP_35, u2_FP_36, u2_FP_37, u2_FP_40, u2_FP_41, u2_FP_42, 
      u2_FP_44, u2_FP_46, u2_FP_47, u2_FP_48, u2_FP_49, u2_FP_51, u2_FP_52, u2_FP_53, u2_FP_54, 
      u2_FP_55, u2_FP_56, u2_FP_57, u2_FP_58, u2_FP_59, u2_FP_60, u2_FP_61, u2_FP_62, u2_FP_63, 
      u2_FP_64, u2_K10_11, u2_K10_17, u2_K10_19, u2_K10_25, u2_K10_26, u2_K10_29, u2_K10_36, u2_K10_42, 
      u2_K10_43, u2_K10_44, u2_K10_5, u2_K10_6, u2_K11_11, u2_K11_13, u2_K11_18, u2_K11_29, u2_K11_37, 
      u2_K11_38, u2_K11_42, u2_K11_45, u2_K11_48, u2_K11_6, u2_K11_7, u2_K12_2, u2_K12_20, u2_K12_22, 
      u2_K12_24, u2_K12_25, u2_K12_26, u2_K12_41, u2_K12_46, u2_K12_47, u2_K12_48, u2_K12_8, u2_K13_14, 
      u2_K13_20, u2_K13_25, u2_K13_26, u2_K13_3, u2_K13_31, u2_K13_32, u2_K13_34, u2_K13_37, u2_K13_40, 
      u2_K13_42, u2_K13_44, u2_K13_45, u2_K13_46, u2_K13_47, u2_K13_8, u2_K14_10, u2_K14_11, u2_K14_12, 
      u2_K14_13, u2_K14_14, u2_K14_16, u2_K14_17, u2_K14_18, u2_K14_3, u2_K14_42, u2_K14_43, u2_K14_48, 
      u2_K14_6, u2_K14_8, u2_K15_1, u2_K15_13, u2_K15_16, u2_K15_18, u2_K15_2, u2_K15_20, u2_K15_29, 
      u2_K15_31, u2_K15_35, u2_K15_37, u2_K15_44, u2_K15_47, u2_K15_48, u2_K15_5, u2_K16_26, u2_K16_31, 
      u2_K16_42, u2_K16_44, u2_K16_47, u2_K16_5, u2_K16_6, u2_K16_8, u2_K1_19, u2_K1_24, u2_K1_30, 
      u2_K1_37, u2_K1_43, u2_K2_1, u2_K2_12, u2_K2_18, u2_K2_20, u2_K2_29, u2_K2_36, u2_K2_43, 
      u2_K2_47, u2_K2_48, u2_K3_13, u2_K3_19, u2_K3_23, u2_K3_26, u2_K3_35, u2_K3_48, u2_K4_13, 
      u2_K4_14, u2_K4_18, u2_K4_19, u2_K4_35, u2_K5_11, u2_K5_13, u2_K5_14, u2_K5_17, u2_K5_18, 
      u2_K5_19, u2_K5_2, u2_K5_29, u2_K5_30, u2_K5_31, u2_K5_32, u2_K5_41, u2_K5_44, u2_K5_48, 
      u2_K5_5, u2_K5_6, u2_K5_8, u2_K6_11, u2_K6_13, u2_K6_19, u2_K6_20, u2_K6_23, u2_K6_24, 
      u2_K6_25, u2_K6_36, u2_K6_48, u2_K6_5, u2_K6_6, u2_K6_8, u2_K7_26, u2_K7_35, u2_K7_37, 
      u2_K7_38, u2_K7_43, u2_K7_44, u2_K7_48, u2_K7_5, u2_K7_7, u2_K8_13, u2_K8_18, u2_K8_24, 
      u2_K8_26, u2_K8_31, u2_K8_41, u2_K8_42, u2_K8_45, u2_K8_5, u2_K8_8, u2_K9_12, u2_K9_14, 
      u2_K9_23, u2_K9_25, u2_K9_29, u2_K9_3, u2_K9_32, u2_K9_36, u2_K9_38, u2_K9_40, u2_K9_45, 
      u2_K9_5, u2_L10_1, u2_L10_10, u2_L10_15, u2_L10_16, u2_L10_17, u2_L10_20, u2_L10_21, u2_L10_23, 
      u2_L10_24, u2_L10_26, u2_L10_27, u2_L10_30, u2_L10_31, u2_L10_5, u2_L10_6, u2_L10_9, u2_L11_1, 
      u2_L11_10, u2_L11_11, u2_L11_12, u2_L11_13, u2_L11_14, u2_L11_15, u2_L11_16, u2_L11_17, u2_L11_18, 
      u2_L11_19, u2_L11_2, u2_L11_20, u2_L11_21, u2_L11_22, u2_L11_23, u2_L11_24, u2_L11_25, u2_L11_26, 
      u2_L11_3, u2_L11_30, u2_L11_31, u2_L11_32, u2_L11_4, u2_L11_5, u2_L11_6, u2_L11_7, u2_L11_8, 
      u2_L11_9, u2_L12_13, u2_L12_15, u2_L12_16, u2_L12_17, u2_L12_18, u2_L12_2, u2_L12_21, u2_L12_23, 
      u2_L12_24, u2_L12_27, u2_L12_28, u2_L12_30, u2_L12_31, u2_L12_5, u2_L12_6, u2_L12_9, u2_L13_13, 
      u2_L13_16, u2_L13_18, u2_L13_2, u2_L13_24, u2_L13_28, u2_L13_30, u2_L13_6, u2_L14_11, u2_L14_12, 
      u2_L14_15, u2_L14_19, u2_L14_21, u2_L14_22, u2_L14_27, u2_L14_29, u2_L14_32, u2_L14_4, u2_L14_5, 
      u2_L14_7, u2_L6_11, u2_L6_14, u2_L6_15, u2_L6_19, u2_L6_21, u2_L6_22, u2_L6_25, u2_L6_27, 
      u2_L6_29, u2_L6_3, u2_L6_32, u2_L6_4, u2_L6_5, u2_L6_7, u2_L6_8, u2_L7_11, u2_L7_12, 
      u2_L7_15, u2_L7_17, u2_L7_19, u2_L7_21, u2_L7_22, u2_L7_23, u2_L7_27, u2_L7_29, u2_L7_31, 
      u2_L7_32, u2_L7_4, u2_L7_5, u2_L7_7, u2_L7_9, u2_L9_12, u2_L9_14, u2_L9_15, u2_L9_21, 
      u2_L9_22, u2_L9_25, u2_L9_27, u2_L9_3, u2_L9_32, u2_L9_5, u2_L9_7, u2_L9_8, u2_R0_1, 
      u2_R0_10, u2_R0_12, u2_R0_13, u2_R0_14, u2_R0_15, u2_R0_17, u2_R0_18, u2_R0_19, u2_R0_20, 
      u2_R0_21, u2_R0_25, u2_R0_28, u2_R0_3, u2_R0_32, u2_R0_4, u2_R0_5, u2_R0_6, u2_R0_7, 
      u2_R0_8, u2_R0_9, u2_R10_1, u2_R10_10, u2_R10_11, u2_R10_12, u2_R10_13, u2_R10_14, u2_R10_15, 
      u2_R10_16, u2_R10_17, u2_R10_19, u2_R10_2, u2_R10_21, u2_R10_28, u2_R10_29, u2_R10_3, u2_R10_30, 
      u2_R10_31, u2_R10_32, u2_R10_4, u2_R10_5, u2_R10_7, u2_R10_8, u2_R10_9, u2_R11_1, u2_R11_10, 
      u2_R11_11, u2_R11_12, u2_R11_13, u2_R11_14, u2_R11_15, u2_R11_16, u2_R11_17, u2_R11_18, u2_R11_19, 
      u2_R11_2, u2_R11_20, u2_R11_21, u2_R11_22, u2_R11_23, u2_R11_24, u2_R11_25, u2_R11_26, u2_R11_27, 
      u2_R11_28, u2_R11_29, u2_R11_3, u2_R11_30, u2_R11_31, u2_R11_32, u2_R11_4, u2_R11_5, u2_R11_6, 
      u2_R11_7, u2_R11_8, u2_R11_9, u2_R12_1, u2_R12_10, u2_R12_11, u2_R12_12, u2_R12_13, u2_R12_17, 
      u2_R12_18, u2_R12_2, u2_R12_20, u2_R12_21, u2_R12_22, u2_R12_23, u2_R12_24, u2_R12_25, u2_R12_27, 
      u2_R12_28, u2_R12_29, u2_R12_3, u2_R12_30, u2_R12_31, u2_R12_32, u2_R12_4, u2_R12_5, u2_R12_6, 
      u2_R12_7, u2_R12_8, u2_R12_9, u2_R13_1, u2_R13_10, u2_R13_11, u2_R13_12, u2_R13_13, u2_R13_17, 
      u2_R13_18, u2_R13_20, u2_R13_22, u2_R13_24, u2_R13_25, u2_R13_27, u2_R13_28, u2_R13_29, u2_R13_30, 
      u2_R13_32, u2_R13_4, u2_R13_5, u2_R13_6, u2_R13_7, u2_R13_8, u2_R13_9, u2_R1_1, u2_R1_12, 
      u2_R1_16, u2_R1_17, u2_R1_19, u2_R1_20, u2_R1_22, u2_R1_24, u2_R1_25, u2_R1_27, u2_R1_3, 
      u2_R1_30, u2_R1_5, u2_R1_8, u2_R1_9, u2_R2_1, u2_R2_11, u2_R2_12, u2_R2_13, u2_R2_16, 
      u2_R2_17, u2_R2_2, u2_R2_20, u2_R2_21, u2_R2_24, u2_R2_28, u2_R2_3, u2_R2_32, u2_R2_6, 
      u2_R2_7, u2_R2_8, u2_R2_9, u2_R3_1, u2_R3_12, u2_R3_13, u2_R3_15, u2_R3_18, u2_R3_20, 
      u2_R3_21, u2_R3_24, u2_R3_28, u2_R3_29, u2_R3_3, u2_R3_30, u2_R3_4, u2_R3_5, u2_R3_8, 
      u2_R3_9, u2_R4_1, u2_R4_12, u2_R4_13, u2_R4_14, u2_R4_16, u2_R4_17, u2_R4_19, u2_R4_20, 
      u2_R4_24, u2_R4_25, u2_R4_26, u2_R4_28, u2_R4_29, u2_R4_4, u2_R4_5, u2_R4_6, u2_R4_7, 
      u2_R4_8, u2_R5_1, u2_R5_10, u2_R5_11, u2_R5_12, u2_R5_13, u2_R5_14, u2_R5_16, u2_R5_17, 
      u2_R5_18, u2_R5_21, u2_R5_23, u2_R5_24, u2_R5_25, u2_R5_26, u2_R5_28, u2_R5_29, u2_R5_32, 
      u2_R5_4, u2_R5_5, u2_R5_8, u2_R5_9, u2_R6_1, u2_R6_10, u2_R6_11, u2_R6_12, u2_R6_13, 
      u2_R6_15, u2_R6_16, u2_R6_17, u2_R6_18, u2_R6_19, u2_R6_2, u2_R6_20, u2_R6_21, u2_R6_22, 
      u2_R6_23, u2_R6_24, u2_R6_25, u2_R6_26, u2_R6_27, u2_R6_28, u2_R6_29, u2_R6_30, u2_R6_31, 
      u2_R6_32, u2_R6_4, u2_R6_5, u2_R6_6, u2_R6_7, u2_R6_8, u2_R6_9, u2_R7_1, u2_R7_11, 
      u2_R7_12, u2_R7_13, u2_R7_14, u2_R7_15, u2_R7_16, u2_R7_17, u2_R7_2, u2_R7_20, u2_R7_21, 
      u2_R7_22, u2_R7_23, u2_R7_24, u2_R7_25, u2_R7_26, u2_R7_27, u2_R7_28, u2_R7_29, u2_R7_3, 
      u2_R7_30, u2_R7_31, u2_R7_32, u2_R7_4, u2_R7_5, u2_R7_6, u2_R7_7, u2_R7_8, u2_R7_9, 
      u2_R8_1, u2_R8_12, u2_R8_13, u2_R8_15, u2_R8_16, u2_R8_17, u2_R8_18, u2_R8_19, u2_R8_20, 
      u2_R8_22, u2_R8_24, u2_R8_25, u2_R8_26, u2_R8_27, u2_R8_28, u2_R8_29, u2_R8_32, u2_R8_4, 
      u2_R8_5, u2_R8_6, u2_R8_8, u2_R8_9, u2_R9_1, u2_R9_12, u2_R9_13, u2_R9_15, u2_R9_16, 
      u2_R9_17, u2_R9_18, u2_R9_19, u2_R9_2, u2_R9_20, u2_R9_21, u2_R9_24, u2_R9_25, u2_R9_26, 
      u2_R9_27, u2_R9_28, u2_R9_29, u2_R9_30, u2_R9_31, u2_R9_32, u2_R9_4, u2_R9_5, u2_R9_8, 
      u2_R9_9, u2_desIn_r_1, u2_desIn_r_11, u2_desIn_r_15, u2_desIn_r_23, u2_desIn_r_25, u2_desIn_r_27, u2_desIn_r_29, u2_desIn_r_3, 
      u2_desIn_r_33, u2_desIn_r_35, u2_desIn_r_37, u2_desIn_r_39, u2_desIn_r_43, u2_desIn_r_45, u2_desIn_r_5, u2_desIn_r_53, u2_desIn_r_55, 
      u2_desIn_r_57, u2_desIn_r_59, u2_desIn_r_61, u2_desIn_r_63, u2_desIn_r_7, u2_desIn_r_9, u2_key_r_0, u2_key_r_10, u2_key_r_11, 
      u2_key_r_12, u2_key_r_14, u2_key_r_16, u2_key_r_17, u2_key_r_19, u2_key_r_21, u2_key_r_22, u2_key_r_23, u2_key_r_24, 
      u2_key_r_25, u2_key_r_26, u2_key_r_28, u2_key_r_29, u2_key_r_3, u2_key_r_30, u2_key_r_31, u2_key_r_32, u2_key_r_33, 
      u2_key_r_34, u2_key_r_35, u2_key_r_36, u2_key_r_37, u2_key_r_40, u2_key_r_41, u2_key_r_42, u2_key_r_43, u2_key_r_44, 
      u2_key_r_46, u2_key_r_47, u2_key_r_48, u2_key_r_51, u2_key_r_53, u2_key_r_55, u2_key_r_6, u2_key_r_7, u2_u0_X_15, 
      u2_u0_X_16, u2_u0_X_28, u2_u0_X_34, u2_u0_X_40, u2_u0_X_45, u2_u0_X_46, u2_u0_X_5, u2_u0_X_7, u2_u0_X_9, 
      u2_u10_X_10, u2_u10_X_15, u2_u10_X_16, u2_u10_X_21, u2_u10_X_33, u2_u10_X_34, u2_u10_X_4, u2_u10_X_9, u2_u11_X_27, 
      u2_u11_X_29, u2_u11_X_31, u2_u11_X_33, u2_u11_X_34, u2_u11_X_35, u2_u11_X_36, u2_u11_X_37, u2_u11_X_38, u2_u11_X_39, 
      u2_u11_X_40, u2_u11_X_9, u2_u13_X_21, u2_u13_X_22, u2_u13_X_23, u2_u13_X_25, u2_u13_X_28, u2_u13_X_39, u2_u14_X_21, 
      u2_u14_X_22, u2_u14_X_23, u2_u14_X_25, u2_u14_X_28, u2_u14_X_3, u2_u14_X_30, u2_u14_X_32, u2_u14_X_34, u2_u14_X_39, 
      u2_u14_X_4, u2_u14_X_46, u2_u15_X_10, u2_u15_X_16, u2_u15_X_18, u2_u15_X_20, u2_u15_X_27, u2_u15_X_9, u2_u1_X_16, 
      u2_u1_X_23, u2_u1_X_25, u2_u1_X_3, u2_u1_X_33, u2_u1_X_34, u2_u1_X_35, u2_u1_X_37, u2_u1_X_39, u2_u1_X_40, 
      u2_u1_X_42, u2_u1_X_44, u2_u1_X_45, u2_u1_X_46, u2_u2_X_1, u2_u2_X_10, u2_u2_X_15, u2_u2_X_16, u2_u2_X_18, 
      u2_u2_X_20, u2_u2_X_21, u2_u2_X_22, u2_u2_X_27, u2_u2_X_3, u2_u2_X_30, u2_u2_X_32, u2_u2_X_34, u2_u2_X_39, 
      u2_u2_X_41, u2_u2_X_42, u2_u2_X_43, u2_u2_X_44, u2_u2_X_46, u2_u2_X_47, u2_u2_X_5, u2_u2_X_7, u2_u2_X_9, 
      u2_u3_X_15, u2_u3_X_21, u2_u3_X_22, u2_u3_X_27, u2_u3_X_28, u2_u3_X_33, u2_u3_X_34, u2_u3_X_36, u2_u3_X_38, 
      u2_u3_X_39, u2_u3_X_40, u2_u3_X_42, u2_u3_X_44, u2_u3_X_45, u2_u3_X_46, u2_u3_X_5, u2_u3_X_6, u2_u3_X_7, 
      u2_u3_X_8, u2_u4_X_1, u2_u4_X_10, u2_u4_X_15, u2_u4_X_16, u2_u4_X_21, u2_u4_X_23, u2_u4_X_24, u2_u4_X_25, 
      u2_u4_X_26, u2_u4_X_28, u2_u4_X_3, u2_u4_X_33, u2_u4_X_34, u2_u4_X_36, u2_u4_X_38, u2_u4_X_39, u2_u4_X_40, 
      u2_u4_X_46, u2_u4_X_47, u2_u4_X_9, u2_u5_X_1, u2_u5_X_12, u2_u5_X_14, u2_u5_X_15, u2_u5_X_16, u2_u5_X_22, 
      u2_u5_X_27, u2_u5_X_3, u2_u5_X_30, u2_u5_X_32, u2_u5_X_33, u2_u5_X_34, u2_u5_X_4, u2_u5_X_40, u2_u5_X_45, 
      u2_u5_X_46, u2_u5_X_47, u2_u6_X_10, u2_u6_X_22, u2_u6_X_28, u2_u6_X_29, u2_u6_X_3, u2_u6_X_31, u2_u6_X_33, 
      u2_u6_X_4, u2_u6_X_40, u2_u6_X_45, u2_u6_X_46, u2_u6_X_9, u2_u7_X_21, u2_u7_X_4, u2_u8_X_15, u2_u8_X_27, 
      u2_u8_X_28, u2_u9_X_10, u2_u9_X_15, u2_u9_X_16, u2_u9_X_21, u2_u9_X_3, u2_u9_X_30, u2_u9_X_32, u2_u9_X_34, 
      u2_u9_X_4, u2_u9_X_45, u2_u9_X_46, u2_uk_K_r0_11, u2_uk_K_r0_15, u2_uk_K_r0_17, u2_uk_K_r0_25, u2_uk_K_r0_32, u2_uk_K_r0_36, 
      u2_uk_K_r0_47, u2_uk_K_r0_49, u2_uk_K_r10_10, u2_uk_K_r10_25, u2_uk_K_r10_27, u2_uk_K_r10_32, u2_uk_K_r10_34, u2_uk_K_r10_4, u2_uk_K_r10_41, 
      u2_uk_K_r10_43, u2_uk_K_r11_10, u2_uk_K_r11_11, u2_uk_K_r11_19, u2_uk_K_r11_20, u2_uk_K_r11_21, u2_uk_K_r11_24, u2_uk_K_r11_25, u2_uk_K_r11_26, 
      u2_uk_K_r11_27, u2_uk_K_r11_28, u2_uk_K_r11_29, u2_uk_K_r11_39, u2_uk_K_r11_47, u2_uk_K_r11_48, u2_uk_K_r11_53, u2_uk_K_r11_6, u2_uk_K_r12_10, 
      u2_uk_K_r12_15, u2_uk_K_r12_16, u2_uk_K_r12_25, u2_uk_K_r12_33, u2_uk_K_r12_41, u2_uk_K_r12_42, u2_uk_K_r13_19, u2_uk_K_r13_25, u2_uk_K_r13_32, 
      u2_uk_K_r13_55, u2_uk_K_r14_10, u2_uk_K_r14_12, u2_uk_K_r14_15, u2_uk_K_r14_16, u2_uk_K_r14_18, u2_uk_K_r14_2, u2_uk_K_r14_3, u2_uk_K_r14_45, 
      u2_uk_K_r14_46, u2_uk_K_r14_50, u2_uk_K_r14_9, u2_uk_K_r1_16, u2_uk_K_r1_21, u2_uk_K_r1_44, u2_uk_K_r2_13, u2_uk_K_r2_18, u2_uk_K_r2_25, 
      u2_uk_K_r2_27, u2_uk_K_r2_28, u2_uk_K_r2_31, u2_uk_K_r2_36, u2_uk_K_r2_49, u2_uk_K_r2_55, u2_uk_K_r3_11, u2_uk_K_r3_19, u2_uk_K_r3_4, 
      u2_uk_K_r3_43, u2_uk_K_r3_9, u2_uk_K_r4_0, u2_uk_K_r4_11, u2_uk_K_r4_17, u2_uk_K_r4_33, u2_uk_K_r4_35, u2_uk_K_r4_38, u2_uk_K_r4_4, 
      u2_uk_K_r4_5, u2_uk_K_r4_55, u2_uk_K_r5_10, u2_uk_K_r5_19, u2_uk_K_r5_41, u2_uk_K_r6_0, u2_uk_K_r6_10, u2_uk_K_r6_14, u2_uk_K_r6_26, 
      u2_uk_K_r6_29, u2_uk_K_r6_3, u2_uk_K_r6_31, u2_uk_K_r6_34, u2_uk_K_r6_37, u2_uk_K_r6_51, u2_uk_K_r6_53, u2_uk_K_r6_7, u2_uk_K_r7_0, 
      u2_uk_K_r7_25, u2_uk_K_r7_26, u2_uk_K_r7_31, u2_uk_K_r7_32, u2_uk_K_r7_37, u2_uk_K_r7_39, u2_uk_K_r7_46, u2_uk_K_r8_13, u2_uk_K_r8_16, 
      u2_uk_K_r8_2, u2_uk_K_r8_22, u2_uk_K_r8_37, u2_uk_K_r8_40, u2_uk_K_r8_41, u2_uk_K_r8_42, u2_uk_K_r8_43, u2_uk_K_r8_48, u2_uk_K_r9_10, 
      u2_uk_K_r9_13, u2_uk_K_r9_15, u2_uk_K_r9_19, u2_uk_K_r9_23, u2_uk_K_r9_25, u2_uk_K_r9_27, u2_uk_K_r9_31, u2_uk_K_r9_4, u2_uk_K_r9_48, 
      u2_uk_K_r9_55, u2_uk_n1001, u2_uk_n1004, u2_uk_n1008, u2_uk_n1020, u2_uk_n1024, u2_uk_n1027, u2_uk_n1028, u2_uk_n1031, 
      u2_uk_n1035, u2_uk_n1036, u2_uk_n1043, u2_uk_n1044, u2_uk_n1046, u2_uk_n1049, u2_uk_n1053, u2_uk_n1058, u2_uk_n1069, 
      u2_uk_n1074, u2_uk_n1075, u2_uk_n1076, u2_uk_n1077, u2_uk_n1079, u2_uk_n1082, u2_uk_n1083, u2_uk_n1084, u2_uk_n1085, 
      u2_uk_n1088, u2_uk_n1089, u2_uk_n1091, u2_uk_n1093, u2_uk_n1095, u2_uk_n1096, u2_uk_n1097, u2_uk_n1100, u2_uk_n1104, 
      u2_uk_n1105, u2_uk_n1107, u2_uk_n1113, u2_uk_n1118, u2_uk_n1120, u2_uk_n1124, u2_uk_n1125, u2_uk_n1127, u2_uk_n1128, 
      u2_uk_n1130, u2_uk_n1131, u2_uk_n1132, u2_uk_n1133, u2_uk_n1134, u2_uk_n1136, u2_uk_n1137, u2_uk_n1140, u2_uk_n1141, 
      u2_uk_n1145, u2_uk_n1188, u2_uk_n1189, u2_uk_n1190, u2_uk_n1194, u2_uk_n1197, u2_uk_n1198, u2_uk_n1199, u2_uk_n1200, 
      u2_uk_n1201, u2_uk_n1203, u2_uk_n1204, u2_uk_n1205, u2_uk_n1206, u2_uk_n1207, u2_uk_n1208, u2_uk_n1209, u2_uk_n1210, 
      u2_uk_n1212, u2_uk_n1213, u2_uk_n1215, u2_uk_n1216, u2_uk_n1217, u2_uk_n1218, u2_uk_n1220, u2_uk_n1221, u2_uk_n1223, 
      u2_uk_n1225, u2_uk_n1226, u2_uk_n1227, u2_uk_n1228, u2_uk_n1230, u2_uk_n1231, u2_uk_n1232, u2_uk_n1234, u2_uk_n1238, 
      u2_uk_n1240, u2_uk_n1243, u2_uk_n1244, u2_uk_n1245, u2_uk_n1246, u2_uk_n1247, u2_uk_n1249, u2_uk_n1259, u2_uk_n1260, 
      u2_uk_n1261, u2_uk_n1265, u2_uk_n1267, u2_uk_n1270, u2_uk_n1275, u2_uk_n1279, u2_uk_n1280, u2_uk_n1282, u2_uk_n1283, 
      u2_uk_n1284, u2_uk_n1285, u2_uk_n1287, u2_uk_n1292, u2_uk_n1293, u2_uk_n1296, u2_uk_n1298, u2_uk_n1300, u2_uk_n1301, 
      u2_uk_n1303, u2_uk_n1305, u2_uk_n1306, u2_uk_n1309, u2_uk_n1310, u2_uk_n1311, u2_uk_n1313, u2_uk_n1314, u2_uk_n1317, 
      u2_uk_n1319, u2_uk_n1322, u2_uk_n1323, u2_uk_n1325, u2_uk_n1326, u2_uk_n1329, u2_uk_n1331, u2_uk_n1333, u2_uk_n1336, 
      u2_uk_n1339, u2_uk_n1341, u2_uk_n1345, u2_uk_n1350, u2_uk_n1353, u2_uk_n1359, u2_uk_n1361, u2_uk_n1363, u2_uk_n1365, 
      u2_uk_n1370, u2_uk_n1375, u2_uk_n1381, u2_uk_n1382, u2_uk_n1403, u2_uk_n1405, u2_uk_n1408, u2_uk_n1411, u2_uk_n1412, 
      u2_uk_n1418, u2_uk_n1420, u2_uk_n1425, u2_uk_n1428, u2_uk_n1430, u2_uk_n1435, u2_uk_n1438, u2_uk_n1439, u2_uk_n1445, 
      u2_uk_n1446, u2_uk_n1447, u2_uk_n1453, u2_uk_n1454, u2_uk_n1456, u2_uk_n1458, u2_uk_n1460, u2_uk_n1462, u2_uk_n1465, 
      u2_uk_n1466, u2_uk_n1470, u2_uk_n1475, u2_uk_n1486, u2_uk_n1488, u2_uk_n1491, u2_uk_n1493, u2_uk_n1494, u2_uk_n1496, 
      u2_uk_n1497, u2_uk_n1498, u2_uk_n1499, u2_uk_n1500, u2_uk_n1502, u2_uk_n1503, u2_uk_n1504, u2_uk_n1506, u2_uk_n1508, 
      u2_uk_n1511, u2_uk_n1513, u2_uk_n1514, u2_uk_n1515, u2_uk_n1517, u2_uk_n1518, u2_uk_n1519, u2_uk_n1521, u2_uk_n1522, 
      u2_uk_n1524, u2_uk_n1525, u2_uk_n1526, u2_uk_n1527, u2_uk_n1529, u2_uk_n1530, u2_uk_n1531, u2_uk_n1532, u2_uk_n1533, 
      u2_uk_n1535, u2_uk_n1536, u2_uk_n1537, u2_uk_n1538, u2_uk_n1542, u2_uk_n1544, u2_uk_n1548, u2_uk_n1549, u2_uk_n1551, 
      u2_uk_n1555, u2_uk_n1556, u2_uk_n1558, u2_uk_n1563, u2_uk_n1565, u2_uk_n1568, u2_uk_n1570, u2_uk_n1571, u2_uk_n1573, 
      u2_uk_n1576, u2_uk_n1577, u2_uk_n1580, u2_uk_n1583, u2_uk_n1585, u2_uk_n1586, u2_uk_n1590, u2_uk_n1591, u2_uk_n1592, 
      u2_uk_n1594, u2_uk_n1599, u2_uk_n1600, u2_uk_n1602, u2_uk_n1604, u2_uk_n1605, u2_uk_n1609, u2_uk_n1610, u2_uk_n1615, 
      u2_uk_n1617, u2_uk_n1622, u2_uk_n1624, u2_uk_n1626, u2_uk_n1629, u2_uk_n1631, u2_uk_n1632, u2_uk_n1634, u2_uk_n1639, 
      u2_uk_n1640, u2_uk_n1642, u2_uk_n1643, u2_uk_n1647, u2_uk_n1652, u2_uk_n1653, u2_uk_n1654, u2_uk_n1657, u2_uk_n1658, 
      u2_uk_n1660, u2_uk_n1665, u2_uk_n1666, u2_uk_n1668, u2_uk_n1672, u2_uk_n1673, u2_uk_n1674, u2_uk_n1675, u2_uk_n1677, 
      u2_uk_n1680, u2_uk_n1681, u2_uk_n1682, u2_uk_n1683, u2_uk_n1684, u2_uk_n1687, u2_uk_n1688, u2_uk_n1689, u2_uk_n1693, 
      u2_uk_n1702, u2_uk_n1707, u2_uk_n1708, u2_uk_n1709, u2_uk_n1720, u2_uk_n1721, u2_uk_n1723, u2_uk_n1724, u2_uk_n1725, 
      u2_uk_n1726, u2_uk_n1727, u2_uk_n1728, u2_uk_n1731, u2_uk_n1732, u2_uk_n1734, u2_uk_n1736, u2_uk_n1737, u2_uk_n1738, 
      u2_uk_n1742, u2_uk_n1743, u2_uk_n1744, u2_uk_n1745, u2_uk_n1746, u2_uk_n1747, u2_uk_n1750, u2_uk_n1753, u2_uk_n1755, 
      u2_uk_n1761, u2_uk_n1762, u2_uk_n1763, u2_uk_n1767, u2_uk_n1769, u2_uk_n1770, u2_uk_n1773, u2_uk_n1776, u2_uk_n1777, 
      u2_uk_n1778, u2_uk_n1781, u2_uk_n1782, u2_uk_n1783, u2_uk_n1785, u2_uk_n1786, u2_uk_n1788, u2_uk_n1789, u2_uk_n1790, 
      u2_uk_n1791, u2_uk_n1792, u2_uk_n1793, u2_uk_n1794, u2_uk_n1796, u2_uk_n1797, u2_uk_n1800, u2_uk_n1801, u2_uk_n1803, 
      u2_uk_n1805, u2_uk_n1807, u2_uk_n1808, u2_uk_n1809, u2_uk_n1811, u2_uk_n1814, u2_uk_n1815, u2_uk_n1816, u2_uk_n1817, 
      u2_uk_n1821, u2_uk_n1823, u2_uk_n1826, u2_uk_n1832, u2_uk_n1833, u2_uk_n1834, u2_uk_n1835, u2_uk_n1837, u2_uk_n1839, 
      u2_uk_n1840, u2_uk_n1843, u2_uk_n1849, u2_uk_n1850, u2_uk_n1851, u2_uk_n1852, u2_uk_n1853, u2_uk_n1855, u2_uk_n238, 
      u2_uk_n240, u2_uk_n251, u2_uk_n257, u2_uk_n299, u2_uk_n301, u2_uk_n305, u2_uk_n308, u2_uk_n313, u2_uk_n319, 
      u2_uk_n363, u2_uk_n369, u2_uk_n373, u2_uk_n376, u2_uk_n379, u2_uk_n385, u2_uk_n407, u2_uk_n408, u2_uk_n415, 
      u2_uk_n421, u2_uk_n443, u2_uk_n456, u2_uk_n467, u2_uk_n500, u2_uk_n503, u2_uk_n504, u2_uk_n520, u2_uk_n526, 
      u2_uk_n551, u2_uk_n586, u2_uk_n608, u2_uk_n665, u2_uk_n677, u2_uk_n682, u2_uk_n689, u2_uk_n692, u2_uk_n694, 
      u2_uk_n702, u2_uk_n931, u2_uk_n933, u2_uk_n939, u2_uk_n942, u2_uk_n943, u2_uk_n944, u2_uk_n946, u2_uk_n947, 
      u2_uk_n948, u2_uk_n954, u2_uk_n955, u2_uk_n956, u2_uk_n961, u2_uk_n967, u2_uk_n970, u2_uk_n972, u2_uk_n984, 
      u2_uk_n986, u2_uk_n991, u2_uk_n994, u2_uk_n997 );
  des_des_die_1 u1 ( u0_K10_25, u0_K10_32, u0_K10_36, u0_K11_48, u0_K13_30, u0_K13_36, u0_K13_38, u0_K14_23, u0_K15_47, 
      u0_L8_17, u0_L8_23, u0_L8_31, u0_L8_9, u0_R11_10, u0_R11_11, u0_R11_12, u0_R11_13, u0_R11_14, 
      u0_R11_15, u0_R11_16, u0_R11_17, u0_R11_20, u0_R11_21, u0_R11_22, u0_R11_23, u0_R11_24, u0_R11_25, 
      u0_R11_28, u0_R11_8, u0_R11_9, u0_R12_12, u0_R12_13, u0_R12_16, u0_R12_19, u0_R12_20, u0_R12_21, 
      u0_R13_1, u0_R13_24, u0_R13_25, u0_R13_26, u0_R13_27, u0_R13_28, u0_R13_29, u0_R13_30, u0_R13_31, 
      u0_R13_32, u0_R6_24, u0_R6_26, u0_R6_27, u0_R6_28, u0_R6_29, u0_R8_1, u0_R8_16, u0_R8_17, 
      u0_R8_19, u0_R8_2, u0_R8_20, u0_R8_21, u0_R8_22, u0_R8_24, u0_R8_25, u0_R8_27, u0_R8_29, 
      u0_R8_3, u0_R8_30, u0_R8_32, u0_R8_4, u0_R8_5, u0_R9_1, u0_R9_28, u0_R9_29, u0_R9_31, 
      u0_R9_32, u0_u10_X_45, u0_u12_X_27, u0_u12_X_28, u0_u12_X_39, u0_u12_X_40, u0_u12_X_42, u0_u13_X_21, u0_u13_X_22, 
      u0_u13_X_24, u0_u13_X_26, u0_u13_X_27, u0_u7_X_38, u0_u9_X_27, u0_u9_X_34, u0_u9_X_39, u0_u9_X_41, u0_u9_X_43, 
      u0_u9_X_46, u0_uk_K_r11_11, u0_uk_K_r11_20, u0_uk_K_r11_27, u0_uk_K_r11_33, u0_uk_K_r11_48, u0_uk_K_r11_6, u0_uk_K_r12_25, u0_uk_K_r12_33, 
      u0_uk_K_r12_44, u0_uk_K_r13_35, u0_uk_K_r6_14, u0_uk_K_r6_22, u0_uk_K_r6_31, u0_uk_K_r6_7, u0_uk_K_r8_16, u0_uk_K_r8_2, u0_uk_K_r8_22, 
      u0_uk_K_r8_37, u0_uk_K_r8_41, u0_uk_K_r9_45, u0_uk_K_r9_9, u0_uk_n10, u0_uk_n100, u0_uk_n1008, u0_uk_n1009, u0_uk_n1012, 
      u0_uk_n1021, u0_uk_n104, u0_uk_n106, u0_uk_n108, u0_uk_n109, u0_uk_n11, u0_uk_n110, u0_uk_n112, u0_uk_n113, 
      u0_uk_n115, u0_uk_n116, u0_uk_n117, u0_uk_n12, u0_uk_n120, u0_uk_n121, u0_uk_n122, u0_uk_n123, u0_uk_n124, 
      u0_uk_n126, u0_uk_n127, u0_uk_n128, u0_uk_n129, u0_uk_n13, u0_uk_n130, u0_uk_n132, u0_uk_n135, u0_uk_n141, 
      u0_uk_n142, u0_uk_n145, u0_uk_n146, u0_uk_n148, u0_uk_n155, u0_uk_n161, u0_uk_n162, u0_uk_n17, u0_uk_n182, 
      u0_uk_n184, u0_uk_n185, u0_uk_n187, u0_uk_n191, u0_uk_n203, u0_uk_n205, u0_uk_n207, u0_uk_n208, u0_uk_n209, 
      u0_uk_n21, u0_uk_n213, u0_uk_n214, u0_uk_n217, u0_uk_n22, u0_uk_n220, u0_uk_n222, u0_uk_n226, u0_uk_n227, 
      u0_uk_n23, u0_uk_n231, u0_uk_n232, u0_uk_n233, u0_uk_n235, u0_uk_n238, u0_uk_n239, u0_uk_n240, u0_uk_n241, 
      u0_uk_n242, u0_uk_n243, u0_uk_n244, u0_uk_n246, u0_uk_n248, u0_uk_n249, u0_uk_n250, u0_uk_n255, u0_uk_n258, 
      u0_uk_n260, u0_uk_n261, u0_uk_n263, u0_uk_n264, u0_uk_n266, u0_uk_n267, u0_uk_n269, u0_uk_n27, u0_uk_n3, 
      u0_uk_n31, u0_uk_n327, u0_uk_n332, u0_uk_n333, u0_uk_n34, u0_uk_n341, u0_uk_n348, u0_uk_n39, u0_uk_n4, 
      u0_uk_n40, u0_uk_n41, u0_uk_n5, u0_uk_n50, u0_uk_n51, u0_uk_n61, u0_uk_n63, u0_uk_n67, u0_uk_n69, 
      u0_uk_n748, u0_uk_n75, u0_uk_n77, u0_uk_n82, u0_uk_n83, u0_uk_n88, u0_uk_n9, u0_uk_n91, u0_uk_n915, 
      u0_uk_n916, u0_uk_n92, u0_uk_n93, u0_uk_n948, u0_uk_n949, u0_uk_n95, u0_uk_n950, u0_uk_n953, u0_uk_n98, 
      u0_uk_n985, u1_FP_46, u1_FP_47, u1_FP_49, u1_FP_50, u1_FP_51, u1_K10_34, u1_K11_1, u1_K11_3, 
      u1_K11_4, u1_K11_45, u1_K11_6, u1_K12_33, u1_K12_34, u1_K12_36, u1_K12_38, u1_K12_39, u1_K12_40, 
      u1_K12_41, u1_K12_43, u1_K12_45, u1_K12_46, u1_K13_8, u1_K13_9, u1_K14_10, u1_K14_12, u1_K14_14, 
      u1_K14_15, u1_K14_16, u1_K14_21, u1_K14_22, u1_K14_27, u1_K14_28, u1_K14_29, u1_K14_31, u1_K14_33, 
      u1_K14_9, u1_K15_10, u1_K15_12, u1_K15_3, u1_K15_33, u1_K15_34, u1_K15_4, u1_K15_5, u1_K15_6, 
      u1_K15_7, u1_K15_9, u1_K16_21, u1_K16_22, u1_K16_24, u1_K16_26, u1_K16_27, u1_K16_28, u1_K1_34, 
      u1_K2_21, u1_K2_22, u1_K2_39, u1_K2_40, u1_K4_15, u1_K4_16, u1_K4_17, u1_K4_18, u1_K4_19, 
      u1_K4_21, u1_K4_22, u1_K4_24, u1_K4_27, u1_K4_28, u1_K4_39, u1_K4_40, u1_K5_15, u1_K5_16, 
      u1_K5_18, u1_K5_21, u1_K5_23, u1_K5_24, u1_K5_25, u1_K5_26, u1_K5_28, u1_K5_29, u1_K5_30, 
      u1_K5_31, u1_K5_32, u1_K5_33, u1_K5_34, u1_K5_37, u1_K5_38, u1_K5_39, u1_K5_40, u1_K5_41, 
      u1_K5_45, u1_K5_46, u1_K7_10, u1_K7_11, u1_K7_14, u1_K7_15, u1_K7_16, u1_K7_17, u1_K7_18, 
      u1_K7_19, u1_K7_21, u1_K7_22, u1_K7_23, u1_K7_26, u1_K7_28, u1_K7_29, u1_K7_3, u1_K7_30, 
      u1_K7_31, u1_K7_33, u1_K7_4, u1_K7_5, u1_K7_7, u1_K7_9, u1_K8_10, u1_K8_11, u1_K8_13, 
      u1_K8_14, u1_K8_16, u1_K8_18, u1_K8_20, u1_K8_21, u1_K8_22, u1_K8_23, u1_K8_25, u1_K8_27, 
      u1_K8_28, u1_K8_4, u1_K8_5, u1_K8_6, u1_K8_7, u1_K8_8, u1_K8_9, u1_K9_13, u1_K9_15, 
      u1_K9_16, u1_K9_17, u1_K9_21, u1_K9_23, u1_K9_24, u1_K9_25, u1_K9_28, u1_R0_14, u1_R0_15, 
      u1_R0_26, u1_R0_27, u1_R10_22, u1_R10_23, u1_R10_25, u1_R10_26, u1_R10_27, u1_R10_28, u1_R10_30, 
      u1_R10_31, u1_R11_5, u1_R11_6, u1_R11_7, u1_R12_10, u1_R12_11, u1_R12_14, u1_R12_15, u1_R12_18, 
      u1_R12_19, u1_R12_20, u1_R12_22, u1_R12_23, u1_R12_6, u1_R12_7, u1_R12_9, u1_R13_2, u1_R13_22, 
      u1_R13_23, u1_R13_3, u1_R13_4, u1_R13_5, u1_R13_6, u1_R13_7, u1_R13_9, u1_R2_10, u1_R2_11, 
      u1_R2_12, u1_R2_13, u1_R2_14, u1_R2_15, u1_R2_16, u1_R2_17, u1_R2_18, u1_R2_19, u1_R2_26, 
      u1_R2_27, u1_R3_10, u1_R3_11, u1_R3_13, u1_R3_14, u1_R3_15, u1_R3_16, u1_R3_17, u1_R3_18, 
      u1_R3_19, u1_R3_20, u1_R3_21, u1_R3_22, u1_R3_23, u1_R3_24, u1_R3_25, u1_R3_26, u1_R3_27, 
      u1_R3_28, u1_R3_30, u1_R3_31, u1_R5_10, u1_R5_11, u1_R5_12, u1_R5_13, u1_R5_14, u1_R5_15, 
      u1_R5_16, u1_R5_17, u1_R5_18, u1_R5_19, u1_R5_2, u1_R5_20, u1_R5_21, u1_R5_22, u1_R5_23, 
      u1_R5_3, u1_R5_4, u1_R5_5, u1_R5_6, u1_R5_7, u1_R5_8, u1_R5_9, u1_R6_10, u1_R6_11, 
      u1_R6_13, u1_R6_14, u1_R6_15, u1_R6_16, u1_R6_18, u1_R6_19, u1_R6_2, u1_R6_3, u1_R6_4, 
      u1_R6_5, u1_R6_6, u1_R6_7, u1_R6_8, u1_R6_9, u1_R7_10, u1_R7_11, u1_R7_12, u1_R7_13, 
      u1_R7_14, u1_R7_15, u1_R7_16, u1_R7_17, u1_R7_18, u1_R7_19, u1_R7_8, u1_R8_22, u1_R8_23, 
      u1_R9_2, u1_R9_3, u1_R9_30, u1_R9_31, u1_R9_32, u1_R9_5, u1_desIn_r_43, u1_desIn_r_51, u1_u0_X_31, 
      u1_u0_X_32, u1_u0_X_35, u1_u0_X_36, u1_u10_X_2, u1_u10_X_43, u1_u10_X_44, u1_u10_X_48, u1_u10_X_5, u1_u11_X_31, 
      u1_u11_X_32, u1_u11_X_35, u1_u11_X_37, u1_u11_X_42, u1_u11_X_44, u1_u11_X_47, u1_u11_X_48, u1_u12_X_11, u1_u12_X_12, 
      u1_u12_X_7, u1_u13_X_11, u1_u13_X_13, u1_u13_X_17, u1_u13_X_18, u1_u13_X_19, u1_u13_X_20, u1_u13_X_23, u1_u13_X_24, 
      u1_u13_X_25, u1_u13_X_26, u1_u13_X_30, u1_u13_X_32, u1_u13_X_35, u1_u13_X_36, u1_u13_X_7, u1_u13_X_8, u1_u14_X_1, 
      u1_u14_X_11, u1_u14_X_2, u1_u14_X_31, u1_u14_X_32, u1_u14_X_35, u1_u14_X_36, u1_u15_X_19, u1_u15_X_20, u1_u15_X_23, 
      u1_u15_X_25, u1_u15_X_29, u1_u15_X_30, u1_u1_X_19, u1_u1_X_20, u1_u1_X_23, u1_u1_X_24, u1_u1_X_37, u1_u1_X_38, 
      u1_u1_X_41, u1_u1_X_42, u1_u3_X_13, u1_u3_X_14, u1_u3_X_29, u1_u3_X_30, u1_u3_X_37, u1_u3_X_38, u1_u3_X_41, 
      u1_u3_X_42, u1_u4_X_13, u1_u4_X_14, u1_u4_X_17, u1_u4_X_19, u1_u4_X_42, u1_u4_X_44, u1_u4_X_47, u1_u4_X_48, 
      u1_u6_X_1, u1_u6_X_2, u1_u6_X_35, u1_u6_X_36, u1_u7_X_1, u1_u7_X_17, u1_u7_X_19, u1_u7_X_2, u1_u7_X_24, 
      u1_u7_X_26, u1_u7_X_29, u1_u7_X_30, u1_u8_X_14, u1_u8_X_29, u1_u8_X_30, u1_u9_X_31, u1_u9_X_32, u1_u9_X_35, 
      u1_u9_X_36, u1_uk_n1011, u1_uk_n1054, u1_uk_n1056, u1_uk_n1057, u1_uk_n1058, u1_uk_n1073, u1_uk_n1074, u1_uk_n1076, 
      u1_uk_n1079, u1_uk_n1080, u1_uk_n1083, u1_uk_n1105, u1_uk_n1106, u1_uk_n1109, u1_uk_n1113, u1_uk_n1114, u1_uk_n1115, 
      u1_uk_n1118, u1_uk_n1119, u1_uk_n1125, u1_uk_n1126, u1_uk_n1128, u1_uk_n1130, u1_uk_n1140, u1_uk_n1153, u1_uk_n1154, 
      u1_uk_n1156, u1_uk_n1157, u1_uk_n1158, u1_uk_n1159, u1_uk_n349, u1_uk_n468, u1_uk_n472, u1_uk_n671, u1_uk_n955, 
      u1_uk_n976, u2_K10_42, u2_K1_19, u2_K1_24, u2_K2_43, u2_K2_47, u2_K2_48, u2_R0_1, u2_R0_28, 
      u2_R0_32, u2_R12_17, u2_R8_24, u2_R8_25, u2_R8_26, u2_R8_27, u2_R8_28, u2_R8_29, u2_desIn_r_15, 
      u2_desIn_r_23, u2_desIn_r_29, u2_desIn_r_3, u2_desIn_r_37, u2_desIn_r_39, u2_desIn_r_45, u2_desIn_r_5, u2_desIn_r_53, u2_desIn_r_55, 
      u2_desIn_r_57, u2_desIn_r_61, u2_desIn_r_63, u2_desIn_r_7, u2_key_r_10, u2_key_r_11, u2_key_r_12, u2_key_r_17, u2_key_r_19, 
      u2_key_r_24, u2_key_r_25, u2_key_r_26, u2_key_r_3, u2_key_r_32, u2_key_r_33, u2_key_r_34, u2_key_r_40, u2_key_r_41, 
      u2_key_r_46, u2_key_r_47, u2_key_r_48, u2_key_r_53, u2_key_r_55, u2_key_r_6, u2_u0_X_15, u2_u0_X_16, u2_u0_X_5, 
      u2_u0_X_7, u2_u0_X_9, u2_u13_X_19, u2_u13_X_20, u2_u13_X_21, u2_u13_X_22, u2_u13_X_23, u2_u1_X_44, u2_u1_X_45, 
      u2_u1_X_46, u2_uk_K_r12_41, u2_uk_K_r8_2, u2_uk_K_r8_22, u2_uk_n10, u2_uk_n100, u2_uk_n109, u2_uk_n11, u2_uk_n1145, 
      u2_uk_n117, u2_uk_n118, u2_uk_n142, u2_uk_n145, u2_uk_n1594, u2_uk_n161, u2_uk_n1622, u2_uk_n17, u2_uk_n1782, 
      u2_uk_n182, u2_uk_n191, u2_uk_n202, u2_uk_n203, u2_uk_n207, u2_uk_n209, u2_uk_n214, u2_uk_n220, u2_uk_n231, 
      u2_uk_n238, u2_uk_n27, u2_uk_n299, u2_uk_n301, u2_uk_n305, u2_uk_n63, u2_uk_n83, u2_uk_n93, u2_uk_n94, 
      u2_uk_n967, u2_uk_n970, u2_uk_n972, u0_N296, u0_N304, u0_N310, u0_N318, u0_out10_15, u0_out10_21, 
      u0_out10_27, u0_out10_5, u0_out12_1, u0_out12_10, u0_out12_11, u0_out12_12, u0_out12_14, u0_out12_16, u0_out12_19, 
      u0_out12_20, u0_out12_22, u0_out12_24, u0_out12_25, u0_out12_26, u0_out12_29, u0_out12_3, u0_out12_30, u0_out12_32, 
      u0_out12_4, u0_out12_6, u0_out12_7, u0_out12_8, u0_out13_1, u0_out13_10, u0_out13_14, u0_out13_20, u0_out13_25, 
      u0_out13_26, u0_out13_3, u0_out13_8, u0_out14_12, u0_out14_15, u0_out14_21, u0_out14_22, u0_out14_27, u0_out14_32, 
      u0_out14_5, u0_out14_7, u0_out7_12, u0_out7_22, u0_out7_32, u0_out7_7, u0_out9_11, u0_out9_12, u0_out9_14, 
      u0_out9_15, u0_out9_19, u0_out9_21, u0_out9_22, u0_out9_25, u0_out9_27, u0_out9_29, u0_out9_3, u0_out9_32, 
      u0_out9_4, u0_out9_5, u0_out9_7, u0_out9_8, u0_uk_n102, u0_uk_n118, u0_uk_n223, u0_uk_n94, u1_out0_11, 
      u1_out0_19, u1_out0_29, u1_out0_4, u1_out10_15, u1_out10_17, u1_out10_21, u1_out10_23, u1_out10_27, u1_out10_31, 
      u1_out10_5, u1_out10_9, u1_out11_11, u1_out11_12, u1_out11_15, u1_out11_19, u1_out11_21, u1_out11_22, u1_out11_27, 
      u1_out11_29, u1_out11_32, u1_out11_4, u1_out11_5, u1_out11_7, u1_out12_13, u1_out12_18, u1_out12_2, u1_out12_28, 
      u1_out13_1, u1_out13_10, u1_out13_11, u1_out13_13, u1_out13_14, u1_out13_16, u1_out13_18, u1_out13_19, u1_out13_2, 
      u1_out13_20, u1_out13_24, u1_out13_25, u1_out13_26, u1_out13_28, u1_out13_29, u1_out13_3, u1_out13_30, u1_out13_4, 
      u1_out13_6, u1_out13_8, u1_out14_11, u1_out14_13, u1_out14_17, u1_out14_18, u1_out14_19, u1_out14_2, u1_out14_23, 
      u1_out14_28, u1_out14_29, u1_out14_31, u1_out14_4, u1_out14_9, u1_out15_1, u1_out15_10, u1_out15_14, u1_out15_20, 
      u1_out15_25, u1_out15_26, u1_out15_3, u1_out15_8, u1_out1_1, u1_out1_10, u1_out1_12, u1_out1_20, u1_out1_22, 
      u1_out1_26, u1_out1_32, u1_out1_7, u1_out3_1, u1_out3_10, u1_out3_12, u1_out3_14, u1_out3_16, u1_out3_20, 
      u1_out3_22, u1_out3_24, u1_out3_25, u1_out3_26, u1_out3_3, u1_out3_30, u1_out3_32, u1_out3_6, u1_out3_7, 
      u1_out3_8, u1_out4_1, u1_out4_10, u1_out4_11, u1_out4_12, u1_out4_14, u1_out4_15, u1_out4_16, u1_out4_19, 
      u1_out4_20, u1_out4_21, u1_out4_22, u1_out4_24, u1_out4_25, u1_out4_26, u1_out4_27, u1_out4_29, u1_out4_3, 
      u1_out4_30, u1_out4_32, u1_out4_4, u1_out4_5, u1_out4_6, u1_out4_7, u1_out4_8, u1_out6_1, u1_out6_10, 
      u1_out6_11, u1_out6_13, u1_out6_14, u1_out6_16, u1_out6_17, u1_out6_18, u1_out6_19, u1_out6_2, u1_out6_20, 
      u1_out6_23, u1_out6_24, u1_out6_25, u1_out6_26, u1_out6_28, u1_out6_29, u1_out6_3, u1_out6_30, u1_out6_31, 
      u1_out6_4, u1_out6_6, u1_out6_8, u1_out6_9, u1_out7_1, u1_out7_10, u1_out7_13, u1_out7_14, u1_out7_16, 
      u1_out7_17, u1_out7_18, u1_out7_2, u1_out7_20, u1_out7_23, u1_out7_24, u1_out7_25, u1_out7_26, u1_out7_28, 
      u1_out7_3, u1_out7_30, u1_out7_31, u1_out7_6, u1_out7_8, u1_out7_9, u1_out8_1, u1_out8_10, u1_out8_14, 
      u1_out8_16, u1_out8_20, u1_out8_24, u1_out8_25, u1_out8_26, u1_out8_3, u1_out8_30, u1_out8_6, u1_out8_8, 
      u1_out9_11, u1_out9_19, u1_out9_29, u1_out9_4, u2_out0_1, u2_out0_10, u2_out0_13, u2_out0_16, u2_out0_17, 
      u2_out0_18, u2_out0_2, u2_out0_20, u2_out0_23, u2_out0_24, u2_out0_26, u2_out0_28, u2_out0_30, u2_out0_31, 
      u2_out0_6, u2_out0_9, u2_out13_1, u2_out13_10, u2_out13_20, u2_out13_26, u2_out1_15, u2_out1_21, u2_out1_27, 
      u2_out1_5, u2_out9_12, u2_out9_22, u2_out9_32, u2_out9_7, u2_uk_n1146, u2_uk_n1161, u2_uk_n1167, u2_uk_n1168, 
      u2_uk_n1179 );
  des_des_die_2 u2 ( u0_K11_25, u0_K11_37, u0_K15_18, u0_K1_13, u0_K1_14, u0_K1_17, u0_K2_17, u0_K3_12, u0_K3_13, 
      u0_K3_14, u0_K3_17, u0_K3_18, u0_K3_19, u0_K3_23, u0_K3_5, u0_K3_6, u0_K5_1, u0_K5_3, 
      u0_K5_31, u0_K5_32, u0_K5_4, u0_K5_41, u0_K5_44, u0_K5_47, u0_K5_48, u0_K8_1, u0_K8_11, 
      u0_K8_13, u0_L13_1, u0_L13_10, u0_L13_13, u0_L13_18, u0_L13_2, u0_L13_20, u0_L13_26, u0_L13_28, 
      u0_L3_15, u0_L3_17, u0_L3_21, u0_L3_23, u0_L3_27, u0_L3_31, u0_L3_5, u0_L3_9, u0_R0_12, 
      u0_R0_14, u0_R0_17, u0_R13_1, u0_R13_11, u0_R13_12, u0_R13_13, u0_R13_14, u0_R13_15, u0_R13_16, 
      u0_R13_17, u0_R13_18, u0_R13_19, u0_R13_2, u0_R13_20, u0_R13_21, u0_R13_22, u0_R13_23, u0_R13_24, 
      u0_R13_25, u0_R13_3, u0_R13_32, u0_R13_4, u0_R13_5, u0_R13_6, u0_R13_7, u0_R13_8, u0_R13_9, 
      u0_R1_1, u0_R1_12, u0_R1_13, u0_R1_16, u0_R1_17, u0_R1_18, u0_R1_19, u0_R1_20, u0_R1_21, 
      u0_R1_22, u0_R1_24, u0_R1_25, u0_R1_26, u0_R1_27, u0_R1_28, u0_R1_29, u0_R1_3, u0_R1_31, 
      u0_R1_32, u0_R1_4, u0_R1_5, u0_R1_8, u0_R1_9, u0_R3_1, u0_R3_2, u0_R3_20, u0_R3_21, 
      u0_R3_22, u0_R3_24, u0_R3_27, u0_R3_28, u0_R3_29, u0_R3_3, u0_R3_30, u0_R3_31, u0_R3_32, 
      u0_R3_4, u0_R3_5, u0_R4_1, u0_R4_22, u0_R4_24, u0_R4_29, u0_R4_30, u0_R6_1, u0_R6_10, 
      u0_R6_11, u0_R6_12, u0_R6_13, u0_R6_2, u0_R6_32, u0_R6_4, u0_R6_5, u0_R6_7, u0_R6_8, 
      u0_R6_9, u0_R9_1, u0_R9_16, u0_R9_17, u0_R9_18, u0_R9_19, u0_R9_2, u0_R9_20, u0_R9_21, 
      u0_R9_22, u0_R9_23, u0_R9_24, u0_R9_25, u0_R9_27, u0_R9_28, u0_R9_29, u0_R9_3, u0_R9_32, 
      u0_R9_4, u0_R9_5, u0_R9_6, u0_R9_7, u0_R9_8, u0_R9_9, u0_desIn_r_15, u0_desIn_r_29, u0_desIn_r_3, 
      u0_desIn_r_31, u0_desIn_r_37, u0_desIn_r_39, u0_desIn_r_45, u0_desIn_r_47, u0_desIn_r_5, u0_desIn_r_53, u0_desIn_r_55, u0_desIn_r_57, 
      u0_desIn_r_63, u0_desIn_r_7, u0_key_r_11, u0_key_r_12, u0_key_r_13, u0_key_r_17, u0_key_r_19, u0_key_r_20, u0_key_r_24, 
      u0_key_r_25, u0_key_r_26, u0_key_r_27, u0_key_r_32, u0_key_r_34, u0_key_r_39, u0_key_r_4, u0_key_r_40, u0_key_r_41, 
      u0_key_r_47, u0_key_r_48, u0_key_r_5, u0_key_r_54, u0_key_r_55, u0_key_r_6, u0_u0_X_15, u0_u0_X_16, u0_u0_X_23, 
      u0_u0_X_4, u0_u10_X_39, u0_u14_X_15, u0_u1_X_13, u0_u1_X_14, u0_u1_X_15, u0_u1_X_16, u0_u1_X_18, u0_u1_X_20, 
      u0_u1_X_22, u0_u1_X_23, u0_u2_X_10, u0_u2_X_15, u0_u2_X_16, u0_u2_X_21, u0_u2_X_22, u0_u2_X_3, u0_u2_X_34, 
      u0_u2_X_45, u0_u2_X_9, u0_u4_X_34, u0_u4_X_36, u0_u4_X_38, u0_u4_X_39, u0_u5_X_1, u0_u5_X_3, u0_u5_X_31, 
      u0_u5_X_32, u0_u5_X_34, u0_u5_X_36, u0_u5_X_38, u0_u5_X_39, u0_u5_X_4, u0_u5_X_40, u0_u5_X_41, u0_u5_X_43, 
      u0_u5_X_46, u0_u5_X_47, u0_u5_X_5, u0_u5_X_6, u0_u7_X_4, u0_u7_X_9, u0_uk_K_r13_0, u0_uk_K_r13_13, u0_uk_K_r13_17, 
      u0_uk_K_r13_22, u0_uk_K_r13_25, u0_uk_K_r13_32, u0_uk_K_r13_38, u0_uk_K_r13_4, u0_uk_K_r13_44, u0_uk_K_r13_55, u0_uk_K_r1_15, u0_uk_K_r1_21, 
      u0_uk_K_r1_22, u0_uk_K_r1_42, u0_uk_K_r1_44, u0_uk_K_r1_7, u0_uk_K_r3_10, u0_uk_K_r3_14, u0_uk_K_r3_15, u0_uk_K_r3_38, u0_uk_K_r3_9, 
      u0_uk_K_r4_38, u0_uk_K_r6_10, u0_uk_K_r6_26, u0_uk_K_r6_27, u0_uk_K_r6_3, u0_uk_K_r6_34, u0_uk_K_r6_46, u0_uk_K_r6_53, u0_uk_K_r9_0, 
      u0_uk_K_r9_1, u0_uk_K_r9_19, u0_uk_K_r9_25, u0_uk_K_r9_31, u0_uk_K_r9_33, u0_uk_K_r9_35, u0_uk_K_r9_45, u0_uk_K_r9_49, u0_uk_K_r9_6, 
      u0_uk_K_r9_9, u0_uk_n1, u0_uk_n10, u0_uk_n100, u0_uk_n1004, u0_uk_n102, u0_uk_n110, u0_uk_n117, u0_uk_n118, 
      u0_uk_n12, u0_uk_n128, u0_uk_n129, u0_uk_n13, u0_uk_n14, u0_uk_n146, u0_uk_n147, u0_uk_n148, u0_uk_n15, 
      u0_uk_n155, u0_uk_n16, u0_uk_n161, u0_uk_n164, u0_uk_n17, u0_uk_n18, u0_uk_n181, u0_uk_n182, u0_uk_n183, 
      u0_uk_n184, u0_uk_n185, u0_uk_n186, u0_uk_n187, u0_uk_n189, u0_uk_n19, u0_uk_n193, u0_uk_n194, u0_uk_n195, 
      u0_uk_n197, u0_uk_n198, u0_uk_n199, u0_uk_n20, u0_uk_n200, u0_uk_n201, u0_uk_n203, u0_uk_n204, u0_uk_n205, 
      u0_uk_n206, u0_uk_n207, u0_uk_n208, u0_uk_n21, u0_uk_n210, u0_uk_n212, u0_uk_n214, u0_uk_n215, u0_uk_n216, 
      u0_uk_n218, u0_uk_n219, u0_uk_n222, u0_uk_n223, u0_uk_n224, u0_uk_n225, u0_uk_n23, u0_uk_n230, u0_uk_n231, 
      u0_uk_n238, u0_uk_n24, u0_uk_n240, u0_uk_n25, u0_uk_n250, u0_uk_n251, u0_uk_n252, u0_uk_n257, u0_uk_n26, 
      u0_uk_n27, u0_uk_n28, u0_uk_n29, u0_uk_n30, u0_uk_n31, u0_uk_n318, u0_uk_n32, u0_uk_n324, u0_uk_n329, 
      u0_uk_n33, u0_uk_n330, u0_uk_n331, u0_uk_n336, u0_uk_n337, u0_uk_n339, u0_uk_n343, u0_uk_n344, u0_uk_n35, 
      u0_uk_n352, u0_uk_n358, u0_uk_n36, u0_uk_n37, u0_uk_n38, u0_uk_n39, u0_uk_n4, u0_uk_n41, u0_uk_n412, 
      u0_uk_n413, u0_uk_n418, u0_uk_n419, u0_uk_n42, u0_uk_n420, u0_uk_n425, u0_uk_n429, u0_uk_n43, u0_uk_n430, 
      u0_uk_n434, u0_uk_n44, u0_uk_n45, u0_uk_n455, u0_uk_n457, u0_uk_n458, u0_uk_n466, u0_uk_n471, u0_uk_n475, 
      u0_uk_n476, u0_uk_n486, u0_uk_n488, u0_uk_n490, u0_uk_n491, u0_uk_n493, u0_uk_n494, u0_uk_n5, u0_uk_n543, 
      u0_uk_n544, u0_uk_n545, u0_uk_n546, u0_uk_n547, u0_uk_n549, u0_uk_n550, u0_uk_n552, u0_uk_n553, u0_uk_n554, 
      u0_uk_n555, u0_uk_n557, u0_uk_n558, u0_uk_n559, u0_uk_n560, u0_uk_n561, u0_uk_n562, u0_uk_n565, u0_uk_n566, 
      u0_uk_n568, u0_uk_n570, u0_uk_n573, u0_uk_n574, u0_uk_n575, u0_uk_n578, u0_uk_n579, u0_uk_n580, u0_uk_n581, 
      u0_uk_n6, u0_uk_n60, u0_uk_n609, u0_uk_n620, u0_uk_n624, u0_uk_n7, u0_uk_n759, u0_uk_n793, u0_uk_n8, 
      u0_uk_n805, u0_uk_n810, u0_uk_n851, u0_uk_n864, u0_uk_n917, u0_uk_n918, u0_uk_n94, u0_uk_n982, u0_uk_n99, 
      u0_uk_n990, u0_uk_n992, u1_FP_42, u1_FP_43, u1_FP_58, u1_FP_59, u1_K10_10, u1_K10_27, u1_K10_28, 
      u1_K13_33, u1_K13_34, u1_K13_35, u1_K13_36, u1_K13_37, u1_K13_38, u1_K13_39, u1_K13_40, u1_K14_3, 
      u1_K14_4, u1_K15_27, u1_K15_28, u1_K15_45, u1_K15_46, u1_K16_15, u1_K16_16, u1_K16_39, u1_K16_40, 
      u1_K1_12, u1_K1_14, u1_K1_15, u1_K1_16, u1_K1_39, u1_K1_40, u1_K1_43, u1_K1_45, u1_K1_46, 
      u1_K1_9, u1_K2_1, u1_K2_3, u1_K2_4, u1_K2_45, u1_K2_46, u1_K2_47, u1_K3_15, u1_K3_16, 
      u1_K3_27, u1_K3_28, u1_K3_39, u1_K3_40, u1_K4_9, u1_K7_39, u1_K7_40, u1_K7_41, u1_K7_43, 
      u1_K7_45, u1_K9_3, u1_K9_34, u1_K9_36, u1_K9_37, u1_K9_38, u1_K9_39, u1_K9_4, u1_K9_40, 
      u1_R0_18, u1_R0_19, u1_R0_2, u1_R0_3, u1_R0_30, u1_R0_31, u1_R0_32, u1_R11_22, u1_R11_23, 
      u1_R11_24, u1_R11_25, u1_R11_26, u1_R11_27, u1_R12_2, u1_R12_3, u1_R13_18, u1_R13_19, u1_R13_30, 
      u1_R13_31, u1_R1_10, u1_R1_11, u1_R1_18, u1_R1_19, u1_R1_26, u1_R1_27, u1_R2_6, u1_R2_7, 
      u1_R5_26, u1_R5_27, u1_R5_28, u1_R5_30, u1_R5_31, u1_R7_2, u1_R7_22, u1_R7_23, u1_R7_24, 
      u1_R7_25, u1_R7_26, u1_R7_27, u1_R7_3, u1_R8_18, u1_R8_19, u1_R8_6, u1_R8_7, u1_desIn_r_13, 
      u1_desIn_r_17, u1_desIn_r_21, u1_desIn_r_25, u1_desIn_r_33, u1_desIn_r_41, u1_desIn_r_47, u1_desIn_r_49, u1_desIn_r_5, u1_desIn_r_55, 
      u1_desIn_r_9, u1_u0_X_11, u1_u0_X_13, u1_u0_X_17, u1_u0_X_18, u1_u0_X_37, u1_u0_X_38, u1_u0_X_47, u1_u0_X_48, 
      u1_u0_X_7, u1_u0_X_8, u1_u12_X_31, u1_u12_X_32, u1_u12_X_41, u1_u12_X_42, u1_u13_X_1, u1_u13_X_2, u1_u13_X_5, 
      u1_u13_X_6, u1_u14_X_25, u1_u14_X_26, u1_u14_X_29, u1_u14_X_30, u1_u14_X_43, u1_u14_X_44, u1_u14_X_47, u1_u14_X_48, 
      u1_u15_X_13, u1_u15_X_14, u1_u15_X_17, u1_u15_X_18, u1_u15_X_37, u1_u15_X_38, u1_u15_X_41, u1_u15_X_42, u1_u1_X_2, 
      u1_u1_X_25, u1_u1_X_26, u1_u1_X_29, u1_u1_X_30, u1_u1_X_43, u1_u1_X_44, u1_u1_X_48, u1_u1_X_5, u1_u1_X_6, 
      u1_u2_X_13, u1_u2_X_14, u1_u2_X_17, u1_u2_X_18, u1_u2_X_25, u1_u2_X_26, u1_u2_X_29, u1_u2_X_30, u1_u2_X_37, 
      u1_u2_X_38, u1_u2_X_41, u1_u2_X_42, u1_u3_X_11, u1_u3_X_12, u1_u3_X_7, u1_u3_X_8, u1_u6_X_37, u1_u6_X_38, 
      u1_u6_X_42, u1_u6_X_44, u1_u6_X_47, u1_u6_X_48, u1_u8_X_1, u1_u8_X_2, u1_u8_X_31, u1_u8_X_32, u1_u8_X_41, 
      u1_u8_X_42, u1_u8_X_5, u1_u8_X_6, u1_u9_X_11, u1_u9_X_12, u1_u9_X_25, u1_u9_X_26, u1_u9_X_29, u1_u9_X_30, 
      u1_u9_X_7, u1_u9_X_8, u1_uk_n1015, u1_uk_n1016, u1_uk_n1017, u1_uk_n1027, u1_uk_n1028, u1_uk_n1050, u1_uk_n1124, 
      u1_uk_n1162, u1_uk_n1163, u1_uk_n376, u1_uk_n996, u2_K15_37, u2_K15_44, u2_K15_47, u2_K15_48, u2_K2_1, 
      u2_K2_12, u2_K2_18, u2_K2_20, u2_K8_13, u2_K8_18, u2_K8_24, u2_K8_5, u2_K8_8, u2_R0_1, 
      u2_R0_10, u2_R0_12, u2_R0_13, u2_R0_14, u2_R0_15, u2_R0_17, u2_R0_3, u2_R0_32, u2_R0_4, 
      u2_R0_5, u2_R0_6, u2_R0_7, u2_R0_8, u2_R0_9, u2_R13_1, u2_R13_24, u2_R13_25, u2_R13_27, 
      u2_R13_28, u2_R13_29, u2_R13_30, u2_R13_32, u2_R6_1, u2_R6_10, u2_R6_11, u2_R6_12, u2_R6_13, 
      u2_R6_15, u2_R6_16, u2_R6_17, u2_R6_2, u2_R6_32, u2_R6_4, u2_R6_5, u2_R6_6, u2_R6_7, 
      u2_R6_8, u2_R6_9, u2_u14_X_39, u2_u14_X_46, u2_u1_X_16, u2_u1_X_23, u2_u1_X_3, u2_u7_X_21, u2_u7_X_4, 
      u2_uk_K_r0_11, u2_uk_K_r0_17, u2_uk_K_r0_25, u2_uk_K_r0_32, u2_uk_K_r0_47, u2_uk_K_r6_10, u2_uk_K_r6_26, u2_uk_K_r6_3, u2_uk_K_r6_34, 
      u2_uk_K_r6_53, u2_uk_n10, u2_uk_n100, u2_uk_n1004, u2_uk_n1097, u2_uk_n110, u2_uk_n1100, u2_uk_n1105, u2_uk_n117, 
      u2_uk_n118, u2_uk_n1231, u2_uk_n1232, u2_uk_n1234, u2_uk_n1238, u2_uk_n1240, u2_uk_n1243, u2_uk_n1244, u2_uk_n1247, 
      u2_uk_n1249, u2_uk_n1260, u2_uk_n1261, u2_uk_n1267, u2_uk_n1270, u2_uk_n1275, u2_uk_n128, u2_uk_n129, u2_uk_n142, 
      u2_uk_n145, u2_uk_n1500, u2_uk_n1502, u2_uk_n1506, u2_uk_n1508, u2_uk_n1513, u2_uk_n1514, u2_uk_n1515, u2_uk_n1518, 
      u2_uk_n1519, u2_uk_n1521, u2_uk_n1522, u2_uk_n1527, u2_uk_n1529, u2_uk_n1535, u2_uk_n155, u2_uk_n161, u2_uk_n162, 
      u2_uk_n164, u2_uk_n17, u2_uk_n1817, u2_uk_n182, u2_uk_n1835, u2_uk_n1837, u2_uk_n1849, u2_uk_n1853, u2_uk_n1855, 
      u2_uk_n187, u2_uk_n188, u2_uk_n191, u2_uk_n202, u2_uk_n208, u2_uk_n209, u2_uk_n213, u2_uk_n220, u2_uk_n230, 
      u2_uk_n231, u2_uk_n238, u2_uk_n27, u2_uk_n31, u2_uk_n63, u2_uk_n83, u2_uk_n92, u2_uk_n93, u2_uk_n94, 
      u2_uk_n943, u2_uk_n944, u2_uk_n99, u2_uk_n991, u2_uk_n994, u0_N132, u0_N136, u0_N142, u0_N144, 
      u0_N148, u0_N150, u0_N154, u0_N158, u0_N448, u0_N449, u0_N457, u0_N460, u0_N465, 
      u0_N467, u0_N473, u0_N475, u0_out0_1, u0_out0_10, u0_out0_13, u0_out0_16, u0_out0_17, u0_out0_18, 
      u0_out0_2, u0_out0_20, u0_out0_23, u0_out0_24, u0_out0_26, u0_out0_28, u0_out0_30, u0_out0_31, u0_out0_6, 
      u0_out0_9, u0_out10_11, u0_out10_12, u0_out10_13, u0_out10_14, u0_out10_17, u0_out10_18, u0_out10_19, u0_out10_2, 
      u0_out10_22, u0_out10_23, u0_out10_25, u0_out10_28, u0_out10_29, u0_out10_3, u0_out10_31, u0_out10_32, u0_out10_4, 
      u0_out10_7, u0_out10_8, u0_out10_9, u0_out14_11, u0_out14_14, u0_out14_16, u0_out14_17, u0_out14_19, u0_out14_23, 
      u0_out14_24, u0_out14_25, u0_out14_29, u0_out14_3, u0_out14_30, u0_out14_31, u0_out14_4, u0_out14_6, u0_out14_8, 
      u0_out14_9, u0_out1_1, u0_out1_10, u0_out1_16, u0_out1_20, u0_out1_24, u0_out1_26, u0_out1_30, u0_out1_6, 
      u0_out2_1, u0_out2_10, u0_out2_11, u0_out2_12, u0_out2_13, u0_out2_14, u0_out2_15, u0_out2_16, u0_out2_17, 
      u0_out2_18, u0_out2_19, u0_out2_2, u0_out2_20, u0_out2_21, u0_out2_22, u0_out2_23, u0_out2_24, u0_out2_25, 
      u0_out2_26, u0_out2_27, u0_out2_28, u0_out2_29, u0_out2_3, u0_out2_30, u0_out2_31, u0_out2_32, u0_out2_4, 
      u0_out2_5, u0_out2_6, u0_out2_7, u0_out2_8, u0_out2_9, u0_out4_11, u0_out4_12, u0_out4_19, u0_out4_22, 
      u0_out4_29, u0_out4_32, u0_out4_4, u0_out4_7, u0_out5_11, u0_out5_12, u0_out5_15, u0_out5_17, u0_out5_19, 
      u0_out5_21, u0_out5_22, u0_out5_23, u0_out5_27, u0_out5_29, u0_out5_31, u0_out5_32, u0_out5_4, u0_out5_5, 
      u0_out5_7, u0_out5_9, u0_out7_13, u0_out7_16, u0_out7_17, u0_out7_18, u0_out7_2, u0_out7_23, u0_out7_24, 
      u0_out7_28, u0_out7_30, u0_out7_31, u0_out7_6, u0_out7_9, u0_uk_n109, u0_uk_n11, u0_uk_n141, u0_uk_n142, 
      u0_uk_n145, u0_uk_n162, u0_uk_n163, u0_uk_n188, u0_uk_n191, u0_uk_n202, u0_uk_n209, u0_uk_n213, u0_uk_n217, 
      u0_uk_n220, u0_uk_n242, u0_uk_n63, u0_uk_n684, u0_uk_n690, u0_uk_n696, u0_uk_n697, u0_uk_n698, u0_uk_n705, 
      u0_uk_n83, u0_uk_n92, u0_uk_n93, u1_out0_12, u1_out0_13, u1_out0_15, u1_out0_16, u1_out0_18, u1_out0_2, 
      u1_out0_21, u1_out0_22, u1_out0_24, u1_out0_27, u1_out0_28, u1_out0_30, u1_out0_32, u1_out0_5, u1_out0_6, 
      u1_out0_7, u1_out12_11, u1_out12_12, u1_out12_19, u1_out12_22, u1_out12_29, u1_out12_32, u1_out12_4, u1_out12_7, 
      u1_out13_17, u1_out13_23, u1_out13_31, u1_out13_9, u1_out14_14, u1_out14_15, u1_out14_21, u1_out14_25, u1_out14_27, 
      u1_out14_3, u1_out14_5, u1_out14_8, u1_out15_12, u1_out15_16, u1_out15_22, u1_out15_24, u1_out15_30, u1_out15_32, 
      u1_out15_6, u1_out15_7, u1_out1_14, u1_out1_15, u1_out1_17, u1_out1_21, u1_out1_23, u1_out1_25, u1_out1_27, 
      u1_out1_3, u1_out1_31, u1_out1_5, u1_out1_8, u1_out1_9, u1_out2_12, u1_out2_14, u1_out2_16, u1_out2_22, 
      u1_out2_24, u1_out2_25, u1_out2_3, u1_out2_30, u1_out2_32, u1_out2_6, u1_out2_7, u1_out2_8, u1_out3_13, 
      u1_out3_18, u1_out3_2, u1_out3_28, u1_out6_12, u1_out6_15, u1_out6_21, u1_out6_22, u1_out6_27, u1_out6_32, 
      u1_out6_5, u1_out6_7, u1_out8_11, u1_out8_12, u1_out8_17, u1_out8_19, u1_out8_22, u1_out8_23, u1_out8_29, 
      u1_out8_31, u1_out8_32, u1_out8_4, u1_out8_7, u1_out8_9, u1_out9_13, u1_out9_14, u1_out9_18, u1_out9_2, 
      u1_out9_25, u1_out9_28, u1_out9_3, u1_out9_8, u2_out14_12, u2_out14_15, u2_out14_21, u2_out14_22, u2_out14_27, 
      u2_out14_32, u2_out14_5, u2_out14_7, u2_out1_1, u2_out1_10, u2_out1_13, u2_out1_16, u2_out1_17, u2_out1_18, 
      u2_out1_2, u2_out1_20, u2_out1_23, u2_out1_24, u2_out1_26, u2_out1_28, u2_out1_30, u2_out1_31, u2_out1_6, 
      u2_out1_9, u2_out7_1, u2_out7_10, u2_out7_13, u2_out7_16, u2_out7_17, u2_out7_18, u2_out7_2, u2_out7_20, 
      u2_out7_23, u2_out7_24, u2_out7_26, u2_out7_28, u2_out7_30, u2_out7_31, u2_out7_6, u2_out7_9 );
  des_des_die_3 u3 ( u0_K2_30, u0_K2_44, u0_K4_24, u0_K4_43, u0_K4_48, u0_K7_2, u0_K7_23, u0_R0_17, u0_R0_18, 
      u0_R0_19, u0_R0_21, u0_R0_22, u0_R0_25, u0_R0_27, u0_R0_28, u0_R0_29, u0_R2_1, u0_R2_12, 
      u0_R2_13, u0_R2_14, u0_R2_15, u0_R2_16, u0_R2_17, u0_R2_20, u0_R2_21, u0_R2_22, u0_R2_23, 
      u0_R2_26, u0_R2_27, u0_R2_28, u0_R2_29, u0_R2_30, u0_R2_31, u0_R2_32, u0_R5_1, u0_R5_11, 
      u0_R5_12, u0_R5_13, u0_R5_14, u0_R5_16, u0_R5_17, u0_R5_18, u0_R5_19, u0_R5_2, u0_R5_20, 
      u0_R5_21, u0_R5_22, u0_R5_23, u0_R5_24, u0_R5_25, u0_R5_26, u0_R5_27, u0_R5_28, u0_R5_29, 
      u0_R5_3, u0_R5_30, u0_R5_31, u0_R5_32, u0_R5_4, u0_R5_5, u0_R5_7, u0_R5_8, u0_R5_9, 
      u0_u1_X_25, u0_u1_X_29, u0_u1_X_31, u0_u1_X_34, u0_u1_X_35, u0_u1_X_37, u0_u1_X_39, u0_u1_X_45, u0_u1_X_46, 
      u0_u1_X_47, u0_u1_X_48, u0_u3_X_27, u0_u3_X_28, u0_u3_X_35, u0_u3_X_36, u0_u3_X_37, u0_u3_X_38, u0_u6_X_15, 
      u0_u6_X_22, u0_u6_X_9, u0_uk_K_r0_15, u0_uk_K_r0_2, u0_uk_K_r0_28, u0_uk_K_r0_31, u0_uk_K_r0_36, u0_uk_K_r0_49, u0_uk_K_r0_7, 
      u0_uk_K_r2_13, u0_uk_K_r2_18, u0_uk_K_r2_28, u0_uk_K_r2_33, u0_uk_K_r2_55, u0_uk_K_r5_10, u0_uk_K_r5_16, u0_uk_K_r5_17, u0_uk_K_r5_19, 
      u0_uk_K_r5_32, u0_uk_K_r5_37, u0_uk_K_r5_39, u0_uk_K_r5_4, u0_uk_K_r5_8, u0_uk_n10, u0_uk_n102, u0_uk_n109, u0_uk_n110, 
      u0_uk_n117, u0_uk_n118, u0_uk_n128, u0_uk_n129, u0_uk_n141, u0_uk_n142, u0_uk_n145, u0_uk_n146, u0_uk_n147, 
      u0_uk_n148, u0_uk_n161, u0_uk_n162, u0_uk_n163, u0_uk_n164, u0_uk_n17, u0_uk_n182, u0_uk_n188, u0_uk_n202, 
      u0_uk_n207, u0_uk_n208, u0_uk_n213, u0_uk_n214, u0_uk_n217, u0_uk_n223, u0_uk_n230, u0_uk_n231, u0_uk_n238, 
      u0_uk_n240, u0_uk_n250, u0_uk_n252, u0_uk_n257, u0_uk_n27, u0_uk_n31, u0_uk_n361, u0_uk_n362, u0_uk_n365, 
      u0_uk_n367, u0_uk_n368, u0_uk_n370, u0_uk_n371, u0_uk_n372, u0_uk_n374, u0_uk_n378, u0_uk_n380, u0_uk_n381, 
      u0_uk_n383, u0_uk_n384, u0_uk_n387, u0_uk_n388, u0_uk_n389, u0_uk_n392, u0_uk_n393, u0_uk_n394, u0_uk_n396, 
      u0_uk_n398, u0_uk_n399, u0_uk_n400, u0_uk_n401, u0_uk_n402, u0_uk_n403, u0_uk_n405, u0_uk_n406, u0_uk_n498, 
      u0_uk_n499, u0_uk_n506, u0_uk_n508, u0_uk_n511, u0_uk_n513, u0_uk_n514, u0_uk_n516, u0_uk_n517, u0_uk_n521, 
      u0_uk_n522, u0_uk_n523, u0_uk_n528, u0_uk_n531, u0_uk_n532, u0_uk_n537, u0_uk_n538, u0_uk_n539, u0_uk_n584, 
      u0_uk_n592, u0_uk_n593, u0_uk_n599, u0_uk_n60, u0_uk_n600, u0_uk_n612, u0_uk_n616, u0_uk_n623, u0_uk_n63, 
      u0_uk_n763, u0_uk_n765, u0_uk_n766, u0_uk_n768, u0_uk_n770, u0_uk_n771, u0_uk_n774, u0_uk_n775, u0_uk_n776, 
      u0_uk_n780, u0_uk_n783, u0_uk_n826, u0_uk_n829, u0_uk_n83, u0_uk_n831, u0_uk_n832, u0_uk_n834, u0_uk_n92, 
      u0_uk_n93, u0_uk_n94, u2_FP_33, u2_FP_34, u2_FP_35, u2_FP_36, u2_FP_37, u2_FP_40, u2_FP_41, 
      u2_FP_42, u2_FP_44, u2_FP_46, u2_FP_47, u2_FP_48, u2_FP_49, u2_FP_51, u2_FP_52, u2_FP_53, 
      u2_FP_64, u2_K10_11, u2_K10_17, u2_K10_19, u2_K10_25, u2_K10_26, u2_K10_29, u2_K10_43, u2_K10_44, 
      u2_K10_5, u2_K10_6, u2_K11_11, u2_K11_13, u2_K11_18, u2_K11_6, u2_K11_7, u2_K12_25, u2_K12_26, 
      u2_K12_8, u2_K14_42, u2_K16_26, u2_K16_5, u2_K16_6, u2_K16_8, u2_K2_29, u2_K2_36, u2_K3_13, 
      u2_K3_19, u2_K3_23, u2_K3_26, u2_K3_35, u2_K3_48, u2_K4_13, u2_K4_14, u2_K4_18, u2_K4_19, 
      u2_K4_35, u2_K5_11, u2_K5_13, u2_K5_14, u2_K5_17, u2_K5_18, u2_K5_19, u2_K5_2, u2_K5_29, 
      u2_K5_30, u2_K5_31, u2_K5_32, u2_K5_41, u2_K5_44, u2_K5_48, u2_K5_5, u2_K5_6, u2_K5_8, 
      u2_K6_11, u2_K6_13, u2_K6_19, u2_K6_20, u2_K6_23, u2_K6_24, u2_K6_25, u2_K6_36, u2_K6_48, 
      u2_K6_5, u2_K6_6, u2_K6_8, u2_K7_26, u2_K7_35, u2_K7_37, u2_K7_38, u2_K7_43, u2_K7_44, 
      u2_K7_48, u2_K7_5, u2_K7_7, u2_K9_12, u2_K9_14, u2_K9_23, u2_K9_25, u2_K9_29, u2_R0_17, 
      u2_R0_18, u2_R0_19, u2_R0_20, u2_R0_21, u2_R0_25, u2_R0_28, u2_R10_16, u2_R10_17, u2_R10_19, 
      u2_R10_21, u2_R10_4, u2_R10_5, u2_R10_7, u2_R10_8, u2_R10_9, u2_R12_17, u2_R12_18, u2_R12_20, 
      u2_R12_21, u2_R12_22, u2_R12_23, u2_R12_24, u2_R12_25, u2_R12_27, u2_R12_28, u2_R12_29, u2_R1_1, 
      u2_R1_12, u2_R1_16, u2_R1_17, u2_R1_19, u2_R1_20, u2_R1_22, u2_R1_24, u2_R1_25, u2_R1_27, 
      u2_R1_3, u2_R1_30, u2_R1_5, u2_R1_8, u2_R1_9, u2_R2_1, u2_R2_11, u2_R2_12, u2_R2_13, 
      u2_R2_16, u2_R2_17, u2_R2_2, u2_R2_20, u2_R2_21, u2_R2_24, u2_R2_28, u2_R2_3, u2_R2_32, 
      u2_R2_6, u2_R2_7, u2_R2_8, u2_R2_9, u2_R3_1, u2_R3_12, u2_R3_13, u2_R3_15, u2_R3_18, 
      u2_R3_20, u2_R3_21, u2_R3_24, u2_R3_28, u2_R3_29, u2_R3_3, u2_R3_30, u2_R3_4, u2_R3_5, 
      u2_R3_8, u2_R3_9, u2_R4_1, u2_R4_12, u2_R4_13, u2_R4_14, u2_R4_16, u2_R4_17, u2_R4_19, 
      u2_R4_20, u2_R4_24, u2_R4_25, u2_R4_26, u2_R4_28, u2_R4_29, u2_R4_4, u2_R4_5, u2_R4_6, 
      u2_R4_7, u2_R4_8, u2_R5_1, u2_R5_10, u2_R5_11, u2_R5_12, u2_R5_13, u2_R5_14, u2_R5_16, 
      u2_R5_17, u2_R5_18, u2_R5_21, u2_R5_23, u2_R5_24, u2_R5_25, u2_R5_26, u2_R5_28, u2_R5_29, 
      u2_R5_32, u2_R5_4, u2_R5_5, u2_R5_8, u2_R5_9, u2_R7_11, u2_R7_12, u2_R7_13, u2_R7_14, 
      u2_R7_15, u2_R7_16, u2_R7_17, u2_R7_20, u2_R7_21, u2_R7_4, u2_R7_5, u2_R7_6, u2_R7_7, 
      u2_R7_8, u2_R7_9, u2_R8_1, u2_R8_12, u2_R8_13, u2_R8_15, u2_R8_16, u2_R8_17, u2_R8_18, 
      u2_R8_19, u2_R8_20, u2_R8_28, u2_R8_29, u2_R8_32, u2_R8_4, u2_R8_5, u2_R8_6, u2_R8_8, 
      u2_R8_9, u2_R9_1, u2_R9_12, u2_R9_13, u2_R9_15, u2_R9_16, u2_R9_17, u2_R9_2, u2_R9_20, 
      u2_R9_21, u2_R9_24, u2_R9_25, u2_R9_32, u2_R9_4, u2_R9_5, u2_R9_8, u2_R9_9, u2_u10_X_10, 
      u2_u10_X_15, u2_u10_X_16, u2_u10_X_21, u2_u10_X_33, u2_u10_X_34, u2_u10_X_4, u2_u10_X_9, u2_u11_X_27, u2_u11_X_29, 
      u2_u11_X_31, u2_u11_X_33, u2_u11_X_34, u2_u11_X_35, u2_u11_X_36, u2_u11_X_9, u2_u13_X_25, u2_u13_X_28, u2_u13_X_39, 
      u2_u15_X_10, u2_u15_X_16, u2_u15_X_18, u2_u15_X_20, u2_u15_X_27, u2_u15_X_9, u2_u1_X_25, u2_u1_X_33, u2_u1_X_34, 
      u2_u1_X_35, u2_u1_X_37, u2_u1_X_39, u2_u1_X_40, u2_u1_X_42, u2_u2_X_1, u2_u2_X_10, u2_u2_X_15, u2_u2_X_16, 
      u2_u2_X_18, u2_u2_X_20, u2_u2_X_21, u2_u2_X_22, u2_u2_X_27, u2_u2_X_3, u2_u2_X_30, u2_u2_X_32, u2_u2_X_34, 
      u2_u2_X_39, u2_u2_X_41, u2_u2_X_42, u2_u2_X_43, u2_u2_X_44, u2_u2_X_46, u2_u2_X_47, u2_u2_X_5, u2_u2_X_7, 
      u2_u2_X_9, u2_u3_X_15, u2_u3_X_21, u2_u3_X_22, u2_u3_X_27, u2_u3_X_28, u2_u3_X_33, u2_u3_X_34, u2_u3_X_36, 
      u2_u3_X_38, u2_u3_X_39, u2_u3_X_40, u2_u3_X_42, u2_u3_X_44, u2_u3_X_45, u2_u3_X_46, u2_u3_X_5, u2_u3_X_6, 
      u2_u3_X_7, u2_u3_X_8, u2_u4_X_1, u2_u4_X_10, u2_u4_X_15, u2_u4_X_16, u2_u4_X_21, u2_u4_X_23, u2_u4_X_24, 
      u2_u4_X_25, u2_u4_X_26, u2_u4_X_28, u2_u4_X_3, u2_u4_X_33, u2_u4_X_34, u2_u4_X_36, u2_u4_X_38, u2_u4_X_39, 
      u2_u4_X_40, u2_u4_X_46, u2_u4_X_47, u2_u4_X_9, u2_u5_X_1, u2_u5_X_12, u2_u5_X_14, u2_u5_X_15, u2_u5_X_16, 
      u2_u5_X_22, u2_u5_X_27, u2_u5_X_3, u2_u5_X_30, u2_u5_X_32, u2_u5_X_33, u2_u5_X_34, u2_u5_X_4, u2_u5_X_40, 
      u2_u5_X_45, u2_u5_X_46, u2_u5_X_47, u2_u6_X_10, u2_u6_X_22, u2_u6_X_28, u2_u6_X_29, u2_u6_X_3, u2_u6_X_31, 
      u2_u6_X_33, u2_u6_X_4, u2_u6_X_40, u2_u6_X_45, u2_u6_X_46, u2_u6_X_9, u2_u8_X_15, u2_u8_X_27, u2_u8_X_28, 
      u2_u9_X_10, u2_u9_X_15, u2_u9_X_16, u2_u9_X_21, u2_u9_X_3, u2_u9_X_30, u2_u9_X_4, u2_u9_X_45, u2_u9_X_46, 
      u2_uk_K_r0_15, u2_uk_K_r0_36, u2_uk_K_r0_49, u2_uk_K_r12_42, u2_uk_K_r14_10, u2_uk_K_r14_12, u2_uk_K_r14_18, u2_uk_K_r14_3, u2_uk_K_r14_45, 
      u2_uk_K_r14_46, u2_uk_K_r1_16, u2_uk_K_r1_21, u2_uk_K_r1_44, u2_uk_K_r2_13, u2_uk_K_r2_18, u2_uk_K_r2_25, u2_uk_K_r2_27, u2_uk_K_r2_28, 
      u2_uk_K_r2_31, u2_uk_K_r2_36, u2_uk_K_r2_49, u2_uk_K_r2_55, u2_uk_K_r3_11, u2_uk_K_r3_19, u2_uk_K_r3_4, u2_uk_K_r3_43, u2_uk_K_r3_9, 
      u2_uk_K_r4_0, u2_uk_K_r4_11, u2_uk_K_r4_17, u2_uk_K_r4_33, u2_uk_K_r4_35, u2_uk_K_r4_38, u2_uk_K_r4_4, u2_uk_K_r4_5, u2_uk_K_r4_55, 
      u2_uk_K_r5_10, u2_uk_K_r5_19, u2_uk_K_r5_41, u2_uk_K_r7_25, u2_uk_K_r7_26, u2_uk_K_r7_32, u2_uk_K_r7_39, u2_uk_K_r7_46, u2_uk_K_r8_13, 
      u2_uk_K_r8_40, u2_uk_K_r8_41, u2_uk_K_r8_43, u2_uk_K_r8_48, u2_uk_K_r9_10, u2_uk_K_r9_13, u2_uk_K_r9_19, u2_uk_K_r9_25, u2_uk_K_r9_27, 
      u2_uk_K_r9_4, u2_uk_K_r9_48, u2_uk_K_r9_55, u2_uk_n1001, u2_uk_n1008, u2_uk_n1020, u2_uk_n1024, u2_uk_n1027, u2_uk_n1028, 
      u2_uk_n1031, u2_uk_n1035, u2_uk_n1036, u2_uk_n1043, u2_uk_n1044, u2_uk_n1046, u2_uk_n1049, u2_uk_n1053, u2_uk_n1058, 
      u2_uk_n1069, u2_uk_n1074, u2_uk_n1075, u2_uk_n1076, u2_uk_n1077, u2_uk_n1079, u2_uk_n1082, u2_uk_n1083, u2_uk_n1084, 
      u2_uk_n1085, u2_uk_n1088, u2_uk_n1089, u2_uk_n1091, u2_uk_n1093, u2_uk_n1095, u2_uk_n1096, u2_uk_n11, u2_uk_n1118, 
      u2_uk_n1120, u2_uk_n1124, u2_uk_n1127, u2_uk_n1128, u2_uk_n1131, u2_uk_n1141, u2_uk_n117, u2_uk_n1189, u2_uk_n1190, 
      u2_uk_n1194, u2_uk_n1197, u2_uk_n1198, u2_uk_n1199, u2_uk_n1204, u2_uk_n1205, u2_uk_n1206, u2_uk_n1207, u2_uk_n1209, 
      u2_uk_n1212, u2_uk_n1213, u2_uk_n1216, u2_uk_n1218, u2_uk_n1221, u2_uk_n1226, u2_uk_n1227, u2_uk_n1228, u2_uk_n1230, 
      u2_uk_n1245, u2_uk_n1246, u2_uk_n1259, u2_uk_n1265, u2_uk_n1279, u2_uk_n1280, u2_uk_n1282, u2_uk_n1283, u2_uk_n1284, 
      u2_uk_n1285, u2_uk_n1287, u2_uk_n1292, u2_uk_n1293, u2_uk_n1296, u2_uk_n1298, u2_uk_n1300, u2_uk_n1301, u2_uk_n1303, 
      u2_uk_n1305, u2_uk_n1306, u2_uk_n1309, u2_uk_n1310, u2_uk_n1311, u2_uk_n1313, u2_uk_n1314, u2_uk_n1317, u2_uk_n1319, 
      u2_uk_n1322, u2_uk_n1323, u2_uk_n1325, u2_uk_n1326, u2_uk_n1329, u2_uk_n1331, u2_uk_n1333, u2_uk_n1336, u2_uk_n1339, 
      u2_uk_n1341, u2_uk_n1345, u2_uk_n1350, u2_uk_n1353, u2_uk_n1359, u2_uk_n1361, u2_uk_n1363, u2_uk_n1365, u2_uk_n1370, 
      u2_uk_n1375, u2_uk_n1381, u2_uk_n1382, u2_uk_n1403, u2_uk_n1405, u2_uk_n1408, u2_uk_n141, u2_uk_n1411, u2_uk_n1412, 
      u2_uk_n1418, u2_uk_n142, u2_uk_n1420, u2_uk_n1425, u2_uk_n1428, u2_uk_n1430, u2_uk_n1435, u2_uk_n1438, u2_uk_n1439, 
      u2_uk_n1445, u2_uk_n1446, u2_uk_n1447, u2_uk_n1453, u2_uk_n1454, u2_uk_n1456, u2_uk_n1458, u2_uk_n1460, u2_uk_n1462, 
      u2_uk_n1465, u2_uk_n1466, u2_uk_n1470, u2_uk_n1475, u2_uk_n1486, u2_uk_n1488, u2_uk_n1491, u2_uk_n1493, u2_uk_n1494, 
      u2_uk_n1496, u2_uk_n1497, u2_uk_n1544, u2_uk_n1548, u2_uk_n1549, u2_uk_n1555, u2_uk_n1568, u2_uk_n1570, u2_uk_n1573, 
      u2_uk_n1580, u2_uk_n1586, u2_uk_n1590, u2_uk_n1591, u2_uk_n1592, u2_uk_n1594, u2_uk_n1599, u2_uk_n1600, u2_uk_n1602, 
      u2_uk_n1604, u2_uk_n1605, u2_uk_n1609, u2_uk_n161, u2_uk_n1610, u2_uk_n1617, u2_uk_n1624, u2_uk_n1626, u2_uk_n1629, 
      u2_uk_n1631, u2_uk_n1639, u2_uk_n1640, u2_uk_n1643, u2_uk_n1652, u2_uk_n1657, u2_uk_n1658, u2_uk_n1660, u2_uk_n1665, 
      u2_uk_n1668, u2_uk_n1673, u2_uk_n1675, u2_uk_n1677, u2_uk_n1680, u2_uk_n1683, u2_uk_n1684, u2_uk_n1688, u2_uk_n1689, 
      u2_uk_n1709, u2_uk_n1720, u2_uk_n1769, u2_uk_n1770, u2_uk_n1776, u2_uk_n1777, u2_uk_n1781, u2_uk_n1785, u2_uk_n1791, 
      u2_uk_n1792, u2_uk_n1793, u2_uk_n1797, u2_uk_n1803, u2_uk_n1807, u2_uk_n1808, u2_uk_n1809, u2_uk_n203, u2_uk_n207, 
      u2_uk_n213, u2_uk_n214, u2_uk_n222, u2_uk_n231, u2_uk_n238, u2_uk_n240, u2_uk_n251, u2_uk_n257, u2_uk_n27, 
      u2_uk_n308, u2_uk_n313, u2_uk_n319, u2_uk_n373, u2_uk_n376, u2_uk_n407, u2_uk_n408, u2_uk_n456, u2_uk_n467, 
      u2_uk_n520, u2_uk_n689, u2_uk_n692, u2_uk_n694, u2_uk_n702, u2_uk_n948, u2_uk_n954, u2_uk_n955, u2_uk_n956, 
      u2_uk_n997, u0_out1_11, u0_out1_12, u0_out1_14, u0_out1_15, u0_out1_19, u0_out1_21, u0_out1_22, u0_out1_25, 
      u0_out1_27, u0_out1_29, u0_out1_3, u0_out1_32, u0_out1_4, u0_out1_5, u0_out1_7, u0_out1_8, u0_out3_1, 
      u0_out3_10, u0_out3_11, u0_out3_12, u0_out3_14, u0_out3_15, u0_out3_19, u0_out3_20, u0_out3_21, u0_out3_22, 
      u0_out3_25, u0_out3_26, u0_out3_27, u0_out3_29, u0_out3_3, u0_out3_32, u0_out3_4, u0_out3_5, u0_out3_7, 
      u0_out3_8, u0_out6_1, u0_out6_10, u0_out6_11, u0_out6_12, u0_out6_13, u0_out6_14, u0_out6_15, u0_out6_16, 
      u0_out6_17, u0_out6_18, u0_out6_19, u0_out6_2, u0_out6_20, u0_out6_21, u0_out6_22, u0_out6_23, u0_out6_24, 
      u0_out6_25, u0_out6_26, u0_out6_27, u0_out6_28, u0_out6_29, u0_out6_3, u0_out6_30, u0_out6_31, u0_out6_32, 
      u0_out6_4, u0_out6_5, u0_out6_6, u0_out6_7, u0_out6_8, u0_out6_9, u2_out10_1, u2_out10_10, u2_out10_11, 
      u2_out10_13, u2_out10_16, u2_out10_17, u2_out10_18, u2_out10_19, u2_out10_2, u2_out10_20, u2_out10_23, u2_out10_24, 
      u2_out10_26, u2_out10_28, u2_out10_29, u2_out10_30, u2_out10_31, u2_out10_4, u2_out10_6, u2_out10_9, u2_out11_11, 
      u2_out11_13, u2_out11_14, u2_out11_18, u2_out11_19, u2_out11_2, u2_out11_25, u2_out11_28, u2_out11_29, u2_out11_3, 
      u2_out11_4, u2_out11_8, u2_out13_11, u2_out13_12, u2_out13_14, u2_out13_19, u2_out13_22, u2_out13_25, u2_out13_29, 
      u2_out13_3, u2_out13_32, u2_out13_4, u2_out13_7, u2_out13_8, u2_out15_1, u2_out15_10, u2_out15_13, u2_out15_14, 
      u2_out15_16, u2_out15_17, u2_out15_18, u2_out15_2, u2_out15_20, u2_out15_23, u2_out15_24, u2_out15_25, u2_out15_26, 
      u2_out15_28, u2_out15_3, u2_out15_30, u2_out15_31, u2_out15_6, u2_out15_8, u2_out15_9, u2_out1_11, u2_out1_12, 
      u2_out1_14, u2_out1_19, u2_out1_22, u2_out1_25, u2_out1_29, u2_out1_3, u2_out1_32, u2_out1_4, u2_out1_7, 
      u2_out1_8, u2_out2_1, u2_out2_10, u2_out2_11, u2_out2_12, u2_out2_13, u2_out2_14, u2_out2_15, u2_out2_16, 
      u2_out2_17, u2_out2_18, u2_out2_19, u2_out2_2, u2_out2_20, u2_out2_21, u2_out2_22, u2_out2_23, u2_out2_24, 
      u2_out2_25, u2_out2_26, u2_out2_27, u2_out2_28, u2_out2_29, u2_out2_3, u2_out2_30, u2_out2_31, u2_out2_32, 
      u2_out2_4, u2_out2_5, u2_out2_6, u2_out2_7, u2_out2_8, u2_out2_9, u2_out3_1, u2_out3_10, u2_out3_11, 
      u2_out3_12, u2_out3_13, u2_out3_14, u2_out3_15, u2_out3_16, u2_out3_17, u2_out3_18, u2_out3_19, u2_out3_2, 
      u2_out3_20, u2_out3_21, u2_out3_22, u2_out3_23, u2_out3_24, u2_out3_25, u2_out3_26, u2_out3_27, u2_out3_28, 
      u2_out3_29, u2_out3_3, u2_out3_30, u2_out3_31, u2_out3_32, u2_out3_4, u2_out3_5, u2_out3_6, u2_out3_7, 
      u2_out3_8, u2_out3_9, u2_out4_1, u2_out4_10, u2_out4_11, u2_out4_12, u2_out4_13, u2_out4_14, u2_out4_15, 
      u2_out4_16, u2_out4_17, u2_out4_18, u2_out4_19, u2_out4_2, u2_out4_20, u2_out4_21, u2_out4_22, u2_out4_23, 
      u2_out4_24, u2_out4_25, u2_out4_26, u2_out4_27, u2_out4_28, u2_out4_29, u2_out4_3, u2_out4_30, u2_out4_31, 
      u2_out4_32, u2_out4_4, u2_out4_5, u2_out4_6, u2_out4_7, u2_out4_8, u2_out4_9, u2_out5_1, u2_out5_10, 
      u2_out5_11, u2_out5_12, u2_out5_13, u2_out5_14, u2_out5_15, u2_out5_16, u2_out5_17, u2_out5_18, u2_out5_19, 
      u2_out5_2, u2_out5_20, u2_out5_21, u2_out5_22, u2_out5_23, u2_out5_24, u2_out5_25, u2_out5_26, u2_out5_27, 
      u2_out5_28, u2_out5_29, u2_out5_3, u2_out5_30, u2_out5_31, u2_out5_32, u2_out5_4, u2_out5_5, u2_out5_6, 
      u2_out5_7, u2_out5_8, u2_out5_9, u2_out6_1, u2_out6_10, u2_out6_11, u2_out6_12, u2_out6_13, u2_out6_14, 
      u2_out6_15, u2_out6_16, u2_out6_17, u2_out6_18, u2_out6_19, u2_out6_2, u2_out6_20, u2_out6_21, u2_out6_22, 
      u2_out6_23, u2_out6_24, u2_out6_25, u2_out6_26, u2_out6_27, u2_out6_28, u2_out6_29, u2_out6_3, u2_out6_30, 
      u2_out6_31, u2_out6_32, u2_out6_4, u2_out6_5, u2_out6_6, u2_out6_7, u2_out6_8, u2_out6_9, u2_out8_1, 
      u2_out8_10, u2_out8_13, u2_out8_14, u2_out8_16, u2_out8_18, u2_out8_2, u2_out8_20, u2_out8_24, u2_out8_25, 
      u2_out8_26, u2_out8_28, u2_out8_3, u2_out8_30, u2_out8_6, u2_out8_8, u2_out9_1, u2_out9_10, u2_out9_13, 
      u2_out9_14, u2_out9_15, u2_out9_16, u2_out9_17, u2_out9_18, u2_out9_2, u2_out9_20, u2_out9_21, u2_out9_23, 
      u2_out9_24, u2_out9_25, u2_out9_26, u2_out9_27, u2_out9_28, u2_out9_3, u2_out9_30, u2_out9_31, u2_out9_5, 
      u2_out9_6, u2_out9_8, u2_out9_9, u2_uk_n10, u2_uk_n100, u2_uk_n102, u2_uk_n109, u2_uk_n110, u2_uk_n118, 
      u2_uk_n128, u2_uk_n129, u2_uk_n145, u2_uk_n146, u2_uk_n147, u2_uk_n148, u2_uk_n155, u2_uk_n162, u2_uk_n163, 
      u2_uk_n164, u2_uk_n17, u2_uk_n182, u2_uk_n187, u2_uk_n188, u2_uk_n191, u2_uk_n202, u2_uk_n208, u2_uk_n209, 
      u2_uk_n217, u2_uk_n220, u2_uk_n223, u2_uk_n230, u2_uk_n31, u2_uk_n60, u2_uk_n63, u2_uk_n83, u2_uk_n92, 
      u2_uk_n93, u2_uk_n94, u2_uk_n99 );
  des_des_die_4 u4 ( n116, u0_FP_33, u0_FP_48, u0_FP_49, u0_FP_50, u0_FP_51, u0_FP_52, u0_FP_53, u0_FP_54, 
      u0_FP_55, u0_FP_56, u0_FP_57, u0_FP_58, u0_FP_59, u0_FP_60, u0_FP_61, u0_FP_62, u0_FP_63, 
      u0_FP_64, u0_K10_10, u0_K10_13, u0_K10_14, u0_K10_18, u0_K10_19, u0_K10_20, u0_K12_19, u0_K12_22, 
      u0_K12_34, u0_K12_35, u0_K12_36, u0_K12_39, u0_K12_40, u0_K12_48, u0_K12_7, u0_K12_9, u0_K14_10, 
      u0_K14_12, u0_K14_13, u0_K14_14, u0_K14_15, u0_K14_18, u0_K14_4, u0_K14_9, u0_K16_26, u0_K16_38, 
      u0_K5_13, u0_K5_14, u0_K5_15, u0_K5_16, u0_K5_18, u0_K5_19, u0_K5_23, u0_K5_24, u0_K5_26, 
      u0_K5_28, u0_K5_9, u0_K9_14, u0_K9_15, u0_K9_32, u0_K9_39, u0_K9_4, u0_K9_40, u0_K9_45, 
      u0_K9_6, u0_L10_1, u0_L10_10, u0_L10_11, u0_L10_12, u0_L10_13, u0_L10_14, u0_L10_15, u0_L10_16, 
      u0_L10_17, u0_L10_18, u0_L10_19, u0_L10_2, u0_L10_20, u0_L10_21, u0_L10_22, u0_L10_23, u0_L10_24, 
      u0_L10_25, u0_L10_26, u0_L10_27, u0_L10_28, u0_L10_29, u0_L10_3, u0_L10_30, u0_L10_31, u0_L10_32, 
      u0_L10_4, u0_L10_5, u0_L10_6, u0_L10_7, u0_L10_8, u0_L10_9, u0_L12_13, u0_L12_16, u0_L12_17, 
      u0_L12_18, u0_L12_2, u0_L12_23, u0_L12_24, u0_L12_28, u0_L12_30, u0_L12_31, u0_L12_6, u0_L12_9, 
      u0_L14_11, u0_L14_12, u0_L14_14, u0_L14_15, u0_L14_19, u0_L14_21, u0_L14_22, u0_L14_25, u0_L14_27, 
      u0_L14_29, u0_L14_3, u0_L14_32, u0_L14_4, u0_L14_5, u0_L14_7, u0_L14_8, u0_L3_1, u0_L3_10, 
      u0_L3_13, u0_L3_14, u0_L3_16, u0_L3_18, u0_L3_2, u0_L3_20, u0_L3_24, u0_L3_25, u0_L3_26, 
      u0_L3_28, u0_L3_3, u0_L3_30, u0_L3_6, u0_L3_8, u0_L7_1, u0_L7_10, u0_L7_11, u0_L7_12, 
      u0_L7_13, u0_L7_14, u0_L7_15, u0_L7_16, u0_L7_17, u0_L7_18, u0_L7_19, u0_L7_2, u0_L7_20, 
      u0_L7_21, u0_L7_22, u0_L7_23, u0_L7_24, u0_L7_25, u0_L7_26, u0_L7_27, u0_L7_28, u0_L7_29, 
      u0_L7_3, u0_L7_30, u0_L7_31, u0_L7_32, u0_L7_4, u0_L7_5, u0_L7_6, u0_L7_7, u0_L7_8, 
      u0_L7_9, u0_L8_1, u0_L8_10, u0_L8_13, u0_L8_16, u0_L8_18, u0_L8_2, u0_L8_20, u0_L8_24, 
      u0_L8_26, u0_L8_28, u0_L8_30, u0_L8_6, u0_R10_1, u0_R10_10, u0_R10_11, u0_R10_12, u0_R10_13, 
      u0_R10_14, u0_R10_15, u0_R10_16, u0_R10_17, u0_R10_18, u0_R10_19, u0_R10_2, u0_R10_20, u0_R10_21, 
      u0_R10_22, u0_R10_23, u0_R10_24, u0_R10_25, u0_R10_26, u0_R10_27, u0_R10_28, u0_R10_29, u0_R10_3, 
      u0_R10_30, u0_R10_31, u0_R10_32, u0_R10_4, u0_R10_5, u0_R10_6, u0_R10_7, u0_R10_8, u0_R10_9, 
      u0_R12_1, u0_R12_10, u0_R12_11, u0_R12_12, u0_R12_13, u0_R12_2, u0_R12_3, u0_R12_32, u0_R12_4, 
      u0_R12_5, u0_R12_6, u0_R12_7, u0_R12_8, u0_R12_9, u0_R3_10, u0_R3_11, u0_R3_12, u0_R3_13, 
      u0_R3_14, u0_R3_15, u0_R3_16, u0_R3_17, u0_R3_18, u0_R3_19, u0_R3_20, u0_R3_21, u0_R3_4, 
      u0_R3_5, u0_R3_6, u0_R3_7, u0_R3_8, u0_R3_9, u0_R7_1, u0_R7_10, u0_R7_11, u0_R7_12, 
      u0_R7_13, u0_R7_14, u0_R7_15, u0_R7_16, u0_R7_17, u0_R7_18, u0_R7_19, u0_R7_2, u0_R7_20, 
      u0_R7_21, u0_R7_22, u0_R7_23, u0_R7_24, u0_R7_25, u0_R7_26, u0_R7_27, u0_R7_28, u0_R7_29, 
      u0_R7_3, u0_R7_30, u0_R7_31, u0_R7_32, u0_R7_4, u0_R7_5, u0_R7_6, u0_R7_7, u0_R7_8, 
      u0_R7_9, u0_R8_10, u0_R8_11, u0_R8_12, u0_R8_13, u0_R8_14, u0_R8_15, u0_R8_16, u0_R8_17, 
      u0_R8_4, u0_R8_5, u0_R8_6, u0_R8_7, u0_R8_8, u0_R8_9, u0_uk_K_r10_10, u0_uk_K_r10_14, u0_uk_K_r10_18, 
      u0_uk_K_r10_23, u0_uk_K_r10_25, u0_uk_K_r10_27, u0_uk_K_r10_28, u0_uk_K_r10_32, u0_uk_K_r10_34, u0_uk_K_r10_37, u0_uk_K_r10_39, u0_uk_K_r10_41, 
      u0_uk_K_r10_42, u0_uk_K_r10_43, u0_uk_K_r10_44, u0_uk_K_r10_47, u0_uk_K_r10_48, u0_uk_K_r10_9, u0_uk_K_r12_10, u0_uk_K_r12_47, u0_uk_K_r14_15, 
      u0_uk_K_r14_16, u0_uk_K_r14_2, u0_uk_K_r14_43, u0_uk_K_r14_45, u0_uk_K_r14_50, u0_uk_K_r14_8, u0_uk_K_r14_9, u0_uk_K_r3_11, u0_uk_K_r3_19, 
      u0_uk_K_r3_24, u0_uk_K_r3_35, u0_uk_K_r3_47, u0_uk_K_r7_0, u0_uk_K_r7_1, u0_uk_K_r7_13, u0_uk_K_r7_15, u0_uk_K_r7_2, u0_uk_K_r7_20, 
      u0_uk_K_r7_22, u0_uk_K_r7_23, u0_uk_K_r7_24, u0_uk_K_r7_25, u0_uk_K_r7_26, u0_uk_K_r7_27, u0_uk_K_r7_30, u0_uk_K_r7_32, u0_uk_K_r7_39, 
      u0_uk_K_r7_48, u0_uk_K_r7_55, u0_uk_K_r7_6, u0_uk_K_r7_8, u0_uk_K_r7_9, u0_uk_K_r8_13, u0_uk_K_r8_17, u0_uk_K_r8_27, u0_uk_K_r8_32, 
      u0_uk_K_r8_40, u0_uk_n1019, u0_uk_n102, u0_uk_n1020, u0_uk_n1024, u0_uk_n109, u0_uk_n11, u0_uk_n110, u0_uk_n118, 
      u0_uk_n136, u0_uk_n137, u0_uk_n139, u0_uk_n140, u0_uk_n141, u0_uk_n142, u0_uk_n143, u0_uk_n144, u0_uk_n145, 
      u0_uk_n147, u0_uk_n149, u0_uk_n150, u0_uk_n151, u0_uk_n152, u0_uk_n153, u0_uk_n154, u0_uk_n155, u0_uk_n156, 
      u0_uk_n157, u0_uk_n159, u0_uk_n162, u0_uk_n163, u0_uk_n164, u0_uk_n165, u0_uk_n166, u0_uk_n167, u0_uk_n168, 
      u0_uk_n169, u0_uk_n17, u0_uk_n170, u0_uk_n171, u0_uk_n172, u0_uk_n173, u0_uk_n174, u0_uk_n175, u0_uk_n176, 
      u0_uk_n177, u0_uk_n178, u0_uk_n179, u0_uk_n180, u0_uk_n188, u0_uk_n191, u0_uk_n202, u0_uk_n207, u0_uk_n209, 
      u0_uk_n213, u0_uk_n217, u0_uk_n220, u0_uk_n222, u0_uk_n223, u0_uk_n228, u0_uk_n229, u0_uk_n230, u0_uk_n231, 
      u0_uk_n234, u0_uk_n238, u0_uk_n242, u0_uk_n245, u0_uk_n250, u0_uk_n252, u0_uk_n253, u0_uk_n254, u0_uk_n257, 
      u0_uk_n259, u0_uk_n262, u0_uk_n266, u0_uk_n267, u0_uk_n268, u0_uk_n272, u0_uk_n273, u0_uk_n274, u0_uk_n275, 
      u0_uk_n276, u0_uk_n278, u0_uk_n280, u0_uk_n281, u0_uk_n282, u0_uk_n283, u0_uk_n285, u0_uk_n288, u0_uk_n289, 
      u0_uk_n290, u0_uk_n293, u0_uk_n296, u0_uk_n300, u0_uk_n303, u0_uk_n304, u0_uk_n307, u0_uk_n309, u0_uk_n31, 
      u0_uk_n310, u0_uk_n311, u0_uk_n314, u0_uk_n315, u0_uk_n316, u0_uk_n451, u0_uk_n453, u0_uk_n459, u0_uk_n46, 
      u0_uk_n462, u0_uk_n463, u0_uk_n464, u0_uk_n465, u0_uk_n473, u0_uk_n475, u0_uk_n479, u0_uk_n480, u0_uk_n481, 
      u0_uk_n483, u0_uk_n484, u0_uk_n485, u0_uk_n489, u0_uk_n53, u0_uk_n54, u0_uk_n57, u0_uk_n60, u0_uk_n62, 
      u0_uk_n63, u0_uk_n632, u0_uk_n633, u0_uk_n635, u0_uk_n638, u0_uk_n64, u0_uk_n641, u0_uk_n642, u0_uk_n643, 
      u0_uk_n647, u0_uk_n648, u0_uk_n649, u0_uk_n650, u0_uk_n655, u0_uk_n657, u0_uk_n658, u0_uk_n663, u0_uk_n666, 
      u0_uk_n669, u0_uk_n670, u0_uk_n69, u0_uk_n719, u0_uk_n72, u0_uk_n720, u0_uk_n725, u0_uk_n726, u0_uk_n728, 
      u0_uk_n731, u0_uk_n732, u0_uk_n735, u0_uk_n736, u0_uk_n739, u0_uk_n740, u0_uk_n75, u0_uk_n78, u0_uk_n80, 
      u0_uk_n813, u0_uk_n815, u0_uk_n83, u0_uk_n84, u0_uk_n85, u0_uk_n87, u0_uk_n897, u0_uk_n898, u0_uk_n904, 
      u0_uk_n92, u0_uk_n93, u0_uk_n94, u0_uk_n963, u0_uk_n981, u1_FP_33, u1_FP_36, u1_FP_40, u1_FP_41, 
      u1_FP_44, u1_FP_45, u1_FP_48, u1_FP_52, u1_FP_53, u1_FP_54, u1_FP_55, u1_FP_56, u1_FP_57, 
      u1_FP_60, u1_FP_61, u1_FP_62, u1_FP_63, u1_FP_64, u1_R0_1, u1_R0_10, u1_R0_11, u1_R0_12, 
      u1_R0_13, u1_R0_16, u1_R0_17, u1_R0_20, u1_R0_21, u1_R0_24, u1_R0_25, u1_R0_28, u1_R0_29, 
      u1_R0_4, u1_R0_5, u1_R0_6, u1_R0_7, u1_R0_8, u1_R0_9, u1_R10_1, u1_R10_12, u1_R10_13, 
      u1_R10_14, u1_R10_15, u1_R10_16, u1_R10_17, u1_R10_18, u1_R10_19, u1_R10_20, u1_R10_21, u1_R10_24, 
      u1_R10_29, u1_R10_32, u1_R10_5, u1_R11_1, u1_R11_10, u1_R11_11, u1_R11_12, u1_R11_13, u1_R11_16, 
      u1_R11_20, u1_R11_21, u1_R11_28, u1_R11_29, u1_R11_4, u1_R11_8, u1_R11_9, u1_R12_1, u1_R12_12, 
      u1_R12_13, u1_R12_16, u1_R12_17, u1_R12_21, u1_R12_24, u1_R12_25, u1_R12_26, u1_R12_27, u1_R12_28, 
      u1_R12_29, u1_R12_30, u1_R12_31, u1_R12_32, u1_R12_4, u1_R12_5, u1_R12_8, u1_R13_1, u1_R13_16, 
      u1_R13_17, u1_R13_20, u1_R13_21, u1_R13_24, u1_R13_25, u1_R13_26, u1_R13_27, u1_R13_28, u1_R13_29, 
      u1_R13_32, u1_R13_8, u1_R1_1, u1_R1_12, u1_R1_13, u1_R1_14, u1_R1_15, u1_R1_16, u1_R1_17, 
      u1_R1_20, u1_R1_21, u1_R1_22, u1_R1_23, u1_R1_24, u1_R1_25, u1_R1_28, u1_R1_29, u1_R1_30, 
      u1_R1_31, u1_R1_32, u1_R1_5, u1_R1_8, u1_R1_9, u1_R2_1, u1_R2_2, u1_R2_20, u1_R2_21, 
      u1_R2_22, u1_R2_23, u1_R2_24, u1_R2_25, u1_R2_28, u1_R2_29, u1_R2_3, u1_R2_32, u1_R2_4, 
      u1_R2_5, u1_R2_8, u1_R2_9, u1_R3_1, u1_R3_12, u1_R3_2, u1_R3_29, u1_R3_3, u1_R3_32, 
      u1_R3_4, u1_R3_5, u1_R3_8, u1_R3_9, u1_R4_10, u1_R4_11, u1_R4_12, u1_R4_13, u1_R4_16, 
      u1_R4_17, u1_R4_18, u1_R4_19, u1_R4_20, u1_R4_21, u1_R4_4, u1_R4_8, u1_R4_9, u1_R5_1, 
      u1_R5_24, u1_R5_25, u1_R5_29, u1_R5_32, u1_R6_1, u1_R6_12, u1_R6_17, u1_R6_20, u1_R6_21, 
      u1_R6_22, u1_R6_23, u1_R6_24, u1_R6_25, u1_R6_26, u1_R6_27, u1_R6_28, u1_R6_29, u1_R6_32, 
      u1_R7_1, u1_R7_20, u1_R7_21, u1_R7_28, u1_R7_29, u1_R7_30, u1_R7_31, u1_R7_32, u1_R7_4, 
      u1_R7_5, u1_R7_9, u1_R8_1, u1_R8_16, u1_R8_17, u1_R8_2, u1_R8_20, u1_R8_21, u1_R8_24, 
      u1_R8_25, u1_R8_26, u1_R8_27, u1_R8_28, u1_R8_29, u1_R8_3, u1_R8_32, u1_R8_4, u1_R8_5, 
      u1_R8_8, u1_R8_9, u1_R9_1, u1_R9_12, u1_R9_13, u1_R9_14, u1_R9_15, u1_R9_16, u1_R9_17, 
      u1_R9_18, u1_R9_19, u1_R9_20, u1_R9_21, u1_R9_22, u1_R9_23, u1_R9_24, u1_R9_25, u1_R9_26, 
      u1_R9_27, u1_R9_28, u1_R9_29, u1_R9_4, u1_desIn_r_1, u1_desIn_r_11, u1_desIn_r_19, u1_desIn_r_27, u1_desIn_r_29, 
      u1_desIn_r_3, u1_desIn_r_31, u1_desIn_r_35, u1_desIn_r_37, u1_desIn_r_39, u1_desIn_r_57, u1_desIn_r_59, u1_desIn_r_61, u1_desIn_r_63, 
      u1_desIn_r_7, u1_key_r_0, u1_key_r_1, u1_key_r_10, u1_key_r_11, u1_key_r_12, u1_key_r_13, u1_key_r_14, u1_key_r_15, 
      u1_key_r_16, u1_key_r_17, u1_key_r_18, u1_key_r_19, u1_key_r_2, u1_key_r_20, u1_key_r_21, u1_key_r_22, u1_key_r_23, 
      u1_key_r_24, u1_key_r_25, u1_key_r_26, u1_key_r_27, u1_key_r_28, u1_key_r_29, u1_key_r_3, u1_key_r_30, u1_key_r_31, 
      u1_key_r_32, u1_key_r_33, u1_key_r_34, u1_key_r_35, u1_key_r_36, u1_key_r_37, u1_key_r_38, u1_key_r_39, u1_key_r_4, 
      u1_key_r_40, u1_key_r_41, u1_key_r_42, u1_key_r_43, u1_key_r_44, u1_key_r_45, u1_key_r_46, u1_key_r_47, u1_key_r_48, 
      u1_key_r_49, u1_key_r_5, u1_key_r_50, u1_key_r_51, u1_key_r_52, u1_key_r_53, u1_key_r_54, u1_key_r_55, u1_key_r_6, 
      u1_key_r_7, u1_key_r_8, u1_key_r_9, u1_uk_K_r0_11, u1_uk_K_r0_13, u1_uk_K_r0_15, u1_uk_K_r0_17, u1_uk_K_r0_19, u1_uk_K_r0_2, 
      u1_uk_K_r0_22, u1_uk_K_r0_25, u1_uk_K_r0_28, u1_uk_K_r0_31, u1_uk_K_r0_32, u1_uk_K_r0_34, u1_uk_K_r0_36, u1_uk_K_r0_47, u1_uk_K_r0_49, 
      u1_uk_K_r0_52, u1_uk_K_r0_55, u1_uk_K_r0_7, u1_uk_K_r10_10, u1_uk_K_r10_11, u1_uk_K_r10_14, u1_uk_K_r10_16, u1_uk_K_r10_18, u1_uk_K_r10_19, 
      u1_uk_K_r10_23, u1_uk_K_r10_25, u1_uk_K_r10_27, u1_uk_K_r10_28, u1_uk_K_r10_32, u1_uk_K_r10_34, u1_uk_K_r10_37, u1_uk_K_r10_39, u1_uk_K_r10_4, 
      u1_uk_K_r10_41, u1_uk_K_r10_42, u1_uk_K_r10_43, u1_uk_K_r10_44, u1_uk_K_r10_47, u1_uk_K_r10_48, u1_uk_K_r10_49, u1_uk_K_r10_52, u1_uk_K_r10_9, 
      u1_uk_K_r11_10, u1_uk_K_r11_11, u1_uk_K_r11_17, u1_uk_K_r11_19, u1_uk_K_r11_20, u1_uk_K_r11_21, u1_uk_K_r11_24, u1_uk_K_r11_25, u1_uk_K_r11_26, 
      u1_uk_K_r11_27, u1_uk_K_r11_28, u1_uk_K_r11_29, u1_uk_K_r11_33, u1_uk_K_r11_34, u1_uk_K_r11_39, u1_uk_K_r11_4, u1_uk_K_r11_46, u1_uk_K_r11_47, 
      u1_uk_K_r11_48, u1_uk_K_r11_5, u1_uk_K_r11_53, u1_uk_K_r11_54, u1_uk_K_r11_6, u1_uk_K_r11_7, u1_uk_K_r11_8, u1_uk_K_r12_1, u1_uk_K_r12_10, 
      u1_uk_K_r12_15, u1_uk_K_r12_16, u1_uk_K_r12_18, u1_uk_K_r12_21, u1_uk_K_r12_22, u1_uk_K_r12_25, u1_uk_K_r12_30, u1_uk_K_r12_33, u1_uk_K_r12_36, 
      u1_uk_K_r12_41, u1_uk_K_r12_42, u1_uk_K_r12_44, u1_uk_K_r12_47, u1_uk_K_r12_7, u1_uk_K_r13_0, u1_uk_K_r13_13, u1_uk_K_r13_17, u1_uk_K_r13_19, 
      u1_uk_K_r13_2, u1_uk_K_r13_22, u1_uk_K_r13_23, u1_uk_K_r13_25, u1_uk_K_r13_31, u1_uk_K_r13_32, u1_uk_K_r13_35, u1_uk_K_r13_36, u1_uk_K_r13_38, 
      u1_uk_K_r13_4, u1_uk_K_r13_44, u1_uk_K_r13_55, u1_uk_K_r14_10, u1_uk_K_r14_11, u1_uk_K_r14_12, u1_uk_K_r14_15, u1_uk_K_r14_16, u1_uk_K_r14_18, 
      u1_uk_K_r14_2, u1_uk_K_r14_23, u1_uk_K_r14_3, u1_uk_K_r14_38, u1_uk_K_r14_39, u1_uk_K_r14_42, u1_uk_K_r14_43, u1_uk_K_r14_45, u1_uk_K_r14_46, 
      u1_uk_K_r14_5, u1_uk_K_r14_50, u1_uk_K_r14_8, u1_uk_K_r14_9, u1_uk_K_r1_10, u1_uk_K_r1_15, u1_uk_K_r1_16, u1_uk_K_r1_17, u1_uk_K_r1_18, 
      u1_uk_K_r1_21, u1_uk_K_r1_22, u1_uk_K_r1_33, u1_uk_K_r1_36, u1_uk_K_r1_41, u1_uk_K_r1_42, u1_uk_K_r1_44, u1_uk_K_r1_47, u1_uk_K_r1_6, 
      u1_uk_K_r1_7, u1_uk_K_r2_13, u1_uk_K_r2_16, u1_uk_K_r2_18, u1_uk_K_r2_20, u1_uk_K_r2_21, u1_uk_K_r2_24, u1_uk_K_r2_25, u1_uk_K_r2_26, 
      u1_uk_K_r2_27, u1_uk_K_r2_28, u1_uk_K_r2_29, u1_uk_K_r2_31, u1_uk_K_r2_33, u1_uk_K_r2_36, u1_uk_K_r2_4, u1_uk_K_r2_41, u1_uk_K_r2_46, 
      u1_uk_K_r2_47, u1_uk_K_r2_49, u1_uk_K_r2_50, u1_uk_K_r2_53, u1_uk_K_r2_55, u1_uk_K_r2_6, u1_uk_K_r2_7, u1_uk_K_r3_10, u1_uk_K_r3_11, 
      u1_uk_K_r3_14, u1_uk_K_r3_15, u1_uk_K_r3_16, u1_uk_K_r3_19, u1_uk_K_r3_24, u1_uk_K_r3_29, u1_uk_K_r3_33, u1_uk_K_r3_34, u1_uk_K_r3_35, 
      u1_uk_K_r3_38, u1_uk_K_r3_4, u1_uk_K_r3_43, u1_uk_K_r3_44, u1_uk_K_r3_47, u1_uk_K_r3_51, u1_uk_K_r3_52, u1_uk_K_r3_9, u1_uk_K_r4_0, 
      u1_uk_K_r4_11, u1_uk_K_r4_17, u1_uk_K_r4_18, u1_uk_K_r4_23, u1_uk_K_r4_27, u1_uk_K_r4_3, u1_uk_K_r4_31, u1_uk_K_r4_33, u1_uk_K_r4_35, 
      u1_uk_K_r4_38, u1_uk_K_r4_4, u1_uk_K_r4_41, u1_uk_K_r4_47, u1_uk_K_r4_48, u1_uk_K_r4_49, u1_uk_K_r4_5, u1_uk_K_r4_54, u1_uk_K_r4_55, 
      u1_uk_K_r5_0, u1_uk_K_r5_1, u1_uk_K_r5_10, u1_uk_K_r5_13, u1_uk_K_r5_16, u1_uk_K_r5_17, u1_uk_K_r5_18, u1_uk_K_r5_19, u1_uk_K_r5_21, 
      u1_uk_K_r5_23, u1_uk_K_r5_26, u1_uk_K_r5_31, u1_uk_K_r5_32, u1_uk_K_r5_35, u1_uk_K_r5_36, u1_uk_K_r5_37, u1_uk_K_r5_39, u1_uk_K_r5_4, 
      u1_uk_K_r5_40, u1_uk_K_r5_41, u1_uk_K_r5_43, u1_uk_K_r5_48, u1_uk_K_r5_5, u1_uk_K_r5_51, u1_uk_K_r5_53, u1_uk_K_r5_7, u1_uk_K_r5_8, 
      u1_uk_K_r6_0, u1_uk_K_r6_10, u1_uk_K_r6_14, u1_uk_K_r6_17, u1_uk_K_r6_19, u1_uk_K_r6_21, u1_uk_K_r6_22, u1_uk_K_r6_26, u1_uk_K_r6_27, 
      u1_uk_K_r6_28, u1_uk_K_r6_29, u1_uk_K_r6_3, u1_uk_K_r6_30, u1_uk_K_r6_31, u1_uk_K_r6_34, u1_uk_K_r6_35, u1_uk_K_r6_37, u1_uk_K_r6_46, 
      u1_uk_K_r6_51, u1_uk_K_r6_53, u1_uk_K_r6_55, u1_uk_K_r6_7, u1_uk_K_r7_0, u1_uk_K_r7_1, u1_uk_K_r7_13, u1_uk_K_r7_15, u1_uk_K_r7_16, 
      u1_uk_K_r7_2, u1_uk_K_r7_20, u1_uk_K_r7_22, u1_uk_K_r7_23, u1_uk_K_r7_24, u1_uk_K_r7_25, u1_uk_K_r7_26, u1_uk_K_r7_27, u1_uk_K_r7_29, 
      u1_uk_K_r7_30, u1_uk_K_r7_31, u1_uk_K_r7_32, u1_uk_K_r7_34, u1_uk_K_r7_37, u1_uk_K_r7_39, u1_uk_K_r7_41, u1_uk_K_r7_46, u1_uk_K_r7_48, 
      u1_uk_K_r7_5, u1_uk_K_r7_53, u1_uk_K_r7_55, u1_uk_K_r7_6, u1_uk_K_r7_7, u1_uk_K_r7_8, u1_uk_K_r7_9, u1_uk_K_r8_10, u1_uk_K_r8_13, 
      u1_uk_K_r8_16, u1_uk_K_r8_17, u1_uk_K_r8_19, u1_uk_K_r8_2, u1_uk_K_r8_21, u1_uk_K_r8_22, u1_uk_K_r8_27, u1_uk_K_r8_28, u1_uk_K_r8_32, 
      u1_uk_K_r8_37, u1_uk_K_r8_39, u1_uk_K_r8_40, u1_uk_K_r8_41, u1_uk_K_r8_42, u1_uk_K_r8_43, u1_uk_K_r8_44, u1_uk_K_r8_48, u1_uk_K_r8_5, 
      u1_uk_K_r8_51, u1_uk_K_r8_52, u1_uk_K_r8_8, u1_uk_K_r9_0, u1_uk_K_r9_1, u1_uk_K_r9_10, u1_uk_K_r9_12, u1_uk_K_r9_13, u1_uk_K_r9_15, 
      u1_uk_K_r9_18, u1_uk_K_r9_19, u1_uk_K_r9_22, u1_uk_K_r9_23, u1_uk_K_r9_25, u1_uk_K_r9_27, u1_uk_K_r9_30, u1_uk_K_r9_31, u1_uk_K_r9_33, 
      u1_uk_K_r9_35, u1_uk_K_r9_38, u1_uk_K_r9_4, u1_uk_K_r9_45, u1_uk_K_r9_48, u1_uk_K_r9_49, u1_uk_K_r9_5, u1_uk_K_r9_54, u1_uk_K_r9_55, 
      u1_uk_K_r9_6, u1_uk_K_r9_7, u1_uk_K_r9_9, u1_uk_n1218, u1_uk_n1219, u1_uk_n1220, u1_uk_n1221, u1_uk_n1222, u1_uk_n1224, 
      u1_uk_n1225, u1_uk_n1227, u1_uk_n1228, u1_uk_n1229, u1_uk_n1230, u1_uk_n1231, u1_uk_n1233, u1_uk_n1234, u1_uk_n1235, 
      u1_uk_n1236, u1_uk_n1237, u1_uk_n1238, u1_uk_n1239, u1_uk_n1240, u1_uk_n1241, u1_uk_n1242, u1_uk_n1243, u1_uk_n1244, 
      u1_uk_n1245, u1_uk_n1246, u1_uk_n1247, u1_uk_n1248, u1_uk_n1249, u1_uk_n1250, u1_uk_n1251, u1_uk_n1252, u1_uk_n1253, 
      u1_uk_n1255, u1_uk_n1256, u1_uk_n1257, u1_uk_n1258, u1_uk_n1259, u1_uk_n1260, u1_uk_n1261, u1_uk_n1262, u1_uk_n1263, 
      u1_uk_n1264, u1_uk_n1265, u1_uk_n1266, u1_uk_n1267, u1_uk_n1268, u1_uk_n1269, u1_uk_n1270, u1_uk_n1271, u1_uk_n1272, 
      u1_uk_n1273, u1_uk_n1274, u1_uk_n1275, u1_uk_n1276, u1_uk_n1277, u1_uk_n1278, u1_uk_n1279, u1_uk_n1281, u1_uk_n1282, 
      u1_uk_n1284, u1_uk_n1286, u1_uk_n1288, u1_uk_n1289, u1_uk_n1290, u1_uk_n1291, u1_uk_n1292, u1_uk_n1293, u1_uk_n1294, 
      u1_uk_n1295, u1_uk_n1296, u1_uk_n1297, u1_uk_n1299, u1_uk_n1300, u1_uk_n1303, u1_uk_n1304, u1_uk_n1305, u1_uk_n1307, 
      u1_uk_n1308, u1_uk_n1309, u1_uk_n1310, u1_uk_n1311, u1_uk_n1312, u1_uk_n1313, u1_uk_n1314, u1_uk_n1315, u1_uk_n1316, 
      u1_uk_n1317, u1_uk_n1318, u1_uk_n1319, u1_uk_n1320, u1_uk_n1321, u1_uk_n1322, u1_uk_n1323, u1_uk_n1324, u1_uk_n1325, 
      u1_uk_n1326, u1_uk_n1327, u1_uk_n1328, u1_uk_n1329, u1_uk_n1330, u1_uk_n1331, u1_uk_n1332, u1_uk_n1333, u1_uk_n1334, 
      u1_uk_n1335, u1_uk_n1336, u1_uk_n1338, u1_uk_n1339, u1_uk_n1340, u1_uk_n1341, u1_uk_n1342, u1_uk_n1343, u1_uk_n1344, 
      u1_uk_n1345, u1_uk_n1346, u1_uk_n1347, u1_uk_n1348, u1_uk_n1349, u1_uk_n1350, u1_uk_n1351, u1_uk_n1352, u1_uk_n1353, 
      u1_uk_n1354, u1_uk_n1355, u1_uk_n1356, u1_uk_n1357, u1_uk_n1358, u1_uk_n1359, u1_uk_n1360, u1_uk_n1361, u1_uk_n1363, 
      u1_uk_n1365, u1_uk_n1366, u1_uk_n1367, u1_uk_n1369, u1_uk_n1371, u1_uk_n1372, u1_uk_n1374, u1_uk_n1375, u1_uk_n1376, 
      u1_uk_n1377, u1_uk_n1378, u1_uk_n1380, u1_uk_n1381, u1_uk_n1382, u1_uk_n1383, u1_uk_n1386, u1_uk_n1389, u1_uk_n1390, 
      u1_uk_n1391, u1_uk_n1393, u1_uk_n1394, u1_uk_n1395, u1_uk_n1396, u1_uk_n1397, u1_uk_n1398, u1_uk_n1399, u1_uk_n1400, 
      u1_uk_n1401, u1_uk_n1402, u1_uk_n1403, u1_uk_n1404, u1_uk_n1405, u1_uk_n1406, u1_uk_n1407, u1_uk_n1408, u1_uk_n1409, 
      u1_uk_n1410, u1_uk_n1411, u1_uk_n1412, u1_uk_n1413, u1_uk_n1414, u1_uk_n1415, u1_uk_n1417, u1_uk_n1418, u1_uk_n1419, 
      u1_uk_n1422, u1_uk_n1423, u1_uk_n1424, u1_uk_n1425, u1_uk_n1426, u1_uk_n1427, u1_uk_n1429, u1_uk_n1430, u1_uk_n1431, 
      u1_uk_n1433, u1_uk_n1435, u1_uk_n1436, u1_uk_n1437, u1_uk_n1438, u1_uk_n1439, u1_uk_n1440, u1_uk_n1441, u1_uk_n1442, 
      u1_uk_n1443, u1_uk_n1444, u1_uk_n1446, u1_uk_n1447, u1_uk_n1448, u1_uk_n1449, u1_uk_n1450, u1_uk_n1452, u1_uk_n1453, 
      u1_uk_n1454, u1_uk_n1455, u1_uk_n1456, u1_uk_n1457, u1_uk_n1458, u1_uk_n1459, u1_uk_n1460, u1_uk_n1461, u1_uk_n1462, 
      u1_uk_n1463, u1_uk_n1464, u1_uk_n1465, u1_uk_n1466, u1_uk_n1468, u1_uk_n1469, u1_uk_n1470, u1_uk_n1471, u1_uk_n1472, 
      u1_uk_n1474, u1_uk_n1475, u1_uk_n1476, u1_uk_n1477, u1_uk_n1478, u1_uk_n1482, u1_uk_n1483, u1_uk_n1484, u1_uk_n1485, 
      u1_uk_n1486, u1_uk_n1487, u1_uk_n1488, u1_uk_n1489, u1_uk_n1490, u1_uk_n1491, u1_uk_n1492, u1_uk_n1494, u1_uk_n1495, 
      u1_uk_n1496, u1_uk_n1498, u1_uk_n1499, u1_uk_n1500, u1_uk_n1501, u1_uk_n1504, u1_uk_n1505, u1_uk_n1507, u1_uk_n1508, 
      u1_uk_n1510, u1_uk_n1514, u1_uk_n1516, u1_uk_n1517, u1_uk_n1518, u1_uk_n1520, u1_uk_n1521, u1_uk_n1523, u1_uk_n1524, 
      u1_uk_n1526, u1_uk_n1527, u1_uk_n1528, u1_uk_n1529, u1_uk_n1530, u1_uk_n1531, u1_uk_n1532, u1_uk_n1533, u1_uk_n1534, 
      u1_uk_n1536, u1_uk_n1537, u1_uk_n1538, u1_uk_n1540, u1_uk_n1541, u1_uk_n1543, u1_uk_n1544, u1_uk_n1545, u1_uk_n1547, 
      u1_uk_n1548, u1_uk_n1549, u1_uk_n1551, u1_uk_n1552, u1_uk_n1554, u1_uk_n1555, u1_uk_n1556, u1_uk_n1557, u1_uk_n1558, 
      u1_uk_n1559, u1_uk_n1560, u1_uk_n1561, u1_uk_n1562, u1_uk_n1563, u1_uk_n1564, u1_uk_n1565, u1_uk_n1566, u1_uk_n1567, 
      u1_uk_n1568, u1_uk_n1570, u1_uk_n1571, u1_uk_n1572, u1_uk_n1573, u1_uk_n1574, u1_uk_n1577, u1_uk_n1578, u1_uk_n1579, 
      u1_uk_n1581, u1_uk_n1584, u1_uk_n1585, u1_uk_n1586, u1_uk_n1588, u1_uk_n1592, u1_uk_n1593, u1_uk_n1595, u1_uk_n1598, 
      u1_uk_n1599, u1_uk_n1600, u1_uk_n1601, u1_uk_n1603, u1_uk_n1604, u1_uk_n1605, u1_uk_n1606, u1_uk_n1607, u1_uk_n1608, 
      u1_uk_n1610, u1_uk_n1612, u1_uk_n1613, u1_uk_n1614, u1_uk_n1615, u1_uk_n1616, u1_uk_n1618, u1_uk_n1619, u1_uk_n1620, 
      u1_uk_n1621, u1_uk_n1622, u1_uk_n1623, u1_uk_n1624, u1_uk_n1625, u1_uk_n1626, u1_uk_n1627, u1_uk_n1628, u1_uk_n1629, 
      u1_uk_n1630, u1_uk_n1632, u1_uk_n1633, u1_uk_n1634, u1_uk_n1635, u1_uk_n1639, u1_uk_n1640, u1_uk_n1641, u1_uk_n1642, 
      u1_uk_n1643, u1_uk_n1644, u1_uk_n1645, u1_uk_n1647, u1_uk_n1649, u1_uk_n1651, u1_uk_n1652, u1_uk_n1653, u1_uk_n1654, 
      u1_uk_n1655, u1_uk_n1656, u1_uk_n1659, u1_uk_n1660, u1_uk_n1661, u1_uk_n1662, u1_uk_n1663, u1_uk_n1664, u1_uk_n1667, 
      u1_uk_n1669, u1_uk_n1670, u1_uk_n1672, u1_uk_n1673, u1_uk_n1676, u1_uk_n1677, u1_uk_n1678, u1_uk_n1682, u1_uk_n1683, 
      u1_uk_n1684, u1_uk_n1687, u1_uk_n1688, u1_uk_n1689, u1_uk_n1690, u1_uk_n1691, u1_uk_n1692, u1_uk_n1693, u1_uk_n1694, 
      u1_uk_n1695, u1_uk_n1696, u1_uk_n1698, u1_uk_n1699, u1_uk_n1702, u1_uk_n1703, u1_uk_n1704, u1_uk_n1705, u1_uk_n1707, 
      u1_uk_n1708, u1_uk_n1709, u1_uk_n1710, u1_uk_n1711, u1_uk_n1712, u1_uk_n1713, u1_uk_n1714, u1_uk_n1715, u1_uk_n1716, 
      u1_uk_n1717, u1_uk_n1718, u1_uk_n1719, u1_uk_n1720, u1_uk_n1721, u1_uk_n1722, u1_uk_n1723, u1_uk_n1728, u1_uk_n1729, 
      u1_uk_n1730, u1_uk_n1731, u1_uk_n1732, u1_uk_n1734, u1_uk_n1735, u1_uk_n1736, u1_uk_n1737, u1_uk_n1738, u1_uk_n1739, 
      u1_uk_n1744, u1_uk_n1745, u1_uk_n1748, u1_uk_n1749, u1_uk_n1750, u1_uk_n1751, u1_uk_n1752, u1_uk_n1753, u1_uk_n1754, 
      u1_uk_n1755, u1_uk_n1756, u1_uk_n1757, u1_uk_n1758, u1_uk_n1761, u1_uk_n1762, u1_uk_n1763, u1_uk_n1764, u1_uk_n1765, 
      u1_uk_n1766, u1_uk_n1767, u1_uk_n1768, u1_uk_n1769, u1_uk_n1772, u1_uk_n1773, u1_uk_n1774, u1_uk_n1775, u1_uk_n1776, 
      u1_uk_n1777, u1_uk_n1780, u1_uk_n1781, u1_uk_n1782, u1_uk_n1783, u1_uk_n1784, u1_uk_n1785, u1_uk_n1787, u1_uk_n1790, 
      u1_uk_n1791, u1_uk_n1792, u1_uk_n1793, u1_uk_n1797, u1_uk_n1798, u1_uk_n1799, u1_uk_n1800, u1_uk_n1801, u1_uk_n1802, 
      u1_uk_n1803, u1_uk_n1804, u1_uk_n1806, u1_uk_n1807, u1_uk_n1808, u1_uk_n1809, u1_uk_n1810, u1_uk_n1811, u1_uk_n1812, 
      u1_uk_n1813, u1_uk_n1814, u1_uk_n1815, u1_uk_n1816, u1_uk_n1817, u1_uk_n1818, u1_uk_n1819, u1_uk_n1820, u1_uk_n1821, 
      u1_uk_n1822, u1_uk_n1823, u1_uk_n1824, u1_uk_n1826, u1_uk_n1827, u1_uk_n1829, u1_uk_n1830, u1_uk_n1831, u1_uk_n1832, 
      u1_uk_n1833, u1_uk_n1834, u1_uk_n1835, u1_uk_n1836, u1_uk_n1837, u1_uk_n1838, u1_uk_n1839, u1_uk_n1840, u1_uk_n1841, 
      u1_uk_n1842, u1_uk_n1843, u1_uk_n1844, u1_uk_n1845, u1_uk_n1846, u1_uk_n1847, u1_uk_n1848, u1_uk_n1849, u1_uk_n1850, 
      u1_uk_n1851, u1_uk_n1852, u1_uk_n1853, u1_uk_n1854, u1_uk_n1855, u1_uk_n1856, u1_uk_n1858, u1_uk_n1859, u1_uk_n1860, 
      u1_uk_n1862, u1_uk_n1863, u1_uk_n1864, u1_uk_n1865, u1_uk_n1866, u1_uk_n1867, u1_uk_n1868, u1_uk_n1869, u1_uk_n1870, 
      u1_uk_n1872, u1_uk_n1873, u1_uk_n1874, u1_uk_n1875, u1_uk_n1876, u1_uk_n1879, u1_uk_n1880, u1_uk_n1881, u1_uk_n1882, 
      u1_uk_n1883, u1_uk_n1884, u1_uk_n1885, u1_uk_n1886, u1_uk_n1887, u2_FP_33, u2_FP_52, u2_FP_53, u2_FP_54, 
      u2_FP_55, u2_FP_56, u2_FP_57, u2_FP_58, u2_FP_59, u2_FP_60, u2_FP_61, u2_FP_62, u2_FP_63, 
      u2_FP_64, u2_K11_29, u2_K11_37, u2_K11_38, u2_K11_42, u2_K11_45, u2_K11_48, u2_K12_2, u2_K12_20, 
      u2_K12_22, u2_K12_24, u2_K12_41, u2_K12_46, u2_K12_47, u2_K12_48, u2_K13_14, u2_K13_20, u2_K13_25, 
      u2_K13_26, u2_K13_3, u2_K13_31, u2_K13_32, u2_K13_34, u2_K13_37, u2_K13_40, u2_K13_42, u2_K13_44, 
      u2_K13_45, u2_K13_46, u2_K13_47, u2_K13_8, u2_K14_10, u2_K14_11, u2_K14_12, u2_K14_13, u2_K14_14, 
      u2_K14_16, u2_K14_17, u2_K14_18, u2_K14_3, u2_K14_43, u2_K14_48, u2_K14_6, u2_K14_8, u2_K15_1, 
      u2_K15_13, u2_K15_16, u2_K15_18, u2_K15_2, u2_K15_20, u2_K15_5, u2_K16_31, u2_K16_42, u2_K16_44, 
      u2_K16_47, u2_K8_26, u2_K8_31, u2_K8_41, u2_K8_42, u2_K8_45, u2_K9_3, u2_K9_32, u2_K9_36, 
      u2_K9_38, u2_K9_40, u2_K9_45, u2_K9_5, u2_L10_1, u2_L10_10, u2_L10_15, u2_L10_16, u2_L10_17, 
      u2_L10_20, u2_L10_21, u2_L10_23, u2_L10_24, u2_L10_26, u2_L10_27, u2_L10_30, u2_L10_31, u2_L10_5, 
      u2_L10_6, u2_L10_9, u2_L11_1, u2_L11_10, u2_L11_11, u2_L11_12, u2_L11_13, u2_L11_14, u2_L11_15, 
      u2_L11_16, u2_L11_17, u2_L11_18, u2_L11_19, u2_L11_2, u2_L11_20, u2_L11_21, u2_L11_22, u2_L11_23, 
      u2_L11_24, u2_L11_25, u2_L11_26, u2_L11_3, u2_L11_30, u2_L11_31, u2_L11_32, u2_L11_4, u2_L11_5, 
      u2_L11_6, u2_L11_7, u2_L11_8, u2_L11_9, u2_L12_13, u2_L12_15, u2_L12_16, u2_L12_17, u2_L12_18, 
      u2_L12_2, u2_L12_21, u2_L12_23, u2_L12_24, u2_L12_27, u2_L12_28, u2_L12_30, u2_L12_31, u2_L12_5, 
      u2_L12_6, u2_L12_9, u2_L13_13, u2_L13_16, u2_L13_18, u2_L13_2, u2_L13_24, u2_L13_28, u2_L13_30, 
      u2_L13_6, u2_L14_11, u2_L14_12, u2_L14_15, u2_L14_19, u2_L14_21, u2_L14_22, u2_L14_27, u2_L14_29, 
      u2_L14_32, u2_L14_4, u2_L14_5, u2_L14_7, u2_L6_11, u2_L6_14, u2_L6_15, u2_L6_19, u2_L6_21, 
      u2_L6_22, u2_L6_25, u2_L6_27, u2_L6_29, u2_L6_3, u2_L6_32, u2_L6_4, u2_L6_5, u2_L6_7, 
      u2_L6_8, u2_L7_11, u2_L7_12, u2_L7_15, u2_L7_17, u2_L7_19, u2_L7_21, u2_L7_22, u2_L7_23, 
      u2_L7_27, u2_L7_29, u2_L7_31, u2_L7_32, u2_L7_4, u2_L7_5, u2_L7_7, u2_L7_9, u2_L9_12, 
      u2_L9_14, u2_L9_15, u2_L9_21, u2_L9_22, u2_L9_25, u2_L9_27, u2_L9_3, u2_L9_32, u2_L9_5, 
      u2_L9_7, u2_L9_8, u2_R10_1, u2_R10_10, u2_R10_11, u2_R10_12, u2_R10_13, u2_R10_14, u2_R10_15, 
      u2_R10_16, u2_R10_17, u2_R10_2, u2_R10_28, u2_R10_29, u2_R10_3, u2_R10_30, u2_R10_31, u2_R10_32, 
      u2_R10_4, u2_R10_5, u2_R10_8, u2_R10_9, u2_R11_1, u2_R11_10, u2_R11_11, u2_R11_12, u2_R11_13, 
      u2_R11_14, u2_R11_15, u2_R11_16, u2_R11_17, u2_R11_18, u2_R11_19, u2_R11_2, u2_R11_20, u2_R11_21, 
      u2_R11_22, u2_R11_23, u2_R11_24, u2_R11_25, u2_R11_26, u2_R11_27, u2_R11_28, u2_R11_29, u2_R11_3, 
      u2_R11_30, u2_R11_31, u2_R11_32, u2_R11_4, u2_R11_5, u2_R11_6, u2_R11_7, u2_R11_8, u2_R11_9, 
      u2_R12_1, u2_R12_10, u2_R12_11, u2_R12_12, u2_R12_13, u2_R12_2, u2_R12_28, u2_R12_29, u2_R12_3, 
      u2_R12_30, u2_R12_31, u2_R12_32, u2_R12_4, u2_R12_5, u2_R12_6, u2_R12_7, u2_R12_8, u2_R12_9, 
      u2_R13_1, u2_R13_10, u2_R13_11, u2_R13_12, u2_R13_13, u2_R13_17, u2_R13_32, u2_R13_4, u2_R13_5, 
      u2_R13_6, u2_R13_7, u2_R13_8, u2_R13_9, u2_R6_1, u2_R6_16, u2_R6_17, u2_R6_18, u2_R6_19, 
      u2_R6_20, u2_R6_21, u2_R6_22, u2_R6_23, u2_R6_24, u2_R6_25, u2_R6_26, u2_R6_27, u2_R6_28, 
      u2_R6_29, u2_R6_30, u2_R6_31, u2_R6_32, u2_R7_1, u2_R7_2, u2_R7_20, u2_R7_21, u2_R7_22, 
      u2_R7_23, u2_R7_24, u2_R7_25, u2_R7_26, u2_R7_27, u2_R7_28, u2_R7_29, u2_R7_3, u2_R7_30, 
      u2_R7_31, u2_R7_32, u2_R7_4, u2_R7_5, u2_R9_1, u2_R9_16, u2_R9_17, u2_R9_18, u2_R9_19, 
      u2_R9_20, u2_R9_21, u2_R9_24, u2_R9_25, u2_R9_26, u2_R9_27, u2_R9_28, u2_R9_29, u2_R9_30, 
      u2_R9_31, u2_R9_32, u2_u11_X_37, u2_u11_X_38, u2_u11_X_39, u2_u11_X_40, u2_u14_X_21, u2_u14_X_22, u2_u14_X_23, 
      u2_u14_X_3, u2_u14_X_4, u2_uk_K_r10_10, u2_uk_K_r10_25, u2_uk_K_r10_27, u2_uk_K_r10_32, u2_uk_K_r10_34, u2_uk_K_r10_4, u2_uk_K_r10_41, 
      u2_uk_K_r10_43, u2_uk_K_r11_10, u2_uk_K_r11_11, u2_uk_K_r11_19, u2_uk_K_r11_20, u2_uk_K_r11_21, u2_uk_K_r11_24, u2_uk_K_r11_25, u2_uk_K_r11_26, 
      u2_uk_K_r11_27, u2_uk_K_r11_28, u2_uk_K_r11_29, u2_uk_K_r11_39, u2_uk_K_r11_47, u2_uk_K_r11_48, u2_uk_K_r11_53, u2_uk_K_r11_6, u2_uk_K_r12_10, 
      u2_uk_K_r12_15, u2_uk_K_r12_16, u2_uk_K_r12_25, u2_uk_K_r12_33, u2_uk_K_r13_19, u2_uk_K_r13_25, u2_uk_K_r13_32, u2_uk_K_r13_55, u2_uk_K_r14_15, 
      u2_uk_K_r14_16, u2_uk_K_r14_2, u2_uk_K_r14_50, u2_uk_K_r14_9, u2_uk_K_r6_0, u2_uk_K_r6_14, u2_uk_K_r6_29, u2_uk_K_r6_31, u2_uk_K_r6_37, 
      u2_uk_K_r6_51, u2_uk_K_r6_7, u2_uk_K_r7_0, u2_uk_K_r7_31, u2_uk_K_r7_37, u2_uk_K_r9_15, u2_uk_K_r9_23, u2_uk_K_r9_31, u2_uk_n10, 
      u2_uk_n100, u2_uk_n102, u2_uk_n109, u2_uk_n110, u2_uk_n1104, u2_uk_n1107, u2_uk_n1113, u2_uk_n1125, u2_uk_n1130, 
      u2_uk_n1132, u2_uk_n1133, u2_uk_n1134, u2_uk_n1136, u2_uk_n1137, u2_uk_n1140, u2_uk_n118, u2_uk_n1188, u2_uk_n1189, 
      u2_uk_n1200, u2_uk_n1201, u2_uk_n1203, u2_uk_n1208, u2_uk_n1209, u2_uk_n1210, u2_uk_n1215, u2_uk_n1217, u2_uk_n1220, 
      u2_uk_n1223, u2_uk_n1225, u2_uk_n1226, u2_uk_n128, u2_uk_n129, u2_uk_n145, u2_uk_n146, u2_uk_n147, u2_uk_n148, 
      u2_uk_n1498, u2_uk_n1499, u2_uk_n1503, u2_uk_n1504, u2_uk_n1511, u2_uk_n1517, u2_uk_n1524, u2_uk_n1525, u2_uk_n1526, 
      u2_uk_n1530, u2_uk_n1531, u2_uk_n1532, u2_uk_n1533, u2_uk_n1536, u2_uk_n1537, u2_uk_n1538, u2_uk_n1542, u2_uk_n1549, 
      u2_uk_n155, u2_uk_n1551, u2_uk_n1555, u2_uk_n1556, u2_uk_n1558, u2_uk_n1563, u2_uk_n1565, u2_uk_n1571, u2_uk_n1576, 
      u2_uk_n1577, u2_uk_n1583, u2_uk_n1585, u2_uk_n162, u2_uk_n163, u2_uk_n1632, u2_uk_n1634, u2_uk_n1642, u2_uk_n1647, 
      u2_uk_n1653, u2_uk_n1654, u2_uk_n1660, u2_uk_n1665, u2_uk_n1666, u2_uk_n1672, u2_uk_n1673, u2_uk_n1674, u2_uk_n1681, 
      u2_uk_n1682, u2_uk_n1683, u2_uk_n1684, u2_uk_n1687, u2_uk_n1688, u2_uk_n1689, u2_uk_n1693, u2_uk_n17, u2_uk_n1702, 
      u2_uk_n1707, u2_uk_n1708, u2_uk_n1720, u2_uk_n1721, u2_uk_n1723, u2_uk_n1724, u2_uk_n1725, u2_uk_n1726, u2_uk_n1727, 
      u2_uk_n1728, u2_uk_n1731, u2_uk_n1732, u2_uk_n1734, u2_uk_n1736, u2_uk_n1737, u2_uk_n1738, u2_uk_n1742, u2_uk_n1743, 
      u2_uk_n1744, u2_uk_n1745, u2_uk_n1746, u2_uk_n1747, u2_uk_n1750, u2_uk_n1753, u2_uk_n1755, u2_uk_n1761, u2_uk_n1762, 
      u2_uk_n1763, u2_uk_n1767, u2_uk_n1773, u2_uk_n1777, u2_uk_n1778, u2_uk_n1783, u2_uk_n1786, u2_uk_n1788, u2_uk_n1789, 
      u2_uk_n1790, u2_uk_n1794, u2_uk_n1796, u2_uk_n1800, u2_uk_n1801, u2_uk_n1805, u2_uk_n1811, u2_uk_n1814, u2_uk_n1815, 
      u2_uk_n1816, u2_uk_n182, u2_uk_n1821, u2_uk_n1823, u2_uk_n1832, u2_uk_n1833, u2_uk_n1834, u2_uk_n1839, u2_uk_n1843, 
      u2_uk_n1850, u2_uk_n1851, u2_uk_n1852, u2_uk_n187, u2_uk_n188, u2_uk_n191, u2_uk_n202, u2_uk_n208, u2_uk_n209, 
      u2_uk_n217, u2_uk_n220, u2_uk_n223, u2_uk_n230, u2_uk_n238, u2_uk_n31, u2_uk_n363, u2_uk_n369, u2_uk_n379, 
      u2_uk_n385, u2_uk_n415, u2_uk_n421, u2_uk_n443, u2_uk_n500, u2_uk_n503, u2_uk_n504, u2_uk_n526, u2_uk_n551, 
      u2_uk_n586, u2_uk_n60, u2_uk_n608, u2_uk_n63, u2_uk_n665, u2_uk_n677, u2_uk_n682, u2_uk_n83, u2_uk_n92, 
      u2_uk_n93, u2_uk_n931, u2_uk_n933, u2_uk_n94, u2_uk_n946, u2_uk_n947, u2_uk_n961, u2_uk_n99, u0_FP_11, 
      u0_FP_12, u0_FP_14, u0_FP_15, u0_FP_19, u0_FP_21, u0_FP_22, u0_FP_25, u0_FP_27, u0_FP_29, 
      u0_FP_3, u0_FP_32, u0_FP_4, u0_FP_5, u0_FP_7, u0_FP_8, u0_N128, u0_N129, u0_N130, 
      u0_N133, u0_N135, u0_N137, u0_N140, u0_N141, u0_N143, u0_N145, u0_N147, u0_N151, 
      u0_N152, u0_N153, u0_N155, u0_N157, u0_N256, u0_N257, u0_N258, u0_N259, u0_N260, 
      u0_N261, u0_N262, u0_N263, u0_N264, u0_N265, u0_N266, u0_N267, u0_N268, u0_N269, 
      u0_N270, u0_N271, u0_N272, u0_N273, u0_N274, u0_N275, u0_N276, u0_N277, u0_N278, 
      u0_N279, u0_N280, u0_N281, u0_N282, u0_N283, u0_N284, u0_N285, u0_N286, u0_N287, 
      u0_N288, u0_N289, u0_N293, u0_N297, u0_N300, u0_N303, u0_N305, u0_N307, u0_N311, 
      u0_N313, u0_N315, u0_N317, u0_N352, u0_N353, u0_N354, u0_N355, u0_N356, u0_N357, 
      u0_N358, u0_N359, u0_N360, u0_N361, u0_N362, u0_N363, u0_N364, u0_N365, u0_N366, 
      u0_N367, u0_N368, u0_N369, u0_N370, u0_N371, u0_N372, u0_N373, u0_N374, u0_N375, 
      u0_N376, u0_N377, u0_N378, u0_N379, u0_N380, u0_N381, u0_N382, u0_N383, u0_N417, 
      u0_N421, u0_N424, u0_N428, u0_N431, u0_N432, u0_N433, u0_N438, u0_N439, u0_N443, 
      u0_N445, u0_N446, u0_uk_n10, u0_uk_n100, u0_uk_n117, u0_uk_n128, u0_uk_n129, u0_uk_n146, u0_uk_n148, 
      u0_uk_n161, u0_uk_n182, u0_uk_n187, u0_uk_n203, u0_uk_n208, u0_uk_n214, u0_uk_n240, u0_uk_n251, u0_uk_n27, 
      u0_uk_n99, u1_K10_10, u1_K10_15, u1_K10_16, u1_K10_17, u1_K10_18, u1_K10_19, u1_K10_20, u1_K10_21, 
      u1_K10_27, u1_K10_28, u1_K10_34, u1_K10_45, u1_K10_46, u1_K11_1, u1_K11_10, u1_K11_11, u1_K11_13, 
      u1_K11_15, u1_K11_16, u1_K11_3, u1_K11_4, u1_K11_45, u1_K11_6, u1_K11_9, u1_K12_10, u1_K12_11, 
      u1_K12_12, u1_K12_13, u1_K12_14, u1_K12_16, u1_K12_33, u1_K12_34, u1_K12_36, u1_K12_38, u1_K12_39, 
      u1_K12_40, u1_K12_41, u1_K12_43, u1_K12_45, u1_K12_46, u1_K12_5, u1_K12_7, u1_K12_9, u1_K13_1, 
      u1_K13_24, u1_K13_26, u1_K13_27, u1_K13_28, u1_K13_3, u1_K13_33, u1_K13_34, u1_K13_35, u1_K13_36, 
      u1_K13_37, u1_K13_38, u1_K13_39, u1_K13_4, u1_K13_40, u1_K13_45, u1_K13_46, u1_K13_47, u1_K13_8, 
      u1_K13_9, u1_K14_10, u1_K14_12, u1_K14_14, u1_K14_15, u1_K14_16, u1_K14_21, u1_K14_22, u1_K14_27, 
      u1_K14_28, u1_K14_29, u1_K14_3, u1_K14_31, u1_K14_33, u1_K14_4, u1_K14_9, u1_K15_10, u1_K15_12, 
      u1_K15_14, u1_K15_15, u1_K15_16, u1_K15_17, u1_K15_18, u1_K15_19, u1_K15_20, u1_K15_21, u1_K15_22, 
      u1_K15_27, u1_K15_28, u1_K15_3, u1_K15_33, u1_K15_34, u1_K15_4, u1_K15_45, u1_K15_46, u1_K15_5, 
      u1_K15_6, u1_K15_7, u1_K15_9, u1_K16_10, u1_K16_15, u1_K16_16, u1_K16_21, u1_K16_22, u1_K16_24, 
      u1_K16_26, u1_K16_27, u1_K16_28, u1_K16_3, u1_K16_39, u1_K16_4, u1_K16_40, u1_K16_6, u1_K16_8, 
      u1_K16_9, u1_K1_12, u1_K1_14, u1_K1_15, u1_K1_16, u1_K1_21, u1_K1_3, u1_K1_34, u1_K1_39, 
      u1_K1_4, u1_K1_40, u1_K1_43, u1_K1_45, u1_K1_46, u1_K1_9, u1_K2_1, u1_K2_21, u1_K2_22, 
      u1_K2_3, u1_K2_33, u1_K2_34, u1_K2_39, u1_K2_4, u1_K2_40, u1_K2_45, u1_K2_46, u1_K2_47, 
      u1_K3_10, u1_K3_15, u1_K3_16, u1_K3_27, u1_K3_28, u1_K3_3, u1_K3_39, u1_K3_4, u1_K3_40, 
      u1_K3_5, u1_K3_7, u1_K3_9, u1_K4_15, u1_K4_16, u1_K4_17, u1_K4_18, u1_K4_19, u1_K4_21, 
      u1_K4_22, u1_K4_24, u1_K4_27, u1_K4_28, u1_K4_39, u1_K4_40, u1_K4_45, u1_K4_46, u1_K4_9, 
      u1_K5_10, u1_K5_15, u1_K5_16, u1_K5_18, u1_K5_21, u1_K5_23, u1_K5_24, u1_K5_25, u1_K5_26, 
      u1_K5_28, u1_K5_29, u1_K5_30, u1_K5_31, u1_K5_32, u1_K5_33, u1_K5_34, u1_K5_37, u1_K5_38, 
      u1_K5_39, u1_K5_40, u1_K5_41, u1_K5_45, u1_K5_46, u1_K5_9, u1_K6_1, u1_K6_22, u1_K6_3, 
      u1_K6_33, u1_K6_34, u1_K6_35, u1_K6_36, u1_K6_37, u1_K6_38, u1_K6_39, u1_K6_40, u1_K6_41, 
      u1_K6_42, u1_K6_43, u1_K6_44, u1_K6_45, u1_K6_46, u1_K6_47, u1_K6_48, u1_K6_6, u1_K6_8, 
      u1_K7_10, u1_K7_11, u1_K7_14, u1_K7_15, u1_K7_16, u1_K7_17, u1_K7_18, u1_K7_19, u1_K7_21, 
      u1_K7_22, u1_K7_23, u1_K7_26, u1_K7_28, u1_K7_29, u1_K7_3, u1_K7_30, u1_K7_31, u1_K7_33, 
      u1_K7_39, u1_K7_4, u1_K7_40, u1_K7_41, u1_K7_43, u1_K7_45, u1_K7_5, u1_K7_7, u1_K7_9, 
      u1_K8_10, u1_K8_11, u1_K8_13, u1_K8_14, u1_K8_16, u1_K8_18, u1_K8_20, u1_K8_21, u1_K8_22, 
      u1_K8_23, u1_K8_25, u1_K8_27, u1_K8_28, u1_K8_4, u1_K8_45, u1_K8_46, u1_K8_5, u1_K8_6, 
      u1_K8_7, u1_K8_8, u1_K8_9, u1_K9_13, u1_K9_15, u1_K9_16, u1_K9_17, u1_K9_21, u1_K9_23, 
      u1_K9_24, u1_K9_25, u1_K9_28, u1_K9_3, u1_K9_34, u1_K9_36, u1_K9_37, u1_K9_38, u1_K9_39, 
      u1_K9_4, u1_K9_40, u1_out0_14, u1_out0_25, u1_out0_3, u1_out0_8, u1_out10_1, u1_out10_10, u1_out10_11, 
      u1_out10_12, u1_out10_14, u1_out10_19, u1_out10_20, u1_out10_22, u1_out10_25, u1_out10_26, u1_out10_29, u1_out10_3, 
      u1_out10_32, u1_out10_4, u1_out10_7, u1_out10_8, u1_out11_1, u1_out11_10, u1_out11_14, u1_out11_20, u1_out11_25, 
      u1_out11_26, u1_out11_3, u1_out11_8, u1_out12_16, u1_out12_24, u1_out12_30, u1_out12_6, u1_out13_12, u1_out13_15, 
      u1_out13_21, u1_out13_22, u1_out13_27, u1_out13_32, u1_out13_5, u1_out13_7, u1_out14_12, u1_out14_22, u1_out14_32, 
      u1_out14_7, u1_out15_11, u1_out15_15, u1_out15_19, u1_out15_21, u1_out15_27, u1_out15_29, u1_out15_4, u1_out15_5, 
      u1_out1_13, u1_out1_16, u1_out1_18, u1_out1_2, u1_out1_24, u1_out1_28, u1_out1_30, u1_out1_6, u1_out2_1, 
      u1_out2_10, u1_out2_11, u1_out2_15, u1_out2_19, u1_out2_20, u1_out2_21, u1_out2_26, u1_out2_27, u1_out2_29, 
      u1_out2_4, u1_out2_5, u1_out3_11, u1_out3_17, u1_out3_19, u1_out3_23, u1_out3_29, u1_out3_31, u1_out3_4, 
      u1_out3_9, u1_out4_17, u1_out4_23, u1_out4_31, u1_out4_9, u1_out5_14, u1_out5_16, u1_out5_24, u1_out5_25, 
      u1_out5_3, u1_out5_30, u1_out5_6, u1_out5_8, u1_out7_11, u1_out7_12, u1_out7_19, u1_out7_22, u1_out7_29, 
      u1_out7_32, u1_out7_4, u1_out7_7, u1_out8_15, u1_out8_21, u1_out8_27, u1_out8_5, u1_out9_12, u1_out9_17, 
      u1_out9_22, u1_out9_23, u1_out9_31, u1_out9_32, u1_out9_7, u1_out9_9, u1_u0_X_1, u1_u0_X_11, u1_u0_X_13, 
      u1_u0_X_17, u1_u0_X_18, u1_u0_X_19, u1_u0_X_2, u1_u0_X_20, u1_u0_X_23, u1_u0_X_24, u1_u0_X_31, u1_u0_X_32, 
      u1_u0_X_35, u1_u0_X_36, u1_u0_X_37, u1_u0_X_38, u1_u0_X_47, u1_u0_X_48, u1_u0_X_5, u1_u0_X_6, u1_u0_X_7, 
      u1_u0_X_8, u1_u10_X_17, u1_u10_X_18, u1_u10_X_2, u1_u10_X_43, u1_u10_X_44, u1_u10_X_48, u1_u10_X_5, u1_u10_X_7, 
      u1_u11_X_1, u1_u11_X_17, u1_u11_X_18, u1_u11_X_2, u1_u11_X_31, u1_u11_X_32, u1_u11_X_35, u1_u11_X_37, u1_u11_X_42, 
      u1_u11_X_44, u1_u11_X_47, u1_u11_X_48, u1_u11_X_6, u1_u11_X_8, u1_u12_X_11, u1_u12_X_12, u1_u12_X_19, u1_u12_X_2, 
      u1_u12_X_20, u1_u12_X_23, u1_u12_X_25, u1_u12_X_29, u1_u12_X_30, u1_u12_X_31, u1_u12_X_32, u1_u12_X_41, u1_u12_X_42, 
      u1_u12_X_43, u1_u12_X_44, u1_u12_X_48, u1_u12_X_5, u1_u12_X_7, u1_u13_X_1, u1_u13_X_11, u1_u13_X_13, u1_u13_X_17, 
      u1_u13_X_18, u1_u13_X_19, u1_u13_X_2, u1_u13_X_20, u1_u13_X_23, u1_u13_X_24, u1_u13_X_25, u1_u13_X_26, u1_u13_X_30, 
      u1_u13_X_32, u1_u13_X_35, u1_u13_X_36, u1_u13_X_5, u1_u13_X_6, u1_u13_X_7, u1_u13_X_8, u1_u14_X_1, u1_u14_X_11, 
      u1_u14_X_13, u1_u14_X_2, u1_u14_X_23, u1_u14_X_24, u1_u14_X_25, u1_u14_X_26, u1_u14_X_29, u1_u14_X_30, u1_u14_X_31, 
      u1_u14_X_32, u1_u14_X_35, u1_u14_X_36, u1_u14_X_43, u1_u14_X_44, u1_u14_X_47, u1_u14_X_48, u1_u15_X_1, u1_u15_X_11, 
      u1_u15_X_12, u1_u15_X_13, u1_u15_X_14, u1_u15_X_17, u1_u15_X_18, u1_u15_X_19, u1_u15_X_2, u1_u15_X_20, u1_u15_X_23, 
      u1_u15_X_25, u1_u15_X_29, u1_u15_X_30, u1_u15_X_37, u1_u15_X_38, u1_u15_X_41, u1_u15_X_42, u1_u15_X_5, u1_u15_X_7, 
      u1_u1_X_19, u1_u1_X_2, u1_u1_X_20, u1_u1_X_23, u1_u1_X_24, u1_u1_X_25, u1_u1_X_26, u1_u1_X_29, u1_u1_X_30, 
      u1_u1_X_31, u1_u1_X_32, u1_u1_X_35, u1_u1_X_36, u1_u1_X_37, u1_u1_X_38, u1_u1_X_41, u1_u1_X_42, u1_u1_X_43, 
      u1_u1_X_44, u1_u1_X_48, u1_u1_X_5, u1_u1_X_6, u1_u2_X_1, u1_u2_X_11, u1_u2_X_12, u1_u2_X_13, u1_u2_X_14, 
      u1_u2_X_17, u1_u2_X_18, u1_u2_X_2, u1_u2_X_25, u1_u2_X_26, u1_u2_X_29, u1_u2_X_30, u1_u2_X_37, u1_u2_X_38, 
      u1_u2_X_41, u1_u2_X_42, u1_u2_X_6, u1_u2_X_8, u1_u3_X_11, u1_u3_X_12, u1_u3_X_13, u1_u3_X_14, u1_u3_X_29, 
      u1_u3_X_30, u1_u3_X_37, u1_u3_X_38, u1_u3_X_41, u1_u3_X_42, u1_u3_X_43, u1_u3_X_44, u1_u3_X_47, u1_u3_X_48, 
      u1_u3_X_7, u1_u3_X_8, u1_u4_X_11, u1_u4_X_12, u1_u4_X_13, u1_u4_X_14, u1_u4_X_17, u1_u4_X_19, u1_u4_X_42, 
      u1_u4_X_44, u1_u4_X_47, u1_u4_X_48, u1_u4_X_7, u1_u4_X_8, u1_u5_X_11, u1_u5_X_12, u1_u5_X_19, u1_u5_X_20, 
      u1_u5_X_23, u1_u5_X_24, u1_u5_X_31, u1_u5_X_32, u1_u5_X_5, u1_u5_X_7, u1_u6_X_1, u1_u6_X_2, u1_u6_X_35, 
      u1_u6_X_36, u1_u6_X_37, u1_u6_X_38, u1_u6_X_42, u1_u6_X_44, u1_u6_X_47, u1_u6_X_48, u1_u7_X_1, u1_u7_X_17, 
      u1_u7_X_19, u1_u7_X_2, u1_u7_X_24, u1_u7_X_26, u1_u7_X_29, u1_u7_X_30, u1_u7_X_43, u1_u7_X_44, u1_u7_X_47, 
      u1_u7_X_48, u1_u8_X_1, u1_u8_X_12, u1_u8_X_14, u1_u8_X_2, u1_u8_X_29, u1_u8_X_30, u1_u8_X_31, u1_u8_X_32, 
      u1_u8_X_41, u1_u8_X_42, u1_u8_X_5, u1_u8_X_6, u1_u8_X_7, u1_u8_X_8, u1_u9_X_11, u1_u9_X_12, u1_u9_X_13, 
      u1_u9_X_14, u1_u9_X_23, u1_u9_X_24, u1_u9_X_25, u1_u9_X_26, u1_u9_X_29, u1_u9_X_30, u1_u9_X_31, u1_u9_X_32, 
      u1_u9_X_35, u1_u9_X_36, u1_u9_X_43, u1_u9_X_44, u1_u9_X_47, u1_u9_X_48, u1_u9_X_7, u1_u9_X_8, u1_uk_n1004, 
      u1_uk_n1011, u1_uk_n1015, u1_uk_n1016, u1_uk_n1017, u1_uk_n1027, u1_uk_n1028, u1_uk_n1050, u1_uk_n1054, u1_uk_n1056, 
      u1_uk_n1057, u1_uk_n1058, u1_uk_n1073, u1_uk_n1074, u1_uk_n1076, u1_uk_n1079, u1_uk_n1080, u1_uk_n1083, u1_uk_n1088, 
      u1_uk_n1092, u1_uk_n1096, u1_uk_n1101, u1_uk_n1104, u1_uk_n1105, u1_uk_n1106, u1_uk_n1109, u1_uk_n1113, u1_uk_n1114, 
      u1_uk_n1115, u1_uk_n1118, u1_uk_n1119, u1_uk_n1124, u1_uk_n1125, u1_uk_n1126, u1_uk_n1128, u1_uk_n1130, u1_uk_n1140, 
      u1_uk_n1147, u1_uk_n1148, u1_uk_n1153, u1_uk_n1154, u1_uk_n1156, u1_uk_n1157, u1_uk_n1158, u1_uk_n1159, u1_uk_n1162, 
      u1_uk_n1163, u1_uk_n1171, u1_uk_n312, u1_uk_n349, u1_uk_n376, u1_uk_n379, u1_uk_n382, u1_uk_n468, u1_uk_n472, 
      u1_uk_n501, u1_uk_n504, u1_uk_n601, u1_uk_n656, u1_uk_n671, u1_uk_n689, u1_uk_n692, u1_uk_n949, u1_uk_n955, 
      u1_uk_n976, u1_uk_n996, u2_FP_11, u2_FP_12, u2_FP_15, u2_FP_19, u2_FP_21, u2_FP_22, u2_FP_27, 
      u2_FP_29, u2_FP_32, u2_FP_4, u2_FP_5, u2_FP_7, u2_N226, u2_N227, u2_N228, u2_N230, 
      u2_N231, u2_N234, u2_N237, u2_N238, u2_N242, u2_N244, u2_N245, u2_N248, u2_N250, 
      u2_N252, u2_N255, u2_N259, u2_N260, u2_N262, u2_N264, u2_N266, u2_N267, u2_N270, 
      u2_N272, u2_N274, u2_N276, u2_N277, u2_N278, u2_N282, u2_N284, u2_N286, u2_N287, 
      u2_N322, u2_N324, u2_N326, u2_N327, u2_N331, u2_N333, u2_N334, u2_N340, u2_N341, 
      u2_N344, u2_N346, u2_N351, u2_N352, u2_N356, u2_N357, u2_N360, u2_N361, u2_N366, 
      u2_N367, u2_N368, u2_N371, u2_N372, u2_N374, u2_N375, u2_N377, u2_N378, u2_N381, 
      u2_N382, u2_N384, u2_N385, u2_N386, u2_N387, u2_N388, u2_N389, u2_N390, u2_N391, 
      u2_N392, u2_N393, u2_N394, u2_N395, u2_N396, u2_N397, u2_N398, u2_N399, u2_N400, 
      u2_N401, u2_N402, u2_N403, u2_N404, u2_N405, u2_N406, u2_N407, u2_N408, u2_N409, 
      u2_N413, u2_N414, u2_N415, u2_N417, u2_N420, u2_N421, u2_N424, u2_N428, u2_N430, 
      u2_N431, u2_N432, u2_N433, u2_N436, u2_N438, u2_N439, u2_N442, u2_N443, u2_N445, 
      u2_N446, u2_N449, u2_N453, u2_N460, u2_N463, u2_N465, u2_N471, u2_N475, u2_N477, 
      u2_out11_12, u2_out11_22, u2_out11_32, u2_out11_7, u2_out12_27, u2_out12_28, u2_out12_29, u2_out14_1, u2_out14_10, 
      u2_out14_17, u2_out14_20, u2_out14_23, u2_out14_26, u2_out14_31, u2_out14_9, u2_out7_12, u2_u13_X_19, u2_u13_X_20, 
      u2_uk_n11, u2_uk_n117, u2_uk_n141, u2_uk_n142, u2_uk_n161, u2_uk_n203, u2_uk_n207, u2_uk_n213, u2_uk_n214, 
      u2_uk_n222, u2_uk_n231, u2_uk_n27 );
  des_des_die_5 u5 ( u0_FP_33, u0_FP_34, u0_FP_36, u0_FP_37, u0_FP_38, u0_FP_39, u0_FP_40, u0_FP_41, u0_FP_42, 
      u0_FP_43, u0_FP_45, u0_FP_48, u0_FP_49, u0_FP_64, u0_K13_8, u0_K14_42, u0_K16_11, u0_K16_18, 
      u0_K16_24, u0_K16_8, u0_K1_31, u0_K1_47, u0_K2_5, u0_K2_6, u0_K2_8, u0_K6_11, u0_K6_13, 
      u0_K6_20, u0_K6_23, u0_K8_19, u0_K8_23, u0_R0_4, u0_R0_5, u0_R11_28, u0_R11_3, u0_R11_32, 
      u0_R11_4, u0_R11_5, u0_R11_6, u0_R11_7, u0_R11_8, u0_R11_9, u0_R12_1, u0_R12_20, u0_R12_21, 
      u0_R12_22, u0_R12_23, u0_R12_24, u0_R12_25, u0_R12_26, u0_R12_28, u0_R12_29, u0_R12_30, u0_R12_32, 
      u0_R2_1, u0_R2_10, u0_R2_11, u0_R2_12, u0_R2_13, u0_R2_3, u0_R2_32, u0_R2_4, u0_R2_6, 
      u0_R2_7, u0_R2_8, u0_R2_9, u0_R4_13, u0_R4_14, u0_R4_16, u0_R4_8, u0_R6_1, u0_R6_12, 
      u0_R6_13, u0_R6_14, u0_R6_16, u0_R6_17, u0_R6_18, u0_R6_20, u0_R6_21, u0_R6_23, u0_R6_24, 
      u0_R6_28, u0_R6_29, u0_R6_32, u0_R9_10, u0_R9_11, u0_R9_12, u0_R9_13, u0_R9_15, u0_R9_16, 
      u0_R9_17, u0_R9_8, u0_R9_9, u0_desIn_r_1, u0_desIn_r_11, u0_desIn_r_25, u0_desIn_r_27, u0_desIn_r_3, u0_desIn_r_33, 
      u0_desIn_r_51, u0_desIn_r_57, u0_desIn_r_59, u0_desIn_r_7, u0_key_r_14, u0_key_r_16, u0_key_r_2, u0_key_r_21, u0_key_r_23, 
      u0_key_r_28, u0_key_r_30, u0_key_r_31, u0_key_r_35, u0_key_r_36, u0_key_r_37, u0_key_r_38, u0_key_r_42, u0_key_r_43, 
      u0_key_r_50, u0_key_r_51, u0_key_r_9, u0_u0_X_25, u0_u0_X_28, u0_u0_X_30, u0_u0_X_32, u0_u0_X_33, u0_u0_X_39, 
      u0_u0_X_40, u0_u0_X_45, u0_u0_X_46, u0_u10_X_21, u0_u12_X_2, u0_u12_X_3, u0_u12_X_44, u0_u12_X_45, u0_u12_X_46, 
      u0_u12_X_48, u0_u13_X_40, u0_u13_X_46, u0_u15_X_17, u0_u15_X_19, u0_u15_X_21, u0_u15_X_22, u0_u15_X_4, u0_u1_X_1, 
      u0_u1_X_10, u0_u1_X_11, u0_u1_X_12, u0_u1_X_2, u0_u1_X_3, u0_u1_X_4, u0_u1_X_9, u0_u3_X_3, u0_u3_X_6, 
      u0_u3_X_8, u0_u5_X_10, u0_u5_X_12, u0_u5_X_14, u0_u5_X_15, u0_u5_X_16, u0_u5_X_17, u0_u5_X_19, u0_u5_X_22, 
      u0_u5_X_24, u0_u5_X_26, u0_u5_X_27, u0_u5_X_28, u0_u5_X_29, u0_u5_X_30, u0_u5_X_7, u0_u5_X_8, u0_u5_X_9, 
      u0_u7_X_22, u0_u7_X_28, u0_u7_X_33, u0_u7_X_36, u0_u7_X_45, u0_u7_X_46, u0_uk_K_r11_17, u0_uk_K_r11_25, u0_uk_K_r11_29, 
      u0_uk_K_r11_34, u0_uk_K_r11_48, u0_uk_K_r11_53, u0_uk_K_r11_54, u0_uk_K_r12_15, u0_uk_K_r12_16, u0_uk_K_r14_11, u0_uk_K_r14_12, u0_uk_K_r14_18, 
      u0_uk_K_r14_46, u0_uk_K_r2_13, u0_uk_K_r2_18, u0_uk_K_r2_20, u0_uk_K_r2_25, u0_uk_K_r2_27, u0_uk_K_r2_53, u0_uk_K_r6_0, u0_uk_K_r6_14, 
      u0_uk_K_r6_21, u0_uk_K_r6_29, u0_uk_K_r9_13, u0_uk_K_r9_19, u0_uk_K_r9_27, u0_uk_n10, u0_uk_n100, u0_uk_n1000, u0_uk_n1001, 
      u0_uk_n1002, u0_uk_n102, u0_uk_n106, u0_uk_n109, u0_uk_n11, u0_uk_n115, u0_uk_n117, u0_uk_n118, u0_uk_n121, 
      u0_uk_n126, u0_uk_n127, u0_uk_n128, u0_uk_n129, u0_uk_n131, u0_uk_n141, u0_uk_n142, u0_uk_n145, u0_uk_n146, 
      u0_uk_n161, u0_uk_n163, u0_uk_n182, u0_uk_n187, u0_uk_n188, u0_uk_n190, u0_uk_n196, u0_uk_n197, u0_uk_n200, 
      u0_uk_n201, u0_uk_n202, u0_uk_n203, u0_uk_n206, u0_uk_n208, u0_uk_n212, u0_uk_n213, u0_uk_n214, u0_uk_n215, 
      u0_uk_n217, u0_uk_n220, u0_uk_n221, u0_uk_n223, u0_uk_n240, u0_uk_n242, u0_uk_n251, u0_uk_n257, u0_uk_n27, 
      u0_uk_n318, u0_uk_n320, u0_uk_n321, u0_uk_n325, u0_uk_n327, u0_uk_n330, u0_uk_n331, u0_uk_n332, u0_uk_n333, 
      u0_uk_n336, u0_uk_n337, u0_uk_n341, u0_uk_n347, u0_uk_n348, u0_uk_n354, u0_uk_n355, u0_uk_n358, u0_uk_n359, 
      u0_uk_n418, u0_uk_n434, u0_uk_n497, u0_uk_n50, u0_uk_n502, u0_uk_n51, u0_uk_n510, u0_uk_n517, u0_uk_n519, 
      u0_uk_n52, u0_uk_n525, u0_uk_n529, u0_uk_n530, u0_uk_n531, u0_uk_n534, u0_uk_n535, u0_uk_n536, u0_uk_n55, 
      u0_uk_n56, u0_uk_n58, u0_uk_n59, u0_uk_n61, u0_uk_n629, u0_uk_n630, u0_uk_n631, u0_uk_n636, u0_uk_n637, 
      u0_uk_n639, u0_uk_n640, u0_uk_n644, u0_uk_n645, u0_uk_n65, u0_uk_n651, u0_uk_n652, u0_uk_n653, u0_uk_n659, 
      u0_uk_n660, u0_uk_n664, u0_uk_n667, u0_uk_n668, u0_uk_n67, u0_uk_n68, u0_uk_n73, u0_uk_n746, u0_uk_n755, 
      u0_uk_n77, u0_uk_n797, u0_uk_n799, u0_uk_n81, u0_uk_n82, u0_uk_n828, u0_uk_n83, u0_uk_n839, u0_uk_n855, 
      u0_uk_n88, u0_uk_n89, u0_uk_n90, u0_uk_n92, u0_uk_n93, u0_uk_n933, u0_uk_n934, u0_uk_n939, u0_uk_n94, 
      u0_uk_n940, u0_uk_n96, u0_uk_n960, u0_uk_n99, u0_uk_n999, u1_FP_34, u1_FP_35, u1_FP_37, u1_FP_38, 
      u1_FP_39, u1_K10_15, u1_K10_16, u1_K10_17, u1_K10_18, u1_K10_19, u1_K10_20, u1_K10_21, u1_K10_45, 
      u1_K10_46, u1_K11_10, u1_K11_11, u1_K11_13, u1_K11_15, u1_K11_16, u1_K11_9, u1_K12_10, u1_K12_11, 
      u1_K12_12, u1_K12_13, u1_K12_14, u1_K12_16, u1_K12_5, u1_K12_7, u1_K12_9, u1_K13_1, u1_K13_24, 
      u1_K13_26, u1_K13_27, u1_K13_28, u1_K13_3, u1_K13_4, u1_K13_45, u1_K13_46, u1_K13_47, u1_K15_14, 
      u1_K15_15, u1_K15_16, u1_K15_17, u1_K15_18, u1_K15_19, u1_K15_20, u1_K15_21, u1_K15_22, u1_K16_10, 
      u1_K16_3, u1_K16_4, u1_K16_6, u1_K16_8, u1_K16_9, u1_K1_21, u1_K1_3, u1_K1_4, u1_K2_33, 
      u1_K2_34, u1_K3_10, u1_K3_3, u1_K3_4, u1_K3_5, u1_K3_7, u1_K3_9, u1_K4_45, u1_K4_46, 
      u1_K5_10, u1_K5_9, u1_K6_1, u1_K6_22, u1_K6_3, u1_K6_33, u1_K6_34, u1_K6_35, u1_K6_36, 
      u1_K6_37, u1_K6_38, u1_K6_39, u1_K6_40, u1_K6_41, u1_K6_42, u1_K6_43, u1_K6_44, u1_K6_45, 
      u1_K6_46, u1_K6_47, u1_K6_48, u1_K6_6, u1_K6_8, u1_K8_45, u1_K8_46, u1_R0_22, u1_R0_23, 
      u1_R10_10, u1_R10_11, u1_R10_2, u1_R10_3, u1_R10_4, u1_R10_6, u1_R10_7, u1_R10_8, u1_R10_9, 
      u1_R11_14, u1_R11_15, u1_R11_17, u1_R11_18, u1_R11_19, u1_R11_2, u1_R11_3, u1_R11_30, u1_R11_31, 
      u1_R11_32, u1_R11_5, u1_R13_10, u1_R13_11, u1_R13_12, u1_R13_13, u1_R13_14, u1_R13_15, u1_R13_9, 
      u1_R1_2, u1_R1_3, u1_R1_4, u1_R1_6, u1_R1_7, u1_R2_30, u1_R2_31, u1_R3_6, u1_R3_7, 
      u1_R4_1, u1_R4_14, u1_R4_15, u1_R4_2, u1_R4_22, u1_R4_23, u1_R4_24, u1_R4_25, u1_R4_26, 
      u1_R4_27, u1_R4_28, u1_R4_29, u1_R4_3, u1_R4_30, u1_R4_31, u1_R4_32, u1_R4_5, u1_R4_6, 
      u1_R4_7, u1_R6_30, u1_R6_31, u1_R7_6, u1_R7_7, u1_R7_8, u1_R8_10, u1_R8_11, u1_R8_12, 
      u1_R8_13, u1_R8_14, u1_R8_15, u1_R8_30, u1_R8_31, u1_R9_10, u1_R9_11, u1_R9_5, u1_R9_6, 
      u1_R9_7, u1_R9_8, u1_R9_9, u1_desIn_r_15, u1_desIn_r_23, u1_desIn_r_45, u1_desIn_r_53, u1_u0_X_1, u1_u0_X_19, 
      u1_u0_X_2, u1_u0_X_20, u1_u0_X_23, u1_u0_X_24, u1_u0_X_5, u1_u0_X_6, u1_u10_X_17, u1_u10_X_18, u1_u10_X_7, 
      u1_u11_X_1, u1_u11_X_17, u1_u11_X_18, u1_u11_X_2, u1_u11_X_6, u1_u11_X_8, u1_u12_X_19, u1_u12_X_2, u1_u12_X_20, 
      u1_u12_X_23, u1_u12_X_25, u1_u12_X_29, u1_u12_X_30, u1_u12_X_43, u1_u12_X_44, u1_u12_X_48, u1_u12_X_5, u1_u14_X_13, 
      u1_u14_X_23, u1_u14_X_24, u1_u15_X_1, u1_u15_X_11, u1_u15_X_12, u1_u15_X_2, u1_u15_X_5, u1_u15_X_7, u1_u1_X_31, 
      u1_u1_X_32, u1_u1_X_35, u1_u1_X_36, u1_u2_X_1, u1_u2_X_11, u1_u2_X_12, u1_u2_X_2, u1_u2_X_6, u1_u2_X_8, 
      u1_u3_X_43, u1_u3_X_44, u1_u3_X_47, u1_u3_X_48, u1_u4_X_11, u1_u4_X_12, u1_u4_X_7, u1_u4_X_8, u1_u5_X_11, 
      u1_u5_X_12, u1_u5_X_19, u1_u5_X_20, u1_u5_X_23, u1_u5_X_24, u1_u5_X_31, u1_u5_X_32, u1_u5_X_5, u1_u5_X_7, 
      u1_u7_X_43, u1_u7_X_44, u1_u7_X_47, u1_u7_X_48, u1_u8_X_12, u1_u8_X_7, u1_u8_X_8, u1_u9_X_13, u1_u9_X_14, 
      u1_u9_X_23, u1_u9_X_24, u1_u9_X_43, u1_u9_X_44, u1_u9_X_47, u1_u9_X_48, u1_uk_n1004, u1_uk_n1088, u1_uk_n1092, 
      u1_uk_n1096, u1_uk_n1101, u1_uk_n1104, u1_uk_n1147, u1_uk_n1148, u1_uk_n1171, u1_uk_n312, u1_uk_n379, u1_uk_n382, 
      u1_uk_n501, u1_uk_n504, u1_uk_n601, u1_uk_n656, u1_uk_n689, u1_uk_n692, u1_uk_n949, u2_K10_36, u2_K15_29, 
      u2_K15_31, u2_K15_35, u2_K1_30, u2_K1_37, u2_K1_43, u2_R13_17, u2_R13_18, u2_R13_20, u2_R13_22, 
      u2_R13_24, u2_R13_25, u2_R8_20, u2_R8_22, u2_R8_24, u2_R8_25, u2_desIn_r_1, u2_desIn_r_11, u2_desIn_r_25, 
      u2_desIn_r_27, u2_desIn_r_3, u2_desIn_r_33, u2_desIn_r_35, u2_desIn_r_43, u2_desIn_r_57, u2_desIn_r_59, u2_desIn_r_61, u2_desIn_r_7, 
      u2_desIn_r_9, u2_key_r_0, u2_key_r_14, u2_key_r_16, u2_key_r_21, u2_key_r_22, u2_key_r_23, u2_key_r_28, u2_key_r_29, 
      u2_key_r_30, u2_key_r_31, u2_key_r_35, u2_key_r_36, u2_key_r_37, u2_key_r_42, u2_key_r_43, u2_key_r_44, u2_key_r_51, 
      u2_key_r_7, u2_u0_X_28, u2_u0_X_34, u2_u0_X_40, u2_u0_X_45, u2_u0_X_46, u2_u14_X_25, u2_u14_X_28, u2_u14_X_30, 
      u2_u14_X_32, u2_u14_X_34, u2_u9_X_32, u2_u9_X_34, u2_uk_K_r8_16, u2_uk_K_r8_2, u2_uk_K_r8_22, u2_uk_K_r8_37, u2_uk_K_r8_42, 
      u2_uk_n10, u2_uk_n100, u2_uk_n102, u2_uk_n109, u2_uk_n117, u2_uk_n118, u2_uk_n128, u2_uk_n142, u2_uk_n155, 
      u2_uk_n1615, u2_uk_n162, u2_uk_n163, u2_uk_n164, u2_uk_n1817, u2_uk_n182, u2_uk_n1826, u2_uk_n1835, u2_uk_n1840, 
      u2_uk_n203, u2_uk_n207, u2_uk_n208, u2_uk_n217, u2_uk_n222, u2_uk_n238, u2_uk_n31, u2_uk_n60, u2_uk_n63, 
      u2_uk_n92, u2_uk_n939, u2_uk_n94, u2_uk_n942, u2_uk_n984, u2_uk_n986, u2_uk_n99, u0_out0_11, u0_out0_12, 
      u0_out0_14, u0_out0_15, u0_out0_19, u0_out0_21, u0_out0_22, u0_out0_25, u0_out0_27, u0_out0_29, u0_out0_3, 
      u0_out0_32, u0_out0_4, u0_out0_5, u0_out0_7, u0_out0_8, u0_out10_1, u0_out10_10, u0_out10_16, u0_out10_20, 
      u0_out10_24, u0_out10_26, u0_out10_30, u0_out10_6, u0_out12_13, u0_out12_15, u0_out12_17, u0_out12_18, u0_out12_2, 
      u0_out12_21, u0_out12_23, u0_out12_27, u0_out12_28, u0_out12_31, u0_out12_5, u0_out12_9, u0_out13_11, u0_out13_12, 
      u0_out13_15, u0_out13_19, u0_out13_21, u0_out13_22, u0_out13_27, u0_out13_29, u0_out13_32, u0_out13_4, u0_out13_5, 
      u0_out13_7, u0_out15_1, u0_out15_10, u0_out15_13, u0_out15_16, u0_out15_17, u0_out15_18, u0_out15_2, u0_out15_20, 
      u0_out15_23, u0_out15_24, u0_out15_26, u0_out15_28, u0_out15_30, u0_out15_31, u0_out15_6, u0_out15_9, u0_out1_13, 
      u0_out1_17, u0_out1_18, u0_out1_2, u0_out1_23, u0_out1_28, u0_out1_31, u0_out1_9, u0_out3_13, u0_out3_16, 
      u0_out3_17, u0_out3_18, u0_out3_2, u0_out3_23, u0_out3_24, u0_out3_28, u0_out3_30, u0_out3_31, u0_out3_6, 
      u0_out3_9, u0_out5_1, u0_out5_10, u0_out5_13, u0_out5_14, u0_out5_16, u0_out5_18, u0_out5_2, u0_out5_20, 
      u0_out5_24, u0_out5_25, u0_out5_26, u0_out5_28, u0_out5_3, u0_out5_30, u0_out5_6, u0_out5_8, u0_out7_1, 
      u0_out7_10, u0_out7_11, u0_out7_14, u0_out7_15, u0_out7_19, u0_out7_20, u0_out7_21, u0_out7_25, u0_out7_26, 
      u0_out7_27, u0_out7_29, u0_out7_3, u0_out7_4, u0_out7_5, u0_out7_8, u0_uk_n110, u0_uk_n147, u0_uk_n155, 
      u0_uk_n164, u0_uk_n17, u0_uk_n207, u0_uk_n222, u0_uk_n230, u0_uk_n231, u0_uk_n238, u0_uk_n250, u0_uk_n252, 
      u0_uk_n31, u0_uk_n60, u0_uk_n687, u0_uk_n707, u1_out0_1, u1_out0_10, u1_out0_17, u1_out0_20, u1_out0_23, 
      u1_out0_26, u1_out0_31, u1_out0_9, u1_out10_13, u1_out10_16, u1_out10_18, u1_out10_2, u1_out10_24, u1_out10_28, 
      u1_out10_30, u1_out10_6, u1_out11_13, u1_out11_16, u1_out11_17, u1_out11_18, u1_out11_2, u1_out11_23, u1_out11_24, 
      u1_out11_28, u1_out11_30, u1_out11_31, u1_out11_6, u1_out11_9, u1_out12_1, u1_out12_10, u1_out12_14, u1_out12_15, 
      u1_out12_17, u1_out12_20, u1_out12_21, u1_out12_23, u1_out12_25, u1_out12_26, u1_out12_27, u1_out12_3, u1_out12_31, 
      u1_out12_5, u1_out12_8, u1_out12_9, u1_out14_1, u1_out14_10, u1_out14_16, u1_out14_20, u1_out14_24, u1_out14_26, 
      u1_out14_30, u1_out14_6, u1_out15_13, u1_out15_17, u1_out15_18, u1_out15_2, u1_out15_23, u1_out15_28, u1_out15_31, 
      u1_out15_9, u1_out1_11, u1_out1_19, u1_out1_29, u1_out1_4, u1_out2_13, u1_out2_17, u1_out2_18, u1_out2_2, 
      u1_out2_23, u1_out2_28, u1_out2_31, u1_out2_9, u1_out3_15, u1_out3_21, u1_out3_27, u1_out3_5, u1_out4_13, 
      u1_out4_18, u1_out4_2, u1_out4_28, u1_out5_1, u1_out5_10, u1_out5_11, u1_out5_12, u1_out5_13, u1_out5_15, 
      u1_out5_17, u1_out5_18, u1_out5_19, u1_out5_2, u1_out5_20, u1_out5_21, u1_out5_22, u1_out5_23, u1_out5_26, 
      u1_out5_27, u1_out5_28, u1_out5_29, u1_out5_31, u1_out5_32, u1_out5_4, u1_out5_5, u1_out5_7, u1_out5_9, 
      u1_out7_15, u1_out7_21, u1_out7_27, u1_out7_5, u1_out8_13, u1_out8_18, u1_out8_2, u1_out8_28, u1_out9_1, 
      u1_out9_10, u1_out9_15, u1_out9_16, u1_out9_20, u1_out9_21, u1_out9_24, u1_out9_26, u1_out9_27, u1_out9_30, 
      u1_out9_5, u1_out9_6, u2_out0_11, u2_out0_12, u2_out0_14, u2_out0_15, u2_out0_19, u2_out0_21, u2_out0_22, 
      u2_out0_25, u2_out0_27, u2_out0_29, u2_out0_3, u2_out0_32, u2_out0_4, u2_out0_5, u2_out0_7, u2_out0_8, 
      u2_out14_11, u2_out14_14, u2_out14_19, u2_out14_25, u2_out14_29, u2_out14_3, u2_out14_4, u2_out14_8, u2_out9_11, 
      u2_out9_19, u2_out9_29, u2_out9_4, u2_uk_n1142, u2_uk_n1152, u2_uk_n1171, u2_uk_n1178 );
endmodule
