module aes_aes_die_8 ( sa01_0, sa01_1, sa01_2, sa01_3, sa01_4, sa01_5, sa01_6, sa01_7, sa01_sr_0, sa01_sr_1, sa01_sr_2, sa01_sr_3, sa01_sr_4, sa01_sr_5, sa01_sr_6, sa01_sr_7 );
  input sa01_0, sa01_1, sa01_2, sa01_3, sa01_4, sa01_5, sa01_6, sa01_7;
  output sa01_sr_0, sa01_sr_1, sa01_sr_2, sa01_sr_3, sa01_sr_4, sa01_sr_5, sa01_sr_6, sa01_sr_7;
  wire us01_n438, us01_n439, us01_n440, us01_n441, us01_n442, us01_n443, us01_n444, us01_n445, us01_n446, 
       us01_n447, us01_n448, us01_n449, us01_n450, us01_n451, us01_n452, us01_n453, us01_n454, us01_n455, 
       us01_n456, us01_n457, us01_n458, us01_n459, us01_n460, us01_n461, us01_n462, us01_n463, us01_n464, 
       us01_n465, us01_n466, us01_n467, us01_n468, us01_n469, us01_n470, us01_n471, us01_n472, us01_n473, 
       us01_n474, us01_n475, us01_n476, us01_n477, us01_n478, us01_n479, us01_n480, us01_n481, us01_n482, 
       us01_n483, us01_n484, us01_n485, us01_n486, us01_n487, us01_n488, us01_n489, us01_n490, us01_n491, 
       us01_n492, us01_n493, us01_n494, us01_n495, us01_n496, us01_n497, us01_n498, us01_n499, us01_n500, 
       us01_n501, us01_n502, us01_n503, us01_n504, us01_n505, us01_n506, us01_n507, us01_n508, us01_n509, 
       us01_n510, us01_n511, us01_n512, us01_n513, us01_n514, us01_n515, us01_n516, us01_n517, us01_n518, 
       us01_n519, us01_n520, us01_n521, us01_n522, us01_n523, us01_n524, us01_n525, us01_n526, us01_n527, 
       us01_n528, us01_n529, us01_n530, us01_n531, us01_n532, us01_n533, us01_n534, us01_n535, us01_n536, 
       us01_n537, us01_n538, us01_n539, us01_n540, us01_n541, us01_n542, us01_n543, us01_n544, us01_n545, 
       us01_n546, us01_n547, us01_n548, us01_n549, us01_n550, us01_n551, us01_n552, us01_n553, us01_n554, 
       us01_n555, us01_n556, us01_n557, us01_n558, us01_n559, us01_n560, us01_n561, us01_n562, us01_n563, 
       us01_n564, us01_n565, us01_n566, us01_n567, us01_n568, us01_n569, us01_n570, us01_n571, us01_n572, 
       us01_n573, us01_n574, us01_n575, us01_n576, us01_n577, us01_n578, us01_n579, us01_n580, us01_n581, 
       us01_n582, us01_n583, us01_n584, us01_n585, us01_n586, us01_n587, us01_n588, us01_n589, us01_n590, 
       us01_n591, us01_n592, us01_n593, us01_n594, us01_n595, us01_n596, us01_n597, us01_n598, us01_n599, 
       us01_n600, us01_n601, us01_n602, us01_n603, us01_n604, us01_n605, us01_n606, us01_n607, us01_n608, 
       us01_n609, us01_n610, us01_n611, us01_n612, us01_n613, us01_n614, us01_n615, us01_n616, us01_n617, 
       us01_n618, us01_n619, us01_n620, us01_n621, us01_n622, us01_n623, us01_n624, us01_n625, us01_n626, 
       us01_n627, us01_n628, us01_n629, us01_n630, us01_n631, us01_n632, us01_n633, us01_n634, us01_n635, 
       us01_n636, us01_n637, us01_n638, us01_n639, us01_n640, us01_n641, us01_n642, us01_n643, us01_n644, 
       us01_n645, us01_n646, us01_n647, us01_n648, us01_n649, us01_n650, us01_n651, us01_n652, us01_n653, 
       us01_n654, us01_n655, us01_n656, us01_n657, us01_n658, us01_n659, us01_n660, us01_n661, us01_n662, 
       us01_n663, us01_n664, us01_n665, us01_n666, us01_n667, us01_n668, us01_n669, us01_n670, us01_n671, 
       us01_n672, us01_n673, us01_n674, us01_n675, us01_n676, us01_n677, us01_n678, us01_n679, us01_n680, 
       us01_n681, us01_n682, us01_n683, us01_n684, us01_n685, us01_n686, us01_n687, us01_n688, us01_n689, 
       us01_n690, us01_n691, us01_n692, us01_n693, us01_n694, us01_n695, us01_n696, us01_n697, us01_n698, 
       us01_n699, us01_n700, us01_n701, us01_n702, us01_n703, us01_n704, us01_n705, us01_n706, us01_n707, 
       us01_n708, us01_n709, us01_n710, us01_n711, us01_n712, us01_n713, us01_n714, us01_n715, us01_n716, 
       us01_n717, us01_n718, us01_n719, us01_n720, us01_n721, us01_n722, us01_n723, us01_n724, us01_n725, 
       us01_n726, us01_n727, us01_n728, us01_n729, us01_n730, us01_n731, us01_n732, us01_n733, us01_n734, 
       us01_n735, us01_n736, us01_n737, us01_n738, us01_n739, us01_n740, us01_n741, us01_n742, us01_n743, 
       us01_n744, us01_n745, us01_n746, us01_n747, us01_n748, us01_n749, us01_n750, us01_n751, us01_n752, 
       us01_n753, us01_n754, us01_n755, us01_n756, us01_n757, us01_n758, us01_n759, us01_n760, us01_n761, 
       us01_n762, us01_n763, us01_n764, us01_n765, us01_n766, us01_n767, us01_n768, us01_n769, us01_n770, 
       us01_n771, us01_n772, us01_n773, us01_n774, us01_n775, us01_n776, us01_n777, us01_n778, us01_n779, 
       us01_n780, us01_n781, us01_n782, us01_n783, us01_n784, us01_n785, us01_n786, us01_n787, us01_n788, 
       us01_n789, us01_n790, us01_n791, us01_n792, us01_n793, us01_n794, us01_n795, us01_n796, us01_n797, 
       us01_n798, us01_n799, us01_n800, us01_n801, us01_n802, us01_n803, us01_n804, us01_n805, us01_n806, 
       us01_n807, us01_n808, us01_n809, us01_n810, us01_n811, us01_n812, us01_n813, us01_n814, us01_n815, 
       us01_n816, us01_n817, us01_n818, us01_n819, us01_n820, us01_n821, us01_n822, us01_n823, us01_n824, 
       us01_n825, us01_n826, us01_n827, us01_n828, us01_n829, us01_n830, us01_n831, us01_n832, us01_n833, 
       us01_n834, us01_n835, us01_n836, us01_n837, us01_n838, us01_n839, us01_n840, us01_n841, us01_n842, 
       us01_n843, us01_n844, us01_n845, us01_n846, us01_n847, us01_n848, us01_n849, us01_n850, us01_n851, 
       us01_n852, us01_n853, us01_n854, us01_n855, us01_n856, us01_n857, us01_n858, us01_n859, us01_n860, 
       us01_n861, us01_n862, us01_n863, us01_n864, us01_n865, us01_n866, us01_n867, us01_n868, us01_n869, 
       us01_n870, us01_n871, us01_n872, us01_n873,  us01_n874;
  NOR2_X1 us01_U10 (.ZN( us01_n573 ) , .A1( us01_n620 ) , .A2( us01_n743 ) );
  AOI211_X1 us01_U100 (.B( us01_n537 ) , .A( us01_n538 ) , .ZN( us01_n549 ) , .C2( us01_n837 ) , .C1( us01_n849 ) );
  NOR4_X1 us01_U101 (.A4( us01_n542 ) , .A3( us01_n543 ) , .A2( us01_n544 ) , .A1( us01_n545 ) , .ZN( us01_n546 ) );
  NOR4_X1 us01_U102 (.A4( us01_n607 ) , .A3( us01_n608 ) , .A2( us01_n609 ) , .A1( us01_n610 ) , .ZN( us01_n617 ) );
  NOR4_X1 us01_U103 (.ZN( us01_n618 ) , .A1( us01_n654 ) , .A3( us01_n664 ) , .A4( us01_n680 ) , .A2( us01_n764 ) );
  NOR4_X1 us01_U104 (.A4( us01_n612 ) , .A3( us01_n613 ) , .A2( us01_n614 ) , .A1( us01_n615 ) , .ZN( us01_n616 ) );
  NOR2_X1 us01_U105 (.ZN( us01_n684 ) , .A1( us01_n829 ) , .A2( us01_n830 ) );
  NAND4_X1 us01_U106 (.A4( us01_n471 ) , .A3( us01_n472 ) , .A2( us01_n473 ) , .A1( us01_n474 ) , .ZN( us01_n676 ) );
  NOR4_X1 us01_U107 (.A4( us01_n468 ) , .ZN( us01_n474 ) , .A3( us01_n554 ) , .A1( us01_n733 ) , .A2( us01_n753 ) );
  NOR4_X1 us01_U108 (.ZN( us01_n473 ) , .A1( us01_n529 ) , .A3( us01_n566 ) , .A4( us01_n598 ) , .A2( us01_n640 ) );
  NOR4_X1 us01_U109 (.ZN( us01_n472 ) , .A1( us01_n504 ) , .A3( us01_n542 ) , .A2( us01_n581 ) , .A4( us01_n714 ) );
  NOR2_X1 us01_U11 (.ZN( us01_n493 ) , .A1( us01_n676 ) , .A2( us01_n692 ) );
  NAND4_X1 us01_U110 (.A4( us01_n689 ) , .A3( us01_n690 ) , .A1( us01_n691 ) , .ZN( us01_n774 ) , .A2( us01_n870 ) );
  INV_X1 us01_U111 (.A( us01_n677 ) , .ZN( us01_n870 ) );
  AOI221_X1 us01_U112 (.A( us01_n679 ) , .ZN( us01_n690 ) , .B2( us01_n838 ) , .C1( us01_n840 ) , .C2( us01_n860 ) , .B1( us01_n863 ) );
  NOR4_X1 us01_U113 (.A4( us01_n685 ) , .A3( us01_n686 ) , .A2( us01_n687 ) , .A1( us01_n688 ) , .ZN( us01_n689 ) );
  NOR2_X1 us01_U114 (.ZN( us01_n731 ) , .A2( us01_n830 ) , .A1( us01_n843 ) );
  NAND4_X1 us01_U115 (.A4( us01_n717 ) , .A3( us01_n718 ) , .A2( us01_n719 ) , .ZN( us01_n739 ) , .A1( us01_n855 ) );
  AOI221_X1 us01_U116 (.A( us01_n708 ) , .ZN( us01_n719 ) , .C2( us01_n842 ) , .B2( us01_n843 ) , .C1( us01_n859 ) , .B1( us01_n860 ) );
  INV_X1 us01_U117 (.A( us01_n707 ) , .ZN( us01_n855 ) );
  NOR4_X1 us01_U118 (.A4( us01_n713 ) , .A3( us01_n714 ) , .A2( us01_n715 ) , .A1( us01_n716 ) , .ZN( us01_n717 ) );
  NOR2_X1 us01_U119 (.ZN( us01_n645 ) , .A1( us01_n852 ) , .A2( us01_n866 ) );
  NOR2_X1 us01_U12 (.A1( us01_n676 ) , .ZN( us01_n691 ) , .A2( us01_n805 ) );
  NAND4_X1 us01_U120 (.A4( us01_n571 ) , .A3( us01_n572 ) , .A1( us01_n573 ) , .ZN( us01_n721 ) , .A2( us01_n872 ) );
  AOI221_X1 us01_U121 (.A( us01_n562 ) , .C2( us01_n563 ) , .ZN( us01_n572 ) , .B2( us01_n843 ) , .B1( us01_n850 ) , .C1( us01_n851 ) );
  NOR4_X1 us01_U122 (.A4( us01_n567 ) , .A3( us01_n568 ) , .A2( us01_n569 ) , .A1( us01_n570 ) , .ZN( us01_n571 ) );
  INV_X1 us01_U123 (.A( us01_n605 ) , .ZN( us01_n872 ) );
  NAND4_X1 us01_U124 (.A4( us01_n491 ) , .A3( us01_n492 ) , .A1( us01_n493 ) , .ZN( us01_n800 ) , .A2( us01_n865 ) );
  AOI221_X1 us01_U125 (.A( us01_n487 ) , .ZN( us01_n492 ) , .B2( us01_n834 ) , .C2( us01_n839 ) , .C1( us01_n849 ) , .B1( us01_n858 ) );
  INV_X1 us01_U126 (.A( us01_n776 ) , .ZN( us01_n865 ) );
  NOR4_X1 us01_U127 (.A2( us01_n489 ) , .A1( us01_n490 ) , .ZN( us01_n491 ) , .A3( us01_n578 ) , .A4( us01_n610 ) );
  NOR4_X1 us01_U128 (.A3( us01_n753 ) , .A2( us01_n754 ) , .A1( us01_n755 ) , .ZN( us01_n756 ) , .A4( us01_n867 ) );
  AOI211_X1 us01_U129 (.B( us01_n743 ) , .A( us01_n744 ) , .ZN( us01_n757 ) , .C1( us01_n830 ) , .C2( us01_n851 ) );
  NOR3_X1 us01_U13 (.ZN( us01_n502 ) , .A2( us01_n677 ) , .A3( us01_n775 ) , .A1( us01_n874 ) );
  NOR3_X1 us01_U130 (.A3( us01_n739 ) , .A2( us01_n740 ) , .A1( us01_n741 ) , .ZN( us01_n758 ) );
  NOR4_X1 us01_U131 (.A4( us01_n732 ) , .A3( us01_n733 ) , .A2( us01_n734 ) , .A1( us01_n735 ) , .ZN( us01_n736 ) );
  AOI211_X1 us01_U132 (.B( us01_n723 ) , .A( us01_n724 ) , .ZN( us01_n737 ) , .C1( us01_n841 ) , .C2( us01_n853 ) );
  NOR3_X1 us01_U133 (.A3( us01_n720 ) , .A1( us01_n721 ) , .ZN( us01_n738 ) , .A2( us01_n739 ) );
  INV_X1 us01_U134 (.A( us01_n760 ) , .ZN( us01_n828 ) );
  NAND4_X1 us01_U135 (.ZN( sa01_sr_3 ) , .A4( us01_n702 ) , .A3( us01_n703 ) , .A2( us01_n704 ) , .A1( us01_n705 ) );
  NOR4_X1 us01_U136 (.A4( us01_n698 ) , .A3( us01_n699 ) , .A2( us01_n700 ) , .A1( us01_n701 ) , .ZN( us01_n702 ) );
  AOI211_X1 us01_U137 (.B( us01_n692 ) , .A( us01_n693 ) , .ZN( us01_n703 ) , .C2( us01_n829 ) , .C1( us01_n849 ) );
  NOR2_X1 us01_U138 (.ZN( us01_n705 ) , .A2( us01_n774 ) , .A1( us01_n798 ) );
  OR4_X1 us01_U139 (.A4( us01_n680 ) , .A3( us01_n681 ) , .A2( us01_n682 ) , .A1( us01_n683 ) , .ZN( us01_n688 ) );
  INV_X1 us01_U14 (.A( us01_n704 ) , .ZN( us01_n874 ) );
  OR4_X1 us01_U140 (.ZN( us01_n464 ) , .A4( us01_n516 ) , .A3( us01_n527 ) , .A2( us01_n576 ) , .A1( us01_n710 ) );
  OR4_X1 us01_U141 (.A4( us01_n564 ) , .A3( us01_n565 ) , .A2( us01_n566 ) , .ZN( us01_n570 ) , .A1( us01_n663 ) );
  OR4_X1 us01_U142 (.A4( us01_n516 ) , .A2( us01_n517 ) , .A1( us01_n518 ) , .ZN( us01_n520 ) , .A3( us01_n819 ) );
  OR4_X1 us01_U143 (.ZN( us01_n490 ) , .A4( us01_n532 ) , .A2( us01_n545 ) , .A1( us01_n557 ) , .A3( us01_n630 ) );
  OR4_X1 us01_U144 (.A4( us01_n578 ) , .A3( us01_n579 ) , .A2( us01_n580 ) , .A1( us01_n581 ) , .ZN( us01_n582 ) );
  INV_X1 us01_U145 (.A( us01_n695 ) , .ZN( us01_n836 ) );
  NAND2_X1 us01_U146 (.ZN( us01_n611 ) , .A2( us01_n835 ) , .A1( us01_n871 ) );
  OR3_X1 us01_U147 (.A3( us01_n504 ) , .A2( us01_n505 ) , .A1( us01_n506 ) , .ZN( us01_n509 ) );
  AOI221_X1 us01_U148 (.A( us01_n711 ) , .B2( us01_n712 ) , .ZN( us01_n718 ) , .C1( us01_n830 ) , .B1( us01_n837 ) , .C2( us01_n861 ) );
  OR2_X1 us01_U149 (.A2( us01_n709 ) , .A1( us01_n710 ) , .ZN( us01_n711 ) );
  INV_X1 us01_U15 (.A( us01_n678 ) , .ZN( us01_n838 ) );
  INV_X1 us01_U150 (.A( us01_n461 ) , .ZN( us01_n862 ) );
  OAI21_X1 us01_U151 (.ZN( us01_n461 ) , .B1( us01_n807 ) , .A( us01_n832 ) , .B2( us01_n849 ) );
  INV_X1 us01_U152 (.A( us01_n752 ) , .ZN( us01_n867 ) );
  OAI21_X1 us01_U153 (.B1( us01_n751 ) , .ZN( us01_n752 ) , .A( us01_n843 ) , .B2( us01_n866 ) );
  INV_X1 us01_U154 (.A( us01_n670 ) , .ZN( us01_n857 ) );
  AOI21_X1 us01_U155 (.A( us01_n668 ) , .B1( us01_n669 ) , .ZN( us01_n670 ) , .B2( us01_n854 ) );
  AOI222_X1 us01_U156 (.ZN( us01_n658 ) , .A2( us01_n837 ) , .B1( us01_n839 ) , .C2( us01_n843 ) , .A1( us01_n858 ) , .C1( us01_n861 ) , .B2( us01_n868 ) );
  INV_X1 us01_U157 (.A( us01_n645 ) , .ZN( us01_n868 ) );
  OAI22_X1 us01_U158 (.ZN( us01_n481 ) , .A1( us01_n706 ) , .B2( us01_n783 ) , .A2( us01_n804 ) , .B1( us01_n810 ) );
  OAI22_X1 us01_U159 (.ZN( us01_n635 ) , .A1( us01_n697 ) , .B2( us01_n726 ) , .A2( us01_n760 ) , .B1( us01_n814 ) );
  NOR4_X1 us01_U16 (.A4( us01_n443 ) , .A3( us01_n444 ) , .A2( us01_n514 ) , .A1( us01_n539 ) , .ZN( us01_n704 ) );
  OAI222_X1 us01_U160 (.ZN( us01_n503 ) , .C2( us01_n623 ) , .B2( us01_n645 ) , .B1( us01_n745 ) , .A2( us01_n746 ) , .C1( us01_n803 ) , .A1( us01_n804 ) );
  OAI222_X1 us01_U161 (.B2( us01_n745 ) , .B1( us01_n746 ) , .A2( us01_n747 ) , .ZN( us01_n755 ) , .C2( us01_n803 ) , .C1( us01_n812 ) , .A1( us01_n815 ) );
  OAI222_X1 us01_U162 (.B2( us01_n706 ) , .ZN( us01_n707 ) , .C2( us01_n722 ) , .B1( us01_n745 ) , .A1( us01_n804 ) , .C1( us01_n812 ) , .A2( us01_n813 ) );
  AOI22_X1 us01_U163 (.ZN( us01_n694 ) , .A1( us01_n828 ) , .B2( us01_n841 ) , .A2( us01_n863 ) , .B1( us01_n866 ) );
  AOI22_X1 us01_U164 (.A2( us01_n780 ) , .ZN( us01_n781 ) , .B2( us01_n829 ) , .A1( us01_n832 ) , .B1( us01_n861 ) );
  INV_X1 us01_U165 (.A( us01_n728 ) , .ZN( us01_n837 ) );
  AOI221_X1 us01_U166 (.A( us01_n762 ) , .ZN( us01_n772 ) , .C2( us01_n808 ) , .B2( us01_n833 ) , .C1( us01_n853 ) , .B1( us01_n864 ) );
  AOI21_X1 us01_U167 (.B2( us01_n761 ) , .ZN( us01_n762 ) , .A( us01_n786 ) , .B1( us01_n790 ) );
  INV_X1 us01_U168 (.A( us01_n759 ) , .ZN( us01_n833 ) );
  INV_X1 us01_U169 (.A( us01_n788 ) , .ZN( us01_n830 ) );
  OR3_X1 us01_U17 (.ZN( us01_n444 ) , .A1( us01_n526 ) , .A3( us01_n575 ) , .A2( us01_n873 ) );
  OAI221_X1 us01_U170 (.A( us01_n725 ) , .C2( us01_n726 ) , .B2( us01_n727 ) , .B1( us01_n728 ) , .ZN( us01_n735 ) , .C1( us01_n815 ) );
  AOI22_X1 us01_U171 (.ZN( us01_n725 ) , .B1( us01_n830 ) , .A2( us01_n836 ) , .A1( us01_n861 ) , .B2( us01_n864 ) );
  NAND2_X1 us01_U172 (.A1( us01_n449 ) , .A2( us01_n451 ) , .ZN( us01_n760 ) );
  OAI22_X1 us01_U173 (.ZN( us01_n622 ) , .B1( us01_n667 ) , .B2( us01_n745 ) , .A1( us01_n813 ) , .A2( us01_n814 ) );
  OAI22_X1 us01_U174 (.A1( us01_n722 ) , .ZN( us01_n724 ) , .B2( us01_n748 ) , .B1( us01_n810 ) , .A2( us01_n814 ) );
  OAI22_X1 us01_U175 (.ZN( us01_n487 ) , .A1( us01_n722 ) , .B2( us01_n726 ) , .B1( us01_n728 ) , .A2( us01_n777 ) );
  OAI22_X1 us01_U176 (.B2( us01_n777 ) , .B1( us01_n778 ) , .ZN( us01_n779 ) , .A2( us01_n812 ) , .A1( us01_n813 ) );
  OAI22_X1 us01_U177 (.B2( us01_n748 ) , .B1( us01_n749 ) , .A1( us01_n750 ) , .ZN( us01_n754 ) , .A2( us01_n804 ) );
  NOR3_X1 us01_U178 (.ZN( us01_n750 ) , .A2( us01_n851 ) , .A1( us01_n861 ) , .A3( us01_n863 ) );
  NOR2_X1 us01_U179 (.ZN( us01_n749 ) , .A2( us01_n850 ) , .A1( us01_n858 ) );
  OR4_X1 us01_U18 (.A4( us01_n440 ) , .A2( us01_n441 ) , .A1( us01_n442 ) , .ZN( us01_n443 ) , .A3( us01_n551 ) );
  INV_X1 us01_U180 (.A( us01_n803 ) , .ZN( us01_n858 ) );
  OAI22_X1 us01_U181 (.B2( us01_n742 ) , .ZN( us01_n744 ) , .A2( us01_n760 ) , .B1( us01_n778 ) , .A1( us01_n790 ) );
  OAI22_X1 us01_U182 (.ZN( us01_n494 ) , .A2( us01_n742 ) , .A1( us01_n778 ) , .B1( us01_n789 ) , .B2( us01_n804 ) );
  OAI22_X1 us01_U183 (.B2( us01_n801 ) , .B1( us01_n802 ) , .A2( us01_n803 ) , .A1( us01_n804 ) , .ZN( us01_n806 ) );
  OAI22_X1 us01_U184 (.ZN( us01_n693 ) , .A2( us01_n728 ) , .A1( us01_n778 ) , .B1( us01_n789 ) , .B2( us01_n815 ) );
  NOR2_X1 us01_U185 (.ZN( us01_n713 ) , .A1( us01_n803 ) , .A2( us01_n815 ) );
  NOR2_X1 us01_U186 (.A1( us01_n697 ) , .ZN( us01_n766 ) , .A2( us01_n811 ) );
  INV_X1 us01_U187 (.A( us01_n786 ) , .ZN( us01_n843 ) );
  NOR2_X1 us01_U188 (.ZN( us01_n539 ) , .A2( us01_n695 ) , .A1( us01_n697 ) );
  INV_X1 us01_U189 (.A( us01_n742 ) , .ZN( us01_n835 ) );
  INV_X1 us01_U19 (.A( us01_n611 ) , .ZN( us01_n873 ) );
  INV_X1 us01_U190 (.A( us01_n814 ) , .ZN( us01_n829 ) );
  INV_X1 us01_U191 (.A( us01_n812 ) , .ZN( us01_n831 ) );
  OAI22_X1 us01_U192 (.B1( us01_n488 ) , .ZN( us01_n489 ) , .A1( us01_n684 ) , .A2( us01_n761 ) , .B2( us01_n815 ) );
  NOR3_X1 us01_U193 (.ZN( us01_n488 ) , .A1( us01_n780 ) , .A2( us01_n848 ) , .A3( us01_n861 ) );
  NOR2_X1 us01_U194 (.A2( us01_n742 ) , .ZN( us01_n753 ) , .A1( us01_n803 ) );
  NOR2_X1 us01_U195 (.ZN( us01_n733 ) , .A2( us01_n801 ) , .A1( us01_n803 ) );
  INV_X1 us01_U196 (.A( us01_n790 ) , .ZN( us01_n849 ) );
  NOR2_X1 us01_U197 (.A2( us01_n742 ) , .ZN( us01_n767 ) , .A1( us01_n810 ) );
  NOR2_X1 us01_U198 (.ZN( us01_n664 ) , .A1( us01_n726 ) , .A2( us01_n801 ) );
  OAI22_X1 us01_U199 (.ZN( us01_n708 ) , .A2( us01_n726 ) , .B2( us01_n727 ) , .A1( us01_n742 ) , .B1( us01_n811 ) );
  AOI222_X1 us01_U20 (.ZN( us01_n561 ) , .B1( us01_n828 ) , .C1( us01_n839 ) , .A2( us01_n841 ) , .A1( us01_n852 ) , .B2( us01_n861 ) , .C2( us01_n871 ) );
  NOR2_X1 us01_U200 (.ZN( us01_n650 ) , .A1( us01_n667 ) , .A2( us01_n812 ) );
  NOR2_X1 us01_U201 (.ZN( us01_n592 ) , .A2( us01_n695 ) , .A1( us01_n726 ) );
  NOR2_X1 us01_U202 (.A1( us01_n667 ) , .ZN( us01_n671 ) , .A2( us01_n742 ) );
  NOR2_X1 us01_U203 (.ZN( us01_n600 ) , .A1( us01_n667 ) , .A2( us01_n801 ) );
  NOR2_X1 us01_U204 (.A1( us01_n667 ) , .ZN( us01_n686 ) , .A2( us01_n814 ) );
  NOR2_X1 us01_U205 (.ZN( us01_n568 ) , .A1( us01_n726 ) , .A2( us01_n804 ) );
  NOR2_X1 us01_U206 (.A1( us01_n667 ) , .ZN( us01_n764 ) , .A2( us01_n811 ) );
  NOR2_X1 us01_U207 (.ZN( us01_n525 ) , .A1( us01_n667 ) , .A2( us01_n777 ) );
  NOR2_X1 us01_U208 (.ZN( us01_n652 ) , .A1( us01_n726 ) , .A2( us01_n811 ) );
  NOR2_X1 us01_U209 (.ZN( us01_n505 ) , .A1( us01_n810 ) , .A2( us01_n815 ) );
  NOR4_X1 us01_U21 (.ZN( us01_n471 ) , .A2( us01_n519 ) , .A4( us01_n592 ) , .A1( us01_n607 ) , .A3( us01_n627 ) );
  NOR2_X1 us01_U210 (.ZN( us01_n659 ) , .A1( us01_n727 ) , .A2( us01_n788 ) );
  NOR2_X1 us01_U211 (.ZN( us01_n544 ) , .A2( us01_n778 ) , .A1( us01_n812 ) );
  NOR2_X1 us01_U212 (.ZN( us01_n575 ) , .A2( us01_n697 ) , .A1( us01_n812 ) );
  NOR2_X1 us01_U213 (.ZN( us01_n507 ) , .A1( us01_n727 ) , .A2( us01_n777 ) );
  NOR2_X1 us01_U214 (.ZN( us01_n716 ) , .A2( us01_n722 ) , .A1( us01_n742 ) );
  INV_X1 us01_U215 (.A( us01_n748 ) , .ZN( us01_n840 ) );
  NOR2_X1 us01_U216 (.ZN( us01_n530 ) , .A2( us01_n747 ) , .A1( us01_n748 ) );
  NOR2_X1 us01_U217 (.ZN( us01_n660 ) , .A2( us01_n695 ) , .A1( us01_n727 ) );
  NOR2_X1 us01_U218 (.ZN( us01_n613 ) , .A1( us01_n783 ) , .A2( us01_n813 ) );
  NOR2_X1 us01_U219 (.ZN( us01_n627 ) , .A2( us01_n726 ) , .A1( us01_n783 ) );
  NOR4_X1 us01_U22 (.ZN( us01_n477 ) , .A1( us01_n518 ) , .A4( us01_n555 ) , .A3( us01_n580 ) , .A2( us01_n628 ) );
  NOR2_X1 us01_U220 (.ZN( us01_n609 ) , .A2( us01_n778 ) , .A1( us01_n804 ) );
  NOR2_X1 us01_U221 (.ZN( us01_n661 ) , .A1( us01_n727 ) , .A2( us01_n783 ) );
  NOR2_X1 us01_U222 (.ZN( us01_n626 ) , .A2( us01_n667 ) , .A1( us01_n783 ) );
  NOR2_X1 us01_U223 (.ZN( us01_n599 ) , .A2( us01_n778 ) , .A1( us01_n801 ) );
  INV_X1 us01_U224 (.A( us01_n745 ) , .ZN( us01_n832 ) );
  NOR2_X1 us01_U225 (.ZN( us01_n554 ) , .A1( us01_n760 ) , .A2( us01_n803 ) );
  NOR2_X1 us01_U226 (.ZN( us01_n529 ) , .A2( us01_n778 ) , .A1( us01_n814 ) );
  NOR2_X1 us01_U227 (.ZN( us01_n526 ) , .A2( us01_n722 ) , .A1( us01_n801 ) );
  NOR2_X1 us01_U228 (.A2( us01_n706 ) , .A1( us01_n748 ) , .ZN( us01_n769 ) );
  NOR2_X1 us01_U229 (.ZN( us01_n597 ) , .A2( us01_n789 ) , .A1( us01_n814 ) );
  NOR4_X1 us01_U23 (.ZN( us01_n454 ) , .A2( us01_n515 ) , .A1( us01_n541 ) , .A3( us01_n577 ) , .A4( us01_n613 ) );
  NOR2_X1 us01_U230 (.ZN( us01_n555 ) , .A1( us01_n790 ) , .A2( us01_n812 ) );
  NOR2_X1 us01_U231 (.ZN( us01_n542 ) , .A2( us01_n783 ) , .A1( us01_n790 ) );
  NOR2_X1 us01_U232 (.A2( us01_n695 ) , .ZN( us01_n714 ) , .A1( us01_n790 ) );
  NOR2_X1 us01_U233 (.ZN( us01_n665 ) , .A1( us01_n748 ) , .A2( us01_n813 ) );
  NOR2_X1 us01_U234 (.ZN( us01_n543 ) , .A1( us01_n747 ) , .A2( us01_n812 ) );
  NOR2_X1 us01_U235 (.ZN( us01_n553 ) , .A1( us01_n748 ) , .A2( us01_n789 ) );
  NOR2_X1 us01_U236 (.ZN( us01_n506 ) , .A2( us01_n778 ) , .A1( us01_n783 ) );
  NOR2_X1 us01_U237 (.ZN( us01_n541 ) , .A2( us01_n706 ) , .A1( us01_n783 ) );
  NOR2_X1 us01_U238 (.ZN( us01_n514 ) , .A1( us01_n706 ) , .A2( us01_n742 ) );
  NOR2_X1 us01_U239 (.ZN( us01_n662 ) , .A1( us01_n783 ) , .A2( us01_n789 ) );
  NOR4_X1 us01_U24 (.A4( us01_n530 ) , .A3( us01_n531 ) , .A2( us01_n532 ) , .ZN( us01_n533 ) , .A1( us01_n818 ) );
  NOR2_X1 us01_U240 (.ZN( us01_n556 ) , .A1( us01_n706 ) , .A2( us01_n814 ) );
  NOR2_X1 us01_U241 (.ZN( us01_n515 ) , .A1( us01_n706 ) , .A2( us01_n801 ) );
  NOR2_X1 us01_U242 (.ZN( us01_n612 ) , .A1( us01_n760 ) , .A2( us01_n810 ) );
  NOR2_X1 us01_U243 (.ZN( us01_n629 ) , .A1( us01_n722 ) , .A2( us01_n811 ) );
  NOR2_X1 us01_U244 (.A1( us01_n747 ) , .ZN( us01_n765 ) , .A2( us01_n801 ) );
  NOR2_X1 us01_U245 (.ZN( us01_n528 ) , .A2( us01_n742 ) , .A1( us01_n790 ) );
  INV_X1 us01_U246 (.A( us01_n804 ) , .ZN( us01_n839 ) );
  OAI22_X1 us01_U247 (.B1( us01_n438 ) , .ZN( us01_n442 ) , .A2( us01_n726 ) , .A1( us01_n742 ) , .B2( us01_n747 ) );
  NOR3_X1 us01_U248 (.ZN( us01_n438 ) , .A2( us01_n834 ) , .A3( us01_n835 ) , .A1( us01_n844 ) );
  INV_X1 us01_U249 (.A( us01_n726 ) , .ZN( us01_n850 ) );
  NOR4_X1 us01_U25 (.A4( us01_n539 ) , .A3( us01_n540 ) , .A2( us01_n541 ) , .ZN( us01_n548 ) , .A1( us01_n686 ) );
  NOR2_X1 us01_U250 (.ZN( us01_n519 ) , .A1( us01_n788 ) , .A2( us01_n810 ) );
  NOR2_X1 us01_U251 (.ZN( us01_n668 ) , .A1( us01_n788 ) , .A2( us01_n803 ) );
  AOI21_X1 us01_U252 (.ZN( us01_n550 ) , .B1( us01_n667 ) , .A( us01_n695 ) , .B2( us01_n803 ) );
  AOI21_X1 us01_U253 (.ZN( us01_n587 ) , .B2( us01_n697 ) , .B1( us01_n813 ) , .A( us01_n815 ) );
  NOR2_X1 us01_U254 (.ZN( us01_n504 ) , .A2( us01_n726 ) , .A1( us01_n760 ) );
  NOR2_X1 us01_U255 (.ZN( us01_n653 ) , .A1( us01_n788 ) , .A2( us01_n813 ) );
  INV_X1 us01_U256 (.A( us01_n801 ) , .ZN( us01_n841 ) );
  NOR2_X1 us01_U257 (.ZN( us01_n628 ) , .A1( us01_n745 ) , .A2( us01_n813 ) );
  NOR2_X1 us01_U258 (.ZN( us01_n545 ) , .A1( us01_n697 ) , .A2( us01_n742 ) );
  INV_X1 us01_U259 (.A( us01_n697 ) , .ZN( us01_n851 ) );
  NOR2_X1 us01_U26 (.ZN( us01_n678 ) , .A2( us01_n832 ) , .A1( us01_n837 ) );
  NOR2_X1 us01_U260 (.ZN( us01_n640 ) , .A2( us01_n786 ) , .A1( us01_n789 ) );
  AOI21_X1 us01_U261 (.ZN( us01_n648 ) , .A( us01_n777 ) , .B1( us01_n790 ) , .B2( us01_n803 ) );
  NOR2_X1 us01_U262 (.ZN( us01_n666 ) , .A2( us01_n706 ) , .A1( us01_n788 ) );
  NOR2_X1 us01_U263 (.A2( us01_n695 ) , .A1( us01_n778 ) , .ZN( us01_n818 ) );
  NOR2_X1 us01_U264 (.A1( us01_n695 ) , .ZN( us01_n768 ) , .A2( us01_n813 ) );
  AOI21_X1 us01_U265 (.ZN( us01_n624 ) , .B2( us01_n667 ) , .A( us01_n788 ) , .B1( us01_n789 ) );
  NOR2_X1 us01_U266 (.ZN( us01_n577 ) , .A2( us01_n706 ) , .A1( us01_n728 ) );
  INV_X1 us01_U267 (.A( us01_n761 ) , .ZN( us01_n864 ) );
  NOR2_X1 us01_U268 (.A2( us01_n706 ) , .A1( us01_n760 ) , .ZN( us01_n792 ) );
  NOR2_X1 us01_U269 (.ZN( us01_n607 ) , .A2( us01_n722 ) , .A1( us01_n815 ) );
  AOI222_X1 us01_U27 (.ZN( us01_n467 ) , .B1( us01_n830 ) , .A1( us01_n837 ) , .C1( us01_n840 ) , .C2( us01_n849 ) , .A2( us01_n853 ) , .B2( us01_n863 ) );
  NOR2_X1 us01_U270 (.ZN( us01_n531 ) , .A2( us01_n722 ) , .A1( us01_n728 ) );
  AOI21_X1 us01_U271 (.ZN( us01_n508 ) , .B2( us01_n667 ) , .A( us01_n728 ) , .B1( us01_n813 ) );
  AOI21_X1 us01_U272 (.ZN( us01_n537 ) , .B2( us01_n810 ) , .A( us01_n812 ) , .B1( us01_n813 ) );
  INV_X1 us01_U273 (.A( us01_n727 ) , .ZN( us01_n866 ) );
  NOR2_X1 us01_U274 (.ZN( us01_n540 ) , .A1( us01_n760 ) , .A2( us01_n789 ) );
  INV_X1 us01_U275 (.A( us01_n810 ) , .ZN( us01_n852 ) );
  AOI21_X1 us01_U276 (.B1( us01_n697 ) , .ZN( us01_n698 ) , .A( us01_n730 ) , .B2( us01_n761 ) );
  NOR2_X1 us01_U277 (.ZN( us01_n579 ) , .A1( us01_n667 ) , .A2( us01_n786 ) );
  AOI21_X1 us01_U278 (.ZN( us01_n589 ) , .B2( us01_n761 ) , .A( us01_n783 ) , .B1( us01_n810 ) );
  NOR2_X1 us01_U279 (.ZN( us01_n654 ) , .A1( us01_n745 ) , .A2( us01_n778 ) );
  NOR4_X1 us01_U28 (.A1( us01_n464 ) , .ZN( us01_n465 ) , .A4( us01_n540 ) , .A2( us01_n552 ) , .A3( us01_n612 ) );
  INV_X1 us01_U280 (.A( us01_n789 ) , .ZN( us01_n871 ) );
  AOI21_X1 us01_U281 (.B1( us01_n623 ) , .ZN( us01_n625 ) , .A( us01_n761 ) , .B2( us01_n812 ) );
  NOR2_X1 us01_U282 (.ZN( us01_n683 ) , .A1( us01_n727 ) , .A2( us01_n814 ) );
  AOI21_X1 us01_U283 (.A( us01_n813 ) , .B2( us01_n814 ) , .B1( us01_n815 ) , .ZN( us01_n816 ) );
  AOI21_X1 us01_U284 (.ZN( us01_n647 ) , .B1( us01_n727 ) , .B2( us01_n761 ) , .A( us01_n811 ) );
  AOI21_X1 us01_U285 (.A( us01_n810 ) , .B2( us01_n811 ) , .B1( us01_n812 ) , .ZN( us01_n817 ) );
  AOI21_X1 us01_U286 (.ZN( us01_n513 ) , .A( us01_n727 ) , .B1( us01_n748 ) , .B2( us01_n801 ) );
  AOI21_X1 us01_U287 (.ZN( us01_n497 ) , .B1( us01_n678 ) , .A( us01_n810 ) , .B2( us01_n814 ) );
  NOR2_X1 us01_U288 (.ZN( us01_n518 ) , .A2( us01_n706 ) , .A1( us01_n812 ) );
  AOI21_X1 us01_U289 (.ZN( us01_n475 ) , .A( us01_n667 ) , .B1( us01_n748 ) , .B2( us01_n804 ) );
  AOI221_X1 us01_U29 (.ZN( us01_n466 ) , .C2( us01_n712 ) , .B2( us01_n829 ) , .C1( us01_n843 ) , .B1( us01_n858 ) , .A( us01_n862 ) );
  NOR2_X1 us01_U290 (.ZN( us01_n566 ) , .A1( us01_n727 ) , .A2( us01_n760 ) );
  NOR2_X1 us01_U291 (.ZN( us01_n580 ) , .A1( us01_n742 ) , .A2( us01_n813 ) );
  AOI21_X1 us01_U292 (.ZN( us01_n591 ) , .B1( us01_n748 ) , .A( us01_n790 ) , .B2( us01_n811 ) );
  NOR2_X1 us01_U293 (.ZN( us01_n564 ) , .A2( us01_n695 ) , .A1( us01_n761 ) );
  AOI21_X1 us01_U294 (.ZN( us01_n512 ) , .A( us01_n777 ) , .B2( us01_n790 ) , .B1( us01_n810 ) );
  NAND2_X2 us01_U295 (.A2( us01_n462 ) , .A1( us01_n463 ) , .ZN( us01_n810 ) );
  AOI21_X1 us01_U296 (.ZN( us01_n637 ) , .B2( us01_n747 ) , .A( us01_n786 ) , .B1( us01_n810 ) );
  NOR2_X1 us01_U297 (.ZN( us01_n557 ) , .A2( us01_n789 ) , .A1( us01_n801 ) );
  NOR2_X1 us01_U298 (.A2( us01_n811 ) , .A1( us01_n813 ) , .ZN( us01_n819 ) );
  NOR2_X1 us01_U299 (.ZN( us01_n527 ) , .A1( us01_n706 ) , .A2( us01_n777 ) );
  NAND2_X2 us01_U3 (.A1( us01_n447 ) , .A2( us01_n462 ) , .ZN( us01_n722 ) );
  NOR4_X1 us01_U30 (.A4( us01_n512 ) , .A3( us01_n513 ) , .A2( us01_n514 ) , .A1( us01_n515 ) , .ZN( us01_n522 ) );
  NOR2_X1 us01_U300 (.ZN( us01_n517 ) , .A2( us01_n697 ) , .A1( us01_n814 ) );
  NOR2_X1 us01_U301 (.ZN( us01_n681 ) , .A2( us01_n697 ) , .A1( us01_n801 ) );
  NOR2_X1 us01_U302 (.ZN( us01_n576 ) , .A1( us01_n706 ) , .A2( us01_n811 ) );
  INV_X1 us01_U303 (.A( us01_n813 ) , .ZN( us01_n853 ) );
  INV_X1 us01_U304 (.A( us01_n811 ) , .ZN( us01_n834 ) );
  AOI21_X1 us01_U305 (.ZN( us01_n448 ) , .B2( us01_n790 ) , .A( us01_n801 ) , .B1( us01_n813 ) );
  AOI21_X1 us01_U306 (.ZN( us01_n538 ) , .A( us01_n761 ) , .B2( us01_n777 ) , .B1( us01_n815 ) );
  AOI21_X1 us01_U307 (.ZN( us01_n496 ) , .A( us01_n722 ) , .B2( us01_n760 ) , .B1( us01_n812 ) );
  AOI21_X1 us01_U308 (.ZN( us01_n687 ) , .B2( us01_n747 ) , .B1( us01_n761 ) , .A( us01_n804 ) );
  AOI21_X1 us01_U309 (.B1( us01_n684 ) , .ZN( us01_n685 ) , .A( us01_n726 ) , .B2( us01_n759 ) );
  AOI222_X1 us01_U31 (.ZN( us01_n523 ) , .A1( us01_n832 ) , .B2( us01_n835 ) , .C1( us01_n842 ) , .C2( us01_n848 ) , .A2( us01_n850 ) , .B1( us01_n864 ) );
  NOR2_X1 us01_U310 (.ZN( us01_n581 ) , .A1( us01_n790 ) , .A2( us01_n815 ) );
  NOR2_X1 us01_U311 (.ZN( us01_n532 ) , .A1( us01_n722 ) , .A2( us01_n786 ) );
  NOR2_X1 us01_U312 (.ZN( us01_n630 ) , .A2( us01_n695 ) , .A1( us01_n722 ) );
  AOI21_X1 us01_U313 (.A( us01_n788 ) , .B2( us01_n789 ) , .B1( us01_n790 ) , .ZN( us01_n791 ) );
  AOI21_X1 us01_U314 (.A( us01_n731 ) , .ZN( us01_n732 ) , .B2( us01_n778 ) , .B1( us01_n790 ) );
  NOR2_X1 us01_U315 (.ZN( us01_n565 ) , .A1( us01_n745 ) , .A2( us01_n803 ) );
  AOI21_X1 us01_U316 (.ZN( us01_n567 ) , .B1( us01_n748 ) , .B2( us01_n760 ) , .A( us01_n778 ) );
  AOI21_X1 us01_U317 (.ZN( us01_n638 ) , .B2( us01_n745 ) , .A( us01_n790 ) , .B1( us01_n801 ) );
  AOI21_X1 us01_U318 (.ZN( us01_n562 ) , .B1( us01_n722 ) , .A( us01_n777 ) , .B2( us01_n789 ) );
  AOI21_X1 us01_U319 (.ZN( us01_n569 ) , .B2( us01_n695 ) , .B1( us01_n804 ) , .A( us01_n810 ) );
  NOR4_X1 us01_U32 (.A3( us01_n519 ) , .A1( us01_n520 ) , .ZN( us01_n521 ) , .A2( us01_n671 ) , .A4( us01_n767 ) );
  NOR2_X1 us01_U320 (.ZN( us01_n663 ) , .A1( us01_n778 ) , .A2( us01_n811 ) );
  NOR2_X1 us01_U321 (.ZN( us01_n578 ) , .A2( us01_n695 ) , .A1( us01_n789 ) );
  NOR2_X1 us01_U322 (.ZN( us01_n682 ) , .A1( us01_n789 ) , .A2( us01_n811 ) );
  NAND2_X2 us01_U323 (.A1( us01_n450 ) , .A2( us01_n463 ) , .ZN( us01_n667 ) );
  NAND2_X1 us01_U324 (.ZN( us01_n751 ) , .A1( us01_n761 ) , .A2( us01_n803 ) );
  NOR2_X1 us01_U325 (.ZN( us01_n709 ) , .A1( us01_n760 ) , .A2( us01_n761 ) );
  AOI21_X1 us01_U326 (.ZN( us01_n476 ) , .B2( us01_n695 ) , .A( us01_n747 ) , .B1( us01_n777 ) );
  NOR2_X1 us01_U327 (.ZN( us01_n680 ) , .A2( us01_n706 ) , .A1( us01_n815 ) );
  INV_X1 us01_U328 (.A( us01_n778 ) , .ZN( us01_n848 ) );
  OAI21_X1 us01_U329 (.A( us01_n729 ) , .B1( us01_n730 ) , .ZN( us01_n734 ) , .B2( us01_n803 ) );
  AOI221_X1 us01_U33 (.A( us01_n779 ) , .ZN( us01_n796 ) , .C2( us01_n835 ) , .B2( us01_n836 ) , .B1( us01_n863 ) , .C1( us01_n864 ) );
  OAI21_X1 us01_U330 (.ZN( us01_n729 ) , .A( us01_n831 ) , .B2( us01_n850 ) , .B1( us01_n871 ) );
  AOI21_X1 us01_U331 (.ZN( us01_n639 ) , .B1( us01_n678 ) , .A( us01_n789 ) , .B2( us01_n815 ) );
  AOI21_X1 us01_U332 (.ZN( us01_n440 ) , .A( us01_n697 ) , .B1( us01_n731 ) , .B2( us01_n748 ) );
  NAND2_X1 us01_U333 (.A1( us01_n697 ) , .A2( us01_n727 ) , .ZN( us01_n780 ) );
  NOR2_X1 us01_U334 (.ZN( us01_n468 ) , .A2( us01_n777 ) , .A1( us01_n813 ) );
  NOR2_X1 us01_U335 (.ZN( us01_n516 ) , .A1( us01_n706 ) , .A2( us01_n786 ) );
  NAND2_X2 us01_U336 (.A2( us01_n447 ) , .A1( us01_n450 ) , .ZN( us01_n761 ) );
  OAI21_X1 us01_U337 (.A( us01_n696 ) , .ZN( us01_n700 ) , .B2( us01_n748 ) , .B1( us01_n802 ) );
  OAI21_X1 us01_U338 (.ZN( us01_n696 ) , .B2( us01_n831 ) , .B1( us01_n836 ) , .A( us01_n858 ) );
  NOR2_X1 us01_U339 (.ZN( us01_n524 ) , .A1( us01_n722 ) , .A2( us01_n748 ) );
  NOR4_X1 us01_U34 (.A4( us01_n791 ) , .A3( us01_n792 ) , .A2( us01_n793 ) , .A1( us01_n794 ) , .ZN( us01_n795 ) );
  AOI21_X1 us01_U340 (.ZN( us01_n441 ) , .B1( us01_n787 ) , .B2( us01_n789 ) , .A( us01_n812 ) );
  AOI21_X1 us01_U341 (.ZN( us01_n495 ) , .A( us01_n777 ) , .B2( us01_n789 ) , .B1( us01_n802 ) );
  NAND2_X1 us01_U342 (.ZN( us01_n712 ) , .A1( us01_n726 ) , .A2( us01_n778 ) );
  NOR2_X1 us01_U343 (.ZN( us01_n482 ) , .A1( us01_n786 ) , .A2( us01_n803 ) );
  NAND2_X1 us01_U344 (.A2( us01_n760 ) , .A1( us01_n804 ) , .ZN( us01_n808 ) );
  OAI21_X1 us01_U345 (.A( us01_n785 ) , .B2( us01_n786 ) , .B1( us01_n787 ) , .ZN( us01_n793 ) );
  OAI21_X1 us01_U346 (.ZN( us01_n785 ) , .A( us01_n837 ) , .B1( us01_n861 ) , .B2( us01_n871 ) );
  INV_X1 us01_U347 (.A( us01_n783 ) , .ZN( us01_n844 ) );
  NOR2_X1 us01_U348 (.ZN( us01_n710 ) , .A2( us01_n722 ) , .A1( us01_n788 ) );
  NAND2_X1 us01_U349 (.ZN( us01_n669 ) , .A1( us01_n804 ) , .A2( us01_n814 ) );
  NOR4_X1 us01_U35 (.A4( us01_n774 ) , .A3( us01_n775 ) , .A1( us01_n776 ) , .ZN( us01_n797 ) , .A2( us01_n799 ) );
  NAND2_X2 us01_U350 (.A2( us01_n446 ) , .A1( us01_n450 ) , .ZN( us01_n727 ) );
  INV_X1 us01_U351 (.A( us01_n722 ) , .ZN( us01_n854 ) );
  NAND2_X2 us01_U352 (.A1( us01_n445 ) , .A2( us01_n463 ) , .ZN( us01_n747 ) );
  INV_X1 us01_U353 (.A( us01_n815 ) , .ZN( us01_n842 ) );
  AND2_X1 us01_U354 (.ZN( us01_n730 ) , .A1( us01_n777 ) , .A2( us01_n783 ) );
  NAND2_X1 us01_U355 (.A1( us01_n445 ) , .A2( us01_n447 ) , .ZN( us01_n803 ) );
  NAND2_X1 us01_U356 (.A1( us01_n449 ) , .A2( us01_n452 ) , .ZN( us01_n812 ) );
  NAND2_X1 us01_U357 (.A1( us01_n453 ) , .A2( us01_n469 ) , .ZN( us01_n801 ) );
  NAND2_X1 us01_U358 (.A1( us01_n453 ) , .A2( us01_n460 ) , .ZN( us01_n748 ) );
  NAND2_X2 us01_U359 (.A2( us01_n446 ) , .A1( us01_n458 ) , .ZN( us01_n726 ) );
  NOR2_X1 us01_U36 (.ZN( us01_n802 ) , .A1( us01_n852 ) , .A2( us01_n859 ) );
  NAND2_X1 us01_U360 (.A2( us01_n451 ) , .A1( us01_n453 ) , .ZN( us01_n804 ) );
  NAND2_X1 us01_U361 (.A1( us01_n449 ) , .A2( us01_n469 ) , .ZN( us01_n814 ) );
  NAND2_X1 us01_U362 (.A1( us01_n452 ) , .A2( us01_n459 ) , .ZN( us01_n811 ) );
  NAND2_X1 us01_U363 (.A1( us01_n451 ) , .A2( us01_n459 ) , .ZN( us01_n742 ) );
  NAND2_X1 us01_U364 (.A1( us01_n451 ) , .A2( us01_n470 ) , .ZN( us01_n783 ) );
  NAND2_X1 us01_U365 (.A2( us01_n452 ) , .A1( us01_n470 ) , .ZN( us01_n777 ) );
  NAND2_X1 us01_U366 (.A2( us01_n459 ) , .A1( us01_n460 ) , .ZN( us01_n745 ) );
  NAND2_X2 us01_U367 (.A2( us01_n446 ) , .A1( us01_n462 ) , .ZN( us01_n813 ) );
  NAND2_X1 us01_U368 (.A1( us01_n460 ) , .A2( us01_n470 ) , .ZN( us01_n786 ) );
  NOR2_X1 us01_U369 (.ZN( us01_n451 ) , .A1( us01_n824 ) , .A2( us01_n825 ) );
  NAND4_X1 us01_U37 (.ZN( sa01_sr_2 ) , .A4( us01_n641 ) , .A3( us01_n642 ) , .A2( us01_n643 ) , .A1( us01_n644 ) );
  NOR2_X1 us01_U370 (.ZN( us01_n449 ) , .A1( us01_n826 ) , .A2( us01_n827 ) );
  NAND2_X1 us01_U371 (.A1( us01_n449 ) , .A2( us01_n460 ) , .ZN( us01_n788 ) );
  NAND2_X2 us01_U372 (.A1( us01_n447 ) , .A2( us01_n458 ) , .ZN( us01_n790 ) );
  NAND2_X2 us01_U373 (.A2( us01_n439 ) , .A1( us01_n450 ) , .ZN( us01_n789 ) );
  NAND2_X1 us01_U374 (.A2( us01_n452 ) , .A1( us01_n453 ) , .ZN( us01_n728 ) );
  NAND2_X2 us01_U375 (.A2( us01_n469 ) , .A1( us01_n470 ) , .ZN( us01_n815 ) );
  NAND2_X1 us01_U376 (.A1( us01_n445 ) , .A2( us01_n446 ) , .ZN( us01_n784 ) );
  NAND2_X2 us01_U377 (.A2( us01_n439 ) , .A1( us01_n445 ) , .ZN( us01_n782 ) );
  NOR2_X1 us01_U378 (.A2( sa01_7 ) , .ZN( us01_n458 ) , .A1( us01_n847 ) );
  NOR2_X1 us01_U379 (.A2( sa01_2 ) , .A1( sa01_3 ) , .ZN( us01_n470 ) );
  AOI222_X1 us01_U38 (.B2( us01_n636 ) , .ZN( us01_n642 ) , .B1( us01_n839 ) , .A1( us01_n840 ) , .C2( us01_n844 ) , .C1( us01_n861 ) , .A2( us01_n863 ) );
  NOR2_X1 us01_U380 (.A2( sa01_1 ) , .ZN( us01_n469 ) , .A1( us01_n824 ) );
  NOR2_X1 us01_U381 (.A2( sa01_0 ) , .ZN( us01_n452 ) , .A1( us01_n825 ) );
  NOR2_X1 us01_U382 (.A2( sa01_0 ) , .A1( sa01_1 ) , .ZN( us01_n460 ) );
  NAND2_X2 us01_U383 (.A1( us01_n439 ) , .A2( us01_n458 ) , .ZN( us01_n697 ) );
  NOR2_X1 us01_U384 (.A2( sa01_3 ) , .ZN( us01_n453 ) , .A1( us01_n826 ) );
  NOR2_X1 us01_U385 (.A2( sa01_2 ) , .ZN( us01_n459 ) , .A1( us01_n827 ) );
  INV_X1 us01_U386 (.A( sa01_3 ) , .ZN( us01_n827 ) );
  INV_X1 us01_U387 (.A( sa01_1 ) , .ZN( us01_n825 ) );
  INV_X1 us01_U388 (.A( sa01_0 ) , .ZN( us01_n824 ) );
  INV_X1 us01_U389 (.A( sa01_2 ) , .ZN( us01_n826 ) );
  NOR4_X1 us01_U39 (.A4( us01_n637 ) , .A3( us01_n638 ) , .A2( us01_n639 ) , .A1( us01_n640 ) , .ZN( us01_n641 ) );
  INV_X1 us01_U390 (.A( sa01_5 ) , .ZN( us01_n846 ) );
  NAND2_X1 us01_U391 (.A1( us01_n727 ) , .A2( us01_n782 ) , .ZN( us01_n809 ) );
  OAI22_X1 us01_U392 (.ZN( us01_n586 ) , .A2( us01_n745 ) , .B2( us01_n760 ) , .A1( us01_n761 ) , .B1( us01_n782 ) );
  AOI21_X1 us01_U393 (.ZN( us01_n590 ) , .B1( us01_n726 ) , .B2( us01_n782 ) , .A( us01_n788 ) );
  AOI21_X1 us01_U394 (.ZN( us01_n646 ) , .A( us01_n760 ) , .B2( us01_n782 ) , .B1( us01_n790 ) );
  AOI21_X1 us01_U395 (.ZN( us01_n621 ) , .B1( us01_n697 ) , .A( us01_n777 ) , .B2( us01_n782 ) );
  OAI22_X1 us01_U396 (.ZN( us01_n679 ) , .A1( us01_n697 ) , .A2( us01_n728 ) , .B2( us01_n782 ) , .B1( us01_n815 ) );
  OAI21_X1 us01_U397 (.A( us01_n611 ) , .ZN( us01_n614 ) , .B1( us01_n623 ) , .B2( us01_n782 ) );
  NOR2_X1 us01_U398 (.ZN( us01_n608 ) , .A1( us01_n782 ) , .A2( us01_n814 ) );
  INV_X2 us01_U399 (.A( us01_n747 ) , .ZN( us01_n861 ) );
  NAND2_X2 us01_U4 (.A1( us01_n439 ) , .A2( us01_n462 ) , .ZN( us01_n706 ) );
  NOR3_X1 us01_U40 (.A2( us01_n605 ) , .A1( us01_n606 ) , .ZN( us01_n644 ) , .A3( us01_n720 ) );
  OAI222_X1 us01_U400 (.A2( us01_n667 ) , .ZN( us01_n672 ) , .B1( us01_n745 ) , .B2( us01_n782 ) , .C2( us01_n786 ) , .C1( us01_n813 ) , .A1( us01_n815 ) );
  NOR2_X1 us01_U401 (.ZN( us01_n649 ) , .A1( us01_n782 ) , .A2( us01_n786 ) );
  NOR2_X1 us01_U402 (.ZN( us01_n598 ) , .A2( us01_n695 ) , .A1( us01_n782 ) );
  NOR2_X1 us01_U403 (.ZN( us01_n551 ) , .A2( us01_n742 ) , .A1( us01_n782 ) );
  INV_X1 us01_U404 (.A( us01_n782 ) , .ZN( us01_n859 ) );
  NAND2_X1 us01_U405 (.A2( us01_n459 ) , .A1( us01_n469 ) , .ZN( us01_n695 ) );
  INV_X1 us01_U406 (.A( sa01_7 ) , .ZN( us01_n856 ) );
  OAI221_X1 us01_U407 (.A( us01_n781 ) , .C2( us01_n782 ) , .B2( us01_n783 ) , .B1( us01_n784 ) , .ZN( us01_n794 ) , .C1( us01_n811 ) );
  AOI21_X1 us01_U408 (.ZN( us01_n498 ) , .A( us01_n695 ) , .B1( us01_n706 ) , .B2( us01_n784 ) );
  OAI221_X1 us01_U409 (.A( us01_n694 ) , .ZN( us01_n701 ) , .C2( us01_n782 ) , .C1( us01_n783 ) , .B1( us01_n784 ) , .B2( us01_n804 ) );
  NAND4_X1 us01_U41 (.ZN( sa01_sr_7 ) , .A4( us01_n820 ) , .A3( us01_n821 ) , .A2( us01_n822 ) , .A1( us01_n823 ) );
  OAI22_X1 us01_U410 (.ZN( us01_n588 ) , .B1( us01_n728 ) , .B2( us01_n747 ) , .A2( us01_n784 ) , .A1( us01_n801 ) );
  AOI222_X1 us01_U411 (.ZN( us01_n511 ) , .C1( us01_n830 ) , .B2( us01_n835 ) , .A2( us01_n841 ) , .C2( us01_n860 ) , .B1( us01_n861 ) , .A1( us01_n864 ) );
  AOI222_X1 us01_U412 (.ZN( us01_n603 ) , .B2( us01_n669 ) , .B1( us01_n751 ) , .C2( us01_n829 ) , .A1( us01_n831 ) , .A2( us01_n860 ) , .C1( us01_n861 ) );
  AOI221_X1 us01_U413 (.A( us01_n481 ) , .ZN( us01_n486 ) , .B1( us01_n829 ) , .C2( us01_n842 ) , .C1( us01_n850 ) , .B2( us01_n860 ) );
  NAND2_X1 us01_U414 (.A2( us01_n747 ) , .A1( us01_n784 ) , .ZN( us01_n807 ) );
  NOR2_X1 us01_U415 (.ZN( us01_n610 ) , .A1( us01_n777 ) , .A2( us01_n784 ) );
  NOR2_X1 us01_U416 (.ZN( us01_n715 ) , .A2( us01_n742 ) , .A1( us01_n784 ) );
  OAI222_X1 us01_U417 (.ZN( us01_n615 ) , .B1( us01_n695 ) , .C1( us01_n722 ) , .C2( us01_n745 ) , .B2( us01_n784 ) , .A2( us01_n790 ) , .A1( us01_n814 ) );
  NOR2_X1 us01_U418 (.ZN( us01_n651 ) , .A1( us01_n760 ) , .A2( us01_n784 ) );
  NOR2_X1 us01_U419 (.ZN( us01_n552 ) , .A1( us01_n784 ) , .A2( us01_n811 ) );
  AOI222_X1 us01_U42 (.C2( us01_n807 ) , .B2( us01_n808 ) , .A2( us01_n809 ) , .ZN( us01_n821 ) , .C1( us01_n830 ) , .A1( us01_n837 ) , .B1( us01_n851 ) );
  NOR2_X1 us01_U420 (.ZN( us01_n787 ) , .A2( us01_n860 ) , .A1( us01_n866 ) );
  NOR2_X1 us01_U421 (.ZN( us01_n699 ) , .A2( us01_n784 ) , .A1( us01_n815 ) );
  NOR2_X1 us01_U422 (.A1( us01_n728 ) , .ZN( us01_n763 ) , .A2( us01_n784 ) );
  INV_X1 us01_U423 (.A( us01_n784 ) , .ZN( us01_n860 ) );
  NOR2_X1 us01_U424 (.A2( sa01_4 ) , .ZN( us01_n447 ) , .A1( us01_n846 ) );
  NOR2_X1 us01_U425 (.ZN( us01_n463 ) , .A2( us01_n845 ) , .A1( us01_n846 ) );
  NOR2_X1 us01_U426 (.A2( sa01_5 ) , .ZN( us01_n446 ) , .A1( us01_n845 ) );
  NOR2_X1 us01_U427 (.A2( sa01_4 ) , .A1( sa01_5 ) , .ZN( us01_n439 ) );
  INV_X1 us01_U428 (.A( sa01_6 ) , .ZN( us01_n847 ) );
  NOR2_X1 us01_U429 (.ZN( us01_n445 ) , .A2( us01_n847 ) , .A1( us01_n856 ) );
  NOR4_X1 us01_U43 (.A4( us01_n816 ) , .A3( us01_n817 ) , .A2( us01_n818 ) , .A1( us01_n819 ) , .ZN( us01_n820 ) );
  NOR2_X1 us01_U430 (.A2( sa01_6 ) , .ZN( us01_n450 ) , .A1( us01_n856 ) );
  NOR2_X1 us01_U431 (.A2( sa01_6 ) , .A1( sa01_7 ) , .ZN( us01_n462 ) );
  AOI221_X1 us01_U432 (.A( us01_n574 ) , .ZN( us01_n585 ) , .B2( us01_n829 ) , .C2( us01_n841 ) , .B1( us01_n852 ) , .C1( us01_n859 ) );
  AOI21_X1 us01_U433 (.ZN( us01_n574 ) , .B2( us01_n722 ) , .B1( us01_n746 ) , .A( us01_n783 ) );
  INV_X1 us01_U434 (.A( sa01_4 ) , .ZN( us01_n845 ) );
  AOI211_X1 us01_U435 (.A( us01_n635 ) , .ZN( us01_n643 ) , .B( us01_n741 ) , .C2( us01_n837 ) , .C1( us01_n852 ) );
  NAND4_X1 us01_U436 (.A4( us01_n631 ) , .A3( us01_n632 ) , .A2( us01_n633 ) , .A1( us01_n634 ) , .ZN( us01_n741 ) );
  NAND3_X1 us01_U437 (.ZN( sa01_sr_6 ) , .A3( us01_n795 ) , .A2( us01_n796 ) , .A1( us01_n797 ) );
  NAND3_X1 us01_U438 (.ZN( sa01_sr_5 ) , .A3( us01_n756 ) , .A2( us01_n757 ) , .A1( us01_n758 ) );
  NAND3_X1 us01_U439 (.ZN( sa01_sr_4 ) , .A3( us01_n736 ) , .A2( us01_n737 ) , .A1( us01_n738 ) );
  AOI211_X1 us01_U44 (.B( us01_n805 ) , .A( us01_n806 ) , .ZN( us01_n822 ) , .C1( us01_n840 ) , .C2( us01_n848 ) );
  NAND3_X1 us01_U440 (.A3( us01_n673 ) , .A2( us01_n674 ) , .A1( us01_n675 ) , .ZN( us01_n805 ) );
  NAND3_X1 us01_U441 (.ZN( us01_n636 ) , .A3( us01_n706 ) , .A2( us01_n722 ) , .A1( us01_n790 ) );
  NAND3_X1 us01_U442 (.A3( us01_n616 ) , .A2( us01_n617 ) , .A1( us01_n618 ) , .ZN( us01_n723 ) );
  NAND3_X1 us01_U443 (.A3( us01_n583 ) , .A2( us01_n584 ) , .A1( us01_n585 ) , .ZN( us01_n619 ) );
  NAND3_X1 us01_U444 (.ZN( us01_n563 ) , .A3( us01_n678 ) , .A2( us01_n748 ) , .A1( us01_n783 ) );
  NAND3_X1 us01_U445 (.A3( us01_n521 ) , .A2( us01_n522 ) , .A1( us01_n523 ) , .ZN( us01_n740 ) );
  NAND3_X1 us01_U446 (.A3( us01_n510 ) , .A1( us01_n511 ) , .ZN( us01_n606 ) , .A2( us01_n869 ) );
  NAND3_X1 us01_U447 (.A3( us01_n465 ) , .A2( us01_n466 ) , .A1( us01_n467 ) , .ZN( us01_n775 ) );
  NAND4_X1 us01_U45 (.ZN( sa01_sr_0 ) , .A4( us01_n499 ) , .A3( us01_n500 ) , .A2( us01_n501 ) , .A1( us01_n502 ) );
  NOR4_X1 us01_U46 (.A4( us01_n496 ) , .A3( us01_n497 ) , .A2( us01_n498 ) , .ZN( us01_n499 ) , .A1( us01_n525 ) );
  AOI221_X1 us01_U47 (.A( us01_n495 ) , .ZN( us01_n500 ) , .B2( us01_n841 ) , .C1( us01_n844 ) , .C2( us01_n858 ) , .B1( us01_n860 ) );
  AOI211_X1 us01_U48 (.A( us01_n494 ) , .ZN( us01_n501 ) , .B( us01_n800 ) , .C2( us01_n837 ) , .C1( us01_n849 ) );
  NOR2_X1 us01_U49 (.ZN( us01_n746 ) , .A1( us01_n859 ) , .A2( us01_n860 ) );
  NAND2_X2 us01_U5 (.A2( us01_n458 ) , .A1( us01_n463 ) , .ZN( us01_n778 ) );
  NAND4_X1 us01_U50 (.ZN( sa01_sr_1 ) , .A4( us01_n593 ) , .A3( us01_n594 ) , .A2( us01_n595 ) , .A1( us01_n596 ) );
  AOI211_X1 us01_U51 (.B( us01_n587 ) , .A( us01_n588 ) , .ZN( us01_n594 ) , .C2( us01_n809 ) , .C1( us01_n831 ) );
  NOR4_X1 us01_U52 (.A4( us01_n589 ) , .A3( us01_n590 ) , .A2( us01_n591 ) , .A1( us01_n592 ) , .ZN( us01_n593 ) );
  AOI211_X1 us01_U53 (.A( us01_n586 ) , .ZN( us01_n595 ) , .B( us01_n619 ) , .C1( us01_n843 ) , .C2( us01_n853 ) );
  NOR2_X1 us01_U54 (.ZN( us01_n623 ) , .A2( us01_n834 ) , .A1( us01_n837 ) );
  NAND4_X1 us01_U55 (.A4( us01_n601 ) , .A3( us01_n602 ) , .A2( us01_n603 ) , .A1( us01_n604 ) , .ZN( us01_n720 ) );
  NOR3_X1 us01_U56 (.A1( us01_n597 ) , .ZN( us01_n602 ) , .A3( us01_n661 ) , .A2( us01_n768 ) );
  NOR4_X1 us01_U57 (.A3( us01_n598 ) , .A2( us01_n599 ) , .A1( us01_n600 ) , .ZN( us01_n601 ) , .A4( us01_n653 ) );
  AOI222_X1 us01_U58 (.ZN( us01_n604 ) , .A1( us01_n828 ) , .C2( us01_n835 ) , .B1( us01_n840 ) , .A2( us01_n854 ) , .B2( us01_n859 ) , .C1( us01_n866 ) );
  NOR4_X1 us01_U59 (.A4( us01_n575 ) , .A3( us01_n576 ) , .A2( us01_n577 ) , .ZN( us01_n584 ) , .A1( us01_n681 ) );
  INV_X1 us01_U6 (.A( us01_n667 ) , .ZN( us01_n863 ) );
  NOR4_X1 us01_U60 (.A1( us01_n582 ) , .ZN( us01_n583 ) , .A3( us01_n650 ) , .A2( us01_n660 ) , .A4( us01_n765 ) );
  NAND4_X1 us01_U61 (.A4( us01_n483 ) , .A3( us01_n484 ) , .A2( us01_n485 ) , .A1( us01_n486 ) , .ZN( us01_n776 ) );
  NOR4_X1 us01_U62 (.A4( us01_n482 ) , .ZN( us01_n485 ) , .A1( us01_n564 ) , .A2( us01_n579 ) , .A3( us01_n600 ) );
  NOR4_X1 us01_U63 (.ZN( us01_n483 ) , .A2( us01_n531 ) , .A1( us01_n556 ) , .A3( us01_n629 ) , .A4( us01_n716 ) );
  NOR4_X1 us01_U64 (.ZN( us01_n484 ) , .A1( us01_n505 ) , .A2( us01_n517 ) , .A4( us01_n544 ) , .A3( us01_n609 ) );
  NOR4_X1 us01_U65 (.A4( us01_n627 ) , .A3( us01_n628 ) , .A2( us01_n629 ) , .A1( us01_n630 ) , .ZN( us01_n631 ) );
  AOI211_X1 us01_U66 (.B( us01_n621 ) , .A( us01_n622 ) , .ZN( us01_n633 ) , .C2( us01_n834 ) , .C1( us01_n861 ) );
  NOR4_X1 us01_U67 (.A4( us01_n624 ) , .A3( us01_n625 ) , .A2( us01_n626 ) , .ZN( us01_n632 ) , .A1( us01_n662 ) );
  NAND4_X1 us01_U68 (.A4( us01_n655 ) , .A3( us01_n656 ) , .A2( us01_n657 ) , .A1( us01_n658 ) , .ZN( us01_n798 ) );
  NOR3_X1 us01_U69 (.A3( us01_n649 ) , .A2( us01_n650 ) , .A1( us01_n651 ) , .ZN( us01_n656 ) );
  NOR3_X1 us01_U7 (.ZN( us01_n596 ) , .A1( us01_n606 ) , .A3( us01_n721 ) , .A2( us01_n740 ) );
  NOR3_X1 us01_U70 (.A3( us01_n652 ) , .A2( us01_n653 ) , .A1( us01_n654 ) , .ZN( us01_n655 ) );
  NOR3_X1 us01_U71 (.A3( us01_n646 ) , .A2( us01_n647 ) , .A1( us01_n648 ) , .ZN( us01_n657 ) );
  NAND4_X1 us01_U72 (.A4( us01_n558 ) , .A3( us01_n559 ) , .A2( us01_n560 ) , .A1( us01_n561 ) , .ZN( us01_n605 ) );
  NOR4_X1 us01_U73 (.ZN( us01_n559 ) , .A1( us01_n651 ) , .A3( us01_n659 ) , .A4( us01_n683 ) , .A2( us01_n766 ) );
  NOR4_X1 us01_U74 (.A4( us01_n550 ) , .A3( us01_n551 ) , .A2( us01_n552 ) , .A1( us01_n553 ) , .ZN( us01_n560 ) );
  NOR4_X1 us01_U75 (.A4( us01_n554 ) , .A3( us01_n555 ) , .A2( us01_n556 ) , .A1( us01_n557 ) , .ZN( us01_n558 ) );
  NAND4_X1 us01_U76 (.A4( us01_n770 ) , .A3( us01_n771 ) , .A2( us01_n772 ) , .A1( us01_n773 ) , .ZN( us01_n799 ) );
  NOR3_X1 us01_U77 (.A3( us01_n763 ) , .A2( us01_n764 ) , .A1( us01_n765 ) , .ZN( us01_n771 ) );
  NOR4_X1 us01_U78 (.A4( us01_n766 ) , .A3( us01_n767 ) , .A2( us01_n768 ) , .A1( us01_n769 ) , .ZN( us01_n770 ) );
  AOI222_X1 us01_U79 (.ZN( us01_n773 ) , .A1( us01_n828 ) , .C1( us01_n832 ) , .B2( us01_n839 ) , .A2( us01_n848 ) , .B1( us01_n859 ) , .C2( us01_n871 ) );
  NOR3_X1 us01_U8 (.A3( us01_n798 ) , .A2( us01_n799 ) , .A1( us01_n800 ) , .ZN( us01_n823 ) );
  NOR4_X1 us01_U80 (.A4( us01_n507 ) , .A2( us01_n508 ) , .A1( us01_n509 ) , .ZN( us01_n510 ) , .A3( us01_n668 ) );
  INV_X1 us01_U81 (.A( us01_n503 ) , .ZN( us01_n869 ) );
  NOR4_X1 us01_U82 (.A4( us01_n663 ) , .A3( us01_n664 ) , .A2( us01_n665 ) , .A1( us01_n666 ) , .ZN( us01_n674 ) );
  NOR4_X1 us01_U83 (.A4( us01_n659 ) , .A3( us01_n660 ) , .A2( us01_n661 ) , .A1( us01_n662 ) , .ZN( us01_n675 ) );
  NOR4_X1 us01_U84 (.A3( us01_n671 ) , .A1( us01_n672 ) , .ZN( us01_n673 ) , .A4( us01_n713 ) , .A2( us01_n857 ) );
  NOR2_X1 us01_U85 (.ZN( us01_n759 ) , .A1( us01_n831 ) , .A2( us01_n832 ) );
  NAND4_X1 us01_U86 (.A4( us01_n454 ) , .A3( us01_n455 ) , .A2( us01_n456 ) , .A1( us01_n457 ) , .ZN( us01_n677 ) );
  NOR3_X1 us01_U87 (.ZN( us01_n455 ) , .A3( us01_n528 ) , .A1( us01_n553 ) , .A2( us01_n568 ) );
  AOI221_X1 us01_U88 (.A( us01_n448 ) , .ZN( us01_n457 ) , .C2( us01_n751 ) , .B1( us01_n830 ) , .C1( us01_n840 ) , .B2( us01_n859 ) );
  NOR4_X1 us01_U89 (.ZN( us01_n456 ) , .A2( us01_n507 ) , .A1( us01_n597 ) , .A4( us01_n626 ) , .A3( us01_n709 ) );
  NOR3_X1 us01_U9 (.A3( us01_n619 ) , .A2( us01_n620 ) , .ZN( us01_n634 ) , .A1( us01_n723 ) );
  NAND4_X1 us01_U90 (.A4( us01_n533 ) , .A3( us01_n534 ) , .A2( us01_n535 ) , .A1( us01_n536 ) , .ZN( us01_n620 ) );
  NOR4_X1 us01_U91 (.A4( us01_n524 ) , .A2( us01_n525 ) , .A1( us01_n526 ) , .ZN( us01_n536 ) , .A3( us01_n699 ) );
  NOR4_X1 us01_U92 (.A1( us01_n529 ) , .ZN( us01_n534 ) , .A2( us01_n652 ) , .A4( us01_n666 ) , .A3( us01_n763 ) );
  NOR4_X1 us01_U93 (.A4( us01_n527 ) , .A3( us01_n528 ) , .ZN( us01_n535 ) , .A2( us01_n682 ) , .A1( us01_n792 ) );
  NAND4_X1 us01_U94 (.A4( us01_n477 ) , .A3( us01_n478 ) , .A2( us01_n479 ) , .A1( us01_n480 ) , .ZN( us01_n692 ) );
  NOR3_X1 us01_U95 (.ZN( us01_n478 ) , .A2( us01_n506 ) , .A3( us01_n599 ) , .A1( us01_n608 ) );
  AOI211_X1 us01_U96 (.B( us01_n475 ) , .A( us01_n476 ) , .ZN( us01_n480 ) , .C2( us01_n831 ) , .C1( us01_n859 ) );
  NOR4_X1 us01_U97 (.ZN( us01_n479 ) , .A3( us01_n530 ) , .A4( us01_n543 ) , .A2( us01_n565 ) , .A1( us01_n715 ) );
  NAND4_X1 us01_U98 (.A4( us01_n546 ) , .A3( us01_n547 ) , .A2( us01_n548 ) , .A1( us01_n549 ) , .ZN( us01_n743 ) );
  NOR3_X1 us01_U99 (.ZN( us01_n547 ) , .A2( us01_n649 ) , .A1( us01_n665 ) , .A3( us01_n769 ) );
endmodule

