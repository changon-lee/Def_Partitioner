module aes_aes_die_15 ( u0_n242, u0_n244, u0_n262, u0_rcon_26, u0_rcon_27, u0_rcon_29, u0_rcon_30, u0_rcon_31, w0_26, 
       w0_27, w0_29, w0_30, w0_31, w3_16, w3_17, w3_18, w3_19, w3_20, 
       w3_21, w3_22, w3_23, w3_26, u0_n1, u0_n11, u0_n164, u0_n172, u0_n3, u0_n5, u0_n80, u0_n82, u0_n9, 
        u0_subword_24, u0_subword_25, u0_subword_28 );
  input u0_n242, u0_n244, u0_n262, u0_rcon_26, u0_rcon_27, u0_rcon_29, u0_rcon_30, u0_rcon_31, w0_26, 
        w0_27, w0_29, w0_30, w0_31, w3_16, w3_17, w3_18, w3_19, w3_20, 
        w3_21, w3_22, w3_23, w3_26;
  output u0_n1, u0_n11, u0_n164, u0_n172, u0_n3, u0_n5, u0_n80, u0_n82, u0_n9, 
        u0_subword_24, u0_subword_25, u0_subword_28;
  wire u0_n226, u0_n228, u0_n230, u0_n234, u0_n236, u0_subword_26, u0_subword_27, u0_subword_29, u0_subword_30, 
       u0_subword_31, u0_u0_n1, u0_u0_n171, u0_u0_n22, u0_u0_n438, u0_u0_n439, u0_u0_n440, u0_u0_n441, u0_u0_n442, 
       u0_u0_n443, u0_u0_n444, u0_u0_n445, u0_u0_n446, u0_u0_n447, u0_u0_n448, u0_u0_n449, u0_u0_n450, u0_u0_n451, 
       u0_u0_n452, u0_u0_n453, u0_u0_n454, u0_u0_n455, u0_u0_n456, u0_u0_n457, u0_u0_n458, u0_u0_n459, u0_u0_n460, 
       u0_u0_n461, u0_u0_n462, u0_u0_n463, u0_u0_n464, u0_u0_n465, u0_u0_n466, u0_u0_n467, u0_u0_n468, u0_u0_n469, 
       u0_u0_n470, u0_u0_n471, u0_u0_n472, u0_u0_n473, u0_u0_n474, u0_u0_n475, u0_u0_n476, u0_u0_n477, u0_u0_n478, 
       u0_u0_n479, u0_u0_n480, u0_u0_n481, u0_u0_n482, u0_u0_n483, u0_u0_n484, u0_u0_n485, u0_u0_n486, u0_u0_n487, 
       u0_u0_n488, u0_u0_n489, u0_u0_n490, u0_u0_n491, u0_u0_n492, u0_u0_n493, u0_u0_n494, u0_u0_n495, u0_u0_n496, 
       u0_u0_n497, u0_u0_n498, u0_u0_n499, u0_u0_n500, u0_u0_n501, u0_u0_n502, u0_u0_n503, u0_u0_n504, u0_u0_n505, 
       u0_u0_n506, u0_u0_n507, u0_u0_n508, u0_u0_n509, u0_u0_n510, u0_u0_n511, u0_u0_n512, u0_u0_n513, u0_u0_n514, 
       u0_u0_n515, u0_u0_n516, u0_u0_n517, u0_u0_n518, u0_u0_n519, u0_u0_n520, u0_u0_n521, u0_u0_n522, u0_u0_n523, 
       u0_u0_n524, u0_u0_n525, u0_u0_n526, u0_u0_n527, u0_u0_n528, u0_u0_n529, u0_u0_n530, u0_u0_n531, u0_u0_n532, 
       u0_u0_n533, u0_u0_n534, u0_u0_n535, u0_u0_n536, u0_u0_n537, u0_u0_n538, u0_u0_n539, u0_u0_n540, u0_u0_n541, 
       u0_u0_n542, u0_u0_n543, u0_u0_n544, u0_u0_n545, u0_u0_n546, u0_u0_n547, u0_u0_n548, u0_u0_n549, u0_u0_n550, 
       u0_u0_n551, u0_u0_n552, u0_u0_n553, u0_u0_n554, u0_u0_n555, u0_u0_n556, u0_u0_n557, u0_u0_n558, u0_u0_n559, 
       u0_u0_n560, u0_u0_n561, u0_u0_n562, u0_u0_n563, u0_u0_n564, u0_u0_n565, u0_u0_n566, u0_u0_n567, u0_u0_n568, 
       u0_u0_n569, u0_u0_n570, u0_u0_n571, u0_u0_n572, u0_u0_n573, u0_u0_n574, u0_u0_n575, u0_u0_n576, u0_u0_n577, 
       u0_u0_n578, u0_u0_n579, u0_u0_n580, u0_u0_n581, u0_u0_n582, u0_u0_n583, u0_u0_n584, u0_u0_n585, u0_u0_n586, 
       u0_u0_n587, u0_u0_n588, u0_u0_n589, u0_u0_n590, u0_u0_n591, u0_u0_n592, u0_u0_n593, u0_u0_n594, u0_u0_n595, 
       u0_u0_n596, u0_u0_n597, u0_u0_n598, u0_u0_n599, u0_u0_n600, u0_u0_n601, u0_u0_n602, u0_u0_n603, u0_u0_n604, 
       u0_u0_n605, u0_u0_n606, u0_u0_n607, u0_u0_n608, u0_u0_n609, u0_u0_n610, u0_u0_n611, u0_u0_n612, u0_u0_n613, 
       u0_u0_n614, u0_u0_n615, u0_u0_n616, u0_u0_n617, u0_u0_n618, u0_u0_n619, u0_u0_n620, u0_u0_n621, u0_u0_n622, 
       u0_u0_n623, u0_u0_n624, u0_u0_n625, u0_u0_n626, u0_u0_n627, u0_u0_n628, u0_u0_n629, u0_u0_n630, u0_u0_n631, 
       u0_u0_n632, u0_u0_n633, u0_u0_n634, u0_u0_n635, u0_u0_n636, u0_u0_n637, u0_u0_n638, u0_u0_n639, u0_u0_n640, 
       u0_u0_n641, u0_u0_n642, u0_u0_n643, u0_u0_n644, u0_u0_n645, u0_u0_n646, u0_u0_n647, u0_u0_n648, u0_u0_n649, 
       u0_u0_n650, u0_u0_n651, u0_u0_n652, u0_u0_n653, u0_u0_n654, u0_u0_n655, u0_u0_n656, u0_u0_n657, u0_u0_n658, 
       u0_u0_n659, u0_u0_n660, u0_u0_n661, u0_u0_n662, u0_u0_n663, u0_u0_n664, u0_u0_n665, u0_u0_n666, u0_u0_n667, 
       u0_u0_n668, u0_u0_n669, u0_u0_n670, u0_u0_n671, u0_u0_n672, u0_u0_n673, u0_u0_n674, u0_u0_n675, u0_u0_n676, 
       u0_u0_n677, u0_u0_n678, u0_u0_n679, u0_u0_n680, u0_u0_n681, u0_u0_n682, u0_u0_n683, u0_u0_n684, u0_u0_n685, 
       u0_u0_n686, u0_u0_n687, u0_u0_n688, u0_u0_n689, u0_u0_n690, u0_u0_n691, u0_u0_n692, u0_u0_n693, u0_u0_n694, 
       u0_u0_n695, u0_u0_n696, u0_u0_n697, u0_u0_n698, u0_u0_n699, u0_u0_n700, u0_u0_n701, u0_u0_n702, u0_u0_n703, 
       u0_u0_n704, u0_u0_n705, u0_u0_n706, u0_u0_n707, u0_u0_n708, u0_u0_n709, u0_u0_n710, u0_u0_n711, u0_u0_n712, 
       u0_u0_n713, u0_u0_n714, u0_u0_n715, u0_u0_n716, u0_u0_n717, u0_u0_n718, u0_u0_n719, u0_u0_n720, u0_u0_n721, 
       u0_u0_n722, u0_u0_n723, u0_u0_n724, u0_u0_n725, u0_u0_n726, u0_u0_n727, u0_u0_n728, u0_u0_n729, u0_u0_n730, 
       u0_u0_n731, u0_u0_n732, u0_u0_n733, u0_u0_n734, u0_u0_n735, u0_u0_n736, u0_u0_n737, u0_u0_n738, u0_u0_n739, 
       u0_u0_n740, u0_u0_n741, u0_u0_n742, u0_u0_n743, u0_u0_n744, u0_u0_n745, u0_u0_n746, u0_u0_n747, u0_u0_n748, 
       u0_u0_n749, u0_u0_n750, u0_u0_n751, u0_u0_n752, u0_u0_n753, u0_u0_n754, u0_u0_n755, u0_u0_n756, u0_u0_n757, 
       u0_u0_n758, u0_u0_n759, u0_u0_n760, u0_u0_n761, u0_u0_n762, u0_u0_n763, u0_u0_n764, u0_u0_n765, u0_u0_n766, 
       u0_u0_n767, u0_u0_n768, u0_u0_n769, u0_u0_n770, u0_u0_n771, u0_u0_n772, u0_u0_n773, u0_u0_n774, u0_u0_n775, 
       u0_u0_n776, u0_u0_n777, u0_u0_n778, u0_u0_n779, u0_u0_n780, u0_u0_n781, u0_u0_n782, u0_u0_n783, u0_u0_n784, 
       u0_u0_n785, u0_u0_n786, u0_u0_n787, u0_u0_n788, u0_u0_n789, u0_u0_n790, u0_u0_n791, u0_u0_n792, u0_u0_n793, 
       u0_u0_n794, u0_u0_n795, u0_u0_n796, u0_u0_n797, u0_u0_n798, u0_u0_n799, u0_u0_n800, u0_u0_n801, u0_u0_n802, 
       u0_u0_n803, u0_u0_n804, u0_u0_n805, u0_u0_n806, u0_u0_n807, u0_u0_n808, u0_u0_n809, u0_u0_n810, u0_u0_n811, 
       u0_u0_n812, u0_u0_n813, u0_u0_n814, u0_u0_n815, u0_u0_n816, u0_u0_n817, u0_u0_n818, u0_u0_n819, u0_u0_n820, 
       u0_u0_n821, u0_u0_n822, u0_u0_n823, u0_u0_n824, u0_u0_n825, u0_u0_n826, u0_u0_n827, u0_u0_n828, u0_u0_n829, 
       u0_u0_n830, u0_u0_n831, u0_u0_n832, u0_u0_n833, u0_u0_n834, u0_u0_n835, u0_u0_n836, u0_u0_n837, u0_u0_n838, 
       u0_u0_n839, u0_u0_n840, u0_u0_n841, u0_u0_n842, u0_u0_n843, u0_u0_n844, u0_u0_n845, u0_u0_n846, u0_u0_n847, 
       u0_u0_n848, u0_u0_n849, u0_u0_n850, u0_u0_n851, u0_u0_n852, u0_u0_n853, u0_u0_n854, u0_u0_n855, u0_u0_n856, 
       u0_u0_n857, u0_u0_n858, u0_u0_n859, u0_u0_n860, u0_u0_n861, u0_u0_n862, u0_u0_n863, u0_u0_n864, u0_u0_n865, 
       u0_u0_n866, u0_u0_n867, u0_u0_n868, u0_u0_n869, u0_u0_n870, u0_u0_n871, u0_u0_n872, u0_u0_n873, u0_u0_n874, 
       u0_u0_n875, u0_u0_n876, u0_u0_n877, u0_u0_n878,  u0_u0_n879;
  XNOR2_X1 u0_U181 (.ZN( u0_n226 ) , .B( u0_subword_31 ) , .A( w0_31 ) );
  XNOR2_X1 u0_U215 (.ZN( u0_n164 ) , .B( u0_n262 ) , .A( u0_n3 ) );
  XNOR2_X1 u0_U260 (.ZN( u0_n230 ) , .B( u0_subword_29 ) , .A( w0_29 ) );
  XNOR2_X1 u0_U287 (.ZN( u0_n236 ) , .A( u0_subword_26 ) , .B( w0_26 ) );
  XOR2_X1 u0_U296 (.Z( u0_n80 ) , .A( u0_n82 ) , .B( w3_26 ) );
  XNOR2_X1 u0_U3 (.A( u0_n11 ) , .ZN( u0_n172 ) , .B( u0_n242 ) );
  XOR2_X1 u0_U356 (.Z( u0_n1 ) , .A( u0_n226 ) , .B( u0_rcon_31 ) );
  XOR2_X1 u0_U358 (.A( u0_n228 ) , .Z( u0_n3 ) , .B( u0_rcon_30 ) );
  XOR2_X1 u0_U360 (.A( u0_n230 ) , .Z( u0_n5 ) , .B( u0_rcon_29 ) );
  XOR2_X1 u0_U364 (.A( u0_n234 ) , .Z( u0_n9 ) , .B( u0_rcon_27 ) );
  XOR2_X1 u0_U366 (.Z( u0_n11 ) , .A( u0_n236 ) , .B( u0_rcon_26 ) );
  XNOR2_X1 u0_U4 (.A( u0_n172 ) , .B( u0_n244 ) , .ZN( u0_n82 ) );
  XNOR2_X1 u0_U6 (.ZN( u0_n234 ) , .B( u0_subword_27 ) , .A( w0_27 ) );
  XNOR2_X1 u0_U7 (.ZN( u0_n228 ) , .B( u0_subword_30 ) , .A( w0_30 ) );
  INV_X1 u0_u0_U10 (.A( u0_u0_n1 ) , .ZN( u0_u0_n440 ) );
  AOI22_X1 u0_u0_U100 (.A2( u0_u0_n787 ) , .ZN( u0_u0_n788 ) , .B2( u0_u0_n836 ) , .A1( u0_u0_n839 ) , .B1( u0_u0_n867 ) );
  INV_X1 u0_u0_U101 (.A( u0_u0_n767 ) , .ZN( u0_u0_n835 ) );
  NOR2_X1 u0_u0_U102 (.ZN( u0_u0_n653 ) , .A1( u0_u0_n859 ) , .A2( u0_u0_n872 ) );
  INV_X1 u0_u0_U103 (.A( u0_u0_n759 ) , .ZN( u0_u0_n873 ) );
  OAI21_X1 u0_u0_U104 (.A( u0_u0_n439 ) , .B1( u0_u0_n758 ) , .ZN( u0_u0_n759 ) , .B2( u0_u0_n872 ) );
  NOR4_X1 u0_u0_U105 (.A4( u0_u0_n671 ) , .A3( u0_u0_n672 ) , .A2( u0_u0_n673 ) , .A1( u0_u0_n674 ) , .ZN( u0_u0_n682 ) );
  NOR4_X1 u0_u0_U106 (.A4( u0_u0_n667 ) , .A3( u0_u0_n668 ) , .A2( u0_u0_n669 ) , .A1( u0_u0_n670 ) , .ZN( u0_u0_n683 ) );
  NOR2_X1 u0_u0_U107 (.ZN( u0_u0_n738 ) , .A2( u0_u0_n837 ) , .A1( u0_u0_n850 ) );
  OR4_X1 u0_u0_U108 (.ZN( u0_u0_n472 ) , .A4( u0_u0_n524 ) , .A3( u0_u0_n535 ) , .A2( u0_u0_n584 ) , .A1( u0_u0_n717 ) );
  OR4_X1 u0_u0_U109 (.A4( u0_u0_n524 ) , .A2( u0_u0_n525 ) , .A1( u0_u0_n526 ) , .ZN( u0_u0_n528 ) , .A3( u0_u0_n826 ) );
  NAND2_X2 u0_u0_U11 (.A1( u0_u0_n455 ) , .A2( u0_u0_n466 ) , .ZN( u0_u0_n797 ) );
  OR4_X1 u0_u0_U110 (.A4( u0_u0_n688 ) , .A3( u0_u0_n689 ) , .A2( u0_u0_n690 ) , .A1( u0_u0_n691 ) , .ZN( u0_u0_n696 ) );
  OR4_X1 u0_u0_U111 (.A4( u0_u0_n572 ) , .A3( u0_u0_n573 ) , .A2( u0_u0_n574 ) , .ZN( u0_u0_n578 ) , .A1( u0_u0_n671 ) );
  OR4_X1 u0_u0_U112 (.ZN( u0_u0_n498 ) , .A4( u0_u0_n540 ) , .A2( u0_u0_n553 ) , .A1( u0_u0_n565 ) , .A3( u0_u0_n638 ) );
  INV_X1 u0_u0_U113 (.A( u0_u0_n442 ) , .ZN( u0_u0_n843 ) );
  OR3_X1 u0_u0_U114 (.A3( u0_u0_n512 ) , .A2( u0_u0_n513 ) , .A1( u0_u0_n514 ) , .ZN( u0_u0_n517 ) );
  INV_X1 u0_u0_U115 (.A( u0_u0_n469 ) , .ZN( u0_u0_n868 ) );
  OAI21_X1 u0_u0_U116 (.ZN( u0_u0_n469 ) , .B1( u0_u0_n814 ) , .A( u0_u0_n839 ) , .B2( u0_u0_n856 ) );
  AOI221_X1 u0_u0_U117 (.A( u0_u0_n718 ) , .B2( u0_u0_n719 ) , .ZN( u0_u0_n725 ) , .C1( u0_u0_n837 ) , .B1( u0_u0_n844 ) , .C2( u0_u0_n867 ) );
  OR2_X1 u0_u0_U118 (.A2( u0_u0_n716 ) , .A1( u0_u0_n717 ) , .ZN( u0_u0_n718 ) );
  NOR4_X1 u0_u0_U119 (.A4( u0_u0_n504 ) , .A3( u0_u0_n505 ) , .A2( u0_u0_n506 ) , .ZN( u0_u0_n507 ) , .A1( u0_u0_n533 ) );
  NAND2_X1 u0_u0_U12 (.A1( u0_u0_n457 ) , .A2( u0_u0_n477 ) , .ZN( u0_u0_n821 ) );
  NOR4_X1 u0_u0_U120 (.A4( u0_u0_n823 ) , .A3( u0_u0_n824 ) , .A2( u0_u0_n825 ) , .A1( u0_u0_n826 ) , .ZN( u0_u0_n827 ) );
  INV_X1 u0_u0_U121 (.A( u0_u0_n754 ) , .ZN( u0_u0_n867 ) );
  AOI221_X1 u0_u0_U122 (.C1( u0_u0_n444 ) , .A( u0_u0_n769 ) , .ZN( u0_u0_n779 ) , .C2( u0_u0_n815 ) , .B2( u0_u0_n840 ) , .B1( u0_u0_n870 ) );
  INV_X1 u0_u0_U123 (.A( u0_u0_n766 ) , .ZN( u0_u0_n840 ) );
  INV_X1 u0_u0_U124 (.A( u0_u0_n735 ) , .ZN( u0_u0_n844 ) );
  INV_X1 u0_u0_U125 (.A( u0_u0_n795 ) , .ZN( u0_u0_n837 ) );
  AOI211_X1 u0_u0_U126 (.B( u0_u0_n595 ) , .A( u0_u0_n596 ) , .ZN( u0_u0_n602 ) , .C2( u0_u0_n816 ) , .C1( u0_u0_n838 ) );
  AOI211_X1 u0_u0_U127 (.A( u0_u0_n502 ) , .ZN( u0_u0_n509 ) , .B( u0_u0_n807 ) , .C2( u0_u0_n844 ) , .C1( u0_u0_n856 ) );
  OAI221_X1 u0_u0_U128 (.A( u0_u0_n732 ) , .C2( u0_u0_n733 ) , .B2( u0_u0_n734 ) , .B1( u0_u0_n735 ) , .ZN( u0_u0_n742 ) , .C1( u0_u0_n822 ) );
  AOI22_X1 u0_u0_U129 (.ZN( u0_u0_n732 ) , .B1( u0_u0_n837 ) , .A2( u0_u0_n843 ) , .A1( u0_u0_n867 ) , .B2( u0_u0_n870 ) );
  NAND2_X1 u0_u0_U13 (.A2( u0_u0_n459 ) , .A1( u0_u0_n461 ) , .ZN( u0_u0_n811 ) );
  NOR4_X1 u0_u0_U130 (.A4( u0_u0_n645 ) , .A3( u0_u0_n646 ) , .A2( u0_u0_n647 ) , .A1( u0_u0_n648 ) , .ZN( u0_u0_n649 ) );
  AOI21_X1 u0_u0_U131 (.ZN( u0_u0_n645 ) , .B2( u0_u0_n754 ) , .A( u0_u0_n793 ) , .B1( u0_u0_n817 ) );
  NOR4_X1 u0_u0_U132 (.A4( u0_u0_n798 ) , .A3( u0_u0_n799 ) , .A2( u0_u0_n800 ) , .A1( u0_u0_n801 ) , .ZN( u0_u0_n802 ) );
  OAI21_X1 u0_u0_U133 (.A( u0_u0_n792 ) , .B2( u0_u0_n793 ) , .B1( u0_u0_n794 ) , .ZN( u0_u0_n800 ) );
  OAI221_X1 u0_u0_U134 (.A( u0_u0_n788 ) , .C2( u0_u0_n789 ) , .B2( u0_u0_n790 ) , .B1( u0_u0_n791 ) , .ZN( u0_u0_n801 ) , .C1( u0_u0_n818 ) );
  NOR3_X1 u0_u0_U135 (.ZN( u0_u0_n496 ) , .A1( u0_u0_n787 ) , .A2( u0_u0_n855 ) , .A3( u0_u0_n867 ) );
  AOI211_X1 u0_u0_U136 (.B( u0_u0_n750 ) , .A( u0_u0_n751 ) , .ZN( u0_u0_n764 ) , .C1( u0_u0_n837 ) , .C2( u0_u0_n858 ) );
  AOI211_X1 u0_u0_U137 (.B( u0_u0_n700 ) , .A( u0_u0_n701 ) , .ZN( u0_u0_n711 ) , .C2( u0_u0_n836 ) , .C1( u0_u0_n856 ) );
  AOI211_X1 u0_u0_U138 (.C2( u0_u0_n444 ) , .B( u0_u0_n730 ) , .A( u0_u0_n731 ) , .ZN( u0_u0_n744 ) , .C1( u0_u0_n848 ) );
  INV_X1 u0_u0_U139 (.A( u0_u0_n793 ) , .ZN( u0_u0_n850 ) );
  NOR3_X1 u0_u0_U14 (.A3( u0_u0_n171 ) , .A1( u0_u0_n622 ) , .A2( u0_u0_n623 ) , .ZN( u0_u0_n624 ) );
  NOR2_X1 u0_u0_U140 (.ZN( u0_u0_n672 ) , .A1( u0_u0_n733 ) , .A2( u0_u0_n808 ) );
  NOR2_X1 u0_u0_U141 (.ZN( u0_u0_n576 ) , .A1( u0_u0_n733 ) , .A2( u0_u0_n811 ) );
  NOR2_X1 u0_u0_U142 (.ZN( u0_u0_n538 ) , .A2( u0_u0_n754 ) , .A1( u0_u0_n755 ) );
  NOR2_X1 u0_u0_U143 (.ZN( u0_u0_n512 ) , .A2( u0_u0_n733 ) , .A1( u0_u0_n767 ) );
  BUF_X2 u0_u0_U144 (.Z( u0_u0_n441 ) , .A( u0_u0_n796 ) );
  CLKBUF_X3 u0_u0_U145 (.Z( u0_u0_n442 ) , .A( u0_u0_n703 ) );
  NOR2_X1 u0_u0_U146 (.ZN( u0_u0_n667 ) , .A1( u0_u0_n734 ) , .A2( u0_u0_n795 ) );
  NOR2_X1 u0_u0_U147 (.ZN( u0_u0_n515 ) , .A1( u0_u0_n734 ) , .A2( u0_u0_n784 ) );
  NOR2_X1 u0_u0_U148 (.ZN( u0_u0_n673 ) , .A1( u0_u0_n755 ) , .A2( u0_u0_n820 ) );
  INV_X1 u0_u0_U149 (.A( u0_u0_n819 ) , .ZN( u0_u0_n838 ) );
  NOR3_X1 u0_u0_U15 (.A3( u0_u0_n438 ) , .A1( u0_u0_n781 ) , .ZN( u0_u0_n804 ) , .A2( u0_u0_n806 ) );
  NOR2_X1 u0_u0_U150 (.A2( u0_u0_n442 ) , .ZN( u0_u0_n668 ) , .A1( u0_u0_n734 ) );
  NOR2_X1 u0_u0_U151 (.ZN( u0_u0_n669 ) , .A1( u0_u0_n734 ) , .A2( u0_u0_n790 ) );
  NOR2_X1 u0_u0_U152 (.ZN( u0_u0_n513 ) , .A1( u0_u0_n817 ) , .A2( u0_u0_n822 ) );
  NOR2_X1 u0_u0_U153 (.ZN( u0_u0_n661 ) , .A1( u0_u0_n795 ) , .A2( u0_u0_n820 ) );
  NOR2_X1 u0_u0_U154 (.ZN( u0_u0_n551 ) , .A1( u0_u0_n754 ) , .A2( u0_u0_n819 ) );
  NOR2_X1 u0_u0_U155 (.ZN( u0_u0_n636 ) , .A1( u0_u0_n752 ) , .A2( u0_u0_n820 ) );
  NOR2_X1 u0_u0_U156 (.A1( u0_u0_n754 ) , .ZN( u0_u0_n772 ) , .A2( u0_u0_n808 ) );
  NOR2_X1 u0_u0_U157 (.A1( u0_u0_n442 ) , .ZN( u0_u0_n775 ) , .A2( u0_u0_n820 ) );
  INV_X1 u0_u0_U158 (.A( u0_u0_n752 ) , .ZN( u0_u0_n839 ) );
  INV_X1 u0_u0_U159 (.A( u0_u0_n755 ) , .ZN( u0_u0_n847 ) );
  OR4_X1 u0_u0_U16 (.A4( u0_u0_n586 ) , .A3( u0_u0_n587 ) , .A2( u0_u0_n588 ) , .A1( u0_u0_n589 ) , .ZN( u0_u0_n590 ) );
  NOR2_X1 u0_u0_U160 (.ZN( u0_u0_n621 ) , .A1( u0_u0_n790 ) , .A2( u0_u0_n820 ) );
  NOR2_X1 u0_u0_U161 (.ZN( u0_u0_n635 ) , .A2( u0_u0_n733 ) , .A1( u0_u0_n790 ) );
  NOR2_X1 u0_u0_U162 (.ZN( u0_u0_n716 ) , .A1( u0_u0_n767 ) , .A2( u0_u0_n768 ) );
  NOR2_X1 u0_u0_U163 (.A2( u0_u0_n442 ) , .ZN( u0_u0_n600 ) , .A1( u0_u0_n733 ) );
  NOR2_X1 u0_u0_U164 (.ZN( u0_u0_n620 ) , .A1( u0_u0_n767 ) , .A2( u0_u0_n817 ) );
  AOI21_X1 u0_u0_U165 (.B1( u0_u0_n631 ) , .ZN( u0_u0_n633 ) , .A( u0_u0_n768 ) , .B2( u0_u0_n819 ) );
  AOI21_X1 u0_u0_U166 (.ZN( u0_u0_n597 ) , .B2( u0_u0_n768 ) , .A( u0_u0_n790 ) , .B1( u0_u0_n817 ) );
  AOI21_X1 u0_u0_U167 (.ZN( u0_u0_n521 ) , .A( u0_u0_n734 ) , .B1( u0_u0_n755 ) , .B2( u0_u0_n808 ) );
  AOI21_X1 u0_u0_U168 (.ZN( u0_u0_n545 ) , .B2( u0_u0_n817 ) , .A( u0_u0_n819 ) , .B1( u0_u0_n820 ) );
  INV_X1 u0_u0_U169 (.A( u0_u0_n808 ) , .ZN( u0_u0_n848 ) );
  NOR2_X1 u0_u0_U17 (.A2( u0_u0_n22 ) , .A1( u0_u0_n590 ) , .ZN( u0_u0_n591 ) );
  AOI21_X1 u0_u0_U170 (.ZN( u0_u0_n546 ) , .A( u0_u0_n768 ) , .B2( u0_u0_n784 ) , .B1( u0_u0_n822 ) );
  NOR2_X1 u0_u0_U171 (.ZN( u0_u0_n574 ) , .A1( u0_u0_n734 ) , .A2( u0_u0_n767 ) );
  AOI21_X1 u0_u0_U172 (.B1( u0_u0_n692 ) , .ZN( u0_u0_n693 ) , .A( u0_u0_n733 ) , .B2( u0_u0_n766 ) );
  NOR2_X1 u0_u0_U173 (.A2( u0_u0_n442 ) , .ZN( u0_u0_n572 ) , .A1( u0_u0_n768 ) );
  INV_X1 u0_u0_U174 (.A( u0_u0_n733 ) , .ZN( u0_u0_n857 ) );
  INV_X1 u0_u0_U175 (.A( u0_u0_n734 ) , .ZN( u0_u0_n872 ) );
  AOI21_X1 u0_u0_U176 (.B2( u0_u0_n442 ) , .ZN( u0_u0_n577 ) , .B1( u0_u0_n811 ) , .A( u0_u0_n817 ) );
  NOR2_X1 u0_u0_U177 (.ZN( u0_u0_n527 ) , .A1( u0_u0_n795 ) , .A2( u0_u0_n817 ) );
  AOI21_X1 u0_u0_U178 (.ZN( u0_u0_n695 ) , .B2( u0_u0_n754 ) , .B1( u0_u0_n768 ) , .A( u0_u0_n811 ) );
  AOI21_X1 u0_u0_U179 (.B2( u0_u0_n442 ) , .ZN( u0_u0_n484 ) , .A( u0_u0_n754 ) , .B1( u0_u0_n784 ) );
  NOR3_X1 u0_u0_U18 (.A3( u0_u0_n805 ) , .A2( u0_u0_n806 ) , .A1( u0_u0_n807 ) , .ZN( u0_u0_n830 ) );
  INV_X1 u0_u0_U180 (.A( u0_u0_n817 ) , .ZN( u0_u0_n859 ) );
  INV_X1 u0_u0_U181 (.A( u0_u0_n811 ) , .ZN( u0_u0_n846 ) );
  INV_X1 u0_u0_U182 (.A( u0_u0_n768 ) , .ZN( u0_u0_n870 ) );
  OAI21_X1 u0_u0_U183 (.A( u0_u0_n704 ) , .ZN( u0_u0_n708 ) , .B2( u0_u0_n755 ) , .B1( u0_u0_n809 ) );
  OAI21_X1 u0_u0_U184 (.ZN( u0_u0_n704 ) , .B2( u0_u0_n838 ) , .B1( u0_u0_n843 ) , .A( u0_u0_n864 ) );
  NOR2_X1 u0_u0_U185 (.ZN( u0_u0_n476 ) , .A2( u0_u0_n784 ) , .A1( u0_u0_n820 ) );
  NAND2_X1 u0_u0_U186 (.A2( u0_u0_n767 ) , .A1( u0_u0_n811 ) , .ZN( u0_u0_n815 ) );
  BUF_X1 u0_u0_U187 (.Z( u0_u0_n443 ) , .A( u0_u0_n818 ) );
  INV_X1 u0_u0_U188 (.A( u0_u0_n790 ) , .ZN( u0_u0_n851 ) );
  INV_X1 u0_u0_U189 (.A( u0_u0_n822 ) , .ZN( u0_u0_n849 ) );
  NOR3_X1 u0_u0_U19 (.ZN( u0_u0_n604 ) , .A1( u0_u0_n614 ) , .A3( u0_u0_n728 ) , .A2( u0_u0_n747 ) );
  OAI22_X1 u0_u0_U190 (.B2( u0_u0_n755 ) , .B1( u0_u0_n756 ) , .A1( u0_u0_n757 ) , .ZN( u0_u0_n761 ) , .A2( u0_u0_n811 ) );
  NOR3_X1 u0_u0_U191 (.ZN( u0_u0_n757 ) , .A2( u0_u0_n858 ) , .A1( u0_u0_n867 ) , .A3( u0_u0_n869 ) );
  NOR2_X1 u0_u0_U192 (.ZN( u0_u0_n756 ) , .A2( u0_u0_n857 ) , .A1( u0_u0_n864 ) );
  AND2_X1 u0_u0_U193 (.ZN( u0_u0_n753 ) , .A1( u0_u0_n789 ) , .A2( u0_u0_n791 ) );
  AND2_X1 u0_u0_U194 (.ZN( u0_u0_n737 ) , .A1( u0_u0_n784 ) , .A2( u0_u0_n790 ) );
  AOI221_X1 u0_u0_U195 (.A( u0_u0_n503 ) , .ZN( u0_u0_n508 ) , .B2( u0_u0_n848 ) , .C1( u0_u0_n851 ) , .C2( u0_u0_n864 ) , .B1( u0_u0_n866 ) );
  AOI221_X1 u0_u0_U196 (.A( u0_u0_n687 ) , .ZN( u0_u0_n698 ) , .B2( u0_u0_n845 ) , .C1( u0_u0_n847 ) , .C2( u0_u0_n866 ) , .B1( u0_u0_n869 ) );
  INV_X1 u0_u0_U197 (.A( u0_u0_n686 ) , .ZN( u0_u0_n845 ) );
  OAI221_X1 u0_u0_U198 (.A( u0_u0_n702 ) , .ZN( u0_u0_n709 ) , .C2( u0_u0_n789 ) , .C1( u0_u0_n790 ) , .B1( u0_u0_n791 ) , .B2( u0_u0_n811 ) );
  AOI22_X1 u0_u0_U199 (.ZN( u0_u0_n702 ) , .A1( u0_u0_n835 ) , .B2( u0_u0_n848 ) , .A2( u0_u0_n869 ) , .B1( u0_u0_n872 ) );
  NOR3_X1 u0_u0_U20 (.A1( u0_u0_n1 ) , .ZN( u0_u0_n510 ) , .A2( u0_u0_n685 ) , .A3( u0_u0_n782 ) );
  OAI222_X1 u0_u0_U200 (.A2( u0_u0_n675 ) , .ZN( u0_u0_n680 ) , .B1( u0_u0_n752 ) , .B2( u0_u0_n789 ) , .C2( u0_u0_n793 ) , .C1( u0_u0_n820 ) , .A1( u0_u0_n822 ) );
  NAND2_X1 u0_u0_U201 (.A2( u0_u0_n454 ) , .A1( u0_u0_n466 ) , .ZN( u0_u0_n733 ) );
  NAND2_X1 u0_u0_U202 (.A2( u0_u0_n454 ) , .A1( u0_u0_n458 ) , .ZN( u0_u0_n734 ) );
  NAND2_X1 u0_u0_U203 (.A2( u0_u0_n455 ) , .A1( u0_u0_n458 ) , .ZN( u0_u0_n768 ) );
  NAND2_X1 u0_u0_U204 (.A2( u0_u0_n454 ) , .A1( u0_u0_n470 ) , .ZN( u0_u0_n820 ) );
  NAND2_X1 u0_u0_U205 (.A2( u0_u0_n466 ) , .A1( u0_u0_n471 ) , .ZN( u0_u0_n785 ) );
  NAND2_X1 u0_u0_U206 (.A1( u0_u0_n453 ) , .A2( u0_u0_n471 ) , .ZN( u0_u0_n754 ) );
  NOR2_X1 u0_u0_U207 (.ZN( u0_u0_n471 ) , .A2( u0_u0_n852 ) , .A1( u0_u0_n853 ) );
  NAND2_X1 u0_u0_U208 (.A2( u0_u0_n467 ) , .A1( u0_u0_n468 ) , .ZN( u0_u0_n752 ) );
  NAND2_X1 u0_u0_U209 (.A1( u0_u0_n468 ) , .A2( u0_u0_n478 ) , .ZN( u0_u0_n793 ) );
  NOR3_X1 u0_u0_U21 (.A2( u0_u0_n613 ) , .A1( u0_u0_n614 ) , .ZN( u0_u0_n652 ) , .A3( u0_u0_n727 ) );
  NOR4_X1 u0_u0_U210 (.A4( u0_u0_n739 ) , .A3( u0_u0_n740 ) , .A2( u0_u0_n741 ) , .A1( u0_u0_n742 ) , .ZN( u0_u0_n743 ) );
  NOR4_X1 u0_u0_U211 (.A4( u0_u0_n706 ) , .A3( u0_u0_n707 ) , .A2( u0_u0_n708 ) , .A1( u0_u0_n709 ) , .ZN( u0_u0_n710 ) );
  NOR4_X1 u0_u0_U212 (.A3( u0_u0_n760 ) , .A2( u0_u0_n761 ) , .A1( u0_u0_n762 ) , .ZN( u0_u0_n763 ) , .A4( u0_u0_n873 ) );
  NOR2_X1 u0_u0_U213 (.ZN( u0_u0_n477 ) , .A1( u0_u0_n831 ) , .A2( w3_17 ) );
  AOI221_X1 u0_u0_U214 (.A( u0_u0_n786 ) , .ZN( u0_u0_n803 ) , .C2( u0_u0_n842 ) , .B2( u0_u0_n843 ) , .B1( u0_u0_n869 ) , .C1( u0_u0_n870 ) );
  NAND4_X1 u0_u0_U215 (.ZN( u0_subword_25 ) , .A4( u0_u0_n601 ) , .A3( u0_u0_n602 ) , .A2( u0_u0_n603 ) , .A1( u0_u0_n604 ) );
  NOR4_X1 u0_u0_U216 (.A4( u0_u0_n597 ) , .A3( u0_u0_n598 ) , .A2( u0_u0_n599 ) , .A1( u0_u0_n600 ) , .ZN( u0_u0_n601 ) );
  NAND4_X1 u0_u0_U217 (.ZN( u0_subword_24 ) , .A4( u0_u0_n507 ) , .A3( u0_u0_n508 ) , .A2( u0_u0_n509 ) , .A1( u0_u0_n510 ) );
  AOI222_X1 u0_u0_U218 (.B2( u0_u0_n644 ) , .ZN( u0_u0_n650 ) , .B1( u0_u0_n846 ) , .A1( u0_u0_n847 ) , .C2( u0_u0_n851 ) , .C1( u0_u0_n867 ) , .A2( u0_u0_n869 ) );
  AND2_X1 u0_u0_U219 (.ZN( u0_u0_n453 ) , .A2( w3_22 ) , .A1( w3_23 ) );
  NOR3_X1 u0_u0_U22 (.A3( u0_u0_n746 ) , .A2( u0_u0_n747 ) , .A1( u0_u0_n748 ) , .ZN( u0_u0_n765 ) );
  NAND4_X1 u0_u0_U220 (.ZN( u0_subword_31 ) , .A4( u0_u0_n827 ) , .A3( u0_u0_n828 ) , .A2( u0_u0_n829 ) , .A1( u0_u0_n830 ) );
  AOI222_X1 u0_u0_U221 (.C2( u0_u0_n814 ) , .B2( u0_u0_n815 ) , .A2( u0_u0_n816 ) , .ZN( u0_u0_n828 ) , .C1( u0_u0_n837 ) , .A1( u0_u0_n844 ) , .B1( u0_u0_n858 ) );
  INV_X1 u0_u0_U222 (.ZN( u0_u0_n853 ) , .A( w3_21 ) );
  NAND4_X1 u0_u0_U223 (.A4( u0_u0_n697 ) , .A3( u0_u0_n698 ) , .A1( u0_u0_n699 ) , .ZN( u0_u0_n781 ) , .A2( u0_u0_n876 ) );
  NAND2_X2 u0_u0_U224 (.A2( u0_u0_n470 ) , .A1( u0_u0_n471 ) , .ZN( u0_u0_n817 ) );
  NAND2_X1 u0_u0_U225 (.A2( u0_u0_n447 ) , .A1( u0_u0_n458 ) , .ZN( u0_u0_n796 ) );
  AOI222_X1 u0_u0_U226 (.ZN( u0_u0_n780 ) , .A1( u0_u0_n835 ) , .C1( u0_u0_n839 ) , .B2( u0_u0_n846 ) , .A2( u0_u0_n855 ) , .B1( u0_u0_n865 ) , .C2( u0_u0_n877 ) );
  OAI21_X1 u0_u0_U227 (.ZN( u0_u0_n736 ) , .A( u0_u0_n838 ) , .B2( u0_u0_n857 ) , .B1( u0_u0_n877 ) );
  AOI222_X1 u0_u0_U228 (.ZN( u0_u0_n569 ) , .B1( u0_u0_n835 ) , .C1( u0_u0_n846 ) , .A2( u0_u0_n848 ) , .A1( u0_u0_n859 ) , .B2( u0_u0_n867 ) , .C2( u0_u0_n877 ) );
  OAI21_X1 u0_u0_U229 (.ZN( u0_u0_n792 ) , .A( u0_u0_n844 ) , .B1( u0_u0_n867 ) , .B2( u0_u0_n877 ) );
  NOR3_X1 u0_u0_U23 (.A3( u0_u0_n727 ) , .A1( u0_u0_n728 ) , .ZN( u0_u0_n745 ) , .A2( u0_u0_n746 ) );
  NAND4_X1 u0_u0_U230 (.A4( u0_u0_n479 ) , .A3( u0_u0_n480 ) , .A2( u0_u0_n481 ) , .A1( u0_u0_n482 ) , .ZN( u0_u0_n684 ) );
  NOR4_X1 u0_u0_U231 (.ZN( u0_u0_n479 ) , .A2( u0_u0_n527 ) , .A4( u0_u0_n600 ) , .A1( u0_u0_n615 ) , .A3( u0_u0_n635 ) );
  NAND2_X1 u0_u0_U232 (.A2( u0_u0_n467 ) , .A1( u0_u0_n477 ) , .ZN( u0_u0_n703 ) );
  NAND2_X1 u0_u0_U233 (.A2( u0_u0_n460 ) , .A1( u0_u0_n461 ) , .ZN( u0_u0_n735 ) );
  NAND2_X1 u0_u0_U234 (.A1( u0_u0_n460 ) , .A2( u0_u0_n467 ) , .ZN( u0_u0_n818 ) );
  NOR2_X1 u0_u0_U235 (.ZN( u0_u0_n461 ) , .A1( u0_u0_n833 ) , .A2( w3_19 ) );
  NAND2_X2 u0_u0_U236 (.A1( u0_u0_n457 ) , .A2( u0_u0_n460 ) , .ZN( u0_u0_n819 ) );
  AOI211_X1 u0_u0_U237 (.B( u0_u0_n812 ) , .A( u0_u0_n813 ) , .ZN( u0_u0_n829 ) , .C1( u0_u0_n847 ) , .C2( u0_u0_n855 ) );
  NOR2_X1 u0_u0_U238 (.A1( u0_u0_n684 ) , .ZN( u0_u0_n699 ) , .A2( u0_u0_n812 ) );
  OAI222_X1 u0_u0_U239 (.B1( u0_u0_n442 ) , .ZN( u0_u0_n623 ) , .C1( u0_u0_n729 ) , .C2( u0_u0_n752 ) , .B2( u0_u0_n791 ) , .A2( u0_u0_n797 ) , .A1( u0_u0_n821 ) );
  NOR2_X1 u0_u0_U24 (.ZN( u0_u0_n581 ) , .A1( u0_u0_n628 ) , .A2( u0_u0_n750 ) );
  AOI21_X1 u0_u0_U240 (.A( u0_u0_n676 ) , .B1( u0_u0_n677 ) , .ZN( u0_u0_n678 ) , .B2( u0_u0_n860 ) );
  AOI21_X1 u0_u0_U241 (.B1( u0_u0_n445 ) , .ZN( u0_u0_n516 ) , .B2( u0_u0_n675 ) , .A( u0_u0_n735 ) );
  INV_X1 u0_u0_U242 (.A( u0_u0_n675 ) , .ZN( u0_u0_n869 ) );
  NOR2_X1 u0_u0_U243 (.ZN( u0_u0_n658 ) , .A1( u0_u0_n675 ) , .A2( u0_u0_n819 ) );
  NOR2_X1 u0_u0_U244 (.ZN( u0_u0_n533 ) , .A1( u0_u0_n675 ) , .A2( u0_u0_n784 ) );
  AOI21_X1 u0_u0_U245 (.ZN( u0_u0_n483 ) , .A( u0_u0_n675 ) , .B1( u0_u0_n755 ) , .B2( u0_u0_n811 ) );
  NOR2_X1 u0_u0_U246 (.ZN( u0_u0_n608 ) , .A1( u0_u0_n675 ) , .A2( u0_u0_n808 ) );
  NOR2_X1 u0_u0_U247 (.ZN( u0_u0_n634 ) , .A2( u0_u0_n675 ) , .A1( u0_u0_n790 ) );
  NOR2_X1 u0_u0_U248 (.ZN( u0_u0_n587 ) , .A1( u0_u0_n675 ) , .A2( u0_u0_n793 ) );
  NAND2_X2 u0_u0_U249 (.A1( u0_u0_n458 ) , .A2( u0_u0_n471 ) , .ZN( u0_u0_n675 ) );
  NOR2_X1 u0_u0_U25 (.ZN( u0_u0_n501 ) , .A1( u0_u0_n684 ) , .A2( u0_u0_n700 ) );
  NAND4_X1 u0_u0_U250 (.A4( u0_u0_n541 ) , .A3( u0_u0_n542 ) , .A2( u0_u0_n543 ) , .A1( u0_u0_n544 ) , .ZN( u0_u0_n628 ) );
  OAI222_X1 u0_u0_U251 (.A2( u0_u0_n445 ) , .B2( u0_u0_n713 ) , .ZN( u0_u0_n714 ) , .C2( u0_u0_n729 ) , .B1( u0_u0_n752 ) , .A1( u0_u0_n811 ) , .C1( u0_u0_n819 ) );
  NOR2_X1 u0_u0_U252 (.ZN( u0_u0_n524 ) , .A1( u0_u0_n713 ) , .A2( u0_u0_n793 ) );
  NOR2_X1 u0_u0_U253 (.ZN( u0_u0_n526 ) , .A2( u0_u0_n713 ) , .A1( u0_u0_n819 ) );
  NOR2_X1 u0_u0_U254 (.A2( u0_u0_n713 ) , .A1( u0_u0_n767 ) , .ZN( u0_u0_n799 ) );
  NOR2_X1 u0_u0_U255 (.A2( u0_u0_n713 ) , .A1( u0_u0_n755 ) , .ZN( u0_u0_n776 ) );
  NOR2_X1 u0_u0_U256 (.ZN( u0_u0_n523 ) , .A1( u0_u0_n713 ) , .A2( u0_u0_n808 ) );
  NOR2_X1 u0_u0_U257 (.ZN( u0_u0_n688 ) , .A2( u0_u0_n713 ) , .A1( u0_u0_n822 ) );
  OAI22_X1 u0_u0_U258 (.ZN( u0_u0_n489 ) , .A1( u0_u0_n713 ) , .B2( u0_u0_n790 ) , .A2( u0_u0_n811 ) , .B1( u0_u0_n817 ) );
  NOR2_X1 u0_u0_U259 (.ZN( u0_u0_n549 ) , .A2( u0_u0_n713 ) , .A1( u0_u0_n790 ) );
  NOR2_X1 u0_u0_U26 (.ZN( u0_u0_n712 ) , .A2( u0_u0_n781 ) , .A1( u0_u0_n805 ) );
  NOR2_X1 u0_u0_U260 (.ZN( u0_u0_n585 ) , .A2( u0_u0_n713 ) , .A1( u0_u0_n735 ) );
  NOR2_X1 u0_u0_U261 (.ZN( u0_u0_n535 ) , .A1( u0_u0_n713 ) , .A2( u0_u0_n784 ) );
  NOR2_X1 u0_u0_U262 (.ZN( u0_u0_n674 ) , .A2( u0_u0_n713 ) , .A1( u0_u0_n795 ) );
  AOI222_X1 u0_u0_U263 (.ZN( u0_u0_n531 ) , .A1( u0_u0_n839 ) , .B2( u0_u0_n842 ) , .C1( u0_u0_n849 ) , .C2( u0_u0_n855 ) , .A2( u0_u0_n857 ) , .B1( u0_u0_n870 ) );
  AOI222_X1 u0_u0_U264 (.ZN( u0_u0_n612 ) , .A1( u0_u0_n835 ) , .C2( u0_u0_n842 ) , .B1( u0_u0_n847 ) , .A2( u0_u0_n860 ) , .B2( u0_u0_n865 ) , .C1( u0_u0_n872 ) );
  NOR3_X1 u0_u0_U265 (.ZN( u0_u0_n446 ) , .A2( u0_u0_n841 ) , .A3( u0_u0_n842 ) , .A1( u0_u0_n851 ) );
  NAND2_X1 u0_u0_U266 (.ZN( u0_u0_n619 ) , .A2( u0_u0_n842 ) , .A1( u0_u0_n877 ) );
  OAI22_X1 u0_u0_U267 (.A1( u0_u0_n445 ) , .B2( u0_u0_n784 ) , .B1( u0_u0_n785 ) , .ZN( u0_u0_n786 ) , .A2( u0_u0_n819 ) );
  NAND4_X1 u0_u0_U268 (.A4( u0_u0_n499 ) , .A3( u0_u0_n500 ) , .A1( u0_u0_n501 ) , .ZN( u0_u0_n807 ) , .A2( u0_u0_n871 ) );
  AOI21_X1 u0_u0_U269 (.ZN( u0_u0_n575 ) , .B1( u0_u0_n755 ) , .B2( u0_u0_n767 ) , .A( u0_u0_n785 ) );
  AOI222_X1 u0_u0_U27 (.ZN( u0_u0_n666 ) , .A2( u0_u0_n844 ) , .B1( u0_u0_n846 ) , .C2( u0_u0_n850 ) , .A1( u0_u0_n864 ) , .C1( u0_u0_n867 ) , .B2( u0_u0_n874 ) );
  NAND2_X1 u0_u0_U270 (.ZN( u0_u0_n719 ) , .A1( u0_u0_n733 ) , .A2( u0_u0_n785 ) );
  OAI22_X1 u0_u0_U271 (.B1( u0_u0_n496 ) , .ZN( u0_u0_n497 ) , .A1( u0_u0_n692 ) , .A2( u0_u0_n768 ) , .B2( u0_u0_n822 ) );
  NOR2_X1 u0_u0_U272 (.ZN( u0_u0_n662 ) , .A1( u0_u0_n752 ) , .A2( u0_u0_n785 ) );
  NOR2_X1 u0_u0_U273 (.A2( u0_u0_n442 ) , .A1( u0_u0_n785 ) , .ZN( u0_u0_n825 ) );
  NOR2_X1 u0_u0_U274 (.ZN( u0_u0_n514 ) , .A2( u0_u0_n785 ) , .A1( u0_u0_n790 ) );
  NOR2_X1 u0_u0_U275 (.ZN( u0_u0_n607 ) , .A2( u0_u0_n785 ) , .A1( u0_u0_n808 ) );
  NOR2_X1 u0_u0_U276 (.ZN( u0_u0_n617 ) , .A2( u0_u0_n785 ) , .A1( u0_u0_n811 ) );
  NOR2_X1 u0_u0_U277 (.ZN( u0_u0_n552 ) , .A2( u0_u0_n785 ) , .A1( u0_u0_n819 ) );
  INV_X1 u0_u0_U278 (.A( u0_u0_n785 ) , .ZN( u0_u0_n855 ) );
  AOI21_X1 u0_u0_U279 (.ZN( u0_u0_n646 ) , .B2( u0_u0_n752 ) , .A( u0_u0_n797 ) , .B1( u0_u0_n808 ) );
  INV_X1 u0_u0_U28 (.A( u0_u0_n653 ) , .ZN( u0_u0_n874 ) );
  AOI21_X1 u0_u0_U280 (.A( u0_u0_n738 ) , .ZN( u0_u0_n739 ) , .B2( u0_u0_n785 ) , .B1( u0_u0_n797 ) );
  NAND4_X1 u0_u0_U281 (.A4( u0_u0_n554 ) , .A3( u0_u0_n555 ) , .A2( u0_u0_n556 ) , .A1( u0_u0_n557 ) , .ZN( u0_u0_n750 ) );
  AOI21_X1 u0_u0_U282 (.ZN( u0_u0_n520 ) , .A( u0_u0_n784 ) , .B2( u0_u0_n797 ) , .B1( u0_u0_n817 ) );
  AOI21_X1 u0_u0_U283 (.B2( u0_u0_n768 ) , .ZN( u0_u0_n769 ) , .A( u0_u0_n793 ) , .B1( u0_u0_n797 ) );
  AOI21_X1 u0_u0_U284 (.ZN( u0_u0_n456 ) , .B2( u0_u0_n797 ) , .A( u0_u0_n808 ) , .B1( u0_u0_n820 ) );
  INV_X1 u0_u0_U285 (.A( u0_u0_n797 ) , .ZN( u0_u0_n856 ) );
  NOR2_X1 u0_u0_U286 (.A2( u0_u0_n442 ) , .ZN( u0_u0_n721 ) , .A1( u0_u0_n797 ) );
  NOR2_X1 u0_u0_U287 (.ZN( u0_u0_n563 ) , .A1( u0_u0_n797 ) , .A2( u0_u0_n819 ) );
  NOR2_X1 u0_u0_U288 (.ZN( u0_u0_n589 ) , .A1( u0_u0_n797 ) , .A2( u0_u0_n822 ) );
  NOR2_X1 u0_u0_U289 (.ZN( u0_u0_n550 ) , .A2( u0_u0_n790 ) , .A1( u0_u0_n797 ) );
  NOR4_X1 u0_u0_U29 (.ZN( u0_u0_n491 ) , .A2( u0_u0_n539 ) , .A1( u0_u0_n564 ) , .A3( u0_u0_n637 ) , .A4( u0_u0_n723 ) );
  INV_X1 u0_u0_U290 (.ZN( u0_u0_n444 ) , .A( u0_u0_n820 ) );
  INV_X1 u0_u0_U291 (.A( u0_u0_n444 ) , .ZN( u0_u0_n445 ) );
  NOR4_X1 u0_u0_U292 (.A2( u0_u0_n497 ) , .A1( u0_u0_n498 ) , .ZN( u0_u0_n499 ) , .A3( u0_u0_n586 ) , .A4( u0_u0_n618 ) );
  INV_X1 u0_u0_U293 (.ZN( u0_u0_n832 ) , .A( w3_17 ) );
  AOI21_X1 u0_u0_U294 (.B1( u0_u0_n445 ) , .ZN( u0_u0_n595 ) , .B2( u0_u0_n705 ) , .A( u0_u0_n822 ) );
  AOI21_X1 u0_u0_U295 (.B1( u0_u0_n705 ) , .ZN( u0_u0_n706 ) , .A( u0_u0_n737 ) , .B2( u0_u0_n768 ) );
  INV_X1 u0_u0_U296 (.A( u0_u0_n705 ) , .ZN( u0_u0_n858 ) );
  AOI21_X1 u0_u0_U297 (.ZN( u0_u0_n448 ) , .A( u0_u0_n705 ) , .B1( u0_u0_n738 ) , .B2( u0_u0_n755 ) );
  NOR2_X1 u0_u0_U298 (.ZN( u0_u0_n583 ) , .A2( u0_u0_n705 ) , .A1( u0_u0_n819 ) );
  NOR2_X1 u0_u0_U299 (.ZN( u0_u0_n689 ) , .A2( u0_u0_n705 ) , .A1( u0_u0_n808 ) );
  OR4_X1 u0_u0_U3 (.ZN( u0_u0_n1 ) , .A4( u0_u0_n451 ) , .A3( u0_u0_n452 ) , .A2( u0_u0_n522 ) , .A1( u0_u0_n547 ) );
  NOR4_X1 u0_u0_U30 (.ZN( u0_u0_n485 ) , .A1( u0_u0_n526 ) , .A4( u0_u0_n563 ) , .A3( u0_u0_n588 ) , .A2( u0_u0_n636 ) );
  NOR2_X1 u0_u0_U300 (.A2( u0_u0_n442 ) , .ZN( u0_u0_n547 ) , .A1( u0_u0_n705 ) );
  NAND2_X1 u0_u0_U301 (.A1( u0_u0_n705 ) , .A2( u0_u0_n734 ) , .ZN( u0_u0_n787 ) );
  NAND2_X2 u0_u0_U302 (.A1( u0_u0_n447 ) , .A2( u0_u0_n466 ) , .ZN( u0_u0_n705 ) );
  NOR4_X1 u0_u0_U303 (.A3( u0_u0_n679 ) , .A1( u0_u0_n680 ) , .ZN( u0_u0_n681 ) , .A4( u0_u0_n720 ) , .A2( u0_u0_n863 ) );
  INV_X1 u0_u0_U304 (.A( u0_u0_n678 ) , .ZN( u0_u0_n863 ) );
  NOR2_X1 u0_u0_U305 (.ZN( u0_u0_n459 ) , .A1( u0_u0_n831 ) , .A2( u0_u0_n832 ) );
  AOI21_X1 u0_u0_U306 (.ZN( u0_u0_n504 ) , .A( u0_u0_n729 ) , .B2( u0_u0_n767 ) , .B1( u0_u0_n819 ) );
  OAI22_X1 u0_u0_U307 (.ZN( u0_u0_n495 ) , .A1( u0_u0_n729 ) , .B2( u0_u0_n733 ) , .B1( u0_u0_n735 ) , .A2( u0_u0_n784 ) );
  NOR2_X1 u0_u0_U308 (.ZN( u0_u0_n717 ) , .A2( u0_u0_n729 ) , .A1( u0_u0_n795 ) );
  NOR2_X1 u0_u0_U309 (.ZN( u0_u0_n534 ) , .A2( u0_u0_n729 ) , .A1( u0_u0_n808 ) );
  NOR4_X1 u0_u0_U31 (.ZN( u0_u0_n462 ) , .A2( u0_u0_n523 ) , .A1( u0_u0_n549 ) , .A3( u0_u0_n585 ) , .A4( u0_u0_n621 ) );
  NOR2_X1 u0_u0_U310 (.ZN( u0_u0_n532 ) , .A1( u0_u0_n729 ) , .A2( u0_u0_n755 ) );
  NOR2_X1 u0_u0_U311 (.ZN( u0_u0_n615 ) , .A2( u0_u0_n729 ) , .A1( u0_u0_n822 ) );
  NOR2_X1 u0_u0_U312 (.A2( u0_u0_n442 ) , .ZN( u0_u0_n638 ) , .A1( u0_u0_n729 ) );
  NOR2_X1 u0_u0_U313 (.ZN( u0_u0_n540 ) , .A1( u0_u0_n729 ) , .A2( u0_u0_n793 ) );
  NOR2_X1 u0_u0_U314 (.ZN( u0_u0_n539 ) , .A2( u0_u0_n729 ) , .A1( u0_u0_n735 ) );
  INV_X1 u0_u0_U315 (.A( u0_u0_n729 ) , .ZN( u0_u0_n860 ) );
  NAND2_X2 u0_u0_U316 (.A1( u0_u0_n447 ) , .A2( u0_u0_n470 ) , .ZN( u0_u0_n713 ) );
  NAND2_X2 u0_u0_U317 (.A1( u0_u0_n455 ) , .A2( u0_u0_n470 ) , .ZN( u0_u0_n729 ) );
  AOI211_X1 u0_u0_U318 (.C1( u0_u0_n439 ) , .C2( u0_u0_n444 ) , .A( u0_u0_n594 ) , .ZN( u0_u0_n603 ) , .B( u0_u0_n627 ) );
  NOR3_X1 u0_u0_U319 (.A2( u0_u0_n627 ) , .A3( u0_u0_n628 ) , .ZN( u0_u0_n642 ) , .A1( u0_u0_n730 ) );
  OR3_X1 u0_u0_U32 (.ZN( u0_u0_n452 ) , .A1( u0_u0_n534 ) , .A3( u0_u0_n583 ) , .A2( u0_u0_n879 ) );
  AOI21_X1 u0_u0_U320 (.B2( u0_u0_n443 ) , .ZN( u0_u0_n599 ) , .B1( u0_u0_n755 ) , .A( u0_u0_n797 ) );
  AOI21_X1 u0_u0_U321 (.A( u0_u0_n817 ) , .B2( u0_u0_n818 ) , .B1( u0_u0_n819 ) , .ZN( u0_u0_n824 ) );
  AOI21_X1 u0_u0_U322 (.A( u0_u0_n443 ) , .ZN( u0_u0_n655 ) , .B1( u0_u0_n734 ) , .B2( u0_u0_n768 ) );
  NOR2_X1 u0_u0_U323 (.A2( u0_u0_n818 ) , .A1( u0_u0_n820 ) , .ZN( u0_u0_n826 ) );
  NOR2_X1 u0_u0_U324 (.A2( u0_u0_n443 ) , .A1( u0_u0_n675 ) , .ZN( u0_u0_n771 ) );
  NOR2_X1 u0_u0_U325 (.ZN( u0_u0_n584 ) , .A1( u0_u0_n713 ) , .A2( u0_u0_n818 ) );
  NOR2_X1 u0_u0_U326 (.ZN( u0_u0_n671 ) , .A1( u0_u0_n785 ) , .A2( u0_u0_n818 ) );
  NAND2_X2 u0_u0_U327 (.A2( u0_u0_n460 ) , .A1( u0_u0_n478 ) , .ZN( u0_u0_n784 ) );
  NOR2_X1 u0_u0_U328 (.A1( u0_u0_n705 ) , .ZN( u0_u0_n773 ) , .A2( u0_u0_n818 ) );
  NOR2_X1 u0_u0_U329 (.A2( u0_u0_n443 ) , .ZN( u0_u0_n660 ) , .A1( u0_u0_n733 ) );
  INV_X1 u0_u0_U33 (.A( u0_u0_n619 ) , .ZN( u0_u0_n879 ) );
  NOR2_X1 u0_u0_U330 (.A2( u0_u0_n443 ) , .ZN( u0_u0_n637 ) , .A1( u0_u0_n729 ) );
  INV_X1 u0_u0_U331 (.A( u0_u0_n818 ) , .ZN( u0_u0_n841 ) );
  NAND2_X2 u0_u0_U332 (.A1( u0_u0_n457 ) , .A2( u0_u0_n459 ) , .ZN( u0_u0_n767 ) );
  NOR2_X1 u0_u0_U333 (.ZN( u0_u0_n478 ) , .A1( w3_18 ) , .A2( w3_19 ) );
  AOI21_X1 u0_u0_U334 (.A( u0_u0_n441 ) , .ZN( u0_u0_n647 ) , .B1( u0_u0_n686 ) , .B2( u0_u0_n822 ) );
  NAND2_X2 u0_u0_U335 (.A1( u0_u0_n453 ) , .A2( u0_u0_n455 ) , .ZN( u0_u0_n810 ) );
  AOI21_X1 u0_u0_U336 (.B2( u0_u0_n441 ) , .A( u0_u0_n795 ) , .B1( u0_u0_n797 ) , .ZN( u0_u0_n798 ) );
  OAI22_X1 u0_u0_U337 (.B1( u0_u0_n441 ) , .ZN( u0_u0_n701 ) , .A2( u0_u0_n735 ) , .A1( u0_u0_n785 ) , .B2( u0_u0_n822 ) );
  AOI21_X1 u0_u0_U338 (.B2( u0_u0_n441 ) , .ZN( u0_u0_n503 ) , .A( u0_u0_n784 ) , .B1( u0_u0_n809 ) );
  AOI21_X1 u0_u0_U339 (.B1( u0_u0_n441 ) , .ZN( u0_u0_n632 ) , .B2( u0_u0_n675 ) , .A( u0_u0_n795 ) );
  NOR4_X1 u0_u0_U34 (.A1( u0_u0_n537 ) , .ZN( u0_u0_n542 ) , .A2( u0_u0_n660 ) , .A4( u0_u0_n674 ) , .A3( u0_u0_n770 ) );
  NAND2_X2 u0_u0_U340 (.A1( u0_u0_n461 ) , .A2( u0_u0_n468 ) , .ZN( u0_u0_n755 ) );
  AOI21_X1 u0_u0_U341 (.B2( u0_u0_n441 ) , .ZN( u0_u0_n570 ) , .B1( u0_u0_n729 ) , .A( u0_u0_n784 ) );
  NAND2_X2 u0_u0_U342 (.A1( u0_u0_n457 ) , .A2( u0_u0_n468 ) , .ZN( u0_u0_n795 ) );
  AOI21_X1 u0_u0_U343 (.B2( u0_u0_n441 ) , .ZN( u0_u0_n449 ) , .B1( u0_u0_n794 ) , .A( u0_u0_n819 ) );
  NOR2_X1 u0_u0_U344 (.A2( u0_u0_n441 ) , .ZN( u0_u0_n670 ) , .A1( u0_u0_n790 ) );
  NOR2_X1 u0_u0_U345 (.A2( u0_u0_n441 ) , .ZN( u0_u0_n561 ) , .A1( u0_u0_n755 ) );
  NOR2_X1 u0_u0_U346 (.A2( u0_u0_n441 ) , .ZN( u0_u0_n565 ) , .A1( u0_u0_n808 ) );
  NOR2_X1 u0_u0_U347 (.A1( u0_u0_n441 ) , .A2( u0_u0_n443 ) , .ZN( u0_u0_n690 ) );
  NOR2_X1 u0_u0_U348 (.A1( u0_u0_n441 ) , .ZN( u0_u0_n648 ) , .A2( u0_u0_n793 ) );
  NAND2_X2 u0_u0_U349 (.A1( u0_u0_n453 ) , .A2( u0_u0_n454 ) , .ZN( u0_u0_n791 ) );
  NOR4_X1 u0_u0_U35 (.A4( u0_u0_n547 ) , .A3( u0_u0_n548 ) , .A2( u0_u0_n549 ) , .ZN( u0_u0_n556 ) , .A1( u0_u0_n694 ) );
  NOR2_X1 u0_u0_U350 (.A2( u0_u0_n441 ) , .ZN( u0_u0_n548 ) , .A1( u0_u0_n767 ) );
  INV_X1 u0_u0_U351 (.A( u0_u0_n796 ) , .ZN( u0_u0_n877 ) );
  NOR2_X1 u0_u0_U352 (.ZN( u0_u0_n586 ) , .A2( u0_u0_n703 ) , .A1( u0_u0_n796 ) );
  NOR2_X1 u0_u0_U353 (.ZN( u0_u0_n467 ) , .A1( u0_u0_n834 ) , .A2( w3_18 ) );
  AOI221_X1 u0_u0_U354 (.A( u0_u0_n582 ) , .ZN( u0_u0_n593 ) , .B2( u0_u0_n836 ) , .C2( u0_u0_n848 ) , .B1( u0_u0_n859 ) , .C1( u0_u0_n865 ) );
  NOR2_X1 u0_u0_U355 (.ZN( u0_u0_n457 ) , .A1( u0_u0_n833 ) , .A2( u0_u0_n834 ) );
  INV_X1 u0_u0_U356 (.ZN( u0_u0_n834 ) , .A( w3_19 ) );
  NAND2_X2 u0_u0_U357 (.A1( u0_u0_n459 ) , .A2( u0_u0_n478 ) , .ZN( u0_u0_n790 ) );
  INV_X1 u0_u0_U358 (.ZN( u0_u0_n833 ) , .A( w3_18 ) );
  AOI222_X1 u0_u0_U359 (.ZN( u0_u0_n611 ) , .B2( u0_u0_n677 ) , .B1( u0_u0_n758 ) , .C2( u0_u0_n836 ) , .A1( u0_u0_n838 ) , .A2( u0_u0_n866 ) , .C1( u0_u0_n867 ) );
  NOR4_X1 u0_u0_U36 (.A4( u0_u0_n583 ) , .A3( u0_u0_n584 ) , .A2( u0_u0_n585 ) , .ZN( u0_u0_n592 ) , .A1( u0_u0_n689 ) );
  AOI222_X1 u0_u0_U360 (.ZN( u0_u0_n519 ) , .C1( u0_u0_n837 ) , .B2( u0_u0_n842 ) , .A2( u0_u0_n848 ) , .C2( u0_u0_n866 ) , .B1( u0_u0_n867 ) , .A1( u0_u0_n870 ) );
  AOI221_X1 u0_u0_U361 (.A( u0_u0_n489 ) , .ZN( u0_u0_n494 ) , .B1( u0_u0_n836 ) , .C2( u0_u0_n849 ) , .C1( u0_u0_n857 ) , .B2( u0_u0_n866 ) );
  NOR2_X1 u0_u0_U362 (.ZN( u0_u0_n794 ) , .A2( u0_u0_n866 ) , .A1( u0_u0_n872 ) );
  INV_X1 u0_u0_U363 (.A( u0_u0_n791 ) , .ZN( u0_u0_n866 ) );
  OAI22_X1 u0_u0_U364 (.ZN( u0_u0_n643 ) , .A1( u0_u0_n705 ) , .B2( u0_u0_n733 ) , .A2( u0_u0_n767 ) , .B1( u0_u0_n821 ) );
  OAI22_X1 u0_u0_U365 (.A1( u0_u0_n729 ) , .ZN( u0_u0_n731 ) , .B2( u0_u0_n755 ) , .B1( u0_u0_n817 ) , .A2( u0_u0_n821 ) );
  AOI21_X1 u0_u0_U366 (.ZN( u0_u0_n505 ) , .B1( u0_u0_n686 ) , .A( u0_u0_n817 ) , .B2( u0_u0_n821 ) );
  AOI21_X1 u0_u0_U367 (.A( u0_u0_n445 ) , .B2( u0_u0_n821 ) , .B1( u0_u0_n822 ) , .ZN( u0_u0_n823 ) );
  OAI22_X1 u0_u0_U368 (.A1( u0_u0_n445 ) , .ZN( u0_u0_n630 ) , .B1( u0_u0_n675 ) , .B2( u0_u0_n752 ) , .A2( u0_u0_n821 ) );
  NOR2_X1 u0_u0_U369 (.A2( u0_u0_n441 ) , .ZN( u0_u0_n605 ) , .A1( u0_u0_n821 ) );
  NOR3_X1 u0_u0_U37 (.ZN( u0_u0_n555 ) , .A2( u0_u0_n657 ) , .A1( u0_u0_n673 ) , .A3( u0_u0_n776 ) );
  NOR2_X1 u0_u0_U370 (.ZN( u0_u0_n537 ) , .A2( u0_u0_n785 ) , .A1( u0_u0_n821 ) );
  NOR2_X1 u0_u0_U371 (.ZN( u0_u0_n525 ) , .A2( u0_u0_n705 ) , .A1( u0_u0_n821 ) );
  NAND2_X2 u0_u0_U372 (.A1( u0_u0_n461 ) , .A2( u0_u0_n477 ) , .ZN( u0_u0_n808 ) );
  NOR2_X1 u0_u0_U373 (.A1( u0_u0_n675 ) , .ZN( u0_u0_n694 ) , .A2( u0_u0_n821 ) );
  NOR2_X1 u0_u0_U374 (.ZN( u0_u0_n564 ) , .A1( u0_u0_n713 ) , .A2( u0_u0_n821 ) );
  NAND2_X2 u0_u0_U375 (.A1( u0_u0_n459 ) , .A2( u0_u0_n467 ) , .ZN( u0_u0_n749 ) );
  NOR2_X1 u0_u0_U376 (.ZN( u0_u0_n691 ) , .A1( u0_u0_n734 ) , .A2( u0_u0_n821 ) );
  INV_X1 u0_u0_U377 (.A( u0_u0_n821 ) , .ZN( u0_u0_n836 ) );
  NAND2_X1 u0_u0_U378 (.ZN( u0_u0_n677 ) , .A1( u0_u0_n811 ) , .A2( u0_u0_n821 ) );
  NOR2_X1 u0_u0_U379 (.ZN( u0_u0_n460 ) , .A1( u0_u0_n832 ) , .A2( w3_16 ) );
  AOI211_X1 u0_u0_U38 (.B( u0_u0_n545 ) , .A( u0_u0_n546 ) , .ZN( u0_u0_n557 ) , .C2( u0_u0_n844 ) , .C1( u0_u0_n856 ) );
  NOR2_X1 u0_u0_U380 (.ZN( u0_u0_n468 ) , .A2( w3_16 ) , .A1( w3_17 ) );
  INV_X1 u0_u0_U381 (.ZN( u0_u0_n831 ) , .A( w3_16 ) );
  AOI211_X1 u0_u0_U382 (.A( u0_u0_n643 ) , .ZN( u0_u0_n651 ) , .B( u0_u0_n748 ) , .C2( u0_u0_n844 ) , .C1( u0_u0_n859 ) );
  NAND4_X1 u0_u0_U383 (.A4( u0_u0_n639 ) , .A3( u0_u0_n640 ) , .A2( u0_u0_n641 ) , .A1( u0_u0_n642 ) , .ZN( u0_u0_n748 ) );
  AOI21_X1 u0_u0_U384 (.ZN( u0_u0_n582 ) , .B2( u0_u0_n729 ) , .B1( u0_u0_n753 ) , .A( u0_u0_n790 ) );
  NAND2_X2 u0_u0_U385 (.A2( u0_u0_n447 ) , .A1( u0_u0_n453 ) , .ZN( u0_u0_n789 ) );
  NOR2_X1 u0_u0_U386 (.ZN( u0_u0_n466 ) , .A1( u0_u0_n854 ) , .A2( w3_23 ) );
  INV_X1 u0_u0_U387 (.ZN( u0_u0_n862 ) , .A( w3_23 ) );
  NOR2_X1 u0_u0_U388 (.ZN( u0_u0_n447 ) , .A2( w3_20 ) , .A1( w3_21 ) );
  NOR2_X1 u0_u0_U389 (.ZN( u0_u0_n454 ) , .A1( u0_u0_n852 ) , .A2( w3_21 ) );
  NOR4_X1 u0_u0_U39 (.A4( u0_u0_n550 ) , .A3( u0_u0_n551 ) , .A2( u0_u0_n552 ) , .A1( u0_u0_n553 ) , .ZN( u0_u0_n554 ) );
  OAI21_X1 u0_u0_U390 (.A( u0_u0_n736 ) , .B1( u0_u0_n737 ) , .ZN( u0_u0_n741 ) , .B2( u0_u0_n810 ) );
  OAI222_X1 u0_u0_U391 (.B2( u0_u0_n752 ) , .B1( u0_u0_n753 ) , .A2( u0_u0_n754 ) , .ZN( u0_u0_n762 ) , .C2( u0_u0_n810 ) , .C1( u0_u0_n819 ) , .A1( u0_u0_n822 ) );
  OAI22_X1 u0_u0_U392 (.B2( u0_u0_n808 ) , .B1( u0_u0_n809 ) , .A2( u0_u0_n810 ) , .A1( u0_u0_n811 ) , .ZN( u0_u0_n813 ) );
  OAI222_X1 u0_u0_U393 (.ZN( u0_u0_n511 ) , .C2( u0_u0_n631 ) , .B2( u0_u0_n653 ) , .B1( u0_u0_n752 ) , .A2( u0_u0_n753 ) , .C1( u0_u0_n810 ) , .A1( u0_u0_n811 ) );
  AOI21_X1 u0_u0_U394 (.ZN( u0_u0_n656 ) , .A( u0_u0_n784 ) , .B1( u0_u0_n797 ) , .B2( u0_u0_n810 ) );
  INV_X1 u0_u0_U395 (.A( u0_u0_n810 ) , .ZN( u0_u0_n864 ) );
  NOR2_X1 u0_u0_U396 (.ZN( u0_u0_n740 ) , .A2( u0_u0_n808 ) , .A1( u0_u0_n810 ) );
  NOR2_X1 u0_u0_U397 (.ZN( u0_u0_n490 ) , .A1( u0_u0_n793 ) , .A2( u0_u0_n810 ) );
  NOR2_X1 u0_u0_U398 (.ZN( u0_u0_n573 ) , .A1( u0_u0_n752 ) , .A2( u0_u0_n810 ) );
  AOI21_X1 u0_u0_U399 (.A( u0_u0_n442 ) , .ZN( u0_u0_n558 ) , .B1( u0_u0_n675 ) , .B2( u0_u0_n810 ) );
  OR4_X1 u0_u0_U4 (.A4( u0_u0_n448 ) , .A2( u0_u0_n449 ) , .A1( u0_u0_n450 ) , .ZN( u0_u0_n451 ) , .A3( u0_u0_n559 ) );
  AOI221_X1 u0_u0_U40 (.A( u0_u0_n495 ) , .ZN( u0_u0_n500 ) , .B2( u0_u0_n841 ) , .C2( u0_u0_n846 ) , .C1( u0_u0_n856 ) , .B1( u0_u0_n864 ) );
  NAND2_X1 u0_u0_U400 (.ZN( u0_u0_n758 ) , .A1( u0_u0_n768 ) , .A2( u0_u0_n810 ) );
  NOR2_X1 u0_u0_U401 (.ZN( u0_u0_n720 ) , .A1( u0_u0_n810 ) , .A2( u0_u0_n822 ) );
  NOR2_X1 u0_u0_U402 (.ZN( u0_u0_n562 ) , .A1( u0_u0_n767 ) , .A2( u0_u0_n810 ) );
  NOR2_X1 u0_u0_U403 (.ZN( u0_u0_n676 ) , .A1( u0_u0_n795 ) , .A2( u0_u0_n810 ) );
  NAND4_X1 u0_u0_U404 (.ZN( u0_subword_27 ) , .A2( u0_u0_n440 ) , .A4( u0_u0_n710 ) , .A3( u0_u0_n711 ) , .A1( u0_u0_n712 ) );
  OAI22_X1 u0_u0_U405 (.B2( u0_u0_n749 ) , .ZN( u0_u0_n751 ) , .A2( u0_u0_n767 ) , .B1( u0_u0_n785 ) , .A1( u0_u0_n797 ) );
  OAI22_X1 u0_u0_U406 (.B1( u0_u0_n441 ) , .ZN( u0_u0_n502 ) , .A2( u0_u0_n749 ) , .A1( u0_u0_n785 ) , .B2( u0_u0_n811 ) );
  NOR2_X1 u0_u0_U407 (.ZN( u0_u0_n522 ) , .A1( u0_u0_n713 ) , .A2( u0_u0_n749 ) );
  OAI22_X1 u0_u0_U408 (.ZN( u0_u0_n715 ) , .A2( u0_u0_n733 ) , .B2( u0_u0_n734 ) , .A1( u0_u0_n749 ) , .B1( u0_u0_n818 ) );
  NOR2_X1 u0_u0_U409 (.A2( u0_u0_n749 ) , .ZN( u0_u0_n774 ) , .A1( u0_u0_n817 ) );
  INV_X1 u0_u0_U41 (.A( u0_u0_n783 ) , .ZN( u0_u0_n871 ) );
  OAI22_X1 u0_u0_U410 (.B1( u0_u0_n446 ) , .ZN( u0_u0_n450 ) , .A2( u0_u0_n733 ) , .A1( u0_u0_n749 ) , .B2( u0_u0_n754 ) );
  NOR2_X1 u0_u0_U411 (.ZN( u0_u0_n553 ) , .A1( u0_u0_n705 ) , .A2( u0_u0_n749 ) );
  NOR2_X1 u0_u0_U412 (.ZN( u0_u0_n536 ) , .A2( u0_u0_n749 ) , .A1( u0_u0_n797 ) );
  NOR2_X1 u0_u0_U413 (.A2( u0_u0_n749 ) , .ZN( u0_u0_n760 ) , .A1( u0_u0_n810 ) );
  NOR2_X1 u0_u0_U414 (.A1( u0_u0_n675 ) , .ZN( u0_u0_n679 ) , .A2( u0_u0_n749 ) );
  NOR2_X1 u0_u0_U415 (.ZN( u0_u0_n723 ) , .A2( u0_u0_n729 ) , .A1( u0_u0_n749 ) );
  NOR2_X1 u0_u0_U416 (.ZN( u0_u0_n588 ) , .A1( u0_u0_n749 ) , .A2( u0_u0_n820 ) );
  INV_X1 u0_u0_U417 (.A( u0_u0_n749 ) , .ZN( u0_u0_n842 ) );
  NAND4_X1 u0_u0_U418 (.ZN( u0_subword_26 ) , .A4( u0_u0_n649 ) , .A3( u0_u0_n650 ) , .A1( u0_u0_n651 ) , .A2( u0_u0_n652 ) );
  OAI22_X1 u0_u0_U419 (.ZN( u0_u0_n594 ) , .A2( u0_u0_n752 ) , .B2( u0_u0_n767 ) , .A1( u0_u0_n768 ) , .B1( u0_u0_n789 ) );
  NOR2_X1 u0_u0_U42 (.ZN( u0_u0_n686 ) , .A2( u0_u0_n839 ) , .A1( u0_u0_n844 ) );
  NAND2_X1 u0_u0_U420 (.A1( u0_u0_n734 ) , .A2( u0_u0_n789 ) , .ZN( u0_u0_n816 ) );
  AOI21_X1 u0_u0_U421 (.ZN( u0_u0_n598 ) , .B1( u0_u0_n733 ) , .B2( u0_u0_n789 ) , .A( u0_u0_n795 ) );
  AOI21_X1 u0_u0_U422 (.ZN( u0_u0_n654 ) , .A( u0_u0_n767 ) , .B2( u0_u0_n789 ) , .B1( u0_u0_n797 ) );
  AOI21_X1 u0_u0_U423 (.ZN( u0_u0_n629 ) , .B1( u0_u0_n705 ) , .A( u0_u0_n784 ) , .B2( u0_u0_n789 ) );
  OAI22_X1 u0_u0_U424 (.ZN( u0_u0_n687 ) , .A1( u0_u0_n705 ) , .A2( u0_u0_n735 ) , .B2( u0_u0_n789 ) , .B1( u0_u0_n822 ) );
  NOR2_X1 u0_u0_U425 (.ZN( u0_u0_n657 ) , .A1( u0_u0_n789 ) , .A2( u0_u0_n793 ) );
  OAI21_X1 u0_u0_U426 (.A( u0_u0_n619 ) , .ZN( u0_u0_n622 ) , .B1( u0_u0_n631 ) , .B2( u0_u0_n789 ) );
  NOR2_X1 u0_u0_U427 (.ZN( u0_u0_n559 ) , .A2( u0_u0_n749 ) , .A1( u0_u0_n789 ) );
  NOR2_X1 u0_u0_U428 (.ZN( u0_u0_n616 ) , .A1( u0_u0_n789 ) , .A2( u0_u0_n821 ) );
  NOR2_X1 u0_u0_U429 (.A2( u0_u0_n442 ) , .ZN( u0_u0_n606 ) , .A1( u0_u0_n789 ) );
  NAND4_X1 u0_u0_U43 (.A4( u0_u0_n609 ) , .A3( u0_u0_n610 ) , .A2( u0_u0_n611 ) , .A1( u0_u0_n612 ) , .ZN( u0_u0_n727 ) );
  INV_X1 u0_u0_U430 (.A( u0_u0_n789 ) , .ZN( u0_u0_n865 ) );
  NOR2_X1 u0_u0_U431 (.ZN( u0_u0_n470 ) , .A2( w3_22 ) , .A1( w3_23 ) );
  NOR2_X1 u0_u0_U432 (.ZN( u0_u0_n458 ) , .A1( u0_u0_n862 ) , .A2( w3_22 ) );
  INV_X1 u0_u0_U433 (.ZN( u0_u0_n854 ) , .A( w3_22 ) );
  AOI21_X1 u0_u0_U434 (.A( u0_u0_n442 ) , .ZN( u0_u0_n506 ) , .B1( u0_u0_n713 ) , .B2( u0_u0_n791 ) );
  OAI22_X1 u0_u0_U435 (.ZN( u0_u0_n596 ) , .B1( u0_u0_n735 ) , .B2( u0_u0_n754 ) , .A2( u0_u0_n791 ) , .A1( u0_u0_n808 ) );
  NOR2_X1 u0_u0_U436 (.ZN( u0_u0_n659 ) , .A1( u0_u0_n767 ) , .A2( u0_u0_n791 ) );
  NAND3_X1 u0_u0_U437 (.ZN( u0_subword_30 ) , .A3( u0_u0_n802 ) , .A2( u0_u0_n803 ) , .A1( u0_u0_n804 ) );
  NAND3_X1 u0_u0_U438 (.ZN( u0_subword_29 ) , .A3( u0_u0_n763 ) , .A2( u0_u0_n764 ) , .A1( u0_u0_n765 ) );
  NAND3_X1 u0_u0_U439 (.ZN( u0_subword_28 ) , .A3( u0_u0_n743 ) , .A2( u0_u0_n744 ) , .A1( u0_u0_n745 ) );
  NOR4_X1 u0_u0_U44 (.A3( u0_u0_n606 ) , .A2( u0_u0_n607 ) , .A1( u0_u0_n608 ) , .ZN( u0_u0_n609 ) , .A4( u0_u0_n661 ) );
  NAND3_X1 u0_u0_U440 (.A3( u0_u0_n681 ) , .A2( u0_u0_n682 ) , .A1( u0_u0_n683 ) , .ZN( u0_u0_n812 ) );
  NAND3_X1 u0_u0_U441 (.ZN( u0_u0_n644 ) , .A3( u0_u0_n713 ) , .A2( u0_u0_n729 ) , .A1( u0_u0_n797 ) );
  NAND3_X1 u0_u0_U442 (.A3( u0_u0_n624 ) , .A2( u0_u0_n625 ) , .A1( u0_u0_n626 ) , .ZN( u0_u0_n730 ) );
  NAND3_X1 u0_u0_U443 (.A1( u0_u0_n591 ) , .A2( u0_u0_n592 ) , .A3( u0_u0_n593 ) , .ZN( u0_u0_n627 ) );
  NAND3_X1 u0_u0_U444 (.ZN( u0_u0_n571 ) , .A3( u0_u0_n686 ) , .A2( u0_u0_n755 ) , .A1( u0_u0_n790 ) );
  NAND3_X1 u0_u0_U445 (.A3( u0_u0_n529 ) , .A2( u0_u0_n530 ) , .A1( u0_u0_n531 ) , .ZN( u0_u0_n747 ) );
  NAND3_X1 u0_u0_U446 (.A3( u0_u0_n518 ) , .A1( u0_u0_n519 ) , .ZN( u0_u0_n614 ) , .A2( u0_u0_n875 ) );
  NAND3_X1 u0_u0_U447 (.A3( u0_u0_n473 ) , .A2( u0_u0_n474 ) , .A1( u0_u0_n475 ) , .ZN( u0_u0_n782 ) );
  NAND2_X1 u0_u0_U448 (.A2( u0_u0_n754 ) , .A1( u0_u0_n791 ) , .ZN( u0_u0_n814 ) );
  NOR2_X1 u0_u0_U449 (.A2( u0_u0_n443 ) , .ZN( u0_u0_n560 ) , .A1( u0_u0_n791 ) );
  NOR3_X1 u0_u0_U45 (.A1( u0_u0_n605 ) , .ZN( u0_u0_n610 ) , .A3( u0_u0_n669 ) , .A2( u0_u0_n775 ) );
  NOR2_X1 u0_u0_U450 (.ZN( u0_u0_n618 ) , .A1( u0_u0_n784 ) , .A2( u0_u0_n791 ) );
  NOR2_X1 u0_u0_U451 (.ZN( u0_u0_n722 ) , .A2( u0_u0_n749 ) , .A1( u0_u0_n791 ) );
  NOR2_X1 u0_u0_U452 (.ZN( u0_u0_n707 ) , .A2( u0_u0_n791 ) , .A1( u0_u0_n822 ) );
  NOR2_X1 u0_u0_U453 (.A1( u0_u0_n735 ) , .ZN( u0_u0_n770 ) , .A2( u0_u0_n791 ) );
  NOR2_X1 u0_u0_U454 (.ZN( u0_u0_n455 ) , .A1( u0_u0_n853 ) , .A2( w3_20 ) );
  INV_X1 u0_u0_U455 (.ZN( u0_u0_n852 ) , .A( w3_20 ) );
  NAND4_X1 u0_u0_U46 (.A4( u0_u0_n566 ) , .A3( u0_u0_n567 ) , .A2( u0_u0_n568 ) , .A1( u0_u0_n569 ) , .ZN( u0_u0_n613 ) );
  NOR4_X1 u0_u0_U47 (.ZN( u0_u0_n567 ) , .A1( u0_u0_n659 ) , .A3( u0_u0_n667 ) , .A4( u0_u0_n691 ) , .A2( u0_u0_n773 ) );
  NOR4_X1 u0_u0_U48 (.A4( u0_u0_n558 ) , .A3( u0_u0_n559 ) , .A2( u0_u0_n560 ) , .A1( u0_u0_n561 ) , .ZN( u0_u0_n568 ) );
  NOR4_X1 u0_u0_U49 (.A4( u0_u0_n562 ) , .A3( u0_u0_n563 ) , .A2( u0_u0_n564 ) , .A1( u0_u0_n565 ) , .ZN( u0_u0_n566 ) );
  OR3_X1 u0_u0_U5 (.ZN( u0_u0_n22 ) , .A3( u0_u0_n658 ) , .A1( u0_u0_n668 ) , .A2( u0_u0_n772 ) );
  NOR4_X1 u0_u0_U50 (.A4( u0_u0_n693 ) , .A3( u0_u0_n694 ) , .A2( u0_u0_n695 ) , .A1( u0_u0_n696 ) , .ZN( u0_u0_n697 ) );
  INV_X1 u0_u0_U51 (.A( u0_u0_n685 ) , .ZN( u0_u0_n876 ) );
  NOR4_X1 u0_u0_U52 (.A4( u0_u0_n532 ) , .A2( u0_u0_n533 ) , .A1( u0_u0_n534 ) , .ZN( u0_u0_n544 ) , .A3( u0_u0_n707 ) );
  NOR4_X1 u0_u0_U53 (.A4( u0_u0_n535 ) , .A3( u0_u0_n536 ) , .ZN( u0_u0_n543 ) , .A2( u0_u0_n690 ) , .A1( u0_u0_n799 ) );
  NOR4_X1 u0_u0_U54 (.A4( u0_u0_n538 ) , .A3( u0_u0_n539 ) , .A2( u0_u0_n540 ) , .ZN( u0_u0_n541 ) , .A1( u0_u0_n825 ) );
  NOR4_X1 u0_u0_U55 (.A4( u0_u0_n520 ) , .A3( u0_u0_n521 ) , .A2( u0_u0_n522 ) , .A1( u0_u0_n523 ) , .ZN( u0_u0_n530 ) );
  NOR4_X1 u0_u0_U56 (.A3( u0_u0_n527 ) , .A1( u0_u0_n528 ) , .ZN( u0_u0_n529 ) , .A2( u0_u0_n679 ) , .A4( u0_u0_n774 ) );
  NOR4_X1 u0_u0_U57 (.A4( u0_u0_n476 ) , .ZN( u0_u0_n482 ) , .A3( u0_u0_n562 ) , .A1( u0_u0_n740 ) , .A2( u0_u0_n760 ) );
  NOR4_X1 u0_u0_U58 (.ZN( u0_u0_n481 ) , .A1( u0_u0_n537 ) , .A3( u0_u0_n574 ) , .A4( u0_u0_n606 ) , .A2( u0_u0_n648 ) );
  NOR4_X1 u0_u0_U59 (.ZN( u0_u0_n480 ) , .A1( u0_u0_n512 ) , .A3( u0_u0_n550 ) , .A2( u0_u0_n589 ) , .A4( u0_u0_n721 ) );
  OR2_X1 u0_u0_U6 (.ZN( u0_u0_n171 ) , .A2( u0_u0_n620 ) , .A1( u0_u0_n621 ) );
  NOR4_X1 u0_u0_U60 (.A4( u0_u0_n635 ) , .A3( u0_u0_n636 ) , .A2( u0_u0_n637 ) , .A1( u0_u0_n638 ) , .ZN( u0_u0_n639 ) );
  NOR4_X1 u0_u0_U61 (.A4( u0_u0_n632 ) , .A3( u0_u0_n633 ) , .A2( u0_u0_n634 ) , .ZN( u0_u0_n640 ) , .A1( u0_u0_n670 ) );
  AOI211_X1 u0_u0_U62 (.B( u0_u0_n629 ) , .A( u0_u0_n630 ) , .ZN( u0_u0_n641 ) , .C2( u0_u0_n841 ) , .C1( u0_u0_n867 ) );
  NAND4_X1 u0_u0_U63 (.A4( u0_u0_n777 ) , .A3( u0_u0_n778 ) , .A2( u0_u0_n779 ) , .A1( u0_u0_n780 ) , .ZN( u0_u0_n806 ) );
  NOR3_X1 u0_u0_U64 (.A3( u0_u0_n770 ) , .A2( u0_u0_n771 ) , .A1( u0_u0_n772 ) , .ZN( u0_u0_n778 ) );
  NOR4_X1 u0_u0_U65 (.A4( u0_u0_n773 ) , .A3( u0_u0_n774 ) , .A2( u0_u0_n775 ) , .A1( u0_u0_n776 ) , .ZN( u0_u0_n777 ) );
  NAND4_X1 u0_u0_U66 (.A4( u0_u0_n663 ) , .A3( u0_u0_n664 ) , .A2( u0_u0_n665 ) , .A1( u0_u0_n666 ) , .ZN( u0_u0_n805 ) );
  NOR3_X1 u0_u0_U67 (.A3( u0_u0_n654 ) , .A2( u0_u0_n655 ) , .A1( u0_u0_n656 ) , .ZN( u0_u0_n665 ) );
  NOR3_X1 u0_u0_U68 (.A3( u0_u0_n657 ) , .A2( u0_u0_n658 ) , .A1( u0_u0_n659 ) , .ZN( u0_u0_n664 ) );
  NOR3_X1 u0_u0_U69 (.A3( u0_u0_n660 ) , .A2( u0_u0_n661 ) , .A1( u0_u0_n662 ) , .ZN( u0_u0_n663 ) );
  OR2_X1 u0_u0_U7 (.ZN( u0_u0_n438 ) , .A1( u0_u0_n782 ) , .A2( u0_u0_n783 ) );
  NOR4_X1 u0_u0_U70 (.A4( u0_u0_n515 ) , .A2( u0_u0_n516 ) , .A1( u0_u0_n517 ) , .ZN( u0_u0_n518 ) , .A3( u0_u0_n676 ) );
  INV_X1 u0_u0_U71 (.A( u0_u0_n511 ) , .ZN( u0_u0_n875 ) );
  NOR2_X1 u0_u0_U72 (.ZN( u0_u0_n809 ) , .A1( u0_u0_n859 ) , .A2( u0_u0_n865 ) );
  NAND4_X1 u0_u0_U73 (.A4( u0_u0_n491 ) , .A3( u0_u0_n492 ) , .A2( u0_u0_n493 ) , .A1( u0_u0_n494 ) , .ZN( u0_u0_n783 ) );
  NOR4_X1 u0_u0_U74 (.A4( u0_u0_n490 ) , .ZN( u0_u0_n493 ) , .A1( u0_u0_n572 ) , .A2( u0_u0_n587 ) , .A3( u0_u0_n608 ) );
  NOR4_X1 u0_u0_U75 (.ZN( u0_u0_n492 ) , .A1( u0_u0_n513 ) , .A2( u0_u0_n525 ) , .A4( u0_u0_n552 ) , .A3( u0_u0_n617 ) );
  NAND4_X1 u0_u0_U76 (.A4( u0_u0_n462 ) , .A3( u0_u0_n463 ) , .A2( u0_u0_n464 ) , .A1( u0_u0_n465 ) , .ZN( u0_u0_n685 ) );
  NOR3_X1 u0_u0_U77 (.ZN( u0_u0_n463 ) , .A3( u0_u0_n536 ) , .A1( u0_u0_n561 ) , .A2( u0_u0_n576 ) );
  AOI221_X1 u0_u0_U78 (.A( u0_u0_n456 ) , .ZN( u0_u0_n465 ) , .C2( u0_u0_n758 ) , .B1( u0_u0_n837 ) , .C1( u0_u0_n847 ) , .B2( u0_u0_n865 ) );
  NOR4_X1 u0_u0_U79 (.ZN( u0_u0_n464 ) , .A2( u0_u0_n515 ) , .A1( u0_u0_n605 ) , .A4( u0_u0_n634 ) , .A3( u0_u0_n716 ) );
  NAND2_X2 u0_u0_U8 (.A2( u0_u0_n477 ) , .A1( u0_u0_n478 ) , .ZN( u0_u0_n822 ) );
  NOR2_X1 u0_u0_U80 (.ZN( u0_u0_n766 ) , .A1( u0_u0_n838 ) , .A2( u0_u0_n839 ) );
  NOR2_X1 u0_u0_U81 (.ZN( u0_u0_n631 ) , .A2( u0_u0_n841 ) , .A1( u0_u0_n844 ) );
  NAND4_X1 u0_u0_U82 (.A4( u0_u0_n485 ) , .A3( u0_u0_n486 ) , .A2( u0_u0_n487 ) , .A1( u0_u0_n488 ) , .ZN( u0_u0_n700 ) );
  NOR3_X1 u0_u0_U83 (.ZN( u0_u0_n486 ) , .A2( u0_u0_n514 ) , .A3( u0_u0_n607 ) , .A1( u0_u0_n616 ) );
  NOR4_X1 u0_u0_U84 (.ZN( u0_u0_n487 ) , .A3( u0_u0_n538 ) , .A4( u0_u0_n551 ) , .A2( u0_u0_n573 ) , .A1( u0_u0_n722 ) );
  AOI211_X1 u0_u0_U85 (.B( u0_u0_n483 ) , .A( u0_u0_n484 ) , .ZN( u0_u0_n488 ) , .C2( u0_u0_n838 ) , .C1( u0_u0_n865 ) );
  AOI222_X1 u0_u0_U86 (.A2( u0_u0_n444 ) , .ZN( u0_u0_n475 ) , .B1( u0_u0_n837 ) , .A1( u0_u0_n844 ) , .C1( u0_u0_n847 ) , .C2( u0_u0_n856 ) , .B2( u0_u0_n869 ) );
  NOR4_X1 u0_u0_U87 (.A1( u0_u0_n472 ) , .ZN( u0_u0_n473 ) , .A4( u0_u0_n548 ) , .A2( u0_u0_n560 ) , .A3( u0_u0_n620 ) );
  AOI221_X1 u0_u0_U88 (.ZN( u0_u0_n474 ) , .C2( u0_u0_n719 ) , .B2( u0_u0_n836 ) , .C1( u0_u0_n850 ) , .B1( u0_u0_n864 ) , .A( u0_u0_n868 ) );
  NAND4_X1 u0_u0_U89 (.A4( u0_u0_n724 ) , .A3( u0_u0_n725 ) , .A2( u0_u0_n726 ) , .ZN( u0_u0_n746 ) , .A1( u0_u0_n861 ) );
  CLKBUF_X1 u0_u0_U9 (.Z( u0_u0_n439 ) , .A( u0_u0_n850 ) );
  INV_X1 u0_u0_U90 (.A( u0_u0_n714 ) , .ZN( u0_u0_n861 ) );
  NOR4_X1 u0_u0_U91 (.A4( u0_u0_n720 ) , .A3( u0_u0_n721 ) , .A2( u0_u0_n722 ) , .A1( u0_u0_n723 ) , .ZN( u0_u0_n724 ) );
  AOI221_X1 u0_u0_U92 (.B2( u0_u0_n439 ) , .A( u0_u0_n715 ) , .ZN( u0_u0_n726 ) , .C2( u0_u0_n849 ) , .C1( u0_u0_n865 ) , .B1( u0_u0_n866 ) );
  NAND4_X1 u0_u0_U93 (.A4( u0_u0_n579 ) , .A3( u0_u0_n580 ) , .A1( u0_u0_n581 ) , .ZN( u0_u0_n728 ) , .A2( u0_u0_n878 ) );
  AOI221_X1 u0_u0_U94 (.A( u0_u0_n570 ) , .C2( u0_u0_n571 ) , .ZN( u0_u0_n580 ) , .B2( u0_u0_n850 ) , .B1( u0_u0_n857 ) , .C1( u0_u0_n858 ) );
  NOR4_X1 u0_u0_U95 (.A4( u0_u0_n575 ) , .A3( u0_u0_n576 ) , .A2( u0_u0_n577 ) , .A1( u0_u0_n578 ) , .ZN( u0_u0_n579 ) );
  INV_X1 u0_u0_U96 (.A( u0_u0_n613 ) , .ZN( u0_u0_n878 ) );
  NOR4_X1 u0_u0_U97 (.A4( u0_u0_n615 ) , .A3( u0_u0_n616 ) , .A2( u0_u0_n617 ) , .A1( u0_u0_n618 ) , .ZN( u0_u0_n625 ) );
  NOR4_X1 u0_u0_U98 (.ZN( u0_u0_n626 ) , .A1( u0_u0_n662 ) , .A3( u0_u0_n672 ) , .A4( u0_u0_n688 ) , .A2( u0_u0_n771 ) );
  NOR2_X1 u0_u0_U99 (.ZN( u0_u0_n692 ) , .A1( u0_u0_n836 ) , .A2( u0_u0_n837 ) );
endmodule

