module des_des ( clk, decrypt, desIn, key1, key2, key3, desOut );
  input clk;
  input decrypt;
  input [63:0] desIn;
  input [55:0] key1;
  input [55:0] key2;
  input [55:0] key3;
  output [63:0] desOut;

  wire u0_FP_33, u0_FP_34, u0_FP_36, u0_FP_37, u0_FP_39, u0_FP_41, u0_FP_42, u0_FP_43, 
       u0_FP_44, u0_FP_45, u0_FP_46, u0_FP_48, u0_FP_49, u0_FP_50, u0_FP_51, u0_FP_52, u0_FP_53, 
       u0_FP_55, u0_FP_56, u0_FP_57, u0_FP_58, u0_FP_59, u0_FP_60, u0_FP_63, u0_FP_64, u0_K10_1, 
       u0_K10_14, u0_K10_17, u0_K10_18, u0_K10_19, u0_K10_20, u0_K10_32, u0_K11_37, u0_K11_42, u0_K11_48, 
       u0_K12_19, u0_K12_25, u0_K12_35, u0_K12_36, u0_K12_48, u0_K12_5, u0_K12_7, u0_K12_8, u0_K13_41, 
       u0_K14_23, u0_K14_24, u0_K14_25, u0_K14_26, u0_K14_29, u0_K14_5, u0_K14_7, u0_K15_13, u0_K16_18, 
       u0_K16_19, u0_K16_24, u0_K16_26, u0_K16_36, u0_K16_38, u0_K16_5, u0_K16_8, u0_K1_13, u0_K1_14, 
       u0_K1_17, u0_K1_30, u0_K1_31, u0_K2_11, u0_K2_12, u0_K2_18, u0_K2_20, u0_K2_29, u0_K2_30, 
       u0_K2_31, u0_K2_5, u0_K3_12, u0_K3_13, u0_K3_14, u0_K3_17, u0_K3_18, u0_K3_19, u0_K3_23, 
       u0_K3_5, u0_K3_6, u0_K4_36, u0_K4_43, u0_K4_48, u0_K4_6, u0_K5_1, u0_K5_18, u0_K5_24, 
       u0_K5_26, u0_K5_29, u0_K5_31, u0_K5_47, u0_K5_8, u0_K6_11, u0_K6_13, u0_K6_19, u0_K6_20, 
       u0_K6_23, u0_K6_24, u0_K6_41, u0_K8_11, u0_K8_13, u0_K8_19, u0_K9_12, u0_K9_13, u0_K9_14, 
       u0_K9_30, u0_K9_32, u0_K9_44, u0_K9_6, u0_R0_1, u0_R0_13, u0_R0_15, u0_R0_18, u0_R0_19, 
       u0_R0_20, u0_R0_21, u0_R0_28, u0_R0_32, u0_R0_4, u0_R0_7, u0_R0_8, u0_R0_9, u0_R10_1, 
       u0_R10_12, u0_R10_14, u0_R10_16, u0_R10_17, u0_R10_18, u0_R10_19, u0_R10_2, u0_R10_20, u0_R10_21, 
       u0_R10_24, u0_R10_25, u0_R10_28, u0_R10_29, u0_R10_3, u0_R10_4, u0_R10_5, u0_R11_10, u0_R11_11, 
       u0_R11_12, u0_R11_13, u0_R11_14, u0_R11_15, u0_R11_16, u0_R11_2, u0_R11_20, u0_R11_28, u0_R11_3, 
       u0_R11_32, u0_R11_5, u0_R11_6, u0_R12_16, u0_R12_17, u0_R12_19, u0_R12_20, u0_R12_22, u0_R12_23, 
       u0_R12_24, u0_R12_30, u0_R12_4, u0_R13_17, u0_R13_18, u0_R13_19, u0_R13_20, u0_R13_21, u0_R13_22, 
       u0_R13_23, u0_R13_24, u0_R13_25, u0_R13_26, u0_R13_27, u0_R13_28, u0_R13_29, u0_R13_30, u0_R13_31, 
       u0_R13_8, u0_R1_1, u0_R1_12, u0_R1_13, u0_R1_14, u0_R1_15, u0_R1_16, u0_R1_19, u0_R1_20, 
       u0_R1_21, u0_R1_22, u0_R1_24, u0_R1_25, u0_R1_26, u0_R1_27, u0_R1_28, u0_R1_29, u0_R1_3, 
       u0_R1_30, u0_R1_32, u0_R1_4, u0_R1_5, u0_R1_8, u0_R1_9, u0_R2_1, u0_R2_10, u0_R2_11, 
       u0_R2_12, u0_R2_13, u0_R2_14, u0_R2_16, u0_R2_2, u0_R2_21, u0_R2_22, u0_R2_25, u0_R2_28, 
       u0_R2_3, u0_R2_32, u0_R2_4, u0_R2_5, u0_R2_6, u0_R2_7, u0_R2_8, u0_R2_9, u0_R3_13, 
       u0_R3_15, u0_R3_17, u0_R3_18, u0_R3_20, u0_R3_22, u0_R3_24, u0_R3_25, u0_R3_32, u0_R3_5, 
       u0_R4_1, u0_R4_12, u0_R4_13, u0_R4_16, u0_R4_17, u0_R4_19, u0_R4_20, u0_R4_21, u0_R4_22, 
       u0_R4_24, u0_R4_25, u0_R4_26, u0_R4_27, u0_R4_28, u0_R4_29, u0_R4_3, u0_R4_30, u0_R4_32, 
       u0_R4_4, u0_R4_5, u0_R4_8, u0_R4_9, u0_R5_12, u0_R5_13, u0_R5_2, u0_R5_25, u0_R5_3, 
       u0_R5_32, u0_R5_4, u0_R5_5, u0_R5_7, u0_R5_8, u0_R5_9, u0_R6_10, u0_R6_11, u0_R6_12, 
       u0_R6_13, u0_R6_14, u0_R6_17, u0_R6_24, u0_R6_26, u0_R6_28, u0_R6_29, u0_R6_4, u0_R6_5, 
       u0_R6_7, u0_R6_8, u0_R6_9, u0_R7_1, u0_R7_12, u0_R7_14, u0_R7_17, u0_R7_20, u0_R7_21, 
       u0_R7_22, u0_R7_23, u0_R7_24, u0_R7_25, u0_R7_28, u0_R7_29, u0_R7_32, u0_R7_4, u0_R7_5, 
       u0_R7_8, u0_R7_9, u0_R8_1, u0_R8_12, u0_R8_13, u0_R8_17, u0_R8_19, u0_R8_20, u0_R8_21, 
       u0_R8_22, u0_R8_27, u0_R8_29, u0_R8_30, u0_R8_32, u0_R8_5, u0_R8_6, u0_R8_9, u0_R9_1, 
       u0_R9_10, u0_R9_11, u0_R9_12, u0_R9_13, u0_R9_16, u0_R9_17, u0_R9_18, u0_R9_19, u0_R9_2, 
       u0_R9_20, u0_R9_21, u0_R9_22, u0_R9_24, u0_R9_25, u0_R9_26, u0_R9_27, u0_R9_29, u0_R9_3, 
       u0_R9_30, u0_R9_31, u0_R9_32, u0_R9_4, u0_R9_5, u0_R9_6, u0_R9_7, u0_R9_8, u0_R9_9, 
       u0_desIn_r_1, u0_desIn_r_11, u0_desIn_r_15, u0_desIn_r_17, u0_desIn_r_23, u0_desIn_r_25, u0_desIn_r_27, u0_desIn_r_29, u0_desIn_r_3, 
       u0_desIn_r_31, u0_desIn_r_35, u0_desIn_r_37, u0_desIn_r_39, u0_desIn_r_47, u0_desIn_r_5, u0_desIn_r_51, u0_desIn_r_55, u0_desIn_r_57, 
       u0_desIn_r_59, u0_desIn_r_63, u0_desIn_r_7, u0_desIn_r_9, u0_key_r_0, u0_key_r_11, u0_key_r_12, u0_key_r_13, u0_key_r_14, 
       u0_key_r_16, u0_key_r_19, u0_key_r_2, u0_key_r_20, u0_key_r_21, u0_key_r_22, u0_key_r_23, u0_key_r_28, u0_key_r_29, 
       u0_key_r_30, u0_key_r_35, u0_key_r_4, u0_key_r_41, u0_key_r_42, u0_key_r_47, u0_key_r_48, u0_key_r_5, u0_key_r_50, 
       u0_key_r_54, u0_key_r_55, u0_key_r_6, u0_key_r_9, u0_out0_1, u0_out0_10, u0_out0_11, u0_out0_12, u0_out0_13, 
       u0_out0_14, u0_out0_15, u0_out0_16, u0_out0_17, u0_out0_18, u0_out0_19, u0_out0_2, u0_out0_20, u0_out0_21, 
       u0_out0_22, u0_out0_23, u0_out0_24, u0_out0_25, u0_out0_26, u0_out0_27, u0_out0_28, u0_out0_29, u0_out0_3, 
       u0_out0_30, u0_out0_31, u0_out0_32, u0_out0_4, u0_out0_5, u0_out0_6, u0_out0_7, u0_out0_8, u0_out0_9, 
       u0_out10_1, u0_out10_10, u0_out10_11, u0_out10_12, u0_out10_13, u0_out10_14, u0_out10_15, u0_out10_16, u0_out10_17, 
       u0_out10_18, u0_out10_19, u0_out10_2, u0_out10_20, u0_out10_21, u0_out10_22, u0_out10_23, u0_out10_24, u0_out10_25, 
       u0_out10_26, u0_out10_27, u0_out10_28, u0_out10_29, u0_out10_3, u0_out10_30, u0_out10_31, u0_out10_32, u0_out10_4, 
       u0_out10_5, u0_out10_6, u0_out10_7, u0_out10_8, u0_out10_9, u0_out11_1, u0_out11_10, u0_out11_11, u0_out11_12, 
       u0_out11_13, u0_out11_14, u0_out11_15, u0_out11_16, u0_out11_17, u0_out11_18, u0_out11_19, u0_out11_2, u0_out11_20, 
       u0_out11_21, u0_out11_22, u0_out11_23, u0_out11_24, u0_out11_25, u0_out11_26, u0_out11_27, u0_out11_28, u0_out11_29, 
       u0_out11_3, u0_out11_30, u0_out11_31, u0_out11_32, u0_out11_4, u0_out11_5, u0_out11_6, u0_out11_7, u0_out11_8, 
       u0_out11_9, u0_out12_1, u0_out12_10, u0_out12_11, u0_out12_12, u0_out12_13, u0_out12_14, u0_out12_15, u0_out12_16, 
       u0_out12_17, u0_out12_18, u0_out12_19, u0_out12_2, u0_out12_20, u0_out12_21, u0_out12_22, u0_out12_23, u0_out12_24, 
       u0_out12_25, u0_out12_26, u0_out12_27, u0_out12_28, u0_out12_29, u0_out12_3, u0_out12_30, u0_out12_31, u0_out12_32, 
       u0_out12_4, u0_out12_5, u0_out12_6, u0_out12_7, u0_out12_8, u0_out12_9, u0_out13_1, u0_out13_10, u0_out13_11, 
       u0_out13_12, u0_out13_13, u0_out13_14, u0_out13_15, u0_out13_17, u0_out13_18, u0_out13_19, u0_out13_2, u0_out13_20, 
       u0_out13_21, u0_out13_22, u0_out13_23, u0_out13_25, u0_out13_26, u0_out13_27, u0_out13_28, u0_out13_29, u0_out13_3, 
       u0_out13_31, u0_out13_32, u0_out13_4, u0_out13_5, u0_out13_7, u0_out13_8, u0_out13_9, u0_out14_1, u0_out14_10, 
       u0_out14_11, u0_out14_12, u0_out14_13, u0_out14_14, u0_out14_15, u0_out14_16, u0_out14_18, u0_out14_19, u0_out14_2, 
       u0_out14_20, u0_out14_21, u0_out14_22, u0_out14_24, u0_out14_25, u0_out14_26, u0_out14_27, u0_out14_28, u0_out14_29, 
       u0_out14_3, u0_out14_30, u0_out14_32, u0_out14_4, u0_out14_5, u0_out14_6, u0_out14_7, u0_out14_8, u0_out15_1, 
       u0_out15_10, u0_out15_11, u0_out15_12, u0_out15_13, u0_out15_14, u0_out15_15, u0_out15_16, u0_out15_17, u0_out15_18, 
       u0_out15_19, u0_out15_2, u0_out15_20, u0_out15_21, u0_out15_22, u0_out15_23, u0_out15_24, u0_out15_25, u0_out15_26, 
       u0_out15_27, u0_out15_28, u0_out15_29, u0_out15_3, u0_out15_30, u0_out15_31, u0_out15_32, u0_out15_4, u0_out15_5, 
       u0_out15_6, u0_out15_7, u0_out15_8, u0_out15_9, u0_out1_1, u0_out1_10, u0_out1_11, u0_out1_12, u0_out1_13, 
       u0_out1_14, u0_out1_16, u0_out1_17, u0_out1_18, u0_out1_19, u0_out1_2, u0_out1_20, u0_out1_22, u0_out1_23, 
       u0_out1_24, u0_out1_25, u0_out1_26, u0_out1_28, u0_out1_29, u0_out1_3, u0_out1_30, u0_out1_31, u0_out1_32, 
       u0_out1_4, u0_out1_6, u0_out1_7, u0_out1_8, u0_out1_9, u0_out2_1, u0_out2_10, u0_out2_11, u0_out2_12, 
       u0_out2_13, u0_out2_14, u0_out2_15, u0_out2_16, u0_out2_17, u0_out2_18, u0_out2_19, u0_out2_2, u0_out2_20, 
       u0_out2_21, u0_out2_22, u0_out2_23, u0_out2_24, u0_out2_25, u0_out2_26, u0_out2_27, u0_out2_28, u0_out2_29, 
       u0_out2_3, u0_out2_30, u0_out2_31, u0_out2_32, u0_out2_4, u0_out2_5, u0_out2_6, u0_out2_7, u0_out2_8, 
       u0_out2_9, u0_out3_1, u0_out3_10, u0_out3_11, u0_out3_12, u0_out3_13, u0_out3_14, u0_out3_15, u0_out3_16, 
       u0_out3_17, u0_out3_18, u0_out3_19, u0_out3_2, u0_out3_20, u0_out3_21, u0_out3_22, u0_out3_23, u0_out3_24, 
       u0_out3_25, u0_out3_26, u0_out3_27, u0_out3_28, u0_out3_29, u0_out3_3, u0_out3_30, u0_out3_31, u0_out3_32, 
       u0_out3_4, u0_out3_5, u0_out3_6, u0_out3_7, u0_out3_8, u0_out3_9, u0_out4_1, u0_out4_10, u0_out4_11, 
       u0_out4_13, u0_out4_14, u0_out4_15, u0_out4_16, u0_out4_17, u0_out4_18, u0_out4_19, u0_out4_2, u0_out4_20, 
       u0_out4_21, u0_out4_23, u0_out4_24, u0_out4_25, u0_out4_26, u0_out4_27, u0_out4_28, u0_out4_29, u0_out4_3, 
       u0_out4_30, u0_out4_31, u0_out4_4, u0_out4_5, u0_out4_6, u0_out4_8, u0_out4_9, u0_out5_1, u0_out5_10, 
       u0_out5_11, u0_out5_12, u0_out5_13, u0_out5_14, u0_out5_15, u0_out5_16, u0_out5_17, u0_out5_18, u0_out5_19, 
       u0_out5_2, u0_out5_20, u0_out5_21, u0_out5_22, u0_out5_23, u0_out5_24, u0_out5_25, u0_out5_26, u0_out5_27, 
       u0_out5_28, u0_out5_29, u0_out5_3, u0_out5_30, u0_out5_31, u0_out5_32, u0_out5_4, u0_out5_5, u0_out5_6, 
       u0_out5_7, u0_out5_8, u0_out5_9, u0_out6_1, u0_out6_10, u0_out6_11, u0_out6_13, u0_out6_16, u0_out6_17, 
       u0_out6_18, u0_out6_19, u0_out6_2, u0_out6_20, u0_out6_23, u0_out6_24, u0_out6_26, u0_out6_28, u0_out6_29, 
       u0_out6_30, u0_out6_31, u0_out6_4, u0_out6_6, u0_out6_9, u0_out7_1, u0_out7_10, u0_out7_11, u0_out7_12, 
       u0_out7_13, u0_out7_14, u0_out7_15, u0_out7_16, u0_out7_17, u0_out7_18, u0_out7_19, u0_out7_2, u0_out7_20, 
       u0_out7_21, u0_out7_22, u0_out7_23, u0_out7_24, u0_out7_25, u0_out7_26, u0_out7_27, u0_out7_28, u0_out7_29, 
       u0_out7_3, u0_out7_30, u0_out7_31, u0_out7_32, u0_out7_4, u0_out7_5, u0_out7_6, u0_out7_7, u0_out7_8, 
       u0_out7_9, u0_out8_1, u0_out8_10, u0_out8_11, u0_out8_12, u0_out8_13, u0_out8_14, u0_out8_15, u0_out8_16, 
       u0_out8_17, u0_out8_18, u0_out8_19, u0_out8_2, u0_out8_20, u0_out8_21, u0_out8_22, u0_out8_23, u0_out8_24, 
       u0_out8_25, u0_out8_26, u0_out8_27, u0_out8_28, u0_out8_29, u0_out8_3, u0_out8_30, u0_out8_31, u0_out8_32, 
       u0_out8_4, u0_out8_5, u0_out8_6, u0_out8_7, u0_out8_8, u0_out8_9, u0_out9_1, u0_out9_10, u0_out9_11, 
       u0_out9_12, u0_out9_13, u0_out9_14, u0_out9_15, u0_out9_16, u0_out9_17, u0_out9_18, u0_out9_19, u0_out9_2, 
       u0_out9_20, u0_out9_21, u0_out9_22, u0_out9_23, u0_out9_24, u0_out9_25, u0_out9_26, u0_out9_27, u0_out9_28, 
       u0_out9_29, u0_out9_3, u0_out9_30, u0_out9_31, u0_out9_32, u0_out9_4, u0_out9_5, u0_out9_6, u0_out9_7, 
       u0_out9_8, u0_out9_9, u0_u0_X_15, u0_u0_X_16, u0_u0_X_21, u0_u0_X_22, u0_u0_X_23, u0_u0_X_25, u0_u0_X_28, 
       u0_u0_X_33, u0_u0_X_42, u0_u0_X_44, u0_u0_X_45, u0_u0_X_46, u0_u10_X_21, u0_u10_X_22, u0_u10_X_34, u0_u10_X_41, 
       u0_u10_X_43, u0_u11_X_1, u0_u11_X_10, u0_u11_X_11, u0_u11_X_12, u0_u11_X_13, u0_u11_X_14, u0_u11_X_15, u0_u11_X_16, 
       u0_u11_X_18, u0_u11_X_20, u0_u11_X_22, u0_u11_X_33, u0_u11_X_34, u0_u11_X_39, u0_u11_X_40, u0_u11_X_45, u0_u11_X_46, 
       u0_u11_X_47, u0_u11_X_9, u0_u12_X_10, u0_u12_X_11, u0_u12_X_12, u0_u12_X_13, u0_u12_X_14, u0_u12_X_2, u0_u12_X_24, 
       u0_u12_X_26, u0_u12_X_27, u0_u12_X_28, u0_u12_X_30, u0_u12_X_32, u0_u12_X_33, u0_u12_X_34, u0_u12_X_35, u0_u12_X_36, 
       u0_u12_X_37, u0_u12_X_38, u0_u12_X_39, u0_u12_X_40, u0_u12_X_42, u0_u12_X_44, u0_u12_X_45, u0_u12_X_46, u0_u12_X_48, 
       u0_u12_X_5, u0_u12_X_7, u0_u13_X_1, u0_u13_X_10, u0_u13_X_11, u0_u13_X_12, u0_u13_X_19, u0_u13_X_2, u0_u13_X_20, 
       u0_u13_X_21, u0_u13_X_22, u0_u13_X_27, u0_u13_X_3, u0_u13_X_30, u0_u13_X_32, u0_u13_X_36, u0_u13_X_38, u0_u13_X_39, 
       u0_u13_X_4, u0_u13_X_40, u0_u13_X_41, u0_u13_X_42, u0_u13_X_43, u0_u13_X_44, u0_u13_X_46, u0_u13_X_47, u0_u13_X_48, 
       u0_u13_X_6, u0_u13_X_8, u0_u13_X_9, u0_u14_X_10, u0_u14_X_12, u0_u14_X_14, u0_u14_X_15, u0_u14_X_16, u0_u14_X_17, 
       u0_u14_X_18, u0_u14_X_19, u0_u14_X_20, u0_u14_X_21, u0_u14_X_22, u0_u14_X_23, u0_u14_X_24, u0_u14_X_25, u0_u14_X_47, 
       u0_u14_X_48, u0_u14_X_7, u0_u14_X_8, u0_u14_X_9, u0_u15_X_11, u0_u15_X_13, u0_u15_X_22, u0_u15_X_33, u0_u15_X_4, 
       u0_u15_X_42, u0_u15_X_44, u0_u15_X_45, u0_u15_X_9, u0_u1_X_15, u0_u1_X_16, u0_u1_X_17, u0_u1_X_19, u0_u1_X_21, 
       u0_u1_X_23, u0_u1_X_24, u0_u1_X_25, u0_u1_X_26, u0_u1_X_3, u0_u1_X_33, u0_u1_X_34, u0_u1_X_35, u0_u1_X_36, 
       u0_u1_X_37, u0_u1_X_38, u0_u1_X_39, u0_u1_X_4, u0_u1_X_40, u0_u1_X_42, u0_u1_X_6, u0_u1_X_8, u0_u1_X_9, 
       u0_u2_X_10, u0_u2_X_15, u0_u2_X_16, u0_u2_X_24, u0_u2_X_26, u0_u2_X_27, u0_u2_X_3, u0_u2_X_34, u0_u2_X_46, 
       u0_u2_X_9, u0_u3_X_22, u0_u3_X_24, u0_u3_X_26, u0_u3_X_27, u0_u3_X_28, u0_u3_X_29, u0_u3_X_31, u0_u3_X_34, 
       u0_u3_X_35, u0_u3_X_37, u0_u3_X_39, u0_u3_X_40, u0_u3_X_42, u0_u3_X_44, u0_u3_X_45, u0_u3_X_46, u0_u4_X_10, 
       u0_u4_X_11, u0_u4_X_12, u0_u4_X_13, u0_u4_X_14, u0_u4_X_15, u0_u4_X_16, u0_u4_X_17, u0_u4_X_19, u0_u4_X_2, 
       u0_u4_X_21, u0_u4_X_23, u0_u4_X_25, u0_u4_X_28, u0_u4_X_3, u0_u4_X_30, u0_u4_X_32, u0_u4_X_34, u0_u4_X_4, 
       u0_u4_X_43, u0_u4_X_44, u0_u4_X_45, u0_u4_X_46, u0_u4_X_48, u0_u4_X_5, u0_u4_X_7, u0_u4_X_9, u0_u5_X_10, 
       u0_u5_X_15, u0_u5_X_16, u0_u5_X_21, u0_u5_X_22, u0_u5_X_27, u0_u5_X_3, u0_u5_X_34, u0_u5_X_46, u0_u5_X_9, 
       u0_u6_X_15, u0_u6_X_16, u0_u6_X_2, u0_u6_X_21, u0_u6_X_22, u0_u6_X_23, u0_u6_X_24, u0_u6_X_31, u0_u6_X_32, 
       u0_u6_X_33, u0_u6_X_34, u0_u6_X_35, u0_u6_X_9, u0_u7_X_1, u0_u7_X_2, u0_u7_X_22, u0_u7_X_23, u0_u7_X_25, 
       u0_u7_X_27, u0_u7_X_28, u0_u7_X_29, u0_u7_X_3, u0_u7_X_30, u0_u7_X_31, u0_u7_X_32, u0_u7_X_33, u0_u7_X_34, 
       u0_u7_X_36, u0_u7_X_38, u0_u7_X_4, u0_u7_X_40, u0_u7_X_45, u0_u7_X_46, u0_u7_X_47, u0_u7_X_48, u0_u7_X_9, 
       u0_u8_X_10, u0_u8_X_15, u0_u8_X_16, u0_u8_X_18, u0_u8_X_20, u0_u8_X_22, u0_u8_X_23, u0_u8_X_25, u0_u8_X_27, 
       u0_u8_X_28, u0_u8_X_3, u0_u8_X_39, u0_u8_X_4, u0_u8_X_40, u0_u8_X_45, u0_u8_X_46, u0_u8_X_9, u0_u9_X_10, 
       u0_u9_X_11, u0_u9_X_13, u0_u9_X_15, u0_u9_X_16, u0_u9_X_21, u0_u9_X_22, u0_u9_X_23, u0_u9_X_25, u0_u9_X_27, 
       u0_u9_X_3, u0_u9_X_34, u0_u9_X_35, u0_u9_X_36, u0_u9_X_37, u0_u9_X_38, u0_u9_X_39, u0_u9_X_4, u0_u9_X_41, 
       u0_u9_X_43, u0_u9_X_46, u0_u9_X_5, u0_u9_X_7, u0_uk_K_r0_15, u0_uk_K_r0_28, u0_uk_K_r0_36, u0_uk_K_r0_49, u0_uk_K_r0_7, 
       u0_uk_K_r10_10, u0_uk_K_r10_18, u0_uk_K_r10_23, u0_uk_K_r10_27, u0_uk_K_r10_28, u0_uk_K_r10_32, u0_uk_K_r10_37, u0_uk_K_r10_41, u0_uk_K_r10_42, 
       u0_uk_K_r10_44, u0_uk_K_r10_9, u0_uk_K_r11_19, u0_uk_K_r11_20, u0_uk_K_r11_24, u0_uk_K_r11_25, u0_uk_K_r11_27, u0_uk_K_r11_29, u0_uk_K_r11_33, 
       u0_uk_K_r11_39, u0_uk_K_r11_4, u0_uk_K_r12_16, u0_uk_K_r13_0, u0_uk_K_r13_25, u0_uk_K_r13_38, u0_uk_K_r13_44, u0_uk_K_r14_10, u0_uk_K_r14_11, 
       u0_uk_K_r14_12, u0_uk_K_r14_15, u0_uk_K_r14_16, u0_uk_K_r14_18, u0_uk_K_r14_2, u0_uk_K_r14_45, u0_uk_K_r14_50, u0_uk_K_r14_8, u0_uk_K_r14_9, 
       u0_uk_K_r1_15, u0_uk_K_r1_16, u0_uk_K_r1_21, u0_uk_K_r1_44, u0_uk_K_r1_7, u0_uk_K_r2_13, u0_uk_K_r2_18, u0_uk_K_r2_20, u0_uk_K_r2_25, 
       u0_uk_K_r2_26, u0_uk_K_r2_27, u0_uk_K_r2_28, u0_uk_K_r2_33, u0_uk_K_r2_4, u0_uk_K_r2_41, u0_uk_K_r2_46, u0_uk_K_r2_50, u0_uk_K_r2_53, 
       u0_uk_K_r2_55, u0_uk_K_r3_10, u0_uk_K_r3_14, u0_uk_K_r4_0, u0_uk_K_r4_23, u0_uk_K_r4_33, u0_uk_K_r4_35, u0_uk_K_r4_38, u0_uk_K_r4_41, 
       u0_uk_K_r4_47, u0_uk_K_r5_10, u0_uk_K_r5_17, u0_uk_K_r5_39, u0_uk_K_r5_4, u0_uk_K_r6_0, u0_uk_K_r6_22, u0_uk_K_r6_26, u0_uk_K_r6_31, 
       u0_uk_K_r6_34, u0_uk_K_r6_46, u0_uk_K_r7_26, u0_uk_K_r8_16, u0_uk_K_r8_40, u0_uk_K_r8_41, u0_uk_K_r9_0, u0_uk_K_r9_1, u0_uk_K_r9_19, 
       u0_uk_K_r9_22, u0_uk_K_r9_25, u0_uk_K_r9_27, u0_uk_K_r9_30, u0_uk_K_r9_33, u0_uk_K_r9_35, u0_uk_K_r9_45, u0_uk_K_r9_6, u0_uk_K_r9_7, 
       u0_uk_K_r9_9, u0_uk_n10, u0_uk_n100, u0_uk_n1000, u0_uk_n1001, u0_uk_n1002, u0_uk_n1004, u0_uk_n1005, u0_uk_n1006, 
       u0_uk_n101, u0_uk_n1012, u0_uk_n102, u0_uk_n1024, u0_uk_n106, u0_uk_n107, u0_uk_n108, u0_uk_n109, u0_uk_n11, 
       u0_uk_n110, u0_uk_n113, u0_uk_n115, u0_uk_n116, u0_uk_n117, u0_uk_n118, u0_uk_n12, u0_uk_n121, u0_uk_n122, 
       u0_uk_n123, u0_uk_n126, u0_uk_n127, u0_uk_n128, u0_uk_n129, u0_uk_n13, u0_uk_n131, u0_uk_n139, u0_uk_n141, 
       u0_uk_n142, u0_uk_n143, u0_uk_n144, u0_uk_n145, u0_uk_n146, u0_uk_n147, u0_uk_n148, u0_uk_n151, u0_uk_n153, 
       u0_uk_n155, u0_uk_n156, u0_uk_n161, u0_uk_n162, u0_uk_n163, u0_uk_n164, u0_uk_n167, u0_uk_n168, u0_uk_n17, 
       u0_uk_n171, u0_uk_n172, u0_uk_n173, u0_uk_n174, u0_uk_n177, u0_uk_n178, u0_uk_n179, u0_uk_n18, u0_uk_n180, 
       u0_uk_n181, u0_uk_n182, u0_uk_n183, u0_uk_n184, u0_uk_n185, u0_uk_n187, u0_uk_n188, u0_uk_n189, u0_uk_n190, 
       u0_uk_n191, u0_uk_n192, u0_uk_n193, u0_uk_n195, u0_uk_n196, u0_uk_n197, u0_uk_n198, u0_uk_n199, u0_uk_n200, 
       u0_uk_n201, u0_uk_n202, u0_uk_n203, u0_uk_n204, u0_uk_n205, u0_uk_n206, u0_uk_n207, u0_uk_n208, u0_uk_n209, 
       u0_uk_n21, u0_uk_n210, u0_uk_n211, u0_uk_n212, u0_uk_n213, u0_uk_n214, u0_uk_n215, u0_uk_n216, u0_uk_n217, 
       u0_uk_n218, u0_uk_n219, u0_uk_n22, u0_uk_n220, u0_uk_n221, u0_uk_n222, u0_uk_n223, u0_uk_n224, u0_uk_n225, 
       u0_uk_n23, u0_uk_n230, u0_uk_n231, u0_uk_n232, u0_uk_n233, u0_uk_n238, u0_uk_n239, u0_uk_n240, u0_uk_n241, 
       u0_uk_n242, u0_uk_n243, u0_uk_n244, u0_uk_n248, u0_uk_n249, u0_uk_n250, u0_uk_n251, u0_uk_n252, u0_uk_n253, 
       u0_uk_n257, u0_uk_n259, u0_uk_n260, u0_uk_n261, u0_uk_n264, u0_uk_n266, u0_uk_n267, u0_uk_n269, u0_uk_n27, 
       u0_uk_n272, u0_uk_n275, u0_uk_n276, u0_uk_n278, u0_uk_n28, u0_uk_n282, u0_uk_n283, u0_uk_n285, u0_uk_n289, 
       u0_uk_n290, u0_uk_n293, u0_uk_n3, u0_uk_n300, u0_uk_n307, u0_uk_n31, u0_uk_n310, u0_uk_n314, u0_uk_n316, 
       u0_uk_n318, u0_uk_n32, u0_uk_n320, u0_uk_n324, u0_uk_n329, u0_uk_n33, u0_uk_n330, u0_uk_n331, u0_uk_n332, 
       u0_uk_n336, u0_uk_n337, u0_uk_n339, u0_uk_n341, u0_uk_n344, u0_uk_n347, u0_uk_n348, u0_uk_n352, u0_uk_n355, 
       u0_uk_n358, u0_uk_n361, u0_uk_n370, u0_uk_n371, u0_uk_n383, u0_uk_n384, u0_uk_n39, u0_uk_n392, u0_uk_n393, 
       u0_uk_n396, u0_uk_n4, u0_uk_n40, u0_uk_n400, u0_uk_n401, u0_uk_n405, u0_uk_n41, u0_uk_n410, u0_uk_n411, 
       u0_uk_n412, u0_uk_n413, u0_uk_n414, u0_uk_n418, u0_uk_n419, u0_uk_n420, u0_uk_n423, u0_uk_n424, u0_uk_n425, 
       u0_uk_n426, u0_uk_n428, u0_uk_n429, u0_uk_n430, u0_uk_n432, u0_uk_n433, u0_uk_n434, u0_uk_n436, u0_uk_n438, 
       u0_uk_n439, u0_uk_n440, u0_uk_n442, u0_uk_n445, u0_uk_n446, u0_uk_n447, u0_uk_n448, u0_uk_n45, u0_uk_n450, 
       u0_uk_n457, u0_uk_n471, u0_uk_n497, u0_uk_n499, u0_uk_n5, u0_uk_n502, u0_uk_n505, u0_uk_n508, u0_uk_n510, 
       u0_uk_n511, u0_uk_n513, u0_uk_n517, u0_uk_n519, u0_uk_n522, u0_uk_n523, u0_uk_n525, u0_uk_n529, u0_uk_n530, 
       u0_uk_n531, u0_uk_n532, u0_uk_n534, u0_uk_n535, u0_uk_n536, u0_uk_n539, u0_uk_n542, u0_uk_n544, u0_uk_n545, 
       u0_uk_n546, u0_uk_n547, u0_uk_n549, u0_uk_n55, u0_uk_n550, u0_uk_n552, u0_uk_n553, u0_uk_n554, u0_uk_n555, 
       u0_uk_n557, u0_uk_n558, u0_uk_n560, u0_uk_n561, u0_uk_n562, u0_uk_n565, u0_uk_n566, u0_uk_n567, u0_uk_n568, 
       u0_uk_n570, u0_uk_n573, u0_uk_n574, u0_uk_n575, u0_uk_n577, u0_uk_n578, u0_uk_n579, u0_uk_n58, u0_uk_n580, 
       u0_uk_n581, u0_uk_n583, u0_uk_n598, u0_uk_n60, u0_uk_n604, u0_uk_n61, u0_uk_n615, u0_uk_n627, u0_uk_n629, 
       u0_uk_n63, u0_uk_n632, u0_uk_n635, u0_uk_n636, u0_uk_n637, u0_uk_n639, u0_uk_n640, u0_uk_n642, u0_uk_n643, 
       u0_uk_n644, u0_uk_n645, u0_uk_n649, u0_uk_n650, u0_uk_n651, u0_uk_n652, u0_uk_n653, u0_uk_n654, u0_uk_n657, 
       u0_uk_n658, u0_uk_n659, u0_uk_n660, u0_uk_n661, u0_uk_n663, u0_uk_n666, u0_uk_n668, u0_uk_n669, u0_uk_n67, 
       u0_uk_n670, u0_uk_n674, u0_uk_n675, u0_uk_n684, u0_uk_n687, u0_uk_n690, u0_uk_n696, u0_uk_n697, u0_uk_n699, 
       u0_uk_n711, u0_uk_n719, u0_uk_n722, u0_uk_n723, u0_uk_n725, u0_uk_n726, u0_uk_n727, u0_uk_n729, u0_uk_n73, 
       u0_uk_n731, u0_uk_n734, u0_uk_n735, u0_uk_n741, u0_uk_n746, u0_uk_n748, u0_uk_n751, u0_uk_n759, u0_uk_n761, 
       u0_uk_n763, u0_uk_n768, u0_uk_n780, u0_uk_n783, u0_uk_n786, u0_uk_n793, u0_uk_n799, u0_uk_n8, u0_uk_n800, 
       u0_uk_n809, u0_uk_n810, u0_uk_n813, u0_uk_n815, u0_uk_n816, u0_uk_n83, u0_uk_n832, u0_uk_n839, u0_uk_n855, 
       u0_uk_n866, u0_uk_n868, u0_uk_n869, u0_uk_n875, u0_uk_n883, u0_uk_n892, u0_uk_n898, u0_uk_n9, u0_uk_n904, 
       u0_uk_n91, u0_uk_n915, u0_uk_n916, u0_uk_n917, u0_uk_n918, u0_uk_n92, u0_uk_n93, u0_uk_n933, u0_uk_n934, 
       u0_uk_n94, u0_uk_n949, u0_uk_n950, u0_uk_n956, u0_uk_n96, u0_uk_n963, u0_uk_n976, u0_uk_n98, u0_uk_n982, 
       u0_uk_n985, u0_uk_n99, u0_uk_n990, u0_uk_n999, u1_FP_33, u1_FP_37, u1_FP_40, u1_FP_41, u1_FP_44, 
       u1_FP_45, u1_FP_52, u1_FP_53, u1_FP_55, u1_FP_56, u1_FP_60, u1_FP_61, u1_K10_1, u1_K10_11, 
       u1_K10_13, u1_K10_14, u1_K10_18, u1_K10_2, u1_K10_20, u1_K10_23, u1_K10_24, u1_K10_25, u1_K10_26, 
       u1_K10_29, u1_K10_30, u1_K10_31, u1_K10_32, u1_K10_36, u1_K10_41, u1_K10_42, u1_K10_43, u1_K10_44, 
       u1_K10_47, u1_K10_48, u1_K10_5, u1_K10_6, u1_K10_7, u1_K10_8, u1_K11_11, u1_K11_13, u1_K11_2, 
       u1_K11_23, u1_K11_25, u1_K11_29, u1_K11_32, u1_K11_35, u1_K11_37, u1_K11_38, u1_K11_48, u1_K11_7, 
       u1_K12_18, u1_K12_19, u1_K12_2, u1_K12_20, u1_K12_24, u1_K12_25, u1_K12_26, u1_K12_35, u1_K12_36, 
       u1_K12_37, u1_K12_38, u1_K12_41, u1_K12_43, u1_K12_47, u1_K12_48, u1_K12_6, u1_K12_8, u1_K13_14, 
       u1_K13_17, u1_K13_18, u1_K13_20, u1_K13_29, u1_K13_30, u1_K13_31, u1_K13_32, u1_K13_35, u1_K13_37, 
       u1_K13_48, u1_K13_8, u1_K14_1, u1_K14_2, u1_K14_29, u1_K14_30, u1_K14_31, u1_K14_32, u1_K14_42, 
       u1_K14_44, u1_K14_47, u1_K14_48, u1_K15_11, u1_K15_12, u1_K15_13, u1_K15_14, u1_K15_18, u1_K15_2, 
       u1_K15_20, u1_K15_23, u1_K15_24, u1_K15_25, u1_K15_29, u1_K15_31, u1_K15_32, u1_K15_35, u1_K15_36, 
       u1_K15_37, u1_K15_41, u1_K15_42, u1_K15_44, u1_K15_48, u1_K15_5, u1_K15_6, u1_K15_7, u1_K16_11, 
       u1_K16_12, u1_K16_13, u1_K16_14, u1_K16_17, u1_K16_18, u1_K16_19, u1_K16_2, u1_K16_20, u1_K16_30, 
       u1_K16_31, u1_K16_32, u1_K16_35, u1_K16_41, u1_K16_42, u1_K16_44, u1_K16_48, u1_K16_6, u1_K16_8, 
       u1_K1_1, u1_K1_17, u1_K1_19, u1_K1_43, u1_K1_47, u1_K1_6, u1_K1_8, u1_K2_1, u1_K2_11, 
       u1_K2_12, u1_K2_13, u1_K2_17, u1_K2_18, u1_K2_2, u1_K2_20, u1_K2_23, u1_K2_24, u1_K2_25, 
       u1_K2_26, u1_K2_29, u1_K2_30, u1_K2_31, u1_K2_42, u1_K2_43, u1_K2_44, u1_K2_47, u1_K2_48, 
       u1_K2_5, u1_K2_6, u1_K2_8, u1_K3_1, u1_K3_12, u1_K3_14, u1_K3_17, u1_K3_18, u1_K3_19, 
       u1_K3_2, u1_K3_20, u1_K3_23, u1_K3_25, u1_K3_26, u1_K3_29, u1_K3_31, u1_K3_35, u1_K3_36, 
       u1_K3_37, u1_K3_38, u1_K3_41, u1_K3_42, u1_K3_43, u1_K3_44, u1_K3_47, u1_K3_48, u1_K3_5, 
       u1_K3_6, u1_K3_7, u1_K3_8, u1_K4_1, u1_K4_11, u1_K4_12, u1_K4_13, u1_K4_14, u1_K4_17, 
       u1_K4_18, u1_K4_19, u1_K4_24, u1_K4_30, u1_K4_32, u1_K4_35, u1_K4_36, u1_K4_37, u1_K4_38, 
       u1_K4_41, u1_K4_42, u1_K4_43, u1_K4_44, u1_K4_47, u1_K4_48, u1_K4_6, u1_K5_1, u1_K5_11, 
       u1_K5_12, u1_K5_13, u1_K5_14, u1_K5_17, u1_K5_18, u1_K5_19, u1_K5_2, u1_K5_23, u1_K5_24, 
       u1_K5_25, u1_K5_26, u1_K5_29, u1_K5_30, u1_K5_31, u1_K5_32, u1_K5_37, u1_K5_38, u1_K5_41, 
       u1_K5_42, u1_K5_44, u1_K5_47, u1_K5_48, u1_K5_5, u1_K5_6, u1_K5_7, u1_K5_8, u1_K6_1, 
       u1_K6_11, u1_K6_12, u1_K6_13, u1_K6_14, u1_K6_20, u1_K6_23, u1_K6_24, u1_K6_25, u1_K6_26, 
       u1_K6_29, u1_K6_30, u1_K6_31, u1_K6_32, u1_K6_35, u1_K6_36, u1_K6_37, u1_K6_38, u1_K6_41, 
       u1_K6_42, u1_K6_43, u1_K6_44, u1_K6_47, u1_K6_48, u1_K6_5, u1_K6_6, u1_K6_7, u1_K6_8, 
       u1_K7_1, u1_K7_11, u1_K7_14, u1_K7_17, u1_K7_18, u1_K7_19, u1_K7_2, u1_K7_23, u1_K7_26, 
       u1_K7_29, u1_K7_30, u1_K7_31, u1_K7_35, u1_K7_37, u1_K7_38, u1_K7_41, u1_K7_43, u1_K7_44, 
       u1_K7_47, u1_K7_48, u1_K7_5, u1_K7_7, u1_K8_1, u1_K8_11, u1_K8_13, u1_K8_14, u1_K8_18, 
       u1_K8_2, u1_K8_20, u1_K8_23, u1_K8_24, u1_K8_25, u1_K8_26, u1_K8_30, u1_K8_31, u1_K8_32, 
       u1_K8_35, u1_K8_36, u1_K8_38, u1_K8_41, u1_K8_42, u1_K8_44, u1_K8_47, u1_K8_48, u1_K8_5, 
       u1_K8_7, u1_K9_12, u1_K9_13, u1_K9_14, u1_K9_17, u1_K9_23, u1_K9_24, u1_K9_25, u1_K9_29, 
       u1_K9_31, u1_K9_36, u1_K9_37, u1_K9_38, u1_K9_43, u1_K9_44, u1_K9_47, u1_K9_5, u1_K9_6, 
       u1_K9_7, u1_K9_8, u1_R0_1, u1_R0_12, u1_R0_13, u1_R0_16, u1_R0_17, u1_R0_20, u1_R0_21, 
       u1_R0_28, u1_R0_29, u1_R0_32, u1_R0_4, u1_R0_5, u1_R0_7, u1_R0_8, u1_R0_9, u1_R10_1, 
       u1_R10_10, u1_R10_12, u1_R10_13, u1_R10_14, u1_R10_16, u1_R10_17, u1_R10_24, u1_R10_25, u1_R10_28, 
       u1_R10_29, u1_R10_32, u1_R10_5, u1_R11_1, u1_R11_10, u1_R11_12, u1_R11_13, u1_R11_20, u1_R11_21, 
       u1_R11_24, u1_R11_4, u1_R11_5, u1_R11_8, u1_R11_9, u1_R12_1, u1_R12_20, u1_R12_21, u1_R12_23, 
       u1_R12_29, u1_R12_32, u1_R13_1, u1_R13_13, u1_R13_16, u1_R13_17, u1_R13_20, u1_R13_21, u1_R13_24, 
       u1_R13_25, u1_R13_28, u1_R13_29, u1_R13_4, u1_R13_5, u1_R13_8, u1_R13_9, u1_R1_1, u1_R1_12, 
       u1_R1_13, u1_R1_16, u1_R1_17, u1_R1_20, u1_R1_24, u1_R1_25, u1_R1_28, u1_R1_29, u1_R1_32, 
       u1_R1_4, u1_R1_5, u1_R1_9, u1_R2_1, u1_R2_12, u1_R2_13, u1_R2_16, u1_R2_17, u1_R2_2, 
       u1_R2_20, u1_R2_21, u1_R2_24, u1_R2_25, u1_R2_28, u1_R2_29, u1_R2_32, u1_R2_5, u1_R2_7, 
       u1_R2_8, u1_R2_9, u1_R3_1, u1_R3_12, u1_R3_13, u1_R3_15, u1_R3_16, u1_R3_17, u1_R3_18, 
       u1_R3_20, u1_R3_21, u1_R3_24, u1_R3_25, u1_R3_28, u1_R3_29, u1_R3_32, u1_R3_4, u1_R3_5, 
       u1_R3_8, u1_R3_9, u1_R4_1, u1_R4_13, u1_R4_14, u1_R4_16, u1_R4_17, u1_R4_20, u1_R4_21, 
       u1_R4_24, u1_R4_25, u1_R4_28, u1_R4_29, u1_R4_3, u1_R4_32, u1_R4_4, u1_R4_5, u1_R4_6, 
       u1_R4_7, u1_R4_8, u1_R4_9, u1_R5_1, u1_R5_12, u1_R5_13, u1_R5_16, u1_R5_17, u1_R5_18, 
       u1_R5_20, u1_R5_21, u1_R5_23, u1_R5_24, u1_R5_25, u1_R5_28, u1_R5_29, u1_R5_31, u1_R5_32, 
       u1_R5_4, u1_R5_5, u1_R5_8, u1_R5_9, u1_R6_1, u1_R6_10, u1_R6_13, u1_R6_16, u1_R6_17, 
       u1_R6_2, u1_R6_20, u1_R6_21, u1_R6_24, u1_R6_25, u1_R6_28, u1_R6_29, u1_R6_32, u1_R6_4, 
       u1_R6_8, u1_R6_9, u1_R7_1, u1_R7_12, u1_R7_13, u1_R7_15, u1_R7_16, u1_R7_17, u1_R7_18, 
       u1_R7_20, u1_R7_24, u1_R7_25, u1_R7_28, u1_R7_29, u1_R7_32, u1_R7_4, u1_R7_5, u1_R7_6, 
       u1_R7_7, u1_R7_8, u1_R7_9, u1_R8_1, u1_R8_13, u1_R8_15, u1_R8_16, u1_R8_17, u1_R8_20, 
       u1_R8_21, u1_R8_22, u1_R8_24, u1_R8_25, u1_R8_28, u1_R8_29, u1_R8_32, u1_R8_4, u1_R8_5, 
       u1_R8_6, u1_R8_8, u1_R8_9, u1_R9_1, u1_R9_12, u1_R9_15, u1_R9_16, u1_R9_20, u1_R9_21, 
       u1_R9_23, u1_R9_24, u1_R9_25, u1_R9_4, u1_R9_8, u1_R9_9, u1_desIn_r_25, u1_desIn_r_29, u1_desIn_r_37, 
       u1_desIn_r_39, u1_desIn_r_57, u1_out0_1, u1_out0_10, u1_out0_11, u1_out0_12, u1_out0_13, u1_out0_14, u1_out0_15, 
       u1_out0_16, u1_out0_17, u1_out0_18, u1_out0_19, u1_out0_2, u1_out0_20, u1_out0_21, u1_out0_22, u1_out0_23, 
       u1_out0_24, u1_out0_25, u1_out0_26, u1_out0_27, u1_out0_28, u1_out0_29, u1_out0_3, u1_out0_30, u1_out0_31, 
       u1_out0_32, u1_out0_4, u1_out0_5, u1_out0_6, u1_out0_7, u1_out0_8, u1_out0_9, u1_out10_1, u1_out10_10, 
       u1_out10_11, u1_out10_12, u1_out10_13, u1_out10_14, u1_out10_15, u1_out10_16, u1_out10_17, u1_out10_18, u1_out10_19, 
       u1_out10_2, u1_out10_20, u1_out10_21, u1_out10_22, u1_out10_23, u1_out10_24, u1_out10_25, u1_out10_26, u1_out10_27, 
       u1_out10_28, u1_out10_29, u1_out10_3, u1_out10_30, u1_out10_31, u1_out10_32, u1_out10_4, u1_out10_5, u1_out10_6, 
       u1_out10_7, u1_out10_8, u1_out10_9, u1_out11_1, u1_out11_10, u1_out11_11, u1_out11_12, u1_out11_13, u1_out11_14, 
       u1_out11_15, u1_out11_16, u1_out11_17, u1_out11_18, u1_out11_19, u1_out11_2, u1_out11_20, u1_out11_21, u1_out11_22, 
       u1_out11_23, u1_out11_24, u1_out11_25, u1_out11_26, u1_out11_27, u1_out11_28, u1_out11_29, u1_out11_3, u1_out11_30, 
       u1_out11_31, u1_out11_32, u1_out11_4, u1_out11_5, u1_out11_6, u1_out11_7, u1_out11_8, u1_out11_9, u1_out12_1, 
       u1_out12_10, u1_out12_11, u1_out12_12, u1_out12_13, u1_out12_14, u1_out12_15, u1_out12_16, u1_out12_17, u1_out12_18, 
       u1_out12_19, u1_out12_2, u1_out12_20, u1_out12_21, u1_out12_22, u1_out12_23, u1_out12_24, u1_out12_25, u1_out12_26, 
       u1_out12_27, u1_out12_28, u1_out12_29, u1_out12_3, u1_out12_30, u1_out12_31, u1_out12_32, u1_out12_4, u1_out12_5, 
       u1_out12_6, u1_out12_7, u1_out12_8, u1_out12_9, u1_out13_1, u1_out13_10, u1_out13_11, u1_out13_12, u1_out13_13, 
       u1_out13_14, u1_out13_15, u1_out13_16, u1_out13_17, u1_out13_18, u1_out13_19, u1_out13_2, u1_out13_20, u1_out13_21, 
       u1_out13_22, u1_out13_23, u1_out13_24, u1_out13_25, u1_out13_26, u1_out13_27, u1_out13_28, u1_out13_29, u1_out13_3, 
       u1_out13_30, u1_out13_31, u1_out13_32, u1_out13_4, u1_out13_5, u1_out13_6, u1_out13_7, u1_out13_8, u1_out13_9, 
       u1_out14_1, u1_out14_10, u1_out14_11, u1_out14_12, u1_out14_13, u1_out14_14, u1_out14_15, u1_out14_16, u1_out14_17, 
       u1_out14_18, u1_out14_19, u1_out14_2, u1_out14_20, u1_out14_21, u1_out14_22, u1_out14_23, u1_out14_24, u1_out14_25, 
       u1_out14_26, u1_out14_27, u1_out14_28, u1_out14_29, u1_out14_3, u1_out14_30, u1_out14_31, u1_out14_32, u1_out14_4, 
       u1_out14_5, u1_out14_6, u1_out14_7, u1_out14_8, u1_out14_9, u1_out15_1, u1_out15_10, u1_out15_11, u1_out15_12, 
       u1_out15_13, u1_out15_14, u1_out15_15, u1_out15_16, u1_out15_17, u1_out15_18, u1_out15_19, u1_out15_2, u1_out15_20, 
       u1_out15_21, u1_out15_22, u1_out15_23, u1_out15_24, u1_out15_25, u1_out15_26, u1_out15_27, u1_out15_28, u1_out15_29, 
       u1_out15_3, u1_out15_30, u1_out15_31, u1_out15_32, u1_out15_4, u1_out15_5, u1_out15_6, u1_out15_7, u1_out15_8, 
       u1_out15_9, u1_out1_1, u1_out1_10, u1_out1_11, u1_out1_12, u1_out1_13, u1_out1_14, u1_out1_15, u1_out1_16, 
       u1_out1_17, u1_out1_18, u1_out1_19, u1_out1_2, u1_out1_20, u1_out1_21, u1_out1_22, u1_out1_23, u1_out1_24, 
       u1_out1_25, u1_out1_26, u1_out1_27, u1_out1_28, u1_out1_29, u1_out1_3, u1_out1_30, u1_out1_31, u1_out1_32, 
       u1_out1_4, u1_out1_5, u1_out1_6, u1_out1_7, u1_out1_8, u1_out1_9, u1_out2_1, u1_out2_10, u1_out2_11, 
       u1_out2_12, u1_out2_13, u1_out2_14, u1_out2_15, u1_out2_16, u1_out2_17, u1_out2_18, u1_out2_19, u1_out2_2, 
       u1_out2_20, u1_out2_21, u1_out2_22, u1_out2_23, u1_out2_24, u1_out2_25, u1_out2_26, u1_out2_27, u1_out2_28, 
       u1_out2_29, u1_out2_3, u1_out2_30, u1_out2_31, u1_out2_32, u1_out2_4, u1_out2_5, u1_out2_6, u1_out2_7, 
       u1_out2_8, u1_out2_9, u1_out3_1, u1_out3_10, u1_out3_11, u1_out3_12, u1_out3_13, u1_out3_14, u1_out3_15, 
       u1_out3_16, u1_out3_17, u1_out3_18, u1_out3_19, u1_out3_2, u1_out3_20, u1_out3_21, u1_out3_22, u1_out3_23, 
       u1_out3_24, u1_out3_25, u1_out3_26, u1_out3_27, u1_out3_28, u1_out3_29, u1_out3_3, u1_out3_30, u1_out3_31, 
       u1_out3_32, u1_out3_4, u1_out3_5, u1_out3_6, u1_out3_7, u1_out3_8, u1_out3_9, u1_out4_1, u1_out4_10, 
       u1_out4_11, u1_out4_12, u1_out4_13, u1_out4_14, u1_out4_15, u1_out4_16, u1_out4_17, u1_out4_18, u1_out4_19, 
       u1_out4_2, u1_out4_20, u1_out4_21, u1_out4_22, u1_out4_23, u1_out4_24, u1_out4_25, u1_out4_26, u1_out4_27, 
       u1_out4_28, u1_out4_29, u1_out4_3, u1_out4_30, u1_out4_31, u1_out4_32, u1_out4_4, u1_out4_5, u1_out4_6, 
       u1_out4_7, u1_out4_8, u1_out4_9, u1_out5_1, u1_out5_10, u1_out5_11, u1_out5_12, u1_out5_13, u1_out5_14, 
       u1_out5_15, u1_out5_16, u1_out5_17, u1_out5_18, u1_out5_19, u1_out5_2, u1_out5_20, u1_out5_21, u1_out5_22, 
       u1_out5_23, u1_out5_24, u1_out5_25, u1_out5_26, u1_out5_27, u1_out5_28, u1_out5_29, u1_out5_3, u1_out5_30, 
       u1_out5_31, u1_out5_32, u1_out5_4, u1_out5_5, u1_out5_6, u1_out5_7, u1_out5_8, u1_out5_9, u1_out6_1, 
       u1_out6_10, u1_out6_11, u1_out6_12, u1_out6_13, u1_out6_14, u1_out6_15, u1_out6_16, u1_out6_17, u1_out6_18, 
       u1_out6_19, u1_out6_2, u1_out6_20, u1_out6_21, u1_out6_22, u1_out6_23, u1_out6_24, u1_out6_25, u1_out6_26, 
       u1_out6_27, u1_out6_28, u1_out6_29, u1_out6_3, u1_out6_30, u1_out6_31, u1_out6_32, u1_out6_4, u1_out6_5, 
       u1_out6_6, u1_out6_7, u1_out6_8, u1_out6_9, u1_out7_1, u1_out7_10, u1_out7_11, u1_out7_12, u1_out7_13, 
       u1_out7_14, u1_out7_15, u1_out7_16, u1_out7_17, u1_out7_18, u1_out7_19, u1_out7_2, u1_out7_20, u1_out7_21, 
       u1_out7_22, u1_out7_23, u1_out7_24, u1_out7_25, u1_out7_26, u1_out7_27, u1_out7_28, u1_out7_29, u1_out7_3, 
       u1_out7_30, u1_out7_31, u1_out7_32, u1_out7_4, u1_out7_5, u1_out7_6, u1_out7_7, u1_out7_8, u1_out7_9, 
       u1_out8_1, u1_out8_10, u1_out8_11, u1_out8_12, u1_out8_13, u1_out8_14, u1_out8_15, u1_out8_16, u1_out8_17, 
       u1_out8_18, u1_out8_19, u1_out8_2, u1_out8_20, u1_out8_21, u1_out8_22, u1_out8_23, u1_out8_24, u1_out8_25, 
       u1_out8_26, u1_out8_27, u1_out8_28, u1_out8_29, u1_out8_3, u1_out8_30, u1_out8_31, u1_out8_32, u1_out8_4, 
       u1_out8_5, u1_out8_6, u1_out8_7, u1_out8_8, u1_out8_9, u1_out9_1, u1_out9_10, u1_out9_11, u1_out9_12, 
       u1_out9_13, u1_out9_14, u1_out9_15, u1_out9_16, u1_out9_17, u1_out9_18, u1_out9_19, u1_out9_2, u1_out9_20, 
       u1_out9_21, u1_out9_22, u1_out9_23, u1_out9_24, u1_out9_25, u1_out9_26, u1_out9_27, u1_out9_28, u1_out9_29, 
       u1_out9_3, u1_out9_30, u1_out9_31, u1_out9_32, u1_out9_4, u1_out9_5, u1_out9_6, u1_out9_7, u1_out9_8, 
       u1_out9_9, u1_u0_X_10, u1_u0_X_11, u1_u0_X_12, u1_u0_X_13, u1_u0_X_14, u1_u0_X_15, u1_u0_X_16, u1_u0_X_2, 
       u1_u0_X_21, u1_u0_X_22, u1_u0_X_23, u1_u0_X_24, u1_u0_X_25, u1_u0_X_26, u1_u0_X_27, u1_u0_X_28, u1_u0_X_29, 
       u1_u0_X_3, u1_u0_X_30, u1_u0_X_31, u1_u0_X_32, u1_u0_X_33, u1_u0_X_34, u1_u0_X_35, u1_u0_X_36, u1_u0_X_37, 
       u1_u0_X_38, u1_u0_X_39, u1_u0_X_4, u1_u0_X_40, u1_u0_X_42, u1_u0_X_44, u1_u0_X_45, u1_u0_X_46, u1_u0_X_48, 
       u1_u0_X_5, u1_u0_X_7, u1_u0_X_9, u1_u10_X_1, u1_u10_X_10, u1_u10_X_15, u1_u10_X_16, u1_u10_X_18, u1_u10_X_20, 
       u1_u10_X_21, u1_u10_X_24, u1_u10_X_26, u1_u10_X_27, u1_u10_X_28, u1_u10_X_3, u1_u10_X_33, u1_u10_X_39, u1_u10_X_4, 
       u1_u10_X_40, u1_u10_X_41, u1_u10_X_42, u1_u10_X_43, u1_u10_X_44, u1_u10_X_45, u1_u10_X_46, u1_u10_X_47, u1_u10_X_6, 
       u1_u10_X_8, u1_u10_X_9, u1_u11_X_10, u1_u11_X_11, u1_u11_X_12, u1_u11_X_13, u1_u11_X_14, u1_u11_X_16, u1_u11_X_22, 
       u1_u11_X_27, u1_u11_X_28, u1_u11_X_29, u1_u11_X_3, u1_u11_X_30, u1_u11_X_31, u1_u11_X_32, u1_u11_X_33, u1_u11_X_34, 
       u1_u11_X_39, u1_u11_X_4, u1_u11_X_40, u1_u11_X_45, u1_u11_X_46, u1_u11_X_5, u1_u11_X_7, u1_u11_X_9, u1_u12_X_1, 
       u1_u12_X_10, u1_u12_X_16, u1_u12_X_21, u1_u12_X_22, u1_u12_X_23, u1_u12_X_24, u1_u12_X_25, u1_u12_X_26, u1_u12_X_27, 
       u1_u12_X_28, u1_u12_X_3, u1_u12_X_33, u1_u12_X_34, u1_u12_X_36, u1_u12_X_38, u1_u12_X_39, u1_u12_X_4, u1_u12_X_40, 
       u1_u12_X_41, u1_u12_X_42, u1_u12_X_43, u1_u12_X_44, u1_u12_X_45, u1_u12_X_46, u1_u12_X_47, u1_u12_X_9, u1_u13_X_10, 
       u1_u13_X_11, u1_u13_X_12, u1_u13_X_13, u1_u13_X_14, u1_u13_X_15, u1_u13_X_16, u1_u13_X_17, u1_u13_X_18, u1_u13_X_19, 
       u1_u13_X_20, u1_u13_X_21, u1_u13_X_22, u1_u13_X_23, u1_u13_X_24, u1_u13_X_25, u1_u13_X_26, u1_u13_X_27, u1_u13_X_28, 
       u1_u13_X_3, u1_u13_X_33, u1_u13_X_35, u1_u13_X_36, u1_u13_X_37, u1_u13_X_38, u1_u13_X_39, u1_u13_X_4, u1_u13_X_40, 
       u1_u13_X_41, u1_u13_X_43, u1_u13_X_45, u1_u13_X_46, u1_u13_X_5, u1_u13_X_6, u1_u13_X_7, u1_u13_X_8, u1_u13_X_9, 
       u1_u14_X_1, u1_u14_X_10, u1_u14_X_15, u1_u14_X_16, u1_u14_X_17, u1_u14_X_19, u1_u14_X_21, u1_u14_X_22, u1_u14_X_27, 
       u1_u14_X_28, u1_u14_X_3, u1_u14_X_33, u1_u14_X_34, u1_u14_X_39, u1_u14_X_4, u1_u14_X_40, u1_u14_X_45, u1_u14_X_46, 
       u1_u14_X_47, u1_u14_X_9, u1_u15_X_1, u1_u15_X_10, u1_u15_X_15, u1_u15_X_16, u1_u15_X_21, u1_u15_X_22, u1_u15_X_23, 
       u1_u15_X_24, u1_u15_X_25, u1_u15_X_26, u1_u15_X_27, u1_u15_X_28, u1_u15_X_3, u1_u15_X_33, u1_u15_X_36, u1_u15_X_38, 
       u1_u15_X_39, u1_u15_X_4, u1_u15_X_40, u1_u15_X_45, u1_u15_X_46, u1_u15_X_47, u1_u15_X_5, u1_u15_X_7, u1_u15_X_9, 
       u1_u1_X_15, u1_u1_X_16, u1_u1_X_21, u1_u1_X_22, u1_u1_X_27, u1_u1_X_28, u1_u1_X_3, u1_u1_X_33, u1_u1_X_34, 
       u1_u1_X_35, u1_u1_X_36, u1_u1_X_37, u1_u1_X_38, u1_u1_X_39, u1_u1_X_4, u1_u1_X_40, u1_u1_X_45, u1_u1_X_46, 
       u1_u1_X_9, u1_u2_X_10, u1_u2_X_11, u1_u2_X_13, u1_u2_X_15, u1_u2_X_16, u1_u2_X_21, u1_u2_X_22, u1_u2_X_27, 
       u1_u2_X_28, u1_u2_X_3, u1_u2_X_30, u1_u2_X_32, u1_u2_X_33, u1_u2_X_34, u1_u2_X_39, u1_u2_X_4, u1_u2_X_40, 
       u1_u2_X_45, u1_u2_X_46, u1_u2_X_9, u1_u3_X_15, u1_u3_X_16, u1_u3_X_21, u1_u3_X_22, u1_u3_X_27, u1_u3_X_28, 
       u1_u3_X_33, u1_u3_X_34, u1_u3_X_39, u1_u3_X_4, u1_u3_X_40, u1_u3_X_45, u1_u3_X_46, u1_u3_X_5, u1_u3_X_7, 
       u1_u3_X_9, u1_u4_X_10, u1_u4_X_15, u1_u4_X_16, u1_u4_X_21, u1_u4_X_28, u1_u4_X_3, u1_u4_X_33, u1_u4_X_34, 
       u1_u4_X_39, u1_u4_X_4, u1_u4_X_40, u1_u4_X_45, u1_u4_X_46, u1_u4_X_9, u1_u5_X_15, u1_u5_X_16, u1_u5_X_17, 
       u1_u5_X_19, u1_u5_X_22, u1_u5_X_27, u1_u5_X_28, u1_u5_X_3, u1_u5_X_33, u1_u5_X_34, u1_u5_X_39, u1_u5_X_40, 
       u1_u5_X_45, u1_u5_X_46, u1_u6_X_10, u1_u6_X_15, u1_u6_X_16, u1_u6_X_21, u1_u6_X_22, u1_u6_X_28, u1_u6_X_3, 
       u1_u6_X_33, u1_u6_X_39, u1_u6_X_4, u1_u6_X_40, u1_u6_X_45, u1_u6_X_9, u1_u7_X_10, u1_u7_X_16, u1_u7_X_17, 
       u1_u7_X_19, u1_u7_X_21, u1_u7_X_22, u1_u7_X_27, u1_u7_X_28, u1_u7_X_33, u1_u7_X_34, u1_u7_X_39, u1_u7_X_4, 
       u1_u7_X_40, u1_u7_X_45, u1_u7_X_46, u1_u7_X_6, u1_u7_X_8, u1_u7_X_9, u1_u8_X_15, u1_u8_X_16, u1_u8_X_21, 
       u1_u8_X_28, u1_u8_X_3, u1_u8_X_30, u1_u8_X_32, u1_u8_X_33, u1_u8_X_34, u1_u8_X_39, u1_u8_X_4, u1_u8_X_40, 
       u1_u8_X_45, u1_u8_X_46, u1_u9_X_10, u1_u9_X_15, u1_u9_X_16, u1_u9_X_17, u1_u9_X_19, u1_u9_X_21, u1_u9_X_27, 
       u1_u9_X_28, u1_u9_X_3, u1_u9_X_34, u1_u9_X_39, u1_u9_X_4, u1_u9_X_40, u1_u9_X_45, u1_u9_X_46, u1_uk_n1002, 
       u1_uk_n1003, u1_uk_n1015, u1_uk_n1021, u1_uk_n1023, u1_uk_n1025, u1_uk_n1029, u1_uk_n1031, u1_uk_n1034, u1_uk_n1038, 
       u1_uk_n1050, u1_uk_n1054, u1_uk_n1056, u1_uk_n1057, u1_uk_n1058, u1_uk_n1060, u1_uk_n1061, u1_uk_n1063, u1_uk_n1065, 
       u1_uk_n1070, u1_uk_n1073, u1_uk_n1074, u1_uk_n1076, u1_uk_n1079, u1_uk_n1080, u1_uk_n1083, u1_uk_n1088, u1_uk_n1090, 
       u1_uk_n1092, u1_uk_n1096, u1_uk_n1101, u1_uk_n1104, u1_uk_n1105, u1_uk_n1106, u1_uk_n1109, u1_uk_n1113, u1_uk_n1114, 
       u1_uk_n1115, u1_uk_n1118, u1_uk_n1119, u1_uk_n1121, u1_uk_n1123, u1_uk_n1124, u1_uk_n1125, u1_uk_n1126, u1_uk_n1128, 
       u1_uk_n1130, u1_uk_n1134, u1_uk_n1138, u1_uk_n1140, u1_uk_n1143, u1_uk_n1147, u1_uk_n1148, u1_uk_n1153, u1_uk_n1154, 
       u1_uk_n1155, u1_uk_n1156, u1_uk_n1157, u1_uk_n1158, u1_uk_n1159, u1_uk_n1160, u1_uk_n1163, u1_uk_n1166, u1_uk_n1167, 
       u1_uk_n1170, u1_uk_n1171, u1_uk_n299, u1_uk_n312, u1_uk_n349, u1_uk_n353, u1_uk_n366, u1_uk_n369, u1_uk_n376, 
       u1_uk_n379, u1_uk_n382, u1_uk_n385, u1_uk_n386, u1_uk_n407, u1_uk_n421, u1_uk_n437, u1_uk_n443, u1_uk_n454, 
       u1_uk_n496, u1_uk_n504, u1_uk_n509, u1_uk_n515, u1_uk_n520, u1_uk_n524, u1_uk_n605, u1_uk_n608, u1_uk_n672, 
       u1_uk_n676, u1_uk_n677, u1_uk_n678, u1_uk_n685, u1_uk_n702, u1_uk_n948, u1_uk_n949, u1_uk_n950, u1_uk_n955, 
       u1_uk_n969, u1_uk_n970, u1_uk_n973, u1_uk_n974, u1_uk_n976, u1_uk_n985, u1_uk_n988, u1_uk_n989, u1_uk_n993, 
       u2_FP_33, u2_FP_36, u2_FP_37, u2_FP_40, u2_FP_41, u2_FP_44, u2_FP_45, u2_FP_48, u2_FP_49, 
       u2_FP_52, u2_FP_53, u2_FP_55, u2_FP_56, u2_FP_57, u2_FP_60, u2_FP_61, u2_FP_64, u2_K10_1, 
       u2_K10_11, u2_K10_13, u2_K10_14, u2_K10_17, u2_K10_18, u2_K10_19, u2_K10_20, u2_K10_23, u2_K10_24, 
       u2_K10_25, u2_K10_26, u2_K10_36, u2_K10_42, u2_K10_43, u2_K10_44, u2_K10_48, u2_K10_5, u2_K10_7, 
       u2_K10_8, u2_K11_11, u2_K11_13, u2_K11_24, u2_K11_26, u2_K11_29, u2_K12_2, u2_K12_20, u2_K12_25, 
       u2_K12_36, u2_K12_38, u2_K12_47, u2_K12_48, u2_K13_32, u2_K13_35, u2_K13_37, u2_K13_48, u2_K14_38, 
       u2_K15_1, u2_K15_12, u2_K15_17, u2_K15_2, u2_K15_23, u2_K15_29, u2_K15_31, u2_K15_35, u2_K15_44, 
       u2_K16_1, u2_K16_11, u2_K16_12, u2_K16_13, u2_K16_14, u2_K16_17, u2_K16_18, u2_K16_19, u2_K16_2, 
       u2_K16_20, u2_K16_23, u2_K16_24, u2_K16_25, u2_K16_26, u2_K16_30, u2_K16_31, u2_K16_32, u2_K16_35, 
       u2_K16_36, u2_K16_38, u2_K16_41, u2_K16_42, u2_K16_44, u2_K16_47, u2_K16_48, u2_K16_5, u2_K16_6, 
       u2_K16_7, u2_K16_8, u2_K1_43, u2_K2_1, u2_K2_11, u2_K2_12, u2_K2_13, u2_K2_17, u2_K2_18, 
       u2_K2_2, u2_K2_20, u2_K2_23, u2_K2_24, u2_K2_25, u2_K2_26, u2_K2_29, u2_K2_30, u2_K2_31, 
       u2_K2_35, u2_K2_36, u2_K2_37, u2_K2_38, u2_K2_42, u2_K2_44, u2_K2_47, u2_K2_48, u2_K2_5, 
       u2_K2_6, u2_K2_8, u2_K3_13, u2_K3_19, u2_K3_20, u2_K3_23, u2_K3_26, u2_K3_42, u2_K3_43, 
       u2_K3_47, u2_K3_48, u2_K4_14, u2_K4_18, u2_K4_19, u2_K4_24, u2_K4_48, u2_K4_6, u2_K4_7, 
       u2_K5_11, u2_K5_13, u2_K5_14, u2_K5_17, u2_K5_18, u2_K5_19, u2_K5_2, u2_K5_23, u2_K5_24, 
       u2_K5_25, u2_K5_26, u2_K5_29, u2_K5_30, u2_K5_31, u2_K5_32, u2_K5_37, u2_K5_38, u2_K5_41, 
       u2_K5_44, u2_K5_48, u2_K5_5, u2_K5_6, u2_K5_8, u2_K6_1, u2_K6_11, u2_K6_13, u2_K6_14, 
       u2_K6_19, u2_K6_20, u2_K6_24, u2_K6_32, u2_K6_47, u2_K6_6, u2_K6_8, u2_K7_26, u2_K7_30, 
       u2_K7_31, u2_K7_35, u2_K7_37, u2_K7_38, u2_K7_43, u2_K7_48, u2_K7_5, u2_K7_7, u2_K8_1, 
       u2_K8_11, u2_K8_13, u2_K8_14, u2_K8_17, u2_K8_18, u2_K8_19, u2_K8_2, u2_K8_20, u2_K8_47, 
       u2_K8_48, u2_K8_5, u2_K8_6, u2_K8_7, u2_K8_8, u2_K9_12, u2_K9_14, u2_K9_23, u2_K9_25, 
       u2_K9_36, u2_K9_37, u2_K9_38, u2_K9_43, u2_K9_5, u2_R0_1, u2_R0_12, u2_R0_13, u2_R0_16, 
       u2_R0_17, u2_R0_19, u2_R0_20, u2_R0_21, u2_R0_24, u2_R0_25, u2_R0_29, u2_R0_32, u2_R0_4, 
       u2_R0_5, u2_R0_7, u2_R0_8, u2_R0_9, u2_R10_1, u2_R10_12, u2_R10_13, u2_R10_16, u2_R10_21, 
       u2_R10_25, u2_R10_29, u2_R10_3, u2_R10_32, u2_R10_4, u2_R10_7, u2_R10_8, u2_R10_9, u2_R11_1, 
       u2_R11_21, u2_R11_24, u2_R11_4, u2_R12_20, u2_R12_21, u2_R12_22, u2_R12_25, u2_R13_1, u2_R13_12, 
       u2_R13_16, u2_R13_17, u2_R13_20, u2_R13_22, u2_R13_24, u2_R13_25, u2_R13_27, u2_R13_29, u2_R13_32, 
       u2_R13_5, u2_R13_9, u2_R1_1, u2_R1_12, u2_R1_13, u2_R1_14, u2_R1_15, u2_R1_16, u2_R1_17, 
       u2_R1_2, u2_R1_25, u2_R1_27, u2_R1_28, u2_R1_29, u2_R1_3, u2_R1_30, u2_R1_31, u2_R1_32, 
       u2_R1_5, u2_R1_6, u2_R1_7, u2_R1_8, u2_R1_9, u2_R2_1, u2_R2_10, u2_R2_11, u2_R2_12, 
       u2_R2_13, u2_R2_16, u2_R2_17, u2_R2_19, u2_R2_2, u2_R2_20, u2_R2_21, u2_R2_25, u2_R2_3, 
       u2_R2_32, u2_R2_4, u2_R2_5, u2_R2_6, u2_R2_7, u2_R2_8, u2_R2_9, u2_R3_1, u2_R3_12, 
       u2_R3_13, u2_R3_16, u2_R3_17, u2_R3_18, u2_R3_20, u2_R3_21, u2_R3_22, u2_R3_24, u2_R3_25, 
       u2_R3_28, u2_R3_29, u2_R3_30, u2_R3_4, u2_R3_5, u2_R3_8, u2_R3_9, u2_R4_1, u2_R4_12, 
       u2_R4_13, u2_R4_14, u2_R4_17, u2_R4_21, u2_R4_22, u2_R4_24, u2_R4_28, u2_R4_29, u2_R4_31, 
       u2_R4_32, u2_R4_4, u2_R4_5, u2_R4_6, u2_R4_8, u2_R4_9, u2_R5_1, u2_R5_10, u2_R5_11, 
       u2_R5_12, u2_R5_13, u2_R5_14, u2_R5_16, u2_R5_17, u2_R5_20, u2_R5_21, u2_R5_23, u2_R5_24, 
       u2_R5_25, u2_R5_26, u2_R5_28, u2_R5_29, u2_R5_32, u2_R5_4, u2_R5_5, u2_R5_8, u2_R5_9, 
       u2_R6_1, u2_R6_12, u2_R6_13, u2_R6_2, u2_R6_28, u2_R6_32, u2_R6_4, u2_R6_5, u2_R6_8, 
       u2_R6_9, u2_R7_1, u2_R7_11, u2_R7_12, u2_R7_13, u2_R7_14, u2_R7_15, u2_R7_16, u2_R7_17, 
       u2_R7_22, u2_R7_24, u2_R7_25, u2_R7_28, u2_R7_29, u2_R7_3, u2_R7_4, u2_R7_5, u2_R7_6, 
       u2_R7_7, u2_R7_8, u2_R7_9, u2_R8_1, u2_R8_12, u2_R8_13, u2_R8_15, u2_R8_16, u2_R8_17, 
       u2_R8_20, u2_R8_22, u2_R8_24, u2_R8_25, u2_R8_26, u2_R8_27, u2_R8_28, u2_R8_29, u2_R8_32, 
       u2_R8_4, u2_R8_5, u2_R8_6, u2_R8_8, u2_R8_9, u2_R9_12, u2_R9_13, u2_R9_17, u2_R9_20, 
       u2_R9_32, u2_R9_8, u2_R9_9, u2_desIn_r_1, u2_desIn_r_25, u2_desIn_r_27, u2_desIn_r_33, u2_desIn_r_57, u2_key_r_14, 
       u2_key_r_23, u2_key_r_30, u2_key_r_7, u2_out0_11, u2_out0_12, u2_out0_13, u2_out0_14, u2_out0_15, u2_out0_18, 
       u2_out0_19, u2_out0_2, u2_out0_21, u2_out0_22, u2_out0_25, u2_out0_27, u2_out0_28, u2_out0_29, u2_out0_3, 
       u2_out0_32, u2_out0_4, u2_out0_5, u2_out0_7, u2_out0_8, u2_out10_1, u2_out10_10, u2_out10_11, u2_out10_12, 
       u2_out10_13, u2_out10_14, u2_out10_15, u2_out10_16, u2_out10_18, u2_out10_19, u2_out10_2, u2_out10_20, u2_out10_21, 
       u2_out10_22, u2_out10_24, u2_out10_25, u2_out10_26, u2_out10_27, u2_out10_28, u2_out10_29, u2_out10_3, u2_out10_30, 
       u2_out10_32, u2_out10_4, u2_out10_5, u2_out10_6, u2_out10_7, u2_out10_8, u2_out11_1, u2_out11_10, u2_out11_11, 
       u2_out11_12, u2_out11_13, u2_out11_14, u2_out11_15, u2_out11_16, u2_out11_17, u2_out11_18, u2_out11_19, u2_out11_2, 
       u2_out11_20, u2_out11_21, u2_out11_22, u2_out11_23, u2_out11_24, u2_out11_25, u2_out11_26, u2_out11_27, u2_out11_28, 
       u2_out11_29, u2_out11_3, u2_out11_30, u2_out11_31, u2_out11_32, u2_out11_4, u2_out11_5, u2_out11_6, u2_out11_7, 
       u2_out11_8, u2_out11_9, u2_out12_11, u2_out12_12, u2_out12_13, u2_out12_14, u2_out12_15, u2_out12_17, u2_out12_18, 
       u2_out12_19, u2_out12_2, u2_out12_21, u2_out12_22, u2_out12_23, u2_out12_25, u2_out12_27, u2_out12_28, u2_out12_29, 
       u2_out12_3, u2_out12_31, u2_out12_32, u2_out12_4, u2_out12_5, u2_out12_7, u2_out12_8, u2_out12_9, u2_out13_11, 
       u2_out13_12, u2_out13_14, u2_out13_15, u2_out13_19, u2_out13_21, u2_out13_22, u2_out13_25, u2_out13_27, u2_out13_29, 
       u2_out13_3, u2_out13_32, u2_out13_4, u2_out13_5, u2_out13_7, u2_out13_8, u2_out14_1, u2_out14_10, u2_out14_11, 
       u2_out14_12, u2_out14_13, u2_out14_14, u2_out14_15, u2_out14_16, u2_out14_17, u2_out14_18, u2_out14_19, u2_out14_2, 
       u2_out14_20, u2_out14_21, u2_out14_22, u2_out14_23, u2_out14_24, u2_out14_25, u2_out14_26, u2_out14_27, u2_out14_28, 
       u2_out14_29, u2_out14_3, u2_out14_30, u2_out14_31, u2_out14_32, u2_out14_4, u2_out14_5, u2_out14_6, u2_out14_7, 
       u2_out14_8, u2_out14_9, u2_out15_1, u2_out15_10, u2_out15_11, u2_out15_12, u2_out15_13, u2_out15_14, u2_out15_15, 
       u2_out15_16, u2_out15_17, u2_out15_18, u2_out15_19, u2_out15_2, u2_out15_20, u2_out15_21, u2_out15_22, u2_out15_23, 
       u2_out15_24, u2_out15_25, u2_out15_26, u2_out15_27, u2_out15_28, u2_out15_29, u2_out15_3, u2_out15_30, u2_out15_31, 
       u2_out15_32, u2_out15_4, u2_out15_5, u2_out15_6, u2_out15_7, u2_out15_8, u2_out15_9, u2_out1_1, u2_out1_10, 
       u2_out1_11, u2_out1_12, u2_out1_13, u2_out1_14, u2_out1_15, u2_out1_16, u2_out1_17, u2_out1_18, u2_out1_19, 
       u2_out1_2, u2_out1_20, u2_out1_21, u2_out1_22, u2_out1_23, u2_out1_24, u2_out1_25, u2_out1_26, u2_out1_27, 
       u2_out1_28, u2_out1_29, u2_out1_3, u2_out1_30, u2_out1_31, u2_out1_32, u2_out1_4, u2_out1_5, u2_out1_6, 
       u2_out1_7, u2_out1_8, u2_out1_9, u2_out2_1, u2_out2_10, u2_out2_11, u2_out2_12, u2_out2_13, u2_out2_14, 
       u2_out2_15, u2_out2_16, u2_out2_17, u2_out2_18, u2_out2_19, u2_out2_2, u2_out2_20, u2_out2_21, u2_out2_22, 
       u2_out2_23, u2_out2_24, u2_out2_25, u2_out2_26, u2_out2_27, u2_out2_28, u2_out2_29, u2_out2_3, u2_out2_30, 
       u2_out2_31, u2_out2_32, u2_out2_4, u2_out2_5, u2_out2_6, u2_out2_7, u2_out2_8, u2_out2_9, u2_out3_1, 
       u2_out3_10, u2_out3_11, u2_out3_13, u2_out3_14, u2_out3_15, u2_out3_16, u2_out3_17, u2_out3_18, u2_out3_19, 
       u2_out3_2, u2_out3_20, u2_out3_21, u2_out3_23, u2_out3_24, u2_out3_25, u2_out3_26, u2_out3_27, u2_out3_28, 
       u2_out3_29, u2_out3_3, u2_out3_30, u2_out3_31, u2_out3_4, u2_out3_5, u2_out3_6, u2_out3_8, u2_out3_9, 
       u2_out4_1, u2_out4_10, u2_out4_11, u2_out4_12, u2_out4_13, u2_out4_14, u2_out4_15, u2_out4_16, u2_out4_17, 
       u2_out4_18, u2_out4_19, u2_out4_2, u2_out4_20, u2_out4_21, u2_out4_22, u2_out4_23, u2_out4_24, u2_out4_25, 
       u2_out4_26, u2_out4_27, u2_out4_28, u2_out4_29, u2_out4_3, u2_out4_30, u2_out4_31, u2_out4_32, u2_out4_4, 
       u2_out4_5, u2_out4_6, u2_out4_7, u2_out4_8, u2_out4_9, u2_out5_1, u2_out5_10, u2_out5_11, u2_out5_12, 
       u2_out5_13, u2_out5_14, u2_out5_15, u2_out5_16, u2_out5_17, u2_out5_18, u2_out5_19, u2_out5_2, u2_out5_20, 
       u2_out5_21, u2_out5_22, u2_out5_23, u2_out5_24, u2_out5_25, u2_out5_26, u2_out5_27, u2_out5_28, u2_out5_29, 
       u2_out5_3, u2_out5_30, u2_out5_31, u2_out5_32, u2_out5_4, u2_out5_5, u2_out5_6, u2_out5_7, u2_out5_8, 
       u2_out5_9, u2_out6_1, u2_out6_10, u2_out6_11, u2_out6_12, u2_out6_13, u2_out6_14, u2_out6_15, u2_out6_16, 
       u2_out6_17, u2_out6_18, u2_out6_19, u2_out6_2, u2_out6_20, u2_out6_21, u2_out6_22, u2_out6_23, u2_out6_24, 
       u2_out6_25, u2_out6_26, u2_out6_27, u2_out6_28, u2_out6_29, u2_out6_3, u2_out6_30, u2_out6_31, u2_out6_32, 
       u2_out6_4, u2_out6_5, u2_out6_6, u2_out6_7, u2_out6_8, u2_out6_9, u2_out7_1, u2_out7_10, u2_out7_13, 
       u2_out7_15, u2_out7_16, u2_out7_17, u2_out7_18, u2_out7_2, u2_out7_20, u2_out7_21, u2_out7_23, u2_out7_24, 
       u2_out7_26, u2_out7_27, u2_out7_28, u2_out7_30, u2_out7_31, u2_out7_5, u2_out7_6, u2_out7_9, u2_out8_1, 
       u2_out8_10, u2_out8_11, u2_out8_12, u2_out8_13, u2_out8_14, u2_out8_15, u2_out8_16, u2_out8_17, u2_out8_18, 
       u2_out8_19, u2_out8_2, u2_out8_20, u2_out8_21, u2_out8_22, u2_out8_23, u2_out8_24, u2_out8_25, u2_out8_26, 
       u2_out8_27, u2_out8_28, u2_out8_29, u2_out8_3, u2_out8_30, u2_out8_31, u2_out8_32, u2_out8_4, u2_out8_5, 
       u2_out8_6, u2_out8_7, u2_out8_8, u2_out8_9, u2_out9_1, u2_out9_10, u2_out9_11, u2_out9_12, u2_out9_13, 
       u2_out9_14, u2_out9_15, u2_out9_16, u2_out9_17, u2_out9_18, u2_out9_19, u2_out9_2, u2_out9_20, u2_out9_21, 
       u2_out9_22, u2_out9_23, u2_out9_24, u2_out9_25, u2_out9_26, u2_out9_27, u2_out9_28, u2_out9_29, u2_out9_3, 
       u2_out9_30, u2_out9_31, u2_out9_32, u2_out9_4, u2_out9_5, u2_out9_6, u2_out9_7, u2_out9_8, u2_out9_9, 
       u2_u0_X_10, u2_u0_X_11, u2_u0_X_12, u2_u0_X_25, u2_u0_X_26, u2_u0_X_27, u2_u0_X_28, u2_u0_X_30, u2_u0_X_32, 
       u2_u0_X_33, u2_u0_X_34, u2_u0_X_35, u2_u0_X_37, u2_u0_X_39, u2_u0_X_40, u2_u0_X_45, u2_u0_X_46, u2_u0_X_48, 
       u2_u0_X_7, u2_u0_X_8, u2_u0_X_9, u2_u10_X_10, u2_u10_X_15, u2_u10_X_16, u2_u10_X_18, u2_u10_X_21, u2_u10_X_22, 
       u2_u10_X_23, u2_u10_X_25, u2_u10_X_27, u2_u10_X_28, u2_u10_X_30, u2_u10_X_32, u2_u10_X_33, u2_u10_X_34, u2_u10_X_35, 
       u2_u10_X_36, u2_u10_X_37, u2_u10_X_38, u2_u10_X_39, u2_u10_X_40, u2_u10_X_41, u2_u10_X_42, u2_u10_X_43, u2_u10_X_44, 
       u2_u10_X_45, u2_u10_X_46, u2_u10_X_48, u2_u10_X_7, u2_u10_X_8, u2_u10_X_9, u2_u11_X_15, u2_u11_X_16, u2_u11_X_21, 
       u2_u11_X_22, u2_u11_X_24, u2_u11_X_26, u2_u11_X_27, u2_u11_X_28, u2_u11_X_29, u2_u11_X_3, u2_u11_X_31, u2_u11_X_33, 
       u2_u11_X_34, u2_u11_X_35, u2_u11_X_37, u2_u11_X_39, u2_u11_X_40, u2_u11_X_41, u2_u11_X_43, u2_u11_X_45, u2_u11_X_46, 
       u2_u11_X_6, u2_u11_X_8, u2_u11_X_9, u2_u12_X_1, u2_u12_X_10, u2_u12_X_11, u2_u12_X_12, u2_u12_X_25, u2_u12_X_26, 
       u2_u12_X_27, u2_u12_X_28, u2_u12_X_29, u2_u12_X_3, u2_u12_X_31, u2_u12_X_33, u2_u12_X_34, u2_u12_X_36, u2_u12_X_38, 
       u2_u12_X_39, u2_u12_X_4, u2_u12_X_40, u2_u12_X_41, u2_u12_X_42, u2_u12_X_43, u2_u12_X_44, u2_u12_X_45, u2_u12_X_46, 
       u2_u12_X_47, u2_u12_X_6, u2_u12_X_8, u2_u12_X_9, u2_u13_X_25, u2_u13_X_26, u2_u13_X_27, u2_u13_X_28, u2_u13_X_34, 
       u2_u13_X_35, u2_u13_X_37, u2_u13_X_39, u2_u13_X_40, u2_u13_X_41, u2_u13_X_42, u2_u13_X_43, u2_u13_X_44, u2_u13_X_45, 
       u2_u13_X_46, u2_u13_X_47, u2_u13_X_48, u2_u14_X_10, u2_u14_X_11, u2_u14_X_13, u2_u14_X_15, u2_u14_X_16, u2_u14_X_18, 
       u2_u14_X_20, u2_u14_X_21, u2_u14_X_22, u2_u14_X_27, u2_u14_X_28, u2_u14_X_3, u2_u14_X_30, u2_u14_X_32, u2_u14_X_34, 
       u2_u14_X_39, u2_u14_X_4, u2_u14_X_41, u2_u14_X_43, u2_u14_X_45, u2_u14_X_46, u2_u14_X_5, u2_u14_X_7, u2_u14_X_9, 
       u2_u15_X_10, u2_u15_X_15, u2_u15_X_16, u2_u15_X_21, u2_u15_X_22, u2_u15_X_27, u2_u15_X_28, u2_u15_X_3, u2_u15_X_33, 
       u2_u15_X_39, u2_u15_X_4, u2_u15_X_40, u2_u15_X_45, u2_u15_X_46, u2_u15_X_9, u2_u1_X_15, u2_u1_X_16, u2_u1_X_21, 
       u2_u1_X_22, u2_u1_X_27, u2_u1_X_3, u2_u1_X_33, u2_u1_X_34, u2_u1_X_39, u2_u1_X_4, u2_u1_X_40, u2_u1_X_41, 
       u2_u1_X_43, u2_u1_X_45, u2_u1_X_46, u2_u1_X_9, u2_u2_X_15, u2_u2_X_16, u2_u2_X_27, u2_u2_X_28, u2_u2_X_29, 
       u2_u2_X_30, u2_u2_X_31, u2_u2_X_32, u2_u2_X_33, u2_u2_X_34, u2_u2_X_35, u2_u2_X_37, u2_u2_X_39, u2_u2_X_5, 
       u2_u2_X_7, u2_u3_X_21, u2_u3_X_22, u2_u3_X_27, u2_u3_X_33, u2_u3_X_34, u2_u3_X_35, u2_u3_X_43, u2_u3_X_44, 
       u2_u3_X_45, u2_u3_X_46, u2_u4_X_1, u2_u4_X_10, u2_u4_X_15, u2_u4_X_16, u2_u4_X_21, u2_u4_X_22, u2_u4_X_28, 
       u2_u4_X_3, u2_u4_X_34, u2_u4_X_39, u2_u4_X_4, u2_u4_X_40, u2_u4_X_46, u2_u4_X_47, u2_u4_X_9, u2_u5_X_10, 
       u2_u5_X_15, u2_u5_X_16, u2_u5_X_22, u2_u5_X_23, u2_u5_X_25, u2_u5_X_27, u2_u5_X_28, u2_u5_X_29, u2_u5_X_3, 
       u2_u5_X_31, u2_u5_X_34, u2_u5_X_36, u2_u5_X_38, u2_u5_X_39, u2_u5_X_4, u2_u5_X_40, u2_u5_X_45, u2_u6_X_10, 
       u2_u6_X_22, u2_u6_X_27, u2_u6_X_28, u2_u6_X_3, u2_u6_X_33, u2_u6_X_4, u2_u6_X_40, u2_u6_X_45, u2_u6_X_46, 
       u2_u6_X_9, u2_u7_X_10, u2_u7_X_15, u2_u7_X_16, u2_u7_X_21, u2_u7_X_22, u2_u7_X_23, u2_u7_X_24, u2_u7_X_4, 
       u2_u7_X_44, u2_u7_X_45, u2_u7_X_46, u2_u7_X_9, u2_u8_X_1, u2_u8_X_15, u2_u8_X_27, u2_u8_X_28, u2_u8_X_29, 
       u2_u8_X_3, u2_u8_X_30, u2_u8_X_31, u2_u8_X_32, u2_u8_X_34, u2_u8_X_39, u2_u8_X_40, u2_u8_X_45, u2_u8_X_46, 
       u2_u8_X_47, u2_u9_X_10, u2_u9_X_15, u2_u9_X_16, u2_u9_X_21, u2_u9_X_27, u2_u9_X_28, u2_u9_X_29, u2_u9_X_3, 
       u2_u9_X_30, u2_u9_X_32, u2_u9_X_34, u2_u9_X_4, u2_u9_X_45, u2_u9_X_46, u2_u9_X_6, u2_uk_K_r11_28, u2_uk_K_r11_48, 
       u2_uk_K_r11_53, u2_uk_K_r13_22, u2_uk_K_r13_32, u2_uk_K_r1_15, u2_uk_K_r1_16, u2_uk_K_r1_18, u2_uk_K_r1_21, u2_uk_K_r1_22, u2_uk_K_r1_47, 
       u2_uk_K_r2_13, u2_uk_K_r2_18, u2_uk_K_r2_21, u2_uk_K_r2_25, u2_uk_K_r2_27, u2_uk_K_r2_28, u2_uk_K_r2_31, u2_uk_K_r2_36, u2_uk_K_r2_49, 
       u2_uk_K_r2_55, u2_uk_K_r3_11, u2_uk_K_r3_14, u2_uk_K_r3_19, u2_uk_K_r3_43, u2_uk_K_r3_9, u2_uk_K_r4_11, u2_uk_K_r4_17, u2_uk_K_r4_33, 
       u2_uk_K_r4_35, u2_uk_K_r4_38, u2_uk_K_r4_4, u2_uk_K_r4_5, u2_uk_K_r4_55, u2_uk_K_r5_10, u2_uk_K_r5_17, u2_uk_K_r5_19, u2_uk_K_r5_39, 
       u2_uk_K_r5_4, u2_uk_K_r5_41, u2_uk_K_r7_0, u2_uk_K_r7_25, u2_uk_K_r7_26, u2_uk_K_r7_32, u2_uk_K_r7_39, u2_uk_K_r7_41, u2_uk_K_r7_48, 
       u2_uk_K_r7_55, u2_uk_K_r8_16, u2_uk_K_r8_2, u2_uk_K_r8_22, u2_uk_K_r8_37, u2_uk_K_r8_41, u2_uk_K_r8_42, u2_uk_K_r9_10, u2_uk_K_r9_4, 
       u2_uk_K_r9_48, u2_uk_n10, u2_uk_n100, u2_uk_n1004, u2_uk_n1008, u2_uk_n102, u2_uk_n1020, u2_uk_n1024, u2_uk_n1027, 
       u2_uk_n1028, u2_uk_n1031, u2_uk_n1035, u2_uk_n1038, u2_uk_n1040, u2_uk_n1043, u2_uk_n1046, u2_uk_n1049, u2_uk_n1050, 
       u2_uk_n1053, u2_uk_n1069, u2_uk_n1074, u2_uk_n1076, u2_uk_n1077, u2_uk_n1079, u2_uk_n1082, u2_uk_n1083, u2_uk_n1084, 
       u2_uk_n1088, u2_uk_n1089, u2_uk_n109, u2_uk_n1091, u2_uk_n1093, u2_uk_n1096, u2_uk_n1098, u2_uk_n11, u2_uk_n110, 
       u2_uk_n1110, u2_uk_n1113, u2_uk_n1120, u2_uk_n1123, u2_uk_n1124, u2_uk_n1128, u2_uk_n1130, u2_uk_n1132, u2_uk_n1133, 
       u2_uk_n1136, u2_uk_n1137, u2_uk_n1140, u2_uk_n1141, u2_uk_n1142, u2_uk_n1152, u2_uk_n117, u2_uk_n1171, u2_uk_n118, 
       u2_uk_n1279, u2_uk_n128, u2_uk_n1280, u2_uk_n1281, u2_uk_n1282, u2_uk_n1283, u2_uk_n1284, u2_uk_n1285, u2_uk_n1286, 
       u2_uk_n1287, u2_uk_n1288, u2_uk_n129, u2_uk_n1290, u2_uk_n1291, u2_uk_n1293, u2_uk_n1295, u2_uk_n1296, u2_uk_n1297, 
       u2_uk_n1300, u2_uk_n1301, u2_uk_n1302, u2_uk_n1305, u2_uk_n1306, u2_uk_n1310, u2_uk_n1311, u2_uk_n1314, u2_uk_n1316, 
       u2_uk_n1317, u2_uk_n1318, u2_uk_n1323, u2_uk_n1324, u2_uk_n1326, u2_uk_n1328, u2_uk_n1329, u2_uk_n1333, u2_uk_n1339, 
       u2_uk_n1341, u2_uk_n1345, u2_uk_n1346, u2_uk_n1350, u2_uk_n1351, u2_uk_n1356, u2_uk_n1359, u2_uk_n1361, u2_uk_n1370, 
       u2_uk_n1375, u2_uk_n1382, u2_uk_n1401, u2_uk_n1405, u2_uk_n1408, u2_uk_n141, u2_uk_n1410, u2_uk_n1413, u2_uk_n142, 
       u2_uk_n1422, u2_uk_n1426, u2_uk_n1428, u2_uk_n1433, u2_uk_n1435, u2_uk_n1438, u2_uk_n1439, u2_uk_n1440, u2_uk_n1441, 
       u2_uk_n1445, u2_uk_n1446, u2_uk_n1447, u2_uk_n145, u2_uk_n1453, u2_uk_n1454, u2_uk_n1456, u2_uk_n1458, u2_uk_n1459, 
       u2_uk_n146, u2_uk_n1462, u2_uk_n1465, u2_uk_n1466, u2_uk_n147, u2_uk_n1470, u2_uk_n1475, u2_uk_n148, u2_uk_n1480, 
       u2_uk_n1486, u2_uk_n1488, u2_uk_n1490, u2_uk_n1493, u2_uk_n1494, u2_uk_n1496, u2_uk_n1497, u2_uk_n1544, u2_uk_n1548, 
       u2_uk_n1549, u2_uk_n155, u2_uk_n1555, u2_uk_n1556, u2_uk_n1563, u2_uk_n1568, u2_uk_n1573, u2_uk_n1580, u2_uk_n1585, 
       u2_uk_n1586, u2_uk_n1592, u2_uk_n1594, u2_uk_n1609, u2_uk_n161, u2_uk_n1615, u2_uk_n162, u2_uk_n1622, u2_uk_n163, 
       u2_uk_n164, u2_uk_n1682, u2_uk_n1683, u2_uk_n1688, u2_uk_n1689, u2_uk_n1693, u2_uk_n17, u2_uk_n1708, u2_uk_n1709, 
       u2_uk_n1720, u2_uk_n1721, u2_uk_n1746, u2_uk_n1769, u2_uk_n1770, u2_uk_n1781, u2_uk_n1785, u2_uk_n1797, u2_uk_n1803, 
       u2_uk_n1807, u2_uk_n1808, u2_uk_n1816, u2_uk_n1817, u2_uk_n1819, u2_uk_n182, u2_uk_n1821, u2_uk_n1824, u2_uk_n1826, 
       u2_uk_n1834, u2_uk_n1840, u2_uk_n1846, u2_uk_n1849, u2_uk_n1851, u2_uk_n1852, u2_uk_n1855, u2_uk_n1856, u2_uk_n187, 
       u2_uk_n188, u2_uk_n191, u2_uk_n202, u2_uk_n203, u2_uk_n207, u2_uk_n208, u2_uk_n209, u2_uk_n213, u2_uk_n214, 
       u2_uk_n217, u2_uk_n220, u2_uk_n222, u2_uk_n223, u2_uk_n230, u2_uk_n231, u2_uk_n238, u2_uk_n240, u2_uk_n257, 
       u2_uk_n27, u2_uk_n299, u2_uk_n301, u2_uk_n305, u2_uk_n308, u2_uk_n31, u2_uk_n313, u2_uk_n319, u2_uk_n335, 
       u2_uk_n373, u2_uk_n386, u2_uk_n408, u2_uk_n415, u2_uk_n421, u2_uk_n454, u2_uk_n456, u2_uk_n467, u2_uk_n503, 
       u2_uk_n504, u2_uk_n515, u2_uk_n520, u2_uk_n60, u2_uk_n63, u2_uk_n665, u2_uk_n682, u2_uk_n689, u2_uk_n83, 
       u2_uk_n92, u2_uk_n93, u2_uk_n939, u2_uk_n94, u2_uk_n942, u2_uk_n943, u2_uk_n945, u2_uk_n946, u2_uk_n955, 
       u2_uk_n958, u2_uk_n959, u2_uk_n963, u2_uk_n985, u2_uk_n986, u2_uk_n987, u2_uk_n99, u2_uk_n991, u2_uk_n993, 
       u2_uk_n995, u2_uk_n998, u2_uk_n999 ;

  des_des_die_0 u0 ( clk, decrypt, desIn, key1, key2, key3, desOut, u0_out0_1, u0_out0_10, u0_out0_11, u0_out0_12, u0_out0_13, u0_out0_14, u0_out0_15, u0_out0_16, 
      u0_out0_17, u0_out0_18, u0_out0_19, u0_out0_2, u0_out0_20, u0_out0_21, u0_out0_22, u0_out0_23, u0_out0_24, 
      u0_out0_25, u0_out0_26, u0_out0_27, u0_out0_28, u0_out0_29, u0_out0_3, u0_out0_30, u0_out0_31, u0_out0_32, 
      u0_out0_4, u0_out0_5, u0_out0_6, u0_out0_7, u0_out0_8, u0_out0_9, u0_out10_1, u0_out10_10, u0_out10_11, 
      u0_out10_12, u0_out10_13, u0_out10_14, u0_out10_15, u0_out10_16, u0_out10_17, u0_out10_18, u0_out10_19, u0_out10_2, 
      u0_out10_20, u0_out10_21, u0_out10_22, u0_out10_23, u0_out10_24, u0_out10_25, u0_out10_26, u0_out10_27, u0_out10_28, 
      u0_out10_29, u0_out10_3, u0_out10_30, u0_out10_31, u0_out10_32, u0_out10_4, u0_out10_5, u0_out10_6, u0_out10_7, 
      u0_out10_8, u0_out10_9, u0_out11_1, u0_out11_10, u0_out11_11, u0_out11_12, u0_out11_13, u0_out11_14, u0_out11_15, 
      u0_out11_16, u0_out11_17, u0_out11_18, u0_out11_19, u0_out11_2, u0_out11_20, u0_out11_21, u0_out11_22, u0_out11_23, 
      u0_out11_24, u0_out11_25, u0_out11_26, u0_out11_27, u0_out11_28, u0_out11_29, u0_out11_3, u0_out11_30, u0_out11_31, 
      u0_out11_32, u0_out11_4, u0_out11_5, u0_out11_6, u0_out11_7, u0_out11_8, u0_out11_9, u0_out12_1, u0_out12_10, 
      u0_out12_11, u0_out12_12, u0_out12_13, u0_out12_14, u0_out12_15, u0_out12_16, u0_out12_17, u0_out12_18, u0_out12_19, 
      u0_out12_2, u0_out12_20, u0_out12_21, u0_out12_22, u0_out12_23, u0_out12_24, u0_out12_25, u0_out12_26, u0_out12_27, 
      u0_out12_28, u0_out12_29, u0_out12_3, u0_out12_30, u0_out12_31, u0_out12_32, u0_out12_4, u0_out12_5, u0_out12_6, 
      u0_out12_7, u0_out12_8, u0_out12_9, u0_out13_1, u0_out13_10, u0_out13_11, u0_out13_12, u0_out13_13, u0_out13_14, 
      u0_out13_15, u0_out13_17, u0_out13_18, u0_out13_19, u0_out13_2, u0_out13_20, u0_out13_21, u0_out13_22, u0_out13_23, 
      u0_out13_25, u0_out13_26, u0_out13_27, u0_out13_28, u0_out13_29, u0_out13_3, u0_out13_31, u0_out13_32, u0_out13_4, 
      u0_out13_5, u0_out13_7, u0_out13_8, u0_out13_9, u0_out14_1, u0_out14_10, u0_out14_11, u0_out14_12, u0_out14_13, 
      u0_out14_14, u0_out14_15, u0_out14_16, u0_out14_18, u0_out14_19, u0_out14_2, u0_out14_20, u0_out14_21, u0_out14_22, 
      u0_out14_24, u0_out14_25, u0_out14_26, u0_out14_27, u0_out14_28, u0_out14_29, u0_out14_3, u0_out14_30, u0_out14_32, 
      u0_out14_4, u0_out14_5, u0_out14_6, u0_out14_7, u0_out14_8, u0_out15_1, u0_out15_10, u0_out15_11, u0_out15_12, 
      u0_out15_13, u0_out15_14, u0_out15_15, u0_out15_16, u0_out15_17, u0_out15_18, u0_out15_19, u0_out15_2, u0_out15_20, 
      u0_out15_21, u0_out15_22, u0_out15_23, u0_out15_24, u0_out15_25, u0_out15_26, u0_out15_27, u0_out15_28, u0_out15_29, 
      u0_out15_3, u0_out15_30, u0_out15_31, u0_out15_32, u0_out15_4, u0_out15_5, u0_out15_6, u0_out15_7, u0_out15_8, 
      u0_out15_9, u0_out1_1, u0_out1_10, u0_out1_11, u0_out1_12, u0_out1_13, u0_out1_14, u0_out1_16, u0_out1_17, 
      u0_out1_18, u0_out1_19, u0_out1_2, u0_out1_20, u0_out1_22, u0_out1_23, u0_out1_24, u0_out1_25, u0_out1_26, 
      u0_out1_28, u0_out1_29, u0_out1_3, u0_out1_30, u0_out1_31, u0_out1_32, u0_out1_4, u0_out1_6, u0_out1_7, 
      u0_out1_8, u0_out1_9, u0_out2_1, u0_out2_10, u0_out2_11, u0_out2_12, u0_out2_13, u0_out2_14, u0_out2_15, 
      u0_out2_16, u0_out2_17, u0_out2_18, u0_out2_19, u0_out2_2, u0_out2_20, u0_out2_21, u0_out2_22, u0_out2_23, 
      u0_out2_24, u0_out2_25, u0_out2_26, u0_out2_27, u0_out2_28, u0_out2_29, u0_out2_3, u0_out2_30, u0_out2_31, 
      u0_out2_32, u0_out2_4, u0_out2_5, u0_out2_6, u0_out2_7, u0_out2_8, u0_out2_9, u0_out3_1, u0_out3_10, 
      u0_out3_11, u0_out3_12, u0_out3_13, u0_out3_14, u0_out3_15, u0_out3_16, u0_out3_17, u0_out3_18, u0_out3_19, 
      u0_out3_2, u0_out3_20, u0_out3_21, u0_out3_22, u0_out3_23, u0_out3_24, u0_out3_25, u0_out3_26, u0_out3_27, 
      u0_out3_28, u0_out3_29, u0_out3_3, u0_out3_30, u0_out3_31, u0_out3_32, u0_out3_4, u0_out3_5, u0_out3_6, 
      u0_out3_7, u0_out3_8, u0_out3_9, u0_out4_1, u0_out4_10, u0_out4_11, u0_out4_13, u0_out4_14, u0_out4_15, 
      u0_out4_16, u0_out4_17, u0_out4_18, u0_out4_19, u0_out4_2, u0_out4_20, u0_out4_21, u0_out4_23, u0_out4_24, 
      u0_out4_25, u0_out4_26, u0_out4_27, u0_out4_28, u0_out4_29, u0_out4_3, u0_out4_30, u0_out4_31, u0_out4_4, 
      u0_out4_5, u0_out4_6, u0_out4_8, u0_out4_9, u0_out5_1, u0_out5_10, u0_out5_11, u0_out5_12, u0_out5_13, 
      u0_out5_14, u0_out5_15, u0_out5_16, u0_out5_17, u0_out5_18, u0_out5_19, u0_out5_2, u0_out5_20, u0_out5_21, 
      u0_out5_22, u0_out5_23, u0_out5_24, u0_out5_25, u0_out5_26, u0_out5_27, u0_out5_28, u0_out5_29, u0_out5_3, 
      u0_out5_30, u0_out5_31, u0_out5_32, u0_out5_4, u0_out5_5, u0_out5_6, u0_out5_7, u0_out5_8, u0_out5_9, 
      u0_out6_1, u0_out6_10, u0_out6_11, u0_out6_13, u0_out6_16, u0_out6_17, u0_out6_18, u0_out6_19, u0_out6_2, 
      u0_out6_20, u0_out6_23, u0_out6_24, u0_out6_26, u0_out6_28, u0_out6_29, u0_out6_30, u0_out6_31, u0_out6_4, 
      u0_out6_6, u0_out6_9, u0_out7_1, u0_out7_10, u0_out7_11, u0_out7_12, u0_out7_13, u0_out7_14, u0_out7_15, 
      u0_out7_16, u0_out7_17, u0_out7_18, u0_out7_19, u0_out7_2, u0_out7_20, u0_out7_21, u0_out7_22, u0_out7_23, 
      u0_out7_24, u0_out7_25, u0_out7_26, u0_out7_27, u0_out7_28, u0_out7_29, u0_out7_3, u0_out7_30, u0_out7_31, 
      u0_out7_32, u0_out7_4, u0_out7_5, u0_out7_6, u0_out7_7, u0_out7_8, u0_out7_9, u0_out8_1, u0_out8_10, 
      u0_out8_11, u0_out8_12, u0_out8_13, u0_out8_14, u0_out8_15, u0_out8_16, u0_out8_17, u0_out8_18, u0_out8_19, 
      u0_out8_2, u0_out8_20, u0_out8_21, u0_out8_22, u0_out8_23, u0_out8_24, u0_out8_25, u0_out8_26, u0_out8_27, 
      u0_out8_28, u0_out8_29, u0_out8_3, u0_out8_30, u0_out8_31, u0_out8_32, u0_out8_4, u0_out8_5, u0_out8_6, 
      u0_out8_7, u0_out8_8, u0_out8_9, u0_out9_1, u0_out9_10, u0_out9_11, u0_out9_12, u0_out9_13, u0_out9_14, 
      u0_out9_15, u0_out9_16, u0_out9_17, u0_out9_18, u0_out9_19, u0_out9_2, u0_out9_20, u0_out9_21, u0_out9_22, 
      u0_out9_23, u0_out9_24, u0_out9_25, u0_out9_26, u0_out9_27, u0_out9_28, u0_out9_29, u0_out9_3, u0_out9_30, 
      u0_out9_31, u0_out9_32, u0_out9_4, u0_out9_5, u0_out9_6, u0_out9_7, u0_out9_8, u0_out9_9, u0_uk_n10, 
      u0_uk_n100, u0_uk_n102, u0_uk_n109, u0_uk_n11, u0_uk_n110, u0_uk_n117, u0_uk_n118, u0_uk_n128, u0_uk_n129, 
      u0_uk_n141, u0_uk_n142, u0_uk_n145, u0_uk_n146, u0_uk_n147, u0_uk_n148, u0_uk_n155, u0_uk_n161, u0_uk_n162, 
      u0_uk_n163, u0_uk_n164, u0_uk_n17, u0_uk_n182, u0_uk_n187, u0_uk_n188, u0_uk_n191, u0_uk_n202, u0_uk_n203, 
      u0_uk_n207, u0_uk_n208, u0_uk_n209, u0_uk_n213, u0_uk_n214, u0_uk_n217, u0_uk_n220, u0_uk_n222, u0_uk_n223, 
      u0_uk_n230, u0_uk_n231, u0_uk_n238, u0_uk_n240, u0_uk_n242, u0_uk_n250, u0_uk_n251, u0_uk_n252, u0_uk_n27, 
      u0_uk_n31, u0_uk_n60, u0_uk_n63, u0_uk_n83, u0_uk_n92, u0_uk_n93, u0_uk_n94, u0_uk_n99, u1_out0_1, 
      u1_out0_10, u1_out0_11, u1_out0_12, u1_out0_13, u1_out0_14, u1_out0_15, u1_out0_16, u1_out0_17, u1_out0_18, 
      u1_out0_19, u1_out0_2, u1_out0_20, u1_out0_21, u1_out0_22, u1_out0_23, u1_out0_24, u1_out0_25, u1_out0_26, 
      u1_out0_27, u1_out0_28, u1_out0_29, u1_out0_3, u1_out0_30, u1_out0_31, u1_out0_32, u1_out0_4, u1_out0_5, 
      u1_out0_6, u1_out0_7, u1_out0_8, u1_out0_9, u1_out10_1, u1_out10_10, u1_out10_11, u1_out10_12, u1_out10_13, 
      u1_out10_14, u1_out10_15, u1_out10_16, u1_out10_17, u1_out10_18, u1_out10_19, u1_out10_2, u1_out10_20, u1_out10_21, 
      u1_out10_22, u1_out10_23, u1_out10_24, u1_out10_25, u1_out10_26, u1_out10_27, u1_out10_28, u1_out10_29, u1_out10_3, 
      u1_out10_30, u1_out10_31, u1_out10_32, u1_out10_4, u1_out10_5, u1_out10_6, u1_out10_7, u1_out10_8, u1_out10_9, 
      u1_out11_1, u1_out11_10, u1_out11_11, u1_out11_12, u1_out11_13, u1_out11_14, u1_out11_15, u1_out11_16, u1_out11_17, 
      u1_out11_18, u1_out11_19, u1_out11_2, u1_out11_20, u1_out11_21, u1_out11_22, u1_out11_23, u1_out11_24, u1_out11_25, 
      u1_out11_26, u1_out11_27, u1_out11_28, u1_out11_29, u1_out11_3, u1_out11_30, u1_out11_31, u1_out11_32, u1_out11_4, 
      u1_out11_5, u1_out11_6, u1_out11_7, u1_out11_8, u1_out11_9, u1_out12_1, u1_out12_10, u1_out12_11, u1_out12_12, 
      u1_out12_13, u1_out12_14, u1_out12_15, u1_out12_16, u1_out12_17, u1_out12_18, u1_out12_19, u1_out12_2, u1_out12_20, 
      u1_out12_21, u1_out12_22, u1_out12_23, u1_out12_24, u1_out12_25, u1_out12_26, u1_out12_27, u1_out12_28, u1_out12_29, 
      u1_out12_3, u1_out12_30, u1_out12_31, u1_out12_32, u1_out12_4, u1_out12_5, u1_out12_6, u1_out12_7, u1_out12_8, 
      u1_out12_9, u1_out13_1, u1_out13_10, u1_out13_11, u1_out13_12, u1_out13_13, u1_out13_14, u1_out13_15, u1_out13_16, 
      u1_out13_17, u1_out13_18, u1_out13_19, u1_out13_2, u1_out13_20, u1_out13_21, u1_out13_22, u1_out13_23, u1_out13_24, 
      u1_out13_25, u1_out13_26, u1_out13_27, u1_out13_28, u1_out13_29, u1_out13_3, u1_out13_30, u1_out13_31, u1_out13_32, 
      u1_out13_4, u1_out13_5, u1_out13_6, u1_out13_7, u1_out13_8, u1_out13_9, u1_out14_1, u1_out14_10, u1_out14_11, 
      u1_out14_12, u1_out14_13, u1_out14_14, u1_out14_15, u1_out14_16, u1_out14_17, u1_out14_18, u1_out14_19, u1_out14_2, 
      u1_out14_20, u1_out14_21, u1_out14_22, u1_out14_23, u1_out14_24, u1_out14_25, u1_out14_26, u1_out14_27, u1_out14_28, 
      u1_out14_29, u1_out14_3, u1_out14_30, u1_out14_31, u1_out14_32, u1_out14_4, u1_out14_5, u1_out14_6, u1_out14_7, 
      u1_out14_8, u1_out14_9, u1_out15_1, u1_out15_10, u1_out15_11, u1_out15_12, u1_out15_13, u1_out15_14, u1_out15_15, 
      u1_out15_16, u1_out15_17, u1_out15_18, u1_out15_19, u1_out15_2, u1_out15_20, u1_out15_21, u1_out15_22, u1_out15_23, 
      u1_out15_24, u1_out15_25, u1_out15_26, u1_out15_27, u1_out15_28, u1_out15_29, u1_out15_3, u1_out15_30, u1_out15_31, 
      u1_out15_32, u1_out15_4, u1_out15_5, u1_out15_6, u1_out15_7, u1_out15_8, u1_out15_9, u1_out1_1, u1_out1_10, 
      u1_out1_11, u1_out1_12, u1_out1_13, u1_out1_14, u1_out1_15, u1_out1_16, u1_out1_17, u1_out1_18, u1_out1_19, 
      u1_out1_2, u1_out1_20, u1_out1_21, u1_out1_22, u1_out1_23, u1_out1_24, u1_out1_25, u1_out1_26, u1_out1_27, 
      u1_out1_28, u1_out1_29, u1_out1_3, u1_out1_30, u1_out1_31, u1_out1_32, u1_out1_4, u1_out1_5, u1_out1_6, 
      u1_out1_7, u1_out1_8, u1_out1_9, u1_out2_1, u1_out2_10, u1_out2_11, u1_out2_12, u1_out2_13, u1_out2_14, 
      u1_out2_15, u1_out2_16, u1_out2_17, u1_out2_18, u1_out2_19, u1_out2_2, u1_out2_20, u1_out2_21, u1_out2_22, 
      u1_out2_23, u1_out2_24, u1_out2_25, u1_out2_26, u1_out2_27, u1_out2_28, u1_out2_29, u1_out2_3, u1_out2_30, 
      u1_out2_31, u1_out2_32, u1_out2_4, u1_out2_5, u1_out2_6, u1_out2_7, u1_out2_8, u1_out2_9, u1_out3_1, 
      u1_out3_10, u1_out3_11, u1_out3_12, u1_out3_13, u1_out3_14, u1_out3_15, u1_out3_16, u1_out3_17, u1_out3_18, 
      u1_out3_19, u1_out3_2, u1_out3_20, u1_out3_21, u1_out3_22, u1_out3_23, u1_out3_24, u1_out3_25, u1_out3_26, 
      u1_out3_27, u1_out3_28, u1_out3_29, u1_out3_3, u1_out3_30, u1_out3_31, u1_out3_32, u1_out3_4, u1_out3_5, 
      u1_out3_6, u1_out3_7, u1_out3_8, u1_out3_9, u1_out4_1, u1_out4_10, u1_out4_11, u1_out4_12, u1_out4_13, 
      u1_out4_14, u1_out4_15, u1_out4_16, u1_out4_17, u1_out4_18, u1_out4_19, u1_out4_2, u1_out4_20, u1_out4_21, 
      u1_out4_22, u1_out4_23, u1_out4_24, u1_out4_25, u1_out4_26, u1_out4_27, u1_out4_28, u1_out4_29, u1_out4_3, 
      u1_out4_30, u1_out4_31, u1_out4_32, u1_out4_4, u1_out4_5, u1_out4_6, u1_out4_7, u1_out4_8, u1_out4_9, 
      u1_out5_1, u1_out5_10, u1_out5_11, u1_out5_12, u1_out5_13, u1_out5_14, u1_out5_15, u1_out5_16, u1_out5_17, 
      u1_out5_18, u1_out5_19, u1_out5_2, u1_out5_20, u1_out5_21, u1_out5_22, u1_out5_23, u1_out5_24, u1_out5_25, 
      u1_out5_26, u1_out5_27, u1_out5_28, u1_out5_29, u1_out5_3, u1_out5_30, u1_out5_31, u1_out5_32, u1_out5_4, 
      u1_out5_5, u1_out5_6, u1_out5_7, u1_out5_8, u1_out5_9, u1_out6_1, u1_out6_10, u1_out6_11, u1_out6_12, 
      u1_out6_13, u1_out6_14, u1_out6_15, u1_out6_16, u1_out6_17, u1_out6_18, u1_out6_19, u1_out6_2, u1_out6_20, 
      u1_out6_21, u1_out6_22, u1_out6_23, u1_out6_24, u1_out6_25, u1_out6_26, u1_out6_27, u1_out6_28, u1_out6_29, 
      u1_out6_3, u1_out6_30, u1_out6_31, u1_out6_32, u1_out6_4, u1_out6_5, u1_out6_6, u1_out6_7, u1_out6_8, 
      u1_out6_9, u1_out7_1, u1_out7_10, u1_out7_11, u1_out7_12, u1_out7_13, u1_out7_14, u1_out7_15, u1_out7_16, 
      u1_out7_17, u1_out7_18, u1_out7_19, u1_out7_2, u1_out7_20, u1_out7_21, u1_out7_22, u1_out7_23, u1_out7_24, 
      u1_out7_25, u1_out7_26, u1_out7_27, u1_out7_28, u1_out7_29, u1_out7_3, u1_out7_30, u1_out7_31, u1_out7_32, 
      u1_out7_4, u1_out7_5, u1_out7_6, u1_out7_7, u1_out7_8, u1_out7_9, u1_out8_1, u1_out8_10, u1_out8_11, 
      u1_out8_12, u1_out8_13, u1_out8_14, u1_out8_15, u1_out8_16, u1_out8_17, u1_out8_18, u1_out8_19, u1_out8_2, 
      u1_out8_20, u1_out8_21, u1_out8_22, u1_out8_23, u1_out8_24, u1_out8_25, u1_out8_26, u1_out8_27, u1_out8_28, 
      u1_out8_29, u1_out8_3, u1_out8_30, u1_out8_31, u1_out8_32, u1_out8_4, u1_out8_5, u1_out8_6, u1_out8_7, 
      u1_out8_8, u1_out8_9, u1_out9_1, u1_out9_10, u1_out9_11, u1_out9_12, u1_out9_13, u1_out9_14, u1_out9_15, 
      u1_out9_16, u1_out9_17, u1_out9_18, u1_out9_19, u1_out9_2, u1_out9_20, u1_out9_21, u1_out9_22, u1_out9_23, 
      u1_out9_24, u1_out9_25, u1_out9_26, u1_out9_27, u1_out9_28, u1_out9_29, u1_out9_3, u1_out9_30, u1_out9_31, 
      u1_out9_32, u1_out9_4, u1_out9_5, u1_out9_6, u1_out9_7, u1_out9_8, u1_out9_9, u2_out0_11, u2_out0_12, 
      u2_out0_13, u2_out0_14, u2_out0_15, u2_out0_18, u2_out0_19, u2_out0_2, u2_out0_21, u2_out0_22, u2_out0_25, 
      u2_out0_27, u2_out0_28, u2_out0_29, u2_out0_3, u2_out0_32, u2_out0_4, u2_out0_5, u2_out0_7, u2_out0_8, 
      u2_out10_1, u2_out10_10, u2_out10_11, u2_out10_12, u2_out10_13, u2_out10_14, u2_out10_15, u2_out10_16, u2_out10_18, 
      u2_out10_19, u2_out10_2, u2_out10_20, u2_out10_21, u2_out10_22, u2_out10_24, u2_out10_25, u2_out10_26, u2_out10_27, 
      u2_out10_28, u2_out10_29, u2_out10_3, u2_out10_30, u2_out10_32, u2_out10_4, u2_out10_5, u2_out10_6, u2_out10_7, 
      u2_out10_8, u2_out11_1, u2_out11_10, u2_out11_11, u2_out11_12, u2_out11_13, u2_out11_14, u2_out11_15, u2_out11_16, 
      u2_out11_17, u2_out11_18, u2_out11_19, u2_out11_2, u2_out11_20, u2_out11_21, u2_out11_22, u2_out11_23, u2_out11_24, 
      u2_out11_25, u2_out11_26, u2_out11_27, u2_out11_28, u2_out11_29, u2_out11_3, u2_out11_30, u2_out11_31, u2_out11_32, 
      u2_out11_4, u2_out11_5, u2_out11_6, u2_out11_7, u2_out11_8, u2_out11_9, u2_out12_11, u2_out12_12, u2_out12_13, 
      u2_out12_14, u2_out12_15, u2_out12_17, u2_out12_18, u2_out12_19, u2_out12_2, u2_out12_21, u2_out12_22, u2_out12_23, 
      u2_out12_25, u2_out12_27, u2_out12_28, u2_out12_29, u2_out12_3, u2_out12_31, u2_out12_32, u2_out12_4, u2_out12_5, 
      u2_out12_7, u2_out12_8, u2_out12_9, u2_out13_11, u2_out13_12, u2_out13_14, u2_out13_15, u2_out13_19, u2_out13_21, 
      u2_out13_22, u2_out13_25, u2_out13_27, u2_out13_29, u2_out13_3, u2_out13_32, u2_out13_4, u2_out13_5, u2_out13_7, 
      u2_out13_8, u2_out14_1, u2_out14_10, u2_out14_11, u2_out14_12, u2_out14_13, u2_out14_14, u2_out14_15, u2_out14_16, 
      u2_out14_17, u2_out14_18, u2_out14_19, u2_out14_2, u2_out14_20, u2_out14_21, u2_out14_22, u2_out14_23, u2_out14_24, 
      u2_out14_25, u2_out14_26, u2_out14_27, u2_out14_28, u2_out14_29, u2_out14_3, u2_out14_30, u2_out14_31, u2_out14_32, 
      u2_out14_4, u2_out14_5, u2_out14_6, u2_out14_7, u2_out14_8, u2_out14_9, u2_out15_1, u2_out15_10, u2_out15_11, 
      u2_out15_12, u2_out15_13, u2_out15_14, u2_out15_15, u2_out15_16, u2_out15_17, u2_out15_18, u2_out15_19, u2_out15_2, 
      u2_out15_20, u2_out15_21, u2_out15_22, u2_out15_23, u2_out15_24, u2_out15_25, u2_out15_26, u2_out15_27, u2_out15_28, 
      u2_out15_29, u2_out15_3, u2_out15_30, u2_out15_31, u2_out15_32, u2_out15_4, u2_out15_5, u2_out15_6, u2_out15_7, 
      u2_out15_8, u2_out15_9, u2_out1_1, u2_out1_10, u2_out1_11, u2_out1_12, u2_out1_13, u2_out1_14, u2_out1_15, 
      u2_out1_16, u2_out1_17, u2_out1_18, u2_out1_19, u2_out1_2, u2_out1_20, u2_out1_21, u2_out1_22, u2_out1_23, 
      u2_out1_24, u2_out1_25, u2_out1_26, u2_out1_27, u2_out1_28, u2_out1_29, u2_out1_3, u2_out1_30, u2_out1_31, 
      u2_out1_32, u2_out1_4, u2_out1_5, u2_out1_6, u2_out1_7, u2_out1_8, u2_out1_9, u2_out2_1, u2_out2_10, 
      u2_out2_11, u2_out2_12, u2_out2_13, u2_out2_14, u2_out2_15, u2_out2_16, u2_out2_17, u2_out2_18, u2_out2_19, 
      u2_out2_2, u2_out2_20, u2_out2_21, u2_out2_22, u2_out2_23, u2_out2_24, u2_out2_25, u2_out2_26, u2_out2_27, 
      u2_out2_28, u2_out2_29, u2_out2_3, u2_out2_30, u2_out2_31, u2_out2_32, u2_out2_4, u2_out2_5, u2_out2_6, 
      u2_out2_7, u2_out2_8, u2_out2_9, u2_out3_1, u2_out3_10, u2_out3_11, u2_out3_13, u2_out3_14, u2_out3_15, 
      u2_out3_16, u2_out3_17, u2_out3_18, u2_out3_19, u2_out3_2, u2_out3_20, u2_out3_21, u2_out3_23, u2_out3_24, 
      u2_out3_25, u2_out3_26, u2_out3_27, u2_out3_28, u2_out3_29, u2_out3_3, u2_out3_30, u2_out3_31, u2_out3_4, 
      u2_out3_5, u2_out3_6, u2_out3_8, u2_out3_9, u2_out4_1, u2_out4_10, u2_out4_11, u2_out4_12, u2_out4_13, 
      u2_out4_14, u2_out4_15, u2_out4_16, u2_out4_17, u2_out4_18, u2_out4_19, u2_out4_2, u2_out4_20, u2_out4_21, 
      u2_out4_22, u2_out4_23, u2_out4_24, u2_out4_25, u2_out4_26, u2_out4_27, u2_out4_28, u2_out4_29, u2_out4_3, 
      u2_out4_30, u2_out4_31, u2_out4_32, u2_out4_4, u2_out4_5, u2_out4_6, u2_out4_7, u2_out4_8, u2_out4_9, 
      u2_out5_1, u2_out5_10, u2_out5_11, u2_out5_12, u2_out5_13, u2_out5_14, u2_out5_15, u2_out5_16, u2_out5_17, 
      u2_out5_18, u2_out5_19, u2_out5_2, u2_out5_20, u2_out5_21, u2_out5_22, u2_out5_23, u2_out5_24, u2_out5_25, 
      u2_out5_26, u2_out5_27, u2_out5_28, u2_out5_29, u2_out5_3, u2_out5_30, u2_out5_31, u2_out5_32, u2_out5_4, 
      u2_out5_5, u2_out5_6, u2_out5_7, u2_out5_8, u2_out5_9, u2_out6_1, u2_out6_10, u2_out6_11, u2_out6_12, 
      u2_out6_13, u2_out6_14, u2_out6_15, u2_out6_16, u2_out6_17, u2_out6_18, u2_out6_19, u2_out6_2, u2_out6_20, 
      u2_out6_21, u2_out6_22, u2_out6_23, u2_out6_24, u2_out6_25, u2_out6_26, u2_out6_27, u2_out6_28, u2_out6_29, 
      u2_out6_3, u2_out6_30, u2_out6_31, u2_out6_32, u2_out6_4, u2_out6_5, u2_out6_6, u2_out6_7, u2_out6_8, 
      u2_out6_9, u2_out7_1, u2_out7_10, u2_out7_13, u2_out7_15, u2_out7_16, u2_out7_17, u2_out7_18, u2_out7_2, 
      u2_out7_20, u2_out7_21, u2_out7_23, u2_out7_24, u2_out7_26, u2_out7_27, u2_out7_28, u2_out7_30, u2_out7_31, 
      u2_out7_5, u2_out7_6, u2_out7_9, u2_out8_1, u2_out8_10, u2_out8_11, u2_out8_12, u2_out8_13, u2_out8_14, 
      u2_out8_15, u2_out8_16, u2_out8_17, u2_out8_18, u2_out8_19, u2_out8_2, u2_out8_20, u2_out8_21, u2_out8_22, 
      u2_out8_23, u2_out8_24, u2_out8_25, u2_out8_26, u2_out8_27, u2_out8_28, u2_out8_29, u2_out8_3, u2_out8_30, 
      u2_out8_31, u2_out8_32, u2_out8_4, u2_out8_5, u2_out8_6, u2_out8_7, u2_out8_8, u2_out8_9, u2_out9_1, 
      u2_out9_10, u2_out9_11, u2_out9_12, u2_out9_13, u2_out9_14, u2_out9_15, u2_out9_16, u2_out9_17, u2_out9_18, 
      u2_out9_19, u2_out9_2, u2_out9_20, u2_out9_21, u2_out9_22, u2_out9_23, u2_out9_24, u2_out9_25, u2_out9_26, 
      u2_out9_27, u2_out9_28, u2_out9_29, u2_out9_3, u2_out9_30, u2_out9_31, u2_out9_32, u2_out9_4, u2_out9_5, 
      u2_out9_6, u2_out9_7, u2_out9_8, u2_out9_9, u2_uk_n10, u2_uk_n100, u2_uk_n102, u2_uk_n109, u2_uk_n11, 
      u2_uk_n110, u2_uk_n117, u2_uk_n118, u2_uk_n128, u2_uk_n129, u2_uk_n141, u2_uk_n142, u2_uk_n145, u2_uk_n146, 
      u2_uk_n147, u2_uk_n148, u2_uk_n155, u2_uk_n161, u2_uk_n162, u2_uk_n163, u2_uk_n164, u2_uk_n17, u2_uk_n182, 
      u2_uk_n187, u2_uk_n188, u2_uk_n191, u2_uk_n202, u2_uk_n203, u2_uk_n207, u2_uk_n208, u2_uk_n209, u2_uk_n213, 
      u2_uk_n214, u2_uk_n217, u2_uk_n220, u2_uk_n222, u2_uk_n223, u2_uk_n230, u2_uk_n231, u2_uk_n27, u2_uk_n31, 
      u2_uk_n60, u2_uk_n63, u2_uk_n83, u2_uk_n92, u2_uk_n93, u2_uk_n94, u2_uk_n99, u0_FP_33, u0_FP_34, 
      u0_FP_36, u0_FP_37, u0_FP_39, u0_FP_41, u0_FP_42, u0_FP_43, u0_FP_44, u0_FP_45, u0_FP_46, 
      u0_FP_48, u0_FP_49, u0_FP_50, u0_FP_51, u0_FP_52, u0_FP_53, u0_FP_55, u0_FP_56, u0_FP_57, 
      u0_FP_58, u0_FP_59, u0_FP_60, u0_FP_63, u0_FP_64, u0_K10_1, u0_K10_14, u0_K10_17, u0_K10_18, 
      u0_K10_19, u0_K10_20, u0_K10_32, u0_K11_37, u0_K11_42, u0_K11_48, u0_K12_19, u0_K12_25, u0_K12_35, 
      u0_K12_36, u0_K12_48, u0_K12_5, u0_K12_7, u0_K12_8, u0_K13_41, u0_K14_23, u0_K14_24, u0_K14_25, 
      u0_K14_26, u0_K14_29, u0_K14_5, u0_K14_7, u0_K15_13, u0_K16_18, u0_K16_19, u0_K16_24, u0_K16_26, 
      u0_K16_36, u0_K16_38, u0_K16_5, u0_K16_8, u0_K1_13, u0_K1_14, u0_K1_17, u0_K1_30, u0_K1_31, 
      u0_K2_11, u0_K2_12, u0_K2_18, u0_K2_20, u0_K2_29, u0_K2_30, u0_K2_31, u0_K2_5, u0_K3_12, 
      u0_K3_13, u0_K3_14, u0_K3_17, u0_K3_18, u0_K3_19, u0_K3_23, u0_K3_5, u0_K3_6, u0_K4_36, 
      u0_K4_43, u0_K4_48, u0_K4_6, u0_K5_1, u0_K5_18, u0_K5_24, u0_K5_26, u0_K5_29, u0_K5_31, 
      u0_K5_47, u0_K5_8, u0_K6_11, u0_K6_13, u0_K6_19, u0_K6_20, u0_K6_23, u0_K6_24, u0_K6_41, 
      u0_K8_11, u0_K8_13, u0_K8_19, u0_K9_12, u0_K9_13, u0_K9_14, u0_K9_30, u0_K9_32, u0_K9_44, 
      u0_K9_6, u0_R0_1, u0_R0_13, u0_R0_15, u0_R0_18, u0_R0_19, u0_R0_20, u0_R0_21, u0_R0_28, 
      u0_R0_32, u0_R0_4, u0_R0_7, u0_R0_8, u0_R0_9, u0_R10_1, u0_R10_12, u0_R10_14, u0_R10_16, 
      u0_R10_17, u0_R10_18, u0_R10_19, u0_R10_2, u0_R10_20, u0_R10_21, u0_R10_24, u0_R10_25, u0_R10_28, 
      u0_R10_29, u0_R10_3, u0_R10_4, u0_R10_5, u0_R11_10, u0_R11_11, u0_R11_12, u0_R11_13, u0_R11_14, 
      u0_R11_15, u0_R11_16, u0_R11_2, u0_R11_20, u0_R11_28, u0_R11_3, u0_R11_32, u0_R11_5, u0_R11_6, 
      u0_R12_16, u0_R12_17, u0_R12_19, u0_R12_20, u0_R12_22, u0_R12_23, u0_R12_24, u0_R12_30, u0_R12_4, 
      u0_R13_17, u0_R13_18, u0_R13_19, u0_R13_20, u0_R13_21, u0_R13_22, u0_R13_23, u0_R13_24, u0_R13_25, 
      u0_R13_26, u0_R13_27, u0_R13_28, u0_R13_29, u0_R13_30, u0_R13_31, u0_R13_8, u0_R1_1, u0_R1_12, 
      u0_R1_13, u0_R1_14, u0_R1_15, u0_R1_16, u0_R1_19, u0_R1_20, u0_R1_21, u0_R1_22, u0_R1_24, 
      u0_R1_25, u0_R1_26, u0_R1_27, u0_R1_28, u0_R1_29, u0_R1_3, u0_R1_30, u0_R1_32, u0_R1_4, 
      u0_R1_5, u0_R1_8, u0_R1_9, u0_R2_1, u0_R2_10, u0_R2_11, u0_R2_12, u0_R2_13, u0_R2_14, 
      u0_R2_16, u0_R2_2, u0_R2_21, u0_R2_22, u0_R2_25, u0_R2_28, u0_R2_3, u0_R2_32, u0_R2_4, 
      u0_R2_5, u0_R2_6, u0_R2_7, u0_R2_8, u0_R2_9, u0_R3_13, u0_R3_15, u0_R3_17, u0_R3_18, 
      u0_R3_20, u0_R3_22, u0_R3_24, u0_R3_25, u0_R3_32, u0_R3_5, u0_R4_1, u0_R4_12, u0_R4_13, 
      u0_R4_16, u0_R4_17, u0_R4_19, u0_R4_20, u0_R4_21, u0_R4_22, u0_R4_24, u0_R4_25, u0_R4_26, 
      u0_R4_27, u0_R4_28, u0_R4_29, u0_R4_3, u0_R4_30, u0_R4_32, u0_R4_4, u0_R4_5, u0_R4_8, 
      u0_R4_9, u0_R5_12, u0_R5_13, u0_R5_2, u0_R5_25, u0_R5_3, u0_R5_32, u0_R5_4, u0_R5_5, 
      u0_R5_7, u0_R5_8, u0_R5_9, u0_R6_10, u0_R6_11, u0_R6_12, u0_R6_13, u0_R6_14, u0_R6_17, 
      u0_R6_24, u0_R6_26, u0_R6_28, u0_R6_29, u0_R6_4, u0_R6_5, u0_R6_7, u0_R6_8, u0_R6_9, 
      u0_R7_1, u0_R7_12, u0_R7_14, u0_R7_17, u0_R7_20, u0_R7_21, u0_R7_22, u0_R7_23, u0_R7_24, 
      u0_R7_25, u0_R7_28, u0_R7_29, u0_R7_32, u0_R7_4, u0_R7_5, u0_R7_8, u0_R7_9, u0_R8_1, 
      u0_R8_12, u0_R8_13, u0_R8_17, u0_R8_19, u0_R8_20, u0_R8_21, u0_R8_22, u0_R8_27, u0_R8_29, 
      u0_R8_30, u0_R8_32, u0_R8_5, u0_R8_6, u0_R8_9, u0_R9_1, u0_R9_10, u0_R9_11, u0_R9_12, 
      u0_R9_13, u0_R9_16, u0_R9_17, u0_R9_18, u0_R9_19, u0_R9_2, u0_R9_20, u0_R9_21, u0_R9_22, 
      u0_R9_24, u0_R9_25, u0_R9_26, u0_R9_27, u0_R9_29, u0_R9_3, u0_R9_30, u0_R9_31, u0_R9_32, 
      u0_R9_4, u0_R9_5, u0_R9_6, u0_R9_7, u0_R9_8, u0_R9_9, u0_desIn_r_1, u0_desIn_r_11, u0_desIn_r_15, 
      u0_desIn_r_17, u0_desIn_r_23, u0_desIn_r_25, u0_desIn_r_27, u0_desIn_r_29, u0_desIn_r_3, u0_desIn_r_31, u0_desIn_r_35, u0_desIn_r_37, 
      u0_desIn_r_39, u0_desIn_r_47, u0_desIn_r_5, u0_desIn_r_51, u0_desIn_r_55, u0_desIn_r_57, u0_desIn_r_59, u0_desIn_r_63, u0_desIn_r_7, 
      u0_desIn_r_9, u0_key_r_0, u0_key_r_11, u0_key_r_12, u0_key_r_13, u0_key_r_14, u0_key_r_16, u0_key_r_19, u0_key_r_2, 
      u0_key_r_20, u0_key_r_21, u0_key_r_22, u0_key_r_23, u0_key_r_28, u0_key_r_29, u0_key_r_30, u0_key_r_35, u0_key_r_4, 
      u0_key_r_41, u0_key_r_42, u0_key_r_47, u0_key_r_48, u0_key_r_5, u0_key_r_50, u0_key_r_54, u0_key_r_55, u0_key_r_6, 
      u0_key_r_9, u0_u0_X_15, u0_u0_X_16, u0_u0_X_21, u0_u0_X_22, u0_u0_X_23, u0_u0_X_25, u0_u0_X_28, u0_u0_X_33, 
      u0_u0_X_42, u0_u0_X_44, u0_u0_X_45, u0_u0_X_46, u0_u10_X_21, u0_u10_X_22, u0_u10_X_34, u0_u10_X_41, u0_u10_X_43, 
      u0_u11_X_1, u0_u11_X_10, u0_u11_X_11, u0_u11_X_12, u0_u11_X_13, u0_u11_X_14, u0_u11_X_15, u0_u11_X_16, u0_u11_X_18, 
      u0_u11_X_20, u0_u11_X_22, u0_u11_X_33, u0_u11_X_34, u0_u11_X_39, u0_u11_X_40, u0_u11_X_45, u0_u11_X_46, u0_u11_X_47, 
      u0_u11_X_9, u0_u12_X_10, u0_u12_X_11, u0_u12_X_12, u0_u12_X_13, u0_u12_X_14, u0_u12_X_2, u0_u12_X_24, u0_u12_X_26, 
      u0_u12_X_27, u0_u12_X_28, u0_u12_X_30, u0_u12_X_32, u0_u12_X_33, u0_u12_X_34, u0_u12_X_35, u0_u12_X_36, u0_u12_X_37, 
      u0_u12_X_38, u0_u12_X_39, u0_u12_X_40, u0_u12_X_42, u0_u12_X_44, u0_u12_X_45, u0_u12_X_46, u0_u12_X_48, u0_u12_X_5, 
      u0_u12_X_7, u0_u13_X_1, u0_u13_X_10, u0_u13_X_11, u0_u13_X_12, u0_u13_X_19, u0_u13_X_2, u0_u13_X_20, u0_u13_X_21, 
      u0_u13_X_22, u0_u13_X_27, u0_u13_X_3, u0_u13_X_30, u0_u13_X_32, u0_u13_X_36, u0_u13_X_38, u0_u13_X_39, u0_u13_X_4, 
      u0_u13_X_40, u0_u13_X_41, u0_u13_X_42, u0_u13_X_43, u0_u13_X_44, u0_u13_X_46, u0_u13_X_47, u0_u13_X_48, u0_u13_X_6, 
      u0_u13_X_8, u0_u13_X_9, u0_u14_X_10, u0_u14_X_12, u0_u14_X_14, u0_u14_X_15, u0_u14_X_16, u0_u14_X_17, u0_u14_X_18, 
      u0_u14_X_19, u0_u14_X_20, u0_u14_X_21, u0_u14_X_22, u0_u14_X_23, u0_u14_X_24, u0_u14_X_25, u0_u14_X_47, u0_u14_X_48, 
      u0_u14_X_7, u0_u14_X_8, u0_u14_X_9, u0_u15_X_11, u0_u15_X_13, u0_u15_X_22, u0_u15_X_33, u0_u15_X_4, u0_u15_X_42, 
      u0_u15_X_44, u0_u15_X_45, u0_u15_X_9, u0_u1_X_15, u0_u1_X_16, u0_u1_X_17, u0_u1_X_19, u0_u1_X_21, u0_u1_X_23, 
      u0_u1_X_24, u0_u1_X_25, u0_u1_X_26, u0_u1_X_3, u0_u1_X_33, u0_u1_X_34, u0_u1_X_35, u0_u1_X_36, u0_u1_X_37, 
      u0_u1_X_38, u0_u1_X_39, u0_u1_X_4, u0_u1_X_40, u0_u1_X_42, u0_u1_X_6, u0_u1_X_8, u0_u1_X_9, u0_u2_X_10, 
      u0_u2_X_15, u0_u2_X_16, u0_u2_X_24, u0_u2_X_26, u0_u2_X_27, u0_u2_X_3, u0_u2_X_34, u0_u2_X_46, u0_u2_X_9, 
      u0_u3_X_22, u0_u3_X_24, u0_u3_X_26, u0_u3_X_27, u0_u3_X_28, u0_u3_X_29, u0_u3_X_31, u0_u3_X_34, u0_u3_X_35, 
      u0_u3_X_37, u0_u3_X_39, u0_u3_X_40, u0_u3_X_42, u0_u3_X_44, u0_u3_X_45, u0_u3_X_46, u0_u4_X_10, u0_u4_X_11, 
      u0_u4_X_12, u0_u4_X_13, u0_u4_X_14, u0_u4_X_15, u0_u4_X_16, u0_u4_X_17, u0_u4_X_19, u0_u4_X_2, u0_u4_X_21, 
      u0_u4_X_23, u0_u4_X_25, u0_u4_X_28, u0_u4_X_3, u0_u4_X_30, u0_u4_X_32, u0_u4_X_34, u0_u4_X_4, u0_u4_X_43, 
      u0_u4_X_44, u0_u4_X_45, u0_u4_X_46, u0_u4_X_48, u0_u4_X_5, u0_u4_X_7, u0_u4_X_9, u0_u5_X_10, u0_u5_X_15, 
      u0_u5_X_16, u0_u5_X_21, u0_u5_X_22, u0_u5_X_27, u0_u5_X_3, u0_u5_X_34, u0_u5_X_46, u0_u5_X_9, u0_u6_X_15, 
      u0_u6_X_16, u0_u6_X_2, u0_u6_X_21, u0_u6_X_22, u0_u6_X_23, u0_u6_X_24, u0_u6_X_31, u0_u6_X_32, u0_u6_X_33, 
      u0_u6_X_34, u0_u6_X_35, u0_u6_X_9, u0_u7_X_1, u0_u7_X_2, u0_u7_X_22, u0_u7_X_23, u0_u7_X_25, u0_u7_X_27, 
      u0_u7_X_28, u0_u7_X_29, u0_u7_X_3, u0_u7_X_30, u0_u7_X_31, u0_u7_X_32, u0_u7_X_33, u0_u7_X_34, u0_u7_X_36, 
      u0_u7_X_38, u0_u7_X_4, u0_u7_X_40, u0_u7_X_45, u0_u7_X_46, u0_u7_X_47, u0_u7_X_48, u0_u7_X_9, u0_u8_X_10, 
      u0_u8_X_15, u0_u8_X_16, u0_u8_X_18, u0_u8_X_20, u0_u8_X_22, u0_u8_X_23, u0_u8_X_25, u0_u8_X_27, u0_u8_X_28, 
      u0_u8_X_3, u0_u8_X_39, u0_u8_X_4, u0_u8_X_40, u0_u8_X_45, u0_u8_X_46, u0_u8_X_9, u0_u9_X_10, u0_u9_X_11, 
      u0_u9_X_13, u0_u9_X_15, u0_u9_X_16, u0_u9_X_21, u0_u9_X_22, u0_u9_X_23, u0_u9_X_25, u0_u9_X_27, u0_u9_X_3, 
      u0_u9_X_34, u0_u9_X_35, u0_u9_X_36, u0_u9_X_37, u0_u9_X_38, u0_u9_X_39, u0_u9_X_4, u0_u9_X_41, u0_u9_X_43, 
      u0_u9_X_46, u0_u9_X_5, u0_u9_X_7, u0_uk_K_r0_15, u0_uk_K_r0_28, u0_uk_K_r0_36, u0_uk_K_r0_49, u0_uk_K_r0_7, u0_uk_K_r10_10, 
      u0_uk_K_r10_18, u0_uk_K_r10_23, u0_uk_K_r10_27, u0_uk_K_r10_28, u0_uk_K_r10_32, u0_uk_K_r10_37, u0_uk_K_r10_41, u0_uk_K_r10_42, u0_uk_K_r10_44, 
      u0_uk_K_r10_9, u0_uk_K_r11_19, u0_uk_K_r11_20, u0_uk_K_r11_24, u0_uk_K_r11_25, u0_uk_K_r11_27, u0_uk_K_r11_29, u0_uk_K_r11_33, u0_uk_K_r11_39, 
      u0_uk_K_r11_4, u0_uk_K_r12_16, u0_uk_K_r13_0, u0_uk_K_r13_25, u0_uk_K_r13_38, u0_uk_K_r13_44, u0_uk_K_r14_10, u0_uk_K_r14_11, u0_uk_K_r14_12, 
      u0_uk_K_r14_15, u0_uk_K_r14_16, u0_uk_K_r14_18, u0_uk_K_r14_2, u0_uk_K_r14_45, u0_uk_K_r14_50, u0_uk_K_r14_8, u0_uk_K_r14_9, u0_uk_K_r1_15, 
      u0_uk_K_r1_16, u0_uk_K_r1_21, u0_uk_K_r1_44, u0_uk_K_r1_7, u0_uk_K_r2_13, u0_uk_K_r2_18, u0_uk_K_r2_20, u0_uk_K_r2_25, u0_uk_K_r2_26, 
      u0_uk_K_r2_27, u0_uk_K_r2_28, u0_uk_K_r2_33, u0_uk_K_r2_4, u0_uk_K_r2_41, u0_uk_K_r2_46, u0_uk_K_r2_50, u0_uk_K_r2_53, u0_uk_K_r2_55, 
      u0_uk_K_r3_10, u0_uk_K_r3_14, u0_uk_K_r4_0, u0_uk_K_r4_23, u0_uk_K_r4_33, u0_uk_K_r4_35, u0_uk_K_r4_38, u0_uk_K_r4_41, u0_uk_K_r4_47, 
      u0_uk_K_r5_10, u0_uk_K_r5_17, u0_uk_K_r5_39, u0_uk_K_r5_4, u0_uk_K_r6_0, u0_uk_K_r6_22, u0_uk_K_r6_26, u0_uk_K_r6_31, u0_uk_K_r6_34, 
      u0_uk_K_r6_46, u0_uk_K_r7_26, u0_uk_K_r8_16, u0_uk_K_r8_40, u0_uk_K_r8_41, u0_uk_K_r9_0, u0_uk_K_r9_1, u0_uk_K_r9_19, u0_uk_K_r9_22, 
      u0_uk_K_r9_25, u0_uk_K_r9_27, u0_uk_K_r9_30, u0_uk_K_r9_33, u0_uk_K_r9_35, u0_uk_K_r9_45, u0_uk_K_r9_6, u0_uk_K_r9_7, u0_uk_K_r9_9, 
      u0_uk_n1000, u0_uk_n1001, u0_uk_n1002, u0_uk_n1004, u0_uk_n1005, u0_uk_n1006, u0_uk_n101, u0_uk_n1012, u0_uk_n1024, 
      u0_uk_n106, u0_uk_n107, u0_uk_n108, u0_uk_n113, u0_uk_n115, u0_uk_n116, u0_uk_n12, u0_uk_n121, u0_uk_n122, 
      u0_uk_n123, u0_uk_n126, u0_uk_n127, u0_uk_n13, u0_uk_n131, u0_uk_n139, u0_uk_n143, u0_uk_n144, u0_uk_n151, 
      u0_uk_n153, u0_uk_n156, u0_uk_n167, u0_uk_n168, u0_uk_n171, u0_uk_n172, u0_uk_n173, u0_uk_n174, u0_uk_n177, 
      u0_uk_n178, u0_uk_n179, u0_uk_n18, u0_uk_n180, u0_uk_n181, u0_uk_n183, u0_uk_n184, u0_uk_n185, u0_uk_n189, 
      u0_uk_n190, u0_uk_n192, u0_uk_n193, u0_uk_n195, u0_uk_n196, u0_uk_n197, u0_uk_n198, u0_uk_n199, u0_uk_n200, 
      u0_uk_n201, u0_uk_n204, u0_uk_n205, u0_uk_n206, u0_uk_n21, u0_uk_n210, u0_uk_n211, u0_uk_n212, u0_uk_n215, 
      u0_uk_n216, u0_uk_n218, u0_uk_n219, u0_uk_n22, u0_uk_n221, u0_uk_n224, u0_uk_n225, u0_uk_n23, u0_uk_n232, 
      u0_uk_n233, u0_uk_n239, u0_uk_n241, u0_uk_n243, u0_uk_n244, u0_uk_n248, u0_uk_n249, u0_uk_n253, u0_uk_n257, 
      u0_uk_n259, u0_uk_n260, u0_uk_n261, u0_uk_n264, u0_uk_n266, u0_uk_n267, u0_uk_n269, u0_uk_n272, u0_uk_n275, 
      u0_uk_n276, u0_uk_n278, u0_uk_n28, u0_uk_n282, u0_uk_n283, u0_uk_n285, u0_uk_n289, u0_uk_n290, u0_uk_n293, 
      u0_uk_n3, u0_uk_n300, u0_uk_n307, u0_uk_n310, u0_uk_n314, u0_uk_n316, u0_uk_n318, u0_uk_n32, u0_uk_n320, 
      u0_uk_n324, u0_uk_n329, u0_uk_n33, u0_uk_n330, u0_uk_n331, u0_uk_n332, u0_uk_n336, u0_uk_n337, u0_uk_n339, 
      u0_uk_n341, u0_uk_n344, u0_uk_n347, u0_uk_n348, u0_uk_n352, u0_uk_n355, u0_uk_n358, u0_uk_n361, u0_uk_n370, 
      u0_uk_n371, u0_uk_n383, u0_uk_n384, u0_uk_n39, u0_uk_n392, u0_uk_n393, u0_uk_n396, u0_uk_n4, u0_uk_n40, 
      u0_uk_n400, u0_uk_n401, u0_uk_n405, u0_uk_n41, u0_uk_n410, u0_uk_n411, u0_uk_n412, u0_uk_n413, u0_uk_n414, 
      u0_uk_n418, u0_uk_n419, u0_uk_n420, u0_uk_n423, u0_uk_n424, u0_uk_n425, u0_uk_n426, u0_uk_n428, u0_uk_n429, 
      u0_uk_n430, u0_uk_n432, u0_uk_n433, u0_uk_n434, u0_uk_n436, u0_uk_n438, u0_uk_n439, u0_uk_n440, u0_uk_n442, 
      u0_uk_n445, u0_uk_n446, u0_uk_n447, u0_uk_n448, u0_uk_n45, u0_uk_n450, u0_uk_n457, u0_uk_n471, u0_uk_n497, 
      u0_uk_n499, u0_uk_n5, u0_uk_n502, u0_uk_n505, u0_uk_n508, u0_uk_n510, u0_uk_n511, u0_uk_n513, u0_uk_n517, 
      u0_uk_n519, u0_uk_n522, u0_uk_n523, u0_uk_n525, u0_uk_n529, u0_uk_n530, u0_uk_n531, u0_uk_n532, u0_uk_n534, 
      u0_uk_n535, u0_uk_n536, u0_uk_n539, u0_uk_n542, u0_uk_n544, u0_uk_n545, u0_uk_n546, u0_uk_n547, u0_uk_n549, 
      u0_uk_n55, u0_uk_n550, u0_uk_n552, u0_uk_n553, u0_uk_n554, u0_uk_n555, u0_uk_n557, u0_uk_n558, u0_uk_n560, 
      u0_uk_n561, u0_uk_n562, u0_uk_n565, u0_uk_n566, u0_uk_n567, u0_uk_n568, u0_uk_n570, u0_uk_n573, u0_uk_n574, 
      u0_uk_n575, u0_uk_n577, u0_uk_n578, u0_uk_n579, u0_uk_n58, u0_uk_n580, u0_uk_n581, u0_uk_n583, u0_uk_n598, 
      u0_uk_n604, u0_uk_n61, u0_uk_n615, u0_uk_n627, u0_uk_n629, u0_uk_n632, u0_uk_n635, u0_uk_n636, u0_uk_n637, 
      u0_uk_n639, u0_uk_n640, u0_uk_n642, u0_uk_n643, u0_uk_n644, u0_uk_n645, u0_uk_n649, u0_uk_n650, u0_uk_n651, 
      u0_uk_n652, u0_uk_n653, u0_uk_n654, u0_uk_n657, u0_uk_n658, u0_uk_n659, u0_uk_n660, u0_uk_n661, u0_uk_n663, 
      u0_uk_n666, u0_uk_n668, u0_uk_n669, u0_uk_n67, u0_uk_n670, u0_uk_n674, u0_uk_n675, u0_uk_n684, u0_uk_n687, 
      u0_uk_n690, u0_uk_n696, u0_uk_n697, u0_uk_n699, u0_uk_n711, u0_uk_n719, u0_uk_n722, u0_uk_n723, u0_uk_n725, 
      u0_uk_n726, u0_uk_n727, u0_uk_n729, u0_uk_n73, u0_uk_n731, u0_uk_n734, u0_uk_n735, u0_uk_n741, u0_uk_n746, 
      u0_uk_n748, u0_uk_n751, u0_uk_n759, u0_uk_n761, u0_uk_n763, u0_uk_n768, u0_uk_n780, u0_uk_n783, u0_uk_n786, 
      u0_uk_n793, u0_uk_n799, u0_uk_n8, u0_uk_n800, u0_uk_n809, u0_uk_n810, u0_uk_n813, u0_uk_n815, u0_uk_n816, 
      u0_uk_n832, u0_uk_n839, u0_uk_n855, u0_uk_n866, u0_uk_n868, u0_uk_n869, u0_uk_n875, u0_uk_n883, u0_uk_n892, 
      u0_uk_n898, u0_uk_n9, u0_uk_n904, u0_uk_n91, u0_uk_n915, u0_uk_n916, u0_uk_n917, u0_uk_n918, u0_uk_n933, 
      u0_uk_n934, u0_uk_n949, u0_uk_n950, u0_uk_n956, u0_uk_n96, u0_uk_n963, u0_uk_n976, u0_uk_n98, u0_uk_n982, 
      u0_uk_n985, u0_uk_n990, u0_uk_n999, u1_FP_33, u1_FP_37, u1_FP_40, u1_FP_41, u1_FP_44, u1_FP_45, 
      u1_FP_52, u1_FP_53, u1_FP_55, u1_FP_56, u1_FP_60, u1_FP_61, u1_K10_1, u1_K10_11, u1_K10_13, 
      u1_K10_14, u1_K10_18, u1_K10_2, u1_K10_20, u1_K10_23, u1_K10_24, u1_K10_25, u1_K10_26, u1_K10_29, 
      u1_K10_30, u1_K10_31, u1_K10_32, u1_K10_36, u1_K10_41, u1_K10_42, u1_K10_43, u1_K10_44, u1_K10_47, 
      u1_K10_48, u1_K10_5, u1_K10_6, u1_K10_7, u1_K10_8, u1_K11_11, u1_K11_13, u1_K11_2, u1_K11_23, 
      u1_K11_25, u1_K11_29, u1_K11_32, u1_K11_35, u1_K11_37, u1_K11_38, u1_K11_48, u1_K11_7, u1_K12_18, 
      u1_K12_19, u1_K12_2, u1_K12_20, u1_K12_24, u1_K12_25, u1_K12_26, u1_K12_35, u1_K12_36, u1_K12_37, 
      u1_K12_38, u1_K12_41, u1_K12_43, u1_K12_47, u1_K12_48, u1_K12_6, u1_K12_8, u1_K13_14, u1_K13_17, 
      u1_K13_18, u1_K13_20, u1_K13_29, u1_K13_30, u1_K13_31, u1_K13_32, u1_K13_35, u1_K13_37, u1_K13_48, 
      u1_K13_8, u1_K14_1, u1_K14_2, u1_K14_29, u1_K14_30, u1_K14_31, u1_K14_32, u1_K14_42, u1_K14_44, 
      u1_K14_47, u1_K14_48, u1_K15_11, u1_K15_12, u1_K15_13, u1_K15_14, u1_K15_18, u1_K15_2, u1_K15_20, 
      u1_K15_23, u1_K15_24, u1_K15_25, u1_K15_29, u1_K15_31, u1_K15_32, u1_K15_35, u1_K15_36, u1_K15_37, 
      u1_K15_41, u1_K15_42, u1_K15_44, u1_K15_48, u1_K15_5, u1_K15_6, u1_K15_7, u1_K16_11, u1_K16_12, 
      u1_K16_13, u1_K16_14, u1_K16_17, u1_K16_18, u1_K16_19, u1_K16_2, u1_K16_20, u1_K16_30, u1_K16_31, 
      u1_K16_32, u1_K16_35, u1_K16_41, u1_K16_42, u1_K16_44, u1_K16_48, u1_K16_6, u1_K16_8, u1_K1_1, 
      u1_K1_17, u1_K1_19, u1_K1_43, u1_K1_47, u1_K1_6, u1_K1_8, u1_K2_1, u1_K2_11, u1_K2_12, 
      u1_K2_13, u1_K2_17, u1_K2_18, u1_K2_2, u1_K2_20, u1_K2_23, u1_K2_24, u1_K2_25, u1_K2_26, 
      u1_K2_29, u1_K2_30, u1_K2_31, u1_K2_42, u1_K2_43, u1_K2_44, u1_K2_47, u1_K2_48, u1_K2_5, 
      u1_K2_6, u1_K2_8, u1_K3_1, u1_K3_12, u1_K3_14, u1_K3_17, u1_K3_18, u1_K3_19, u1_K3_2, 
      u1_K3_20, u1_K3_23, u1_K3_25, u1_K3_26, u1_K3_29, u1_K3_31, u1_K3_35, u1_K3_36, u1_K3_37, 
      u1_K3_38, u1_K3_41, u1_K3_42, u1_K3_43, u1_K3_44, u1_K3_47, u1_K3_48, u1_K3_5, u1_K3_6, 
      u1_K3_7, u1_K3_8, u1_K4_1, u1_K4_11, u1_K4_12, u1_K4_13, u1_K4_14, u1_K4_17, u1_K4_18, 
      u1_K4_19, u1_K4_24, u1_K4_30, u1_K4_32, u1_K4_35, u1_K4_36, u1_K4_37, u1_K4_38, u1_K4_41, 
      u1_K4_42, u1_K4_43, u1_K4_44, u1_K4_47, u1_K4_48, u1_K4_6, u1_K5_1, u1_K5_11, u1_K5_12, 
      u1_K5_13, u1_K5_14, u1_K5_17, u1_K5_18, u1_K5_19, u1_K5_2, u1_K5_23, u1_K5_24, u1_K5_25, 
      u1_K5_26, u1_K5_29, u1_K5_30, u1_K5_31, u1_K5_32, u1_K5_37, u1_K5_38, u1_K5_41, u1_K5_42, 
      u1_K5_44, u1_K5_47, u1_K5_48, u1_K5_5, u1_K5_6, u1_K5_7, u1_K5_8, u1_K6_1, u1_K6_11, 
      u1_K6_12, u1_K6_13, u1_K6_14, u1_K6_20, u1_K6_23, u1_K6_24, u1_K6_25, u1_K6_26, u1_K6_29, 
      u1_K6_30, u1_K6_31, u1_K6_32, u1_K6_35, u1_K6_36, u1_K6_37, u1_K6_38, u1_K6_41, u1_K6_42, 
      u1_K6_43, u1_K6_44, u1_K6_47, u1_K6_48, u1_K6_5, u1_K6_6, u1_K6_7, u1_K6_8, u1_K7_1, 
      u1_K7_11, u1_K7_14, u1_K7_17, u1_K7_18, u1_K7_19, u1_K7_2, u1_K7_23, u1_K7_26, u1_K7_29, 
      u1_K7_30, u1_K7_31, u1_K7_35, u1_K7_37, u1_K7_38, u1_K7_41, u1_K7_43, u1_K7_44, u1_K7_47, 
      u1_K7_48, u1_K7_5, u1_K7_7, u1_K8_1, u1_K8_11, u1_K8_13, u1_K8_14, u1_K8_18, u1_K8_2, 
      u1_K8_20, u1_K8_23, u1_K8_24, u1_K8_25, u1_K8_26, u1_K8_30, u1_K8_31, u1_K8_32, u1_K8_35, 
      u1_K8_36, u1_K8_38, u1_K8_41, u1_K8_42, u1_K8_44, u1_K8_47, u1_K8_48, u1_K8_5, u1_K8_7, 
      u1_K9_12, u1_K9_13, u1_K9_14, u1_K9_17, u1_K9_23, u1_K9_24, u1_K9_25, u1_K9_29, u1_K9_31, 
      u1_K9_36, u1_K9_37, u1_K9_38, u1_K9_43, u1_K9_44, u1_K9_47, u1_K9_5, u1_K9_6, u1_K9_7, 
      u1_K9_8, u1_R0_1, u1_R0_12, u1_R0_13, u1_R0_16, u1_R0_17, u1_R0_20, u1_R0_21, u1_R0_28, 
      u1_R0_29, u1_R0_32, u1_R0_4, u1_R0_5, u1_R0_7, u1_R0_8, u1_R0_9, u1_R10_1, u1_R10_10, 
      u1_R10_12, u1_R10_13, u1_R10_14, u1_R10_16, u1_R10_17, u1_R10_24, u1_R10_25, u1_R10_28, u1_R10_29, 
      u1_R10_32, u1_R10_5, u1_R11_1, u1_R11_10, u1_R11_12, u1_R11_13, u1_R11_20, u1_R11_21, u1_R11_24, 
      u1_R11_4, u1_R11_5, u1_R11_8, u1_R11_9, u1_R12_1, u1_R12_20, u1_R12_21, u1_R12_23, u1_R12_29, 
      u1_R12_32, u1_R13_1, u1_R13_13, u1_R13_16, u1_R13_17, u1_R13_20, u1_R13_21, u1_R13_24, u1_R13_25, 
      u1_R13_28, u1_R13_29, u1_R13_4, u1_R13_5, u1_R13_8, u1_R13_9, u1_R1_1, u1_R1_12, u1_R1_13, 
      u1_R1_16, u1_R1_17, u1_R1_20, u1_R1_24, u1_R1_25, u1_R1_28, u1_R1_29, u1_R1_32, u1_R1_4, 
      u1_R1_5, u1_R1_9, u1_R2_1, u1_R2_12, u1_R2_13, u1_R2_16, u1_R2_17, u1_R2_2, u1_R2_20, 
      u1_R2_21, u1_R2_24, u1_R2_25, u1_R2_28, u1_R2_29, u1_R2_32, u1_R2_5, u1_R2_7, u1_R2_8, 
      u1_R2_9, u1_R3_1, u1_R3_12, u1_R3_13, u1_R3_15, u1_R3_16, u1_R3_17, u1_R3_18, u1_R3_20, 
      u1_R3_21, u1_R3_24, u1_R3_25, u1_R3_28, u1_R3_29, u1_R3_32, u1_R3_4, u1_R3_5, u1_R3_8, 
      u1_R3_9, u1_R4_1, u1_R4_13, u1_R4_14, u1_R4_16, u1_R4_17, u1_R4_20, u1_R4_21, u1_R4_24, 
      u1_R4_25, u1_R4_28, u1_R4_29, u1_R4_3, u1_R4_32, u1_R4_4, u1_R4_5, u1_R4_6, u1_R4_7, 
      u1_R4_8, u1_R4_9, u1_R5_1, u1_R5_12, u1_R5_13, u1_R5_16, u1_R5_17, u1_R5_18, u1_R5_20, 
      u1_R5_21, u1_R5_23, u1_R5_24, u1_R5_25, u1_R5_28, u1_R5_29, u1_R5_31, u1_R5_32, u1_R5_4, 
      u1_R5_5, u1_R5_8, u1_R5_9, u1_R6_1, u1_R6_10, u1_R6_13, u1_R6_16, u1_R6_17, u1_R6_2, 
      u1_R6_20, u1_R6_21, u1_R6_24, u1_R6_25, u1_R6_28, u1_R6_29, u1_R6_32, u1_R6_4, u1_R6_8, 
      u1_R6_9, u1_R7_1, u1_R7_12, u1_R7_13, u1_R7_15, u1_R7_16, u1_R7_17, u1_R7_18, u1_R7_20, 
      u1_R7_24, u1_R7_25, u1_R7_28, u1_R7_29, u1_R7_32, u1_R7_4, u1_R7_5, u1_R7_6, u1_R7_7, 
      u1_R7_8, u1_R7_9, u1_R8_1, u1_R8_13, u1_R8_15, u1_R8_16, u1_R8_17, u1_R8_20, u1_R8_21, 
      u1_R8_22, u1_R8_24, u1_R8_25, u1_R8_28, u1_R8_29, u1_R8_32, u1_R8_4, u1_R8_5, u1_R8_6, 
      u1_R8_8, u1_R8_9, u1_R9_1, u1_R9_12, u1_R9_15, u1_R9_16, u1_R9_20, u1_R9_21, u1_R9_23, 
      u1_R9_24, u1_R9_25, u1_R9_4, u1_R9_8, u1_R9_9, u1_desIn_r_25, u1_desIn_r_29, u1_desIn_r_37, u1_desIn_r_39, 
      u1_desIn_r_57, u1_u0_X_10, u1_u0_X_11, u1_u0_X_12, u1_u0_X_13, u1_u0_X_14, u1_u0_X_15, u1_u0_X_16, u1_u0_X_2, 
      u1_u0_X_21, u1_u0_X_22, u1_u0_X_23, u1_u0_X_24, u1_u0_X_25, u1_u0_X_26, u1_u0_X_27, u1_u0_X_28, u1_u0_X_29, 
      u1_u0_X_3, u1_u0_X_30, u1_u0_X_31, u1_u0_X_32, u1_u0_X_33, u1_u0_X_34, u1_u0_X_35, u1_u0_X_36, u1_u0_X_37, 
      u1_u0_X_38, u1_u0_X_39, u1_u0_X_4, u1_u0_X_40, u1_u0_X_42, u1_u0_X_44, u1_u0_X_45, u1_u0_X_46, u1_u0_X_48, 
      u1_u0_X_5, u1_u0_X_7, u1_u0_X_9, u1_u10_X_1, u1_u10_X_10, u1_u10_X_15, u1_u10_X_16, u1_u10_X_18, u1_u10_X_20, 
      u1_u10_X_21, u1_u10_X_24, u1_u10_X_26, u1_u10_X_27, u1_u10_X_28, u1_u10_X_3, u1_u10_X_33, u1_u10_X_39, u1_u10_X_4, 
      u1_u10_X_40, u1_u10_X_41, u1_u10_X_42, u1_u10_X_43, u1_u10_X_44, u1_u10_X_45, u1_u10_X_46, u1_u10_X_47, u1_u10_X_6, 
      u1_u10_X_8, u1_u10_X_9, u1_u11_X_10, u1_u11_X_11, u1_u11_X_12, u1_u11_X_13, u1_u11_X_14, u1_u11_X_16, u1_u11_X_22, 
      u1_u11_X_27, u1_u11_X_28, u1_u11_X_29, u1_u11_X_3, u1_u11_X_30, u1_u11_X_31, u1_u11_X_32, u1_u11_X_33, u1_u11_X_34, 
      u1_u11_X_39, u1_u11_X_4, u1_u11_X_40, u1_u11_X_45, u1_u11_X_46, u1_u11_X_5, u1_u11_X_7, u1_u11_X_9, u1_u12_X_1, 
      u1_u12_X_10, u1_u12_X_16, u1_u12_X_21, u1_u12_X_22, u1_u12_X_23, u1_u12_X_24, u1_u12_X_25, u1_u12_X_26, u1_u12_X_27, 
      u1_u12_X_28, u1_u12_X_3, u1_u12_X_33, u1_u12_X_34, u1_u12_X_36, u1_u12_X_38, u1_u12_X_39, u1_u12_X_4, u1_u12_X_40, 
      u1_u12_X_41, u1_u12_X_42, u1_u12_X_43, u1_u12_X_44, u1_u12_X_45, u1_u12_X_46, u1_u12_X_47, u1_u12_X_9, u1_u13_X_10, 
      u1_u13_X_11, u1_u13_X_12, u1_u13_X_13, u1_u13_X_14, u1_u13_X_15, u1_u13_X_16, u1_u13_X_17, u1_u13_X_18, u1_u13_X_19, 
      u1_u13_X_20, u1_u13_X_21, u1_u13_X_22, u1_u13_X_23, u1_u13_X_24, u1_u13_X_25, u1_u13_X_26, u1_u13_X_27, u1_u13_X_28, 
      u1_u13_X_3, u1_u13_X_33, u1_u13_X_35, u1_u13_X_36, u1_u13_X_37, u1_u13_X_38, u1_u13_X_39, u1_u13_X_4, u1_u13_X_40, 
      u1_u13_X_41, u1_u13_X_43, u1_u13_X_45, u1_u13_X_46, u1_u13_X_5, u1_u13_X_6, u1_u13_X_7, u1_u13_X_8, u1_u13_X_9, 
      u1_u14_X_1, u1_u14_X_10, u1_u14_X_15, u1_u14_X_16, u1_u14_X_17, u1_u14_X_19, u1_u14_X_21, u1_u14_X_22, u1_u14_X_27, 
      u1_u14_X_28, u1_u14_X_3, u1_u14_X_33, u1_u14_X_34, u1_u14_X_39, u1_u14_X_4, u1_u14_X_40, u1_u14_X_45, u1_u14_X_46, 
      u1_u14_X_47, u1_u14_X_9, u1_u15_X_1, u1_u15_X_10, u1_u15_X_15, u1_u15_X_16, u1_u15_X_21, u1_u15_X_22, u1_u15_X_23, 
      u1_u15_X_24, u1_u15_X_25, u1_u15_X_26, u1_u15_X_27, u1_u15_X_28, u1_u15_X_3, u1_u15_X_33, u1_u15_X_36, u1_u15_X_38, 
      u1_u15_X_39, u1_u15_X_4, u1_u15_X_40, u1_u15_X_45, u1_u15_X_46, u1_u15_X_47, u1_u15_X_5, u1_u15_X_7, u1_u15_X_9, 
      u1_u1_X_15, u1_u1_X_16, u1_u1_X_21, u1_u1_X_22, u1_u1_X_27, u1_u1_X_28, u1_u1_X_3, u1_u1_X_33, u1_u1_X_34, 
      u1_u1_X_35, u1_u1_X_36, u1_u1_X_37, u1_u1_X_38, u1_u1_X_39, u1_u1_X_4, u1_u1_X_40, u1_u1_X_45, u1_u1_X_46, 
      u1_u1_X_9, u1_u2_X_10, u1_u2_X_11, u1_u2_X_13, u1_u2_X_15, u1_u2_X_16, u1_u2_X_21, u1_u2_X_22, u1_u2_X_27, 
      u1_u2_X_28, u1_u2_X_3, u1_u2_X_30, u1_u2_X_32, u1_u2_X_33, u1_u2_X_34, u1_u2_X_39, u1_u2_X_4, u1_u2_X_40, 
      u1_u2_X_45, u1_u2_X_46, u1_u2_X_9, u1_u3_X_15, u1_u3_X_16, u1_u3_X_21, u1_u3_X_22, u1_u3_X_27, u1_u3_X_28, 
      u1_u3_X_33, u1_u3_X_34, u1_u3_X_39, u1_u3_X_4, u1_u3_X_40, u1_u3_X_45, u1_u3_X_46, u1_u3_X_5, u1_u3_X_7, 
      u1_u3_X_9, u1_u4_X_10, u1_u4_X_15, u1_u4_X_16, u1_u4_X_21, u1_u4_X_28, u1_u4_X_3, u1_u4_X_33, u1_u4_X_34, 
      u1_u4_X_39, u1_u4_X_4, u1_u4_X_40, u1_u4_X_45, u1_u4_X_46, u1_u4_X_9, u1_u5_X_15, u1_u5_X_16, u1_u5_X_17, 
      u1_u5_X_19, u1_u5_X_22, u1_u5_X_27, u1_u5_X_28, u1_u5_X_3, u1_u5_X_33, u1_u5_X_34, u1_u5_X_39, u1_u5_X_40, 
      u1_u5_X_45, u1_u5_X_46, u1_u6_X_10, u1_u6_X_15, u1_u6_X_16, u1_u6_X_21, u1_u6_X_22, u1_u6_X_28, u1_u6_X_3, 
      u1_u6_X_33, u1_u6_X_39, u1_u6_X_4, u1_u6_X_40, u1_u6_X_45, u1_u6_X_9, u1_u7_X_10, u1_u7_X_16, u1_u7_X_17, 
      u1_u7_X_19, u1_u7_X_21, u1_u7_X_22, u1_u7_X_27, u1_u7_X_28, u1_u7_X_33, u1_u7_X_34, u1_u7_X_39, u1_u7_X_4, 
      u1_u7_X_40, u1_u7_X_45, u1_u7_X_46, u1_u7_X_6, u1_u7_X_8, u1_u7_X_9, u1_u8_X_15, u1_u8_X_16, u1_u8_X_21, 
      u1_u8_X_28, u1_u8_X_3, u1_u8_X_30, u1_u8_X_32, u1_u8_X_33, u1_u8_X_34, u1_u8_X_39, u1_u8_X_4, u1_u8_X_40, 
      u1_u8_X_45, u1_u8_X_46, u1_u9_X_10, u1_u9_X_15, u1_u9_X_16, u1_u9_X_17, u1_u9_X_19, u1_u9_X_21, u1_u9_X_27, 
      u1_u9_X_28, u1_u9_X_3, u1_u9_X_34, u1_u9_X_39, u1_u9_X_4, u1_u9_X_40, u1_u9_X_45, u1_u9_X_46, u1_uk_n1002, 
      u1_uk_n1003, u1_uk_n1015, u1_uk_n1021, u1_uk_n1023, u1_uk_n1025, u1_uk_n1029, u1_uk_n1031, u1_uk_n1034, u1_uk_n1038, 
      u1_uk_n1050, u1_uk_n1054, u1_uk_n1056, u1_uk_n1057, u1_uk_n1058, u1_uk_n1060, u1_uk_n1061, u1_uk_n1063, u1_uk_n1065, 
      u1_uk_n1070, u1_uk_n1073, u1_uk_n1074, u1_uk_n1076, u1_uk_n1079, u1_uk_n1080, u1_uk_n1083, u1_uk_n1088, u1_uk_n1090, 
      u1_uk_n1092, u1_uk_n1096, u1_uk_n1101, u1_uk_n1104, u1_uk_n1105, u1_uk_n1106, u1_uk_n1109, u1_uk_n1113, u1_uk_n1114, 
      u1_uk_n1115, u1_uk_n1118, u1_uk_n1119, u1_uk_n1121, u1_uk_n1123, u1_uk_n1124, u1_uk_n1125, u1_uk_n1126, u1_uk_n1128, 
      u1_uk_n1130, u1_uk_n1134, u1_uk_n1138, u1_uk_n1140, u1_uk_n1143, u1_uk_n1147, u1_uk_n1148, u1_uk_n1153, u1_uk_n1154, 
      u1_uk_n1155, u1_uk_n1156, u1_uk_n1157, u1_uk_n1158, u1_uk_n1159, u1_uk_n1160, u1_uk_n1163, u1_uk_n1166, u1_uk_n1167, 
      u1_uk_n1170, u1_uk_n1171, u1_uk_n299, u1_uk_n312, u1_uk_n349, u1_uk_n353, u1_uk_n366, u1_uk_n369, u1_uk_n376, 
      u1_uk_n379, u1_uk_n382, u1_uk_n385, u1_uk_n386, u1_uk_n407, u1_uk_n421, u1_uk_n437, u1_uk_n443, u1_uk_n454, 
      u1_uk_n496, u1_uk_n504, u1_uk_n509, u1_uk_n515, u1_uk_n520, u1_uk_n524, u1_uk_n605, u1_uk_n608, u1_uk_n672, 
      u1_uk_n676, u1_uk_n677, u1_uk_n678, u1_uk_n685, u1_uk_n702, u1_uk_n948, u1_uk_n949, u1_uk_n950, u1_uk_n955, 
      u1_uk_n969, u1_uk_n970, u1_uk_n973, u1_uk_n974, u1_uk_n976, u1_uk_n985, u1_uk_n988, u1_uk_n989, u1_uk_n993, 
      u2_FP_33, u2_FP_36, u2_FP_37, u2_FP_40, u2_FP_41, u2_FP_44, u2_FP_45, u2_FP_48, u2_FP_49, 
      u2_FP_52, u2_FP_53, u2_FP_55, u2_FP_56, u2_FP_57, u2_FP_60, u2_FP_61, u2_FP_64, u2_K10_1, 
      u2_K10_11, u2_K10_13, u2_K10_14, u2_K10_17, u2_K10_18, u2_K10_19, u2_K10_20, u2_K10_23, u2_K10_24, 
      u2_K10_25, u2_K10_26, u2_K10_36, u2_K10_42, u2_K10_43, u2_K10_44, u2_K10_48, u2_K10_5, u2_K10_7, 
      u2_K10_8, u2_K11_11, u2_K11_13, u2_K11_24, u2_K11_26, u2_K11_29, u2_K12_2, u2_K12_20, u2_K12_25, 
      u2_K12_36, u2_K12_38, u2_K12_47, u2_K12_48, u2_K13_32, u2_K13_35, u2_K13_37, u2_K13_48, u2_K14_38, 
      u2_K15_1, u2_K15_12, u2_K15_17, u2_K15_2, u2_K15_23, u2_K15_29, u2_K15_31, u2_K15_35, u2_K15_44, 
      u2_K16_1, u2_K16_11, u2_K16_12, u2_K16_13, u2_K16_14, u2_K16_17, u2_K16_18, u2_K16_19, u2_K16_2, 
      u2_K16_20, u2_K16_23, u2_K16_24, u2_K16_25, u2_K16_26, u2_K16_30, u2_K16_31, u2_K16_32, u2_K16_35, 
      u2_K16_36, u2_K16_38, u2_K16_41, u2_K16_42, u2_K16_44, u2_K16_47, u2_K16_48, u2_K16_5, u2_K16_6, 
      u2_K16_7, u2_K16_8, u2_K1_43, u2_K2_1, u2_K2_11, u2_K2_12, u2_K2_13, u2_K2_17, u2_K2_18, 
      u2_K2_2, u2_K2_20, u2_K2_23, u2_K2_24, u2_K2_25, u2_K2_26, u2_K2_29, u2_K2_30, u2_K2_31, 
      u2_K2_35, u2_K2_36, u2_K2_37, u2_K2_38, u2_K2_42, u2_K2_44, u2_K2_47, u2_K2_48, u2_K2_5, 
      u2_K2_6, u2_K2_8, u2_K3_13, u2_K3_19, u2_K3_20, u2_K3_23, u2_K3_26, u2_K3_42, u2_K3_43, 
      u2_K3_47, u2_K3_48, u2_K4_14, u2_K4_18, u2_K4_19, u2_K4_24, u2_K4_48, u2_K4_6, u2_K4_7, 
      u2_K5_11, u2_K5_13, u2_K5_14, u2_K5_17, u2_K5_18, u2_K5_19, u2_K5_2, u2_K5_23, u2_K5_24, 
      u2_K5_25, u2_K5_26, u2_K5_29, u2_K5_30, u2_K5_31, u2_K5_32, u2_K5_37, u2_K5_38, u2_K5_41, 
      u2_K5_44, u2_K5_48, u2_K5_5, u2_K5_6, u2_K5_8, u2_K6_1, u2_K6_11, u2_K6_13, u2_K6_14, 
      u2_K6_19, u2_K6_20, u2_K6_24, u2_K6_32, u2_K6_47, u2_K6_6, u2_K6_8, u2_K7_26, u2_K7_30, 
      u2_K7_31, u2_K7_35, u2_K7_37, u2_K7_38, u2_K7_43, u2_K7_48, u2_K7_5, u2_K7_7, u2_K8_1, 
      u2_K8_11, u2_K8_13, u2_K8_14, u2_K8_17, u2_K8_18, u2_K8_19, u2_K8_2, u2_K8_20, u2_K8_47, 
      u2_K8_48, u2_K8_5, u2_K8_6, u2_K8_7, u2_K8_8, u2_K9_12, u2_K9_14, u2_K9_23, u2_K9_25, 
      u2_K9_36, u2_K9_37, u2_K9_38, u2_K9_43, u2_K9_5, u2_R0_1, u2_R0_12, u2_R0_13, u2_R0_16, 
      u2_R0_17, u2_R0_19, u2_R0_20, u2_R0_21, u2_R0_24, u2_R0_25, u2_R0_29, u2_R0_32, u2_R0_4, 
      u2_R0_5, u2_R0_7, u2_R0_8, u2_R0_9, u2_R10_1, u2_R10_12, u2_R10_13, u2_R10_16, u2_R10_21, 
      u2_R10_25, u2_R10_29, u2_R10_3, u2_R10_32, u2_R10_4, u2_R10_7, u2_R10_8, u2_R10_9, u2_R11_1, 
      u2_R11_21, u2_R11_24, u2_R11_4, u2_R12_20, u2_R12_21, u2_R12_22, u2_R12_25, u2_R13_1, u2_R13_12, 
      u2_R13_16, u2_R13_17, u2_R13_20, u2_R13_22, u2_R13_24, u2_R13_25, u2_R13_27, u2_R13_29, u2_R13_32, 
      u2_R13_5, u2_R13_9, u2_R1_1, u2_R1_12, u2_R1_13, u2_R1_14, u2_R1_15, u2_R1_16, u2_R1_17, 
      u2_R1_2, u2_R1_25, u2_R1_27, u2_R1_28, u2_R1_29, u2_R1_3, u2_R1_30, u2_R1_31, u2_R1_32, 
      u2_R1_5, u2_R1_6, u2_R1_7, u2_R1_8, u2_R1_9, u2_R2_1, u2_R2_10, u2_R2_11, u2_R2_12, 
      u2_R2_13, u2_R2_16, u2_R2_17, u2_R2_19, u2_R2_2, u2_R2_20, u2_R2_21, u2_R2_25, u2_R2_3, 
      u2_R2_32, u2_R2_4, u2_R2_5, u2_R2_6, u2_R2_7, u2_R2_8, u2_R2_9, u2_R3_1, u2_R3_12, 
      u2_R3_13, u2_R3_16, u2_R3_17, u2_R3_18, u2_R3_20, u2_R3_21, u2_R3_22, u2_R3_24, u2_R3_25, 
      u2_R3_28, u2_R3_29, u2_R3_30, u2_R3_4, u2_R3_5, u2_R3_8, u2_R3_9, u2_R4_1, u2_R4_12, 
      u2_R4_13, u2_R4_14, u2_R4_17, u2_R4_21, u2_R4_22, u2_R4_24, u2_R4_28, u2_R4_29, u2_R4_31, 
      u2_R4_32, u2_R4_4, u2_R4_5, u2_R4_6, u2_R4_8, u2_R4_9, u2_R5_1, u2_R5_10, u2_R5_11, 
      u2_R5_12, u2_R5_13, u2_R5_14, u2_R5_16, u2_R5_17, u2_R5_20, u2_R5_21, u2_R5_23, u2_R5_24, 
      u2_R5_25, u2_R5_26, u2_R5_28, u2_R5_29, u2_R5_32, u2_R5_4, u2_R5_5, u2_R5_8, u2_R5_9, 
      u2_R6_1, u2_R6_12, u2_R6_13, u2_R6_2, u2_R6_28, u2_R6_32, u2_R6_4, u2_R6_5, u2_R6_8, 
      u2_R6_9, u2_R7_1, u2_R7_11, u2_R7_12, u2_R7_13, u2_R7_14, u2_R7_15, u2_R7_16, u2_R7_17, 
      u2_R7_22, u2_R7_24, u2_R7_25, u2_R7_28, u2_R7_29, u2_R7_3, u2_R7_4, u2_R7_5, u2_R7_6, 
      u2_R7_7, u2_R7_8, u2_R7_9, u2_R8_1, u2_R8_12, u2_R8_13, u2_R8_15, u2_R8_16, u2_R8_17, 
      u2_R8_20, u2_R8_22, u2_R8_24, u2_R8_25, u2_R8_26, u2_R8_27, u2_R8_28, u2_R8_29, u2_R8_32, 
      u2_R8_4, u2_R8_5, u2_R8_6, u2_R8_8, u2_R8_9, u2_R9_12, u2_R9_13, u2_R9_17, u2_R9_20, 
      u2_R9_32, u2_R9_8, u2_R9_9, u2_desIn_r_1, u2_desIn_r_25, u2_desIn_r_27, u2_desIn_r_33, u2_desIn_r_57, u2_key_r_14, 
      u2_key_r_23, u2_key_r_30, u2_key_r_7, u2_u0_X_10, u2_u0_X_11, u2_u0_X_12, u2_u0_X_25, u2_u0_X_26, u2_u0_X_27, 
      u2_u0_X_28, u2_u0_X_30, u2_u0_X_32, u2_u0_X_33, u2_u0_X_34, u2_u0_X_35, u2_u0_X_37, u2_u0_X_39, u2_u0_X_40, 
      u2_u0_X_45, u2_u0_X_46, u2_u0_X_48, u2_u0_X_7, u2_u0_X_8, u2_u0_X_9, u2_u10_X_10, u2_u10_X_15, u2_u10_X_16, 
      u2_u10_X_18, u2_u10_X_21, u2_u10_X_22, u2_u10_X_23, u2_u10_X_25, u2_u10_X_27, u2_u10_X_28, u2_u10_X_30, u2_u10_X_32, 
      u2_u10_X_33, u2_u10_X_34, u2_u10_X_35, u2_u10_X_36, u2_u10_X_37, u2_u10_X_38, u2_u10_X_39, u2_u10_X_40, u2_u10_X_41, 
      u2_u10_X_42, u2_u10_X_43, u2_u10_X_44, u2_u10_X_45, u2_u10_X_46, u2_u10_X_48, u2_u10_X_7, u2_u10_X_8, u2_u10_X_9, 
      u2_u11_X_15, u2_u11_X_16, u2_u11_X_21, u2_u11_X_22, u2_u11_X_24, u2_u11_X_26, u2_u11_X_27, u2_u11_X_28, u2_u11_X_29, 
      u2_u11_X_3, u2_u11_X_31, u2_u11_X_33, u2_u11_X_34, u2_u11_X_35, u2_u11_X_37, u2_u11_X_39, u2_u11_X_40, u2_u11_X_41, 
      u2_u11_X_43, u2_u11_X_45, u2_u11_X_46, u2_u11_X_6, u2_u11_X_8, u2_u11_X_9, u2_u12_X_1, u2_u12_X_10, u2_u12_X_11, 
      u2_u12_X_12, u2_u12_X_25, u2_u12_X_26, u2_u12_X_27, u2_u12_X_28, u2_u12_X_29, u2_u12_X_3, u2_u12_X_31, u2_u12_X_33, 
      u2_u12_X_34, u2_u12_X_36, u2_u12_X_38, u2_u12_X_39, u2_u12_X_4, u2_u12_X_40, u2_u12_X_41, u2_u12_X_42, u2_u12_X_43, 
      u2_u12_X_44, u2_u12_X_45, u2_u12_X_46, u2_u12_X_47, u2_u12_X_6, u2_u12_X_8, u2_u12_X_9, u2_u13_X_25, u2_u13_X_26, 
      u2_u13_X_27, u2_u13_X_28, u2_u13_X_34, u2_u13_X_35, u2_u13_X_37, u2_u13_X_39, u2_u13_X_40, u2_u13_X_41, u2_u13_X_42, 
      u2_u13_X_43, u2_u13_X_44, u2_u13_X_45, u2_u13_X_46, u2_u13_X_47, u2_u13_X_48, u2_u14_X_10, u2_u14_X_11, u2_u14_X_13, 
      u2_u14_X_15, u2_u14_X_16, u2_u14_X_18, u2_u14_X_20, u2_u14_X_21, u2_u14_X_22, u2_u14_X_27, u2_u14_X_28, u2_u14_X_3, 
      u2_u14_X_30, u2_u14_X_32, u2_u14_X_34, u2_u14_X_39, u2_u14_X_4, u2_u14_X_41, u2_u14_X_43, u2_u14_X_45, u2_u14_X_46, 
      u2_u14_X_5, u2_u14_X_7, u2_u14_X_9, u2_u15_X_10, u2_u15_X_15, u2_u15_X_16, u2_u15_X_21, u2_u15_X_22, u2_u15_X_27, 
      u2_u15_X_28, u2_u15_X_3, u2_u15_X_33, u2_u15_X_39, u2_u15_X_4, u2_u15_X_40, u2_u15_X_45, u2_u15_X_46, u2_u15_X_9, 
      u2_u1_X_15, u2_u1_X_16, u2_u1_X_21, u2_u1_X_22, u2_u1_X_27, u2_u1_X_3, u2_u1_X_33, u2_u1_X_34, u2_u1_X_39, 
      u2_u1_X_4, u2_u1_X_40, u2_u1_X_41, u2_u1_X_43, u2_u1_X_45, u2_u1_X_46, u2_u1_X_9, u2_u2_X_15, u2_u2_X_16, 
      u2_u2_X_27, u2_u2_X_28, u2_u2_X_29, u2_u2_X_30, u2_u2_X_31, u2_u2_X_32, u2_u2_X_33, u2_u2_X_34, u2_u2_X_35, 
      u2_u2_X_37, u2_u2_X_39, u2_u2_X_5, u2_u2_X_7, u2_u3_X_21, u2_u3_X_22, u2_u3_X_27, u2_u3_X_33, u2_u3_X_34, 
      u2_u3_X_35, u2_u3_X_43, u2_u3_X_44, u2_u3_X_45, u2_u3_X_46, u2_u4_X_1, u2_u4_X_10, u2_u4_X_15, u2_u4_X_16, 
      u2_u4_X_21, u2_u4_X_22, u2_u4_X_28, u2_u4_X_3, u2_u4_X_34, u2_u4_X_39, u2_u4_X_4, u2_u4_X_40, u2_u4_X_46, 
      u2_u4_X_47, u2_u4_X_9, u2_u5_X_10, u2_u5_X_15, u2_u5_X_16, u2_u5_X_22, u2_u5_X_23, u2_u5_X_25, u2_u5_X_27, 
      u2_u5_X_28, u2_u5_X_29, u2_u5_X_3, u2_u5_X_31, u2_u5_X_34, u2_u5_X_36, u2_u5_X_38, u2_u5_X_39, u2_u5_X_4, 
      u2_u5_X_40, u2_u5_X_45, u2_u6_X_10, u2_u6_X_22, u2_u6_X_27, u2_u6_X_28, u2_u6_X_3, u2_u6_X_33, u2_u6_X_4, 
      u2_u6_X_40, u2_u6_X_45, u2_u6_X_46, u2_u6_X_9, u2_u7_X_10, u2_u7_X_15, u2_u7_X_16, u2_u7_X_21, u2_u7_X_22, 
      u2_u7_X_23, u2_u7_X_24, u2_u7_X_4, u2_u7_X_44, u2_u7_X_45, u2_u7_X_46, u2_u7_X_9, u2_u8_X_1, u2_u8_X_15, 
      u2_u8_X_27, u2_u8_X_28, u2_u8_X_29, u2_u8_X_3, u2_u8_X_30, u2_u8_X_31, u2_u8_X_32, u2_u8_X_34, u2_u8_X_39, 
      u2_u8_X_40, u2_u8_X_45, u2_u8_X_46, u2_u8_X_47, u2_u9_X_10, u2_u9_X_15, u2_u9_X_16, u2_u9_X_21, u2_u9_X_27, 
      u2_u9_X_28, u2_u9_X_29, u2_u9_X_3, u2_u9_X_30, u2_u9_X_32, u2_u9_X_34, u2_u9_X_4, u2_u9_X_45, u2_u9_X_46, 
      u2_u9_X_6, u2_uk_K_r11_28, u2_uk_K_r11_48, u2_uk_K_r11_53, u2_uk_K_r13_22, u2_uk_K_r13_32, u2_uk_K_r1_15, u2_uk_K_r1_16, u2_uk_K_r1_18, 
      u2_uk_K_r1_21, u2_uk_K_r1_22, u2_uk_K_r1_47, u2_uk_K_r2_13, u2_uk_K_r2_18, u2_uk_K_r2_21, u2_uk_K_r2_25, u2_uk_K_r2_27, u2_uk_K_r2_28, 
      u2_uk_K_r2_31, u2_uk_K_r2_36, u2_uk_K_r2_49, u2_uk_K_r2_55, u2_uk_K_r3_11, u2_uk_K_r3_14, u2_uk_K_r3_19, u2_uk_K_r3_43, u2_uk_K_r3_9, 
      u2_uk_K_r4_11, u2_uk_K_r4_17, u2_uk_K_r4_33, u2_uk_K_r4_35, u2_uk_K_r4_38, u2_uk_K_r4_4, u2_uk_K_r4_5, u2_uk_K_r4_55, u2_uk_K_r5_10, 
      u2_uk_K_r5_17, u2_uk_K_r5_19, u2_uk_K_r5_39, u2_uk_K_r5_4, u2_uk_K_r5_41, u2_uk_K_r7_0, u2_uk_K_r7_25, u2_uk_K_r7_26, u2_uk_K_r7_32, 
      u2_uk_K_r7_39, u2_uk_K_r7_41, u2_uk_K_r7_48, u2_uk_K_r7_55, u2_uk_K_r8_16, u2_uk_K_r8_2, u2_uk_K_r8_22, u2_uk_K_r8_37, u2_uk_K_r8_41, 
      u2_uk_K_r8_42, u2_uk_K_r9_10, u2_uk_K_r9_4, u2_uk_K_r9_48, u2_uk_n1004, u2_uk_n1008, u2_uk_n1020, u2_uk_n1024, u2_uk_n1027, 
      u2_uk_n1028, u2_uk_n1031, u2_uk_n1035, u2_uk_n1038, u2_uk_n1040, u2_uk_n1043, u2_uk_n1046, u2_uk_n1049, u2_uk_n1050, 
      u2_uk_n1053, u2_uk_n1069, u2_uk_n1074, u2_uk_n1076, u2_uk_n1077, u2_uk_n1079, u2_uk_n1082, u2_uk_n1083, u2_uk_n1084, 
      u2_uk_n1088, u2_uk_n1089, u2_uk_n1091, u2_uk_n1093, u2_uk_n1096, u2_uk_n1098, u2_uk_n1110, u2_uk_n1113, u2_uk_n1120, 
      u2_uk_n1123, u2_uk_n1124, u2_uk_n1128, u2_uk_n1130, u2_uk_n1132, u2_uk_n1133, u2_uk_n1136, u2_uk_n1137, u2_uk_n1140, 
      u2_uk_n1141, u2_uk_n1142, u2_uk_n1152, u2_uk_n1171, u2_uk_n1279, u2_uk_n1280, u2_uk_n1281, u2_uk_n1282, u2_uk_n1283, 
      u2_uk_n1284, u2_uk_n1285, u2_uk_n1286, u2_uk_n1287, u2_uk_n1288, u2_uk_n1290, u2_uk_n1291, u2_uk_n1293, u2_uk_n1295, 
      u2_uk_n1296, u2_uk_n1297, u2_uk_n1300, u2_uk_n1301, u2_uk_n1302, u2_uk_n1305, u2_uk_n1306, u2_uk_n1310, u2_uk_n1311, 
      u2_uk_n1314, u2_uk_n1316, u2_uk_n1317, u2_uk_n1318, u2_uk_n1323, u2_uk_n1324, u2_uk_n1326, u2_uk_n1328, u2_uk_n1329, 
      u2_uk_n1333, u2_uk_n1339, u2_uk_n1341, u2_uk_n1345, u2_uk_n1346, u2_uk_n1350, u2_uk_n1351, u2_uk_n1356, u2_uk_n1359, 
      u2_uk_n1361, u2_uk_n1370, u2_uk_n1375, u2_uk_n1382, u2_uk_n1401, u2_uk_n1405, u2_uk_n1408, u2_uk_n1410, u2_uk_n1413, 
      u2_uk_n1422, u2_uk_n1426, u2_uk_n1428, u2_uk_n1433, u2_uk_n1435, u2_uk_n1438, u2_uk_n1439, u2_uk_n1440, u2_uk_n1441, 
      u2_uk_n1445, u2_uk_n1446, u2_uk_n1447, u2_uk_n1453, u2_uk_n1454, u2_uk_n1456, u2_uk_n1458, u2_uk_n1459, u2_uk_n1462, 
      u2_uk_n1465, u2_uk_n1466, u2_uk_n1470, u2_uk_n1475, u2_uk_n1480, u2_uk_n1486, u2_uk_n1488, u2_uk_n1490, u2_uk_n1493, 
      u2_uk_n1494, u2_uk_n1496, u2_uk_n1497, u2_uk_n1544, u2_uk_n1548, u2_uk_n1549, u2_uk_n1555, u2_uk_n1556, u2_uk_n1563, 
      u2_uk_n1568, u2_uk_n1573, u2_uk_n1580, u2_uk_n1585, u2_uk_n1586, u2_uk_n1592, u2_uk_n1594, u2_uk_n1609, u2_uk_n1615, 
      u2_uk_n1622, u2_uk_n1682, u2_uk_n1683, u2_uk_n1688, u2_uk_n1689, u2_uk_n1693, u2_uk_n1708, u2_uk_n1709, u2_uk_n1720, 
      u2_uk_n1721, u2_uk_n1746, u2_uk_n1769, u2_uk_n1770, u2_uk_n1781, u2_uk_n1785, u2_uk_n1797, u2_uk_n1803, u2_uk_n1807, 
      u2_uk_n1808, u2_uk_n1816, u2_uk_n1817, u2_uk_n1819, u2_uk_n1821, u2_uk_n1824, u2_uk_n1826, u2_uk_n1834, u2_uk_n1840, 
      u2_uk_n1846, u2_uk_n1849, u2_uk_n1851, u2_uk_n1852, u2_uk_n1855, u2_uk_n1856, u2_uk_n238, u2_uk_n240, u2_uk_n257, 
      u2_uk_n299, u2_uk_n301, u2_uk_n305, u2_uk_n308, u2_uk_n313, u2_uk_n319, u2_uk_n335, u2_uk_n373, u2_uk_n386, 
      u2_uk_n408, u2_uk_n415, u2_uk_n421, u2_uk_n454, u2_uk_n456, u2_uk_n467, u2_uk_n503, u2_uk_n504, u2_uk_n515, 
      u2_uk_n520, u2_uk_n665, u2_uk_n682, u2_uk_n689, u2_uk_n939, u2_uk_n942, u2_uk_n943, u2_uk_n945, u2_uk_n946, 
      u2_uk_n955, u2_uk_n958, u2_uk_n959, u2_uk_n963, u2_uk_n985, u2_uk_n986, u2_uk_n987, u2_uk_n991, u2_uk_n993, 
      u2_uk_n995, u2_uk_n998, u2_uk_n999 );
  des_des_die_1 u1 ( u0_K10_1, u0_K10_14, u0_K10_17, u0_K10_18, u0_K10_19, u0_K10_20, u0_K10_32, u0_K14_23, u0_K14_24, 
      u0_K14_25, u0_K14_26, u0_K14_29, u0_K14_5, u0_K14_7, u0_K4_36, u0_K4_43, u0_K4_48, u0_K4_6, 
      u0_K5_1, u0_K5_18, u0_K5_24, u0_K5_26, u0_K5_29, u0_K5_31, u0_K5_47, u0_K5_8, u0_K8_11, 
      u0_K8_13, u0_K8_19, u0_R11_16, u0_R11_20, u0_R12_16, u0_R12_17, u0_R12_19, u0_R12_20, u0_R12_22, 
      u0_R12_23, u0_R12_24, u0_R12_4, u0_R13_17, u0_R13_18, u0_R13_19, u0_R13_20, u0_R13_21, u0_R13_22, 
      u0_R13_23, u0_R13_24, u0_R13_25, u0_R13_26, u0_R13_27, u0_R13_28, u0_R13_29, u0_R13_30, u0_R13_31, 
      u0_R2_1, u0_R2_10, u0_R2_11, u0_R2_12, u0_R2_13, u0_R2_14, u0_R2_16, u0_R2_2, u0_R2_21, 
      u0_R2_22, u0_R2_25, u0_R2_28, u0_R2_3, u0_R2_32, u0_R2_4, u0_R2_5, u0_R2_6, u0_R2_7, 
      u0_R2_8, u0_R2_9, u0_R3_13, u0_R3_15, u0_R3_17, u0_R3_18, u0_R3_20, u0_R3_22, u0_R3_24, 
      u0_R3_25, u0_R3_32, u0_R3_5, u0_R5_12, u0_R5_13, u0_R5_2, u0_R5_25, u0_R5_3, u0_R5_32, 
      u0_R5_4, u0_R5_5, u0_R5_7, u0_R5_8, u0_R5_9, u0_R6_10, u0_R6_11, u0_R6_12, u0_R6_13, 
      u0_R6_14, u0_R6_17, u0_R6_4, u0_R6_5, u0_R6_7, u0_R6_8, u0_R6_9, u0_R8_1, u0_R8_12, 
      u0_R8_13, u0_R8_17, u0_R8_19, u0_R8_20, u0_R8_21, u0_R8_22, u0_R8_27, u0_R8_29, u0_R8_30, 
      u0_R8_32, u0_R8_5, u0_R8_6, u0_R8_9, u0_u12_X_26, u0_u12_X_27, u0_u12_X_28, u0_u12_X_30, u0_u12_X_32, 
      u0_u12_X_33, u0_u12_X_34, u0_u12_X_35, u0_u12_X_36, u0_u13_X_1, u0_u13_X_10, u0_u13_X_11, u0_u13_X_12, u0_u13_X_19, 
      u0_u13_X_2, u0_u13_X_20, u0_u13_X_21, u0_u13_X_22, u0_u13_X_27, u0_u13_X_3, u0_u13_X_30, u0_u13_X_32, u0_u13_X_36, 
      u0_u13_X_38, u0_u13_X_39, u0_u13_X_4, u0_u13_X_40, u0_u13_X_41, u0_u13_X_42, u0_u13_X_6, u0_u13_X_8, u0_u13_X_9, 
      u0_u14_X_25, u0_u14_X_47, u0_u14_X_48, u0_u3_X_22, u0_u3_X_24, u0_u3_X_26, u0_u3_X_27, u0_u3_X_28, u0_u3_X_29, 
      u0_u3_X_31, u0_u3_X_34, u0_u3_X_35, u0_u3_X_37, u0_u3_X_39, u0_u3_X_40, u0_u3_X_42, u0_u3_X_44, u0_u3_X_45, 
      u0_u3_X_46, u0_u4_X_10, u0_u4_X_11, u0_u4_X_12, u0_u4_X_13, u0_u4_X_14, u0_u4_X_15, u0_u4_X_16, u0_u4_X_17, 
      u0_u4_X_19, u0_u4_X_2, u0_u4_X_21, u0_u4_X_23, u0_u4_X_25, u0_u4_X_28, u0_u4_X_3, u0_u4_X_30, u0_u4_X_32, 
      u0_u4_X_34, u0_u4_X_4, u0_u4_X_43, u0_u4_X_44, u0_u4_X_45, u0_u4_X_46, u0_u4_X_48, u0_u4_X_5, u0_u4_X_7, 
      u0_u4_X_9, u0_u6_X_15, u0_u6_X_16, u0_u6_X_2, u0_u6_X_21, u0_u6_X_22, u0_u6_X_23, u0_u6_X_24, u0_u6_X_31, 
      u0_u6_X_32, u0_u6_X_33, u0_u6_X_34, u0_u6_X_35, u0_u6_X_9, u0_u7_X_1, u0_u7_X_2, u0_u7_X_22, u0_u7_X_23, 
      u0_u7_X_3, u0_u7_X_4, u0_u7_X_9, u0_u9_X_10, u0_u9_X_11, u0_u9_X_13, u0_u9_X_15, u0_u9_X_16, u0_u9_X_21, 
      u0_u9_X_22, u0_u9_X_23, u0_u9_X_25, u0_u9_X_27, u0_u9_X_3, u0_u9_X_34, u0_u9_X_35, u0_u9_X_36, u0_u9_X_37, 
      u0_u9_X_38, u0_u9_X_39, u0_u9_X_4, u0_u9_X_41, u0_u9_X_43, u0_u9_X_46, u0_u9_X_5, u0_u9_X_7, u0_uk_K_r13_0, 
      u0_uk_K_r13_38, u0_uk_K_r13_44, u0_uk_K_r2_13, u0_uk_K_r2_18, u0_uk_K_r2_20, u0_uk_K_r2_25, u0_uk_K_r2_26, u0_uk_K_r2_27, u0_uk_K_r2_28, 
      u0_uk_K_r2_33, u0_uk_K_r2_4, u0_uk_K_r2_41, u0_uk_K_r2_46, u0_uk_K_r2_50, u0_uk_K_r2_53, u0_uk_K_r2_55, u0_uk_K_r3_10, u0_uk_K_r3_14, 
      u0_uk_K_r5_10, u0_uk_K_r5_17, u0_uk_K_r5_39, u0_uk_K_r5_4, u0_uk_K_r6_26, u0_uk_K_r6_34, u0_uk_K_r6_46, u0_uk_K_r8_16, u0_uk_K_r8_40, 
      u0_uk_K_r8_41, u0_uk_n10, u0_uk_n100, u0_uk_n1005, u0_uk_n1006, u0_uk_n1012, u0_uk_n102, u0_uk_n1024, u0_uk_n109, 
      u0_uk_n11, u0_uk_n110, u0_uk_n113, u0_uk_n116, u0_uk_n117, u0_uk_n118, u0_uk_n12, u0_uk_n123, u0_uk_n128, 
      u0_uk_n129, u0_uk_n13, u0_uk_n141, u0_uk_n142, u0_uk_n145, u0_uk_n146, u0_uk_n147, u0_uk_n148, u0_uk_n155, 
      u0_uk_n161, u0_uk_n162, u0_uk_n163, u0_uk_n164, u0_uk_n17, u0_uk_n18, u0_uk_n182, u0_uk_n187, u0_uk_n188, 
      u0_uk_n202, u0_uk_n203, u0_uk_n207, u0_uk_n208, u0_uk_n209, u0_uk_n21, u0_uk_n214, u0_uk_n217, u0_uk_n22, 
      u0_uk_n220, u0_uk_n23, u0_uk_n230, u0_uk_n231, u0_uk_n232, u0_uk_n233, u0_uk_n238, u0_uk_n239, u0_uk_n240, 
      u0_uk_n241, u0_uk_n242, u0_uk_n243, u0_uk_n244, u0_uk_n248, u0_uk_n249, u0_uk_n250, u0_uk_n251, u0_uk_n252, 
      u0_uk_n253, u0_uk_n257, u0_uk_n259, u0_uk_n260, u0_uk_n261, u0_uk_n264, u0_uk_n266, u0_uk_n267, u0_uk_n269, 
      u0_uk_n27, u0_uk_n28, u0_uk_n3, u0_uk_n31, u0_uk_n318, u0_uk_n32, u0_uk_n324, u0_uk_n329, u0_uk_n33, 
      u0_uk_n330, u0_uk_n331, u0_uk_n336, u0_uk_n337, u0_uk_n339, u0_uk_n344, u0_uk_n352, u0_uk_n358, u0_uk_n361, 
      u0_uk_n370, u0_uk_n371, u0_uk_n383, u0_uk_n384, u0_uk_n39, u0_uk_n392, u0_uk_n393, u0_uk_n396, u0_uk_n4, 
      u0_uk_n40, u0_uk_n400, u0_uk_n401, u0_uk_n405, u0_uk_n41, u0_uk_n45, u0_uk_n457, u0_uk_n471, u0_uk_n497, 
      u0_uk_n499, u0_uk_n5, u0_uk_n502, u0_uk_n505, u0_uk_n508, u0_uk_n510, u0_uk_n511, u0_uk_n513, u0_uk_n517, 
      u0_uk_n519, u0_uk_n522, u0_uk_n523, u0_uk_n525, u0_uk_n529, u0_uk_n530, u0_uk_n531, u0_uk_n532, u0_uk_n534, 
      u0_uk_n535, u0_uk_n536, u0_uk_n539, u0_uk_n55, u0_uk_n60, u0_uk_n61, u0_uk_n63, u0_uk_n67, u0_uk_n73, 
      u0_uk_n759, u0_uk_n761, u0_uk_n763, u0_uk_n768, u0_uk_n780, u0_uk_n783, u0_uk_n809, u0_uk_n810, u0_uk_n813, 
      u0_uk_n815, u0_uk_n816, u0_uk_n83, u0_uk_n832, u0_uk_n839, u0_uk_n9, u0_uk_n915, u0_uk_n916, u0_uk_n917, 
      u0_uk_n918, u0_uk_n92, u0_uk_n93, u0_uk_n933, u0_uk_n934, u0_uk_n94, u0_uk_n98, u0_uk_n99, u2_K10_1, 
      u2_K10_36, u2_K10_42, u2_K10_43, u2_K10_44, u2_K10_48, u2_K10_5, u2_K11_24, u2_K11_26, u2_K11_29, 
      u2_K12_2, u2_K12_20, u2_K12_25, u2_K12_36, u2_K12_38, u2_K12_47, u2_K12_48, u2_K13_32, u2_K13_35, 
      u2_K13_37, u2_K13_48, u2_K14_38, u2_K15_1, u2_K15_12, u2_K15_17, u2_K15_2, u2_K15_23, u2_K15_29, 
      u2_K15_31, u2_K15_35, u2_K15_44, u2_K1_43, u2_K3_13, u2_K3_19, u2_K3_20, u2_K3_23, u2_K3_26, 
      u2_K3_42, u2_K3_43, u2_K3_47, u2_K3_48, u2_K4_14, u2_K4_18, u2_K4_19, u2_K4_24, u2_K4_48, 
      u2_K4_6, u2_K4_7, u2_K5_11, u2_K5_13, u2_K5_14, u2_K5_17, u2_K5_18, u2_K5_19, u2_K5_2, 
      u2_K5_23, u2_K5_24, u2_K5_25, u2_K5_26, u2_K5_29, u2_K5_30, u2_K5_31, u2_K5_32, u2_K5_37, 
      u2_K5_38, u2_K5_41, u2_K5_44, u2_K5_48, u2_K5_5, u2_K5_6, u2_K5_8, u2_K6_1, u2_K6_11, 
      u2_K6_13, u2_K6_14, u2_K6_19, u2_K6_20, u2_K6_24, u2_K6_32, u2_K6_47, u2_K6_6, u2_K6_8, 
      u2_K7_26, u2_K7_30, u2_K7_31, u2_K7_35, u2_K7_37, u2_K7_38, u2_K7_43, u2_K7_48, u2_K7_5, 
      u2_K7_7, u2_K9_12, u2_K9_14, u2_K9_23, u2_K9_25, u2_K9_5, u2_R10_1, u2_R10_12, u2_R10_13, 
      u2_R10_16, u2_R10_21, u2_R10_25, u2_R10_29, u2_R10_3, u2_R10_32, u2_R10_4, u2_R10_7, u2_R10_8, 
      u2_R10_9, u2_R11_1, u2_R11_21, u2_R11_24, u2_R11_4, u2_R12_20, u2_R12_21, u2_R12_22, u2_R12_25, 
      u2_R13_1, u2_R13_12, u2_R13_16, u2_R13_17, u2_R13_20, u2_R13_22, u2_R13_24, u2_R13_25, u2_R13_27, 
      u2_R13_29, u2_R13_32, u2_R13_5, u2_R13_9, u2_R1_1, u2_R1_12, u2_R1_13, u2_R1_14, u2_R1_15, 
      u2_R1_16, u2_R1_17, u2_R1_2, u2_R1_25, u2_R1_27, u2_R1_28, u2_R1_29, u2_R1_3, u2_R1_30, 
      u2_R1_31, u2_R1_32, u2_R1_5, u2_R1_6, u2_R1_7, u2_R1_8, u2_R1_9, u2_R2_1, u2_R2_10, 
      u2_R2_11, u2_R2_12, u2_R2_13, u2_R2_16, u2_R2_17, u2_R2_19, u2_R2_2, u2_R2_20, u2_R2_21, 
      u2_R2_25, u2_R2_3, u2_R2_32, u2_R2_4, u2_R2_5, u2_R2_6, u2_R2_7, u2_R2_8, u2_R2_9, 
      u2_R3_1, u2_R3_12, u2_R3_13, u2_R3_16, u2_R3_17, u2_R3_18, u2_R3_20, u2_R3_21, u2_R3_22, 
      u2_R3_24, u2_R3_25, u2_R3_28, u2_R3_29, u2_R3_30, u2_R3_4, u2_R3_5, u2_R3_8, u2_R3_9, 
      u2_R4_1, u2_R4_12, u2_R4_13, u2_R4_14, u2_R4_17, u2_R4_21, u2_R4_22, u2_R4_24, u2_R4_28, 
      u2_R4_29, u2_R4_31, u2_R4_32, u2_R4_4, u2_R4_5, u2_R4_6, u2_R4_8, u2_R4_9, u2_R5_1, 
      u2_R5_10, u2_R5_11, u2_R5_12, u2_R5_13, u2_R5_14, u2_R5_16, u2_R5_17, u2_R5_20, u2_R5_21, 
      u2_R5_23, u2_R5_24, u2_R5_25, u2_R5_26, u2_R5_28, u2_R5_29, u2_R5_32, u2_R5_4, u2_R5_5, 
      u2_R5_8, u2_R5_9, u2_R7_1, u2_R7_11, u2_R7_12, u2_R7_13, u2_R7_14, u2_R7_15, u2_R7_16, 
      u2_R7_17, u2_R7_3, u2_R7_4, u2_R7_5, u2_R7_6, u2_R7_7, u2_R7_8, u2_R7_9, u2_R8_1, 
      u2_R8_20, u2_R8_22, u2_R8_24, u2_R8_25, u2_R8_26, u2_R8_27, u2_R8_28, u2_R8_29, u2_R8_32, 
      u2_R8_4, u2_R9_12, u2_R9_13, u2_R9_17, u2_R9_20, u2_R9_32, u2_desIn_r_1, u2_desIn_r_25, u2_desIn_r_27, 
      u2_desIn_r_33, u2_desIn_r_57, u2_key_r_14, u2_key_r_23, u2_key_r_30, u2_key_r_7, u2_u0_X_10, u2_u0_X_11, u2_u0_X_12, 
      u2_u0_X_25, u2_u0_X_26, u2_u0_X_27, u2_u0_X_28, u2_u0_X_30, u2_u0_X_32, u2_u0_X_33, u2_u0_X_34, u2_u0_X_35, 
      u2_u0_X_37, u2_u0_X_39, u2_u0_X_40, u2_u0_X_45, u2_u0_X_46, u2_u0_X_48, u2_u0_X_7, u2_u0_X_8, u2_u0_X_9, 
      u2_u10_X_21, u2_u10_X_22, u2_u10_X_23, u2_u10_X_25, u2_u10_X_27, u2_u10_X_28, u2_u10_X_30, u2_u10_X_32, u2_u10_X_33, 
      u2_u10_X_34, u2_u10_X_35, u2_u10_X_36, u2_u10_X_37, u2_u10_X_38, u2_u10_X_39, u2_u10_X_40, u2_u10_X_41, u2_u10_X_42, 
      u2_u10_X_43, u2_u10_X_44, u2_u10_X_45, u2_u10_X_46, u2_u10_X_48, u2_u11_X_15, u2_u11_X_16, u2_u11_X_21, u2_u11_X_22, 
      u2_u11_X_24, u2_u11_X_26, u2_u11_X_27, u2_u11_X_28, u2_u11_X_29, u2_u11_X_3, u2_u11_X_31, u2_u11_X_33, u2_u11_X_34, 
      u2_u11_X_35, u2_u11_X_37, u2_u11_X_39, u2_u11_X_40, u2_u11_X_41, u2_u11_X_43, u2_u11_X_45, u2_u11_X_46, u2_u11_X_6, 
      u2_u11_X_8, u2_u11_X_9, u2_u12_X_1, u2_u12_X_10, u2_u12_X_11, u2_u12_X_12, u2_u12_X_25, u2_u12_X_26, u2_u12_X_27, 
      u2_u12_X_28, u2_u12_X_29, u2_u12_X_3, u2_u12_X_31, u2_u12_X_33, u2_u12_X_34, u2_u12_X_36, u2_u12_X_38, u2_u12_X_39, 
      u2_u12_X_4, u2_u12_X_40, u2_u12_X_41, u2_u12_X_42, u2_u12_X_43, u2_u12_X_44, u2_u12_X_45, u2_u12_X_46, u2_u12_X_47, 
      u2_u12_X_6, u2_u12_X_8, u2_u12_X_9, u2_u13_X_25, u2_u13_X_26, u2_u13_X_27, u2_u13_X_28, u2_u13_X_34, u2_u13_X_35, 
      u2_u13_X_37, u2_u13_X_39, u2_u13_X_40, u2_u13_X_41, u2_u13_X_42, u2_u13_X_43, u2_u13_X_44, u2_u13_X_45, u2_u13_X_46, 
      u2_u13_X_47, u2_u13_X_48, u2_u14_X_10, u2_u14_X_11, u2_u14_X_13, u2_u14_X_15, u2_u14_X_16, u2_u14_X_18, u2_u14_X_20, 
      u2_u14_X_21, u2_u14_X_22, u2_u14_X_27, u2_u14_X_28, u2_u14_X_3, u2_u14_X_30, u2_u14_X_32, u2_u14_X_34, u2_u14_X_39, 
      u2_u14_X_4, u2_u14_X_41, u2_u14_X_43, u2_u14_X_45, u2_u14_X_46, u2_u14_X_5, u2_u14_X_7, u2_u14_X_9, u2_u2_X_15, 
      u2_u2_X_16, u2_u2_X_27, u2_u2_X_28, u2_u2_X_29, u2_u2_X_30, u2_u2_X_31, u2_u2_X_32, u2_u2_X_33, u2_u2_X_34, 
      u2_u2_X_35, u2_u2_X_37, u2_u2_X_39, u2_u2_X_5, u2_u2_X_7, u2_u3_X_21, u2_u3_X_22, u2_u3_X_27, u2_u3_X_33, 
      u2_u3_X_34, u2_u3_X_35, u2_u3_X_43, u2_u3_X_44, u2_u3_X_45, u2_u3_X_46, u2_u4_X_1, u2_u4_X_10, u2_u4_X_15, 
      u2_u4_X_16, u2_u4_X_21, u2_u4_X_22, u2_u4_X_28, u2_u4_X_3, u2_u4_X_34, u2_u4_X_39, u2_u4_X_4, u2_u4_X_40, 
      u2_u4_X_46, u2_u4_X_47, u2_u4_X_9, u2_u5_X_10, u2_u5_X_15, u2_u5_X_16, u2_u5_X_22, u2_u5_X_23, u2_u5_X_25, 
      u2_u5_X_27, u2_u5_X_28, u2_u5_X_29, u2_u5_X_3, u2_u5_X_31, u2_u5_X_34, u2_u5_X_36, u2_u5_X_38, u2_u5_X_39, 
      u2_u5_X_4, u2_u5_X_40, u2_u5_X_45, u2_u6_X_10, u2_u6_X_22, u2_u6_X_27, u2_u6_X_28, u2_u6_X_3, u2_u6_X_33, 
      u2_u6_X_4, u2_u6_X_40, u2_u6_X_45, u2_u6_X_46, u2_u6_X_9, u2_u8_X_1, u2_u8_X_15, u2_u8_X_27, u2_u8_X_28, 
      u2_u8_X_29, u2_u8_X_3, u2_u8_X_30, u2_u9_X_3, u2_u9_X_32, u2_u9_X_34, u2_u9_X_4, u2_u9_X_45, u2_u9_X_46, 
      u2_u9_X_6, u2_uk_K_r11_28, u2_uk_K_r11_48, u2_uk_K_r11_53, u2_uk_K_r13_22, u2_uk_K_r13_32, u2_uk_K_r1_15, u2_uk_K_r1_16, u2_uk_K_r1_18, 
      u2_uk_K_r1_21, u2_uk_K_r1_22, u2_uk_K_r1_47, u2_uk_K_r2_13, u2_uk_K_r2_18, u2_uk_K_r2_21, u2_uk_K_r2_25, u2_uk_K_r2_27, u2_uk_K_r2_28, 
      u2_uk_K_r2_31, u2_uk_K_r2_36, u2_uk_K_r2_49, u2_uk_K_r2_55, u2_uk_K_r3_11, u2_uk_K_r3_14, u2_uk_K_r3_19, u2_uk_K_r3_43, u2_uk_K_r3_9, 
      u2_uk_K_r4_11, u2_uk_K_r4_17, u2_uk_K_r4_33, u2_uk_K_r4_35, u2_uk_K_r4_38, u2_uk_K_r4_4, u2_uk_K_r4_5, u2_uk_K_r4_55, u2_uk_K_r5_10, 
      u2_uk_K_r5_17, u2_uk_K_r5_19, u2_uk_K_r5_39, u2_uk_K_r5_4, u2_uk_K_r5_41, u2_uk_K_r7_25, u2_uk_K_r7_26, u2_uk_K_r7_32, u2_uk_K_r7_39, 
      u2_uk_K_r7_41, u2_uk_K_r7_48, u2_uk_K_r7_55, u2_uk_K_r8_16, u2_uk_K_r8_2, u2_uk_K_r8_22, u2_uk_K_r8_37, u2_uk_K_r8_41, u2_uk_K_r8_42, 
      u2_uk_K_r9_10, u2_uk_K_r9_4, u2_uk_K_r9_48, u2_uk_n1008, u2_uk_n1020, u2_uk_n1024, u2_uk_n1027, u2_uk_n1028, u2_uk_n1031, 
      u2_uk_n1035, u2_uk_n1038, u2_uk_n1040, u2_uk_n1043, u2_uk_n1046, u2_uk_n1049, u2_uk_n1050, u2_uk_n1053, u2_uk_n1069, 
      u2_uk_n1074, u2_uk_n1076, u2_uk_n1077, u2_uk_n1079, u2_uk_n1082, u2_uk_n1083, u2_uk_n1084, u2_uk_n1088, u2_uk_n1089, 
      u2_uk_n1091, u2_uk_n1093, u2_uk_n1096, u2_uk_n1120, u2_uk_n1123, u2_uk_n1124, u2_uk_n1128, u2_uk_n1130, u2_uk_n1141, 
      u2_uk_n1142, u2_uk_n1152, u2_uk_n1171, u2_uk_n1279, u2_uk_n1280, u2_uk_n1281, u2_uk_n1282, u2_uk_n1283, u2_uk_n1284, 
      u2_uk_n1285, u2_uk_n1286, u2_uk_n1287, u2_uk_n1288, u2_uk_n1290, u2_uk_n1291, u2_uk_n1293, u2_uk_n1295, u2_uk_n1296, 
      u2_uk_n1297, u2_uk_n1300, u2_uk_n1301, u2_uk_n1302, u2_uk_n1305, u2_uk_n1306, u2_uk_n1310, u2_uk_n1311, u2_uk_n1314, 
      u2_uk_n1316, u2_uk_n1317, u2_uk_n1318, u2_uk_n1323, u2_uk_n1324, u2_uk_n1326, u2_uk_n1328, u2_uk_n1329, u2_uk_n1333, 
      u2_uk_n1339, u2_uk_n1341, u2_uk_n1345, u2_uk_n1346, u2_uk_n1350, u2_uk_n1351, u2_uk_n1356, u2_uk_n1359, u2_uk_n1361, 
      u2_uk_n1370, u2_uk_n1375, u2_uk_n1382, u2_uk_n1401, u2_uk_n1405, u2_uk_n1408, u2_uk_n1410, u2_uk_n1413, u2_uk_n1422, 
      u2_uk_n1426, u2_uk_n1428, u2_uk_n1433, u2_uk_n1435, u2_uk_n1438, u2_uk_n1439, u2_uk_n1440, u2_uk_n1441, u2_uk_n1445, 
      u2_uk_n1446, u2_uk_n1447, u2_uk_n1453, u2_uk_n1454, u2_uk_n1456, u2_uk_n1458, u2_uk_n1459, u2_uk_n1462, u2_uk_n1465, 
      u2_uk_n1466, u2_uk_n1470, u2_uk_n1475, u2_uk_n1480, u2_uk_n1486, u2_uk_n1488, u2_uk_n1490, u2_uk_n1493, u2_uk_n1494, 
      u2_uk_n1496, u2_uk_n1497, u2_uk_n1544, u2_uk_n1548, u2_uk_n1549, u2_uk_n1555, u2_uk_n1556, u2_uk_n1563, u2_uk_n1568, 
      u2_uk_n1573, u2_uk_n1580, u2_uk_n1586, u2_uk_n1592, u2_uk_n1594, u2_uk_n1609, u2_uk_n1615, u2_uk_n1622, u2_uk_n1682, 
      u2_uk_n1683, u2_uk_n1688, u2_uk_n1689, u2_uk_n1693, u2_uk_n1708, u2_uk_n1709, u2_uk_n1720, u2_uk_n1721, u2_uk_n1746, 
      u2_uk_n1769, u2_uk_n1770, u2_uk_n1781, u2_uk_n1785, u2_uk_n1797, u2_uk_n1803, u2_uk_n1807, u2_uk_n1808, u2_uk_n1816, 
      u2_uk_n1817, u2_uk_n1819, u2_uk_n1821, u2_uk_n1824, u2_uk_n1826, u2_uk_n1834, u2_uk_n1840, u2_uk_n1846, u2_uk_n1849, 
      u2_uk_n1851, u2_uk_n1852, u2_uk_n1855, u2_uk_n1856, u2_uk_n238, u2_uk_n299, u2_uk_n301, u2_uk_n305, u2_uk_n373, 
      u2_uk_n386, u2_uk_n408, u2_uk_n415, u2_uk_n421, u2_uk_n454, u2_uk_n456, u2_uk_n467, u2_uk_n503, u2_uk_n504, 
      u2_uk_n515, u2_uk_n520, u2_uk_n665, u2_uk_n682, u2_uk_n689, u2_uk_n939, u2_uk_n942, u2_uk_n943, u2_uk_n945, 
      u2_uk_n946, u2_uk_n985, u2_uk_n986, u2_uk_n987, u0_out12_11, u0_out12_14, u0_out12_19, u0_out12_25, u0_out12_29, 
      u0_out12_3, u0_out12_4, u0_out12_8, u0_out13_1, u0_out13_10, u0_out13_11, u0_out13_12, u0_out13_13, u0_out13_14, 
      u0_out13_17, u0_out13_18, u0_out13_19, u0_out13_2, u0_out13_20, u0_out13_22, u0_out13_23, u0_out13_25, u0_out13_26, 
      u0_out13_28, u0_out13_29, u0_out13_3, u0_out13_31, u0_out13_32, u0_out13_4, u0_out13_7, u0_out13_8, u0_out13_9, 
      u0_out14_11, u0_out14_12, u0_out14_14, u0_out14_15, u0_out14_19, u0_out14_21, u0_out14_22, u0_out14_25, u0_out14_27, 
      u0_out14_29, u0_out14_3, u0_out14_32, u0_out14_4, u0_out14_5, u0_out14_7, u0_out14_8, u0_out3_1, u0_out3_10, 
      u0_out3_11, u0_out3_12, u0_out3_13, u0_out3_14, u0_out3_15, u0_out3_16, u0_out3_17, u0_out3_18, u0_out3_19, 
      u0_out3_2, u0_out3_20, u0_out3_21, u0_out3_22, u0_out3_23, u0_out3_24, u0_out3_25, u0_out3_26, u0_out3_27, 
      u0_out3_28, u0_out3_29, u0_out3_3, u0_out3_30, u0_out3_31, u0_out3_32, u0_out3_4, u0_out3_5, u0_out3_6, 
      u0_out3_7, u0_out3_8, u0_out3_9, u0_out4_1, u0_out4_10, u0_out4_11, u0_out4_13, u0_out4_14, u0_out4_15, 
      u0_out4_16, u0_out4_17, u0_out4_18, u0_out4_19, u0_out4_2, u0_out4_20, u0_out4_21, u0_out4_23, u0_out4_24, 
      u0_out4_25, u0_out4_26, u0_out4_27, u0_out4_28, u0_out4_29, u0_out4_3, u0_out4_30, u0_out4_31, u0_out4_4, 
      u0_out4_5, u0_out4_6, u0_out4_8, u0_out4_9, u0_out6_1, u0_out6_10, u0_out6_11, u0_out6_13, u0_out6_16, 
      u0_out6_17, u0_out6_18, u0_out6_19, u0_out6_2, u0_out6_20, u0_out6_23, u0_out6_24, u0_out6_26, u0_out6_28, 
      u0_out6_29, u0_out6_30, u0_out6_31, u0_out6_4, u0_out6_6, u0_out6_9, u0_out7_1, u0_out7_10, u0_out7_13, 
      u0_out7_16, u0_out7_17, u0_out7_18, u0_out7_2, u0_out7_20, u0_out7_23, u0_out7_24, u0_out7_26, u0_out7_28, 
      u0_out7_30, u0_out7_31, u0_out7_6, u0_out7_9, u0_out9_1, u0_out9_10, u0_out9_11, u0_out9_12, u0_out9_13, 
      u0_out9_14, u0_out9_15, u0_out9_16, u0_out9_17, u0_out9_18, u0_out9_19, u0_out9_2, u0_out9_20, u0_out9_21, 
      u0_out9_22, u0_out9_23, u0_out9_24, u0_out9_25, u0_out9_26, u0_out9_27, u0_out9_28, u0_out9_29, u0_out9_3, 
      u0_out9_30, u0_out9_31, u0_out9_32, u0_out9_4, u0_out9_5, u0_out9_6, u0_out9_7, u0_out9_8, u0_out9_9, 
      u0_uk_n213, u0_uk_n223, u2_out0_11, u2_out0_12, u2_out0_13, u2_out0_14, u2_out0_15, u2_out0_18, u2_out0_19, 
      u2_out0_2, u2_out0_21, u2_out0_22, u2_out0_25, u2_out0_27, u2_out0_28, u2_out0_29, u2_out0_3, u2_out0_32, 
      u2_out0_4, u2_out0_5, u2_out0_7, u2_out0_8, u2_out10_1, u2_out10_10, u2_out10_11, u2_out10_12, u2_out10_14, 
      u2_out10_15, u2_out10_19, u2_out10_20, u2_out10_21, u2_out10_22, u2_out10_25, u2_out10_26, u2_out10_27, u2_out10_29, 
      u2_out10_3, u2_out10_32, u2_out10_4, u2_out10_5, u2_out10_7, u2_out10_8, u2_out11_1, u2_out11_10, u2_out11_11, 
      u2_out11_12, u2_out11_13, u2_out11_14, u2_out11_15, u2_out11_16, u2_out11_17, u2_out11_18, u2_out11_19, u2_out11_2, 
      u2_out11_20, u2_out11_21, u2_out11_22, u2_out11_23, u2_out11_24, u2_out11_25, u2_out11_26, u2_out11_27, u2_out11_28, 
      u2_out11_29, u2_out11_3, u2_out11_30, u2_out11_31, u2_out11_32, u2_out11_4, u2_out11_5, u2_out11_6, u2_out11_7, 
      u2_out11_8, u2_out11_9, u2_out12_11, u2_out12_12, u2_out12_13, u2_out12_14, u2_out12_15, u2_out12_17, u2_out12_18, 
      u2_out12_19, u2_out12_2, u2_out12_21, u2_out12_22, u2_out12_23, u2_out12_25, u2_out12_27, u2_out12_28, u2_out12_29, 
      u2_out12_3, u2_out12_31, u2_out12_32, u2_out12_4, u2_out12_5, u2_out12_7, u2_out12_8, u2_out12_9, u2_out13_11, 
      u2_out13_12, u2_out13_14, u2_out13_15, u2_out13_19, u2_out13_21, u2_out13_22, u2_out13_25, u2_out13_27, u2_out13_29, 
      u2_out13_3, u2_out13_32, u2_out13_4, u2_out13_5, u2_out13_7, u2_out13_8, u2_out14_1, u2_out14_10, u2_out14_11, 
      u2_out14_12, u2_out14_13, u2_out14_14, u2_out14_15, u2_out14_16, u2_out14_17, u2_out14_18, u2_out14_19, u2_out14_2, 
      u2_out14_20, u2_out14_21, u2_out14_22, u2_out14_23, u2_out14_24, u2_out14_25, u2_out14_26, u2_out14_27, u2_out14_28, 
      u2_out14_29, u2_out14_3, u2_out14_30, u2_out14_31, u2_out14_32, u2_out14_4, u2_out14_5, u2_out14_6, u2_out14_7, 
      u2_out14_8, u2_out14_9, u2_out2_1, u2_out2_10, u2_out2_11, u2_out2_12, u2_out2_13, u2_out2_14, u2_out2_15, 
      u2_out2_16, u2_out2_17, u2_out2_18, u2_out2_19, u2_out2_2, u2_out2_20, u2_out2_21, u2_out2_22, u2_out2_23, 
      u2_out2_24, u2_out2_25, u2_out2_26, u2_out2_27, u2_out2_28, u2_out2_29, u2_out2_3, u2_out2_30, u2_out2_31, 
      u2_out2_32, u2_out2_4, u2_out2_5, u2_out2_6, u2_out2_7, u2_out2_8, u2_out2_9, u2_out3_1, u2_out3_10, 
      u2_out3_11, u2_out3_13, u2_out3_14, u2_out3_15, u2_out3_16, u2_out3_17, u2_out3_18, u2_out3_19, u2_out3_2, 
      u2_out3_20, u2_out3_21, u2_out3_23, u2_out3_24, u2_out3_25, u2_out3_26, u2_out3_27, u2_out3_28, u2_out3_29, 
      u2_out3_3, u2_out3_30, u2_out3_31, u2_out3_4, u2_out3_5, u2_out3_6, u2_out3_8, u2_out3_9, u2_out4_1, 
      u2_out4_10, u2_out4_11, u2_out4_12, u2_out4_13, u2_out4_14, u2_out4_15, u2_out4_16, u2_out4_17, u2_out4_18, 
      u2_out4_19, u2_out4_2, u2_out4_20, u2_out4_21, u2_out4_22, u2_out4_23, u2_out4_24, u2_out4_25, u2_out4_26, 
      u2_out4_27, u2_out4_28, u2_out4_29, u2_out4_3, u2_out4_30, u2_out4_31, u2_out4_32, u2_out4_4, u2_out4_5, 
      u2_out4_6, u2_out4_7, u2_out4_8, u2_out4_9, u2_out5_1, u2_out5_10, u2_out5_11, u2_out5_12, u2_out5_13, 
      u2_out5_14, u2_out5_15, u2_out5_16, u2_out5_17, u2_out5_18, u2_out5_19, u2_out5_2, u2_out5_20, u2_out5_21, 
      u2_out5_22, u2_out5_23, u2_out5_24, u2_out5_25, u2_out5_26, u2_out5_27, u2_out5_28, u2_out5_29, u2_out5_3, 
      u2_out5_30, u2_out5_31, u2_out5_32, u2_out5_4, u2_out5_5, u2_out5_6, u2_out5_7, u2_out5_8, u2_out5_9, 
      u2_out6_1, u2_out6_10, u2_out6_11, u2_out6_12, u2_out6_13, u2_out6_14, u2_out6_15, u2_out6_16, u2_out6_17, 
      u2_out6_18, u2_out6_19, u2_out6_2, u2_out6_20, u2_out6_21, u2_out6_22, u2_out6_23, u2_out6_24, u2_out6_25, 
      u2_out6_26, u2_out6_27, u2_out6_28, u2_out6_29, u2_out6_3, u2_out6_30, u2_out6_31, u2_out6_32, u2_out6_4, 
      u2_out6_5, u2_out6_6, u2_out6_7, u2_out6_8, u2_out6_9, u2_out8_1, u2_out8_10, u2_out8_13, u2_out8_14, 
      u2_out8_16, u2_out8_17, u2_out8_18, u2_out8_2, u2_out8_20, u2_out8_23, u2_out8_24, u2_out8_25, u2_out8_26, 
      u2_out8_28, u2_out8_3, u2_out8_30, u2_out8_31, u2_out8_6, u2_out8_8, u2_out8_9, u2_out9_11, u2_out9_12, 
      u2_out9_15, u2_out9_17, u2_out9_19, u2_out9_21, u2_out9_22, u2_out9_23, u2_out9_27, u2_out9_29, u2_out9_31, 
      u2_out9_32, u2_out9_4, u2_out9_5, u2_out9_7, u2_out9_9, u2_uk_n10, u2_uk_n100, u2_uk_n102, u2_uk_n109, 
      u2_uk_n11, u2_uk_n110, u2_uk_n117, u2_uk_n118, u2_uk_n128, u2_uk_n129, u2_uk_n141, u2_uk_n142, u2_uk_n145, 
      u2_uk_n146, u2_uk_n147, u2_uk_n148, u2_uk_n155, u2_uk_n161, u2_uk_n162, u2_uk_n163, u2_uk_n164, u2_uk_n17, 
      u2_uk_n182, u2_uk_n187, u2_uk_n188, u2_uk_n191, u2_uk_n202, u2_uk_n203, u2_uk_n207, u2_uk_n208, u2_uk_n209, 
      u2_uk_n213, u2_uk_n214, u2_uk_n217, u2_uk_n220, u2_uk_n222, u2_uk_n223, u2_uk_n230, u2_uk_n231, u2_uk_n27, 
      u2_uk_n31, u2_uk_n60, u2_uk_n63, u2_uk_n83, u2_uk_n92, u2_uk_n93, u2_uk_n94, u2_uk_n99 );
  des_des_die_2 u2 ( u0_FP_33, u0_FP_34, u0_FP_36, u0_FP_37, u0_FP_39, u0_FP_41, u0_FP_42, u0_FP_43, u0_FP_44, 
      u0_FP_45, u0_FP_46, u0_FP_48, u0_FP_49, u0_FP_50, u0_FP_51, u0_FP_52, u0_FP_53, u0_FP_55, 
      u0_FP_56, u0_FP_57, u0_FP_60, u0_FP_63, u0_FP_64, u0_K11_37, u0_K11_42, u0_K11_48, u0_K12_25, 
      u0_K12_48, u0_K12_5, u0_K12_7, u0_K12_8, u0_K16_18, u0_K16_19, u0_K16_24, u0_K16_26, u0_K16_36, 
      u0_K16_5, u0_K16_8, u0_K1_30, u0_K1_31, u0_K2_11, u0_K2_12, u0_K2_18, u0_K2_20, u0_K2_5, 
      u0_K3_19, u0_K3_23, u0_K9_12, u0_K9_13, u0_K9_14, u0_K9_30, u0_K9_32, u0_K9_44, u0_K9_6, 
      u0_R0_1, u0_R0_13, u0_R0_15, u0_R0_32, u0_R0_4, u0_R0_7, u0_R0_8, u0_R0_9, u0_R10_1, 
      u0_R10_16, u0_R10_17, u0_R10_18, u0_R10_19, u0_R10_2, u0_R10_20, u0_R10_21, u0_R10_28, u0_R10_29, 
      u0_R10_3, u0_R10_4, u0_R10_5, u0_R1_1, u0_R1_12, u0_R1_13, u0_R1_14, u0_R1_15, u0_R1_16, 
      u0_R1_19, u0_R1_20, u0_R1_21, u0_R1_22, u0_R1_24, u0_R1_25, u0_R1_26, u0_R1_27, u0_R1_28, 
      u0_R1_29, u0_R1_30, u0_R1_32, u0_R6_17, u0_R6_24, u0_R6_26, u0_R6_28, u0_R6_29, u0_R7_1, 
      u0_R7_12, u0_R7_14, u0_R7_17, u0_R7_20, u0_R7_21, u0_R7_22, u0_R7_23, u0_R7_24, u0_R7_25, 
      u0_R7_28, u0_R7_29, u0_R7_32, u0_R7_4, u0_R7_5, u0_R7_8, u0_R7_9, u0_R9_1, u0_R9_16, 
      u0_R9_17, u0_R9_18, u0_R9_19, u0_R9_2, u0_R9_20, u0_R9_21, u0_R9_22, u0_R9_24, u0_R9_25, 
      u0_R9_26, u0_R9_27, u0_R9_29, u0_R9_3, u0_R9_30, u0_R9_31, u0_R9_32, u0_R9_4, u0_R9_5, 
      u0_desIn_r_1, u0_desIn_r_11, u0_desIn_r_17, u0_desIn_r_25, u0_desIn_r_27, u0_desIn_r_3, u0_desIn_r_35, u0_desIn_r_51, u0_desIn_r_57, 
      u0_desIn_r_59, u0_desIn_r_7, u0_desIn_r_9, u0_key_r_0, u0_key_r_14, u0_key_r_16, u0_key_r_2, u0_key_r_21, u0_key_r_22, 
      u0_key_r_23, u0_key_r_28, u0_key_r_29, u0_key_r_30, u0_key_r_35, u0_key_r_42, u0_key_r_50, u0_key_r_9, u0_u0_X_25, 
      u0_u0_X_28, u0_u0_X_33, u0_u0_X_42, u0_u0_X_44, u0_u0_X_45, u0_u0_X_46, u0_u10_X_34, u0_u10_X_41, u0_u10_X_43, 
      u0_u11_X_1, u0_u11_X_10, u0_u11_X_11, u0_u11_X_12, u0_u11_X_45, u0_u11_X_46, u0_u11_X_47, u0_u11_X_9, u0_u15_X_11, 
      u0_u15_X_13, u0_u15_X_22, u0_u15_X_33, u0_u15_X_4, u0_u15_X_44, u0_u15_X_45, u0_u15_X_9, u0_u1_X_15, u0_u1_X_16, 
      u0_u1_X_17, u0_u1_X_19, u0_u1_X_21, u0_u1_X_23, u0_u1_X_24, u0_u1_X_3, u0_u1_X_4, u0_u1_X_6, u0_u1_X_8, 
      u0_u1_X_9, u0_u2_X_24, u0_u2_X_26, u0_u2_X_27, u0_u2_X_34, u0_u2_X_46, u0_u7_X_25, u0_u7_X_27, u0_u7_X_28, 
      u0_u7_X_29, u0_u7_X_30, u0_u7_X_31, u0_u7_X_32, u0_u7_X_33, u0_u7_X_34, u0_u7_X_36, u0_u7_X_38, u0_u7_X_40, 
      u0_u7_X_45, u0_u7_X_46, u0_u7_X_47, u0_u7_X_48, u0_u8_X_10, u0_u8_X_15, u0_u8_X_16, u0_u8_X_18, u0_u8_X_20, 
      u0_u8_X_22, u0_u8_X_23, u0_u8_X_25, u0_u8_X_27, u0_u8_X_28, u0_u8_X_3, u0_u8_X_39, u0_u8_X_4, u0_u8_X_40, 
      u0_u8_X_45, u0_u8_X_46, u0_u8_X_9, u0_uk_K_r10_10, u0_uk_K_r10_18, u0_uk_K_r10_23, u0_uk_K_r10_27, u0_uk_K_r10_37, u0_uk_K_r10_42, 
      u0_uk_K_r14_10, u0_uk_K_r14_11, u0_uk_K_r14_12, u0_uk_K_r14_16, u0_uk_K_r14_18, u0_uk_K_r14_2, u0_uk_K_r14_45, u0_uk_K_r14_8, u0_uk_K_r14_9, 
      u0_uk_K_r1_15, u0_uk_K_r1_16, u0_uk_K_r1_21, u0_uk_K_r1_44, u0_uk_K_r1_7, u0_uk_K_r6_0, u0_uk_K_r6_22, u0_uk_K_r6_31, u0_uk_K_r7_26, 
      u0_uk_K_r9_0, u0_uk_K_r9_1, u0_uk_K_r9_19, u0_uk_K_r9_22, u0_uk_K_r9_25, u0_uk_K_r9_30, u0_uk_K_r9_35, u0_uk_K_r9_45, u0_uk_K_r9_7, 
      u0_uk_K_r9_9, u0_uk_n10, u0_uk_n102, u0_uk_n11, u0_uk_n110, u0_uk_n117, u0_uk_n129, u0_uk_n139, u0_uk_n142, 
      u0_uk_n144, u0_uk_n145, u0_uk_n147, u0_uk_n151, u0_uk_n156, u0_uk_n162, u0_uk_n163, u0_uk_n167, u0_uk_n168, 
      u0_uk_n171, u0_uk_n172, u0_uk_n174, u0_uk_n177, u0_uk_n178, u0_uk_n181, u0_uk_n182, u0_uk_n183, u0_uk_n184, 
      u0_uk_n185, u0_uk_n189, u0_uk_n192, u0_uk_n193, u0_uk_n195, u0_uk_n198, u0_uk_n199, u0_uk_n200, u0_uk_n201, 
      u0_uk_n202, u0_uk_n203, u0_uk_n204, u0_uk_n205, u0_uk_n207, u0_uk_n208, u0_uk_n210, u0_uk_n211, u0_uk_n213, 
      u0_uk_n215, u0_uk_n216, u0_uk_n217, u0_uk_n218, u0_uk_n219, u0_uk_n220, u0_uk_n222, u0_uk_n223, u0_uk_n224, 
      u0_uk_n231, u0_uk_n238, u0_uk_n242, u0_uk_n251, u0_uk_n252, u0_uk_n257, u0_uk_n272, u0_uk_n275, u0_uk_n276, 
      u0_uk_n278, u0_uk_n282, u0_uk_n283, u0_uk_n285, u0_uk_n289, u0_uk_n290, u0_uk_n293, u0_uk_n300, u0_uk_n307, 
      u0_uk_n31, u0_uk_n310, u0_uk_n314, u0_uk_n316, u0_uk_n320, u0_uk_n332, u0_uk_n341, u0_uk_n347, u0_uk_n348, 
      u0_uk_n355, u0_uk_n542, u0_uk_n544, u0_uk_n545, u0_uk_n546, u0_uk_n549, u0_uk_n550, u0_uk_n553, u0_uk_n554, 
      u0_uk_n555, u0_uk_n558, u0_uk_n560, u0_uk_n561, u0_uk_n562, u0_uk_n566, u0_uk_n567, u0_uk_n568, u0_uk_n570, 
      u0_uk_n574, u0_uk_n575, u0_uk_n577, u0_uk_n579, u0_uk_n580, u0_uk_n581, u0_uk_n583, u0_uk_n598, u0_uk_n60, 
      u0_uk_n604, u0_uk_n615, u0_uk_n627, u0_uk_n629, u0_uk_n632, u0_uk_n635, u0_uk_n636, u0_uk_n637, u0_uk_n639, 
      u0_uk_n640, u0_uk_n642, u0_uk_n643, u0_uk_n644, u0_uk_n645, u0_uk_n649, u0_uk_n650, u0_uk_n651, u0_uk_n652, 
      u0_uk_n653, u0_uk_n654, u0_uk_n657, u0_uk_n658, u0_uk_n659, u0_uk_n660, u0_uk_n661, u0_uk_n663, u0_uk_n666, 
      u0_uk_n668, u0_uk_n669, u0_uk_n670, u0_uk_n675, u0_uk_n687, u0_uk_n711, u0_uk_n719, u0_uk_n722, u0_uk_n723, 
      u0_uk_n725, u0_uk_n726, u0_uk_n727, u0_uk_n729, u0_uk_n731, u0_uk_n734, u0_uk_n735, u0_uk_n741, u0_uk_n746, 
      u0_uk_n748, u0_uk_n751, u0_uk_n855, u0_uk_n866, u0_uk_n868, u0_uk_n875, u0_uk_n883, u0_uk_n904, u0_uk_n963, 
      u0_uk_n985, u0_uk_n990, u1_FP_33, u1_FP_37, u1_FP_40, u1_FP_41, u1_FP_56, u1_FP_60, u1_FP_61, 
      u1_K10_1, u1_K10_11, u1_K10_13, u1_K10_14, u1_K10_18, u1_K10_2, u1_K10_20, u1_K10_23, u1_K10_24, 
      u1_K10_25, u1_K10_26, u1_K10_29, u1_K10_30, u1_K10_5, u1_K10_6, u1_K10_7, u1_K10_8, u1_K11_23, 
      u1_K11_25, u1_K11_29, u1_K12_18, u1_K12_19, u1_K12_2, u1_K12_20, u1_K12_24, u1_K12_25, u1_K12_26, 
      u1_K12_35, u1_K12_36, u1_K12_37, u1_K12_38, u1_K12_41, u1_K12_43, u1_K12_47, u1_K12_48, u1_K12_6, 
      u1_K12_8, u1_K13_29, u1_K13_30, u1_K13_31, u1_K13_32, u1_K13_35, u1_K13_37, u1_K14_29, u1_K14_30, 
      u1_K14_31, u1_K14_32, u1_K16_11, u1_K16_12, u1_K16_2, u1_K16_41, u1_K16_42, u1_K16_44, u1_K16_48, 
      u1_K16_6, u1_K16_8, u1_K1_17, u1_K1_19, u1_K2_1, u1_K2_11, u1_K2_12, u1_K2_13, u1_K2_17, 
      u1_K2_18, u1_K2_2, u1_K2_31, u1_K2_5, u1_K2_6, u1_K2_8, u1_K3_12, u1_K3_14, u1_K3_17, 
      u1_K3_18, u1_K3_19, u1_K3_20, u1_K3_23, u1_K3_25, u1_K3_26, u1_K3_29, u1_K3_31, u1_K3_35, 
      u1_K3_36, u1_K3_7, u1_K3_8, u1_K4_13, u1_K4_14, u1_K4_17, u1_K4_18, u1_K4_19, u1_K4_24, 
      u1_K4_30, u1_K4_32, u1_K4_35, u1_K4_36, u1_K4_37, u1_K4_38, u1_K4_41, u1_K4_42, u1_K4_43, 
      u1_K4_44, u1_K4_47, u1_K4_48, u1_K5_1, u1_K5_11, u1_K5_12, u1_K5_13, u1_K5_14, u1_K5_17, 
      u1_K5_18, u1_K5_2, u1_K5_25, u1_K5_26, u1_K5_29, u1_K5_30, u1_K5_31, u1_K5_32, u1_K5_37, 
      u1_K5_38, u1_K5_41, u1_K5_42, u1_K5_44, u1_K5_47, u1_K5_48, u1_K5_5, u1_K5_6, u1_K5_7, 
      u1_K5_8, u1_K6_1, u1_K6_11, u1_K6_12, u1_K6_13, u1_K6_14, u1_K6_20, u1_K6_23, u1_K6_24, 
      u1_K6_37, u1_K6_38, u1_K6_41, u1_K6_42, u1_K6_43, u1_K6_44, u1_K6_47, u1_K6_48, u1_K6_5, 
      u1_K6_6, u1_K6_7, u1_K6_8, u1_K7_19, u1_K7_23, u1_K7_26, u1_K7_29, u1_K7_30, u1_K7_31, 
      u1_K7_35, u1_K8_1, u1_K8_11, u1_K8_13, u1_K8_14, u1_K8_18, u1_K8_2, u1_K8_20, u1_K8_23, 
      u1_K8_24, u1_K8_25, u1_K8_26, u1_K8_30, u1_K8_31, u1_K8_32, u1_K8_35, u1_K8_36, u1_K8_38, 
      u1_K8_41, u1_K8_42, u1_K8_44, u1_K8_47, u1_K8_48, u1_K8_5, u1_K8_7, u1_K9_12, u1_K9_13, 
      u1_K9_14, u1_K9_17, u1_K9_7, u1_K9_8, u1_R0_1, u1_R0_12, u1_R0_13, u1_R0_20, u1_R0_21, 
      u1_R0_32, u1_R0_4, u1_R0_5, u1_R0_7, u1_R0_8, u1_R0_9, u1_R10_1, u1_R10_10, u1_R10_12, 
      u1_R10_13, u1_R10_14, u1_R10_16, u1_R10_17, u1_R10_24, u1_R10_25, u1_R10_28, u1_R10_29, u1_R10_32, 
      u1_R10_5, u1_R11_20, u1_R11_21, u1_R11_24, u1_R12_20, u1_R12_21, u1_R12_23, u1_R1_12, u1_R1_13, 
      u1_R1_16, u1_R1_17, u1_R1_20, u1_R1_24, u1_R1_25, u1_R1_4, u1_R1_5, u1_R1_9, u1_R2_1, 
      u1_R2_12, u1_R2_13, u1_R2_16, u1_R2_17, u1_R2_20, u1_R2_21, u1_R2_24, u1_R2_25, u1_R2_28, 
      u1_R2_29, u1_R2_32, u1_R2_8, u1_R2_9, u1_R3_1, u1_R3_12, u1_R3_13, u1_R3_16, u1_R3_17, 
      u1_R3_18, u1_R3_20, u1_R3_21, u1_R3_24, u1_R3_25, u1_R3_28, u1_R3_29, u1_R3_32, u1_R3_4, 
      u1_R3_5, u1_R3_8, u1_R3_9, u1_R4_1, u1_R4_13, u1_R4_14, u1_R4_16, u1_R4_17, u1_R4_24, 
      u1_R4_25, u1_R4_28, u1_R4_29, u1_R4_3, u1_R4_32, u1_R4_4, u1_R4_5, u1_R4_6, u1_R4_7, 
      u1_R4_8, u1_R4_9, u1_R5_12, u1_R5_13, u1_R5_16, u1_R5_17, u1_R5_18, u1_R5_20, u1_R5_21, 
      u1_R5_23, u1_R5_24, u1_R5_25, u1_R6_1, u1_R6_10, u1_R6_13, u1_R6_16, u1_R6_17, u1_R6_2, 
      u1_R6_20, u1_R6_21, u1_R6_24, u1_R6_25, u1_R6_28, u1_R6_29, u1_R6_32, u1_R6_4, u1_R6_8, 
      u1_R6_9, u1_R7_12, u1_R7_13, u1_R7_4, u1_R7_5, u1_R7_6, u1_R7_7, u1_R7_8, u1_R7_9, 
      u1_R8_1, u1_R8_13, u1_R8_15, u1_R8_16, u1_R8_17, u1_R8_20, u1_R8_21, u1_R8_32, u1_R8_4, 
      u1_R8_5, u1_R8_6, u1_R8_8, u1_R8_9, u1_R9_12, u1_R9_15, u1_R9_16, u1_R9_20, u1_R9_21, 
      u1_desIn_r_29, u1_desIn_r_37, u1_u0_X_13, u1_u0_X_14, u1_u0_X_15, u1_u0_X_16, u1_u0_X_21, u1_u0_X_22, u1_u0_X_23, 
      u1_u0_X_24, u1_u0_X_25, u1_u0_X_26, u1_u0_X_27, u1_u0_X_28, u1_u0_X_29, u1_u0_X_30, u1_u10_X_20, u1_u10_X_21, 
      u1_u10_X_24, u1_u10_X_26, u1_u10_X_27, u1_u10_X_28, u1_u11_X_10, u1_u11_X_11, u1_u11_X_12, u1_u11_X_13, u1_u11_X_14, 
      u1_u11_X_16, u1_u11_X_22, u1_u11_X_27, u1_u11_X_28, u1_u11_X_29, u1_u11_X_3, u1_u11_X_30, u1_u11_X_31, u1_u11_X_32, 
      u1_u11_X_33, u1_u11_X_34, u1_u11_X_39, u1_u11_X_4, u1_u11_X_40, u1_u11_X_45, u1_u11_X_46, u1_u11_X_5, u1_u11_X_7, 
      u1_u11_X_9, u1_u12_X_25, u1_u12_X_26, u1_u12_X_27, u1_u12_X_28, u1_u12_X_33, u1_u12_X_34, u1_u12_X_36, u1_u12_X_38, 
      u1_u12_X_39, u1_u12_X_40, u1_u12_X_41, u1_u12_X_42, u1_u13_X_13, u1_u13_X_14, u1_u13_X_15, u1_u13_X_16, u1_u13_X_17, 
      u1_u13_X_18, u1_u13_X_19, u1_u13_X_20, u1_u13_X_21, u1_u13_X_22, u1_u13_X_23, u1_u13_X_24, u1_u13_X_25, u1_u13_X_26, 
      u1_u13_X_27, u1_u13_X_28, u1_u13_X_33, u1_u13_X_35, u1_u13_X_36, u1_u15_X_1, u1_u15_X_10, u1_u15_X_3, u1_u15_X_38, 
      u1_u15_X_39, u1_u15_X_4, u1_u15_X_40, u1_u15_X_45, u1_u15_X_46, u1_u15_X_47, u1_u15_X_5, u1_u15_X_7, u1_u15_X_9, 
      u1_u1_X_15, u1_u1_X_16, u1_u1_X_3, u1_u1_X_33, u1_u1_X_34, u1_u1_X_35, u1_u1_X_36, u1_u1_X_4, u1_u1_X_9, 
      u1_u2_X_10, u1_u2_X_11, u1_u2_X_13, u1_u2_X_15, u1_u2_X_16, u1_u2_X_21, u1_u2_X_22, u1_u2_X_27, u1_u2_X_28, 
      u1_u2_X_30, u1_u2_X_32, u1_u2_X_33, u1_u2_X_34, u1_u2_X_9, u1_u3_X_15, u1_u3_X_16, u1_u3_X_21, u1_u3_X_22, 
      u1_u3_X_27, u1_u3_X_28, u1_u3_X_33, u1_u3_X_34, u1_u3_X_39, u1_u3_X_40, u1_u3_X_45, u1_u3_X_46, u1_u4_X_10, 
      u1_u4_X_15, u1_u4_X_16, u1_u4_X_28, u1_u4_X_3, u1_u4_X_33, u1_u4_X_34, u1_u4_X_39, u1_u4_X_4, u1_u4_X_40, 
      u1_u4_X_45, u1_u4_X_46, u1_u4_X_9, u1_u5_X_15, u1_u5_X_16, u1_u5_X_17, u1_u5_X_19, u1_u5_X_22, u1_u5_X_3, 
      u1_u5_X_39, u1_u5_X_40, u1_u5_X_45, u1_u5_X_46, u1_u6_X_21, u1_u6_X_22, u1_u6_X_28, u1_u6_X_33, u1_u7_X_10, 
      u1_u7_X_16, u1_u7_X_17, u1_u7_X_19, u1_u7_X_21, u1_u7_X_22, u1_u7_X_27, u1_u7_X_28, u1_u7_X_33, u1_u7_X_34, 
      u1_u7_X_39, u1_u7_X_4, u1_u7_X_40, u1_u7_X_45, u1_u7_X_46, u1_u7_X_6, u1_u7_X_8, u1_u7_X_9, u1_u8_X_15, 
      u1_u8_X_16, u1_u9_X_10, u1_u9_X_15, u1_u9_X_16, u1_u9_X_17, u1_u9_X_19, u1_u9_X_21, u1_u9_X_27, u1_u9_X_28, 
      u1_u9_X_3, u1_u9_X_4, u1_uk_n1002, u1_uk_n1003, u1_uk_n1021, u1_uk_n1023, u1_uk_n1029, u1_uk_n1034, u1_uk_n1038, 
      u1_uk_n1054, u1_uk_n1056, u1_uk_n1057, u1_uk_n1058, u1_uk_n1060, u1_uk_n1063, u1_uk_n1076, u1_uk_n1079, u1_uk_n1080, 
      u1_uk_n1083, u1_uk_n1088, u1_uk_n1090, u1_uk_n1092, u1_uk_n1096, u1_uk_n1101, u1_uk_n1104, u1_uk_n1109, u1_uk_n1113, 
      u1_uk_n1114, u1_uk_n1115, u1_uk_n1118, u1_uk_n1119, u1_uk_n1121, u1_uk_n1128, u1_uk_n1130, u1_uk_n1134, u1_uk_n1138, 
      u1_uk_n1140, u1_uk_n1143, u1_uk_n1147, u1_uk_n1148, u1_uk_n1153, u1_uk_n1171, u1_uk_n299, u1_uk_n312, u1_uk_n376, 
      u1_uk_n386, u1_uk_n407, u1_uk_n421, u1_uk_n504, u1_uk_n509, u1_uk_n515, u1_uk_n520, u1_uk_n524, u1_uk_n605, 
      u1_uk_n608, u1_uk_n955, u1_uk_n989, u1_uk_n993, u2_K10_11, u2_K10_13, u2_K10_14, u2_K10_17, u2_K10_18, 
      u2_K10_19, u2_K10_20, u2_K10_23, u2_K10_24, u2_K10_25, u2_K10_26, u2_K10_7, u2_K10_8, u2_K2_1, 
      u2_K2_11, u2_K2_12, u2_K2_13, u2_K2_17, u2_K2_18, u2_K2_2, u2_K2_20, u2_K2_23, u2_K2_24, 
      u2_K2_25, u2_K2_26, u2_K2_29, u2_K2_30, u2_K2_31, u2_K2_35, u2_K2_36, u2_K2_37, u2_K2_38, 
      u2_K2_42, u2_K2_44, u2_K2_47, u2_K2_48, u2_K2_5, u2_K2_6, u2_K2_8, u2_R0_1, u2_R0_12, 
      u2_R0_13, u2_R0_16, u2_R0_17, u2_R0_19, u2_R0_20, u2_R0_21, u2_R0_24, u2_R0_25, u2_R0_29, 
      u2_R0_32, u2_R0_4, u2_R0_5, u2_R0_7, u2_R0_8, u2_R0_9, u2_R8_12, u2_R8_13, u2_R8_15, 
      u2_R8_16, u2_R8_17, u2_R8_4, u2_R8_5, u2_R8_6, u2_R8_8, u2_R8_9, u2_u1_X_15, u2_u1_X_16, 
      u2_u1_X_21, u2_u1_X_22, u2_u1_X_27, u2_u1_X_3, u2_u1_X_33, u2_u1_X_34, u2_u1_X_39, u2_u1_X_4, u2_u1_X_40, 
      u2_u1_X_41, u2_u1_X_43, u2_u1_X_45, u2_u1_X_46, u2_u1_X_9, u2_u9_X_10, u2_u9_X_15, u2_u9_X_16, u2_u9_X_21, 
      u2_u9_X_27, u2_u9_X_28, u2_u9_X_29, u2_u9_X_30, u2_uk_n1004, u2_uk_n240, u2_uk_n257, u2_uk_n308, u2_uk_n991, 
      u2_uk_n993, u2_uk_n995, u2_uk_n998, u2_uk_n999, u0_out0_11, u0_out0_12, u0_out0_14, u0_out0_15, u0_out0_19, 
      u0_out0_21, u0_out0_22, u0_out0_25, u0_out0_27, u0_out0_29, u0_out0_3, u0_out0_32, u0_out0_4, u0_out0_5, 
      u0_out0_7, u0_out0_8, u0_out10_11, u0_out10_12, u0_out10_14, u0_out10_15, u0_out10_17, u0_out10_19, u0_out10_21, 
      u0_out10_22, u0_out10_23, u0_out10_25, u0_out10_27, u0_out10_29, u0_out10_3, u0_out10_31, u0_out10_32, u0_out10_4, 
      u0_out10_5, u0_out10_7, u0_out10_8, u0_out10_9, u0_out11_13, u0_out11_14, u0_out11_15, u0_out11_17, u0_out11_18, 
      u0_out11_2, u0_out11_21, u0_out11_23, u0_out11_25, u0_out11_27, u0_out11_28, u0_out11_3, u0_out11_31, u0_out11_5, 
      u0_out11_8, u0_out11_9, u0_out15_1, u0_out15_10, u0_out15_11, u0_out15_13, u0_out15_14, u0_out15_15, u0_out15_16, 
      u0_out15_17, u0_out15_18, u0_out15_19, u0_out15_2, u0_out15_20, u0_out15_21, u0_out15_23, u0_out15_24, u0_out15_25, 
      u0_out15_26, u0_out15_27, u0_out15_28, u0_out15_29, u0_out15_3, u0_out15_30, u0_out15_31, u0_out15_4, u0_out15_5, 
      u0_out15_6, u0_out15_8, u0_out15_9, u0_out1_1, u0_out1_10, u0_out1_13, u0_out1_16, u0_out1_17, u0_out1_18, 
      u0_out1_2, u0_out1_20, u0_out1_23, u0_out1_24, u0_out1_26, u0_out1_28, u0_out1_30, u0_out1_31, u0_out1_6, 
      u0_out1_9, u0_out2_1, u0_out2_10, u0_out2_11, u0_out2_12, u0_out2_14, u0_out2_15, u0_out2_19, u0_out2_20, 
      u0_out2_21, u0_out2_22, u0_out2_25, u0_out2_26, u0_out2_27, u0_out2_29, u0_out2_3, u0_out2_32, u0_out2_4, 
      u0_out2_5, u0_out2_7, u0_out2_8, u0_out7_11, u0_out7_12, u0_out7_14, u0_out7_15, u0_out7_19, u0_out7_21, 
      u0_out7_22, u0_out7_25, u0_out7_27, u0_out7_29, u0_out7_3, u0_out7_32, u0_out7_4, u0_out7_5, u0_out7_7, 
      u0_out7_8, u0_out8_1, u0_out8_10, u0_out8_11, u0_out8_12, u0_out8_13, u0_out8_14, u0_out8_15, u0_out8_16, 
      u0_out8_17, u0_out8_18, u0_out8_19, u0_out8_2, u0_out8_20, u0_out8_21, u0_out8_22, u0_out8_23, u0_out8_24, 
      u0_out8_25, u0_out8_26, u0_out8_27, u0_out8_28, u0_out8_29, u0_out8_3, u0_out8_30, u0_out8_31, u0_out8_32, 
      u0_out8_4, u0_out8_5, u0_out8_6, u0_out8_7, u0_out8_8, u0_out8_9, u0_uk_n100, u0_uk_n109, u0_uk_n118, 
      u0_uk_n128, u0_uk_n146, u0_uk_n148, u0_uk_n155, u0_uk_n161, u0_uk_n164, u0_uk_n17, u0_uk_n187, u0_uk_n188, 
      u0_uk_n191, u0_uk_n209, u0_uk_n214, u0_uk_n230, u0_uk_n240, u0_uk_n27, u0_uk_n63, u0_uk_n83, u0_uk_n92, 
      u0_uk_n93, u0_uk_n94, u0_uk_n99, u1_out0_1, u1_out0_10, u1_out0_14, u1_out0_16, u1_out0_20, u1_out0_24, 
      u1_out0_25, u1_out0_26, u1_out0_3, u1_out0_30, u1_out0_6, u1_out0_8, u1_out10_1, u1_out10_10, u1_out10_14, 
      u1_out10_20, u1_out10_25, u1_out10_26, u1_out10_3, u1_out10_8, u1_out11_1, u1_out11_10, u1_out11_11, u1_out11_12, 
      u1_out11_13, u1_out11_14, u1_out11_15, u1_out11_16, u1_out11_17, u1_out11_18, u1_out11_19, u1_out11_2, u1_out11_20, 
      u1_out11_21, u1_out11_22, u1_out11_23, u1_out11_24, u1_out11_25, u1_out11_26, u1_out11_27, u1_out11_28, u1_out11_29, 
      u1_out11_3, u1_out11_30, u1_out11_31, u1_out11_32, u1_out11_4, u1_out11_5, u1_out11_6, u1_out11_7, u1_out11_8, 
      u1_out11_9, u1_out12_11, u1_out12_12, u1_out12_14, u1_out12_19, u1_out12_22, u1_out12_25, u1_out12_29, u1_out12_3, 
      u1_out12_32, u1_out12_4, u1_out12_7, u1_out12_8, u1_out13_1, u1_out13_10, u1_out13_11, u1_out13_14, u1_out13_16, 
      u1_out13_19, u1_out13_20, u1_out13_24, u1_out13_25, u1_out13_26, u1_out13_29, u1_out13_3, u1_out13_30, u1_out13_4, 
      u1_out13_6, u1_out13_8, u1_out15_12, u1_out15_13, u1_out15_15, u1_out15_17, u1_out15_18, u1_out15_2, u1_out15_21, 
      u1_out15_22, u1_out15_23, u1_out15_27, u1_out15_28, u1_out15_31, u1_out15_32, u1_out15_5, u1_out15_7, u1_out15_9, 
      u1_out1_11, u1_out1_13, u1_out1_16, u1_out1_17, u1_out1_18, u1_out1_19, u1_out1_2, u1_out1_23, u1_out1_24, 
      u1_out1_28, u1_out1_29, u1_out1_30, u1_out1_31, u1_out1_4, u1_out1_6, u1_out1_9, u1_out2_1, u1_out2_10, 
      u1_out2_11, u1_out2_13, u1_out2_14, u1_out2_16, u1_out2_18, u1_out2_19, u1_out2_2, u1_out2_20, u1_out2_24, 
      u1_out2_25, u1_out2_26, u1_out2_28, u1_out2_29, u1_out2_3, u1_out2_30, u1_out2_4, u1_out2_6, u1_out2_8, 
      u1_out3_1, u1_out3_10, u1_out3_11, u1_out3_12, u1_out3_14, u1_out3_15, u1_out3_16, u1_out3_19, u1_out3_20, 
      u1_out3_21, u1_out3_22, u1_out3_24, u1_out3_25, u1_out3_26, u1_out3_27, u1_out3_29, u1_out3_3, u1_out3_30, 
      u1_out3_32, u1_out3_4, u1_out3_5, u1_out3_6, u1_out3_7, u1_out3_8, u1_out4_11, u1_out4_12, u1_out4_13, 
      u1_out4_14, u1_out4_15, u1_out4_16, u1_out4_17, u1_out4_18, u1_out4_19, u1_out4_2, u1_out4_21, u1_out4_22, 
      u1_out4_23, u1_out4_24, u1_out4_25, u1_out4_27, u1_out4_28, u1_out4_29, u1_out4_3, u1_out4_30, u1_out4_31, 
      u1_out4_32, u1_out4_4, u1_out4_5, u1_out4_6, u1_out4_7, u1_out4_8, u1_out4_9, u1_out5_1, u1_out5_10, 
      u1_out5_12, u1_out5_13, u1_out5_15, u1_out5_16, u1_out5_17, u1_out5_18, u1_out5_2, u1_out5_20, u1_out5_21, 
      u1_out5_22, u1_out5_23, u1_out5_24, u1_out5_26, u1_out5_27, u1_out5_28, u1_out5_30, u1_out5_31, u1_out5_32, 
      u1_out5_5, u1_out5_6, u1_out5_7, u1_out5_9, u1_out6_1, u1_out6_10, u1_out6_11, u1_out6_14, u1_out6_19, 
      u1_out6_20, u1_out6_25, u1_out6_26, u1_out6_29, u1_out6_3, u1_out6_4, u1_out6_8, u1_out7_1, u1_out7_10, 
      u1_out7_11, u1_out7_12, u1_out7_13, u1_out7_14, u1_out7_15, u1_out7_16, u1_out7_17, u1_out7_18, u1_out7_19, 
      u1_out7_2, u1_out7_20, u1_out7_21, u1_out7_22, u1_out7_23, u1_out7_24, u1_out7_25, u1_out7_26, u1_out7_27, 
      u1_out7_28, u1_out7_29, u1_out7_3, u1_out7_30, u1_out7_31, u1_out7_32, u1_out7_4, u1_out7_5, u1_out7_6, 
      u1_out7_7, u1_out7_8, u1_out7_9, u1_out8_13, u1_out8_16, u1_out8_18, u1_out8_2, u1_out8_24, u1_out8_28, 
      u1_out8_30, u1_out8_6, u1_out9_1, u1_out9_10, u1_out9_13, u1_out9_14, u1_out9_16, u1_out9_17, u1_out9_18, 
      u1_out9_2, u1_out9_20, u1_out9_23, u1_out9_24, u1_out9_25, u1_out9_26, u1_out9_28, u1_out9_3, u1_out9_30, 
      u1_out9_31, u1_out9_6, u1_out9_8, u1_out9_9, u2_out1_1, u2_out1_10, u2_out1_11, u2_out1_12, u2_out1_13, 
      u2_out1_14, u2_out1_15, u2_out1_16, u2_out1_17, u2_out1_18, u2_out1_19, u2_out1_2, u2_out1_20, u2_out1_21, 
      u2_out1_22, u2_out1_23, u2_out1_24, u2_out1_25, u2_out1_26, u2_out1_27, u2_out1_28, u2_out1_29, u2_out1_3, 
      u2_out1_30, u2_out1_31, u2_out1_32, u2_out1_4, u2_out1_5, u2_out1_6, u2_out1_7, u2_out1_8, u2_out1_9, 
      u2_out9_1, u2_out9_10, u2_out9_13, u2_out9_14, u2_out9_16, u2_out9_18, u2_out9_2, u2_out9_20, u2_out9_24, 
      u2_out9_25, u2_out9_26, u2_out9_28, u2_out9_3, u2_out9_30, u2_out9_6, u2_out9_8 );
  des_des_die_3 u3 ( u0_FP_56, u0_FP_57, u0_FP_58, u0_FP_59, u0_FP_60, u0_K12_19, u0_K12_35, u0_K12_36, u0_K13_41, 
      u0_K15_13, u0_K16_38, u0_K1_13, u0_K1_14, u0_K1_17, u0_K2_29, u0_K2_30, u0_K2_31, u0_K3_12, 
      u0_K3_13, u0_K3_14, u0_K3_17, u0_K3_18, u0_K3_5, u0_K3_6, u0_K6_11, u0_K6_13, u0_K6_19, 
      u0_K6_20, u0_K6_23, u0_K6_24, u0_K6_41, u0_R0_18, u0_R0_19, u0_R0_20, u0_R0_21, u0_R0_28, 
      u0_R10_12, u0_R10_14, u0_R10_16, u0_R10_17, u0_R10_20, u0_R10_21, u0_R10_24, u0_R10_25, u0_R10_28, 
      u0_R10_29, u0_R11_10, u0_R11_11, u0_R11_12, u0_R11_13, u0_R11_14, u0_R11_15, u0_R11_16, u0_R11_2, 
      u0_R11_28, u0_R11_3, u0_R11_32, u0_R11_5, u0_R11_6, u0_R12_30, u0_R13_8, u0_R1_1, u0_R1_12, 
      u0_R1_13, u0_R1_3, u0_R1_32, u0_R1_4, u0_R1_5, u0_R1_8, u0_R1_9, u0_R4_1, u0_R4_12, 
      u0_R4_13, u0_R4_16, u0_R4_17, u0_R4_19, u0_R4_20, u0_R4_21, u0_R4_22, u0_R4_24, u0_R4_25, 
      u0_R4_26, u0_R4_27, u0_R4_28, u0_R4_29, u0_R4_3, u0_R4_30, u0_R4_32, u0_R4_4, u0_R4_5, 
      u0_R4_8, u0_R4_9, u0_R9_10, u0_R9_11, u0_R9_12, u0_R9_13, u0_R9_16, u0_R9_17, u0_R9_4, 
      u0_R9_5, u0_R9_6, u0_R9_7, u0_R9_8, u0_R9_9, u0_desIn_r_15, u0_desIn_r_23, u0_desIn_r_29, u0_desIn_r_3, 
      u0_desIn_r_31, u0_desIn_r_37, u0_desIn_r_39, u0_desIn_r_47, u0_desIn_r_5, u0_desIn_r_55, u0_desIn_r_57, u0_desIn_r_63, u0_desIn_r_7, 
      u0_key_r_11, u0_key_r_12, u0_key_r_13, u0_key_r_19, u0_key_r_20, u0_key_r_4, u0_key_r_41, u0_key_r_47, u0_key_r_48, 
      u0_key_r_5, u0_key_r_54, u0_key_r_55, u0_key_r_6, u0_u0_X_15, u0_u0_X_16, u0_u0_X_21, u0_u0_X_22, u0_u0_X_23, 
      u0_u10_X_21, u0_u10_X_22, u0_u11_X_13, u0_u11_X_14, u0_u11_X_15, u0_u11_X_16, u0_u11_X_18, u0_u11_X_20, u0_u11_X_22, 
      u0_u11_X_33, u0_u11_X_34, u0_u11_X_39, u0_u11_X_40, u0_u12_X_10, u0_u12_X_11, u0_u12_X_12, u0_u12_X_13, u0_u12_X_14, 
      u0_u12_X_2, u0_u12_X_24, u0_u12_X_37, u0_u12_X_38, u0_u12_X_39, u0_u12_X_40, u0_u12_X_42, u0_u12_X_44, u0_u12_X_45, 
      u0_u12_X_46, u0_u12_X_48, u0_u12_X_5, u0_u12_X_7, u0_u13_X_43, u0_u13_X_44, u0_u13_X_46, u0_u13_X_47, u0_u13_X_48, 
      u0_u14_X_10, u0_u14_X_12, u0_u14_X_14, u0_u14_X_15, u0_u14_X_16, u0_u14_X_17, u0_u14_X_18, u0_u14_X_19, u0_u14_X_20, 
      u0_u14_X_21, u0_u14_X_22, u0_u14_X_23, u0_u14_X_24, u0_u14_X_7, u0_u14_X_8, u0_u14_X_9, u0_u15_X_42, u0_u1_X_25, 
      u0_u1_X_26, u0_u1_X_33, u0_u1_X_34, u0_u1_X_35, u0_u1_X_36, u0_u1_X_37, u0_u1_X_38, u0_u1_X_39, u0_u1_X_40, 
      u0_u1_X_42, u0_u2_X_10, u0_u2_X_15, u0_u2_X_16, u0_u2_X_3, u0_u2_X_9, u0_u5_X_10, u0_u5_X_15, u0_u5_X_16, 
      u0_u5_X_21, u0_u5_X_22, u0_u5_X_27, u0_u5_X_3, u0_u5_X_34, u0_u5_X_46, u0_u5_X_9, u0_uk_K_r0_15, u0_uk_K_r0_28, 
      u0_uk_K_r0_36, u0_uk_K_r0_49, u0_uk_K_r0_7, u0_uk_K_r10_18, u0_uk_K_r10_23, u0_uk_K_r10_28, u0_uk_K_r10_32, u0_uk_K_r10_41, u0_uk_K_r10_44, 
      u0_uk_K_r10_9, u0_uk_K_r11_19, u0_uk_K_r11_20, u0_uk_K_r11_24, u0_uk_K_r11_25, u0_uk_K_r11_27, u0_uk_K_r11_29, u0_uk_K_r11_33, u0_uk_K_r11_39, 
      u0_uk_K_r11_4, u0_uk_K_r12_16, u0_uk_K_r13_25, u0_uk_K_r14_15, u0_uk_K_r14_2, u0_uk_K_r14_50, u0_uk_K_r4_0, u0_uk_K_r4_23, u0_uk_K_r4_33, 
      u0_uk_K_r4_35, u0_uk_K_r4_38, u0_uk_K_r4_41, u0_uk_K_r4_47, u0_uk_K_r9_25, u0_uk_K_r9_27, u0_uk_K_r9_33, u0_uk_K_r9_6, u0_uk_n100, 
      u0_uk_n1000, u0_uk_n1001, u0_uk_n1002, u0_uk_n1004, u0_uk_n101, u0_uk_n106, u0_uk_n107, u0_uk_n108, u0_uk_n109, 
      u0_uk_n115, u0_uk_n118, u0_uk_n121, u0_uk_n122, u0_uk_n126, u0_uk_n127, u0_uk_n128, u0_uk_n131, u0_uk_n139, 
      u0_uk_n143, u0_uk_n144, u0_uk_n146, u0_uk_n148, u0_uk_n153, u0_uk_n155, u0_uk_n161, u0_uk_n164, u0_uk_n172, 
      u0_uk_n173, u0_uk_n179, u0_uk_n180, u0_uk_n187, u0_uk_n188, u0_uk_n190, u0_uk_n191, u0_uk_n195, u0_uk_n196, 
      u0_uk_n197, u0_uk_n200, u0_uk_n201, u0_uk_n206, u0_uk_n212, u0_uk_n213, u0_uk_n214, u0_uk_n215, u0_uk_n221, 
      u0_uk_n225, u0_uk_n230, u0_uk_n240, u0_uk_n257, u0_uk_n410, u0_uk_n411, u0_uk_n412, u0_uk_n413, u0_uk_n414, 
      u0_uk_n418, u0_uk_n419, u0_uk_n420, u0_uk_n423, u0_uk_n424, u0_uk_n425, u0_uk_n426, u0_uk_n428, u0_uk_n429, 
      u0_uk_n430, u0_uk_n432, u0_uk_n433, u0_uk_n434, u0_uk_n436, u0_uk_n438, u0_uk_n439, u0_uk_n440, u0_uk_n442, 
      u0_uk_n445, u0_uk_n446, u0_uk_n447, u0_uk_n448, u0_uk_n450, u0_uk_n547, u0_uk_n552, u0_uk_n557, u0_uk_n562, 
      u0_uk_n565, u0_uk_n568, u0_uk_n573, u0_uk_n578, u0_uk_n58, u0_uk_n63, u0_uk_n632, u0_uk_n643, u0_uk_n657, 
      u0_uk_n670, u0_uk_n674, u0_uk_n684, u0_uk_n690, u0_uk_n696, u0_uk_n697, u0_uk_n699, u0_uk_n786, u0_uk_n793, 
      u0_uk_n799, u0_uk_n8, u0_uk_n800, u0_uk_n83, u0_uk_n869, u0_uk_n892, u0_uk_n898, u0_uk_n91, u0_uk_n92, 
      u0_uk_n93, u0_uk_n94, u0_uk_n949, u0_uk_n950, u0_uk_n956, u0_uk_n96, u0_uk_n976, u0_uk_n982, u0_uk_n99, 
      u0_uk_n999, u1_FP_40, u1_FP_41, u1_FP_44, u1_FP_45, u1_FP_52, u1_FP_53, u1_FP_55, u1_FP_56, 
      u1_K10_31, u1_K10_32, u1_K10_36, u1_K10_41, u1_K10_42, u1_K10_43, u1_K10_44, u1_K10_47, u1_K10_48, 
      u1_K11_11, u1_K11_13, u1_K11_2, u1_K11_32, u1_K11_35, u1_K11_37, u1_K11_38, u1_K11_48, u1_K11_7, 
      u1_K13_14, u1_K13_17, u1_K13_18, u1_K13_20, u1_K13_48, u1_K13_8, u1_K14_1, u1_K14_2, u1_K14_42, 
      u1_K14_44, u1_K14_47, u1_K14_48, u1_K15_11, u1_K15_12, u1_K15_13, u1_K15_14, u1_K15_18, u1_K15_2, 
      u1_K15_20, u1_K15_23, u1_K15_24, u1_K15_25, u1_K15_29, u1_K15_31, u1_K15_32, u1_K15_35, u1_K15_36, 
      u1_K15_37, u1_K15_41, u1_K15_42, u1_K15_44, u1_K15_48, u1_K15_5, u1_K15_6, u1_K15_7, u1_K16_13, 
      u1_K16_14, u1_K16_17, u1_K16_18, u1_K16_19, u1_K16_20, u1_K16_30, u1_K16_31, u1_K16_32, u1_K16_35, 
      u1_K1_1, u1_K1_43, u1_K1_47, u1_K1_6, u1_K1_8, u1_K2_20, u1_K2_23, u1_K2_24, u1_K2_25, 
      u1_K2_26, u1_K2_29, u1_K2_30, u1_K2_42, u1_K2_43, u1_K2_44, u1_K2_47, u1_K2_48, u1_K3_1, 
      u1_K3_2, u1_K3_37, u1_K3_38, u1_K3_41, u1_K3_42, u1_K3_43, u1_K3_44, u1_K3_47, u1_K3_48, 
      u1_K3_5, u1_K3_6, u1_K4_1, u1_K4_11, u1_K4_12, u1_K4_6, u1_K5_19, u1_K5_23, u1_K5_24, 
      u1_K6_25, u1_K6_26, u1_K6_29, u1_K6_30, u1_K6_31, u1_K6_32, u1_K6_35, u1_K6_36, u1_K7_1, 
      u1_K7_11, u1_K7_14, u1_K7_17, u1_K7_18, u1_K7_2, u1_K7_37, u1_K7_38, u1_K7_41, u1_K7_43, 
      u1_K7_44, u1_K7_47, u1_K7_48, u1_K7_5, u1_K7_7, u1_K9_23, u1_K9_24, u1_K9_25, u1_K9_29, 
      u1_K9_31, u1_K9_36, u1_K9_37, u1_K9_38, u1_K9_43, u1_K9_44, u1_K9_47, u1_K9_5, u1_K9_6, 
      u1_R0_1, u1_R0_12, u1_R0_13, u1_R0_16, u1_R0_17, u1_R0_20, u1_R0_21, u1_R0_28, u1_R0_29, 
      u1_R0_32, u1_R11_1, u1_R11_10, u1_R11_12, u1_R11_13, u1_R11_4, u1_R11_5, u1_R11_8, u1_R11_9, 
      u1_R12_1, u1_R12_29, u1_R12_32, u1_R13_1, u1_R13_13, u1_R13_16, u1_R13_17, u1_R13_20, u1_R13_21, 
      u1_R13_24, u1_R13_25, u1_R13_28, u1_R13_29, u1_R13_4, u1_R13_5, u1_R13_8, u1_R13_9, u1_R1_1, 
      u1_R1_24, u1_R1_25, u1_R1_28, u1_R1_29, u1_R1_32, u1_R1_4, u1_R1_5, u1_R2_1, u1_R2_2, 
      u1_R2_32, u1_R2_5, u1_R2_7, u1_R2_8, u1_R2_9, u1_R3_12, u1_R3_13, u1_R3_15, u1_R3_16, 
      u1_R3_17, u1_R4_16, u1_R4_17, u1_R4_20, u1_R4_21, u1_R4_24, u1_R4_25, u1_R5_1, u1_R5_12, 
      u1_R5_13, u1_R5_24, u1_R5_25, u1_R5_28, u1_R5_29, u1_R5_31, u1_R5_32, u1_R5_4, u1_R5_5, 
      u1_R5_8, u1_R5_9, u1_R7_1, u1_R7_12, u1_R7_13, u1_R7_15, u1_R7_16, u1_R7_17, u1_R7_18, 
      u1_R7_20, u1_R7_24, u1_R7_25, u1_R7_28, u1_R7_29, u1_R7_32, u1_R7_4, u1_R7_5, u1_R8_1, 
      u1_R8_20, u1_R8_21, u1_R8_22, u1_R8_24, u1_R8_25, u1_R8_28, u1_R8_29, u1_R8_32, u1_R9_1, 
      u1_R9_12, u1_R9_20, u1_R9_21, u1_R9_23, u1_R9_24, u1_R9_25, u1_R9_4, u1_R9_8, u1_R9_9, 
      u1_desIn_r_25, u1_desIn_r_39, u1_desIn_r_57, u1_u0_X_10, u1_u0_X_11, u1_u0_X_12, u1_u0_X_2, u1_u0_X_3, u1_u0_X_31, 
      u1_u0_X_32, u1_u0_X_33, u1_u0_X_34, u1_u0_X_35, u1_u0_X_36, u1_u0_X_37, u1_u0_X_38, u1_u0_X_39, u1_u0_X_4, 
      u1_u0_X_40, u1_u0_X_42, u1_u0_X_44, u1_u0_X_45, u1_u0_X_46, u1_u0_X_48, u1_u0_X_5, u1_u0_X_7, u1_u0_X_9, 
      u1_u10_X_1, u1_u10_X_10, u1_u10_X_15, u1_u10_X_16, u1_u10_X_18, u1_u10_X_3, u1_u10_X_33, u1_u10_X_39, u1_u10_X_4, 
      u1_u10_X_40, u1_u10_X_41, u1_u10_X_42, u1_u10_X_43, u1_u10_X_44, u1_u10_X_45, u1_u10_X_46, u1_u10_X_47, u1_u10_X_6, 
      u1_u10_X_8, u1_u10_X_9, u1_u12_X_1, u1_u12_X_10, u1_u12_X_16, u1_u12_X_21, u1_u12_X_22, u1_u12_X_23, u1_u12_X_24, 
      u1_u12_X_3, u1_u12_X_4, u1_u12_X_43, u1_u12_X_44, u1_u12_X_45, u1_u12_X_46, u1_u12_X_47, u1_u12_X_9, u1_u13_X_10, 
      u1_u13_X_11, u1_u13_X_12, u1_u13_X_3, u1_u13_X_37, u1_u13_X_38, u1_u13_X_39, u1_u13_X_4, u1_u13_X_40, u1_u13_X_41, 
      u1_u13_X_43, u1_u13_X_45, u1_u13_X_46, u1_u13_X_5, u1_u13_X_6, u1_u13_X_7, u1_u13_X_8, u1_u13_X_9, u1_u14_X_1, 
      u1_u14_X_10, u1_u14_X_15, u1_u14_X_16, u1_u14_X_17, u1_u14_X_19, u1_u14_X_21, u1_u14_X_22, u1_u14_X_27, u1_u14_X_28, 
      u1_u14_X_3, u1_u14_X_33, u1_u14_X_34, u1_u14_X_39, u1_u14_X_4, u1_u14_X_40, u1_u14_X_45, u1_u14_X_46, u1_u14_X_47, 
      u1_u14_X_9, u1_u15_X_15, u1_u15_X_16, u1_u15_X_21, u1_u15_X_22, u1_u15_X_23, u1_u15_X_24, u1_u15_X_25, u1_u15_X_26, 
      u1_u15_X_27, u1_u15_X_28, u1_u15_X_33, u1_u15_X_36, u1_u1_X_21, u1_u1_X_22, u1_u1_X_27, u1_u1_X_28, u1_u1_X_37, 
      u1_u1_X_38, u1_u1_X_39, u1_u1_X_40, u1_u1_X_45, u1_u1_X_46, u1_u2_X_3, u1_u2_X_39, u1_u2_X_4, u1_u2_X_40, 
      u1_u2_X_45, u1_u2_X_46, u1_u3_X_4, u1_u3_X_5, u1_u3_X_7, u1_u3_X_9, u1_u4_X_21, u1_u5_X_27, u1_u5_X_28, 
      u1_u5_X_33, u1_u5_X_34, u1_u6_X_10, u1_u6_X_15, u1_u6_X_16, u1_u6_X_3, u1_u6_X_39, u1_u6_X_4, u1_u6_X_40, 
      u1_u6_X_45, u1_u6_X_9, u1_u8_X_21, u1_u8_X_28, u1_u8_X_3, u1_u8_X_30, u1_u8_X_32, u1_u8_X_33, u1_u8_X_34, 
      u1_u8_X_39, u1_u8_X_4, u1_u8_X_40, u1_u8_X_45, u1_u8_X_46, u1_u9_X_34, u1_u9_X_39, u1_u9_X_40, u1_u9_X_45, 
      u1_u9_X_46, u1_uk_n1015, u1_uk_n1025, u1_uk_n1031, u1_uk_n1050, u1_uk_n1061, u1_uk_n1065, u1_uk_n1070, u1_uk_n1073, 
      u1_uk_n1074, u1_uk_n1105, u1_uk_n1106, u1_uk_n1123, u1_uk_n1124, u1_uk_n1125, u1_uk_n1126, u1_uk_n1154, u1_uk_n1155, 
      u1_uk_n1156, u1_uk_n1157, u1_uk_n1158, u1_uk_n1159, u1_uk_n1160, u1_uk_n1163, u1_uk_n1166, u1_uk_n1167, u1_uk_n1170, 
      u1_uk_n349, u1_uk_n353, u1_uk_n366, u1_uk_n369, u1_uk_n379, u1_uk_n382, u1_uk_n385, u1_uk_n437, u1_uk_n443, 
      u1_uk_n454, u1_uk_n496, u1_uk_n672, u1_uk_n676, u1_uk_n677, u1_uk_n678, u1_uk_n685, u1_uk_n702, u1_uk_n948, 
      u1_uk_n949, u1_uk_n950, u1_uk_n969, u1_uk_n970, u1_uk_n973, u1_uk_n974, u1_uk_n976, u1_uk_n985, u1_uk_n988, 
      u2_FP_33, u2_FP_36, u2_FP_37, u2_FP_40, u2_FP_41, u2_FP_44, u2_FP_45, u2_FP_48, u2_FP_49, 
      u2_FP_52, u2_FP_53, u2_FP_55, u2_FP_56, u2_FP_57, u2_FP_60, u2_FP_61, u2_FP_64, u2_K11_11, 
      u2_K11_13, u2_K16_1, u2_K16_11, u2_K16_12, u2_K16_13, u2_K16_14, u2_K16_17, u2_K16_18, u2_K16_19, 
      u2_K16_2, u2_K16_20, u2_K16_23, u2_K16_24, u2_K16_25, u2_K16_26, u2_K16_30, u2_K16_31, u2_K16_32, 
      u2_K16_35, u2_K16_36, u2_K16_38, u2_K16_41, u2_K16_42, u2_K16_44, u2_K16_47, u2_K16_48, u2_K16_5, 
      u2_K16_6, u2_K16_7, u2_K16_8, u2_K8_1, u2_K8_11, u2_K8_13, u2_K8_14, u2_K8_17, u2_K8_18, 
      u2_K8_19, u2_K8_2, u2_K8_20, u2_K8_47, u2_K8_48, u2_K8_5, u2_K8_6, u2_K8_7, u2_K8_8, 
      u2_K9_36, u2_K9_37, u2_K9_38, u2_K9_43, u2_R6_1, u2_R6_12, u2_R6_13, u2_R6_2, u2_R6_28, 
      u2_R6_32, u2_R6_4, u2_R6_5, u2_R6_8, u2_R6_9, u2_R7_1, u2_R7_22, u2_R7_24, u2_R7_25, 
      u2_R7_28, u2_R7_29, u2_R9_12, u2_R9_8, u2_R9_9, u2_u10_X_10, u2_u10_X_15, u2_u10_X_16, u2_u10_X_18, 
      u2_u10_X_7, u2_u10_X_8, u2_u10_X_9, u2_u15_X_10, u2_u15_X_15, u2_u15_X_16, u2_u15_X_21, u2_u15_X_22, u2_u15_X_27, 
      u2_u15_X_28, u2_u15_X_3, u2_u15_X_33, u2_u15_X_39, u2_u15_X_4, u2_u15_X_40, u2_u15_X_45, u2_u15_X_46, u2_u15_X_9, 
      u2_u7_X_10, u2_u7_X_15, u2_u7_X_16, u2_u7_X_21, u2_u7_X_22, u2_u7_X_23, u2_u7_X_24, u2_u7_X_4, u2_u7_X_44, 
      u2_u7_X_45, u2_u7_X_46, u2_u7_X_9, u2_u8_X_31, u2_u8_X_32, u2_u8_X_34, u2_u8_X_39, u2_u8_X_40, u2_u8_X_45, 
      u2_u8_X_46, u2_u8_X_47, u2_uk_K_r7_0, u2_uk_n1098, u2_uk_n1110, u2_uk_n1113, u2_uk_n1132, u2_uk_n1133, u2_uk_n1136, 
      u2_uk_n1137, u2_uk_n1140, u2_uk_n155, u2_uk_n1585, u2_uk_n214, u2_uk_n313, u2_uk_n319, u2_uk_n335, u2_uk_n955, 
      u2_uk_n958, u2_uk_n959, u2_uk_n963, u0_out0_1, u0_out0_10, u0_out0_13, u0_out0_16, u0_out0_17, u0_out0_18, 
      u0_out0_2, u0_out0_20, u0_out0_23, u0_out0_24, u0_out0_26, u0_out0_28, u0_out0_30, u0_out0_31, u0_out0_6, 
      u0_out0_9, u0_out10_1, u0_out10_10, u0_out10_13, u0_out10_16, u0_out10_18, u0_out10_2, u0_out10_20, u0_out10_24, 
      u0_out10_26, u0_out10_28, u0_out10_30, u0_out10_6, u0_out11_1, u0_out11_10, u0_out11_11, u0_out11_12, u0_out11_16, 
      u0_out11_19, u0_out11_20, u0_out11_22, u0_out11_24, u0_out11_26, u0_out11_29, u0_out11_30, u0_out11_32, u0_out11_4, 
      u0_out11_6, u0_out11_7, u0_out12_1, u0_out12_10, u0_out12_12, u0_out12_13, u0_out12_15, u0_out12_16, u0_out12_17, 
      u0_out12_18, u0_out12_2, u0_out12_20, u0_out12_21, u0_out12_22, u0_out12_23, u0_out12_24, u0_out12_26, u0_out12_27, 
      u0_out12_28, u0_out12_30, u0_out12_31, u0_out12_32, u0_out12_5, u0_out12_6, u0_out12_7, u0_out12_9, u0_out13_15, 
      u0_out13_21, u0_out13_27, u0_out13_5, u0_out14_1, u0_out14_10, u0_out14_13, u0_out14_16, u0_out14_18, u0_out14_2, 
      u0_out14_20, u0_out14_24, u0_out14_26, u0_out14_28, u0_out14_30, u0_out14_6, u0_out15_12, u0_out15_22, u0_out15_32, 
      u0_out15_7, u0_out1_11, u0_out1_12, u0_out1_14, u0_out1_19, u0_out1_22, u0_out1_25, u0_out1_29, u0_out1_3, 
      u0_out1_32, u0_out1_4, u0_out1_7, u0_out1_8, u0_out2_13, u0_out2_16, u0_out2_17, u0_out2_18, u0_out2_2, 
      u0_out2_23, u0_out2_24, u0_out2_28, u0_out2_30, u0_out2_31, u0_out2_6, u0_out2_9, u0_out5_1, u0_out5_10, 
      u0_out5_11, u0_out5_12, u0_out5_13, u0_out5_14, u0_out5_15, u0_out5_16, u0_out5_17, u0_out5_18, u0_out5_19, 
      u0_out5_2, u0_out5_20, u0_out5_21, u0_out5_22, u0_out5_23, u0_out5_24, u0_out5_25, u0_out5_26, u0_out5_27, 
      u0_out5_28, u0_out5_29, u0_out5_3, u0_out5_30, u0_out5_31, u0_out5_32, u0_out5_4, u0_out5_5, u0_out5_6, 
      u0_out5_7, u0_out5_8, u0_out5_9, u0_uk_n10, u0_uk_n102, u0_uk_n11, u0_uk_n110, u0_uk_n117, u0_uk_n129, 
      u0_uk_n141, u0_uk_n142, u0_uk_n145, u0_uk_n147, u0_uk_n162, u0_uk_n163, u0_uk_n182, u0_uk_n202, u0_uk_n203, 
      u0_uk_n207, u0_uk_n208, u0_uk_n217, u0_uk_n220, u0_uk_n222, u0_uk_n231, u0_uk_n238, u0_uk_n242, u0_uk_n250, 
      u0_uk_n251, u0_uk_n252, u0_uk_n31, u0_uk_n60, u1_out0_11, u1_out0_12, u1_out0_13, u1_out0_15, u1_out0_17, 
      u1_out0_18, u1_out0_19, u1_out0_2, u1_out0_21, u1_out0_22, u1_out0_23, u1_out0_27, u1_out0_28, u1_out0_29, 
      u1_out0_31, u1_out0_32, u1_out0_4, u1_out0_5, u1_out0_7, u1_out0_9, u1_out10_11, u1_out10_12, u1_out10_13, 
      u1_out10_15, u1_out10_16, u1_out10_17, u1_out10_18, u1_out10_19, u1_out10_2, u1_out10_21, u1_out10_22, u1_out10_23, 
      u1_out10_24, u1_out10_27, u1_out10_28, u1_out10_29, u1_out10_30, u1_out10_31, u1_out10_32, u1_out10_4, u1_out10_5, 
      u1_out10_6, u1_out10_7, u1_out10_9, u1_out12_1, u1_out12_10, u1_out12_13, u1_out12_15, u1_out12_16, u1_out12_17, 
      u1_out12_18, u1_out12_2, u1_out12_20, u1_out12_21, u1_out12_23, u1_out12_24, u1_out12_26, u1_out12_27, u1_out12_28, 
      u1_out12_30, u1_out12_31, u1_out12_5, u1_out12_6, u1_out12_9, u1_out13_12, u1_out13_13, u1_out13_15, u1_out13_17, 
      u1_out13_18, u1_out13_2, u1_out13_21, u1_out13_22, u1_out13_23, u1_out13_27, u1_out13_28, u1_out13_31, u1_out13_32, 
      u1_out13_5, u1_out13_7, u1_out13_9, u1_out14_1, u1_out14_10, u1_out14_11, u1_out14_12, u1_out14_13, u1_out14_14, 
      u1_out14_15, u1_out14_16, u1_out14_17, u1_out14_18, u1_out14_19, u1_out14_2, u1_out14_20, u1_out14_21, u1_out14_22, 
      u1_out14_23, u1_out14_24, u1_out14_25, u1_out14_26, u1_out14_27, u1_out14_28, u1_out14_29, u1_out14_3, u1_out14_30, 
      u1_out14_31, u1_out14_32, u1_out14_4, u1_out14_5, u1_out14_6, u1_out14_7, u1_out14_8, u1_out14_9, u1_out15_1, 
      u1_out15_10, u1_out15_11, u1_out15_14, u1_out15_16, u1_out15_19, u1_out15_20, u1_out15_24, u1_out15_25, u1_out15_26, 
      u1_out15_29, u1_out15_3, u1_out15_30, u1_out15_4, u1_out15_6, u1_out15_8, u1_out1_1, u1_out1_10, u1_out1_12, 
      u1_out1_14, u1_out1_15, u1_out1_20, u1_out1_21, u1_out1_22, u1_out1_25, u1_out1_26, u1_out1_27, u1_out1_3, 
      u1_out1_32, u1_out1_5, u1_out1_7, u1_out1_8, u1_out2_12, u1_out2_15, u1_out2_17, u1_out2_21, u1_out2_22, 
      u1_out2_23, u1_out2_27, u1_out2_31, u1_out2_32, u1_out2_5, u1_out2_7, u1_out2_9, u1_out3_13, u1_out3_17, 
      u1_out3_18, u1_out3_2, u1_out3_23, u1_out3_28, u1_out3_31, u1_out3_9, u1_out4_1, u1_out4_10, u1_out4_20, 
      u1_out4_26, u1_out5_11, u1_out5_14, u1_out5_19, u1_out5_25, u1_out5_29, u1_out5_3, u1_out5_4, u1_out5_8, 
      u1_out6_12, u1_out6_13, u1_out6_15, u1_out6_16, u1_out6_17, u1_out6_18, u1_out6_2, u1_out6_21, u1_out6_22, 
      u1_out6_23, u1_out6_24, u1_out6_27, u1_out6_28, u1_out6_30, u1_out6_31, u1_out6_32, u1_out6_5, u1_out6_6, 
      u1_out6_7, u1_out6_9, u1_out8_1, u1_out8_10, u1_out8_11, u1_out8_12, u1_out8_14, u1_out8_15, u1_out8_17, 
      u1_out8_19, u1_out8_20, u1_out8_21, u1_out8_22, u1_out8_23, u1_out8_25, u1_out8_26, u1_out8_27, u1_out8_29, 
      u1_out8_3, u1_out8_31, u1_out8_32, u1_out8_4, u1_out8_5, u1_out8_7, u1_out8_8, u1_out8_9, u1_out9_11, 
      u1_out9_12, u1_out9_15, u1_out9_19, u1_out9_21, u1_out9_22, u1_out9_27, u1_out9_29, u1_out9_32, u1_out9_4, 
      u1_out9_5, u1_out9_7, u2_out10_13, u2_out10_16, u2_out10_18, u2_out10_2, u2_out10_24, u2_out10_28, u2_out10_30, 
      u2_out10_6, u2_out15_1, u2_out15_10, u2_out15_11, u2_out15_12, u2_out15_13, u2_out15_14, u2_out15_15, u2_out15_16, 
      u2_out15_17, u2_out15_18, u2_out15_19, u2_out15_2, u2_out15_20, u2_out15_21, u2_out15_22, u2_out15_23, u2_out15_24, 
      u2_out15_25, u2_out15_26, u2_out15_27, u2_out15_28, u2_out15_29, u2_out15_3, u2_out15_30, u2_out15_31, u2_out15_32, 
      u2_out15_4, u2_out15_5, u2_out15_6, u2_out15_7, u2_out15_8, u2_out15_9, u2_out7_1, u2_out7_10, u2_out7_13, 
      u2_out7_15, u2_out7_16, u2_out7_17, u2_out7_18, u2_out7_2, u2_out7_20, u2_out7_21, u2_out7_23, u2_out7_24, 
      u2_out7_26, u2_out7_27, u2_out7_28, u2_out7_30, u2_out7_31, u2_out7_5, u2_out7_6, u2_out7_9, u2_out8_11, 
      u2_out8_12, u2_out8_15, u2_out8_19, u2_out8_21, u2_out8_22, u2_out8_27, u2_out8_29, u2_out8_32, u2_out8_4, 
      u2_out8_5, u2_out8_7 );
endmodule
