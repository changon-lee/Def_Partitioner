module aes_aes_die_10 ( sa30_6, sa30_7, us30_n441, us30_n447, us30_n448, us30_n449, us30_n452, us30_n460, us30_n465, 
       us30_n697, us30_n730, us30_n744, us30_n747, us30_n750, us30_n762, us30_n779, us30_n785, us30_n788, 
       us30_n790, us30_n803, us30_n806, us30_n813, us30_n814, us30_n816, us30_n817, sa31_sr_0, sa31_sr_1, sa31_sr_2, sa31_sr_3, sa31_sr_4, sa31_sr_5, sa31_sr_6, sa31_sr_7 );
  input sa30_6, sa30_7, us30_n441, us30_n447, us30_n448, us30_n449, us30_n452, us30_n460, us30_n465, 
        us30_n697, us30_n730, us30_n744, us30_n747, us30_n750, us30_n762, us30_n779, us30_n785, us30_n788, 
        us30_n790, us30_n803, us30_n806, us30_n813, us30_n814, us30_n816, us30_n817;
  output sa31_sr_0, sa31_sr_1, sa31_sr_2, sa31_sr_3, sa31_sr_4, sa31_sr_5, sa31_sr_6, sa31_sr_7;
  wire us30_n438, us30_n439, us30_n440, us30_n442, us30_n443, us30_n444, us30_n445, us30_n446, us30_n450, 
       us30_n456, us30_n457, us30_n458, us30_n459, us30_n463, us30_n464, us30_n466, us30_n467, us30_n468, 
       us30_n469, us30_n470, us30_n473, us30_n474, us30_n475, us30_n476, us30_n477, us30_n478, us30_n479, 
       us30_n480, us30_n481, us30_n482, us30_n483, us30_n484, us30_n485, us30_n486, us30_n487, us30_n488, 
       us30_n489, us30_n490, us30_n491, us30_n492, us30_n493, us30_n494, us30_n495, us30_n496, us30_n497, 
       us30_n498, us30_n499, us30_n500, us30_n501, us30_n502, us30_n503, us30_n504, us30_n505, us30_n506, 
       us30_n507, us30_n508, us30_n509, us30_n510, us30_n511, us30_n512, us30_n513, us30_n514, us30_n515, 
       us30_n516, us30_n517, us30_n518, us30_n519, us30_n520, us30_n521, us30_n522, us30_n523, us30_n524, 
       us30_n525, us30_n526, us30_n527, us30_n528, us30_n529, us30_n530, us30_n531, us30_n532, us30_n533, 
       us30_n534, us30_n535, us30_n536, us30_n537, us30_n538, us30_n539, us30_n540, us30_n541, us30_n542, 
       us30_n543, us30_n544, us30_n545, us30_n546, us30_n547, us30_n548, us30_n549, us30_n550, us30_n551, 
       us30_n552, us30_n553, us30_n554, us30_n555, us30_n556, us30_n557, us30_n558, us30_n559, us30_n560, 
       us30_n561, us30_n562, us30_n563, us30_n564, us30_n565, us30_n566, us30_n567, us30_n568, us30_n569, 
       us30_n570, us30_n571, us30_n572, us30_n573, us30_n574, us30_n575, us30_n576, us30_n577, us30_n578, 
       us30_n579, us30_n580, us30_n581, us30_n582, us30_n583, us30_n584, us30_n585, us30_n586, us30_n587, 
       us30_n588, us30_n589, us30_n590, us30_n591, us30_n592, us30_n593, us30_n594, us30_n595, us30_n596, 
       us30_n597, us30_n598, us30_n599, us30_n600, us30_n601, us30_n602, us30_n603, us30_n604, us30_n605, 
       us30_n606, us30_n607, us30_n608, us30_n609, us30_n610, us30_n611, us30_n612, us30_n613, us30_n614, 
       us30_n615, us30_n616, us30_n617, us30_n618, us30_n619, us30_n620, us30_n621, us30_n622, us30_n623, 
       us30_n624, us30_n625, us30_n626, us30_n627, us30_n628, us30_n629, us30_n630, us30_n631, us30_n632, 
       us30_n633, us30_n634, us30_n635, us30_n636, us30_n637, us30_n638, us30_n639, us30_n640, us30_n641, 
       us30_n642, us30_n643, us30_n644, us30_n645, us30_n646, us30_n647, us30_n648, us30_n649, us30_n650, 
       us30_n651, us30_n652, us30_n653, us30_n654, us30_n655, us30_n656, us30_n657, us30_n658, us30_n659, 
       us30_n660, us30_n661, us30_n662, us30_n663, us30_n664, us30_n665, us30_n666, us30_n667, us30_n668, 
       us30_n669, us30_n670, us30_n671, us30_n672, us30_n673, us30_n674, us30_n675, us30_n676, us30_n677, 
       us30_n678, us30_n679, us30_n680, us30_n681, us30_n682, us30_n683, us30_n684, us30_n685, us30_n686, 
       us30_n687, us30_n688, us30_n689, us30_n690, us30_n691, us30_n692, us30_n693, us30_n694, us30_n695, 
       us30_n696, us30_n698, us30_n699, us30_n700, us30_n701, us30_n702, us30_n703, us30_n704, us30_n705, 
       us30_n706, us30_n707, us30_n708, us30_n709, us30_n710, us30_n711, us30_n712, us30_n713, us30_n714, 
       us30_n715, us30_n716, us30_n717, us30_n718, us30_n719, us30_n720, us30_n721, us30_n722, us30_n723, 
       us30_n724, us30_n725, us30_n726, us30_n727, us30_n728, us30_n729, us30_n731, us30_n732, us30_n733, 
       us30_n734, us30_n735, us30_n736, us30_n737, us30_n738, us30_n739, us30_n740, us30_n741, us30_n742, 
       us30_n743, us30_n745, us30_n746, us30_n748, us30_n749, us30_n751, us30_n752, us30_n753, us30_n754, 
       us30_n755, us30_n756, us30_n757, us30_n758, us30_n759, us30_n760, us30_n761, us30_n763, us30_n764, 
       us30_n765, us30_n766, us30_n767, us30_n768, us30_n769, us30_n770, us30_n771, us30_n772, us30_n773, 
       us30_n774, us30_n775, us30_n776, us30_n777, us30_n778, us30_n780, us30_n781, us30_n782, us30_n783, 
       us30_n784, us30_n786, us30_n787, us30_n789, us30_n791, us30_n792, us30_n793, us30_n794, us30_n795, 
       us30_n796, us30_n797, us30_n798, us30_n799, us30_n800, us30_n801, us30_n802, us30_n804, us30_n805, 
       us30_n807, us30_n808, us30_n809, us30_n810, us30_n811, us30_n812, us30_n815, us30_n818, us30_n819, 
       us30_n820, us30_n821, us30_n822, us30_n823, us30_n824, us30_n825, us30_n830, us30_n831, us30_n832, 
       us30_n833, us30_n834, us30_n835, us30_n836, us30_n837, us30_n838, us30_n839, us30_n840, us30_n841, 
       us30_n842, us30_n843, us30_n844, us30_n845, us30_n846, us30_n850, us30_n851, us30_n852, us30_n853, 
       us30_n854, us30_n855, us30_n856, us30_n857, us30_n859, us30_n860, us30_n861, us30_n862, us30_n863, 
       us30_n864, us30_n865, us30_n866, us30_n867, us30_n868, us30_n869, us30_n870, us30_n871, us30_n872, 
       us30_n873, us30_n874, us30_n875,  us30_n876;
  NOR2_X1 us30_U10 (.ZN( us30_n575 ) , .A1( us30_n622 ) , .A2( us30_n745 ) );
  NOR2_X1 us30_U100 (.ZN( us30_n647 ) , .A1( us30_n854 ) , .A2( us30_n868 ) );
  NAND4_X1 us30_U101 (.A4( us30_n479 ) , .A3( us30_n480 ) , .A2( us30_n481 ) , .A1( us30_n482 ) , .ZN( us30_n694 ) );
  NOR3_X1 us30_U102 (.ZN( us30_n480 ) , .A2( us30_n508 ) , .A3( us30_n601 ) , .A1( us30_n610 ) );
  AOI211_X1 us30_U103 (.B( us30_n477 ) , .A( us30_n478 ) , .ZN( us30_n482 ) , .C2( us30_n833 ) , .C1( us30_n861 ) );
  NOR4_X1 us30_U104 (.ZN( us30_n481 ) , .A3( us30_n532 ) , .A4( us30_n545 ) , .A2( us30_n567 ) , .A1( us30_n717 ) );
  NAND4_X1 us30_U105 (.A4( us30_n548 ) , .A3( us30_n549 ) , .A2( us30_n550 ) , .A1( us30_n551 ) , .ZN( us30_n745 ) );
  NOR3_X1 us30_U106 (.ZN( us30_n549 ) , .A2( us30_n651 ) , .A1( us30_n667 ) , .A3( us30_n771 ) );
  AOI211_X1 us30_U107 (.B( us30_n539 ) , .A( us30_n540 ) , .ZN( us30_n551 ) , .C2( us30_n839 ) , .C1( us30_n851 ) );
  NOR4_X1 us30_U108 (.A4( us30_n544 ) , .A3( us30_n545 ) , .A2( us30_n546 ) , .A1( us30_n547 ) , .ZN( us30_n548 ) );
  NOR4_X1 us30_U109 (.ZN( us30_n620 ) , .A1( us30_n656 ) , .A3( us30_n666 ) , .A4( us30_n682 ) , .A2( us30_n766 ) );
  NOR2_X1 us30_U11 (.ZN( us30_n495 ) , .A1( us30_n678 ) , .A2( us30_n694 ) );
  NOR4_X1 us30_U110 (.A4( us30_n609 ) , .A3( us30_n610 ) , .A2( us30_n611 ) , .A1( us30_n612 ) , .ZN( us30_n619 ) );
  NOR4_X1 us30_U111 (.A4( us30_n614 ) , .A3( us30_n615 ) , .A2( us30_n616 ) , .A1( us30_n617 ) , .ZN( us30_n618 ) );
  NOR2_X1 us30_U112 (.ZN( us30_n686 ) , .A1( us30_n831 ) , .A2( us30_n832 ) );
  NAND4_X1 us30_U113 (.A4( us30_n485 ) , .A3( us30_n486 ) , .A2( us30_n487 ) , .A1( us30_n488 ) , .ZN( us30_n778 ) );
  NOR4_X1 us30_U114 (.A4( us30_n484 ) , .ZN( us30_n487 ) , .A1( us30_n566 ) , .A2( us30_n581 ) , .A3( us30_n602 ) );
  NOR4_X1 us30_U115 (.ZN( us30_n486 ) , .A1( us30_n507 ) , .A2( us30_n519 ) , .A4( us30_n546 ) , .A3( us30_n611 ) );
  NOR4_X1 us30_U116 (.ZN( us30_n485 ) , .A2( us30_n533 ) , .A1( us30_n558 ) , .A3( us30_n631 ) , .A4( us30_n718 ) );
  NAND4_X1 us30_U117 (.A4( us30_n691 ) , .A3( us30_n692 ) , .A1( us30_n693 ) , .ZN( us30_n776 ) , .A2( us30_n872 ) );
  AOI221_X1 us30_U118 (.A( us30_n681 ) , .ZN( us30_n692 ) , .B2( us30_n840 ) , .C1( us30_n842 ) , .C2( us30_n862 ) , .B1( us30_n865 ) );
  INV_X1 us30_U119 (.A( us30_n679 ) , .ZN( us30_n872 ) );
  NOR2_X1 us30_U12 (.A1( us30_n678 ) , .ZN( us30_n693 ) , .A2( us30_n807 ) );
  NOR4_X1 us30_U120 (.A4( us30_n687 ) , .A3( us30_n688 ) , .A2( us30_n689 ) , .A1( us30_n690 ) , .ZN( us30_n691 ) );
  NAND4_X1 us30_U121 (.A4( us30_n719 ) , .A3( us30_n720 ) , .A2( us30_n721 ) , .ZN( us30_n741 ) , .A1( us30_n857 ) );
  INV_X1 us30_U122 (.A( us30_n709 ) , .ZN( us30_n857 ) );
  AOI221_X1 us30_U123 (.A( us30_n710 ) , .ZN( us30_n721 ) , .C2( us30_n844 ) , .B2( us30_n845 ) , .C1( us30_n861 ) , .B1( us30_n862 ) );
  NOR4_X1 us30_U124 (.A4( us30_n715 ) , .A3( us30_n716 ) , .A2( us30_n717 ) , .A1( us30_n718 ) , .ZN( us30_n719 ) );
  NAND4_X1 us30_U125 (.A4( us30_n473 ) , .A3( us30_n474 ) , .A2( us30_n475 ) , .A1( us30_n476 ) , .ZN( us30_n678 ) );
  NOR4_X1 us30_U126 (.ZN( us30_n475 ) , .A1( us30_n531 ) , .A3( us30_n568 ) , .A4( us30_n600 ) , .A2( us30_n642 ) );
  NOR4_X1 us30_U127 (.A4( us30_n470 ) , .ZN( us30_n476 ) , .A3( us30_n556 ) , .A1( us30_n735 ) , .A2( us30_n755 ) );
  NOR4_X1 us30_U128 (.ZN( us30_n474 ) , .A1( us30_n506 ) , .A3( us30_n544 ) , .A2( us30_n583 ) , .A4( us30_n716 ) );
  NOR2_X1 us30_U129 (.ZN( us30_n733 ) , .A2( us30_n832 ) , .A1( us30_n845 ) );
  NOR3_X1 us30_U13 (.ZN( us30_n504 ) , .A2( us30_n679 ) , .A3( us30_n777 ) , .A1( us30_n876 ) );
  NOR2_X1 us30_U130 (.ZN( us30_n789 ) , .A2( us30_n862 ) , .A1( us30_n868 ) );
  NAND4_X1 us30_U131 (.A4( us30_n573 ) , .A3( us30_n574 ) , .A1( us30_n575 ) , .ZN( us30_n723 ) , .A2( us30_n874 ) );
  AOI221_X1 us30_U132 (.A( us30_n564 ) , .C2( us30_n565 ) , .ZN( us30_n574 ) , .B2( us30_n845 ) , .B1( us30_n852 ) , .C1( us30_n853 ) );
  NOR4_X1 us30_U133 (.A4( us30_n569 ) , .A3( us30_n570 ) , .A2( us30_n571 ) , .A1( us30_n572 ) , .ZN( us30_n573 ) );
  INV_X1 us30_U134 (.A( us30_n607 ) , .ZN( us30_n874 ) );
  NAND4_X1 us30_U135 (.A4( us30_n633 ) , .A3( us30_n634 ) , .A2( us30_n635 ) , .A1( us30_n636 ) , .ZN( us30_n743 ) );
  AOI211_X1 us30_U136 (.B( us30_n623 ) , .A( us30_n624 ) , .ZN( us30_n635 ) , .C2( us30_n836 ) , .C1( us30_n863 ) );
  NOR4_X1 us30_U137 (.A4( us30_n629 ) , .A3( us30_n630 ) , .A2( us30_n631 ) , .A1( us30_n632 ) , .ZN( us30_n633 ) );
  NOR4_X1 us30_U138 (.A4( us30_n626 ) , .A3( us30_n627 ) , .A2( us30_n628 ) , .ZN( us30_n634 ) , .A1( us30_n664 ) );
  NAND4_X1 us30_U139 (.A4( us30_n493 ) , .A3( us30_n494 ) , .A1( us30_n495 ) , .ZN( us30_n802 ) , .A2( us30_n867 ) );
  INV_X1 us30_U14 (.A( us30_n706 ) , .ZN( us30_n876 ) );
  AOI221_X1 us30_U140 (.A( us30_n489 ) , .ZN( us30_n494 ) , .B2( us30_n836 ) , .C2( us30_n841 ) , .C1( us30_n851 ) , .B1( us30_n860 ) );
  INV_X1 us30_U141 (.A( us30_n778 ) , .ZN( us30_n867 ) );
  NOR4_X1 us30_U142 (.A2( us30_n491 ) , .A1( us30_n492 ) , .ZN( us30_n493 ) , .A3( us30_n580 ) , .A4( us30_n612 ) );
  NOR4_X1 us30_U143 (.A4( us30_n734 ) , .A3( us30_n735 ) , .A2( us30_n736 ) , .A1( us30_n737 ) , .ZN( us30_n738 ) );
  AOI211_X1 us30_U144 (.B( us30_n725 ) , .A( us30_n726 ) , .ZN( us30_n739 ) , .C1( us30_n843 ) , .C2( us30_n855 ) );
  NOR3_X1 us30_U145 (.A3( us30_n722 ) , .A1( us30_n723 ) , .ZN( us30_n740 ) , .A2( us30_n741 ) );
  INV_X1 us30_U146 (.A( us30_n762 ) , .ZN( us30_n830 ) );
  OR4_X1 us30_U147 (.A4( us30_n566 ) , .A3( us30_n567 ) , .A2( us30_n568 ) , .ZN( us30_n572 ) , .A1( us30_n665 ) );
  OR4_X1 us30_U148 (.A4( us30_n682 ) , .A3( us30_n683 ) , .A2( us30_n684 ) , .A1( us30_n685 ) , .ZN( us30_n690 ) );
  OR4_X1 us30_U149 (.ZN( us30_n466 ) , .A4( us30_n518 ) , .A3( us30_n529 ) , .A2( us30_n578 ) , .A1( us30_n712 ) );
  INV_X1 us30_U15 (.A( us30_n680 ) , .ZN( us30_n840 ) );
  OR4_X1 us30_U150 (.A4( us30_n518 ) , .A2( us30_n519 ) , .A1( us30_n520 ) , .ZN( us30_n522 ) , .A3( us30_n821 ) );
  OR4_X1 us30_U151 (.ZN( us30_n492 ) , .A4( us30_n534 ) , .A2( us30_n547 ) , .A1( us30_n559 ) , .A3( us30_n632 ) );
  OR4_X1 us30_U152 (.A4( us30_n580 ) , .A3( us30_n581 ) , .A2( us30_n582 ) , .A1( us30_n583 ) , .ZN( us30_n584 ) );
  INV_X1 us30_U153 (.A( us30_n697 ) , .ZN( us30_n838 ) );
  NAND2_X1 us30_U154 (.ZN( us30_n613 ) , .A2( us30_n837 ) , .A1( us30_n873 ) );
  OR3_X1 us30_U155 (.A3( us30_n506 ) , .A2( us30_n507 ) , .A1( us30_n508 ) , .ZN( us30_n511 ) );
  INV_X1 us30_U156 (.A( us30_n754 ) , .ZN( us30_n869 ) );
  OAI21_X1 us30_U157 (.B1( us30_n753 ) , .ZN( us30_n754 ) , .A( us30_n845 ) , .B2( us30_n868 ) );
  INV_X1 us30_U158 (.A( us30_n463 ) , .ZN( us30_n864 ) );
  OAI21_X1 us30_U159 (.ZN( us30_n463 ) , .B1( us30_n809 ) , .A( us30_n834 ) , .B2( us30_n851 ) );
  NOR4_X1 us30_U16 (.A4( us30_n445 ) , .A3( us30_n446 ) , .A2( us30_n516 ) , .A1( us30_n541 ) , .ZN( us30_n706 ) );
  INV_X1 us30_U160 (.A( us30_n672 ) , .ZN( us30_n859 ) );
  AOI21_X1 us30_U161 (.A( us30_n670 ) , .B1( us30_n671 ) , .ZN( us30_n672 ) , .B2( us30_n856 ) );
  OAI222_X1 us30_U162 (.B2( us30_n747 ) , .B1( us30_n748 ) , .A2( us30_n749 ) , .ZN( us30_n757 ) , .C2( us30_n805 ) , .C1( us30_n814 ) , .A1( us30_n817 ) );
  OAI222_X1 us30_U163 (.ZN( us30_n505 ) , .C2( us30_n625 ) , .B2( us30_n647 ) , .B1( us30_n747 ) , .A2( us30_n748 ) , .C1( us30_n805 ) , .A1( us30_n806 ) );
  OAI222_X1 us30_U164 (.B2( us30_n708 ) , .ZN( us30_n709 ) , .C2( us30_n724 ) , .B1( us30_n747 ) , .A1( us30_n806 ) , .C1( us30_n814 ) , .A2( us30_n815 ) );
  NAND2_X1 us30_U165 (.A1( us30_n447 ) , .A2( us30_n465 ) , .ZN( us30_n749 ) );
  AOI22_X1 us30_U166 (.ZN( us30_n696 ) , .A1( us30_n830 ) , .B2( us30_n843 ) , .A2( us30_n865 ) , .B1( us30_n868 ) );
  AOI22_X1 us30_U167 (.A2( us30_n782 ) , .ZN( us30_n783 ) , .B2( us30_n831 ) , .A1( us30_n834 ) , .B1( us30_n863 ) );
  INV_X1 us30_U168 (.A( us30_n730 ) , .ZN( us30_n839 ) );
  AOI221_X1 us30_U169 (.A( us30_n764 ) , .ZN( us30_n774 ) , .C2( us30_n810 ) , .B2( us30_n835 ) , .C1( us30_n855 ) , .B1( us30_n866 ) );
  OR3_X1 us30_U17 (.ZN( us30_n446 ) , .A1( us30_n528 ) , .A3( us30_n577 ) , .A2( us30_n875 ) );
  AOI21_X1 us30_U170 (.B2( us30_n763 ) , .ZN( us30_n764 ) , .A( us30_n788 ) , .B1( us30_n792 ) );
  INV_X1 us30_U171 (.A( us30_n761 ) , .ZN( us30_n835 ) );
  AOI221_X1 us30_U172 (.A( us30_n483 ) , .ZN( us30_n488 ) , .B1( us30_n831 ) , .C2( us30_n844 ) , .C1( us30_n852 ) , .B2( us30_n862 ) );
  OAI22_X1 us30_U173 (.ZN( us30_n483 ) , .A1( us30_n708 ) , .B2( us30_n785 ) , .A2( us30_n806 ) , .B1( us30_n812 ) );
  INV_X1 us30_U174 (.A( us30_n790 ) , .ZN( us30_n832 ) );
  OAI221_X1 us30_U176 (.A( us30_n727 ) , .C2( us30_n728 ) , .B2( us30_n729 ) , .B1( us30_n730 ) , .ZN( us30_n737 ) , .C1( us30_n817 ) );
  AOI22_X1 us30_U177 (.ZN( us30_n727 ) , .B1( us30_n832 ) , .A2( us30_n838 ) , .A1( us30_n863 ) , .B2( us30_n866 ) );
  INV_X1 us30_U178 (.A( us30_n786 ) , .ZN( us30_n862 ) );
  OAI22_X1 us30_U179 (.ZN( us30_n710 ) , .A2( us30_n728 ) , .B2( us30_n729 ) , .A1( us30_n744 ) , .B1( us30_n813 ) );
  OR4_X1 us30_U18 (.A4( us30_n442 ) , .A2( us30_n443 ) , .A1( us30_n444 ) , .ZN( us30_n445 ) , .A3( us30_n553 ) );
  INV_X1 us30_U180 (.A( us30_n816 ) , .ZN( us30_n831 ) );
  OAI22_X1 us30_U181 (.ZN( us30_n489 ) , .A1( us30_n724 ) , .B2( us30_n728 ) , .B1( us30_n730 ) , .A2( us30_n779 ) );
  OAI22_X1 us30_U182 (.ZN( us30_n624 ) , .B1( us30_n669 ) , .B2( us30_n747 ) , .A1( us30_n815 ) , .A2( us30_n816 ) );
  INV_X1 us30_U183 (.A( us30_n744 ) , .ZN( us30_n837 ) );
  INV_X1 us30_U184 (.A( us30_n788 ) , .ZN( us30_n845 ) );
  OAI22_X1 us30_U185 (.B2( us30_n779 ) , .B1( us30_n780 ) , .ZN( us30_n781 ) , .A2( us30_n814 ) , .A1( us30_n815 ) );
  OAI22_X1 us30_U186 (.A1( us30_n724 ) , .ZN( us30_n726 ) , .B2( us30_n750 ) , .B1( us30_n812 ) , .A2( us30_n816 ) );
  INV_X1 us30_U187 (.A( us30_n805 ) , .ZN( us30_n860 ) );
  INV_X1 us30_U188 (.A( us30_n814 ) , .ZN( us30_n833 ) );
  INV_X1 us30_U189 (.A( us30_n669 ) , .ZN( us30_n865 ) );
  INV_X1 us30_U19 (.A( us30_n613 ) , .ZN( us30_n875 ) );
  OAI22_X1 us30_U190 (.B2( us30_n744 ) , .ZN( us30_n746 ) , .A2( us30_n762 ) , .B1( us30_n780 ) , .A1( us30_n792 ) );
  OAI22_X1 us30_U191 (.ZN( us30_n496 ) , .A2( us30_n744 ) , .A1( us30_n780 ) , .B1( us30_n791 ) , .B2( us30_n806 ) );
  OAI22_X1 us30_U192 (.B2( us30_n803 ) , .B1( us30_n804 ) , .A2( us30_n805 ) , .A1( us30_n806 ) , .ZN( us30_n808 ) );
  AOI211_X1 us30_U193 (.A( us30_n637 ) , .ZN( us30_n645 ) , .B( us30_n743 ) , .C2( us30_n839 ) , .C1( us30_n854 ) );
  OAI22_X1 us30_U194 (.ZN( us30_n637 ) , .A1( us30_n699 ) , .B2( us30_n728 ) , .A2( us30_n762 ) , .B1( us30_n816 ) );
  OAI22_X1 us30_U195 (.B1( us30_n490 ) , .ZN( us30_n491 ) , .A1( us30_n686 ) , .A2( us30_n763 ) , .B2( us30_n817 ) );
  NOR3_X1 us30_U196 (.ZN( us30_n490 ) , .A1( us30_n782 ) , .A2( us30_n850 ) , .A3( us30_n863 ) );
  INV_X1 us30_U197 (.A( us30_n750 ) , .ZN( us30_n842 ) );
  OAI22_X1 us30_U198 (.ZN( us30_n695 ) , .A2( us30_n730 ) , .A1( us30_n780 ) , .B1( us30_n791 ) , .B2( us30_n817 ) );
  NOR2_X1 us30_U199 (.ZN( us30_n715 ) , .A1( us30_n805 ) , .A2( us30_n817 ) );
  INV_X1 us30_U20 (.A( us30_n749 ) , .ZN( us30_n863 ) );
  NOR2_X1 us30_U200 (.ZN( us30_n666 ) , .A1( us30_n728 ) , .A2( us30_n803 ) );
  NOR2_X1 us30_U201 (.ZN( us30_n594 ) , .A2( us30_n697 ) , .A1( us30_n728 ) );
  NOR2_X1 us30_U202 (.ZN( us30_n570 ) , .A1( us30_n728 ) , .A2( us30_n806 ) );
  NOR2_X1 us30_U203 (.A2( us30_n744 ) , .ZN( us30_n755 ) , .A1( us30_n805 ) );
  NOR2_X1 us30_U204 (.ZN( us30_n735 ) , .A2( us30_n803 ) , .A1( us30_n805 ) );
  NOR2_X1 us30_U205 (.ZN( us30_n546 ) , .A2( us30_n780 ) , .A1( us30_n814 ) );
  NOR2_X1 us30_U206 (.ZN( us30_n577 ) , .A2( us30_n699 ) , .A1( us30_n814 ) );
  NOR2_X1 us30_U207 (.ZN( us30_n654 ) , .A1( us30_n728 ) , .A2( us30_n813 ) );
  NOR2_X1 us30_U208 (.ZN( us30_n718 ) , .A2( us30_n724 ) , .A1( us30_n744 ) );
  NOR2_X1 us30_U209 (.ZN( us30_n532 ) , .A2( us30_n749 ) , .A1( us30_n750 ) );
  AOI222_X1 us30_U21 (.ZN( us30_n605 ) , .B2( us30_n671 ) , .B1( us30_n753 ) , .C2( us30_n831 ) , .A1( us30_n833 ) , .A2( us30_n862 ) , .C1( us30_n863 ) );
  NOR2_X1 us30_U210 (.ZN( us30_n615 ) , .A1( us30_n785 ) , .A2( us30_n815 ) );
  NOR2_X1 us30_U211 (.ZN( us30_n629 ) , .A2( us30_n728 ) , .A1( us30_n785 ) );
  NOR2_X1 us30_U212 (.ZN( us30_n611 ) , .A2( us30_n780 ) , .A1( us30_n806 ) );
  NOR2_X1 us30_U213 (.ZN( us30_n628 ) , .A2( us30_n669 ) , .A1( us30_n785 ) );
  INV_X1 us30_U214 (.A( us30_n747 ) , .ZN( us30_n834 ) );
  INV_X1 us30_U215 (.A( us30_n728 ) , .ZN( us30_n852 ) );
  NOR2_X1 us30_U216 (.ZN( us30_n652 ) , .A1( us30_n669 ) , .A2( us30_n814 ) );
  NOR2_X1 us30_U217 (.A1( us30_n669 ) , .ZN( us30_n673 ) , .A2( us30_n744 ) );
  NOR2_X1 us30_U218 (.ZN( us30_n602 ) , .A1( us30_n669 ) , .A2( us30_n803 ) );
  NOR2_X1 us30_U219 (.A1( us30_n669 ) , .ZN( us30_n688 ) , .A2( us30_n816 ) );
  AOI222_X1 us30_U22 (.ZN( us30_n563 ) , .B1( us30_n830 ) , .C1( us30_n841 ) , .A2( us30_n843 ) , .A1( us30_n854 ) , .B2( us30_n863 ) , .C2( us30_n873 ) );
  NOR2_X1 us30_U220 (.A2( us30_n744 ) , .ZN( us30_n769 ) , .A1( us30_n812 ) );
  NOR2_X1 us30_U221 (.ZN( us30_n531 ) , .A2( us30_n780 ) , .A1( us30_n816 ) );
  INV_X1 us30_U222 (.A( us30_n792 ) , .ZN( us30_n851 ) );
  NOR2_X1 us30_U223 (.A2( us30_n708 ) , .A1( us30_n750 ) , .ZN( us30_n771 ) );
  NOR2_X1 us30_U224 (.ZN( us30_n599 ) , .A2( us30_n791 ) , .A1( us30_n816 ) );
  NOR2_X1 us30_U225 (.A1( us30_n669 ) , .ZN( us30_n766 ) , .A2( us30_n813 ) );
  NOR2_X1 us30_U226 (.ZN( us30_n601 ) , .A2( us30_n780 ) , .A1( us30_n803 ) );
  NOR2_X1 us30_U227 (.A1( us30_n699 ) , .ZN( us30_n768 ) , .A2( us30_n813 ) );
  NOR2_X1 us30_U228 (.ZN( us30_n541 ) , .A2( us30_n697 ) , .A1( us30_n699 ) );
  NOR2_X1 us30_U229 (.ZN( us30_n527 ) , .A1( us30_n669 ) , .A2( us30_n779 ) );
  AOI222_X1 us30_U23 (.ZN( us30_n660 ) , .A2( us30_n839 ) , .B1( us30_n841 ) , .C2( us30_n845 ) , .A1( us30_n860 ) , .C1( us30_n863 ) , .B2( us30_n870 ) );
  NOR2_X1 us30_U230 (.ZN( us30_n667 ) , .A1( us30_n750 ) , .A2( us30_n815 ) );
  NOR2_X1 us30_U231 (.ZN( us30_n555 ) , .A1( us30_n750 ) , .A2( us30_n791 ) );
  NOR2_X1 us30_U232 (.ZN( us30_n508 ) , .A2( us30_n780 ) , .A1( us30_n785 ) );
  NOR2_X1 us30_U233 (.ZN( us30_n543 ) , .A2( us30_n708 ) , .A1( us30_n785 ) );
  NOR2_X1 us30_U234 (.ZN( us30_n528 ) , .A2( us30_n724 ) , .A1( us30_n803 ) );
  NOR2_X1 us30_U235 (.ZN( us30_n664 ) , .A1( us30_n785 ) , .A2( us30_n791 ) );
  NOR2_X1 us30_U236 (.ZN( us30_n556 ) , .A1( us30_n762 ) , .A2( us30_n805 ) );
  INV_X1 us30_U237 (.A( us30_n806 ) , .ZN( us30_n841 ) );
  NOR2_X1 us30_U238 (.ZN( us30_n661 ) , .A1( us30_n729 ) , .A2( us30_n790 ) );
  OAI22_X1 us30_U239 (.B1( us30_n440 ) , .ZN( us30_n444 ) , .A2( us30_n728 ) , .A1( us30_n744 ) , .B2( us30_n749 ) );
  INV_X1 us30_U24 (.A( us30_n647 ) , .ZN( us30_n870 ) );
  NOR3_X1 us30_U240 (.ZN( us30_n440 ) , .A2( us30_n836 ) , .A3( us30_n837 ) , .A1( us30_n846 ) );
  NOR2_X1 us30_U241 (.ZN( us30_n507 ) , .A1( us30_n812 ) , .A2( us30_n817 ) );
  NOR2_X1 us30_U242 (.ZN( us30_n557 ) , .A1( us30_n792 ) , .A2( us30_n814 ) );
  NOR2_X1 us30_U243 (.ZN( us30_n545 ) , .A1( us30_n749 ) , .A2( us30_n814 ) );
  NOR2_X1 us30_U244 (.ZN( us30_n509 ) , .A1( us30_n729 ) , .A2( us30_n779 ) );
  NOR2_X1 us30_U245 (.ZN( us30_n662 ) , .A2( us30_n697 ) , .A1( us30_n729 ) );
  OAI22_X1 us30_U246 (.B2( us30_n750 ) , .B1( us30_n751 ) , .A1( us30_n752 ) , .ZN( us30_n756 ) , .A2( us30_n806 ) );
  NOR2_X1 us30_U247 (.ZN( us30_n751 ) , .A2( us30_n852 ) , .A1( us30_n860 ) );
  NOR3_X1 us30_U248 (.ZN( us30_n752 ) , .A2( us30_n853 ) , .A1( us30_n863 ) , .A3( us30_n865 ) );
  NOR2_X1 us30_U249 (.ZN( us30_n544 ) , .A2( us30_n785 ) , .A1( us30_n792 ) );
  NOR4_X1 us30_U25 (.ZN( us30_n473 ) , .A2( us30_n521 ) , .A4( us30_n594 ) , .A1( us30_n609 ) , .A3( us30_n629 ) );
  NOR2_X1 us30_U250 (.ZN( us30_n663 ) , .A1( us30_n729 ) , .A2( us30_n785 ) );
  NOR2_X1 us30_U251 (.ZN( us30_n530 ) , .A2( us30_n744 ) , .A1( us30_n792 ) );
  NOR2_X1 us30_U252 (.ZN( us30_n506 ) , .A2( us30_n728 ) , .A1( us30_n762 ) );
  NOR2_X1 us30_U253 (.ZN( us30_n631 ) , .A1( us30_n724 ) , .A2( us30_n813 ) );
  NOR2_X1 us30_U254 (.ZN( us30_n614 ) , .A1( us30_n762 ) , .A2( us30_n812 ) );
  NOR2_X1 us30_U255 (.A1( us30_n749 ) , .ZN( us30_n767 ) , .A2( us30_n803 ) );
  NOR2_X1 us30_U256 (.ZN( us30_n516 ) , .A1( us30_n708 ) , .A2( us30_n744 ) );
  NOR2_X1 us30_U257 (.ZN( us30_n670 ) , .A1( us30_n790 ) , .A2( us30_n805 ) );
  NOR2_X1 us30_U258 (.ZN( us30_n558 ) , .A1( us30_n708 ) , .A2( us30_n816 ) );
  NOR2_X1 us30_U259 (.A2( us30_n697 ) , .ZN( us30_n716 ) , .A1( us30_n792 ) );
  NOR4_X1 us30_U26 (.ZN( us30_n479 ) , .A1( us30_n520 ) , .A4( us30_n557 ) , .A3( us30_n582 ) , .A2( us30_n630 ) );
  NOR2_X1 us30_U260 (.ZN( us30_n517 ) , .A1( us30_n708 ) , .A2( us30_n803 ) );
  NOR2_X1 us30_U261 (.ZN( us30_n521 ) , .A1( us30_n790 ) , .A2( us30_n812 ) );
  NOR2_X1 us30_U262 (.ZN( us30_n630 ) , .A1( us30_n747 ) , .A2( us30_n815 ) );
  NOR2_X1 us30_U263 (.ZN( us30_n655 ) , .A1( us30_n790 ) , .A2( us30_n815 ) );
  INV_X1 us30_U264 (.A( us30_n763 ) , .ZN( us30_n866 ) );
  AOI21_X1 us30_U265 (.ZN( us30_n552 ) , .B1( us30_n669 ) , .A( us30_n697 ) , .B2( us30_n805 ) );
  NOR2_X1 us30_U266 (.ZN( us30_n668 ) , .A2( us30_n708 ) , .A1( us30_n790 ) );
  NOR2_X1 us30_U267 (.ZN( us30_n542 ) , .A1( us30_n762 ) , .A2( us30_n791 ) );
  NOR2_X1 us30_U268 (.ZN( us30_n656 ) , .A1( us30_n747 ) , .A2( us30_n780 ) );
  NOR2_X1 us30_U269 (.ZN( us30_n609 ) , .A2( us30_n724 ) , .A1( us30_n817 ) );
  NOR4_X1 us30_U27 (.A4( us30_n532 ) , .A3( us30_n533 ) , .A2( us30_n534 ) , .ZN( us30_n535 ) , .A1( us30_n820 ) );
  INV_X1 us30_U270 (.A( us30_n729 ) , .ZN( us30_n868 ) );
  AOI21_X1 us30_U271 (.B1( us30_n625 ) , .ZN( us30_n627 ) , .A( us30_n763 ) , .B2( us30_n814 ) );
  AOI21_X1 us30_U272 (.ZN( us30_n650 ) , .A( us30_n779 ) , .B1( us30_n792 ) , .B2( us30_n805 ) );
  AOI21_X1 us30_U273 (.A( us30_n815 ) , .B2( us30_n816 ) , .B1( us30_n817 ) , .ZN( us30_n818 ) );
  NOR2_X1 us30_U274 (.ZN( us30_n579 ) , .A2( us30_n708 ) , .A1( us30_n730 ) );
  NOR2_X1 us30_U275 (.ZN( us30_n533 ) , .A2( us30_n724 ) , .A1( us30_n730 ) );
  NOR2_X1 us30_U276 (.ZN( us30_n642 ) , .A2( us30_n788 ) , .A1( us30_n791 ) );
  AOI21_X1 us30_U277 (.A( us30_n812 ) , .B2( us30_n813 ) , .B1( us30_n814 ) , .ZN( us30_n819 ) );
  NOR2_X1 us30_U278 (.A2( us30_n708 ) , .A1( us30_n762 ) , .ZN( us30_n794 ) );
  NOR2_X1 us30_U279 (.A2( us30_n697 ) , .A1( us30_n780 ) , .ZN( us30_n820 ) );
  NOR4_X1 us30_U28 (.ZN( us30_n456 ) , .A2( us30_n517 ) , .A1( us30_n543 ) , .A3( us30_n579 ) , .A4( us30_n615 ) );
  AOI21_X1 us30_U280 (.ZN( us30_n626 ) , .B2( us30_n669 ) , .A( us30_n790 ) , .B1( us30_n791 ) );
  AOI21_X1 us30_U281 (.ZN( us30_n499 ) , .B1( us30_n680 ) , .A( us30_n812 ) , .B2( us30_n816 ) );
  NOR2_X1 us30_U282 (.ZN( us30_n520 ) , .A2( us30_n708 ) , .A1( us30_n814 ) );
  AOI21_X1 us30_U283 (.ZN( us30_n477 ) , .A( us30_n669 ) , .B1( us30_n750 ) , .B2( us30_n806 ) );
  NOR2_X1 us30_U284 (.ZN( us30_n582 ) , .A1( us30_n744 ) , .A2( us30_n815 ) );
  AOI21_X1 us30_U285 (.ZN( us30_n593 ) , .B1( us30_n750 ) , .A( us30_n792 ) , .B2( us30_n813 ) );
  AOI21_X1 us30_U286 (.ZN( us30_n515 ) , .A( us30_n729 ) , .B1( us30_n750 ) , .B2( us30_n803 ) );
  NOR2_X1 us30_U287 (.A1( us30_n697 ) , .ZN( us30_n770 ) , .A2( us30_n815 ) );
  AOI21_X1 us30_U288 (.ZN( us30_n510 ) , .B2( us30_n669 ) , .A( us30_n730 ) , .B1( us30_n815 ) );
  NOR2_X1 us30_U289 (.ZN( us30_n519 ) , .A2( us30_n699 ) , .A1( us30_n816 ) );
  NOR4_X1 us30_U29 (.A4( us30_n541 ) , .A3( us30_n542 ) , .A2( us30_n543 ) , .ZN( us30_n550 ) , .A1( us30_n688 ) );
  NOR2_X1 us30_U290 (.ZN( us30_n559 ) , .A2( us30_n791 ) , .A1( us30_n803 ) );
  NOR2_X1 us30_U291 (.ZN( us30_n581 ) , .A1( us30_n669 ) , .A2( us30_n788 ) );
  INV_X1 us30_U292 (.A( us30_n813 ) , .ZN( us30_n836 ) );
  NOR2_X1 us30_U293 (.ZN( us30_n683 ) , .A2( us30_n699 ) , .A1( us30_n803 ) );
  AOI21_X1 us30_U294 (.ZN( us30_n589 ) , .B2( us30_n699 ) , .B1( us30_n815 ) , .A( us30_n817 ) );
  AOI21_X1 us30_U295 (.ZN( us30_n539 ) , .B2( us30_n812 ) , .A( us30_n814 ) , .B1( us30_n815 ) );
  AOI21_X1 us30_U296 (.ZN( us30_n540 ) , .A( us30_n763 ) , .B2( us30_n779 ) , .B1( us30_n817 ) );
  AOI21_X1 us30_U297 (.B1( us30_n699 ) , .ZN( us30_n700 ) , .A( us30_n732 ) , .B2( us30_n763 ) );
  AOI21_X1 us30_U298 (.ZN( us30_n591 ) , .B2( us30_n763 ) , .A( us30_n785 ) , .B1( us30_n812 ) );
  AOI21_X1 us30_U299 (.ZN( us30_n498 ) , .A( us30_n724 ) , .B2( us30_n762 ) , .B1( us30_n814 ) );
  NAND2_X1 us30_U3 (.A2( us30_n448 ) , .A1( us30_n464 ) , .ZN( us30_n815 ) );
  AOI221_X1 us30_U30 (.A( us30_n713 ) , .B2( us30_n714 ) , .ZN( us30_n720 ) , .C1( us30_n832 ) , .B1( us30_n839 ) , .C2( us30_n863 ) );
  NOR2_X1 us30_U300 (.ZN( us30_n547 ) , .A1( us30_n699 ) , .A2( us30_n744 ) );
  INV_X1 us30_U301 (.A( us30_n791 ) , .ZN( us30_n873 ) );
  AOI21_X1 us30_U302 (.ZN( us30_n649 ) , .B1( us30_n729 ) , .B2( us30_n763 ) , .A( us30_n813 ) );
  NOR2_X1 us30_U303 (.ZN( us30_n685 ) , .A1( us30_n729 ) , .A2( us30_n816 ) );
  AOI21_X1 us30_U304 (.B1( us30_n686 ) , .ZN( us30_n687 ) , .A( us30_n728 ) , .B2( us30_n761 ) );
  AOI21_X1 us30_U305 (.ZN( us30_n569 ) , .B1( us30_n750 ) , .B2( us30_n762 ) , .A( us30_n780 ) );
  AOI21_X1 us30_U306 (.ZN( us30_n571 ) , .B2( us30_n697 ) , .B1( us30_n806 ) , .A( us30_n812 ) );
  NOR2_X1 us30_U307 (.ZN( us30_n568 ) , .A1( us30_n729 ) , .A2( us30_n762 ) );
  NOR2_X1 us30_U308 (.ZN( us30_n566 ) , .A2( us30_n697 ) , .A1( us30_n763 ) );
  AOI21_X1 us30_U309 (.ZN( us30_n640 ) , .B2( us30_n747 ) , .A( us30_n792 ) , .B1( us30_n803 ) );
  OR2_X1 us30_U31 (.A2( us30_n711 ) , .A1( us30_n712 ) , .ZN( us30_n713 ) );
  INV_X1 us30_U310 (.A( us30_n699 ) , .ZN( us30_n853 ) );
  AOI21_X1 us30_U311 (.ZN( us30_n514 ) , .A( us30_n779 ) , .B2( us30_n792 ) , .B1( us30_n812 ) );
  AOI21_X1 us30_U312 (.ZN( us30_n639 ) , .B2( us30_n749 ) , .A( us30_n788 ) , .B1( us30_n812 ) );
  NAND2_X1 us30_U313 (.ZN( us30_n753 ) , .A1( us30_n763 ) , .A2( us30_n805 ) );
  NOR2_X1 us30_U314 (.ZN( us30_n665 ) , .A1( us30_n780 ) , .A2( us30_n813 ) );
  AOI21_X1 us30_U315 (.ZN( us30_n564 ) , .B1( us30_n724 ) , .A( us30_n779 ) , .B2( us30_n791 ) );
  AOI21_X1 us30_U316 (.ZN( us30_n497 ) , .A( us30_n779 ) , .B2( us30_n791 ) , .B1( us30_n804 ) );
  AOI21_X1 us30_U317 (.ZN( us30_n689 ) , .B2( us30_n749 ) , .B1( us30_n763 ) , .A( us30_n806 ) );
  AOI21_X1 us30_U318 (.ZN( us30_n450 ) , .B2( us30_n792 ) , .A( us30_n803 ) , .B1( us30_n815 ) );
  NOR2_X1 us30_U319 (.ZN( us30_n567 ) , .A1( us30_n747 ) , .A2( us30_n805 ) );
  NOR2_X1 us30_U32 (.ZN( us30_n680 ) , .A2( us30_n834 ) , .A1( us30_n839 ) );
  NOR2_X1 us30_U320 (.ZN( us30_n529 ) , .A1( us30_n708 ) , .A2( us30_n779 ) );
  NOR2_X1 us30_U321 (.ZN( us30_n578 ) , .A1( us30_n708 ) , .A2( us30_n813 ) );
  AOI21_X1 us30_U322 (.ZN( us30_n478 ) , .B2( us30_n697 ) , .A( us30_n749 ) , .B1( us30_n779 ) );
  AOI21_X1 us30_U323 (.A( us30_n790 ) , .B2( us30_n791 ) , .B1( us30_n792 ) , .ZN( us30_n793 ) );
  NOR2_X1 us30_U324 (.ZN( us30_n684 ) , .A1( us30_n791 ) , .A2( us30_n813 ) );
  AOI21_X1 us30_U325 (.A( us30_n733 ) , .ZN( us30_n734 ) , .B2( us30_n780 ) , .B1( us30_n792 ) );
  NOR2_X1 us30_U326 (.A2( us30_n813 ) , .A1( us30_n815 ) , .ZN( us30_n821 ) );
  AOI21_X1 us30_U327 (.ZN( us30_n641 ) , .B1( us30_n680 ) , .A( us30_n791 ) , .B2( us30_n817 ) );
  NOR2_X1 us30_U328 (.ZN( us30_n711 ) , .A1( us30_n762 ) , .A2( us30_n763 ) );
  NOR2_X1 us30_U329 (.ZN( us30_n583 ) , .A1( us30_n792 ) , .A2( us30_n817 ) );
  AOI222_X1 us30_U33 (.ZN( us30_n469 ) , .B1( us30_n832 ) , .A1( us30_n839 ) , .C1( us30_n842 ) , .C2( us30_n851 ) , .A2( us30_n855 ) , .B2( us30_n865 ) );
  NOR2_X1 us30_U330 (.ZN( us30_n534 ) , .A1( us30_n724 ) , .A2( us30_n788 ) );
  NOR2_X1 us30_U331 (.ZN( us30_n632 ) , .A2( us30_n697 ) , .A1( us30_n724 ) );
  NOR2_X1 us30_U332 (.ZN( us30_n682 ) , .A2( us30_n708 ) , .A1( us30_n817 ) );
  NOR2_X1 us30_U333 (.ZN( us30_n580 ) , .A2( us30_n697 ) , .A1( us30_n791 ) );
  INV_X1 us30_U334 (.A( us30_n815 ) , .ZN( us30_n855 ) );
  AOI21_X1 us30_U335 (.ZN( us30_n442 ) , .A( us30_n699 ) , .B1( us30_n733 ) , .B2( us30_n750 ) );
  INV_X1 us30_U336 (.A( us30_n780 ) , .ZN( us30_n850 ) );
  INV_X1 us30_U337 (.A( us30_n785 ) , .ZN( us30_n846 ) );
  NAND2_X1 us30_U338 (.ZN( us30_n714 ) , .A1( us30_n728 ) , .A2( us30_n780 ) );
  NAND2_X1 us30_U339 (.A2( us30_n762 ) , .A1( us30_n806 ) , .ZN( us30_n810 ) );
  NOR4_X1 us30_U34 (.A1( us30_n466 ) , .ZN( us30_n467 ) , .A4( us30_n542 ) , .A2( us30_n554 ) , .A3( us30_n614 ) );
  AOI21_X1 us30_U340 (.ZN( us30_n443 ) , .B1( us30_n789 ) , .B2( us30_n791 ) , .A( us30_n814 ) );
  NAND2_X1 us30_U341 (.ZN( us30_n671 ) , .A1( us30_n806 ) , .A2( us30_n816 ) );
  NOR2_X1 us30_U342 (.ZN( us30_n484 ) , .A1( us30_n788 ) , .A2( us30_n805 ) );
  NOR2_X1 us30_U343 (.ZN( us30_n470 ) , .A2( us30_n779 ) , .A1( us30_n815 ) );
  NOR2_X1 us30_U344 (.ZN( us30_n712 ) , .A2( us30_n724 ) , .A1( us30_n790 ) );
  OAI21_X1 us30_U345 (.A( us30_n787 ) , .B2( us30_n788 ) , .B1( us30_n789 ) , .ZN( us30_n795 ) );
  OAI21_X1 us30_U346 (.ZN( us30_n787 ) , .A( us30_n839 ) , .B1( us30_n863 ) , .B2( us30_n873 ) );
  NOR2_X1 us30_U347 (.ZN( us30_n526 ) , .A1( us30_n724 ) , .A2( us30_n750 ) );
  NAND2_X1 us30_U348 (.A1( us30_n699 ) , .A2( us30_n729 ) , .ZN( us30_n782 ) );
  NOR2_X1 us30_U349 (.ZN( us30_n518 ) , .A1( us30_n708 ) , .A2( us30_n788 ) );
  AOI221_X1 us30_U35 (.ZN( us30_n468 ) , .C2( us30_n714 ) , .B2( us30_n831 ) , .C1( us30_n845 ) , .B1( us30_n860 ) , .A( us30_n864 ) );
  OAI21_X1 us30_U350 (.A( us30_n698 ) , .ZN( us30_n702 ) , .B2( us30_n750 ) , .B1( us30_n804 ) );
  OAI21_X1 us30_U351 (.ZN( us30_n698 ) , .B2( us30_n833 ) , .B1( us30_n838 ) , .A( us30_n860 ) );
  OAI21_X1 us30_U352 (.A( us30_n731 ) , .B1( us30_n732 ) , .ZN( us30_n736 ) , .B2( us30_n805 ) );
  OAI21_X1 us30_U353 (.ZN( us30_n731 ) , .A( us30_n833 ) , .B2( us30_n852 ) , .B1( us30_n873 ) );
  INV_X1 us30_U354 (.A( us30_n817 ) , .ZN( us30_n844 ) );
  INV_X1 us30_U355 (.A( us30_n724 ) , .ZN( us30_n856 ) );
  AND2_X1 us30_U356 (.ZN( us30_n732 ) , .A1( us30_n779 ) , .A2( us30_n785 ) );
  NAND2_X1 us30_U357 (.A1( us30_n447 ) , .A2( us30_n449 ) , .ZN( us30_n805 ) );
  NAND2_X1 us30_U359 (.A1( us30_n452 ) , .A2( us30_n465 ) , .ZN( us30_n669 ) );
  NOR4_X1 us30_U36 (.A4( us30_n514 ) , .A3( us30_n515 ) , .A2( us30_n516 ) , .A1( us30_n517 ) , .ZN( us30_n524 ) );
  NAND2_X1 us30_U360 (.A2( us30_n448 ) , .A1( us30_n460 ) , .ZN( us30_n728 ) );
  NAND2_X1 us30_U369 (.A2( us30_n464 ) , .A1( us30_n465 ) , .ZN( us30_n812 ) );
  AOI222_X1 us30_U37 (.ZN( us30_n525 ) , .A1( us30_n834 ) , .B2( us30_n837 ) , .C1( us30_n844 ) , .C2( us30_n850 ) , .A2( us30_n852 ) , .B1( us30_n866 ) );
  NAND2_X1 us30_U370 (.A1( us30_n441 ) , .A2( us30_n460 ) , .ZN( us30_n699 ) );
  NAND2_X1 us30_U371 (.A2( us30_n449 ) , .A1( us30_n452 ) , .ZN( us30_n763 ) );
  NAND2_X1 us30_U372 (.A2( us30_n448 ) , .A1( us30_n452 ) , .ZN( us30_n729 ) );
  NAND2_X1 us30_U379 (.A2( us30_n441 ) , .A1( us30_n447 ) , .ZN( us30_n784 ) );
  NOR4_X1 us30_U38 (.A3( us30_n521 ) , .A1( us30_n522 ) , .ZN( us30_n523 ) , .A2( us30_n673 ) , .A4( us30_n769 ) );
  NAND2_X2 us30_U381 (.A1( us30_n449 ) , .A2( us30_n464 ) , .ZN( us30_n724 ) );
  NAND2_X2 us30_U382 (.A1( us30_n449 ) , .A2( us30_n460 ) , .ZN( us30_n792 ) );
  NAND2_X2 us30_U383 (.A2( us30_n460 ) , .A1( us30_n465 ) , .ZN( us30_n780 ) );
  NAND2_X1 us30_U385 (.A1( us30_n447 ) , .A2( us30_n448 ) , .ZN( us30_n786 ) );
  NOR2_X1 us30_U386 (.A2( sa30_6 ) , .A1( sa30_7 ) , .ZN( us30_n464 ) );
  AOI221_X1 us30_U39 (.A( us30_n781 ) , .ZN( us30_n798 ) , .C2( us30_n837 ) , .B2( us30_n838 ) , .B1( us30_n865 ) , .C1( us30_n866 ) );
  NAND2_X1 us30_U4 (.A1( us30_n441 ) , .A2( us30_n464 ) , .ZN( us30_n708 ) );
  NOR4_X1 us30_U40 (.A4( us30_n793 ) , .A3( us30_n794 ) , .A2( us30_n795 ) , .A1( us30_n796 ) , .ZN( us30_n797 ) );
  OAI221_X1 us30_U407 (.A( us30_n783 ) , .C2( us30_n784 ) , .B2( us30_n785 ) , .B1( us30_n786 ) , .ZN( us30_n796 ) , .C1( us30_n813 ) );
  NAND2_X1 us30_U408 (.A1( us30_n729 ) , .A2( us30_n784 ) , .ZN( us30_n811 ) );
  OAI22_X1 us30_U409 (.ZN( us30_n588 ) , .A2( us30_n747 ) , .B2( us30_n762 ) , .A1( us30_n763 ) , .B1( us30_n784 ) );
  NOR4_X1 us30_U41 (.A4( us30_n776 ) , .A3( us30_n777 ) , .A1( us30_n778 ) , .ZN( us30_n799 ) , .A2( us30_n801 ) );
  AOI21_X1 us30_U410 (.ZN( us30_n592 ) , .B1( us30_n728 ) , .B2( us30_n784 ) , .A( us30_n790 ) );
  AOI21_X1 us30_U411 (.ZN( us30_n623 ) , .B1( us30_n699 ) , .A( us30_n779 ) , .B2( us30_n784 ) );
  AOI21_X1 us30_U412 (.ZN( us30_n648 ) , .A( us30_n762 ) , .B2( us30_n784 ) , .B1( us30_n792 ) );
  OAI22_X1 us30_U413 (.ZN( us30_n681 ) , .A1( us30_n699 ) , .A2( us30_n730 ) , .B2( us30_n784 ) , .B1( us30_n817 ) );
  OAI21_X1 us30_U414 (.A( us30_n613 ) , .ZN( us30_n616 ) , .B1( us30_n625 ) , .B2( us30_n784 ) );
  NOR2_X1 us30_U415 (.ZN( us30_n610 ) , .A1( us30_n784 ) , .A2( us30_n816 ) );
  OAI222_X1 us30_U416 (.A2( us30_n669 ) , .ZN( us30_n674 ) , .B1( us30_n747 ) , .B2( us30_n784 ) , .C2( us30_n788 ) , .C1( us30_n815 ) , .A1( us30_n817 ) );
  NOR2_X1 us30_U417 (.ZN( us30_n651 ) , .A1( us30_n784 ) , .A2( us30_n788 ) );
  NOR2_X1 us30_U418 (.ZN( us30_n600 ) , .A2( us30_n697 ) , .A1( us30_n784 ) );
  NOR2_X1 us30_U419 (.ZN( us30_n553 ) , .A2( us30_n744 ) , .A1( us30_n784 ) );
  NOR4_X1 us30_U42 (.A3( us30_n755 ) , .A2( us30_n756 ) , .A1( us30_n757 ) , .ZN( us30_n758 ) , .A4( us30_n869 ) );
  INV_X1 us30_U420 (.A( us30_n784 ) , .ZN( us30_n861 ) );
  AOI21_X1 us30_U421 (.ZN( us30_n500 ) , .A( us30_n697 ) , .B1( us30_n708 ) , .B2( us30_n786 ) );
  OAI221_X1 us30_U422 (.A( us30_n696 ) , .ZN( us30_n703 ) , .C2( us30_n784 ) , .C1( us30_n785 ) , .B1( us30_n786 ) , .B2( us30_n806 ) );
  OAI22_X1 us30_U423 (.ZN( us30_n590 ) , .B1( us30_n730 ) , .B2( us30_n749 ) , .A2( us30_n786 ) , .A1( us30_n803 ) );
  NOR2_X1 us30_U424 (.ZN( us30_n612 ) , .A1( us30_n779 ) , .A2( us30_n786 ) );
  NAND2_X1 us30_U425 (.A2( us30_n749 ) , .A1( us30_n786 ) , .ZN( us30_n809 ) );
  OAI222_X1 us30_U426 (.ZN( us30_n617 ) , .B1( us30_n697 ) , .C1( us30_n724 ) , .C2( us30_n747 ) , .B2( us30_n786 ) , .A2( us30_n792 ) , .A1( us30_n816 ) );
  NOR2_X1 us30_U427 (.ZN( us30_n717 ) , .A2( us30_n744 ) , .A1( us30_n786 ) );
  NOR2_X1 us30_U428 (.ZN( us30_n653 ) , .A1( us30_n762 ) , .A2( us30_n786 ) );
  NOR2_X1 us30_U429 (.ZN( us30_n554 ) , .A1( us30_n786 ) , .A2( us30_n813 ) );
  AOI211_X1 us30_U43 (.B( us30_n745 ) , .A( us30_n746 ) , .ZN( us30_n759 ) , .C1( us30_n832 ) , .C2( us30_n853 ) );
  NOR2_X1 us30_U430 (.ZN( us30_n701 ) , .A2( us30_n786 ) , .A1( us30_n817 ) );
  NOR2_X1 us30_U431 (.A1( us30_n730 ) , .ZN( us30_n765 ) , .A2( us30_n786 ) );
  AND2_X1 us30_U432 (.ZN( us30_n438 ) , .A2( us30_n831 ) , .A1( us30_n854 ) );
  AND2_X1 us30_U433 (.ZN( us30_n439 ) , .A2( us30_n843 ) , .A1( us30_n861 ) );
  NOR3_X1 us30_U434 (.A1( us30_n438 ) , .A2( us30_n439 ) , .A3( us30_n576 ) , .ZN( us30_n587 ) );
  NAND4_X1 us30_U435 (.ZN( sa31_sr_2 ) , .A4( us30_n643 ) , .A3( us30_n644 ) , .A2( us30_n645 ) , .A1( us30_n646 ) );
  INV_X1 us30_U436 (.A( us30_n812 ) , .ZN( us30_n854 ) );
  NAND3_X1 us30_U437 (.ZN( sa31_sr_6 ) , .A3( us30_n797 ) , .A2( us30_n798 ) , .A1( us30_n799 ) );
  NAND3_X1 us30_U438 (.ZN( sa31_sr_5 ) , .A3( us30_n758 ) , .A2( us30_n759 ) , .A1( us30_n760 ) );
  NAND3_X1 us30_U439 (.ZN( sa31_sr_4 ) , .A3( us30_n738 ) , .A2( us30_n739 ) , .A1( us30_n740 ) );
  NOR3_X1 us30_U44 (.A3( us30_n741 ) , .A2( us30_n742 ) , .A1( us30_n743 ) , .ZN( us30_n760 ) );
  NAND3_X1 us30_U440 (.A3( us30_n675 ) , .A2( us30_n676 ) , .A1( us30_n677 ) , .ZN( us30_n807 ) );
  NAND3_X1 us30_U441 (.ZN( us30_n638 ) , .A3( us30_n708 ) , .A2( us30_n724 ) , .A1( us30_n792 ) );
  NAND3_X1 us30_U442 (.A3( us30_n618 ) , .A2( us30_n619 ) , .A1( us30_n620 ) , .ZN( us30_n725 ) );
  NAND3_X1 us30_U443 (.A3( us30_n585 ) , .A2( us30_n586 ) , .A1( us30_n587 ) , .ZN( us30_n621 ) );
  NAND3_X1 us30_U444 (.ZN( us30_n565 ) , .A3( us30_n680 ) , .A2( us30_n750 ) , .A1( us30_n785 ) );
  NAND3_X1 us30_U445 (.A3( us30_n523 ) , .A2( us30_n524 ) , .A1( us30_n525 ) , .ZN( us30_n742 ) );
  NAND3_X1 us30_U446 (.A3( us30_n512 ) , .A1( us30_n513 ) , .ZN( us30_n608 ) , .A2( us30_n871 ) );
  NAND3_X1 us30_U447 (.A3( us30_n467 ) , .A2( us30_n468 ) , .A1( us30_n469 ) , .ZN( us30_n777 ) );
  INV_X1 us30_U448 (.A( us30_n803 ) , .ZN( us30_n843 ) );
  AOI21_X1 us30_U449 (.ZN( us30_n576 ) , .B2( us30_n724 ) , .B1( us30_n748 ) , .A( us30_n785 ) );
  NAND4_X1 us30_U45 (.ZN( sa31_sr_3 ) , .A4( us30_n704 ) , .A3( us30_n705 ) , .A2( us30_n706 ) , .A1( us30_n707 ) );
  NOR4_X1 us30_U46 (.A4( us30_n700 ) , .A3( us30_n701 ) , .A2( us30_n702 ) , .A1( us30_n703 ) , .ZN( us30_n704 ) );
  AOI211_X1 us30_U47 (.B( us30_n694 ) , .A( us30_n695 ) , .ZN( us30_n705 ) , .C2( us30_n831 ) , .C1( us30_n851 ) );
  NOR2_X1 us30_U48 (.ZN( us30_n707 ) , .A2( us30_n776 ) , .A1( us30_n800 ) );
  AOI222_X1 us30_U49 (.B2( us30_n638 ) , .ZN( us30_n644 ) , .B1( us30_n841 ) , .A1( us30_n842 ) , .C2( us30_n846 ) , .C1( us30_n863 ) , .A2( us30_n865 ) );
  NAND2_X1 us30_U5 (.A2( us30_n441 ) , .A1( us30_n452 ) , .ZN( us30_n791 ) );
  NOR4_X1 us30_U50 (.A4( us30_n639 ) , .A3( us30_n640 ) , .A2( us30_n641 ) , .A1( us30_n642 ) , .ZN( us30_n643 ) );
  NOR3_X1 us30_U51 (.A2( us30_n607 ) , .A1( us30_n608 ) , .ZN( us30_n646 ) , .A3( us30_n722 ) );
  NOR2_X1 us30_U52 (.ZN( us30_n804 ) , .A1( us30_n854 ) , .A2( us30_n861 ) );
  NAND4_X1 us30_U53 (.ZN( sa31_sr_7 ) , .A4( us30_n822 ) , .A3( us30_n823 ) , .A2( us30_n824 ) , .A1( us30_n825 ) );
  NOR4_X1 us30_U54 (.A4( us30_n818 ) , .A3( us30_n819 ) , .A2( us30_n820 ) , .A1( us30_n821 ) , .ZN( us30_n822 ) );
  AOI222_X1 us30_U55 (.C2( us30_n809 ) , .B2( us30_n810 ) , .A2( us30_n811 ) , .ZN( us30_n823 ) , .C1( us30_n832 ) , .A1( us30_n839 ) , .B1( us30_n853 ) );
  AOI211_X1 us30_U56 (.B( us30_n807 ) , .A( us30_n808 ) , .ZN( us30_n824 ) , .C1( us30_n842 ) , .C2( us30_n850 ) );
  NAND4_X1 us30_U57 (.ZN( sa31_sr_0 ) , .A4( us30_n501 ) , .A3( us30_n502 ) , .A2( us30_n503 ) , .A1( us30_n504 ) );
  AOI221_X1 us30_U58 (.A( us30_n497 ) , .ZN( us30_n502 ) , .B2( us30_n843 ) , .C1( us30_n846 ) , .C2( us30_n860 ) , .B1( us30_n862 ) );
  NOR4_X1 us30_U59 (.A4( us30_n498 ) , .A3( us30_n499 ) , .A2( us30_n500 ) , .ZN( us30_n501 ) , .A1( us30_n527 ) );
  AOI211_X1 us30_U60 (.A( us30_n496 ) , .ZN( us30_n503 ) , .B( us30_n802 ) , .C2( us30_n839 ) , .C1( us30_n851 ) );
  NAND4_X1 us30_U61 (.ZN( sa31_sr_1 ) , .A4( us30_n595 ) , .A3( us30_n596 ) , .A2( us30_n597 ) , .A1( us30_n598 ) );
  NOR4_X1 us30_U62 (.A4( us30_n591 ) , .A3( us30_n592 ) , .A2( us30_n593 ) , .A1( us30_n594 ) , .ZN( us30_n595 ) );
  AOI211_X1 us30_U63 (.B( us30_n589 ) , .A( us30_n590 ) , .ZN( us30_n596 ) , .C2( us30_n811 ) , .C1( us30_n833 ) );
  AOI211_X1 us30_U64 (.A( us30_n588 ) , .ZN( us30_n597 ) , .B( us30_n621 ) , .C1( us30_n845 ) , .C2( us30_n855 ) );
  NOR2_X1 us30_U65 (.ZN( us30_n748 ) , .A1( us30_n861 ) , .A2( us30_n862 ) );
  NOR2_X1 us30_U66 (.ZN( us30_n625 ) , .A2( us30_n836 ) , .A1( us30_n839 ) );
  NAND4_X1 us30_U67 (.A4( us30_n603 ) , .A3( us30_n604 ) , .A2( us30_n605 ) , .A1( us30_n606 ) , .ZN( us30_n722 ) );
  NOR3_X1 us30_U68 (.A1( us30_n599 ) , .ZN( us30_n604 ) , .A3( us30_n663 ) , .A2( us30_n770 ) );
  NOR4_X1 us30_U69 (.A3( us30_n600 ) , .A2( us30_n601 ) , .A1( us30_n602 ) , .ZN( us30_n603 ) , .A4( us30_n655 ) );
  NOR3_X1 us30_U7 (.ZN( us30_n598 ) , .A1( us30_n608 ) , .A3( us30_n723 ) , .A2( us30_n742 ) );
  AOI222_X1 us30_U70 (.ZN( us30_n606 ) , .A1( us30_n830 ) , .C2( us30_n837 ) , .B1( us30_n842 ) , .A2( us30_n856 ) , .B2( us30_n861 ) , .C1( us30_n868 ) );
  NAND4_X1 us30_U71 (.A4( us30_n657 ) , .A3( us30_n658 ) , .A2( us30_n659 ) , .A1( us30_n660 ) , .ZN( us30_n800 ) );
  NOR3_X1 us30_U72 (.A3( us30_n648 ) , .A2( us30_n649 ) , .A1( us30_n650 ) , .ZN( us30_n659 ) );
  NOR3_X1 us30_U73 (.A3( us30_n651 ) , .A2( us30_n652 ) , .A1( us30_n653 ) , .ZN( us30_n658 ) );
  NOR3_X1 us30_U74 (.A3( us30_n654 ) , .A2( us30_n655 ) , .A1( us30_n656 ) , .ZN( us30_n657 ) );
  NAND4_X1 us30_U75 (.A4( us30_n560 ) , .A3( us30_n561 ) , .A2( us30_n562 ) , .A1( us30_n563 ) , .ZN( us30_n607 ) );
  NOR4_X1 us30_U76 (.ZN( us30_n561 ) , .A1( us30_n653 ) , .A3( us30_n661 ) , .A4( us30_n685 ) , .A2( us30_n768 ) );
  NOR4_X1 us30_U77 (.A4( us30_n552 ) , .A3( us30_n553 ) , .A2( us30_n554 ) , .A1( us30_n555 ) , .ZN( us30_n562 ) );
  NOR4_X1 us30_U78 (.A4( us30_n556 ) , .A3( us30_n557 ) , .A2( us30_n558 ) , .A1( us30_n559 ) , .ZN( us30_n560 ) );
  NAND4_X1 us30_U79 (.A4( us30_n772 ) , .A3( us30_n773 ) , .A2( us30_n774 ) , .A1( us30_n775 ) , .ZN( us30_n801 ) );
  NOR3_X1 us30_U8 (.A3( us30_n800 ) , .A2( us30_n801 ) , .A1( us30_n802 ) , .ZN( us30_n825 ) );
  NOR3_X1 us30_U80 (.A3( us30_n765 ) , .A2( us30_n766 ) , .A1( us30_n767 ) , .ZN( us30_n773 ) );
  NOR4_X1 us30_U81 (.A4( us30_n768 ) , .A3( us30_n769 ) , .A2( us30_n770 ) , .A1( us30_n771 ) , .ZN( us30_n772 ) );
  AOI222_X1 us30_U82 (.ZN( us30_n775 ) , .A1( us30_n830 ) , .C1( us30_n834 ) , .B2( us30_n841 ) , .A2( us30_n850 ) , .B1( us30_n861 ) , .C2( us30_n873 ) );
  NOR4_X1 us30_U83 (.A4( us30_n665 ) , .A3( us30_n666 ) , .A2( us30_n667 ) , .A1( us30_n668 ) , .ZN( us30_n676 ) );
  NOR4_X1 us30_U84 (.A4( us30_n661 ) , .A3( us30_n662 ) , .A2( us30_n663 ) , .A1( us30_n664 ) , .ZN( us30_n677 ) );
  NOR4_X1 us30_U85 (.A3( us30_n673 ) , .A1( us30_n674 ) , .ZN( us30_n675 ) , .A4( us30_n715 ) , .A2( us30_n859 ) );
  NOR2_X1 us30_U86 (.ZN( us30_n761 ) , .A1( us30_n833 ) , .A2( us30_n834 ) );
  NOR4_X1 us30_U87 (.A4( us30_n577 ) , .A3( us30_n578 ) , .A2( us30_n579 ) , .ZN( us30_n586 ) , .A1( us30_n683 ) );
  NOR4_X1 us30_U88 (.A1( us30_n584 ) , .ZN( us30_n585 ) , .A3( us30_n652 ) , .A2( us30_n662 ) , .A4( us30_n767 ) );
  AOI222_X1 us30_U89 (.ZN( us30_n513 ) , .C1( us30_n832 ) , .B2( us30_n837 ) , .A2( us30_n843 ) , .C2( us30_n862 ) , .B1( us30_n863 ) , .A1( us30_n866 ) );
  NOR3_X1 us30_U9 (.A3( us30_n621 ) , .A2( us30_n622 ) , .ZN( us30_n636 ) , .A1( us30_n725 ) );
  NOR4_X1 us30_U90 (.A4( us30_n509 ) , .A2( us30_n510 ) , .A1( us30_n511 ) , .ZN( us30_n512 ) , .A3( us30_n670 ) );
  INV_X1 us30_U91 (.A( us30_n505 ) , .ZN( us30_n871 ) );
  NAND4_X1 us30_U92 (.A4( us30_n456 ) , .A3( us30_n457 ) , .A2( us30_n458 ) , .A1( us30_n459 ) , .ZN( us30_n679 ) );
  NOR3_X1 us30_U93 (.ZN( us30_n457 ) , .A3( us30_n530 ) , .A1( us30_n555 ) , .A2( us30_n570 ) );
  AOI221_X1 us30_U94 (.A( us30_n450 ) , .ZN( us30_n459 ) , .C2( us30_n753 ) , .B1( us30_n832 ) , .C1( us30_n842 ) , .B2( us30_n861 ) );
  NOR4_X1 us30_U95 (.ZN( us30_n458 ) , .A2( us30_n509 ) , .A1( us30_n599 ) , .A4( us30_n628 ) , .A3( us30_n711 ) );
  NAND4_X1 us30_U96 (.A4( us30_n535 ) , .A3( us30_n536 ) , .A2( us30_n537 ) , .A1( us30_n538 ) , .ZN( us30_n622 ) );
  NOR4_X1 us30_U97 (.A4( us30_n526 ) , .A2( us30_n527 ) , .A1( us30_n528 ) , .ZN( us30_n538 ) , .A3( us30_n701 ) );
  NOR4_X1 us30_U98 (.A1( us30_n531 ) , .ZN( us30_n536 ) , .A2( us30_n654 ) , .A4( us30_n668 ) , .A3( us30_n765 ) );
  NOR4_X1 us30_U99 (.A4( us30_n529 ) , .A3( us30_n530 ) , .ZN( us30_n537 ) , .A2( us30_n684 ) , .A1( us30_n794 ) );
endmodule

