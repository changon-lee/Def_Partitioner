module des_des_die_11 ( u0_K14_4, u0_K14_42, u0_K14_46, u0_K15_18, u0_L12_12, u0_L12_15, u0_L12_17, u0_L12_21, u0_L12_22, 
       u0_L12_23, u0_L12_27, u0_L12_31, u0_L12_32, u0_L12_5, u0_L12_7, u0_L12_9, u0_L13_13, u0_L13_16, 
       u0_L13_17, u0_L13_18, u0_L13_2, u0_L13_23, u0_L13_24, u0_L13_28, u0_L13_30, u0_L13_31, u0_L13_6, 
       u0_L13_9, u0_L4_15, u0_L4_21, u0_L4_27, u0_L4_5, u0_R12_1, u0_R12_2, u0_R12_24, u0_R12_25, 
       u0_R12_26, u0_R12_27, u0_R12_28, u0_R12_29, u0_R12_3, u0_R12_30, u0_R12_31, u0_R12_32, u0_R12_4, 
       u0_R12_5, u0_R13_1, u0_R13_10, u0_R13_11, u0_R13_12, u0_R13_13, u0_R13_2, u0_R13_3, u0_R13_32, 
       u0_R13_4, u0_R13_5, u0_R13_6, u0_R13_7, u0_R13_8, u0_R13_9, u0_R4_1, u0_R4_28, u0_R4_29, 
       u0_R4_30, u0_R4_31, u0_R4_32, u0_uk_K_r12_10, u0_uk_K_r12_15, u0_uk_K_r12_16, u0_uk_K_r12_21, u0_uk_K_r12_47, u0_uk_K_r13_13, 
       u0_uk_K_r13_17, u0_uk_K_r13_19, u0_uk_K_r13_25, u0_uk_K_r13_32, u0_uk_K_r13_4, u0_uk_K_r13_55, u0_uk_K_r4_23, u0_uk_n1, u0_uk_n10, 
       u0_uk_n100, u0_uk_n109, u0_uk_n11, u0_uk_n110, u0_uk_n117, u0_uk_n118, u0_uk_n128, u0_uk_n14, u0_uk_n141, 
       u0_uk_n146, u0_uk_n15, u0_uk_n155, u0_uk_n16, u0_uk_n17, u0_uk_n187, u0_uk_n19, u0_uk_n20, u0_uk_n203, 
       u0_uk_n208, u0_uk_n213, u0_uk_n214, u0_uk_n217, u0_uk_n220, u0_uk_n222, u0_uk_n230, u0_uk_n24, u0_uk_n240, 
       u0_uk_n242, u0_uk_n25, u0_uk_n250, u0_uk_n251, u0_uk_n252, u0_uk_n26, u0_uk_n27, u0_uk_n29, u0_uk_n30, 
       u0_uk_n35, u0_uk_n36, u0_uk_n37, u0_uk_n38, u0_uk_n411, u0_uk_n412, u0_uk_n417, u0_uk_n418, u0_uk_n425, 
       u0_uk_n429, u0_uk_n43, u0_uk_n430, u0_uk_n434, u0_uk_n439, u0_uk_n44, u0_uk_n445, u0_uk_n450, u0_uk_n46, 
       u0_uk_n52, u0_uk_n56, u0_uk_n57, u0_uk_n58, u0_uk_n59, u0_uk_n6, u0_uk_n60, u0_uk_n62, u0_uk_n63, 
       u0_uk_n64, u0_uk_n65, u0_uk_n67, u0_uk_n68, u0_uk_n73, u0_uk_n75, u0_uk_n77, u0_uk_n78, u0_uk_n8, 
       u0_uk_n80, u0_uk_n81, u0_uk_n82, u0_uk_n85, u0_uk_n90, u0_uk_n92, u0_uk_n94, u1_L10_14, u1_L10_25, 
       u1_L10_3, u1_L10_8, u1_L12_1, u1_L12_10, u1_L12_20, u1_L12_26, u1_L1_12, u1_L1_15, u1_L1_21, 
       u1_L1_22, u1_L1_27, u1_L1_32, u1_L1_5, u1_L1_7, u1_L2_14, u1_L2_25, u1_L2_3, u1_L2_8, 
       u1_L3_1, u1_L3_10, u1_L3_20, u1_L3_26, u1_L6_1, u1_L6_10, u1_L6_20, u1_L6_26, u1_L8_1, 
       u1_L8_10, u1_L8_20, u1_L8_26, u1_R10_16, u1_R10_17, u1_R10_18, u1_R10_19, u1_R10_20, u1_R10_21, 
       u1_R12_12, u1_R12_13, u1_R12_14, u1_R12_15, u1_R12_16, u1_R12_17, u1_R1_1, u1_R1_24, u1_R1_25, 
       u1_R1_26, u1_R1_27, u1_R1_28, u1_R1_29, u1_R1_30, u1_R1_31, u1_R1_32, u1_R2_16, u1_R2_17, 
       u1_R2_18, u1_R2_19, u1_R2_20, u1_R2_21, u1_R3_12, u1_R3_13, u1_R3_14, u1_R3_15, u1_R3_16, 
       u1_R3_17, u1_R6_12, u1_R6_13, u1_R6_14, u1_R6_15, u1_R6_16, u1_R6_17, u1_R8_12, u1_R8_13, 
       u1_R8_14, u1_R8_15, u1_R8_16, u1_R8_17, u1_uk_K_r10_23, u1_uk_K_r10_42, u1_uk_K_r12_25, u1_uk_K_r12_33, u1_uk_K_r12_41, 
       u1_uk_K_r1_15, u1_uk_K_r1_16, u1_uk_K_r1_21, u1_uk_K_r1_22, u1_uk_K_r2_16, u1_uk_K_r2_21, u1_uk_K_r2_28, u1_uk_K_r2_31, u1_uk_K_r2_36, 
       u1_uk_K_r2_49, u1_uk_K_r2_7, u1_uk_K_r3_24, u1_uk_K_r3_33, u1_uk_K_r3_47, u1_uk_K_r8_13, u1_uk_K_r8_19, u1_uk_K_r8_27, u1_uk_K_r8_40, 
       u1_uk_K_r8_5, u1_uk_n10, u1_uk_n100, u1_uk_n102, u1_uk_n109, u1_uk_n11, u1_uk_n117, u1_uk_n118, u1_uk_n128, 
       u1_uk_n1307, u1_uk_n1313, u1_uk_n1314, u1_uk_n1318, u1_uk_n1322, u1_uk_n1327, u1_uk_n1328, u1_uk_n1330, u1_uk_n1334, 
       u1_uk_n1335, u1_uk_n1338, u1_uk_n1342, u1_uk_n1350, u1_uk_n1375, u1_uk_n1376, u1_uk_n1381, u1_uk_n1398, u1_uk_n1402, 
       u1_uk_n1409, u1_uk_n1415, u1_uk_n142, u1_uk_n1424, u1_uk_n1427, u1_uk_n1429, u1_uk_n1435, u1_uk_n145, u1_uk_n146, 
       u1_uk_n147, u1_uk_n148, u1_uk_n1530, u1_uk_n1538, u1_uk_n1543, u1_uk_n1545, u1_uk_n1548, u1_uk_n155, u1_uk_n1551, 
       u1_uk_n1552, u1_uk_n1557, u1_uk_n1558, u1_uk_n1559, u1_uk_n1565, u1_uk_n1570, u1_uk_n161, u1_uk_n162, u1_uk_n1620, 
       u1_uk_n1629, u1_uk_n163, u1_uk_n1633, u1_uk_n1643, u1_uk_n1659, u1_uk_n1660, u1_uk_n17, u1_uk_n1710, u1_uk_n1714, 
       u1_uk_n1717, u1_uk_n1720, u1_uk_n1721, u1_uk_n1729, u1_uk_n1734, u1_uk_n1744, u1_uk_n1749, u1_uk_n1802, u1_uk_n1809, 
       u1_uk_n1812, u1_uk_n1813, u1_uk_n1814, u1_uk_n1819, u1_uk_n182, u1_uk_n1840, u1_uk_n187, u1_uk_n191, u1_uk_n202, 
       u1_uk_n203, u1_uk_n207, u1_uk_n209, u1_uk_n214, u1_uk_n217, u1_uk_n220, u1_uk_n222, u1_uk_n230, u1_uk_n231, 
       u1_uk_n238, u1_uk_n242, u1_uk_n251, u1_uk_n252, u1_uk_n27, u1_uk_n271, u1_uk_n277, u1_uk_n279, u1_uk_n286, 
       u1_uk_n291, u1_uk_n292, u1_uk_n294, u1_uk_n298, u1_uk_n31, u1_uk_n60, u1_uk_n83, u1_uk_n92, u1_uk_n93, 
       u1_uk_n94, u2_K2_20, u2_K2_43, u2_K2_44, u2_K2_45, u2_K2_46, u2_K2_47, u2_K2_48, u2_K5_31, 
       u2_K5_32, u2_K5_34, u2_K5_38, u2_K5_41, u2_K8_45, u2_L0_1, u2_L0_10, u2_L0_15, u2_L0_20, 
       u2_L0_21, u2_L0_26, u2_L0_27, u2_L0_5, u2_L3_11, u2_L3_12, u2_L3_19, u2_L3_22, u2_L3_29, 
       u2_L3_32, u2_L3_4, u2_L3_7, u2_L6_15, u2_L6_21, u2_L6_27, u2_L6_5, u2_R0_1, u2_R0_12, 
       u2_R0_13, u2_R0_14, u2_R0_15, u2_R0_16, u2_R0_17, u2_R0_28, u2_R0_29, u2_R0_30, u2_R0_31, 
       u2_R0_32, u2_R3_20, u2_R3_21, u2_R3_22, u2_R3_23, u2_R3_24, u2_R3_25, u2_R3_26, u2_R3_27, 
       u2_R3_28, u2_R3_29, u2_R6_1, u2_R6_28, u2_R6_29, u2_R6_30, u2_R6_31, u2_R6_32, u2_uk_K_r0_11, 
       u2_uk_K_r0_47, u2_uk_K_r3_14, u2_uk_K_r3_16, u2_uk_K_r3_29, u2_uk_K_r3_52, u2_uk_K_r3_9, u2_uk_K_r6_0, u2_uk_K_r6_37, u2_uk_n102, 
       u2_uk_n1049, u2_uk_n1113, u2_uk_n117, u2_uk_n1234, u2_uk_n1238, u2_uk_n1243, u2_uk_n1248, u2_uk_n1249, u2_uk_n1260, 
       u2_uk_n1269, u2_uk_n128, u2_uk_n1365, u2_uk_n1376, u2_uk_n1382, u2_uk_n1383, u2_uk_n1400, u2_uk_n1401, u2_uk_n1403, 
       u2_uk_n142, u2_uk_n146, u2_uk_n147, u2_uk_n1504, u2_uk_n1511, u2_uk_n1531, u2_uk_n1532, u2_uk_n1537, u2_uk_n1538, 
       u2_uk_n155, u2_uk_n161, u2_uk_n162, u2_uk_n17, u2_uk_n182, u2_uk_n191, u2_uk_n202, u2_uk_n203, u2_uk_n217, 
       u2_uk_n222, u2_uk_n223, u2_uk_n230, u2_uk_n231, u2_uk_n31, u2_uk_n60, u2_uk_n63, u2_uk_n92, u2_uk_n94, u0_N164, u0_N174, u0_N180, u0_N186, u0_N420, u0_N422, u0_N424, u0_N427, u0_N430, 
        u0_N432, u0_N436, u0_N437, u0_N438, u0_N442, u0_N446, u0_N447, u0_N449, u0_N453, 
        u0_N456, u0_N460, u0_N463, u0_N464, u0_N465, u0_N470, u0_N471, u0_N475, u0_N477, 
        u0_N478, u0_uk_n163, u0_uk_n188, u0_uk_n231, u0_uk_n83, u0_uk_n93, u1_N103, u1_N109, u1_N120, 
        u1_N128, u1_N137, u1_N147, u1_N153, u1_N224, u1_N233, u1_N243, u1_N249, u1_N288, 
        u1_N297, u1_N307, u1_N313, u1_N354, u1_N359, u1_N365, u1_N376, u1_N416, u1_N425, 
        u1_N435, u1_N441, u1_N68, u1_N70, u1_N75, u1_N78, u1_N84, u1_N85, u1_N90, 
        u1_N95, u1_N98, u2_N131, u2_N134, u2_N138, u2_N139, u2_N146, u2_N149, u2_N156, 
        u2_N159, u2_N228, u2_N238, u2_N244, u2_N250, u2_N32, u2_N36, u2_N41, u2_N46, 
        u2_N51, u2_N52, u2_N57, u2_N58 );
  input u0_K14_4, u0_K14_42, u0_K14_46, u0_K15_18, u0_L12_12, u0_L12_15, u0_L12_17, u0_L12_21, u0_L12_22, 
        u0_L12_23, u0_L12_27, u0_L12_31, u0_L12_32, u0_L12_5, u0_L12_7, u0_L12_9, u0_L13_13, u0_L13_16, 
        u0_L13_17, u0_L13_18, u0_L13_2, u0_L13_23, u0_L13_24, u0_L13_28, u0_L13_30, u0_L13_31, u0_L13_6, 
        u0_L13_9, u0_L4_15, u0_L4_21, u0_L4_27, u0_L4_5, u0_R12_1, u0_R12_2, u0_R12_24, u0_R12_25, 
        u0_R12_26, u0_R12_27, u0_R12_28, u0_R12_29, u0_R12_3, u0_R12_30, u0_R12_31, u0_R12_32, u0_R12_4, 
        u0_R12_5, u0_R13_1, u0_R13_10, u0_R13_11, u0_R13_12, u0_R13_13, u0_R13_2, u0_R13_3, u0_R13_32, 
        u0_R13_4, u0_R13_5, u0_R13_6, u0_R13_7, u0_R13_8, u0_R13_9, u0_R4_1, u0_R4_28, u0_R4_29, 
        u0_R4_30, u0_R4_31, u0_R4_32, u0_uk_K_r12_10, u0_uk_K_r12_15, u0_uk_K_r12_16, u0_uk_K_r12_21, u0_uk_K_r12_47, u0_uk_K_r13_13, 
        u0_uk_K_r13_17, u0_uk_K_r13_19, u0_uk_K_r13_25, u0_uk_K_r13_32, u0_uk_K_r13_4, u0_uk_K_r13_55, u0_uk_K_r4_23, u0_uk_n1, u0_uk_n10, 
        u0_uk_n100, u0_uk_n109, u0_uk_n11, u0_uk_n110, u0_uk_n117, u0_uk_n118, u0_uk_n128, u0_uk_n14, u0_uk_n141, 
        u0_uk_n146, u0_uk_n15, u0_uk_n155, u0_uk_n16, u0_uk_n17, u0_uk_n187, u0_uk_n19, u0_uk_n20, u0_uk_n203, 
        u0_uk_n208, u0_uk_n213, u0_uk_n214, u0_uk_n217, u0_uk_n220, u0_uk_n222, u0_uk_n230, u0_uk_n24, u0_uk_n240, 
        u0_uk_n242, u0_uk_n25, u0_uk_n250, u0_uk_n251, u0_uk_n252, u0_uk_n26, u0_uk_n27, u0_uk_n29, u0_uk_n30, 
        u0_uk_n35, u0_uk_n36, u0_uk_n37, u0_uk_n38, u0_uk_n411, u0_uk_n412, u0_uk_n417, u0_uk_n418, u0_uk_n425, 
        u0_uk_n429, u0_uk_n43, u0_uk_n430, u0_uk_n434, u0_uk_n439, u0_uk_n44, u0_uk_n445, u0_uk_n450, u0_uk_n46, 
        u0_uk_n52, u0_uk_n56, u0_uk_n57, u0_uk_n58, u0_uk_n59, u0_uk_n6, u0_uk_n60, u0_uk_n62, u0_uk_n63, 
        u0_uk_n64, u0_uk_n65, u0_uk_n67, u0_uk_n68, u0_uk_n73, u0_uk_n75, u0_uk_n77, u0_uk_n78, u0_uk_n8, 
        u0_uk_n80, u0_uk_n81, u0_uk_n82, u0_uk_n85, u0_uk_n90, u0_uk_n92, u0_uk_n94, u1_L10_14, u1_L10_25, 
        u1_L10_3, u1_L10_8, u1_L12_1, u1_L12_10, u1_L12_20, u1_L12_26, u1_L1_12, u1_L1_15, u1_L1_21, 
        u1_L1_22, u1_L1_27, u1_L1_32, u1_L1_5, u1_L1_7, u1_L2_14, u1_L2_25, u1_L2_3, u1_L2_8, 
        u1_L3_1, u1_L3_10, u1_L3_20, u1_L3_26, u1_L6_1, u1_L6_10, u1_L6_20, u1_L6_26, u1_L8_1, 
        u1_L8_10, u1_L8_20, u1_L8_26, u1_R10_16, u1_R10_17, u1_R10_18, u1_R10_19, u1_R10_20, u1_R10_21, 
        u1_R12_12, u1_R12_13, u1_R12_14, u1_R12_15, u1_R12_16, u1_R12_17, u1_R1_1, u1_R1_24, u1_R1_25, 
        u1_R1_26, u1_R1_27, u1_R1_28, u1_R1_29, u1_R1_30, u1_R1_31, u1_R1_32, u1_R2_16, u1_R2_17, 
        u1_R2_18, u1_R2_19, u1_R2_20, u1_R2_21, u1_R3_12, u1_R3_13, u1_R3_14, u1_R3_15, u1_R3_16, 
        u1_R3_17, u1_R6_12, u1_R6_13, u1_R6_14, u1_R6_15, u1_R6_16, u1_R6_17, u1_R8_12, u1_R8_13, 
        u1_R8_14, u1_R8_15, u1_R8_16, u1_R8_17, u1_uk_K_r10_23, u1_uk_K_r10_42, u1_uk_K_r12_25, u1_uk_K_r12_33, u1_uk_K_r12_41, 
        u1_uk_K_r1_15, u1_uk_K_r1_16, u1_uk_K_r1_21, u1_uk_K_r1_22, u1_uk_K_r2_16, u1_uk_K_r2_21, u1_uk_K_r2_28, u1_uk_K_r2_31, u1_uk_K_r2_36, 
        u1_uk_K_r2_49, u1_uk_K_r2_7, u1_uk_K_r3_24, u1_uk_K_r3_33, u1_uk_K_r3_47, u1_uk_K_r8_13, u1_uk_K_r8_19, u1_uk_K_r8_27, u1_uk_K_r8_40, 
        u1_uk_K_r8_5, u1_uk_n10, u1_uk_n100, u1_uk_n102, u1_uk_n109, u1_uk_n11, u1_uk_n117, u1_uk_n118, u1_uk_n128, 
        u1_uk_n1307, u1_uk_n1313, u1_uk_n1314, u1_uk_n1318, u1_uk_n1322, u1_uk_n1327, u1_uk_n1328, u1_uk_n1330, u1_uk_n1334, 
        u1_uk_n1335, u1_uk_n1338, u1_uk_n1342, u1_uk_n1350, u1_uk_n1375, u1_uk_n1376, u1_uk_n1381, u1_uk_n1398, u1_uk_n1402, 
        u1_uk_n1409, u1_uk_n1415, u1_uk_n142, u1_uk_n1424, u1_uk_n1427, u1_uk_n1429, u1_uk_n1435, u1_uk_n145, u1_uk_n146, 
        u1_uk_n147, u1_uk_n148, u1_uk_n1530, u1_uk_n1538, u1_uk_n1543, u1_uk_n1545, u1_uk_n1548, u1_uk_n155, u1_uk_n1551, 
        u1_uk_n1552, u1_uk_n1557, u1_uk_n1558, u1_uk_n1559, u1_uk_n1565, u1_uk_n1570, u1_uk_n161, u1_uk_n162, u1_uk_n1620, 
        u1_uk_n1629, u1_uk_n163, u1_uk_n1633, u1_uk_n1643, u1_uk_n1659, u1_uk_n1660, u1_uk_n17, u1_uk_n1710, u1_uk_n1714, 
        u1_uk_n1717, u1_uk_n1720, u1_uk_n1721, u1_uk_n1729, u1_uk_n1734, u1_uk_n1744, u1_uk_n1749, u1_uk_n1802, u1_uk_n1809, 
        u1_uk_n1812, u1_uk_n1813, u1_uk_n1814, u1_uk_n1819, u1_uk_n182, u1_uk_n1840, u1_uk_n187, u1_uk_n191, u1_uk_n202, 
        u1_uk_n203, u1_uk_n207, u1_uk_n209, u1_uk_n214, u1_uk_n217, u1_uk_n220, u1_uk_n222, u1_uk_n230, u1_uk_n231, 
        u1_uk_n238, u1_uk_n242, u1_uk_n251, u1_uk_n252, u1_uk_n27, u1_uk_n271, u1_uk_n277, u1_uk_n279, u1_uk_n286, 
        u1_uk_n291, u1_uk_n292, u1_uk_n294, u1_uk_n298, u1_uk_n31, u1_uk_n60, u1_uk_n83, u1_uk_n92, u1_uk_n93, 
        u1_uk_n94, u2_K2_20, u2_K2_43, u2_K2_44, u2_K2_45, u2_K2_46, u2_K2_47, u2_K2_48, u2_K5_31, 
        u2_K5_32, u2_K5_34, u2_K5_38, u2_K5_41, u2_K8_45, u2_L0_1, u2_L0_10, u2_L0_15, u2_L0_20, 
        u2_L0_21, u2_L0_26, u2_L0_27, u2_L0_5, u2_L3_11, u2_L3_12, u2_L3_19, u2_L3_22, u2_L3_29, 
        u2_L3_32, u2_L3_4, u2_L3_7, u2_L6_15, u2_L6_21, u2_L6_27, u2_L6_5, u2_R0_1, u2_R0_12, 
        u2_R0_13, u2_R0_14, u2_R0_15, u2_R0_16, u2_R0_17, u2_R0_28, u2_R0_29, u2_R0_30, u2_R0_31, 
        u2_R0_32, u2_R3_20, u2_R3_21, u2_R3_22, u2_R3_23, u2_R3_24, u2_R3_25, u2_R3_26, u2_R3_27, 
        u2_R3_28, u2_R3_29, u2_R6_1, u2_R6_28, u2_R6_29, u2_R6_30, u2_R6_31, u2_R6_32, u2_uk_K_r0_11, 
        u2_uk_K_r0_47, u2_uk_K_r3_14, u2_uk_K_r3_16, u2_uk_K_r3_29, u2_uk_K_r3_52, u2_uk_K_r3_9, u2_uk_K_r6_0, u2_uk_K_r6_37, u2_uk_n102, 
        u2_uk_n1049, u2_uk_n1113, u2_uk_n117, u2_uk_n1234, u2_uk_n1238, u2_uk_n1243, u2_uk_n1248, u2_uk_n1249, u2_uk_n1260, 
        u2_uk_n1269, u2_uk_n128, u2_uk_n1365, u2_uk_n1376, u2_uk_n1382, u2_uk_n1383, u2_uk_n1400, u2_uk_n1401, u2_uk_n1403, 
        u2_uk_n142, u2_uk_n146, u2_uk_n147, u2_uk_n1504, u2_uk_n1511, u2_uk_n1531, u2_uk_n1532, u2_uk_n1537, u2_uk_n1538, 
        u2_uk_n155, u2_uk_n161, u2_uk_n162, u2_uk_n17, u2_uk_n182, u2_uk_n191, u2_uk_n202, u2_uk_n203, u2_uk_n217, 
        u2_uk_n222, u2_uk_n223, u2_uk_n230, u2_uk_n231, u2_uk_n31, u2_uk_n60, u2_uk_n63, u2_uk_n92, u2_uk_n94;
  output u0_N164, u0_N174, u0_N180, u0_N186, u0_N420, u0_N422, u0_N424, u0_N427, u0_N430, 
        u0_N432, u0_N436, u0_N437, u0_N438, u0_N442, u0_N446, u0_N447, u0_N449, u0_N453, 
        u0_N456, u0_N460, u0_N463, u0_N464, u0_N465, u0_N470, u0_N471, u0_N475, u0_N477, 
        u0_N478, u0_uk_n163, u0_uk_n188, u0_uk_n231, u0_uk_n83, u0_uk_n93, u1_N103, u1_N109, u1_N120, 
        u1_N128, u1_N137, u1_N147, u1_N153, u1_N224, u1_N233, u1_N243, u1_N249, u1_N288, 
        u1_N297, u1_N307, u1_N313, u1_N354, u1_N359, u1_N365, u1_N376, u1_N416, u1_N425, 
        u1_N435, u1_N441, u1_N68, u1_N70, u1_N75, u1_N78, u1_N84, u1_N85, u1_N90, 
        u1_N95, u1_N98, u2_N131, u2_N134, u2_N138, u2_N139, u2_N146, u2_N149, u2_N156, 
        u2_N159, u2_N228, u2_N238, u2_N244, u2_N250, u2_N32, u2_N36, u2_N41, u2_N46, 
        u2_N51, u2_N52, u2_N57, u2_N58;
  wire u0_K14_1, u0_K14_2, u0_K14_3, u0_K14_37, u0_K14_38, u0_K14_39, u0_K14_40, u0_K14_41, u0_K14_43, 
       u0_K14_44, u0_K14_45, u0_K14_47, u0_K14_48, u0_K14_5, u0_K14_6, u0_K15_1, u0_K15_10, u0_K15_11, 
       u0_K15_12, u0_K15_13, u0_K15_14, u0_K15_15, u0_K15_16, u0_K15_17, u0_K15_2, u0_K15_3, u0_K15_4, 
       u0_K15_5, u0_K15_6, u0_K15_7, u0_K15_8, u0_K15_9, u0_K6_43, u0_K6_44, u0_K6_45, u0_K6_46, 
       u0_K6_47, u0_K6_48, u0_out13_12, u0_out13_15, u0_out13_17, u0_out13_21, u0_out13_22, u0_out13_23, u0_out13_27, 
       u0_out13_31, u0_out13_32, u0_out13_5, u0_out13_7, u0_out13_9, u0_out14_13, u0_out14_16, u0_out14_17, u0_out14_18, 
       u0_out14_2, u0_out14_23, u0_out14_24, u0_out14_28, u0_out14_30, u0_out14_31, u0_out14_6, u0_out14_9, u0_out5_15, 
       u0_out5_21, u0_out5_27, u0_out5_5, u0_u13_X_1, u0_u13_X_2, u0_u13_X_3, u0_u13_X_37, u0_u13_X_38, u0_u13_X_39, 
       u0_u13_X_4, u0_u13_X_40, u0_u13_X_41, u0_u13_X_42, u0_u13_X_43, u0_u13_X_44, u0_u13_X_45, u0_u13_X_46, u0_u13_X_47, 
       u0_u13_X_48, u0_u13_X_5, u0_u13_X_6, u0_u13_u0_n100, u0_u13_u0_n101, u0_u13_u0_n102, u0_u13_u0_n103, u0_u13_u0_n104, u0_u13_u0_n105, 
       u0_u13_u0_n106, u0_u13_u0_n107, u0_u13_u0_n108, u0_u13_u0_n109, u0_u13_u0_n110, u0_u13_u0_n111, u0_u13_u0_n112, u0_u13_u0_n113, u0_u13_u0_n114, 
       u0_u13_u0_n115, u0_u13_u0_n116, u0_u13_u0_n117, u0_u13_u0_n118, u0_u13_u0_n119, u0_u13_u0_n120, u0_u13_u0_n121, u0_u13_u0_n122, u0_u13_u0_n123, 
       u0_u13_u0_n124, u0_u13_u0_n125, u0_u13_u0_n126, u0_u13_u0_n127, u0_u13_u0_n128, u0_u13_u0_n129, u0_u13_u0_n130, u0_u13_u0_n131, u0_u13_u0_n132, 
       u0_u13_u0_n133, u0_u13_u0_n134, u0_u13_u0_n135, u0_u13_u0_n136, u0_u13_u0_n137, u0_u13_u0_n138, u0_u13_u0_n139, u0_u13_u0_n140, u0_u13_u0_n141, 
       u0_u13_u0_n142, u0_u13_u0_n143, u0_u13_u0_n144, u0_u13_u0_n145, u0_u13_u0_n146, u0_u13_u0_n147, u0_u13_u0_n148, u0_u13_u0_n149, u0_u13_u0_n150, 
       u0_u13_u0_n151, u0_u13_u0_n152, u0_u13_u0_n153, u0_u13_u0_n154, u0_u13_u0_n155, u0_u13_u0_n156, u0_u13_u0_n157, u0_u13_u0_n158, u0_u13_u0_n159, 
       u0_u13_u0_n160, u0_u13_u0_n161, u0_u13_u0_n162, u0_u13_u0_n163, u0_u13_u0_n164, u0_u13_u0_n165, u0_u13_u0_n166, u0_u13_u0_n167, u0_u13_u0_n168, 
       u0_u13_u0_n169, u0_u13_u0_n170, u0_u13_u0_n171, u0_u13_u0_n172, u0_u13_u0_n173, u0_u13_u0_n174, u0_u13_u0_n88, u0_u13_u0_n89, u0_u13_u0_n90, 
       u0_u13_u0_n91, u0_u13_u0_n92, u0_u13_u0_n93, u0_u13_u0_n94, u0_u13_u0_n95, u0_u13_u0_n96, u0_u13_u0_n97, u0_u13_u0_n98, u0_u13_u0_n99, 
       u0_u13_u6_n100, u0_u13_u6_n101, u0_u13_u6_n102, u0_u13_u6_n103, u0_u13_u6_n104, u0_u13_u6_n105, u0_u13_u6_n106, u0_u13_u6_n107, u0_u13_u6_n108, 
       u0_u13_u6_n109, u0_u13_u6_n110, u0_u13_u6_n111, u0_u13_u6_n112, u0_u13_u6_n113, u0_u13_u6_n114, u0_u13_u6_n115, u0_u13_u6_n116, u0_u13_u6_n117, 
       u0_u13_u6_n118, u0_u13_u6_n119, u0_u13_u6_n120, u0_u13_u6_n121, u0_u13_u6_n122, u0_u13_u6_n123, u0_u13_u6_n124, u0_u13_u6_n125, u0_u13_u6_n126, 
       u0_u13_u6_n127, u0_u13_u6_n128, u0_u13_u6_n129, u0_u13_u6_n130, u0_u13_u6_n131, u0_u13_u6_n132, u0_u13_u6_n133, u0_u13_u6_n134, u0_u13_u6_n135, 
       u0_u13_u6_n136, u0_u13_u6_n137, u0_u13_u6_n138, u0_u13_u6_n139, u0_u13_u6_n140, u0_u13_u6_n141, u0_u13_u6_n142, u0_u13_u6_n143, u0_u13_u6_n144, 
       u0_u13_u6_n145, u0_u13_u6_n146, u0_u13_u6_n147, u0_u13_u6_n148, u0_u13_u6_n149, u0_u13_u6_n150, u0_u13_u6_n151, u0_u13_u6_n152, u0_u13_u6_n153, 
       u0_u13_u6_n154, u0_u13_u6_n155, u0_u13_u6_n156, u0_u13_u6_n157, u0_u13_u6_n158, u0_u13_u6_n159, u0_u13_u6_n160, u0_u13_u6_n161, u0_u13_u6_n162, 
       u0_u13_u6_n163, u0_u13_u6_n164, u0_u13_u6_n165, u0_u13_u6_n166, u0_u13_u6_n167, u0_u13_u6_n168, u0_u13_u6_n169, u0_u13_u6_n170, u0_u13_u6_n171, 
       u0_u13_u6_n172, u0_u13_u6_n173, u0_u13_u6_n174, u0_u13_u6_n88, u0_u13_u6_n89, u0_u13_u6_n90, u0_u13_u6_n91, u0_u13_u6_n92, u0_u13_u6_n93, 
       u0_u13_u6_n94, u0_u13_u6_n95, u0_u13_u6_n96, u0_u13_u6_n97, u0_u13_u6_n98, u0_u13_u6_n99, u0_u13_u7_n100, u0_u13_u7_n101, u0_u13_u7_n102, 
       u0_u13_u7_n103, u0_u13_u7_n104, u0_u13_u7_n105, u0_u13_u7_n106, u0_u13_u7_n107, u0_u13_u7_n108, u0_u13_u7_n109, u0_u13_u7_n110, u0_u13_u7_n111, 
       u0_u13_u7_n112, u0_u13_u7_n113, u0_u13_u7_n114, u0_u13_u7_n115, u0_u13_u7_n116, u0_u13_u7_n117, u0_u13_u7_n118, u0_u13_u7_n119, u0_u13_u7_n120, 
       u0_u13_u7_n121, u0_u13_u7_n122, u0_u13_u7_n123, u0_u13_u7_n124, u0_u13_u7_n125, u0_u13_u7_n126, u0_u13_u7_n127, u0_u13_u7_n128, u0_u13_u7_n129, 
       u0_u13_u7_n130, u0_u13_u7_n131, u0_u13_u7_n132, u0_u13_u7_n133, u0_u13_u7_n134, u0_u13_u7_n135, u0_u13_u7_n136, u0_u13_u7_n137, u0_u13_u7_n138, 
       u0_u13_u7_n139, u0_u13_u7_n140, u0_u13_u7_n141, u0_u13_u7_n142, u0_u13_u7_n143, u0_u13_u7_n144, u0_u13_u7_n145, u0_u13_u7_n146, u0_u13_u7_n147, 
       u0_u13_u7_n148, u0_u13_u7_n149, u0_u13_u7_n150, u0_u13_u7_n151, u0_u13_u7_n152, u0_u13_u7_n153, u0_u13_u7_n154, u0_u13_u7_n155, u0_u13_u7_n156, 
       u0_u13_u7_n157, u0_u13_u7_n158, u0_u13_u7_n159, u0_u13_u7_n160, u0_u13_u7_n161, u0_u13_u7_n162, u0_u13_u7_n163, u0_u13_u7_n164, u0_u13_u7_n165, 
       u0_u13_u7_n166, u0_u13_u7_n167, u0_u13_u7_n168, u0_u13_u7_n169, u0_u13_u7_n170, u0_u13_u7_n171, u0_u13_u7_n172, u0_u13_u7_n173, u0_u13_u7_n174, 
       u0_u13_u7_n175, u0_u13_u7_n176, u0_u13_u7_n177, u0_u13_u7_n178, u0_u13_u7_n179, u0_u13_u7_n180, u0_u13_u7_n91, u0_u13_u7_n92, u0_u13_u7_n93, 
       u0_u13_u7_n94, u0_u13_u7_n95, u0_u13_u7_n96, u0_u13_u7_n97, u0_u13_u7_n98, u0_u13_u7_n99, u0_u14_X_1, u0_u14_X_10, u0_u14_X_11, 
       u0_u14_X_12, u0_u14_X_13, u0_u14_X_14, u0_u14_X_15, u0_u14_X_16, u0_u14_X_17, u0_u14_X_18, u0_u14_X_2, u0_u14_X_3, 
       u0_u14_X_4, u0_u14_X_5, u0_u14_X_6, u0_u14_X_7, u0_u14_X_8, u0_u14_X_9, u0_u14_u0_n100, u0_u14_u0_n101, u0_u14_u0_n102, 
       u0_u14_u0_n103, u0_u14_u0_n104, u0_u14_u0_n105, u0_u14_u0_n106, u0_u14_u0_n107, u0_u14_u0_n108, u0_u14_u0_n109, u0_u14_u0_n110, u0_u14_u0_n111, 
       u0_u14_u0_n112, u0_u14_u0_n113, u0_u14_u0_n114, u0_u14_u0_n115, u0_u14_u0_n116, u0_u14_u0_n117, u0_u14_u0_n118, u0_u14_u0_n119, u0_u14_u0_n120, 
       u0_u14_u0_n121, u0_u14_u0_n122, u0_u14_u0_n123, u0_u14_u0_n124, u0_u14_u0_n125, u0_u14_u0_n126, u0_u14_u0_n127, u0_u14_u0_n128, u0_u14_u0_n129, 
       u0_u14_u0_n130, u0_u14_u0_n131, u0_u14_u0_n132, u0_u14_u0_n133, u0_u14_u0_n134, u0_u14_u0_n135, u0_u14_u0_n136, u0_u14_u0_n137, u0_u14_u0_n138, 
       u0_u14_u0_n139, u0_u14_u0_n140, u0_u14_u0_n141, u0_u14_u0_n142, u0_u14_u0_n143, u0_u14_u0_n144, u0_u14_u0_n145, u0_u14_u0_n146, u0_u14_u0_n147, 
       u0_u14_u0_n148, u0_u14_u0_n149, u0_u14_u0_n150, u0_u14_u0_n151, u0_u14_u0_n152, u0_u14_u0_n153, u0_u14_u0_n154, u0_u14_u0_n155, u0_u14_u0_n156, 
       u0_u14_u0_n157, u0_u14_u0_n158, u0_u14_u0_n159, u0_u14_u0_n160, u0_u14_u0_n161, u0_u14_u0_n162, u0_u14_u0_n163, u0_u14_u0_n164, u0_u14_u0_n165, 
       u0_u14_u0_n166, u0_u14_u0_n167, u0_u14_u0_n168, u0_u14_u0_n169, u0_u14_u0_n170, u0_u14_u0_n171, u0_u14_u0_n172, u0_u14_u0_n173, u0_u14_u0_n174, 
       u0_u14_u0_n88, u0_u14_u0_n89, u0_u14_u0_n90, u0_u14_u0_n91, u0_u14_u0_n92, u0_u14_u0_n93, u0_u14_u0_n94, u0_u14_u0_n95, u0_u14_u0_n96, 
       u0_u14_u0_n97, u0_u14_u0_n98, u0_u14_u0_n99, u0_u14_u1_n100, u0_u14_u1_n101, u0_u14_u1_n102, u0_u14_u1_n103, u0_u14_u1_n104, u0_u14_u1_n105, 
       u0_u14_u1_n106, u0_u14_u1_n107, u0_u14_u1_n108, u0_u14_u1_n109, u0_u14_u1_n110, u0_u14_u1_n111, u0_u14_u1_n112, u0_u14_u1_n113, u0_u14_u1_n114, 
       u0_u14_u1_n115, u0_u14_u1_n116, u0_u14_u1_n117, u0_u14_u1_n118, u0_u14_u1_n119, u0_u14_u1_n120, u0_u14_u1_n121, u0_u14_u1_n122, u0_u14_u1_n123, 
       u0_u14_u1_n124, u0_u14_u1_n125, u0_u14_u1_n126, u0_u14_u1_n127, u0_u14_u1_n128, u0_u14_u1_n129, u0_u14_u1_n130, u0_u14_u1_n131, u0_u14_u1_n132, 
       u0_u14_u1_n133, u0_u14_u1_n134, u0_u14_u1_n135, u0_u14_u1_n136, u0_u14_u1_n137, u0_u14_u1_n138, u0_u14_u1_n139, u0_u14_u1_n140, u0_u14_u1_n141, 
       u0_u14_u1_n142, u0_u14_u1_n143, u0_u14_u1_n144, u0_u14_u1_n145, u0_u14_u1_n146, u0_u14_u1_n147, u0_u14_u1_n148, u0_u14_u1_n149, u0_u14_u1_n150, 
       u0_u14_u1_n151, u0_u14_u1_n152, u0_u14_u1_n153, u0_u14_u1_n154, u0_u14_u1_n155, u0_u14_u1_n156, u0_u14_u1_n157, u0_u14_u1_n158, u0_u14_u1_n159, 
       u0_u14_u1_n160, u0_u14_u1_n161, u0_u14_u1_n162, u0_u14_u1_n163, u0_u14_u1_n164, u0_u14_u1_n165, u0_u14_u1_n166, u0_u14_u1_n167, u0_u14_u1_n168, 
       u0_u14_u1_n169, u0_u14_u1_n170, u0_u14_u1_n171, u0_u14_u1_n172, u0_u14_u1_n173, u0_u14_u1_n174, u0_u14_u1_n175, u0_u14_u1_n176, u0_u14_u1_n177, 
       u0_u14_u1_n178, u0_u14_u1_n179, u0_u14_u1_n180, u0_u14_u1_n181, u0_u14_u1_n182, u0_u14_u1_n183, u0_u14_u1_n184, u0_u14_u1_n185, u0_u14_u1_n186, 
       u0_u14_u1_n187, u0_u14_u1_n188, u0_u14_u1_n95, u0_u14_u1_n96, u0_u14_u1_n97, u0_u14_u1_n98, u0_u14_u1_n99, u0_u14_u2_n100, u0_u14_u2_n101, 
       u0_u14_u2_n102, u0_u14_u2_n103, u0_u14_u2_n104, u0_u14_u2_n105, u0_u14_u2_n106, u0_u14_u2_n107, u0_u14_u2_n108, u0_u14_u2_n109, u0_u14_u2_n110, 
       u0_u14_u2_n111, u0_u14_u2_n112, u0_u14_u2_n113, u0_u14_u2_n114, u0_u14_u2_n115, u0_u14_u2_n116, u0_u14_u2_n117, u0_u14_u2_n118, u0_u14_u2_n119, 
       u0_u14_u2_n120, u0_u14_u2_n121, u0_u14_u2_n122, u0_u14_u2_n123, u0_u14_u2_n124, u0_u14_u2_n125, u0_u14_u2_n126, u0_u14_u2_n127, u0_u14_u2_n128, 
       u0_u14_u2_n129, u0_u14_u2_n130, u0_u14_u2_n131, u0_u14_u2_n132, u0_u14_u2_n133, u0_u14_u2_n134, u0_u14_u2_n135, u0_u14_u2_n136, u0_u14_u2_n137, 
       u0_u14_u2_n138, u0_u14_u2_n139, u0_u14_u2_n140, u0_u14_u2_n141, u0_u14_u2_n142, u0_u14_u2_n143, u0_u14_u2_n144, u0_u14_u2_n145, u0_u14_u2_n146, 
       u0_u14_u2_n147, u0_u14_u2_n148, u0_u14_u2_n149, u0_u14_u2_n150, u0_u14_u2_n151, u0_u14_u2_n152, u0_u14_u2_n153, u0_u14_u2_n154, u0_u14_u2_n155, 
       u0_u14_u2_n156, u0_u14_u2_n157, u0_u14_u2_n158, u0_u14_u2_n159, u0_u14_u2_n160, u0_u14_u2_n161, u0_u14_u2_n162, u0_u14_u2_n163, u0_u14_u2_n164, 
       u0_u14_u2_n165, u0_u14_u2_n166, u0_u14_u2_n167, u0_u14_u2_n168, u0_u14_u2_n169, u0_u14_u2_n170, u0_u14_u2_n171, u0_u14_u2_n172, u0_u14_u2_n173, 
       u0_u14_u2_n174, u0_u14_u2_n175, u0_u14_u2_n176, u0_u14_u2_n177, u0_u14_u2_n178, u0_u14_u2_n179, u0_u14_u2_n180, u0_u14_u2_n181, u0_u14_u2_n182, 
       u0_u14_u2_n183, u0_u14_u2_n184, u0_u14_u2_n185, u0_u14_u2_n186, u0_u14_u2_n187, u0_u14_u2_n188, u0_u14_u2_n95, u0_u14_u2_n96, u0_u14_u2_n97, 
       u0_u14_u2_n98, u0_u14_u2_n99, u0_u5_X_43, u0_u5_X_44, u0_u5_X_45, u0_u5_X_46, u0_u5_X_47, u0_u5_X_48, u0_u5_u7_n100, 
       u0_u5_u7_n101, u0_u5_u7_n102, u0_u5_u7_n103, u0_u5_u7_n104, u0_u5_u7_n105, u0_u5_u7_n106, u0_u5_u7_n107, u0_u5_u7_n108, u0_u5_u7_n109, 
       u0_u5_u7_n110, u0_u5_u7_n111, u0_u5_u7_n112, u0_u5_u7_n113, u0_u5_u7_n114, u0_u5_u7_n115, u0_u5_u7_n116, u0_u5_u7_n117, u0_u5_u7_n118, 
       u0_u5_u7_n119, u0_u5_u7_n120, u0_u5_u7_n121, u0_u5_u7_n122, u0_u5_u7_n123, u0_u5_u7_n124, u0_u5_u7_n125, u0_u5_u7_n126, u0_u5_u7_n127, 
       u0_u5_u7_n128, u0_u5_u7_n129, u0_u5_u7_n130, u0_u5_u7_n131, u0_u5_u7_n132, u0_u5_u7_n133, u0_u5_u7_n134, u0_u5_u7_n135, u0_u5_u7_n136, 
       u0_u5_u7_n137, u0_u5_u7_n138, u0_u5_u7_n139, u0_u5_u7_n140, u0_u5_u7_n141, u0_u5_u7_n142, u0_u5_u7_n143, u0_u5_u7_n144, u0_u5_u7_n145, 
       u0_u5_u7_n146, u0_u5_u7_n147, u0_u5_u7_n148, u0_u5_u7_n149, u0_u5_u7_n150, u0_u5_u7_n151, u0_u5_u7_n152, u0_u5_u7_n153, u0_u5_u7_n154, 
       u0_u5_u7_n155, u0_u5_u7_n156, u0_u5_u7_n157, u0_u5_u7_n158, u0_u5_u7_n159, u0_u5_u7_n160, u0_u5_u7_n161, u0_u5_u7_n162, u0_u5_u7_n163, 
       u0_u5_u7_n164, u0_u5_u7_n165, u0_u5_u7_n166, u0_u5_u7_n167, u0_u5_u7_n168, u0_u5_u7_n169, u0_u5_u7_n170, u0_u5_u7_n171, u0_u5_u7_n172, 
       u0_u5_u7_n173, u0_u5_u7_n174, u0_u5_u7_n175, u0_u5_u7_n176, u0_u5_u7_n177, u0_u5_u7_n178, u0_u5_u7_n179, u0_u5_u7_n180, u0_u5_u7_n91, 
       u0_u5_u7_n92, u0_u5_u7_n93, u0_u5_u7_n94, u0_u5_u7_n95, u0_u5_u7_n96, u0_u5_u7_n97, u0_u5_u7_n98, u0_u5_u7_n99, u0_uk_n789, 
       u0_uk_n912, u0_uk_n913, u0_uk_n922, u0_uk_n923, u0_uk_n924, u0_uk_n925, u0_uk_n927, u0_uk_n929, u0_uk_n930, 
       u0_uk_n931, u0_uk_n932, u1_K10_19, u1_K10_20, u1_K10_21, u1_K10_22, u1_K10_23, u1_K10_24, u1_K12_25, 
       u1_K12_26, u1_K12_27, u1_K12_28, u1_K12_29, u1_K12_30, u1_K14_19, u1_K14_20, u1_K14_21, u1_K14_22, 
       u1_K14_23, u1_K14_24, u1_K3_37, u1_K3_38, u1_K3_39, u1_K3_40, u1_K3_41, u1_K3_42, u1_K3_43, 
       u1_K3_44, u1_K3_45, u1_K3_46, u1_K3_47, u1_K3_48, u1_K4_25, u1_K4_26, u1_K4_27, u1_K4_28, 
       u1_K4_29, u1_K4_30, u1_K5_19, u1_K5_20, u1_K5_21, u1_K5_22, u1_K5_23, u1_K5_24, u1_K8_19, 
       u1_K8_20, u1_K8_21, u1_K8_22, u1_K8_23, u1_K8_24, u1_out11_14, u1_out11_25, u1_out11_3, u1_out11_8, 
       u1_out13_1, u1_out13_10, u1_out13_20, u1_out13_26, u1_out2_12, u1_out2_15, u1_out2_21, u1_out2_22, u1_out2_27, 
       u1_out2_32, u1_out2_5, u1_out2_7, u1_out3_14, u1_out3_25, u1_out3_3, u1_out3_8, u1_out4_1, u1_out4_10, 
       u1_out4_20, u1_out4_26, u1_out7_1, u1_out7_10, u1_out7_20, u1_out7_26, u1_out9_1, u1_out9_10, u1_out9_20, 
       u1_out9_26, u1_u11_X_25, u1_u11_X_26, u1_u11_X_27, u1_u11_X_28, u1_u11_X_29, u1_u11_X_30, u1_u11_u4_n100, u1_u11_u4_n101, 
       u1_u11_u4_n102, u1_u11_u4_n103, u1_u11_u4_n104, u1_u11_u4_n105, u1_u11_u4_n106, u1_u11_u4_n107, u1_u11_u4_n108, u1_u11_u4_n109, u1_u11_u4_n110, 
       u1_u11_u4_n111, u1_u11_u4_n112, u1_u11_u4_n113, u1_u11_u4_n114, u1_u11_u4_n115, u1_u11_u4_n116, u1_u11_u4_n117, u1_u11_u4_n118, u1_u11_u4_n119, 
       u1_u11_u4_n120, u1_u11_u4_n121, u1_u11_u4_n122, u1_u11_u4_n123, u1_u11_u4_n124, u1_u11_u4_n125, u1_u11_u4_n126, u1_u11_u4_n127, u1_u11_u4_n128, 
       u1_u11_u4_n129, u1_u11_u4_n130, u1_u11_u4_n131, u1_u11_u4_n132, u1_u11_u4_n133, u1_u11_u4_n134, u1_u11_u4_n135, u1_u11_u4_n136, u1_u11_u4_n137, 
       u1_u11_u4_n138, u1_u11_u4_n139, u1_u11_u4_n140, u1_u11_u4_n141, u1_u11_u4_n142, u1_u11_u4_n143, u1_u11_u4_n144, u1_u11_u4_n145, u1_u11_u4_n146, 
       u1_u11_u4_n147, u1_u11_u4_n148, u1_u11_u4_n149, u1_u11_u4_n150, u1_u11_u4_n151, u1_u11_u4_n152, u1_u11_u4_n153, u1_u11_u4_n154, u1_u11_u4_n155, 
       u1_u11_u4_n156, u1_u11_u4_n157, u1_u11_u4_n158, u1_u11_u4_n159, u1_u11_u4_n160, u1_u11_u4_n161, u1_u11_u4_n162, u1_u11_u4_n163, u1_u11_u4_n164, 
       u1_u11_u4_n165, u1_u11_u4_n166, u1_u11_u4_n167, u1_u11_u4_n168, u1_u11_u4_n169, u1_u11_u4_n170, u1_u11_u4_n171, u1_u11_u4_n172, u1_u11_u4_n173, 
       u1_u11_u4_n174, u1_u11_u4_n175, u1_u11_u4_n176, u1_u11_u4_n177, u1_u11_u4_n178, u1_u11_u4_n179, u1_u11_u4_n180, u1_u11_u4_n181, u1_u11_u4_n182, 
       u1_u11_u4_n183, u1_u11_u4_n184, u1_u11_u4_n185, u1_u11_u4_n186, u1_u11_u4_n94, u1_u11_u4_n95, u1_u11_u4_n96, u1_u11_u4_n97, u1_u11_u4_n98, 
       u1_u11_u4_n99, u1_u13_X_19, u1_u13_X_20, u1_u13_X_21, u1_u13_X_22, u1_u13_X_23, u1_u13_X_24, u1_u13_u3_n100, u1_u13_u3_n101, 
       u1_u13_u3_n102, u1_u13_u3_n103, u1_u13_u3_n104, u1_u13_u3_n105, u1_u13_u3_n106, u1_u13_u3_n107, u1_u13_u3_n108, u1_u13_u3_n109, u1_u13_u3_n110, 
       u1_u13_u3_n111, u1_u13_u3_n112, u1_u13_u3_n113, u1_u13_u3_n114, u1_u13_u3_n115, u1_u13_u3_n116, u1_u13_u3_n117, u1_u13_u3_n118, u1_u13_u3_n119, 
       u1_u13_u3_n120, u1_u13_u3_n121, u1_u13_u3_n122, u1_u13_u3_n123, u1_u13_u3_n124, u1_u13_u3_n125, u1_u13_u3_n126, u1_u13_u3_n127, u1_u13_u3_n128, 
       u1_u13_u3_n129, u1_u13_u3_n130, u1_u13_u3_n131, u1_u13_u3_n132, u1_u13_u3_n133, u1_u13_u3_n134, u1_u13_u3_n135, u1_u13_u3_n136, u1_u13_u3_n137, 
       u1_u13_u3_n138, u1_u13_u3_n139, u1_u13_u3_n140, u1_u13_u3_n141, u1_u13_u3_n142, u1_u13_u3_n143, u1_u13_u3_n144, u1_u13_u3_n145, u1_u13_u3_n146, 
       u1_u13_u3_n147, u1_u13_u3_n148, u1_u13_u3_n149, u1_u13_u3_n150, u1_u13_u3_n151, u1_u13_u3_n152, u1_u13_u3_n153, u1_u13_u3_n154, u1_u13_u3_n155, 
       u1_u13_u3_n156, u1_u13_u3_n157, u1_u13_u3_n158, u1_u13_u3_n159, u1_u13_u3_n160, u1_u13_u3_n161, u1_u13_u3_n162, u1_u13_u3_n163, u1_u13_u3_n164, 
       u1_u13_u3_n165, u1_u13_u3_n166, u1_u13_u3_n167, u1_u13_u3_n168, u1_u13_u3_n169, u1_u13_u3_n170, u1_u13_u3_n171, u1_u13_u3_n172, u1_u13_u3_n173, 
       u1_u13_u3_n174, u1_u13_u3_n175, u1_u13_u3_n176, u1_u13_u3_n177, u1_u13_u3_n178, u1_u13_u3_n179, u1_u13_u3_n180, u1_u13_u3_n181, u1_u13_u3_n182, 
       u1_u13_u3_n183, u1_u13_u3_n184, u1_u13_u3_n185, u1_u13_u3_n186, u1_u13_u3_n94, u1_u13_u3_n95, u1_u13_u3_n96, u1_u13_u3_n97, u1_u13_u3_n98, 
       u1_u13_u3_n99, u1_u2_X_37, u1_u2_X_38, u1_u2_X_39, u1_u2_X_40, u1_u2_X_41, u1_u2_X_42, u1_u2_X_43, u1_u2_X_44, 
       u1_u2_X_45, u1_u2_X_46, u1_u2_X_47, u1_u2_X_48, u1_u2_u6_n100, u1_u2_u6_n101, u1_u2_u6_n102, u1_u2_u6_n103, u1_u2_u6_n104, 
       u1_u2_u6_n105, u1_u2_u6_n106, u1_u2_u6_n107, u1_u2_u6_n108, u1_u2_u6_n109, u1_u2_u6_n110, u1_u2_u6_n111, u1_u2_u6_n112, u1_u2_u6_n113, 
       u1_u2_u6_n114, u1_u2_u6_n115, u1_u2_u6_n116, u1_u2_u6_n117, u1_u2_u6_n118, u1_u2_u6_n119, u1_u2_u6_n120, u1_u2_u6_n121, u1_u2_u6_n122, 
       u1_u2_u6_n123, u1_u2_u6_n124, u1_u2_u6_n125, u1_u2_u6_n126, u1_u2_u6_n127, u1_u2_u6_n128, u1_u2_u6_n129, u1_u2_u6_n130, u1_u2_u6_n131, 
       u1_u2_u6_n132, u1_u2_u6_n133, u1_u2_u6_n134, u1_u2_u6_n135, u1_u2_u6_n136, u1_u2_u6_n137, u1_u2_u6_n138, u1_u2_u6_n139, u1_u2_u6_n140, 
       u1_u2_u6_n141, u1_u2_u6_n142, u1_u2_u6_n143, u1_u2_u6_n144, u1_u2_u6_n145, u1_u2_u6_n146, u1_u2_u6_n147, u1_u2_u6_n148, u1_u2_u6_n149, 
       u1_u2_u6_n150, u1_u2_u6_n151, u1_u2_u6_n152, u1_u2_u6_n153, u1_u2_u6_n154, u1_u2_u6_n155, u1_u2_u6_n156, u1_u2_u6_n157, u1_u2_u6_n158, 
       u1_u2_u6_n159, u1_u2_u6_n160, u1_u2_u6_n161, u1_u2_u6_n162, u1_u2_u6_n163, u1_u2_u6_n164, u1_u2_u6_n165, u1_u2_u6_n166, u1_u2_u6_n167, 
       u1_u2_u6_n168, u1_u2_u6_n169, u1_u2_u6_n170, u1_u2_u6_n171, u1_u2_u6_n172, u1_u2_u6_n173, u1_u2_u6_n174, u1_u2_u6_n88, u1_u2_u6_n89, 
       u1_u2_u6_n90, u1_u2_u6_n91, u1_u2_u6_n92, u1_u2_u6_n93, u1_u2_u6_n94, u1_u2_u6_n95, u1_u2_u6_n96, u1_u2_u6_n97, u1_u2_u6_n98, 
       u1_u2_u6_n99, u1_u2_u7_n100, u1_u2_u7_n101, u1_u2_u7_n102, u1_u2_u7_n103, u1_u2_u7_n104, u1_u2_u7_n105, u1_u2_u7_n106, u1_u2_u7_n107, 
       u1_u2_u7_n108, u1_u2_u7_n109, u1_u2_u7_n110, u1_u2_u7_n111, u1_u2_u7_n112, u1_u2_u7_n113, u1_u2_u7_n114, u1_u2_u7_n115, u1_u2_u7_n116, 
       u1_u2_u7_n117, u1_u2_u7_n118, u1_u2_u7_n119, u1_u2_u7_n120, u1_u2_u7_n121, u1_u2_u7_n122, u1_u2_u7_n123, u1_u2_u7_n124, u1_u2_u7_n125, 
       u1_u2_u7_n126, u1_u2_u7_n127, u1_u2_u7_n128, u1_u2_u7_n129, u1_u2_u7_n130, u1_u2_u7_n131, u1_u2_u7_n132, u1_u2_u7_n133, u1_u2_u7_n134, 
       u1_u2_u7_n135, u1_u2_u7_n136, u1_u2_u7_n137, u1_u2_u7_n138, u1_u2_u7_n139, u1_u2_u7_n140, u1_u2_u7_n141, u1_u2_u7_n142, u1_u2_u7_n143, 
       u1_u2_u7_n144, u1_u2_u7_n145, u1_u2_u7_n146, u1_u2_u7_n147, u1_u2_u7_n148, u1_u2_u7_n149, u1_u2_u7_n150, u1_u2_u7_n151, u1_u2_u7_n152, 
       u1_u2_u7_n153, u1_u2_u7_n154, u1_u2_u7_n155, u1_u2_u7_n156, u1_u2_u7_n157, u1_u2_u7_n158, u1_u2_u7_n159, u1_u2_u7_n160, u1_u2_u7_n161, 
       u1_u2_u7_n162, u1_u2_u7_n163, u1_u2_u7_n164, u1_u2_u7_n165, u1_u2_u7_n166, u1_u2_u7_n167, u1_u2_u7_n168, u1_u2_u7_n169, u1_u2_u7_n170, 
       u1_u2_u7_n171, u1_u2_u7_n172, u1_u2_u7_n173, u1_u2_u7_n174, u1_u2_u7_n175, u1_u2_u7_n176, u1_u2_u7_n177, u1_u2_u7_n178, u1_u2_u7_n179, 
       u1_u2_u7_n180, u1_u2_u7_n91, u1_u2_u7_n92, u1_u2_u7_n93, u1_u2_u7_n94, u1_u2_u7_n95, u1_u2_u7_n96, u1_u2_u7_n97, u1_u2_u7_n98, 
       u1_u2_u7_n99, u1_u3_X_25, u1_u3_X_26, u1_u3_X_27, u1_u3_X_28, u1_u3_X_29, u1_u3_X_30, u1_u3_u4_n100, u1_u3_u4_n101, 
       u1_u3_u4_n102, u1_u3_u4_n103, u1_u3_u4_n104, u1_u3_u4_n105, u1_u3_u4_n106, u1_u3_u4_n107, u1_u3_u4_n108, u1_u3_u4_n109, u1_u3_u4_n110, 
       u1_u3_u4_n111, u1_u3_u4_n112, u1_u3_u4_n113, u1_u3_u4_n114, u1_u3_u4_n115, u1_u3_u4_n116, u1_u3_u4_n117, u1_u3_u4_n118, u1_u3_u4_n119, 
       u1_u3_u4_n120, u1_u3_u4_n121, u1_u3_u4_n122, u1_u3_u4_n123, u1_u3_u4_n124, u1_u3_u4_n125, u1_u3_u4_n126, u1_u3_u4_n127, u1_u3_u4_n128, 
       u1_u3_u4_n129, u1_u3_u4_n130, u1_u3_u4_n131, u1_u3_u4_n132, u1_u3_u4_n133, u1_u3_u4_n134, u1_u3_u4_n135, u1_u3_u4_n136, u1_u3_u4_n137, 
       u1_u3_u4_n138, u1_u3_u4_n139, u1_u3_u4_n140, u1_u3_u4_n141, u1_u3_u4_n142, u1_u3_u4_n143, u1_u3_u4_n144, u1_u3_u4_n145, u1_u3_u4_n146, 
       u1_u3_u4_n147, u1_u3_u4_n148, u1_u3_u4_n149, u1_u3_u4_n150, u1_u3_u4_n151, u1_u3_u4_n152, u1_u3_u4_n153, u1_u3_u4_n154, u1_u3_u4_n155, 
       u1_u3_u4_n156, u1_u3_u4_n157, u1_u3_u4_n158, u1_u3_u4_n159, u1_u3_u4_n160, u1_u3_u4_n161, u1_u3_u4_n162, u1_u3_u4_n163, u1_u3_u4_n164, 
       u1_u3_u4_n165, u1_u3_u4_n166, u1_u3_u4_n167, u1_u3_u4_n168, u1_u3_u4_n169, u1_u3_u4_n170, u1_u3_u4_n171, u1_u3_u4_n172, u1_u3_u4_n173, 
       u1_u3_u4_n174, u1_u3_u4_n175, u1_u3_u4_n176, u1_u3_u4_n177, u1_u3_u4_n178, u1_u3_u4_n179, u1_u3_u4_n180, u1_u3_u4_n181, u1_u3_u4_n182, 
       u1_u3_u4_n183, u1_u3_u4_n184, u1_u3_u4_n185, u1_u3_u4_n186, u1_u3_u4_n94, u1_u3_u4_n95, u1_u3_u4_n96, u1_u3_u4_n97, u1_u3_u4_n98, 
       u1_u3_u4_n99, u1_u4_X_19, u1_u4_X_20, u1_u4_X_21, u1_u4_X_22, u1_u4_X_23, u1_u4_X_24, u1_u4_u3_n100, u1_u4_u3_n101, 
       u1_u4_u3_n102, u1_u4_u3_n103, u1_u4_u3_n104, u1_u4_u3_n105, u1_u4_u3_n106, u1_u4_u3_n107, u1_u4_u3_n108, u1_u4_u3_n109, u1_u4_u3_n110, 
       u1_u4_u3_n111, u1_u4_u3_n112, u1_u4_u3_n113, u1_u4_u3_n114, u1_u4_u3_n115, u1_u4_u3_n116, u1_u4_u3_n117, u1_u4_u3_n118, u1_u4_u3_n119, 
       u1_u4_u3_n120, u1_u4_u3_n121, u1_u4_u3_n122, u1_u4_u3_n123, u1_u4_u3_n124, u1_u4_u3_n125, u1_u4_u3_n126, u1_u4_u3_n127, u1_u4_u3_n128, 
       u1_u4_u3_n129, u1_u4_u3_n130, u1_u4_u3_n131, u1_u4_u3_n132, u1_u4_u3_n133, u1_u4_u3_n134, u1_u4_u3_n135, u1_u4_u3_n136, u1_u4_u3_n137, 
       u1_u4_u3_n138, u1_u4_u3_n139, u1_u4_u3_n140, u1_u4_u3_n141, u1_u4_u3_n142, u1_u4_u3_n143, u1_u4_u3_n144, u1_u4_u3_n145, u1_u4_u3_n146, 
       u1_u4_u3_n147, u1_u4_u3_n148, u1_u4_u3_n149, u1_u4_u3_n150, u1_u4_u3_n151, u1_u4_u3_n152, u1_u4_u3_n153, u1_u4_u3_n154, u1_u4_u3_n155, 
       u1_u4_u3_n156, u1_u4_u3_n157, u1_u4_u3_n158, u1_u4_u3_n159, u1_u4_u3_n160, u1_u4_u3_n161, u1_u4_u3_n162, u1_u4_u3_n163, u1_u4_u3_n164, 
       u1_u4_u3_n165, u1_u4_u3_n166, u1_u4_u3_n167, u1_u4_u3_n168, u1_u4_u3_n169, u1_u4_u3_n170, u1_u4_u3_n171, u1_u4_u3_n172, u1_u4_u3_n173, 
       u1_u4_u3_n174, u1_u4_u3_n175, u1_u4_u3_n176, u1_u4_u3_n177, u1_u4_u3_n178, u1_u4_u3_n179, u1_u4_u3_n180, u1_u4_u3_n181, u1_u4_u3_n182, 
       u1_u4_u3_n183, u1_u4_u3_n184, u1_u4_u3_n185, u1_u4_u3_n186, u1_u4_u3_n94, u1_u4_u3_n95, u1_u4_u3_n96, u1_u4_u3_n97, u1_u4_u3_n98, 
       u1_u4_u3_n99, u1_u7_X_19, u1_u7_X_20, u1_u7_X_21, u1_u7_X_22, u1_u7_X_23, u1_u7_X_24, u1_u7_u3_n100, u1_u7_u3_n101, 
       u1_u7_u3_n102, u1_u7_u3_n103, u1_u7_u3_n104, u1_u7_u3_n105, u1_u7_u3_n106, u1_u7_u3_n107, u1_u7_u3_n108, u1_u7_u3_n109, u1_u7_u3_n110, 
       u1_u7_u3_n111, u1_u7_u3_n112, u1_u7_u3_n113, u1_u7_u3_n114, u1_u7_u3_n115, u1_u7_u3_n116, u1_u7_u3_n117, u1_u7_u3_n118, u1_u7_u3_n119, 
       u1_u7_u3_n120, u1_u7_u3_n121, u1_u7_u3_n122, u1_u7_u3_n123, u1_u7_u3_n124, u1_u7_u3_n125, u1_u7_u3_n126, u1_u7_u3_n127, u1_u7_u3_n128, 
       u1_u7_u3_n129, u1_u7_u3_n130, u1_u7_u3_n131, u1_u7_u3_n132, u1_u7_u3_n133, u1_u7_u3_n134, u1_u7_u3_n135, u1_u7_u3_n136, u1_u7_u3_n137, 
       u1_u7_u3_n138, u1_u7_u3_n139, u1_u7_u3_n140, u1_u7_u3_n141, u1_u7_u3_n142, u1_u7_u3_n143, u1_u7_u3_n144, u1_u7_u3_n145, u1_u7_u3_n146, 
       u1_u7_u3_n147, u1_u7_u3_n148, u1_u7_u3_n149, u1_u7_u3_n150, u1_u7_u3_n151, u1_u7_u3_n152, u1_u7_u3_n153, u1_u7_u3_n154, u1_u7_u3_n155, 
       u1_u7_u3_n156, u1_u7_u3_n157, u1_u7_u3_n158, u1_u7_u3_n159, u1_u7_u3_n160, u1_u7_u3_n161, u1_u7_u3_n162, u1_u7_u3_n163, u1_u7_u3_n164, 
       u1_u7_u3_n165, u1_u7_u3_n166, u1_u7_u3_n167, u1_u7_u3_n168, u1_u7_u3_n169, u1_u7_u3_n170, u1_u7_u3_n171, u1_u7_u3_n172, u1_u7_u3_n173, 
       u1_u7_u3_n174, u1_u7_u3_n175, u1_u7_u3_n176, u1_u7_u3_n177, u1_u7_u3_n178, u1_u7_u3_n179, u1_u7_u3_n180, u1_u7_u3_n181, u1_u7_u3_n182, 
       u1_u7_u3_n183, u1_u7_u3_n184, u1_u7_u3_n185, u1_u7_u3_n186, u1_u7_u3_n94, u1_u7_u3_n95, u1_u7_u3_n96, u1_u7_u3_n97, u1_u7_u3_n98, 
       u1_u7_u3_n99, u1_u9_X_19, u1_u9_X_20, u1_u9_X_21, u1_u9_X_22, u1_u9_X_23, u1_u9_X_24, u1_u9_u3_n100, u1_u9_u3_n101, 
       u1_u9_u3_n102, u1_u9_u3_n103, u1_u9_u3_n104, u1_u9_u3_n105, u1_u9_u3_n106, u1_u9_u3_n107, u1_u9_u3_n108, u1_u9_u3_n109, u1_u9_u3_n110, 
       u1_u9_u3_n111, u1_u9_u3_n112, u1_u9_u3_n113, u1_u9_u3_n114, u1_u9_u3_n115, u1_u9_u3_n116, u1_u9_u3_n117, u1_u9_u3_n118, u1_u9_u3_n119, 
       u1_u9_u3_n120, u1_u9_u3_n121, u1_u9_u3_n122, u1_u9_u3_n123, u1_u9_u3_n124, u1_u9_u3_n125, u1_u9_u3_n126, u1_u9_u3_n127, u1_u9_u3_n128, 
       u1_u9_u3_n129, u1_u9_u3_n130, u1_u9_u3_n131, u1_u9_u3_n132, u1_u9_u3_n133, u1_u9_u3_n134, u1_u9_u3_n135, u1_u9_u3_n136, u1_u9_u3_n137, 
       u1_u9_u3_n138, u1_u9_u3_n139, u1_u9_u3_n140, u1_u9_u3_n141, u1_u9_u3_n142, u1_u9_u3_n143, u1_u9_u3_n144, u1_u9_u3_n145, u1_u9_u3_n146, 
       u1_u9_u3_n147, u1_u9_u3_n148, u1_u9_u3_n149, u1_u9_u3_n150, u1_u9_u3_n151, u1_u9_u3_n152, u1_u9_u3_n153, u1_u9_u3_n154, u1_u9_u3_n155, 
       u1_u9_u3_n156, u1_u9_u3_n157, u1_u9_u3_n158, u1_u9_u3_n159, u1_u9_u3_n160, u1_u9_u3_n161, u1_u9_u3_n162, u1_u9_u3_n163, u1_u9_u3_n164, 
       u1_u9_u3_n165, u1_u9_u3_n166, u1_u9_u3_n167, u1_u9_u3_n168, u1_u9_u3_n169, u1_u9_u3_n170, u1_u9_u3_n171, u1_u9_u3_n172, u1_u9_u3_n173, 
       u1_u9_u3_n174, u1_u9_u3_n175, u1_u9_u3_n176, u1_u9_u3_n177, u1_u9_u3_n178, u1_u9_u3_n179, u1_u9_u3_n180, u1_u9_u3_n181, u1_u9_u3_n182, 
       u1_u9_u3_n183, u1_u9_u3_n184, u1_u9_u3_n185, u1_u9_u3_n186, u1_u9_u3_n94, u1_u9_u3_n95, u1_u9_u3_n96, u1_u9_u3_n97, u1_u9_u3_n98, 
       u1_u9_u3_n99, u1_uk_n1044, u1_uk_n1045, u1_uk_n1046, u1_uk_n1047, u1_uk_n1057, u1_uk_n1058, u1_uk_n1059, u1_uk_n1060, 
       u1_uk_n1062, u1_uk_n1073, u1_uk_n1074, u1_uk_n308, u1_uk_n312, u1_uk_n313, u1_uk_n319, u1_uk_n526, u1_uk_n951, 
       u1_uk_n952, u2_K2_19, u2_K2_21, u2_K2_22, u2_K2_23, u2_K2_24, u2_K5_33, u2_K5_35, u2_K5_36, 
       u2_K5_37, u2_K5_39, u2_K5_40, u2_K5_42, u2_K8_43, u2_K8_44, u2_K8_46, u2_K8_47, u2_K8_48, 
       u2_out1_1, u2_out1_10, u2_out1_15, u2_out1_20, u2_out1_21, u2_out1_26, u2_out1_27, u2_out1_5, u2_out4_11, 
       u2_out4_12, u2_out4_19, u2_out4_22, u2_out4_29, u2_out4_32, u2_out4_4, u2_out4_7, u2_out7_15, u2_out7_21, 
       u2_out7_27, u2_out7_5, u2_u1_X_19, u2_u1_X_20, u2_u1_X_21, u2_u1_X_22, u2_u1_X_23, u2_u1_X_24, u2_u1_X_43, 
       u2_u1_X_44, u2_u1_X_45, u2_u1_X_46, u2_u1_X_47, u2_u1_X_48, u2_u1_u3_n100, u2_u1_u3_n101, u2_u1_u3_n102, u2_u1_u3_n103, 
       u2_u1_u3_n104, u2_u1_u3_n105, u2_u1_u3_n106, u2_u1_u3_n107, u2_u1_u3_n108, u2_u1_u3_n109, u2_u1_u3_n110, u2_u1_u3_n111, u2_u1_u3_n112, 
       u2_u1_u3_n113, u2_u1_u3_n114, u2_u1_u3_n115, u2_u1_u3_n116, u2_u1_u3_n117, u2_u1_u3_n118, u2_u1_u3_n119, u2_u1_u3_n120, u2_u1_u3_n121, 
       u2_u1_u3_n122, u2_u1_u3_n123, u2_u1_u3_n124, u2_u1_u3_n125, u2_u1_u3_n126, u2_u1_u3_n127, u2_u1_u3_n128, u2_u1_u3_n129, u2_u1_u3_n130, 
       u2_u1_u3_n131, u2_u1_u3_n132, u2_u1_u3_n133, u2_u1_u3_n134, u2_u1_u3_n135, u2_u1_u3_n136, u2_u1_u3_n137, u2_u1_u3_n138, u2_u1_u3_n139, 
       u2_u1_u3_n140, u2_u1_u3_n141, u2_u1_u3_n142, u2_u1_u3_n143, u2_u1_u3_n144, u2_u1_u3_n145, u2_u1_u3_n146, u2_u1_u3_n147, u2_u1_u3_n148, 
       u2_u1_u3_n149, u2_u1_u3_n150, u2_u1_u3_n151, u2_u1_u3_n152, u2_u1_u3_n153, u2_u1_u3_n154, u2_u1_u3_n155, u2_u1_u3_n156, u2_u1_u3_n157, 
       u2_u1_u3_n158, u2_u1_u3_n159, u2_u1_u3_n160, u2_u1_u3_n161, u2_u1_u3_n162, u2_u1_u3_n163, u2_u1_u3_n164, u2_u1_u3_n165, u2_u1_u3_n166, 
       u2_u1_u3_n167, u2_u1_u3_n168, u2_u1_u3_n169, u2_u1_u3_n170, u2_u1_u3_n171, u2_u1_u3_n172, u2_u1_u3_n173, u2_u1_u3_n174, u2_u1_u3_n175, 
       u2_u1_u3_n176, u2_u1_u3_n177, u2_u1_u3_n178, u2_u1_u3_n179, u2_u1_u3_n180, u2_u1_u3_n181, u2_u1_u3_n182, u2_u1_u3_n183, u2_u1_u3_n184, 
       u2_u1_u3_n185, u2_u1_u3_n186, u2_u1_u3_n94, u2_u1_u3_n95, u2_u1_u3_n96, u2_u1_u3_n97, u2_u1_u3_n98, u2_u1_u3_n99, u2_u1_u7_n100, 
       u2_u1_u7_n101, u2_u1_u7_n102, u2_u1_u7_n103, u2_u1_u7_n104, u2_u1_u7_n105, u2_u1_u7_n106, u2_u1_u7_n107, u2_u1_u7_n108, u2_u1_u7_n109, 
       u2_u1_u7_n110, u2_u1_u7_n111, u2_u1_u7_n112, u2_u1_u7_n113, u2_u1_u7_n114, u2_u1_u7_n115, u2_u1_u7_n116, u2_u1_u7_n117, u2_u1_u7_n118, 
       u2_u1_u7_n119, u2_u1_u7_n120, u2_u1_u7_n121, u2_u1_u7_n122, u2_u1_u7_n123, u2_u1_u7_n124, u2_u1_u7_n125, u2_u1_u7_n126, u2_u1_u7_n127, 
       u2_u1_u7_n128, u2_u1_u7_n129, u2_u1_u7_n130, u2_u1_u7_n131, u2_u1_u7_n132, u2_u1_u7_n133, u2_u1_u7_n134, u2_u1_u7_n135, u2_u1_u7_n136, 
       u2_u1_u7_n137, u2_u1_u7_n138, u2_u1_u7_n139, u2_u1_u7_n140, u2_u1_u7_n141, u2_u1_u7_n142, u2_u1_u7_n143, u2_u1_u7_n144, u2_u1_u7_n145, 
       u2_u1_u7_n146, u2_u1_u7_n147, u2_u1_u7_n148, u2_u1_u7_n149, u2_u1_u7_n150, u2_u1_u7_n151, u2_u1_u7_n152, u2_u1_u7_n153, u2_u1_u7_n154, 
       u2_u1_u7_n155, u2_u1_u7_n156, u2_u1_u7_n157, u2_u1_u7_n158, u2_u1_u7_n159, u2_u1_u7_n160, u2_u1_u7_n161, u2_u1_u7_n162, u2_u1_u7_n163, 
       u2_u1_u7_n164, u2_u1_u7_n165, u2_u1_u7_n166, u2_u1_u7_n167, u2_u1_u7_n168, u2_u1_u7_n169, u2_u1_u7_n170, u2_u1_u7_n171, u2_u1_u7_n172, 
       u2_u1_u7_n173, u2_u1_u7_n174, u2_u1_u7_n175, u2_u1_u7_n176, u2_u1_u7_n177, u2_u1_u7_n178, u2_u1_u7_n179, u2_u1_u7_n180, u2_u1_u7_n91, 
       u2_u1_u7_n92, u2_u1_u7_n93, u2_u1_u7_n94, u2_u1_u7_n95, u2_u1_u7_n96, u2_u1_u7_n97, u2_u1_u7_n98, u2_u1_u7_n99, u2_u4_X_31, 
       u2_u4_X_32, u2_u4_X_33, u2_u4_X_34, u2_u4_X_35, u2_u4_X_36, u2_u4_X_37, u2_u4_X_38, u2_u4_X_39, u2_u4_X_40, 
       u2_u4_X_41, u2_u4_X_42, u2_u4_u5_n100, u2_u4_u5_n101, u2_u4_u5_n102, u2_u4_u5_n103, u2_u4_u5_n104, u2_u4_u5_n105, u2_u4_u5_n106, 
       u2_u4_u5_n107, u2_u4_u5_n108, u2_u4_u5_n109, u2_u4_u5_n110, u2_u4_u5_n111, u2_u4_u5_n112, u2_u4_u5_n113, u2_u4_u5_n114, u2_u4_u5_n115, 
       u2_u4_u5_n116, u2_u4_u5_n117, u2_u4_u5_n118, u2_u4_u5_n119, u2_u4_u5_n120, u2_u4_u5_n121, u2_u4_u5_n122, u2_u4_u5_n123, u2_u4_u5_n124, 
       u2_u4_u5_n125, u2_u4_u5_n126, u2_u4_u5_n127, u2_u4_u5_n128, u2_u4_u5_n129, u2_u4_u5_n130, u2_u4_u5_n131, u2_u4_u5_n132, u2_u4_u5_n133, 
       u2_u4_u5_n134, u2_u4_u5_n135, u2_u4_u5_n136, u2_u4_u5_n137, u2_u4_u5_n138, u2_u4_u5_n139, u2_u4_u5_n140, u2_u4_u5_n141, u2_u4_u5_n142, 
       u2_u4_u5_n143, u2_u4_u5_n144, u2_u4_u5_n145, u2_u4_u5_n146, u2_u4_u5_n147, u2_u4_u5_n148, u2_u4_u5_n149, u2_u4_u5_n150, u2_u4_u5_n151, 
       u2_u4_u5_n152, u2_u4_u5_n153, u2_u4_u5_n154, u2_u4_u5_n155, u2_u4_u5_n156, u2_u4_u5_n157, u2_u4_u5_n158, u2_u4_u5_n159, u2_u4_u5_n160, 
       u2_u4_u5_n161, u2_u4_u5_n162, u2_u4_u5_n163, u2_u4_u5_n164, u2_u4_u5_n165, u2_u4_u5_n166, u2_u4_u5_n167, u2_u4_u5_n168, u2_u4_u5_n169, 
       u2_u4_u5_n170, u2_u4_u5_n171, u2_u4_u5_n172, u2_u4_u5_n173, u2_u4_u5_n174, u2_u4_u5_n175, u2_u4_u5_n176, u2_u4_u5_n177, u2_u4_u5_n178, 
       u2_u4_u5_n179, u2_u4_u5_n180, u2_u4_u5_n181, u2_u4_u5_n182, u2_u4_u5_n183, u2_u4_u5_n184, u2_u4_u5_n185, u2_u4_u5_n186, u2_u4_u5_n187, 
       u2_u4_u5_n188, u2_u4_u5_n189, u2_u4_u5_n190, u2_u4_u5_n191, u2_u4_u5_n192, u2_u4_u5_n193, u2_u4_u5_n194, u2_u4_u5_n195, u2_u4_u5_n196, 
       u2_u4_u5_n99, u2_u4_u6_n100, u2_u4_u6_n101, u2_u4_u6_n102, u2_u4_u6_n103, u2_u4_u6_n104, u2_u4_u6_n105, u2_u4_u6_n106, u2_u4_u6_n107, 
       u2_u4_u6_n108, u2_u4_u6_n109, u2_u4_u6_n110, u2_u4_u6_n111, u2_u4_u6_n112, u2_u4_u6_n113, u2_u4_u6_n114, u2_u4_u6_n115, u2_u4_u6_n116, 
       u2_u4_u6_n117, u2_u4_u6_n118, u2_u4_u6_n119, u2_u4_u6_n120, u2_u4_u6_n121, u2_u4_u6_n122, u2_u4_u6_n123, u2_u4_u6_n124, u2_u4_u6_n125, 
       u2_u4_u6_n126, u2_u4_u6_n127, u2_u4_u6_n128, u2_u4_u6_n129, u2_u4_u6_n130, u2_u4_u6_n131, u2_u4_u6_n132, u2_u4_u6_n133, u2_u4_u6_n134, 
       u2_u4_u6_n135, u2_u4_u6_n136, u2_u4_u6_n137, u2_u4_u6_n138, u2_u4_u6_n139, u2_u4_u6_n140, u2_u4_u6_n141, u2_u4_u6_n142, u2_u4_u6_n143, 
       u2_u4_u6_n144, u2_u4_u6_n145, u2_u4_u6_n146, u2_u4_u6_n147, u2_u4_u6_n148, u2_u4_u6_n149, u2_u4_u6_n150, u2_u4_u6_n151, u2_u4_u6_n152, 
       u2_u4_u6_n153, u2_u4_u6_n154, u2_u4_u6_n155, u2_u4_u6_n156, u2_u4_u6_n157, u2_u4_u6_n158, u2_u4_u6_n159, u2_u4_u6_n160, u2_u4_u6_n161, 
       u2_u4_u6_n162, u2_u4_u6_n163, u2_u4_u6_n164, u2_u4_u6_n165, u2_u4_u6_n166, u2_u4_u6_n167, u2_u4_u6_n168, u2_u4_u6_n169, u2_u4_u6_n170, 
       u2_u4_u6_n171, u2_u4_u6_n172, u2_u4_u6_n173, u2_u4_u6_n174, u2_u4_u6_n88, u2_u4_u6_n89, u2_u4_u6_n90, u2_u4_u6_n91, u2_u4_u6_n92, 
       u2_u4_u6_n93, u2_u4_u6_n94, u2_u4_u6_n95, u2_u4_u6_n96, u2_u4_u6_n97, u2_u4_u6_n98, u2_u4_u6_n99, u2_u7_X_43, u2_u7_X_44, 
       u2_u7_X_45, u2_u7_X_46, u2_u7_X_47, u2_u7_X_48, u2_u7_u7_n100, u2_u7_u7_n101, u2_u7_u7_n102, u2_u7_u7_n103, u2_u7_u7_n104, 
       u2_u7_u7_n105, u2_u7_u7_n106, u2_u7_u7_n107, u2_u7_u7_n108, u2_u7_u7_n109, u2_u7_u7_n110, u2_u7_u7_n111, u2_u7_u7_n112, u2_u7_u7_n113, 
       u2_u7_u7_n114, u2_u7_u7_n115, u2_u7_u7_n116, u2_u7_u7_n117, u2_u7_u7_n118, u2_u7_u7_n119, u2_u7_u7_n120, u2_u7_u7_n121, u2_u7_u7_n122, 
       u2_u7_u7_n123, u2_u7_u7_n124, u2_u7_u7_n125, u2_u7_u7_n126, u2_u7_u7_n127, u2_u7_u7_n128, u2_u7_u7_n129, u2_u7_u7_n130, u2_u7_u7_n131, 
       u2_u7_u7_n132, u2_u7_u7_n133, u2_u7_u7_n134, u2_u7_u7_n135, u2_u7_u7_n136, u2_u7_u7_n137, u2_u7_u7_n138, u2_u7_u7_n139, u2_u7_u7_n140, 
       u2_u7_u7_n141, u2_u7_u7_n142, u2_u7_u7_n143, u2_u7_u7_n144, u2_u7_u7_n145, u2_u7_u7_n146, u2_u7_u7_n147, u2_u7_u7_n148, u2_u7_u7_n149, 
       u2_u7_u7_n150, u2_u7_u7_n151, u2_u7_u7_n152, u2_u7_u7_n153, u2_u7_u7_n154, u2_u7_u7_n155, u2_u7_u7_n156, u2_u7_u7_n157, u2_u7_u7_n158, 
       u2_u7_u7_n159, u2_u7_u7_n160, u2_u7_u7_n161, u2_u7_u7_n162, u2_u7_u7_n163, u2_u7_u7_n164, u2_u7_u7_n165, u2_u7_u7_n166, u2_u7_u7_n167, 
       u2_u7_u7_n168, u2_u7_u7_n169, u2_u7_u7_n170, u2_u7_u7_n171, u2_u7_u7_n172, u2_u7_u7_n173, u2_u7_u7_n174, u2_u7_u7_n175, u2_u7_u7_n176, 
       u2_u7_u7_n177, u2_u7_u7_n178, u2_u7_u7_n179, u2_u7_u7_n180, u2_u7_u7_n91, u2_u7_u7_n92, u2_u7_u7_n93, u2_u7_u7_n94, u2_u7_u7_n95, 
       u2_u7_u7_n96, u2_u7_u7_n97, u2_u7_u7_n98, u2_u7_u7_n99, u2_uk_n1048, u2_uk_n1050, u2_uk_n1051, u2_uk_n1052, u2_uk_n1114, 
       u2_uk_n1115,  u2_uk_n995;
  XOR2_X1 u0_U100 (.B( u0_L12_27 ) , .Z( u0_N442 ) , .A( u0_out13_27 ) );
  XOR2_X1 u0_U105 (.B( u0_L12_23 ) , .Z( u0_N438 ) , .A( u0_out13_23 ) );
  XOR2_X1 u0_U106 (.B( u0_L12_22 ) , .Z( u0_N437 ) , .A( u0_out13_22 ) );
  XOR2_X1 u0_U107 (.B( u0_L12_21 ) , .Z( u0_N436 ) , .A( u0_out13_21 ) );
  XOR2_X1 u0_U111 (.B( u0_L12_17 ) , .Z( u0_N432 ) , .A( u0_out13_17 ) );
  XOR2_X1 u0_U113 (.B( u0_L12_15 ) , .Z( u0_N430 ) , .A( u0_out13_15 ) );
  XOR2_X1 u0_U117 (.B( u0_L12_12 ) , .Z( u0_N427 ) , .A( u0_out13_12 ) );
  XOR2_X1 u0_U120 (.B( u0_L12_9 ) , .Z( u0_N424 ) , .A( u0_out13_9 ) );
  XOR2_X1 u0_U122 (.B( u0_L12_7 ) , .Z( u0_N422 ) , .A( u0_out13_7 ) );
  XOR2_X1 u0_U124 (.B( u0_L12_5 ) , .Z( u0_N420 ) , .A( u0_out13_5 ) );
  XOR2_X1 u0_U385 (.B( u0_L4_27 ) , .Z( u0_N186 ) , .A( u0_out5_27 ) );
  XOR2_X1 u0_U391 (.B( u0_L4_21 ) , .Z( u0_N180 ) , .A( u0_out5_21 ) );
  XOR2_X1 u0_U398 (.B( u0_L4_15 ) , .Z( u0_N174 ) , .A( u0_out5_15 ) );
  XOR2_X1 u0_U409 (.B( u0_L4_5 ) , .Z( u0_N164 ) , .A( u0_out5_5 ) );
  XOR2_X1 u0_U61 (.B( u0_L13_31 ) , .Z( u0_N478 ) , .A( u0_out14_31 ) );
  XOR2_X1 u0_U62 (.B( u0_L13_30 ) , .Z( u0_N477 ) , .A( u0_out14_30 ) );
  XOR2_X1 u0_U64 (.B( u0_L13_28 ) , .Z( u0_N475 ) , .A( u0_out14_28 ) );
  XOR2_X1 u0_U68 (.B( u0_L13_24 ) , .Z( u0_N471 ) , .A( u0_out14_24 ) );
  XOR2_X1 u0_U69 (.B( u0_L13_23 ) , .Z( u0_N470 ) , .A( u0_out14_23 ) );
  XOR2_X1 u0_U75 (.B( u0_L13_18 ) , .Z( u0_N465 ) , .A( u0_out14_18 ) );
  XOR2_X1 u0_U76 (.B( u0_L13_17 ) , .Z( u0_N464 ) , .A( u0_out14_17 ) );
  XOR2_X1 u0_U77 (.B( u0_L13_16 ) , .Z( u0_N463 ) , .A( u0_out14_16 ) );
  XOR2_X1 u0_U80 (.B( u0_L13_13 ) , .Z( u0_N460 ) , .A( u0_out14_13 ) );
  XOR2_X1 u0_U85 (.B( u0_L13_9 ) , .Z( u0_N456 ) , .A( u0_out14_9 ) );
  XOR2_X1 u0_U88 (.B( u0_L13_6 ) , .Z( u0_N453 ) , .A( u0_out14_6 ) );
  XOR2_X1 u0_U93 (.B( u0_L13_2 ) , .Z( u0_N449 ) , .A( u0_out14_2 ) );
  XOR2_X1 u0_U95 (.B( u0_L12_32 ) , .Z( u0_N447 ) , .A( u0_out13_32 ) );
  XOR2_X1 u0_U96 (.B( u0_L12_31 ) , .Z( u0_N446 ) , .A( u0_out13_31 ) );
  XOR2_X1 u0_u13_U10 (.B( u0_K14_45 ) , .A( u0_R12_30 ) , .Z( u0_u13_X_45 ) );
  XOR2_X1 u0_u13_U11 (.B( u0_K14_44 ) , .A( u0_R12_29 ) , .Z( u0_u13_X_44 ) );
  XOR2_X1 u0_u13_U12 (.B( u0_K14_43 ) , .A( u0_R12_28 ) , .Z( u0_u13_X_43 ) );
  XOR2_X1 u0_u13_U13 (.B( u0_K14_42 ) , .A( u0_R12_29 ) , .Z( u0_u13_X_42 ) );
  XOR2_X1 u0_u13_U14 (.B( u0_K14_41 ) , .A( u0_R12_28 ) , .Z( u0_u13_X_41 ) );
  XOR2_X1 u0_u13_U15 (.B( u0_K14_40 ) , .A( u0_R12_27 ) , .Z( u0_u13_X_40 ) );
  XOR2_X1 u0_u13_U16 (.B( u0_K14_3 ) , .A( u0_R12_2 ) , .Z( u0_u13_X_3 ) );
  XOR2_X1 u0_u13_U17 (.B( u0_K14_39 ) , .A( u0_R12_26 ) , .Z( u0_u13_X_39 ) );
  XOR2_X1 u0_u13_U18 (.B( u0_K14_38 ) , .A( u0_R12_25 ) , .Z( u0_u13_X_38 ) );
  XOR2_X1 u0_u13_U19 (.B( u0_K14_37 ) , .A( u0_R12_24 ) , .Z( u0_u13_X_37 ) );
  XOR2_X1 u0_u13_U27 (.B( u0_K14_2 ) , .A( u0_R12_1 ) , .Z( u0_u13_X_2 ) );
  XOR2_X1 u0_u13_U38 (.B( u0_K14_1 ) , .A( u0_R12_32 ) , .Z( u0_u13_X_1 ) );
  XOR2_X1 u0_u13_U4 (.B( u0_K14_6 ) , .A( u0_R12_5 ) , .Z( u0_u13_X_6 ) );
  XOR2_X1 u0_u13_U5 (.B( u0_K14_5 ) , .A( u0_R12_4 ) , .Z( u0_u13_X_5 ) );
  XOR2_X1 u0_u13_U6 (.B( u0_K14_4 ) , .A( u0_R12_3 ) , .Z( u0_u13_X_4 ) );
  XOR2_X1 u0_u13_U7 (.B( u0_K14_48 ) , .A( u0_R12_1 ) , .Z( u0_u13_X_48 ) );
  XOR2_X1 u0_u13_U8 (.B( u0_K14_47 ) , .A( u0_R12_32 ) , .Z( u0_u13_X_47 ) );
  XOR2_X1 u0_u13_U9 (.B( u0_K14_46 ) , .A( u0_R12_31 ) , .Z( u0_u13_X_46 ) );
  AND3_X1 u0_u13_u0_U10 (.A2( u0_u13_u0_n112 ) , .ZN( u0_u13_u0_n127 ) , .A3( u0_u13_u0_n130 ) , .A1( u0_u13_u0_n148 ) );
  NAND2_X1 u0_u13_u0_U11 (.ZN( u0_u13_u0_n113 ) , .A1( u0_u13_u0_n139 ) , .A2( u0_u13_u0_n149 ) );
  AND2_X1 u0_u13_u0_U12 (.ZN( u0_u13_u0_n107 ) , .A1( u0_u13_u0_n130 ) , .A2( u0_u13_u0_n140 ) );
  AND2_X1 u0_u13_u0_U13 (.A2( u0_u13_u0_n129 ) , .A1( u0_u13_u0_n130 ) , .ZN( u0_u13_u0_n151 ) );
  AND2_X1 u0_u13_u0_U14 (.A1( u0_u13_u0_n108 ) , .A2( u0_u13_u0_n125 ) , .ZN( u0_u13_u0_n145 ) );
  INV_X1 u0_u13_u0_U15 (.A( u0_u13_u0_n143 ) , .ZN( u0_u13_u0_n173 ) );
  NOR2_X1 u0_u13_u0_U16 (.A2( u0_u13_u0_n136 ) , .ZN( u0_u13_u0_n147 ) , .A1( u0_u13_u0_n160 ) );
  INV_X1 u0_u13_u0_U17 (.ZN( u0_u13_u0_n172 ) , .A( u0_u13_u0_n88 ) );
  OAI222_X1 u0_u13_u0_U18 (.C1( u0_u13_u0_n108 ) , .A1( u0_u13_u0_n125 ) , .B2( u0_u13_u0_n128 ) , .B1( u0_u13_u0_n144 ) , .A2( u0_u13_u0_n158 ) , .C2( u0_u13_u0_n161 ) , .ZN( u0_u13_u0_n88 ) );
  NOR2_X1 u0_u13_u0_U19 (.A1( u0_u13_u0_n163 ) , .A2( u0_u13_u0_n164 ) , .ZN( u0_u13_u0_n95 ) );
  AOI21_X1 u0_u13_u0_U20 (.B1( u0_u13_u0_n103 ) , .ZN( u0_u13_u0_n132 ) , .A( u0_u13_u0_n165 ) , .B2( u0_u13_u0_n93 ) );
  INV_X1 u0_u13_u0_U21 (.A( u0_u13_u0_n142 ) , .ZN( u0_u13_u0_n165 ) );
  OAI221_X1 u0_u13_u0_U22 (.C1( u0_u13_u0_n121 ) , .ZN( u0_u13_u0_n122 ) , .B2( u0_u13_u0_n127 ) , .A( u0_u13_u0_n143 ) , .B1( u0_u13_u0_n144 ) , .C2( u0_u13_u0_n147 ) );
  OAI22_X1 u0_u13_u0_U23 (.B1( u0_u13_u0_n125 ) , .ZN( u0_u13_u0_n126 ) , .A1( u0_u13_u0_n138 ) , .A2( u0_u13_u0_n146 ) , .B2( u0_u13_u0_n147 ) );
  OAI22_X1 u0_u13_u0_U24 (.B1( u0_u13_u0_n131 ) , .A1( u0_u13_u0_n144 ) , .B2( u0_u13_u0_n147 ) , .A2( u0_u13_u0_n90 ) , .ZN( u0_u13_u0_n91 ) );
  AND3_X1 u0_u13_u0_U25 (.A3( u0_u13_u0_n121 ) , .A2( u0_u13_u0_n125 ) , .A1( u0_u13_u0_n148 ) , .ZN( u0_u13_u0_n90 ) );
  INV_X1 u0_u13_u0_U26 (.A( u0_u13_u0_n136 ) , .ZN( u0_u13_u0_n161 ) );
  NOR2_X1 u0_u13_u0_U27 (.A1( u0_u13_u0_n120 ) , .ZN( u0_u13_u0_n143 ) , .A2( u0_u13_u0_n167 ) );
  OAI221_X1 u0_u13_u0_U28 (.C1( u0_u13_u0_n112 ) , .ZN( u0_u13_u0_n120 ) , .B1( u0_u13_u0_n138 ) , .B2( u0_u13_u0_n141 ) , .C2( u0_u13_u0_n147 ) , .A( u0_u13_u0_n172 ) );
  AOI211_X1 u0_u13_u0_U29 (.B( u0_u13_u0_n115 ) , .A( u0_u13_u0_n116 ) , .C2( u0_u13_u0_n117 ) , .C1( u0_u13_u0_n118 ) , .ZN( u0_u13_u0_n119 ) );
  INV_X1 u0_u13_u0_U3 (.A( u0_u13_u0_n113 ) , .ZN( u0_u13_u0_n166 ) );
  AOI22_X1 u0_u13_u0_U30 (.B2( u0_u13_u0_n109 ) , .A2( u0_u13_u0_n110 ) , .ZN( u0_u13_u0_n111 ) , .B1( u0_u13_u0_n118 ) , .A1( u0_u13_u0_n160 ) );
  INV_X1 u0_u13_u0_U31 (.A( u0_u13_u0_n118 ) , .ZN( u0_u13_u0_n158 ) );
  AOI21_X1 u0_u13_u0_U32 (.ZN( u0_u13_u0_n104 ) , .B1( u0_u13_u0_n107 ) , .B2( u0_u13_u0_n141 ) , .A( u0_u13_u0_n144 ) );
  AOI21_X1 u0_u13_u0_U33 (.B1( u0_u13_u0_n127 ) , .B2( u0_u13_u0_n129 ) , .A( u0_u13_u0_n138 ) , .ZN( u0_u13_u0_n96 ) );
  AOI21_X1 u0_u13_u0_U34 (.ZN( u0_u13_u0_n116 ) , .B2( u0_u13_u0_n142 ) , .A( u0_u13_u0_n144 ) , .B1( u0_u13_u0_n166 ) );
  NAND2_X1 u0_u13_u0_U35 (.A1( u0_u13_u0_n100 ) , .A2( u0_u13_u0_n103 ) , .ZN( u0_u13_u0_n125 ) );
  NAND2_X1 u0_u13_u0_U36 (.A1( u0_u13_u0_n101 ) , .A2( u0_u13_u0_n102 ) , .ZN( u0_u13_u0_n150 ) );
  INV_X1 u0_u13_u0_U37 (.A( u0_u13_u0_n138 ) , .ZN( u0_u13_u0_n160 ) );
  NAND2_X1 u0_u13_u0_U38 (.A1( u0_u13_u0_n102 ) , .ZN( u0_u13_u0_n128 ) , .A2( u0_u13_u0_n95 ) );
  NAND2_X1 u0_u13_u0_U39 (.A1( u0_u13_u0_n100 ) , .ZN( u0_u13_u0_n129 ) , .A2( u0_u13_u0_n95 ) );
  AOI21_X1 u0_u13_u0_U4 (.B1( u0_u13_u0_n114 ) , .ZN( u0_u13_u0_n115 ) , .B2( u0_u13_u0_n129 ) , .A( u0_u13_u0_n161 ) );
  NAND2_X1 u0_u13_u0_U40 (.A2( u0_u13_u0_n100 ) , .ZN( u0_u13_u0_n131 ) , .A1( u0_u13_u0_n92 ) );
  NAND2_X1 u0_u13_u0_U41 (.A2( u0_u13_u0_n100 ) , .A1( u0_u13_u0_n101 ) , .ZN( u0_u13_u0_n139 ) );
  NAND2_X1 u0_u13_u0_U42 (.ZN( u0_u13_u0_n148 ) , .A1( u0_u13_u0_n93 ) , .A2( u0_u13_u0_n95 ) );
  NAND2_X1 u0_u13_u0_U43 (.A2( u0_u13_u0_n102 ) , .A1( u0_u13_u0_n103 ) , .ZN( u0_u13_u0_n149 ) );
  NAND2_X1 u0_u13_u0_U44 (.A2( u0_u13_u0_n102 ) , .ZN( u0_u13_u0_n114 ) , .A1( u0_u13_u0_n92 ) );
  NAND2_X1 u0_u13_u0_U45 (.A2( u0_u13_u0_n101 ) , .ZN( u0_u13_u0_n121 ) , .A1( u0_u13_u0_n93 ) );
  NAND2_X1 u0_u13_u0_U46 (.ZN( u0_u13_u0_n112 ) , .A2( u0_u13_u0_n92 ) , .A1( u0_u13_u0_n93 ) );
  OR3_X1 u0_u13_u0_U47 (.A3( u0_u13_u0_n152 ) , .A2( u0_u13_u0_n153 ) , .A1( u0_u13_u0_n154 ) , .ZN( u0_u13_u0_n155 ) );
  AOI21_X1 u0_u13_u0_U48 (.B2( u0_u13_u0_n150 ) , .B1( u0_u13_u0_n151 ) , .ZN( u0_u13_u0_n152 ) , .A( u0_u13_u0_n158 ) );
  AOI21_X1 u0_u13_u0_U49 (.A( u0_u13_u0_n144 ) , .B2( u0_u13_u0_n145 ) , .B1( u0_u13_u0_n146 ) , .ZN( u0_u13_u0_n154 ) );
  AOI21_X1 u0_u13_u0_U5 (.B2( u0_u13_u0_n131 ) , .ZN( u0_u13_u0_n134 ) , .B1( u0_u13_u0_n151 ) , .A( u0_u13_u0_n158 ) );
  AOI21_X1 u0_u13_u0_U50 (.A( u0_u13_u0_n147 ) , .B2( u0_u13_u0_n148 ) , .B1( u0_u13_u0_n149 ) , .ZN( u0_u13_u0_n153 ) );
  INV_X1 u0_u13_u0_U51 (.ZN( u0_u13_u0_n171 ) , .A( u0_u13_u0_n99 ) );
  OAI211_X1 u0_u13_u0_U52 (.C2( u0_u13_u0_n140 ) , .C1( u0_u13_u0_n161 ) , .A( u0_u13_u0_n169 ) , .B( u0_u13_u0_n98 ) , .ZN( u0_u13_u0_n99 ) );
  AOI211_X1 u0_u13_u0_U53 (.C1( u0_u13_u0_n118 ) , .A( u0_u13_u0_n123 ) , .B( u0_u13_u0_n96 ) , .C2( u0_u13_u0_n97 ) , .ZN( u0_u13_u0_n98 ) );
  INV_X1 u0_u13_u0_U54 (.ZN( u0_u13_u0_n169 ) , .A( u0_u13_u0_n91 ) );
  NOR2_X1 u0_u13_u0_U55 (.A2( u0_u13_X_6 ) , .ZN( u0_u13_u0_n100 ) , .A1( u0_u13_u0_n162 ) );
  NOR2_X1 u0_u13_u0_U56 (.A2( u0_u13_X_4 ) , .A1( u0_u13_X_5 ) , .ZN( u0_u13_u0_n118 ) );
  NOR2_X1 u0_u13_u0_U57 (.A2( u0_u13_X_2 ) , .ZN( u0_u13_u0_n103 ) , .A1( u0_u13_u0_n164 ) );
  NOR2_X1 u0_u13_u0_U58 (.A2( u0_u13_X_1 ) , .A1( u0_u13_X_2 ) , .ZN( u0_u13_u0_n92 ) );
  NOR2_X1 u0_u13_u0_U59 (.A2( u0_u13_X_1 ) , .ZN( u0_u13_u0_n101 ) , .A1( u0_u13_u0_n163 ) );
  NOR2_X1 u0_u13_u0_U6 (.A1( u0_u13_u0_n108 ) , .ZN( u0_u13_u0_n123 ) , .A2( u0_u13_u0_n158 ) );
  NAND2_X1 u0_u13_u0_U60 (.A2( u0_u13_X_4 ) , .A1( u0_u13_X_5 ) , .ZN( u0_u13_u0_n144 ) );
  NOR2_X1 u0_u13_u0_U61 (.A2( u0_u13_X_5 ) , .ZN( u0_u13_u0_n136 ) , .A1( u0_u13_u0_n159 ) );
  NAND2_X1 u0_u13_u0_U62 (.A1( u0_u13_X_5 ) , .ZN( u0_u13_u0_n138 ) , .A2( u0_u13_u0_n159 ) );
  AND2_X1 u0_u13_u0_U63 (.A2( u0_u13_X_3 ) , .A1( u0_u13_X_6 ) , .ZN( u0_u13_u0_n102 ) );
  AND2_X1 u0_u13_u0_U64 (.A1( u0_u13_X_6 ) , .A2( u0_u13_u0_n162 ) , .ZN( u0_u13_u0_n93 ) );
  INV_X1 u0_u13_u0_U65 (.A( u0_u13_X_4 ) , .ZN( u0_u13_u0_n159 ) );
  INV_X1 u0_u13_u0_U66 (.A( u0_u13_X_1 ) , .ZN( u0_u13_u0_n164 ) );
  INV_X1 u0_u13_u0_U67 (.A( u0_u13_X_2 ) , .ZN( u0_u13_u0_n163 ) );
  INV_X1 u0_u13_u0_U68 (.A( u0_u13_u0_n126 ) , .ZN( u0_u13_u0_n168 ) );
  AOI211_X1 u0_u13_u0_U69 (.B( u0_u13_u0_n133 ) , .A( u0_u13_u0_n134 ) , .C2( u0_u13_u0_n135 ) , .C1( u0_u13_u0_n136 ) , .ZN( u0_u13_u0_n137 ) );
  OAI21_X1 u0_u13_u0_U7 (.B1( u0_u13_u0_n150 ) , .B2( u0_u13_u0_n158 ) , .A( u0_u13_u0_n172 ) , .ZN( u0_u13_u0_n89 ) );
  INV_X1 u0_u13_u0_U70 (.ZN( u0_u13_u0_n174 ) , .A( u0_u13_u0_n89 ) );
  AOI211_X1 u0_u13_u0_U71 (.B( u0_u13_u0_n104 ) , .A( u0_u13_u0_n105 ) , .ZN( u0_u13_u0_n106 ) , .C2( u0_u13_u0_n113 ) , .C1( u0_u13_u0_n160 ) );
  OR4_X1 u0_u13_u0_U72 (.ZN( u0_out13_17 ) , .A4( u0_u13_u0_n122 ) , .A2( u0_u13_u0_n123 ) , .A1( u0_u13_u0_n124 ) , .A3( u0_u13_u0_n170 ) );
  AOI21_X1 u0_u13_u0_U73 (.B2( u0_u13_u0_n107 ) , .ZN( u0_u13_u0_n124 ) , .B1( u0_u13_u0_n128 ) , .A( u0_u13_u0_n161 ) );
  INV_X1 u0_u13_u0_U74 (.A( u0_u13_u0_n111 ) , .ZN( u0_u13_u0_n170 ) );
  OR4_X1 u0_u13_u0_U75 (.ZN( u0_out13_31 ) , .A4( u0_u13_u0_n155 ) , .A2( u0_u13_u0_n156 ) , .A1( u0_u13_u0_n157 ) , .A3( u0_u13_u0_n173 ) );
  AOI21_X1 u0_u13_u0_U76 (.A( u0_u13_u0_n138 ) , .B2( u0_u13_u0_n139 ) , .B1( u0_u13_u0_n140 ) , .ZN( u0_u13_u0_n157 ) );
  AOI21_X1 u0_u13_u0_U77 (.B2( u0_u13_u0_n141 ) , .B1( u0_u13_u0_n142 ) , .ZN( u0_u13_u0_n156 ) , .A( u0_u13_u0_n161 ) );
  AOI21_X1 u0_u13_u0_U78 (.B1( u0_u13_u0_n132 ) , .ZN( u0_u13_u0_n133 ) , .A( u0_u13_u0_n144 ) , .B2( u0_u13_u0_n166 ) );
  OAI22_X1 u0_u13_u0_U79 (.ZN( u0_u13_u0_n105 ) , .A2( u0_u13_u0_n132 ) , .B1( u0_u13_u0_n146 ) , .A1( u0_u13_u0_n147 ) , .B2( u0_u13_u0_n161 ) );
  AND2_X1 u0_u13_u0_U8 (.A1( u0_u13_u0_n114 ) , .A2( u0_u13_u0_n121 ) , .ZN( u0_u13_u0_n146 ) );
  NAND2_X1 u0_u13_u0_U80 (.ZN( u0_u13_u0_n110 ) , .A2( u0_u13_u0_n132 ) , .A1( u0_u13_u0_n145 ) );
  INV_X1 u0_u13_u0_U81 (.A( u0_u13_u0_n119 ) , .ZN( u0_u13_u0_n167 ) );
  NAND2_X1 u0_u13_u0_U82 (.A2( u0_u13_u0_n103 ) , .ZN( u0_u13_u0_n140 ) , .A1( u0_u13_u0_n94 ) );
  NAND2_X1 u0_u13_u0_U83 (.A1( u0_u13_u0_n101 ) , .ZN( u0_u13_u0_n130 ) , .A2( u0_u13_u0_n94 ) );
  NAND2_X1 u0_u13_u0_U84 (.ZN( u0_u13_u0_n108 ) , .A1( u0_u13_u0_n92 ) , .A2( u0_u13_u0_n94 ) );
  NAND2_X1 u0_u13_u0_U85 (.ZN( u0_u13_u0_n142 ) , .A1( u0_u13_u0_n94 ) , .A2( u0_u13_u0_n95 ) );
  INV_X1 u0_u13_u0_U86 (.A( u0_u13_X_3 ) , .ZN( u0_u13_u0_n162 ) );
  NOR2_X1 u0_u13_u0_U87 (.A2( u0_u13_X_3 ) , .A1( u0_u13_X_6 ) , .ZN( u0_u13_u0_n94 ) );
  NAND3_X1 u0_u13_u0_U88 (.ZN( u0_out13_23 ) , .A3( u0_u13_u0_n137 ) , .A1( u0_u13_u0_n168 ) , .A2( u0_u13_u0_n171 ) );
  NAND3_X1 u0_u13_u0_U89 (.A3( u0_u13_u0_n127 ) , .A2( u0_u13_u0_n128 ) , .ZN( u0_u13_u0_n135 ) , .A1( u0_u13_u0_n150 ) );
  AND2_X1 u0_u13_u0_U9 (.A1( u0_u13_u0_n131 ) , .ZN( u0_u13_u0_n141 ) , .A2( u0_u13_u0_n150 ) );
  NAND3_X1 u0_u13_u0_U90 (.ZN( u0_u13_u0_n117 ) , .A3( u0_u13_u0_n132 ) , .A2( u0_u13_u0_n139 ) , .A1( u0_u13_u0_n148 ) );
  NAND3_X1 u0_u13_u0_U91 (.ZN( u0_u13_u0_n109 ) , .A2( u0_u13_u0_n114 ) , .A3( u0_u13_u0_n140 ) , .A1( u0_u13_u0_n149 ) );
  NAND3_X1 u0_u13_u0_U92 (.ZN( u0_out13_9 ) , .A3( u0_u13_u0_n106 ) , .A2( u0_u13_u0_n171 ) , .A1( u0_u13_u0_n174 ) );
  NAND3_X1 u0_u13_u0_U93 (.A2( u0_u13_u0_n128 ) , .A1( u0_u13_u0_n132 ) , .A3( u0_u13_u0_n146 ) , .ZN( u0_u13_u0_n97 ) );
  AOI22_X1 u0_u13_u6_U10 (.A2( u0_u13_u6_n151 ) , .B2( u0_u13_u6_n161 ) , .A1( u0_u13_u6_n167 ) , .B1( u0_u13_u6_n170 ) , .ZN( u0_u13_u6_n89 ) );
  AOI21_X1 u0_u13_u6_U11 (.B1( u0_u13_u6_n107 ) , .B2( u0_u13_u6_n132 ) , .A( u0_u13_u6_n158 ) , .ZN( u0_u13_u6_n88 ) );
  AOI21_X1 u0_u13_u6_U12 (.B2( u0_u13_u6_n147 ) , .B1( u0_u13_u6_n148 ) , .ZN( u0_u13_u6_n149 ) , .A( u0_u13_u6_n158 ) );
  AOI21_X1 u0_u13_u6_U13 (.ZN( u0_u13_u6_n106 ) , .A( u0_u13_u6_n142 ) , .B2( u0_u13_u6_n159 ) , .B1( u0_u13_u6_n164 ) );
  INV_X1 u0_u13_u6_U14 (.A( u0_u13_u6_n155 ) , .ZN( u0_u13_u6_n161 ) );
  INV_X1 u0_u13_u6_U15 (.A( u0_u13_u6_n128 ) , .ZN( u0_u13_u6_n164 ) );
  NAND2_X1 u0_u13_u6_U16 (.ZN( u0_u13_u6_n110 ) , .A1( u0_u13_u6_n122 ) , .A2( u0_u13_u6_n129 ) );
  NAND2_X1 u0_u13_u6_U17 (.ZN( u0_u13_u6_n124 ) , .A2( u0_u13_u6_n146 ) , .A1( u0_u13_u6_n148 ) );
  INV_X1 u0_u13_u6_U18 (.A( u0_u13_u6_n132 ) , .ZN( u0_u13_u6_n171 ) );
  AND2_X1 u0_u13_u6_U19 (.A1( u0_u13_u6_n100 ) , .ZN( u0_u13_u6_n130 ) , .A2( u0_u13_u6_n147 ) );
  INV_X1 u0_u13_u6_U20 (.A( u0_u13_u6_n127 ) , .ZN( u0_u13_u6_n173 ) );
  INV_X1 u0_u13_u6_U21 (.A( u0_u13_u6_n121 ) , .ZN( u0_u13_u6_n167 ) );
  INV_X1 u0_u13_u6_U22 (.A( u0_u13_u6_n100 ) , .ZN( u0_u13_u6_n169 ) );
  INV_X1 u0_u13_u6_U23 (.A( u0_u13_u6_n123 ) , .ZN( u0_u13_u6_n170 ) );
  INV_X1 u0_u13_u6_U24 (.A( u0_u13_u6_n113 ) , .ZN( u0_u13_u6_n168 ) );
  AND2_X1 u0_u13_u6_U25 (.A1( u0_u13_u6_n107 ) , .A2( u0_u13_u6_n119 ) , .ZN( u0_u13_u6_n133 ) );
  AND2_X1 u0_u13_u6_U26 (.A2( u0_u13_u6_n121 ) , .A1( u0_u13_u6_n122 ) , .ZN( u0_u13_u6_n131 ) );
  AND3_X1 u0_u13_u6_U27 (.ZN( u0_u13_u6_n120 ) , .A2( u0_u13_u6_n127 ) , .A1( u0_u13_u6_n132 ) , .A3( u0_u13_u6_n145 ) );
  INV_X1 u0_u13_u6_U28 (.A( u0_u13_u6_n146 ) , .ZN( u0_u13_u6_n163 ) );
  AOI222_X1 u0_u13_u6_U29 (.ZN( u0_u13_u6_n114 ) , .A1( u0_u13_u6_n118 ) , .A2( u0_u13_u6_n126 ) , .B2( u0_u13_u6_n151 ) , .C2( u0_u13_u6_n159 ) , .C1( u0_u13_u6_n168 ) , .B1( u0_u13_u6_n169 ) );
  INV_X1 u0_u13_u6_U3 (.A( u0_u13_u6_n110 ) , .ZN( u0_u13_u6_n166 ) );
  NOR2_X1 u0_u13_u6_U30 (.A1( u0_u13_u6_n162 ) , .A2( u0_u13_u6_n165 ) , .ZN( u0_u13_u6_n98 ) );
  AOI211_X1 u0_u13_u6_U31 (.B( u0_u13_u6_n134 ) , .A( u0_u13_u6_n135 ) , .C1( u0_u13_u6_n136 ) , .ZN( u0_u13_u6_n137 ) , .C2( u0_u13_u6_n151 ) );
  AOI21_X1 u0_u13_u6_U32 (.B2( u0_u13_u6_n132 ) , .B1( u0_u13_u6_n133 ) , .ZN( u0_u13_u6_n134 ) , .A( u0_u13_u6_n158 ) );
  AOI21_X1 u0_u13_u6_U33 (.B1( u0_u13_u6_n131 ) , .ZN( u0_u13_u6_n135 ) , .A( u0_u13_u6_n144 ) , .B2( u0_u13_u6_n146 ) );
  NAND4_X1 u0_u13_u6_U34 (.A4( u0_u13_u6_n127 ) , .A3( u0_u13_u6_n128 ) , .A2( u0_u13_u6_n129 ) , .A1( u0_u13_u6_n130 ) , .ZN( u0_u13_u6_n136 ) );
  NAND2_X1 u0_u13_u6_U35 (.A1( u0_u13_u6_n144 ) , .ZN( u0_u13_u6_n151 ) , .A2( u0_u13_u6_n158 ) );
  NAND2_X1 u0_u13_u6_U36 (.ZN( u0_u13_u6_n132 ) , .A1( u0_u13_u6_n91 ) , .A2( u0_u13_u6_n97 ) );
  AOI22_X1 u0_u13_u6_U37 (.B2( u0_u13_u6_n110 ) , .B1( u0_u13_u6_n111 ) , .A1( u0_u13_u6_n112 ) , .ZN( u0_u13_u6_n115 ) , .A2( u0_u13_u6_n161 ) );
  NAND4_X1 u0_u13_u6_U38 (.A3( u0_u13_u6_n109 ) , .ZN( u0_u13_u6_n112 ) , .A4( u0_u13_u6_n132 ) , .A2( u0_u13_u6_n147 ) , .A1( u0_u13_u6_n166 ) );
  NOR2_X1 u0_u13_u6_U39 (.ZN( u0_u13_u6_n109 ) , .A1( u0_u13_u6_n170 ) , .A2( u0_u13_u6_n173 ) );
  INV_X1 u0_u13_u6_U4 (.A( u0_u13_u6_n142 ) , .ZN( u0_u13_u6_n174 ) );
  NOR2_X1 u0_u13_u6_U40 (.A2( u0_u13_u6_n126 ) , .ZN( u0_u13_u6_n155 ) , .A1( u0_u13_u6_n160 ) );
  NAND2_X1 u0_u13_u6_U41 (.ZN( u0_u13_u6_n146 ) , .A2( u0_u13_u6_n94 ) , .A1( u0_u13_u6_n99 ) );
  AOI21_X1 u0_u13_u6_U42 (.A( u0_u13_u6_n144 ) , .B2( u0_u13_u6_n145 ) , .B1( u0_u13_u6_n146 ) , .ZN( u0_u13_u6_n150 ) );
  INV_X1 u0_u13_u6_U43 (.A( u0_u13_u6_n111 ) , .ZN( u0_u13_u6_n158 ) );
  NAND2_X1 u0_u13_u6_U44 (.ZN( u0_u13_u6_n127 ) , .A1( u0_u13_u6_n91 ) , .A2( u0_u13_u6_n92 ) );
  NAND2_X1 u0_u13_u6_U45 (.ZN( u0_u13_u6_n129 ) , .A2( u0_u13_u6_n95 ) , .A1( u0_u13_u6_n96 ) );
  INV_X1 u0_u13_u6_U46 (.A( u0_u13_u6_n144 ) , .ZN( u0_u13_u6_n159 ) );
  NAND2_X1 u0_u13_u6_U47 (.ZN( u0_u13_u6_n145 ) , .A2( u0_u13_u6_n97 ) , .A1( u0_u13_u6_n98 ) );
  NAND2_X1 u0_u13_u6_U48 (.ZN( u0_u13_u6_n148 ) , .A2( u0_u13_u6_n92 ) , .A1( u0_u13_u6_n94 ) );
  NAND2_X1 u0_u13_u6_U49 (.ZN( u0_u13_u6_n108 ) , .A2( u0_u13_u6_n139 ) , .A1( u0_u13_u6_n144 ) );
  NAND2_X1 u0_u13_u6_U5 (.A2( u0_u13_u6_n143 ) , .ZN( u0_u13_u6_n152 ) , .A1( u0_u13_u6_n166 ) );
  NAND2_X1 u0_u13_u6_U50 (.ZN( u0_u13_u6_n121 ) , .A2( u0_u13_u6_n95 ) , .A1( u0_u13_u6_n97 ) );
  NAND2_X1 u0_u13_u6_U51 (.ZN( u0_u13_u6_n107 ) , .A2( u0_u13_u6_n92 ) , .A1( u0_u13_u6_n95 ) );
  AND2_X1 u0_u13_u6_U52 (.ZN( u0_u13_u6_n118 ) , .A2( u0_u13_u6_n91 ) , .A1( u0_u13_u6_n99 ) );
  NAND2_X1 u0_u13_u6_U53 (.ZN( u0_u13_u6_n147 ) , .A2( u0_u13_u6_n98 ) , .A1( u0_u13_u6_n99 ) );
  NAND2_X1 u0_u13_u6_U54 (.ZN( u0_u13_u6_n128 ) , .A1( u0_u13_u6_n94 ) , .A2( u0_u13_u6_n96 ) );
  NAND2_X1 u0_u13_u6_U55 (.ZN( u0_u13_u6_n119 ) , .A2( u0_u13_u6_n95 ) , .A1( u0_u13_u6_n99 ) );
  NAND2_X1 u0_u13_u6_U56 (.ZN( u0_u13_u6_n123 ) , .A2( u0_u13_u6_n91 ) , .A1( u0_u13_u6_n96 ) );
  NAND2_X1 u0_u13_u6_U57 (.ZN( u0_u13_u6_n100 ) , .A2( u0_u13_u6_n92 ) , .A1( u0_u13_u6_n98 ) );
  NAND2_X1 u0_u13_u6_U58 (.ZN( u0_u13_u6_n122 ) , .A1( u0_u13_u6_n94 ) , .A2( u0_u13_u6_n97 ) );
  INV_X1 u0_u13_u6_U59 (.A( u0_u13_u6_n139 ) , .ZN( u0_u13_u6_n160 ) );
  AOI22_X1 u0_u13_u6_U6 (.B2( u0_u13_u6_n101 ) , .A1( u0_u13_u6_n102 ) , .ZN( u0_u13_u6_n103 ) , .B1( u0_u13_u6_n160 ) , .A2( u0_u13_u6_n161 ) );
  NAND2_X1 u0_u13_u6_U60 (.ZN( u0_u13_u6_n113 ) , .A1( u0_u13_u6_n96 ) , .A2( u0_u13_u6_n98 ) );
  NOR2_X1 u0_u13_u6_U61 (.A2( u0_u13_X_40 ) , .A1( u0_u13_X_41 ) , .ZN( u0_u13_u6_n126 ) );
  NOR2_X1 u0_u13_u6_U62 (.A2( u0_u13_X_39 ) , .A1( u0_u13_X_42 ) , .ZN( u0_u13_u6_n92 ) );
  NOR2_X1 u0_u13_u6_U63 (.A2( u0_u13_X_39 ) , .A1( u0_u13_u6_n156 ) , .ZN( u0_u13_u6_n97 ) );
  NOR2_X1 u0_u13_u6_U64 (.A2( u0_u13_X_38 ) , .A1( u0_u13_u6_n165 ) , .ZN( u0_u13_u6_n95 ) );
  NOR2_X1 u0_u13_u6_U65 (.A2( u0_u13_X_41 ) , .ZN( u0_u13_u6_n111 ) , .A1( u0_u13_u6_n157 ) );
  NOR2_X1 u0_u13_u6_U66 (.A2( u0_u13_X_37 ) , .A1( u0_u13_u6_n162 ) , .ZN( u0_u13_u6_n94 ) );
  NOR2_X1 u0_u13_u6_U67 (.A2( u0_u13_X_37 ) , .A1( u0_u13_X_38 ) , .ZN( u0_u13_u6_n91 ) );
  NAND2_X1 u0_u13_u6_U68 (.A1( u0_u13_X_41 ) , .ZN( u0_u13_u6_n144 ) , .A2( u0_u13_u6_n157 ) );
  NAND2_X1 u0_u13_u6_U69 (.A2( u0_u13_X_40 ) , .A1( u0_u13_X_41 ) , .ZN( u0_u13_u6_n139 ) );
  NOR2_X1 u0_u13_u6_U7 (.A1( u0_u13_u6_n118 ) , .ZN( u0_u13_u6_n143 ) , .A2( u0_u13_u6_n168 ) );
  AND2_X1 u0_u13_u6_U70 (.A1( u0_u13_X_39 ) , .A2( u0_u13_u6_n156 ) , .ZN( u0_u13_u6_n96 ) );
  AND2_X1 u0_u13_u6_U71 (.A1( u0_u13_X_39 ) , .A2( u0_u13_X_42 ) , .ZN( u0_u13_u6_n99 ) );
  INV_X1 u0_u13_u6_U72 (.A( u0_u13_X_40 ) , .ZN( u0_u13_u6_n157 ) );
  INV_X1 u0_u13_u6_U73 (.A( u0_u13_X_37 ) , .ZN( u0_u13_u6_n165 ) );
  INV_X1 u0_u13_u6_U74 (.A( u0_u13_X_38 ) , .ZN( u0_u13_u6_n162 ) );
  INV_X1 u0_u13_u6_U75 (.A( u0_u13_X_42 ) , .ZN( u0_u13_u6_n156 ) );
  NAND4_X1 u0_u13_u6_U76 (.ZN( u0_out13_32 ) , .A4( u0_u13_u6_n103 ) , .A3( u0_u13_u6_n104 ) , .A2( u0_u13_u6_n105 ) , .A1( u0_u13_u6_n106 ) );
  AOI22_X1 u0_u13_u6_U77 (.ZN( u0_u13_u6_n105 ) , .A2( u0_u13_u6_n108 ) , .A1( u0_u13_u6_n118 ) , .B2( u0_u13_u6_n126 ) , .B1( u0_u13_u6_n171 ) );
  AOI22_X1 u0_u13_u6_U78 (.ZN( u0_u13_u6_n104 ) , .A1( u0_u13_u6_n111 ) , .B1( u0_u13_u6_n124 ) , .B2( u0_u13_u6_n151 ) , .A2( u0_u13_u6_n93 ) );
  NAND4_X1 u0_u13_u6_U79 (.ZN( u0_out13_12 ) , .A4( u0_u13_u6_n114 ) , .A3( u0_u13_u6_n115 ) , .A2( u0_u13_u6_n116 ) , .A1( u0_u13_u6_n117 ) );
  OAI21_X1 u0_u13_u6_U8 (.A( u0_u13_u6_n159 ) , .B1( u0_u13_u6_n169 ) , .B2( u0_u13_u6_n173 ) , .ZN( u0_u13_u6_n90 ) );
  OAI22_X1 u0_u13_u6_U80 (.B2( u0_u13_u6_n111 ) , .ZN( u0_u13_u6_n116 ) , .B1( u0_u13_u6_n126 ) , .A2( u0_u13_u6_n164 ) , .A1( u0_u13_u6_n167 ) );
  OAI21_X1 u0_u13_u6_U81 (.A( u0_u13_u6_n108 ) , .ZN( u0_u13_u6_n117 ) , .B2( u0_u13_u6_n141 ) , .B1( u0_u13_u6_n163 ) );
  OAI211_X1 u0_u13_u6_U82 (.ZN( u0_out13_7 ) , .B( u0_u13_u6_n153 ) , .C2( u0_u13_u6_n154 ) , .C1( u0_u13_u6_n155 ) , .A( u0_u13_u6_n174 ) );
  NOR3_X1 u0_u13_u6_U83 (.A1( u0_u13_u6_n141 ) , .ZN( u0_u13_u6_n154 ) , .A3( u0_u13_u6_n164 ) , .A2( u0_u13_u6_n171 ) );
  AOI211_X1 u0_u13_u6_U84 (.B( u0_u13_u6_n149 ) , .A( u0_u13_u6_n150 ) , .C2( u0_u13_u6_n151 ) , .C1( u0_u13_u6_n152 ) , .ZN( u0_u13_u6_n153 ) );
  OAI211_X1 u0_u13_u6_U85 (.ZN( u0_out13_22 ) , .B( u0_u13_u6_n137 ) , .A( u0_u13_u6_n138 ) , .C2( u0_u13_u6_n139 ) , .C1( u0_u13_u6_n140 ) );
  AOI22_X1 u0_u13_u6_U86 (.B1( u0_u13_u6_n124 ) , .A2( u0_u13_u6_n125 ) , .A1( u0_u13_u6_n126 ) , .ZN( u0_u13_u6_n138 ) , .B2( u0_u13_u6_n161 ) );
  AND4_X1 u0_u13_u6_U87 (.A3( u0_u13_u6_n119 ) , .A1( u0_u13_u6_n120 ) , .A4( u0_u13_u6_n129 ) , .ZN( u0_u13_u6_n140 ) , .A2( u0_u13_u6_n143 ) );
  NAND3_X1 u0_u13_u6_U88 (.A2( u0_u13_u6_n123 ) , .ZN( u0_u13_u6_n125 ) , .A1( u0_u13_u6_n130 ) , .A3( u0_u13_u6_n131 ) );
  NAND3_X1 u0_u13_u6_U89 (.A3( u0_u13_u6_n133 ) , .ZN( u0_u13_u6_n141 ) , .A1( u0_u13_u6_n145 ) , .A2( u0_u13_u6_n148 ) );
  INV_X1 u0_u13_u6_U9 (.ZN( u0_u13_u6_n172 ) , .A( u0_u13_u6_n88 ) );
  NAND3_X1 u0_u13_u6_U90 (.ZN( u0_u13_u6_n101 ) , .A3( u0_u13_u6_n107 ) , .A2( u0_u13_u6_n121 ) , .A1( u0_u13_u6_n127 ) );
  NAND3_X1 u0_u13_u6_U91 (.ZN( u0_u13_u6_n102 ) , .A3( u0_u13_u6_n130 ) , .A2( u0_u13_u6_n145 ) , .A1( u0_u13_u6_n166 ) );
  NAND3_X1 u0_u13_u6_U92 (.A3( u0_u13_u6_n113 ) , .A1( u0_u13_u6_n119 ) , .A2( u0_u13_u6_n123 ) , .ZN( u0_u13_u6_n93 ) );
  NAND3_X1 u0_u13_u6_U93 (.ZN( u0_u13_u6_n142 ) , .A2( u0_u13_u6_n172 ) , .A3( u0_u13_u6_n89 ) , .A1( u0_u13_u6_n90 ) );
  AND3_X1 u0_u13_u7_U10 (.A3( u0_u13_u7_n110 ) , .A2( u0_u13_u7_n127 ) , .A1( u0_u13_u7_n132 ) , .ZN( u0_u13_u7_n92 ) );
  OAI21_X1 u0_u13_u7_U11 (.A( u0_u13_u7_n161 ) , .B1( u0_u13_u7_n168 ) , .B2( u0_u13_u7_n173 ) , .ZN( u0_u13_u7_n91 ) );
  AOI211_X1 u0_u13_u7_U12 (.A( u0_u13_u7_n117 ) , .ZN( u0_u13_u7_n118 ) , .C2( u0_u13_u7_n126 ) , .C1( u0_u13_u7_n177 ) , .B( u0_u13_u7_n180 ) );
  OAI22_X1 u0_u13_u7_U13 (.B1( u0_u13_u7_n115 ) , .ZN( u0_u13_u7_n117 ) , .A2( u0_u13_u7_n133 ) , .A1( u0_u13_u7_n137 ) , .B2( u0_u13_u7_n162 ) );
  INV_X1 u0_u13_u7_U14 (.A( u0_u13_u7_n116 ) , .ZN( u0_u13_u7_n180 ) );
  NOR3_X1 u0_u13_u7_U15 (.ZN( u0_u13_u7_n115 ) , .A3( u0_u13_u7_n145 ) , .A2( u0_u13_u7_n168 ) , .A1( u0_u13_u7_n169 ) );
  OAI211_X1 u0_u13_u7_U16 (.B( u0_u13_u7_n122 ) , .A( u0_u13_u7_n123 ) , .C2( u0_u13_u7_n124 ) , .ZN( u0_u13_u7_n154 ) , .C1( u0_u13_u7_n162 ) );
  AOI222_X1 u0_u13_u7_U17 (.ZN( u0_u13_u7_n122 ) , .C2( u0_u13_u7_n126 ) , .C1( u0_u13_u7_n145 ) , .B1( u0_u13_u7_n161 ) , .A2( u0_u13_u7_n165 ) , .B2( u0_u13_u7_n170 ) , .A1( u0_u13_u7_n176 ) );
  INV_X1 u0_u13_u7_U18 (.A( u0_u13_u7_n133 ) , .ZN( u0_u13_u7_n176 ) );
  NOR3_X1 u0_u13_u7_U19 (.A2( u0_u13_u7_n134 ) , .A1( u0_u13_u7_n135 ) , .ZN( u0_u13_u7_n136 ) , .A3( u0_u13_u7_n171 ) );
  NOR2_X1 u0_u13_u7_U20 (.A1( u0_u13_u7_n130 ) , .A2( u0_u13_u7_n134 ) , .ZN( u0_u13_u7_n153 ) );
  INV_X1 u0_u13_u7_U21 (.A( u0_u13_u7_n101 ) , .ZN( u0_u13_u7_n165 ) );
  NOR2_X1 u0_u13_u7_U22 (.ZN( u0_u13_u7_n111 ) , .A2( u0_u13_u7_n134 ) , .A1( u0_u13_u7_n169 ) );
  AOI21_X1 u0_u13_u7_U23 (.ZN( u0_u13_u7_n104 ) , .B2( u0_u13_u7_n112 ) , .B1( u0_u13_u7_n127 ) , .A( u0_u13_u7_n164 ) );
  AOI21_X1 u0_u13_u7_U24 (.ZN( u0_u13_u7_n106 ) , .B1( u0_u13_u7_n133 ) , .B2( u0_u13_u7_n146 ) , .A( u0_u13_u7_n162 ) );
  AOI21_X1 u0_u13_u7_U25 (.A( u0_u13_u7_n101 ) , .ZN( u0_u13_u7_n107 ) , .B2( u0_u13_u7_n128 ) , .B1( u0_u13_u7_n175 ) );
  INV_X1 u0_u13_u7_U26 (.A( u0_u13_u7_n138 ) , .ZN( u0_u13_u7_n171 ) );
  INV_X1 u0_u13_u7_U27 (.A( u0_u13_u7_n131 ) , .ZN( u0_u13_u7_n177 ) );
  INV_X1 u0_u13_u7_U28 (.A( u0_u13_u7_n110 ) , .ZN( u0_u13_u7_n174 ) );
  NAND2_X1 u0_u13_u7_U29 (.A1( u0_u13_u7_n129 ) , .A2( u0_u13_u7_n132 ) , .ZN( u0_u13_u7_n149 ) );
  OAI21_X1 u0_u13_u7_U3 (.ZN( u0_u13_u7_n159 ) , .A( u0_u13_u7_n165 ) , .B2( u0_u13_u7_n171 ) , .B1( u0_u13_u7_n174 ) );
  NAND2_X1 u0_u13_u7_U30 (.A1( u0_u13_u7_n113 ) , .A2( u0_u13_u7_n124 ) , .ZN( u0_u13_u7_n130 ) );
  INV_X1 u0_u13_u7_U31 (.A( u0_u13_u7_n112 ) , .ZN( u0_u13_u7_n173 ) );
  INV_X1 u0_u13_u7_U32 (.A( u0_u13_u7_n128 ) , .ZN( u0_u13_u7_n168 ) );
  INV_X1 u0_u13_u7_U33 (.A( u0_u13_u7_n148 ) , .ZN( u0_u13_u7_n169 ) );
  INV_X1 u0_u13_u7_U34 (.A( u0_u13_u7_n127 ) , .ZN( u0_u13_u7_n179 ) );
  NOR2_X1 u0_u13_u7_U35 (.ZN( u0_u13_u7_n101 ) , .A2( u0_u13_u7_n150 ) , .A1( u0_u13_u7_n156 ) );
  AOI211_X1 u0_u13_u7_U36 (.B( u0_u13_u7_n154 ) , .A( u0_u13_u7_n155 ) , .C1( u0_u13_u7_n156 ) , .ZN( u0_u13_u7_n157 ) , .C2( u0_u13_u7_n172 ) );
  INV_X1 u0_u13_u7_U37 (.A( u0_u13_u7_n153 ) , .ZN( u0_u13_u7_n172 ) );
  AOI211_X1 u0_u13_u7_U38 (.B( u0_u13_u7_n139 ) , .A( u0_u13_u7_n140 ) , .C2( u0_u13_u7_n141 ) , .ZN( u0_u13_u7_n142 ) , .C1( u0_u13_u7_n156 ) );
  NAND4_X1 u0_u13_u7_U39 (.A3( u0_u13_u7_n127 ) , .A2( u0_u13_u7_n128 ) , .A1( u0_u13_u7_n129 ) , .ZN( u0_u13_u7_n141 ) , .A4( u0_u13_u7_n147 ) );
  INV_X1 u0_u13_u7_U4 (.A( u0_u13_u7_n111 ) , .ZN( u0_u13_u7_n170 ) );
  AOI21_X1 u0_u13_u7_U40 (.A( u0_u13_u7_n137 ) , .B1( u0_u13_u7_n138 ) , .ZN( u0_u13_u7_n139 ) , .B2( u0_u13_u7_n146 ) );
  OAI22_X1 u0_u13_u7_U41 (.B1( u0_u13_u7_n136 ) , .ZN( u0_u13_u7_n140 ) , .A1( u0_u13_u7_n153 ) , .B2( u0_u13_u7_n162 ) , .A2( u0_u13_u7_n164 ) );
  AOI21_X1 u0_u13_u7_U42 (.ZN( u0_u13_u7_n123 ) , .B1( u0_u13_u7_n165 ) , .B2( u0_u13_u7_n177 ) , .A( u0_u13_u7_n97 ) );
  AOI21_X1 u0_u13_u7_U43 (.B2( u0_u13_u7_n113 ) , .B1( u0_u13_u7_n124 ) , .A( u0_u13_u7_n125 ) , .ZN( u0_u13_u7_n97 ) );
  INV_X1 u0_u13_u7_U44 (.A( u0_u13_u7_n125 ) , .ZN( u0_u13_u7_n161 ) );
  INV_X1 u0_u13_u7_U45 (.A( u0_u13_u7_n152 ) , .ZN( u0_u13_u7_n162 ) );
  AOI22_X1 u0_u13_u7_U46 (.A2( u0_u13_u7_n114 ) , .ZN( u0_u13_u7_n119 ) , .B1( u0_u13_u7_n130 ) , .A1( u0_u13_u7_n156 ) , .B2( u0_u13_u7_n165 ) );
  NAND2_X1 u0_u13_u7_U47 (.A2( u0_u13_u7_n112 ) , .ZN( u0_u13_u7_n114 ) , .A1( u0_u13_u7_n175 ) );
  AND2_X1 u0_u13_u7_U48 (.ZN( u0_u13_u7_n145 ) , .A2( u0_u13_u7_n98 ) , .A1( u0_u13_u7_n99 ) );
  NOR2_X1 u0_u13_u7_U49 (.ZN( u0_u13_u7_n137 ) , .A1( u0_u13_u7_n150 ) , .A2( u0_u13_u7_n161 ) );
  INV_X1 u0_u13_u7_U5 (.A( u0_u13_u7_n149 ) , .ZN( u0_u13_u7_n175 ) );
  AOI21_X1 u0_u13_u7_U50 (.ZN( u0_u13_u7_n105 ) , .B2( u0_u13_u7_n110 ) , .A( u0_u13_u7_n125 ) , .B1( u0_u13_u7_n147 ) );
  NAND2_X1 u0_u13_u7_U51 (.ZN( u0_u13_u7_n146 ) , .A1( u0_u13_u7_n95 ) , .A2( u0_u13_u7_n98 ) );
  NAND2_X1 u0_u13_u7_U52 (.A2( u0_u13_u7_n103 ) , .ZN( u0_u13_u7_n147 ) , .A1( u0_u13_u7_n93 ) );
  NAND2_X1 u0_u13_u7_U53 (.A1( u0_u13_u7_n103 ) , .ZN( u0_u13_u7_n127 ) , .A2( u0_u13_u7_n99 ) );
  OR2_X1 u0_u13_u7_U54 (.ZN( u0_u13_u7_n126 ) , .A2( u0_u13_u7_n152 ) , .A1( u0_u13_u7_n156 ) );
  NAND2_X1 u0_u13_u7_U55 (.A2( u0_u13_u7_n102 ) , .A1( u0_u13_u7_n103 ) , .ZN( u0_u13_u7_n133 ) );
  NAND2_X1 u0_u13_u7_U56 (.ZN( u0_u13_u7_n112 ) , .A2( u0_u13_u7_n96 ) , .A1( u0_u13_u7_n99 ) );
  NAND2_X1 u0_u13_u7_U57 (.A2( u0_u13_u7_n102 ) , .ZN( u0_u13_u7_n128 ) , .A1( u0_u13_u7_n98 ) );
  NAND2_X1 u0_u13_u7_U58 (.A1( u0_u13_u7_n100 ) , .ZN( u0_u13_u7_n113 ) , .A2( u0_u13_u7_n93 ) );
  NAND2_X1 u0_u13_u7_U59 (.A2( u0_u13_u7_n102 ) , .ZN( u0_u13_u7_n124 ) , .A1( u0_u13_u7_n96 ) );
  INV_X1 u0_u13_u7_U6 (.A( u0_u13_u7_n154 ) , .ZN( u0_u13_u7_n178 ) );
  NAND2_X1 u0_u13_u7_U60 (.ZN( u0_u13_u7_n110 ) , .A1( u0_u13_u7_n95 ) , .A2( u0_u13_u7_n96 ) );
  INV_X1 u0_u13_u7_U61 (.A( u0_u13_u7_n150 ) , .ZN( u0_u13_u7_n164 ) );
  AND2_X1 u0_u13_u7_U62 (.ZN( u0_u13_u7_n134 ) , .A1( u0_u13_u7_n93 ) , .A2( u0_u13_u7_n98 ) );
  NAND2_X1 u0_u13_u7_U63 (.A1( u0_u13_u7_n100 ) , .A2( u0_u13_u7_n102 ) , .ZN( u0_u13_u7_n129 ) );
  NAND2_X1 u0_u13_u7_U64 (.A2( u0_u13_u7_n103 ) , .ZN( u0_u13_u7_n131 ) , .A1( u0_u13_u7_n95 ) );
  NAND2_X1 u0_u13_u7_U65 (.A1( u0_u13_u7_n100 ) , .ZN( u0_u13_u7_n138 ) , .A2( u0_u13_u7_n99 ) );
  NAND2_X1 u0_u13_u7_U66 (.ZN( u0_u13_u7_n132 ) , .A1( u0_u13_u7_n93 ) , .A2( u0_u13_u7_n96 ) );
  NAND2_X1 u0_u13_u7_U67 (.A1( u0_u13_u7_n100 ) , .ZN( u0_u13_u7_n148 ) , .A2( u0_u13_u7_n95 ) );
  NOR2_X1 u0_u13_u7_U68 (.A2( u0_u13_X_47 ) , .ZN( u0_u13_u7_n150 ) , .A1( u0_u13_u7_n163 ) );
  NOR2_X1 u0_u13_u7_U69 (.A2( u0_u13_X_43 ) , .A1( u0_u13_X_44 ) , .ZN( u0_u13_u7_n103 ) );
  AOI211_X1 u0_u13_u7_U7 (.ZN( u0_u13_u7_n116 ) , .A( u0_u13_u7_n155 ) , .C1( u0_u13_u7_n161 ) , .C2( u0_u13_u7_n171 ) , .B( u0_u13_u7_n94 ) );
  NOR2_X1 u0_u13_u7_U70 (.A2( u0_u13_X_48 ) , .A1( u0_u13_u7_n166 ) , .ZN( u0_u13_u7_n95 ) );
  NOR2_X1 u0_u13_u7_U71 (.A2( u0_u13_X_45 ) , .A1( u0_u13_X_48 ) , .ZN( u0_u13_u7_n99 ) );
  NOR2_X1 u0_u13_u7_U72 (.A2( u0_u13_X_44 ) , .A1( u0_u13_u7_n167 ) , .ZN( u0_u13_u7_n98 ) );
  NOR2_X1 u0_u13_u7_U73 (.A2( u0_u13_X_46 ) , .A1( u0_u13_X_47 ) , .ZN( u0_u13_u7_n152 ) );
  AND2_X1 u0_u13_u7_U74 (.A1( u0_u13_X_47 ) , .ZN( u0_u13_u7_n156 ) , .A2( u0_u13_u7_n163 ) );
  NAND2_X1 u0_u13_u7_U75 (.A2( u0_u13_X_46 ) , .A1( u0_u13_X_47 ) , .ZN( u0_u13_u7_n125 ) );
  AND2_X1 u0_u13_u7_U76 (.A2( u0_u13_X_45 ) , .A1( u0_u13_X_48 ) , .ZN( u0_u13_u7_n102 ) );
  AND2_X1 u0_u13_u7_U77 (.A2( u0_u13_X_43 ) , .A1( u0_u13_X_44 ) , .ZN( u0_u13_u7_n96 ) );
  AND2_X1 u0_u13_u7_U78 (.A1( u0_u13_X_44 ) , .ZN( u0_u13_u7_n100 ) , .A2( u0_u13_u7_n167 ) );
  AND2_X1 u0_u13_u7_U79 (.A1( u0_u13_X_48 ) , .A2( u0_u13_u7_n166 ) , .ZN( u0_u13_u7_n93 ) );
  OAI222_X1 u0_u13_u7_U8 (.C2( u0_u13_u7_n101 ) , .B2( u0_u13_u7_n111 ) , .A1( u0_u13_u7_n113 ) , .C1( u0_u13_u7_n146 ) , .A2( u0_u13_u7_n162 ) , .B1( u0_u13_u7_n164 ) , .ZN( u0_u13_u7_n94 ) );
  INV_X1 u0_u13_u7_U80 (.A( u0_u13_X_46 ) , .ZN( u0_u13_u7_n163 ) );
  INV_X1 u0_u13_u7_U81 (.A( u0_u13_X_43 ) , .ZN( u0_u13_u7_n167 ) );
  INV_X1 u0_u13_u7_U82 (.A( u0_u13_X_45 ) , .ZN( u0_u13_u7_n166 ) );
  NAND4_X1 u0_u13_u7_U83 (.ZN( u0_out13_27 ) , .A4( u0_u13_u7_n118 ) , .A3( u0_u13_u7_n119 ) , .A2( u0_u13_u7_n120 ) , .A1( u0_u13_u7_n121 ) );
  OAI21_X1 u0_u13_u7_U84 (.ZN( u0_u13_u7_n121 ) , .B2( u0_u13_u7_n145 ) , .A( u0_u13_u7_n150 ) , .B1( u0_u13_u7_n174 ) );
  OAI21_X1 u0_u13_u7_U85 (.ZN( u0_u13_u7_n120 ) , .A( u0_u13_u7_n161 ) , .B2( u0_u13_u7_n170 ) , .B1( u0_u13_u7_n179 ) );
  NAND4_X1 u0_u13_u7_U86 (.ZN( u0_out13_21 ) , .A4( u0_u13_u7_n157 ) , .A3( u0_u13_u7_n158 ) , .A2( u0_u13_u7_n159 ) , .A1( u0_u13_u7_n160 ) );
  OAI21_X1 u0_u13_u7_U87 (.B1( u0_u13_u7_n145 ) , .ZN( u0_u13_u7_n160 ) , .A( u0_u13_u7_n161 ) , .B2( u0_u13_u7_n177 ) );
  AOI22_X1 u0_u13_u7_U88 (.B2( u0_u13_u7_n149 ) , .B1( u0_u13_u7_n150 ) , .A2( u0_u13_u7_n151 ) , .A1( u0_u13_u7_n152 ) , .ZN( u0_u13_u7_n158 ) );
  NAND4_X1 u0_u13_u7_U89 (.ZN( u0_out13_15 ) , .A4( u0_u13_u7_n142 ) , .A3( u0_u13_u7_n143 ) , .A2( u0_u13_u7_n144 ) , .A1( u0_u13_u7_n178 ) );
  OAI221_X1 u0_u13_u7_U9 (.C1( u0_u13_u7_n101 ) , .C2( u0_u13_u7_n147 ) , .ZN( u0_u13_u7_n155 ) , .B2( u0_u13_u7_n162 ) , .A( u0_u13_u7_n91 ) , .B1( u0_u13_u7_n92 ) );
  OR2_X1 u0_u13_u7_U90 (.A2( u0_u13_u7_n125 ) , .A1( u0_u13_u7_n129 ) , .ZN( u0_u13_u7_n144 ) );
  AOI22_X1 u0_u13_u7_U91 (.A2( u0_u13_u7_n126 ) , .ZN( u0_u13_u7_n143 ) , .B2( u0_u13_u7_n165 ) , .B1( u0_u13_u7_n173 ) , .A1( u0_u13_u7_n174 ) );
  NAND4_X1 u0_u13_u7_U92 (.ZN( u0_out13_5 ) , .A4( u0_u13_u7_n108 ) , .A3( u0_u13_u7_n109 ) , .A1( u0_u13_u7_n116 ) , .A2( u0_u13_u7_n123 ) );
  AOI22_X1 u0_u13_u7_U93 (.ZN( u0_u13_u7_n109 ) , .A2( u0_u13_u7_n126 ) , .B2( u0_u13_u7_n145 ) , .B1( u0_u13_u7_n156 ) , .A1( u0_u13_u7_n171 ) );
  NOR4_X1 u0_u13_u7_U94 (.A4( u0_u13_u7_n104 ) , .A3( u0_u13_u7_n105 ) , .A2( u0_u13_u7_n106 ) , .A1( u0_u13_u7_n107 ) , .ZN( u0_u13_u7_n108 ) );
  NAND3_X1 u0_u13_u7_U95 (.A3( u0_u13_u7_n146 ) , .A2( u0_u13_u7_n147 ) , .A1( u0_u13_u7_n148 ) , .ZN( u0_u13_u7_n151 ) );
  NAND3_X1 u0_u13_u7_U96 (.A3( u0_u13_u7_n131 ) , .A2( u0_u13_u7_n132 ) , .A1( u0_u13_u7_n133 ) , .ZN( u0_u13_u7_n135 ) );
  XOR2_X1 u0_u14_U1 (.B( u0_K15_9 ) , .A( u0_R13_6 ) , .Z( u0_u14_X_9 ) );
  XOR2_X1 u0_u14_U16 (.B( u0_K15_3 ) , .A( u0_R13_2 ) , .Z( u0_u14_X_3 ) );
  XOR2_X1 u0_u14_U2 (.B( u0_K15_8 ) , .A( u0_R13_5 ) , .Z( u0_u14_X_8 ) );
  XOR2_X1 u0_u14_U27 (.B( u0_K15_2 ) , .A( u0_R13_1 ) , .Z( u0_u14_X_2 ) );
  XOR2_X1 u0_u14_U3 (.B( u0_K15_7 ) , .A( u0_R13_4 ) , .Z( u0_u14_X_7 ) );
  XOR2_X1 u0_u14_U38 (.B( u0_K15_1 ) , .A( u0_R13_32 ) , .Z( u0_u14_X_1 ) );
  XOR2_X1 u0_u14_U4 (.B( u0_K15_6 ) , .A( u0_R13_5 ) , .Z( u0_u14_X_6 ) );
  XOR2_X1 u0_u14_U40 (.B( u0_K15_18 ) , .A( u0_R13_13 ) , .Z( u0_u14_X_18 ) );
  XOR2_X1 u0_u14_U41 (.B( u0_K15_17 ) , .A( u0_R13_12 ) , .Z( u0_u14_X_17 ) );
  XOR2_X1 u0_u14_U42 (.B( u0_K15_16 ) , .A( u0_R13_11 ) , .Z( u0_u14_X_16 ) );
  XOR2_X1 u0_u14_U43 (.B( u0_K15_15 ) , .A( u0_R13_10 ) , .Z( u0_u14_X_15 ) );
  XOR2_X1 u0_u14_U44 (.B( u0_K15_14 ) , .A( u0_R13_9 ) , .Z( u0_u14_X_14 ) );
  XOR2_X1 u0_u14_U45 (.B( u0_K15_13 ) , .A( u0_R13_8 ) , .Z( u0_u14_X_13 ) );
  XOR2_X1 u0_u14_U46 (.B( u0_K15_12 ) , .A( u0_R13_9 ) , .Z( u0_u14_X_12 ) );
  XOR2_X1 u0_u14_U47 (.B( u0_K15_11 ) , .A( u0_R13_8 ) , .Z( u0_u14_X_11 ) );
  XOR2_X1 u0_u14_U48 (.B( u0_K15_10 ) , .A( u0_R13_7 ) , .Z( u0_u14_X_10 ) );
  XOR2_X1 u0_u14_U5 (.B( u0_K15_5 ) , .A( u0_R13_4 ) , .Z( u0_u14_X_5 ) );
  XOR2_X1 u0_u14_U6 (.B( u0_K15_4 ) , .A( u0_R13_3 ) , .Z( u0_u14_X_4 ) );
  AND3_X1 u0_u14_u0_U10 (.A2( u0_u14_u0_n112 ) , .ZN( u0_u14_u0_n127 ) , .A3( u0_u14_u0_n130 ) , .A1( u0_u14_u0_n148 ) );
  NAND2_X1 u0_u14_u0_U11 (.ZN( u0_u14_u0_n113 ) , .A1( u0_u14_u0_n139 ) , .A2( u0_u14_u0_n149 ) );
  AND2_X1 u0_u14_u0_U12 (.ZN( u0_u14_u0_n107 ) , .A1( u0_u14_u0_n130 ) , .A2( u0_u14_u0_n140 ) );
  AND2_X1 u0_u14_u0_U13 (.A2( u0_u14_u0_n129 ) , .A1( u0_u14_u0_n130 ) , .ZN( u0_u14_u0_n151 ) );
  AND2_X1 u0_u14_u0_U14 (.A1( u0_u14_u0_n108 ) , .A2( u0_u14_u0_n125 ) , .ZN( u0_u14_u0_n145 ) );
  INV_X1 u0_u14_u0_U15 (.A( u0_u14_u0_n143 ) , .ZN( u0_u14_u0_n173 ) );
  NOR2_X1 u0_u14_u0_U16 (.A2( u0_u14_u0_n136 ) , .ZN( u0_u14_u0_n147 ) , .A1( u0_u14_u0_n160 ) );
  NOR2_X1 u0_u14_u0_U17 (.A1( u0_u14_u0_n163 ) , .A2( u0_u14_u0_n164 ) , .ZN( u0_u14_u0_n95 ) );
  AOI21_X1 u0_u14_u0_U18 (.B1( u0_u14_u0_n103 ) , .ZN( u0_u14_u0_n132 ) , .A( u0_u14_u0_n165 ) , .B2( u0_u14_u0_n93 ) );
  INV_X1 u0_u14_u0_U19 (.A( u0_u14_u0_n142 ) , .ZN( u0_u14_u0_n165 ) );
  OAI221_X1 u0_u14_u0_U20 (.C1( u0_u14_u0_n121 ) , .ZN( u0_u14_u0_n122 ) , .B2( u0_u14_u0_n127 ) , .A( u0_u14_u0_n143 ) , .B1( u0_u14_u0_n144 ) , .C2( u0_u14_u0_n147 ) );
  OAI22_X1 u0_u14_u0_U21 (.B1( u0_u14_u0_n125 ) , .ZN( u0_u14_u0_n126 ) , .A1( u0_u14_u0_n138 ) , .A2( u0_u14_u0_n146 ) , .B2( u0_u14_u0_n147 ) );
  OAI22_X1 u0_u14_u0_U22 (.B1( u0_u14_u0_n131 ) , .A1( u0_u14_u0_n144 ) , .B2( u0_u14_u0_n147 ) , .A2( u0_u14_u0_n90 ) , .ZN( u0_u14_u0_n91 ) );
  AND3_X1 u0_u14_u0_U23 (.A3( u0_u14_u0_n121 ) , .A2( u0_u14_u0_n125 ) , .A1( u0_u14_u0_n148 ) , .ZN( u0_u14_u0_n90 ) );
  NAND2_X1 u0_u14_u0_U24 (.A1( u0_u14_u0_n100 ) , .A2( u0_u14_u0_n103 ) , .ZN( u0_u14_u0_n125 ) );
  INV_X1 u0_u14_u0_U25 (.A( u0_u14_u0_n136 ) , .ZN( u0_u14_u0_n161 ) );
  NOR2_X1 u0_u14_u0_U26 (.A1( u0_u14_u0_n120 ) , .ZN( u0_u14_u0_n143 ) , .A2( u0_u14_u0_n167 ) );
  OAI221_X1 u0_u14_u0_U27 (.C1( u0_u14_u0_n112 ) , .ZN( u0_u14_u0_n120 ) , .B1( u0_u14_u0_n138 ) , .B2( u0_u14_u0_n141 ) , .C2( u0_u14_u0_n147 ) , .A( u0_u14_u0_n172 ) );
  AOI211_X1 u0_u14_u0_U28 (.B( u0_u14_u0_n115 ) , .A( u0_u14_u0_n116 ) , .C2( u0_u14_u0_n117 ) , .C1( u0_u14_u0_n118 ) , .ZN( u0_u14_u0_n119 ) );
  AOI22_X1 u0_u14_u0_U29 (.B2( u0_u14_u0_n109 ) , .A2( u0_u14_u0_n110 ) , .ZN( u0_u14_u0_n111 ) , .B1( u0_u14_u0_n118 ) , .A1( u0_u14_u0_n160 ) );
  INV_X1 u0_u14_u0_U3 (.A( u0_u14_u0_n113 ) , .ZN( u0_u14_u0_n166 ) );
  NAND2_X1 u0_u14_u0_U30 (.A1( u0_u14_u0_n100 ) , .ZN( u0_u14_u0_n129 ) , .A2( u0_u14_u0_n95 ) );
  INV_X1 u0_u14_u0_U31 (.A( u0_u14_u0_n118 ) , .ZN( u0_u14_u0_n158 ) );
  AOI21_X1 u0_u14_u0_U32 (.ZN( u0_u14_u0_n104 ) , .B1( u0_u14_u0_n107 ) , .B2( u0_u14_u0_n141 ) , .A( u0_u14_u0_n144 ) );
  AOI21_X1 u0_u14_u0_U33 (.B1( u0_u14_u0_n127 ) , .B2( u0_u14_u0_n129 ) , .A( u0_u14_u0_n138 ) , .ZN( u0_u14_u0_n96 ) );
  AOI21_X1 u0_u14_u0_U34 (.ZN( u0_u14_u0_n116 ) , .B2( u0_u14_u0_n142 ) , .A( u0_u14_u0_n144 ) , .B1( u0_u14_u0_n166 ) );
  NAND2_X1 u0_u14_u0_U35 (.A2( u0_u14_u0_n100 ) , .A1( u0_u14_u0_n101 ) , .ZN( u0_u14_u0_n139 ) );
  NAND2_X1 u0_u14_u0_U36 (.A2( u0_u14_u0_n100 ) , .ZN( u0_u14_u0_n131 ) , .A1( u0_u14_u0_n92 ) );
  NAND2_X1 u0_u14_u0_U37 (.A1( u0_u14_u0_n101 ) , .A2( u0_u14_u0_n102 ) , .ZN( u0_u14_u0_n150 ) );
  INV_X1 u0_u14_u0_U38 (.A( u0_u14_u0_n138 ) , .ZN( u0_u14_u0_n160 ) );
  NAND2_X1 u0_u14_u0_U39 (.A1( u0_u14_u0_n102 ) , .ZN( u0_u14_u0_n128 ) , .A2( u0_u14_u0_n95 ) );
  AOI21_X1 u0_u14_u0_U4 (.B1( u0_u14_u0_n114 ) , .ZN( u0_u14_u0_n115 ) , .B2( u0_u14_u0_n129 ) , .A( u0_u14_u0_n161 ) );
  NAND2_X1 u0_u14_u0_U40 (.ZN( u0_u14_u0_n148 ) , .A1( u0_u14_u0_n93 ) , .A2( u0_u14_u0_n95 ) );
  NAND2_X1 u0_u14_u0_U41 (.A2( u0_u14_u0_n102 ) , .A1( u0_u14_u0_n103 ) , .ZN( u0_u14_u0_n149 ) );
  NAND2_X1 u0_u14_u0_U42 (.A2( u0_u14_u0_n102 ) , .ZN( u0_u14_u0_n114 ) , .A1( u0_u14_u0_n92 ) );
  NAND2_X1 u0_u14_u0_U43 (.A2( u0_u14_u0_n101 ) , .ZN( u0_u14_u0_n121 ) , .A1( u0_u14_u0_n93 ) );
  INV_X1 u0_u14_u0_U44 (.ZN( u0_u14_u0_n172 ) , .A( u0_u14_u0_n88 ) );
  OAI222_X1 u0_u14_u0_U45 (.C1( u0_u14_u0_n108 ) , .A1( u0_u14_u0_n125 ) , .B2( u0_u14_u0_n128 ) , .B1( u0_u14_u0_n144 ) , .A2( u0_u14_u0_n158 ) , .C2( u0_u14_u0_n161 ) , .ZN( u0_u14_u0_n88 ) );
  NAND2_X1 u0_u14_u0_U46 (.ZN( u0_u14_u0_n112 ) , .A2( u0_u14_u0_n92 ) , .A1( u0_u14_u0_n93 ) );
  OR3_X1 u0_u14_u0_U47 (.A3( u0_u14_u0_n152 ) , .A2( u0_u14_u0_n153 ) , .A1( u0_u14_u0_n154 ) , .ZN( u0_u14_u0_n155 ) );
  AOI21_X1 u0_u14_u0_U48 (.B2( u0_u14_u0_n150 ) , .B1( u0_u14_u0_n151 ) , .ZN( u0_u14_u0_n152 ) , .A( u0_u14_u0_n158 ) );
  AOI21_X1 u0_u14_u0_U49 (.A( u0_u14_u0_n144 ) , .B2( u0_u14_u0_n145 ) , .B1( u0_u14_u0_n146 ) , .ZN( u0_u14_u0_n154 ) );
  AOI21_X1 u0_u14_u0_U5 (.B2( u0_u14_u0_n131 ) , .ZN( u0_u14_u0_n134 ) , .B1( u0_u14_u0_n151 ) , .A( u0_u14_u0_n158 ) );
  AOI21_X1 u0_u14_u0_U50 (.A( u0_u14_u0_n147 ) , .B2( u0_u14_u0_n148 ) , .B1( u0_u14_u0_n149 ) , .ZN( u0_u14_u0_n153 ) );
  INV_X1 u0_u14_u0_U51 (.ZN( u0_u14_u0_n171 ) , .A( u0_u14_u0_n99 ) );
  OAI211_X1 u0_u14_u0_U52 (.C2( u0_u14_u0_n140 ) , .C1( u0_u14_u0_n161 ) , .A( u0_u14_u0_n169 ) , .B( u0_u14_u0_n98 ) , .ZN( u0_u14_u0_n99 ) );
  AOI211_X1 u0_u14_u0_U53 (.C1( u0_u14_u0_n118 ) , .A( u0_u14_u0_n123 ) , .B( u0_u14_u0_n96 ) , .C2( u0_u14_u0_n97 ) , .ZN( u0_u14_u0_n98 ) );
  INV_X1 u0_u14_u0_U54 (.ZN( u0_u14_u0_n169 ) , .A( u0_u14_u0_n91 ) );
  NOR2_X1 u0_u14_u0_U55 (.A2( u0_u14_X_4 ) , .A1( u0_u14_X_5 ) , .ZN( u0_u14_u0_n118 ) );
  NOR2_X1 u0_u14_u0_U56 (.A2( u0_u14_X_2 ) , .ZN( u0_u14_u0_n103 ) , .A1( u0_u14_u0_n164 ) );
  NOR2_X1 u0_u14_u0_U57 (.A2( u0_u14_X_1 ) , .A1( u0_u14_X_2 ) , .ZN( u0_u14_u0_n92 ) );
  NOR2_X1 u0_u14_u0_U58 (.A2( u0_u14_X_1 ) , .ZN( u0_u14_u0_n101 ) , .A1( u0_u14_u0_n163 ) );
  NAND2_X1 u0_u14_u0_U59 (.A2( u0_u14_X_4 ) , .A1( u0_u14_X_5 ) , .ZN( u0_u14_u0_n144 ) );
  NOR2_X1 u0_u14_u0_U6 (.A1( u0_u14_u0_n108 ) , .ZN( u0_u14_u0_n123 ) , .A2( u0_u14_u0_n158 ) );
  NOR2_X1 u0_u14_u0_U60 (.A2( u0_u14_X_5 ) , .ZN( u0_u14_u0_n136 ) , .A1( u0_u14_u0_n159 ) );
  NAND2_X1 u0_u14_u0_U61 (.A1( u0_u14_X_5 ) , .ZN( u0_u14_u0_n138 ) , .A2( u0_u14_u0_n159 ) );
  AND2_X1 u0_u14_u0_U62 (.A2( u0_u14_X_3 ) , .A1( u0_u14_X_6 ) , .ZN( u0_u14_u0_n102 ) );
  AND2_X1 u0_u14_u0_U63 (.A1( u0_u14_X_6 ) , .A2( u0_u14_u0_n162 ) , .ZN( u0_u14_u0_n93 ) );
  INV_X1 u0_u14_u0_U64 (.A( u0_u14_X_4 ) , .ZN( u0_u14_u0_n159 ) );
  INV_X1 u0_u14_u0_U65 (.A( u0_u14_X_1 ) , .ZN( u0_u14_u0_n164 ) );
  INV_X1 u0_u14_u0_U66 (.A( u0_u14_X_2 ) , .ZN( u0_u14_u0_n163 ) );
  INV_X1 u0_u14_u0_U67 (.A( u0_u14_X_3 ) , .ZN( u0_u14_u0_n162 ) );
  INV_X1 u0_u14_u0_U68 (.A( u0_u14_u0_n126 ) , .ZN( u0_u14_u0_n168 ) );
  AOI211_X1 u0_u14_u0_U69 (.B( u0_u14_u0_n133 ) , .A( u0_u14_u0_n134 ) , .C2( u0_u14_u0_n135 ) , .C1( u0_u14_u0_n136 ) , .ZN( u0_u14_u0_n137 ) );
  OAI21_X1 u0_u14_u0_U7 (.B1( u0_u14_u0_n150 ) , .B2( u0_u14_u0_n158 ) , .A( u0_u14_u0_n172 ) , .ZN( u0_u14_u0_n89 ) );
  INV_X1 u0_u14_u0_U70 (.ZN( u0_u14_u0_n174 ) , .A( u0_u14_u0_n89 ) );
  AOI211_X1 u0_u14_u0_U71 (.B( u0_u14_u0_n104 ) , .A( u0_u14_u0_n105 ) , .ZN( u0_u14_u0_n106 ) , .C2( u0_u14_u0_n113 ) , .C1( u0_u14_u0_n160 ) );
  OR4_X1 u0_u14_u0_U72 (.ZN( u0_out14_31 ) , .A4( u0_u14_u0_n155 ) , .A2( u0_u14_u0_n156 ) , .A1( u0_u14_u0_n157 ) , .A3( u0_u14_u0_n173 ) );
  AOI21_X1 u0_u14_u0_U73 (.A( u0_u14_u0_n138 ) , .B2( u0_u14_u0_n139 ) , .B1( u0_u14_u0_n140 ) , .ZN( u0_u14_u0_n157 ) );
  AOI21_X1 u0_u14_u0_U74 (.B2( u0_u14_u0_n141 ) , .B1( u0_u14_u0_n142 ) , .ZN( u0_u14_u0_n156 ) , .A( u0_u14_u0_n161 ) );
  OR4_X1 u0_u14_u0_U75 (.ZN( u0_out14_17 ) , .A4( u0_u14_u0_n122 ) , .A2( u0_u14_u0_n123 ) , .A1( u0_u14_u0_n124 ) , .A3( u0_u14_u0_n170 ) );
  AOI21_X1 u0_u14_u0_U76 (.B2( u0_u14_u0_n107 ) , .ZN( u0_u14_u0_n124 ) , .B1( u0_u14_u0_n128 ) , .A( u0_u14_u0_n161 ) );
  INV_X1 u0_u14_u0_U77 (.A( u0_u14_u0_n111 ) , .ZN( u0_u14_u0_n170 ) );
  AOI21_X1 u0_u14_u0_U78 (.B1( u0_u14_u0_n132 ) , .ZN( u0_u14_u0_n133 ) , .A( u0_u14_u0_n144 ) , .B2( u0_u14_u0_n166 ) );
  OAI22_X1 u0_u14_u0_U79 (.ZN( u0_u14_u0_n105 ) , .A2( u0_u14_u0_n132 ) , .B1( u0_u14_u0_n146 ) , .A1( u0_u14_u0_n147 ) , .B2( u0_u14_u0_n161 ) );
  AND2_X1 u0_u14_u0_U8 (.A1( u0_u14_u0_n114 ) , .A2( u0_u14_u0_n121 ) , .ZN( u0_u14_u0_n146 ) );
  NAND2_X1 u0_u14_u0_U80 (.ZN( u0_u14_u0_n110 ) , .A2( u0_u14_u0_n132 ) , .A1( u0_u14_u0_n145 ) );
  INV_X1 u0_u14_u0_U81 (.A( u0_u14_u0_n119 ) , .ZN( u0_u14_u0_n167 ) );
  NAND2_X1 u0_u14_u0_U82 (.A2( u0_u14_u0_n103 ) , .ZN( u0_u14_u0_n140 ) , .A1( u0_u14_u0_n94 ) );
  NAND2_X1 u0_u14_u0_U83 (.A1( u0_u14_u0_n101 ) , .ZN( u0_u14_u0_n130 ) , .A2( u0_u14_u0_n94 ) );
  NAND2_X1 u0_u14_u0_U84 (.ZN( u0_u14_u0_n108 ) , .A1( u0_u14_u0_n92 ) , .A2( u0_u14_u0_n94 ) );
  NAND2_X1 u0_u14_u0_U85 (.ZN( u0_u14_u0_n142 ) , .A1( u0_u14_u0_n94 ) , .A2( u0_u14_u0_n95 ) );
  NOR2_X1 u0_u14_u0_U86 (.A2( u0_u14_X_6 ) , .ZN( u0_u14_u0_n100 ) , .A1( u0_u14_u0_n162 ) );
  NOR2_X1 u0_u14_u0_U87 (.A2( u0_u14_X_3 ) , .A1( u0_u14_X_6 ) , .ZN( u0_u14_u0_n94 ) );
  NAND3_X1 u0_u14_u0_U88 (.ZN( u0_out14_23 ) , .A3( u0_u14_u0_n137 ) , .A1( u0_u14_u0_n168 ) , .A2( u0_u14_u0_n171 ) );
  NAND3_X1 u0_u14_u0_U89 (.A3( u0_u14_u0_n127 ) , .A2( u0_u14_u0_n128 ) , .ZN( u0_u14_u0_n135 ) , .A1( u0_u14_u0_n150 ) );
  AND2_X1 u0_u14_u0_U9 (.A1( u0_u14_u0_n131 ) , .ZN( u0_u14_u0_n141 ) , .A2( u0_u14_u0_n150 ) );
  NAND3_X1 u0_u14_u0_U90 (.ZN( u0_u14_u0_n117 ) , .A3( u0_u14_u0_n132 ) , .A2( u0_u14_u0_n139 ) , .A1( u0_u14_u0_n148 ) );
  NAND3_X1 u0_u14_u0_U91 (.ZN( u0_u14_u0_n109 ) , .A2( u0_u14_u0_n114 ) , .A3( u0_u14_u0_n140 ) , .A1( u0_u14_u0_n149 ) );
  NAND3_X1 u0_u14_u0_U92 (.ZN( u0_out14_9 ) , .A3( u0_u14_u0_n106 ) , .A2( u0_u14_u0_n171 ) , .A1( u0_u14_u0_n174 ) );
  NAND3_X1 u0_u14_u0_U93 (.A2( u0_u14_u0_n128 ) , .A1( u0_u14_u0_n132 ) , .A3( u0_u14_u0_n146 ) , .ZN( u0_u14_u0_n97 ) );
  AOI21_X1 u0_u14_u1_U10 (.ZN( u0_u14_u1_n106 ) , .A( u0_u14_u1_n112 ) , .B1( u0_u14_u1_n154 ) , .B2( u0_u14_u1_n156 ) );
  NAND3_X1 u0_u14_u1_U100 (.ZN( u0_u14_u1_n113 ) , .A1( u0_u14_u1_n120 ) , .A3( u0_u14_u1_n133 ) , .A2( u0_u14_u1_n155 ) );
  INV_X1 u0_u14_u1_U11 (.A( u0_u14_u1_n101 ) , .ZN( u0_u14_u1_n184 ) );
  AOI21_X1 u0_u14_u1_U12 (.ZN( u0_u14_u1_n107 ) , .B1( u0_u14_u1_n134 ) , .B2( u0_u14_u1_n149 ) , .A( u0_u14_u1_n174 ) );
  NAND2_X1 u0_u14_u1_U13 (.ZN( u0_u14_u1_n140 ) , .A2( u0_u14_u1_n150 ) , .A1( u0_u14_u1_n155 ) );
  NAND2_X1 u0_u14_u1_U14 (.A1( u0_u14_u1_n131 ) , .ZN( u0_u14_u1_n147 ) , .A2( u0_u14_u1_n153 ) );
  AOI22_X1 u0_u14_u1_U15 (.B2( u0_u14_u1_n136 ) , .A2( u0_u14_u1_n137 ) , .ZN( u0_u14_u1_n143 ) , .A1( u0_u14_u1_n171 ) , .B1( u0_u14_u1_n173 ) );
  INV_X1 u0_u14_u1_U16 (.A( u0_u14_u1_n147 ) , .ZN( u0_u14_u1_n181 ) );
  INV_X1 u0_u14_u1_U17 (.A( u0_u14_u1_n139 ) , .ZN( u0_u14_u1_n174 ) );
  INV_X1 u0_u14_u1_U18 (.A( u0_u14_u1_n112 ) , .ZN( u0_u14_u1_n171 ) );
  NAND2_X1 u0_u14_u1_U19 (.ZN( u0_u14_u1_n141 ) , .A1( u0_u14_u1_n153 ) , .A2( u0_u14_u1_n156 ) );
  AND2_X1 u0_u14_u1_U20 (.A1( u0_u14_u1_n123 ) , .ZN( u0_u14_u1_n134 ) , .A2( u0_u14_u1_n161 ) );
  NAND2_X1 u0_u14_u1_U21 (.A2( u0_u14_u1_n115 ) , .A1( u0_u14_u1_n116 ) , .ZN( u0_u14_u1_n148 ) );
  NAND2_X1 u0_u14_u1_U22 (.A2( u0_u14_u1_n133 ) , .A1( u0_u14_u1_n135 ) , .ZN( u0_u14_u1_n159 ) );
  NAND2_X1 u0_u14_u1_U23 (.A2( u0_u14_u1_n115 ) , .A1( u0_u14_u1_n120 ) , .ZN( u0_u14_u1_n132 ) );
  INV_X1 u0_u14_u1_U24 (.A( u0_u14_u1_n154 ) , .ZN( u0_u14_u1_n178 ) );
  AOI22_X1 u0_u14_u1_U25 (.B2( u0_u14_u1_n113 ) , .A2( u0_u14_u1_n114 ) , .ZN( u0_u14_u1_n125 ) , .A1( u0_u14_u1_n171 ) , .B1( u0_u14_u1_n173 ) );
  NAND2_X1 u0_u14_u1_U26 (.ZN( u0_u14_u1_n114 ) , .A1( u0_u14_u1_n134 ) , .A2( u0_u14_u1_n156 ) );
  INV_X1 u0_u14_u1_U27 (.A( u0_u14_u1_n151 ) , .ZN( u0_u14_u1_n183 ) );
  AND2_X1 u0_u14_u1_U28 (.A1( u0_u14_u1_n129 ) , .A2( u0_u14_u1_n133 ) , .ZN( u0_u14_u1_n149 ) );
  INV_X1 u0_u14_u1_U29 (.A( u0_u14_u1_n131 ) , .ZN( u0_u14_u1_n180 ) );
  INV_X1 u0_u14_u1_U3 (.A( u0_u14_u1_n159 ) , .ZN( u0_u14_u1_n182 ) );
  AOI221_X1 u0_u14_u1_U30 (.B1( u0_u14_u1_n140 ) , .ZN( u0_u14_u1_n167 ) , .B2( u0_u14_u1_n172 ) , .C2( u0_u14_u1_n175 ) , .C1( u0_u14_u1_n178 ) , .A( u0_u14_u1_n188 ) );
  INV_X1 u0_u14_u1_U31 (.ZN( u0_u14_u1_n188 ) , .A( u0_u14_u1_n97 ) );
  AOI211_X1 u0_u14_u1_U32 (.A( u0_u14_u1_n118 ) , .C1( u0_u14_u1_n132 ) , .C2( u0_u14_u1_n139 ) , .B( u0_u14_u1_n96 ) , .ZN( u0_u14_u1_n97 ) );
  AOI21_X1 u0_u14_u1_U33 (.B2( u0_u14_u1_n121 ) , .B1( u0_u14_u1_n135 ) , .A( u0_u14_u1_n152 ) , .ZN( u0_u14_u1_n96 ) );
  OAI221_X1 u0_u14_u1_U34 (.A( u0_u14_u1_n119 ) , .C2( u0_u14_u1_n129 ) , .ZN( u0_u14_u1_n138 ) , .B2( u0_u14_u1_n152 ) , .C1( u0_u14_u1_n174 ) , .B1( u0_u14_u1_n187 ) );
  INV_X1 u0_u14_u1_U35 (.A( u0_u14_u1_n148 ) , .ZN( u0_u14_u1_n187 ) );
  AOI211_X1 u0_u14_u1_U36 (.B( u0_u14_u1_n117 ) , .A( u0_u14_u1_n118 ) , .ZN( u0_u14_u1_n119 ) , .C2( u0_u14_u1_n146 ) , .C1( u0_u14_u1_n159 ) );
  NOR2_X1 u0_u14_u1_U37 (.A1( u0_u14_u1_n168 ) , .A2( u0_u14_u1_n176 ) , .ZN( u0_u14_u1_n98 ) );
  AOI211_X1 u0_u14_u1_U38 (.B( u0_u14_u1_n162 ) , .A( u0_u14_u1_n163 ) , .C2( u0_u14_u1_n164 ) , .ZN( u0_u14_u1_n165 ) , .C1( u0_u14_u1_n171 ) );
  AOI21_X1 u0_u14_u1_U39 (.A( u0_u14_u1_n160 ) , .B2( u0_u14_u1_n161 ) , .ZN( u0_u14_u1_n162 ) , .B1( u0_u14_u1_n182 ) );
  AOI221_X1 u0_u14_u1_U4 (.A( u0_u14_u1_n138 ) , .C2( u0_u14_u1_n139 ) , .C1( u0_u14_u1_n140 ) , .B2( u0_u14_u1_n141 ) , .ZN( u0_u14_u1_n142 ) , .B1( u0_u14_u1_n175 ) );
  OR2_X1 u0_u14_u1_U40 (.A2( u0_u14_u1_n157 ) , .A1( u0_u14_u1_n158 ) , .ZN( u0_u14_u1_n163 ) );
  OAI21_X1 u0_u14_u1_U41 (.B2( u0_u14_u1_n123 ) , .ZN( u0_u14_u1_n145 ) , .B1( u0_u14_u1_n160 ) , .A( u0_u14_u1_n185 ) );
  INV_X1 u0_u14_u1_U42 (.A( u0_u14_u1_n122 ) , .ZN( u0_u14_u1_n185 ) );
  AOI21_X1 u0_u14_u1_U43 (.B2( u0_u14_u1_n120 ) , .B1( u0_u14_u1_n121 ) , .ZN( u0_u14_u1_n122 ) , .A( u0_u14_u1_n128 ) );
  NAND2_X1 u0_u14_u1_U44 (.A1( u0_u14_u1_n128 ) , .ZN( u0_u14_u1_n146 ) , .A2( u0_u14_u1_n160 ) );
  NAND2_X1 u0_u14_u1_U45 (.A2( u0_u14_u1_n112 ) , .ZN( u0_u14_u1_n139 ) , .A1( u0_u14_u1_n152 ) );
  NAND2_X1 u0_u14_u1_U46 (.A1( u0_u14_u1_n105 ) , .ZN( u0_u14_u1_n156 ) , .A2( u0_u14_u1_n99 ) );
  NOR2_X1 u0_u14_u1_U47 (.ZN( u0_u14_u1_n117 ) , .A1( u0_u14_u1_n121 ) , .A2( u0_u14_u1_n160 ) );
  AOI21_X1 u0_u14_u1_U48 (.A( u0_u14_u1_n128 ) , .B2( u0_u14_u1_n129 ) , .ZN( u0_u14_u1_n130 ) , .B1( u0_u14_u1_n150 ) );
  NAND2_X1 u0_u14_u1_U49 (.ZN( u0_u14_u1_n112 ) , .A1( u0_u14_u1_n169 ) , .A2( u0_u14_u1_n170 ) );
  AOI211_X1 u0_u14_u1_U5 (.ZN( u0_u14_u1_n124 ) , .A( u0_u14_u1_n138 ) , .C2( u0_u14_u1_n139 ) , .B( u0_u14_u1_n145 ) , .C1( u0_u14_u1_n147 ) );
  NAND2_X1 u0_u14_u1_U50 (.ZN( u0_u14_u1_n129 ) , .A2( u0_u14_u1_n95 ) , .A1( u0_u14_u1_n98 ) );
  NAND2_X1 u0_u14_u1_U51 (.A1( u0_u14_u1_n102 ) , .ZN( u0_u14_u1_n154 ) , .A2( u0_u14_u1_n99 ) );
  NAND2_X1 u0_u14_u1_U52 (.A2( u0_u14_u1_n100 ) , .ZN( u0_u14_u1_n135 ) , .A1( u0_u14_u1_n99 ) );
  AOI21_X1 u0_u14_u1_U53 (.A( u0_u14_u1_n152 ) , .B2( u0_u14_u1_n153 ) , .B1( u0_u14_u1_n154 ) , .ZN( u0_u14_u1_n158 ) );
  INV_X1 u0_u14_u1_U54 (.A( u0_u14_u1_n160 ) , .ZN( u0_u14_u1_n175 ) );
  NAND2_X1 u0_u14_u1_U55 (.A1( u0_u14_u1_n100 ) , .ZN( u0_u14_u1_n116 ) , .A2( u0_u14_u1_n95 ) );
  NAND2_X1 u0_u14_u1_U56 (.A1( u0_u14_u1_n102 ) , .ZN( u0_u14_u1_n131 ) , .A2( u0_u14_u1_n95 ) );
  NAND2_X1 u0_u14_u1_U57 (.A2( u0_u14_u1_n104 ) , .ZN( u0_u14_u1_n121 ) , .A1( u0_u14_u1_n98 ) );
  NAND2_X1 u0_u14_u1_U58 (.A1( u0_u14_u1_n103 ) , .ZN( u0_u14_u1_n153 ) , .A2( u0_u14_u1_n98 ) );
  NAND2_X1 u0_u14_u1_U59 (.A2( u0_u14_u1_n104 ) , .A1( u0_u14_u1_n105 ) , .ZN( u0_u14_u1_n133 ) );
  NOR2_X1 u0_u14_u1_U6 (.A1( u0_u14_u1_n112 ) , .A2( u0_u14_u1_n116 ) , .ZN( u0_u14_u1_n118 ) );
  NAND2_X1 u0_u14_u1_U60 (.ZN( u0_u14_u1_n150 ) , .A2( u0_u14_u1_n98 ) , .A1( u0_u14_u1_n99 ) );
  NAND2_X1 u0_u14_u1_U61 (.A1( u0_u14_u1_n105 ) , .ZN( u0_u14_u1_n155 ) , .A2( u0_u14_u1_n95 ) );
  OAI21_X1 u0_u14_u1_U62 (.ZN( u0_u14_u1_n109 ) , .B1( u0_u14_u1_n129 ) , .B2( u0_u14_u1_n160 ) , .A( u0_u14_u1_n167 ) );
  NAND2_X1 u0_u14_u1_U63 (.A2( u0_u14_u1_n100 ) , .A1( u0_u14_u1_n103 ) , .ZN( u0_u14_u1_n120 ) );
  NAND2_X1 u0_u14_u1_U64 (.A1( u0_u14_u1_n102 ) , .A2( u0_u14_u1_n104 ) , .ZN( u0_u14_u1_n115 ) );
  NAND2_X1 u0_u14_u1_U65 (.A2( u0_u14_u1_n100 ) , .A1( u0_u14_u1_n104 ) , .ZN( u0_u14_u1_n151 ) );
  NAND2_X1 u0_u14_u1_U66 (.A2( u0_u14_u1_n103 ) , .A1( u0_u14_u1_n105 ) , .ZN( u0_u14_u1_n161 ) );
  INV_X1 u0_u14_u1_U67 (.A( u0_u14_u1_n152 ) , .ZN( u0_u14_u1_n173 ) );
  INV_X1 u0_u14_u1_U68 (.A( u0_u14_u1_n128 ) , .ZN( u0_u14_u1_n172 ) );
  NAND2_X1 u0_u14_u1_U69 (.A2( u0_u14_u1_n102 ) , .A1( u0_u14_u1_n103 ) , .ZN( u0_u14_u1_n123 ) );
  OAI21_X1 u0_u14_u1_U7 (.ZN( u0_u14_u1_n101 ) , .B1( u0_u14_u1_n141 ) , .A( u0_u14_u1_n146 ) , .B2( u0_u14_u1_n183 ) );
  NOR2_X1 u0_u14_u1_U70 (.A2( u0_u14_X_7 ) , .A1( u0_u14_X_8 ) , .ZN( u0_u14_u1_n95 ) );
  NOR2_X1 u0_u14_u1_U71 (.A1( u0_u14_X_12 ) , .A2( u0_u14_X_9 ) , .ZN( u0_u14_u1_n100 ) );
  NOR2_X1 u0_u14_u1_U72 (.A2( u0_u14_X_8 ) , .A1( u0_u14_u1_n177 ) , .ZN( u0_u14_u1_n99 ) );
  NOR2_X1 u0_u14_u1_U73 (.A2( u0_u14_X_12 ) , .ZN( u0_u14_u1_n102 ) , .A1( u0_u14_u1_n176 ) );
  NOR2_X1 u0_u14_u1_U74 (.A2( u0_u14_X_9 ) , .ZN( u0_u14_u1_n105 ) , .A1( u0_u14_u1_n168 ) );
  NAND2_X1 u0_u14_u1_U75 (.A1( u0_u14_X_10 ) , .ZN( u0_u14_u1_n160 ) , .A2( u0_u14_u1_n169 ) );
  NAND2_X1 u0_u14_u1_U76 (.A2( u0_u14_X_10 ) , .A1( u0_u14_X_11 ) , .ZN( u0_u14_u1_n152 ) );
  NAND2_X1 u0_u14_u1_U77 (.A1( u0_u14_X_11 ) , .ZN( u0_u14_u1_n128 ) , .A2( u0_u14_u1_n170 ) );
  AND2_X1 u0_u14_u1_U78 (.A2( u0_u14_X_7 ) , .A1( u0_u14_X_8 ) , .ZN( u0_u14_u1_n104 ) );
  AND2_X1 u0_u14_u1_U79 (.A1( u0_u14_X_8 ) , .ZN( u0_u14_u1_n103 ) , .A2( u0_u14_u1_n177 ) );
  AOI21_X1 u0_u14_u1_U8 (.B2( u0_u14_u1_n155 ) , .B1( u0_u14_u1_n156 ) , .ZN( u0_u14_u1_n157 ) , .A( u0_u14_u1_n174 ) );
  INV_X1 u0_u14_u1_U80 (.A( u0_u14_X_10 ) , .ZN( u0_u14_u1_n170 ) );
  INV_X1 u0_u14_u1_U81 (.A( u0_u14_X_9 ) , .ZN( u0_u14_u1_n176 ) );
  INV_X1 u0_u14_u1_U82 (.A( u0_u14_X_11 ) , .ZN( u0_u14_u1_n169 ) );
  INV_X1 u0_u14_u1_U83 (.A( u0_u14_X_12 ) , .ZN( u0_u14_u1_n168 ) );
  INV_X1 u0_u14_u1_U84 (.A( u0_u14_X_7 ) , .ZN( u0_u14_u1_n177 ) );
  NAND4_X1 u0_u14_u1_U85 (.ZN( u0_out14_28 ) , .A4( u0_u14_u1_n124 ) , .A3( u0_u14_u1_n125 ) , .A2( u0_u14_u1_n126 ) , .A1( u0_u14_u1_n127 ) );
  OAI21_X1 u0_u14_u1_U86 (.ZN( u0_u14_u1_n127 ) , .B2( u0_u14_u1_n139 ) , .B1( u0_u14_u1_n175 ) , .A( u0_u14_u1_n183 ) );
  OAI21_X1 u0_u14_u1_U87 (.ZN( u0_u14_u1_n126 ) , .B2( u0_u14_u1_n140 ) , .A( u0_u14_u1_n146 ) , .B1( u0_u14_u1_n178 ) );
  NAND4_X1 u0_u14_u1_U88 (.ZN( u0_out14_18 ) , .A4( u0_u14_u1_n165 ) , .A3( u0_u14_u1_n166 ) , .A1( u0_u14_u1_n167 ) , .A2( u0_u14_u1_n186 ) );
  AOI22_X1 u0_u14_u1_U89 (.B2( u0_u14_u1_n146 ) , .B1( u0_u14_u1_n147 ) , .A2( u0_u14_u1_n148 ) , .ZN( u0_u14_u1_n166 ) , .A1( u0_u14_u1_n172 ) );
  OR4_X1 u0_u14_u1_U9 (.A4( u0_u14_u1_n106 ) , .A3( u0_u14_u1_n107 ) , .ZN( u0_u14_u1_n108 ) , .A1( u0_u14_u1_n117 ) , .A2( u0_u14_u1_n184 ) );
  INV_X1 u0_u14_u1_U90 (.A( u0_u14_u1_n145 ) , .ZN( u0_u14_u1_n186 ) );
  NAND4_X1 u0_u14_u1_U91 (.ZN( u0_out14_2 ) , .A4( u0_u14_u1_n142 ) , .A3( u0_u14_u1_n143 ) , .A2( u0_u14_u1_n144 ) , .A1( u0_u14_u1_n179 ) );
  OAI21_X1 u0_u14_u1_U92 (.B2( u0_u14_u1_n132 ) , .ZN( u0_u14_u1_n144 ) , .A( u0_u14_u1_n146 ) , .B1( u0_u14_u1_n180 ) );
  INV_X1 u0_u14_u1_U93 (.A( u0_u14_u1_n130 ) , .ZN( u0_u14_u1_n179 ) );
  OR4_X1 u0_u14_u1_U94 (.ZN( u0_out14_13 ) , .A4( u0_u14_u1_n108 ) , .A3( u0_u14_u1_n109 ) , .A2( u0_u14_u1_n110 ) , .A1( u0_u14_u1_n111 ) );
  AOI21_X1 u0_u14_u1_U95 (.ZN( u0_u14_u1_n111 ) , .A( u0_u14_u1_n128 ) , .B2( u0_u14_u1_n131 ) , .B1( u0_u14_u1_n135 ) );
  AOI21_X1 u0_u14_u1_U96 (.ZN( u0_u14_u1_n110 ) , .A( u0_u14_u1_n116 ) , .B1( u0_u14_u1_n152 ) , .B2( u0_u14_u1_n160 ) );
  NAND3_X1 u0_u14_u1_U97 (.A3( u0_u14_u1_n149 ) , .A2( u0_u14_u1_n150 ) , .A1( u0_u14_u1_n151 ) , .ZN( u0_u14_u1_n164 ) );
  NAND3_X1 u0_u14_u1_U98 (.A3( u0_u14_u1_n134 ) , .A2( u0_u14_u1_n135 ) , .ZN( u0_u14_u1_n136 ) , .A1( u0_u14_u1_n151 ) );
  NAND3_X1 u0_u14_u1_U99 (.A1( u0_u14_u1_n133 ) , .ZN( u0_u14_u1_n137 ) , .A2( u0_u14_u1_n154 ) , .A3( u0_u14_u1_n181 ) );
  OAI22_X1 u0_u14_u2_U10 (.ZN( u0_u14_u2_n109 ) , .A2( u0_u14_u2_n113 ) , .B2( u0_u14_u2_n133 ) , .B1( u0_u14_u2_n167 ) , .A1( u0_u14_u2_n168 ) );
  NAND3_X1 u0_u14_u2_U100 (.A2( u0_u14_u2_n100 ) , .A1( u0_u14_u2_n104 ) , .A3( u0_u14_u2_n138 ) , .ZN( u0_u14_u2_n98 ) );
  OAI22_X1 u0_u14_u2_U11 (.B1( u0_u14_u2_n151 ) , .A2( u0_u14_u2_n152 ) , .A1( u0_u14_u2_n153 ) , .ZN( u0_u14_u2_n160 ) , .B2( u0_u14_u2_n168 ) );
  NOR3_X1 u0_u14_u2_U12 (.A1( u0_u14_u2_n150 ) , .ZN( u0_u14_u2_n151 ) , .A3( u0_u14_u2_n175 ) , .A2( u0_u14_u2_n188 ) );
  AOI21_X1 u0_u14_u2_U13 (.ZN( u0_u14_u2_n144 ) , .B2( u0_u14_u2_n155 ) , .A( u0_u14_u2_n172 ) , .B1( u0_u14_u2_n185 ) );
  AOI21_X1 u0_u14_u2_U14 (.B2( u0_u14_u2_n143 ) , .ZN( u0_u14_u2_n145 ) , .B1( u0_u14_u2_n152 ) , .A( u0_u14_u2_n171 ) );
  AOI21_X1 u0_u14_u2_U15 (.B2( u0_u14_u2_n120 ) , .B1( u0_u14_u2_n121 ) , .ZN( u0_u14_u2_n126 ) , .A( u0_u14_u2_n167 ) );
  INV_X1 u0_u14_u2_U16 (.A( u0_u14_u2_n156 ) , .ZN( u0_u14_u2_n171 ) );
  INV_X1 u0_u14_u2_U17 (.A( u0_u14_u2_n120 ) , .ZN( u0_u14_u2_n188 ) );
  NAND2_X1 u0_u14_u2_U18 (.A2( u0_u14_u2_n122 ) , .ZN( u0_u14_u2_n150 ) , .A1( u0_u14_u2_n152 ) );
  INV_X1 u0_u14_u2_U19 (.A( u0_u14_u2_n153 ) , .ZN( u0_u14_u2_n170 ) );
  INV_X1 u0_u14_u2_U20 (.A( u0_u14_u2_n137 ) , .ZN( u0_u14_u2_n173 ) );
  NAND2_X1 u0_u14_u2_U21 (.A1( u0_u14_u2_n132 ) , .A2( u0_u14_u2_n139 ) , .ZN( u0_u14_u2_n157 ) );
  INV_X1 u0_u14_u2_U22 (.A( u0_u14_u2_n113 ) , .ZN( u0_u14_u2_n178 ) );
  INV_X1 u0_u14_u2_U23 (.A( u0_u14_u2_n139 ) , .ZN( u0_u14_u2_n175 ) );
  INV_X1 u0_u14_u2_U24 (.A( u0_u14_u2_n155 ) , .ZN( u0_u14_u2_n181 ) );
  INV_X1 u0_u14_u2_U25 (.A( u0_u14_u2_n119 ) , .ZN( u0_u14_u2_n177 ) );
  INV_X1 u0_u14_u2_U26 (.A( u0_u14_u2_n116 ) , .ZN( u0_u14_u2_n180 ) );
  INV_X1 u0_u14_u2_U27 (.A( u0_u14_u2_n131 ) , .ZN( u0_u14_u2_n179 ) );
  INV_X1 u0_u14_u2_U28 (.A( u0_u14_u2_n154 ) , .ZN( u0_u14_u2_n176 ) );
  NAND2_X1 u0_u14_u2_U29 (.A2( u0_u14_u2_n116 ) , .A1( u0_u14_u2_n117 ) , .ZN( u0_u14_u2_n118 ) );
  NOR2_X1 u0_u14_u2_U3 (.ZN( u0_u14_u2_n121 ) , .A2( u0_u14_u2_n177 ) , .A1( u0_u14_u2_n180 ) );
  INV_X1 u0_u14_u2_U30 (.A( u0_u14_u2_n132 ) , .ZN( u0_u14_u2_n182 ) );
  INV_X1 u0_u14_u2_U31 (.A( u0_u14_u2_n158 ) , .ZN( u0_u14_u2_n183 ) );
  OAI21_X1 u0_u14_u2_U32 (.A( u0_u14_u2_n156 ) , .B1( u0_u14_u2_n157 ) , .ZN( u0_u14_u2_n158 ) , .B2( u0_u14_u2_n179 ) );
  NOR2_X1 u0_u14_u2_U33 (.ZN( u0_u14_u2_n156 ) , .A1( u0_u14_u2_n166 ) , .A2( u0_u14_u2_n169 ) );
  NOR2_X1 u0_u14_u2_U34 (.A2( u0_u14_u2_n114 ) , .ZN( u0_u14_u2_n137 ) , .A1( u0_u14_u2_n140 ) );
  NOR2_X1 u0_u14_u2_U35 (.A2( u0_u14_u2_n138 ) , .ZN( u0_u14_u2_n153 ) , .A1( u0_u14_u2_n156 ) );
  AOI211_X1 u0_u14_u2_U36 (.ZN( u0_u14_u2_n130 ) , .C1( u0_u14_u2_n138 ) , .C2( u0_u14_u2_n179 ) , .B( u0_u14_u2_n96 ) , .A( u0_u14_u2_n97 ) );
  OAI22_X1 u0_u14_u2_U37 (.B1( u0_u14_u2_n133 ) , .A2( u0_u14_u2_n137 ) , .A1( u0_u14_u2_n152 ) , .B2( u0_u14_u2_n168 ) , .ZN( u0_u14_u2_n97 ) );
  OAI221_X1 u0_u14_u2_U38 (.B1( u0_u14_u2_n113 ) , .C1( u0_u14_u2_n132 ) , .A( u0_u14_u2_n149 ) , .B2( u0_u14_u2_n171 ) , .C2( u0_u14_u2_n172 ) , .ZN( u0_u14_u2_n96 ) );
  OAI221_X1 u0_u14_u2_U39 (.A( u0_u14_u2_n115 ) , .C2( u0_u14_u2_n123 ) , .B2( u0_u14_u2_n143 ) , .B1( u0_u14_u2_n153 ) , .ZN( u0_u14_u2_n163 ) , .C1( u0_u14_u2_n168 ) );
  INV_X1 u0_u14_u2_U4 (.A( u0_u14_u2_n134 ) , .ZN( u0_u14_u2_n185 ) );
  OAI21_X1 u0_u14_u2_U40 (.A( u0_u14_u2_n114 ) , .ZN( u0_u14_u2_n115 ) , .B1( u0_u14_u2_n176 ) , .B2( u0_u14_u2_n178 ) );
  OAI221_X1 u0_u14_u2_U41 (.A( u0_u14_u2_n135 ) , .B2( u0_u14_u2_n136 ) , .B1( u0_u14_u2_n137 ) , .ZN( u0_u14_u2_n162 ) , .C2( u0_u14_u2_n167 ) , .C1( u0_u14_u2_n185 ) );
  AND3_X1 u0_u14_u2_U42 (.A3( u0_u14_u2_n131 ) , .A2( u0_u14_u2_n132 ) , .A1( u0_u14_u2_n133 ) , .ZN( u0_u14_u2_n136 ) );
  AOI22_X1 u0_u14_u2_U43 (.ZN( u0_u14_u2_n135 ) , .B1( u0_u14_u2_n140 ) , .A1( u0_u14_u2_n156 ) , .B2( u0_u14_u2_n180 ) , .A2( u0_u14_u2_n188 ) );
  AOI21_X1 u0_u14_u2_U44 (.ZN( u0_u14_u2_n149 ) , .B1( u0_u14_u2_n173 ) , .B2( u0_u14_u2_n188 ) , .A( u0_u14_u2_n95 ) );
  AND3_X1 u0_u14_u2_U45 (.A2( u0_u14_u2_n100 ) , .A1( u0_u14_u2_n104 ) , .A3( u0_u14_u2_n156 ) , .ZN( u0_u14_u2_n95 ) );
  OAI21_X1 u0_u14_u2_U46 (.A( u0_u14_u2_n141 ) , .B2( u0_u14_u2_n142 ) , .ZN( u0_u14_u2_n146 ) , .B1( u0_u14_u2_n153 ) );
  OAI21_X1 u0_u14_u2_U47 (.A( u0_u14_u2_n140 ) , .ZN( u0_u14_u2_n141 ) , .B1( u0_u14_u2_n176 ) , .B2( u0_u14_u2_n177 ) );
  NOR3_X1 u0_u14_u2_U48 (.ZN( u0_u14_u2_n142 ) , .A3( u0_u14_u2_n175 ) , .A2( u0_u14_u2_n178 ) , .A1( u0_u14_u2_n181 ) );
  OAI21_X1 u0_u14_u2_U49 (.A( u0_u14_u2_n101 ) , .B2( u0_u14_u2_n121 ) , .B1( u0_u14_u2_n153 ) , .ZN( u0_u14_u2_n164 ) );
  INV_X1 u0_u14_u2_U5 (.A( u0_u14_u2_n150 ) , .ZN( u0_u14_u2_n184 ) );
  NAND2_X1 u0_u14_u2_U50 (.A2( u0_u14_u2_n100 ) , .A1( u0_u14_u2_n107 ) , .ZN( u0_u14_u2_n155 ) );
  NAND2_X1 u0_u14_u2_U51 (.A2( u0_u14_u2_n105 ) , .A1( u0_u14_u2_n108 ) , .ZN( u0_u14_u2_n143 ) );
  NAND2_X1 u0_u14_u2_U52 (.A1( u0_u14_u2_n104 ) , .A2( u0_u14_u2_n106 ) , .ZN( u0_u14_u2_n152 ) );
  NAND2_X1 u0_u14_u2_U53 (.A1( u0_u14_u2_n100 ) , .A2( u0_u14_u2_n105 ) , .ZN( u0_u14_u2_n132 ) );
  INV_X1 u0_u14_u2_U54 (.A( u0_u14_u2_n140 ) , .ZN( u0_u14_u2_n168 ) );
  INV_X1 u0_u14_u2_U55 (.A( u0_u14_u2_n138 ) , .ZN( u0_u14_u2_n167 ) );
  INV_X1 u0_u14_u2_U56 (.ZN( u0_u14_u2_n187 ) , .A( u0_u14_u2_n99 ) );
  OAI21_X1 u0_u14_u2_U57 (.B1( u0_u14_u2_n137 ) , .B2( u0_u14_u2_n143 ) , .A( u0_u14_u2_n98 ) , .ZN( u0_u14_u2_n99 ) );
  NAND2_X1 u0_u14_u2_U58 (.A1( u0_u14_u2_n102 ) , .A2( u0_u14_u2_n106 ) , .ZN( u0_u14_u2_n113 ) );
  NAND2_X1 u0_u14_u2_U59 (.A1( u0_u14_u2_n106 ) , .A2( u0_u14_u2_n107 ) , .ZN( u0_u14_u2_n131 ) );
  NOR4_X1 u0_u14_u2_U6 (.A4( u0_u14_u2_n124 ) , .A3( u0_u14_u2_n125 ) , .A2( u0_u14_u2_n126 ) , .A1( u0_u14_u2_n127 ) , .ZN( u0_u14_u2_n128 ) );
  NAND2_X1 u0_u14_u2_U60 (.A1( u0_u14_u2_n103 ) , .A2( u0_u14_u2_n107 ) , .ZN( u0_u14_u2_n139 ) );
  NAND2_X1 u0_u14_u2_U61 (.A1( u0_u14_u2_n103 ) , .A2( u0_u14_u2_n105 ) , .ZN( u0_u14_u2_n133 ) );
  NAND2_X1 u0_u14_u2_U62 (.A1( u0_u14_u2_n102 ) , .A2( u0_u14_u2_n103 ) , .ZN( u0_u14_u2_n154 ) );
  NAND2_X1 u0_u14_u2_U63 (.A2( u0_u14_u2_n103 ) , .A1( u0_u14_u2_n104 ) , .ZN( u0_u14_u2_n119 ) );
  NAND2_X1 u0_u14_u2_U64 (.A2( u0_u14_u2_n107 ) , .A1( u0_u14_u2_n108 ) , .ZN( u0_u14_u2_n123 ) );
  NAND2_X1 u0_u14_u2_U65 (.A1( u0_u14_u2_n104 ) , .A2( u0_u14_u2_n108 ) , .ZN( u0_u14_u2_n122 ) );
  INV_X1 u0_u14_u2_U66 (.A( u0_u14_u2_n114 ) , .ZN( u0_u14_u2_n172 ) );
  NAND2_X1 u0_u14_u2_U67 (.A2( u0_u14_u2_n100 ) , .A1( u0_u14_u2_n102 ) , .ZN( u0_u14_u2_n116 ) );
  NAND2_X1 u0_u14_u2_U68 (.A1( u0_u14_u2_n102 ) , .A2( u0_u14_u2_n108 ) , .ZN( u0_u14_u2_n120 ) );
  NAND2_X1 u0_u14_u2_U69 (.A2( u0_u14_u2_n105 ) , .A1( u0_u14_u2_n106 ) , .ZN( u0_u14_u2_n117 ) );
  AOI21_X1 u0_u14_u2_U7 (.B2( u0_u14_u2_n119 ) , .ZN( u0_u14_u2_n127 ) , .A( u0_u14_u2_n137 ) , .B1( u0_u14_u2_n155 ) );
  NOR2_X1 u0_u14_u2_U70 (.A2( u0_u14_X_16 ) , .ZN( u0_u14_u2_n140 ) , .A1( u0_u14_u2_n166 ) );
  NOR2_X1 u0_u14_u2_U71 (.A2( u0_u14_X_13 ) , .A1( u0_u14_X_14 ) , .ZN( u0_u14_u2_n100 ) );
  NOR2_X1 u0_u14_u2_U72 (.A2( u0_u14_X_16 ) , .A1( u0_u14_X_17 ) , .ZN( u0_u14_u2_n138 ) );
  NOR2_X1 u0_u14_u2_U73 (.A2( u0_u14_X_15 ) , .A1( u0_u14_X_18 ) , .ZN( u0_u14_u2_n104 ) );
  NOR2_X1 u0_u14_u2_U74 (.A2( u0_u14_X_14 ) , .ZN( u0_u14_u2_n103 ) , .A1( u0_u14_u2_n174 ) );
  NOR2_X1 u0_u14_u2_U75 (.A2( u0_u14_X_15 ) , .ZN( u0_u14_u2_n102 ) , .A1( u0_u14_u2_n165 ) );
  NOR2_X1 u0_u14_u2_U76 (.A2( u0_u14_X_17 ) , .ZN( u0_u14_u2_n114 ) , .A1( u0_u14_u2_n169 ) );
  AND2_X1 u0_u14_u2_U77 (.A1( u0_u14_X_15 ) , .ZN( u0_u14_u2_n105 ) , .A2( u0_u14_u2_n165 ) );
  AND2_X1 u0_u14_u2_U78 (.A2( u0_u14_X_15 ) , .A1( u0_u14_X_18 ) , .ZN( u0_u14_u2_n107 ) );
  AND2_X1 u0_u14_u2_U79 (.A1( u0_u14_X_14 ) , .ZN( u0_u14_u2_n106 ) , .A2( u0_u14_u2_n174 ) );
  AOI21_X1 u0_u14_u2_U8 (.ZN( u0_u14_u2_n124 ) , .B1( u0_u14_u2_n131 ) , .B2( u0_u14_u2_n143 ) , .A( u0_u14_u2_n172 ) );
  AND2_X1 u0_u14_u2_U80 (.A1( u0_u14_X_13 ) , .A2( u0_u14_X_14 ) , .ZN( u0_u14_u2_n108 ) );
  INV_X1 u0_u14_u2_U81 (.A( u0_u14_X_16 ) , .ZN( u0_u14_u2_n169 ) );
  INV_X1 u0_u14_u2_U82 (.A( u0_u14_X_17 ) , .ZN( u0_u14_u2_n166 ) );
  INV_X1 u0_u14_u2_U83 (.A( u0_u14_X_13 ) , .ZN( u0_u14_u2_n174 ) );
  INV_X1 u0_u14_u2_U84 (.A( u0_u14_X_18 ) , .ZN( u0_u14_u2_n165 ) );
  NAND4_X1 u0_u14_u2_U85 (.ZN( u0_out14_30 ) , .A4( u0_u14_u2_n147 ) , .A3( u0_u14_u2_n148 ) , .A2( u0_u14_u2_n149 ) , .A1( u0_u14_u2_n187 ) );
  NOR3_X1 u0_u14_u2_U86 (.A3( u0_u14_u2_n144 ) , .A2( u0_u14_u2_n145 ) , .A1( u0_u14_u2_n146 ) , .ZN( u0_u14_u2_n147 ) );
  AOI21_X1 u0_u14_u2_U87 (.B2( u0_u14_u2_n138 ) , .ZN( u0_u14_u2_n148 ) , .A( u0_u14_u2_n162 ) , .B1( u0_u14_u2_n182 ) );
  NAND4_X1 u0_u14_u2_U88 (.ZN( u0_out14_24 ) , .A4( u0_u14_u2_n111 ) , .A3( u0_u14_u2_n112 ) , .A1( u0_u14_u2_n130 ) , .A2( u0_u14_u2_n187 ) );
  AOI221_X1 u0_u14_u2_U89 (.A( u0_u14_u2_n109 ) , .B1( u0_u14_u2_n110 ) , .ZN( u0_u14_u2_n111 ) , .C1( u0_u14_u2_n134 ) , .C2( u0_u14_u2_n170 ) , .B2( u0_u14_u2_n173 ) );
  AOI21_X1 u0_u14_u2_U9 (.B2( u0_u14_u2_n123 ) , .ZN( u0_u14_u2_n125 ) , .A( u0_u14_u2_n171 ) , .B1( u0_u14_u2_n184 ) );
  AOI21_X1 u0_u14_u2_U90 (.ZN( u0_u14_u2_n112 ) , .B2( u0_u14_u2_n156 ) , .A( u0_u14_u2_n164 ) , .B1( u0_u14_u2_n181 ) );
  NAND4_X1 u0_u14_u2_U91 (.ZN( u0_out14_16 ) , .A4( u0_u14_u2_n128 ) , .A3( u0_u14_u2_n129 ) , .A1( u0_u14_u2_n130 ) , .A2( u0_u14_u2_n186 ) );
  AOI22_X1 u0_u14_u2_U92 (.A2( u0_u14_u2_n118 ) , .ZN( u0_u14_u2_n129 ) , .A1( u0_u14_u2_n140 ) , .B1( u0_u14_u2_n157 ) , .B2( u0_u14_u2_n170 ) );
  INV_X1 u0_u14_u2_U93 (.A( u0_u14_u2_n163 ) , .ZN( u0_u14_u2_n186 ) );
  OR4_X1 u0_u14_u2_U94 (.ZN( u0_out14_6 ) , .A4( u0_u14_u2_n161 ) , .A3( u0_u14_u2_n162 ) , .A2( u0_u14_u2_n163 ) , .A1( u0_u14_u2_n164 ) );
  OR3_X1 u0_u14_u2_U95 (.A2( u0_u14_u2_n159 ) , .A1( u0_u14_u2_n160 ) , .ZN( u0_u14_u2_n161 ) , .A3( u0_u14_u2_n183 ) );
  AOI21_X1 u0_u14_u2_U96 (.B2( u0_u14_u2_n154 ) , .B1( u0_u14_u2_n155 ) , .ZN( u0_u14_u2_n159 ) , .A( u0_u14_u2_n167 ) );
  NAND3_X1 u0_u14_u2_U97 (.A2( u0_u14_u2_n117 ) , .A1( u0_u14_u2_n122 ) , .A3( u0_u14_u2_n123 ) , .ZN( u0_u14_u2_n134 ) );
  NAND3_X1 u0_u14_u2_U98 (.ZN( u0_u14_u2_n110 ) , .A2( u0_u14_u2_n131 ) , .A3( u0_u14_u2_n139 ) , .A1( u0_u14_u2_n154 ) );
  NAND3_X1 u0_u14_u2_U99 (.A2( u0_u14_u2_n100 ) , .ZN( u0_u14_u2_n101 ) , .A1( u0_u14_u2_n104 ) , .A3( u0_u14_u2_n114 ) );
  XOR2_X1 u0_u5_U10 (.B( u0_K6_45 ) , .A( u0_R4_30 ) , .Z( u0_u5_X_45 ) );
  XOR2_X1 u0_u5_U11 (.B( u0_K6_44 ) , .A( u0_R4_29 ) , .Z( u0_u5_X_44 ) );
  XOR2_X1 u0_u5_U12 (.B( u0_K6_43 ) , .A( u0_R4_28 ) , .Z( u0_u5_X_43 ) );
  XOR2_X1 u0_u5_U7 (.B( u0_K6_48 ) , .A( u0_R4_1 ) , .Z( u0_u5_X_48 ) );
  XOR2_X1 u0_u5_U8 (.B( u0_K6_47 ) , .A( u0_R4_32 ) , .Z( u0_u5_X_47 ) );
  XOR2_X1 u0_u5_U9 (.B( u0_K6_46 ) , .A( u0_R4_31 ) , .Z( u0_u5_X_46 ) );
  AND3_X1 u0_u5_u7_U10 (.A3( u0_u5_u7_n110 ) , .A2( u0_u5_u7_n127 ) , .A1( u0_u5_u7_n132 ) , .ZN( u0_u5_u7_n92 ) );
  OAI21_X1 u0_u5_u7_U11 (.A( u0_u5_u7_n161 ) , .B1( u0_u5_u7_n168 ) , .B2( u0_u5_u7_n173 ) , .ZN( u0_u5_u7_n91 ) );
  AOI211_X1 u0_u5_u7_U12 (.A( u0_u5_u7_n117 ) , .ZN( u0_u5_u7_n118 ) , .C2( u0_u5_u7_n126 ) , .C1( u0_u5_u7_n177 ) , .B( u0_u5_u7_n180 ) );
  OAI22_X1 u0_u5_u7_U13 (.B1( u0_u5_u7_n115 ) , .ZN( u0_u5_u7_n117 ) , .A2( u0_u5_u7_n133 ) , .A1( u0_u5_u7_n137 ) , .B2( u0_u5_u7_n162 ) );
  INV_X1 u0_u5_u7_U14 (.A( u0_u5_u7_n116 ) , .ZN( u0_u5_u7_n180 ) );
  NOR3_X1 u0_u5_u7_U15 (.ZN( u0_u5_u7_n115 ) , .A3( u0_u5_u7_n145 ) , .A2( u0_u5_u7_n168 ) , .A1( u0_u5_u7_n169 ) );
  OAI211_X1 u0_u5_u7_U16 (.B( u0_u5_u7_n122 ) , .A( u0_u5_u7_n123 ) , .C2( u0_u5_u7_n124 ) , .ZN( u0_u5_u7_n154 ) , .C1( u0_u5_u7_n162 ) );
  AOI222_X1 u0_u5_u7_U17 (.ZN( u0_u5_u7_n122 ) , .C2( u0_u5_u7_n126 ) , .C1( u0_u5_u7_n145 ) , .B1( u0_u5_u7_n161 ) , .A2( u0_u5_u7_n165 ) , .B2( u0_u5_u7_n170 ) , .A1( u0_u5_u7_n176 ) );
  INV_X1 u0_u5_u7_U18 (.A( u0_u5_u7_n133 ) , .ZN( u0_u5_u7_n176 ) );
  NOR3_X1 u0_u5_u7_U19 (.A2( u0_u5_u7_n134 ) , .A1( u0_u5_u7_n135 ) , .ZN( u0_u5_u7_n136 ) , .A3( u0_u5_u7_n171 ) );
  NOR2_X1 u0_u5_u7_U20 (.A1( u0_u5_u7_n130 ) , .A2( u0_u5_u7_n134 ) , .ZN( u0_u5_u7_n153 ) );
  INV_X1 u0_u5_u7_U21 (.A( u0_u5_u7_n101 ) , .ZN( u0_u5_u7_n165 ) );
  NOR2_X1 u0_u5_u7_U22 (.ZN( u0_u5_u7_n111 ) , .A2( u0_u5_u7_n134 ) , .A1( u0_u5_u7_n169 ) );
  AOI21_X1 u0_u5_u7_U23 (.ZN( u0_u5_u7_n104 ) , .B2( u0_u5_u7_n112 ) , .B1( u0_u5_u7_n127 ) , .A( u0_u5_u7_n164 ) );
  AOI21_X1 u0_u5_u7_U24 (.ZN( u0_u5_u7_n106 ) , .B1( u0_u5_u7_n133 ) , .B2( u0_u5_u7_n146 ) , .A( u0_u5_u7_n162 ) );
  AOI21_X1 u0_u5_u7_U25 (.A( u0_u5_u7_n101 ) , .ZN( u0_u5_u7_n107 ) , .B2( u0_u5_u7_n128 ) , .B1( u0_u5_u7_n175 ) );
  INV_X1 u0_u5_u7_U26 (.A( u0_u5_u7_n138 ) , .ZN( u0_u5_u7_n171 ) );
  INV_X1 u0_u5_u7_U27 (.A( u0_u5_u7_n131 ) , .ZN( u0_u5_u7_n177 ) );
  INV_X1 u0_u5_u7_U28 (.A( u0_u5_u7_n110 ) , .ZN( u0_u5_u7_n174 ) );
  NAND2_X1 u0_u5_u7_U29 (.A1( u0_u5_u7_n129 ) , .A2( u0_u5_u7_n132 ) , .ZN( u0_u5_u7_n149 ) );
  OAI21_X1 u0_u5_u7_U3 (.ZN( u0_u5_u7_n159 ) , .A( u0_u5_u7_n165 ) , .B2( u0_u5_u7_n171 ) , .B1( u0_u5_u7_n174 ) );
  NAND2_X1 u0_u5_u7_U30 (.A1( u0_u5_u7_n113 ) , .A2( u0_u5_u7_n124 ) , .ZN( u0_u5_u7_n130 ) );
  INV_X1 u0_u5_u7_U31 (.A( u0_u5_u7_n112 ) , .ZN( u0_u5_u7_n173 ) );
  INV_X1 u0_u5_u7_U32 (.A( u0_u5_u7_n128 ) , .ZN( u0_u5_u7_n168 ) );
  INV_X1 u0_u5_u7_U33 (.A( u0_u5_u7_n148 ) , .ZN( u0_u5_u7_n169 ) );
  INV_X1 u0_u5_u7_U34 (.A( u0_u5_u7_n127 ) , .ZN( u0_u5_u7_n179 ) );
  NOR2_X1 u0_u5_u7_U35 (.ZN( u0_u5_u7_n101 ) , .A2( u0_u5_u7_n150 ) , .A1( u0_u5_u7_n156 ) );
  AOI211_X1 u0_u5_u7_U36 (.B( u0_u5_u7_n154 ) , .A( u0_u5_u7_n155 ) , .C1( u0_u5_u7_n156 ) , .ZN( u0_u5_u7_n157 ) , .C2( u0_u5_u7_n172 ) );
  INV_X1 u0_u5_u7_U37 (.A( u0_u5_u7_n153 ) , .ZN( u0_u5_u7_n172 ) );
  AOI211_X1 u0_u5_u7_U38 (.B( u0_u5_u7_n139 ) , .A( u0_u5_u7_n140 ) , .C2( u0_u5_u7_n141 ) , .ZN( u0_u5_u7_n142 ) , .C1( u0_u5_u7_n156 ) );
  NAND4_X1 u0_u5_u7_U39 (.A3( u0_u5_u7_n127 ) , .A2( u0_u5_u7_n128 ) , .A1( u0_u5_u7_n129 ) , .ZN( u0_u5_u7_n141 ) , .A4( u0_u5_u7_n147 ) );
  INV_X1 u0_u5_u7_U4 (.A( u0_u5_u7_n111 ) , .ZN( u0_u5_u7_n170 ) );
  AOI21_X1 u0_u5_u7_U40 (.A( u0_u5_u7_n137 ) , .B1( u0_u5_u7_n138 ) , .ZN( u0_u5_u7_n139 ) , .B2( u0_u5_u7_n146 ) );
  OAI22_X1 u0_u5_u7_U41 (.B1( u0_u5_u7_n136 ) , .ZN( u0_u5_u7_n140 ) , .A1( u0_u5_u7_n153 ) , .B2( u0_u5_u7_n162 ) , .A2( u0_u5_u7_n164 ) );
  AOI21_X1 u0_u5_u7_U42 (.ZN( u0_u5_u7_n123 ) , .B1( u0_u5_u7_n165 ) , .B2( u0_u5_u7_n177 ) , .A( u0_u5_u7_n97 ) );
  AOI21_X1 u0_u5_u7_U43 (.B2( u0_u5_u7_n113 ) , .B1( u0_u5_u7_n124 ) , .A( u0_u5_u7_n125 ) , .ZN( u0_u5_u7_n97 ) );
  INV_X1 u0_u5_u7_U44 (.A( u0_u5_u7_n125 ) , .ZN( u0_u5_u7_n161 ) );
  INV_X1 u0_u5_u7_U45 (.A( u0_u5_u7_n152 ) , .ZN( u0_u5_u7_n162 ) );
  AOI22_X1 u0_u5_u7_U46 (.A2( u0_u5_u7_n114 ) , .ZN( u0_u5_u7_n119 ) , .B1( u0_u5_u7_n130 ) , .A1( u0_u5_u7_n156 ) , .B2( u0_u5_u7_n165 ) );
  NAND2_X1 u0_u5_u7_U47 (.A2( u0_u5_u7_n112 ) , .ZN( u0_u5_u7_n114 ) , .A1( u0_u5_u7_n175 ) );
  AND2_X1 u0_u5_u7_U48 (.ZN( u0_u5_u7_n145 ) , .A2( u0_u5_u7_n98 ) , .A1( u0_u5_u7_n99 ) );
  NOR2_X1 u0_u5_u7_U49 (.ZN( u0_u5_u7_n137 ) , .A1( u0_u5_u7_n150 ) , .A2( u0_u5_u7_n161 ) );
  INV_X1 u0_u5_u7_U5 (.A( u0_u5_u7_n149 ) , .ZN( u0_u5_u7_n175 ) );
  AOI21_X1 u0_u5_u7_U50 (.ZN( u0_u5_u7_n105 ) , .B2( u0_u5_u7_n110 ) , .A( u0_u5_u7_n125 ) , .B1( u0_u5_u7_n147 ) );
  NAND2_X1 u0_u5_u7_U51 (.ZN( u0_u5_u7_n146 ) , .A1( u0_u5_u7_n95 ) , .A2( u0_u5_u7_n98 ) );
  NAND2_X1 u0_u5_u7_U52 (.A2( u0_u5_u7_n103 ) , .ZN( u0_u5_u7_n147 ) , .A1( u0_u5_u7_n93 ) );
  NAND2_X1 u0_u5_u7_U53 (.A1( u0_u5_u7_n103 ) , .ZN( u0_u5_u7_n127 ) , .A2( u0_u5_u7_n99 ) );
  OR2_X1 u0_u5_u7_U54 (.ZN( u0_u5_u7_n126 ) , .A2( u0_u5_u7_n152 ) , .A1( u0_u5_u7_n156 ) );
  NAND2_X1 u0_u5_u7_U55 (.A2( u0_u5_u7_n102 ) , .A1( u0_u5_u7_n103 ) , .ZN( u0_u5_u7_n133 ) );
  NAND2_X1 u0_u5_u7_U56 (.ZN( u0_u5_u7_n112 ) , .A2( u0_u5_u7_n96 ) , .A1( u0_u5_u7_n99 ) );
  NAND2_X1 u0_u5_u7_U57 (.A2( u0_u5_u7_n102 ) , .ZN( u0_u5_u7_n128 ) , .A1( u0_u5_u7_n98 ) );
  NAND2_X1 u0_u5_u7_U58 (.A1( u0_u5_u7_n100 ) , .ZN( u0_u5_u7_n113 ) , .A2( u0_u5_u7_n93 ) );
  NAND2_X1 u0_u5_u7_U59 (.A2( u0_u5_u7_n102 ) , .ZN( u0_u5_u7_n124 ) , .A1( u0_u5_u7_n96 ) );
  INV_X1 u0_u5_u7_U6 (.A( u0_u5_u7_n154 ) , .ZN( u0_u5_u7_n178 ) );
  NAND2_X1 u0_u5_u7_U60 (.ZN( u0_u5_u7_n110 ) , .A1( u0_u5_u7_n95 ) , .A2( u0_u5_u7_n96 ) );
  INV_X1 u0_u5_u7_U61 (.A( u0_u5_u7_n150 ) , .ZN( u0_u5_u7_n164 ) );
  AND2_X1 u0_u5_u7_U62 (.ZN( u0_u5_u7_n134 ) , .A1( u0_u5_u7_n93 ) , .A2( u0_u5_u7_n98 ) );
  NAND2_X1 u0_u5_u7_U63 (.A1( u0_u5_u7_n100 ) , .A2( u0_u5_u7_n102 ) , .ZN( u0_u5_u7_n129 ) );
  NAND2_X1 u0_u5_u7_U64 (.A2( u0_u5_u7_n103 ) , .ZN( u0_u5_u7_n131 ) , .A1( u0_u5_u7_n95 ) );
  NAND2_X1 u0_u5_u7_U65 (.A1( u0_u5_u7_n100 ) , .ZN( u0_u5_u7_n138 ) , .A2( u0_u5_u7_n99 ) );
  NAND2_X1 u0_u5_u7_U66 (.ZN( u0_u5_u7_n132 ) , .A1( u0_u5_u7_n93 ) , .A2( u0_u5_u7_n96 ) );
  NAND2_X1 u0_u5_u7_U67 (.A1( u0_u5_u7_n100 ) , .ZN( u0_u5_u7_n148 ) , .A2( u0_u5_u7_n95 ) );
  NOR2_X1 u0_u5_u7_U68 (.A2( u0_u5_X_47 ) , .ZN( u0_u5_u7_n150 ) , .A1( u0_u5_u7_n163 ) );
  NOR2_X1 u0_u5_u7_U69 (.A2( u0_u5_X_43 ) , .A1( u0_u5_X_44 ) , .ZN( u0_u5_u7_n103 ) );
  AOI211_X1 u0_u5_u7_U7 (.ZN( u0_u5_u7_n116 ) , .A( u0_u5_u7_n155 ) , .C1( u0_u5_u7_n161 ) , .C2( u0_u5_u7_n171 ) , .B( u0_u5_u7_n94 ) );
  NOR2_X1 u0_u5_u7_U70 (.A2( u0_u5_X_48 ) , .A1( u0_u5_u7_n166 ) , .ZN( u0_u5_u7_n95 ) );
  NOR2_X1 u0_u5_u7_U71 (.A2( u0_u5_X_45 ) , .A1( u0_u5_X_48 ) , .ZN( u0_u5_u7_n99 ) );
  NOR2_X1 u0_u5_u7_U72 (.A2( u0_u5_X_44 ) , .A1( u0_u5_u7_n167 ) , .ZN( u0_u5_u7_n98 ) );
  NOR2_X1 u0_u5_u7_U73 (.A2( u0_u5_X_46 ) , .A1( u0_u5_X_47 ) , .ZN( u0_u5_u7_n152 ) );
  AND2_X1 u0_u5_u7_U74 (.A1( u0_u5_X_47 ) , .ZN( u0_u5_u7_n156 ) , .A2( u0_u5_u7_n163 ) );
  NAND2_X1 u0_u5_u7_U75 (.A2( u0_u5_X_46 ) , .A1( u0_u5_X_47 ) , .ZN( u0_u5_u7_n125 ) );
  AND2_X1 u0_u5_u7_U76 (.A2( u0_u5_X_45 ) , .A1( u0_u5_X_48 ) , .ZN( u0_u5_u7_n102 ) );
  AND2_X1 u0_u5_u7_U77 (.A2( u0_u5_X_43 ) , .A1( u0_u5_X_44 ) , .ZN( u0_u5_u7_n96 ) );
  AND2_X1 u0_u5_u7_U78 (.A1( u0_u5_X_44 ) , .ZN( u0_u5_u7_n100 ) , .A2( u0_u5_u7_n167 ) );
  AND2_X1 u0_u5_u7_U79 (.A1( u0_u5_X_48 ) , .A2( u0_u5_u7_n166 ) , .ZN( u0_u5_u7_n93 ) );
  OAI222_X1 u0_u5_u7_U8 (.C2( u0_u5_u7_n101 ) , .B2( u0_u5_u7_n111 ) , .A1( u0_u5_u7_n113 ) , .C1( u0_u5_u7_n146 ) , .A2( u0_u5_u7_n162 ) , .B1( u0_u5_u7_n164 ) , .ZN( u0_u5_u7_n94 ) );
  INV_X1 u0_u5_u7_U80 (.A( u0_u5_X_46 ) , .ZN( u0_u5_u7_n163 ) );
  INV_X1 u0_u5_u7_U81 (.A( u0_u5_X_43 ) , .ZN( u0_u5_u7_n167 ) );
  INV_X1 u0_u5_u7_U82 (.A( u0_u5_X_45 ) , .ZN( u0_u5_u7_n166 ) );
  NAND4_X1 u0_u5_u7_U83 (.ZN( u0_out5_27 ) , .A4( u0_u5_u7_n118 ) , .A3( u0_u5_u7_n119 ) , .A2( u0_u5_u7_n120 ) , .A1( u0_u5_u7_n121 ) );
  OAI21_X1 u0_u5_u7_U84 (.ZN( u0_u5_u7_n121 ) , .B2( u0_u5_u7_n145 ) , .A( u0_u5_u7_n150 ) , .B1( u0_u5_u7_n174 ) );
  OAI21_X1 u0_u5_u7_U85 (.ZN( u0_u5_u7_n120 ) , .A( u0_u5_u7_n161 ) , .B2( u0_u5_u7_n170 ) , .B1( u0_u5_u7_n179 ) );
  NAND4_X1 u0_u5_u7_U86 (.ZN( u0_out5_21 ) , .A4( u0_u5_u7_n157 ) , .A3( u0_u5_u7_n158 ) , .A2( u0_u5_u7_n159 ) , .A1( u0_u5_u7_n160 ) );
  OAI21_X1 u0_u5_u7_U87 (.B1( u0_u5_u7_n145 ) , .ZN( u0_u5_u7_n160 ) , .A( u0_u5_u7_n161 ) , .B2( u0_u5_u7_n177 ) );
  AOI22_X1 u0_u5_u7_U88 (.B2( u0_u5_u7_n149 ) , .B1( u0_u5_u7_n150 ) , .A2( u0_u5_u7_n151 ) , .A1( u0_u5_u7_n152 ) , .ZN( u0_u5_u7_n158 ) );
  NAND4_X1 u0_u5_u7_U89 (.ZN( u0_out5_15 ) , .A4( u0_u5_u7_n142 ) , .A3( u0_u5_u7_n143 ) , .A2( u0_u5_u7_n144 ) , .A1( u0_u5_u7_n178 ) );
  OAI221_X1 u0_u5_u7_U9 (.C1( u0_u5_u7_n101 ) , .C2( u0_u5_u7_n147 ) , .ZN( u0_u5_u7_n155 ) , .B2( u0_u5_u7_n162 ) , .A( u0_u5_u7_n91 ) , .B1( u0_u5_u7_n92 ) );
  OR2_X1 u0_u5_u7_U90 (.A2( u0_u5_u7_n125 ) , .A1( u0_u5_u7_n129 ) , .ZN( u0_u5_u7_n144 ) );
  AOI22_X1 u0_u5_u7_U91 (.A2( u0_u5_u7_n126 ) , .ZN( u0_u5_u7_n143 ) , .B2( u0_u5_u7_n165 ) , .B1( u0_u5_u7_n173 ) , .A1( u0_u5_u7_n174 ) );
  NAND4_X1 u0_u5_u7_U92 (.ZN( u0_out5_5 ) , .A4( u0_u5_u7_n108 ) , .A3( u0_u5_u7_n109 ) , .A1( u0_u5_u7_n116 ) , .A2( u0_u5_u7_n123 ) );
  AOI22_X1 u0_u5_u7_U93 (.ZN( u0_u5_u7_n109 ) , .A2( u0_u5_u7_n126 ) , .B2( u0_u5_u7_n145 ) , .B1( u0_u5_u7_n156 ) , .A1( u0_u5_u7_n171 ) );
  NOR4_X1 u0_u5_u7_U94 (.A4( u0_u5_u7_n104 ) , .A3( u0_u5_u7_n105 ) , .A2( u0_u5_u7_n106 ) , .A1( u0_u5_u7_n107 ) , .ZN( u0_u5_u7_n108 ) );
  NAND3_X1 u0_u5_u7_U95 (.A3( u0_u5_u7_n146 ) , .A2( u0_u5_u7_n147 ) , .A1( u0_u5_u7_n148 ) , .ZN( u0_u5_u7_n151 ) );
  NAND3_X1 u0_u5_u7_U96 (.A3( u0_u5_u7_n131 ) , .A2( u0_u5_u7_n132 ) , .A1( u0_u5_u7_n133 ) , .ZN( u0_u5_u7_n135 ) );
  OAI21_X1 u0_uk_U1020 (.ZN( u0_K14_44 ) , .B1( u0_uk_n163 ) , .B2( u0_uk_n81 ) , .A( u0_uk_n930 ) );
  NAND2_X1 u0_uk_U1021 (.A1( u0_uk_K_r12_15 ) , .A2( u0_uk_n203 ) , .ZN( u0_uk_n930 ) );
  OAI21_X1 u0_uk_U1042 (.ZN( u0_K14_40 ) , .B1( u0_uk_n27 ) , .B2( u0_uk_n65 ) , .A( u0_uk_n931 ) );
  NAND2_X1 u0_uk_U1043 (.A1( u0_uk_K_r12_21 ) , .A2( u0_uk_n110 ) , .ZN( u0_uk_n931 ) );
  OAI21_X1 u0_uk_U1044 (.ZN( u0_K15_14 ) , .B2( u0_uk_n37 ) , .B1( u0_uk_n92 ) , .A( u0_uk_n923 ) );
  NAND2_X1 u0_uk_U1045 (.A1( u0_uk_K_r13_32 ) , .A2( u0_uk_n11 ) , .ZN( u0_uk_n923 ) );
  OAI22_X1 u0_uk_U109 (.ZN( u0_K14_41 ) , .A1( u0_uk_n230 ) , .B2( u0_uk_n77 ) , .A2( u0_uk_n82 ) , .B1( u0_uk_n93 ) );
  INV_X1 u0_uk_U11 (.A( u0_uk_n231 ) , .ZN( u0_uk_n83 ) );
  OAI21_X1 u0_uk_U120 (.ZN( u0_K6_47 ) , .B1( u0_uk_n11 ) , .B2( u0_uk_n439 ) , .A( u0_uk_n789 ) );
  NAND2_X1 u0_uk_U121 (.A1( u0_uk_K_r4_23 ) , .ZN( u0_uk_n789 ) , .A2( u0_uk_n93 ) );
  OAI21_X1 u0_uk_U147 (.ZN( u0_K15_15 ) , .B2( u0_uk_n15 ) , .B1( u0_uk_n163 ) , .A( u0_uk_n922 ) );
  NAND2_X1 u0_uk_U148 (.A1( u0_uk_K_r13_19 ) , .A2( u0_uk_n208 ) , .ZN( u0_uk_n922 ) );
  OAI22_X1 u0_uk_U237 (.ZN( u0_K14_39 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n163 ) , .A2( u0_uk_n52 ) , .B2( u0_uk_n56 ) );
  OAI22_X1 u0_uk_U254 (.ZN( u0_K14_48 ) , .B1( u0_uk_n128 ) , .A1( u0_uk_n230 ) , .A2( u0_uk_n52 ) , .B2( u0_uk_n90 ) );
  OAI22_X1 u0_uk_U268 (.ZN( u0_K6_44 ) , .A1( u0_uk_n109 ) , .B1( u0_uk_n231 ) , .A2( u0_uk_n412 ) , .B2( u0_uk_n430 ) );
  OAI22_X1 u0_uk_U269 (.ZN( u0_K6_48 ) , .A1( u0_uk_n242 ) , .A2( u0_uk_n418 ) , .B2( u0_uk_n425 ) , .B1( u0_uk_n60 ) );
  BUF_X1 u0_uk_U27 (.Z( u0_uk_n163 ) , .A( u0_uk_n217 ) );
  INV_X1 u0_uk_U284 (.ZN( u0_K15_8 ) , .A( u0_uk_n913 ) );
  AOI22_X1 u0_uk_U285 (.B2( u0_uk_K_r13_13 ) , .A2( u0_uk_K_r13_17 ) , .B1( u0_uk_n146 ) , .A1( u0_uk_n230 ) , .ZN( u0_uk_n913 ) );
  OAI22_X1 u0_uk_U337 (.ZN( u0_K15_4 ) , .A1( u0_uk_n100 ) , .B1( u0_uk_n222 ) , .B2( u0_uk_n38 ) , .A2( u0_uk_n8 ) );
  BUF_X1 u0_uk_U36 (.Z( u0_uk_n188 ) , .A( u0_uk_n230 ) );
  OAI22_X1 u0_uk_U387 (.ZN( u0_K14_1 ) , .A1( u0_uk_n118 ) , .B1( u0_uk_n240 ) , .A2( u0_uk_n75 ) , .B2( u0_uk_n80 ) );
  OAI21_X1 u0_uk_U402 (.ZN( u0_K15_9 ) , .B2( u0_uk_n15 ) , .A( u0_uk_n912 ) , .B1( u0_uk_n93 ) );
  NAND2_X1 u0_uk_U403 (.A1( u0_uk_K_r13_4 ) , .A2( u0_uk_n10 ) , .ZN( u0_uk_n912 ) );
  OAI22_X1 u0_uk_U425 (.ZN( u0_K15_1 ) , .A2( u0_uk_n1 ) , .B2( u0_uk_n20 ) , .A1( u0_uk_n230 ) , .B1( u0_uk_n83 ) );
  OAI22_X1 u0_uk_U434 (.ZN( u0_K15_16 ) , .A2( u0_uk_n14 ) , .A1( u0_uk_n188 ) , .B2( u0_uk_n29 ) , .B1( u0_uk_n92 ) );
  OAI22_X1 u0_uk_U451 (.ZN( u0_K14_37 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n231 ) , .A2( u0_uk_n67 ) , .B2( u0_uk_n73 ) );
  OAI22_X1 u0_uk_U488 (.ZN( u0_K14_2 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n231 ) , .A2( u0_uk_n57 ) , .B2( u0_uk_n64 ) );
  BUF_X1 u0_uk_U49 (.Z( u0_uk_n231 ) , .A( u0_uk_n250 ) );
  OAI22_X1 u0_uk_U518 (.ZN( u0_K15_12 ) , .A1( u0_uk_n118 ) , .B1( u0_uk_n231 ) , .B2( u0_uk_n25 ) , .A2( u0_uk_n43 ) );
  OAI22_X1 u0_uk_U529 (.ZN( u0_K15_2 ) , .A2( u0_uk_n1 ) , .A1( u0_uk_n128 ) , .B1( u0_uk_n188 ) , .B2( u0_uk_n30 ) );
  OAI22_X1 u0_uk_U537 (.ZN( u0_K15_17 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n220 ) , .B2( u0_uk_n26 ) , .A2( u0_uk_n44 ) );
  OAI21_X1 u0_uk_U572 (.ZN( u0_K15_10 ) , .B1( u0_uk_n128 ) , .B2( u0_uk_n19 ) , .A( u0_uk_n925 ) );
  NAND2_X1 u0_uk_U573 (.A1( u0_uk_K_r13_55 ) , .A2( u0_uk_n10 ) , .ZN( u0_uk_n925 ) );
  INV_X1 u0_uk_U6 (.A( u0_uk_n231 ) , .ZN( u0_uk_n93 ) );
  OAI21_X1 u0_uk_U624 (.ZN( u0_K15_11 ) , .B1( u0_uk_n163 ) , .B2( u0_uk_n8 ) , .A( u0_uk_n924 ) );
  NAND2_X1 u0_uk_U625 (.A1( u0_uk_K_r13_25 ) , .A2( u0_uk_n251 ) , .ZN( u0_uk_n924 ) );
  OAI22_X1 u0_uk_U650 (.ZN( u0_K14_43 ) , .B1( u0_uk_n203 ) , .A2( u0_uk_n56 ) , .B2( u0_uk_n59 ) , .A1( u0_uk_n60 ) );
  OAI21_X1 u0_uk_U662 (.ZN( u0_K14_45 ) , .B1( u0_uk_n217 ) , .B2( u0_uk_n58 ) , .A( u0_uk_n929 ) );
  NAND2_X1 u0_uk_U663 (.A1( u0_uk_K_r12_16 ) , .A2( u0_uk_n252 ) , .ZN( u0_uk_n929 ) );
  OAI22_X1 u0_uk_U679 (.ZN( u0_K15_7 ) , .A1( u0_uk_n155 ) , .B1( u0_uk_n17 ) , .A2( u0_uk_n19 ) , .B2( u0_uk_n35 ) );
  OAI22_X1 u0_uk_U842 (.ZN( u0_K15_6 ) , .B1( u0_uk_n17 ) , .A1( u0_uk_n187 ) , .B2( u0_uk_n24 ) , .A2( u0_uk_n6 ) );
  OAI22_X1 u0_uk_U850 (.ZN( u0_K15_3 ) , .A1( u0_uk_n155 ) , .B1( u0_uk_n17 ) , .A2( u0_uk_n20 ) , .B2( u0_uk_n36 ) );
  OAI21_X1 u0_uk_U856 (.ZN( u0_K14_3 ) , .B1( u0_uk_n17 ) , .B2( u0_uk_n46 ) , .A( u0_uk_n932 ) );
  NAND2_X1 u0_uk_U857 (.A1( u0_uk_K_r12_47 ) , .A2( u0_uk_n63 ) , .ZN( u0_uk_n932 ) );
  OAI22_X1 u0_uk_U889 (.ZN( u0_K6_45 ) , .A1( u0_uk_n213 ) , .A2( u0_uk_n429 ) , .B2( u0_uk_n434 ) , .B1( u0_uk_n60 ) );
  OAI22_X1 u0_uk_U893 (.ZN( u0_K14_6 ) , .A1( u0_uk_n230 ) , .B2( u0_uk_n78 ) , .A2( u0_uk_n85 ) , .B1( u0_uk_n92 ) );
  OAI22_X1 u0_uk_U902 (.ZN( u0_K15_13 ) , .B2( u0_uk_n16 ) , .A1( u0_uk_n230 ) , .A2( u0_uk_n44 ) , .B1( u0_uk_n92 ) );
  OAI22_X1 u0_uk_U947 (.ZN( u0_K14_47 ) , .A1( u0_uk_n17 ) , .B1( u0_uk_n231 ) , .A2( u0_uk_n58 ) , .B2( u0_uk_n68 ) );
  OAI22_X1 u0_uk_U95 (.ZN( u0_K15_5 ) , .B1( u0_uk_n220 ) , .A2( u0_uk_n26 ) , .B2( u0_uk_n29 ) , .A1( u0_uk_n94 ) );
  OAI22_X1 u0_uk_U951 (.ZN( u0_K6_46 ) , .A1( u0_uk_n109 ) , .B1( u0_uk_n203 ) , .B2( u0_uk_n417 ) , .A2( u0_uk_n445 ) );
  OAI21_X1 u0_uk_U96 (.ZN( u0_K14_5 ) , .B1( u0_uk_n203 ) , .B2( u0_uk_n62 ) , .A( u0_uk_n927 ) );
  OAI22_X1 u0_uk_U966 (.ZN( u0_K14_38 ) , .A1( u0_uk_n141 ) , .B1( u0_uk_n250 ) , .B2( u0_uk_n65 ) , .A2( u0_uk_n81 ) );
  NAND2_X1 u0_uk_U97 (.A1( u0_uk_K_r12_10 ) , .A2( u0_uk_n251 ) , .ZN( u0_uk_n927 ) );
  OAI22_X1 u0_uk_U977 (.ZN( u0_K6_43 ) , .A1( u0_uk_n109 ) , .B1( u0_uk_n214 ) , .A2( u0_uk_n411 ) , .B2( u0_uk_n450 ) );
  XOR2_X1 u1_U101 (.B( u1_L12_26 ) , .Z( u1_N441 ) , .A( u1_out13_26 ) );
  XOR2_X1 u1_U108 (.B( u1_L12_20 ) , .Z( u1_N435 ) , .A( u1_out13_20 ) );
  XOR2_X1 u1_U119 (.B( u1_L12_10 ) , .Z( u1_N425 ) , .A( u1_out13_10 ) );
  XOR2_X1 u1_U12 (.B( u1_L1_27 ) , .Z( u1_N90 ) , .A( u1_out2_27 ) );
  XOR2_X1 u1_U129 (.B( u1_L12_1 ) , .Z( u1_N416 ) , .A( u1_out13_1 ) );
  XOR2_X1 u1_U174 (.B( u1_L10_25 ) , .Z( u1_N376 ) , .A( u1_out11_25 ) );
  XOR2_X1 u1_U18 (.B( u1_L1_22 ) , .Z( u1_N85 ) , .A( u1_out2_22 ) );
  XOR2_X1 u1_U186 (.B( u1_L10_14 ) , .Z( u1_N365 ) , .A( u1_out11_14 ) );
  XOR2_X1 u1_U19 (.B( u1_L1_21 ) , .Z( u1_N84 ) , .A( u1_out2_21 ) );
  XOR2_X1 u1_U193 (.B( u1_L10_8 ) , .Z( u1_N359 ) , .A( u1_out11_8 ) );
  XOR2_X1 u1_U198 (.B( u1_L10_3 ) , .Z( u1_N354 ) , .A( u1_out11_3 ) );
  XOR2_X1 u1_U243 (.B( u1_L8_26 ) , .Z( u1_N313 ) , .A( u1_out9_26 ) );
  XOR2_X1 u1_U250 (.B( u1_L8_20 ) , .Z( u1_N307 ) , .A( u1_out9_20 ) );
  XOR2_X1 u1_U26 (.B( u1_L1_15 ) , .Z( u1_N78 ) , .A( u1_out2_15 ) );
  XOR2_X1 u1_U262 (.B( u1_L8_10 ) , .Z( u1_N297 ) , .A( u1_out9_10 ) );
  XOR2_X1 u1_U272 (.B( u1_L8_1 ) , .Z( u1_N288 ) , .A( u1_out9_1 ) );
  XOR2_X1 u1_U29 (.B( u1_L1_12 ) , .Z( u1_N75 ) , .A( u1_out2_12 ) );
  XOR2_X1 u1_U315 (.B( u1_L6_26 ) , .Z( u1_N249 ) , .A( u1_out7_26 ) );
  XOR2_X1 u1_U321 (.B( u1_L6_20 ) , .Z( u1_N243 ) , .A( u1_out7_20 ) );
  XOR2_X1 u1_U332 (.B( u1_L6_10 ) , .Z( u1_N233 ) , .A( u1_out7_10 ) );
  XOR2_X1 u1_U34 (.B( u1_L1_7 ) , .Z( u1_N70 ) , .A( u1_out2_7 ) );
  XOR2_X1 u1_U342 (.B( u1_L6_1 ) , .Z( u1_N224 ) , .A( u1_out7_1 ) );
  XOR2_X1 u1_U37 (.B( u1_L1_5 ) , .Z( u1_N68 ) , .A( u1_out2_5 ) );
  XOR2_X1 u1_U4 (.B( u1_L2_3 ) , .Z( u1_N98 ) , .A( u1_out3_3 ) );
  XOR2_X1 u1_U421 (.B( u1_L3_26 ) , .Z( u1_N153 ) , .A( u1_out4_26 ) );
  XOR2_X1 u1_U428 (.B( u1_L3_20 ) , .Z( u1_N147 ) , .A( u1_out4_20 ) );
  XOR2_X1 u1_U439 (.B( u1_L3_10 ) , .Z( u1_N137 ) , .A( u1_out4_10 ) );
  XOR2_X1 u1_U449 (.B( u1_L3_1 ) , .Z( u1_N128 ) , .A( u1_out4_1 ) );
  XOR2_X1 u1_U457 (.B( u1_L2_25 ) , .Z( u1_N120 ) , .A( u1_out3_25 ) );
  XOR2_X1 u1_U470 (.B( u1_L2_14 ) , .Z( u1_N109 ) , .A( u1_out3_14 ) );
  XOR2_X1 u1_U476 (.B( u1_L2_8 ) , .Z( u1_N103 ) , .A( u1_out3_8 ) );
  XOR2_X1 u1_U7 (.B( u1_L1_32 ) , .Z( u1_N95 ) , .A( u1_out2_32 ) );
  XOR2_X1 u1_u11_U26 (.B( u1_K12_30 ) , .A( u1_R10_21 ) , .Z( u1_u11_X_30 ) );
  XOR2_X1 u1_u11_U28 (.B( u1_K12_29 ) , .A( u1_R10_20 ) , .Z( u1_u11_X_29 ) );
  XOR2_X1 u1_u11_U29 (.B( u1_K12_28 ) , .A( u1_R10_19 ) , .Z( u1_u11_X_28 ) );
  XOR2_X1 u1_u11_U30 (.B( u1_K12_27 ) , .A( u1_R10_18 ) , .Z( u1_u11_X_27 ) );
  XOR2_X1 u1_u11_U31 (.B( u1_K12_26 ) , .A( u1_R10_17 ) , .Z( u1_u11_X_26 ) );
  XOR2_X1 u1_u11_U32 (.B( u1_K12_25 ) , .A( u1_R10_16 ) , .Z( u1_u11_X_25 ) );
  OAI22_X1 u1_u11_u4_U10 (.B2( u1_u11_u4_n135 ) , .ZN( u1_u11_u4_n137 ) , .B1( u1_u11_u4_n153 ) , .A1( u1_u11_u4_n155 ) , .A2( u1_u11_u4_n171 ) );
  AND3_X1 u1_u11_u4_U11 (.A2( u1_u11_u4_n134 ) , .ZN( u1_u11_u4_n135 ) , .A3( u1_u11_u4_n145 ) , .A1( u1_u11_u4_n157 ) );
  NAND2_X1 u1_u11_u4_U12 (.ZN( u1_u11_u4_n132 ) , .A2( u1_u11_u4_n170 ) , .A1( u1_u11_u4_n173 ) );
  AOI21_X1 u1_u11_u4_U13 (.B2( u1_u11_u4_n160 ) , .B1( u1_u11_u4_n161 ) , .ZN( u1_u11_u4_n162 ) , .A( u1_u11_u4_n170 ) );
  AOI21_X1 u1_u11_u4_U14 (.ZN( u1_u11_u4_n107 ) , .B2( u1_u11_u4_n143 ) , .A( u1_u11_u4_n174 ) , .B1( u1_u11_u4_n184 ) );
  AOI21_X1 u1_u11_u4_U15 (.B2( u1_u11_u4_n158 ) , .B1( u1_u11_u4_n159 ) , .ZN( u1_u11_u4_n163 ) , .A( u1_u11_u4_n174 ) );
  AOI21_X1 u1_u11_u4_U16 (.A( u1_u11_u4_n153 ) , .B2( u1_u11_u4_n154 ) , .B1( u1_u11_u4_n155 ) , .ZN( u1_u11_u4_n165 ) );
  AOI21_X1 u1_u11_u4_U17 (.A( u1_u11_u4_n156 ) , .B2( u1_u11_u4_n157 ) , .ZN( u1_u11_u4_n164 ) , .B1( u1_u11_u4_n184 ) );
  INV_X1 u1_u11_u4_U18 (.A( u1_u11_u4_n138 ) , .ZN( u1_u11_u4_n170 ) );
  AND2_X1 u1_u11_u4_U19 (.A2( u1_u11_u4_n120 ) , .ZN( u1_u11_u4_n155 ) , .A1( u1_u11_u4_n160 ) );
  INV_X1 u1_u11_u4_U20 (.A( u1_u11_u4_n156 ) , .ZN( u1_u11_u4_n175 ) );
  NAND2_X1 u1_u11_u4_U21 (.A2( u1_u11_u4_n118 ) , .ZN( u1_u11_u4_n131 ) , .A1( u1_u11_u4_n147 ) );
  NAND2_X1 u1_u11_u4_U22 (.A1( u1_u11_u4_n119 ) , .A2( u1_u11_u4_n120 ) , .ZN( u1_u11_u4_n130 ) );
  NAND2_X1 u1_u11_u4_U23 (.ZN( u1_u11_u4_n117 ) , .A2( u1_u11_u4_n118 ) , .A1( u1_u11_u4_n148 ) );
  NAND2_X1 u1_u11_u4_U24 (.ZN( u1_u11_u4_n129 ) , .A1( u1_u11_u4_n134 ) , .A2( u1_u11_u4_n148 ) );
  AND3_X1 u1_u11_u4_U25 (.A1( u1_u11_u4_n119 ) , .A2( u1_u11_u4_n143 ) , .A3( u1_u11_u4_n154 ) , .ZN( u1_u11_u4_n161 ) );
  AND2_X1 u1_u11_u4_U26 (.A1( u1_u11_u4_n145 ) , .A2( u1_u11_u4_n147 ) , .ZN( u1_u11_u4_n159 ) );
  OR3_X1 u1_u11_u4_U27 (.A3( u1_u11_u4_n114 ) , .A2( u1_u11_u4_n115 ) , .A1( u1_u11_u4_n116 ) , .ZN( u1_u11_u4_n136 ) );
  AOI21_X1 u1_u11_u4_U28 (.A( u1_u11_u4_n113 ) , .ZN( u1_u11_u4_n116 ) , .B2( u1_u11_u4_n173 ) , .B1( u1_u11_u4_n174 ) );
  AOI21_X1 u1_u11_u4_U29 (.ZN( u1_u11_u4_n115 ) , .B2( u1_u11_u4_n145 ) , .B1( u1_u11_u4_n146 ) , .A( u1_u11_u4_n156 ) );
  NOR2_X1 u1_u11_u4_U3 (.ZN( u1_u11_u4_n121 ) , .A1( u1_u11_u4_n181 ) , .A2( u1_u11_u4_n182 ) );
  OAI22_X1 u1_u11_u4_U30 (.ZN( u1_u11_u4_n114 ) , .A2( u1_u11_u4_n121 ) , .B1( u1_u11_u4_n160 ) , .B2( u1_u11_u4_n170 ) , .A1( u1_u11_u4_n171 ) );
  INV_X1 u1_u11_u4_U31 (.A( u1_u11_u4_n158 ) , .ZN( u1_u11_u4_n182 ) );
  INV_X1 u1_u11_u4_U32 (.ZN( u1_u11_u4_n181 ) , .A( u1_u11_u4_n96 ) );
  INV_X1 u1_u11_u4_U33 (.A( u1_u11_u4_n144 ) , .ZN( u1_u11_u4_n179 ) );
  INV_X1 u1_u11_u4_U34 (.A( u1_u11_u4_n157 ) , .ZN( u1_u11_u4_n178 ) );
  NAND2_X1 u1_u11_u4_U35 (.A2( u1_u11_u4_n154 ) , .A1( u1_u11_u4_n96 ) , .ZN( u1_u11_u4_n97 ) );
  INV_X1 u1_u11_u4_U36 (.ZN( u1_u11_u4_n186 ) , .A( u1_u11_u4_n95 ) );
  OAI221_X1 u1_u11_u4_U37 (.C1( u1_u11_u4_n134 ) , .B1( u1_u11_u4_n158 ) , .B2( u1_u11_u4_n171 ) , .C2( u1_u11_u4_n173 ) , .A( u1_u11_u4_n94 ) , .ZN( u1_u11_u4_n95 ) );
  AOI222_X1 u1_u11_u4_U38 (.B2( u1_u11_u4_n132 ) , .A1( u1_u11_u4_n138 ) , .C2( u1_u11_u4_n175 ) , .A2( u1_u11_u4_n179 ) , .C1( u1_u11_u4_n181 ) , .B1( u1_u11_u4_n185 ) , .ZN( u1_u11_u4_n94 ) );
  INV_X1 u1_u11_u4_U39 (.A( u1_u11_u4_n113 ) , .ZN( u1_u11_u4_n185 ) );
  INV_X1 u1_u11_u4_U4 (.A( u1_u11_u4_n117 ) , .ZN( u1_u11_u4_n184 ) );
  INV_X1 u1_u11_u4_U40 (.A( u1_u11_u4_n143 ) , .ZN( u1_u11_u4_n183 ) );
  NOR2_X1 u1_u11_u4_U41 (.ZN( u1_u11_u4_n138 ) , .A1( u1_u11_u4_n168 ) , .A2( u1_u11_u4_n169 ) );
  NOR2_X1 u1_u11_u4_U42 (.A1( u1_u11_u4_n150 ) , .A2( u1_u11_u4_n152 ) , .ZN( u1_u11_u4_n153 ) );
  NOR2_X1 u1_u11_u4_U43 (.A2( u1_u11_u4_n128 ) , .A1( u1_u11_u4_n138 ) , .ZN( u1_u11_u4_n156 ) );
  AOI22_X1 u1_u11_u4_U44 (.B2( u1_u11_u4_n122 ) , .A1( u1_u11_u4_n123 ) , .ZN( u1_u11_u4_n124 ) , .B1( u1_u11_u4_n128 ) , .A2( u1_u11_u4_n172 ) );
  INV_X1 u1_u11_u4_U45 (.A( u1_u11_u4_n153 ) , .ZN( u1_u11_u4_n172 ) );
  NAND2_X1 u1_u11_u4_U46 (.A2( u1_u11_u4_n120 ) , .ZN( u1_u11_u4_n123 ) , .A1( u1_u11_u4_n161 ) );
  AOI22_X1 u1_u11_u4_U47 (.B2( u1_u11_u4_n132 ) , .A2( u1_u11_u4_n133 ) , .ZN( u1_u11_u4_n140 ) , .A1( u1_u11_u4_n150 ) , .B1( u1_u11_u4_n179 ) );
  NAND2_X1 u1_u11_u4_U48 (.ZN( u1_u11_u4_n133 ) , .A2( u1_u11_u4_n146 ) , .A1( u1_u11_u4_n154 ) );
  NAND2_X1 u1_u11_u4_U49 (.A1( u1_u11_u4_n103 ) , .ZN( u1_u11_u4_n154 ) , .A2( u1_u11_u4_n98 ) );
  NOR4_X1 u1_u11_u4_U5 (.A4( u1_u11_u4_n106 ) , .A3( u1_u11_u4_n107 ) , .A2( u1_u11_u4_n108 ) , .A1( u1_u11_u4_n109 ) , .ZN( u1_u11_u4_n110 ) );
  NAND2_X1 u1_u11_u4_U50 (.A1( u1_u11_u4_n101 ) , .ZN( u1_u11_u4_n158 ) , .A2( u1_u11_u4_n99 ) );
  AOI21_X1 u1_u11_u4_U51 (.ZN( u1_u11_u4_n127 ) , .A( u1_u11_u4_n136 ) , .B2( u1_u11_u4_n150 ) , .B1( u1_u11_u4_n180 ) );
  INV_X1 u1_u11_u4_U52 (.A( u1_u11_u4_n160 ) , .ZN( u1_u11_u4_n180 ) );
  NAND2_X1 u1_u11_u4_U53 (.A2( u1_u11_u4_n104 ) , .A1( u1_u11_u4_n105 ) , .ZN( u1_u11_u4_n146 ) );
  NAND2_X1 u1_u11_u4_U54 (.A2( u1_u11_u4_n101 ) , .A1( u1_u11_u4_n102 ) , .ZN( u1_u11_u4_n160 ) );
  NAND2_X1 u1_u11_u4_U55 (.ZN( u1_u11_u4_n134 ) , .A1( u1_u11_u4_n98 ) , .A2( u1_u11_u4_n99 ) );
  NAND2_X1 u1_u11_u4_U56 (.A1( u1_u11_u4_n103 ) , .A2( u1_u11_u4_n104 ) , .ZN( u1_u11_u4_n143 ) );
  NAND2_X1 u1_u11_u4_U57 (.A2( u1_u11_u4_n105 ) , .ZN( u1_u11_u4_n145 ) , .A1( u1_u11_u4_n98 ) );
  NAND2_X1 u1_u11_u4_U58 (.A1( u1_u11_u4_n100 ) , .A2( u1_u11_u4_n105 ) , .ZN( u1_u11_u4_n120 ) );
  NAND2_X1 u1_u11_u4_U59 (.A1( u1_u11_u4_n102 ) , .A2( u1_u11_u4_n104 ) , .ZN( u1_u11_u4_n148 ) );
  AOI21_X1 u1_u11_u4_U6 (.ZN( u1_u11_u4_n106 ) , .B2( u1_u11_u4_n146 ) , .B1( u1_u11_u4_n158 ) , .A( u1_u11_u4_n170 ) );
  NAND2_X1 u1_u11_u4_U60 (.A2( u1_u11_u4_n100 ) , .A1( u1_u11_u4_n103 ) , .ZN( u1_u11_u4_n157 ) );
  INV_X1 u1_u11_u4_U61 (.A( u1_u11_u4_n150 ) , .ZN( u1_u11_u4_n173 ) );
  INV_X1 u1_u11_u4_U62 (.A( u1_u11_u4_n152 ) , .ZN( u1_u11_u4_n171 ) );
  NAND2_X1 u1_u11_u4_U63 (.A1( u1_u11_u4_n100 ) , .ZN( u1_u11_u4_n118 ) , .A2( u1_u11_u4_n99 ) );
  NAND2_X1 u1_u11_u4_U64 (.A2( u1_u11_u4_n100 ) , .A1( u1_u11_u4_n102 ) , .ZN( u1_u11_u4_n144 ) );
  NAND2_X1 u1_u11_u4_U65 (.A2( u1_u11_u4_n101 ) , .A1( u1_u11_u4_n105 ) , .ZN( u1_u11_u4_n96 ) );
  INV_X1 u1_u11_u4_U66 (.A( u1_u11_u4_n128 ) , .ZN( u1_u11_u4_n174 ) );
  NAND2_X1 u1_u11_u4_U67 (.A2( u1_u11_u4_n102 ) , .ZN( u1_u11_u4_n119 ) , .A1( u1_u11_u4_n98 ) );
  NAND2_X1 u1_u11_u4_U68 (.A2( u1_u11_u4_n101 ) , .A1( u1_u11_u4_n103 ) , .ZN( u1_u11_u4_n147 ) );
  NAND2_X1 u1_u11_u4_U69 (.A2( u1_u11_u4_n104 ) , .ZN( u1_u11_u4_n113 ) , .A1( u1_u11_u4_n99 ) );
  AOI21_X1 u1_u11_u4_U7 (.ZN( u1_u11_u4_n108 ) , .B2( u1_u11_u4_n134 ) , .B1( u1_u11_u4_n155 ) , .A( u1_u11_u4_n156 ) );
  NOR2_X1 u1_u11_u4_U70 (.A2( u1_u11_X_28 ) , .ZN( u1_u11_u4_n150 ) , .A1( u1_u11_u4_n168 ) );
  NOR2_X1 u1_u11_u4_U71 (.A2( u1_u11_X_29 ) , .ZN( u1_u11_u4_n152 ) , .A1( u1_u11_u4_n169 ) );
  NOR2_X1 u1_u11_u4_U72 (.A2( u1_u11_X_26 ) , .ZN( u1_u11_u4_n100 ) , .A1( u1_u11_u4_n177 ) );
  NOR2_X1 u1_u11_u4_U73 (.A2( u1_u11_X_30 ) , .ZN( u1_u11_u4_n105 ) , .A1( u1_u11_u4_n176 ) );
  NOR2_X1 u1_u11_u4_U74 (.A2( u1_u11_X_28 ) , .A1( u1_u11_X_29 ) , .ZN( u1_u11_u4_n128 ) );
  NOR2_X1 u1_u11_u4_U75 (.A2( u1_u11_X_25 ) , .A1( u1_u11_X_26 ) , .ZN( u1_u11_u4_n98 ) );
  NOR2_X1 u1_u11_u4_U76 (.A2( u1_u11_X_27 ) , .A1( u1_u11_X_30 ) , .ZN( u1_u11_u4_n102 ) );
  AND2_X1 u1_u11_u4_U77 (.A2( u1_u11_X_25 ) , .A1( u1_u11_X_26 ) , .ZN( u1_u11_u4_n104 ) );
  AND2_X1 u1_u11_u4_U78 (.A1( u1_u11_X_30 ) , .A2( u1_u11_u4_n176 ) , .ZN( u1_u11_u4_n99 ) );
  AND2_X1 u1_u11_u4_U79 (.A1( u1_u11_X_26 ) , .ZN( u1_u11_u4_n101 ) , .A2( u1_u11_u4_n177 ) );
  AOI21_X1 u1_u11_u4_U8 (.ZN( u1_u11_u4_n109 ) , .A( u1_u11_u4_n153 ) , .B1( u1_u11_u4_n159 ) , .B2( u1_u11_u4_n184 ) );
  AND2_X1 u1_u11_u4_U80 (.A1( u1_u11_X_27 ) , .A2( u1_u11_X_30 ) , .ZN( u1_u11_u4_n103 ) );
  INV_X1 u1_u11_u4_U81 (.A( u1_u11_X_28 ) , .ZN( u1_u11_u4_n169 ) );
  INV_X1 u1_u11_u4_U82 (.A( u1_u11_X_29 ) , .ZN( u1_u11_u4_n168 ) );
  INV_X1 u1_u11_u4_U83 (.A( u1_u11_X_25 ) , .ZN( u1_u11_u4_n177 ) );
  INV_X1 u1_u11_u4_U84 (.A( u1_u11_X_27 ) , .ZN( u1_u11_u4_n176 ) );
  NAND4_X1 u1_u11_u4_U85 (.ZN( u1_out11_25 ) , .A4( u1_u11_u4_n139 ) , .A3( u1_u11_u4_n140 ) , .A2( u1_u11_u4_n141 ) , .A1( u1_u11_u4_n142 ) );
  OAI21_X1 u1_u11_u4_U86 (.A( u1_u11_u4_n128 ) , .B2( u1_u11_u4_n129 ) , .B1( u1_u11_u4_n130 ) , .ZN( u1_u11_u4_n142 ) );
  OAI21_X1 u1_u11_u4_U87 (.B2( u1_u11_u4_n131 ) , .ZN( u1_u11_u4_n141 ) , .A( u1_u11_u4_n175 ) , .B1( u1_u11_u4_n183 ) );
  NAND4_X1 u1_u11_u4_U88 (.ZN( u1_out11_14 ) , .A4( u1_u11_u4_n124 ) , .A3( u1_u11_u4_n125 ) , .A2( u1_u11_u4_n126 ) , .A1( u1_u11_u4_n127 ) );
  AOI22_X1 u1_u11_u4_U89 (.B2( u1_u11_u4_n117 ) , .ZN( u1_u11_u4_n126 ) , .A1( u1_u11_u4_n129 ) , .B1( u1_u11_u4_n152 ) , .A2( u1_u11_u4_n175 ) );
  AOI211_X1 u1_u11_u4_U9 (.B( u1_u11_u4_n136 ) , .A( u1_u11_u4_n137 ) , .C2( u1_u11_u4_n138 ) , .ZN( u1_u11_u4_n139 ) , .C1( u1_u11_u4_n182 ) );
  AOI22_X1 u1_u11_u4_U90 (.ZN( u1_u11_u4_n125 ) , .B2( u1_u11_u4_n131 ) , .A2( u1_u11_u4_n132 ) , .B1( u1_u11_u4_n138 ) , .A1( u1_u11_u4_n178 ) );
  NAND4_X1 u1_u11_u4_U91 (.ZN( u1_out11_8 ) , .A4( u1_u11_u4_n110 ) , .A3( u1_u11_u4_n111 ) , .A2( u1_u11_u4_n112 ) , .A1( u1_u11_u4_n186 ) );
  NAND2_X1 u1_u11_u4_U92 (.ZN( u1_u11_u4_n112 ) , .A2( u1_u11_u4_n130 ) , .A1( u1_u11_u4_n150 ) );
  AOI22_X1 u1_u11_u4_U93 (.ZN( u1_u11_u4_n111 ) , .B2( u1_u11_u4_n132 ) , .A1( u1_u11_u4_n152 ) , .B1( u1_u11_u4_n178 ) , .A2( u1_u11_u4_n97 ) );
  AOI22_X1 u1_u11_u4_U94 (.B2( u1_u11_u4_n149 ) , .B1( u1_u11_u4_n150 ) , .A2( u1_u11_u4_n151 ) , .A1( u1_u11_u4_n152 ) , .ZN( u1_u11_u4_n167 ) );
  NOR4_X1 u1_u11_u4_U95 (.A4( u1_u11_u4_n162 ) , .A3( u1_u11_u4_n163 ) , .A2( u1_u11_u4_n164 ) , .A1( u1_u11_u4_n165 ) , .ZN( u1_u11_u4_n166 ) );
  NAND3_X1 u1_u11_u4_U96 (.ZN( u1_out11_3 ) , .A3( u1_u11_u4_n166 ) , .A1( u1_u11_u4_n167 ) , .A2( u1_u11_u4_n186 ) );
  NAND3_X1 u1_u11_u4_U97 (.A3( u1_u11_u4_n146 ) , .A2( u1_u11_u4_n147 ) , .A1( u1_u11_u4_n148 ) , .ZN( u1_u11_u4_n149 ) );
  NAND3_X1 u1_u11_u4_U98 (.A3( u1_u11_u4_n143 ) , .A2( u1_u11_u4_n144 ) , .A1( u1_u11_u4_n145 ) , .ZN( u1_u11_u4_n151 ) );
  NAND3_X1 u1_u11_u4_U99 (.A3( u1_u11_u4_n121 ) , .ZN( u1_u11_u4_n122 ) , .A2( u1_u11_u4_n144 ) , .A1( u1_u11_u4_n154 ) );
  XOR2_X1 u1_u13_U33 (.B( u1_K14_24 ) , .A( u1_R12_17 ) , .Z( u1_u13_X_24 ) );
  XOR2_X1 u1_u13_U34 (.B( u1_K14_23 ) , .A( u1_R12_16 ) , .Z( u1_u13_X_23 ) );
  XOR2_X1 u1_u13_U35 (.B( u1_K14_22 ) , .A( u1_R12_15 ) , .Z( u1_u13_X_22 ) );
  XOR2_X1 u1_u13_U36 (.B( u1_K14_21 ) , .A( u1_R12_14 ) , .Z( u1_u13_X_21 ) );
  XOR2_X1 u1_u13_U37 (.B( u1_K14_20 ) , .A( u1_R12_13 ) , .Z( u1_u13_X_20 ) );
  XOR2_X1 u1_u13_U39 (.B( u1_K14_19 ) , .A( u1_R12_12 ) , .Z( u1_u13_X_19 ) );
  OAI22_X1 u1_u13_u3_U10 (.B1( u1_u13_u3_n113 ) , .A2( u1_u13_u3_n135 ) , .A1( u1_u13_u3_n150 ) , .B2( u1_u13_u3_n164 ) , .ZN( u1_u13_u3_n98 ) );
  OAI211_X1 u1_u13_u3_U11 (.B( u1_u13_u3_n106 ) , .ZN( u1_u13_u3_n119 ) , .C2( u1_u13_u3_n128 ) , .C1( u1_u13_u3_n167 ) , .A( u1_u13_u3_n181 ) );
  AOI221_X1 u1_u13_u3_U12 (.C1( u1_u13_u3_n105 ) , .ZN( u1_u13_u3_n106 ) , .A( u1_u13_u3_n131 ) , .B2( u1_u13_u3_n132 ) , .C2( u1_u13_u3_n133 ) , .B1( u1_u13_u3_n169 ) );
  INV_X1 u1_u13_u3_U13 (.ZN( u1_u13_u3_n181 ) , .A( u1_u13_u3_n98 ) );
  NAND2_X1 u1_u13_u3_U14 (.ZN( u1_u13_u3_n105 ) , .A2( u1_u13_u3_n130 ) , .A1( u1_u13_u3_n155 ) );
  AOI22_X1 u1_u13_u3_U15 (.B1( u1_u13_u3_n115 ) , .A2( u1_u13_u3_n116 ) , .ZN( u1_u13_u3_n123 ) , .B2( u1_u13_u3_n133 ) , .A1( u1_u13_u3_n169 ) );
  NAND2_X1 u1_u13_u3_U16 (.ZN( u1_u13_u3_n116 ) , .A2( u1_u13_u3_n151 ) , .A1( u1_u13_u3_n182 ) );
  NOR2_X1 u1_u13_u3_U17 (.ZN( u1_u13_u3_n126 ) , .A2( u1_u13_u3_n150 ) , .A1( u1_u13_u3_n164 ) );
  AOI21_X1 u1_u13_u3_U18 (.ZN( u1_u13_u3_n112 ) , .B2( u1_u13_u3_n146 ) , .B1( u1_u13_u3_n155 ) , .A( u1_u13_u3_n167 ) );
  NAND2_X1 u1_u13_u3_U19 (.A1( u1_u13_u3_n135 ) , .ZN( u1_u13_u3_n142 ) , .A2( u1_u13_u3_n164 ) );
  NAND2_X1 u1_u13_u3_U20 (.ZN( u1_u13_u3_n132 ) , .A2( u1_u13_u3_n152 ) , .A1( u1_u13_u3_n156 ) );
  AND2_X1 u1_u13_u3_U21 (.A2( u1_u13_u3_n113 ) , .A1( u1_u13_u3_n114 ) , .ZN( u1_u13_u3_n151 ) );
  INV_X1 u1_u13_u3_U22 (.A( u1_u13_u3_n133 ) , .ZN( u1_u13_u3_n165 ) );
  INV_X1 u1_u13_u3_U23 (.A( u1_u13_u3_n135 ) , .ZN( u1_u13_u3_n170 ) );
  NAND2_X1 u1_u13_u3_U24 (.A1( u1_u13_u3_n107 ) , .A2( u1_u13_u3_n108 ) , .ZN( u1_u13_u3_n140 ) );
  NAND2_X1 u1_u13_u3_U25 (.ZN( u1_u13_u3_n117 ) , .A1( u1_u13_u3_n124 ) , .A2( u1_u13_u3_n148 ) );
  NAND2_X1 u1_u13_u3_U26 (.ZN( u1_u13_u3_n143 ) , .A1( u1_u13_u3_n165 ) , .A2( u1_u13_u3_n167 ) );
  INV_X1 u1_u13_u3_U27 (.A( u1_u13_u3_n130 ) , .ZN( u1_u13_u3_n177 ) );
  INV_X1 u1_u13_u3_U28 (.A( u1_u13_u3_n128 ) , .ZN( u1_u13_u3_n176 ) );
  INV_X1 u1_u13_u3_U29 (.A( u1_u13_u3_n155 ) , .ZN( u1_u13_u3_n174 ) );
  INV_X1 u1_u13_u3_U3 (.A( u1_u13_u3_n129 ) , .ZN( u1_u13_u3_n183 ) );
  INV_X1 u1_u13_u3_U30 (.A( u1_u13_u3_n139 ) , .ZN( u1_u13_u3_n185 ) );
  NOR2_X1 u1_u13_u3_U31 (.ZN( u1_u13_u3_n135 ) , .A2( u1_u13_u3_n141 ) , .A1( u1_u13_u3_n169 ) );
  OAI222_X1 u1_u13_u3_U32 (.C2( u1_u13_u3_n107 ) , .A2( u1_u13_u3_n108 ) , .B1( u1_u13_u3_n135 ) , .ZN( u1_u13_u3_n138 ) , .B2( u1_u13_u3_n146 ) , .C1( u1_u13_u3_n154 ) , .A1( u1_u13_u3_n164 ) );
  NOR4_X1 u1_u13_u3_U33 (.A4( u1_u13_u3_n157 ) , .A3( u1_u13_u3_n158 ) , .A2( u1_u13_u3_n159 ) , .A1( u1_u13_u3_n160 ) , .ZN( u1_u13_u3_n161 ) );
  AOI21_X1 u1_u13_u3_U34 (.B2( u1_u13_u3_n152 ) , .B1( u1_u13_u3_n153 ) , .ZN( u1_u13_u3_n158 ) , .A( u1_u13_u3_n164 ) );
  AOI21_X1 u1_u13_u3_U35 (.A( u1_u13_u3_n154 ) , .B2( u1_u13_u3_n155 ) , .B1( u1_u13_u3_n156 ) , .ZN( u1_u13_u3_n157 ) );
  AOI21_X1 u1_u13_u3_U36 (.A( u1_u13_u3_n149 ) , .B2( u1_u13_u3_n150 ) , .B1( u1_u13_u3_n151 ) , .ZN( u1_u13_u3_n159 ) );
  AOI211_X1 u1_u13_u3_U37 (.ZN( u1_u13_u3_n109 ) , .A( u1_u13_u3_n119 ) , .C2( u1_u13_u3_n129 ) , .B( u1_u13_u3_n138 ) , .C1( u1_u13_u3_n141 ) );
  AOI211_X1 u1_u13_u3_U38 (.B( u1_u13_u3_n119 ) , .A( u1_u13_u3_n120 ) , .C2( u1_u13_u3_n121 ) , .ZN( u1_u13_u3_n122 ) , .C1( u1_u13_u3_n179 ) );
  INV_X1 u1_u13_u3_U39 (.A( u1_u13_u3_n156 ) , .ZN( u1_u13_u3_n179 ) );
  INV_X1 u1_u13_u3_U4 (.A( u1_u13_u3_n140 ) , .ZN( u1_u13_u3_n182 ) );
  OAI22_X1 u1_u13_u3_U40 (.B1( u1_u13_u3_n118 ) , .ZN( u1_u13_u3_n120 ) , .A1( u1_u13_u3_n135 ) , .B2( u1_u13_u3_n154 ) , .A2( u1_u13_u3_n178 ) );
  AND3_X1 u1_u13_u3_U41 (.ZN( u1_u13_u3_n118 ) , .A2( u1_u13_u3_n124 ) , .A1( u1_u13_u3_n144 ) , .A3( u1_u13_u3_n152 ) );
  INV_X1 u1_u13_u3_U42 (.A( u1_u13_u3_n121 ) , .ZN( u1_u13_u3_n164 ) );
  NAND2_X1 u1_u13_u3_U43 (.ZN( u1_u13_u3_n133 ) , .A1( u1_u13_u3_n154 ) , .A2( u1_u13_u3_n164 ) );
  OAI211_X1 u1_u13_u3_U44 (.B( u1_u13_u3_n127 ) , .ZN( u1_u13_u3_n139 ) , .C1( u1_u13_u3_n150 ) , .C2( u1_u13_u3_n154 ) , .A( u1_u13_u3_n184 ) );
  INV_X1 u1_u13_u3_U45 (.A( u1_u13_u3_n125 ) , .ZN( u1_u13_u3_n184 ) );
  AOI221_X1 u1_u13_u3_U46 (.A( u1_u13_u3_n126 ) , .ZN( u1_u13_u3_n127 ) , .C2( u1_u13_u3_n132 ) , .C1( u1_u13_u3_n169 ) , .B2( u1_u13_u3_n170 ) , .B1( u1_u13_u3_n174 ) );
  OAI22_X1 u1_u13_u3_U47 (.A1( u1_u13_u3_n124 ) , .ZN( u1_u13_u3_n125 ) , .B2( u1_u13_u3_n145 ) , .A2( u1_u13_u3_n165 ) , .B1( u1_u13_u3_n167 ) );
  NOR2_X1 u1_u13_u3_U48 (.A1( u1_u13_u3_n113 ) , .ZN( u1_u13_u3_n131 ) , .A2( u1_u13_u3_n154 ) );
  NAND2_X1 u1_u13_u3_U49 (.A1( u1_u13_u3_n103 ) , .ZN( u1_u13_u3_n150 ) , .A2( u1_u13_u3_n99 ) );
  INV_X1 u1_u13_u3_U5 (.A( u1_u13_u3_n117 ) , .ZN( u1_u13_u3_n178 ) );
  NAND2_X1 u1_u13_u3_U50 (.A2( u1_u13_u3_n102 ) , .ZN( u1_u13_u3_n155 ) , .A1( u1_u13_u3_n97 ) );
  INV_X1 u1_u13_u3_U51 (.A( u1_u13_u3_n141 ) , .ZN( u1_u13_u3_n167 ) );
  AOI21_X1 u1_u13_u3_U52 (.B2( u1_u13_u3_n114 ) , .B1( u1_u13_u3_n146 ) , .A( u1_u13_u3_n154 ) , .ZN( u1_u13_u3_n94 ) );
  AOI21_X1 u1_u13_u3_U53 (.ZN( u1_u13_u3_n110 ) , .B2( u1_u13_u3_n142 ) , .B1( u1_u13_u3_n186 ) , .A( u1_u13_u3_n95 ) );
  INV_X1 u1_u13_u3_U54 (.A( u1_u13_u3_n145 ) , .ZN( u1_u13_u3_n186 ) );
  AOI21_X1 u1_u13_u3_U55 (.B1( u1_u13_u3_n124 ) , .A( u1_u13_u3_n149 ) , .B2( u1_u13_u3_n155 ) , .ZN( u1_u13_u3_n95 ) );
  INV_X1 u1_u13_u3_U56 (.A( u1_u13_u3_n149 ) , .ZN( u1_u13_u3_n169 ) );
  NAND2_X1 u1_u13_u3_U57 (.ZN( u1_u13_u3_n124 ) , .A1( u1_u13_u3_n96 ) , .A2( u1_u13_u3_n97 ) );
  NAND2_X1 u1_u13_u3_U58 (.A2( u1_u13_u3_n100 ) , .ZN( u1_u13_u3_n146 ) , .A1( u1_u13_u3_n96 ) );
  NAND2_X1 u1_u13_u3_U59 (.A1( u1_u13_u3_n101 ) , .ZN( u1_u13_u3_n145 ) , .A2( u1_u13_u3_n99 ) );
  AOI221_X1 u1_u13_u3_U6 (.A( u1_u13_u3_n131 ) , .C2( u1_u13_u3_n132 ) , .C1( u1_u13_u3_n133 ) , .ZN( u1_u13_u3_n134 ) , .B1( u1_u13_u3_n143 ) , .B2( u1_u13_u3_n177 ) );
  NAND2_X1 u1_u13_u3_U60 (.A1( u1_u13_u3_n100 ) , .ZN( u1_u13_u3_n156 ) , .A2( u1_u13_u3_n99 ) );
  NAND2_X1 u1_u13_u3_U61 (.A2( u1_u13_u3_n101 ) , .A1( u1_u13_u3_n104 ) , .ZN( u1_u13_u3_n148 ) );
  NAND2_X1 u1_u13_u3_U62 (.A1( u1_u13_u3_n100 ) , .A2( u1_u13_u3_n102 ) , .ZN( u1_u13_u3_n128 ) );
  NAND2_X1 u1_u13_u3_U63 (.A2( u1_u13_u3_n101 ) , .A1( u1_u13_u3_n102 ) , .ZN( u1_u13_u3_n152 ) );
  NAND2_X1 u1_u13_u3_U64 (.A2( u1_u13_u3_n101 ) , .ZN( u1_u13_u3_n114 ) , .A1( u1_u13_u3_n96 ) );
  NAND2_X1 u1_u13_u3_U65 (.ZN( u1_u13_u3_n107 ) , .A1( u1_u13_u3_n97 ) , .A2( u1_u13_u3_n99 ) );
  NAND2_X1 u1_u13_u3_U66 (.A2( u1_u13_u3_n100 ) , .A1( u1_u13_u3_n104 ) , .ZN( u1_u13_u3_n113 ) );
  NAND2_X1 u1_u13_u3_U67 (.A1( u1_u13_u3_n104 ) , .ZN( u1_u13_u3_n153 ) , .A2( u1_u13_u3_n97 ) );
  NAND2_X1 u1_u13_u3_U68 (.A2( u1_u13_u3_n103 ) , .A1( u1_u13_u3_n104 ) , .ZN( u1_u13_u3_n130 ) );
  NAND2_X1 u1_u13_u3_U69 (.A2( u1_u13_u3_n103 ) , .ZN( u1_u13_u3_n144 ) , .A1( u1_u13_u3_n96 ) );
  OAI22_X1 u1_u13_u3_U7 (.B2( u1_u13_u3_n147 ) , .A2( u1_u13_u3_n148 ) , .ZN( u1_u13_u3_n160 ) , .B1( u1_u13_u3_n165 ) , .A1( u1_u13_u3_n168 ) );
  NAND2_X1 u1_u13_u3_U70 (.A1( u1_u13_u3_n102 ) , .A2( u1_u13_u3_n103 ) , .ZN( u1_u13_u3_n108 ) );
  NOR2_X1 u1_u13_u3_U71 (.A2( u1_u13_X_19 ) , .A1( u1_u13_X_20 ) , .ZN( u1_u13_u3_n99 ) );
  NOR2_X1 u1_u13_u3_U72 (.A2( u1_u13_X_21 ) , .A1( u1_u13_X_24 ) , .ZN( u1_u13_u3_n103 ) );
  NOR2_X1 u1_u13_u3_U73 (.A2( u1_u13_X_24 ) , .A1( u1_u13_u3_n171 ) , .ZN( u1_u13_u3_n97 ) );
  NOR2_X1 u1_u13_u3_U74 (.A2( u1_u13_X_23 ) , .ZN( u1_u13_u3_n141 ) , .A1( u1_u13_u3_n166 ) );
  NOR2_X1 u1_u13_u3_U75 (.A2( u1_u13_X_19 ) , .A1( u1_u13_u3_n172 ) , .ZN( u1_u13_u3_n96 ) );
  NAND2_X1 u1_u13_u3_U76 (.A1( u1_u13_X_22 ) , .A2( u1_u13_X_23 ) , .ZN( u1_u13_u3_n154 ) );
  NAND2_X1 u1_u13_u3_U77 (.A1( u1_u13_X_23 ) , .ZN( u1_u13_u3_n149 ) , .A2( u1_u13_u3_n166 ) );
  NOR2_X1 u1_u13_u3_U78 (.A2( u1_u13_X_22 ) , .A1( u1_u13_X_23 ) , .ZN( u1_u13_u3_n121 ) );
  AND2_X1 u1_u13_u3_U79 (.A1( u1_u13_X_24 ) , .ZN( u1_u13_u3_n101 ) , .A2( u1_u13_u3_n171 ) );
  AND3_X1 u1_u13_u3_U8 (.A3( u1_u13_u3_n144 ) , .A2( u1_u13_u3_n145 ) , .A1( u1_u13_u3_n146 ) , .ZN( u1_u13_u3_n147 ) );
  AND2_X1 u1_u13_u3_U80 (.A1( u1_u13_X_19 ) , .ZN( u1_u13_u3_n102 ) , .A2( u1_u13_u3_n172 ) );
  AND2_X1 u1_u13_u3_U81 (.A1( u1_u13_X_21 ) , .A2( u1_u13_X_24 ) , .ZN( u1_u13_u3_n100 ) );
  AND2_X1 u1_u13_u3_U82 (.A2( u1_u13_X_19 ) , .A1( u1_u13_X_20 ) , .ZN( u1_u13_u3_n104 ) );
  INV_X1 u1_u13_u3_U83 (.A( u1_u13_X_22 ) , .ZN( u1_u13_u3_n166 ) );
  INV_X1 u1_u13_u3_U84 (.A( u1_u13_X_21 ) , .ZN( u1_u13_u3_n171 ) );
  INV_X1 u1_u13_u3_U85 (.A( u1_u13_X_20 ) , .ZN( u1_u13_u3_n172 ) );
  NAND4_X1 u1_u13_u3_U86 (.ZN( u1_out13_26 ) , .A4( u1_u13_u3_n109 ) , .A3( u1_u13_u3_n110 ) , .A2( u1_u13_u3_n111 ) , .A1( u1_u13_u3_n173 ) );
  INV_X1 u1_u13_u3_U87 (.ZN( u1_u13_u3_n173 ) , .A( u1_u13_u3_n94 ) );
  OAI21_X1 u1_u13_u3_U88 (.ZN( u1_u13_u3_n111 ) , .B2( u1_u13_u3_n117 ) , .A( u1_u13_u3_n133 ) , .B1( u1_u13_u3_n176 ) );
  NAND4_X1 u1_u13_u3_U89 (.ZN( u1_out13_20 ) , .A4( u1_u13_u3_n122 ) , .A3( u1_u13_u3_n123 ) , .A1( u1_u13_u3_n175 ) , .A2( u1_u13_u3_n180 ) );
  INV_X1 u1_u13_u3_U9 (.A( u1_u13_u3_n143 ) , .ZN( u1_u13_u3_n168 ) );
  INV_X1 u1_u13_u3_U90 (.A( u1_u13_u3_n112 ) , .ZN( u1_u13_u3_n175 ) );
  INV_X1 u1_u13_u3_U91 (.A( u1_u13_u3_n126 ) , .ZN( u1_u13_u3_n180 ) );
  NAND4_X1 u1_u13_u3_U92 (.ZN( u1_out13_1 ) , .A4( u1_u13_u3_n161 ) , .A3( u1_u13_u3_n162 ) , .A2( u1_u13_u3_n163 ) , .A1( u1_u13_u3_n185 ) );
  NAND2_X1 u1_u13_u3_U93 (.ZN( u1_u13_u3_n163 ) , .A2( u1_u13_u3_n170 ) , .A1( u1_u13_u3_n176 ) );
  AOI22_X1 u1_u13_u3_U94 (.B2( u1_u13_u3_n140 ) , .B1( u1_u13_u3_n141 ) , .A2( u1_u13_u3_n142 ) , .ZN( u1_u13_u3_n162 ) , .A1( u1_u13_u3_n177 ) );
  OR4_X1 u1_u13_u3_U95 (.ZN( u1_out13_10 ) , .A4( u1_u13_u3_n136 ) , .A3( u1_u13_u3_n137 ) , .A1( u1_u13_u3_n138 ) , .A2( u1_u13_u3_n139 ) );
  OAI222_X1 u1_u13_u3_U96 (.C1( u1_u13_u3_n128 ) , .ZN( u1_u13_u3_n137 ) , .B1( u1_u13_u3_n148 ) , .A2( u1_u13_u3_n150 ) , .B2( u1_u13_u3_n154 ) , .C2( u1_u13_u3_n164 ) , .A1( u1_u13_u3_n167 ) );
  OAI221_X1 u1_u13_u3_U97 (.A( u1_u13_u3_n134 ) , .B2( u1_u13_u3_n135 ) , .ZN( u1_u13_u3_n136 ) , .C1( u1_u13_u3_n149 ) , .B1( u1_u13_u3_n151 ) , .C2( u1_u13_u3_n183 ) );
  NAND3_X1 u1_u13_u3_U98 (.A1( u1_u13_u3_n114 ) , .ZN( u1_u13_u3_n115 ) , .A2( u1_u13_u3_n145 ) , .A3( u1_u13_u3_n153 ) );
  NAND3_X1 u1_u13_u3_U99 (.ZN( u1_u13_u3_n129 ) , .A2( u1_u13_u3_n144 ) , .A1( u1_u13_u3_n153 ) , .A3( u1_u13_u3_n182 ) );
  XOR2_X1 u1_u2_U10 (.B( u1_K3_45 ) , .A( u1_R1_30 ) , .Z( u1_u2_X_45 ) );
  XOR2_X1 u1_u2_U11 (.B( u1_K3_44 ) , .A( u1_R1_29 ) , .Z( u1_u2_X_44 ) );
  XOR2_X1 u1_u2_U12 (.B( u1_K3_43 ) , .A( u1_R1_28 ) , .Z( u1_u2_X_43 ) );
  XOR2_X1 u1_u2_U13 (.B( u1_K3_42 ) , .A( u1_R1_29 ) , .Z( u1_u2_X_42 ) );
  XOR2_X1 u1_u2_U14 (.B( u1_K3_41 ) , .A( u1_R1_28 ) , .Z( u1_u2_X_41 ) );
  XOR2_X1 u1_u2_U15 (.B( u1_K3_40 ) , .A( u1_R1_27 ) , .Z( u1_u2_X_40 ) );
  XOR2_X1 u1_u2_U17 (.B( u1_K3_39 ) , .A( u1_R1_26 ) , .Z( u1_u2_X_39 ) );
  XOR2_X1 u1_u2_U18 (.B( u1_K3_38 ) , .A( u1_R1_25 ) , .Z( u1_u2_X_38 ) );
  XOR2_X1 u1_u2_U19 (.B( u1_K3_37 ) , .A( u1_R1_24 ) , .Z( u1_u2_X_37 ) );
  XOR2_X1 u1_u2_U7 (.B( u1_K3_48 ) , .A( u1_R1_1 ) , .Z( u1_u2_X_48 ) );
  XOR2_X1 u1_u2_U8 (.B( u1_K3_47 ) , .A( u1_R1_32 ) , .Z( u1_u2_X_47 ) );
  XOR2_X1 u1_u2_U9 (.B( u1_K3_46 ) , .A( u1_R1_31 ) , .Z( u1_u2_X_46 ) );
  OAI21_X1 u1_u2_u6_U10 (.A( u1_u2_u6_n159 ) , .B1( u1_u2_u6_n169 ) , .B2( u1_u2_u6_n173 ) , .ZN( u1_u2_u6_n90 ) );
  INV_X1 u1_u2_u6_U11 (.ZN( u1_u2_u6_n172 ) , .A( u1_u2_u6_n88 ) );
  AOI22_X1 u1_u2_u6_U12 (.A2( u1_u2_u6_n151 ) , .B2( u1_u2_u6_n161 ) , .A1( u1_u2_u6_n167 ) , .B1( u1_u2_u6_n170 ) , .ZN( u1_u2_u6_n89 ) );
  AOI21_X1 u1_u2_u6_U13 (.ZN( u1_u2_u6_n106 ) , .A( u1_u2_u6_n142 ) , .B2( u1_u2_u6_n159 ) , .B1( u1_u2_u6_n164 ) );
  INV_X1 u1_u2_u6_U14 (.A( u1_u2_u6_n155 ) , .ZN( u1_u2_u6_n161 ) );
  INV_X1 u1_u2_u6_U15 (.A( u1_u2_u6_n128 ) , .ZN( u1_u2_u6_n164 ) );
  NAND2_X1 u1_u2_u6_U16 (.ZN( u1_u2_u6_n110 ) , .A1( u1_u2_u6_n122 ) , .A2( u1_u2_u6_n129 ) );
  NAND2_X1 u1_u2_u6_U17 (.ZN( u1_u2_u6_n124 ) , .A2( u1_u2_u6_n146 ) , .A1( u1_u2_u6_n148 ) );
  INV_X1 u1_u2_u6_U18 (.A( u1_u2_u6_n132 ) , .ZN( u1_u2_u6_n171 ) );
  AND2_X1 u1_u2_u6_U19 (.A1( u1_u2_u6_n100 ) , .ZN( u1_u2_u6_n130 ) , .A2( u1_u2_u6_n147 ) );
  INV_X1 u1_u2_u6_U20 (.A( u1_u2_u6_n127 ) , .ZN( u1_u2_u6_n173 ) );
  INV_X1 u1_u2_u6_U21 (.A( u1_u2_u6_n121 ) , .ZN( u1_u2_u6_n167 ) );
  INV_X1 u1_u2_u6_U22 (.A( u1_u2_u6_n100 ) , .ZN( u1_u2_u6_n169 ) );
  INV_X1 u1_u2_u6_U23 (.A( u1_u2_u6_n123 ) , .ZN( u1_u2_u6_n170 ) );
  INV_X1 u1_u2_u6_U24 (.A( u1_u2_u6_n113 ) , .ZN( u1_u2_u6_n168 ) );
  AND2_X1 u1_u2_u6_U25 (.A1( u1_u2_u6_n107 ) , .A2( u1_u2_u6_n119 ) , .ZN( u1_u2_u6_n133 ) );
  AND2_X1 u1_u2_u6_U26 (.A2( u1_u2_u6_n121 ) , .A1( u1_u2_u6_n122 ) , .ZN( u1_u2_u6_n131 ) );
  AND3_X1 u1_u2_u6_U27 (.ZN( u1_u2_u6_n120 ) , .A2( u1_u2_u6_n127 ) , .A1( u1_u2_u6_n132 ) , .A3( u1_u2_u6_n145 ) );
  INV_X1 u1_u2_u6_U28 (.A( u1_u2_u6_n146 ) , .ZN( u1_u2_u6_n163 ) );
  AOI222_X1 u1_u2_u6_U29 (.ZN( u1_u2_u6_n114 ) , .A1( u1_u2_u6_n118 ) , .A2( u1_u2_u6_n126 ) , .B2( u1_u2_u6_n151 ) , .C2( u1_u2_u6_n159 ) , .C1( u1_u2_u6_n168 ) , .B1( u1_u2_u6_n169 ) );
  INV_X1 u1_u2_u6_U3 (.A( u1_u2_u6_n110 ) , .ZN( u1_u2_u6_n166 ) );
  NOR2_X1 u1_u2_u6_U30 (.A1( u1_u2_u6_n162 ) , .A2( u1_u2_u6_n165 ) , .ZN( u1_u2_u6_n98 ) );
  NAND2_X1 u1_u2_u6_U31 (.A1( u1_u2_u6_n144 ) , .ZN( u1_u2_u6_n151 ) , .A2( u1_u2_u6_n158 ) );
  NAND2_X1 u1_u2_u6_U32 (.ZN( u1_u2_u6_n132 ) , .A1( u1_u2_u6_n91 ) , .A2( u1_u2_u6_n97 ) );
  AOI22_X1 u1_u2_u6_U33 (.B2( u1_u2_u6_n110 ) , .B1( u1_u2_u6_n111 ) , .A1( u1_u2_u6_n112 ) , .ZN( u1_u2_u6_n115 ) , .A2( u1_u2_u6_n161 ) );
  NAND4_X1 u1_u2_u6_U34 (.A3( u1_u2_u6_n109 ) , .ZN( u1_u2_u6_n112 ) , .A4( u1_u2_u6_n132 ) , .A2( u1_u2_u6_n147 ) , .A1( u1_u2_u6_n166 ) );
  NOR2_X1 u1_u2_u6_U35 (.ZN( u1_u2_u6_n109 ) , .A1( u1_u2_u6_n170 ) , .A2( u1_u2_u6_n173 ) );
  NOR2_X1 u1_u2_u6_U36 (.A2( u1_u2_u6_n126 ) , .ZN( u1_u2_u6_n155 ) , .A1( u1_u2_u6_n160 ) );
  NAND2_X1 u1_u2_u6_U37 (.ZN( u1_u2_u6_n146 ) , .A2( u1_u2_u6_n94 ) , .A1( u1_u2_u6_n99 ) );
  AOI21_X1 u1_u2_u6_U38 (.A( u1_u2_u6_n144 ) , .B2( u1_u2_u6_n145 ) , .B1( u1_u2_u6_n146 ) , .ZN( u1_u2_u6_n150 ) );
  INV_X1 u1_u2_u6_U39 (.A( u1_u2_u6_n111 ) , .ZN( u1_u2_u6_n158 ) );
  INV_X1 u1_u2_u6_U4 (.A( u1_u2_u6_n142 ) , .ZN( u1_u2_u6_n174 ) );
  NAND2_X1 u1_u2_u6_U40 (.ZN( u1_u2_u6_n127 ) , .A1( u1_u2_u6_n91 ) , .A2( u1_u2_u6_n92 ) );
  NAND2_X1 u1_u2_u6_U41 (.ZN( u1_u2_u6_n129 ) , .A2( u1_u2_u6_n95 ) , .A1( u1_u2_u6_n96 ) );
  INV_X1 u1_u2_u6_U42 (.A( u1_u2_u6_n144 ) , .ZN( u1_u2_u6_n159 ) );
  NAND2_X1 u1_u2_u6_U43 (.ZN( u1_u2_u6_n145 ) , .A2( u1_u2_u6_n97 ) , .A1( u1_u2_u6_n98 ) );
  NAND2_X1 u1_u2_u6_U44 (.ZN( u1_u2_u6_n148 ) , .A2( u1_u2_u6_n92 ) , .A1( u1_u2_u6_n94 ) );
  NAND2_X1 u1_u2_u6_U45 (.ZN( u1_u2_u6_n108 ) , .A2( u1_u2_u6_n139 ) , .A1( u1_u2_u6_n144 ) );
  NAND2_X1 u1_u2_u6_U46 (.ZN( u1_u2_u6_n121 ) , .A2( u1_u2_u6_n95 ) , .A1( u1_u2_u6_n97 ) );
  NAND2_X1 u1_u2_u6_U47 (.ZN( u1_u2_u6_n107 ) , .A2( u1_u2_u6_n92 ) , .A1( u1_u2_u6_n95 ) );
  AND2_X1 u1_u2_u6_U48 (.ZN( u1_u2_u6_n118 ) , .A2( u1_u2_u6_n91 ) , .A1( u1_u2_u6_n99 ) );
  NAND2_X1 u1_u2_u6_U49 (.ZN( u1_u2_u6_n147 ) , .A2( u1_u2_u6_n98 ) , .A1( u1_u2_u6_n99 ) );
  NAND2_X1 u1_u2_u6_U5 (.A2( u1_u2_u6_n143 ) , .ZN( u1_u2_u6_n152 ) , .A1( u1_u2_u6_n166 ) );
  NAND2_X1 u1_u2_u6_U50 (.ZN( u1_u2_u6_n128 ) , .A1( u1_u2_u6_n94 ) , .A2( u1_u2_u6_n96 ) );
  AOI211_X1 u1_u2_u6_U51 (.B( u1_u2_u6_n134 ) , .A( u1_u2_u6_n135 ) , .C1( u1_u2_u6_n136 ) , .ZN( u1_u2_u6_n137 ) , .C2( u1_u2_u6_n151 ) );
  AOI21_X1 u1_u2_u6_U52 (.B2( u1_u2_u6_n132 ) , .B1( u1_u2_u6_n133 ) , .ZN( u1_u2_u6_n134 ) , .A( u1_u2_u6_n158 ) );
  AOI21_X1 u1_u2_u6_U53 (.B1( u1_u2_u6_n131 ) , .ZN( u1_u2_u6_n135 ) , .A( u1_u2_u6_n144 ) , .B2( u1_u2_u6_n146 ) );
  NAND4_X1 u1_u2_u6_U54 (.A4( u1_u2_u6_n127 ) , .A3( u1_u2_u6_n128 ) , .A2( u1_u2_u6_n129 ) , .A1( u1_u2_u6_n130 ) , .ZN( u1_u2_u6_n136 ) );
  NAND2_X1 u1_u2_u6_U55 (.ZN( u1_u2_u6_n119 ) , .A2( u1_u2_u6_n95 ) , .A1( u1_u2_u6_n99 ) );
  NAND2_X1 u1_u2_u6_U56 (.ZN( u1_u2_u6_n123 ) , .A2( u1_u2_u6_n91 ) , .A1( u1_u2_u6_n96 ) );
  NAND2_X1 u1_u2_u6_U57 (.ZN( u1_u2_u6_n100 ) , .A2( u1_u2_u6_n92 ) , .A1( u1_u2_u6_n98 ) );
  NAND2_X1 u1_u2_u6_U58 (.ZN( u1_u2_u6_n122 ) , .A1( u1_u2_u6_n94 ) , .A2( u1_u2_u6_n97 ) );
  INV_X1 u1_u2_u6_U59 (.A( u1_u2_u6_n139 ) , .ZN( u1_u2_u6_n160 ) );
  AOI22_X1 u1_u2_u6_U6 (.B2( u1_u2_u6_n101 ) , .A1( u1_u2_u6_n102 ) , .ZN( u1_u2_u6_n103 ) , .B1( u1_u2_u6_n160 ) , .A2( u1_u2_u6_n161 ) );
  NAND2_X1 u1_u2_u6_U60 (.ZN( u1_u2_u6_n113 ) , .A1( u1_u2_u6_n96 ) , .A2( u1_u2_u6_n98 ) );
  NOR2_X1 u1_u2_u6_U61 (.A2( u1_u2_X_40 ) , .A1( u1_u2_X_41 ) , .ZN( u1_u2_u6_n126 ) );
  NOR2_X1 u1_u2_u6_U62 (.A2( u1_u2_X_39 ) , .A1( u1_u2_X_42 ) , .ZN( u1_u2_u6_n92 ) );
  NOR2_X1 u1_u2_u6_U63 (.A2( u1_u2_X_39 ) , .A1( u1_u2_u6_n156 ) , .ZN( u1_u2_u6_n97 ) );
  NOR2_X1 u1_u2_u6_U64 (.A2( u1_u2_X_38 ) , .A1( u1_u2_u6_n165 ) , .ZN( u1_u2_u6_n95 ) );
  NOR2_X1 u1_u2_u6_U65 (.A2( u1_u2_X_41 ) , .ZN( u1_u2_u6_n111 ) , .A1( u1_u2_u6_n157 ) );
  NOR2_X1 u1_u2_u6_U66 (.A2( u1_u2_X_37 ) , .A1( u1_u2_u6_n162 ) , .ZN( u1_u2_u6_n94 ) );
  NOR2_X1 u1_u2_u6_U67 (.A2( u1_u2_X_37 ) , .A1( u1_u2_X_38 ) , .ZN( u1_u2_u6_n91 ) );
  NAND2_X1 u1_u2_u6_U68 (.A1( u1_u2_X_41 ) , .ZN( u1_u2_u6_n144 ) , .A2( u1_u2_u6_n157 ) );
  NAND2_X1 u1_u2_u6_U69 (.A2( u1_u2_X_40 ) , .A1( u1_u2_X_41 ) , .ZN( u1_u2_u6_n139 ) );
  NOR2_X1 u1_u2_u6_U7 (.A1( u1_u2_u6_n118 ) , .ZN( u1_u2_u6_n143 ) , .A2( u1_u2_u6_n168 ) );
  AND2_X1 u1_u2_u6_U70 (.A1( u1_u2_X_39 ) , .A2( u1_u2_u6_n156 ) , .ZN( u1_u2_u6_n96 ) );
  AND2_X1 u1_u2_u6_U71 (.A1( u1_u2_X_39 ) , .A2( u1_u2_X_42 ) , .ZN( u1_u2_u6_n99 ) );
  INV_X1 u1_u2_u6_U72 (.A( u1_u2_X_40 ) , .ZN( u1_u2_u6_n157 ) );
  INV_X1 u1_u2_u6_U73 (.A( u1_u2_X_37 ) , .ZN( u1_u2_u6_n165 ) );
  INV_X1 u1_u2_u6_U74 (.A( u1_u2_X_38 ) , .ZN( u1_u2_u6_n162 ) );
  INV_X1 u1_u2_u6_U75 (.A( u1_u2_X_42 ) , .ZN( u1_u2_u6_n156 ) );
  NAND4_X1 u1_u2_u6_U76 (.ZN( u1_out2_32 ) , .A4( u1_u2_u6_n103 ) , .A3( u1_u2_u6_n104 ) , .A2( u1_u2_u6_n105 ) , .A1( u1_u2_u6_n106 ) );
  AOI22_X1 u1_u2_u6_U77 (.ZN( u1_u2_u6_n105 ) , .A2( u1_u2_u6_n108 ) , .A1( u1_u2_u6_n118 ) , .B2( u1_u2_u6_n126 ) , .B1( u1_u2_u6_n171 ) );
  AOI22_X1 u1_u2_u6_U78 (.ZN( u1_u2_u6_n104 ) , .A1( u1_u2_u6_n111 ) , .B1( u1_u2_u6_n124 ) , .B2( u1_u2_u6_n151 ) , .A2( u1_u2_u6_n93 ) );
  NAND4_X1 u1_u2_u6_U79 (.ZN( u1_out2_12 ) , .A4( u1_u2_u6_n114 ) , .A3( u1_u2_u6_n115 ) , .A2( u1_u2_u6_n116 ) , .A1( u1_u2_u6_n117 ) );
  AOI21_X1 u1_u2_u6_U8 (.B1( u1_u2_u6_n107 ) , .B2( u1_u2_u6_n132 ) , .A( u1_u2_u6_n158 ) , .ZN( u1_u2_u6_n88 ) );
  OAI22_X1 u1_u2_u6_U80 (.B2( u1_u2_u6_n111 ) , .ZN( u1_u2_u6_n116 ) , .B1( u1_u2_u6_n126 ) , .A2( u1_u2_u6_n164 ) , .A1( u1_u2_u6_n167 ) );
  OAI21_X1 u1_u2_u6_U81 (.A( u1_u2_u6_n108 ) , .ZN( u1_u2_u6_n117 ) , .B2( u1_u2_u6_n141 ) , .B1( u1_u2_u6_n163 ) );
  OAI211_X1 u1_u2_u6_U82 (.ZN( u1_out2_7 ) , .B( u1_u2_u6_n153 ) , .C2( u1_u2_u6_n154 ) , .C1( u1_u2_u6_n155 ) , .A( u1_u2_u6_n174 ) );
  NOR3_X1 u1_u2_u6_U83 (.A1( u1_u2_u6_n141 ) , .ZN( u1_u2_u6_n154 ) , .A3( u1_u2_u6_n164 ) , .A2( u1_u2_u6_n171 ) );
  AOI211_X1 u1_u2_u6_U84 (.B( u1_u2_u6_n149 ) , .A( u1_u2_u6_n150 ) , .C2( u1_u2_u6_n151 ) , .C1( u1_u2_u6_n152 ) , .ZN( u1_u2_u6_n153 ) );
  OAI211_X1 u1_u2_u6_U85 (.ZN( u1_out2_22 ) , .B( u1_u2_u6_n137 ) , .A( u1_u2_u6_n138 ) , .C2( u1_u2_u6_n139 ) , .C1( u1_u2_u6_n140 ) );
  AOI22_X1 u1_u2_u6_U86 (.B1( u1_u2_u6_n124 ) , .A2( u1_u2_u6_n125 ) , .A1( u1_u2_u6_n126 ) , .ZN( u1_u2_u6_n138 ) , .B2( u1_u2_u6_n161 ) );
  AND4_X1 u1_u2_u6_U87 (.A3( u1_u2_u6_n119 ) , .A1( u1_u2_u6_n120 ) , .A4( u1_u2_u6_n129 ) , .ZN( u1_u2_u6_n140 ) , .A2( u1_u2_u6_n143 ) );
  NAND3_X1 u1_u2_u6_U88 (.A2( u1_u2_u6_n123 ) , .ZN( u1_u2_u6_n125 ) , .A1( u1_u2_u6_n130 ) , .A3( u1_u2_u6_n131 ) );
  NAND3_X1 u1_u2_u6_U89 (.A3( u1_u2_u6_n133 ) , .ZN( u1_u2_u6_n141 ) , .A1( u1_u2_u6_n145 ) , .A2( u1_u2_u6_n148 ) );
  AOI21_X1 u1_u2_u6_U9 (.B2( u1_u2_u6_n147 ) , .B1( u1_u2_u6_n148 ) , .ZN( u1_u2_u6_n149 ) , .A( u1_u2_u6_n158 ) );
  NAND3_X1 u1_u2_u6_U90 (.ZN( u1_u2_u6_n101 ) , .A3( u1_u2_u6_n107 ) , .A2( u1_u2_u6_n121 ) , .A1( u1_u2_u6_n127 ) );
  NAND3_X1 u1_u2_u6_U91 (.ZN( u1_u2_u6_n102 ) , .A3( u1_u2_u6_n130 ) , .A2( u1_u2_u6_n145 ) , .A1( u1_u2_u6_n166 ) );
  NAND3_X1 u1_u2_u6_U92 (.A3( u1_u2_u6_n113 ) , .A1( u1_u2_u6_n119 ) , .A2( u1_u2_u6_n123 ) , .ZN( u1_u2_u6_n93 ) );
  NAND3_X1 u1_u2_u6_U93 (.ZN( u1_u2_u6_n142 ) , .A2( u1_u2_u6_n172 ) , .A3( u1_u2_u6_n89 ) , .A1( u1_u2_u6_n90 ) );
  AND3_X1 u1_u2_u7_U10 (.A3( u1_u2_u7_n110 ) , .A2( u1_u2_u7_n127 ) , .A1( u1_u2_u7_n132 ) , .ZN( u1_u2_u7_n92 ) );
  OAI21_X1 u1_u2_u7_U11 (.A( u1_u2_u7_n161 ) , .B1( u1_u2_u7_n168 ) , .B2( u1_u2_u7_n173 ) , .ZN( u1_u2_u7_n91 ) );
  AOI211_X1 u1_u2_u7_U12 (.A( u1_u2_u7_n117 ) , .ZN( u1_u2_u7_n118 ) , .C2( u1_u2_u7_n126 ) , .C1( u1_u2_u7_n177 ) , .B( u1_u2_u7_n180 ) );
  OAI22_X1 u1_u2_u7_U13 (.B1( u1_u2_u7_n115 ) , .ZN( u1_u2_u7_n117 ) , .A2( u1_u2_u7_n133 ) , .A1( u1_u2_u7_n137 ) , .B2( u1_u2_u7_n162 ) );
  INV_X1 u1_u2_u7_U14 (.A( u1_u2_u7_n116 ) , .ZN( u1_u2_u7_n180 ) );
  NOR3_X1 u1_u2_u7_U15 (.ZN( u1_u2_u7_n115 ) , .A3( u1_u2_u7_n145 ) , .A2( u1_u2_u7_n168 ) , .A1( u1_u2_u7_n169 ) );
  OAI211_X1 u1_u2_u7_U16 (.B( u1_u2_u7_n122 ) , .A( u1_u2_u7_n123 ) , .C2( u1_u2_u7_n124 ) , .ZN( u1_u2_u7_n154 ) , .C1( u1_u2_u7_n162 ) );
  AOI222_X1 u1_u2_u7_U17 (.ZN( u1_u2_u7_n122 ) , .C2( u1_u2_u7_n126 ) , .C1( u1_u2_u7_n145 ) , .B1( u1_u2_u7_n161 ) , .A2( u1_u2_u7_n165 ) , .B2( u1_u2_u7_n170 ) , .A1( u1_u2_u7_n176 ) );
  INV_X1 u1_u2_u7_U18 (.A( u1_u2_u7_n133 ) , .ZN( u1_u2_u7_n176 ) );
  NOR3_X1 u1_u2_u7_U19 (.A2( u1_u2_u7_n134 ) , .A1( u1_u2_u7_n135 ) , .ZN( u1_u2_u7_n136 ) , .A3( u1_u2_u7_n171 ) );
  NOR2_X1 u1_u2_u7_U20 (.A1( u1_u2_u7_n130 ) , .A2( u1_u2_u7_n134 ) , .ZN( u1_u2_u7_n153 ) );
  INV_X1 u1_u2_u7_U21 (.A( u1_u2_u7_n101 ) , .ZN( u1_u2_u7_n165 ) );
  NOR2_X1 u1_u2_u7_U22 (.ZN( u1_u2_u7_n111 ) , .A2( u1_u2_u7_n134 ) , .A1( u1_u2_u7_n169 ) );
  AOI21_X1 u1_u2_u7_U23 (.ZN( u1_u2_u7_n104 ) , .B2( u1_u2_u7_n112 ) , .B1( u1_u2_u7_n127 ) , .A( u1_u2_u7_n164 ) );
  AOI21_X1 u1_u2_u7_U24 (.ZN( u1_u2_u7_n106 ) , .B1( u1_u2_u7_n133 ) , .B2( u1_u2_u7_n146 ) , .A( u1_u2_u7_n162 ) );
  AOI21_X1 u1_u2_u7_U25 (.A( u1_u2_u7_n101 ) , .ZN( u1_u2_u7_n107 ) , .B2( u1_u2_u7_n128 ) , .B1( u1_u2_u7_n175 ) );
  INV_X1 u1_u2_u7_U26 (.A( u1_u2_u7_n138 ) , .ZN( u1_u2_u7_n171 ) );
  INV_X1 u1_u2_u7_U27 (.A( u1_u2_u7_n131 ) , .ZN( u1_u2_u7_n177 ) );
  INV_X1 u1_u2_u7_U28 (.A( u1_u2_u7_n110 ) , .ZN( u1_u2_u7_n174 ) );
  NAND2_X1 u1_u2_u7_U29 (.A1( u1_u2_u7_n129 ) , .A2( u1_u2_u7_n132 ) , .ZN( u1_u2_u7_n149 ) );
  OAI21_X1 u1_u2_u7_U3 (.ZN( u1_u2_u7_n159 ) , .A( u1_u2_u7_n165 ) , .B2( u1_u2_u7_n171 ) , .B1( u1_u2_u7_n174 ) );
  NAND2_X1 u1_u2_u7_U30 (.A1( u1_u2_u7_n113 ) , .A2( u1_u2_u7_n124 ) , .ZN( u1_u2_u7_n130 ) );
  INV_X1 u1_u2_u7_U31 (.A( u1_u2_u7_n112 ) , .ZN( u1_u2_u7_n173 ) );
  INV_X1 u1_u2_u7_U32 (.A( u1_u2_u7_n128 ) , .ZN( u1_u2_u7_n168 ) );
  INV_X1 u1_u2_u7_U33 (.A( u1_u2_u7_n148 ) , .ZN( u1_u2_u7_n169 ) );
  INV_X1 u1_u2_u7_U34 (.A( u1_u2_u7_n127 ) , .ZN( u1_u2_u7_n179 ) );
  NOR2_X1 u1_u2_u7_U35 (.ZN( u1_u2_u7_n101 ) , .A2( u1_u2_u7_n150 ) , .A1( u1_u2_u7_n156 ) );
  AOI211_X1 u1_u2_u7_U36 (.B( u1_u2_u7_n154 ) , .A( u1_u2_u7_n155 ) , .C1( u1_u2_u7_n156 ) , .ZN( u1_u2_u7_n157 ) , .C2( u1_u2_u7_n172 ) );
  INV_X1 u1_u2_u7_U37 (.A( u1_u2_u7_n153 ) , .ZN( u1_u2_u7_n172 ) );
  AOI211_X1 u1_u2_u7_U38 (.B( u1_u2_u7_n139 ) , .A( u1_u2_u7_n140 ) , .C2( u1_u2_u7_n141 ) , .ZN( u1_u2_u7_n142 ) , .C1( u1_u2_u7_n156 ) );
  NAND4_X1 u1_u2_u7_U39 (.A3( u1_u2_u7_n127 ) , .A2( u1_u2_u7_n128 ) , .A1( u1_u2_u7_n129 ) , .ZN( u1_u2_u7_n141 ) , .A4( u1_u2_u7_n147 ) );
  INV_X1 u1_u2_u7_U4 (.A( u1_u2_u7_n111 ) , .ZN( u1_u2_u7_n170 ) );
  AOI21_X1 u1_u2_u7_U40 (.A( u1_u2_u7_n137 ) , .B1( u1_u2_u7_n138 ) , .ZN( u1_u2_u7_n139 ) , .B2( u1_u2_u7_n146 ) );
  OAI22_X1 u1_u2_u7_U41 (.B1( u1_u2_u7_n136 ) , .ZN( u1_u2_u7_n140 ) , .A1( u1_u2_u7_n153 ) , .B2( u1_u2_u7_n162 ) , .A2( u1_u2_u7_n164 ) );
  AOI21_X1 u1_u2_u7_U42 (.ZN( u1_u2_u7_n123 ) , .B1( u1_u2_u7_n165 ) , .B2( u1_u2_u7_n177 ) , .A( u1_u2_u7_n97 ) );
  AOI21_X1 u1_u2_u7_U43 (.B2( u1_u2_u7_n113 ) , .B1( u1_u2_u7_n124 ) , .A( u1_u2_u7_n125 ) , .ZN( u1_u2_u7_n97 ) );
  INV_X1 u1_u2_u7_U44 (.A( u1_u2_u7_n125 ) , .ZN( u1_u2_u7_n161 ) );
  INV_X1 u1_u2_u7_U45 (.A( u1_u2_u7_n152 ) , .ZN( u1_u2_u7_n162 ) );
  AOI22_X1 u1_u2_u7_U46 (.A2( u1_u2_u7_n114 ) , .ZN( u1_u2_u7_n119 ) , .B1( u1_u2_u7_n130 ) , .A1( u1_u2_u7_n156 ) , .B2( u1_u2_u7_n165 ) );
  NAND2_X1 u1_u2_u7_U47 (.A2( u1_u2_u7_n112 ) , .ZN( u1_u2_u7_n114 ) , .A1( u1_u2_u7_n175 ) );
  AND2_X1 u1_u2_u7_U48 (.ZN( u1_u2_u7_n145 ) , .A2( u1_u2_u7_n98 ) , .A1( u1_u2_u7_n99 ) );
  NOR2_X1 u1_u2_u7_U49 (.ZN( u1_u2_u7_n137 ) , .A1( u1_u2_u7_n150 ) , .A2( u1_u2_u7_n161 ) );
  INV_X1 u1_u2_u7_U5 (.A( u1_u2_u7_n149 ) , .ZN( u1_u2_u7_n175 ) );
  AOI21_X1 u1_u2_u7_U50 (.ZN( u1_u2_u7_n105 ) , .B2( u1_u2_u7_n110 ) , .A( u1_u2_u7_n125 ) , .B1( u1_u2_u7_n147 ) );
  NAND2_X1 u1_u2_u7_U51 (.ZN( u1_u2_u7_n146 ) , .A1( u1_u2_u7_n95 ) , .A2( u1_u2_u7_n98 ) );
  NAND2_X1 u1_u2_u7_U52 (.A2( u1_u2_u7_n103 ) , .ZN( u1_u2_u7_n147 ) , .A1( u1_u2_u7_n93 ) );
  NAND2_X1 u1_u2_u7_U53 (.A1( u1_u2_u7_n103 ) , .ZN( u1_u2_u7_n127 ) , .A2( u1_u2_u7_n99 ) );
  OR2_X1 u1_u2_u7_U54 (.ZN( u1_u2_u7_n126 ) , .A2( u1_u2_u7_n152 ) , .A1( u1_u2_u7_n156 ) );
  NAND2_X1 u1_u2_u7_U55 (.A2( u1_u2_u7_n102 ) , .A1( u1_u2_u7_n103 ) , .ZN( u1_u2_u7_n133 ) );
  NAND2_X1 u1_u2_u7_U56 (.ZN( u1_u2_u7_n112 ) , .A2( u1_u2_u7_n96 ) , .A1( u1_u2_u7_n99 ) );
  NAND2_X1 u1_u2_u7_U57 (.A2( u1_u2_u7_n102 ) , .ZN( u1_u2_u7_n128 ) , .A1( u1_u2_u7_n98 ) );
  NAND2_X1 u1_u2_u7_U58 (.A1( u1_u2_u7_n100 ) , .ZN( u1_u2_u7_n113 ) , .A2( u1_u2_u7_n93 ) );
  NAND2_X1 u1_u2_u7_U59 (.A2( u1_u2_u7_n102 ) , .ZN( u1_u2_u7_n124 ) , .A1( u1_u2_u7_n96 ) );
  INV_X1 u1_u2_u7_U6 (.A( u1_u2_u7_n154 ) , .ZN( u1_u2_u7_n178 ) );
  NAND2_X1 u1_u2_u7_U60 (.ZN( u1_u2_u7_n110 ) , .A1( u1_u2_u7_n95 ) , .A2( u1_u2_u7_n96 ) );
  INV_X1 u1_u2_u7_U61 (.A( u1_u2_u7_n150 ) , .ZN( u1_u2_u7_n164 ) );
  AND2_X1 u1_u2_u7_U62 (.ZN( u1_u2_u7_n134 ) , .A1( u1_u2_u7_n93 ) , .A2( u1_u2_u7_n98 ) );
  NAND2_X1 u1_u2_u7_U63 (.A1( u1_u2_u7_n100 ) , .A2( u1_u2_u7_n102 ) , .ZN( u1_u2_u7_n129 ) );
  NAND2_X1 u1_u2_u7_U64 (.A2( u1_u2_u7_n103 ) , .ZN( u1_u2_u7_n131 ) , .A1( u1_u2_u7_n95 ) );
  NAND2_X1 u1_u2_u7_U65 (.A1( u1_u2_u7_n100 ) , .ZN( u1_u2_u7_n138 ) , .A2( u1_u2_u7_n99 ) );
  NAND2_X1 u1_u2_u7_U66 (.ZN( u1_u2_u7_n132 ) , .A1( u1_u2_u7_n93 ) , .A2( u1_u2_u7_n96 ) );
  NAND2_X1 u1_u2_u7_U67 (.A1( u1_u2_u7_n100 ) , .ZN( u1_u2_u7_n148 ) , .A2( u1_u2_u7_n95 ) );
  NOR2_X1 u1_u2_u7_U68 (.A2( u1_u2_X_47 ) , .ZN( u1_u2_u7_n150 ) , .A1( u1_u2_u7_n163 ) );
  NOR2_X1 u1_u2_u7_U69 (.A2( u1_u2_X_43 ) , .A1( u1_u2_X_44 ) , .ZN( u1_u2_u7_n103 ) );
  AOI211_X1 u1_u2_u7_U7 (.ZN( u1_u2_u7_n116 ) , .A( u1_u2_u7_n155 ) , .C1( u1_u2_u7_n161 ) , .C2( u1_u2_u7_n171 ) , .B( u1_u2_u7_n94 ) );
  NOR2_X1 u1_u2_u7_U70 (.A2( u1_u2_X_48 ) , .A1( u1_u2_u7_n166 ) , .ZN( u1_u2_u7_n95 ) );
  NOR2_X1 u1_u2_u7_U71 (.A2( u1_u2_X_45 ) , .A1( u1_u2_X_48 ) , .ZN( u1_u2_u7_n99 ) );
  NOR2_X1 u1_u2_u7_U72 (.A2( u1_u2_X_44 ) , .A1( u1_u2_u7_n167 ) , .ZN( u1_u2_u7_n98 ) );
  NOR2_X1 u1_u2_u7_U73 (.A2( u1_u2_X_46 ) , .A1( u1_u2_X_47 ) , .ZN( u1_u2_u7_n152 ) );
  AND2_X1 u1_u2_u7_U74 (.A1( u1_u2_X_47 ) , .ZN( u1_u2_u7_n156 ) , .A2( u1_u2_u7_n163 ) );
  NAND2_X1 u1_u2_u7_U75 (.A2( u1_u2_X_46 ) , .A1( u1_u2_X_47 ) , .ZN( u1_u2_u7_n125 ) );
  AND2_X1 u1_u2_u7_U76 (.A2( u1_u2_X_45 ) , .A1( u1_u2_X_48 ) , .ZN( u1_u2_u7_n102 ) );
  AND2_X1 u1_u2_u7_U77 (.A2( u1_u2_X_43 ) , .A1( u1_u2_X_44 ) , .ZN( u1_u2_u7_n96 ) );
  AND2_X1 u1_u2_u7_U78 (.A1( u1_u2_X_44 ) , .ZN( u1_u2_u7_n100 ) , .A2( u1_u2_u7_n167 ) );
  AND2_X1 u1_u2_u7_U79 (.A1( u1_u2_X_48 ) , .A2( u1_u2_u7_n166 ) , .ZN( u1_u2_u7_n93 ) );
  OAI222_X1 u1_u2_u7_U8 (.C2( u1_u2_u7_n101 ) , .B2( u1_u2_u7_n111 ) , .A1( u1_u2_u7_n113 ) , .C1( u1_u2_u7_n146 ) , .A2( u1_u2_u7_n162 ) , .B1( u1_u2_u7_n164 ) , .ZN( u1_u2_u7_n94 ) );
  INV_X1 u1_u2_u7_U80 (.A( u1_u2_X_46 ) , .ZN( u1_u2_u7_n163 ) );
  INV_X1 u1_u2_u7_U81 (.A( u1_u2_X_43 ) , .ZN( u1_u2_u7_n167 ) );
  INV_X1 u1_u2_u7_U82 (.A( u1_u2_X_45 ) , .ZN( u1_u2_u7_n166 ) );
  NAND4_X1 u1_u2_u7_U83 (.ZN( u1_out2_5 ) , .A4( u1_u2_u7_n108 ) , .A3( u1_u2_u7_n109 ) , .A1( u1_u2_u7_n116 ) , .A2( u1_u2_u7_n123 ) );
  AOI22_X1 u1_u2_u7_U84 (.ZN( u1_u2_u7_n109 ) , .A2( u1_u2_u7_n126 ) , .B2( u1_u2_u7_n145 ) , .B1( u1_u2_u7_n156 ) , .A1( u1_u2_u7_n171 ) );
  NOR4_X1 u1_u2_u7_U85 (.A4( u1_u2_u7_n104 ) , .A3( u1_u2_u7_n105 ) , .A2( u1_u2_u7_n106 ) , .A1( u1_u2_u7_n107 ) , .ZN( u1_u2_u7_n108 ) );
  NAND4_X1 u1_u2_u7_U86 (.ZN( u1_out2_27 ) , .A4( u1_u2_u7_n118 ) , .A3( u1_u2_u7_n119 ) , .A2( u1_u2_u7_n120 ) , .A1( u1_u2_u7_n121 ) );
  OAI21_X1 u1_u2_u7_U87 (.ZN( u1_u2_u7_n121 ) , .B2( u1_u2_u7_n145 ) , .A( u1_u2_u7_n150 ) , .B1( u1_u2_u7_n174 ) );
  OAI21_X1 u1_u2_u7_U88 (.ZN( u1_u2_u7_n120 ) , .A( u1_u2_u7_n161 ) , .B2( u1_u2_u7_n170 ) , .B1( u1_u2_u7_n179 ) );
  NAND4_X1 u1_u2_u7_U89 (.ZN( u1_out2_21 ) , .A4( u1_u2_u7_n157 ) , .A3( u1_u2_u7_n158 ) , .A2( u1_u2_u7_n159 ) , .A1( u1_u2_u7_n160 ) );
  OAI221_X1 u1_u2_u7_U9 (.C1( u1_u2_u7_n101 ) , .C2( u1_u2_u7_n147 ) , .ZN( u1_u2_u7_n155 ) , .B2( u1_u2_u7_n162 ) , .A( u1_u2_u7_n91 ) , .B1( u1_u2_u7_n92 ) );
  OAI21_X1 u1_u2_u7_U90 (.B1( u1_u2_u7_n145 ) , .ZN( u1_u2_u7_n160 ) , .A( u1_u2_u7_n161 ) , .B2( u1_u2_u7_n177 ) );
  AOI22_X1 u1_u2_u7_U91 (.B2( u1_u2_u7_n149 ) , .B1( u1_u2_u7_n150 ) , .A2( u1_u2_u7_n151 ) , .A1( u1_u2_u7_n152 ) , .ZN( u1_u2_u7_n158 ) );
  NAND4_X1 u1_u2_u7_U92 (.ZN( u1_out2_15 ) , .A4( u1_u2_u7_n142 ) , .A3( u1_u2_u7_n143 ) , .A2( u1_u2_u7_n144 ) , .A1( u1_u2_u7_n178 ) );
  OR2_X1 u1_u2_u7_U93 (.A2( u1_u2_u7_n125 ) , .A1( u1_u2_u7_n129 ) , .ZN( u1_u2_u7_n144 ) );
  AOI22_X1 u1_u2_u7_U94 (.A2( u1_u2_u7_n126 ) , .ZN( u1_u2_u7_n143 ) , .B2( u1_u2_u7_n165 ) , .B1( u1_u2_u7_n173 ) , .A1( u1_u2_u7_n174 ) );
  NAND3_X1 u1_u2_u7_U95 (.A3( u1_u2_u7_n146 ) , .A2( u1_u2_u7_n147 ) , .A1( u1_u2_u7_n148 ) , .ZN( u1_u2_u7_n151 ) );
  NAND3_X1 u1_u2_u7_U96 (.A3( u1_u2_u7_n131 ) , .A2( u1_u2_u7_n132 ) , .A1( u1_u2_u7_n133 ) , .ZN( u1_u2_u7_n135 ) );
  XOR2_X1 u1_u3_U26 (.B( u1_K4_30 ) , .A( u1_R2_21 ) , .Z( u1_u3_X_30 ) );
  XOR2_X1 u1_u3_U28 (.B( u1_K4_29 ) , .A( u1_R2_20 ) , .Z( u1_u3_X_29 ) );
  XOR2_X1 u1_u3_U29 (.B( u1_K4_28 ) , .A( u1_R2_19 ) , .Z( u1_u3_X_28 ) );
  XOR2_X1 u1_u3_U30 (.B( u1_K4_27 ) , .A( u1_R2_18 ) , .Z( u1_u3_X_27 ) );
  XOR2_X1 u1_u3_U31 (.B( u1_K4_26 ) , .A( u1_R2_17 ) , .Z( u1_u3_X_26 ) );
  XOR2_X1 u1_u3_U32 (.B( u1_K4_25 ) , .A( u1_R2_16 ) , .Z( u1_u3_X_25 ) );
  OAI22_X1 u1_u3_u4_U10 (.B2( u1_u3_u4_n135 ) , .ZN( u1_u3_u4_n137 ) , .B1( u1_u3_u4_n153 ) , .A1( u1_u3_u4_n155 ) , .A2( u1_u3_u4_n171 ) );
  AND3_X1 u1_u3_u4_U11 (.A2( u1_u3_u4_n134 ) , .ZN( u1_u3_u4_n135 ) , .A3( u1_u3_u4_n145 ) , .A1( u1_u3_u4_n157 ) );
  NAND2_X1 u1_u3_u4_U12 (.ZN( u1_u3_u4_n132 ) , .A2( u1_u3_u4_n170 ) , .A1( u1_u3_u4_n173 ) );
  AOI21_X1 u1_u3_u4_U13 (.B2( u1_u3_u4_n160 ) , .B1( u1_u3_u4_n161 ) , .ZN( u1_u3_u4_n162 ) , .A( u1_u3_u4_n170 ) );
  AOI21_X1 u1_u3_u4_U14 (.ZN( u1_u3_u4_n107 ) , .B2( u1_u3_u4_n143 ) , .A( u1_u3_u4_n174 ) , .B1( u1_u3_u4_n184 ) );
  AOI21_X1 u1_u3_u4_U15 (.B2( u1_u3_u4_n158 ) , .B1( u1_u3_u4_n159 ) , .ZN( u1_u3_u4_n163 ) , .A( u1_u3_u4_n174 ) );
  AOI21_X1 u1_u3_u4_U16 (.A( u1_u3_u4_n153 ) , .B2( u1_u3_u4_n154 ) , .B1( u1_u3_u4_n155 ) , .ZN( u1_u3_u4_n165 ) );
  AOI21_X1 u1_u3_u4_U17 (.A( u1_u3_u4_n156 ) , .B2( u1_u3_u4_n157 ) , .ZN( u1_u3_u4_n164 ) , .B1( u1_u3_u4_n184 ) );
  INV_X1 u1_u3_u4_U18 (.A( u1_u3_u4_n138 ) , .ZN( u1_u3_u4_n170 ) );
  AND2_X1 u1_u3_u4_U19 (.A2( u1_u3_u4_n120 ) , .ZN( u1_u3_u4_n155 ) , .A1( u1_u3_u4_n160 ) );
  INV_X1 u1_u3_u4_U20 (.A( u1_u3_u4_n156 ) , .ZN( u1_u3_u4_n175 ) );
  NAND2_X1 u1_u3_u4_U21 (.A2( u1_u3_u4_n118 ) , .ZN( u1_u3_u4_n131 ) , .A1( u1_u3_u4_n147 ) );
  NAND2_X1 u1_u3_u4_U22 (.A1( u1_u3_u4_n119 ) , .A2( u1_u3_u4_n120 ) , .ZN( u1_u3_u4_n130 ) );
  NAND2_X1 u1_u3_u4_U23 (.ZN( u1_u3_u4_n117 ) , .A2( u1_u3_u4_n118 ) , .A1( u1_u3_u4_n148 ) );
  NAND2_X1 u1_u3_u4_U24 (.ZN( u1_u3_u4_n129 ) , .A1( u1_u3_u4_n134 ) , .A2( u1_u3_u4_n148 ) );
  AND3_X1 u1_u3_u4_U25 (.A1( u1_u3_u4_n119 ) , .A2( u1_u3_u4_n143 ) , .A3( u1_u3_u4_n154 ) , .ZN( u1_u3_u4_n161 ) );
  AND2_X1 u1_u3_u4_U26 (.A1( u1_u3_u4_n145 ) , .A2( u1_u3_u4_n147 ) , .ZN( u1_u3_u4_n159 ) );
  OR3_X1 u1_u3_u4_U27 (.A3( u1_u3_u4_n114 ) , .A2( u1_u3_u4_n115 ) , .A1( u1_u3_u4_n116 ) , .ZN( u1_u3_u4_n136 ) );
  AOI21_X1 u1_u3_u4_U28 (.A( u1_u3_u4_n113 ) , .ZN( u1_u3_u4_n116 ) , .B2( u1_u3_u4_n173 ) , .B1( u1_u3_u4_n174 ) );
  AOI21_X1 u1_u3_u4_U29 (.ZN( u1_u3_u4_n115 ) , .B2( u1_u3_u4_n145 ) , .B1( u1_u3_u4_n146 ) , .A( u1_u3_u4_n156 ) );
  NOR2_X1 u1_u3_u4_U3 (.ZN( u1_u3_u4_n121 ) , .A1( u1_u3_u4_n181 ) , .A2( u1_u3_u4_n182 ) );
  OAI22_X1 u1_u3_u4_U30 (.ZN( u1_u3_u4_n114 ) , .A2( u1_u3_u4_n121 ) , .B1( u1_u3_u4_n160 ) , .B2( u1_u3_u4_n170 ) , .A1( u1_u3_u4_n171 ) );
  INV_X1 u1_u3_u4_U31 (.A( u1_u3_u4_n158 ) , .ZN( u1_u3_u4_n182 ) );
  INV_X1 u1_u3_u4_U32 (.ZN( u1_u3_u4_n181 ) , .A( u1_u3_u4_n96 ) );
  INV_X1 u1_u3_u4_U33 (.A( u1_u3_u4_n144 ) , .ZN( u1_u3_u4_n179 ) );
  INV_X1 u1_u3_u4_U34 (.A( u1_u3_u4_n157 ) , .ZN( u1_u3_u4_n178 ) );
  NAND2_X1 u1_u3_u4_U35 (.A2( u1_u3_u4_n154 ) , .A1( u1_u3_u4_n96 ) , .ZN( u1_u3_u4_n97 ) );
  INV_X1 u1_u3_u4_U36 (.ZN( u1_u3_u4_n186 ) , .A( u1_u3_u4_n95 ) );
  OAI221_X1 u1_u3_u4_U37 (.C1( u1_u3_u4_n134 ) , .B1( u1_u3_u4_n158 ) , .B2( u1_u3_u4_n171 ) , .C2( u1_u3_u4_n173 ) , .A( u1_u3_u4_n94 ) , .ZN( u1_u3_u4_n95 ) );
  AOI222_X1 u1_u3_u4_U38 (.B2( u1_u3_u4_n132 ) , .A1( u1_u3_u4_n138 ) , .C2( u1_u3_u4_n175 ) , .A2( u1_u3_u4_n179 ) , .C1( u1_u3_u4_n181 ) , .B1( u1_u3_u4_n185 ) , .ZN( u1_u3_u4_n94 ) );
  INV_X1 u1_u3_u4_U39 (.A( u1_u3_u4_n113 ) , .ZN( u1_u3_u4_n185 ) );
  INV_X1 u1_u3_u4_U4 (.A( u1_u3_u4_n117 ) , .ZN( u1_u3_u4_n184 ) );
  INV_X1 u1_u3_u4_U40 (.A( u1_u3_u4_n143 ) , .ZN( u1_u3_u4_n183 ) );
  NOR2_X1 u1_u3_u4_U41 (.ZN( u1_u3_u4_n138 ) , .A1( u1_u3_u4_n168 ) , .A2( u1_u3_u4_n169 ) );
  NOR2_X1 u1_u3_u4_U42 (.A1( u1_u3_u4_n150 ) , .A2( u1_u3_u4_n152 ) , .ZN( u1_u3_u4_n153 ) );
  NOR2_X1 u1_u3_u4_U43 (.A2( u1_u3_u4_n128 ) , .A1( u1_u3_u4_n138 ) , .ZN( u1_u3_u4_n156 ) );
  AOI22_X1 u1_u3_u4_U44 (.B2( u1_u3_u4_n122 ) , .A1( u1_u3_u4_n123 ) , .ZN( u1_u3_u4_n124 ) , .B1( u1_u3_u4_n128 ) , .A2( u1_u3_u4_n172 ) );
  INV_X1 u1_u3_u4_U45 (.A( u1_u3_u4_n153 ) , .ZN( u1_u3_u4_n172 ) );
  NAND2_X1 u1_u3_u4_U46 (.A2( u1_u3_u4_n120 ) , .ZN( u1_u3_u4_n123 ) , .A1( u1_u3_u4_n161 ) );
  AOI22_X1 u1_u3_u4_U47 (.B2( u1_u3_u4_n132 ) , .A2( u1_u3_u4_n133 ) , .ZN( u1_u3_u4_n140 ) , .A1( u1_u3_u4_n150 ) , .B1( u1_u3_u4_n179 ) );
  NAND2_X1 u1_u3_u4_U48 (.ZN( u1_u3_u4_n133 ) , .A2( u1_u3_u4_n146 ) , .A1( u1_u3_u4_n154 ) );
  NAND2_X1 u1_u3_u4_U49 (.A1( u1_u3_u4_n103 ) , .ZN( u1_u3_u4_n154 ) , .A2( u1_u3_u4_n98 ) );
  NOR4_X1 u1_u3_u4_U5 (.A4( u1_u3_u4_n106 ) , .A3( u1_u3_u4_n107 ) , .A2( u1_u3_u4_n108 ) , .A1( u1_u3_u4_n109 ) , .ZN( u1_u3_u4_n110 ) );
  NAND2_X1 u1_u3_u4_U50 (.A1( u1_u3_u4_n101 ) , .ZN( u1_u3_u4_n158 ) , .A2( u1_u3_u4_n99 ) );
  AOI21_X1 u1_u3_u4_U51 (.ZN( u1_u3_u4_n127 ) , .A( u1_u3_u4_n136 ) , .B2( u1_u3_u4_n150 ) , .B1( u1_u3_u4_n180 ) );
  INV_X1 u1_u3_u4_U52 (.A( u1_u3_u4_n160 ) , .ZN( u1_u3_u4_n180 ) );
  NAND2_X1 u1_u3_u4_U53 (.A2( u1_u3_u4_n104 ) , .A1( u1_u3_u4_n105 ) , .ZN( u1_u3_u4_n146 ) );
  NAND2_X1 u1_u3_u4_U54 (.A2( u1_u3_u4_n101 ) , .A1( u1_u3_u4_n102 ) , .ZN( u1_u3_u4_n160 ) );
  NAND2_X1 u1_u3_u4_U55 (.ZN( u1_u3_u4_n134 ) , .A1( u1_u3_u4_n98 ) , .A2( u1_u3_u4_n99 ) );
  NAND2_X1 u1_u3_u4_U56 (.A1( u1_u3_u4_n103 ) , .A2( u1_u3_u4_n104 ) , .ZN( u1_u3_u4_n143 ) );
  NAND2_X1 u1_u3_u4_U57 (.A2( u1_u3_u4_n105 ) , .ZN( u1_u3_u4_n145 ) , .A1( u1_u3_u4_n98 ) );
  NAND2_X1 u1_u3_u4_U58 (.A1( u1_u3_u4_n100 ) , .A2( u1_u3_u4_n105 ) , .ZN( u1_u3_u4_n120 ) );
  NAND2_X1 u1_u3_u4_U59 (.A1( u1_u3_u4_n102 ) , .A2( u1_u3_u4_n104 ) , .ZN( u1_u3_u4_n148 ) );
  AOI21_X1 u1_u3_u4_U6 (.ZN( u1_u3_u4_n106 ) , .B2( u1_u3_u4_n146 ) , .B1( u1_u3_u4_n158 ) , .A( u1_u3_u4_n170 ) );
  NAND2_X1 u1_u3_u4_U60 (.A2( u1_u3_u4_n100 ) , .A1( u1_u3_u4_n103 ) , .ZN( u1_u3_u4_n157 ) );
  INV_X1 u1_u3_u4_U61 (.A( u1_u3_u4_n150 ) , .ZN( u1_u3_u4_n173 ) );
  INV_X1 u1_u3_u4_U62 (.A( u1_u3_u4_n152 ) , .ZN( u1_u3_u4_n171 ) );
  NAND2_X1 u1_u3_u4_U63 (.A1( u1_u3_u4_n100 ) , .ZN( u1_u3_u4_n118 ) , .A2( u1_u3_u4_n99 ) );
  NAND2_X1 u1_u3_u4_U64 (.A2( u1_u3_u4_n100 ) , .A1( u1_u3_u4_n102 ) , .ZN( u1_u3_u4_n144 ) );
  NAND2_X1 u1_u3_u4_U65 (.A2( u1_u3_u4_n101 ) , .A1( u1_u3_u4_n105 ) , .ZN( u1_u3_u4_n96 ) );
  INV_X1 u1_u3_u4_U66 (.A( u1_u3_u4_n128 ) , .ZN( u1_u3_u4_n174 ) );
  NAND2_X1 u1_u3_u4_U67 (.A2( u1_u3_u4_n102 ) , .ZN( u1_u3_u4_n119 ) , .A1( u1_u3_u4_n98 ) );
  NAND2_X1 u1_u3_u4_U68 (.A2( u1_u3_u4_n101 ) , .A1( u1_u3_u4_n103 ) , .ZN( u1_u3_u4_n147 ) );
  NAND2_X1 u1_u3_u4_U69 (.A2( u1_u3_u4_n104 ) , .ZN( u1_u3_u4_n113 ) , .A1( u1_u3_u4_n99 ) );
  AOI21_X1 u1_u3_u4_U7 (.ZN( u1_u3_u4_n109 ) , .A( u1_u3_u4_n153 ) , .B1( u1_u3_u4_n159 ) , .B2( u1_u3_u4_n184 ) );
  NOR2_X1 u1_u3_u4_U70 (.A2( u1_u3_X_28 ) , .ZN( u1_u3_u4_n150 ) , .A1( u1_u3_u4_n168 ) );
  NOR2_X1 u1_u3_u4_U71 (.A2( u1_u3_X_29 ) , .ZN( u1_u3_u4_n152 ) , .A1( u1_u3_u4_n169 ) );
  NOR2_X1 u1_u3_u4_U72 (.A2( u1_u3_X_30 ) , .ZN( u1_u3_u4_n105 ) , .A1( u1_u3_u4_n176 ) );
  NOR2_X1 u1_u3_u4_U73 (.A2( u1_u3_X_26 ) , .ZN( u1_u3_u4_n100 ) , .A1( u1_u3_u4_n177 ) );
  NOR2_X1 u1_u3_u4_U74 (.A2( u1_u3_X_28 ) , .A1( u1_u3_X_29 ) , .ZN( u1_u3_u4_n128 ) );
  NOR2_X1 u1_u3_u4_U75 (.A2( u1_u3_X_27 ) , .A1( u1_u3_X_30 ) , .ZN( u1_u3_u4_n102 ) );
  NOR2_X1 u1_u3_u4_U76 (.A2( u1_u3_X_25 ) , .A1( u1_u3_X_26 ) , .ZN( u1_u3_u4_n98 ) );
  AND2_X1 u1_u3_u4_U77 (.A2( u1_u3_X_25 ) , .A1( u1_u3_X_26 ) , .ZN( u1_u3_u4_n104 ) );
  AND2_X1 u1_u3_u4_U78 (.A1( u1_u3_X_30 ) , .A2( u1_u3_u4_n176 ) , .ZN( u1_u3_u4_n99 ) );
  AND2_X1 u1_u3_u4_U79 (.A1( u1_u3_X_26 ) , .ZN( u1_u3_u4_n101 ) , .A2( u1_u3_u4_n177 ) );
  AOI21_X1 u1_u3_u4_U8 (.ZN( u1_u3_u4_n108 ) , .B2( u1_u3_u4_n134 ) , .B1( u1_u3_u4_n155 ) , .A( u1_u3_u4_n156 ) );
  AND2_X1 u1_u3_u4_U80 (.A1( u1_u3_X_27 ) , .A2( u1_u3_X_30 ) , .ZN( u1_u3_u4_n103 ) );
  INV_X1 u1_u3_u4_U81 (.A( u1_u3_X_28 ) , .ZN( u1_u3_u4_n169 ) );
  INV_X1 u1_u3_u4_U82 (.A( u1_u3_X_29 ) , .ZN( u1_u3_u4_n168 ) );
  INV_X1 u1_u3_u4_U83 (.A( u1_u3_X_25 ) , .ZN( u1_u3_u4_n177 ) );
  INV_X1 u1_u3_u4_U84 (.A( u1_u3_X_27 ) , .ZN( u1_u3_u4_n176 ) );
  NAND4_X1 u1_u3_u4_U85 (.ZN( u1_out3_25 ) , .A4( u1_u3_u4_n139 ) , .A3( u1_u3_u4_n140 ) , .A2( u1_u3_u4_n141 ) , .A1( u1_u3_u4_n142 ) );
  OAI21_X1 u1_u3_u4_U86 (.A( u1_u3_u4_n128 ) , .B2( u1_u3_u4_n129 ) , .B1( u1_u3_u4_n130 ) , .ZN( u1_u3_u4_n142 ) );
  OAI21_X1 u1_u3_u4_U87 (.B2( u1_u3_u4_n131 ) , .ZN( u1_u3_u4_n141 ) , .A( u1_u3_u4_n175 ) , .B1( u1_u3_u4_n183 ) );
  NAND4_X1 u1_u3_u4_U88 (.ZN( u1_out3_14 ) , .A4( u1_u3_u4_n124 ) , .A3( u1_u3_u4_n125 ) , .A2( u1_u3_u4_n126 ) , .A1( u1_u3_u4_n127 ) );
  AOI22_X1 u1_u3_u4_U89 (.B2( u1_u3_u4_n117 ) , .ZN( u1_u3_u4_n126 ) , .A1( u1_u3_u4_n129 ) , .B1( u1_u3_u4_n152 ) , .A2( u1_u3_u4_n175 ) );
  AOI211_X1 u1_u3_u4_U9 (.B( u1_u3_u4_n136 ) , .A( u1_u3_u4_n137 ) , .C2( u1_u3_u4_n138 ) , .ZN( u1_u3_u4_n139 ) , .C1( u1_u3_u4_n182 ) );
  AOI22_X1 u1_u3_u4_U90 (.ZN( u1_u3_u4_n125 ) , .B2( u1_u3_u4_n131 ) , .A2( u1_u3_u4_n132 ) , .B1( u1_u3_u4_n138 ) , .A1( u1_u3_u4_n178 ) );
  NAND4_X1 u1_u3_u4_U91 (.ZN( u1_out3_8 ) , .A4( u1_u3_u4_n110 ) , .A3( u1_u3_u4_n111 ) , .A2( u1_u3_u4_n112 ) , .A1( u1_u3_u4_n186 ) );
  NAND2_X1 u1_u3_u4_U92 (.ZN( u1_u3_u4_n112 ) , .A2( u1_u3_u4_n130 ) , .A1( u1_u3_u4_n150 ) );
  AOI22_X1 u1_u3_u4_U93 (.ZN( u1_u3_u4_n111 ) , .B2( u1_u3_u4_n132 ) , .A1( u1_u3_u4_n152 ) , .B1( u1_u3_u4_n178 ) , .A2( u1_u3_u4_n97 ) );
  AOI22_X1 u1_u3_u4_U94 (.B2( u1_u3_u4_n149 ) , .B1( u1_u3_u4_n150 ) , .A2( u1_u3_u4_n151 ) , .A1( u1_u3_u4_n152 ) , .ZN( u1_u3_u4_n167 ) );
  NOR4_X1 u1_u3_u4_U95 (.A4( u1_u3_u4_n162 ) , .A3( u1_u3_u4_n163 ) , .A2( u1_u3_u4_n164 ) , .A1( u1_u3_u4_n165 ) , .ZN( u1_u3_u4_n166 ) );
  NAND3_X1 u1_u3_u4_U96 (.ZN( u1_out3_3 ) , .A3( u1_u3_u4_n166 ) , .A1( u1_u3_u4_n167 ) , .A2( u1_u3_u4_n186 ) );
  NAND3_X1 u1_u3_u4_U97 (.A3( u1_u3_u4_n146 ) , .A2( u1_u3_u4_n147 ) , .A1( u1_u3_u4_n148 ) , .ZN( u1_u3_u4_n149 ) );
  NAND3_X1 u1_u3_u4_U98 (.A3( u1_u3_u4_n143 ) , .A2( u1_u3_u4_n144 ) , .A1( u1_u3_u4_n145 ) , .ZN( u1_u3_u4_n151 ) );
  NAND3_X1 u1_u3_u4_U99 (.A3( u1_u3_u4_n121 ) , .ZN( u1_u3_u4_n122 ) , .A2( u1_u3_u4_n144 ) , .A1( u1_u3_u4_n154 ) );
  XOR2_X1 u1_u4_U33 (.B( u1_K5_24 ) , .A( u1_R3_17 ) , .Z( u1_u4_X_24 ) );
  XOR2_X1 u1_u4_U34 (.B( u1_K5_23 ) , .A( u1_R3_16 ) , .Z( u1_u4_X_23 ) );
  XOR2_X1 u1_u4_U35 (.B( u1_K5_22 ) , .A( u1_R3_15 ) , .Z( u1_u4_X_22 ) );
  XOR2_X1 u1_u4_U36 (.B( u1_K5_21 ) , .A( u1_R3_14 ) , .Z( u1_u4_X_21 ) );
  XOR2_X1 u1_u4_U37 (.B( u1_K5_20 ) , .A( u1_R3_13 ) , .Z( u1_u4_X_20 ) );
  XOR2_X1 u1_u4_U39 (.B( u1_K5_19 ) , .A( u1_R3_12 ) , .Z( u1_u4_X_19 ) );
  OAI22_X1 u1_u4_u3_U10 (.B1( u1_u4_u3_n113 ) , .A2( u1_u4_u3_n135 ) , .A1( u1_u4_u3_n150 ) , .B2( u1_u4_u3_n164 ) , .ZN( u1_u4_u3_n98 ) );
  OAI211_X1 u1_u4_u3_U11 (.B( u1_u4_u3_n106 ) , .ZN( u1_u4_u3_n119 ) , .C2( u1_u4_u3_n128 ) , .C1( u1_u4_u3_n167 ) , .A( u1_u4_u3_n181 ) );
  AOI221_X1 u1_u4_u3_U12 (.C1( u1_u4_u3_n105 ) , .ZN( u1_u4_u3_n106 ) , .A( u1_u4_u3_n131 ) , .B2( u1_u4_u3_n132 ) , .C2( u1_u4_u3_n133 ) , .B1( u1_u4_u3_n169 ) );
  INV_X1 u1_u4_u3_U13 (.ZN( u1_u4_u3_n181 ) , .A( u1_u4_u3_n98 ) );
  NAND2_X1 u1_u4_u3_U14 (.ZN( u1_u4_u3_n105 ) , .A2( u1_u4_u3_n130 ) , .A1( u1_u4_u3_n155 ) );
  AOI22_X1 u1_u4_u3_U15 (.B1( u1_u4_u3_n115 ) , .A2( u1_u4_u3_n116 ) , .ZN( u1_u4_u3_n123 ) , .B2( u1_u4_u3_n133 ) , .A1( u1_u4_u3_n169 ) );
  NAND2_X1 u1_u4_u3_U16 (.ZN( u1_u4_u3_n116 ) , .A2( u1_u4_u3_n151 ) , .A1( u1_u4_u3_n182 ) );
  NOR2_X1 u1_u4_u3_U17 (.ZN( u1_u4_u3_n126 ) , .A2( u1_u4_u3_n150 ) , .A1( u1_u4_u3_n164 ) );
  AOI21_X1 u1_u4_u3_U18 (.ZN( u1_u4_u3_n112 ) , .B2( u1_u4_u3_n146 ) , .B1( u1_u4_u3_n155 ) , .A( u1_u4_u3_n167 ) );
  NAND2_X1 u1_u4_u3_U19 (.A1( u1_u4_u3_n135 ) , .ZN( u1_u4_u3_n142 ) , .A2( u1_u4_u3_n164 ) );
  NAND2_X1 u1_u4_u3_U20 (.ZN( u1_u4_u3_n132 ) , .A2( u1_u4_u3_n152 ) , .A1( u1_u4_u3_n156 ) );
  AND2_X1 u1_u4_u3_U21 (.A2( u1_u4_u3_n113 ) , .A1( u1_u4_u3_n114 ) , .ZN( u1_u4_u3_n151 ) );
  INV_X1 u1_u4_u3_U22 (.A( u1_u4_u3_n133 ) , .ZN( u1_u4_u3_n165 ) );
  INV_X1 u1_u4_u3_U23 (.A( u1_u4_u3_n135 ) , .ZN( u1_u4_u3_n170 ) );
  NAND2_X1 u1_u4_u3_U24 (.A1( u1_u4_u3_n107 ) , .A2( u1_u4_u3_n108 ) , .ZN( u1_u4_u3_n140 ) );
  NAND2_X1 u1_u4_u3_U25 (.ZN( u1_u4_u3_n117 ) , .A1( u1_u4_u3_n124 ) , .A2( u1_u4_u3_n148 ) );
  NAND2_X1 u1_u4_u3_U26 (.ZN( u1_u4_u3_n143 ) , .A1( u1_u4_u3_n165 ) , .A2( u1_u4_u3_n167 ) );
  INV_X1 u1_u4_u3_U27 (.A( u1_u4_u3_n130 ) , .ZN( u1_u4_u3_n177 ) );
  INV_X1 u1_u4_u3_U28 (.A( u1_u4_u3_n128 ) , .ZN( u1_u4_u3_n176 ) );
  INV_X1 u1_u4_u3_U29 (.A( u1_u4_u3_n155 ) , .ZN( u1_u4_u3_n174 ) );
  INV_X1 u1_u4_u3_U3 (.A( u1_u4_u3_n129 ) , .ZN( u1_u4_u3_n183 ) );
  INV_X1 u1_u4_u3_U30 (.A( u1_u4_u3_n139 ) , .ZN( u1_u4_u3_n185 ) );
  NOR2_X1 u1_u4_u3_U31 (.ZN( u1_u4_u3_n135 ) , .A2( u1_u4_u3_n141 ) , .A1( u1_u4_u3_n169 ) );
  OAI222_X1 u1_u4_u3_U32 (.C2( u1_u4_u3_n107 ) , .A2( u1_u4_u3_n108 ) , .B1( u1_u4_u3_n135 ) , .ZN( u1_u4_u3_n138 ) , .B2( u1_u4_u3_n146 ) , .C1( u1_u4_u3_n154 ) , .A1( u1_u4_u3_n164 ) );
  NOR4_X1 u1_u4_u3_U33 (.A4( u1_u4_u3_n157 ) , .A3( u1_u4_u3_n158 ) , .A2( u1_u4_u3_n159 ) , .A1( u1_u4_u3_n160 ) , .ZN( u1_u4_u3_n161 ) );
  AOI21_X1 u1_u4_u3_U34 (.B2( u1_u4_u3_n152 ) , .B1( u1_u4_u3_n153 ) , .ZN( u1_u4_u3_n158 ) , .A( u1_u4_u3_n164 ) );
  AOI21_X1 u1_u4_u3_U35 (.A( u1_u4_u3_n149 ) , .B2( u1_u4_u3_n150 ) , .B1( u1_u4_u3_n151 ) , .ZN( u1_u4_u3_n159 ) );
  AOI21_X1 u1_u4_u3_U36 (.A( u1_u4_u3_n154 ) , .B2( u1_u4_u3_n155 ) , .B1( u1_u4_u3_n156 ) , .ZN( u1_u4_u3_n157 ) );
  AOI211_X1 u1_u4_u3_U37 (.ZN( u1_u4_u3_n109 ) , .A( u1_u4_u3_n119 ) , .C2( u1_u4_u3_n129 ) , .B( u1_u4_u3_n138 ) , .C1( u1_u4_u3_n141 ) );
  AOI211_X1 u1_u4_u3_U38 (.B( u1_u4_u3_n119 ) , .A( u1_u4_u3_n120 ) , .C2( u1_u4_u3_n121 ) , .ZN( u1_u4_u3_n122 ) , .C1( u1_u4_u3_n179 ) );
  INV_X1 u1_u4_u3_U39 (.A( u1_u4_u3_n156 ) , .ZN( u1_u4_u3_n179 ) );
  INV_X1 u1_u4_u3_U4 (.A( u1_u4_u3_n140 ) , .ZN( u1_u4_u3_n182 ) );
  OAI22_X1 u1_u4_u3_U40 (.B1( u1_u4_u3_n118 ) , .ZN( u1_u4_u3_n120 ) , .A1( u1_u4_u3_n135 ) , .B2( u1_u4_u3_n154 ) , .A2( u1_u4_u3_n178 ) );
  AND3_X1 u1_u4_u3_U41 (.ZN( u1_u4_u3_n118 ) , .A2( u1_u4_u3_n124 ) , .A1( u1_u4_u3_n144 ) , .A3( u1_u4_u3_n152 ) );
  INV_X1 u1_u4_u3_U42 (.A( u1_u4_u3_n121 ) , .ZN( u1_u4_u3_n164 ) );
  NAND2_X1 u1_u4_u3_U43 (.ZN( u1_u4_u3_n133 ) , .A1( u1_u4_u3_n154 ) , .A2( u1_u4_u3_n164 ) );
  OAI211_X1 u1_u4_u3_U44 (.B( u1_u4_u3_n127 ) , .ZN( u1_u4_u3_n139 ) , .C1( u1_u4_u3_n150 ) , .C2( u1_u4_u3_n154 ) , .A( u1_u4_u3_n184 ) );
  INV_X1 u1_u4_u3_U45 (.A( u1_u4_u3_n125 ) , .ZN( u1_u4_u3_n184 ) );
  AOI221_X1 u1_u4_u3_U46 (.A( u1_u4_u3_n126 ) , .ZN( u1_u4_u3_n127 ) , .C2( u1_u4_u3_n132 ) , .C1( u1_u4_u3_n169 ) , .B2( u1_u4_u3_n170 ) , .B1( u1_u4_u3_n174 ) );
  OAI22_X1 u1_u4_u3_U47 (.A1( u1_u4_u3_n124 ) , .ZN( u1_u4_u3_n125 ) , .B2( u1_u4_u3_n145 ) , .A2( u1_u4_u3_n165 ) , .B1( u1_u4_u3_n167 ) );
  NOR2_X1 u1_u4_u3_U48 (.A1( u1_u4_u3_n113 ) , .ZN( u1_u4_u3_n131 ) , .A2( u1_u4_u3_n154 ) );
  NAND2_X1 u1_u4_u3_U49 (.A1( u1_u4_u3_n103 ) , .ZN( u1_u4_u3_n150 ) , .A2( u1_u4_u3_n99 ) );
  INV_X1 u1_u4_u3_U5 (.A( u1_u4_u3_n117 ) , .ZN( u1_u4_u3_n178 ) );
  NAND2_X1 u1_u4_u3_U50 (.A2( u1_u4_u3_n102 ) , .ZN( u1_u4_u3_n155 ) , .A1( u1_u4_u3_n97 ) );
  INV_X1 u1_u4_u3_U51 (.A( u1_u4_u3_n141 ) , .ZN( u1_u4_u3_n167 ) );
  AOI21_X1 u1_u4_u3_U52 (.B2( u1_u4_u3_n114 ) , .B1( u1_u4_u3_n146 ) , .A( u1_u4_u3_n154 ) , .ZN( u1_u4_u3_n94 ) );
  AOI21_X1 u1_u4_u3_U53 (.ZN( u1_u4_u3_n110 ) , .B2( u1_u4_u3_n142 ) , .B1( u1_u4_u3_n186 ) , .A( u1_u4_u3_n95 ) );
  INV_X1 u1_u4_u3_U54 (.A( u1_u4_u3_n145 ) , .ZN( u1_u4_u3_n186 ) );
  AOI21_X1 u1_u4_u3_U55 (.B1( u1_u4_u3_n124 ) , .A( u1_u4_u3_n149 ) , .B2( u1_u4_u3_n155 ) , .ZN( u1_u4_u3_n95 ) );
  INV_X1 u1_u4_u3_U56 (.A( u1_u4_u3_n149 ) , .ZN( u1_u4_u3_n169 ) );
  NAND2_X1 u1_u4_u3_U57 (.ZN( u1_u4_u3_n124 ) , .A1( u1_u4_u3_n96 ) , .A2( u1_u4_u3_n97 ) );
  NAND2_X1 u1_u4_u3_U58 (.A2( u1_u4_u3_n100 ) , .ZN( u1_u4_u3_n146 ) , .A1( u1_u4_u3_n96 ) );
  NAND2_X1 u1_u4_u3_U59 (.A1( u1_u4_u3_n101 ) , .ZN( u1_u4_u3_n145 ) , .A2( u1_u4_u3_n99 ) );
  AOI221_X1 u1_u4_u3_U6 (.A( u1_u4_u3_n131 ) , .C2( u1_u4_u3_n132 ) , .C1( u1_u4_u3_n133 ) , .ZN( u1_u4_u3_n134 ) , .B1( u1_u4_u3_n143 ) , .B2( u1_u4_u3_n177 ) );
  NAND2_X1 u1_u4_u3_U60 (.A1( u1_u4_u3_n100 ) , .ZN( u1_u4_u3_n156 ) , .A2( u1_u4_u3_n99 ) );
  NAND2_X1 u1_u4_u3_U61 (.A2( u1_u4_u3_n101 ) , .A1( u1_u4_u3_n104 ) , .ZN( u1_u4_u3_n148 ) );
  NAND2_X1 u1_u4_u3_U62 (.A1( u1_u4_u3_n100 ) , .A2( u1_u4_u3_n102 ) , .ZN( u1_u4_u3_n128 ) );
  NAND2_X1 u1_u4_u3_U63 (.A2( u1_u4_u3_n101 ) , .A1( u1_u4_u3_n102 ) , .ZN( u1_u4_u3_n152 ) );
  NAND2_X1 u1_u4_u3_U64 (.A2( u1_u4_u3_n101 ) , .ZN( u1_u4_u3_n114 ) , .A1( u1_u4_u3_n96 ) );
  NAND2_X1 u1_u4_u3_U65 (.ZN( u1_u4_u3_n107 ) , .A1( u1_u4_u3_n97 ) , .A2( u1_u4_u3_n99 ) );
  NAND2_X1 u1_u4_u3_U66 (.A2( u1_u4_u3_n100 ) , .A1( u1_u4_u3_n104 ) , .ZN( u1_u4_u3_n113 ) );
  NAND2_X1 u1_u4_u3_U67 (.A1( u1_u4_u3_n104 ) , .ZN( u1_u4_u3_n153 ) , .A2( u1_u4_u3_n97 ) );
  NAND2_X1 u1_u4_u3_U68 (.A2( u1_u4_u3_n103 ) , .A1( u1_u4_u3_n104 ) , .ZN( u1_u4_u3_n130 ) );
  NAND2_X1 u1_u4_u3_U69 (.A2( u1_u4_u3_n103 ) , .ZN( u1_u4_u3_n144 ) , .A1( u1_u4_u3_n96 ) );
  OAI22_X1 u1_u4_u3_U7 (.B2( u1_u4_u3_n147 ) , .A2( u1_u4_u3_n148 ) , .ZN( u1_u4_u3_n160 ) , .B1( u1_u4_u3_n165 ) , .A1( u1_u4_u3_n168 ) );
  NAND2_X1 u1_u4_u3_U70 (.A1( u1_u4_u3_n102 ) , .A2( u1_u4_u3_n103 ) , .ZN( u1_u4_u3_n108 ) );
  NOR2_X1 u1_u4_u3_U71 (.A2( u1_u4_X_19 ) , .A1( u1_u4_X_20 ) , .ZN( u1_u4_u3_n99 ) );
  NOR2_X1 u1_u4_u3_U72 (.A2( u1_u4_X_21 ) , .A1( u1_u4_X_24 ) , .ZN( u1_u4_u3_n103 ) );
  NOR2_X1 u1_u4_u3_U73 (.A2( u1_u4_X_24 ) , .A1( u1_u4_u3_n171 ) , .ZN( u1_u4_u3_n97 ) );
  NOR2_X1 u1_u4_u3_U74 (.A2( u1_u4_X_23 ) , .ZN( u1_u4_u3_n141 ) , .A1( u1_u4_u3_n166 ) );
  NOR2_X1 u1_u4_u3_U75 (.A2( u1_u4_X_19 ) , .A1( u1_u4_u3_n172 ) , .ZN( u1_u4_u3_n96 ) );
  NAND2_X1 u1_u4_u3_U76 (.A1( u1_u4_X_22 ) , .A2( u1_u4_X_23 ) , .ZN( u1_u4_u3_n154 ) );
  NAND2_X1 u1_u4_u3_U77 (.A1( u1_u4_X_23 ) , .ZN( u1_u4_u3_n149 ) , .A2( u1_u4_u3_n166 ) );
  NOR2_X1 u1_u4_u3_U78 (.A2( u1_u4_X_22 ) , .A1( u1_u4_X_23 ) , .ZN( u1_u4_u3_n121 ) );
  AND2_X1 u1_u4_u3_U79 (.A1( u1_u4_X_24 ) , .ZN( u1_u4_u3_n101 ) , .A2( u1_u4_u3_n171 ) );
  AND3_X1 u1_u4_u3_U8 (.A3( u1_u4_u3_n144 ) , .A2( u1_u4_u3_n145 ) , .A1( u1_u4_u3_n146 ) , .ZN( u1_u4_u3_n147 ) );
  AND2_X1 u1_u4_u3_U80 (.A1( u1_u4_X_19 ) , .ZN( u1_u4_u3_n102 ) , .A2( u1_u4_u3_n172 ) );
  AND2_X1 u1_u4_u3_U81 (.A1( u1_u4_X_21 ) , .A2( u1_u4_X_24 ) , .ZN( u1_u4_u3_n100 ) );
  AND2_X1 u1_u4_u3_U82 (.A2( u1_u4_X_19 ) , .A1( u1_u4_X_20 ) , .ZN( u1_u4_u3_n104 ) );
  INV_X1 u1_u4_u3_U83 (.A( u1_u4_X_22 ) , .ZN( u1_u4_u3_n166 ) );
  INV_X1 u1_u4_u3_U84 (.A( u1_u4_X_21 ) , .ZN( u1_u4_u3_n171 ) );
  INV_X1 u1_u4_u3_U85 (.A( u1_u4_X_20 ) , .ZN( u1_u4_u3_n172 ) );
  NAND4_X1 u1_u4_u3_U86 (.ZN( u1_out4_26 ) , .A4( u1_u4_u3_n109 ) , .A3( u1_u4_u3_n110 ) , .A2( u1_u4_u3_n111 ) , .A1( u1_u4_u3_n173 ) );
  INV_X1 u1_u4_u3_U87 (.ZN( u1_u4_u3_n173 ) , .A( u1_u4_u3_n94 ) );
  OAI21_X1 u1_u4_u3_U88 (.ZN( u1_u4_u3_n111 ) , .B2( u1_u4_u3_n117 ) , .A( u1_u4_u3_n133 ) , .B1( u1_u4_u3_n176 ) );
  NAND4_X1 u1_u4_u3_U89 (.ZN( u1_out4_20 ) , .A4( u1_u4_u3_n122 ) , .A3( u1_u4_u3_n123 ) , .A1( u1_u4_u3_n175 ) , .A2( u1_u4_u3_n180 ) );
  INV_X1 u1_u4_u3_U9 (.A( u1_u4_u3_n143 ) , .ZN( u1_u4_u3_n168 ) );
  INV_X1 u1_u4_u3_U90 (.A( u1_u4_u3_n126 ) , .ZN( u1_u4_u3_n180 ) );
  INV_X1 u1_u4_u3_U91 (.A( u1_u4_u3_n112 ) , .ZN( u1_u4_u3_n175 ) );
  NAND4_X1 u1_u4_u3_U92 (.ZN( u1_out4_1 ) , .A4( u1_u4_u3_n161 ) , .A3( u1_u4_u3_n162 ) , .A2( u1_u4_u3_n163 ) , .A1( u1_u4_u3_n185 ) );
  NAND2_X1 u1_u4_u3_U93 (.ZN( u1_u4_u3_n163 ) , .A2( u1_u4_u3_n170 ) , .A1( u1_u4_u3_n176 ) );
  AOI22_X1 u1_u4_u3_U94 (.B2( u1_u4_u3_n140 ) , .B1( u1_u4_u3_n141 ) , .A2( u1_u4_u3_n142 ) , .ZN( u1_u4_u3_n162 ) , .A1( u1_u4_u3_n177 ) );
  OR4_X1 u1_u4_u3_U95 (.ZN( u1_out4_10 ) , .A4( u1_u4_u3_n136 ) , .A3( u1_u4_u3_n137 ) , .A1( u1_u4_u3_n138 ) , .A2( u1_u4_u3_n139 ) );
  OAI222_X1 u1_u4_u3_U96 (.C1( u1_u4_u3_n128 ) , .ZN( u1_u4_u3_n137 ) , .B1( u1_u4_u3_n148 ) , .A2( u1_u4_u3_n150 ) , .B2( u1_u4_u3_n154 ) , .C2( u1_u4_u3_n164 ) , .A1( u1_u4_u3_n167 ) );
  OAI221_X1 u1_u4_u3_U97 (.A( u1_u4_u3_n134 ) , .B2( u1_u4_u3_n135 ) , .ZN( u1_u4_u3_n136 ) , .C1( u1_u4_u3_n149 ) , .B1( u1_u4_u3_n151 ) , .C2( u1_u4_u3_n183 ) );
  NAND3_X1 u1_u4_u3_U98 (.A1( u1_u4_u3_n114 ) , .ZN( u1_u4_u3_n115 ) , .A2( u1_u4_u3_n145 ) , .A3( u1_u4_u3_n153 ) );
  NAND3_X1 u1_u4_u3_U99 (.ZN( u1_u4_u3_n129 ) , .A2( u1_u4_u3_n144 ) , .A1( u1_u4_u3_n153 ) , .A3( u1_u4_u3_n182 ) );
  XOR2_X1 u1_u7_U33 (.B( u1_K8_24 ) , .A( u1_R6_17 ) , .Z( u1_u7_X_24 ) );
  XOR2_X1 u1_u7_U34 (.B( u1_K8_23 ) , .A( u1_R6_16 ) , .Z( u1_u7_X_23 ) );
  XOR2_X1 u1_u7_U35 (.B( u1_K8_22 ) , .A( u1_R6_15 ) , .Z( u1_u7_X_22 ) );
  XOR2_X1 u1_u7_U36 (.B( u1_K8_21 ) , .A( u1_R6_14 ) , .Z( u1_u7_X_21 ) );
  XOR2_X1 u1_u7_U37 (.B( u1_K8_20 ) , .A( u1_R6_13 ) , .Z( u1_u7_X_20 ) );
  XOR2_X1 u1_u7_U39 (.B( u1_K8_19 ) , .A( u1_R6_12 ) , .Z( u1_u7_X_19 ) );
  OAI22_X1 u1_u7_u3_U10 (.B1( u1_u7_u3_n113 ) , .A2( u1_u7_u3_n135 ) , .A1( u1_u7_u3_n150 ) , .B2( u1_u7_u3_n164 ) , .ZN( u1_u7_u3_n98 ) );
  OAI211_X1 u1_u7_u3_U11 (.B( u1_u7_u3_n106 ) , .ZN( u1_u7_u3_n119 ) , .C2( u1_u7_u3_n128 ) , .C1( u1_u7_u3_n167 ) , .A( u1_u7_u3_n181 ) );
  AOI221_X1 u1_u7_u3_U12 (.C1( u1_u7_u3_n105 ) , .ZN( u1_u7_u3_n106 ) , .A( u1_u7_u3_n131 ) , .B2( u1_u7_u3_n132 ) , .C2( u1_u7_u3_n133 ) , .B1( u1_u7_u3_n169 ) );
  INV_X1 u1_u7_u3_U13 (.ZN( u1_u7_u3_n181 ) , .A( u1_u7_u3_n98 ) );
  NAND2_X1 u1_u7_u3_U14 (.ZN( u1_u7_u3_n105 ) , .A2( u1_u7_u3_n130 ) , .A1( u1_u7_u3_n155 ) );
  AOI22_X1 u1_u7_u3_U15 (.B1( u1_u7_u3_n115 ) , .A2( u1_u7_u3_n116 ) , .ZN( u1_u7_u3_n123 ) , .B2( u1_u7_u3_n133 ) , .A1( u1_u7_u3_n169 ) );
  NAND2_X1 u1_u7_u3_U16 (.ZN( u1_u7_u3_n116 ) , .A2( u1_u7_u3_n151 ) , .A1( u1_u7_u3_n182 ) );
  NOR2_X1 u1_u7_u3_U17 (.ZN( u1_u7_u3_n126 ) , .A2( u1_u7_u3_n150 ) , .A1( u1_u7_u3_n164 ) );
  AOI21_X1 u1_u7_u3_U18 (.ZN( u1_u7_u3_n112 ) , .B2( u1_u7_u3_n146 ) , .B1( u1_u7_u3_n155 ) , .A( u1_u7_u3_n167 ) );
  NAND2_X1 u1_u7_u3_U19 (.A1( u1_u7_u3_n135 ) , .ZN( u1_u7_u3_n142 ) , .A2( u1_u7_u3_n164 ) );
  NAND2_X1 u1_u7_u3_U20 (.ZN( u1_u7_u3_n132 ) , .A2( u1_u7_u3_n152 ) , .A1( u1_u7_u3_n156 ) );
  AND2_X1 u1_u7_u3_U21 (.A2( u1_u7_u3_n113 ) , .A1( u1_u7_u3_n114 ) , .ZN( u1_u7_u3_n151 ) );
  INV_X1 u1_u7_u3_U22 (.A( u1_u7_u3_n133 ) , .ZN( u1_u7_u3_n165 ) );
  INV_X1 u1_u7_u3_U23 (.A( u1_u7_u3_n135 ) , .ZN( u1_u7_u3_n170 ) );
  NAND2_X1 u1_u7_u3_U24 (.A1( u1_u7_u3_n107 ) , .A2( u1_u7_u3_n108 ) , .ZN( u1_u7_u3_n140 ) );
  NAND2_X1 u1_u7_u3_U25 (.ZN( u1_u7_u3_n117 ) , .A1( u1_u7_u3_n124 ) , .A2( u1_u7_u3_n148 ) );
  NAND2_X1 u1_u7_u3_U26 (.ZN( u1_u7_u3_n143 ) , .A1( u1_u7_u3_n165 ) , .A2( u1_u7_u3_n167 ) );
  INV_X1 u1_u7_u3_U27 (.A( u1_u7_u3_n130 ) , .ZN( u1_u7_u3_n177 ) );
  INV_X1 u1_u7_u3_U28 (.A( u1_u7_u3_n128 ) , .ZN( u1_u7_u3_n176 ) );
  INV_X1 u1_u7_u3_U29 (.A( u1_u7_u3_n155 ) , .ZN( u1_u7_u3_n174 ) );
  INV_X1 u1_u7_u3_U3 (.A( u1_u7_u3_n129 ) , .ZN( u1_u7_u3_n183 ) );
  INV_X1 u1_u7_u3_U30 (.A( u1_u7_u3_n139 ) , .ZN( u1_u7_u3_n185 ) );
  NOR2_X1 u1_u7_u3_U31 (.ZN( u1_u7_u3_n135 ) , .A2( u1_u7_u3_n141 ) , .A1( u1_u7_u3_n169 ) );
  OAI222_X1 u1_u7_u3_U32 (.C2( u1_u7_u3_n107 ) , .A2( u1_u7_u3_n108 ) , .B1( u1_u7_u3_n135 ) , .ZN( u1_u7_u3_n138 ) , .B2( u1_u7_u3_n146 ) , .C1( u1_u7_u3_n154 ) , .A1( u1_u7_u3_n164 ) );
  NOR4_X1 u1_u7_u3_U33 (.A4( u1_u7_u3_n157 ) , .A3( u1_u7_u3_n158 ) , .A2( u1_u7_u3_n159 ) , .A1( u1_u7_u3_n160 ) , .ZN( u1_u7_u3_n161 ) );
  AOI21_X1 u1_u7_u3_U34 (.B2( u1_u7_u3_n152 ) , .B1( u1_u7_u3_n153 ) , .ZN( u1_u7_u3_n158 ) , .A( u1_u7_u3_n164 ) );
  AOI21_X1 u1_u7_u3_U35 (.A( u1_u7_u3_n154 ) , .B2( u1_u7_u3_n155 ) , .B1( u1_u7_u3_n156 ) , .ZN( u1_u7_u3_n157 ) );
  AOI21_X1 u1_u7_u3_U36 (.A( u1_u7_u3_n149 ) , .B2( u1_u7_u3_n150 ) , .B1( u1_u7_u3_n151 ) , .ZN( u1_u7_u3_n159 ) );
  AOI211_X1 u1_u7_u3_U37 (.ZN( u1_u7_u3_n109 ) , .A( u1_u7_u3_n119 ) , .C2( u1_u7_u3_n129 ) , .B( u1_u7_u3_n138 ) , .C1( u1_u7_u3_n141 ) );
  AOI211_X1 u1_u7_u3_U38 (.B( u1_u7_u3_n119 ) , .A( u1_u7_u3_n120 ) , .C2( u1_u7_u3_n121 ) , .ZN( u1_u7_u3_n122 ) , .C1( u1_u7_u3_n179 ) );
  INV_X1 u1_u7_u3_U39 (.A( u1_u7_u3_n156 ) , .ZN( u1_u7_u3_n179 ) );
  INV_X1 u1_u7_u3_U4 (.A( u1_u7_u3_n140 ) , .ZN( u1_u7_u3_n182 ) );
  OAI22_X1 u1_u7_u3_U40 (.B1( u1_u7_u3_n118 ) , .ZN( u1_u7_u3_n120 ) , .A1( u1_u7_u3_n135 ) , .B2( u1_u7_u3_n154 ) , .A2( u1_u7_u3_n178 ) );
  AND3_X1 u1_u7_u3_U41 (.ZN( u1_u7_u3_n118 ) , .A2( u1_u7_u3_n124 ) , .A1( u1_u7_u3_n144 ) , .A3( u1_u7_u3_n152 ) );
  INV_X1 u1_u7_u3_U42 (.A( u1_u7_u3_n121 ) , .ZN( u1_u7_u3_n164 ) );
  NAND2_X1 u1_u7_u3_U43 (.ZN( u1_u7_u3_n133 ) , .A1( u1_u7_u3_n154 ) , .A2( u1_u7_u3_n164 ) );
  OAI211_X1 u1_u7_u3_U44 (.B( u1_u7_u3_n127 ) , .ZN( u1_u7_u3_n139 ) , .C1( u1_u7_u3_n150 ) , .C2( u1_u7_u3_n154 ) , .A( u1_u7_u3_n184 ) );
  INV_X1 u1_u7_u3_U45 (.A( u1_u7_u3_n125 ) , .ZN( u1_u7_u3_n184 ) );
  AOI221_X1 u1_u7_u3_U46 (.A( u1_u7_u3_n126 ) , .ZN( u1_u7_u3_n127 ) , .C2( u1_u7_u3_n132 ) , .C1( u1_u7_u3_n169 ) , .B2( u1_u7_u3_n170 ) , .B1( u1_u7_u3_n174 ) );
  OAI22_X1 u1_u7_u3_U47 (.A1( u1_u7_u3_n124 ) , .ZN( u1_u7_u3_n125 ) , .B2( u1_u7_u3_n145 ) , .A2( u1_u7_u3_n165 ) , .B1( u1_u7_u3_n167 ) );
  NOR2_X1 u1_u7_u3_U48 (.A1( u1_u7_u3_n113 ) , .ZN( u1_u7_u3_n131 ) , .A2( u1_u7_u3_n154 ) );
  NAND2_X1 u1_u7_u3_U49 (.A1( u1_u7_u3_n103 ) , .ZN( u1_u7_u3_n150 ) , .A2( u1_u7_u3_n99 ) );
  INV_X1 u1_u7_u3_U5 (.A( u1_u7_u3_n117 ) , .ZN( u1_u7_u3_n178 ) );
  NAND2_X1 u1_u7_u3_U50 (.A2( u1_u7_u3_n102 ) , .ZN( u1_u7_u3_n155 ) , .A1( u1_u7_u3_n97 ) );
  INV_X1 u1_u7_u3_U51 (.A( u1_u7_u3_n141 ) , .ZN( u1_u7_u3_n167 ) );
  AOI21_X1 u1_u7_u3_U52 (.B2( u1_u7_u3_n114 ) , .B1( u1_u7_u3_n146 ) , .A( u1_u7_u3_n154 ) , .ZN( u1_u7_u3_n94 ) );
  AOI21_X1 u1_u7_u3_U53 (.ZN( u1_u7_u3_n110 ) , .B2( u1_u7_u3_n142 ) , .B1( u1_u7_u3_n186 ) , .A( u1_u7_u3_n95 ) );
  INV_X1 u1_u7_u3_U54 (.A( u1_u7_u3_n145 ) , .ZN( u1_u7_u3_n186 ) );
  AOI21_X1 u1_u7_u3_U55 (.B1( u1_u7_u3_n124 ) , .A( u1_u7_u3_n149 ) , .B2( u1_u7_u3_n155 ) , .ZN( u1_u7_u3_n95 ) );
  INV_X1 u1_u7_u3_U56 (.A( u1_u7_u3_n149 ) , .ZN( u1_u7_u3_n169 ) );
  NAND2_X1 u1_u7_u3_U57 (.ZN( u1_u7_u3_n124 ) , .A1( u1_u7_u3_n96 ) , .A2( u1_u7_u3_n97 ) );
  NAND2_X1 u1_u7_u3_U58 (.A2( u1_u7_u3_n100 ) , .ZN( u1_u7_u3_n146 ) , .A1( u1_u7_u3_n96 ) );
  NAND2_X1 u1_u7_u3_U59 (.A1( u1_u7_u3_n101 ) , .ZN( u1_u7_u3_n145 ) , .A2( u1_u7_u3_n99 ) );
  AOI221_X1 u1_u7_u3_U6 (.A( u1_u7_u3_n131 ) , .C2( u1_u7_u3_n132 ) , .C1( u1_u7_u3_n133 ) , .ZN( u1_u7_u3_n134 ) , .B1( u1_u7_u3_n143 ) , .B2( u1_u7_u3_n177 ) );
  NAND2_X1 u1_u7_u3_U60 (.A1( u1_u7_u3_n100 ) , .ZN( u1_u7_u3_n156 ) , .A2( u1_u7_u3_n99 ) );
  NAND2_X1 u1_u7_u3_U61 (.A2( u1_u7_u3_n101 ) , .A1( u1_u7_u3_n104 ) , .ZN( u1_u7_u3_n148 ) );
  NAND2_X1 u1_u7_u3_U62 (.A1( u1_u7_u3_n100 ) , .A2( u1_u7_u3_n102 ) , .ZN( u1_u7_u3_n128 ) );
  NAND2_X1 u1_u7_u3_U63 (.A2( u1_u7_u3_n101 ) , .A1( u1_u7_u3_n102 ) , .ZN( u1_u7_u3_n152 ) );
  NAND2_X1 u1_u7_u3_U64 (.A2( u1_u7_u3_n101 ) , .ZN( u1_u7_u3_n114 ) , .A1( u1_u7_u3_n96 ) );
  NAND2_X1 u1_u7_u3_U65 (.ZN( u1_u7_u3_n107 ) , .A1( u1_u7_u3_n97 ) , .A2( u1_u7_u3_n99 ) );
  NAND2_X1 u1_u7_u3_U66 (.A2( u1_u7_u3_n100 ) , .A1( u1_u7_u3_n104 ) , .ZN( u1_u7_u3_n113 ) );
  NAND2_X1 u1_u7_u3_U67 (.A1( u1_u7_u3_n104 ) , .ZN( u1_u7_u3_n153 ) , .A2( u1_u7_u3_n97 ) );
  NAND2_X1 u1_u7_u3_U68 (.A2( u1_u7_u3_n103 ) , .A1( u1_u7_u3_n104 ) , .ZN( u1_u7_u3_n130 ) );
  NAND2_X1 u1_u7_u3_U69 (.A2( u1_u7_u3_n103 ) , .ZN( u1_u7_u3_n144 ) , .A1( u1_u7_u3_n96 ) );
  OAI22_X1 u1_u7_u3_U7 (.B2( u1_u7_u3_n147 ) , .A2( u1_u7_u3_n148 ) , .ZN( u1_u7_u3_n160 ) , .B1( u1_u7_u3_n165 ) , .A1( u1_u7_u3_n168 ) );
  NAND2_X1 u1_u7_u3_U70 (.A1( u1_u7_u3_n102 ) , .A2( u1_u7_u3_n103 ) , .ZN( u1_u7_u3_n108 ) );
  NOR2_X1 u1_u7_u3_U71 (.A2( u1_u7_X_19 ) , .A1( u1_u7_X_20 ) , .ZN( u1_u7_u3_n99 ) );
  NOR2_X1 u1_u7_u3_U72 (.A2( u1_u7_X_21 ) , .A1( u1_u7_X_24 ) , .ZN( u1_u7_u3_n103 ) );
  NOR2_X1 u1_u7_u3_U73 (.A2( u1_u7_X_24 ) , .A1( u1_u7_u3_n171 ) , .ZN( u1_u7_u3_n97 ) );
  NOR2_X1 u1_u7_u3_U74 (.A2( u1_u7_X_23 ) , .ZN( u1_u7_u3_n141 ) , .A1( u1_u7_u3_n166 ) );
  NOR2_X1 u1_u7_u3_U75 (.A2( u1_u7_X_19 ) , .A1( u1_u7_u3_n172 ) , .ZN( u1_u7_u3_n96 ) );
  NAND2_X1 u1_u7_u3_U76 (.A1( u1_u7_X_22 ) , .A2( u1_u7_X_23 ) , .ZN( u1_u7_u3_n154 ) );
  NAND2_X1 u1_u7_u3_U77 (.A1( u1_u7_X_23 ) , .ZN( u1_u7_u3_n149 ) , .A2( u1_u7_u3_n166 ) );
  NOR2_X1 u1_u7_u3_U78 (.A2( u1_u7_X_22 ) , .A1( u1_u7_X_23 ) , .ZN( u1_u7_u3_n121 ) );
  AND2_X1 u1_u7_u3_U79 (.A1( u1_u7_X_24 ) , .ZN( u1_u7_u3_n101 ) , .A2( u1_u7_u3_n171 ) );
  AND3_X1 u1_u7_u3_U8 (.A3( u1_u7_u3_n144 ) , .A2( u1_u7_u3_n145 ) , .A1( u1_u7_u3_n146 ) , .ZN( u1_u7_u3_n147 ) );
  AND2_X1 u1_u7_u3_U80 (.A1( u1_u7_X_19 ) , .ZN( u1_u7_u3_n102 ) , .A2( u1_u7_u3_n172 ) );
  AND2_X1 u1_u7_u3_U81 (.A1( u1_u7_X_21 ) , .A2( u1_u7_X_24 ) , .ZN( u1_u7_u3_n100 ) );
  AND2_X1 u1_u7_u3_U82 (.A2( u1_u7_X_19 ) , .A1( u1_u7_X_20 ) , .ZN( u1_u7_u3_n104 ) );
  INV_X1 u1_u7_u3_U83 (.A( u1_u7_X_22 ) , .ZN( u1_u7_u3_n166 ) );
  INV_X1 u1_u7_u3_U84 (.A( u1_u7_X_21 ) , .ZN( u1_u7_u3_n171 ) );
  INV_X1 u1_u7_u3_U85 (.A( u1_u7_X_20 ) , .ZN( u1_u7_u3_n172 ) );
  OR4_X1 u1_u7_u3_U86 (.ZN( u1_out7_10 ) , .A4( u1_u7_u3_n136 ) , .A3( u1_u7_u3_n137 ) , .A1( u1_u7_u3_n138 ) , .A2( u1_u7_u3_n139 ) );
  OAI222_X1 u1_u7_u3_U87 (.C1( u1_u7_u3_n128 ) , .ZN( u1_u7_u3_n137 ) , .B1( u1_u7_u3_n148 ) , .A2( u1_u7_u3_n150 ) , .B2( u1_u7_u3_n154 ) , .C2( u1_u7_u3_n164 ) , .A1( u1_u7_u3_n167 ) );
  OAI221_X1 u1_u7_u3_U88 (.A( u1_u7_u3_n134 ) , .B2( u1_u7_u3_n135 ) , .ZN( u1_u7_u3_n136 ) , .C1( u1_u7_u3_n149 ) , .B1( u1_u7_u3_n151 ) , .C2( u1_u7_u3_n183 ) );
  NAND4_X1 u1_u7_u3_U89 (.ZN( u1_out7_26 ) , .A4( u1_u7_u3_n109 ) , .A3( u1_u7_u3_n110 ) , .A2( u1_u7_u3_n111 ) , .A1( u1_u7_u3_n173 ) );
  INV_X1 u1_u7_u3_U9 (.A( u1_u7_u3_n143 ) , .ZN( u1_u7_u3_n168 ) );
  INV_X1 u1_u7_u3_U90 (.ZN( u1_u7_u3_n173 ) , .A( u1_u7_u3_n94 ) );
  OAI21_X1 u1_u7_u3_U91 (.ZN( u1_u7_u3_n111 ) , .B2( u1_u7_u3_n117 ) , .A( u1_u7_u3_n133 ) , .B1( u1_u7_u3_n176 ) );
  NAND4_X1 u1_u7_u3_U92 (.ZN( u1_out7_20 ) , .A4( u1_u7_u3_n122 ) , .A3( u1_u7_u3_n123 ) , .A1( u1_u7_u3_n175 ) , .A2( u1_u7_u3_n180 ) );
  INV_X1 u1_u7_u3_U93 (.A( u1_u7_u3_n126 ) , .ZN( u1_u7_u3_n180 ) );
  INV_X1 u1_u7_u3_U94 (.A( u1_u7_u3_n112 ) , .ZN( u1_u7_u3_n175 ) );
  NAND4_X1 u1_u7_u3_U95 (.ZN( u1_out7_1 ) , .A4( u1_u7_u3_n161 ) , .A3( u1_u7_u3_n162 ) , .A2( u1_u7_u3_n163 ) , .A1( u1_u7_u3_n185 ) );
  NAND2_X1 u1_u7_u3_U96 (.ZN( u1_u7_u3_n163 ) , .A2( u1_u7_u3_n170 ) , .A1( u1_u7_u3_n176 ) );
  AOI22_X1 u1_u7_u3_U97 (.B2( u1_u7_u3_n140 ) , .B1( u1_u7_u3_n141 ) , .A2( u1_u7_u3_n142 ) , .ZN( u1_u7_u3_n162 ) , .A1( u1_u7_u3_n177 ) );
  NAND3_X1 u1_u7_u3_U98 (.A1( u1_u7_u3_n114 ) , .ZN( u1_u7_u3_n115 ) , .A2( u1_u7_u3_n145 ) , .A3( u1_u7_u3_n153 ) );
  NAND3_X1 u1_u7_u3_U99 (.ZN( u1_u7_u3_n129 ) , .A2( u1_u7_u3_n144 ) , .A1( u1_u7_u3_n153 ) , .A3( u1_u7_u3_n182 ) );
  XOR2_X1 u1_u9_U33 (.B( u1_K10_24 ) , .A( u1_R8_17 ) , .Z( u1_u9_X_24 ) );
  XOR2_X1 u1_u9_U34 (.B( u1_K10_23 ) , .A( u1_R8_16 ) , .Z( u1_u9_X_23 ) );
  XOR2_X1 u1_u9_U35 (.B( u1_K10_22 ) , .A( u1_R8_15 ) , .Z( u1_u9_X_22 ) );
  XOR2_X1 u1_u9_U36 (.B( u1_K10_21 ) , .A( u1_R8_14 ) , .Z( u1_u9_X_21 ) );
  XOR2_X1 u1_u9_U37 (.B( u1_K10_20 ) , .A( u1_R8_13 ) , .Z( u1_u9_X_20 ) );
  XOR2_X1 u1_u9_U39 (.B( u1_K10_19 ) , .A( u1_R8_12 ) , .Z( u1_u9_X_19 ) );
  OAI22_X1 u1_u9_u3_U10 (.B1( u1_u9_u3_n113 ) , .A2( u1_u9_u3_n135 ) , .A1( u1_u9_u3_n150 ) , .B2( u1_u9_u3_n164 ) , .ZN( u1_u9_u3_n98 ) );
  OAI211_X1 u1_u9_u3_U11 (.B( u1_u9_u3_n106 ) , .ZN( u1_u9_u3_n119 ) , .C2( u1_u9_u3_n128 ) , .C1( u1_u9_u3_n167 ) , .A( u1_u9_u3_n181 ) );
  AOI221_X1 u1_u9_u3_U12 (.C1( u1_u9_u3_n105 ) , .ZN( u1_u9_u3_n106 ) , .A( u1_u9_u3_n131 ) , .B2( u1_u9_u3_n132 ) , .C2( u1_u9_u3_n133 ) , .B1( u1_u9_u3_n169 ) );
  INV_X1 u1_u9_u3_U13 (.ZN( u1_u9_u3_n181 ) , .A( u1_u9_u3_n98 ) );
  NAND2_X1 u1_u9_u3_U14 (.ZN( u1_u9_u3_n105 ) , .A2( u1_u9_u3_n130 ) , .A1( u1_u9_u3_n155 ) );
  AOI22_X1 u1_u9_u3_U15 (.B1( u1_u9_u3_n115 ) , .A2( u1_u9_u3_n116 ) , .ZN( u1_u9_u3_n123 ) , .B2( u1_u9_u3_n133 ) , .A1( u1_u9_u3_n169 ) );
  NAND2_X1 u1_u9_u3_U16 (.ZN( u1_u9_u3_n116 ) , .A2( u1_u9_u3_n151 ) , .A1( u1_u9_u3_n182 ) );
  NOR2_X1 u1_u9_u3_U17 (.ZN( u1_u9_u3_n126 ) , .A2( u1_u9_u3_n150 ) , .A1( u1_u9_u3_n164 ) );
  AOI21_X1 u1_u9_u3_U18 (.ZN( u1_u9_u3_n112 ) , .B2( u1_u9_u3_n146 ) , .B1( u1_u9_u3_n155 ) , .A( u1_u9_u3_n167 ) );
  NAND2_X1 u1_u9_u3_U19 (.A1( u1_u9_u3_n135 ) , .ZN( u1_u9_u3_n142 ) , .A2( u1_u9_u3_n164 ) );
  NAND2_X1 u1_u9_u3_U20 (.ZN( u1_u9_u3_n132 ) , .A2( u1_u9_u3_n152 ) , .A1( u1_u9_u3_n156 ) );
  AND2_X1 u1_u9_u3_U21 (.A2( u1_u9_u3_n113 ) , .A1( u1_u9_u3_n114 ) , .ZN( u1_u9_u3_n151 ) );
  INV_X1 u1_u9_u3_U22 (.A( u1_u9_u3_n133 ) , .ZN( u1_u9_u3_n165 ) );
  INV_X1 u1_u9_u3_U23 (.A( u1_u9_u3_n135 ) , .ZN( u1_u9_u3_n170 ) );
  NAND2_X1 u1_u9_u3_U24 (.A1( u1_u9_u3_n107 ) , .A2( u1_u9_u3_n108 ) , .ZN( u1_u9_u3_n140 ) );
  NAND2_X1 u1_u9_u3_U25 (.ZN( u1_u9_u3_n117 ) , .A1( u1_u9_u3_n124 ) , .A2( u1_u9_u3_n148 ) );
  NAND2_X1 u1_u9_u3_U26 (.ZN( u1_u9_u3_n143 ) , .A1( u1_u9_u3_n165 ) , .A2( u1_u9_u3_n167 ) );
  INV_X1 u1_u9_u3_U27 (.A( u1_u9_u3_n130 ) , .ZN( u1_u9_u3_n177 ) );
  INV_X1 u1_u9_u3_U28 (.A( u1_u9_u3_n128 ) , .ZN( u1_u9_u3_n176 ) );
  INV_X1 u1_u9_u3_U29 (.A( u1_u9_u3_n155 ) , .ZN( u1_u9_u3_n174 ) );
  INV_X1 u1_u9_u3_U3 (.A( u1_u9_u3_n129 ) , .ZN( u1_u9_u3_n183 ) );
  INV_X1 u1_u9_u3_U30 (.A( u1_u9_u3_n139 ) , .ZN( u1_u9_u3_n185 ) );
  NOR2_X1 u1_u9_u3_U31 (.ZN( u1_u9_u3_n135 ) , .A2( u1_u9_u3_n141 ) , .A1( u1_u9_u3_n169 ) );
  OAI222_X1 u1_u9_u3_U32 (.C2( u1_u9_u3_n107 ) , .A2( u1_u9_u3_n108 ) , .B1( u1_u9_u3_n135 ) , .ZN( u1_u9_u3_n138 ) , .B2( u1_u9_u3_n146 ) , .C1( u1_u9_u3_n154 ) , .A1( u1_u9_u3_n164 ) );
  NOR4_X1 u1_u9_u3_U33 (.A4( u1_u9_u3_n157 ) , .A3( u1_u9_u3_n158 ) , .A2( u1_u9_u3_n159 ) , .A1( u1_u9_u3_n160 ) , .ZN( u1_u9_u3_n161 ) );
  AOI21_X1 u1_u9_u3_U34 (.B2( u1_u9_u3_n152 ) , .B1( u1_u9_u3_n153 ) , .ZN( u1_u9_u3_n158 ) , .A( u1_u9_u3_n164 ) );
  AOI21_X1 u1_u9_u3_U35 (.A( u1_u9_u3_n154 ) , .B2( u1_u9_u3_n155 ) , .B1( u1_u9_u3_n156 ) , .ZN( u1_u9_u3_n157 ) );
  AOI21_X1 u1_u9_u3_U36 (.A( u1_u9_u3_n149 ) , .B2( u1_u9_u3_n150 ) , .B1( u1_u9_u3_n151 ) , .ZN( u1_u9_u3_n159 ) );
  AOI211_X1 u1_u9_u3_U37 (.ZN( u1_u9_u3_n109 ) , .A( u1_u9_u3_n119 ) , .C2( u1_u9_u3_n129 ) , .B( u1_u9_u3_n138 ) , .C1( u1_u9_u3_n141 ) );
  AOI211_X1 u1_u9_u3_U38 (.B( u1_u9_u3_n119 ) , .A( u1_u9_u3_n120 ) , .C2( u1_u9_u3_n121 ) , .ZN( u1_u9_u3_n122 ) , .C1( u1_u9_u3_n179 ) );
  INV_X1 u1_u9_u3_U39 (.A( u1_u9_u3_n156 ) , .ZN( u1_u9_u3_n179 ) );
  INV_X1 u1_u9_u3_U4 (.A( u1_u9_u3_n140 ) , .ZN( u1_u9_u3_n182 ) );
  OAI22_X1 u1_u9_u3_U40 (.B1( u1_u9_u3_n118 ) , .ZN( u1_u9_u3_n120 ) , .A1( u1_u9_u3_n135 ) , .B2( u1_u9_u3_n154 ) , .A2( u1_u9_u3_n178 ) );
  AND3_X1 u1_u9_u3_U41 (.ZN( u1_u9_u3_n118 ) , .A2( u1_u9_u3_n124 ) , .A1( u1_u9_u3_n144 ) , .A3( u1_u9_u3_n152 ) );
  INV_X1 u1_u9_u3_U42 (.A( u1_u9_u3_n121 ) , .ZN( u1_u9_u3_n164 ) );
  NAND2_X1 u1_u9_u3_U43 (.ZN( u1_u9_u3_n133 ) , .A1( u1_u9_u3_n154 ) , .A2( u1_u9_u3_n164 ) );
  OAI211_X1 u1_u9_u3_U44 (.B( u1_u9_u3_n127 ) , .ZN( u1_u9_u3_n139 ) , .C1( u1_u9_u3_n150 ) , .C2( u1_u9_u3_n154 ) , .A( u1_u9_u3_n184 ) );
  INV_X1 u1_u9_u3_U45 (.A( u1_u9_u3_n125 ) , .ZN( u1_u9_u3_n184 ) );
  AOI221_X1 u1_u9_u3_U46 (.A( u1_u9_u3_n126 ) , .ZN( u1_u9_u3_n127 ) , .C2( u1_u9_u3_n132 ) , .C1( u1_u9_u3_n169 ) , .B2( u1_u9_u3_n170 ) , .B1( u1_u9_u3_n174 ) );
  OAI22_X1 u1_u9_u3_U47 (.A1( u1_u9_u3_n124 ) , .ZN( u1_u9_u3_n125 ) , .B2( u1_u9_u3_n145 ) , .A2( u1_u9_u3_n165 ) , .B1( u1_u9_u3_n167 ) );
  NOR2_X1 u1_u9_u3_U48 (.A1( u1_u9_u3_n113 ) , .ZN( u1_u9_u3_n131 ) , .A2( u1_u9_u3_n154 ) );
  NAND2_X1 u1_u9_u3_U49 (.A1( u1_u9_u3_n103 ) , .ZN( u1_u9_u3_n150 ) , .A2( u1_u9_u3_n99 ) );
  INV_X1 u1_u9_u3_U5 (.A( u1_u9_u3_n117 ) , .ZN( u1_u9_u3_n178 ) );
  NAND2_X1 u1_u9_u3_U50 (.A2( u1_u9_u3_n102 ) , .ZN( u1_u9_u3_n155 ) , .A1( u1_u9_u3_n97 ) );
  INV_X1 u1_u9_u3_U51 (.A( u1_u9_u3_n141 ) , .ZN( u1_u9_u3_n167 ) );
  AOI21_X1 u1_u9_u3_U52 (.B2( u1_u9_u3_n114 ) , .B1( u1_u9_u3_n146 ) , .A( u1_u9_u3_n154 ) , .ZN( u1_u9_u3_n94 ) );
  AOI21_X1 u1_u9_u3_U53 (.ZN( u1_u9_u3_n110 ) , .B2( u1_u9_u3_n142 ) , .B1( u1_u9_u3_n186 ) , .A( u1_u9_u3_n95 ) );
  INV_X1 u1_u9_u3_U54 (.A( u1_u9_u3_n145 ) , .ZN( u1_u9_u3_n186 ) );
  AOI21_X1 u1_u9_u3_U55 (.B1( u1_u9_u3_n124 ) , .A( u1_u9_u3_n149 ) , .B2( u1_u9_u3_n155 ) , .ZN( u1_u9_u3_n95 ) );
  INV_X1 u1_u9_u3_U56 (.A( u1_u9_u3_n149 ) , .ZN( u1_u9_u3_n169 ) );
  NAND2_X1 u1_u9_u3_U57 (.ZN( u1_u9_u3_n124 ) , .A1( u1_u9_u3_n96 ) , .A2( u1_u9_u3_n97 ) );
  NAND2_X1 u1_u9_u3_U58 (.A2( u1_u9_u3_n100 ) , .ZN( u1_u9_u3_n146 ) , .A1( u1_u9_u3_n96 ) );
  NAND2_X1 u1_u9_u3_U59 (.A1( u1_u9_u3_n101 ) , .ZN( u1_u9_u3_n145 ) , .A2( u1_u9_u3_n99 ) );
  AOI221_X1 u1_u9_u3_U6 (.A( u1_u9_u3_n131 ) , .C2( u1_u9_u3_n132 ) , .C1( u1_u9_u3_n133 ) , .ZN( u1_u9_u3_n134 ) , .B1( u1_u9_u3_n143 ) , .B2( u1_u9_u3_n177 ) );
  NAND2_X1 u1_u9_u3_U60 (.A1( u1_u9_u3_n100 ) , .ZN( u1_u9_u3_n156 ) , .A2( u1_u9_u3_n99 ) );
  NAND2_X1 u1_u9_u3_U61 (.A2( u1_u9_u3_n101 ) , .A1( u1_u9_u3_n104 ) , .ZN( u1_u9_u3_n148 ) );
  NAND2_X1 u1_u9_u3_U62 (.A1( u1_u9_u3_n100 ) , .A2( u1_u9_u3_n102 ) , .ZN( u1_u9_u3_n128 ) );
  NAND2_X1 u1_u9_u3_U63 (.A2( u1_u9_u3_n101 ) , .A1( u1_u9_u3_n102 ) , .ZN( u1_u9_u3_n152 ) );
  NAND2_X1 u1_u9_u3_U64 (.A2( u1_u9_u3_n101 ) , .ZN( u1_u9_u3_n114 ) , .A1( u1_u9_u3_n96 ) );
  NAND2_X1 u1_u9_u3_U65 (.ZN( u1_u9_u3_n107 ) , .A1( u1_u9_u3_n97 ) , .A2( u1_u9_u3_n99 ) );
  NAND2_X1 u1_u9_u3_U66 (.A2( u1_u9_u3_n100 ) , .A1( u1_u9_u3_n104 ) , .ZN( u1_u9_u3_n113 ) );
  NAND2_X1 u1_u9_u3_U67 (.A1( u1_u9_u3_n104 ) , .ZN( u1_u9_u3_n153 ) , .A2( u1_u9_u3_n97 ) );
  NAND2_X1 u1_u9_u3_U68 (.A2( u1_u9_u3_n103 ) , .A1( u1_u9_u3_n104 ) , .ZN( u1_u9_u3_n130 ) );
  NAND2_X1 u1_u9_u3_U69 (.A2( u1_u9_u3_n103 ) , .ZN( u1_u9_u3_n144 ) , .A1( u1_u9_u3_n96 ) );
  OAI22_X1 u1_u9_u3_U7 (.B2( u1_u9_u3_n147 ) , .A2( u1_u9_u3_n148 ) , .ZN( u1_u9_u3_n160 ) , .B1( u1_u9_u3_n165 ) , .A1( u1_u9_u3_n168 ) );
  NAND2_X1 u1_u9_u3_U70 (.A1( u1_u9_u3_n102 ) , .A2( u1_u9_u3_n103 ) , .ZN( u1_u9_u3_n108 ) );
  NOR2_X1 u1_u9_u3_U71 (.A2( u1_u9_X_19 ) , .A1( u1_u9_X_20 ) , .ZN( u1_u9_u3_n99 ) );
  NOR2_X1 u1_u9_u3_U72 (.A2( u1_u9_X_21 ) , .A1( u1_u9_X_24 ) , .ZN( u1_u9_u3_n103 ) );
  NOR2_X1 u1_u9_u3_U73 (.A2( u1_u9_X_24 ) , .A1( u1_u9_u3_n171 ) , .ZN( u1_u9_u3_n97 ) );
  NOR2_X1 u1_u9_u3_U74 (.A2( u1_u9_X_23 ) , .ZN( u1_u9_u3_n141 ) , .A1( u1_u9_u3_n166 ) );
  NOR2_X1 u1_u9_u3_U75 (.A2( u1_u9_X_19 ) , .A1( u1_u9_u3_n172 ) , .ZN( u1_u9_u3_n96 ) );
  NAND2_X1 u1_u9_u3_U76 (.A1( u1_u9_X_22 ) , .A2( u1_u9_X_23 ) , .ZN( u1_u9_u3_n154 ) );
  NAND2_X1 u1_u9_u3_U77 (.A1( u1_u9_X_23 ) , .ZN( u1_u9_u3_n149 ) , .A2( u1_u9_u3_n166 ) );
  NOR2_X1 u1_u9_u3_U78 (.A2( u1_u9_X_22 ) , .A1( u1_u9_X_23 ) , .ZN( u1_u9_u3_n121 ) );
  AND2_X1 u1_u9_u3_U79 (.A1( u1_u9_X_24 ) , .ZN( u1_u9_u3_n101 ) , .A2( u1_u9_u3_n171 ) );
  AND3_X1 u1_u9_u3_U8 (.A3( u1_u9_u3_n144 ) , .A2( u1_u9_u3_n145 ) , .A1( u1_u9_u3_n146 ) , .ZN( u1_u9_u3_n147 ) );
  AND2_X1 u1_u9_u3_U80 (.A1( u1_u9_X_19 ) , .ZN( u1_u9_u3_n102 ) , .A2( u1_u9_u3_n172 ) );
  AND2_X1 u1_u9_u3_U81 (.A1( u1_u9_X_21 ) , .A2( u1_u9_X_24 ) , .ZN( u1_u9_u3_n100 ) );
  AND2_X1 u1_u9_u3_U82 (.A2( u1_u9_X_19 ) , .A1( u1_u9_X_20 ) , .ZN( u1_u9_u3_n104 ) );
  INV_X1 u1_u9_u3_U83 (.A( u1_u9_X_22 ) , .ZN( u1_u9_u3_n166 ) );
  INV_X1 u1_u9_u3_U84 (.A( u1_u9_X_21 ) , .ZN( u1_u9_u3_n171 ) );
  INV_X1 u1_u9_u3_U85 (.A( u1_u9_X_20 ) , .ZN( u1_u9_u3_n172 ) );
  OR4_X1 u1_u9_u3_U86 (.ZN( u1_out9_10 ) , .A4( u1_u9_u3_n136 ) , .A3( u1_u9_u3_n137 ) , .A1( u1_u9_u3_n138 ) , .A2( u1_u9_u3_n139 ) );
  OAI222_X1 u1_u9_u3_U87 (.C1( u1_u9_u3_n128 ) , .ZN( u1_u9_u3_n137 ) , .B1( u1_u9_u3_n148 ) , .A2( u1_u9_u3_n150 ) , .B2( u1_u9_u3_n154 ) , .C2( u1_u9_u3_n164 ) , .A1( u1_u9_u3_n167 ) );
  OAI221_X1 u1_u9_u3_U88 (.A( u1_u9_u3_n134 ) , .B2( u1_u9_u3_n135 ) , .ZN( u1_u9_u3_n136 ) , .C1( u1_u9_u3_n149 ) , .B1( u1_u9_u3_n151 ) , .C2( u1_u9_u3_n183 ) );
  NAND4_X1 u1_u9_u3_U89 (.ZN( u1_out9_26 ) , .A4( u1_u9_u3_n109 ) , .A3( u1_u9_u3_n110 ) , .A2( u1_u9_u3_n111 ) , .A1( u1_u9_u3_n173 ) );
  INV_X1 u1_u9_u3_U9 (.A( u1_u9_u3_n143 ) , .ZN( u1_u9_u3_n168 ) );
  INV_X1 u1_u9_u3_U90 (.ZN( u1_u9_u3_n173 ) , .A( u1_u9_u3_n94 ) );
  OAI21_X1 u1_u9_u3_U91 (.ZN( u1_u9_u3_n111 ) , .B2( u1_u9_u3_n117 ) , .A( u1_u9_u3_n133 ) , .B1( u1_u9_u3_n176 ) );
  NAND4_X1 u1_u9_u3_U92 (.ZN( u1_out9_20 ) , .A4( u1_u9_u3_n122 ) , .A3( u1_u9_u3_n123 ) , .A1( u1_u9_u3_n175 ) , .A2( u1_u9_u3_n180 ) );
  INV_X1 u1_u9_u3_U93 (.A( u1_u9_u3_n126 ) , .ZN( u1_u9_u3_n180 ) );
  INV_X1 u1_u9_u3_U94 (.A( u1_u9_u3_n112 ) , .ZN( u1_u9_u3_n175 ) );
  NAND4_X1 u1_u9_u3_U95 (.ZN( u1_out9_1 ) , .A4( u1_u9_u3_n161 ) , .A3( u1_u9_u3_n162 ) , .A2( u1_u9_u3_n163 ) , .A1( u1_u9_u3_n185 ) );
  NAND2_X1 u1_u9_u3_U96 (.ZN( u1_u9_u3_n163 ) , .A2( u1_u9_u3_n170 ) , .A1( u1_u9_u3_n176 ) );
  AOI22_X1 u1_u9_u3_U97 (.B2( u1_u9_u3_n140 ) , .B1( u1_u9_u3_n141 ) , .A2( u1_u9_u3_n142 ) , .ZN( u1_u9_u3_n162 ) , .A1( u1_u9_u3_n177 ) );
  NAND3_X1 u1_u9_u3_U98 (.A1( u1_u9_u3_n114 ) , .ZN( u1_u9_u3_n115 ) , .A2( u1_u9_u3_n145 ) , .A3( u1_u9_u3_n153 ) );
  NAND3_X1 u1_u9_u3_U99 (.ZN( u1_u9_u3_n129 ) , .A2( u1_u9_u3_n144 ) , .A1( u1_u9_u3_n153 ) , .A3( u1_u9_u3_n182 ) );
  OAI21_X1 u1_uk_U1018 (.ZN( u1_K3_45 ) , .A( u1_uk_n1046 ) , .B2( u1_uk_n1335 ) , .B1( u1_uk_n161 ) );
  NAND2_X1 u1_uk_U1019 (.A1( u1_uk_K_r1_16 ) , .ZN( u1_uk_n1046 ) , .A2( u1_uk_n17 ) );
  OAI21_X1 u1_uk_U1024 (.ZN( u1_K10_21 ) , .B2( u1_uk_n1660 ) , .A( u1_uk_n308 ) , .B1( u1_uk_n60 ) );
  NAND2_X1 u1_uk_U1025 (.A1( u1_uk_K_r8_19 ) , .ZN( u1_uk_n308 ) , .A2( u1_uk_n31 ) );
  OAI21_X1 u1_uk_U1052 (.ZN( u1_K4_28 ) , .A( u1_uk_n1059 ) , .B2( u1_uk_n1381 ) , .B1( u1_uk_n148 ) );
  NAND2_X1 u1_uk_U1053 (.A1( u1_uk_K_r2_21 ) , .A2( u1_uk_n10 ) , .ZN( u1_uk_n1059 ) );
  OAI21_X1 u1_uk_U1109 (.ZN( u1_K3_40 ) , .A( u1_uk_n1044 ) , .B2( u1_uk_n1330 ) , .B1( u1_uk_n209 ) );
  NAND2_X1 u1_uk_U1110 (.A1( u1_uk_K_r1_21 ) , .ZN( u1_uk_n1044 ) , .A2( u1_uk_n292 ) );
  OAI22_X1 u1_uk_U122 (.ZN( u1_K3_41 ) , .A2( u1_uk_n1313 ) , .B2( u1_uk_n1318 ) , .A1( u1_uk_n147 ) , .B1( u1_uk_n207 ) );
  INV_X1 u1_uk_U159 (.ZN( u1_K14_19 ) , .A( u1_uk_n951 ) );
  AOI22_X1 u1_uk_U160 (.B2( u1_uk_K_r12_25 ) , .A2( u1_uk_K_r12_33 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n231 ) , .ZN( u1_uk_n951 ) );
  OAI22_X1 u1_uk_U172 (.ZN( u1_K8_19 ) , .B2( u1_uk_n1538 ) , .A2( u1_uk_n1545 ) , .A1( u1_uk_n277 ) , .B1( u1_uk_n92 ) );
  OAI22_X1 u1_uk_U173 (.ZN( u1_K10_19 ) , .A1( u1_uk_n117 ) , .B2( u1_uk_n1633 ) , .A2( u1_uk_n1643 ) , .B1( u1_uk_n238 ) );
  INV_X1 u1_uk_U177 (.ZN( u1_K12_30 ) , .A( u1_uk_n526 ) );
  AOI22_X1 u1_uk_U178 (.B2( u1_uk_K_r10_23 ) , .A2( u1_uk_K_r10_42 ) , .A1( u1_uk_n182 ) , .B1( u1_uk_n271 ) , .ZN( u1_uk_n526 ) );
  OAI21_X1 u1_uk_U192 (.ZN( u1_K10_24 ) , .B2( u1_uk_n1629 ) , .B1( u1_uk_n17 ) , .A( u1_uk_n319 ) );
  NAND2_X1 u1_uk_U193 (.A1( u1_uk_K_r8_40 ) , .A2( u1_uk_n27 ) , .ZN( u1_uk_n319 ) );
  OAI21_X1 u1_uk_U201 (.ZN( u1_K14_24 ) , .B1( u1_uk_n100 ) , .B2( u1_uk_n1812 ) , .A( u1_uk_n952 ) );
  NAND2_X1 u1_uk_U202 (.A1( u1_uk_K_r12_41 ) , .A2( u1_uk_n10 ) , .ZN( u1_uk_n952 ) );
  OAI21_X1 u1_uk_U213 (.ZN( u1_K4_30 ) , .A( u1_uk_n1062 ) , .B2( u1_uk_n1375 ) , .B1( u1_uk_n252 ) );
  NAND2_X1 u1_uk_U214 (.A1( u1_uk_K_r2_28 ) , .ZN( u1_uk_n1062 ) , .A2( u1_uk_n230 ) );
  OAI21_X1 u1_uk_U283 (.ZN( u1_K3_44 ) , .A( u1_uk_n1045 ) , .B2( u1_uk_n1314 ) , .B1( u1_uk_n161 ) );
  NAND2_X1 u1_uk_U284 (.A1( u1_uk_K_r1_15 ) , .ZN( u1_uk_n1045 ) , .A2( u1_uk_n17 ) );
  OAI22_X1 u1_uk_U285 (.ZN( u1_K3_48 ) , .B2( u1_uk_n1307 ) , .A2( u1_uk_n1342 ) , .A1( u1_uk_n148 ) , .B1( u1_uk_n207 ) );
  INV_X1 u1_uk_U317 (.ZN( u1_K4_26 ) , .A( u1_uk_n1058 ) );
  AOI22_X1 u1_uk_U318 (.B2( u1_uk_K_r2_16 ) , .A2( u1_uk_K_r2_7 ) , .ZN( u1_uk_n1058 ) , .B1( u1_uk_n162 ) , .A1( u1_uk_n207 ) );
  OAI22_X1 u1_uk_U331 (.ZN( u1_K12_26 ) , .A1( u1_uk_n118 ) , .A2( u1_uk_n1710 ) , .B2( u1_uk_n1720 ) , .B1( u1_uk_n271 ) );
  OAI21_X1 u1_uk_U340 (.ZN( u1_K3_46 ) , .A( u1_uk_n1047 ) , .B2( u1_uk_n1327 ) , .B1( u1_uk_n292 ) );
  NAND2_X1 u1_uk_U341 (.A1( u1_uk_K_r1_22 ) , .ZN( u1_uk_n1047 ) , .A2( u1_uk_n251 ) );
  OAI22_X1 u1_uk_U391 (.ZN( u1_K12_28 ) , .A1( u1_uk_n142 ) , .B2( u1_uk_n1710 ) , .A2( u1_uk_n1714 ) , .B1( u1_uk_n242 ) );
  OAI22_X1 u1_uk_U479 (.ZN( u1_K3_37 ) , .B2( u1_uk_n1322 ) , .A2( u1_uk_n1328 ) , .A1( u1_uk_n292 ) , .B1( u1_uk_n94 ) );
  INV_X1 u1_uk_U501 (.ZN( u1_K4_29 ) , .A( u1_uk_n1060 ) );
  AOI22_X1 u1_uk_U502 (.B2( u1_uk_K_r2_31 ) , .A2( u1_uk_K_r2_36 ) , .ZN( u1_uk_n1060 ) , .A1( u1_uk_n109 ) , .B1( u1_uk_n214 ) );
  OAI22_X1 u1_uk_U503 (.ZN( u1_K12_29 ) , .B1( u1_uk_n100 ) , .B2( u1_uk_n1721 ) , .A2( u1_uk_n1744 ) , .A1( u1_uk_n286 ) );
  INV_X1 u1_uk_U603 (.ZN( u1_K10_22 ) , .A( u1_uk_n312 ) );
  AOI22_X1 u1_uk_U604 (.B2( u1_uk_K_r8_27 ) , .A2( u1_uk_K_r8_5 ) , .B1( u1_uk_n148 ) , .A1( u1_uk_n279 ) , .ZN( u1_uk_n312 ) );
  OAI22_X1 u1_uk_U607 (.ZN( u1_K8_22 ) , .B2( u1_uk_n1559 ) , .A2( u1_uk_n1565 ) , .A1( u1_uk_n217 ) , .B1( u1_uk_n60 ) );
  INV_X1 u1_uk_U608 (.ZN( u1_K5_22 ) , .A( u1_uk_n1074 ) );
  AOI22_X1 u1_uk_U609 (.B2( u1_uk_K_r3_24 ) , .A2( u1_uk_K_r3_33 ) , .ZN( u1_uk_n1074 ) , .B1( u1_uk_n222 ) , .A1( u1_uk_n31 ) );
  OAI22_X1 u1_uk_U658 (.ZN( u1_K3_43 ) , .B2( u1_uk_n1334 ) , .A2( u1_uk_n1338 ) , .A1( u1_uk_n286 ) , .B1( u1_uk_n94 ) );
  OAI22_X1 u1_uk_U695 (.ZN( u1_K12_25 ) , .A1( u1_uk_n128 ) , .B2( u1_uk_n1729 ) , .A2( u1_uk_n1734 ) , .B1( u1_uk_n298 ) );
  INV_X1 u1_uk_U715 (.ZN( u1_K4_25 ) , .A( u1_uk_n1057 ) );
  AOI22_X1 u1_uk_U716 (.B2( u1_uk_K_r2_16 ) , .A2( u1_uk_K_r2_49 ) , .ZN( u1_uk_n1057 ) , .A1( u1_uk_n17 ) , .B1( u1_uk_n292 ) );
  OAI22_X1 u1_uk_U738 (.ZN( u1_K3_42 ) , .B2( u1_uk_n1307 ) , .A2( u1_uk_n1334 ) , .A1( u1_uk_n292 ) , .B1( u1_uk_n94 ) );
  OAI22_X1 u1_uk_U750 (.ZN( u1_K12_27 ) , .A1( u1_uk_n118 ) , .B2( u1_uk_n1717 ) , .A2( u1_uk_n1749 ) , .B1( u1_uk_n286 ) );
  OAI22_X1 u1_uk_U765 (.ZN( u1_K14_21 ) , .A1( u1_uk_n145 ) , .B2( u1_uk_n1814 ) , .A2( u1_uk_n1840 ) , .B1( u1_uk_n220 ) );
  OAI22_X1 u1_uk_U769 (.ZN( u1_K5_21 ) , .A1( u1_uk_n118 ) , .B2( u1_uk_n1409 ) , .A2( u1_uk_n1429 ) , .B1( u1_uk_n202 ) );
  OAI22_X1 u1_uk_U776 (.ZN( u1_K4_27 ) , .B1( u1_uk_n109 ) , .B2( u1_uk_n1350 ) , .A2( u1_uk_n1376 ) , .A1( u1_uk_n286 ) );
  OAI22_X1 u1_uk_U830 (.ZN( u1_K8_20 ) , .B1( u1_uk_n147 ) , .B2( u1_uk_n1551 ) , .A2( u1_uk_n1557 ) , .A1( u1_uk_n222 ) );
  INV_X1 u1_uk_U839 (.ZN( u1_K5_20 ) , .A( u1_uk_n1073 ) );
  AOI22_X1 u1_uk_U840 (.B2( u1_uk_K_r3_24 ) , .A2( u1_uk_K_r3_47 ) , .ZN( u1_uk_n1073 ) , .A1( u1_uk_n202 ) , .B1( u1_uk_n83 ) );
  OAI22_X1 u1_uk_U867 (.ZN( u1_K14_22 ) , .B1( u1_uk_n109 ) , .B2( u1_uk_n1802 ) , .A2( u1_uk_n1840 ) , .A1( u1_uk_n277 ) );
  OAI22_X1 u1_uk_U873 (.ZN( u1_K14_23 ) , .B1( u1_uk_n102 ) , .A2( u1_uk_n1802 ) , .B2( u1_uk_n1809 ) , .A1( u1_uk_n291 ) );
  OAI22_X1 u1_uk_U874 (.ZN( u1_K5_23 ) , .B1( u1_uk_n11 ) , .B2( u1_uk_n1415 ) , .A2( u1_uk_n1424 ) , .A1( u1_uk_n242 ) );
  OAI22_X1 u1_uk_U877 (.ZN( u1_K3_47 ) , .B2( u1_uk_n1327 ) , .A2( u1_uk_n1335 ) , .A1( u1_uk_n251 ) , .B1( u1_uk_n94 ) );
  OAI21_X1 u1_uk_U90 (.ZN( u1_K10_23 ) , .B2( u1_uk_n1620 ) , .B1( u1_uk_n294 ) , .A( u1_uk_n313 ) );
  OAI22_X1 u1_uk_U904 (.ZN( u1_K5_19 ) , .A2( u1_uk_n1398 ) , .B2( u1_uk_n1435 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n217 ) );
  OAI22_X1 u1_uk_U905 (.ZN( u1_K5_24 ) , .B2( u1_uk_n1402 ) , .A2( u1_uk_n1427 ) , .B1( u1_uk_n145 ) , .A1( u1_uk_n242 ) );
  OAI22_X1 u1_uk_U908 (.ZN( u1_K8_21 ) , .B2( u1_uk_n1552 ) , .A2( u1_uk_n1558 ) , .B1( u1_uk_n17 ) , .A1( u1_uk_n252 ) );
  NAND2_X1 u1_uk_U91 (.A1( u1_uk_K_r8_13 ) , .A2( u1_uk_n271 ) , .ZN( u1_uk_n313 ) );
  OAI22_X1 u1_uk_U92 (.ZN( u1_K8_23 ) , .B2( u1_uk_n1543 ) , .A2( u1_uk_n1548 ) , .A1( u1_uk_n279 ) , .B1( u1_uk_n93 ) );
  OAI22_X1 u1_uk_U925 (.ZN( u1_K3_38 ) , .A2( u1_uk_n1314 ) , .B2( u1_uk_n1330 ) , .A1( u1_uk_n207 ) , .B1( u1_uk_n94 ) );
  OAI22_X1 u1_uk_U926 (.ZN( u1_K3_39 ) , .B2( u1_uk_n1338 ) , .A2( u1_uk_n1342 ) , .A1( u1_uk_n203 ) , .B1( u1_uk_n94 ) );
  OAI22_X1 u1_uk_U939 (.ZN( u1_K14_20 ) , .A1( u1_uk_n146 ) , .B2( u1_uk_n1813 ) , .A2( u1_uk_n1819 ) , .B1( u1_uk_n220 ) );
  OAI22_X1 u1_uk_U943 (.ZN( u1_K8_24 ) , .B2( u1_uk_n1530 ) , .A1( u1_uk_n155 ) , .A2( u1_uk_n1570 ) , .B1( u1_uk_n286 ) );
  OAI22_X1 u1_uk_U963 (.ZN( u1_K10_20 ) , .B2( u1_uk_n1629 ) , .A1( u1_uk_n163 ) , .A2( u1_uk_n1659 ) , .B1( u1_uk_n191 ) );
  XOR2_X1 u2_U136 (.B( u2_L0_10 ) , .Z( u2_N41 ) , .A( u2_out1_10 ) );
  XOR2_X1 u2_U192 (.B( u2_L0_5 ) , .Z( u2_N36 ) , .A( u2_out1_5 ) );
  XOR2_X1 u2_U236 (.B( u2_L0_1 ) , .Z( u2_N32 ) , .A( u2_out1_1 ) );
  XOR2_X1 u2_U313 (.B( u2_L6_27 ) , .Z( u2_N250 ) , .A( u2_out7_27 ) );
  XOR2_X1 u2_U320 (.B( u2_L6_21 ) , .Z( u2_N244 ) , .A( u2_out7_21 ) );
  XOR2_X1 u2_U327 (.B( u2_L6_15 ) , .Z( u2_N238 ) , .A( u2_out7_15 ) );
  XOR2_X1 u2_U338 (.B( u2_L6_5 ) , .Z( u2_N228 ) , .A( u2_out7_5 ) );
  XOR2_X1 u2_U415 (.B( u2_L3_32 ) , .Z( u2_N159 ) , .A( u2_out4_32 ) );
  XOR2_X1 u2_U418 (.B( u2_L3_29 ) , .Z( u2_N156 ) , .A( u2_out4_29 ) );
  XOR2_X1 u2_U426 (.B( u2_L3_22 ) , .Z( u2_N149 ) , .A( u2_out4_22 ) );
  XOR2_X1 u2_U429 (.B( u2_L3_19 ) , .Z( u2_N146 ) , .A( u2_out4_19 ) );
  XOR2_X1 u2_U437 (.B( u2_L3_12 ) , .Z( u2_N139 ) , .A( u2_out4_12 ) );
  XOR2_X1 u2_U438 (.B( u2_L3_11 ) , .Z( u2_N138 ) , .A( u2_out4_11 ) );
  XOR2_X1 u2_U442 (.B( u2_L3_7 ) , .Z( u2_N134 ) , .A( u2_out4_7 ) );
  XOR2_X1 u2_U445 (.B( u2_L3_4 ) , .Z( u2_N131 ) , .A( u2_out4_4 ) );
  XOR2_X1 u2_U48 (.B( u2_L0_27 ) , .Z( u2_N58 ) , .A( u2_out1_27 ) );
  XOR2_X1 u2_U49 (.B( u2_L0_26 ) , .Z( u2_N57 ) , .A( u2_out1_26 ) );
  XOR2_X1 u2_U54 (.B( u2_L0_21 ) , .Z( u2_N52 ) , .A( u2_out1_21 ) );
  XOR2_X1 u2_U55 (.B( u2_L0_20 ) , .Z( u2_N51 ) , .A( u2_out1_20 ) );
  XOR2_X1 u2_U81 (.B( u2_L0_15 ) , .Z( u2_N46 ) , .A( u2_out1_15 ) );
  XOR2_X1 u2_u1_U10 (.B( u2_K2_45 ) , .A( u2_R0_30 ) , .Z( u2_u1_X_45 ) );
  XOR2_X1 u2_u1_U11 (.B( u2_K2_44 ) , .A( u2_R0_29 ) , .Z( u2_u1_X_44 ) );
  XOR2_X1 u2_u1_U12 (.B( u2_K2_43 ) , .A( u2_R0_28 ) , .Z( u2_u1_X_43 ) );
  XOR2_X1 u2_u1_U33 (.B( u2_K2_24 ) , .A( u2_R0_17 ) , .Z( u2_u1_X_24 ) );
  XOR2_X1 u2_u1_U34 (.B( u2_K2_23 ) , .A( u2_R0_16 ) , .Z( u2_u1_X_23 ) );
  XOR2_X1 u2_u1_U35 (.B( u2_K2_22 ) , .A( u2_R0_15 ) , .Z( u2_u1_X_22 ) );
  XOR2_X1 u2_u1_U36 (.B( u2_K2_21 ) , .A( u2_R0_14 ) , .Z( u2_u1_X_21 ) );
  XOR2_X1 u2_u1_U37 (.B( u2_K2_20 ) , .A( u2_R0_13 ) , .Z( u2_u1_X_20 ) );
  XOR2_X1 u2_u1_U39 (.B( u2_K2_19 ) , .A( u2_R0_12 ) , .Z( u2_u1_X_19 ) );
  XOR2_X1 u2_u1_U7 (.B( u2_K2_48 ) , .A( u2_R0_1 ) , .Z( u2_u1_X_48 ) );
  XOR2_X1 u2_u1_U8 (.B( u2_K2_47 ) , .A( u2_R0_32 ) , .Z( u2_u1_X_47 ) );
  XOR2_X1 u2_u1_U9 (.B( u2_K2_46 ) , .A( u2_R0_31 ) , .Z( u2_u1_X_46 ) );
  OAI22_X1 u2_u1_u3_U10 (.B1( u2_u1_u3_n113 ) , .A2( u2_u1_u3_n135 ) , .A1( u2_u1_u3_n150 ) , .B2( u2_u1_u3_n164 ) , .ZN( u2_u1_u3_n98 ) );
  OAI211_X1 u2_u1_u3_U11 (.B( u2_u1_u3_n106 ) , .ZN( u2_u1_u3_n119 ) , .C2( u2_u1_u3_n128 ) , .C1( u2_u1_u3_n167 ) , .A( u2_u1_u3_n181 ) );
  AOI221_X1 u2_u1_u3_U12 (.C1( u2_u1_u3_n105 ) , .ZN( u2_u1_u3_n106 ) , .A( u2_u1_u3_n131 ) , .B2( u2_u1_u3_n132 ) , .C2( u2_u1_u3_n133 ) , .B1( u2_u1_u3_n169 ) );
  INV_X1 u2_u1_u3_U13 (.ZN( u2_u1_u3_n181 ) , .A( u2_u1_u3_n98 ) );
  NAND2_X1 u2_u1_u3_U14 (.ZN( u2_u1_u3_n105 ) , .A2( u2_u1_u3_n130 ) , .A1( u2_u1_u3_n155 ) );
  AOI22_X1 u2_u1_u3_U15 (.B1( u2_u1_u3_n115 ) , .A2( u2_u1_u3_n116 ) , .ZN( u2_u1_u3_n123 ) , .B2( u2_u1_u3_n133 ) , .A1( u2_u1_u3_n169 ) );
  NAND2_X1 u2_u1_u3_U16 (.ZN( u2_u1_u3_n116 ) , .A2( u2_u1_u3_n151 ) , .A1( u2_u1_u3_n182 ) );
  NOR2_X1 u2_u1_u3_U17 (.ZN( u2_u1_u3_n126 ) , .A2( u2_u1_u3_n150 ) , .A1( u2_u1_u3_n164 ) );
  AOI21_X1 u2_u1_u3_U18 (.ZN( u2_u1_u3_n112 ) , .B2( u2_u1_u3_n146 ) , .B1( u2_u1_u3_n155 ) , .A( u2_u1_u3_n167 ) );
  NAND2_X1 u2_u1_u3_U19 (.A1( u2_u1_u3_n135 ) , .ZN( u2_u1_u3_n142 ) , .A2( u2_u1_u3_n164 ) );
  NAND2_X1 u2_u1_u3_U20 (.ZN( u2_u1_u3_n132 ) , .A2( u2_u1_u3_n152 ) , .A1( u2_u1_u3_n156 ) );
  AND2_X1 u2_u1_u3_U21 (.A2( u2_u1_u3_n113 ) , .A1( u2_u1_u3_n114 ) , .ZN( u2_u1_u3_n151 ) );
  INV_X1 u2_u1_u3_U22 (.A( u2_u1_u3_n133 ) , .ZN( u2_u1_u3_n165 ) );
  INV_X1 u2_u1_u3_U23 (.A( u2_u1_u3_n135 ) , .ZN( u2_u1_u3_n170 ) );
  NAND2_X1 u2_u1_u3_U24 (.A1( u2_u1_u3_n107 ) , .A2( u2_u1_u3_n108 ) , .ZN( u2_u1_u3_n140 ) );
  NAND2_X1 u2_u1_u3_U25 (.ZN( u2_u1_u3_n117 ) , .A1( u2_u1_u3_n124 ) , .A2( u2_u1_u3_n148 ) );
  NAND2_X1 u2_u1_u3_U26 (.ZN( u2_u1_u3_n143 ) , .A1( u2_u1_u3_n165 ) , .A2( u2_u1_u3_n167 ) );
  INV_X1 u2_u1_u3_U27 (.A( u2_u1_u3_n130 ) , .ZN( u2_u1_u3_n177 ) );
  INV_X1 u2_u1_u3_U28 (.A( u2_u1_u3_n128 ) , .ZN( u2_u1_u3_n176 ) );
  INV_X1 u2_u1_u3_U29 (.A( u2_u1_u3_n155 ) , .ZN( u2_u1_u3_n174 ) );
  INV_X1 u2_u1_u3_U3 (.A( u2_u1_u3_n129 ) , .ZN( u2_u1_u3_n183 ) );
  INV_X1 u2_u1_u3_U30 (.A( u2_u1_u3_n139 ) , .ZN( u2_u1_u3_n185 ) );
  NOR2_X1 u2_u1_u3_U31 (.ZN( u2_u1_u3_n135 ) , .A2( u2_u1_u3_n141 ) , .A1( u2_u1_u3_n169 ) );
  OAI222_X1 u2_u1_u3_U32 (.C2( u2_u1_u3_n107 ) , .A2( u2_u1_u3_n108 ) , .B1( u2_u1_u3_n135 ) , .ZN( u2_u1_u3_n138 ) , .B2( u2_u1_u3_n146 ) , .C1( u2_u1_u3_n154 ) , .A1( u2_u1_u3_n164 ) );
  NOR4_X1 u2_u1_u3_U33 (.A4( u2_u1_u3_n157 ) , .A3( u2_u1_u3_n158 ) , .A2( u2_u1_u3_n159 ) , .A1( u2_u1_u3_n160 ) , .ZN( u2_u1_u3_n161 ) );
  AOI21_X1 u2_u1_u3_U34 (.B2( u2_u1_u3_n152 ) , .B1( u2_u1_u3_n153 ) , .ZN( u2_u1_u3_n158 ) , .A( u2_u1_u3_n164 ) );
  AOI21_X1 u2_u1_u3_U35 (.A( u2_u1_u3_n154 ) , .B2( u2_u1_u3_n155 ) , .B1( u2_u1_u3_n156 ) , .ZN( u2_u1_u3_n157 ) );
  AOI21_X1 u2_u1_u3_U36 (.A( u2_u1_u3_n149 ) , .B2( u2_u1_u3_n150 ) , .B1( u2_u1_u3_n151 ) , .ZN( u2_u1_u3_n159 ) );
  AOI211_X1 u2_u1_u3_U37 (.ZN( u2_u1_u3_n109 ) , .A( u2_u1_u3_n119 ) , .C2( u2_u1_u3_n129 ) , .B( u2_u1_u3_n138 ) , .C1( u2_u1_u3_n141 ) );
  AOI211_X1 u2_u1_u3_U38 (.B( u2_u1_u3_n119 ) , .A( u2_u1_u3_n120 ) , .C2( u2_u1_u3_n121 ) , .ZN( u2_u1_u3_n122 ) , .C1( u2_u1_u3_n179 ) );
  INV_X1 u2_u1_u3_U39 (.A( u2_u1_u3_n156 ) , .ZN( u2_u1_u3_n179 ) );
  INV_X1 u2_u1_u3_U4 (.A( u2_u1_u3_n140 ) , .ZN( u2_u1_u3_n182 ) );
  OAI22_X1 u2_u1_u3_U40 (.B1( u2_u1_u3_n118 ) , .ZN( u2_u1_u3_n120 ) , .A1( u2_u1_u3_n135 ) , .B2( u2_u1_u3_n154 ) , .A2( u2_u1_u3_n178 ) );
  AND3_X1 u2_u1_u3_U41 (.ZN( u2_u1_u3_n118 ) , .A2( u2_u1_u3_n124 ) , .A1( u2_u1_u3_n144 ) , .A3( u2_u1_u3_n152 ) );
  INV_X1 u2_u1_u3_U42 (.A( u2_u1_u3_n121 ) , .ZN( u2_u1_u3_n164 ) );
  NAND2_X1 u2_u1_u3_U43 (.ZN( u2_u1_u3_n133 ) , .A1( u2_u1_u3_n154 ) , .A2( u2_u1_u3_n164 ) );
  OAI211_X1 u2_u1_u3_U44 (.B( u2_u1_u3_n127 ) , .ZN( u2_u1_u3_n139 ) , .C1( u2_u1_u3_n150 ) , .C2( u2_u1_u3_n154 ) , .A( u2_u1_u3_n184 ) );
  INV_X1 u2_u1_u3_U45 (.A( u2_u1_u3_n125 ) , .ZN( u2_u1_u3_n184 ) );
  AOI221_X1 u2_u1_u3_U46 (.A( u2_u1_u3_n126 ) , .ZN( u2_u1_u3_n127 ) , .C2( u2_u1_u3_n132 ) , .C1( u2_u1_u3_n169 ) , .B2( u2_u1_u3_n170 ) , .B1( u2_u1_u3_n174 ) );
  OAI22_X1 u2_u1_u3_U47 (.A1( u2_u1_u3_n124 ) , .ZN( u2_u1_u3_n125 ) , .B2( u2_u1_u3_n145 ) , .A2( u2_u1_u3_n165 ) , .B1( u2_u1_u3_n167 ) );
  NOR2_X1 u2_u1_u3_U48 (.A1( u2_u1_u3_n113 ) , .ZN( u2_u1_u3_n131 ) , .A2( u2_u1_u3_n154 ) );
  NAND2_X1 u2_u1_u3_U49 (.A1( u2_u1_u3_n103 ) , .ZN( u2_u1_u3_n150 ) , .A2( u2_u1_u3_n99 ) );
  INV_X1 u2_u1_u3_U5 (.A( u2_u1_u3_n117 ) , .ZN( u2_u1_u3_n178 ) );
  NAND2_X1 u2_u1_u3_U50 (.A2( u2_u1_u3_n102 ) , .ZN( u2_u1_u3_n155 ) , .A1( u2_u1_u3_n97 ) );
  INV_X1 u2_u1_u3_U51 (.A( u2_u1_u3_n141 ) , .ZN( u2_u1_u3_n167 ) );
  AOI21_X1 u2_u1_u3_U52 (.B2( u2_u1_u3_n114 ) , .B1( u2_u1_u3_n146 ) , .A( u2_u1_u3_n154 ) , .ZN( u2_u1_u3_n94 ) );
  AOI21_X1 u2_u1_u3_U53 (.ZN( u2_u1_u3_n110 ) , .B2( u2_u1_u3_n142 ) , .B1( u2_u1_u3_n186 ) , .A( u2_u1_u3_n95 ) );
  INV_X1 u2_u1_u3_U54 (.A( u2_u1_u3_n145 ) , .ZN( u2_u1_u3_n186 ) );
  AOI21_X1 u2_u1_u3_U55 (.B1( u2_u1_u3_n124 ) , .A( u2_u1_u3_n149 ) , .B2( u2_u1_u3_n155 ) , .ZN( u2_u1_u3_n95 ) );
  INV_X1 u2_u1_u3_U56 (.A( u2_u1_u3_n149 ) , .ZN( u2_u1_u3_n169 ) );
  NAND2_X1 u2_u1_u3_U57 (.ZN( u2_u1_u3_n124 ) , .A1( u2_u1_u3_n96 ) , .A2( u2_u1_u3_n97 ) );
  NAND2_X1 u2_u1_u3_U58 (.A2( u2_u1_u3_n100 ) , .ZN( u2_u1_u3_n146 ) , .A1( u2_u1_u3_n96 ) );
  NAND2_X1 u2_u1_u3_U59 (.A1( u2_u1_u3_n101 ) , .ZN( u2_u1_u3_n145 ) , .A2( u2_u1_u3_n99 ) );
  AOI221_X1 u2_u1_u3_U6 (.A( u2_u1_u3_n131 ) , .C2( u2_u1_u3_n132 ) , .C1( u2_u1_u3_n133 ) , .ZN( u2_u1_u3_n134 ) , .B1( u2_u1_u3_n143 ) , .B2( u2_u1_u3_n177 ) );
  NAND2_X1 u2_u1_u3_U60 (.A1( u2_u1_u3_n100 ) , .ZN( u2_u1_u3_n156 ) , .A2( u2_u1_u3_n99 ) );
  NAND2_X1 u2_u1_u3_U61 (.A2( u2_u1_u3_n101 ) , .A1( u2_u1_u3_n104 ) , .ZN( u2_u1_u3_n148 ) );
  NAND2_X1 u2_u1_u3_U62 (.A1( u2_u1_u3_n100 ) , .A2( u2_u1_u3_n102 ) , .ZN( u2_u1_u3_n128 ) );
  NAND2_X1 u2_u1_u3_U63 (.A2( u2_u1_u3_n101 ) , .A1( u2_u1_u3_n102 ) , .ZN( u2_u1_u3_n152 ) );
  NAND2_X1 u2_u1_u3_U64 (.A2( u2_u1_u3_n101 ) , .ZN( u2_u1_u3_n114 ) , .A1( u2_u1_u3_n96 ) );
  NAND2_X1 u2_u1_u3_U65 (.ZN( u2_u1_u3_n107 ) , .A1( u2_u1_u3_n97 ) , .A2( u2_u1_u3_n99 ) );
  NAND2_X1 u2_u1_u3_U66 (.A2( u2_u1_u3_n100 ) , .A1( u2_u1_u3_n104 ) , .ZN( u2_u1_u3_n113 ) );
  NAND2_X1 u2_u1_u3_U67 (.A1( u2_u1_u3_n104 ) , .ZN( u2_u1_u3_n153 ) , .A2( u2_u1_u3_n97 ) );
  NAND2_X1 u2_u1_u3_U68 (.A2( u2_u1_u3_n103 ) , .A1( u2_u1_u3_n104 ) , .ZN( u2_u1_u3_n130 ) );
  NAND2_X1 u2_u1_u3_U69 (.A2( u2_u1_u3_n103 ) , .ZN( u2_u1_u3_n144 ) , .A1( u2_u1_u3_n96 ) );
  OAI22_X1 u2_u1_u3_U7 (.B2( u2_u1_u3_n147 ) , .A2( u2_u1_u3_n148 ) , .ZN( u2_u1_u3_n160 ) , .B1( u2_u1_u3_n165 ) , .A1( u2_u1_u3_n168 ) );
  NAND2_X1 u2_u1_u3_U70 (.A1( u2_u1_u3_n102 ) , .A2( u2_u1_u3_n103 ) , .ZN( u2_u1_u3_n108 ) );
  NOR2_X1 u2_u1_u3_U71 (.A2( u2_u1_X_19 ) , .A1( u2_u1_X_20 ) , .ZN( u2_u1_u3_n99 ) );
  NOR2_X1 u2_u1_u3_U72 (.A2( u2_u1_X_21 ) , .A1( u2_u1_X_24 ) , .ZN( u2_u1_u3_n103 ) );
  NOR2_X1 u2_u1_u3_U73 (.A2( u2_u1_X_24 ) , .A1( u2_u1_u3_n171 ) , .ZN( u2_u1_u3_n97 ) );
  NOR2_X1 u2_u1_u3_U74 (.A2( u2_u1_X_23 ) , .ZN( u2_u1_u3_n141 ) , .A1( u2_u1_u3_n166 ) );
  NOR2_X1 u2_u1_u3_U75 (.A2( u2_u1_X_19 ) , .A1( u2_u1_u3_n172 ) , .ZN( u2_u1_u3_n96 ) );
  NAND2_X1 u2_u1_u3_U76 (.A1( u2_u1_X_22 ) , .A2( u2_u1_X_23 ) , .ZN( u2_u1_u3_n154 ) );
  NAND2_X1 u2_u1_u3_U77 (.A1( u2_u1_X_23 ) , .ZN( u2_u1_u3_n149 ) , .A2( u2_u1_u3_n166 ) );
  NOR2_X1 u2_u1_u3_U78 (.A2( u2_u1_X_22 ) , .A1( u2_u1_X_23 ) , .ZN( u2_u1_u3_n121 ) );
  AND2_X1 u2_u1_u3_U79 (.A1( u2_u1_X_24 ) , .ZN( u2_u1_u3_n101 ) , .A2( u2_u1_u3_n171 ) );
  AND3_X1 u2_u1_u3_U8 (.A3( u2_u1_u3_n144 ) , .A2( u2_u1_u3_n145 ) , .A1( u2_u1_u3_n146 ) , .ZN( u2_u1_u3_n147 ) );
  AND2_X1 u2_u1_u3_U80 (.A1( u2_u1_X_19 ) , .ZN( u2_u1_u3_n102 ) , .A2( u2_u1_u3_n172 ) );
  AND2_X1 u2_u1_u3_U81 (.A1( u2_u1_X_21 ) , .A2( u2_u1_X_24 ) , .ZN( u2_u1_u3_n100 ) );
  AND2_X1 u2_u1_u3_U82 (.A2( u2_u1_X_19 ) , .A1( u2_u1_X_20 ) , .ZN( u2_u1_u3_n104 ) );
  INV_X1 u2_u1_u3_U83 (.A( u2_u1_X_22 ) , .ZN( u2_u1_u3_n166 ) );
  INV_X1 u2_u1_u3_U84 (.A( u2_u1_X_21 ) , .ZN( u2_u1_u3_n171 ) );
  INV_X1 u2_u1_u3_U85 (.A( u2_u1_X_20 ) , .ZN( u2_u1_u3_n172 ) );
  OR4_X1 u2_u1_u3_U86 (.ZN( u2_out1_10 ) , .A4( u2_u1_u3_n136 ) , .A3( u2_u1_u3_n137 ) , .A1( u2_u1_u3_n138 ) , .A2( u2_u1_u3_n139 ) );
  OAI222_X1 u2_u1_u3_U87 (.C1( u2_u1_u3_n128 ) , .ZN( u2_u1_u3_n137 ) , .B1( u2_u1_u3_n148 ) , .A2( u2_u1_u3_n150 ) , .B2( u2_u1_u3_n154 ) , .C2( u2_u1_u3_n164 ) , .A1( u2_u1_u3_n167 ) );
  OAI221_X1 u2_u1_u3_U88 (.A( u2_u1_u3_n134 ) , .B2( u2_u1_u3_n135 ) , .ZN( u2_u1_u3_n136 ) , .C1( u2_u1_u3_n149 ) , .B1( u2_u1_u3_n151 ) , .C2( u2_u1_u3_n183 ) );
  NAND4_X1 u2_u1_u3_U89 (.ZN( u2_out1_26 ) , .A4( u2_u1_u3_n109 ) , .A3( u2_u1_u3_n110 ) , .A2( u2_u1_u3_n111 ) , .A1( u2_u1_u3_n173 ) );
  INV_X1 u2_u1_u3_U9 (.A( u2_u1_u3_n143 ) , .ZN( u2_u1_u3_n168 ) );
  INV_X1 u2_u1_u3_U90 (.ZN( u2_u1_u3_n173 ) , .A( u2_u1_u3_n94 ) );
  OAI21_X1 u2_u1_u3_U91 (.ZN( u2_u1_u3_n111 ) , .B2( u2_u1_u3_n117 ) , .A( u2_u1_u3_n133 ) , .B1( u2_u1_u3_n176 ) );
  NAND4_X1 u2_u1_u3_U92 (.ZN( u2_out1_20 ) , .A4( u2_u1_u3_n122 ) , .A3( u2_u1_u3_n123 ) , .A1( u2_u1_u3_n175 ) , .A2( u2_u1_u3_n180 ) );
  INV_X1 u2_u1_u3_U93 (.A( u2_u1_u3_n112 ) , .ZN( u2_u1_u3_n175 ) );
  INV_X1 u2_u1_u3_U94 (.A( u2_u1_u3_n126 ) , .ZN( u2_u1_u3_n180 ) );
  NAND4_X1 u2_u1_u3_U95 (.ZN( u2_out1_1 ) , .A4( u2_u1_u3_n161 ) , .A3( u2_u1_u3_n162 ) , .A2( u2_u1_u3_n163 ) , .A1( u2_u1_u3_n185 ) );
  NAND2_X1 u2_u1_u3_U96 (.ZN( u2_u1_u3_n163 ) , .A2( u2_u1_u3_n170 ) , .A1( u2_u1_u3_n176 ) );
  AOI22_X1 u2_u1_u3_U97 (.B2( u2_u1_u3_n140 ) , .B1( u2_u1_u3_n141 ) , .A2( u2_u1_u3_n142 ) , .ZN( u2_u1_u3_n162 ) , .A1( u2_u1_u3_n177 ) );
  NAND3_X1 u2_u1_u3_U98 (.A1( u2_u1_u3_n114 ) , .ZN( u2_u1_u3_n115 ) , .A2( u2_u1_u3_n145 ) , .A3( u2_u1_u3_n153 ) );
  NAND3_X1 u2_u1_u3_U99 (.ZN( u2_u1_u3_n129 ) , .A2( u2_u1_u3_n144 ) , .A1( u2_u1_u3_n153 ) , .A3( u2_u1_u3_n182 ) );
  AND3_X1 u2_u1_u7_U10 (.A3( u2_u1_u7_n110 ) , .A2( u2_u1_u7_n127 ) , .A1( u2_u1_u7_n132 ) , .ZN( u2_u1_u7_n92 ) );
  OAI21_X1 u2_u1_u7_U11 (.A( u2_u1_u7_n161 ) , .B1( u2_u1_u7_n168 ) , .B2( u2_u1_u7_n173 ) , .ZN( u2_u1_u7_n91 ) );
  AOI211_X1 u2_u1_u7_U12 (.A( u2_u1_u7_n117 ) , .ZN( u2_u1_u7_n118 ) , .C2( u2_u1_u7_n126 ) , .C1( u2_u1_u7_n177 ) , .B( u2_u1_u7_n180 ) );
  OAI22_X1 u2_u1_u7_U13 (.B1( u2_u1_u7_n115 ) , .ZN( u2_u1_u7_n117 ) , .A2( u2_u1_u7_n133 ) , .A1( u2_u1_u7_n137 ) , .B2( u2_u1_u7_n162 ) );
  INV_X1 u2_u1_u7_U14 (.A( u2_u1_u7_n116 ) , .ZN( u2_u1_u7_n180 ) );
  NOR3_X1 u2_u1_u7_U15 (.ZN( u2_u1_u7_n115 ) , .A3( u2_u1_u7_n145 ) , .A2( u2_u1_u7_n168 ) , .A1( u2_u1_u7_n169 ) );
  OAI211_X1 u2_u1_u7_U16 (.B( u2_u1_u7_n122 ) , .A( u2_u1_u7_n123 ) , .C2( u2_u1_u7_n124 ) , .ZN( u2_u1_u7_n154 ) , .C1( u2_u1_u7_n162 ) );
  AOI222_X1 u2_u1_u7_U17 (.ZN( u2_u1_u7_n122 ) , .C2( u2_u1_u7_n126 ) , .C1( u2_u1_u7_n145 ) , .B1( u2_u1_u7_n161 ) , .A2( u2_u1_u7_n165 ) , .B2( u2_u1_u7_n170 ) , .A1( u2_u1_u7_n176 ) );
  INV_X1 u2_u1_u7_U18 (.A( u2_u1_u7_n133 ) , .ZN( u2_u1_u7_n176 ) );
  NOR3_X1 u2_u1_u7_U19 (.A2( u2_u1_u7_n134 ) , .A1( u2_u1_u7_n135 ) , .ZN( u2_u1_u7_n136 ) , .A3( u2_u1_u7_n171 ) );
  NOR2_X1 u2_u1_u7_U20 (.A1( u2_u1_u7_n130 ) , .A2( u2_u1_u7_n134 ) , .ZN( u2_u1_u7_n153 ) );
  INV_X1 u2_u1_u7_U21 (.A( u2_u1_u7_n101 ) , .ZN( u2_u1_u7_n165 ) );
  NOR2_X1 u2_u1_u7_U22 (.ZN( u2_u1_u7_n111 ) , .A2( u2_u1_u7_n134 ) , .A1( u2_u1_u7_n169 ) );
  AOI21_X1 u2_u1_u7_U23 (.ZN( u2_u1_u7_n104 ) , .B2( u2_u1_u7_n112 ) , .B1( u2_u1_u7_n127 ) , .A( u2_u1_u7_n164 ) );
  AOI21_X1 u2_u1_u7_U24 (.ZN( u2_u1_u7_n106 ) , .B1( u2_u1_u7_n133 ) , .B2( u2_u1_u7_n146 ) , .A( u2_u1_u7_n162 ) );
  AOI21_X1 u2_u1_u7_U25 (.A( u2_u1_u7_n101 ) , .ZN( u2_u1_u7_n107 ) , .B2( u2_u1_u7_n128 ) , .B1( u2_u1_u7_n175 ) );
  INV_X1 u2_u1_u7_U26 (.A( u2_u1_u7_n138 ) , .ZN( u2_u1_u7_n171 ) );
  INV_X1 u2_u1_u7_U27 (.A( u2_u1_u7_n131 ) , .ZN( u2_u1_u7_n177 ) );
  INV_X1 u2_u1_u7_U28 (.A( u2_u1_u7_n110 ) , .ZN( u2_u1_u7_n174 ) );
  NAND2_X1 u2_u1_u7_U29 (.A1( u2_u1_u7_n129 ) , .A2( u2_u1_u7_n132 ) , .ZN( u2_u1_u7_n149 ) );
  OAI21_X1 u2_u1_u7_U3 (.ZN( u2_u1_u7_n159 ) , .A( u2_u1_u7_n165 ) , .B2( u2_u1_u7_n171 ) , .B1( u2_u1_u7_n174 ) );
  NAND2_X1 u2_u1_u7_U30 (.A1( u2_u1_u7_n113 ) , .A2( u2_u1_u7_n124 ) , .ZN( u2_u1_u7_n130 ) );
  INV_X1 u2_u1_u7_U31 (.A( u2_u1_u7_n112 ) , .ZN( u2_u1_u7_n173 ) );
  INV_X1 u2_u1_u7_U32 (.A( u2_u1_u7_n128 ) , .ZN( u2_u1_u7_n168 ) );
  INV_X1 u2_u1_u7_U33 (.A( u2_u1_u7_n148 ) , .ZN( u2_u1_u7_n169 ) );
  INV_X1 u2_u1_u7_U34 (.A( u2_u1_u7_n127 ) , .ZN( u2_u1_u7_n179 ) );
  NOR2_X1 u2_u1_u7_U35 (.ZN( u2_u1_u7_n101 ) , .A2( u2_u1_u7_n150 ) , .A1( u2_u1_u7_n156 ) );
  AOI211_X1 u2_u1_u7_U36 (.B( u2_u1_u7_n154 ) , .A( u2_u1_u7_n155 ) , .C1( u2_u1_u7_n156 ) , .ZN( u2_u1_u7_n157 ) , .C2( u2_u1_u7_n172 ) );
  INV_X1 u2_u1_u7_U37 (.A( u2_u1_u7_n153 ) , .ZN( u2_u1_u7_n172 ) );
  AOI211_X1 u2_u1_u7_U38 (.B( u2_u1_u7_n139 ) , .A( u2_u1_u7_n140 ) , .C2( u2_u1_u7_n141 ) , .ZN( u2_u1_u7_n142 ) , .C1( u2_u1_u7_n156 ) );
  NAND4_X1 u2_u1_u7_U39 (.A3( u2_u1_u7_n127 ) , .A2( u2_u1_u7_n128 ) , .A1( u2_u1_u7_n129 ) , .ZN( u2_u1_u7_n141 ) , .A4( u2_u1_u7_n147 ) );
  INV_X1 u2_u1_u7_U4 (.A( u2_u1_u7_n111 ) , .ZN( u2_u1_u7_n170 ) );
  AOI21_X1 u2_u1_u7_U40 (.A( u2_u1_u7_n137 ) , .B1( u2_u1_u7_n138 ) , .ZN( u2_u1_u7_n139 ) , .B2( u2_u1_u7_n146 ) );
  OAI22_X1 u2_u1_u7_U41 (.B1( u2_u1_u7_n136 ) , .ZN( u2_u1_u7_n140 ) , .A1( u2_u1_u7_n153 ) , .B2( u2_u1_u7_n162 ) , .A2( u2_u1_u7_n164 ) );
  AOI21_X1 u2_u1_u7_U42 (.ZN( u2_u1_u7_n123 ) , .B1( u2_u1_u7_n165 ) , .B2( u2_u1_u7_n177 ) , .A( u2_u1_u7_n97 ) );
  AOI21_X1 u2_u1_u7_U43 (.B2( u2_u1_u7_n113 ) , .B1( u2_u1_u7_n124 ) , .A( u2_u1_u7_n125 ) , .ZN( u2_u1_u7_n97 ) );
  INV_X1 u2_u1_u7_U44 (.A( u2_u1_u7_n125 ) , .ZN( u2_u1_u7_n161 ) );
  INV_X1 u2_u1_u7_U45 (.A( u2_u1_u7_n152 ) , .ZN( u2_u1_u7_n162 ) );
  AOI22_X1 u2_u1_u7_U46 (.A2( u2_u1_u7_n114 ) , .ZN( u2_u1_u7_n119 ) , .B1( u2_u1_u7_n130 ) , .A1( u2_u1_u7_n156 ) , .B2( u2_u1_u7_n165 ) );
  NAND2_X1 u2_u1_u7_U47 (.A2( u2_u1_u7_n112 ) , .ZN( u2_u1_u7_n114 ) , .A1( u2_u1_u7_n175 ) );
  AND2_X1 u2_u1_u7_U48 (.ZN( u2_u1_u7_n145 ) , .A2( u2_u1_u7_n98 ) , .A1( u2_u1_u7_n99 ) );
  NOR2_X1 u2_u1_u7_U49 (.ZN( u2_u1_u7_n137 ) , .A1( u2_u1_u7_n150 ) , .A2( u2_u1_u7_n161 ) );
  INV_X1 u2_u1_u7_U5 (.A( u2_u1_u7_n149 ) , .ZN( u2_u1_u7_n175 ) );
  AOI21_X1 u2_u1_u7_U50 (.ZN( u2_u1_u7_n105 ) , .B2( u2_u1_u7_n110 ) , .A( u2_u1_u7_n125 ) , .B1( u2_u1_u7_n147 ) );
  NAND2_X1 u2_u1_u7_U51 (.ZN( u2_u1_u7_n146 ) , .A1( u2_u1_u7_n95 ) , .A2( u2_u1_u7_n98 ) );
  NAND2_X1 u2_u1_u7_U52 (.A2( u2_u1_u7_n103 ) , .ZN( u2_u1_u7_n147 ) , .A1( u2_u1_u7_n93 ) );
  NAND2_X1 u2_u1_u7_U53 (.A1( u2_u1_u7_n103 ) , .ZN( u2_u1_u7_n127 ) , .A2( u2_u1_u7_n99 ) );
  OR2_X1 u2_u1_u7_U54 (.ZN( u2_u1_u7_n126 ) , .A2( u2_u1_u7_n152 ) , .A1( u2_u1_u7_n156 ) );
  NAND2_X1 u2_u1_u7_U55 (.A2( u2_u1_u7_n102 ) , .A1( u2_u1_u7_n103 ) , .ZN( u2_u1_u7_n133 ) );
  NAND2_X1 u2_u1_u7_U56 (.ZN( u2_u1_u7_n112 ) , .A2( u2_u1_u7_n96 ) , .A1( u2_u1_u7_n99 ) );
  NAND2_X1 u2_u1_u7_U57 (.A2( u2_u1_u7_n102 ) , .ZN( u2_u1_u7_n128 ) , .A1( u2_u1_u7_n98 ) );
  NAND2_X1 u2_u1_u7_U58 (.A1( u2_u1_u7_n100 ) , .ZN( u2_u1_u7_n113 ) , .A2( u2_u1_u7_n93 ) );
  NAND2_X1 u2_u1_u7_U59 (.A2( u2_u1_u7_n102 ) , .ZN( u2_u1_u7_n124 ) , .A1( u2_u1_u7_n96 ) );
  INV_X1 u2_u1_u7_U6 (.A( u2_u1_u7_n154 ) , .ZN( u2_u1_u7_n178 ) );
  NAND2_X1 u2_u1_u7_U60 (.ZN( u2_u1_u7_n110 ) , .A1( u2_u1_u7_n95 ) , .A2( u2_u1_u7_n96 ) );
  INV_X1 u2_u1_u7_U61 (.A( u2_u1_u7_n150 ) , .ZN( u2_u1_u7_n164 ) );
  AND2_X1 u2_u1_u7_U62 (.ZN( u2_u1_u7_n134 ) , .A1( u2_u1_u7_n93 ) , .A2( u2_u1_u7_n98 ) );
  NAND2_X1 u2_u1_u7_U63 (.A1( u2_u1_u7_n100 ) , .A2( u2_u1_u7_n102 ) , .ZN( u2_u1_u7_n129 ) );
  NAND2_X1 u2_u1_u7_U64 (.A2( u2_u1_u7_n103 ) , .ZN( u2_u1_u7_n131 ) , .A1( u2_u1_u7_n95 ) );
  NAND2_X1 u2_u1_u7_U65 (.A1( u2_u1_u7_n100 ) , .ZN( u2_u1_u7_n138 ) , .A2( u2_u1_u7_n99 ) );
  NAND2_X1 u2_u1_u7_U66 (.ZN( u2_u1_u7_n132 ) , .A1( u2_u1_u7_n93 ) , .A2( u2_u1_u7_n96 ) );
  NAND2_X1 u2_u1_u7_U67 (.A1( u2_u1_u7_n100 ) , .ZN( u2_u1_u7_n148 ) , .A2( u2_u1_u7_n95 ) );
  NOR2_X1 u2_u1_u7_U68 (.A2( u2_u1_X_47 ) , .ZN( u2_u1_u7_n150 ) , .A1( u2_u1_u7_n163 ) );
  NOR2_X1 u2_u1_u7_U69 (.A2( u2_u1_X_43 ) , .A1( u2_u1_X_44 ) , .ZN( u2_u1_u7_n103 ) );
  AOI211_X1 u2_u1_u7_U7 (.ZN( u2_u1_u7_n116 ) , .A( u2_u1_u7_n155 ) , .C1( u2_u1_u7_n161 ) , .C2( u2_u1_u7_n171 ) , .B( u2_u1_u7_n94 ) );
  NOR2_X1 u2_u1_u7_U70 (.A2( u2_u1_X_48 ) , .A1( u2_u1_u7_n166 ) , .ZN( u2_u1_u7_n95 ) );
  NOR2_X1 u2_u1_u7_U71 (.A2( u2_u1_X_45 ) , .A1( u2_u1_X_48 ) , .ZN( u2_u1_u7_n99 ) );
  NOR2_X1 u2_u1_u7_U72 (.A2( u2_u1_X_44 ) , .A1( u2_u1_u7_n167 ) , .ZN( u2_u1_u7_n98 ) );
  NOR2_X1 u2_u1_u7_U73 (.A2( u2_u1_X_46 ) , .A1( u2_u1_X_47 ) , .ZN( u2_u1_u7_n152 ) );
  AND2_X1 u2_u1_u7_U74 (.A1( u2_u1_X_47 ) , .ZN( u2_u1_u7_n156 ) , .A2( u2_u1_u7_n163 ) );
  NAND2_X1 u2_u1_u7_U75 (.A2( u2_u1_X_46 ) , .A1( u2_u1_X_47 ) , .ZN( u2_u1_u7_n125 ) );
  AND2_X1 u2_u1_u7_U76 (.A2( u2_u1_X_45 ) , .A1( u2_u1_X_48 ) , .ZN( u2_u1_u7_n102 ) );
  AND2_X1 u2_u1_u7_U77 (.A2( u2_u1_X_43 ) , .A1( u2_u1_X_44 ) , .ZN( u2_u1_u7_n96 ) );
  AND2_X1 u2_u1_u7_U78 (.A1( u2_u1_X_44 ) , .ZN( u2_u1_u7_n100 ) , .A2( u2_u1_u7_n167 ) );
  AND2_X1 u2_u1_u7_U79 (.A1( u2_u1_X_48 ) , .A2( u2_u1_u7_n166 ) , .ZN( u2_u1_u7_n93 ) );
  OAI222_X1 u2_u1_u7_U8 (.C2( u2_u1_u7_n101 ) , .B2( u2_u1_u7_n111 ) , .A1( u2_u1_u7_n113 ) , .C1( u2_u1_u7_n146 ) , .A2( u2_u1_u7_n162 ) , .B1( u2_u1_u7_n164 ) , .ZN( u2_u1_u7_n94 ) );
  INV_X1 u2_u1_u7_U80 (.A( u2_u1_X_46 ) , .ZN( u2_u1_u7_n163 ) );
  INV_X1 u2_u1_u7_U81 (.A( u2_u1_X_43 ) , .ZN( u2_u1_u7_n167 ) );
  INV_X1 u2_u1_u7_U82 (.A( u2_u1_X_45 ) , .ZN( u2_u1_u7_n166 ) );
  NAND4_X1 u2_u1_u7_U83 (.ZN( u2_out1_27 ) , .A4( u2_u1_u7_n118 ) , .A3( u2_u1_u7_n119 ) , .A2( u2_u1_u7_n120 ) , .A1( u2_u1_u7_n121 ) );
  OAI21_X1 u2_u1_u7_U84 (.ZN( u2_u1_u7_n121 ) , .B2( u2_u1_u7_n145 ) , .A( u2_u1_u7_n150 ) , .B1( u2_u1_u7_n174 ) );
  OAI21_X1 u2_u1_u7_U85 (.ZN( u2_u1_u7_n120 ) , .A( u2_u1_u7_n161 ) , .B2( u2_u1_u7_n170 ) , .B1( u2_u1_u7_n179 ) );
  NAND4_X1 u2_u1_u7_U86 (.ZN( u2_out1_15 ) , .A4( u2_u1_u7_n142 ) , .A3( u2_u1_u7_n143 ) , .A2( u2_u1_u7_n144 ) , .A1( u2_u1_u7_n178 ) );
  OR2_X1 u2_u1_u7_U87 (.A2( u2_u1_u7_n125 ) , .A1( u2_u1_u7_n129 ) , .ZN( u2_u1_u7_n144 ) );
  AOI22_X1 u2_u1_u7_U88 (.A2( u2_u1_u7_n126 ) , .ZN( u2_u1_u7_n143 ) , .B2( u2_u1_u7_n165 ) , .B1( u2_u1_u7_n173 ) , .A1( u2_u1_u7_n174 ) );
  NAND4_X1 u2_u1_u7_U89 (.ZN( u2_out1_5 ) , .A4( u2_u1_u7_n108 ) , .A3( u2_u1_u7_n109 ) , .A1( u2_u1_u7_n116 ) , .A2( u2_u1_u7_n123 ) );
  OAI221_X1 u2_u1_u7_U9 (.C1( u2_u1_u7_n101 ) , .C2( u2_u1_u7_n147 ) , .ZN( u2_u1_u7_n155 ) , .B2( u2_u1_u7_n162 ) , .A( u2_u1_u7_n91 ) , .B1( u2_u1_u7_n92 ) );
  AOI22_X1 u2_u1_u7_U90 (.ZN( u2_u1_u7_n109 ) , .A2( u2_u1_u7_n126 ) , .B2( u2_u1_u7_n145 ) , .B1( u2_u1_u7_n156 ) , .A1( u2_u1_u7_n171 ) );
  NOR4_X1 u2_u1_u7_U91 (.A4( u2_u1_u7_n104 ) , .A3( u2_u1_u7_n105 ) , .A2( u2_u1_u7_n106 ) , .A1( u2_u1_u7_n107 ) , .ZN( u2_u1_u7_n108 ) );
  NAND4_X1 u2_u1_u7_U92 (.ZN( u2_out1_21 ) , .A4( u2_u1_u7_n157 ) , .A3( u2_u1_u7_n158 ) , .A2( u2_u1_u7_n159 ) , .A1( u2_u1_u7_n160 ) );
  OAI21_X1 u2_u1_u7_U93 (.B1( u2_u1_u7_n145 ) , .ZN( u2_u1_u7_n160 ) , .A( u2_u1_u7_n161 ) , .B2( u2_u1_u7_n177 ) );
  AOI22_X1 u2_u1_u7_U94 (.B2( u2_u1_u7_n149 ) , .B1( u2_u1_u7_n150 ) , .A2( u2_u1_u7_n151 ) , .A1( u2_u1_u7_n152 ) , .ZN( u2_u1_u7_n158 ) );
  NAND3_X1 u2_u1_u7_U95 (.A3( u2_u1_u7_n146 ) , .A2( u2_u1_u7_n147 ) , .A1( u2_u1_u7_n148 ) , .ZN( u2_u1_u7_n151 ) );
  NAND3_X1 u2_u1_u7_U96 (.A3( u2_u1_u7_n131 ) , .A2( u2_u1_u7_n132 ) , .A1( u2_u1_u7_n133 ) , .ZN( u2_u1_u7_n135 ) );
  XOR2_X1 u2_u4_U13 (.B( u2_K5_42 ) , .A( u2_R3_29 ) , .Z( u2_u4_X_42 ) );
  XOR2_X1 u2_u4_U14 (.B( u2_K5_41 ) , .A( u2_R3_28 ) , .Z( u2_u4_X_41 ) );
  XOR2_X1 u2_u4_U15 (.B( u2_K5_40 ) , .A( u2_R3_27 ) , .Z( u2_u4_X_40 ) );
  XOR2_X1 u2_u4_U17 (.B( u2_K5_39 ) , .A( u2_R3_26 ) , .Z( u2_u4_X_39 ) );
  XOR2_X1 u2_u4_U18 (.B( u2_K5_38 ) , .A( u2_R3_25 ) , .Z( u2_u4_X_38 ) );
  XOR2_X1 u2_u4_U19 (.B( u2_K5_37 ) , .A( u2_R3_24 ) , .Z( u2_u4_X_37 ) );
  XOR2_X1 u2_u4_U20 (.B( u2_K5_36 ) , .A( u2_R3_25 ) , .Z( u2_u4_X_36 ) );
  XOR2_X1 u2_u4_U21 (.B( u2_K5_35 ) , .A( u2_R3_24 ) , .Z( u2_u4_X_35 ) );
  XOR2_X1 u2_u4_U22 (.B( u2_K5_34 ) , .A( u2_R3_23 ) , .Z( u2_u4_X_34 ) );
  XOR2_X1 u2_u4_U23 (.B( u2_K5_33 ) , .A( u2_R3_22 ) , .Z( u2_u4_X_33 ) );
  XOR2_X1 u2_u4_U24 (.B( u2_K5_32 ) , .A( u2_R3_21 ) , .Z( u2_u4_X_32 ) );
  XOR2_X1 u2_u4_U25 (.B( u2_K5_31 ) , .A( u2_R3_20 ) , .Z( u2_u4_X_31 ) );
  NOR2_X1 u2_u4_u5_U10 (.ZN( u2_u4_u5_n135 ) , .A1( u2_u4_u5_n173 ) , .A2( u2_u4_u5_n176 ) );
  NOR3_X1 u2_u4_u5_U100 (.A3( u2_u4_u5_n141 ) , .A1( u2_u4_u5_n142 ) , .ZN( u2_u4_u5_n143 ) , .A2( u2_u4_u5_n191 ) );
  NAND4_X1 u2_u4_u5_U101 (.ZN( u2_out4_4 ) , .A4( u2_u4_u5_n112 ) , .A2( u2_u4_u5_n113 ) , .A1( u2_u4_u5_n114 ) , .A3( u2_u4_u5_n195 ) );
  AOI211_X1 u2_u4_u5_U102 (.A( u2_u4_u5_n110 ) , .C1( u2_u4_u5_n111 ) , .ZN( u2_u4_u5_n112 ) , .B( u2_u4_u5_n118 ) , .C2( u2_u4_u5_n177 ) );
  INV_X1 u2_u4_u5_U103 (.A( u2_u4_u5_n102 ) , .ZN( u2_u4_u5_n195 ) );
  NAND3_X1 u2_u4_u5_U104 (.A2( u2_u4_u5_n154 ) , .A3( u2_u4_u5_n158 ) , .A1( u2_u4_u5_n161 ) , .ZN( u2_u4_u5_n99 ) );
  INV_X1 u2_u4_u5_U11 (.A( u2_u4_u5_n121 ) , .ZN( u2_u4_u5_n177 ) );
  NOR2_X1 u2_u4_u5_U12 (.ZN( u2_u4_u5_n160 ) , .A2( u2_u4_u5_n173 ) , .A1( u2_u4_u5_n177 ) );
  INV_X1 u2_u4_u5_U13 (.A( u2_u4_u5_n150 ) , .ZN( u2_u4_u5_n174 ) );
  AOI21_X1 u2_u4_u5_U14 (.A( u2_u4_u5_n160 ) , .B2( u2_u4_u5_n161 ) , .ZN( u2_u4_u5_n162 ) , .B1( u2_u4_u5_n192 ) );
  INV_X1 u2_u4_u5_U15 (.A( u2_u4_u5_n159 ) , .ZN( u2_u4_u5_n192 ) );
  AOI21_X1 u2_u4_u5_U16 (.A( u2_u4_u5_n156 ) , .B2( u2_u4_u5_n157 ) , .B1( u2_u4_u5_n158 ) , .ZN( u2_u4_u5_n163 ) );
  AOI21_X1 u2_u4_u5_U17 (.B2( u2_u4_u5_n139 ) , .B1( u2_u4_u5_n140 ) , .ZN( u2_u4_u5_n141 ) , .A( u2_u4_u5_n150 ) );
  OAI21_X1 u2_u4_u5_U18 (.A( u2_u4_u5_n133 ) , .B2( u2_u4_u5_n134 ) , .B1( u2_u4_u5_n135 ) , .ZN( u2_u4_u5_n142 ) );
  OAI21_X1 u2_u4_u5_U19 (.ZN( u2_u4_u5_n133 ) , .B2( u2_u4_u5_n147 ) , .A( u2_u4_u5_n173 ) , .B1( u2_u4_u5_n188 ) );
  NAND2_X1 u2_u4_u5_U20 (.A2( u2_u4_u5_n119 ) , .A1( u2_u4_u5_n123 ) , .ZN( u2_u4_u5_n137 ) );
  INV_X1 u2_u4_u5_U21 (.A( u2_u4_u5_n155 ) , .ZN( u2_u4_u5_n194 ) );
  NAND2_X1 u2_u4_u5_U22 (.A1( u2_u4_u5_n121 ) , .ZN( u2_u4_u5_n132 ) , .A2( u2_u4_u5_n172 ) );
  NAND2_X1 u2_u4_u5_U23 (.A2( u2_u4_u5_n122 ) , .ZN( u2_u4_u5_n136 ) , .A1( u2_u4_u5_n154 ) );
  NAND2_X1 u2_u4_u5_U24 (.A2( u2_u4_u5_n119 ) , .A1( u2_u4_u5_n120 ) , .ZN( u2_u4_u5_n159 ) );
  INV_X1 u2_u4_u5_U25 (.A( u2_u4_u5_n156 ) , .ZN( u2_u4_u5_n175 ) );
  INV_X1 u2_u4_u5_U26 (.A( u2_u4_u5_n158 ) , .ZN( u2_u4_u5_n188 ) );
  INV_X1 u2_u4_u5_U27 (.A( u2_u4_u5_n152 ) , .ZN( u2_u4_u5_n179 ) );
  INV_X1 u2_u4_u5_U28 (.A( u2_u4_u5_n140 ) , .ZN( u2_u4_u5_n182 ) );
  INV_X1 u2_u4_u5_U29 (.A( u2_u4_u5_n151 ) , .ZN( u2_u4_u5_n183 ) );
  NOR2_X1 u2_u4_u5_U3 (.ZN( u2_u4_u5_n134 ) , .A1( u2_u4_u5_n183 ) , .A2( u2_u4_u5_n190 ) );
  INV_X1 u2_u4_u5_U30 (.A( u2_u4_u5_n123 ) , .ZN( u2_u4_u5_n185 ) );
  INV_X1 u2_u4_u5_U31 (.A( u2_u4_u5_n161 ) , .ZN( u2_u4_u5_n184 ) );
  INV_X1 u2_u4_u5_U32 (.A( u2_u4_u5_n139 ) , .ZN( u2_u4_u5_n189 ) );
  INV_X1 u2_u4_u5_U33 (.A( u2_u4_u5_n157 ) , .ZN( u2_u4_u5_n190 ) );
  INV_X1 u2_u4_u5_U34 (.A( u2_u4_u5_n120 ) , .ZN( u2_u4_u5_n193 ) );
  NAND2_X1 u2_u4_u5_U35 (.ZN( u2_u4_u5_n111 ) , .A1( u2_u4_u5_n140 ) , .A2( u2_u4_u5_n155 ) );
  INV_X1 u2_u4_u5_U36 (.A( u2_u4_u5_n117 ) , .ZN( u2_u4_u5_n196 ) );
  OAI221_X1 u2_u4_u5_U37 (.A( u2_u4_u5_n116 ) , .ZN( u2_u4_u5_n117 ) , .B2( u2_u4_u5_n119 ) , .C1( u2_u4_u5_n153 ) , .C2( u2_u4_u5_n158 ) , .B1( u2_u4_u5_n172 ) );
  AOI222_X1 u2_u4_u5_U38 (.ZN( u2_u4_u5_n116 ) , .B2( u2_u4_u5_n145 ) , .C1( u2_u4_u5_n148 ) , .A2( u2_u4_u5_n174 ) , .C2( u2_u4_u5_n177 ) , .B1( u2_u4_u5_n187 ) , .A1( u2_u4_u5_n193 ) );
  INV_X1 u2_u4_u5_U39 (.A( u2_u4_u5_n115 ) , .ZN( u2_u4_u5_n187 ) );
  INV_X1 u2_u4_u5_U4 (.A( u2_u4_u5_n138 ) , .ZN( u2_u4_u5_n191 ) );
  NOR2_X1 u2_u4_u5_U40 (.ZN( u2_u4_u5_n100 ) , .A1( u2_u4_u5_n170 ) , .A2( u2_u4_u5_n180 ) );
  OAI221_X1 u2_u4_u5_U41 (.A( u2_u4_u5_n101 ) , .ZN( u2_u4_u5_n102 ) , .C2( u2_u4_u5_n115 ) , .C1( u2_u4_u5_n126 ) , .B1( u2_u4_u5_n134 ) , .B2( u2_u4_u5_n160 ) );
  OAI21_X1 u2_u4_u5_U42 (.ZN( u2_u4_u5_n101 ) , .B1( u2_u4_u5_n137 ) , .A( u2_u4_u5_n146 ) , .B2( u2_u4_u5_n147 ) );
  AOI22_X1 u2_u4_u5_U43 (.B2( u2_u4_u5_n131 ) , .A2( u2_u4_u5_n146 ) , .ZN( u2_u4_u5_n169 ) , .B1( u2_u4_u5_n174 ) , .A1( u2_u4_u5_n185 ) );
  NOR2_X1 u2_u4_u5_U44 (.A1( u2_u4_u5_n146 ) , .ZN( u2_u4_u5_n150 ) , .A2( u2_u4_u5_n173 ) );
  AOI21_X1 u2_u4_u5_U45 (.A( u2_u4_u5_n118 ) , .B2( u2_u4_u5_n145 ) , .ZN( u2_u4_u5_n168 ) , .B1( u2_u4_u5_n186 ) );
  INV_X1 u2_u4_u5_U46 (.A( u2_u4_u5_n122 ) , .ZN( u2_u4_u5_n186 ) );
  NOR2_X1 u2_u4_u5_U47 (.A1( u2_u4_u5_n146 ) , .ZN( u2_u4_u5_n152 ) , .A2( u2_u4_u5_n176 ) );
  NOR2_X1 u2_u4_u5_U48 (.A1( u2_u4_u5_n115 ) , .ZN( u2_u4_u5_n118 ) , .A2( u2_u4_u5_n153 ) );
  NOR2_X1 u2_u4_u5_U49 (.A2( u2_u4_u5_n145 ) , .ZN( u2_u4_u5_n156 ) , .A1( u2_u4_u5_n174 ) );
  OAI21_X1 u2_u4_u5_U5 (.B2( u2_u4_u5_n136 ) , .B1( u2_u4_u5_n137 ) , .ZN( u2_u4_u5_n138 ) , .A( u2_u4_u5_n177 ) );
  NOR2_X1 u2_u4_u5_U50 (.ZN( u2_u4_u5_n121 ) , .A2( u2_u4_u5_n145 ) , .A1( u2_u4_u5_n176 ) );
  AOI22_X1 u2_u4_u5_U51 (.ZN( u2_u4_u5_n114 ) , .A2( u2_u4_u5_n137 ) , .A1( u2_u4_u5_n145 ) , .B2( u2_u4_u5_n175 ) , .B1( u2_u4_u5_n193 ) );
  OAI211_X1 u2_u4_u5_U52 (.B( u2_u4_u5_n124 ) , .A( u2_u4_u5_n125 ) , .C2( u2_u4_u5_n126 ) , .C1( u2_u4_u5_n127 ) , .ZN( u2_u4_u5_n128 ) );
  NOR3_X1 u2_u4_u5_U53 (.ZN( u2_u4_u5_n127 ) , .A1( u2_u4_u5_n136 ) , .A3( u2_u4_u5_n148 ) , .A2( u2_u4_u5_n182 ) );
  OAI21_X1 u2_u4_u5_U54 (.ZN( u2_u4_u5_n124 ) , .A( u2_u4_u5_n177 ) , .B2( u2_u4_u5_n183 ) , .B1( u2_u4_u5_n189 ) );
  OAI21_X1 u2_u4_u5_U55 (.ZN( u2_u4_u5_n125 ) , .A( u2_u4_u5_n174 ) , .B2( u2_u4_u5_n185 ) , .B1( u2_u4_u5_n190 ) );
  AOI21_X1 u2_u4_u5_U56 (.A( u2_u4_u5_n153 ) , .B2( u2_u4_u5_n154 ) , .B1( u2_u4_u5_n155 ) , .ZN( u2_u4_u5_n164 ) );
  AOI21_X1 u2_u4_u5_U57 (.ZN( u2_u4_u5_n110 ) , .B1( u2_u4_u5_n122 ) , .B2( u2_u4_u5_n139 ) , .A( u2_u4_u5_n153 ) );
  INV_X1 u2_u4_u5_U58 (.A( u2_u4_u5_n153 ) , .ZN( u2_u4_u5_n176 ) );
  INV_X1 u2_u4_u5_U59 (.A( u2_u4_u5_n126 ) , .ZN( u2_u4_u5_n173 ) );
  AOI222_X1 u2_u4_u5_U6 (.ZN( u2_u4_u5_n113 ) , .A1( u2_u4_u5_n131 ) , .C1( u2_u4_u5_n148 ) , .B2( u2_u4_u5_n174 ) , .C2( u2_u4_u5_n178 ) , .A2( u2_u4_u5_n179 ) , .B1( u2_u4_u5_n99 ) );
  AND2_X1 u2_u4_u5_U60 (.A2( u2_u4_u5_n104 ) , .A1( u2_u4_u5_n107 ) , .ZN( u2_u4_u5_n147 ) );
  AND2_X1 u2_u4_u5_U61 (.A2( u2_u4_u5_n104 ) , .A1( u2_u4_u5_n108 ) , .ZN( u2_u4_u5_n148 ) );
  NAND2_X1 u2_u4_u5_U62 (.A1( u2_u4_u5_n105 ) , .A2( u2_u4_u5_n106 ) , .ZN( u2_u4_u5_n158 ) );
  NAND2_X1 u2_u4_u5_U63 (.A2( u2_u4_u5_n108 ) , .A1( u2_u4_u5_n109 ) , .ZN( u2_u4_u5_n139 ) );
  NAND2_X1 u2_u4_u5_U64 (.A1( u2_u4_u5_n106 ) , .A2( u2_u4_u5_n108 ) , .ZN( u2_u4_u5_n119 ) );
  NAND2_X1 u2_u4_u5_U65 (.A2( u2_u4_u5_n103 ) , .A1( u2_u4_u5_n105 ) , .ZN( u2_u4_u5_n140 ) );
  NAND2_X1 u2_u4_u5_U66 (.A2( u2_u4_u5_n104 ) , .A1( u2_u4_u5_n105 ) , .ZN( u2_u4_u5_n155 ) );
  NAND2_X1 u2_u4_u5_U67 (.A2( u2_u4_u5_n106 ) , .A1( u2_u4_u5_n107 ) , .ZN( u2_u4_u5_n122 ) );
  NAND2_X1 u2_u4_u5_U68 (.A2( u2_u4_u5_n100 ) , .A1( u2_u4_u5_n106 ) , .ZN( u2_u4_u5_n115 ) );
  NAND2_X1 u2_u4_u5_U69 (.A2( u2_u4_u5_n100 ) , .A1( u2_u4_u5_n103 ) , .ZN( u2_u4_u5_n161 ) );
  INV_X1 u2_u4_u5_U7 (.A( u2_u4_u5_n135 ) , .ZN( u2_u4_u5_n178 ) );
  NAND2_X1 u2_u4_u5_U70 (.A1( u2_u4_u5_n105 ) , .A2( u2_u4_u5_n109 ) , .ZN( u2_u4_u5_n154 ) );
  INV_X1 u2_u4_u5_U71 (.A( u2_u4_u5_n146 ) , .ZN( u2_u4_u5_n172 ) );
  NAND2_X1 u2_u4_u5_U72 (.A1( u2_u4_u5_n103 ) , .A2( u2_u4_u5_n108 ) , .ZN( u2_u4_u5_n123 ) );
  NAND2_X1 u2_u4_u5_U73 (.A2( u2_u4_u5_n103 ) , .A1( u2_u4_u5_n107 ) , .ZN( u2_u4_u5_n151 ) );
  NAND2_X1 u2_u4_u5_U74 (.A2( u2_u4_u5_n107 ) , .A1( u2_u4_u5_n109 ) , .ZN( u2_u4_u5_n120 ) );
  NAND2_X1 u2_u4_u5_U75 (.A2( u2_u4_u5_n100 ) , .A1( u2_u4_u5_n109 ) , .ZN( u2_u4_u5_n157 ) );
  AND2_X1 u2_u4_u5_U76 (.A2( u2_u4_u5_n100 ) , .A1( u2_u4_u5_n104 ) , .ZN( u2_u4_u5_n131 ) );
  NOR2_X1 u2_u4_u5_U77 (.A2( u2_u4_X_34 ) , .A1( u2_u4_X_35 ) , .ZN( u2_u4_u5_n145 ) );
  NOR2_X1 u2_u4_u5_U78 (.A2( u2_u4_X_34 ) , .ZN( u2_u4_u5_n146 ) , .A1( u2_u4_u5_n171 ) );
  NOR2_X1 u2_u4_u5_U79 (.A2( u2_u4_X_31 ) , .A1( u2_u4_X_32 ) , .ZN( u2_u4_u5_n103 ) );
  OAI22_X1 u2_u4_u5_U8 (.B2( u2_u4_u5_n149 ) , .B1( u2_u4_u5_n150 ) , .A2( u2_u4_u5_n151 ) , .A1( u2_u4_u5_n152 ) , .ZN( u2_u4_u5_n165 ) );
  NOR2_X1 u2_u4_u5_U80 (.A2( u2_u4_X_36 ) , .ZN( u2_u4_u5_n105 ) , .A1( u2_u4_u5_n180 ) );
  NOR2_X1 u2_u4_u5_U81 (.A2( u2_u4_X_33 ) , .ZN( u2_u4_u5_n108 ) , .A1( u2_u4_u5_n170 ) );
  NOR2_X1 u2_u4_u5_U82 (.A2( u2_u4_X_33 ) , .A1( u2_u4_X_36 ) , .ZN( u2_u4_u5_n107 ) );
  NOR2_X1 u2_u4_u5_U83 (.A2( u2_u4_X_31 ) , .ZN( u2_u4_u5_n104 ) , .A1( u2_u4_u5_n181 ) );
  NAND2_X1 u2_u4_u5_U84 (.A2( u2_u4_X_34 ) , .A1( u2_u4_X_35 ) , .ZN( u2_u4_u5_n153 ) );
  NAND2_X1 u2_u4_u5_U85 (.A1( u2_u4_X_34 ) , .ZN( u2_u4_u5_n126 ) , .A2( u2_u4_u5_n171 ) );
  AND2_X1 u2_u4_u5_U86 (.A1( u2_u4_X_31 ) , .A2( u2_u4_X_32 ) , .ZN( u2_u4_u5_n106 ) );
  AND2_X1 u2_u4_u5_U87 (.A1( u2_u4_X_31 ) , .ZN( u2_u4_u5_n109 ) , .A2( u2_u4_u5_n181 ) );
  INV_X1 u2_u4_u5_U88 (.A( u2_u4_X_33 ) , .ZN( u2_u4_u5_n180 ) );
  INV_X1 u2_u4_u5_U89 (.A( u2_u4_X_35 ) , .ZN( u2_u4_u5_n171 ) );
  NOR3_X1 u2_u4_u5_U9 (.A2( u2_u4_u5_n147 ) , .A1( u2_u4_u5_n148 ) , .ZN( u2_u4_u5_n149 ) , .A3( u2_u4_u5_n194 ) );
  INV_X1 u2_u4_u5_U90 (.A( u2_u4_X_36 ) , .ZN( u2_u4_u5_n170 ) );
  INV_X1 u2_u4_u5_U91 (.A( u2_u4_X_32 ) , .ZN( u2_u4_u5_n181 ) );
  NAND4_X1 u2_u4_u5_U92 (.ZN( u2_out4_29 ) , .A4( u2_u4_u5_n129 ) , .A3( u2_u4_u5_n130 ) , .A2( u2_u4_u5_n168 ) , .A1( u2_u4_u5_n196 ) );
  AOI221_X1 u2_u4_u5_U93 (.A( u2_u4_u5_n128 ) , .ZN( u2_u4_u5_n129 ) , .C2( u2_u4_u5_n132 ) , .B2( u2_u4_u5_n159 ) , .B1( u2_u4_u5_n176 ) , .C1( u2_u4_u5_n184 ) );
  AOI222_X1 u2_u4_u5_U94 (.ZN( u2_u4_u5_n130 ) , .A2( u2_u4_u5_n146 ) , .B1( u2_u4_u5_n147 ) , .C2( u2_u4_u5_n175 ) , .B2( u2_u4_u5_n179 ) , .A1( u2_u4_u5_n188 ) , .C1( u2_u4_u5_n194 ) );
  NAND4_X1 u2_u4_u5_U95 (.ZN( u2_out4_19 ) , .A4( u2_u4_u5_n166 ) , .A3( u2_u4_u5_n167 ) , .A2( u2_u4_u5_n168 ) , .A1( u2_u4_u5_n169 ) );
  AOI22_X1 u2_u4_u5_U96 (.B2( u2_u4_u5_n145 ) , .A2( u2_u4_u5_n146 ) , .ZN( u2_u4_u5_n167 ) , .B1( u2_u4_u5_n182 ) , .A1( u2_u4_u5_n189 ) );
  NOR4_X1 u2_u4_u5_U97 (.A4( u2_u4_u5_n162 ) , .A3( u2_u4_u5_n163 ) , .A2( u2_u4_u5_n164 ) , .A1( u2_u4_u5_n165 ) , .ZN( u2_u4_u5_n166 ) );
  NAND4_X1 u2_u4_u5_U98 (.ZN( u2_out4_11 ) , .A4( u2_u4_u5_n143 ) , .A3( u2_u4_u5_n144 ) , .A2( u2_u4_u5_n169 ) , .A1( u2_u4_u5_n196 ) );
  AOI22_X1 u2_u4_u5_U99 (.A2( u2_u4_u5_n132 ) , .ZN( u2_u4_u5_n144 ) , .B2( u2_u4_u5_n145 ) , .B1( u2_u4_u5_n184 ) , .A1( u2_u4_u5_n194 ) );
  AOI22_X1 u2_u4_u6_U10 (.A2( u2_u4_u6_n151 ) , .B2( u2_u4_u6_n161 ) , .A1( u2_u4_u6_n167 ) , .B1( u2_u4_u6_n170 ) , .ZN( u2_u4_u6_n89 ) );
  AOI21_X1 u2_u4_u6_U11 (.B1( u2_u4_u6_n107 ) , .B2( u2_u4_u6_n132 ) , .A( u2_u4_u6_n158 ) , .ZN( u2_u4_u6_n88 ) );
  AOI21_X1 u2_u4_u6_U12 (.B2( u2_u4_u6_n147 ) , .B1( u2_u4_u6_n148 ) , .ZN( u2_u4_u6_n149 ) , .A( u2_u4_u6_n158 ) );
  AOI21_X1 u2_u4_u6_U13 (.ZN( u2_u4_u6_n106 ) , .A( u2_u4_u6_n142 ) , .B2( u2_u4_u6_n159 ) , .B1( u2_u4_u6_n164 ) );
  INV_X1 u2_u4_u6_U14 (.A( u2_u4_u6_n155 ) , .ZN( u2_u4_u6_n161 ) );
  INV_X1 u2_u4_u6_U15 (.A( u2_u4_u6_n128 ) , .ZN( u2_u4_u6_n164 ) );
  NAND2_X1 u2_u4_u6_U16 (.ZN( u2_u4_u6_n110 ) , .A1( u2_u4_u6_n122 ) , .A2( u2_u4_u6_n129 ) );
  NAND2_X1 u2_u4_u6_U17 (.ZN( u2_u4_u6_n124 ) , .A2( u2_u4_u6_n146 ) , .A1( u2_u4_u6_n148 ) );
  INV_X1 u2_u4_u6_U18 (.A( u2_u4_u6_n132 ) , .ZN( u2_u4_u6_n171 ) );
  AND2_X1 u2_u4_u6_U19 (.A1( u2_u4_u6_n100 ) , .ZN( u2_u4_u6_n130 ) , .A2( u2_u4_u6_n147 ) );
  INV_X1 u2_u4_u6_U20 (.A( u2_u4_u6_n127 ) , .ZN( u2_u4_u6_n173 ) );
  INV_X1 u2_u4_u6_U21 (.A( u2_u4_u6_n121 ) , .ZN( u2_u4_u6_n167 ) );
  INV_X1 u2_u4_u6_U22 (.A( u2_u4_u6_n100 ) , .ZN( u2_u4_u6_n169 ) );
  INV_X1 u2_u4_u6_U23 (.A( u2_u4_u6_n123 ) , .ZN( u2_u4_u6_n170 ) );
  INV_X1 u2_u4_u6_U24 (.A( u2_u4_u6_n113 ) , .ZN( u2_u4_u6_n168 ) );
  AND2_X1 u2_u4_u6_U25 (.A1( u2_u4_u6_n107 ) , .A2( u2_u4_u6_n119 ) , .ZN( u2_u4_u6_n133 ) );
  AND2_X1 u2_u4_u6_U26 (.A2( u2_u4_u6_n121 ) , .A1( u2_u4_u6_n122 ) , .ZN( u2_u4_u6_n131 ) );
  AND3_X1 u2_u4_u6_U27 (.ZN( u2_u4_u6_n120 ) , .A2( u2_u4_u6_n127 ) , .A1( u2_u4_u6_n132 ) , .A3( u2_u4_u6_n145 ) );
  INV_X1 u2_u4_u6_U28 (.A( u2_u4_u6_n146 ) , .ZN( u2_u4_u6_n163 ) );
  AOI222_X1 u2_u4_u6_U29 (.ZN( u2_u4_u6_n114 ) , .A1( u2_u4_u6_n118 ) , .A2( u2_u4_u6_n126 ) , .B2( u2_u4_u6_n151 ) , .C2( u2_u4_u6_n159 ) , .C1( u2_u4_u6_n168 ) , .B1( u2_u4_u6_n169 ) );
  INV_X1 u2_u4_u6_U3 (.A( u2_u4_u6_n110 ) , .ZN( u2_u4_u6_n166 ) );
  NOR2_X1 u2_u4_u6_U30 (.A1( u2_u4_u6_n162 ) , .A2( u2_u4_u6_n165 ) , .ZN( u2_u4_u6_n98 ) );
  NAND2_X1 u2_u4_u6_U31 (.A1( u2_u4_u6_n144 ) , .ZN( u2_u4_u6_n151 ) , .A2( u2_u4_u6_n158 ) );
  NAND2_X1 u2_u4_u6_U32 (.ZN( u2_u4_u6_n132 ) , .A1( u2_u4_u6_n91 ) , .A2( u2_u4_u6_n97 ) );
  AOI22_X1 u2_u4_u6_U33 (.B2( u2_u4_u6_n110 ) , .B1( u2_u4_u6_n111 ) , .A1( u2_u4_u6_n112 ) , .ZN( u2_u4_u6_n115 ) , .A2( u2_u4_u6_n161 ) );
  NAND4_X1 u2_u4_u6_U34 (.A3( u2_u4_u6_n109 ) , .ZN( u2_u4_u6_n112 ) , .A4( u2_u4_u6_n132 ) , .A2( u2_u4_u6_n147 ) , .A1( u2_u4_u6_n166 ) );
  NOR2_X1 u2_u4_u6_U35 (.ZN( u2_u4_u6_n109 ) , .A1( u2_u4_u6_n170 ) , .A2( u2_u4_u6_n173 ) );
  NOR2_X1 u2_u4_u6_U36 (.A2( u2_u4_u6_n126 ) , .ZN( u2_u4_u6_n155 ) , .A1( u2_u4_u6_n160 ) );
  NAND2_X1 u2_u4_u6_U37 (.ZN( u2_u4_u6_n146 ) , .A2( u2_u4_u6_n94 ) , .A1( u2_u4_u6_n99 ) );
  AOI21_X1 u2_u4_u6_U38 (.A( u2_u4_u6_n144 ) , .B2( u2_u4_u6_n145 ) , .B1( u2_u4_u6_n146 ) , .ZN( u2_u4_u6_n150 ) );
  AOI211_X1 u2_u4_u6_U39 (.B( u2_u4_u6_n134 ) , .A( u2_u4_u6_n135 ) , .C1( u2_u4_u6_n136 ) , .ZN( u2_u4_u6_n137 ) , .C2( u2_u4_u6_n151 ) );
  INV_X1 u2_u4_u6_U4 (.A( u2_u4_u6_n142 ) , .ZN( u2_u4_u6_n174 ) );
  NAND4_X1 u2_u4_u6_U40 (.A4( u2_u4_u6_n127 ) , .A3( u2_u4_u6_n128 ) , .A2( u2_u4_u6_n129 ) , .A1( u2_u4_u6_n130 ) , .ZN( u2_u4_u6_n136 ) );
  AOI21_X1 u2_u4_u6_U41 (.B2( u2_u4_u6_n132 ) , .B1( u2_u4_u6_n133 ) , .ZN( u2_u4_u6_n134 ) , .A( u2_u4_u6_n158 ) );
  AOI21_X1 u2_u4_u6_U42 (.B1( u2_u4_u6_n131 ) , .ZN( u2_u4_u6_n135 ) , .A( u2_u4_u6_n144 ) , .B2( u2_u4_u6_n146 ) );
  INV_X1 u2_u4_u6_U43 (.A( u2_u4_u6_n111 ) , .ZN( u2_u4_u6_n158 ) );
  NAND2_X1 u2_u4_u6_U44 (.ZN( u2_u4_u6_n127 ) , .A1( u2_u4_u6_n91 ) , .A2( u2_u4_u6_n92 ) );
  NAND2_X1 u2_u4_u6_U45 (.ZN( u2_u4_u6_n129 ) , .A2( u2_u4_u6_n95 ) , .A1( u2_u4_u6_n96 ) );
  INV_X1 u2_u4_u6_U46 (.A( u2_u4_u6_n144 ) , .ZN( u2_u4_u6_n159 ) );
  NAND2_X1 u2_u4_u6_U47 (.ZN( u2_u4_u6_n145 ) , .A2( u2_u4_u6_n97 ) , .A1( u2_u4_u6_n98 ) );
  NAND2_X1 u2_u4_u6_U48 (.ZN( u2_u4_u6_n148 ) , .A2( u2_u4_u6_n92 ) , .A1( u2_u4_u6_n94 ) );
  NAND2_X1 u2_u4_u6_U49 (.ZN( u2_u4_u6_n108 ) , .A2( u2_u4_u6_n139 ) , .A1( u2_u4_u6_n144 ) );
  NAND2_X1 u2_u4_u6_U5 (.A2( u2_u4_u6_n143 ) , .ZN( u2_u4_u6_n152 ) , .A1( u2_u4_u6_n166 ) );
  NAND2_X1 u2_u4_u6_U50 (.ZN( u2_u4_u6_n121 ) , .A2( u2_u4_u6_n95 ) , .A1( u2_u4_u6_n97 ) );
  NAND2_X1 u2_u4_u6_U51 (.ZN( u2_u4_u6_n107 ) , .A2( u2_u4_u6_n92 ) , .A1( u2_u4_u6_n95 ) );
  AND2_X1 u2_u4_u6_U52 (.ZN( u2_u4_u6_n118 ) , .A2( u2_u4_u6_n91 ) , .A1( u2_u4_u6_n99 ) );
  NAND2_X1 u2_u4_u6_U53 (.ZN( u2_u4_u6_n147 ) , .A2( u2_u4_u6_n98 ) , .A1( u2_u4_u6_n99 ) );
  NAND2_X1 u2_u4_u6_U54 (.ZN( u2_u4_u6_n128 ) , .A1( u2_u4_u6_n94 ) , .A2( u2_u4_u6_n96 ) );
  NAND2_X1 u2_u4_u6_U55 (.ZN( u2_u4_u6_n119 ) , .A2( u2_u4_u6_n95 ) , .A1( u2_u4_u6_n99 ) );
  NAND2_X1 u2_u4_u6_U56 (.ZN( u2_u4_u6_n123 ) , .A2( u2_u4_u6_n91 ) , .A1( u2_u4_u6_n96 ) );
  NAND2_X1 u2_u4_u6_U57 (.ZN( u2_u4_u6_n100 ) , .A2( u2_u4_u6_n92 ) , .A1( u2_u4_u6_n98 ) );
  NAND2_X1 u2_u4_u6_U58 (.ZN( u2_u4_u6_n122 ) , .A1( u2_u4_u6_n94 ) , .A2( u2_u4_u6_n97 ) );
  INV_X1 u2_u4_u6_U59 (.A( u2_u4_u6_n139 ) , .ZN( u2_u4_u6_n160 ) );
  AOI22_X1 u2_u4_u6_U6 (.B2( u2_u4_u6_n101 ) , .A1( u2_u4_u6_n102 ) , .ZN( u2_u4_u6_n103 ) , .B1( u2_u4_u6_n160 ) , .A2( u2_u4_u6_n161 ) );
  NAND2_X1 u2_u4_u6_U60 (.ZN( u2_u4_u6_n113 ) , .A1( u2_u4_u6_n96 ) , .A2( u2_u4_u6_n98 ) );
  NOR2_X1 u2_u4_u6_U61 (.A2( u2_u4_X_40 ) , .A1( u2_u4_X_41 ) , .ZN( u2_u4_u6_n126 ) );
  NOR2_X1 u2_u4_u6_U62 (.A2( u2_u4_X_39 ) , .A1( u2_u4_X_42 ) , .ZN( u2_u4_u6_n92 ) );
  NOR2_X1 u2_u4_u6_U63 (.A2( u2_u4_X_39 ) , .A1( u2_u4_u6_n156 ) , .ZN( u2_u4_u6_n97 ) );
  NOR2_X1 u2_u4_u6_U64 (.A2( u2_u4_X_38 ) , .A1( u2_u4_u6_n165 ) , .ZN( u2_u4_u6_n95 ) );
  NOR2_X1 u2_u4_u6_U65 (.A2( u2_u4_X_41 ) , .ZN( u2_u4_u6_n111 ) , .A1( u2_u4_u6_n157 ) );
  NOR2_X1 u2_u4_u6_U66 (.A2( u2_u4_X_37 ) , .A1( u2_u4_u6_n162 ) , .ZN( u2_u4_u6_n94 ) );
  NOR2_X1 u2_u4_u6_U67 (.A2( u2_u4_X_37 ) , .A1( u2_u4_X_38 ) , .ZN( u2_u4_u6_n91 ) );
  NAND2_X1 u2_u4_u6_U68 (.A1( u2_u4_X_41 ) , .ZN( u2_u4_u6_n144 ) , .A2( u2_u4_u6_n157 ) );
  NAND2_X1 u2_u4_u6_U69 (.A2( u2_u4_X_40 ) , .A1( u2_u4_X_41 ) , .ZN( u2_u4_u6_n139 ) );
  NOR2_X1 u2_u4_u6_U7 (.A1( u2_u4_u6_n118 ) , .ZN( u2_u4_u6_n143 ) , .A2( u2_u4_u6_n168 ) );
  AND2_X1 u2_u4_u6_U70 (.A1( u2_u4_X_39 ) , .A2( u2_u4_u6_n156 ) , .ZN( u2_u4_u6_n96 ) );
  AND2_X1 u2_u4_u6_U71 (.A1( u2_u4_X_39 ) , .A2( u2_u4_X_42 ) , .ZN( u2_u4_u6_n99 ) );
  INV_X1 u2_u4_u6_U72 (.A( u2_u4_X_40 ) , .ZN( u2_u4_u6_n157 ) );
  INV_X1 u2_u4_u6_U73 (.A( u2_u4_X_37 ) , .ZN( u2_u4_u6_n165 ) );
  INV_X1 u2_u4_u6_U74 (.A( u2_u4_X_38 ) , .ZN( u2_u4_u6_n162 ) );
  INV_X1 u2_u4_u6_U75 (.A( u2_u4_X_42 ) , .ZN( u2_u4_u6_n156 ) );
  NAND4_X1 u2_u4_u6_U76 (.ZN( u2_out4_32 ) , .A4( u2_u4_u6_n103 ) , .A3( u2_u4_u6_n104 ) , .A2( u2_u4_u6_n105 ) , .A1( u2_u4_u6_n106 ) );
  AOI22_X1 u2_u4_u6_U77 (.ZN( u2_u4_u6_n105 ) , .A2( u2_u4_u6_n108 ) , .A1( u2_u4_u6_n118 ) , .B2( u2_u4_u6_n126 ) , .B1( u2_u4_u6_n171 ) );
  AOI22_X1 u2_u4_u6_U78 (.ZN( u2_u4_u6_n104 ) , .A1( u2_u4_u6_n111 ) , .B1( u2_u4_u6_n124 ) , .B2( u2_u4_u6_n151 ) , .A2( u2_u4_u6_n93 ) );
  NAND4_X1 u2_u4_u6_U79 (.ZN( u2_out4_12 ) , .A4( u2_u4_u6_n114 ) , .A3( u2_u4_u6_n115 ) , .A2( u2_u4_u6_n116 ) , .A1( u2_u4_u6_n117 ) );
  INV_X1 u2_u4_u6_U8 (.ZN( u2_u4_u6_n172 ) , .A( u2_u4_u6_n88 ) );
  OAI22_X1 u2_u4_u6_U80 (.B2( u2_u4_u6_n111 ) , .ZN( u2_u4_u6_n116 ) , .B1( u2_u4_u6_n126 ) , .A2( u2_u4_u6_n164 ) , .A1( u2_u4_u6_n167 ) );
  OAI21_X1 u2_u4_u6_U81 (.A( u2_u4_u6_n108 ) , .ZN( u2_u4_u6_n117 ) , .B2( u2_u4_u6_n141 ) , .B1( u2_u4_u6_n163 ) );
  OAI211_X1 u2_u4_u6_U82 (.ZN( u2_out4_22 ) , .B( u2_u4_u6_n137 ) , .A( u2_u4_u6_n138 ) , .C2( u2_u4_u6_n139 ) , .C1( u2_u4_u6_n140 ) );
  AOI22_X1 u2_u4_u6_U83 (.B1( u2_u4_u6_n124 ) , .A2( u2_u4_u6_n125 ) , .A1( u2_u4_u6_n126 ) , .ZN( u2_u4_u6_n138 ) , .B2( u2_u4_u6_n161 ) );
  AND4_X1 u2_u4_u6_U84 (.A3( u2_u4_u6_n119 ) , .A1( u2_u4_u6_n120 ) , .A4( u2_u4_u6_n129 ) , .ZN( u2_u4_u6_n140 ) , .A2( u2_u4_u6_n143 ) );
  OAI211_X1 u2_u4_u6_U85 (.ZN( u2_out4_7 ) , .B( u2_u4_u6_n153 ) , .C2( u2_u4_u6_n154 ) , .C1( u2_u4_u6_n155 ) , .A( u2_u4_u6_n174 ) );
  NOR3_X1 u2_u4_u6_U86 (.A1( u2_u4_u6_n141 ) , .ZN( u2_u4_u6_n154 ) , .A3( u2_u4_u6_n164 ) , .A2( u2_u4_u6_n171 ) );
  AOI211_X1 u2_u4_u6_U87 (.B( u2_u4_u6_n149 ) , .A( u2_u4_u6_n150 ) , .C2( u2_u4_u6_n151 ) , .C1( u2_u4_u6_n152 ) , .ZN( u2_u4_u6_n153 ) );
  NAND3_X1 u2_u4_u6_U88 (.A2( u2_u4_u6_n123 ) , .ZN( u2_u4_u6_n125 ) , .A1( u2_u4_u6_n130 ) , .A3( u2_u4_u6_n131 ) );
  NAND3_X1 u2_u4_u6_U89 (.A3( u2_u4_u6_n133 ) , .ZN( u2_u4_u6_n141 ) , .A1( u2_u4_u6_n145 ) , .A2( u2_u4_u6_n148 ) );
  OAI21_X1 u2_u4_u6_U9 (.A( u2_u4_u6_n159 ) , .B1( u2_u4_u6_n169 ) , .B2( u2_u4_u6_n173 ) , .ZN( u2_u4_u6_n90 ) );
  NAND3_X1 u2_u4_u6_U90 (.ZN( u2_u4_u6_n101 ) , .A3( u2_u4_u6_n107 ) , .A2( u2_u4_u6_n121 ) , .A1( u2_u4_u6_n127 ) );
  NAND3_X1 u2_u4_u6_U91 (.ZN( u2_u4_u6_n102 ) , .A3( u2_u4_u6_n130 ) , .A2( u2_u4_u6_n145 ) , .A1( u2_u4_u6_n166 ) );
  NAND3_X1 u2_u4_u6_U92 (.A3( u2_u4_u6_n113 ) , .A1( u2_u4_u6_n119 ) , .A2( u2_u4_u6_n123 ) , .ZN( u2_u4_u6_n93 ) );
  NAND3_X1 u2_u4_u6_U93 (.ZN( u2_u4_u6_n142 ) , .A2( u2_u4_u6_n172 ) , .A3( u2_u4_u6_n89 ) , .A1( u2_u4_u6_n90 ) );
  XOR2_X1 u2_u7_U10 (.B( u2_K8_45 ) , .A( u2_R6_30 ) , .Z( u2_u7_X_45 ) );
  XOR2_X1 u2_u7_U11 (.B( u2_K8_44 ) , .A( u2_R6_29 ) , .Z( u2_u7_X_44 ) );
  XOR2_X1 u2_u7_U12 (.B( u2_K8_43 ) , .A( u2_R6_28 ) , .Z( u2_u7_X_43 ) );
  XOR2_X1 u2_u7_U7 (.B( u2_K8_48 ) , .A( u2_R6_1 ) , .Z( u2_u7_X_48 ) );
  XOR2_X1 u2_u7_U8 (.B( u2_K8_47 ) , .A( u2_R6_32 ) , .Z( u2_u7_X_47 ) );
  XOR2_X1 u2_u7_U9 (.B( u2_K8_46 ) , .A( u2_R6_31 ) , .Z( u2_u7_X_46 ) );
  OAI21_X1 u2_u7_u7_U10 (.A( u2_u7_u7_n161 ) , .B1( u2_u7_u7_n168 ) , .B2( u2_u7_u7_n173 ) , .ZN( u2_u7_u7_n91 ) );
  AOI211_X1 u2_u7_u7_U11 (.A( u2_u7_u7_n117 ) , .ZN( u2_u7_u7_n118 ) , .C2( u2_u7_u7_n126 ) , .C1( u2_u7_u7_n177 ) , .B( u2_u7_u7_n180 ) );
  OAI22_X1 u2_u7_u7_U12 (.B1( u2_u7_u7_n115 ) , .ZN( u2_u7_u7_n117 ) , .A2( u2_u7_u7_n133 ) , .A1( u2_u7_u7_n137 ) , .B2( u2_u7_u7_n162 ) );
  INV_X1 u2_u7_u7_U13 (.A( u2_u7_u7_n116 ) , .ZN( u2_u7_u7_n180 ) );
  NOR3_X1 u2_u7_u7_U14 (.ZN( u2_u7_u7_n115 ) , .A3( u2_u7_u7_n145 ) , .A2( u2_u7_u7_n168 ) , .A1( u2_u7_u7_n169 ) );
  INV_X1 u2_u7_u7_U15 (.A( u2_u7_u7_n133 ) , .ZN( u2_u7_u7_n176 ) );
  NOR3_X1 u2_u7_u7_U16 (.A2( u2_u7_u7_n134 ) , .A1( u2_u7_u7_n135 ) , .ZN( u2_u7_u7_n136 ) , .A3( u2_u7_u7_n171 ) );
  NOR2_X1 u2_u7_u7_U17 (.A1( u2_u7_u7_n130 ) , .A2( u2_u7_u7_n134 ) , .ZN( u2_u7_u7_n153 ) );
  AOI21_X1 u2_u7_u7_U18 (.ZN( u2_u7_u7_n104 ) , .B2( u2_u7_u7_n112 ) , .B1( u2_u7_u7_n127 ) , .A( u2_u7_u7_n164 ) );
  AOI21_X1 u2_u7_u7_U19 (.ZN( u2_u7_u7_n106 ) , .B1( u2_u7_u7_n133 ) , .B2( u2_u7_u7_n146 ) , .A( u2_u7_u7_n162 ) );
  AOI21_X1 u2_u7_u7_U20 (.A( u2_u7_u7_n101 ) , .ZN( u2_u7_u7_n107 ) , .B2( u2_u7_u7_n128 ) , .B1( u2_u7_u7_n175 ) );
  INV_X1 u2_u7_u7_U21 (.A( u2_u7_u7_n101 ) , .ZN( u2_u7_u7_n165 ) );
  NOR2_X1 u2_u7_u7_U22 (.ZN( u2_u7_u7_n111 ) , .A2( u2_u7_u7_n134 ) , .A1( u2_u7_u7_n169 ) );
  INV_X1 u2_u7_u7_U23 (.A( u2_u7_u7_n138 ) , .ZN( u2_u7_u7_n171 ) );
  INV_X1 u2_u7_u7_U24 (.A( u2_u7_u7_n131 ) , .ZN( u2_u7_u7_n177 ) );
  INV_X1 u2_u7_u7_U25 (.A( u2_u7_u7_n110 ) , .ZN( u2_u7_u7_n174 ) );
  NAND2_X1 u2_u7_u7_U26 (.A1( u2_u7_u7_n129 ) , .A2( u2_u7_u7_n132 ) , .ZN( u2_u7_u7_n149 ) );
  NAND2_X1 u2_u7_u7_U27 (.A1( u2_u7_u7_n113 ) , .A2( u2_u7_u7_n124 ) , .ZN( u2_u7_u7_n130 ) );
  INV_X1 u2_u7_u7_U28 (.A( u2_u7_u7_n112 ) , .ZN( u2_u7_u7_n173 ) );
  INV_X1 u2_u7_u7_U29 (.A( u2_u7_u7_n128 ) , .ZN( u2_u7_u7_n168 ) );
  OAI21_X1 u2_u7_u7_U3 (.ZN( u2_u7_u7_n159 ) , .A( u2_u7_u7_n165 ) , .B2( u2_u7_u7_n171 ) , .B1( u2_u7_u7_n174 ) );
  INV_X1 u2_u7_u7_U30 (.A( u2_u7_u7_n148 ) , .ZN( u2_u7_u7_n169 ) );
  INV_X1 u2_u7_u7_U31 (.A( u2_u7_u7_n127 ) , .ZN( u2_u7_u7_n179 ) );
  NOR2_X1 u2_u7_u7_U32 (.ZN( u2_u7_u7_n101 ) , .A2( u2_u7_u7_n150 ) , .A1( u2_u7_u7_n156 ) );
  AOI211_X1 u2_u7_u7_U33 (.B( u2_u7_u7_n139 ) , .A( u2_u7_u7_n140 ) , .C2( u2_u7_u7_n141 ) , .ZN( u2_u7_u7_n142 ) , .C1( u2_u7_u7_n156 ) );
  NAND4_X1 u2_u7_u7_U34 (.A3( u2_u7_u7_n127 ) , .A2( u2_u7_u7_n128 ) , .A1( u2_u7_u7_n129 ) , .ZN( u2_u7_u7_n141 ) , .A4( u2_u7_u7_n147 ) );
  AOI21_X1 u2_u7_u7_U35 (.A( u2_u7_u7_n137 ) , .B1( u2_u7_u7_n138 ) , .ZN( u2_u7_u7_n139 ) , .B2( u2_u7_u7_n146 ) );
  OAI22_X1 u2_u7_u7_U36 (.B1( u2_u7_u7_n136 ) , .ZN( u2_u7_u7_n140 ) , .A1( u2_u7_u7_n153 ) , .B2( u2_u7_u7_n162 ) , .A2( u2_u7_u7_n164 ) );
  INV_X1 u2_u7_u7_U37 (.A( u2_u7_u7_n125 ) , .ZN( u2_u7_u7_n161 ) );
  AOI21_X1 u2_u7_u7_U38 (.ZN( u2_u7_u7_n123 ) , .B1( u2_u7_u7_n165 ) , .B2( u2_u7_u7_n177 ) , .A( u2_u7_u7_n97 ) );
  AOI21_X1 u2_u7_u7_U39 (.B2( u2_u7_u7_n113 ) , .B1( u2_u7_u7_n124 ) , .A( u2_u7_u7_n125 ) , .ZN( u2_u7_u7_n97 ) );
  INV_X1 u2_u7_u7_U4 (.A( u2_u7_u7_n149 ) , .ZN( u2_u7_u7_n175 ) );
  INV_X1 u2_u7_u7_U40 (.A( u2_u7_u7_n152 ) , .ZN( u2_u7_u7_n162 ) );
  AOI22_X1 u2_u7_u7_U41 (.A2( u2_u7_u7_n114 ) , .ZN( u2_u7_u7_n119 ) , .B1( u2_u7_u7_n130 ) , .A1( u2_u7_u7_n156 ) , .B2( u2_u7_u7_n165 ) );
  NAND2_X1 u2_u7_u7_U42 (.A2( u2_u7_u7_n112 ) , .ZN( u2_u7_u7_n114 ) , .A1( u2_u7_u7_n175 ) );
  NOR2_X1 u2_u7_u7_U43 (.ZN( u2_u7_u7_n137 ) , .A1( u2_u7_u7_n150 ) , .A2( u2_u7_u7_n161 ) );
  AND2_X1 u2_u7_u7_U44 (.ZN( u2_u7_u7_n145 ) , .A2( u2_u7_u7_n98 ) , .A1( u2_u7_u7_n99 ) );
  AOI21_X1 u2_u7_u7_U45 (.ZN( u2_u7_u7_n105 ) , .B2( u2_u7_u7_n110 ) , .A( u2_u7_u7_n125 ) , .B1( u2_u7_u7_n147 ) );
  NAND2_X1 u2_u7_u7_U46 (.ZN( u2_u7_u7_n146 ) , .A1( u2_u7_u7_n95 ) , .A2( u2_u7_u7_n98 ) );
  NAND2_X1 u2_u7_u7_U47 (.A2( u2_u7_u7_n103 ) , .ZN( u2_u7_u7_n147 ) , .A1( u2_u7_u7_n93 ) );
  NAND2_X1 u2_u7_u7_U48 (.A1( u2_u7_u7_n103 ) , .ZN( u2_u7_u7_n127 ) , .A2( u2_u7_u7_n99 ) );
  NAND2_X1 u2_u7_u7_U49 (.A2( u2_u7_u7_n102 ) , .A1( u2_u7_u7_n103 ) , .ZN( u2_u7_u7_n133 ) );
  INV_X1 u2_u7_u7_U5 (.A( u2_u7_u7_n154 ) , .ZN( u2_u7_u7_n178 ) );
  OR2_X1 u2_u7_u7_U50 (.ZN( u2_u7_u7_n126 ) , .A2( u2_u7_u7_n152 ) , .A1( u2_u7_u7_n156 ) );
  NAND2_X1 u2_u7_u7_U51 (.ZN( u2_u7_u7_n112 ) , .A2( u2_u7_u7_n96 ) , .A1( u2_u7_u7_n99 ) );
  NAND2_X1 u2_u7_u7_U52 (.A2( u2_u7_u7_n102 ) , .ZN( u2_u7_u7_n128 ) , .A1( u2_u7_u7_n98 ) );
  NAND2_X1 u2_u7_u7_U53 (.A1( u2_u7_u7_n100 ) , .ZN( u2_u7_u7_n113 ) , .A2( u2_u7_u7_n93 ) );
  NAND2_X1 u2_u7_u7_U54 (.ZN( u2_u7_u7_n110 ) , .A1( u2_u7_u7_n95 ) , .A2( u2_u7_u7_n96 ) );
  INV_X1 u2_u7_u7_U55 (.A( u2_u7_u7_n150 ) , .ZN( u2_u7_u7_n164 ) );
  AND2_X1 u2_u7_u7_U56 (.ZN( u2_u7_u7_n134 ) , .A1( u2_u7_u7_n93 ) , .A2( u2_u7_u7_n98 ) );
  NAND2_X1 u2_u7_u7_U57 (.A2( u2_u7_u7_n102 ) , .ZN( u2_u7_u7_n124 ) , .A1( u2_u7_u7_n96 ) );
  NAND2_X1 u2_u7_u7_U58 (.A1( u2_u7_u7_n100 ) , .A2( u2_u7_u7_n102 ) , .ZN( u2_u7_u7_n129 ) );
  NAND2_X1 u2_u7_u7_U59 (.A2( u2_u7_u7_n103 ) , .ZN( u2_u7_u7_n131 ) , .A1( u2_u7_u7_n95 ) );
  AOI211_X1 u2_u7_u7_U6 (.ZN( u2_u7_u7_n116 ) , .A( u2_u7_u7_n155 ) , .C1( u2_u7_u7_n161 ) , .C2( u2_u7_u7_n171 ) , .B( u2_u7_u7_n94 ) );
  NAND2_X1 u2_u7_u7_U60 (.A1( u2_u7_u7_n100 ) , .ZN( u2_u7_u7_n138 ) , .A2( u2_u7_u7_n99 ) );
  NAND2_X1 u2_u7_u7_U61 (.ZN( u2_u7_u7_n132 ) , .A1( u2_u7_u7_n93 ) , .A2( u2_u7_u7_n96 ) );
  NAND2_X1 u2_u7_u7_U62 (.A1( u2_u7_u7_n100 ) , .ZN( u2_u7_u7_n148 ) , .A2( u2_u7_u7_n95 ) );
  AOI211_X1 u2_u7_u7_U63 (.B( u2_u7_u7_n154 ) , .A( u2_u7_u7_n155 ) , .C1( u2_u7_u7_n156 ) , .ZN( u2_u7_u7_n157 ) , .C2( u2_u7_u7_n172 ) );
  INV_X1 u2_u7_u7_U64 (.A( u2_u7_u7_n153 ) , .ZN( u2_u7_u7_n172 ) );
  NOR2_X1 u2_u7_u7_U65 (.A2( u2_u7_X_47 ) , .ZN( u2_u7_u7_n150 ) , .A1( u2_u7_u7_n163 ) );
  NOR2_X1 u2_u7_u7_U66 (.A2( u2_u7_X_43 ) , .A1( u2_u7_X_44 ) , .ZN( u2_u7_u7_n103 ) );
  NOR2_X1 u2_u7_u7_U67 (.A2( u2_u7_X_48 ) , .A1( u2_u7_u7_n166 ) , .ZN( u2_u7_u7_n95 ) );
  NOR2_X1 u2_u7_u7_U68 (.A2( u2_u7_X_45 ) , .A1( u2_u7_X_48 ) , .ZN( u2_u7_u7_n99 ) );
  NOR2_X1 u2_u7_u7_U69 (.A2( u2_u7_X_44 ) , .A1( u2_u7_u7_n167 ) , .ZN( u2_u7_u7_n98 ) );
  OAI222_X1 u2_u7_u7_U7 (.C2( u2_u7_u7_n101 ) , .B2( u2_u7_u7_n111 ) , .A1( u2_u7_u7_n113 ) , .C1( u2_u7_u7_n146 ) , .A2( u2_u7_u7_n162 ) , .B1( u2_u7_u7_n164 ) , .ZN( u2_u7_u7_n94 ) );
  NOR2_X1 u2_u7_u7_U70 (.A2( u2_u7_X_46 ) , .A1( u2_u7_X_47 ) , .ZN( u2_u7_u7_n152 ) );
  NAND2_X1 u2_u7_u7_U71 (.A2( u2_u7_X_46 ) , .A1( u2_u7_X_47 ) , .ZN( u2_u7_u7_n125 ) );
  AND2_X1 u2_u7_u7_U72 (.A1( u2_u7_X_47 ) , .ZN( u2_u7_u7_n156 ) , .A2( u2_u7_u7_n163 ) );
  AND2_X1 u2_u7_u7_U73 (.A2( u2_u7_X_45 ) , .A1( u2_u7_X_48 ) , .ZN( u2_u7_u7_n102 ) );
  AND2_X1 u2_u7_u7_U74 (.A2( u2_u7_X_43 ) , .A1( u2_u7_X_44 ) , .ZN( u2_u7_u7_n96 ) );
  AND2_X1 u2_u7_u7_U75 (.A1( u2_u7_X_44 ) , .ZN( u2_u7_u7_n100 ) , .A2( u2_u7_u7_n167 ) );
  AND2_X1 u2_u7_u7_U76 (.A1( u2_u7_X_48 ) , .A2( u2_u7_u7_n166 ) , .ZN( u2_u7_u7_n93 ) );
  INV_X1 u2_u7_u7_U77 (.A( u2_u7_X_46 ) , .ZN( u2_u7_u7_n163 ) );
  INV_X1 u2_u7_u7_U78 (.A( u2_u7_X_43 ) , .ZN( u2_u7_u7_n167 ) );
  INV_X1 u2_u7_u7_U79 (.A( u2_u7_X_45 ) , .ZN( u2_u7_u7_n166 ) );
  OAI221_X1 u2_u7_u7_U8 (.C1( u2_u7_u7_n101 ) , .C2( u2_u7_u7_n147 ) , .ZN( u2_u7_u7_n155 ) , .B2( u2_u7_u7_n162 ) , .A( u2_u7_u7_n91 ) , .B1( u2_u7_u7_n92 ) );
  NAND4_X1 u2_u7_u7_U80 (.ZN( u2_out7_5 ) , .A4( u2_u7_u7_n108 ) , .A3( u2_u7_u7_n109 ) , .A1( u2_u7_u7_n116 ) , .A2( u2_u7_u7_n123 ) );
  AOI22_X1 u2_u7_u7_U81 (.ZN( u2_u7_u7_n109 ) , .A2( u2_u7_u7_n126 ) , .B2( u2_u7_u7_n145 ) , .B1( u2_u7_u7_n156 ) , .A1( u2_u7_u7_n171 ) );
  NOR4_X1 u2_u7_u7_U82 (.A4( u2_u7_u7_n104 ) , .A3( u2_u7_u7_n105 ) , .A2( u2_u7_u7_n106 ) , .A1( u2_u7_u7_n107 ) , .ZN( u2_u7_u7_n108 ) );
  NAND4_X1 u2_u7_u7_U83 (.ZN( u2_out7_27 ) , .A4( u2_u7_u7_n118 ) , .A3( u2_u7_u7_n119 ) , .A2( u2_u7_u7_n120 ) , .A1( u2_u7_u7_n121 ) );
  OAI21_X1 u2_u7_u7_U84 (.ZN( u2_u7_u7_n121 ) , .B2( u2_u7_u7_n145 ) , .A( u2_u7_u7_n150 ) , .B1( u2_u7_u7_n174 ) );
  OAI21_X1 u2_u7_u7_U85 (.ZN( u2_u7_u7_n120 ) , .A( u2_u7_u7_n161 ) , .B2( u2_u7_u7_n170 ) , .B1( u2_u7_u7_n179 ) );
  NAND4_X1 u2_u7_u7_U86 (.ZN( u2_out7_21 ) , .A4( u2_u7_u7_n157 ) , .A3( u2_u7_u7_n158 ) , .A2( u2_u7_u7_n159 ) , .A1( u2_u7_u7_n160 ) );
  OAI21_X1 u2_u7_u7_U87 (.B1( u2_u7_u7_n145 ) , .ZN( u2_u7_u7_n160 ) , .A( u2_u7_u7_n161 ) , .B2( u2_u7_u7_n177 ) );
  AOI22_X1 u2_u7_u7_U88 (.B2( u2_u7_u7_n149 ) , .B1( u2_u7_u7_n150 ) , .A2( u2_u7_u7_n151 ) , .A1( u2_u7_u7_n152 ) , .ZN( u2_u7_u7_n158 ) );
  NAND4_X1 u2_u7_u7_U89 (.ZN( u2_out7_15 ) , .A4( u2_u7_u7_n142 ) , .A3( u2_u7_u7_n143 ) , .A2( u2_u7_u7_n144 ) , .A1( u2_u7_u7_n178 ) );
  AND3_X1 u2_u7_u7_U9 (.A3( u2_u7_u7_n110 ) , .A2( u2_u7_u7_n127 ) , .A1( u2_u7_u7_n132 ) , .ZN( u2_u7_u7_n92 ) );
  OR2_X1 u2_u7_u7_U90 (.A2( u2_u7_u7_n125 ) , .A1( u2_u7_u7_n129 ) , .ZN( u2_u7_u7_n144 ) );
  AOI22_X1 u2_u7_u7_U91 (.A2( u2_u7_u7_n126 ) , .ZN( u2_u7_u7_n143 ) , .B2( u2_u7_u7_n165 ) , .B1( u2_u7_u7_n173 ) , .A1( u2_u7_u7_n174 ) );
  OAI211_X1 u2_u7_u7_U92 (.B( u2_u7_u7_n122 ) , .A( u2_u7_u7_n123 ) , .C2( u2_u7_u7_n124 ) , .ZN( u2_u7_u7_n154 ) , .C1( u2_u7_u7_n162 ) );
  AOI222_X1 u2_u7_u7_U93 (.ZN( u2_u7_u7_n122 ) , .C2( u2_u7_u7_n126 ) , .C1( u2_u7_u7_n145 ) , .B1( u2_u7_u7_n161 ) , .A2( u2_u7_u7_n165 ) , .B2( u2_u7_u7_n170 ) , .A1( u2_u7_u7_n176 ) );
  INV_X1 u2_u7_u7_U94 (.A( u2_u7_u7_n111 ) , .ZN( u2_u7_u7_n170 ) );
  NAND3_X1 u2_u7_u7_U95 (.A3( u2_u7_u7_n146 ) , .A2( u2_u7_u7_n147 ) , .A1( u2_u7_u7_n148 ) , .ZN( u2_u7_u7_n151 ) );
  NAND3_X1 u2_u7_u7_U96 (.A3( u2_u7_u7_n131 ) , .A2( u2_u7_u7_n132 ) , .A1( u2_u7_u7_n133 ) , .ZN( u2_u7_u7_n135 ) );
  OAI21_X1 u2_uk_U1015 (.ZN( u2_K8_46 ) , .A( u2_uk_n1115 ) , .B2( u2_uk_n1532 ) , .B1( u2_uk_n182 ) );
  NAND2_X1 u2_uk_U1016 (.A1( u2_uk_K_r6_37 ) , .ZN( u2_uk_n1115 ) , .A2( u2_uk_n155 ) );
  OAI21_X1 u2_uk_U1037 (.ZN( u2_K5_42 ) , .A( u2_uk_n1052 ) , .B2( u2_uk_n1382 ) , .B1( u2_uk_n17 ) );
  NAND2_X1 u2_uk_U1038 (.A1( u2_uk_K_r3_9 ) , .ZN( u2_uk_n1052 ) , .A2( u2_uk_n60 ) );
  OAI21_X1 u2_uk_U1078 (.ZN( u2_K5_39 ) , .A( u2_uk_n1051 ) , .B2( u2_uk_n1376 ) , .B1( u2_uk_n162 ) );
  NAND2_X1 u2_uk_U1079 (.A1( u2_uk_K_r3_16 ) , .ZN( u2_uk_n1051 ) , .A2( u2_uk_n155 ) );
  INV_X1 u2_uk_U1126 (.ZN( u2_K5_35 ) , .A( u2_uk_n1049 ) );
  INV_X1 u2_uk_U1139 (.ZN( u2_K8_43 ) , .A( u2_uk_n1113 ) );
  OAI22_X1 u2_uk_U116 (.ZN( u2_K8_47 ) , .B2( u2_uk_n1531 ) , .A2( u2_uk_n1537 ) , .B1( u2_uk_n17 ) , .A1( u2_uk_n223 ) );
  INV_X1 u2_uk_U156 (.ZN( u2_K2_19 ) , .A( u2_uk_n995 ) );
  AOI22_X1 u2_uk_U157 (.B2( u2_uk_K_r0_11 ) , .A2( u2_uk_K_r0_47 ) , .A1( u2_uk_n128 ) , .B1( u2_uk_n231 ) , .ZN( u2_uk_n995 ) );
  OAI21_X1 u2_uk_U264 (.ZN( u2_K8_44 ) , .B1( u2_uk_n102 ) , .A( u2_uk_n1114 ) , .B2( u2_uk_n1538 ) );
  NAND2_X1 u2_uk_U265 (.A1( u2_uk_K_r6_0 ) , .ZN( u2_uk_n1114 ) , .A2( u2_uk_n31 ) );
  OAI22_X1 u2_uk_U266 (.ZN( u2_K8_48 ) , .A2( u2_uk_n1504 ) , .B2( u2_uk_n1511 ) , .B1( u2_uk_n217 ) , .A1( u2_uk_n92 ) );
  OAI21_X1 u2_uk_U374 (.ZN( u2_K5_33 ) , .A( u2_uk_n1048 ) , .B2( u2_uk_n1401 ) , .B1( u2_uk_n202 ) );
  NAND2_X1 u2_uk_U375 (.A1( u2_uk_K_r3_14 ) , .ZN( u2_uk_n1048 ) , .A2( u2_uk_n203 ) );
  OAI22_X1 u2_uk_U470 (.ZN( u2_K5_37 ) , .B2( u2_uk_n1365 ) , .A2( u2_uk_n1403 ) , .B1( u2_uk_n147 ) , .A1( u2_uk_n92 ) );
  INV_X1 u2_uk_U561 (.ZN( u2_K5_36 ) , .A( u2_uk_n1050 ) );
  AOI22_X1 u2_uk_U562 (.B2( u2_uk_K_r3_29 ) , .A2( u2_uk_K_r3_52 ) , .ZN( u2_uk_n1050 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n191 ) );
  OAI22_X1 u2_uk_U764 (.ZN( u2_K2_21 ) , .A2( u2_uk_n1234 ) , .B2( u2_uk_n1238 ) , .B1( u2_uk_n142 ) , .A1( u2_uk_n94 ) );
  OAI22_X1 u2_uk_U79 (.ZN( u2_K2_23 ) , .B2( u2_uk_n1248 ) , .A2( u2_uk_n1269 ) , .B1( u2_uk_n222 ) , .A1( u2_uk_n94 ) );
  OAI22_X1 u2_uk_U884 (.ZN( u2_K2_24 ) , .A2( u2_uk_n1234 ) , .B2( u2_uk_n1249 ) , .A1( u2_uk_n161 ) , .B1( u2_uk_n63 ) );
  OAI22_X1 u2_uk_U949 (.ZN( u2_K5_40 ) , .B2( u2_uk_n1383 ) , .A2( u2_uk_n1400 ) , .B1( u2_uk_n146 ) , .A1( u2_uk_n92 ) );
  OAI22_X1 u2_uk_U950 (.ZN( u2_K2_22 ) , .B2( u2_uk_n1243 ) , .A2( u2_uk_n1260 ) , .B1( u2_uk_n230 ) , .A1( u2_uk_n94 ) );
endmodule

