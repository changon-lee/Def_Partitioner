module des_des_die_7 ( u0_K1_13, u0_K1_14, u0_K1_15, u0_K1_16, u0_K1_17, u0_K5_1, u0_K5_3, u0_K5_4, u0_K5_44, 
       u0_K5_47, u0_K5_48, u0_K8_28, u0_K8_33, u0_K8_36, u0_K9_14, u0_K9_15, u0_K9_32, u0_K9_39, 
       u0_K9_4, u0_K9_40, u0_K9_6, u0_L3_15, u0_L3_17, u0_L3_21, u0_L3_23, u0_L3_27, u0_L3_31, 
       u0_L3_5, u0_L3_9, u0_L6_11, u0_L6_12, u0_L6_14, u0_L6_19, u0_L6_22, u0_L6_25, u0_L6_29, 
       u0_L6_3, u0_L6_32, u0_L6_4, u0_L6_7, u0_L6_8, u0_L7_11, u0_L7_12, u0_L7_13, u0_L7_16, 
       u0_L7_17, u0_L7_18, u0_L7_19, u0_L7_2, u0_L7_22, u0_L7_23, u0_L7_24, u0_L7_28, u0_L7_29, 
       u0_L7_30, u0_L7_31, u0_L7_32, u0_L7_4, u0_L7_6, u0_L7_7, u0_L7_9, u0_R3_1, u0_R3_2, 
       u0_R3_28, u0_R3_29, u0_R3_3, u0_R3_30, u0_R3_31, u0_R3_32, u0_R3_4, u0_R3_5, u0_R6_16, 
       u0_R6_17, u0_R6_18, u0_R6_19, u0_R6_20, u0_R6_21, u0_R6_22, u0_R6_23, u0_R6_24, u0_R6_25, 
       u0_R6_26, u0_R6_27, u0_R6_28, u0_R6_29, u0_R7_1, u0_R7_10, u0_R7_11, u0_R7_12, u0_R7_13, 
       u0_R7_2, u0_R7_20, u0_R7_21, u0_R7_22, u0_R7_23, u0_R7_24, u0_R7_25, u0_R7_26, u0_R7_27, 
       u0_R7_28, u0_R7_29, u0_R7_3, u0_R7_32, u0_R7_4, u0_R7_5, u0_R7_6, u0_R7_7, u0_R7_8, 
       u0_R7_9, u0_desIn_r_13, u0_desIn_r_21, u0_desIn_r_29, u0_desIn_r_37, u0_desIn_r_40, u0_desIn_r_46, u0_desIn_r_5, u0_desIn_r_58, 
       u0_desIn_r_60, u0_desIn_r_63, u0_key_r_10, u0_key_r_45, u0_key_r_5, u0_key_r_55, u0_uk_K_r10_19, u0_uk_K_r12_18, u0_uk_K_r14_3, 
       u0_uk_K_r14_5, u0_uk_K_r3_10, u0_uk_K_r3_15, u0_uk_K_r3_38, u0_uk_K_r6_14, u0_uk_K_r6_21, u0_uk_K_r6_22, u0_uk_K_r6_29, u0_uk_K_r6_31, 
       u0_uk_K_r6_51, u0_uk_K_r6_55, u0_uk_K_r6_7, u0_uk_K_r7_1, u0_uk_K_r7_13, u0_uk_K_r7_15, u0_uk_K_r7_20, u0_uk_K_r7_22, u0_uk_K_r7_23, 
       u0_uk_K_r7_24, u0_uk_K_r7_25, u0_uk_K_r7_26, u0_uk_K_r7_27, u0_uk_K_r7_30, u0_uk_K_r7_32, u0_uk_K_r7_48, u0_uk_K_r7_55, u0_uk_K_r7_6, 
       u0_uk_K_r7_8, u0_uk_n100, u0_uk_n102, u0_uk_n109, u0_uk_n11, u0_uk_n110, u0_uk_n117, u0_uk_n128, u0_uk_n129, 
       u0_uk_n142, u0_uk_n145, u0_uk_n147, u0_uk_n148, u0_uk_n155, u0_uk_n161, u0_uk_n162, u0_uk_n17, u0_uk_n182, 
       u0_uk_n191, u0_uk_n202, u0_uk_n207, u0_uk_n208, u0_uk_n213, u0_uk_n214, u0_uk_n220, u0_uk_n222, u0_uk_n223, 
       u0_uk_n230, u0_uk_n231, u0_uk_n238, u0_uk_n240, u0_uk_n242, u0_uk_n250, u0_uk_n251, u0_uk_n257, u0_uk_n272, 
       u0_uk_n275, u0_uk_n276, u0_uk_n278, u0_uk_n283, u0_uk_n285, u0_uk_n289, u0_uk_n290, u0_uk_n300, u0_uk_n303, 
       u0_uk_n307, u0_uk_n309, u0_uk_n31, u0_uk_n310, u0_uk_n311, u0_uk_n314, u0_uk_n315, u0_uk_n316, u0_uk_n320, 
       u0_uk_n321, u0_uk_n322, u0_uk_n325, u0_uk_n327, u0_uk_n328, u0_uk_n332, u0_uk_n333, u0_uk_n341, u0_uk_n347, 
       u0_uk_n348, u0_uk_n354, u0_uk_n355, u0_uk_n359, u0_uk_n457, u0_uk_n466, u0_uk_n471, u0_uk_n486, u0_uk_n488, 
       u0_uk_n490, u0_uk_n491, u0_uk_n494, u0_uk_n60, u0_uk_n63, u0_uk_n725, u0_uk_n726, u0_uk_n736, u0_uk_n739, 
       u0_uk_n740, u0_uk_n748, u0_uk_n755, u0_uk_n805, u0_uk_n93, u0_uk_n99, u2_K10_25, u2_K10_26, u2_K10_30, 
       u2_K10_4, u2_K10_43, u2_K10_44, u2_K10_46, u2_K10_6, u2_K14_21, u2_K5_44, u2_K5_47, u2_K5_48, 
       u2_L12_1, u2_L12_10, u2_L12_20, u2_L12_26, u2_L3_15, u2_L3_21, u2_L3_27, u2_L3_5, u2_L8_14, 
       u2_L8_15, u2_L8_17, u2_L8_21, u2_L8_23, u2_L8_25, u2_L8_27, u2_L8_3, u2_L8_31, u2_L8_5, 
       u2_L8_8, u2_L8_9, u2_R12_12, u2_R12_13, u2_R12_14, u2_R12_15, u2_R12_16, u2_R12_17, u2_R3_1, 
       u2_R3_28, u2_R3_29, u2_R3_30, u2_R3_31, u2_R3_32, u2_R8_1, u2_R8_16, u2_R8_17, u2_R8_18, 
       u2_R8_19, u2_R8_2, u2_R8_20, u2_R8_21, u2_R8_28, u2_R8_29, u2_R8_3, u2_R8_30, u2_R8_31, 
       u2_R8_32, u2_R8_4, u2_R8_5, u2_uk_K_r12_25, u2_uk_K_r12_33, u2_uk_K_r12_41, u2_uk_K_r3_15, u2_uk_K_r3_38, u2_uk_K_r3_43, 
       u2_uk_K_r8_41, u2_uk_K_r8_43, u2_uk_n100, u2_uk_n102, u2_uk_n109, u2_uk_n117, u2_uk_n128, u2_uk_n1364, u2_uk_n1370, 
       u2_uk_n1401, u2_uk_n141, u2_uk_n146, u2_uk_n148, u2_uk_n155, u2_uk_n1592, u2_uk_n1594, u2_uk_n1595, u2_uk_n1597, 
       u2_uk_n1598, u2_uk_n1600, u2_uk_n1602, u2_uk_n1603, u2_uk_n1609, u2_uk_n1610, u2_uk_n1612, u2_uk_n1614, u2_uk_n1617, 
       u2_uk_n162, u2_uk_n1623, u2_uk_n1625, u2_uk_n1626, u2_uk_n163, u2_uk_n164, u2_uk_n17, u2_uk_n1772, u2_uk_n1779, 
       u2_uk_n1782, u2_uk_n1783, u2_uk_n1789, u2_uk_n1810, u2_uk_n182, u2_uk_n202, u2_uk_n207, u2_uk_n220, u2_uk_n223, 
       u2_uk_n230, u2_uk_n231, u2_uk_n251, u2_uk_n27, u2_uk_n63, u2_uk_n83, u2_uk_n92, u2_uk_n93, u2_uk_n94, 
       u2_uk_n99, u0_N132, u0_N136, u0_N142, u0_N144, u0_N148, u0_N15, u0_N150, u0_N154, u0_N158, 
        u0_N226, u0_N227, u0_N23, u0_N230, u0_N231, u0_N234, u0_N235, u0_N237, u0_N242, 
        u0_N245, u0_N248, u0_N252, u0_N255, u0_N257, u0_N259, u0_N261, u0_N262, u0_N264, 
        u0_N266, u0_N267, u0_N268, u0_N271, u0_N272, u0_N273, u0_N274, u0_N277, u0_N278, 
        u0_N279, u0_N283, u0_N284, u0_N285, u0_N286, u0_N287, u0_N29, u0_N5, u0_uk_n10, 
        u0_uk_n141, u0_uk_n27, u0_uk_n756, u0_uk_n762, u0_uk_n880, u0_uk_n888, u0_uk_n894, u0_uk_n906, u0_uk_n926, 
        u0_uk_n961, u2_N132, u2_N142, u2_N148, u2_N154, u2_N290, u2_N292, u2_N295, u2_N296, 
        u2_N301, u2_N302, u2_N304, u2_N308, u2_N310, u2_N312, u2_N314, u2_N318, u2_N416, 
        u2_N425, u2_N435, u2_N441 );
  input u0_K1_13, u0_K1_14, u0_K1_15, u0_K1_16, u0_K1_17, u0_K5_1, u0_K5_3, u0_K5_4, u0_K5_44, 
        u0_K5_47, u0_K5_48, u0_K8_28, u0_K8_33, u0_K8_36, u0_K9_14, u0_K9_15, u0_K9_32, u0_K9_39, 
        u0_K9_4, u0_K9_40, u0_K9_6, u0_L3_15, u0_L3_17, u0_L3_21, u0_L3_23, u0_L3_27, u0_L3_31, 
        u0_L3_5, u0_L3_9, u0_L6_11, u0_L6_12, u0_L6_14, u0_L6_19, u0_L6_22, u0_L6_25, u0_L6_29, 
        u0_L6_3, u0_L6_32, u0_L6_4, u0_L6_7, u0_L6_8, u0_L7_11, u0_L7_12, u0_L7_13, u0_L7_16, 
        u0_L7_17, u0_L7_18, u0_L7_19, u0_L7_2, u0_L7_22, u0_L7_23, u0_L7_24, u0_L7_28, u0_L7_29, 
        u0_L7_30, u0_L7_31, u0_L7_32, u0_L7_4, u0_L7_6, u0_L7_7, u0_L7_9, u0_R3_1, u0_R3_2, 
        u0_R3_28, u0_R3_29, u0_R3_3, u0_R3_30, u0_R3_31, u0_R3_32, u0_R3_4, u0_R3_5, u0_R6_16, 
        u0_R6_17, u0_R6_18, u0_R6_19, u0_R6_20, u0_R6_21, u0_R6_22, u0_R6_23, u0_R6_24, u0_R6_25, 
        u0_R6_26, u0_R6_27, u0_R6_28, u0_R6_29, u0_R7_1, u0_R7_10, u0_R7_11, u0_R7_12, u0_R7_13, 
        u0_R7_2, u0_R7_20, u0_R7_21, u0_R7_22, u0_R7_23, u0_R7_24, u0_R7_25, u0_R7_26, u0_R7_27, 
        u0_R7_28, u0_R7_29, u0_R7_3, u0_R7_32, u0_R7_4, u0_R7_5, u0_R7_6, u0_R7_7, u0_R7_8, 
        u0_R7_9, u0_desIn_r_13, u0_desIn_r_21, u0_desIn_r_29, u0_desIn_r_37, u0_desIn_r_40, u0_desIn_r_46, u0_desIn_r_5, u0_desIn_r_58, 
        u0_desIn_r_60, u0_desIn_r_63, u0_key_r_10, u0_key_r_45, u0_key_r_5, u0_key_r_55, u0_uk_K_r10_19, u0_uk_K_r12_18, u0_uk_K_r14_3, 
        u0_uk_K_r14_5, u0_uk_K_r3_10, u0_uk_K_r3_15, u0_uk_K_r3_38, u0_uk_K_r6_14, u0_uk_K_r6_21, u0_uk_K_r6_22, u0_uk_K_r6_29, u0_uk_K_r6_31, 
        u0_uk_K_r6_51, u0_uk_K_r6_55, u0_uk_K_r6_7, u0_uk_K_r7_1, u0_uk_K_r7_13, u0_uk_K_r7_15, u0_uk_K_r7_20, u0_uk_K_r7_22, u0_uk_K_r7_23, 
        u0_uk_K_r7_24, u0_uk_K_r7_25, u0_uk_K_r7_26, u0_uk_K_r7_27, u0_uk_K_r7_30, u0_uk_K_r7_32, u0_uk_K_r7_48, u0_uk_K_r7_55, u0_uk_K_r7_6, 
        u0_uk_K_r7_8, u0_uk_n100, u0_uk_n102, u0_uk_n109, u0_uk_n11, u0_uk_n110, u0_uk_n117, u0_uk_n128, u0_uk_n129, 
        u0_uk_n142, u0_uk_n145, u0_uk_n147, u0_uk_n148, u0_uk_n155, u0_uk_n161, u0_uk_n162, u0_uk_n17, u0_uk_n182, 
        u0_uk_n191, u0_uk_n202, u0_uk_n207, u0_uk_n208, u0_uk_n213, u0_uk_n214, u0_uk_n220, u0_uk_n222, u0_uk_n223, 
        u0_uk_n230, u0_uk_n231, u0_uk_n238, u0_uk_n240, u0_uk_n242, u0_uk_n250, u0_uk_n251, u0_uk_n257, u0_uk_n272, 
        u0_uk_n275, u0_uk_n276, u0_uk_n278, u0_uk_n283, u0_uk_n285, u0_uk_n289, u0_uk_n290, u0_uk_n300, u0_uk_n303, 
        u0_uk_n307, u0_uk_n309, u0_uk_n31, u0_uk_n310, u0_uk_n311, u0_uk_n314, u0_uk_n315, u0_uk_n316, u0_uk_n320, 
        u0_uk_n321, u0_uk_n322, u0_uk_n325, u0_uk_n327, u0_uk_n328, u0_uk_n332, u0_uk_n333, u0_uk_n341, u0_uk_n347, 
        u0_uk_n348, u0_uk_n354, u0_uk_n355, u0_uk_n359, u0_uk_n457, u0_uk_n466, u0_uk_n471, u0_uk_n486, u0_uk_n488, 
        u0_uk_n490, u0_uk_n491, u0_uk_n494, u0_uk_n60, u0_uk_n63, u0_uk_n725, u0_uk_n726, u0_uk_n736, u0_uk_n739, 
        u0_uk_n740, u0_uk_n748, u0_uk_n755, u0_uk_n805, u0_uk_n93, u0_uk_n99, u2_K10_25, u2_K10_26, u2_K10_30, 
        u2_K10_4, u2_K10_43, u2_K10_44, u2_K10_46, u2_K10_6, u2_K14_21, u2_K5_44, u2_K5_47, u2_K5_48, 
        u2_L12_1, u2_L12_10, u2_L12_20, u2_L12_26, u2_L3_15, u2_L3_21, u2_L3_27, u2_L3_5, u2_L8_14, 
        u2_L8_15, u2_L8_17, u2_L8_21, u2_L8_23, u2_L8_25, u2_L8_27, u2_L8_3, u2_L8_31, u2_L8_5, 
        u2_L8_8, u2_L8_9, u2_R12_12, u2_R12_13, u2_R12_14, u2_R12_15, u2_R12_16, u2_R12_17, u2_R3_1, 
        u2_R3_28, u2_R3_29, u2_R3_30, u2_R3_31, u2_R3_32, u2_R8_1, u2_R8_16, u2_R8_17, u2_R8_18, 
        u2_R8_19, u2_R8_2, u2_R8_20, u2_R8_21, u2_R8_28, u2_R8_29, u2_R8_3, u2_R8_30, u2_R8_31, 
        u2_R8_32, u2_R8_4, u2_R8_5, u2_uk_K_r12_25, u2_uk_K_r12_33, u2_uk_K_r12_41, u2_uk_K_r3_15, u2_uk_K_r3_38, u2_uk_K_r3_43, 
        u2_uk_K_r8_41, u2_uk_K_r8_43, u2_uk_n100, u2_uk_n102, u2_uk_n109, u2_uk_n117, u2_uk_n128, u2_uk_n1364, u2_uk_n1370, 
        u2_uk_n1401, u2_uk_n141, u2_uk_n146, u2_uk_n148, u2_uk_n155, u2_uk_n1592, u2_uk_n1594, u2_uk_n1595, u2_uk_n1597, 
        u2_uk_n1598, u2_uk_n1600, u2_uk_n1602, u2_uk_n1603, u2_uk_n1609, u2_uk_n1610, u2_uk_n1612, u2_uk_n1614, u2_uk_n1617, 
        u2_uk_n162, u2_uk_n1623, u2_uk_n1625, u2_uk_n1626, u2_uk_n163, u2_uk_n164, u2_uk_n17, u2_uk_n1772, u2_uk_n1779, 
        u2_uk_n1782, u2_uk_n1783, u2_uk_n1789, u2_uk_n1810, u2_uk_n182, u2_uk_n202, u2_uk_n207, u2_uk_n220, u2_uk_n223, 
        u2_uk_n230, u2_uk_n231, u2_uk_n251, u2_uk_n27, u2_uk_n63, u2_uk_n83, u2_uk_n92, u2_uk_n93, u2_uk_n94, 
        u2_uk_n99;
  output u0_N132, u0_N136, u0_N142, u0_N144, u0_N148, u0_N15, u0_N150, u0_N154, u0_N158, 
        u0_N226, u0_N227, u0_N23, u0_N230, u0_N231, u0_N234, u0_N235, u0_N237, u0_N242, 
        u0_N245, u0_N248, u0_N252, u0_N255, u0_N257, u0_N259, u0_N261, u0_N262, u0_N264, 
        u0_N266, u0_N267, u0_N268, u0_N271, u0_N272, u0_N273, u0_N274, u0_N277, u0_N278, 
        u0_N279, u0_N283, u0_N284, u0_N285, u0_N286, u0_N287, u0_N29, u0_N5, u0_uk_n10, 
        u0_uk_n141, u0_uk_n27, u0_uk_n756, u0_uk_n762, u0_uk_n880, u0_uk_n888, u0_uk_n894, u0_uk_n906, u0_uk_n926, 
        u0_uk_n961, u2_N132, u2_N142, u2_N148, u2_N154, u2_N290, u2_N292, u2_N295, u2_N296, 
        u2_N301, u2_N302, u2_N304, u2_N308, u2_N310, u2_N312, u2_N314, u2_N318, u2_N416, 
        u2_N425, u2_N435, u2_N441;
  wire u0_K1_18, u0_K5_2, u0_K5_43, u0_K5_45, u0_K5_46, u0_K5_5, u0_K5_6, u0_K8_25, u0_K8_26, 
       u0_K8_27, u0_K8_29, u0_K8_30, u0_K8_31, u0_K8_32, u0_K8_34, u0_K8_35, u0_K8_37, u0_K8_38, 
       u0_K8_39, u0_K8_40, u0_K8_41, u0_K8_42, u0_K9_1, u0_K9_10, u0_K9_11, u0_K9_12, u0_K9_13, 
       u0_K9_16, u0_K9_17, u0_K9_18, u0_K9_2, u0_K9_3, u0_K9_31, u0_K9_33, u0_K9_34, u0_K9_35, 
       u0_K9_36, u0_K9_37, u0_K9_38, u0_K9_41, u0_K9_42, u0_K9_5, u0_K9_7, u0_K9_8, u0_K9_9, 
       u0_out0_16, u0_out0_24, u0_out0_30, u0_out0_6, u0_out4_15, u0_out4_17, u0_out4_21, u0_out4_23, u0_out4_27, 
       u0_out4_31, u0_out4_5, u0_out4_9, u0_out7_11, u0_out7_12, u0_out7_14, u0_out7_19, u0_out7_22, u0_out7_25, 
       u0_out7_29, u0_out7_3, u0_out7_32, u0_out7_4, u0_out7_7, u0_out7_8, u0_out8_11, u0_out8_12, u0_out8_13, 
       u0_out8_16, u0_out8_17, u0_out8_18, u0_out8_19, u0_out8_2, u0_out8_22, u0_out8_23, u0_out8_24, u0_out8_28, 
       u0_out8_29, u0_out8_30, u0_out8_31, u0_out8_32, u0_out8_4, u0_out8_6, u0_out8_7, u0_out8_9, u0_u0_X_13, 
       u0_u0_X_14, u0_u0_X_15, u0_u0_X_16, u0_u0_X_17, u0_u0_X_18, u0_u0_u2_n1, u0_u0_u2_n10, u0_u0_u2_n11, u0_u0_u2_n12, 
       u0_u0_u2_n13, u0_u0_u2_n14, u0_u0_u2_n15, u0_u0_u2_n16, u0_u0_u2_n17, u0_u0_u2_n18, u0_u0_u2_n19, u0_u0_u2_n2, u0_u0_u2_n20, 
       u0_u0_u2_n21, u0_u0_u2_n22, u0_u0_u2_n23, u0_u0_u2_n24, u0_u0_u2_n25, u0_u0_u2_n26, u0_u0_u2_n27, u0_u0_u2_n28, u0_u0_u2_n29, 
       u0_u0_u2_n3, u0_u0_u2_n30, u0_u0_u2_n31, u0_u0_u2_n32, u0_u0_u2_n33, u0_u0_u2_n34, u0_u0_u2_n35, u0_u0_u2_n36, u0_u0_u2_n37, 
       u0_u0_u2_n38, u0_u0_u2_n39, u0_u0_u2_n4, u0_u0_u2_n40, u0_u0_u2_n41, u0_u0_u2_n42, u0_u0_u2_n43, u0_u0_u2_n44, u0_u0_u2_n45, 
       u0_u0_u2_n46, u0_u0_u2_n47, u0_u0_u2_n48, u0_u0_u2_n49, u0_u0_u2_n5, u0_u0_u2_n50, u0_u0_u2_n51, u0_u0_u2_n52, u0_u0_u2_n53, 
       u0_u0_u2_n54, u0_u0_u2_n55, u0_u0_u2_n56, u0_u0_u2_n57, u0_u0_u2_n58, u0_u0_u2_n59, u0_u0_u2_n6, u0_u0_u2_n60, u0_u0_u2_n61, 
       u0_u0_u2_n62, u0_u0_u2_n63, u0_u0_u2_n64, u0_u0_u2_n65, u0_u0_u2_n66, u0_u0_u2_n67, u0_u0_u2_n68, u0_u0_u2_n69, u0_u0_u2_n7, 
       u0_u0_u2_n70, u0_u0_u2_n71, u0_u0_u2_n72, u0_u0_u2_n73, u0_u0_u2_n74, u0_u0_u2_n75, u0_u0_u2_n76, u0_u0_u2_n77, u0_u0_u2_n78, 
       u0_u0_u2_n79, u0_u0_u2_n8, u0_u0_u2_n80, u0_u0_u2_n81, u0_u0_u2_n82, u0_u0_u2_n83, u0_u0_u2_n84, u0_u0_u2_n85, u0_u0_u2_n86, 
       u0_u0_u2_n87, u0_u0_u2_n88, u0_u0_u2_n89, u0_u0_u2_n9, u0_u0_u2_n90, u0_u0_u2_n91, u0_u0_u2_n92, u0_u0_u2_n93, u0_u0_u2_n94, 
       u0_u4_X_1, u0_u4_X_2, u0_u4_X_3, u0_u4_X_4, u0_u4_X_43, u0_u4_X_44, u0_u4_X_45, u0_u4_X_46, u0_u4_X_47, 
       u0_u4_X_48, u0_u4_X_5, u0_u4_X_6, u0_u4_u0_n100, u0_u4_u0_n101, u0_u4_u0_n102, u0_u4_u0_n103, u0_u4_u0_n104, u0_u4_u0_n105, 
       u0_u4_u0_n106, u0_u4_u0_n107, u0_u4_u0_n108, u0_u4_u0_n109, u0_u4_u0_n110, u0_u4_u0_n111, u0_u4_u0_n112, u0_u4_u0_n113, u0_u4_u0_n114, 
       u0_u4_u0_n115, u0_u4_u0_n116, u0_u4_u0_n117, u0_u4_u0_n118, u0_u4_u0_n119, u0_u4_u0_n120, u0_u4_u0_n121, u0_u4_u0_n122, u0_u4_u0_n123, 
       u0_u4_u0_n124, u0_u4_u0_n125, u0_u4_u0_n126, u0_u4_u0_n127, u0_u4_u0_n128, u0_u4_u0_n129, u0_u4_u0_n130, u0_u4_u0_n131, u0_u4_u0_n132, 
       u0_u4_u0_n133, u0_u4_u0_n134, u0_u4_u0_n135, u0_u4_u0_n136, u0_u4_u0_n137, u0_u4_u0_n138, u0_u4_u0_n139, u0_u4_u0_n140, u0_u4_u0_n141, 
       u0_u4_u0_n142, u0_u4_u0_n143, u0_u4_u0_n144, u0_u4_u0_n145, u0_u4_u0_n146, u0_u4_u0_n147, u0_u4_u0_n148, u0_u4_u0_n149, u0_u4_u0_n150, 
       u0_u4_u0_n151, u0_u4_u0_n152, u0_u4_u0_n153, u0_u4_u0_n154, u0_u4_u0_n155, u0_u4_u0_n156, u0_u4_u0_n157, u0_u4_u0_n158, u0_u4_u0_n159, 
       u0_u4_u0_n160, u0_u4_u0_n161, u0_u4_u0_n162, u0_u4_u0_n163, u0_u4_u0_n164, u0_u4_u0_n165, u0_u4_u0_n166, u0_u4_u0_n167, u0_u4_u0_n168, 
       u0_u4_u0_n169, u0_u4_u0_n170, u0_u4_u0_n171, u0_u4_u0_n172, u0_u4_u0_n173, u0_u4_u0_n174, u0_u4_u0_n88, u0_u4_u0_n89, u0_u4_u0_n90, 
       u0_u4_u0_n91, u0_u4_u0_n92, u0_u4_u0_n93, u0_u4_u0_n94, u0_u4_u0_n95, u0_u4_u0_n96, u0_u4_u0_n97, u0_u4_u0_n98, u0_u4_u0_n99, 
       u0_u4_u7_n100, u0_u4_u7_n101, u0_u4_u7_n102, u0_u4_u7_n103, u0_u4_u7_n104, u0_u4_u7_n105, u0_u4_u7_n106, u0_u4_u7_n107, u0_u4_u7_n108, 
       u0_u4_u7_n109, u0_u4_u7_n110, u0_u4_u7_n111, u0_u4_u7_n112, u0_u4_u7_n113, u0_u4_u7_n114, u0_u4_u7_n115, u0_u4_u7_n116, u0_u4_u7_n117, 
       u0_u4_u7_n118, u0_u4_u7_n119, u0_u4_u7_n120, u0_u4_u7_n121, u0_u4_u7_n122, u0_u4_u7_n123, u0_u4_u7_n124, u0_u4_u7_n125, u0_u4_u7_n126, 
       u0_u4_u7_n127, u0_u4_u7_n128, u0_u4_u7_n129, u0_u4_u7_n130, u0_u4_u7_n131, u0_u4_u7_n132, u0_u4_u7_n133, u0_u4_u7_n134, u0_u4_u7_n135, 
       u0_u4_u7_n136, u0_u4_u7_n137, u0_u4_u7_n138, u0_u4_u7_n139, u0_u4_u7_n140, u0_u4_u7_n141, u0_u4_u7_n142, u0_u4_u7_n143, u0_u4_u7_n144, 
       u0_u4_u7_n145, u0_u4_u7_n146, u0_u4_u7_n147, u0_u4_u7_n148, u0_u4_u7_n149, u0_u4_u7_n150, u0_u4_u7_n151, u0_u4_u7_n152, u0_u4_u7_n153, 
       u0_u4_u7_n154, u0_u4_u7_n155, u0_u4_u7_n156, u0_u4_u7_n157, u0_u4_u7_n158, u0_u4_u7_n159, u0_u4_u7_n160, u0_u4_u7_n161, u0_u4_u7_n162, 
       u0_u4_u7_n163, u0_u4_u7_n164, u0_u4_u7_n165, u0_u4_u7_n166, u0_u4_u7_n167, u0_u4_u7_n168, u0_u4_u7_n169, u0_u4_u7_n170, u0_u4_u7_n171, 
       u0_u4_u7_n172, u0_u4_u7_n173, u0_u4_u7_n174, u0_u4_u7_n175, u0_u4_u7_n176, u0_u4_u7_n177, u0_u4_u7_n178, u0_u4_u7_n179, u0_u4_u7_n180, 
       u0_u4_u7_n91, u0_u4_u7_n92, u0_u4_u7_n93, u0_u4_u7_n94, u0_u4_u7_n95, u0_u4_u7_n96, u0_u4_u7_n97, u0_u4_u7_n98, u0_u4_u7_n99, 
       u0_u7_X_25, u0_u7_X_26, u0_u7_X_27, u0_u7_X_28, u0_u7_X_29, u0_u7_X_30, u0_u7_X_31, u0_u7_X_32, u0_u7_X_33, 
       u0_u7_X_34, u0_u7_X_35, u0_u7_X_36, u0_u7_X_37, u0_u7_X_38, u0_u7_X_39, u0_u7_X_40, u0_u7_X_41, u0_u7_X_42, 
       u0_u7_u4_n100, u0_u7_u4_n101, u0_u7_u4_n102, u0_u7_u4_n103, u0_u7_u4_n104, u0_u7_u4_n105, u0_u7_u4_n106, u0_u7_u4_n107, u0_u7_u4_n108, 
       u0_u7_u4_n109, u0_u7_u4_n110, u0_u7_u4_n111, u0_u7_u4_n112, u0_u7_u4_n113, u0_u7_u4_n114, u0_u7_u4_n115, u0_u7_u4_n116, u0_u7_u4_n117, 
       u0_u7_u4_n118, u0_u7_u4_n119, u0_u7_u4_n120, u0_u7_u4_n121, u0_u7_u4_n122, u0_u7_u4_n123, u0_u7_u4_n124, u0_u7_u4_n125, u0_u7_u4_n126, 
       u0_u7_u4_n127, u0_u7_u4_n128, u0_u7_u4_n129, u0_u7_u4_n130, u0_u7_u4_n131, u0_u7_u4_n132, u0_u7_u4_n133, u0_u7_u4_n134, u0_u7_u4_n135, 
       u0_u7_u4_n136, u0_u7_u4_n137, u0_u7_u4_n138, u0_u7_u4_n139, u0_u7_u4_n140, u0_u7_u4_n141, u0_u7_u4_n142, u0_u7_u4_n143, u0_u7_u4_n144, 
       u0_u7_u4_n145, u0_u7_u4_n146, u0_u7_u4_n147, u0_u7_u4_n148, u0_u7_u4_n149, u0_u7_u4_n150, u0_u7_u4_n151, u0_u7_u4_n152, u0_u7_u4_n153, 
       u0_u7_u4_n154, u0_u7_u4_n155, u0_u7_u4_n156, u0_u7_u4_n157, u0_u7_u4_n158, u0_u7_u4_n159, u0_u7_u4_n160, u0_u7_u4_n161, u0_u7_u4_n162, 
       u0_u7_u4_n163, u0_u7_u4_n164, u0_u7_u4_n165, u0_u7_u4_n166, u0_u7_u4_n167, u0_u7_u4_n168, u0_u7_u4_n169, u0_u7_u4_n170, u0_u7_u4_n171, 
       u0_u7_u4_n172, u0_u7_u4_n173, u0_u7_u4_n174, u0_u7_u4_n175, u0_u7_u4_n176, u0_u7_u4_n177, u0_u7_u4_n178, u0_u7_u4_n179, u0_u7_u4_n180, 
       u0_u7_u4_n181, u0_u7_u4_n182, u0_u7_u4_n183, u0_u7_u4_n184, u0_u7_u4_n185, u0_u7_u4_n186, u0_u7_u4_n94, u0_u7_u4_n95, u0_u7_u4_n96, 
       u0_u7_u4_n97, u0_u7_u4_n98, u0_u7_u4_n99, u0_u7_u5_n100, u0_u7_u5_n101, u0_u7_u5_n102, u0_u7_u5_n103, u0_u7_u5_n104, u0_u7_u5_n105, 
       u0_u7_u5_n106, u0_u7_u5_n107, u0_u7_u5_n108, u0_u7_u5_n109, u0_u7_u5_n110, u0_u7_u5_n111, u0_u7_u5_n112, u0_u7_u5_n113, u0_u7_u5_n114, 
       u0_u7_u5_n115, u0_u7_u5_n116, u0_u7_u5_n117, u0_u7_u5_n118, u0_u7_u5_n119, u0_u7_u5_n120, u0_u7_u5_n121, u0_u7_u5_n122, u0_u7_u5_n123, 
       u0_u7_u5_n124, u0_u7_u5_n125, u0_u7_u5_n126, u0_u7_u5_n127, u0_u7_u5_n128, u0_u7_u5_n129, u0_u7_u5_n130, u0_u7_u5_n131, u0_u7_u5_n132, 
       u0_u7_u5_n133, u0_u7_u5_n134, u0_u7_u5_n135, u0_u7_u5_n136, u0_u7_u5_n137, u0_u7_u5_n138, u0_u7_u5_n139, u0_u7_u5_n140, u0_u7_u5_n141, 
       u0_u7_u5_n142, u0_u7_u5_n143, u0_u7_u5_n144, u0_u7_u5_n145, u0_u7_u5_n146, u0_u7_u5_n147, u0_u7_u5_n148, u0_u7_u5_n149, u0_u7_u5_n150, 
       u0_u7_u5_n151, u0_u7_u5_n152, u0_u7_u5_n153, u0_u7_u5_n154, u0_u7_u5_n155, u0_u7_u5_n156, u0_u7_u5_n157, u0_u7_u5_n158, u0_u7_u5_n159, 
       u0_u7_u5_n160, u0_u7_u5_n161, u0_u7_u5_n162, u0_u7_u5_n163, u0_u7_u5_n164, u0_u7_u5_n165, u0_u7_u5_n166, u0_u7_u5_n167, u0_u7_u5_n168, 
       u0_u7_u5_n169, u0_u7_u5_n170, u0_u7_u5_n171, u0_u7_u5_n172, u0_u7_u5_n173, u0_u7_u5_n174, u0_u7_u5_n175, u0_u7_u5_n176, u0_u7_u5_n177, 
       u0_u7_u5_n178, u0_u7_u5_n179, u0_u7_u5_n180, u0_u7_u5_n181, u0_u7_u5_n182, u0_u7_u5_n183, u0_u7_u5_n184, u0_u7_u5_n185, u0_u7_u5_n186, 
       u0_u7_u5_n187, u0_u7_u5_n188, u0_u7_u5_n189, u0_u7_u5_n190, u0_u7_u5_n191, u0_u7_u5_n192, u0_u7_u5_n193, u0_u7_u5_n194, u0_u7_u5_n195, 
       u0_u7_u5_n196, u0_u7_u5_n99, u0_u7_u6_n100, u0_u7_u6_n101, u0_u7_u6_n102, u0_u7_u6_n103, u0_u7_u6_n104, u0_u7_u6_n105, u0_u7_u6_n106, 
       u0_u7_u6_n107, u0_u7_u6_n108, u0_u7_u6_n109, u0_u7_u6_n110, u0_u7_u6_n111, u0_u7_u6_n112, u0_u7_u6_n113, u0_u7_u6_n114, u0_u7_u6_n115, 
       u0_u7_u6_n116, u0_u7_u6_n117, u0_u7_u6_n118, u0_u7_u6_n119, u0_u7_u6_n120, u0_u7_u6_n121, u0_u7_u6_n122, u0_u7_u6_n123, u0_u7_u6_n124, 
       u0_u7_u6_n125, u0_u7_u6_n126, u0_u7_u6_n127, u0_u7_u6_n128, u0_u7_u6_n129, u0_u7_u6_n130, u0_u7_u6_n131, u0_u7_u6_n132, u0_u7_u6_n133, 
       u0_u7_u6_n134, u0_u7_u6_n135, u0_u7_u6_n136, u0_u7_u6_n137, u0_u7_u6_n138, u0_u7_u6_n139, u0_u7_u6_n140, u0_u7_u6_n141, u0_u7_u6_n142, 
       u0_u7_u6_n143, u0_u7_u6_n144, u0_u7_u6_n145, u0_u7_u6_n146, u0_u7_u6_n147, u0_u7_u6_n148, u0_u7_u6_n149, u0_u7_u6_n150, u0_u7_u6_n151, 
       u0_u7_u6_n152, u0_u7_u6_n153, u0_u7_u6_n154, u0_u7_u6_n155, u0_u7_u6_n156, u0_u7_u6_n157, u0_u7_u6_n158, u0_u7_u6_n159, u0_u7_u6_n160, 
       u0_u7_u6_n161, u0_u7_u6_n162, u0_u7_u6_n163, u0_u7_u6_n164, u0_u7_u6_n165, u0_u7_u6_n166, u0_u7_u6_n167, u0_u7_u6_n168, u0_u7_u6_n169, 
       u0_u7_u6_n170, u0_u7_u6_n171, u0_u7_u6_n172, u0_u7_u6_n173, u0_u7_u6_n174, u0_u7_u6_n88, u0_u7_u6_n89, u0_u7_u6_n90, u0_u7_u6_n91, 
       u0_u7_u6_n92, u0_u7_u6_n93, u0_u7_u6_n94, u0_u7_u6_n95, u0_u7_u6_n96, u0_u7_u6_n97, u0_u7_u6_n98, u0_u7_u6_n99, u0_u8_X_1, 
       u0_u8_X_10, u0_u8_X_11, u0_u8_X_12, u0_u8_X_13, u0_u8_X_14, u0_u8_X_15, u0_u8_X_16, u0_u8_X_17, u0_u8_X_18, 
       u0_u8_X_2, u0_u8_X_3, u0_u8_X_31, u0_u8_X_32, u0_u8_X_33, u0_u8_X_34, u0_u8_X_35, u0_u8_X_36, u0_u8_X_37, 
       u0_u8_X_38, u0_u8_X_39, u0_u8_X_4, u0_u8_X_40, u0_u8_X_41, u0_u8_X_42, u0_u8_X_5, u0_u8_X_6, u0_u8_X_7, 
       u0_u8_X_8, u0_u8_X_9, u0_u8_u0_n100, u0_u8_u0_n101, u0_u8_u0_n102, u0_u8_u0_n103, u0_u8_u0_n104, u0_u8_u0_n105, u0_u8_u0_n106, 
       u0_u8_u0_n107, u0_u8_u0_n108, u0_u8_u0_n109, u0_u8_u0_n110, u0_u8_u0_n111, u0_u8_u0_n112, u0_u8_u0_n113, u0_u8_u0_n114, u0_u8_u0_n115, 
       u0_u8_u0_n116, u0_u8_u0_n117, u0_u8_u0_n118, u0_u8_u0_n119, u0_u8_u0_n120, u0_u8_u0_n121, u0_u8_u0_n122, u0_u8_u0_n123, u0_u8_u0_n124, 
       u0_u8_u0_n125, u0_u8_u0_n126, u0_u8_u0_n127, u0_u8_u0_n128, u0_u8_u0_n129, u0_u8_u0_n130, u0_u8_u0_n131, u0_u8_u0_n132, u0_u8_u0_n133, 
       u0_u8_u0_n134, u0_u8_u0_n135, u0_u8_u0_n136, u0_u8_u0_n137, u0_u8_u0_n138, u0_u8_u0_n139, u0_u8_u0_n140, u0_u8_u0_n141, u0_u8_u0_n142, 
       u0_u8_u0_n143, u0_u8_u0_n144, u0_u8_u0_n145, u0_u8_u0_n146, u0_u8_u0_n147, u0_u8_u0_n148, u0_u8_u0_n149, u0_u8_u0_n150, u0_u8_u0_n151, 
       u0_u8_u0_n152, u0_u8_u0_n153, u0_u8_u0_n154, u0_u8_u0_n155, u0_u8_u0_n156, u0_u8_u0_n157, u0_u8_u0_n158, u0_u8_u0_n159, u0_u8_u0_n160, 
       u0_u8_u0_n161, u0_u8_u0_n162, u0_u8_u0_n163, u0_u8_u0_n164, u0_u8_u0_n165, u0_u8_u0_n166, u0_u8_u0_n167, u0_u8_u0_n168, u0_u8_u0_n169, 
       u0_u8_u0_n170, u0_u8_u0_n171, u0_u8_u0_n172, u0_u8_u0_n173, u0_u8_u0_n174, u0_u8_u0_n88, u0_u8_u0_n89, u0_u8_u0_n90, u0_u8_u0_n91, 
       u0_u8_u0_n92, u0_u8_u0_n93, u0_u8_u0_n94, u0_u8_u0_n95, u0_u8_u0_n96, u0_u8_u0_n97, u0_u8_u0_n98, u0_u8_u0_n99, u0_u8_u1_n100, 
       u0_u8_u1_n101, u0_u8_u1_n102, u0_u8_u1_n103, u0_u8_u1_n104, u0_u8_u1_n105, u0_u8_u1_n106, u0_u8_u1_n107, u0_u8_u1_n108, u0_u8_u1_n109, 
       u0_u8_u1_n110, u0_u8_u1_n111, u0_u8_u1_n112, u0_u8_u1_n113, u0_u8_u1_n114, u0_u8_u1_n115, u0_u8_u1_n116, u0_u8_u1_n117, u0_u8_u1_n118, 
       u0_u8_u1_n119, u0_u8_u1_n120, u0_u8_u1_n121, u0_u8_u1_n122, u0_u8_u1_n123, u0_u8_u1_n124, u0_u8_u1_n125, u0_u8_u1_n126, u0_u8_u1_n127, 
       u0_u8_u1_n128, u0_u8_u1_n129, u0_u8_u1_n130, u0_u8_u1_n131, u0_u8_u1_n132, u0_u8_u1_n133, u0_u8_u1_n134, u0_u8_u1_n135, u0_u8_u1_n136, 
       u0_u8_u1_n137, u0_u8_u1_n138, u0_u8_u1_n139, u0_u8_u1_n140, u0_u8_u1_n141, u0_u8_u1_n142, u0_u8_u1_n143, u0_u8_u1_n144, u0_u8_u1_n145, 
       u0_u8_u1_n146, u0_u8_u1_n147, u0_u8_u1_n148, u0_u8_u1_n149, u0_u8_u1_n150, u0_u8_u1_n151, u0_u8_u1_n152, u0_u8_u1_n153, u0_u8_u1_n154, 
       u0_u8_u1_n155, u0_u8_u1_n156, u0_u8_u1_n157, u0_u8_u1_n158, u0_u8_u1_n159, u0_u8_u1_n160, u0_u8_u1_n161, u0_u8_u1_n162, u0_u8_u1_n163, 
       u0_u8_u1_n164, u0_u8_u1_n165, u0_u8_u1_n166, u0_u8_u1_n167, u0_u8_u1_n168, u0_u8_u1_n169, u0_u8_u1_n170, u0_u8_u1_n171, u0_u8_u1_n172, 
       u0_u8_u1_n173, u0_u8_u1_n174, u0_u8_u1_n175, u0_u8_u1_n176, u0_u8_u1_n177, u0_u8_u1_n178, u0_u8_u1_n179, u0_u8_u1_n180, u0_u8_u1_n181, 
       u0_u8_u1_n182, u0_u8_u1_n183, u0_u8_u1_n184, u0_u8_u1_n185, u0_u8_u1_n186, u0_u8_u1_n187, u0_u8_u1_n188, u0_u8_u1_n95, u0_u8_u1_n96, 
       u0_u8_u1_n97, u0_u8_u1_n98, u0_u8_u1_n99, u0_u8_u2_n100, u0_u8_u2_n101, u0_u8_u2_n102, u0_u8_u2_n103, u0_u8_u2_n104, u0_u8_u2_n105, 
       u0_u8_u2_n106, u0_u8_u2_n107, u0_u8_u2_n108, u0_u8_u2_n109, u0_u8_u2_n110, u0_u8_u2_n111, u0_u8_u2_n112, u0_u8_u2_n113, u0_u8_u2_n114, 
       u0_u8_u2_n115, u0_u8_u2_n116, u0_u8_u2_n117, u0_u8_u2_n118, u0_u8_u2_n119, u0_u8_u2_n120, u0_u8_u2_n121, u0_u8_u2_n122, u0_u8_u2_n123, 
       u0_u8_u2_n124, u0_u8_u2_n125, u0_u8_u2_n126, u0_u8_u2_n127, u0_u8_u2_n128, u0_u8_u2_n129, u0_u8_u2_n130, u0_u8_u2_n131, u0_u8_u2_n132, 
       u0_u8_u2_n133, u0_u8_u2_n134, u0_u8_u2_n135, u0_u8_u2_n136, u0_u8_u2_n137, u0_u8_u2_n138, u0_u8_u2_n139, u0_u8_u2_n140, u0_u8_u2_n141, 
       u0_u8_u2_n142, u0_u8_u2_n143, u0_u8_u2_n144, u0_u8_u2_n145, u0_u8_u2_n146, u0_u8_u2_n147, u0_u8_u2_n148, u0_u8_u2_n149, u0_u8_u2_n150, 
       u0_u8_u2_n151, u0_u8_u2_n152, u0_u8_u2_n153, u0_u8_u2_n154, u0_u8_u2_n155, u0_u8_u2_n156, u0_u8_u2_n157, u0_u8_u2_n158, u0_u8_u2_n159, 
       u0_u8_u2_n160, u0_u8_u2_n161, u0_u8_u2_n162, u0_u8_u2_n163, u0_u8_u2_n164, u0_u8_u2_n165, u0_u8_u2_n166, u0_u8_u2_n167, u0_u8_u2_n168, 
       u0_u8_u2_n169, u0_u8_u2_n170, u0_u8_u2_n171, u0_u8_u2_n172, u0_u8_u2_n173, u0_u8_u2_n174, u0_u8_u2_n175, u0_u8_u2_n176, u0_u8_u2_n177, 
       u0_u8_u2_n178, u0_u8_u2_n179, u0_u8_u2_n180, u0_u8_u2_n181, u0_u8_u2_n182, u0_u8_u2_n183, u0_u8_u2_n184, u0_u8_u2_n185, u0_u8_u2_n186, 
       u0_u8_u2_n187, u0_u8_u2_n188, u0_u8_u2_n95, u0_u8_u2_n96, u0_u8_u2_n97, u0_u8_u2_n98, u0_u8_u2_n99, u0_u8_u5_n100, u0_u8_u5_n101, 
       u0_u8_u5_n102, u0_u8_u5_n103, u0_u8_u5_n104, u0_u8_u5_n105, u0_u8_u5_n106, u0_u8_u5_n107, u0_u8_u5_n108, u0_u8_u5_n109, u0_u8_u5_n110, 
       u0_u8_u5_n111, u0_u8_u5_n112, u0_u8_u5_n113, u0_u8_u5_n114, u0_u8_u5_n115, u0_u8_u5_n116, u0_u8_u5_n117, u0_u8_u5_n118, u0_u8_u5_n119, 
       u0_u8_u5_n120, u0_u8_u5_n121, u0_u8_u5_n122, u0_u8_u5_n123, u0_u8_u5_n124, u0_u8_u5_n125, u0_u8_u5_n126, u0_u8_u5_n127, u0_u8_u5_n128, 
       u0_u8_u5_n129, u0_u8_u5_n130, u0_u8_u5_n131, u0_u8_u5_n132, u0_u8_u5_n133, u0_u8_u5_n134, u0_u8_u5_n135, u0_u8_u5_n136, u0_u8_u5_n137, 
       u0_u8_u5_n138, u0_u8_u5_n139, u0_u8_u5_n140, u0_u8_u5_n141, u0_u8_u5_n142, u0_u8_u5_n143, u0_u8_u5_n144, u0_u8_u5_n145, u0_u8_u5_n146, 
       u0_u8_u5_n147, u0_u8_u5_n148, u0_u8_u5_n149, u0_u8_u5_n150, u0_u8_u5_n151, u0_u8_u5_n152, u0_u8_u5_n153, u0_u8_u5_n154, u0_u8_u5_n155, 
       u0_u8_u5_n156, u0_u8_u5_n157, u0_u8_u5_n158, u0_u8_u5_n159, u0_u8_u5_n160, u0_u8_u5_n161, u0_u8_u5_n162, u0_u8_u5_n163, u0_u8_u5_n164, 
       u0_u8_u5_n165, u0_u8_u5_n166, u0_u8_u5_n167, u0_u8_u5_n168, u0_u8_u5_n169, u0_u8_u5_n170, u0_u8_u5_n171, u0_u8_u5_n172, u0_u8_u5_n173, 
       u0_u8_u5_n174, u0_u8_u5_n175, u0_u8_u5_n176, u0_u8_u5_n177, u0_u8_u5_n178, u0_u8_u5_n179, u0_u8_u5_n180, u0_u8_u5_n181, u0_u8_u5_n182, 
       u0_u8_u5_n183, u0_u8_u5_n184, u0_u8_u5_n185, u0_u8_u5_n186, u0_u8_u5_n187, u0_u8_u5_n188, u0_u8_u5_n189, u0_u8_u5_n190, u0_u8_u5_n191, 
       u0_u8_u5_n192, u0_u8_u5_n193, u0_u8_u5_n194, u0_u8_u5_n195, u0_u8_u5_n196, u0_u8_u5_n99, u0_u8_u6_n100, u0_u8_u6_n101, u0_u8_u6_n102, 
       u0_u8_u6_n103, u0_u8_u6_n104, u0_u8_u6_n105, u0_u8_u6_n106, u0_u8_u6_n107, u0_u8_u6_n108, u0_u8_u6_n109, u0_u8_u6_n110, u0_u8_u6_n111, 
       u0_u8_u6_n112, u0_u8_u6_n113, u0_u8_u6_n114, u0_u8_u6_n115, u0_u8_u6_n116, u0_u8_u6_n117, u0_u8_u6_n118, u0_u8_u6_n119, u0_u8_u6_n120, 
       u0_u8_u6_n121, u0_u8_u6_n122, u0_u8_u6_n123, u0_u8_u6_n124, u0_u8_u6_n125, u0_u8_u6_n126, u0_u8_u6_n127, u0_u8_u6_n128, u0_u8_u6_n129, 
       u0_u8_u6_n130, u0_u8_u6_n131, u0_u8_u6_n132, u0_u8_u6_n133, u0_u8_u6_n134, u0_u8_u6_n135, u0_u8_u6_n136, u0_u8_u6_n137, u0_u8_u6_n138, 
       u0_u8_u6_n139, u0_u8_u6_n140, u0_u8_u6_n141, u0_u8_u6_n142, u0_u8_u6_n143, u0_u8_u6_n144, u0_u8_u6_n145, u0_u8_u6_n146, u0_u8_u6_n147, 
       u0_u8_u6_n148, u0_u8_u6_n149, u0_u8_u6_n150, u0_u8_u6_n151, u0_u8_u6_n152, u0_u8_u6_n153, u0_u8_u6_n154, u0_u8_u6_n155, u0_u8_u6_n156, 
       u0_u8_u6_n157, u0_u8_u6_n158, u0_u8_u6_n159, u0_u8_u6_n160, u0_u8_u6_n161, u0_u8_u6_n162, u0_u8_u6_n163, u0_u8_u6_n164, u0_u8_u6_n165, 
       u0_u8_u6_n166, u0_u8_u6_n167, u0_u8_u6_n168, u0_u8_u6_n169, u0_u8_u6_n170, u0_u8_u6_n171, u0_u8_u6_n172, u0_u8_u6_n173, u0_u8_u6_n174, 
       u0_u8_u6_n88, u0_u8_u6_n89, u0_u8_u6_n90, u0_u8_u6_n91, u0_u8_u6_n92, u0_u8_u6_n93, u0_u8_u6_n94, u0_u8_u6_n95, u0_u8_u6_n96, 
       u0_u8_u6_n97, u0_u8_u6_n98, u0_u8_u6_n99, u0_uk_n718, u0_uk_n722, u0_uk_n723, u0_uk_n727, u0_uk_n729, u0_uk_n734, 
       u0_uk_n737, u0_uk_n741, u0_uk_n742, u0_uk_n747, u0_uk_n750, u0_uk_n751, u0_uk_n752, u0_uk_n753, u0_uk_n803, 
       u0_uk_n806, u0_uk_n887, u2_K10_1, u2_K10_2, u2_K10_27, u2_K10_28, u2_K10_29, u2_K10_3, u2_K10_45, 
       u2_K10_47, u2_K10_48, u2_K10_5, u2_K14_19, u2_K14_20, u2_K14_22, u2_K14_23, u2_K14_24, u2_K5_43, 
       u2_K5_45, u2_K5_46, u2_out13_1, u2_out13_10, u2_out13_20, u2_out13_26, u2_out4_15, u2_out4_21, u2_out4_27, 
       u2_out4_5, u2_out9_14, u2_out9_15, u2_out9_17, u2_out9_21, u2_out9_23, u2_out9_25, u2_out9_27, u2_out9_3, 
       u2_out9_31, u2_out9_5, u2_out9_8, u2_out9_9, u2_u13_X_19, u2_u13_X_20, u2_u13_X_21, u2_u13_X_22, u2_u13_X_23, 
       u2_u13_X_24, u2_u13_u3_n100, u2_u13_u3_n101, u2_u13_u3_n102, u2_u13_u3_n103, u2_u13_u3_n104, u2_u13_u3_n105, u2_u13_u3_n106, u2_u13_u3_n107, 
       u2_u13_u3_n108, u2_u13_u3_n109, u2_u13_u3_n110, u2_u13_u3_n111, u2_u13_u3_n112, u2_u13_u3_n113, u2_u13_u3_n114, u2_u13_u3_n115, u2_u13_u3_n116, 
       u2_u13_u3_n117, u2_u13_u3_n118, u2_u13_u3_n119, u2_u13_u3_n120, u2_u13_u3_n121, u2_u13_u3_n122, u2_u13_u3_n123, u2_u13_u3_n124, u2_u13_u3_n125, 
       u2_u13_u3_n126, u2_u13_u3_n127, u2_u13_u3_n128, u2_u13_u3_n129, u2_u13_u3_n130, u2_u13_u3_n131, u2_u13_u3_n132, u2_u13_u3_n133, u2_u13_u3_n134, 
       u2_u13_u3_n135, u2_u13_u3_n136, u2_u13_u3_n137, u2_u13_u3_n138, u2_u13_u3_n139, u2_u13_u3_n140, u2_u13_u3_n141, u2_u13_u3_n142, u2_u13_u3_n143, 
       u2_u13_u3_n144, u2_u13_u3_n145, u2_u13_u3_n146, u2_u13_u3_n147, u2_u13_u3_n148, u2_u13_u3_n149, u2_u13_u3_n150, u2_u13_u3_n151, u2_u13_u3_n152, 
       u2_u13_u3_n153, u2_u13_u3_n154, u2_u13_u3_n155, u2_u13_u3_n156, u2_u13_u3_n157, u2_u13_u3_n158, u2_u13_u3_n159, u2_u13_u3_n160, u2_u13_u3_n161, 
       u2_u13_u3_n162, u2_u13_u3_n163, u2_u13_u3_n164, u2_u13_u3_n165, u2_u13_u3_n166, u2_u13_u3_n167, u2_u13_u3_n168, u2_u13_u3_n169, u2_u13_u3_n170, 
       u2_u13_u3_n171, u2_u13_u3_n172, u2_u13_u3_n173, u2_u13_u3_n174, u2_u13_u3_n175, u2_u13_u3_n176, u2_u13_u3_n177, u2_u13_u3_n178, u2_u13_u3_n179, 
       u2_u13_u3_n180, u2_u13_u3_n181, u2_u13_u3_n182, u2_u13_u3_n183, u2_u13_u3_n184, u2_u13_u3_n185, u2_u13_u3_n186, u2_u13_u3_n94, u2_u13_u3_n95, 
       u2_u13_u3_n96, u2_u13_u3_n97, u2_u13_u3_n98, u2_u13_u3_n99, u2_u4_X_43, u2_u4_X_44, u2_u4_X_45, u2_u4_X_46, u2_u4_X_47, 
       u2_u4_X_48, u2_u4_u7_n100, u2_u4_u7_n101, u2_u4_u7_n102, u2_u4_u7_n103, u2_u4_u7_n104, u2_u4_u7_n105, u2_u4_u7_n106, u2_u4_u7_n107, 
       u2_u4_u7_n108, u2_u4_u7_n109, u2_u4_u7_n110, u2_u4_u7_n111, u2_u4_u7_n112, u2_u4_u7_n113, u2_u4_u7_n114, u2_u4_u7_n115, u2_u4_u7_n116, 
       u2_u4_u7_n117, u2_u4_u7_n118, u2_u4_u7_n119, u2_u4_u7_n120, u2_u4_u7_n121, u2_u4_u7_n122, u2_u4_u7_n123, u2_u4_u7_n124, u2_u4_u7_n125, 
       u2_u4_u7_n126, u2_u4_u7_n127, u2_u4_u7_n128, u2_u4_u7_n129, u2_u4_u7_n130, u2_u4_u7_n131, u2_u4_u7_n132, u2_u4_u7_n133, u2_u4_u7_n134, 
       u2_u4_u7_n135, u2_u4_u7_n136, u2_u4_u7_n137, u2_u4_u7_n138, u2_u4_u7_n139, u2_u4_u7_n140, u2_u4_u7_n141, u2_u4_u7_n142, u2_u4_u7_n143, 
       u2_u4_u7_n144, u2_u4_u7_n145, u2_u4_u7_n146, u2_u4_u7_n147, u2_u4_u7_n148, u2_u4_u7_n149, u2_u4_u7_n150, u2_u4_u7_n151, u2_u4_u7_n152, 
       u2_u4_u7_n153, u2_u4_u7_n154, u2_u4_u7_n155, u2_u4_u7_n156, u2_u4_u7_n157, u2_u4_u7_n158, u2_u4_u7_n159, u2_u4_u7_n160, u2_u4_u7_n161, 
       u2_u4_u7_n162, u2_u4_u7_n163, u2_u4_u7_n164, u2_u4_u7_n165, u2_u4_u7_n166, u2_u4_u7_n167, u2_u4_u7_n168, u2_u4_u7_n169, u2_u4_u7_n170, 
       u2_u4_u7_n171, u2_u4_u7_n172, u2_u4_u7_n173, u2_u4_u7_n174, u2_u4_u7_n175, u2_u4_u7_n176, u2_u4_u7_n177, u2_u4_u7_n178, u2_u4_u7_n179, 
       u2_u4_u7_n180, u2_u4_u7_n91, u2_u4_u7_n92, u2_u4_u7_n93, u2_u4_u7_n94, u2_u4_u7_n95, u2_u4_u7_n96, u2_u4_u7_n97, u2_u4_u7_n98, 
       u2_u4_u7_n99, u2_u9_X_1, u2_u9_X_2, u2_u9_X_25, u2_u9_X_26, u2_u9_X_27, u2_u9_X_28, u2_u9_X_29, u2_u9_X_3, 
       u2_u9_X_30, u2_u9_X_4, u2_u9_X_43, u2_u9_X_44, u2_u9_X_45, u2_u9_X_46, u2_u9_X_47, u2_u9_X_48, u2_u9_X_5, 
       u2_u9_X_6, u2_u9_u0_n100, u2_u9_u0_n101, u2_u9_u0_n102, u2_u9_u0_n103, u2_u9_u0_n104, u2_u9_u0_n105, u2_u9_u0_n106, u2_u9_u0_n107, 
       u2_u9_u0_n108, u2_u9_u0_n109, u2_u9_u0_n110, u2_u9_u0_n111, u2_u9_u0_n112, u2_u9_u0_n113, u2_u9_u0_n114, u2_u9_u0_n115, u2_u9_u0_n116, 
       u2_u9_u0_n117, u2_u9_u0_n118, u2_u9_u0_n119, u2_u9_u0_n120, u2_u9_u0_n121, u2_u9_u0_n122, u2_u9_u0_n123, u2_u9_u0_n124, u2_u9_u0_n125, 
       u2_u9_u0_n126, u2_u9_u0_n127, u2_u9_u0_n128, u2_u9_u0_n129, u2_u9_u0_n130, u2_u9_u0_n131, u2_u9_u0_n132, u2_u9_u0_n133, u2_u9_u0_n134, 
       u2_u9_u0_n135, u2_u9_u0_n136, u2_u9_u0_n137, u2_u9_u0_n138, u2_u9_u0_n139, u2_u9_u0_n140, u2_u9_u0_n141, u2_u9_u0_n142, u2_u9_u0_n143, 
       u2_u9_u0_n144, u2_u9_u0_n145, u2_u9_u0_n146, u2_u9_u0_n147, u2_u9_u0_n148, u2_u9_u0_n149, u2_u9_u0_n150, u2_u9_u0_n151, u2_u9_u0_n152, 
       u2_u9_u0_n153, u2_u9_u0_n154, u2_u9_u0_n155, u2_u9_u0_n156, u2_u9_u0_n157, u2_u9_u0_n158, u2_u9_u0_n159, u2_u9_u0_n160, u2_u9_u0_n161, 
       u2_u9_u0_n162, u2_u9_u0_n163, u2_u9_u0_n164, u2_u9_u0_n165, u2_u9_u0_n166, u2_u9_u0_n167, u2_u9_u0_n168, u2_u9_u0_n169, u2_u9_u0_n170, 
       u2_u9_u0_n171, u2_u9_u0_n172, u2_u9_u0_n173, u2_u9_u0_n174, u2_u9_u0_n88, u2_u9_u0_n89, u2_u9_u0_n90, u2_u9_u0_n91, u2_u9_u0_n92, 
       u2_u9_u0_n93, u2_u9_u0_n94, u2_u9_u0_n95, u2_u9_u0_n96, u2_u9_u0_n97, u2_u9_u0_n98, u2_u9_u0_n99, u2_u9_u4_n100, u2_u9_u4_n101, 
       u2_u9_u4_n102, u2_u9_u4_n103, u2_u9_u4_n104, u2_u9_u4_n105, u2_u9_u4_n106, u2_u9_u4_n107, u2_u9_u4_n108, u2_u9_u4_n109, u2_u9_u4_n110, 
       u2_u9_u4_n111, u2_u9_u4_n112, u2_u9_u4_n113, u2_u9_u4_n114, u2_u9_u4_n115, u2_u9_u4_n116, u2_u9_u4_n117, u2_u9_u4_n118, u2_u9_u4_n119, 
       u2_u9_u4_n120, u2_u9_u4_n121, u2_u9_u4_n122, u2_u9_u4_n123, u2_u9_u4_n124, u2_u9_u4_n125, u2_u9_u4_n126, u2_u9_u4_n127, u2_u9_u4_n128, 
       u2_u9_u4_n129, u2_u9_u4_n130, u2_u9_u4_n131, u2_u9_u4_n132, u2_u9_u4_n133, u2_u9_u4_n134, u2_u9_u4_n135, u2_u9_u4_n136, u2_u9_u4_n137, 
       u2_u9_u4_n138, u2_u9_u4_n139, u2_u9_u4_n140, u2_u9_u4_n141, u2_u9_u4_n142, u2_u9_u4_n143, u2_u9_u4_n144, u2_u9_u4_n145, u2_u9_u4_n146, 
       u2_u9_u4_n147, u2_u9_u4_n148, u2_u9_u4_n149, u2_u9_u4_n150, u2_u9_u4_n151, u2_u9_u4_n152, u2_u9_u4_n153, u2_u9_u4_n154, u2_u9_u4_n155, 
       u2_u9_u4_n156, u2_u9_u4_n157, u2_u9_u4_n158, u2_u9_u4_n159, u2_u9_u4_n160, u2_u9_u4_n161, u2_u9_u4_n162, u2_u9_u4_n163, u2_u9_u4_n164, 
       u2_u9_u4_n165, u2_u9_u4_n166, u2_u9_u4_n167, u2_u9_u4_n168, u2_u9_u4_n169, u2_u9_u4_n170, u2_u9_u4_n171, u2_u9_u4_n172, u2_u9_u4_n173, 
       u2_u9_u4_n174, u2_u9_u4_n175, u2_u9_u4_n176, u2_u9_u4_n177, u2_u9_u4_n178, u2_u9_u4_n179, u2_u9_u4_n180, u2_u9_u4_n181, u2_u9_u4_n182, 
       u2_u9_u4_n183, u2_u9_u4_n184, u2_u9_u4_n185, u2_u9_u4_n186, u2_u9_u4_n94, u2_u9_u4_n95, u2_u9_u4_n96, u2_u9_u4_n97, u2_u9_u4_n98, 
       u2_u9_u4_n99, u2_u9_u7_n100, u2_u9_u7_n101, u2_u9_u7_n102, u2_u9_u7_n103, u2_u9_u7_n104, u2_u9_u7_n105, u2_u9_u7_n106, u2_u9_u7_n107, 
       u2_u9_u7_n108, u2_u9_u7_n109, u2_u9_u7_n110, u2_u9_u7_n111, u2_u9_u7_n112, u2_u9_u7_n113, u2_u9_u7_n114, u2_u9_u7_n115, u2_u9_u7_n116, 
       u2_u9_u7_n117, u2_u9_u7_n118, u2_u9_u7_n119, u2_u9_u7_n120, u2_u9_u7_n121, u2_u9_u7_n122, u2_u9_u7_n123, u2_u9_u7_n124, u2_u9_u7_n125, 
       u2_u9_u7_n126, u2_u9_u7_n127, u2_u9_u7_n128, u2_u9_u7_n129, u2_u9_u7_n130, u2_u9_u7_n131, u2_u9_u7_n132, u2_u9_u7_n133, u2_u9_u7_n134, 
       u2_u9_u7_n135, u2_u9_u7_n136, u2_u9_u7_n137, u2_u9_u7_n138, u2_u9_u7_n139, u2_u9_u7_n140, u2_u9_u7_n141, u2_u9_u7_n142, u2_u9_u7_n143, 
       u2_u9_u7_n144, u2_u9_u7_n145, u2_u9_u7_n146, u2_u9_u7_n147, u2_u9_u7_n148, u2_u9_u7_n149, u2_u9_u7_n150, u2_u9_u7_n151, u2_u9_u7_n152, 
       u2_u9_u7_n153, u2_u9_u7_n154, u2_u9_u7_n155, u2_u9_u7_n156, u2_u9_u7_n157, u2_u9_u7_n158, u2_u9_u7_n159, u2_u9_u7_n160, u2_u9_u7_n161, 
       u2_u9_u7_n162, u2_u9_u7_n163, u2_u9_u7_n164, u2_u9_u7_n165, u2_u9_u7_n166, u2_u9_u7_n167, u2_u9_u7_n168, u2_u9_u7_n169, u2_u9_u7_n170, 
       u2_u9_u7_n171, u2_u9_u7_n172, u2_u9_u7_n173, u2_u9_u7_n174, u2_u9_u7_n175, u2_u9_u7_n176, u2_u9_u7_n177, u2_u9_u7_n178, u2_u9_u7_n179, 
       u2_u9_u7_n180, u2_u9_u7_n91, u2_u9_u7_n92, u2_u9_u7_n93, u2_u9_u7_n94, u2_u9_u7_n95, u2_u9_u7_n96, u2_u9_u7_n97, u2_u9_u7_n98, 
       u2_u9_u7_n99, u2_uk_n1053, u2_uk_n1054, u2_uk_n279, u2_uk_n286, u2_uk_n685,  u2_uk_n686;
  XOR2_X1 u0_U270 (.Z( u0_N29 ) , .B( u0_desIn_r_40 ) , .A( u0_out0_30 ) );
  XOR2_X1 u0_U273 (.B( u0_L7_32 ) , .Z( u0_N287 ) , .A( u0_out8_32 ) );
  XOR2_X1 u0_U274 (.B( u0_L7_31 ) , .Z( u0_N286 ) , .A( u0_out8_31 ) );
  XOR2_X1 u0_U275 (.B( u0_L7_30 ) , .Z( u0_N285 ) , .A( u0_out8_30 ) );
  XOR2_X1 u0_U276 (.B( u0_L7_29 ) , .Z( u0_N284 ) , .A( u0_out8_29 ) );
  XOR2_X1 u0_U277 (.B( u0_L7_28 ) , .Z( u0_N283 ) , .A( u0_out8_28 ) );
  XOR2_X1 u0_U282 (.B( u0_L7_24 ) , .Z( u0_N279 ) , .A( u0_out8_24 ) );
  XOR2_X1 u0_U283 (.B( u0_L7_23 ) , .Z( u0_N278 ) , .A( u0_out8_23 ) );
  XOR2_X1 u0_U284 (.B( u0_L7_22 ) , .Z( u0_N277 ) , .A( u0_out8_22 ) );
  XOR2_X1 u0_U287 (.B( u0_L7_19 ) , .Z( u0_N274 ) , .A( u0_out8_19 ) );
  XOR2_X1 u0_U288 (.B( u0_L7_18 ) , .Z( u0_N273 ) , .A( u0_out8_18 ) );
  XOR2_X1 u0_U289 (.B( u0_L7_17 ) , .Z( u0_N272 ) , .A( u0_out8_17 ) );
  XOR2_X1 u0_U290 (.B( u0_L7_16 ) , .Z( u0_N271 ) , .A( u0_out8_16 ) );
  XOR2_X1 u0_U294 (.B( u0_L7_13 ) , .Z( u0_N268 ) , .A( u0_out8_13 ) );
  XOR2_X1 u0_U295 (.B( u0_L7_12 ) , .Z( u0_N267 ) , .A( u0_out8_12 ) );
  XOR2_X1 u0_U296 (.B( u0_L7_11 ) , .Z( u0_N266 ) , .A( u0_out8_11 ) );
  XOR2_X1 u0_U298 (.B( u0_L7_9 ) , .Z( u0_N264 ) , .A( u0_out8_9 ) );
  XOR2_X1 u0_U300 (.B( u0_L7_7 ) , .Z( u0_N262 ) , .A( u0_out8_7 ) );
  XOR2_X1 u0_U301 (.B( u0_L7_6 ) , .Z( u0_N261 ) , .A( u0_out8_6 ) );
  XOR2_X1 u0_U304 (.B( u0_L7_4 ) , .Z( u0_N259 ) , .A( u0_out8_4 ) );
  XOR2_X1 u0_U306 (.B( u0_L7_2 ) , .Z( u0_N257 ) , .A( u0_out8_2 ) );
  XOR2_X1 u0_U308 (.B( u0_L6_32 ) , .Z( u0_N255 ) , .A( u0_out7_32 ) );
  XOR2_X1 u0_U311 (.B( u0_L6_29 ) , .Z( u0_N252 ) , .A( u0_out7_29 ) );
  XOR2_X1 u0_U316 (.B( u0_L6_25 ) , .Z( u0_N248 ) , .A( u0_out7_25 ) );
  XOR2_X1 u0_U319 (.B( u0_L6_22 ) , .Z( u0_N245 ) , .A( u0_out7_22 ) );
  XOR2_X1 u0_U322 (.B( u0_L6_19 ) , .Z( u0_N242 ) , .A( u0_out7_19 ) );
  XOR2_X1 u0_U328 (.B( u0_L6_14 ) , .Z( u0_N237 ) , .A( u0_out7_14 ) );
  XOR2_X1 u0_U330 (.B( u0_L6_12 ) , .Z( u0_N235 ) , .A( u0_out7_12 ) );
  XOR2_X1 u0_U331 (.B( u0_L6_11 ) , .Z( u0_N234 ) , .A( u0_out7_11 ) );
  XOR2_X1 u0_U334 (.B( u0_L6_8 ) , .Z( u0_N231 ) , .A( u0_out7_8 ) );
  XOR2_X1 u0_U335 (.B( u0_L6_7 ) , .Z( u0_N230 ) , .A( u0_out7_7 ) );
  XOR2_X1 u0_U336 (.Z( u0_N23 ) , .B( u0_desIn_r_58 ) , .A( u0_out0_24 ) );
  XOR2_X1 u0_U339 (.B( u0_L6_4 ) , .Z( u0_N227 ) , .A( u0_out7_4 ) );
  XOR2_X1 u0_U340 (.B( u0_L6_3 ) , .Z( u0_N226 ) , .A( u0_out7_3 ) );
  XOR2_X1 u0_U416 (.B( u0_L3_31 ) , .Z( u0_N158 ) , .A( u0_out4_31 ) );
  XOR2_X1 u0_U420 (.B( u0_L3_27 ) , .Z( u0_N154 ) , .A( u0_out4_27 ) );
  XOR2_X1 u0_U424 (.B( u0_L3_23 ) , .Z( u0_N150 ) , .A( u0_out4_23 ) );
  XOR2_X1 u0_U425 (.Z( u0_N15 ) , .B( u0_desIn_r_60 ) , .A( u0_out0_16 ) );
  XOR2_X1 u0_U427 (.B( u0_L3_21 ) , .Z( u0_N148 ) , .A( u0_out4_21 ) );
  XOR2_X1 u0_U431 (.B( u0_L3_17 ) , .Z( u0_N144 ) , .A( u0_out4_17 ) );
  XOR2_X1 u0_U433 (.B( u0_L3_15 ) , .Z( u0_N142 ) , .A( u0_out4_15 ) );
  XOR2_X1 u0_U440 (.B( u0_L3_9 ) , .Z( u0_N136 ) , .A( u0_out4_9 ) );
  XOR2_X1 u0_U444 (.B( u0_L3_5 ) , .Z( u0_N132 ) , .A( u0_out4_5 ) );
  XOR2_X1 u0_U57 (.Z( u0_N5 ) , .B( u0_desIn_r_46 ) , .A( u0_out0_6 ) );
  XOR2_X1 u0_u0_U40 (.B( u0_K1_18 ) , .A( u0_desIn_r_37 ) , .Z( u0_u0_X_18 ) );
  XOR2_X1 u0_u0_U41 (.B( u0_K1_17 ) , .A( u0_desIn_r_29 ) , .Z( u0_u0_X_17 ) );
  XOR2_X1 u0_u0_U42 (.B( u0_K1_16 ) , .A( u0_desIn_r_21 ) , .Z( u0_u0_X_16 ) );
  XOR2_X1 u0_u0_U43 (.B( u0_K1_15 ) , .A( u0_desIn_r_13 ) , .Z( u0_u0_X_15 ) );
  XOR2_X1 u0_u0_U44 (.B( u0_K1_14 ) , .A( u0_desIn_r_5 ) , .Z( u0_u0_X_14 ) );
  XOR2_X1 u0_u0_U45 (.B( u0_K1_13 ) , .A( u0_desIn_r_63 ) , .Z( u0_u0_X_13 ) );
  OAI22_X1 u0_u0_u2_U10 (.B2( u0_u0_u2_n21 ) , .ZN( u0_u0_u2_n29 ) , .A1( u0_u0_u2_n36 ) , .A2( u0_u0_u2_n37 ) , .B1( u0_u0_u2_n38 ) );
  NAND3_X1 u0_u0_u2_U100 (.A3( u0_u0_u2_n51 ) , .A1( u0_u0_u2_n85 ) , .A2( u0_u0_u2_n89 ) , .ZN( u0_u0_u2_n91 ) );
  NOR3_X1 u0_u0_u2_U11 (.A2( u0_u0_u2_n1 ) , .A3( u0_u0_u2_n14 ) , .ZN( u0_u0_u2_n38 ) , .A1( u0_u0_u2_n39 ) );
  AOI21_X1 u0_u0_u2_U12 (.A( u0_u0_u2_n18 ) , .B1( u0_u0_u2_n5 ) , .ZN( u0_u0_u2_n64 ) , .B2( u0_u0_u2_n66 ) );
  INV_X1 u0_u0_u2_U13 (.A( u0_u0_u2_n39 ) , .ZN( u0_u0_u2_n5 ) );
  AOI21_X1 u0_u0_u2_U14 (.A( u0_u0_u2_n17 ) , .B2( u0_u0_u2_n34 ) , .B1( u0_u0_u2_n4 ) , .ZN( u0_u0_u2_n45 ) );
  AOI21_X1 u0_u0_u2_U15 (.A( u0_u0_u2_n18 ) , .B1( u0_u0_u2_n37 ) , .ZN( u0_u0_u2_n44 ) , .B2( u0_u0_u2_n46 ) );
  INV_X1 u0_u0_u2_U16 (.ZN( u0_u0_u2_n18 ) , .A( u0_u0_u2_n33 ) );
  INV_X1 u0_u0_u2_U17 (.ZN( u0_u0_u2_n1 ) , .A( u0_u0_u2_n69 ) );
  NAND2_X1 u0_u0_u2_U18 (.A1( u0_u0_u2_n37 ) , .ZN( u0_u0_u2_n39 ) , .A2( u0_u0_u2_n67 ) );
  INV_X1 u0_u0_u2_U19 (.ZN( u0_u0_u2_n19 ) , .A( u0_u0_u2_n36 ) );
  INV_X1 u0_u0_u2_U20 (.ZN( u0_u0_u2_n16 ) , .A( u0_u0_u2_n52 ) );
  NAND2_X1 u0_u0_u2_U21 (.ZN( u0_u0_u2_n32 ) , .A2( u0_u0_u2_n50 ) , .A1( u0_u0_u2_n57 ) );
  INV_X1 u0_u0_u2_U22 (.ZN( u0_u0_u2_n11 ) , .A( u0_u0_u2_n76 ) );
  INV_X1 u0_u0_u2_U23 (.ZN( u0_u0_u2_n14 ) , .A( u0_u0_u2_n50 ) );
  INV_X1 u0_u0_u2_U24 (.A( u0_u0_u2_n34 ) , .ZN( u0_u0_u2_n8 ) );
  INV_X1 u0_u0_u2_U25 (.ZN( u0_u0_u2_n12 ) , .A( u0_u0_u2_n70 ) );
  INV_X1 u0_u0_u2_U26 (.A( u0_u0_u2_n73 ) , .ZN( u0_u0_u2_n9 ) );
  INV_X1 u0_u0_u2_U27 (.ZN( u0_u0_u2_n10 ) , .A( u0_u0_u2_n58 ) );
  INV_X1 u0_u0_u2_U28 (.ZN( u0_u0_u2_n13 ) , .A( u0_u0_u2_n35 ) );
  NAND2_X1 u0_u0_u2_U29 (.ZN( u0_u0_u2_n71 ) , .A1( u0_u0_u2_n72 ) , .A2( u0_u0_u2_n73 ) );
  NOR2_X1 u0_u0_u2_U3 (.A2( u0_u0_u2_n12 ) , .ZN( u0_u0_u2_n68 ) , .A1( u0_u0_u2_n9 ) );
  INV_X1 u0_u0_u2_U30 (.A( u0_u0_u2_n57 ) , .ZN( u0_u0_u2_n7 ) );
  INV_X1 u0_u0_u2_U31 (.A( u0_u0_u2_n31 ) , .ZN( u0_u0_u2_n6 ) );
  OAI21_X1 u0_u0_u2_U32 (.B2( u0_u0_u2_n10 ) , .ZN( u0_u0_u2_n31 ) , .B1( u0_u0_u2_n32 ) , .A( u0_u0_u2_n33 ) );
  NOR2_X1 u0_u0_u2_U33 (.A2( u0_u0_u2_n20 ) , .A1( u0_u0_u2_n23 ) , .ZN( u0_u0_u2_n33 ) );
  NOR2_X1 u0_u0_u2_U34 (.A1( u0_u0_u2_n49 ) , .ZN( u0_u0_u2_n52 ) , .A2( u0_u0_u2_n75 ) );
  NOR2_X1 u0_u0_u2_U35 (.A1( u0_u0_u2_n33 ) , .ZN( u0_u0_u2_n36 ) , .A2( u0_u0_u2_n51 ) );
  AOI211_X1 u0_u0_u2_U36 (.C2( u0_u0_u2_n10 ) , .C1( u0_u0_u2_n51 ) , .ZN( u0_u0_u2_n59 ) , .A( u0_u0_u2_n92 ) , .B( u0_u0_u2_n93 ) );
  OAI22_X1 u0_u0_u2_U37 (.B2( u0_u0_u2_n21 ) , .A1( u0_u0_u2_n37 ) , .A2( u0_u0_u2_n52 ) , .B1( u0_u0_u2_n56 ) , .ZN( u0_u0_u2_n92 ) );
  OAI221_X1 u0_u0_u2_U38 (.C2( u0_u0_u2_n17 ) , .B2( u0_u0_u2_n18 ) , .A( u0_u0_u2_n40 ) , .C1( u0_u0_u2_n57 ) , .B1( u0_u0_u2_n76 ) , .ZN( u0_u0_u2_n93 ) );
  OAI221_X1 u0_u0_u2_U39 (.C1( u0_u0_u2_n21 ) , .ZN( u0_u0_u2_n26 ) , .B1( u0_u0_u2_n36 ) , .B2( u0_u0_u2_n46 ) , .C2( u0_u0_u2_n66 ) , .A( u0_u0_u2_n74 ) );
  INV_X1 u0_u0_u2_U4 (.ZN( u0_u0_u2_n4 ) , .A( u0_u0_u2_n55 ) );
  OAI21_X1 u0_u0_u2_U40 (.B2( u0_u0_u2_n11 ) , .B1( u0_u0_u2_n13 ) , .ZN( u0_u0_u2_n74 ) , .A( u0_u0_u2_n75 ) );
  OAI221_X1 u0_u0_u2_U41 (.C2( u0_u0_u2_n22 ) , .ZN( u0_u0_u2_n27 ) , .C1( u0_u0_u2_n4 ) , .B1( u0_u0_u2_n52 ) , .B2( u0_u0_u2_n53 ) , .A( u0_u0_u2_n54 ) );
  AND3_X1 u0_u0_u2_U42 (.ZN( u0_u0_u2_n53 ) , .A1( u0_u0_u2_n56 ) , .A2( u0_u0_u2_n57 ) , .A3( u0_u0_u2_n58 ) );
  AOI22_X1 u0_u0_u2_U43 (.A2( u0_u0_u2_n1 ) , .A1( u0_u0_u2_n33 ) , .B1( u0_u0_u2_n49 ) , .ZN( u0_u0_u2_n54 ) , .B2( u0_u0_u2_n9 ) );
  AOI21_X1 u0_u0_u2_U44 (.B2( u0_u0_u2_n1 ) , .B1( u0_u0_u2_n16 ) , .ZN( u0_u0_u2_n40 ) , .A( u0_u0_u2_n94 ) );
  AND3_X1 u0_u0_u2_U45 (.A3( u0_u0_u2_n33 ) , .A1( u0_u0_u2_n85 ) , .A2( u0_u0_u2_n89 ) , .ZN( u0_u0_u2_n94 ) );
  OAI21_X1 u0_u0_u2_U46 (.B1( u0_u0_u2_n36 ) , .ZN( u0_u0_u2_n43 ) , .B2( u0_u0_u2_n47 ) , .A( u0_u0_u2_n48 ) );
  OAI21_X1 u0_u0_u2_U47 (.B2( u0_u0_u2_n12 ) , .B1( u0_u0_u2_n13 ) , .ZN( u0_u0_u2_n48 ) , .A( u0_u0_u2_n49 ) );
  NOR3_X1 u0_u0_u2_U48 (.A2( u0_u0_u2_n11 ) , .A3( u0_u0_u2_n14 ) , .ZN( u0_u0_u2_n47 ) , .A1( u0_u0_u2_n8 ) );
  OAI21_X1 u0_u0_u2_U49 (.ZN( u0_u0_u2_n25 ) , .B1( u0_u0_u2_n36 ) , .B2( u0_u0_u2_n68 ) , .A( u0_u0_u2_n88 ) );
  NOR4_X1 u0_u0_u2_U5 (.ZN( u0_u0_u2_n61 ) , .A1( u0_u0_u2_n62 ) , .A2( u0_u0_u2_n63 ) , .A3( u0_u0_u2_n64 ) , .A4( u0_u0_u2_n65 ) );
  NAND2_X1 u0_u0_u2_U50 (.ZN( u0_u0_u2_n34 ) , .A1( u0_u0_u2_n82 ) , .A2( u0_u0_u2_n89 ) );
  NAND2_X1 u0_u0_u2_U51 (.ZN( u0_u0_u2_n46 ) , .A1( u0_u0_u2_n81 ) , .A2( u0_u0_u2_n84 ) );
  NAND2_X1 u0_u0_u2_U52 (.ZN( u0_u0_u2_n37 ) , .A2( u0_u0_u2_n83 ) , .A1( u0_u0_u2_n85 ) );
  NAND2_X1 u0_u0_u2_U53 (.ZN( u0_u0_u2_n57 ) , .A2( u0_u0_u2_n84 ) , .A1( u0_u0_u2_n89 ) );
  INV_X1 u0_u0_u2_U54 (.ZN( u0_u0_u2_n21 ) , .A( u0_u0_u2_n49 ) );
  INV_X1 u0_u0_u2_U55 (.ZN( u0_u0_u2_n22 ) , .A( u0_u0_u2_n51 ) );
  NAND2_X1 u0_u0_u2_U56 (.ZN( u0_u0_u2_n76 ) , .A2( u0_u0_u2_n83 ) , .A1( u0_u0_u2_n87 ) );
  NAND2_X1 u0_u0_u2_U57 (.ZN( u0_u0_u2_n58 ) , .A2( u0_u0_u2_n82 ) , .A1( u0_u0_u2_n83 ) );
  NAND2_X1 u0_u0_u2_U58 (.ZN( u0_u0_u2_n50 ) , .A2( u0_u0_u2_n82 ) , .A1( u0_u0_u2_n86 ) );
  NAND2_X1 u0_u0_u2_U59 (.ZN( u0_u0_u2_n56 ) , .A2( u0_u0_u2_n84 ) , .A1( u0_u0_u2_n86 ) );
  AOI21_X1 u0_u0_u2_U6 (.B1( u0_u0_u2_n34 ) , .A( u0_u0_u2_n52 ) , .ZN( u0_u0_u2_n62 ) , .B2( u0_u0_u2_n70 ) );
  NAND2_X1 u0_u0_u2_U60 (.ZN( u0_u0_u2_n35 ) , .A2( u0_u0_u2_n86 ) , .A1( u0_u0_u2_n87 ) );
  NAND2_X1 u0_u0_u2_U61 (.ZN( u0_u0_u2_n70 ) , .A1( u0_u0_u2_n85 ) , .A2( u0_u0_u2_n86 ) );
  NAND2_X1 u0_u0_u2_U62 (.ZN( u0_u0_u2_n66 ) , .A1( u0_u0_u2_n81 ) , .A2( u0_u0_u2_n82 ) );
  NAND2_X1 u0_u0_u2_U63 (.ZN( u0_u0_u2_n67 ) , .A2( u0_u0_u2_n81 ) , .A1( u0_u0_u2_n85 ) );
  INV_X1 u0_u0_u2_U64 (.ZN( u0_u0_u2_n17 ) , .A( u0_u0_u2_n75 ) );
  NAND2_X1 u0_u0_u2_U65 (.ZN( u0_u0_u2_n73 ) , .A1( u0_u0_u2_n87 ) , .A2( u0_u0_u2_n89 ) );
  NAND2_X1 u0_u0_u2_U66 (.ZN( u0_u0_u2_n69 ) , .A2( u0_u0_u2_n81 ) , .A1( u0_u0_u2_n87 ) );
  NAND2_X1 u0_u0_u2_U67 (.ZN( u0_u0_u2_n72 ) , .A1( u0_u0_u2_n83 ) , .A2( u0_u0_u2_n84 ) );
  INV_X1 u0_u0_u2_U68 (.ZN( u0_u0_u2_n2 ) , .A( u0_u0_u2_n90 ) );
  OAI21_X1 u0_u0_u2_U69 (.B2( u0_u0_u2_n46 ) , .B1( u0_u0_u2_n52 ) , .ZN( u0_u0_u2_n90 ) , .A( u0_u0_u2_n91 ) );
  AOI21_X1 u0_u0_u2_U7 (.A( u0_u0_u2_n17 ) , .B2( u0_u0_u2_n46 ) , .B1( u0_u0_u2_n58 ) , .ZN( u0_u0_u2_n65 ) );
  NOR2_X1 u0_u0_u2_U70 (.A2( u0_u0_X_16 ) , .A1( u0_u0_u2_n23 ) , .ZN( u0_u0_u2_n49 ) );
  NOR2_X1 u0_u0_u2_U71 (.A2( u0_u0_X_13 ) , .A1( u0_u0_X_14 ) , .ZN( u0_u0_u2_n89 ) );
  NOR2_X1 u0_u0_u2_U72 (.A2( u0_u0_X_16 ) , .A1( u0_u0_X_17 ) , .ZN( u0_u0_u2_n51 ) );
  NOR2_X1 u0_u0_u2_U73 (.A2( u0_u0_X_15 ) , .A1( u0_u0_X_18 ) , .ZN( u0_u0_u2_n85 ) );
  NOR2_X1 u0_u0_u2_U74 (.A2( u0_u0_X_14 ) , .A1( u0_u0_u2_n15 ) , .ZN( u0_u0_u2_n86 ) );
  NOR2_X1 u0_u0_u2_U75 (.A2( u0_u0_X_15 ) , .A1( u0_u0_u2_n24 ) , .ZN( u0_u0_u2_n87 ) );
  NOR2_X1 u0_u0_u2_U76 (.A2( u0_u0_X_17 ) , .A1( u0_u0_u2_n20 ) , .ZN( u0_u0_u2_n75 ) );
  AND2_X1 u0_u0_u2_U77 (.A1( u0_u0_X_15 ) , .A2( u0_u0_u2_n24 ) , .ZN( u0_u0_u2_n84 ) );
  AND2_X1 u0_u0_u2_U78 (.A2( u0_u0_X_15 ) , .A1( u0_u0_X_18 ) , .ZN( u0_u0_u2_n82 ) );
  AND2_X1 u0_u0_u2_U79 (.A1( u0_u0_X_14 ) , .A2( u0_u0_u2_n15 ) , .ZN( u0_u0_u2_n83 ) );
  AOI21_X1 u0_u0_u2_U8 (.A( u0_u0_u2_n22 ) , .ZN( u0_u0_u2_n63 ) , .B1( u0_u0_u2_n68 ) , .B2( u0_u0_u2_n69 ) );
  AND2_X1 u0_u0_u2_U80 (.A1( u0_u0_X_13 ) , .A2( u0_u0_X_14 ) , .ZN( u0_u0_u2_n81 ) );
  INV_X1 u0_u0_u2_U81 (.A( u0_u0_X_16 ) , .ZN( u0_u0_u2_n20 ) );
  INV_X1 u0_u0_u2_U82 (.A( u0_u0_X_17 ) , .ZN( u0_u0_u2_n23 ) );
  INV_X1 u0_u0_u2_U83 (.A( u0_u0_X_13 ) , .ZN( u0_u0_u2_n15 ) );
  INV_X1 u0_u0_u2_U84 (.A( u0_u0_X_18 ) , .ZN( u0_u0_u2_n24 ) );
  NAND4_X1 u0_u0_u2_U85 (.ZN( u0_out0_30 ) , .A1( u0_u0_u2_n2 ) , .A2( u0_u0_u2_n40 ) , .A3( u0_u0_u2_n41 ) , .A4( u0_u0_u2_n42 ) );
  NOR3_X1 u0_u0_u2_U86 (.ZN( u0_u0_u2_n42 ) , .A1( u0_u0_u2_n43 ) , .A2( u0_u0_u2_n44 ) , .A3( u0_u0_u2_n45 ) );
  AOI21_X1 u0_u0_u2_U87 (.A( u0_u0_u2_n27 ) , .ZN( u0_u0_u2_n41 ) , .B2( u0_u0_u2_n51 ) , .B1( u0_u0_u2_n7 ) );
  NAND4_X1 u0_u0_u2_U88 (.ZN( u0_out0_24 ) , .A2( u0_u0_u2_n2 ) , .A1( u0_u0_u2_n59 ) , .A3( u0_u0_u2_n77 ) , .A4( u0_u0_u2_n78 ) );
  AOI221_X1 u0_u0_u2_U89 (.B2( u0_u0_u2_n16 ) , .C2( u0_u0_u2_n19 ) , .C1( u0_u0_u2_n55 ) , .ZN( u0_u0_u2_n78 ) , .B1( u0_u0_u2_n79 ) , .A( u0_u0_u2_n80 ) );
  OAI22_X1 u0_u0_u2_U9 (.A1( u0_u0_u2_n21 ) , .B1( u0_u0_u2_n22 ) , .B2( u0_u0_u2_n56 ) , .A2( u0_u0_u2_n76 ) , .ZN( u0_u0_u2_n80 ) );
  AOI21_X1 u0_u0_u2_U90 (.A( u0_u0_u2_n25 ) , .B2( u0_u0_u2_n33 ) , .ZN( u0_u0_u2_n77 ) , .B1( u0_u0_u2_n8 ) );
  NAND4_X1 u0_u0_u2_U91 (.ZN( u0_out0_16 ) , .A2( u0_u0_u2_n3 ) , .A1( u0_u0_u2_n59 ) , .A3( u0_u0_u2_n60 ) , .A4( u0_u0_u2_n61 ) );
  AOI22_X1 u0_u0_u2_U92 (.B2( u0_u0_u2_n19 ) , .B1( u0_u0_u2_n32 ) , .A1( u0_u0_u2_n49 ) , .ZN( u0_u0_u2_n60 ) , .A2( u0_u0_u2_n71 ) );
  INV_X1 u0_u0_u2_U93 (.A( u0_u0_u2_n26 ) , .ZN( u0_u0_u2_n3 ) );
  OR4_X1 u0_u0_u2_U94 (.ZN( u0_out0_6 ) , .A1( u0_u0_u2_n25 ) , .A2( u0_u0_u2_n26 ) , .A3( u0_u0_u2_n27 ) , .A4( u0_u0_u2_n28 ) );
  OR3_X1 u0_u0_u2_U95 (.ZN( u0_u0_u2_n28 ) , .A1( u0_u0_u2_n29 ) , .A2( u0_u0_u2_n30 ) , .A3( u0_u0_u2_n6 ) );
  AOI21_X1 u0_u0_u2_U96 (.A( u0_u0_u2_n22 ) , .ZN( u0_u0_u2_n30 ) , .B1( u0_u0_u2_n34 ) , .B2( u0_u0_u2_n35 ) );
  NAND3_X1 u0_u0_u2_U97 (.ZN( u0_u0_u2_n55 ) , .A3( u0_u0_u2_n66 ) , .A1( u0_u0_u2_n67 ) , .A2( u0_u0_u2_n72 ) );
  NAND3_X1 u0_u0_u2_U98 (.A1( u0_u0_u2_n35 ) , .A3( u0_u0_u2_n50 ) , .A2( u0_u0_u2_n58 ) , .ZN( u0_u0_u2_n79 ) );
  NAND3_X1 u0_u0_u2_U99 (.A3( u0_u0_u2_n75 ) , .A1( u0_u0_u2_n85 ) , .ZN( u0_u0_u2_n88 ) , .A2( u0_u0_u2_n89 ) );
  XOR2_X1 u0_u4_U10 (.B( u0_K5_45 ) , .A( u0_R3_30 ) , .Z( u0_u4_X_45 ) );
  XOR2_X1 u0_u4_U11 (.B( u0_K5_44 ) , .A( u0_R3_29 ) , .Z( u0_u4_X_44 ) );
  XOR2_X1 u0_u4_U12 (.B( u0_K5_43 ) , .A( u0_R3_28 ) , .Z( u0_u4_X_43 ) );
  XOR2_X1 u0_u4_U16 (.B( u0_K5_3 ) , .A( u0_R3_2 ) , .Z( u0_u4_X_3 ) );
  XOR2_X1 u0_u4_U27 (.B( u0_K5_2 ) , .A( u0_R3_1 ) , .Z( u0_u4_X_2 ) );
  XOR2_X1 u0_u4_U38 (.B( u0_K5_1 ) , .A( u0_R3_32 ) , .Z( u0_u4_X_1 ) );
  XOR2_X1 u0_u4_U4 (.B( u0_K5_6 ) , .A( u0_R3_5 ) , .Z( u0_u4_X_6 ) );
  XOR2_X1 u0_u4_U5 (.B( u0_K5_5 ) , .A( u0_R3_4 ) , .Z( u0_u4_X_5 ) );
  XOR2_X1 u0_u4_U6 (.B( u0_K5_4 ) , .A( u0_R3_3 ) , .Z( u0_u4_X_4 ) );
  XOR2_X1 u0_u4_U7 (.B( u0_K5_48 ) , .A( u0_R3_1 ) , .Z( u0_u4_X_48 ) );
  XOR2_X1 u0_u4_U8 (.B( u0_K5_47 ) , .A( u0_R3_32 ) , .Z( u0_u4_X_47 ) );
  XOR2_X1 u0_u4_U9 (.B( u0_K5_46 ) , .A( u0_R3_31 ) , .Z( u0_u4_X_46 ) );
  AND3_X1 u0_u4_u0_U10 (.A2( u0_u4_u0_n112 ) , .ZN( u0_u4_u0_n127 ) , .A3( u0_u4_u0_n130 ) , .A1( u0_u4_u0_n148 ) );
  NAND2_X1 u0_u4_u0_U11 (.ZN( u0_u4_u0_n113 ) , .A1( u0_u4_u0_n139 ) , .A2( u0_u4_u0_n149 ) );
  AND2_X1 u0_u4_u0_U12 (.ZN( u0_u4_u0_n107 ) , .A1( u0_u4_u0_n130 ) , .A2( u0_u4_u0_n140 ) );
  AND2_X1 u0_u4_u0_U13 (.A2( u0_u4_u0_n129 ) , .A1( u0_u4_u0_n130 ) , .ZN( u0_u4_u0_n151 ) );
  AND2_X1 u0_u4_u0_U14 (.A1( u0_u4_u0_n108 ) , .A2( u0_u4_u0_n125 ) , .ZN( u0_u4_u0_n145 ) );
  INV_X1 u0_u4_u0_U15 (.A( u0_u4_u0_n143 ) , .ZN( u0_u4_u0_n173 ) );
  NOR2_X1 u0_u4_u0_U16 (.A2( u0_u4_u0_n136 ) , .ZN( u0_u4_u0_n147 ) , .A1( u0_u4_u0_n160 ) );
  INV_X1 u0_u4_u0_U17 (.ZN( u0_u4_u0_n172 ) , .A( u0_u4_u0_n88 ) );
  OAI222_X1 u0_u4_u0_U18 (.C1( u0_u4_u0_n108 ) , .A1( u0_u4_u0_n125 ) , .B2( u0_u4_u0_n128 ) , .B1( u0_u4_u0_n144 ) , .A2( u0_u4_u0_n158 ) , .C2( u0_u4_u0_n161 ) , .ZN( u0_u4_u0_n88 ) );
  AOI21_X1 u0_u4_u0_U19 (.B1( u0_u4_u0_n103 ) , .ZN( u0_u4_u0_n132 ) , .A( u0_u4_u0_n165 ) , .B2( u0_u4_u0_n93 ) );
  INV_X1 u0_u4_u0_U20 (.A( u0_u4_u0_n142 ) , .ZN( u0_u4_u0_n165 ) );
  OAI221_X1 u0_u4_u0_U21 (.C1( u0_u4_u0_n112 ) , .ZN( u0_u4_u0_n120 ) , .B1( u0_u4_u0_n138 ) , .B2( u0_u4_u0_n141 ) , .C2( u0_u4_u0_n147 ) , .A( u0_u4_u0_n172 ) );
  AOI211_X1 u0_u4_u0_U22 (.B( u0_u4_u0_n115 ) , .A( u0_u4_u0_n116 ) , .C2( u0_u4_u0_n117 ) , .C1( u0_u4_u0_n118 ) , .ZN( u0_u4_u0_n119 ) );
  OAI22_X1 u0_u4_u0_U23 (.B1( u0_u4_u0_n125 ) , .ZN( u0_u4_u0_n126 ) , .A1( u0_u4_u0_n138 ) , .A2( u0_u4_u0_n146 ) , .B2( u0_u4_u0_n147 ) );
  OAI22_X1 u0_u4_u0_U24 (.B1( u0_u4_u0_n131 ) , .A1( u0_u4_u0_n144 ) , .B2( u0_u4_u0_n147 ) , .A2( u0_u4_u0_n90 ) , .ZN( u0_u4_u0_n91 ) );
  AND3_X1 u0_u4_u0_U25 (.A3( u0_u4_u0_n121 ) , .A2( u0_u4_u0_n125 ) , .A1( u0_u4_u0_n148 ) , .ZN( u0_u4_u0_n90 ) );
  INV_X1 u0_u4_u0_U26 (.A( u0_u4_u0_n136 ) , .ZN( u0_u4_u0_n161 ) );
  AOI22_X1 u0_u4_u0_U27 (.B2( u0_u4_u0_n109 ) , .A2( u0_u4_u0_n110 ) , .ZN( u0_u4_u0_n111 ) , .B1( u0_u4_u0_n118 ) , .A1( u0_u4_u0_n160 ) );
  INV_X1 u0_u4_u0_U28 (.A( u0_u4_u0_n118 ) , .ZN( u0_u4_u0_n158 ) );
  AOI21_X1 u0_u4_u0_U29 (.ZN( u0_u4_u0_n104 ) , .B1( u0_u4_u0_n107 ) , .B2( u0_u4_u0_n141 ) , .A( u0_u4_u0_n144 ) );
  INV_X1 u0_u4_u0_U3 (.A( u0_u4_u0_n113 ) , .ZN( u0_u4_u0_n166 ) );
  AOI21_X1 u0_u4_u0_U30 (.B1( u0_u4_u0_n127 ) , .B2( u0_u4_u0_n129 ) , .A( u0_u4_u0_n138 ) , .ZN( u0_u4_u0_n96 ) );
  AOI21_X1 u0_u4_u0_U31 (.ZN( u0_u4_u0_n116 ) , .B2( u0_u4_u0_n142 ) , .A( u0_u4_u0_n144 ) , .B1( u0_u4_u0_n166 ) );
  NAND2_X1 u0_u4_u0_U32 (.A1( u0_u4_u0_n102 ) , .ZN( u0_u4_u0_n128 ) , .A2( u0_u4_u0_n95 ) );
  NAND2_X1 u0_u4_u0_U33 (.A1( u0_u4_u0_n100 ) , .A2( u0_u4_u0_n103 ) , .ZN( u0_u4_u0_n125 ) );
  NAND2_X1 u0_u4_u0_U34 (.ZN( u0_u4_u0_n148 ) , .A1( u0_u4_u0_n93 ) , .A2( u0_u4_u0_n95 ) );
  NAND2_X1 u0_u4_u0_U35 (.A1( u0_u4_u0_n101 ) , .A2( u0_u4_u0_n102 ) , .ZN( u0_u4_u0_n150 ) );
  INV_X1 u0_u4_u0_U36 (.A( u0_u4_u0_n138 ) , .ZN( u0_u4_u0_n160 ) );
  NAND2_X1 u0_u4_u0_U37 (.A1( u0_u4_u0_n100 ) , .ZN( u0_u4_u0_n129 ) , .A2( u0_u4_u0_n95 ) );
  NAND2_X1 u0_u4_u0_U38 (.A2( u0_u4_u0_n102 ) , .A1( u0_u4_u0_n103 ) , .ZN( u0_u4_u0_n149 ) );
  NAND2_X1 u0_u4_u0_U39 (.A2( u0_u4_u0_n100 ) , .A1( u0_u4_u0_n101 ) , .ZN( u0_u4_u0_n139 ) );
  AOI21_X1 u0_u4_u0_U4 (.B1( u0_u4_u0_n114 ) , .ZN( u0_u4_u0_n115 ) , .B2( u0_u4_u0_n129 ) , .A( u0_u4_u0_n161 ) );
  NAND2_X1 u0_u4_u0_U40 (.A2( u0_u4_u0_n100 ) , .ZN( u0_u4_u0_n131 ) , .A1( u0_u4_u0_n92 ) );
  NAND2_X1 u0_u4_u0_U41 (.A2( u0_u4_u0_n102 ) , .ZN( u0_u4_u0_n114 ) , .A1( u0_u4_u0_n92 ) );
  NAND2_X1 u0_u4_u0_U42 (.A2( u0_u4_u0_n101 ) , .ZN( u0_u4_u0_n121 ) , .A1( u0_u4_u0_n93 ) );
  NAND2_X1 u0_u4_u0_U43 (.ZN( u0_u4_u0_n112 ) , .A2( u0_u4_u0_n92 ) , .A1( u0_u4_u0_n93 ) );
  OR3_X1 u0_u4_u0_U44 (.A3( u0_u4_u0_n152 ) , .A2( u0_u4_u0_n153 ) , .A1( u0_u4_u0_n154 ) , .ZN( u0_u4_u0_n155 ) );
  AOI21_X1 u0_u4_u0_U45 (.B2( u0_u4_u0_n150 ) , .B1( u0_u4_u0_n151 ) , .ZN( u0_u4_u0_n152 ) , .A( u0_u4_u0_n158 ) );
  AOI21_X1 u0_u4_u0_U46 (.A( u0_u4_u0_n144 ) , .B2( u0_u4_u0_n145 ) , .B1( u0_u4_u0_n146 ) , .ZN( u0_u4_u0_n154 ) );
  AOI21_X1 u0_u4_u0_U47 (.A( u0_u4_u0_n147 ) , .B2( u0_u4_u0_n148 ) , .B1( u0_u4_u0_n149 ) , .ZN( u0_u4_u0_n153 ) );
  INV_X1 u0_u4_u0_U48 (.ZN( u0_u4_u0_n171 ) , .A( u0_u4_u0_n99 ) );
  OAI211_X1 u0_u4_u0_U49 (.C2( u0_u4_u0_n140 ) , .C1( u0_u4_u0_n161 ) , .A( u0_u4_u0_n169 ) , .B( u0_u4_u0_n98 ) , .ZN( u0_u4_u0_n99 ) );
  AOI21_X1 u0_u4_u0_U5 (.B2( u0_u4_u0_n131 ) , .ZN( u0_u4_u0_n134 ) , .B1( u0_u4_u0_n151 ) , .A( u0_u4_u0_n158 ) );
  AOI211_X1 u0_u4_u0_U50 (.C1( u0_u4_u0_n118 ) , .A( u0_u4_u0_n123 ) , .B( u0_u4_u0_n96 ) , .C2( u0_u4_u0_n97 ) , .ZN( u0_u4_u0_n98 ) );
  INV_X1 u0_u4_u0_U51 (.ZN( u0_u4_u0_n169 ) , .A( u0_u4_u0_n91 ) );
  NOR2_X1 u0_u4_u0_U52 (.A2( u0_u4_X_6 ) , .ZN( u0_u4_u0_n100 ) , .A1( u0_u4_u0_n162 ) );
  NOR2_X1 u0_u4_u0_U53 (.A2( u0_u4_X_4 ) , .A1( u0_u4_X_5 ) , .ZN( u0_u4_u0_n118 ) );
  NOR2_X1 u0_u4_u0_U54 (.A2( u0_u4_X_2 ) , .ZN( u0_u4_u0_n103 ) , .A1( u0_u4_u0_n164 ) );
  NOR2_X1 u0_u4_u0_U55 (.A2( u0_u4_X_1 ) , .A1( u0_u4_X_2 ) , .ZN( u0_u4_u0_n92 ) );
  NOR2_X1 u0_u4_u0_U56 (.A2( u0_u4_X_1 ) , .ZN( u0_u4_u0_n101 ) , .A1( u0_u4_u0_n163 ) );
  NAND2_X1 u0_u4_u0_U57 (.A2( u0_u4_X_4 ) , .A1( u0_u4_X_5 ) , .ZN( u0_u4_u0_n144 ) );
  NOR2_X1 u0_u4_u0_U58 (.A2( u0_u4_X_5 ) , .ZN( u0_u4_u0_n136 ) , .A1( u0_u4_u0_n159 ) );
  NAND2_X1 u0_u4_u0_U59 (.A1( u0_u4_X_5 ) , .ZN( u0_u4_u0_n138 ) , .A2( u0_u4_u0_n159 ) );
  NOR2_X1 u0_u4_u0_U6 (.A1( u0_u4_u0_n108 ) , .ZN( u0_u4_u0_n123 ) , .A2( u0_u4_u0_n158 ) );
  AND2_X1 u0_u4_u0_U60 (.A2( u0_u4_X_3 ) , .A1( u0_u4_X_6 ) , .ZN( u0_u4_u0_n102 ) );
  AND2_X1 u0_u4_u0_U61 (.A1( u0_u4_X_6 ) , .A2( u0_u4_u0_n162 ) , .ZN( u0_u4_u0_n93 ) );
  INV_X1 u0_u4_u0_U62 (.A( u0_u4_X_4 ) , .ZN( u0_u4_u0_n159 ) );
  INV_X1 u0_u4_u0_U63 (.A( u0_u4_X_1 ) , .ZN( u0_u4_u0_n164 ) );
  INV_X1 u0_u4_u0_U64 (.A( u0_u4_X_2 ) , .ZN( u0_u4_u0_n163 ) );
  INV_X1 u0_u4_u0_U65 (.A( u0_u4_X_3 ) , .ZN( u0_u4_u0_n162 ) );
  INV_X1 u0_u4_u0_U66 (.A( u0_u4_u0_n126 ) , .ZN( u0_u4_u0_n168 ) );
  AOI211_X1 u0_u4_u0_U67 (.B( u0_u4_u0_n133 ) , .A( u0_u4_u0_n134 ) , .C2( u0_u4_u0_n135 ) , .C1( u0_u4_u0_n136 ) , .ZN( u0_u4_u0_n137 ) );
  OR4_X1 u0_u4_u0_U68 (.ZN( u0_out4_17 ) , .A4( u0_u4_u0_n122 ) , .A2( u0_u4_u0_n123 ) , .A1( u0_u4_u0_n124 ) , .A3( u0_u4_u0_n170 ) );
  AOI21_X1 u0_u4_u0_U69 (.B2( u0_u4_u0_n107 ) , .ZN( u0_u4_u0_n124 ) , .B1( u0_u4_u0_n128 ) , .A( u0_u4_u0_n161 ) );
  OAI21_X1 u0_u4_u0_U7 (.B1( u0_u4_u0_n150 ) , .B2( u0_u4_u0_n158 ) , .A( u0_u4_u0_n172 ) , .ZN( u0_u4_u0_n89 ) );
  INV_X1 u0_u4_u0_U70 (.A( u0_u4_u0_n111 ) , .ZN( u0_u4_u0_n170 ) );
  OR4_X1 u0_u4_u0_U71 (.ZN( u0_out4_31 ) , .A4( u0_u4_u0_n155 ) , .A2( u0_u4_u0_n156 ) , .A1( u0_u4_u0_n157 ) , .A3( u0_u4_u0_n173 ) );
  AOI21_X1 u0_u4_u0_U72 (.A( u0_u4_u0_n138 ) , .B2( u0_u4_u0_n139 ) , .B1( u0_u4_u0_n140 ) , .ZN( u0_u4_u0_n157 ) );
  AOI21_X1 u0_u4_u0_U73 (.B2( u0_u4_u0_n141 ) , .B1( u0_u4_u0_n142 ) , .ZN( u0_u4_u0_n156 ) , .A( u0_u4_u0_n161 ) );
  INV_X1 u0_u4_u0_U74 (.ZN( u0_u4_u0_n174 ) , .A( u0_u4_u0_n89 ) );
  AOI211_X1 u0_u4_u0_U75 (.B( u0_u4_u0_n104 ) , .A( u0_u4_u0_n105 ) , .ZN( u0_u4_u0_n106 ) , .C2( u0_u4_u0_n113 ) , .C1( u0_u4_u0_n160 ) );
  NOR2_X1 u0_u4_u0_U76 (.A2( u0_u4_X_3 ) , .A1( u0_u4_X_6 ) , .ZN( u0_u4_u0_n94 ) );
  NOR2_X1 u0_u4_u0_U77 (.A1( u0_u4_u0_n163 ) , .A2( u0_u4_u0_n164 ) , .ZN( u0_u4_u0_n95 ) );
  OAI221_X1 u0_u4_u0_U78 (.C1( u0_u4_u0_n121 ) , .ZN( u0_u4_u0_n122 ) , .B2( u0_u4_u0_n127 ) , .A( u0_u4_u0_n143 ) , .B1( u0_u4_u0_n144 ) , .C2( u0_u4_u0_n147 ) );
  NOR2_X1 u0_u4_u0_U79 (.A1( u0_u4_u0_n120 ) , .ZN( u0_u4_u0_n143 ) , .A2( u0_u4_u0_n167 ) );
  AND2_X1 u0_u4_u0_U8 (.A1( u0_u4_u0_n114 ) , .A2( u0_u4_u0_n121 ) , .ZN( u0_u4_u0_n146 ) );
  AOI21_X1 u0_u4_u0_U80 (.B1( u0_u4_u0_n132 ) , .ZN( u0_u4_u0_n133 ) , .A( u0_u4_u0_n144 ) , .B2( u0_u4_u0_n166 ) );
  OAI22_X1 u0_u4_u0_U81 (.ZN( u0_u4_u0_n105 ) , .A2( u0_u4_u0_n132 ) , .B1( u0_u4_u0_n146 ) , .A1( u0_u4_u0_n147 ) , .B2( u0_u4_u0_n161 ) );
  NAND2_X1 u0_u4_u0_U82 (.ZN( u0_u4_u0_n110 ) , .A2( u0_u4_u0_n132 ) , .A1( u0_u4_u0_n145 ) );
  INV_X1 u0_u4_u0_U83 (.A( u0_u4_u0_n119 ) , .ZN( u0_u4_u0_n167 ) );
  NAND2_X1 u0_u4_u0_U84 (.A2( u0_u4_u0_n103 ) , .ZN( u0_u4_u0_n140 ) , .A1( u0_u4_u0_n94 ) );
  NAND2_X1 u0_u4_u0_U85 (.A1( u0_u4_u0_n101 ) , .ZN( u0_u4_u0_n130 ) , .A2( u0_u4_u0_n94 ) );
  NAND2_X1 u0_u4_u0_U86 (.ZN( u0_u4_u0_n108 ) , .A1( u0_u4_u0_n92 ) , .A2( u0_u4_u0_n94 ) );
  NAND2_X1 u0_u4_u0_U87 (.ZN( u0_u4_u0_n142 ) , .A1( u0_u4_u0_n94 ) , .A2( u0_u4_u0_n95 ) );
  NAND3_X1 u0_u4_u0_U88 (.ZN( u0_out4_23 ) , .A3( u0_u4_u0_n137 ) , .A1( u0_u4_u0_n168 ) , .A2( u0_u4_u0_n171 ) );
  NAND3_X1 u0_u4_u0_U89 (.A3( u0_u4_u0_n127 ) , .A2( u0_u4_u0_n128 ) , .ZN( u0_u4_u0_n135 ) , .A1( u0_u4_u0_n150 ) );
  AND2_X1 u0_u4_u0_U9 (.A1( u0_u4_u0_n131 ) , .ZN( u0_u4_u0_n141 ) , .A2( u0_u4_u0_n150 ) );
  NAND3_X1 u0_u4_u0_U90 (.ZN( u0_u4_u0_n117 ) , .A3( u0_u4_u0_n132 ) , .A2( u0_u4_u0_n139 ) , .A1( u0_u4_u0_n148 ) );
  NAND3_X1 u0_u4_u0_U91 (.ZN( u0_u4_u0_n109 ) , .A2( u0_u4_u0_n114 ) , .A3( u0_u4_u0_n140 ) , .A1( u0_u4_u0_n149 ) );
  NAND3_X1 u0_u4_u0_U92 (.ZN( u0_out4_9 ) , .A3( u0_u4_u0_n106 ) , .A2( u0_u4_u0_n171 ) , .A1( u0_u4_u0_n174 ) );
  NAND3_X1 u0_u4_u0_U93 (.A2( u0_u4_u0_n128 ) , .A1( u0_u4_u0_n132 ) , .A3( u0_u4_u0_n146 ) , .ZN( u0_u4_u0_n97 ) );
  OAI21_X1 u0_u4_u7_U10 (.A( u0_u4_u7_n161 ) , .B1( u0_u4_u7_n168 ) , .B2( u0_u4_u7_n173 ) , .ZN( u0_u4_u7_n91 ) );
  AOI211_X1 u0_u4_u7_U11 (.A( u0_u4_u7_n117 ) , .ZN( u0_u4_u7_n118 ) , .C2( u0_u4_u7_n126 ) , .C1( u0_u4_u7_n177 ) , .B( u0_u4_u7_n180 ) );
  OAI22_X1 u0_u4_u7_U12 (.B1( u0_u4_u7_n115 ) , .ZN( u0_u4_u7_n117 ) , .A2( u0_u4_u7_n133 ) , .A1( u0_u4_u7_n137 ) , .B2( u0_u4_u7_n162 ) );
  INV_X1 u0_u4_u7_U13 (.A( u0_u4_u7_n116 ) , .ZN( u0_u4_u7_n180 ) );
  NOR3_X1 u0_u4_u7_U14 (.ZN( u0_u4_u7_n115 ) , .A3( u0_u4_u7_n145 ) , .A2( u0_u4_u7_n168 ) , .A1( u0_u4_u7_n169 ) );
  INV_X1 u0_u4_u7_U15 (.A( u0_u4_u7_n133 ) , .ZN( u0_u4_u7_n176 ) );
  NOR3_X1 u0_u4_u7_U16 (.A2( u0_u4_u7_n134 ) , .A1( u0_u4_u7_n135 ) , .ZN( u0_u4_u7_n136 ) , .A3( u0_u4_u7_n171 ) );
  NOR2_X1 u0_u4_u7_U17 (.A1( u0_u4_u7_n130 ) , .A2( u0_u4_u7_n134 ) , .ZN( u0_u4_u7_n153 ) );
  AOI21_X1 u0_u4_u7_U18 (.ZN( u0_u4_u7_n104 ) , .B2( u0_u4_u7_n112 ) , .B1( u0_u4_u7_n127 ) , .A( u0_u4_u7_n164 ) );
  AOI21_X1 u0_u4_u7_U19 (.ZN( u0_u4_u7_n106 ) , .B1( u0_u4_u7_n133 ) , .B2( u0_u4_u7_n146 ) , .A( u0_u4_u7_n162 ) );
  AOI21_X1 u0_u4_u7_U20 (.A( u0_u4_u7_n101 ) , .ZN( u0_u4_u7_n107 ) , .B2( u0_u4_u7_n128 ) , .B1( u0_u4_u7_n175 ) );
  INV_X1 u0_u4_u7_U21 (.A( u0_u4_u7_n101 ) , .ZN( u0_u4_u7_n165 ) );
  NOR2_X1 u0_u4_u7_U22 (.ZN( u0_u4_u7_n111 ) , .A2( u0_u4_u7_n134 ) , .A1( u0_u4_u7_n169 ) );
  INV_X1 u0_u4_u7_U23 (.A( u0_u4_u7_n138 ) , .ZN( u0_u4_u7_n171 ) );
  INV_X1 u0_u4_u7_U24 (.A( u0_u4_u7_n131 ) , .ZN( u0_u4_u7_n177 ) );
  INV_X1 u0_u4_u7_U25 (.A( u0_u4_u7_n110 ) , .ZN( u0_u4_u7_n174 ) );
  NAND2_X1 u0_u4_u7_U26 (.A1( u0_u4_u7_n129 ) , .A2( u0_u4_u7_n132 ) , .ZN( u0_u4_u7_n149 ) );
  NAND2_X1 u0_u4_u7_U27 (.A1( u0_u4_u7_n113 ) , .A2( u0_u4_u7_n124 ) , .ZN( u0_u4_u7_n130 ) );
  INV_X1 u0_u4_u7_U28 (.A( u0_u4_u7_n112 ) , .ZN( u0_u4_u7_n173 ) );
  INV_X1 u0_u4_u7_U29 (.A( u0_u4_u7_n128 ) , .ZN( u0_u4_u7_n168 ) );
  OAI21_X1 u0_u4_u7_U3 (.ZN( u0_u4_u7_n159 ) , .A( u0_u4_u7_n165 ) , .B2( u0_u4_u7_n171 ) , .B1( u0_u4_u7_n174 ) );
  INV_X1 u0_u4_u7_U30 (.A( u0_u4_u7_n148 ) , .ZN( u0_u4_u7_n169 ) );
  INV_X1 u0_u4_u7_U31 (.A( u0_u4_u7_n127 ) , .ZN( u0_u4_u7_n179 ) );
  NOR2_X1 u0_u4_u7_U32 (.ZN( u0_u4_u7_n101 ) , .A2( u0_u4_u7_n150 ) , .A1( u0_u4_u7_n156 ) );
  AOI211_X1 u0_u4_u7_U33 (.B( u0_u4_u7_n139 ) , .A( u0_u4_u7_n140 ) , .C2( u0_u4_u7_n141 ) , .ZN( u0_u4_u7_n142 ) , .C1( u0_u4_u7_n156 ) );
  AOI21_X1 u0_u4_u7_U34 (.A( u0_u4_u7_n137 ) , .B1( u0_u4_u7_n138 ) , .ZN( u0_u4_u7_n139 ) , .B2( u0_u4_u7_n146 ) );
  NAND4_X1 u0_u4_u7_U35 (.A3( u0_u4_u7_n127 ) , .A2( u0_u4_u7_n128 ) , .A1( u0_u4_u7_n129 ) , .ZN( u0_u4_u7_n141 ) , .A4( u0_u4_u7_n147 ) );
  OAI22_X1 u0_u4_u7_U36 (.B1( u0_u4_u7_n136 ) , .ZN( u0_u4_u7_n140 ) , .A1( u0_u4_u7_n153 ) , .B2( u0_u4_u7_n162 ) , .A2( u0_u4_u7_n164 ) );
  INV_X1 u0_u4_u7_U37 (.A( u0_u4_u7_n125 ) , .ZN( u0_u4_u7_n161 ) );
  AOI21_X1 u0_u4_u7_U38 (.ZN( u0_u4_u7_n123 ) , .B1( u0_u4_u7_n165 ) , .B2( u0_u4_u7_n177 ) , .A( u0_u4_u7_n97 ) );
  AOI21_X1 u0_u4_u7_U39 (.B2( u0_u4_u7_n113 ) , .B1( u0_u4_u7_n124 ) , .A( u0_u4_u7_n125 ) , .ZN( u0_u4_u7_n97 ) );
  INV_X1 u0_u4_u7_U4 (.A( u0_u4_u7_n149 ) , .ZN( u0_u4_u7_n175 ) );
  INV_X1 u0_u4_u7_U40 (.A( u0_u4_u7_n152 ) , .ZN( u0_u4_u7_n162 ) );
  AOI22_X1 u0_u4_u7_U41 (.A2( u0_u4_u7_n114 ) , .ZN( u0_u4_u7_n119 ) , .B1( u0_u4_u7_n130 ) , .A1( u0_u4_u7_n156 ) , .B2( u0_u4_u7_n165 ) );
  NAND2_X1 u0_u4_u7_U42 (.A2( u0_u4_u7_n112 ) , .ZN( u0_u4_u7_n114 ) , .A1( u0_u4_u7_n175 ) );
  NOR2_X1 u0_u4_u7_U43 (.ZN( u0_u4_u7_n137 ) , .A1( u0_u4_u7_n150 ) , .A2( u0_u4_u7_n161 ) );
  AND2_X1 u0_u4_u7_U44 (.ZN( u0_u4_u7_n145 ) , .A2( u0_u4_u7_n98 ) , .A1( u0_u4_u7_n99 ) );
  AOI21_X1 u0_u4_u7_U45 (.ZN( u0_u4_u7_n105 ) , .B2( u0_u4_u7_n110 ) , .A( u0_u4_u7_n125 ) , .B1( u0_u4_u7_n147 ) );
  NAND2_X1 u0_u4_u7_U46 (.ZN( u0_u4_u7_n146 ) , .A1( u0_u4_u7_n95 ) , .A2( u0_u4_u7_n98 ) );
  NAND2_X1 u0_u4_u7_U47 (.A2( u0_u4_u7_n103 ) , .ZN( u0_u4_u7_n147 ) , .A1( u0_u4_u7_n93 ) );
  NAND2_X1 u0_u4_u7_U48 (.A1( u0_u4_u7_n103 ) , .ZN( u0_u4_u7_n127 ) , .A2( u0_u4_u7_n99 ) );
  NAND2_X1 u0_u4_u7_U49 (.A2( u0_u4_u7_n102 ) , .A1( u0_u4_u7_n103 ) , .ZN( u0_u4_u7_n133 ) );
  INV_X1 u0_u4_u7_U5 (.A( u0_u4_u7_n154 ) , .ZN( u0_u4_u7_n178 ) );
  OR2_X1 u0_u4_u7_U50 (.ZN( u0_u4_u7_n126 ) , .A2( u0_u4_u7_n152 ) , .A1( u0_u4_u7_n156 ) );
  NAND2_X1 u0_u4_u7_U51 (.ZN( u0_u4_u7_n112 ) , .A2( u0_u4_u7_n96 ) , .A1( u0_u4_u7_n99 ) );
  NAND2_X1 u0_u4_u7_U52 (.A2( u0_u4_u7_n102 ) , .ZN( u0_u4_u7_n128 ) , .A1( u0_u4_u7_n98 ) );
  NAND2_X1 u0_u4_u7_U53 (.A1( u0_u4_u7_n100 ) , .ZN( u0_u4_u7_n113 ) , .A2( u0_u4_u7_n93 ) );
  NAND2_X1 u0_u4_u7_U54 (.ZN( u0_u4_u7_n110 ) , .A1( u0_u4_u7_n95 ) , .A2( u0_u4_u7_n96 ) );
  INV_X1 u0_u4_u7_U55 (.A( u0_u4_u7_n150 ) , .ZN( u0_u4_u7_n164 ) );
  AND2_X1 u0_u4_u7_U56 (.ZN( u0_u4_u7_n134 ) , .A1( u0_u4_u7_n93 ) , .A2( u0_u4_u7_n98 ) );
  NAND2_X1 u0_u4_u7_U57 (.A2( u0_u4_u7_n102 ) , .ZN( u0_u4_u7_n124 ) , .A1( u0_u4_u7_n96 ) );
  NAND2_X1 u0_u4_u7_U58 (.A1( u0_u4_u7_n100 ) , .A2( u0_u4_u7_n102 ) , .ZN( u0_u4_u7_n129 ) );
  NAND2_X1 u0_u4_u7_U59 (.A2( u0_u4_u7_n103 ) , .ZN( u0_u4_u7_n131 ) , .A1( u0_u4_u7_n95 ) );
  AOI211_X1 u0_u4_u7_U6 (.ZN( u0_u4_u7_n116 ) , .A( u0_u4_u7_n155 ) , .C1( u0_u4_u7_n161 ) , .C2( u0_u4_u7_n171 ) , .B( u0_u4_u7_n94 ) );
  NAND2_X1 u0_u4_u7_U60 (.A1( u0_u4_u7_n100 ) , .ZN( u0_u4_u7_n138 ) , .A2( u0_u4_u7_n99 ) );
  NAND2_X1 u0_u4_u7_U61 (.ZN( u0_u4_u7_n132 ) , .A1( u0_u4_u7_n93 ) , .A2( u0_u4_u7_n96 ) );
  NAND2_X1 u0_u4_u7_U62 (.A1( u0_u4_u7_n100 ) , .ZN( u0_u4_u7_n148 ) , .A2( u0_u4_u7_n95 ) );
  AOI211_X1 u0_u4_u7_U63 (.B( u0_u4_u7_n154 ) , .A( u0_u4_u7_n155 ) , .C1( u0_u4_u7_n156 ) , .ZN( u0_u4_u7_n157 ) , .C2( u0_u4_u7_n172 ) );
  INV_X1 u0_u4_u7_U64 (.A( u0_u4_u7_n153 ) , .ZN( u0_u4_u7_n172 ) );
  NOR2_X1 u0_u4_u7_U65 (.A2( u0_u4_X_47 ) , .ZN( u0_u4_u7_n150 ) , .A1( u0_u4_u7_n163 ) );
  NOR2_X1 u0_u4_u7_U66 (.A2( u0_u4_X_43 ) , .A1( u0_u4_X_44 ) , .ZN( u0_u4_u7_n103 ) );
  NOR2_X1 u0_u4_u7_U67 (.A2( u0_u4_X_48 ) , .A1( u0_u4_u7_n166 ) , .ZN( u0_u4_u7_n95 ) );
  NOR2_X1 u0_u4_u7_U68 (.A2( u0_u4_X_45 ) , .A1( u0_u4_X_48 ) , .ZN( u0_u4_u7_n99 ) );
  NOR2_X1 u0_u4_u7_U69 (.A2( u0_u4_X_44 ) , .A1( u0_u4_u7_n167 ) , .ZN( u0_u4_u7_n98 ) );
  OAI222_X1 u0_u4_u7_U7 (.C2( u0_u4_u7_n101 ) , .B2( u0_u4_u7_n111 ) , .A1( u0_u4_u7_n113 ) , .C1( u0_u4_u7_n146 ) , .A2( u0_u4_u7_n162 ) , .B1( u0_u4_u7_n164 ) , .ZN( u0_u4_u7_n94 ) );
  NOR2_X1 u0_u4_u7_U70 (.A2( u0_u4_X_46 ) , .A1( u0_u4_X_47 ) , .ZN( u0_u4_u7_n152 ) );
  NAND2_X1 u0_u4_u7_U71 (.A2( u0_u4_X_46 ) , .A1( u0_u4_X_47 ) , .ZN( u0_u4_u7_n125 ) );
  AND2_X1 u0_u4_u7_U72 (.A1( u0_u4_X_47 ) , .ZN( u0_u4_u7_n156 ) , .A2( u0_u4_u7_n163 ) );
  AND2_X1 u0_u4_u7_U73 (.A2( u0_u4_X_45 ) , .A1( u0_u4_X_48 ) , .ZN( u0_u4_u7_n102 ) );
  AND2_X1 u0_u4_u7_U74 (.A2( u0_u4_X_43 ) , .A1( u0_u4_X_44 ) , .ZN( u0_u4_u7_n96 ) );
  AND2_X1 u0_u4_u7_U75 (.A1( u0_u4_X_44 ) , .ZN( u0_u4_u7_n100 ) , .A2( u0_u4_u7_n167 ) );
  AND2_X1 u0_u4_u7_U76 (.A1( u0_u4_X_48 ) , .A2( u0_u4_u7_n166 ) , .ZN( u0_u4_u7_n93 ) );
  INV_X1 u0_u4_u7_U77 (.A( u0_u4_X_46 ) , .ZN( u0_u4_u7_n163 ) );
  INV_X1 u0_u4_u7_U78 (.A( u0_u4_X_43 ) , .ZN( u0_u4_u7_n167 ) );
  INV_X1 u0_u4_u7_U79 (.A( u0_u4_X_45 ) , .ZN( u0_u4_u7_n166 ) );
  OAI221_X1 u0_u4_u7_U8 (.C1( u0_u4_u7_n101 ) , .C2( u0_u4_u7_n147 ) , .ZN( u0_u4_u7_n155 ) , .B2( u0_u4_u7_n162 ) , .A( u0_u4_u7_n91 ) , .B1( u0_u4_u7_n92 ) );
  NAND4_X1 u0_u4_u7_U80 (.ZN( u0_out4_5 ) , .A4( u0_u4_u7_n108 ) , .A3( u0_u4_u7_n109 ) , .A1( u0_u4_u7_n116 ) , .A2( u0_u4_u7_n123 ) );
  AOI22_X1 u0_u4_u7_U81 (.ZN( u0_u4_u7_n109 ) , .A2( u0_u4_u7_n126 ) , .B2( u0_u4_u7_n145 ) , .B1( u0_u4_u7_n156 ) , .A1( u0_u4_u7_n171 ) );
  NOR4_X1 u0_u4_u7_U82 (.A4( u0_u4_u7_n104 ) , .A3( u0_u4_u7_n105 ) , .A2( u0_u4_u7_n106 ) , .A1( u0_u4_u7_n107 ) , .ZN( u0_u4_u7_n108 ) );
  NAND4_X1 u0_u4_u7_U83 (.ZN( u0_out4_27 ) , .A4( u0_u4_u7_n118 ) , .A3( u0_u4_u7_n119 ) , .A2( u0_u4_u7_n120 ) , .A1( u0_u4_u7_n121 ) );
  OAI21_X1 u0_u4_u7_U84 (.ZN( u0_u4_u7_n121 ) , .B2( u0_u4_u7_n145 ) , .A( u0_u4_u7_n150 ) , .B1( u0_u4_u7_n174 ) );
  OAI21_X1 u0_u4_u7_U85 (.ZN( u0_u4_u7_n120 ) , .A( u0_u4_u7_n161 ) , .B2( u0_u4_u7_n170 ) , .B1( u0_u4_u7_n179 ) );
  NAND4_X1 u0_u4_u7_U86 (.ZN( u0_out4_21 ) , .A4( u0_u4_u7_n157 ) , .A3( u0_u4_u7_n158 ) , .A2( u0_u4_u7_n159 ) , .A1( u0_u4_u7_n160 ) );
  OAI21_X1 u0_u4_u7_U87 (.B1( u0_u4_u7_n145 ) , .ZN( u0_u4_u7_n160 ) , .A( u0_u4_u7_n161 ) , .B2( u0_u4_u7_n177 ) );
  AOI22_X1 u0_u4_u7_U88 (.B2( u0_u4_u7_n149 ) , .B1( u0_u4_u7_n150 ) , .A2( u0_u4_u7_n151 ) , .A1( u0_u4_u7_n152 ) , .ZN( u0_u4_u7_n158 ) );
  NAND4_X1 u0_u4_u7_U89 (.ZN( u0_out4_15 ) , .A4( u0_u4_u7_n142 ) , .A3( u0_u4_u7_n143 ) , .A2( u0_u4_u7_n144 ) , .A1( u0_u4_u7_n178 ) );
  AND3_X1 u0_u4_u7_U9 (.A3( u0_u4_u7_n110 ) , .A2( u0_u4_u7_n127 ) , .A1( u0_u4_u7_n132 ) , .ZN( u0_u4_u7_n92 ) );
  OR2_X1 u0_u4_u7_U90 (.A2( u0_u4_u7_n125 ) , .A1( u0_u4_u7_n129 ) , .ZN( u0_u4_u7_n144 ) );
  AOI22_X1 u0_u4_u7_U91 (.A2( u0_u4_u7_n126 ) , .ZN( u0_u4_u7_n143 ) , .B2( u0_u4_u7_n165 ) , .B1( u0_u4_u7_n173 ) , .A1( u0_u4_u7_n174 ) );
  OAI211_X1 u0_u4_u7_U92 (.B( u0_u4_u7_n122 ) , .A( u0_u4_u7_n123 ) , .C2( u0_u4_u7_n124 ) , .ZN( u0_u4_u7_n154 ) , .C1( u0_u4_u7_n162 ) );
  AOI222_X1 u0_u4_u7_U93 (.ZN( u0_u4_u7_n122 ) , .C2( u0_u4_u7_n126 ) , .C1( u0_u4_u7_n145 ) , .B1( u0_u4_u7_n161 ) , .A2( u0_u4_u7_n165 ) , .B2( u0_u4_u7_n170 ) , .A1( u0_u4_u7_n176 ) );
  INV_X1 u0_u4_u7_U94 (.A( u0_u4_u7_n111 ) , .ZN( u0_u4_u7_n170 ) );
  NAND3_X1 u0_u4_u7_U95 (.A3( u0_u4_u7_n146 ) , .A2( u0_u4_u7_n147 ) , .A1( u0_u4_u7_n148 ) , .ZN( u0_u4_u7_n151 ) );
  NAND3_X1 u0_u4_u7_U96 (.A3( u0_u4_u7_n131 ) , .A2( u0_u4_u7_n132 ) , .A1( u0_u4_u7_n133 ) , .ZN( u0_u4_u7_n135 ) );
  XOR2_X1 u0_u7_U13 (.B( u0_K8_42 ) , .A( u0_R6_29 ) , .Z( u0_u7_X_42 ) );
  XOR2_X1 u0_u7_U14 (.B( u0_K8_41 ) , .A( u0_R6_28 ) , .Z( u0_u7_X_41 ) );
  XOR2_X1 u0_u7_U15 (.B( u0_K8_40 ) , .A( u0_R6_27 ) , .Z( u0_u7_X_40 ) );
  XOR2_X1 u0_u7_U17 (.B( u0_K8_39 ) , .A( u0_R6_26 ) , .Z( u0_u7_X_39 ) );
  XOR2_X1 u0_u7_U18 (.B( u0_K8_38 ) , .A( u0_R6_25 ) , .Z( u0_u7_X_38 ) );
  XOR2_X1 u0_u7_U19 (.B( u0_K8_37 ) , .A( u0_R6_24 ) , .Z( u0_u7_X_37 ) );
  XOR2_X1 u0_u7_U20 (.B( u0_K8_36 ) , .A( u0_R6_25 ) , .Z( u0_u7_X_36 ) );
  XOR2_X1 u0_u7_U21 (.B( u0_K8_35 ) , .A( u0_R6_24 ) , .Z( u0_u7_X_35 ) );
  XOR2_X1 u0_u7_U22 (.B( u0_K8_34 ) , .A( u0_R6_23 ) , .Z( u0_u7_X_34 ) );
  XOR2_X1 u0_u7_U23 (.B( u0_K8_33 ) , .A( u0_R6_22 ) , .Z( u0_u7_X_33 ) );
  XOR2_X1 u0_u7_U24 (.B( u0_K8_32 ) , .A( u0_R6_21 ) , .Z( u0_u7_X_32 ) );
  XOR2_X1 u0_u7_U25 (.B( u0_K8_31 ) , .A( u0_R6_20 ) , .Z( u0_u7_X_31 ) );
  XOR2_X1 u0_u7_U26 (.B( u0_K8_30 ) , .A( u0_R6_21 ) , .Z( u0_u7_X_30 ) );
  XOR2_X1 u0_u7_U28 (.B( u0_K8_29 ) , .A( u0_R6_20 ) , .Z( u0_u7_X_29 ) );
  XOR2_X1 u0_u7_U29 (.B( u0_K8_28 ) , .A( u0_R6_19 ) , .Z( u0_u7_X_28 ) );
  XOR2_X1 u0_u7_U30 (.B( u0_K8_27 ) , .A( u0_R6_18 ) , .Z( u0_u7_X_27 ) );
  XOR2_X1 u0_u7_U31 (.B( u0_K8_26 ) , .A( u0_R6_17 ) , .Z( u0_u7_X_26 ) );
  XOR2_X1 u0_u7_U32 (.B( u0_K8_25 ) , .A( u0_R6_16 ) , .Z( u0_u7_X_25 ) );
  OAI22_X1 u0_u7_u4_U10 (.B2( u0_u7_u4_n135 ) , .ZN( u0_u7_u4_n137 ) , .B1( u0_u7_u4_n153 ) , .A1( u0_u7_u4_n155 ) , .A2( u0_u7_u4_n171 ) );
  AND3_X1 u0_u7_u4_U11 (.A2( u0_u7_u4_n134 ) , .ZN( u0_u7_u4_n135 ) , .A3( u0_u7_u4_n145 ) , .A1( u0_u7_u4_n157 ) );
  OR3_X1 u0_u7_u4_U12 (.A3( u0_u7_u4_n114 ) , .A2( u0_u7_u4_n115 ) , .A1( u0_u7_u4_n116 ) , .ZN( u0_u7_u4_n136 ) );
  AOI21_X1 u0_u7_u4_U13 (.A( u0_u7_u4_n113 ) , .ZN( u0_u7_u4_n116 ) , .B2( u0_u7_u4_n173 ) , .B1( u0_u7_u4_n174 ) );
  AOI21_X1 u0_u7_u4_U14 (.ZN( u0_u7_u4_n115 ) , .B2( u0_u7_u4_n145 ) , .B1( u0_u7_u4_n146 ) , .A( u0_u7_u4_n156 ) );
  OAI22_X1 u0_u7_u4_U15 (.ZN( u0_u7_u4_n114 ) , .A2( u0_u7_u4_n121 ) , .B1( u0_u7_u4_n160 ) , .B2( u0_u7_u4_n170 ) , .A1( u0_u7_u4_n171 ) );
  NAND2_X1 u0_u7_u4_U16 (.ZN( u0_u7_u4_n132 ) , .A2( u0_u7_u4_n170 ) , .A1( u0_u7_u4_n173 ) );
  AOI21_X1 u0_u7_u4_U17 (.B2( u0_u7_u4_n160 ) , .B1( u0_u7_u4_n161 ) , .ZN( u0_u7_u4_n162 ) , .A( u0_u7_u4_n170 ) );
  AOI21_X1 u0_u7_u4_U18 (.ZN( u0_u7_u4_n107 ) , .B2( u0_u7_u4_n143 ) , .A( u0_u7_u4_n174 ) , .B1( u0_u7_u4_n184 ) );
  AOI21_X1 u0_u7_u4_U19 (.B2( u0_u7_u4_n158 ) , .B1( u0_u7_u4_n159 ) , .ZN( u0_u7_u4_n163 ) , .A( u0_u7_u4_n174 ) );
  AOI21_X1 u0_u7_u4_U20 (.A( u0_u7_u4_n153 ) , .B2( u0_u7_u4_n154 ) , .B1( u0_u7_u4_n155 ) , .ZN( u0_u7_u4_n165 ) );
  AOI21_X1 u0_u7_u4_U21 (.A( u0_u7_u4_n156 ) , .B2( u0_u7_u4_n157 ) , .ZN( u0_u7_u4_n164 ) , .B1( u0_u7_u4_n184 ) );
  INV_X1 u0_u7_u4_U22 (.A( u0_u7_u4_n138 ) , .ZN( u0_u7_u4_n170 ) );
  AND2_X1 u0_u7_u4_U23 (.A2( u0_u7_u4_n120 ) , .ZN( u0_u7_u4_n155 ) , .A1( u0_u7_u4_n160 ) );
  INV_X1 u0_u7_u4_U24 (.A( u0_u7_u4_n156 ) , .ZN( u0_u7_u4_n175 ) );
  NAND2_X1 u0_u7_u4_U25 (.A2( u0_u7_u4_n118 ) , .ZN( u0_u7_u4_n131 ) , .A1( u0_u7_u4_n147 ) );
  NAND2_X1 u0_u7_u4_U26 (.A1( u0_u7_u4_n119 ) , .A2( u0_u7_u4_n120 ) , .ZN( u0_u7_u4_n130 ) );
  NAND2_X1 u0_u7_u4_U27 (.ZN( u0_u7_u4_n117 ) , .A2( u0_u7_u4_n118 ) , .A1( u0_u7_u4_n148 ) );
  NAND2_X1 u0_u7_u4_U28 (.ZN( u0_u7_u4_n129 ) , .A1( u0_u7_u4_n134 ) , .A2( u0_u7_u4_n148 ) );
  AND3_X1 u0_u7_u4_U29 (.A1( u0_u7_u4_n119 ) , .A2( u0_u7_u4_n143 ) , .A3( u0_u7_u4_n154 ) , .ZN( u0_u7_u4_n161 ) );
  NOR2_X1 u0_u7_u4_U3 (.ZN( u0_u7_u4_n121 ) , .A1( u0_u7_u4_n181 ) , .A2( u0_u7_u4_n182 ) );
  AND2_X1 u0_u7_u4_U30 (.A1( u0_u7_u4_n145 ) , .A2( u0_u7_u4_n147 ) , .ZN( u0_u7_u4_n159 ) );
  INV_X1 u0_u7_u4_U31 (.A( u0_u7_u4_n158 ) , .ZN( u0_u7_u4_n182 ) );
  INV_X1 u0_u7_u4_U32 (.ZN( u0_u7_u4_n181 ) , .A( u0_u7_u4_n96 ) );
  INV_X1 u0_u7_u4_U33 (.A( u0_u7_u4_n144 ) , .ZN( u0_u7_u4_n179 ) );
  INV_X1 u0_u7_u4_U34 (.A( u0_u7_u4_n157 ) , .ZN( u0_u7_u4_n178 ) );
  NAND2_X1 u0_u7_u4_U35 (.A2( u0_u7_u4_n154 ) , .A1( u0_u7_u4_n96 ) , .ZN( u0_u7_u4_n97 ) );
  INV_X1 u0_u7_u4_U36 (.ZN( u0_u7_u4_n186 ) , .A( u0_u7_u4_n95 ) );
  OAI221_X1 u0_u7_u4_U37 (.C1( u0_u7_u4_n134 ) , .B1( u0_u7_u4_n158 ) , .B2( u0_u7_u4_n171 ) , .C2( u0_u7_u4_n173 ) , .A( u0_u7_u4_n94 ) , .ZN( u0_u7_u4_n95 ) );
  AOI222_X1 u0_u7_u4_U38 (.B2( u0_u7_u4_n132 ) , .A1( u0_u7_u4_n138 ) , .C2( u0_u7_u4_n175 ) , .A2( u0_u7_u4_n179 ) , .C1( u0_u7_u4_n181 ) , .B1( u0_u7_u4_n185 ) , .ZN( u0_u7_u4_n94 ) );
  INV_X1 u0_u7_u4_U39 (.A( u0_u7_u4_n113 ) , .ZN( u0_u7_u4_n185 ) );
  INV_X1 u0_u7_u4_U4 (.A( u0_u7_u4_n117 ) , .ZN( u0_u7_u4_n184 ) );
  INV_X1 u0_u7_u4_U40 (.A( u0_u7_u4_n143 ) , .ZN( u0_u7_u4_n183 ) );
  NOR2_X1 u0_u7_u4_U41 (.ZN( u0_u7_u4_n138 ) , .A1( u0_u7_u4_n168 ) , .A2( u0_u7_u4_n169 ) );
  NOR2_X1 u0_u7_u4_U42 (.A1( u0_u7_u4_n150 ) , .A2( u0_u7_u4_n152 ) , .ZN( u0_u7_u4_n153 ) );
  NOR2_X1 u0_u7_u4_U43 (.A2( u0_u7_u4_n128 ) , .A1( u0_u7_u4_n138 ) , .ZN( u0_u7_u4_n156 ) );
  AOI22_X1 u0_u7_u4_U44 (.B2( u0_u7_u4_n122 ) , .A1( u0_u7_u4_n123 ) , .ZN( u0_u7_u4_n124 ) , .B1( u0_u7_u4_n128 ) , .A2( u0_u7_u4_n172 ) );
  NAND2_X1 u0_u7_u4_U45 (.A2( u0_u7_u4_n120 ) , .ZN( u0_u7_u4_n123 ) , .A1( u0_u7_u4_n161 ) );
  INV_X1 u0_u7_u4_U46 (.A( u0_u7_u4_n153 ) , .ZN( u0_u7_u4_n172 ) );
  AOI22_X1 u0_u7_u4_U47 (.B2( u0_u7_u4_n132 ) , .A2( u0_u7_u4_n133 ) , .ZN( u0_u7_u4_n140 ) , .A1( u0_u7_u4_n150 ) , .B1( u0_u7_u4_n179 ) );
  NAND2_X1 u0_u7_u4_U48 (.ZN( u0_u7_u4_n133 ) , .A2( u0_u7_u4_n146 ) , .A1( u0_u7_u4_n154 ) );
  NAND2_X1 u0_u7_u4_U49 (.A1( u0_u7_u4_n103 ) , .ZN( u0_u7_u4_n154 ) , .A2( u0_u7_u4_n98 ) );
  NOR4_X1 u0_u7_u4_U5 (.A4( u0_u7_u4_n106 ) , .A3( u0_u7_u4_n107 ) , .A2( u0_u7_u4_n108 ) , .A1( u0_u7_u4_n109 ) , .ZN( u0_u7_u4_n110 ) );
  NAND2_X1 u0_u7_u4_U50 (.A1( u0_u7_u4_n101 ) , .ZN( u0_u7_u4_n158 ) , .A2( u0_u7_u4_n99 ) );
  AOI21_X1 u0_u7_u4_U51 (.ZN( u0_u7_u4_n127 ) , .A( u0_u7_u4_n136 ) , .B2( u0_u7_u4_n150 ) , .B1( u0_u7_u4_n180 ) );
  INV_X1 u0_u7_u4_U52 (.A( u0_u7_u4_n160 ) , .ZN( u0_u7_u4_n180 ) );
  NAND2_X1 u0_u7_u4_U53 (.A2( u0_u7_u4_n104 ) , .A1( u0_u7_u4_n105 ) , .ZN( u0_u7_u4_n146 ) );
  NAND2_X1 u0_u7_u4_U54 (.A2( u0_u7_u4_n101 ) , .A1( u0_u7_u4_n102 ) , .ZN( u0_u7_u4_n160 ) );
  NAND2_X1 u0_u7_u4_U55 (.ZN( u0_u7_u4_n134 ) , .A1( u0_u7_u4_n98 ) , .A2( u0_u7_u4_n99 ) );
  NAND2_X1 u0_u7_u4_U56 (.A1( u0_u7_u4_n103 ) , .A2( u0_u7_u4_n104 ) , .ZN( u0_u7_u4_n143 ) );
  NAND2_X1 u0_u7_u4_U57 (.A2( u0_u7_u4_n105 ) , .ZN( u0_u7_u4_n145 ) , .A1( u0_u7_u4_n98 ) );
  NAND2_X1 u0_u7_u4_U58 (.A1( u0_u7_u4_n100 ) , .A2( u0_u7_u4_n105 ) , .ZN( u0_u7_u4_n120 ) );
  NAND2_X1 u0_u7_u4_U59 (.A1( u0_u7_u4_n102 ) , .A2( u0_u7_u4_n104 ) , .ZN( u0_u7_u4_n148 ) );
  AOI21_X1 u0_u7_u4_U6 (.ZN( u0_u7_u4_n106 ) , .B2( u0_u7_u4_n146 ) , .B1( u0_u7_u4_n158 ) , .A( u0_u7_u4_n170 ) );
  NAND2_X1 u0_u7_u4_U60 (.A2( u0_u7_u4_n100 ) , .A1( u0_u7_u4_n103 ) , .ZN( u0_u7_u4_n157 ) );
  INV_X1 u0_u7_u4_U61 (.A( u0_u7_u4_n150 ) , .ZN( u0_u7_u4_n173 ) );
  INV_X1 u0_u7_u4_U62 (.A( u0_u7_u4_n152 ) , .ZN( u0_u7_u4_n171 ) );
  NAND2_X1 u0_u7_u4_U63 (.A1( u0_u7_u4_n100 ) , .ZN( u0_u7_u4_n118 ) , .A2( u0_u7_u4_n99 ) );
  NAND2_X1 u0_u7_u4_U64 (.A2( u0_u7_u4_n100 ) , .A1( u0_u7_u4_n102 ) , .ZN( u0_u7_u4_n144 ) );
  NAND2_X1 u0_u7_u4_U65 (.A2( u0_u7_u4_n101 ) , .A1( u0_u7_u4_n105 ) , .ZN( u0_u7_u4_n96 ) );
  INV_X1 u0_u7_u4_U66 (.A( u0_u7_u4_n128 ) , .ZN( u0_u7_u4_n174 ) );
  NAND2_X1 u0_u7_u4_U67 (.A2( u0_u7_u4_n102 ) , .ZN( u0_u7_u4_n119 ) , .A1( u0_u7_u4_n98 ) );
  NAND2_X1 u0_u7_u4_U68 (.A2( u0_u7_u4_n101 ) , .A1( u0_u7_u4_n103 ) , .ZN( u0_u7_u4_n147 ) );
  NAND2_X1 u0_u7_u4_U69 (.A2( u0_u7_u4_n104 ) , .ZN( u0_u7_u4_n113 ) , .A1( u0_u7_u4_n99 ) );
  AOI21_X1 u0_u7_u4_U7 (.ZN( u0_u7_u4_n108 ) , .B2( u0_u7_u4_n134 ) , .B1( u0_u7_u4_n155 ) , .A( u0_u7_u4_n156 ) );
  NOR2_X1 u0_u7_u4_U70 (.A2( u0_u7_X_28 ) , .ZN( u0_u7_u4_n150 ) , .A1( u0_u7_u4_n168 ) );
  NOR2_X1 u0_u7_u4_U71 (.A2( u0_u7_X_29 ) , .ZN( u0_u7_u4_n152 ) , .A1( u0_u7_u4_n169 ) );
  NOR2_X1 u0_u7_u4_U72 (.A2( u0_u7_X_26 ) , .ZN( u0_u7_u4_n100 ) , .A1( u0_u7_u4_n177 ) );
  NOR2_X1 u0_u7_u4_U73 (.A2( u0_u7_X_30 ) , .ZN( u0_u7_u4_n105 ) , .A1( u0_u7_u4_n176 ) );
  NOR2_X1 u0_u7_u4_U74 (.A2( u0_u7_X_28 ) , .A1( u0_u7_X_29 ) , .ZN( u0_u7_u4_n128 ) );
  NOR2_X1 u0_u7_u4_U75 (.A2( u0_u7_X_25 ) , .A1( u0_u7_X_26 ) , .ZN( u0_u7_u4_n98 ) );
  NOR2_X1 u0_u7_u4_U76 (.A2( u0_u7_X_27 ) , .A1( u0_u7_X_30 ) , .ZN( u0_u7_u4_n102 ) );
  AND2_X1 u0_u7_u4_U77 (.A2( u0_u7_X_25 ) , .A1( u0_u7_X_26 ) , .ZN( u0_u7_u4_n104 ) );
  AND2_X1 u0_u7_u4_U78 (.A1( u0_u7_X_30 ) , .A2( u0_u7_u4_n176 ) , .ZN( u0_u7_u4_n99 ) );
  AND2_X1 u0_u7_u4_U79 (.A1( u0_u7_X_26 ) , .ZN( u0_u7_u4_n101 ) , .A2( u0_u7_u4_n177 ) );
  AOI21_X1 u0_u7_u4_U8 (.ZN( u0_u7_u4_n109 ) , .A( u0_u7_u4_n153 ) , .B1( u0_u7_u4_n159 ) , .B2( u0_u7_u4_n184 ) );
  AND2_X1 u0_u7_u4_U80 (.A1( u0_u7_X_27 ) , .A2( u0_u7_X_30 ) , .ZN( u0_u7_u4_n103 ) );
  INV_X1 u0_u7_u4_U81 (.A( u0_u7_X_28 ) , .ZN( u0_u7_u4_n169 ) );
  INV_X1 u0_u7_u4_U82 (.A( u0_u7_X_29 ) , .ZN( u0_u7_u4_n168 ) );
  INV_X1 u0_u7_u4_U83 (.A( u0_u7_X_25 ) , .ZN( u0_u7_u4_n177 ) );
  INV_X1 u0_u7_u4_U84 (.A( u0_u7_X_27 ) , .ZN( u0_u7_u4_n176 ) );
  NAND4_X1 u0_u7_u4_U85 (.ZN( u0_out7_25 ) , .A4( u0_u7_u4_n139 ) , .A3( u0_u7_u4_n140 ) , .A2( u0_u7_u4_n141 ) , .A1( u0_u7_u4_n142 ) );
  OAI21_X1 u0_u7_u4_U86 (.A( u0_u7_u4_n128 ) , .B2( u0_u7_u4_n129 ) , .B1( u0_u7_u4_n130 ) , .ZN( u0_u7_u4_n142 ) );
  OAI21_X1 u0_u7_u4_U87 (.B2( u0_u7_u4_n131 ) , .ZN( u0_u7_u4_n141 ) , .A( u0_u7_u4_n175 ) , .B1( u0_u7_u4_n183 ) );
  NAND4_X1 u0_u7_u4_U88 (.ZN( u0_out7_14 ) , .A4( u0_u7_u4_n124 ) , .A3( u0_u7_u4_n125 ) , .A2( u0_u7_u4_n126 ) , .A1( u0_u7_u4_n127 ) );
  AOI22_X1 u0_u7_u4_U89 (.B2( u0_u7_u4_n117 ) , .ZN( u0_u7_u4_n126 ) , .A1( u0_u7_u4_n129 ) , .B1( u0_u7_u4_n152 ) , .A2( u0_u7_u4_n175 ) );
  AOI211_X1 u0_u7_u4_U9 (.B( u0_u7_u4_n136 ) , .A( u0_u7_u4_n137 ) , .C2( u0_u7_u4_n138 ) , .ZN( u0_u7_u4_n139 ) , .C1( u0_u7_u4_n182 ) );
  AOI22_X1 u0_u7_u4_U90 (.ZN( u0_u7_u4_n125 ) , .B2( u0_u7_u4_n131 ) , .A2( u0_u7_u4_n132 ) , .B1( u0_u7_u4_n138 ) , .A1( u0_u7_u4_n178 ) );
  NAND4_X1 u0_u7_u4_U91 (.ZN( u0_out7_8 ) , .A4( u0_u7_u4_n110 ) , .A3( u0_u7_u4_n111 ) , .A2( u0_u7_u4_n112 ) , .A1( u0_u7_u4_n186 ) );
  NAND2_X1 u0_u7_u4_U92 (.ZN( u0_u7_u4_n112 ) , .A2( u0_u7_u4_n130 ) , .A1( u0_u7_u4_n150 ) );
  AOI22_X1 u0_u7_u4_U93 (.ZN( u0_u7_u4_n111 ) , .B2( u0_u7_u4_n132 ) , .A1( u0_u7_u4_n152 ) , .B1( u0_u7_u4_n178 ) , .A2( u0_u7_u4_n97 ) );
  AOI22_X1 u0_u7_u4_U94 (.B2( u0_u7_u4_n149 ) , .B1( u0_u7_u4_n150 ) , .A2( u0_u7_u4_n151 ) , .A1( u0_u7_u4_n152 ) , .ZN( u0_u7_u4_n167 ) );
  NOR4_X1 u0_u7_u4_U95 (.A4( u0_u7_u4_n162 ) , .A3( u0_u7_u4_n163 ) , .A2( u0_u7_u4_n164 ) , .A1( u0_u7_u4_n165 ) , .ZN( u0_u7_u4_n166 ) );
  NAND3_X1 u0_u7_u4_U96 (.ZN( u0_out7_3 ) , .A3( u0_u7_u4_n166 ) , .A1( u0_u7_u4_n167 ) , .A2( u0_u7_u4_n186 ) );
  NAND3_X1 u0_u7_u4_U97 (.A3( u0_u7_u4_n146 ) , .A2( u0_u7_u4_n147 ) , .A1( u0_u7_u4_n148 ) , .ZN( u0_u7_u4_n149 ) );
  NAND3_X1 u0_u7_u4_U98 (.A3( u0_u7_u4_n143 ) , .A2( u0_u7_u4_n144 ) , .A1( u0_u7_u4_n145 ) , .ZN( u0_u7_u4_n151 ) );
  NAND3_X1 u0_u7_u4_U99 (.A3( u0_u7_u4_n121 ) , .ZN( u0_u7_u4_n122 ) , .A2( u0_u7_u4_n144 ) , .A1( u0_u7_u4_n154 ) );
  INV_X1 u0_u7_u5_U10 (.A( u0_u7_u5_n121 ) , .ZN( u0_u7_u5_n177 ) );
  NOR3_X1 u0_u7_u5_U100 (.A3( u0_u7_u5_n141 ) , .A1( u0_u7_u5_n142 ) , .ZN( u0_u7_u5_n143 ) , .A2( u0_u7_u5_n191 ) );
  NAND4_X1 u0_u7_u5_U101 (.ZN( u0_out7_4 ) , .A4( u0_u7_u5_n112 ) , .A2( u0_u7_u5_n113 ) , .A1( u0_u7_u5_n114 ) , .A3( u0_u7_u5_n195 ) );
  AOI211_X1 u0_u7_u5_U102 (.A( u0_u7_u5_n110 ) , .C1( u0_u7_u5_n111 ) , .ZN( u0_u7_u5_n112 ) , .B( u0_u7_u5_n118 ) , .C2( u0_u7_u5_n177 ) );
  AOI222_X1 u0_u7_u5_U103 (.ZN( u0_u7_u5_n113 ) , .A1( u0_u7_u5_n131 ) , .C1( u0_u7_u5_n148 ) , .B2( u0_u7_u5_n174 ) , .C2( u0_u7_u5_n178 ) , .A2( u0_u7_u5_n179 ) , .B1( u0_u7_u5_n99 ) );
  NAND3_X1 u0_u7_u5_U104 (.A2( u0_u7_u5_n154 ) , .A3( u0_u7_u5_n158 ) , .A1( u0_u7_u5_n161 ) , .ZN( u0_u7_u5_n99 ) );
  NOR2_X1 u0_u7_u5_U11 (.ZN( u0_u7_u5_n160 ) , .A2( u0_u7_u5_n173 ) , .A1( u0_u7_u5_n177 ) );
  INV_X1 u0_u7_u5_U12 (.A( u0_u7_u5_n150 ) , .ZN( u0_u7_u5_n174 ) );
  AOI21_X1 u0_u7_u5_U13 (.A( u0_u7_u5_n160 ) , .B2( u0_u7_u5_n161 ) , .ZN( u0_u7_u5_n162 ) , .B1( u0_u7_u5_n192 ) );
  INV_X1 u0_u7_u5_U14 (.A( u0_u7_u5_n159 ) , .ZN( u0_u7_u5_n192 ) );
  AOI21_X1 u0_u7_u5_U15 (.A( u0_u7_u5_n156 ) , .B2( u0_u7_u5_n157 ) , .B1( u0_u7_u5_n158 ) , .ZN( u0_u7_u5_n163 ) );
  AOI21_X1 u0_u7_u5_U16 (.B2( u0_u7_u5_n139 ) , .B1( u0_u7_u5_n140 ) , .ZN( u0_u7_u5_n141 ) , .A( u0_u7_u5_n150 ) );
  OAI21_X1 u0_u7_u5_U17 (.A( u0_u7_u5_n133 ) , .B2( u0_u7_u5_n134 ) , .B1( u0_u7_u5_n135 ) , .ZN( u0_u7_u5_n142 ) );
  OAI21_X1 u0_u7_u5_U18 (.ZN( u0_u7_u5_n133 ) , .B2( u0_u7_u5_n147 ) , .A( u0_u7_u5_n173 ) , .B1( u0_u7_u5_n188 ) );
  NAND2_X1 u0_u7_u5_U19 (.A2( u0_u7_u5_n119 ) , .A1( u0_u7_u5_n123 ) , .ZN( u0_u7_u5_n137 ) );
  INV_X1 u0_u7_u5_U20 (.A( u0_u7_u5_n155 ) , .ZN( u0_u7_u5_n194 ) );
  NAND2_X1 u0_u7_u5_U21 (.A1( u0_u7_u5_n121 ) , .ZN( u0_u7_u5_n132 ) , .A2( u0_u7_u5_n172 ) );
  NAND2_X1 u0_u7_u5_U22 (.A2( u0_u7_u5_n122 ) , .ZN( u0_u7_u5_n136 ) , .A1( u0_u7_u5_n154 ) );
  NAND2_X1 u0_u7_u5_U23 (.A2( u0_u7_u5_n119 ) , .A1( u0_u7_u5_n120 ) , .ZN( u0_u7_u5_n159 ) );
  INV_X1 u0_u7_u5_U24 (.A( u0_u7_u5_n156 ) , .ZN( u0_u7_u5_n175 ) );
  INV_X1 u0_u7_u5_U25 (.A( u0_u7_u5_n158 ) , .ZN( u0_u7_u5_n188 ) );
  INV_X1 u0_u7_u5_U26 (.A( u0_u7_u5_n152 ) , .ZN( u0_u7_u5_n179 ) );
  INV_X1 u0_u7_u5_U27 (.A( u0_u7_u5_n140 ) , .ZN( u0_u7_u5_n182 ) );
  INV_X1 u0_u7_u5_U28 (.A( u0_u7_u5_n151 ) , .ZN( u0_u7_u5_n183 ) );
  INV_X1 u0_u7_u5_U29 (.A( u0_u7_u5_n123 ) , .ZN( u0_u7_u5_n185 ) );
  NOR2_X1 u0_u7_u5_U3 (.ZN( u0_u7_u5_n134 ) , .A1( u0_u7_u5_n183 ) , .A2( u0_u7_u5_n190 ) );
  INV_X1 u0_u7_u5_U30 (.A( u0_u7_u5_n161 ) , .ZN( u0_u7_u5_n184 ) );
  INV_X1 u0_u7_u5_U31 (.A( u0_u7_u5_n139 ) , .ZN( u0_u7_u5_n189 ) );
  INV_X1 u0_u7_u5_U32 (.A( u0_u7_u5_n157 ) , .ZN( u0_u7_u5_n190 ) );
  INV_X1 u0_u7_u5_U33 (.A( u0_u7_u5_n120 ) , .ZN( u0_u7_u5_n193 ) );
  NAND2_X1 u0_u7_u5_U34 (.ZN( u0_u7_u5_n111 ) , .A1( u0_u7_u5_n140 ) , .A2( u0_u7_u5_n155 ) );
  NOR2_X1 u0_u7_u5_U35 (.ZN( u0_u7_u5_n100 ) , .A1( u0_u7_u5_n170 ) , .A2( u0_u7_u5_n180 ) );
  INV_X1 u0_u7_u5_U36 (.A( u0_u7_u5_n117 ) , .ZN( u0_u7_u5_n196 ) );
  OAI221_X1 u0_u7_u5_U37 (.A( u0_u7_u5_n116 ) , .ZN( u0_u7_u5_n117 ) , .B2( u0_u7_u5_n119 ) , .C1( u0_u7_u5_n153 ) , .C2( u0_u7_u5_n158 ) , .B1( u0_u7_u5_n172 ) );
  AOI222_X1 u0_u7_u5_U38 (.ZN( u0_u7_u5_n116 ) , .B2( u0_u7_u5_n145 ) , .C1( u0_u7_u5_n148 ) , .A2( u0_u7_u5_n174 ) , .C2( u0_u7_u5_n177 ) , .B1( u0_u7_u5_n187 ) , .A1( u0_u7_u5_n193 ) );
  INV_X1 u0_u7_u5_U39 (.A( u0_u7_u5_n115 ) , .ZN( u0_u7_u5_n187 ) );
  INV_X1 u0_u7_u5_U4 (.A( u0_u7_u5_n138 ) , .ZN( u0_u7_u5_n191 ) );
  AOI22_X1 u0_u7_u5_U40 (.B2( u0_u7_u5_n131 ) , .A2( u0_u7_u5_n146 ) , .ZN( u0_u7_u5_n169 ) , .B1( u0_u7_u5_n174 ) , .A1( u0_u7_u5_n185 ) );
  NOR2_X1 u0_u7_u5_U41 (.A1( u0_u7_u5_n146 ) , .ZN( u0_u7_u5_n150 ) , .A2( u0_u7_u5_n173 ) );
  AOI21_X1 u0_u7_u5_U42 (.A( u0_u7_u5_n118 ) , .B2( u0_u7_u5_n145 ) , .ZN( u0_u7_u5_n168 ) , .B1( u0_u7_u5_n186 ) );
  INV_X1 u0_u7_u5_U43 (.A( u0_u7_u5_n122 ) , .ZN( u0_u7_u5_n186 ) );
  NOR2_X1 u0_u7_u5_U44 (.A1( u0_u7_u5_n146 ) , .ZN( u0_u7_u5_n152 ) , .A2( u0_u7_u5_n176 ) );
  NOR2_X1 u0_u7_u5_U45 (.A1( u0_u7_u5_n115 ) , .ZN( u0_u7_u5_n118 ) , .A2( u0_u7_u5_n153 ) );
  NOR2_X1 u0_u7_u5_U46 (.A2( u0_u7_u5_n145 ) , .ZN( u0_u7_u5_n156 ) , .A1( u0_u7_u5_n174 ) );
  NOR2_X1 u0_u7_u5_U47 (.ZN( u0_u7_u5_n121 ) , .A2( u0_u7_u5_n145 ) , .A1( u0_u7_u5_n176 ) );
  AOI22_X1 u0_u7_u5_U48 (.ZN( u0_u7_u5_n114 ) , .A2( u0_u7_u5_n137 ) , .A1( u0_u7_u5_n145 ) , .B2( u0_u7_u5_n175 ) , .B1( u0_u7_u5_n193 ) );
  OAI211_X1 u0_u7_u5_U49 (.B( u0_u7_u5_n124 ) , .A( u0_u7_u5_n125 ) , .C2( u0_u7_u5_n126 ) , .C1( u0_u7_u5_n127 ) , .ZN( u0_u7_u5_n128 ) );
  OAI21_X1 u0_u7_u5_U5 (.B2( u0_u7_u5_n136 ) , .B1( u0_u7_u5_n137 ) , .ZN( u0_u7_u5_n138 ) , .A( u0_u7_u5_n177 ) );
  NOR3_X1 u0_u7_u5_U50 (.ZN( u0_u7_u5_n127 ) , .A1( u0_u7_u5_n136 ) , .A3( u0_u7_u5_n148 ) , .A2( u0_u7_u5_n182 ) );
  OAI21_X1 u0_u7_u5_U51 (.ZN( u0_u7_u5_n124 ) , .A( u0_u7_u5_n177 ) , .B2( u0_u7_u5_n183 ) , .B1( u0_u7_u5_n189 ) );
  OAI21_X1 u0_u7_u5_U52 (.ZN( u0_u7_u5_n125 ) , .A( u0_u7_u5_n174 ) , .B2( u0_u7_u5_n185 ) , .B1( u0_u7_u5_n190 ) );
  AOI21_X1 u0_u7_u5_U53 (.A( u0_u7_u5_n153 ) , .B2( u0_u7_u5_n154 ) , .B1( u0_u7_u5_n155 ) , .ZN( u0_u7_u5_n164 ) );
  AOI21_X1 u0_u7_u5_U54 (.ZN( u0_u7_u5_n110 ) , .B1( u0_u7_u5_n122 ) , .B2( u0_u7_u5_n139 ) , .A( u0_u7_u5_n153 ) );
  INV_X1 u0_u7_u5_U55 (.A( u0_u7_u5_n153 ) , .ZN( u0_u7_u5_n176 ) );
  INV_X1 u0_u7_u5_U56 (.A( u0_u7_u5_n126 ) , .ZN( u0_u7_u5_n173 ) );
  AND2_X1 u0_u7_u5_U57 (.A2( u0_u7_u5_n104 ) , .A1( u0_u7_u5_n107 ) , .ZN( u0_u7_u5_n147 ) );
  AND2_X1 u0_u7_u5_U58 (.A2( u0_u7_u5_n104 ) , .A1( u0_u7_u5_n108 ) , .ZN( u0_u7_u5_n148 ) );
  NAND2_X1 u0_u7_u5_U59 (.A1( u0_u7_u5_n105 ) , .A2( u0_u7_u5_n106 ) , .ZN( u0_u7_u5_n158 ) );
  INV_X1 u0_u7_u5_U6 (.A( u0_u7_u5_n135 ) , .ZN( u0_u7_u5_n178 ) );
  NAND2_X1 u0_u7_u5_U60 (.A2( u0_u7_u5_n108 ) , .A1( u0_u7_u5_n109 ) , .ZN( u0_u7_u5_n139 ) );
  NAND2_X1 u0_u7_u5_U61 (.A1( u0_u7_u5_n106 ) , .A2( u0_u7_u5_n108 ) , .ZN( u0_u7_u5_n119 ) );
  NAND2_X1 u0_u7_u5_U62 (.A2( u0_u7_u5_n103 ) , .A1( u0_u7_u5_n105 ) , .ZN( u0_u7_u5_n140 ) );
  NAND2_X1 u0_u7_u5_U63 (.A2( u0_u7_u5_n104 ) , .A1( u0_u7_u5_n105 ) , .ZN( u0_u7_u5_n155 ) );
  NAND2_X1 u0_u7_u5_U64 (.A2( u0_u7_u5_n106 ) , .A1( u0_u7_u5_n107 ) , .ZN( u0_u7_u5_n122 ) );
  NAND2_X1 u0_u7_u5_U65 (.A2( u0_u7_u5_n100 ) , .A1( u0_u7_u5_n106 ) , .ZN( u0_u7_u5_n115 ) );
  NAND2_X1 u0_u7_u5_U66 (.A2( u0_u7_u5_n100 ) , .A1( u0_u7_u5_n103 ) , .ZN( u0_u7_u5_n161 ) );
  NAND2_X1 u0_u7_u5_U67 (.A1( u0_u7_u5_n105 ) , .A2( u0_u7_u5_n109 ) , .ZN( u0_u7_u5_n154 ) );
  INV_X1 u0_u7_u5_U68 (.A( u0_u7_u5_n146 ) , .ZN( u0_u7_u5_n172 ) );
  NAND2_X1 u0_u7_u5_U69 (.A1( u0_u7_u5_n103 ) , .A2( u0_u7_u5_n108 ) , .ZN( u0_u7_u5_n123 ) );
  OAI22_X1 u0_u7_u5_U7 (.B2( u0_u7_u5_n149 ) , .B1( u0_u7_u5_n150 ) , .A2( u0_u7_u5_n151 ) , .A1( u0_u7_u5_n152 ) , .ZN( u0_u7_u5_n165 ) );
  NAND2_X1 u0_u7_u5_U70 (.A2( u0_u7_u5_n103 ) , .A1( u0_u7_u5_n107 ) , .ZN( u0_u7_u5_n151 ) );
  NAND2_X1 u0_u7_u5_U71 (.A2( u0_u7_u5_n107 ) , .A1( u0_u7_u5_n109 ) , .ZN( u0_u7_u5_n120 ) );
  NAND2_X1 u0_u7_u5_U72 (.A2( u0_u7_u5_n100 ) , .A1( u0_u7_u5_n109 ) , .ZN( u0_u7_u5_n157 ) );
  AND2_X1 u0_u7_u5_U73 (.A2( u0_u7_u5_n100 ) , .A1( u0_u7_u5_n104 ) , .ZN( u0_u7_u5_n131 ) );
  INV_X1 u0_u7_u5_U74 (.A( u0_u7_u5_n102 ) , .ZN( u0_u7_u5_n195 ) );
  OAI221_X1 u0_u7_u5_U75 (.A( u0_u7_u5_n101 ) , .ZN( u0_u7_u5_n102 ) , .C2( u0_u7_u5_n115 ) , .C1( u0_u7_u5_n126 ) , .B1( u0_u7_u5_n134 ) , .B2( u0_u7_u5_n160 ) );
  OAI21_X1 u0_u7_u5_U76 (.ZN( u0_u7_u5_n101 ) , .B1( u0_u7_u5_n137 ) , .A( u0_u7_u5_n146 ) , .B2( u0_u7_u5_n147 ) );
  NOR2_X1 u0_u7_u5_U77 (.A2( u0_u7_X_34 ) , .A1( u0_u7_X_35 ) , .ZN( u0_u7_u5_n145 ) );
  NOR2_X1 u0_u7_u5_U78 (.A2( u0_u7_X_34 ) , .ZN( u0_u7_u5_n146 ) , .A1( u0_u7_u5_n171 ) );
  NOR2_X1 u0_u7_u5_U79 (.A2( u0_u7_X_31 ) , .A1( u0_u7_X_32 ) , .ZN( u0_u7_u5_n103 ) );
  NOR3_X1 u0_u7_u5_U8 (.A2( u0_u7_u5_n147 ) , .A1( u0_u7_u5_n148 ) , .ZN( u0_u7_u5_n149 ) , .A3( u0_u7_u5_n194 ) );
  NOR2_X1 u0_u7_u5_U80 (.A2( u0_u7_X_36 ) , .ZN( u0_u7_u5_n105 ) , .A1( u0_u7_u5_n180 ) );
  NOR2_X1 u0_u7_u5_U81 (.A2( u0_u7_X_33 ) , .ZN( u0_u7_u5_n108 ) , .A1( u0_u7_u5_n170 ) );
  NOR2_X1 u0_u7_u5_U82 (.A2( u0_u7_X_33 ) , .A1( u0_u7_X_36 ) , .ZN( u0_u7_u5_n107 ) );
  NOR2_X1 u0_u7_u5_U83 (.A2( u0_u7_X_31 ) , .ZN( u0_u7_u5_n104 ) , .A1( u0_u7_u5_n181 ) );
  NAND2_X1 u0_u7_u5_U84 (.A2( u0_u7_X_34 ) , .A1( u0_u7_X_35 ) , .ZN( u0_u7_u5_n153 ) );
  NAND2_X1 u0_u7_u5_U85 (.A1( u0_u7_X_34 ) , .ZN( u0_u7_u5_n126 ) , .A2( u0_u7_u5_n171 ) );
  AND2_X1 u0_u7_u5_U86 (.A1( u0_u7_X_31 ) , .A2( u0_u7_X_32 ) , .ZN( u0_u7_u5_n106 ) );
  AND2_X1 u0_u7_u5_U87 (.A1( u0_u7_X_31 ) , .ZN( u0_u7_u5_n109 ) , .A2( u0_u7_u5_n181 ) );
  INV_X1 u0_u7_u5_U88 (.A( u0_u7_X_33 ) , .ZN( u0_u7_u5_n180 ) );
  INV_X1 u0_u7_u5_U89 (.A( u0_u7_X_35 ) , .ZN( u0_u7_u5_n171 ) );
  NOR2_X1 u0_u7_u5_U9 (.ZN( u0_u7_u5_n135 ) , .A1( u0_u7_u5_n173 ) , .A2( u0_u7_u5_n176 ) );
  INV_X1 u0_u7_u5_U90 (.A( u0_u7_X_36 ) , .ZN( u0_u7_u5_n170 ) );
  INV_X1 u0_u7_u5_U91 (.A( u0_u7_X_32 ) , .ZN( u0_u7_u5_n181 ) );
  NAND4_X1 u0_u7_u5_U92 (.ZN( u0_out7_29 ) , .A4( u0_u7_u5_n129 ) , .A3( u0_u7_u5_n130 ) , .A2( u0_u7_u5_n168 ) , .A1( u0_u7_u5_n196 ) );
  AOI221_X1 u0_u7_u5_U93 (.A( u0_u7_u5_n128 ) , .ZN( u0_u7_u5_n129 ) , .C2( u0_u7_u5_n132 ) , .B2( u0_u7_u5_n159 ) , .B1( u0_u7_u5_n176 ) , .C1( u0_u7_u5_n184 ) );
  AOI222_X1 u0_u7_u5_U94 (.ZN( u0_u7_u5_n130 ) , .A2( u0_u7_u5_n146 ) , .B1( u0_u7_u5_n147 ) , .C2( u0_u7_u5_n175 ) , .B2( u0_u7_u5_n179 ) , .A1( u0_u7_u5_n188 ) , .C1( u0_u7_u5_n194 ) );
  NAND4_X1 u0_u7_u5_U95 (.ZN( u0_out7_19 ) , .A4( u0_u7_u5_n166 ) , .A3( u0_u7_u5_n167 ) , .A2( u0_u7_u5_n168 ) , .A1( u0_u7_u5_n169 ) );
  AOI22_X1 u0_u7_u5_U96 (.B2( u0_u7_u5_n145 ) , .A2( u0_u7_u5_n146 ) , .ZN( u0_u7_u5_n167 ) , .B1( u0_u7_u5_n182 ) , .A1( u0_u7_u5_n189 ) );
  NOR4_X1 u0_u7_u5_U97 (.A4( u0_u7_u5_n162 ) , .A3( u0_u7_u5_n163 ) , .A2( u0_u7_u5_n164 ) , .A1( u0_u7_u5_n165 ) , .ZN( u0_u7_u5_n166 ) );
  NAND4_X1 u0_u7_u5_U98 (.ZN( u0_out7_11 ) , .A4( u0_u7_u5_n143 ) , .A3( u0_u7_u5_n144 ) , .A2( u0_u7_u5_n169 ) , .A1( u0_u7_u5_n196 ) );
  AOI22_X1 u0_u7_u5_U99 (.A2( u0_u7_u5_n132 ) , .ZN( u0_u7_u5_n144 ) , .B2( u0_u7_u5_n145 ) , .B1( u0_u7_u5_n184 ) , .A1( u0_u7_u5_n194 ) );
  INV_X1 u0_u7_u6_U10 (.ZN( u0_u7_u6_n172 ) , .A( u0_u7_u6_n88 ) );
  OAI21_X1 u0_u7_u6_U11 (.A( u0_u7_u6_n159 ) , .B1( u0_u7_u6_n169 ) , .B2( u0_u7_u6_n173 ) , .ZN( u0_u7_u6_n90 ) );
  AOI22_X1 u0_u7_u6_U12 (.A2( u0_u7_u6_n151 ) , .B2( u0_u7_u6_n161 ) , .A1( u0_u7_u6_n167 ) , .B1( u0_u7_u6_n170 ) , .ZN( u0_u7_u6_n89 ) );
  AOI21_X1 u0_u7_u6_U13 (.ZN( u0_u7_u6_n106 ) , .A( u0_u7_u6_n142 ) , .B2( u0_u7_u6_n159 ) , .B1( u0_u7_u6_n164 ) );
  INV_X1 u0_u7_u6_U14 (.A( u0_u7_u6_n155 ) , .ZN( u0_u7_u6_n161 ) );
  INV_X1 u0_u7_u6_U15 (.A( u0_u7_u6_n128 ) , .ZN( u0_u7_u6_n164 ) );
  NAND2_X1 u0_u7_u6_U16 (.ZN( u0_u7_u6_n110 ) , .A1( u0_u7_u6_n122 ) , .A2( u0_u7_u6_n129 ) );
  NAND2_X1 u0_u7_u6_U17 (.ZN( u0_u7_u6_n124 ) , .A2( u0_u7_u6_n146 ) , .A1( u0_u7_u6_n148 ) );
  INV_X1 u0_u7_u6_U18 (.A( u0_u7_u6_n132 ) , .ZN( u0_u7_u6_n171 ) );
  AND2_X1 u0_u7_u6_U19 (.A1( u0_u7_u6_n100 ) , .ZN( u0_u7_u6_n130 ) , .A2( u0_u7_u6_n147 ) );
  INV_X1 u0_u7_u6_U20 (.A( u0_u7_u6_n127 ) , .ZN( u0_u7_u6_n173 ) );
  INV_X1 u0_u7_u6_U21 (.A( u0_u7_u6_n121 ) , .ZN( u0_u7_u6_n167 ) );
  INV_X1 u0_u7_u6_U22 (.A( u0_u7_u6_n100 ) , .ZN( u0_u7_u6_n169 ) );
  INV_X1 u0_u7_u6_U23 (.A( u0_u7_u6_n123 ) , .ZN( u0_u7_u6_n170 ) );
  INV_X1 u0_u7_u6_U24 (.A( u0_u7_u6_n113 ) , .ZN( u0_u7_u6_n168 ) );
  AND2_X1 u0_u7_u6_U25 (.A1( u0_u7_u6_n107 ) , .A2( u0_u7_u6_n119 ) , .ZN( u0_u7_u6_n133 ) );
  AND2_X1 u0_u7_u6_U26 (.A2( u0_u7_u6_n121 ) , .A1( u0_u7_u6_n122 ) , .ZN( u0_u7_u6_n131 ) );
  AND3_X1 u0_u7_u6_U27 (.ZN( u0_u7_u6_n120 ) , .A2( u0_u7_u6_n127 ) , .A1( u0_u7_u6_n132 ) , .A3( u0_u7_u6_n145 ) );
  INV_X1 u0_u7_u6_U28 (.A( u0_u7_u6_n146 ) , .ZN( u0_u7_u6_n163 ) );
  AOI222_X1 u0_u7_u6_U29 (.ZN( u0_u7_u6_n114 ) , .A1( u0_u7_u6_n118 ) , .A2( u0_u7_u6_n126 ) , .B2( u0_u7_u6_n151 ) , .C2( u0_u7_u6_n159 ) , .C1( u0_u7_u6_n168 ) , .B1( u0_u7_u6_n169 ) );
  INV_X1 u0_u7_u6_U3 (.A( u0_u7_u6_n110 ) , .ZN( u0_u7_u6_n166 ) );
  NOR2_X1 u0_u7_u6_U30 (.A1( u0_u7_u6_n162 ) , .A2( u0_u7_u6_n165 ) , .ZN( u0_u7_u6_n98 ) );
  NAND2_X1 u0_u7_u6_U31 (.A1( u0_u7_u6_n144 ) , .ZN( u0_u7_u6_n151 ) , .A2( u0_u7_u6_n158 ) );
  NAND2_X1 u0_u7_u6_U32 (.ZN( u0_u7_u6_n132 ) , .A1( u0_u7_u6_n91 ) , .A2( u0_u7_u6_n97 ) );
  AOI22_X1 u0_u7_u6_U33 (.B2( u0_u7_u6_n110 ) , .B1( u0_u7_u6_n111 ) , .A1( u0_u7_u6_n112 ) , .ZN( u0_u7_u6_n115 ) , .A2( u0_u7_u6_n161 ) );
  NAND4_X1 u0_u7_u6_U34 (.A3( u0_u7_u6_n109 ) , .ZN( u0_u7_u6_n112 ) , .A4( u0_u7_u6_n132 ) , .A2( u0_u7_u6_n147 ) , .A1( u0_u7_u6_n166 ) );
  NOR2_X1 u0_u7_u6_U35 (.ZN( u0_u7_u6_n109 ) , .A1( u0_u7_u6_n170 ) , .A2( u0_u7_u6_n173 ) );
  NOR2_X1 u0_u7_u6_U36 (.A2( u0_u7_u6_n126 ) , .ZN( u0_u7_u6_n155 ) , .A1( u0_u7_u6_n160 ) );
  NAND2_X1 u0_u7_u6_U37 (.ZN( u0_u7_u6_n146 ) , .A2( u0_u7_u6_n94 ) , .A1( u0_u7_u6_n99 ) );
  AOI21_X1 u0_u7_u6_U38 (.A( u0_u7_u6_n144 ) , .B2( u0_u7_u6_n145 ) , .B1( u0_u7_u6_n146 ) , .ZN( u0_u7_u6_n150 ) );
  AOI211_X1 u0_u7_u6_U39 (.B( u0_u7_u6_n134 ) , .A( u0_u7_u6_n135 ) , .C1( u0_u7_u6_n136 ) , .ZN( u0_u7_u6_n137 ) , .C2( u0_u7_u6_n151 ) );
  INV_X1 u0_u7_u6_U4 (.A( u0_u7_u6_n142 ) , .ZN( u0_u7_u6_n174 ) );
  NAND4_X1 u0_u7_u6_U40 (.A4( u0_u7_u6_n127 ) , .A3( u0_u7_u6_n128 ) , .A2( u0_u7_u6_n129 ) , .A1( u0_u7_u6_n130 ) , .ZN( u0_u7_u6_n136 ) );
  AOI21_X1 u0_u7_u6_U41 (.B2( u0_u7_u6_n132 ) , .B1( u0_u7_u6_n133 ) , .ZN( u0_u7_u6_n134 ) , .A( u0_u7_u6_n158 ) );
  AOI21_X1 u0_u7_u6_U42 (.B1( u0_u7_u6_n131 ) , .ZN( u0_u7_u6_n135 ) , .A( u0_u7_u6_n144 ) , .B2( u0_u7_u6_n146 ) );
  INV_X1 u0_u7_u6_U43 (.A( u0_u7_u6_n111 ) , .ZN( u0_u7_u6_n158 ) );
  NAND2_X1 u0_u7_u6_U44 (.ZN( u0_u7_u6_n127 ) , .A1( u0_u7_u6_n91 ) , .A2( u0_u7_u6_n92 ) );
  NAND2_X1 u0_u7_u6_U45 (.ZN( u0_u7_u6_n129 ) , .A2( u0_u7_u6_n95 ) , .A1( u0_u7_u6_n96 ) );
  INV_X1 u0_u7_u6_U46 (.A( u0_u7_u6_n144 ) , .ZN( u0_u7_u6_n159 ) );
  NAND2_X1 u0_u7_u6_U47 (.ZN( u0_u7_u6_n145 ) , .A2( u0_u7_u6_n97 ) , .A1( u0_u7_u6_n98 ) );
  NAND2_X1 u0_u7_u6_U48 (.ZN( u0_u7_u6_n148 ) , .A2( u0_u7_u6_n92 ) , .A1( u0_u7_u6_n94 ) );
  NAND2_X1 u0_u7_u6_U49 (.ZN( u0_u7_u6_n108 ) , .A2( u0_u7_u6_n139 ) , .A1( u0_u7_u6_n144 ) );
  NAND2_X1 u0_u7_u6_U5 (.A2( u0_u7_u6_n143 ) , .ZN( u0_u7_u6_n152 ) , .A1( u0_u7_u6_n166 ) );
  NAND2_X1 u0_u7_u6_U50 (.ZN( u0_u7_u6_n121 ) , .A2( u0_u7_u6_n95 ) , .A1( u0_u7_u6_n97 ) );
  NAND2_X1 u0_u7_u6_U51 (.ZN( u0_u7_u6_n107 ) , .A2( u0_u7_u6_n92 ) , .A1( u0_u7_u6_n95 ) );
  AND2_X1 u0_u7_u6_U52 (.ZN( u0_u7_u6_n118 ) , .A2( u0_u7_u6_n91 ) , .A1( u0_u7_u6_n99 ) );
  NAND2_X1 u0_u7_u6_U53 (.ZN( u0_u7_u6_n147 ) , .A2( u0_u7_u6_n98 ) , .A1( u0_u7_u6_n99 ) );
  NAND2_X1 u0_u7_u6_U54 (.ZN( u0_u7_u6_n128 ) , .A1( u0_u7_u6_n94 ) , .A2( u0_u7_u6_n96 ) );
  NAND2_X1 u0_u7_u6_U55 (.ZN( u0_u7_u6_n119 ) , .A2( u0_u7_u6_n95 ) , .A1( u0_u7_u6_n99 ) );
  NAND2_X1 u0_u7_u6_U56 (.ZN( u0_u7_u6_n123 ) , .A2( u0_u7_u6_n91 ) , .A1( u0_u7_u6_n96 ) );
  NAND2_X1 u0_u7_u6_U57 (.ZN( u0_u7_u6_n100 ) , .A2( u0_u7_u6_n92 ) , .A1( u0_u7_u6_n98 ) );
  NAND2_X1 u0_u7_u6_U58 (.ZN( u0_u7_u6_n122 ) , .A1( u0_u7_u6_n94 ) , .A2( u0_u7_u6_n97 ) );
  INV_X1 u0_u7_u6_U59 (.A( u0_u7_u6_n139 ) , .ZN( u0_u7_u6_n160 ) );
  AOI22_X1 u0_u7_u6_U6 (.B2( u0_u7_u6_n101 ) , .A1( u0_u7_u6_n102 ) , .ZN( u0_u7_u6_n103 ) , .B1( u0_u7_u6_n160 ) , .A2( u0_u7_u6_n161 ) );
  NAND2_X1 u0_u7_u6_U60 (.ZN( u0_u7_u6_n113 ) , .A1( u0_u7_u6_n96 ) , .A2( u0_u7_u6_n98 ) );
  NOR2_X1 u0_u7_u6_U61 (.A2( u0_u7_X_40 ) , .A1( u0_u7_X_41 ) , .ZN( u0_u7_u6_n126 ) );
  NOR2_X1 u0_u7_u6_U62 (.A2( u0_u7_X_39 ) , .A1( u0_u7_X_42 ) , .ZN( u0_u7_u6_n92 ) );
  NOR2_X1 u0_u7_u6_U63 (.A2( u0_u7_X_39 ) , .A1( u0_u7_u6_n156 ) , .ZN( u0_u7_u6_n97 ) );
  NOR2_X1 u0_u7_u6_U64 (.A2( u0_u7_X_38 ) , .A1( u0_u7_u6_n165 ) , .ZN( u0_u7_u6_n95 ) );
  NOR2_X1 u0_u7_u6_U65 (.A2( u0_u7_X_41 ) , .ZN( u0_u7_u6_n111 ) , .A1( u0_u7_u6_n157 ) );
  NOR2_X1 u0_u7_u6_U66 (.A2( u0_u7_X_37 ) , .A1( u0_u7_u6_n162 ) , .ZN( u0_u7_u6_n94 ) );
  NOR2_X1 u0_u7_u6_U67 (.A2( u0_u7_X_37 ) , .A1( u0_u7_X_38 ) , .ZN( u0_u7_u6_n91 ) );
  NAND2_X1 u0_u7_u6_U68 (.A1( u0_u7_X_41 ) , .ZN( u0_u7_u6_n144 ) , .A2( u0_u7_u6_n157 ) );
  NAND2_X1 u0_u7_u6_U69 (.A2( u0_u7_X_40 ) , .A1( u0_u7_X_41 ) , .ZN( u0_u7_u6_n139 ) );
  NOR2_X1 u0_u7_u6_U7 (.A1( u0_u7_u6_n118 ) , .ZN( u0_u7_u6_n143 ) , .A2( u0_u7_u6_n168 ) );
  AND2_X1 u0_u7_u6_U70 (.A1( u0_u7_X_39 ) , .A2( u0_u7_u6_n156 ) , .ZN( u0_u7_u6_n96 ) );
  AND2_X1 u0_u7_u6_U71 (.A1( u0_u7_X_39 ) , .A2( u0_u7_X_42 ) , .ZN( u0_u7_u6_n99 ) );
  INV_X1 u0_u7_u6_U72 (.A( u0_u7_X_40 ) , .ZN( u0_u7_u6_n157 ) );
  INV_X1 u0_u7_u6_U73 (.A( u0_u7_X_37 ) , .ZN( u0_u7_u6_n165 ) );
  INV_X1 u0_u7_u6_U74 (.A( u0_u7_X_38 ) , .ZN( u0_u7_u6_n162 ) );
  INV_X1 u0_u7_u6_U75 (.A( u0_u7_X_42 ) , .ZN( u0_u7_u6_n156 ) );
  NAND4_X1 u0_u7_u6_U76 (.ZN( u0_out7_32 ) , .A4( u0_u7_u6_n103 ) , .A3( u0_u7_u6_n104 ) , .A2( u0_u7_u6_n105 ) , .A1( u0_u7_u6_n106 ) );
  AOI22_X1 u0_u7_u6_U77 (.ZN( u0_u7_u6_n105 ) , .A2( u0_u7_u6_n108 ) , .A1( u0_u7_u6_n118 ) , .B2( u0_u7_u6_n126 ) , .B1( u0_u7_u6_n171 ) );
  AOI22_X1 u0_u7_u6_U78 (.ZN( u0_u7_u6_n104 ) , .A1( u0_u7_u6_n111 ) , .B1( u0_u7_u6_n124 ) , .B2( u0_u7_u6_n151 ) , .A2( u0_u7_u6_n93 ) );
  NAND4_X1 u0_u7_u6_U79 (.ZN( u0_out7_12 ) , .A4( u0_u7_u6_n114 ) , .A3( u0_u7_u6_n115 ) , .A2( u0_u7_u6_n116 ) , .A1( u0_u7_u6_n117 ) );
  AOI21_X1 u0_u7_u6_U8 (.B1( u0_u7_u6_n107 ) , .B2( u0_u7_u6_n132 ) , .A( u0_u7_u6_n158 ) , .ZN( u0_u7_u6_n88 ) );
  OAI22_X1 u0_u7_u6_U80 (.B2( u0_u7_u6_n111 ) , .ZN( u0_u7_u6_n116 ) , .B1( u0_u7_u6_n126 ) , .A2( u0_u7_u6_n164 ) , .A1( u0_u7_u6_n167 ) );
  OAI21_X1 u0_u7_u6_U81 (.A( u0_u7_u6_n108 ) , .ZN( u0_u7_u6_n117 ) , .B2( u0_u7_u6_n141 ) , .B1( u0_u7_u6_n163 ) );
  OAI211_X1 u0_u7_u6_U82 (.ZN( u0_out7_22 ) , .B( u0_u7_u6_n137 ) , .A( u0_u7_u6_n138 ) , .C2( u0_u7_u6_n139 ) , .C1( u0_u7_u6_n140 ) );
  AOI22_X1 u0_u7_u6_U83 (.B1( u0_u7_u6_n124 ) , .A2( u0_u7_u6_n125 ) , .A1( u0_u7_u6_n126 ) , .ZN( u0_u7_u6_n138 ) , .B2( u0_u7_u6_n161 ) );
  AND4_X1 u0_u7_u6_U84 (.A3( u0_u7_u6_n119 ) , .A1( u0_u7_u6_n120 ) , .A4( u0_u7_u6_n129 ) , .ZN( u0_u7_u6_n140 ) , .A2( u0_u7_u6_n143 ) );
  OAI211_X1 u0_u7_u6_U85 (.ZN( u0_out7_7 ) , .B( u0_u7_u6_n153 ) , .C2( u0_u7_u6_n154 ) , .C1( u0_u7_u6_n155 ) , .A( u0_u7_u6_n174 ) );
  NOR3_X1 u0_u7_u6_U86 (.A1( u0_u7_u6_n141 ) , .ZN( u0_u7_u6_n154 ) , .A3( u0_u7_u6_n164 ) , .A2( u0_u7_u6_n171 ) );
  AOI211_X1 u0_u7_u6_U87 (.B( u0_u7_u6_n149 ) , .A( u0_u7_u6_n150 ) , .C2( u0_u7_u6_n151 ) , .C1( u0_u7_u6_n152 ) , .ZN( u0_u7_u6_n153 ) );
  NAND3_X1 u0_u7_u6_U88 (.A2( u0_u7_u6_n123 ) , .ZN( u0_u7_u6_n125 ) , .A1( u0_u7_u6_n130 ) , .A3( u0_u7_u6_n131 ) );
  NAND3_X1 u0_u7_u6_U89 (.A3( u0_u7_u6_n133 ) , .ZN( u0_u7_u6_n141 ) , .A1( u0_u7_u6_n145 ) , .A2( u0_u7_u6_n148 ) );
  AOI21_X1 u0_u7_u6_U9 (.B2( u0_u7_u6_n147 ) , .B1( u0_u7_u6_n148 ) , .ZN( u0_u7_u6_n149 ) , .A( u0_u7_u6_n158 ) );
  NAND3_X1 u0_u7_u6_U90 (.ZN( u0_u7_u6_n101 ) , .A3( u0_u7_u6_n107 ) , .A2( u0_u7_u6_n121 ) , .A1( u0_u7_u6_n127 ) );
  NAND3_X1 u0_u7_u6_U91 (.ZN( u0_u7_u6_n102 ) , .A3( u0_u7_u6_n130 ) , .A2( u0_u7_u6_n145 ) , .A1( u0_u7_u6_n166 ) );
  NAND3_X1 u0_u7_u6_U92 (.A3( u0_u7_u6_n113 ) , .A1( u0_u7_u6_n119 ) , .A2( u0_u7_u6_n123 ) , .ZN( u0_u7_u6_n93 ) );
  NAND3_X1 u0_u7_u6_U93 (.ZN( u0_u7_u6_n142 ) , .A2( u0_u7_u6_n172 ) , .A3( u0_u7_u6_n89 ) , .A1( u0_u7_u6_n90 ) );
  XOR2_X1 u0_u8_U1 (.B( u0_K9_9 ) , .A( u0_R7_6 ) , .Z( u0_u8_X_9 ) );
  XOR2_X1 u0_u8_U13 (.B( u0_K9_42 ) , .A( u0_R7_29 ) , .Z( u0_u8_X_42 ) );
  XOR2_X1 u0_u8_U14 (.B( u0_K9_41 ) , .A( u0_R7_28 ) , .Z( u0_u8_X_41 ) );
  XOR2_X1 u0_u8_U15 (.B( u0_K9_40 ) , .A( u0_R7_27 ) , .Z( u0_u8_X_40 ) );
  XOR2_X1 u0_u8_U16 (.B( u0_K9_3 ) , .A( u0_R7_2 ) , .Z( u0_u8_X_3 ) );
  XOR2_X1 u0_u8_U17 (.B( u0_K9_39 ) , .A( u0_R7_26 ) , .Z( u0_u8_X_39 ) );
  XOR2_X1 u0_u8_U18 (.B( u0_K9_38 ) , .A( u0_R7_25 ) , .Z( u0_u8_X_38 ) );
  XOR2_X1 u0_u8_U19 (.B( u0_K9_37 ) , .A( u0_R7_24 ) , .Z( u0_u8_X_37 ) );
  XOR2_X1 u0_u8_U2 (.B( u0_K9_8 ) , .A( u0_R7_5 ) , .Z( u0_u8_X_8 ) );
  XOR2_X1 u0_u8_U20 (.B( u0_K9_36 ) , .A( u0_R7_25 ) , .Z( u0_u8_X_36 ) );
  XOR2_X1 u0_u8_U21 (.B( u0_K9_35 ) , .A( u0_R7_24 ) , .Z( u0_u8_X_35 ) );
  XOR2_X1 u0_u8_U22 (.B( u0_K9_34 ) , .A( u0_R7_23 ) , .Z( u0_u8_X_34 ) );
  XOR2_X1 u0_u8_U23 (.B( u0_K9_33 ) , .A( u0_R7_22 ) , .Z( u0_u8_X_33 ) );
  XOR2_X1 u0_u8_U24 (.B( u0_K9_32 ) , .A( u0_R7_21 ) , .Z( u0_u8_X_32 ) );
  XOR2_X1 u0_u8_U25 (.B( u0_K9_31 ) , .A( u0_R7_20 ) , .Z( u0_u8_X_31 ) );
  XOR2_X1 u0_u8_U27 (.B( u0_K9_2 ) , .A( u0_R7_1 ) , .Z( u0_u8_X_2 ) );
  XOR2_X1 u0_u8_U3 (.B( u0_K9_7 ) , .A( u0_R7_4 ) , .Z( u0_u8_X_7 ) );
  XOR2_X1 u0_u8_U38 (.B( u0_K9_1 ) , .A( u0_R7_32 ) , .Z( u0_u8_X_1 ) );
  XOR2_X1 u0_u8_U4 (.B( u0_K9_6 ) , .A( u0_R7_5 ) , .Z( u0_u8_X_6 ) );
  XOR2_X1 u0_u8_U40 (.B( u0_K9_18 ) , .A( u0_R7_13 ) , .Z( u0_u8_X_18 ) );
  XOR2_X1 u0_u8_U41 (.B( u0_K9_17 ) , .A( u0_R7_12 ) , .Z( u0_u8_X_17 ) );
  XOR2_X1 u0_u8_U42 (.B( u0_K9_16 ) , .A( u0_R7_11 ) , .Z( u0_u8_X_16 ) );
  XOR2_X1 u0_u8_U43 (.B( u0_K9_15 ) , .A( u0_R7_10 ) , .Z( u0_u8_X_15 ) );
  XOR2_X1 u0_u8_U44 (.B( u0_K9_14 ) , .A( u0_R7_9 ) , .Z( u0_u8_X_14 ) );
  XOR2_X1 u0_u8_U45 (.B( u0_K9_13 ) , .A( u0_R7_8 ) , .Z( u0_u8_X_13 ) );
  XOR2_X1 u0_u8_U46 (.B( u0_K9_12 ) , .A( u0_R7_9 ) , .Z( u0_u8_X_12 ) );
  XOR2_X1 u0_u8_U47 (.B( u0_K9_11 ) , .A( u0_R7_8 ) , .Z( u0_u8_X_11 ) );
  XOR2_X1 u0_u8_U48 (.B( u0_K9_10 ) , .A( u0_R7_7 ) , .Z( u0_u8_X_10 ) );
  XOR2_X1 u0_u8_U5 (.B( u0_K9_5 ) , .A( u0_R7_4 ) , .Z( u0_u8_X_5 ) );
  XOR2_X1 u0_u8_U6 (.B( u0_K9_4 ) , .A( u0_R7_3 ) , .Z( u0_u8_X_4 ) );
  AND3_X1 u0_u8_u0_U10 (.A2( u0_u8_u0_n112 ) , .ZN( u0_u8_u0_n127 ) , .A3( u0_u8_u0_n130 ) , .A1( u0_u8_u0_n148 ) );
  NAND2_X1 u0_u8_u0_U11 (.ZN( u0_u8_u0_n113 ) , .A1( u0_u8_u0_n139 ) , .A2( u0_u8_u0_n149 ) );
  AND2_X1 u0_u8_u0_U12 (.ZN( u0_u8_u0_n107 ) , .A1( u0_u8_u0_n130 ) , .A2( u0_u8_u0_n140 ) );
  AND2_X1 u0_u8_u0_U13 (.A2( u0_u8_u0_n129 ) , .A1( u0_u8_u0_n130 ) , .ZN( u0_u8_u0_n151 ) );
  AND2_X1 u0_u8_u0_U14 (.A1( u0_u8_u0_n108 ) , .A2( u0_u8_u0_n125 ) , .ZN( u0_u8_u0_n145 ) );
  INV_X1 u0_u8_u0_U15 (.A( u0_u8_u0_n143 ) , .ZN( u0_u8_u0_n173 ) );
  NOR2_X1 u0_u8_u0_U16 (.A2( u0_u8_u0_n136 ) , .ZN( u0_u8_u0_n147 ) , .A1( u0_u8_u0_n160 ) );
  AOI21_X1 u0_u8_u0_U17 (.B1( u0_u8_u0_n103 ) , .ZN( u0_u8_u0_n132 ) , .A( u0_u8_u0_n165 ) , .B2( u0_u8_u0_n93 ) );
  INV_X1 u0_u8_u0_U18 (.A( u0_u8_u0_n142 ) , .ZN( u0_u8_u0_n165 ) );
  OAI22_X1 u0_u8_u0_U19 (.B1( u0_u8_u0_n125 ) , .ZN( u0_u8_u0_n126 ) , .A1( u0_u8_u0_n138 ) , .A2( u0_u8_u0_n146 ) , .B2( u0_u8_u0_n147 ) );
  OAI22_X1 u0_u8_u0_U20 (.B1( u0_u8_u0_n131 ) , .A1( u0_u8_u0_n144 ) , .B2( u0_u8_u0_n147 ) , .A2( u0_u8_u0_n90 ) , .ZN( u0_u8_u0_n91 ) );
  AND3_X1 u0_u8_u0_U21 (.A3( u0_u8_u0_n121 ) , .A2( u0_u8_u0_n125 ) , .A1( u0_u8_u0_n148 ) , .ZN( u0_u8_u0_n90 ) );
  INV_X1 u0_u8_u0_U22 (.A( u0_u8_u0_n136 ) , .ZN( u0_u8_u0_n161 ) );
  AOI22_X1 u0_u8_u0_U23 (.B2( u0_u8_u0_n109 ) , .A2( u0_u8_u0_n110 ) , .ZN( u0_u8_u0_n111 ) , .B1( u0_u8_u0_n118 ) , .A1( u0_u8_u0_n160 ) );
  INV_X1 u0_u8_u0_U24 (.A( u0_u8_u0_n118 ) , .ZN( u0_u8_u0_n158 ) );
  AOI21_X1 u0_u8_u0_U25 (.ZN( u0_u8_u0_n104 ) , .B1( u0_u8_u0_n107 ) , .B2( u0_u8_u0_n141 ) , .A( u0_u8_u0_n144 ) );
  AOI21_X1 u0_u8_u0_U26 (.B1( u0_u8_u0_n127 ) , .B2( u0_u8_u0_n129 ) , .A( u0_u8_u0_n138 ) , .ZN( u0_u8_u0_n96 ) );
  AOI21_X1 u0_u8_u0_U27 (.ZN( u0_u8_u0_n116 ) , .B2( u0_u8_u0_n142 ) , .A( u0_u8_u0_n144 ) , .B1( u0_u8_u0_n166 ) );
  NOR2_X1 u0_u8_u0_U28 (.A1( u0_u8_u0_n120 ) , .ZN( u0_u8_u0_n143 ) , .A2( u0_u8_u0_n167 ) );
  OAI221_X1 u0_u8_u0_U29 (.C1( u0_u8_u0_n112 ) , .ZN( u0_u8_u0_n120 ) , .B1( u0_u8_u0_n138 ) , .B2( u0_u8_u0_n141 ) , .C2( u0_u8_u0_n147 ) , .A( u0_u8_u0_n172 ) );
  INV_X1 u0_u8_u0_U3 (.A( u0_u8_u0_n113 ) , .ZN( u0_u8_u0_n166 ) );
  AOI211_X1 u0_u8_u0_U30 (.B( u0_u8_u0_n115 ) , .A( u0_u8_u0_n116 ) , .C2( u0_u8_u0_n117 ) , .C1( u0_u8_u0_n118 ) , .ZN( u0_u8_u0_n119 ) );
  NAND2_X1 u0_u8_u0_U31 (.A1( u0_u8_u0_n100 ) , .A2( u0_u8_u0_n103 ) , .ZN( u0_u8_u0_n125 ) );
  NAND2_X1 u0_u8_u0_U32 (.A2( u0_u8_u0_n103 ) , .ZN( u0_u8_u0_n140 ) , .A1( u0_u8_u0_n94 ) );
  NAND2_X1 u0_u8_u0_U33 (.A1( u0_u8_u0_n101 ) , .A2( u0_u8_u0_n102 ) , .ZN( u0_u8_u0_n150 ) );
  INV_X1 u0_u8_u0_U34 (.A( u0_u8_u0_n138 ) , .ZN( u0_u8_u0_n160 ) );
  NAND2_X1 u0_u8_u0_U35 (.A2( u0_u8_u0_n102 ) , .A1( u0_u8_u0_n103 ) , .ZN( u0_u8_u0_n149 ) );
  NAND2_X1 u0_u8_u0_U36 (.A2( u0_u8_u0_n100 ) , .A1( u0_u8_u0_n101 ) , .ZN( u0_u8_u0_n139 ) );
  NAND2_X1 u0_u8_u0_U37 (.A2( u0_u8_u0_n100 ) , .ZN( u0_u8_u0_n131 ) , .A1( u0_u8_u0_n92 ) );
  NAND2_X1 u0_u8_u0_U38 (.ZN( u0_u8_u0_n108 ) , .A1( u0_u8_u0_n92 ) , .A2( u0_u8_u0_n94 ) );
  NAND2_X1 u0_u8_u0_U39 (.A2( u0_u8_u0_n102 ) , .ZN( u0_u8_u0_n114 ) , .A1( u0_u8_u0_n92 ) );
  AOI21_X1 u0_u8_u0_U4 (.B1( u0_u8_u0_n114 ) , .ZN( u0_u8_u0_n115 ) , .B2( u0_u8_u0_n129 ) , .A( u0_u8_u0_n161 ) );
  NAND2_X1 u0_u8_u0_U40 (.A1( u0_u8_u0_n101 ) , .ZN( u0_u8_u0_n130 ) , .A2( u0_u8_u0_n94 ) );
  NAND2_X1 u0_u8_u0_U41 (.A2( u0_u8_u0_n101 ) , .ZN( u0_u8_u0_n121 ) , .A1( u0_u8_u0_n93 ) );
  INV_X1 u0_u8_u0_U42 (.ZN( u0_u8_u0_n172 ) , .A( u0_u8_u0_n88 ) );
  OAI222_X1 u0_u8_u0_U43 (.C1( u0_u8_u0_n108 ) , .A1( u0_u8_u0_n125 ) , .B2( u0_u8_u0_n128 ) , .B1( u0_u8_u0_n144 ) , .A2( u0_u8_u0_n158 ) , .C2( u0_u8_u0_n161 ) , .ZN( u0_u8_u0_n88 ) );
  NAND2_X1 u0_u8_u0_U44 (.ZN( u0_u8_u0_n112 ) , .A2( u0_u8_u0_n92 ) , .A1( u0_u8_u0_n93 ) );
  OR3_X1 u0_u8_u0_U45 (.A3( u0_u8_u0_n152 ) , .A2( u0_u8_u0_n153 ) , .A1( u0_u8_u0_n154 ) , .ZN( u0_u8_u0_n155 ) );
  AOI21_X1 u0_u8_u0_U46 (.A( u0_u8_u0_n144 ) , .B2( u0_u8_u0_n145 ) , .B1( u0_u8_u0_n146 ) , .ZN( u0_u8_u0_n154 ) );
  AOI21_X1 u0_u8_u0_U47 (.B2( u0_u8_u0_n150 ) , .B1( u0_u8_u0_n151 ) , .ZN( u0_u8_u0_n152 ) , .A( u0_u8_u0_n158 ) );
  AOI21_X1 u0_u8_u0_U48 (.A( u0_u8_u0_n147 ) , .B2( u0_u8_u0_n148 ) , .B1( u0_u8_u0_n149 ) , .ZN( u0_u8_u0_n153 ) );
  INV_X1 u0_u8_u0_U49 (.ZN( u0_u8_u0_n171 ) , .A( u0_u8_u0_n99 ) );
  AOI21_X1 u0_u8_u0_U5 (.B2( u0_u8_u0_n131 ) , .ZN( u0_u8_u0_n134 ) , .B1( u0_u8_u0_n151 ) , .A( u0_u8_u0_n158 ) );
  OAI211_X1 u0_u8_u0_U50 (.C2( u0_u8_u0_n140 ) , .C1( u0_u8_u0_n161 ) , .A( u0_u8_u0_n169 ) , .B( u0_u8_u0_n98 ) , .ZN( u0_u8_u0_n99 ) );
  INV_X1 u0_u8_u0_U51 (.ZN( u0_u8_u0_n169 ) , .A( u0_u8_u0_n91 ) );
  AOI211_X1 u0_u8_u0_U52 (.C1( u0_u8_u0_n118 ) , .A( u0_u8_u0_n123 ) , .B( u0_u8_u0_n96 ) , .C2( u0_u8_u0_n97 ) , .ZN( u0_u8_u0_n98 ) );
  NOR2_X1 u0_u8_u0_U53 (.A2( u0_u8_X_2 ) , .ZN( u0_u8_u0_n103 ) , .A1( u0_u8_u0_n164 ) );
  NOR2_X1 u0_u8_u0_U54 (.A2( u0_u8_X_4 ) , .A1( u0_u8_X_5 ) , .ZN( u0_u8_u0_n118 ) );
  NOR2_X1 u0_u8_u0_U55 (.A2( u0_u8_X_1 ) , .A1( u0_u8_X_2 ) , .ZN( u0_u8_u0_n92 ) );
  NOR2_X1 u0_u8_u0_U56 (.A2( u0_u8_X_1 ) , .ZN( u0_u8_u0_n101 ) , .A1( u0_u8_u0_n163 ) );
  NOR2_X1 u0_u8_u0_U57 (.A2( u0_u8_X_3 ) , .A1( u0_u8_X_6 ) , .ZN( u0_u8_u0_n94 ) );
  NOR2_X1 u0_u8_u0_U58 (.A2( u0_u8_X_6 ) , .ZN( u0_u8_u0_n100 ) , .A1( u0_u8_u0_n162 ) );
  NAND2_X1 u0_u8_u0_U59 (.A2( u0_u8_X_4 ) , .A1( u0_u8_X_5 ) , .ZN( u0_u8_u0_n144 ) );
  NOR2_X1 u0_u8_u0_U6 (.A1( u0_u8_u0_n108 ) , .ZN( u0_u8_u0_n123 ) , .A2( u0_u8_u0_n158 ) );
  NOR2_X1 u0_u8_u0_U60 (.A2( u0_u8_X_5 ) , .ZN( u0_u8_u0_n136 ) , .A1( u0_u8_u0_n159 ) );
  NAND2_X1 u0_u8_u0_U61 (.A1( u0_u8_X_5 ) , .ZN( u0_u8_u0_n138 ) , .A2( u0_u8_u0_n159 ) );
  AND2_X1 u0_u8_u0_U62 (.A2( u0_u8_X_3 ) , .A1( u0_u8_X_6 ) , .ZN( u0_u8_u0_n102 ) );
  AND2_X1 u0_u8_u0_U63 (.A1( u0_u8_X_6 ) , .A2( u0_u8_u0_n162 ) , .ZN( u0_u8_u0_n93 ) );
  INV_X1 u0_u8_u0_U64 (.A( u0_u8_X_4 ) , .ZN( u0_u8_u0_n159 ) );
  INV_X1 u0_u8_u0_U65 (.A( u0_u8_X_2 ) , .ZN( u0_u8_u0_n163 ) );
  INV_X1 u0_u8_u0_U66 (.A( u0_u8_X_3 ) , .ZN( u0_u8_u0_n162 ) );
  INV_X1 u0_u8_u0_U67 (.A( u0_u8_u0_n126 ) , .ZN( u0_u8_u0_n168 ) );
  AOI211_X1 u0_u8_u0_U68 (.B( u0_u8_u0_n133 ) , .A( u0_u8_u0_n134 ) , .C2( u0_u8_u0_n135 ) , .C1( u0_u8_u0_n136 ) , .ZN( u0_u8_u0_n137 ) );
  OR4_X1 u0_u8_u0_U69 (.ZN( u0_out8_17 ) , .A4( u0_u8_u0_n122 ) , .A2( u0_u8_u0_n123 ) , .A1( u0_u8_u0_n124 ) , .A3( u0_u8_u0_n170 ) );
  OAI21_X1 u0_u8_u0_U7 (.B1( u0_u8_u0_n150 ) , .B2( u0_u8_u0_n158 ) , .A( u0_u8_u0_n172 ) , .ZN( u0_u8_u0_n89 ) );
  AOI21_X1 u0_u8_u0_U70 (.B2( u0_u8_u0_n107 ) , .ZN( u0_u8_u0_n124 ) , .B1( u0_u8_u0_n128 ) , .A( u0_u8_u0_n161 ) );
  INV_X1 u0_u8_u0_U71 (.A( u0_u8_u0_n111 ) , .ZN( u0_u8_u0_n170 ) );
  OR4_X1 u0_u8_u0_U72 (.ZN( u0_out8_31 ) , .A4( u0_u8_u0_n155 ) , .A2( u0_u8_u0_n156 ) , .A1( u0_u8_u0_n157 ) , .A3( u0_u8_u0_n173 ) );
  AOI21_X1 u0_u8_u0_U73 (.A( u0_u8_u0_n138 ) , .B2( u0_u8_u0_n139 ) , .B1( u0_u8_u0_n140 ) , .ZN( u0_u8_u0_n157 ) );
  AOI21_X1 u0_u8_u0_U74 (.B2( u0_u8_u0_n141 ) , .B1( u0_u8_u0_n142 ) , .ZN( u0_u8_u0_n156 ) , .A( u0_u8_u0_n161 ) );
  INV_X1 u0_u8_u0_U75 (.ZN( u0_u8_u0_n174 ) , .A( u0_u8_u0_n89 ) );
  AOI211_X1 u0_u8_u0_U76 (.B( u0_u8_u0_n104 ) , .A( u0_u8_u0_n105 ) , .ZN( u0_u8_u0_n106 ) , .C2( u0_u8_u0_n113 ) , .C1( u0_u8_u0_n160 ) );
  INV_X1 u0_u8_u0_U77 (.A( u0_u8_X_1 ) , .ZN( u0_u8_u0_n164 ) );
  NOR2_X1 u0_u8_u0_U78 (.A1( u0_u8_u0_n163 ) , .A2( u0_u8_u0_n164 ) , .ZN( u0_u8_u0_n95 ) );
  OAI221_X1 u0_u8_u0_U79 (.C1( u0_u8_u0_n121 ) , .ZN( u0_u8_u0_n122 ) , .B2( u0_u8_u0_n127 ) , .A( u0_u8_u0_n143 ) , .B1( u0_u8_u0_n144 ) , .C2( u0_u8_u0_n147 ) );
  AND2_X1 u0_u8_u0_U8 (.A1( u0_u8_u0_n114 ) , .A2( u0_u8_u0_n121 ) , .ZN( u0_u8_u0_n146 ) );
  AOI21_X1 u0_u8_u0_U80 (.B1( u0_u8_u0_n132 ) , .ZN( u0_u8_u0_n133 ) , .A( u0_u8_u0_n144 ) , .B2( u0_u8_u0_n166 ) );
  OAI22_X1 u0_u8_u0_U81 (.ZN( u0_u8_u0_n105 ) , .A2( u0_u8_u0_n132 ) , .B1( u0_u8_u0_n146 ) , .A1( u0_u8_u0_n147 ) , .B2( u0_u8_u0_n161 ) );
  NAND2_X1 u0_u8_u0_U82 (.ZN( u0_u8_u0_n110 ) , .A2( u0_u8_u0_n132 ) , .A1( u0_u8_u0_n145 ) );
  INV_X1 u0_u8_u0_U83 (.A( u0_u8_u0_n119 ) , .ZN( u0_u8_u0_n167 ) );
  NAND2_X1 u0_u8_u0_U84 (.ZN( u0_u8_u0_n148 ) , .A1( u0_u8_u0_n93 ) , .A2( u0_u8_u0_n95 ) );
  NAND2_X1 u0_u8_u0_U85 (.A1( u0_u8_u0_n100 ) , .ZN( u0_u8_u0_n129 ) , .A2( u0_u8_u0_n95 ) );
  NAND2_X1 u0_u8_u0_U86 (.A1( u0_u8_u0_n102 ) , .ZN( u0_u8_u0_n128 ) , .A2( u0_u8_u0_n95 ) );
  NAND2_X1 u0_u8_u0_U87 (.ZN( u0_u8_u0_n142 ) , .A1( u0_u8_u0_n94 ) , .A2( u0_u8_u0_n95 ) );
  NAND3_X1 u0_u8_u0_U88 (.ZN( u0_out8_23 ) , .A3( u0_u8_u0_n137 ) , .A1( u0_u8_u0_n168 ) , .A2( u0_u8_u0_n171 ) );
  NAND3_X1 u0_u8_u0_U89 (.A3( u0_u8_u0_n127 ) , .A2( u0_u8_u0_n128 ) , .ZN( u0_u8_u0_n135 ) , .A1( u0_u8_u0_n150 ) );
  AND2_X1 u0_u8_u0_U9 (.A1( u0_u8_u0_n131 ) , .ZN( u0_u8_u0_n141 ) , .A2( u0_u8_u0_n150 ) );
  NAND3_X1 u0_u8_u0_U90 (.ZN( u0_u8_u0_n117 ) , .A3( u0_u8_u0_n132 ) , .A2( u0_u8_u0_n139 ) , .A1( u0_u8_u0_n148 ) );
  NAND3_X1 u0_u8_u0_U91 (.ZN( u0_u8_u0_n109 ) , .A2( u0_u8_u0_n114 ) , .A3( u0_u8_u0_n140 ) , .A1( u0_u8_u0_n149 ) );
  NAND3_X1 u0_u8_u0_U92 (.ZN( u0_out8_9 ) , .A3( u0_u8_u0_n106 ) , .A2( u0_u8_u0_n171 ) , .A1( u0_u8_u0_n174 ) );
  NAND3_X1 u0_u8_u0_U93 (.A2( u0_u8_u0_n128 ) , .A1( u0_u8_u0_n132 ) , .A3( u0_u8_u0_n146 ) , .ZN( u0_u8_u0_n97 ) );
  AOI21_X1 u0_u8_u1_U10 (.B2( u0_u8_u1_n155 ) , .B1( u0_u8_u1_n156 ) , .ZN( u0_u8_u1_n157 ) , .A( u0_u8_u1_n174 ) );
  NAND3_X1 u0_u8_u1_U100 (.ZN( u0_u8_u1_n113 ) , .A1( u0_u8_u1_n120 ) , .A3( u0_u8_u1_n133 ) , .A2( u0_u8_u1_n155 ) );
  NAND2_X1 u0_u8_u1_U11 (.ZN( u0_u8_u1_n140 ) , .A2( u0_u8_u1_n150 ) , .A1( u0_u8_u1_n155 ) );
  NAND2_X1 u0_u8_u1_U12 (.A1( u0_u8_u1_n131 ) , .ZN( u0_u8_u1_n147 ) , .A2( u0_u8_u1_n153 ) );
  AOI22_X1 u0_u8_u1_U13 (.B2( u0_u8_u1_n136 ) , .A2( u0_u8_u1_n137 ) , .ZN( u0_u8_u1_n143 ) , .A1( u0_u8_u1_n171 ) , .B1( u0_u8_u1_n173 ) );
  INV_X1 u0_u8_u1_U14 (.A( u0_u8_u1_n147 ) , .ZN( u0_u8_u1_n181 ) );
  INV_X1 u0_u8_u1_U15 (.A( u0_u8_u1_n139 ) , .ZN( u0_u8_u1_n174 ) );
  OR4_X1 u0_u8_u1_U16 (.A4( u0_u8_u1_n106 ) , .A3( u0_u8_u1_n107 ) , .ZN( u0_u8_u1_n108 ) , .A1( u0_u8_u1_n117 ) , .A2( u0_u8_u1_n184 ) );
  AOI21_X1 u0_u8_u1_U17 (.ZN( u0_u8_u1_n106 ) , .A( u0_u8_u1_n112 ) , .B1( u0_u8_u1_n154 ) , .B2( u0_u8_u1_n156 ) );
  AOI21_X1 u0_u8_u1_U18 (.ZN( u0_u8_u1_n107 ) , .B1( u0_u8_u1_n134 ) , .B2( u0_u8_u1_n149 ) , .A( u0_u8_u1_n174 ) );
  INV_X1 u0_u8_u1_U19 (.A( u0_u8_u1_n101 ) , .ZN( u0_u8_u1_n184 ) );
  INV_X1 u0_u8_u1_U20 (.A( u0_u8_u1_n112 ) , .ZN( u0_u8_u1_n171 ) );
  NAND2_X1 u0_u8_u1_U21 (.ZN( u0_u8_u1_n141 ) , .A1( u0_u8_u1_n153 ) , .A2( u0_u8_u1_n156 ) );
  AND2_X1 u0_u8_u1_U22 (.A1( u0_u8_u1_n123 ) , .ZN( u0_u8_u1_n134 ) , .A2( u0_u8_u1_n161 ) );
  NAND2_X1 u0_u8_u1_U23 (.A2( u0_u8_u1_n115 ) , .A1( u0_u8_u1_n116 ) , .ZN( u0_u8_u1_n148 ) );
  NAND2_X1 u0_u8_u1_U24 (.A2( u0_u8_u1_n133 ) , .A1( u0_u8_u1_n135 ) , .ZN( u0_u8_u1_n159 ) );
  NAND2_X1 u0_u8_u1_U25 (.A2( u0_u8_u1_n115 ) , .A1( u0_u8_u1_n120 ) , .ZN( u0_u8_u1_n132 ) );
  INV_X1 u0_u8_u1_U26 (.A( u0_u8_u1_n154 ) , .ZN( u0_u8_u1_n178 ) );
  INV_X1 u0_u8_u1_U27 (.A( u0_u8_u1_n151 ) , .ZN( u0_u8_u1_n183 ) );
  AND2_X1 u0_u8_u1_U28 (.A1( u0_u8_u1_n129 ) , .A2( u0_u8_u1_n133 ) , .ZN( u0_u8_u1_n149 ) );
  INV_X1 u0_u8_u1_U29 (.A( u0_u8_u1_n131 ) , .ZN( u0_u8_u1_n180 ) );
  INV_X1 u0_u8_u1_U3 (.A( u0_u8_u1_n159 ) , .ZN( u0_u8_u1_n182 ) );
  AOI221_X1 u0_u8_u1_U30 (.B1( u0_u8_u1_n140 ) , .ZN( u0_u8_u1_n167 ) , .B2( u0_u8_u1_n172 ) , .C2( u0_u8_u1_n175 ) , .C1( u0_u8_u1_n178 ) , .A( u0_u8_u1_n188 ) );
  INV_X1 u0_u8_u1_U31 (.ZN( u0_u8_u1_n188 ) , .A( u0_u8_u1_n97 ) );
  AOI211_X1 u0_u8_u1_U32 (.A( u0_u8_u1_n118 ) , .C1( u0_u8_u1_n132 ) , .C2( u0_u8_u1_n139 ) , .B( u0_u8_u1_n96 ) , .ZN( u0_u8_u1_n97 ) );
  AOI21_X1 u0_u8_u1_U33 (.B2( u0_u8_u1_n121 ) , .B1( u0_u8_u1_n135 ) , .A( u0_u8_u1_n152 ) , .ZN( u0_u8_u1_n96 ) );
  OAI221_X1 u0_u8_u1_U34 (.A( u0_u8_u1_n119 ) , .C2( u0_u8_u1_n129 ) , .ZN( u0_u8_u1_n138 ) , .B2( u0_u8_u1_n152 ) , .C1( u0_u8_u1_n174 ) , .B1( u0_u8_u1_n187 ) );
  INV_X1 u0_u8_u1_U35 (.A( u0_u8_u1_n148 ) , .ZN( u0_u8_u1_n187 ) );
  AOI211_X1 u0_u8_u1_U36 (.B( u0_u8_u1_n117 ) , .A( u0_u8_u1_n118 ) , .ZN( u0_u8_u1_n119 ) , .C2( u0_u8_u1_n146 ) , .C1( u0_u8_u1_n159 ) );
  NOR2_X1 u0_u8_u1_U37 (.A1( u0_u8_u1_n168 ) , .A2( u0_u8_u1_n176 ) , .ZN( u0_u8_u1_n98 ) );
  AOI211_X1 u0_u8_u1_U38 (.B( u0_u8_u1_n162 ) , .A( u0_u8_u1_n163 ) , .C2( u0_u8_u1_n164 ) , .ZN( u0_u8_u1_n165 ) , .C1( u0_u8_u1_n171 ) );
  AOI21_X1 u0_u8_u1_U39 (.A( u0_u8_u1_n160 ) , .B2( u0_u8_u1_n161 ) , .ZN( u0_u8_u1_n162 ) , .B1( u0_u8_u1_n182 ) );
  AOI221_X1 u0_u8_u1_U4 (.A( u0_u8_u1_n138 ) , .C2( u0_u8_u1_n139 ) , .C1( u0_u8_u1_n140 ) , .B2( u0_u8_u1_n141 ) , .ZN( u0_u8_u1_n142 ) , .B1( u0_u8_u1_n175 ) );
  OR2_X1 u0_u8_u1_U40 (.A2( u0_u8_u1_n157 ) , .A1( u0_u8_u1_n158 ) , .ZN( u0_u8_u1_n163 ) );
  NAND2_X1 u0_u8_u1_U41 (.A1( u0_u8_u1_n128 ) , .ZN( u0_u8_u1_n146 ) , .A2( u0_u8_u1_n160 ) );
  NAND2_X1 u0_u8_u1_U42 (.A2( u0_u8_u1_n112 ) , .ZN( u0_u8_u1_n139 ) , .A1( u0_u8_u1_n152 ) );
  NAND2_X1 u0_u8_u1_U43 (.A1( u0_u8_u1_n105 ) , .ZN( u0_u8_u1_n156 ) , .A2( u0_u8_u1_n99 ) );
  NOR2_X1 u0_u8_u1_U44 (.ZN( u0_u8_u1_n117 ) , .A1( u0_u8_u1_n121 ) , .A2( u0_u8_u1_n160 ) );
  OAI21_X1 u0_u8_u1_U45 (.B2( u0_u8_u1_n123 ) , .ZN( u0_u8_u1_n145 ) , .B1( u0_u8_u1_n160 ) , .A( u0_u8_u1_n185 ) );
  INV_X1 u0_u8_u1_U46 (.A( u0_u8_u1_n122 ) , .ZN( u0_u8_u1_n185 ) );
  AOI21_X1 u0_u8_u1_U47 (.B2( u0_u8_u1_n120 ) , .B1( u0_u8_u1_n121 ) , .ZN( u0_u8_u1_n122 ) , .A( u0_u8_u1_n128 ) );
  AOI21_X1 u0_u8_u1_U48 (.A( u0_u8_u1_n128 ) , .B2( u0_u8_u1_n129 ) , .ZN( u0_u8_u1_n130 ) , .B1( u0_u8_u1_n150 ) );
  NAND2_X1 u0_u8_u1_U49 (.ZN( u0_u8_u1_n112 ) , .A1( u0_u8_u1_n169 ) , .A2( u0_u8_u1_n170 ) );
  AOI211_X1 u0_u8_u1_U5 (.ZN( u0_u8_u1_n124 ) , .A( u0_u8_u1_n138 ) , .C2( u0_u8_u1_n139 ) , .B( u0_u8_u1_n145 ) , .C1( u0_u8_u1_n147 ) );
  NAND2_X1 u0_u8_u1_U50 (.ZN( u0_u8_u1_n129 ) , .A2( u0_u8_u1_n95 ) , .A1( u0_u8_u1_n98 ) );
  NAND2_X1 u0_u8_u1_U51 (.A1( u0_u8_u1_n102 ) , .ZN( u0_u8_u1_n154 ) , .A2( u0_u8_u1_n99 ) );
  NAND2_X1 u0_u8_u1_U52 (.A2( u0_u8_u1_n100 ) , .ZN( u0_u8_u1_n135 ) , .A1( u0_u8_u1_n99 ) );
  AOI21_X1 u0_u8_u1_U53 (.A( u0_u8_u1_n152 ) , .B2( u0_u8_u1_n153 ) , .B1( u0_u8_u1_n154 ) , .ZN( u0_u8_u1_n158 ) );
  INV_X1 u0_u8_u1_U54 (.A( u0_u8_u1_n160 ) , .ZN( u0_u8_u1_n175 ) );
  NAND2_X1 u0_u8_u1_U55 (.A1( u0_u8_u1_n100 ) , .ZN( u0_u8_u1_n116 ) , .A2( u0_u8_u1_n95 ) );
  NAND2_X1 u0_u8_u1_U56 (.A1( u0_u8_u1_n102 ) , .ZN( u0_u8_u1_n131 ) , .A2( u0_u8_u1_n95 ) );
  NAND2_X1 u0_u8_u1_U57 (.A2( u0_u8_u1_n104 ) , .ZN( u0_u8_u1_n121 ) , .A1( u0_u8_u1_n98 ) );
  NAND2_X1 u0_u8_u1_U58 (.A1( u0_u8_u1_n103 ) , .ZN( u0_u8_u1_n153 ) , .A2( u0_u8_u1_n98 ) );
  NAND2_X1 u0_u8_u1_U59 (.A2( u0_u8_u1_n104 ) , .A1( u0_u8_u1_n105 ) , .ZN( u0_u8_u1_n133 ) );
  AOI22_X1 u0_u8_u1_U6 (.B2( u0_u8_u1_n113 ) , .A2( u0_u8_u1_n114 ) , .ZN( u0_u8_u1_n125 ) , .A1( u0_u8_u1_n171 ) , .B1( u0_u8_u1_n173 ) );
  NAND2_X1 u0_u8_u1_U60 (.ZN( u0_u8_u1_n150 ) , .A2( u0_u8_u1_n98 ) , .A1( u0_u8_u1_n99 ) );
  NAND2_X1 u0_u8_u1_U61 (.A1( u0_u8_u1_n105 ) , .ZN( u0_u8_u1_n155 ) , .A2( u0_u8_u1_n95 ) );
  OAI21_X1 u0_u8_u1_U62 (.ZN( u0_u8_u1_n109 ) , .B1( u0_u8_u1_n129 ) , .B2( u0_u8_u1_n160 ) , .A( u0_u8_u1_n167 ) );
  NAND2_X1 u0_u8_u1_U63 (.A2( u0_u8_u1_n100 ) , .A1( u0_u8_u1_n103 ) , .ZN( u0_u8_u1_n120 ) );
  NAND2_X1 u0_u8_u1_U64 (.A1( u0_u8_u1_n102 ) , .A2( u0_u8_u1_n104 ) , .ZN( u0_u8_u1_n115 ) );
  NAND2_X1 u0_u8_u1_U65 (.A2( u0_u8_u1_n100 ) , .A1( u0_u8_u1_n104 ) , .ZN( u0_u8_u1_n151 ) );
  NAND2_X1 u0_u8_u1_U66 (.A2( u0_u8_u1_n103 ) , .A1( u0_u8_u1_n105 ) , .ZN( u0_u8_u1_n161 ) );
  INV_X1 u0_u8_u1_U67 (.A( u0_u8_u1_n152 ) , .ZN( u0_u8_u1_n173 ) );
  INV_X1 u0_u8_u1_U68 (.A( u0_u8_u1_n128 ) , .ZN( u0_u8_u1_n172 ) );
  NAND2_X1 u0_u8_u1_U69 (.A2( u0_u8_u1_n102 ) , .A1( u0_u8_u1_n103 ) , .ZN( u0_u8_u1_n123 ) );
  NAND2_X1 u0_u8_u1_U7 (.ZN( u0_u8_u1_n114 ) , .A1( u0_u8_u1_n134 ) , .A2( u0_u8_u1_n156 ) );
  NOR2_X1 u0_u8_u1_U70 (.A2( u0_u8_X_7 ) , .A1( u0_u8_X_8 ) , .ZN( u0_u8_u1_n95 ) );
  NOR2_X1 u0_u8_u1_U71 (.A1( u0_u8_X_12 ) , .A2( u0_u8_X_9 ) , .ZN( u0_u8_u1_n100 ) );
  NOR2_X1 u0_u8_u1_U72 (.A2( u0_u8_X_8 ) , .A1( u0_u8_u1_n177 ) , .ZN( u0_u8_u1_n99 ) );
  NOR2_X1 u0_u8_u1_U73 (.A2( u0_u8_X_12 ) , .ZN( u0_u8_u1_n102 ) , .A1( u0_u8_u1_n176 ) );
  NOR2_X1 u0_u8_u1_U74 (.A2( u0_u8_X_9 ) , .ZN( u0_u8_u1_n105 ) , .A1( u0_u8_u1_n168 ) );
  NAND2_X1 u0_u8_u1_U75 (.A1( u0_u8_X_10 ) , .ZN( u0_u8_u1_n160 ) , .A2( u0_u8_u1_n169 ) );
  NAND2_X1 u0_u8_u1_U76 (.A2( u0_u8_X_10 ) , .A1( u0_u8_X_11 ) , .ZN( u0_u8_u1_n152 ) );
  NAND2_X1 u0_u8_u1_U77 (.A1( u0_u8_X_11 ) , .ZN( u0_u8_u1_n128 ) , .A2( u0_u8_u1_n170 ) );
  AND2_X1 u0_u8_u1_U78 (.A2( u0_u8_X_7 ) , .A1( u0_u8_X_8 ) , .ZN( u0_u8_u1_n104 ) );
  AND2_X1 u0_u8_u1_U79 (.A1( u0_u8_X_8 ) , .ZN( u0_u8_u1_n103 ) , .A2( u0_u8_u1_n177 ) );
  NOR2_X1 u0_u8_u1_U8 (.A1( u0_u8_u1_n112 ) , .A2( u0_u8_u1_n116 ) , .ZN( u0_u8_u1_n118 ) );
  INV_X1 u0_u8_u1_U80 (.A( u0_u8_X_10 ) , .ZN( u0_u8_u1_n170 ) );
  INV_X1 u0_u8_u1_U81 (.A( u0_u8_X_9 ) , .ZN( u0_u8_u1_n176 ) );
  INV_X1 u0_u8_u1_U82 (.A( u0_u8_X_11 ) , .ZN( u0_u8_u1_n169 ) );
  INV_X1 u0_u8_u1_U83 (.A( u0_u8_X_12 ) , .ZN( u0_u8_u1_n168 ) );
  INV_X1 u0_u8_u1_U84 (.A( u0_u8_X_7 ) , .ZN( u0_u8_u1_n177 ) );
  NAND4_X1 u0_u8_u1_U85 (.ZN( u0_out8_28 ) , .A4( u0_u8_u1_n124 ) , .A3( u0_u8_u1_n125 ) , .A2( u0_u8_u1_n126 ) , .A1( u0_u8_u1_n127 ) );
  OAI21_X1 u0_u8_u1_U86 (.ZN( u0_u8_u1_n127 ) , .B2( u0_u8_u1_n139 ) , .B1( u0_u8_u1_n175 ) , .A( u0_u8_u1_n183 ) );
  OAI21_X1 u0_u8_u1_U87 (.ZN( u0_u8_u1_n126 ) , .B2( u0_u8_u1_n140 ) , .A( u0_u8_u1_n146 ) , .B1( u0_u8_u1_n178 ) );
  NAND4_X1 u0_u8_u1_U88 (.ZN( u0_out8_18 ) , .A4( u0_u8_u1_n165 ) , .A3( u0_u8_u1_n166 ) , .A1( u0_u8_u1_n167 ) , .A2( u0_u8_u1_n186 ) );
  AOI22_X1 u0_u8_u1_U89 (.B2( u0_u8_u1_n146 ) , .B1( u0_u8_u1_n147 ) , .A2( u0_u8_u1_n148 ) , .ZN( u0_u8_u1_n166 ) , .A1( u0_u8_u1_n172 ) );
  OAI21_X1 u0_u8_u1_U9 (.ZN( u0_u8_u1_n101 ) , .B1( u0_u8_u1_n141 ) , .A( u0_u8_u1_n146 ) , .B2( u0_u8_u1_n183 ) );
  INV_X1 u0_u8_u1_U90 (.A( u0_u8_u1_n145 ) , .ZN( u0_u8_u1_n186 ) );
  NAND4_X1 u0_u8_u1_U91 (.ZN( u0_out8_2 ) , .A4( u0_u8_u1_n142 ) , .A3( u0_u8_u1_n143 ) , .A2( u0_u8_u1_n144 ) , .A1( u0_u8_u1_n179 ) );
  OAI21_X1 u0_u8_u1_U92 (.B2( u0_u8_u1_n132 ) , .ZN( u0_u8_u1_n144 ) , .A( u0_u8_u1_n146 ) , .B1( u0_u8_u1_n180 ) );
  INV_X1 u0_u8_u1_U93 (.A( u0_u8_u1_n130 ) , .ZN( u0_u8_u1_n179 ) );
  OR4_X1 u0_u8_u1_U94 (.ZN( u0_out8_13 ) , .A4( u0_u8_u1_n108 ) , .A3( u0_u8_u1_n109 ) , .A2( u0_u8_u1_n110 ) , .A1( u0_u8_u1_n111 ) );
  AOI21_X1 u0_u8_u1_U95 (.ZN( u0_u8_u1_n111 ) , .A( u0_u8_u1_n128 ) , .B2( u0_u8_u1_n131 ) , .B1( u0_u8_u1_n135 ) );
  AOI21_X1 u0_u8_u1_U96 (.ZN( u0_u8_u1_n110 ) , .A( u0_u8_u1_n116 ) , .B1( u0_u8_u1_n152 ) , .B2( u0_u8_u1_n160 ) );
  NAND3_X1 u0_u8_u1_U97 (.A3( u0_u8_u1_n149 ) , .A2( u0_u8_u1_n150 ) , .A1( u0_u8_u1_n151 ) , .ZN( u0_u8_u1_n164 ) );
  NAND3_X1 u0_u8_u1_U98 (.A3( u0_u8_u1_n134 ) , .A2( u0_u8_u1_n135 ) , .ZN( u0_u8_u1_n136 ) , .A1( u0_u8_u1_n151 ) );
  NAND3_X1 u0_u8_u1_U99 (.A1( u0_u8_u1_n133 ) , .ZN( u0_u8_u1_n137 ) , .A2( u0_u8_u1_n154 ) , .A3( u0_u8_u1_n181 ) );
  OAI22_X1 u0_u8_u2_U10 (.B1( u0_u8_u2_n151 ) , .A2( u0_u8_u2_n152 ) , .A1( u0_u8_u2_n153 ) , .ZN( u0_u8_u2_n160 ) , .B2( u0_u8_u2_n168 ) );
  NAND3_X1 u0_u8_u2_U100 (.A2( u0_u8_u2_n100 ) , .A1( u0_u8_u2_n104 ) , .A3( u0_u8_u2_n138 ) , .ZN( u0_u8_u2_n98 ) );
  NOR3_X1 u0_u8_u2_U11 (.A1( u0_u8_u2_n150 ) , .ZN( u0_u8_u2_n151 ) , .A3( u0_u8_u2_n175 ) , .A2( u0_u8_u2_n188 ) );
  AOI21_X1 u0_u8_u2_U12 (.B2( u0_u8_u2_n123 ) , .ZN( u0_u8_u2_n125 ) , .A( u0_u8_u2_n171 ) , .B1( u0_u8_u2_n184 ) );
  INV_X1 u0_u8_u2_U13 (.A( u0_u8_u2_n150 ) , .ZN( u0_u8_u2_n184 ) );
  AOI21_X1 u0_u8_u2_U14 (.ZN( u0_u8_u2_n144 ) , .B2( u0_u8_u2_n155 ) , .A( u0_u8_u2_n172 ) , .B1( u0_u8_u2_n185 ) );
  AOI21_X1 u0_u8_u2_U15 (.B2( u0_u8_u2_n143 ) , .ZN( u0_u8_u2_n145 ) , .B1( u0_u8_u2_n152 ) , .A( u0_u8_u2_n171 ) );
  INV_X1 u0_u8_u2_U16 (.A( u0_u8_u2_n156 ) , .ZN( u0_u8_u2_n171 ) );
  INV_X1 u0_u8_u2_U17 (.A( u0_u8_u2_n120 ) , .ZN( u0_u8_u2_n188 ) );
  NAND2_X1 u0_u8_u2_U18 (.A2( u0_u8_u2_n122 ) , .ZN( u0_u8_u2_n150 ) , .A1( u0_u8_u2_n152 ) );
  INV_X1 u0_u8_u2_U19 (.A( u0_u8_u2_n153 ) , .ZN( u0_u8_u2_n170 ) );
  INV_X1 u0_u8_u2_U20 (.A( u0_u8_u2_n137 ) , .ZN( u0_u8_u2_n173 ) );
  NAND2_X1 u0_u8_u2_U21 (.A1( u0_u8_u2_n132 ) , .A2( u0_u8_u2_n139 ) , .ZN( u0_u8_u2_n157 ) );
  INV_X1 u0_u8_u2_U22 (.A( u0_u8_u2_n113 ) , .ZN( u0_u8_u2_n178 ) );
  INV_X1 u0_u8_u2_U23 (.A( u0_u8_u2_n139 ) , .ZN( u0_u8_u2_n175 ) );
  INV_X1 u0_u8_u2_U24 (.A( u0_u8_u2_n155 ) , .ZN( u0_u8_u2_n181 ) );
  INV_X1 u0_u8_u2_U25 (.A( u0_u8_u2_n119 ) , .ZN( u0_u8_u2_n177 ) );
  INV_X1 u0_u8_u2_U26 (.A( u0_u8_u2_n116 ) , .ZN( u0_u8_u2_n180 ) );
  INV_X1 u0_u8_u2_U27 (.A( u0_u8_u2_n131 ) , .ZN( u0_u8_u2_n179 ) );
  INV_X1 u0_u8_u2_U28 (.A( u0_u8_u2_n154 ) , .ZN( u0_u8_u2_n176 ) );
  NAND2_X1 u0_u8_u2_U29 (.A2( u0_u8_u2_n116 ) , .A1( u0_u8_u2_n117 ) , .ZN( u0_u8_u2_n118 ) );
  NOR2_X1 u0_u8_u2_U3 (.ZN( u0_u8_u2_n121 ) , .A2( u0_u8_u2_n177 ) , .A1( u0_u8_u2_n180 ) );
  INV_X1 u0_u8_u2_U30 (.A( u0_u8_u2_n132 ) , .ZN( u0_u8_u2_n182 ) );
  INV_X1 u0_u8_u2_U31 (.A( u0_u8_u2_n158 ) , .ZN( u0_u8_u2_n183 ) );
  OAI21_X1 u0_u8_u2_U32 (.A( u0_u8_u2_n156 ) , .B1( u0_u8_u2_n157 ) , .ZN( u0_u8_u2_n158 ) , .B2( u0_u8_u2_n179 ) );
  NOR2_X1 u0_u8_u2_U33 (.ZN( u0_u8_u2_n156 ) , .A1( u0_u8_u2_n166 ) , .A2( u0_u8_u2_n169 ) );
  NOR2_X1 u0_u8_u2_U34 (.A2( u0_u8_u2_n114 ) , .ZN( u0_u8_u2_n137 ) , .A1( u0_u8_u2_n140 ) );
  NOR2_X1 u0_u8_u2_U35 (.A2( u0_u8_u2_n138 ) , .ZN( u0_u8_u2_n153 ) , .A1( u0_u8_u2_n156 ) );
  AOI211_X1 u0_u8_u2_U36 (.ZN( u0_u8_u2_n130 ) , .C1( u0_u8_u2_n138 ) , .C2( u0_u8_u2_n179 ) , .B( u0_u8_u2_n96 ) , .A( u0_u8_u2_n97 ) );
  OAI22_X1 u0_u8_u2_U37 (.B1( u0_u8_u2_n133 ) , .A2( u0_u8_u2_n137 ) , .A1( u0_u8_u2_n152 ) , .B2( u0_u8_u2_n168 ) , .ZN( u0_u8_u2_n97 ) );
  OAI221_X1 u0_u8_u2_U38 (.B1( u0_u8_u2_n113 ) , .C1( u0_u8_u2_n132 ) , .A( u0_u8_u2_n149 ) , .B2( u0_u8_u2_n171 ) , .C2( u0_u8_u2_n172 ) , .ZN( u0_u8_u2_n96 ) );
  OAI221_X1 u0_u8_u2_U39 (.A( u0_u8_u2_n115 ) , .C2( u0_u8_u2_n123 ) , .B2( u0_u8_u2_n143 ) , .B1( u0_u8_u2_n153 ) , .ZN( u0_u8_u2_n163 ) , .C1( u0_u8_u2_n168 ) );
  INV_X1 u0_u8_u2_U4 (.A( u0_u8_u2_n134 ) , .ZN( u0_u8_u2_n185 ) );
  OAI21_X1 u0_u8_u2_U40 (.A( u0_u8_u2_n114 ) , .ZN( u0_u8_u2_n115 ) , .B1( u0_u8_u2_n176 ) , .B2( u0_u8_u2_n178 ) );
  OAI221_X1 u0_u8_u2_U41 (.A( u0_u8_u2_n135 ) , .B2( u0_u8_u2_n136 ) , .B1( u0_u8_u2_n137 ) , .ZN( u0_u8_u2_n162 ) , .C2( u0_u8_u2_n167 ) , .C1( u0_u8_u2_n185 ) );
  AND3_X1 u0_u8_u2_U42 (.A3( u0_u8_u2_n131 ) , .A2( u0_u8_u2_n132 ) , .A1( u0_u8_u2_n133 ) , .ZN( u0_u8_u2_n136 ) );
  AOI22_X1 u0_u8_u2_U43 (.ZN( u0_u8_u2_n135 ) , .B1( u0_u8_u2_n140 ) , .A1( u0_u8_u2_n156 ) , .B2( u0_u8_u2_n180 ) , .A2( u0_u8_u2_n188 ) );
  AOI21_X1 u0_u8_u2_U44 (.ZN( u0_u8_u2_n149 ) , .B1( u0_u8_u2_n173 ) , .B2( u0_u8_u2_n188 ) , .A( u0_u8_u2_n95 ) );
  AND3_X1 u0_u8_u2_U45 (.A2( u0_u8_u2_n100 ) , .A1( u0_u8_u2_n104 ) , .A3( u0_u8_u2_n156 ) , .ZN( u0_u8_u2_n95 ) );
  OAI21_X1 u0_u8_u2_U46 (.A( u0_u8_u2_n141 ) , .B2( u0_u8_u2_n142 ) , .ZN( u0_u8_u2_n146 ) , .B1( u0_u8_u2_n153 ) );
  OAI21_X1 u0_u8_u2_U47 (.A( u0_u8_u2_n140 ) , .ZN( u0_u8_u2_n141 ) , .B1( u0_u8_u2_n176 ) , .B2( u0_u8_u2_n177 ) );
  NOR3_X1 u0_u8_u2_U48 (.ZN( u0_u8_u2_n142 ) , .A3( u0_u8_u2_n175 ) , .A2( u0_u8_u2_n178 ) , .A1( u0_u8_u2_n181 ) );
  OAI21_X1 u0_u8_u2_U49 (.A( u0_u8_u2_n101 ) , .B2( u0_u8_u2_n121 ) , .B1( u0_u8_u2_n153 ) , .ZN( u0_u8_u2_n164 ) );
  NOR4_X1 u0_u8_u2_U5 (.A4( u0_u8_u2_n124 ) , .A3( u0_u8_u2_n125 ) , .A2( u0_u8_u2_n126 ) , .A1( u0_u8_u2_n127 ) , .ZN( u0_u8_u2_n128 ) );
  NAND2_X1 u0_u8_u2_U50 (.A2( u0_u8_u2_n100 ) , .A1( u0_u8_u2_n107 ) , .ZN( u0_u8_u2_n155 ) );
  NAND2_X1 u0_u8_u2_U51 (.A2( u0_u8_u2_n105 ) , .A1( u0_u8_u2_n108 ) , .ZN( u0_u8_u2_n143 ) );
  NAND2_X1 u0_u8_u2_U52 (.A1( u0_u8_u2_n104 ) , .A2( u0_u8_u2_n106 ) , .ZN( u0_u8_u2_n152 ) );
  NAND2_X1 u0_u8_u2_U53 (.A1( u0_u8_u2_n100 ) , .A2( u0_u8_u2_n105 ) , .ZN( u0_u8_u2_n132 ) );
  INV_X1 u0_u8_u2_U54 (.A( u0_u8_u2_n140 ) , .ZN( u0_u8_u2_n168 ) );
  INV_X1 u0_u8_u2_U55 (.A( u0_u8_u2_n138 ) , .ZN( u0_u8_u2_n167 ) );
  NAND2_X1 u0_u8_u2_U56 (.A1( u0_u8_u2_n102 ) , .A2( u0_u8_u2_n106 ) , .ZN( u0_u8_u2_n113 ) );
  NAND2_X1 u0_u8_u2_U57 (.A1( u0_u8_u2_n106 ) , .A2( u0_u8_u2_n107 ) , .ZN( u0_u8_u2_n131 ) );
  NAND2_X1 u0_u8_u2_U58 (.A1( u0_u8_u2_n103 ) , .A2( u0_u8_u2_n107 ) , .ZN( u0_u8_u2_n139 ) );
  NAND2_X1 u0_u8_u2_U59 (.A1( u0_u8_u2_n103 ) , .A2( u0_u8_u2_n105 ) , .ZN( u0_u8_u2_n133 ) );
  AOI21_X1 u0_u8_u2_U6 (.B2( u0_u8_u2_n119 ) , .ZN( u0_u8_u2_n127 ) , .A( u0_u8_u2_n137 ) , .B1( u0_u8_u2_n155 ) );
  NAND2_X1 u0_u8_u2_U60 (.A1( u0_u8_u2_n102 ) , .A2( u0_u8_u2_n103 ) , .ZN( u0_u8_u2_n154 ) );
  NAND2_X1 u0_u8_u2_U61 (.A2( u0_u8_u2_n103 ) , .A1( u0_u8_u2_n104 ) , .ZN( u0_u8_u2_n119 ) );
  NAND2_X1 u0_u8_u2_U62 (.A2( u0_u8_u2_n107 ) , .A1( u0_u8_u2_n108 ) , .ZN( u0_u8_u2_n123 ) );
  NAND2_X1 u0_u8_u2_U63 (.A1( u0_u8_u2_n104 ) , .A2( u0_u8_u2_n108 ) , .ZN( u0_u8_u2_n122 ) );
  INV_X1 u0_u8_u2_U64 (.A( u0_u8_u2_n114 ) , .ZN( u0_u8_u2_n172 ) );
  NAND2_X1 u0_u8_u2_U65 (.A2( u0_u8_u2_n100 ) , .A1( u0_u8_u2_n102 ) , .ZN( u0_u8_u2_n116 ) );
  NAND2_X1 u0_u8_u2_U66 (.A1( u0_u8_u2_n102 ) , .A2( u0_u8_u2_n108 ) , .ZN( u0_u8_u2_n120 ) );
  NAND2_X1 u0_u8_u2_U67 (.A2( u0_u8_u2_n105 ) , .A1( u0_u8_u2_n106 ) , .ZN( u0_u8_u2_n117 ) );
  INV_X1 u0_u8_u2_U68 (.ZN( u0_u8_u2_n187 ) , .A( u0_u8_u2_n99 ) );
  OAI21_X1 u0_u8_u2_U69 (.B1( u0_u8_u2_n137 ) , .B2( u0_u8_u2_n143 ) , .A( u0_u8_u2_n98 ) , .ZN( u0_u8_u2_n99 ) );
  AOI21_X1 u0_u8_u2_U7 (.ZN( u0_u8_u2_n124 ) , .B1( u0_u8_u2_n131 ) , .B2( u0_u8_u2_n143 ) , .A( u0_u8_u2_n172 ) );
  NOR2_X1 u0_u8_u2_U70 (.A2( u0_u8_X_16 ) , .ZN( u0_u8_u2_n140 ) , .A1( u0_u8_u2_n166 ) );
  NOR2_X1 u0_u8_u2_U71 (.A2( u0_u8_X_13 ) , .A1( u0_u8_X_14 ) , .ZN( u0_u8_u2_n100 ) );
  NOR2_X1 u0_u8_u2_U72 (.A2( u0_u8_X_16 ) , .A1( u0_u8_X_17 ) , .ZN( u0_u8_u2_n138 ) );
  NOR2_X1 u0_u8_u2_U73 (.A2( u0_u8_X_15 ) , .A1( u0_u8_X_18 ) , .ZN( u0_u8_u2_n104 ) );
  NOR2_X1 u0_u8_u2_U74 (.A2( u0_u8_X_14 ) , .ZN( u0_u8_u2_n103 ) , .A1( u0_u8_u2_n174 ) );
  NOR2_X1 u0_u8_u2_U75 (.A2( u0_u8_X_15 ) , .ZN( u0_u8_u2_n102 ) , .A1( u0_u8_u2_n165 ) );
  NOR2_X1 u0_u8_u2_U76 (.A2( u0_u8_X_17 ) , .ZN( u0_u8_u2_n114 ) , .A1( u0_u8_u2_n169 ) );
  AND2_X1 u0_u8_u2_U77 (.A1( u0_u8_X_15 ) , .ZN( u0_u8_u2_n105 ) , .A2( u0_u8_u2_n165 ) );
  AND2_X1 u0_u8_u2_U78 (.A2( u0_u8_X_15 ) , .A1( u0_u8_X_18 ) , .ZN( u0_u8_u2_n107 ) );
  AND2_X1 u0_u8_u2_U79 (.A1( u0_u8_X_14 ) , .ZN( u0_u8_u2_n106 ) , .A2( u0_u8_u2_n174 ) );
  AOI21_X1 u0_u8_u2_U8 (.B2( u0_u8_u2_n120 ) , .B1( u0_u8_u2_n121 ) , .ZN( u0_u8_u2_n126 ) , .A( u0_u8_u2_n167 ) );
  AND2_X1 u0_u8_u2_U80 (.A1( u0_u8_X_13 ) , .A2( u0_u8_X_14 ) , .ZN( u0_u8_u2_n108 ) );
  INV_X1 u0_u8_u2_U81 (.A( u0_u8_X_16 ) , .ZN( u0_u8_u2_n169 ) );
  INV_X1 u0_u8_u2_U82 (.A( u0_u8_X_17 ) , .ZN( u0_u8_u2_n166 ) );
  INV_X1 u0_u8_u2_U83 (.A( u0_u8_X_13 ) , .ZN( u0_u8_u2_n174 ) );
  INV_X1 u0_u8_u2_U84 (.A( u0_u8_X_18 ) , .ZN( u0_u8_u2_n165 ) );
  NAND4_X1 u0_u8_u2_U85 (.ZN( u0_out8_30 ) , .A4( u0_u8_u2_n147 ) , .A3( u0_u8_u2_n148 ) , .A2( u0_u8_u2_n149 ) , .A1( u0_u8_u2_n187 ) );
  NOR3_X1 u0_u8_u2_U86 (.A3( u0_u8_u2_n144 ) , .A2( u0_u8_u2_n145 ) , .A1( u0_u8_u2_n146 ) , .ZN( u0_u8_u2_n147 ) );
  AOI21_X1 u0_u8_u2_U87 (.B2( u0_u8_u2_n138 ) , .ZN( u0_u8_u2_n148 ) , .A( u0_u8_u2_n162 ) , .B1( u0_u8_u2_n182 ) );
  NAND4_X1 u0_u8_u2_U88 (.ZN( u0_out8_24 ) , .A4( u0_u8_u2_n111 ) , .A3( u0_u8_u2_n112 ) , .A1( u0_u8_u2_n130 ) , .A2( u0_u8_u2_n187 ) );
  AOI221_X1 u0_u8_u2_U89 (.A( u0_u8_u2_n109 ) , .B1( u0_u8_u2_n110 ) , .ZN( u0_u8_u2_n111 ) , .C1( u0_u8_u2_n134 ) , .C2( u0_u8_u2_n170 ) , .B2( u0_u8_u2_n173 ) );
  OAI22_X1 u0_u8_u2_U9 (.ZN( u0_u8_u2_n109 ) , .A2( u0_u8_u2_n113 ) , .B2( u0_u8_u2_n133 ) , .B1( u0_u8_u2_n167 ) , .A1( u0_u8_u2_n168 ) );
  AOI21_X1 u0_u8_u2_U90 (.ZN( u0_u8_u2_n112 ) , .B2( u0_u8_u2_n156 ) , .A( u0_u8_u2_n164 ) , .B1( u0_u8_u2_n181 ) );
  NAND4_X1 u0_u8_u2_U91 (.ZN( u0_out8_16 ) , .A4( u0_u8_u2_n128 ) , .A3( u0_u8_u2_n129 ) , .A1( u0_u8_u2_n130 ) , .A2( u0_u8_u2_n186 ) );
  AOI22_X1 u0_u8_u2_U92 (.A2( u0_u8_u2_n118 ) , .ZN( u0_u8_u2_n129 ) , .A1( u0_u8_u2_n140 ) , .B1( u0_u8_u2_n157 ) , .B2( u0_u8_u2_n170 ) );
  INV_X1 u0_u8_u2_U93 (.A( u0_u8_u2_n163 ) , .ZN( u0_u8_u2_n186 ) );
  OR4_X1 u0_u8_u2_U94 (.ZN( u0_out8_6 ) , .A4( u0_u8_u2_n161 ) , .A3( u0_u8_u2_n162 ) , .A2( u0_u8_u2_n163 ) , .A1( u0_u8_u2_n164 ) );
  OR3_X1 u0_u8_u2_U95 (.A2( u0_u8_u2_n159 ) , .A1( u0_u8_u2_n160 ) , .ZN( u0_u8_u2_n161 ) , .A3( u0_u8_u2_n183 ) );
  AOI21_X1 u0_u8_u2_U96 (.B2( u0_u8_u2_n154 ) , .B1( u0_u8_u2_n155 ) , .ZN( u0_u8_u2_n159 ) , .A( u0_u8_u2_n167 ) );
  NAND3_X1 u0_u8_u2_U97 (.A2( u0_u8_u2_n117 ) , .A1( u0_u8_u2_n122 ) , .A3( u0_u8_u2_n123 ) , .ZN( u0_u8_u2_n134 ) );
  NAND3_X1 u0_u8_u2_U98 (.ZN( u0_u8_u2_n110 ) , .A2( u0_u8_u2_n131 ) , .A3( u0_u8_u2_n139 ) , .A1( u0_u8_u2_n154 ) );
  NAND3_X1 u0_u8_u2_U99 (.A2( u0_u8_u2_n100 ) , .ZN( u0_u8_u2_n101 ) , .A1( u0_u8_u2_n104 ) , .A3( u0_u8_u2_n114 ) );
  NOR2_X1 u0_u8_u5_U10 (.ZN( u0_u8_u5_n135 ) , .A1( u0_u8_u5_n173 ) , .A2( u0_u8_u5_n176 ) );
  NOR3_X1 u0_u8_u5_U100 (.A3( u0_u8_u5_n141 ) , .A1( u0_u8_u5_n142 ) , .ZN( u0_u8_u5_n143 ) , .A2( u0_u8_u5_n191 ) );
  NAND4_X1 u0_u8_u5_U101 (.ZN( u0_out8_4 ) , .A4( u0_u8_u5_n112 ) , .A2( u0_u8_u5_n113 ) , .A1( u0_u8_u5_n114 ) , .A3( u0_u8_u5_n195 ) );
  AOI211_X1 u0_u8_u5_U102 (.A( u0_u8_u5_n110 ) , .C1( u0_u8_u5_n111 ) , .ZN( u0_u8_u5_n112 ) , .B( u0_u8_u5_n118 ) , .C2( u0_u8_u5_n177 ) );
  INV_X1 u0_u8_u5_U103 (.A( u0_u8_u5_n102 ) , .ZN( u0_u8_u5_n195 ) );
  NAND3_X1 u0_u8_u5_U104 (.A2( u0_u8_u5_n154 ) , .A3( u0_u8_u5_n158 ) , .A1( u0_u8_u5_n161 ) , .ZN( u0_u8_u5_n99 ) );
  INV_X1 u0_u8_u5_U11 (.A( u0_u8_u5_n121 ) , .ZN( u0_u8_u5_n177 ) );
  NOR2_X1 u0_u8_u5_U12 (.ZN( u0_u8_u5_n160 ) , .A2( u0_u8_u5_n173 ) , .A1( u0_u8_u5_n177 ) );
  INV_X1 u0_u8_u5_U13 (.A( u0_u8_u5_n150 ) , .ZN( u0_u8_u5_n174 ) );
  AOI21_X1 u0_u8_u5_U14 (.A( u0_u8_u5_n160 ) , .B2( u0_u8_u5_n161 ) , .ZN( u0_u8_u5_n162 ) , .B1( u0_u8_u5_n192 ) );
  INV_X1 u0_u8_u5_U15 (.A( u0_u8_u5_n159 ) , .ZN( u0_u8_u5_n192 ) );
  AOI21_X1 u0_u8_u5_U16 (.A( u0_u8_u5_n156 ) , .B2( u0_u8_u5_n157 ) , .B1( u0_u8_u5_n158 ) , .ZN( u0_u8_u5_n163 ) );
  AOI21_X1 u0_u8_u5_U17 (.B2( u0_u8_u5_n139 ) , .B1( u0_u8_u5_n140 ) , .ZN( u0_u8_u5_n141 ) , .A( u0_u8_u5_n150 ) );
  OAI21_X1 u0_u8_u5_U18 (.A( u0_u8_u5_n133 ) , .B2( u0_u8_u5_n134 ) , .B1( u0_u8_u5_n135 ) , .ZN( u0_u8_u5_n142 ) );
  OAI21_X1 u0_u8_u5_U19 (.ZN( u0_u8_u5_n133 ) , .B2( u0_u8_u5_n147 ) , .A( u0_u8_u5_n173 ) , .B1( u0_u8_u5_n188 ) );
  NAND2_X1 u0_u8_u5_U20 (.A2( u0_u8_u5_n119 ) , .A1( u0_u8_u5_n123 ) , .ZN( u0_u8_u5_n137 ) );
  INV_X1 u0_u8_u5_U21 (.A( u0_u8_u5_n155 ) , .ZN( u0_u8_u5_n194 ) );
  NAND2_X1 u0_u8_u5_U22 (.A1( u0_u8_u5_n121 ) , .ZN( u0_u8_u5_n132 ) , .A2( u0_u8_u5_n172 ) );
  NAND2_X1 u0_u8_u5_U23 (.A2( u0_u8_u5_n122 ) , .ZN( u0_u8_u5_n136 ) , .A1( u0_u8_u5_n154 ) );
  NAND2_X1 u0_u8_u5_U24 (.A2( u0_u8_u5_n119 ) , .A1( u0_u8_u5_n120 ) , .ZN( u0_u8_u5_n159 ) );
  INV_X1 u0_u8_u5_U25 (.A( u0_u8_u5_n156 ) , .ZN( u0_u8_u5_n175 ) );
  INV_X1 u0_u8_u5_U26 (.A( u0_u8_u5_n158 ) , .ZN( u0_u8_u5_n188 ) );
  INV_X1 u0_u8_u5_U27 (.A( u0_u8_u5_n152 ) , .ZN( u0_u8_u5_n179 ) );
  INV_X1 u0_u8_u5_U28 (.A( u0_u8_u5_n140 ) , .ZN( u0_u8_u5_n182 ) );
  INV_X1 u0_u8_u5_U29 (.A( u0_u8_u5_n151 ) , .ZN( u0_u8_u5_n183 ) );
  NOR2_X1 u0_u8_u5_U3 (.ZN( u0_u8_u5_n134 ) , .A1( u0_u8_u5_n183 ) , .A2( u0_u8_u5_n190 ) );
  INV_X1 u0_u8_u5_U30 (.A( u0_u8_u5_n123 ) , .ZN( u0_u8_u5_n185 ) );
  INV_X1 u0_u8_u5_U31 (.A( u0_u8_u5_n161 ) , .ZN( u0_u8_u5_n184 ) );
  INV_X1 u0_u8_u5_U32 (.A( u0_u8_u5_n139 ) , .ZN( u0_u8_u5_n189 ) );
  INV_X1 u0_u8_u5_U33 (.A( u0_u8_u5_n157 ) , .ZN( u0_u8_u5_n190 ) );
  INV_X1 u0_u8_u5_U34 (.A( u0_u8_u5_n120 ) , .ZN( u0_u8_u5_n193 ) );
  NAND2_X1 u0_u8_u5_U35 (.ZN( u0_u8_u5_n111 ) , .A1( u0_u8_u5_n140 ) , .A2( u0_u8_u5_n155 ) );
  NOR2_X1 u0_u8_u5_U36 (.ZN( u0_u8_u5_n100 ) , .A1( u0_u8_u5_n170 ) , .A2( u0_u8_u5_n180 ) );
  INV_X1 u0_u8_u5_U37 (.A( u0_u8_u5_n117 ) , .ZN( u0_u8_u5_n196 ) );
  OAI221_X1 u0_u8_u5_U38 (.A( u0_u8_u5_n116 ) , .ZN( u0_u8_u5_n117 ) , .B2( u0_u8_u5_n119 ) , .C1( u0_u8_u5_n153 ) , .C2( u0_u8_u5_n158 ) , .B1( u0_u8_u5_n172 ) );
  AOI222_X1 u0_u8_u5_U39 (.ZN( u0_u8_u5_n116 ) , .B2( u0_u8_u5_n145 ) , .C1( u0_u8_u5_n148 ) , .A2( u0_u8_u5_n174 ) , .C2( u0_u8_u5_n177 ) , .B1( u0_u8_u5_n187 ) , .A1( u0_u8_u5_n193 ) );
  INV_X1 u0_u8_u5_U4 (.A( u0_u8_u5_n138 ) , .ZN( u0_u8_u5_n191 ) );
  INV_X1 u0_u8_u5_U40 (.A( u0_u8_u5_n115 ) , .ZN( u0_u8_u5_n187 ) );
  OAI221_X1 u0_u8_u5_U41 (.A( u0_u8_u5_n101 ) , .ZN( u0_u8_u5_n102 ) , .C2( u0_u8_u5_n115 ) , .C1( u0_u8_u5_n126 ) , .B1( u0_u8_u5_n134 ) , .B2( u0_u8_u5_n160 ) );
  OAI21_X1 u0_u8_u5_U42 (.ZN( u0_u8_u5_n101 ) , .B1( u0_u8_u5_n137 ) , .A( u0_u8_u5_n146 ) , .B2( u0_u8_u5_n147 ) );
  AOI22_X1 u0_u8_u5_U43 (.B2( u0_u8_u5_n131 ) , .A2( u0_u8_u5_n146 ) , .ZN( u0_u8_u5_n169 ) , .B1( u0_u8_u5_n174 ) , .A1( u0_u8_u5_n185 ) );
  NOR2_X1 u0_u8_u5_U44 (.A1( u0_u8_u5_n146 ) , .ZN( u0_u8_u5_n150 ) , .A2( u0_u8_u5_n173 ) );
  AOI21_X1 u0_u8_u5_U45 (.A( u0_u8_u5_n118 ) , .B2( u0_u8_u5_n145 ) , .ZN( u0_u8_u5_n168 ) , .B1( u0_u8_u5_n186 ) );
  INV_X1 u0_u8_u5_U46 (.A( u0_u8_u5_n122 ) , .ZN( u0_u8_u5_n186 ) );
  NOR2_X1 u0_u8_u5_U47 (.A1( u0_u8_u5_n146 ) , .ZN( u0_u8_u5_n152 ) , .A2( u0_u8_u5_n176 ) );
  NOR2_X1 u0_u8_u5_U48 (.A1( u0_u8_u5_n115 ) , .ZN( u0_u8_u5_n118 ) , .A2( u0_u8_u5_n153 ) );
  NOR2_X1 u0_u8_u5_U49 (.A2( u0_u8_u5_n145 ) , .ZN( u0_u8_u5_n156 ) , .A1( u0_u8_u5_n174 ) );
  OAI21_X1 u0_u8_u5_U5 (.B2( u0_u8_u5_n136 ) , .B1( u0_u8_u5_n137 ) , .ZN( u0_u8_u5_n138 ) , .A( u0_u8_u5_n177 ) );
  NOR2_X1 u0_u8_u5_U50 (.ZN( u0_u8_u5_n121 ) , .A2( u0_u8_u5_n145 ) , .A1( u0_u8_u5_n176 ) );
  AOI22_X1 u0_u8_u5_U51 (.ZN( u0_u8_u5_n114 ) , .A2( u0_u8_u5_n137 ) , .A1( u0_u8_u5_n145 ) , .B2( u0_u8_u5_n175 ) , .B1( u0_u8_u5_n193 ) );
  OAI211_X1 u0_u8_u5_U52 (.B( u0_u8_u5_n124 ) , .A( u0_u8_u5_n125 ) , .C2( u0_u8_u5_n126 ) , .C1( u0_u8_u5_n127 ) , .ZN( u0_u8_u5_n128 ) );
  NOR3_X1 u0_u8_u5_U53 (.ZN( u0_u8_u5_n127 ) , .A1( u0_u8_u5_n136 ) , .A3( u0_u8_u5_n148 ) , .A2( u0_u8_u5_n182 ) );
  OAI21_X1 u0_u8_u5_U54 (.ZN( u0_u8_u5_n124 ) , .A( u0_u8_u5_n177 ) , .B2( u0_u8_u5_n183 ) , .B1( u0_u8_u5_n189 ) );
  OAI21_X1 u0_u8_u5_U55 (.ZN( u0_u8_u5_n125 ) , .A( u0_u8_u5_n174 ) , .B2( u0_u8_u5_n185 ) , .B1( u0_u8_u5_n190 ) );
  AOI21_X1 u0_u8_u5_U56 (.A( u0_u8_u5_n153 ) , .B2( u0_u8_u5_n154 ) , .B1( u0_u8_u5_n155 ) , .ZN( u0_u8_u5_n164 ) );
  AOI21_X1 u0_u8_u5_U57 (.ZN( u0_u8_u5_n110 ) , .B1( u0_u8_u5_n122 ) , .B2( u0_u8_u5_n139 ) , .A( u0_u8_u5_n153 ) );
  INV_X1 u0_u8_u5_U58 (.A( u0_u8_u5_n153 ) , .ZN( u0_u8_u5_n176 ) );
  INV_X1 u0_u8_u5_U59 (.A( u0_u8_u5_n126 ) , .ZN( u0_u8_u5_n173 ) );
  AOI222_X1 u0_u8_u5_U6 (.ZN( u0_u8_u5_n113 ) , .A1( u0_u8_u5_n131 ) , .C1( u0_u8_u5_n148 ) , .B2( u0_u8_u5_n174 ) , .C2( u0_u8_u5_n178 ) , .A2( u0_u8_u5_n179 ) , .B1( u0_u8_u5_n99 ) );
  AND2_X1 u0_u8_u5_U60 (.A2( u0_u8_u5_n104 ) , .A1( u0_u8_u5_n107 ) , .ZN( u0_u8_u5_n147 ) );
  AND2_X1 u0_u8_u5_U61 (.A2( u0_u8_u5_n104 ) , .A1( u0_u8_u5_n108 ) , .ZN( u0_u8_u5_n148 ) );
  NAND2_X1 u0_u8_u5_U62 (.A1( u0_u8_u5_n105 ) , .A2( u0_u8_u5_n106 ) , .ZN( u0_u8_u5_n158 ) );
  NAND2_X1 u0_u8_u5_U63 (.A2( u0_u8_u5_n108 ) , .A1( u0_u8_u5_n109 ) , .ZN( u0_u8_u5_n139 ) );
  NAND2_X1 u0_u8_u5_U64 (.A1( u0_u8_u5_n106 ) , .A2( u0_u8_u5_n108 ) , .ZN( u0_u8_u5_n119 ) );
  NAND2_X1 u0_u8_u5_U65 (.A2( u0_u8_u5_n103 ) , .A1( u0_u8_u5_n105 ) , .ZN( u0_u8_u5_n140 ) );
  NAND2_X1 u0_u8_u5_U66 (.A2( u0_u8_u5_n104 ) , .A1( u0_u8_u5_n105 ) , .ZN( u0_u8_u5_n155 ) );
  NAND2_X1 u0_u8_u5_U67 (.A2( u0_u8_u5_n106 ) , .A1( u0_u8_u5_n107 ) , .ZN( u0_u8_u5_n122 ) );
  NAND2_X1 u0_u8_u5_U68 (.A2( u0_u8_u5_n100 ) , .A1( u0_u8_u5_n106 ) , .ZN( u0_u8_u5_n115 ) );
  NAND2_X1 u0_u8_u5_U69 (.A2( u0_u8_u5_n100 ) , .A1( u0_u8_u5_n103 ) , .ZN( u0_u8_u5_n161 ) );
  INV_X1 u0_u8_u5_U7 (.A( u0_u8_u5_n135 ) , .ZN( u0_u8_u5_n178 ) );
  NAND2_X1 u0_u8_u5_U70 (.A1( u0_u8_u5_n105 ) , .A2( u0_u8_u5_n109 ) , .ZN( u0_u8_u5_n154 ) );
  INV_X1 u0_u8_u5_U71 (.A( u0_u8_u5_n146 ) , .ZN( u0_u8_u5_n172 ) );
  NAND2_X1 u0_u8_u5_U72 (.A1( u0_u8_u5_n103 ) , .A2( u0_u8_u5_n108 ) , .ZN( u0_u8_u5_n123 ) );
  NAND2_X1 u0_u8_u5_U73 (.A2( u0_u8_u5_n103 ) , .A1( u0_u8_u5_n107 ) , .ZN( u0_u8_u5_n151 ) );
  NAND2_X1 u0_u8_u5_U74 (.A2( u0_u8_u5_n107 ) , .A1( u0_u8_u5_n109 ) , .ZN( u0_u8_u5_n120 ) );
  NAND2_X1 u0_u8_u5_U75 (.A2( u0_u8_u5_n100 ) , .A1( u0_u8_u5_n109 ) , .ZN( u0_u8_u5_n157 ) );
  AND2_X1 u0_u8_u5_U76 (.A2( u0_u8_u5_n100 ) , .A1( u0_u8_u5_n104 ) , .ZN( u0_u8_u5_n131 ) );
  NOR2_X1 u0_u8_u5_U77 (.A2( u0_u8_X_34 ) , .A1( u0_u8_X_35 ) , .ZN( u0_u8_u5_n145 ) );
  NOR2_X1 u0_u8_u5_U78 (.A2( u0_u8_X_34 ) , .ZN( u0_u8_u5_n146 ) , .A1( u0_u8_u5_n171 ) );
  NOR2_X1 u0_u8_u5_U79 (.A2( u0_u8_X_31 ) , .A1( u0_u8_X_32 ) , .ZN( u0_u8_u5_n103 ) );
  OAI22_X1 u0_u8_u5_U8 (.B2( u0_u8_u5_n149 ) , .B1( u0_u8_u5_n150 ) , .A2( u0_u8_u5_n151 ) , .A1( u0_u8_u5_n152 ) , .ZN( u0_u8_u5_n165 ) );
  NOR2_X1 u0_u8_u5_U80 (.A2( u0_u8_X_36 ) , .ZN( u0_u8_u5_n105 ) , .A1( u0_u8_u5_n180 ) );
  NOR2_X1 u0_u8_u5_U81 (.A2( u0_u8_X_33 ) , .ZN( u0_u8_u5_n108 ) , .A1( u0_u8_u5_n170 ) );
  NOR2_X1 u0_u8_u5_U82 (.A2( u0_u8_X_33 ) , .A1( u0_u8_X_36 ) , .ZN( u0_u8_u5_n107 ) );
  NOR2_X1 u0_u8_u5_U83 (.A2( u0_u8_X_31 ) , .ZN( u0_u8_u5_n104 ) , .A1( u0_u8_u5_n181 ) );
  NAND2_X1 u0_u8_u5_U84 (.A2( u0_u8_X_34 ) , .A1( u0_u8_X_35 ) , .ZN( u0_u8_u5_n153 ) );
  NAND2_X1 u0_u8_u5_U85 (.A1( u0_u8_X_34 ) , .ZN( u0_u8_u5_n126 ) , .A2( u0_u8_u5_n171 ) );
  AND2_X1 u0_u8_u5_U86 (.A1( u0_u8_X_31 ) , .A2( u0_u8_X_32 ) , .ZN( u0_u8_u5_n106 ) );
  AND2_X1 u0_u8_u5_U87 (.A1( u0_u8_X_31 ) , .ZN( u0_u8_u5_n109 ) , .A2( u0_u8_u5_n181 ) );
  INV_X1 u0_u8_u5_U88 (.A( u0_u8_X_33 ) , .ZN( u0_u8_u5_n180 ) );
  INV_X1 u0_u8_u5_U89 (.A( u0_u8_X_35 ) , .ZN( u0_u8_u5_n171 ) );
  NOR3_X1 u0_u8_u5_U9 (.A2( u0_u8_u5_n147 ) , .A1( u0_u8_u5_n148 ) , .ZN( u0_u8_u5_n149 ) , .A3( u0_u8_u5_n194 ) );
  INV_X1 u0_u8_u5_U90 (.A( u0_u8_X_36 ) , .ZN( u0_u8_u5_n170 ) );
  INV_X1 u0_u8_u5_U91 (.A( u0_u8_X_32 ) , .ZN( u0_u8_u5_n181 ) );
  NAND4_X1 u0_u8_u5_U92 (.ZN( u0_out8_29 ) , .A4( u0_u8_u5_n129 ) , .A3( u0_u8_u5_n130 ) , .A2( u0_u8_u5_n168 ) , .A1( u0_u8_u5_n196 ) );
  AOI221_X1 u0_u8_u5_U93 (.A( u0_u8_u5_n128 ) , .ZN( u0_u8_u5_n129 ) , .C2( u0_u8_u5_n132 ) , .B2( u0_u8_u5_n159 ) , .B1( u0_u8_u5_n176 ) , .C1( u0_u8_u5_n184 ) );
  AOI222_X1 u0_u8_u5_U94 (.ZN( u0_u8_u5_n130 ) , .A2( u0_u8_u5_n146 ) , .B1( u0_u8_u5_n147 ) , .C2( u0_u8_u5_n175 ) , .B2( u0_u8_u5_n179 ) , .A1( u0_u8_u5_n188 ) , .C1( u0_u8_u5_n194 ) );
  NAND4_X1 u0_u8_u5_U95 (.ZN( u0_out8_19 ) , .A4( u0_u8_u5_n166 ) , .A3( u0_u8_u5_n167 ) , .A2( u0_u8_u5_n168 ) , .A1( u0_u8_u5_n169 ) );
  AOI22_X1 u0_u8_u5_U96 (.B2( u0_u8_u5_n145 ) , .A2( u0_u8_u5_n146 ) , .ZN( u0_u8_u5_n167 ) , .B1( u0_u8_u5_n182 ) , .A1( u0_u8_u5_n189 ) );
  NOR4_X1 u0_u8_u5_U97 (.A4( u0_u8_u5_n162 ) , .A3( u0_u8_u5_n163 ) , .A2( u0_u8_u5_n164 ) , .A1( u0_u8_u5_n165 ) , .ZN( u0_u8_u5_n166 ) );
  NAND4_X1 u0_u8_u5_U98 (.ZN( u0_out8_11 ) , .A4( u0_u8_u5_n143 ) , .A3( u0_u8_u5_n144 ) , .A2( u0_u8_u5_n169 ) , .A1( u0_u8_u5_n196 ) );
  AOI22_X1 u0_u8_u5_U99 (.A2( u0_u8_u5_n132 ) , .ZN( u0_u8_u5_n144 ) , .B2( u0_u8_u5_n145 ) , .B1( u0_u8_u5_n184 ) , .A1( u0_u8_u5_n194 ) );
  AOI22_X1 u0_u8_u6_U10 (.A2( u0_u8_u6_n151 ) , .B2( u0_u8_u6_n161 ) , .A1( u0_u8_u6_n167 ) , .B1( u0_u8_u6_n170 ) , .ZN( u0_u8_u6_n89 ) );
  AOI21_X1 u0_u8_u6_U11 (.B1( u0_u8_u6_n107 ) , .B2( u0_u8_u6_n132 ) , .A( u0_u8_u6_n158 ) , .ZN( u0_u8_u6_n88 ) );
  AOI21_X1 u0_u8_u6_U12 (.B2( u0_u8_u6_n147 ) , .B1( u0_u8_u6_n148 ) , .ZN( u0_u8_u6_n149 ) , .A( u0_u8_u6_n158 ) );
  AOI21_X1 u0_u8_u6_U13 (.ZN( u0_u8_u6_n106 ) , .A( u0_u8_u6_n142 ) , .B2( u0_u8_u6_n159 ) , .B1( u0_u8_u6_n164 ) );
  INV_X1 u0_u8_u6_U14 (.A( u0_u8_u6_n155 ) , .ZN( u0_u8_u6_n161 ) );
  INV_X1 u0_u8_u6_U15 (.A( u0_u8_u6_n128 ) , .ZN( u0_u8_u6_n164 ) );
  NAND2_X1 u0_u8_u6_U16 (.ZN( u0_u8_u6_n110 ) , .A1( u0_u8_u6_n122 ) , .A2( u0_u8_u6_n129 ) );
  NAND2_X1 u0_u8_u6_U17 (.ZN( u0_u8_u6_n124 ) , .A2( u0_u8_u6_n146 ) , .A1( u0_u8_u6_n148 ) );
  INV_X1 u0_u8_u6_U18 (.A( u0_u8_u6_n132 ) , .ZN( u0_u8_u6_n171 ) );
  AND2_X1 u0_u8_u6_U19 (.A1( u0_u8_u6_n100 ) , .ZN( u0_u8_u6_n130 ) , .A2( u0_u8_u6_n147 ) );
  INV_X1 u0_u8_u6_U20 (.A( u0_u8_u6_n127 ) , .ZN( u0_u8_u6_n173 ) );
  INV_X1 u0_u8_u6_U21 (.A( u0_u8_u6_n121 ) , .ZN( u0_u8_u6_n167 ) );
  INV_X1 u0_u8_u6_U22 (.A( u0_u8_u6_n100 ) , .ZN( u0_u8_u6_n169 ) );
  INV_X1 u0_u8_u6_U23 (.A( u0_u8_u6_n123 ) , .ZN( u0_u8_u6_n170 ) );
  INV_X1 u0_u8_u6_U24 (.A( u0_u8_u6_n113 ) , .ZN( u0_u8_u6_n168 ) );
  AND2_X1 u0_u8_u6_U25 (.A1( u0_u8_u6_n107 ) , .A2( u0_u8_u6_n119 ) , .ZN( u0_u8_u6_n133 ) );
  AND2_X1 u0_u8_u6_U26 (.A2( u0_u8_u6_n121 ) , .A1( u0_u8_u6_n122 ) , .ZN( u0_u8_u6_n131 ) );
  AND3_X1 u0_u8_u6_U27 (.ZN( u0_u8_u6_n120 ) , .A2( u0_u8_u6_n127 ) , .A1( u0_u8_u6_n132 ) , .A3( u0_u8_u6_n145 ) );
  INV_X1 u0_u8_u6_U28 (.A( u0_u8_u6_n146 ) , .ZN( u0_u8_u6_n163 ) );
  AOI222_X1 u0_u8_u6_U29 (.ZN( u0_u8_u6_n114 ) , .A1( u0_u8_u6_n118 ) , .A2( u0_u8_u6_n126 ) , .B2( u0_u8_u6_n151 ) , .C2( u0_u8_u6_n159 ) , .C1( u0_u8_u6_n168 ) , .B1( u0_u8_u6_n169 ) );
  INV_X1 u0_u8_u6_U3 (.A( u0_u8_u6_n110 ) , .ZN( u0_u8_u6_n166 ) );
  NOR2_X1 u0_u8_u6_U30 (.A1( u0_u8_u6_n162 ) , .A2( u0_u8_u6_n165 ) , .ZN( u0_u8_u6_n98 ) );
  AOI211_X1 u0_u8_u6_U31 (.B( u0_u8_u6_n134 ) , .A( u0_u8_u6_n135 ) , .C1( u0_u8_u6_n136 ) , .ZN( u0_u8_u6_n137 ) , .C2( u0_u8_u6_n151 ) );
  AOI21_X1 u0_u8_u6_U32 (.B2( u0_u8_u6_n132 ) , .B1( u0_u8_u6_n133 ) , .ZN( u0_u8_u6_n134 ) , .A( u0_u8_u6_n158 ) );
  NAND4_X1 u0_u8_u6_U33 (.A4( u0_u8_u6_n127 ) , .A3( u0_u8_u6_n128 ) , .A2( u0_u8_u6_n129 ) , .A1( u0_u8_u6_n130 ) , .ZN( u0_u8_u6_n136 ) );
  AOI21_X1 u0_u8_u6_U34 (.B1( u0_u8_u6_n131 ) , .ZN( u0_u8_u6_n135 ) , .A( u0_u8_u6_n144 ) , .B2( u0_u8_u6_n146 ) );
  NAND2_X1 u0_u8_u6_U35 (.A1( u0_u8_u6_n144 ) , .ZN( u0_u8_u6_n151 ) , .A2( u0_u8_u6_n158 ) );
  NAND2_X1 u0_u8_u6_U36 (.ZN( u0_u8_u6_n132 ) , .A1( u0_u8_u6_n91 ) , .A2( u0_u8_u6_n97 ) );
  AOI22_X1 u0_u8_u6_U37 (.B2( u0_u8_u6_n110 ) , .B1( u0_u8_u6_n111 ) , .A1( u0_u8_u6_n112 ) , .ZN( u0_u8_u6_n115 ) , .A2( u0_u8_u6_n161 ) );
  NAND4_X1 u0_u8_u6_U38 (.A3( u0_u8_u6_n109 ) , .ZN( u0_u8_u6_n112 ) , .A4( u0_u8_u6_n132 ) , .A2( u0_u8_u6_n147 ) , .A1( u0_u8_u6_n166 ) );
  NOR2_X1 u0_u8_u6_U39 (.ZN( u0_u8_u6_n109 ) , .A1( u0_u8_u6_n170 ) , .A2( u0_u8_u6_n173 ) );
  INV_X1 u0_u8_u6_U4 (.A( u0_u8_u6_n142 ) , .ZN( u0_u8_u6_n174 ) );
  NOR2_X1 u0_u8_u6_U40 (.A2( u0_u8_u6_n126 ) , .ZN( u0_u8_u6_n155 ) , .A1( u0_u8_u6_n160 ) );
  NAND2_X1 u0_u8_u6_U41 (.ZN( u0_u8_u6_n146 ) , .A2( u0_u8_u6_n94 ) , .A1( u0_u8_u6_n99 ) );
  AOI21_X1 u0_u8_u6_U42 (.A( u0_u8_u6_n144 ) , .B2( u0_u8_u6_n145 ) , .B1( u0_u8_u6_n146 ) , .ZN( u0_u8_u6_n150 ) );
  INV_X1 u0_u8_u6_U43 (.A( u0_u8_u6_n111 ) , .ZN( u0_u8_u6_n158 ) );
  NAND2_X1 u0_u8_u6_U44 (.ZN( u0_u8_u6_n127 ) , .A1( u0_u8_u6_n91 ) , .A2( u0_u8_u6_n92 ) );
  NAND2_X1 u0_u8_u6_U45 (.ZN( u0_u8_u6_n129 ) , .A2( u0_u8_u6_n95 ) , .A1( u0_u8_u6_n96 ) );
  INV_X1 u0_u8_u6_U46 (.A( u0_u8_u6_n144 ) , .ZN( u0_u8_u6_n159 ) );
  NAND2_X1 u0_u8_u6_U47 (.ZN( u0_u8_u6_n145 ) , .A2( u0_u8_u6_n97 ) , .A1( u0_u8_u6_n98 ) );
  NAND2_X1 u0_u8_u6_U48 (.ZN( u0_u8_u6_n148 ) , .A2( u0_u8_u6_n92 ) , .A1( u0_u8_u6_n94 ) );
  NAND2_X1 u0_u8_u6_U49 (.ZN( u0_u8_u6_n108 ) , .A2( u0_u8_u6_n139 ) , .A1( u0_u8_u6_n144 ) );
  NAND2_X1 u0_u8_u6_U5 (.A2( u0_u8_u6_n143 ) , .ZN( u0_u8_u6_n152 ) , .A1( u0_u8_u6_n166 ) );
  NAND2_X1 u0_u8_u6_U50 (.ZN( u0_u8_u6_n121 ) , .A2( u0_u8_u6_n95 ) , .A1( u0_u8_u6_n97 ) );
  NAND2_X1 u0_u8_u6_U51 (.ZN( u0_u8_u6_n107 ) , .A2( u0_u8_u6_n92 ) , .A1( u0_u8_u6_n95 ) );
  AND2_X1 u0_u8_u6_U52 (.ZN( u0_u8_u6_n118 ) , .A2( u0_u8_u6_n91 ) , .A1( u0_u8_u6_n99 ) );
  NAND2_X1 u0_u8_u6_U53 (.ZN( u0_u8_u6_n147 ) , .A2( u0_u8_u6_n98 ) , .A1( u0_u8_u6_n99 ) );
  NAND2_X1 u0_u8_u6_U54 (.ZN( u0_u8_u6_n128 ) , .A1( u0_u8_u6_n94 ) , .A2( u0_u8_u6_n96 ) );
  NAND2_X1 u0_u8_u6_U55 (.ZN( u0_u8_u6_n119 ) , .A2( u0_u8_u6_n95 ) , .A1( u0_u8_u6_n99 ) );
  NAND2_X1 u0_u8_u6_U56 (.ZN( u0_u8_u6_n123 ) , .A2( u0_u8_u6_n91 ) , .A1( u0_u8_u6_n96 ) );
  NAND2_X1 u0_u8_u6_U57 (.ZN( u0_u8_u6_n100 ) , .A2( u0_u8_u6_n92 ) , .A1( u0_u8_u6_n98 ) );
  NAND2_X1 u0_u8_u6_U58 (.ZN( u0_u8_u6_n122 ) , .A1( u0_u8_u6_n94 ) , .A2( u0_u8_u6_n97 ) );
  INV_X1 u0_u8_u6_U59 (.A( u0_u8_u6_n139 ) , .ZN( u0_u8_u6_n160 ) );
  AOI22_X1 u0_u8_u6_U6 (.B2( u0_u8_u6_n101 ) , .A1( u0_u8_u6_n102 ) , .ZN( u0_u8_u6_n103 ) , .B1( u0_u8_u6_n160 ) , .A2( u0_u8_u6_n161 ) );
  NAND2_X1 u0_u8_u6_U60 (.ZN( u0_u8_u6_n113 ) , .A1( u0_u8_u6_n96 ) , .A2( u0_u8_u6_n98 ) );
  NOR2_X1 u0_u8_u6_U61 (.A2( u0_u8_X_40 ) , .A1( u0_u8_X_41 ) , .ZN( u0_u8_u6_n126 ) );
  NOR2_X1 u0_u8_u6_U62 (.A2( u0_u8_X_39 ) , .A1( u0_u8_X_42 ) , .ZN( u0_u8_u6_n92 ) );
  NOR2_X1 u0_u8_u6_U63 (.A2( u0_u8_X_39 ) , .A1( u0_u8_u6_n156 ) , .ZN( u0_u8_u6_n97 ) );
  NOR2_X1 u0_u8_u6_U64 (.A2( u0_u8_X_38 ) , .A1( u0_u8_u6_n165 ) , .ZN( u0_u8_u6_n95 ) );
  NOR2_X1 u0_u8_u6_U65 (.A2( u0_u8_X_41 ) , .ZN( u0_u8_u6_n111 ) , .A1( u0_u8_u6_n157 ) );
  NOR2_X1 u0_u8_u6_U66 (.A2( u0_u8_X_37 ) , .A1( u0_u8_u6_n162 ) , .ZN( u0_u8_u6_n94 ) );
  NOR2_X1 u0_u8_u6_U67 (.A2( u0_u8_X_37 ) , .A1( u0_u8_X_38 ) , .ZN( u0_u8_u6_n91 ) );
  NAND2_X1 u0_u8_u6_U68 (.A1( u0_u8_X_41 ) , .ZN( u0_u8_u6_n144 ) , .A2( u0_u8_u6_n157 ) );
  NAND2_X1 u0_u8_u6_U69 (.A2( u0_u8_X_40 ) , .A1( u0_u8_X_41 ) , .ZN( u0_u8_u6_n139 ) );
  NOR2_X1 u0_u8_u6_U7 (.A1( u0_u8_u6_n118 ) , .ZN( u0_u8_u6_n143 ) , .A2( u0_u8_u6_n168 ) );
  AND2_X1 u0_u8_u6_U70 (.A1( u0_u8_X_39 ) , .A2( u0_u8_u6_n156 ) , .ZN( u0_u8_u6_n96 ) );
  AND2_X1 u0_u8_u6_U71 (.A1( u0_u8_X_39 ) , .A2( u0_u8_X_42 ) , .ZN( u0_u8_u6_n99 ) );
  INV_X1 u0_u8_u6_U72 (.A( u0_u8_X_40 ) , .ZN( u0_u8_u6_n157 ) );
  INV_X1 u0_u8_u6_U73 (.A( u0_u8_X_37 ) , .ZN( u0_u8_u6_n165 ) );
  INV_X1 u0_u8_u6_U74 (.A( u0_u8_X_38 ) , .ZN( u0_u8_u6_n162 ) );
  INV_X1 u0_u8_u6_U75 (.A( u0_u8_X_42 ) , .ZN( u0_u8_u6_n156 ) );
  NAND4_X1 u0_u8_u6_U76 (.ZN( u0_out8_32 ) , .A4( u0_u8_u6_n103 ) , .A3( u0_u8_u6_n104 ) , .A2( u0_u8_u6_n105 ) , .A1( u0_u8_u6_n106 ) );
  AOI22_X1 u0_u8_u6_U77 (.ZN( u0_u8_u6_n105 ) , .A2( u0_u8_u6_n108 ) , .A1( u0_u8_u6_n118 ) , .B2( u0_u8_u6_n126 ) , .B1( u0_u8_u6_n171 ) );
  AOI22_X1 u0_u8_u6_U78 (.ZN( u0_u8_u6_n104 ) , .A1( u0_u8_u6_n111 ) , .B1( u0_u8_u6_n124 ) , .B2( u0_u8_u6_n151 ) , .A2( u0_u8_u6_n93 ) );
  NAND4_X1 u0_u8_u6_U79 (.ZN( u0_out8_12 ) , .A4( u0_u8_u6_n114 ) , .A3( u0_u8_u6_n115 ) , .A2( u0_u8_u6_n116 ) , .A1( u0_u8_u6_n117 ) );
  OAI21_X1 u0_u8_u6_U8 (.A( u0_u8_u6_n159 ) , .B1( u0_u8_u6_n169 ) , .B2( u0_u8_u6_n173 ) , .ZN( u0_u8_u6_n90 ) );
  OAI22_X1 u0_u8_u6_U80 (.B2( u0_u8_u6_n111 ) , .ZN( u0_u8_u6_n116 ) , .B1( u0_u8_u6_n126 ) , .A2( u0_u8_u6_n164 ) , .A1( u0_u8_u6_n167 ) );
  OAI21_X1 u0_u8_u6_U81 (.A( u0_u8_u6_n108 ) , .ZN( u0_u8_u6_n117 ) , .B2( u0_u8_u6_n141 ) , .B1( u0_u8_u6_n163 ) );
  OAI211_X1 u0_u8_u6_U82 (.ZN( u0_out8_7 ) , .B( u0_u8_u6_n153 ) , .C2( u0_u8_u6_n154 ) , .C1( u0_u8_u6_n155 ) , .A( u0_u8_u6_n174 ) );
  NOR3_X1 u0_u8_u6_U83 (.A1( u0_u8_u6_n141 ) , .ZN( u0_u8_u6_n154 ) , .A3( u0_u8_u6_n164 ) , .A2( u0_u8_u6_n171 ) );
  AOI211_X1 u0_u8_u6_U84 (.B( u0_u8_u6_n149 ) , .A( u0_u8_u6_n150 ) , .C2( u0_u8_u6_n151 ) , .C1( u0_u8_u6_n152 ) , .ZN( u0_u8_u6_n153 ) );
  OAI211_X1 u0_u8_u6_U85 (.ZN( u0_out8_22 ) , .B( u0_u8_u6_n137 ) , .A( u0_u8_u6_n138 ) , .C2( u0_u8_u6_n139 ) , .C1( u0_u8_u6_n140 ) );
  AOI22_X1 u0_u8_u6_U86 (.B1( u0_u8_u6_n124 ) , .A2( u0_u8_u6_n125 ) , .A1( u0_u8_u6_n126 ) , .ZN( u0_u8_u6_n138 ) , .B2( u0_u8_u6_n161 ) );
  AND4_X1 u0_u8_u6_U87 (.A3( u0_u8_u6_n119 ) , .A1( u0_u8_u6_n120 ) , .A4( u0_u8_u6_n129 ) , .ZN( u0_u8_u6_n140 ) , .A2( u0_u8_u6_n143 ) );
  NAND3_X1 u0_u8_u6_U88 (.A2( u0_u8_u6_n123 ) , .ZN( u0_u8_u6_n125 ) , .A1( u0_u8_u6_n130 ) , .A3( u0_u8_u6_n131 ) );
  NAND3_X1 u0_u8_u6_U89 (.A3( u0_u8_u6_n133 ) , .ZN( u0_u8_u6_n141 ) , .A1( u0_u8_u6_n145 ) , .A2( u0_u8_u6_n148 ) );
  INV_X1 u0_u8_u6_U9 (.ZN( u0_u8_u6_n172 ) , .A( u0_u8_u6_n88 ) );
  NAND3_X1 u0_u8_u6_U90 (.ZN( u0_u8_u6_n101 ) , .A3( u0_u8_u6_n107 ) , .A2( u0_u8_u6_n121 ) , .A1( u0_u8_u6_n127 ) );
  NAND3_X1 u0_u8_u6_U91 (.ZN( u0_u8_u6_n102 ) , .A3( u0_u8_u6_n130 ) , .A2( u0_u8_u6_n145 ) , .A1( u0_u8_u6_n166 ) );
  NAND3_X1 u0_u8_u6_U92 (.A3( u0_u8_u6_n113 ) , .A1( u0_u8_u6_n119 ) , .A2( u0_u8_u6_n123 ) , .ZN( u0_u8_u6_n93 ) );
  NAND3_X1 u0_u8_u6_U93 (.ZN( u0_u8_u6_n142 ) , .A2( u0_u8_u6_n172 ) , .A3( u0_u8_u6_n89 ) , .A1( u0_u8_u6_n90 ) );
  OAI22_X1 u0_uk_U101 (.ZN( u0_K9_5 ) , .A1( u0_uk_n142 ) , .B1( u0_uk_n155 ) , .A2( u0_uk_n272 ) , .B2( u0_uk_n278 ) );
  NAND2_X1 u0_uk_U1011 (.A1( u0_key_r_10 ) , .A2( u0_uk_n27 ) , .ZN( u0_uk_n888 ) );
  OAI22_X1 u0_uk_U103 (.ZN( u0_K5_5 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n182 ) , .B2( u0_uk_n466 ) , .A2( u0_uk_n490 ) );
  OAI21_X1 u0_uk_U1032 (.ZN( u0_K8_41 ) , .B2( u0_uk_n341 ) , .B1( u0_uk_n63 ) , .A( u0_uk_n748 ) );
  NAND2_X1 u0_uk_U1039 (.A1( u0_uk_K_r6_51 ) , .A2( u0_uk_n10 ) , .ZN( u0_uk_n756 ) );
  OAI21_X1 u0_uk_U1054 (.ZN( u0_K8_42 ) , .B1( u0_uk_n31 ) , .B2( u0_uk_n348 ) , .A( u0_uk_n747 ) );
  NAND2_X1 u0_uk_U1055 (.A1( u0_uk_K_r6_22 ) , .A2( u0_uk_n10 ) , .ZN( u0_uk_n747 ) );
  OAI21_X1 u0_uk_U1095 (.ZN( u0_K8_39 ) , .B1( u0_uk_n191 ) , .B2( u0_uk_n332 ) , .A( u0_uk_n750 ) );
  NAND2_X1 u0_uk_U1096 (.A1( u0_uk_K_r6_31 ) , .A2( u0_uk_n208 ) , .ZN( u0_uk_n750 ) );
  INV_X1 u0_uk_U1105 (.ZN( u0_K1_18 ) , .A( u0_uk_n887 ) );
  AOI22_X1 u0_uk_U1106 (.A2( u0_key_r_5 ) , .B2( u0_key_r_55 ) , .B1( u0_uk_n145 ) , .A1( u0_uk_n240 ) , .ZN( u0_uk_n887 ) );
  INV_X1 u0_uk_U1129 (.ZN( u0_K9_41 ) , .A( u0_uk_n723 ) );
  AOI22_X1 u0_uk_U1130 (.B2( u0_uk_K_r7_23 ) , .A2( u0_uk_K_r7_30 ) , .B1( u0_uk_n129 ) , .A1( u0_uk_n148 ) , .ZN( u0_uk_n723 ) );
  INV_X1 u0_uk_U1133 (.ZN( u0_K9_42 ) , .A( u0_uk_n722 ) );
  AOI22_X1 u0_uk_U1134 (.B2( u0_uk_K_r7_15 ) , .A2( u0_uk_K_r7_22 ) , .B1( u0_uk_n129 ) , .A1( u0_uk_n220 ) , .ZN( u0_uk_n722 ) );
  AOI22_X1 u0_uk_U1149 (.B2( u0_uk_K_r3_15 ) , .A2( u0_uk_K_r3_38 ) , .B1( u0_uk_n141 ) , .A1( u0_uk_n230 ) , .ZN( u0_uk_n806 ) );
  INV_X1 u0_uk_U1150 (.ZN( u0_K5_43 ) , .A( u0_uk_n806 ) );
  OAI21_X1 u0_uk_U1151 (.ZN( u0_K5_6 ) , .B1( u0_uk_n109 ) , .B2( u0_uk_n471 ) , .A( u0_uk_n803 ) );
  NAND2_X1 u0_uk_U1152 (.A1( u0_uk_K_r3_10 ) , .ZN( u0_uk_n803 ) , .A2( u0_uk_n93 ) );
  AOI22_X1 u0_uk_U1153 (.B2( u0_uk_K_r7_24 ) , .A2( u0_uk_K_r7_6 ) , .B1( u0_uk_n10 ) , .A1( u0_uk_n242 ) , .ZN( u0_uk_n734 ) );
  INV_X1 u0_uk_U1154 (.ZN( u0_K9_1 ) , .A( u0_uk_n734 ) );
  AOI22_X1 u0_uk_U1162 (.B2( u0_uk_K_r7_20 ) , .A2( u0_uk_K_r7_27 ) , .B1( u0_uk_n129 ) , .A1( u0_uk_n238 ) , .ZN( u0_uk_n729 ) );
  INV_X1 u0_uk_U1163 (.ZN( u0_K9_2 ) , .A( u0_uk_n729 ) );
  OAI21_X1 u0_uk_U173 (.ZN( u0_K8_30 ) , .B1( u0_uk_n250 ) , .B2( u0_uk_n333 ) , .A( u0_uk_n753 ) );
  NAND2_X1 u0_uk_U174 (.A1( u0_uk_K_r6_29 ) , .A2( u0_uk_n207 ) , .ZN( u0_uk_n753 ) );
  NAND2_X1 u0_uk_U202 (.A1( u0_key_r_45 ) , .A2( u0_uk_n27 ) , .ZN( u0_uk_n880 ) );
  OAI22_X1 u0_uk_U215 (.ZN( u0_K8_31 ) , .A1( u0_uk_n102 ) , .B1( u0_uk_n223 ) , .A2( u0_uk_n321 ) , .B2( u0_uk_n359 ) );
  INV_X1 u0_uk_U23 (.ZN( u0_uk_n10 ) , .A( u0_uk_n148 ) );
  OAI22_X1 u0_uk_U235 (.ZN( u0_K9_31 ) , .A1( u0_uk_n257 ) , .B1( u0_uk_n27 ) , .A2( u0_uk_n275 ) , .B2( u0_uk_n316 ) );
  OAI22_X1 u0_uk_U318 (.ZN( u0_K8_26 ) , .A1( u0_uk_n102 ) , .B1( u0_uk_n222 ) , .B2( u0_uk_n348 ) , .A2( u0_uk_n355 ) );
  OAI22_X1 u0_uk_U325 (.ZN( u0_K5_46 ) , .A1( u0_uk_n100 ) , .B1( u0_uk_n214 ) , .A2( u0_uk_n457 ) , .B2( u0_uk_n494 ) );
  NAND2_X1 u0_uk_U336 (.A1( u0_uk_K_r14_3 ) , .A2( u0_uk_n10 ) , .ZN( u0_uk_n894 ) );
  OAI22_X1 u0_uk_U363 (.ZN( u0_K8_40 ) , .A1( u0_uk_n162 ) , .B1( u0_uk_n27 ) , .A2( u0_uk_n327 ) , .B2( u0_uk_n333 ) );
  OAI22_X1 u0_uk_U395 (.ZN( u0_K9_16 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n231 ) , .A2( u0_uk_n303 ) , .B2( u0_uk_n310 ) );
  NAND2_X1 u0_uk_U405 (.A1( u0_uk_K_r12_18 ) , .A2( u0_uk_n10 ) , .ZN( u0_uk_n926 ) );
  INV_X1 u0_uk_U414 (.ZN( u0_K8_37 ) , .A( u0_uk_n751 ) );
  AOI22_X1 u0_uk_U415 (.B2( u0_uk_K_r6_14 ) , .A2( u0_uk_K_r6_7 ) , .B1( u0_uk_n141 ) , .A1( u0_uk_n240 ) , .ZN( u0_uk_n751 ) );
  INV_X1 u0_uk_U418 (.ZN( u0_K9_9 ) , .A( u0_uk_n718 ) );
  AOI22_X1 u0_uk_U419 (.B2( u0_uk_K_r7_13 ) , .A1( u0_uk_K_r7_6 ) , .A2( u0_uk_n128 ) , .B1( u0_uk_n207 ) , .ZN( u0_uk_n718 ) );
  INV_X1 u0_uk_U437 (.ZN( u0_K9_33 ) , .A( u0_uk_n727 ) );
  AOI22_X1 u0_uk_U438 (.B2( u0_uk_K_r7_1 ) , .A2( u0_uk_K_r7_8 ) , .B1( u0_uk_n129 ) , .A1( u0_uk_n238 ) , .ZN( u0_uk_n727 ) );
  OAI21_X1 u0_uk_U459 (.ZN( u0_K9_37 ) , .B1( u0_uk_n17 ) , .B2( u0_uk_n307 ) , .A( u0_uk_n725 ) );
  OAI21_X1 u0_uk_U497 (.ZN( u0_K9_12 ) , .B1( u0_uk_n17 ) , .B2( u0_uk_n315 ) , .A( u0_uk_n740 ) );
  INV_X1 u0_uk_U5 (.ZN( u0_uk_n141 ) , .A( u0_uk_n191 ) );
  OAI21_X1 u0_uk_U504 (.ZN( u0_K9_17 ) , .B2( u0_uk_n290 ) , .A( u0_uk_n737 ) , .B1( u0_uk_n99 ) );
  NAND2_X1 u0_uk_U505 (.A1( u0_uk_K_r7_26 ) , .A2( u0_uk_n10 ) , .ZN( u0_uk_n737 ) );
  INV_X1 u0_uk_U506 (.ZN( u0_K8_29 ) , .A( u0_uk_n755 ) );
  OAI22_X1 u0_uk_U530 (.ZN( u0_K5_2 ) , .A1( u0_uk_n109 ) , .B1( u0_uk_n222 ) , .B2( u0_uk_n486 ) , .A2( u0_uk_n491 ) );
  OAI22_X1 u0_uk_U536 (.ZN( u0_K9_36 ) , .A1( u0_uk_n142 ) , .B1( u0_uk_n161 ) , .A2( u0_uk_n283 ) , .B2( u0_uk_n289 ) );
  OAI22_X1 u0_uk_U557 (.ZN( u0_K9_38 ) , .A1( u0_uk_n145 ) , .B1( u0_uk_n155 ) , .A2( u0_uk_n276 ) , .B2( u0_uk_n283 ) );
  INV_X1 u0_uk_U579 (.ZN( u0_K9_10 ) , .A( u0_uk_n742 ) );
  AOI22_X1 u0_uk_U580 (.B2( u0_uk_K_r7_25 ) , .A2( u0_uk_K_r7_32 ) , .B1( u0_uk_n128 ) , .A1( u0_uk_n242 ) , .ZN( u0_uk_n742 ) );
  OAI22_X1 u0_uk_U605 (.ZN( u0_K8_35 ) , .A1( u0_uk_n242 ) , .B1( u0_uk_n31 ) , .A2( u0_uk_n341 ) , .B2( u0_uk_n347 ) );
  INV_X1 u0_uk_U616 (.ZN( u0_K9_35 ) , .A( u0_uk_n726 ) );
  INV_X1 u0_uk_U62 (.ZN( u0_K8_34 ) , .A( u0_uk_n752 ) );
  AOI22_X1 u0_uk_U63 (.B2( u0_uk_K_r6_14 ) , .A2( u0_uk_K_r6_21 ) , .A1( u0_uk_n141 ) , .B1( u0_uk_n202 ) , .ZN( u0_uk_n752 ) );
  NAND2_X1 u0_uk_U632 (.A1( u0_uk_K_r6_55 ) , .A2( u0_uk_n10 ) , .ZN( u0_uk_n762 ) );
  INV_X1 u0_uk_U637 (.ZN( u0_K9_11 ) , .A( u0_uk_n741 ) );
  AOI22_X1 u0_uk_U638 (.B2( u0_uk_K_r7_48 ) , .A2( u0_uk_K_r7_55 ) , .A1( u0_uk_n251 ) , .ZN( u0_uk_n741 ) , .B1( u0_uk_n99 ) );
  OAI21_X1 u0_uk_U673 (.ZN( u0_K5_45 ) , .B1( u0_uk_n10 ) , .B2( u0_uk_n488 ) , .A( u0_uk_n805 ) );
  NAND2_X1 u0_uk_U681 (.A1( u0_uk_K_r10_19 ) , .A2( u0_uk_n27 ) , .ZN( u0_uk_n961 ) );
  INV_X1 u0_uk_U7 (.A( u0_uk_n147 ) , .ZN( u0_uk_n27 ) );
  OAI22_X1 u0_uk_U701 (.ZN( u0_K8_25 ) , .A1( u0_uk_n161 ) , .A2( u0_uk_n320 ) , .B2( u0_uk_n325 ) , .B1( u0_uk_n60 ) );
  OAI22_X1 u0_uk_U718 (.ZN( u0_K8_32 ) , .A1( u0_uk_n213 ) , .B1( u0_uk_n27 ) , .A2( u0_uk_n325 ) , .B2( u0_uk_n332 ) );
  OAI22_X1 u0_uk_U749 (.ZN( u0_K8_27 ) , .B1( u0_uk_n128 ) , .A1( u0_uk_n257 ) , .A2( u0_uk_n354 ) , .B2( u0_uk_n359 ) );
  OAI21_X1 u0_uk_U757 (.ZN( u0_K9_13 ) , .B2( u0_uk_n309 ) , .B1( u0_uk_n63 ) , .A( u0_uk_n739 ) );
  NAND2_X1 u0_uk_U816 (.A1( u0_uk_K_r14_5 ) , .A2( u0_uk_n10 ) , .ZN( u0_uk_n906 ) );
  INV_X1 u0_uk_U825 (.ZN( u0_K9_18 ) , .A( u0_uk_n736 ) );
  OAI22_X1 u0_uk_U895 (.ZN( u0_K9_3 ) , .A1( u0_uk_n161 ) , .B1( u0_uk_n27 ) , .B2( u0_uk_n311 ) , .A2( u0_uk_n315 ) );
  OAI22_X1 u0_uk_U896 (.ZN( u0_K9_7 ) , .A1( u0_uk_n257 ) , .B1( u0_uk_n27 ) , .B2( u0_uk_n310 ) , .A2( u0_uk_n314 ) );
  OAI22_X1 u0_uk_U921 (.ZN( u0_K8_38 ) , .A1( u0_uk_n223 ) , .B1( u0_uk_n27 ) , .A2( u0_uk_n322 ) , .B2( u0_uk_n328 ) );
  OAI22_X1 u0_uk_U937 (.ZN( u0_K9_8 ) , .A1( u0_uk_n100 ) , .B1( u0_uk_n147 ) , .A2( u0_uk_n278 ) , .B2( u0_uk_n285 ) );
  OAI22_X1 u0_uk_U950 (.ZN( u0_K9_34 ) , .A1( u0_uk_n11 ) , .B1( u0_uk_n161 ) , .A2( u0_uk_n300 ) , .B2( u0_uk_n307 ) );
  XOR2_X1 u2_U101 (.B( u2_L12_26 ) , .Z( u2_N441 ) , .A( u2_out13_26 ) );
  XOR2_X1 u2_U108 (.B( u2_L12_20 ) , .Z( u2_N435 ) , .A( u2_out13_20 ) );
  XOR2_X1 u2_U119 (.B( u2_L12_10 ) , .Z( u2_N425 ) , .A( u2_out13_10 ) );
  XOR2_X1 u2_U129 (.B( u2_L12_1 ) , .Z( u2_N416 ) , .A( u2_out13_1 ) );
  XOR2_X1 u2_U238 (.B( u2_L8_31 ) , .Z( u2_N318 ) , .A( u2_out9_31 ) );
  XOR2_X1 u2_U242 (.B( u2_L8_27 ) , .Z( u2_N314 ) , .A( u2_out9_27 ) );
  XOR2_X1 u2_U244 (.B( u2_L8_25 ) , .Z( u2_N312 ) , .A( u2_out9_25 ) );
  XOR2_X1 u2_U246 (.B( u2_L8_23 ) , .Z( u2_N310 ) , .A( u2_out9_23 ) );
  XOR2_X1 u2_U249 (.B( u2_L8_21 ) , .Z( u2_N308 ) , .A( u2_out9_21 ) );
  XOR2_X1 u2_U253 (.B( u2_L8_17 ) , .Z( u2_N304 ) , .A( u2_out9_17 ) );
  XOR2_X1 u2_U255 (.B( u2_L8_15 ) , .Z( u2_N302 ) , .A( u2_out9_15 ) );
  XOR2_X1 u2_U256 (.B( u2_L8_14 ) , .Z( u2_N301 ) , .A( u2_out9_14 ) );
  XOR2_X1 u2_U263 (.B( u2_L8_9 ) , .Z( u2_N296 ) , .A( u2_out9_9 ) );
  XOR2_X1 u2_U264 (.B( u2_L8_8 ) , .Z( u2_N295 ) , .A( u2_out9_8 ) );
  XOR2_X1 u2_U267 (.B( u2_L8_5 ) , .Z( u2_N292 ) , .A( u2_out9_5 ) );
  XOR2_X1 u2_U269 (.B( u2_L8_3 ) , .Z( u2_N290 ) , .A( u2_out9_3 ) );
  XOR2_X1 u2_U420 (.B( u2_L3_27 ) , .Z( u2_N154 ) , .A( u2_out4_27 ) );
  XOR2_X1 u2_U427 (.B( u2_L3_21 ) , .Z( u2_N148 ) , .A( u2_out4_21 ) );
  XOR2_X1 u2_U433 (.B( u2_L3_15 ) , .Z( u2_N142 ) , .A( u2_out4_15 ) );
  XOR2_X1 u2_U444 (.B( u2_L3_5 ) , .Z( u2_N132 ) , .A( u2_out4_5 ) );
  XOR2_X1 u2_u13_U33 (.B( u2_K14_24 ) , .A( u2_R12_17 ) , .Z( u2_u13_X_24 ) );
  XOR2_X1 u2_u13_U34 (.B( u2_K14_23 ) , .A( u2_R12_16 ) , .Z( u2_u13_X_23 ) );
  XOR2_X1 u2_u13_U35 (.B( u2_K14_22 ) , .A( u2_R12_15 ) , .Z( u2_u13_X_22 ) );
  XOR2_X1 u2_u13_U36 (.B( u2_K14_21 ) , .A( u2_R12_14 ) , .Z( u2_u13_X_21 ) );
  XOR2_X1 u2_u13_U37 (.B( u2_K14_20 ) , .A( u2_R12_13 ) , .Z( u2_u13_X_20 ) );
  XOR2_X1 u2_u13_U39 (.B( u2_K14_19 ) , .A( u2_R12_12 ) , .Z( u2_u13_X_19 ) );
  OAI22_X1 u2_u13_u3_U10 (.B1( u2_u13_u3_n113 ) , .A2( u2_u13_u3_n135 ) , .A1( u2_u13_u3_n150 ) , .B2( u2_u13_u3_n164 ) , .ZN( u2_u13_u3_n98 ) );
  OAI211_X1 u2_u13_u3_U11 (.B( u2_u13_u3_n106 ) , .ZN( u2_u13_u3_n119 ) , .C2( u2_u13_u3_n128 ) , .C1( u2_u13_u3_n167 ) , .A( u2_u13_u3_n181 ) );
  AOI221_X1 u2_u13_u3_U12 (.C1( u2_u13_u3_n105 ) , .ZN( u2_u13_u3_n106 ) , .A( u2_u13_u3_n131 ) , .B2( u2_u13_u3_n132 ) , .C2( u2_u13_u3_n133 ) , .B1( u2_u13_u3_n169 ) );
  INV_X1 u2_u13_u3_U13 (.ZN( u2_u13_u3_n181 ) , .A( u2_u13_u3_n98 ) );
  NAND2_X1 u2_u13_u3_U14 (.ZN( u2_u13_u3_n105 ) , .A2( u2_u13_u3_n130 ) , .A1( u2_u13_u3_n155 ) );
  AOI22_X1 u2_u13_u3_U15 (.B1( u2_u13_u3_n115 ) , .A2( u2_u13_u3_n116 ) , .ZN( u2_u13_u3_n123 ) , .B2( u2_u13_u3_n133 ) , .A1( u2_u13_u3_n169 ) );
  NAND2_X1 u2_u13_u3_U16 (.ZN( u2_u13_u3_n116 ) , .A2( u2_u13_u3_n151 ) , .A1( u2_u13_u3_n182 ) );
  NOR2_X1 u2_u13_u3_U17 (.ZN( u2_u13_u3_n126 ) , .A2( u2_u13_u3_n150 ) , .A1( u2_u13_u3_n164 ) );
  AOI21_X1 u2_u13_u3_U18 (.ZN( u2_u13_u3_n112 ) , .B2( u2_u13_u3_n146 ) , .B1( u2_u13_u3_n155 ) , .A( u2_u13_u3_n167 ) );
  NAND2_X1 u2_u13_u3_U19 (.A1( u2_u13_u3_n135 ) , .ZN( u2_u13_u3_n142 ) , .A2( u2_u13_u3_n164 ) );
  NAND2_X1 u2_u13_u3_U20 (.ZN( u2_u13_u3_n132 ) , .A2( u2_u13_u3_n152 ) , .A1( u2_u13_u3_n156 ) );
  AND2_X1 u2_u13_u3_U21 (.A2( u2_u13_u3_n113 ) , .A1( u2_u13_u3_n114 ) , .ZN( u2_u13_u3_n151 ) );
  INV_X1 u2_u13_u3_U22 (.A( u2_u13_u3_n133 ) , .ZN( u2_u13_u3_n165 ) );
  INV_X1 u2_u13_u3_U23 (.A( u2_u13_u3_n135 ) , .ZN( u2_u13_u3_n170 ) );
  NAND2_X1 u2_u13_u3_U24 (.A1( u2_u13_u3_n107 ) , .A2( u2_u13_u3_n108 ) , .ZN( u2_u13_u3_n140 ) );
  NAND2_X1 u2_u13_u3_U25 (.ZN( u2_u13_u3_n117 ) , .A1( u2_u13_u3_n124 ) , .A2( u2_u13_u3_n148 ) );
  NAND2_X1 u2_u13_u3_U26 (.ZN( u2_u13_u3_n143 ) , .A1( u2_u13_u3_n165 ) , .A2( u2_u13_u3_n167 ) );
  INV_X1 u2_u13_u3_U27 (.A( u2_u13_u3_n130 ) , .ZN( u2_u13_u3_n177 ) );
  INV_X1 u2_u13_u3_U28 (.A( u2_u13_u3_n128 ) , .ZN( u2_u13_u3_n176 ) );
  INV_X1 u2_u13_u3_U29 (.A( u2_u13_u3_n155 ) , .ZN( u2_u13_u3_n174 ) );
  INV_X1 u2_u13_u3_U3 (.A( u2_u13_u3_n129 ) , .ZN( u2_u13_u3_n183 ) );
  INV_X1 u2_u13_u3_U30 (.A( u2_u13_u3_n139 ) , .ZN( u2_u13_u3_n185 ) );
  NOR2_X1 u2_u13_u3_U31 (.ZN( u2_u13_u3_n135 ) , .A2( u2_u13_u3_n141 ) , .A1( u2_u13_u3_n169 ) );
  OAI222_X1 u2_u13_u3_U32 (.C2( u2_u13_u3_n107 ) , .A2( u2_u13_u3_n108 ) , .B1( u2_u13_u3_n135 ) , .ZN( u2_u13_u3_n138 ) , .B2( u2_u13_u3_n146 ) , .C1( u2_u13_u3_n154 ) , .A1( u2_u13_u3_n164 ) );
  NOR4_X1 u2_u13_u3_U33 (.A4( u2_u13_u3_n157 ) , .A3( u2_u13_u3_n158 ) , .A2( u2_u13_u3_n159 ) , .A1( u2_u13_u3_n160 ) , .ZN( u2_u13_u3_n161 ) );
  AOI21_X1 u2_u13_u3_U34 (.B2( u2_u13_u3_n152 ) , .B1( u2_u13_u3_n153 ) , .ZN( u2_u13_u3_n158 ) , .A( u2_u13_u3_n164 ) );
  AOI21_X1 u2_u13_u3_U35 (.A( u2_u13_u3_n154 ) , .B2( u2_u13_u3_n155 ) , .B1( u2_u13_u3_n156 ) , .ZN( u2_u13_u3_n157 ) );
  AOI21_X1 u2_u13_u3_U36 (.A( u2_u13_u3_n149 ) , .B2( u2_u13_u3_n150 ) , .B1( u2_u13_u3_n151 ) , .ZN( u2_u13_u3_n159 ) );
  AOI211_X1 u2_u13_u3_U37 (.ZN( u2_u13_u3_n109 ) , .A( u2_u13_u3_n119 ) , .C2( u2_u13_u3_n129 ) , .B( u2_u13_u3_n138 ) , .C1( u2_u13_u3_n141 ) );
  AOI211_X1 u2_u13_u3_U38 (.B( u2_u13_u3_n119 ) , .A( u2_u13_u3_n120 ) , .C2( u2_u13_u3_n121 ) , .ZN( u2_u13_u3_n122 ) , .C1( u2_u13_u3_n179 ) );
  INV_X1 u2_u13_u3_U39 (.A( u2_u13_u3_n156 ) , .ZN( u2_u13_u3_n179 ) );
  INV_X1 u2_u13_u3_U4 (.A( u2_u13_u3_n140 ) , .ZN( u2_u13_u3_n182 ) );
  OAI22_X1 u2_u13_u3_U40 (.B1( u2_u13_u3_n118 ) , .ZN( u2_u13_u3_n120 ) , .A1( u2_u13_u3_n135 ) , .B2( u2_u13_u3_n154 ) , .A2( u2_u13_u3_n178 ) );
  AND3_X1 u2_u13_u3_U41 (.ZN( u2_u13_u3_n118 ) , .A2( u2_u13_u3_n124 ) , .A1( u2_u13_u3_n144 ) , .A3( u2_u13_u3_n152 ) );
  INV_X1 u2_u13_u3_U42 (.A( u2_u13_u3_n121 ) , .ZN( u2_u13_u3_n164 ) );
  NAND2_X1 u2_u13_u3_U43 (.ZN( u2_u13_u3_n133 ) , .A1( u2_u13_u3_n154 ) , .A2( u2_u13_u3_n164 ) );
  OAI211_X1 u2_u13_u3_U44 (.B( u2_u13_u3_n127 ) , .ZN( u2_u13_u3_n139 ) , .C1( u2_u13_u3_n150 ) , .C2( u2_u13_u3_n154 ) , .A( u2_u13_u3_n184 ) );
  INV_X1 u2_u13_u3_U45 (.A( u2_u13_u3_n125 ) , .ZN( u2_u13_u3_n184 ) );
  AOI221_X1 u2_u13_u3_U46 (.A( u2_u13_u3_n126 ) , .ZN( u2_u13_u3_n127 ) , .C2( u2_u13_u3_n132 ) , .C1( u2_u13_u3_n169 ) , .B2( u2_u13_u3_n170 ) , .B1( u2_u13_u3_n174 ) );
  OAI22_X1 u2_u13_u3_U47 (.A1( u2_u13_u3_n124 ) , .ZN( u2_u13_u3_n125 ) , .B2( u2_u13_u3_n145 ) , .A2( u2_u13_u3_n165 ) , .B1( u2_u13_u3_n167 ) );
  NOR2_X1 u2_u13_u3_U48 (.A1( u2_u13_u3_n113 ) , .ZN( u2_u13_u3_n131 ) , .A2( u2_u13_u3_n154 ) );
  NAND2_X1 u2_u13_u3_U49 (.A1( u2_u13_u3_n103 ) , .ZN( u2_u13_u3_n150 ) , .A2( u2_u13_u3_n99 ) );
  INV_X1 u2_u13_u3_U5 (.A( u2_u13_u3_n117 ) , .ZN( u2_u13_u3_n178 ) );
  NAND2_X1 u2_u13_u3_U50 (.A2( u2_u13_u3_n102 ) , .ZN( u2_u13_u3_n155 ) , .A1( u2_u13_u3_n97 ) );
  INV_X1 u2_u13_u3_U51 (.A( u2_u13_u3_n141 ) , .ZN( u2_u13_u3_n167 ) );
  AOI21_X1 u2_u13_u3_U52 (.B2( u2_u13_u3_n114 ) , .B1( u2_u13_u3_n146 ) , .A( u2_u13_u3_n154 ) , .ZN( u2_u13_u3_n94 ) );
  AOI21_X1 u2_u13_u3_U53 (.ZN( u2_u13_u3_n110 ) , .B2( u2_u13_u3_n142 ) , .B1( u2_u13_u3_n186 ) , .A( u2_u13_u3_n95 ) );
  INV_X1 u2_u13_u3_U54 (.A( u2_u13_u3_n145 ) , .ZN( u2_u13_u3_n186 ) );
  AOI21_X1 u2_u13_u3_U55 (.B1( u2_u13_u3_n124 ) , .A( u2_u13_u3_n149 ) , .B2( u2_u13_u3_n155 ) , .ZN( u2_u13_u3_n95 ) );
  INV_X1 u2_u13_u3_U56 (.A( u2_u13_u3_n149 ) , .ZN( u2_u13_u3_n169 ) );
  NAND2_X1 u2_u13_u3_U57 (.ZN( u2_u13_u3_n124 ) , .A1( u2_u13_u3_n96 ) , .A2( u2_u13_u3_n97 ) );
  NAND2_X1 u2_u13_u3_U58 (.A2( u2_u13_u3_n100 ) , .ZN( u2_u13_u3_n146 ) , .A1( u2_u13_u3_n96 ) );
  NAND2_X1 u2_u13_u3_U59 (.A1( u2_u13_u3_n101 ) , .ZN( u2_u13_u3_n145 ) , .A2( u2_u13_u3_n99 ) );
  AOI221_X1 u2_u13_u3_U6 (.A( u2_u13_u3_n131 ) , .C2( u2_u13_u3_n132 ) , .C1( u2_u13_u3_n133 ) , .ZN( u2_u13_u3_n134 ) , .B1( u2_u13_u3_n143 ) , .B2( u2_u13_u3_n177 ) );
  NAND2_X1 u2_u13_u3_U60 (.A1( u2_u13_u3_n100 ) , .ZN( u2_u13_u3_n156 ) , .A2( u2_u13_u3_n99 ) );
  NAND2_X1 u2_u13_u3_U61 (.A2( u2_u13_u3_n101 ) , .A1( u2_u13_u3_n104 ) , .ZN( u2_u13_u3_n148 ) );
  NAND2_X1 u2_u13_u3_U62 (.A1( u2_u13_u3_n100 ) , .A2( u2_u13_u3_n102 ) , .ZN( u2_u13_u3_n128 ) );
  NAND2_X1 u2_u13_u3_U63 (.A2( u2_u13_u3_n101 ) , .A1( u2_u13_u3_n102 ) , .ZN( u2_u13_u3_n152 ) );
  NAND2_X1 u2_u13_u3_U64 (.A2( u2_u13_u3_n101 ) , .ZN( u2_u13_u3_n114 ) , .A1( u2_u13_u3_n96 ) );
  NAND2_X1 u2_u13_u3_U65 (.ZN( u2_u13_u3_n107 ) , .A1( u2_u13_u3_n97 ) , .A2( u2_u13_u3_n99 ) );
  NAND2_X1 u2_u13_u3_U66 (.A2( u2_u13_u3_n100 ) , .A1( u2_u13_u3_n104 ) , .ZN( u2_u13_u3_n113 ) );
  NAND2_X1 u2_u13_u3_U67 (.A1( u2_u13_u3_n104 ) , .ZN( u2_u13_u3_n153 ) , .A2( u2_u13_u3_n97 ) );
  NAND2_X1 u2_u13_u3_U68 (.A2( u2_u13_u3_n103 ) , .A1( u2_u13_u3_n104 ) , .ZN( u2_u13_u3_n130 ) );
  NAND2_X1 u2_u13_u3_U69 (.A2( u2_u13_u3_n103 ) , .ZN( u2_u13_u3_n144 ) , .A1( u2_u13_u3_n96 ) );
  OAI22_X1 u2_u13_u3_U7 (.B2( u2_u13_u3_n147 ) , .A2( u2_u13_u3_n148 ) , .ZN( u2_u13_u3_n160 ) , .B1( u2_u13_u3_n165 ) , .A1( u2_u13_u3_n168 ) );
  NAND2_X1 u2_u13_u3_U70 (.A1( u2_u13_u3_n102 ) , .A2( u2_u13_u3_n103 ) , .ZN( u2_u13_u3_n108 ) );
  NOR2_X1 u2_u13_u3_U71 (.A2( u2_u13_X_19 ) , .A1( u2_u13_X_20 ) , .ZN( u2_u13_u3_n99 ) );
  NOR2_X1 u2_u13_u3_U72 (.A2( u2_u13_X_21 ) , .A1( u2_u13_X_24 ) , .ZN( u2_u13_u3_n103 ) );
  NOR2_X1 u2_u13_u3_U73 (.A2( u2_u13_X_24 ) , .A1( u2_u13_u3_n171 ) , .ZN( u2_u13_u3_n97 ) );
  NOR2_X1 u2_u13_u3_U74 (.A2( u2_u13_X_23 ) , .ZN( u2_u13_u3_n141 ) , .A1( u2_u13_u3_n166 ) );
  NOR2_X1 u2_u13_u3_U75 (.A2( u2_u13_X_19 ) , .A1( u2_u13_u3_n172 ) , .ZN( u2_u13_u3_n96 ) );
  NAND2_X1 u2_u13_u3_U76 (.A1( u2_u13_X_22 ) , .A2( u2_u13_X_23 ) , .ZN( u2_u13_u3_n154 ) );
  NAND2_X1 u2_u13_u3_U77 (.A1( u2_u13_X_23 ) , .ZN( u2_u13_u3_n149 ) , .A2( u2_u13_u3_n166 ) );
  NOR2_X1 u2_u13_u3_U78 (.A2( u2_u13_X_22 ) , .A1( u2_u13_X_23 ) , .ZN( u2_u13_u3_n121 ) );
  AND2_X1 u2_u13_u3_U79 (.A1( u2_u13_X_24 ) , .ZN( u2_u13_u3_n101 ) , .A2( u2_u13_u3_n171 ) );
  AND3_X1 u2_u13_u3_U8 (.A3( u2_u13_u3_n144 ) , .A2( u2_u13_u3_n145 ) , .A1( u2_u13_u3_n146 ) , .ZN( u2_u13_u3_n147 ) );
  AND2_X1 u2_u13_u3_U80 (.A1( u2_u13_X_19 ) , .ZN( u2_u13_u3_n102 ) , .A2( u2_u13_u3_n172 ) );
  AND2_X1 u2_u13_u3_U81 (.A1( u2_u13_X_21 ) , .A2( u2_u13_X_24 ) , .ZN( u2_u13_u3_n100 ) );
  AND2_X1 u2_u13_u3_U82 (.A2( u2_u13_X_19 ) , .A1( u2_u13_X_20 ) , .ZN( u2_u13_u3_n104 ) );
  INV_X1 u2_u13_u3_U83 (.A( u2_u13_X_22 ) , .ZN( u2_u13_u3_n166 ) );
  INV_X1 u2_u13_u3_U84 (.A( u2_u13_X_21 ) , .ZN( u2_u13_u3_n171 ) );
  INV_X1 u2_u13_u3_U85 (.A( u2_u13_X_20 ) , .ZN( u2_u13_u3_n172 ) );
  NAND4_X1 u2_u13_u3_U86 (.ZN( u2_out13_26 ) , .A4( u2_u13_u3_n109 ) , .A3( u2_u13_u3_n110 ) , .A2( u2_u13_u3_n111 ) , .A1( u2_u13_u3_n173 ) );
  INV_X1 u2_u13_u3_U87 (.ZN( u2_u13_u3_n173 ) , .A( u2_u13_u3_n94 ) );
  OAI21_X1 u2_u13_u3_U88 (.ZN( u2_u13_u3_n111 ) , .B2( u2_u13_u3_n117 ) , .A( u2_u13_u3_n133 ) , .B1( u2_u13_u3_n176 ) );
  NAND4_X1 u2_u13_u3_U89 (.ZN( u2_out13_20 ) , .A4( u2_u13_u3_n122 ) , .A3( u2_u13_u3_n123 ) , .A1( u2_u13_u3_n175 ) , .A2( u2_u13_u3_n180 ) );
  INV_X1 u2_u13_u3_U9 (.A( u2_u13_u3_n143 ) , .ZN( u2_u13_u3_n168 ) );
  INV_X1 u2_u13_u3_U90 (.A( u2_u13_u3_n112 ) , .ZN( u2_u13_u3_n175 ) );
  INV_X1 u2_u13_u3_U91 (.A( u2_u13_u3_n126 ) , .ZN( u2_u13_u3_n180 ) );
  NAND4_X1 u2_u13_u3_U92 (.ZN( u2_out13_1 ) , .A4( u2_u13_u3_n161 ) , .A3( u2_u13_u3_n162 ) , .A2( u2_u13_u3_n163 ) , .A1( u2_u13_u3_n185 ) );
  NAND2_X1 u2_u13_u3_U93 (.ZN( u2_u13_u3_n163 ) , .A2( u2_u13_u3_n170 ) , .A1( u2_u13_u3_n176 ) );
  AOI22_X1 u2_u13_u3_U94 (.B2( u2_u13_u3_n140 ) , .B1( u2_u13_u3_n141 ) , .A2( u2_u13_u3_n142 ) , .ZN( u2_u13_u3_n162 ) , .A1( u2_u13_u3_n177 ) );
  OR4_X1 u2_u13_u3_U95 (.ZN( u2_out13_10 ) , .A4( u2_u13_u3_n136 ) , .A3( u2_u13_u3_n137 ) , .A1( u2_u13_u3_n138 ) , .A2( u2_u13_u3_n139 ) );
  OAI222_X1 u2_u13_u3_U96 (.C1( u2_u13_u3_n128 ) , .ZN( u2_u13_u3_n137 ) , .B1( u2_u13_u3_n148 ) , .A2( u2_u13_u3_n150 ) , .B2( u2_u13_u3_n154 ) , .C2( u2_u13_u3_n164 ) , .A1( u2_u13_u3_n167 ) );
  OAI221_X1 u2_u13_u3_U97 (.A( u2_u13_u3_n134 ) , .B2( u2_u13_u3_n135 ) , .ZN( u2_u13_u3_n136 ) , .C1( u2_u13_u3_n149 ) , .B1( u2_u13_u3_n151 ) , .C2( u2_u13_u3_n183 ) );
  NAND3_X1 u2_u13_u3_U98 (.A1( u2_u13_u3_n114 ) , .ZN( u2_u13_u3_n115 ) , .A2( u2_u13_u3_n145 ) , .A3( u2_u13_u3_n153 ) );
  NAND3_X1 u2_u13_u3_U99 (.ZN( u2_u13_u3_n129 ) , .A2( u2_u13_u3_n144 ) , .A1( u2_u13_u3_n153 ) , .A3( u2_u13_u3_n182 ) );
  XOR2_X1 u2_u4_U10 (.B( u2_K5_45 ) , .A( u2_R3_30 ) , .Z( u2_u4_X_45 ) );
  XOR2_X1 u2_u4_U11 (.B( u2_K5_44 ) , .A( u2_R3_29 ) , .Z( u2_u4_X_44 ) );
  XOR2_X1 u2_u4_U12 (.B( u2_K5_43 ) , .A( u2_R3_28 ) , .Z( u2_u4_X_43 ) );
  XOR2_X1 u2_u4_U7 (.B( u2_K5_48 ) , .A( u2_R3_1 ) , .Z( u2_u4_X_48 ) );
  XOR2_X1 u2_u4_U8 (.B( u2_K5_47 ) , .A( u2_R3_32 ) , .Z( u2_u4_X_47 ) );
  XOR2_X1 u2_u4_U9 (.B( u2_K5_46 ) , .A( u2_R3_31 ) , .Z( u2_u4_X_46 ) );
  AND3_X1 u2_u4_u7_U10 (.A3( u2_u4_u7_n110 ) , .A2( u2_u4_u7_n127 ) , .A1( u2_u4_u7_n132 ) , .ZN( u2_u4_u7_n92 ) );
  OAI21_X1 u2_u4_u7_U11 (.A( u2_u4_u7_n161 ) , .B1( u2_u4_u7_n168 ) , .B2( u2_u4_u7_n173 ) , .ZN( u2_u4_u7_n91 ) );
  AOI211_X1 u2_u4_u7_U12 (.A( u2_u4_u7_n117 ) , .ZN( u2_u4_u7_n118 ) , .C2( u2_u4_u7_n126 ) , .C1( u2_u4_u7_n177 ) , .B( u2_u4_u7_n180 ) );
  OAI22_X1 u2_u4_u7_U13 (.B1( u2_u4_u7_n115 ) , .ZN( u2_u4_u7_n117 ) , .A2( u2_u4_u7_n133 ) , .A1( u2_u4_u7_n137 ) , .B2( u2_u4_u7_n162 ) );
  INV_X1 u2_u4_u7_U14 (.A( u2_u4_u7_n116 ) , .ZN( u2_u4_u7_n180 ) );
  NOR3_X1 u2_u4_u7_U15 (.ZN( u2_u4_u7_n115 ) , .A3( u2_u4_u7_n145 ) , .A2( u2_u4_u7_n168 ) , .A1( u2_u4_u7_n169 ) );
  NOR3_X1 u2_u4_u7_U16 (.A2( u2_u4_u7_n134 ) , .A1( u2_u4_u7_n135 ) , .ZN( u2_u4_u7_n136 ) , .A3( u2_u4_u7_n171 ) );
  NOR2_X1 u2_u4_u7_U17 (.A1( u2_u4_u7_n130 ) , .A2( u2_u4_u7_n134 ) , .ZN( u2_u4_u7_n153 ) );
  NOR2_X1 u2_u4_u7_U18 (.ZN( u2_u4_u7_n111 ) , .A2( u2_u4_u7_n134 ) , .A1( u2_u4_u7_n169 ) );
  AOI21_X1 u2_u4_u7_U19 (.ZN( u2_u4_u7_n104 ) , .B2( u2_u4_u7_n112 ) , .B1( u2_u4_u7_n127 ) , .A( u2_u4_u7_n164 ) );
  AOI21_X1 u2_u4_u7_U20 (.ZN( u2_u4_u7_n106 ) , .B1( u2_u4_u7_n133 ) , .B2( u2_u4_u7_n146 ) , .A( u2_u4_u7_n162 ) );
  AOI21_X1 u2_u4_u7_U21 (.A( u2_u4_u7_n101 ) , .ZN( u2_u4_u7_n107 ) , .B2( u2_u4_u7_n128 ) , .B1( u2_u4_u7_n175 ) );
  INV_X1 u2_u4_u7_U22 (.A( u2_u4_u7_n101 ) , .ZN( u2_u4_u7_n165 ) );
  INV_X1 u2_u4_u7_U23 (.A( u2_u4_u7_n138 ) , .ZN( u2_u4_u7_n171 ) );
  INV_X1 u2_u4_u7_U24 (.A( u2_u4_u7_n131 ) , .ZN( u2_u4_u7_n177 ) );
  INV_X1 u2_u4_u7_U25 (.A( u2_u4_u7_n110 ) , .ZN( u2_u4_u7_n174 ) );
  NAND2_X1 u2_u4_u7_U26 (.A1( u2_u4_u7_n129 ) , .A2( u2_u4_u7_n132 ) , .ZN( u2_u4_u7_n149 ) );
  NAND2_X1 u2_u4_u7_U27 (.A1( u2_u4_u7_n113 ) , .A2( u2_u4_u7_n124 ) , .ZN( u2_u4_u7_n130 ) );
  INV_X1 u2_u4_u7_U28 (.A( u2_u4_u7_n128 ) , .ZN( u2_u4_u7_n168 ) );
  INV_X1 u2_u4_u7_U29 (.A( u2_u4_u7_n148 ) , .ZN( u2_u4_u7_n169 ) );
  INV_X1 u2_u4_u7_U3 (.A( u2_u4_u7_n149 ) , .ZN( u2_u4_u7_n175 ) );
  INV_X1 u2_u4_u7_U30 (.A( u2_u4_u7_n112 ) , .ZN( u2_u4_u7_n173 ) );
  INV_X1 u2_u4_u7_U31 (.A( u2_u4_u7_n127 ) , .ZN( u2_u4_u7_n179 ) );
  NOR2_X1 u2_u4_u7_U32 (.ZN( u2_u4_u7_n101 ) , .A2( u2_u4_u7_n150 ) , .A1( u2_u4_u7_n156 ) );
  AOI211_X1 u2_u4_u7_U33 (.B( u2_u4_u7_n154 ) , .A( u2_u4_u7_n155 ) , .C1( u2_u4_u7_n156 ) , .ZN( u2_u4_u7_n157 ) , .C2( u2_u4_u7_n172 ) );
  INV_X1 u2_u4_u7_U34 (.A( u2_u4_u7_n153 ) , .ZN( u2_u4_u7_n172 ) );
  AOI211_X1 u2_u4_u7_U35 (.B( u2_u4_u7_n139 ) , .A( u2_u4_u7_n140 ) , .C2( u2_u4_u7_n141 ) , .ZN( u2_u4_u7_n142 ) , .C1( u2_u4_u7_n156 ) );
  NAND4_X1 u2_u4_u7_U36 (.A3( u2_u4_u7_n127 ) , .A2( u2_u4_u7_n128 ) , .A1( u2_u4_u7_n129 ) , .ZN( u2_u4_u7_n141 ) , .A4( u2_u4_u7_n147 ) );
  AOI21_X1 u2_u4_u7_U37 (.A( u2_u4_u7_n137 ) , .B1( u2_u4_u7_n138 ) , .ZN( u2_u4_u7_n139 ) , .B2( u2_u4_u7_n146 ) );
  OAI22_X1 u2_u4_u7_U38 (.B1( u2_u4_u7_n136 ) , .ZN( u2_u4_u7_n140 ) , .A1( u2_u4_u7_n153 ) , .B2( u2_u4_u7_n162 ) , .A2( u2_u4_u7_n164 ) );
  INV_X1 u2_u4_u7_U39 (.A( u2_u4_u7_n125 ) , .ZN( u2_u4_u7_n161 ) );
  INV_X1 u2_u4_u7_U4 (.A( u2_u4_u7_n154 ) , .ZN( u2_u4_u7_n178 ) );
  AOI21_X1 u2_u4_u7_U40 (.ZN( u2_u4_u7_n123 ) , .B1( u2_u4_u7_n165 ) , .B2( u2_u4_u7_n177 ) , .A( u2_u4_u7_n97 ) );
  AOI21_X1 u2_u4_u7_U41 (.B2( u2_u4_u7_n113 ) , .B1( u2_u4_u7_n124 ) , .A( u2_u4_u7_n125 ) , .ZN( u2_u4_u7_n97 ) );
  INV_X1 u2_u4_u7_U42 (.A( u2_u4_u7_n152 ) , .ZN( u2_u4_u7_n162 ) );
  AOI22_X1 u2_u4_u7_U43 (.A2( u2_u4_u7_n114 ) , .ZN( u2_u4_u7_n119 ) , .B1( u2_u4_u7_n130 ) , .A1( u2_u4_u7_n156 ) , .B2( u2_u4_u7_n165 ) );
  NAND2_X1 u2_u4_u7_U44 (.A2( u2_u4_u7_n112 ) , .ZN( u2_u4_u7_n114 ) , .A1( u2_u4_u7_n175 ) );
  AOI22_X1 u2_u4_u7_U45 (.B2( u2_u4_u7_n149 ) , .B1( u2_u4_u7_n150 ) , .A2( u2_u4_u7_n151 ) , .A1( u2_u4_u7_n152 ) , .ZN( u2_u4_u7_n158 ) );
  NOR2_X1 u2_u4_u7_U46 (.ZN( u2_u4_u7_n137 ) , .A1( u2_u4_u7_n150 ) , .A2( u2_u4_u7_n161 ) );
  AND2_X1 u2_u4_u7_U47 (.ZN( u2_u4_u7_n145 ) , .A2( u2_u4_u7_n98 ) , .A1( u2_u4_u7_n99 ) );
  AOI21_X1 u2_u4_u7_U48 (.ZN( u2_u4_u7_n105 ) , .B2( u2_u4_u7_n110 ) , .A( u2_u4_u7_n125 ) , .B1( u2_u4_u7_n147 ) );
  NAND2_X1 u2_u4_u7_U49 (.ZN( u2_u4_u7_n146 ) , .A1( u2_u4_u7_n95 ) , .A2( u2_u4_u7_n98 ) );
  INV_X1 u2_u4_u7_U5 (.A( u2_u4_u7_n111 ) , .ZN( u2_u4_u7_n170 ) );
  NAND2_X1 u2_u4_u7_U50 (.A2( u2_u4_u7_n103 ) , .ZN( u2_u4_u7_n147 ) , .A1( u2_u4_u7_n93 ) );
  NAND2_X1 u2_u4_u7_U51 (.A1( u2_u4_u7_n103 ) , .ZN( u2_u4_u7_n127 ) , .A2( u2_u4_u7_n99 ) );
  NAND2_X1 u2_u4_u7_U52 (.A2( u2_u4_u7_n102 ) , .A1( u2_u4_u7_n103 ) , .ZN( u2_u4_u7_n133 ) );
  OR2_X1 u2_u4_u7_U53 (.ZN( u2_u4_u7_n126 ) , .A2( u2_u4_u7_n152 ) , .A1( u2_u4_u7_n156 ) );
  NAND2_X1 u2_u4_u7_U54 (.ZN( u2_u4_u7_n112 ) , .A2( u2_u4_u7_n96 ) , .A1( u2_u4_u7_n99 ) );
  NAND2_X1 u2_u4_u7_U55 (.A2( u2_u4_u7_n102 ) , .ZN( u2_u4_u7_n128 ) , .A1( u2_u4_u7_n98 ) );
  INV_X1 u2_u4_u7_U56 (.A( u2_u4_u7_n150 ) , .ZN( u2_u4_u7_n164 ) );
  AND2_X1 u2_u4_u7_U57 (.ZN( u2_u4_u7_n134 ) , .A1( u2_u4_u7_n93 ) , .A2( u2_u4_u7_n98 ) );
  NAND2_X1 u2_u4_u7_U58 (.ZN( u2_u4_u7_n110 ) , .A1( u2_u4_u7_n95 ) , .A2( u2_u4_u7_n96 ) );
  NAND2_X1 u2_u4_u7_U59 (.A2( u2_u4_u7_n102 ) , .ZN( u2_u4_u7_n124 ) , .A1( u2_u4_u7_n96 ) );
  AOI211_X1 u2_u4_u7_U6 (.ZN( u2_u4_u7_n116 ) , .A( u2_u4_u7_n155 ) , .C1( u2_u4_u7_n161 ) , .C2( u2_u4_u7_n171 ) , .B( u2_u4_u7_n94 ) );
  NAND2_X1 u2_u4_u7_U60 (.ZN( u2_u4_u7_n132 ) , .A1( u2_u4_u7_n93 ) , .A2( u2_u4_u7_n96 ) );
  NAND2_X1 u2_u4_u7_U61 (.A2( u2_u4_u7_n103 ) , .ZN( u2_u4_u7_n131 ) , .A1( u2_u4_u7_n95 ) );
  NOR2_X1 u2_u4_u7_U62 (.A2( u2_u4_X_47 ) , .ZN( u2_u4_u7_n150 ) , .A1( u2_u4_u7_n163 ) );
  NOR2_X1 u2_u4_u7_U63 (.A2( u2_u4_X_43 ) , .A1( u2_u4_X_44 ) , .ZN( u2_u4_u7_n103 ) );
  NOR2_X1 u2_u4_u7_U64 (.A2( u2_u4_X_48 ) , .A1( u2_u4_u7_n166 ) , .ZN( u2_u4_u7_n95 ) );
  NOR2_X1 u2_u4_u7_U65 (.A2( u2_u4_X_44 ) , .A1( u2_u4_u7_n167 ) , .ZN( u2_u4_u7_n98 ) );
  NOR2_X1 u2_u4_u7_U66 (.A2( u2_u4_X_45 ) , .A1( u2_u4_X_48 ) , .ZN( u2_u4_u7_n99 ) );
  NOR2_X1 u2_u4_u7_U67 (.A2( u2_u4_X_46 ) , .A1( u2_u4_X_47 ) , .ZN( u2_u4_u7_n152 ) );
  AND2_X1 u2_u4_u7_U68 (.A1( u2_u4_X_47 ) , .ZN( u2_u4_u7_n156 ) , .A2( u2_u4_u7_n163 ) );
  NAND2_X1 u2_u4_u7_U69 (.A2( u2_u4_X_46 ) , .A1( u2_u4_X_47 ) , .ZN( u2_u4_u7_n125 ) );
  OAI222_X1 u2_u4_u7_U7 (.C2( u2_u4_u7_n101 ) , .B2( u2_u4_u7_n111 ) , .A1( u2_u4_u7_n113 ) , .C1( u2_u4_u7_n146 ) , .A2( u2_u4_u7_n162 ) , .B1( u2_u4_u7_n164 ) , .ZN( u2_u4_u7_n94 ) );
  AND2_X1 u2_u4_u7_U70 (.A2( u2_u4_X_43 ) , .A1( u2_u4_X_44 ) , .ZN( u2_u4_u7_n96 ) );
  AND2_X1 u2_u4_u7_U71 (.A2( u2_u4_X_45 ) , .A1( u2_u4_X_48 ) , .ZN( u2_u4_u7_n102 ) );
  AND2_X1 u2_u4_u7_U72 (.A1( u2_u4_X_48 ) , .A2( u2_u4_u7_n166 ) , .ZN( u2_u4_u7_n93 ) );
  INV_X1 u2_u4_u7_U73 (.A( u2_u4_X_46 ) , .ZN( u2_u4_u7_n163 ) );
  AND2_X1 u2_u4_u7_U74 (.A1( u2_u4_X_44 ) , .ZN( u2_u4_u7_n100 ) , .A2( u2_u4_u7_n167 ) );
  INV_X1 u2_u4_u7_U75 (.A( u2_u4_X_45 ) , .ZN( u2_u4_u7_n166 ) );
  INV_X1 u2_u4_u7_U76 (.A( u2_u4_X_43 ) , .ZN( u2_u4_u7_n167 ) );
  NAND4_X1 u2_u4_u7_U77 (.ZN( u2_out4_5 ) , .A4( u2_u4_u7_n108 ) , .A3( u2_u4_u7_n109 ) , .A1( u2_u4_u7_n116 ) , .A2( u2_u4_u7_n123 ) );
  AOI22_X1 u2_u4_u7_U78 (.ZN( u2_u4_u7_n109 ) , .A2( u2_u4_u7_n126 ) , .B2( u2_u4_u7_n145 ) , .B1( u2_u4_u7_n156 ) , .A1( u2_u4_u7_n171 ) );
  NOR4_X1 u2_u4_u7_U79 (.A4( u2_u4_u7_n104 ) , .A3( u2_u4_u7_n105 ) , .A2( u2_u4_u7_n106 ) , .A1( u2_u4_u7_n107 ) , .ZN( u2_u4_u7_n108 ) );
  INV_X1 u2_u4_u7_U8 (.A( u2_u4_u7_n133 ) , .ZN( u2_u4_u7_n176 ) );
  NAND4_X1 u2_u4_u7_U80 (.ZN( u2_out4_27 ) , .A4( u2_u4_u7_n118 ) , .A3( u2_u4_u7_n119 ) , .A2( u2_u4_u7_n120 ) , .A1( u2_u4_u7_n121 ) );
  OAI21_X1 u2_u4_u7_U81 (.ZN( u2_u4_u7_n121 ) , .B2( u2_u4_u7_n145 ) , .A( u2_u4_u7_n150 ) , .B1( u2_u4_u7_n174 ) );
  OAI21_X1 u2_u4_u7_U82 (.ZN( u2_u4_u7_n120 ) , .A( u2_u4_u7_n161 ) , .B2( u2_u4_u7_n170 ) , .B1( u2_u4_u7_n179 ) );
  NAND4_X1 u2_u4_u7_U83 (.ZN( u2_out4_21 ) , .A4( u2_u4_u7_n157 ) , .A3( u2_u4_u7_n158 ) , .A2( u2_u4_u7_n159 ) , .A1( u2_u4_u7_n160 ) );
  OAI21_X1 u2_u4_u7_U84 (.B1( u2_u4_u7_n145 ) , .ZN( u2_u4_u7_n160 ) , .A( u2_u4_u7_n161 ) , .B2( u2_u4_u7_n177 ) );
  OAI21_X1 u2_u4_u7_U85 (.ZN( u2_u4_u7_n159 ) , .A( u2_u4_u7_n165 ) , .B2( u2_u4_u7_n171 ) , .B1( u2_u4_u7_n174 ) );
  NAND4_X1 u2_u4_u7_U86 (.ZN( u2_out4_15 ) , .A4( u2_u4_u7_n142 ) , .A3( u2_u4_u7_n143 ) , .A2( u2_u4_u7_n144 ) , .A1( u2_u4_u7_n178 ) );
  OR2_X1 u2_u4_u7_U87 (.A2( u2_u4_u7_n125 ) , .A1( u2_u4_u7_n129 ) , .ZN( u2_u4_u7_n144 ) );
  AOI22_X1 u2_u4_u7_U88 (.A2( u2_u4_u7_n126 ) , .ZN( u2_u4_u7_n143 ) , .B2( u2_u4_u7_n165 ) , .B1( u2_u4_u7_n173 ) , .A1( u2_u4_u7_n174 ) );
  NAND2_X1 u2_u4_u7_U89 (.A1( u2_u4_u7_n100 ) , .ZN( u2_u4_u7_n148 ) , .A2( u2_u4_u7_n95 ) );
  OAI221_X1 u2_u4_u7_U9 (.C1( u2_u4_u7_n101 ) , .C2( u2_u4_u7_n147 ) , .ZN( u2_u4_u7_n155 ) , .B2( u2_u4_u7_n162 ) , .A( u2_u4_u7_n91 ) , .B1( u2_u4_u7_n92 ) );
  NAND2_X1 u2_u4_u7_U90 (.A1( u2_u4_u7_n100 ) , .ZN( u2_u4_u7_n113 ) , .A2( u2_u4_u7_n93 ) );
  NAND2_X1 u2_u4_u7_U91 (.A1( u2_u4_u7_n100 ) , .ZN( u2_u4_u7_n138 ) , .A2( u2_u4_u7_n99 ) );
  NAND2_X1 u2_u4_u7_U92 (.A1( u2_u4_u7_n100 ) , .A2( u2_u4_u7_n102 ) , .ZN( u2_u4_u7_n129 ) );
  OAI211_X1 u2_u4_u7_U93 (.B( u2_u4_u7_n122 ) , .A( u2_u4_u7_n123 ) , .C2( u2_u4_u7_n124 ) , .ZN( u2_u4_u7_n154 ) , .C1( u2_u4_u7_n162 ) );
  AOI222_X1 u2_u4_u7_U94 (.ZN( u2_u4_u7_n122 ) , .C2( u2_u4_u7_n126 ) , .C1( u2_u4_u7_n145 ) , .B1( u2_u4_u7_n161 ) , .A2( u2_u4_u7_n165 ) , .B2( u2_u4_u7_n170 ) , .A1( u2_u4_u7_n176 ) );
  NAND3_X1 u2_u4_u7_U95 (.A3( u2_u4_u7_n146 ) , .A2( u2_u4_u7_n147 ) , .A1( u2_u4_u7_n148 ) , .ZN( u2_u4_u7_n151 ) );
  NAND3_X1 u2_u4_u7_U96 (.A3( u2_u4_u7_n131 ) , .A2( u2_u4_u7_n132 ) , .A1( u2_u4_u7_n133 ) , .ZN( u2_u4_u7_n135 ) );
  XOR2_X1 u2_u9_U10 (.B( u2_K10_45 ) , .A( u2_R8_30 ) , .Z( u2_u9_X_45 ) );
  XOR2_X1 u2_u9_U11 (.B( u2_K10_44 ) , .A( u2_R8_29 ) , .Z( u2_u9_X_44 ) );
  XOR2_X1 u2_u9_U12 (.B( u2_K10_43 ) , .A( u2_R8_28 ) , .Z( u2_u9_X_43 ) );
  XOR2_X1 u2_u9_U16 (.B( u2_K10_3 ) , .A( u2_R8_2 ) , .Z( u2_u9_X_3 ) );
  XOR2_X1 u2_u9_U26 (.B( u2_K10_30 ) , .A( u2_R8_21 ) , .Z( u2_u9_X_30 ) );
  XOR2_X1 u2_u9_U27 (.B( u2_K10_2 ) , .A( u2_R8_1 ) , .Z( u2_u9_X_2 ) );
  XOR2_X1 u2_u9_U28 (.B( u2_K10_29 ) , .A( u2_R8_20 ) , .Z( u2_u9_X_29 ) );
  XOR2_X1 u2_u9_U29 (.B( u2_K10_28 ) , .A( u2_R8_19 ) , .Z( u2_u9_X_28 ) );
  XOR2_X1 u2_u9_U30 (.B( u2_K10_27 ) , .A( u2_R8_18 ) , .Z( u2_u9_X_27 ) );
  XOR2_X1 u2_u9_U31 (.B( u2_K10_26 ) , .A( u2_R8_17 ) , .Z( u2_u9_X_26 ) );
  XOR2_X1 u2_u9_U32 (.B( u2_K10_25 ) , .A( u2_R8_16 ) , .Z( u2_u9_X_25 ) );
  XOR2_X1 u2_u9_U38 (.B( u2_K10_1 ) , .A( u2_R8_32 ) , .Z( u2_u9_X_1 ) );
  XOR2_X1 u2_u9_U4 (.B( u2_K10_6 ) , .A( u2_R8_5 ) , .Z( u2_u9_X_6 ) );
  XOR2_X1 u2_u9_U5 (.B( u2_K10_5 ) , .A( u2_R8_4 ) , .Z( u2_u9_X_5 ) );
  XOR2_X1 u2_u9_U6 (.B( u2_K10_4 ) , .A( u2_R8_3 ) , .Z( u2_u9_X_4 ) );
  XOR2_X1 u2_u9_U7 (.B( u2_K10_48 ) , .A( u2_R8_1 ) , .Z( u2_u9_X_48 ) );
  XOR2_X1 u2_u9_U8 (.B( u2_K10_47 ) , .A( u2_R8_32 ) , .Z( u2_u9_X_47 ) );
  XOR2_X1 u2_u9_U9 (.B( u2_K10_46 ) , .A( u2_R8_31 ) , .Z( u2_u9_X_46 ) );
  AND3_X1 u2_u9_u0_U10 (.A2( u2_u9_u0_n112 ) , .ZN( u2_u9_u0_n127 ) , .A3( u2_u9_u0_n130 ) , .A1( u2_u9_u0_n148 ) );
  NAND2_X1 u2_u9_u0_U11 (.ZN( u2_u9_u0_n113 ) , .A1( u2_u9_u0_n139 ) , .A2( u2_u9_u0_n149 ) );
  AND2_X1 u2_u9_u0_U12 (.ZN( u2_u9_u0_n107 ) , .A1( u2_u9_u0_n130 ) , .A2( u2_u9_u0_n140 ) );
  AND2_X1 u2_u9_u0_U13 (.A2( u2_u9_u0_n129 ) , .A1( u2_u9_u0_n130 ) , .ZN( u2_u9_u0_n151 ) );
  AND2_X1 u2_u9_u0_U14 (.A1( u2_u9_u0_n108 ) , .A2( u2_u9_u0_n125 ) , .ZN( u2_u9_u0_n145 ) );
  INV_X1 u2_u9_u0_U15 (.A( u2_u9_u0_n143 ) , .ZN( u2_u9_u0_n173 ) );
  NOR2_X1 u2_u9_u0_U16 (.A2( u2_u9_u0_n136 ) , .ZN( u2_u9_u0_n147 ) , .A1( u2_u9_u0_n160 ) );
  OAI221_X1 u2_u9_u0_U17 (.C1( u2_u9_u0_n112 ) , .ZN( u2_u9_u0_n120 ) , .B1( u2_u9_u0_n138 ) , .B2( u2_u9_u0_n141 ) , .C2( u2_u9_u0_n147 ) , .A( u2_u9_u0_n172 ) );
  AOI211_X1 u2_u9_u0_U18 (.B( u2_u9_u0_n115 ) , .A( u2_u9_u0_n116 ) , .C2( u2_u9_u0_n117 ) , .C1( u2_u9_u0_n118 ) , .ZN( u2_u9_u0_n119 ) );
  OAI22_X1 u2_u9_u0_U19 (.B1( u2_u9_u0_n125 ) , .ZN( u2_u9_u0_n126 ) , .A1( u2_u9_u0_n138 ) , .A2( u2_u9_u0_n146 ) , .B2( u2_u9_u0_n147 ) );
  OAI22_X1 u2_u9_u0_U20 (.B1( u2_u9_u0_n131 ) , .A1( u2_u9_u0_n144 ) , .B2( u2_u9_u0_n147 ) , .A2( u2_u9_u0_n90 ) , .ZN( u2_u9_u0_n91 ) );
  AND3_X1 u2_u9_u0_U21 (.A3( u2_u9_u0_n121 ) , .A2( u2_u9_u0_n125 ) , .A1( u2_u9_u0_n148 ) , .ZN( u2_u9_u0_n90 ) );
  NOR2_X1 u2_u9_u0_U22 (.A1( u2_u9_u0_n163 ) , .A2( u2_u9_u0_n164 ) , .ZN( u2_u9_u0_n95 ) );
  INV_X1 u2_u9_u0_U23 (.A( u2_u9_u0_n136 ) , .ZN( u2_u9_u0_n161 ) );
  AOI22_X1 u2_u9_u0_U24 (.B2( u2_u9_u0_n109 ) , .A2( u2_u9_u0_n110 ) , .ZN( u2_u9_u0_n111 ) , .B1( u2_u9_u0_n118 ) , .A1( u2_u9_u0_n160 ) );
  INV_X1 u2_u9_u0_U25 (.A( u2_u9_u0_n118 ) , .ZN( u2_u9_u0_n158 ) );
  AOI21_X1 u2_u9_u0_U26 (.ZN( u2_u9_u0_n104 ) , .B1( u2_u9_u0_n107 ) , .B2( u2_u9_u0_n141 ) , .A( u2_u9_u0_n144 ) );
  AOI21_X1 u2_u9_u0_U27 (.B1( u2_u9_u0_n127 ) , .B2( u2_u9_u0_n129 ) , .A( u2_u9_u0_n138 ) , .ZN( u2_u9_u0_n96 ) );
  AOI21_X1 u2_u9_u0_U28 (.ZN( u2_u9_u0_n116 ) , .B2( u2_u9_u0_n142 ) , .A( u2_u9_u0_n144 ) , .B1( u2_u9_u0_n166 ) );
  NAND2_X1 u2_u9_u0_U29 (.A1( u2_u9_u0_n100 ) , .A2( u2_u9_u0_n103 ) , .ZN( u2_u9_u0_n125 ) );
  INV_X1 u2_u9_u0_U3 (.A( u2_u9_u0_n113 ) , .ZN( u2_u9_u0_n166 ) );
  NAND2_X1 u2_u9_u0_U30 (.A2( u2_u9_u0_n103 ) , .ZN( u2_u9_u0_n140 ) , .A1( u2_u9_u0_n94 ) );
  NAND2_X1 u2_u9_u0_U31 (.A1( u2_u9_u0_n101 ) , .A2( u2_u9_u0_n102 ) , .ZN( u2_u9_u0_n150 ) );
  INV_X1 u2_u9_u0_U32 (.A( u2_u9_u0_n138 ) , .ZN( u2_u9_u0_n160 ) );
  NAND2_X1 u2_u9_u0_U33 (.A2( u2_u9_u0_n102 ) , .A1( u2_u9_u0_n103 ) , .ZN( u2_u9_u0_n149 ) );
  NAND2_X1 u2_u9_u0_U34 (.A2( u2_u9_u0_n100 ) , .A1( u2_u9_u0_n101 ) , .ZN( u2_u9_u0_n139 ) );
  NAND2_X1 u2_u9_u0_U35 (.A2( u2_u9_u0_n100 ) , .ZN( u2_u9_u0_n131 ) , .A1( u2_u9_u0_n92 ) );
  NAND2_X1 u2_u9_u0_U36 (.ZN( u2_u9_u0_n108 ) , .A1( u2_u9_u0_n92 ) , .A2( u2_u9_u0_n94 ) );
  NAND2_X1 u2_u9_u0_U37 (.A2( u2_u9_u0_n102 ) , .ZN( u2_u9_u0_n114 ) , .A1( u2_u9_u0_n92 ) );
  NAND2_X1 u2_u9_u0_U38 (.A1( u2_u9_u0_n101 ) , .ZN( u2_u9_u0_n130 ) , .A2( u2_u9_u0_n94 ) );
  NAND2_X1 u2_u9_u0_U39 (.A2( u2_u9_u0_n101 ) , .ZN( u2_u9_u0_n121 ) , .A1( u2_u9_u0_n93 ) );
  AOI21_X1 u2_u9_u0_U4 (.B1( u2_u9_u0_n114 ) , .ZN( u2_u9_u0_n115 ) , .B2( u2_u9_u0_n129 ) , .A( u2_u9_u0_n161 ) );
  INV_X1 u2_u9_u0_U40 (.ZN( u2_u9_u0_n172 ) , .A( u2_u9_u0_n88 ) );
  OAI222_X1 u2_u9_u0_U41 (.C1( u2_u9_u0_n108 ) , .A1( u2_u9_u0_n125 ) , .B2( u2_u9_u0_n128 ) , .B1( u2_u9_u0_n144 ) , .A2( u2_u9_u0_n158 ) , .C2( u2_u9_u0_n161 ) , .ZN( u2_u9_u0_n88 ) );
  NAND2_X1 u2_u9_u0_U42 (.ZN( u2_u9_u0_n112 ) , .A2( u2_u9_u0_n92 ) , .A1( u2_u9_u0_n93 ) );
  OR3_X1 u2_u9_u0_U43 (.A3( u2_u9_u0_n152 ) , .A2( u2_u9_u0_n153 ) , .A1( u2_u9_u0_n154 ) , .ZN( u2_u9_u0_n155 ) );
  AOI21_X1 u2_u9_u0_U44 (.A( u2_u9_u0_n144 ) , .B2( u2_u9_u0_n145 ) , .B1( u2_u9_u0_n146 ) , .ZN( u2_u9_u0_n154 ) );
  AOI21_X1 u2_u9_u0_U45 (.B2( u2_u9_u0_n150 ) , .B1( u2_u9_u0_n151 ) , .ZN( u2_u9_u0_n152 ) , .A( u2_u9_u0_n158 ) );
  AOI21_X1 u2_u9_u0_U46 (.A( u2_u9_u0_n147 ) , .B2( u2_u9_u0_n148 ) , .B1( u2_u9_u0_n149 ) , .ZN( u2_u9_u0_n153 ) );
  AOI21_X1 u2_u9_u0_U47 (.B1( u2_u9_u0_n103 ) , .ZN( u2_u9_u0_n132 ) , .A( u2_u9_u0_n165 ) , .B2( u2_u9_u0_n93 ) );
  INV_X1 u2_u9_u0_U48 (.A( u2_u9_u0_n142 ) , .ZN( u2_u9_u0_n165 ) );
  INV_X1 u2_u9_u0_U49 (.ZN( u2_u9_u0_n171 ) , .A( u2_u9_u0_n99 ) );
  AOI21_X1 u2_u9_u0_U5 (.B2( u2_u9_u0_n131 ) , .ZN( u2_u9_u0_n134 ) , .B1( u2_u9_u0_n151 ) , .A( u2_u9_u0_n158 ) );
  OAI211_X1 u2_u9_u0_U50 (.C2( u2_u9_u0_n140 ) , .C1( u2_u9_u0_n161 ) , .A( u2_u9_u0_n169 ) , .B( u2_u9_u0_n98 ) , .ZN( u2_u9_u0_n99 ) );
  INV_X1 u2_u9_u0_U51 (.ZN( u2_u9_u0_n169 ) , .A( u2_u9_u0_n91 ) );
  AOI211_X1 u2_u9_u0_U52 (.C1( u2_u9_u0_n118 ) , .A( u2_u9_u0_n123 ) , .B( u2_u9_u0_n96 ) , .C2( u2_u9_u0_n97 ) , .ZN( u2_u9_u0_n98 ) );
  NOR2_X1 u2_u9_u0_U53 (.A2( u2_u9_X_2 ) , .ZN( u2_u9_u0_n103 ) , .A1( u2_u9_u0_n164 ) );
  NOR2_X1 u2_u9_u0_U54 (.A2( u2_u9_X_4 ) , .A1( u2_u9_X_5 ) , .ZN( u2_u9_u0_n118 ) );
  NOR2_X1 u2_u9_u0_U55 (.A2( u2_u9_X_1 ) , .A1( u2_u9_X_2 ) , .ZN( u2_u9_u0_n92 ) );
  NOR2_X1 u2_u9_u0_U56 (.A2( u2_u9_X_1 ) , .ZN( u2_u9_u0_n101 ) , .A1( u2_u9_u0_n163 ) );
  NOR2_X1 u2_u9_u0_U57 (.A2( u2_u9_X_3 ) , .A1( u2_u9_X_6 ) , .ZN( u2_u9_u0_n94 ) );
  NOR2_X1 u2_u9_u0_U58 (.A2( u2_u9_X_6 ) , .ZN( u2_u9_u0_n100 ) , .A1( u2_u9_u0_n162 ) );
  NAND2_X1 u2_u9_u0_U59 (.A2( u2_u9_X_4 ) , .A1( u2_u9_X_5 ) , .ZN( u2_u9_u0_n144 ) );
  NOR2_X1 u2_u9_u0_U6 (.A1( u2_u9_u0_n108 ) , .ZN( u2_u9_u0_n123 ) , .A2( u2_u9_u0_n158 ) );
  NOR2_X1 u2_u9_u0_U60 (.A2( u2_u9_X_5 ) , .ZN( u2_u9_u0_n136 ) , .A1( u2_u9_u0_n159 ) );
  NAND2_X1 u2_u9_u0_U61 (.A1( u2_u9_X_5 ) , .ZN( u2_u9_u0_n138 ) , .A2( u2_u9_u0_n159 ) );
  AND2_X1 u2_u9_u0_U62 (.A2( u2_u9_X_3 ) , .A1( u2_u9_X_6 ) , .ZN( u2_u9_u0_n102 ) );
  AND2_X1 u2_u9_u0_U63 (.A1( u2_u9_X_6 ) , .A2( u2_u9_u0_n162 ) , .ZN( u2_u9_u0_n93 ) );
  INV_X1 u2_u9_u0_U64 (.A( u2_u9_X_4 ) , .ZN( u2_u9_u0_n159 ) );
  INV_X1 u2_u9_u0_U65 (.A( u2_u9_X_1 ) , .ZN( u2_u9_u0_n164 ) );
  INV_X1 u2_u9_u0_U66 (.A( u2_u9_X_2 ) , .ZN( u2_u9_u0_n163 ) );
  INV_X1 u2_u9_u0_U67 (.A( u2_u9_X_3 ) , .ZN( u2_u9_u0_n162 ) );
  INV_X1 u2_u9_u0_U68 (.A( u2_u9_u0_n126 ) , .ZN( u2_u9_u0_n168 ) );
  AOI211_X1 u2_u9_u0_U69 (.B( u2_u9_u0_n133 ) , .A( u2_u9_u0_n134 ) , .C2( u2_u9_u0_n135 ) , .C1( u2_u9_u0_n136 ) , .ZN( u2_u9_u0_n137 ) );
  OAI21_X1 u2_u9_u0_U7 (.B1( u2_u9_u0_n150 ) , .B2( u2_u9_u0_n158 ) , .A( u2_u9_u0_n172 ) , .ZN( u2_u9_u0_n89 ) );
  OR4_X1 u2_u9_u0_U70 (.ZN( u2_out9_17 ) , .A4( u2_u9_u0_n122 ) , .A2( u2_u9_u0_n123 ) , .A1( u2_u9_u0_n124 ) , .A3( u2_u9_u0_n170 ) );
  AOI21_X1 u2_u9_u0_U71 (.B2( u2_u9_u0_n107 ) , .ZN( u2_u9_u0_n124 ) , .B1( u2_u9_u0_n128 ) , .A( u2_u9_u0_n161 ) );
  INV_X1 u2_u9_u0_U72 (.A( u2_u9_u0_n111 ) , .ZN( u2_u9_u0_n170 ) );
  OR4_X1 u2_u9_u0_U73 (.ZN( u2_out9_31 ) , .A4( u2_u9_u0_n155 ) , .A2( u2_u9_u0_n156 ) , .A1( u2_u9_u0_n157 ) , .A3( u2_u9_u0_n173 ) );
  AOI21_X1 u2_u9_u0_U74 (.A( u2_u9_u0_n138 ) , .B2( u2_u9_u0_n139 ) , .B1( u2_u9_u0_n140 ) , .ZN( u2_u9_u0_n157 ) );
  AOI21_X1 u2_u9_u0_U75 (.B2( u2_u9_u0_n141 ) , .B1( u2_u9_u0_n142 ) , .ZN( u2_u9_u0_n156 ) , .A( u2_u9_u0_n161 ) );
  INV_X1 u2_u9_u0_U76 (.ZN( u2_u9_u0_n174 ) , .A( u2_u9_u0_n89 ) );
  AOI211_X1 u2_u9_u0_U77 (.B( u2_u9_u0_n104 ) , .A( u2_u9_u0_n105 ) , .ZN( u2_u9_u0_n106 ) , .C2( u2_u9_u0_n113 ) , .C1( u2_u9_u0_n160 ) );
  OAI221_X1 u2_u9_u0_U78 (.C1( u2_u9_u0_n121 ) , .ZN( u2_u9_u0_n122 ) , .B2( u2_u9_u0_n127 ) , .A( u2_u9_u0_n143 ) , .B1( u2_u9_u0_n144 ) , .C2( u2_u9_u0_n147 ) );
  NOR2_X1 u2_u9_u0_U79 (.A1( u2_u9_u0_n120 ) , .ZN( u2_u9_u0_n143 ) , .A2( u2_u9_u0_n167 ) );
  AND2_X1 u2_u9_u0_U8 (.A1( u2_u9_u0_n114 ) , .A2( u2_u9_u0_n121 ) , .ZN( u2_u9_u0_n146 ) );
  AOI21_X1 u2_u9_u0_U80 (.B1( u2_u9_u0_n132 ) , .ZN( u2_u9_u0_n133 ) , .A( u2_u9_u0_n144 ) , .B2( u2_u9_u0_n166 ) );
  OAI22_X1 u2_u9_u0_U81 (.ZN( u2_u9_u0_n105 ) , .A2( u2_u9_u0_n132 ) , .B1( u2_u9_u0_n146 ) , .A1( u2_u9_u0_n147 ) , .B2( u2_u9_u0_n161 ) );
  NAND2_X1 u2_u9_u0_U82 (.ZN( u2_u9_u0_n110 ) , .A2( u2_u9_u0_n132 ) , .A1( u2_u9_u0_n145 ) );
  INV_X1 u2_u9_u0_U83 (.A( u2_u9_u0_n119 ) , .ZN( u2_u9_u0_n167 ) );
  NAND2_X1 u2_u9_u0_U84 (.ZN( u2_u9_u0_n148 ) , .A1( u2_u9_u0_n93 ) , .A2( u2_u9_u0_n95 ) );
  NAND2_X1 u2_u9_u0_U85 (.A1( u2_u9_u0_n100 ) , .ZN( u2_u9_u0_n129 ) , .A2( u2_u9_u0_n95 ) );
  NAND2_X1 u2_u9_u0_U86 (.A1( u2_u9_u0_n102 ) , .ZN( u2_u9_u0_n128 ) , .A2( u2_u9_u0_n95 ) );
  NAND2_X1 u2_u9_u0_U87 (.ZN( u2_u9_u0_n142 ) , .A1( u2_u9_u0_n94 ) , .A2( u2_u9_u0_n95 ) );
  NAND3_X1 u2_u9_u0_U88 (.ZN( u2_out9_23 ) , .A3( u2_u9_u0_n137 ) , .A1( u2_u9_u0_n168 ) , .A2( u2_u9_u0_n171 ) );
  NAND3_X1 u2_u9_u0_U89 (.A3( u2_u9_u0_n127 ) , .A2( u2_u9_u0_n128 ) , .ZN( u2_u9_u0_n135 ) , .A1( u2_u9_u0_n150 ) );
  AND2_X1 u2_u9_u0_U9 (.A1( u2_u9_u0_n131 ) , .ZN( u2_u9_u0_n141 ) , .A2( u2_u9_u0_n150 ) );
  NAND3_X1 u2_u9_u0_U90 (.ZN( u2_u9_u0_n117 ) , .A3( u2_u9_u0_n132 ) , .A2( u2_u9_u0_n139 ) , .A1( u2_u9_u0_n148 ) );
  NAND3_X1 u2_u9_u0_U91 (.ZN( u2_u9_u0_n109 ) , .A2( u2_u9_u0_n114 ) , .A3( u2_u9_u0_n140 ) , .A1( u2_u9_u0_n149 ) );
  NAND3_X1 u2_u9_u0_U92 (.ZN( u2_out9_9 ) , .A3( u2_u9_u0_n106 ) , .A2( u2_u9_u0_n171 ) , .A1( u2_u9_u0_n174 ) );
  NAND3_X1 u2_u9_u0_U93 (.A2( u2_u9_u0_n128 ) , .A1( u2_u9_u0_n132 ) , .A3( u2_u9_u0_n146 ) , .ZN( u2_u9_u0_n97 ) );
  OAI22_X1 u2_u9_u4_U10 (.B2( u2_u9_u4_n135 ) , .ZN( u2_u9_u4_n137 ) , .B1( u2_u9_u4_n153 ) , .A1( u2_u9_u4_n155 ) , .A2( u2_u9_u4_n171 ) );
  AND3_X1 u2_u9_u4_U11 (.A2( u2_u9_u4_n134 ) , .ZN( u2_u9_u4_n135 ) , .A3( u2_u9_u4_n145 ) , .A1( u2_u9_u4_n157 ) );
  NAND2_X1 u2_u9_u4_U12 (.ZN( u2_u9_u4_n132 ) , .A2( u2_u9_u4_n170 ) , .A1( u2_u9_u4_n173 ) );
  AOI21_X1 u2_u9_u4_U13 (.B2( u2_u9_u4_n160 ) , .B1( u2_u9_u4_n161 ) , .ZN( u2_u9_u4_n162 ) , .A( u2_u9_u4_n170 ) );
  AOI21_X1 u2_u9_u4_U14 (.ZN( u2_u9_u4_n107 ) , .B2( u2_u9_u4_n143 ) , .A( u2_u9_u4_n174 ) , .B1( u2_u9_u4_n184 ) );
  AOI21_X1 u2_u9_u4_U15 (.B2( u2_u9_u4_n158 ) , .B1( u2_u9_u4_n159 ) , .ZN( u2_u9_u4_n163 ) , .A( u2_u9_u4_n174 ) );
  AOI21_X1 u2_u9_u4_U16 (.A( u2_u9_u4_n153 ) , .B2( u2_u9_u4_n154 ) , .B1( u2_u9_u4_n155 ) , .ZN( u2_u9_u4_n165 ) );
  AOI21_X1 u2_u9_u4_U17 (.A( u2_u9_u4_n156 ) , .B2( u2_u9_u4_n157 ) , .ZN( u2_u9_u4_n164 ) , .B1( u2_u9_u4_n184 ) );
  INV_X1 u2_u9_u4_U18 (.A( u2_u9_u4_n138 ) , .ZN( u2_u9_u4_n170 ) );
  AND2_X1 u2_u9_u4_U19 (.A2( u2_u9_u4_n120 ) , .ZN( u2_u9_u4_n155 ) , .A1( u2_u9_u4_n160 ) );
  INV_X1 u2_u9_u4_U20 (.A( u2_u9_u4_n156 ) , .ZN( u2_u9_u4_n175 ) );
  NAND2_X1 u2_u9_u4_U21 (.A2( u2_u9_u4_n118 ) , .ZN( u2_u9_u4_n131 ) , .A1( u2_u9_u4_n147 ) );
  NAND2_X1 u2_u9_u4_U22 (.A1( u2_u9_u4_n119 ) , .A2( u2_u9_u4_n120 ) , .ZN( u2_u9_u4_n130 ) );
  NAND2_X1 u2_u9_u4_U23 (.ZN( u2_u9_u4_n117 ) , .A2( u2_u9_u4_n118 ) , .A1( u2_u9_u4_n148 ) );
  NAND2_X1 u2_u9_u4_U24 (.ZN( u2_u9_u4_n129 ) , .A1( u2_u9_u4_n134 ) , .A2( u2_u9_u4_n148 ) );
  AND3_X1 u2_u9_u4_U25 (.A1( u2_u9_u4_n119 ) , .A2( u2_u9_u4_n143 ) , .A3( u2_u9_u4_n154 ) , .ZN( u2_u9_u4_n161 ) );
  AND2_X1 u2_u9_u4_U26 (.A1( u2_u9_u4_n145 ) , .A2( u2_u9_u4_n147 ) , .ZN( u2_u9_u4_n159 ) );
  OR3_X1 u2_u9_u4_U27 (.A3( u2_u9_u4_n114 ) , .A2( u2_u9_u4_n115 ) , .A1( u2_u9_u4_n116 ) , .ZN( u2_u9_u4_n136 ) );
  AOI21_X1 u2_u9_u4_U28 (.A( u2_u9_u4_n113 ) , .ZN( u2_u9_u4_n116 ) , .B2( u2_u9_u4_n173 ) , .B1( u2_u9_u4_n174 ) );
  AOI21_X1 u2_u9_u4_U29 (.ZN( u2_u9_u4_n115 ) , .B2( u2_u9_u4_n145 ) , .B1( u2_u9_u4_n146 ) , .A( u2_u9_u4_n156 ) );
  NOR2_X1 u2_u9_u4_U3 (.ZN( u2_u9_u4_n121 ) , .A1( u2_u9_u4_n181 ) , .A2( u2_u9_u4_n182 ) );
  OAI22_X1 u2_u9_u4_U30 (.ZN( u2_u9_u4_n114 ) , .A2( u2_u9_u4_n121 ) , .B1( u2_u9_u4_n160 ) , .B2( u2_u9_u4_n170 ) , .A1( u2_u9_u4_n171 ) );
  INV_X1 u2_u9_u4_U31 (.A( u2_u9_u4_n158 ) , .ZN( u2_u9_u4_n182 ) );
  INV_X1 u2_u9_u4_U32 (.ZN( u2_u9_u4_n181 ) , .A( u2_u9_u4_n96 ) );
  INV_X1 u2_u9_u4_U33 (.A( u2_u9_u4_n144 ) , .ZN( u2_u9_u4_n179 ) );
  INV_X1 u2_u9_u4_U34 (.A( u2_u9_u4_n157 ) , .ZN( u2_u9_u4_n178 ) );
  NAND2_X1 u2_u9_u4_U35 (.A2( u2_u9_u4_n154 ) , .A1( u2_u9_u4_n96 ) , .ZN( u2_u9_u4_n97 ) );
  INV_X1 u2_u9_u4_U36 (.ZN( u2_u9_u4_n186 ) , .A( u2_u9_u4_n95 ) );
  OAI221_X1 u2_u9_u4_U37 (.C1( u2_u9_u4_n134 ) , .B1( u2_u9_u4_n158 ) , .B2( u2_u9_u4_n171 ) , .C2( u2_u9_u4_n173 ) , .A( u2_u9_u4_n94 ) , .ZN( u2_u9_u4_n95 ) );
  AOI222_X1 u2_u9_u4_U38 (.B2( u2_u9_u4_n132 ) , .A1( u2_u9_u4_n138 ) , .C2( u2_u9_u4_n175 ) , .A2( u2_u9_u4_n179 ) , .C1( u2_u9_u4_n181 ) , .B1( u2_u9_u4_n185 ) , .ZN( u2_u9_u4_n94 ) );
  INV_X1 u2_u9_u4_U39 (.A( u2_u9_u4_n113 ) , .ZN( u2_u9_u4_n185 ) );
  INV_X1 u2_u9_u4_U4 (.A( u2_u9_u4_n117 ) , .ZN( u2_u9_u4_n184 ) );
  INV_X1 u2_u9_u4_U40 (.A( u2_u9_u4_n143 ) , .ZN( u2_u9_u4_n183 ) );
  NOR2_X1 u2_u9_u4_U41 (.ZN( u2_u9_u4_n138 ) , .A1( u2_u9_u4_n168 ) , .A2( u2_u9_u4_n169 ) );
  NOR2_X1 u2_u9_u4_U42 (.A1( u2_u9_u4_n150 ) , .A2( u2_u9_u4_n152 ) , .ZN( u2_u9_u4_n153 ) );
  NOR2_X1 u2_u9_u4_U43 (.A2( u2_u9_u4_n128 ) , .A1( u2_u9_u4_n138 ) , .ZN( u2_u9_u4_n156 ) );
  AOI22_X1 u2_u9_u4_U44 (.B2( u2_u9_u4_n122 ) , .A1( u2_u9_u4_n123 ) , .ZN( u2_u9_u4_n124 ) , .B1( u2_u9_u4_n128 ) , .A2( u2_u9_u4_n172 ) );
  INV_X1 u2_u9_u4_U45 (.A( u2_u9_u4_n153 ) , .ZN( u2_u9_u4_n172 ) );
  NAND2_X1 u2_u9_u4_U46 (.A2( u2_u9_u4_n120 ) , .ZN( u2_u9_u4_n123 ) , .A1( u2_u9_u4_n161 ) );
  AOI22_X1 u2_u9_u4_U47 (.B2( u2_u9_u4_n132 ) , .A2( u2_u9_u4_n133 ) , .ZN( u2_u9_u4_n140 ) , .A1( u2_u9_u4_n150 ) , .B1( u2_u9_u4_n179 ) );
  NAND2_X1 u2_u9_u4_U48 (.ZN( u2_u9_u4_n133 ) , .A2( u2_u9_u4_n146 ) , .A1( u2_u9_u4_n154 ) );
  NAND2_X1 u2_u9_u4_U49 (.A1( u2_u9_u4_n103 ) , .ZN( u2_u9_u4_n154 ) , .A2( u2_u9_u4_n98 ) );
  NOR4_X1 u2_u9_u4_U5 (.A4( u2_u9_u4_n106 ) , .A3( u2_u9_u4_n107 ) , .A2( u2_u9_u4_n108 ) , .A1( u2_u9_u4_n109 ) , .ZN( u2_u9_u4_n110 ) );
  NAND2_X1 u2_u9_u4_U50 (.A1( u2_u9_u4_n101 ) , .ZN( u2_u9_u4_n158 ) , .A2( u2_u9_u4_n99 ) );
  AOI21_X1 u2_u9_u4_U51 (.ZN( u2_u9_u4_n127 ) , .A( u2_u9_u4_n136 ) , .B2( u2_u9_u4_n150 ) , .B1( u2_u9_u4_n180 ) );
  INV_X1 u2_u9_u4_U52 (.A( u2_u9_u4_n160 ) , .ZN( u2_u9_u4_n180 ) );
  NAND2_X1 u2_u9_u4_U53 (.A2( u2_u9_u4_n104 ) , .A1( u2_u9_u4_n105 ) , .ZN( u2_u9_u4_n146 ) );
  NAND2_X1 u2_u9_u4_U54 (.A2( u2_u9_u4_n101 ) , .A1( u2_u9_u4_n102 ) , .ZN( u2_u9_u4_n160 ) );
  NAND2_X1 u2_u9_u4_U55 (.ZN( u2_u9_u4_n134 ) , .A1( u2_u9_u4_n98 ) , .A2( u2_u9_u4_n99 ) );
  NAND2_X1 u2_u9_u4_U56 (.A1( u2_u9_u4_n103 ) , .A2( u2_u9_u4_n104 ) , .ZN( u2_u9_u4_n143 ) );
  NAND2_X1 u2_u9_u4_U57 (.A2( u2_u9_u4_n105 ) , .ZN( u2_u9_u4_n145 ) , .A1( u2_u9_u4_n98 ) );
  NAND2_X1 u2_u9_u4_U58 (.A1( u2_u9_u4_n100 ) , .A2( u2_u9_u4_n105 ) , .ZN( u2_u9_u4_n120 ) );
  NAND2_X1 u2_u9_u4_U59 (.A1( u2_u9_u4_n102 ) , .A2( u2_u9_u4_n104 ) , .ZN( u2_u9_u4_n148 ) );
  AOI21_X1 u2_u9_u4_U6 (.ZN( u2_u9_u4_n106 ) , .B2( u2_u9_u4_n146 ) , .B1( u2_u9_u4_n158 ) , .A( u2_u9_u4_n170 ) );
  NAND2_X1 u2_u9_u4_U60 (.A2( u2_u9_u4_n100 ) , .A1( u2_u9_u4_n103 ) , .ZN( u2_u9_u4_n157 ) );
  INV_X1 u2_u9_u4_U61 (.A( u2_u9_u4_n150 ) , .ZN( u2_u9_u4_n173 ) );
  INV_X1 u2_u9_u4_U62 (.A( u2_u9_u4_n152 ) , .ZN( u2_u9_u4_n171 ) );
  NAND2_X1 u2_u9_u4_U63 (.A1( u2_u9_u4_n100 ) , .ZN( u2_u9_u4_n118 ) , .A2( u2_u9_u4_n99 ) );
  NAND2_X1 u2_u9_u4_U64 (.A2( u2_u9_u4_n100 ) , .A1( u2_u9_u4_n102 ) , .ZN( u2_u9_u4_n144 ) );
  NAND2_X1 u2_u9_u4_U65 (.A2( u2_u9_u4_n101 ) , .A1( u2_u9_u4_n105 ) , .ZN( u2_u9_u4_n96 ) );
  INV_X1 u2_u9_u4_U66 (.A( u2_u9_u4_n128 ) , .ZN( u2_u9_u4_n174 ) );
  NAND2_X1 u2_u9_u4_U67 (.A2( u2_u9_u4_n102 ) , .ZN( u2_u9_u4_n119 ) , .A1( u2_u9_u4_n98 ) );
  NAND2_X1 u2_u9_u4_U68 (.A2( u2_u9_u4_n101 ) , .A1( u2_u9_u4_n103 ) , .ZN( u2_u9_u4_n147 ) );
  NAND2_X1 u2_u9_u4_U69 (.A2( u2_u9_u4_n104 ) , .ZN( u2_u9_u4_n113 ) , .A1( u2_u9_u4_n99 ) );
  AOI21_X1 u2_u9_u4_U7 (.ZN( u2_u9_u4_n108 ) , .B2( u2_u9_u4_n134 ) , .B1( u2_u9_u4_n155 ) , .A( u2_u9_u4_n156 ) );
  NOR2_X1 u2_u9_u4_U70 (.A2( u2_u9_X_28 ) , .ZN( u2_u9_u4_n150 ) , .A1( u2_u9_u4_n168 ) );
  NOR2_X1 u2_u9_u4_U71 (.A2( u2_u9_X_29 ) , .ZN( u2_u9_u4_n152 ) , .A1( u2_u9_u4_n169 ) );
  NOR2_X1 u2_u9_u4_U72 (.A2( u2_u9_X_30 ) , .ZN( u2_u9_u4_n105 ) , .A1( u2_u9_u4_n176 ) );
  NOR2_X1 u2_u9_u4_U73 (.A2( u2_u9_X_26 ) , .ZN( u2_u9_u4_n100 ) , .A1( u2_u9_u4_n177 ) );
  NOR2_X1 u2_u9_u4_U74 (.A2( u2_u9_X_28 ) , .A1( u2_u9_X_29 ) , .ZN( u2_u9_u4_n128 ) );
  NOR2_X1 u2_u9_u4_U75 (.A2( u2_u9_X_27 ) , .A1( u2_u9_X_30 ) , .ZN( u2_u9_u4_n102 ) );
  NOR2_X1 u2_u9_u4_U76 (.A2( u2_u9_X_25 ) , .A1( u2_u9_X_26 ) , .ZN( u2_u9_u4_n98 ) );
  AND2_X1 u2_u9_u4_U77 (.A2( u2_u9_X_25 ) , .A1( u2_u9_X_26 ) , .ZN( u2_u9_u4_n104 ) );
  AND2_X1 u2_u9_u4_U78 (.A1( u2_u9_X_30 ) , .A2( u2_u9_u4_n176 ) , .ZN( u2_u9_u4_n99 ) );
  AND2_X1 u2_u9_u4_U79 (.A1( u2_u9_X_26 ) , .ZN( u2_u9_u4_n101 ) , .A2( u2_u9_u4_n177 ) );
  AOI21_X1 u2_u9_u4_U8 (.ZN( u2_u9_u4_n109 ) , .A( u2_u9_u4_n153 ) , .B1( u2_u9_u4_n159 ) , .B2( u2_u9_u4_n184 ) );
  AND2_X1 u2_u9_u4_U80 (.A1( u2_u9_X_27 ) , .A2( u2_u9_X_30 ) , .ZN( u2_u9_u4_n103 ) );
  INV_X1 u2_u9_u4_U81 (.A( u2_u9_X_28 ) , .ZN( u2_u9_u4_n169 ) );
  INV_X1 u2_u9_u4_U82 (.A( u2_u9_X_29 ) , .ZN( u2_u9_u4_n168 ) );
  INV_X1 u2_u9_u4_U83 (.A( u2_u9_X_25 ) , .ZN( u2_u9_u4_n177 ) );
  INV_X1 u2_u9_u4_U84 (.A( u2_u9_X_27 ) , .ZN( u2_u9_u4_n176 ) );
  NAND4_X1 u2_u9_u4_U85 (.ZN( u2_out9_25 ) , .A4( u2_u9_u4_n139 ) , .A3( u2_u9_u4_n140 ) , .A2( u2_u9_u4_n141 ) , .A1( u2_u9_u4_n142 ) );
  OAI21_X1 u2_u9_u4_U86 (.A( u2_u9_u4_n128 ) , .B2( u2_u9_u4_n129 ) , .B1( u2_u9_u4_n130 ) , .ZN( u2_u9_u4_n142 ) );
  OAI21_X1 u2_u9_u4_U87 (.B2( u2_u9_u4_n131 ) , .ZN( u2_u9_u4_n141 ) , .A( u2_u9_u4_n175 ) , .B1( u2_u9_u4_n183 ) );
  NAND4_X1 u2_u9_u4_U88 (.ZN( u2_out9_14 ) , .A4( u2_u9_u4_n124 ) , .A3( u2_u9_u4_n125 ) , .A2( u2_u9_u4_n126 ) , .A1( u2_u9_u4_n127 ) );
  AOI22_X1 u2_u9_u4_U89 (.B2( u2_u9_u4_n117 ) , .ZN( u2_u9_u4_n126 ) , .A1( u2_u9_u4_n129 ) , .B1( u2_u9_u4_n152 ) , .A2( u2_u9_u4_n175 ) );
  AOI211_X1 u2_u9_u4_U9 (.B( u2_u9_u4_n136 ) , .A( u2_u9_u4_n137 ) , .C2( u2_u9_u4_n138 ) , .ZN( u2_u9_u4_n139 ) , .C1( u2_u9_u4_n182 ) );
  AOI22_X1 u2_u9_u4_U90 (.ZN( u2_u9_u4_n125 ) , .B2( u2_u9_u4_n131 ) , .A2( u2_u9_u4_n132 ) , .B1( u2_u9_u4_n138 ) , .A1( u2_u9_u4_n178 ) );
  NAND4_X1 u2_u9_u4_U91 (.ZN( u2_out9_8 ) , .A4( u2_u9_u4_n110 ) , .A3( u2_u9_u4_n111 ) , .A2( u2_u9_u4_n112 ) , .A1( u2_u9_u4_n186 ) );
  NAND2_X1 u2_u9_u4_U92 (.ZN( u2_u9_u4_n112 ) , .A2( u2_u9_u4_n130 ) , .A1( u2_u9_u4_n150 ) );
  AOI22_X1 u2_u9_u4_U93 (.ZN( u2_u9_u4_n111 ) , .B2( u2_u9_u4_n132 ) , .A1( u2_u9_u4_n152 ) , .B1( u2_u9_u4_n178 ) , .A2( u2_u9_u4_n97 ) );
  AOI22_X1 u2_u9_u4_U94 (.B2( u2_u9_u4_n149 ) , .B1( u2_u9_u4_n150 ) , .A2( u2_u9_u4_n151 ) , .A1( u2_u9_u4_n152 ) , .ZN( u2_u9_u4_n167 ) );
  NOR4_X1 u2_u9_u4_U95 (.A4( u2_u9_u4_n162 ) , .A3( u2_u9_u4_n163 ) , .A2( u2_u9_u4_n164 ) , .A1( u2_u9_u4_n165 ) , .ZN( u2_u9_u4_n166 ) );
  NAND3_X1 u2_u9_u4_U96 (.ZN( u2_out9_3 ) , .A3( u2_u9_u4_n166 ) , .A1( u2_u9_u4_n167 ) , .A2( u2_u9_u4_n186 ) );
  NAND3_X1 u2_u9_u4_U97 (.A3( u2_u9_u4_n146 ) , .A2( u2_u9_u4_n147 ) , .A1( u2_u9_u4_n148 ) , .ZN( u2_u9_u4_n149 ) );
  NAND3_X1 u2_u9_u4_U98 (.A3( u2_u9_u4_n143 ) , .A2( u2_u9_u4_n144 ) , .A1( u2_u9_u4_n145 ) , .ZN( u2_u9_u4_n151 ) );
  NAND3_X1 u2_u9_u4_U99 (.A3( u2_u9_u4_n121 ) , .ZN( u2_u9_u4_n122 ) , .A2( u2_u9_u4_n144 ) , .A1( u2_u9_u4_n154 ) );
  AND3_X1 u2_u9_u7_U10 (.A3( u2_u9_u7_n110 ) , .A2( u2_u9_u7_n127 ) , .A1( u2_u9_u7_n132 ) , .ZN( u2_u9_u7_n92 ) );
  OAI21_X1 u2_u9_u7_U11 (.A( u2_u9_u7_n161 ) , .B1( u2_u9_u7_n168 ) , .B2( u2_u9_u7_n173 ) , .ZN( u2_u9_u7_n91 ) );
  AOI211_X1 u2_u9_u7_U12 (.A( u2_u9_u7_n117 ) , .ZN( u2_u9_u7_n118 ) , .C2( u2_u9_u7_n126 ) , .C1( u2_u9_u7_n177 ) , .B( u2_u9_u7_n180 ) );
  OAI22_X1 u2_u9_u7_U13 (.B1( u2_u9_u7_n115 ) , .ZN( u2_u9_u7_n117 ) , .A2( u2_u9_u7_n133 ) , .A1( u2_u9_u7_n137 ) , .B2( u2_u9_u7_n162 ) );
  INV_X1 u2_u9_u7_U14 (.A( u2_u9_u7_n116 ) , .ZN( u2_u9_u7_n180 ) );
  NOR3_X1 u2_u9_u7_U15 (.ZN( u2_u9_u7_n115 ) , .A3( u2_u9_u7_n145 ) , .A2( u2_u9_u7_n168 ) , .A1( u2_u9_u7_n169 ) );
  OAI211_X1 u2_u9_u7_U16 (.B( u2_u9_u7_n122 ) , .A( u2_u9_u7_n123 ) , .C2( u2_u9_u7_n124 ) , .ZN( u2_u9_u7_n154 ) , .C1( u2_u9_u7_n162 ) );
  AOI222_X1 u2_u9_u7_U17 (.ZN( u2_u9_u7_n122 ) , .C2( u2_u9_u7_n126 ) , .C1( u2_u9_u7_n145 ) , .B1( u2_u9_u7_n161 ) , .A2( u2_u9_u7_n165 ) , .B2( u2_u9_u7_n170 ) , .A1( u2_u9_u7_n176 ) );
  INV_X1 u2_u9_u7_U18 (.A( u2_u9_u7_n133 ) , .ZN( u2_u9_u7_n176 ) );
  NOR3_X1 u2_u9_u7_U19 (.A2( u2_u9_u7_n134 ) , .A1( u2_u9_u7_n135 ) , .ZN( u2_u9_u7_n136 ) , .A3( u2_u9_u7_n171 ) );
  NOR2_X1 u2_u9_u7_U20 (.A1( u2_u9_u7_n130 ) , .A2( u2_u9_u7_n134 ) , .ZN( u2_u9_u7_n153 ) );
  INV_X1 u2_u9_u7_U21 (.A( u2_u9_u7_n101 ) , .ZN( u2_u9_u7_n165 ) );
  NOR2_X1 u2_u9_u7_U22 (.ZN( u2_u9_u7_n111 ) , .A2( u2_u9_u7_n134 ) , .A1( u2_u9_u7_n169 ) );
  AOI21_X1 u2_u9_u7_U23 (.ZN( u2_u9_u7_n104 ) , .B2( u2_u9_u7_n112 ) , .B1( u2_u9_u7_n127 ) , .A( u2_u9_u7_n164 ) );
  AOI21_X1 u2_u9_u7_U24 (.ZN( u2_u9_u7_n106 ) , .B1( u2_u9_u7_n133 ) , .B2( u2_u9_u7_n146 ) , .A( u2_u9_u7_n162 ) );
  AOI21_X1 u2_u9_u7_U25 (.A( u2_u9_u7_n101 ) , .ZN( u2_u9_u7_n107 ) , .B2( u2_u9_u7_n128 ) , .B1( u2_u9_u7_n175 ) );
  INV_X1 u2_u9_u7_U26 (.A( u2_u9_u7_n138 ) , .ZN( u2_u9_u7_n171 ) );
  INV_X1 u2_u9_u7_U27 (.A( u2_u9_u7_n131 ) , .ZN( u2_u9_u7_n177 ) );
  INV_X1 u2_u9_u7_U28 (.A( u2_u9_u7_n110 ) , .ZN( u2_u9_u7_n174 ) );
  NAND2_X1 u2_u9_u7_U29 (.A1( u2_u9_u7_n129 ) , .A2( u2_u9_u7_n132 ) , .ZN( u2_u9_u7_n149 ) );
  OAI21_X1 u2_u9_u7_U3 (.ZN( u2_u9_u7_n159 ) , .A( u2_u9_u7_n165 ) , .B2( u2_u9_u7_n171 ) , .B1( u2_u9_u7_n174 ) );
  NAND2_X1 u2_u9_u7_U30 (.A1( u2_u9_u7_n113 ) , .A2( u2_u9_u7_n124 ) , .ZN( u2_u9_u7_n130 ) );
  INV_X1 u2_u9_u7_U31 (.A( u2_u9_u7_n112 ) , .ZN( u2_u9_u7_n173 ) );
  INV_X1 u2_u9_u7_U32 (.A( u2_u9_u7_n128 ) , .ZN( u2_u9_u7_n168 ) );
  INV_X1 u2_u9_u7_U33 (.A( u2_u9_u7_n148 ) , .ZN( u2_u9_u7_n169 ) );
  INV_X1 u2_u9_u7_U34 (.A( u2_u9_u7_n127 ) , .ZN( u2_u9_u7_n179 ) );
  NOR2_X1 u2_u9_u7_U35 (.ZN( u2_u9_u7_n101 ) , .A2( u2_u9_u7_n150 ) , .A1( u2_u9_u7_n156 ) );
  AOI211_X1 u2_u9_u7_U36 (.B( u2_u9_u7_n154 ) , .A( u2_u9_u7_n155 ) , .C1( u2_u9_u7_n156 ) , .ZN( u2_u9_u7_n157 ) , .C2( u2_u9_u7_n172 ) );
  INV_X1 u2_u9_u7_U37 (.A( u2_u9_u7_n153 ) , .ZN( u2_u9_u7_n172 ) );
  AOI211_X1 u2_u9_u7_U38 (.B( u2_u9_u7_n139 ) , .A( u2_u9_u7_n140 ) , .C2( u2_u9_u7_n141 ) , .ZN( u2_u9_u7_n142 ) , .C1( u2_u9_u7_n156 ) );
  NAND4_X1 u2_u9_u7_U39 (.A3( u2_u9_u7_n127 ) , .A2( u2_u9_u7_n128 ) , .A1( u2_u9_u7_n129 ) , .ZN( u2_u9_u7_n141 ) , .A4( u2_u9_u7_n147 ) );
  INV_X1 u2_u9_u7_U4 (.A( u2_u9_u7_n111 ) , .ZN( u2_u9_u7_n170 ) );
  AOI21_X1 u2_u9_u7_U40 (.A( u2_u9_u7_n137 ) , .B1( u2_u9_u7_n138 ) , .ZN( u2_u9_u7_n139 ) , .B2( u2_u9_u7_n146 ) );
  OAI22_X1 u2_u9_u7_U41 (.B1( u2_u9_u7_n136 ) , .ZN( u2_u9_u7_n140 ) , .A1( u2_u9_u7_n153 ) , .B2( u2_u9_u7_n162 ) , .A2( u2_u9_u7_n164 ) );
  AOI21_X1 u2_u9_u7_U42 (.ZN( u2_u9_u7_n123 ) , .B1( u2_u9_u7_n165 ) , .B2( u2_u9_u7_n177 ) , .A( u2_u9_u7_n97 ) );
  AOI21_X1 u2_u9_u7_U43 (.B2( u2_u9_u7_n113 ) , .B1( u2_u9_u7_n124 ) , .A( u2_u9_u7_n125 ) , .ZN( u2_u9_u7_n97 ) );
  INV_X1 u2_u9_u7_U44 (.A( u2_u9_u7_n125 ) , .ZN( u2_u9_u7_n161 ) );
  INV_X1 u2_u9_u7_U45 (.A( u2_u9_u7_n152 ) , .ZN( u2_u9_u7_n162 ) );
  AOI22_X1 u2_u9_u7_U46 (.A2( u2_u9_u7_n114 ) , .ZN( u2_u9_u7_n119 ) , .B1( u2_u9_u7_n130 ) , .A1( u2_u9_u7_n156 ) , .B2( u2_u9_u7_n165 ) );
  NAND2_X1 u2_u9_u7_U47 (.A2( u2_u9_u7_n112 ) , .ZN( u2_u9_u7_n114 ) , .A1( u2_u9_u7_n175 ) );
  AND2_X1 u2_u9_u7_U48 (.ZN( u2_u9_u7_n145 ) , .A2( u2_u9_u7_n98 ) , .A1( u2_u9_u7_n99 ) );
  NOR2_X1 u2_u9_u7_U49 (.ZN( u2_u9_u7_n137 ) , .A1( u2_u9_u7_n150 ) , .A2( u2_u9_u7_n161 ) );
  INV_X1 u2_u9_u7_U5 (.A( u2_u9_u7_n149 ) , .ZN( u2_u9_u7_n175 ) );
  AOI21_X1 u2_u9_u7_U50 (.ZN( u2_u9_u7_n105 ) , .B2( u2_u9_u7_n110 ) , .A( u2_u9_u7_n125 ) , .B1( u2_u9_u7_n147 ) );
  NAND2_X1 u2_u9_u7_U51 (.ZN( u2_u9_u7_n146 ) , .A1( u2_u9_u7_n95 ) , .A2( u2_u9_u7_n98 ) );
  NAND2_X1 u2_u9_u7_U52 (.A2( u2_u9_u7_n103 ) , .ZN( u2_u9_u7_n147 ) , .A1( u2_u9_u7_n93 ) );
  NAND2_X1 u2_u9_u7_U53 (.A1( u2_u9_u7_n103 ) , .ZN( u2_u9_u7_n127 ) , .A2( u2_u9_u7_n99 ) );
  OR2_X1 u2_u9_u7_U54 (.ZN( u2_u9_u7_n126 ) , .A2( u2_u9_u7_n152 ) , .A1( u2_u9_u7_n156 ) );
  NAND2_X1 u2_u9_u7_U55 (.A2( u2_u9_u7_n102 ) , .A1( u2_u9_u7_n103 ) , .ZN( u2_u9_u7_n133 ) );
  NAND2_X1 u2_u9_u7_U56 (.ZN( u2_u9_u7_n112 ) , .A2( u2_u9_u7_n96 ) , .A1( u2_u9_u7_n99 ) );
  NAND2_X1 u2_u9_u7_U57 (.A2( u2_u9_u7_n102 ) , .ZN( u2_u9_u7_n128 ) , .A1( u2_u9_u7_n98 ) );
  NAND2_X1 u2_u9_u7_U58 (.A1( u2_u9_u7_n100 ) , .ZN( u2_u9_u7_n113 ) , .A2( u2_u9_u7_n93 ) );
  NAND2_X1 u2_u9_u7_U59 (.A2( u2_u9_u7_n102 ) , .ZN( u2_u9_u7_n124 ) , .A1( u2_u9_u7_n96 ) );
  INV_X1 u2_u9_u7_U6 (.A( u2_u9_u7_n154 ) , .ZN( u2_u9_u7_n178 ) );
  NAND2_X1 u2_u9_u7_U60 (.ZN( u2_u9_u7_n110 ) , .A1( u2_u9_u7_n95 ) , .A2( u2_u9_u7_n96 ) );
  INV_X1 u2_u9_u7_U61 (.A( u2_u9_u7_n150 ) , .ZN( u2_u9_u7_n164 ) );
  AND2_X1 u2_u9_u7_U62 (.ZN( u2_u9_u7_n134 ) , .A1( u2_u9_u7_n93 ) , .A2( u2_u9_u7_n98 ) );
  NAND2_X1 u2_u9_u7_U63 (.A1( u2_u9_u7_n100 ) , .A2( u2_u9_u7_n102 ) , .ZN( u2_u9_u7_n129 ) );
  NAND2_X1 u2_u9_u7_U64 (.A2( u2_u9_u7_n103 ) , .ZN( u2_u9_u7_n131 ) , .A1( u2_u9_u7_n95 ) );
  NAND2_X1 u2_u9_u7_U65 (.A1( u2_u9_u7_n100 ) , .ZN( u2_u9_u7_n138 ) , .A2( u2_u9_u7_n99 ) );
  NAND2_X1 u2_u9_u7_U66 (.ZN( u2_u9_u7_n132 ) , .A1( u2_u9_u7_n93 ) , .A2( u2_u9_u7_n96 ) );
  NAND2_X1 u2_u9_u7_U67 (.A1( u2_u9_u7_n100 ) , .ZN( u2_u9_u7_n148 ) , .A2( u2_u9_u7_n95 ) );
  NOR2_X1 u2_u9_u7_U68 (.A2( u2_u9_X_47 ) , .ZN( u2_u9_u7_n150 ) , .A1( u2_u9_u7_n163 ) );
  NOR2_X1 u2_u9_u7_U69 (.A2( u2_u9_X_43 ) , .A1( u2_u9_X_44 ) , .ZN( u2_u9_u7_n103 ) );
  AOI211_X1 u2_u9_u7_U7 (.ZN( u2_u9_u7_n116 ) , .A( u2_u9_u7_n155 ) , .C1( u2_u9_u7_n161 ) , .C2( u2_u9_u7_n171 ) , .B( u2_u9_u7_n94 ) );
  NOR2_X1 u2_u9_u7_U70 (.A2( u2_u9_X_48 ) , .A1( u2_u9_u7_n166 ) , .ZN( u2_u9_u7_n95 ) );
  NOR2_X1 u2_u9_u7_U71 (.A2( u2_u9_X_45 ) , .A1( u2_u9_X_48 ) , .ZN( u2_u9_u7_n99 ) );
  NOR2_X1 u2_u9_u7_U72 (.A2( u2_u9_X_44 ) , .A1( u2_u9_u7_n167 ) , .ZN( u2_u9_u7_n98 ) );
  NOR2_X1 u2_u9_u7_U73 (.A2( u2_u9_X_46 ) , .A1( u2_u9_X_47 ) , .ZN( u2_u9_u7_n152 ) );
  AND2_X1 u2_u9_u7_U74 (.A1( u2_u9_X_47 ) , .ZN( u2_u9_u7_n156 ) , .A2( u2_u9_u7_n163 ) );
  NAND2_X1 u2_u9_u7_U75 (.A2( u2_u9_X_46 ) , .A1( u2_u9_X_47 ) , .ZN( u2_u9_u7_n125 ) );
  AND2_X1 u2_u9_u7_U76 (.A2( u2_u9_X_45 ) , .A1( u2_u9_X_48 ) , .ZN( u2_u9_u7_n102 ) );
  AND2_X1 u2_u9_u7_U77 (.A2( u2_u9_X_43 ) , .A1( u2_u9_X_44 ) , .ZN( u2_u9_u7_n96 ) );
  AND2_X1 u2_u9_u7_U78 (.A1( u2_u9_X_44 ) , .ZN( u2_u9_u7_n100 ) , .A2( u2_u9_u7_n167 ) );
  AND2_X1 u2_u9_u7_U79 (.A1( u2_u9_X_48 ) , .A2( u2_u9_u7_n166 ) , .ZN( u2_u9_u7_n93 ) );
  OAI222_X1 u2_u9_u7_U8 (.C2( u2_u9_u7_n101 ) , .B2( u2_u9_u7_n111 ) , .A1( u2_u9_u7_n113 ) , .C1( u2_u9_u7_n146 ) , .A2( u2_u9_u7_n162 ) , .B1( u2_u9_u7_n164 ) , .ZN( u2_u9_u7_n94 ) );
  INV_X1 u2_u9_u7_U80 (.A( u2_u9_X_46 ) , .ZN( u2_u9_u7_n163 ) );
  INV_X1 u2_u9_u7_U81 (.A( u2_u9_X_43 ) , .ZN( u2_u9_u7_n167 ) );
  INV_X1 u2_u9_u7_U82 (.A( u2_u9_X_45 ) , .ZN( u2_u9_u7_n166 ) );
  NAND4_X1 u2_u9_u7_U83 (.ZN( u2_out9_27 ) , .A4( u2_u9_u7_n118 ) , .A3( u2_u9_u7_n119 ) , .A2( u2_u9_u7_n120 ) , .A1( u2_u9_u7_n121 ) );
  OAI21_X1 u2_u9_u7_U84 (.ZN( u2_u9_u7_n121 ) , .B2( u2_u9_u7_n145 ) , .A( u2_u9_u7_n150 ) , .B1( u2_u9_u7_n174 ) );
  OAI21_X1 u2_u9_u7_U85 (.ZN( u2_u9_u7_n120 ) , .A( u2_u9_u7_n161 ) , .B2( u2_u9_u7_n170 ) , .B1( u2_u9_u7_n179 ) );
  NAND4_X1 u2_u9_u7_U86 (.ZN( u2_out9_21 ) , .A4( u2_u9_u7_n157 ) , .A3( u2_u9_u7_n158 ) , .A2( u2_u9_u7_n159 ) , .A1( u2_u9_u7_n160 ) );
  OAI21_X1 u2_u9_u7_U87 (.B1( u2_u9_u7_n145 ) , .ZN( u2_u9_u7_n160 ) , .A( u2_u9_u7_n161 ) , .B2( u2_u9_u7_n177 ) );
  AOI22_X1 u2_u9_u7_U88 (.B2( u2_u9_u7_n149 ) , .B1( u2_u9_u7_n150 ) , .A2( u2_u9_u7_n151 ) , .A1( u2_u9_u7_n152 ) , .ZN( u2_u9_u7_n158 ) );
  NAND4_X1 u2_u9_u7_U89 (.ZN( u2_out9_15 ) , .A4( u2_u9_u7_n142 ) , .A3( u2_u9_u7_n143 ) , .A2( u2_u9_u7_n144 ) , .A1( u2_u9_u7_n178 ) );
  OAI221_X1 u2_u9_u7_U9 (.C1( u2_u9_u7_n101 ) , .C2( u2_u9_u7_n147 ) , .ZN( u2_u9_u7_n155 ) , .B2( u2_u9_u7_n162 ) , .A( u2_u9_u7_n91 ) , .B1( u2_u9_u7_n92 ) );
  OR2_X1 u2_u9_u7_U90 (.A2( u2_u9_u7_n125 ) , .A1( u2_u9_u7_n129 ) , .ZN( u2_u9_u7_n144 ) );
  AOI22_X1 u2_u9_u7_U91 (.A2( u2_u9_u7_n126 ) , .ZN( u2_u9_u7_n143 ) , .B2( u2_u9_u7_n165 ) , .B1( u2_u9_u7_n173 ) , .A1( u2_u9_u7_n174 ) );
  NAND4_X1 u2_u9_u7_U92 (.ZN( u2_out9_5 ) , .A4( u2_u9_u7_n108 ) , .A3( u2_u9_u7_n109 ) , .A1( u2_u9_u7_n116 ) , .A2( u2_u9_u7_n123 ) );
  AOI22_X1 u2_u9_u7_U93 (.ZN( u2_u9_u7_n109 ) , .A2( u2_u9_u7_n126 ) , .B2( u2_u9_u7_n145 ) , .B1( u2_u9_u7_n156 ) , .A1( u2_u9_u7_n171 ) );
  NOR4_X1 u2_u9_u7_U94 (.A4( u2_u9_u7_n104 ) , .A3( u2_u9_u7_n105 ) , .A2( u2_u9_u7_n106 ) , .A1( u2_u9_u7_n107 ) , .ZN( u2_u9_u7_n108 ) );
  NAND3_X1 u2_u9_u7_U95 (.A3( u2_u9_u7_n146 ) , .A2( u2_u9_u7_n147 ) , .A1( u2_u9_u7_n148 ) , .ZN( u2_u9_u7_n151 ) );
  NAND3_X1 u2_u9_u7_U96 (.A3( u2_u9_u7_n131 ) , .A2( u2_u9_u7_n132 ) , .A1( u2_u9_u7_n133 ) , .ZN( u2_u9_u7_n135 ) );
  OAI22_X1 u2_uk_U115 (.ZN( u2_K10_47 ) , .A2( u2_uk_n1594 ) , .B2( u2_uk_n1609 ) , .B1( u2_uk_n164 ) , .A1( u2_uk_n93 ) );
  INV_X1 u2_uk_U147 (.ZN( u2_K14_19 ) , .A( u2_uk_n685 ) );
  AOI22_X1 u2_uk_U148 (.B2( u2_uk_K_r12_25 ) , .A2( u2_uk_K_r12_33 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n207 ) , .ZN( u2_uk_n685 ) );
  OAI21_X1 u2_uk_U192 (.ZN( u2_K14_24 ) , .B1( u2_uk_n100 ) , .B2( u2_uk_n1782 ) , .A( u2_uk_n686 ) );
  NAND2_X1 u2_uk_U193 (.A1( u2_uk_K_r12_41 ) , .A2( u2_uk_n17 ) , .ZN( u2_uk_n686 ) );
  OAI22_X1 u2_uk_U261 (.ZN( u2_K10_48 ) , .A1( u2_uk_n148 ) , .B2( u2_uk_n1610 ) , .A2( u2_uk_n1626 ) , .B1( u2_uk_n83 ) );
  OAI22_X1 u2_uk_U321 (.ZN( u2_K5_46 ) , .B2( u2_uk_n1364 ) , .A2( u2_uk_n1401 ) , .B1( u2_uk_n146 ) , .A1( u2_uk_n92 ) );
  OAI22_X1 u2_uk_U378 (.ZN( u2_K10_28 ) , .B2( u2_uk_n1610 ) , .A2( u2_uk_n1617 ) , .B1( u2_uk_n182 ) , .A1( u2_uk_n92 ) );
  OAI21_X1 u2_uk_U384 (.ZN( u2_K10_1 ) , .B1( u2_uk_n109 ) , .B2( u2_uk_n1600 ) , .A( u2_uk_n251 ) );
  OAI22_X1 u2_uk_U489 (.ZN( u2_K10_29 ) , .B2( u2_uk_n1597 ) , .A2( u2_uk_n1625 ) , .B1( u2_uk_n202 ) , .A1( u2_uk_n92 ) );
  OAI21_X1 u2_uk_U497 (.ZN( u2_K10_2 ) , .B2( u2_uk_n1592 ) , .B1( u2_uk_n220 ) , .A( u2_uk_n286 ) );
  NAND2_X1 u2_uk_U498 (.A1( u2_uk_K_r8_41 ) , .A2( u2_uk_n230 ) , .ZN( u2_uk_n286 ) );
  INV_X1 u2_uk_U663 (.ZN( u2_K5_43 ) , .A( u2_uk_n1053 ) );
  AOI22_X1 u2_uk_U664 (.B2( u2_uk_K_r3_15 ) , .A2( u2_uk_K_r3_38 ) , .ZN( u2_uk_n1053 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n155 ) );
  OAI22_X1 u2_uk_U673 (.ZN( u2_K10_45 ) , .B2( u2_uk_n1598 ) , .A2( u2_uk_n1614 ) , .A1( u2_uk_n223 ) , .B1( u2_uk_n83 ) );
  OAI21_X1 u2_uk_U744 (.ZN( u2_K10_27 ) , .B1( u2_uk_n102 ) , .B2( u2_uk_n1602 ) , .A( u2_uk_n279 ) );
  NAND2_X1 u2_uk_U745 (.A1( u2_uk_K_r8_43 ) , .ZN( u2_uk_n279 ) , .A2( u2_uk_n94 ) );
  OAI22_X1 u2_uk_U846 (.ZN( u2_K14_22 ) , .A1( u2_uk_n162 ) , .B2( u2_uk_n1772 ) , .A2( u2_uk_n1810 ) , .B1( u2_uk_n83 ) );
  OAI22_X1 u2_uk_U847 (.ZN( u2_K10_5 ) , .B2( u2_uk_n1595 ) , .A2( u2_uk_n1612 ) , .A1( u2_uk_n231 ) , .B1( u2_uk_n83 ) );
  OAI22_X1 u2_uk_U852 (.ZN( u2_K14_23 ) , .A1( u2_uk_n163 ) , .A2( u2_uk_n1772 ) , .B2( u2_uk_n1779 ) , .B1( u2_uk_n63 ) );
  OAI22_X1 u2_uk_U871 (.ZN( u2_K10_3 ) , .A1( u2_uk_n148 ) , .B2( u2_uk_n1603 ) , .A2( u2_uk_n1623 ) , .B1( u2_uk_n63 ) );
  OAI22_X1 u2_uk_U917 (.ZN( u2_K14_20 ) , .B1( u2_uk_n141 ) , .B2( u2_uk_n1783 ) , .A2( u2_uk_n1789 ) , .A1( u2_uk_n99 ) );
  OAI21_X1 u2_uk_U995 (.ZN( u2_K5_45 ) , .A( u2_uk_n1054 ) , .B2( u2_uk_n1370 ) , .B1( u2_uk_n27 ) );
  NAND2_X1 u2_uk_U996 (.A1( u2_uk_K_r3_43 ) , .ZN( u2_uk_n1054 ) , .A2( u2_uk_n17 ) );
endmodule

